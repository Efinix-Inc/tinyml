//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2022 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = tinyml_accelerator_v2_0
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Wed Oct 26 10:04:16 2022
// ***************************************************************************************
`define IP_UUID _fc770eb8d5cc46df9bede998a24cd569
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)

`include "defines.v"

module tinyml_accelerator #(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 5,
    parameter                       ADD_MODE                        = `ADD_MODE,          //Only supported "STANDARD" / "LITE".
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,      //Only supported "STANDARD" / "LITE".
    parameter                       MULT_MODE                       = `MULT_MODE,         //Only supported "STANDARD" / "LITE".
    parameter                       FC_MODE                         = `FC_MODE,           //Only supported "STANDARD" / "LITE".
    //Convolution & Depthwise Convolution OP Parameter          
    parameter                       CONV_DEPTH_MODE                 = `CONV_DEPTH_MODE,    //Only supported "STANDARD" / "LITE".    
    parameter                       CONV_DEPTH_LITE_PARALLEL        = `CONV_DEPTH_LITE_PARALLEL,        
    parameter                       CONV_DEPTH_LITE_AW              = `CONV_DEPTH_LITE_AW,        
    parameter                       CONV_DEPTH_STD_IN_PARALLEL      = `CONV_DEPTH_STD_IN_PARALLEL,        
    parameter                       CONV_DEPTH_STD_OUT_PARALLEL     = `CONV_DEPTH_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTH_STD_OUT_CH_FIFO_A    = `CONV_DEPTH_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTH_STD_FILTER_FIFO_A    = `CONV_DEPTH_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTH_STD_CNT_DTH          = `CONV_DEPTH_STD_CNT_DTH,
    //FC OP Parameter         
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,  
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE   
)(
input                           clk,
input                           rstn,
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
input                           m_axi_clk,
input                           m_axi_rstn,
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);
`IP_MODULE_NAME(tinyml_accelerator_v2_0) #(
 .AXI_DW(AXI_DW),
 .OP_CNT(OP_CNT),
 .ADD_MODE(ADD_MODE),          //Only supported "STANDARD" / "LITE".
 .MIN_MAX_MODE(MIN_MAX_MODE),      //Only supported "STANDARD" / "LITE".
 .MULT_MODE(MULT_MODE),         //Only supported "STANDARD" / "LITE".
 .FC_MODE(FC_MODE),           //Only supported "STANDARD" / "LITE".         
 .CONV_DEPTH_MODE(CONV_DEPTH_MODE),    //Only supported "STANDARD" / "LITE".    
 .CONV_DEPTH_LITE_PARALLEL(CONV_DEPTH_LITE_PARALLEL),        
 .CONV_DEPTH_LITE_AW(CONV_DEPTH_LITE_AW),        
 .CONV_DEPTH_STD_IN_PARALLEL(CONV_DEPTH_STD_IN_PARALLEL),        
 .CONV_DEPTH_STD_OUT_PARALLEL(CONV_DEPTH_STD_OUT_PARALLEL),
 .CONV_DEPTH_STD_OUT_CH_FIFO_A(CONV_DEPTH_STD_OUT_CH_FIFO_A),
 .CONV_DEPTH_STD_FILTER_FIFO_A(CONV_DEPTH_STD_FILTER_FIFO_A),
 .CONV_DEPTH_STD_CNT_DTH(CONV_DEPTH_STD_CNT_DTH),
 .FC_MAX_IN_NODE(FC_MAX_IN_NODE),  
 .FC_MAX_OUT_NODE(FC_MAX_OUT_NODE)   
) u_tinyml_accelerator_v2_0 (
.clk(clk),
.rstn(rstn),
.cmd_valid(cmd_valid),
.cmd_function_id(cmd_function_id),
.cmd_inputs_0(cmd_inputs_0),
.cmd_inputs_1(cmd_inputs_1),
.cmd_ready(cmd_ready),
.cmd_int(cmd_int),
.rsp_valid(rsp_valid),
.rsp_outputs_0(rsp_outputs_0),
.rsp_ready(rsp_ready),
.m_axi_clk(m_axi_clk),
.m_axi_rstn(m_axi_rstn),
.m_axi_awvalid(m_axi_awvalid),
.m_axi_awaddr(m_axi_awaddr),
.m_axi_awlen(m_axi_awlen),
.m_axi_awsize(m_axi_awsize),
.m_axi_awburst(m_axi_awburst),
.m_axi_awprot(m_axi_awprot),
.m_axi_awlock(m_axi_awlock),
.m_axi_awcache(m_axi_awcache),
.m_axi_awready(m_axi_awready),
.m_axi_wdata(m_axi_wdata),
.m_axi_wstrb(m_axi_wstrb),
.m_axi_wlast(m_axi_wlast),
.m_axi_wvalid(m_axi_wvalid),
.m_axi_wready(m_axi_wready),
.m_axi_bresp(m_axi_bresp),
.m_axi_bvalid(m_axi_bvalid),
.m_axi_bready(m_axi_bready),
.m_axi_arvalid(m_axi_arvalid),
.m_axi_araddr(m_axi_araddr),
.m_axi_arlen(m_axi_arlen),
.m_axi_arsize(m_axi_arsize),
.m_axi_arburst(m_axi_arburst),
.m_axi_arprot(m_axi_arprot),
.m_axi_arlock(m_axi_arlock),
.m_axi_arcache(m_axi_arcache),
.m_axi_arready(m_axi_arready),
.m_axi_rvalid(m_axi_rvalid),
.m_axi_rdata(m_axi_rdata),
.m_axi_rlast(m_axi_rlast),
.m_axi_rresp(m_axi_rresp),
.m_axi_rready(m_axi_rready)
);
endmodule

//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
OkW1wxqwM4vhQV8ylRifsIg4EixFtA8cw6WIblte0qNggC7px2KjCibDb8pBPhD2
mRjZePC3oJsUypO0tgS5Q23sq+y3xywZzqrYGPya9vZdOSoxr6iTh5li+O7EDciT
WhVOwnb/sCU9uXFvGuHmnY+0WHQJ47g5LF6IEsFaJACybP7FyFILV5tGVrgxQ1GI
gSLMU11ue/+59ePZcht5cp/I3OE/Xaeu73x/SbXWnBV08Q0IyfzhcruIplGm1tmo
zjYc2/uBNPO0JZ8FRhNR/X9KsyVRHZ+jX7P2HxRGqfnbhICeuiJpktawZ2PdJwvL
db5gbhxwBoV0t41twbmTeA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1200 )
`pragma protect data_block
DxBZUselblb6uRSTjUQWAqVa35cNQIDnatVMOT3Nf+wxTa5i/uhSOj1Jq+65wsM7
8eGnKHENcAb6rC+81I8Uxzc2ub0zUS1Sc/53yW4ZY7hcfYUmzEXq99xAO1b+vEMU
orBplWQuyDmPASvC+BGRIAats4a1UZDQydVMWG5cE+xZ6wL5CpbZgeIMrnBUyJvY
MA38grqtmMApnmpkWuq7Li7Kh5dlXqm935uqJYvwE1jstII0Pxglfc5pTR3OBYgn
BrjIi+vrOA34ZS034GP8jEgGuLJG//gk5zGkWcAGpF3mKyM1NYF2ZjLS67mMhwZR
GBryzhSh7vb4xlebgOhuZkyxviXZhyFU8EuF6sTb8LrUAaXj7bAOlR3vphmWdcmg
CX5rhFHPMCeu1v2iAm3UJl3uObLdWgpi/ps+HOrOmgfnkvYHy8rWmWz/8o2qKf+v
+rp2ryUFHF9/4dIDStYxMOVU+33KCGLFc9+lVofvcFsCvdDcvIxAQIy+zq9790HM
t1mvui39UyokBBYhfyjdnTn6gBvVYXsCyuOSbCQAfnloEJJqa+QVq1u1bFf9t7Jn
/KLW24G9OBxAKkX6TLDAQlVJYCs5YNozoImG6CmeXuhmbOn3Ue/h956a3s3LLYdh
d0LJA+hs9XbGN4n8AsB3JzRDzoQofsC3lFbLUQEaOm0FJ7hqgLz3kMHXQ4WMpm9r
BFzFZJPFuq7L4ZHp4z5U8po+Y0s4ybSwWY5aVp9IgFXuR5JJtiKvnL5cv1Xq2/7W
ePSTsIhyb8ZDLDAhWAWvZgkaJSQlHu//7faSf++vY8/mI96hvbL5ZpdoNwyhycVH
pSpqQON5RRX2UBhZgdPmeMdpSotj4BWzf4QOm5nUoG/dU4OpOCRGSxTc1n1Cu+tb
0n3MMkdvC91rZqY0I0YMeRPUoOsaLhclpz4zOtaqRjyrXw6mY2jyLfyGwFSxstbM
V8HzlAG15e9bPS8boFkt3RKIcglnY33aR/F1KFhMEW0/MPFJaxXlCr9Z3LhFR6FC
nj400UeZz32Ts+i1UzkMPsa8jIiyy3XR44z8eijqGSyQQ5mBFt9DFsSep2Anlxf3
PocwrRBl4C8xNtjdaetT+KDQBMPZQg39Un/j+vt9VNcHdoL+n4DZciEmAh7Q9Ej7
3r6RBVEmkrmCTbTBqJnV2OTOp/4L8asD3rmf0vIYiiPxMacBhXG3SGNB4vGNXYAO
9NEnOGuOaZe+AlwIj3a4DcVztlgMXRtEMaqly0+8YnnFesI4Ll1ed1afH80MA3Pt
ofaxVJTqBpeaiOVvhVGJDycEHk+6Uw+eFKJDt6+fzyJxFEJrturj+KkqeG4rotND
M5lGGzz8gVNX4Bn8OBb86N1Tp3qAe3vBhFiDVbDxFUGcnfzC+EjuQqlY68UD/Udt
HyzLMuxP3WtzG+z4V6bMbSISOnrEN63pB4bp7rbC91hF17dZYATvA/HN7O2wKwCE
4dR+mVx0jLoSLKuRiDucGpFTjyJshmyegt2s2H1bjWDy4tx+7DRh/x9lnsodj2Ar
SoxaB10uB/GOsnIqthf3bGBYsGQ4la3dNvmWFpxe9W2NC7WFSXJizkCSckJHrTKX
`pragma protect end_protected

//pragma protect end
`include "defines.v"
`timescale 1 ns / 1 ns
module `IP_MODULE_NAME(tinyml_accelerator_v2_0)#(
    parameter                       AXI_DW                          = 128,
    parameter                       OP_CNT                          = 5,
    parameter                       ADD_MODE                        = `ADD_MODE,          
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,      
    parameter                       MULT_MODE                       = `MULT_MODE,         
    parameter                       FC_MODE                         = `FC_MODE,           
    parameter                       CONV_DEPTH_MODE                 = `CONV_DEPTH_MODE,    
    parameter                       CONV_DEPTH_LITE_PARALLEL        = `CONV_DEPTH_LITE_PARALLEL,
    parameter                       CONV_DEPTH_LITE_AW              = `CONV_DEPTH_LITE_AW,
    parameter                       CONV_DEPTH_STD_IN_PARALLEL      = `CONV_DEPTH_STD_IN_PARALLEL,
    parameter                       CONV_DEPTH_STD_OUT_PARALLEL     = `CONV_DEPTH_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTH_STD_OUT_CH_FIFO_A    = `CONV_DEPTH_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTH_STD_FILTER_FIFO_A    = `CONV_DEPTH_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTH_STD_CNT_DTH          = `CONV_DEPTH_STD_CNT_DTH,
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE
)
(
input                           clk,
input                           rstn,
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
input                           m_axi_clk,
input                           m_axi_rstn,
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SV8mbATU6655QCuR7h4KhGX7pkXHeKasGxMBOUEl9ID241n5AhgHd9K4hclyJjvX
xeL/JXgRdOvVcUYmIZQyYhaYqpzrNy1qTfBHgMSCUNptYTpgdSXcSWkRNYfwYY/q
v2N+obJCB6FQFydHIf4L1ZXcfAbHRHr32AhNSdRbyMffnRdfdFNn/pg4p+lo7ldi
FhmY2Ihj8komclKto0yL0+Yh7k7/2o1grfYDJhBI6m+FI722vDwo7HKK8LJI1XZF
/1gA1wFDkD7f5JZ5+pQtt4bPc25+HNC44nqpx9FxypteEJZn8WFpzgD2dkrHGc8q
/Ek4FzvQUpo7eIo/pGtD8A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 40336 )
`pragma protect data_block
yey4YoSUPrTibRZHmXR2/YHr4QUwUP1jdnZNOqI+PQ3FnQAOgphJlDMSdCuWn0sq
5pj6YJxFuotDLTXUvr7EQi8rDemtqlkPYzQH8S/V4etl/2kN+57Dg9+ejP6i6twY
sfAXg6NrPIt5HmnE/nJPPWZYPjpGrk2qRP/+g1Y1v0wPr+24r7EgQcL6k/A/DGbN
jCJ4NBmVkYndSuGREbN70cxQvbzih+KXbhX6VPLbOHmaw5s24Qc/Za4iqfY9E8yW
TOjqUSv5XRr42jl/HuXbYl5/lDo1tT4Jv7hRcL4i/G04p8/XROd2zCxFRmFq/3kq
rCV1eLDMAf3UMa5X/YRldDrfHWrvCuM7Ej9EhD0Lzsy+7Tl1AGj8/HZtVsAmdXdN
30wVcxX+4yfjMh52z6C46BdqLe0wUUuy1Tkt/k/vN0TZ+Pz4z6+vTw6tPuXdRlqE
5X2xav5hJCCyqryAGXZ+Yi/IQiPSGStbOHkr21Zn2Q+JMpl/TNNosAJVpPmYts5/
5F8akL4ADKJbOBEDaHF8exI2efsDTg/N3/rvF7oLYTtiYPb4FURylYytVHql6xat
8RbKJ7d7UNa3MaGuYk/yEGemG3UCZEJEFWKAyRoyy+IKy70cFnBL2xfI5VALEa5s
v2dMmVOM/wV+a2aqqXU2aiJYZEZB6QpplVrhVT035Tr+ZNZb5M6X2VuWFLuIlowN
qZPOADjCvzfR7Dk4VZcnJqP5RcVK87+DZ2rbIIAniQ0PolQzcXsdyikk8jkgLZ/C
OBDnKoPSUbtrf2BA8jqWnxWwfJ1eVYlq/FNrSvaoHwfD2SSvH/HBtml5mq4b2Zf9
c0j3h2rKl8sDwzn7Uu9MYc4Sl6Rg+pmRxUP2VG0Y4R22uh7wcDZXy1VnoLPHtMjM
yMn11ZsDrfezc73VGZ7UjCTfhKqe5HWg6Cn3MiKFFXZJFjt6UvHzrplzPO8Iok0H
nWC8CXsH6Hmt1vWc8vdA7HZbAGIBzRc7Fs1pAd71WBmI4gode+9IxgbImCTQry2w
/HRkjsZBoE/FO8dYWxWpGqUPjaz1yPtcT0fn4CEAxdvF/HjKTl3aHGFTJSx9gLe4
H+OQVB/phWg41KIhqQn5XQ+86XWlhNBMXDrYuZlAokAgpScThGTtHVEJJMwidK5p
USPPfqtaS8xzHWdS1SdrH/VZP97ljYQDjsv7ogAMVeaodO73qzq/liBSZr/R8LND
sFJ8S4e18eYmCIwy6yYyuk++i8RAwXoLhqcJnRZjirk6zWxrLwHY3CGE+EghimH7
J1cpCbZPcRQfZMrZ2IF3bcFoshSVP1P+IbRUJZET4UyC6UJr8y06BNpq6dJuN1jm
7Ac0epfv6eV1+/3IYrykdWwV1HH2uOjM+6fbZ6HpBH9QSR+S+BV2rPC80sZ5Uxzt
kD4OHtN6TR5I6ByfuNFy5sSW9/zBBGnXoZedvp/NxQj/HGltrmTcYbJ2TlXFxXi7
syAE2oWDKEMNm8o4dlwW/a/U62wgihmN9p0msHiIagPqDdxo1F9cEkVQZoIhF2de
ScNVOfuRAi5JRzdW+4gs6RPxeVhinEFnf7T4wv97Yj5WpztWJ5gR/KSVINNk2tj6
OZY/k2EDLVF1e3vSxbfn2zWVIEV0fKa57clN+ZHcNkZjpF6FZK6W9poJZ+yqfADJ
5pzqxG2VLXH9LWYcP3f6joANrmVUuJlLmbxOffqucNXkTLO8qIKWPRh8UgMliGTH
iop0rjYERgFNZlGDH4XYmOS7M9L85KbXBVu0a1PaSREkF7aFJ7/nMx5krrHKwuIG
/OgC1Ao0MmTEPRDuI1DBx4NCH5T8Okn1+/QREu5+BxaGXB2NEoAnE5m4TUhMBU7D
YUGogfMhYeYI8pnJpweN0FJ2i/P307MC3oTe3Ch0C5tMn3eT3qzM06NRS1ko7mRI
xGaAPUFy1vJ7e499X+E/Cg2iABsA9i87Qyrqs803BFCcGE0N6YNi+zxGNpae5rhZ
Vgzf6YFVQetWSYHoKnYKx1buaryNDb31WYROaqouvzd6PK1Q/8tQgWcy822PfrvP
UYlAQ1NKsvuW7IbWTUsOZloHRuByBcZAahwSJBqek38TvM+wJpmeZjBgkoaRuWBn
WVQUC60TrkEiOWyiOFAD00zcHIx32euqSoX5TH4NivDH4nKvH+WZlyLr+vKsBA+7
NSs0nCwctNYdj8avmMcysxFfv3gFUdHVrkhQCRgv/8aMWWSagtn+nZJi89GWGRC9
ZPxG4Iilyjy1TBLJeuRVx3PIPEycjSt67CcXTW0sK/C5Zp85CCOcRfrzzU9iS8Dp
WsN1nLfkIv4xrnHzp80P0X+PagO+AsFE7J/p49nWFg2ohSpKz/3zMqosrdSFeE2z
Jl2NFnwEyLECxo0AJ6d6p7ZQ3sPXaUyuy9tWSJoUKmeKlXSVE7E7YLr/GBG2Zac6
XiGCXYhfopQbS+JQCaeYRqumwyGYL+isb+fBjGMP9YfpZp5nLvKIYT1WQj2bPBUl
gPfE2lB71+nO6dxe/qcrxe0bOD2kMg4gpdesJdhSedRqeaR0FsIHMjsdnDyPokiL
uT2qQPbk2o4b1vAstnOjzvjWxUjLeuLjbgpUS9kf3ZRRGzBU5DDzRuRj4p7WuwVh
xQNF71ha4P/HLFoVzz4E2UExItoRyGcOHHR7SA3FZ3XsL5k4Ea2MZCfMEpvaa6Lc
URk1cMsKMaW8LG23bLV04P30PRNcX8LFjd3JR2YbQgCJbLJlAnjASkegrqbQU+Rp
OjpZN5aH9vkwHaYNYVCS1g+drycWVpOsbT7+jt5wuRCCZjHxLrdrUUDYZPdrE+Ss
O3yOAFOWU4wJk9Nxyk5ifVJNf7EpIUTUYJC0WI7qccdJk6m3Bhabjn/CcTvrcwjd
Ty9djm8lM3Ydfxf6PAPRTZOvYCPf6wFHwCplv8jkFWhQ6UFnd0iFUagPB4R1ts+7
gIupJLoFxNlSiXdUmK1WBSaEUoGU+cSPs8vV9+3w745NlY9yuf79JPzI8w3fijkq
PlHQu9yn+KlALr5oW2UVicrT1gwjIwlQoXkkOYpeJEVJJDbSrDDkOS94RQ2hHPyI
2M8u8bWt/lcYdAAL9IrZXUqSezxrPo7BPIQiZqFs3XWbTaIYnjmxXW94rBWWV0Tc
jkZz/HAR8sHTym+CXvUUnU3DCtDKuMKeQ1iuLFzaAl0hynWYcobvUO18gd4ODaeS
24rJLCoSCsqw0H6NuTE7La0J0HLbyG+Ak7OeADoBIREI38t56NZf5r1AnQRLveSD
8kvueyKSa7eYIt1yUYo0u8M+GWCBuLGckKjQ8EDpS1gHmbKaWwKBBTp9LYxBOxdb
sw+sbyjuXOe6r2WtetkQ5HR+XwboLpYdorjKMYj8YxNa/xSe1EkOznHZhXXHZGSs
VmH4v2QhiyDrXstpa4FOt1C5DZ17JOTt4TCd2oGIVBnWoGa0cC3UY5yRX2b388J1
ko5xcU189VV7XFYuN83lkS80qBb/XEF1+9y80M2j5R7IulFF7lZ5vWt4nCtCx3sN
HvB4UGwjowovODPOFeiSlhDpkF5dIhWzNZgaV4n2yltRTqx6140GcdADGwo9mwEQ
gzmZRMkc76Y6er2htiJ+vklUBrvFhjJaCWO9TYzW33KJKoIPRuJXak9MSN6ZufxD
MIH8SkQlGcr/1siOGl3WfRz8TONKzM1wESpOy/tdW0Cx2aLwmjKqIRC29aBAO61U
ZrLdtKQm2D6QJEt2WecOs1wdErn3bqeiu1rVowenULefDMwEriNh/9lSlAEqShx4
6QzmBDfdpbcHPWTZ2fyXUu9n6jYETtE6cf+FMCL+k4yyVl+yZzcL8tdw2BWhkiuY
5kVYAqBHrXJcyyDLFHpoanwM8SCCElEx36sax3NIQQA66WmZ4emp0hY/3E4vJuLw
5TLkYhITFtbe5BCQuESHK/OSFP+4bpLDGAi1RDfe7yfiagioxYdNNwsi4bWZol/j
4W2th2MtN2OLfMlKkk+MjYClxD0+zYL28zJu7tylLoxyhFvZItxs6sXcXVVY+c7j
PK7HUh7pu4GhbocD0UgoMSkR2kkJa4P+HEaJgk2HsiN3plgOm1+7tEkPExatgtXY
Te2vbSSNA/yWC88WgbYoe36E9haYJLH9mJLD/jBeTvjSoPjvNoDQqX0H9/ArWFHb
sENPnoSu0MJN4Pp/jMQEZv/JtWoP1vtDXNyAB3WsJvRtjt4p9O1UCthRp2PkZvt2
FS/Pm9IBgqzeNmVLB+Xe5gxZLOqz7Xa4MBNr+jwHdVmwCfstRupOWe2dKa26buo5
fSTlcyGxCFacr7KD5sfI0CuGa66C06RaePp02S/Gby6JGo7OB2la22HAx7d4yFn/
TRO9kq/yvFpfqQLl0T/2A0TL1LDsV35/xvOL1ulrvy0Kf4sYsz/tQwTh7Xuhe2q9
s/6kH6SUmq+FwydBWH9JgMJt6ePq1VnEFcqR2s3OBGvubDRbz/8gr3oNzhnDN4xw
855fSDC0zLS3ScgG9DUuiuP0w/hd4nHnOzH+xCYsoRr2A5w2ddrHBKZZohtFk51E
Wjh07s2nJhp11aIC8VeEv2TcQK4sPbdd2SAHzK3EJnK1Wwr1yYOzR+GkCWuMZNuX
uufYi8yfB7C7/NvTxuwdxwwaGYvDN3Lv/aos3cS4K4Y8ieYwkNKbtr4X8+NPuzxM
u7JxpTBPfa9XvIySVCE8PZYnmfbYv5ipB0C5EXEkKskNXj32Zr+6BCuIyKr2JYCV
Wukqm1xIEJNNn0fUnTas/YmZeb0Y53KgSx3jLvF3eEhIWNO1odzpN3xQ2OWHi0VI
qr94nK3q0ECJRwxT6gN76LGSHcyHGL+oYWxpbaa2co7sU1e11nAPnA7ptwcQvhJT
3lbzLChL5gqp7jkcnnhJ+9PTn7hZnP3aD1GyUyWGzSZDSB+6AvpB70KYioBbVahe
eD5q+olcatm4oy5uB7ZZtyih1tbp1JfinbV9aYRWSsmuddP4Gwo52aeCTyVALxY0
Q3MCpzOuZeQbMDzO5A13GU3+TzJo3ula7Rjz0cPwitSHiUPQKfyzsZO1w5ZWowku
U+GPA4PV5E+uYULvj0OnlVqzu15RiUnkE8I8WCEHq/i+Wvnn4pENA9No/hcyP0ZT
+Do5s67FxKNSSxpvgHpDQoGsQneqiQdTO43uVtg4+SDXWt/FzZ/Jku4+Nn0mBCEo
FD68A0To39Okb5C45U0MuhiRgErfFdaMX6yUfsAZbcfo4y5Tmg9+pGlPbUAZL/7I
fQPa0WehL1YvzWASej5u7YuZ8oM2QaTIoFlsk94AMhge4X9A0OX6M9+wzDOGmek2
3gzQIkQ/DzWCgXpeX/j/u3m8B95nUz6dEtI/Q2djFvb7MelhxskYRnkn8dr/pkau
NOybWjRcSNXmbZH9u9kH7T06uORKrefzx4dgPk9iTsyenmxTyqKC+v8vUP5oNoIq
tu+QuX+KYRWfSJkDcFu4BZKs7gCxhosDFI2orV5UxNriK5v1ikNRi3KvYifgVVRp
iELh/HM8KjNFO++MGVKRnAW23TBNwbSMPbkZIusD4v+qcXVY0S6OqRRMTItIpF8M
aD96HrEdAPBIStDdxEeKz3QU+XYlRX9U3LauD0nxUYLW8qnsc83UvrclN9pJRUu2
B4NevcYNvwJGgIIfVXbTcdpMQYlkMYoK+gXUvf54V9EQNSICk7h+9jeI2vW/siR+
+hkGu8jFmI4Yh1IRfMJgWipBw15x/7knbevfFMYcn6i1DQivxqzLQpvLVq1VfGFj
lFVso0zpTAdY72gRw2wRCghLZf4fQZw+YbWiUBKr8867f8LgzIGDBG+snJtqpEd/
WxAPr+I4wxWJeBXPNXhUalcYRLbpRwI25dvyaE+QaZRB6zlNPeqDtdQpe22TIbp/
85LNXAatDa7h3euEu/q0O8W09CsA42bMCO25g5XvV3rfHeQf64b/OmXgvvyjL2AD
vmHhBa43eUpvPEfn1mZAsi5/5V1M7IrCee/VnMKs0MqMO1tzvgmzsY+4672T0lAN
bBOSD6yTJvtmcep1A+7o/9bzOJ5k00pETJdBfKJ1oaqf236zvGs10qZy0WjTGHLm
zMEaWaho7SzyJPdMiy5bq5FCvWAFCNk6HqckpHUEQybhexNlfv2hdGJ+AKZ7pQx9
VfHlz+GANdMBEGKB4ECRgnP6gSx0K4FZ74Run7c9vgClmE4tLq6FGnwzFvarZkl2
c565Y22njwZU+JfQL7vDPKSYN2AF3BzTh1dSguud3zgxyVFg+f5oX62XWdM+1rJ2
inBp9qSsI09eNZLrAt3bLN4gI2UyCfn9NhdmFXfoHdvREg1u1bamqJLZ4s7XqDWI
3R/Zv/kZnCaS5Z3iMpinU8txb2hZ8KQzrxlsJp/74TZbIY1X8mS3T/yJLiHikUWb
FdBPgnZcQrpMIQ255CvXUTd9qVaz8GpcVyT9pRugxc144WyEcXqtD4NSqWIGZa9X
Y14YAuBkEfhP8OOLf6Ad7hxX5Azz/TcGhJQToUu2y/3rfrdzQMs13VTpvlXoxEUM
HwiSsfg1bzqO9Vx6O5NsnOIrEDWsT14e4AfvzCNn/CUHSaJdhmHbrA1cKz0t5aF4
B9STnob3JIO+gxPrYi+MJjXzbH1UB7XwDQTXBG3h/CQJydwqUaEgkmuynh+uzT1o
/J92EpDJGYBCb8pJjEMyOl42lQfpBIDBitZYyhJrF7hAK/3MuxAy2sQefxtdCIYW
cfXiBjTqXFGFvBVM3zetKwUz8BYJZ1/TFlLXR/eaqFW61MzvJ3TwKiAu3Mjywlzf
QTMYZX8D48VtexynflpHBrqzE/kKPfeCYmFGaaTjUL9DglyRgleUZ6p33ZCPLlRF
7K28Hy+0EGkzXhUKkOVmq6JoBxvK/drUkwi05gvafM4ReKxKtcY/+fKndC8jkm7j
lXCwjPhfKHCSd6qojrMOX6oiet3PE/gyCvvyvUnlKSPXN+us/mv9RVAW/Aimrt6S
62+A8TwaI937q50F0rohyMKB48VUr1bbER4IGFJb4FDxJPBJfvbQFizNPGNGjBaw
FtSk9V9EOnlthUocwTDK7WVQ3cPTlJMyAOJgMEbTOMtrEKyitFp/o2gUWWNIBM6x
5CqnURBCmwinYiEbAXyJSgko0GDNjb87WMgtY6Lu/UO7YzZZcdrX8dl0IUVEZV2e
+qQ0vDS+Yq8I0byn2MEO/+L6vTlOaZDaT79rLOK1IpwgmJACPt3eUT4BMb64RfId
puLn9gitM7A8G/9RkoP4USkiELfAdelI+uCMvNItINjgpjXZosSN4VLr/Ow3UdsT
1/iBIT2MpEbA1lZZ6FvVl/olaO/xac0qG8jbQxLzFWLEdkrqeoFt2gs/E+mWk9cf
7Y4dGUZq6Ut7jlXAQ9vQpUJbrXU0Uf3GcX0KVDM2kxv79bPT6aN3QuLxhc1uET1a
+ohwhwSNhadRl4jYZz97FQhGucgElGDgQUQCMB4pVToOqdCRN6cmBLfsAuOCZ//V
kn3SS3add4Fm1WQqYY6X8XgUO9yBd4rnwZCE9v+m1fZumrTM/VTbd6n2b7OFplmo
PK0HCAAE8kNlSDw3iOISEb7XjvcIi19JfMqIaUx5ZAeGRVpOZd2IOXsya5CDDZgV
WgZlc9fZO2FNx9sDMLmQLxmI3Y6U11M/LPbfD7mUFs9UANUYimrAb9XCsqSbzFLC
sW2V2s9jyGU3GvIwrsK2FqqfynQgTcMn8z4iwWHe2mspKCLNHOBdN+9O8XBCILuo
M5tvPzV4ZCKkeMDKM6HnTOzRD8OY6wXhX9Z1w/Swxcy85/96gsduoXZiyA0ieWzH
0Lkjb9MQyV6R0v4NECRLdaY7Ixt4mJPa/jVmfXKa9Wx6CA1a7qiI8ddzwMThjwHR
sBPol4H7gtvITM4eQl+dRfVa1kzLM32aPjWyqQUD40BOsSBjfDKRa5+UgEwQzgEr
TUY5z0ryPTHdH/Jx3/pQVOGcoiKQeL0VmIaxzGNp0NFBoTji50ohOlUcKhyXKShC
p45kBGC/0WMJDLPN6iv26+9JiQcuyCnkc3ZI8KA+QYU+mhW071CcVw7Np8sWpomg
GVg9GFUgHgLGIupbfnCD/vf5zr41RMe6gsBp5kJXJtdfibGPJBbKhBKu7AI50GZm
gPMlgbUhCwmMk/7k/xQQDVvNdUg5QeY9RgFzTz+9ZO5o85nPnZ0SR3cMim8ciYjl
kARGk6YglGn40FEnEojcUN4chaAvHQpJYF+gqXh2P4q/+XM3r9WYTyDW+zjXK3Gx
koNkPCIn4pQMUKHfuDfbYDX6O7UU2ulaYkK/vLORuoz+xGfSrHcewf//WhUzcywT
UzItfywp7OK8uXCq1mIrJOPp8gBVvR/rTo2B6hCvhBap5BzDNA4Z0Jlegc7/nYOv
b/bu7IbQrwit/JCrBMwCubKvdSU5x9oqOldru9sdlTn37CM9dmcl5Mf9B54VF6HQ
CICz7e2Uqi1SrRdQ81PP/tq1qFf68mcARNWH8Jh3ZPMmjXcoWhysIhZVw/8xcfDB
Fy+y/JV76P6j4EQXYATSZekVn6qRt/vzmmOgZFOXFzCSwegguOyYKVn0MkXSIRj1
oiT5RbBibMEazihwjXKEfnwH8VRXlfjxOwNpZdbYMhRovROd/LWEd4+/lPUby3u6
g0zpXlDkBsSRuOZnS3/uT2jblP+lm9gwLMM9oykFAoIQFq/pQGmAmAANq77iQOKG
/MuNcQj2dRanhagvw6s1FDeLOrk0lAPozIZdyYRRwpK6Sz3IRSQZGuAmUUEVKoAU
VuDdrV1ZWgfUE4ueKgrl/uj7w310o96PPXH8V5oCL0LSviDqqtVLxrVo8B4sgURo
ybkLW7roSyILYkcsG/uDryLn/YTtk9C1NkJwjhzN2u2hNI53bEv+JndM/V0KYjJN
LaGzEnm8WMxjtka192ItRDAYjdjDsvng1UHPnF7fgmN7HMfHV7QYOUUruZcjZ51e
2Bp4absv3D4WkUEkEykei4qHkkZl/KQ90YM5sAL0ojzEfYqqGn0kGidhLo2j4mm1
Q1jFV5vSjAn1KNPZ6cge73ZWIHQzLF69WDdQGtxoalDVmXeC5EKJfTE7FJVY8ImS
UC5wBg/U87/Im739L8jbFQuP2MDUAHHJcdAgksM9HZgr5EQOI+miF6ZNnsMNMzLL
4soreoeCAZybnubgUDYIEI05VIDYW1bbm9xO7ygBrWgFlPOAGvMnAwitf3eUctK2
vzqIsN+6WIjsZ6zE6jQ3HbXEkQBXmm3/tSU77jlTjIbrrJ1G5A5lDB3VULBGkBlL
SOFRyHUs7FUXXW1DwhW3yV8mF09B9958V3SC+IUXTKuVtOE44s8+0jHCfCSO56wQ
Oz6d+/I1jr969yXsO2XRzA99N1zvkPzracruUzdIXVMbdXr/Op9grnJCBzRj4JYU
pvlzJkKRctHCtnPLvwz3e0IjPyCeudnI6xDpwAIdEe8/+S0XgXRa6vhrB+rCtNDV
3uJvhVnT5LnTbcQQd1LvrZ287wgu7zo+AQ/pQL1kwLPKUMIa0XEHjtdaVAD4BXOJ
OTY/sOcBBUQclDc4x7KAZCekOKMPF3YVsM8Ex3yFRKMvO8jvJ1ilZlxUsxh/X0UE
qaD+DSX4PCgRFbmPMv0sgAEfUPuRff2s98JFqsKyxoXT323nUzYXoCRbXya85bXY
Gl2zPwxNUOOvuQjJ1sYUZK1DGktEqOoNXxmYs2/l9rGRaaFroDNpfdIkWT6ZVzb0
fH6cMpqEftrnKfa8rT04/IYa2uxBBYHeWyD/Vv5slqCCfuGaQwYaC/9tXhlFELs1
Kz19jVlIfCz0aNx042H0fLKYv/uxdMqfU3d9N6veZCUVnNBrUYIJLDLV1Oni+EEh
2NhApCd/83FUWtYmBRyxgw4mnmPEE+O5CmKMeav5a2t1KJgRfOKbEuBdCDRG859V
oRV3nDUIWYk4sd6bw2gyhTAWYEX6h9EGdxlwFDwQie2pt6LpYM/xAKPohlFGbP5V
UarkS6Vq6AwTDbJfcXRdgmTzM6pGCcZbf3oInHSn+5vZlMNpXsKruhe+MiPZwshl
haITcdWNQdsOiU3yojgO+3GCiMdOUuDQ2M4X1nMo/GjJoD4o/5n+sIgmuuRqnP+a
um66SVMgIt89oumSM7ZxcAfFwJ3cTz9FK+xiDyeTbe2jVK1OvzaVOAXM7ssZ6MXL
eEu+QaduG23TCQ1csA06OnIrCpV6WdAdSee8qzrMsRWx9GTWKt1r7EAvLQAiUj1j
bigqvy1EZWdFPtpOywRJvhaNMM16xVS0DpMViOdqf1G86qXaU8ErXlHQLQPYvrh/
Mf/k9dA8BqRk3lG/EnK7aD1gcVc1HZSq6cL1HSSEUgs8fmrgxfn7Pw19GTTT0wGZ
CZEvO9WGj4SXd95hkTBRaMC1GMQSkCv3U+gXTn3nCATcd9pZZYGmGT5b/B2DjXS8
0lazrCGEXFFnWR3AG0XOLITrdCg2MmRqD+0ahUK7hK2M34uYb1eLdnyd76XyMC+B
gPYyPK0edbtJhsQ13ohm3MBm616huCsJUCWmXttGosajFgwgK8+F/qZQlfqL59pU
hrMJRduj8DNb4EQvJ/CwRd2sQX6Q27O0z5hUbz1InbjdJkrTNSPC5IesZdH9baWC
62CUe8gWK0Regpm5SS7ZcvWZqt2HflTzYZBA+Dq8MOprLEGK0YtNbLfQ+hLrYuXH
jeEy8U6pn0SHQXmC2oZWWEgeQgENrCZZGoOhts3owoS/6Jyxk/AQIpbvOnrN6vuU
8iKi3coI8YQ601nXF6oOZhrdYLC9sVSfWgIEK/pG8EGWrEWtx1Z39mtBd2BWHDGa
9jG8NiaEmYXVglABeW32SRIIWdMxDYeVeKa2mJFh3Ud6rLm5VJ9WlADzL4jGfLXq
g649EYJFu58HgvX1o96KyAfiuCfkFx7qabMGUROT5Yx3G6foFb6QkEZIZNrtufzo
9JbthJQyFZcm7iWwhECkqjsowVHbxAzEJVGbxy7vv7/ATNQWkF0m4MptIYITzwpl
ZE+0s6EjjD5pun1sfIvFLd15HYSzIk7c3JpjoJjPfJC4L8KH1rqL6D0peUpC2krK
Yc0WhRXmh8gWx7ZD7HoZZcyLf2GA9gQhhccirPFjXEotvOk062RwhHFYEtoPBsaL
RTPIcXT73KCNTAdNOdZSgU5MHQjrd0/efXbtAXbS7zQAD3XCZwMZN89w1kNo8H5N
MFtoFW4uVI0RXBE8KgaQwFvfmi8tEBLMcDwz/Ojm1yrwutY5eq2v0TMGplc2rAQ/
W25tDAyg2wDuI4tXAAZj7xjxQasSJdVQo4+IhCFPf3Pk4Sm8XjtIWUDfUga7vbHL
TMfNNgpuB3gf1RhWAQ5Z2uWM1Th0yngI6vR+8XoDgr3cKT4pEHoNG6HXSCMTOebX
kOSqdtUpYuDY8Q1lPu6mH/fFnj+TsZqbjq55DcqYkNb1GTeatKlllRhCXV53ypGu
HCo+ZxxwAs5ql6E4G05Vxu2GFd4M1ghjP6P3JACfbmrG8+JIwK/y9pDahO7djzHd
Q/FC/S4zg/BBpgla7+fXJpvkd3tjsi8BYQaxB9PFzEHMlxdcyVqDE7FNVibgrNBE
KXQ5KSb4L8PW1XaoOuR49iPEUrmO0gckPNO6Vs/zHZtrZGP34dn3xW2eg7PnI85y
UHAKwM2bShoshY6Um5WZPFFaLWoElZmvboFZ8RbzmxhWUACdAztlH8sWAgB4KX2U
IzosRjMQqfymdJFAqSucGurx8KFnSqSa3lbS2Nvv4T4MsDE8/wDra3yA1LgTJoxr
gx4fQQ4UCzTCkggG1waHBC/7e9mGMaxBn2/pHpI+Pi7f4X5va/aBdRy4m1rDgMtK
rwRJ5Qoae0a3Z9UcUASGuTWnGo2hneqzbV9PaXhl4J/4rZX54N4+DIL6HnzSWoQO
+qjFTIPeXUtyH5kNm1Zi8vcfBoG9QHl4ap+YJAgTu6FBSW6OP8cip3hDIgIYrrin
KeabpqE3GXpjtJG0cGSkhJLeGaYK2MsWnH4Y+A0TPsbbfhk8qfg904rNaj58ZcWE
b1V7a6Zpre5/YX88s1z8EUHR3ko1oO6z62cry+mIlb6MH+xK/OtFfasE7X3bD79x
rvK4z+McnrAorRPO3XBQCCUrEtX+UdaQ5IROnbTkghQclPl1DmG9zRwO+ED9hRHt
2fqcYVKfP5yS2g4uge8UNyG41RbFNhDl71MpM5imDvMhR/parCsdKKmyJ5Jt1sNq
pphtmoZqgHkga+jB9l30gCSXsTemRj13dxcpc5Lsbo64EilGLkm19dOJcdIIQScZ
9F8vdYdwF/dd1YkKdd+0hap3hjqmqfDGgL6zXLne5OrPrEJL/QyeW0SXgHrAQE2w
kBAae7I7M0FzJqNW8e2ismBZIOTqeeuFgGp/Ri+TZgn7Mv9/SP5NDuqDZQ4RsF7a
g2uvqPAYoZc1PEGYLfs1d49bgxzaMLo3xbYBLikFpokUss0n2YZnvdKUb6IGf430
TLzJqDbfT4iqnlGjisdGAsCfp/2x5wWjOPFCtYsgLX3WCbtUaWeWRBTbY/hUI3Ps
6mBuNGSsrKBnglbLYbpBqoC57YuVTsoUIEk+YiqhkOPhm1U2nQE1gPk2SwsBiMUr
/a22vibvS86OdHj2WbYeVktcxmhIIVwN+SF5sV3c0OZ+FQ5t1RKVwzP9p6unhYnc
6EEQpB+uPuXkTU8SbIanK2iBSF7YbxHKlHLaNNfjOrl1SyrNIeCcGMgufzdnsfPJ
zs+pclXlRmrd6E5zTSWvPEG1TgaDBPQqfs2NxWSDMmE8eBjaeSRNNCX5YRldWKLJ
Fp0HOdhb2sj7yB85FuwF9yD8/yUNNvQxAAiER74J9BOVir6UjvjBn7SOWSG0Q/I+
uVWIpo93FQ1AuGz8kpjP/gc3X5FMN9M1R7/DAx6X2pJRRZm575iP6GObOKPNIAFz
WF2ElK4ZhTEm6v7RotKQknbrtSEeSMa4N7RoNjdFPhrzWFiCncqmtHxm4IjYuYIV
yT9reeuSkabPtP4mPfpJP3F8T+1iXPAvjieTZEyNXcKxsynQKh4mTtGFJp3aFxvn
f4n+rBnX3tuvd0f9RRvECcCqzypzyafnWOGyWSaIHokL1ghgbrl6MydVFAeI02o1
RyPCrjSIKd/qvKRg4qvXVxztIJz11vpj/6ZQazRxHpHJOwzxZMIRaktYjjWfkkky
l7YHFDOc7D9S0IbfI+1t3KNHuRRCM5amQ4I8XtgGq4J+keVBE3d2YfOcj2mMZfsA
H2lgBbD4jNwLJkMH2lEfTbv54VVoJSkwqsBINszslw1pjzD9wnkA1HRihwa302w7
chnc05OuaOp9DuT8sxsqWeZka1YBr0gFGzUJtOGXVAGKfLB4YPinNAb9C+QO5gf0
shGsGFFRD02k/ZFrBIdA79M44dXx1lOo6YrUtf3VnHty1MiALcR+8xaNO97SX/AM
iR5D86GGwarwposRrB4H6dFLJjZkHxgFujPT3qWDRBg1ZEftqeBZUEbvohSJvGVD
ngc67H0uG7uUVsgwphnDUnV8GSJ5BipTEeqbvwvFKsycfiyXVxF1NQJrja7j4y8F
9/HsRremIhmuNEmUFVRLnbWAvy9C6BSBlpEBeYk9Zdu23NRhcdFcB07aAWFeAI5I
UvxQJl7tLtYbag1sjB53q1fhZeRgRxXlIlkfBpRg2d/zqwS7sCzC4ZsSW9y/mYJE
oOBsgBqN/QPdMVmUub2uxAx+dKCsJQvfAv43D1m6OzXrJt8wb6VhnErlSvh4tHi3
neYjNc41QXuy/xsosVuPlNn+Cf3PtXMu4ccvJVdTJf+2qDCLp+FUcSOtiRxI9PiD
Re1z0HyJv7PmDU5q9/tCegBcixHdMe3h8j/0D1ezhbRsSuBa9dfqy/L/ag8103hT
Za3WHzw2tPU+FkX8ISA7A1wPeFMGFPjmdRC3QdgE/rV7rBCG9rSVs/yM+ErPy3Z3
d8Fa+lAXL/dehk+A+RXtCK7yNwnm75K2KwBZX2AquAhFWep79I9E2O49WMtbntqr
rnhRNqun20IuhBkW+JxeNbwAGUjdzdbl+UUZ44dX/WkNqR1PJe51RoEWipWhAJxZ
X6MaRqxtSaP9JYlmj3xK0QLdiynbJshEyJ9/fxWA/esiLq3POmfa2neLnioTs4fu
WDT1Turey3LiMffRhOXJsofU9Dquoa+HeIGe9vCWCmx00cYTY5nu+1JLksFVfyl3
BC90+Lfc8pDO6EFBg01Tl56i1MgxWtTHRQdOnxJTJniBjIZ6OYgJpjoHSDpO7L/z
Ue+Gk6dCry3Wq79T5Dw/7FaVsQgdm/sYo0sVDnUXOlrsYqYs+Cv9Eb+OUNAtMhTH
e6Ah7Q8HG+rD0Wk6hP7JMbWAeKQSuLef5+jMQ6ZnhoBtqssQc1DACpouqeuiuf0S
PMRezSV1mh/VcNXbKIM86/uCvd/jyADx1n3tMlp9XFL72IXIJdgMA+ZpjQwkXbpA
eglVBqkedOECtuSJ6neNTf0MeOKp5t2IXPSfctkF1zzNx2PheWEikJ4glrHU1EMC
KmCc1SFHhQiXqOKGq+fVLZlTYKndx5o1WKefaqJ92+0hBR4b2zUkATCXMz+5Q/qA
qn++iEeLHxwPKv2zPTSq0s7fICSBhqRoXdQYEtcQ67i2YNEBoeazf422jJXdve4g
71Tmew1N25GUmd+MoubAj3oSchKrnpr0MccU5CbfZBvFeY2qanv9vwqVLF3Nqdkm
bU4dhC2QXacl8K7a5U3FWDaiRsK+J9rtYpt7Hrcmv9Xdux4lEsdwDVNnCbxKaeYH
sRdXfYeCEx9yMQL2qu1iAtfA8W4nSwOFE8DKw+gaSWBjWj+MFk8Wx0F9qP8yi6dd
+96q+Ere8Xf+wm39+uVunD0rqJ+c4vO8zqunmGP99/PNZDqgjs5hRXO5UIS17Jc4
Og9aKqJPtFrArlj+pmmdc2WAwIa7BxfIP0GV7BidnxdlUwywFBhhwtEiiy9u6v1I
o4G8gNiJcamRYbpOmb4KxkQ5kUuGnSYiJBV5R2h4N5racblfNiJ/qrnh3M7aXcSB
BnZ9gmTbG9TaJXmIW7yyUlqrtgjKCxmbM3rzqfYSWwiQLTaNwzJsN21gr+Q3l2ZN
8VqhbcSTNSVDwRyPRYNIpmTC/fV28gum7JyUTdBDTWOYTjRHJgE8k3gO4qK3PfNU
LySmp7hkKqKHxU78kYOi8lw2gWgwjnmQN0j0X6m9lybAkm6oHFJpKxK2Za18ma2v
ux8OKfvWew7qZW+r4nYqmVJ+5f9GudzcjnbS+gX8Z+XIylRH4avgaCmoe1w5ZY72
Xt9NK5Q8gmsB7+wXIEizntDBTUcrCGOvEBkE7uyqP7OuK78H/vea6sMgOQH1+ikm
JNUG3Y3EJSc6WWa8CTxW1J35C4iEDIj3NvjOg1hEraBqfy7xkzgujcnTpaizw121
fcvU3gofBEfwAtUJbi+Meie9CjYZryUdUqgH8E8AGm50NeqyN6vwzDTZxqCCqGlU
RZBg/RsWBp9Bch7uu0DP3KCVXclk0jN0K+pTQRUuoXxnTu3grrxLxrEUop7UN5qn
n7nK+84xloSunOL2/LMb3lPE+kJ8d9vOBHM89Ssm4vO0cUdd8mKAETac+hUWoo75
jPBpolKfAisvKDzRYOm/trxP3wwTDtiQcFTcyIPfGEqBILY7Fs/5OuGDWtZhgg+h
fEMs162nXU/CTGTvDqH//OwnebOEAdkEyZn5dJOvqJhhrrqvrutRdB7HvLFgpZmd
rRVbo9bE5Y0zFVKsXN5rvAzn1JMCamIld3BlE15fIeWf9/guJMQFHZHAZmXXMkjM
wdNv1ToQ24wbveqrIm0qDnHBDFelhFijI6aWc9mQys/Iumm5ontKhpk7e3YTTcUP
PWEHnTNxR+90AN5WGFE6A/vpu7Vn/h3ya5U0o5RtoNlOTeqjzLfcuOFpnboQLY/e
G9rZgt016Q+hOnG9QMfN7OW5IpaEZFOoz/qGISbLdqmTriRU7n+Ky/4qxDIlruSC
LV2i5QyFymA7lH6H31xsexfyN1W99scd34Vu256iyexWrXgdmNAnRT8SmeHKEnHb
HaAj3gGFf54HVfNYaOuBQosmfKzu6T2poqSRRmJnFrabD6aQYLIDu7cDQV7LjvjQ
qRLyebX6cpz7dXNHu3sCqBhaECzpcCdBR1weMu4pmIcwVvaAcKkFCttm3Qj8IVbT
A14KmbokxxOZASho0sUoRvpViQS9V6qJSt6EzSoMONrJcp859c60mJjQnug1WdYZ
pR4yzkV5I3aolnUZ2ss3VUZk5uiW2vrAZ3adkuC8iZXVI+CiUSFUQ4N4s/Kzcxd9
HsbnpsRm82z9GwDLpwseB54ZDtpmkemQf0RpCrwEl7/7FSWuNu96ki1yh2r/Mnqr
2e+v1onWx2fTKfnghgiaU0kDyDcS2WTARwnt5DUtwqoL87VHoU59uHVpSsb09eOA
06sgqEFsoO5lPT1YJ8RG3xmuA+KA0PXoA6dVgaAog2WcLQs8T5HZi5iyRFxN/p1i
/5bTK0K5zGOEcLIVYnpBt5+d0vdCMLMzQDG/a2EN5LjWqitMzaozYUQQG0E0Rg2o
drVhnr7giJx53t1L3fJyXutNw1Xii57OYSiZwOrbwrnXp56rmQrHjEzX6elQKjzU
hru2XA4VBOxqI3LET7IZ0YpZdXQEBg5QWe0R6nJmd83nigr8q9X7dnj98jZ/9blv
8uJJIs4zC5yJulrJJ77SILrcHNvFrKqh311M/auAbz7NG1KNtIU/XP/I2Wc0mNsB
8fxD2SpfW4ycGD2tLdbdZ5rcfJNVIIDebi9BZAw1bz/wRniM7hPu14AI9y/FIoO7
uvIEO//ZC+OsYMpAmI0ZqpQ7PQkGMUw+h9Nz6zCpgwf5sDP+YKPF9O4y1L0tvY+J
cpVmf9EB3+4z9Rjiida3gkG83zSknjRr2D4ewVvz6CVWOCJ5m1UlcFl+mCDBDbi1
0PpuBlK+5BTIYrO8PFyxN2Njq1q4MjJhg8F/Pb3Ma0KB9qeY3V+dwDQyJRAr79jb
luqh7KeMzTnVTpcRbgOf4LlSfewLpt2wTJvKGfqnwcUegETh6Y/Zhas6xwa2hdt6
1nJD0jK+GOQ8bWrFFHrTPwUnzeM+Q3OCqoWqcZ8gessiRU0vFY1/fyGbwdl+Gmvs
kaQbNTYs/ck/60deHBUqffdCiMk/4yxFKiWtooaUtRiffdLWY8EP9jcPmUDxOQzv
Sz2KJCAO9d8grkkIzW0zZ2MY5PpkIFNm3fhGckslAmMTD+tzttFOq51f7aSbwTy6
p6FttvwbzKzjoQXzyqS+hxLPamVQ0gB93bGE81qlfqarIPh503ynLlFW4qZQjL9e
HBTsteXQhRz7n23Y4RjS42DxjG1P7kiJwZAC9LmxHnI98sjKslCD6FXplw0HxayX
+VZNlnSccz3BZOoBlPrZWWMmfoCu0kmoCNG6ColSsGkonI7+jmDK/TtzH1aLJr74
+MKDS7JMNp9dIITLYWk3rdPdGMOdSG8DT3YNiGT4E6yiyn3qjYcfpxBh6acy3h6s
nIKQjxn835B8u5bmqr3pQMAljbhZphY1H4HueoaA+Hy2SXlt6aiVDzqo2PTx+1g1
jfO3dyUKotJ8Th4h8Mg5Ny9CDZjLcDlJfIYe+rENXrFJIkOGsrKFINwFWDO6bAJm
5hHA2TSW4W5+A36g2jQ1wagxdn1eZU2KCJmGyEunzJMDbMbHBq+4UYrHdTt3o0j1
Iaq4LDuVLlC8ONYJ73+MhqWe+ujPJEwNMdtQAvAfVmyY27A//i+p2ILTNYd/81kk
WOCoTVYR00u/q6LgtnqbQv1i3f0pyTRHaSL9lLCvtnO21zWPuj34K6tmKLo/jZkj
ziWnW768MRkm0YtmC9vYLYnlFAFnqEEx5XwU4wWE+JVGzA3JxWppTzGRYEpfLA/i
sJACv4s6kcsQBfZPvzV5f9MjGmd64EnHZm+7tXZjaPEv17NbHpYgVbE+7CQswFXS
mMVkj/YZQTTmDM9L8yHgeohAE52MG2SZWKL438KvTNVsp8OnpBeE/j8N5GjW+Cum
Mn3+/xQdwgGZ3yH3E3USMJrjGSSg9tKfHA6yVSXBbqvV2QhEwhHrSZli3mSgluBb
D/jiWrOHYYLN2+cKNil7i0dg7y1RZFxJwLa1C8n8YpcdPIbpzs5n+abBkkPKpFI4
gp07poMNPQrpZyy1aVOMnUzyAnV6NWy27/e66LMIbK4SCs3SQUlfzPMUjKH7zxnj
svknh0gsBCwnuOQnojxiYUZHHY49KnUP1DbPzKd5anPhleUvUs2n52mFLgNAwi7+
yeVLveoAeG1EeD01nmvXbp5V3AxYBFd+ulWK3Dq9h/9bap7/GQ75N7g3B+Q4t7Hg
KcFHEPt/hOx3B7AkwUftQMKBZDbvfpCR41PV4dqEicFNhpkp/q7OQyQpfliTctrW
dni+ioYvS74sOI3ozOu1Zn0kBaU81QbTK3TsYWtSEz1BtoCux8J1qttock0yC3Bo
GJHTqPT3AfI4PnnhiQrnSfwQTef1OinXgDzjmaTtLVFr5GUJiKULk3a1EBeokjw5
wxxHHNGDuQs6hUAxY1nWYhzZzQnaBvyMFGdspjqWqAn6jcUu/aBybVoa15ZgTDct
iB9wkGmLHHW9YQzhVpeQDW+6/f5bF7EeXpOrdRTXLvtrAaBQoP43I3Omcd6V5qjk
EHSgXXTHIf4IFP0qo+znWDKonUqyw/JKRUXNkQgsJjFeLgw1WXSDo58AYow9hjM+
pC5FhtfFkGND79sD8gZVUNdCiHA/cq04Y1PpVtVMtC89ly+uqK8fIdABdY439B/N
an1IjsobrCXqGt5KeHCe6d3sO7CU1EMcQPk0slpBhER6zGA5TS7/ID6txQbpk85X
UmBScxoUAuerLReWPDu1gtXLfS8N3Klo6PimLA1TiqQkQO1aj/pCeYaOnDRHpZmu
ynUyDeMaNE2MMs4ZRTlYDjrEAaPEuJJNXIkGT/BIFABsgyM60zVnaOrIW9I4YDLa
/Lj2qBblkpBNzCPeLYh/PECSTPrWqunihdHb1kTRS1NvDN1+tBiFqegejPB/poJm
bRvAvwJuDMuI1cS2XIapfAG8sLkd514uskm0omOeEbHutMZeUqDGQy8b0X0ZZPX/
gbEBeDSm4XxafRc5MWjckBpSSoMIvoRcfArVJCap9pkk3hkPkAgGJ8lsTNKBTEyD
amrA/HTij3CFWtdPfb3AMYeW98tLgKiMyWZIFtlJD3v/0d0Dj956MD/oQaaIiU0D
5S3KXLUsKnurCtPel+XDnQDyQ/VyYHL5BJxy1cXlVZwkQkfNOGsfjqOvVbUHIFND
O1s7qI6ZrqcvQayg07UHPNYgGbRRKUnZuibkg6fPGjkBAFa9LPqSEDzP8wAqTS3H
fCWSPYwpxN5xkXFUKyzNuPqrXdI/BZwNyLq1VavpOIY+K0mSN4UhoQMqJu6JPaey
p+bp7ZlOQyi3YCZIdx9jFsWeJQKYa6f6n5Q66XdwAKTDrqUAiohXwXQr/nDUspBb
145IFT9Sq3oRQHhD8A1ckAuxobbNvO7Wq/LvafzsjOzc6KGJkUbDxss2PKwf5emT
hbOCKsnocc9qb4WKs1CzkemFk1Jjn1ghpArUcAS7rFUtxS2slM1GdpwxQiGDgWhZ
zzDCEl+OasgPWZAaiNzlUFjgKHT/yBedpa2S/+/j1YAmExOcKL8nrcWqWkFgCLaL
OZz1moz+N9aRTpwdIjiaCwVS9WLeEzbVuHJGurTs8XDyD7bM6DHCJskpF3R35pi0
8VUzeM3PacLngQbTe6NUJ+cWiGgFvQREOr6YVHjX2pQ/D6ESqkxv/AsYTLU/YuR+
vce3v3oisMDeLBOymMh8PbuZF6UUBMz3tjCp9V2/QbNm9WmiFmXWI8CqP5g+xjzQ
CGXzuIXyB1UDqefq0AcT9vrpRUV+kIenXYCXXf3lQK5mfhOjlK+yomjU6aK9PWHq
b3vmzG0QkbrW8ffbSpdUxNi5kr7TQd934IydI+IShFpMVC/YJmTDXexNVVdAgHxR
hGUxOP2Lu8W4LJ0ISQTT7QQ/BPYqeKGAFGwPVLM0od0alKhJyu3pAqIu0YzebMVy
oC8XLWqoU0vkWBPs32rdZT2W65QCaJ/FsOVh6lkwUCzAzigcCniLowmciCAYMtk9
O3sNXOdWQ+J8c4tbddoXRJ+UCLyz0aPqBAMCbCM0Aa8B9Cm0/7SZgXlEfbkKWeeU
Z63MbRPspQSF45MYjI6ta1+4R6z1s8OGv5BtXCP1Mr/fNE7grhtCc3CE6i9e4EDT
ZR6A1w+tl1omOVQ3DcSNxpDkAPQjkvo74GiDWXoDNvFoZ2A0Zu6YOP+wOqKrPFuQ
p1i7vmoHEz4oFjJYB3ecX6GovE1mRSC3DKfUTIf9uRd8FTeCCXVcQbjLBlMqg+mZ
aU+zy2Ru6l0h95H5/8DlYguwwGxPWwAcXGoXwKiqNS0OfMR9M8JAx/7DIeL6xhdH
V7kLxjWLXrwiNlUynBV8HZ7C12CMf5qdzhY/rU6ubcNUYCnW9Vyd5WrVprnuaJmT
gpSOMeQFIuU+1ucRILVwkI1yBO71r3ARzjOJnZ9FFCjb7hWFbI11eTuTzPfcGKdk
7y7Zbl52TyGmex9b6FbdTY7mZp0bUEbKmLbMd2vQ0LLkCUegWLrq5jVQrmy6wzh5
YYsc5p0tHC9JA3zcuAOTwQJL2IRkGYAtm4+oeI2luqHvBqeXQopCe1UwnYFqOv2j
estvRPONio6HfPYyY643vWFRuh8cuNokgZWnqDW1TR9r1/kHUQZEHvF1XzjNSnRi
Uhbs27smQRB6pVs1Y2z57Tn1jwt6U0fKZyJlNUYBFL4Pc9SqNpzJhb5ltVRu9N9N
3dqCbXDUt1WHAQpWXmNB/EfsaQLdRNsqamg/QpUxvLMmrQfs2rHsbhhOrJt4dKMC
/4GpeRKpm4mWl+lvgG/gLdPc3/T6UquSdXTaHCNYbie9T94X7n8HgVkGye2GxNs5
KiXlRvBTWdITjBQOhFaM2vZe4W/cUhlWrP4R/93IZ51xfQtbc8dGAy51rKf1PtqJ
o21TKU8n0EVeOs5PQOufLUHKipEmUo6ZSibz0Nl8JOhU7t6DfAI51cs0rAJSUECH
Lu5Gj7W7nxUVdY+tvU+7R2wddaPflE140ZdziGG/m6QQ/+ovY3lteCJMyZ7pWQUs
9EejrEs0jLGmrbxhYBXlhv9wBQCsvU+RftIpu0lAf3nRQE1tGcW/PgUL06CDYBxf
80GxOG8AuQRHNNKfRqOgbEa3+f6X/C3G8pr5OXQAIypOEMQc0KYoi4nb/bFjuBM+
kEOM8JR5raZy21k5KaA8eUXKs48eGcWKmfIinTx3AOvR6oJVl+4ahfB+n0zRnOzd
UtcOTjsCb91OjchoIiuKz27CNvPum87t/YnUj7xJnt++KTIxaTsmZlztvO876OGD
7blaIXBA5D+YsyfYDxdtQRbunKvUyMlPaBkOj88qWh7jL0FQLTaN6d9oDflDCbDs
UKv6nJY5+jNYbpsxj/D6cpG+Hko1CsD2vKwkVxsidiURUC2mIOzUKoaxXZSQXnbO
IHLxmBSzVpE2+WUBi3Gf/fRm6m6nm5gN1rMuohMdbHrrr02Xf1sU+3osy/75tmoZ
iM1OE5XVCtv/g3Jip/Wt7RfoTiN4AiAi9TChdfeC28kRORmbqbnvV/A+4sF5pRTi
CuiBFC+oTDWHdwXuoKU5lDYS2QsmELm7u55xj5lySv61cPjoe59Y32v5+tq7y8Ri
M10BES0R6Aaskd9tbPyVL7HWG2FDMwtTIAbnrU0OreQAW8RsV1VNmIns/dLRZ3or
AgdtqlIgia3au0pILEYEqF1KHHppRhkZBZ91/CTG1Cp3Lcp+p1O67IFnVaMb7A9R
ayuCZ3EVwicGlBBQlHFPDilMDH+CSkgCYHIqOX81gYUEFUb2d1KLcLQTa+1h7l9+
Mjga4QI6BWl+Yai6LSMFWj+edRfaMI6sm6mcIuNo47wL8C4gJnguiC5gl4Gys/vW
WqCFhDUrryA+d3Z4kwSosllYrIwycHbmp9N2w6lS0XykqURJ/5lNVLyxb8W0a/cT
4S1XYaTaN/qgpjROplwzWYru2pjupgeUwLRzakS27e4GvQyewKsPdLcAcltLxAim
L9jA8VyYyQR7fm5telh8F7odY869hPYaIbOKSLkzIIx/pXHUmXTi5qXRW1pjbqRR
ofTjmju9X4eOmOTnIJO78IXW6DetBE0k85RLqk+m1Ya8fKyRRUHgqK1n/KjIINeT
gE8zrxgeSUfZZy9q800zFl4u2oLPHtUhvE+Eq/tX+RwXTxZ8c+nkJBHggO4nbZ4f
wzRt1MgWsluAoXF75N6iZDH3gorLEIXaaTagWab3bxOVGf91uYzSqALCAvaN4AdG
fhp5/g18BHkSht/myhaubxM93+MfOzBU+Ulfsta/JEf8UZRd6bs93W3H0PN1cuCs
oBmFOsJy9JPCOZ5SbZ0lhr2Bgmy6Vdls6XCi+gZQXaurkqmv4H3KPm1fp9zqLaHq
OGHJmIH9TJXWHWKt4RJpHdQoE7Qosht5hsoNMrGWPvuIyMyon1SqeScfd1Q9v/oa
xW653tBG+n1MdYUQx+cXTXKnQvYDbVLC8t1y5nurqVHOEv2GdogQ3J9Kq7366KWJ
pGx56aS1+sSddHNQt2uJlIBKY/Z98VnR8g4TS38kvQLUuOXuEJukIVeyof/VJlL1
K0rElx22Rq5DQFBHYe/bvvjiZw2Zm0t/EqjJjkddQvvRERPseqY1h2FALg8YbgTz
ST8Nd6HIGzy9SR/+OhXGRrH8NTmpAiEW5K4Vl1gkN5BDHsCsURX271vFrJerybus
j8AJ4WKRNTkalVwtwZg07w/7pOdBkZofh/iB0iIZmq10vlEEpL1l1cJBwqD+n8CB
m5ew4+3x6sqZ2dMVnrWEOeH80zLSPIWYyl4tBXZIqrdeAE44qEBzdhkQNGTPUDpB
nryoHONtmhY1s+dXKShl7sNgEiv6gvQeM839kgZ82KAhyyBoKxSzU7IzgB/YvKmQ
5xnaPwFVNYttjmoILK0WFm7PfqSfaYjW+5BRvbEDSwSl5NL1fMzBKqYfJW5I41ic
1je/OgjXFCKtubcn/WPZ/8WtUEvUbcosBD7fLXS9Njz5wIskmKWLgV7fdc2583C8
f0WibKDwepD83zWYbTLEa5aOEBm98m4TzvjdEKFsr2FO9EduOlZzBBzdWtdzft5u
KofccqH0M0Tibs8eAaP3/XbL9PbYmKRJBkhEHDReEmPao2BzyvRpmu7KuzAFO/Qv
d/lCQYmUIdstfcOd59iWiJP6KuEalwcDs6Ap/mE1rzfFzA8qZo8ZvSg4gvM3HLlL
cEMZT39cMfQJ6X7GsG21k9Eh55DAWsgdqL8JpeHPv90pMpbLjPKCbCyPpMLCS74m
9yZYXCZ+VlkXQVQtyiigXbJpVP2rAeUzu9VS7yH6APNLC37VdDbav1cH9yoS8qZ1
rpq/ifBwkEk4ePeUbXD0Q/5Hg7DtIaXTyqbnxy6xW4Z2zjAUC33y8DA6qzGfgOKX
8sj+AfD2AcHiIiFfGYTXffyQcndbPqY72TCDl/bUCujhHVAQAY917MoEUtIJfvpq
re5NfkQ/+3NW+PB3VlLM5vAnkHLlAT6Ico4PQD3OP5yfX/wgTiFKhq8ynvESlLWh
blNf7fObSHZvIlu1Y/rKbMnf1VuIOYBUACeodp7r+UhEHhZehNaew2R3mpdpOY2B
RBb4+uNQGABTbwS8dMP0FUUCYOsGpZv0JEG3jY5vOu16HQGnm4+JeypvkRnf/md4
bOHd8TQcobUorwbni/m91qBUxV6E0qEpvjVcxFuC/RhXB5F6nW+fM2Por32JbCOc
uCwd0PghzisStglsmkRJdjuD6g9r12ZyISeGXGnNgOX3Lv93BEm6gZqnj3EJk4kK
P9gInW6062ChrXWCOYTetudab2kmf8kf6zNvw06A7y0lTSQjZ/XCROq8IsT4gj/I
S0ZclPcYo4DmVIB6/0J4Q3VwYSIf5hkOQI22NQ2hqGZuWdNZ6bPknAileJCSj5J3
sRB1lDwLNptL76yb90HyQQGGixaw2LfsY+OzWD34YWbdKtGQsY5dTEKMWRfLBoaB
NG3T43fpunY3zgObtKCjANviTbBT+OY7elSSk8+0T7y/FfeFTvTqwgCVnlc+rMAv
upmO35bOg48DEzISBVX9LSMGiLy0AWJH2zyAM77MZNLXBq6ppmF3p8G/fMZWHcEL
Vjr/TAfNzgX2hHuZYKsE6jxLz6lgwMJ/bKlfdeIlGIfxRhesFVUBVx2AZ5V+jl3H
PLzuJoScQ/4acqRy1gO9tU19OVMQm0BX2Gk4yt2hZWPaKJNwWiUu2UikA1FhxcQf
S0gv371dTHTaYAurtyGdknXA8wAbvGqqKjXtiW2y5myJ61B1GO9+ENdid4H7whtw
wBY5xPDJFJeAlEGczomRoNiwbkwND5CmJbPphYRbr7I+lQIJOn+zFSRL2sRhr/fB
i47ftaq/awz2oJFXA0l93Paa+677IaKuHOUEh5Lfl3ZEEFXk/hm3Ou2HKe7kR0Nw
pCp5HPDguB+rqPJnlk6EL5eib5bRSO7vKpmhF5zmUU2FiY4y1aKIYN5LQZf3pJKc
S/FhDJqaYyt1aEmLtsa578qs0kmKlJd5vS28NdD8plTM7qHPFgY9wd5xFvYsePsG
8QNF/DrVpvHkS4zBYGaKzDOmlT3+9H5ggXFbKVwy/9mjbocFU+9twSn/8lGpWS6d
ewiBzlB5yhSDcP+5m+0xayWP4pGm+BHmrAJcb+HTmZOLRBfz4aPeWwGsJEpWDBAJ
kwsXUokqy+zg6edY/MZMcw+QLXPpiwzB5neay8VGTwCZn8zA7ZlUllnnAj98Ekgt
EMUr0/FYE2XFuhkTVuPOf4TtKMPZMhcLVYWF2y2YwqYZ4wAjZcEZsuxhC5+32us1
sZkZ2WN2HFVcIFXFkW/ALR1eao2Ce9m3SBo/naTqY1RcVP5C6vCd36XgzclpTZNr
+vhmwLmcZqY9qpRU6QPJ866+4zueSjtiNFeIF0WbXQx6OlbhVbgH6tsqOqWifUi2
J63BF3ZcJpeLxP/5wtKhnUWGMhCx46wxGBDDsGwHr3SK0ImMw1wELEhq0j174gET
YSk20yNhq1NbKB3c6jFmE/KoqeMxjGZL0G+KfcYTWDQGO/klZR5dG/d/FrYugN1j
72uu/iKW3H0P5egJxPp6VJpY5PjIZsd3RrxA3mJ28XzAUixoThwzQ4vJQKCo8e/N
Ax20Iko8+qid7FYS+Es38vmmZ67V7Kzdppx4DUzA/6iL/4RM/wZhXKkiQCfVSrQt
AybzCgAwe+2Ydq2R8KXImER4A/YiV5MBsMU3sZm55DwhGxHI0m4XKZy+yrgHHbU6
59v0zweo5p5q70yUHf+OWoqjiXjBaVUaYXqZs1PUHcqSIRP+NP7FO6GZyKJAzI7v
3aRFgrQ57F5pMREIZKYQyBkCUZh+dVqvg+NJzmnbJSCjw6OdburqZxzwA16WZhUm
o05NyEZLhOsqlDfWiC8D9VApvrV4ieP7SyHYhPDVClAhlP2H2l6Ozsmc38Zi7ESs
vCHdZyy/pSwmtYg2rSrl4yiphm3daQldgC1NOzwXkErbPpL3+S+fB0JshuCd1iWe
fZCw0KrHAxtc3FkO2G8FEv/23QCrIy9L6zIHfeLJeYi0vF+joDkC3UVoUDSTVjTu
WtVn8hIMMMiOrXEgSQ37FO5sgCbagCiAkEGFducA7viP7TDIT0gOmUBCLcqlwP6/
dAHo2mPrtVGmpy5s71Uz0zlG4rKFpQvI2QrFdR7naUCStp7QF0SAqw9EFkHElSuX
PaaaxhdVyCLoAsjr5+oyK35dx44+965zcorck+2RaW94vioTaGjEf/bbWFJtAUez
jMvK9XHPZqFE3GH6cK3bEp2C5MQ4MKfLAQVYseWQql88BWWiKZ01IO0vQ/v2evVu
ZsKHa0okvrjFeacaK0pJQnaJhY/Ys2uS+Lq2JvquKZ2Bu8+I6TxBmXChVXE0HcwU
nd6wcCDoix+Y/IPYBAgAbQZKE3Cdk26xpyZATJjte6nuJBnehp40y0DmSkYuRHtg
8+EVdIoyziqgtTGfMU6HhtdRvd9jqF/9Uaiov5HItBAyEBJXS1WWd0fFZXYzxBBw
dZE42iSVjmxNqT3NW6xhVnEtXyikhI9L/d0cGXnYtNi4ZXbSfTtoWrT0nWIj+YjQ
rTS+YJ0yfPbBJkpwOOSB5a5p+f/lX2QB49R5xz9eEJ99nDjAQh1K/nU9mUslXkmO
LIwQ2T6Nk3gtQ8c5TCToUBv/nI7LffOTG/kHfAOn7mQbpMmUjB2Ck0FmWXSMYsDg
hjcq5z5zCtvqrB4/Xs3xgOFta2RXfs6e7lZRN9mvDNfklo3srVhtksY83hzFv7We
qR1/dy9trF+c6/JqWXi2AFAMDNXW6GRzhloYCA2QZfeEmBnqLl3vG9NShwdAitki
/JIIZL4WFIMWWWetGgYRwWCJKlPE9Td/chDVH31H5UhsvzD0XDheJYDaO7dkwnTm
WyTwpYRg5nlboirDNPfSksYPul6BvR+QboEI7SXJJ8MNCIz0dA/FNeliKHkgJCz5
be6x++HKjvo40pmTYRIInxXss79txgUMLwucUOvGmPMKnbKH1D2uS9K2ivWKdO1q
P8uLd4K70JBFWlNloh+N0gVy9yJWseAnsyHA4ZxRmXHr42y+rIDSRGFWeQNzfe9d
vB/XWYRGPvnuXwe3vFiD1qJ8WwVjAkuYmFA6/Qv6Sk3ELSxFGXK2Wd0oiQZ0tQKM
UPHu2SjBwcaD/arfLnLl4CRJT8fqBephRlo0ldIbES2ld+Md/fdglkaSaMgtRmro
LTksYKTf+S/eQmmtU8qazzQ3JIaSwFbfhwDVt9A9QQrsXU6DIFOKz5coQQGxV+sQ
zjTf5gkX/f4wpZgPZy2QsZ5nMGVYMc0f9Sd6zzD7rJV9OwrDNNrWVvvlWPUHv4S2
bcMX6ZO4tf56ANRxrwn1SITTvdMyA0mk6wSfgGBt6HtkmWcrhRjATjQIh92hsviN
/vmIEUCpYIMgMqfyzuLXQSNQJ20wFXkxTuxiSgmPvWlmEL0YDJDgqJvxla46Zab5
MBeWzoww9jtUV0hWRSeaID11KBuQBsfLu8Q+AmXOLDSbcpEGu3OsZal5MoT+mBVU
yEaKVF3uJj+eo58Ducr+o9IrZJGNvcrTbANMbk7bzr7qD+0RcrLUQvHwyKNmdMby
WY8jDRSo/eLOpFdnXF/upGBlv+iCJpFqgv6+4Bp3NH+BuGja/cGZSE19S3zZv4i8
b1HW9rO/9Xxv8ysDAl7fub+5rzlx2+UDC9xN2K4n9hz/2osBnU6VpArrw6//U+Zu
iLvO/MmnJNTLJ8WqcXVSn5mP/TbhE1tAHwRIONiNGsJywRVjxbhfJrOg8dtueSeh
bdN1Ccv4Jd5WjLcd/W+tGi2FjRzmm7ypuG8JK+YcT5sDHj1VNldhV3q5PcRnncvl
8AedlEYDcXPnX3dx5IkTgi+ORN+DGAamSwk9AkLJ89SXPFT2RCENNnDh+mpPlHjo
o90ADCmYhRc3UEYg88JHrmDxQaXzPepm90zAwtS7JhXGQFKkwCVetE44yLwkKkJa
3OVl/lieMCKqOzX6O5RYw+ZT+FVFHkHSXtyecJpgu5BRVzj4eUuW8iYuv/HH3JFy
mDgWQxGHsykVVA2N7cnUcTXpGxY5fYrKAgUP/b3JvDNhPuPtBGo1bnj1Gcqd/nv9
cptex9beSNAuQhSKoxW2lI4je7FcEX0c5xMsab2cYSBGDi4EvlAdjuPZU9XQp/a2
Zfz7frpD/HhFNIpKT72Nsq2IaUhpKQ1bBE1sBZtMBrnUFePhbX5hcuRrXVhe+oZx
U4I2NAFwDwP0g7sMsPpvSIh1RqfNBi56h6Snc0Bp4SdY7TQth5rS4TNwuxvnM4ZM
JpW2gn070xnHlJi1djJHRv6IQmhcCO+zATX6+TEM8KEoThMu2unCItjv+RBCQInT
ICVS4AAPwBDDqTurM6L564vWmZ6iT4TVTMGxuIClzU3jBp1UcFqazx5Imm+sFFJ+
lrZrjMEyV6/FGrFzBGEHCfs7TW8rW9LFjNtWsBoz5LMlWS1HQ+pAlorFKVTfNgiR
9KeVhDm5P2IGvYUtAXOYg6ix+B52vzvXEUhy46+xXSpsPOpiigeE1WuYYc2qdXNM
Soq7FcoqMEoSfKzclAzlon28+Jt/N9D/x61uvFSRXOS3JrpW67YW7ee1fRMSbYAo
f4++qkqK4Z82U4IuWqdEBY2BNtvuebBaIUNsqUr4XHw+5qckpeHbToKqgZlY816H
tsXB9ipaiYWAuKNH4UVy83mS8nqOPPyQ04suYesWRysBs+K1X4df+i6nW7gx2TmO
C0gPwOmQ4m9CK8u9KitDd2qFz15qhXiP++SHyGFC6smS1UL4SF3iuJAbTMj3zscG
A4jdGiRX3g6SQvWSVCpl0/7JBhHOa+0Nuf9tKv/7mbxeCCngWHwYnnbpWu50iDHa
wmkf0LM5RlJp2lK4+XpykS1FTOzszihf1fZEB5x742HgWr6m9Geiwl7xuwz5qNkK
lfFCEDCWWmCNxhyJWVSSJUTRVsMbULp0Hpax/7OH3ZH9pd0hfgOZtvqL4MeDF3JK
49ie2UvhupEZP9BZ4dGphvVIjP8CmFdFzGOjBDvWZkszbYHNx6qVJWL4x7P5VlM/
3awUTzOxfi9BRl5fmftwR1jKXHHmvfeGJtgjaordll99FdJuiu+du3rAU3R8/MA7
Zrbi+nZuqMNiENaoh7QYQp2dafrNR8PC0a4xGB03S388ScbX6vE7E4th/fRDPL51
ydfRYUC4HN3NgWlJZ9/y0N7u0HJ9G10oZpizAr7uGXP0CnbRWB2lvD/sxVADghxd
g7mP947qZIbeOX6bAlweWVq664ddeioebQLeh+MNFgRjo/GwyoJho3gk50DiqPPS
SVDi7zrXvpbB7/eqZBeH+Ys0Xn4Ga92CVSmhSUk7yDNmOwKML4zVQHvGP0lIfAw4
fRZY+Ph6Jn65U33/Z1ZTzuwpbWXPoCpfnKVhmTAta2gX/7aCsg1CiE2S4ZY+5lcf
1/E+r5G/OQueGRBR9OmyA3nIljsRGWEKlSs23LIOZkjYwVf8dmtuSFHafRyL1g2a
8GTlSU05Au7ZFq8HWHfav9fhiwWlhuSKETYrJUOapikSki2IBRkwP6Eom3uvD9ve
oJymUwPNTgi7AtZvmEk4noJO0bnZhQZj/JWOVHbcLR2jwUygFmM4fDjmSSj6QCFf
yecLcB74NYGwLGODYjGrwg6SIIN/51vkjMFSI4ebAcoyZjH6/DCo8eMl+Jb5HJ4+
h3oZrqvJvW4M9Xn5qqe9RCaERbzp9XV5SIZjH/Ga1cpthsVt3dQeMcqTXVNpIpCZ
GrDIVBkX1y0ovRGeZrDO7yVP+CrZIqZz1+wk4+JAzZEz6cSD9HSzzjSevkXKbZ2z
Z7jWfEtM0/86y5ub7dCm8KE36wHPfB4BNo7HNXeV/DdcfBjPHk1kyEQetBW00DgP
2P7IFiBDrh/9AuJCgWMmtEfRgKwBQvm7ryzc+mLuUqM4xvhh03aZtcU/zH9UUK1l
VjsgK/gysn1oB5BEKipQoriMrl1VQuvJNyt1nGvH5rUeiiTJM7nE4l5CcqASw33h
BOtrmwqRqja+B5BNFDwo3VacnfxiUPqo5hrkVfJ5yYvqEux+GpcE1uWzr+uq4T22
3Me+LveJ5pV+ZYgR7sKpIdzSD3942AQIQ65OFD6SwBUNDSxAZrIE7KqvACTXvZZ0
9jogYYtEEwsf1oSoc7fhixPZNssTE6BpCDLKtmPEXTJnDgC4nY9+kp5yX6950TjK
YILxR+DkSJGKqJaCZyn3K0Hku9HU0X4DAJwgTThE0mzvOKuQ4Kb1DnAj8pc3PE0J
XlZAlBosb8uPIsjv7hf794dYp8w/z/eVl9pTfPBb1nPicYaTow4PbUs+G+U51dPu
+SoNL84De3+PDVWb0XuKj9mtAiqjA0djL5errEJgBY4ISe3+mUzCMkXVtpAgMwHY
Mk5tQG/2RQWw8wnJPVUikYMgTB1dLnlTCBXhuogqkdJPoAg3gPiHamqQoUvDFoeg
9Dz9AI9pHg2o2G+WdAuFuNBeFRVjLhuC9JDL/mXuaMvuyHjf4rMOQvwc5Yoex+7S
6SKwmQbNWI7OxcUepkrQUfZNt3eHzv9hQ09V1oi9POMlo7UFj4urCwDuJcuGO6uJ
RRdFNDauONzCaVAyakncvdC710ONklAcD3YXAvT20UIHuiCRG+jjwFNt/uR4DvUO
C4XZA5yV7r94S/j8Yq8nQNYTEjyA716cXBGNkkAaBovU5Oi5UVI17bh+tWsXP2HJ
LBkIx3kZZTdBEnMEEgy0zPd9QaN++f8DV14CzyAbr2S5/q1dRnxywZ8eac35mWd7
JnlTVVJg1+t0ezvLfTKucqFF0pXstU0QrQ3ApK4qEPwhBerVT1ZWHGvkP1V5dbrr
xyJKlWs+STdhXtG0zSGHKRCWhGd8BBz+DMifTpBj7piOAbRXDEuey6mM9RMq23jz
XxSpe2BnXi2gauvQND4YJvmQYJ9mrTB619+bi5Q2xGBoktjVD8/16igdALHJp7cg
rk9PiaguH77Rd2Hh0rmIZ8JdYRztewwzCIVEjPI+cqE9ilHWNqIvGwJIKIocxnhB
a/g5130cvN8xUhGIulkkbsnakEEgp4HXgnEIGX61EPtDh+fgu3GdXAKb23ziwLv2
82r9ivD0WysSDGadIU+MB2IwtsznJSfKylEfeVTdWxEsuf+HXq1UOKSvsd42kiil
Wl670493VWI3yCbDMQnN01TKHJohGe3r0ah9kB9WLlPnP6EoQHdkNYFDyiWR285h
uG0EvHmlwhLZaj7ZzudBMh4RHOnzEkSjsuJ8dvAwXzHRpbPgKOB75JeStzn60uaY
+jDckrTlk3RdFKU/8yisVcTWBLufGYZKJJ+L6t04nQqF6tHoqgbjnF66ndtHVjAK
xtthS7Uel4QT8ohN1ZQqi+w5GjPGk77ducgv9Yk5Ioj6qQcQDdFis1dfvP1uQaxt
AfJGQBezRce5Kf63hDdkXqheZ+sF6jOUhErEKto8UNNXhdphJXFz6HuoGI7eISV1
W9Lm334Nt6ktPTBbR5J+J/8Xh2g2fMGQClgSBC/MQ1lj258Wgpbbhd/GsD1D5wYB
P+NJmENcIbjLHidJuO64TSL0pvqfT2UtPudEaw1D9t+L12x7IcOgdZu6vxVp3GbB
VxiUJjE6hbkzEghzbJ/SMQOGvzCjW3/bhjf6ijRjWndasxEClU6m4whvvTxFoRoq
rhOcGuzf+SpGbguJAUkSnjFRJwxy6CEzT5VJZApzaYn007Pl8PDMzZqO7+6e1HeK
G7kKIFdruC5/i9Ktacm9AGLzoQ306Ig0vPydSiDBi9+hNldR0Dfz4JChcCTm6OgS
/HZPILGJ/mKWB1b6ADeKrj+ptxtgaFPNmR2dOMAMt9PHkPtSa2oxoHiXoVLJADO5
5K9D8Td2X/9hL0yMBRwsP4zBtxfYvR55LG6dwVB4XF2J8yZM8oJOYeuHvcSES9RS
rt4RWHDXEdoESfXgDsHDspTdpOtiDVlHzSx9jQMlCBihd9ovdd4560+68L3tZtHd
5+PkcuMJaJ3YA1/ckXsFolSgwy9dTV6RpAN4Po/bVI1PYYcY17kgasb1LTHhpfJu
AGU51kx569irU4cOe5UbmR3i1IdZcrSU5Had+ukZvHiVcY4cxkF9kX+b6Ozj9wWp
hdICrlaf5ybOMUu7qsUNDeu5FMzZ2ez2s864pmEfS+2ebnEeZG8lBz6u7wOxQqUO
HQ8JgCux4M4odWJSW+8l6ARdEtUBjxZGBUPsL1qoEl/GYI4gp5lWqMu5ZsD7qqio
qoBmW0RRptV1weVRRSlXe1u3GeI8Kp+d0n51j4ASrTFbHNUFsCNlPT7z9Ymv+l5E
/jSKZacSgVSOas+19DAVuemxZvO3k4cSSIFVXJZPdBsWF6v5YjPw5VJsHP2YeXbf
kive0nJHIN9vbaxSbvaYFOlYDXLmq0X4fNQdat8a0NVSiHGSkxqH0Txn2q/hk7Kk
SQgUxsGX87PWo+oBJAxZOBAdAHQmp1qq2x5BYFDpHjMsY/y+L5GBr2jZUzrKT0VR
+hAATDpuWs7VdUtC77CGrlBtNXoG0dlEhIAML0+qVJ+omDApOnw73hb0DIPq0fMj
Dzm31NBRg+XKuxkrrwYgvGvEO6k6pt3PZ38UmI9fl0xTirGLucoPF4kxdIbc5N/B
FNkxLzi7EK9wGaoqV0et3ex+LKfq3mFwS/YJhwKHuNoAK/K4Bs8ZpXMnre2l4Q17
CDlvbDDycw33lj9lvBBTeF/fQ3p4VLHPK/JD5Quxu7vXi3bdFJkRC7jjopGfTR3k
76fn8O9yVo1LZkr3LWLwQvCzkgRFi+V8KDxW53RaQfRrx+7jeGAwAdaf6xFByFSo
u3s97+3ngoySpMTAmDJthWc57pvHQ4hSNVq4dAYagRTDGJ53LobDdSXW/XXMSxmF
oMmrLLlj+yq1MpstObZuCrwbKwtUUX/d0imFBhwzvuQjrgW2/fKvO445O/Q2pEJp
+dzqTfyLMJ+MWYyeAwiNqXzi6N7iqdsar7T1h1gNL0IKNJjUjr6D7ZrUsFXBo4fD
3vKxsm0ki/iTDgj+3jlyOMeT1NK/cnaKYCfd6KT4Fo3CD5PSY3s8t03r3TZsvNVc
NXDOWOgiznXAUp3X/ICVGCNe0x2Z9qvHmiX8jyV64Q2ERXSR+AVbmzg2f/J6ZQtB
dhDRe3UT+vri4yJ5DYqT/qll2vukKRbPFPrQkNml5lrXFbUQ101rlWVikqIr5Hv5
9grML411PBiZcpPXICYNeQWEgGuRGGylCj1RxgPqXTOUKlWzwXoBvZ+mragPwefZ
sr6XbJHO5p1OiUwqk2SLjmChGaS0JFLuEo5A90yWL0Otwgn/0gpZ+66Zy9xPiacg
I1tEACNKUYsQX3hg9aK7YeICQ8hILh21r77iOtNKnBn/ms7LBCYDlCeaRlNXfQU4
v2Wj7+9XVEHmyapNSck765Io8Vx6AOnurk8xgyJlbnt+rUD6xkRVkEwnjuQibgBW
hcAOx0f+2+kc8ifpFLVr6UU9LOWtBs5Md/G9Jw8/8VjDL2sEim1KHsx2/YD0DSxd
ZbpoJYCD81YJm1M7fCfUNsnqWoFebI5wvawrVIXjtshIExIGSavMwH0ZEnhVz4ix
RJvhm5r/VAb9fOW0q7C0cEcLdC9zO/uDYTtMdxvMuBNgtDZ7pukMbSzQaS1a5EKU
Nkc7pzI9YLj/C1nZo3p7+RzHpCdC1gYIy6Mmgj+RPpP1eetOct+IlFJxnRslbik1
GiRU6nrKRKvDQV4UQXHjM1vEoy8xjKLSjI8M6KAjJ8TvGQ/2MMFS7CjAdbEmMhjw
HMeS7HayEnY482ZJDOv3xaSUiKXe/CDztgKa4BOTGol3brpivFbU3iVPB25IxCvA
eIcihPG/Y1Gey7eZOhGa3h35lU/EZo/PGyijSY75Sm5PkhlwuUqpakjuIirLmQ+X
wanlUqeGFqioypdFMN8WzYYdCoB9uCPKbRhDBTu+cuDnhYyc+4tXvjIBbsJeIS3n
UCQE4Q3PMRgAB2LtehlQqLxpI55MTgjX07FLMw07Xq5RNM9U89GBpSYmp1EIOwtq
XX9wkI58GJZdHJTuIa2tLn0CMuN7M61+ojVA+5l42f+g2/BBKwGR3BsFDqtzOZmN
W6ng+rE19KI5C3bfTt/FKW46hizzxP52Gr+VRhD/RAuQiDoLp+52LU4+FHZTx4Ft
3oIn4kgt0s7waIe6K3/GC05NBwlTXCff45NBPXnmtFm4nj5xCVdhjZWkvi+JvmgM
dVlOZkLtO503bUsEmYdXry57XGzJpWpx058/X5GGSPFO8d1wVhixTR77YQBHTLvw
6VvrTdP6kqVKLKS7J79OmJ7LUbnkXPuHb7mnRkg30nBVPixZqalhc91yqiW7R+1+
tMJMgZcBJmqYdHhtE/FPH/3yrg2E53QIEgFmhqd/Gx1vAqrV/O9aPfyc1dJ+l0x/
qiasRHywgxT+qH+fLehlTL+U4TWUJ2dY800RIxx9R0jsWS/EKb0ZskgmQMSEGDDX
EnTVRDiZkbwWmaXfYnuw2KlQ8bsLRQFcpTUQFYYHPJVIjv0BPbdJ/1ZV8kqHDfM8
ucMstBG5zsdCm5UJjNboIEJjPy11QgVGxlnlR6u/iSO07rfFfV2rRjQ28ZalIKFr
tufH/6JRxRcpuLGI7nrssIKb8czfU/xn5N2bM5jEd5/esbe0DjngIE5gg5p4H2S1
l+KX0IO+XHaAEGDce77A/oSIlbCV6JusNixJ3P3db9jm3xXJ7mgkLU9Gbn+d7Xvo
VcU8e91hT5I557arcbhgJfEXpa4pIl/iYdk9EupZPYSX9zZo/EJyIYCm22FKjC9u
IuWbBbWXdFTElIr8GWQaqm96goWxG0dPW3Iva5L5MksUtoX+t+8zUuG2fVCNMxyb
5GyQWtGqPhRlq0dLtjgNTA/KePkTSn0TWQIXuJmKUYLhftRajnmsyYU2OJfCNlst
HkwnWC9LdDY52pJQ404i4Cl8XOPjeXam1upmncFGIyB08ZkhVtaKu7FxyCxaXoUP
HQK7oRVRUtazbP3WQ/bst8nY2vK1M+AGPQqoqdXXMPaVFZQ1qZFnOQS1hwAc/pEQ
1oHXa4P18aiqVmhspaw7BBQXxEEC8UmeGbwj7zzwlyGaKS3rZ6rwXu20tHqWUPDn
j6ITUPqzT/x00e59ZP7e4FW/AvqueW+/gOqA9pfl4G2tYn2om4QGEjoTDYBWLeqk
Q3qegqxpoVQJ+eh9HW5REwoqg5UNjqP3OyMWo3uy64LKOVqpxLg9Of0JTzUtCok1
XX1gqXF6K7Ou40GJ8JPXGE7gy83XMw9SLxM68GNfFAUKDk7xhfScBKfLwtMoooS4
FaghwtmIios7msS7qgp9Wl984LIQoEUINeVUgHW5gOu4KbzznZH6ydyBGvrnodiG
sKNu+E84XdrrhOLwg2flrQQk2VYmiFRPI4Ui8C5M2YvM7LkgBgvTPxGZ2PoNA3gX
fdOXSwSv+lBledNhbaY5J+iQTuj2G/GRUhFbLTANtgGNWHkqIaHXASUktlAuMfth
wtNDF+j6r2C8HVTEcNoxuUFK2uXOSHneL5i+K+qVU1bVXd7jn5L3LMBnSV70izbm
vvdRBIfchoBAVxMv2YARQ998RRBY6kWdMZGYZgwiEjiY4faeLZbMxmvsOUfQn3HG
QwW9aZ0vCIQsJOepdjDVYE9xQ2lTj3wpt+8p2zk8rsK+yGkTssqwSQcqMwT3klnR
gaQkFLheUN/K78J0VCNv6mplTCpU6xig+FxmiE/sTHVbs4TtABARCfstq7x4wRE2
Y8b9xiiXt7cFu9sd1Qek2QVT0faw6xoTLE8rBo2nf861fEjyzA0+/UNR4w6Zwmya
5I4qE4SiGSECF09xzJAUPhi1KW/b/lO8jx84uNlqXUl0acboSe0kSN13El1LgM91
sCeTdrT4V3KcRQcawp18ivVTT2wAtDWNNRwmkkqLbTkCY+esuxYez9zndsh7Aukf
V5GavQz1JGkVOOabM2D7XEiO9EYyfRFCghTsEwnQE6tapv2XFK1oc7HaLMajSj6b
DMYpgeXLmpqfoVusajnv5RvfXoq5TefinD8ZYJo/54PFJf4scvQSsRXfooo06T4d
tNyFbM+hpV4mTCD+L0+5OBiF0O4+nr0Kzf4VEYWyW1gdYlzHz6go4tY0Nc6qqwYh
AhuqKmUQUfFRVveWFzPEHqf1rHLRkANh9hHIXx53ug6diLwOkuYNnZTGKeKEFsOn
jEjjWWakWPXUPws80iS0HqqvpeDMZS8t8nGZrkCZCxsm6hA1HD4Oe9DGtA8IMwRD
unevSWvNIXqKVCr6o7kwnQTP9b61pdRvzGrxDmipiY4MpGoJx3WkvfYNA8gH2eFt
sQssd0pj+dLubSyKiEK2U70PzOo2ZgfsH0quQAo9br2M86vhV/CRmwwEis3iWMuG
SAZ/qW9rUc0jrUSRtRlGk4iEYZ33idGlb36kVnoTnBk88neCqeStjuAvu2D0RT2A
OCjdeaPZmiup+lGSnnzVhcl75lGxvYSIeA+QopML9N7NCE7cbrsgOZW5dzTEwMsQ
FQfhF3BpFMe22oldo5hhkWuxYjP5uFzLLuD/0zRgwPwVR3vsyPSofIxrv0FxIYgL
LllPCDqe5q5zrOrnYZS+/wXAa/YlKK6cGmp3Rp75Q69utnBHQwKzAqT8HrvNAb0B
cnveFzzvoedQdnS6glegt7H+m6FFiQUFAwCkk9Ev7yMACnhoKO0k4TV0lH+nf/rD
o4ExvvVxJivsF3NSxH5w/6C6qnK7WRRwgA8gKQRAXi+3nwZcwk9G4f+Na4BISxNE
uei2gnOYuoguTZ6L26bU9a8odwji8t6hjqJB1UzOJxGaYAu7iLNejlzSVo2AgaM3
M36g+dHy2MK65S6Xk4LEaDpCeRp0trnZr/W4p9pxFnLg7ZIyNPaxBnk7hSHEP+RY
ScWfRJtnYcRd56OjCdMThFC4ULNpWdqHhYlHocSFALv0PYE+YoewBSd6d+Qpz3rb
UWK/wboiJrus66CjHE9s161JOgvgQvtqIdTjPHho+lzmQk+mVVJ78bs0rhe5jbNG
mJZuioajbqX0kcInavVutIr+SfMBAufa0dIBfvsVJD8kdUpyli6csXeBacOeaVop
ihKzIbx7KkWJ1MyBP3BwzqN/35pzuHQ0TOiZlGmiItejbC/dpgiM023EJxvz4ckx
f13D1+iW12N5jb+KGtz+cZ5DOh7W8eZiGW+J4fm/081vhqlhfPz4FUgQSMq2KN0r
to8U6A9BjefqG9p3wuR3gT3/5UYJ0cH5oei3sA/7B8pHBvu2N86IAUrbcVy2HNVs
tWU7tUxqV8CdRJO5xwuFeB5KACyC5nfVsR46fze1emR1U4bYB0Lg50TR0pvWnZaS
lPNlE/flKlq7nRnKwIuX/ONreG/P6K8Xb9DYvG7ajGJgRWbpjc/+zV5gywwUy7YK
RELJxwbTwg9kq25IYmDDhvky5oOQN5uAA68HbQV3zaYnB08Of0saRl5A1ZVR5CVH
xX8S7rUgoinAjU5mOHMovkywIVv07QcNW7yMnfcEVhLyr4h+UlmTy1D6fpjzU1O1
ynM4zjJ1FUG9z2q03gJYUl2aw0nYZPLda1ePwHS/Go3fqpXjxFDf/3GekrV5Q+Fr
5TpXZiZ7Cwe5P+44ZwTc/4iRilxmSyZgFBSnc4rN79oB69Eb/8kuorfaU8LkMohh
jqy11BwRtM5xP9FGTldD6jyk2chuXBJrY9mAxzkvfEfkjqhS5OGPfCOg8BoKyTKw
vHpXxODGzRirUC7zETas1DFXriHRKCdkmdiHLBzUspo5OJoMyghMSo/6y4WAfyPU
zEBZ2CKR6z6N33T4X0jFbpTvXK1cAQLra90Zjj/CRbkex+AOpNRoS1OIK7gvOv2J
DindtwH6DdiUhZsXG172ar2PYjSZO8x56aTs0g18DUKF64HndyexUOHvLoORx8Oi
WfLJYynwvRUTUscpz+LPQo4VZa3YgRM8lCyc0py5FDtj3yaYTGAqEnooi+2MNcAB
okCoSzKScus/s7B5VjLl8ePhUu2ZF1qw35PdQuHZaebIDkLwJez/dbZ4x2yCNRy1
S8FEaJWktNeGZXE7Cp59IBDWKQGVb2g9QX9DIJgrrjDOaK90z6zPf1kjJ4b176E1
ZSvk2XP9oHQDT30B6VNnHj9oxugTxbGLaHoNnJjBrS2zXP6u5dJ71HFmwTnDeilV
obUAGUXxA2rEpJb4PBNF39JgjUH+GaN3wIOR6VoxV6xh0bDRCoUhIHezfRKtV25G
z5ZvGTJW7yNz69S0L3n/bJns678aZTeNdebqiXK9vqaiVYUWM4Ip0bFXTcU5NyuG
Z2bhKimWuXfFJsD0/pLZ8gV4/MCyVImUU1756pHsSyVJ+uTCTQw7r5ZeOBi3VZl2
RDXtyDtGebvLLlVwRp5ArRTHiFZseT2rH9rIw2F1o/cl1RzY0BzmQGXfTgaRF2gh
M+43F9lkYVjEzn1JBWjVoyrrxSkqDPchKO6/ODLHVSKFAEYKHkOjrMrhu4VNFYq0
NG44Ofd0UJ6j7gH74rmFVSRLFyzEp39jqDSeXao7n2xj4n59ZLW9Ui/dPvJclFs0
ogjd503X7PHGxSSYqBa06v3BdWRTrWt1FNuZjI8hfaLN6LttBhHC/Gc7ocWXB/YI
03DnzdtYmhfXP2rD17Ub5Y38eDpIG8k63ZnS+XSCbLSNwkWqvbacMNF7pwxpQQY2
+McFqRwbP/ubC5MoBvlZmhbhrq5HDPWVZzUTRSl9ruAJXHA7JingbOJpbnx0kgHJ
lrgP66kQxoqQb419T75bdIOBisBB6XaRS1rpcPFkYr6CtuonQjFTzshp3h/pM3aO
8HYVqe20hUgkPK8GHv//IWRqiwcl8NoB0JZX0fXqSx2r3xO6xXNbhvk3hEI14iCf
wV7wRmPVgbHzGV2LWIKeduKlC4C08IYfZYjSDAwEES8ayFxTuUnw/2GrgO/HHj5W
JgTRqXx7Mry7T2IU3MU2crgIVjFShhxJdYC7Tk8LBTjcKsuUbG/O5xVKhR/+NfLN
4Kx0qEcsS+0tOq3Ujju7BfF2HNg/wb/XQ5pk9H8XcODe+EKizDBQpJoj25JoBgVC
eFgLkdxuGNzsLmRabNCXnm1HP9g4Pz4/a8TsZX6NEAQGYZTHqkR7HITAaklJMreV
V2QKIcFPafy7YqQZM7jZRdBc1wD5txx3fw9Tc9HoCLjuoLa+ox2gnu5irQJF26Ip
1cAkHxeeHBsNlkyRwOAwC88smE71a/4KgcVq5mfBV/KidIKDoxPR+M2mG1EvDgqI
lDWQ1QuZYiAVoErtFjY1akwEfZ2ruPM2+YAm6eXLPqgutgyTtsoA6kOy+Qbgzpzv
I+GYze8PX8vyF1Y7E20wFHsfpvd31L4K97Oz/OdvTn6KQnoFhjzQlNB5UFX4mRRm
9exRMe9efR+UGWs6s7BxBF+K/ZDvFjCYUnNRlgFHjsbIcbxJ/3FLHAR2kSjKjpnB
ZSiWJR5Hpw7LxNoIRmkSX/DBKzSXMZWQOskKtaNYBx+A1htH+NRKgR+ubg90jqme
pGWNX6hlM8DZvmcJ8evCgIHp+UxE+c59HwB4RCGPPbu8Q+lTqiotH5HHhagP8zS6
Dmg+GFoRqUSb2gONUJkI+ozcmKlFunmTJyU54VYJzq+tqcoNt/mGYRn7KicaREC0
2VFWWsILZzfYm6f5+QAEnzCG9tRtHqG8FYnTPoEqF6XxHlewYOE9DX+rAJIfJ0A7
INvNiBzuspsX+/UqKFvXBMAjrvBckh7pijpOtgrtLnbLXjrYySGpCQ3w2eHblZM4
kQSeobF62lI+TnZZ/05juXT9cHVDnpaWombAwrJsrotls6snkj0WOhd8GrcItPJm
i6SReknblyKm877TSfyhWnbUZgPsFzYOBMtzcTj93mO7ysSMymnCnDCkpUPMAmM6
Yo7uxW7tHKM2JO3RegJmscKozU2cNR+ZT91QalapaL2qOCb+uIoYRyRqsowd4THv
wbuWpU2PmmFssW4LUQ536TJ/gxHJLDEM88Iysu9qr71DWXR7T0ANoA3DmY16Q3Le
8V4zMTNYt7AA2dwS9rdsNfYiGKhCEjyMt5LhXIh23FVoAAKPx7H2evkESLkMlIyc
A83PDRocm5RswogpWdndAJQ0Af+8tdeF87Wb0k5+dRUC7WLG32TGmQn0SY+7FdJY
26zD74rLDI9nrTCf2atWeQFgdwbf0VhXxgNP3KFB3Jz7h+df2j1uYEWMHxUKd4R8
kFgvXVlU0uJcPUyFP0PQtdde4AsRl0tqKB9f9U7rLgX7oMdZ0rf8xO/Dwh/q/471
6YKlctHnVY4IMs8eMCOEjg/TGdgPM8mAZ9Y85+efeO5ufNfvjubEK0nmVZj1VuyM
ZKda3DM/WvgscGrCG/yBK+1I7tMTtnRtRAKeBMVKS5YuV9qFgzzDQZvnO88bv4Zk
LQTsmxQXEJH33vUt+227Co97S685qyZpDOzSrh7CJYSeFL6xTJLV06k7TIcO8juy
0/2j44snFpk8t6MGBayw5ougXNtku7IGbVa9kb9ynDWJlTmBbldsN6Nc4dGQlUNI
2gTocNSfdo1cvws24WaOx7RQRJvXLNy/GfouCTFc5rxbwQ1lXMVINcryOyld/m7x
z1EnsbcyNf8Nk9T5UOvqjZhSEYi8WsBBWCsR/OHngOZqBnHkjuCzmBfAV+5IRlUu
OP7XIO5/EdsCJj1IrucnDY7/tYrsPMQ5V15Z4Aa4wuFKaS6rY6moxdg7uyu2lNp5
Jrle0kXuaUKY9IHtTzBap4tXmQ7WKD7kUtz1X1U3aazyggpIXq8QEwzT6cs9bRiA
UUSEOr9mJMU6RMpWFgCqG+Af6a2p/VLkxoLbTdn9z61CdFjZ4cWj3aqL0NlqFlbv
LTiWZOrS/5rDQQjKthVM02Lhj+894g78wDTZaHgctCPqJy+9LXOvbXP3kuHDDLV6
VfK2k+hd5keaPUvN2hMOllxJNkkZnQa2kh/QWUHR3ghWYvOg4iVAOdg2SGCGGlaA
xUrWxJlc/RAXOfTFrMXhfmyjX1sUTmC3Nx0bmmrQByCYQea5HKyUBWGIYVFM5Scx
EN4J5V8EAllRSq+k5qelxlcexXxqpsX5V9NMRmvtnHd9ZOQqfGNoFMTq4Y0W47/7
LaVEJHV/VGqpTl2e/n0aH+88Qx9LwCpn6ozGJxBkW0KEB0rejFOTxSHmlh+oY8Gk
/phzHQob1HOOwgcZBLYLmmWWTH7skFQgvwr3WB1wyOXGO0iy5gc5sz/uemZSaKv5
KEqJv2PsUl5i0idaPhuqrWALx6kzUpWcSShDsX/9Ob+CmQn0Gc46PFZec2df8RIJ
9RssQjJSWqyClEBp2gWfTv1AE6tYkfdXtsyKdtTXqUG6oSg7+GtJmp6KLZ0LB2n0
YZ8LaSCOhUY/n8lZALBDc0B9wNfbgoM8lyKJXCLBeBxD3irT8TryxMuARO8hAW9p
33IHQpfxitiGsopmtA+xS/xKqM47VoZ0Q3uNOoe5UNBUCQJ7PRyZ5DXNq+ZZF+y1
/rxqt3OG9a6W5ulp1zT+5v1z/u4ewc/6IMLi3YPOBSiVT+BO7PC4DWoBJhNKUTKn
OTZaJqVyj1iV8KsS3JUg1PgFE7CzRKdiYpU5Ci5QhLzCp6V0K8qsm9SQYWUaA8lO
gx24A0HRUMmaGyLL5TAMHjS5hTT7D7ETW/jWBpADaHizlrs73D7wHYxQvfFmiF2e
+d9GWLz99FuWclBBRBU/j/tsFK+0fV3w9X64vDq2sN9ACif03UMpxi1Nlhduh4hY
OzKkK208zZgZIufRpHmPBPnxu2X0PQjv4V1TTTnb3UP+5dlzRUIMjrvDTgtS//1X
U4qvU2iYuWdoUF0zIHWUWhzRH+7NDF2Md2jV+YyMdtooXRVUB+swz03b6u3mPz54
OzF5nK8FLXE3icCuH3KCRJsoV5+/uY/b00Poi7TXxYw/auTbtVRu9U/VMTHrkzV+
+RKFnizxHnRZnnoiu5p6xVtqJiwkl15x99977jDFKEb6gZ118UiBVPnQkz54uIt/
nbCvpj6DWk24CSrsdEomqo2O2Fc1wmBBDhf5DNcUiWHZhhDYLzP4OLxW04s5RpVH
9THMVkw2Zdv4KI1FPbwnfkyPKM+tsmndloyR4WWgLmkOzfpjbEwDaBbi6BexxQmG
+VEEkjC7O6fuTOsfBQkR7MiRWPRxtcfMTKxyqAl0P8S0Ez+Sp/P2AIiKnWUj8hN0
HpnASLzihLmI4/6rCbT8TtsLaAVWuwVRftTZ9TCsOAipEALpqSlvKj/sCcDJ/YNs
KUdm3A2/d4l1AwsuGk2cWeYGOx3q9Dr3rKz1g/fuTp2utawHJX6PyEAxzVTCmHd5
dD4S/07DYUDE7tAzhcTwlkSTjCTSCuGNYn28Fr0Xx2byn+fPRhLWAflrLtB6oxgT
xBTypkJWp6Qw9SWIOjH9JYf2x0uTmDsqn7c1E6Z+QFdmcMu5I5EiTnbzZEhHNful
5vdONm7jBTaiA+8kJvqNA1MoCTMaKhLLsv8AkJAXQiqh0D7o4VukVipsFJeuuaZR
P+35dnhH1Oisv1XgQglW5I9nBzIugC5AfsXWFp9S2p0KfsF/+MjARSFguqtRjfVQ
jiphrvCgcb8PcVts/F9xvLiw0oTt8bDBVynkpYk6cgglF2jnV6CuqKPprBprIjb3
1wYZD/IjOdyLZw0R5CPhV7sPXWiLUWw9MYG6UqN41G+gkBYErnfISYjozUz9MI4W
VJ6KYQJxXq5SUg9pt0PzCMk/isP3mo9HZdnOhulUoH+iwYLU65LR+a0JYxn5WJt3
W5Em1zxkXWpAFcTSyWHBCQSeg4uODhPYGM28VC48jVkoh4DflxPN4aN9kslOr1+3
QvPVh2ACrEEoUZ9lo/UV52NXbMEfM2EWb9vQ+hd1ZkkHh270JfFsfBLe05kzKoPI
jl7fbUWOJLNP3q3X+GG89Wd3uTOmXGYBoFyvH/uczE8R5j/FDB7y+XFxIGt76Wn3
dMslKjqAB2ou7AjAF3aK/KHh50UBADXaAFJV6B9CXbiYzLVThpu5pRhpWuAksV5H
qfUqnHLZnbz+uTjCDh38QWNlOImapuufYeI8uL5bUBpsyhE5c/k/OPhL6L1h1QNf
R0km2Hnu1rR+MkJTBur4MnTODIqWSiB5pls3aQq/+a69R8a/vO87BnZvuiv5n/LK
/fxrwrb9373y2IhaQsvNpgVTQ8WU+JiB/C1KWcZFNl/w/+kBsDrePIlWT154qMsh
rV3ETSj87oHvvbwOMa1fiPq6x8O9ChSAY9UJjJTUnETp0ss89uUs2ud4d8SNWYAj
uwqSu9i9mxfT2nDoK6jMrm5oo6YOESaznarf4fOIQJGjyeun5sKH9CXRXXl5ua5Y
eeWAP6sMzzSfNEKW7E2vxZr6h0nyxtHy3lkC3Rkvg7TMUw1EZYWRPTFf46N+bZRP
cyB3rSA/yO/7FZv8butdOfNRpBjq+4pG6X8wz+bUlta9DcXGIk/wYPVhUUiJKbTP
kNYO4eRSAWmH9STg3skIZi5t21vE3PLa+zKckrIQLlRKJhYzH8sBD64QXn1KaPSL
a+PM0qUxv+H0LLfNf2IKxJqV8AAqpw6PKgngHFb9vlMShTPNQ7E79k1z8c2nqxvY
rmCVgPfTMp0mxw53YPcRKRe9demXt8WvOnQI2WFsMD37XfkT6FWtdIERgBRAIM6C
8/Q6F0s0JVJ9UVONvHawaAU0KHGyQ8KBt/p/SX6xY63ACGxkSryKTrAsEpP4Xmni
LUJJQauACgi+1NuKBIB+AbZQUTOXWP3F6lT6Aw+0l3CKA/dZByaUHE4IUR9/4T7N
xOlhrLAImWly0hWBph7KcX4y3Vd+SU6fmfHMxMfQ8u1urzbUFfgX7uD2Jd9fqKNN
19C55Cfrd+sEftO8ISYBgBnfRFvavrOHwQkDkCO8x6jBVA3w+h0fdwzyDQBX9Zq0
mRb/oL8MX/5hU/MxZTLj8pLHtc+W4IEyCk3AQGLWBQM/CIOl2AX9kPZTOpoiLXyg
Yj9jimI/YWtxyTWRzdJz9Gms2fcdKzUNIdWQH6TrksIVgtzNByMdS+VX2KqbklxZ
8kkNLh9LKnnY/D917CaTkTKqLdLyrZZZs7ErxtXeLZCq5caEuQEzwowqip2+nsNW
GJlutVny6y5PBzeEX2hd7GRBE8cWqz7hWsRGug/0/+/sE9LlL/Y92uLsAkr8tLIH
Llf4jEkrVUcyHR0rcwxG1qzbrdMPs06dA+ii2EQ9p/joRAiX2rksnEQt34sdo1rQ
RN5yLVuvRVUaChsKEunTCDRAbD4ElBrFsj2OM36ETX3z/++s//WeZImwtKF39xoJ
6a7VBeFxmb6DlFasb5eXQnWocTjyt1M2c9rRBEYSGK+kUhqHMUnkM/ZhVRiBQimz
SlwjUYTU/YuXGLPfMKm6ZhFUYqnvQHQUhoBg7aKugF88jQir3aux+/YHihxfIrkY
ok4dFkYUT/wyvd41XwBidRCFrpHAbzTZfJ/sEnZeSAzv9qzojN0B+ecmiLklpz2z
hGd6L6jyB4uyEfXnk4tvAoySFCpQ6kXXAd0eL5bdqBiOF1N4Yqd/dKUzFWbla3pA
JcpmgC9FImxlRnH7PvWXELVruI5dz8cmOC9Foj+NQcf+HNUIgaTcfZDitAMbJD1p
CM7p47k2r7gTlkKStWKZqJ2kDCC2I+tql40iVwMYEgZAp3UpD3WVvyukKUSdGgCf
m0vL03h3XRNslqcjXfpvWNOQf5SxYMtJY7sQ1vlVMM3nY19J/tbtvGfpjJq6IxyS
pvtwb9ccDWoH5ezkReTNvPqoSIfD3k+HWBnjJhtksNGIyVeTGw0apgb3CHWFhgkd
uXSG5D3/ra33299aZdYQ3+rgBlH3/+VyQjWJnXnQLWsLVSzHzpfYjLm6F0HTqQFV
fSSU7qNV8HFOnwW6pi+jGXAMLYeK05LV6Okky3s/H+pvsE8L+/o71msX1vbCf2tz
HqXn5t1wOG5QglwTt5B4qGpxo6U5reSu9UyFDgG08n0Zfv0ouHAXvcbcYWA/noxE
2UmA5c89fDGNGoiw/zECT9Tum8KHGtgvrOZRmU7fyYJXOXmTpkpsXUhCyRWh+aoT
okfXQWcZgr2QI/nQeMKGNXpbKAHDl/q6jFBnsBuQZpaAYaJcZ0L8HEY5Ko7krIpP
tB4iu5T3wLXL57iaHUkq9NETFqi6k1ogYT1n+Nhjwuge91qngw7o4EJ7WBhUQFq8
L5NSpc0SoyQPuZpprTjM7wijHeIT+rIqnjhR23/Td2hzwFb/v00EoGLymG6+t6fh
QSbiqfsAZwOYwuXLofg4USeRNH4LR4hV0RiQTAsLyOLnL3RI9Mg/nRrExotEwBCl
SqSwK7Az6u1WUQORgRF88RTCMKXFy8/6rjckkpRvnuTEryu+Bx3nNTVElAht/gCU
4zWFei9KknbMqqsWuGLtQKWjmuf1Gh2f8WpSulvQS81bC9CcoggjGVRW5wPKfh+o
jzKrPZMejKZZsWh16PeqaLdD4rMGiMn5V69OwjaCNtRsppQp8d8qLdIB8Y4kfzmj
uhrYkvCrUNhqogPHsNdWUif/WlFXFHiFlHebbRvrixb6XXG0lWgtufyCdyWidbBM
7biy4FPm9Bp1AeN11jteRyAXugTwpCetfJnSmtSDf9jrsQDTU1EqAxx4uTF7dcKT
fp7Nf0AW0F9vd/hcAtjMZHIOON+EsjiKE1KP4A5JqIA/11XVMYSUuLVOGaMvh75w
WacvhZkS229gO0n9v2IXxXJvf+UO7VqCQVWtacl49bvA3RzWS+fgWKx7BIMUg9hB
nCVpYwGUHysOiH2G0NE9R+YpsDPyWlaX1cZaEo/sOf/STpWqn2jzINjmwS6dRmQX
PrRAefv501xvA0UrpTIGjkRqAdxCXyQ8eKRwJXYmcOQut+oC4IN7fG/5Pu/gL3Pz
jwlDHtdlLusDlRzHPHUYCoueIg2eTnSwB5XAmip3u7SCMnT03GLlN+KAMf7czpdL
XMM8ydqkto24MK/rlWwwrOxpgwlFsc+mTq7Z+I+KRRLXH6picKQ0VDM+FAlFfACu
AdfupIrodPSMg1HYklQ9pZ/lbG+/rB7UCr5gIWhONOdiZhDchWtQMc0/Kz2TKi9W
YOkY5dTNniUjBfMdM9lMmuhrnMnNhKcsgw42V29oJ0Zx9qJyz6iyoFgvk6zK6Jcy
DLA7fprZ3RjU2BXrMx9Ozp/MPBRQNXq3RTxBkz3n4fxiIWJl6iPxvfoyp5iwwIP+
tlBO0laKE/WE/wHHYolWG/+Q2aA+TtL1CXZWtRXpLF4//PpMwTykB3QAGJlx4Khj
n5rx8BE8PKmsggrJQbSC2J5091x/5XGaIBE4rA6zm7YlU2EnFlK/8reBQjBFUy5c
eOVoOSEnAH3/0oALtwA8OhmEt/WClskmRgYGdTs+s+xeBv/P6gEfCbZmnqcsgHBW
n7Hw+9H+YcX4Pvgqsgg1NC7B0V3Ds30+vh+QNmUYP68Zvhzt3moiO3+ZmXRwBnzE
hyvWJUp773s6CyjCPLVX2eML6b8wC462xU43PMWPr45ssjNae9S41FGoilwhRmKa
XsVdqQXW7fbJd9NQMMKQ+HOadZYYKyDlw9oiHxWvWY5SdStbGDN9XMd4yeqF7KFw
HsPaR2406plckebZQsgvmIlzDRhXivW+i0/serY8OtzKYRAM+pYHia252+vQtMIe
u8U8TMUw7RKTvc5oSOyXK3UqZpsWihy++D3xd6jwa+oMqHeb/PyWcnrfdoSMKX+J
tayTvQ4m1kRfKjGCMzTsD4VM7TOYqJe165FIQlvRzOsnle1oFXrhPNx8vnBi/bEc
Vpmjp9Ua2uBgieoKs0ofaZGcOC4l1LGkdEimUN1jQWStN5SbR2qRUTEwZHhNNoWV
HPdN8koPAMZdFhSWayJGvpjAu+OTNT/PZtDakHvFyQIgoGmd5kQq7rOzsWHzGG9J
9fLj2nF3kY+P8OLGOLfN2NerHS59EaDqhTNUjIat0eE9F8isKyFZj9/PXDq594EY
D8Ay7yqMVhT6cT90snPsclzvz/7yY3cSgg4v3Jxz077sRYc+WU173+LxRGuzgaML
7SDSOJp/Y5IYr1QQ5nswKgxqjAUAZdDaCvP58zjrvfhHyI0rjxKuXIAK9dFOc1tR
fLqxPkBkNBLuc+l3ircdCnev0/lp4q9XhELYOLhpNGNZ8NufL0bR0g8RQ5bB3Pv8
of2pB+47oj5I/Km9ACJhoVSz+XQaX+UlM9UZwKJWmPIoaF3GBjJwh4M3BtgJrp45
T7OZ7uwA9/a871OwEvitlf0DPotetHPCiFQgnUyB0TXUNZ3Kr0kXqDHWd07rEhut
F8mykCsy4fbu5IYF+hWAyAZ1mKo8cCLf6q8MTKlTB/WdksEQeH0e1SmMNvMQDNuy
YUiaHYlbLeCvmBPW1Cy5CuXAWXgBfCIi+pFX45tBpV/NeX/R/akLi3GkW7I/r9Qu
ySxfpsPJEWKGGKdsV3H4b3OcC/4TiaRgDP4t7YiJLA7YAEeRdSxaUI4CHM6uMziv
57R37duQW7TZ4i57U7TyuZKUeGgzK3QzE5e9IjYpSaAHASGZ4QjNRWYJn34UoCsy
lestvTHWaDvo45L4sFedwMmH0i8R/yZKkkGVJpvs9Iq1gRPfty2EYZf3AiNjSK9r
EXIRL15QfEwseONyfffZHz+e7/kWiKfxUrHb0xW3oYCZmEfbt3p7Rj1MD++Yy5UT
knYtpyiQu4Q42byG3v8Bha1KtNQOVW0XnrhFgSG1Qud8iDt0lSQcK+arcawPlJ+p
xWpSmkdo9+eqnBNzUetT0rTHC0llexwypEPcoclD1P9ymavbt//6SO04SvhSxkxv
NbRLi0SuE0znNjYR9fOKbBkUe/KHOKHOkNDvNRARU4GOVtgW2Fav246Gr1wnZZfl
ohsSvLYdCfnp+lhri6yWi8hEowZdYm8UAHySqIt6Db5uMSKd1g5vPXYzX2/tsMqJ
FuucOrPt0k6kOCgKMXWh7jrGZBkLgauaLdVGER90yqJHGE/CNep5PvbTrkeBq6Zx
KQOU4qC88wN2LUvHT+3yQ5CgnBQV18Ek3JDfB8ORn+W1mQ9gGrfzXi8fpu6S+voc
CBxQ9+0Tz2RyqbDKYrKnslYXMpj4jl67OM2pmEcC9IZowG8Zrrghsynp66isxpbr
20C/mjTl9SJ4zyGUfX9dy5nyCe94D/1UbEU8VR+p21LctPyEv78fjHxqtFqJtWXJ
8Vhtitwd6EMt7BrJTlmeEYHtBbo1kVqN/h3+23OcXiE23X0bvc+5BOLOe6lbZ0Cf
jV3XTWZ++bj05cI4oBRiZEo9kDYdaMzOFu9Pu/uLKICZa9HrUxVyGsZqvh4pkzIw
Rm8KVgMdiUrWkeoYHaRiLXSPpS13JHQuL64U919lc7LHNRriWINawok3wYp+vFVk
/L/mFw4ARfL5rIKzb9YVFCmAlVZCHlrsCfDwsLZYCFntODEDAoyTSJXkuwJc5fQU
39AXPVL6PJllNoJyF1w9M0lxufzefK5PDK/+G7pvnSQi797bdjuMCxcw5ZCTBJaw
RiYgNPc9HWoWNmwIncroCgjkAriH52j+kxIUTv47ZGJdQbqR7dTS5AgGgGSXWOwW
O3R8wM82985AypXrbaOuiewVD1EbR5VaPuQxUvqCvXOAv60fZ2GQDAryMlGYhBdH
dh/EkrwNkFcq4esdEmGkWVqOfUgQd4TgezJqIg2t/CA641Zh904XfiwpsD4hHlts
ZWpWlNwKTWXEd/Zo9cBtK6Td6UT/ED5zVdkDrfrWXt8ykhOdFot+KNseqB7W9kGZ
q+GMJ5Vj0IuWda9xYxzFDIYVY9s6JXJ5a/5CxPoswaTsIi1xAyFgYfbQhsN/Alhy
8P/JMLkKQO97VQFNKxXcOX1mEwxs8UIYzq2M334rJtGKptrHVFrSI223Ri4Odaa+
2YyCpQDzhJ+FRD1OlgaQ23EeOdAnfzq7CD76iz+4gK7ogl++8FeAL9qg5s3AQVE1
tYtEZUIu3cZS1pdr/77gV/lluhjd9gU3N5q4FGWS6ZQCOHoikfmqnocOovpFexGd
ufSWLciTYwblKkS7JMy0cfsLmtFZXp+sG46LhJeyw1W/gPqY5UsyRUAnjTlX3nGS
S/d1vUKWqZubHd1YpSdJfc4f5EgYrDPpm46CjBdEki0Ly+VPWtrsbL317CEB5Cre
TgVswq3ycxr33W10/8qi1l02+ATU54yugBe2yBzObFMXV7L7fgJW2B4GrMmrAt16
EQJXgbPSttY4KA1JhAlx0GN5+fV7ciqT+ERvNImqIzm6oqyh4u7GEduvSOJQLzxy
JBoJE40KI1YoWk7wp0OSsBLOfGSJ9Q31UiHYjfXX/c3D4EG3VGj4pVDUmaYN5bdm
/WI0NpFbsF6ng9YVvsWN+eSj8eKJ8KMd8SArMLIpB151gPJtILhXtP8CVY5kqS3Y
rvdOxUnZParyzb46n5iGHTT3y2QoMAfPIsbAqdrgcptvoG5ELy5uUVkNkfJWpsVS
tChymvw3rY/3RrSGnMyfIVB0H/Gu3jKZKgrWMFB0g0a2wcUBP4+YFOFxyugSetPE
tIMDDBbFDfqvtypRWG167mDb+xFNfDp5LRuG6g4nhN0kkVsxjasD5CoTXZCPKMBx
WC/F5cjotiu4aDhrCiq+Xv2AaMZXDEEGAuW+CSbQo06HlfRDOFjILLbf8hPEFYOf
rvq9DjOFH2RHqRXnxgdvjJS6KypCGXhwzImK/fL/4x8u2TuI2Gydk9k8QrbxqPlg
9FNfu6xRY1BufjGk3QmpnqFZ7KpTUzs+0Q3f1CNJSYX6tUrChtXAPUXMAoI8FdRK
9FG0qLO3GGRQ9fkogDDSfJPExLNEgg9fAyk8TsBigAWDeS2VH8lFVIaN7rSdS1QC
K0e0V8fEGm45rKbig/417FGLj6akPuLlKqzsibsPLHSOewovpQoMVQjKPGlni089
SmhOOG//MuPFRWWbh+O9DWy+fCPFHUHHJMNfWO59MI3DcYYcZPn2lLZm406/b4tz
U5Jm1IlhbMwYEv5WIjV0dIDxpwSAG3PAUK6ONEUP0fBNtL7QhLPV7bhFIBC+Nhz+
eOPtGu4DVXe6QtLGReO6sSL/t7ra+gopk/OGhmQzm+2wSWMg9GNKjY3q/x5KqmVy
FxPB1WKZ2dlXp5xkodh0zLVL3pXzhLLbNQ4CoT/5sWAGo5LqguWYmUJryzLp6kTN
lRWr07Q6RXg7XZhGVXRW4QN6yI00FKvfR+s1pJn7wOYcyxzkkRVnbFdkUaq9AZCu
jTaJLRy4pR1mQhTljUTmtgw7jPPflhEcRj3D+QT601I9Am9z/53rvvZUIoi83eoA
ZkuuqLgvLsXMIVlDHvd+iJTIXCD2aOgKRYcRX/EmKfCgybTea4hL0dk3JLNi8jXt
lFyGHMxCSTrJp/4vPVfez5wmu1AVLfdexMI95PPAflc0nWX5+eRLdbFu2iU1dyU7
RlScAqNFZ2hI0tnLOADJU0ZNk93zpyvf14Vb+NcAWhrCTnYPGHJjPOaJKot7kzgO
vanaBs+M1c/On/kfFie5UwnHt7HPznTeXlon/YCNpgb6wgKBALjQYKZ9Gtr2ztku
pOrtWnzAhT6ECTX/7t9oBfZcEK/DLj0DQWJihV5gTm/DoXQJ9EnP/0DvGbIEy630
bCXFSM5G6kiyRfRZYD0fmDNbnXp3JxSenTsfRMz+YPvTMyGkyjWFqWVT0inn+3P7
0925ET9rLsLvtm2wIOx2UbcaLBtnF6VBYzz6YDT9vh9mBk2K57DjnI+4vhQaWS/G
w9/o6PAY2oSC+TZQe8qCEdoKNHKT1nBaBIMv18pRYsJpqSZBUtttGEw1PJa1FHlK
S1co4AwevcWoeeyoKuL9vOzvKO3UH+Rus/zcIEzciwhzu/sYsR5FVVxpWOgzvvZC
0oIYPcs3yLIufzKvUhKM3XN4oeTT0BBFw7hi9kr0bjqs/8OsVjnvUEsbdCjvVpIo
cxvIJVVxFC0nFoE6+M9HgcikI03yJu3g1x9V761b1BV4cvs6Ar97q+Kt9zh4xguW
KDvMLVq6ttG+DxjvKFx7VSo3Q+8vGrTe+s6lxKK2aEEcvfFI/mszohY6mq7/aP+t
bmhJeeO77Fu94TvFsQ5HwV6ZTFE5+j2mcWcIMr5iV/ODUJNGf+h8Hnw/PV9SYfs5
2mCn3P0Oz9aGemVBQZpZwBA3DTncN+nt+y+jF7GWP2X7e42vgfUH68iUK/wsurcq
6KUJK6BJ7xUNEevgP0aSEKZnRSTswciIIO7Rb4ctbXWE51N9vhXnTeY1Sxd89bBa
iDIGUUE9BJwiTZJb+A/U30bIojzPlVAkN0O7JfX8F0GI6dDuDjqnJ6AzfBaOIrer
/FhfL2pkGPSbpZAlU4u0Z9+9yCDl9vWS/m3UpSd7g5FQ2Y0OLE0EXHqdpV4DGaIy
Bh+bUeNNrYFRXR3GGt1JIrTJd9ysAZS2avc5plIOnrzy1SgUjbylLjBR2TUdQ9Cr
eddQIGiEumkbybOHO5TnfC/UAqSSNfI+2gYnVdN12IehPLQ+ryLtCXw8+WTpmxWl
+YM2Le5DyB3eV5bboApy7IVvou+3U6tQjJgvSqieOtFOkVTDMICPsNtJZFQFzhwa
ZaSHdSoOsSyAzf5Q7xu4MSHwDq9uuY4NdbyJZfL8tz+TRdu1dJoDvRZHFJ1zMXAr
3P082x+dyMuqY4QLxG96JZm+kaVp+U0DAGWvR7EIZDNtUddgKYIzHL/eeTIjWZeZ
XRdm8JxYoPeNioeDZUDNICHzFD2/GbVnpZ8H5F+dDXODZladNtwkTIMw1nV/TD6b
iKVgrvI2HjtaiELVBoZJcLwQgNfyEi6ZVskHZYwm2GK1UBYDBxmcyGzWOgCPM5l+
fENm+jWR036y0EmocH6gZbCxXhgmLeQVldNZszy0DR04QhkLftkd1/LKD21s/inI
fVUZQ0wssSdjvs5Xw9NSEkfEDOzizboTQ5kcaUgJwxUmZs/iqhYG6uQVSgXlNOYN
HUi1vZE5v1mjHAklLxtIWtmdSVG7bEM17zL2mn9tMNHiztR9JioGEYDuJfccVU7/
re5UARZOfsDq4kKVU8P3NTFjompxQ+3SHZDUE3qpxlaBgq0r6JIffAIjz7AunJe0
MCR2B3AjB1TcO7OVsoacidXUy2+/c2tJbpMrmcvArx93jPgMJCVci4645JHeWs35
WLPcv0FCvEroRCIHrLkvH3jughHS3YTqG/8eu6AyjN5yxmDcUiqG2asfgohcC0Mq
arsu31KvIFhzzLhBtZfld4/QiH8a3l4L2kaA3ugt8hMuDbzpLJNrBHN3alqwqXoX
3kl9FU5cg9ZymhYalB8SJjjy6CnkuB8X/UMayMZMDGS1tGMAQHPT9wQ2iPdIha/+
lW4br4UXlXaWtsMGn/a7G2ZTQ+qAFUySP696XLgkNxL/5EROTWUeiq1gyAS93HXX
yALh3pFh0WOp6gbGGGLvYzZ20W5vERSBx3zzjpsX6kPmHOYS4fN8DmeGd+R3xGZk
K1LgFUPijKLTq0r69zNrs7IfNgTv1Ud2ivFNC4FquGtXtNzqigbsJkypD5z8W3vq
rTx23Qy6FCMHmhPiVyu5+CHWBk4sK9MoyvZGAxgea1hPMGEOZWZ+FavJXrqcAmRs
wIiZSd3cgY49JCHgUPdiQDBU/nBcOnH4V2yupRiOYWSviHcsh6btaYetvONwQqUc
aXcGbNa5ktb+Noja5gC9zWWNZCqA7WvSHN0clH4ncID+U3x3oC9mhUirj5qVUAEm
spGYsE4cGGxu8y8sTE5/I+tDmdT1+wPxK5GLOVZcrznN7Nwj6JV4Tc1lDYGrBe0q
vaorAYtgo68C8iOwiIj0PQofMPH2rzPUgtgYG3ZVPXYbvgtGeWORj2ORO6y0Zcf+
yBom4/vwRTSU7alDcDTSNOUiklVsuTtf7GNdHkdKH/kxyYimkDnUbaba6hxJAWEt
oxYe1HJTUVc7Wq0FCf559ai1HH/D9GR1+l/KWHtfsHKOMwkPhLSx9Hv/sSO3cjgS
T0inRXU/hL/B05Nr61k2sxkUjvien/kV4xigyaf+IbEQD84Nbv7HS18V8wK8+bkT
bOPjAyui23/77sdYVQyQTozGYBghj80Aiaun4pn+enAH1vfBiz4lDEU2Q4VHMG0R
MbKaMvXEEnC2vblcd6sfNwoFJ35YDeSqE33FJOIxhOdX0RmMEoDxKitP4uQ0MnhJ
muawkCOvktvr1yvqMgC1vGMLXwnKSlkIHy2kqpG4ZzyWkEuBHedJRateFJOMcLMJ
WVJ/kmXTI/wUN7c2vU5ZRz2Ea+2sYHo15pqWc0vm144mE4BkXCBbXNG5pMiHcBPY
TYcwvrJ1x7oJVbk8uhBMlpSeqR8g6KzV4znHUKQBVfP8HN83ccVCDtjzwfIJHaSF
PloApbK8r0DFzv0dUAzW5YX+aTQqu9qsvpVz6qULZ4dnGoB2f0Xk1Tx6E5Y/5Jwn
Ss+ZFgFNwGka7TDDnv1zVYnnrq27XNdjXAx3VZc8RtfiOgEtBzknWhYPCb465Pm8
FWkvxmjmHMex9qTk7b0MJ/dHk+ZWxcJlLdau5a7MC5iH7RlJjx+iKC3Zw+kIWHY1
noEh2xq2aE88DcLI/OKKvF2xTVy/QTxHeDrBTuFlN/Xtr29m6S4PcjRjd0ZJ3936
GTsQfa64c1PUQDoxtdlTi3mbiA2iy4JP747UTJSd9IyBJ4450l9TAc9+FIgcOLHV
gRFDaB+ONSSY2VLDIVuvdyz2tA/oupXEfDh4EyrlmQ8wPfeOPPP2E6ONJqgguuDE
QtAybrI9UDh3fZkZzTmnmqmxKdYoza6pGWhXzElM6q0mKWPUjOUetAc1l9tnTE9C
K6wJbMRF+Fx2wldLeCG25PlbDujdkd+ZZlvfK0+BtCjDmwN5x8YbngBNvEjHh8/s
KhAMSbXyIr9zKw3q3uzC8IO3J9efIPAdbzIughQZVzirfO4PV3zkmv4XKZbYKePc
YL28sA7uIYtjZ/hzJvhdgmM936L+ddXm/KqAHtPLlp5ZN2ncDvGrE02vyxP8nAs1
oy09QNUo/u2wsU/kEBYQ1Q==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
mld/aEnKvN2/n+d4Ba5C9t/gfO+GBdMLXoN2uJkkBpY5y9rmEqPECFanlVli3ul3
gLKLqJNm9+Qhd6SgkVlIOWtsh7XRE5iKr2YbI/uTUJ6N32oAzxCkrTtW2vSjFd1E
M6PHYkGj/rTDzqC7ymapjgVtTsBIph6/31qVM1bXErTGPoARKHDFEx7fHqs2Kr1a
nUQczTiuETwwPeBu+fv+YZdeeFAgY2zyMgNphIuLifrwV9FeOaJ/XtXrjQ4v7uII
zcdSHBTfEzst5WMYkWxpraWkD5FGQvwPWneDUr1wvY93VzzvTrC7LQTqM/093ryv
6YyfA/2u85kthAk30UMs4Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4672 )
`pragma protect data_block
mdRJ0/G/BhQ5LnE7rg2d4U5A4QtZeQLm/E2SF4IlLLovVk7YueURX1Rh4P+BYz2T
t2rMkCMaObJGb1W6WzZW6U4+69esMDWi0N8/UWvhEgLlUzmjlfd4rjHcGoaPTtK3
LFheB4ljEl9PCwp4k2SQz+tHORzH1Idd/XxOFQUFb+j2gElN+ZsXFhhhbAzxdFgB
6FNZSI8ehL55ibSiI/K8MqwWi5z0hx2btCuVmsoQwu5RCvPLKQ3CWptph7P7Y2QR
mgZC6fM4umL+39Hy4AE9T6J7crKZMlH6S7/7VCC+LfP6HwhcGJU45ZJBLIF+NdJ+
1eLlbJKr/7qQFPRMNnZRzrnKgo7MKeixuGfyvnuAYGl0M79ftVY/tw9/YlGN3SMo
5vrgXZlZW7dnFi44JC0fOBXCNMCdZYhzbWSkVN2h75zkSV7jSSHItHDJcVd7Fspj
yx1uyEelWdZjxWNpdr/DSr9swDgTa/vNhgR8pvdqi8TxoHE33wd3it49CgBhbuSt
+RRZ0kCJmg+hm3GMA5FR/qUtUoX0gF2YfLm/jyuqfPvo7BgLBXS66KkUYQFwc663
j//do9snfZRH3lXCUL6IGRih5Qqo1EfKqjMqTn2ViaIOvgw6p1sgqQbDHDmxRIZ/
VLZtfccvRTi8LIr2CaKdA+xSKOKzZxdmSqXsFDN+wQ7o1xF/cBtyTWoYlx8L21Or
6OLUtdRYdVNX6cpPkmwvcNB9WVaKYGUrcUPq6F1KPVawlNtz3S0Z2MiXdOVLy1u5
Ri3kktTWSkD4EAjYpHdzJpHNYRC4huckExxedYoZo0yJMCgMD5L7S5wZuW9yNCHg
4u7FGMeSH2z6MkGstHiXtqvmoAWav/pT/E14uu4PBMLNSMWD4ts3vVHE6UvJAC9S
yuZtr6FE/q0uLlfp5QLHRIuvSEuYZqV0T3CN75xVDs3SMsp22FITB3AyhO8FFPdz
UTQBhb23DziQNd2XXAfwxBxDb3zbMUD2gM5fgC8qFL/t0AFxqLPq6oeXgBw9CUtb
3TkruzdTlFC6nyDvaXY782kt5AkrkmE98oIIo1ZJaPR7aq56UizQRhpuarlKU2xI
ey686uY4E9v/fUiZa6j39YVNUW2IxkrLSf3QaTrRl8/v+l0lJgRGyByhb3YU7wyu
JCArHrYX0AnMeO4aolUdWIIjhL7x9rAyR3tz+EpKBGCMCZVdioBM23rgO2ed9+mH
qY1S8E/pgPXe/qIxueKrVsmCH7oXPmFEjkIvId00gcuhs1TtiLtCpE3X49q3/7z1
vjRsvXOn/v7fKsJqdRu3mfhoKlYSnyv0nzk10dFpqmSOmDIUVFQn2eCmbgdWm3jp
Eu2nXLikMhA7NVWIgwa7PP44PiFCBACIIbcXXfcge+UJTBAxmMXHlYPp0PGHs6wm
ia8axv+b83tveL7y8uFVZGAjacUPT4xNdR6LNeqj9rUJmIkdancAIRflBvTnHxdb
wrpiB5Mx5I0l85eYwR1kVSTZYeikMj+Goi+RlhuUUMU6WC/k3y0487s0sWDZcR6Q
rrtirYQoKJMSVodce1++9EW/BQfqixZoZM40qPu5DWvke2Yh4o7Eu9blsFgPv1XF
zpAKC+9/ZXk7kEL3xeexd4MGQ89H2R4FGnArl0lhjQHwrP45m4h0Jdn2MK0IxMGK
+AKLSUuoxlG67T4zUQNXv2g1CvQkTPSEOlOV1YXwTsiKrkTH0WWO63IVNnt9ibGF
B5VL5mbnbmPefC+Dv8Ry7blMo07LTo+YV1nb0XdAoTomyzcQ6beihOiY+kTebQMq
VeQdreVLPZTXKxTPUQzG2V0AXbHmsMvYKIE5OmnPpvEbOiLmHUg+vmeNIntnoe+X
maj7OXAMb41lBm/B6CHG4Vb4r/GlXuqyLPOtR4+4Oc9KP0rahdi5ObGyr9E7kfYV
GM1CjBlJ4Tj8+Knx6Uap6nZGgRCD+aC5QcbjHC6QEO6FfyIUjRwMWhne/6HeBw59
OvG36ESbBUHSIdslWed5QS4krzhfvanu35+Q0wYnn/GPR/pXfKMi3us/EJP28nS6
CuD4jY5g43sNLVFV8p/YE4ugFO806qi4vQP5puOJx/+AgvGyHRg03l6s8QG7FYGK
0zWy5wJmBSLePgYDM4RgP9B4D+b3HxOgS3rQZGGl69MV/RWlXN25q6tbTJnnS5Ow
f52cE/JCJ4tDfELUFRCx+RNaY4K8RncvdIi+6PUOnrdXxBJyHfov2++Jbt2e6kwo
aDKHxG9JwJnDqLQZiDHONLMKhCkzj1mi3UfBeJgR7+i3GpKviwuA/N1G48tJDSyS
dkwbfWoOOND01sne/6BKP1eCYSdx5W2C3knnSGGF7vRm2GcbpL/4hAT28QTJ8VtP
60TvQGsM/y/Jsr7GyTyDrofzQjRtBw+LB5hSgIgqJSPDT093xQWmFfDqZVU2N0K1
dKi24MzMeEnd4/yc20Jn6jYgmXOeLPTSxLFWsziybdVXKtOw2vIMEYx038KJ3XcG
5TTAMIdgCV2ZZHRAif7lcBlzohAp5GSbiv+9KekxX02ao11U7Ao18je8WSeM0XB2
Mdzw4/1vRIWJqdBSJkW3X6HFuFa93vJ5/Du69ONwLptR5ModvjFRvIOkqC00JE3Z
fPnpRnZnHwsu4wXNMi7k92JVNv7Ywo3e3QHDDXB3qj7lcwi5uw8Z3NDlOMa8YFgi
e/mBinAEtTZ3NsFkfBLBoSv4rugNhsbOPwJKPBgEjuPS9wQOs4vZFKteZi0AbAau
HSXEJ/SVzQI16+WTh7zCb9m5HQWjVITWShwOkcnrwQrUD8VjGm3FD6PQFlEyNCNy
tyJlc2EYMrKGJ4lATeQ5EA94VOU6QygU5J/C+eCDJSX+ph0rfFwN9VN+veBtQRmL
BtbSJJ3mp3Oi6nCwABEuwSX01p8xWE/3EONrJP81RKKDDBGUW6cJYVHPHTkoN5QW
k3DEds+h6b65gF69pvCq1uOjc6F/Apl6088yBLgBp+20270B0C3Iyj0L6Ak8tZZr
q1zo3tP0H47o66l2AjqPmTxFlJl/+ZBmq82BBBx7QFuLCWVpkgEh2orE3k+tyZYl
r6E/4S2EOMOCAM/9ynSDUDZqdFiIxxHZRmwIKOoXk+wGL5nh9POEw7aPd2osa3c+
CAY7Q6EGLAqQaVOE5q0EzFW/snm4+GXLIpTzJrIEvaXV4XwDAKsUCrnVq7sT0JB6
8Gkw/NdRh6/7vGVf8xJjKG82ng/KltGpM6t7Uw/HzfXC7xNAgA+ZLxN2YmIoNOZN
BKJqWPCfGOMcuUBAeENjxw/wvzuM9Gk9iQkwJoJrKoFqAwrUSQxdKgNSaT7Hrasf
DH+19px9zUZojDX8f/iZZEArK1DiVYv8XQGrvyvISlSD0R5VThOFxrg8Lk7/5+QL
i+R0rUyFjxggCWc2Vi1e//KgMVOhIiMmhXw4fVaYqgbYyUnqxkHEbQXjQ7QqsVyG
XHCsK2+/ayntKg8eB9CVBggBabDCGAphF2PSv+EqHXq6cjQMwZuX/B9feKNrvtqn
WMcSiX44gQMyortR/kXRKf89QyZ/+eaoKATxALaS0RycciG9xB8ykPBcAsWd57i9
q6HJ4x3FNGh1plhQOsbjIbzbZ8jta6g+WHo6KawcauezReBzyJHc+soPbkQoBX4C
ibaxYJ8XUREgUXWfGbWtD8x+paqKgKbjUWSC6Q0pcUCgfJG6HfuNNFbRxqq9Gs/H
w/8pGKG1IHknhCQ5UieEYmQqnxZyqqb7tAb8Ju1ee+zyZKFHS/m6f7Jz3BJV37OL
QLidp+kg7mMObaWQOre35ua35dmoXXrSdo62t2OF3W7p5y1YC1ZDh+bIjvO4m3/4
M+cTSW9NejtQ8xg8tNZfVbxClm7M6Py844No+69h/2ubdan2zEANGzDJnW+3xMVX
g6CTX/n7oRJWgahBEIMXhfOyJpVnWR1Ek+Z6qFUgSvQIYYjhumsqa4lphkbNv+uc
HQaQTlzofTMamwtstm6tDiJz75e84SL7hf15M/d01ruDWILL9Bp1B6G4WsYZP/57
WAg683nGLUNT2Bjn9mshsRMjcAe7vlil/rUJkl8TRHZcTDr87LnVPrKoQfPqf7eF
t3SahkmuC45UyxLhLASewEQMdNkzYMpenXO9lVxJIjXsIRQXQowYEYVedGBwWjgn
NXdAApRib+wcvQgvZEToGA+/zI8g4p0hyE0uNQV5PlEVBsRNHs9otlfn+U+GLn5Y
vpW9BOV1RQyNJXjaRxSzeTxTzdX5J8XVHl/3F0zTHo6SZ/dU8PdgP57pvm4gt9zn
IE9GMFF6LSwPgRhtJVK8Fp7LBGjZtSaQ+laNKPhQgLCVto2fSkNuUup7zBNhoaNr
E4Vb9OBLp53/qtrbmK1XCNcLbPAprVKo81R2POlip0kJIkaRc0VJkOMtGhxw9/Vm
df5DtbEFVhbhrSgT6hY5pWmjFSTChBEfoOqj/nUdtS10A+UEQeGu5H4pvKJrmjXe
4bKfX4JuSq5NOWT5y9iJl6c89Nu5/432FjTpl7QJqbAU6KEY4ilmkvtDzx1FRyPE
Op8kXvpJGVlnP/46iHYIl+sPwOdDcWPAtu1Mrf1edxescBPZSSOpwcE4qUQy9S1V
n1JposUEyuv0d4d/Utv8M2M6yKNKTqFDbba5xWP19uL6sl5QipOCasDG0e8JTPEz
U2MkWqMGK4IImfoHexl5xWhLy66UJ+jOMFAB8P/eMJ31K7N1f0cWNvyrh+INWwkv
loDGgTF1JGSdigDFBhB/9BpDbPQSPimgxw6yyAB1sVSoxWdJ8lRegWwDLLGwEoF5
C2hY6fEodN0iAxGLcPPOsEFZJQObGwK+nyXUraRwi7NtHqrAEbq0RBrMoZuOyCHh
1u4tu2YvhwgHFy4uUDB7hSb7Lmv5mu0scGiWyYzcjLij8ogPsRrlFYgyANxtfM+V
WGEsez3CvsUl2OiDqvtR4uiRzmIdUX1pl2wYWzJtQ3UXaMBCqGgACfiTW7n1DBSo
XQuWmv5oOReLszTrRlO7S/ZhKfqADBa8bMz9Y+Ta/wXwX/zvrtC18Og7yQm2ef2e
ZapG/v98Q9z1e7xX+KqHDA5fV3a3AABv3SWy+5JndM/vhTsr5laoguogGZjJfvhS
3oq1fGGe14x3Is25lqbX/hQ5lUQ4pSLcGV7hQjwWUQvHSVS727x7NO4xbjYZuFnp
NLKpOIV2DdQHthpqgU/CtI6wq2zLbZaMj9eDAPcU3xhirhJwqhKINj561aJwtka6
QvOJDo3tD/kyHsNwv+bBN4nCdeDpVvnY98T0mqZy4u672ysy7wGb0EUtMlYbO46t
rG4kOi+ztLcscnve7iW0WlaDlGSdZSi6HNMA62A8p9ILKmlgaZljLh6N6gamao+3
Q5HilqMqnboFM4Q1wzrz7matOGTebH+HQSXlC9nu7PuZ0DrmnyKf79mYRuUmgckx
4BLRBNsgHV1/t5gyVbqBrATIpT+ynXoujIenqTeZO8DfFIYrdM9Jggk5p8kWS3kt
nYRYEnaHOxFFUNx+bboN2VM/qGHTa1d9psuSGPO4fNvm/VIVgsSHbP28yM1p+bo1
X6rMGFjAlQFWYDJzRB8Kt7mqrXyJhAWjoPpg/PNRjXYX9cJ1FwCIXXjqi0i0Gi9x
ZLRUH3FtU3za8Eu4O3LjGXXjGuB2ZOBcio7NvUGvUDJEiAxwwNYHKSv+vg9ORJZj
CTHoe8sCmeciqLg7K+VEmly5HVTMbA6nOH5j/20E3Lu6P0oZaJeJqoDb71Auap+L
Ch80b6CF4cxKPI2x3xyydVjL52/pHGccnd5LODTjiZJFnQKYiGrToFo1Nq71nlHH
kGsemZ0s5THwZf/1Bq3BRzL5SYI101J8TNapY1MlJEJAtW09V/aHGJEv/X84EP52
RcdoPmThH8k5PbdE6HsENxgjfcqLLyiCGZYmdQBQxuxsrnoIzsjsihZLvQC6P/Oz
ZmRCyHNOw/rF3EenToh+bE3vNcN2U/Xd3jxQnGSOz1qygj0lDQ4+y8DI3I1p9lyj
i5DpoqJKvPd3ndlETpWDDHzal86vtoIhDi0hVlUptX1T6odZZ7Qk5eKTQIConYCB
BySTxaTy+JBfPaSyI6tipYrys4SEwNuKVwgAAMZEjMbgtGsig19IPIS42vhOzTjc
gLk7/re2w5nXW+3E728PDT3WCir3bIt9017ppkgvMXgmnsJDIJRpK7JdIMRiTa0H
VvniT1iybLnsHKCeP2iBYg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UvZaLE5wxJnQywTB1HfurwdJ1FKNJNheBLTtvNgiZehyz/AVGbhOEKJFMsvi2hKX
cXchMmn5MIEAohr+dcc4S7nNN6sa+vWUUQ76Lm5MCh74xP4cGF6ZyeaO1Rr32YQL
9Ehw0q7B/HA/W+t/5f5DVCGzLp53Fs1tItUPIlCt3bHAs+VFLOzxOxlvs816Plgn
3To3mYDLjr434Hb7sn84Ml9sZPi0rfwEUaFt1AW2Jzm6Vg9UqsIBnghNYlTHKFvy
dgjp/fvx3h+blED65HdGoTIlMqvEdwWwCITFrkGas64/Uom6CfFhkm37PKK+SZew
fTPLNp0VdUZuX2CyF8qUZQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9344 )
`pragma protect data_block
0RGGy72iKZ7oQkr9KLk5awACZvO0r4RGozVzwRA0s3v9T/HzqD5WmWCm2AsI/uDN
la6HWMhr1vo8AErpxPDB8k2LBbJRTBz/yVqCccm1/tC8Yd8OJdLJfuCX4lazATB+
m+W1GOreD6gA99Pv9SNGHtivS8LHEwfpw6/7VI30p5JiGYrX4qzldYMtiVSRfikV
etC9q4vToIwES118TxpvlV0tdx8S1IXP7/TOhOQErn3NRqEFY9oqp37z4PhxpMxm
YwWert6q4gKLKdc/Sz36BqQAktMCVNTcQcK+56RWwFsstOwlXAhivFDEE/3CEv4/
I2+a3lSUPzjqE3/ykg1+wg8vVKlOUezJ5ddqL4x4GqHY6oLIAbPy5WvGsr9ggVdi
WpWX4aW3lS2QbzJxt46IcGFfzeuVxXuIhO84RTvdicIo6czTwaV8cqGBJVe5ha24
e74MA24bjOGw5lo26lpJ3+Yo712qd2Ir1P2dG84NIUpymtQE9DJrP12xmhT8oq39
uNKqKqeWbM2N9yX7QMJnzlBcpgykmGLMCAhJFI8uRZX1Nn7XbL0IumEHVC4UneNL
FehvpGTplckj6ZMSO3ZOp22jJWEB+Ni3I+gw/Wif5IiE5rMhNkuIOsgDES2q4y3N
PuliUS2LGPh+Loo674u0Cl0nyJq/v87kAJTVo80fdCntoAaZraKwq7WD3bebHNJw
zWlvsl8xtJeWypk8O0fTqXohzlJfWU+qrNpWQdloGC/y8HNBeVj+yqQB1j/52Drh
p/UFvuhOY22Fb+iQJ4rjIspCodh2gJaZBXXh6KEuDvdeLUYGk/HqSI2kGDfpGBot
JzzUdHXpjxBcY4XRgbFrtEkzV2gS2XgHvoUA71A7on/28QqpxXwMrJEZkOq2DGxH
LlgFP3yIvU2A3sZkAHM01UAorDNEFVnmEG1MqNcXUiQwR6G4NmOb15jKBAVGnVUQ
7YPzgfb6F34NASvVgctuuN7IFIONR7IPyudDAVckoTKF7QioYdqzv3otI8HeqxzZ
cpxkSkybV0GHekS02a6YDmtt1CVPwmwZbcOv9jDDG6wud7EAi5NDxq2/ZOaXAmuG
Rtqv9XyPMc0fehWkE0GKGHtxuv6ah0vpEa8LmI92ZqmDpMS+Q09awHSj/uOjlNbn
BI12CwCRtXkvvD7BLYym+9VM5Lc9433NQAKSZT5UcQLEGrdqkaMLWXBBffDWhsZn
xpbAm3pfFY3Ax/CUyLDlpFtNNdOOcs4BUG619vTGGCEahxcgsGUbrrCv+SUOEaSP
Qi/CYKL8ct1CGPN5fo6zRYXFLyRapAIfbcVMkw5Zo8RD62pYxvrNXEEBmk7e1aoK
21AibNDnqyTwJUH9Z8mzB35Jwzlt/bY7E+zReR80CEmYS4ax9hfKs1BNvLkn+mF0
AC+gAv4ykRkOpK8G5CWsI7ukzhYMi0T7zXVCHsNeWzvkC6jZVHyHYFWbi5DqM3u5
g/3qCWxReOU0mdVwzCMI5+c3jcnTGDnE7SWwM13en9LH4m1x4QOpHIlf8hkUoiTc
6bCvUiWRFVdACE33VftN707jC+JhCSH1Ifoalt9HUcs2NV3MuJGibcdEq0xgjl5k
dDvUuLpzxo2kxHkEMO71cjdas02N0oJ7zsN0P7ANgUhIdzZlyXG0/aMSJYSyEiQX
AtTtJnM5k30ZIZiB7xRTgfx5nmsJm7MvxJfrkfb0EO2QGlGGzLRBit/KJJkFF4/l
iC6rKtmIy8NgnzCdlD9h/MEDK4XShqPZg/g7jx4GmEEUjBBUTzm023GA9QxtuKuu
eJ4K0lm6SJjgW4WQlu6tsCca/xVPRNeVYenvc+EUNHZWoX98ZRAtpFEEnyp4qsUB
pzN4VSyGKsJg3WFHwIAhdNgJ6O+OQHhwkAGn7hq7mvTbg40RIy9+WXqh5gM6b2sT
xT8vBy1jnrQFKAZvfwFmh/lw/gthomrJCQeE1DzTFkJz/uPo+t+f0fXykQa+uzAo
ZxiBdV8uYMwA2mzSFCOR6qz2HysaT0zCIiPCXgLH+2RKWEza5FsSqKdsSQarECOb
Z0BjuhQb8L1CDOIJkEuxYpyav6u7BEtHgfyGWBbX8axJkMANjMjn6JeU9YI2VVxM
L1yMXRBmuVwW2W+I/rP+7y/FP3m0tCAjEnMaUJrojmvsZLPHTsv/mMApw+qadFPh
sH8zKiRFSmbxzdeinINEtYCCdXozb3Bz/vKCSoaJDLhR+35j23mFT3Y4dC2FdOut
VY2dOzOtBymvuDX9NlgDQWrlLN8JNqJEwhmQxnTCT3z+iv80iw8RdK8zGfeC1ud+
01Eak1Mfu5tXzVM41lSIhhV8tc7bW9W4B7M1UV/dUv+g7G/2SVDP7ado42aocOJv
+LCBWvir+PfRoVtIEIl4CJORhe7vqfuKiMst+UJBUq8Lxen2dStlOeO/zOI1nKFc
tbeqou/Ryk86/15EMatqSIzZBLsVNmJKCSS3c6igvI6Nmxssk3MfthGnJE4ILgUw
QWbKjBXGDvMcczjLJZabL/N/hga3Fx0pzioeGh8cdhuuJYf0OcxK1XjbKwIqrvF8
NRIdFFpVC4kAGyDSHGu4OrjPy480tQv65yuODkjFfBnc2aTZT4XAm+LGYHu7Xq0q
kivXjUaqdD1+zGiDkaYR22XPbFIddA/wAmZhUNZnVCXTLpJXpSZ5nqgwogW3byel
u3zS0lzR1VNCoOK7Sw23fnkSlf5n9JMLN99oaDaMDU7EvL+IGaWMLwvmIBD6KXdB
tMck2koWhV9+09JAB1UmqMNtl5NqmmOKrRRHCQHdpHD+5s7+o/M4IhJChnraOxcm
s92yOuL18i9W4frS7sPUUMMA//pCUKhDUYkfyA6Pp+hDT9z6fDalPTFWwl1xGo6/
PodZiXRrxQuG0vOBE/qE4G/y+lfXe5sU1iw3a1NFOSI/QSmbAsc7C3dAe5dIlWdo
1HkMv74T1KIyJIry5cOBdfLr2NcnVtNivUAh2KYCC3K7xhXEsb3VPpwHFO0HwrcI
XFTr8P4Uak8JYmtNny+rnb0ZgYyX32xkInKHuLcqS2bCMH67NQVviY/QEwOsEGEH
5aON6lwVjTZAwkS+1cPS1P/Kt5glp6n19mAIMQsEzRU842XrLGmkhZHoQxtW/Azc
CQ5RTc2YvZvs/lAlqE8dyIfCadILiOtH658GcylzNNlrz1bhJTe8QPSn7kmB6vs3
3KZpoUwPMIArY+Y5dIdhRmZtcsJyUg0+ulPoQ1fBmSbPaUUy8J7QCG8Fv3z75d15
p8fx2YdrfSKpyYqfaeSCRA85lM70Bnd7j31OmpBeaDUhNhPn0uPpEcuuO850+rm0
PaTIQd4ETuQp4SbFhQeTAYG8KAEAMb9UvGOQe638aUsjPie/wqz7BRzGzkIvAj7g
29AtS4R3GgN3L37l9SNfiqpPQSifQ9qHSICYtZdktJHau1og0okF9zQ/0dO1a3pe
3UR4UpOcpyHurWXyYVYXwf1b+z9A3u3aKRhvVPQto7/Gx0XueFYldKjvYu4DbcoK
I5i5yifgzEjJ4G0OB82q12gialpo1nnhXyctepcNFpBA/mv4dKQWBaEUCyB6iPzT
zafXM6QurgZJPImEUwYSWPrNoeFsBDZK/QrB9WXXNc5W0MGYV1Z62mtXXCTF9+K3
dy/M0iPH2TLXx7gXtbOVyI3A1TlENf5opvu8/MAdpGLWRA3uwzFt96x+VZwS72xe
M6ahLj87itS4bYNTVRQvcOkl5Iea99qaTn29SzS9ouNNWTisJQwr+lnesFcKuQbj
4Gj3nvjAaMwzJHrj2W0/SroCi7sMIyxjp7FCdWcDeA8JCGJu2HD1JM+FyIMrj6XJ
PScqq1YiDs858I0VaUYyB4SBjjmx2Zh2eOQLJHKsXj0c6eajbHZR4ipYokstwtbe
AZ8j/8jWeema3V5JbufpiXLgM7JseQHOgfWpQ0R+Nn67uR5O42gvIDqGYQ0lRtGl
FASFLaqsdvc3YQ/Yxm70cvWO47531Nzc4MHPJ38BxBUtlH/BN+fSnl7V+0onM9Xo
aStWtncDhE/3KNsIeVPdHH5FVv//Kxrkbc/9Le6c+d0b1KZjSglkmLkqRoUzL03E
Wjckn0YwRrlqO6H8+q8xFa78Zp9RSzy9D18ZyEwY97WFeymFN6iQJM/ZYfMwh3gA
GHkqviR96iOTZ1cySErDo/4ot7y9H8W0iBxrCkuSEG3uN0zZCHcV09cTu+kSIjQ4
KpBqV02HTCika1oeW6jj5tz3wHV0cy2sE/153PZJNqsNc2ZcYEe9IImPA/sdOOJj
h5/thtd/3l6jkMaY5NvASjaXtecqW2Nl28zf3KgZMp6Z+dxQ0xVJmwuc4Qd/eOYq
8x4l+GjujpAern0XcdmOUyY/pY57/L6FCZBt+6alX4wvxV75pnpSG/JcweOoV7Ae
MuPNpn8nziF0hm924zptlZ8PTJuXP4NeVE7TfdQbyGCl0mZF2972a9JEnQRjxxHa
Zx22bXwdsZddMYLVnU0XHoXCDdzlobXAA5nIKYFn/23RiZgmxvCmoCCrcGJg+wwD
rbUPa+RpNRnidTZcFwwsggLUrcIPuk8lEuJ+ZYo+Gr9hfklxi8sfr1BU5VdItioP
mr9wJ9zoMspYfZPkpYqtaShLudaUsNS8V+kHHcfd0A4K6EIBcMfsFnG3nPXoQ3Ca
QLRLoJOFKP1O5PbM3+Es6x6Hzjtbsf0JsLsjO5Jb+G9z7Vf0DZa90BWxZTL84taD
C9WnBGC9fu2uJnzt/J7yCf8Qxu8BS4DLxS20VY//A/179iBUpZ2pRX99V7MxNAmD
loJOn8dvOlBmoUa/JOapDOCZow+jFOnt7NrYjgan8tloQMcAY29v4Cqf22qGy3hu
zviB8ET4enfUFa/ZGk5RMaX4GEJlvgfDGHqBA2KpjPwdxhmXPyimoU6FPnCBcy1W
LtkQ90KwKpBVPhkGnkmo+BI19f5RqygRBWIjNBdHYGJXabCqQVa14wU2NGZ1T+uK
3ULVsbfSWMJSrGtxTm9flFa/zSyJ/qrNzMdc5QTX0KIrA143I3kMeRsWkEz73lCm
3xtX0Qd8wuAfiYhAgZ0DGbH5NzJYErQEbrwJJtz6WI9tFVm5Vn2ATbSZ5qssj74y
kF+GN1DRPw/IjH8yIXyZYfRe/8a3Hh9q3qLuOS/ry7zKGCd6ByPPq19PqQQmiQcJ
FxyjVeKnZVKb3JvUefO/6SmrkzhCAIVXuCaUhzzdGbsB+l5J4H7Eyv5zpjUeeVgh
pnRxG21n+d0ZSUfJXUYRvV0kpseV+3z2QsQQcBAgit6ugeJYiyH0KAH8ZasJouo3
QnCy7IPH6A2lIKexAEDueIhN5hFmp2AK09iOToKV9K3nBO0nzDeRPt2L6749dkx7
f+SowRyJLgh6JIGZnkQWNkXNWPc9f1zYdCvzrYZRZzqlCyqa6XHb6CQuiUFIoKI9
WqfLbSkAdT4QL28XENuwiSkGsWAZ9lrzEjsqojiFZAl74e6Wmw3DK471Uy0UJkxZ
p8bYiVr2/D9CLL2Thwp+iAhr7eUnPcYCUyXYqnb7RHNJObjEIzjxM5jps8W58DIN
orU66EvlFasxXpoBA1dDT0DvO90oqj+bdHqsn1mrojhVlESyMn1nTlUfp7ijEUvv
unlg6V3cexmh8gsBG2vFeYsWUFlPN2jw/XIRyw8iDYxjGJgJWkoCTRxfPF1lsF5i
tjm1MpZXRzrecCsl+fv8UTg6A6wP2ZJgiB0CSvdChp8B+736DauOJS4dV9m+Cuqk
LjfttRU26nyqcU0hVTjEEJ5Aqbsixf5eW5sNvq6v438QxlMeWF8yVWcQoZv4UnHK
GfrMYzTzUsgqlMXQPyqqmDidESx6+9uMtMVyTNvVKFaGx08egePpv9hlPEISPOGN
XqnIAjEgwfMrS8SfxVNgLK/fbVZvmsdTjeT3dsTrpypLe+m9PgrSRncFTb0mJ4GG
Se6BujGnv/Gevw8as9KLPNTj6oy3XcH666bwkGBD9fKc7b2qKWI/qBnZXvq4lT3t
gjePKZ4/MTqx1yOgtXkRgP4MnUe6B3kdfBFXma/NyM+uRQvJrH7fP11xthdvD6eg
Sd/WLv0W1P64I0C5iigf8K75jxkIVsk3d7Lyx3NcC/wm4FW0ZOuOhettJ2xTKdLH
mah+alvc6fiaBFYf1jWQMuKq/Gpoz7znhcNyVe8AhJQ+9nclrHWwgF/yx+ZHg2d2
ObuiZj322yCNmOUnOw0ERqK+vu33FpyTnZDVtAS1Iaou/rR7ToKygFXKNkAlTn6b
eFc5vIXWEf4KdnHQtRr5IpeYEcbpYG6ovl6/Z7ZzK+qKe4rLkGGL5iZRnfEyQX0S
Te6EjszasqckA/hpvsCorffG0wSHcKXbac4jSVZTY/FSqlVSeIvbpNUotHHowkxq
PSeW47EfEUaPSiAmF4ngfI+UJJS1Az8XXo1qBHDdpk0P8RcDzvXz8rnppWB0jo1F
6BXGGjKOkilP08p84O3ZA/zLF39D2CbI3LEQBSRRpCP0v7vxIyKRt7hpHw6Xq0Pn
XVLy+o2hjXzyjYPnuklv7+X+I5fNUZ2vSv4EtyeNnKGzGvZdnpoWING4oaz3fP+W
JbOQaVBqPVPbzgJUQdxbGPYv9qFIjIX0ZBrfE4U8X2xRrBIWt17U2qWEIVYIWGdx
PqIe8Qr+PcBxrLDf8I/jQc813lybTvjMGTIJ5b4No5glY8HXB1zMDlXisixPOAik
PzzPfE6c7QvrEFYTuYfeZ7XInX4F1pvTwJzhY9KFQLrYBrfdJD5XsDq0RHZ5oW1k
0FMY7g6PGCTWgBUir3ZuVMCNW62Huekw6vdr1oTqh4vrKPIS1DwLnR8XvMaAPXeg
o4rsGtZ5EHK517z0O45GkSNI3F27u7amSd7zJaiw+5IPAQ1Z1WKS7UoH0+Y/0k6T
Xpipf+eLf+nn7ATIkFX9Kb/hZU5zfHNgizSqPw+RFjvoYZa4t/UmvcMhitwVXzQJ
tgZbJGd/ZtuJTiQ0D+p9KXKuDF2aJSMzevXYhlnPOSmCbK7x42tDxfgtdE/adO2G
eBEf05bBU7VqgIiLJBU2dvFySeiKMLNYjOZKLH+Z31DTmxuWIbZs8TvIGPt5goEV
G54sTAW20f1CWtE33bRRYs+Pt7lahNOi0i1UVy/0MjRhhJDmpq7QvJOMa6vZztI0
w3vTMVOgCfiuFjA5yHruybxB6ElQdGYDtON5xzaFvz+6yh/mkIK9eW2nAjdxsNrU
PbMxB/3TLZehYnCEsCuhVUom/hARskfljwieo8u/T3nQYVhX9CiRZ0SbLN2+Is1G
F1B9cMgK6GmjSqv7ew9soXhabY/1GWpQzU2M3y3f1NkVRP2mNs7+IE1KGxQd3fMB
Kj1jg7FmNt4rloGeyq2kn/2Q4hoKCZYOjbSoeTaSmSmHZusZtblGFH/yXazYo9xr
y0fQaCqGXoEBnK2nfUKt3qUdNzykHExZKT0jaPhyEL6lHjmqJG2m2tNZg2S7BryS
jcOuVC6jQHUdEdyO5gjEt4e0GZ7w7IRlTQYjvqwHnHIihdqoa46AWGuTCB7GawnL
/zUACj+WtY2KA79Luu72rmWAhlWqzycL5t+nfvSysLkoDq1zDmVH2bZ4WzQCF8Sm
vBhG/LeBW4sa6iZyn8C4pep3bMWuVRu9ICJ2dD1E8M2gt3RP5wYE2YvfIJBKwqNh
54EYZFgL5MSxI0m0gxL6cgSstQfn48cbHBrudLmqf3LFy0q0GZNj4uscGT3QbWR9
ZFi0/nf1uJEVmE6KdrxEkAhewKF1SvB/Vpu5schaX9ZeiJdVa4zkZjpO6s5HElwQ
RZjQoFomxIx1mnd08ySKTel+zCW28Tv+6UGe4SIpj6hcWE+V9yBEX+hxXHzzSuJg
399E69kQzDkHaEOn/avP3ddiLU4ziw+pho4oyfGDVEoccqWWs4L2VWhNrFBDNIVB
pFoqsaCRZqtDeiNPudg/KSUhMZ/uJpoPrpTgxw6EdSJHB5W9RT1DerhFvDLzZYjO
RTz9UDHQt9koBktsMskphswjgIbMADnqNFZyATyX7dwMZTW4ibxBviOzCB06NLS4
PhcEVwmLSR1eo74ZthAqfcAmjP7HCAhmyw5neqQsvV4DQul/se4g95Qb2+Gk/rXF
WlNGZcNBgKAUV6RCPh+bG9zVKM8N1Y3QqQEjOLiOybeT6YbqN/SnlC2VARrWL5pV
b+r3AWOfQ47V7ueAHJ9Vu9iq/4YraxnmdwzKsIMR+r0tl7v5RzuRzWReAKPLGIAq
sP/gBcPCogeMWFKMLsHDo2jB/lDFSE6xCrLh+T4Ljc+wnk/gkzGenOCUc9ffGvJX
nTUv2Lr3wAxfqeUkT9bsdWnsUviiy5shzr8xz+tMBNzDcxLQIb+dJb64LgxSI9ew
51I6kviBXDUB4kWxlM1bVsr+XfiHBVVV9QUpfk1WusjGnepCPe7dOLFrQoAyJDqe
6Qs2fRL0K2vmMSYIVKG08stOw8m/NC7LKO5NfCcgYiLziYOpREy7dKRltbsWhx79
/zzRBIvKs8AqJcv1GLna7xVwDkwwpLafWAGfM6ngk1N1PIHQlWpVKyGnRsWt9pZE
kpQeohBwsD6XQCFiIW25M/SZfgtXq5KW3axTaQ1uuwma3buWaWOGVwxoS7qm8qkz
LNg69WEkQyMZFI+UtgKaqz966SHtuR3u+PB6F/s5rnrlWg+7B79JrXlcUyck4VEG
erltIa12mVzfOR7dfQW+PTxoYChEtdNd7k11LK592CKVszoDv/GURSSCN/FWaMo/
mtRxdo/9V+EXzfiVrXO/NeKQD0Pg459exz343zz1yOW02kU2jZfn2qnTWK8DbkWG
D7M84g39CnZPAFDRC9hogSV8TpeueYE5pYzgO+Z3Me2aNoKuil0ZVln1Dbrb52MZ
NEq37QkJLF/oD0JTQ4Rjr4mBtnBw8Kac7B8b8T4z/Fo9+DTGQnfyNI859/n1Br+U
5Z9c+7cIslr3tiPbUASV2F4gPg9PoGBgPTwMvsN4eT6LdnoP2BdgJq4/4aFTNzv9
J0vkvm0d97J16mEu6tqj2/0hinKAAyGGTF3tHEneXARxlaJ0P1M693ROvklXcHrX
rNKw/mMMVGyOu4ORxmo665PbzLvVan527coAVOxoH8H/R3e7GE4Z0fmpqgqAAT8i
z9STEg633zXcwJ5LvgIQkq6i/5FEGtEBf7EPPcVm9mte8zc5+M5ojJdZR3iIEqtl
V4huJmnIqCVcpvKNXGY08iVGKhbj4TYPDi4AaygkURSvCLdvr3IsjTPuvhWcB0mf
K6rCKiBhip2ZwAKkQXQufJd6WTHHVI3Se6P2/FNf+93xkSdhfIaRg+9YIeeg+0b8
I7HuXh4LGFRwZvH/pqw5D1RwgYaudTh2V8D2RW0G5w8BV0P0uACWN9knFB0OdJwl
Noo+wVv7FR2M2Zd7mM6Mxj7eA8EmZozegS9LFAKIoro74OvpwNXL4xeLPZ8jUJJ1
AkUfIKIUp75EJsDycZcJVK0tmEXZoo62Rhx6kdVl0lqFTvtxELHX7tzYierPryxr
nMYIHwyJDd97wFyqR65dsdVm4rbdrKcOnNxDEpUh5FB4HLhIfd/QlzkxWVc3mYzy
ZwOGvjj14JgxkzbzZ3ABK8D7pqjQFdexBDw53/2x5OHXNrA5H4bw989Lg9Pw1i7b
ctDBrJNUc9NpIQclFP7s/m+tZiuHMLMOipLHi6vpKMeB4z4bodaN/WKv0FcgwDVi
P2ptawZ5g/X4rXd3kUnwl47H9mpcTov61duGsmS4yu5hlhfy+qDYiGg5JWWid6ga
npUuAQl+QtOrCMOMAaB7Vld+Vc4a61hkjr4uIRZ3W42FmSG6tvPAz/Nsi8tCBNdU
Wv/hIlg3qz7YkJB7xc2P3pn7zEt+JoSnrjeoohHNNeO00lZ4HNHe+r8SpZVphGMU
+BMNC/c9QABydlzkKIXAXR9tOh4JQHPCIrLDP4LxwLhuO71SPTDKvBi+0y7gw+1S
oeVIc1ii7s0ybNAHrJcWxsegYiN64htyUhwuhOoV1jp6G2GSN5jytW5MbR7U8xK1
kEWdYSemfbbByO/D/zr1OpHQqNpgCu6nR6hkRBILb2mTxL630HDOUzgtOfqvmLpq
P8xyPEv+QbrNwE/WbiZUo1MZIiSLVz3akylzMPVOOaaf6axKgVo3Ptv9BuAThkwv
ApuCjJsFKUA8O2WPpbfYZKERaCaipSAQAFI6HIhezKStT9i698gZtaxQM0J6R1dt
SAO5PITvGFE5FJlIPSC63w8QBxvibNoknjd8ylm3NeSKOSiQ14SpI6IrVT8reRS0
+aNZcSjzERmsNHilwLEDYTulMwZVQySoSX0j77ops08bS7HmppFXeRcOFoz2c2QP
AlOJDFPR5gp8dvhld/ZSFy1QfZms/3Z9I373sS4SGK9mw/WOTzXNI60Yh2aiz8g4
C3Q3NsSWETpIsA0YrwBv7O7X4jN3i0OPXMJHffwl2QM8X/FGDT9erbOmiHc60jtP
ij9T8n3u5tx6SJZr8Ob4rNpdrUVBdYjSJtrqxNKTmhjuzIFAYU5AIztZZ8cCmKVs
mhf795DU6gOOo+AStp6LZ/ezecU1a3rcvOeMcXYBbb22Ol0+dsaMkdl5NrRQRqQv
T8q0MlKy2533LNmx5kW8Sx8jT7PiB3jS2vQhWyzHhIjiW9VdP1LeqBP8BeAhvAOC
X9Su+OPAZ6NUsofb7B0HbC3CtxfqZ7JTkrBu6F5vFFDyRhnBL7yLoSZJJAi75omz
KbNaQWs9n08ZvF3vQQCAREfCZ/6yBadG+T6yrZQU/z2Nbj5RJ3yZqahEygM86TJr
L92eGlIM4t+8ZZ9qgNlY6cNc4mZZ6+6VJkvsfG3DZ5PFmb+QhYgOWbYLjtDYirnc
HmzNNx3PcQIs+3rnCPguZicbfOT92Tneq8UEdw5ej65qa24I1PgNyTI8+n0r+z1q
ddYfYW6CbjMExyJljMoIbT1Q2XFPCHTa7cmpOd5KiK8o6NBa2kd/d4ngABn5zmDE
6TJfZ/3Sa9l4U35haINSSbqLdK3xgBz5b4WPP5U42GGm9q4nIDjJ7SZpETvWM4Le
+3n/OhV8H3BXuqZbyB5DGl5KMD9nKkgmlwNjY1pRaelzQbrhvY/GOwgddK62JL7X
/qfgMmVd1nilL+zEdC3NU9sUPke7J0kbB3UEfuTHa4KEmYQXJLp3+P/oKlfwnabN
AvYx9x/wR+ZjAY/zgunE1E/UuLmRcPOb1czxqhh4BGY2jom8BsjjWvsbbAMXHeBl
bdn/loImWQkR/UKMgMTuc95wbeijkdKeKxck3BqbCYNxze3JAN1get53CnzuuQOG
gQSZf04r7BTDdvldlyTsrbNdSu7RTvi7YHhod15zHA+EtqutR41fPBYB4kzwk9F7
FWYZldi4JUNuOy7VZ2cTQTxLy9RFiIYI0qUJ+XAtLhlIWHqpRO5zXK+XbJHUR2jY
SJ0PFg6RFX1VW2x4TCOxDz3RMogvd6Fmpzo0kenwsgW7IjA3+Wh1Y6A2vLabv431
4YI0ptsVAYspaanD+/4f3hQJOkLO4gVSwdSohfHad2w81Ic71HX1JiyfqebK2UMA
LhH1eKy9yrdCGVg0DpvNYRy0o131pOibj64NKzlP+YlxoIEJ7aa2E573ta6dTI3t
6CxK+FPIZNcNNHgXJiPukk1YfTUeECk9qHsCW4bQfJRt4se5xP3YFI8RGZAhdLoL
EJQAMmpxBMAwLXzQsIeNdN+otZuL5NcmZGE8idcI8J+ThGT2lUisdV1zQof9S8vZ
5XZWS1/hnjyZ5ZB4JamqcNxN4nI6GvFQj/o3LBV4WKUmDmjOqs5A35pGQQn1UYQr
nN+xxMT3uyAbf0p6vJOpP9AC1OHjl8+B1kHX2KTNEHvdFad19z1druscWgULc2FO
OJqGo+XhZ88ek3lel7yTZEnvpS0VuqAvNx+O8gSN5PrMSuHJEiAMKygFr43d3zHO
rpJjHW0+fWtGtNLYZekhMQwYOAe3EmK0WSChobauhd21I6RjLHTzNyBO1fZEbyP1
w/EGAbXKYAm7S2qxYtCor6XXbJIC47nrWRPBmfL+FjkN1jtCIwgbtFmt0efD83j5
hgvy1IPIlNnYYkmuoTI7N9rO/0aYazON77///1YEZfk41cKqy4qjHJleZyyjZpWz
0mA3aGY7W8rpLPzkkgfaOcw2xHOCwXffWYXCLNE3VAy06p79PZZ2e/qWgYcoe1E2
IR8JSdi/R9QUxAZnAka4JtplNd40fmbw9BHBRdZ6esGdJXIFC0w87U4lbh7gPlY6
AVrsu8QEPqYeuGPaPeoByKAHMs5Dda3M/pCUchdqwGRIMafbeOTz4eG5CTQX7Qg/
cYzu0h6sju7lOpdUBdn9CWCR84zl4rS0WEhQ+shdHEWokcx6nWaVzYYULKwuLH9u
GBdk5crt6lsKhFMqUtSABdyQMajGbfmh+SMzB5f7NPQ=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
T+1Qgam+gIPRN078LCtNONXHjpjKQ76mF4ELSwJZwIUIbiXSwgcnvUpgmUhPewzq
OJjLSkScottG/7UNE65v7OXD9h9VhYFwDPFlATIOv+s9DONr76+0q2tZgvpszhdI
TXQBZRV3xmNeNEDf/tWqe/dZM1gI88n6JMTpabBustxyn9oO0CTHV64uHOl6IkJd
Prfx2dUaeH10+4SmqwwKmazhObJEntKbkbV9xlI1QA4TpTAmtPoeSIkABKYP41/3
NkJgZrk0B0PRmKEcL/4bYYliw3/cZmhIP4SX3H0D1HyUtogZCSRzXPy4KpKZNxS3
7hciY7WMOYayziXL578aEw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
JXzBxXIKNsM90qq/Gr9CCipwudJjCK/mGU+J883dwm8kVQtfFK7nUgiYX2WJqtG8
OgpL8sWCj02jCvYjVtCqVJLfg2dLpatsqU3PlchB22Z3A2p5z2JqKZLyeALOrFgx
kya8bWydekepZSvUlfQlVBXrVSGTbZaue4OQexizbYAf/FKJqNmm3nFnm1MfH3jK
sQR5i7/yCkupn4deH+xm8jIj+2zrGRZbdx7IRBODBg7O5b72bi8EmJw35agR2QT/
VFhctw54mGMxRJ/1Sp6JnBS9hA4bdoMJxzz5WuF+Z7DHNPYp0UIjvugOHMM6y0eO
ZXOuWo4yX1m2LgRJ0RdQjxBrGo2UYuHyXxfX8WvCxiggakg6306SDPpqWwW27MdB
9Inckw7VSvYegOaexbe1O7/YlNblUcA7PJbDTMwtVqJuEilHLO9R6E+/BKWBqzlO
71YPZhg1EF8NwPWkjsXnjBfo06gwdfEgtAUE1GHLsJysW3/ow6Da9AFW+rM0ehyL
9eacw/y4NLBbCGC+hPwVWWpdpJM0914HWYbeMEFn28K9aAXgje2sBN11Zf1rHSqT
9nA99mP23DAbhj8WJdkzCT9V0CWNLXBq1SoVcWz2YCsfXKNuuHiWoMhqcvjz7KlI
bg14fe4RC+DYdpu/gPUjlwVDCqmGVqYFI5YJbCjS7BDUlUSkUMTEZJAV6/Hio47h
oJ0L8rxaJhf5anTAoPIXtbj5YZAfwQaO9rm5bWwdGeaTI5sMc0qDg3PDpVJhDpIu
VkNq1/oznTIjIcbTZycUaEV8BpnH8guB88dIqC2I4eL5Id+cACKLz0LnyMfysxLH
RXP43LjO+0wYXpzC3jSjOUpI/2TKtdbz90kMYGeGUXjLpe9Gm8cEoUx75EpIEj4N
IYwqyXVNeGlBDEsCj9093oDEv5ICtC9usHgR5+xorigt87DSrGk4C6erOhlUgUSM
x/3FZuwomAmDA5MTElEwe6icP4alN+f9GwVh1QYDlwXY8nI9nbyx1vXDY/7pn5e3
QW7NJdR9PsWI6B/j4T5TbyV9dqmnUOY2FoTnrmuNZvrUKcKMuuL8DlCA25Bc5J6G
YRQLTt0RFLGaNVq649z6ImZkCxtw2A3cIvUHqmM7B8iNUfwxQhJlJZdfzo5e0BRk
GzX+gZEXjzWSUzzklCNwGO2XxZlXnEI7BGCFW7YHx3BfgnHxV/U2uudqXQLnVb7F
eX2shkvjxJ9N/uhBVMYXUiZrvZCVoEkSak2zFhV9VK0OPEJceKLBVUADNtQ6PQtp
m8+Qw+KZNgdf1Ku7nMU+CAjgMoyZrEYjHlfbsPk+snEQSD3eVpqgDrzOjCYNQg46
ZwSytbJ/GrLUgBV+4bxa12LClbUhuDjwe3BLrUN1QoFkL9g2ckh2M1g64Lo8sNjF
r8AO0DtER51TEG21I1fEiEB1axgymuLdImUIiu1aZQx5metw5PFue2dUWI2Dub9V
Pr8WkDdyE5WQSW0JPJBQm56dBv2/Ws5CaoAqVg1yO4gtceZFhtnwmtK/AQqc9h5z
PHnk/twk/GFs+lhDukgxXflvkKS3lUWySeHS6O2rdVXq2kIZLf8ARRhubAvc8vcZ
U3Ecb/9LJyONBcyqW4mnBO9ixgmQ00pCMSZwrdHhhp9UV99eDl+rAFqgHWO+7bTz
+IkTld49FWeUfogafMzRPPfoUTcmpsi/S8h2rx8fjucaFs/fg8WcZ4XZKl9EZeEp
y2ne+B0zK/RwAsruyGzfSItd8UoRlYtbJXnEaAhBmhDpJxGdn/e1QEI9QXa7hT+s
ael07lvsRsyir2wHj6/REvO2Jmv8xWiwInwJn0Fu/UKqiy+bO5058d1Jfm2rzVL8
xTkt2mpWCa7T2x5LgOsOdM7q1rmjoHXZZ1HTQ2IlfAcB1cpD1bws/+6d5QAD2BLV
45Etve/Simb3cqYL5qnbYNFSdyhWHqahU1j+VXan1Mt1uN9HTHIu+fhmoW5eJL6j
jbPnWfbV0QDGX0JhFQNHjYcBIF1COgZQcWP70b1hPEUpck/ClUCwRHaeyVhj0C3f
QJsI8aClWw2MDwVYlJxCdXVW9tSkpSZ/c1E+wS9/UjKkfeonIeueEp4sDfgQtYOU
mo9/IZeNDjEjeYtzlULgdflDdubO6YoE0qHM5nXPqmqV4k6ZEr2keJfoy9O1P6v7
bFw5SX2GvLjbrvNcyK+joj5x6zkNRK10CNBiE33E0Ose20l+wHSTX0jfIj2hvTA/
Vg02hYcU3qQWduDh5TI7/UWoipkj96GAqPyYayw0EhGxOFtIuZ5eK5wTFv67XiYu
lFcqLWEXxXbpnp5Q8LqUd/08aMulBsksi8mHuDv6bPxXaBxiQp0VRugjpmyjhpUk
elBV4ZGLhEfbQMfp88z7QFx8gRxFBaAnzOX02yusAArc+ddpcdxBVGetRPhUridY
3Jfgz1mc6mtvapHeOkgYX/rEagLGmTL5aWV64cAuN794fWS2weJaBKnLtVsiXwdK
FpE+3kc80G/cSUNfhJacUwCGET8oajBTIpzCbShOlBb4D9NHRT/DIY1y1Xh1MvVZ
gHS0QQcbvGhRhFTtMHLnDDkOQ/8mx3fV8ZfFODi9+KshtVGOgt3MkL3onljLbD+g
+gWIDrGll/SR/br2zZk0mihRWMjgiY/XAJJlBIbHUt+QEY36dqyyDrxu4bGo7uQp
0s2uvG+hBmH84XEaOUjjH+IXAcQh0GYlkYgvSV00qiOHOzm9mlOgzTsAJNmxwjpW
u7ih2/pfm3/cvSVGVO6G4uckn3YY8fNfAhG94TBaGMN6ZLdnEF3todWPJaYHQzvS
NZMr+/4cYSnHW33gVQZB0Ohb74fws4ZuLcbI3cKkMnZMmJTsUepQpNyMJszrfFPF
Uvo+8QgGysF4HKTpNvKEEzV0Tn7hl2FW0n9GSH2y5kArCD/78Tyqw+v+uu+wLMPQ
m1Bovkybz2bviSSnBCr5h/+mP9nee2ED5HKuPiZ5birK9P62zWVQbjnVqkBkaux1
iFx3IbStLbha2dH60bc9J7AvmLTxfllbhzF65J/QlPYtrzYQZueyQPr4YKIWKTc7
L15k9CtWGm08IPVKPt/DglyQDEH5TsacmpylPjm1KlmcrVG5wd1q+WwjXHfYZ1wm
Mj4DyUBZpUEMuQACpGTJHS34vgamJMxqKY1A3Z7DhGTQkUAp//vD5g3QQxyPVRy8
Bfsc7IjDr4KvUzR/+qB41nyozPbOWrXLrNQw2NzI9ld+oCC838Qvdq/Dpv1MFf9L
KOOauDSTiUkeZ81s5Zh/NKc0JrbqUemaBdii3Eze3j+mxEVQeCYWttGXKN3rStge
miIGgrEfH+34kT0E4jOmgoRsnq+25NvCb83zk1Xx6lg2pRMFVd/8yD7Vm5WsEkBO
+yiC+pXwD5CZSOvgrh8nFxnoaLVt9S5P8nSRELqLa0e1vmuYtbWrQK9xjIo4DEq2
oLxTAX0/UAoG2hbEE4D4AwPR2mjDV0x9+evd622xYHSLAfPF6x7CIvd2b/YanCPt
j23pd4gHlsyBkevMsccPNfWMsaG4qcWqM5n9ZEq2Vj6ghVTP6POuWGLJsTM5UMgy
BYMlBhMFO2Sz96EIKhuVeW8MZc0MgHs+Hg/2WOSzqw88B5PRoHQUPnQhH4XpxXOZ
A0jtdRbZKXFOM5lhVV4oIJWkXeKcfcl8uYZiiqWY4R8zir8pPAPvUg3lyP5g8EKs
QnLtwofPW6uuAPqytKuMM8M693YwpNpxGIxF/qU/SODzX0joyxATYlx9UhU8R0+V
cKB5Y5Y2QoVzK3DmB2vp7/mgBQmnjYdser0asnkmZO5q3NcSuRiMhWw+S4/6UrAQ
h7FncH9WsfTCHGrb6EE9w/m9cy3WMet3ua9htpzqwCx6YOfpFXStfNdwIRmLRLmn
HO4BwMayCwAXk6veKJyihIx6mAmxUhZCTNi5rydPL1flURpJgd9GaNP/G4zruPMk
ZO3sKM1ENzOLjcoRoSwttA6i9vOrmEt6nIWlcK6eSaPdiHHqp2YIOxRXXqRu9thl
yxzyzF8yA09O/X07sHhwh/rTYyWKxPiKwbEHgHdMKpBEDgjvbnMwLbxgv6KN2OfT
oZf2K2eqN7OsiAp8fBoAKp4p++GzQbUIMZC0OuZVHQS2+ySjcWN7k4ut2EteJyhK
IcUbaVNPzDoTBMfYCqf3w9v9y5CiT4IMEDnEkwPkVsuAHlPFZZa0bsOJdKI/JrvL
5gcVgCRFHxeUzLrG89WY/7NQKTON67p8mklaytKllHWE5mqxsowqQvqLLC7L2qOH
L+efN2282i9EjixBG0h7uVSGcxdWM5btUaHDrcfdhMka7xrCxb/KStq8ZO4pTb2p
1WhXF8u3gQE57OQZOlTvG9/ylCZ/zyaei8wArUpMJzuKn99iFoJy939hwLq43GTb
kOOqERp8nG5rJLS3cOkJjOozYzNqj9TmH+jBZWz/sJvArlmGqKZWYSpl8a8X2SfF
kuLzBzEtUbD16mtfUhx+gOk8uf6wD5gLEruukedxqeYgrizF9u32nvvNvxw3y23U
EGgTr98UkXqweiZfL5uKAnO5dAGDRaPkhgrdJbqTX5xaL0j5DHkFaprvEmzMOLLe
t49b8qrDAx3QLBfNf1UOTizU7yXUlJi4FRAcjtbgu/4NXvMqQQJqkfUfDG8S6L1k
vuWW8aHKzQ1Ju0yW8U/rbnQw3YZEl7fk5xlMqK6z/lbXKXHK9Jv6xnSvHPochkfY
2hadxT+BgNG3KoOX5U8ilfhVdQ38vfHEwS7iP9rMOvfNd9lQONtw8S2s1OfeYZrO
Cwa9aRoEnXf16gaLaTgvLcxjoz2gIQuqBn5+xXR6vj9eK/AXRJhDQ7/1TVH6Dy0r
jCJOOc1RCHnrqdSEM/kwmjQDvydHPuIkBTIDhAa6pxdYtCTsiCtm8jnWXOxr+BDE
6Lbono8noJkk0I2mtO4CDy2wMITeEsFWnUf6TMppw9aRROhwhh9hlUBsCW+B6yIo
DQALAUIUScg02Jj/X62cD6UkMiq8VTIH5VVN/+EaQD5K4P5AY8uhgRMX/VMuo+6K
yB5lWNcdWAa1GKJTGuuoDy4U8orhT6aa0uSjvGUmyKG1AYYy76kK+oU7rhVpgybO
dWLiekJH8Nb1hI5VbTCkn/4TZM8xhyYKeZAEHzyg3oj7NAxQ+yMMplaWAv5czgac
0mtsbsk/7xqB1KOkalITOYNktQsezyLuI03kucMr55ntJr9DLfTXDS9hDLg6btMJ
nwdtKil74gwkpL6htGpg07xNbgw6WMaBlYAUBcoYlpgOV92PwxEe389i0yZsrZs8
3JNuStdhJmAFPkZczXYGnbSKFd+7nfde/3Ffa2rTRN2h3RHFM2jkzMFdizkZWeLV
Lsa4orlDSStA4iGDdQVU3HpbGGqnNwP2t6FASw00k6UvXprDo5CedeySN+X0Mryn
IUmvI+oRgmKWA9OaCyx0bL+x/T1JaRF10oOv5mhluX0mTK9GMR0+t6WRkYFB41mc
tuF2Yb1abUjo9zCvUYjKUQVvNOkCRNHQRgGrqQaRSsbfSdrAtvDuBH1hljI/0yCm
GqI0W9hNRnstCjXKnzwey/m6PkjVp8vVbKmQ3Fw9WIW/RXc6OinqQoC8XgzA20/o
IFcW2R83g8Cw9t1XbEsc6Wz3f0p0w590Gwh34Xwpx/8HuNXDyRXxwPu4yfLcqUxG
jBQGTizTselnz7IKvSdjYMiSH6r/yhSRt/kcHx07bpzXPbG4OYrxaqRFwwTNyIia
aVs2elU5H+z5UZrcIRpI/PhMv1eFobE8O9e5svfa5nR+4Xgu5T9kR3S2aoah3zXE
TJa141LSySkMB62WsUac/Y3pZkBwOcC1gqzsQEAxBxN8N8WXltBPFoEV4uHrmvV3
DCg6hcfkYErpicOJEeA74ikcfLhX4xfgWC6+zp4Jpg7iIsMTSlOmvFF3mgMr6Je0
QY6d5CJi9sDWH5m/cYhvHYuIFEQZP+dSqcfCWFGg4wBb52nAn2zYP4voOchbjCWl
lUuVtn8Q56qVxBOSKcyiHxA7U3r+6GNzO9OH6XyJFju1gXqYiKhRbgWQBdcMEMZg
9/hcedznWY/lndCVA34Y3gFn6yqDdA6tZGOq4eKAvEM5+CSNhA2aWXfOKX2hXgWA
t7muXJP9unq4MFdm9AkmYjZsIwx0iIDBKALkfpeWtzp+KKG3/xpnAnQOF4QQVggf
gOBxp6mg1bfymO9jPv7RZpWBYxUhthXMX8B9TcOm6G+T0nxIID22RhGEoG5isiyk
X2pNNERyPvKelXchypv/RfUff+/Jnhsd8hn6y4dtGTJZ/gZ65onFUf5dMAw0b/ea
BhlXBl31WqhZMiCxlR0XaVpfRkNF/h55h2yBhGbm2iaxrinWC9FsJ8+P3RIk62LO
pvIgpxC3v1Ro12Q51K4c7ka5k0C681ylaw7Ng2M3Sd73DPsbbyXyOijf8iOw97fO
wFNKf2jJ+10KcmaTRgFbqJ+deOvX9rZZcUBDtQccv8M0Fz3XL8RPT4K9mYOZUCPZ
Vtha4vBv53J0hxBQOkFRyYSxAmvgxH5q+P4z9U3R4m4/8suYZ+41EcACJxaVWZ8E
U6fHwrldp0cjAnzExSGs09KmRYRWBKGKm1lObMxVR/S72uMBRzhqOGB290n82m6Q
sVKDYYQ4nQZgWFBi3vwcELHbZEt331hJJNLraU6IZZVXcX/9QLPnjJYyWwiPhbZx
rnTiO14LRqT+8YGeRdaQ0xJ/ZQ0JymsKIPyh/UtNu4MNNM1Xf2vAO46RCfS3L7R9
508sYvxzOIcswKqEtWRSziuko36tAjw/y0aIh7/YteIBt3eUBdN0FbrSgrfxJlNy
Me7Vg1yxG8O03qhDRLxMYU3WYUhbF5DIb8KJrL65f6Oe1bIdpsMkIibLSm2JUhcz
37fK328KCDTv10pAU26PKvspZxCRawaiXbncoVuaCS0UDhEm5liTFEfe2HL+O5Cr
4ziPr/0kuJQk8l7Wi5LL2r21QwIOpu68AFuKE8t5atCL4RunsVKofHTnnRKG63cd
sue8AEuufI877/JUA6pTKMZr6XiaAmG8+5BgpYqtlF5aKfyUatg6IR1RO4OIN1rz
Ixk9okvPICCxsmpOMTKgI8+5dBa8syLFiamwFiRO5kuSBbD3EEBWoPVHXpQM0itf
Pf/lIUD+/8Z5OwI1l2X0ICUGzX83NtTJtaTJIv0Y/CUjkY3KcVzdKZJlNG7IL5h+
VFvp26FXlXPqidB5Akqd/jWzHW2jrsnc7azh3ybi8sdnUpzVPc47VWLpBh0FI6CV
BWg6aGHh34NsQiuiUtwUmTFEWjPw8DH6RXaDPRVBdrQhre5mMrZNt/Y6KoaDARvr
ESuw5MJwJVPLvDYmRM//3AgzEUXnDMj7tWYq3G75oC1ejjGYEf0kuYolZcLxzSld
SJyhp1SaLX9I1pVd+xwxFjAuQd1zKblLsUacJgMLRPYVnas8wKl37whiN+SYA4rE
7gTEsf/KqGpQPo3v6O+Xq4wS7fPyBz/F4Kn1hlRmBk5pc+18jKLR4h8uBIza9u00
6kwgR1cNz9d9cK4Js2dattNGFd5nX3ubtOIbWH1igJY6jgq6mF6dgpUtaJ5Q8WSP
a8/rtYjuB+kK2VfjrkFRQKYtpmoRyV5SaBCb+03tro3so1F4Fg2zs85fFfDXsgVv
4uuXBE7uxiJcGbqMuJzz/xlG/1S/JQ6u7URQO3tzvYRG3q+im0bJ2qFoYK3GsLio
Yj7ix8W3ZYbsPjPtFLaSREhW0pUExgtwSL0jg6SSKXY/ITFgOziOSENF8B5TRJo5
jcOBdjAXeDHRyDECvQb76C4kUKdymrED9Ib7IW0jFbJTyQzyas3xYeavzKg8C7d5
0+Ju9FcLKA2iJ1BguYYhEwXJy/xTRHQg2RJsc33VGZTo7AbCpe62zfnBEVfIsmD2
vIcbOyT4xnFt0232cLuDrvQ0+HOy7prCb2HSqAtWb2hLHedERFSGhNjxZ6FHwTKp
i1CEi4pdJV+ll5wOVVQ8ep1eZRcI1zdguTXG/hRJLnzOQGG1cFmpPs8s5tqdNtyE
Vyb1EFQ6+uGBhhjIL0kE54C5gFrHKwysUrgDzzrUSBxJaIJmsufZP/XlaqJnDwwz
UQnWLfgNrrEhDXVd7oAt0HdOuKBpAkqLmokVbzeL0bqA/mR9GEpxwq4NykLE2xGX
uT5sDMrz7Ek2Z6FPAiqNYACUkJU7wu5UVSpTJq8Hq2uXmGUVVOnpuvkoQcKYwuQj
zoiI57QddaVSRLvKD0fwJNqm/dPWkF4QwtSrWUhimYy2sLxwx2HiYaziXYJtDLmM
gclXEnCmchubjHL2eNE1dLtW9cRPnexd+K2H/dxlTOyvaZxKWglcyMDNINyh9xkh
0E7S7pdcwaMTuytaKm2L/wEYimSmkBvQbmltp9YpuscTDKiFz4STjx/EBVAJUy2P
VjxzxqNMcOWxaU3hAKjf89/kGgR19pbE9r2IVzotX2jqoX0AuzWEFxyGXEXcPHR+
Mz/mw9NF6my0s75lLJvGKxCCuSTTGVxeQgS6ZHP8ssAHrb1qq6RYTrL+QYUhfHw5
j2oEYbp6VqPYQl2a+GKfcQR9mTtPZINw6Ps8s6rdr2aFRMEImD9P0rn5lppXwUIB
ILOtM+POmQkSjctb+Ow/T72G9h6ZTulSz+JX6LQw1/uHQjuDK59sxr6+8cmdSJ5f
EUAdjXOX4lrLt11jvHOph2vY/szSnazVPijKfxI3O/kFMvLr2sCPtRJPA8TrIPEU
3b+eTiCT1U65QanDj2Ko32CuE6RVprnNA36uFx/Pqa5wv/SuNG3IJbcKhmzpbEzS
prsDjlqkmq/vjd5LJScYok84jVctHV21f3WZ3kF89YHfI6vI0QgEr8MoNyh1fNqI
xAappAIeRekiUmJyyhjx7WvMPctZhmikUzQreLWJIebiOumBUEurFzG6gTOuJNeu
x6G42QcG44R/eG6sDX2LniC2waOjlYvz62dYVUk28y2Z089kXVbgtwATIuLqscjU
9UbeAWlA1D1Wjd69MtIe3MCz0q4lliGcoa0ElOZXe7FJxUvHfT6AW3dOwTF4urLB
sVIXKbM4/nysikHVPK5KhakhWXe90e27dNe7EUYfqd4ukf/m+0lluo+PtUNFHndy
K62/l45J75jMINLyGh5PoslfSN6SJfYOfjSEnOxlYl3W8t3hkgL7Clh3Wpef4Dqe
UU+aF/7BoF7pY3duLyJEfgpWDljUCmZWfJPPQ0bHPMTtzzLCrTh2p0aHOOtLfrii
VvWjh59EMOZ5oHybZZKx7EQn9YwKfINv4pAHWVN1dinPM2yyz1wyWzdXlfksA0WH
O/Rj7KK/wYkd0+Aoqk1dlOAFs35bVFrVrPdgZJ9V7eZ9N27uPbIRGPUq8BWjR8iv
Se8EGmb9WrNLFpRI05dTs5nFG9FQRx3seHxeOLOaW6gDvbDkUalEjh7lNMGPElZG
R+8YdBPWX+egis4GrwhHgJS9VB4wT2byc0xf/E/hBCrxvnPXX5q6Ta+9Pm1LT72F
FBcIPSvUGpPPVz9r3tBTL8rHG1y54Od8yr5E8X5d9Sk4IaMnBGy9A4DxW/BhQUGR
JkKQTCeQ5qDatP9exnON6M+e2qhaqShyMcmjlblewfh1KeK8SsRl1Fwds12XoqZW
mmw/x5E0Bw6FWUuNN9SHWPppv2xKCKT6NH4HTRSxxS0vHmCBm8aCogSvBFYhOeUg
GbURb6x3IzvlHhdpn2M848kGDdQfWqza/1dybnBzhlsk/Lej66D2H/OdIOU4b2pd
YZscVs+DpZsHaMTpi2QlrOsw2qytEJczx8Yi/ruxSRODjI5uywL/xTP14MiXghuK
zbeGF2D/HzIgRBbu18smT0KDrNkbiF5MpCWmQg74FVgS4mVe6Yot7pi5WDP7KRDk
qS1sOU4XnAEKWYdugu3VL+eFft7JvzrybGLqNwrekkqBRRU+FvX4lQwjh06+niH8
M6ehyDVzeiG8IBBcGO0W7pOD46gNI6xvRfpR1ZY2n6Gui4qWnyjgdlpW/LAjC/cQ
q5OHgm2s8ArHdjD58cgocUp9IoElcZDgzBXMUJBqzfbW0av4JDouswPDjOitzQKz
ZW9GByuuYyEKzPMk3KvSVO7E4hB6/d2uWjuEbNclD985yXCNfR8VNJVG77fZskQv
kv+Fw59cPFT1EmZIBWBTFpqtv8wljXbg1G1dA45rTARCwyIwRmHv8LetxuQ+PX0a
CrUXhMnd+Uwn1DhfcUryrf5KJ5Y3Y4PppFPtKPgurvy5lkap1o8jdYeZsV6IDR8U
MU5JW4H9pQ8qVsTMxzMqNn//jiPAT4YPiohDkwx4ElZy0S2cMZMF9A59AkscfyzZ
P72QfB/qC3k15LzLARnrEiEx42JnQWi1CKDYJsf4Egq07PMG7HEVBvWBBUuZbkpM
9hKER237WWtcJ1x5hFWMoxkJQHRcYP37KpwwBkyRax86f7cW4OLh+nsx166Rh356
h7ARO46eXjJj+fIMQRCGQY403Wa6x1lvlRtOKMcu1XBByprVn+n3NeHPAcddZc42
0HN0iT7denBcwA5mrucQ+leYIkDn2UZSyCwKjJ2wVGzDGIQ/vzXXvEK1fyvf5ncl
mKAp7zC7GvNy4vdIVrCVmg0E0oTXf2aNcDwehZ7vrgM+2Wg+zEM1ap1vRAYLksyO
JAgylVJjYqJhrRPc9QyaHLC8JoebP4pUP3gS5UpcucMuO2hXyUquFXmelVXqHPo0
0S0sSeJIMfMNjmxCfGSHXqjHuMNE2VvjpHCXkFYby0yHDNBgRzmynv1xjMbkWUzG
rY1ITRkLQ3mLL6tLu+dgYR2TrIN8WtQAv+R9CTow/9Ig8Mxni+M/DWoPsQiKGWEU
jzCjqhOD6pfkzlEEn1uOqYSGkApLxSmd/Rl5cYV1Nq3QWB/xcJVzCiRsKsCqeXb4
+Ac4la7tMgJZWK0WRwaEcbBIyKVJTO06Ivh1+OfHM6KY7X8rRciPrIU76LP29dTM
Whmew5mNHe2Fuh7FJdeZwyC7jMtd+MRoWmzskpStzEVjbrhi0wvYS1mHuGyWB8uG
YnbGGQnoK1hcv1Xhb3fOhdYQSVEzxV/+UPCCEXjNDBiB6AKebMRv7k2s3Iuvob0f
1b4pxrECIzIocremPkHcyQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ccWX6ATTtVLANB4G3vJibBraY7RrOHBxA+jEbSPLUWIRTmvoEB/nLYSeL6+8lCoC
k5gKUFalqs25lzlNY+1DQJnun4/XH6wi+RMX+B4E2dFjaRmc4HJD0bESk+CnN2E7
ved/IBooBSDxGvVxYknE8hUTUR3Rl6L+cZBd4IBGrpluLUTcHTATU0ZdN7TstU8n
/e+NWMBsUHzv7tSSiNIfSDz+hZCpPV/xTnPEfyoCRqDru1+520bw39Q1lCrnSiTp
spWO+IAtd4McfAIoPEDCyi/DPNvXaPcFkXGtJ1cfuW7dhqa5ksBPyHNTXNYY/9kE
inixnVigFUtK0ql1tVSPig==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11840 )
`pragma protect data_block
n9duB6tYmw7rB/ibV+NQrLOaUlxru7+iFjEJTc6OviXWI1vQMtv5uM4ReNnE0XDY
vdGp+dgbanTGxRjsIw3Z3vgs88Bb3NX/0cgSQOyJ4zGupmRdyv331kfOuHsrkPXM
ZGR2X9ECs4xLP9h4khvBG0warpcD7dgVswbL1xd4OS/Kkdl17iDRCy/uiuMDOvm8
06kbrSHevaP4PgCOTIzFHVizaDZeg+Zdruzo/acyTXA9Rp1t80VwufrLp307eNCK
uzrESnIRvEySVNnVXfu/Pa08BzOR3LIt2bdpes4rsckC5kOkOM7F/ZV2/ffYvify
GI30Tb0rzMrQC47fphwSS+7FEcuKb7UbSyXM3ckhM7AP7dwH77Wkqh/eRfOnSada
Vrm174s8FsY5UmYXKdvJdlC2/83e6sDUB5xcJLGAwMzrh4cjNdaUCUfeWyZd4Tvq
KZY4y5Ma5wFtd8HXz6iqEoHjWgVaU27aciRhHnqjxWOIkr+uUlnBCAEbS2Kk8xo+
Gc2JbWt28k7kFxgs6ho+Osr4ZMkpfwm3gWEPn2PFwierHnLF3NypIZgF9rhPJcoq
snJJU2qYMmRAhD6RHkqv4X+M8iDtTMs/dxrb1dJnpuXq2QZfkAZ3WjgRHT7cJqSX
dNfujBPY/+kg7Gpa5bg6yX3UP6iIozXR3IM46LFntf0TSYtAT4lqDRsbX3UUz6Ma
bkz5RA5UF1DwvBTfIIO7UpqS4Le90BIK1PJRDrTNyCmWrwZ83lpQ6EROFMy3Gxex
wMh0scFTbmCMI8Uk3rNzZJVpgyXUBKxwiY80jCNB9C4aOrMgs8ut0m1RgyLdKo4h
4ipWhoTn8FU2rGMj/f2l0M6oOkayXUS7s/FVPP9uZ+ma2pQSbZqwHVkGfHCR2Eim
7pRG15HonwOp8Cw4UnrELQ6wLWjQVaJsfuANfCzHJxNG8UN4E7GRBQkc6NgTJOWb
WtFpm3e0iNis0UDx9nu0X/1O5twvyi87OYMv4qLOqSMG9eLiavKpiQaHoJgGqmhf
4aQmzKTEZRwo+mSVE/PyYOXZRaIAie4Xs8woS5cyAAIad+b2JcSnlPtY3CJ20eyB
1AJJRpqRITvDP1oy0wELiKX3vzlczG1AdBMR/gC3rc96KKvlGeKDhpUmOgjxOvHy
DVPQTBjV63hoJamqU5Z8ce+Btumb+7DGulPYScm9AgDSe1/BRqc+fa9+dDTZ8MMy
FwsfYG+hO4gEUOVTo6oo4EnP40A2rR4ZH6YvduQ52VeZxePE2NyGZutJ/2ggi+ug
pKOfE9ZGeLVLlYXwukVa4hBz0do5QmKomIiqRUNot1+E9cngOgEbpQ5wn/mQxruL
tDX/IijXuvZuCfC3PnedoBvXAm/C49Q8GMzNyxd/TU2xaKD1HWN/3h+eXJMkXo7p
ZhnbRQaEFz01vyeRx9XGTEfNFJJVwlNxTPuB1NfMVM8y0c+hBMtjwyPsMEuSuekb
kb41+CmysRaSpUqg3qmOHD9noxNwQU5Ok1v5RPEGmgakd7k8n+C0iJ9NWTrI6uZi
zYfZckmFewXNxzWb+c1GvSVyeeoF5GaIYz+0IBc6nZwEJVB1cWbI+TPV2u4SnPx/
+4XDEw7kiv4IK75gORcbs9WG/wiNLgmsDJ3DwWqvrni+SDwt6E68JjjoyGPGjkPD
Y+pNGAYmAuO/lnCLIVJ3Pxd/jTdO8Zfp1tI8aHPVCiDKEsDMrDfERnMrfzmUUft7
sUreSjsHi/AnVEyrhhInLx5afZC1GX6eosdZJWkHWMEZ6dE6aduetinTrAOGDMON
OeikZSU/i5cxEL74zVHlWpuGRtbbPOXDdUz5q8UKHwXY5uo/z9uPEBbIBQlDUOTD
XphIdyEO1NcjGII8a+8ta3uujcvJ5RDDP5jOH2Q1PjDY44j2eTImCpapQDUEUIqw
mMVG5OD03RgtnMT6GGjae1U/QSSHVBr8Pndg+KVqPpFVjhCwiR+TbiSwiX6bVbwD
3M9+nQzGVmyfX8FtrUbXuatE3U1t1mdWG9bxDZUPCEj7Z/0oMIYVGWhTSsC8Edvn
BqTjQwvmi0qVTIbtRmnp/f2/T4IPszy4/nokKUD8MupniRpgc96xa0XV2OsYiSiU
mnYcvh5u++p61A+oMRLkgEfhyG7Blu8MoqMMDaDZlZtYSQAtwoZcmP9YVVOYw1aT
yyLy6mbJYH1ibl3ttkPDA5i8vcrl87KfJ/GuYf0zefMQ9Te0Re4tLVkCu+4ekiM0
jxxfposlehkgrQMM609GtssGPoqsTkLMSkZuLfpYi6Rs/dMQJt6yXnBbE8wfyPHq
t/tQuh+7YM7gnxHdFoU3++dCAkOAtTCQQ3XCEA9x4tuXPW35uG7pe9cRkjSSbJz4
DTETWdkdNdWLVN9Q4OV5ujVgfoDTDVMolOFlDxd6pb42BddwTxmp856swZ/yNbDN
zjSAh1mJNWJ5LlSrCBhcYe0QZgbxi/2a56ZEaWtZ3tU2v8gOdfdG7TBVWCm90qeR
a2GqpOw5ntpYDy0DpV+3RL+OAizotB3Xaela8ck6LrYJLQ5wSis6hkAqODCXSUJx
MmaCa2t28emjPxFDHDTb3i0zx6LWiD1PkF7l1iqB5cluZA6pb2Tb5TB8MdVPl4Wr
fOS8MTZUx1zFm4bvKWn7zgvYIUEmgt1EEnnDVoNigMaipNE71wRcQ8Au8U1Qcrop
rJiXp+g4tnxn2QFc8c9uqMrAAWdOSU3z1S/SZfhbSVLqeTvyT4N6vID4IYbZ7bSS
oLUOKmJbxzX/nCtKOZcaE4iZiGvKP/P8LJ4LBRCUfO6l5tbBvkrxVFFhH7y9Q+Sl
Y5mVNGCzzNaDetZiWiP9DVmg4kF3fD6UVh8p2yrzPjmL3jRbsqtvms8qjDbvskyy
2wEWXgL0VPrNvLmy3gFQNu4oUAyqUxWrfJVAg1DvC3lPPfSBZfaHaedOoakse8jN
M/5L0mv9dfdmsvaCqlrAVJuNLEu6HARIZgML+Kv39ktmNAx1oLhpshwTAIGPSZXr
n+iUXLeI+KPvHOmCzlaeEetZ1DMSsEC4lVLMFkX4Bm0R5Ej95GtMhcl50oGTgJLZ
dQyol8RPdCGRG8aFYvRQFWW9YEeKx6gKohIrqMFFpcPwj6PGqXbZf91SFgK+5SmH
aB+db1lMQiiLa2OKYhvJzErv4BGQHFbtEsFM+yI0VkGuVBnNVJndKTjYdMNygZS2
MfxHcM2PcUXpzeIoL6Z+b6MV5jrwcLMXUXppYD5RiLyNMd7Q0+nN149/jMjk7x61
cor05TR3Ink4Wz42ravuU1XHo/tIkxu39Xi7RIzhM9Tp+AEHu6zOvZRf+qBeaMpM
GZRhz7Wtr8SD/AOztPT/DtXQ7RoLOE5bBNMk1RevVcmcvIUOn0J845LB7leSdo1w
S81HhgnOU9tjsWgGHWhZWPmsJ1IMzrLmnWIXPx3i3KbDkg4Gl0pGrhr3wZ4Ei7lU
sYzAY17MgRZN500Dui1TKmytMTgxFJ2bXdO0DKlkIooN2M+WvhcSVyRtCkrxKSQE
M1EcbwnU0rKKxaGGhuxlMjy9xlj/YMRs0VRsGbn13ihf5dlVM2qSr8rWuhzivtG/
D0ikoSzwPumbhKywwHZ1NIzIkQuvRXjHCY03+O11eSdRndz0L3sJBOD/WYC3HfS1
XTssncQNX9+w2kP6qbfHAovUmau3zfg4ajI0DJ5woIfGXXte/mlvOqipebKeAqgq
ncbUnOQRmGgRxQPIxxxAT7PepII+6ceRUY4hnEKVbp5ZkRQiS7c9n2xQgnTnA0Av
bk719RZLcsUlPXKJJCPO/16TYCKBM0sYyOpJyV84eaJA099qof7Xy2FyH6lzkSXS
S7Nd46pqW1zZ3fn5VZLFkv+cVck8aBrUOYmdgBHi/qxoZ3ohf/EVeSaiDWCzO90N
2F8DjVpBT4MilW9ia+qc+r2yEy489mhL+6ufVz2Tm3oofwNOJ0+LAZ1svbB/FXGU
a98hza4aeGRPKcW1AWIuWm1JbsNabKg7lWsZFt2WzDBF7MAfQFu8ocmTuPzgi/S5
ilkNw78MCwE9IKHRES4xX6R3dC9LIA8SO9hkyKBttUuSJGkwcXCSkG+1vymwiRXe
A5kJTlPdUbZoRq1fzuUaWf8iyDZRs3bzN7MIB/FY8lQa9NVRwDeCPbog+pTeQwI6
HNj0xZn5w4eYjLPVdEKb1WGFcuQgUwlLWo2ewcCIE3LzwGOQR4987ueR/I2jZCHo
/hMKzA00kS1gYjkayHHbhN4APOSjcXjsiXjbKFOlfEXZP0M5COq3kUWLz8p6k00A
3Uxfm3nkBrsIRlvmoYoQ7mZ+xHBJVTnEJNowyN8Z93eTDkjaPC/wI7XS2WWZA07l
VqqWeuk1XX3W6EXiXPIfPbUAuL6RwGrR80xCHtW8wpxbj60U2MKkYcKnhMy2LB2p
BDvcZmSnyjU2ISoxaTL70MTP05kqIjawPRteUo0JsOKbAVuw64zNiTnw5d1O8Ca+
2veVjwU4ITtrSS2xMsQxqItapkfZcqoyUQ9pYQGBDGG1+g63j3R2KF8n77FIQOiL
mqPh9DxcB9ZrRa6VMy/1V8EG8tjCA+X3TIB+CncOojdBW0nIdghntJD0jQGfVu8Y
EcxXU6LHezLRnxD7zbYUpteabRRHmVEUGtr7mjvC24myfWe+1xo4wXUmH/K2PgOd
YycXhIXX60N40YsFEy/uoWsNodt10C+1liit6Ho4+LqOSAFMA0kTD65csWa+dWRs
R4QtV4E2I7hC74Pxn5vCRDT1M8w7261KZJnq+QpbmCEAukDsGSK+oBoljQa+xRE2
dXGFgvvHMKx3T+RWUDqu3v4Q/hUsS4NUcFukqbIy2uJ8sav06eYVd+H2VH7dHRNF
crC+wzk1MKlkwm57LJBFExlWvobHjiApP3pssve9uQFRULkj+Z/voXv08YlNl6Vz
jsVmxzCdsX4Mpm3nW6/xuWjIpuDYUW0/IKXrv/BV/txY6NvYQqydYiL1HjtGO1Kz
upjOLSox0ypZQPYhGhebW7P+IrySz8FUqppz2JkarxYQY5cy12T+roX+hF24Ddg+
FtHh7Q+IeJ2drSM3PxeoRi1oH1LUn0WxNXjC+/max3dIC6pprOOjuTk1NGi4+qxh
m7x26A+CkI9LCsSIi1+bJik+3Mqg58WgLznRpPYVQeIXgE7+P+qZlLKP2WUr25JL
Cvxky1ZAuZbtrxABiZx0sJ5MlBBrsr3HczaJIRz8IAWgNJzLPXjl5W9bvhcSiTI0
h9dfMXHlRv9ZGT0iT8Npx62lH9vfUIsfQMGwDgWRfrsvXaScmZghjQdPGBgsDh97
dS2U+lhDC5CSVioGtmrEth0ASTzvML9Boo0Wq26QK2NOrD99CPYYcjH1KkfQYqFl
hiU6Znn0uLoQzdp61mcsRJi5QnwjrFm3g0bshU3VhQhX1CYl/uRL00aObLfj8KCo
QQYkkvvht+dDPHeDb4aPGyNNBsCE3JBhpDu4wU5J0A7JfsWCzc9uIas45woDo85T
TIJWoDCBT/d73pvRFDP9KrPZ44ga24rgX+zbuZ7HZ0qDGgkJP89BKDZvdyo7w046
/HDPR+xXjw8YE8mJi//JGcM4Jpki3esJ7POjA7L8NG+jFqBTYGuHz5+LdxP366WL
gFc9KRWUaakrftropQ5ENqed43P3FkL7TkMaTuLLhHHLE4hRudJmBdPbOK2JbFQZ
Yqa1/U//tE6zmRPU+wEem0kc/CvOywoAAVdFqnEo467UTrGnTyG5pi9qLTLIQ/hQ
O6SVsJRPWfp6ctA7jCoHvOYfrO0ERA4IT3L/MKqZXGH+QbJ/j+HoFP4il88MW+T/
IbYvcX1G/6DcxuYNX4hVJVSRXf8Q4sh2gImCNvo7LI4SAQOtEmkQttN51EQ1zcgO
9iV2Pp/QfU2izPkFWGioHW6qJYmrzmEvUfc5P4r5q6O4appGJB56lLIgZdygEO2b
dGZsaTMwI2bZ0CO5k68i+/kRf9Tl8TJJyz/j+/+Pv1o3ziMKqkD4Roh7EHbkWawu
luU7QIApLvlUxJ57atrw8AxMzHzo4+uPkeNFjOR6OBn3pGUgd33FRn+HdlsREziH
GnHx2mMNjI6Uxfr4XIEOk7ruIe8wvlFC1XCakr/O/y/2+lO044fwIOiL9MYsqBmu
C3cjJeyM+0F84ed763ZzKoONfR5dLQX7gGj1h94Pt87KAhMGhhkemKsEMY+4vWE5
b0MGGKrVUEJdChWqN6upopvq7wtfPFrcslBxpEhM8wwfMCpYP3dPsjV3LodHZiGO
fxEaXzxa1ICSg8fKK9FntaynAq7EqtJDIhMQd87FLjW2qUMyC+xJnwpxKCe0Be4l
qwx86wB+VWa130LqIbRnr9DntJK0TvU8sU9FUznevd7FrMOIEXnjN9k/sdNd3LcR
6e0kODePd80iCEujLkrUFJxaFMKb+PcrHw1ojadZDftyJ7MBaRYuWoDoJ4CdQpzP
rWBKLl6w80cm7BJGW0rnA3aqDDrf2Yles6VkTSk5tKNxl9PU4EnxpwgkAj86mcQk
MlfgotoZYu+KnK8paObfnuAu7gLVb/NAHLp+rDbkLA6grBtgDIAfxngmrqNl+kmc
7uBgKqJQ3c6El8XXqLWNwyzNhtaReM7/5ICVdN6zfkbUZzFaNOZg/qdjJcZa5AzX
QA168jO3qViiOz+xEIl0HPA7CZnGKMtFP5FnQHC3DKSbZcu5C4kvHxVA0hmvxGb4
4lQLwa84xp5AwoDH0UI5urr51rF6s0OT/hrx4psaIPuOri9wyF2K1N3JcUMeuneq
VWQwkE2kAsc36FYF0M7DzjwMRiC+9XAqJNM+2ebi1zVNcyBZBhk+VgxTKLNt45bz
38oCoWS7mUzCL+XPxybOH9hU0518zA35oH2rLCoKJbiicIZPY1FOu9ZzNd7bx1qd
l+cDVPIHytGicv+pkuzWYA9RXeb3Y/5tBtxiJLFltjQft5uuWTy8FdxCXIBoAxZk
hgqkiYyhw5K8tpfgpkAmawKWDP0BOOO4R4aVd5mJpqWKiZ3yrEUPPHhDVeAPhDrj
Dez0uWHgzVJ23vSzEnY2M/ztcemH8p2+VSakkeJ8zApGyYZTHd+NFbmlhkAGzMGL
VwDK2tC6KUFNjlE/WQI1SZbliG5/+XsS4ufKn3ipLLR8I1pqTgP+D319rZjRUYoQ
EHbpW3Pb0fshoBbOukmfPSpCvdxkQKN5wJHSJWP6HcugVDdOF51vtXl3Jugv07Gm
gpF99bYdd2xA/PjihDa/hQS892867VXtd0h7l65FrOjh/73uoDdkyxSDY3WclpGH
xkY/kgFkTCYLYRvFSOw/AaJg912nwCV8kQmqcTxveTlL2jJ59jdZMkHg9iEP4qEw
QXIdvPYUF6NmC15r5FKeNw4BZXrIjRF2Og464VEdOwHjxeXJzJ8yDwuomISLxQLw
8WS709mgpn/lidKxv1DAQNcYZvYdzyaBHQdJ2/Yh4dCoZ+ZHI4d4wGv9WwvcxB3F
f7aPSrpOhihBkvbyxJEnBeyK4yhcCJkC8GCGv5rPT5yhAA/YTkxEHrRjrcHpU2af
SzRSSvL3io84MearsUipSrfrjy7Ih702PeS6VqY45BrZxyI3TEppHVIighx6M92q
Kd+Nta2TH/Rn//sDkwMa52hdo0IVxsKaDfBA8wHULnn367QWZs+C7jItGo8MFLgF
axHO17ei3njCHPGtDIkm+xV0SKETm3n8ORQdyTBeC43w5kdRJtUFXPpEiKa/xA5S
h2cA4/Zn5dfE5qetHqWFNvIU16W7fUqWaFl6wK9NfRNe5fMtivqaz5L1tO347Fsa
sc7J9v4G0xwbc613Yu7l/lazlEkIU6p9WKVxp+4hFCbRakKbRS2jYjFmM8jrBeKt
RHKCOqIOlxrT6GiyZSUYVcpMWZBIADJhbmDrblWclQ2Xky8o7Bh8pB2z6SmYPTHj
asUCob3HgTCgZ04B2IfrLluUDSinoCQNHmfnrZZtUa++v9SeGnV8pOQ/8aK+aduy
1Cr+91vqyEqSj9yaW3OiqWxWzb1ps6GeaTurcZWE3yADQOpdjjxMprBK8aA5elp5
YlU75ipGnvefV3GKYI9KvYWyzc58YT4cHCdsjH+fUXOEitRzzLfmuEmWDzVyF39Y
doMGAE1zcGWiycYlxz0HKKI7/yVE0fKEP3OnqvnDAFyT6b2+5cZExNBqVt/T+3RZ
XeYQZPKRjwWQEKgbOZWr9OMywDZIpv32bcQW2b/iWCsA7iEBdCmllFcSl8Gz8oME
hTExJnaVwCDTv+LV7Pv4Zf1MpbArKTnlUKM+Ml5B15GXd9BnZXvqolvoYhxnlCtf
p18im7oO6Sw+M4rxOIu9GP7/8kF4npL/jo+2w6Rr17Dh5dI9jKlw+IpwTsM+e5o2
vTIEn0n6ALhrazv5t7+IcGKEABrR7Y0H2o1VjmQI8rJZY6UJEwLidJAMY8/961h4
asWvRLwr7/DNZeUuO9VRvRVXR0TGh2GyzMDCIFOJWVVGFWeOCMbSkrv5EemkBqXS
veTkRxCZgeeU/l6qhCPxcIaNPjM0/qdfofb6RGadffngibzB+3SQ4y3LNWlLYM70
3Yr+hOt4U8nTJxSKg6/i5HiN9vMeJXRyYM/h0Fyb5srrUomIAEpYY0cJYW7MZhYo
67ObOKZwHrnun13mFJ1A/G5xIzJMfvitDRIJLKMZYoyH11iObzSA9CxGemb96ytx
1g7jnWfUA1Pvsv7jNTXLaN4XI9J4bRuP4pfwke0SHPCRACQPgUxavww2t3B8lSG8
5luUI4/Ueyf8pPF26GdBuAHfbEaH/RN87RQOUt96VXbW6hGyNpp2bg/FCXryZ5F7
+4a1/VLRlTqs8twaeB4GmYyWH+kjpZFtEE2K3UKm7qo0pUeJRgKFNRmkGfEaLM/x
vSU5JeXJBvUSkQUgruhd759COg+B8IKUvNKe6mHb1FNuZuGWE1Pe5zAhN4yBSevc
eTWNevwbvPwxn4CL4jn0SqmRqm2qAN8mBL7kRyFhZBQtyIxRv2tZ1OEsi6kDxcHg
p9hrunIBXpV0iIsGvLxPOrCDYktTzwO4hq0euPrEGyqhBG4BQxgcq9/sGRdKlAdX
I/PgSwm0mGIhUYi2CLX4lDtZ199kyfSguBgEeZzrVxZ1bB9+PIkI1Z2Y3dMqmIRC
bdJryPPI60VLK5UyXY5x9iKZQi94bwNeE3yEW7whOxAAlHuF5vRcCs6dbK9Hnjqz
Txfu+pOMap1C5Yqv+G85pM9gZBmpEOcxo1lsXotMMJuJy6ZqmHC+CM+CnmHKZ+ke
VKH459tINjpCSzmtUSvAvcF68YUt1cuhwejwAEv/4GOFM+ZgPQCm4beSYhHX2L9q
NCmVJgyV64V2BFaD8o2IBEnYaPh2VgOxEBc0b487V5lFzS94FIlTm7WS9799KukA
YeyCBn9bSz6F1STdRNFge5U4cTFMPbUpsZNJf5aROwIh4mVXQr+D6dGz/auc9RM6
I77Izz/CFCPJ3JXhtzopAh/7G96fBM2ItZF8S4M3S/PWdS43Wek/AM3ORIkCxnny
rGYaujaSG080fxM3v8k5K164P15urP/791fa/aAhPKtaDymhNZqmSIST5rR0To/8
8igrwYUICSrGMFIccWnjFagtDmxz1A55DGjkjPhdLwtWagXhFnjhk767Lu2zFRVw
tMFt1woRkNilbf1BSgMb90i4h1O5NX63Ker1paKIU40gIHkPZL0wZbL4VGdG8n/h
0OI36Eavq7LePjiOtNWc1S3FcFgAldZxLPTftg/oEZ6cRhgzY2fte0DZXAB2Tjdb
dwNMzuf2nglv+Vg3TCSkNOfUXJ6ztrQl0+Yd6/UOdDjNp5nbult/B0KqGVC0uiHk
OLkVv+NzHqkmr94YSiyuwO6WkTEQ49Ogz3lAgd7lJg8B4EvOTYjtRBTyd9uTY3fd
Dx0EcVCEXStnjKR2Qnc8R6/+428KW8rV2QlG/zlYPmwEWNblCBzKwqpjD3sT41kO
5YK5t5mEzzww/ACIOZvdyAPdu/EFXg2H44TumtgkSKpi5JhG7SX4YukKKxkq2wGq
c4u/3QsbFrRLLelbQrwtUwHeKLoHf++kGBriH5mIGftffANrbuNRykiglNYnHlRn
weAgYOcujXfzz7jwRhfu5gseoh/oyUHNW5vMJ0Mem4ivEmExrfpNsIsI6JFZlMsu
AED3JDFGR9bom2FaA5ENfKHIFKe/QQvTGqyyhar0Er746bI/hqRwbWiW2kthvtlN
daK+QYzeH8PY+d79G6lZNEvxphgQ7O5fB0DyvUf3x9jRSqjwp+KGy65uFw+UrPku
BU+YJy3nrnRBJ+vBO1a9WC15Uq0IM711wPnvlbjc5BgTF9xcwroRJYkcORcCVx9C
Fl8J7YYoKb53v4/7uzAEFsSp+3V2q4/Ajfx44rcx5KT4CAm/4zPaqEiEh/RDZbbf
9M7o7KaVkFoMhdWhMfffHZgW/EOjCr7zxYZkkK2eFO7ICttkmHh4rjgEVSwiTQZ3
Dy0PdOYz+T/BqMTA5SKeWwbOjxKrmlSuUi4xl6O1TMP0WuM9erdfhawegDgN+G9d
UU/R2u22nAwa/zT/k+8sHxjE4Gg8ii3TXK3fgMelo4QZ/JQtWwSxLX/iHtEnIyzz
hdwQyH828E4Yum3rVsZ2kbaAK3KPwcOtp1a6iju1c8LNRcenI+VgPFm1JlDyzC8V
Vn+3Ps031yJIllvxHtpVDW+wM/0WF72Eq9L0tmf5M0lNlCNY3oMEMggzXMRROoT/
g5PIQzh6XnvIS2GgQwnm35suaCiQQS0q+PC4poaLttP53t5JJj016ZNwbGpYvUzV
e7gqLp9Y1A9VBZu/5XfbdyPJVfOOakKCzxR2NLIAQiWfrCfqfYW+udiTn27JbSly
FQgz8nh19cKgvaBVlnbJReyslFvKJmAGemQqK1QCI4EwFjourTwTu5P1NhoS5t09
WL9L0x9FBT7gLzM00QzXkbwBspWkPJ39LgO/3rumq6Eej7i3gSja5macmJ6/CT82
lSMVIxhF5g6yDH8PXQXwm7ycOZpPaoCU4rkHcfYm4wzv/2Y6t5Zi9V78tZWA3q+Q
CxTMRMTVtwOfTDPOlUxoneBBvdnfD+yNXdy4qURFzsmOUNr1NhvMTPuZEoOc5MKE
mgd5UtV3PJJNGN0OK07FA47nyatTxwIJsO0e+flkiSWc5nXjBT3umGdPkewdeftl
xqFTr9kFifMZGs47CWIUkxcTLAt3ZK98fu0yh5XPmUSReayDXGXuKfAJyiGewJQe
6czmR6qsFIAFjTq2VrYA0CiunowzhjuBUa51YPfOezX2tz/FmUUBoUryfdGXfXmk
1C+BUtO/8SP1PXoWh0bTU4POVKBfsK3+xI51p7/r5npbAbUpVbJs6QZOe8eQdDfu
9XspFuRBDczRgpeJYcOSZSlyiP1b9nxVZgFf7AVBeDhz1OZNeINZwKvE/HODVv1G
dk+62wDjPOzttJNlErRoyPtsQzKRLN2AYjg1E8y9XGQ74RP4wWMNFkrzlenpAKyk
38EtcWMFCmuXabbLjtnzNdBCgIaz/Vtz8qSjRKm/1aN0bNfy/N4dmGTwVDVq0hfT
cGGoWZ3ZrcqAbs0zzFylBupF5zk9db66iBeL/WcWZeSLT85pyttpD42OglcSUct2
enIMaDucmWtRd9tBFmghchk3vhuwEWWS8GQ5RjiCZkRFNrKEWagMqZRgHGl8HWag
2ayRK7uQaAjUZJLwQlqtm9WPASrWVl8XzlGMWHE61f8kbaRmhNPL5fjxHuBlveIU
7Z3ZU+hTNzcdJ9k4PkY4HHdCTiFTKulHgLmptgTuT94+c0grHViuaM70MIc1S1cl
g0JrLlVgfVMLF9CVTADZZXgdhB9G/6UriDsTimeZkXZzipSlsCGDvC7M0MDGmkDd
sg++GEN7AplwzdjeZsEvRBEaQgTR8j9uB+1wSu/C0j/XXNf3/BqKQ6dknnJXskrY
QDeHtiMbqqSlU7pDccvw4v5VicBEyTHiDxje3Nqya4ZqLPb9qssSmIJaglW70GIS
PT0KDWEkN96QAxt5Au7IZZWO+i63zZBJRDm4ofY1HVOPQrQhzurHDtQwiIOH3a00
pjPaS4knrMhpqucqjsQEEja9OeZQZvBbqF45CoYtVzVuL2UFPJxXd/JAV4QQn0PC
1fyb1/HwyWW4sUHSO2JY2yQZfecXScdhfgLQcjEHh1ZQGNjYeOW4tcY28uLB61l2
A7kUaHIqKvVX8eTmT5PxYVfDCDGdraTDQd6ryiIDHAVGmHR1hhG0KX/zly0S3A8c
6MsS0SUNoDv3j5thvylzbasqSeEDJMpkqOWSVatYELCHFAsEKKQrew65rgN2QXIB
htjOXH5DNFAilPXj/dtvMk9OIGZRepzmy5D52jSyW1FWQkldUaOkDZNyWE5of0y8
SAxQ3gH+RPz8MkfhalA4ZIrpcgpfWSGGtzDsqGLbZ8Lm9ezSc/PxG+NvaMX2YHpn
nXXFaxXLBDRc+3rMoFMjqlsFKzN7oWTJ33kdxHfLLTpOxUYXL0r347Um4v9ifhLk
GpN0dmEzRCG+1IySfWCcX7sAApOkWwsLBSHyALm7TMqoYlBrbbIQHswTSWunzQa/
0oSCMP2k/FCTmjI8iAKvGs1eiTjPdHc0FQoloznIlUJYAgbGsnSIgUNPsvmlWZrg
/NF9Dhnq4p44MCECtxvnLShXz0g2DjWXpVdTJRzbZy0HbqZtG5tmmyD6YBm+YqzL
yn7Cp2Jic4MnLsMGSlEC3hKaVWwrf1NQjakrsgLf6+WgLDKHZT5K71JzFGhHHnvP
Dh75NORpvpQK1bkn/QrmuzUQmUXx/PMeUN8r4yMh7S9FghMPFrPUTuXbz6A9g2Dt
Q6ArVTKKYE7SrSc4zyt6ozUXuoNN0KoTLv81do2wSGX0BOHBUOT5heBne6RZEuxo
/sGzGkUElIieOiPB5Bd+/qcbto0FR2lKMaEcBXuacpSqBeUO7m9q5pzXgMNSucrc
fefw2pQlGsPlS0OoP7W0E5QIuQEldlBaGEWwULNIxob/9TRFcashPQAvuHjiBS3t
O1bSGKoylPcbEMFmebzN/HN1HyiitbedwD8AVvInQp2AiSqaX++5bWRKWjcsKsd4
JQPIPTeuS2YFeRxNZNT/55dozOCkrqKvwnV2mq88Ww7jsRVDu0ILRv5iuLc2Mjwa
qPXQiy/5XkiQQoLAa1U11DDUrdMnrPpXYYhHRnOB8vSQJg63pR3uXTj5P1B5mSBf
5w5jYqaDUAGYXx/9xT4gshryC8u25pBZRGMSYbE7YuQynV5yBxecgV1ptAx+HGCR
Ry+ia1Ckw3NT0sRfuna9ru0yOodXs+CkXphYRLy0Xer0jDMkeL3MPWWwWdK/ItAj
urus4zCY7rrFMwv32PW/r1iGiqHkztn8DOqx0C8o5kieE2u5RUOqruLv9x64pIzh
L2BBWHYaliCSQNwc8hHKuCFdQdw+n2mmEW8sd73jGDMSIfPD8yqDXHnKKHmzD5Zv
cuEVnrDdrrAlT7TCNAnhMzCoi1pbrA1XFb7BxARhL61mUe5A8a5sZx0jErY4l5es
3ypcHVY/idruJ43ghl9bchA5fiVq/9OGkAF4vfFkK0JR9zOlazzEOiAY/yXWPd8H
Q142f6FS8MPDzJ+NzttPvedxInNUb/DMfgkIT+NYSQQH4y7xxv+aQfErpWM1Iouv
kfQ7D0UHt//WFIXwvUu5EzWNybLifZWbkm8sQvruU6Tjpzm7lP0Qe6UG42c3qHGi
IO1i0W4HSmSkJ2JyQOpcIkMpcBMIrDhjDyoRCG0ZmJMNestoazGOMi9L4z8UB2Qu
xNGqugs6gKtt+lieb0LHyNcL7C8W0pMw3adHIVg2IPa7AcPDGSESCt4n9Yu1Hbl5
PQ6001EH6Vxlhx4sSl729na/nD7hXf7F9X84+HkQFSPopvRfJoKsENqYJj9rxIJo
ceT2ZCw/tbHTUgaBGe3/NmvJbQQT4sBR9fGmY4JjWQDNFYsCrd+NHVGXtGSYT/gV
YHc/Gl5XZS0JNbOKE6/KUquonzin+wr9bKwdkw5ux+Grrb6QGEfJBijiVCpNmA/3
pFoQwTEzkMCmmyCnccghxL1x2h4oe3q5zFqsdlEZmX2xA/xD74kMC2AmRu/4StTX
x9RX5ovF5/bdzc2jZcbuA/VvrVcrEWWOHeu8O/q+k6J6WSDZtrjVsz1a7KYGYJkh
JIlG/x8Ah/OMGfXpur52EqRzOMbufaLtp1Nut1OpLqaYKhlXdsJtcVVmClbzFki8
eAeVDbI9Q3WGOQuU+v1xu2qd0KU3jckF875Wx8KLv7DXbw6KlNkmuU5uuKe/jZUq
EVX4uxS1k0ReAajHe/RBiaLkC2KhpucwITB4W+T5M0ezkL+mE5CS6oZjZdixfPKR
zSszmQAAra0fRtrJHc+yNL1n9gkCWuSmfXDbkl6XgsTerKyHpNUOidN2Bs0AjSQP
Yf/aIXTJ6x5CAhj6ejTNSYEdDRR+gdWxC7L9+TFi8fV3eaiq0VONo/YAqjHauFPB
1qwKvf7g24Yen/6yoXYyZRu+tSwrWyNciFsEk8CxVkfGRzpC/YkH8IZTixbXGcKz
Y1ad6sONDjq+82478lysbZ02srgCGjhr9uJGWsrD21R9Aa8HNRcsgXj/Avg6iQs8
+g7EeMucWqE/0owM9PjFTXVPKugQDoZwHdZEll5OCSUK/lKxDFUAaIMEd0JvuFNI
SakrcmMmu5AhJUlyR2zpp3nuRnGHa3ZNTzW9kPxaKtz96Ul6utO2J1nokZMR+B8I
7ypL6eLJbZ70HRizN9+5aid90SDVsyyql74LtSovUhhuwmugarjPepxsZfYFmKir
P1F2gSCMcq5Dq2yPBelCylyr2dQxl5avTfeCI6g1+SflSN97fZx977UPvwASef9A
lGDMyqnUXdbkeiOthQ1KOUx48x8Ace8IqZIhOoV+i6ukevAK+eyHZXiU/8NoSqC+
QFkT2POVj5SUjnJdAYeax8IkMQXeIWrFb3FU5ncL2K4Z3M1ZauD6zkzkAsHdrUhc
00oYVvgS+28rpYw6yvm1t0Y3BYY5LEa8WwEpFWF6FqxsNVoBe+kY03XFsG9NCq/9
7i3JLOl/ijwVvG2MPz3TDkx+/TLW09rNh8eMVdjnLG9BRG8Ae3hC1XA4lQNs4g7n
baPtkjpXwrieqEJJxgaB9a96rt4jeDUPzaSPCwEDiCwZrz4cuiB3pgGaUSye+GjC
MwlGZeyXKeryCjJ8Ho2pjXpNRRP0nKfR8jyViZY/Sp7snDruuZg/FgT4KMFNZD1g
TJLtOJTXcroAzwDUYd02SkmcDtB3zv6b5keTVzk5wm9MuDeHo+wOM1ATiwY7WpeO
rBbSiTcf26fDYv98lkBwMu1HSSraivYDP70tsGZ6A9TrnChZLOiAC4i1m87fXS4P
MBKC/hAbJnGi9rmQLEVriG8YVl8cUFt62Z3jg1zikSrCOEfGuTUMPygpwdGAE9c5
2ex86Bzr31f7WHICtiY1mt/69S9dTdPVOzvJTx8ia1OxD3CI1lXDYsa/UCEBLGAV
5vjEWWKSe2LJ55gZvdStofD4p4r8tfKXoqQ17VTMpMVSapPIKxGAsDYt1dM5p1tD
ccPCsIzzZA/5OL82rP2gQLKDtvyLcL0CIf3oU31YxEe8GS1Ug7jEEhu/AWa3WpGw
2ZSuGTn+7buLDZM2tUaXMJCsRrOkfLMOgfl022nP6ucbLSjyztLiJa1uEoA6xLpw
54SAHxoMTk7oImCeU10tWFB1uhIuIFkKZ66Zi5nEdsE=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FLcvNZtQAChwZRjZtG48k0vR2S2dLiDNnt5bI+UY+z65lyLWd3+ak2qWWi+UucGI
5OCacMUUmK9q8qbvGSqxC9KYqUJseRaxQ0o5F1k51sJGBvcICz7usZOjvAhNTAtE
2RpHaZJvevbxQqzQ6cn9dR1tMfg/XMYQ52r+QJfCDGv+dXXNzjiBDFrH6KIR9S2C
BKdCEuYdzHFyPdpkYcvhb38yaXw9d2olNemFdHYO6jZKTPlaoI5uSFI+E6lzZpNh
xi7SL0ztKxtMHh0f23HP5EW66SpLtN56hcGkNnjgTHR4KmYpatuUQ5CGF3iUmyyl
x+LsQeJvRnVZuDJKERxVFg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17376 )
`pragma protect data_block
2vaEDtFpsT/O2lNt8+9S3kS28tG4VXyE8Mz7UV5trubwQWhpvysy19k8ChB/uEdH
K2f4GSDKYu1LIjjgSPfSAR+QbpUiySi0D9yc8CN1u7eVOKX/8ESLy2i7SmWf2vjy
IDoI/aVa303udfxbGvfDU68zhPc5VNLP77igz7WciNxms0wrlE504lM0wvusAD8S
6Rr3a5dUfAqyyt7uY1NQWKoLcVBkV90anBxPOjZscMjDknwcmn78jW8+qvOLKk0Q
eZt3DlXVHyG0PsD55VctTQZoBspMr7wBlfCPrm4Cp2n0gOgOgFz1iIlpDsPtW8PY
ff4M9e/b0ieeP15RrKDJu5D25tfPa+nmLuBhLSUZ1m5pNjfJ/LZGlVdI0WB/UzJR
VfuWskGZ8ugnD9895JEi25sAOC9cGojk/sasjKcRHv52GIVbt1+xTwhmddRLiH/l
Eg2c8Ei2prO+m3YSqPNEaNbUEUCWe/BRimLTtmGZrIOyJ0sfmgoFBTSr5L4zdd/x
DWqVHCuJ31Ci0E+HCVnSz7cwz9ffmiidvNv4xuBtGxvDF4pwfE8GO6ZLx6qsPCfn
eB7sWp7Hme0o3Rw7uh98dQFWCHxkCknxNTHuQizWfSO3fXJJRPn6zc7YXCY5C7Ok
NAe/b01Ae/ohOX6EXspozGG0zTSlkopVIqIKMRWn6LTuRoqDWbOQEurZQOJxvG+0
u6pHBOzxOtmmt76SvHhCdeSb4T9GnCW6X4AnyB7wlFZmfLl6CVNLE8ogwytgNfVd
PmE409gDdZghSs6Ac06dKSee+naeKzazlYTc/mIAesD9YKn13fkQo9ZY8R17GbI1
/aReJx8CmIRFKR2LljHoUvF+p6f805ypjZMWI2X8MRL+wZlgCdwD0s2sUCio3riE
J2L89dXqDLP8OmlgQaVa2T6KnTToHo6GGVdnWaFoILlMhdpNqaikdZ9vYQnxlDCP
hajM5HnaBKhdSTvVOHoNiAtRPWLym2Us5QVcBBxOyqqI8wUIBhbVnV5ABEQBQmLv
HO71LVwlLbIs67c8SLTEcGRybMVt20M2A9/8iTBDZkjIhgPQf5nwKl64w+GZ+7dQ
gigSKHBNtytAgfovfSytSGexmBsukRZj/zYVQz1hKf/AzuYeNC6CvChdlj4D5vP9
P1ijAPRlUICyfmZAmEhhIFUEll7QoFhIUDp6j6dGZ2OQMWm5Sq4K7lMZ/uROWWSw
nqU8RYXCd3ohgYYKQr4YATS3XX1Uxjk4C7fTvvxxGfICJhlpjzUx+OT0CmjIc5BV
eIA74dK5c0r0UUZV0d+AmOIm54YuxdEoJFG6ZJa5UeecwuvswIb5Y2nY36uE1KuD
hpkaIpCJWNrEDNRmRE20E+GNRJPhR1is14cmAWX0VlHBdKp/3bMw0gVjpixq4yaM
trHa9EntbCIhdh9oDmQkDCzaxpEW3Z740cRUviCmWF6XRc0ZHWUN1tvTFbX/vC0j
bD0c2g/CEMm+qzUet/4YKegZ/U8JQERPekdK5ahMEWoR6CF0uALm3LoprOlzw4NO
0Chf57E+XIQV7GFHpTaXrdrRTAGQ0qIfRaPxVCU8Xa8cSP6DI+v3JKxLWTvGQgKm
vMxRCUPlapywDUrs7zXkfdJ5XzVpIcP54GdeTiEmUiJWEqSgErsmJUNvgqY32RBc
mG2oWpbNcuax920w9Rt2MlENgAfV4Gwhz0/rT8j0HpEVmM4wFChNNd+T33kTRgf1
Df7r8taf1BD9sbCQC6Sh6aGRXU+C7pMICV0zC9CUOL0hugMXfNVKTQf2LAh5fJyo
/xDN8LQ1glsIQEY8+LO+f/M/dJFS465x1GLviQORxR5Pp61tktCd2w6lIS2D2irE
bjbIBR8xjzEPSjHneeyoNfyL2jQ4Tp7WsZ7VZ1JuJ2wo+8zx8zoT8ndvbUwF7e9n
L3iQy8MC7IxjC+r4NvCFCl9qv5NRd9nG0JgsPzJb8D3CF/v3XQTV6QMrOxREom7i
40+cGfc1mgY93w9Z9tSTxilzhDd4dPMRX2UINZS+yDxv0UkjKf9ddA7SHBaGJ4qG
qAVwZ4B4epAIoLJ8b3LKgzweGumG+q/lYDgIZETBsZyGeNZBI0TcVfOfa8j9gxSx
5AZXmTkx1OljdeKaGOkOVsjSSW0ovTxa64CGNst7F9eQm9ymQZ+EF1/zC1kLXobY
lHUnIkKdO8wuGnZIsDWykO2zDbAKYKHpf9sKnOlT8ofFd7ypBqftKUvIJJC+fuA2
QYwlG4V1j7ul5cz439QXtkWBJuOhC5j+VK5hWkSvuJTx488akP1auvWvQxm0tVEd
auo7X3f0vgJWbwE/ypslKlT17wCYNjVImZxL1vIdESGabMsvl987LD6Dxl4EUa5T
SDGyb138t1uFVf2FC8hWlEmjN4J6+CVCCph30KvXiLEzku6/yL4mmA4Wy36loLGN
1LBYCnM5nRl1PSqXTWvgEmiF5JEM9zNsLHM5BT3VPGV9zo794kVqFs+N+I00Fsec
JjfqYoYbZWbjSJKAjtIv/iViUJlsPDtfIDK5TWKpOhl7MRg5fSimWVM2o7N+RSld
5KbuUKDuKFhiSA090xyA47gYirMyG0mjDiXlfXbQb8XPE98JkTO1IqeqndwM/fZE
MDuh++z+b9H/E4REIdQBrS2CKo5YbOWq0pOpToitrec9C1YeClB6He2H7ps0tL0V
PoNj5jFNxEOArMl2HsbwOwwvNwQcergWQ2CiRzgV+567ov619GXc9oGh6IJyssHA
XgUQCOfnI7x8lycAQkkqmB10Py/RYTlhFzUIoYLYM8XI+d0ggTy7moEmm8GtiEmq
fOqRO10IHRU2Ijtka4XilRO7UcRzDE4RQJeYARMqOIxYk2s4EG7/5O/gSXHMD8TM
WSG5I63UDnM35AVM7iUiMdxARJXyE6R5ztQqR8myo5eHNuiHqi7rFb1SEhWjL/Fq
PdcUMMrI5U2jqKJRoAPZXy1xP0FdUMgwd2vzHbIyIgL9nxkfx8ksBtMfX99mFU3n
1L8ai/zDHzWrwBP6O5Ue2e/4NJqIDL0gs4iP18wGgLgSIRCefOU8nT39JPlozXdR
iNMJ4dstmi266fz/iy1pHBjozB7Zg+CO7gGgmDyyixZkgq5/Ib91U5X+wke/VCIf
BbN8NG108m/SeSAOGqPFHxBGICvqm4fFwODh2M6AOUM+W8WqQ0LcoN821nq/Ntfi
TJ27ryD2xerCT8LS9gf08pm48CDc0vk9aQKI7y+MpgAOrmF8myV8y8KGnAyyB9ML
YqKbkBhlrEx7MpeDsniZCXvARSOQ+lU6eIPn5mjNAC/6bUMIPe0+Lb7CwxRZQF71
8VxNo87JSHfAhUMiRhp8Xx2nchNBNd2lT1yAYJldWDi+Oat19i6c8aSO+lPf6fk3
xM/pAktQQzVXkF4LqWCaqJJNXA6FhDp2dVW9Skp/otbkLT+CqpaLWx2fPKXuBWg8
xetVGm/fo+1gKNltiVBu643Eh4oKWgnW17cSolkp6n8M2Ryl2AT7woVBPOvXlfDj
HzYb+qiCrpmx8tR4RqyOz/FWNm0WcFIeo6vLUsaBeQeZNtfZtzR1nSI4PZoGxmGc
Td3atVc9FX9FbMyqdhuuzPZRJ+mFJgAF7y4CZccPX2DHwwqt0OarARDOfNdwXkr3
a0eGl8y435dll/0jn9TitTWWKrAYX73S2Y6RFKRVqdc71KGLX6YWT9z09ORurTz9
CE0TCFeSRzjGhbPCyrCQrT4ozPeO1l5EBNsM1GL3R1N3YVcZt0npnXEJe1ogRycy
RMg6FI/3o7ro40gYx8Zw66gP1DgIeThHfVn4MD3TmkLqpS2W/ybDY6fA39c3NuY/
tPlL0b7Czi82/PmOoJVjkF99joqe28x/+Ls9atRaW1B+KWHSCvEfTCG+StOqpOMD
Oz+tTB8qqvglHHu6pJktO3ggqtoKW/rkeV527W6D+cg5n1woMvcAq43PcZnzNXrt
RSqPfqJAS5RWWCtZJsv5M5H3fkFTn4HoAVKJu4PIgajrBhqFnkd0sEyTM7Vdl4O5
ql6yI/u2oWoWHpr2RDb7ncg4Hox5Fe1hK9CUbvX6KUiVZJsPaOP4pmsNJDZJy2Ja
nmkFCb9SRitN1q/KCkkWr31LY+z1CrBL20KkuvwQjqz9t75PuyAS8SOfSKpn5eUs
c7ELj/szVMDsCwWagg17lgOBJRYvPimEGGWXQLsuOcYQDQvxdHk/AD8IefcnKamj
TG6APSSEPMD6uENBbbfx99gjUzhapcsjuFTlXYKhp7b4xiODfk3KyT9DzPP6RQu5
mBOFt+k/Y+EhY4tOrp8iVY0beFVKYRZCBulrrHmEZhjSISQyUrTxZWtpxBe17R/O
4DgAz/SyWpMtiuAqckzATHjq237OomXnFtGSPk+xZ6bS00Px7d/gyObdzosrUYor
NvkI2ZN3zeseP1NAD7B+JGcBnd2ZqMV5jdh4ijo+ydCUI5Z/Tazi2YcQkXv+dhhN
b5i997B7bjCWXyruBGC6CtzR8mPItDGKFVwcCV3lgdOT6GZohvY/gIuunvkmBP57
7LalbQGE+nfmZkt4UCumvvcD+dhyAwcdR1YCCOHJ3B2QUJEjf5k8daom90KCeHTG
hKOjoKI0Ykmm4g0wvx4RJvxT78yDC6CjGYJvpWtsIQ3FcUDxKu7IRK6mzheZJs72
XWORVnmVCMXzkmUv4oL1gGMOHnrdenuoSWNZvqBeI46DsXFENPjnkqJuS5jgqomW
mWFkM+hCp2wtFniEIav/UoGmRzoHPYwZCuWO78BOije+dm4xxqyELM64g/f5tyC6
V5snE7fFtDW7wNsn1B6OK4bX/h0BHR2CkC6cHdwyAGSjQDMWHx9gzjX+RTXlwizU
Mn/BLWVU7VPGgXnfItStdoitwWsgaIi1ErhxaxhbNI8S1mpanSdWqL5XOWn7A+VO
Igj6kQ4rj9JFZAv2AriywlK7FJLzizdDoBQg+WmM9/1mcj+iTFZJL2Ai5IaXXMaP
qPMZcOtLnwu2R5QZurKWAInIMTLd1izMMrspAFkfFn/PWTfOlS1xpDSuO60WLRpw
CgSgLZKjq1EBZwDPFKWuYxqd+F35hJAbOCXqY/N21dgcvOS9vGGsq1l4TrHg+n0j
sQdpcqZ24NxPVpKeE5NMvgCMy5KubZg13LMj6am/3oNtQQZLYHOJGpe6364p8+ku
t1wiWrjvDFJtXeylty812z+V8myrZQBa4N+lTUha+kartYHPzAnJgmrVD5g5yKoS
grtYTcK84LYiXrRp8z++hbGQF08+N9xnBI6YXk5vZfFPr8s93DUnSbVRwH0fTZ3z
IaoLFzxUy0mbjvrzwswKPzKox+ootuXthvm+Mg85p/8Mq5a9XWqbi/Bfk25DyJZQ
X3cU7JIXK0iqTEwSnv9B9CMqGxKiP76bb6M6M3AVhh2b9C7VC2jvMdGbQEbA/cGY
GeuNj3swmYOEL2jdP65J9POwxGHsltD99YkPjl4KXhBi1/6c60lUGekvGvtxTptH
E++JSVEbuQO5Pz81//C42arWVwshnfoUe6QoInzSIEeBvHT5B+koJAbS2O2AGswE
mohn5jrLMUYAD5NyeFPOhZm/tJuvNufj1++3Nsit9VqDQ3tIcHlOBpOQGDWfeD5O
iOWRsidp2zgNtTaBMgxw3wcUQ14OzRhzJATFJvA0hdRNph92ju+NyDp5KY2SZjmg
TN6vJWGG+aCKrbgdDO5PQwf2m2+z7+DBDKkeUTdBf9Nk7r/88bpzrgeg7DqXvaRr
nIydw5MacKl1R5+Ccok+FY0EpRY6oyJsOT0lmop/eNWdEpm3bUVIXzQFTKZycUOr
LWtmjIKP32qjeCXwEBEP9xRVE+YdQiUv5HlPaQ96qS4atfTpuWnn276ix6bI1xj7
e0tP+V18i4gAiCleXScu/pNGJl6Zn5LLhfmL1GEShHNLDttcCFvw714NHeE29x4l
ay2Xy0h/oyoD68s5n/0H50wceBkBJQwfo91hFKwkQk0AN6rswKYeZFr60ESQjaKJ
Az5WTTGCdDEOZlAwG4hDR7Mpc4qxH29hZI8/IKS6AuvvpRzCIFKpaT2pIbIv7dlH
IscudfPQfZ4k3WfK1M1l/IkVr8Oh7R9IztPhdZLmvxZ2oPEF27Ngc2hs3UGkZ8nH
nvfGRFUAZr5Zq60RZEw5SQVgRzPl2K7b/375uaCBSjYJd/rJbrkIXW9V8SxBZf7Z
tlUYzmTAaGuIlr3RB+EPkOn3NLyN989wK6LWbb/5PbZmHUDeQzsJbNp+WC/81IQZ
f2WSHdEI4MH5ot8jd2M2Dn50hzJXEG3ddkWaGQVhGCH8CJU6JJissPlaIfbztGJI
6ZyGrtbkH9qeq249NcQMiQ8sO6tbQqxEqb55Of2yItIaxWlRyHMnUBrLXBudrFZl
KvcjEp5AkzfFcLUUkzfhQqD6KIQWJwyoylCwydTiNqGZg7q6Q6cbAGyFK+AHoUOO
NVNFh8N+AJUru1TSIKK12bTkNeEBDLaVh+vr0abuJXKhJ9Wl6WSFQYL9TcaDBLPX
21L6xOwApTjVUjIp5Jkojci2EsYIM/cLAVK9qHCDVloJfRIaIpTSu87ZeQmjMwH+
p3a+UQlfo4ATu2JhOH1lX2Z4mEkjrtNwbDkJfx3Ixx21sNIlbamIzkxY8sG+1Bb6
qXpsD936HLNPajWEk85dsEVhtcs09OCUGq0bK+l00Sei2PFRQxfc78nASNh8Ht9s
H8HdJgnsvyRdWcWwQfcPc9fuYAB5gkxP1inR/vgMTe0f1YuLMrZqJU52BOLkThxr
2s1qt0eeCrNuoVkOr68IXchgM7Ce+BYlItbLQ9aT6ejWbZ4sG6awviIRuxL/vyjS
DFpesfJwO54utCxVmV3gQsfZwzJ43VH/OdB5pwXSpg1QbuuDuImlByK/a9QKDtSZ
v7NTilLhhCWkARErOICTt3qIqoh3oe+1m7FV/T3fluUQQap49cgD7zKpHqA89ac8
Ewl26vUsxWHLbZuqaHTFSZgZ36nvqOAadDWLPFDEfmVG13mESjoK9Txur7avW52c
jz/LM4VczMwQmi3bZt4aHVaH1eLazUr8z+hRdx5pKu0KBYPRomd4WjEueX1Vt5PU
r8i4TorTjZ2ifQProIMcIv4QCw+lU8iwS86uNV6hN3izRq194OMccuaHUF7IMImI
H9+BA47tmHSyHFzcXJ3A+d7vp80826XeIkuyLF6UIvkZE3T1aXFgV/hFUteWKlzr
N+RWzo5MtGwwkAKfFuhDusgojbN6Gdjj7Wgmw1goLLjYF9oqjK4A4jYvothlBdIQ
TbnZenbaSDdclrYoQuVKKObkn5sRNVlAT2wn14ZOebn12S2nJlki6/bQhvL+88ld
6UZ11NZM/Aurh54AwW89dMPGaZZqNzukUUkpLzgi2CMHnBQ/a/ZInX5KfXmgkFRE
HEGaNhSO0l3xFxeTcY79gYD6thp5LxqQ4gXuU3ZI0TTUV+Ep2f3YvSk20lzUgL2d
qNLQSuMUp2OPZ++fK4ExIpe7Q+WbjP8ygPdtnJA3mshH1+YluNn1YDm/XTp2UB/q
2oKWqbukx1DxPixS3tTt1Nj0BaTTz8eFwQnhSRvXTwx0L2rnjChU7SQ1eQu5HG9v
CU0udIFZYIPFob5cIjSE1KVcVptwC+E4FgU0ez9XCsu268kI2CrisvBsxluZHi/H
k1uE+ay433vhVHO52Y2GMPqFRCrGEeIKqryR3oayk0m2jzi01lZuY8PqXf3fdAgD
eXrIiYN8X6UdX45a2bnRehGbHzg/B4KOp5K+Ov1CxLRJMygx02TJLhZBDNWBmfpd
H0fpARYze2z3bPWyTl5b0NQFj3611ATwc0sKC/jz8jXcaVy1vNwlLkN+VUJS1Hux
F8gtdWHbfEFbWhopZgTO6dcuNVVxPyG8GXvq2GkG2xzZ0bqx7rsHaT1DV74gEsBa
czZ4ojEZriOxqDPFRq78gob3p4ElON6gZHVUjnO+DWMEam37gD2boPMzykXXbzGQ
EpHe+ghKUOaGq1ZUnSLCMxCKvFZK8hkJtzVe+/b118cxIB1sPZrVKSroqQBZq8XZ
9mposLc6wbJkN9nML7U7IGYESIW5vnpc0T7kayzdQdo1xVAVTfn5vBPxammOBXOQ
QSR4aOvqI9o49nc8OTenR/GaPRgnIOymS5gGUADkCj+s85EfRyWOdlodIrzBo6UC
s/FsmWx9+FhOQNJRFXAZo9PaHTGtBFCzDiJ1fUf8fXC1MUsz2B4/R57FuMee0zKV
AOatgc1cqZXc8pSmjd64D+cJ7OfvlxRMAN0JQxrCMrF+mFAHZFMYkWgrRyxi/AEg
tfZ/bfAlAmZzwlkx39MFwhuUsuQQmAgHIkitje2th2+WExrXQiBQlw/ST8pnRk2T
exAdtc+b9fe3AUaeX9IL+r+T6OJer3rVTeKrEuwymvcAtW4fKdZD2MecGOrfLyKn
0kO0miHSgpPE+MzigYxlxvKkhrgYiR6wfVVkPtPb0eJHCEbsAHvTKs49+o1qFuPH
SZrr2gtTE9hKK3Zn7ZezsgTtrVgh4t3AieLJeNyABcwYlYIUU3exbi/znb/MbgY7
RBpSNepNV/BgC33ZZRNwYZwO9dioE3cU76pLjOYyTMVmIZW/8qIg9xzdxQvpaQZw
wi1P0+ojd3SCzP3bq+hcHx47TKKOAmFeOHBwXJZlLuu2FtcwU8OV4Mb+MuRArJaX
kBtHAybzdNVA8hJ85yu4e6TSH5heutmdIIU9ZNQaRhj8Y0z9hwYeWGX9bI4mtyPG
QdSxVZwSuD3Km2AOScetJnNLO9TN3igSD9IAEPEYBr1OcQjU1dukKed65jBK6DWW
YebCANXrPXamE9AyFDevN3XzpxxjAEMUe7lWHZTR8jXITv4CqUhGMDtiC0w7e4/4
bcBZXceQ/+0lyxFZghC+xSvd9SeKvQvQRoYZH93vSB374sqeFuRbVd/u/+kGISFV
1qpmRzAHFllg/VaCpX8H+5tsIpyWNHye4XsoUSyBI+MPHQZCeT5e+/fSR8OI3x5b
PzQBXfplPJefXYsb5S4OdbU8w1Z2vEj8mPqezFFhHh/cvCEkFEx3k3dv6EbiJ/FX
g2wch+hpvMDBeqEM+JciaN+ZSNK4iyaqnSc6mt6qIxXXiOn+bPsKj7c3fsxL+VrM
v58jvHCoo/BeU3O/xricFlwlJnEjJVdQ6LYetbWmLYO0+JuDSzNj/rvHdeJK7sgO
ykojyH/z/tigT2NqlzzIkpzLJv/sJL4u+cqS9aQR05K1OYbEPO08dKJ62TiF3Bi1
T2KiyblU9IQPV4xtx9YYtG89DXiKmEvB/LAz8EIF8Pj9/gnW97fSbVp+ZOEETVbk
50G5GwvCsQiYn5BpMKj2le4M//BH4TJlMSXQF3O3PFpg7LznlPk3fp2xsjlnHVeO
kAVJQaISiGy7GDnUoC8EkHq7V1tgMspGcx/LZKXLl0hER6hzf/DgGwC4LtXsJuSD
ySiWtR62HwX5MeVMAX9N+RKkhFGVx+Yj9mnch6VbI3oeYy2uScYmh41JCWVfg2wc
herhq8dduvi0EmMBk0wAlOd3dv7PyS9oA8GJ4HgXiF+FM5sLCiiXXWR8YnobD3gi
A9TKsUDop0FmJtp3yl5mzvw1aF/c71OZ2Qen8NAfoOArlxofBHAq5/fiGbcuDaJO
mZir18xuFXpcweV3/mO+qQ1LIkW93s0YUCW+gYeOkq/+a/avRrpZ8CFjn98KKwl5
7q5HaJkNSWPRKOGYevKRQWdBnvZOmEP0SSIyjCob03XNK0F5oJppGwUBC73MrlP4
nUEPnI98VkMsd/2nyGVCnEh0i1Q88stPYxk/lqeHGf6s8Tw+QgKAzNwpUee9A0vb
HhPnb78s04p1qvXt9Z6oO0hpfSS8AF4Q4iga9gV/O+489hizAnUNe27BWmsdyrUZ
RlKUzXSZxMuZr3cC5UAB0ztYyF0eMZZzsyU5T26N5w8Uw7Y1XSPyuq1+zaMfqrvg
qghZObcTEdbHIsUn0oKAEv+1pSkMo4lwSKyvIqLYBkLzbDxAlkX7NwPZkKE48Zh3
6qB+Y5N3xBhHg+xxB1wnQAKZbaetEghFu82MIIotR4Rw7SnkKmWEy6QmAeOhYM0W
bpZIe8rE8Y2P7xRYhBG0VCrFSCMvF8Tvn54DCQVehG5GfKCidzFbA0xe4GFrtuUs
mq/qhjh4pEL6xXfZ9uhvrj+QE7Yn+6iOUqUeviZIt9JpqGBiEKLdLgbzOTS1GtkQ
n37ciM3Y/6m6IrTSGHkLin2vMotrbrt8sdcuLfDqmD7OZ73+4HqOKf/ZmjntECdm
w7PhXRIsKnwnmBzHSuqEH54LP3dQiUZbtGS3/C4wYO1HESZpNBhCTRD73ZOM3xuP
U/tL+HMoWASElXzkecBXf8xGWuCu44weVXMABUt2+xGeqKtczj9FKXXmqLej3dKZ
Pcsbso1l3Bq3m1Y0EkH60pRzXGj9RtHYlo72KzLzJPiT0wutv8ofyMhPAYaLq9N1
sKFNmrC4GIwqkqM01zEfBpIb2aT35ZGCWwGEcj3SyHyHdzKPJzZGuQX4ljIJ/0JV
UgQSHFvCcGZqCsdvC5Nm4WmKEi0G6oviTunUgjYKf6EBplmu8kZETUaPlfbwokJG
/lHSF/4WrDQ3uZAxjtr1GhXFF01W0byowFgtN7uUSYH2V/NaUGc9ZziRMJWUIFSN
sk0GxNPS5S1EXktrTHetOwO+WHrEfStsCR+REpLHeR3cZ8yp1WEEAQeB/tCI7zkO
09X+5XkCJZtx/NMTrrzg4YN67EWlXCJGeVFvECsyr/zRgputlQte1+/13bo4CI8I
RNXKXzmEJSrK/teVs/NkKsYrgFe9bApAQ7g7QZRcWPQfXGZ3OckPBMhfAT+sYoKL
sBHxq2WhsK8W4l5JxkAcXM/+qUtQUiz8k0yjTipYQJDrpMMqpLmftYlJEu1xFQ1E
GQ+f7VVIaE/4bxHP0jERI9CwEM0zR0Zp0X2Sk2CY7eLwofFHud3COl/RhUC3KNUK
3tC0ZCwUb5wywe6wrUamyuBfdqsPtyrcM28kzj2Pgafp5i8kBB1CQ/lXEEOA+vhf
0rEZ7CY4rRlwvDyP+jydiqegZdEny9mq1ied82S8N/T7NPVzHK0M0efJlqmCO/4D
lafiQ3yCEgcEULx05abU/GSO20/KFV/54utcTACYxWgp6z1GY3azy2yT1IjmWmw4
pXGuxz7LNVZZ5o5fuBb2qbQ+aMk+iSpXBbFCPGZS3PqF1aauW75Z83wUPprvW+f8
8J1Gr/Azb5FD4o6heeUwEY04c5/Bbv0T6V3yeF89lH3eesv/2glS+XUNeQchkcKp
Mt9hk/AJUrnEANf4L+LLgJWMI7Y5gIn8ZMVKCEcP36Id99hfgJf2x7F2Q4c8NCNM
FM1G0GbxiBcr/WpsXGMWYQkW14s2y55Il/rEU1LYq4B7Liz1Tde5mynijo5kEFSB
o4mW4S/V4FBZipevOiX7bFB7Dl+MdyCSePhY2RiAccBNL+aSEUn4JBNhLa7Ynuum
mZtXMXERmMpMzjqLBH7VahnRbEEF1qdniW01ldmbys9RmRjzMVCE8PrHugrmsByO
buwRTwHLOs/RAoZUufYKg5HPoCP0FdoUH2MJSHc/OgrkgsnvQeLUdGreqqPinw7D
jfML/RcFA7cMYbT1g7ZUUBC9ll5oQB4I9K4IEIcbJHV51wwDeL6hjCMKKBuSP9rh
FOwcaw44z5wNOXYxlsKZ+TWonymYD8m0quD7lFnv9zurWjDtxLLn0cTagMa2aCIU
t0v4+XKD54UsHpttPS8mZOYmn18hJ0TZeXb+0ci5pQ0SvSk5rRECIMxxchbeGgE4
UeAgDSeu6bmt1Dglftu0ZK/T5all0lnayLeje+kLLcIsGm8UC/IP0JowiDQfH3MO
ztC4kNalpFervckkrZcirwLskVNOFKnnROfnesd2axr2IT88+Gz9S4WL5hX9pIpV
qtdmB0Qwx1arsJHBwyFpocFnRfwQh2tjyhp6tAbokNHt4dIuURTTGu/VwgkXUgKj
YlO0VRAVEps9EjQGir+aKozh4DC0P3uuA9Q4VSwlAqd6+VgZUlhy9thToK2P5Mq1
XcDxK+PV67B3/ZGIPd+5/nHjJjTEa/GC0JojmFFDBEOGMenvuGw2yst70izeDCQJ
ZVh+Zs5NoNvAKUYiKUcl3kQKQQqjCN64glafRnRRY2JxV/43hYm5PnjP1LVQ9uFf
fgDAp1KtYA3IR+VAZiGJPmpD269RV2OQdaMxcQN0yjtwJgtTKUxp9VM4K/6mSpV0
yprZYqvrv73HhC0qhGtdhkPQ64FaPIDmAPydL72Cp4MImxtyVtkjItJ7xdjf2CaH
kmhPm1ZJMnB78SF+Ysi+3RO506J+YAbR6jQitahfqvwy/uoRJViOi98Zh8xTSNSH
7gWoM6kY6KVrbgYqWl+VDdSbass4eFW1dvIfOdue8a7pkr74DJXgN7b3alU0pr7S
I26G6RDj6kB9Mtqaod52eVCwldU/BwUIIJEWfLLRpN28/eXG6mBQ0sfd4ZZfmwFr
iyHnHHbg1PQlAUId3FnM1sOYOC7BSBCsKOhqpRzuhuSPJqiw3L0HzSK03pWHZ8et
plDjl5ksh4PY+ToMlNLk9F5/r3xTvXCAGIxj/VzBRKPYuo/gLdI269a2KhTlfhrC
p8iUGqw+ftPNzjJ9FbIEs2jP3PdEOSCxR6mrSIOVcsBGh4NKqyLYYmZHUcGNaB0w
ZUfGJN4ic21fLr3H7goEwNFuLFL5FZrczAFGC8eeNHtdc/kZjlhn4oLeu6LyfQlJ
5VXFO+Ig6SdldPqBw8ZfJcA+Oc1WHosL/4zVWsPXaNCJmOIazXrlzODMKY425ezO
j82Y4PXuyMSEFOqXUI9RxBzv52U0Vgl7L+EnLI9xhcMjKvxfEq/rR3N2c+2K6g8a
aVoBy2kXpdL6n377kAgC8CCGR989R8PkS1geBmjeNKDNKhtrEpODG0RLapZ0C2mP
6oXSehVkcg/XQaniBK7wyIcwkG5AVsAXtxOhyauzxChXUxP6lB2lT7yADdtp23KF
pNc4gHX/gjId3wQsM66NOAWXI0KB1D2EyWIUGBCzJsZA7QxOjT5r4dxCuVW6N2nA
qJ3AjNjOMZ/4t8f3JX+KNFDDRfCtLyy1stPTF31g5CnbDpS8pkn0DJJAndtKVJSS
XBz0K0keW04LzW/7FP043DWGWT1g58gpdFJrk5GKRDGjlkUPn2tST4cOU3jC20p/
7HmVKerXMPfrPY/FX2kb2kT+1uig/DrxcI4kgesflCBlbMmDBgIm/qXUjxsHKyem
yNDv3MlboWV9JvDUUlWtS5egxrlfhG+AWk0k4btANwPW4hqV8dS5ey+GIBvoxNO5
mvR6YXoPr3aMnGxvbT2Ayiev5F0V0gb7OdorRhXFpiPLfZjxZvPuF/5vzcTyW15v
/kOci8rdw7eTozK1fG+EtsNKoa44VYmBQ48yNNSnl3M1nfSFduvvFVWyCGcp3O3b
QvSsFgGtVgwjeR/wA5GoYyil8v4yNWVwyukSG45mn4JAhh4hwoyRfWd7dRi0UDg7
O5P4CG0EFn8SgWLqFLqViPqlOi5TQwUuAdKhXAvCDFuAweZWQkg8LsH+Yko860IL
RY2VPPp7ctX7ouBmLH50oY52MKoXraDkgmztM1Jqeqk514S1vZtQ5DoCFdj4gz9i
mgS5qnKF2j+9FswHWpyH5M2el7EmCL89WMo3JQhmyC+Blbuw0Zv9Qf/UGo7enBtS
TIE1XR8Vkga8l1nBKaqp8ADYx+UkWpITbveNc4ldmUbGpYgzekIARz1ZqtsqTAZb
A40pRD+kOVSSv6Epg7DXk+nPb+y/qobu09c4WAb365uZJ7zicNWLMEWoLZ04E/XB
FB+3RjnyauzZsXanVEus8mpjbayzWGcw+Vkjj7tzSHDCET0yc2IcASTCu0Gk0KZe
FeAOqNGtHstKxrjGVO0uuclj9cwvelCWlpTJWaok3h4rk1ujXmTFY/bO6zrlIy66
43ugWHIJTcYpY8j5l+vyxqsyj+ucC9rLWk8orbfuKnvtDUq8b7i52vwL9yt2mkh5
XHN1+0tYa7T5QLTfxgfGjKjKHOBccl/uILY+TGbSUFyQGAs46yOLAe3wMoiRmmqa
UN+91Q+PhwyBYgD6FejJL65QarPc9gopzh8bi9e9BiVD9vve6rO86dqQXW+3lbEa
w+QCZhneN5KyosFD9ENJ7x10ufF1pTwaCDAgbwii7D2LtBXZP/5Wq7Rx04MgRYMC
w6mu8WIInH76Lt///UhTTEuNibVqbBkMbwrNFN3JXkC0OkatzkW9XJd+t4q0BpDa
kBNGzHoZ0wzGj49VdK0a8fM1PwwNYpaMmC/uBS+FuOt7zFIReygjwMQ9MbB82hco
75c49RS9UCCvw9sa+M9ILJWN7KDChsoGbMcZwiaaBUBDFgjf1JdJULjcUIBr/T/4
kODwnz9UF4k1P6Cne3svK9F4pOMToipe0JBuptV/s6kYjXCpRr0obx/hn0z0in3H
yk812iPrPj5bBhCfVNLZ5XDzotAGp2/s9BzJ/CCrIKpVJbCoeoUCF2b9XeV2eV45
LTqqzReQBR/ZUwo4VaFeS6SsAP46UT49JkOEAhP45M6VOAjK2ieC/WuT0gqcmEW9
6pcuKOlF9iB3/eJykJRa8Kuxnx93dGKJ+y2/E5cIXGxoyUfYAiNu5TJpVSEf3CCG
Kes8J3DpBQnNGOljmj9nlctqH+w7vAWx3KPk20imVegdWIYL7wdF7URq4zNbrn9s
wLGw9Ufd6FoX3P3pRcysplGObio4iYh7mHewwRKB1R7PErDwrktrea9Jn/3uvQUP
Pr3LadvC59R2SCJ8hJMEnmi9BYD0UqPgjOzBCdlVYj3VelTgQcaJva1Cv+eo6r4H
20G+N6BxW0xGniRy8QdsXXPCMRLV4kBRzGrXwc4w9wBjh4OhZMoZaMynx55c8eAi
ltyC1eDdpiSey5KrGkU3ZkZaQ3X5kYOFWueKEh04bv/Q08p068D+WQ8oqjiSW2Ur
kF/84Cc0NuVX2/vfUZzImmwSoLRMtAw6vsm9mMm0+G4bM98hB0ng9UnzRoE2RGDs
nF72ZFWkojb8zDHaOfKOQGOEzYO/RlLOvcNlufutB00oQ0sj8+sHsiGc8I2rJmN1
jgIYTHThpXpZMifsDMy/nA+98a6BgAObwm28Y2vKvcgPXUqzcHNzeK9pZq3fcBUv
5MW++uv8wjYJpzxfuFRDftSSNEom3p1DW/j6s9cCjfPta7ybvaeBcpmPvnflTj5A
5V2FpJy8ygYa/yflk3JMIt3VDoaVe+7unD64IhPGCcuOyY88BIu/WPE13vEtFKrB
5Be4/m6+ScE/7nV1at7xsbQpL3y49ULHpvjvdSz3UZ7ayxGCq6WfL2kvzuHrLEQ4
mwkdozLIt76VMPO1n5Jqjn3O9w8g9xdN64yGnBmSFd8rHd0j3illiGWiruHFbC9j
LvlHN3kwz+LRjlvJr1aLWQmjsxAgyLrUKVZRe/dMOWeHJjWz5c2jMTxfuZZBgoT5
Ho+5pPGSgf7jsb5zZrA9rpH7bYFgJDCkKzrys21EUW86Tvxp21ZIXf95QrelaHDT
ntr2D3NniJtqZeyK1Q4Vdq4jp9DW2P/sM2UJnNN7ns1pRGiD2hUl1BVrrnstQGVw
GZyQMYGuHdDmKBewdOPj/MignVJMQorHcBvu3sLMLR3mlMoR8kN5QaKsT6mp37JA
ait5x3jvZzBLJCflkRGKQO+FuuQsRIvEEm3EEbucJW1D8um8RfwRP6ps60PV+VRR
Auui1s938O8li9ffuGuzlStG43cA1429rnl0f3O0RK0hCNkPr3RPTgj/GNZlbXCl
0hssPEjFYy9ebqDxoabzKQFr65Dt0aSM2Y5rml2JNzmwgeZL3/NrW/fRKCFXrAQ5
Ke1eSGBu7BDV/En/nLsIIA2cMgzKQmFgIC3xh/9y0KeIcJpiFiuuG7NkS9dzA97J
VnGsrnJ3G59fP7g+YhSCTPwjkutd9pmTUmIpk0d1SYGMxFFXFyhZXLqNu/o8HvcO
vWlNzjxQ/PMGXKdw0yHT1vTujHwf5TGRdfqz3eKFZZg+kYCp0BwW1HgarE4C+4cg
ZxiBXkQdQ8fW5+Hhzfk+vg8jrCQhKOvoTfd26UZI5Wvz0fFsVI79uRS2WVFc01oW
ggZ3CZLDtCKQuSa68LGV5d7BWDi65ZOTcbkDAczQhjQZ/j7YkMRTChWeTGxFZo5M
hYVcuBFQZLvQcJansc6mtutTFckLk1ujmfPEYTCflZPxQiTJAOI7XhqNYRoiYa6O
oZYu8oTIJgYL+vu43nNGaNR3oQ1Qu42tuKEcqv6AXjox7EkQnAmy7/YMZ8JCUf47
9bGN2hZqZ0qFQcGhZ1p630hhHkRKh/Vprg1tXG0rKD1Lgb/w7YLnYMHFQkEdUg5V
eoisDv3Uulc/1308zECanBtss648wjH/oxUJCdx+ERms3Qb7ly8YUs3qPWSEA0J9
AKiqcU0j+MWSOqUBYH1Fn4qFo5kgAc1VYA1XcvNqWDQiGwzzi+omRqeUb61TVB1h
ZyojCZIbtTLtKcUgTeBbf1+nCOlrgNXor5/nxP0FefYzMVnh5l7PguQ7QSFRScp1
9ehA1y9jhv+XprWlboE4JvN8k2lbJBY9jq6heqnbMJDsuAGWSbuUiJieGnfvfmPM
njfEbQO437Y4/dslmUOcZ+yoX1JrO/oGI9eisQgZtfKQaOblIceQtffsNRb/XdDm
CziAGQS2kG7RPoyrrXyYkVOg85yOcT03yEtyK/UAVqKF/uV0sCvRhgZm/fmx9gWl
eu1JtQGyZRvmqoaytUMPIcpgGKMSNxVmMSmt4FN1ta86HpVDcboy8eJfL3pp1ulE
TaiqQoOHVxQ1Q18TREEyE9NS8ImETgPGWwaV5fdmoC5qMGO6avkvRWKn614vBrp7
5SOFb30jQnttbSLkRxShCEiJBLGVGkgz+JBBJXRaEQWDng6xXVHSAQgaNy3BHi+S
onApzkYpFKxS6KTKGVe/oOmunTdHkVBDE7yyrvqn4Ugjk9pCu0Y8FPlHEMILepiq
DV5XiOLtIdtP9zog5fE/ecnfd2p38RRZoSk2d+7Nw1QsJj1Xwx/fZsiV3esKof7B
yp6fTO3NG1UwvsfnsT2DFgfb7ntm97PxkCi4G/SMxB0KduJIQrZmCv7S21DzLXMs
wJy9myTxTVkc1aoYGg3WiPfHh1uV/NhdMEA3PmC5La6KqGP/Tc7kjCTXMvemCMJn
Bk7eIaSiux49EJUbwMNZCZCVDQoGyuaIZr4ZCQuzvRhEgvFGKJUX2L2mEhYUVE67
7Qmq7E9H6H9kCih9kOO9KQszrCaoIRnYk4LWCFdUoJJoo26f0mlfpoISj1LUSEwS
9K+ZkNKtcHJybVZAIIOhHCnMnmLm4yNewCYXw44PyeiIuTTCiQKBIO0F24t/Xs1L
yHcC//mtgIGe3lqjaap45adgGeCE2O0vb8Z81RJq6M5vskKXfiehWYgbtQuNFrpM
uNNVRLDZsmDVLdRrcaGOOyYn517nlF0zzBxfoK3tWMxsDstl9R6LFuw8SkC8UUg9
bAJUZ68Wt9+eWhnhgCK3jVYuSZse3HlX/g0JB8Ua87QZPcpLgQtk5t2k0YMwwL5l
TAmXiYvJ8O4zzjv0KIvQ10+OFSEi042Qxv31oGjJJRRvu6rYnxWeGFza8cHSZocL
jSFsW9TJQZbzpgRwzjKo9AQZ3d3wh9rGQde2ImGMv6/MWUMaO0s6ADes9xbuH8Eb
vLFY5UE8lCdvi0AeGK440kpKPZS2uLiNG9xr9+Yr9L8aqc0qgFWDA2xSQsk6CGRs
+xce0aQRG52S8cmmJD2fUqH0bbC/051RdG++36phj9kGmk6akAXHLSsLRbLI4k8i
UXhm+zxsx/bWHQ7Shfko01x00thK8o+fN8lOl8DdNLnDd7kST6uZv3hQid6UtYp4
r8mSLkJo83Lb6c7OfrRX4qkIgJhvFVjB+BIkv2VHySwOU3nFgL89IZmC8GPpsJsZ
aZ4W1IDPu1kd74bt29hh4yypsMl+10xaJosreKNiCtMLSLFvcuNY8Pdty/ZKpT0e
Em51j1qf5AF0tR0mJyiVO4DVkl8NncGTg+Qta98sy2uHxqIV0vZzkZChySYxU9oo
6+b7wKN+1RFkTSQE26IUYjL/UJ93WEH82qURnFEFFHTn8IeWqYMAan5tCHwpAKn0
uqcBQGp5YYzHFjx2vHH6HAc5q8aSrp5sTEC6Y1Bm0/tFRXq6YWmjwspbDBQQiQw0
hMP8G/poFYEFI24dBvTyYuWvwaOzJ1J5obxilnNz6V7L+swbi6qXUrsvAvY4AHMS
QFcrrem7KieaCjKPd1obYUxsrf66fx6CS4HwkcJl5NNlPY1J2J7TYVwWJhjP/6TV
0T0LjUoTuzqoHLNEsm6EyKFkNJggxqkKOVlJ5PNvsQGFDkSKaPBoWjqB+qZE0F1z
RJoJra8Jb7E+hF8KzJIUt7YJ4FVFV2ERILnzDvoJaQ0GXB1SkrncAITMe5l7sq4x
bQ4IXvIqjXtGNwfQA+Uv3jbgjA8QvHmJFbcySRIalgNijSPkYWQQZhlopTYTUtWE
2+hXCuUKlgjMitO0mxHtH28IIx+7oz2cP8dYjUwUIN/4Q4FVfH7afn9nsJRgBTzC
j9i3ojQBosuDMZ7CN1efdaagQhaecpG00IeiS4bdPNbMD2sJkkOf4Rfkn8xBTqjl
u45W/2MWbVk3xHctubgsWMuR/Tg3o/YJHlmvRE4FxrfQ7CH8VB8O7LROBs+sZOdt
JnePgmFVcjExEbARgLblEn0uX1EE34bbLNMPa5vq4gQG+sF+fM2w0a5JyRpb4zHj
kEuQ1o3UECWwiC2Eq9QstDucg+RTNdg0WtNc49Gxpj1egcVJslDtT/cBztGwRf8T
x1x0/67j0FkWkQEaaB0EjzYQbSqC1uoeoRZCc9x9Or75CzrJECLURJx7FL8fpD4C
ldZ7FvK2isnnp6E+vATiVf8Di8x368wZ3bORxhCs5ToRj8QeqSRQCHZyqu5OLavJ
aYnoAtKYFC9arcZB4/L9NrScGeLIlVIBMVgioFUBHsxO2COwSgBEBMmk38boZI04
1VqJoo2re3hgU6/IWY99VzGbdvbuam/OLoHPRIlTxKnkUUdaG5lU6NtBNlW7ljSB
DOuCnQiwJvsUuW0tdUJOToxLspJJw4cxVtmhedCrazRb95KRHPTS3cLG/3cQ7E8x
trMGHRaQY1xx/ItKWR22VcBa5Q+qOKgATUxFEuj7ofWZYy9eXhJF7S+/CWHoJwbD
YDDLEBeTI/HMeN2PM/JFQlqRg9EdKNtuGf4NHm/RzlufPEODdE43Z5MkYfV/SJP+
qQ6jZ+pHla1KVj5OoDmDIX1Ogcj4hMXLASlnLsP6T2apBtaJarS1rP3L3y6nJrsS
xDNASuBDW6hsyB74rw21tqz03rjrQf+97MqjPBVe71mVKIppuBaIn/BBiPVBm/VC
giOCTaG3j6tuxmIz/BNQNvQwpV22l0jdGYs3U42jDJaAsB9xCB85w5xqcfaJdyH9
YDN2raVwi93QJCsUQfEc8w7DC40vXMisFJlkaUyyovQ+1H+l2CjmYAKJdmPahFNt
+kqHMFUsUDrApCGInIDUvPPJSIA3h/M9L9UE38tuPWvWxVfmWLuVZIEESje7zouQ
AGKkiA2dTiKBhRBJ2uP8cKx9sbP0C38lnbfFx7+P7a9Xd5FDoRCfNXTafzGPrTzx
h0ffVT7r+kdhRnT0Z4KOtZEuhvA1xMW7LhsiVzzAbjvMU2vjpr+YmsgfCCxZN1E0
fCxTKgXdiEPga6BTzJevh3rfwLiEwy1zTRpASrm0JCRWWzfGhoN0vxFtFtDZuUOT
YO5AakLvv4t0lMZd7GhvunjBHyMUAYF2JPQFKXFiKMfoeNHJu3BUBEnpRXosD9A3
mzdkCXMDCKTC47T5pzcFq9ZyzS3f6cuBR0ON3nb7C05LDUTxvAGwpJsiT3jYkOm6
XqdvayR/1Sx9erSMjuRh9MFDqeV8tXXPu+wI2maUNWTSp16YVS0rvvxM/t99TRGd
vpPuTmuZqmrAfktpIM38L53zv+elT2cQlyK0vl2+mOUb/2fDzbSC2S/E0UdCMhmD
kDw6Z8NgAI5MVmLhRvkdsC06ZoLqN0jdckhc9xXHZdwK8fHRLKxHO6vuBbLBVqQs
hUXUtVEHpZt+Pl6SNpmMZ5S1w2HbClgAhYbwldMBSPoztF4Bei52JkxYFnk4jaop
D1t5jAGpWd7S/Wek96A5f3oK6BXp1WOooIjzYZELErK/Osu1lFpjNsmDgPpSHqyn
0676XVRlKRkZT5qcJrzD+JfTJwl+iXyyLrL2oJZa7jTfSZEUoF4fs8DNpsQ8X0qR
0Id3RA5EozQrjCF8tOWI1mapUJ+Z7crEctFuPMjosK65X3PCBaBHimkuKHklwupt
Vh0voXLHkGGI2iXjt8pD8SWhG445TO/hRncdoSNxFlID+oBZrw8EmtVavwPacoI5
JvV9JoIVdn4r93wppJQ0mAMsMIfHsdBs8eDgNOykYdUxhfQau1HQLO85VouoxSiP
8ulmTbHD70/8BxLtMHZn7UE45y+YIMhQUC5+7YZifn9rn6fYwsmsMASP7NIhjvLX
idzTF2AXf73zwj4L82YhYSKU41tiU5lRhAGEocAGt8+mYdIQqrcBAvirGgGlOTRb
pT0HdbEAPgUxhgdxXmCXO1NXflq41NT+B5e+cnFtuB3VNC4hiXQb33xezEJcL4qC
go05kIpQ3SEOEdqUGqyX1DbKgMPCqma9CeVawd3Cp/Mtra3Snm3jxP0G9YhNEp6B
LMhKQl+dNMZLsU5M8bYA278LQRbMEB7VQG0SU+g3dlpI2k6o/w9y30eun0cbIXKP
lk5S953KNaNgHKae5XMqcVbQSdaEhfAPUQkBYHFU1NWshGMV5vGFLmohGz9j8Zgf
BVu0Gk/vxXjR7zBfrlE3W44rUxb+bJgMXCFJRxETIcot0WOYQemekCskuVX7Zp7F
RIbkKxydqRXTVV8YA1nSK0BUweEQfmROA+cTGj0P2Fc90IIXQzqsb16FvABaKsKn
h4Xra8AnzBWXgWbOEU3FXVfXWDoyyOFQOiXgEi/DrXFHEYUfPWjOkIkFiUvoJ04+
OJwD7Q39eoTF/zjSTk2tt/deDD1CYmqCY7Bp+HPXDgmy2gFVClY2SnmkLEBAluqr
ZmcnGgE+VsLRYDXElwXrr/5qlRXRLbG2wHvwSA/i7t1Goo+sASK3vvWE+ciQi97A
LTPJNJ4uGV/D+h0aQVadFJ220rOsSSewpXdM2wL4bkp1eBT8I3ZnXXQLeoNyEr+r
HS9PvpKXvkOT3F4klFhOldRCGo7LE5FvUqIfKfZ4pSq+2cKNYgUBja3Bk/CFySyz
estZ3kYTgWdEGHo5HAxw1IBlHIB0sv4M5qIKfFhyxrAtLWvBVabfGdXxtQDFgEej
hTQlW1rxeENEqW/pkzb8LABN1WTWCFT+tUNuTdpSV6lY6Xq0SmdoALAit/+Gw9/G
Uyl1iXTCrUm4Jyz6TdtVoD6qsC3kMSGae05RQQjdrFqDUfcHRMjCfmvglYFnWcEA
oZ/e8CnJtHgW1DHncO5sKIIYxfhkjlYsX7PrOEf2rrsVW63y7DFSXzv1Wa3syG+2
Yn8Kvk33++Jw0+gcgc4jiakpEtQeIwfppmML48X78p2JuYjR4WvfiCZlPBjhnM7b
hu7iMp+7YlNFSSmwDxx2Mj744F4frwa+g2lcOoBtdNzDMpYtpd5hWsyAHfdzDw9o
gR2tW1mkRa6lBUBxU+R3DskKt9LmsD7/RHzhdsMgKj3f9CkDaR5gUcRkJijlB3KO
XgSAOhb0PIwN9vBVaaogVNgFByqSOSya+Eu8FtcmL6IQEoA1ApI43XFbVoAY3/He
VYqOnsow4FHJZ6uEYrkkV1FgrWyrnIcTuiWUZIOW7zkIeZdY6SzUAo5v6bjHUt3a
3pPA2NsHvr9zKEscLVgdgMO/Y8FUNFTEPdgL0gopguqgDkTAmu/wCFxUi2Mkl5XA
PN60Qh8LAI9N82fXP0Ld8j9ohgT6oXnE9t6PTTLWH6Pc2vECjJUC13Jb3y+0eloI
UBqsP6hT56r/eM66B5dCnrGZ5yRhAvq/qC41LcYr4SPtTHJXaKdc/jxCmcxOX/1N
jPa5+icxva25WOL+on/yHNFd4w6Vx3bIe4iReKv0oID4oHXDlv8pBHwQ6yLiAxhu
XXmOr5dv7d9IlqR7BNQerjIyPbfaExQeaY8XZ9mmh+BxVKd9cntmvtQ9k4JPases
yr+S2rIDjapD1tGWpV/f6HwZLnUDZkwew6wZKIjWV8eCQQ7eme5PB8jDLxD76h0i
Y4vCrSaRHJsmqpw9zEmgsK1t99ouQObS6NtFg17acOaR8en1hCiIIKTlV/wL222e
YlGDq10dl2MKcq1oy7Z1X6LBMk4LWfoXXT9tHl6tpiUL6KKOeTDfyPZE5MZ4Q+g3
m7fixMjlk/WYheokaq6jH1zE73bl4TsUOSHO0GJ/UU2c7GON0HQLfiRh/bfs61/A
IF5npTUpt4LhucuVfa6wiAEjTPaG3e+rh4S3WpYbI6WWCx38/6Hsas7UqyhYRmAy
mrJNVmpg3gAIRoNCKvIL71YSWuIEz2HXGK5sQJF0cIXGKo+2LMUT5uoBhdSPQcoT
HRaM6jAdOLMYitmfLiBzNVqrVES70ASO+043CoGXnF7fyTyJz/1p6nuy0Zx6AKqK
SedHQWeMFsJ6xS4/IrqAXWHkopXkSkYbCJMlArGUz8AbWvKLr2XkI+dysh6am7Z5
msIL1jQSibVscohhS6v4eka5/j46OYpsoMA7z2F0Buabx7Yo11BJm35mCA8htTO0
zUfCtURYuOmMxLex4bYkH8lPonmmcA0cCtwgwrXf8KK6Nfx7J7l16LST4OAPZDn+
5wBuc7FP4ARqwTdxFSXEi5gKWdVnQEvMR4yuiTVhkJiFHME+iJXXgAWVKtoQ4cRQ
pjQTy8/DHSFKMJ4AG8Ikc8x0aUyR4V27oqQdu1NL7GK3is3ZQE5c3JPg4kSb4jyG
Mkvfh1c1iaaOYRTB3BWho64TApMWUyuueJWdDbadYEfHyXyeGULlLODKDLIr56ya
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ge8S3o9zLKrtOFJg4PI4Fq/94Kgaj6Fpp5aGOr4ZN9kVIJlRm8VLJkps5ohjFyv1
IaJY5cm45pJsFjCh1OZf8CI6drKBeXzaRVbDTp74dz3/95wsvrDH0xtsDjHjudZb
GPDpLIW7Jphxpyy5WzRnLzEU36BMdNH40efKtVbxAlvptxZcdIJApHATt4GJk61w
47eWiFPE6hZiLJ8K16gO1TlRGi7x1+bGUlPPFPG1ILcJGT3ArdSGrNudB47sNiB3
++0FMbvNPIr3U4aBBQCrf4jhr40W/ZgDVULeb4Z3yJC6N5n23p1opc6Uf7ewTR83
K2qM/Kq/DvNT/iJh83GIvg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 20400 )
`pragma protect data_block
SeSAYOxIRy+Lzwl+Wghpx2b4P6ceH2X+QjH3Xs5dJsDzUj3djix/ChiUP6YoOBKv
LqKZv7jMNbBij78n6QQEAIjW6FFcRvrz711gmhezbguMqG5c/Saha1DZCjrBY4i2
x3zDojlJr9jmWFHwnvalFf85//ACBTDCSSjduOESCUT3kVmMbZmrT2zI7EhsTuq3
ZAfhKr9MupRTxLh6jpGPewEgbFPHGQK9GKy2c84OzRBhsR6MzEgeW5Ic/NX9+05A
4d5XsmNpTuhM3NkS0kQ4L1K5F2FTSLV3NDHAF3m9CmTJ97QGPEPunOulTNsElkZP
C18iyxu+AHHP4Rpb0lckSS+NKnxmYmqIm9yu41W6nPg88+3lcXGLx6h0qSGmAHL5
S0q7FUfPr2qXVp5Fcy9h93WeCBAz5gMwufmf5Zr/qb5sK+j3Ubh9SBlFNgQrxMIp
vmAJRbNQJGnMQf7iOt5F+kHORrvqarwahvO6AE+gq9CjIMQgKzMvoHKkqW0XL9OP
RK2qxhxfQBp5KDFRGliaEwaAp4ziIuRmT3DdGKbndnTzz3OXEYL3NWouuIRTiSKE
ng1G6v/NDcG4K2zmzxekE5q598KBTWQik1Ax+SDwPWlbc9kceiBVeh8zTUjTaNrP
MGY/ZDlneLry6YbOJaIGANBffPKjfteX9u0yyeyL4QV79rWYs4dvuhCYQwtN6GBQ
PmzxfKioV/ZbZRJ+0zYTGy8QdesDj2XPfrmve84azeoa/aSTJL+XWSvXyKZK/vLg
24bOW6jxoqh6/iGsNomu87x1JFrUaxV2C9zI0kZp/EpB/DlQDiuLSWhftLayzh1Y
iSEuNf1x+yYgtVix4OGWIfa7iWis2XrDsh7xd+DK8C2rTQbvN9S2gmy1hh/AfCMA
KViSQN1+pGNPB73OS293ybXYJDS5cR3JGyf1XNUO9o8m84SMyjXUGQlGQnzaK/6q
uSZ7h8CebbSrY6NBp9deVW7fqRGLGeQjt/LbAMu4bVJGEUMsnjDNU9JE1QhSU/ZY
5LrJo0OzBSpYc+Z9NetlT+yAvBiQsBudFcN/vsQ3kn2nh+gvlIc+Y8w+NA9sEe/h
/vnFHCm+5I/snYSsstRhVz089yCjOBcmTlPWYW1b6QZdit1IjTNNz9h6B0SH+I5c
jU/nohVc8EAdkWbQOWo31FLc7RyvB9ZoVVU1U9gl1HcsvKxfhbsfWkpy9IYJGZgQ
ZpsXFNMZKNXtO94ahwS6GZSNrZi5I7BziVZ01N61f7LGbWu4A2L2GNxllA4FJIgc
xPN7I/b0GU/uvEC8vgVZpY1RA7+amRbEH3vwR9spwCPbL55NEdfQwQZjf8jwmlcv
xQgNJFUkibMOk7hNfEGH67gZLVTr8ng34GxUF3Gp43XQhKunVUCB/5WIXoP5sOyF
ZAadQAFDR002amNt6em0/rtOjXudXAyvBQ3WU6O46bWAWszNnGZxIYdRM5BoKpqN
CbPL0U1f6kQ4SPNmeKCZfixNAX+wJc48RO/GxS4NsvRlAhAQbtdCW566ztL+bojr
tL4RbNDzSX+mmzEc1GpNXpbLCaJ7AH1dTCw/cBPHbfUmYqP1efdKrQdD/ApiR8dh
QhTlEXwuGoXMTpL21otNlU/W6HGJ5lC5MIo24wIXB/YnyqsHo1WUgoxzQuU1HGmZ
r8AbsB0M4vLYb00k0mEOe+iWyg6czv6LYW5mD/Wwc5y9eqR1txrpGgnUlTH6Njry
V2HiEDTQkcNLyNe1yFxByqIi2jcKeWXvEtiPVzYUeblDePWZCKBRXPFZDqaGbmyX
eD/Hs4nze9QrqTmdTp5NRDGKAqi8is22MrYjEbVFDHwGqajR1xUQR/zoXCZ+9yo/
Q/kC/wyESxJ+5zf4cwCzCgfFbhY70QjU7eMgLPWfTr5itIOc92EMwhHojbxaMAea
KRnzv3cv1KjexSDOg4/haWIn46t/5YXk3oJMfIzRCcyAdcH8DqWpT33FotOZnfLf
+JsZxtXFvn/73UaLUN+lCHJ1WNoYHn1rSAedVnu/NbJ6pG1PDTTpqrVeHf3vzU7/
vqCVKoE8BinQvIga7n9eS6jFd7jVreLrFL8VqSLq7K1jtQo3m8iNMTkBLfR2E1oH
Uiyn2iRzHkYvIEqP8iM95zXjtHfDr9VKYZEJQKPOauu3J+XkBCMzLzPqyWQw8qbj
VxFu+4whvfxOxcKt7oIQotlzvQsYuXCGysb36o5sAg/hwStXP8AW7FI5b2dWclUn
VtaoipfKD3uKNcPcK5f/Gu+WHaN+xrGK94InELxswu2rj16ucYp8lpgwo4T9ISKt
0G7pe6VhZ2eprTdS9tuTgG55/tfJYFbScP6fNUF0SwcYbQFagzHOw8Dh2WrfwTAi
QfRijueZwxi34YpMF9kBfuLcy9K0XU69Sa6QKC6ZxV1+vLkCMExZM/WzZNY1K+54
aWuaTu4uJgKXae4kHYc07+a2n0z2Gro+ZwRm8voQA6nKW1boZL6eYolVi9vB9LFv
DkTVn1U7fIiuEwRWKnBjy/oG8a1o1XlOb9C2KbpD/Rc5Rp68hiZuuBX2juVaFRMH
83COO8uMa5WglZAhtsojB9pOYzzxGV1UwhKNn3K5VV1nKVCX3q0ZeD38h/anqhw+
JtagkYnJJe52Ae5mnd+KdcUSrL+YgYCDbt3MeUuNlN9CulvNylWnx87aXeATu8FB
dfZAvIFdIF3aiY5ttXRFlR7rgMv3UdAWxDQdQnNzyQnYsK5NkuhMl3/E8bECbkOD
HcAH2ESafgkoj1OYbaqoq9owIftTJSNkRzOHJV++N4c9pOSGCiZ0sEuRMKOC2TCO
lEB8Sc6irvPOhi/18u+MWt1Bnnimge3walpNP/z8jJxzvoGIODct/AeAK/l+R7v8
qofnbTjRtQxWNjXq8cf6ZtMEgl9jMJGxJV2oJKo4yGlRDQViXGC7Z9IgCYd9Aojk
zzvAKiwFBJ2l6uyIK/wKLuqcfO816iYHQXBIlJX/PwvkNE/T0o5ndwbfa5d5net8
RYoGWANe6RBpA52EjUdAUXhypUwbDZSA3O4Af8i9ourYu+1DF3ZuX8/cIJh+VsO0
IL/xJw/qjeD1z+EqHfyIf/sUU7iMj8xMK73hDs5JUWR9vXp5SrUwUlz+D6d/F55F
yZmZURvDDioQAd9bYmluZXTSGl7tevqnnVde4hGrVRv50bAxzPEMohKt06J8zOx9
eDl/HtW+QT5TrWGn0CbHF4Cej1tXaGxsytCpQloKNu1jSoxZTjysZgq+LEb88pLg
odfzTvepDN59WtCT+93jMLZzvzbn7YpZbE6/gRoIJ4eRtqikLuCo7gkXyt6ahpD0
r9gG9D9+jv9+0ChA+ZuOe10U05YsHYTALFZipo9f3QFo4Gh10M0wa7WwLsgZISxL
ccl4KA07Aqke5I3hlCsklDmcoDD7nw0A38DbnplXrBvT8wntMrRf9aa3dAhiS0L/
24H+jhFTDhY8KN9HJ/AUDlJojZ6gG7IJnuDy2jockbyhSXOneZ8TiJdUzIYPHeXh
RFm4BmUiW1oMA0fGsuvxUg7L9tZzHidZaQcmUuTpJqon80NXIWdAmm8EP60AV1C/
apacUhOpQgcNh6jNXrg5YmRpDlFXpngmDg+sC0zc87AL9bkrwvIpfHxD/gL6r6kW
Rz0hdEc9m2D5ympeP7q5nMWbxPuWAJqOpe2XD5r9w/xwfOwW6sUKshBpxFkfALbl
uxiLYmBWs/J8EdZDE7fzT7/zxron9I872/BlWbckZaq9ZZ5ndtJb34alc2o1ZKvA
i0fdxH4RjrVw4G4UrpbXgPkfwIGpZnCC3FjmwsQ4wsk6OeLW2YBT8yEF0lCnx/QD
m99nOh67ZqSOkhkYXiOBJQRpEWcDg16T71jjiOSrmSyUmiauXlUollkPoE0K33n/
U/tE9N9Mb7da4lSSZV2hYxAPPiIy941qXkZT1nCd+kuDYCpk+xEo48dPetg80BqT
yVKQ/INKGt3h02rlCE7zoexngZfUCW3eWVb91o8X5aWzyLU2GpWFUAmQ+kCbCIJW
MVyE2HV9FLdLTwcU8n5W+nYXuOxPsoeX34sMkfM280nDXX4d0iCuPcO8FQDdwa58
+Zc9Yd+DjyQhV4oEgoAFLmzpBVznCOqbF8eDACTFTPEhUxYt0gy5VkUTtgc7YsKM
MO0eyIE00t02rc1W47FqtwMfzaRn939MudEcqCVYs3BnHkyeE7N9vq7ewj0Hjklg
YkS1tFu83UoozSkKIw7bd/PBTjU5isarhdrCKLjSiGpVijs8BBiTy4hW9hbOPoeJ
YPZvdzv+IRymJpxjmyZnIuMQaCK/+CEFwZJxfpHzys/ivPariJjVCjjLbSGpLMa3
O9Fv/zXUNuQydeJ9UPhZrG2Dc5IWT0DphOmEVIyGkPnXfrqvDbOemlFNR7Y/diae
7e8Sd0MeutGFEEJ9a3J7QT6cpbajWnHGLXI3qsx+MBmI37pg9XxaAuAm8/3s3onC
dQAtPTflOxF0hvK/6S7zhfbI6D8IjalTzO2LpEdlNIkrggD9UVUSb/uCjc+URZmz
PrpXzxv3mYBiQ/NJDoGQ+c9Xt6CjPfJiTxe1G7LxpCBtrF484K7NhIpwsSL6J2Wm
Lx3FqSG8he3jhZkyTiXITOcd6mVrEcw+AWVPgic2INOym+yzgbcpTTR7tEQ3rFn/
VjOMnvtphBBg1Kki3pRHDSbQ0QhszPsr9xQXMegT6O//JUQ/E98UFTxI2X/yvKDT
XKUS5YDe30G0YHzaZHgGajW5qdWWJ/EzTM4lpBRYOQ1GxiB6fAIn9vp4iq43Iurg
OZaClsQk3bqy4kSaV2U/S0yntnfefu6cqmuOXXDeaDztIM/s6N9Qa6euWr/obELg
qpCYNCscNS6nKQKmhzNp2v3JWEB6uikZBrO1oqWCeXsgcM7DZ3h755RniuhQA43J
ktxho8My8E8bu9UmEkcU/84ihyDZzL6bWo678wqEuiMOKxKzZkzkogiPUllcIZVD
hmZc/Xcbp3tnrfYB8sZx1yRzbq1zleAWrCAzT7iCejY0aL9jppASvzHxNc1XEhD/
q1hKXvIcSln5BuQhUByGLVOqpVXeVdzTv95ryTf6MrSKQqU09A4+gyyr4bHsiyEd
sc/ua4PTGBLVsvEPZUUvFnox+fH4siscBe4SGM3SQBAkdSKrGWvO52XjjoZ+wghh
NuQUqfzAPb7dvI3sQKhGvf9ww2yYCeCKCISW1lThAubz0nOLUEOZrXLGrAUZ294F
i6wAQzGYnUevbuCyhGGSlqYtRZoSmjkxvbDC9VD24f2fu4WTBizPpVPUGqHcVrA0
YDcbeqOAZx3+ahhRoM3xf1rxQbkLVWS1VxtQSabAhB0JVeFxIXZ1vT8JyuXMVYRT
B/I3Unvk0/HKRLauMBMJNGkDvcY1We42Q318K3sj4M5wrTQdsTKC6ZBXF45QklQH
WPF/hYTXRT3EIS7or/0WioOn90aNjfHLn7YqRmjMT+KvVGTvuON/7n3nfPPLRwY6
q+Tb/Xztz5rjhOvaOvQBrypLZ3MTJ5CCC5LGKUDT37FsrDV8jRmK2FsDpuu8xkMO
IgBMKY+B6dti+vlgLh8lt7lwwyL6W0TwBOMP+eF72XMK0MeEzM4n+dSCM/sj7LFZ
Y3KwexkvBAjspSHP8ReGZkrQlpaBs2lG5a/+iCbyKJIJTPP0sH8R5BU7sX9pM5AL
4sryLL1z2CAsGLjERqjHulfuBuDJYTZCrUz6cS4QNxV6Nf62JRboxLJectPA5WyR
/9ZqQY73WPMD849zWn5rPHmgKTF3s17mbv6NiaVvWECnM1rXpSHQYBHTXc8dTAhq
CoL0mS7HRsJMXTEtyllE0Gpfyx9Cm1nhJiRAxHrut0tzesTcH4cZ9xvA+Turxfjz
igPpi0lpIxukZzT/wLaygyMhvbwAWIk7iHB+kYIywyBuUtYcSOgj+dmRSlBc9YE3
NrCNJUhrDslpG3R8L+gV2DlOpWREbUNx5kzoRr8uPdj+Pim4J7c7ZMVNe+hnpKh+
RtA1ySayL7SqgO/0HvpB1IS2sobJs8hgtAyqbzffPu4zM0ABJak0Q+XAOuonCj9d
d96gJZKUyHhOEn73iZDgDeXffRGrbxW3y0eXGyZ47pz3d/jpUP5JYBW3LEjngv7j
Fa3QM1vZb3F88LlQISfXdhWonnsFWMuRRe7D4MoDMpAGvZ5vGf9zXvCWBSZjs1bw
jupTlEv+cwGFk6iHGiPemRf9b3pA/UuucI0d9Nqid9zxoHJAZoh4QYu5Nw5+urGE
BFHeeiYRBIOHdFxuTsrdcYsQpax0+L3cMOPfRdJJ82Ip/i4FcatDPD6uqeQxECkA
XHsQWh50Sy2MA2erPloGkc0ic7FYM5cFV2+jKo1mnliEG6t1CuNo2AvoSCvNfAht
tjPN89R07AcDt9bupyMi0XyXdc5sZ78nWaro7RrWblEm1PPnFY1hgInM+KbwE1UM
rgLyMRqtA/CJYrXZuFMC74kZEhvnVzeorglkQLVx0XiSok9cXRKXi+d6NIeaJdDu
xNCbqkpGRL33lNmDPidds3VPk7vMlCTG8UrGcCVlxM/XrUewxhOSVWME02fsHAtl
jcNn/gPd27lmjqHrxcwZYcCQxYuDLi8ydGNex/hmLBsSrfklvnU+HzAotZ5fGZsx
YHg8KwRQCRlAXvtlR5xcMSknRjYuPGU6VHgA9jJfj7ClkyhglUwi1OICQGJKlVd8
R7HS75jGErgZDsyllJjhI4vtXzzc/Z0fm6a/jGqlh1e0W7FEpMtqCgh1CO/4hN99
qdAe2SBKluYy6Ca6ne6V8VLuCkE+fWo5XwIO5rulyWSyEONd5AGYZ6BvuGXz5olv
r3+F7u8GjeUco1JgxFfsHHHw4AUfdfjJjv4a1IgzScHtJXxg6Wj/c7oVMLAQe+7P
EWoxn6JXv+xWWVkv2/6IwkLytLo7G56j0PH5VMt7DkxxKVYq8jZqHsykT6WcI9wn
rmEo4feds2bVgZ7o6hwYKwc++J7jSIx4U3h+zhsTCvjR7uas6Z4740TXIUeMMTR4
fNVyXjtSm/6Txhl+FMUwTfSywRX4MvRUsQ1oU9CNSH0W5o1GoVbANVujXKFjTNdB
HMh634M4SYNhZqncWhXXvKdLzDMhiEZuFMGaEsx12KEVePIIT6IQJFZsdxvL87wZ
v3+aoQZgVHeHpRmRqBfB4b/GIQ9OoiCnDq0a9cCwvQaJIy/2+B8LBoCEOZL656u5
PJujMvVR0lGJsz0hROZ6HWzNNTU3+R9PwtxU2BX20TQUhk9SbuwAkt2PUraUjgm7
qpOm/8OhrYkJbCDJHvWAaoBpCz5orNejSMK7k/Q7TJIGwuctmUJvS3MLUoHyJYir
EqUDJuaADpKNhWUtYHKWms2RsqjABE3VEtXmjmFxoDcWvHMJk4s5idpZ/21HnuTn
V0HouSNuFw2WlJ1qBEgt6PZDY7Ln2S/FUPeQXrbJrmxCddAoRY1JmRy1j5qSgVPl
NGRd+yQscZUtVemn+1rZP9+n4FsIWP0DGi4dGiSKL3XdEOHNqi1Yj5ljF49mn9ml
yXQDK54jT7ZVmeCp+sC0VK7YaVS56wKUsonPbzr5mdOJsOAHSp+e5FyzOVQTyNTd
1lPy0VANE+Z5QlAnY70EJogNb1JGGu7BOF8El2z7gVXMLd0T9TdPdJr6N8QdmwRD
3y2dznl29bGk0vBFbFEMemkOphMexj3zQPedqlwpEc6au32lXXsEGTQskqIVCoK9
H+/ocpJQwWa0G6J+jDUJo2JA1nfEm3T55WyjorygcLEi5XiV1v9DSyxavDRFi9My
j8ROpSNnqlRoZe+8Ba61Ow3GX+rZVp+w6yUyJjgAQkc8OHHpCZ6oQZUl7AmB7L9f
ty4cX4XTZzV8WCg1NvtbUGvioxXAKnMNh/mTwB1WnR2MT/LtHh66q2rgkv4sXn3O
QvG1SbvxzjWLuQ3qPiurmgqibjf0B7M4DWL6nRoy69kV5KYVoRjgfkbbJTgQ61tq
5ylgCeSYEsS2+tZJNOD1DDqjYwniSIF8A1Obn2/EsPUCPKaM0XcAMqJc7XiWKMzJ
dpakh+ly1UGeKEDJpEbtByG1UrKjf1VSd8kGAVOiKK8LzFotvnJXDbaidWENLb8T
cv7FZClFQwH7UDloxeAdwXxgo8tLgwEXL5IwpIGbYts8l8UfU745QbzAy+pFt99O
8rElop+moD8tcMjEiz34YPDqO1EN/czrKI/p7GWKsL1VAE45kHrFCRZHYBzGd/e/
LdJse+ngCAyWhv1WTySfmst5CfzJZqhOYPD4zcCRa9L/HRqRLjlOUVJR95+TLSsn
Qe8xqr3i6JVeZZ8zzBVWn1cvp3mt+LMLRtjR+l6XHB8YuO0YbXTWLw+ERjo9+q1T
sMRXNSGZPzHObh/Qo0HvH9BTTCAgVABmXsEeuLsXbgxqVWw+PSZGFo7AQN3POMnv
+aD/oVHEVWGTf2yfMMsVXipvYfou5e4JcELkYb7QmA1N6N9im+MuPLv+rJQOvzCD
sr7pSg6jtAjlHABkAL5XvWhPBiklwCU3ST5lSTf6mXz3ORtA/c5jC9/ID47KcfY6
n7NSDB1UusZqjzn+KhaUW2Utq6b7eemeI5WpEY61rO9dFLnk8kk0uBJaIDlQExur
JdHAke2+NnpH3BjzFNBIfZ0gppnvrBONNukBpBtKkT0hAKk6sY4SW6i/clIABOam
SZfuz+9TVCUm1/VcqW6tRLz30RzMkxJTRBUQoZjXG+i/hxdx13VWgerLU4gdIA7O
U3QwvhffVxNOOhEtxBplCCmIbiqC43hnJ6c2siBOluqiCVJy7TuOhk0m3miCL7zj
ad8mHqIRvUPIiha2CQTNforKTZb7EMWYDd8Xo/ED+w1X8hdlE1C9uhlT95XzI0+g
2qqVLINt4+9TyLWiAEtejMk3GT5iHpz+XPpmHbnHE2aTGfoTlQejNk31VBijiKuS
fpU+4LBrxD5Yb0fvkFaQrhtuaYIoyzCjo/cA+teF6oIQp5MRdZyvzgBdReaYzxEm
9sc/x19vtgdKKcRxNzyrgovErgl8pACRNOV9du8Aocl1wQMM3gzoGRijSpRmlz0v
Rgqi3ujLu4ra5IekOJ+GmRM8VDYGGYJGWXr/Ut2gvdCqOFHrqPS0BZ/4q259ai5W
ER3avGwONHg0WhiU4gDV4WJzpkSnwWgbo4VkWEIL4tgk70c+1gxPWnyR7cuirAxn
/Yrx6FV1ofb7pFSle8WbVmjWC6Y+xSB2Bl3DVDdRgr5WefczJyVyC+Ps+BVnWZCj
J87Or1dTBVH/97/K1ggBBSlUBXWwpeJ1ij5DrQdDE0rMM6cZaOrL/C8D+0Vrw5AR
nrjp00oRFkfM7+JWn20PN+6awWYvze6A4MQ20N5pDJypGuhnVdzPQgG0Af4d00f7
ErMaUDdzntTIdMn8wn0PCz0VYG5VVPTVLsY3vPho/oLgxCRx3Ngo7A35vlfJlXmr
bJAZSDNlxY7NZb7aNrpWEaw79bdZoYdsuTM6A8K4R3CEd0HceLaa9kU8R4ktLdvP
2MLHgFf417HFBdt6eFqWUVUj3pVjmtccVjXWg720Iii13KixZpK68N29E1Reiakl
5+1BovLA5sZ+E9jntDEg8LfyTUiIJp3Jhs+/uWaX0vcTCxsEeeSATLTh0vCDfcJr
c2HbRKdtOQ0TXX0quhIC16r1uhNJtg71vSLPu+LJfRsGpTvtejnEHBsLo1TZxkJg
XSNchw/rJfkb/rPMVn9YZOp+PDJdl9S165JTkT6rEOlVU4kvh/SIXuscDmbf9BmC
5LK6Th51/B1tJDsH5hmWFb5IppmwQir+P9pxmjX5dR6KSIeJGygAJ0Up5LVtchdF
ekpHc08s9WGv3jF/mGlkR2bk85cmt5D43lfDVlMTGBurlMI9RREIGL02fkgdM1+Q
HdqBaKNfkslLlj93zJTzu4PkQdPWYBPWnSAvfElp3CTuJ06ohZeRA82DJgo2uKNR
4swrpKV4WBcaO5c4qRhFKNEJTI4LFCJSUhlk1+u9FukGyy2fSpmYvhPXm03emlIx
mZHHDevAD1h4oq5PnhfKCPHOAglovrG7wIgpi/J9VVoA9Dt3Sz1XlC02jLLEyCqQ
9zTsKwtdrt2wmvUrgLUbfSoTBDw7Br49vixKgYMvP0kYyJuokSdqbrV31LmQLDyp
kGkcASQd2Lg1XKGusOvywKR2Z3jLHj/IDUvDqXGPsQUb1L8kgDkm0h2FU4y+h2ae
Hbmkahd7SSiQPkMvwWTx/TB+JzPPpYO4/amj8fiAuYD02lB598niZbWhtb+p1HTV
+gCa5+awC0qVHxmZo0yMOANGF21/psEQxWYOA1I3FhrD+MdspysCrwwJpHK+T859
kV1qAkNrerJHiHK0aGqUe/DlwU6dGkcO4ugFiBjSvzpR1WBCqxTzUTKty9zk+XyZ
Bl4ddvSLtXBjeetkUAJflp944cPF2K1br52PXShP+3h/rXCoTkNS5E38z0NvX1ru
1x5uSoIdUdcJ8nJWHthw3Y9BAJ2lW7hnmqjBKB1UwuFqmEwV2I52w9HJLqZpFivJ
o9xVryGXFpLROYljrPW0+tl4sjpziU9AW10xzAXaWI0neXsyy0fjyJd0VG/4i0L7
EE0tV9Lbz0A2gUZ+bDlOBRcIejtw9T0sHWp0BZsUU9X9hH47t1pwlEtfWM8re98A
RyBJMpzGejnwJBPS8GHofeJBCaWRFImNgvTtrCC880VLEWStiGcf8d+/SVadsIVb
MZNvi0d1UDzzMTRL0XrX5E+QRFPOnsbzqZ5bXOgWIlGnxxlUpn2srWOkEI1DVUgN
88ay6mI+WdesTogMQHNsjA06jUbJHzXNNrO6Iz07WUsg7zx3wi/5hLaHzpix6Cu8
tpzZPN1kIJtxyrJilh5nSLvLCO/0Bk2CSzSsEKySlfkghEYRYuSJBgPufAzUSwhB
OMplBz3lCDfvA6KLNuffOxCXQN4dXb3qrNfFAYLi7BpS0Jm9p2Zj2Z2peHt1P2yg
4SqkfUro38bD9gEc5MMwPGj5UGd4kGLZ1fWcnCa6wNaeWsmyhi+9z6suKhdbftTJ
LYrbjbYcK9nr556eicVOuoix5wkZ4dyArI+MQxHmK12kTNQ4TvbuMINMG/UbcbmS
Qze5cY0W4dwNBXIv24epOogla7ffajzZh4YMuJFqJLTs/8e+Cw/vOETVo0rljnYd
YXF39atMsblGxY03STDQlkxjb4jJXO0h3N4u2suVpnWFf3mjwGkRHauUPlw+yLLe
3l3ACBcDC3szXzq8LVzbNzDRd0zEv/qfDhM3oTiIiAa20s+frhFEcGapr0E2H/8b
+au4oE5G+8Liq18t04vAF5lYKhTcu5LFBniCO1A5DsyfzcmU7IxzIDkiJ1MoEn8A
Q2+xPQ1PCckw0Hn9AltZio5JnbHy3LQ+PN9nw6BSDMv+xWi+t2GTa5skn8YmKGwu
n2fN7J+g5UrJtumwfMcDr4LiZRjakBedd5jRE+xCNHBMB/FZr+nErEmiXpvuH4Z/
4dg20CtYBWhDXKtJ9/5FFxBIu3Rq+id/R/Dvyn5l8B6QDRIHF7moOMlnx1qOxiQc
b+0OmJRCvF5qe3qqov9CNX4CHcqfHqf+o/z2VBoYDWXSpckDDGa5rC9ZHYXtlvO4
EXEKGMJiHNS0BVx/iitSfspWIXkEpKTiT/eGgzuJPgw+fUWEkv74VxZgMmTNZ+T1
c8hjZvV3SVh/FvY4IuVeeTdgVdZRIk8s5M6Dy77eS9IlxiZgu3eFGu95PGyzTpSR
GfUeTzaH9GYStK03ory9lyWTVrNdroN2OrLY+/wzSPwpwGV8juxkFvbJJ1aeuvFw
/Sd9bazc7LdcflKlDHKMWLgUnRRRcA4ZUiJAlTENvlrZHEsJuGM/o0q4hYMngi/I
p5Xj5Gwlc0KiKsS7gvvn4UkrELRB6B9LCvkjKUhvrE61561wXhu9HVyfyB++9VqG
MH1VM3yy/P4MhyV/JCvbS5dgmeKDrbmPQaML2baHtl8x0PGYGd7E1o1cL76xFjog
E0wHe4LjKUal4RCY/ESaMSU21276xh+zG0thBVb6wjlchZvi2ib+4psM213pYOM7
G5DyPvFaVKsni8ZqPePIJRCNIR4LIcRbV87qIeYCoOVweDvvxzG6kTWuO503XBmO
xWIxOpctJJfr2+lHTDDLHBs4dUjDSbbCtFlHv2Cxs5sGZtD2mgr4hDN/SIQcWABK
Ywe4jtRH9Sr+ai7LFLvHnC3rZp3riDgERgT2wiDRSbW6jV6HrixoV0MUaIAo45LU
H6vyydM9FLTbfzRiKcpQeqlMAiThU1VcopDhMUTvpwK2Hubzrn79oSk4VWufy3Xm
dYUsranp5mnSuqSiB2VUCOpDkyI/iG1Tiq7GLV5LKGOCn81uzj9bf5xR2rAO+rN5
6cvGuoOrOSn+9iA/Fmb3NSj9CJ3yB59oaolqsX10X4v6IAE+rUcCwdM9utpf5TBH
YB8ey4hsZ3y8lgx8TmgwnbVuGRV5+oLwtEO3RBcwIRISPR+2MNzk/Db9KSE4CjUm
cbHcWVwxXvo0jmEWcUML+dY/4X2jsuO5mDGj8btkflYq+1DcI4So57k5vd3+pEeu
r5EJ/guQDeYGFYItgi/XQFnqh3Qs3olpaNGQqETA4anZlq7fY3+zsW4BiHNywB14
9761fYjf2dsdhcWryvijrDeWXmaAOiEsJuaU2cmqYf7HUCHA3baXyQ5nDpbwx7KI
GkeC8DpznHdpUCpoYLP8sB6j08BUIf1vzvJigDPsg98JH7UIQV1r+7LFyKwkYvMr
fSE/goDLDRihKlkdG7gxy++LwnjmQMp8ltuDORUOmhFig2LcklLlbZ5018RmoE/i
L2bvU89ETe4wbpo/51BucdWjOGCtbtzayQY7lKGkVZxYRMs9q5Kno3YWw4lW64s/
Id9RYMU+qLi9EMcHd2mVQwqAV23nYAXItAwqzGGRXscmT+SjQvxR7CMAY1/qN1iy
2jcjdxgkIQ+2WY+bmwvG1h/iyMCQ4G9cPZr6G0NUNmf2tm3bRL70aKbRGawOaIqQ
ExiTaMQZLLqWOG7mqohQe5gWr5tgImly66NNmpC4Kps/r7yAwtWVO32iJDFSd0xV
T6FKX1ayfKmB9D7L8a7d6suCgPKcPyNbUPdwXNtseS+8uS/+qiMa+LRASPYhPPKB
E7DJ659/4HnSiibSSyE9AG74ldUmCgrgVr6MypZvtf8v6SPeHSPq8g352lXbt5CH
pr3/L18YasLSW80jysO+pKA04OQ3US+acyU5gEUmoxhq7nDGE/xxT1wZjv95O/wA
vJvxAv1KVZXN06r1BNY+gKbSNUNi1V4zb4sYiWYVG5bLuVrZEPqo9WaOePQbrYY1
ProfYsOSOnuhotoF/oZE6SvVcNkPS9JyusCr90iMHOnhZ3QgjYUq2AlN6orCj3Zx
8KZ6lQQUT/wMgogIABwjzPCCDvmiWMX7eYW7WdkGAf2vJQZeyCdfpz1NdB4tMY5J
V98YvJqzfiYN8fQm2yTqBEId1UUNU1/IUD5ZMk/7vqk1MEojaaOtXBvapa1vKHmY
pqYv3eNoR7i7daFy85Vfb1vuo8Q8updeOmTQkCG9FycFEkcpeXwwvgaYAMca5WiY
DYszI1OH/4n4w8d8KjzrjhHZF2LREaMbK1Bwm5Y53KlFBleuvsI4Mlj3CxOdytTt
3HvYvCPcGCjejEDMorPeDem6FQ2cuLUdmrSYaaSssuyAK9VMC1/DoYR1LJ7Bu2NH
urCYWDYyGy3o+D/xkE5FW2h0vr83JjQ1ynqKBAzFcSr7PtdW5xXzvAdbnAoZyO3F
9SAll2D7n3ufcPg2rvu4IGsMjE7NSgi4Aue0AYUQOnOcxeTgVCvjNTR7yqhqUhfz
yIQg2cyvSMntB3ZY9kMpcWMBgFJj6aP/VhiDcWjP+yl0v4HEji6PeM9LUblnb5wl
9Tb2WI6fHwy+nR03wZsS498z8EbtyHhH5nJwGzWHV5FdphzXnj2Q9RlRfFQR9tVA
0FdH/VwsImKmGBzgZabEpspBQH4xy103v0Ooo1668RX/zxdqcBwdqFZQEXwqiPhQ
57EZrkJd5CiM0pWGBSAxgHXlUT8rbMewaH/Hb8u33e02LvfjFUKpNKvbjx0fgqHF
WJwVG7PLYp7zje0qZV4q8WCg9W9i/2opAo5tx700h2HJQXEvXD2yL9Ut3HWOaIo0
Ry+w2HcwsKJ4b7nnXJSuuCmHjStUrx1q4cYlRZgPAuHjDmIjzprmvzzpXGAFd5fv
N8/TlBc2zE4sA8uBaPeNIl9vzZwUd9NxLR7HvjA3cQJYp+mbODRLBycBcZ85Uxsd
yUFO6z1V/dCPaqsU4tDWjANYGCSNV4ah2+zf0o2vZtRLZX2ijDeGplNj0xm/mWmN
TioFi6EQwaLAmNTrnWF9ubms7eYAGYiNl7yRAhwvlnczCO66YLIaN1JNyE4LZPtd
6KR4kLFyuew8jSE1ioK6VX5ckpmSgmIlj3bGealaRwqx8MqXmkkozMrZlEV9dOay
F7RH9DaoY6duocl1HngL5XdCe+oczUI6LsiZqnnz/RkwZn0yr1R9JEJkLZxl/OtN
1e6fiy+Lb45w2AlqfP6SmOColD9VfkAUKM/+xh2YRVJZcW7Gi5PGsw84pFM8PguU
jPm1YOHQigzkrtTZtaexAVosTJqgnW8jQECRoR3WWUGi1Ev/RYaLvKMPkWRX8idn
Jpvidim0DomG/OzcBitlV4vR2e3g4m2m9C6oVWVklIce/gFeHos1uQduzTSw9wbP
nR42EAREKkkjnQBZTfhn8GiaQEAmg2aXCc1+4ki7p0jUFQ6MGiJomogfZAqy01CQ
DyjtVbAb9oBs8QAAyOlpKohtZPFJogUHnnUq8NJYfJh5Keg5LjdVfRpKxWWMh3ni
YQ8UwR+yi5P5lAhq8qoGvgs9l9a+M+SFvcyMN+CUR5zxl1c/S08Cfd57jK42DbnO
yWC6NlG5kN82KfAs32NTMma+d0hjyYpBDG8tw4Vr/rKOz72L7U/COFtg37OlFqLL
uBBLsYoe7EiMkamPdNQzqFdmW+vHa7t96e7wqObWy+tAN2IEItqnxmfWYFFE2u7S
aGXk4ItbnftCQKe+6sqkJKxHluLtnBrLesgsqFU9rzwRZ0gJRBnQlZ3kfhnTNjp7
NTuXAn4lYa1dxYaNbk29lPQJI3fw9A94L/gtVtrXcfc+RpxfiiSsNgN8uchdfDd8
b06w3CVuVlS31tUbrj0MTqhKGJfF0pdClm404asxdm9wisMs7M7utnho1Jfz3oZJ
VCgy9DA/pPnEXffkGTr9mQsl7ernBcIQoZumSlaSJLH5J1SDZBD2xt2bsV6AmKE4
oCGvhBmF3I+ttaPf6ZK2qcfEVs7UhNGvxTYII2dIF/rChozR1fQsnV4yjjmhRT1D
viWwk15mxAmyJbamwqfHiKtnNEaS57hKKYEbHu1PryZJsSdjzntgCP/ix+89OuWQ
Q0YPxjxrvKVcWGsUl9rrNIAU02864HdZy5jAOJAYPAc1fnAhbRz52r5pOPrBB4xK
Emw32SqO1pe+SbcpMJjp3C3vG8i+mnUEtPLkMfEb4ApNWlkuvr5u6wVQkEVwIwra
mr5AoJtH6GN0iYd7ajMK5FIoKDJuwn2SSkQXGfLBwq+F4J9u/fyAXVyaBjojgIKK
XvBNLwSpwp4bpikbADqBoyW3b2ZatqITYOkeSzkYhUEcAcQibjWhOiU2zGtctTUX
tmQJRz4IzUy10JoRSc5lQ8PhEH/c7bvx7pOfml2L0uM65WugCRDVU68g9EBNn2KD
7G5sT+p2zE1z7hAcDurkRnYe5Q3X3U2ecxETLi2W9O/gJFrpXifqMpxtRVYjIBLa
NoVfTygB655rZYyhJHaNB+k6OIgnlKY/dgH48Pz0owl/KLaeOAKkq97GsBrMA+IZ
E2wmT7INyL0w26QRU0vAE6I+eRT5M1Y/Ayl/Vku7v3r9EerQL3bK/qRP1pN2BDiQ
2lLojP1rVOMev69IXCGqLrh5LnHmuMCbr7FK0cy8wCCaoIV2rvEpLBlci6/ie9Uv
0AdgJFmJZcFjjcAbqtj+capcomuQc2AZQoLTPHATIR085av/oAtmFx/jug3gO28H
aBdpiu6zDH3gVVa+GLNkJAAAsuy8sy4VpH1H9CcLGS5rX1xTuabgUjRuHrBwo4fR
pPdYidL0koBZja9O3ImfsNxiso3G5K68jyYd64vwpn/ab5NB1UZrq/bBhJHGkWbd
a6csNGjbHn0Sgy7sG5nQ3VEtLTFKf/HqM59+7+DVBeWDB/K6JL5XOXNkeM8/fh8z
d3ABUaYN3s8khwdQagfwtSN2KT0CUiTAAR3XL+yNJ6B5FM2Maw3AeCR39OIh7OXE
osAhct7KXWGiW/EOvvrl+EVAtdo5UOAxl5ABGBFLGWhSgzdkReqNST45KdCMU9V6
N0FBi2CAmQv1khPOhTaGeaOYlWfRm1e+p0RadD5Ys2coczmwMHFtNrqTiMAM+T2M
umqTQzuGhxGv7/JZIhWaL90bwhcxB8C3KhCnyWh90nwSzMkSq8ol+nAbtm4RdbY8
9+1+DsK96HMZEJlF292lrqMr+YsQBOz3FIdC3306rzDd/1PDxXZd8kiFu5Ai7u+o
Ih5iR9/mLHF5QsbRVTPCVyMMmyOO/9UNzWIUqopWbKLr3uzhtKOTzcG/iGTjXGeZ
tmlPFdquvtL0FKuVrHRsIHCewyJ0fyBJMH/sB8TF91yCzcpCdEQxn+FDmqfjkXPZ
HDj1tLZ1JN7kTiCb11nDoPy7Gzl/EJiv6PGrsXhabOeZGW6GBH32QRWZpfPIBBLE
oat7QyS6OUeEyhbL/MXqfbFTCxyDQnCr9IqMqakB2HISj+8QKljNNYciP3NbiXV0
fJYLyZ5X/KwcjaFFMf+t7kGGNNwp3jrT00reNNz0EDKE8+4Uo1plYPzYJUu9MZNE
HDvxTft59H+Vhg3oG8LR37ENxTGEZwTbi69oM7ldc+1JMmwsoXdSG/q7cEm2RcdJ
Bv9ygotW5yc0mF6d97HsbWKB20xqoRar0brYcXnKt6TWFkfcQhNM3oN5GrFlX1yy
iQmisjMJWnOPp3OUV/fZGAU2sluMdwD8VGbGNYaDGHphyeIJGxXUIUm+Ly3ruVjD
i1Th642XYVsRv19BahX4KIyHxN9xFF7jEc2aWA/Ze21MSCWp3VEsf3lhSlRQ/jRz
dqFdMcF3j0HtOY54uF8pHp8Zsx0KNxqchf1argGrao69K33z+0MAXSGu7LjtosGg
EzpRw2aKWYlQ82jZkv8CJYkDEU4TOkWmLr2WK0mJCV4V+gnmcQnHSzyjdcP78COb
ek5YJVa1VGGjJX2rpjsXSYjoy9JZ9C/Q93gZSN8jZ6MGDEIskuE5VyxLhIn4lycL
gC6j9jm28RvZmL24Qy4+fsx8L3gQhhzypYGI8PEPib/6JS0DYjCKnaZqU7sfa6fU
tn1HBDWKZYUcZQtmOyhy5g0I8QQ99CaJrn7EOPO7dkHR83suMYEuxUsOjnvZxL7B
VgyICdHwC2sjiYgexFM3h0Nq7JyH5nfAplYKuZM6FIV/RYrSJpRE//82cQPw1ytx
ADSobROrNads4yFUgHoiW7oKlVogwtbVa/jIMQYPXMjcVKWcEk1J/LylZktsSnBw
G/f2Hbam5EPn+Tt1g1rL+Yb228YUYKBoFSKDU5wqftOTJLXTnevDpupTbNNbnvol
hZiBCLwaJ515kU43IVsPYqyvMV3IT9itVmMZsUpXN3JiR9L2dQHLnB90arBiAVNe
VY6/zLdjURBG2+Jm0G1CZX2eZXg/8kapxbq0jUhEhU1kA3qXepGolfgukI9xmU2p
7+q/d5wH+KK/JQZ9JqqFC1gaYVrX2/0vG6kSpbIuLPhbMVOjICiexx8PwrJ6JsKk
mBY7bfCVOaaXhBrEjScE79722Rg10AzTF3T/1DMQjLED8KKW1KYoLYjBl12qLftI
EPcdsaMO82UCjk1Idj+qTxM5wwXoxs2tjoqggQT7rSioEYGegul5eBXnSV/l+FYz
yAv8VD5pzVmP2LmhtQ0bhEj72ipoYpI61lnLoea8911wSIwHJvMm/ioyfdL//hBM
t26ZOz7YPWZCeoAcB18BnklMNpYTmv//2Pykzvbw1Dqbn72cePtLsPNN2XOQh65R
8jasINqWMFpqhYsF4nWl+XjncQpJpvygOoS2xyFNjyMDkDEnNrjqKxScdorPa9VX
GSfRLKOjHNfQw5xXOJg32Cv5s8ZfVlEPN/NtumIDgt9B/eSP9WCCcskAYrxlrkuI
nEmP7RjU1Fe77TRsCXjktXIEmyw+mW+iCj6T2JtEYeMlB0RLma6bHi/3cpw/CFxo
s69R4X8T/AUp/lZAxqRkSPbNKgwDZwcBwhG4FuBqftfvuwXhaQpdbaJPSSLV+c6d
w/tijUrVCspsdNezp0VkViJHAuAKj6sZBI4V68XpA6wFHUb252JKU+9+C7zb4p8x
502ZScvxR/wB9X/AvLFFfVYZIkuRAANW7JfIqiKPUgJvFtq2v7I7GiCrzeEarxuj
LM/J0drTBf5T2u7Yh2qe8/vwEs4BlPGZXTXW4CBPVMLBJ/vYo9aJuGhlQb00JKue
fKFNlCZJ23p69JnTVlNEdNKYeGiYpdEGqI2CUn54KM1FY9ChaOfUmsHZisgOasGa
fpG0gYllweK1eGAjhOyRZSKN9mz007XWrI99WCeig49t05IxSZLhoQFdUYzrJ3qC
XSafEKa51WddCQy8kBhwi5Gj7YAnP9OY4oqFCCugVoDXCWMS7jmdTUNpvbQU4iWN
wInoz00SzhGcM6Npzr0cjmp6UcO+4/TJnA0bAzfvy91jhJE+QpVTuHebAI2TH71v
RpQgho2HJtQIgTKXy+vF4xfOiX6v8Se0pEYeBWOnBHMGgYsj0OmAw4shYPHaN4Pz
9HQI9kxZr/33NPRkUMAyKlfFQd3syn3+lMnTK9nS6Am4njaxtvSS0lgOSd3jSCvJ
14c2+t/PyABeBJec19RqsbxlOBAvxP1+ZQ1f8ILG9vuhpSdNPpiCD4FBru7Nmft6
6wlfBaJ+Uq+RspE1mcprlPb2xZJhK97t+SIxKNSQ6N7Kg7PsOZlqEtJtTyKjNvxC
hbqqivdY2p3EQpDKYEbSq2hR1m5MZxwupFlaMjrVFuEtmBKRfVahHHvQ4CFPm+o+
m7fevBXDlQnpSr70dA8N5GWn4yvWJw7Mq7QCQdPprLOxo+de7/4V/IbsUTyUEEVt
jm5tZOU3rZBR9PO9EKynATdPlXjn+JOFT8aKOV55O1KfDeLg8pTeQ50mXTIOXy9J
Aj7QPYU44aFxN5rNWUXKC3GRSgBIO3ujYXQrTxTAvnR9yN28r4+LxgWyV5Ng+3yN
efQMEallNf519JOPZubjs7gXK2m5EsZkttzMeb2ZtU8FfLtbxMvlZSE+R0BgEkSU
3D9jp+4pkO/R4BM6p1TByHAhRw6Z3/0nRERlWO9b/wMN/XPvqAxUAqcQf7aFD3JJ
xONEWUwIJDpFb6T3ZdF4qPGuJU42QMhGAQuYEHWZXYye/WSgWMnOk9zkQ76dfDUK
Yge8fHAeUkGP2f6hbcq0Oq+HM4kLfBWgNzAfVL4pVMItbM6EZs+yGNXKBSKQ4VTq
9V1PVVXuEJkBdIcqKQN5SjCUZ3ijZPdATl1F31B2tKZBwuTD5/qmPD40YDO+R161
OaHbXfALVKRcP2PYfbWcqkzP1onEyZmobtE8GveOT1bsuU7hwx4WYxH5dEeaBbbR
hXDqLeR4wlb2g+4ebpXUx/eqoV3uays2lcxsSxNuc4BOl6vBIjyG3J1zsYb4qF7j
N1SAM5eogPPbWPOpYrKWXfej5/LRNNui79ia4rtEU2RLm8Nh0uCnaKuKu4XMoxC9
Luv51KdxsGijdzR/2HHazCQEWKJ2b64ZlkleM7i1tKuJ1npgyS6KucJ+vO0U/mJ9
ijA7oKjf7m5GrulGaVivw9ZlleDtmhwKPxbGRbD+Pu3y5hQ9QLJDNNRejJ6kzAVd
VBAk5LQUh7s7Zgk6U2jFOK4qXRiJga8Wdu3CcjRALWjJI8GpIObpegi+jqbUhZPO
JC1GKn2B1jz4o5OpeZIKn0SnCUTZOqqB68YJ4E9aXzuu/7cPPOiOWGq5fS99ApK+
eZQuKrFhA63XKT6879nNOEHNV/fGo9rBnWSy1wJQtKL+igJE/Guon6voIT0fz0Lg
awKUrHiAZ96N5QCow0nHq8RUKHWGdagPaJbcAi+McwQnTEHsqEktiCdQvWbZvMqK
N8mXfh03Ldv6SW3Ea19J+BgtpuNjNSEQUGkaJ6a2PMQNWpQ5LcEm8xmn60tpiNDl
bXj1DTXtdNr1xzhgWcQEEhm9K/uayBKLVL23/LSPIl26zxFL96maaR9HFNB39z3m
buhlWSRd90Eek9eSABd9ITPv9O8fbdn4/m85SzC5pPMOkVkUX4c6Vg83ASL4yohe
FJhp6wd4M0nod1gv560Se/+VBhNb0w7Sk5Bv7ISkkmJBxO1V9BOH+AvDVj7mvo7t
dAr06YZoN1f/6+s5+Rz+/9v/paL751OEEZ8WfMqTRs5NLub49c4Q8+bUSx2/5Q74
kx0QBw0b4BeCxK5KTtnaNEa/5y41OTPQQmsFCy4ri3wVLaJtiegJts77nhn/d8f3
UOLAND+nfLgEhcKV2mCxpdc2Um7njQdHeWl4GnOGCirTW31oDjamf8x1J1PDRqcV
MEtOqLU8DdsnUWCn7LIDMakxmqXy8dStK/PdoWxSkTFUayzxftdeFL3BCSkf8aWb
TRZFkG527aGiw6MeWwhrYFD8t4iiogpjnA/r2fxf0Xv3trA7j71BmzLfaE3gTsmF
eYzDYFST/iRqSrqcM4nkGuJ2CcNGShgNkRMTKw3GJ+8l8cITBa9eQLPIafQMPyCR
dk1DdxTQqHpcwdFpl5pojt7YNmWCS7w7G88hV/cdNYNE0f0TMflkV8G5wLEJD1Bn
SezyPy0TNHaAxsCGbUB+e8ZwQhygEbByk6L8nt2v47co3h9Tzy7T/Mwxb0xY1pvD
f7tJOM04g3XhkHoEH8jLRnvIervAFttrC9dyjV/pDs5IvNiS+qywNd87XunWcijt
UFX19KwLla7RtHLfPD1CMClAk9SlGuTAE0ZhlfSq7UId/oWITd4f/MyFSnc4U5rm
jeTuaqCil+WvDUlBnhj3aoetPxzRMZ6SHcz7mfWJtX3v0PJZ3V1PEH9Xkg4RJCjt
rSbxxnDGweQ8swfuYpTpbauky4GF8JPq7iQM24rExVndWtaJcvq3ZMf5XWxF6iZV
VZCXyFJ6vhbSaNEnVLJbf7sET+s09cRXOzczstdPLtkcRszkMjFtGaA4+S+LzPWp
71pXx6N/doFiBIN4sA6W6RdAMzRdYJOiMFXHg74xC7l39hdlkQEoEHqtd0HdDXI4
VV+3IZGDXNWn+ve/ndSf9+yQe/EcG8D2zuMIshAMgzPMV00+kJzk0UYljPxo+rVD
w0EfigE0egu7JilbF4ve3q/cfKMcXyy8DR3O8LfWpIHPF6VCdy3O13OBbMu5LScU
OH0AaSfZwfHP4beOXtKvw/gQKa+k2h6tw42XKpau6ZcuuGGKSDGAD7AsWXxL5X9x
KkKSdjZ6pgdORBsTdX3TlyiTuJkv6+vm0T3jpejoTdlHwmsOPL5jl60S7DtNwZS8
RCXo9oKPPA483We+OIgDCn/AHPPuBdt8M9CQTyf9vbQn7U3nZ2M1JjOVltyINO6J
uZFPi7xFDXZpLMSEK8qArXWn6YjzER3qSERBIHccHHvxlQ8Kr7Xl0ihwiux3v+l+
6qZk7qhGJweDTRF1jdIb0UYjSnKt3fZ1OPaZp3MBKfBGiu6kInLg9gaEpGugyakl
QtRHkPiNFrdWpB9Ly8P7BKjMLxC7WiZRdrd3/zxNyuLbSNs7MdH8MEioGkOlCD+F
y2/5bNu3j3dkvmMBiAHTDIdLQVB/6XfkdtcdsFnQh4WDGUKylN/w+DCyFBAYCiNO
yoZ/+ci883+7JnQU/TGEJDuTUR4YHS0NiWafZN3f8H0GmDsEWoh1lJo3uw4LubdS
Fz9X70M3Y65hMkxK9meEOq91ovvjcjZpjqr5D7XskOV68fXmHhaGQMIBbEfCQKdu
ebWLfsOvB+v2VRAOW6gcGDgpx2gKkIdCfUC6/nQv0rC3vbC1WLDqDBAL7SxE5F4q
hy4NiaDMCNfuiwyGJLnDD5vpzIdgwbWa5nEuI7qW+F/+lXLTm1ePFAO+EttfheCS
uMcxAnYwz6fgT/d27FNFZJ1a9qqZ6QPNhxRfrEw6Uo8nxfc2uapDaAofNUYOAiXH
nGHplIsKinsoiyBZCPB6SYGehNuKVVCCq54qincP0eJjyTge8EdiWBHv39yEgcs7
czNhPHJJ3wZHuEunxHAD8TQeB+l8kSlCO0x3jJ5YXv7c7tivxV1th3n/j8mVOomO
AuG6QGY7xahNi8wrF37rESs49/P/YbWMhuTbsXl9h/f6OZprknsrItu1H5bgNmB/
lFx2uRphcJk5PT6Ox1UMu4aZpEOHxPE/jAQ7dcm43h1ZayJmQc1EE7lbvzr1eSDJ
7Dc0TwPWrMhmJDsHXym9QNyh+ajQ8GTtsYOEFHBgSq0bk4+qo0y+RqKDIjaYvqyl
NVHc7THElKa1MjFcwCUFlLGIGAvClr0Yc+u5K5TppglNMvtmPGI0gBuijwfIDo9f
XT/5+EFFvngPNmt1uWmhupAH19H7h8M5+8gnqBXB6+ymu6cd0Mlo2sL0kqKCT0qM
15wPxqP9EWNW2Wy+0nAvQt1pU0PwjTsdsX1spXm/DvpEGXaDLAzBfTBiD5EPtCmX
5AzEL28PdPhCtUc1v2gEngGOyLRShV5+GGvPbNDpzY3jZtA/kRkN7CuBs8X+ZKxe
t3BURPlMvCtUDslMOCuxq/IOatb1KVvhb50WstGEreBRJ2qw16A3pfdo37FApqf6
zIPaAYntNB1XuoVFLTTgyz+2vycuFnutCpIso4GPalU/0CFJEuGNSVrB9IJj7EGU
2RuQQ3mEOwWh5VsGZo5xjSIUb7xKvSFQ9tBJAmpAAVKZr/U2XojmCRH4Lg0sUoEz
t30yEkeSYMCEPRXMKBEkM6eRLGCpp5wvXLBtIdsLrjDwhbQj9AubncKcZubgHckd
6YQ8f15UoKeF6/PMv1X5emDHpbJKpH+B7iP7NzdkzAEyL98rpb1AxbuyWpOkqAHA
1ZRxQJPG1MHt2kEEsfniS2SUK9ItM3SDIiCIweZK2bjCZHJpKA7fB7ZUjM/9PM93
C62SYPV1xIAAKYBr5j+effFiHHLGzAeLucTgSaECoG5HeNoqFdOggtkNRcFfo9rA
X4zQWfu9eIbpj0vyBte6pwUgoBZpT+tII1PpZY+TJP5LvCO7SqTp42oLmdIgcTGu
sCcnoCG5YjkAJyKhKdnpJzoez8kt6H5L36w0NovDLWuQw6T2WFKSwvP6KGqCwmHU
X0fUE1v0pHO+qZbxyfAlYaAUt2FlAKgDZtPJ2eMGHs+Hlp04i3QSpe4qNXmaCu36
7lfS6nyo6Sx9j7+cTAiTZYOsxfIUkS9PNAI8kj6oiBse7887crXXtgRr56OOKvuJ
En0AtJmJqDr6YiZny4xL64m3Bb5akyvZr0YSo676pM08GOdwGrcOwRkjv+uy/7/w
VDdshrR8vtyqNzvq9B1kvHoT4Ze2E+Ux4sGTnfQ0lJoqHupP/qzBzrJMyfCu0AyO
pI879ITVaPllxzx4/JHXznE17/8NKKDjslkpcH9VmgFVAU3agWFWei8C7iuYVtiX
9SdlrFdkVh9iC4N+V4OcTdYLKIj3lwk0JJ0qJOefMwM5svpjOqHp+NpXtVgGdCKI
1WV3nz5cNcMzcL/2o5h4UIMx8AFPQDo6uwHDmVwOUQdXwfoOOKKbfqyK6BCDte1U
7Bq6NuJJRdARZJPBj11EhMamMiHuDvm+JNdAyQGXimGMhEZo9CsbVgh/gU7PxwbC
Q1qPT3uDhbc7QaFP28sPPeuZhpObalYej7k/GMQgX0KxJZ4wSU4VP9jpdhU1TQnR
fhFKP2pA8CRxYdUqzpgzj5+iDpZl3C5jNvafmbjicTmovdnGfZzJ9N5ovrmOrAiL
WGMZPLK5dXWQorO7Q3kjKHRsPreHvsyOKHekyAmFmmVRj+mMD1ENFMqaYSC0fo2r
r6i05zZct4ZrOBrkMnodJEEcPXFhEvO+VsNm+30fMeb7mtHNRrPWjivot//lm2uv
Ppp9UP+MdP1NnvK071jNHz31MFouOUiSq7HCQ4MKOJN0bVzsFFhfob4da47RrACw
X+mWH9Wq5EtdhrvKDcVEh7xRYWJZQ1ddSnQD/Jc7Bbyr5Jf9Jogb4ZEZomx8aR6+
IYAvQYS0INaOGWdo3akeay0Zsx2jSj+aEaBNzjfTRSPiPNlEe+qrKzMIbY261VWM
mXcosywLh1dY8nQ1YlGjTjkXjCK8XDckNO+QGZLEcuciNjtbRdbXiuzYrmcqAWGa
lFSNFp8CMNB3bHLoC27AZi20m5peCKoqV4zq1vkT7+EhBjAIMleG6ifSKh79LFDk
76xZlxQueS1GL9njlj/V7XDM2VImfmhjX6fceXkQ9JC17hAT07k0oB9Bs11yMrJ1
Wcm9uivuCakkHUw+Nc2T/uUfz26Lm8596mfl7fBYYH33aLOCS0bOwFf7xnGmj6/D
2GhKkwIbcSxFQXrik51qKyAWaXLhHQf6oMuPYUqE2QtZ+j/iNh1Ldsc8aT57CXt3
q4s5KKd+Bvj2giZ6QmSjobF9pLWcOAltrclW2WmZWyvmQjwfCGXYXDWqQE93paz/
pdJhK5zFqR9t7kNbJ1iCQgnrw44k9IgH1vl2XKFm/eqIKKhVEbJe0RxpdY3rJZUy
LNNlfwiuureppmO+AJD3/g6cqTSPaUd3OFc9nlo99uCUclc2WOTniLRgp4qT0jEw
PpAwZPLddwaG96CDDyzvfAB7/7Ch44nptWMeiIJZG+JmjH6edJmOV/I+nszK0mey
pXNt1twXWZzXLFuAo1gA2rIXXia2LO8fN7SgjV6CrAPd5+PO/K14bETiHu4muTV/
G/fG3AgAePqcY9meg/MvMlSV1SrNoPSP2Q3SnwQKfxi8RH1aPdtT/vVdb48MVLRN
PwDlkPGfnKLXwS4jULpauOicPfVxKhJeHVBa6e8h1S5PhSwtJfKtxNlVHjy14hbG
2nvI+E6TBFnReLKByIUU5vTcYDy+ktblpND6c5SRTqbLjhMTZx3734UpEnFtU6hg
uuHgbGz+TfAwSIVJuRxRn/jwRQB++lZ9OXYEuqSBThjWk+OfCwCRhDWA8IgVB/AM
0MTLzmhauDFvqLlUifZyS4Mbf6KtCJ8HCMbYMKL00YFspsC887fJ9aOyiYIEKwEL
E3hvAt1EgmXvCaFCAXFumDOgh2jb1V/FS1E0PW6nHTQSc1A0o0BOklrNsnv70Q1p
TrrEfulG8qWhptXZKVGeJ/JPMCd7sX0f4TTw1DRVJytrJlgvmde37vGiGYh8zr05
qE2szpl6z9jG7nb+sO8Ug3TP7VNp9cJ5Tc1ZD3iIzjg74LrFYoPHG6/wbNmaSLZx
8caUnBKUChn1FwWFJJ5dzFHEzFcOdlSLJByV6mKL8EMhMkNzkUThAnWJkKIvWyTb
I30DQsJIx2YNPUOmgLHxHMzFo+LJDOu+je8vtVT6cc8cjeob3qZJRsYpg345j+79
NktWfi32Zd6+g02DHhL8j3p7btTq4ckcg8j7Q2Mw6swLwW6+op5/mMskC7liUEZh
8Jg2iujIk0x/ONMZ/pYYKNpXnWI3Bn3VpTTu+nNHaslKTm73wYLTbRpPa9usmGQY
GSvYTYwLIrn4Ef8/GehES9WOy2kmazZzy+I5t1GG2NMYtWWCESgA6o5Ox95z2+J4
rirVDxQ4w3fAmjK4C4lbbDg5TSNxcrWqnUttsIV57sQBD9C1IPKHUzcUQDqTb7YC
A1d7reGx80/EXJdxe6kfgH4X9JgkM3tLya/wZGotAtDX9BlSA/8+/4cHXpPEVz+Z
R7zlXNhy4T2fE3cUDmb8v96zJFAKIuWDeie2Geah+YyK2OtuMSMPCjhshdyn0mW6
1TGnMACk1LFAJLdDiINVxFogyRFSLz+9XBTaahBOfYBCS1E6nAkkM/zz8Aq0+j8/
afDxp4Wzz53yGWzpQKdwjgD5hEQQ3d2u7z/tZfSXZhQs5Z6cn2C895Pk35zqP4XY
qNAmcMQ4C3E7teX2BqDpHb6maQlUigP9JNdGG1UE6IOyFYsSSjVQ9NzroAyuWbRk
b8TEa4KjpVJGS3uKXUtTwFkDLZ63tL7NG68ClHIFwx0kDYlFq+3VQuXYbeu/nuD3
XWQ4vxKLAX5LwuBLRI0PiR2tYElBte7d6cCkn/ErxChT61l2HAl291id7avLMYXU
p+JCfPsgXQooDnEdjBkVlgzUqnq3lQ8aX1eJhPOjC1AGg2VCB5Z3FkMtHkd6d3fE
XWD5D8QhkHu4+x1u9qg3v5/K62DK11MJDEdNW+hKK5dayzZqPXUXGt70EMm/Dag9
DkFWY8gINrIz9eW4vuCQrZ2Tv6jA1giB5//Q8m2sy+X+z1jmZHSaT7KScpyPv8Ve
E1lPsjJtxSJPDwSl3JxeYsYEZ1MtwzB0YQ7A6JV4sVVMEiqLPvtd3zcz6EVLQrnx
025vjXYSAE2J4ZnzCfbFGuvvPGNBOF5M+h9dEVcu/weSF+RL9a7iH66Olfqts9Pm
bTFMkblLJUaRbG1SCTagE0/H86ewANmEKtVFZSU86A8MnnHkmJ40QhQC4iDmPywX
NEnudArFsz1YRBy2cs0tj/3Qm7IvcrjvWU5SKnqUBxbLRc0aOpV6D/s1Bls6WtqN
29vC4qysjV+jtap65ZnHZlsZHh/i98HcJtpc82cl94LKTeXsrmgITbnjiitV5u69
ce7GuWYf6RNGThOnhaOb66kOvic6AKqoDohd5KAmpqapd+7zpUTxNMWyRfDJog5T
orAirE89KBnU4cKPX1DYL2uPtjSRTdNNU4XiO5ENuJYVn3z8P466jS0bVer0BUaC
2rNnzVYLj2P72araUbZiVirYpwcBVi0A+h2A47AMPvZZbCQ49AlZ274nLoOmbaNt
B6ukK1stt9wXv0fuz6ENCuEBO6HJoJRhYqhVM83JoB7Qhr3oGbs3Qi0M2a55ZcJn
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RPnaGZQ2HOBA+Yi0bstOF6wQhR9qdb9d5ispve3fvrUPbVqwiBpBuuzkiwP7zKZ9
zbK46PsqXKr0aCQegFUAN8zZv43c3s2htN61P2e/sbPBokHdKde5jGiZoywsPmn7
QO9ote8RhjoMwKQBivYXyIT8mQiCGMjeg/D7ewrqe0F/Gl5V91IpilFHOdYcZq2D
SxQiUSVOp2AIiJ1H0UlMwDUBwLH846on/JA9T46GU0kUiphQpVyLbbhhwxz6Zkbr
36K+tu8POLGCtj8KXRgQmtCMFNRyO42m5YhfQkLe8djco3Jle2leJ6y+QZH+xxgU
3Epgg2W8IgoyTZEI9Zxzag==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 784 )
`pragma protect data_block
XKoCRSy8xhOiUpvM+qmXH6gd3GZN4OpUGDOruTptXra5NG6v+uQDMGFKz5Naixfz
40GL9DIhYQyZ8MIgOk0KeALgMMLOOCXFBlhhdiqZlwTgk/qitfGwrrMYSZIlBptw
1D/F+4ORidzqD6EP1frwwKqjfNDVALmviQoBCTTlKV9xqC7BorU9izfDLROrs6uB
USm192kGwlloUHbvuXpd9if7K+F8X6v1zJZ72wi/r3abdqldku6b7ftIffm2Hm8V
bDoWC3w3kZcHdl66nivxlGDQyBtothz0pZfMR/iWH6Wx/I35hfxVEW4BfoIO+AtG
7Veb94xlGj30+tdILpFKku4+qXJH5TKMHVAYCW0yxj8yp7prIXfwk5NoS3I0da80
1EZ5YtCShizuMRNkpznYBHfzxuanaTEXPRgrQtYUZnUWK9Tt8gWodr6PQhREvZkX
wWPyY31En7fX7O3/HhEsSS3n/+9yBxRKD2gk3iPNGFDxASoMnOwON+1t1fC4n7AQ
l57ZZSjkqEFCHs7X2gQfVzq3Cl1SzGWpuG9/JIUlWKO40pd0XWeH2xWfyVv/kn/+
rOMbE9T+gmCOiLHgREl97vZMuuuB7MEaPUAaegHrZOg0EZcIbLQznzUwvjqTtPZe
RDvzeyFwKDRFRkKM0uJEeLTzGT4aGyJd+C3wrLKEZPu6h1QsqUZpMiDZd+74xlUJ
ysblMvfk3AgrSX9EL9pCwGDtJWLxOwd74y072m2Xla+G9MwfxU9+9SUlvKxo+jRr
0+PhT0TVvT3W25e1YOPIqyoNaMlsFq5JiyLmKnpwCq3bWrY1MQRhDwlY3Dc7i4LN
/7kUW78E5hQ3cuZyYM2xrZRU3kd4qP2wj96XEb44iGoWCzkfbROIyGUqOr4lz6JY
aIH7iOFCMXqTFbozkgkpo2OaCJWZmaoPVFDYCSmrfsBrZySfmZHoLv/qrMrCtAFN
wzAY1/6u513lszN7V1EJVfwtq2wg5I9tT/yk4fFKJVYJk4eY+75FTYCBxcIL7wM8
0Wt1PW24DL77MnqamBV27A==
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
O0JYBNuR+aR9Me5KzkCN2K9PxAIr1CJqtzXrA3CmHDjN3PhyUOLT+ZchtUMZLZzA
6h8PPoc+TtZemz6XWE/TfsN9HLXcAEezJqaqxFo+mJnd843ZZxqd5IVz+oiPb5Fc
dH1wodU4SmzA8fqJRqyJEqJg6bE+82YVMGGMBNz6/bC6k1GKJbGZxBdThcYC15O1
MWbbLBXMMH/ob1RkA4t1DMopiz/iOL2oBtvXVuocWivYcnbv2Rpzis3zwYcqh2Ui
1/Lh9/khLj57PxcMKXISJ4mlrw8IPK7Beu4u6gU81cSDBm1wPdLaqdR4KeVIoUjd
tKrmfhUQqlWWet3kQp0Fnw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7536 )
`pragma protect data_block
BA5ooFcYbott5dD6gadqUiCrwf3/04aTUhHnRvrNNEKIwZQbnm8T2a6YAxq8rfw8
wOAYneldYHL1qmkShszQJNc4DfjL5c+XfWPfkf36BLE2b8ZU9O6YGYIC+CRsBXDx
4Oga7P5ZgPZKWBMKGmaxLc1AzxmeFWp4LNgkG6FaDvq63V60CTH9Z1BnZQH92D+j
yXdNbBlu/CVPwAcgNrqbVREyIUkCwu7OUL4vof6IFXp7iuDCCyzK6ujESQF7vEaq
7u+Wh38p31lutQSREcvw3SjzFQhVswomxzOMzwFx6ej2UiyCOLyyXbf6qAnaY0NQ
H5pyez/cbSF1FGOT0wFO0oABcH3I1m8oUtisI9ZVAuAAzrSfQs2iA7in4zdtE/Zq
QH+2/13kptusIKifH3dNJJ+0WIHefSaDXMvppBFURjk6xHPoaoZoY0MQouhiypfN
OUJudldKoxKLHECJsp/DqoTjL1xEsgC/nCrIg7l66arKBGE5wXfcF4AyrLdPRxwi
gmnhUczzNAv4wTA6EG7geilzV9XnL/x44oefkf8tJiPWAulvROtdgX1WAap61J8o
DoQfiE43zQYdoyx2dDNUT1J0nEPImZFfixyfgZ6WVHrVN1WGl/G/ko+VT82FnMmO
DDGDwvp7NiW68LLIHIL5COfBUuhi+Rc//J4aq22vHvcRQKNrTlf6glUyxoEX50Je
O8ibT4PUwff8POYqQolUAeC/I4/BPJaYzxy1adVcDW1li67KOrjuY78QpEaJT+Ic
hoMeu3LWfSDZJn0loQA1fD0H8BkT/AjtZiOabxUhAa9WzWMS26Hpu+WjyjaFtPzB
6qxkqiWqUMXnI+HVd+JXVxcBdTinc4/80A8QLrKRfEn/Y3FuiRBoB2D6q/tERs7W
agMfraJG2yTjKKzX/6qSsq1Hna8jiSepEFKG69MeKpMJt1UazGaJyJ5OdrvTZpp0
e44bN6S8IXgOyFDy/Tca9ixueULlOSkbDuZpFwHh/bAk6kzaP+bM39dQWfysCmxF
W/7Kml3OHuhMxnMqnZSANMlPIx3ELtOquY6T7AGHHX5/N36JtyZ9Npz0de4CfvCt
/pLKgETH9wyuN5BVEo/zt/PQ7LlwuAFzHlS5gtNJ+b1rsvW/YkZVFUfeJ6uqUp6W
SnXa0lx1dIFkPZ8Hpfw4hrN4oQrALObQe43SoFs7+YLjn0uh4TG6ee0QW6QKi1xW
jVwZoYoPYx5O0BnmlqkBeA60e/v7+J/Acn9YDlOhjpMxcxdTtT4Bczf8GRkkqsW8
biIztzfO0MQHUdMMpVtA3rh3c4teYCjmWxYb63Jky+1GwwGxd/HDuWk/NwEAX0jp
FdtbdAjR0cz8v1NvpkESU0AQAwUQX2EMmRrc34X7oK67edlSTjFI1AHGEXTjAech
5HP/YbXkcROcAcGiwuzFen/UCGr9XxW2H7LLjByraSDSPmGM9EElv9IzBqf0DZAG
qbHAEPpCfTDHxUeT2eu1zTwkTzITyU9mada80P+x7ZXmTHimOGymtTvPZau1QIQQ
VT8+6fEP/+I1x0Jz/zVu7neKNb6UpXX2hOKXAErkVuyTiTIRyvMS7BRNWR+el0HB
pmb7A4HMNLxn3xx881Ro6FU4zO1c6l+XG0VWsu2ozDLT9ZTThz7J2P+z/5QM1w6e
X40crAikPdAlXMw08nUwwSooJ+xMUczwLdrxzYtPiTCQzZiwBWY3sP3VK9h29FDq
5ohv3PVxRVkLzeaEU7JXbdRo2138OCJOCCjzj6tELLbdGA3lPt7WiWPe9NXE81GS
7rwFKFgJIlHkSbOpwmPZuPSHX/hGG/VFXK6IfsPaMN7t00wPO355bPNtWa2lBfLV
YHt/yw/CDJ+hMO4Gyb2IB/lAGhhI3rGWHaY8oGZdur5Arkc5i4lKcjvbsuInbuu3
WTJ2y9u6fx8hvz9hSNqcMnQw4wE8g8D75K2wSyur24dKou9cSztWUGStm7U1n+xn
qCNYZmPgk6xbDKgfVuQxlrKNdmY7A6eA2zSMFuChDIIxw7x7CHvWIOEs7h3UX8L0
0EhNzc0kiEAaCql0sIepfAmX8j2RCUNZm7xh2bGe4VN9VOx1OxKfNppZwRkOWota
n7ep8vDKcZNJ+KtDJv2f1YzgqKrh/ef1tDSbx4Rj++n3FDF04UEiqnWZjzqo93Gv
4B0BoW8RZtORXGjKHYeAM7VRUn9Mr1nb7ae4LRyDF2Biqi1eZxWYCOipVHlJrLWP
1XMTPHnU/BjVCuGOc4T/PwW2xtsf37333gQ/ApibTTDQ8kqaJBheLxJ7LYt0pF7y
8wlFSWkvthILvGM8nQfRqoalB0potWy8e7lkJUlhJsqUdnG6TI0jns48Kr5UQyFc
9BfcYfdxcrJuvB5T0YHGm3u4k/N9VBBx6F4b9t+b+91L+d0wz1X2fEhRP3QPCEgW
hpTee9yEqjxgUhY5K+yooi15rL0vqRlqPtNvEeMAjtyV1WjQGc7l8LYX4XTF0C+h
dJpeUJWPNqJr8lVeA4+HdSptrWcbCRNYNbJ5w+lm3rDre5oCwFrWDoqVhQjhDJcY
jsNBdN7yWtg2d9ToC8gpPgDKEVZ+mZirZyt/61jmJINtODJS6HfuKhZ5xMMU0ogl
7+fU7jBmAUd65+9cLkffRNZ3fJdyr+w/6RQqUqtpYfRGkCXWU5IZDK9+CX7h1aDn
9jGYl0fsWdVAsfX1yrkIkZVSbVmghak39tcBvOzVKKmX5TJ+T8BMAPjAZlDUvvtj
TWqqRxRGYfY2b/RyaTD8gzGi5mJvCP/BF/kRViQ5qtmL4f1Am2FTM7EuwLlCXWET
3JgIF4TnoYmqIHYWXYbg6KWF0O2vwZc4WyYHtssc/Korv8WHxo5h9HNyIPQW+LMf
chzZrYTO4datbjuEz4psEJhOVURWkkZwVwB9CKduYHrH2zbafy8RI+6LwZBeAXRX
YXOoALdeSlWb1mXbQaJvQ9UU0yC1cwOqkyQjPq+Reboc805Sw8ifBStYA8VDV2sA
LcrQsbPcWk7Q9/ezwANP2Za9l37O2tu6qcWTonZQAr7a4QVMMhp8d1kDFpCVivtf
OPnYDRDIs4n4Se4W+vjn6q7bYK7NCXirQVW5XwD9yGVE9Tb2MrmYUw19zy7XobJ8
6Hw3Zvy7kefUh7OK5ob4IokugYG1ALE8qJ7/Q3RGyq7BpfFICa/hGtwsB0UOjcSH
iJwT0RN8bhbC69GIZHhSAqyN1rkvovof0Unh2fG3uGIjZYaIaeQOgjU3QBAzAocs
mBApQCIuIY7dqmt0IWNlmxqubEyGebbq3AIHuMZwNlr/840t+J1N9Nf6d+mFZ8XF
lkvm1dH/K8I9vBN+TsentF5E0sfPb0Vh0a27PtFhDwmG0PLTobQGDUXOGT1b/7zV
pAKFb52S870Vsy6sRtxwY8wykDmtE6kBmRyGVxSwjuucaX5Lf9Fm+Qd0GijE9eCs
H8oxsQ6im8AJDqMbBXDeN7p5s2NVVkSowoxVKnypYZf6k7RwtoqtCCRo5nWONdbC
+cQAmFp2gtBjjbxI89g3YRL4HQDVQr3aAikzFzJc8JRxsw8xsg+C1zl/TiCKqOAa
gNQJd5WemFxS8h7sfCncXwPxbRmT3jMwgWOjpg49+MxVf0+PW5DgbTuQhdDKYiP5
w8YnVUEMXhZlgDTvQlHmBwJ0xrO28cAeWCn8/q0OkCTYzLRcYkf5vXN0/K9NImy3
IqHu3fi0kNZ38aAW04lL7WNxsKMiBSRYO75AONMPdn/f1v3ymdXUXV1j5OGbqgIe
qBf/fKrxzxmWUsU3hNVh+SGIRyY1iDGYpmjA91n2YkzCMoksdlq6Rx7En74Pv75U
/ltg+UMQJ5VOw8Y7kACpWook1bFb0kEjU5h61Uxvx2Xlr42wMGKH1hMC7FIRTX/9
ISG9ZhFs5NFj9fD4JRpR6fN8HsgXb0OzU8OX9LZfbcy5NkycTW9rBudhTdmRjc4o
i7/ueKgs0rX92rCZfSso4BkeX/xOmPs2pNdUc4MvtCCgU7kOZgCsvpTuGCglQQHS
FcmUtahX2M0gKU8VNGcaMs3EKPngV/AvtbafjGg6xX7fdMM7HXnd1CZM5jUJUbE6
iYkVF7olDIXFBrET7lmQManVgNa7XJUSAS8Kzu/MlMzrXomqGSU8lvUdgS9MK+iM
5LE3fneiP781aGXxLVpj2FUmJw/ATmROTLbkOh+SdBqmmjPX4m75MPR0sAkRCn21
r0Fo0EeZvBJJfL/dERpSXfmevlLZByUU6Apn30s3iSIUUd1znzAduPPVp8tTRoa3
rF5bgISPM1GBHHszfVG/mJXWSwu0iRvzBLW4wRn6Dq7MhJKS4NE0obM7IPUgcnhX
tL8DHd6ZVA0uuhkXxTKymR/xn9n9wyZ156w7AY5weWRUihJgSEm7QyxmJwdqJY8p
6qksbybomtQN3UGsRpq+xL3pXyeYw10i762Se2tw4rlTlcleJ9JSX3K38U0P8wZp
HWXGG/O31mR2MDmAFCVxKdJqMpPveF1hgfo3NMfapB9GbJcXUVNyewljq/XYTfT2
UOSiU5NWsWzVe0lGx9kfSu8UUaLP3XEjMj8Z4lgZVuWJxi0ke06l43+HHpOSa9lj
p6TukUHBzs8M+YpncF6pU3kpEKLxqdeaw653FJB8TA5Q0XOLDmYfV+/I18lI8Hp9
Wm2Xx5edkmcMmjRF+hjujLUF+ceBnqYpTJ9qldQSfDBFwJaCGjSgzJBFfuZu0c6M
2q8wvXWs30xapmQ0DRNknJYzkC6QX0f2xzS04X5wgXUHr62pjMqcLdHfasoYlK4C
lc17geaug7GKbygTUX+oP2DOJzOd9/jDcILnAOkOAb0HLRGG/drHUaJRX2zYLi4Q
aZyUSlx9WRNIUjhBZPdNGl0FDS9edbyia8dNhgIcM3GMnFNuUDSrNkYD2YIpvVcq
orSxUoBRFy2jm8mFnLY67833lV41NwGiEhwxM/8l3pvG6Wq2F99YaloUeiQPImUf
jgjT9/17LTiRmKJstrDRrxyu0sFhm3H3aw3ukZqhIIusYCMKdnPQQ+mryV/2PiKw
5v/g5c7Cdp8eNZ4ABMHc47kjEJEO7R05rBHnwZmPkSARhNefzxYkXBMrQffu5yU4
HXoG4JaGrIwZAtlFkVFW2hJKw9dy1Df1Uv78CIMepRNtJMIsyzO0ZT0AtXEVabqY
KQ8qYfhw37Z74+qyMRyom4GK0xpbxoEsRMaDYfRI8l4aQZW7opnrCJ9NkiKnb8iH
L4sWF85DkxjgtFVLBmCIATIfKHGCcz7LiPYyKJ/50T+Fu2D0WsvqaGa1imI57/on
sQRf0qD8Mfafslgsy4WeC8kDisgq2M29RGIOxjNmRW429VutG3wiXSrNipKJK1v0
hXHfOFAzudKMVSZR5psBQPcfYKwFrFIi0ZTu8JZWv1hX/0q1jhr2pomQfiIgPGAQ
6cOCcwYWidBEMCgjFnFJrRscFiMnIKdV7/jKA2B3U+dOgtapx/msKMOfALR1oQfF
9ex6CQUdv9RF5n77Leu5lmiqYvg1UD5J5MnhlmpJ9FIjbLM6H52O6SFz09g6UXiE
55qDEhmOx18e4KDlvsgdGpXpz+cwYXCfyOjfXGpo/ypMRj2fwckvOs4F0M6yaQ5o
bL2W1G/2SGjIzfB5u0Ktw2IHO/SYE//fWMkIhbCggznxQ9hkqu+5Qvm9tGiSE8P3
AVNkmDwaHUCP21UgkQe0e4nN3Wgg0RhHtKluLrMcMMrozuz9fhgz2vcmSE/3Q71Y
a0oorEVUZlPudYpfYxWXh7Q3RKksyK5pioqixdpFziriv2OvNq89SOKtExcxM94s
ZrtHTz5xDGQL9d0iQRzFP9XrmZU7liICeePKFjCuTPHsIVRajmmzG8fUVlSO8qhE
Mharhosxr4aRyu4RYjjRwM6fLxSGQB6pIfY9TOJ4IYmt6pVVHS6pYTUjXW3qE9Pn
JlKSE5TPVzdyQjWRvHe3nRg7S/SrxU7ESI5/HygIC+X/LRf/4n9b2tFQVAHeTRe4
FajN+iiF1ZpDDdaZEyxpby270Eh75UhN2vHxtarts1YQmH7AsrEYQ7Y9p6C26Rjz
edXbcBMteMIpuCHK3oMdJNibY2/yvXBKDxjao7nEyLwlpX6NyxrATAs/aTvp7P4h
SR8r/rBSFLwPoeHsQtDFS/V4iC4trOeTxhtnDoEj91oaRCXlMJE0uPB1qH5B6Xre
SZa3ksnk31DrhcUO9IAUFzvpFe9RhNTI/Ptx5Oe0Vzzn2GcY/MkHDV8dKeG+ZeGX
Hv7UF6sMdoFd4FH1Jcf539DKY4A2lvLaAtPqCGAEv6rKXRR5Vp/V6j3PG5fQ97zp
uAbs4pBVYHRVCHNcIC1H5pN5yVjWNR9b/jjYfA77L+7+SxHReNUMt9ZS7cjJjuDZ
44O5nQPiVs0XsP9oFHw5KwMC50w+q1Ebeo2V/jazgLVDLNKnBlEyNO6udnEcTNbH
MSW7JmoS2AgP3qSVT9EjpwQ5iWJ9ENxfqTA8JNcmQLHSx3awsVfsFIPMLZ9VI9zQ
19pPQypBqz89t/VFeicsb4rjwWfgcDvs6dy7fXaQQOXi+htPqyeNn0DrBn+f7l+5
pSZj3QOYGD8ob+0C3RAESVDAkZo+N8H7c+7xTOQ6wW43xypYgpvaH+Bagn3hoLHo
zq/3ewh5Gbs8Y8mm5LEpGhY+Anw+QlSMz2iufP0fY7qnUe9PKI0wQ/6aPj35IJNu
WOHzSMQhHvroTL/xFNfbgQKlxbvrlEZTCSdLrKXiHjR0e7CQLYUBKO77yPvDKCjq
JX3lyHx2Ne7hJkZ7EDGrKcGyLj/EUXwkmTHANxLE51VMeUuiA6YKLsrVbMpr+EZI
9Dlm2Wa2UAtzsctahNm1HYRMHpUDVp9dbDLv55FrUIgRduWBt/ClUXzyJdkTOrmm
YAYkbewPJfqiG4gESDFvvLyJOOllUYbkiE9PtI24KqviQVh/oJyACU2zIdEIBKvY
jiaEIO+Q4gpiv1ggcAgeUfCNHFjC+R1Vnftv2zK878izzON9G5GXs4A9YJjJ2N6M
wmdVVyysjh5us2ne0GMA0evVF+bmohkSYLmf+RSxHFzR5AAmlTzPBYcE7werkqaC
1hTDUy05d0rEpGE6CBQm3SuRW4MM6Qc8JuhARDvaNQKA6mKQQhmcNIdYznSpjwPt
yWy7yZ7Co6za8A7UGTSaxGijCrBav6bhTEd8gVwkpAgtPIPupxc/E4dx/Ubx0/Nj
0aU8IzkVeS51grj0LOJCRn6g/oCNBNVuFWtESaNmtT+PZIZCk7jH9hrpNW6k/a66
KgRuW7lg5H0QqV9NdvGG8QgsFWz4HLtOCmiCaUNyxX4KUiIpomcE5GYdm2j356gh
dvyN6UPTVLYLHKc7QbDLW0DfgVs3lMo1cSo7gE4EzgNdwJJ/yM0tfzSiGpTRc+Cz
CV+0QKMmFku/lop3ALdbHYVKzQ6Y1YQEgd4ZwvAvWaGWb4jUsedIwDsOskEE9NnS
8ohATBs/RkJAr+vKhYQQC/gd3ajCqe553s0IYzpdsp84N22ChbzO6orX5l4s24yC
lKgL476YWU+oJWV9LS7vlOwYMRZ1GdNNx9W2lZwTSrSYlZLOeLXDhVy1RknCKOkD
kv2XZ24Fr82A1awaCZnsZ4L39dVN2/T1OifJQUmN4FvJ9hUb21On2Jy90woP/PWf
cYX7/gbHjnLQyndhRIBKTz/nRO6E2qKshwywRlcZ5O8ak2xwXa3LNkHfKuNGyse8
NDvo8W+/LS2DZE3XSFqgQq4Miwdu++/yRp34qcvFgBLbPRqlTFMdJ+R5yuMFW3Kf
bvMelU6SjAhzYwZtSTcxLQskZLmD6X7vrP2o9t9pzQmTxxazyQjgyTRKgrwf4/2M
DMxueSCvnufyli+fGUr/VwfiDX+wBdQqPAD4+BGJoiFifF9nBkFNQ0CVmAIkFE6u
4I1ui072kiGKnjoBjFjMoxdGPOXvcMICEKqeTZrigdH8fYUqzML1W3ETjG2DKPrb
hz2RQqZjz+2WBg1DPg1raGSG99zhIYxb5tKuWgiBl50D0KPtIkrj2lK8jJgblECT
/RYcKKBjQNDoEjuAw83NXUn0v/jKKFitphkbrVshyIEJQRs/tQly0xU2OfH9eF4S
YPW/fKF30gypGXIB+a3JR2yOyPe6b/4dcc4gINinBXQx3u5/7F8VgCo3JRZI/CdE
RTPvoKbb29AUAMdET9B2TRQ/+Kej9ImJJFerW78lRF3bOeJdb+4Nrbcj5pjyL3A8
dbmlQMgqGWRyMjIhwdMmUfk/FhyoBXoRc35v3hFpOj76jG80+LFrh3iylzVDuNAZ
zNB2m9/qYdrC2CsozKhcalMbGsCTOlYZ6w5TE9kgZv/syHSvCirgFR/Ccr5z534E
8nOiBTAJEdcg+bLJwULnjLlJo+66RVsfi4GqyjDVSUvGUE16RCWls3VcF/d+98L5
7Qno31edHJRH2cqV7folLoi+C3cFuwy2J4eBg1C4gtHGOm7cbXJakQHX53aPjm45
FiV5fJ4VS4oCqUvVLtWJroOyhNVSUUrXoAYAmaNGJGBWwO/kbMUX08+vjdSxj+o+
V/dhMbqo99jwTkFtBI/PzXArwBUL36q7BGLGtvcOTgCgiXpp0IR59WL//B5PnnbB
z7z7n5L792I+FtqA8R51trFOcEJsh3PQZACesTzH4FSefb3DnSZdjhFZ5fpreUgr
J9jDf45383FGLb4bnXIkZuBfV+nj9TDWTWVQ5dvkR6hgk2Jgb0VxqELHbWFcIULe
gUv/Bfhoi4SuRLy3pDwzFuAYMGDfon5yP1RxSoTY0B90JJlIPpKQxeiLLq+YVzfG
tU2GbqrH/FoJQUCb+gGlvLNQvOAriEnXaXTvHQ3Sr0m9RilLaj2TRulxHjrnCPkn
jVudawFBX7DqEad+2/JK0XMJyw00ai3h5MpWhzmTW8SdzA33tiOrZGpt54VUo30m
l9eSOhCBVcpwJ412Gfl5EOiCTaOqQ00gyaIqAhjx28/UBotR6IUSWrBz2aBrVaCY
nroGwYjsyJDDPRecjgzTMRq0oqcRkPzFsrrUsMPBPBdZDKOegLx0gvEFdZ30fV15
Me6Euj6Br3J66cEcagQG1GNqGTHFbGWvyPXV/oMKmysWRu3glVkrCGov1AbHKADp
iP/fiCBbofDj1rQD6JoTTQhSI6iCXrgRvtwsefPjLKQy0ziCGI3EUlS+jhu574Iu
7dzmdIQc/o1X9CxLT1Dn1dMBPUJRWazKUOjNGGwsnG+JIcl8vT7nK2OR8Bibj99b
p0w6bpmnoUZJCZUuTPs3xhApgUSIztadbXgWVD7IBuuDSrwb3+9P8WwuVm8lkN6Z
AHu2op9Nhdg5BsTrNi/AfF5ZW7Z5+00+b6iBgWNPfPYPyt/5Gx+DKk7RPOCh9Pz3
fCiFqnUHEyBUTIQ2MOMLY3LE2NwGIK0sXPzaZCPGjXIElmOGWWA8V9jYV9Kp5K/e
AXvIHku6QqvmGuzrDWMv21wSK4YuXyHjEWVYa+Rfn+n1ISzKLIa7HcDyedgwF/ZP
SYw36rim7wOj4cNK12D4QnBcwzLgt5vUR9mwFND91F4nny1IM0hWxpOpGqeUK8rI
OKNQtQJSfFnHYqafULtsPdTzlEv3mlZ+/rFg1kL/5A0/k9YtflcY4XUISrpgum89
ZwQgKfWBbki3qQoe4eKDLsGca8wCyznDzrWkYoN+Z1980MilzTjz1qLaZhS3oPwI
5HVyn2I/MCovCMejL/iUEKiXM7m9a4/cmC/j3Y5xNLxxxaTYThVSQY7nENR7+kp7
5bNbPL97+QxAxYMH5y2S9S5Eyai99Qiv9xqROwjsmr6s/MbvHHkvC01y+1BzrpAw
ZNsNNknkJd28Bjqtf7v6UF4KaOhYf164CTYfs7K194uKecvSGDnXh0ANA21Ilxol
ze4q0dyNAhpmECtteFAxCKGEfQwjyHVB/Rkpq2eqbBquqKOMzVLBkrCkKPge821J
W3mQR2smPZ+ZkmjoJA+8KCH3W1hp+u//OPWCfwpTNRnGEhOklIwhdzTQu+yzczbx
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
llLNGEeKGaShHo0IX+Or9EbCYJ1nwiDdjtxguSJfvb7hAiGiBsoZ8FtOdRGh3Y/p
mS/ts+ZWIMiXeKVDtDrL1JyDnj+jUdu/fMDc5COXzzmclH+FrMrCPO2nFIXXd+7p
qFUOLmNERUbWATIRmM8fkmPgoTrbAl9zssgFvRSwKdzKDAABS181326q+uD0q4KJ
7SFlyaEpN0CBjGa4oLRyQUnC7AfHrLBtkbHmVn8nyybqqkuHtm8pUQHh4cjYfpMX
UMejsrdtzl7eLPl1Gaxz0bF7H/fWP8Us8+lw3psUOrjYQvRw6RWnGJrgaqXqeDpl
hwFo3oJJZopGGiLrECIruQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9200 )
`pragma protect data_block
KG1qTpXD6ytvnjyIYfnjlXlmGr3JLqPWG+JawCND4zgaVxXPuxukDKeGJS/pejmY
iPqn3YGEBekaivsUWNN5EG3NFwkR/Czw7JCTKS1fMJY2o9TSwvxy8PYDAHyI6E5b
gv4Fk9mr7WxMx+dg9c7rjCtmVRq+cHRju94b1ODiiTx3Aan1B+P0XbxNvjF/a/v7
6uiB7MhG6/juWBA/ZKASfD6W2WKe20l4aWiu5LIKHteN3ybhLeYRcVA9bHR0bhY1
xCB/vssHEkr0lUpikEBaN+pR0kXntNvC5t2++dvOJO3jMFNi+Sp6zjKvQK+s11yV
Th/pGp6XMPUyEffrAGk3VDbYXfXDZK0W/FVIvaOPLKlEqxFYyDEqMdj+XbewlVMN
EojbbzDg8Hc8CkL0gyvta5DzjhjDJgqibbl+F5p5szEio2o79bjxrxSUNw9MyFRa
Eu/HjRFmczD0HFyWWGHqwuG7SbtSIGt0A5nvDrJNXwzE36+n1LZjF1w/FDPSj91D
SBxlm5ju26lM5tPnYl4KTW4B/Bn6ktcp9ddn3SskNy1r+LlWP3NC/l6N88r0GfPZ
waGe1BH1Ggm484SLHK03fwSKftdauIHwvh6ZaoxiIk88T1fTT29s3IvztZBx/sr1
gV8XssUG44aG5P0jD2jMhGAyXt47doB5y7uYyiN+bRugL7aPbTr8dFNwHYojC6UH
BbxSCBunM4fbIIeohVwFVLL2Ps9kbsZmPyZnxxK18IurojbmKZVYSiNg4ibpwcwT
/bNMnO7wCDzhucXqWerTICIFtN2p5QaTAavjqwpZEdg17Q9wt7XUgPFVv2Q0zidb
haNTb8pUsWWlCsrevWhlnsd0DkyzzV3Z/8GzjJtm67lSqA3aG/XUQUQVt4nEnxZ4
NPyWlVCW2FxhsIMvxhVmqIk7+xgvFx9HVoil/Nt4+vrIrNvSWS4fYIReDkEVL8Pz
VdH5rK+MnTgE9938RU302VPz8CSNgn//kAhCpnN74YmTucLocQwCTPzfXEwhbUJa
9Yv20Adri95IxlajCmKxucmR6asq8Txh7b/5qFRjloOf2fJqZpWtFwdIva0SFopc
GB4jdbZqZJnB6jQFNkFZq7bEcEICaqjPMxvs1u4gYxLx/yWh1aQXFlXqVJLDSYU+
ibCnSa6y+f9pfZlEWAC50rpaRiNHqqFAIDGdPx1e0Ch/yYXmBcAcRSZNLVzbZyrp
q8L0r87iR09rb1YwaXbL3TZrpUtr4NOHzE/ZDiikdRPgJmO+rUFUbaRHwMK9/AVK
pQLHUknKq0UPsIw0IxH/TPXTMylZ6INoadEWN1xFNxQpmzIP7oy4ZUKOpkvPagFT
qohxTU3DGRjKA+DP/sdGDbQ1prNXHLIfmMIO+IfGaUA4ba7pMxHQbDMfjVQ+7sKf
NBnOs4C2wtGrgxs8Iyp41TxKhvK59ROA614v8LYvPpn7TfEIr+EcEs+GunogGD/k
hnS23j3HKPn7MNx5GW444rkdAP/6A4DB/DYmchyoVco1A+DUbdAYjKCHMZQ+Q184
gAVK8e8cyXOEDecqJI9VtKh8zGx8mhDo7tZ25BojBzJuu/96gMmkYbZ9JuzBV78b
ZFN8NNPj+1wqQh5O7UQjWva5pW3uq1Eo6glia1TbmIYcaNaE4A3q+Asq4IPVceIV
xC+j1MjGKgr1GHH+lYLW8LKlK2f9INlTQKvW5MxwvyhIEcA1bmfQU+jYWYIS+ycr
OKPzCMHl26mZ/mSecf1jnJ/08I7UBMSwejsKhpNaumjzj3gSwYqmSwcPk8pa5c4i
ziqGD/cFANxzpdF/IYuwwKXw+lB0QCL9nt4LENvKmZbaN3INCj/W/Ox0/ElC5ZX9
MrCmetDHgBqebDGe/bahHFmRPtIPSmsfXUw8ucqW2m7LJpkQ/nN1mNldK2XfhBwN
nMHFjY/QYxNt2cFUOeOf04WN4ax8nV/kl+J6aNssJNfzyp4wIsNxK2bX0rc+iDCm
aXGVyIfktxz21EMhLhQyWGO8AIoXMcc0XZkASZACOarZpyFKFYaEaKwBiuLaelW9
/VsjUano6FMJMSiEkIxx0ROjuai1fVkQxDl+3l/teB3PL9XIWaVsKi9UG79aDrE/
F4omHceKA8xyTmzA0l/Y/eKi5L3KUnrsbkqFFqGeik1gur9zDfcsksGXQKsK17Tt
MIijG1pgFUW7oqh85DjNDlOqdqIzUXCpLFYJdgnBw0er5sEoo3Tmo4TG5CVooO+Y
JnZm7tEyJFcQ3Q1CSil5qAU4rRyRWhhXKK5oCTCVvljasdy+6fiSFMRefdgdDDgO
4wOi4uYZGfm2Q0S9q9sQE0TloouIWcx9ppUy167/BQmDgDrupArYxFJ9OiAf6pXk
jZ/vWOBEYR7+wUGX8g/0k26DVr0G32aYMfVhdt2RzR4Iv+adSkTwu8Dxbu3CO6Tf
/4Jrw9sJ1uL8yY7hTG1T2Ku+/re/IBrkUfqZ6muurj4woHcpArvhnaeBogyeLNIW
t+MecPuMnx/ewcUiS+DF/lGAHgJ0r5ulvWH0gj86W4YzSymb+xy9vp6c2nE7pKKC
OkDPr9COygqxBqmHx8/fPW9O1ax3ZS0TR4XxdLiH8ohGIDYunJ5bHl0MCSqD1SZI
bGKLmqaHNxvAEkqFgv46PIHFR2H9PpYyt34DGaNbvJBCuU9ok8Mj/4bCPs8IptTh
6bPh61K7/77YsdvX+IdA6rXi/ehef0a26lm5nW/h78sCNMAsCaXOTou7HBMVdHlo
by1ajt9OcnXvssVPy+Yf6/AfezqH4WWgG0oRXtYebS/PImSHJIW0OH1q/2jtFEeX
9v//ja7wjo0D9/QYZPrCZf8T0Pz5p5WX2AU3crg8rMonHVhMkBf20/ex5pz0lstd
C0tFT12OMinXKibtWZ48UphxjN987Fr5nrLCy+iIp3szHfeQW8qAvoDxR5Ha69FF
rlTaHJ300i9uxT26Tn88OVOaQPTqEfLA1hEX6qUXJyzZhtitsoUoVEGn2TM03AWl
V9XzQMre6BSDsPmhbkv3vYsKB0JwUENAC/BgW/6UQTnkAyaDoOe12B3AYii6ZS3u
Tu9m+DbTWHVgBAqQmcIL6sCYrWSRyBDzGKbgucTx47j3VrlkVBncFel+zhHExJT5
0ea7jndAznlf/TsRSraXeqUhH1C0qQ8cstbW4s1U61Gzi8B1ofLWTkJEgGeK4hmk
/Uj49plUF63nxqU9SgcOUTeu4Abs/MeYm2zJtizCVqfjm3f6VSljitmYNYh+UK/K
7QirjDvKqUz9nSL1V6Y0E3/L5T6XOD3y60Qbt732wer4YdGi41S1rQmxv7ntI74v
O2fdOJsApdsV3FWfEuEoBr0YT++D+03xEklpA4bvrkzxpPSl7wZyr75Nlo3IeKjH
U46h2Z+ltadlee/U45F+02cw+g3ShSnNG0OB2hYvJCXHHNqRWqNC9yOdXVEyvLuW
yKdwj3Iz9j0V2AleRXXeEuXIwAZ+1bnve9Lw9AppSqneIM73SSEKpjHgdSAQuib7
sbB+orPurvWB5iE+tny2Jna4L6OR8hUSb2FHlbxYdCxCF7mcCv8csbeZ2vxvwpDw
nKakG7+gMNtDAgfv/fk4Ki3ycuBroiFKGJrhKVz7wMbcOmpJSI1cJMz0UX7KQSBs
YWltSAV7zAcRVWH3TOVkoVu9lYppLgfu3R5qWKYbOurjoUDORWmwktutl9ll/SiI
5Pa7A+JsFtVMYGiYRca/TMJ66c26NXoUacGxhRb8Doe5U/FJbtB8rjE1QAnuE0xo
KXAgdI30y0ROAFVBktRYT/Qfr9VbiQxb2ksB3vomhmS3SJJeKpffs5D4PEP8NqYN
RGPBlB7SMkJpEhx8Cp0kYQQKnost8GLGacafKXbEwF6VNBW7lHojWRjqB+ubpvIu
KKhuFnH5o/kWDaLkVLIRApT708Dg8THHCyE4crj0gV3njYPlUuH2E2jdqFJ7+Kf5
n9Ye9xtJ5Z4owB8bHsvt24Yh4Qth+jqTk1mHagzTwhcxPvqBdNsieafZvNjhIHQ5
nHu8cz2+kTiHpz5ZQthVp+s7KV286puIdpeijHeWc9tb5TwwD29Uq9Q5g+X71aRD
UWxc8SCqWRI9SdUukVmgQSNJVj7WqqKA4yF/o5u1+P64a5jxg2J3syWENn/YUV6b
wr8pY/G8q5rSQeoFwrzls1VesEAVzz7PLH1fTmYvWuhZBgAkE6XNRfBsxwLZ21mh
Hch4b+ZzM0nrjPTn6xlRh/TXkWhIc+8JOQ9hDy/ZiKKdz3G3+chm6gqRKcDp4mOM
SnQZy2Y5dGMdJtTslxsXSlczTZoSvXtv+88TvO+aV+RzGMUa/o9pADaE1SNtIyLn
DMsqAItO/ZdCGD8/BDsz9tceagVAcfm3mwjYhIJHFlSIFsoOpPvlYNKaRfH7uOdQ
+b9QgRU2o0E1lzetHqPEKIX25SaTBc40hXqFlBhnCtStKlbVOtqtk/zAlUkVhacN
JFT4iZa2v5wFj3wF9UE4mVf4cfFyDXoZasoD93j4H3nyfgzzjVs5JP4wheNptCN1
RTiRTXPDvNpSSa38r4VsUY5PTn6fpbY2My9VYedYIZlAInvR34PFfRjL2MRTkFbT
OVwaxxwXaxpEZDIxu+SdY+Z+Quz2TKw8YWivLhVvDMUVm4eaEj0LqAFwxGKNBBrF
oQlTziHvcDZ6Y9lPm75ZdxHh7cNf2koZLBYFqfP3WhClKr9IcvRC01XC/dGLYsN9
86b3+XQqADEgasEzqwCnBtRoP6kbl28lVcZpImUvKEJGLurHdLFOuk0/qDFFMoPI
MNm4jPKtl20AfQJOqif4PWqqzb3JUDDXLgP62y802KUqj5mkahDTHt4uvfs8qoMf
GsQvmQWDHJibRMBKFPUluPKEIs8pg+vnPWJpEKgZmA0QDFtbKwi5oa/8xI3DhK1G
WCB+qeeJoz8IPbWaPyXyp0skAv1i4kSOMDzJ2xdV1JksVq/HlwHHmSZV1zpljs7R
c5Xlc7RrOJNzxsDOaQpAjkpkVLOnsCqGVGICewrm7+6zX0JAXAji5JEMjbQEUbM/
NLZ95uMvEkT8QDblt+JXrP9+S+Qpdk8ruUFj1tfryjMuVJPIpp3ihlT+SHyudr8P
AarDlLbIdvbd1MExqzJU2+tJMyRuPrsA1lTVRvM7FGkM5d/j6g9+mn8D18CaGPzK
PbalriG13lMSU68ZRMXJnaj5Fjz8RfVSOw2SbezBOgEPeZgQUMHa6x5LCMOAC2Rw
DX9Wp2dCvAjXUgZy16An2YmAhJiGVkKm2o4VuKniTsaC8rmAJ8kh3HeYj77WxgCE
xcyTHxu2B5jsYZKrBCmaHpzzO9j9P6Q2JPFtoK4JUNslcodqFiVe/2QHM1SmK1J0
ik5++RA6SOuzfPaT4lzahqG2wZ/Os8ahrSzxB4sH5iP+uITue7PxDmLvmSnr8/fd
BURJmomMKIjb1lmN2Ygk8YV+eG/+G5+UPEuV1IG+60A1iCwdv0EtUJDA5OBUIiKD
uBkSvhA1VfSqunfd+JyEwy1ANZuBHqXU6QTOzulVf/p6SxMcCBkoDmhfONAix918
BNxUptSyo1ERXtcayAZMVvwrwlBlSMB4qok7AqrCvwiIpKMWfnQvMOA4gnUfqIVn
lqoy7UZY/WOiz59OQbgGL+ONQLMSqFaOWATo2F5wSkeReKZu0UOu1Ewe6FIB+brU
ayCmZ3FXhqsUgOaTmysSgGJ6SKg7/SUOOdW+HLXEn8M8pTHx1DLtyKqcpDCk0N8I
0srR4Boq9cSrQF5Z+UF3HRD84xORSQZLS85dmf22Wgz6FcBgpQIZjILAHUlENFAn
sTltW/4RmbU1BeAmVL+0A0RL2Cso7CWChk4E/txNoA8lP9AkksQr1Q3A5HYKmv/M
qfKLyj1M4ryd/c0QEHCifxMcTwSGx0p4Vw1T58K0GEjt/MviJtjT1i1jXQYWpU/B
oioxmUr0XXiDnxJADb4Hct8uxlAJeHYEi4UENHVkvV4BNRlfWJsKeu7/mucmUkBK
XMJ5YksnENYeUcAtk1wYD6GD+5xkxJx+fAquRfiXwwudmQigiLYDr3MZgUgh1wzf
+p7gVwE9qoPHoLG/hS4PyC/UDw6LDF9XtdMfl3ArVdwbO8gI695JNM6XqYQXgYIY
L40PNYY0zOdFCsXaFAeg9taSoPUVduHyEZFcb6Sp85m0GUfc2Pkh5SMlTZXsQrjl
usFJg3MF4d4ni8wF1/1xlBuSYFrMQ4XKNtsPmVkwjpkkMH/88gvOeh7ctPpYFle3
aVXehj1m45MLYCUwBv4eG0keA+falMDO0Fsz3eWSMlihMD+VYej8dlzlBxm+RORz
tP7mTyXUFSkM6T6fezTZuXWD83zDijT1EdLqaYU905QbDhXMqwO+0yQw8BWvksZL
kuGCr8c1Y9voW92yJ/APqXWUDzUi7I2gMW05eyZJGpkbhMbx6bS231VEjg/6jxLj
QIsr9DKKQ2V2e7VEsRAED6BN5CIVeeH5v7acWslFSZj+zMDONRkUO52jFdnhXkbH
c1qQue6YGfTln3cznP8iiX1C3fPIU1hw6HwttTyw1FV1K9hbzWkRlMGF+wxKWWn3
HD5GjhKop8tL9hVtOJA4pclI2hPmIjIFYZlNKLx+FhHii+jPJRp17Itt2WvBbfBL
ZG9nAbwssGarQbsTVRgFx+UCfsdC9rRItPwiGNkXqg7e4nhblFJBjlS7ToxaNuvl
AbgOue0wCe8gM4PDjAwiGtC+F5OT6Qg3ihEmUKFTkgV9cBhCsM6KLBT2Ignrc3X3
nW78TuX+VKBefKc5FS7X+FYkXIcGzv2pdBLUaypR7sRDcSKmO9zvheL3dSuBzFau
0bovTvMQsuscxYawfSA75L83tlYaR0LlIABXJzKYzDpgM7cUYBHSGcbMNXtXcMia
FFJtdoJP19WJMnT0HyS2CjB40zpXZxLhMWsAhjaeKp6AsBJtaH3QO26ufjyLj9qX
XsLM6cxjXoQwWdruFJnrIVej6V2nFcBdRvu44ijcybVdTvd7Kgr7u6TgLUqsclWD
vh6TlcbjhqPiosRd69lubpYGGjeqWBdhMDAa3lTaqNbsev22STq6Sug8QSJ67HtL
2AHB6ctW/QGRB227J3VHMHVWwm/D3LYSi0ScaM4kn1suGsqF8P9+MNQonv01hrIO
TWLeNMmlju2rj5m+CYEIPTZgnyglakU9L/6HxtxGLtPCIRDhF7mKzv9bx0BI2SC4
ihCF3udRs1iZ2HLBog4IX1CDc7qJXgkdA+Pxnlk0a+CUifu0Tlbcouv5/OF3qBR7
xv7PNKdkw/ZBc199yEViSinchyj0Hmkg0vRc88UO6Sxf7ADUhbD62/AwnSDj+f2a
08coe65SMfAq3I0eLlQ8rpsVdezUmMFfu1rL+puizA9yxleuHx50ur0xGoM8VnOJ
vfWEKi98TvbyLKM0uQjNM+1pAaHK72bt0mr8Wmk/MDllNB5WS0weATYNMUt8b7At
OXmQQhIHyWtwi8Mdd036C61sX74fqvebwwWafBGrCIPWVjw30/VLrowWEynAX1OT
jMkUqq2ydMPGw4EAzHUCgAad7qpM7Or3Q8KEWfKkUAbGWBUWV7IRGfBF6MZYkXhO
xVY0iVT8mtjSBI/4vvEht2QdBW6cbtmDw6qy4N8gaDKxPaYcdYeIe8Z6iaMApm6J
as8VpBSsPjRCXAcoX4tEkucSfip5M01ftsOh+TxVGOWMyOHb0U8nloaZA0EG33KT
L+3OAMl5YzKk7UklvZiUwgqvG9He615OFxkAFO0si//s8aeu0c06ECsjkWfYHi5u
PDzwh+lwKDOZhuRWCEnBmD8ofVwKNF33rpKMRU0E6d44IWvbh0KcRqcV6zS4yR6z
Tad9gW3Y6G4EIle6e7RNIA2N29dBkfJSd1/o4ylIMg3wohqGgQVNytucQSKXQsIM
+6VKhndd7sRtdJFMkv0df9jYA6JyW6M8PS0sXJA21P/WANgskuvNcm6AuEazVVeS
6ZJkvI+22aRvViRQB4PVsfKzvgjr2RhAe4mVFcl1tcQYrA7cRqDSmNJaCoWwnlQW
YygmiIVxSkTkYFy/ge8aIAvshYwNT0Ub07riqDlon7uFoRTtaLAVkgG0Y7rZxlJ3
e7yB0PoV939c6zeexf+QHdhUeVZ2ijI/hrJuoksdexAJVTQ/GbYIgBhs3sHlvOpu
T8FmTh0RA6aRAfk4kmfV54agXP3iC8fyWomGq6d4S+0160noqAWbv7IEzBF92G+K
T1lCDw4c4gMrmvY4Ekl6vH8mS2H+xJ1/N8eie3NiwaKBAi/ofmgZ9O5+dQJytAjh
LcQssZ+24noOtSixm3dq9IcUBE07/HnHHY70vMm3mhCyoUnLvTzHh2S3KUGS7kBk
9zkRRzw9vunGyCmWYCI0zNfN+9m8MLwSuCfmMXYJRPyGl2lTkx0gKl00a21bSv9Z
VuTOvHO9tHYDMAlMYNOWY/BmghL7OwK4bRi4bY3oYg+jp9w+X/pk0+QaOKrJFXj3
Bg0P7uP6lZrupDysLMaU+pTxuawl9oW6CJWCBcsiauPdWfJwkLyjCCHRE8OdXFod
ukXmKNhM8oBAiZQuyP2df8jzA1S4na21OFfmxHCZW7luJRWguo2KZZyWNGp/0F2U
y6/buO44AYxj7pjvvTuglyQ6wUgzkhIITkRRwTpYxXS69ObdzETvfeuJdJ5CXV8W
f6yhKDfaPcRL7PsCCaeWrYC+3kBJ89EeilNyUIGzMZn7U08fUAGXPpCdk0+plT1T
EgeIFx36cDhUD9qqCqUjSUhncB2uraFA67fXeZ7E5cszU2TEoTvjhpLapBNVygw8
hXzUvLPC7OR+tuUYAMMVLYKfmFCnu4ilkRJ/SSGL7twrg/Ds/FHi6FTffH96thC2
HSgR0ozCxsWdjGvhYTZ6jzOPNjHX9def824xHo3WLseafmJWbfno5lgsEJNPom8z
KiI/SSt7L3CGsjjkJSaPkEEuAKE8pJbKYBOUVA8Kzmxx8Xvv1H3EeR+qZM2bVhvv
ASsBLWfDd2Z/31Sq7nirP1TXTqOvR8OT3ekbEtBOVGRXIo6HKzWYs446DlF+jy1z
IXk/OW80isT1PBy1bFs1XV0wYTIfNZvvCfP4Nj2q2Y1AfI2xslkZ8AP3d59JyEa6
VH/HdfbueeVq6igMw7irfETd3/mA81prUCCRIGqQw7cSmn8vcrs00o8fLyJ1srmx
iBYut5kkjCsYcz4DLK197pMOPHwBl5SHvfrps6YJynapiCeio4CPvKoxLP0XrtcO
M09+nB1TRKfia0Pywt8+dr0RX9HBt3ZSOMBAphKRrCBpapd8kjV3sidMd8NGvf9P
YrFnvja9EKr/sy1bi2Rcj03ThB7ppq7l/AdU63tiPz3Gzr4CUxnjksXaSG1yYlP2
k7EnyBPJYc2wRsDwGvWfiB3r+vZOajlrEkZn+PvQ/1z3d9kJoc6urghKeRv6XXda
XufCVX2LHRsV37lMb2A6JhjSpqf5IKQfJFupmEKTnseXknIZyYqYzzxgq9qMsKDP
rycjDq/Vtxv/AIrQQbl7Jz38m/ahTjLcILHemvQuAzmkUX6EZ0Hb7KEcVuQst9Lc
hZKCbdY3RfYTK2h/MrSA2g8w+WoZLSlBLQyZHb/+TWHrLUyB5SraU/DXpDDL5hBA
6AjVhz9HnabCaJ0+g9nye7gb2Nd1xUfx4iEESl2CKVNBWEMEMDPnRwy2oInoQrjj
YOuqgl6D/xhu63o/0YCEkrl65rDlOFtFlI7IHS6Q7KpuseV3rG77YhG1s5xugRvl
A0ILhj3Fsfp75f36D3vLhLim1YQhKpsUPmOzWXhLNrLt4PE24e3YsJWvVVa+M5Y8
g48Is2qdbMqrfbU1ISpZC6Zv3+sJaj0LrpfONfqU2tYl2tHrMW/j/SuLZ7rbZJ1l
45J0AWY27aFCywzN0GkXGMlivhQop+/totINWj0T7hJ+IMvii7WYGnNkiGvoIINr
kDCAIPx45vg8B7HS+TwgVy+lFEd/evoYf2i8EMj+OFeilJDYsFr4x2ZQyF65XKfk
osonaT1X3uZcXJz6pGJcKojaSjGlDewy2ILDK0CMVrnwu9bPsRWGOgqXYl5WCXsj
h0BU1K08Br7qBa59+a41LwYSLMG5CpnPTZrDdFLERdOP3pQwagKlTJt5Kut2STq7
Dn1ozh7YLFJU+g0qpIZ1TWhGH6frQLBhOfVGD0CUxWstze860ug6FZVsuldFUWAb
y8/Bx6ngiaxEGTGSc7u+8M0E4tVVnwCqTptJYy6EvsTNNT5GLGwZgvsF45sSXeDh
VyzcCt7E3hx+Tjg8yQLHrRzOSBVTowN/Wt0s7MXecwAaTT/Pv1xteBd+ZxIfEH9E
ZgUSNildLWg13KDMyU406olefjUk3ejDvg0LcZwW3rRhhIs9wZAcAs5JlAejTx6Y
uqAUfcaKk4fQDc79H58eV+rQuJcDNpZ1JupCyBk8u/ow8tihCDeG6w/3JxfPvCPY
fjagdkxQ7MF4kY7/D2RjpPqUJya/Byz3ZXjQec3mZusO3MOljLkw4WDW28z3nCMW
Zg3wmYXKP+aH41KZm7Pb8eem0s+Qs0aTKoaDzn79YMXzKUfAPFeP1jdFiY359R92
lni+6j3sgLidJIP3AJj4BlVnUr1LJ0irxyPf445LkGRlBLrvxl0dTlmEl89MUeE3
JqQPeAseTIlw8g5j7+4vFX/7kwQNRRvVtEWIGrwlqynRfE07nOfdeSMQ+pYyowzb
FwoG+RZzYymE126wfnJIbxF0BKwe+aoCzo4cCAEyWyUfTqWasIDtOeLgZ0kWPvYX
otIhnzVRrkd7JTNhCv7NGpEQmjGbEC0YiliZ3I4aMM9yPLw0F7zBHhiLAhMU/x8v
ADHhCYuqjPrwE+ys6UA9/83FSCf8ReAx9mIQkeozerUkTUbvyg1kG7ECENyxp45Q
XRNm/IafFIkC9HdJtUH6m/gHMDrbeQQAObB3e4CW0FuSChePtRBGC3hUb7CCgXBy
qM8nKkhmmq7TTYExYH1A25ced0NDg80BxK4njztdG5JlJdZvdJ4E7hEX8zCd522q
ohBCo1uiQf0FK49a0hR3jN6HzlZujaatQ7JDMcM525lZxA4KK5CcAHaUqzNTynYZ
QcBtYZT/aJI7NkX5gki2xK5fZekcpqcAR9y52hQqSh6ZvkWs4ctBVctxs435JQZ2
BC/n+LGPFJ/KD1b75KOr6qOOb6HWQyCleUCCiSnUVE4F9I0deQ7o6rheGGjx7u1i
F9RcJU94hWs4Ctc+u4nxmEgQ3cAyOUq6Gr2R8coI9PpnnAWYi9UHQrCmxr3ER0OS
YFMnT3q0uq0ltPg3WSOogI1uaaPn80pLjDy3RQ9N36nzFLB4aWcCvk3ZU6+XKcBZ
jkwlvu5yIu4SpZCIeRfJ85sXuvOTYRqdZXIg0XyWKkuw2ioLVRVHdY0uJ5jutn2R
Wmd9MUzANuk/VLyVDcwcpfaKWKUBWHH9xZBHONaFIJm7eapJIPumeGd9j1Ing7DD
9DpeNw5T/vw9crG3pl/8dthoiIdrcMPOeZoTkNdEkNT/ztpA3F4c27nw9S/r+id/
2QRIyrfW8L5FPzvdn30iTEaPR7R5rCADqXoKCyVoB+YatLvCLel73BJZdwGg273j
Th9qbREzDmCvu3ILYIW+kAsCpG48wfz3MKIF6XCpxCEVbbFQdbOKZi1Yzo1acbxS
gasXoAVl6uF3ycuQakt6nQtYpQgtBKhQGUCxoQih1qNFPziJ3UyoPjEK2NN3Xv8n
vnxsIVQ382nVNecxelCEnOgrvNQ/iZkqWbEXmE4c3Mt8ssUCr1dmSwyKLtyal2HA
HMtfjZ+6UKtXS0MssOxs7MeoYKQplyUPkfUQX8B7M9bEHMr/uaelNp0BzAIeytHf
wsvHKlwa2o5W7lo6YV4CmELm6VToDscB0eTyMmep00hCYqb08CO8vdgI9iR/vEN7
3vL14FSMKwYzqOG6vRRjd6Wv/yVR100dM+pr7hAybavCiekxtObBDgejwfKAGHLO
pvTpUP5w01WKU6b+w5G8Y1B87TdJgP+41ewLMNKIf5bIEK4I+0/pXyQX68VQolVj
lk065p2Bdml687lDy+shYAUCY47WwWT9RHGWhgq7sbrj5/oCI35pKp7oPZ4DCSjR
NJb5FwFwBUhTRh9o1nicp1T0PXs/AEAqaVQG0hU84lY0o6RTnIDyZT3hQ9nP7Ekm
Ze8BHtUXfxIQESFcT0bgV1nOUDyDJOObQuEA9T2VNwI=
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BUYFKmoXOugT/rCKrKW+aD9ZxbRyABebcZt9KuZAUbxeQI1gDyKg0typOlvcMwJC
f+kA8Oy0I4iPZY5bB22IdLPWwx3z4cquui8MWaGRODVLAWYAuPxhWv0nU314Oahs
c+de21/1hYmJ+ZM9LDsdFTZ9qJomSX/gVTE32XjdYBL345JDPdnlke/dy3arFsId
aY2yIxYNfXcwJ532W6okBJKzmfA5UHQ1R4xsYLqPIHosP4Hhv4qjctCiGJKVPQPz
MFLWLDxZdX0T/69FDYYlcEZ/xCk7tWRt3I/QXLLr9cH2YXG+jhG8JWikWIVpXW3s
M/rVUf2a/uZz2Njfm4HWTw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 752 )
`pragma protect data_block
a/fYe+3Y50MIvyC63wIYccDSzE5DP2JWcV5MnozbjiLhJsqoRu7Y8k+PlptjDGQe
Qke5FqAdWUtDjFKw4jHJupeJ5VWbrBKKccB9AYJl73Uft39myq6W1ZbE8hnUpXAO
dKR1Wrvd6vxGNgZXzBUZyJt6gUo+BE4EqfWJPoj1Cnq2pWsdW0vyC532j0ToblGI
5p+bmsANflmYEVbawFXk3j7mR8WDu62Vx/exFv0ZHLP/KfztVqnFqpFK5FGp0L6S
oL1Nej6mhogsuZa8rph2HvhJWzGeC6O2JZwCnGE8xjFHVnu5HtmY6PuMKorAbycw
S2jbvnHn7n7Wde1Q8cWgSftojkzg1f0UkEqlOfVv+y1kOos3eS4fdqroLehBErE8
NXav+Bxia03a8+m43w8JcNrJImFwAyBvpDLq7Qsl5RaK7v00XqCm3DMsE/prf2E4
pEXpRAiwQT9W8UGmQDhd/BmQUOFdwy5gezHgfWbgDK/LC0px5iJowWFUq5K358+M
2nEcmhLkhuSQ88u2v7wa8MQaseM1deIdms5XmcMsdwRBPqD7/BNeSchpXVtL3ZTI
RQayX6vMigqaqW1neufjwes6WN/jQW2Q1W4/r2Ru2tFICavOeo+T8DXwxumDUJRo
cCj4AiAD7IC0YyFyjJctR2TstWQKi84EX4aAy4RHMXcgh3WeqhUzVooF7MQcKfD9
Emd8+/d08VQJoTwViEFTJR2q6tZLYNkMWi2e2iQEk+YdvtKcgq2oiF2ZsYzOGD6V
jK14OxQPaaR+V1EN5UhHhzFFMx3S0jfvn5MfcYd4Aegb/8cunUjEYyPf2vf0VMgC
cUmRO/8/J7FgJ1JHkyLH7WQOWF6r1rAIcx1lmOMPSrofFxOgNxTB34h0mFxUv6fQ
cGJjoe8txVyPLZD4iwIi+ZIvgeFWHhBn7WQTF2pfafj3rE/lOpaIwk1mtE8SIgAr
rU2zqMjjbf4Eaffx0S5N/BwjYjcr9jnVWCef79xvCZQ=
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ceAuXH4LUuJqtquMv6Jhru/xHZ8OuH4f+0BoPSpNAR1NGDnvdM5pN1nVDf89m2YU
jyBIWxg4gvmJlDVELNa8scK+SwNs26SpM6aurcKfjkbePmebijdxx2gqr8EImdvi
xzFjg2EcZNt73Y2HUjfvfUNrzcdfSLn+LRd45ZmhKDh43CDtNRJiNg1Bi1aMnlHe
4t1qKFNA8kG0v/5OvnXEVGXYjbZqS60Kqctzo4SnR/hcNKqFwVTo09WFe7EhwgB8
JCNaZ2qJc5v82zYk7h8DQ8tP7geVXQ0M/RoZUrmapglcdS/PXqzTpfNi/SQLjgfD
n/5Z/lNqsjPXSZCqrx73PQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 624 )
`pragma protect data_block
XRTJiQA8snVEAc8zOobMyF0nXFk7SJE3s3CvHuVu5GcmAIHf1T7IjEi1erJ1hMNa
J7KY5X7C3Q4QRIsT92Dsek98PeqjB/E/I+Ja4VobddwpaCJSy7pAlb38cHA3w+MY
CtqiAIkS3xKO9bpD8AoRfwDDnIXz6JpBSTTJNTmpGn7//wg45wauRbk4Ia2nKYuQ
yNH/OwwHrhLY+VRVMN159ZLVkuYXgTsGcI6sIXrfxyLGUd8Sk5jbUqYYYcTBwBKK
l2LRiLnm6vQJS8r4DeFXve3rSJlPfZbZPGhFf+jPVMaJcEht4qmw/elXCRy3/QV4
RNxs5z49GHkqPedjITtPlswiOzn+rpWeeDIi/+s1s7KFmKadjhYNr7QDdmIukniz
JS6rgVaaWkLetce+OoHKmLozEsDkRlcuTSwlJuWeFFpz2NMOkmTgGVM0Ky5SHO98
I0Z21NDs4HdvB9NWvZd9UX0DuiWm/YYmxgVoAhut7kNyJtZ3bnKcoUrTiE5mZ3I+
58tCAe1TtZCo1sX4h28yua7CR1xcQS9vYd8EBlpktQd31MiI+N5pIqzfHCgIq6Hg
Cqc2ORb4t+aEFtEYQomIx5n+rKIYpeJupdHqJazc3QgkwKJJaQWwR+0uRv48p6IJ
6LTZm8bNhvR7CU+Cl9Av5uYeXato2PUoj77uz5iVXmxg+T/z9WckGpK3cLcwSJWP
aObnbYSgv3E4RLuyQr+IoX3K7rdgDuXW6GO6tTBFkva29FckvoUEwjR+3Hf/JJeq
NZwtBQRiKgEdocBlvd8cosMmsZPS0IjCAsw1ezeWrIxd67qmJIImd3loHBkbzQbx
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VeuJuZUSpWjZ8en4TtZaqy1e4K+Qg6eYCtvQ53vqd+UxA/A/kdApZ9zxZWv1DAPb
iQT+bcrGbb/QIVsoaiSx/CrAteDVyEbMsIX+L03qjj8QuDMD4zVGn30tOCYfMTNp
JrBbLUdrbson+V6bEMxHZ+W1ADVX+vC7slXDGIfUuXWQUIxVUlEDa++1uv/JdiAt
eWkgraJfnDejTPSf6E+Q18Kug6hR/l3QO7a0p9F3exQnBxZnQvJokc06i/52djJP
Wx+xwygsBeVQtGOBX7i3nArg0IKVsOZd9L6QeHV78bxyvpXFnATp9BcZWb5GV52s
xcbF4dXCZ5r3o2wdMcZiZw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2592 )
`pragma protect data_block
GVO314/Rigu9JdkOPfn40Ygf2EGSEOmt6Y3n3+5LEVX3424ZoDHCx4uVRYN0MpE0
KZAl5nNzrvZD5cGldJjxX89gJST58M+89GGKQfABdoBL547W3B3YnL8cDco4FHOw
0cgWyStEOE23u3R8t+9z2QIC1jhZuJ3HNsMwK4gdryc9SJ0uELhH0eP7P6AhgdBn
2vpu4wYKh01y7UmzZZ2kZ4aVXVgCBO2KOov72BEwOxcLpP0x+u//e0o+XLahlYqO
OqXJI8jztaBGfiZKIPnN4yCPVhHgM7lmCYPTmFPlqW7W6EHA0YhMzbj1zFQQ3oGI
Erw2sDOoWtQQXbnB6Qspv5R+o6IdTwQ1lF4veeKhPdj5JSNeWur+xrwabpuqCNFs
s1jJBt56jchCp9QtSdYc6dzz6MV4VRKU0tjnmB4qd1mzsAOqBZhIbN5XOQ+1p7Ag
Jcv/O9bCgKixEuy5P1Flnas5jIaxvYQCFfIIdz8FhC1IMSDYZA+awbRwz+OyZad5
Xqu3YSYv/TJre5OURMcZHmq3hruIbgYMXpfqZq3h5jCVgD+dmwwx8MjSPO0qZs15
U2o7XKkX4oRGTRSE5+ySj1S3R7g09goEgeKo6GZHqjw9Gi9tgRc0uEzo8qixCFPw
3eqjFuJhe+8hbMznpneZkL989cTZO+bmaWLTaFMS91uexgkFJYaKHchlJLl+KCQs
1dXcnbF4TVwEejDXev51DtvhEZl7CEqO4QetLuzJI4JToiUfQ3iLSS9APiyQLGVY
0RICdhkjmRoT2hoIyVmpRqsWSWvsHg9YNGrzl5odZeHPJ41w58WwDLkw55lDA4Ii
VxMc9cXfxzsCc5r9ZohZMqVuEPVKUxxqnskxVX1170PGu6gY1cghMKrR8YXcBKTb
LjOPgWTE5J/6xwRj8lJiADwHcrPsdf/yEoCOzHvecAvwkvWxZnC42Hny1YlaTA3F
jbn4orcZVOY60hkiXR2InibXJJukDX1Iv2Uu+HwWAPU5My233HHpCGhS2mPmfZEo
fNdpLJ0z27pdAzgzcjIMrLEQDb0swDZJNQqg8hUcxMr2cFOgqKozMVjITBwVu6s7
dAT89CE+1gQiHvJbrky7gZxmEToXJslXfnURj5C/5RvFgZbkxSItku0YpmkYD2XQ
PQYYqhZ4E7VVZcoE4kKQY/Ks+RRJ4GK+AnGsSl6sftlwSsuMYC093fyrqUdqLGND
+5Svy2RyXt4e+njCbYESr5WZz7uxiEesEu+P87pbua8i0dKpBIcsXMOvCxIe92yf
K3AZbcM+vNogjNnZsF5mNKImIZTmePmX+5qGlOpi1kDR48CG7WyFlolsFoHHm+rg
j9c5rHIqYoz8a+xj7WFvnUFysqTu7DH17fE0l6dDYMuk9+SAfm7IYtVF03QH//fW
T/ge54xMluEzR9jb6F0s7EhFJ7N/Hf/gVyP3+vNO5jlqv+bSXDSmMtQ9ak5ZJP+M
N5/XLqeczWw4UqFFerREd9x8PbpOgzrxXO+GnA+QQznZEis8hyglqUCvb+P9jBTR
zKtqmCeFV2xEgIT+pUtFX8F64miKv88lpZfNRngkXTUks4tEnB7MtM/fXyqxWsvt
1NXi+IqT9PbV2heDqrhtzfaoSls+UA4j3gxqhN17NawoWyZ7Wy/WVBG9KJLO1DHj
LO0rLtHwAbrADMuRcuL2Ewt39i8F4iLvA6TzkscVtUZU1BEqSCZuL+xscaCxrJGV
GVev6QKpKTY1CN3yBuUNokG05TTyq8Rz9kJ6XPmO0WqoP3yIW4drU3oHJiGxPmbw
aI6WQrN4rbUr3bYLGZLps/N6t4KU+pqhk5PElAUc/ilnuCUS3IvxwBPSBt9r5rRZ
+pYE3be6pwburhcgav1G00LvDLBxgaQoQwO92XWZOMqiLg+4t6Y1kd7yoztEy8XR
+ziTrP7I2FwKgz7ISb8TNKfSCzz+i5SgL84p1RKpEqb2X+uMsTqCnc4FfYTl4CG0
ib60I0zgyKlcHT0gfdIpOWZ+dDIkYpPXawTPrCsQWT7miKFkz7k4SRpaBMyQUet7
DtzTaKn594IMsgUvaD676DdaSAh9MmNkvIyv968I2GeIAp8oJWXzQL44l7uAg6qm
H8sbKO0hRTdXgk6Wk+JOyMPcgom0YPZ8mS4hVh+AR5DjOMFPcv+DdZsdYAucHMWM
Oov0QfciMOokYNhsxWRzpAIdZJpbLATuinelk0P2j12kJjwq63S8s6Kw5gt7xKHs
uScm/1kVYr7iwQP8dmJhv6nS+fCXYe7qxw8JRi4iGtuNi+T2sb+w817cHIi1Zskm
wYlmG2Pkx8gNi5LiDPxb3FRXpd42tY/QMr7C8pWLQYpXIFCSNhIybwTfYnK1qApa
I+DR7tXIM4mL6SG/aBbsIA5hS4IUOf2jdChLvVeWxcig8yQCEBNylOIJ97H7DkNI
WhhQAR33qb5RmeUfOZh16KIXPqd0ufZisnnLjHxpOo07MdQJ1lRhEMRDhQW5TxuD
RoM/62qd8yxpJmnCdlVFepn7WSHUCTnDmhXPELBQfIJPcKcuHM7RVL+gwzIfgRHF
T/3eYP8hu+GTXGSd3UBGdqyUIpVOb+WeUbOyCtjo2wI0syBKSA3mRtcDNwbj+TtB
/VHYElpXMfPs2HYl3wYIIJPIK6r/Zlx7hXAin6bD2S8ibmAlaHKckWcVidmg8X7F
6JE0nhTfurNWH+P7saL6A/uxr5LWVM9jZfUd/89TO0a0Lt5P97p+vuTGv+aUC2Hx
oBux4HQNzlTm52YcVqSVodigYe2t71YliTNhc36Tp1w2uWer+VMJ8FIZxQe/rqPp
gCvONi9pMOY/2b5TW1VANJ/viP0kMvcfMYoxqvxmtoX9WbvnXX0xdGw/HcKI80RR
18gSiv45nGRyQl/7wphtvCyDTk1tEOsYG+95p8iujFXfINqsUPb2KcqUqdBaW6zA
bqSQzNV7fxvejlYIEKzFkgPLL/2ulaEPwptDJEgjDP+XsnPnbOBsYd9jr0waBd4L
2wliTTugdpBScs+05PQOs/p5LDSqINIdGY5m21ggmzvJe0zfTnds5TLouvjz6Xcd
I61FB9JV1WHIeyrrZtO5wUfMtoBYsBNvInwMXJ8hcsHa/XEvi8LXmFOvKMI6SAyJ
AKokWasfZKrihU1vlYVofBjNJrbQw7HLi91pQl7PdkqJ0/q8SUdiSQYc9oGC2kd7
Xzl8of8eGlo7ErWfQnkUo9Al5goel+B05oFnsVNV9dnicAokOHz/HXWPg20BINjY
TSyXcvkQvZc3Y4ASZNyfyyrWfylujKudNqsmSx2DCvkgfsBuLxh5tv6MqLzWdHG2
6z4lQdwUmuecUXDvUf5binN5BPPmX7nfqz2WzKQV4HqED1oho0ul3fyD/16XCSso
UFZpHg0de8p1HwPyPkKufbFsNZVmzKyHlrwFrVmuIrgQS8lzmcvwTwaGSow1HsNV
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
oJgV7+82mBgnjhTlaa8Y4sOjkZxjPkcyZPQFkaUC3g4Q3G/iKO4jY4K9H5zg8seM
TrLHOXdNWMEm9u/py8veoxd2v+RBz1gkoAHA0OBKeff2kAJmiLGC3UGjD/fyd7fF
/5I38KlnLGA2de6J4FtMTM0eYjG3EhyBUd5hCz1pMmFm0ttLF0loPBL/D0esn4P1
JWAuUNFB+nN73YpwpPz5/GCYRTbLx/S7jRA3cVsLIhRglp5fBSwGOT1DgxZP9ycT
fdVomH2gdSbqp12stK5fhgnMPTCdc9wV+uudWV74pE/jxdWSAOs56IqCCsz6yF9g
CM8xaJtujgZTY0IkEEuSFA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
Kk3FLTUmZJrM4hdNiQT9IGjr7ap9jctt843KKcKoqE82CZQeauAwF/nOw2c8wBLR
nCqoKpfwMvLnKOtT1cd9fDnJ1NH7BEMkP7Ulvb2FSqxJYoOqjA0OVA/Yig8wt5aM
/YjmPMA9C4Xu7cEvefzzce4K7rIMI2L/lRaHdLpgvRe19ALbgsR3bBgCQkh+pqSK
P0Job6L4QkbNubGGW8udZyyquY9RilBAPNpwAtc4w44nAfbZhzOliYta6Ffxxb6S
4SbQOO5qwJy0gJhPfVOIbTkI3TR++F54jVPNBpWwQ2CQejo368PCuHZWAud5Z5JJ
rsbS6IEpPhZUAaDknnjAIfNxJHtshUYL/i0PYt2sVRhYKFEfACMLWuiQzXV45NtR
bTDiqQYjB7P1zujIREtUPjjIWYcRG/5qT9Ye3ZiEc0t4iXpO3LXX7ovWLZjJfNlT
xvKL0PVZIWEIetEk8GhEoPoFOKYSa9NF7I2UVihzpkWeGlCn0EQXuz3CsgcSISd8
AutrcaZg3/2722dss+IAIuuZsKNWHbg7XsK3JZkEvb+u1RXOGgBgrNg3N9dNN97o
iE3CjWgL7us4D6YNlVHPuJA0UwejQCg2xXVEbw3QV48GZi/EoBItezVxv/O9YWQg
j8AObsSbX+blPscRm3NVIRdUM188ALxwx+JfaAJgKBeUfcbzsHzaMEw/qLtCXGJx
x99aFUly1hjPs25OdxUYqDIPouXxqr07wE7ZpqB/9fLyvqnYVBUV64bjzbKXew59
Xq4vEWQVhlFmA/lf5M3oZ7beoQQaw5Yu6bXXvV5fjFjTejYorzuP1Rq+UGDwYCTE
1vKbPkxAnsKJL/Al9x06FqYKW1J93lqMY1Y1HRQ5ypqegJpFBuru30u8fh+3JUtm
Z1qaLpue1ALCOzV+cBSYm6v1/Qjhv2Bnju/XoYeuIxLVIJYHYslBg6E/Vh3f5IJD
oNl90ZxCFx0+jQ00+DpzVkCq9zb3DFW8IJV4O5BwXcVppxjJbsSZsbEFm4qz45j4
acCacGDcqKQI2efIc9510WL+JwXIzc0n3U9jMDNyzCuMdKf7cI7h7lIAU+c9i5vF
Q6IgdRkn2hoPMZwnC065KOok4pdAHit7q1dR+U0jHx2cUpcSLIVn6vBREYZN1PQd
xNouqJ+IbEBla7l+VlMgK/OvhvvM8DiaZiItjBUM4yq6zIkPyEFX8IwL1v0pthDi
pu69u3jdntDFI5e36nIPv/asF6IxVPK7tMyfcLvQ/b39a9IRQLmlaP01IwTJyl72
ihNEUUPRCvtX8O1mgwvdErEMLWiC95Vn9ZTx+HBUs2CoSsQDPAlrdL48+M2b7Je2
5+mvZ5qbRIwJv4q4IvxgXd/XH83T4QRnuW6k9B5KULBvOWxUa6veRhf4c+aNyTtj
fMIG/5zMr/ReEe//KBkQucBDlJ/NdahV1bMWVFMV+0mVIYlXuFdBa55SMRmt9fXB
pOeq0BArrAEoIdMNKd70KAQolxCx/CUJPVYbRhE8iWnVFBZtGTLk7jc8LRo8KT9x
kxsf0PBuQaiJZcomww4CoNaz7mCGrR/p+rr89DBd6kVmIss5jOO08Q8y+9+JeWCw
8iwRa/wWva3K0uSsN/dePVs+WyKjtSOK5Z6day8PJm91Eg9u9bIwdyQR9XMhR20Y
tRHRZsAdFpKr07AKzhH06fvRvbyUXseHlrXswrvGoMBEUVBKoAekb5rEfHZfKS1s
T9y8nSTflW65ebAk92r6yLqw2U6r9XakdH1dRFOTs/pgbWTkhc4GXL+6r6UGEBjM
QC9Mjjpcb9YXDfDtGzLuRAhbw47OS1cyBOCJxT9z/1IC6iJLxcjEwG6cik7o0pMK
nrqjeqnOQF+4O2xmyA6XBD/JSWHV6l7xJsa9qouEJ/AL6XwRDudq2qW30+5u+M4n
aVvsSK2I4X7qKdxex7NCs2WD+kc6o2Hnjr0t/7BVW2hxD5IgxCn2DxO+mKOI+pPA
/R/KIisYhK9pYDViNIoquncuOz1VwjrbJhNQeU+slkymoOw/s/9qw3DEwbzJ9lZP
yppe+NnF5UhlAntTymTLrKC9zy9EfFMZQ7KIBgJ6HqoELe4lhRFiLILLiQRcrlEc
t/yPktcfrImRcbzCjrOaFcWBT2MdSrfDzQ90uRzhr23ZIeYMZD8TEUTYjHaY6oo8
+FIEF4ASyXzuIaOl1TO6M/lCKoWNJv5TWhy0PuwtTI2b1T5/tIXOHsXo91qMMdZ+
hvRVFujELht1Q6ly/m53kh/HDahsjWyzekA89ejA6qU696/LgvfLB6lMUWtrzgGi
v8oNPNcBmz6EHEAag/DfcNW0VUlzuK/g17f88vvyDiL/uhGCBg3UzYAZ2b/k8Nzb
A3R+I8AysnikoWmOTnG4AUibAYazbghU5vTm08QQzu4MGTKUUs6ranqCDefdgQL8
AkqOpdNhTck02TcrtY66/w6LpNLw4fdxlroMAk053I6rp9wNC5SbT26Saq39R9oe
9sM9F0JMlL7+vj1OMFnTMuxXCv/VRZ317uN1tPFyNs6ypKvwl4UASRFkztbRvstS
OAfaz1eKYOIEmwhKVHub+csyFhWRmhr9BLcfz+64AD7+6GTl5N6JnHz/COOXmFiu
GWXH7uQ1+shbz+cI5DIEurx/psb3vTnyCretVn376jvqNwNUirTkqHLvXP4jxMGJ
G4LatlmjSTc336lE6nMIHhcvH/2d0yKgWA3+SuFtoz1fBh0RPtLUfJC45dznNQ9A
RhDAXWnmU9aWmgcI/Mv9e8L2kEbANzTMFYOOoJeIytP7qJsEvfyFbjlGTWCjlsbi
RR50bMjbUqR+OIVG2tj5vNY41NK9ut6IJIrSKKnmuz6zm63bYFat+sqX93UYOpx2
kNQ2xsBjxuCB/xabQcW7f9H70tFljJMe59RDIyxzH9PIQJNIHM56XRJdUXEwDiKL
j/FMCwU8pPq9DbaNUIIRFYqr5hcZpYV5vKkforKyYnZFqFfTXN7yLCo3HtZ4BCM6
/oXkB2kI3s9ctnHKdrNP4l5qAAULHGGTRVug+iA2bN/q52nhTQ/TwCFmjABiPr11
xbs0c57kY/Xk+4Scdm9bBqNf/oK+pCbFog5K5bEDNCYDedhk0SU08wV5AtMBgrfl
zqtZSv4ZAQSzgXqXjLVXGIXaWuOr+4zQxnC/To+27YP+7mQgqh5/SnMAr80nHzdB
zTSMwoeK050KaVjHRXe73wegqksjzVNicDVhVaIyJOpOjlheVGH8t4j0DsCLtFeO
Fr6NoFUITX6c3nzxEECYpXsOEG/KK9oi3l4gQre841PtCfiahotOGpwqSI2QnQy+
KCRN3WRLf0QYyG5ybQyBSIXmtvsMf8Ch7+GJtFH2tQI0eQQKI6rUu/9LZIWuWXau
TLMCVSo1B/gZgH57XZiyoat7x4jWvE0YjZMYFwJFHG0t0j6xiqXpcho2A/xrLBFl
9bVLdVGTrt+w94ohL7/uEYyOkW3g2LCT/RVdGPGnv3v6TBznO2GWDeLRc2rohrQG
7JP8WLUPABYaDuyTZQL13ufu/ueBw/tQJnF0i764kT5FxuwNl5mcDdKEee4qCOy3
8+4PyLhj/M9pCQxrwrzTyepiK8n+Jihp3nCm0hBan/DSeevH8isolfoUCud61iUh
A4iW1hiUc4OEaJiGD1xlVtRNtOH9hYuHKWKUPsi4CFvNkj42TN0cWcu9pXLfRQhd
cht21sY+GAiWPrjnnddyI/rXe6pmKRmMfuZjxfwgOLiX/VilotwjmuVEUSBapkXA
A1OaDrMgReUoIfTbvgAeDjLY6ZwWMGM/0lY5a6mVRkAUxa7IjV+a2DGowK52SB2j
ep3FEod7Qo1p00LMChdtwhmqUReGr0Jwa4iJ9ovyPXvPmw3/tZvtJCxrn/eMhwk3
jiDFfs95PUTqe9WOQbJtMw2AZ2OeKDQ3CFfMhRrnzRdjf+ndhOplJeabqcxDw3CY
uDJ3xKzfqUobTgRFNdQ5cidHxBlKIwAToFnH3FAG+oBttgdTfgQAJoc+h8Eou1pL
bGE3ahkVVCDldH70fNQp1B6PgmK3KqTHR50AROlyLS/h49GO1cWLOYTT9MAlCeYj
96fKhMZ5Yk/MxvrEInZL6lwy/1DZYycT0T3w0xpaD0KWK/zobxnYr3f4nQjmxXfe
C7TbtlMuE4cWQb6Ckub4sJNxdoeVJzC3saJzh8r5gojle8kJaADvr24+WjhA4LvQ
CA6yzZ8Ob3F7NIUhHlc7I9X2bwg9irNLAVGb7WOgeGikTBnDBqzv/pecu5xZwJ+7
rLI/L17ty1TV5WgV1Z4i5FrWNSwa0c3dxljicy65ANC81tPS33FRy0VZQKmqWesL
6pqi7rrsOvMtebNNY9fPRkfA3E7paNIsXYq78TcqjYva4CFV8ULiZKWY+FtLwJI1
yFfNS4KykIute+IKFmdP10IJrChAY/cAFvEO21xWES8LpKvv1xN7FOybbkCw3Ict
ZJolyuf6Y568w8n1PegwQEbbFHqw6VznNDh0o5X4NwHOfSk++hNhvUfe5MzMVGiB
DgAmG82GZ8VI+XtZRxZ76yfT6qjWxgMBP4O4CdBNM/fCb+jvOC8ocUdd4O+pFoZ1
gzVC60FvBGF7qTOJRzo17zNSnPEwcKnIie+QoE00Euku0MGcpzEaixiFkDoup4gi
WjibuXXVZlH7aZtbJg8qPgzex2gTxhHod9+583I8zKDHTuktqEkJ0QqgyRFCFMZ4
MFzX+4YtyBz7a4AjuJV0kzNN/9Mh/rYhYeL8kSG3n8LCO+j8UyB2oDrtX1ZtbJqD
uOynJidQpuZBJol9HLhzobJxF9qBCPLASf2Hk/INXXkNlmEDVbzIKNf3aaMEL0wV
wZ4peKEkjRrfStCoKhCoGgjKPeBg5ZRHeGZbE+30waoRcAvArjnUaPllwyGuPatq
dS8vghGBK6/7R/P2VSKxiVwzERvspuB8ewke/aN4nPdRO5VxSDfy1/fkz3nyS3ka
LNeILQuAOLjx12UYfJQ9fSvuqnNzewzwFj7F0FBL/K8j9MxAoSuDZkq0epaqyvvI
Jueokgm6TF7KzAZG9fuycSG9vnkWQBuu3DXRaTpSksX3t1kc9LpyESr1XTH6vuVo
oOvWwboaaUr1Vq2gIDEQdPULcYqdPd4oD/2gu0HfLZ151GiJr/W4gxzLZ5l2MhAi
6LoDcxvsO5LAd5hPYinn1LLt6G+6H1LFt/JFrIuHwGEtsCLuAzFPh6F5HwjaTn4Q
P+Dsn42EHj8rbe3Vh2Z8QX0ykdhcPqvoSwbHiiTnwBZ6NTYJqwYe63FNGdTXig4i
7jrRn9sEqeHFBfJwsluyjCoFx+1q9Oy9Qljvltze7L52UpaJ4smLBWmo9mSvjQIH
RJPoMvPmCd7q5g61LTaxeJeIjV/MMp0qX7vXOdY+W+N52xmjUzr2HNe4YfQl9MUm
0RFXNHLIFTTkAjsOYQONU1yNLszFa/4Cq6VIvvqYgsAVAWXqHA+eYJaGGyfp7PG8
IFDVQYIwgJBptYLe+N4onOg1r1KDI19qU1c+cDH7YbDxW1sspBwbaQVd7os99DDM
Yla6BoSnHD+fw3e3CwUIHyu3GtS0RdO0Sabjd9xaw/85oCLvVMuMWCzdOQnWwVcz
Uby/oH/6r3Gxb68sw2+SvcJI0QPiMQwo9cidsgpn9UUSatBbJyGEbnz4wXMxyz0m
2SDT2wmV0xtuMlCfBs3oyHQ3SocYWaTsPCldLlb8IKJqVQUlkENiIGG7XgLGOgGN
UDTMdwMBiAnuhkcBA1NPPFeUbgso1qQGq1QaaoS87LPgVl2DRtfATwTQ0xVomMiU
x+ZrtTxVN9mAiW7MJGgxrJLkJN5+JQ8fP2kixVp1Naske7LpB3oMpLHUy+fE63EH
704Sozd45pyoCTy4TImT372HE023FzvIroCqWuf0sFy5nMCnQwiqcvOZi63Codvt
vHXQIEyxfeGz7gyIGPkiJgtHyI2qxepbL5JbyU8N1q+1R4otlzv3sBpgTBmG6589
BYKTz95Wf64Fi80a/ViE7+kklmXlMcmIH0WuBJhTJ5isQRyeiOGpfNFvIJx9DQvG
gs/XbknxFoTWBgke6wgDzTuTH2kzx7HTB+uSNCUL2YBvpsIjECYoP+njU5fmQzD3
Ew+f6ftGzpIdStEVyO2Wa2wFFj4ltLV2+qrX3CPM/jtNXTcFgcx7LWqNuhUYb+tI
bIKrEjdTTPo/B20TI1xUWYG7wRwFfZoUac6nqiJ0F53VgLQSrvFwpibMZ/m+XJD/
+INyTsvL9cjcHVZ6x0G+l+ZHd4GVrGKqZRAjfP0LYVxR0GpiBk9AeIphCUX6OjH6
NBmR0rbTdHzurxWPZpEo/yb5eSrY9VCZSCC3sGJ0cUxobOEkyZoZpCfvSbz6QKjS
yPlHKTJCmgltbAix01fb3HIUjgx0c3mkxhmkPkoZIRO9gWL8CT0K8Rk9Gh6f+i+n
chk4Uk5YA+MU/bzhqBwOWEpteQN0B62DJUpcz1ftsAlQNi1bLcrr7ftlXb6omrjA
f4KYcnkdXX0qdwD3oa8sNqQa6Q49qciPCyYsZ9wt20k45rDex1QYQ4Qq2Bwh7q1y
zwm88dWtsXaCAmV3ai3zSWYfx0jIv1RZ1gOrVaGeZB6TC/Zk9ceJLLFMqHPsDEuN
NQ2wdhk4/wlqXJG6mdeFJP7hkMNuzIKpm9SDcOQ8Ov7ff40Xej2qd/2qoclDxAGE
kVeHzIazhJ3eJiZ2kxY2H0WgJ+F+sfpY2ODT6vgnL2vpTdUgRkMP6aarMx1IKXEI
qtRTwCmH2RDvhB/uRykFThgQJW58tqx1XxzltjKoKCN0QiDMiOdR03umBVexLt7/
Q+4kJ42e/R4pHLiOyyHZV/tPyHqNIUHV/jUHSjhDONR9skirKREouOgF1Qq4R5AT
HWMbB+FCajW2eUy9+EcVaiMaJtBJMw2dS7S9EBKU6d7wBKCcaBKntbUuUxSRTt8i
b2CtMMerss93R7v/ggOmQDTT0CNgQQtsC+CsIntkJ+9JZBhvmXJQQOCOweqCDrul
PxFjWo5YfpowtCISkP+PsNmOpCstkDPUCB1AQjH73XOOd1A4OzYH5gE0yyGrA5Nl
BaLWqrgSKIAj8fUBIrpjRrxlPI1y6lwXjVLHDWpxD0GgWdNSkfRm2vS8f20hDt/l
m6Pvk5N1msXkD5wKC11wkx6L2rkRNcfX7uPhavxRIEGouly2KDc7BtO+eEATpKSb
bC90K6EyaAX8EfnLW40/voEJG1gH0ksC0l5TtuFM5873kv8PgGtYeLScPJdFtioM
cEf/uGlhcfFV8x+sovACmuAjKDKeD6mfWg+YpIt/xvJCeACV7dQ+xU41+2Lul2nK
FOglB0RSeSfCcMTjt88IUbqoxUqo6OmdiKZHxnx6TSjhmMQMFxoUagTjypl98roq
gGAYMbNnxXO2xeUP4U4cOtRy4pmUZMkM/D14fqsDnjB2OOPV/EGa0N//9WfbXYb8
LrP1AtqF7FLJZuOPKEKTFxd8hf4xjPG9Wg+CIYL8bDYs6/L9xYu1l4BpTl7fValX
TZRgVkIshUxSRJpoiLMzlV9KeBl0KIwLYyGLE1TNs1w91CImeQQN1cutiC37J/1m
hcRsoceNNZ1q7dqq7PrfXs7RIhxuuwW1xo34MVEM5fmOyFb1oZRC0QiHXvNvKXmu
auNtY53Bi2X7OSdhjUm8SBmfO9b2fgL45FTLXRwTdLfFKHAWQt7pQS306ZsMUDbV
aL/wwfhf2HghBHCABIl9ULTlUBota2OdUNgJph8AF0GPOJPKwJ2mEu7KCifN0vAH
S1jUS3F4GoB8j2fdcA9KzfZHHMpJeSGFGnXfLQ97fO3V7XDFkB3LQYWUHXu3e9w+
vUuLXJccoK1WjPA6riaaGkboHWSrIactPAO/cmVWiqfXCCTTiKPWRY0kY2+4CPzy
xPphjd3Uyy1LF9gNUrxXaHD4GjqlQTa7a/i9NaIBKuyQ2pVb2vLo9+hxLbTGfQ7B
WsJXUvp++TFCNdS+Q6PKjkgXS1xJCwmKWCMsH84HB4mUubxA7i3ugxLCow/4x/DZ
1ekiumXjavQJhPcZuTkK1RLXBi2m/rs0s7hLvXxMRp3+nuWvqUqdEyf1eTm4kJKq
JyfQLGpgC0+H4z0p2gv7ByhKFbFLUV4rlB/rzdZSc0OMCDvDRL5752VL+HCkhSNP
PDUxpESksFoxrIcMl+0jO9KvAow6zzrogiAXDhgxFvsVlepGTM1gEMiGlDAhPATd
IgVhQoMLDk/sllVYmdIaD98NBqu4UkZUZlRFbSFrsfF7WwZIMGoUhYFLQnHHaTpb
s6WayqLExkga0zYRIDqC4sKffT3Cu0A7akHzocuQJObOZXxmypNr8MwnZ6Hzu7Jz
3Lkz7FLJCnWQQ4w5yWNVguuwjc16zybsqZXUA29oi5UQuaHJQAYIwWXpaQLspLb1
vW9cfXNvI4GhcoLUlbSwIIuOFcKyUmjhCnYZK3mzLMqlMQ6MGcyT9UyQGNtfDlv0
FFe2nYEev9Mm3l2BHKtf4GHrS7pp4vJOmZgshYWstnDk7+oQT+F4mLSwf8EOnwBR
t/MVSwM5M/vA6g95dMzRD/HnvvOh8LXfAEcI0dBb7QNvscYrqCQthTCQK+OlO98q
V51u2VNZ27nwBIAShyI27mYeceBXZSQ1nZkENeyaqyt/uBTfCGlX64+VRGhUeMot
RB5c579leEspbyLRhQF2LkRDEpR2Xkd5qGgOm6tHMoXfzkEvXTPmNiEAhIUphr2f
hmm+fjpGPBmSqCGOyje5jO0sWMPJrJ9oXDRWhdN/S47dr+QZ03RG0yvKAxejR91v
vC3LUWRd/SbhibXPbKM7D8MyKjNdKl5Y+8cbvtSH+8HpbzoHu0vv7qhesn2rbr3n
6d8+qS2+ILFFPI7csCQc1mTHTVVAfWFQsZ3v6YEz0d+zeO045UimgzCnrk7IGFeR
gYCyNZQKEshOdg7CWVDgrxjM3Ey7rw7MUxNE5a2iVeiCaH+EhOFP0H91GLUfGD68
ySJR8w5t2Lq/g1HMl/oFhCMDWAarUG1d3woNqO313grR/3gUK9IFrT5T/odspc4e
oEpfoUoJXHy+jbpE2XjAo4bGzovBsIH2iOol3EEa1fbLShKdkQEfzXIuKj3hqlyH
4HZr4LajrqgUQOmDzOH4z408F9LweAjpg0UoAGQH+sMODahBJ3QKS+eioEeB0kX/
2HF14B+F+WGrjyvVViyGGr6LLUBmNtLjLK277NebyyazaPSAucRjXlsifJgBn6o/
XRAkVzWQFITjeKBGRc8IwOmjUJic4XCTELsOaAvJznxxmB0wRZMHfclDprXwTe/+
W6dgBKDMhaH2gGnBOZ8+0DkbnLE5ovxqlENYiUH4jQe/GjaR1+H/zpK/Ur6/PPq/
ZqCjzK+E39ZdSGzMwMXqe7sDj/AWv8QuTDu4vrICIGpySrjSSLE6UvxY/CBO1VF5
7vwtu/oJhB6oCm5k8c/nG6f7xI5Hd/tdrWblPKSPrxLQUpjNLcjDJa4aqdkzoaC+
vh5Wmig2zFNt7FA4pbvGm29ajUn+jHw+V+sqT6K5mT0k5wbKi89Mq2iCJMOmtcte
mi7xzBj0rLDVKcNkDJBDlIlrgQpdQ2qYfizMHSp2VhNkMhMoKXOAZUcCovds6Tvi
kCKZ6CdsufWN5DAFXz2W/HBZHR/ASyuuFwevchaSPHWMJI7rv7+VTElQAMiyxx42
nCFBfiN9jP+Le1xe4Gw7c7+NBTDVRHZHLhC1vYB/+0usMaHJR6R/4l9QaXhUFV/t
gWh3T2QkEJ1AuG83TzpLrWWoyEzcubS1lzArTKGj+UbqQFbRpvnOgZdqmONB4AXj
hqaWjV9/yyqREyfLE1yQh+vhX/lFjJeMnmf1nPLOpMcP7mBz+Ro1pHQjt6XQIdy4
ooIk1Muul/69uWPitghQzc/84kPlfwA1EHajCCiMqu49sIxhQwNTUjWa6Kc5HELe
B0XvCU0k6fk5jpvJwR4719geB29YFumY4X59w1Um/AOmAE6oNepa48DdEXgRssgp
f0/428VKKnYAEFWNJgBYOUTo0Oz97oqDswNbuQdC1prDRFPeKmnu9Uezw7X1/UsY
cGoFNoc7lGoMdp26/b5Fiks6fIWvaBM9AqYXpBQBiISyF/EkT3VVboP17Hp5DO1J
fKwxJ7VekbHaVywbgivJDwNXy65WGr77KGoQGINcky+P70x0aRFIZIj/jpkTHlVG
+D1Uxx0Mu/Cbzflk3C/SDjCQERGVA8L+//G5+RGIRMDDvbDxLXFxrs1lFgGVfoqd
eEj1bdR4VzH4WOgqqV+aEG9CSYxXWoZBGFQ3V4vf7fcC9mfpmP7z6DE2jC3s22oL
uKLmCZqYo8HM5cFCYvn1KNdUTrexGpsRSMb8I9VMZHdxJbP3Xj3dlJp9mxEG8ySt
07wvubJmWuDA6LMgmOMsH95/GlTe9TF+Ydg09Dqhwjq7phjeV7uGHMOGTIQCfhOP
EMaZpyIhjr025L1k6g3TD1Wjyze4mKFHg0DpCrgz3ZkiJ5jfcc52RKcZdJ3xlI15
FNK9tfL4r6E0D5yfqZXjHT9Yn1/yXlhWmNVBdH4A+t0BNx1MmZu1kqXXCvtAPbJG
akAyvyYybI7TxOaKGhdrD22762B///JjkD6fFBXwKQaXsExFNvnDqhX65clrWwQn
NU9HMQlMz7cGwYYNYsOvA6ykFNgL5X2h6NiG0mDp5OA+BF4pL4UDe+tEiIlDiBb4
jVNb81Dg01eh/I58GZQkIXhtJgeL8YLiBmMvN+t5kiya2rjaBbjFgYV54BgjwrQO
uxfpoP18muQrZ0n8K9dljty0qnnK/frJ0FrTI6fYt3Z8KzJmO6fu23cDh8Mn+w9x
ZAj3rRXaUai/Xabv7W73C3yRfYAcciR9Ph34jS4vsSMI26aBgXxdbFsMBfdukqop
x0LausJiXALZhjfbWQR2kNBuWIXQBLsBZlqellKDGKkxgB9rsp9eZfBC0oSll+u7
6h2l/SghC3+EDbb+YmdCtpj14B9m4G3x1p3u+sdoRI2o4CIoB+ISHBAIeIEP7ovY
KapU3S6MA3QQHbIW0UJ5UU5pceQqdMzgrwC/NBTp5vHT1CNwNRAFbHbTuVRIzsAO
+FVjwu0t31Btf1spKlNfOnIc3RQqqFLvjCHV2NL1rS1dAQnHjG4FGz7d32/SWHsy
nFZXQtYNMZ8eEb7yav2A6Q==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UTSuumVgtnA6TOMeSeGLJwUpivxvTre7CZLrmwT1F52ZXqlW4zcyIwb/mPtq0SSJ
HLa4+Ke7aK76QEDhce38KXgUPZkWsajirperJDUOtNRRbXtwcbv1HkrWpNJGy9P+
HAVEy/k/cot1rHFC9eDK1Lz77oTtd9Eeu83qctlGJzAVnhScXODAzFtzsSk4HbxT
aw0yyVxJSmaFJT59dPOxqr5lxtMNZYBXIsmvV2/CsKH64ycQ8JfgiisQyZfWBbdp
47QUqr1shR2qrWuyg/ElKgpPyzMnF75AK/AkQw2VSfpRcl8v4ZUD7kofQV+B6qAm
Nq8tmd+B6x5dpWEmKHEpvw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2544 )
`pragma protect data_block
vW7DtYOCACKsGIZ7paay6fUC4Seq8u6wUZoLGH1Hk4ouF2dmNtEisO+b01ltVHLT
Choy5LhDJZiv2rtQ1Mn11COXVDRTCT0985Z/xWV5/V/hGl1gUt7kgWkJzoDMo7l/
r06eFUZmLwTELjlzfEVX5Mx0BXVDx+ZSTPobtX1KoSOvMlwmpOw8ihaMR0rtons1
Bu1FsJ0qAtr4VIobFpWX27DE8gxtt40xfFE4DvtrQaqZSacLJ94vi7BmWodgGcde
k9j0DH+IbBfpKVXFv4Df2vqAHrHMl0mnJbXsoNZFkHP7l9mLh2CJDooU2lbBMsTM
0LYYf38J6jj5yexEEwIZ8QdLhpuOVlgLE6PzDHXL+oR9GolPjZbxyYcVDoD8lwfU
5Ol2GTRXf9omxsYxbOyorB8yJqF60tURCozp5zFQ85cNOZ7ymGaGJBqZlUmEgqSa
hoigV8P1na3KprZs+cT2DG9pMckdmeZwjHMZwQAkgmunv6clVBLYzoFGAHJV+Ok/
9/Z+UM/ptcIx2c4NAOFqGvuYvdYFg3cKQtaeaBFzRuMN+TP/tJgN4/KJEqv+NV8w
EAew0q8Z60QAXOTYCmj0MEnMd1AgI6Zt62U4nvFIQTn2yAcrkR8X+ehGoJZsUoCW
/2IcPb9Pf239o+NG2fErQ80YnUt/8c5bzwrJcelM2fwgRnUTjEwEOybAPmOO0R4z
q/kUgO2RosAm9C0nPxMyi00mfltdSag6OgdlLxvPht0kltQ08A9WY0PTgV12EfqF
d9m2Tdw5SdHuVi77x0BNEeoi4v6pbUiowq1ZeyW9ebnsxc7cxq4dGvDu7uRJ67ia
NL821yt6c9JiEJd0m5b8DnAXYj0nSRwab7XIbVPDlDf1mVoF4FjO8/b3F8UT+eUD
uTtjogdw8p75T2D1POEIvEvZITUEefX/Oso/qq5Qdh+SkCBNxb72b41lrmbGBukn
A/biLgEnL6DC2Es5Mb0wO/P8QfCWC7m4g6jjqduxUb62QFQsGIk1F00ZgDtZmfGK
MaPrWniEQ0l3Awy3aCj+ExxqtLDdpFZlnOYZej5QWTeAqca+5boTLMV3ydR7Jn6s
Vm5znbO6lQ/KFpMAIDmU8U1xP0HFHIKmFh+0xzOFQAtMnfXLrV+x8vDUEETuVlmE
Xr1DLAkLvG/4li5/XfUsSAvbW+/LWbY9MGznVpTkbcdOp/LBOSGqHtw8DEoQlhFX
DTKm/WVOCkZDez3g2PNL0WAIQ7rMc+IWNrJwWrDCt+mH2/7sQKGZvVXMZLDG2vU6
8qQC2K2CER1ssFk1Z0OgE+7nZ+2ul276Q6bXsyQU+0+GpukVipQURxh65Feloehl
836tfR+QaQyeqG/1qYWpDU0dMED5Y71Qj92SHt2aoPmlOpJNrCTdpgZt0SEIoXxz
eDQN1uYSkrmTm5L158hufQ+Y8aotf7saYVl0u1QCP6dS2Jgm31DGXciu1qeDU1ug
z5d6Ey+l60fmtcs8UtQCldkryQLlfdO5HD+YUVxt2Z8Wi9q6nonc27Gbeko46lo8
5EpYP6CwdtU/58z/u/rhq00erZvX4tdGYjXNUbU2mgsPCEP0axNGiRnAbJneqePX
h1RrGnaR02Goa+AcZdmz8qvvvLK1b0duoX3g7RkB2MCEv/e1YPOmBqKGJG+H3s9w
0oTRggqTN6MisL0XtoCc7totuEB842HOgpR+CjNxXfLEQrP88T5TUTWJVbX70AZi
IvfenbrmEi61w1yvTJauRx3TiTHZkGe776a02LTlJ+qIF3wR5vBZbIT1Oe7IjSyi
w99+EC2K2UHeUfo/TKDarMZg8eHMPOTHgNOXZgM+uZUHOCNeDAJOSG79LMsrasOf
opDowW4GL0RAgm7QQ+EhUBqLc8IhWALHytPw1cBNkEjE4A6VX1tl94eSj/lAUaQf
M3RutUC551n5DsPmaKYOi4b3z5C6jcDn+5RQ8EFwE0Oee8G0LkKAMzXrMZJM9Zgu
R6sgfn52/Nd5kpxVThuNnS49TU21nTPpMaCyAoJpTaAm8n+ZvZUb3UQBOuwPBASJ
gwd4kLZeye4jpATPI/7p192bTko0dN+U7+RGbpk1BGrAstgXj+xksGiJxDl/UPwc
VCHMzLB3jv8/CuF+IuhgVvF9RqhV3OcA3ovpmNewgF0mG/9MIW3lHxSVTELRRj8I
RGgVMDIWYAfCi5QQBxsTK4E3DSLGo7lphSCCoHlqVncoMPQcNO1GpWh/3FQ+wTJi
0DSUovgsPIVUckZqa86QGjB6WL1FLHaWKMCU6v/5I0r3NWEOMhWxytbqVIBcO6HA
KaNKYwEX2M1owX3aenBp2YVPv/fxNF7D06pQchg9yHT3uH2OyFzjgF10bMD5NCUb
5xLPlc6T37676vCYommsON9F0r97aLD816Qffb4ABNwuFyUMYqXO98DOSDBiNkB8
HCHYxaxilynrT+3foKaCQfssTG7nTiNWvh/8bQVcLra/u/u+i5K4ELdoaq7USLqM
QFLJvdG2jwnEY3p2kOcA+vCwispO9l7Ib8+xVv+oTJaZQJ7JqKxi6IfT6nMNi8iv
6JwdLS4rt5aNt0XCCP5OP3zo7Q8J+niz57HX+GaNJae7M9EJ0dCXnMATwSklD4Ni
nepq2vrf3PiKpUiKVGZgv/Bhx67lrA4J30E59etqtI6RxeWR6iaNy3l1idaZvcpl
NWvTp9W557Fp7ICIkVNRn6kDQvPeuSK5t19iyRQCkrfv/Eh1GLPGJo9F2A+PhmCp
O/jzrPlAKSAwaD3+4SzP/RDEV6Taxy6Q485IOTZ5QuFThafQgSzH+oYuFCcMnnFi
JdpNt8hD10CUIqnA1yjQ4ISg+IeDno5z3rbU8VEwNCggbRC2gcVqrveOk6N7I54f
PPhKJA9q1+JtJcmxr8QX8lIfN5h/WHqK/QzxGMBN2TRKTWbCYgUVdelD80a6MW+B
fpxdz1VBYH8xPzbYVoaj339/xUUzBdwsnsg3wfSwrwW3r/g94OKZ6qsokXKUxSE+
vIyDiuIoSKZFYXFNKghzs6m0IMYr+GJVl5J1PZSpJK3In18pYqJPpLNjmPt6wqET
amkEVg8qpt6EzVws5a99wfa1RzhH2DrXXPbzXPqQOPzIS5b19+CmDLhR/BcOjRqv
h/UBwNQ8+aTv/jXiMSQBI0HPnxp9uWLikur0sE8uzvT6pdwKRMBdk1lr/Z8pnXnC
XoTwIYB22g7Hte4fZsh5x3eSrQR0s3YI3ULYxi0sSk9QMnQC3uW3L5nCOuotQRYL
SVg+zKaRGIOldYpez8NaPUsFVOtuBo3rK2ibQVPO2+at+P+xS6gfZpY7iDkD9FpH
bftLQXwrKpLqEqJPXdqB8wTMogKWRUV4MtKK7EHpt9Dy0AzYTbnTgJ5aj1Krklnt
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EMJG3FhAMCnsMFpG0kTT5as0p7Mk3TSD7Me5c2mYJj9hKB5iDt5K2HSAnew8tMy6
GMu63/4vZFpK+MN9XLfT+dmhxzQW+C/h8oWsAJU08ohyLxMBEd0KC5EnJeMdjqOn
t5+Wf0Ui1SJnplwIGHvF9UzSfAvC9SO5tdcaXpk2VW6d6Nvvo/d99OZVCUB3Zd1o
xtsZpWo+6SiYOi2yMhkO+86OkpnEODylHg7qquSZBICjht69SR6OO2VOebXa5CbW
Wh49XQuaFtTLOC77T1fLhqP+R+r6KpGP2Cni0S3NcLMPkyfeBNIULhTQm30iy3D4
vxbP2xdYm2DWsqf15GzOmA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8432 )
`pragma protect data_block
TNjRY8/3bnaI4FGXpcRxDcSScdvvYrUak8OIL0MkESx/lFwc5tDtkSJ7t4zoRgsY
ljRqAL/ePNLX9Ofjz7tH2ifFQXpv1TZCChB00wAwCJlCfq4xIl+TXKZqhseRRUhZ
WW52zWVEOSD1Yh/yTHynWM/MxMgmlCMZbvIHOOvbgIBPp1mdqfIzyVKCPymwgo6p
uOtTKFMRzvANtfgRTtIPEUDubCo0NjxPEfepLj2vUVAnUUmcnLLC3mfv09d87jpf
FoYHgYk/5XjfPzFunrV3u2fuUZCGhDqlsprhJrAxFCuqsOnyKOG1dP+cvbPhcgod
vXFLadv1EKD6VdEXTu1e6GUc5GtzeQ9fvbu0er5K8/5ayC3P57TPbsyDAF5gGKxW
Hs/EgjP4XRpcOQrpt6HRVoAS8Ky7v0S1DdaHXg1JJ3oAyRZqZ1yim+oOv2jO/yCv
3Jp1ujTy0AZ4H/QVXYlRVqwFAwIiKmZzg1U+sLPA102hbE/xyNaoDTNaRxJ+pD3g
/pA92xRWR7bzJt5DAkLxz0asPxXg5lbupwPdGPTzTCR2cE04d9eEC5LT/JuKzjqR
69aOzhWeYCkBvj3JfUGnaYBFkEtRgAeomdgOle1IkjYO1GZAkvd3zkFfJS0swnUw
KQ8+25zfcx2QTsLRx0EjrmcoH/43aS0hejP+Dq2Jg4ZnrPZ/IogcVcAeA38svaC/
PyOdkT8uxVzIWbrluis5kdK0uNG/DuOX9tTPSzmoGF6Fl6KOQj0zF4d/L0EZZWM0
2O5ojcfUWgDVuX0dAUv7CYS0T2uXbdjrf31QI97xsGyCYsyfHOrPOyjYCsbH821g
bV4WAUSP3cAYLRStNHsacSrakYh1BiwZOjJshDOYmM75LxCjdXhmU0gmhIdZSUHz
n/S38zjHP2v0Q7hKTkiGrZcON1WfTJdQC4nguxPvgwcojY0PZNvCezp+e6ZYJRic
4WoRZHX/4Rq+w5CrAwRB+eAZgxUh8heT5ZSm96rWrd0Gr5tBCyst2weZKrIh/hwz
5pZweF/z9+yQfaiiIOhlGBq+hUL+cZFmecwBwLWN3U9IAUchI/+x2O6NvwQpGhPj
mhluOKa3R2isl3DkKigjPzv+YOmVG4gcS/1pLTPLoOrOvFk2ZPlUL2LKVLiCTGV5
deRx+9OdD20foeyJ/cs6q1nLJw7vo8dsswPLq5TUPr2Z4gk+6PUX2pdLhiWt2KF1
wcmm5ER1hlVKdKbmLKn0/6qOoj/DhGkxkEwWHKFvJxsb3+DVo2KIJ/3w8EeCKL9R
SvGyiIR8O9zXbUao5JfgWwu6W+zOeYzkgectaQptrhC3TEyz0n33y9Y7UQyBURWN
H7o72CQGhtivUy9hrsVcrVLL/ov+n1IRkxQTUYGjdFl3vkzT65cUjTvUMkOVFlM3
FAwcUxghx3SGh6V+TMhJFRltiFY203hMN5byF8fQGMX/FM6aRzHAHhrRqWM5mZUe
/rB/nvw/WZX2Zn7K6610egzC3RiEghDVV9QPmMTxUBLJg24wfIJAoOO7XAbpb1yA
wd9B9b2vRPA5VKDKduH0Nr6XBnEKl8GzKu2HRsPcY2btCHkKhWK1SUCDax+7nInv
DQMWh8WbvSv2pfRoHS5OHyMQ4PsDuqqv60FTcNJ+UKOC7ztqRn/dSU5tvNzuSOrA
9R2GHkMiEJeaG6ZKJxdlXsf8DQ6LYcTzBYtcfL7e60jbkbBAn09P8dNZ/8yxsFrt
evRpq69yJv12Y2qFGK78ww6l7RPEV17iEnbiyAejtvkZsC413oByyvts5BQWCm+W
hiUujrCwwQS9x8SE/+s00C1GV9YnqyBHA7Hoew3tjy147tgr5G5C7dvpUAOXRZtM
tiZe1xyhSpK4+Wv4mRK8AhQH+9OSp+Qd/6YFzjBTTTezIiaUEyLe+RQJCXXJGgH1
61R7RItV7ouMSCRvZoaTh3afnCfU0GUoIrFvRyu5I7D7SZnuEvQdNrWXUEJfmW5g
wBvXu8DewWB4ebsKiM8HeqxygFKY8ye+aCL+9RCPSW8NFNhR8mgPehgm55GTZs9T
03Wz31tJLwT1x1RPvF2tc1Uv5oWvYP691pqPoTX3VcSd0tndELfbPz4L1fGS0hgX
UszlOix1WLigmyLCfDof8XqyFAsG6kCJuiZicUnKKF7mgBexLiJwjWyuwpbSuvVl
90Xb3Y5yLr4bEZzwl3dQzfwclAmy02ZKOk6ZXU+VBm0fYk2++OnYEVtkG5q5zhrU
srbQyb1bVMJQlEBGsrNF4FnoEbKEvFU6tHsQ8OHiIdmoTKnJazaUAgh+10r7B1q4
x/69RGlVEQtWEyzRBlF7jJVrUZU3z06k9tw8j6mtKRmvUsjRAAx9EjW27ubT+hMo
QNVywPJGKBYFKjaOO91rV3V3f1e/ck4MmvaT1NKPmSgkJcgBHIiWm8UUl9gPrfiZ
Nb/9cZlS7l7FY9qy0DAB0gsGKKcSxCAsxStSlS3pT7I/4zjKTsGkEfw9FANvvUd+
d+bd6bEoq7Sn0OPRdGtvC+5PwQh45olKRGQCR2JEdlU48kPxzxRbvj2SQ49sEnym
W+r7875gJQVqCfNFagQCbsQ4RtCeLJMgrEuz5zp0rK42mjQPbpOTt50obSidMa5P
HLDBVZROo4N56sok4iK3EDdXgxp2KFmCUBEFEe6X29R5qIhiCUAauJ2uSbvIPkBR
vziK/Ha/WsnYQQ8uIdF6IjYbfF+zs0g34/jxOBtHJLyFW0ipes3eeRdsUNkiNSRB
fbB9LINAWlbVSzXNsx2NLioB01b4wrqe5Y4yKWESsoWLnK7GakSD87gwZFXWq/Xg
oR7Rkw9f12NkTXJeigwPmpHduEfGH8P+T/8KDr9NKTkAp8qVbmQcxuDfP5EbFhQT
h+NME5xnsBjEjx3L7FiDBsQXUkAwCUoReaxbXbwLBW9XooTIrcZHF9YqOkpKOsZq
2evcK7LpZfcUpBnOJF6G5Ep9HF06sslxUT9s8Z/LS2BxmRFgTgkmjSwY2B/kphPj
U2nlG3nmReQVqsTmmBXKnWZ2I+omid1sI+LAAsdYNx2jxtzD5y7ogXeOkgWsjjNp
YYlt/4kf+4VbSPhYeOOIQz6dnStdh2+SObeXLsOUq2SvEYYoo2UWeMbRpkH/ZdAp
CNMVcjXvhZLI3WV3MrHiNgtNQ5vVhDqlQjwvLRi+st4IGUIKkdyetLlnNchB2Djw
pZywZVh4n9ijx3qsfQajkNm7ZDc77JQAiyCpKib/6BrOD4qTSrgjtEf1yWIij6Qm
CkSKK8WpqICdH8yhyA4wSTKVY6TlDGg2iTT7mzxdA1W84yGLzYFTDSHwJwl6ncqZ
lva23cHlqvNFtwLZ/jbhhSyqRlI1vbWMQqQyvXhUv6e5cOyrYm5+r85z38eqM2L7
Nm+i5oS0L5jobu9RQUVqNb1ibPUPbXfpmLf4WJGp0xcf/AxfU0LOxk5yG42jJssg
qJjNLfwbKVBBeYZPrzLsUzxE8aM0jshIPqt7OdDg07su5WX16Na9HCcwvsT0c7PG
J3VESB2WOGz+OuzRCZiM5PkRbFsSUVqYpsyoEYQOetD3pH7nrMYBENnljRUAc9Xl
T7UeehZ6dZZ9ggRRf1c4bQxv88HvmBzH35Z009dscFKFcbqZoCVxKkVRLDLp1ufH
dQfNkvkS05yid718F7RVFQEkL6x07fq561IgPmFDIfoturGmQWFkX8mKriyZ8m5X
ClacWS6yWh1XcFgtbG1/gx0yW/F7dhh1oOGT0mNeCunmFfTEbFXXlGYrqeYrNPXN
aHc44DKTSAsUBbI4puiYjrxqEXnc12Qq7S1nf1GZ2Puli0h9E8J+qDYfkpbLjKj9
+b6WWqa4mDNXEq+gpu8pOBX1FVQH0h8iMhc8kYeb74J2ePT5yytjwpiaAAIefV+y
Ct6C+ru5CrOOZ2w1soU+cyD5bGatE45q+AuqhROfX/hH0n8f/nJfIe7Os8FqPzEU
YQpYCmQq4IH9WYGWvLDkrCg7fowRIfm+u1wPaTSBLTxDiLfIWhc2zCPQdVg82qbl
riPcU449yoqsf+1ERhZAAEr8b4VGixIQXbTQqsiWnZoS2wuMpD3EWa8t2LbHfPq+
b9iRLDUsppTXz1sziC8XEHFo+r4YdVE1RpoYqjo5DbD1jAhmoKOeAh6U32D/rdKc
JMVy1tmvDrTDQX6C8Y7bdP5IIjbUSvNTJUoALg3vqO/kpA9Czt3eLGDupQGgoWE+
4QdnFsc74K5lxogEXBevOxFrGwMuDN1haaj+vvTg71DQHuFsVrkgNw9XtxPSuKvV
hEei5R0LBDYPsAC473WprXvAolkMfgCmWYK9l1M5hBcLHgqLBwxjIcjjuLBWFJ7N
Q/7rkTkDsFJCE8hefVPeYPsMgFt4k1mZOqPGJiseKS/hvdccBhHwczFn3ibQutG/
54kPVMzu7MzxQw/NYN57YWyOYWhIYaxWBhkkBtgzhVhNsKFUw18NKC156jzZKmoo
Jrge4++l1z2MRano/hR3aMZ7cm541+t1EV8WbYtaR3vXgkmoqW9Iux8zVdv/CsNU
ifAB0S2e7wNAWePuUy/noGI/U+kSvhXIvWbk7rf5lFU1g55WGevvWSDkFi1iUeiP
mQK8RFY6RI4ZEZbKWIoUj+ZbMaryIAYtIGZj1XJTOAq22TKMSVX1mgv+S0BRAKjz
f08pxSoIhCaW3z632aIM9DoCxVNI4v2NqIAPaGF+3YMydVcGnhMSl0+fmholBJkN
7JlXsw4RYT0BXGxcLR+9kQOspaYIUJP37VtJ3LOe5RNuYD2E66C+jsBHnK3gJqs9
JuH+OMa20HO4AojyTSYfsaNLNxqYuF/tXXzBs8uu4xHX/eaaD7wFX+5F0K3F0Ygg
PWvxZ9Mx0tnuBHGQYw/cTz5RFgw9A3bCu0E6vowoXiRK274a3Gg1OSOJ37pawIOt
6UXkyyGz3HoY9TnsBMPs1KCQ3sPo6Afq/fvEapjtNyPi5V88QlXCpTWhdX8FrnAz
+sywbOMcY19rRfJ8tfXh+K4bmks7u29j1ovbsqjCxDLVnJ5873nvFehFfY9HjkV5
Pm7ljvyB5v6JhiSTmYlKvaQor3dCfSn6tamuXRGrhArBfVQy/RXGgSS76zF6To5C
+zrm4NiC1PUte4JhiRnNEMhaD8j1z2G5h3MgEcLaskWf1IE+Xa+csKFdAOiJK4o3
pkl+DXtj+pL+pVVNBPQASXnKarEJOknAzv1MhzpGvU4pkHj6GHKcSYw1uggtxYzN
jwByiuN7jmbIRby0pKopbQMA7TTcJ8Vp4bbojz+nI8XVkB7p8nbB46lh2Y4eY/h7
mSWvwbVQcVynmxDymyG+IUOmkmJw829r8Elry7rGV5rOIyKDlJE3r8X1A9TSsg6b
3GLMezu5yhtT+FXMtmJ3TiV5sdvXmdvTjLFZserC0SufQ8kaEf4DDc4FKvnoJdCU
4dxCVCiR9aABvSLnoBcyhMfVbFmOISLlpU+MbJXCgWaqdeBzXz8mTQbDEm3pltWy
xa0+PHELaWo3zRBCfVzfIIyUq13Wt1W7dEHAOCNQ+qpQMWX5/t1+uzqy0rNIhsdh
KGUEoWsvDj+d7ij5V8w7S2O/BffjhYKD4WTpRZW5UKPWePfdhZoLHZvaUWTkIjq9
4nWEYbVtDr9zjnTZAS87HvkHbWHvUHLyRJB2ViJKZFFz4Ctb857LyfKwND29vQSo
wC2JFiEL4M3wOeBRS4hJyc4d9pzuGI68c2p0xkJkaIIf8TRO+oxd6D+NCvFwgG+f
pLPp0E7gi2u6lpmwHTjKN2mnGRK+mjFuKvqJWCGJqVGM2HexqV+35p8CzKrtNwBP
hh4rKGUUbtrTG4G4vtzbxM3EkgAQnpJR5I8Yf7GNTDIfEmE1gfxJyXWbusnWgftb
EePXEZ+CWFb2FHk9Tg7m4wWevsaljBl+iKJ4N17QvDDPQzfWLFYtfA9voE6kZ/A+
poKlpnmWfpYIUUyikafqlfQFOTGP1lOoXjM1pvWnu9pYrODYijVXvoODcLjKM6H8
4FaepKBNnQoPydI9LclfIupF/YPOwZzeSOFsDMnObt3XErrR+mkbgIuJBFm6E57L
r0jI6e2/KTj+3WtF7VZZ+ZoriKDlO9NjJHznUEfI0mSpV/DyFR2kWf3EYSODw9sg
YGaAmmTeEoZz3zZ3HIrJ2r6Eq7i8Of2QcV22tg2qiHoQqrFT9RBj2o/LW8YiskJi
kSW3JQCfwyyHcbe6eRsSYXIRABvOc/AeAWoPsPyBJwTSoXPL54wwVw04Zv0mSEEi
5t5yBDriX8XIbnFwMTJh6tA/+HLm+rimfpg/hV29vyFddOa5hDWuZJ+t+PDmLQ8q
oF5276jVMtAD8oby16C+Tyf602Nq9Uw6LgPe+O+zB0FBx1pIwLuOsLOqqi0AFrBl
bkn/dM000pMnWQM16yPCZyID/bKZSsQtTRrLjqg9bKzAD8fp21xVA4HiSq5shAJX
yGxxUI92C3Yu/TvhggYtkJpBsdn/MZfU2ogOL7rJT5xWS0BzXq6LSUMQUGC8ef5S
5syp5b8Vgz9nAC0lI5wBCQ7OkwiGSUnjhUhVc8XKkL4TB2RgBamrgnoG3D+ZbHGm
0yO13zErXY0z1InOAPQJuCG9sjj5gD/FHx6OK0uNBV9B+jzvC0dgfvuXM8M7xauw
boiCyHG+vsFkkjLWC8n519XOhD64earAzilz6aUwwaxPYM9ZGTAw/VpzL9892IuB
iELIQcVzbdwYtY6OjLz4NxT6bfToeEZ3S3SfgkUWKlqr/FvfAZk5rSVwwdu/mjts
F1QF3LvfsSMejx1C5/iyczCcw3h6gH4gabZ/S+quXPwMrGvIOjPQ32qdkhfP6pmC
rlz4tQWLxBUKT+jKrOPzh+jqZ33KN0V10ePNyBNzuJkfI1uEDJwzvVj6Lr+En30P
m56tCi/Wh0UTR4ntswB6LqCmRpmaJGT/SLAnzha27ExKqN232Ko62eQLGzg1OxxU
AwQp9+RWwYdHNSSLjk7T9TladWewSnpKSCKXIZuRZTu0RI24ohPB8j3yU8ImB3CB
pAbtORio1PyIKrfl96RABF6IoXe0p4D7ft1bewunW0kv1kJm3aIrOcYePi/KwRu3
s8+Ja7Q357okNah/X1z6Pq/nZinW2PgJg4BC4TLLxnvtDPjvQ8euR4i0mwuwmXrk
nIzJDPCbdaxOAX6sUmgZoW5IKEMKT/GJZqn0J2JlxwVDbREh9W/H/qpwE3WxVh1B
1EgbWwLsWHFp1/xqGGlqVTdYdK0OiMNggbO+t6k+lROwGtleJ7rPxOmayaZRSPoU
vDAKcR7os7nL40PvDhGhDYGurqGZBGKdZ2eNRxWykOPGSEVdkS6AX1FoqXWJhu7G
HECYhGasR14ZBQqm1OBcR1HhDti0p7YPdf1Y5TocnJ2qRH2weuP2lSONe7/03t2P
VqLHzC7LB0FcwfWjoPeLeE6R1o4BBHmTfCXk6Htufyr1Xsk+R3sWVF7QZs4BrCHM
9HGiqEr/5o+bnFU8jm6xbwFF4K2tCrZk+nr6srh8F4KXQfyeDyeTEZ9YO94PUjpG
O/XCZSVgHKX81eM4RmNONNDIq6E73Z1x4U+v1hhC5J1OOvIAug9vHcyWhHGrztGu
7zByu4LKAnlWInYtVuk3n85apYRwfBpJO6sYzJVsOXJkq3adBakvThVI+A1sftHy
n5pzaPGX2sCLMu5e4j+vBHtpcSaah0pBO7KciBhfSYiMMyWCVb84b+4bNHDSKzih
KoG5DUAnwljinvEQCtLBj1SEQVX8MDqrTwewE0oJaGQwslxOHALpi09wKDjS2MtC
/Hk12ThSiEZ31Iexs9udNjnFaRCtPbJ20cC7tkqgh84QZPTLootxXiCUsMz4Hggw
egtoEaqYqN6bx4myZ+3m6uXuNdSzwUm45rvTiyAhzOifvPDXmOGGNamkRaXQLEzc
PaW2HpGDF9ZIYnqVFtQ+SBHSPsctYHnPjeNkM/oZlNYOIJvGQPQgDbaiuEzMmtNX
SS9k9Y4axmN2YBolOFDvw51nZgtOgfJnf8zIypooYrvmTKZPB+dU60MtxsUAwgXu
JvHVj+KrgTE5FcBj+Zod79nZk++EdRvKEjJ65T0SDp/xGiQg4GlborjYXLBg7Qdw
/7DMzz+liMCalMW1FtaPNPDggRXu3PBKHk1TZCN8AXXpltf5xlagYMjUInlLNudV
EVjd4fmK2vQCFv0KVgT0PTggZnyl7EoVlKbfPHHU3sKaxgn6pNJ3r8sM05VAHLz6
mqazGfamxKBgfXFeg/LFuq1c3Yhl3ScN7zJJH3PffzfhlTotghI/+QQqXCeGpMUR
dpdFgO9c/NSziZuZP2Iqws8GizjEFVqyPNb39U+HqNRSwzN+jLZQAiibx3sMTU2a
O9rNjXUv2hPjn9gz5XqttAQPnq54Nhone3q5jX4JOijvqkGDy+2QSCMKbufnJe3M
39lEIBAjRLzXz49E8obuhdBF4l1D9OIab9otOzy+I/UG5Ww4SujSYteRtrtPdSRT
7a6353YzdSfT1AuC8CrOrRbWpNGwDwqy0iy10zOExRgom+NGy+jPIKKwsR+4bOTy
iK663A6VUOx2acS5oAHDzZv0NyWuD/RuFiULLi2mUTAoOiMv8gUxA5JdvxyW1Nv5
XVtsJY/T3nsqmXrG9L9qou/LMZ1+LkRMUm1qo/cX5y938QwefFoLhQYra3Qa8WaD
kghqQm3U62tJ/UBG360hEWnA6bOPi+D08jWFtHbbpq4k+EwrBY04Pr+03a60iFi2
czGNDSm4kQN4eY9V5Ru8s3tzuWrjUxtv7HY0gP44KF70HTd2Z7L/kgzthRbw5XEE
l1crABvu7lKUYglS55j7QcX5IzDle2SYvoJEQyk5poMxaJwK4JIiuq9x7ofU+1PU
DbfkJNeAq+F5Gw+aKAc5sgcpLgd/KqTm0DTl//iwAB1W7FWyHwFSTjyCViwOVFit
fUK/sl2ZCbVkEJE1hFEl4eXR3XXpGs1U9H/D8zQOondEOPurqo9q2AsnwSpoQuDu
J5jEgdqXnB3BVRNU02wOOmRpfLP5BRzemCZ3EjvY5s28JNpdc53zc06T4XywmTAg
pYvvi+FJqBZe99pJyxMfgRQ7UfnfB9SP+0N0JVC99GE4WkTn1WIB3YflnBFhWYS7
slQgjdtRV6nQXrIcb8eFYP9o89vp5bTD5QEke6GZtu1RSrkJ/S1Z4uWixUpbWE+8
tIiEmUcwF7WG/nzwKsoXkTVND+SIt2osNbwA9B7iDD9HtE/R3tee84tzYaHvlUyq
eRBxG/xxReZyyFQHSMVSTXzCuRptWIUSLKie0zNTUqKZV8E/qjaQ3/6RIaijgdhd
lzkcc/CZMppTtMQm5w4aq1abUvKQKjb9nz5kfT0o3x7+ZJob5ZHPgwCScqVMdfls
jsGBzQ2ZK8uRcGJiA8fK+B82VpKW9dEwx7gAdpBzUj/fDN7MOrloJq9Z7Q+WrH8k
+rYeMkLTeYjZonLydkSacCBazWNieN2eGraOgf69AEX2BWlgL8lNbIjna3PYL6dG
U/EfO8azXucqNOLdSLO1I0tYm//pca9XUW9d0DRmTRUjnGlAsY6t9UpE+mUaFNtX
sBtox2vC3L1G1+sgQjrJJBQcdPnXg641F2iowNRY1U4lrIuCoMc0kqzk4HR1hWFV
Oe+SH987gOwJgZV5m6sQfaTfENk/SjSAjvxPKdJTm++G0tO0hfnTVdwEZjJrRfOD
tMy34KUIJAxM55R6LoQ1N/2TynFh74LrbaVCHyR1TW4OdtPQENX74AJeni+uD4kI
i0G8Rd7IQy4cVtOPQnXMzmT+OzrcNN/I9YSqAVfOjvla6tJoReUxaS0ZBQiZkS7N
R/R4zfwUgFfx0Vy9pA3i/q5a/uPDLLxtc2FLjxo3dlR26RiBK+KJJZdoiJUbCtCe
rnRZPi8IyNcjLKPa8/rObE+JAYMKs8k5+gbTkuSyqzJkq8iqxTT6GjvcZPM29VFO
yHu3o8oy2mnhahOJ2uO8trsBN/9mIwZoxTQrWVOgHHZ9x1Y/Nxi1+P58tiLLQ+A4
bSqLzPhJpXQ+MnXrMgi2ql3Jj+dNb8doUGDvsQuRmLxnF+IcQLN84YGI3g6l6JXi
u2DlZ+NDRnW4M2lI7fGobOGWnaP3S43acOpP7hzIHR1SbxQvKHmAgx/uopUCLPfK
apT/lyw8xuCnsgJ4ykAR5Ro9b8bT/jYkrZa1GIlNWby+qDKF9T7W+x4IwBSBsFjA
JljhpCFMO8oyYj7H8tyALHWBJMBGU4pjxqIOu0VEN52N7Fv4E0AoH0pQpWc3Lmau
X7UotKozjJTrsdYpmv2TfTI0ukkpfD54qi2/dz9uVNjJlY7Gizx5FGVkXXZQfvxk
eI8mXZmOCUUwZAzajJiJ2WIZJeQJ0HjLgF1IfhcuUlOxibnrgNAwSEsZbmwpB8QL
OFGK6b4ov6/cPrCvbtUiWEuoP+Oqruwun5Ie8BFlisG31OfPlk/xyEvyOjDcNi8M
y2l7uIc6OBs4MMcA+1PZhnMxX7jBvCrg7PHRTgJVKPRHyUpf+7E5Nrk1ESFrIZlN
hF6iiIOnztBqd53yERqwl3IcJDJjP5eH4X5+EAZDgcJurTz4FcWlZKJkfe11CuXd
Nq1TD1hmoolEfwGwh/eJYA+WKcIiguG04AdRotO/TkLilM/qZkFFPnGfoTADYiPL
hDCIxK2frAeguI9fg5JnQ8vj3huBOkdatR/0BcTqVFpeA1o/HZhRVZ8fIhZ9Ih2S
dxSVJAaHQZAu4T1pUtlQTsTpwUzTV2eXRe5z+BMlQr3I2d6X/MNQ8LB9lQcJzCOe
50K4+v0veGAURes2TxaOz4ynGpAIz1/JJHYiahlRYluy5CRf7+wq5TRzTygF1spg
jworphToocQ9duKDMIgfYhRYFBzPT9UP+HZYrBA+l1Vp5tT35ynE0Q1/p0eVyq44
djdC4bC5oEJs40z8w5oU0W5/9EZtSIMVi5szx87BC+fEaun41T1X3s7NmcclaeIK
WQH4JQjadY7esLG7Wg34yE86d4PaP3XwzMWNIIvtnxZkxU+DolHR6bm4I5+VLMnE
zWZTgkDShoIA5djDPXb/C6JuQQW2skkT9bABonPDZ24/EmvOQUoOXi8xH6kcIz39
MaxS0YQNbdNlIzWaIAZ3gwnhlPycVSvsrOQtKuI/9ZWaS4OL4wkYbpvBoufG7JuJ
40Ad//hzEPo3jhpQQ1iRGM4r6BStbyk7YpLS25tA5Jg=
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dMrjhunXqWWWEXOnDM+/QAk5esXE7qjFOKOyY4O8K3a3hoQ2XeFA9z0KOfDIH49M
dDtH8B7/bL1VvqGFMDwIvjIsHYXKxigUmcpJKLNxIjaZIlJZ1+Dg7BVU5kvMlXFz
lPlFvde9cbabQSm1NBZLdnXVmgc2bpzXfFtNQ1RuSKsVy6oRIeu40cyA0KY0zN2V
SJuzXUolU0S+CxNo2ME4pc2neCrhXZbUl5uOVYn8f36rzpbJvXry2Q1moU9LQSI3
AHzQ7YEKa0hRBTKEBKyARKo6jYxiNSmAlnaWWPAFFVawgxvZLkFpZRtbfpG43YGV
2B9+B9H+IYOdb3vDOa0Xng==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7216 )
`pragma protect data_block
q3ibSugmaLxuNpduO9IBIoDXKHPEDxTB9lHxSYpn4yArKhZ+OBspFZCWpZFVdqhN
FNUfUGHawVJGjTSlC92B3rqW3kgzyBQWdccXFzsx7PjFlfssdkG8UbMAV5YAccHW
MH/zdobI407eHHdOgDswWL0a4R5MAdIZH0i2yFVpGTpnVsJBHtW7M1n2obpXHkLU
2Sa1X6O+TcIKJa4nLy7KW4jmziZyMROb1UB22K0h3x19+QLC9GBl70z1HInEo1QU
gs9X4HSeaegI2K9SG9jrTV5VHat6yZozmWCVnxo93Utmnu0aQgNTPytSq5jQhWXB
cY8t9obKkdaG3ye9QwgINRivtmrUhc+PHE7DmQRMXSW3v0oQNaYT232et6nkG6rj
7RzdvLva8C/ObvrXAF/z4N0T4z59lsEQxgcp+vC4/puz5+T/KfxvaJVuf/S79050
Ju/IG7OI+P/J/RxIvF6Jy3FFJGNOyz+gFckf9HpftnOjKxPslmIOT0Rsfl8vbr5Z
g52oSKA33l7DiA+HoSts9A4tcDEcsStGv74QQ8a2z6LZIsIGqpmy3tUQd+3UXJ+0
/i5e/59ZdeeTC0vcJg38xuf0PfPMlDnf0O21QmIhWeJibxKzmEf4eVVM43mZt42V
x9EJNm5ybgrm0wmgN8sxSwjGcrF6o5arAkkTl4Q4de84nrfRQP7Hpov8+X1wER1H
F0ePOt2VE9eCnKrbjYb3KBszjR7oWUDg8pGb06+wdjpdiUkVJPbQghtgtaE1G4Fb
2yi2dNs34OSpG2EI0dypVJF8cvqjQ7opye6i4GDfyt+7mwtnbu/CiXjbNLf4e2uI
3za4xmxOaDbiLsg40692lc00eE+n3q348vmTCWr2EiR4PU1ZgxactBF49/UYAbOt
TMaldFKZM2Ow+4ZZE8ecxOKbdAMnbYBgnJJpsjvcQs4A9h1opw98v50RCNXfbzoX
MWDN2jdroAE2riou2BWO0mOWXbu5JQwqAoe5z09saTrpobdGuAx+cUMIwXEXwa0R
6ByEdbBcq0hslnzzCVND8XqYPcNbodw2DVvLojDZfB1g64Rln/GDbXkEb+NXiTfO
XT0xTCEDR/CP/j1W95yxxTnvzHtsuLx1UIUnqZ2dTzbrQlj6qeL53LcgyX96bNH2
VvIeBnMRh+HnoSO25lTfdT8Mfu/rmRrhXI5PzN1QQk7l48oucSw2gRdsJmvQ3cK2
NdOPYivHitcypiHkK5KB7FmL8Tv6z8zEnxj7s/f9VuQdkX11sw/Miv0BfAuHIiuW
7DJybFBN6V0Gf/rlPU7ws/N2dDQedUd18H96gsu6CoQkScl2BU/QJljuSbAShLX6
xnkJPPZNLMLm+KwAQlccs6O/DY0Xx2WWvrrRtmk+vtCvCk3x8LB/Fv0W4PDP6lEB
3YDbJd4TsbaUWbm0meNcaeHAVPPzGVk+g6WKMCjz5JTfl9cyR8RKPUzC3wJqCn7k
+iTpntc9W0MjfzDE9G7aDl1fCtTKpOLJr01xPRXx/Cn4Eo3WbgWfy3fCWl/zso8D
s3ZjAo2Up5PatHUMt30L1fReFEUSUYVeGV1atnGew1vd06//9Gv4fFCh3gPVXYkW
MpYPBjhTC4erkbzutu7Ilp/JDXHYFKAHni1M2jn1WF7TQkpleuQMdHG9C66Hq7Nh
d2ZNwYLGw9Hr1GZLAgWiWfUv61sqzO0/A1elNtvOPKtw3evrjIi4SoSbWX2u9wvC
/We57g/N1HNS/4iAJ3+YX4ZBXC7dlBpfi5wijWlfjNGjUR4/TATnyAFDUvZdTJO3
KXTjcQHn3UJXPHuqxwbzLP+69QUE9DoEvB2f9qWs5qf1xwJJKx0WmNrPPsQw2b8w
6bLalWcQljokM+7d7jqK5hbI4A8Pktnf5fOpNSMKNoRQKgdfPkNGgZ7kmnTOMaQ0
agOoz7jCL7+gBB9a+b5EmE7oFTpgco5z3eLMm+QkYDedbJSMZhxRVmV2Aalckjb9
Lkt5JP38pWD+Vfz+TFT3mi6s1jonvJR+NVQE/izGRli4QugspLSVbOcmFBHQ0YZL
YRy7Bg6ssl/1YdnwYcjf7jYfDSv4vv2sRzUCZf5Z8Fs+BfTy5LGTf6uK+194QNls
MKYOwyTs31Xy4WRy6BgHje5vDrB4Qvrq8jM4HgIBCzoH0gvHeGumenQhVOo9cLLo
LlcO4EoiXq3NRxY70+IkhD9PithUyktzLkwYR6LUMGtbW0X1nJxWoNT0IOMcYUfM
q3SkJgKZWUTk37QLYt5D6qk9lpUgC+yS4krmyWfj/d8oaAiS07Si5kFDUqv4JBUr
fqzV2X07y29yjVAoB/8+Tg6e4/roylpvSngbzVTyraQJhFcrxr3MHcYQo0sPiPHE
Dr/NK/9PlUL9sy35yUTZ70d7J7utOshj5/9xusUx0LX7TiNh05MKm2zQuU6yKtj+
ujOVhZVqcqleZ6rKwy4pPjB6msqX79vzhTOAIwRX4OB9rFsDAHFPogPNnUeGNwea
08TnswCoxzjrACciX4MkFiXTfAQWn/n/+HNTDeojrCN6dZV2ETASeJ90niw4/Dq1
F6xvwx0d6mNsexjhSC1fbAkGf6jBS8XdCTO2cafEuVILjosQtkTfwEO6F90c6z3A
GIgIw2PBrkI3SufpHaKlMJ5gNKRdGLWpVOWZ9mHXQ1p1IiBZof0nP5m0+R6ixZ11
4EJuaMwzNZCWU2610FsyCePGqiZnoLDI/Hgu/f+Yswr+TkaqNmPX/VUjm2wPAIKT
fDxNPLWfiy0bfYaG5kxIrbiCcnQtO1jK8twOzpyBhj1/mIXP5mZN32GsQaC6zzP0
k6dFsg8bQ/Q0BTEWySHhhjW6nOSnpQ+WROpOqpPp96WNZPOf9XnMCQakBl/rOT4A
xjGxa+WJsKcEowczzT8tC5TTuZrGtoOcDnCfcN+U+Wf9073IouPkeOILSy7VKNX0
SeiZUNTGTPfiB+G3y70fdy8uMf9seIl+SnL3Ri8K9LlcuhvI9JMzCP4EqTxcB7UY
Ngh0DasN8NsUtdQnwEGEwyDE9p0lTe9zyvYOe0BrjLKjXmiE/2HkLhWMrsCkq8WC
fwQIDHBGaSgmXoNq8gDg4sOizJFcGDo87Bl/B/sZX+WtxkIszldRwEqrlpQW5azD
Nf6Cy/6rXXkFIfEM1rQ+jLjZc9O0kieuaYopswWzvPGg+uivPXB8mgbg5dyWj5Xa
SpUcGj5zf3T8/93XzXQTk/novjT1Bh5EkpW+3CNWycXg1iwDSrkVu4K/ozFzKdCP
fqLn9PnOxd6Z7dYo5T47R6DK59vGYMXjTR9VOx4TN49TQrXS4hZULEjBbA0+bm1c
9dN3srIXIN/SYn+RMwqqM1+mXeEr9MqMD/c6WArbtp8lNBmLbgawUrDx5oJeW6n5
Neme6VXw0rKuCxQdLAX5g4OkrmSUMjqf0s4tv0+HpGZXp4pm5B2ba1kuMBpzBCB6
AENomw9QGOQ6TOPmLQYdZqUqJM3qrN2YsnIa0qJcq4AKlk7QMzpGjvMkwukPYJkx
qLCb5OcevNjapGCOPqoGWrr7dz9lRlVQ8cdRG0Fd0QCmgsCmu8D36SvbGVaANqvV
hTWFltd9g6EMXS6NO78RgCCDPjIEBVkr5LPhMBKZCLkRwKF6iOXWNPqtVSJ1SmpM
ih6ED2zvx3RQwkQSuUht88s1uuYCTvK/Lrwltct5Nma2I3Y3nW8G2yUkYezKKROW
9YqMMHCoQ4fyyDlxcH9cJwVkfR3D6XwTfA+4aIXoK17CYL+4ds0dvS8+Dh2ZBJ7C
RFgmQpRQb/oJzIcOilT5n4/tIELsr5aPqEQEbdWmZ/ZpPXJugS0ZkFiJ+6GiKXQm
lrcy/H0SjHkJTvJs5cVzrDLreKxCqpq82j1JK2Qz00VFqM1bhmEOxUevLVoKW7yv
tqyCebkFbK4zeXVy1a25Nigr2HD9qiZK5QlvK53xtdGEBAARMtbZ9MEMQqx7gQq+
1wWhHpuuieSmQprg/oF8YgT1OLMCx+enWsqBBMxfCBGqK/PyK0fbeclA2X+ax8Vc
9/xWluFdkrQq54KXVefgICLWjhia3zv/pYE3kOmGYroH/hbjB82dXYSZuYx5ZVFN
TCr3iX4aRjiVgQ+ZwZhOl/mVfqMCQVPLKDw/OrKNxeAQVOS2bNII0rgdQ3Ks2Lsv
T6JMrdcqMYJANmZrXjYEjh5mNI/EicdXTXU3pU9DGb0vARhKFbWMOhrEiGDJDI9M
vx1fle+mG0eVYUrgbpbgY18k6uWh0vyJZ82etfC2L7o6nG45xu2k89Alx6vVUgG8
XowP+ofdZQG3k6D8TdmuELiOzbZuDEf+iakN8hNKcg/pJP64g5UUN5j7Sv5+AdNo
JgfYl9znlZX5SkE9tKxQc5O+5qvc4mYO9HhgqY1DnP8ORlyvCfhSm52qNOIDiiPU
ENHCWYSkBmnMxkmfBRiFskOz9rSKTKriNA5RCVrdxmbaQbFbVk7lqhGDGEtcRM5B
C/EeTlJ9phajBodF+vmzSneMlj/WQp6Qdlrl3WRLUme6Fz9ZIiJ38dJg7vAcE14n
rns8JtNIPx7lo5wk3SY2O3iyAR8JKtU3QK+/TCcARk0g486nV1QfSX8rTL6fsqOM
5otkpuJdiUSGK+PbyBem3SOnR1/iP+RrcisydyeHIL3PubFyV88M34p1y7jzIW36
o4jklSxDiFUAhXJug8BWkAgo76sNfAZPE5dMn08RKOvvR/eEmun6cdDOZtRzOgKr
F9A+yfREdbwPeEESilKo1xtKOLiX/r0T9/zzroToTt7SAybsew/B30g6Yzx/wPJl
F/aPymMP8792xIUISTzQLXO7KjHXFfeJHgz+3JHoutu40MTdhmEL6ouTSVF29Rlc
bqoRslpZ8/SJaUtD8x3Cvs5Xw9IrB1K/eWQfozmayu6ocbElL1CkGIx272K8MCaD
0dWOV+o4FBVAdwaTEv5ZtVyY9gWb8QyMW5rFsFM71w9Y0ehEUcseA9uxxDF8bVha
PSNEf28zkPIw0Nloi94u7wCPWKcy3d6EJJQMuaL/S3Y18/hPsj+WH2gZefHgb194
78aZvpYo2akPvgUIuD7koj59PHPk28UYbAjqpNWDOcBooTHyJ1SBfw0Xku2BXph3
lV0n1FzRFTIneltqLOf0QAYBZR8xjyEKK8UI5P4WgPeIco8PrH+Cz46RdoBQdBv7
c/LTKyebtm7qudp0sAZEDRhVcVj//RsCIeGFjBd3r63o/7eOGQ4ostv5XDoXPiq/
Pxjxbfqj2NprZnOnB5XTwi+lapyD4D4fbpE4klLfBiHmIfyrlqgH6TuxVegP2h8s
LnVhO8uixyZVLYsWCHHY6SgWS9FZezZlcQWt1XWvNnui8uibqZny5G1kuc9mm5Qr
XjQUBCVw7qVh7Pz/vJYFGsFY6ZzhGgWEJmqGASwmNO41v/tjCiXSykasA24b4UQp
IbM3gvE/SCiGDWIyEgtV8aVf1d4sw4ZyNha8ZElDyNmJNZlfZD9kg9MJhrAflEtB
E7Jg5crWPHuEKFuZZakyvf6dzJ01QGZ/NL/oV9B8cHtbHfi3GAv7it25FAfND9t9
MT2lqGpVKO8kku09WBr9p7kqYBmefJoCnvCLdAleEi/t1lXgnhiaay1i17TX2R/s
wAULfNGv0NO7wxB0nokHYuM/w4tvojoFg38seczPu5fvUh+j92V9eSJYKIwdDGz4
wo4G9DYcg+OYYwVGSxi1w4PDsEVLc31MopLi0dhhqi+QaIgmpEqVfkDajw7HIBMO
yDNjvZrROxIq0as9F+gXIu445w2pBh/4UXthDQO8nen29DGpm/A2xUR/AoUu6g0r
5N075LSyTGlBi5i/AiZv685yn0AOybKeAKk9nNC2S4CCtdRrgVb9BXw8lU4YP6bT
PBIrryldadm3jSarj2k/XjsJaYsc4khsGsUkd9Rlc/RR1J/SWZeqVILGV3LL153o
zYP4llglz4LCahlxLus1jylK9Y68I9xB+OfY1VXkc+wzlnrg+0DuBl1RV3ujogK5
ac77p1iLVgDSxFB+GAQWL8/WKWcGvAbAXLcMIxsErCLlbrd8HaKxnWNRsEeF4uKy
NcVul/D2Mki6mZbf9MwHedwaMwQT3njMH94cHJYd9xcJjT8XuLmTaP4pJPwz+HCA
FIAe8vmBPmoD9rfbZjeDc1o/PwaaQTyQnF6IdmGcnsq7USVGDgjgrNm7O0BJB0xP
4CQo9n0tt15GJIZoa91Q+It83aVe/fzaaVWvQp2fP+rfvtfJY+AfEg4I6JVW6SEH
tYR+WUbu7StAOHL76y5v/gcbGMCb6fLiA0CDf19MLfPjclaS292GUyMA87TApD5g
oJBKjFGH1QApcbYhnkLAtrZ/26F4LxovSd9xABqp0oaTdghLBED9QsAk+w6XIWfl
hdxPNen5hxrXVet4/XJ68kLJC3zfLTDuUvhTNjEAWLGTQiV0kBAVR9RDOC4qU7l3
4shem4VeQQk2hgxJxzigmqCBK3jcdELzA8ad3bW+JjmxRq3LLGCTE2QDLEOsmpQk
q03dAYiu06r1bSBb7vPM3uYrh7WmVnoolh+TckQWbG2n36Neg7gsHsu/yH4LmiFb
O5icdwMv38SJ7+w6laIxjqNznaWvXuwKOrDROSWuZXu7bOt+0hKwti4j4fh/luJe
D6PW8tBIh++Iyx+/oY1ckopjCdbYnl46gqgClezau8/aTbZgixThERyxgjk9lkXF
o10c8VmSt+P0uvXInT+mowXaHzqswDg4FZQeVY+N143IiiAeCohPMP91ZMEQv4LF
oDj1vTr/r3LrdF8qB0YW6Yxk1i2fCWZRUnCgxhr2lgw2zW85vZWxsibGmd/n8+5H
BjUa9UOYF5rMD70UV9fWr4wmiaQppXmdGTKLo3WM7vm6m+piPKvll3NVE09PIiQJ
L59m5HE6QG27K+biPDWG/EWFu7IpWhxNi73hPX2eD1MxlzkB7Og4v3vg2fO8QQMS
fOA4JuixGf+BrEfcNnZ3Mn1asI/a9ECDDLcKI1C/A5gpeBL27sxKG7TItzWMTsnu
F2HOnqt47DE4z1oT1/cbWWadRj9/rJ77TqDOIXeAKtgLAHe7MJUCM0Mdbpe0u5EO
+VmPmSqXEj+qZS1ncrp8yWNI/DJehOcL3pTXbEDqDab3byvKCVPrbnj6iJZLu8IN
akSfStIFGgTmO73z5c0shhOgPGEWf8wPn6gpWwhpDKL0nMMmKUxo7z197m1PydEv
CFALS2jNQ/ss8a3HlBPTjXWOsNsvEjTwg0m6SLjcBOtAB6bX6s+c5RfxHLzrZ94u
fNY1S5hhSI8b0Tnd5/dIHk9ft48xwxLzXf01D3rwolAxzs7y0K0lADAfz21Yf/AY
XOwn0+7AVYoP5Tk56ege9KdNikP9WTPEhqmWKulkcF6944ILRBAmDDWxheVkWXl0
RQR2VdldE3aDI/di1ixdfwuxGUIRsWiG1wsZZCP23weByx6+w5PMB+c6DRqmM/fY
4qM+tiDOb7TgIEWcLI/G7lbA8bhahnGY9LGYKE7THiS7EzxiZf3kaUiz8udCwjHN
y+UeNqQx9AeaCZ9dU8ZZ0u/czr7VPd0pkj7k8VvgbZoI1JGCjL/FIS26rZZnskpe
vYemuabdfd6r5nF4uEHv4gSOjUmqYY4SjnwEZlVI7zVV94ZjUkShWmatSdJGPyW2
Ig8Bdq/EPSLUfJnTeyfMxhiY2PNxnFmOU1RVgGZ6pHrHwrATGba15jad9mzaYMKZ
vsGMui7cqHKd/zIJ5XHRb7HLtU/YAIJJaIBvPsq45x6SxnSEGtCXUi2yC9wbGdvl
jkc3BfF5aipwv6rBHa3yCNTelMJipILrwBqMtULOPREE+yG9tUcu2Gl1aYNPqZSE
wE9crBJT3YCsYldoFcvYa1cZaN7JnMeVIrSOVX8gx43RBdPANT789c+1U4toKgFQ
y3xU8gkMuqZvEidPryokEQjFc1s/uXcQaPudmhHELpyruLJTqn105qpYhXvVsyJF
ILc7BtvKFEj/06NG1PA3syMUiubwBuGMIfeCyHBdc+8ta+p2z9l4iJIhqZhObppU
QRwljoO621meEnIfbzh8e8sRxf1vRzWuiS4Hvb5+8Li2uHB/lDgnpU49v22JH+5n
R1kMxVylkG0Bp2EzfZcfKZ0sdzUq9K0aJrelA86u8s7zxviFrU6+qJFn+WeCMYuA
S4sA7udJzT7o/VaTzx0cfyz8m5JHDqRHJX049ZL2/Zrx1inY0UcCu17hYXQmkrpn
dY43i0aMb+jTnpRWbkKX467+NwxomTAhRRCy04eadZ1+ws2qEquFa1TNmspoznTO
Flsni8KaTtth7Uy+FYtlfuxzrTa7ZC8ajzmzDEnk28CWWhFwQ7NhPCqDg/pl+804
ghQD43xeZUVP9SZ4ZjwEeZajEiCkXsLNC+Hrc7eOjyV4ItoDYjfxXeUmssXyM3+F
Wq/6OjeotZvvC0jS7LV8qaPFv1pvzfzujqMez9zp4/A5MbbuJaUG0Jt1jPujdsW+
SFJaIddWCd9fvav1TF3t5QqzGSHWia5NhsPIUTWg+KvfxHa8SxEvpFy4EuhS8yba
0R6Sedytqg/BwIy46WsYmKIduhAYy2iJx0LZ8IxjqiMoEMYZuN8RXn6oTo59yDxv
zYWpF9QMBtfK3kqSMTaLN2ujmqybqeVGXCk+q9gugvqWj7MZhLyJVDanZ2aee8Lw
z/FgIy3ZZL+wKI4gjNsLy+7lJ1j4HVvSqqZS13IMWI/wX6fp63oHcv06m9Bw7Ai6
1fZHRH9SDz9IlvCCsRj/UNsq/JzK4OcGd/nBqPSBggQLe1HLbzXaSRCQxs5+uLK0
ZrErj/VFSYF1IR2i2pJkR7d71is1DOokm+qVWrBFVrXil6moe740pOS9NEVE8G81
MsoW2jnPk17ZPhi+LrcB59LHEvXmqASPTvyIvm/ZHGcwaGacZ6Itjux6x6zCCyEq
a8kNsOJPz9O8zzGaiOY7kgJx8c+PgGSJrIysAKkdp6FapJAibCb2yunhTpnAlelz
CVBIAmOQvnSMlaSoLatbGrAzjvxF2DnJ0iI2fChnK18w1AiY3WzY0H7ImUgSvj56
RHHXzretaSn8qK8vHyB3B3L1B17xFaLoioIYtIUj1MTID4b5vahMnIF+A4yny5V7
ez0vmVmfNyqLufFx1zS2DFQJE/iNJHXs08ovX2f7Upf01APujbncfFasT4Ce6BA+
r4P8s/N5zZthA0Cxrrei2km+I2NrdjBBkvwlYl7bHUqrjsKK3pcvnLK9ZNfJ4e2e
Vd2D4JFOXU4xK2ZiMOZcnFRXgb+qtZio4v9jkv0PdUvYJks9zaANad1FxTiYc2ET
KF8KTD0H17F8EbUugLNcvRIQp+JuclLdUkKh3gM17C55yFH0FX92XLi1UvebUj0+
7RCkXn9iAYkVi4/s+iOtt0gu/gviXVKl/PbBDr37jind9euzLPH5FCvso3QYMp5U
Ne+epjz65qIjXkUuN7NrN2HB35DPseo8HX4g9HLqLQroxXe51CpzR1+C789ghjTJ
qDia9x3OvwLHZq0WLuJsfnRJ3Cr+Gh0Iwndb0T/lnJ0pXVKvrJYiaF+vUG0BvOLP
jbFvgQ4BX8nKlUazzxyKzw==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
d7wchxpMLuyXhO/b3AAb8DaVjRjitjVrYZHE1GpHEQqObg0H7LUcmZSngcu6U2Mk
aAS+/vq4QgSVoWgYbAdwKl02TGZmFvz1jLkjluommtIHSGBSDYP+jLG/jrvf+aJj
KXSvUwe1qhbczxEOuqrsrv0UfSGPUgjTfHCNI8l3aO7KS16YJS1yYnjdMpe2FR7w
LDKZ1RsLofaFVn2n/MO0I+Bl63TgygOwNSuYTJKydefqUzEVCxZJ0Dl4vZB01TvM
PP5nal0hqx2WO4JlIak2b97NecLqU0LAiM4EydLJyjIKrlMMkqSmpmQlyiRygMy+
KI7vpZ0wT++iPGuDwQNfaQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2016 )
`pragma protect data_block
MYnzFIBWSOphgdDAxJMe3ksa5RvJrWkOKPdYcQvV9/dWuqzVVSnbggzc5NsgHb51
EGCFUGLf3oRqFyaVEHPRL/3aObsl46KlGxF7QXb0RwtlquTVjNKVPDko22TpMrcT
R5ZYgSgB9XQHJZiYtITCk2pYK026S6Wf7IQygGCbKzlTpijiHotTWV/Va4pdG0J2
KWaJ/EJml0SjogoNrcZBi+XWZNwiXBvVU89cPb1r/Vi/IhYCo+RUiGwTitE5Wvrs
SCQvOGvanEiD2RUgHJbTB7S70ARNVfCLmjx7+x6FlagpY9kwXw3govTLYIvUmQ8y
dm4BryPUE24XqWvxAih+5pYWUSwL7BFH4K4W9DK2/3vuDJSCZ0N7Lmgtycf/6QsO
QYQiACkMeBTcid+TauaMLfY1jMggn9s7l35Qk+VxpLt+dcuS0VDeMI8yZDWOTCsJ
+vvCyhoNZ2uzXTJ8jh0WREtL9iUGQogmn2u26RJOMXMIuivPhG5QzJWbIITixyYd
9lHAVFDrEwJxT2AinkZZ2x31Bn8s5WNwJc37KM2iB1u03xTgB+3uOFa8MOBzFRkl
iNGr+Rr6S7/Ibi5+M/ZoYO4kYU/7Yq7GxOi+yaTH3ikJHS0xqicrVhD33bUeMATU
pPTTerSyKnGaNBZPkRGgBmNjzZBll10c9UqSG6yvNTBIrD/3oxRyKDKycy/tsJUS
E3yqJtlYo/DuolAjdkWxLabMv6GZLm+QY7N0Pi+JZYC43wvIS6iaQls5ORw1PQLx
WjGur8DhEcNi7HhDzO3dbA+qR/DVqpqFBz4GdkM8T6U51R/lXMRnAtKDftlVrkqe
6lHlYpe4c6QWbmCxvfxCDeLfEj30YAoA0KJx7Cqwe3gaTsmUJtDhbktjGEeyXFuO
k+VOdMb5WdOxToD8AZq+Yy923DGBrkFK5P0Kz+B0e0jxmxFQZBDeUFWs5hh+f1Fn
x1KxIUxOtJexkNwH9dmD4SpIFi9p59ooBttTzPydp8bO/7ydZuSqTa57e7dWfT2W
ARglhp6gFMynUxv0XLtLSmnkBe56OyqTbwYtNIyQQc1NISUSEW+ghVgHyb+osORh
JOL22AsEK/o1BGvajnQWDKpNbt87sV6ZoPr/v7m+9dkdMm05rjHjB5ctFRqVp5G2
cKUnI3xafddrql8knHkAfWvwXc9d/SJXrxg7n/ZOzSfoZK6Tyad15172cjEismhS
vUhAbSPPsWEIQQ/pMq2s40PhpHZOwHvP3rO5fLibb2rw7acjizULQq6hgCPnyccB
06NDC6tZ5rEbQj2FdSREsVku78UpmijkdQJ0+sfpu3VEER9/qc8es+XGDIJcEC61
GzZJguvHajMf2v3/081Q9W9VEfYClcU+CLTpjH7GkDeekw0B8nlLnlv7rAu9lJnF
HVm9MgUbdk6zawa7ZMCm/+osPDKmD/RwfO8DeEzhO3a9+kuEyDIlGqhKWLBRXSgY
lPkcFu8YFFQ3LlKBWmv2oc/PIEUd7GojjpucyqMW5HJ+bYQUNOfEyQFuvXWt7Coi
azsk4DqdJp/ejdQy6thTiLaJabG+5XQbtNO7hccAGTyq1G1E6FAegHD+zRMoR57O
zDQefoyjENKhisiB6wFEJUJ9riYKoOrePZ3xfzIX7RqnkAdmYXTEXlhOdWFp6Rxu
b8bSt31ryY6xnK04QXgDuEwY2dKmSf5darzd4CwiXtTD6zqoo9dfbQmL64QglB77
+pxIqR2np2p3f2iLVe0ieUMwk8CSbke8fr/OwcYjHfSJGCNnbSSbyLDULtCdh2ur
bWhovqlwX1otPsbmv8jxV2L3Ka6nQJsGylkYIPSOqhzW7E/XEyqgsv2EP8QuxOBM
34AO1IxCX/Xc0OOaSEUY+r88jQrLhMxI7vl395tB6QfcQJ2hA+AvQBw5M3gI5Ode
25QGApqlttkh6SUHpi/kfs1D2YmTiXzNVuNew6EkcgNkkB4fondQimYJnQTLuu8d
mwbaS7ngCOe1v40FHwOZyEuXTfIVmgrgz1jWX33vhiPLkQ0q5HHMraKX6I2wR5EP
m4r3xnc+m+X2hfsY8IyZyC+Z/Qxd390cwjdzvkLgVTN0ff2HUU4s4v1Dj51Jf/9g
y/retZDO0d00i9icKBelmmrO2S50y7PdcxODTEDQa/jIvophe6T46VpF89Q8Dajh
N6JKzoGv1dCdXrWbtRG+iOCLASvvz7R/FWWsDcIEgYuZZk30qgkn6l6KUYJCxOfx
KQpz63HLSUel420ZUrnRYHYm6LIys2V+Q0ZdfvDIQPDkV/K2xv6VrBYpRVecToQK
ntcYaWxJsm/gJWDqUOPBUPhGimBRaMY4KAfaOYhiVC8sLvzdPK+YxKVgVHsT7SUt
5/jTLH/MwnwdQj3hRzOPBCuRY+5LVsXN6tWz5NQB63f3Ka3p9/LLkmAL1UsWaG2d
DWVX8IwEqjhHOPDGYWh+qpOhhIx8FxZXaItqAnHId/HWyNRTVruBR+86DGFrga/y
spheT+9Dm2alncKCWU8UUr9uoHAfdrJ/WiL3xG0fH+oA3zu0u5tudokkQtiY3kYx
c9V0Rg88p1wBzZmim+wTg4JAiMPH5mscbFTbkabJV4pSsHkpkt7xk3s9Qk2MhjmN
T09HHBzzA1GOJaeWUxGF43HTnTK1vj05E21cogABqJQ/LyksWHpQZx3HvgQpT3mb
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
b+LVkkviLg5hMtH/Z1h8LI3gjocI8dwDWI8Sj++TYOuD/H/eNdUcwDp3nXmJ06Tk
A5dLu/+nXVaX3eBrG/QKG+YfAfofAyhgMowzWGPaH6G6XWtI+97RxIMR/AFhDS1J
vUT7aW7CR94DLjoUng2KhJY8HyazLa/2beSlR57XwDIZgEsMbeSHUqN8tB7eqZqA
70gcv+8Uk5LbC/MrAv/Hxdqd1UcXfZb79Dlb9ECEPRd6KnEw3u3W9n6s4j4O1qjR
PXTjNX44QafUuhJc/FSG3JJgeaLSbDUDEONvX09G8Fmk1z+/u22WO6e8MyAyxif9
/7dr+SEv0accMgDr68a+Ig==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10976 )
`pragma protect data_block
3ChofW+o2k6kBdPfFrdKMKKCTzonuSYyaFYh+64Kl9dVj6dciDan3FAP+tC4KZZ/
5AaQzaOaYwQUkJxQeSLLRK4qFwbKv3zO8jl9rFCvksMSp7n1VqTUeJA+ouV1AxIu
R+d7mu6baqgck6/nwrtI18vGm1ItfcRHpdeRj1P3JRYp6OET5g7nchxOzqoBRCuM
2poyVMFKpxkNQi8XRQf0X+wFi+a2u70by0YA/rfT+uqjN7vR978X3SoQOrA4DGDK
BNhA82IJy/rUnox2zDVUw4G1HmB+0I9wr1D9g+jChfJ+Cp0P/OlAikPjDMVLcmuk
0hR+mhJN/p3Wi0GQjnhKvwZQD7RizcjP/BPBZvy9COoJfnJIv1HmVXIk7XyRUx7U
GXElVArzagXTahbel/D9FjIspyu/bq6FEH4VE35LgU1Zp3hLDktEHC9o85ag4/Nh
KsNiFgRbhBElfO2boDysr2N3Dj5R0KdcNmMJm23uUbFxzYPdUdK+hUpTP2xEArXY
1NwvprNmzkvFBog4qbvy/+cDPFDS4q42fUPMQHc/LpGc772iTn54ioeAPapnQfjK
iiLbkg0av048InETQw8JgSqTnu/lSck8FXPrEl2liH3Q5xohq/YZYP5X0k7sW7Rf
hUKnNkt81vPZHJhKWlZq1L05lvFhsQ35Db4eHN8yDKGKzplrfLefHjAh9L7c7T99
IPMj/uPuTq0a5puTTHvIbeengA1TW3afOdmx+0dFE/14IyO9c5Cije3/rXoybZPk
ejjZx0AW4EV2QDLz9SHfSiSwDYA/8e7m+EGVjOYu9k/FlzEcr8M984X1nLBKBIQX
mry7o5CTNxMdqEFy32e0eWBaSdEOpQdKJmChSzmw2vXPY5E0HFP993TjmsuGiIys
bzlAwW8UwstN3Mt9EpkE4yc6rpGNUObg7uLWWgxIKv3iurG05HjvZzA9CailJc0q
2/dipTde/XPYEK8VdgbWT9/OLtOLT4rslCjkxfS4HrMk63xAT6DaYikPz8V7k0Gx
GEybafu/Yy6CO6NB9UD8utVG/cW8ykfGWw84oqP+NK4vsUq91rPLU3oY4ECN6QKT
b/51Ch9yo4GThT1h2KWRRu/sD851wDhtHjqOfgr38o0ZKGAUHvNJxzeAm8RyDn8e
i5npnnLw/cl8ObRIrNy9TmCSjJB88sYw2Pio1RibRrd0GV7+lIwLHEMv7y64YX+W
4m+XFe8HXoIIfo3pzc31qu5r/dKZ8ej44rOmonjJZvTmIPCHfrVe/SbXZspo6Ywv
rGv5xJZLHn7XoE0bHiX0uCY6rP/fOLbsYL0Ys4QUOyrB3HT9sTu5+k6wgVZdwtzm
hxqP2Gi/jDyMJ+rClSKiT7Yj/Wt18A+P+D1SNwdu95UK/fieI8aTBUe6NY6bX03P
F0SoKrctsDURYVp9BmhFq6k6U/dt3i88EXO0d7V+z6CiJSW9PfMagO24jVlUg4AL
mQ5zz4uSIa98bQqo2bJyivHyHv8Q1osTsoWhfsqzCf4dTxVBfhoIjc9LW9wimPK8
jMA1P2MddT5/Dgx/DdL6DmkEdkWk2/8JlfYDhN3WInGHFhe2N0qYLp44D4q16ltp
IIMYzAubk6VompAnOSi8Fu/a/AJhmRWZNqZRfzPC0oAPMhdLil2Q2hPPYlvNmRDK
SNw1lyVqGOAo5pQZs26P/6IVvV1RO28v/FovVOvChBgGh2zdjhhkdZJL2wQZgLDW
72tRNfkIfJKqj2VMLaqQkUPDgUYthlX97Y5IusYO1MAH8iF3zSOgHO/M9QmpofQx
gz1aXP6DAasDW+aothG43a1pEhlhRmUXPzlsi3FdatJtLn2KwsHvjj9tVZx6bsSP
iMCRp4NZzHFXs8hNAooh4g/omTLZ40nM1Ig6G5jpWY70dsiL2rREAoLO0lODalit
XbAWAtpT7mUznpmRx46T2CEazbJujj/nuLqTksO9HdgWRKkw1RZFrCr0+JYrMcsu
AEbeSmOjbpkobXa4wp7QMOEl7zwTP0RZmEmyfjyRHdAbIWQlXKQogoCVLR3IIe51
oIBXJ/6XmsZz+jgIkKvDyauL2DH075sPEiwgTiWDEQM2xbXHZV5qjTMWbjsfyOQv
C+DqX87qM5u9+eKLXoY5AN58QOjRBrKWMpuP36nIwyIGJUCQnFzKXJND+DPzDWA2
V0IlBUWDmAnPGWS9z/xkVbqZULY1BL+cQ65NkDxxDvFcHbg3XnvFfBrmnEPKNzz5
FtC21abMDRWa6ytCaRV6zf7d+BVvTZHuUIxvbLVUAxSyjm3q8GsT35n7KV1TPHsw
/IrIHtp/b70cIHkMrdhmxvu5QOvPcXG1gEUs8FV2r5XOXsHQGQjX+s0JKTljjeB3
qC3wdrdkIie4JdL+UhBcZb3b+ctjZYyVrpBmQYI/tjOQ3DCkQVKTmrLVQ1wxoXUe
YPFC15ddyZuaZDpZK/jP6/tuNjHVD5yhpN29avLMbXhcmLQInyWAs5Iks4dKRb0r
hcpjZ8fgpD8gBNeKdTi5om9T87MWJpROaKRJ+2CxPLjQtJcGw5zoDYG1ghb8UNaa
r8kjivvKG4wFD5lq2T88A7pvWQ/wFzR7Y9FTmsJK4hAEIT7faVpljmbqC9RxUoi5
k1aKWcJSdP8eD+zxZMIRT0ucobyWV8/QbCmD7SwGYVwaSyypINXvi68BjH6tXBmk
JPd7e6/HZWxaMFcNdAXn0I33elLuma/EVaSg3aCHBYma/ZQTzcGIbOJsXvH/fn5G
Ey+yi8b1pWP2Fjr7YVJlzOudmxsTgcePWFeHysWQaMd7h1sXWCoihqQIivTzu8/D
8Op+oqjHc/ORXOZuEwsQcxziCtA51egN2686E0E4dVnPDA4dYTilDaMpX5RpANdz
3jDNKTqxZR6C+CX28tlZ6EMiFfCRXmdDUNAZ6F+y1Jrgm8HGvMauIHmWLkUfr58L
6SjTEcoXCyYNM4PjTW1itVRcb59YI0QtZ67GBnFG5UmcvgfdM4qhxpbrK83rLhSP
4wB141EDC+nsF6KvNmwTdG74wfDpUYuTLryaBIZo4ouxZhK+IotLux8JfqGTK7X5
06LvZuhPJKa8AMIUgFBiKpzYdzfaAJCdLb74PfWtHGXmdCV6vaA04hJ9Te+/7Z+3
X2xrrq7wA9ptGz+49JogLAsSLmAWNxYsgZwZc6NqJ5jhRBq1GWWZ6+vX9rr2wR5S
vfRfwyMNcFLgMBDPgb3ecTSVhKzFkAx0zatPystF+NEcO/hSLbym5MxuFNaAfB18
YTcj0f/UTWjQijWZOtm9T3e9qNRkqHlc/5PAx2mCzL+CB/EyljXsBstFG0BGhxwm
YPPsgUOtc7eSnBAjM93koG/ASZg+RwcMEXcr4e6PsKsiQ2qyb7VyEsUui2d1L/ze
GCjtjdH7jAoU+23OuwV+hdyNKxNI9llWLdBBonj3/jT78T8Xiq2RFYGBrf3EDFsz
w/E25bI5o8InF/RBm0UASynTzuOAnIq+ALEcSoAdXOQP1YKMzkLSuRSPmx5B62YI
eICFW3fN4HyI+U1Ywtwof3loqGPh2dJPjDBARkVZB9ZS5+GEMxI9BJ5h7rBi9INv
bkKH2nnpQ06N5LyvMCD4vz23lQPjnwoKfD+I4gFcKWv60dlfV4MKGbGgXJear4VN
84j2ei7LzznphsKQueO+OVLJC0xA69SUEDy6jerxtd6bBGuzVfCB+SCin4VEr9xm
vFsDaRM7pIL5L5AZoD4RnZAetIDpSwEODNaGjpID/MD/46KWoFd/IvClHiaMgFfb
k6o9IU+husBFkP4AwpQXyHHePfo6jUmcCpuWQ18olo6OoCFQv3RC1QWlCvwmN6cT
rU5gU1gxDyHqQhIyNAu9Oq494cSoWoMX2VFdxPjeYh/c8zF2b1wm7I6774ZEomKS
4da7evmUacnR5L8+1VWq24tt2jVRSPC17UCQOBpxY32IqhhFmcwy4NJSLnZHZ0Qp
wPNdH7t3hg76d4vferJrSTTgUzgfTk6tmfiFwpo0ZhdE2Bc4BqsDqqAACYPUCimK
qpZvzsZozr9UdKf796GeLBJR61K+Y01DMEFSebbhk4MCkNLcllA8jqxKBRCKxjgb
H51I/o6Xz91PTkf1ezHKJQ9h4DaemvURUf4xaK5Z4BA4dDSEwSYoCJJRSew/AoDh
LBBtrCS1dphSID5q4+epmt6uH6uGNs/Ajrlxc8+sqGr38TGTrN2OfIJCTUc1MwvC
4vdCrtUtOkJkFDJbg6Sp798UwWe/hD9QlFO78udqPRE3UF81PmWSncdhL9IY0AjF
YozvOFrVmyFtfkOlpxB87U71UCmQt4PQnv7RLtStttotN+IpFaWT4UHexmFW9nJI
dJy467A2iml97Fd+8zyWiO2uZI3WjY/EyuXjJS9hxv234dkN/i5hFca/+/dustmH
2F0oOL1KU2Q51Rf7GP2NM9MYyGXiz1F8mWsIbvSv8K/do2fJkFZlxARY3+UNdDtb
I75XHFmXiVhVELO755bjnCEKwNGev77+HLkRl79Dosup2RgkRghzsZt4lqGfZ1TC
Qo+DSy6gQ95M08z8/5sgVN2e12HUYWEfgQQcc5yxqoxYEbLoAcF5JvSYD96/adL2
OJc0T2Md6mLQhOpahw1OakULyPjotovaqXI1XUjXDLb/Nl7kjsOu7mBdQ+vudJeW
4mS1fPdEI5/BM6gppCaTmq8iARryVxoRm5VcEJy4ACdP+CfREXV8RmbrPeUoTs++
mXmuKadIq2px84qv25QeNe+CosZ9f+r2Vy6u+8Lzz+2dZB/hfJ6K7dLwe7zHflsq
krn1wcBuDLpmZ1OQE5RJ9w7n+7tDLkCm8ULG0V3MDNnN0BZ2RxsPU/8FgVkWQ54S
UDTcum377pGtUvRoiZZtnh8nJUwlpocj8msfOO+ZzL8b+yYH6Y2G9Fg3VQH++tq4
76d3fdIr/9F/dfpca3dHP3e5wnOtQ7MEuYovXBfixuH+x05nuLmPewCMl2XDZla8
b7+j8yehXDXPikdqcPIfbV34v345Z3d6ro4CvZ7DJ3VvlaTMhi8BrMS16zGut/T5
CjZoTNXXuwkkYWv7R10j2yqH8mntNgSyLXm4bi/VEdo41JtAwL2bolFhL5exbOKB
smwFp1A5ostt9NvTyxFMdygIxOqUCnB69HekAo0inntMnqEyHFQ+iwVyLCyq4ILO
pxP7PHhrroV+RGVvm9h8LVzaGkqvmBpoUgk80ws18dFh5nD7z2/XB1sEGJ7sXkGY
E6S6UfbfhpgPXWgXyV5+6G/BCKmltvchGJiWkS6lIYPwP4TUdbpKuFUumjSj7FyF
F1ijHhc+roj8SnmQI3JqgvJLNhnORlua6AtlSVxABsj5uFj6r6KLSy64XatFDv+p
dxDlgN5L+rzhroFyiZQ0KwYRgIP68tojzA/Vbvd9x40a9qrGIcTMGw62l/ieg5rZ
OnJy4+JF5sKihzG3c2G1+Y+m/cLsr5b0LvMeAYUOeFRum3exYW5kGtvOmabCmdc/
BdBN27zRw9KeIyzZOBOGa0GZjewGASnJlc6UKM/6fhbofTd0lt4B9C4IA7mJoFhc
dIN5ZW66otwzUnxzHjQz82nIFLPpykZPhBDgweryXxvjmctC8yH8b3oU9FT1PKZa
BqKrkN09Y5EWg2HLmlkw38ymINb4l+yeEc/wMuCpfK4vckbvIIiAHp88R3mIiZIK
0hvc8P0obN00FKIhaI605mhJdorI0QHcICYq7NGRIWGoR7ZtMjlKVsRwccMv/rWi
aEBdgmRyXKNAJaPwuUQrrwqJSGlEjHOOh5LkWv3GjydGbx6SAyQ2Ky7FGSLr4jVS
vCiOI94HDJiC7zN4KDWbWlikLjf5AloRL4Kad8YKOEKlJijCtSexuxEXfifGXBAJ
W28WoM5jvlpDIAQA+5p3qEJ6zW8t0s5sWRHAsLkkGqYFQNsg9PQ1p6NCMLAJWCoR
FjnfyuLghFjaLZpeJGfnNTBkDZvciwg2PoreGKfc86gm/6cU6JyInWygXdj6hRYm
GQoY7p2RZ9ghwssXXioHwsK0r3BzhcfYwNXMYWRPGH25kU1TzGRD3kdVrFz7DtvF
QM3PvwSM0yuD6WFPfSeLwtLqedUjc1dBfeydmYgpOfFx/hpoKyIaLC8k1PePzz8D
Ejc0qwuCduJUpwW0nrx9YIWglsiyLhPcBBCjlMHCy/8Uo60xGQts9J0XcRXoypk4
F18qc/IrmSKMn+K6D8QUGF6qJcDeMa910RXekIDDPxFY6Fa+IzZT/gYFtATCpibC
rl0bTdglaHufO7Nx5XCumvkrXYm3oemlhwtUp7FNd0bS0rtn8OmO/sMEWDXRoU9j
RlAYjFsHpVlzXg6dey5FJOgY6Tr8OehZ6Dr5oOdiDSVjXQZ3IIJPEZqwXJFe0fOV
o0/uOm0NyTLFuhl8gd/y2755hJNYGmMJgRm9FXQR84IeiSdD4AMavP+NOWovkbxW
NU1Bpoa24+0KPteyIF26mJIjvXeNfkZWhq9yV8r5KCsGq7N0gmgTmq3BvfbMajbb
QJlztq1APiRONjdZ5tUy3Cl9Sl7Wlg+4c4AW+EpuzYLAznhIzFKQ/xlzFonVOSAR
1+zHsZ6Y/0vCq6+Gwjmlguaw4IfG1xMO3yJ5HBQWF4mvgqXQz1v84hURKZlU4q7h
XIBd52WgZuEdaj45b5TCFuFHP+CFVdXDLpBpaSKWNDZ9hRddpSWfNn5y0nRrTpMi
YRhq2jVXyR1qlWOyiuBzD7bFKsAA63OtMRlc+EOrBC8+OXKpOpN6qp0rhYGyV3tA
6fDRz/ON5DlIO1SF6zRyNDXWWIu68vASfw/0mS8hLYS5C6boqSkDJxVDIkZnTabd
TytR3Cde6+wBoch4f+aMP85trDOpL4W6euqcNfer20Bl2Lt8p5capW4vtJRLNwd4
JZCO6L/5is0EL1j1ZcsbOKP4QY9jjtgANEvBQtMWO7+07Y3ml7ynGdA5pYKUpItE
YCmvmGqfNnCx9K0xV+luNWn0BZDfI6nw7cyaRZi4+WFS42WYXcNsDIH6G67maHZH
uw2LICpL8YQndfmEEjsWmkjHR2VMunsmzvpQYd6DQlblipN3hsW1stuGon+lYiZb
tD1CRuAhNe1H1DSKe6n7tsaJE6CdGwYAngZgLTT8Z7kaIL4T0hHmLaoMjH9eSU0r
bJzWhBBj3IjXntN2DOxquo0+510zE3Y1d/wFjPfD5tI0oKF8eLe42ERNAUSfkLDg
I0Ytd+v563uNeIG5qot3mzt/AlgEd5g6v5LZplL4fan1WHiVM6uLad+j6M0G5XJA
g6Bur3ONpX1/jLL8yDi+XyqkzAjB2cuagtegtieni+EfS1UCs846QPPa2PAGQ2tr
t3Fbl4vjcjttEc8tjsrfmhE07xmykGz1d9CrK/68cBYpo+xwMFWEfrU3XHm3huFm
ef0PA3gYl1n9aqMnwuAk0xooB52MOdMvjhpopp8TE9m748naQDRzHUsdJib85WaD
a50U5S0XRwGWXMTA2GHc59YbIr/E56iLViIP5zNHJ9DjQn3Vd5hWeVjgrrMdIYVL
GUMU6gZkqkNYbfoalXk8J1h0dEakFZW20N3ogqDSuCRxwz+pOJ9+wWGPQmwUrDq/
CeEA30kO8BK+g8iBMZK4KkuWmiE2f1DP+LTEFJ1IQ0Sq0HKlFJvhGZYiA+LvwV4E
R1EOcqpsl750HphPyF1/OexMBUSvZ0fXvh7sKcoB55TfABH2gNsu0tQ8LlBIT0xy
fOtSuHDgqOULam2fC3RjcjsJHDtA5kozcYecglVn1Mh4JoJDQLulIA0saMxHzwrp
/Bs64qtGfPiwhAHiGqefuAITii+vA9YIH2VeMvaffBmhzlFSmPX8judOUk54FL6C
gaVdPB00Pkr1b/CpbvXTPWwb/3J1oczoVzl4de9Pdzsb4HoGXJEgtlsiJ/cGDHfz
tfO74TG4csaZMM2BYHdW72HQLgfVIJ+drxk4BAhB38Fow5KP+jI8XLDslXD4hWDq
5J4tVJnB8ac/rtZ3ExnRch4gWAzHhIleKuDWZ8wTB8xYojxTzTlul2JTnaAPbLwT
CXuxnBzO2WXEVigxq5cyYkdaAmeJHouA3ucnXNsxfLKb+4RfKQmrYnS+pudmT7VO
ufoFy6Kc4LWkFyDBuBpL6rdquTppj5p1DFck0XBsfbeb7hCXAtprXAX0duxHcqCr
xDx1qaPvhLM25BBFL3uis+fjO7LJUjOyk0NbnIxA6rHSf+7W2csFAG+p91Nb0X9P
1V9jlDZsaWwPWM+4xe7QNXtThlRpNxJJlxDJcHNMkBgQtghWGsDB2nZE4BKTiqg3
XzYCf1E+60BcyN9UwBdtXEcuIumqRgWcUG1TR6+bEBUNKQQDUYUEYnIx9E0XXVGL
/kyungn7G5O2BSDx6g7eSNCruzQnIZQpd+P2Hyl4Jrh1+3yDxLYmlBFohIEv7rgQ
hxElauPox6kjrTQeJ8SL9gSDYoLcUA4j0RC0dvdSVgLjaldjhGIOOKRRS0wnzOjf
dndsZejvMsFltsTJYND0ffPMqpr50pPTZBJYd1t7wPXACEudMiU3nfUs/aj2nNVc
2G9AUt3e6uDQkPVG9JMMjpYo2ezello/ht4YLgm9DxoqQM5Dz8aoyK/fN3HwEeDi
yFI5E+YlgnUOv6jRZnD6yj6jDcHzoXqdg2DG2+S0LPzze4VM5WgCkX2q01Ff2Di/
AeyXeVX/H68yS74ODakIaOah/RUugjsO9N1ep0sx5IxHDI/419ONFDJjv/9IlPuC
Rm28D17zZoo4TTZ+I7gbrTwRhapLwBpHJK+JstyySZxITeqSNgF4VicE6ikIaeKG
vkcDKTBAKeWL5twO7DY3xXgUpX6FNCQMU6gZaE3Xcel66B+oCWZJTtBtmqUhlvAJ
sCM+dvwDAPsVtgAaEbiQSnfnkTNdqUjXGOrhJ3m2l4gNPqakJXNekydsdC0+AI+t
rBv2fJnGVBK0QTEi+JVCQiGFBIPMnn6kENSNCpjHPWEMaR8EmSA952x32PSrBL4V
WCfxbyJDEg8S5vyMWPmlzTsDwnl06qEiRQIHrKGiRcE3gsM+KXylR4GLuhPo2Hfx
uQH1epnu9DU/LIsu0etV4r5cvFIBUawaIolk0hfu3E3TFuDaSXl47oWsvsYXz7HY
7UorsnwGozh22kEnS9/16aJp3z5FGhHsawplKsx3hFkOs7+HwZDxa8T3YzkoLSna
oKR1Gym9RBS0pCTBkkV/OiSejISCywHtfV3+f6UmlY+XzFUzGfFg3HMnOjWXFbWM
puPwYKAHhwPrH9pbQu4JwBv70Pkfszb6+VPVb1CHRrjwGrksrLPPMHBhmQNEs9xL
8VyCM0m5eU3y79Hk/eyXj0T0AlGZF5rXpwRFC6JwnrrEMz+6tHlIgH0u4AIgao6U
V69ZxX2yEQ39nQdDQKwJ3mGqqDsGP9/Qk6poHCxOCrZt3wbVj1psfK3zYRyAEUOL
wJlraLOiv4U0JKIjJ/8mIG3G8p7FlSL+WwQu6p2hvsVV9uKB68cOSIp0CEt6DGWI
YSdnML6FHpbwOb7akDO3iQuKrea5nujQ53vZC0Bz1LPNYvhC7zfYtVrMCg6sbBKt
ZbshQgG+ZmKnNHheSQgcClS8KBf5/y2hpP49JpAr3T99ytvEhEAbLWf/nPBbSdIs
0fTdg3Ov6sU+CQ/SSSU1cy4N/jS79lB5m2MLzAZfyRi5zzfaunKRaLTAndZ3XDvI
dBXPt3P2iY/5lcFZAc5dC91oT1ZIiBORLq17QQ7kYK2sjjWda/xEGaCePgKq65FF
Wdg6EM9Lq1CkykKQ+fcbx343utXkRpF27TXdx5w6GDA95z1SWPnV6sPQvTyCz2Cn
/1kLEUn//qzLVJnQbjlnGi6R6LU559CPEP374bMTkzDEg1ozbksNwRX1qOznh5Nh
AeD7U6SzytAFouy6jrh5++idAVdtRBBe1Fkxg11/eyyy0TgV4v+trDJfAan820vL
ZAfKksUEr3llk/oipKqombpge/nvf4dZzDfE/oCnhU1mg8zu8hLnPWbD6W8tiMAr
77QGU7klpN36D7+NGEiU8L6VQorD4VLq7iSl+vKmN4kCBybzV+GWgRUBoeQu/OA4
adb8RWtH9RDvD+35j+L1T+6TgytxDWRe5S0Wuq5j2LvrF3XYEy1q8VGzjeRdJuhF
eI0xOlrrIwhiHXL7PwdYfttm+++Yn0+GczvRSXnVf3zQTjle64HgnDAq18/VuE0H
FVVchYLAsVA/9JaHJFQgdNmYv3fs/x4JblNt0IPhPrZnxPXfZ2nkghvRII+/lgjs
Uh+8eDPY/bog6LdhnmoJOx4PK4pZxpdxZYiBkckIfCnhNgTu4URR89MeCjY4l2JA
gsStwGfEeIDverR1bUx2s4CPgEqr1hEvkuqDpKn6X/J1s2hV56rqUnL2M0QM/2KT
JEitTg31sTEYMCETgLYZywcVbl/r4FfjLu/3eWQ07qmQmZyzh5OqeJmTOpRCmezT
3mXO+a/ku4LqlcCHnOqPhTAUAj671rryWDJGw4e6zjLq2el+IYu0cNu7K3lOWcLe
DXX5jA77epzhaQYmSdr5UqocwRTb50c0Ze6QYz2c1wqooAP0ct+gbiVF+psr0Li1
hmyzZZG/8aQbe/a6SxwdBDzG0IR1FmyNvFJHTAqIYnTnCz+fnsKr0N0vEP3MB/4q
8wwv552/mWRxJwcqDQ64if2Odpx6vQ3MYseozEk+Xvc4jVyjSpetcIMzTJ+1eVZO
yiCUxcDEJ1vU5u/DexIu3N3U8PWzZ/H3G21RsUkJZ1tcMvNNN8E5pNzzUQ0AsaZr
U/1xL3+AaLXJK3djPrr/8Wu7xbN9+0BNMEa+Z2Ssv2aF0A9q0ewbkpi3WR8QIEJg
QXr8kn/G29L82O0SpGOHEHtqpTGkvzBnRoOEIerJ92d5GnzJSygosZvxVi9nfYY2
QaB0Gpx2SlwfSEfLZjDWs6ChVne7U4elwS+BpacyQ43Je8pMPoyLn19qeqJlAgzL
PeqnZpoF+IZ/ORsiqfyLUWvP6TeaPDAx/0BCzzYcAq6sEAapfZN25QwP0fZAJe/T
NXObhUvzkQEfLIyEliBocLWwK7D1B2P6urazGCnEU/fc10BVKIieckZVacwEAtWd
NOvQrdcmCrLlgI5kTDG4sZOsTySiCTkncCXD369rnIQ9Az9izqRaGvZ9ogzrl8hs
B5zw54MnnYiju4663XaPR8a0B/jjaqUQ4kwWtWNrV7BVhvFvGJJKkv7jQolYm1wb
ORaVAExja3fHGh33ZpxU6zzzOvPMs6FSkgAdT71tfJyAmvuwXI0dM3WCHdDSfglR
bM+SOmeb2xZiUEuWbb+WfM0HV80E/oH6fOxn6mw5ifbl9iIjaIvxMmAeiUPT1hgB
7JjPhIyoD7YY/2yKCiC6QfHSst6yKN4JG8MMkSbFxZucai3UaAwdrq6BA5kzLSkW
nJ1tRV9PTW0uj8ff2+5y11DyPZlx4fBvJP/MQdJvFDSC6Rkkms1fkxQE9nEW8mtn
VnTljGtwac8+k6un1/80hSfy5V6opkDxFKx3GtwKrGjfI8oXN529HCmMir1C4N5K
NNsRRihzY01azjHJgVAI8U6dGsmViN4Y+/WzlKXkR9VsJUWuYUhr4fC3G1Z7QcG3
R+Ki2w3VU+mZOG061Ni8HCpNJ3HLJPNgoeDsS6Ja7qgSdf0hCD3vNX1Qt8simRlw
CA5VULlHiUd2G2Y+OK8SGtdaqiSyhOpZrp4+LqGnk8dboUMmgkPQzaC1RCbRQ7kD
BvRDdUI9Q+/Cgf+ARJ6Qsid9/C5bSDhfOrawIp5ziS84HQCdZ3DakiANz3+/hKwv
NMdc1xBc3uYSOoxjdPzbpma2wDYUh0bNSV0ZjS1SK/6qjBAbg6BNfHDIfQqpmc2P
76mYNIgwPV1zWHy/g+6wlXD16G6WMWYDcGVXPbmi+OcEappeosdZqvUAmccyiBut
ZqiSv1DhL3VD5LFNDI0E+Ec/JL/PZqNSkppuBkpTeHPqz8oXPtJxj446iPDzTir2
bzBQr7GtXQjUPDN10rXA22JBIS6uMeH4uKzZdrxl6duCTbE1SmwEf32iSVd9oylb
OYAsuNDvU/U7Y3YjywEGqwt0GeiMeuYVkN8Knhb/D3kEOD1efgn2msBCaLT67fQ3
ioc2a2/Tf6ifXJMyyyFtR7x2TNHMhRjBGU2o9tKMWEu8EHC9lnF6jk1XN/v6X8JF
BQlfhxIcL0Wy9cWFpLkKfdkLnhaQS1RRaUPLBokYmXSH+FPFoYyzz1904UAYBFex
H/6z1YpRnOfbbXk1cmgM6jmR/Ay8H/cjFfxbTKGYfUo6vDETA+PLcozvcDY3Lz0P
avrb43x6/iWGrS3pkT6OF+84s4dCiHQ6x/yuaGYRZ5XdLXdbc4WECVhhHnbwtj5I
DroOpI8kZpZaT/PnLidjS0AJUXsaVYrwLWWUAzuQ5gFo1wYHbLn41dzAjPWXciZ6
ITMWN2IEzgtVOZLa7w92v8mftKNfrTBTa7VXYT40lh5O2arRcaq7QIC8Xa5Mjpwn
SWyl3yWT/yZ8fAoY2KxQLfRlj/2/pq2Em0QyHFwBII3uMvg4IZnw36reAFSX/WVd
GcS9i6Q1ryMaRPU8f73MpaxN9IoQWS826gsDY6vanf0txwrs2J5pOwJHR3y8RI3+
flknUXIYv2VJ4GIGPB29y1cFoFspNChtY6P7X3lt/wzv9wgur1EB86xAsWh9Gb6H
/0UqhgKgALtxYylBTlXASBew+mZaKQG0//Tdh5gIsjDQ/alA9PpuuaZLzGlQvopr
dCShIDq4R7c9MfNTJ4RUoVCWwOHElYCJTKnUXCVLkvnExJDe4ueZs0+zcA1KDB0E
3G00DlS8AFZGUYGEbejm5OR/1OMXbsuAKxC3kpfX2AOLAYzIwCAAXMypS+UCuRxb
0A+ADbUzB7NwGr3amPYPHW8g3RYn1C6q5Vq7lZ6U0YBqLR+kOihxwAexW3LmSuaH
HtoJMKnvDwp7+/0po1yR8VN7qpFHE8UalBJZ1RRQrjI8ImojYxFAXlqSf1Mr05yn
0Ym7j4uQxrHKSk9XYz8zwxwk2e3uS/EN5ikMD2wJaGpUlHxZsjvVKIZqze/MGsvZ
EsRhdQCkBh1+ghYLGcazBebKn8jxyhHarApMsvdM3ovkPkMZYM+Z+mPyA+wSmn4b
2zo6hT9CqJK9bT64KPl+pJu1fTVwRU1SDPJlJPFNu5IZvXGerl15mHczE/adiHqz
yQdqdJfGPI8CbSXkk2joyZOztqf8xYFdBt0qhRcqYj1JABxgblOzy22x3v40KJP9
2wut7QpGnxGFLWo7hzwQzVmX7QTBOoAH1aUh+0J7el4bKws8eMTHOvptEERFvv9G
9VcrzZX17Q3i4LK49XAKeRCsAG3mn0MeyxEZpxhngholDVndL1nJNVFVnmlD8TBl
6vkxa1EJphHBWsEkgDb6Lyn4TBdu9skV/xcq3U0MBrYxcuC5BXXh330VMPuIByOM
1HNls7FBCaOXubJaNP6uOk3TQDXBQ1iloDvgWyhGB/Wjdmfn4ya4K9TDot7C1if8
lxxElsE9yD1kxR2SgIIioGhh66n6P3hNTfdmTdIuGqXY17u0QZqN+f+KCoFnaI6p
7Eg4DqN/VllwgHew1TeAroH3f2mz0yjNDzzV+0VJUjrrY1O9NVSphQjNIvXGzV9O
5iZtJSi7oKxXWRIG1TWfUSHTbP8IDmHfAGZ3CJ+755Erd8EjfNzvPw2Cpvbwlw+n
Uk8BvhdyabUBTXd+q0BkVlFeXwi7tnAsMqIWr+744eq6moeG/oMadCHntiSrNrw4
o90cVXfOAg19MmRJCyXZ6ltV+x+JTKwlWAQdBhR587YjNP6yEq2m9Zf9MQwgV82u
DI9jhpFC4duBxhrA89MuqpCGW6R9jMk3LlCmVySN3Hnen8uPu8erXPOqKJsHKEwn
GKcp2VR5LTwjfAyY1Vn0RU7PL9QG9KCh18uDYH53+ETQ0z9r/grJYF16S5kcy0Vh
KDFKRj1+YXhJHo1UctGIu4qIcXXLS6IfJKkmxgjdEs73N6a8Hzr0CDuEKtPabLgQ
w/NWFaXEVn6Y/xbtYUaFGfvMXFrMmjKt9UXGWbf0p9MSYMKHRlmc2OcQ4AhpU+00
vGG0i9g4MvDyMBmVKYzM/dK2aUf0JG+mw9jx4O+/1QCus/vUKNd6BHL/S6CnAMnA
TLFsCoOzS5Au8j87GQscOpRsQPeFOx7IsO+w42zgf7zODerYKCz8gksxKIqnNEbT
pztAYS4CKk+3zFynWalBoePYtTpL91NEaa5w+ggwtah5+W1XD+YMeykOrIV4P11s
c2+RXKkGMZNbv4W13PAOzGAv+9a9/4fhqoYm/YBfCmmiJaP5hTDGClYk7hGiFZko
Wfb0TjVyjZa3SkGl8+zjlA+PNOsE/h9OtiOd/jvdYtjC1gyTj9mXVcifkiJM+7Lt
zQFHsUiS5O0PTv+EKVjhWpxC86eUN8w5fIwgEZ0exMx2iIRoSwl6rFVmWem41Koo
1jnNUdb/hjScpZdwnwNif0wJmx38/6KtH2cjJ6JqhotBXW0j8OFGugD5CZvRNjI2
FaQsgAsF5ABil6XtUgB+geK4hO1tFh5XhiAssMUK9tM=
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hP4hCdCmmYRca5XvxUUkSv372dZno4oozOYiJAmuxV8m0BjQtUZQVjlQ31ApMdtX
JKpkGIXVyZbZBHfwBm3MAeLqGMYaN+powbhEnH4u6eL/IuhoIyZQa1eu9UVZwYh3
9t7dGfsVKxrBLeBnuBIbVYF/scFbKuv3V4Bslg6zIUQG1aiT/vIdNxT/NoUxJje0
gm+Rq3r1m7Vp9oPbPWl2Pc8w6/t9A7UA/gYq7rvSxBECf/y3h9Z/OkchTX5RRyNx
sKoV55o38WsdeugIkyXkynO5950DXGQkGeK60ARm6GefMBMPSOgQ0zBanrHmzD5x
oWnn2NlKSPunZfYLMBQ4UQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5040 )
`pragma protect data_block
cBt/46kDPBkH2Xh4JyRdbJX/OLz2uoyyF77d35viuIb9q2ofomb7IZ7S3x4sQir+
uoQpi1lZzG1aAhsTZ1wzy8PgLLRuPpQ+94xGu1pQNy9l3yuyItcwOSIO6X7KLXzO
CBgWD9OhC0EMp+gj6FTlHSvj2t4GMVZTXZ/wm3hpk62Ra8EiW/T3D/lzjRASsBTm
TiCDPj/xE7qsE3Vzlk5m5nQeK/0Wm+XAVj8+E90cOAIotZY21zyP+lNaHwerXp4H
LDgNCWgW4cjXnD9zM8KpZDdGi5aDX9Dr4YaoyPvOrbq7Es73lfiY3zOd4Qlt7DXN
nSxv4yxb3uSxSTUZvudAwUjaqCJAQoMOzFkCJ/F2K3WxB4851UyA0jM5nBdA8yxe
80KrdgopA7X1vfK51YmC2DP+POeAk7lH10W6IFtZb+zrFx0A+SQyFZjbEW6ZFzex
XuJ03EDKE/ziD8tfOemHo5RyJJ6S0IKo64QHTIz4HV/ys6+muyFYezbaOv2qdIn9
N035RVgP8qXvBW4l8d2Fd82/mUbILlceUYpjG82UGyRzqkzMCIvg/LyiaZbdrZLU
F0uARNj5cMOi1V6OP9U1kcp0e/bu8bvhJjIM/cn7CvVys/ifX7KE1NLHo+SiW/2L
uT0rDUyn8TraWqD8hKOuKojwSHellgeZZ8ELKe4D0n6K0wHy4H1xe4rddzCb9mCp
OZeORjyW+dBmWUZiEkX2lBlLpyq4YXxTwF+GwNt5JK+SMySFDX2arcXnc+5hmuAF
CxNwNG39/jxzXps4+etvCt58rU7uZ7C4LR6TqNd/J4lwXJ4Hb+FqrvRGJtpbw6mZ
2S+Gf76q8fmjTDaVKb6ig3yF3IMvs1g3c+72n1gGV8SiZAxpKFNVVNjo+u8WpAa3
gLg0OKGYTOBu0Yo+ZnEeqw9TGLX1cyEJRnNH1by/uydzV2Jg6SdClcmAnutYGic/
guV8LIHunINEz7JfLECHQ9cepQGHxZmgxgTUc96eCz36O8GNBMN0urvRxc555Ak3
0pDubL+ErPY2Cc/Kel7Yev94QN34TNU24QWAut4hwujrKUhqiJlXIEawCdldQLUl
NJCeXN7peRLSSeOg9YZxjsa832AnbsDaf4ZDAMeCBvG2rjwSCgCw/5wdt0Ob36oD
bQqwmuN5n/q/mHOkv5EcJBvCy/Oa5t2byD90931abxjQPBVnvvuATDXyMuSAWJNW
lOdxhyLwe79SrIR2pgKlRM11di1a3wCzSEUB77/cUfx4RnKLquhkdDrUiXIt5uyG
htLs7Y9RLhqqKxXN5Gvq3WmJh/6NVpXkCA+EzpXbV1Y+49YUDT3D06XCrkNav2wR
7+eptuA1bFrYMZzfjLzxxSMEvITptCs5MbPVKCyXDXBobUgtsHfbDFy5oVwIckbO
EEYQva+RXcFOiOz5i6NUQm4tDFTT6LFOR06KR3VJpvRZvi74WOsJLQHFIJhBNZDw
2bbT1HTy36+pMtiv61DlDmEK2YPYcROtQEWWxVipxSRn/kJ6bxR/swY1NEaFOtRC
Kyz8oBV9FQUXkDSXNET9FspYUcymmErI6vAqgs3fm0sURnqpb/I9DN8+HMSoW9X/
hjq/kwukCuaMI0HumsgojRH9RM1yxA6uWBAKE4EOMC2o/CqzPJm9NIb5JH3Cz1im
xrpmr4FNYNeX/lbgpbd6Xql5klWDTZ+2jUIDyQNnAFu7BPry1uAJCI9Xsaf88CX0
yL3gHAA4Nxt2jhjVTGNJK/4UTTkqJKZZLBMKoZjFnYSLdvnKlXR+d1u7y/cmJ8SJ
w5Q/VG1gWSEubv5e1sAFT9rSobLQy8Y02yQ4DoteIVsV6HF5oPoHqxcaYWY+A9V3
T5SYZvfmTNQs2uq7hCM8+sS1lNGn6xJw8mpXnDUBXO4Wu0JVsWIxNzluhmVzDfho
Z/S9gFmsTgcFgTyeznNgsNptObvOfWkWAMJBFgJ8YaLqqoU1Y5jOIHJWtedhmt64
UZdqSxJpdUpNmhUVeGIWHOiwSE8r6/IwLNErOPU64WV6kNaULPc/jtrkprzzc4Zw
IXk7I4yaqQNxCKrvI1e37/wtUYFgAeGpaPaSK1F/JzoGLshR9QSJBNyIXs5/fBNM
ZzXNEGhkHoWCr153EtKQbds8A/Sv5d+gLguwny7kmclR66PZ40iPhTzt7XlRcurR
gktWXrYttUwEqc0vmbFBZjcrX4Og/lV3uMsOxNFCpqE8LQGb+On9/q7GrcGLJcye
dwo+lB3cWSrb413D4FlWAUZlWwjMfcQgQ5BTbiPp7t4nACN4STQj6ASZ8QnAnf0P
1eOirfdeG41vEtWGR92cmtt07sjSgjq9pJ7Kvu2kTgCn1oVvPYiBnHb4NcAVctM5
xPDXkl4A4tn7hN1QBni4IKxP1dby8ZHT/2ckBjGXIfJeUj3cv2AvfG9jL1VEnG3G
aWjKaF9czmZaIs14xv4gtE+o6bnn/B8aTHosSFogEygkpYVdhM+xy48vQJ/gMQR/
WY6CocMZB1PeLAnTbDKbow3IF7z+HYtgKrGiaQdJmC7/Oe2VYQL1iOUCM+boNAHj
Ia2ka8JtULyxfPireoZc4JTmpTLPREjVFDCL80UeXyzHIaa6ljV+xOF3iGW0gIS/
LHNLy7cBr3O1btoIEVaqXWcuZGrhwFRee2M5xu+A9o2S9mnvgHDpS8O49xINsJCE
PB8lo8l5MnCudhVH9bBENGl4wRojYqQDghwRI3dlGU8tc44m9ITuupVvMwQrqpyH
QmKrSghgPtrXZhVntbhqDmxfCypfG205x54UmkAmlHkDIEXiojqCYtzuaonS6dZK
A3mZXfVVAehMjjdMccxODY+yRkvdehn5SvwiFdZqDVdpB/hJlG27FXGzDuJE+p84
Cs0Imi7ajq1F94siSs7R5eHVMRiKy8Rt/H/rIAwfOWmAZ26dejeZ3sID+lhCaw4D
SXg4frGEYprwZjphdGskuNRY1xy0M0ebfpWJ6aKPNgVd5wzS5gsi7rpGChw8WlVb
x7UDpnfoK55I+CQzY37K0Unm59ruoRCVil87Kqrun0iFxtiUgzBdikEB5gFXFxCX
KFzqWE8aAT8RDkitHfXkf+uUPr+W5vtJ+DMvTaO30qHEPQCOpNCadl6cumhenaw6
pNb1YLCaJ+sWrphcudVaB1vGMtMzco00rJvoMb37bnOR7IOu30tjosd2xuVCvzXh
6+eG4YRYImwq+HlgxJVoq52zmyXmJGt+EzCrQgDDyBld6s6c0GWwJJakHqM/2T4i
1npVM/YgsfktaX6atD3A//H0yXZd4M6fAcRtamRAQcXYcl73F7KSFEFJ9fckuAZH
OQwQL4bzzhKwiVduHSa7J/EWg6GyOPbpnWEYqsj0OWLhtI+EDnncOV+9mJFtL9de
EoXnmS/JKfunZ4xpzjeWJ9mOEryx2OO8d4i8X+aBkuNnFKc/G6i9dzPac+QJ322b
2Rh1pFFs0EWLs/n5iGk33S/6fz2NIdW36U5niPnNHd62tpSeh+mVilnrpemTnBIW
tqlokph8XflYYJsT5ZDr3hBSg36lK6OgE3YVqZHONjnmIW1Nnmf2eUv5y5qDzD+i
U+hmau1Suq1vHdJyk0fgLWjmJkd3uzPGDRM4isesnt70SwHmTZ78fpOmcEzQLesi
f54KYOX/dod6sI1s6WqEFCM4L59G0KR7EKF5NtQmCqaVpN0A+OfD3SQjpzJU6V5v
rjhcyVN/qbCOLkwCPDNpVmVprptORz6cKkiDGcXec6hYEhoNGu3i+rMu/1vP4fOJ
rlh11SsojR2XINr2AXLBggJoe/I+JojT6iwLj4d65UIh6Uc4el1UncVR9jwlc6Sn
AHDyLl+f9wa2pXbqAkrH4Pov/p8Vvh78PfeaOZ8CN+GXznBpasBBZeQjriLyrmTf
jXOfeiFl+fVlfcnAR7wSdg5nPZSp7MpeCooAu/vXx+RcAh/uSvkW1TDeOaaNjgiB
OtfUtIQ1opC0tcEcdQoZv+MMwJoyW4FLHl08y/dTc8snbjH9xRHV5Usm4xhOhKm1
uNuzdcPXAG6iM3c7XFmrYORFejcjkCNpdHvPSRVfkFunpdupLQqn2qMt4aTNkYYh
g3avmscAq526+n9zz2PW8WJfDqOFjviMBd1T/39SkCjuTdo3a2H8XRBF83vOTLQt
/fOMyxWuhWP/TN9M+Vy6QqpDXAGI458W5hOawbn4eYTQlyTB1AEzCvOV1OIsEydI
EZJRmhsju/IJmdNfqf5QewbII2MitIkoZ8UCM49l4Dd0N/xIqGqTN5QOjiX0+cCJ
TS9toTgQdxj7KChDZUdT79cxaRH9EJsGOPeslDTIYMe3bxJnDlmWDVclATntrosj
oNT4PTYP82Onzrg7TLFxVhiodgqZdaTYpBRXa2F17ErnVKZnuT8/leF7ndGSISGf
zbq0xL/mokzTuCJcp4dF/PanvqN0DJ20gdLkRfQXgoqnJ/JxxoHr/95rYmHyLzNo
pZl9NMyQoWrjqT2BvRn6RS4LGNQIDeqU3tCKk+l6RdksSAGYnrMrFgFBNCxzoWrT
RRHG/WS/15Eckj9o28Uw5jTeUbLh6k8E3l1OkHKRj8vQTJsEb3LZZHXDYiNZTCSh
7r41edrri3xdClNJYg+UD354Sq0vANBIc9f987g+js8lpxyLxb5FRSiTT9c5eEeg
lpq6orAUlcykbYI76W1MRnf1NjsNmeIa6NjyUbRxhdulrbeembsShg2C0MSj5WLU
KTAnzp4SsybJdvwoAt0qh9D637EOwTwERWC9+f+hoUzDCXds9lDkhfZDKUFauMd1
6e+0qnMBr5Y0KmmA4v7luZB1uJ/OrpKVDDU1e/4h8+aGtqnYSNZCZcg5mHkiaX+s
xi9+MjTlZaQvxUmeIn/waa1xbtc8USlfOnWW5AIWrpU0ReDH7tatUs300ZHFxxcU
xg/T/UAe3d8f4fDl3C6fBj80B2YZhJHGIK1ENk1hPbWm6zvrf0lrr9Vj3hpOCOOL
7XSYiax2lrmB5UzE8ByHtiigZFMFEpopxXQAT296KY0jJIgrYBKK4XbLT+SoLU4o
5AzheuG7MF4KmwO2kex/CRlrbI7x3p1TXDJJvRGDrqXsWzA3OmAYYM/Zu7cKc0Ti
1BSBZ06OBpNl9yFsWJmZ947mwUfqsiTZv5U3KqBNAM30sygx189ILDekmJNUgj92
sJMPjL3h/0hAOc5at3qRqp/DJ0tcdWEaMG7iTbtbewx2kQJ5B75wrUA9jhsJiOz/
hopAxW0duIUG4rM9ZIMRsT8M8cSeu/IFQBfiPlC0Sa99LFKM21HCLtBV46VrFOHe
UiiZiZgEJHJ3vHxgeUO2gSomPl/+iLK2BhSLc+yD87NIOJTcL2/pjYc+6KKZo2gg
BteoDdJPK8jxJyX2xqTLzFJxHG2bD4cglQCC4R2i8hpQzg6PuihNF11zDldLwZaX
LmyR1JmutnbfcFPNKvTIcE/TtaBW+VvCqwJHDeq8aTFZX9qd7EVq2t2RMIevWKoW
QlNGf8CCmERnqiamtCGfzfHpW/2DsmF7x7oVrRdUbXBr7EKj2JG7FU0ylhgXhSYu
/fIcTaqK0S3ADIpxz3O+kwd+wOXQoB/1EY9s9JeXkkTt0NqI+PbWxCSOpPkuS0YC
w/FLyWr2LU0Fj9uPuXz9Dw0esx+vD2t3unSRsZrLQvv3FbL0iQwxQa3W+e58Pawg
/dB9F7MtNXVvZOdy27d+RfPCzuqNDMH+a3/vtN9ksqZHdSQtcc/BF+csZ8M2UQM9
RJ3TH8ixr0LgOmZSrx2VuQn914Sperj6G0NovxsyG28dljS3Q3ham2hp1KXTSMzL
B5g0KfxUKsWBuU0gRMcN2aBPj6Hg7lWyVM+IDTtr3UetxotMhAoNCPATLZ2Xw1Vl
UiSEXldiGUcIz2GlG/t709dxuR4F7nWuEyB65CGGNGBpPgeQEq/H8RGF0T5mM8F0
oWodwQ/24Fw9EjpdbdKc4Fc0rmB7NzwSbyOH42RqFP0BZ0WQQVBCWcbXA++Jioup
TS15q82JikL/ZeLiv7qB0FRKiwQutYJPc5lhD68Y/gHv4zcqQpsQ2gOZRFPFLpRt
e7R8eF7i0uzDgzWjYomLzv+zA1WRmyAw6Iwd+WDnRmgO3SwWLkduktjBsfpCYxmI
dK2FGCOuJV5NKXWZeqQxGXiR5Bnq5xg5J2a3HpzbzyfC1DWBc1x6GdUU9L/z4rEY
FVg6VbLuAsS0OMaHdI187HFoNB/qoCzkTGUXXQv1hlqeFoqI346FK0AuHP9zI/O3
IsrvK8/WOWdDlOv1lFaOplUYuxxlfpfUTVkJ8469yI+4uK84Qr7xA+GB/JLITHYN
7YJgvscE6a+TV+ZDrPJ7vkl/5WIdd2frZftgAWnFT/tZymW8OxAQxKP+HPKeaY8l
HcYF0UfVsgpKR2Kd2zLpQaU0ksU+suCKhlNMx+wqgZCdBwYMFUjxExGs67Rh6SVD
1LeT3vZDRQz9uTYOPsS7xWCk0KSMwxoixzQid8DWS6W/8kw8ZqnXURnmvS+OL7Ha
uT7efY3I4WDxj+07ihqVHerwvuChULsASy+W/GWK6y57gFaCpK7fIL3dNDIzA7eP
2QpWkJQCa6/Ww5S4NMYSwBhXFGmaKAujbveXfE2T9QCJ8cCGLRwXEYTkJit7GvlM
BEB3FHWTm8aoZDBc2zEuR53Xl37hR99Rt0ouEuR2TrEIRkpnqZjVbgoFF3Xs877M
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TvvysXBVJ7JCnn6V82ZHuDYo8obtENE1GFoG+AFT3qc0h3+B7qFtXDqyBgHLcgpx
691x/6jP5onWvF/J0vJsomG0m3EHo+cVRIdmrmHAHqs9jjO11dfYQKpAFGF798qv
r5xQ9KCjCYPkJenLyNy1mpGNqlxPptVTWAbnpc1hc5RRF8o+zjZJPrufYrkL+sBR
ETXpHK579Whx3oEv2MxU15LAe7GzNNX0+H5F6upGB0jx3D/8M/+1dUOWRyv0c8a5
Yxa8ZOkBiEVqxiTmc+zmEprKDQfUDr+aiPeY5zKbp0oPSF3h/U76DdKl1cDScYNM
yIQJUmexxYoWAAl93WMsCw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
7s69ai3ctxicJSRvTv6EJl1Xk7M+6AcuEXlSmJ4JLHbZVjHbKYVXm2DVhCKOtJH/
e2zU1iLiEKvRsTNewHfO0RLIxAwqcJvhZtNt4KQldDHlpU4JRFAwm4QMdNHzEMSd
hFgZ2wy7QEo1RKIT93HTlcUQ3hhjf0E6gIEeLwMFJMkX3UNPmYbaZ8EOhI+Pg8oM
M7+Yi0hd99JFDBois8t9NYkaHKfMFFtXEyQsLzQbFyDVP25xQJaoD+xmwyg6kuUw
paOjqdum2DydCRka5aN0Fi+/1/HtKDknkujfOiCbfzOncDGFvZ6EP+5s7LFysd40
R+fQbCBRfnCo4XgjwZ2j5ltGxtd5AsC6bL/r/Z7Qm6sWNz7/WUfNtoCGq3hscu5N
1FRaauvEHoImZ8DOLT+HmbZxprH7luxIDvA0UR4bnUmxuf8SVWXnvUavuHgeGgZZ
LnzHncx2fGfP8oAYJplJx9suElWNfcuwRH5TzG9lRzwsFXj6JP0vpXNx1sAB8s7o
z4CgnYnXRluQb4/qIA8tF4GTS5bPKT/d/KKC1VPdcm+jycKn94KxJanO5nch3kkj
jByygawWEFpFBR1XhBK6NamtjJfayovDZBDndaFJVk7NJ5wtfXnCtn73FrfGmUGS
qz6mxzBE+fV7C93L8BdEVHG2ld1Qt3l1yczFaSQIxgG2NQHJJRd+kKRZpyfh0VJ/
j0P4ULcBA8koZ/2KUe2A0NSLayLMhImSWvsFNd4QvLcx7+MJ5T/ZaGw4E44Wmm5J
f0A9ulNCSK+h+QcvvBIvt7fNZ/0VRz5xg2xSPs8QW2b2UG+Td31hnVeUzG1C0yoS
OB4GLWSzroJKrnGlVwiSEkUi21QZn6kXN+mCvHSgPwlcPdVINhUqjL8V+XrVnDIs
8P8M1Ydkwy6qBw8qkEYm9BMzo5x65yyBIeH0KoU8Fec=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
kSujr8ws6TrbNV6SdfYFmLHUIptHxwyzt5W+KXXlNOOHN2Ps3cYuq2JdGPaLRIrn
ZjxK4ur+mtBCQ9pU62R+ij32rZPnMm9aEjTwucSqowTwVHZa88AtHcOocXZPPB0z
S0d6yqLIhQ8z1teUW9VrTSy+DKMcSMBTf+X0ZKYa5hxXaHQTmCvib122aklKlKt8
123gEOfdnpEEr5PDonuWEoG1xdPEr3VzNBPhM7rwuvsK8PpCaGY+HfEGflLOnWvb
bXVY4zqiMjwB23w9/XNxTx6MXgXh45zVFkm+lPxpCEpAG0RBgbGKZktlpvJNtu/t
84wH1oFHq5yhQBSJBp1f+A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1792 )
`pragma protect data_block
oaPJ0bpIxDU9i6kBvEFEyoPFcsoXKe1BehqsUQwt3LOCYkrhzX8x1DvEG6hKlx/j
ZGWlg0OTvAVwdQjiRVVLXYaMcuGIv2dna+jiQhUnbxjaxYShNOcREs7131Cnj9qd
huivY3LLDV+ZY3/HqdtJjvmu1zLg6TDTZLkJtdhGQkvBO48zWC4VgFJfYz2lLBNc
33A2/TErCAhanVrVGuOxM5S2uNNZ1EyKkvYoqRgUMA1VQPF7TK0QOEQF3aEBahcn
hynljhSpM7Ck3Yq/m4qA93sQ1QuI9ctVpiQe4FLaQwAUW+5sIYRBYtch29W9PhnM
LpJBaZcyOvPwRssBvflZsKPc72A/z57PdHcuo9G1tDzReEOnt4SQ+3fW8bZ+SeXK
m1ucdKCMtUOS8y/MUx0fHw7YXOe7KWva9+OCMmpT5tETeQc2NhyPyxy1dVrq7D+W
GzYA9+Rf6Mih5Phquu0mR8yABEnax0H/ryqpGcCyZ6J5FCKtAV75dLvXK/TfzZGt
2ocsiURiX16dQ/it9UV1YR7tD+1WNnlCtj5gyYJ2yBorpEOjg/6uIcJBB2nrPl46
TtRewu9Gt7pf5QnQxBRMa+LcK9+rrBa4vl5cqhwN3Hqhh4SVKSbSKLbjOjKRKgSi
U4FpZFRN3mHCmre3MbzGgWY/wDGu8e+Q9upniNt8T+3MN9q0spG2NONfeS6slu4R
kT7b0wKjzhhAtxg0XFcE0DjQjyZgGkEHCbiZiLGx5JQdoHJQXY7f0p+DhKct1tnm
Fy0NQyZvRNk+0kX6GkclI90/tASH7ioI8I6wtWr6a1qtIj1gjmh75NxeEcoxjab0
53viH21hKFCJ44q7s+8W4RiGY1WGOgrMnLYy3D2a6VFSwn1wVGEEZSZwThPtlaNH
ccYPer30Tb/X9iTkP+Ij+ZAnSl28WKsxA6DDiKxg6fke6b0v71kT42EyDlqujU1Q
4tzEgaaWuMiWemma6liBleI/drcGrKsRFolqH3gFf+IpogI5wU/t6BXpE5B0BPmi
2G6uIywZKvPY67WVs5uwQPLY513TnmiDT7Z5c9PGcMC/QRX3XwzxhjRtzdvBE4ZJ
SYsa+IiXV8d5PH79RLs7p2CYBdyooDWbsIBr9KI8qnbdAWsevMCH0P96FwzkTDI/
W60ieYZVOF/9sFo7gr5kPaqidy3JuJQMLriP+LA6E3wVkfoQRAIw7VfxfQ4e0s2K
oXhOwvTkKq97CFxNQQ0hFrTEG7zoJ5Xl9FOoRustup2/mNTP6Bx6x1PLj/iY0KL7
PyEaOiTOV9AOtJMqwOFs5KNPhnSCGa/iWAF57m3uFDXI8znzG3jDLL+M5qO6wcgz
BA03ALwri7MC7z7eKK784lCfutl56hK+O5FhfHjdTAIwDh00/I0xJHRoaHLj5j6W
wEZVsFvJpttW4q92wxpmH7afbjRIG7LW3i5CbkjAqqjIfwO1R4JHhvWsaHutjwet
RwBfOubRNoqM+4B6X6QzBH/8P3mxlCgXh9+zFDFIPElFetBe3gZg45IOhRQcm7p7
+EBtBrM63eRNwG8eMQFbipTuQaz8KukwvlXLa0xMK1ZQZpSFULxZ/p//OMKV/dxs
7NTqfCZPQW1nTA+Nq9a/kV3Z4es2akUwvdKYwqA9WQk5NtqVX6o079BvsPHkA5cB
c0FvOcHEvyRujrvpFhPPkZjRdBvOKJBJSnlZQzReNDgYSpFxcbflQmsnaKG5XGsv
yVJenYkcjon7dM7Kh7VnBfMd4G3HYZrS2fntvNWWsQSpOoV+UudZE4ZZ0JjkS6lc
7KljxMQfzoKEdENPEC6mzG8xJe/agnd5SH18D25gGVwRC10oR2120exHIdfqzW6t
k3Pm7DFIaS4o+x+SI5NFG9RhVdN3xaUn0gx1YstwcUTOaHnbI1iJbBAxvYdoovV/
4WgfzRT7CetrOOQI6nhW+sUj1fg511HCnU/Kn7SvYWxoGYxUBsZvYi7NuqEzRJgb
YAtMZPQxkN3gzzt/x3oWx+GbQVcaTBhhscj4Y8sd35URLJDef40pomXPpnp9n5nX
GXQaIIvdwUMfPZtC84T4AjUdanx0fn4+ZeG8CTJnH5sT6h4Ig0WOaIfAAAZS1wQy
KkTCRUv2+6+RPAC7PVmIOdTJ44uZEPiozx6IQQWn9P459j1f6JNizZEOduvt2VV5
Ugdog3PJKrqR9CVpx+SsAjplJ75iyOKf74llUg34MET7gHTBguD377uxT+7XKHKr
rMJOsfuZGfNUX/nw7WJ+NzhOWZ8RvO4OW0vTbbUJi5P5hvF+x+ONU4i5XXs4jORz
DkVo/v279SinoBWQewVLjZxYqufGlBAOy8maoRRDiDYC1lc22ZN8QdL1GZSMEqLi
Q7zackKR/bnpcqb4tzIj8A==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JCkXbenfEWxp4ZNQMwlXOjZY/UqcEXlDgT/kgx/tVqSxkhWM56oFtQG70xPkySkp
N9Y2QNZU4bdg8SeVtNwOAxMndl4m/UdjAIvzna4OdWa0ViKGoAxId8gJ+q5Gju3t
hpahuHMrNRa+vkIhIRzbq6eoB3dnR9fFLmea/TmmetIPO39E2lZ5U1ZO+SEcAUmf
5CJHo1VfOnKFSRDaZPSJxSOAXc48tVeevH6+RfZJ8bgQUBS93MqpYeQONLzzri8z
0gpeAlM7jhzIE1Zp0dvzYSNBOh9HRgLcKyA+gDvXh5m/JMTFfvqDgArNE+f1gFW/
a0YxAF5NGTVshoBUaDFE0g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 30544 )
`pragma protect data_block
bzT81RNqrrVqXjTciPdCqmv/Iqr5MuvEvElOvftOg3oxhBbKwexL8wqmdn23ShQb
nYVI4/IzvX6lbWrF9AymXf1MySl5gNGk6TIduLLO+4UhnYdyRoT2EOE2xJbTZbzi
yd9xzNEXtXmzYE4nA2vlWnkE2m0ghKbfd95/EG464eUQ0EGMMg9o2ef+gi0DgUle
cUTNFkbZ7bajYgfUWn6e2puG/aiMp/QQUnqRI91/Nvdgcp4SANn2AzaQ1uE7tIGR
9La2WVolnp1uGuqSwm/uon/+J41+pcZEFiYMy4BNxwQU9RZV2mKWWLgs4Ci503ZX
cfcAi3EGOeRtko1xxv/XaA6XvtpXcj870ynGIh2xhkrxWG9hGoeCWMHp680i6xRu
ZmTMfLHd56GMbwPcqoaa8xc0MOtfR36iQnKjyG5gXjWnOfw+4ivICZh9gzWG+FF7
DINaP9udrlPtIJ5eoelKNazotuMN6mCnU5+lYARZTu6DMbIobYFh3fANkWRd94Mh
QkAT5UfsrwyYLzhFb4vezOplA+C0zvS+KGkfbt0xqQ2VYEemi6zOsmA0l+vob2jx
9B194YIsfbzgrrPRlY2f97qq87qpfaLO4OtDfbkP5K4tGtT5R4UFewtED8a2bNM4
6mdFgi6NwSRqbDDBALcFOXPohptxawgQPkrkwtC0YJmhPkvEHAT6HNm/0Kznjo4n
DvZC9M/1jfEtzb9vvZQj2mtfCEeAH63U08VMFELz/v6F4Xm5yhkVGAqF0Mqcll1E
HtXg6PA/zkWq/QwEaLy/OPBsuGd9KaMQayLXO1waBZKTdBnUVg2UDjLmA9WEMhlh
tec3Pdrhu+C8Dgbkhh5dYWVqZtKK+lYFdHt1uzznHS0/+FYJjurcEceG4bempmyO
hQXXutYiFu+nt5olHisg2M+AKHZr0XHPs8tiRVjvZVUT2FhGNx40wYSNJ8uJvoU5
tUNh1kCc3Oedk/Vs9F43iHka8YzEyeUKW+DsBi/mXWu9n057Zkv8NHNaj5ryhDvD
q/ZyfSCicIXjFR36iMDJsyv9xZrFMK6RZY1iZ83/I7fn7+NP/AqPmRSuvnV0PHCc
UAiYEusVOUpEzTtk9YYqs6Kt+XWl1ip6KqGzZlA3KMbspV4du/HX9V+jVSA3qZqi
4eyZkAx/a3suPiRkUYFN3uvULGpfGcX+y3knOoKb+sknqDzTW6XvdtprFCFyiP6W
IJB/POo6/jfWWes2d7RwtMj6/HKty/RdRBM+R2Cs1dF6Fy0Q0PditmGrqS57ajuB
g3CezZP0qsx4Rit5SLTjESkjTIa2joPdv4Yv70bMLGnNydKP9ebnF+Ljnk+52Mrn
CrirYbGt1ot8zbZgXSoksK5gyYoi6Yx2LRInBiwLu0ycZydIjQqP3B7lyRAEiXjv
zgxucNFxdAUJHqx5/YIYeNSigBMJHin3+NC/fRqxXLZZAtUzRmuCL1ZhAwJfe76O
7Xw7ACSYvS5OUCULvwezcMCNrYXKLWGTM+v+4AcxkPdzEpt42p3zKbGNJzTYpU2g
YS8BWp27aiX/OOQEmf/2gGS3dc03RbhmcwQA7aT2D9cFCkJ0scwfCoSy+HHuwMUp
Oqxf9ZrBwN/W/rFWrNFGlEkd9pslIOIzNP3zGfJZpiDItZaWGHyB3aCNJmy0Ssqo
ERhQAHUV5dOGkQ9bfqCkBYu5WY52NkVgNZjdQYOIEhPf72xvID07DjxCVx32AcBX
M8xGo6VtpmYF5QO2dJ+fFNp17LhvXStsZWvKBoFushXPB3LzZUxxf/S2YboMWYvu
iG4F3YegI9+Uf+UvDxqYzdKV7iGudhg0ZmGPhguEfOyRVNiOv2tpmuK/OYxwRun0
Zz/+7IcbV5/ON7kzpj4hra1UT93vMgr+Pd/Wexisn2uGvLp0crqAJOs5UAK9QGM+
P5Qu+rqY2mo4dxt/ehq3D/cgDBvbUKdbMMKDRifmdTtTzIz7oQjaYJaCbXuTO7hn
ASBPgm1GjEc5BqLE27jhSN1QpR7gdeOSRuwFBDdTm1qi7Fja/xIWxYSqotf3wVqW
Sw5LAFNzvbJtT8zAd/MMZTD6CEDjqqqtU7BFs/y1/bQ/b0orprDt7+V/9cRRioNS
usivzczwFClhCWI6eNgtSK5dFGgzVXMiBN2PqurY6/X+w01njZWrwTdUK51+cQhy
iJ1iBTuqbml+yHD9RLurAAVueBldc2Q8060AT60kh9qmKROsOq7R69g4uMfVBbUI
xe+lcvhK64Z5rShKwA0PufjY7L1i9Xd1xz2bjQhuTV/F26TKeWzW/RIJ9tfCSGWB
o342BwBDksD3LjxdpFsyHq+ceTQMD8rCyJe/IADtiTHT07asNIkqwNNMFC6f5f21
ZbJmaqHntHBhU+BvThst/zddZlXlwVIKfsJNTIgaNCckDQWqekFPtAl+9FXwACNz
39ZX9aw1rm76SWMLK1vlFfl+lj5GB3IAoZBrzposS9i09SSZtvjzakBPxfxiHrsM
1O8AlD1jTeQ++oLDWJTIHoumxJJEJfDUmrsL0GU5Huz0P4XyWB/sKSwbvH7BjKEX
AAITBUceX1ykwgHRKgjuk588kuz3l//dzRf0kG3hDDIOvuGcbqaeJU5jZlE4Guj+
4RjT81GEdxTYu/vxL0UT0y6NS+Frinw4OfBi5opCyM7tp9Kzx7rMKcBCbjOtOHSn
318qdL7K7ZM0tM2K0nsoHBtDUgFINfz511MM+O+C0KM4MqfrUgv5MTW18GURMsvR
eLV35HoxNh+jC0a1DpDjb8I6tewle5wyZVHQwD6+lqPBje5KoQfo5VU8CnKXjT/5
7BPYB/k4OeUXPwW1m1ZeJw7uVGaG6NFtfzLV2yNIF0pueWSPeSj8eIgL43tHiHCz
DwavF8Lor5wJiSsBWMNbodEKlgPtyrJ5zp+9LRMzTjcd9qVDWhk4FDRc2hvt8Z8F
JZF0o2l3kNnjFKuQVpA2kEG+INPGZkW1pqQXOT/cQl1h7yo7DdlGWTTs5G0XF4c4
/B7Q1kmW1Sg4zxI+ipMidwFj+tVvxwPWclAO92XGlEEF6mlusNtapwlFSMbkLToh
4XucVToNW12JIlNRz0Fbl8pHtUILcey9rDlZMe8cBDteFlFaszUZU7cnv758/fTY
998Khc4ep3Sc7Vts8vBVpViYYdcUccuZLAxdJJauLeDq+LGFDU8K+CqBbUZYUR4T
JXRMCAGzoabuG+rAfIL+e/8/k7I5C9smk40le2DVG8ZQffBsGJ/LvuM9DrEwacPG
JQM7qD8rt8ICbQoo5iZq3kidhNLHtDVEpBJ+F9pEKRe70SE4rvRqyyIDrJxRou2s
9EUW9h0ojkayLnk7vR/x0wJLwV0qNdWxibOh/ZPS5wV9vrXJYH5bgQwdfzXQ8zQO
9U4ziMTaT/XqdGBl8kqsEkuyROa5P1Ld2JqWz+LUk88u7Qc2G4C5aEiTR3OwZL6L
lQVyYz6sPk1jr6oueZ+SN7QfDhZXD56GPFxVLUh+cQTaXupa3/Xbrw3IX7/yiplg
ATZ8geVA3WYw/5Ha+j5/NtN8JRhhe1zU+eeY8sgUVeebzX73XHUr/tv5ryU45pP6
NLwCQaeR4p6Zy1b/CE8Uans7Ol7LsUDg/3iZ9RSHDFQs3ek/H+NDDGJtHeXwwe9G
GaPrEUMeQ2lMTFCqpfAwTSWemrGw1q3GEJLD7wGkOR+uZjKf9VmCRUpIoD+eoF+b
mLp4bMyOOev7TwD6v4HhmV5G1kSjQKx7VsLlh0Yh4pW1J8Ce7jm9D03sMfk0GZPi
awDdAtyXbk/e3CCJiPOm9zJQn2ywd4UQ7Qux/B73vi92o7xa/yavJNCN0AmYQ/rU
HkBuqbNIY3qNpQhZp8Ulgb4NRGE2nQTa6Mzf4T9Xj8dIahv2WD65QsMDDzp9xFfG
ZsMI08z/EzfgEC8PX8LD832VGeHhvh1/EVK8yB1FW0erX9mzlg3cpik0iSB5Pw+A
LV/cLayQJoiq9PbH3JEMTivTAb45wAAU8ILPT8RRMa7NlCNglALaTjo/JUgyIx3X
wy1hvoMuC/Ks2Da32AzP88ez1pcKqlQfwXExST1pTuwZQvGliSTkG4/Z+fT+EtDc
gcr5BVLge5KgfLWh4qJL1V2UUKE4gtLm8MLKpY9TJ93JS4W+XVmkA+Zarb2D/sbY
BsCOUHc4W3GaORNUNpYZJH6IOC/YS2pJqS7oBXfylXxbSB4tep0HtFqi3e8TVEFb
f3juYFp/8xCyXN+tdDPho837lW4f1sNnbikaeCDwBDbyfKX1GlrD6awEZh6I6wKg
m+Z3Za0WoG/Rh7OdVKCIH9BbsmhYQp3KkdnplmFGe1sdu+MpUwQx5yWgXypXMNYf
SwjQ00slc3RrHYW7hTpKFYWlq2sO8QIRz08xI9XW24DKSwDNuMuDqVX7MTqIc1V7
iNty6g+G3tJ2sYNXB+F9ZD5M/4TkwKZHPEKjq4W1aVx7NCLTEDwMXH6wM340oph9
uxuygFhIkXspnsPgLdy/Xi3AgJWnXtmxvUSg+fe0nZSDpZc24nWWI7emAAcCuGcX
NbxECDt9zWjxlWqh0Ctok5f1AgO9LnkwLr/AtUHEe6dVHInT2/NlMoxavaTPp3k6
ecGP/iI8hvpiUhNR4vuHRuddIGossXMD3sf3cIyteoW3mteG6MKaYpEJprK8u9WQ
ECI3S1Y7SwQph+Uug7X5dE7oZ8rhM0VOCCQ0+pH365qnMFVSEou1eUtrZIVDXlrF
O1EL6+47PjCwJYDraTJnF3P/xadM6ddsgCHJSXGXn/2lIPpdr5cHreQ2EWx0Zotr
VCOd+CLokKLseFbxjIk0Wp9D7s0o0LA+y2F8Zh6p1YRuRmCHytWcOpiaUC/eqUAi
f/arSNKLHsu8DC7CL9egsTAV/P4wn+igUzF+Cftr1aWzyx2alP8AnaiBkwW12LkP
QHL5nBs3t364LLoB2X2snJCx2TWZqx9j/4LzTbqBJzzx69bdgLypMWVC60/Q3yi1
2RmylvV/wE1PRnBBxKTc+c/qMrIoSTVqJy5l96hOR6mn+U763pZTZKvMI21RGAXa
+pavvwya4CmQLBHcBKvepssfyzYcIrjDn0B5qZuJjb2+594/5MSeMJymvxivA/VH
5wZ5RGfHX5dJA+192R6eWHllB505SFnVKLW8a5Hl5rV/N0O9pWXTrJzwNLpZfTa8
90gqiUdSvi96QajTck/II/k04XsTGH+ywCO2RYVD8K2kHwbau93WIW7D9FYFwp9C
IPWyQ0c7q7UDHJjwi6r1ar8xMJJQG9kxK9WO3u+Qy4ShbLIVC9paI+BkQ4Eq2YLG
tUdL7JnKh4g58DbvM7/7xmVTkSpj+/eRy684ROXlRxKEaJWP9nuPX/G1/bbGDq6V
KMCaSOdduDpkNdb7lcfNWPRkG8XK9FVHnLjhHOCNR6u3LH733tXYBSSX8g015G/Q
gBQq4LvipoGCskcEzv8y6YOoXwKhUQvstqMc0SDLX/uAgn7wX6qsO2WHL/uoIDqG
4vvOg7W60l2i+tvy5DUYlw6ldwjbM4PRtBcaMxiGjK785Sk/KwylcjyYiZn63N9Q
Om/MwnYTSdksUOZlg5i54UjH8/bwdin0zdtrHKB192N2BBq6r1iFqfP+vGuw7G9Q
70O8wbj9qoFqX4+iVhPNbQVFqR4ylLYxHomF+SnGvTGpmWtD6UmPQkNxEa1hl++U
7pRd9eOkYJM9W79o7Q5CNR/gpIxZRwu3KYJsJv2jn0n/W6WUd89DBD+2My2CMnfw
lxvYRA7oMo9MZqCsNiphaMxSeTy3jT0T7/1CGCgnEJO8IMnFWETlJ+33BuD8rAd8
OvFEGx3CN38bCbaxexR3HIk0JrGci9FaA/7LAbfgOr1eQCyEaghkWCU3/G+CmcBh
AQJwBV5LKOq36iawL+qXMx1T67E2ZZQJh0zIwI79LtZ+n1qWCv58Si6HZv6gOM+V
aaXUpb4ZKausOfNSVN42XtAfRQHrd5OzUQgFWuPRc2RfLHz8P4gWcMQx3jRdtky6
dhHU3bk69xmYnwrhlLuyCwdd9/nrk6ntX+W0f66Z2k6O4pCWoVvb/fLbnJ8UZ2zX
Ox/kCwbQiyPXTL/T3K+wvZ1wbnuw1aLWYCmpCrIblpvxRVj2RubeHIlRtVAnTvJN
i3c0GIlOtbkNLXvXnFkW4S8nzPhlxmFnFa4W+Kc7yxp8T4WG+KhItT0Y+fp5cf2X
QMGp2T9HLfAPN/+UYDt8WdT3cdITPVtP/Kf4fvVezUDlky6Ww7vo4NwdN48e+M4t
GT8X+5KPD42dEMsvHy9y91+eeiCJWREq0I9t7WNKIxk2Dtw9SbNNFBw+RkIHDBqb
CCkNolMAaT9Aiuwz6YIM/16lR1yz6rvM9B5Jf0Kvo6kYljYd45waEWZM1Wy0AGZg
ZAJXU5VICUtN1aVlcPzM5VG2yt0zvxSDw3gPlG6vSIrgr4YFMoni3m2MHPZ1Ysil
78IEbFPhpnoyNk/z/nST0HmUWP4ipXHzU6EkgNKRIJfF9GAuurgYwDkJt7VDEqcD
esX38ytgA9Ui5XoIOVesgikQiuzk8O5HtL30krOsVqUFe1xpw7ribDG5FoLXWIB9
g29kk3OSqXMIB737qKMu71weJCtZnAQV40rfLSDVLarRclzQopXR58QeThFQZFLP
0pvi8JkryVlE6ObPlr+drSjWZHqRmXyLKBOyRDp0KfvK6Q1aMHAJD4Bo+lPNLeVi
jkEHozKWrilgx5lTKRXKP4aMCv1Q1g6Bnvh9+yIqXI6yAGdndS3kFaGKXpaK5vLs
WgW0xar2eQ2jd2f7p2YzZ9fqg+jgkkcF3BRMSntvbKtu/BajAm6v1SHj9zJSKWzd
WfLY9NGzhvhCwdc23lYxtk1y/wNNQqRcaPPQgE2lpOZowEW8Yr43eK8HXvVpaGxR
w0cwvLPN71LesXaBSG7UtXh4RQbPgZQgNaFvs1GOXg6TpAuF9POFNmbTpYEMjJks
VYef+Xu7EUy7qOnhfjjimU7nQWpx9HUD+uUg/5LvpdY69NZzaFwPCvWjweWrR8UG
dnx6uMGoY1mNaCPEFGYj+2TBg3dEJhxNKJIQyenQlj2qY40bNvZjopPv4uCpsg36
7OV8I8L3JtqL9e3ILge1iG/cL2gxRkd3ZcySY5HUYEWfzKVV5azskp5zERs3P3ma
wRhaHOE+8q5PFm3YiLurPelXzWSDtlctIAQj8QjQz7Pi1PHVD5pltmr1vJ0GyAlb
NOaAPkYVvi9EPL3wQvVsigSrbEjCpAwyGKnfWb3yMO5tFUUQM4D1V6s+TgNqGNmO
jj6YeOhlbXkoIhrVsFaTbd74Z6eRQ7+m9JmHuQ4Ex26Vew4klq/gkf6dtHEY6fRS
OJbEAqyOb4GtKrXfAX+2hqTvqLrnjtoZWYAYN4wG9vIS7iesAviIK5Yvw5nuYPZB
iNywxrTKUZ96dw1EaRCq76MRtEVZyTB8YJUfBH8eIVM3sy01w95sUo0P6nMNlEnL
NWeGSGhJ/OSLXASnn+Zdiv7Xfv3CaLqRG1o8JjpQVq9wACbDwlpKTM47RYBOr4UQ
s7MWdsvsk7CtKTOIJgEeKf0fhYOeOtKrmH7yYP2RrGbtI0Nd+LQ/aYttTGkFEbAI
XBKQA5DK0j9mDOwK24Z3UJSnA0VncOVLL9EXSYg6Pv63nasXtUe24lGQdEzfaCgy
hzAuOVd/1kkPKqLYU3PM2gqEnIlAKQIFKhkIwUKl2GDeSFoGFSnUgHTnmf+qpg+x
yHIQ4eMI8tsdtaydJc9sxgv8rfyqIpiDZ8A7IpJAE12t5aM1EjKVjyfCome/8fbz
tT3O/2vkgkc5IOPcIZ50AIFvlHIuUh1h+N2NtC+kSlhniYQMJ0v86WQ9f1gRLwnG
BmzC/oQ+gbdifnOu/dl3v7t2WyhImJBN10mapbnc+pW2SDLtn0G+YpZhk8zA22h4
Ibc0BsYywkF00epxNukvbKR7tRRQIsojfurT+cTpy1V4D2OZJlxYrS8TB5zGWxeJ
gaKqjKFN+ZNVi06k/K8L/85AV8Zmxo8+e8hv83exWEMQguO+zML+PrSnKsbJbW5N
KF06tybPt4QkJyMbna3sWTzpJLdnFl2M0DJUjwKA73AMWW9dJObQLcikLOvaQMWo
ywxQje0wzTYbUUUmcYHn6ztNtXWO6a5sOIxVq3kzGLQ7DdI8OXExSoyBCNaqHDwE
FHA+Hp4OljTNe9zkeyniqT6pfD0QM2i4q6PzXQD+N3doNjJzdt/H/cJg+w+IM4qj
FXOYJbo35mZGRsvakkbnqwAKBAQm2QX7EcOH1ucBsg+882i+ij/9+jc6fneqmw6H
AUC8DJenL6gZZ9rInoX8uqDq/ZUcu+1Kk1Gjcgt3QY4Lh6EElr2XZJkD7dmUdYI4
qiYyZJS9a7G6zHyr2j15RXJhI4h/Itq8yULJA524xjBfq4UU+AVKK2vF3Ep2Rnjp
YHLJz+zv51ucAUW3ky+Y5L0OsoMLd88CpcY7W1nBWf4rWV9oW4YId6wmV0lfhxeM
g0IkIMS9XmF2Bu/tQAlz/LW5RBXGU0c/jZxEERCnKCf4pUGmEdOcUA3ra832YYtf
i7sqyahEhc0oUCLLwKSMhAiK/PS8IraUaaxx8FBYzqtFpO1NuWzlKbz+x7K+YVIY
QNXbDxIf+VgDv961tr0ro9qyHAp1M6MhBmMfTqNaKh+Mepdb0/KffSd4Zh0QbVfs
tjKK/jsaM0JPUU8Wgybq/wrwILzSXKnBOmfzsaNhDL2GTrmLgQoWKCHGH/wpOpAh
QBmabRHo8I2pKwx+caoEr2G6x4GwO0QfCVl/VsfbevmQPSd4qBn/nqibZHbH9+di
zq+4y38hHmzfnF0xGiM21y5PhxFyjMZyG/MF4/nZm3QkNWi/ZiMSsUBG7QZ4D0F1
cIFeXXnR+SGQpL36xHFVuaP132jzipRHbTm/yDWXnIsRVrpvy95f+kU24B5Jnknt
SywAAPt8UyvTHKIJqxfLaTC7/DPkLBFnt385fB+s2reB53hOo16L8lZjqYUe01x9
bU8RmrDkMKwA0pHPK+dKQF1RKeSqxLa56O3cVwWgTL6zMeARZyPuPwTZj5UDGweb
/q/sGGn+GaobPYK0v+lLd4+146orjU0c6Zh/Hfq3mvEg1XJdmgS9qxVnqh9n0oFU
LHe62KHPvCzPmqGYaPqYu3WScxoRrE0r5bNgqAd/TvOM/SzghRSOO2OI9zYGdIaK
8eF4QGws4TCymCXg0VjsR0a075ZWFH8bo5pkWLfT7fPLPfZOei2u0KLgy6FY9Nx5
5tKKzwbhcb8XCWpgEEwNfDx8RsT5+QZ32rHmzzTEHFgNCe2XjgV4bCYc/fG84dx8
RmRdSBrsaC9UPpALC8bOjGYziXH+DxnUdt/6uOKOWwDFe3z5lnICklevTEhVdjT7
0a+iH1+acQXPaaj4Ms0iFdjMdaZGovEEsUtAs454VPklwq8HnTo02zj4i88187Rp
Fu+6/I4SUfbptQZDMXU5Gl6nc8MjjczUE/9ZKHnJzuNrWhoRKM1aUs/SImLfyD8F
QYrOqUZNtCxYeMLEfnBzMv5PhM4OzgGEPIjIUxaa542OIjJQbVRNAjnHXEdq/xxr
A1re1Xu1N3qO0BbfU6liFng0IJDvNJF4292As9g+Ch84chTbp2++TLr57hz9XuXN
cPFLB5TP/XmVMBjPPS8kkdDQYV5FdX5hCWupnhT5N2lOGpnvKcUucQ3p7intxPp+
PYsKEy4u2QTITU1lfLpbDtdXYLYppfvav2OSxAH/EhS3+HM4EUje3al90O2hjMpE
nHbT/OgaHzHZwblXPWidGwLRoo0uLjTgcDWlmiWjaba7bd03lytnQvOjDCF3V8d/
B/NthBxUaXPpQy+YOtpDhGdUQtURLSWk7PSdS6A0/pRO3nUvTCIHU8UlyQSMd6Ik
LUmhh1C1XY/aqmT1Aa2BQ/ZINHjDIeuQOUYcAZsUp7SIdfo1EkUBtwvgoUSiL06s
s8xuonvqOmXDttMYPFOngGU6jp6/FLJDm2jgXd77RxlViUeIaBZosLOa4EyDksEY
iE09Yd9LWfaQBJthA2Gw/4chBV5InecFD1oLjp0FQ23JXDphyAcdlDvcM3mJi/Mo
0cUTzlXIOx9zGU2IlPoJeSGUqavVPbwVA4XRyBMSfQQruGjf60zXNgV7rdel/EDY
NJ1WW2tI+7DR3qUPD7SizP9dbxxfUvAu7PwNW1Nc0RPqiwMYAtzVu8UGEnaQK38Z
Fvq1YONQ6qXKb/Ejf3dj5e5/05P+jrFvHJ1h/5CdT0Y+CcGJBNBSVvFd9hWXz9UH
yW3npc1kkkNt4yZ9IOfH8+XnE3ThO+sFKZtuALyrfPHWVbKeiKarY2kgp3/FzDa/
VZcfHNbtg2uz0k01mWwuyXEtBp9EFCyF3XP8HEi4EdVCkRVf1Z+SHDJV2l+8L51P
AltcsbJ+X++VRZE4TczvSPL55H1G1rzjJ2zpiffwxlXp1biAlzHTAXfDLU8iz6At
o3QJ6GgifPNyqlKSRl24jWyws6z0mUOwB7gI8/HH5Dn9to2BZyb+/JSGhNC2dlpA
XcQuSKYEdandpWvhIu7zRlADzs4WX2RIKwxdy5k+3fTSBxJixw2jNapQ5s//2ceg
dwkAYJbPT/8Jb8sZRe0JyCqmtlTTLt8jC4WK16Tr+1uaptRbVrK0IShFBnvykHkU
7uJLV/K/ehokwiq+9qpakSV8RQUZyvV/bg+FDtRZdzQMVEQO6bB9jQGnNp3fsW9J
YbrOa1Jy0156Kv61cVsHELeuJ8z6MpQuMa1EjyDdy9+tFV+JC0I3gIS1ynCFs1Po
8bwqhk+2e7m2GEP37bGtKkNRH70QCHZvlmp8yjT2kTBjZuur7gAFzLZeLc30Y85m
A8eS2t8mtKM74ugf4FwQdg6+WhrPKZb85KO/gFVFV3aSr06R1upauYOwOOqrgpAC
vA3gxhBf6wX4sZWMX+GCmcEEZ781xyo3xEFIRGIWGLXMmpDlngT4b5E0e8q2j1uS
Dtyxpb+ODIo9YLxzcPAkJH231wMvUksx3UCJnZsKYn9UxXO2ZWyKw1E8zd0jPg/e
DoTvuvuJSIEsWR20I8VWDCXCuRzXA5vSH2CGwbXOQRXA87X+he/8f5CXR98epqxL
UkSaQNDVtVf1MuXn06CVQeaeGPmexF+UNJcGNolJflvyX1ykuRm2pzCroKFGC+xD
/vMNlQk+nVlAaBm8kvQ7WiAd0OtYnhbQiSQUHPH7RLsyuOV1Exknz4xj4/bQK51Y
3XCD3KANFzeW0/2O6zq2ziUyrTtNPyQtB36P8AidvtQrgV4dsRWyrfC++HRtuGWH
E2pY/iKiSDQ7qRcqeUwiSxeu+geA8Se4vjqpg8Rt3WfV2XxVaOhurw7RkrvCtObd
y3X8AImbGijXwOYnUMeea+OXgS+XjGD+MeuacWHYPuVYVwiRN+NzqqwnshbX883r
3nts19iiPPWlXUcTok0r/HMaydZ2/v/yu+2GWI2+ebA3MjbkfE6E48LOD5ZaXDIN
z+RalebWjUtYmG5jCcAZE2/OB2wdyURf9PZLweO2Nc8IZSOiS84EDuBQJpH3bcOl
h5cPm4ToLES4QxIIXAd4H9gFP234eARlTsS4QtnMN0RzQN8/qMESazGvQ5tJ+zeh
4eaN2vQLGEZQM57qeYkUqNcHrFWK7NGweIRH4bp8qJl5RvXOaaL6zyQiXEN/Xx5+
Q7kl9bYOb8heD+bEtcxzmZQkHwjZgWGgEcBQT9lNPCwhbQqIv5MGBdqVSp35kPil
I1UDSBp3mJz6OUOZ8YUxy/IG7ouBgDcFLRk8271n7JM0qEOomhc1FAnfVnmnzfJk
ZwjWiR787Ku8RTjQFPIF8kTsa72hlesi22hxxzyXGjV//q3oU1laRPo715nS3N2A
2e4q0dAilckfreg3+7Eh0KjR8HZiv0vyH+TW+0WHlXXPRh8VN/NK54riKY23yhAL
BcmB/B5/rh5HEWfYpVl/Uq68HUrLApprcqFKMU4yC/DFbu+3MsPdBzL4x1orVTRr
qet3eysvECrGutbkbIPhNC1IU/Op9s2FyZr1MeA/bgTnQIaP5kUVdiTlytXJGO49
PIYYzFyB274TGEfIAY2M7Dwth7jXDd039wQcTCe41m87rBgSlpO9JSXT9B5MbH7v
SQN9IIn9zErPx++vtiKdyZNWHi7UXnK3wuXsBlQ0uzjNisZPkNR2Vglayn1oUr4c
lNo4MKFyGQbXkU2qltB0yh3S88F8cLyqHDicEyNM2K/O63cp86wXaNqDbo2IAov/
cQAsPUPm0xgwhQD/Vw1mMY3AgpI3Jrmp3nizXE3OuoMHBjyrQQmnI8igzgLyrpKh
JTgQw4l3dvr3OBkB5eL3OqaLER+HTVgJCzNquTzcrDG7vrN5foUs7jv5PaIDced/
KNV5HU94q9WBxe2qcB+CnAw/fiMkaDP66v7F9I17szQaYAurmXEQvavgyuWoy4VG
MP8fG7IbKq7Hndm0DLeubliBhh4AFJu1QX5eIfOhR/X2rAFuLR8qAhUO6lRWWrTW
Nx0tmUTvNqANnuaLsIe1AVGVtjdBcMIYaVKP2LpuiSWzlN8Jel2YTBdJdjwy+utp
Evi0PDrfCiROwAlGJUkoVirD+/b94nViHyxviSJ8Lmypnhc/ydcl00QEJM3/GGDz
lkPwNH4bKYw92bpEkwPwN3ovnUX+w8iWWAvc+LyYok2cXXj8jxSWUrWhdGqOQ7Ap
IdQeZ+fVoYh78Xq8C7zzqCNrFBpcbqhVWyJQmoDg6S7sqNKaLitwGs2/iAiHDhq7
bgyfF1lyfuElzosTcv/NpDYuVDhSaWXIkHi+mj6gQZcknt/Zejc2DjCqnX1kRof0
Th7Ntuuuco2jXbLH2uwjZS1ObYrpVwNY9KDvye502FhloD4nR/ezVu75/yw5utJ6
2qsK6vGLtLjzH0H6AESqOlWJo5W2VgTEqIkp71yJZGobQDFrv3Adqqtq5pptE/kN
ncCxaoLlanWcXBJFbkCMDAeJn4KExLhTVW2/eVw3atYJvGvZ/K9ZtwRGGBXdrNTF
z/7n77t7fVc3gwQdWgkiolL6SUIdqoZqhl9XdR7CE7h8EpaIZU0nT6a0F6aPAC+m
2jSTD+eQUm96QtEadfzU505zFrx+Fp2j8et7WlzzwUN+qH6ZXG89sQc8J9Zb42vB
54GsRFWZMMS4aTSq5TLg2ixsvemODJcSCWLkwNqpwOgjShy/ybiWeycSQKEIoLl4
UIIvim+R9DOqD3QWCOmSs7MRQwPe9PRMFI1TgvFDXIF3P+z577yd4BEaOxu1M4yY
qhSqSuFvFssFV9VOJXqP+fJQmYfJ/WEghKaOpbno9oGNdb5TaTrB5qAvDyCvYywx
egeLNe+9J6lmecHA8j0AsfV6exN/kN420JY6Y0OOSaL7waI3I3PlysbuMoUD8Aky
RLgEYr0Wpww2SqLKatJBScrJlqaRIpjPs5ZcyrGMrsw+KnyzYq1lAPTgZJTpTH6G
cwcHKrAwJs65+q3Qva6ZTVypf+y/tTaL+jeX0DR73MU+bz/FbimZ4lbm/ZrIhNV3
sUqxSC79I0PnreR6gkuRa6ldmbrVPW4C39PbdN9zm8WDNoccenCxTdh9vvBtDa5F
iDiCUl+fZBnsIp/kwygW1trHSBjjw5Hp5VHyrP3i7e7VZpiVwt4YaW5C/H+06l1e
FeW87iAGS/2JQDVVdmzqyVQ9CyGE7M0gPbA3GmuWuT5d+cvr4fvurKL6wH77BpDf
nRq/9uPazz6sl45HxNtBvkfptqH6JnLphiSVAId3PE1om+M9m1BePUrsRF3ujRwg
7WrcjXVjhQW9Rw+5QHiQUaBE/S3BrwQagWUp4GHqOf6ViHMZ1YJZDLsehqijxpeY
wFX6Gt1qcMI2x+P0YzthwBYFrefmUfeVZOcin/be4v+KLmHpyeOhyKS41djGn5rV
VNUUq0wv44kKckHXIYB1IjOUx68a4gICDf7Yw9nJ5aG9gsto+UEZsmpVmxCpvYO2
/fcuyaXX0pLZs8wiXgyST8W7UWbZVeV/cnC/KQKoUHeE9zD5bcIBWwRVaddQmoEN
J3DhYNF2j0NPmc99mf1ojEEcGtv3aD3KxmNDcE1U+DOoftGuJf3bMMy+56qFix26
HPlqzSB3vqU/7oQW2XAMRM5OIRoWkr911Zl7QbG1uFmGmE+No5P43Dgp01fVv5cl
LSr8Rmhxm6M5I1DGe1nhl3WQpTS2wAgV4RRghcjABPQqqX9NSl9vFv6R3yWykknA
/hsJWWC5JUnWudKa/0//hx7aAdCErRAokYhkm3B/l+DdqPxaaNS522S28dsdCOv6
7PdRbYincx2rTGDxpaQ2C37dLYogfe0jHMY2kiSMl6AWbdrZOn3aRD/WvNY71edq
//LW2yON0Bgsp7nfVgJ5f0chdetG3Vfb3yYo0oVa/HdjqmQHyq3N5IETHnHfCqZe
4DXopi43gsRy7k9vFHatBn0a61hTrcjPYQ9TfXkp2gl2iayQgyk/whPT1g7CAthb
0nu7bQW4rK9pYbVHUbq1gUGs4uI9QjI2QntpPt8dGxrXujucvUtbjauMgh8C+2qw
ajAibaZvzOriJ6Qq3F6zdpSNAM64C56bC7Q2Bq1yfRh68BOwXOKTys3xICQYQGAM
9Mu6tE9xSvSR1HATomq0H7mb09AKJuRhyYphjJN2289RqAooxAAJJ/hBi6Jgp+uO
IYGHfwuU7wTdhNH5YHuY4gLL3BYnvXHqWkGBd9zqY32FZ62TATmXiGR7e0PCzvk9
gPikoCqSWgQWZnMrW1hXktiJhVmEuOLaWRWBGdzBKiPXH6HY/aD03RVg9e6gNz2f
15S4vwv8XlubiqjlK+40OtffORJ8xHhcPqjzUVj5hdjDBDnko0GYuKp/bz75qBkw
L5bs6RtSWbUwAqTPHR09/EIc0oZgVCYuH7JnAAMGm2kWg6ZsPsRsOnaSceJ3yEw7
FicAQFcq1xHTRdkBHvnN5mHGKLpghlvgH3ycE/iSaDB030tMizAYcN0aPSsJn1cA
mGiE7DpG3Y8Z6FhmMt0loLOB4roCKtIhoyaVPIpa1V1LUTN1QQUbxgg4yY3EbcUb
JBSy3gBJw9E8DJPpSn3MyjujzRIE4MBhSwoKVTB/ALP27+eYuzlGPzEnlxotYFQL
PktzEcdv63uO+yuuKFPWB1gGPd06xbaTvb6ZAO8hSud1O+ptm8h5NC197IZmXLkO
w/QQT/0k9euygLJtzOoY7yCuM3pjpku8mleWI/+ggwEd+liMl/gCjV99cTaMCDYx
R22EentLhXjM8uFusDM+mMWIJs4zOJKh6ihmZwa/UQekhIJa8MMaiS8KZw97TjbD
eLHfYdRsjmi8K0Bj0lJcJc3nuOONEsFDwpr++4V/Jpwuv1fCRstPeJ2O+CdPJWSC
1KJPRYfipgOKr6y1zH+4LRJDXq+05eyALsTKFTZpbmUvLXGXQlNg4qFhUU3atAiT
8M7ZUTydYLFchK31T5NK0RhmqfcUmOaSrcrIAeQAHUGdrDQOETtJHOu65ZBdeRPu
Z2R4W4zovdN5rQptj54D+gTtkZMoewYHl2qxBHdMdBZ4DlwhgK3uo7W+CrNq2mH0
ySFg2ut41mNWplLx6NYmaI2GoQsRaZBrOPp6o1kgt3se1t9ndeJ+9g63shxGnWUI
gBzHtZDGDBy7QMn76XlimznmjZY3Hu5agqzuU3uvvSJW5nlSoERmNdCuK6zwVnJM
hnzqWPuHlPuyYEzw3RwxRDnoXclIHjVYvCHHLHCdn4F64z2rNu9YtDtFXPTFjB6P
sLPIJ6Pqinl3sVJlgzBOc+GKAvoO8TKl1n6GLLLZ40BuJA70K1yTuDEnpjuIyhUb
tu/aOUSliUek2dOrmdLN3SgdTFda0/UXChruHeqT5OYhQ0IOHMBdM3eUR4wNPhta
HDUF3envPWUPhPHIPqzuTFbahClOyar8IjuvWGJwvgGllv3VOOYYitcJU880WB4t
fB6MvQlCBnkGvgDQ7snFtaYR0SNtJu+XnhM5jXAti4MGhe/cnNByv06I8CDsUUur
DRgWwihvUpi0nwAcPWroCIW4JdPC3+LKElu9EiGFQRt9xdcLQc7qOLQxIByYSB9R
NE5mGNLa2OPy1wC9cuDAmnEk7hhByiY9Rit/cOOAPyGR+J1l+dpuKQirqb/KIlbm
lbmvX059vPV2SrlX7LTrrUTP1wD/kLIGo0s8il+VoIFXh/F68f+66siReTjPAREu
u2uy9ffffXlcD6grOqAqUaxD/MEc2baGgNpX5RC4phQOxSvOKYvD9+wXF/havt3C
yEOo8Oo+FbY6dqgsjZ3ZNA09Ep6Zh9byrCk4q+TbBUFAXSuYj8caDd6RG/VsHFcR
Nc+UJoiEsZIDVC8CfzU353J2bhUvnus09IZ4LmToeiov8cO7bX4oZFIEUaQgqDXU
2HCFDirHQG8ecZ8GHvJYdijB5zXwZrvXiAUIPipbPqwxMAHQGKIpk8adQaVZrc4v
F6zSQxSCifmus7JQHXR65R5GzgBJdnaINxMDZzmCLNO0BnuIwXJk9jDChx8yZOKX
zFpB6MsUPV8LaaqFTTG+g2W54zUA90UoL0nsE+7ntrnu+14UIXRjYCvab46eiZjR
B/J7we/dmOHge14OdFe+xwy6i12RECIMZuYFTs0E3Cc0Wy9B/c6P5hcWyjunhjwR
Em1/VigK9uFEellNr9HungBC9NmUorWtIz8VYE7CGEOWjOptrR6RBt7EZ5p6a8jY
GglRsS4By5lI012TEUuMXPp73qdRqt7ZuFKrnZ2eLBE0NQvNj5c3q5Eww0SD5dzE
gNm6+2GUP2Wh96ElOg//xx1vdDXY2mfV/5iRIN9K9/h+kTXrR+l6wiQi5zn0K/rl
mmxXcqhnXpN13zelaz95aJWlr/5QtC3OuOGT4xKX8G+rtrubD0oY8O/agIaAYma7
78Z81HnkhW153M+OdT5KxGi4EkNFG5VUUKN3IfGJDQa/Hdt/mGYy3Xryn4BRg7ai
J7XYUFF8uHwkmdAjvpQfT6b/sWogSHAku6xHjsNsgwkmC5rPkZWhIQk00qWPVnAt
9C4Ag0KL1poeovuEq+HcSAyWvxeqHzjdl1dwDi5+zLNMY0Fze06K/UO+HV1oiPGl
QqUALdSZzi/PXDvA25JwQI9OzG50voQdGUDtLQM4v9nt/vMH+qAtAiorYElAgOCD
R6i3sacG2BKmmRL4HOI4OSt9aXTpfMP7Qt6DvKfRolrbBf1XiVHhQ0gGW68VGxRE
U3N8qkrRG/Mnrz82oKIRoaM83pfGcMz7Mexq7YWg8z3+Pr48JrXHjGfcs/buCc8C
PuTCjzXL7gzc/NdjLYMb12JyiRYbfrj4ig8TInhD7Crg9UwZAaAe5Aeid04hf2lE
tRFlzt9vBrZsZzctWPZRJlHITGH5ATz5QNxaRiXL7L5BIWrdcj9xo7oGxucSNsrb
2dSwq/Hb2BkCkUaLuUg4nBosgsvPG1qpot3Z7ilTePU3OcUL2V3miO6VGwefad+W
xhGoJNmlTJ8rR/SV43xtyJ3v2By1+kLIFPkm0RkBkYM63Lncw9TpYcupstiLcO2q
HQgqp4XQuzBSi+qzVr9q38qhhyWCtpGrYen3FvdjQA797Jd2tET4fCBJXB6xDh7c
jLwNEP1h1fWMsZvJzDxvVMlFiRUSXuPANhdzS1S/yMq9VmxV0uuRkgD6JAQ1YtKS
G/4Nb3KZzCXZhbMgCXpORYYIhwUrT4U5p/Oc/aNioxT8hDRZG+9KPu4+yT4xzitN
I9S4Hz1NPWLbWvNN1TM1zKGZn8fV0rJOeuUXx5tCiEVsoFLLLH2GM5OeIw6juvaC
Zcb/DKaYIPJR0nCQSGKYeuQbKXmSCTmfXQgo2jLGu+EMSKnVGMH3Y1PbuJrshrsg
cXOC4O3bHE5b6l1zayl4VJBqFmmz/2/pm/wU6aGcRgFDUguGYBt1k6AeAYH8Ty3Q
ZdIvuXpeifcdkQiloV0GHxb9bx4YsiFdrBJ5ZAwxTvjdou6kOGn86p8puc3CS7+G
UDQQ1Fni7bt8WWideSBU3VZ9MiomFIAyYZ7RwEDOKToJmdnUhRYrtEsyPycW8W1y
Wx7a1kvVvi6x5ozHhQm0BupKJbyS9hyApmYYmIHaXaMtI6ZTgeh7O90RGv56yX9U
XzSXY2l0W6kRzuJN6xPOhgU7kZjzWPv+ww8s4/lYt/e+EQgEDr2IU5JII/tPPup5
SVTALNbb1jnRHEvwpQFen1zYjij8UapsK3Fhcbp3O1xwtng9Svvvypw2Xus5A6ni
kRCgwQmotJoHUDvPxcUw+HUzza2SMU4AG/FYqVrcU6luYMDZ58THFSiG5oFTqKXc
9/sdNWPd8cVSiEOi7V5JZ4Nj23xCjj1n+VqvYPVqA2XiAHbkSTVPIPp7OQAbTPN6
U6uvhaewzF6lXg1T07XyVQFbN7QyS8C1k27thlZ+3a8Zsp3Sqz29Fkus18lqnZ4h
pGS/vZ6zGk8r0xbeira0zdRCCJ77owkYRXf0ATVKKu+KNlWUQm14VM6ePl/XEvL9
fFrhI4CGlHtyEWtOF5xc87vTjad9qBdtS2D9jX3PAd44Bf2KEv6odckuijB3BcyB
a6LcUpmjQzrnXYJ6fIQgvQYG2YMCGiuceDwCSL2vGrV+B9F9ivHtokFNWzfjlRR/
Xl1Lm+vngJEm1Sp9Ppw7weV8ocwZXU36Dx0zvhc7pccX7aePw4IKAScHnKHJw2s7
NVDciNHUMiDBY2xmEopmgUiSKw2WDJeOG3V+lzLpNqQ0dnBuWJmxyr/QA2jU+c7c
yOQv9e6xs+Tp3UDIXGMZD0Z7fFHzAogM9KbQKcQzVPWBCHOuaE6eKQBf2WugVaBN
yR0miHgpUseNSaFhijYccjKClzUv2cCLSt6Dj2YKl48UZXVlkpYF8bnPVtNSOLAA
8YwUS7osntRfM35mj8my8N7wqmba834KOU6pF/UfQhtjbNvkmdGnU6qDgngo3niW
8U7hmgtzWM6ulh3ZO7qbTGoJZkw83ExMHkV66hursXqezgo2i1XIpBa2gACixW4I
pmZrexwHV6A8U5iLO4CKrtc01YkY7fN+v2ODE5fGejo6jEN+FuPoyIpgrZjZnEaC
mwb01gfj6dmDDvvtb+X7Cz0WbAbC1i7nJTbQwEEph6cFQwIUtaLDwXZBX9ijCYz4
GEq4umY3/6PWZUboR8bj46XodL/xyPtMNmXKjJPq1FT8m9ETCrOuy8+y8zHDfCxU
+Nxd9uScRm0FG9vcBOGwhK29X8Ms1UQ37jmmhUqXVdTbVLyZbcu5HdKefH/SSPFP
+L0VBTAonqqnqHUJhjhc0BKXc2DN+8jhZ7DD6ZxqmeF1oJwGNluJxOuffv+yZXX4
GhdxwHkPZzPy0xixKGQXs7WxOX40WvDrD6vuGxmQopyg4l6sICtWjrwGrNNGktAs
AZXwly6iaAM28IEddoSLYlAbKb+xg3FzG4lEIg6L5AhmAH7tdBLyxF4JUi85t9Hf
XeVSSAwT1s78OdgtJ3FYXc5q4eKbFH26+dKm46x2IQbNi1hAECJyXzJldCMqw6d2
FL5C9Z4QcEzMVY4p3hVVxbzpGBrXN9qZ2hICW8Q1oqFftTfW9DtAPX9+TeTD42xy
kQNgL9BQ7NEALLuzsmptc2epUnIRghcp6rRr/6zTPfuN8QUJKOp4FHCRVDPotg9C
rL7Q727wcHrw7x6Nh+LzG9M2Gq/duRdF8TMxJWdY5KuBWouP6uBzWRjVnIAYaHCC
91wZ05uDZl7ENHELFqg9/6bRPzdwywZtjaT/HwVL52XEmElXlZ7naOCkhU6CJ91L
f90fD91kHSOczn+jDdsmqWPWjRHkyeRFOoyytfLMwId0UhPcbw6fm8anmfIFL2yk
14f62Vxljg61GBYKj/Rn3UcCB0JoE15TV/zK/ymrJnlfw1ZG59bHsJuohVo9Bgc0
GJzA1n1PO87VGVZ0fuKEiAZar+iFwciDDWWevFVfIJ1bvYtJZQqC6E50J1QdNdIE
UCP4aAenKPPZeXzFz/ugHHIMPRNAcke6axN5L+3TN4uWM2ywp289PQdY9zDNQyyb
dTmMAuEiSvhz9Zrxq9WKthOjTvUZa+AAoE0kucNJaWPMMi1szObI0uXFfJTv1CcQ
6JB8s1cWe/yhNRkCD+GsSfK+nlAJAAy+xL8SqjLW1oQ3L8Pd5AHj/smYq0+iosbL
jJqU6daI4Zzuvu0DYU5SbONJI5CpIR57GXbm6pb5buEkKMb6pNyJSXykl+it8nhI
JHNgEWlpn4r9bQilf2GzNmMUKO/PIg9nNlg0kbnPiM5FiyWM5Jo2CG8LoxjIaXGH
eJgs+CZMaeGn8CxU2Dz0kQe/t9wPRtpfNTq3OsxGwFAvPO3Jo0T3bAjpcTnUs0EF
9plIbDrk73BVjU4DegE99dB5ih+Jf1CuL1PuwkeQY6GiYMhs+Y8xWblw/wgA73ME
YM0DlDM5RFTXNAArHWSYI+N77vaHd2KyA5BeyOVy824EpdHuvlwmAZiTCG+7YZKK
Xa5aFw/V4FY1PXv+r9eekhUvBnwx5lp+hm8r4PH2KKRjKCawOiQRl6kPtz/zwQxO
UV5/NwXeeCV7iP08uC5rmow+YNgjKksc1rQNn+R6GBCQ6oxoFHM23CGC8Br4QRiq
/v3MmlrHZOb34Vmw7JVhxRuy1PwEtD9/5UTr9wbq3vctSSEYPeDCTsgjEJ+4Psft
lSyfXr3Vktu64mrNElAjfHRTmmvY2rvs2dkYQ6rGSZfGKDflxoma9kginbjBgmI1
WNNVBJGAQvU72a+SED5mflRHnsnNANndIowuEbyhI53L9pf9i+ifTWAB7zv/MiHr
RxdWkzQ7tGCL+ulWE/8BZRnlZPTL8krznjODmUTc0L4VJ4pO17HHuaovrZCcCBOM
2SDyCkh68LOuDR4uaIFToG/Hu2veMz0jpmWMWxyBFkl/1jePDDqhS9WO5qu5z28A
rk1IAKdwAz4wFTy9mGGCPTm7FAo4sP4oKf3uUEGHl+L6mUrekYmWM9pqegqeLvHG
qgbLvLnKfsBrOJzd6isuUbgndy+WJFWt7aCWozUpqGdEDzxIl+AkWqYRwb+dxufH
ETzp8A2ubQepgTUakSi2xWjxSDtbMdrQAN6t0MCiBNiBbj6iXJEFEZSOWyDp/qmH
1f5vQn2IDwDXF3nW9PR1EsxhEHxmAHqXU8Arw+367M81rPAz0a964Kc/hevw6m3M
dw85R8U2geBL/A6Vzd+jxsfi21ks5W6umE3yqrzpnkuhtKP8HwAtgMvSgaUO7ySD
vg8QO80Lwou8l04j/FiT0MMa/RDi0SKJRnt9JS9Nkjmn5e1D55ihBQsWt2ghl3+N
/8cY+kfM50LuvtTFvuHqUSQaRR8056n804q0tOwK1Fya68SHUFHasYzXVB3Iaq7G
3+773a8DKL1tqJwZwI73tqXM6WY+Y8di4nC23EFUlHkowg/iuMDL6jgPp8xwaDba
DT986xwga9SNCQ4X6FIb9eDgkmbNCBjH5dO5XM3zo4nRdD1h+FHsZ8cLFluzuOpl
tqRKch84zO/JtCMvzJ0aRgbZ5kw+gIg04Cf9i4jsNhFPGiRPOYJGk8gacoVzyZPf
KKUOEMGxQBaoRMTha05mWPisOtkL211CPnFxYuNs48p44umZFhGk2cu6gDGeivhs
txEoMlZKVBKUSJR28sa55sHZYzplwujXe/yx+kSrNnZ4BcRZhOMunnu7KGYcJ+4P
Ae24goX1ThYj35ucMg8I8+ZN9hI0wChSkcjVvblpmKNfwFCMj6AHULvUuoS35H4m
2zuHMNU971P+QrpLBYMfzvCZnqOkRX32ouPdaspP3mDafaesMnkDhXdxIFmTeD5x
CXIzBBOsD8jup3r1N1xelBGl60l7u4tA5f+Kv120jOlu2aHLYdZ984xS9NaeXhgM
wuT1u7/DE61E272FAYsZ29uwYFnd1VTb2l8za1Hym66sADN+jdVG3vWb0QAI0jDI
/zE2qEaLKaoVgWZEG0VPq6sCeqt0fmdbp1pgX0aeUPDOGkw6Jc40rOeGjk4usUqU
Zvdz7aAtiRdgaCtU7UBmCWKi8aXd6GsAEd9qOBdzj4IP4rb6mWerx5Q7TKBKaddM
BqNASZRAuVptnJNEp5vSzLs+FE5jM8YOLN8EiASSrW3/YLjP8H4HK8zh3iItXwfv
dpkn2c95XfrrVyOGe77RHtVvscfKB99+WJWjQpwrcUfek7dyGc0sEblybH7/fVtY
+R+vHWlxBfeAQNAk+/jNJOU0tw2GZCl+Nd6U1RGgc+yf1vlIaG65Spf+lR7YAfgc
q5HIVxYtOkT9N3cV3LESf+pnch2pjAmCpcGavgzlAEdO0TBR0Y3wAACKVz0RP8Od
64uRpNLGjSTJCs1MJfvV6UDGrKp0rA2Ks+OTpEyESEZml4XuQkKs1ksl8m9vW0wu
l6oZf8dzqA0doZlnp5h4YM72NnVNv93/S0R/3DRfOvdYd9KDfq5/CQBx6EX1tMHt
pjOq6l7zFrtLKqldNRpoSkOzSP+bJHEj/kUfetuk4yvwn/VG5AQShNEolfG7CuK0
IRZQcacJNtnZ907WmHxsG0hf+B/ralhapR03QCwWrKq+qgB1SQHYaZ2RIDer6QfG
5oa5xYwYVwLYDR2U08qQqYpsPWl5vGzjXgmMarzIVHrTow5Ct9/XRbEYKBe+LGnd
qDue5gmvGzHarwnQCwGCGJ3vLkLa8JgJil63Dvk9zvAGVduVFQpRkEC/Mznwu0MV
HNW2UW3F6K8If1nvkdCV/jGtHGGqMoDsA5H3AoLjhJ7sl0I0OFUS+PY5w4RVu5G4
EN+cjm1NfXlIL0hP8fh8OwhsTnS0I+DJa1+ip9OpWqxylZhuQNr6+GQ9wsVpHraD
+YToC3m4A35zSkeJYTRX4MvDk0SUpOPSpQs2NQjUvwWGy7uWi4rRilFmcI3nSs97
MaPsgd0uQIvJJy1Om9rpejsne0VjVHH+tdomD1e6twuQpiFfFvr5eiLUVOAhGyJ8
bs1PC1pQkezlA9edf4icv83c+apcAIhxgrWWtVugDlIhJ+OOGN8QYgCzbKf9y2QK
RCvmPYvJcWoCGuK/+XAPwBOYAaOid7ViiOVQB3AEtTLj1bIALLSeCR/SnW1vjz8w
x/K0PQwuiQZ+sA6DZY+cJBJk9npjtSJIXUSyO63Qhs67BHF7jk0A2Mfw4hqWZZfP
HABMZn85Yf9OG0uZpQesdN2dQtJI1ABSjCpTPKadGAmpWNHn3PVZXb8sdhNXqXwX
ZxRnTwHH9VwCuUsLrs1Tcj91jnbOo1imTZ4268By0lvPFfrSpX2ARgqET+aFeZKS
DWQrxDA9U9ag8uQsmpElGzuSluNt5sQIzx68NiGcbRQptHEq8QwrUPjlzwrJiup2
3XMH9hkdG5XxJNfXSaTR7/7GHz2oe+d8+EeJID00iR0ImnBpgYjP8QrxGd5O9i+j
xOsAudVLcQKAxcHnMfTwYcMzBQE3hhpWq/xIu8d0zcJ4Kj88N5N7NFRH88FWQCS9
xzlUfZdAYQbrRRnYBp6uGRm71as5VjjrT0Beng+F86ulYZWnTvW6a9CgNcr3Suem
/v3BPxvS8V1p3Y1gS/uJlr++pM0WISVfbGqXtFaLMS/uIRwHjTgkYiuXRneIJPYz
hV9jRuPg3zTMc+ruOwQH5tPnOnW6vBl49DUZtsmmzW8aSf58G+Zqv9peV1c9ATmK
IFEbs7T7mibsgm0qwnJYYmR6Uk0OHjEc8Pj3aCx4FfSv2s/p+2VXkStV/lcbJHJ9
kswgY9rF7fPby91zKAeWrmL8eRk7vc2eRcpxdN7sMPaQCdKW1tDqQvpuy+2nMj61
ZKZeTosl32YpNsPf3EfqXU3Qjo9gyFGzIIN+FX4f33rbi1BTNmKVni+EaX0eNa43
vm6MwmzHNVi7w+3tbsbXuSsaW83L9cL90l15JbZzcK29Vm45do6xso+epSgtikNQ
D4aRDgm09XcqmXSWA6+oGCEfFRjYv8cX2I4Szb+ZhXQ5eu3CyVnyR0i7YDqaDxvi
u+m0ffJax53X1qlq1Hc6k7yxNqQ1rE3jOHgyprBRhHI5AjxXAziRthajyX2Smcyo
m2V96yBQ7Lhs/ldGWMPeIjbwh94B7Sv83NF/yVyOPaB2pvXbitXNEL1LtavR7c/t
vH0KGzI2nzJLM/JgPbCx0iS27RKj/4PRwNzJILcUYDWp65d8K3YTUFNAIjDGmhWK
GnTf1WAOMp8qrMydPbaiAppAFBsBEO9r10BHxJNR9H1toU+fM27fNdG8vBwl1dNP
AkbGGRNv749azQXE28ctpU/EpJ/DqKRF7MoHLTvgBt5wxlOvj44piwCEMlAELN2d
WcrCvkkIUg9Gy3khS3KE7uq10cLWIgY6RMgNSKwJyGeChPQNbtaDyYbJxohzEZ5u
zv5ze9aXRk8xGcVfxL3hx8rOcCrSX6GH4fL2wyXMqSf5g9l0qPhykP6ECd//lDpH
b5Y3Hl35AiJS/PO9Yp6elDiEcZ3bscw3MDXJ39Z2I2VXsakhil24oBA9KjPlGeZK
Ino9bt0ZhAS8GXm1lA+lZCsWYeLL2ET1QmMrW0Mv4skU6pz67a3F1s7SLxjoqrMf
e1XE0rCjGtYv7ctgfm+8z2MbYMqTds66qqCp9JaW8vfPVsnKJksB9Pl0OVk3ewlv
+pwpRtRBmDWWiPy7sdMHaIG0lm5b8DXIs9zaKA1u78w1ScF0Dkh//1XvrKfKGeiG
GzD/4Zd+cp4YaEdjWI0IIR1d7X+BhVRZBYGI+hPiwMvxo9T4TEKBgAWMpUM/HeUd
vbr+VnNG/JmN3p3P17yt13OZTZ81ClH4b0AExX7vqP0JTpBNI3Qus1WBKqTnaomh
TfIj/VNmupjqjl00D+gg3P7iHTom+eEtusHytg7V8ZWrMF7Kwct83qzaKyzgbBw8
HJXPqMQGucbmyF6+qcQLWFYfkatiOIOCRsq0Kpb/FAXmnT3U+NGhRJsyTko5cTsF
n2Mfz45TkZ7vaW/YFbd5G/8mcH7/73uz8HhiuYYF4Yre+ZYfWQeStFjZv6KaGm8W
JzvVp9mOkgS5RmpHkdFxvVnQH1CeV4ybpdCTKQaI3CRaiK5CAGw+C1iKjS709SrA
9AunIILbpWG3JXqHjH/z8Fo3elkf9HTmF/tq+U7WyaiRuPVLMgFAhdv/57Cum4Hc
bDrJsVIHKvmFy3jNFAhoIklyx7Psq0yWL5/2fGjLvaz6cqvlsTTvCrCpfGIjd7+U
ERSp5KPRuyOI3Df/meIvfcKNI6edmu8dbXSIgsaIO80c0WLohCsts2NGAXy2apdH
7pLBfycnFWDRMXJHrEkgnhfiSroJpr1tMspD4d0u4Jx5+zUCR4BKOiukcVVkdpuG
Px5wFvfDE8nRAB37j2oO5RGK7dWP7Oj+vzB3LSoVRxX9HHNMKEWndYMsEOcaLPkO
7bhdukPAsmKyczE9tY9aXOTzbE4njS20dskZz95cNktCBSayCnJ/Jn7JDP5RjK/l
eR/eY0i4ZfM4L7RNoC/mmE+luEwcWf02t+yvWfjRtnid49xlSyw/jrArRg1BSreX
KlDgP1//kyozht4cetae6VhUZZD6SsH8draSPXj9GaR+zb2h+G/PmA7eN+qUXUs+
2XoHWna7qY3RrGQfBc5JGwTTrOfkd02LqVzv9sxsdo0+ZBwU/10ao3BsTHuS35QW
u6OXXTFtyzs8ENkb1WF9ivW74VPC1Fk33x5rE0yxa/Zv0+mbYrvNKAycdwy+HTfQ
CzALF8No0kH7mwSI5pgBJ4wyio1JC8l5HKPk/Lm+M1oSvozVqw4MJ9fWo79TzOk7
R2eZAjttTDrclwesapsPTkw1TCQa9V7VJwL1I8jFfkTrugHSWZQhB97vvsKCME4Z
neIZMZ9zvMjxI4tBGOkgQBSE8ghHQH7zmjpdpZXHJkZLxMLrWuqef39GMER/Dwvc
KHE1CSDGcK7hoCs4LkLCr4aAGhLyyqzFnqOm26IOffZtoS+vtTkmh804eCVVWMIu
lBqnG9Be93fTeSFu2PxzfdjYtFY22ra7NzLOKhRR09lJYgKiWKYWcIUVmpi0Cq3H
MWZUFH2WyhQeXmelVlKaIWZipMyr/vkReI4jDnqZaSJdspfroAT7BYWnQxj+ohVb
5dJysa1GpoAf8fFG+mEFyNH0emGrbT8WJndfEEsLy/iPubmu0XsnSPQomc2SeA+2
VQ2WxpWBXIPDffZVgFPCZsGLXHJuefuNjUz5K9z/26CueJQi/A3no+tKXrO9Xvxl
BqJwFBJvugvrC7E/fALDtbaobro0H81wy9GWLpmFUzoiGY2+yaamwIv/MiIPA0A3
9GDEs9anuzxA7T58nF+QAnw7Djz3o1ddan7hegdcEwy280NdHM/fxEoDoT1nZMZ0
CU7IDcdFoQS9KifsZtyNUXnCtjZMV54k/v+Kfv/wh8gnPm144KYD2QqV/T20DbnG
SwkwF9+e78lg8raitIPwMQJfzdFiNxRurgtmVUDLbCS17lVRkQ+5Ylnge+LMR5hj
b7IMYuiE8i/odt6Xl/kMYlo0YyytmsaKXb7gXxaGO1rkE3GosxKbHIG6vcpvM4WF
VXoCKcAyvq/6XlaFpaox4v/5gnqEzqXvGBslWhBXep2P8+vy6CCUPMlxQ0v6H9mk
JueHu/EJlinG6a4a77mnxPYN4Ya7+H7rFfnPudGkRB7rR1uI4mfQrE3Pl9GEasI5
vURiJ903e2/uc3g3FvQjukvZkmxvwhON4ro2jRLG4oQhx36ZhNWtOsviNmA8Wpom
wJ4k+R3L/z4q59jF9xASS2WBpKno1MAtxH5iUowTnNZY92eXpJ/ux3/obHs7ha76
lXo29aM6d8NyPn3ossb3ilYAzXpQUExsVcx7vEOm7J0fTjUdaSjoKRj3zQ4QNvKL
+j6oDmjHNbpAT2E+oPmQZRQ+0zreVZ2t6MzMIjc1N4h8RKiMqIT/vE1P+/VVMoMD
f8j40D0Cz552TGx1c/C4+0qTtgrIdkHdf8+BYX4WqSRxvjakKZhBLQCXAQx4Kkj6
YxQC9ez5/EXQnfNGnHYtDKWCs/Q0hfLhv6OhvW0NperRItpKVPdUsl3VC59xN13J
onhYsoWAWdjpZgopGXhLxkmGavrPO8mWHvQzr66/xtK32gz8SI15caU8zuVXiYix
9j+nk/hXFE58wvwJTGJNt2zVzH/Z/FO2gMQKJr6JRIZU2HyNX8DWqwyctJeIgMdn
8g1tJXkb5kwDw5tii74E0hxteHB36wRFL23D8NRyT3vmhdLv+V7oHq2xkL21i1d/
cCCGfrTjDZ4hCzk7D6ckj6THKTyudiJ3Oo4nIHGHqvPQH9ubsy2AKiamZNGCYjzQ
l0kbxWfffNi7HRkgTDm/rAyXY+7IzKVv9armlyN5cgcLq5TvJ+peNPilZxpyJLig
qf3XAb5aBZH4vf0DWSdXNJzcXuPqavD6Uyob37heVesT+AkQLV4qsepMpG4h06EZ
xflKULF2qQnyNlbbYY26AVGUwZbpJT4mj3U+RyhfJVNaSWnNkvSuSDkpSJQrmZkI
wujPJn1Yv/+Q9HPObj7wqwimFA2i/LofQS47CgEwtzVKbA++nfkoP4eHX+W6IPED
+SAEdgXwl5dep3dszpJk9mnipEAtEbzsXiiGElbys5AC4n9lvqa1csEkkBvzD19W
0/pS4Dy40NRyG3rLQa+miKEp3e9e0MXrdyNv/3WuRfjM49RKJQ4sLvDB46J/DXDF
47brbch2Lxg4wNFQjVkM6Qmm+bunvdztHecWqJks0/N0DThOxa8K+f8a2FnWt8xZ
uSOPOw088Y6/HG4N7hisbM+WGJ4EwqUpNYnL0SXTammGVTT2AAfeYimR/MHvP1em
faeC6RygMTYOfFQlmQkd1i+OiCacIbguPXI2zwHxDawBGeA35zm2ZOXG3OdWKYsg
xXYWax6uWhCH3SaOppH6ufWiq0StzaU9iHgyE4gEFgd5BLZux7mB8IB9armqKLVO
4rADMvBYvBZF7m6j4PR9mGGdWbRnynVBOjTcUyQ0fLiYKoRwyVD6VrCGcn8txAK3
X3v826OUg1n/F1UKRMA8IuSO0nLHyJ/LOMLnFKuK9h2gB4D9L+C3GCXllMIFvEYy
BYvPPkP9r3f7O0tySpHf/G8mkvRZb0ovNJz8Bz0hKoG0QRUmDQ67NfkMXIgCxwDs
wi5b/qY2zVwh8WokD/YEdgoiQJSNku+mdeEz7woIb3QA46mBTwFx3of0OU7sfyJU
kKVnT87qH3cHCfaogV4eRVHPwRJYjS8gVmLGUG5NN6/tuCcEiSp6XI52MvE5+cmp
iawk/P1CSIWrpxk8VMwNl+uBp1UXFhTTCX5RYLt4Xqz+Stfr7cOep8H9V94nrlYn
qlw92knozvojqVGN0x5in590sK0WecUZrpd6/2+CeDYmICF2dsQPj59BNk718FPE
6opQIcpqB27UrL4GEhgY9jocZ2KrQY2Ev0rKj1dNEX+lJPdqOX94EvUYehYanCy1
xmruvMOfpDIYvAcAie9DiO9R0vVedjNopf+gZPcD3X6KlWHL6ZX37roJ0Rld257J
3LTaFsuKAGxcPfE1NATwK6X5Um3k3uevcDOr+ciD7zFxbblPxvkgqyRcMLPJ+nj+
qdZolCYnbGxlM2KMT+ofc8t0ZzurmhdXjyo8w6hnO5EChIWe4DvWykcf5O6PH4ZG
d/DnCHvPvIVu4WozCWECTESvKXCgEacGffNApAUKYrNfKwPFNJvDKsM4lmxQIZcJ
nhkf0q+OxOf3m2csnViDy+l7/nLdZjKIE8rMiSEmKhsCugQ+DGpqT7LywvgNCbz5
IS3dJKLNcJ3X75a22yZ6ocPSecUe4s5ZZcnfZaZs7WWPB+6L9aJlcRVUL9eIQqBt
sTeZ3oUhtPuF02yfvRV4zBu8GajnxDCOp+/XQSDuGr4XOQYjHt6zEauDl239nhox
SOkmXhHzjZPLh7WVenjJtjASTGJRIZWFfkhwMLkACLz1wuLc++aPtxwI+aZF5781
46EfFr7SyuhsshGIjIlKdw4r1n4iVj9Upd6LBHycObI9CU1UBh367UjPeGq3trcf
2ncsJfeSpCWoAiVpiSnmB2kJUxOudi+kODOlw6u0SoQjD/lhq1fyPOW/vddKC5/r
CAMOgBNrKt0LEsgkMzSZPWmVTbQPWD7U8uJP1tv7cuTgjtLkhaSrQTdeARCZvWch
z/iYSjcVq2bucei0iuS+heRZbZhGvu7Slu0A8rmkbi4CRkqXL1p6KfWotYnrfJpT
ubhyuJ2hxAQhSmUy7jSrYISs2wv4LaTY9AfExixeV9q8JFZhidYws2pWRWH9Iy4V
cb0rwIdRdmSFHx0A+xxHK3n5+ZUnsjDIUdqICYVwRCucCkG50LIvBV4nuLIEeaXQ
6Th/8qGMP9peObd7TEJhHTEaYq5fCKL8wY3vk0nONlVL6ElHpwRX10Gsy/B5iEwU
QMYRVRAjXnfYzxqoswSncByE1Z39zvM31XU4QDmYN7W6dgynSm0PM4Rd6L0jy3Zl
i16XYSZG8x7FSddz8acpESw8WHzH4T620bNzvhNp3b2SXksl/dvIpybjcHFQgujI
jpJ9QMJKtULkRMmV9rZfHdvcJT710sKpobGOChtCoGri0O2uH0CwxN1MbuAH/RYN
HswEQn5BSaHbJUs2bwjFyo7a1rycGY12hnd8sJ0bzgW+xjw6ijPxYloSwaaKmMK/
aM3uWHvX1yVw+bpACDelSayRLCaIlZB0+UGMfQq8dFVT+1ys1gi9PQ+ZAVxrXqji
SZurprD+Kks29cWwfHu0fTpRC7Lgq3f/apE1n/DmaHWCIxUeZ5aE5ydEXDqV7Gkr
IZGS3R2/pmr/k29v3l8pkLWCgEcf547cZBzC36+Z1T1ZBv9FZj0WR8h8RmOfYgrG
F3sx+OoHPoz8NqGh3HpwVnCNYMOuKwbCY/P16M9JUxXvdrVl+kmsW6ZdcX6rPckY
FWoA97sUxXFbXBmAGfuOUMm0j9tXKQgohF7dpVGOmhSlBpIMx+/FxTz/TNNmWo8F
OYDr9d2juyELMTf/tHUF/CoYE8P74BkmYW8XFNJJnBvllgte/xXovXrZlYZsddT3
gQwsTHxsbchYXdSCM5fQtQWFuC5h0COhufkCV1i9hoR63LbpvwVxBrpW3geVpshG
/CR49SqCbWV+bspNFnytPDjJgRH6YE9ZueworR5EBct7QTM2o/yrAYGFDC3HWW7C
NnqWdySMoZt2lHSzz+x8zkZASlniCdEyyQVrcfulfe8pSAIe1fku58aMsWCJJgcq
37nuXbxmtcWO+qh0jE3HWeVgcHWnLdSXffl3EC3vk+4oOrgm4UOkLTwqlkESaZ9X
pTueqPo9wDPgJcosgHYbATDDJ0TnjDBI9yZweTJCVuTHIpB98dhgCFSfWf1t2Rym
VQymCl+kd1aUkgM1Q5+k1CS2Dd4jE6PJQx8EGlML/6mczPE/clqchWpCqLdJiF2A
cLwlhPcJTgglD9aBQ+4ZHyeXxUCV6i5jrp9bzV7JghhvxPrPNw9qy7YwTf07H5Zt
0pOJNGI4bzK0bXL1JMAWsEQ7e+RlJfznudHHBwPhiUm0kZvvbNZsOFJoCaYBbTtC
Jt1srzV3VZW1Hfi6IMMF2Np7aBXnWfLczSTmZT7jV/HDFeoaD6gRDvFOLrn3fLBT
UhcxMYyDToywh9XltAtsbafM9xHiqdWhXmIsJUWMXVseZwspU+FgQXmG+rbEvZFB
FjFbmLNGS2xjjhSR1OmM6lboPRhRHCWw3I/uAEfX7a+M5h2RnVyDRxKEX7rtCEmA
yussMPenuxnWRdk2/Jr+94ZEcUZvpjR3VcSc2tJdk0l1Ts+M9dsefHgBpUMgRPTH
hJWwZaovCHwx7jqJUMczUZllXK9y8885+cG/DDhA2YOPKAHl22KFmXfAMphuUV+p
mmP5jb5SPPtygTiOEp9zmJ+ugMHGy724CpoadVW2qHjohQoLPsUuKkHJAMvLzK5q
+6VlsUzVXbIL16+G8LQ92mqOUCmaFEgU/j/H0TEA8BFYjPMByr79eOfcOdYcbUFC
FipXXQmVtjPKcZG0sOloc7TfDPWCT3q8wZ35u/sYz1r57/vJjrBcy5aYpqr+MQUn
i1xDSoYnAr6sVDHcK8nmDWxrFAU9hCWlRN/tEiRn4aYdyZYBFSaXGB8RRidgfHve
QGtsW9crr+GlEJB2v2NO15Amayd77ZnE0H13SuIkzqrS7AnE95b8xpOk0WQa3iO+
dc28CCbrgCeA7Tqt4mTmTeEHPG6AfoDl0hAPMXL+lTeYeUWGc6++qoAab9w4PyZp
8+i0UeOu9gbHGAk808mvKgiZ1rAYxeNTDFRgO4xgzfCo0PIb7DOp5pnhiTH0lPDc
/2E68SEXD6onk6cRc7ApvTn+2dxkgzNOyjaHjovnPfY9Hw+ZlOZZX/d36HTgCmQ3
AUNBkEoX+WNEpS4/x7C3WkLnqV0OcbjWMmQCHaS0ADfDgeqmOfYCTXrdgtKZQZOf
2n7z6KXOxYiSRr9nqMQCy76t7yPEzgicK72xuPf12Bjp1vwPCxIEINxNziNQlGY3
dTytnfIPB1m9BjY55PSVHYnxpiU+rdBxMlGfmC04pNEpgEK0gfh9arzYNDjwW2ZI
dH6dfoTuqA46DRnPGI994oi0FUj7SCDP2HmMy40QgPQpBC2ODddm9jkAUgjnYJM0
xOPOVZvenjqPBcDZDnOXO5f6ioeORL8fNe3hXeb04Ur5KYSAFSeQDJ0+8ppBT5bp
P030khgTBnACWHiZcPGzqxocO8epHRiRdV2tw2H75FIILrhYIAz/Zqre4bzIESWT
0BsO4quy1mU6WHQNY5hc0bCQL2CLDdV/B+EInWSbw+uJg37F22WFawJbClvqQvKF
1I5bUXDORSG1prZJEC31wqw2fmlkyrY1H53tzdaKMcU9xo/tcSXxccJvg7PUONmV
oESabygdXIFj2iziZVYqVpqri98chDVaRYXH3A6mJ2RvYEKvnQ8Ej0RPzUTGcq2t
uG5ZhUL1ifV4I1rYbxCYyqEO3ARqQMr8meNcyRruQsMA3+bKxD25nvvrZXDbAT8i
8MiFnw7bjxl4GznTZ8fNEoAPMRg5nzZPS7TPwiMct2SplirSoACOOLfmJAj1OfZ+
gojZ3V6oFgyQkNPyixZlNp70YkoyHboapsG59KSRTlwqF5zvO3w8pJcpXGKRLGeB
8gpOXy0ZTFyphxeH4tk+4mgPnAzU/Uhu7MpkLFueNnh3bCeKWqadlUJ8xuDLnNnc
MUq0lmp4DEbn3jYeS8pyjOuufYi1gXgV0VJRDFMkdHRIUmLTTCt8uJxG0kgfcjfv
uB50teNex5+7DWXS/Mi4R7mQ6cuWxrT5wbxpu4H1afwp/wJfJHfrgi2cYkTjyS5b
iyPcayzF9vrJFg+YeHyVESi14SeBnADH81PkiDLbRU+5O8mLeAjPhqhu/mrhyd69
ZPeWmjLmLrapfXxz+aX6mpmPqyKTwzsX0TKRZA34aiY3pIGdXHAmSJybTbFEgcwL
Ov/u8lGFV6vHA87ECW0l8YvnqPFtMFMk6TuuMVzF1JZCKHm5tWvqONIHbuE4iRMT
E2MCMgo1sqF8BsgOs7zz4PGyiqAfxH83wv4g2V/37zFnsnRQUjRoW7wXJhH/ac0j
CPscaRnYDE3eLmelzfZ3ANbM+RALI90Y/matX9qlluLgU60d8bHfgTpBfjlIrBLj
g4AGoui9oyu/oKU26G9E2RuryfDVFHWyMhaF4JjPBV0/ng4aIS7EtbaSZJ6nYb+t
BGiJIuSSNK0M9p6Q2rL2hYYmGu+LG+Yaxm2Os/y7rjqfvuP7RN6aG4xVtv72j1Ta
AaLyXxY0NIFSJ8sCfcdCpI+z20QsI1apTW45+dgKEvVsdX7DDpJVPsWp5lCsBscW
NClFLK+Miz4U3a8OIHA7nzkDbk5863aQsqwYryfT6YaFS656pW7thLu5Z7uID1wW
rQ+8rhZ/jlc5CW7yJ+9KTpTt2CRoPFF4481bqxTEmJyuF1tRLBsbA1eq8h6zIdkv
d8o1rJB/skIKVlZO49WB2b6kFXtHlGXAseUaXGJayuXEH1PHX4b7qNvYRalmPDBU
4rpqMak7uPplIzXIikJM2oIt3+8oLK/pgELnQ/ntzMwsjXWFVhqtBwEfPEWGc2sS
Sgy2nl/i/i1j7Uj9MI5F42Hy97twnxfu/ldH/Llb/21OrEpaIkThEw2pbkgYOc+6
OCTBhN3EMrcAA8VAVGlDYW5Co9f0nPSoupgykTyJmraBog+N3VuK0JiikxnNixt/
hFpnsR5MmGjD8jtoCPnigu9v+eJ/1NIopG6w9aZHmj3mgGUHjzfrg3YeJ1kw3Yp1
M8o0ldS6HkoaNvy3YaYvdjdHnX2w0w7zfoGJR+FqCpzi+vp+v7rWcIqcv8D5E4/3
y9R6Nrqmxmi2y7qzt+7N0LJHqMXMGB4F8BRSSNHR38GTeXfOaMb/FsqCbUPfYzRW
QO5ZhM7ufLS0mpa0GTi5TQYOrDq+ssKz0Meo3VF65jO6SxL4XeEjZ+kNCGZj9PyC
pC/lQZPU7glWg/pihy+kc9+Eh4E7aPvuabW2HZ6WeDpK7YSPC3lUHiemY1Ci95KB
TZza+90Zbdw82/b/oZsSWfDMS3J7PHVFeqgdgMASsG3y/kqWy+N15iFYyiuw8G3s
Qa4gJRtlWETQyHegQluoHGdeWADUiXLvQpKBG6P92p6y9w+aru9lQb4iabHasINr
qB6WdK+5p4GBGeFeRwvifvB/3DEPQLn9inL483TxDvOZ7sHNu0KlsQzoymWilW/y
YFtMbEr+ItW0p1Tt0fkmFb3CNa9YWVKeujhGym0y7nQnkABQL8VSHC39NaxF15d+
A7taD0mn3YEL2TYegCtH1Olabn7JNC3ASFDaj6Kh0mqyKodZOOphkCQqtrf9KhSW
5iD9WtQprns8a3wNy+/pHlVsm8qOCRO4AbPSLBRg+6+xZVA/a20IS0u83zzsIiRl
Dr7FuZWwMheRtAnYbOvAGPM1tvs86lKrdOitpKQhH5Yd32q1WOCXBHSRRzgWV0EN
hhzOLjb4zZwesA3nqcu1PptEUbhe9QLILpzz/ucGjeKJ838iG/vtSOCuc0768Tf5
wLhxW/dEBxiBxByjydedwv7gED4IkrQoq8c7Rd9ib8OL5/GG/Wwj7btmluxggPwL
s34JPVH3AfGeP990IT4yKy6k9dhldi5EDXx/lsGmZixyx/XG0585at9eW4tMmct6
EnXZJ+TL7h7K3Rm2UM52e2dO0ZoANMZS1OzWOgcq2cUYhgohjmFgtHYgEXUWwjOp
nxhJEzmME/P9lau+K+sdyOZnMZpGhXsId2xOiBqeHplObIDlv9jLWZG+KvGwgvfR
fmx5OSxOr8Sy/sYBfvKrNJQvSzBHNhoL76/CnoWZ0Cxxa8leKmrPLBx/sxIT1zWB
hoUe+lYnLGoB1fA+8+1AHm5XpG9UOxrez4QhIhR/WKkKZ41hDC2mUXv/NBag9Jdx
dNmHwROVbd4v0qxAX5WK93k6sMF9q/QCX/o7vgiaHgiKbw4v+ZjoTteziXYVdM2O
2i5s0CI10DqjoHh/utm1nWHfWBTVEONKfv/ksfT/oyHcS5x/5Q6E/GAy91Yt63hm
QcumFJbmwEBlSYEzyYDgFOTG6gueEJU2pbYpbBDbi7a6GC1l6q0RbwHlFzS+BFYA
Rk7m2V27UTdUFTu8ApEo0n1OxhbZMSJx4VF6nb5sP9d/gWA5VIoH7Gqo126+ZtZb
Xn+7TlsqB4VmRnRqHiSbBSRsenIInK9GR7gWVOdOoWk7kwJ5JmVDDQMhB0ZiG1Ov
WXWPr33f9rjvV58k0OXspQIdlP7cJgZlKESoRbJvNDqTsO9IOrFh7aD8RqfcEki2
eIp3CaAsBlDXKLLv2xD7i0uYOV+ngEX0Ku2gKjhx8r5i1wI9XvR+KyGyj4UKsTZX
t7bmaMUaBfUY0NG/PnqcBDP1fWw7bu9tz3lw3R02WEgftJillaCmJ77qwZHBNlSt
9baNYKFaam4zFA+6CPg4G6lmMfWPD96bQSAF52ECltW3i6OOV9YYWViE/ahk4Qzl
IQ7405uVzRMSoI4SlCWsvkMMG8MfNGTQPAxkmXs4uITccylahHEb2W1zGkmYsjtN
c60XYh/6YvpzqG3DR6y4B6bw9JO0GhuP/Wy8lKpi7klu2z5uRbU9PS19KfuxLh95
VwL2EN9veQi1nUz4ey7Epy1JGE5bF17LRAvwRZ9K5kEYlEWx1QLIDA+lPG1HgZDd
SHEwYFQVbZgatfg4/11ebE79mVHcB0d3J8Ntb0oeR3gc70jXDIEANVZM2LrECP9C
XJixAEcFYdZk6xtbz2HRMApou4Ub5RIxbD88VhAGA6hy9nehDHyackTgIG0swe+j
j5ZrseQbU9L76cjeuYx6IbJ7ZJugq/ou0VgfjUD6xGdO/qspQFQxaqh9dqaFnKiq
CZdzlIxtN2CtnsMSF27x9uCS0/D7vogIepnhBmwEnxIJqHl0TPzLOk89Nrcpqe8g
3lUvZyX+upG/xzEOcS1kOnf0wQDNTyE//pOwxtAsc4mavQl1MudVfYC6lmbzNBi+
3nwxEW6m3FuIZ3RcyxuZoLtVCcBIjxSWJal8dVShenrvnuGo9LPUlvyh6sHlu5jZ
PXg/7GZpjTfJeE3/tzlUswRVTPXxsNy3NHcVxU2gVmicqhH6tpM9svgI8N1os+/5
5+vs+3BHRuJglonBeRmAi4qROFpM5MnUGxHmfQSBkm7nOpVkS51tIpBlXurAYnGl
m4eNFhFmucvtpQs9nhwROQ3MEOVED88hf2TlxJsVoJseII9a5KRMKYW8f5mWrIwK
cEcKDUPe+eFIskTth8Up5XX8z/rSiBlOPSNHMK45yoShAymb6h0k4M8XC++vi70E
wvour1poPrB5XOaO0CSKH/dGFqQIYQONBmg6KyP/0f7FvzUEXZ67NzqWKhIPPfY4
IgMtq4/lCzAUPt7Je3h0fPsvGMaX1i5UURNkMG9BMn5PXXBYMBWQzKDUWwdoKD8e
50/NGoZW2G1BV4MaTdob9QCvYO9fieU41PdOKQry+TEe1QUnNBeu11g0829rpqgT
/NwfExh7gjMX29b8v+0rm7vx/K5iKpl30o+xH/n/ohvhybiI6Q55+nQlBwL0grBF
JBzLidAcbNsFdZII++C/bpWG02jqyKT7CdZMF03IyFWwQ8YjOgZ0cVFXmBLHYOwd
6IGRI7jlEMS8tsS+3fbBRwuL+uCK4aMBdfdhgvmLZJFQShlD6e/SiAoO7EL5heJe
nTp6CEFcijO1y3ks1Bv0YWkCI/s8n35qGWfVV+ramagrMkxPgiNPJAZTGRspphiR
BKEZ/7IEYNGQKjryULCcndAKR6N4kO0ei48pxI6agyNml3S3Wpr2XaJbT3ekWsu6
xDNVwyQOgrqPOCxvfnVNKQ4wCR43AK2hTfvUQS05SS/a7CKuvVxkE9V9Xx4CXGik
DaN0TrG4YqfU56oIqdRsxoQ3afsiL+dBnpQR+mtOGh2BLVxuky457Ugkq52s/7E8
bRHS7Z7pkD9TfBlq7i0pfwPFyOzhkkkdYdl9nNU83N7DhMXVng2jRyJO1dT0dOW9
D1dHvSfLDybnggjk3302Q+KpEFImGrSxGiSxUxy2Gl8UbBmQZ+CaTGKBkDZXywup
Uaer+xfplNd/C63zg8e18nnwGo++YUQW6vBiCQihTHnf2WDFJtD9JUHsf73qcZFD
yC67nbuOOfMn6KsJIx9zV7nDAPyOswJnA5IXwQOG8P4wFbL5yMefdzMqx5qHC/oE
kSqhtSNAsB0CR4T4MjK0GOWFhDZNID67W7b91WLXQXkr6KdreOrHEseCG9JkOFvL
Vi3sVCnY7vFvO3oOMTBST3TdxMSisVjHpjWFZNWLSsPyIw3lDqM7jvrtNftNByrF
5g0S6xYGMLwPpe7uPy0eU9CAEJ9TSQxNbgO+uXx34noJ8dGZ0ZDqkwVgEG5kJy0j
AcbFqznM2MVkeZHwlc/J8/IdALd8DSpfaCbKaOsuGbylwLlv5Sl22wCW8N0xex0v
lWcPYOvwzjydVV0z1hh1BvfsbKzV0FdFhXGMsCXr/GZAi0X2E88+PPddO+njn8l8
uQV9rmca8V9ZQCOmIw/xeuQZpi5yKj1hbiGD3Kgs/Y9YNGb/nKdQv6QGnWpCJMY2
z9HAT5qR0EgOCKZGUmcGVq8B+gyDc26s6EsEP8eZxz9zpG8v+vD+D/BMKV/PWw6J
sqQL3HB+P2m1cE8n3nGXd2GyhfZCfr22rU+z5BOST0VqLXV5QuSm3MZgKv725gId
zMCMuccv3QvYdcjm3aWCRtELZyIKnqE9zP4iEKFjYpS4rHqJKSl+kJOc+U4ghFys
Rda1uAKtBI5h9JQx9aecJ7ljzoMZmDoyOcE43NdcaGYr8juV1VGSMCWUDw+t55Cn
r+Whdm7asUGomWvYZ15S0qfCWZs5DPEFUulBhe+6ClSuzBV56aUyMNM1MwRKyHIq
Aq4quI3IuSHooFHuY6JYktVL+37Tw4WrDvzIGYXNQI3Fsw3Y2PfB3Qjl0EwLYsiy
50pwuDcBjni9L3ZDuz+WAiwp6lu63L8odrpV7kOo73nVuZK7B+zod6LuLvuN1cN9
qYtkPmDd5jJeZ4NrmVV8powi86+S8di/Ablzm6D6OfQ86a2B9Qld657Ew3Y+Uu8C
16Pqi1lQVaPQ98R4VxzAqsH6j/wuGZ+tK3xDkstG+bTPYYzkIv1Mp7eq2SYz7ScL
11HSVtUD0kqly7SpYMwm92BBi9c2IYeTaV/9QUJVVc0gCVlr4GY5J5au8v+ooHyO
D/RmK/+1pBD2jg1u3hrcB6eZWzMkse7Mr0JCDYSs4SX8vHFSV1iypxIS4bpMcBFg
Pw0zmoV/lJnw8+gLuWO0ebuNsxitL4S21VFet0CHDgcid1NM1IhqJsbkEXulTkSI
0ZwKF4sOEYNQhnQx50Pp44NO7Q/6X9C/O+Sq4idj07W04Yi/jyXcF4URf1A8jw2z
KcW5+gLfzPMxje53xdNXLyOpicR5GJEM3dz4jYe0YNlBmQOWGGfB84VOiw6sZ5AD
3qACcnXVJ4FqkXKQeGJQ4pBE1NBe4HaICAeHj897WsA8KcNkKWK/U1qeWf8BQrwi
4/j7nKkI/XCNZiOUoqv3Jz4DaMDZLI59oEYs5sIRljLawCHKoFLaKTI0Cc0tzUjE
gC2G566dpMv7PK8SZrAPoBVEa43NvSVjRxw3AKySY/6cdXSM3vFYzmD8h0/Efbm0
SInf/ChNGuDjK6MHHMErn+GkO9zkxPJeoF5bfza5SKJa3b9ja4C2owZbSa+w1tDn
PAJ/KTqNzGKQbYfkzBeH3b8F2iF5eTd/14eV4FtZENTPeF55fxQV48IDOShqMRGY
/l2ngPqcn9Nvz7wyliz8j0Y3mQ4K4wWIgiOSmqBvNFbz2yIblywyOpZ4pkvOYJnA
j/155n/q+/QAU/yUWk12omeEx3Lf/egtJWroNndZh/cTuFiMM10O8PuIL4C34uMr
6f2sI7aCy1s+K/Fnve3HCqIDxsYH8HNvT5AtoN/Fbr8Y6EFkYfH2ykYqpGUX+RaG
ss2ovKQYf4vd9otkA5FRShZXekBiXzGlqTUvMS6TyZuQnfvn5XYJrWiBeoNEABH4
f0cd+lp2JB39ElSLYcBGtEm2R23v75hNByyqbQoNUwrDHi7gNik7RfG+clb4mYoX
aikpcswBM/NSCay7e7P2eQZffpi3OqYdpnDHrwiF6TJIndScCT8W280KvDMs5o+1
JYlf9DL8wM2aUmL5QjBAsCMVc72y3V+Squ8J1IBACfzfKJm8KqYxGSpbbuwTdK6x
/rC9LfXSClEGagrnvNidlBP+e5rPa/ptYg+vfWZKwLU74PlUyBcpjFc2raO8GFwM
DlvkapLJmvQTW7sdLhhXnMBCC26QLbAaSc8qmo1wrs8CIK1ICQ55FbxcCTTIBBa1
UvN+f1TgR/HbiGEKMBzzLDKw+I+5nMiLYIojselLVoXYlwKmMow3WGttdIIbp4Yq
gBimVU6Y6vr8z/aJJKh7UCT/cX2RPBESghreuU69/yUoJYpn8bKntB9BMRtLcq6y
mvm0RFV96yX+O3T+FTRi+OYFVAi80lMCU5wuNyvHtNK+Ke8viGpRPSsR8CcqkVGx
gD/6EL96QL7P1Mq057uQ5Bm+Kosa5vzg8l61IfXLeveDpRcJp00/obJ9Y7MGI7uG
cs2+taLDejC7BztbH0AHYxEI9v6jibS6Zlj7y12IlmuEVABCXapHWvttDINNJjkr
KLy6XOE6j/Ao6IgSdqeOlLN3nce3zJRiKMflYT3fQd+ZrYUG3nHig0RaLJ4o9ecK
bZ5ozKLGWM5zLRo3TEYzmE7BCz7X35ga2tY8LIM3AHk/Z0ylbxWQHUSyjkCNqx2c
6L/s+vOh99M5mFpZQm1v+h5NzdfP9LyUNYO4YFrN/kWu9PK11X7x2lMe+t6YOefa
lwxQ06uUw0MXXMYSnmTDGStzEHSJ3AOMZNuYDcHgzZZRufsrAzkjq8f6xChlRfjn
ZUu9yMRy+FlXI+/TntccQrn1+r6YOajnka6M5ORznb7xsUF8QqQdLn6v/F9TNPi/
98ND1v60QSS0m/4eXjzlF/KVJg5kAXzQRzr6fm6Niw9Iyslg2jR03Fujiy9znezP
Bq78HseSgQkabdlUMgzZpKEU039s7pMGshG2ic1J8bwrOt8Xhd5uA+D7VaZJpgg9
LsoRUhe5JYqxd3LOZhW4Ej7JGJyPLo+Kadj3L18vEwdqxLThx5SjB+AiSevFOECJ
dm3dLVDRiG6b9LKYRAA/hfcFY4P0YbIRXNtxFsz9ZZLhLTRo/RkUpSF4ItFn/zNQ
r1/2kEEXfvn5LjlZeG+Lyuk2LMlnLMlZs81pSN3WVLla2cyV1vTOe1T9EiJUjnkH
NP1AYHBOEESyMGt8B1wtO/ldp6+l5sfUy6gJU/OwCZ3prUZ0CnQFUu6dR5+0Kw76
61JlzHzWtlSDu4HLMxIVRZfXTXRHJJMP2egQSq0MdcRPpRHCYu2G8X+enaBpqgL6
kWe8ZTYkcUMy5mf3rEfWQeY8L46JyDOczEGlzx6YxSAMZJDnrNT2XRBivLowf5Yf
oedtCdHcAvQBX44dJfwy2zNSiQxH3oYc9BthJC4gGy9EWRxXq4G6Pp+BSp6wfwf6
6w0degtoiS9uCbMXnLCRAdKPyP9cRTFPlZhj62/RJBRXDHwVlSCYdwgIMc8RKGZS
rY3j/2e+d5VlXOSEZnpHqyqlNApV6uPP/EmL77cMr51BoDDDUIcO5Mp+7NeGk78N
C3a7KMhDnAHuTTWdYgRMTWQ2AynTkvijckWTtw/wnot4oq63B7iJtrKz/eo1Coo4
qFLr4+p2Z/cc90KwHYyTaWQu0YcDDrsgCv6VMubcO1RgNiR0Wna7vL97X72xvV4+
M9xbqEr1C5IIrMLa+667f2lqsXoQbzyBS5vDhtEEqLjQs7apuogk6UUH8GqrAXMb
CU0dgykERDTIJg+iLrrzgSJ5XDNwy77tzcwGIztuAPl8lbwMmMLO8r9Iv+hPHzCx
1KRHdKIVK2m6RHTXzRSTpGF4T069YeqzmzjRD9bynKpNchLdKrKLM4wTUKvo+24g
j3wDYCjTA2+WxYBVArG2UQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cFmj5GcGam88r09u76JJNzSo5ghiT8LaVnGuOSSkHbIPBNxtcgtjaKh+/nCunDv0
9RHfpGYU1YAnPPxr4Aw9z4Re55vTX3unGAhPY02ZLlo9i5XYuUyOGw+0U6yyMxYK
Fpl+dS0M1lBbpJjI4vRzrz1d9QkwpPyMJY8WWavBKhWw8B674z+/JqCblA+JAnrn
HW7JaWKJ2BjwuNyTHewByMDkNyEaI6zly5XqeEKK6dkt/eycp0q/Mkb/fe1xNZYm
fi3N4WuLUWhfaXw6ZU+XxrjO/58+HoSK+tk/YfQ6dsQpXS80AUPpZIpVXtf6yF7r
KxG4GqXXjTtpKzJg6vZulA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2864 )
`pragma protect data_block
ES6tOWgm6/wSC91xu7OuLJLeS/IfiiSw9ROyfdVUvA5JgDFXkYRiKrddssl6d/KK
xqwJjDPzL9G666M3h9LZQw1O6IpAVWFUHYISW3bLAP3I9jaG6KcHnRB1P8F7TsR9
rrAXmrnZcy5PtqJ51gG4/MLxzKYG2bzM5/pTHg5Kub4VMyLmT9GCZw/rjpsuzn/2
ZCawKEUU6PU+KIfVHVTljydVvtrjyR7aakuAo54YtLTo49oleWkRpAGgpeKQdn/u
NnJXB2OxGVV2EltqSF/wF/BDDpql0SpGUMPtLHk/gVZwid3comK/lb3ndVaCl7ER
6pZQAyiLoWo7jxFWPNMvoK2DDtA9PkFEdqKoe/VIPv/4dWVCWHoNBaNvYPtPN251
jmmOdwl1QBBUkw9w1CMWfkL6mMxqFMT4eIDYDA2mfjGGefuS48B1EWxuHBipQSfe
JTRsqjid2K3zzXZGae4i8xCQmqorWa97hB+ui3zs3QUNASNV3zuNoyIMbZswnm+8
R1h1lxXfq5b3uYLnfdK1DO4N1Sy5Ak7vuIUNL1yvPeCtp7UoYLkkIt2W3AtGhyQW
e43Qp0le/HFfDx4jwYVo7xIZG5MVnddDKN68U0Sg6zNEXRy2LaR0SjvaTdM5q6bF
M1QY82aSj9YCVsKsECsY4QxNEZpMYoJ63JnVXV+Z+3vlv5lhQSAGe911kHk98jRp
HufCOtwzy6gzjoF1VvBNdG8h4tFVXYp36K/0hC9GtGYiaJRaSXO1LUlR2tnFi9fC
gBgFpHPv/ZVufyGIlxWnUyqDdMckLoJUfn1uUmcKmwDH4JZ3b8NfdTqLL2wR6LWf
CwQjsFRAj6/+jo+3ZIn+2dybPEF91MoJx85FNnILeYjUu1PlZ7gQxo+BPq+FCaue
GoQrFg37J/SAli8kFIVKZHepyIVmJ3fkWx3j3nF7gvuYgCxUL8E1kBoQx8TTWY7/
DXpL4VybH/2tqPdXcXd99pwJJKNkZPNIjs7vLKpJjPibcj8JuIcqNDmxIu/9mxoe
LXtaXasUQcw3HA/Dd6OMGa8uTv+H+zNuFPRFUiy8hrCZSy27dS2Errw5FPnWw8Cv
FjvDVAHdxjpCxzCG1G1q3K++D3UsQn07wpjNwkDTPrbkaPohSl7ZH+5B+DRs/FeH
lZnx8TNY9iSnUjQ8yX4FmZvnq18f4SrOJzbUg7e5F9vPAtqMwpaKHnUmwIUAxUX9
l4zjWJj5EjKf61yyOyfrGcRdu0pzN1FRW3YRgtzrENzmcTUZVp5vhqX4mUsUHF1c
cZCdJylg9HLcS530OwIXsOQIIbw+OuiM64NZvTxDYlWt0BloMxOB4Mn7KxN2GR8A
HTnQMz4OheiQNFo+u2Rs65oYSGWQGZ/YDomGNH3ithaAiB13yI0ScjAb2eazJESm
oh3HWctGP9WmCDbU/+dOBr9/Cww/0mc/BzEhwV3EWSNXOD4pIsX0Pq64yk4izlnl
bjwEqQ5wQkfiQV4VNRctj/y9gQCKdFAG73O3Q6iqLuaPTo55uSU5+MzJQNFVxENm
+or5vN/qdHb4TQckCmNViiuqneLM39GHn2TYMQKPfWK9v7NPKLK+Y7j/DGZWQ4oY
ZYe6MzvV5q2ZtLWitm+46WgJmxjqHXf6CxxneSyNzlXJJA0+u6QDmmvoM1sfYEYt
ZH+WYmXkPC4IuI6jr6Kfq2Pktya40srPqysDaBSnO36kF8ODnt+JSAMRRb15FpIA
tWAIGX/o/T9lNBIQU3gEmZXCCGuCEvXRfKm4HhGQ0jf0gem/HVJgBbaXUCRh5Z2L
JLNlybx9kNPIu2aiCIG9SxG93AlfobOc+ZXmOb8BxaSGqccFbFwq7rMPVX/ZSigr
9oByD/wsIN6lyeY2157TUoToO7/r+j5nn1xoEMBoPwNXfh2nXMW6Yt5Dcb+kVsG7
dSb+5Njo80CFCc7tMJCaiCv9c4I0rNEGM2zaMt4O89ACdb12KafauwUa0qyMFEkS
25QXKbp8IvpNlcJp1y/Lx78sjfq2gKjjms/ADf+KlMBMwmjQRglfJrOR2S1tuS+k
4Z0UbAGK13Q46crA0odaGQj2cApzAU3R3VinEq0jqdANlDyyZmqSjzynWvZOYCo+
axDTFKysjkXTP4dqiYKudVwZUSirnQhKtF/sjnDwliDrHKHVPArIF08Bu1ydA5v2
hPapJSGdF29QxsNEKinOcBFrM0dB28kW7YXpEFd/or3oDdP4Y56B3qusTKZ0ioyQ
6IqD7+qa45nLpG3E8Yvix+G073JeNxmAvOVS6q1nwtYrPee+esq82wWBGKN7nIhU
ZAbH29YQO4xVG98WL0XlHpwoJg1uhd3YZKSdX7nfpVSUNvdM4mWs+QjCTBTLc/YM
726Bw4xJk1WccZm2GNaYdmyPXKhbDZReFkochyZHuN+6VjOCkWFS1c1tFTCgUq6S
X++EL6wKtqtQcbV72faIoEMJhF203NgSaTUYBsmpI86bEBZvypWF3YskjsNwEW9c
9i++vrIVakuUpSvwJm3hbSgZGESOWoz470Zvhx2xakhlJlWuZbv1aDrH8akl/6s4
ALi0lgCnfdO4jpu1LuJR8KOEZ4KI8loA/hfyBzAuFtyAor3N0s7UzhcbhJtR4rrt
2w7uMten3nvZptzVFtkuAKOs/kGCAfpc8ki4t2yrnN14kE6IDT0bx9pkiXMVGvSL
PFLI99XMLXk/3LY1a4avEdLOSdM6lPc0czawczqSqmAUOcuXgURCDk54t+EtNFqJ
O3AZotYMQd7DiyL3o2CbrLHATJi60PZeUGrZngkv9W9cmbJVKIszoiDeL8iEDA9D
FgrU0pm/ld16hbib/uQwXw+Ye0eG0bGN08T2fvIFBM1eL75HKe84Soid+07Ho5XU
OAonfgiZpdzf1eDc94p7MAHQCfj2qxGTh6yrEHqtN5YpfJC9ZrV5hzrQHYIcPVZ6
XTXNvWujpwwuH0Boq2EY9FzPccPeV8cSMhva7WO2XU/UU+M54CrSV7iDNGD99T95
0CgyqN+7kphOCTUF+nQaaiz6s9Oab2Tk4TrvxdOxcatVOGKeYXXAzW5uBop+Ql1O
RBjRmkooLv5IkG2zEdDkfLdtavkzFyUvRT646+iEOEbzXecJbsxkdn6dv6DByY66
Jp5MLTweftxHpuzmAh6UZ1wiYEF/1lqxGhefmCITnBkmqwu8qPU52BU1BWycMPq/
5Cpa7X/rb+Wco5k9bYNvInogFvnClKZZ4Kx1o3iV1VFEY+NTkZ9geKwkjpVjWcgS
0yisjtzBKRq3wyqJksEQbcpBlc019M8Bl3ag+5KdjlBmd9rXLlHX1bMXJ8XStR/R
nD8WbazTha+OjelN9ATtqIDF7rtVyqXFMCjoNn94o77JXzvFlsdMWY1ZUqgqbWyv
bOgO9K1vxWOX4mklaYYUpyWfHow/kSzNpN7BYoonUVS46w4FzO2ZMYEZDVx+ZOQQ
46jW8rUTnzoRrOGhg/htpvS3CLDpvJPiS8biq/Hy3/ygIF9G5MV1cNAxW28GN3NH
QIodPHXUEqznJsd1wBmXOWT790dZ8LGaQzc2Dt1C2AKaJmBGAvqkH3ZxhbQICGwe
mXbES7lymmhva1cUVS9rKM698ub67mw4uskGj+JbcpQe4ccRHXqCvTLuLU17Zv3G
qI6Yet8Al8/42xfrqZzZ+by5nTCs1ndp5h2ZFfS4c/4FT8welmrcj3IGcCht32FK
oalkmK6zMAJTIt8UO9vRMDqr6pQ1SYzO9PXD4tmE2BruNWlYwvXL0Bw2XId9CEuc
iyXUM/eQomV+3jVnHomfBckdTICFBqM/KnM3wbCiPEU=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
H/qNCw80s94a7WBIPhiFe5lgDSEqnyIXuSvX39w5jyy0R0mpIweN4jqkvatrMuQX
wF2MFCGiN9KJ/0J4zllmiPeHjsW9QTmYTuttc3KRPgJbo7dStDVIqOB4iz1Bhqup
icmnU+AudkMVRHchY/KSvMM+53Ti8uoZUUXrr+5Jzx8ZqkY7aWahF1lZB32QTVoY
0wDdhlYOO701kzMl0HH/OSEs2A1VmX7Sy1PioHVf7s4K9SD45bqNsG/bdT+hbMkE
93QgI16VPq9p93g7z3S7i3m9802JOpgMs9AEIAK1MPRgxSXzPGHG8yV/TueP0Fbh
LvGRanRRZBzLBGLzP/y9Nw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8720 )
`pragma protect data_block
NdJqYay/u/xOtyJaSyFfdfdmNza7RxOv6VKePahae/wVOPe6QTfelR1u3yaLzJT1
jz4f2ZiIV1PYA1VjSeoVrMEzRxYeqSabDeMyU4HtP3m4NXovDIzxLcxZ/CvmQ6If
7ezgVr8GOghPQJvJ76kfCHEkIQlSSfg608Kvc/lWBPjB0ih/1yaB98Km0Xs8WZNd
QC+ujUzFbTz6R86yWJVuKDK7MUKqBAOuWF3CgD3nCT57ccImEKylh+bGZF2ATdv2
8rangKFEfHaITJdskSKkqZ5C2pGRHM4ulSllBg6+3qiQ6Yccovv+dX7Kc/k64W5Y
b08UHc+vtDI+QlyjfHDj8E4iM2qtBuV+cdor8FEo6QLiwis+ZAprzsEoBchL84cG
ZIWSI1ff31Agm47fItgnX+t/BiMkZd5CH5JgvQSwPSqLmU3/NxySGEeYvuFhoCUa
+nqvk2tG/O2sRPDFBqcWe/FYpBpCKXW1cvKDtKmGtsYYTMyEN2dEedFActWCDWKX
zl6IK05R2xLpidaoVpYXEbSOok19w9tArFH+eOo4huLZObrc2uos6meNWJrkOjs2
bl4gghGKEtYPkwyyfhw3JLh1E1IGIkcRpjJp6vZcsSD7RINAfNhMcUP8x1Ooejm2
mYAS00sm+wOrvSs41N6GV2Ri/W/erSd2m6svOqOW7rvIMWr+TO6Ldv2ragzOPauG
wImB5cXAuh4SIsai8MFJLWK8WzVMFJjK8xMsA2ri1pJxeoPtomdr6FJF09wToy1f
SxIfjw2N6eGBLqaSfEvzGYgiH3JOacKyPE0YdYHn40jHEC1je3cWH4mlqyOkN74l
d8bnqcQbN+RyegndYe9JnkQQgfvXN7fYExSCZLvnviAto0wTnk+GhAvyXPitSuFW
0gMm12SQYRtl9F8bhiWHBp2X5bU6nLuySyGoyM7X8n6fw8QsfR8s7JK4H3vM790W
/sgcl+Uyaf8rVVIPYpEznXAvxFrRYrk1Ta27MtLcwgkzgOuO/HQxW/JuzqCgdCIk
5sU9xd6sCE5N+8dD7uT/gWFeGlbeRUDT0uANBTO1T4YGS0Ysb9PvXEcd+xzbSMCV
1G+XMO0kw5cc+/o6TwxrLQdLl+7n2ZmRvb8YCcbifKbmrdpu+VauunuFO7pRCw1h
Z7sV0S7bA/4/AGLKmyjf231KX60GLE/ye16WRxb8mVOszkw4TZt2IjX+7ElGsfWT
lL4zO+Th+EdMY46gaKIgUMiJI40fpcGvLj6QZ0Rbo7cvCQ5DCHuPTVkYDaPMnf7K
bCj6veYUClkJb/I1MLeMmAHhQ/aH33wp825hGm5Du1hWmuY0gb9NgCGR6teBeeTn
KFiYF0JG9MaLGnqQDMBE2Vi9rB8CvuLX598nzk1Qy+BUoXNjkiOaH+cA4LjBB9Ay
F8AxGS2qaQrtHqhe1530dxDVvJhqXln7vh6f+LBBgVK4OZHmpzxbouG7z43gmGjo
NVQ79EjM2Ryr+VZtkx+HEAANvdf9Vg3zlR/oHcl9nBYSOr+OiGojLiwnycO4p/IB
zw+Y8IelB5czu/ZOeHsA3+8n4zZ2+3Xccw63P4jCZJ4fPNdv1Y0ZAQmvLCgNCII1
LwMpB6ZGsVMPeVH1Gf9gyqPjaNyy0lrMgZV43bdAmXEOCmJpyFTI8abCGg1odLQX
yRPuwM8CTz4vvRwrjrTEngqWlXVvoeUGeAnC9LnHPBe3mqJPuMrleGEcN2y60E/R
Ttdq4bNvtpUyZlV2xprxAFu+xTV66YTZBNwgGcleUPKAQ1+09dV5DS1b9K0Hg5uU
Csc3FhBKtoekHPDBnVsAiPy8Xk0CnLjIIAlN8nNqLCngIIgGkQ/ddhbytU5KGCF1
MosGqdXzeI0crveUNZfTdABBuOGA3JT9TqSfRgbcY1fR9gXRB62f/1ZBo5lUjfFf
XICpfqeL0CcVLPj2nEc1eqgId8iGYPCkjrptIGTTeRNIt7kWLF4sYzHtxnf5H6ur
/00Khl+fmrQEhiotS6Hvlf5UAYfQORmGjPk0t86Ey6uw8yeKc4DwOyJlpKlrdIrH
fkZAaysn6Yui9Vifh0tKlkOqfzRIz/Mj2iYi58RBbJzWFTJkeD/QLf8dG4ukF0Tx
LUgJqgo/JXUiJsRj54rjQdx9D9LIna198LNpzDKZfiBhRsPeB/kQbI4uigzCYpyC
bT9J/njCi9wvnhcGXAhNxTDaS17jH3g1uAdbOYgA830x26D9p3Vk/2PHY+/y+rfj
oRfYUGgLsCYkFIR6Rz8B49bXaBbWqMeEdNdSWSRLT3c11iQO7N7u3HUIHi5iVMtp
oUup9Gz4A2fI0n6NzsUuxCd/BNOIGEkqaGJupxWwiXKcD+ggg0b1cbuHa006XTvN
TggLysin76wtThfacflpSOBf9qwQYgYJXPsUTlsbyg79a43XUtjphqfwMeXlLejM
7+qDxLUEyBLFign2UcfdW/y62Dt8ENh2euuB2EEQMC0l2GYbRBoR703Tbi6+eJcO
1gdWG89uL67r6ktj9Q+X6nogTmiTf4D7izhV1sL3Z2N3iimx6IQ1QDIoQke9GBCg
VlNnWmQXAKljjjiFiXgLhc5gz7kUot1bzNRs+b1vfBYk8VV6AR+yvDC+IV/DKCvW
fLf7tQw9is/UkPI62THaSMksQp+zzInpmlctJhgTcc8yu4nOWEp8i48zhmSj9aj7
7+SwWiHQPqB8ISkKjRAH2Jl+8DULF5LbIWApJbkwV4qAGIc5JWzJ9kfNJQ1TY8XC
HPE6Mh0hxLbQS0s90iOU+iUzPFmHcuLfN0AIRU+bmnE0t3CkwdBfx2YSIOFM3wbk
G0er68fqGK9ghiTm+XQ/KOxDnB8d8ERcpHdyztuer1qWyzJQY2AveGgc1J063nea
YneCwDKHHe5PGEXr/XLSXRir/JWlHTuK0tKQHqkckG6lAD8zny1T502Uod6Pg+Zs
goebu0CqEjFuTPWaHV6BMBTVx3MNd4wQM5ZQlkCHkJC5vAAjleyIe3MKjW7LYvLJ
FiYJJ2Xx4IsRwVZk3xcZP0MMvkylshn6V7LD6hwdHsIXoEEgEsjfrYk8O7s9air1
cD1ro9+oCwRFEOPgxcQQi+ESaURe9JNDcF4rqZH4ALsynLERpWtslonIg5ZpGqC4
wcWRv7Q0dK41/F3KV9MAMUoF0mXAKLM1qfZDRA5mPZ4YABrzjxTW5eOB7bf2Yye0
8o61c8Bb3ZCKfGD2Ehqk0CKxhz6gOo4+n240fCDnbmkCTu6VHovzO2igHa4Z02O/
HqJMl85aaFjwrC5+cEFg6dV9e2kUGNhbKCVSimVjGXYvn8A4J1tz3CA3u5YHZ1nP
Ggfyswb2aFTXhHLY5+HYla0zXufZb/NxX7zEElQ8PLaxVw5LUdPPKjuWVwcV5y3w
EcMFuOXZvyumuWD7CIoJ7i/q0wgqgvBK1puHY4IkivqKNCjF/iYfQ0GFvKJ9GfaQ
zq9r3kTDOjqZNqZcZKloRzPZddGsFAuctUCdzLJrj73SnOj+chBJUcNSXun+IiLE
9cRBTgqpb/dUez1Bnk809ra6lntpZ0gsolV547WSneEgPQz1mHV56mtNAqf5wvY0
keq9gKvAOvGVP1wZWDj2T13Eur5WD2ryhGZ9NiArKgxTvhlN9ilcGR6QH48UhPy1
Znr0bTl0Ql+TG0m9fJI6R+FItRmcNPR7/GXaZ+LBdmUWyZ43IM3fGh9bCdMuwg57
Mlfu7oaEzczUxa/POvgzgpexHzrUTHiJzJ0nA3VQMmKcMhY9IJlOP6oDhIX4y9Nb
Hl3N3CyKLXMeCoBuslyN1sYhuFkF5VoMrFIALJ1ZUKD2CyuKJrnpWtEBrKHKy5X8
zMv4m2nND1QCsJIbVg8pBk8jqyDGkaX25SRcYFsrT4TyFk4YPx71VQFkKRF8Aktd
pUO2YH53N6TK9JUWt+GnX67wG41QnHaVUdLcGPrAsI3HngctQkhYJBjIRdv14dJb
7W2KcwVLSjBwFaW+ROA9ZizOXMM1LYTipAQnrA0fg6hw04K1wK4F+0RaJElfCRmS
BM7wGh6ivatT9RResilpnhM2oV0xl030C/R5jPzDQqTgazv57q9mVRuzp6v+ZZx9
widur/dHjvxAyPD28xrrVUj5YHPtsnMqTPNxqRLqMIEGnk4ALgH3eSzDtV9N93dk
vscKNNBkHI5mJaKntxsTgOaM9tLUfcsRUkuqZyM60S+kKDdWwJD915+BXqSKmPSW
m6FVOzyMWl6ZTrixiKfpjiXLZBCRUGFiNkTAjhignC+HV3KJi+/H6ts+c4zlD4BR
+pEjMp6XlBXQcXLBsbsOJ6h0kWBuXbPfK9FRW1QPMWvDl26MrkmncRUcIXExoWKv
O3aUMo2qgBowCicATNdhXhuWPxzYb+RA09/EtA6mZSrXeZmsWUrn7sQHT6Zm7v7l
yGrjoAMe9Y8cgoKQ26Y6G99bQVBJrWfOAx2nqkDOvnC8qeIgezGLp78j9GKuHDUa
wGQTJj9Yv1w+jA+8jnn5m7kfced3PBwr4yPAe5t1gNpuvSxTw37bjXc4eABrxZ7q
zerrh6fnF0C6azULa2cFq0g+4ztNpRMkwBnfWdUpfEFhGGUQClzcq/S/avFvoSC2
28N3ssNnobUQL8CfOCT7XdlxtO53hc0GsX16JpMANzskMdlsTS7aqW4F86zakAxB
mbdT8pWmLcFV3YiXtDGovdRKonrEn2HNUVPLIubxWghj0HxOcdiKNmIJMgnJK754
APieLyOX2HdP+AgIpwcKmvG14yFWGIX5Nu0PWEw7LJmUFytwLElZ7XUrZwcb8qoA
dunF2d6V9z06sHzkganUYXqpXxwnMhzZ4ZKmSsOUtHmwGQnJE+IjYSw9ivOGo9K1
RQiyNBvzoFo500h8KaZGLwI3T3zug/8kzftKrENewwgvb06fJs4DxQ28Q0fb1MiM
x8Pck6yddS00V23FsMtWdkP7x+BZylYJBOWaOrEP6mukp0RA8m/GdRF1DlTybQ6n
QwFnyiec0yVMaU3QVyXI67Ar/gWSKXmGMIW61tx0IO2S+DSl/uIa8GH1YpB21ORp
UOgvofBUuujYVoPPyZwnYlr76RkJK270URhc8YS1m55+yz2iCDsCN9dskx82fXh0
N7g4Hd8H35T/kmSKupzWsqzNszIsF3tICLEVweqSNLrSgKTPXr3xHcWngb73IRy4
qqFAFWX5npBg1z9tmzzycJzOEsXqIPjl348ImTEZkgEQv1ZWH/h8wPg4T452eOTQ
MFmFlJ5os01t6HaTzxIreZ8nVxWP4bCllnoMX41nysc0qg99TUK4qb9rHiVnnu5S
opN+45Y6L6Q0Nl23o4yJryfPsSSgZh802WM54V2TxTt0dmgjymKSCuTM89cymQrW
t6UHQilvXjieGol3irOrFvVMls4jatH/6DvJrjZkUUE0Eqp7bjHXEl191Cq4cqlO
G4hexYySS7XeJrDA7XCZehJW/sNzS1WZvMNi89zbFjE7ucMp/gb41t+30c5YubSX
wIHV4BTlEAaQPRpafJQayHQ6teDLEEiR3H9MFwmAYctcssvAIeRqzNczkwWqNsX5
cDFztpJNWV9sC6Q9ovmXwfZqGErCBu9A9/m46pAL006T+LzR5Ga9v3rFpfqfvKJO
S3rnvCioxxPRv7M0aycjr6M2YVJ/bTcwRWy4EQdONv8YJHllkX1LgTAkAU5ITG4t
frzl+I71GjNVz5Gzkn02dDHYbY4x/04Z7Mwtd5pDRogIYvRZtmo0NBw6QIJA+X6S
9xhFS8ptb/ajXrrD8ihFTsPvkDOOB79u5jOVKu5osQ5RO2bced7LVvHn19twTHM8
T8A5PFZf4H1kZ8bxRJd4ingDaZfGUXiRDq8hBHhf0GVLvfTQLVGt1yiqIQGhUfC8
QvEzvN9JF5bn5O8VA/pUffsnVfmkNsa3mVqcY+Rk3i1AgWfFSGUO/wTtTwLsI1TV
6P5im3ciFeE/vNh0z6IPIRoRBtktQpKOmzPSu7vH/dlcBr4ZB8ptJmpNN6YXbva+
HbMJxp/om+rgFMprbZf0lkmAxfCsuhi85O82rUkagQ8lF76wUIigL+QqdIAPMVh+
iwKaC9QCcFKDt2u5YzpfrheAf1qBTZ4tNzqc78NazdWMTNgic836fsE7HWveMr9O
0RlZ7fF/1yrvww78G5bogJ4ucR49ZgjWaQla3tlIOZwNO+P3Y54Nn+VT4gdqFACX
hv+ih2u9kCLsSAIVL+jVjwCmaG9TyokJCa2GkDyJcmYvz2JPmKR4Hby5QwKmdLhO
5+hPo4mwkJupWpNqs3yDB7nkuXAh0XsFP1GqCWUAOznD612i/gth6AGc5WbF44qT
Mr8bI7udraqh1M184K/1BByKm9PoU3UPEGT6WxbDsUlTugwyYe4gYc2dpGlsfeI2
vD/ridkfhNY5xZWsr1FgJt5ddpqV098bJBTgZz/6wfgMVPjnMiTqpjYtWiD8iFij
NExcGLIVWkeMh93UDyRbHswvTNvNowdzUKY4NW5wvpkt8z9GvZi3azs98ipDLdd5
7akTmZrlcK0gWm0XS9AwReeheWCHcIMiVzHr8q0Kb7EeJxtPAlPkW7QEMx55Lxfk
QDGt1zNciMqqM5UuCCQwotJPSSrWHBqL8alNG0IVK3yC+MUqP25FAZjbLDbb3knT
K+GJC/dRvbKSYMXT9i87K5iG3P7NRIqj9XfCy3h2q0HfITmQr6iLKVjR+8BVT3Eb
OVnFYeNvt+g2+FVa/gApHEfYqsHinCuvjTzz4mrG5cQvwpH94AL5G0nb9Pn+r5l4
LR2sQX5bRmVM2SjC7dEOfi7Nq5Bf962Lz1yfXuqn7R/h/qorZo9xtL42ZKNlnwEh
B6xLLdcAve3pqwr3D3F3f8yjy5N25+gsctlXL8zzIMW5A4GI033VgFJPx0lnPXpt
i+h/y6OntY0bYFKi71Mk+/h3eWkcHG55B6U86rlyayJlU4CsgHj+o+KI5uOIbOkv
pXTbiKkcgJW9wH53HrDoI+nM6Bpedb4quu1Y91D1I3j4ShY8yyrGcPhx9FkfVByN
0ShRdoIG1VLv8mBIP9irB8SltpNSwXJ8NtfDkM94njYXA2iff3UW9MHRD9k/7aV4
YgGIqjJz73RkOHU9SsNFyKcoW+6owqwSO8d0mrtvZu8Jmc/NxQ/QXZ/+i5qwdtXh
KVOY00XjFjoYkH9/cQOJxezowh/YdylbmBY4BGXrZ1Ioji3SQRgkhQkNN36OVKcD
pcAHJLqwUeXCDrjM0rx3oZGNeAdy2G7dJApxAxunczFZrPKcpm7nPB3LT7oNxDE1
zbprn+yhbwfNdPUsxzH+Y0tWra+G5sKR5EN3MoFDSC0UZMbk6bTOqrm81IeU/+d9
InBpKDLukV3yuKc18Ltx6dXbGasnZM8ILEKpoTZ0sXu1cPiW/zMgCI7YJyk8EFuY
vkh+VSKpJpaj08Q85Vfd0Up6eQ0arJ/BT2nXl6zjNSPGvpFK3j25sXjtrLRDqMFB
AiZxjBmd5w8uVRfb8rgQn16y0hpa8lrz5klQctjrdeRQIcdFCplpcQC9pR53UCcc
Lqph41Wp1RWcGIAwS16gV7srktNgPVZAjTp8JrP0g3M9NxB7cV41uYfAWciXR7Zu
CpdYRgPU+fDDT/fADjq15n8W3dtWgTbs9NqIyI18eOpT/uMKcFzs8+RtR/6BZKVF
WjTwwK+Ko6q5x3Aj7/VhtcN1F0QCEu3SBO8oY22eOJd4ZHhjfndmwXp6fadEDXck
eSLpEoAbsHk28RsbUxQOFnZdb6eGTcLxHsg8kjZQo35l+aIbZS7jbMi0XehqAyfo
dVKOazlVlRPbjDAzQ17odvQOo6/Tqy7VZbWSu3/38R0aSvcBgrFrVPCygChoAl8t
0fJ4tK3Y8+dbzOdYrSwn+gT6UJS2LqW+lQZX0+tCZfOXRgFYFI29FJZ0ji1HCE9P
wAidxpuRZI6F00OzR2spvFyVl15zC43trzQPKFY0vJu7kQe4kQJBWNiJh6RlldcP
MHoWlBoVnYda1wjK+qw2pwQXEMd/egaQI8NQL4d1z4BcIi/nUuT3EFkc+bTPn07S
pKSjllFdsFhZ3j8RLev2gtuA9LASfqYtVqf+4EonBp2v/Vz7CwNxEkP8KZUTpO4f
xXqfRgDQNPnn87GedygzyGMER4VOfaf/zi2oVwGCehxGuUKaMRqgvb+ZJqNGYYy3
jL1kXcKtatCr6Jak5Qu0RPrtvEpt5p3o0fWPtyKSpntGTmU2RuOVb/G0P2vdRdWM
dc2jGUOiuDsNSoI0l+clXvnAoTVuBg5PVepmoppuMmHcWWGI+ZEtLOvu8+rtJET7
yvditxlfCFvND8/LgbYYTUdkXd/h9mw/1Roy2yxWgVMMuj4NOMrKyk63VeZSrNNG
ToIZa0cSzrD9ZASlcu5wzw9+MFEQrIMI9dsTYEL4vqQuQpzuUt6KNOKFdk0nbH1i
FhN4z/EvbfBGHJw6qEKf1lKshRPOv6YV1M2MB6I+/QbsNRNXWeQV9lrQMxc6/g+4
M4IPCMNlIsF6BbdBUHOnIevA/DPjw/6bhlYma5m2PQURon/H+OpSh2iJJUM9zaFM
wUgOBUcBsfdXf372LbhY0HSJtPwi9VX6sR75iGqjr6dGTAld5NakvkmI3gPkEYCE
5ahfyOswzWor0kEAmvQnjOl7KgICEHQ5ZEGz5QHogxpzJgDOeuoB3dFSVr9ipSBY
NfETtogDIOKNWiED2EJ2SIhnfWNsS6MVepQyqUO4cCgk0R8OX36gMHjMzjQeFB6o
teaJeDr7+86CUvWzCAuIw8210OXaVZfiFh6PaA/gH8/dbJ2so98EoMbhZutWxjp0
kzbOlqk/GXgFUYboEognAhMky/qdZPFYvyCnW5KcL2oD1WOn6Adi33WpcSuIm4UJ
mfp2PytirEss9viD7OAUfFOa/Zv4SMZeIQvUHCmWu5zES7EgMKMd/lWOc54vjwRn
bc1CM3A7G83Rzx2dDgUDyuulkcME7FvbDnB6N9JdKcFmlUFvFTM7iEdWRAPC+RUz
BVus+80OukEmkaAJQgxaoGoZUVikU2XXF1X5j+USxPUdFvL9E4gKv1gXZgDspEOb
5qtl5l/Y5ixnvFZSV4UjeP1owqpS7cpJK1MhjxlMk874qqwnEqyS1pice7TWGlfL
9+L1Q2ynd1pTm+prt1W5HFMXfvO8kTAMkqb1mRWs8hTv0bBbwJ8DJVCB9Y0tpl1S
bfXPee4tUksZfL0IQA0Uu/CQQLkPhKweXFGETQgdBaILVSfFXuoPXQV1FvF5Ok25
FwwqeIyxSiPA67cNefqHKEEKhXHD9o7SLD7ERW8oZnkfDy9fZ497BdlFZ9Or4fHH
VYwW5VUSc3b72g/9IlaWmp9rMNe8NzdviMaeJxW5XrX16ugm3f6dCqZ4lb0d2dxL
e+4R7Mh9td8x1bioSG9SspdvSfbISxFhAkWMRVZo9r+20n6ITavYkm/xHYYnLUGE
rYGlMff6/maTWY6XNV7YeIt2OJ25uXnT/KMod0VC7qjh6Ws/XFmoJKBneUNK/2Dn
BinwRkMROJ8i2+SSAs6PE/P0SeowOPu/u1KgOz1Hn3m3rDtJdcpsL9SKB1CEVQeY
AqQWQxeImTTPI4En+8A8R3xjY3vfOYtiCspfYjd1Eoutqa0VqSj2FWB7kxp5HVv+
M0eevfIRUwHHRCCLhy2tX5DFZxZfkJh5pHeOhtI9AR7oJQvGsYz2ZPxuNbChIIQ4
3R2SQGIsYwmlrz06+FadG3NBrLduy+006/fB+RxV8GD4dOVZtBdYaYyth8l2cWw5
LXxb0982HKs8X4KqUYDtQuzaTh6KhkA39weBf1pzBmlfJUALXo44+O3siDvxF2xv
0OSwd7Ismk+ccgfQyWvBuHN+1aHF+L8hWt4bYqTJrgL+W7p29qkNmr7yZ+Up8AOs
Mvt8JKgPdQqJjR+pBVbBrv1Dnn5+aDdgsC/4f2jzmG2n8CnWqfn/hoVOAhGA1Y+y
1lXRWV0DPzJsLEvZE9SaSSZzpJ7k/5BrZxi/H61Ru0+6jybL11Z3QboIVwXF8qWl
6PbORO8lsrqMNrg9G4CamFlHi6EWVI0r8E1GAdq6Wt2k9HNuDwvxUC6pHOGvpUF1
nX3H5klK+cYqB/s0I8A/QjnznETwUlZVdNdvoHRG+Yd07HD/q5u58wSdm/IglrsK
vzTGsjQqARK8DxbuJwm2jTJ+v73MQFKibJAY1YTb7aND90/8LXUupFRyg+QfRMm4
FNhQpuvJ07bzEOYseNU0Zna8k1rtsGm1g+6kC2KlFxsLJqAf/x/tRbua6bs/DiJX
Cq7fGxGB6M2qTQCIg2hMyhy/tbg3A3TigyxOnnRpaU44yHKPq0CnXCG93SEi7+Pp
J/FEk88W79X2VwC502Va4eUG20AnL6bOqDoQ0l+6LAsHr96hZJdMM6s1SzKPhhAp
3Y27LmHPZPqJ2gRshLkkTfVXQa3oKlK5q0m9O06qoqm2tNr0npGsxOQ4fln1V5Qm
Q1Slre3IFSGLHYPZHn0Ji6XETERxztlXhWOQKdxu63SBx7SHsuk1SH0E0pQaSdQ5
g3dq7EfwjFLpqvA2GeteeMovcP342zjq/nFB6IMggv41CvPf9ggh6sz7hZhnBX5+
35ja2yIIc5S8EZ5JgxGKNHUAK1eXJGn9S4AaJnZ46ZI+cHq4cs2u7JCRD3ZWkQ01
EqoKw9gw5e97sNZSs2b1jU0RCCK5S5IqgVJTN6Ahhe6R+Vw9HwDTcGkOFwPV00BB
p8uQS6MmZD8Bw1pcH8tM6xfExqEzK8SOpfEOEDd7wdJscrCOBoWCZ7UU3Q/AiKgK
thrpDY79wRM9ET619TmFyUo0CGl53ScKOusbMJVFwp1xnB6XUU+b+39ro/LCglCW
LRZBLPs9o8XpK92GSgOQD+GUgs0CAMrT150md2022rHdkztwgy356V3RUyxYHGe3
EuQHV8sSE1KoFWxsl0k7MxybuVKWf6+sNlWK4ExFPhcmjKlLbnX3yr8oH234bBHy
oNE04lQ0jBovmn0XrbA1wRBzmjEUmNHX6BwsBQS08ZMaqmTvuqILxaGIH+tFJuV8
NSqoOl3PmW3MS2NMzj4DAsXa45POsir0OLVB/WgEwus1+wao7p+Lf65wYGVPJSoO
rxu/m75w1TJua+N2o7++D9WwAWvCtQE/eOuozBvYkYnKn/3eNqqOthF08kzrheXK
h4hTcRQD6HTvAuSPrhY1vKx0ZQGcCsQqUBIG/mVjSvViUUbLUjBHHaUUIgRzuPUF
+WG+gprvVOaMowjNTfM+nyt+OMitj6rKS4I7wjT1uVY5g5Q60kM01F0sQp9kPjhv
qXDqKcArEvbmq2AR1Smc2CZPvKxyF9ouSTZjvsh81tR4EaWiS+vZJ8JsXJ16wUu9
aEPqA81D3il8+LlH7I+VUTAfSxHmABrtFIVj9wp8C+SbrUkYLssOJZY61ua2FQ4H
nRlQCkEEx/5gOnU6h90rNSmOUCuB66W1h1ADBEUpsYTdqysfE02TilFdTpEsigvV
0vd/+/onVTMRHr416GE5NGJcqdQRTO8L/TBrbMDzfDzEfKoJFH9vIecev+wJoZdf
P4IAcBx9HHEUlrrTC7mY5pdsSRyHOaHY8i74QMPhFi4=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hebxek3V0dVVGIDwNF/aiTT1+VJwkIyr7uvReNDI/SSU6fkIScYm1lqiBj8F/Exf
j50QtjNfBREAiu7GyLHzfy6URI2+7gTHlvNd0prOSbZ3QdXJMd7KvS/hEf+sCTL1
6DgQ9hdjkYkiSjojgdZWeCEAcE97Zfzk7I5ZrPoEqwQt/e69vJ+ByZSGUHmTVvRy
Z6B9ZIoUcZc4rWkRrcjvs7Rc879UyeDEFzGOFe6mda2Dt2MBzSLDaH/6zfMUKOGa
z1nEc8S0ReP9jtpgEu7WiAyAZf+i5a3pnzvgWsgP8kMfS+u4rkAwbHq7hoR96azZ
pIbzDpaawZwzB1U69y4txQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8400 )
`pragma protect data_block
Xw3kKp7oSyp1o/9wBOKyxpKMcdPvRZbLL2ke3D6MhD5YahZkRR0YAttMOxxi9Ewo
C5LKhtZlI8WuPZSgjlPHGDvHQC0MaPmFDne1g8yxxuw/PGW4JAyDnD5+0sgYWDvb
mXSgYAakdL4LHWTDjhbXJ8nv3p9fztCTzmcWYsIJAvUdpzbMvhW7T5y60mTxIXHV
ztK7e/AbcDhVOK88FlvvWN0uEOTLEyATaJicnQ9RUzhtA3OL0seh3VfLjkgk3f7H
y68y1/3RLllwyojmHj85UJBpYUxrWKKnIA4j6eEFZoGdN+Da/6ule40Bzx4nW9uS
xtmsyS1jl+/hpnUwYvAvfU6CcozhkdFA3s4bRsYAFW0IHpWaF4lrCrZb0JbgbShj
44fjFOw4fAG8Ovi6l8xmf3QQ6MiikSdUw16SCqK/TboN1uWMAQctAMUSAOJKFd+e
vYqLqU+2xG1m1PFd5qnp9MFrc+1On6/kD0Cja5eZAheBzepRldpRCbYH36EdXIBo
Amdqfl2sTRt+EdjezPjz4LBtZfN2VQMI+rbJj1n0ttmzzdW57tkYkJ4EWp7b02Lj
mlGRQGpE8uAdalzcQLwsKiFHV40GBCghGHy6ulYSL/nTj6nCc8hrZlvQD05Q4X5l
KSFWQ8mpUKsW1JWZPpXOKYS5dUe/pRCzb0hoQlxF6j9xMguji0b5P0K2YDdRNtQf
CK2ELIba4BC2EzTy/H0jsdNIS1IijWKdo9Ci9TuMG1IavP4jsp96x7FOGAMi+8tU
tOnZleHAycYNZhhHYq4q4EIPBRnFErGdSr+pFXtbHc09AhApX5/90coQ3ev08/qj
VAX2L1ZzslIGdfi0rt1wiP/P5k2PBXKFFT2VPaWTW90iXLQa++0pccgovoVnWlvE
KdBz6y1Wv0a2KzvFk/z96QPTDC9ZCVcnP3Y/FT5NvOcS7T2EsLd/gXZUf+TbqKxr
ExQRw996tOy0XQufvINY/FP06aXNVTSp5hH2HLcXayNTah5BT+VTD16ENCr272N2
oqndFBb8pMA3eixWD+hGebbpaPvIvw/TyVqjlgLDocJix55h8Vdg7DojBYQ4EhsA
sMyPBovrIrHtui4GECaqOA4CTCpDqL0Ivo+ewdn0XQM6DKze4YdCE/rgq6/eyEkH
Gy6yW+nWaWnCIy6oikHbQnkxTFX2ihAKmkeXb0heMNVYlNA8ZDt6nCgy5fxnmWuK
kxI3OMDro9SFdW8jYj4VH2tOvJAnYjaeEBO/Y2dyv8efmmAs5Zbf2iH8qPiFpPhQ
Iw8N/6Occ4UZSN6O70zlbDn95D8QcVr6gEuki4ZCAmOuodbhEXrwK+rCvvZae/cG
Uyibw1jIV0/N23AG5kC2C+i0krRQtYwI7arTz62/NDMjwLi2T8k0DLmQo2IJTPDN
EoIlf1l4W0yhJqpNA3rBlIR38uabRll72icc4I0AJAzUoQfWnVmqBBOLGzYTwtAw
ji6vvFyyym/AA8SYvXogEn7A4xbV74P8CnmpFTacpvlKB66yilB0jAYOdEWs6jvf
uvaQTGoJ/VWVKId+zi64Y0Yulj3s6DCVdVO4f+j67elqDA4XG8W6KPqaQ2TZkA1Q
reL7kyP0pUL6kCyEMpeIRj/ATRAGw29l/N1ZO71UqjKC1oEzc1WuMBGArleWGfNW
jAQCtu9B8veqp6UJUHYHpr9k+DqRUSxJ0W3jA7VHvpct9FLRGrAI5+opxpWkLgaN
ZFUczQAteXBppR1VRuqTyIUTN4ZCf+EPZH41A1//i0UaCjX3XibbRVAVOit5vqDz
SFc4tv1W3lrEscas1WfK3arrxSSLqxZZJkUcqXvox7f1TMRFBvVWH5rC86gqI2Xv
T8qtjnxlb+tuSqdBEOsEsR/M66O2XdnR/wh3FKDGH3SHVnvuJE4UNavvMfTbEpKE
Fng2aQmmNdu0U9PL5LAlzg3wzEGqBDVcWIyffzNBIfmMbjdtq/Zq+cjNJ3ZxHear
84fS8PFGfGWa9PdT2pqX0vVNPs5tY2H8syqCD/Lx5cAiFhyZRc9mgyFPLCxP95Ns
G2/dMr2fn/0XEBC03T63hLqWgzGvk0gFzGUe6mSpYArUWV0hkoc1PKufXaEvo1Gy
TwcXD8hoenumOoYs1EcM/XYl1bWWH4QeFAqTn+T64eVF+0St9tj52YPRGfpBd56O
IyyGpmEbdtFNvfdbpCtzzDF1P2ppNyXKWTqy+vWdiYy8MTPjYdUMCc2cxyxMBwqg
78BR2hacemdpPfgmUFBsxh+EXnPHzLGweqFZsOIbYrB2k4+CLpeTUqvlf/HiKetj
4wNi+8zhwVLI4W4myNH73mGiT0zFjA7HepzoYi/W7U6XojFSiwBccLSHexWA3JMg
mnSh2WPAA5oFm/FzmUFbr+ScZ8qRFTSolGwLZ81b8pQerqYQFOaXkB2Cu7nMHsXV
hxFAavHBishcaudoD/lQ5sBsBp6sFzVeBP0WGoaHNW+RLQLQfZK/AtlirvJpWPl7
oKGma1uE6RxjHW8yCAJYx/91Z9gNHPSR801Jpk5dNQnTKeD8OI7I/kyIME2n1Hr1
hZe0RfuERH5e7ZVNw8SI3BSYsUWCjK8bO9JCL3V5abjlxjzg5Q80DrAx3vrVF5xN
8OWcW567msuKOgtu9zpC77neXTJeWY1mevc5xRtggU37qi66jeZg8OgMntSCpGIw
RQoeCOhGGhBNpO7HkQUy5NB73Aqbj+Ka2/nerq29Cjh2wt0LA2tRmi9GkBoaIVaI
tUGrYuKytgFFnEkoLcryGPOdJ0iMDesx6O+vnF38bJm3YH/hzePsnhTeWjQc2WUs
W4KQviq7uG3SP1gZkrl6pP8qrfG+yOlqzXfaGfrh87rLUlLbH+MwGWMirkgYO1J5
TW+zMlGzx0/1L27SHOKoPDf0WZW7aj33bnh5vm0WF+zQccOYgif2mBDvYci4zg8f
NmBNXvX51FXCRsuLzzdU15oZsiPA/ZaGNZQ4pCz5BZcMUgofkBG6PH9R+pmSS5fX
sZi9I6GU1ZVMjz1v2DrRAGm5KZI3EUeyQHvsHrh3nRH8gIT69rVMrfwruHSRnns5
2lBheZKU492rMZM+uyZbPTuvwNEOcy+kLtX23wNPJeaagHjTnPI7Lh4tW/W3f0QQ
xGjFfZISNp2SH48Os/C7xSpsoUjHBQf+FZ2+IfZtfEQFiZ5tlINDoBT48wPxkc/B
Oy5UG2MEpsVQsPIj9ECBFP3JSTA5QkykXopdDI781yeVRS+PTx9/Y+cas6I5w4uh
eiqEdcWoOfMLw8ZMRdInOazXfE3VpAYlgeW+R/8iq0sElOJbCvnzSTI5+4tiHEhd
I4UoUqec3EoftwShP2X2Nj0oboGiNdyPW/jgY00Cxtew0HQYnIit6miwr7054vuJ
78GErsWjt4d0qAtAmCz4+W2xypo8j8wuVkmC/mtUwAReGLT5NLFSAzZ8pa1NBGqK
jjy5AJ8Y8/XetM3HvuYF5IlHd3NR29E4L9NWug7jMNkusFS9Q2wr1jVXRH8j6qMy
SLiyKR7/TtqQZjsw2i/2iTlMamGq2xJ79GHFczsfNha0xRT8llAdG/BWjZlaONMc
botDUKnkS1wnsc2aKraXXJTTDRas2qltS9KR9Zz62ANkJ0E1dvKajbdMkicsFGvm
ttQ+CdeknPlTqvMEfYQCpuUWeUjHpKI37T7eb7aty202QEk3ywXOl+1GExZzYhs8
SO2zbd36ekzSukF5jJtqfcQRV9n5VE8bQ2o8LQmoubA40zu42dNMBN64tfnrVPir
IwOQ2GYTQ/iKeUu6sVp+LsHd+N1yGfYPqEatvtalkk00/r3422jQ8GSo6W4NFWNz
JJ1u4WDFot+GCCRmGDfXBQOElv3KvgHYwqgHcRTHCrXRsBD1My6prmBxORkJoQyd
eXJ5qWCsqW/3CCxSz/LaNpffCQLv9SYXeA+y2JOOz9UZIUGUwkteRDiZY7rgXDQ4
fAoaftPiLPhzZ0lzeG1tGDmqenxk1TrXpyDBBrhvWws0lH4yzNQN+cAOIKMYrveU
aLWPsuKALx8iz7WW+goHa4UVYx/o9+tJlyuXTsd9HIzo1Ln09H80/NAttMAite0Z
JjHDklQzsCTBQMzWSJuk50yZgFaI6D8rrkrEOXd43CRNDDcODiiy5w3NZogUe46+
XKYl2suEOcAnLlCFMX72Dmjrd148SgERO+t7dNiPFuX+6jDPmurfPBD8X7V2q9s+
DQp19fB8p4sW72FOm8IfNyusqpMu3HUqewh4yiXqk8O6cIEXiF/tLsyrFN2Yt+Yw
467rCId5z2iK7SxCIKRuRFpxnP4dneTFpK7LY4+sSUvWXmVnvo8JVnY64C8VgBke
amIVf0L16r018dVFO322MoNi31/HOPJW8OLXE0x1oXmmDJjfi8SBOxWHxt53/fsE
/nwfw9wq+7ZuPKWonreX/l4z4V9Sb4lUbBOuDM4IyWkL5QbmpZfRrrK4uQqhf60N
5sgbXPRcXSYCXhaOHoupvHTkK9c1oJ7GD4omgO+405Bto0nNk1dgnFOJbdTN/jpq
nQ8uz+AzKRA+PwvZiE9f5XRFN4FH6HjFRMQaUtXnyKpk6W1ptxnWywrZsIEd/Vzl
Ns93lPAOYVrx9VcXo+AXqvp664hI5kdX73K28ZVMjMgRPulofAofixo1yIrBL003
nfXf2cSyTilnLwOnTTNI57dzCJ3omdUuk2Qc3uSXTX1hNQKEUYHxHMub0htvFPAT
7eECAyjB3X8wc/ezdlAY1OTVVwlPrJnYXzXAP0jAoZ93VmTgrYNSjf5SZer/B2B2
T2mj9MBbvMeYDQmGvWihxRG//G53Zn/GmkI/OquqYFQF+hEPt9/ZwjMDEElyw2Sk
v/YLyJjMPQdRqXyolKZTUvXRBzDTv6yu5Q4tKlaUjyDQ2/OtJXmUht7iPkCOV6F2
SL/vuWZwKc4kkncVJfQLlQUzvohyEGuBfFfayKqcU9PlwMZAQg8yvqEzVroAWcQY
uOWQ2ns5N0Rt1DH0DiEacAm+lPhm4E+ZZD2mHI/DHOe48v69OWjxwKhnrPHXTsLz
WSaFjm+wJTKPsYH5MpxMOfF3/aBl8uwdRSqDrr1ZugCVHlVnDNJ48CEpLxEDbF3W
7F8C7BExLEDJb6vqhRRLjdmW/5n5x128vaEWrdU54wgmpiQmMp04MCtEh5dE/amn
lBK9mSQsPb3vKhtY6VVBKYZpFX/5klAwQa2+vqrtrkTJ7ufaou3MxUckiiwXDuW1
92WrdPVqxdD2Wd5gB8g9iLDuFrcYbdBaEcTptCxth/GSMSW7fd9A1VZ64pC97zuI
Xo+UttVW8gwx4sMWZET5OmubMKjYV6hZknWH7XrwQqheiR7C/2b8rWNkDlN27wse
EN82VLCOe8vFlfmHdTFzOi84RJajTySeVLzGMaWO1UQSU/TXgN9XHT3gSKcgXgfM
HAo4lSOtQ9LIlBaZutfpngcAcmvaHagsVlf88VjBDhiKh51J43mAwRnQilwj/tLM
zmZR0IakgixVdWBhWiqtGC95vcNxDYIewAESDfQvE6Pk8rHCOMpq7Prab1uRFV2s
vRWT1wvlsO+r1S/QGV6Pwv0bmjUtMVZqNdwtcTrVjdpOkwz8VY7wi8Z2ZEGrjCZm
xdirGkLSj2MP5IF+1rPpoCXbqsDi2OezS0RuysFi4wCrsM6qeBjfChIKyhVSdsgO
K7ZzlWBNMCi8DLqOnqbcjJJdJX2v5yk2wRoUBiM6RBVFkn2adsUO8TbYK+cltZIF
12hG1N13on3NCNJph/hVZyhpl5dHjoa7nutJ1GBZt9THJn2qV63Bklm89l8WNTcV
ef80t4rSZw3M4yaPrS06L+LyiwNqxbte1tPYuRF8YjE8SZ4cq6FsqkRMjhTkKJTZ
NafWgiMuX18eAk3dEJtINwYiMSUWWDhlR+oRcsUO1mIsv8fCRAO2lhqFWYeA0V4a
JWjSiQ7PwX7wxwPwiV5gQ1RcIQmir5RMMzEUg72wxVMc5igQ0tpZYgACeEFFwoqJ
bZQbd4OTTmA1zxxd+pl673Jm4whk+6IW3H4zu8kWt1fDs+qEeDd/8sY310NgMTQE
rTHjNg/SbZBtePczeNO7UUFb99Rvxwj9gTNxaBpmJJzsuDPbf4zANjyqxyGT0KE3
9KGxvVblOERuhkxW3eYmUn4Okbp/BNnBUpKI6AwCfJqL/aE4jfO8j9HkUdLNBNUh
crUTwgSmmMuPIPTMA3rID/v+eJRmst/YqVhK8JJA9leP0clKa1pjxzVL0VMLkHgk
+S0Ah4rpnYrXBWc4yW4FiK9aspalYqv862xSfCMxq6qTYtiDoaIJ/1/w9ZnvmVI2
svcKXKr4eRrBenDhnqnnXpbHYxh5+f6mbDYMmp59Y8Io8uWNf/H8znhHxVX5GzfR
I7omID5aZNcSNaTBWk9sD2pAjq2tb5QYhB9XJ+vXKKhEMNUoEqUzLwxQYV0SARJ8
LUxLDv+oawAAv5/aDjafYMt1gUe5f2Wy82b+8aAO0T3eBmhD4PxftqhLVMPIuWAA
pbRjCgR7QToOhdXhdrx26DpEqkj5kcVpqILJiVhNk4J6QhsHp2v3G2a4ow0ghmYJ
2HKgqHJW0jjXBC4kIeFVXaEoi0Ci6g0gwWLWZVPsGNrlYobPdSWHtUOQCKdIFVQf
2D+T5vwVpdkm+nRp/idsO4hfjzcI8MdylM8qDQGu4Q4yLG4p5w6z0VsZUdCUy4yG
yvmaGjFznFkoKb7D6zsL0QxLhsH7ua/A9tATLryCMfytA1pLT8gpAQKsbdVta6oe
jyWOI3cSYz8Qb8eq3gAQzwVeBdob8h5tqOLfNneVdeAbmG/3JFaBZFJmSYwl1cJz
jE0FFYsoXBHcwr71SPbt97pNuN6MZF8DCgIL1lBWHU5jfQxVkorNuUwIqDC6Wd3D
rWfkCoFO8dUbfUBvBS3tpiyqQp/jGYClvJVNum62WeHl7f7MCpi0CnR3DqEVb+pI
9k1ot0mKAMe7KVsMTQquWyg42uezKkR2C9gi5/gjYa6KUdriXs2zkX/1fiJXhK0U
UeJN7sRdFj5b6eXe7VzGvXddBzlgzRkqrIRHofNXC7D2Ds1WSNQVbrBf9M0JXgbh
MuptNl2twMZvCJRJjwm1yy4CE///RmrAxPxXrqnunWNWEqAs+669qkToYFS06gaT
5Poypm3lwWhjC6cKWuoFSlugBTP6OXZT5tIgcnBhOuy6xhdJjHYIjVEHxjhtMkcs
G4sFzCHD2ednSwX5CZGC9SfOZznN506j9ulULSTazd6qnFltAjN+Dr5OMmDtwYvO
B7mA9ESt0bdJW1tGMi++ClWP966TPBYO46nJgLf9v2Y3RiGIbNG5a6omH3Bc4GvI
D0EbwX8ty3/koKfWxaDRTzHft4v6jO+Z1SYF8YOZuwj8sA0eVnQ6PFnwmuu+QRwY
yHlxl1OXuEjzJRfa95JHXnXzPd81IhyydM2/Sx29gN4fBOqbMhr9PjE1Ki8GOCUo
IqQ3OpD6ftvk3HD/RE0LYrxZOgkdkaOMIP4U1pvqp6zE6uUgiCiF48j0jfo4ilrG
N2Z+Udx+2VBiyUbAk2jSHTW1Bdse8XlrAIAH0knLfvnQx/dufxAiB7wR3RhUpyLy
nMj/JFg1yv/gj+Ersf632B2Io+xo0+4YjzExFZwFx09WDPeMNPLlt1B7WxWYjvOX
ushJYiyYuxVfF1Z2BbzCs6vw01f58NhsCNsDoF5UUISq3/znBQftUx8FB5UmGHec
WYuuS2ivszEDGSm3Iwimoq6yFyiZgFAs83YfAWwBnavKga1EMAxT7aumGWPSNYvO
MnpskTvGFCvr7N240W4uIH17oyMMGtIEfcLJNVE/BLDyQcI5G5I2hkBYtbeZ3EEI
HB08hClnh34h/hLDKI7/DbNwOfTAmTcjDzVY6uiBghjxEiCbiSmqwmu3GMXuf5/O
RM6gQB2hWAuaUgSh0QxHvFbld4PASxbNXgqdl/R4N8pBj3gti+gS6gmy+9MPB6b+
Coky1olGZ4yWhj+sZrHqvazNr+3EoBHQme7vFUF3lO339kXwJnNkMKyDQHeX+rSf
jZgRIGHN1rhyTcsqE+eMB8tzJVxxV97Jbfcp7Y3fnHP8FjTHEuZlisealXoVr7af
QoOlz8Ak0QLCge3vN7DsOz0eXcZH9p8DYMDKkbGm1qzwtml3E5cKlGzcJUimuQXV
NjPmUzihhZUXlhRXsGPVFVCMbtuXuVBB229hIgbXNwL5cG5/wPwWknUAB7ekmRBX
qo9sQbz0Cf8QaFtYZ/dAxgByMsZlf6f9ACABDK3GaIqsJPLMF0h4ydDtj6JV2okh
LSHuxZvHVeBnfgBySltFYws3f7gf41URSmmaJipV2izoUg2YRem5EkZ0aZLcxrqR
pWUcOnW2c6SUuOIekSinRkRXg8OxOpOP2mnPCt4XvJa0ND5jireK7cOe9FgoDTqh
UQw/J9BwGLlt8UpKwg1OOZB4wNAhgKQMw+LuXnNaoTB2lNzDmV/cZsPBN6UlneWl
7Efl00eenr7uZSS1iyanqPfwqXq5f+v6QnB01eYk6y/WjaD1JInfLwF/BrLlboSk
Fjlj+lfrVvcfAw3lkDEFGVs3T7R8wUbi/XlmAZMBXLXDr2yhVMpykYbnaacQN4Rv
moy1E3g7Avc0vu+qDFnW8lZIOyQj0trjVBfPf5fV2KtRl+nl0SB3vCpE/cNXiIPf
heN1JmsnM2J5zlJIPqmReQa3ioScmT4vstc4d/YZRio+ib3qNM3Z5fRovjxv8xZM
fBE8IiFOOqpoNWpos2Z5NFcJpiqjkiVXog8b2mKljSINtTBSqT8A7M3RSo/tEgRs
DNUGfx/debgTlqV1ezx0Z46Rvm9X/Td4O4HywZ5y2VU8lY79xv+X+OS3FIDxFfL7
JrnctX3giDfUhVsgWbbr+HRrho0/ku7Sgo9t4Tg3RGPZLHFmeb8oGdlW+rmOJ0d5
xLT4VIJIA/MZraa1Y3d+1+76q9ruo5l4S1PPt5p5ZZA3d9Z93xI+H0zI5cOkgWiL
H1NKq2ojw681ueK9JZOVG7gVYmEQKSuLfdC72KobFdAnGA+Mm7jMdOdPkW+k2fOc
ratDeyVGmHiCKIeQFznqiQE7pOU3fsAZin4KKQe9hvoshI1RvHPoa2/UDWeC2mqb
fX/cJ1VwOLKca/EwxgYLIVwimuHWiMKGI6RAK4n7ZxkxvhR0IYypBoSM0ETVyagQ
yWnBOM3lNkXvGrRc7NNbCJ0lfVbeFO0vI7Assl14N9J/G+2cO59ctqB0AsNlwnpR
fioTDIHPYfJuOZnGvzWR/mTqO4IQwmkmD+kxiyN92EOGJEsJuMkljjtIKHcFG6XM
j6kbf4AMQjrdj5+1gsHBeptLP4ElLjao5JBdTlVP7s59q2KM349dAU/UUjVRVVRX
t2eMftx5/QLi8wp/kD8luHKSQkkZCz5NdH71hZuJqWr9ZX50ydRLlsTvZFamNeGE
YpD6FVRhsa1hgujEb1Rkq8ti3UHlfe/oAnA+thSLU9wkk/1Z53Np90eoksllT4kX
O5MvlEkPe5xkDeAM8Qyjo+mSBzXY34zBAGruaGptNIj8zv5SIsspKv355EkeTZek
bEl1V4wxkxQia0LDBUAx/r/qiQ5z5eWPqvXuDxlHL0K6e5cvA/UOUDYLAoQsY1tu
gsIxOCwHdZnm8AyAKnk3JUNoDVdf3X5dZVGnI9U3pBjZI2HJYELvvvn+5dIjEu+3
R9kzC+SocRmSO8Qn1TgikRZaXdwtEozwJcpmrA3k5aiMkjEMPcoxXCNlTB+mUSrV
uWNv9rFTIfntGeN7XsWpdqslnGecRmMR2Uj8bUN83Ym1W9gjJU11/p6ohL6K4h9q
rYcMGj6RxU/tNQizCtn+z1BuuMM/h34ra6XAAqvrzh+sLh4daw4yNDwew43qkRHy
VSYwmTdTD9sbsrf8uHByEHavqlBdWRSlTdOFPP+/7gNpRlv/+0fmfSI8uaKbc+Bk
9Q798reqCIUthO5LnxPdE1FYA2oegLJGnIzKlqucMqMtM59cx6APE+11hgxvYKdx
3mF0kK+9oenFEHUna5LHcwB2iPNEbp4Bo+lkDM/BAcXzxwIO2g+qfuInVKxcjISn
+8ncq+yfrTDo3pqwLRMju+sm3DDj72Orh3YlcTS7Rf3nCcnZ7Kq6u24RX0a4aBcK
t0CJF1TMj9WOtsPEk2k4W2ILXwhfVhvXTT3k3D4wy4Mo3ybiUXXrxNgkFD6Or7xL
eRqJI4sKlds65VAhZGOPqifJHY+xpFDVNn2MnUX6lPibqCXysKbMdG5jbA6YLy+k
Pl9z15D4DZztfgb/YfERTHyaKa0cNSXKg0tt/iOca16eWRPyyCbRjNmdR92V+dxy
jMWXgU8cbDMyWAmZ5ZhgykE8RgqWauEENuQDi+wF6tksFVDB8tayF/I/sdFzxHnL
XldN/dk55MJUrVkNz2xWdNxKjwXQ0x/jOAciu9asVjsYm+/FFtIIRzkmnrA89T9w
ZC8SdR7Fp0aE/82DCEcpnTA8tM3lQwghPBNOJ7qIc4yKa7+rlhmAqwISXONNJrBM
OvrmzYvddzfcceBXZevF0MpAAIE/hUBVy3VsYHdQCLb9px7QyYnjMo0m8svM9CNv
HO802itBNk8onWolyCFBT/43lZwixNoM0ZIxeb45N6R6BwA/0mcQomrTZAvt9FDO
0VrpgwRBEKDt0fvOFktHUYI8EQ/MqsPnSGNksYQ8OhiZJk5NEsYpmIl3hH0QblyT
oGeFkxK0XlIPQFTkCplHho5vFatXo2sOW5ofKXcfZUEFxy2WQsleRkd2Gli5qpD9
5WPZHVsgXOb1CJig5ngYwk3K8trxQDfyG//EuY3SO5bV5coWGRwCsMKw17+qTIdQ
Npagj3+8sSnZSjZX8M8uP9XVgYbN2AUzFnpSQobFyFcWiJDSr9Wsuyn9EbMnIa8c
0W4GwoOsCbRcqsrT1H/mPz9fuNE9V8wSAZRTW8n18s7CxcgUUKhURmBJCzzNcE8M
vQ05vVXrDmaj4WwfS/L+NVo4K8q4EOFT5uJZf0Pkb5jXET7i5faixnx/g9reGyLa
f894vZ9m/hC6OF6c1lbV2OcS9+yERsfBXKmKs6Ay4Gyt6QP6wK/VkFaGvzKaoaDd
FdD9k8+6/t9KxWa9CSJw0zIa9eR0ek7M9BAwd7qw6pFuroKGbxn2M+6Ts92d4f/7
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Fgqs/LvfA8OsF6VQiZy0xiiAzJVJLen7w4T1t7EbGjY7bRd7rdjLqi7W4i7vHqvB
ZqUIwrVG2xkqTh1EQ83yhrhjPzJoH6qKZRiyk4oBWDFYJIbxTga+DMj6rjoTRt5o
jrJ7Cq4nSQpn/xrR2kPURBd7kq2uZHukmByLtzhRZthwPAknhi68X41xPrfk4iC1
ExoDHsyRkRziIOPumWjOfvE3a0tmt31FAUppXImo5f9WDsxpy8Mk6aAavelfNUL4
vVMpnNa0K5F0KWHYeIFZbRhEkXM4m4riD5uQajGTe372TjLrspcxb6iP9bR3PJFL
1PYTrOPmNEOngxmFO+7QOA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9280 )
`pragma protect data_block
6mEELEsBJ6Rwv85C9LEpEZctLvs7hBS/DI+pYnwKjH3SMVdznNEI6ePWNBkXCYRQ
w+GCUdbDgjvQ9n2k1PQqUJ/vB1ZVLppcRfmpPSsJ+4iH/7eDea0nBGhIwsR5hOG7
EbRCKzIUSGz0SS5Tgn4M75fDxyOv0kZIlAftsd3b8JJFFIJWj2D6lKDu1G+qPbv3
ahu48wIaHDeoKuSZpM+EciP6tHlxg/84RTtfl5WEmeGHwTtF1OFkvbRBEL6qsbTU
jkITOr1atPYKW/OSanXCxMVk3yYYPO43QYq6fRB5C8rEU/wB3wnI3ELTs5WerlOl
+jnv/6tkS3/uaBRjkDxt/EfCKiiRQtL9PUzlTGuCZ9lABqRUpfGOaqPJPdQ9Bkp6
IKjxLmdV2r3ZD7Sv9riK4WN8kbBtywMudZMEIQTv/PdwbLZXiHgcqdwj9Jnhqkjg
mzJQrO0YWE6Z9tzwaT0fD2yKeHxD3fWtJWbTMcvJw6iUzOPLM2Ei6y7ZUV+O3lIX
/2mVf8saeE/X1Q8D+iL57s8y9TbJJIxK9SehY8rboEThAahLzoQauSt3+Pz6fKzL
ceVLzbqCO5j5LKF/P+s3d7Fz+eIv/OIGD21AjSIcMm+R78YxWdOHjC0G7KkugUG3
Tw61Kgt9ZTV2DG4MUrLh1rFBq1XhvWRE2IFK/5SX7iScFXuFKy48b4YE6ovDCF3E
zdfJTV6n0shCvFGkOXU8UpZkWILnL3BNSARV/t/jNSVNdTeh40lVLvvOpTyecSB6
8lnW8mgqL/QzkvKS4GRm6h8ZN+myCDcZdGaN/VT1+i5bcuGS5fuGlRePSlt50Mk5
La35wm42E/VSdh3iNagH82yT7LibQi7BmtMU+x9/u+vQ4jTlH1+twknjjiAuQjOt
1t48uF33q5dO0mIJlAdhZOYPOOhXv4webM0qlUE98OaxOglzUi4i9ql9REmxTSH4
3ERSvdPiDlu5wMNBq+cQBfDT809DUCprqxoXt/SWbzLsS5mXgCPwdVXVTH+oOdl/
GkFzORIE8COvjzZ5JG9WVIe57Ym4C31fm6TyB3gpOvU7ZF/b0LkgGp0aJWBPpGH4
Wm51XAMqURN1EbtWGCTMQke/SmJUf01q3JCF5eDT3I/CvpW3CN6ZoAB/wPEZKIJq
Nlek5G7VtBCHntn8C12sdYwBEahayc+ayQH8FtZZpqqahn7ygq6LnJvm9PHYizBf
b19pYO04f1ItSKTzFWhm1kAVs0bIAJ/EzmSdJJl+Sg2Ma0PjfbFb4JWdRvKqYXkH
VDjrgVT81xnC5/ZPYK75Hs9stz3eVp2OTrqtBpPDx4r9cIJEtADc9W1j0ihZz1NS
5UPJSZX4Uoi56zburIyPRvls79Zo/6aqGCx0UcsQEDyL4FWoy8UhgAe7PymwwPp/
yBrMsc7kr8yfxtkhesiRvdBCUEiHdLhKWFUiExmBO355iUHXXYh+qY8Awhp4lGut
WeosYCiwaNW/2CjIlbpJVRvfFCvJwze4HVAksH05u2qkbfKGbdCm9b4JLHUOnvou
0CqmYNo4jumV6m/oquDoxMDVHKSNmdfC1jaRC1tHztrobeeTKvLDw32LhnkJNuPh
n74xgR+9SHW+leNVbMhhqBAjiCm95hRO9bPo0q6kY2C8GPp9DgkTNkmV3MaDHWOn
53jjNNTlC0SOwb6KEQ12l3hofJ2OdeCmSIizyZRaxtUdmD8ZlI1IFsSQfzXqyZGt
jwikc14S1U5bKJkijUs2p47BOqpxfLTADHGDPpp5f74zakuJp0iHFIUZOUThv30q
iug1BLmvOkv1DnMgs2xkwi7dDRz/BHhCLTngPvjPSkdYXZjSVzRhdXLs49s8sLXg
oxrVD1kuupPhjoLmRKNJGs993AnoYEsV0ahBSPcEyldTGHj6kcLVloizu4nDt8hV
qVd3tbZS4LQNCBkGHxa1RUgDwmMLAyBKJ22285kwef7h8ix6JnPl0BXyoe0Kipfp
WL4OK3HIafg21PbvGIe6Jv2b6bt7ybMfOYWQRclhgB7ODuxMduaqofZVM0S15W89
6z0LfJWrUcbPyQkKi9U9vPEaF6wfkjFg/tLwLQFfl1tNP4et7MHtZ1/PE1wlkyEi
tSN95cd9CLl919sH+UJHS4vU5qI5cSo9QWHs5JgyODtClYftDPtf6IbF+RmCEzTY
fqRFRC0GMG3hqXNgNVK1abkrllpfkPXSSe4GK+eOdKrKHngVMEY3mGQqGBs4LwGa
z05LymeXGhDKnAQ1VBl3Xrt/4weC2BbUVEXHFF1Ko/0ai1kWsoUPgOCBf7ZIrlWN
s5pmfygDBkOHEyuj3Si0B56oD6Z2+qjhZu8O988S4kjs1QCS3uch9pooriNJNDeR
/ObzrTCAvhRmu2TUMQWSTDVMt4CWZHcVuONhUqmSyQ73vgBzYfymGv4QOtxhH2jz
2ps2egMa3qXbokAVoJdAOsi8OSFgg7cwB+8bp+M9W4KGMcs6noZe9Kr92of03sYq
8k32gjmtYKzubQbfRQw5O5KHZ3M8ahKGwi8CeewhjitOxuDfzm8b+NfdicHt1gBW
ekgaGPtpeBRvuy18ScIrsowPvbGluYJGZZfyFeKODEOt6ETF+PG9TVZI3YC3OsXa
hsFa6OyZAjsyvpqZeQ+T/rD0+tTixG4Fu1y15KpoSwWnZeHCopvbAEiOQD97iWPU
R0pbvUn/oXe6XhLODPB4q4h72PocXFNCwkobmKItM8ZX2xJM3FVsDuvTQ/3q7xOJ
Fp9bxBnKLcgYawYUSXGVRTIbRNI7/4VgHKnIo/fqN7YAwYCTQcTef+WKqu91XQxa
NtNWWkV4s7uMGpoZhzm8xi3PvanDk9IJC428tv+BkZHeDIfeI3IeboMhgKdI7LIX
GJKazkjIESzbyLINoKMFrB0ezFGeuqZEbZQ5t3PH+PSPSmlhNZX5VyTgv2Gb3Nul
V+cGlMl/zAjnAhJ4zCYkj2+AOzkqTd32tHZL78lhAlZU/kwAEJELETe5JmbsUreM
M0g0odA2PajdR/O4GX0NtKpyqp1srT5ZqXEWoWaZwjG8L77q9M7jX4Z18ByoooqH
fareL+6fupsVTGJWiJbnP5vIbwnz8EX6NECJkvS0glah+p6ue8XQdGRSM++/yh1i
Uz/yTJfukc6PZelz+Q8dbalx2iccVoLy3T0cpPZx6PM5GI7EJSgkFURejbb6q9A5
bJRZUNM4kz7pss7JlpnZE+IdtmqTuGO1r1Rb7OqFmsXJpf1GmfjelWxyIJi8xNvP
WfJFv4YnccNgOd9fLYMstUjoevdL4/3KR6O1ExaHZ2txU87OWtt26GeNW+pt5raI
NqREodjYzpuxu1r8pMOHd5TkvFYPzqGL4Jx2nyZMyvXE9h/0UdaPY78nQQFlQYww
OmDDlaFpMvnaUnVP/l/aYw8hWO1XXOcozxXtPw6424ET83kuLzWydoJqC2lHTis0
ZmxBjhfhcM8kF47ZJF8TEyYI4YTL0IGe4evL2ttx+LBIjApqdwhFY6YL/NCYGHOa
uQAv9vTSI8Tx558/WEWwy7ttGFR3Q7HQskb54D6x3tUjlM3UTaboaj5ug4D+wlYj
Fl3HrF2KcA2nnUdPD55yKbt8CQZjchH/QIRaIFMgOuVGYrjABw6rZW37e3+tCmTn
JvWXejg5F0FBIz21hXrleSdISmPnMd/EBLl6KM2pPrKr3mlFU2azoWxfGFPo58Fs
gE5rty39n5NTn7KYUcdPqg1GdPC85O4a2uAI2sIIpyHcgnMU+JQ7hG3scfA6TKyO
luM++kHyqjCLNoofVgqyazvbN6hHSKHr91Tc95/JaI7asOSsCuBQNb/oyUFFiIkA
uaASSmdlmIpg/J3bSnbw1Gn3aJC9sVY0w99A3/Ehh4uCOfMWTFSNoEHy44/u2QjN
J1mdSApEZO+lZiZ7rUO7z0bMd9qOXgcpOeb6yZPsFYCm/ns5b0GLgv2uNa/AcO9q
z6g46X4g2wYg4eqjun733wBGOuphb2MNAQXCtEvyseQaEtbF6YsWBa7B3HOiR7xh
Xi/1Y+GfN+GkDw4VGTfmfVXK9/mHf/wdkkas/5cL9AbrW1/G5UD3kt9pBtxeaP9P
F6TlSsh6nwH+V1KMB3iHktRFXTs0/XQPW4HahIQwJlBPjmmaWNI3hxbIvm+clu4q
EVw5cfwx8SMZ2VwPDAD2+ykiLSE4EbE6AVztqnaPkRaVABbI2I8aWcwD9aU5FIlM
78YPMCNtGhfw3QWfTYu00Ic+WOyPhA7zC+VfhhxPoH/MfW0UqimzJ90zLVYA8i5M
ycsLN04UWve74Prv9ZrCopYC9TwcvVPQtZQdF3nZNRoygbWFqKTQAa8Zgfv56nR6
GXwBJ9D2TWoutxP7nNUgF8tamZxBdM1GN60cwihun7pchis0aVinfYvqG6St/mx9
Slu0S6VJiiFxGreUWlyJetQXINlFYxl7C81y51PNeoUR3IWdt5bdPkp/ld2hbaQ1
DVOefNwFyZnhKFp8DAjrriLjFseMRYUrN11MPZaaVSifjIgZmFp9aSFjW1Epkp0d
3xTMw1nQUNNKXPubrBKhxw2MM1/k3CxAugaoJBCy9DhSq+DiKfC5ODYozsMY7Qly
mNMl2/XBP1lxxzP0+CKvKTfClvYnJQoX9sukbQs4Ck7/ZEkT2LccUY2pVFmf5u9O
wa276X4WCmHpJRB9Z2CpmEWLwV638NByFxFGzCfeCTDjNA7NFe1WgxHwPZ4GVEbC
KSQ3Uc73CSgMdbE1xim20UJHKPk25c/CB9j6WvR1+/yGuwVzWaMmsnb6KPdzYAm+
UNlECJLpHc0EufMIsyBcHAqVenbP+sq94HOJ81l1KXeCq6nhbjFf3DtQWJpDcAtT
81RDhL9vu0F9V64R/rHRtZPF1ZfEBs2B4obUlktv/3uNUtC3RAE/CKQkvRYOlaA6
6VC3ukbUDO4h5gcfHsl36QTTm/I9VQo5Iquq4kb1WRGtz6TsRswnxgX7Xty+pNmU
1hNPh674M8WkgDZTgtAxMTT85t06Con2/3U1RXFhKfuRUHzDvlf4AkmSkmPHjE8q
b8XpIhTxl445EZp4Fkh7gJS96L8iZzB2X3carQqJqgrkh0lW112ROq9krQYvwC7j
Hmg7Sjxhbdzv2O1MwKNfrrP50Cj1tQJni08KXgJBzvWrwxtPimeYQNBvg8RlBq21
umn0Vu3Aa8w6mm7UIplnvMwUCmShV3MCyLjw8L3zpCFsdgF3LjRkq/fgIvgI+xdM
6xz6TMzg1scdTifECOyu/TmVQ9+1kqEU5GHK8kI4SL6WKCHoasJH3Q0KwZGuilJD
slu7UbDrVyVXr+O0R8sZoX0cZP7EEH2DkAFfvGcWxuEMuRpbOzBC9I01msH/nqt6
30aXXfA1HDPytiNXlj3gFKQlwwB42lTp6MK61brhCDypCZ1HG/l+Gzw6DJILKQP+
Nu8PO6uIuSW/y+p4lRJDFYZYW2GV9LTq5r+2e7lCbq9RC3Th5FYQ9xqlbOtJNeN7
+WY/7grETl2F6kKi/wLEnohKYd8UvF/6qHggKfBl0TCbA6YpU8cZlw8+YIGqW/Hc
rKGYdIz63tpas++kuAMrFqb1Eo/H4rfdvxgmAlMzNlAgCjmBHe9BB21Njnqc+2uB
TXAn7neSFFem/wFbhbVYkPATgiowZuZa9ZETdtVlj3WnIGtKS2z2qCzLjHJDbttM
K+W8izeDImsYkFwNBUh6ZqZ2WpK6s4AcQwK1UuadOgerD+wnDzFicGtblcM1oU8y
TL83BCRy9Ee5Pp/rDyMh/ne3OElOHT9rr9+xwETlitDKXz3IrCKNnNgMzPoan9GH
jiaojQmCbED9VWfm8j9wL+6VlwZFtG6Tj9tntpKptCTjunYixd6CE99rvfBWiFUU
Rahx+BW+vVfgOM69wD0biD2XsznSD6tqyBdsqjwI66hQ+Id4vMa9r3rJNjav35Nd
qB5XjIbG1Qr4lybx+izM8nRzFL5Ith2WIo/8awnLPmoaOpmzlMxnrPnoRIxIw6y5
Ssj9u/NcX47w2/7HRGW4gjMqcGahDby82PeDTx8Oa9UFiGI23+5lCXL3AiU3o8i5
PN6OHgOfrbmVtu8LacuSzbXd3SJ3Myriz1ZMDucIWV+p1wmfuK/KKhm9hzJujWKs
w+1CP9IOPrtmjlaZa3UwWJGIO59BwcnATbTIX4bVArd2zZfQNXcpzfJhQqF7dpD7
3NUCDQYwsyfsQf9v+PpnPQHIZrxJQ08l6bwOHFU2B20/HM9nmd680ur0WvZ7lpiq
KO3BGzuye3aOSGZwEpv9Y98veYADwnURKJrVm89NbUEjUixmvCVRwiRGXAvFXFUk
kAAy6LeqSg4P+KRpe5iNZqkLLUGozOU4uolqfW6zEbhl25UJvaXp43khzvjmFnKv
VaakTbOP9AtbqQNb1R28u+A0gpv3B5nXmXyAAzWbs0Wj6ip/TfF0wrZZuzYJKVNp
CaIqeNvVsIdiBuYqjVOGKSogsRCyM5/GTGQBr8DDplgXCAZ61sFjSFGxkZZK5/+S
Otn5E+0JlzTpt9294WR/BGCmzG43jFlXezt/jaV5Hfjp1/C+EJ0qnkYbRGkm2JI5
cO7Lnp4WOkpyHqlvmy6k6zKTUVSQSPdKx1BvAQIVdTIbDyUgKuUEY96jSagvWkfA
33Nx4NiNfEfS5huP2Kp8Ms7NYpPW66Bj79jps7+nV+CLblUZz2H8ZMYohmLvmcoV
vMI5/OD9kwhE8C1Ii3VLNdb/TUxO5ZQo/A+7dysITOsWKsmOEuFl/cvt1dCtgZSt
iSx1hre6uCPh/AzvD7LyX+Man7SRyzZpHJj15xBfb2LVH/LgEAz2kuHgopgjF3IW
ol4I+eio0ASL7EYp7nSf3EcP5Nq9ZKlK6rDqTujx0NvnQulBfHhyNuoW7Cy+oLjI
yYNCoWd4nlWwgEKTHb+1eGT9XZRISB2j5gnpi4Higx7SkaSojFTTSrgjUs4CZi6F
D9D4xHr19ndMTA8SzeVwNGMQGdyZOHBssqorRWb27C3cAaBWbBspf6KY8N7W12XQ
1pRQUpuJ6Ew5k8Ts9I0q25TKe+8inwoPDI24swELWSydDUaIY17CFas0Dvu4ENVk
kaP4PXqbOohlppVikIVw7o65yEn8sypzjrYHMx8wQPAeVMoK4QO9cbhsLdkc882y
N6OU21R4z81zYtbHL33Rf0QaMVgowknW55htdEBT0JgwtUj/BMMOHh6VbNhkDph7
zGHCK+2McbuEZpGrjGhx/NZWLb6Vv/6Km78y/xbUABF2ofObIoazfpAIIb02Jzh/
0CddKfJn8Xpk3uCT6p0mrhBsB6HAzOlaCBMqAn7pobndhZ565+MTpPTV/tGLKocQ
n05COydRNMkAYvFoFxKlrDTmlaLjNMsNdB8CgkD0yidLryGwKeLYJQNrb5BmZrDM
xqBpvvjCiHNvxYxA5KRJpY7vM349WA+ZgXsemKKKNwaunAIriMFie6YbPSSXZLHR
RCfyzAZjBNtw3exVKIoFG3DbatGDTiFtY4b0qadUwQXIYVmOHrFfTPOuCF4uPclS
n4sQfiOuNrKD3onpiOAY68Ogm2jMp3ENzlvSvBUndEK909fcb2PLn8D4EIzNNUaz
p5CaSdcur9SNlDI0sO7qvSrE49/0Klal+/gF0SlkuD2Z9MAjb15nuLa4Iwsx0E1P
mMyIqjgqnwnNJZNdd+5uTvtnqHJb20R0l0FbvXPMKCtA2LGUoxD0KvId4jMEvN8w
ZQTZPh23OI4Nq+WTHf8XRA3O7cu0vSmqBL3XCd1u933ECn7yI/P7JamE0/7Q6gzK
P+l5+gYyjrjN9T6VDLctB6DAbGqjhE0sa38HWCacKo6MAit6OpNXPLRxbfptBPKe
e0pvlOP8ehV/OIB8UXVXcP9dRiovl0jqcLrmafqgawa0o0pWpQTXEjOPVgCmYITg
AR1sifEiX0n+USDR1aTeIVaJ3rLWeZOf3o0v5yTll16nWo2/rwkWVaxiIxARNmaO
EEBFF5/jDwym3sAKmCIq/PZDXTBmvSoq83ubcrh6tIevNVrUynOQ2exOx3tiwh8R
dDHvuPRGZBvBkP+8e5m3pG+smLF2DJXjPKyvrtpJ0CuauBQWy4/4FqXTPhPeZTpj
838Sw5z52WKo9eu2UuuPA5Bo28FIoFMfnsEi+339nTNyEZyABrSvV2jBOSOWb7Xu
GifyE5NcoqnLUpLEdqT58Q+xzPDEPywu/Ywoy6RBRsN0JcDSahthGVIF4IuUf/dm
rinlHRhszc90aTLgZNb79tCuhjqxdjJ3L2EhADD2Kq2avNOkTYbFNV9AqFqEf1XU
1yozXEv/w5T3vzr0Hed8l3D4UmZGIB1+xjwyK2nmXQZrDnwn1kFnRj0LCbDuRxOs
naeow+aGGYvGwxMS7v5nZ3SiADtmFbv7CbppnkL6zI67aM+Q9tF/sRkFhgSRF8MU
DjvJ37mGzioBaacJDJ+6LoJvIhcWoqZ/0WAFuR/crx4unODtop0PEnH6L9ieAynB
mIWPZh5XSjCk1yyU4zPk9sYU4Bt12EziMvA8DMXxttz8UA6fWy6BzWSji6kSz/UU
9bII9Nu0f6lIOI93draocKSIBiU70uECE9v4Ad7tH9GKOw3SrDdZpz7yRseACLOf
8C5EOMPzGUr0VEJlDVRr2cJYhbw/jT5t4IP4Sni2Q9Z3foBR77UQJTgeyI1EFLol
ppn+g/jQX25chHsRjw/380jWOsN3BUFxifR1Sxa0Qld9bN4HIC0qTL5U/mIXFGqh
uMbrVgbZBrVe5Bm7H7Sww6OuNsEGaATUCEBoI5RPkuhzu7OC6BTfOWiAAuqFaNXD
z3/Tl9kukvsAgsk7Pm4MZUwlJy9+aRibXJ04rK/wBohp/lNf7tpNue7IoVxXn0bd
JkItZEjtsRXjW6NYBr9hcPaM5cbAZS2+yasZ9FWJD4d9gxvClTyZp2yyMPMbQoD2
STo1gMKKGIosHGyTMdY2dw//px8IyxcI0uDjGWHzIuYC8WahERmlF3bzMUHyT43J
ECVVbjHidwV6pQHmbTf4jHhYmp74cKi3jYzVWGx/p9JSPKCqLRZTF2KWND+bhpom
X2smlkSU6+Kwks+8+IWjjJU0UdekzjdaLZ5ZQYgFPE6gkLF6GOi+lSRQBc/ct2PG
H+BTLawmJ2JV8Ga8IWmrwl5f2XjEGDAwlbAWHwPYmH6CLajEUm1VTI1ATtH8peWa
/D5S6Hhx8klWOBB/88+Be7oVFxaw8d66FwUI3f/3XJPTn8yYyM3c/SOvx0IX8Qnd
Hq+k6RWPkMnQ9Dqz/XR3jiUjEEGh0X6q8KNs8bUQEr28lt37Lya/IMSsx2UHsJvV
A4XkBIPKmi5mO5UUHwgiPgyINUNHPXKIHjdzugRfFx8+ZQHAM013APdTnFlwj1ck
ZRe5Uq9se33pSozhlU0mE2psm/Q+ukb4Vm9hcdFtH48vd/QJ2aTxM1NY9R73yOiC
lyB0JLb6yOK4WmI+lvyTdAzryd46BkrONKudZOUh05UjU10Mvfo1nwCqb/t2+S7b
4fN7JeX5Yrv+JQ7QpDzV+7YyAr20WPYgMbpyPjR/HKXUfAPPzig3iyw0obTCC8ZK
2GiT+KSqu4eKRifJPXyni/3u+XmY05vkWqzhwH00XVU/sbEbcdaWq+SFocooceHq
wNPCH+4raywIgunAmfCphJorNkaw6pxzfbWYut5CV4Jrjb3ZIECnf8o7Ztk2soeQ
Nx+oyNjlxlnA6UvozS9twqWtQcg5nJR73nse4QkgWfIkHsKRHN+8x2v3A1JGCbXu
raVomYEfAM9Z3PGC7G2U3CAAT2R3FAnyfqN5sy/xGfkrxm1Gbjo6axs3JTXsn2d5
ld+7KVEchWyB9/YpCNMPEY74iGkyUrxszNWJ3IQD5QrUszq2LF0aZO6zT6TuSsZi
BwAoXvJmeL3XEsu1Al024Dkc0VSOeRT9EqYLyJVFylZGd9xAgBSabHxLedMBNJui
21A6UFsYf0nJzpZwT+jrPmt1mlhoXF4oJMbrHa72OaE+XSH/TAPa5/SAPOOLGb+n
YZWrCE0jsFucMCGS7W27Em9+TdloXjdQcVlDZeK8ffYKXDRHDRyOAF2AXV+tXs7U
ttMhIGC9RYn65mTnSrUP2bqHa3obR8WZobde4PK0599s2WtUZNT8kW8uCaNpn4ID
69DoirWQRqj/rpqV4tyreymMD+yZoQTxQAtlvUCfYK+v+y3iLcBCoUtZXf02hEIm
XL7+d4YnzcVqxW52B8sq23iNWTDINcK8I45ZrZtuhvnQYLauWXQJxn3BQ2JaKuWk
LAC2h/yfkbWnTMo0Cpo9HFrdObf1JGK7xkdr7Kk2aUTaygW6sJwl6LtRoVOlrdRb
nzc6Kp2JowB67sbfYnG/98YseDB2MEp/5YUqk1h2PuQOlkDnR8JI+Lj64sHQpsaU
HR9zFJwJFvVSmMf4ob3n9XxkBXZt1bTEPCmMCMHVx0umABIHSOPmVFqPMrujbDHq
5RyOGnkIOZhCdNxstDrg3pGkqgst8/DKDhfI9becAqAFM37wYybXPhZmq3tHJZwV
PQ3GbPxUQgJ+WvtvVzvgNH/vq0N8Z2Bq/lwFkTgwgipKRNiSs6J8Lc45+q/3l/hy
w/+z11Tjzllwa3xpVniMw29TvxbjfOHJ+2pSRE6R3UX8YHxts6/Db1/O5k6cGCfO
FT9M/3OJmE5DjgZZE/AtnLESrdgt2qaJkhLp02YjOlffeZaMur94gViSzgcDUfB8
jJojgK449gqZKOYQjiKQZsVHxYMGH0aaMP4qceK0nM2tjL7I/0J1bZfYHpw8NKZM
f7YtMkKDWdWqsthdZt7m9GhIkhFcMrwtl4NZXihMhfH1Crwo2MFTQODEj7UD4mbe
Zz2/tBlrTmDJxWsgNivAzr1DQQp/jBjYAcWttFRUCVG0iTBK1MwGuAPIsj9+7Anz
IrRxnR3i0dVY0hIafzp2oNFi67Qsx1X/mQ5REjK2z/V/LLJdZG8UY04lp0TV6xn0
4A2VCaFMwj/R88Wnc65TvzqRs+bIhbIvhabrFFenOvRx6OubgHovOiPzpsAIf+Nh
Mdt6ILUvFL67C0ymLDQZCiMxzC6fgIJDqUy8BcQNB1RFJzJkj/O5hZ8tJ0+6MKgW
E9cg14vIn/yP4U72dLRrp3zZz5V2S+1Oohev/DWNEgAxm+WYXng3zT7RuUBQRuyL
GIElERq9i8yygMgPR5OiOFgq85URA6MkNJMN/2h7ZPnR3s55gRBc4M2+pv2IgDTl
m5+mXlgp4uV5FOmLTTWdybFb1rmnRvCY33ObVgHXqh2YHVHpNl0bnxYBcI7HHath
xcYd3LKAMRC6Mb+Rc2kCNcsbY1v02UUyxRNFe2X77c0TlpGH0QQAl5At7oVYh1TN
6BO5/OKs4bM3FbiXa9rykq2RCZUClCtURye9jt1pZixpiKhhrFXkJsTRAcTr3lmy
ssiX6wVnj0JZXIGMD2QqKDm2S2H49+3dWZrtKonMebhdJ4qzGHAQFXvTeDlgSkKL
Ulul7co5C7H0UUS5j3k++9Lv+RyVwgcMqPCvh4W1acR4PVRWLd9ne4mHkscUpOS2
cdDB6rhTLTkzDlzgLmXsMNk5QGMvLDzGuqj14GSYiRJgAkxVkcU9h3LBPTbBgiGA
HCoaGy3fOCHkds/9aQC8+C6BkMt9wCTnwEWt3LMx8QzdR9910/20irGKgFyTmCEU
CzPEEyD+5kICXM7Eczag1EYGP1DpHGzKBYUdImHuEDykzPHOADFl9QsKGiSQSiq2
xRzrA3v1tRylF0zsDdBNfj0bYaS5fIgruYkyAqj5hT82wXdovjC69M26917MKmBV
elUTs7pqprgZYzZm22HdkO1KJ4gpjFdit+dk8zkl0okeWnQlB2KInrQq/E3uMChb
BSlICieKGe16T7qCB1yEGCK3OnK3AEodaevMbPj8qz93zrgGUkSDIOj2sAAhwJ4R
v0MeGUumeu9q8O/xsYYOqPqaAK3/GCtJwjy1lLnmRJofVkWCklGVMnHjuMW4R6XP
RJcCJUD2CapP+EnsgelkWK/+lA78eKEXkqEWddBbJW4NFfC6YK5R5cHDrxzRMCB8
SCjENmXpJckNbP+QKM1sTpeyWinR1QRi77H2Eg72cjStjPCJEfrKp5mq02fGzr6Y
+DugMXJ1dVdrjjNqYqZehwqCJQTgbZGBRBYJwV55ZrFUbtqngFctYV+WaPdFr7oG
mVMmxqZdFZx5YHypY0aTfLWq66miDMHNaFcHsRFWoUDRyxHJgmn5LTmXp3dpIjKY
lEM9xKr75CnABts+nXefhAh6uJtfZEjxL+5IyrvlkWyGCI7uURgj1xa/khTAgZqs
yTMY0G9XBIAvNMSbP+bEGQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ObJ5bVa0Sgv7NY+C3u/f8VJow7ise/JRO3pe+QsPFPEvAPxgqswyrZJ22gbX9mrE
zn7j5ONoX55ay5jzRoo9xw9cT7PnLu+K1YJ65Pbss1vPcalcOwlSjg1ggzBiY2NQ
2A337zAFghHdoCo3tavZ84wdsmDtbA4EXHRxH3iHWVWLVyirWag7HjhFsZ6N6gzF
MGYX3bRqcOTxYLQRVAlYygR4X4SVCV1AeqsT/vLHeyfl2kdg2yvBKsIbOSGUVdrg
17YOivsJ4cVUENGv942dmsTuBm0oJN8w19rUcldkNc1eRmE17tp+oe+plHeTk54l
ZCvM4zI/z3WllFW91mZs5w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
3qbDHz7VirKCV356im4OiRe7j984iA5p6kMsReGCv29/wZBOY55FaqfvELOVNePE
eoXSRwGl8B7rEGf0wAlnFRvcx5KCs9EZPixpn/kbRVf/jjPieEz/nQFLLJa2MbuI
kOOZjJH3oq1bFk0JGFW37SR7w9RsslpsR0eFJ6/W/qfcCi4QIrM/07Gqw0t7ZWc1
AvRj5IbEBMcLEVIsfF4EpGqoo0PjQ8TnTk1Bsx6zOyKcHgH1KGZNQaOkM078wqNT
+Chv4d9ufqnEN+Upc8Bt/DIAx75tdGg2fwMxmn5LCt+Dt5un773GqMlT5PPVsg62
Fy3kOlcuzeCjn/AciQSDCLiQ1y+PGSRaoxUgf53PxtF4eAYRsp8az0dNWKn50m25
k3v8ho5nJU5R54PSNHJ/o7T2pCHqRe+c1UQBIPKzNfAqAi5/ZAGEbwf4aZXoxr3c
iFB/QsUAqAarRs5UDeCUeIdu2iIfIjrHGphkMEs9ftQxwQtFwPjH5dE0+5BuyiHz
BcuYHQm0AX0efKujKDNQ31ejSLjSCjPhvjh9+1UjdXIrSrWI0jI4PG4vkWXpWFct
Wq4qxXVtdqMROI/t5TxPZGo3lelbYauZp2ew06kWlUzdwqBwMJf0J5pxtlHK4JXA
LE/fauiXAIW16ZPiq4GL33bEsmV69jHM6cMssEh2udFW6/wTgHXi/Mnkr8C45hiL
818uaCWs0BwXLuscQPuOv0NFm6tIMWQPn8s5wgwX3NH+KYPaXF4KnZDfJ7V5V67s
MT/V5JqPAuXuRHnf+4XBsvfbdqc++e7C2o0EX7FEPdn5NfIrPTS7qLQOOSmg24Bo
r40eSVnvSBHlnUYMsTjqFOD1uiMv0CwmFOS0+xOT8nklK4BULGi+L0axZMq7US9f
SZJQx1cmx7zZ6u7XsruCFhdHPY3GxRN5cwVRGI8Br2D093s+JioWsVl++ItHDi04
RRF4RMatlwtEogHXMnMR3VXQRWN2GcnFgdywyuLoqV7tQSMS6pXGMZcx+tdvNbnv
er1rUEreY6MqBaDYJQ9tpmBMRvFVTr2xIBY6DgWNM468SOiHQfqB67G7QtlKUUIw
k0Tr2PLxJ+/hpN8ThBST1KW1JmbHQoSTspQgK9x5STx9MeAUIA1aJ9guUoNEd2gi
ZK9eVpr40gVSR6mQvI+jue14cLdeyNyKKnLCZ0xilZfXruk75h6rPaZLtf87+CcR
JmdkaxXu/xdU8BSzFwjlghDVZiwlAYVLdegnsFAv/xoQMm+Zg7r3ay569WcgaVCr
JOBfk+IWN7vWmgO1l/toJCOVoSKgmVTUghT/2OZjhsr1VAaL5CaD5Z7EOm+fT2DD
sdVlLKo6oSJe8SoOCgMKTM/njVV7DDevtkXxXfYgK52U8uSgYoHpgWa9AhUdwUql
CdjqaoeTp3skyOA1cbyRuxalwjGirY+Dezw759F0VEd94yEWJuYIHtNHR3epc0Wg
Pk1EaRX6iYLx/fBg9GqmhxFfyRii/ePF8qtDOK42W3nZrstYwo58yVFIP470HJGj
7AEMANN2uAKjBWGqBvNDmjMMnIvHZt52gw0VrGZUPtd4Rt1VmPAcFlk2FYcpu80M
mjP5OO7O4564ZL/BZQAwW33h/7vqquGJI5/YoUH9ujHcrjNNOIvz5ERSpPoTqwgU
jJBxyHPk4oJP/+MFShT1HG1xFRUx1Z+Z45xHroXo7YLxAF54vpNCdNI86YQNxA3H
pcmd5lLN67vbQNcStl9kg8ZfnFzUL4eROO3CLG7BUxjQ43HrxG313nwDptPibSR3
bV5pofeYWm4tkF7bFk/Hfpey+ZXfo3fQ7ad1KbolZ/nc5WEsRu1oIb9H/r0giXJ1
hIJ/N1zdjLZLbxk7ghCkB0675yDaJVkaoqaluWM2tFfBi/K5+YTKfsmOimXSCPmN
P0UAUFZY8Xph7yQlvGnN+r8bJBitwV161TObT3nJm3i8IUm5hp3mwHuUjP6NaOhB
6p02a2SCpz8AxG6I4UZg+YHdM4mf+g2ZTq2rUafjLxrJDIfRi106N4KINnZgamR2
DddeyZP9YhTbKksyOzKVRzytIzFAvdpnZujTS3q83yWSi1L362LeZxjHTgcfcm+K
SvXuykfL8rFgfN/kg8OgKrYS6zjXgBJO1Nh4nEmaQY8sBlwJsa5wuw9NqupjtFTj
MR0Mq1YcM03ZugWivj+jxAWLpyJ7apwm6fD72F7tnFGTYRjZfD75aIK6ma7v4e/4
zEUmd9p2SeHoQelqiX09bDgNokE/6SgwJyUZDWryNXV9vu/wpMiKb//ii5tZDW8Z
lNfheszaImU2EeypXtY4eV7g16qiHzurtElIwJx+HyWY5RJvMrJEOhmE5jpqMoH0
MmIXFNCeVIv3pRZskAuJA3x9gGCZXiKsuL45ZatsxjxKLaKRuMDhG7dqoI9GRYzN
jXgC1rETcTMouMPjBIFxnJtvXqsLblG5krQYe0WU0LbPEpvlb9eiRaUxy9U6gnKw
qrL+KIsd4R+9/qXSXKxv8wyATn9G8+MIAyn0SfxRUOiaPC8El6pL03+fkt3eJu5E
CYC/NUVvHmAiPdAxJRE9SeYacv/QWCqHo30uE4UrY8KR3mmlJn5XR00amQGD56tX
v9UwPzotRg+1g1T0Ql4Ey7/s1xBKcI8mbzBYSRfPNk595EHpvpoQfh0MgD323Lb3
4o08sG7O1SaPKe8EyNrAeneuEORplAi6+IhyuXxsxwkq45yrX4HB1ME6XAIV48BU
L+zvWCaIzu6gHqel/B/+fYHl4YlprGKTZBWo3rXptrI+zJxQ5Y1nvyKWnBL8AaVR
Ax7TM1JT9gIgbCt6Bnc+mRwAgopPoOmumYQFYWlh4aTJmuvyuwaMcle8+KPL70MZ
oTUfHqy7qBzmAlwvkGUAbr3PyqvnF6mmLw6/gD/oaffj9HAg8C0/t2ZsT9OAKrVT
Vq9D7CKnQ8YheaI3V+Fe3W+4Aa7MFKha5D55/TdqLYt77/TQ+BvDcqsUzb/rsrED
5tfrDlHNkgpWz2dhnmbj3c4mIQW57NfbtbMH25GrUFtzdkmTSfDDnsnV+74OB/Zq
LaTgnswA6aZ/97y/rFtpuaiYBKQLQRMjzo97ZVmJUGsrDpyyC89EuDfrZRZKfzgo
uSt0pmFGK40OBCXqUBA1gGQkilWqv8DsWWhxRz4VYW+s+guVHMuB3tpsR154f1i4
2l600bRkj0UbPEGxWXS9X9Iu+DDu2dkk/JjRjnO9szmosYguO0HSmNw3F+dxR+aa
KtsH+t+O3PrRLGGLpVa8mGJP7kqLCYp1GXtD4N3HMTNzK2SBWwLmy5Nx6JceIvKr
nuS1Kse0o95XGLGb2SU3pEk5A9RdVNxELflmBLLvku0it7UzFhzP7juFIChOewbD
TqaCB0pLJuqDjm8VmGfFKQsZqJIjSDpQpRzKMgzTYudNrZb771GIudwReVpFHKOm
PKNvDxmYemmIFbAHWXRA1RMxRJtZF8RTyAaQl4rplijGo5IUGWJ8xm+ZTecnq6E0
nAtSL3q6mHSlN6+IMa1J8WVrCpTs1MnpG/W8E61BtOfb+mUjbCvoUdx8zyAoJRr9
qU4OTTf6E+WQMJcd+hRj/oK/AM0NcQi/3AqDRzp8CHJ7k4jtm351tO1THuZa7fuJ
4MqqdQegxPHwsV82710MxgHmIUIrUuSZdG6X2kmQzXnUtIsX6PL0DlKhnm9S6wt/
G8H058j/xpMM0KDhj4ryIYC3ZY1ZFaYAu6SLgq51RcOfZ90fqeGzprPRzB2EES9w
Szq0uw9zJOOBDjBNbBYS+sM/OpaH9tP54TYbI3b5LzpB74jGvClMJVHkqqlKGdzF
HPhn7LeVRMy8r9744P03aIGXqrXcOHILEktCe42Mo/L9A/XpJ5dCZ+RvnkZZlpJQ
Zoc/CjGBrMIt/5I3eY2LMrhG1RBU2QeXhz8EegKZqr2HT5E/WZLMySzRLBx9tRWM
oACKRaEgYAVdp3YosZ+JpH0gP+7CzEOzU/tjqj6fQezuJLkq62zCj/FHKL44hToY
Dbi4UwYaNVM8zcA9t1+eDxlOJJPHC0p5z+KKEPzgSGlVjipUgeyI2+1aOvPBMLCg
wjzB27gdTSkUji8KMupSW754O3G4Zubo2Pasm3giizW/bku9SG8i0nTLGNu8cPYQ
+ffWHw3L3mcL+X4JZ5O9k3EHFslgPdb/7BgP2H8fbaWDVd+gdOFJMky01oIwFWRj
6HjBt434W1nWz644wn9TebU+N8iK30giVRHFxeXue1Hs9xoWUGHe+iiN9gBaMt1v
mL5GSnrjwB1JCFyQRJhv48P0rRCgYZp7Hkd+jDce1zGk9l17v974U/eXmhkekvpy
AbOTRxOX8CSSxA1XbhCwoAX++2vnl0reJ2yDdOXUxiXo5La8X5szSzDoQ6VrwOwT
4BhQJ5+eVjQ8ClF4Cf6ZA+2JdxluSNc3goploS9hMi3p/xeeIC3P30+nt6qZIjPg
nDCf9pRuWoiiDmlOMV5UNit+78Oegu95TnzPpUHKShWj9kq8l8QKO9LKXaS8J/2H
HlvQ9u9NRaEj70tujT2HpaHZmEmYI0JclM/q+3+UhnGlI9ljH7+bSLDn/2On5sSN
ZaF8uz+RsiDqiFKbfkEeehXtyfzL1/dsYXsszaKmUE1l3OF0HHFrOQHow28GRNtE
24QcDlZw23qyN9jKZlmAHQoJUqjtR2nWrInfXNme/hexmbaNi/DbzZMDki7krbD4
QWdUOPaTgXIRjArc4V7vksT2dIkZtbZveAOoKOZr5kg9MMwj+O6J3EbF6h4zKnIu
W11Bv2xN3L15Bc2xhrtczUpGGtMrEK1H890uqTbFf0doLOTWfGknOlvFc1vp2Has
id3qKqqclGEnVAoQGGfj3V63z7NW+W5gRpdPrugD9ou1qpOHkeUnEP28AVjsHuck
a4JQHDvj5gX76ZVeNAqmmHUtvnbOdsOfrBgIZ1ja2BYU8Xe4rtCktSYuvwIizrRX
n/8VnXmjqSt1158SYPNYsG5xc8woHNADgF7kr358BJv7YK38dtiESFsdQL4DLN60
YSZd6kgtXgIsXuJHYF/Wwu5RBAXtJaNdPjCJZG6ZLuZNfkZ12E6KR9IeVXxnVKWn
b86mTmuiicSZ2nRl9BLiIPSUtcNVWqEJo/fbuRU5c/UCA9Sn51NvJLC38toPhxWM
PRbFHG0vVrOmdb+cV7jyKVQ2Sf4vW7ZBQsyhkD++nZhpCQ0m/DdqrE5n7LLSb2Jx
B674oGvA/FmwIEERc8brjVrFD5GOA93ETGShjqs+uOO45R3+PgRCS+Kz0KTODmcR
sKfMHeT3Fb8dLru9FWP198x0cQvPPvm2ibjTfShaEndE1PD3wJyhOL0FPtD05Em8
S5wbVSi9FP+tDeZgQmavwV7ScwZHD/6b07tOtbFld3fKkDwo3eNqTc4K2NerBexP
s96WtYvZt8d4okXWHA0UyvMJmLfZCD4XaU/PGMoWkr5DBdGFqjoQfVgHv2LevNed
wkgWnt2tjwy9hHsrbGvWwdXDbd65FNwofi3MiNE65FpzS6Gbaa/Gn24ziq8H1vPG
880JQBXvn/7hYHb0Y5DK2SQYr9lRvb5DTM0fCfjKk8NleYpHniyK8X8/qB/+8si+
gn3gaRmfg/QBkOko7plYzmJ374dI6PdLmyzamcWy8DX2Y7bUNjPBeaDsQBwEl6xP
ugFJfxu4pStTO8RGYrs9aAezCfDjKnbcePIt3ZACwliPP0HZPQDyDb0WhKgb0SIs
KG3r3Urb7JKLpf0WPcSgHi12F7chtEQcM4woLEUAG8XHhpltvAOBDzKeEk9CguZE
GSr73M1Fu8dGQr6DXvcM5EdMKI+KVjo31gj0dZwL4hdkmv+4ULA8KA7DQ27FStT5
kezDlCTtsn1j6yxGV5gIot4PJWE0yrd3qiqMbB2QOUy1LiUrKdPOTqLunROD1I62
YGm1qbU5rYrvOs7S99PI9v8PSmJRBIR+qicw9BS4PSLcVZOPJW7hpftprm3SjS3A
1Pb+/pLc4W+bufOa5V+WPHBktsEQfez+s2aOqTT6wzt2FyfhyTMELPTDmK1RL6bH
B7s01rtk78elBv1JjBQ+zy11iP3heddbuoTGe/wAvj5t7aUq29/GJpTVXVBk3JYx
wqfkvXYwoojcog726b2nYiCJQ/g64uwPa4rz1PoI3czimHc5wmFBidJbaO3cc0FV
GWNaLcCBx24BKxPRi2RTosi+r+9rtSz46sC8wk8shIqLhAk7GaHx6KA8ICzU2hO3
z6h9Ron+LhGB9xy8mS/rRSKG4b85ialdsgOWLsIKOU7Yx/6GHXcLTF0xG3Prc26g
3Vw6FqZxixrNpfIIfp75klDZtkxjBHPr/LaUfIwPSPnCkxn8Aq60VsOKbycZmVOd
MMfc+t+ssi8OnQmKF7Z5B/5dNIO1uN5a0BoO3ad9Ufv04OSJxmK4sAM7Ktz+hGIL
0fLWb4oehK73KGcDl8/HkQf+wJmkuIxPcPkMWZIVqmZaGeJohXcddeEuE9cEA6Pu
RcMI+BbFFB3XL3bG/aSkENxQ08lWROuxnyfoj/cbC/BATchz1VHLp+UbsUR9koNd
DX8qOqbh4zEz8R9upqWi7Ts0c1Qq0YgHTY2W8FgCNqeE2PiJHnNzGCXZthQ4NKKh
nIWWk2oguZO0/TNNuNhT4HfPN2EVFvUD40VfWLvnM2dI7uP5kD+QiuXZQeU7slS+
sSvPtZQjVpzybyga0/lw+UHY4PVVXrqpvyw4m2MOWSEBdCg/hAHvbryvi38hdqd3
1rVxNQ0mrLYbRaTcFGwTe2+RZg0V26/is+WVSkjBIQLlupzzUYH8lKky1OQW0gzp
pm+YIMfAuQ5MdyGlMMcVCArFguesEqFP3EgxrmjA6tDxRikMEW0QNHR9+5UbYHTB
Xi05qgIklA8bwkDzYvuvujNrAuoqS87rKrpIwHrmcZYgji/okDrI2wj6HoUOr+dF
I69Hrj0Jdg3qLJJZIe4vNi6Y/L4KKjbQtAR3ORb+ho8XifPjZf5xqrgiobHT9Uv1
46+TiNerM92wbfwOm30NKNf+oGyeRir8+O1zGQKP4oHFIKaG21f/Q3EPD5ivP4+i
FsgXjRB8yJMvcJqJC1QNLzvQqTjPlYmkgvYU9nHpPernD1oiaFVoZKqHJuGg07mL
/x2y/u4/HDCroZ4aIX87iGp/9J2UJel7E/T9djKAUwZ3Yd05BwEu/Ca+QaScCs1z
YvmLYiWuBFCN1kYgwKfkT5gZfWFJk5c9UDa00a/gzGT5+UzQSZmLh17ZXBRjTn+S
Gd1ftICK8m7nYHNBxRgV3kVOTqRENxINKTZWrLCyfOErKqxbI9LhCQ3GoMa1Ir7g
3gDJiw5T5g4l71MEpUhnLD8u/ji/QCZddv8MrLSgEC9RjdZQatOOKs3DPYLPYJga
89HzfzAR1HlB5tfqo+Mt43WrvEXwihZCR+74peehVsbHeRv7gzB+Oxyzxdi8KcDZ
If7kaADVTsbhiqq+vX/RGLRCb6cbnsO7ZDiuHqX4qJbTFqYkxblE7gHbFd2/5AH5
QJdkKA2idpnZ3niCCQG0izntBfaQhe4FBHr04vvj5an10tn8Sp8gE7FzarcQxOez
WmRYEmHBbgqC3MiNCOHYTKjqlAUshyraQyesPRyt7IYswUoZSu6gk9rMxk7Opxdd
rm/Q3yCVup7MwqLpsMdLH+nodEGyS/GO8EA0FD987Eth6s5ZOnyn066Q7aNCsWcr
Ifp9iTkH3OvwANbfnqH1pk5ICBtrPybBB1uw9IDFTnYzrmxE4fk2ae9E3Uvf9qQa
c7QYT8QaIFnwj7U9aig2o45pKT3O7dKwZ0d5sculCRbe17Eo8i4vwA2rd1UZYSh3
WkD7pbLtax0Uq5RWN40V0e+z3o12bjwGZeQWEcS9dsNrqYscpVVlgtD1Qki7vDUB
VpRG9hOcf6nx6Y9V1jmPcGoJxMD+mME/cZEmJM7SlQZBZ0pAaKl/nHxDPTgy0qTt
sGMfj/WoJm+YI4bjel9mzQDM5IkJPUnvqjKHnKhpPTufRMxqANkhgOEuHG0RHSL/
d7hKNOXH2iqt6sVDpQwIQdMZlHIQHAdXMwZsA90P8I98xjeEm8AejBSkz7ENTYuQ
+35Rk/FvwONlikbC5FKBLWiQSn/+iN+DMcku001wkHIog/lKeeI+ex0yQuXZAadD
UhRh83Np4BTYDpTn/lAgV9mNc0YRhRjiFvAVhU/gaDDtG0GuDklQ/8jrk54Dwt+8
/QHJh/JHVqyexWkhACHAH/G44m69+lKJiUROd+0TreoOo66XIhlBjmf46PfNylDS
29EteFiScPxPW/TlfOVBWwn4zor66TjsVArdzm5w2V/DU/tw2aHzZ+zHhVSyfvf5
T8QkX0K323q/jF6Z6Jrv8qivAgetFsPOTw/tW6XWWhOdlQul2hC6aMBLFBC+412I
xxo3vAeCmGOM6H5bf/VcD59IgXxwmbmaizxt/zRQa+Gtx3p4TG5ebAVs+3+9kJUT
FZ2r/SfcRDzSn9ckSmiRK4Km2omGec71zfv1UMP2bRw0ay2OixAnh8H+gyWwxrf1
uHT59qlrMX8/1sP+ozd05Cv9RKYddNT+M7E1EiMmKIDsiLpggOTWQdAatf0wqtu9
g711f1CnUoQaAFtDyasv4/l84eqmdohwN7yJZgWzkfJR0TmMyt5Dwu6HMOC1nEK9
3Bkqiyw/vp+G97+rBRLBeBVV9HjXfe+E9mJP1IVJKJs7QvCw/k7YRGzxUvfdzTmG
Q69CdrJ75m2UD66fXV7ico/IOG45TyyEcMNG0avBf14xjPEKVabgRYbOQ5jwHn/R
NjJswn8DjawCIqwozd9jyFH9r5bcXR924skVE4WIjrwU6J+AKypY6u53gFDeXeKX
NFSAEelDDHGSO70ryhSEWGDMNpV6KiZ6husAw4gfz3MzfAodwplihBmPzB46xHl5
06uq5/uLBsm9On+r/2HrIobj9iqt0pXvPRHQg8BsgSpWIjoLdRa9+mJit6xIPimo
WLZtRIl2r25a14AZfIKmqvLBNZW2ZG6SbO2TXacwoMFTqXoJndCiOcRNCaj3K0Fp
F56yZf1kXdJp1bbSTo4iuk8En6DMPl0IsG26bw5jInv/+itGdA+7LjWPeNfkRLS3
5M0wR2KjGYmtnWSvh2qNNLOVCRmKOxlEOp/ZnTdmq5bShGdP4rpm5WgMW4P0P7jC
CXPm4h6OWvpK5tBeRvz3NNsnxqlaPc3WG9ZCBp6nbjTUQJNvyu0/kD8pX9wttRN+
qqMSgP+c0xEl8MANeuod3r0zuIj8EzTdYXR5IMB9lwiHo9JwBb2/VrltFwd4N/rw
Xsaaa6op/rjidcX+AMXdwheTYmqYykelTttBjtWmAB7ytdOf5bykFTaQZ98WG7ca
v6Utu3U1w7sQ0s2FJS6KG7fcw0EigtXl5eL+7Kn/uKytTx3qxzmzAJJ1cp9C0Us9
ONC31WRO2oJ2a6WA466rYQdRnqzTj8BhwAKwdjeupjjaJnyx4Tx6F9bxFV0l6RjQ
ZruJjHsabP7x6B9O5kvdX5J6l3xlP5k2kFo+WCOYsO3ocouWrKf9cCBJFe25ohlW
qM9svCHklruO2fuQeVl+DiLRdnvhV5wfJ1IkUrRWMonBsf8ylQG9fUoSU38v99cY
RhkM/KbAAF/98gUNvyi3W5S/uPDoOuZaZqD8ykJ5VeHhrsetGVdzbkVRMzMuV9J2
QLeRT7cECdLcFodbb+2hPkbEGAG0VFZBjLhMOO5JPAAJpq+lvmum5uFlxxkMVZB+
CVp2Vr0vV5MaXXSIlfECIAt3s6PWe9AKHd4vqETZgsriYhmWkolTlG/i92+RMSuu
Gw9ZUSfSOIa/E39wL43sudNh6zeJ4BBkHOy1z6uaOmvtUuBM0wWbcmrTIi47xIiP
mJ9QlfzBgy7S+EniR3RK/vcM33DxuQlft4Y5/I/Hrvvno3Fu0kSTyYZeLdfLU6Uf
/mAPsrD1DCMK3Ov2SwpWeE5as+H/d7HVq7y6zpObrZAFFxTcdsvgM/lZF9Tw2VYe
8/vOLIaJOnJ7MdRrgRvCzVP/RFTYZ4kV+DcHfioWWlna6oeSrzE9ScS0Ze2LvJaS
cKR+3FD57VqOdzq8TbD5pHwgAGCO+QH/Avs4zTmboa0LnsLjRBqdYdemCem9NUia
u5owP1SwK02X+Q9YgmsmkLZelkfKsICAikREeOnY1T8mSoH39Lcv4nxPumxng/68
v+ErnRrrfXPXV/HdxyrSoN/36VfxL9cF8YUdIDsRsU4crwzF6DWKCAfx8D2RsU40
ZE19awh6qbVkZDjc/utmBXmGFdTQyXoiPVwmV18uWxVx+7IaYTh0hpuAlBDFgBDo
f28Mm3zQVZ3lEy3hRCC/z056J+34qivAhUcg+3Or1xXDpVQyf+a+Uh7pL8ONmVot
0kQNnUpUC4ygazz10kq3fSAApQmmpnlcKrIE6dDO7NcMHeLlflJagdXdJURtBHdP
GZB9A0S+hkytRCZgfIsIQr/Dp0F3F+UNdDuhS9k3HI52eq/Agecb2ZB7gBKEE2wu
aPsfvv5Gd9BlmizH4mRua3wBgoKVhb0HbMjfsV4z0AQi1fWxE0XvzKsxLFV6APSN
obNDAgsKjcUbifMdF9s/7R/BFfQLCBVQeJChkO8nlX4zZHqtl6lqn5EdG0r6uTy8
uwDxu4b43wnyAXUkrynU6zh9QS1h+N028Eb7HX576AiIw2IO8xWN3Sz8L2B2LafD
qoD6F2XAMx0TzgfZege60M8oK33vK7qhA05ZOJNPZqZR2ItHdh9j24bGaK2j5Dfk
ufpqBbT7r6ZlPRT/FZD56qDdQfeRSTn+yPSW3tZ5ImCtqYC0kJokwGlpvecRra89
+7awLy7bOe9eDDRj+c7TnPxPYkR/zTBUPZ3dTc2tV3UEDloUe5mRWih+NC+60MtQ
mL1hV3H78dvMUchUudH5L6JEjEZwo9K7Sf899aXyXpySfQd19ibF8fthSRcU0TaA
nL8wLwqcS2pU5+TSo/JQh9NVkrLWmAog4HGdyWUAFXVrvJlljpFCJV9NlIoxf+ER
xM4x/3lnGzBSSQDJzP3Txjy18xX+GJ+6Gh/MNIb3ZMCEqU9pziFGrf8Jrg6v1Bi/
JofNHJZ1xQDhLh1wFIk5eSVzTzot49p5YWyJIheKdaFlKHxxRU3SawhdhSkqK0In
QwfovakBy3eGBwZja8wXXg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
KX08CUVSmcZ2vrgF/P5qbcYgWLcmWU7xwpGEeb4BuXw13RWGur+emPlFydW2gH8n
KdqrtgT2Ya80x5bGJeKcuAhvb5F6HTGUlpAH4e/zUW3ZHXKz7tOW5Nqzgxqip3QS
d89FnheulCRragxmJtFDLHZj50DfZ0Cj0fuKezrcoKnT9WSRfXmpiIkLKk/DPs/8
R/B3/PaXS7WE8DE09FXtBqL+17jPS+eXqzh28ir81I1YNGdlgT+OwtLFWnc+3TCc
NJmCA+9F3ftZwPTK5nspPEb3CezWWMplSOwHTJT7F1nvJWRfbnafTjMoYvoRZLoK
jExNp2gLTN6EUmJBKXFoWA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 27200 )
`pragma protect data_block
+RsVZm0zSwghb6TNayuEBoOYkrKRynr7/wIIk3Q5tqOETpuO7x/7sQ95J2hitVuc
R/2gYj1ed/eRQzkQdHVAOkOdQ0bUfMxsCepvuzxiODE1Bw+AgPSF61bFRx1sMTTY
bITbFCZwuLWNN+bD84S2eJ3BLjXAO0B7nTVa9LDslQQKqZEy7p8JpiMI6tZXOmsw
RGdzjwEIShRTeyt4moTTY5qyT0Qw5rk0AFTO0gCS416QCGYKh7qA9VAt4BN13bcT
OljLuAZpyx6COGnGqjOmMLFlJHW3Kxu7l0zNHDOx5ubewUi48ZiB/Jcg4HNBSZ0f
jCYxQW/bqCPpJ0MEI+BQRV+lNUwxDeZhWIIBbtOx1mXp62UsbjV8YTGCXziP4gto
a8nHtUk5NS1YL0CwJSXPtHYHYFw/ddlpwPi/pMY3kABL2Sq7wp6bmPRkPTV29F59
A6OZ8I7B9TkulK9BDD6rsAg2YZYVYWfogLfuZ1SjRl29C+U5PidS3AVW2+RZBEoQ
dX15JjxMDXGlrEmroaMbw6Vziog6pK+9cczoPBdr3vpi3VBFKY6TbMiXQ2dWjXli
Pds2NijNiR2/9oOlkx67xwEH/nGTTHE9L4CaCg72K8DwGtLjjFHdkv7PjC30kPPz
er9rW4vUQg+P/JOKz58YKlIJc34YdjXHyVUmqV9jrSBXVlIkxsPlOMycggYzL7zI
mTUD9n8FK/ljycR20YI1jNXbBL4vSYqAKsW6et4L/llo42xLDJ+oFgABtxgGOnrg
gLGHwJ1V0rrmwAdnpKIrn2kGQ4naZ1sdqqFnISnFkep67zgXufzz2LMYPcghWUM8
9ZfopgbZKbV02bj5oqgkd8ojQ3NPAIpg5ZF8GOQB6abpshcTo+y77lA9NunDUFxO
bvfl5JjkYpfZ/Onq4yznORYcVd72Bw5Ver5xW7vN8HfXGZTglTdTkx0mIphhSkaP
iUsZ8TIe2Gb7UmB6tPrnsvxAADi7II3K1msKWZyXQk9KLELc0xQtvTI/brQP+PCN
kBVGj9bg9yS+EPUFdccDBCiD99z13osVUEixFZBw4JivyI6vZuRXE+2jbHfR+Z6S
JAq9LZOvVqQiJov9dfA8qXMSpA1YW6L5Zeq6Ueq/NSnJ4MX0RihIq103t+5UQU+s
RUIq+gxhtcFccersvRRRF4/KGqP1l9Ex3+fYNfw0DJSKqxo16lofe3tYWrWbux3N
GCco3hpFLT8HrQnnKkZgSVml3BZHw/xhknP50larQID2GS8xoX0IjUaqs7E3QnNA
vb4kXzEi5cB4+maGwuDMVgSGRG2w46zgQndsYGc3BYu4x9d5P9/Ysz90UnjMT8QE
wyqXTalcEBDDmfF4JvxE+Hz0K28nNuk5v4WpY/n/NdCPQUSLjc8vsSAo8eIrWCog
JDkjlCBpBrEmPa54U5+tmJEoj86T6/XyrCsjY/NqZepKK2EvUvWLKi2FKDN5uO2e
oQGUX0TNGROJ7GxR2kORSLLZC3/uQZhkXigxwb4i7nN/NFRmCCcADQBbd9IflUYE
u6JhXLeBR9aqNddVb9uBvDZAVaCQC4aRvHVLXYGs2jzoSm28j2R2pPJHnj5eyYs5
4IKV81vptpOzA9OSA/VGEQ+B4K7E0KtdlUOSXto9kadctYGLCwqnd89awfkmsJUM
cjPQZcz1+Iv5OT7qxIFXCnE2swyurfyre5awcYDseW+Tt6xEfWksmRlp9ZQpAMdB
VzQY3Bgm9tSl2GrGcaD/tAf5czhsBIbj9rN1K4SSXccNkV1aRTh8CJeh6ObjGXT+
5mMcOH2QalhJO+uEHtjgRklMgOdt0QPTll9+dpgpl9O3CMVmDfQlBKT6kjrZ/Orl
cNJCkOLNSVyibFwhZY2VxOu6QVePht7K4CetTJJizVhKhkmHq7vIdpl4xc3KE67j
u0tyI4o6WE6g9X4P9SJupymKEPHrNw5+lduuTGVmra2fT+47nHfftB8FOshwjjPO
O6v1fg41CsO5q2tEZeHKJfg8WotvDWZOUxikHncfzZ1svoR1csjLi63gkaNZKVdn
CoiZPVDi50G3Kxs8oql7BBcT3Yt2XRkRjFaY2SIJ8A9oTmkhtSmx+UZ71SnF8EaB
jFRT1KS+DkMQzUXmjqA+/b3gOm6dzMyknnsahS2iKEUTkUdnp7g8LsJWWke1iPqm
gjhbhobxsNwDVD1qkLTvlSlKtKDEXKgSmMlzvc63SiaypDa2nFs7Ik8AguIuNOAn
hPJQsBIFDEZkFXOeZsyuCJ+QbClusLQCiVQWfFUK9VdJFLcUxoLdHBg/APoiGnhe
5IxKNDUUS4ik7TNzipt7pgyNraqy6tEa6H0Ri0dGehTbrMkp/N3MKisMpKD5I6+o
XwQhvegfKorM/F3SjqHPSSseC/3MuhIXQzOnSGK7eWSUZW6BE8Cxg19MRHcNDZVi
M0XylFCEBq+cwGNchWc2jP6UUqMmhCsan/JmoI9rkG45Aebke3+V7S1O/kf9/xhT
u0ZveAtvCqGzs0CuLKc/hW423GZ4UcAmfCU1iSm/K4pElkWIvSHB/ydxC/E1rrwd
pCunuLt6QXhjwraB7tyvgEi/OaJziVPN5oeax+8lwPpuiCv3mwOhFlNgx4Eo312J
/Fdr2888iaNO46kA7D64RO8KEmirGSJfUXaadK55Cnf47/5twJfJCVwvuC8qa0zP
aZRIgUaN/ZrkSDJ2/7IV6UpAfyM9xFgo9O0onnNs5x8ojn2fkIm4RLlFtd7kKqKe
uZvHw3oqnDXewbOAVxtc+qAs3wMigNyGkLyLkgtfodY5Oi1lIxzg4lU+Rp2Xkw6E
Ht4PlI+iLZTiYG4WF8/DVJo44hFNd7dixegHBx+HYSnRM+S0fDi3oiuW6l/93Luj
PTjMzhwUq/y7MxkPQMMnVMhgxHKFw+Fm+c2pb2cInrNTClb6VGeMShunossYMSsb
Bdhb6e54YeUhUi+tECWcnZsmvJpyQUb1MDin6JwsYmoo4GxQHBrFz0AznYdefMMN
xduAmTYy/dxI2tlDql7lF+/YM+oy7+lOQqApx+Q+bNmNTpY/dLW0GBc4MCHZOtnh
9v3ZN5569yEGj+wEUbSmti9YcYnfFjlaCUbXxYS/OfbYUAYZdl4e4XDtCbPYvHny
bPN9E4gQFAIms78nl9TI0MMxKnTvYqLrvqdctA0Yh7vBjxDn5zO8+goFfCEq+1vr
06SQcpRKIRiINuRdEOxuWbFic9cq1a09XDDXjGf95mIPeDDJ0j86ggxnw6eXYwkm
Xw9scEf4GLmAX3kdgWif6uaM4jGx/PbJIuhzeqI9T8SepvzXlIaEe+2LPLN+K2E2
m5H1ZHKCJHydmbJG7xqWFgLTIDFEWj1qqgxHerZybNCG85oiODOU/tOXFlOhk26b
J1Z7IBkUGW8ydGsgtr4sc3c3fmTgM52ueXYNjTszywzR8/53UeBgnDAp87G1PQci
jHUWdFaVrjwRuAgBk4mcYVL/m+3jQjACHJibz1qGILRwMZvf3KPXRktrrvKEokOu
qOdXkvnZjbElJikzrTW7Fn/bpqJHP7T13pRQy4WKBjYzQtiCdLuB+94ikKcRiWs3
Nn4Stg/kBycrw9Ipoo+GNxSqp8wadXO396M8ZteqkP/nS5dV2Y6I0zNFis1aLKp6
tE10ibNANNaHMEOpgy6Guudm0rO//4Ss1pfHTaMje3ze22+3LD/9dnfDAD3u0IMe
Q+DqUppgmkF8hnVJhjcLx3oIYfdBoPPr2EQIo/z4yw7/GMKxy66p/vNh4nl146Ij
IXOj9dZz28xpMVPETaKcE0yqmUi/jQzldMV6+XrfwGGV8ZQkFi8WpaURNEdSjIUh
sngmdXiMtUQ1zsBusxYpZISpxnt12oNiFlC+zEwP2OUJfn+OXbyia1+VIs01NIhj
nnjnG/BA4sMvPB8Zlhm0rePRbKHtlSM+uEsZ6qyPlgoEDQ8a74JpP2hsbVFQAsuM
iU1ynSmW5qJfcV4s8BeFvV6ZRTi8MQQ4sSwE68j/tGvzx7EmPKM84bzm/O382GrD
4SO//GKEe8vIL6PgQSQ3lQCivX7mYo+CFRlxoyVnwKkz4V2MKOwOYKWnjhSWcPWf
D/go4nJ78MbNAKkZ6zIsX6dDgCQ2XBVIxjemPJ9BlJYXppuCHo6UNVj4wyuCVGy7
AFvVk2sloD1g+E1LcCBUbgB6jS4YzW/r448uLgYznSIDVxp7/WhLIBtezmaVnyQS
zsqKMdIY3AqyFRcYuYyQ2WNNKy9l4Ck0orjR3ZzVX/EC0tSYAlfFNptR7dGbHmW3
FowrVjU1x6StMO1+/+8u7kbdC07nsjBeiijYG9cYlDIeQtOSPZSEqIJBTlhtKaYa
h+V/0X6A2DJBNXlXKQHnxL7gpsmObZZF0gU8tLFaDcxgwsBDgYPYTg4yYNPbpljC
Cbgk4HQVhTJ1wuTmG3yQRhZKmD9/7YMNf4niubS3LSi5S/kj91zIDZHYY0Rcz4gE
O5io4M9GwWCvi32IPvI/0kFgo1HNdTHQU90jFJUy3l6XVdkXUU94ulsy7+jXjp00
EC4gi6Arhn0y3Pcc20AgRMN1xscZyDRFU1KS1KuFvfhBNXnl9IaxCkMphq0iCXkp
Cm8tO0ml83S1g0ECCVEBgJQFBbnR7e7sVatXC3kcoAPZXKHYyhHOGTPvPxEC5BNX
BKY9lpRoo6/LxZpmkGNM1M4xY/Ozeng6YXJA5KfvfU5Zo6RyuBbPgKvehRMa2yfZ
od6FFrT61w+WU4JM+4XJ7+Nr+HC/nzOaEc0pKjNAnHGBtvALrGmtlaLkppr0EwIB
RtwbZHa9eBYTk20fHj9l+XAXavSnr/Q6eMCDIkSgusrx8nzH2ie1DlF1aHjWmZ7t
JASWu2dAa67g6CekSCd1TT0ybPK6nC+NQK+1EGtfEJ0ZBX7AN5TVlmcgPY1aGOye
pAl9gEa23/KfGRn6LQMCwuFeMICmHqLotm2h1cQloJnRxsV36rGU+BHew6T97p0S
Zz21KboVKuEwWF8TApXZQ+tDqrLx1ndU1NJbwC68mLb9JW0JaUw1sQZ0BGLf8iW1
w8DVpJq1VlKp3+MHdcs6wrgp22Ddo5iRbgAjusENdaSgYsWKKaIp6i6T3ScDbJ8D
zaWPibYf8PZPyvTEWtUfHFvI7/RX1gCfeEJX4K4NoEKO9a5nfqZt1FuvcdnX6NW3
/nqKkzoD2vv8efn+O9wxKW5VBue42Qn30+3WOHDQnyvV1LOApihAytub0vQWqxjx
emZC8TCDFm7CEugSK+C/guRsgf9lNrhgRFQsrzeNK/s4Eb4691o+e7fqEd/tOnJ/
9MKxIIByJqBkf/frr5zFGAaadaoUGuhfkdqcJzrNqm2o2KlAb+6X8wwOrclVc7J3
OluIK27n8YGAh9vZG959XgzXgIFTtR3P2GP/Pg/mu8P00Bm9yXohyBAZAiUGo+SK
tf+FCzdSvkAv/ZMMfuiZR+vdGaZcq9CzCcXttWSXx8oA8vOXwHWSUGEagloOSpA6
cKOB55PeWQKnW92krbu4Dq7owicy4FUpx27xEPaUlhtejs4FrhMIDy5spfSDQT3T
WtkI1hH/ZhtbDy0TgDiATmVLRXc9oZxScb11a0MocKPz+dY8rOAj5PV+dKbboYTh
f/yS5gM6ymFRDvcfJqufcYrDCKKaw+Pwzt4LwN0ZBOy5viNeuD5UiCQ5hnVQ1LZ4
Fil9OBwDxYA/4xntKw5yOzjvOg3ua6S71m0tJw5VFhyFYCD8lNYZMNU1VHTJmjLH
Gcoj96QUs2QfTpLjgNtE2vos9YXVFqWc+sJ2NnV3JQHW0GbrfaypOb16henGcVvY
fHPc7CR+P1TgPTyijmJ0hHw1nd4BNDAdvDnkSkTrAv7LxAUa81FtW0DPLhJBccS5
w8k/n2v6w6gt22MnaQTxH2b1VoZecu3dtzRy7nRGmszQMpd1ZktcIvNXJbns+PDQ
1G258Aw/1ZYv4/UIXNdoSP9aXft7hfzvB2D7FWU1T6cm6V+gpxvecM0Sp5si4w53
kRPdorL3BPYN1EJlZDwxIy6e/djKQ3mCC29jQaQv9CPZ/ylLYh03Jrp4cBkctmpQ
JRT8UzBPTiCS37aKMFUibb4+Pfkko52jm5eljkN3rZjWtVMrZgKQIJWuEMhyVZlL
2rzwwEXSt+rUEceNhkqQEkTJPgNdecx6FYT9kPXZYygaZ8KGobgprhXifeRC3y//
Ku7LnX7WI1Q5v0a7Olx4uneMPRqmHzdnWgbIcbCtTF6TN+WpDlO0qjYzOtlAGMf2
w0owC/NhU7CkUQBcwB9M5CqKbAO6Aj5ytSV2N6Wr5l/8sTWKCpnZuP+LO4m2YTJm
QXiirH5/WYsQvJ8piXa7/ABIgbEhStNqJ0Vp421ArA9IvwQiNfiU8AcjkvWVD9eo
lAqNKa6mXMq/HyFbpxv/0nfcm8NhAg6VQDmO9uLRa0ftnUUqpRc1EQl168fbAy1m
h98N0fFJ/9wikc1aYnCBzHzvUtiG/Eeb/sAdyk69luVuHo5bWxNMgsV0kJdiew1a
pG8NppenLcSEckfmRcuqOSzZzLr4q9vbXNh5xkxakF3x/4D8NQNSihnVBkpqvWEw
Tvop92h49s40wh/lJsKJ8MiLI2p2yAb3UqVBzRLByXNuqEp8AGnO5iKtRIrgDVVk
RJNQb1Qc62XIJ1/I1jDfBel8wLESlZxt2LbuQV+4yOjiA5f6MXtzWbqShPjt26Jb
xU1ORKkhdP0GAlgYHHZvr+W/KcId6n1yHuKPE0wcdmz8dWI8aJBnbhZhYKElJYrA
OaCh4rkBoJle50WPdvyjXAbzxNj/z1dlL7Goy+0NX6ld9HB56qg6JQQkF7021VPn
NNkeYjPJQEOiXckUytwG6EM+fmYPrNfbDHSmAQJbAG4BaTcfd6Bnhx/ZhJ73NmB0
/Vz47va0s26qScaQf/jqWAnETFBJs/omAliydP8stjg4buPKgFJOeY6xEt3c5jBm
y0OaeaiG50FLLzbfG7KpdaKd+bdXYMzm1Ica2VDuS15oztVgxMerbtkQrtoRXboT
rLNNacjGLYw0EIwD6KJdvafymG4DHTWkpJl+QZ1Yv5wx8E2wkbcio+Sbrsb7mSc6
cCUCPCBU1rq+92PMCSyoqU2VfUeO59jj0iLYD99ujp4r8xb1rvAztVtvfgyO6XtJ
kIBqZfp+o1nJzyzpljOtJUtqjGuR52qpy+lx/ZRuASs2cyXPtCFjcSE4vnpHkIOZ
E4F/mYXOwKw1w0072Zr/7GK938Acb73w5ZAJclnOpwUuJ2Frz0LhNzimx1pOO7+m
g62NGi9jxaK5PcNp31cvgx0qculZp5baY75EXObMUR6lZp6ImE5egiHTD8VjwWmv
p970LiambniFHQFVwmExeRUHJRD5KT3tzeuvTVQroXQcEuOGjVE6NWdjJzIzEXFi
G8CFJs/vmKNRUVolduS2L78l+S/IH6pbCfC0Phgw5p+9wnEPk1Sybt23pkMICibq
NRmK/8zvahwi9WxfkuSPvclfmAasoP5hSHgXu/oMWxO1irl3QxSl0pHwwOw80J2s
FQGdMyrC/+0XHpTdgQRyrORq2M2lxi4CwGL86C+DyNGsiXYl/abcDoj4H3/BUQr9
b0tmfWvv8P7LzTJKzkCVWYWydYd6CduUMevp9ZlUDlxtxAg/6t7PYXwYNGeyATRq
2BBIEuAX4OjtWqJAo+ae/NnXDXg8c3JxkjDtpNzfORwpziBBdXykE0hO4cdYpDKE
5qDBqAK3ZbubTWT/Ekdy2tavICaGMjWoTkYtjFzRjzSBvj3neTTOw0EEHrRIEfNv
fwQWAemeWI5hdQN+Ycs6NsmlEYxi9fqK9vWmy+CSxksIF2xrHCxDWiojRRCZdyT6
7y9EdY2vcDZcjhDPVZ6vs/V72bpS061EapBAFoVeaIh1R2+/JaYpJI2ETC+jbgpL
BY7F3A4r5/pO/YtUa5DpLUzHHO9N5L25I95p1CKLpyJtzGwUsiXH5vCwuJCGsUnL
A9CDMSazaERd+b+tJj9W0J2xVgo8s5OA9WwBJDPjnHPAn/Xb+mYe1c7lmNbyphQi
9lRghgsS9UX3eNQe9wqey1khCG3Lq7zRFQVS7HqmZ8PqCK+d0X6FBCDB1YswH+9/
kUQBqJY8xv+Ph3RLKl6/ZG3+tILUWtxmAqlq7oHHm+7nBG4qHR2Pa4qCeE7RiA5i
27Ya54KiNSf1fYHwADKG3+UNSPHGyqtw0vEHS6sBY+e9TBcJkVOJVedsNh0CY471
vHcPdMBamJBAwexAkd2ZG2qEiuK5rsJkm/gROaJ3vAH76Iu81L/Ns6+svIocJ0In
fzHyaaY8LuJk7VmHT+EdSVLNEkZ9mE1JcEa7JVK4gWLGZOanBqEju89lJzz1J7Fq
ayEGQuBKNSS1ScDhi0N4zLmFzDx782ZFp2vM2I3c3L8G51bPQNOBQdt3ZPXjXWpK
z2AvxDsKnTSiNgGqKDnH6ISO55zLn0p3FwsGYt0QApomIzK/2aj8qxT72MQsObG/
f3It5HOLb3EQfF6eAT5VkFbTgswkLmjRYgVL2BlPU9sngpRw3cE5Rlnbkwccy+dy
V3nyYVu2/01O8Ywd7xNLkwRVrZeL1B6fQIiZPCs/ddgHuNewZmDbUxsUsfbTqkmU
FOqDS7P68l0c968+SjGU2Wn6qgHWYGreJ2jjmkekq5b9NFbZX2bUIoop+tMWFKw0
la21cosJjitt0cgp5ltCd/EVkaZT3JlhZEBfNnZyxtBsyvEkS2OF7Ks6evg3kVy1
TzyM5Uxx8b4NIQ/ZQFzpBq8C+oU3HSV0bBrjnQnfvrksTN3OiVzhjkb7lblnvgZ+
B3ir6EWm8d1MnVKomA9PKJaZSl9Ws+riggwXNMrw28EXHtlBxizzxQedOWwDssQ6
NzSY06Ua7eGuVsp0OFyybUS3B4tYQjoSOBUPn/HCsLNvyKhoFNav8vRJsG3kfH3B
PPvHL30aJmX9/rxrGoV0WeW/vQD8taQKrPAZ8rOQd7ITXGP8W2nNoP4DO8QvfbgY
kxDfpADCL0pAd2tXu0WW7EVSIuBrukrrNyNQ3OhuHEj8Lu2P8s6l2dpuuxff7YZp
ejMxnqklhUcb3I98YCt+78w1NdBFJIpqLVhxEYAZMXmtADjgZbfF2p7FAQsp6q5M
kLvfH0oiqGPd2pjuhg7aJY6VSZWBf/KFIsMQ8Tt6kTPNdE9AqBV0LYf6OsEypC4l
DJGDaNaDkuS+8dO16wQG7T/mSmRKyquJwN4TTj8HjQQEblCs89Gjic+IkJi3xxqX
4SgKYjuKrYT3OmTTwCR96H9lTYxQ8zofwr01nMwNy8bl7xH/mCZtr0B8o2aBUcSz
McIQpmpQM1iY55nCFNdFoVxPGFIBu8Cli1Lfl8EUqjc/Fp9NMbz3K5ZBdT5bwD0j
AWrFZEMfDiYNO79mXD3ppOUXdTqzGZQnnhA7tiapbmnuKsikBC8YTPP4yyBII+qm
oyiqKdnLOVhbZWoEAbuGTeAxKoeY/6ZJj00HPnlImA1QWctlLwWaWGqRxI7HaDzW
PMNUbqH6yUap2rBeaAm6zvk8bP13GpmKf39sz+mO9hvyPLyI3zzKtonp4mWdDOQF
F/b+I9CsxqI4TOKndMWVQZ0wX5rLzrb19xObSSAatuBcxvVpCxXhy3jOLFFu/Ybu
3OQqEeaD3vnxKYqlbWQ5pfKpTEAX6hwbSp11Qlr40X0Jo9f/TLAVUBwYSiz/DWaR
CXT5fMtppvWYMi/ciZbooZp9DPteik3cZdeSZLO5KcY8SHfWsEwcHMKC6FtCfnHG
r54TQ3phom56iGwEX0ybd2FKlLhug9x6ZVb93U4fDzdlni0TJUEbLzvEwxDZUuaf
x6XL2abdzK+BlVEiJQMeUzsEidyt8W10vhVdGNUC/x1gML2EL/z+DXf64N9sXP04
rS2Vl759DR3au5WdWw36XI2588akUpywctWp5RJOaCmDcnBBpBPRv958ketYjQri
/3biKOsv5+iZhaGJ6MmmQf9vUT8OGqomgUn/4JaJSa2n+6o8b5uFtlHXi3Px07+B
2jUoSyqItdSRQOppWbsaVWF4M1y+OEJhPYAzF0/LIOVoQTMKdVVeKZnlJ6t6hopx
I7v5e/WoqQg7RY1AdFLMvgnW8ozF6L6/Ty3v07erPjKnIqUOf+W9KdmnwrjnybvK
iUha9UdBRivg+l+QjrMH3S/qQ8JoTov7Xx24IOaHsIyLH2VKY+bui8fn9WANH/50
PGvg3i3LzvZp5tbDApzm0u6TyTCJqi9LLRAd5ZUnymAs5Nt4iuS7JhTmy6GHwXW7
prDJ4G1IcEpjKTVwhX2X/DMMAZedutd4M5N4/CWQOlmS7YvpDIirKEbxdLo+yNfc
jH8FCDAkGWWMbkAV49ZIHK6IoTvE1qYqDpAEsu1y8ZTrlyAgkH/g1PQzXeHQBfRg
ErKoj8dSmPIKZbymOkZ+7LpkVCxoCOtMya4gXyIfOaZypn15busf2xMm44GlizUG
Dd2G3/7BOOASsJkmnw3Jp0eZn526SjfSUlTmhclyI0BTYk0q9fdcAVzbERUsyFpt
obTFoPESjNbgqDKLnE3rjpjkyhKc9+mraORwAMPhHdL11ZrW6I31pKB+gXntcpGR
6eUMgEIxhurBqlWFpeGrkJx5b5rlIFyly7QblS4nNOTaqDA7sRcsBd8yjn1hftQB
jszMANaMLD0Wz7jyScjLM+GIuKjhNqm3cVkkUziTcV15c0DLEWjQnquZ3DbveLxa
hO2Mp04ug8Z+4FJvm6lvoowOcUriktbFng9Sd+X7zl/J34txwsjyQgpN/P/fWGp5
bZ9I6V28/OQDPyj443ies5mbnoqpLCC9z0NzXZd2h5yfWum0l4zL6zxBt/L2nscl
vwWvgUFNDJTm8Z+Qvf7tkL3F6jPdWhZ1VWSnFR4ItoNae1X85nr11Iz5hANbtk3U
9oNAp9k4AGdbU/fHeKl/KHYv0Fo5ePENO1z9fwBZy/s0glK3p8pSUaFJu6WfYNjF
TM8k0jO3mV14IxAlDDYdRpgprSVQojvEgS86SRNwKBzpvlKTN0uPYGnhygYvvq7f
V5CkM0PwuoiABi27RUS/19hsLhv33XrZ0oa26ai4o29eMTvsnrYYB/QEy9VZmaZ8
gM/3AY3MY8dunhWHtWyoWvzuYYC9n6fHBPcZG9t/1FqMjhAbtP97uY8KhJTE7Fgt
Q/pIJIp/ukHZ3LombGRvMtTryfWT6yC7xZHvsSNXsrks3mj3AIg377o8XuAt5kii
it7tSzkJ441TqvtYNrmgjX6sLJwXsTCxYgylFetgYc4fnuYVwPfp6om7FfXtIXE6
3VIh8acm8ng7lA/HGmuJ3pDykNxolemvukdsjIITYgtTVUCIZpGDQgmswKJ7SbEe
bV0EdpeLCFf+BIpOALwAE1LBFsvHhd4CEbBen3rpUnmQXmo4T6N88hacs2E2oXOJ
nt3Wre1dCQhsZa4PQJrEGPDtHnPK5NVzwQxEjt8AYvkgexFWJ2WBeIFIKL3dNrwN
Vw4T1jurxAT8McZOZoc5ymGMyt2LJD4hSRr0eTx6jd9ApXuXal/kcMkZUl52yqcD
fJ0xVcSdlSGucUTBkrQZCq3JGN0bC+FSSDffPiUWTksRuRO0NnfeL9+ECXO9t7tp
gMSbmGrs3gNTb9eNq/cL+IjCtM7duQpp0vllEy7sx3RhSGU82j4S+AaIaUHvlbmC
sdSIX9wmFSUIb4vcL7Ul6Iosk3cy3PfFfLBXQ3IElbKyG/LLs8Vj2odaMFwusuRn
rP691dFlMaevhJ4qNrvw+7FvvoPzy+FWUXSag1yAuGy3NN3cFQPoSaYmnt/74XnN
V7NxMahzAnUb9+6KDO2YjwhAnHYsomemD3UZspzzsZl76FuMx8fbxI1TZEO/SA0K
cFC774X4v4f5rEbPa9AAE+OG7MYOTBVaMU+4jYDpgzOgfgZPs4emn9xqfBpGqFdW
VT7XNPNsZgK1tswOR55lYUSNkvMJhwkEvHhGeM7DYdbyZdWtBKASyooRCTBhy+0G
kaPOTm7GSFERah18GUR2uiGjFLeK6B8fJ/mgoMo+CWhi1xn6bQdnzgIT86rodG5r
k++xaQwBGvL/WJWvGCKf5603aggCbfw0z06u+V0aOZPkSIDFoV2pAO83pUaa+3hV
K/84JdhSvcuInKDNwyH8RkEyHs/+Yy/7yuMXEniGiEwI11byiLkgbc0ABp1Oi/pD
bvoLA7lDwSEsNTCXlUf3KKsG9GnRUbKvSB/ybDba2RqCsVWG0VgOl6ijy5xW/CX5
6oVwDiyJogrbReVd83kTQO+ujBBMqKzRnIDHhIAWXb7jFmLrEPY3UokJJDlFfQLL
uW8C61hlaLc7SohhSeXp2Iw18eSe32mlPxuMsjDbnN3H7x+P+tsRIBHjSC5EvjRm
qSBF9UvOqQi2DqRP5O1V5EiD+AFAlwLvmIK7BFAYIxTEOj8xGA1iaDvkEVTuEiuF
NnsAcTWa/gXJAdPU+5pDfrhPtZPSFFvuDy6nLciSAUBQFPcTRiXQvTt8H9/yOXCj
0s0LWsjpncWGLTda6U0CWWrYvJuUlGt28Y5yR7f4O+Vr8YbejtzaFXZo/g9LJTPO
gz9HFncEE4N+GLB3CBdA3wtN2d9wl8JDrAfTejTYfkhaObKPzfgYQr59tISahW3i
cYGs1CjHxg/Z1kCugonHE669fhemmECRjbd4/YoZyMH3Y3Qxm8BZAl/l5ZiCv2iX
6vSVKLDtHIPAUXCLNv2djltVyE9IQ3OQPV7QocYlBx/tnQD58tJiBiDnVH/ZJXlD
VwtztKX79/oUB4TkVennOSc+RhhEaciKdwlKzYKJ6aAyapzfCf5FqJ9GY+RY+EZK
k4Dx8VKywcHfYzQgmzpx1heGoFSIlAFnmwTpvUclwA9317AVGoOmCHtJgJdOV5Kl
D0TjLyU8YwY98E1z0jKISuLMzT5gkifU6PodTPvyaRSmpnEjVpKLIyl94MMlw0ry
ysryc5jtJBg3p/yjVfMt2BHKHkAh52Hb1IwHyS4wBaJZBDF3bQg9GDR4KwImy7AG
qXd8TVhI/mPaTPkbihSeNopxnuFmXhYEpnUxBZGKOajyqahRuBCaIHYRSoOxSasy
C1mlsiKVI/2KT7jmx97xpyuQzSPxaqHSqmcg/euD6fmyaDtIwAWzsvmf6r2nX0g+
b1lAWTw0RtACE/VXyVeSCLukV01cFkE4pnkSlPIxekppzRv8t6Trk/m1iQeW9GhB
K8YSztnKJpYE4zWORMcnb+2mx3kblXT8fEPVBxoCPuntKWZiKAkJ4a9pK15oqbOu
l2Jx3pjVjqT2Q08Vd2l+gnokYcoFrqm7ekLCL96lWgTORgEcSetyhHHZsnIHz5Ao
5Ox5txlAi+o/JzJlJmRySzMSF3F72Cwvl0esustZW34NS7R4JgaddrLEswP9IzHI
LnMZIoayuYwfPwArKkdbaLPLkYFGlsG4t9d/A9mru+bAgwusn1nK5UydbDsx1qKl
Puz72dEdUDClxAtoSk+jQxqwiEejsrIMLH5DlUTBgNZe0g6rFlC2IDOd0t4DvYUy
jBIJIzSPOArT33a8DIpz3TS+RNE/P4AO32prz4CMiqKISWGGGtm64XuT3kbePRbx
Ua9Ik849WRtjCKJfSAI71oTxf9jyDWwkilBBqptjj39oUJSyMX73xgCfBDLDgXmM
hNK0kmDqxONc73FBviq5GUd7vtwnjeTXIDthnKB0hwEbongep9Zo+HpzzMOnY4Xx
uz4upuh6C7mIZDrd8nCsknqte65Ikx/mqpOZoGd9JmNAc2pe7wxMTRpHv8wUjZyS
PXhxLmUInDavtbYLmpLj41HFUkzevgx8jred51iBJeZ4mSNSqBkAvZKoIs0wQ79X
PlPKhWFfNVpmKPy1PAwzXNJ/YgxgSx2zI+mDm6DzGbEg+3WGMSDsJ2ZX2LLPuIm1
X2EptReP8drZJ7L45fw9v3eeKsN1vEOTlOi/hI5xE+UEsG4d9qKCt92yz3glUnFX
lhMk6wzxn9wnlOC2Jy4Z1c//+4zAwz8rR412AfQJytDPzytEGpGdRg54se16plW7
/fS575eVEdvOEiDa4riXpUMzoTAFsZWTXet8DGAh+jeLLtNDXrlKBmJjoC5nz4jZ
954k6+SCnaJp7i+ZNKAGO1ovNglQxJ5j7bGFr9/+O+zh8Rdg2czG61T+jzIQTBbn
3CwnVRda4LzteiOyjFAdX05Jb0OXndRf0eovyfR1t+EgrAoxT4NPiTmHl5ANo6yy
u7kR+yeZgNgJSab3TOPWsKIydWMIEuF1/PaRDDdJemcJ1e85fGMtW0RX9Fr1+J6z
0CdvOnOrDQ9qP4qts0SdpiOKG8iqNWiAFsopYOsG8jc3sG2BPrHDy46anhpzRjIo
6eSZr4bT+4NPGP5xNXBbKvNRc+wJnfJ65tRK4F2IhXEp6ZZVRoEyO2gegvLTJTZd
f5WGFRFh50IrU37GyftqDsBrSJxjjCJ3mLi4Fr4M5t7rA8YTYV7fRMaOgj5MGoJU
dJZE/SCNvBeiWOZOAHxVUiuTGwmPZrbJVp6Mju5c1GtXf/5D5eUjNBRcwyMyZL9J
g9dHBAZyhTmvZyb/StoA/MtC3dxlL2mdzF9r/44db5YbyJU7Vu3pvelHWAPMJi3K
GcrrDIDNqAgAEEqsMwOJKsLgjSTxGWJQcjmcqQcczYvGgiQ7nalXi01FGuTQ0ByP
Q+vXkjy/dXjX+YACqqaEeTuL0dyx8vKij3vmGQI9muHp0b8rBvMD/jzoOqwWupPX
CSf+xNV3a/T9hF5HZBj+rfPSjCg7Rklm/v+XCFU+9XVg5I3vIpYbNZzVy5tKMmiZ
aEVpE6kc+nm89gqj+QeKEzYTfOuF/1w/afiGHf7ehhrVmj87Dx4bO2+rNI4y+GGa
z49TWAgIY64vEJiDrKj/rymIPwZmQVn2jWxakOxIfvSGDdTi3UdmBw/5vB+Ym/Y4
AQSNIyZOrzKYdwBwrGb53VjhEYWPDpZ5vN5X+rb86SVP60u0t4e5hqrAilYuH0NA
hdM5Z9va0qMbIVlYCMBo3eU9X8GmauRAOwOKmL0CHPtrxvIEufb6dP3TlB8ZlRFF
NMatXMaOHdqTzkOlCEL34PlXZpdyB8qQc0f0an1rg9eEcYt0p2uRNMCJE4k/DV0k
DO588s1Kr7ZAESlwnSi7c7BCKfX8fw/Qe9XbRHZ9ARHkTR7g2qhhBrShbz0I2qM+
HGZ+stIgsd1bib63VECC35DX2tok9JgBKkLyR2i70HoRaiXqA11hy0TPHZphFh8m
BSVdCzafShRNvHR3U8zX9ovHGXblW0xUAzzww5fBx9qSK1p44LesMKnnbXpkOpQb
dP+bRNXvwItU8NuT/cHLFGTRU03+3+vPGWDqlECMac5lFpkeOwnzzVUiT3udU6kR
txs583gOh1genJyZhtMPmLDEV3q7Z2S+dDflXKYOSNoU1rMyeG+W20IIDtUEAGg4
OoPSR/y3RXXCBwfiDGky8Olj9g/ick0SDcWVC0VoDJ+sGWyH16PcrU+BtEXoMhQv
z32cZ1LbzR6vqpUBBav8l1QeFQHGxuCllTjyP9+eR7u95737gSdDg3JNwcaFVI4w
0Ny1NN4NWc1enauBqjnSnoANetlb4AidaldcNYssJOg2ELLCYrclsCBCNAOCqO4+
hwzftOkkkP2RF30D+CWyMvYAkRN5/CoIaZc7WNzYJNRnla0V2xqimJAydctGokRr
nyc9pwuG/GGBf5ODR7glLLHSyoB/oCEFEkAkiy2zZemnUj3UFaNC+IwVvzDOwHGj
RbzSX6t62/DtmpXz16T7m289muUMzDVY2/j5nWJ3PhXBijXEblbDhqRk5AS3E3aO
5bdEyatyX3/nFSa8LQkO55g36yUDnsKWDvY2Gekuk1Ql3vJB2srKPf+BrKli4cMS
l4DcW3YiOcQQJdD42nI6PyLrlJhtIMHTn06h6Y74l9aYoRh3OdwgtigtcCck9kaU
D24xch2d16rB+iLa8rQs8yXokfGWiB4nRok1U32GArSbj4Vo+XEXAhXBc0nkixk6
BiIkZ57JMSZDmqOvh4RrPZg9Oc4RNFqbuaYI0wT6PH6P/IrdKIBRw7l3p9dFlEaO
tXq6IzgoK4Ouvx8PM73zcvwHoe56dGdUhXo9ZF/kk8+q/Qkjj46Vmz8cAETiI5Rn
OXqeX4mfQA/9QOh8BHAnpzmceoiX0rhb/Ep/xldNTmjTuwtMH7edHKrE+Quql/L5
j90ykgWe0f6XWXo5VAwn0LxwBHRvcG9fz4muh2tmhB7Y94ck64UIpt4+ROS1S9II
xCKy/ibUF97D03F1hVIQWMCutjP4CBNWTHYine+3mrVWh2yb2zlcbfc4r20UHKYJ
888u/b2FJtWtmQ6wgi4Pj88WMX0x8rR8S/jjV85ftJMtLgbvtz4tHtjp4WKns3vX
qQzRb/dgQfKUoQg002cccxb/0wKCvHE/unGS+Rj7Fbmy7l9D9clN3yDSdm4YBH1o
q+N62xpx6HytfhCBMJT5STxRPhh+kw5gL5Yf9dGhvT044fqs/QdjKwZ+M/QG0FNq
DZEhdLRs5lXAXwGImmzZGC6aXexaeGFTiP79XJZWNKotS5DlBnpjZLbkN5m0F35L
BvQf6xRL35OfgeZM6A1KALc2JX6a4iSeelCYOqahK79eiw51xt2PHcsuHFZXQBac
miUr2mFJu6iez95YMS+rBV+DSmu1xKO299oMYjRf51O35Ky9JmuJRYXT4bLlWVxo
d8+C+w1LtbGaipjFHRSgF0K9jA/V90sNsH+x9wPV49/xHXg4ZxD38Eoo1xSoyBzd
SU3e3jccSB5N3oa7HhDiByJj9qeE2zsLA1Hi3D3uToJS3nXJLwR8TV0hMRIKBhOp
MdqSpt3EY0E/LsS9HLRdSuhfew598tOxHQDN1hlcLSEYudjnVBEwXGccT1m4PGli
KUAYgPqOC3YlWaQofsCCFpFGdMbHlp68WTW33srb8OT0vcgOBqRkW1YTFxh6LZnM
+d6VnGGS+Vu5zzJg8Qb1XOWgVpU9G+VjwF9OW2tx8GsgyH5ft+xBse7a61Rejg3f
8UIqZHYqak8m7hA9KqHgnssFfaqHSt8sCG5jQb5Dra6eb5L8bjs+bN4mpnMJjzA3
mvEMI59nitzZBNDlm/jgzbfN/8fvZhmbcAMmWL+TDq2Yl/DROgVjNxJHhVWEpuMd
MDTmiaxSSgmvyvoq1UOjEfx5BWID1umULTNJXFFstuLqZwuNk9M21nVpqm9AWHMS
VqmHBWfNpPymu7LXqbEF+8d+GAKx4j8qOtl2+W4P0CNfpxJ7r/L42b5pzv8iLUd4
3XXK7+soUSxrQ3Ugka1RMs8gagUB7L8ErdLieXCrAYZfDvFj+HH3TP7CLnIfb27g
JZMR2oWbWnVpbPSeQ+u55oTINg3/CC95VcdnA8ZwiFaEU68qOiGdJG9BFSqJGPwC
k/NooQU6SRXx4WOpFcEonFq+sqT5z8T+Y7hzqbb5Tjf45Z5W7KOmtOsO75ScC51H
qvjeKtC/9hu3/wDwIY/L7qoL+m3t4Yp1hmrhU+ikDzVCoHpZGiI4tlAVbR+8NmDa
XR7RnQ0ywt6fNNMSLK2AFP6JUoR+y5FvNTHbDa93AlANIfSixeTXG6fAKXxk/CBZ
5ie02xWX8LE/hu4AkndKMkAQLVCbGxY1L9jGYqBKoELbFkZwfqo8soDQtJPoPTFN
4AmuXqpW1UxEdSiLpN/VaE9V2gqi1l7EpxgaBV3MGz7ELJcGqhLbUy/O0D5FzR9i
8V2M+YskOyblHJEsczOn0h+lg1rJ5Yr2dF4Hy9s7dhjz+eRnS2eiouUftjqTNZMV
p+tkLUuHISvjLGwJBjlLG1E/SdoQSyInHOr/QSch2sN+9QY+Ujm6TLPgTbrEI3ib
xAQrR+wedbcU3yUt/SBcypmq4ykZVW04SLG9CGGvRX+hpBkCa+llen75BfZjLRQk
BxpLcxR8JU2la26wDOBauf9wLokYr+J/pLxzEv1PiwsogYU1cc4etb5VKA6+kBYM
QhUuPvQmLwmsm4uwECBZt/hVEID/P1mcze4eG52Z4uK3n8up1H4OCNkvo7acGUle
anP7mZi7uKoKLBZTuFmFVzvo79EjrGiNXgqA8IXvuCT2k3Ds30MKGek9KIKKyEu9
46bLNQJX+VsfaST63DZBX6dH6I5mlOUbrN2lSTHhGH30c941If75LslDU1t3RQQg
sI9rGQ11zGtH+feGAN2FrpbZAcWyJ9MUvhj5pbg9mCebbBPrmFWdtwDyEdpDkIUQ
zbbaZCe1dCZDpAzvNLETfOxs/s69ML52mvg0ud0oH2ZM5xa7QqBwKq5+aih7YP0h
hOG2Fw0MJ9XDx/HlSvH2C1YdbZFDbYkHb6wW975lPwkwLe+Cb1hArZfhQPPL6Glj
8/CFjTP76IO54P5qaguYqBtmEyuB0EZ0bn7l78kxVbsMcNxPl4XgiTMkRnlmv/Po
ajlFxbXsFlT/joLtkKVJG5q3v1EuD5MSjIjytBwYqqzZAjNo983wD/YFy89Ifd0V
vlBtGg2DtuTf+/vXmfTtH4+wBNUhDj+R8yyUQpGfg/E3uQZ8dmYr1J7U+B+FFIya
/TEhFcu3OxKeztc1XevSh1YqPim90WTKxSCu765aUE6S1NBxaBmZQ0pu420HZin7
d6MG1ktrj8ivMPnak5vJtYkZuy+qOUROO/qBQrSXF5BCXYN6Mz1I0Gg9na4aVgEq
rjbfRlFAIMrmV59P7hZ9zTUrLFZ2ya4CtOJZuYybev+vE3OA8fKlQguBK0niU7Wz
7HMdFrlvhX7GffcKowA6RpPGDvu7jIAGGqoPczoQAzzHBfqq2L3r1rpwXYFIhpui
IlRkb232hbuv1s7TRtbRse+s7GJ3+reWQWx+iOSD335kbJ+SExPjyiDwclOwkJrr
1knzroRRlJ5nRU2fSbsYtTzL1yKlQa4kGxjfhMHNQ9WuYdrnOX1q4xDO7yXr8BYH
OXox5JX8mCsjz7uWiHw8zgckmzqWfAhtrtFKALAe4foxNNGdCe80TNJTS82Y/tzU
CTggT/n+fqNuD2cV/1y683/9jo5TgLWQhsQoh17kC/Ehu0xyOQ/Zb4qY5E8uZn3a
zaftVnSrB4miyWieeJ1KlL+rrzI93LJ0P+iyXRqN+60Kr6a7pzlwNbQe0d2c72qw
sxLVh8rH2nIBRYmsLMxLb9v1pAy3euT8AH0h4jegtox8Lqp/FZJpceydDFkyV1M0
lyKIvXD+3RkTlrAylWGeWKMc7NImE1kMxaXQuIFwnpitTsRaD7Q7H2sG3Z7nD4cc
0pa8HI3vf5azjLEf9fgHygAd2OkLkf+q4WGs0LvC7rkt3r6sRNu87Nt28DG/A5zi
2fIC9vgvFT2mnsn+wViDNmwdSX4KeYPRKzBVhJGV8vHjBISFog235Zgz3msAcsVQ
FWcEwXIghwgzCR2QG3H1ppZ618jXPFT0bd15L/GcwviMACUWMspHSrzLHkhwjzl2
5tIVO62vcXPsxI4bxJ78Jkq5xT36UNaUOBJNrNci1yXjE8Krf1sD20kdSjqBycJT
IkYi9vHkYtUOL5gW6gRIKHA4K77r8cjdP3qQ2xiKUoN4eg2L1n0LWgwj653Y5Oy2
gd3lxizFQL2DkoFAl6q9++uWi5Nstzra5ma3+gT/o2ftcGWDvPX0Dke7Ac4FBhZq
Q40hmL14IQLvMixJrBKBU6CnArCOeWvd8rf2kJlhzRHwnLTzx7hZcijP0yYt9otb
aHbhWjrp3xsHi/747ZQHG+xGvKjxfGyLMEahLH8b0OtYIVJtkcAf843j4XhqQ535
eeY/kSWaB0QBZpk2dAh4wAGAiBx1ksRgRax8qt/d6dp+5UfuPrMppNrS4W6JCFTq
m+C210gxkzF80HYRoANrCBphm35Ynb4/dTrW5YICx9Yck2sSxdNskrSekFWUzVZ/
75gA1esC1xrQmseBIIz3aX7DBLMj3egiXmpazas3N3uWQGsuiNi66AJxEMUrTUNw
QM32oXryRCH8SykP+q9qBNr5/EQ/1W7LIsCWCSdbbZpwJj9OPo7glRHq9DY1aU/E
+wYRfomGfA3ZiH0Q1AxxSOgO/GZ+7DMZeAjm94rpCVrhepS0fjocg5SxIGSqiken
B8YSL1bhTKCr+38wyIMWWZGyts7Zr23zsulLT3yywKQDh4tdafSMFe/IizqMOMGG
gGT5iVeSMFWEjTSvknuoptHbfAiqf10nGuyLGsKAgLpCiHCKYzud57qMf3o5jZVY
Ue9LYAnxv9kOF/7kLpcz8rNdrdtAvj2ZYeVyE5GhPuXIivB7tadQ+FPAjayUePTX
cMlp3BQMBgtBvFL9Tfvb0nND74e9rglsrKqZp9T3HziBhx6O3wXNm63mlH2EWeZO
0i5ktdo7vcQbuxTNs+gT+GpW08Qv6Vs/6TilQ8YS+OfiE33ffIzXSjS2l9CXKrVV
2ZIvYZzptw5/PT+F9M9n08DNrsHFSVUrEGm9HLMhHGryI0wRi4doqW4ZGSOQ/yRl
gFUS6ZvkVEFVEh25XgPPHklsPx8xpv32Lj0c3p8tZNOokV4iZhIjB2VSVRQ7/FsG
GJ/bPQGCZnXtMowUlsM3W931OrZSnepgOmq7SqfEdbXGJzNcjVQX7fFLmdwqP6Si
ll1V5/aAtyCc5LnropZlV5D+D/PSl1sJZQlpa6ojeA8kFoDL2Z1aBFflm7yyTiIR
b0B9lZqnMo4EEzgWMNSVOT/LyIabPumZ3EtrUjYYHxueExGBW4Dv3U28QgdDODJ7
E4kGaCQtpde1mtNkn881prQNLKbDAWrj9UfKdl0uYjX35YVYF77y40m8khWaEKwW
Cy3LO7WBL98rRfw6zzpYiQPO7sVTsievBCQMJ9cKA6flkR4tXfcgJfNIlC7X/RyN
hHT+yVgW4ab9fUNy0/yAbNT1Z4FB7IT5H80m8t5p4NVEKHgUWv117jeynAd3SeGP
7Wfd6w7XQboyPO4/R5lfgKP0Ouz/G15lvXGzByLN10d8rJfg8vLn7HshfZMY/PI+
phXSnrw8tE/oYZtsiI+Kf2QeIKLVzp77mMgsbsdZTkjtUXFRvaB2xfAiFdTh3bA0
v4WK/ZQGOGJsKTC8Kbptus/bMAVijXQvk59fdQMh6rvazPUY0E8Zf2r1I+L8IL7X
ANmpfHwf4aIRMSJoRIXCOFm5Y3ZuM9rKTD42GWq7O+i/kUebsHBmqCblBRxxskg2
tQ8PK2VdMKg2BLk9Jok5Q+iPD5/Bv8bek2IrgzoR4CBymAWAe00pDzkLj96WvZom
s4XDRkB+LL1qDJATMZw1UbdN3zHz5lKt97zjvJPGwzmTfEmA/9O4bMGe+9CyECxP
Zks543DpJlLxRUs/szqtwGsZgrZZu0rnA5mjng9EUwPwfLDCMrrybCEfIv5YVaQm
Cy9erj5KQxWxWMCcs/EDDAwsciGnpGkUQflFx576G8kDn0XLr+A+cS5a6Qn8Qv3Y
T41Bqqkw2PJofRs+7W8Lnh2kJi0mQR+G9spDwicmWzj7m4iCZtDmw5mWFYiDMP2y
R164zNO3M+nuTZIn96vXDHJCsqxvGpCvQIOu0HmCes6k8+5w52MaLtlMZc+1iNTB
pFofjNBDrhxYGoAl8UM5a/lAUJZDOcW2hLuzG+89szJomziB6w1U8NDGZ2aHqRH3
rlruD4BqvGvvBKGRdFjdqzVlaCFi6bB+XYAvyGLJjWNnrQQwc7mxsXYhXr/UCPrd
gsrBozBamgbkE3QO0R73yvSc9ZdZPZNXRURA+MkB+eidznVvmshjOofJiv5eFeC4
A1ISNsV8JXF+KzDIoYiuV9a8AScy2adGrlVVN6rwlvCY1fJhwkD1lH9z81Zdj+S2
uKIJvghHMliMi3jHCFYyvdGVhR10ixCbVSZjh32x0dC20nxAEuNIKW6e/FkVw0Hg
ssG/ro7d7A9H2m64RyRzjYs0Xkb/X1b2v2CVAQ1PYXG5OocuDr3eG3UJDtxoo6cL
8nXgLyPN9oTfOjVGbOV1fUHTtfAsysdJR4V0RN0g4j4ek8cbvV4mXAsR1gH4YkiL
21GwRLJcEo6UXumKnSKSlsFsZwX6UDCMUsNrPjnEVheI6hWD6O3Smn4+V5wqL8+t
s4O0kBzn/maUOcW/PUGtJeiUXYTjevshdciuL/gYC6Ozue4b2YGj/1vorvdUej5p
Kd3sNiErZGfM7rvQvlbH5yIExkhLanbTdi5q1SyDY6l1DoQWKQ329qKNzA7l9snx
1zNNgnsBpesgLICH5RWFTXBUM8WpYFHgeZUn77q+sKgMHGpNtjlFNeYEDftt52pq
YHQr1MC68MgAeau3/bjjDKcMQD7dyPZ5O1jKZ9fXQLAlisUzfZ/gTkVtzUMB7C8Y
yCPxnq/3lZWkAQX92lPNSkSzRUpPTstLlC1aMAJFqWAVDThT/19lN1CRtpCCWlTS
fPeU49LxDljwgiSaDjLe2kn7v8zXND6U4gI/TYiJkiA5fPQzn33HGXO+90D3dn7k
j1UaXUSEYLj9GE0myUPNkOdTaj+AlMwWDpbcVQsFoR9y6niFUxJAIimFvH1vi7IQ
TfDI02hNoeJc7AxpE5oooyV5vGTkp/ITKeJR8EuBh9G5oIsSr8t3666B1rh7iUFD
P8fV9hT5PEEuio4uGoM3up9be8z7/KDsicg12EG7jyOUbIutJY3jCBWzCYv+6jmk
FxpiFSHm7Mnf9rPxYxqmBKOYUtUnv9MR+B3KnQdH6F1nHS6HENDgYEbdZs7YMQz6
vaLBSacbc8t1RbccfxLbgbqxxX95kW7QqlToHIq+3y606AYBWeHtWXaqSUqULhTH
+4J7JgmG9OXdoplQp5YfmoC2YHHLA1UtdHbvF2C1lHaKm6wOtFFQIQ76K8LSvEqx
poRMBuLdKpVPIJe3M1BEW3ccUaH08D4o/+B2u8dJRUgjuYSNwPy8xT3OTGDRTtNO
acgDzXd5J6HDoaZk/zNJ24vvJ6M5Ka0alf5xuodF19m2/JxnYZKrwkH5Qzi10fcm
ika1GA3CbU+vXWKJ0hLUGsb3TX/BNCRen8SfM/okILLYO70W7IJTK82PkER7iV9Q
LLNRiT3VM3DpRQ64h0nzarbsiOzs5KbnJbrZcqeXTomSSwybSuxzWw+H99lS4nfl
95IaYwQhcqZMxdketyfUAzxSfw3lggGfdFcItdiy/L9cHy+9joB4CmysDJW6K5A2
kkvPg49fRrJesF1VMWXDBkss1RjCft0JMj1XpqDfgG3a+n6OHkF6XZvSqJStrmSC
FOmYrFHaZH7StMtRg6fhRVpX10y4PdaSuNzmYCyvkJd9rcFT+drBMqu4wzi4NLJ3
d5nGrAwfpkvXrt8RFDbfTU1yCmit8W3qKeftOqHvHNdfBIHbNJ8pt7NO8Bsmt3Zh
/sYGy5aL4y0TlQWZbjm8i7A9Gre5P9K+Dk+0iSQlHuaas1YsZFr9W29G35S8DXEL
w85KwXWDa38fa1vdn3OLzon40hc8fsCiQUuWWRg+Us3eAkWjuLTSJLt6jOjo7+Pb
91uA76+FdxP0kIRsa06ijncYSafR4h0JBLBrhSDWcs55YBPyTTPXiRhy/K7WnFl+
oAuCbIPJ7NfURMNv4YJqXJAjLykV5HcbCnpmqYeT6ZPj1KlgMC5st0an8pNkjd+C
Gm14vpTiqCMekXEul4vwavyr4hiFEwPEjgpgbEBMyt/qZJfDRJzbJuYVdB4qOUHd
OGfvcFFlmjzQmghl+otLGh4s1lJRrkqCnXEtj0x8PKdko6xNXnKKU/zC3Miy2mmg
Uvg1Lmh0JaPEz58nxFd6+4SBThAM/B4ihGSjEJkyWQXj2OkOdGy/p34L0ww3zcXb
sE/fzCiaQ53zb3bV1iRWPWVAhxpdm9byiclYiovwdSDFv77V0h6bMEu/GPQS+vsF
GVcVp2+vOyChnbVp5q2YqbOUkiBuQCAd6/BZIM0xRQ7ai+SToWmcS0lRSRABoVJm
Dy1FSwmZ2zWY7mzYowZX3HgjHT9Tdk6dhYcy+/rM/0LQFGKdIVBBaZTZgRZ7MaMU
R3qMQ5cKz0eOAj1AR81Fn1NEeXBTNjl/iMFUTxIZ6mpXaEqMbmwdLq7zJKQsVTtl
PFax7Ghi61BoY7YQa2pG4JFSJdzcLF7UWiCjkEaLP8GH1/PHcSEObrbHLwqHvj+t
7faiyJrDCKmqiGhtf+TxWnuKNfzXCZ+nKYYgdaW4whJo14jN2glFwoiWzJK9jC9q
B/Ktjm2I7toSvqbaHcMOTqej3ZwGUWsVt0bO04GEBsWYWflavBbmLP7sCBVhKlXQ
YRPCEu7QLaa5pXLhniDGcbx0+Q7gp5aLp4H7PWrvVIvXiLfH/KJkE48RkmAgrA3L
bgMR/GONEo0W8MCnhE5GaQnLB7jbR5vvP6IkSF7QSsCqGsR9x2BfZYHXdVpud/3K
yVbaWYbZ2SyIDeX6kNpZ4ta1CxQ7bAeMVwKzyDhKaLe/U0XOGTVQmjeSHfjMBWbl
MKsJGWF0o14mjvorAxKueFWffMrh88ELd2mGFyOjrx3lTnslrepnK27MPC6bMrjj
XRYpjqLghYmIsN1hcPYs0xVId0jakaFNHGzX7ZYznhDFFc/dWbX7KfLR+8ai3WAn
gP0WC4ns7sYmuh6xMeLpSg6Ep+U9Vp5xvT8i7o2HpilB7ivduPcKKzvxRTZtewl1
ayA21b7HCH0AERcmYxl1NoogvcmGv3C+lfsW7x5mVzSnzLPCL6Vwxx0t1Cw4pNfu
Yqn5DcggmCbjy/GEZY688NU5TGnFLgf4/q2L63HLEWtCvF75Q0izHb9DtGwSp/q3
F0s7FMc//nIoxIjXnZG4hJddgl74BHuO8XMhsU4I9yDSGT2OUDx5itUbOGjUAXl0
0MGOnT7LqI/5ORlDClQ4TbPmLG2ZWI6tcAsGpisMxK/g66KONoo57IDEuP0l865P
oaeI5wjYw9nZpgoeDmccBd6TOCB7fRa9MibMHQq4JEJgQ/I1oaJLix+dc1/fXLsK
DkqIfGor7bMFTJDS88VZJThqmsVG4idpunzCWJDVT6jTc4oyqQWpDURp0WQdOEeQ
TGm5KHhQJD3Z1YlSLcqXMhgxVhFQjVoPZkNV/RxflidnQA5BLO3I9u7BbJ2CeeTo
wcG/Vwn4zC1kJjOPd+reRjff3lmkyk0WXIhfp8Gz5QGu0UQXpiPRn8wEUDFwHmS8
EVU2sMFL7su1NMX9D7Zqfv5eQtuFaJJCBmYLGOGA8KlchvS5cvBYxYgyWcO/feGj
XS5VdCV3GQXja0ylDWqcV6d8C3jg/TRydKKaZveppikRzghOzq/X+Jw2OhjrLWfq
LbCJ72j+K0YrfC2lbrjQo215+BVVfbUpE9Iig5CnzZTaRyDlbFJq0+t927wfFqer
8k0iHly+0tpclhY6YpAsJaFdo7MwtPU0jcYnUtlIUbu1bAVoRXcMwIzLR7mFlA2U
jewB4W/HfjovVUqSVtCLwX3HR/3IRNZFM9e7Sbz5xp+VZNAgiIVZwOey6TM1hXzy
spnI28HAoUTBUB9Jqv3wbtjQwao4CQ/0EnkBodKl0/5ZKjOTnR4ZeCAFpT9SIRdC
DFszpxaTeyAdPqPF7Rp7SIyn2VeVkggA41GER2nLDqFhTWW+5uEPoOP4PmoFpQaI
R/Ypbp2MhKGU0VgV0vopQCzxzufvdrqydGUIrMXOa0K8Jhbzcq8IdSwiNirSikBh
B5Vi9X6+/Ne8RFPOl6NsOcqhiHavwtZDLFgaG2tBnCinLggAMciT8v2uX2/um7IS
UiD9W2SSbi9ww1SOClZIp1HtCzEVWsPvLZnT7Dd0ry+Nn9uje66ButpqW8RPCh5N
LBscsMToF0qEhmIOyH29HTsFiCdyfKqTW7ZlN+cou8am9xJPsH83FYq/lbzs9D8L
bs0tPMQKm3E06wIFtB6sm/g1Ny1niai2kmXQvwtUC+43u5BDoUqeAaAEBHQfq2rf
id/Wy0+troWpKj0LrBfkNY6f3FgG8V/yCgt4f7PAqtv43x0v0rtQp84H1GEsjhEf
DXj8Agz0UJ9v0Y/u0Dbk9iSUHYj+dB7pgXvJV3Jf0pPj1FXV4az8XTb4tu11Yrj3
tJdj4vSas6tNzxEbLfIEgKr9Qiv1FydpR4VX7J/uK9m47JTtq0JS64UC2sK9H8L3
pMvg1yDRO3ifYvvymlY3tbj6f5QOhh5JNeqZ6SN7eEGarDbx8gxwkCf7cm9MhhwA
nGt26N4DUydGj4ZKBrGJNQJfq5mm7atDIRMtSseNqRwuVODOJPtGvMpwbPVF++qZ
vUXXv22lAMEKBAGZc+awXQ+HVez3fyxXFsiqDrLROyUE5AhstQnO0OsWQGOUtfTo
C5AT6zMbKgzCyewwm5YaZ7TIxt1hqXnv5MVy6sfP0PIUk2vzpbi8UV5QJgIUTvOE
d+JjF3QmVyu1oI9yPigmGlNno8aKoFDE+DgrINUDaoE0ZxRxELu7vDtjC0OaWpET
wq2iON9P3ODf2dcKt5rexqwE5vcR09eH2Ti95ggyXc+LDR8q/lT0QN9L/Kt47kgX
qc1914NXIXXR3wJ609AkqWZg2uEWKe/eWNYxTWGv/1XAcScXRdIkSA+9gVPC9b2A
Ir7nJgOH8UagxY2l8UjZtLoRqfMYVMU/NpUuGQ8Yj31Og15aBmJ3uX4FAxPlmsCf
GFH9WN1sIPvlIXq2Ghc4GiGtYM7rRVY8b95ecLXfm4HNp0QAmSTXi0XkbuPVmg8/
6We6AIeoes4fSDWIu/xMOyadW8piz249JFyODocx9jZHnb8cE1Sg53H0e+N5ZdZa
J29zADe0EUT67HjnBZ+OOieUqaGfEU7AiwNzf1Y1n7R+kEAi0xXSipFSYW/L+tgO
fdkTcPWUqKN+FwaHYjVgMw9cP/S9278jGcLDXSyetJyUBr68b14lt/ZhF1QSsIz8
78gneNsP/QzfzpNtSqsb3NBoHyUNMfSV2Dr7F7IAjir1ZTOjQxus3u6PAqcKMCZc
/qtjrET4OZQFH6zD8ovd+hvcotrltgYFl7cm6LHCoTRTwcekpHpWiZo7eHJ9ZRjB
Qe2L493Wf+sX8XeHUyeLchYwW4Qt98qc9PUk+ouHWWp5VLMjrlVG1BdrHZAnDVp8
YUvmqLXa1QqyYcsNFMzOvbLBzILoezkL00WzEAQ6eEAS0qsbIWGrAuTTmYe8JfOB
6lThlQdC8FzNH7Q/QEd4H0jRp3B3wJ689kY65RcW+tOAndWIYslW67jHz2xwn6+3
zmFsoWwMRv2mV6PvK6RuTiy+y5ltgVV2y46prqVdEBlx5J6Q1n4/d1aaQJkOUSZD
SzmqJvKhiH7xmFnoJ4NrZ4WcQChp4qEJ0+fot+9tFlHrrHkkuhGb6ygkLHo7fbgB
ltav/z4U0RS733U3nzDuGHBHrK7MH6kJ2awNqhEowslfYKB3chcyERVZ9/vy/r+t
WN0zYlC0MGBqP8Onv29DHYPfVu3uWQ26mEzh11YlPxSIglQh4Ttzl2yt6yoRbcIZ
vgdKNpuUiaumyaZaX+9rZ0C/nXTKNbi8hve8+HPYxymVsPHIqNpDfTL6mufnZvWi
v06RYhBnO/wTapBytc74/rQ+GO0OdDeNlmtwjDMloktoHJLtbdV7kEdtR/ykMTsm
+c0yaxRTpfcEsfMX3MjBf7Y2GEIfvzfOQz4Ldaj92edSzT+3RyC0EpoF3ESZox34
5AU6DzCUZ+bRtZByqRnmnIUJ4sZXnERtW3+dCt7/JWL57jK+p/CKPyr1p0FZ9AEe
qsMNKPCkcZYolY0ZZjOShpVSdPLogjY+OlzIP247JyoScKXDKsAFtgVYdLLNo/hB
tHnGbCWXwhajJfHI5/tpyhxoNqk9uQjq2QZMiFgP/E09v5f9YEzOyL6EajIClgpJ
SLOLw3dK6WQYAzWp8y3IpomkW9NPrYiyjS6CC+w8tB+DJyyWhLJXXMR5aRsXzU19
g7ahOpc+ClY98dud/XXqZJulmpm7/lL1HUoiISCqb1oSE1d8npF46Hkgon8zaHYw
lumg1VLpb09sct487HuqUMb0252fedWdCRSdJhh5oK7nJsBARKOZmFGI3avYb81o
d32TJgEjaB3sXsAo3xzB1Rkb8wGEbI8B8VGwehF18cb7GbKiny/X/HBjUsAslWvO
16fyAGnSCfEDmyXsZTQqUOImQ0FBlOMnIhJqGMuhR6HWTiytSWQBfm5oGybQFreT
oRreGjHlVj5v3qeC94Sc5SC/ZFZwKY8CT7J5Fw5BJTk9FFQMyk94XZ3qkV7Yphir
T3PgvlSdlA99XAQVxRXlah/jsgs/gt6d3zmUwvXA7akAlc8xTQL6/3h6Jd854KCp
KcQaNQqGi7hH6h5oQYppJVM80jxOu7l5c3HT3y9QwRRtUPTTK4nQnt2bik7v2YNx
vHS02X1Ux5FDnwnZGp1j3qCODKn+qPB0GfnKFunKbV0n1Tyb86gs7Y+QdKfc1r6p
2gQS2D73kH+hZa4PPTVul0BLelqWBLBuAVwLqKjqqlYGRWbaR4z1bjSpoMAYrzUF
2jrF14c0bT3NppZQBc4iqEE40Yq0lA8t/VBtJyBtVtNlsOCoe8DPUTul+P1Qrdpx
GExRLz53ASVtA9UzScwtRRdrxxpdA20QJ31ayyR/L5ladh/QXH/Eqzj4/wUTVCCn
TWSx+pSmmoDUMb7IVbtcYxWqE0jSQFv5D1e1Ob4er5onHiwBw6ajMPhmCwB57YJT
gs5nbNmSyvziYqFwbXtqJ1hD2karF1I6UgL4nzF5bD8QierPHdvWXwqp+bskIE54
I+uTkLQ5iGq5U9lW5ofsbAgpkSCGRzhOuT6t/hIlIzGnhUXPEtM9FLhTtiPSXdoG
eelKLKL1qFlsdX/1UrSRKfmqK7qRSceV2YJQHf8RjwOOGw0jVx8/T8dujHVndrDn
w9lmxC2N4oUUbHU3JBE6gPguJklYfkY9gPYqhaQZqt1HNMjZkanP26xYgCfnm5lr
MOQ6QeAfZfBqnl4CU5wmATHzSQq941TcRfGaajwH3Lo9mmn9c+Hd5+VOdBB7XSw/
ldWF+RNZ2XuUrjLBHfgjz28ettQjdGFO2OCAamLTOpRqqfxRHYVlQs624qECXL0p
r6nmWc8omFNM/4KvcyQjIGEHAbMKh8v1y7BSCMm0c9wGFC9AKj/l/WIAp84IyR4Z
1Cz1BUtymbsdWeIs12cXV51AdAB4EJLH4QD8dZ0brsOpLvcw04co3CBMrv6ThIFF
zruviHtAoi6mARSvnxeBkgVEONFY00n0DqRyg/4QLmqkyPMSud3c7BTG8F4qnKTZ
gbSHWWEotsNCyts/E8PjYCSJmxAKosN9B25USC/fjzMrhkvu357k9fU753UfmHJR
Z8Th1/2ue4b4qA/ORKEinHz4Gc42/XEwMCYH6tT7GmAwcPmF3Uv/NzOHYcuDjIr6
Gdu/HidxLAFXaC+yxRJSGz4/KcYO+uO09lhI6Uns4Oh8FZQRtUI5l5ANNfZJ4+VS
Dxkt0Ng77qJGf+4ji5IeC7Dh7IvQzyPJcnSQsUjCKWXxR0y2BEYnaxYoKzc7rTLQ
+G3Ger4Ao7p6zFhHWWfZyy9J8TRPzura1P9CXbqzOgu9KMAKJ1OvJyM8g7N5kWzh
GI0G57Sv0rMnCQbp++EUys9mYhphkaGV/fhO3lBf4mJkypwC+p1kcDKdalyb6uo+
tyuUl7TDnMPQ8bu7vIwnGFWqYoxT/tE6tkdakMYibsYslI7OpT+iWuWK4C9AX7fB
MhNXKpi/9ef1SutozQV7TXUFaJDWLmE3vUmgr7tbjFhNk4ot4wo2Q3BX5mO6iRaH
l+iz5C8QQ+nynclRAcEJ8JASxz8/gyo7XWtuimIG5HF5vSAHwV2cCsMgiMC0hdnY
/DSixs7lQmwggTn8z93eHIjxrAH2EDWgTRFqCIOdYeckPrP+3k6NCie9N11MHmgG
H9Rvdu+Xg4squJmldDghHgVTW+mBXQ1W+KqmID/nIrwPKZnVdyqzo2CWXVN1wGKU
ofqexKH+AwIOmGkoaski83XhKPRnjDlzkITYXuhn/gtxF84PFjpjL5v9ZfWK1azg
tJbg14/e55KNsMnrE2zL2nenPBs4pTo8nsSqpg/MPhvkd4L5xgWkaUu0mnBZFKbt
KHlb8S91ya3eclqdLVoMpgCS8IIQUrqBxHrbB6gQb0rD4u6saPcBumxitmQ0xJbp
rKPPAyj7NhFjYrA6ksjoY12bz2ifoQRlrNw+R3d/VdfFZ1XAm3rLTKt4C+ew3dgI
2WpEhuD+ALJ6jbn8aAuCFGgy7Zdo83ov55gJA6RBtCqmw50dq4oEacc80KeJFVoH
JAud+XmT63abjJNFNVxovJcaTjgbTmazbCTDgBgKoKG/15yzUJKeGBSkKZ3SQBUA
in/5dev89zTcThqLw1FG/xneOxrfbsUh//mWSFn1LkM+DNO0arxDI7xArVIb3R04
MDmitordG3xwnAWuyZAZKDohNGqFKboiefjj7MVDQyWIiVVTLIvtOW1pRscrqoce
d404tT1OboGZI/FmuN01c0r26ERqqytXIZxg0DVyEusk02qTBuNTOaSBfKuzRpfS
YPyBg+jjQDXGJ0GO17M49BGKQz4ey1XX0aG01M75s2/zTRZ4IaaOgBRh2iBTk5iH
lI8l/ML1XGEM+gC1Ssxk1Qb1egN+EBiOFJd1dsNqx4SUVOgWlwv9flzH0hsu1Wzp
JVeLd3Hv/fILhefN5TUB7ywjxo0N4EpRnandGrNBLeTnzmP0G7URSzI8jnGkwTS2
lzx4xQnGWuO+isZt9DfFi8ydAMPJsx+sOIQaRSZUtSJH33ZNwUomN0eLsFkW+TPO
anR51/9tc5lTgo4+56lc32rGTbvdQifnqzjuumbpVTvyrggK5TgAgp75jm3JouXr
Ykq6BwtF8jj+eAnk+/I5gByli6O0ntxSYoXpCZSkvVqlA0O0kcZsAeXWZ98DaB6y
Uv7TUiStf2zzXTBaaqiNmpOzDR/myz9t5FA1iKqPiEUI5ifBE8sw4v7sVrRWbX+e
PKLDM6aQDvBP2ZrovLJz54LukJN0FXSMXAznSS7N8TZ9XR7Trhf8PbH1/df7sGsM
EIbArgxMiFfVMCS2XXPSh+K+HR3Bx91eLvsQFQZ02QBZZ6AqNHenQSltp7509UZT
OTO0/7fw1zBA1GObIF//5tuepUpsZOs5Ho6fo0r4wNnqrUL8HAuVfwvVss9tGHnU
8SLiDBIxhCp4EuC0E8ItS8dP/Ku1o2RC1woRVQGpYSufn5vcz3naYR7W4q31x7ll
tWAUqppjV1UwvNmo3csdQcij2Yj0ULNht/JJbUgsD1mh4Vjs+3UD1+cGmbaw00VX
jYixckeHKSCaSls3EjaFF7TTvXDRQu2uselu5vVz47/G2S3TQGOAT9fUb+ihZMe6
83TMxzzHNoX5CDYNqdN3cG2pKv4HOYuuNe88kcWEAEe0bOoUfyQUUVzA75juviF6
gX15ZCrkY5PG0XBehoqVJSVg+4CnDfAfcnyD7m/rt2YJP0j4kX6sIXN4wJqE5oJh
lASDtuNOmlSl/Sax7zdNAyo9Sz214bRd8hIhO88cw2Q2iL44XQ7SkWldF/tCdrqR
uA02qxwTlAG4qsrhhJdL4xDjoL0wDZqqlTGrrhoguk26Got4OD+5KOj3dBgCLv8I
g4C4LcoGWbSyZEfUhmHqhxHav4GhBFuoOkRyYvTNo8A8Zsd1XtHLC5i898l7j6/q
roz2mlmBIcOtyDQQ+hK2HVay55ASxMr46NzPllL92ZQVTjLUI/N8H+IyITxhGWlu
HbieBBO2pihuC3tKkuMynhcom+0RHcLzZ4b6yOkDOa1sFHGkrhiM/7wQ7wJy8cNe
KZcQteWTXg4oFiNTRsF7zMHDbFj8qSQhVUycwfkk3w8etmXkcS9xqkvU8VRF3NUv
6AJCqecntrTd6kZz9iuPiRxkgbEJ3YdCGZOiNZci/mYjNdewF/bjWM+vsHwQFD6w
Q57katwn75mZJSB8wK4Yz9vvttKpRw+ETFnKF9bksHQk46ZzRbqBHhaexglLvBlf
NfgrikgMmvVGOCl26lH9qfXufUR/tJ1fmKgCVpI4iQ/xADsfP1lUhDuEJxw7pVjM
9FYdVsOU3mXEgyf3OZ6TuJHsA4Id7SnZZTfxhmWpMfpe8WzCYlr3kb6qj/uJ3soC
2bDR5E0jmoF4ooJA/KY977asSTY+W583b5Hga2cxA61KeolEFD4GgEw3RJKfj0j6
shHWnS3OCOufa34D/YTueeUGRH9Ac7tzIxhwN9DS352b7EJRq19oVFirwWo0/ObA
x/vA9/Uv2pCSqjpXsPpJ5rw1pHwjyumUvhr0p4jDlfpZB6Wqm3MFyodSWnnL0nFN
AVFan2A3ZV0sll4PVGHeyGl87YlJNQyYQA1Lm1NxStd88ufenjNcEvNuWQuMwHky
0PYQEYP5fa+DEJL1g1rfHvyVz7mURYIMpaOJKUY06eWeL7RiR4PEO6sRjK7e5AQt
T6yLn7+khPBMHc6MKwUOAx567l3qBV55E9LIC7XCqFNnw8gnOi3NDFB2aGXrVMZE
npqvVnyLcb/8DhusANXO2ZiPMx16AI+++VgVsBII6WPWyTR9bDAYW+spWrRMZSgB
dBq4mxMrsjyUgslP4KshTC7gHzGwrowTT1lcETnUkG2G/eS32RZOTfyjzCFkD/RM
MTW5vg6rWPYTnAVHrMuJl7gzlgEafwhoUPeEDhDdi226JzfcIqXCpzbK3daTyU4M
TXRpZrpscKzxpafN60rh9k9BY4Eod845tC+crZbtlVAbjnbY9UCe5wKPyF6skLJj
+rbd0D/nsOJnMGLZ5LetvsKaGsIZIc/MzZrcW9GbNXTw/98W4n92FJNDSWh9hTgO
Dd8JrZbv+aZxwWzl2lUoAHKlq9BqX9Z5bPo/E9ywx/+ASL/LrgX0TCyjL0cCqah1
JP0dW93UR/9qmpPp91u291BTwqr6wVls9PJs30NYX3l6pofekPIQYMr2of2+Pg+V
wZcTzQzR2SLDBTeRuTp8wQxKU/fdFBb4C7nwpuf9z9O3HjXAmDOaF4faqCnoR1HO
7bMxlLsOG1kM1Y89bQRalDR7Eoon0eRIo5SZ1hEkr7537hAIQkizYY/3jEJv2Vcu
0rpe3Kgq8KrTPbbK4hmcdS7aw2pNMsCXL1z397fjswFOGvBzrfCs0Puuf6QFCUbo
KZp7baDqesI67Jqjslb/QrlLlNTXYEYLMFkU2J0P1J7KC9JsVawOdUsrEZNi2dGf
dsBnh9A+LnhVR7m5YPAcuczOuxK/QMYla8z+TrloAiYNsjvOTd//5usPc1cHcRtK
atiDCR+OEOFIkkQSkSxZoTXFUhqx1HOG/gCLfB/t1+I4rQqAJNCBfS8NnLtYQv2W
OzguYMFYdYT/JlxQw0aJFLPeVF7dj1wm6LOxHQ6N8ymKgeu+wLulbRrRhQRQD3aR
Of1I6DYbXMvMr1ylwZ7JWSRnBIUdqJuQzqTNjIBD1zgGTcTSTS1Pzx+WRXyUV78i
b6ugu+y//DQ8x21ajwDXtDIW7zXwSfxfaiX5y7NG6ylo2B2E1vf1v8JiWNbyo6WS
rX+SUSW0/b48LBAx3bT/B2yG67vd6DNo7eY2gWy3mA0SWG1fgx2rv/RSU5SuuZwT
ANQKex7oF2Y8qm78sT3u4bMPv5fd/vhAWY0gxBRjuTouBPG7mJ9qJHdeBHFafjLk
OpQ9Jyp5dz8KIZCrwzptUJUOjiBQTcxjziTbBOj8xDa+ohbgDfYSGY7en+CIxdXN
CjU2eDxPBCAKhBjELAuYes6XhQaGKNBc60mF0dth7HAiPERxvD4mkECUdVcCnKUg
Jc8MJLz9KVy3PwmwjN3r2vzIDlBNn7Q8Nz6HDO8mrJhjg/5MgPkmqSPo+PcZ+IWP
gj9aMnxP5FzkVdxzO/gz6rhHpIQ1d9DZQlUYhCBtTGlm2CHOCGcwfB+MmAtFsqd1
k0gMlLls0XCVcx1DhlcxUQ7Vr2jmfIARXPNNc+OL7Tz6UWqpKlzDrR1FO9vV7TLq
ohvjwpT+zjiHIOrVY6yriyd2YoyAd4qamC/Lxnyqu1rGhu2Hv9ldc99ByWtAtjkG
XQAoyCuh9h92TnwRr0fR6RzzUGTQNjzWKzzZtpl2oLuWWbpAMoWuZy6CeAux3ZMm
5AJ2f4Vb9Maspo3tSPp53NMOv4wf49VQi8stY24UXkole0jlduzDBiU64dNTaUeo
fYkt3cFlkqUk/oIplyTgsyPrExN0NXcBi4Bp8CY8Rg2Smti1EyhJNFt/A/aJu3xQ
8Z/UzeIKvvGl8wW7T0PjEGECNpDUDpzORq4zm/q4kEI2seClEMMd3Gf9Xi2Lbr7s
wkCqbDPve7xBMYm2tyFhx2W/H/cP0WwyNjzSCD8GgXVHqJb8bIkEim3ZvRnCZXzI
6Wvnudxo9vATibgsewcrQTuRW5u16PR6iRP8dL+wYsE7W/R5uJJK7+Do5b2sddYr
SqQx7LzGuTpv/o1nkd+y8jMLvVXavYWfaM1PPQkN3v+EtWMxxKjwN5ZsTMQTpICr
IcddexWC/NUopwGt/neHUtLcebP8sA8a3HiNc/xSFHII8NYhzHnM2uL1ZOtuc9Ds
hPjUmBHFRMgChm0evHOFKyKrHoTBu99eKQxz0esjH0Lkwz4j923aq3azV+BzAmEr
vqinZpnY2xoBlS9iLF6HUfAXVL3hxhESVaBX8PAcXfwG/PFgd0p/7W9ehKwXR8yb
1z56ZavFqd1DVomnD2XwO+uyEYN7dGDuAYU87a2eCb4wGLqfgEGx0AkKhbFU1zdN
nr+ZIQgxY7jUD8zVKihlzIMiQAu2Bw+sEwLxGAAez75Xr/YNupI42N6FxyVtHG+l
If7bL0tTm2Q1XqPRIE/zCY7KQFvPDLNdv3fWsJk6Zoet/D9x1l9j7R3ZsnKeofd1
M+Ddc0ewxj1sLQW/+Q/YVeIyM872dtOAqlTYlCLhSiFKR0E+mJeAy0qpxgyJ+BPu
DbpGrTWnnb+scLqMQ5uzqx3cpqwiWixGUwFfFOggWqIUSQp5GfF0hS0VG/JFs30T
QAf94p+vbhLyF25BF2a8LanE1ilY9ruhzZhTw02Htz7lESubsXPg2DYXKLxH/xBa
y2bIRpxcmxKKTK4Mbnh8fmK/X7osw6Kdwjk/GNQo7whzjlWtVAUVj2wwVyKfOvc0
U+o7n+Phz/bNpPix9FxlrcehmECWdVElBbsO6zNAXYubhEch8Flg2dXCHl+Wd40m
9M52roPakClpR5P51mPDJqJtOPH0+UA+aCN1V8EtRzNH1DR8AZOxpB1y1VWf6ZzR
ph3ftUuW6jSPhDZ0PrsVIKH4V2szsVaINpLM3ORmNrzEAk+ywcsB/qy3hcpKbpBb
Kb0xnG4vYiHCuZn8Xxax7rY0KFqHQGh//DcvvRXkSPwc0Jm368r3buZ1tu4MlZix
giIhXWJ/sP2HJ73KfinYgqdWgnvw4KjEb0p0mqe56LB4Wmzg5m72+LJq4PJqia+c
keIh9Ag0x7xqfw6eWg3M4pQ6WC5Ufc7yy0kFssfSgFuH104liFcJ/55cS1HT1oMy
yAyCdjNjOtMA1zPy92meKrKFNov0JMPkv/ceVFjgcH62kKH2FDsLTuw3WiCX0ztq
dD7CwQEbZ3M6Il5GKV6IHYSuk7RoYhYLHV88iQAQrXpCRmyQJDGZcT9VLb1Pu/9Q
DjtNh4NcYG3KA7TolAZ2b7NefhkFdwYmWHJZvC10ovTb216UELkQdz1moeWMO1N9
xL2ywCg40NlMbpOJFaMg0T+a5VRTbVmHxIOfAraWv3AjcVdAbrRW2TQGAiYZq4Fv
+KmGSNYKCx23K9NKZT6kTlY0DDHpIND2Ue54NQmlJ+eVRal7aIu4IxnYVE0JuA1p
/48QWVPXZasQMmNsPs4weo+p+6qPlQs2xsCCNKCsaLwmmn0S8WT+vTUJLNtm1VUd
k02Ko3adZ3TTJ6xKOY/sb3+iCLdVphnKZM/KuWTBz7I+T0OtOd2QxYECYb7XkVzz
0NFko8ZivoZU/9QGlR/MNJAUhfhE3xt0S/3e/SqH2Jpr/LJ3cMQZ1Jt/7VAJS3HX
ZDJBF4KfU+ADfJWgpfBOPhcN8+D9ddEwFvgtHa9vbtHdWZGX30zLsMiJKhytgJe6
hzae78WYyIswW/s19YTB1peceuWYqYz5qefqTMw9ej+XamPsA0FG3kfJ360zIlud
3XbWPLhM/haHhZsj4C51O/jmrICQ6LTwOT4a8Hbj02A=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ThbPrp3NR3J/ug3dJeixhZJaXkrARx0vFOFA3v4YXuMZRPof+VoaohDHdVJXfWnp
eX8aNEpIL6JhC+3Q6zKLoPqOrKFqiTnQj+BrF7VI0w2id3fx68ebY/QoaEAbxnub
vLqOKL/unlTcevVA6dfqVZ5m1msa0ux60Wc1RMjOdwHVd7TEf1zfLPTdExIteHJl
oaOSomEArp5yVHaullZX9ovOtW3LmE//aa4K8Qv4C6y5jLQDAXUaRAWWN7hk93+O
vDdQ0T/aEVqbp9l/0RKhu4A5NlTqKvzUXlPF9QH41tytMJ8NxYkrrqAysGn8F6Ee
Yz7eQHUPxmcP+9JPPCMagw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9232 )
`pragma protect data_block
ukffgPlJGYZAqahMqqrPYIdaTV4DqE/TtSqPbBO5XGgMWdQkYPwlCqUeIQuH+mM1
ZADmMh5yVGcgLoxNNiBLZIyinTuz9e7udQ2DwOjSshNPnwVe/8+AAiTg3lX++8H6
BCXSQ5JRzsCxt2bGVtCUKbUv4HaHDDMJEBJb7ohDK6k4hQmpFb4Mav1hUE0G6Cag
aSniYxC1qVx6Z1IynKceRdCDciK73y6q1TQNWwjYwnej2IUUaXe2HBupRyBc6DA0
4CuX3EDzo+cO4yA8o4dIvTDUjOdesQ/s5Vk7LTyLU64D+Yn9jGIFO+rPbzFeEVUE
BhyXGLltlPkm6GObPEjmXK16TiA0X10RR58XEVl4yFRDjxnoNQVWisf1krSRJOk0
zQ/ub0QJ+OzgiOUtG42Yrhl2TB8t+4g1lIfTcUDm171JLPQHVy1MrERranl3pCf3
ftbUqC736FHx4FYgdeiWxkcmHa4Vrnr+HcNKgGJeL0o6RmxsmdjSycPLZKI89yp/
OwbIx39WSJTobAAq929w4XLAeIcdrDvTXql6Gfl9cSN9JnYk7Pu3Fgl2Lw3YU8Hj
WbYx97kx0GK+63a2CLXL7lw681ivl4iGOFx22buzNhSRohKEVD8NiuhWcOwZisDs
PP6YPwV5xkE0qVAUxDoHjfe0MAvUKhAjDgTQ2BUhadd93w21LGZaTjbcdKypj0q1
N5tBm4t7i1kOtqZw1xuQKDNRLePBW1bQGcb/84cLsm6V3GcJeJXTNIeGlDF4bEpo
bpP+O0jJ/NaBlPZiZjPj+/7PFCCL71b+aU7Vp9f1QYD0r9zG4BSLY2G9JR5wm50P
8m08FgUiYWqSDjFSK/KjiqfsWkY90hoaOw8695vdLR6ZZ6VEo/EZVGPOZnu0p7Dv
U0fNIl2KTIFwXmtaHU+9iqFaq+WAF2hktaqiFJdNe/ONQK/Bux6Ms8b3+WskiAV8
x4TKwR++n2hZiyptvUHYNdmHRCd1FIaWoijRKghmvCIgTpeJZgOQbA+IQOtfU7UU
s5bsvRi1zU/sbQrZJIae4w5kFfLOOvs1rTA1t36DAfgtE1gxhdRVTDhVFA5mPjdJ
APGq5RSDmZAZ/yuM7IUc184u+V3fGbnoWwFGTiMICSFDbf6Iav6UHEr+OljJkUoE
HewpaigPukXiB8ELzrv5FsVbmJGqE2QQITcSiXoz7PuJ569BIn37vHDQHlc5xsTp
izPF79DnUtiy02jzQ1CSuVwgAoNL1IOsZTyeICrjWbQOnQnEcKGpNs7b9o25JmC4
6ehiiPGflCN3hPQqGqmjF/jrPTWXMhtFWtbSoUYSDwUPu2PtNrIHOaAozer4mtxf
eCivxWUIjknqoNf/R93HVQcx8mjxODjexHH5cUYta6IDzTmIUx9lyuIaQpfomZis
b0hwcMnxEoX7lyR9VpLh/XKSEv4/pOAeXMUXqQc9H7ruFLY3YLm58oLKPA13htHC
3Mvto09oDZHHZROCuH2Bd+mGuNd0eZfX5TsUt1lA/qooa4tTeRFUadjDYr+cEMzL
ADtjEbmz0Ei9tkf9B2mi5FhoiYpRgKefwuhWlCBFzqvDrlcyqF65pK7ZA3OiOMGc
7lphBCic7+o2OPMB2s6MvFscVfuNYLzbs2gCodZmitTrDRLtUtWLcvsV3NRCxuMU
wRRmWz4L9sRJk5OvsZmC3ZRSplSuPh/pwBertorM1fCqrCASknTo8v0rG6bOkKGw
iLxmqa1GtDXy90mgYqzLcE79JZfZWS47qSmyJi3Qnvg/7uI42JiqeM/gfgrJGMLU
WYtKhZkZJvkbRp6JA9S0GUyl2d36y9d1cr3rM8xzUJ727nbxAIp/7jgV2lNghuhw
wupvgWS8W/Sipc7XEe+4OJjO1pwl8G/T9Gf8Shc0fAUs9VLCWHHdYzNle5Kpw/ul
S2WM4zCK8EVZeKw5Dga4xmCUM3TOYgeTgn/cen753JpLjEFqnal+3jICdjFoSnxn
ztB7Jch7EyDOH4qToMMlsuWM1FAoBhYZW8tkNEMMYS+HB4Az91K/+fmkyeynl+95
Hx7keAa5Nu9lh5X8s9VcH+k6gyTaWe/Png7dBEoAerqSu1QH29OInR70Wwf9nU/1
fDvfbUMVyHgfYCOLxiZLxzJ4haEN22e8R94TdarysLl2FKlcLGW6OCgVdx9Z1Gl5
IDi//UUKGknJA0736VI9JEubU/Sgfdz3vVRcEYwRatMltLvY6w/FyF3sbS+gdsbp
QzxfHIt6S8vk+lsKZXzglA+oikqtc5T9JEOCFVt0MS76XbX8afOBLuUljB0N6RKD
mrXHAbtNrAW+i1adoa+kK3Tfa6aR6ad87jipn5O1BGq8dTeXjmREiFFQ9l6WEJQ2
Yg9ixLFyuwShZ90X4cDYlkWW6gEaLHYOp52KV6NI2p3qxCbIV44DJ5oB5b6xxpMK
TuX7w5PcXvFJBrq3r4ltpzw2r12yduqCWRaPz6ToihO3xuNqTvCxaWqnMlPbgAYu
wasi4uyhdT5DYeNC/oov/vFhMkVXmojM8AtCK9wfl/7DyPDa2f21fNirX10I4Qut
3HCKpL3tJRXy1t2mFBvGl4ExqQRQuRnZBfeEg4o8bQsCE+3sdQNLq1oxsIWn4Jmt
3866GEslCMiBaiIYW16npNZvGNpEwTuvtkXM/u7TKMU2lodpypJ28nx2mSglC9ZQ
lZ8SZVDI1OSG8rlCGfBUCWa7vbx62zBK1KqvimzvMAY4ppwiqsaK4xfPVdlE+JNb
MkQxSKti/GqgjXmPTVf/gJdh1hokVntoZT8eWTjGqfYbq1MRDxnbQgQn0hzdEsej
wf5WbwanZsklJp8GXDnHByzP3LdVfbzUAhJMc7XwAKU1VXy52esrkCseQCU/OyEL
XNeb4AhPnXFx2VkDFGCookV405DaFBlmUDyWIeRz4gK/3Iv0Pd9VL0JbPWK5ZL55
s7jiby8sY5L5u6uioKn/aOWYZC5O0PRfrQOehQpqnB/e0TkBZMOuBszyM7b96wm+
sFrDSwpuH60HCijIN7VmitBoeFfXbiT5cBJEi2xfjSVtYSrsVMpvRG//VoOH2JCo
bPsff13t2vrMnpABupkSPe1q6aw7rCYiSNs0yD1JRhTX/6tzTOSboRdmElXIx6Et
vok5KyQwA/xZ0ChPrVdEbVfXVD+dU3e82Sdma+rnNvYnKOrlZsnA0g6lKkIZaEr6
riPNLeCs/W5BQXwk5RMG0CxKMiTdkFbk76WnPwcfq8Aqyw+8WnK+4J7glQzS+Qus
CWPe61czLYr+ZRQOZ4qFHGpIBDJPT2PLyCF7F410JE4cmih+32k8/hcH0D2Fg1CL
Ucqq+7TnFGBCXSqn30mOorAxoL4jG7iaV4FG+0LN/Q/CmQ20Zq1wx1fZKAdxsUAq
KmAbO9z5iGKEfwMMRG+ehl/OXXwmFRYXcHcNkLzil0Kg5eHej8MSWMAbu301OZLU
GZD79swQtLXQE4MLkO/iD6Q0kmaa1u/I5OxL8iKfIlHSWQvTJT8qnm8piTUeHtCI
KJzRyfCbjbzbMxA3g7EaBKonsDMyH6pUWVn4BSvg2p8K5zujUilPo12fjarNIUFv
g750AkkorQgGewXj2AgzmK9BvGMcz1oyH45YANfIt8PFUKystmO/Qry4rNDlCMiw
D+7wvF3o2wD0XkB1TP/c02AbrVrn7K6qBJhPpKW3+OqGENwDNhwPDRmVKDzvVeI4
1APVfjWACeCUJseInZNur3oOoc7BuPj1Oxv7aDAvD+90HpoR0WjlU8fZIYYQ8BFv
bvprk6Az6MSd7teOsoLjzXfTk4REMtvunwq9XWOaVOFmC+DY6dcHAco4Ru82KHdz
L0HxUjyNWXhR2i3NzrbU2bi1wAYcQUDGVOQl5T6r1yl6b4vdkl5JQwibRclaO8o7
OjQVhMpfpgwD8PtLnRSBQdv85vChcxId6PS+OzWZCQ5hsWEI43JlOBdzDZaIueGa
tu5T/9J47VT7ASGhZi1/B9DewOvFjqES7fIDki48UYPJFz4W7nFKXvmgH1CUSYoS
6PMZqr72wVc1vBOFPEuTO/qBj38rXJ8HvqIa6LMRHnfc6TxykzZHozuArbXqBQH4
SXSc+EW3qO9XgMViv1OG8xEj+gZhaw1x1JjmVipA6yq2Lm5cedmvbkggOjmJQFey
HevgwSyasADbXCj9CdzU3Jly9pI90ZYPgCJx0t+wBeySG3GDmYifwJCtnQQhyIXi
dElCse9Km0uvAD9r1RqkB8DrGiV/w5qljxTQOOe7oNhVguUn+dZvCiRYfQt8m9ic
+IAXTNRlu1vo2R/aG2ell65pX4aB5rOosfLTnILC/JM3pkteiejRqAcwoU7QQvmj
b9gpn31S09g6Vp0tpi+PfsFHe9MvJ1hpqCU/OTXBfSiupVfs0Ju62vm3Ya3LcfHH
mOH2Xcx2HDKavEqzBDdYmhsTJwvANBIjWVUMvhk4inqbDEBfLHbz2g7KCbgRyaeL
eYSJJ2TLKbFdIfUgdhOY7q3174HurfwHGraLl8kDzs1Q30GjPtejW47vIxux5lBg
iZdDNMWUGnW7vmuyo9ZBu7sHMtENupPbGZSgDVu/RVg0g5fjJy+Lp00vQBDZH9pH
SVC/AKeiSDvDdrBHxEUp9G1EONf1ZUL0UBywUbexnKF+K8gt97CxxuHXirxbKRbJ
gOjt1ZCsuh9Hcfk2QussSE3I+mXLaWRoD4/CuxHluXTRelIcgm9YYdDrmxUQ0kEI
Eq4x8TsWpTvQQh+hw3IO3L6fCL3VNtsqJtFQpTA6UbwqXeOZ/4vQPc8AWeb+v58R
T7C0iC866YhtsPNjxj9Q/FsIprLXPzIN8nil3lCDxa8Vi72iyBBWreodtkzht29Q
jr0ML2xeTNMfSKn5a8vLeR/0YiP0foF87c+Gj8XCHCIO/dhw0T5dLvLGx53ya3dR
S/Y7dCcb37Ij++B15T+6F18rwHsMHM3wI8QLtzfDQA/9jGCJvjWo6v8FJEbk7VYb
TWNDjyGHw6njn5hryhv71HIImzXT4hEflf2fohxnYvr+ubXwtV5Tia8r6rx+mnrE
nAI02+T8pqzVR1BBbCPXT7DuaMXAkPSvluX907b/FQIt2MtVv+2ifHdCDNwnyQSH
2Yt2Q0j4l63fXJREz0vS1nGqgI85eipKiPRHxrprlDpjA6/TP5aVi6CEpui7Lr/l
4y05ALd1fRzH8juzqeiY5RZ/7zeUmh8eFhcsIOCY+9xPazquPs0jE/QMVZ2YDD7I
ZxA0RcJIJUwQcN+QT3hufEAe1IQr2ZtetsTHAeoFchoUfe6XLslwAwgqSfLoHjcM
1UKizvaaBxLYjVjbkzv9gy9FTz3NtaJhljDh6CPUPa4yg+UPluODNbw1qUUCku9m
CU3pJberTpg4mdbKz/h4uFraUtZ0wZMpKygwXFRRV6rk3shedxcdBlYdZ+DoaD4Z
jZQPCaFmKM7tuL3gXgajKkOPHf6Fce3oynuLsjyYRtj2syRQH0ttkLWgnEQ9M1fh
6XAmMYVjXpd4TUOEZ5/kTIZtzbmAk9yh6K2/nGi+xlLWJSzvdk4+dmm/vcY7J86f
5oYTirW+ZU7EoBiiD9WixD6/pzet7qG39uEXygwB+5CoQDCTKzw+FboJ/OrJKN6z
u6Ax/aQjefUBi/uWj23lgoOvBoKoj06baAxuTlgAti+i387Jgl4Qcgq9t7Y5B9Vp
84OcdzxkLErbF9Unvm3T1HsLcNw2FgbE6wvKivyk5UaY9o2RbFVL95UG1cFygx6f
wmYRhmREtUeUDpZRMJcupW2MOBeIvMjJceKy+ong0J6cK3xBlpdeaKqdMdUlVTMq
7zzctw98kZdqdggh1jbdxd2LNY5EROtE7sZw9naLFpXRt67pJ4RZC4b3sfoiv4HY
eUJWFGoOLhyqQXYj2N/ZP1njuzgXzSiUe+fxJdjRJQkpHuBNc9N/yLmISuSFJZok
crL6BEnx/eszUvuE9+dM+kiTLxWDw2ZUEiUkomsBLvFaCbl+bG/Mz3Es44KGaBpY
OTDiYbBKJt82aG5Dwe1MCGOunpXe525IAfCGk3Chy9/NVd+WajjakVrGoptBqF+c
VHORMUgVYILqtHUqDhn2KpiDbxcSbb4tY+iVmssq3Dxn+5A6aAcW9JvFVEw43vsg
BT04lWGwoWW1+VBxQF3F37VRPRNQ2JFCvCR2/70YlUJnevlfK1PJBut2cvb6K4lX
OV/T9oJAi7xMS8yzxAX+IaHBWjClekz5tktB9xsrs6rCEfpC1m3bTo56j719/Zo8
n93Cw5fnVRZPXMwtnP9Nfnq4AdNJbH/zhHHCLqYa5E71M9UTjc+0UrhvZC9qkhyZ
0VO+TneNYB4oR2+GfQCiy1OX4TW7ZLYi6f97P/RabBa3XHdJQyoXVe4dcOk8RyfU
zA1qay9DHg8d0zuXlQ/fwH8S4QAc7hqAWFq3BQLJWJqmohxwsg19oI5n+EUSm2PU
Cyd4lurVCd5tV119ioMGHFo+YbUzQVx+eo5uHpFP1f/6swrzzHhVmWAZVxlQhmx3
5VtOmEWnOaSS/eWaxeGpwGJl0CsmY6xnpoPWNHgkpfN0woD+XRIkpZuujEi4tm4i
TGExAmP74FL9riWin7WWg3Rxi/Noh+ujqK/+KC6SJGiVVSFoK8i8bJh3Smlz8PLI
VbjCiYveKaF4fpQ8UvkPThfbae7g9JVl6QUsAkTC4aO9oAcjwPXhBPZ7sVkMQej7
96tAZoTJULbWesmgV7fsVn31WjstpVoNsZV+obOxEQLtegWTkfu7v+jiLytRhsbv
3gF2/cvUeGRuLOFt81g1LWhErpUg4vc2BgOLpB7t4Z+2SDkhqcaHSVsgZm41+KsB
dS/Gp6EswG8cX98/IiSaGkVSdCnEk2QCs7/yuZB9hUpI/mH0TmaZRo5aD1c16Lj6
5kWDtYI/gyeO6mgQW6FWAsPlK4FMVaIzhhDx472+kSEAQ6ZfqnMAU3ipeGcyCU8y
4tngsBiItqhmjF0EnX+Umv+pamIYRaScUrzF6KLE9Cj6XZAGq1KmVSxH9MRvOgLe
OYTfZr/yKyb5jqt/kOzi58smbmoXsDDFnW88vr1T0UnePyson+jnkMYrEMQwYlhr
9wR0a7xdv7ElSSkHiGscfuYlTdErTxzXBYZLLCemJiHQqXGsmkcBptUZ6sI084jL
mcUVZCHZGzwxEbOom7kNT1glEBO2iDQcc+KsjxK3waWnxe1w9BAoAbFPPkOIJNLa
L7QmMgWec3IcBX27tC6Dnspkk+A5URB1hFaL8KgdJj8mQVxvh0UgrwA4u5pOvHjC
gPDTVj7683i5aymFJo40Z/7M6TYDbN3wjo+jamcl3P+hMh9oJ4eRtZ/L/z3RjSmS
5HHf43drZsGdm5PZKaxSzkLfnlrFDqQHFsFOA+wukemiu23XM47O6/yvxXfISY0h
0NJB4vFHhXp7lNo2/TPihqIqNwxfRK5Fg3NJXG9Zfn6Y2q9aSV5FXL/HIuNZY/9k
3oiULCBROM5lBFhPhaqXQPDLE2zTqB05Xj9P6qyBpnfJbA+9rGsHQHq3/muzHIGV
nz5rEb8IugN4snxhUxr9E7tvdWMYQBBrhy/cEtxB9DbKTH5QXBc5kLAfrn8ZLpus
WYHCRRIZ01S2+WBwPUXHaIxQnOAWiS7D6WXPJj3Bi+rO38/UeaJb0Mdo6CswE/iL
yi9qUqvtXf1sFaVnGO2pYCqRygR1ElJOVL26p046vhsxkkCIe1XazbS8NMXxZiN2
+UDNwvmYkbznk2zWghBU4Bn45IriRe7coPW6RMySmLzNB/WB2mXeMDFuclXgc3qh
LqgZqIMK78seiEfRQXEQvSIVRiXYwYNGZhGRQhEp/WdBHxddF0W3X58QS5dIroFC
ZU4C5OWNsRBlhyIDxcUTsLcr6hun741uS5bpYw6kdhZ8Q90Gm404fREjS52+9Zkj
Bi+yOtGFHk2pzM0bz1kPfkH8xl8TbGOtF3EzR6fz0+KjviGe+CyQR2WJYqLxv7iM
zO390j2W6gjj8yOQpHRlOGlAPMAaM6jsXbKvL5LA0/BxIan9aVOea+qPzr6mk/W7
GTLQeu43H6EpXSwtojoLqO/WXfv/hU+8LG/wiQotlT6789NhDRY+FVeFcyCcWGEs
4LMl/f4Xn7h1fBb5lfoZnu5M/cjsC3FF563paBPM9GP32CpxXDoa40TOWrxYYmw2
hMPSA6JQzdNK1/iYMJhoiZNvnq1/50eJwoZ442PlkYuom8qd8C61tUEz8UvIicfD
gSfKyIePD//h7DjVbRWRtEhaqP3PlKNgRYgKH1MlWDfoVVJdnRHCXxxDo4sFbh2T
TY5Lc5Zp2sQogwXjja8ZePbN5ZJJhwcFtXCiD0v4GepiO3mZtDgHl6OmpoIqmZ6l
QLbc+dY4fSVEA1uuwVecy8M1ogUNSMemSo6EcJB+0HCLjbXzhh4WFNvErWPKNvF0
Dhckn9p+/YhC8SYB01I+lKhUebbbzxTk7yaj6uZxUuweRZ1MkWSgIP8KJmFenbD3
vA9h7DUKAo9fv1gZTisIE+NUixt/muzluh7ornFoLYMc6G6veLWEPmcd2mz+gmeu
VwPpQVTLcMjlG0uzvOj0EOElN8awCK3w1qqxC6SXZH51+ovCg8h3aw5hYjF13MpS
g9OXfTYR4Xg+RjI+CuqZMFqOdh5O94j5sQ/HumM7LrkGVNeDXLgNKS8GEP/YG114
IiVIaDOp7VRjB4NhR6/I+7FjiB2qbxN9kUZL0WL0SGqEbQ4Dyw6kK/fPPmF21ObO
mnHUPsl+uZ3SjwtAQ5kPeVDob5qVr+5d5rT1cNBT+wM7j9/rIYkVZBfful1neODW
epS8Nh8zGcRGv4xDOgeOtIieSWNCRw69dmB1wy3O2u6F6MFjwg7hp+/yNCpDPMRI
KFx8sIrLazclx6rsLA9KJklbRxc5QCzhv4RF/f2IwAkR6ajbq704LFSZj7vb9gHa
r7OOEtT1S4xnpzseaPiEa4I68ORt0jLcle7B39k43HQ3fNRG4ozN1B89klcVbxXG
sWQNbPGOtf+ONhLvZtPqpy7dIltHQi+V3nJwUlwrkZMBSAHJl1VrW42TSC2Gwu94
HzrlbajCdd/7wYuib0PGPZ1ow20Wuyw23m1dLlBasjsokiCqmQGg0W3RnpVEI+Hu
XJkvEc91EXrIQfkZmJO3JAJI6qH2uQT32wc3/ZxDQAd+ehjX9xajsMJL/gyPH+l4
ypF0SuDLtHYObojrNY8+pBICaFF4OMMFfvx6OjuAIXO+FZF9koi4EZCHMtZf1IBu
ps5+SwSKCBVG1iHVqAzf5cJEyRJDCfirbmVUBmSl7gdbdMrP2WJ8g4knNCZBuuIG
NT2qABJfzqbHVhUgtAqfxaYngxIgeQ3sBhzoMxoKRLR+OlSha6yyevHArHvDEP+D
VVz9F+Zxafc2DLw6qhs8fnu57nKXJZUKbAz5luV1D3bEGl4O/EeSimLsHOHzrUF2
79/zbgJsreyMCX7oDdxEC2IbNRohTMcWIb/9UsQl+cUls+IsHMeKlkGdwb6HWofa
VmzOVkOeDPzAMQPV3pq17mIqLQSCKrUNILw2blp4yADZh9A3wRzNeOLBVAlKXwih
2XUZjy1TqXgxD63PirRipFv8SXsBi7tUR7P1+4E4ONdkLYyo1K4zrtKQoil0KgHn
RZZlJYMTLpx6PNEJ7LTp28qdssWu5RXXXn32GW9I2/LjdSd3BSy2NqcIz+oT0QA3
ZKzjkgMNqa2QEl98Vs6PqIHKrvoRfndQ/kqh6damOrVB/5fjeMkvwLlqnkQ8F5Bn
n46hCe9Uythc75XMCPFhZmXZRMc7ZotBu9JHvy5VgKo1+08C+7raxExP4fzMNR7+
YTdmDd1QzNP13WZ71Nro7mf/L9AGGIisz1ductYwhs+RJqBxSGa4YS+ooadxpejV
ht1jWmrYD+VdOhIYF7Vd6VQ2T44wpl0LRJkdNs4SX7Ngmj2fOenmS0zM6Lnkywx/
aym52UZRONah1oadH00kAy+9N6ZDMylDvHdoE/CM8FS0OTII+IqwBAgMMWe/DEdn
/Mjrizc/mrFPkKx+mciykJHu1iYjuPbHX8zYzcMbFotIakpWo5CA5tEvZRMpyQx+
obdwNW05Wajsh0MZfPGIxd2+hMrvW0znltPPEAVOEBtp0ILHGD304fs5KALWkc1y
5gffdAFHdDD2k6DRBw9Dn6ZNW5Z/if2mziuUiDtJX9q3thuftN3FZZxKu2NVCcW7
dFu0iXqKyjVdGHrruH/QINeTe+/O2g5G8ANbCg4ceOikkCrBMdroWpBrxzH7V/+E
E5VfRZ9n+Tsy08+qZ0gjn5XgDuCnXQ5msIKVNN1Sy+sJKkXo77AOEe2OPTMbqK1I
LNLsNbkEAqZIKgtJOZz0RlJbcXqcGKvp33aILX8iOOsC9wSDuHp7miifzse9jfdE
J1mEc1F5Eg7vaqGBoKqLEj6LHo1yrfZBkNVZkeOwXO8DAQallOVtcqPcfUHAg+1N
ocggMnTuGN1d4OAo6bVyIzsth88CO97tVFpWXsT87ELTR3UcXjBcgz/KOJZQu+I9
pPKwjJvjtETObShEiXXSUFpY5vKDPF+WBQ7m7Pp3oLmZNm/Lm2R063PRqieIk3lm
/rieh0zd7wmypWvwElk1cc7VBJmvFOOGSmSI7R2B4ItP4RKSWklNguWjKMktVHcZ
evp0HK0btRN70rE6E4/Y1NUuZKh2hGhVULBZanFjYdF2mxYAAYZmyK5zvMxPufQz
s2cUz5WzpyMWlUdIeN7D9Lo2uaK92hKiVLckNwswAiJV+aH1sCVzTnqxKh9IJXkn
2+HD+VRYlHazs8kGaxcLb/na0Xh8ND4guBH220TkFLMCdSUKtQg2ae1JH5sRotOk
3+AlvErRUz55buhIecT4MPKkFDb88NWa4HRagBy6utv9vLvqz3NRt90bmlQuxhZE
wt03+Z8veaXbTjyAYTJqRfLetyih02ynSNbdqNwlToOu9dxNfs76xDI3ysfT2abt
UScAEsoUfpascMvUjo692uLsVqsxtUjJ30erUgtEi+y8xbWXjZRUYHkK6HREdlB+
wbDXMC21ZP4PyxvXu2FvJSadpOzjszi0/JqtTZvZpXTkhbRUkb6i4IdPWipeGdzo
X5Utvy8V4L4Jv2NHngUxYJbAibS2y3mLZIN9AxFazTHkbpNpWY6dHe7skZ+Oh2dr
/ZbvtBX6xz0UssLoL82X25gDRDCXFnQDLWYRLtsMawziiX40a4asuOBZEyp3+cyM
qHRJP2abqXoPSLOYmz2mqUULZhVZrp3v+u5sS0TK+WWU7LWd0MS+TC7BnIZP5Rzp
2ISIvChZnZ1H/ejpj32MhD8kk+jNUBmAM5tl4ja4/UrBvFAJJUzC/7lJlrbTCah9
smu+Sh5e9N071XuvvZG4L2O8JZRllSqYl6B3ibw6Yh4FE/pkrI5yw/3x9EZ/3hFB
4fa7gSLARgPdzsz39lesXuAKM2pjxzrwpn+0sQmD9kW1c/3U2+zpHfWQZCGujFk6
Dp5DJ9cezJBy9yssCKpT3A5lU1Rp573K/NfwLlGwLU0im4NEbR9S11N6QYJdx4KN
IC2iLBldHvUUWGTGdYEAp+WMwKcsm5yvmsxXjyS0QJTBAj+P6ou33kLJgVNCyQ9k
ULy9pnW3FfPwwVY+HT+kTmqebk52eK6ldYmjQFKOt/cVYIdiNwsvA/YWW7bUp9U4
4EPn4U3nDWGI1BpdSBMmuqF9q2oyGOkNZTngwOtrbq7qMj06a1APSZjHYCs2wwkW
bzr7IP4O4c5HQS9P+hL7m/7AiTtooGonZsjGr6vhYPsnWso+a3fFxo/VbLR1WHAk
G0E2M41gDMSEUlbBHc1CuZOZV1NHBSoNJ5LWrxKniePGBqmJB/2dhF+xhzdnmRKY
WEudoKuSzwJaustVbb09Cs9bw64L2u0GPXUoAEr0r1miRJqhiw/zj8XIDOUKf+tl
7fwP6gLilPuGN0I8G3EaLN90SdaX8J4SbunP1gOFGyuQeToGJ1JPgrmqS8iInZ2N
1uqjuhaNXAUEZyJUJt/1DgfPT1luIdTSxP/VKdJ61ZSpjkAVGTGd5n3OZJ3MbFuL
Z2Fzb1bT+V5lHGh2/GKriLEARd2X6AosusSB5DBXmv9BwiVl5DZiw1D/9GmA6AW9
rieSWcmyBNFj0ZMOiWxpDX624vOnncvYmj/ZfsTjjvQcTQQfadNxulXg7iWJcRuz
QqlGm+jWV4C+fXLdxoSpBMBT+Ii+qz9UjSZEcZzk70QKCZck1Cs3td9IBB3GoMBb
s4s6m+XwrOwvm809T+b3eA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
B6N8EYt0yae3AamB82DXAWeFT8GV4YyN2I6FcF1r87TMndNWFXcxs4zjtNsKh4sa
5J3W8E6RiZyUowHKgcSs2jSGak9mploEHGkFfWWdgbj/Su38hBbcFE68IN4XHQBY
IJi55siC/CcYbiaDizYxLYouTKjmPoHMnLUGFmiJzKa23J3MeAuxObIwIKjM+oO5
yEVmvy/40GVF+ccUv4HpC7XaUWAji0XcRr12FKhj9hyvaQBHYL8QB39uQ2KdvuYt
SwrOgTeJO6X9YdTazhLEFSwNHGLL/zkHAMuGe/3LvQpMGNxfCcLI/TOl1skm/wAG
DUuyILcV49zNbrNzu3VEsg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14640 )
`pragma protect data_block
Js7LhHOiAhcv4HM2C7Kmk1rdMcuSJ1erVx2mkmOUPsZEk9OA4t3gs3A35xoamzZy
69id3dXKXn+hPdBZvFLYWPjItf+6LbkBYmy6uQuEedkKhTrr5i+RW3iQE926y+CC
fVyS1OPgzTZBP8H+eb1Q23+KQEEQfUUDlcPqc/zctk/VfHZ85lqoZfXcPdrK4LiY
/WZHC7YmPfFCCuFl43FdJMqUM68W0y0+Az66eV1HcAsJTz7hD4Rf2drJFrtaZUvr
s/AjbMvDU5wT0jNLox2wWK4EueTIpZ2DQiB3kXEq0If+C7B/eE0doLcMBGSg1Qlz
cddUj7rsuT1O8ZNYRk5DRxUGJtaWmq/XVdFLpeUc5GEVEb6XFH4YYyVudAnEqJ4e
QgHCQ2m0PFX8VAgvUd1f5nszh8dteSc/SZnojo3NeXQl8LdESe3ENAnO7IW44Q8T
j3Jg/gK4/H0pSQw5dftQ0iyRBJzujPn1uwMP+daH5yXolbe1VnwpjNXM2VJRlscB
TrqeQSrK1dQlRRtYreQ3/oru5XXTlrV4voN2QXvwGhLn0Aa8+wZPBdZuIUxbJsRq
HG/sx7tanMaNFjR1dFiiM3WnH9c4hqLaIk6p2rusty5l04GPn1iXvR6XBIetknm+
wIg8G2hDdqd6/r0CRgFXz5hFoSiM1/S7Yrxdr61PzipLsrUa77pDNvCu/9OHqZzb
VogTtpRgGtudgokkPHqcJ73WyyQuwndDm9DJKoStLvN9YWHq9fRb06wIMp0Bn0fH
zRkyNAXbrir4y+1FbJRNWk55JX1UEe/Uyaku+Qcvjfa+h0ZVTZcMX71vz+NdLeRz
MfZlMxn0/AElAkDcFaLtMBbu9sjRyTAZz1B/tOMQv8Np0E/B7PAZL1fGn5qQYriB
E6Z113k7sFHgZgNiF2buFlsYMzX+MeKPFlXHFZINXX1ie9v2SEcvngM5ZkcjYAaE
1inyUzpcYRp+xDp/KaeUM0ilW45eXwwObmKIoFAN/+f/lZq1/pYGYnYs9n09zTaa
NG3XoBVAvpvsYGHt+Lo0MGO7yzXqlr6lLBVKuNHZU81asxW9DW8iiQcrMPX08/m4
YnOD9AG2bjsVE+2wYovI4ExXJvIrwUl34diDgorr4Xj2Rs+COM8iU/fT++8SxlAn
zdEmU/AWkTeOVaNluTpuPGSqgyV+nTZJFLNc33TwX7TeGy9K8l2/2WrRmwZSzBo/
B4054+Y7ioYlNHV6qiid8fJZHw39bvoqoEUQXc5yh/qlSmpGq+Ygf2QTObHNiD76
la72kE6Hn/ViHGZDxzBZe73SGKNzVtM0xgUFj2j0/fODJxJFwFwziytC1Dxx1uJc
BOvytEico+Qzkot5oVyW8wYtUuPul3ZwLd5EXArpVxkEWnfPgD0Lo2OYkUC/j1qI
PsVaTx6gLwa+rDuynpKHKudG7I1PhwgG+iYLiad40dgLlQ/KQ6LgYbGuEhhgg+B/
LFAPQoad9HiHk5IXlXMdQ18jvFN1rQjdakJC4pJO0qXjERG/urK4yX5fwAsl8j9a
AXrrNVdfGmEZnyC7/W8IjM4Ur2cwOzMLUeBxTspibbwF1mylz3TJIKkPUluJG7AD
2jfyhT1nFG6/w3s40LiO162qZZBUrsQ1fgrq2aZxk2VuAE1HY4LgDRMmQ496u5Ta
3TjVHFw85kwTMOYjhNjyrDcpAIedaVgkiB/sReUY5d2otcbWwWXQXuruuGjdPvjf
vgz9aqqGvd0IUQWUof5Su53QjT/bA6v8R9gRbPU0PtIb4JrURccvWHl2UYWrZExL
1JWps9/Y1s2Cn9/BTt7uSIwhD2P/JLRwK7xXP3aZzqzeYc6fM9IGtdepUD86eQPc
nS8EfeX755kXuryjfDqP8We+eGH9K0ylzOif0AUCTXmHbFiQRIPt12d3+aEMT5xr
qA2bz3mHyxoXszNyR/mAHPWdBTYaD8ub8TjfhX853MFKzokjHCL58qgJsR2E07mp
xU9KMLL3FSyd8jM5xL2DHjUkqAjB3laEveUJOKMolrhWuhtONv5OPvRiIMcpMl9t
8b5R2RyUEdlBIy0/QowD5/1Af6jZwOpONNUrkpxTuEMTDhmS8XosL8S8yTDbjDAJ
AUKSkjCoxGmapYqlqDSfqaGaIKhDchBXZkUcxxqmGiR7wPEgqEvlIpH1CllDv08p
/78lB/h1Z0dDoK+9Nm9+l7nzaJQ1egvj+tGGugI00s4+IAdR4w+cMmCUrpxDdqP4
q8n4lZsKINwi/ssWpqno16IPVXjjV4SMtIM1wNbExubcNOJJ9x3M0oi/MqK/R2L9
f3De4N/5ODOXwvf5YefrHgidn5QB750I8mVLxBzNKLyfs2W9Vr95/2/ppGxoOtdO
iT25TaDG0N8K0Z+WgBDRqTtw7eF6TgH1blgxlJALXy2576TSDKNh4vAZ0gj/U2OB
4Hk0Ex93n3EDaBM1QKztus8muMLBBr7tjM2cmvDmTSYZXW41T84nApiZGUgsNxOg
xpL4/OTMyHlmHWjxc8r4rAolZosmP9HSPyF6gtqm6+lyBitQt0E772Ikxi3WeQKy
5dDWTQVh3QHSn+0AznDVxL/kcivW2uOkEGYByfMxMLLYMwyd8YNN9b0ZTISylEV8
OgdGSsnwS+uxO7/UtuqKfMAKmyzU+danuPJsbVkXmi7i2Yq3y/6HLyjBkFCo6iul
6iaIJkezhE8QQeqOfh+hW5zAf9mmE3/RuTzu7sLW+EhA1PsnSdZcEEprKMRlXc09
dENvngVDX8zhwcuuuVL4LxZ9kaJ2LdPYx5yBydprkr1bJhvxD1lgn69uyy4XyRMF
Lqt3z2r8+yNnepF3AiqLn9W9BX1hK0p41IK9ujVxJ6ScApB5r/UjDwGh+LUSLnhp
CassvLCZQZoYIv/yJxhJK5p4CnTtA82C0XbGt0SYX+PQ9e18P3NCrLOIRlWAMSDJ
kIWVY6t50s2jof8/X2yDr0tUUBx0rauc7hV8NiW+82YUblXyA0vj9dR4pfroiWnO
hfMudbsbUVbB4vHbwKzhEz6xbL0XxDquYLWIa1lD+W2Wpm1iURDzGcbYKu8A0Ycp
XEo9vKWOgZWLxQfZgR6eSmxelfcSS1XKXEM+PMfnXdBkPl2TgLAHFkTl/o0xbhHE
gmfkL9ENwq1vr5vtqlpRkzFpIuc6TIY1x6RZjKGT/DGfZve8hTNd5ZHX6WO+50UN
yYlEJJ+qycTEpooxaTmDYzzBLnahiDJ4/sZ+9N5mAo9MP0Ub1OcWjyEgsHvsbI2i
JskC9XmeoZa9JdVQnitjmr+t3g2lBe5to33J1nTrFOI6dRUqOjsyrBgLBhlHQx/E
GrguefYMVQPNPQa+LPhZS+XSgutDpnTUP3g4/v9MmQlJyZa3+R7rQaIR9p53kEuE
f+FGmem4s+hpP+ejxCr32yTfdCE08dN7b2mUPgUrGOkIcBHVh1ovKX2nxoVHzECe
GCZBip3O5Dd+Fj2CMr+Gpn8agAI/oLSBH3bbWLDbF27bG3d3WVRvlJSkMqJ1M4PO
xd2D9dE9agAu+l27bBoJtbgwm4QPiL8YIoXXg46DeGjIZpjkjHuteYtoPBIeBpXs
fyEZQ4kcLQdPsGNdmnTjNdutAFar4A4WW6fjdPPEgOU4HPzuFeYUGXEUAjNk+RM4
crQRnjFcECc0t4LzeKsGirU3YEQdBYvqysVWCExMXqzX1nRtFn7LVnyI8ztzO5u0
d2uc0xOjZ20RqF/8VT5yTt09Mku5DikfPtz4eb8Vfn+PgDB4rWBQ961e2qWozv1b
3zeZZZERnvspqVRGPTPix2rAm3ZAh44GaXFzSQ0088ywGOuOw0Br2QaXn6TMdwlE
FTDDiE65U2Z9nTqfzJl1wIJ9Y3RM9fh6GSuqp7FepVm5G3iOExlGbbZjGNajDSZS
fpKVaOWxCp40FqPlca771oSh06fHkNuGf+lkslZYDRFpqF0SijlL8A3jbevdGiMV
wuzCqm2mzIS7c1infs5XqupQzfxr9gbKoOxS76KTAk5WAJUy+OHjNz53wr0lssnn
j6oIUsH7nY0mqvQrdg209NTK8y9jqlW+nUsiS0sbLtF6sOZeS4Cz3zRMFtVskxaX
hqAo64f5oz9L4enmLVd3hUi5xeVxUwr2M6yjqQZQeIqXRSqI/Zw1qEhLTG1VJozj
dUiIKUTaitegBBfzVrUxJ0+ju83Oj/U7TgxwkRRv0jR9LPjyTe4VuhPF/Av1umiN
37EbA5MBFC40zj6iFT3uOGJIhSjST5tGnC8Zw9FSpqrTIjC7EHA2I8vfh46egK6f
kO4Hj5BO2x0EkBB57AvUekRwP92jPfEjSHLDo/s5POwpnXMNR5+UrfjLRJve68EQ
Sorr1fn70oy3KbDxFFurgmfVn2VJ2ANIHtRnu0/gTK59baVGtyzuMbMPpK8IbKhh
tAkdbVF4R1e2EG+x81T4sNLmbFTSBsePfBpRG/M6P2ifSR6IGjPHR0FuCxDhwKJw
AcEQaMUOxwa1TpCscIjYxkXYtb2eVcI3ZqVVRy/29bhKU6uhZylHWleWTwLyhXBp
9X/3+7KVl9tD3KjohmVMBqIvsG9fvq2+/4uiWpPK7td0ZrbCJAmUpBHeppr9sRWq
4dDs5a1N06JnRitBOx9YPud8pVDKJzjLsqfX/v9qcsW8VmylpcG9z9jG9nXRGAdL
43Ii/W5Tzw1KGw5hPr4sHCQbPFNOF6XXwGSLqASfRHiLivyfvD3OOpdn6l9aALiy
0tgTyJpLaiHGM8swdsn/nIid8uZr0eX7C3ngLX5Kvo3mH20T1z3G0GE61yrEgOqE
f8ikg4ERWe/kUBvPbv1GfN+wKCRkedMWh6DDV2yq7fDGRL60LVyeNCPeTythaMFU
ff0pJfsjL8Qa0J423C9kKP0QxmITdUjBnJc+teSuvNQD6Kh72aJseWPvxP8gp0qs
zuAKsZ3YE4Pfmq09k2/hrcUp7hKGOlBYEbvS0L4YMD4a32+wW2JmXTWxjCNyz22K
7r1pU4BcMLYbvlKQ4YMEFulScqv1A97NiaU8a4CbB5Olwy4k35j45Rqzg4lxpCcI
U3bMp7wv2u2vdsazVe8za56ijYKddN8fjHUVQTGakM3OyDEvSoh/aRjLxKi8e9X2
2/q+L6JTPxf00UW7YmLBTH2duaFoqToJsB7EEUMDZSKwzaGdXZlmszcqgz1w8vn5
HaLYOk7aBMAvrz1eZTfUekm63C1TuWk5bmCLwn32djrHM4xoaiuiaHlXpdr5WKMJ
hRdnTkUcZaVIk/I4eT1uj1REyfDZHKyOAB+1ASYB/si9czI8db+IYoIlo136YouQ
F9cTgX6IW4VidkTNJYOZLiYFUrA84t88yaw2U1oOIv9MXzsi0mYAt2lLWFaRTfWT
h++dXeWGbqTkz30g6aCVNgaMhHqfp3qURnwKRpjAdx0op25tKeHX7B0R+lmzyD4G
AGj9/Ie09W9KLaeTlPa8c1NDUniS3QMW5GW1QazuOtVSNDoLXHOADbtChv340N4M
yGmeZyelZHoRm3hRFYl0ymqmbgEyhzrv9v7XtwcE6Ak7VxgH2bDjNrXdxw/2iBJX
9fuw7JNSdVKYqjcpOusMwYVLVnzV8PeyNAcRnqJUUJlXXEpg74VWinKyYJ8rfVUb
1hPWsrNUCLR165EjdIx6u8G5SEGyEEKXJRBDROjBeFB6dj1cTagW42UbGmG0xIU6
WB8/xC3nHmIt2+0j0xcFccCXyfzLQXzIHAopUga4Xx7kAzUb2H9+iqxfiDRX0IuV
8vN5OgHLweACb3PrtuuYcyhZZl3RjCcHxzq5LhuSdUZNMM50Wj5YrfEb+oMcQSKK
C4SbSxZ7+o9rqqt/7VO+qp4V2OYIjaDZV3+EiMcQFjanUBN7gEIQ6LAXtbrTQsYn
ClkY3Eb+omXk7uviIaiJaFM7IWhGtRw9eljFFqxGWL3psrqv7VY6ELy04CcdJ5BV
aDo3WL9CXSByM0nI6SjQmS6MubhoEiICaWgCLcU6Y0m7t+Tbw3Zr6Gf9b/Up5xQI
hKBC86qOXe82ma8CjPzP3AOGNw4Ty7auKAScTrksjsfxaZss9oE6TpY/rvbKtJJF
oVgMmAhk4gjXtyRhtdd1AYDf0jIiMxdJcJaSz6dpcObly/TATcgDnz7RIwTsUZLA
0MNRRqGEoCV4Xsatw4QRQ3/6sQPXjOu3Xgdyd4J6xZZYnddmJ+s0OUIeABtJ1aQ3
/4s85LPS3zQHOz08A0QIDqU1CjpF9wzyoq6yaEYTV9fY9pEdWUkLeJPvHLeta1nA
QsNogzk/8tRpskUcDM+SSWIphjGE0pEurXB75RQbnRVNv95MJc6RcecNVqpeBSTl
+KZ3PRJC/9FV8ENANPnmVoSqqf0e1g3XUcKLqAqYL7GkdeuOoNO0NVuBp/ytZY7U
2MlfWZeTga60PVurnjfuaCNFYy2j5S3QdYB8fdxYOZdfAqTIbf9kNTfXKdSKi7y4
qQzCtPfn9v3gKQ4JOhxe5MdepfghjvlMvwG/QgJ+yuvGyay6O6+eQ4ZICuIFoq29
IrDTGLiv9Q9EPW7zhjm4r3U5EvQkCPJg8w2HGsuqeQRBrzelI1Uy2rogTv871RXH
pEu6EFD5U0/03nr1/OcVBFZ2CMEx4dBJ2bu0stekvy5Y/uz/GZDsCjH5hLS+ka6r
z6pk114cxDjLwvq6R969ZGWVLF6xbbdtPobeoPCcM1uu/sj8i8q93lVaagRJvi86
SZb9BlkWdaPq633cIYWwyEqdVXJgLtZ3BSazIDKANWT6z/bohPDRxwHNBLU8DRb7
ysM0Q3gRIr7lNcxvcAV9nrNHr0p8Qb/1OCz0TxXkrJTRMiU06/aE/QUj0LqvtZ5M
cMVDD1zxOevow5eGCsq+WNeAAiFepd70RGC4uHZBVGBxTAWqBfx5A7Ycta6YNQU3
KovUSS/zBg7hlA4Q7h2kuAG6xrcony6AjwT/j2CpSoW5VFNxWXrpPiB8QJJCPxkq
XW1TnOxLAj7B7afBGool5A03GGtO5KZQHxQHfSiAkT/NhpzPEQmPGeugP/nf1dEQ
BhJ9Xmie8wWkvzxRdDGMz7ZHHLi56hACi5Fek2XopzaOlbohEXkIHhJcBDmcmSfY
u//gJeCrb6sfx2IDztTF+L28Pn40DKSsj1F718MxOJOBLsT02UB0ox2DLPrEOlSm
xTqy3FBIW2T7LGfLPLRbh7Mu19wkFQ00FRvmIFwRGXY6ICr/4Dz86OWVLrmzcvEG
U70okxmZVCQRmn+olLcGKT/QF64y8itqoSflpXJhw9kar5ORoKx4dBmgYGJtagNY
HpsvP4zJW56klsKQDJCjhC7FOxKkmTFcz8/0IiWgBSt1Vkqd3BIASbvaVUuuE9m0
FygJcQD8RdNWpj9yzbZ0z4h7gYoXO612wxyCCK0dSZpP17/As9AxOLgJuUoDwTOG
1WbjHyLaiIj9q7u9XWQJRTlEiXFWwNRmd/kecVMnq5jb12yZySiMXWK9qkL1AMm0
Kw3V9nayGOnWKPEOmBNv6ocWPgMiKsL8yNnt2QY3KWB9Gl96DyyfQQ4ovD+1h3NX
/qmuB8nItTS+VxkgoFHv99E9OhhnNTmaTmuM/oSavvMJ3aghKD+k3aFX/elVcHYD
YV5Yfp1bDciGeKfupKyCaHbW/8dK5wbrAh2OPjYTFw1YriIAgXWuy2rTYjmJ1ZXU
uBfVDQv4GSt33req4DqDorG8LvoCqcqw446/PrqfZA7shLongSr1gxyOkvOJAd5o
sbqe/oTqhbN5NQoRUfpgm7gssCwiBrrqxLWXaGB0QIzj+yvv0IddDpMHKLcsdiVO
vY40vL6tw6ATL4x1xiDbnJYtftM/pOD30xM0pY1D+TYGFQHgjenWyev6++XBVZ1Y
LRW8Zx5bPKQumtvAV/K7HhSFs2uQEjsuabA/MaLDXYLgRMMhZuCdcGa10Tuiqj2u
9mcK1lWV/14siZEVhkbgc+gZWaSnAO1MDWP/ylihpqb7+jupEzAbgyzElWE0NOLt
ZW3ThWNJ48RUP4kqaQUMI6zRKFgrVRKKqnN0Mya2SD+KyH0M308xHMQNOl+BUIkn
ZKoCF3gmAS2m7rmafBdBXFC0mn2m3jLCe0R4CQaivGGRmJv8YJDi/gz+S9J0oxbI
5QieuDW1J+iEjDW0xQxggsrO+lHveAqhK+hqTRLIEs7VL2/OQRI7dCbJBIEr3Bvv
nSD+trJXR12pn2PJV7Zt+F5DBNQ88YF+5R0dme292JrYNGsJA2+BIwnv+CSd/Wp9
Fb1zxl5Z5n+nxtnUGJRFOM1d5M/jVirvShWcS3+WTiR93WhumEqZdsdEsQJNVZF+
6iTNEeNM0PZKVtu5E+V5l1RsEk2+M7UHrzCARcUgm+K8QRbuMmfJQ0bqDm+LfQEk
xOmDMRPtR61hTmkhBT8Ra5JvZXo+mVxaxJEBgK3Yhh1rMetmbTZW5LflNVfys4hX
lQBQLAtThUKkhYhxKyEnPngH42ZPHB9jM9YTv2lya1/Ma1455hAtF4l0WWAgt5F8
R0w9R2H6+EKXBwXy0N3KfZPZ/wXaJ/2/HvO/okVUWpAVtiMv1a/jc8y3CKRi84kA
VYwRsfQzerioalOH+kxSfovmxlZ/0nQxtSAo1zkymIU/eNgFF3+rrfMKtijXJo/u
7ddgD31usLEeNb0F5yUrnjxygqNxI2Tn0l8ReEj6NyBoXtQpFv6XNIFznIQ2/A0q
Oiok8r//idGWyw4y/hlDfA7DP6p26pEyIGJYXUz0BL6RhLbRWe0qFtw0LWIXj38l
wYBFsKapElZsVSwN0wqjE/IlR86SEgyrYQ1nnErD+9Q8Bm3OM2XmOjdyhJJ2S9mv
Ju7EKZZrCXOAtDB2FhxEoG5PkXqyhD0OPiDPpipzhSBTHL8/0xQyQ5Ezdj4m202v
h8ETa2ucaBpqhBAoFcIPkFawYggnfRj9uwXWJqWItWNEWInjxoYGAlM9XKTva6c0
jYTlo2gI3gk0z4ogJqgNZG7VmLcwccA29OyHxDrZBRxkgBWPBEu9Hd9rU81EyPcH
8qMgGzbobZFWJ4BSl8As6ugtauJKtgdcALg9tlI7CFjFGObGKh2fz51KZfX206Dy
lhvInbdrsaZ9wnw0NMwW0Rdfs6dllFMjg2e63b68dkNPrvkUNOueF7p3g8pSRfML
EDtBnKux3xEmj/5O/rIK6cTzk09/Cig4+aRBxSd5IrmzOW9H9RyjZm+MMXCyhA87
PyhcSfXC3QRHNwZTZA5MlDN8g/3WmFDZ6HGswoGp8bbVAHBY3lS9OgAs146tpQAv
EDn1YFbwi/HRVV3MRL14ZGMgNNpAg6NiFWzTgJ7gNhGM/8CrD8Ml/CvBACtklW9+
+S0U2tTGa72upthBvp46QONv9HHrRnG3w7ITFZGfnUWXN7d4CRI3BFNS2MwnvFjX
Ge+xw1XiWvq9YbVSrkGBE3e+z0CYFc95lxF6r7MjUILmq28cf4hRQfA3ZPMCKdvb
gQ/+6CrJvCPLwnVIINiDdGyYWDo5cvYAGKeMLeHf9DIOaIGpL4xBmT6yZEQj3pW5
vOgEbNP0cBw0gfBnSyJlOLaM9IKZUyYxICvZQ2heeUZM72xuJ8i3vvBo2wSC3Vap
mPwP+gu4c/bb77i8q4gFDt2JMD7ZLAiCOYNm2iuNjHDt2Pxnc57cbCFG0OYUPgiD
KFJanCvWxHtjbAqsBELRHviVvEuv4WO+fZ2RAhjNL6UzGm4uca5oeCN6nmQOJdYT
BwlPqZSAWSJCWNUnNtna5iQL+6/HUa4rl/pYCfWbspK9fX5Kla5nmsKfXIiVFiDZ
5KIMKQkakX+ig82D5XPhovMAlTGFadFwJsHXddBoNnJKtZ8fSluGjkCXSDfz1/sa
fRgmphjrZGvKejf1mEWEgb6bezpBPViFNr8ofgST/2fNFMv4zwJP/lPBGINyKG5R
uKgG20li5LKTdNh1vd6aqASzVhJbjP2sEjR6bDGb7nGMRV7Q5tkcvHnHolOmCDxe
CP3L8zUsK7kbUt2RWKdOANDH5BSQPNLbSDGkZtFoQPYh8BznJ9vAIKqqBLGibiSN
nNDbvBgE2Ft6ESfqBLS408XQ4Ugk4ZMnL2BW7MBJhuC0HeO5N7cLGp6IdTsM4mTF
w/B+YBWryWgcs7OZjuBrFfwyJqMYaplyR50yycstzPN3oSLg2cfJyJBTD2pMOMf+
tRCmWZOrNkna6fv4kuH+7aNeK7gBOK8+7rlkhwFQUrONJUzHyCArJ3qy98ZqrJWI
VNM7iyf4U1vCbaUMbX9Fki1T5Dbo3CRsxTTfKSo/RW8u25L4eiHmLNn/Z5MAuv5o
G+UVL/095RWJ3ZAsjc2s/X5yrrq9uSmvhAMrUmLKCJYckv4fkR+vVrXWLrZDsUgD
nxwmI1H5H/SqPcXC1b6YFJpzUnK2iGrejdQDOy+CeHmp3ruAA9a7L+1ky/qJ3syn
evLOJgUEsMS/Auu6elc9C36OovMttYo6lkgbpWpbJfmwuW0qzQPBFlI191VsW/MI
pwfZhvSE3ILBakqcfh+N5mfJesp2SFUeSG1ZNPtTMRj+pnwkkZIwEOhJu8miDJon
NkXW8qvFFQQ5CAB34pUkyin7gOp1+ro9jQNAQOOP4Fd516y4uwKYXkAElPEiZRTZ
kJT2eMfjrj3Mu23ic6d9OTLWOK6EmNrlbX+AtimHyRq39r/QIg/IysZSzwxqbopm
stFlgYlReFJXod7ZuzAwFvqpTUSZtGNB7o4fATQyAZd/atLRgMbDepA0U+FHTjLa
4giRDUZuP/iZBmpWWm+a88yTg9dly3n4lEC1PvUaju/4G4dDivk5tXEo8/zS6odq
PfMawErQo66bKRiHZfMIZ227S2SBxtHk6pwyMgP443zYuq4kEmeL8OJHh9+uM+SS
q1O5jJ7WS1Sbnv7m2QRz/hXc78iZosk/75p+9LxfVIGYa1+eYwH/wOORApt6H5eW
IRqJlHlHNAnlPvr+GfCkqiKIS9lW6hb3eIPLbK+LYCzr5GaPDSAbeLc0nyENZgAa
5A645DpLj65eCBcIYx93cq8bRG/6z6FeLekI9y3QGWbpa2npusrwB0OdXRCXLzWj
6nSIehs643bDrz6Oh2XTcW6xy8pPVbt15lLqKXfBQAMHiU9neOSroCnQVsIEB7CT
+ORUER+XIRCoXV3yF2cp9bLWxefhmilSyPtkCOwKoXtObFnlUbESGaa7wVzLJLBh
4aC7SObsrH9nZsmg1W9zrW3LfkSbcq2g+bCFuLbDqk39VQ5UjEU2gWCihyk4oYZU
m3zAoIzIX7FBJhpsneO0p21bFHFe1//XpN1VGdLfeHdqTnh+Oooc6qrZDY09Hpi0
TKSVDdtimU7UIavVhja+u3qVlmkW6tlWGVaui2rjMZKYEun43AlpPflYYolRawLY
fs5O6d4ioZgd85MhmAFBLL961uccTFTTPyx9+e2wrhSoQVikrlk7Kt3iTnjqCGbW
99nvMRpx5qO4hA+OyS/FsNqs+M+OoeozQOtp5bv44xtkmVF8JnwrRotg6J3bz4Ww
hGs2UBhxsPJvlHBlITtRTy5SBUUEHhFUw3A0RA/sFo7lfsfKuqb/KzpLvu79StnH
HD77dM1ygCBAPKkb6t6I3odASEqrNbj2YIYKcb6tVc4tXRWlNzQ/oIlRYGJ2aNcO
2vDNcmf12CVtdpnT9OOsDDxPmeUN/GksF1iBD+fm4rfNj37xZSh9y2E8DDmFR0W6
SdYXC/eBTDOOjcbYoKpQZuci8ZRlTICwvUvVY6R80NNe/nFHmfySJmIDvjYv2lnq
FZKsol6PrRvLTagyz947BNsVlDVtfBvHVjylqbvHdMjzhGVAZMEaBlE4/gvfMQmF
gj0slqGDAzgZ0s4vPGkSfCAjFEbzRAXwIei/AROxlwVej/2sh8UKYpmp7pfVC5ID
fTofTrpIv4dgj5THYEhl/vpJl/Lua8eJ9XYBSiTDDOTIzQ4PAhdmUormwOWnApgS
ptNvfLvo4KCwSv4m2ZBIOTfyBhQjLIb2HCF4xYae6gwiaH6jK6iPMkTxcud6qCvf
9fRXeUFHKlUX+ASYg+Opue7So0A9gvkf0+rtVOpMTEzYazCDnT6n0Tc3omdCbsTC
Xl7tsxlvmq8Gn7mlNKkPLEALl6jdTJFvpdZbiBbx/3M2G5xF9uo0TBvdjXczvFC3
uqJlEWKtC6kw0e6kXuLINmll7n+dGXrCBsI1JQ6YxcMtLAYLuvUBBtSYI+lMeALT
N6twRvbjSbCoiNky8I9egpuegz5qHq+KcmTM3j/88tHPgsLqjc86Zev+XtY05XwX
b7OzSOgXaEFuOl3GXJh9f3wicsrmVG0aOz92mF06v3Z21pv4B9yzThINGG7t57AF
Z6GkdmYah/iTQljT4Fwa3nxb5kocqyGGKwMcZ86dVOxLIosf7CQtXYto9Bx5Dnnc
wobcadRj5ekH34t6nUWrNdpf6Kio1ynb7/2Syl0/p3Iwgr3JgQP3T+rC5lj5klYK
rH/MO5GZKPtciDuOCNcGua5d4AS8EWv1BtGlS8lNqiUALzaAIfF5Vzb23fkHR2UM
ZtuqhZfSoJtDrHItOgrWrbZ20Qy/O2J3ijXzJwKps0vs2sjxwadGqrumu/9z6idO
c6ZbzI0tKLcDKvYtdX99EIP3kYxd0xIrXxISdWicpng6IePkh57JUPZ0T648WSI6
GEnHHDWWldvMBPiitPZxgUKzRN6pvXwit4iC/cqoTwUtV35eRiiMauP1gJWkrhMc
CL0Gp8d32RsrgYb1SIOXJwcSLlBOUm3fdoCWFN1iz0NOoFj76BWA/6rMFuWJfVxz
qhi4f0fhczaKU9JstVzE/0YfT0IHLzexLnPMLDf655c84k3jymmec0JPTBY09czx
FzERdSjjgO5TKtk8tIYNQObLah2xLRwDv6c7NkBqJFhMqSFLKIB5iiSXWV0Po7oD
gsdrfWkkVfDI2vfavWg04YvGbmaztpfInPPB980vlRVAQWnpoj8wRUz6go7sW5BT
vLljIydcqEwnVYpFpfh26jWNKhJ/FkHvme15cf2Rn5zRa10DbNF6rfZ+P59GuB1u
n4eyf8mH6TZQMZbCm7qFCmgj6ZKct6YniO3qzskGqZEHlCW0gy7j7xAE0Dojqqcf
V7ineeTp46JY5eDVUcUVZgQQtsAQuxfPCkeOmX8ut1nSQGE2kkybI9gwB60wnV3L
6pgNHnrfDJZo7mmmfOEnUYy974i6DramNzQKVZgLKuXPJMCCf0TLXVq6A5UT0jKY
OfjnC1VJoJQxXid7ySM5RVbFFkIXqnVCRaoMtw0NRk3MFIp+Nvy4nZIIxE9JCXVX
mIk58qMHHC6M09mfUqH9m2XoBKwBYwc5Er0teCAjxwO2Yol7ACs6w6Km6FMzpJQZ
Uysfv4Ijl/3lcIUCWzo3ynMZiH3hUC12N7RfltKSZeZvANdtnvPIg+ApixUl40vQ
ugZfZsm2DJ+KvJXIgsWeTy9445TL89SHZS97AcBKp2Mp6MXuuOcrLy0G04m1wiKg
RksTCJQAu7ubBX91ARh84amr5YBCziTOdbgrmNn5AiFO3rT2UFtt7/ckDTJGOE6m
J4FfRM2hqSyVBZneq3dQQ2AF09vVUXcDGKA4UaWhU/Sgbh5Lj9X9TofnnUbexWIy
uyxQhz/O1cCr5bNeg7gGQbxWKWGuBjOTlBwRcBQc7ERwapuB6/u7aK6CKCel5bx6
l/7LxRNcX23BZyfSH3srEXNFlbvoXoUJn519T1DaUsB+yvebrtRc47YHVmH+V0bE
1WFGTQwk0P0zrI0eLUW0a/oz6u+T9gUQckKUx6cm7w47iv3IgiQg+BtcpejJuCj6
8l1ouK49YD+IvChcOnnH1skq+Kp6MzOXF8fG3SjQuCmfZFgxjkbv+29MreI2ddv0
RTNkuPCBIVW3TPz1zgB2TLKGaPqUQSE7f2oOUp/2hMij0Uzio/Ehj9I4AMDPEvWW
hGNd6Wzk4uYFdhleIS8VXIRmf+fZCZYLCePkOwzC6iRyt0zUZHOVL/1O30NNMefB
tcJjMjBv+ewJRG1e/pqyXdSb+nG2b6yOa2X72Q9IYLn5pC+BxWdi7c1c9uqaOnpM
2ebFZ9mydOfubHesRtk/gYbC5JPTk4r4X6Iw86pLvBx6JthXNva3e9Q+x2Qa4EYy
QNhlHkrZktTNI7Bxov/EOENWdETTN4lZsvdfG39DWQn/oZz+91lds5VicoKy/hXg
NH0NgRLPCI1M9Sj/FysWXFAIqIS3T7ypSSdlrxQeUh0UKbEJYfyX+f97f3zfCHqQ
PWdOCgJdOKME38E6cmOdImNnFwQfCCvi29X2GK8eUWC5hpjFeQxLSkVXYFMcFIXQ
RcbJGH/OWhmqhqJ3Gcn6xqCzTU4mZ/qEH1P0TBwbl92TjX3JOacfwZQnDHAz2T20
fza7yuuRVnABDrgyv0WS6h2jXS83L/bzZW8U0P1p3p8aChsGsjOIEpZVrhcET08y
7wvGSUxRLh0QIeXcZaWCZDA3mb89pUAp+CeL8hCjto+rXJWkOBONxzRtwK3KGyOm
zJAe9NlmdNRDVWaTBnhlouVAjsoG6XqZA1Ixp4sXj6h/spummMmCbkME5PVoqJ4n
GwW4R1Hjb1l1m2UeneJDKVTngEKieNwTkzQTr+fXuoAE0Wnb1Up71WOOvrcunjYL
5eB9SV+EvS2++uFoL0dirSyb5Ub2ioODkzqjGJ76+EFZwSsu1/ka6/zzG4huRnaT
6yL/9BgSAYC8bX+vRT2uLoC+IICdxoTsHuL+4IDyigw9naQC8xNXt6bkZ1cmOs3Y
FidkHis1k8tO/eM/widBfA4qxbdgKmu077GRWhPux/26M7N02Q0ucEe8diKdwD0Z
xAgHyFvCl+3AMHhSDbiEkwfhoWdPPANgrfP+CaFvQqjIovcZG8/Qd6JcrBeeJb40
SAo0RPipO+iuXq0/J86YJqNOec7aV4G5MJgakdLyVQ2ek85dqiCbvt/WcPY0LjXo
ebBhqWiCdYN19OwPgKu6Bs3Fg3ke3q5qZDBkHL+g7CyMbQNOm9ztefqt/LYQN89O
eDYEDcxgUZLkNSrywCEzVWtqE0U2CVUgqHfUG6dSV0xTvTHDvClVx1fD7isJ4e1/
boCXMkCc4z3yLU4Yh/HJvOqk6POXJ/x3g2jE+nAzT0sZegB0+FpAx0uU9oH5YRCu
G6Vx+yPf9v1We2+3So0XZmHBMLfvsZ0C8ClLlhlsjwmv0x5mKicsi5Cow5S8Ma8O
rOmEU137oTW8LL4WnIOehMG139OHOdLXugS/GgoWr6f+4QzVMA05RiF244X6hb6u
4AhPR2G+3JPGBuCRjCAkzNq/RxDD4DjKqQ+nTfIQjHYmaCQLAo+e0/LQunT//i73
SfGDBf8hEi4mcr9H/GQIiZmzbRVk+TMDNEPKKuJikKO46VcuRtjNqZFEUCYRKonW
UtXQddvhjvXRtowOlkl8/Pkw+xqowrxrti61/NiRHN1ktM2dxzoEHBGntEbZYQ9u
aJawJZTbWksmeQTdL04UQ2wwnT1dE+wYA97zD8iycquS5PtWLLNcDZFvRTRk3re2
HAdQB8iw79IH8txYM8WX8f6uyQWfNPQcvk/YW5/7DhZHcGrbgjLbV9S7yZXCoGrB
PF8U8GY5QPjfqi29USYnpRLLvLpcBKKO8cp7+CP/F0XBnH/+OMjEfFaaTAkKsMM7
f0i2ShzD0pBoiClzeZ3iUMVJ1uuRPWpCv36jKjJggPKJWSno8qnagsaPmitOMM19
CNP9hkkLDU3U/v2SjGMuksYgkSE4DOH2OOUN57AOuL5RXM2jH4h0CzR1lBgJwhUn
YK35NkEPPDBiToKKKpqVmeYHZN8cjToZkNY5lYFK+2nJsN99gMfjoMEMw+KZXrzR
rac+qSWaKqGPNcn75rDwet353hCNb1zsYyHQhJt9tpZHB/LrLpHoX3TGduecj9nm
xr7vwSM3+4UjXGjGXYxTQ29CwN7Ep5gMdUAeofC1Ot4lG0v8zu77xGBPeT9gVyL3
QLg4YNJiiViIsUb6fK4f+EMAdZJhXDlL2flIinmbC04YK8/I6cQuPEPBYMrYlyMg
W5p6C8a22ICQxCIwLCj2PcmzhAAgBam/Isj045BNAnW4yStHAf3PAhqt3Lrs78FI
WtLs/A336yTJhUdmKgio6MkcYMtBkOLjEz5T3lUbtPcIBurTdpxzUeZkXXWw1Iq9
pR7KGHClK/glZyGINYQ51suruEFhzn2krhZG8EfnpeuFgknaP0azFG1tdN+/S7pW
u0TxQRB931O5MN+2XtXWrLp9rl0QtLb3jFO1jxHy3vDk6Hd4VeVBtJbU1wO7EEmF
6mWfBz8uIM9la+xUeVzSFcSIcCLFDY9++GrBxaT1p1x65Hn/vcb2i4WmLHnP3Qzx
IOVNMktYs41xNiFY0xweR7eZz/vLyGITHFiMBRiZHv61Ml9XdFDquZIr1LAsqB5y
vMYA5j4CMxcaBMBS1eqCV5lPi1os98Sda2FiKGLxV01ElRC5GQ6+XH/bhMyx+eV7
ffhv5/xCKspzi9avz0qKezP8Y6aztkfa0dwZWPIX8CNxaB+dmyx+Tjp9I17jxLLi
w75eneTKAf1z1gIfAnfPRKDkTY3wBsbP9iH/+KQ7A0BwtbSbFfvfZ5nfL0Iuu7Pv
ZSUzGZTrNgstq7bQnD4ryXZNatwuF8kdiskvbIs6FsbAL8RBbDKANOc8fG5TzWql
N64ge+dgte463UFuyAEmrUfRTZ26HySolGs3bXaoyIrAhdnyaeqdj9E03ws4TVtK
0I6Wd0401aJkrYZTU4ERzVY+XtP/O4d8IPFw1vHBRuFJz/CXnk5MRhjwSPvnNNAV
7J4X7RlTWTlXEYXN1xlNTqnB+lfPjPUx1dluyFxiQeXFhrbIrrcWQINHHJEDBbAX
leiQsAw4lK5IhK3AClqx4nnyjZqI/T56tAzIIIWcacuBX8KkMl+EZLAVOkqe4iFe
5cQ+7LHvNw7LnH0t/fSsflzoEWeVZv1JpgGNYorH1a+UorKW4c7cB6QexGQpTRf6
ek1ndyQvKJIrrw5F7pOHf5tcH3RUKwWGIsFxKIuDxyFeNnPkLYqTkRslRhShi3nC
zZbaoBMEBQVcXdA+24aJn5KEnf+YorWH3Yi78ey5X1TD1a/FurLFGb5WWW6Hhb0N
jiEZcIukSkGYvDkbCCXE1H8o1+nuQTVBMaXDYWAQuD7dHnw3eo89x5wlkzfG0ygo
bOKgTXBqEI1kKW5ZyEb9SKz29g7uznwrq9HQSeCIIrjhHB+nTlB2mO1LDkceTACJ
mCoiC9/CVdNEfFZxsm1EHVE20gtDaj31PXEieagibmS2EYZ/aJr0cJ2i3mf5CIOC
ygnEA2LbNF2IoKeY8XxIrORKf4EebaQ9a4O0RjiwB/FK6/NDwZ7cLZH58dcNFO4j
hQrt4Ic76MMU454F5fviei/TytuHRE+TNPBZ2ALGiOKOoDsFOf2gIKDXjVsqoM2A
1PZyLcXbg5p6gU2e/tuon8eh4vaBjz0gxgBJQo3X41xhEqlk7iO9keHXuKXBsH9e
cJlVW7jaAKq3Qd+WfqetJyP9D9Uoh8oLu6OziR6D0WI6zXGlpev6hVW85cu5BAqc
gimFk4EoScnjsQdVS9no2Gv4pbp1D5NfI1cVdrbpiTWMXBbbMCCySu/EP30vtDpU
csPeTDzdEdqUZPnQEI+XZIOqjJRqFTP9XSgK9vM73ulBBAK1ZQ0gPXM7e9FvPhJy
91XGHPwRrtDm5edlB3q3fsJIMnNjOEZEDw6QWDuW6kRKQy4R+jRgZ0aOJeVJPrSZ
Wo8ZhBeejuBQAOWI123foyBMBPzAsGL2aCBxgop2mQiTC6zHFuTb+1qa7xXJ2Kck
fyXRTNcrCbe7KyppMne4LIe6uAeOU3aO5pJlet8F7etPtaSLcsn7BlfxbW+MDm+e
DOojdSxKOhXndkzm002P+us9t4zv4IFBZYc1wleUiGSsD0Oyr4cboY0URkuASlmL
z8JEACXr15lIY8vYreytQPuFDVjrdJ9oyjJdPC2u+EiR3pEb3v0PqhAR82r/t6OL
t3tv4wNnEmAMkHovFSc62Nzjuqgphs/nohMrR/ehK8iRKELqPKYprb70PzM+uE8O
WVsi2OCEQUB9TNC1gOPT7811Jol9mIisPab+2dYud1cpDF0Qo5ou2VYaK0pzghvp
qcCq0LKh9dVe5mI4mkCzXznnAGqbW2R8y4upsm6mGDjHQ0yovgUqnJ3/5c466uA6
ADUIhZI3IQlxhNyLGXMQm9lFmfXUCNYMd7sjULNR9GPhTB87a+ku4xO2YyYI8+qr
sq7bLIXZBgan3i5xRQADU8u8y6PCMnVfh3Ho0vxqFQ125tRKZqn5UZX9uzycKoRz
37d5CYwUNng1Iw7zoEpH07jooItiuVNkj+mDtouXLIMm8fdBz60x9lTRcqGaIyeD
KLbmXj0vJC+xaGSmGPE+hvFJcuVbZs/zVNPoBg1jWDYVDjNHOK/b1z+x1neixAmL
Rij56nZ3P8uRx3z7Bw54rzuvSQgB+GAjp3W4HxPoa/dazj8FNPtAIZHBGIVKEpxT
mKfjtv/u2r2OTwESZd6mSDfOMnKfVem5Z9CJRpbBtugR69H8dNrgOtFMyYCC+RTN
K/IB15W8crx/fsrfsn1ZLPj8LkLA8pg+JiDYUqTXh49JOvLJTH0OTQzBQK/HfZC5
nhnYFz5iWPLLGp3kiHfyWk9m8+kalQkIsyzLYC7iM3iQdm4Qwpg1zPd6C4yfqvNy
dgm9rfe0G7Z0+ixmfkTBvCBr/R08a86PJR4MJLHfbQoF2+dhplmTdEqp0/jm6aq1
t0P02qVd774KTbFKhmnlS8AXYfdt/KWg+oHl/ObQYlD7tVUsLRM+hzRI4lu3dhtd
a8QTH887Tzsk4grPTsM4sHDe8hCu9d5c4kQfxNeHYTJlJWeLpJYV0Kt4fhTGBCWm
nk178nd1SqYCPyDwWF1eisz+v1NVLuQKvvROEKqhs5IZEXq6mair57hBlplGbpog
5lPywEScRJMxwVY1QYLfxc2h1eO/u16Xi+E0EAsy9B17aAnm1FN+AjHP3IG35j6L
xPBjJewdy1IuhncLNmFaTXluxlZcPAObtjx+QBDEhXA8b9Pqr/i5hbaPx4lwr1BW
eQZBj7MUqVz2UPZlLv4s+rX2D45iGWWCDPbBUMAQ34JJ5YCyyPmIT/73A+CorBj0
aUSHCXtRagSJSLegrMCaraTmKs5C66cKbZIVrhj+mRjTx7zxcvZkEtQI44fUidZy
iAkXWcqM5P0oDJj3qgTwilSD70/8AI7Wsqox8AAOHyfxKy4wRbL4I1m/MJlGJhxA
4kxzoC4zj4MvLwYE+2On+QqO/X6Bo4yEn+El4UC+ex5Rh/T41qrRDEGoRpVJz2zg
8lZsm+HN/6xiuXHpfd88aoO2HY1sIZnLS/hLJauOvI1n+8q8gyBoYVNT6eUD/uky
PWJOsjQ7IuKbgxwvm84FArmWbtruWLqmFEMB8FEj1fP5OItH4GVmg/Zlt2OEu+Fy
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TE57uAUnGU8Nmex0vhsZmTXfQvOJ6Hrpfwo7Su3/M08V7e+v+4A3zY2q1zKYwqpl
vdXPLpsibyRNX72+f6jqGbV6LBgC9L0s5Y2TZZ7xJC+lfsvIHG6ADhuZNMLVarDh
Upfa8hrnoYnFiddFXnRw1t70UO23zr2/hcAnG029pxJclOi2SDfleLfKusb0Rxnl
jQ8yeADBsZTbfqcGjRynIzCOF243OqIWfa8N4XZSMJb15zHFdSuSgLdIIvSfEWDQ
d3rdxl8VjeTtKQUVrWsSGo/sTYfQztWO2tdzjEpfsOWeK6+M78rJPx9u8DccmtX1
qFUKvp5BYxDuYl/e6ogf9w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 21648 )
`pragma protect data_block
JGanKDhyh7CeGNbXeM2Dk4vuOoZGFJVbBezidqVpQvMBlvuvGFbEuTCs54e3C7ul
AFB5YLKpyxuP8kUqN3kilnowJPAWkTDMYLN0f2PYsSjIXI2fgxMHZAH1e/+gmnQo
PJKHfQtRQt20MQVppC/SMuBdtawvGvCwIMiJ0ULx579JHXqJWXZyn3eGd8dP9i4l
WCArjAcd56WTDNajHrmHJdtoL9d7gge9MwyVqlDfcho9b1/di2vvIdrNkLx4S48S
86MSsiYjdRLiwvP/Utb2+AyZ12koEunEnwrCgCz2aA1WlmUEXs9xr0HL8zgYcbpv
z/ZynAcAe+mScqvB+sImtWbpubQA2WY+KyVoTU02hTYwBvNst+K0KNTiomQecP0P
YqolUHVuvkHEUvPHpAb6Q00dK+3moblC6Xe9CLHlJs347sKqstCVuVhqk9Aeqx2R
2I9PIPKdy6CwtwjIKJ/h/QWfbu9LX49ZLWWvk4QVrpbPRjccuFYxut2fzWXwz6L7
KNtwtaL3ncOlC+Et9Ge91JQnepfapn+SNRzFHOq4E4Z4yScZWSN9KdTqtq0CzIUX
sIuoBtM9gHFpmbCLpzNPy2FlDJ5SCXWuRejdvd8UCIoBlB9bn3kvigH4B0/VYeAJ
Okc+1zat0opUHF3u6BoOc7GRHXeAEFiIWirUqzDuw5cSJe6MKN3VIDaVFczbxhP+
TMsVFCPhxUj05qtiBV/FJQ07yvR2YDrIzZmbdLmBJzIQOa0FVoJ8gv5L2sVyj6Lu
EyMyw+3njVhD7BLaxOJ8lvmKjrgIzUEPrUDMDhQtvbn6WOix/k0Dg3YZkut/xo2E
90/DISdiabtPIa6VqsWgL2cfOc2CKM9uUDQ8Fn8eZwWw3R24jwKT8TRPntTRxZXB
SxVzOnZLT4G45JwoR5BteMaFzSSIx5hldNLx7LJLzU7UGyvaV600dhZZmzDyMgA+
Fv/8mGrQz0ZoPBP27jkL2VtQKb8WUvCj21xwUh7Qk07WZRSOBJu+RLq9tU4S7SNi
KwMkFfdFsFsxvCHSG1X5ANMdua/K0mf1ZmDG2baL4YoccX39XzsL5LyqIVsQiM8N
a0SBiYOK87fY1hOtW0wQZgnFOEQMJj8HKJI9G5MfRpuIFpJ+0hKtmCXTV09sBKRv
fRCRXeZuWGdwLRREup9WRAu016scLTvEaPLg0Br+gh4CbB1zKSSJrnu2uq7d+EOs
rtYBMyKPm6tLJmO6Y5HqI3oidLBKEfIhalOG3lE6JOtp6WgPG1zXJpzOKirEWGeV
GySmZbfLAJ/U98A4XDmtW5CNyJY5TTRbjgFyNGHiBk+skWaTowCEmDXO3bDNYyxG
8MSVxeZizrWE29uxIm0k090PcHSNhHDE4jU2gSSSgOKdVIXfBxnvEm3AHZJqSULg
UL+nEwEoIaqYvBAvyYTw7Lgu5MOz9LzJHvLqIOwXlrOQvwKY1B4N8DySyT/xdne8
cRG602LKt5PxFSrt8F+3loPjqQDc7ZcrDclpxgz032otZrRnh3bNV45gWwzubcEu
f+mJuh/PZXqaqTQ1LyW2vmYmaVZubuFpbSt5W02eT2Ib8qTaNA4MpT88sGSEGSLq
vCcfbPffgtPkMaFmNFCQwYTuXe74AnPXGw6YAAGzYYgc595/LXbfXZaxDDmHIveu
x958/s86J7qtRIT6HQqR+5hebzDMPZUR+FMufQodrRToJLCr5kcqEgPnKTaoYwtx
Cl6HbPM/Pw+tiWpvwHiUG5U5Aj0rwMFOZDyyhUtbQb5mqridpxVzooO3wgVT1DMI
FP1tBGcR2juH0quXEJhvBTAmu7uqdL4u/caHOieqCD7rKJODLbHpdqOlPWlQ+sMR
dXxWB8m5ipAT0EwKVrWixTXa1oxcu66RrTLOfSmT8dVwCKRromKFF5CuMB6Clrys
w3guXxnbjvQ30nYiaFwpLruF1rHTuXRdhf9um67vWWwTBn4m/JyMcvQFvWMdYzFB
fsbzsYceejY/+COCRfSfgce5y78ZL7ficEmlTW51ESgEKfnBl+6JVIjysO8vpMkM
n1R6tF7VSWQHxgX5NTUR90Z7gApbDpVwQFHIP9QmUbLySGopMZUDhMwDqBJSutlB
2HL1OAw0mwzvVNy+qMy5ddCltACLxAxkiMnwVOdKShYaHGnP/qT5F6VtVzJ5nOeY
Znda4gUi9zjs2RvAt8KO6rMr4WH4l86wFOmoNctRmVwXu+5YoLkYcLmL4NUKsbAi
+ExpA4yznmMDdw0Q8G8usyYUapCTFWYQC6pKcoei3BePtfTcDEXLeNec6Ju6cWAS
CKVTo+bgzyprIweMgOd+sDLPxCOP5X/nJt4IuhVxw1p33hWeTl4WcJUuERExivd2
mKweKozTr7iWJcLBnRUDNTcZBHRkYZLSPUMuhfmHkKuvDxPW4bVpRHnLd179p7vb
Ow3WWy9Nosl7DDZt0yVcXFX/k8LoOJVBhJkMV3DA7tKKcC3S3DvWlDID94N0GDbE
faUspHg6dmC22f60sPWU8fqdxxySwFpCS6TtRw7MoHORDh/0EeQgtsWK/AlLZsr7
LiJ4doZ0DPkjmRmOu4L/TQzkhuBWRCBYczaDBJ4IsrOsIloVLi/KU5gmUg83QiN2
stJ4emaiiPnx0ws6bDzH9R20cdMY3DaASRXzaHQFJGRgq0T6s+du6IeXjvgp+BAu
UNoMlAk2+AFZ2JDrG5CIOARcWYfYdBP994rjXEmOo8a+RlXEs/1eSLdPq3mP/M7o
KhDKeLu8sfQC8mqTbVxQ7bEY2IMmwqYA1MsJMGbDZKcHnE40nPiP01a/UVxY9nF0
p4HvaI/FYRQQ3/gqf+4wubTQ6gpkQUhirZFKkfbGPeD54YovV3nry8miRaTYKEto
p3SXApEWLzbm94rIqpVygqy4if1bRK7owcr7fzFxpyFigB7LTTOXnMgCJhWG6Viu
eBC8mqHMlM29kb8WmxSnsdHBohbMlOTp8z/dPKezZ+t+S72kSk+5lcE0fL/tijOl
T6f9DRK4odnNo6UK6iQK2Ud2qaLhuvRcVUVe3fRBrnfCn2OuhdNIWOOCraFE24at
/n4/cPQScKbGswHup00B2Qyi1w2cslwBbwFFNGz8I797R2+ZUQE3ODPXAl+XSJZZ
lucaSdbcdLiEVZWUrFHqQCZ2supaZ5aqJoc9db3MeujAhMbxsvPgjtCpj0JfqEit
2KN8/WMvmU9lW9x6QV68rrwiq0CJ+3thn50ODmklsEDzZ+uTqWxdhkldmU8z5x4E
ssNArd/deeAUWpJikoqmKxvXc/40ByTMBG6Owkxno7jTLn1HGcFukV8ehV1JyykZ
Ot4QhxoXR4e0yVO1Kwc741E/41ln5c+vNWZN6WmjiGlVKfpqsx3u0bEq12BR9EdP
0hop9gEw0KfXpeFcKTyw3cfB/Of6a8rzw4z/Ifi6aNLIDhLzuVhkfEKqewHrMBLy
8PIXSIxtPXq9MAZQ3py75RTpeexF0WmDKYYsz/5p5RgL6Vq1A8UEbIMkwcrBuglA
TR6G2e3odoz6mGZkpzuzvhzQyjecpWj62Fn/pCx58oTxaIHyZSYUUwFupm0E9NCI
tBH4MRMMdfI/CrJdxpvSggRKWjYbuSkP07wUNy758iBgFl2sd5q+mFy1IW6L/03N
54spWrPf/g+7wl06avB/1etFaWXHnKjZqbdZnC3bxS+rk2df3DP6GaeW4nJM/LmS
ERFgPVsij91b6ZO2k/fkbS0N1HCdNMWScb+kplF0IYT+6EezkOD86VAatTpAPYuC
oQi4NojzGXi8TwNVgj4HkqCfVJ4F5Dcp0vbU9/pfh6C+dtZ5n4RYtb7CDc/KMqZH
XHeaU27B5Cll3uBkZP2C1f4gWS1sNSjRaYcwHuT/lbDFLAXi8pO+0pZe1T/sbK8W
oYn1f/zKx/igVtIyYYLJfnaYbsD6QWlGszx5x5H/Ktk6DCqKczZmpxmBzaBCGtVI
VluU+mIbUhg5At02R1Ulu/ufzil8N80H6MZXkaMMrLR4nNCob/GxRPlkxGjfR4KS
64Pe+4AvtZ9MS9v8AzvFRW/NkNyT3ie41+GXyc4+yWWr4NhJHwPCawFz8pG9goLP
GvV7PtZVbIHNOMavOq3A+UQXF769onSIPiIZMCHpbHLTrFfJgvE4uc5941NFbfas
zmdhy3WZw12N50sFVdM8VHQWy1eWqHMVzl9Q1VFu6IqtMExeSDmE2OAIgJ4Dggmt
4JGUlDDPZvKwTj6rWyWszR+3MOWqI2nTrkr5CEtk/I2ZunnFBcRyDioSEfI7RnfW
bq50kbuOihjBW0MrlpSfQieFJKbXMoeTMocXVc7zUN+f2d2fWdVMT5J5UUjuGXPm
2ixOhWP1el60ACu9Su6xG0P2JuV67w/B8msSXaQXk1igpkPWIBtCaMuLYV3vtDuu
xA257Vt8jfsdMvnO8PyjnwwTlwdczipCfLdg5+feKyp8TO8VbwkHTTekKQ2eWhI+
95PAbaVtTnNC+A2q+5vGCwXNGDFBCQjAjlTSKmF8P9Ni1bWlVQcRFYsHkbp755IX
ArqoQNMqahlHPpByB8evYiIeKesccys0Q5RU5Kxe9QWQVpFx05bkSjgC9+eeHHn/
6rUGRUmt6dO3hz7BJzjdv/pKXvsXO3c39RCJbADTG++tB0lBEr8Mp/bkhF2SmE5l
8qAjW7q1suhT37OMORMDcO8HQP7e7kxFi0Lf5e7RROjVI8iFiMfsS0+sYnkKyBXA
+5LIQdtoHY2mdmnRDd27ECSJtCaykse/O97QFcuIWZEddNaHolZg+csa32q3e0rO
1ALg5eEgMJzfAU/zVhlva7g+f5tCNe6CeVO07n+Uwcfxgrthjzr+gjX4wseEGvhv
EyOYRoqZKd+h+Y+EMZ6B9iW+4Pp5ODkKCD/loDfyz6YSvkJYgpGMPZKM1ugtHPl7
cVT3mtrQcGatlnMbDUmu7fLAtVb2136W35jwLLYxOZP8vHZidzORFgJj/6Km/pnP
ISZzG9tx854ODa3BocqzeV/cxUti6LAfuuDE/LegnN6kPLqy/Qt9Waq6Nxmfx8sS
smvseGmg4L1+cNqRQ8TS7RMcURAvp8GBpKYvDWJWhD9hAp+/lwGg7M/yMmTpLO8Q
n+igvUWFxerB/rA2si0yPhPlMjO6Bdyl3GiAAcAHGukdANhI2HC7rSi2ZEsQDcCX
0l8E/1lO8MijdKA3r7vKnJsIlNOJ58PiUaiN4aYB8XnTO71YEoJJ1m3nrbzemnDo
HVpzlpslaYabNpZ4fegmwyQMPwz+BsD0p7Gzf35SXoJ9ePiFHkXeBZmU77WlQ1Dy
JpzGhdrU6GctVVl7aI1lFMRh8y6NjK0pOD0sxfChysi14fy7h4q2OOsSD30Q5uB/
/z/9cK1P1+kzNnyBcyDFdiufVCi8MqCJzIu/o8Xgkmb2jiXU/2ALoLPu0E4ICpwG
kJz0uJMkaEWPFU16TVu0i5xmEAyTemc/XW0gFD1L9WQmduMvT/2Cv6DzJ6MwcWGZ
TPNqWSOFEOH8ZlbJedARx7zEO3ZOVnheY9aBiyAkFNycOs3A+BUsZW+/WaH6pzI2
3ID95sDsBPoBpsLQ6k90xqdxOhaepIMcj4weM+zbRDzlOCrjZHIXgaKx9O4P395q
gr1sr9eN1DdMMxZGhPk1EIYbD5WNyQmEyWCKSwMQ9hMt3k/JMrDbwvVdap/4ACFh
uYoRZEvHRt2Io6zAdyvfu37kktDdzTCipHkEYLwZ6ps4fVWEHgd8AVp7y1lnlCvk
OWweU40fhgclqc301UjC7uPEcu3VaiMifTngQn3b6LBB7GIsDRcmQelxycMLt9ai
9+dpz7FzpWQ+NPZ4OH/Uyk23B1n43LR8FqVje/dHEcxAmV96tO4MEUHUlMFm+q1L
RdcB3D2HpgfgBL5qaasfSSou7um0HQQdjeyM0llwahNev7i7rGwU3wiNfy3RRyUD
npvNs+8hcKk9rF4ey+LCA9+8nlI75v5tO0xykfobQJS1IN2ERQCKTOJrFzJs/lHx
YlucVpERsc06SbcEQs4hW2m+gi7af0F7ce/e0H/F4rnaeWkMZiIoU7NiYe2oH7V0
f1a2vSt6uzAjYdc2ePvVXrjGrSwl9Gqh7K4gUKMZ/QowiSfmT0KxXdV5MpsADbDX
paJ6zepeOToFRxcLC7P1AYqxikeXLCprcJDYY4gyQtBphgnhv07Il2BbsH5iklkq
b7BzIFBVCZ99LuC+luY/ZFLVHMQSGvIYjq3dbaATOWt3DbVb1fuMi+1jkT5tgkfn
QrUS/N6MFT4oiMPRCU6YI6yAHQeft8pg8DrjOsaJ/gQw0aUqJEa/cgRTM/agIPg1
bQ0ZT8GNtgiNUi/4x8IsZ4BYaDQkmeb3LZG5IQ6kbDO9IOQwjLxejemoPtTg2Ypx
eulokZB4dbzxBbOKWzPw7hJwXcun3D9vpPU2Mp68DhRYeOQKHOLvj08FlqIs/RHO
7Im/yZ6b7eO/BnRgQzO0rNkIxevR1Ttj/vtG+aj9H4xViU78sIX0Xgf5sNYciO2B
D0564SfljqK8ATnmNIk5kxgCK5DuGGOUKnmqGTFvChUY5XPh9Cu6MRjtOqd81vK3
LqExxwBozGulArbO/sIiS+PFk4/R6vv3AiBk+qSvI0Y4AhJxWqEFAJZLO0SrYy/l
MIAt+TzduwNRXpJ1P/G1LLcpGqgq3Fd9c/9QZwkD5P0Q/EWFjF9Zn99mbSZGCFl6
26WhvqUv+ta8v3JVJlEn5atSFlZ9fHKvhoz9xS7CBBfzsTEkvzZ7rbgpL4O20eHD
M8BFsulaw7JsjzPCkke1fhwPcWbr+HcAstJEnUjHj1pMeI5T5dtTsVnP5B21OPL0
2xvr200ggPD3dDwgbomkYLrcAnKS4yXg4heCKw6SzevXH8TjeRPU4HLpZ7J/6lmj
Ssi8ojqKe8UGaX1JL/SaoAhSu19SHu8/GTTl+tGczgxLQ1NEviCei/EKWN/k+kr8
44nMOPovKaEDm+4Iwt5jj3Oq1CkiqpsPRt5fmXr593mgt5FGbrSRUzOCX/KrwgyS
gk/lRUjtte3J2cpQkaO7btsfEYye+FV+GrB66DpzEuu3LHWFBI6P5K2JI+feZjLA
kq0exETayumsu9olSPpw6foDsTwPCzw+6eeqzqGY+nqYBcetxXUCZqrdI8yig1r1
RtkZHedBVJLdnlUfOGh5liCnqvOaYPVKqJoKUCWOzMLAqOJ68SP8c6HaLSbBHk9o
aFhAd0ADC8fw8rTXysiHbLDqw4MKGaFxlVeV8+nSJzTSWMpyUcY3hRdTc+Gi+CO+
9qY91bHRCYKOYT+mdGuTqW4GHYcdvl/aKFnC1tmRjTnEjYTy+tjbSvCobnZXMz/L
njDjTJjbjx5UbigL1FkYT+HBEmx4bXQQjvqgxx8labD55KEZ7gsqX8IaByMi1DxB
yKyidWLakiK5YsgSuCMf48g0M+SmVSbEiZsoq1or/iQSlUGIqDIk45CNEEsaHetM
dSwpavnYOY20CuFMvPB8LRAmUVdjVwFZKWW0Gob/DJhntwSix8aPE1pQ3q8NjfCs
FVfO2FlyKYCo6OYRUC6evREyr4OD0X63LdyKfDaO9RgKioTTJD3tuCOpysxBC4Ws
nwMasZgwyWJRJedaG5xqMw0Xeb0nOF+hnALbqc6blDQtewjuN/hnBMpyt01QdFDp
s9UGn3N7AGM/B6TE1/H9jw5H5QSRjlBkMtgTj41dnfmygjmUB+RJyRCQSDpZIE5V
4u1pRFVQVho+F/mXvQtWW6Mw4qqpBzfHA3LNVv8yGQnFr11CKYSNsDUJySWNR90v
czKXIyLQWXL+TWtVjCzOHdAehVn2B7oDSC3nudSu+uIOceTwgwDmUGv//xMekd0J
02ssfWaVnieg4HwuE+SbaJtX05rHHERBtcco/7aL6aYJHMO9rWrWlvTitdzXJr+m
wzBw/C3dNK+0l2k7By5ANzlXm1Zwpu2hdm7yxPhtKXewLwLoBaiIyIDXNNf5aC6q
KkjqW+jlmWD83BrCO1GwmbBggz/svxm05XD1ki788VxOYym8FDiyqX9HxjVC8NOd
Q92LiCDk3fKeslS3d+i9/GP3qSc60PsvE9cXu2FMuuuPkyY3Rz3YpNxllzS4WAUS
r7dSBb+9JDshahmjvcioRDkm9CoyZjx6FZnSrSp5CG1AQ57lYDe1/G4BJetsLjoP
b0hdPGxQ5LUpdGZ+5Egi65dmcf3SH1TpykAL2Oa3zLdLfj7dVnZ0QX4WZDaH+JvK
9kej1jFPGoFIUQmhp/Zri+FCMJFssmmf/wz8ek9Y7afS0rAMwBl62XR/cEXA9xRY
+WKaEfJoiWqojHAA0flLPUs3IJTIeb1v+48lUdyVRVqJ5/XaaO4Cw5wEZl+J5nJ3
lFu+bcZlLu2YQ8zo2JHpHcjueAMUNNW2jkjMR2F0kZXbnr8TmpnDjTynfpvGDBZM
EUd0e/nRHDQP4C9VitTn4gRF6WdPrNxyI8uwwszWLIwJoVOMZeP/6BSvYj1Ik4D0
PUrwOtY6CdSJyRfNJWWK0SOWft6XWnoVI+DAl7x1BQ2ni9/hIgiVb6e6gm5P7tP4
M059nTrWPkyStAXKDccRF2pAQ38jucyIrngQ/izAwtmN39Kw7n99zMn3LdAx6cLx
5ClBbc5r0+ch3kK0CusEXYcAuWq/p1SJNEJv9I+jMdPiTZoxfd0LXpPmD5bk8zia
eVRPlSB/eUosMsG3yAIp8mki7QV6GCIOl4tNvfJoY6jhUqJ5rQrzoMPVALSpqBRb
R2eECzhMYN5vi7JoFk4XXc7b4LukZXN7CuRsCjWiOt6dhptTOzv4A4PNHbym/WVE
yyaXuQZGaMhpYtBWJWK3/t/IniGbnB0agsyaF6DlwOEVT0getZ+SklNxdKhdtefg
AFFABYpoLwWEX5KzsrfnEH6g/6bnuAxj3lbKKJRa5Ilz0pVIAel3Ds0wR5tj2uIn
67y8IZgMh2gVgEl7SmsAwEtBed4mVDVzhv1p3coj2EAhmIpU1Qp3BGQdpssJGSaJ
jc6sUz9qiqvJaXDAsFdOY5WU/PuhidLUc3/W3/D2pn8/oXdjFl0l6spm2Z4CK+C9
FCDfL92s+F9Z+xkbjCHqUp/f+KLtUej2EL3Nc8XtB7k66F4AlOXvCSCL+nAbE1ae
UrC1O2KlZhXZ+CxcD1w79i0uJ7Tibv+waQKW+xQJS3eLH2WdLVSGGVniB/fUJuLO
ZTnW+oK8VDiuKLEHrvybZNe2jJ9YeyigbcmKUwnugXaqS+I933qv9szuN5qL6uHJ
ce1APsikVLrXXFsmsTeysJ380NeSksb+sA1NIwoRyE15p7p5hZ8TmmDgFU6CEiKU
V164GDlarMw/KOD+Vpfr0wTvF2fMXQVbXWM32ItTDc6rsyJ2n3iJ78rBIep8PkTQ
+uTIHgt9+nkrBoGAoPsLdXg4qgVK//sEsLMS/SiM9K4kk7RRAFtDA9LRwWcdxeNE
v9Mpy52lZTLJobjB57HVengi5RBb5U6gc1mADaj9C5Y49HvpRoqUu2tyy0TyP0vP
EsPNG8Z3m28ep29tayuLpTJWtbk/xi2iDlvvWY90xb9pia+E89h2vJZ0ZP90M6pt
uJi6WgqqNDWBDFfXNcQuRvd/vjw+QxKd+pL3tpf0NYsp6gWdbr3ZwM9HJgQgHpew
iYnVEuFu5NP4mapCmYtdVVNlf7mkl4YKoEmYifUpdNAFiiv4z6a5OF/dJTamU+1F
Fn2OHqUkSOgRgQ7VBE9nKIPclPo2wiM1kSc+hwbslK+eV4lklAaOrcNIxsyYvqoo
DrQTlQWJj3cd5g1uOHuQKbcHQY3LuJgRlIWDEtQki6fsAmVgpLcXvFOdDxpbCaNo
olSzIFmkJJ51I5jHFKpjhywnabfncJMYu7FJZSYz0bhUSMtsXsziheMyGUGNKgPU
j8tFH4rDlpmzRpaEiNnAuCrePA/nlAGhxuokUe2DIuWXFKDu4XMV4vKHTg2iSocD
3B4VKtKoEkTe0jTcqYS87iCO/LepJLe5/iwr1xoXr85WxYuuQrNxp+1DwTvqOvK6
dqitjw0BoRZqlTcJFRhjPkNMJWJF1vYgoabFPS/lBQ7QGx+N8Y7uFGa9sd8lslse
WxDYJZkmb3hhVFYS+VnRFq1ZUwgXxL6tv5c9JVTcRfICWgcz50PtUPVlVf9wGyPA
nX6xUxT8EFnwDui31Bz6VymoC9vX2L/grNyu5sbV1cazWs9WfXL3BKzqoDShSpvs
j0IMHO+yeI32QIoV4CFBuBhMngYIHIuuAVGjNFlZbSKsC4j6iwH2PKw/dLDzgf0a
jrfxnMuO8YCPK7/wDj1OZ0JhHIMsDEZO0Gpf0mjbtTS0ZveOz598sdAQBeRWbACz
fS6SVlvFIc7VI+wl04zahiRkMF6Cebh8rMEN+4ahRFPJ5pITeZC5ENrFc+sCZ3sU
mvySQdROEEBttPy5sSHDWq2/EJDWd5+PcCiJW0QhYNK2HE7YS1EqxoYlWKEpMiGu
Rjg8gbxkjosvaueZ680baGtRhbP6hQQ4cPloNqcNgihQ7s/jDMDZ2ISX6+oAifCk
KK5z7WS6CmudrTgMEkZv3UqrhxgoH25gQsjxLV2Y4o7UK9+mgAWdlRZrM76gg6LY
42Ni6cIdrVlKwdE98MNjnnbxQwWC95ekgjDRbF+/TZlhR44okXuXPHUYbCkUL9fk
yyYSqgIfJCI50HgBeARx6Pe/9nduFNJN/0F90Vk1VV4wf5ML8+FRJV1AxjgfdylK
9qGaFVRHVTGIywbpmVXG5asy6dwhRmPP7EL86cTZpito+ongBZ2D/lnCPUkiJGkh
FPFtF7oOfoe/5gVBEhR98oVzg8Aqa4u98pfOCCa6mQVwXuy5nDn2PvEF79rqpfKt
aYXXHpsV5BuDFhDIdAvL3iSWb9yabLhmqiYSdqgK7QLCKHV3Ze2eyDwLBA7q4NoA
cpXAub4MA7I5FmqedntO7WhyVc6gORt3azT8Zc2Qj79Z6xfUIwBqx9Gfa6IcIj71
y1WfaMWaTSNKBqjCC+NfNehzPiNAFc9SWn4Qj6JvBk5VBcfm2unG1d0C0rC/jxjT
mD0k/bWWou9l23s0OtOYXO3ffV3pi+D9lszADKjQoH4yiEBhXnrV59ULaqC378S0
pPWvpKAP2LsoLN6tMKAQlXxeRFNo5ewm4vk1ZQXSzAmhT3ghFEbu0ZhUxm0KB4zn
XgA7nc5m8whTEwkDyay0r8NRyHVUyRlQhPaiaK91EEiRq2ElJHtNOlPZZkGxqsYF
yV0WC+HfyAAeT8msvBUsf+gi6p8JP2VqJ3U1OmaBmJOjSA5YoszQ6V2xC3Kkba6B
ChgRXsR2sNn9ix7Y3TC6L9yMV5SCTOeh6FZo2yf8Xhbe2wdZRMDmeVTBlvvmLvZo
Lvl9LZGbUMU922X37kC6R+yiec2d/ZhqGIpYnDJFuWr//p7cvbJIacrMg6Z7R6DG
NC1KVIVcnCguj+Nsdp7GUw7lKhVtLuhXhL9hYZ7um7AWbsQ0ZDrfVEZdbrWh4/PO
RVOx/s8ah3hC4dpjOFnSh+Q3YUCbstOy0sg2Te4Xl4D/MJ1Jiu+pFTc7QeJaVtB4
kNGR86jyGDCt770lMrn7b+xQXd4j6v7CYosFxyoebJG1vaNbMMVJNid+x692n4jo
IGYQPZemHKbTQRWbI2mbbztIKBMF+iGInEXqaODKDIA9tQZrkZbtL8VbBpfiHvOx
x8dJ1ZwH2O2DDkskhe+gePYkQZdwrDUEdDB2WOhOlKcx4KKL7DrDi3xcQmGx9PTR
RZocYwrnXBAOymoATlWOdrP5xQbPaQgb4ZBUZo76dRMgFzPayE6lmOHeRPvaBUPi
CqELQGER83HHxpBOckwx/yu9EQPNkcuKWIHOegVvN08CXVCrufU6GoFmlmdNmNM9
SQoFtMRd9IFCljcPtjvJb330C2n0uX4aB8Pwifq+8oiH8vAnN/2edqpF8RY/IhBW
PLSm5v9K7cYtvKYo6Scqc6v3IfNrXqvamzYYLLXA1tdwEZ3W4Yc6xqZmZBLfh9y+
JFopVHd5RqhrqbW51cF/qScrd9gkQ5mejisBVT0cEeEZmG885JUZIQ5vcVMGfmN0
yoR8dE6jytvnB56UFtkbKb7kGPGoqDDKGW2AdcYUsvdqI3fOoKf02u5s35KIHnIh
CDvb3su8qbpjjLwejSgTuFQ5/cPJwL3ZCPsn0ECKzwoGiiV8e4vw8TM4qElp8M2h
vNsJFMY9x2gzuaGFqwcg5zhZ9QyQyrS09mYwcehq/Q1jHzRV9TuoSATNsZo1qqsh
gyfkCpX8Ts2JS0ERqmWLVWvXcJSTDHp1bnfVQAIbVTdHiq1fcWl2N7fX7T8jelFQ
bK6h+5N889jw7VrZ+ZtyufIHAS7khUpg5HitIOhvH8obmalQSo44jfFyFilOe0nN
cPALJR7LGX33vvK+CxKujwwAu7FB6+TbsIVJpo84b+m3jAl/nWD9RA+GOatvmyho
IZ5bqye1X6rx65rAznrLwJYJAR6tbYuM1KZFFYpPO6a2oO8cqP9CkyGCMaR9OH7R
BQHiTkQ0CdTBxt3SllwGsFWWhCWh3HbUpqyWaRkVHvjMjofKEPeY0CyzrO8iRNyG
Rhphu6I0VguQ73xAUzRwx+5BGv/f9Io/HBItB18x44Awk3zfv7VjZ17KX0NLCxgq
tO0NeRV/4ASorCCNni8JM8Tc+Z7so/lfFe2lwkhKp83UUBQP/2lWC7Ez5GhH5I/M
+FeH04EjND9A4sJm8KRUKb2QWnuGKxeHzE0KiI4dPrNQusIdWTHWPdrq3vquWzjf
N7bzQDCVVTduJaw7DDLsIPqLqoSfm/UpdPq8SPgV5KKRagJl0EsylvL1jDIHx45k
8LnFDT2hLc7eUjZy+m2WiJJPk96z3znYlyxGuERMvFpM8TsknTySMw+Pb20rxD7C
p/pYCldqmUO4JcaeDo5SLjZsvxwQVN6J69CA6KTr4m02OZrqzQwVccNZomnv6tLW
t8wr6teEmGI71tDKUbVTAPNiWwrPc4Vq1GGyUIIRJ2W2OnHVRDNH9V3KQcnGn0vq
uEbBoDYTNO3VSXRFLF4AWwW/t4rHaWtIyj4J68YR4LOQkfU/jNQqU+9CrGZs1+s2
cw4Ur6596iP2JHQSuVqAr5moTlwBmtKxXCbAiGkIuGcILZpP4seCFsNDip52qPLw
DZiY0gQakGxo/BUdXvEJYU7YjcziN6uXgnbnkPb2zTI4Jreock+1u3e36srmMW+x
5ANYUuJnT2GAbBUWOwIhqiIIAB4YwvJaF7yI7OlBDXuzgB/ckR35Or08svveA9R/
zEbJFyeuf5Mosu+uGtDou5dzJMNcX+SAacZ3C6plQMGbYkEADLblSIQQHBL5fKZB
yyHtSWQ3SefyCmYl8ArmxXto0SV00Ai/YWujH7hY4Nal6dls8QvySR8QsZvDRiKQ
rCA50T+ZdBZgOwMU1T0Y0veRY5+xRpXNVKZwNOVZqWk59Wn8vSVN+UNCg/xAKMBZ
ccyJRBdpVvfhJBUG3Q8+uwAx49tJWy7ELWwu/TxQZaOQZOxowceT5I85q4intWeo
vGZt8CXReKLBZARxejpp656hs5pLWvofbi1HeR12qqnZsLhkvBAEsa62ZX+voDzM
N0N8MpbRV/UICwFzhTO+jMbUVcnCY9u0tiVUPZTVRKTdGUC/CQZxSotGMTOg6xij
tpY/GpqwRYeiOH12haClpc7ihtyIAGFW043Zp8vNgen2AbGoJuvREeFxysGSkMdm
1x7oXxEImnfifURi259Hjud0k6+9M6w7xG5AmRzAC8rkUTyUUOW47TO0IIroNcs2
S+xcXvAh3PeqbFrwBP+ls1mswwxu/bsDuL8zcrhcXMynxyVej2ElXASaFDZJ+IOF
63TbSPlfQgfnQ0qYu7DrJFWnrBG99kBm1HwcDHaq7sGkaj8is2n8vZ99lc/2ptrl
U0WNPO5jmjFL/DKSIMIcw8Qy1wSPCsh2GCLdBDbzytjxLONTKEb/VcZEwXUq+hAT
IBAr2SVrtgsesks2vug1AujUZ46tuDqRgAhZG+bDBnMfFWUXmOBKi5g5vpmWviGk
W8wbtXYcpzF0tyouqTa6uDS1ko+MRyCOaDe5mFpsBEusO2yIU453z4baXAnIIfJc
lDnHbbdtqdvW9eDccnOrT+IBtU8chhoATydZ659XB1bMfBBsk1KhPHF0GWMTrYI6
/oJjgsLQqKsE8VtVV8cAqME5Jc2iASRh4xg1vlh4FF9PBGgY96La1DWpZtq4IWoy
EFFEqB/OpZacaE8KZu/xO19bw2ZUMzQCYmGoXQW+riygwUQygfPQJ2rRivi4iocE
1hmLqIjgvXIXnSSDvV2IzO2Y7J8LbpmMM1kNs/OA+Dl3QnGN4T//S8AqAK2MKzyG
VIaorP4ip5ZXUDtFR49ZWxMzoptUWdep2m1hAhMmZeEKoEXzvwPSQnzF+wJWvtqM
3PR5XlQgQjMOvX4nfphewVVdOrSjDeut/25NOjFtYFxbxsRt8Qd/rfPCle5itwhU
DqHozNMwIg84+7AkpGXtpw233w6o4DZo/e2OtXRG+c+AjD7QQ3OSsqHBRcw3/W5+
rmSPd4o2xf5hidTftKIESfYVxNIChKkMi/vd7r7ZNPkKOqdigvul7VD5kx9nUYdt
sSSdMc1f2IFm5xOcZyY+3YHaSUd/Mdl8oXbMg2UgnZmiJWO6GznFDz3Ku3nTvIEa
e38GiJ8Kw4dWPaknrFPd8P9XjaD4htIFd2HOhOVUPm23vt8E6HDU1xD/FBIkT+gJ
Zms2YbNLfP45ULoPi1XW5w9+6+juvZL30LXnl9U5SzI0MBJlwc3puLrom1K1i/J9
Y48dTVHXtX7V+NsvWPduT8RzhLyczEXOWaAR+MKgDJOZ27LDik79//y3CqX3mWCp
o3EPfxUESk4ca46Tr/39Lcr45WtgcSx1Ssi0TkuI0VbATMH/GUUg8ZjlqhlKKU8L
KodtPlYgg64WvrD/4BMA/u4G8B1oHBT4wACcEJwgh7SJXt9Uc/Z7N3M4TbmG6ubv
1HmXI7tEC7vu0x2SEX97N4/NVSI5RnYwcAjFWb1pWPFAIIbI/flDqFEP6Z5TM2xm
DPSpNVNDId9Sz7BnhwjEmhOj1aoP/QbjADSn1GujruGk01f36ZyLvGEXcvpX7S0P
vR0HHm6ErVAQBR21YzspvAOR8AMA7hMa4KBpUmwtiZmsfsSPNG3Aq+l2PMIJSAfc
D1WE5WHmNzG8vriVUsppcZj5BgJZ4sip5oM+Lr9UpKotWmINUDW41ts1fPHBd/Xm
Lg0zsvDIu/J6QqXOsE+wNYLomNk9FuVqtSAUcWFGI4Aq15ivmD/b6DMkFffhhQnH
u2oFI65YZTE2iU9A7MBbMYSqLJSWxGF3UP2GyRkUhDoNAkv0lN8Ze7LQMAYHb7x8
BQ0pNHygFTFXacKiRm1lB9+ZDmVao9ZXUZMuk5AGw5PN3eM5m3VXxd9u5jV5NlGL
Ek4YX/Ry2B3UgY0YtD89haElJiXmr12VVh1QPnw77kNM5jMcNJSzfrto98VnOYyP
5zL+Z3dLTZm+VDAAq9516sK+7508CZdThncHXB4SqKAGItwhPI5CdbEPyDpo0CCB
sOkrpWKto5uJKehBmM+1rtIHKqA9LqjRDx2664Wh/oLcAsrhO2KJLYMjTQAASD1P
Kn36Noq+7unCPxzfx3Nes1DufNg8bBebbEYbQizp6UirbrJry47uNK5RzqDo/hyF
NAKTB5kKUkETiMGh581gse2vFfiYA20SAwvFBSf26fsn0COBAJgJMdlEyxMsXGw+
6d7MJqGjGyXZQ5JMonyqf7BtiNBBLeBZFbmtS64saqpYy9TzVu06rDA5GfZUgLD0
rrlSKhBPD7U5nyKWfqxImvKMqCCFqGW6RX6mi+btqc2cCX5I8FGne1ZuLQiN0x/u
5koOxI8beu2skGOl+WIRQH/17iQCU6KB+6wFAF30KBr230RXcvGAePlkaaH8sw3W
nVbche4B/Y9++F5WNEWCzJK8FGDy3oqLjk0DDteac0icIx9urnRhveXypOeUaEfR
0uTcdrNIooOYH/1oU2WQaShnQCp35Y/D7UQqVqEaXPVvCk7iUxmFgNkAiYQtsFTd
PRIKWMOyGmAerxrcDRfOYFV50avPmPt9c5j1XmuIhKA0UhU72XzoL0bogIp3fRCp
jzOjOOTzlD1ebvQHEohyHwPwa/YP+WTerF3Ui9UmuMrfEc3R8nylQmezVjRz+qFW
DrYqPJvasfs97kEyjxp5JzzsF3LarwC3mJAuc0DZm7MKiIMz6iipPAz4DizVlCxe
E8Cxi4KsGUrsK7tRt1/t2JAb+d3kUw9zWKKna/8n13vWiVJX2uquiISFxAbx/kyK
SIEch7+NoqFhPf3dMT+7deigkQXHgpgygpo5AVDFRuBkxlWQliJFXHE9EW8cCY3a
xDMo+bfOgG/CnHadWlxv514deZ8w/j3Gr01jkPCWC4vxw7xACLqjlNmFeXiGHCUp
LX4iCiEhxau0q9LYyS7Gt2rJMEwmyWNNQ5tH4cXn3Lym+JBKYwYZaIKDQlSzcnLk
FvDanKdHTWjE8jIvLWfqghLtevtC8Hgps9nxztFVxira9bhZAxu+UcYWZEvoV4Ho
ivN94y6JkkfhURfURAFSmIiP9CoUc68Lwdygv0TnGNFR2OWN2BuIhQrmEseMz77x
z9UKAdsXOUfepOYATAtnfkv/sjIVpspQnSeJPGfmT+0Oz077HDuns6UtgIVlu18w
a/NUT+BKCVbOTNz64SsAL1/YdcOw2kX0h+jGijfxQP2j5NJPWCnW2n4Gf11X8yZ+
y2gmn+geFQvAJh+oVMVsPjRmsN64EODrr2adwkh0VTKACCAvihFBD+IC/FyjtcYQ
K1Eoo+iw41i0nr+iax5+ccG/5prgM07KCvMbemYqUGPqS5lG/Yw2FdvuGsAx9kkT
Bwjvonyqwbuy/GvWHSeaZp7Zs3CQ9e+v/wbXBGoVgnTjMHhkeM3GkhRWrRIpdlbz
bo36Njq1DA8iSg0wU2Bm27ADHoRaQo6R+CmL1MUPnaRVIywGgWRkGibWQuRGNoI7
t0wy274DNEtXT7iGUSJqnEDojGUyCz8QbGoSXpngq1K0Pk/sZiAbCvAQbs3fsUdw
Ey48NU5cX/R1x7rbx9kAy167R1UbC0xISIlHFcXnbnl5XsJWp3SYDUh01m/agFvo
Dh3HldUFecxQZQAIPlipr0oEeHCUu/UrDcyfI46b+dpAIZt99xoUkT/IgnN1eP2+
k9GPHKoy0tS4xqFe0XMDhznL8NvsaBNUpYcdswALOUss64h9wEhn4bNBV4fmJXvf
fLqonytK9ry1YdOx6o0k7Rcf4Q8rFNlE5zvGsLLthubCv+jvR+mvCz/4epkoE3Aj
/MABnF/ufdy0X6QpXxKgLMtowkvPU+WMSIjlzduR43YDJI1Si+K2oqbupdH21G78
vbmq2Z7/9sKVaM1JS/rEDhzAipb/UBcjYvIwFY/IkTdopeXRCT81EAXyT9uDYFnD
2qTjyDYQkH1X9cO6CQxWqa6MPwRD/f+coBPLWjrH9mramccLfPEn3T+4hMkq67g1
kDvov4ugXftGNTK8p+30jJ1wEndxhAYK8/DwPOoChX06XVfkhEcgPsuXFxZFDAA1
CPMTIW9NXcNmMlD7kfGSE27GCJJII8EbyNN6gTeqp1qycLaRsHseUnM9fn1lGEQC
ob60YNTOd9FelsbdD7Ap7n+AwHcD4PS5gGg78BL3Avco4PBRcuJPCv0LvAv/k54F
7cZozIgUa6kru+RdJPKFEGG55MoHCX+nU3bUlm8OmWTJIsQWB+PDAvB+3hpc/KZg
35gS+OvkOHSpNR4lQxZF/y9cnDcWrqCYu4yYTQKZtWqXtvhCZM3SkDMtGj0B9OUN
Cb1x2emLUGeccHLkN97HuJxQ/AKkMzx87/NORh8+FMv8075MWa+8J8WoIHwhMaiE
SKt43cMNKh2wHk0Td6A1WhLN5ZxDmR/CGrrnvlnyRau+sBaCCie71RH16noZ9mgY
6pQSQ+sya3dHmUOuYjed/1r7YKKDx5zRfs0xelgj1/8bMHHpRya7ReDajqz0ozjO
fzi/nOlfy8s3A8fL926YSsNMUoT2Z4H2CL0GGWwC7TttbFgqzjX/6Qtaw5EG8nPS
W8KSbRaKBO+SWLlIncbaOQ1GkPV4YV6TKikuj68IasTYNj0FQzAPdzaNuYiT5tLy
9Sz1Eh49ks5qlv8nbb/86t+KvjPYcrtncdcGKblYlWwCnEZ8ngrIrF2blhcYrKHN
BwdaIDFKNeG55Q4mACuGKlinMXAoVr0UlYlmj/OkgvR1Ea/X6FE47sA5YT4OBTXw
pCX3b8SMr7BAeW5LQ9DkJZznqUqV6cqA9RtEGicVq4j2KXOyQpEnnbqtuJwJ7aTF
kZzMi7PFIFd52vraKpXj9oYEYtj4nCRYNIDVCmvuPCcmfgQYdHsTMEFaUtE5BIVQ
eB9hq++JsGmHzgxIv8BRsxdnfkcuWFpeSqnnpwGpZDxSjN1mQoul4FjMKNmXC3yq
ETqndlerq31fqH3sR079BvEXNw1wYv2piEABwOwl/qLZZ25cxyp1Rzqzx42JrJ4K
tIy2XRG+MQB+l1cQiUA91ssACgxps0Ne5+I/uVXXPxjYBBLPXk3Cc6UUKRYHuhWP
LzfBFdPacnDYxTpXqeV9Z2Bt3w9TIOyJlRD/pkNlvlaRp1c4DVguaTmDiOlHLwKA
ytTG+S4PKlXpc6br80VCtV98JyTLy8pF55tnHf9yS7UawQVHZQaAtdx5J/oTVx+6
KwRC+bYI+wG/wUZEtc8sCLSEnVUP5guDgKm/OhQVNab8QM8ifP+lJP6FaIAzlhs2
+e32xn4S3D+7++gjDVfzD5BjIE/JImJGytrijQEiDmTmKTz0UldUVmGa22fSnT+x
KLmdBFSZ8kS5LjpJQcwFaGG2WCGnLZ7UxeiYb4zO1ptxPM/ZTm1EaQT8/tTM9KAz
saT86FLp64bgDAmgEZ5K9I4oD7YRs4hw69f1tWb1ab3nNV7rIfi+OcwwKUF8DEFb
JX6T0gvlGl573Dmuufg5BpQG3OK3XLUJaH0gUHeccINi2UbjwKZZIbqvqfw3219L
LY6K0RAS42Wzxs2eF/ojpM27ZJf4nvRNJfS1Hi7yIs6pVXqkrCg4KXnIsbo6wrw9
FjiVvMJDI5KnodrF0K51qakCMnD66hv6M38a8iueq4a7Vmkhlx4DyXNbPgO9Wsoe
Xlg8GNjfov5HldBM6qwaRUg3fVObOtr59TqQVgKSZhleypMTihN4y9M/9AkpX8/v
YCr1oPs05k/qOVg4UJ9bbxZTf6I4nkrX/+d1zcHsxRxkjThBnJ+0f34q8H6vIjud
sVnJTNyKQIkojS56RsHCOJEPLk0pfI9rLBs3juMNZJpIFIDIPQcppwIRdoP+7mdM
fHB886e482+Uevy7OPawRgSVpu7Jyb61lIctlTbboJCyEn8cGA4CD2dhW8NVc/Au
KgBYPvm1WVnQaxaYMgEKI+PYEcLRZzc/4pW94/NQrBWJ7xLK4Q84JC1Zq2Zn5lL4
uR+F2P+cOQXf0W6m7SBPk9Lh0NQe+ZqKB91dhqwT6HTLivbnj3G/QndrVxAwJvi0
/8tn0gIHzpCb1y+ME9+QRs8zRe4EGugQvivfU3Goh7boIw48SGidWgaP4SAT+AMO
hq4ndF+YKZYzHbLrgYa8m4oVNVhY+9KJlhDjqss9cOcVxGZlI0qehmy2xxErYJoY
JGR7WteAz0e8lEp1/41cWYU5hZVk01O5tnUJTKjhJVw3/YhtpTpr4p6Sy/Q3I6hN
IM57uPRfKJCbdIxlFauPut72ThN0bLBNbXChOGN5v1/F1bS9EYwoV0a1zSVFUe9t
IKYQzsVOvOhPpkoAhs3GW17WdJj7IcH2Xu2M8TwsUalIHeMRs6br9Ve9DULE68VH
JFlqrdmHXm2b+QO+CTRS89pWuIz3xCTejf3m+xvKR4pJ9rLE78X2AAmkpJUNTD//
1zsi7MZHSHg3IFw5ia802FEvGnKzAq13o39+WJje0m0b1vdC3V/Oco/OQt5UkToE
39p91zLeIzlFzFV0GSdNZKaZhAv/iwUY0EwL1wZEYccOWdSm83zRyK2jO+A7Znfl
uvPIjmQJ9swkvBeFboQJmIIeSSYKp8Mkzin2vdspmQvx9xjj87p2haP+2wGn4FL/
R/PZfDZLK/bBmmNPUmddL4tzLMwdsgwi0fsOiiQEfE6WIKe8LTkzRhtRP8M7dBn7
6HA+Ek7Oie/vkWGWiClEiHzeD1ho8CMTNf1MySCgjOMreRk+P9GIsFYuTitPqJMs
mAtiwSZX17j+4jDwGZCCyi4P8YVvp1rt+hydZX01+OyOuS/vz++Vxy8VtXyWMtnq
1thZEOAAmBCAFwh4MVzAlrSI0X7Vfh33RVPqFXce0SFAh8X2MsCnXxvbWTBq/olR
KYTR51hmXcg+RDOxtrt6vAzLILr5UCps4HIPghxX49lm/N/ZHKBeiMQQC8Z96ad3
4dn9l4cHIkDWw9sk9M69zsJKGXgceHP6ZX2Rvo78ABG9Mv3r6ADIAI4ry9IwnLjV
wR2SKczkZyxpMujveMjdnys9mhRnNhem+ovEs1Xpm5AQ4SCWMXKime6zVK7TVSvN
QLgnRVG9r081VQo4v0k0dgt1SI3QWoUpf+mXz0cLBUAYTtPTnE9ZFnITxD3U0LIV
TqtXD/PVeUQ//7rWbfLEimQAnMNWyUU74WcvY2DsTF/S1eCSagfHKMdekMyqzMsB
uZDXDbKJaNT8C6aUslh0wcgg9GRmOrjS93YBvOcNgPKeYEim5JqTWLSrPnarFzaq
VCjeI2m1d0WLBwyfved/3uy8jtx+AOw2o7mk8GJHLo7EcqE8SAW2qjcYqJEvgLX6
SbwPHKKlwLzYxwnsHA05gPKHHwGoqpjI9PpAkzyj245l0WT6JSirCmbuagEFW52P
j/TjswyMiW6zzJrgM5EkNMZodRwD7OCu8guS4ycKR87qdEmW9cZQ2evzAPPpgLC2
M+hgoJAnJtaWdX61ogDhpUXgBxBFDdSymIpzBjVpsrdJsjSpWRyebidZlYXa8BGO
+p3OmRha8+2Kz4d/gexSfjyuBdmeUxxUSwxxl2PjYwVbG/Ap1HarXu55U3xqeiGM
/cKoUC9kAd/yPMh1VMh4kBeCM4qNCrIriTyqtAErwStUcZ2VGXFCVjQr3WvzoFD0
0PlVlYtJMV+/cwuFN5ypj3U/lIC9+DF2xvdQrk/upBTCW3tglVRo7BDVqJtmBqdi
4YQvYVE3B8BJr+UFsAyrW2cachUHyLt/djDkmc+kNq1Eh83G0ZdMfyUculii8mYu
a3eezDQo751wb42TnDhqhCr9WVsq2tMbWK2tnyMt3+TMExLgDVM8b6HCtM43Mb2/
OZlqZgFewuB2ocnUU5qEKDFiCOwugW1NjyliUItJlGbj5JfJvjXD1z6gxx8uxewQ
JvKy//ldi96vWLF3ZyBNc9JK0w9dAuxXK8Gt/awXW8q8mq2bn1/i4XpSjNdKDHA5
0Ya1Qpw2gvDKGqXDdBxP+InTJJuJ+mNUnSXZy6iYjZ5szVjc+XdzlLeZMBMc9QW4
940+UaV0t7xI5avbAKKDx2CMLqJnVc7M5J6jzZcDVPNqHLLGFrQ7Kse+J0mSIY37
OuYzDrpAJ60MbCyBw+Pqk4WyqG4GDhj3l0kKbkkksNIcuUJV524RrmGmGnAMuOcH
EIX3B8RYF8v4suQpTygehbmu+jbg68nsfbag0Uop5uuWgfrOe5xFYpK7Bl7TKXQx
ePr1HeHsaS+6Mz9viFkCHlWgslpAF60VTnxOxpbP2pXg+f0ClccUszBthyG+7th2
dFW4Yb85mHB0VXdPnwwwmzISqvgGN6jqdwZFokr4YIy8FHRlGkG5ocJ0PlqQuLhA
g0XDre8TODsmGxBMEEgu97h6UKiF+oBfXCJwCrMD7/92oSVlmQydNYLeqPbDmJwX
Rs77bz/0P6HtKw4xn/WtmtV5sCTNLf2zfQYKsbKpejbv3bm5eXkEQc5wi1rY+lOB
dg0nW0Rjle8+eKWc07nOKoo+B/yZQHpn8tj1MWDt6qdykKqcYZ1/VgckyLCAQSat
ZBbepKiUfXG1WnAO2OWWp9DaR3rl/6oMDS5jV5TJw1WuUx6rl7XyrodLY/qzYFIi
1BuBQOjVtMpGwFEf123EPZpmxuYQuGtrNNs3T/1feLfuAQAOpdEXgNsJNvSlCZrR
D1ERzhhARTLkuzE7wgGcU/haJCyXWCYteWiwPTpBSqyyzUw3CfL0IhgwRBR1vRMT
G5P6uEQBn589hyhopNhm3g4uk4zcNtoNRKK6YFLvKXLA/opfnCE8uOJqZwGBp8f8
iP4qpu+v03h129tXEU3niqONJ621X95KB6VtTKAQE6vychGg762I9mWw7oHzzjTV
9vSEVC/pvxuAiqH3pPkYhDrcJMOzjJjRNieo8qehoMoI5t5Ej5D+ggmENwaRGN6Y
lWkybRgCcfDsgbfpLK4fTUinVUfiJsKlwB/5Bc2qkQgSPeK6shEmBU4v2lenD1z9
Zn0bT049vfsskuVaCMiwSk1pkja6paWw63UI0S+Krf+xYv4/hEWmxPpxgw4I4d5W
NRIKoK8EWCsw29hf3H0PF/8TokIio0Qw3V7h8IhGSrmkzR078rR5ZChDOk0pXZs5
G+zZBHnCb8p9lwXHDAZ9nfkESymWhQ+wDtooRkTXbZp9XECanO8npg9AQ+HH/JXr
7bjfZUpLcQ/3VrwMwcpQu51o1SXhlNERXgXAAcERi7tEKNt9etWe84W/fcZsmVNZ
oz+7d3qdBMrt921eTnqevUsOGWfLHVTnjnDQCrgsmnY7G4nGgETC3/ZMZxV4o+L3
ygQqeuvbuBAvLgIBYichvipMn84wl4azjszM5EIn9UBjiCoYjpe/NIqqw6WqZgkF
atkFz7/eEpuHcgMbTpMlG7TQcadLAaMaUoNqqqT4GPRzgnbrVd1/632Bp/kMljDX
IXwbkuMm7vJ4LSu1Z0rGkXNQn1SjtsJTiZFgsBlgdUtKRBh4XmYLEO0Sz+kwCHIv
4OttSGZl74SgRzjKs3brgvooiFtHa6kF07vAMWDdvR94D3Z8N7WRYMGpahI6A4NU
Wfs5jdDsaDWr8dLumIII5cY4U4S/CilBcNBzDhX2wBTt3D8ZoVJDf2Iijv3faSHb
NxcrLobzHlgsJVTiWG7rHyZhYso/wdJRjRT5ZN49jFjFWfbPT2HG1sIpjBFzoSa2
MCRJFzJdgi2Kt11VJfJfXrfj1GpdsYWqc/D+Jmzi9OPqQ9SeUn8kKqpGwVPNfeK3
ekZHWOhdeR4DV9GOjWu/nd8PkfTCTO/DZPMuOWuUefQ0eRef0N/uI4IoiXEcUu6i
1Twp6CDYsLWVCabxe72hg0gMiP8x54cBgKb8gwnoEoDVulZtTWR44+0NnsjoroPo
RUwtWDIgZS4aCzP0BF3ymwQOWUCgpfRIQSxDhSColC60twNg15O+jRbXgbCgK2i6
zpa45FufJXmWL3fkFyk3OBHltWe96j/uLtf9I5D30xvaBslw0XLdS7Qq50it1Q8V
rKS8JzAcIh+I3RifMWE0+RUYsTZaoXpHGZu0KwtEKlTvXqjA3I90qs0Ep8Z3AV8v
GBldIRkNb3aU/Ipc7+pH62QGrtT+OEF+/yzsFQCJr7z8ktXpfme8CoXcSBaIJgij
fKenVIuJsvP89yCyhaG5EUIL/KBW4Yz+Slj4wMlv28gDur/jWZEOVeu3ZhBTC/ri
bOFhm7mtCim4vl2N/aQh9DqdqHjiP3W1T0FD4BhE7vE0X2ewM1SgGqI5jPe4zTrY
+lOt7mRMvcLlllcW5RglMzwkW+sqt1gr6V4y+NcdyrPa+YHD25SWMG7jfJvHG0xA
Ev8pK5rjDo6Uk91RwnFmrhvBxCsZWHhdpj/73fqs/+9v3SlX4ZyArOmK39a7c1VR
5xQ686Qbf2CYmAdqVKL/Xj7UOcttWUNjXWQr93+v0MgWM6SA0vufG2jCC+UkHCdQ
0CnFpEidZkzWm6KYIpwNVhUazn/u12CHZglzGU7ozbDOkptRJ1xCqt8pYMruIpzL
21N3kwTqrxvaTEmOk8N/ADW+e644jJq54E7gPn1D7IMrwWA9bGsxHJidx9RO6BKW
tMjFGojSZYjaWpLaBQOC9uLLSVBWTzTIKsQl45BqCxmc5rgosXd1ScAOErkGEd9N
XNvZCbfWLm3g7KfymlNnqEETPHx1/y8cLrPdHAj2wvSJA+Z/7LsLwSelbvtN9j60
74AMA7kVUxhXs5rQuW/5VbeJD1BdlrBbN2JEg/Tfc6aOh1f+IdcedBL7B/UH46eH
P1m3hScaEttOVKeoIexqLWL+16LPdO4m62S+YgmIiLHLImhMhAFz7Atv3WSqJEJX
+/sBR4pnA/P1QLYykXE9pW4QFZudKw9oSloGom/mtGkkN3nnslEYCv8lEY+aHwpI
c7QTyxgWCqF+GSNCGfEUj8q7ENRz+pvtHsk6dQHuCMIwlo8RwoA9ixsrvYz7wND1
wjdiP4rmQphSnXh9iH8836wqLkxMxQY2v3ziOvFqw+xydUR6SZJpyvqOXVyFfFgK
tsauK4beK1O9ia4V2QWdvX9ZNQ/eTj1uuHMx4550wvZC0ZEIJDtqeAhC2n6TCJG/
CRoeHxwsgolDKlFEBekAq/ShChW3Ab/RADkO7pyiiCbcojxv8F/YHr/Uce2VSC1Z
DgXcB9lsDXe7ZyXpKWnNTxTCSSTzDg8OA0i9FaEFXnfldAg49g1jEB99z0cjC+qf
Zj94XZLww56KfBJ9a6ipdFhrWDa7oNy5EsO17e0q2XO62o8IjZIy1RB87gevN/HP
ErdRLDTnt+jxdwplyrWbuZBjHo4aK1l3+l19MoB6D2wJcjCnr9GmQeVEzY40hIn4
yOrX2oCdwjqYX/Lw3pciJYU26ls8sutNu1/HgEaBuk1cANr8Mx5vMsaLsuM99VcZ
pHV30if6IFqmxYP5hbI6kRYyoVu9q0KCcBJhwnC8UgTcIqwE7h9sS+1EXc/PaKx7
VUyF99XQZtdpSgZBFdw0qtz+9v2vBMW+P+ilQr/5vFN4045jM40Pki2PyBoDudoh
X/L8pd3gtsJhbI85Qn3pP1QdG92rZOBmyG2xu8DX1LMPO30XEaqFtJEsf9DqdlQ+
QyAwr2PMY6f1q0oLhTHxPQeELC98L/AXs9IwZwcmJumdCuXkbEA/IES9Bk01SQDm
OC0RuoTeGr/f+a2hN+PHV2+gncei/9rlLFRf2PolEXVAHSw4LZ1drVTdKEBvDfXX
GQ4kzkcW9U4hyxc4DqhpkyObg2Rw6VTf7WCZAORLnk4mbe78z33vikOW6PB6Qdoe
U8ANLdgmhjJAp00OJ1we53s32AbvriYLE4jgBuguu+/Zu4Q9DF8KCB8VeSBhHtfI
cWTuBN6iNcvNNnioOqVBTYRXLMRhW16wAVeapWmscgYQfSkz3ja/MP2aY6xoklmN
kesFVfgqaMICMlJW4+nXqpar02CcPRVc6b4ORNTLqbkLju7CMNLB0VWuYuquDOK2
4uVwZ6/kdjcqHnRGmHE6NcORBsBNsM/gdRwM6ufsLb0pCBbz2n5B9kygXMVPiDIp
R6KQYd6OWZgMEoaX72j9pyQq13XI+ec/nDCgUzFYuEGp/yE+z24wKymTOophGeh9
35bpHGNECDee0cbSfBOPTxkeUWNS01qFpm42/l+voVTdhadTI5+7yB2OjyhLf042
0p7BXZfKmUhOZehowREr2250ep9yRYCjTfPtwhvtuTIOzu7CBhdDzJkqAgo5fj25
gM07enK48CRS/PC/hwZ9OcgajjCBdRlZvDIYoylAFlYon/Del1VF1grunkFZv+qj
a6ciJdOFXvvLCjnrXA6IrWXiICUIYGxGS8+Decx93aV95vvJn+heQkFjhiopGaQ2
7SI9U6uptMsKvHBStZ0qR+iYw+B8kqa168IoiR8vdDmC8HZKo6gAvv0nekzw+3PZ
vLyC8mzYC8XGJO9NQKSk5IhtxveUhMIqRG1CnXbKIUq5AFDBbvruwEmXehvsrx3a
Muq3J/9dhGamWoh0bLaEylQ8xDk9D4pGIyPpm/QEh1eSX5MgRti0ZS4gNSIwqpla
8pu8vDqj9ocNCxlvBAzc3Ng+1mjzrAVi/BmR6YC+5w2UTJQgHqU/lw5Dydlaz2cL
oRWYC44QxAlgnTAm1NQ47xStB10QwERBoiZgYykh4Dd6rgV3BvBzqTYnGvTlSmVp
w0xc9Ew1q6fNAH7SMgGXndV1Ck+8wrK0yFm7iDB590gKNColylGWxjpv/v46sTQ0
CTPaMVghdGHzGtX57UXMAyShlCXG1pOfL2ZZURSnBJpqBbVC0gsZ+nllvftbXA3N
f/Ijs9hXVtnTXRX6TkfUvCsHhGB15yklf+LFDU6v89UIQdrGOwN2DMKNTinTOhdN
VcBZjU3Wc/PsFCE8bOyZbNWjmI8x1ByrUCRjEjN7gu7MOmL85XM+WQCcqvF5DUkz
rQ8LWhDMvr7izFLItJ4drucofylf1NXj5ijU0FLjOzIGtGS6zcQIECLqZsXU5aJ5
TKDSn/nNUw+N8c3Xxm6Gi2cxMRrNNbX0WIQdaXZrICaMBylU5PP336uZbxO8ZcUP
JZVFLQM53RHBT0tAgMdA+NSFYXiHvk8O0LqzT6KBgHhTsvIf1WEW3cd7SFJnQys9
p6iiHlVy5dh1JKkLn+XRxxt0dBe9dETqp4MTixNAR+gdM1a/hrfpQhWrtsboT17V
KVtqk6OTo1e9F/MaH841YRz1vIp7Pjx1VTI6hFDrwzOsckeZuG2wIZgdOY/lqaOB
/cBbleM0hviKoKj2jbrd8hi11XIeu5Vauz0rhBJ5LNluIwzKsygNyICPMgi3TFQV
MY3K7zSm1RDoifNwfemBGqke1CTe/W+CH+byeMXRdeED9GJMPdkuPEk5SlRK9Iar
OTuanV45dARspm2k9FukkbzMN2JEmyYzH00rA05Ksra3+E7LQBSO2U3PN/uH5rED
5Cf3nejwBpdNm/SbeRDWKNbL2u68DkzdwQ9kMkPtnOGVOMpAUIVmaYdax1RzZySC
umD4nr9VZeUmqCmXlcA8exM1l6VbWxyKPfJCE72wJQRKmp8FHBLQy0GMI9HHOPKL
Qa4KUmimj/yI5Iq089bLaGLEnJDPBYHjAJl0fRNd6QvHfx3GnlLTsjukCzvAIVCx
zal+UUKecqeGXewUmRS1lU8bUT81FwFwVsaivKERqimY/Vw+fgOHa1SgZZ4tJ4jt
0rOelrgKj+LAjI9PDWBfgFyYFTrcK1VDmeQW9Cs8mq8AWdUt00TF+L2IHMA5YVvy
N6+pS8uXKlhD6rLmv8FsMuavKGoSGC4GX28GbtAQieKQwqpydhBDiQ9sKuiQhRMh
GJEklL0HQBbmbLL8T8XxibICHTEZ+U3/J5nwAunmOCWiEiNdkxR/ldoXyjZGBa10
FVgy5qcPK5oGzNR7hFAzT7T6n3dDXvwXwf1RWz3S+JBqDMbfZkKgg1pScWqCvQLr
ybt/xnmcmmnP+lqIoeBGlw2VxZlW6x2usE/uMNkwP3KDmqLe2PE6/5QLhRMa/QaI
aVmfRdfVrwaONMEAcb2jPYfyFhTWC1/8fOFpDkY+l7VyaxWjynr4LXjQTB4EEVrT
WBfOs9p+gdgxOjPl9wIJNBdx2pzgVGGKkv4rlNzJeAz7YgrD9xX/6wumdZoPHVMo
1+ExmtOSsuHCp7zgekCEtrnyoksz80XdJ+kbjUZb6PgKfGlwG408T6nQ3iG6aBdG
f29GVZkNXMQhaeUBpRspGD+aRGGRi3Bly9P6Pz62vJjoCshJ+1SqbIPdlZ4z0VPi
uh4SOMYcWBtvUovhtJJSB6dU6KS4/A3len4r5wXPv//McGM69nBxwsjstdHGvvC7
ZenRVAqax5KecVpBcRfCLJueNbrBoAewsvWf1xiu3NL5JNfyXRekH8fh4bftkhOT
vMB1e4ToOfTu9Y6xsDPji65x729zKk0KQ6dSmboH/HLVb0qaC3irz6nHgYXSgSa5
gRJff6qES65RswdnsMiB4QeXNnnc3rNC2QgbwapWEDSW56uasUFA1GVNnXMRPg1M
zTGbtrqgObNKGRWZMrU3t7UaSHThkDnqbym/BSPR0GmSf0/9iNUhgQt2mRHm/viA
AFGuZBIEBgYcrmYRPf1t8pjRGJua/5IzwhdPQXftYLq5vAWTWg/oBxQm5SZwO5iK
nhXd225WHE8VXehFBnBDyd9xB7SnvH4aqKkEuhObcziSe8tFo3QTlynSzHAihkFr
RKm4UaiYWoIOTu5LrVNfp3LXp5uvfQNw4USC58hV8kNioGG69WPN0FhytINA+JER
FaxBsQgEzQqkZWWbY4Ivue0bKH34uMRiEeYoczY+2WwSoovm27pFCfApk+iVOsiR
2YgxfzTzoC/CB4blAs9xv0NFZLbjydf/bfE7A0T/cGey5IpQohJ/kC55LlafwEtr
AyuQ0K9CGE7diD1nKgtOTxy1sfq9Dx2urjPB48MTJbkY7TNJr2/ohoZyeq8+G9tg
BcIS/drcbbB8rNjCoz0QIlpfEgCYJIt0jLU9EkeBIUwYP+nnuNDWlXcdTgN0hbKB
yuaH1ebwuMzs4jQj1QgeeBpIK1yXwJ2oAAvMKxACR5us8seZPzhKZVRhALpoWwmy
q6ryqR8PoftJVSEivwFLDjTG6hW7MTzu2XSFSw/nlWwzwpfNowZTGgcQuVFvQiH3
UHRMO8D2w0D/02j+6lw+OJ/DXiCDaFnazKC4TlL9a1sqAfCmRlnuVetEfRPX4/YD
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ezbEJhVQmXlDkRGnJpOoNlcHZzZn1z0uzu41vDyirCe9Ks/mBKCk1DsMj4hPvhXL
55jm0POMPUNjLUUAVJFoXGHBX7kuYFlZ2GrPsuSZgiePqpkNSPNpjs/f70KEhBF6
TaDxr8pq2s4FdsHdo6h5DuoUdd6AWOUKkwHPEpjSR76zMB4a9D8/IdSQRgV8MohA
xNKgQiZx6PADli/gsGvFq7bN4/aXuq55Z1eoa2Q7YUJ0FtZ95Gx1Yk9DHKlu3Fcy
MRs73A7O6zQASzhbrrzWNXXXnN8EhL6SDXFtYQT9726yO0Qg5rQN4+PQ6HWwQDGp
aJdhM9hibsUdApUCgi8NAQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6496 )
`pragma protect data_block
A0clq0xm8AEmgaELhr4My0DkJb2TrXSy1IIQkbAjLL4KiQdmlyS2CIjSb0yh4nhi
d9nJBJEh35XtZWftUQCVjI2ZIGrE8KoSrWzyo8D/IIXV+jeeRqhW6oQ6VlE8DBeY
xH/IU6zKoutN8WVQnDC/Q2f68atdwyUe5dEJMbfp6OmDt36eTwGFf27UPZFSK8rZ
/QitAYyPVq/67TRRKrMx2HW8gCTW3ES5yfr6W1JaKCspmIFHj7MBlc8/GcKY2fUd
MzzARt7po5gcH4VpeI8sDlFkdvR7kl2lvpQmc/4Z2SAPUcKItbMflG/qFGeF5SD5
HSJhSzbAFdMit9O5CMO3FLpV2mfNvmzBFzbC/TrJbhj6oNqor8ZJIBhagX8MNK37
S2apBjUCXeYFy0LknSllDJ3EqlQAJiUj00QpX360M5Wag5Cvsjw+ZGmSuQxW0LEF
On17TKX4trWhlVqvUqEsEfHsDzmM/8sVJy7b8PexDcuvFQs5OKmSk9o9RE2chjbm
h4vCeD3QdSbBlM1qIcZXfE2pEvOiBdNawa5HY/Lv5Ps/j3UKqRC8sjrM1EWCay+S
FpViXNldLWawE7wyVrGE7HjWtHSmiv79izkzmpadW9JIb9uL7QocIOQH+9A+mwOr
OfGh5HQxGm7VRYHWAMxHcNTg9eGirIA7FsFrMXbxXlId5uQJgUpkSmYMmYMucWuB
oalai7b+PF/lgaEj1+HmLc0EEeVIYZqB5+OVCkRVypDbRRZTgLPbT9Kqo6lC4pzV
b3c3rvHmNytelg/To4FthHmN2UWRlVFEi2lyuM0jb0sTspifeSjrIHQSmVFcIT0m
mrnm11Eo2OsFzHHWC7Wj6USU/3fQuj7t/16DFvzZkfyetbW34FurPl5tmaezpKVd
tX908pPaTde3jejurkuq7L5dA1P2IQWNl6cJ69HGzYvZPklEwHH9t8To1lnZjXp7
ywMIu9Bc4+dcgTNiyNOidSz6c/6AmyqmM3l22xpFoEjsBCiOy0OPYtmvOdbtAY2C
MG0k+5Q2w4yULipG2n7DXmkFf1oyII8IXA/nGUt+JAV/EVEeEr1l7xmQ04HJtiXA
EysXfRA0lp6REGeJR3FVPjWSAAH+6Vh0HlRsHArmrg2KfSLKywnVPEvDQD3LO1L+
zwIPdik6119dNqN17W7Et0YnxX6USjEI4Ap2W5qCh6C8XBa3lJmYfHx5abJ+nCHr
nI7PiR64ao7brKw8uOtrBRxgS8yJBRYdZoGht5e3zknFzutoQjUbPi/LjNYAHXfP
Vq7agmLDsHjDiF7sc6K5YEsYmHoH7Rz4AjY4buFrQXirTA5YQGf9EsYi1zDGYYtk
RzXxdlG6Sn78Z81HIcEpDpBnkKpcQW4Jq05cW4F82dI/8cPFIFv4p6bN4Dyc6dOu
KS5Wo6oii/sAb0+OcuQql5G31VrtTNd0bPj5ZsoR3J+KIhGYQViTauvpDBdbx3+i
qkVLdcxz+sagV7B4cvtkyxxMrMQS1gAAsFzm0SaMjG+8CCSVyKLufcWkwWArgVhC
izPKeVFG4E7UvmlZPCnN7/CFrSYdXvjVczYxMQJYUHrBxkg2mBsf6L5EY5cPtZZq
wr/wUTxOUOQ19mO3/8+q4d0DLdZKwUB9jI6ODrcKvqv6iez3xKzPu4MwOpbwwy+p
sxg1xlnJAXHrTk3UTuRCuOuqM6hp2ZBVSDvcJnDDYzeLb8UILPjH0SnDEJaCWuhy
ctgN52+a3EAmFH+68M02Xi1flzyaRP8n376qpMKt2rDIMBmURgY9uPhrXQTeuB55
JLLp7cdFYAVYSTE3Z0j9wtafOUY4a6YvF27LQg7Ou24dPQqdVNvQkqxFAGXOly87
x9UK1R0npFHrX8qOxDvFwblmFREsVSoU/8KHhrK+2+ihgZLE1mFoLqo2SvFxmoJ8
hufnxHmu0g459o5a8SHRIvO5NLgF2oDzD1xy6gRIOEBjvCSidj73otiqiDf919wE
UB7kbwsiz3Cr3zB2gOMS7UZDva62+RWB4XH9UGHxtap8/X6FViIhsS1RCXhLuOKh
DPwvjD5g9Q0QPEoX7FWlJ6OSC3ai0lP5I87uv7zEmplBzymNsF1KYBGsBuqWQmL0
yOEq+XUaaPiYzCGUZ7qioGeGyrF+qmJidnUirwCYf51VAFIZZ4Pg4yFvK0rftv+N
zf4HN5+Iq7FmvNZLXJiqruqHvH6CqbKr7BfhivTdlqteVpJIA1PEsYrLD4RLzjjK
rwHa+Raks924l6rtjdFo9GYybXa1ER3KDJsUjGD5mDbL9nyqU68rRUG8rn2IHd5J
houAECkgUj6lciZdv4MQptDdnBldix6e6Jck8q5Aamgz2jTcKMkyyi1eCtA7YXBR
bvCPs6JZ1GMkFk1RpDvapBR8jEWPQ1YTeBDamC6Yb+ONK4y5CGBFAKO2090fDaE5
zHhFbcsWs/rejvHMivn/4nd7fHeApkZQeOunN2zbUstCzegHkHC6PEwj/XgLyNTH
xGo19brP8M8/53SqJ9VlD37w+JiBj7Qi/LaO+0z5jcexnkGiUj+JBzpe8dpU4wMH
WQSwwN8h8PgNPA4oXDy2YBpFHFP6/fbr16YwIQck5VECgGjZBQe2h99fS9TjnBTr
8sdN/9/MvX2ovi0LWHFGn/XMrhIHsWvR9wgjV951MdXpZZwrRGIrVJQ+gEtwul0c
ahU2KX2b7hoAgEbre9ePHPPfZnomE34z5imXFpuAy2tRZSOxkVdnmXbt0+Flk6ip
g/T/bn/7Mwnru3Z5W054tpNX4pTq9AZueAf0Xwm3WIMfqQEi3SiuGh8YtIcOqOlG
ghdqOLzDyBXETSY/XiFlEa92tnhDVfughR3PhLJjx9w4F/ET9YiXwUCUgHPJZ89f
Mj3D6kbcAl64POQT6nFsbxaTTXzT3yqVNl4wi1bQBdB5GM2ZGbOEJrls+dtTXu1C
xua7aLIFCnyGXwAnYwnKuooO7Wi4bHXGS+4VVEHjacFsvzdh51tlYzBqLIm2XfPm
+9i0s9h/d310v8YHaMUMjJXn8SPWaDurFJh9051sqHMDLm9rlp9WzWljYNKJDJ+f
JTCcPvILFk31f/zAYMN5jtEJkfUUMTJHv0/qvDWQ02wtmZON5XMj7EtYg951/Bkd
HvACC1zo408EOdvodJXj9L4tQZgRIWiG4jlOnpwZEyWp8kgpUcIaTc+T4rpnD76+
byY9IplK5qQqsbo+6+FwjoV98ciKoRWZj+Dz+0qOhgyg3db1+OxYHeuzPZcPVP67
YXQMbRU+/g89xFJgtey7mYJS6UeNt12wuO4RmQN12EwqR8qCFL8FjGlo0n2gjyRN
YK0HU/tNSdyuXHmpPuPsXOu25XUf5KxFGQtf4UemvU+S0aVWLJ9NW/r14rsevwfX
F1hCKi2NCqEfXTnEaiVQyVgjO11CCrVzt2ozBoiNjP7d2BVip22aSqS0r3m6Ep5b
WE/XP4f4ZzhE4mmomCXnymwhAHG3uJPqmjNFWUMakTOEh37Ad8j/AmTmBTPsNqkU
NTaRco5NysKxIEtgtgPc0lXpV2xKJm5zkTSQ0cS8/2XETVyrZeYDlBV04M82L1ov
OjY36Rj/qdyy2W3Nl6Z0x3qAbKUKPEJAmjYZCQhkfGkX114/HsFk8g3LfDAJt0BM
HHQF6cjh89GC2mXdQFhQ8HGDRDyC9cS0skUGXul+8tQj7ei74lHnPXZPmP9wvlUB
vLLCK6cAxJ8t2uw+Cx8zrL7ln5d0JjrqTGTi5IsK4SbFc5huXjsUOF2Ge7jhsTFN
6pA9lYdgJPtkASqUbO1qXfE9uCD6pNUeh173zVk6tb9n6l80zUjlPX6KMmqfO/I+
4++JyBUopqNCHEFGGK5F0o+8QGkRmCjqD8gnOnCuJ08J8BylP85CyUqYRAjsgTT6
Vx8PZxYA2Rx/6EoWP9jnX4nJKg3dve1ghoQ9FuZAotph/C1+j/zQ0Enszru4Wrm9
E+SkFZkBoubrc/wdk3LbzaPfsfmswHF8IPMibNqjUzjSpbhVn6RN62uNVot0Z8Rc
MEhazbvfhrESnLCpTrPR0h7TuIJsPbym0d1sPm3s54dq5uQ22jJbbu5Rjv3zfASN
gMSNsw4dqpV+xPhkeLTCKhfiM5wZ71GDWGIiY5Gca8LWZOppFpBNMEW/Ulan+Tof
7ZeO1lrexKcgIwkZuNveW52fjxzAstgstKXYRXuiirE1VpxNPjOM0an4iw5cbYVd
uMtdfKazKIqSv1UBHNYOKlV8B/i8tjg5x2pG25Rz/YmmxN2dQGgcfKu5BXj7d3Uf
v4IHGm0jxyfvJEhKM7JcpjlrdCx1uZi7ylIx96hTXjZ00hN0jO2ICPnSI6OJ/Akk
2Lliv0RbbrTkA2U7u/fKGlQMmW9euV5s8HDUTQbZlphHZ+2/HF69Tj1WhUkGm2GL
Ty2oebl9fJjtYb0Pu/CVeLLmiVlfcdX0Ov5ODBeYuqHeHNiZuwbSw8pN8NAaemrO
kr84CxlDaLJn+JynJrsmjmG38wtwSnKBF9eguGlYfZTpZA9tg5dYyW7hM6zi3RVc
5yEzjNCzMs6o9R1MDxPpElijCecb4kfcS9SamW+aTkyN1/RuMD9zKsPIG7oWP8zB
pEZHq4xpaNgn3lu1xkLmvigdOAnfiyI/BIS+/PvGEY1+bmDr5ErNhtInWEc4EOIW
piRHOOxPwelYZW9JwkaZnEHJhaiv8Gj4Ns1O2AvEIIOZ49NC7aDd4trE4p4B3znw
ztjMkpMLXMX+fZ3xbCNoIYxe5P6lD+UivFu1Qbgwzc+YT6CRWMlfIZJgWyK2pSs2
2vtsajIq2X4u1GBTRDsUWIXeH0DPbeCbT6ogFqMmV+xbwUtTnZEQdT31iNh4qKtM
LRaxRtLXygW6gzijwi1dIDAxoE2i+SI67gAbTP0SjOWvccmUZiMcsYjG9Jc9U/5o
ILCmMHVtr4xwgPUx8Fygzi+hTF7TeUgIYSjqScf+ybTEuoMUMibceO42P7kA1Np0
4pL+HmUwIS3qtbmrEc6b4Euzcfy24TAcMVYPNeD1S6MPS1I3mI4Rpgb9Ka+KdSOn
KCNk8zhcWuHsBgC5AmDvcc03Ygyzm8MRU96OnFK362GYHIgyVKeECvEFU3irwwFG
QtVe7noqUYw3AKjw+FW6ZniwhtOamzJNVwywo6CDJ2lmWunzVhXgKE84YUG71YDC
SxdVSwmgORukMP2WoJ8jVVtQvbyWGM7hmBINQqjVDrivyXslkoFCdPvWKK1VZaiW
ybdTqYqnRB+ikLa9u8kpG34dZpsLanuCsnZGnG6zoZG8lhL2VQuEbkNqN/COErhL
HmKNOb67wH2Urtm3IddmN9JoOBSWFWLPstqyf10s5a5lOqua+Exbag+lK3Pocjvb
tDz9ds35xktELPECCP52kmXIXSYUfe8hqp6D8j6NnOzmE7Ie553PnzPltEdHs0sC
17tDYvZ4shac1lzY58KMq381AkgiXJoO0iDD7jOIZMrPtPQXn57LAoAlpJ+M5EUV
E8k+eY/aaRB6qqfAr8y76yBrIkxR70HANB03Kq/EOq79XLhHsf9RSgaBNjENPDuI
2Sy+kthJfmZ7PrS1nMaz/kR+ZaqW8iPtpOgzf63eqN869uiRFdyvDQAW7A7ka1Wi
IEQy55Nm4f0uIDkotDyDCbwEFYXbopFAf4sHPMuAo1HVJfypWXELwYudQuqBHTc4
AyM80gTVhVpAcwLXDnnzzwcFD1m9BL+MSCHLYuECj5i22W1/0iCpih6tfrvkPvee
BTJ+1EJU/FsveAtPNFUF2MjH+yuSKIVlMAMVRpr2bwsik0TavwldPKRzlE6En/dr
0uhRzWRhfFtWe9Tyqk9xXh4TwwZToCxDmXEvdIZNUVKsZZp9wfTOuEqOK7WDc7Nk
h9rvVjAc6TS4SeZNb5qNSAvFl75G906re6lSV5gXxr30hFyFaixvQA087Gd4u94j
V7A/qV1dEw7wyRH0G9OGCKMeG/OKm7CZJM1IICVEh2bE690hrm68q0FMT4FxDNYI
5AeVTDXmR/jK+VgN+gynip8kOcv+hBDwL7Ov/SPtbFGUt58WDj3xmhDi2WiuTIg3
TiRBhf012/FvMmMFCfUVtSgwZpeu/AhZDEp9PNuODxbHJQfx8+k+iKWvAbksCgMX
6lrkerWcSjOrifWh7ZhuGnmYR0lPf1ZIXz4IHozbgfeeCr8RbjqbvC7q/FhwKzri
2iKgWaDwqHqDq6T9nU9MvcFpqH9qyxXpY95rvh36S6dxQbwee3WZH/YxPb0ZSVvA
OWHuUTmxzjrCxZMcEpQkoCWPUWBWr7L9XRE5yxcqZp8vlT5WpUeyg17L/XJKImz6
B22vPvKuW0DoqnaNgjm6zIxqhkSC5nAEeWutsX+6rK6YkBThCGNWTz9lnC8t4n2Z
qzB/bAM5XYVDS1jUb39a/8FjHi1GhQHuW9tJ89F1bdg8OlsnTz7Y/E0tpCT6bTHf
rmGpHIZG2phlhGxHyVZmzg5cYanAZBS/NV3GDSxGuOtvHPabPh6NsBFJbNDLPfs1
IGSkU+m8ONTNCYEH59rs9stKZ2JwL5Naf7rPHpMfpVTlJ3POq4HbIKOL929NUidv
vD5imtfAonjKrAJGhFc98Y9TgfC03BNuhHgyvAll67ByP54leEtBkkDubvWXM+nl
HFbqOBNxGER0TdOXSwCq63khqb3at1UoWutv0LdWteolOa/Jh3k2EcrZNYY6QNHQ
pWHbglGezmGK91NTuHQN6W9CN8PiSDBL00RIqvfUw1RHLfwpperuLRMBT6mvPU+4
QroXqbtQ+Rv3hAmDF1hkHPsf/zpx4xrE0PQs/2oOJr4kjiwy8ZYwQ4rMVOxtm8PZ
4P2MyfHU90OW2DgiL6ME3WHfPqcl0G/1vsEP/S+1vsRE5Pnw8PFTpWV8HxOyhBDl
rj55wphImQxJ41Dn6iFLTccBk5EuiUPSR5CkANP8sgl1WI0b4IzCXcsvMs0Me/om
oP/tVBa0lDlm1tlftdvUZ++7u76rUiZe5ltFTSOOvuSe/n7vg/MVzexSxgAZnBrI
Jk/1wBOjYoNfiXqdim8jE8UDGom6pveb/mzemJbDo4/rqvvybEeCBpbjTdZUJ6Ls
W0XcvdJIdG/0Hi/8kQGEMlnxQK9RNXe9DjA+ISmKK1T3r5ekQ/4B92w5q0w46jt8
3n3L913Ozt3Lwr+JJwpNVX1Ly6Quf5snx9ebadDgnEAbL+gAiQUB6p4YMFQs3iMk
I4Ywpa3uDTDeojZPfQsHaN8zWtwQMklfBUzSGcmNirrYg11Xmuh3+CF4q3Em5jED
5cSwn+X8Fjg+g+ZOBWpPIx3ThaB8nNap3Q+FJwoEsAXj+P7eX1aYy5iA9QPuycTB
iBzOgB8pNFVNEF5U02MMIT/zOJptRpDymF82Bw7R1QP6GrLHYA7rB3XNT1kj7n8X
TxV5mSE/N4UKk5j7FwTXb+84mREEgkJdnpWkNLxzubenvQhcap88YYi+p2Eh7MTb
2UaSzi9ogy9eFTN+3lXwLkstIjNGGUE8VHGjz/crVp69THRUXEnbFYFhJtiouGO+
WOXZEW+yGRo54dpB7vm8xdgoxNeJdSxUIUZmigkEY93IN0rMNRnpUY+64Tc/M4OD
FG4dJhcF2hEuRV7PI5oNAkltMeKnIjZEz+Kchxl/CIjwxB8zctV1j/OUi5LTrNvv
4fZC7emCSBra9D41y801bgZ/bm3b55hhkLO9M4DDskWhYGVCLYDCF+pMx32Dr3Fc
M/uqEJagwZWtb/qgNSy8455I1gvuor18ker+bZ66/svUTg6AKX0j0+Crx2Vr5xph
0wvPMCbOq+JV2Xo5zxeHvfZt3xBWUaTziU7LSi6JUGTAn8+uELbNYoY32323t20L
nUzaVn9obpg1fsfAu7HT4dXjQbEt1kh6XnwRghS6CPTRD95LfP+E2vQfNu6a/uzi
TluGNQaHbExZQuExipTh1/yQC/KHF2gh6kta9IJgYQE1cNjES8AYdsqzC2czE7GP
uwCwQp9nqmm2ODoQFg+6HEYJusm2TXXLJOhxxds6SBDktdHjL9QVv5IAKlilk29g
9BQJ73YZXQWLSbl5cl8nJChGACIW9uD67AO4jA6gq2AfejUDhmmJZJ9wKG0vt+Au
7RL+DRsHHm9GAk2Gu998gb1ZUdWZD8lFWouKykVragQv15QjKntSRSXHIBpckrfJ
lct2sR96CPipzODYpkBsE1g/I9uQUMLBa81wJQIaihTh4Mozw+09zq48RJuohONp
BP87OgtFc1XjZv8aMe8zG7McbKRpF1RbJmKzX+yRSGoJKNnppRsEJFsMI9BIixeO
N8Uxm0EysXYkMII34GFtsSfi/crm032fJjUzarnzb+uZtG+uypFuQ8vTy6t0C9B7
qnQcOT4I304yJMOx7DkWcGd7NCCJiaX8ZwVsUHOfoNXBw1VNhzCDMyI6bQuc59lG
p4/0e1mzT8OkIQAUQIR3b7tcncvKek+vqdALdNMVzbMFBYZG2gSUUxQ3Vnvw0N6V
3pWX1dQQ0jdlRhbt0CyX5quq6p0xvyat0odg3XXh2ysYOyh91yCEYCDQIcI4N1Qf
ORpjjIKzFtWokOatLPwsGyAaYcneA/1mO9z6qadldD19RGve9FERoPz8w/U9QZt4
g+4wDZbT1EdBLX8q83NBvw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RO4AOkjXNeI6bmJEtIMV0UqeZPf3vuKopJMy/8VSeiK0G0i6MiCpUn+piq8HtkQk
P+iqmu4PJ6pDhwPQ2uIFWDjZIon0YU3zySOWePJyoSnAE9x2gOvirBNlp64OJ43O
Pn3wecZOyJHnja2KFjgG8zABTknuLB4W1HEZVd/5Bsz2Mp3JmRC0nsI+lIDXtp0c
NhXFcxOimND5muvNxIlAS8By+Mr/nt1INOw5/GUyX++TH9Rlx+CoH+VQgroFNEC1
UxIFxX5zZJxATA3weq+Oex+LzAcGSdZTWsMlyIy11P4i7q02fTYv8uV9TiJA9fRJ
hk6QRFEOTvqibX/Barwl3A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 23792 )
`pragma protect data_block
rJE5zogtdRE9SA//GORjIHkyIlgliCvSqJlhQVOXUTfMPvgKZqswkNJRxrYeFmcE
JDeKwgArEygrcxvskss8A1dwLn5t288fCyQDjKq78lWuomeDNCSfwXjCJ2wYFOEA
GIxeyVymzYSmFkwqTPbM+6saEzCrYTpEZVfR+42jHX2xNC2jAxv8vrcnbLAQJGg+
pAO3fVXzNUGePXTVOXfiRJv5Ff1o/43enqjZl0zrEUx7qN9MkH4aHoVUb8f82Jia
9gWsRGtq0cf89noM0zaCl4hmj/QIpW6KDQ+mR9umdDqysGJNY8on8WFAwzLmTZR8
NwNgNpf4CDDn+Cf9mVlppX0K8Emx9IReDqbsLznv9ASJAM3oyYUK3H/eLuMnw9Ze
gNex50JR5RsghCcodtv7FbDQya5d0mgCOx+u5TZKKUB4j3WljKXxX1FVUlC/idPK
C+fxxQjDLiziBNlhWg1m+s5IudOs+i7ic0bACxI9fFUfsjseyko0JHVdnpyoE+iE
G85y/1UfpygVnexGsENtx4wX9HgSR41Q2y8j1CX7BjsPGaBSr4XTlByaG0aL7Fix
wjgz2uG0JfNVfds2fuBGja+HyiZ/gN3dXffYjevxw66iZys74mqtth1eWL7QNkGk
Z03gYPViuPjv40+PbWKO1IhN99bBqQZIbiYfv1r1r4YsVOgwY+DXhN2LGEirST0E
cE6q1JqFYsDdmfH+qsW6z0vuo0S7cX0AMRSr/OdFN/u3cAazUfJktOv2Djqg5uf2
ITSf4WI3RwMXLYTEzlFos4UQ0DZpJj/WD3P43+yqJ4sbNCulUrynD7xtYDitrnIV
4jDqojE7JCNDSV0CE3VqrPpWYis1Jyz2xoARP+M9wG1iABnzWQtJH6dPm6yFYywh
IISIbiMAfU4qwrzhysUriM5joECilokM4BZdFRQYr16V13DXRbL3wf56kEB9oZYz
BfomiwM+JCo+bs83FtQy4JoMbvUmYt3F29XzhoY3gB7NixbzbJpMGqUiM6W8AiOQ
hHjP3F90m9vxHW4U2/2Ipz+MguSI+aFX1V5ZmiF9N66IYikpAMVkNASGpIDWpJ0I
ufQaYncYQyVDmsaR2zFLgf3sHKi7qOFhSSTPcE8kAotw//sv7V5CYIPUKlc02Xt9
47yrKc+KPgVKH/mwMkwdjM+Lt8+M+nmmklsTmtkhm2MyJ7hThIGtQsqbiRRb1GLo
AsXP8C51zFXbKNApa7/GFXIaLMoTMZi38BfH2GlcWamf7EEZRxLzEovQtmZFWMqf
eE+Th/8psbBLmD27HcwS3apeAy5OGIxsuCoVTr9caaYCGFiogWgsEgQkupYavcpu
eysb6bUH9HjVdIxAvR0FfWQp4VOsFXCtpq0dvjCrCTHW5vhJI7/7Ex0rBmxy/pCI
yFWSJRJIsoSDn0hIRk3eTj4LFLuiRLtQUzxCiur2Vp4sBQb7Rh1h861+yCiRVA+U
6/t89kjb6/LS4chAYqtTJtQS+9gqglKLjVXyyO69fPqu/nBikhuWzYZtWIwcj/VQ
n3IZtkUzzkFofG6fthDHeyqYL1n6I0tcsJB2ZviluV8G8tndmlH4X+Hh9XsP4oCG
cLArcFOBM4/PCIPmYPnUA7FLPzVNlAJJrs3HZ68rM1ivHphhwSQRv8Djz2LOiE20
USdFVRrUzyg5TEsq0HEEzqfK2Yw4RvYPBU93nn4THA483Fafv+oceLiW6zrZy74D
qLYG8tIxhwle5xYJsNrghhB7do5YM7heqNWfT6C63XzaWUZy5ungdimETMMZYX48
4eGG7oN4Kc4WjLwFO96AQrcn1PZBCVkz8qDa4kUpFc6U/i3qmlIzBrhLqSAqXiUr
EqBu+bfFnEn/3AL8915gVnGxb4e24z2I9+EUN4mnZF4hnkN1YMQ51YyK7TW95CLU
MZAwXhUnX0l/SeQPmjcCTwWBzgyKQh3OAax1absnyI63GXipYy+IRmh2qFnTxzsU
NBKgUVJVaPCo9WS+OFxd7X4T8uoeZKv1PEfUbTSZA2r6cK01NaUNmQ4GprNSOOHc
XuvwWqs9cywmWFo8XzfpawDzXg+1+rTe4xZcVXrTdN3VvjKDIN/L3z4KPb+wn9sL
frPPBSYWD4dTX3/b1gsaxSrRlvgJ4eW/Wwp4heKFwcgFa0QdPIkOq4RkwjnwlaSm
mpSluVNIgNymEXXsalVHhhOy90c5r6aft7VuqAfz4y1jdIkAS4cvhI2xPQUvWIWw
wOaJjEm6BJnqZyUrRIvkCIIie/ce64jGTLBsrdeqCpTY2Ixd/UFKLdGxkPi0bn8Y
ecEBaZFFsXvz/URZAwf9wnGH66oP3ad2kij0XvDcwx2jMi3BbVewhpGXgpA/NmNf
h1ba4KZUC+zYD39mMXaFHLDTIfc+9RXsMAzuNBIX873d1z3bm+ZOfQyz6eUcTR3T
XCPXtCNNgsf0YDH+h4AFwIYsoGqtF1tyh/8kz2gbKyv3Km3wPd8f4cy/jhfcpjLF
9yfgBfPBuTVJ48Su/UDFRxkKswZ3JlXbwlmvJknJgd+IkQzaOvBTTUEzWVCaf4ZB
kEUavxiISAJq2xACfnikDa4bgeyU1Nrv1AgnwQyqIOPdfBY3j5D8g2bILONeO8ud
wd0bzKYl6OC9pI/wlvDR95GDSNSe5F8TpsCFc7OwFliDDSMZt7/uj8cYYjT2aWZe
FSWhFTsTjFNUHJbwc6Ly37NeqinbDyir9EXjtuHes6TI7rsKRqAfL4+LemE7cUyQ
nyQIQIqGZ6Yj3ys77jcf72n6wblviayY+aV6kcs3ix1n2iEX7In1A81hyDD5a9lg
/mYsKiEgd4+iBpvAW+C8XACposX85y6XgLQ2xpRmK2s6gY+0a+5psmEhByIHrx9A
GTpzoyw2oDVqs9YMwLnd1PTzXam6PINAES2aIQyqm1I1psAoOVHj5SQNm6a+t+80
kKyW0DdEx6oSYtN61t3Zu5O8LO4tWST2cZtoTRz5hfAUpMN57aVGE8QzaBfCw2Dt
6epb2NCFSXLfllHA42OV3s4N1WqaQ06rmhaqaaIF9WvKpwIiIjpDXOeMqo+cTTaC
83bvev2NFjabaPQMLzRnM07PNWvjfaZpD1xD3qrm++fyaof+JVw0p8xjW3P7kzJM
tNpz1iycKpv/5ATOKexSzzZvJWlf0xg+rOLQUqwE0mxb5ukM+1+HNxiSofb/tG2R
whk/x5sG5R3lLwDIt/YybZwnqCNXSzEhGJq4RhhHMf2dp+cDvLb69K3E+eXDhjfA
FeJht4DCLmqjBH7v5anFH0fkP+hEuZsu5KA6FxRI6QoyjmoQtln1ezcH3noM5GpM
Yb81XvNJtodijku7L4fzt6dM6C8PrmkQZnnXsZuq5OzioOy0pSoBJf9b5Aew2lhj
zt+h0NbDlRUdPYs/TzEQ49l40HvsmVUmydPgIcD6x4tlO+XnOBQgGEBUCjI1KPNL
bS1fiRMy/7dmxrXNf9RplCpJc9pmOF0LSPfzRtHuxnX6hyL0BhhDawXhPwZfWDiw
56Ot6bQlu29O0cwXMm4GLbfISNiE85bVix+10ucuQyBaF2I1+CTV1EWndU/3D5JN
mNRiQYCW1rNRsNqe4lRZixU3OpFLbRsJZZXkOLJ/KNm/2qS9zdbPxkgcbCmCnDCS
Fgdr9L7OyA8XxqNSaR61qbDUCEGMEtd/f27T/I3+55OEjyIPx2F9XmZv3KCdXK+Y
meAronzm7dHdpfyuMabTjiq3G/QeTcytp6Tg6it36EQz2D/G21byibZ0bJQvV21x
uuERK/XgiHWjKWNRktEScw17/lT+YC+ZnvDNK/x+KUNnjC7iXFS+EXNJzziHO3xX
kShsl3GqFiuhNzTGjj2mTXf64gBYe4/s8iAnhbJLtPtgI1KLZ5Xi94zE8AmO1bBu
6Yh+vDwQ3ZzQYKdhdycg+vxnKgLoxsf+lEjLnoNh+AP8hGCrSoPfUyREanCmdbmD
EAHgoN1iOQKOx0XTYqVrPR2oWE6q+iyn4OlmJ7yV0Hxju4GjrCDHBCiuqlx/UYJK
skpJyTo/by1tWFKt8BndkzAKS9hR/44KCJmsuI/UO/sWHRm5XKvAsuKcs72rM4Ks
5eKTOsYGLSTsJDmcDIckOSREZoRAc8U3n1eFGgkwJCWJHzPAg9AwqK+T4bKZaLHZ
QT6l6YdgZUhZ5IOevD8P/wVJJlDj/XFEbmbRjrVNxcgfn/2EncAGwbCnjF/N3Rqx
vjhjYT/3bTkl0/GLgqJTPdfCDS4EUt5MI2cksmo2pCPwg3zdhV6rw+vUzXlf7XPl
AwRb9nBxwpfwdHu8FntOf+1OngZ1vhaIl5EaxELQ/YnxcQgjsA1W3rdIME6EC2dE
7JQ69/HxddSXY/uEWiYM2YEGHw64oTQejtIGT5M3f7PpaDw7Un2TlXiysmHsxcMt
DUPcJvcyQM2p0VPhVlXRJdFVSEXe76nNkjEBt6EKT4T2TApRkOZ5KnG60j0SgS3v
amnTgCsIVO2a8J09yoQhIPa06hlT4nOKIu14CuJVZX0SBXsD4/0vmWNgj8lsvtAB
KMDKq+J6lBAPL3ToL8ymqnGVpjIO9lMYjWR9gJR+GtUVWN9dkE9C5AQImTYcbmvn
eehIxLsF6vTsFrxM5K0he7zNAQsbFMjlP9Pz88L83LfRn0DQ2/t97xEZdoHOFczW
A1e/LHNoEkwoMq7Dzndd14YCjaqvWZy5ir8Xw1ZWZehMSZPK07bw3C3qjBhkoHzF
42jzmePMHxhLDDANmiapjCh5KC6/EhQwXF+/gHMkgHGjKjg0yZj3LOcEq6H0Y7sh
kWCQAy9NUbLtXKKaXcAsTVIiHqOVJkX4EHOg7kmpagAoPgJ9A7fENFmfs0ARKOFn
4OJEEHC59vgq3DgtoU56gmyisKalP+zj46hSuYpmAP+qduP+1CkuRvgKNsPZ3NMU
pKDKqb+PSmM2nnLINDnbWeN0nZnMHBzqpyeBjlLn2Mmesow3mTzRBM+o3nGWS4Bi
F76+faORAOuTt71tj2bu8HJLzdoiZ5VykO6pq4L/o5c1y+G2voDBcZGSqTNaSCmJ
NWyWwhF/XH03CFmLd6uN+GuMxhLa7Dvocef3qNHPHRXNciWypjvjwjz5Zs5paFhT
cD6H4ptUtz/x8FpiMsM6CuW06dUO2EGuaxlllzpx4/SPuECu4Rf6CjvYMnq7YJ0B
lX8IEtKPpNb3Yxjw+O34qCKHRL81nA3HC4AmGiWCpVgok6FbwkhP968562c3JWS5
NX/Y+Aik83dLlq8FLOogCFrDzF6NAVTY3vDjgB25DuIeiegPrf2eeTxJAZ6NXaz6
65yzNG+2p7618Qo1z0I7BFcyq5cv1nzWJYX/VXy/fpDczNAbymePOOiJ5O90LBYC
lbesTX+VoFycR7+lwhT+5+F4kedDO/HEBn1iyUOQa+PKOLZ8LOUfM7hLkQj3zbae
wvLHGqj7BQDuSGiFAmIbPUuWl1slibe1lPahV/PdD4MpkY+zgYT0eOHBtsje01fp
eVSBu548xA5pcAu/jN7sCLJXWCGrlICFPoyBUCuwTqC0S47N+xSaWby4WetGu8ux
dlY0g2GwUzOYtt2CC6hWRb2oxNLgGBrCcioom/I5uZv4REc0UdTRoZSDK6gMSpzK
ai/SgZOmbQLh4koTpnc3wLyt2zKZLHccrI4bfyDbUwokcUFHnmXQsMv/ayxIFvnO
2+mjZK/KlcfAe+wye0HXlLAaHXWb3VpFPlgEdhOgJ9uXIgCWC5hZorr/Vir4evUa
I2Fq0OXmppn0NGpE2bgPICH5ap/vDsU3TZlW8oqlBMNTRR/jb5bi7gmt30kOUtHh
Yh3DUuxzJqwwkg61XDrBUwQJH/dHqb7LR3a8ngRogygyoEQzEg8D12dGTCQ+KBUX
Fi4S6WWle8E9h3dUigglJ+nKStA0yG4DzpTq5Y+0bSaz+Cwx4TqaN9QBHj4764js
fjcO65ndaPJEb2RGdheW2OPPR+/jAamtlWD5/cPSVW2j9H9fEvAM0Bh5F8pE7sdX
1LIvjrYGtalymkBrnAb/trwYYfKz7T7FP1ANquNfzjCf3ThiFUwLGZmFUMRxbvy2
XiJiJDV003x5qGE3+/YhmaLdkHgFvCVFTmUvfAl7UHWaMSHgbEcyTUW3TwNbF57U
ifyTdTpHiIVnCkePhYMTTgYCMK9gReeN/ztgiHSLj0LL4bW4/aJI9XmCoEmgMtm8
dNA2lzU2km+GWwHFPL4TaPNoevAu7u9IzMqFTsVWshmvMiJha4g1sHPNKrqG9g/P
TeRfnkQxeCMgOvhfDgmyJxzuKi636FsVZ7S63uwcHpK4y27ycGXrRGpplukTaXzD
Fs4vnFJiiZREN5OvI+v7bc3pi9jP/IC4W/O4ZOn6S1G0g0LO5oFEsvZvqSTwSCgw
LjyDLCWshKRrqWsX5tkkwbekZLy2IWXiroGmamLOpALj3eeo5GxobK3uBSzVF1v+
UVkBWkcZrI0KRB9bQVr7mlExuYv2uZoqTGqHtOnjxSyz1kKAYmYEyH8K/mhfWkWy
Cc+HSrAgmpGGMFs6pBIWP2Nxx3t5XiQf8oXWE9wybhrE67tordr9FRWDoGsBB9r+
F5EFg0t3VeWe0m1bJFmRZJIK+6InNyeVn0jzjdeCHClie/l+fBfzlA5rQvw9aPe5
LM2AzHg3mTog6Y+5+KKwrFauUJiJifISXiekLT2hIReZsTFp8/LUhoutrAEiv1fg
S8ah5IvPcoprk+u3H1pud6irSAz6dZBLhhaj1VrKr8FD5Cj1Ea3CZOSG9SVtGSxx
VuDPTg1jydQtRw49NY+lu/kh5y3yFYnuhD896kAicUlVahrpxbTvOjTynM7lPMUN
vENoqJrsl0VkMO02+g0AONtwaQdUJx+ODmwVUhpIJbbs3EKTRh9OL6VeVdS4DZL9
FfHyQo6blGzwD+IvLwhsDt4IZmUzQCiooHvfv9o/lqWbPDe9u7UehTl8qTPgwF8h
wA7ufyS0GyyfvtvbbR0FvDM0MI71WaGDPtXNC1QtDxCtbTuFbQNUmggeruwWpByz
EY1HDDv9aNNNQaLMuTpggRk1hq1T4ihbbbPTOkGmvaETggvFsDzOblZdtY1t/7MQ
9FYoMf6wth13slhp54mQvfpXjBUNZUB4ZKGmOPD/bjdu5vBNChYGwEpM06fEyTEq
AnkQzaZNSw8NChFATQXh63Gld87ReGkdGvju9zCwRom2/8/l4ELiCNUgKKLo5J39
nVEK7Hdv44YE3sQlFJbxZ5ZrOnqlFFvX6Y+SFuaBmVROmWn3rvAgvRKvd2Bo1iU/
fVMueovEnINS0J+pjNG+US/Y2hBUkUDM3dHafF8piZEfYR8ZRDkekw7h+D6k0gN9
mKRmedKmw3BsOXlFI536j+FY8SdtQTskwjrZGFtc8WRuNGFv6EfanFeUj90KGgpy
qVlpKE1+Wz6CsyG/FDZsBcLCWh0OmPIRreiuZvN0tYyYmnxqEKteJrEx/8Z44IsT
VjJNHh3hCY83NmmSCFjgZbLXz1pzdcEmJevCNAfLuC27Y6ytIEy4Wn70OVDB6M8V
L8RiqL57wstgK0IjAB+JT9zJP5YnfhI+nA/pZ8KLKXFMBufWXKehKCxnMUBwF9Be
mDFCWwq23Dzc8vTmb7mSoCfUod+azqHn4VmSOmD+uwJKsX2ysLGzfvnPhNmgm0pL
W6t/ISzUrNuqVpUpn21KFwcVNFXSTMCwgKTTYRbsPAa2f2f2ZUPk1Yy8hvuztRIM
rgcy+zloyu4SFdM4xe+/HjcnNsNCT2MMS/3rFuv0nqJa9OjwK+/3nfK5hsWDpQnF
8+WjcKVOxosxadJP2oyb/j2kIti62knoPbqeVltN8Lw3Cu+f9IHU1dHK3GMXQLkM
U1F1Ab7+3u/mCDv1WT28ZysnpZi+CnWBWl3RXYDjQ4ElXaPoo/dteHQlTZsqZAk6
gJC82oO4tGTrvLfSB28QYkFB4eehEaXwqI37RNrmX3D7hPmLdGGdf97MX7fkY9cy
9p+hs9iWeM4j4bQyqoBGpOZRDvlckskQymS6WA7cGGxINLkGoVPd39EkGbPI1i3I
B0YIq0MevkujkZU9i4Gto6G7Zk5UA/6rMnaZ1qQvtiDql8iOLOUp0tcOxmEX0Kkc
L6cuR4nizrr8A8NTXrD/EwCFA0wkAah4rxz2AkrCLlXLx5k0qPQqkQLOZQ43rtTK
dz88yGF3JIpoCd4kEW4pOueC2bAc2LjjegCBJzifnkpYdKF3wePDkyvFa0DZ7gbM
vyrEDU+2qcguvnEWb3ZMS/RaMeAgJwme411S3b0jCvLd+uY8FEaKsrd0xVL6I2zo
IydtujftXjVirce6juxVudZbQf0uRRAwT43bvrLSU6CS413ivs8VHYGUlAa1XtuX
xeEjCY0swN4uOwvFvk/Qi1ekQIovKFC0gD5sh0SXlz8fGW+skS88mR1Q6rzhrB0h
e3PgzQgKsUpn7vCWo+x47QIBiH8CBPpS2E4xJYQaxaBbsFhuP0BGoowaGotgznBC
AMJpFbG/qeNZ2/TFjqOb5lj5GG8PePCPJStCVamtnpWzvRjus6IR7XPjGt/6SSDr
rVZO/d+0gKYLBnltVoict4O3QanTkPm5VYfPOWYrV/HK7Qry5LhdwILjHkzyiXWM
wbRFzp4pl+Imee7Ob5OxRct7geTROrSSyLS3N9sEjgudPVnXYx8VWIjQ0fKPF8yG
IaOgU/hVw5G+OgZignsb02dCpldtWJEs83BlNuVd6x9T6zH3mpHxNodr06U8Nix1
Zc7pxsiEE+tGxBgkn6aGd3jKNwk81sd+jp2YdpVZeHNx31R6iOdLD0KuQH3+lKC4
Yu5vNlPGZBXX9NJHady+dOEKrXTHUTYhxDamfdSDQzg8kXpJ0zu6E60q2044jiKk
7RoVVL35KqJkBFJzYvsNRRbf+AvfwaWx3RY8Dg3ZOPS6MQcnJECtJZwtjTOAbsT+
K4OBbQDcG/SCf1LtXVgT9Sb6FLD1MnCX4w3nUG0S9HfZVL+pB/XnwKt8IKfk15gn
vGU/0rPhzf+qhHBNXGd+TzSeJ1+W2JVHX7QiUUS8pLHiYAChvJoMNtdYAG0CAhN6
++kM99gMzHdKHMsm9oJNEdZcxqWzxm6muvekA+yr+5fLXVW/YV5/yrPsuAKS+aL6
odkbXrZYUAGLsR+zlBfvsklIXAmtYPrZINVrnzVI0Sd5f+YdDeJqroAZifWpQDcW
F+12HGzmTVk/l5geUD3VihMgZAc3jvEF6lc2eOH1ET4B+RyupPALEtScfBKH0FWl
TWZMDe+BPxM/M9ppDXApCJMkyoQmUHLzE1ZJVpqGxGfoatDFWfAwJV9VsA1LMVrc
OR06Ep60X59GYkj+NQuadlUtcL7RljG+LhicZJslpsyOo3quuJQEfwiejRZ2TD/L
nb3GW8QJbfb5VPhlxK6Am9a/9fFnrDNNy7PPjtTQP5pqe/XZN5ONBs+mZ1SKhczN
ust0BQjdLzmwan3cnPq8BRexCm39ygCXAliGwlJKEetyWRUsmhACvRAm7YmZqqMr
hCT9UlZwCi61Zu7JBuwwg1LDyZHWEG8a7b77DR8QWZ1MwuHxb5UnYM1l/jsUigxD
64kBsUWKSxj1JVIcoO4D5hOfc7vmyUfNDXesKkzKGaNAF+2VpXJKJO+HBGRmdP6w
J/TKkeoFdWYbS6wXT+L/LFaLG7EhtnDVI7DDC9BLRPgsy6REDmmGHtwtJHV3MUaD
sFDMTGEAy2pi2bGz7WdwjbWQm3VVKKpoXoCjeJ9DaUsMR4W6/kVcn0ZmGALlEdQY
KwsWKj0CfVbfP1NYuKDdny7TccgI/lZZqNrprypmGKrE+InGxXIy5h1Iqyt/USqV
Z7Stb2+GxOQ8K4V3TOXCrGYD+sxqvpxzmcJFMXTrE+XN0el4zk0ezRDBwHbAf6pi
EwyhroVm02TQfCS4xU4G2OOKbppReSIZYscVLllYIl2Cza7T+u+0Q/a57LcfdKA9
9Al1O9PMKWde8k6w74Psy7mWA7Li9VzK7l4CsvfZWlPb2cSABSB5uh1pB6JxSBDe
ZFBjEuveQlET2m85z4UcoflnTVzT6RYbagJkhd9X5M6GH3OafH0AabYJQP+D0Ca2
Lqi2c0E5KBhODHE0cKpbdkygcmwtrna+a9rAczt2JbZX2l4enTwqvx1FVlrW6nJl
uYL9oGOhK60R/JppQMcXBe/ew2gIDBHTKlez+kczBFyHGc2OYU+RS21iWxMXpcej
TMXY8ytO68dNUNEb0uP7Tc2lB9XwholyE/GN1Hz/RU7E1hy6NwW4+87Eq185gRim
IfDq2DG0dDLgJHyagNcortwcqy+TafWHrcUlg+zaPyXgW/RAbq080/eLNPkIAG0H
XR66HYr+JqqP+dBasDGJAX26gifeTA6ZB/py7BIDy4GOBL6Do9ARfiNXnblPpG9+
8Kwmy70KKj1RCWbTXzFwKlWhFFsaUbvyPtiPfI0DiRqMC3hPiYQTveMZMa3AFNwb
9TvUu8l46aOCzu13ez1hlaYWb8BeD7BHsestDlgGmVQ6HNAhcY7DHCqV1ht9VaNU
xA1ao1NEbHMjYTY8zLZaY1lt/8CA70StAKCcdfLg94umanjgVOrKFaTUaa2TW4x6
NVuEAAwH12+OuNAVIlu9K7X4hHsch74GMK6p/BhpptvF9AyRZLXAsuzEUHfQw+NW
x7TUs7Ka4lj6o7p6fuIdNJTNdj6ke2dRlm7jyzIUznykWMgC+S2rkBE4hWNJ3gHs
0nICBLfh/pTp7gdGrhuMdfqM9CA/vx/7guTawgGQ47ODIKIOApbKgovcq6uhQgSM
bIHmYp0xQWnobZBOqRlD79LpkMM1CyTWrSokD8HzWaHauu8T2/+oTXURj8ISjYF8
9fADiSrF3PECAhJmaOh0fdRWbBed6GzlY1r748QUewd7hM81Eb2XQ6MRQpAcdyot
asYYfwEVvNpODb2G88BloqkoasXdOk38lxu1UUjb0V4BojlHqOwHzgoXZjSbygPH
c3e4124jzJFme1VdLedlTvDaGG2tYXfeFbv2einbOPdwMepyNCVa9x6NwU3NDm8I
eUzMZ48e+0/y7wHxRi17D18jw7UXexjg9uRnlZvu+Gm74NnFlX/mYaO5tWp0DxMf
tOd4B9dkJC3FiMtbpr0wi/ycmYmlm93QJvH0NuDJjxLfTNaiwneae/IOepdDSjqp
NthA8Fj+Tf76RYEaeLk11O60R3317nk9hrOW1Gnbn1iVrbo6jTjfQXFrGPEFvWDK
cV+Rzr7WMu21MLVBXhcVglfEpLSEGLj0fCCX9+rzCcXhREF8Ipe3ZcdoYiDhNsZj
JER07zUiz9QHcFx5WYS9RjN/HOuqasVcJ9r42+gFsU6JI28pNl3wOXwD5lZ5devN
GHC8RtmKwqrRuv2vDOZK8CMjRmn5kdQgDGyGuxeUaA6u4LYuPplRlqZ9di+9r3OD
1qAN1XHKxXswExx11ahMO3QlMz/ioPMAat4ZPjBHyXxY81/3OyfOt/51czGYpu6p
9dhQmQbL+I2cbda8i0wzXpqqjFCPZWdcs8v49vcoG0wS9p1sojF9AghuCMaLr9Z2
OzwEDi7G4G6AZ0tdkCXjy2yptV9FCNABkeaBORJLCLwgGlk6TFzZglh9Dg/83/7j
HizfEoDePiyMQBdcaz577Ehmx3jnaETQfOBdkjRCCgy6W1dlIwx0sjcdS0w1gQ8W
s5jTR8Js14nF3xC+xF0RCLpU6/MV/wm2su1hsF8TrGiHglyzESuA1fR8XL1WznI9
hb5wCqNyVZ5xJY0KBS1dnkHiCdPFqTE3H3/kLmVWUDamHIN9VXE7nGdLekrNhhZ7
kSRD846XtlPEMLmM/MazJF2Y1GVPe+yYRDsiBzDEBANphIrbqiiA0WmvXpJFXSdL
fzUqR9yempAueTch+Be/tDopiA8JtGd2fctKZUVfInto1CCfrJaX19V18LjD0StW
UGefZVCvsW16iPMAnubFp2b9TjVWkpCAL14BeqKwFkrTn2iMuoe5wY1N6VqWAI5p
BOi2DZqj96mM1sZFxwgctaIHYvT57jLRma9KPVCWlKlOS1An3f9WmOrxWelaJQTt
W2XmO/gFY3/exLuCRL3ipvY7uvmKry29yS4XxUayXi6IZRrRQBv5CWRkGaczX9Vq
Afw3/w8YxU3u8iZxcsmvTlwMLbqibUch4joQEC0euvHnM0BFDvQBpt++tBgeauPp
CRLNOv8MGlooCFrWDs4BmgAJKYcjuu+VJY0m8hlQDx8J28pFPsazPd9+6PEsbsxr
plxGgcphYKpPL3lY2yJEOynABOW3Vp14E0T/tpcSpCmz2eNuoGSRHesPbgWEn3Nu
dzajocdMuFWIfVi4GzL0QuGIPApR6kLgT0MGHMZovwqJ02d84sFY7aWO2CauKynK
ssegumFVt6NaVfj3DbGLfkxQwikZ4t2zVOStGClJERT3MQBz/VycNAfCR2xA8RTO
CiVbq/tELjzJGGXON2EBzWcCzmMRAx7sHOaeK3PHajRHjvFYS2b1d1fZ429DR/bw
tf/E7pmglBYk+cZ514398b7I1Zd7/Fx9eBpKRrSiRFd8lsbVFqAy7lNuH+NClSDS
fOG4wuwTATi4LFnbySrdKYHHQfkmOzv9+TYHp2nwcsoKRsfsPJcXsmu1geKQDJa4
8/i/S9Z+1l83KN+7zToUhT4D+IZWMbB3Zu4GRhXAGRLBbTjgQWt9NwFTY4Zs6LsL
62uHYRa/4vk3L6UcYGX5JAvMLHMJI6u2/PhJWZEIlaR8EEMgU5+YyvIEPH73kHr4
B6/i5AYdKGHQA416f2JWRSVu5wT64iiJy7u/mRue/+MfxR0jdVvH2Yi9SHkvo0R5
4W63OwMP6jk45DI+DQUM0TevDbYChauXYtGtIjCeSU398qqdhwqVDledTJ6cE5Es
VO4uQXtc4+UQcCSbX+lGwRp+TFsiY2pJpY89Dr2IHlsrzih4MAMauk0XElotuJim
phApZrVL2QJSBDFd5LYWmEsW1QH3OChJdwpmzP1OXecStstUC0J8V2Y9mNbkx0nF
Isw+EZAe5u4s5ktR3BJ50HUkyUhODrS9JjhX7CAooTzyW7QjN3viD6tE5JXmhuQe
vCKgtF9INBF4rYjdB464S8M869PdwJzHvidKY8TZ3D++MtnITz6ZybQmb4Sg3D5z
7l+JJZlzrOLP+ZMnMJnVpnbqBjg3UlL9YDsCSo3yzvQVwnw2CniUUAjjlo0gRJrK
Lt3pW4Fpp+GE9eXK/MukJbblzJewcogXM1Sh7IU4CdkdOTG3CiFp8hp1nWAMBfUi
O3sqUBcer+yl+KNFG7JZoT6dx7CSoMfi70pXthBxPzlrAIwuhEsMApMSt66HIQET
Y+IhfKZXSfzRgnO5TNVGBUIcRsguDci4YtuMpBfhpkKH8blBrl7gDlebhP3syFZN
PTPXLtmk3O/FJ0EzR3AN18FfzJNepGGhPPhhZdPhYRxASrHZmaEhqK0vVbmFc/tB
TDaWcVwqhz0TdjgeZEu4mfxl08Oet10A86XyJxdFELr4ZfhExD8J2n5HTjCRxSmX
ww53zLgnYV0Q447UntTVrRcvdc/JAh3odDwqr6gBI/b/r2ymjG+gNguqR4TKU45O
TO/dxwaD2XlpStFr0kFyD6rMJLSYgEh3kFZgY9D/gJRRr/pOSozmwuGIoE3l54wS
MMZCqtiRbeJ9/2gbht8NPeXOVP88n0+CnvHEdCi4UL5CDgpSHU28fYuGHK03Akdq
ntW9glO7iliBazEtP2gciUauD7Chy46zLfBqj+9PfAHOHiLOIhcQRcCksygPirYd
A1x2piILC4nLZdZzmmAUtMjyy9THPmgO8YZ+4M0bRe5Cc1jXvmgYQAO8GZXSqTUt
oYL3ZqsgM6dbW3AAuNbKScEHKDG9PQtyLMkdGpt/GzGj/lBXM5sMmIfAZJHgDAq5
9nhQLUviLasa4NmR7n1y6kZbyVTW6DDcdKWhV55iPl2z3hbuPIz9cFq1doABuBqe
hZjUxUQzmXo3Zb6goP0o8uXA7MJNgglmSqvVKW302UNETOxmDQQhn+v6O0RUPJGI
+X/EnvyrNRInuoOctn3MH3GUs1V8uqzGwKnVXUUVFrWrdI9sE+rIyoxLYIUMWQZY
jJNaURhFtALFcTcn7kJitELiPzN6YjZ0hxdRi59uroabLHJgrEo86cjnj5Aq/SUM
ddm3wYXkmZC7aY5TYzE6SJ/vACwMqr/5IAG1u9NXIud11KDXWQHVxtmsdHlOeMK0
EbSHPI03GK2GO+K4zqKuC/xC210rClmchcbOfU8vVLiu7axwMh1MfXvd+kodAPcb
f/J3B1aZTY0DB23t+MM7z8wr6xcED6p/Hn88J6XXAeEO85YmSlD9S4ZhwXMRG5SI
WXVmrJriazbkyjD8RBokjNKX++uFgHekb+Vi/e4oSI/O0+H3kMfOpft2kyUvwBsv
ouynQvY8j4c9NdA1Y5DB8C8lZc/rZLW1YeDGhCAvWXYqxRR8RaHdImlvPCFnGN/s
MKkxE0DxG8o0/+I4IFRbba6O375gGgb72JkvTtUbTxPtiQXNGDYp//EEA2fpOcYf
bbnEK5hISJ6BiPDaFNho5zduEWwQqOW89JNBCUtITniiOmSBSfCfCX3OHfGxdSTu
avW+pGQheRFE3uDZU+ZQqUNyDPsF9T6p37xZFYaWxtgfe/VJoIOcyNFGVkm7E3EQ
q4AXoDDBw4EomcWaHC+Edfxu1d3ubgTCRkN3xwT+WtCtYbOicisQ0GLx220lCHq9
ue5Glz5RHdGl8eBFKXNnSm0xYVt4C+oIteEeSmQ8Eu77L1mpu6yCeStKosJ0qAHn
MaASq63Ng4Fk7tAgzhM9O9Urzox19nRrhwAGNOIwLNKR6xbmMzImMrJ7h+uxmpsV
BH7CCCWnxyK2zE5kCOoe+bpkg2YB3NVtUMZ/E8dk7ezKhkVL8Ld5fjE2EqeQY6UM
QzV9mwL/bGMl0CnnZCu8xITyxWgaOv0ktzYu7AELMiCSBpcfS27qjP/sg5hr6sTw
JM7zK2swRpU43QOghdCSHggdW0aGHGqq3zL74JEU15rFzifm5QktH6M2qcFaQzUk
8Ru81yOvyUwnn9rlkPX/AJvPeriv81Qk4e73vH1kqSXXtH8n9OJvoJOhAWyyBajy
p+uijYpiO4xgYwCyGm1vmhKu/15sR1cupp9XFqvFuBRCNsK56jMzRTDr61kEI41R
0jp043bBFEHdbYzPOQbMZOvq/PjQVtOi0cj5AUp/fODb4cgAe+kY8oWJMVQ3kfCb
Dih1nV5BuDgvm+YMJ9Rfb6fzJxeZDsxZvHJs/7A4WDa+M4hR2w6oDCziABQlQENE
stxfWCI2Vu3zSWTAUivPj88NwQP+vELhcBqyUrwpRjXxMeOtw9joH/oU69KyR7c3
zQoJQ8wRtwyniq40rrOCtHti8vf2aqBNf4dHkAtfhpVcvYtuaYujVJ+1eqiYrXeo
X9YQusi9mF8XBG1VctZuXeJ17hG4oHpZDM0CcxdnyGd4Jo+npFwjgn1OWTB21yYf
dMVh6X3XTzmESWfby+Ufx217uoeGn1GGmeM3kff8w3fftRlzO7PwKiuANTZLGK+X
XseQjPUiD0N2VH+7B2Il9q+kJ3m0CxXWKw2jUMW5kLZoJdnjqQ+rB4CCk792eqrh
C2RCt2/twVx97erC8f3SoYcOI/VtmHO5TLX7Zfs0VzCGJMLSTIozlgx0yG2EQP8E
1a5YAAKrZfiErD1veMEk2WdCf7GHtgP31qcyCIpNQGyoJlmv4l8FHsCLPwFDlBIv
T/s75ZxYs8iS3JDDZKf7crqTSCDJbfrH0Pk9jdSh9IiNo+aT40SKNR607wqi1h+y
BG0eRS7ebbSCx5BjvOdvP8hq3fyWfV5rLUCYmYZbtfQHOPSDr98aKIA7z7dcZruC
nl3I2SfqP6ILn5HZF1kOozqJ/gI6VLnNB5oNdAGDxVDR9hwk0h+LXRtdby6ACfj6
wMy2adEfNa95CI21hyjlzFJc+DHiF2WXQDBX2QcsLf6Dbe0vy426QjDBeiWiQLVV
J2o2xr06xSfjzE+GQ4ceteV1iPOSKy63oRGxJ3khb/xfyZGCONRta/VSiiAGxpCj
UJlRJoFmbf21sIt4qPrgLoXVnN8TdSYaF01eI2TDe6pnmMFt7ufzz9oQfmF44xy0
KUpIU3VqDvdjMs3tQ3TMbGZDDeqS5xp164G9xxE9eTELd2yupbA3LBaYJIZIDOzc
gqTXS6aIXeHYLSvcC3s/5duGmv9bLp7EA1X6f1Q67l17JrUw7naeUL3oBowltP4Y
ZQkP1gzoHa1N3Mzhj3QBwZQiiCSQkAacrSW3XTXH1qCB2ZGqNE5eq5MP08cy1GC5
R/ZA2S8io72Z/k/R0kIcEi3azDaOkD6vZW+hgj1yuEWSayLnsH5dovSiK4wN6Nwi
5Q5C+JcGd1QA2Y4Yqis0ro4LVsC5AseQIzGrE3qi6VlN6MEHulUUYcH9Bs8EYRHb
L+IDb+AgRx6S8+XFh2H5KVSYPQvgfGTjksdTZ4qZ0Kj1YB/MMR0oxyKeFIrzcj4d
yvFrjrnWpUiYS5wn/1iv/93k1BAx/v2ovvis6PuFwmm9YDH2H1p5I60OfIOBJSFx
geptU//JLYy+O6SQM1aq4f1PbzGIbb+7Cxd3Ty9+IBB4XdF+XmTuZCvpVgUxrElN
AGL9SH2r3DHKRtLF8AkC9wjrC9WJh2xOL3ywrGXzuFjDmL3q0/3xdL9cM1aG9icn
6wtV0w3IqKJk6NyjcaPC+C7rvdeX48D/wqhl1v43ZULw3IKWTl28etFPlFRHGMAv
V7sMwCTCHhB+yXh1MBm31EZd3bMlxmgqitiy4zRUGFg5id2SXdykOn1fmxqwlsGV
Qy8mxhqqPZY9IFMkafhp5UQj+1xkRL8UWvLE7h+2epgoGFkfpff7bCu0rYn6+cV9
85Kv/nRKMLfW61Koi3NAs1yzzsFN4A34GJWQ0hEg6nG8ltp0BrA+b0m0KGqf/6Lj
IJAtAsJ8fj0kFAzcPMKATvRZjMiUC92swl1aCTirvDRygGc9bkK3vqKoWAdjQ8eB
sEmYJL0J0B6eNeIbe4B4vxyZRhnghVAhNvPmbNfeF4wmC1nfugIxF6Ik2ONCz6k5
z3Kur/f4+SHZRJkYeO5YxCMCUudsPe8hL10yLSRnWkWv4BvYpXDZsrPYPPd4cVjI
Q3Lb1dxaLSEDTu6DDuFaVt3qKF1OLgmI2+nYMbzRLQncYY26T8rqBbYNUT19jPJY
QvfwMgtpUNX2cj6yuCts3uTz+M9WZV/HrSX0eBsmbP5rW/tWeN85FLYKVSbjDp83
roIW2hbDb64MVwYKobr5K/W3HL1ZIhJ0H+3SA/ixdBtjY3O3Jb80kJ+2CDcd9EB0
5hOMqbL41BlfcLKb4U1v/GF+bwd2TtyFCp+Xv1E+yMJTmJ+rpls+7FXlcbxANsFB
Sc+SVNFdCSm5lGeY5nktnHLRat0t5PRqBjAQAwsVmsStEpzBSGF9ozPLDM2Oy9nC
eqo9yKvmi8Zp3hUpef/1q/crwUroQQKmQnv+9Q36ca9EXTs/onxne4dtysojIc9w
L5WafRNuwmfB/0CWkHZ03fwjMcaENmNTGgzL2ykhrQOn77/ae27rXH5UDlHGR9AI
262n02q5M42uPhFNfj5Dd3xyxLIItmTzL40Y6yhxY/oJ2lxsnQoF7FLLL4Sw+Lp4
2GG440p6LNxket59aXOk+tpOiEtlrgkO40UH/bp3t2ul/3nnFOFb0hcbeXlpwXfk
9cP7u2EPanq+9DHnPiUwPkAK1X5GxS9mEYw0lz9y9kYYt49VfTPqdtivOLY0mSgJ
jgqxn3Rxaov09wH7hMWnumEVD3PJxAfqZ/j5tRlzEeX8gw4MjGkZM2383pOm3SwC
SJJ4SykT6eHXyJT8l6+1QDSJLNZnE4oWcQCNeMYLv8TA7K4YUYD02ZmjDl45Hr0b
mB0LBBNvmCSfkknuR/7I7eO7D1ANcgSX8NGDicHd5HPlpukpyG+4GsX3w6l7uR1u
iiZfkd3RXbgni+shSqgbww92nLDpukfAzuZP7H8FEOrPM3lcHmn2nNoNQugYy9un
thjcur1S3fVcDDMohCwyB6j8fyCg+08HBXcpXzLgVZDVmde5m6Oe0Nc7kt5tp4dQ
jYZcfvOHMACWlYu1/CgN5766hV3CSMS59xoK5Z8tVuhkz45ZdMVZ6qD7wf/nkKmS
2gg94qblHJJ9utepgxqDqfpiO002POFgddPM40F7hYtP1dQ7Xvi+PS2/otBpmK2h
Z7MAzS/2L4y4IviFKHlTGwfP7dOMT55JBNsU//XqJqfeeOaXkF+dm6ohesRF6NuK
kZjRd6DmtsKKiPt3dzg/ONY0P/hSv3e79aj3x/itsTZnhy14WAf+PJeECtbyCmI6
CtXlow55c4WfihBKPEwU/JQD9+u8IZiZo8NdVwAC7eEpVigzbk5iiyRLkDZSpmd0
kKVT365JP6IGHx2VUlF7kELdfWfl01Z5fsPWHMlX+A3s8ISm+vhhMRFPo/H0zFOz
C/7TDqkZ32r9DQpbCeSwoVcE5whwsftYYPxPhU+VL1y2BL5HTioAjv/GyWeR3GjJ
Gz2QnfWNMnzWPuTnYLhDUurf+RjRXB30byhvFkkCcmXGhUE+/y3BygMFhbjoBaga
rdD0MoKNPbzk0S4QOWWq0BC35+nvC3bycYR8FDntfdspYgVyXSdPRn5dbezdvaOY
ZANyX5rEcTFsjMp18figrzz5juYXcuZLaVIioLKz3EZl87l5LnpjRLf1dTqQ0r42
IFjSB4RoxmBaPwvCkjcqN06D1pk9MU0YTeViwVr2J4aOTUUE/wKZ6PnvWFgJRfDP
gx5FMPDpfnnz4iv1yz7ik5kqXnfHQFC5gWqUCcGyGK5IHWyr52mkkFgAtVwHA8Yy
d11FnwO5NjLmZ0SmEB8qDuAvkrhLlp3xB/K5rivLZKj2ROHSp6DQqzLziLAGTj0I
qmoz3TPqN3liglcX1mh9iy3L+barnLY0cacxNEnE1K0+vcmTzv9DDt6vN4ZVNeGb
gjsGZvoZqezIrQMYErJ03bOe8jdwgL/XhFfTZzRRyuqK7pfUZePp/Yk4MwjBHm6J
Kp5N+QOGm6um3+bbTcU0ozk9nM9qDbW3ttweIw4fX9h2XH1MVfaQA7breXIN1Blr
GUZkMAoVZEd1sIuLhiIP41HAMh0OKCt8uqN8MIKB25cQo4ui1jGsj6XwZ2k8Sygq
EOfyLVISYxY4O6FL8KTaV2Q56un6axIBcGG8lD+bwgJbuCspQFxCP4j1Qe+AvML1
wtQk4+m4ihEJbui/We3ZDiL8TQE8E0s0aWmJyC5hyVdqA98xyRENCnBXDrAAvPQB
GZTyB66iaIFYJdtQZioe9jY++iTdXysGKi3fs2iaKdEed2GaqUeWSj+k51JTYkbK
yrNfz1k07asVu2DHMgBM0Cb6RJnp81R8qe8fMobY8NRN3+KbYxSHU7I3QKA0T2wX
T2tE/OvKUZ1JE4eahFAIHsA2Sbi4+zy0cccmsAjSFfGexcrKPss41Rt0L6ocIijE
Hfwmlo1cvQS92jGQZbOWmuhBlRRktMCl6O//8TVYhmefshNkpdCjSSMgWnsj3zFH
tBS50D3uHXqt4nP0dH0ztjFW9WshzSVNE9JAzuLpn1WL1aBkbsGaTRf9pCsqVdJ8
AM+qOVH9hJ50wU+TfHq/5Z525t77aEmVFscr49xE5uM8qmArMMCY3xqJknAtdjam
NYIJUA1SbdICQbC9xYZ36fxGvJLLHYIfVnuKp6oCtCVrax1joAPoC/32GDvVTyMe
ObFlfbkG9rjbDcqeyQfIGemAUv4NH7fvuGy8X5Cx8U5VAKIgEVcmOXujNii9K00k
eJVjmXqNW72zRlga9O0PMr5GmGGmGIj4VSR6MmIAjQcVr8U+RGmi9Tq9FXKoPgKE
ZRwSm5bIQRAS0aEgQ6TSADsV/NOMYbH8TKlUQXRgiDCXRiBfVYR4AyhiKG8UlXaM
dpTCa7LWPgePqb5OTri5xTPeKqinRG6iVvjCDT7pY5yttK895P06BqWkyIXG8Ofl
txdakCV1btEu0wPJnJNdixduE2ErNkuPQAyizOLrkwqOl+UkiqhyK5kCBGBfZTsT
5i/QpQ0RBVtwfmyvxlXfA7bs2XtX1Gn31Tufq+exroTaMkG5QVFwPtioKE4vZygc
zC0Rjrv7esHUJdhYBu3VOIOXHAQnj4XtMmfdutLkw/vchejMD+MhjdPLEuPT/38b
wI1giwHFEFCYGqn4FF82b5O9YUbma9YfiFGMs51daUWZkjnlhNoiRMz1N+b802w0
oxf6u3nlq0ZpscyWQ+jm4n62Tm9qd6cNKxW26pyYgXjmvai/5TKe28QeJMOXg79C
SEG8B3hoTj0DTeqzAZIy9LPSs9oGm+FwzAqmxNXy6BfaZJwqrbJqZQyL5ttUbMLr
8JfVonxEKppQbAAZvMmMAb/4mVsFjT9MyX6+Moyccem9KRTI8kuWMFY1CTB/LOF1
AZWjJCqbLMzmGdIEbkS26TzGgxaQVOT9lvXOX62Fd4j/sqDx470UE5JuBnv/xmES
lPdexb0BIOu0d1wiNS4dm+rtsO/4B9cKPEOToailITYyKXymiMGy+RRO6xXe56re
O7YB4OFEVePn6NMcpxEfJVp0u9Mfp3kNj1uIq/r2z144HKJxbhgy4Rt9QMs939Nj
IAzhRIsz403oyb3MbEKB8Zgfo+3vX3LfiSwiq2Yh7OaGyub1ThGLjeQ+ViiQP7x5
cx/p6UmEYJTvXlgJrWp5hkEuonvuzKA5mSWfdiTuxhvipddJLDwFI1+NYqUjQvek
2XdBgDcW6OOOXUV3tZBgMOoQkVa9JyZuWvBxPMDlJHuYJpTf3JGdJIR5F0Hzg+Oz
SB1kReKpcmFs4xvRP04YXP0qol+BvUkzRApV+kH26w5e+kCprbOWXmC2a5NNiBix
qOv4J6/wDCRwP08fvDYUlAm3iK7GH0uLWYvX7FoYB9zgbb6WadBg9CQZFSMjdecV
JAw8o9n37wpRnddmAvX02zICjabkxa2surBPyuiyRNjrktXDEabZ9kbnFaLHc/c+
0+nMvh0j8cswPNWhO2tZB0Lse5ENfjXOgiEZaRypuJ6lBuNM93IxcZOEwnbEsWgz
YUQ8/Ild2J+RGYmizDDPMlNl68RJr2GBLC619LpFNY4SQzGwrJJ7oNEd+OXr8T/E
EWb+CsaGXDyjHJ6dfCYCgtlOnsE+Tud3RsqR1038ZytyhwHzinoHmWElUPSBF14d
bR0jAiEAffBr8qKMWrEshFIvRcQIc29nAHsTL2H/Phczb4vOjaO/d/kKyWUW0fQr
lQOtRPF3HY4PeD5tFbvSTu4iYTK27uO/l/OfXk1wkuQlZqoAS5biqL58Y/w3Qtoj
iZg2g0OksKfNJLYVNrAuMD4w0NpfE6Yr11J+YAQ86uK0BPlx0NIEa8tMnleR8ZTU
pWR3DCD3hIo/0hIH3emTB8slR9ynbzxsGu70+QCFhcpbn4IRpHjuBDhsx3VQM5Ck
G69UrTqkiuk3fcohZUFjbNRrnWU2FifAMyvbYkuRm8hljzgvNThsBAxaOGJb+F2r
WxtZpZYTGvbE+IyZTkY/OcXfFZlG/99QWuNju8sBUfu0Z/iF5tyzzYqvrY8eZwxN
LIhQ0ZXf+k33Ie5QlTWWvGMH82cDMrDf90x2DECf/E5pprQGDKRDxpLQR1qUi13A
AfN+HssHKtuorvSTiYEoyryqNWSvfWh4GKE/ClsmyEhh8+SZPj1YqubkM7Mh5mYU
Qv2KAcT8WHg28n9ZgW49MQkoCBIb5NpiDv9jKLHMxq3ZrCs2R8sEWIEZq0ty66yA
7T027tEqtu54QWCyjcN+Obg5eylOACC+vhf9zl2w5gmgJQekmiVb6l0Uw6pExQBW
FNTrNTHfysRMhOE6Wov407kccXoSq/159zBZYn9sYGgwm0BbsToigSDxJwg/hMne
F5+H9mM/2v7dsfxlRpl7P7FQYSIKHqHWjmt9b0x92u9M2x4k7fnQg+OBlrY6qzm/
I0oP3AkRfz0XZHM9dTFWgPbh2rI1Monoul9EMcZb+qNeFtY+/RmhtuLNqFy1vbPr
UyBshW8wvcXErSbx/Yyx5baUXDgAXY8cxHXMw2KypHPEl6M5OJGWhx5O/E5IZmIW
TCt3qhoNhvUvHscj4vEfZ0/ykH0Yib0JnaOyrz3ZTnxsu7NOvznmQNJIMbPUJBZB
YKls5DZX+RUV7iLl3Vk31wf1PpccCKX1xX6lm/r35W8gmSBVImVfXi2brvp5hyQD
e3Do80OiSyedHVjOTqf6d979RkqI1sDH+lfy+NNGaFrPse/nFAvN8C0NPXOYFw/j
gAgDmiZ9EBfu/muKABz3o6d7i80VpNDL6C3bOHbo6DvNEw9zgVV+8brWNtmZUoiO
dN1+ow7JvKqcvpkdqySjtZCGUPp3SpvLjrH132VaWkFra360N3VWD5P4IJSVxXdV
jK+808IM/eEPCSdlaul8lFUu/oomL9zkeWwSi4FwbBYloeUe02kcFKEnXnW3V/Gd
o9ww8R4wbFxTzzz1cJ7hR0tifxKw9WbGbj9Xxcz0hfagB8eJ/WD2COqhwI9t18C2
V3HPu7AMFic5SSr9GJ6CBL7chilkB+Z5F+oSapvRlHbGNqx6GHoqQgriPPBVIBzP
tD/dy/uTkFl/PHANUbyvZfl+THLvh9ecckn2Kw0B03T2VDmvoVCuMH0TSNuerrOk
6y4m2jCQY+WpLC2GM5xnK8kloIeTbC3fyRxiuMOYKsELKsYWSC5kH+aLEjJBtRdI
0tkl1LP4C7SAM/j4kYc3GPP7RPVy9V6mO4e7flRxud1rMtfctguRRDW7sBRifLmh
HX8r5YC4WcM0O/ovg664kDne7LGj/qjGSST5IadiyCGx9jYF9AwKERgDT3PMZIIq
mzkBYEruhrCRcbcPmpt+06mCqXs/jNVCoRTX029MmGBLQUrN/1opJNFGvYhdMpkw
UYHmemA9WaU8DW40J8sVaL/p6CEqVssoBRC+lps2Uxynigb7xKw8mvx7NVYtgTYm
ZTRv1DtkHRtREKp5EIizPfXOvHp1YnURzc3uEfMIxNDEq4TL/spLI1Wv8Y7irlft
NB6wB6SUCgiP2SNH3uXhojtZjMWWgEm7AKYzqQxJtZLTCJVOtl8/HRLdDYk5cyv9
zwYzmB6LkGXhIiURZxYhjvbJVeOdxpURMTO1bGn2KrkVFnKKB6Xh6JBJLULOsJL/
XLFD6aCB0oIL2Dhxp55DPzeGVh9RJs+hkI0q4Fg8/A66mF9+cQ5yuhrJ6M7YFkZA
z49z84E5CtiP3w3IhEM888YXGYH6kFD73yEBWrG8PiWTYA+mNfoZnFeK4dpBds36
2k1HkdWrKwsTYSLX9KQR8HnA+D62K6z2Av1WHUZyOA+324a3w8Wl3zfFowgVXYnx
zFOcoEgTJwjtDg7V8XzhkCxzFmJd3BNno8qIX6S/zAPKOO5c7gpK3f1MCCbE21x7
b8pYKk/o+c5ltAF6zX5plZoBa7ivlSNWpUyc8R74+LfK5RDCvv/rNX6RcSyjHdDW
OY0yp2p8t6XvzUF8EoD1uj0fQyz2f2/4GFpTkanwIffwMajReRWn26DlG60Sqv/X
cklxzIJsZW9nyGWkN4r15QDo3HFVY/+2cxIY+MBrpjS1M4U6DjjMeQ+PwfPxwCGC
WKrF0PiiOa5k4fvXewyz3uD3tPbXdnfBFfByzb66O8IjYNFFkvZRTbpRZBV0dJW0
LdctqJ+MdfgTjqzyMr8rn27kd6/IKSGso5xRYMA28shHF0Jho8sBtCYOgTPZCX0P
j+ZjBo/ykr0knPS5IizJuokWsx3El/Wygov+y1arKexBuCvch1pZh66p0YYKVb+P
BQpKxJcOAcFyZfpj9MGnrV6jqAqW/U4fMJEkkR4Cwt3pSlN1KxAMbOE1jrhVMkSz
C3DR/WHn+EYpR0N1Kudk31fu828NqUP6f0QjBiKpwY5/5qMAIxcb5UDbHvu/tWDv
jHipRgcDRo+P47a36repa/9z7bQLprz6yK/LELG1W0xvV0fQIlvced/A0JxwwazS
H/ahj3ZSC04Ghox9zSmrqToLV7t739N0n/RcC1edynbZnH6+i//SYe26HKTgrE0R
ETroyiCzWG6GCiyqqaTJfcBLO59nY26nBFmxZUdGDCU9qDjeXTV44I5+lMm93eyy
/dQuxQ8rE5uvcVv3Qxh2QRS0ssJ1kkIhROomarKddmSsAjArexevW0ICFI0WGiAA
sf/1jpQVKmBPCnd5LciYWi1YY1/95D+eQ2rg+AVHcc0BbPwPAQAN95WstMapab+4
3iuBH9AAISVcT5Ollitl8ivw8odrthO2mbbEg0WVSdyoZ4q3w8jRSPmZ1+hQtZeV
c1VlR04yJN4k8DAekMmK1ZId3h7+n7UitNlT/en0X6egpZQxht88EOmB2TCie6s3
4phch/m40TmHO6fiB/+NjA+SNGn0rs9JFF6DEcrKbpU6Gl0CM3+AHCy6+BHSxOG1
dZ/naVetOFVOSMQL54m5OrDjoyzLxmow39V+bYSF2cNLfSn85LcBVz95SaRMHKqJ
ZkVgoOG2CmqQVkdFOANvsmcsJriTEj+v6dEUXpOKuP2g81+2LuX0yfu9IG//+rPp
/T5LY5PHThT9qrQumV2u1qfh/tFB7oOInKIUtSlA21Bych1PMRMBvF0CJRcp65JU
5uKWN5jFZ5X/z8OT5i7QZiUTv4CPkShCrZWoMoAMt5qw/GNdCddQSj0rbvSf2Yje
kkpmeoTHPdgqpYn7j0Le4lmUrEosQ3MDdX6NZAme6Xx7lpYO2nf1U6HGJNflA1eG
Q7YSM0Phengs5l9AqI6vRJSpkOgemRdpOqOIsDW0IMDfI86eL4d8mYVRdKPUc807
1l+ppOgX5iGSM6W2pjoWFmh3CpUnXQcwoScvYw/Y/nD9B1P4gy7C+/wpt3pCJ2Ft
yRpScjYErVT/zvAuaex7cG5X81Wqsjsm2/WNzF/jm7qFSBOyPvaf0TsmnFcKTnkN
SYVLu4sLejPTSruQ8g/1CqSUlHuxeumLZfiGaCtzkYxrZIXdoQgZx1eb8dF7qmCy
vJ62cL6kaaWjGp1B0oNlTSE+i1Y7mb4VO2y379D7tri4i6VLHLJeRwnAMvsQZ/43
sFTIcMfRHQE0VsU2Rk3Lp737E0NMjQTr4dwSBef3KFNCyiKhhlcjx0VbmKa7Pi6q
PkZclhm8MeamA8HXzgrWzWCz9tMOGRXigJmajM3jEzCsV57ivuwbgknDwog5csvi
ewa4Q6XGc4DRl2xHF41Dg90e7s6eASKFhJWjO6LPBVtR2mTpKOguZL3dDCKuAZTW
ibQvnoBj4pkRFeyLEDl9/zlFHQ4PwLyCr+d5KCFbcEZoCAi5ZlPM0pkMinX3tDyb
dpAg8rEOY+XPPGZk+wBvO/Zehc49GlUsiRKuW/NLSXjEWxzuqjE4KZg7vCuNLMI9
9OB1gA/9kqIDE5SsfjFStm5UVpe4y1+EqWGVPXM5mAaZnSh1gmp/f0bUOJ6n22zE
2kakW9HOq7FCID8Xw1ylyWEdyCL7Kgyx4mP1KCW19d+j5gifYu4SanV82x2PnW2n
kgelOnoGsWWfS+1Pobev6zav0BwSrwiIMe4QrQoah/Fo0C+SaxuGbN566/7aIHjx
nknbhEnlgzt8UF/L/XF9fkh/in/I1ERUMAc22p3njbY+qj0007BoGprU72NltAqe
tRr0j608uDaGuuto78sF8drwi85e33XFpxxd+BKl3/BBrslWO1vgYNATQDKrsoVT
dIAsKroRD5tly8S+JrpvaZjJs8yELAadHu9GA4dAWh2aJuvZ/LYWflaaUiW+Mg16
fT8o0N9GemfzgHo+/c0fQYxbDY+lFryBa0P85B3an63T87qUUFgiH6l4/bQBUXnB
frCrZt9ZyQeUMDPgGtxWIoKeHt3pTM/Vr5J9grWpYdFdcldBts+e2mG5RuVcoQt4
LJjMaQlR2ejNDLpvbDzeuLwGcWn51l5bfXjXtVQ+R82Z0jN4jXeARg/JRVkx5DGQ
fVc6pV6jWS7eQeMv2pj0c03IwKmWc+H5zD2hhpyxnDgniF4S9o/tCOdQ+y+ui/jY
8iJRers9fVF8ajvWCO0EhPQMBYWtR2zVruwvpld5R7yDEoEI7tgNjcJmv3FrScsO
tGvnxZ4DXxx1XJ2eLUOHtM9DgeRlrYwU8ynxA19Zy/iwntJRYRd0GwI7oyixmNBb
vLaO31amQgGMeHS8kbSL9jiXGDFnJexbsqMoWbFiIbQmavXXvp2ozOr5EFXzZ3A3
xqqCX+ViX5lHy393+kjCvr7PQWZTt8XUGqWyxWhZXUr0gJ2I514YWu1H7z3OE3n2
C2jeayb+DyzsoPq9Fw/Dkh9KBbXRn5WQ7x6g61+WhEzUv7qySM/+CUI4lXHLs/sY
b8JH/HntMfn/kK5cJ99NXbaV6esunROUA7Q9nR84QpS6h7W1Mh/6ijDQmHdu5RK/
Rqy8biR5oqZQK/0D0FYdUktJoG5PCIyTY0U6KfA6FnqkXZ1ue10XXEBx1dr6ldq6
QPW01hFOZE7lnRF6hgrrnWnvTewJ2N1X/QaamN/TxwlA59JZ5T9k+J6qnrhcIP56
JZoAYhA7hk2PfZZ//Ln6aGYs5oSnPvAJ057pXG8BXlzQ2JEUXphf8VlhqkHLNuDH
cyPnVmN//oFFPDUFioCjMQPNTt7y/mn9WZgYN8toYS1ceW1DwWWZWfbWxXSlFI/M
Q2ld+V5PvaOJLofg/OnyTsuELf6uBN7b84PcoHNDqSU4PyWk5CHJmTUBHLVPHuex
0YAEZvR/dIDmXawkyBxZIubZypaS/cjiI9BH9A7ZWoBwMbuDkIvyEQuKQwQgIdpG
ymUh1ji44JA+xMl7Kzqe+krehtRezAd0AjwNgEwYR37BQ/eLt6SVzx6N5nLHdaiD
xX6y4x6qTwU4Y74jNfQ3a2H3bhksl1emMbHFDlD8E3Mw8H8yESQf8gfNhcQwohnN
NXXlkZFSqrkonT9Zzw9z9mJDDd/NVN6o3LbW0xiJNABH0iXEMPnD9fdZpgniUGr+
YCA6HVcrYK60RIPzDEIB/yIgubpAk4fUEUaRO5EBmwEb+vyQQWLfsgKb+1OBDEdO
dQOd6U+fCmvT4HPm5S0ddm5IibfQNCgudTjd2AthoQxtJaDkVJu6d7gzzdqa84nK
7yhnsJNHz2X4oirrrxdKprbTYAkQyysEsvLTVEz8Favhzoiz5E7LeWeUevASAk6h
VHvhCiBEseZxuFaKKveo5dlimDaLn6oLHdmNZrYTJe2lph60nwY5Wr0G6MUtN/me
cb4smFXB4yNS95MCxcfYZgyNbjgzXz2ZxEp93/8ETyM0FRtiZ86Yy9tR7UkeZ0Dj
fqmYccqtSm7vJON89n3AsgTj5V0E/t9UNH5pWrNc8dqrAkGMW1B+ycNHdFCAs0ex
+rNdI3Im86PjiCV3q7a8YIx+cWRaFRY/Jq/A8V8BsWkmTvFiu9FaBjzwfLojaYrr
1/16g+/ucYtNrpQsOig1/ij5Mi3UkVVMnxAugHK+Ue9fyNX2bXugmumac5Kkn4YM
Dox45QW9/LwVtncZRwzhF62P+DEW//iFAchyB8js9fzFvjDzqZjd/y3wbeBpyua4
CYwB5ViGv0LRQpsVREfNGApU7JCDFvQOU7TOfUdsc8drk0wxWFmzO1tsYNfYyvF3
v5YeyXvsyxq+woo1nsHxTHKyOC9Jvf5/7YRfsGyCHXq7ZfLnP1DnTzQyvQmnxitR
OdMbieHBhhUGBR6xa8mH0bb1zmS6lPGLu/iaIqrIyDJbWC6YhdwMcQFypKWYS2we
blUa6vqBqcC98RJJ2tnytEuKej+y9bG/t4cB9SMl7qVcE96aOXhG5hgmm6IJzA5Z
VewLE67Jajsbg22k2cYXQqop7U633P+EorQHttW0YWKb5m4WA+Z6HrhTF7DzRaYX
yvmnMK798EGNtaoR0hNJ2H/U4UBFrrBwQHpD3RKkdPTZ+x+qnARvjnVap99xeuiU
tcVzfMgMvnUsADJzJZMxlw0IbF0QsMdGOB9bXC/R7qjqAi3zeE7QllPeZahe2B1k
mJvcQaHtflhP+SPMNSJan4umazTN6GKDZwGyIkV4pYQMA+mRjwcOKOII6z55Qadc
jwtkhmLZ6+3ZlKV/pVLcefm8pzFqEPlJyAb37uTtgg2sIgPIVJKj7p7LmnoO30Zj
h1pTJjwso5WW1OE7fFsbMnbd20ULcA69SdnwjWTmWkgOxILhNOpzxuxy/VE0pzXL
Sx+xW1zONP/hRvZZPFLYkCRMVHtFNbU/PAwfvBPDNdKpgCgdDSk7xBO/qTP/rsbc
a3yjUzisdSWnd5b8JnC1hvirtXWPw8dNubBr13ildiKCZUgSzVW4RGg8113z2tk7
+MVN5vyYCIvld8k3abH7o8xJ1DkiNbw7dCBgPBQ9cmBJvyknbqHvbNsaMpPx0Muu
r/uKZIpjZ8G6CFtP4uBe+JhDfZZwxFSVcMs/m2jtSZFjzPGfrYes3XydM/v1IdU+
xt7NrLapTe8qlOg9ScsGI1NpbIGr/vHdxe9HBssOLCMjn0A5X5mraPqtQ1FcOAY3
rMTZDJcy4rPbFZxPcvJapZTJNvLZmD85tGPY8CORoTLpJI7X9t6aJ0QYFdSAau8U
CQVC7+5+khz1wzzzmQ4pZmpFsxF9eE9Wv/PDyqd5FqBMlLYHFdhwSUHwe/wB0o3p
XaBokQtyRA5hHXY5wDf2sWI3EXRSeGvmPfHuBeFY0q0DIkfNGOtsRSIhQZnPy78Z
SpDk1KKGS+To91ySVNJkEVimJJ0dHYQ5y3Kz0mCvA6jNmlQwOtzEn0B5bvAEv7aJ
S3u0WF1gfcunb68qI7Qlwe1vMlMAwWi6f//aOdgYq02qkYRivf/wkI50KYQOSlEI
QK8p+/GljKi8eu5UJ3e793GISfsG0oB//YTO097020NMpKF9YgFYnsHtTebwRhJZ
zLElAbMKg1MmEoyRAMdiOGtDK3fchyFPPGCeM9nutftCjNWbp8pantMgHsK/lIKW
gjTquZ4JbzIClgDfLAlAvZfsWO5C6kMji7Tazxc3B9brdr0LkX0heDbvi8zrCxyZ
fQ7LJJdtCkAqyBcu4dAeu9sH3rk1O/fNp/rtdauuvm8n98Q/ovxiSfMLk+xa+JUl
0o0FzcnyAVvKbkbGzXL2UNwCZFZ4HNFdC0mRMztHS804QgWM05vMYHrhW/nVMJea
U4/2y29Ig6zLKrsnounS8LIzYQaheqmewXEX0zF+ROcZx5nTelQnHOMedv8tcGeH
jrhpUj2PXp06UY4cs3q/yNNgswXFlg7+1J4uNw9bnp1h0Q8nt2X5AakPiDM7Ov6K
JhhUujhcsY6Kn+HcFUy2dz5SIy9lAWs9u6K/2BgBFaInAl2pyN9bcHDHQgbq/wfW
j/yIVqNMO3bKt8oje4h+pMha86Weq0ne9mU5u51+EKibj99krOXLvsLXNwP7qdtZ
Whpqu+WhVVTX7Pv+OnDfFN4qm7WFRzCViXSl+WNVHzEIDHJ1qrSIACNZk2tUZZ03
R/WRG+ntXsTsnc+hwKz8lEDRGD+NvHUpwIYGb7cUPjs6KyUk3w2lqLkHz/z5Xs6L
popeiueeSl2HaxuQoRwd9/wReGgCuCo6gPDa7DElWV2HffUM3lXrQ3Hf3FJUapX1
glNinFbwQ4Xl2MdA1H9Lj3HFRebJTycJPRwRT9rJZp8D8HCPkM8sE0/DJSziePAJ
fkBYe9g3SoOQ2TYtHWOZc6D2alALGfhl2ep9TJ7V7WXnaYCof3OAH3S1ULkeQ/yI
UH5GVVF0PG4cNvKYOi8rh9VtikNS29QHM6FDHew/l0tfVDGo8bJXEG0QTfA/4Vuj
F/SJZQ5+b+xwj01cXfvQBURRXh6jgjH+XIGKDjFCMQEdhYMH9laefv6xP4FnmMBG
OaReVFug7/2uzdCVlMtmcpS5QdL2kLxiiUO/UOQTsaCmobNjYbWAu5h5b5NfqeNZ
z1j+hRPlxOGkS5HzBG87qLjqYNSHOCLVodPKBMIi+LNO2ModtckkXbs3TW404pP/
uDdltnlMxTIC7iMoQoLFQ6t2GV1crMxzxAemPjbrc14B0CO7LDSX8VsUChbE6Ptj
uYTQtS/hxwZ78stVm8UvHHvZvd1fMF4YWm677DwQEgs1Dnpvnv6Jqy0PdcbjombQ
vT8UFqndEm1OViujJraQGlwYSNLEQ0IfQZYGvJnNtT8+7RkWgyMM5IgY4xRbsz7D
dwiU9ddexEZYLg2J04QJysgZi/vCWrCQeOEW9xfauM5dcNFLYHPQCCgyWhAMDPM1
FrUJsFb6PGnSyn9FYLSRp/ydJX/H2aZpPwPPgbKQztN7J8NLuRyB/edWnwbjYmgj
BYXFSVMnyPt14TsVXa67n4OSqeOvz3akSXjYHlUF2EbqxcQ3ifMRslw1dyEKY7zY
JFBYPnr+h3ZNn3E4iGGH6OfW1HYoApIBDnK/tK0UgKA8yUm4gv3si5PGTmG1u4Gj
iEPiMrt/60YUUY92vw1ByhmRniXoAwn+AJgtvl+I5coyFIzqVG6rk6PZ8ZcKbVX6
N8mdtNnLNYrZ0L1tPTwZS6UiHdjhUmnIcorVtotaPbc1qRb2Bt+5CtJubw2TlSIk
MG5YyXbYG/m6uXHwXRLmXgus5yYUXQOo7isVp6mcBUmLTduB1G/nyHvAUiuA0Ozz
FDIahrgLNdI8KYovIJMqdhOiXEfoMMf5Cdt+/Yt2TFTafKkDKsMlqMLH8i7eLepH
++PppihEutHRoMOf++iNkLPbtrYzkCeTz274EzBs3ICjtyy4zy+4eR5RrV7rQWI6
zcV9pDVNaOBCPqGKNQbyvy+fqFDwU6Vw6yLVt8urtiVE6FYEiNxbVJFluOUBAtmI
XDZbeJHQRAJOaDDRZLFyne8jsY4CtY7rBI0Q3E2337pT5h0U3Mt/yR0Mn9Mq3SoP
opDDMIeJyDKyRqwMyJQlr0bNx0jQtPSFKUBj+dfSdNCYeQoo0+SURyPnOM8uzwsu
WckpOvAhPdlMSjXOtp5qjGhbf1rzsVF04vCmFbaSlzTubKjvGXjqwDOyfluI47id
5gCIdMzrTFjl3dh5DaJNdDB8Kaslwu2TzIEjmsz5IPqkW/ENmaq6r8IkWnLgFrI8
ssnODO/LzByD7Cvf0M8x3Bod/ahjZ39v8pNgkXwn/3qPgAcqzp9Q1berl3G0MNFZ
zhxJH9wC6vRxoxAiu6TRw7/Lw35pV00c0DADuIcSYf5Fzf1Gg/MYKK0798ONIhel
d4Y4KFAHpNKxe3X7HIbZ2JLM+Q87vfh9klq9OWxcGTh9MjYuMQhIdTWcG+gqyLe+
Dl/KBHEnOypE/2K5c2JK7NHB9yttTXElc5Q1d3ODO1MPIIhGs4NRWB0GFhZcSBp8
31XOutl7akUqG0FQ+Tr/LOrV4klg9qtkCMa3EzEHBq2rWAU0f4F3b0zHKG6z7Hg1
upTvdel75tnfGvKsZWAiZPH8Sf1GqRGzv7apNzG0MoBFZR47coHKISnh+3iFr8fK
87TzpGEo0BwYJpFz1/cjR59+jwFS1QwpA3yQ41HIj9K7u3BhbI8HaJFBIbAbPGgr
0dVpB5HY199gSLoREQOZWdF4SYT0XKxJOuUcGrkVtJo=
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HopnTa/mSoS7wywrH5ULNp1/lNzOaoXM/Q5HU9hRFq/e6hCUGdUM8TAbigipLP+9
IWXheAhXRgAk/nYWH5Y8EuWZy0Dhdr4f/BJk5r0FcBQZ91FIUdTXiGWDcMGWdlMk
d7vHMCzEsrcyFehM0oPpm98u1NuP1LWabB+1FqR9nWEaoxMp+RQH9dRDn6300CIu
08nGuT1lGvnujMy3iTE6uY+DeTWUzwGRNqb7tWKGOJPCctT5dfAyIChESfs7EOS8
ycwViExbN0syXWJERa2+hWqjGuWgHrXSZ8D7XHv5WYK9TsIXI7VLXbw8ADRlCDUm
/RtracKsXfw52tN9ZM0fYQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5104 )
`pragma protect data_block
d63NiPduO6Ui3hWZgBgCIZsCgzHCFq1P6oyWNfJpbmpZPicUx7ZV0TnV1utIdIH5
CTZbCPbsHAeO0EY4lEuKcllSmS3CPEEMRpCCzi6h6nn1yVHf//ePBReXXZ9r3Lu4
/5eeTsTMF00M73V3zol8bexqdkDOsWTSQaWvLtx/oGlV2TS2t5X+C+jls9N7yBpo
zzXFj1LJaUElQ7+2MeLRSm1/M/R8wF+1yTAofoSr0pnp5mYLQZ6DfpztYu/UzSnD
TKy/3AU7zYmrZpdunHC7fP8mE41opJrk3/ykNbH4bswzs55oVPCLFcR/89JoMGYY
slQVBbupEEGsl+Dop640BAbdxDRuSRssPHJBPkRRyBmMxEidjnNiF2VkQhytTW1J
EKQO8n/O5wpiG+csH7DHUC3lYFGjlQ08Jd10vxo51kL4lc0FwvL2vXKx+rXLsTKR
XBL2cxYI5MYt1pLko6jD4FTb3kVfPwLXnHuXIZphCcG3HxecVzbVEZFZcpQ+ZXMd
J7yQvztILR3lLgPuSgLhd4Yp7f4cEwOMwa4aIFitaY1xRoSNGr0B/lLg/z/pXyoi
qtnn0tJOnB7ZaFMAoRAHSuejeGVRc/eu4C03gUK1LfZdzszePttQQnNWc4qyCjn9
wbMqBgsyF8R/iBi1xJFysjF9OEeHshEKhuMb1YnzbjfqFMGnAW2OW62ZjsbN7rIN
MZgOxkrRjgf6dei3w9Yng1SYcIthxHUrmhRAdG4H5t2Z7wTx8r8HLCQDa+qpEt1c
l6bPcbvQSdWjsx1ryAvsr7+A8ccf5YFoo3rTfYV/0fPGqJEV4rbOjYwuU0x/iYd5
bfzMPIqbHsq3BuOom+/i0AF557Wno8KC+gaIECPYssJuX4DBeRtKPHh2yakNnfja
z2BPXzfR1iRESIfatvgqrPRPkWW/MN9WLqk4o4styMF85O9Af6J7N1QZSF2vdHe8
4MJldfGZL8RzBFE9zxR2H4ilRaqwxKyJfAQq3huhb7GMkiMqUUcpmHpblfrFPMDU
kaSY744rGC3p3AuS13MLtw9wW/ZSgq7y0A08G6rvHfWw+6yyk311rqGoLDgBf2Vd
gRH7ByqDii68rZqd8JX2WXxqB+kmtVUl+G5yjHrmcIrd+ZhYU/Wvnc/BtahmnzUK
7FNxioW8JWDnR+4HLVHcnr1TGaDvZ/K8YmmZRbP1IncI+uugPB0/wnjcL32py4m5
6AkXVMKXgsBnSUHQM0l152cKLYjcy41UOXS056Lgt5GXaHvXQhKDstaK+vDejgHl
nY8e8g8E5mtOHICWqF8yjCmvQrU47pG9YjzFwV88r8Dk3A88qxb8H+E2SfK/36UE
ezl5Sr0H58Dbkr9HMMYQRmy9nWAzxwHwHQ6rVsI/KiZ5qAHFeU0bM4joG1vPAcr/
98b03onLCRTmhYO3au6VzsYFnsySTCJ+b3Bq9rxwu23TwLMeJksdrEV8ZZlqyRYc
byset/zqN27Apy1IaqUe2mb5DZ/NwzKkKGRYJzxeNo6cDZSf//eYGL7FvBrselpc
j3Ub5O04yoagYdP4p3H9VYiVnvwmWlA+ESneK6Kkx4fS+y816VDg4EJbr8OhWvEv
9lzM06/ZraYPl5wtt3VowYAY7w+EqgkWY2RxkhdeH08B5Ar0KrxalTjr9Jot/LeB
nXtS1PF8zzL7b8vXm169IQdgVEM7yZfmeXWmuHNCSplptDZ6VbEjkRivyMeHdYbi
r9539z8XH3U/nq3y7iDhSUKWqklPhoKI60hbahAbj5jU64rpqHyK2DaLAGiRSMM2
YpU1Ds6FPnGPNjXuF1O0zEvWMTpOunW1H+z4OrD8ocXaKl2tTIruSGrGN5oV2Nps
an90KC2Y/0MveKJBfG1uEA5O0exNkYAvxK2dh3lfBSQyoaTMqVxN0P5nZxLBKDJf
pN0GobHB2HIt+zVi1Bb+eBV1XhJUWiuN9BmdLBSwabTZd5/+qR0uhvPmnOubSMns
vk1k5a97SB/Aeka1Qo4cA2QnJD3CXAejgKr+6AvtPdmhH78bEa5vF87umih27bwK
VSWJY+8hn9Cp7aRrd24/X7HNknhoWwTftgVc6VGpxP0rKrmqB4LhDmOT3DkfN5qa
kKiZ7DS7uhu8YZXo6xE46LjeEpRYmAkt4pI95zA0Wux1QCufmiZ44a0ahRNrpdJ/
SfGX7/9FYEG5wf0qRThQltDv7acV9l/akBPVKZeVJewljN4v2mmI3cecx+bV/TKZ
3l9OHGPO5vlNDkiULbqJUkqBibB02csrD9ef91TM/sold7EkEjNv2K1DDvSJntTF
v7yvRVQJ/VzBuvvcEFgZHt64pvg1Jy/qLDBdq/eXF+cxkxROvTfEdChRsevJeZey
46fHLtqXczmyfspcNb0PHbfSl+yHfhKTbJfvWHAUKwOrmRUhacE2zStnIfxR4nj0
NhDTX4VAtr01CN4dOMl5xLdC4Zl8/9HPkfwlLH6U0AzlXxJq0OgkDBmx6MOtHXm7
n+EL1g+zCBdI/CYr1tSc9t9xIa8vvEMlxnHkZ91miFUje2FEgGNtmJdVxmPcvEVT
9V27RpuqVB+hGlbxvaetnsOy1VmiQiSpI31CTEF73Du2acL0lljUzxGwH0sJwuRX
xN7ncOPNAUlXlv4QFsmXPiCQ9bGjBcGMdoCpT6SRXdNGX0fWe98n+BIqM68098/A
YXia3T8qlMhVMBQxpadNoVSq1KPqQ2cEgDNl7C3v3If8iNVNO5vjaepjzq8afK7D
gEIm2QcW4boN6ShfCpjONMNY8laKX+DmdoZumWkf8gW14H0kiPr0y4x8CY1yVx5u
TSkWQJl8vYi0T9iU1dvvRP4tSgSL7a43tz39XdhHRPO+W3oTRkJwe2KmeJkV3Ghj
j5zAlAA0dwZ+tXMMf/Z+ZII3hN66nBW3BiHJFG+PVeq0BCW4pVuLor/Anw0+bkwS
OpkPQbrOdpoUsWr7OyWk6UV7iaQd6SZriZVEXkW2O3QrSNhw7f7H2DHR9UCXwiql
Bj3xO6WSrjfQwztwqwMhsCWwEOri+k57GaWJoH9mi4oVo4S2Pnrzy7YVlPSZEIwF
LrclJUWP09+DfMR9N8RCIokXMWZjNfkpp6B63y3ZN+9d9jVijE9S11YGC4KyKll4
FzHlEmBwkcV7jFKT47boOCEBP8AEEFLPlm0h2MOJDR/PmInso7qcLhuM8nKxILgi
d3J7MHry7IviAizamBH4Q4SaMbOujjroi/yV5vpVRi15L1JjcvZpkRx1P8JuZk70
lEDvA2/cnVh7xALEPHb5d8HeFbqVB0vnepFw31JiqOf5ATZO74DWQIFU+S6scBno
4vWHpi/iVsckyw3b5y4YapTDZAgzDNnk58HN/8dk40KbYHfy7LwJybqR+tIMBAcY
3/bGjaH5WQWNBI1MkuzZ9btbMbHPzWZ+AklUWV2S5tLjnGoo7YEYPJOY+vzpLJIh
cdRZpyVLlAQtwY5Kh640juyWY4iEur4tS0QPeyGIle0TsOWfAgTWDX5FwJ/bj6QF
kpfPSGr3gsoM/ZpnuE6om6WGyct0SsR64b2BSuiUPxcCIMTOrlkB3x723NHlYwrA
cM+XGaagCbsKgqRYzRn2UdXPkqdCrKFAyZzDqOArTA4sBIuWbsG09MtXgWrwdzmM
B3EKFi6B3TJjYMo2G9hJginNUY2Y636pxkj8f/HFiECjYL5UrUZPDTAM/jAErziL
gdVkdjjN5Wj8IMkBnRpnrv6FmQELsiCaAJQ5tUMTo7d9mExT61aK/qpXG2BNOgcO
erft72qK6cK3f5eRkFry6ibFf3k3itZr1BYifRAWSqcRqx5oYFZHRn9t71q/muLf
aQwxfSNJnbmfVIlZuSGFW3FvaPKCBpJxPOwuBJPDQMMw94FEJMFrI94uVhyBxdrP
3Ll/i8BShx9uRT+Tnhs2Wwvn2ZInxCsnUx3dAlAYLwS54UwqcDyhpMmsmAZR7iR3
jLpjlWbTfCNuuC8ODPexc56ZsAu9Xx1WQKejjeCmDsqacmx4uSTYnoQ6DcqL/tpA
/zycZaHfMM11llPzWX8CbPmvqNzwpKGkH3k2VbW65Ey2AzJxdtXgDX7Sga4IzdDm
N5fQYP15QA5fSE2iCDPcv7GFN0R0n56jcz/5lYMcBlOFO5vwS/zF5vyqfe3NM1xv
RK7LdrlO67I8bOW7xA6lqY6GVbSogm1CpkZs7X+wZFr82/BInd7UvakaW9E1pfqr
h2eS7mGThsbznTE8AEGJ9dnA/X8UVblcbs9sEHTecoXjRg+SVgBs8has8owUJzzT
JTzZWaYTpLrLIhXaNcsB8q6/aPV8b4X+GSKuNJN9QnTPeL0+Wtqr536UJuuvVZ4b
UQp+E3kdr3v9XF6PWPSFFRHufKLR2JA108q7O00GImFUyKWwvwL2RTOysYgUDyZc
VmPE2IESLK3FvRbyNF51yK8YwRltQZhprPUvolSonKMsH2tmC2aNrK6U80zZVu/O
R/AOAWCMbPWzMQ7ssRc4/L2J/K0xs5Y4AQUHGWkVtb0ESzq8YLfZJEqzv0JGovd4
3pEI6dipEnKos0EKIxao06YcvmRxV1S5u5PQrHmV1PcZU+HUq4j1BUHdX+MJyKWn
z4ju5kMIxMtO2Xz5UQItYHEhvqfFPMrhPRVYue46/8thCmn8TmQFc0Mos3udg5oA
Z1xqHThDlcQ/YSqVeKS6kwKqksBwq9q26gQlqmrL2U+6m/KwFAv+XnSsmuL7FnNO
gi/j7dteFa8FkrGMYjOkhFqrPo8vUo6z48jp1nvrIpoLOtju/a/hIskMEqAZjiAR
egGQVfq7ZaUXdd+AQRXv0TtSCrgKk5IzgmTai+lhbaoU9dsbRi6waFWNcLah2evG
5TAOXSgOQDZ14vaenkmvnL7Vc122X4Y4uJtnscb+3wWTS7/4u0+Q7liL4thtMvdg
/TxRg2K+yIHGRlMM19n1hKRJ9kA/Qd2svasEY8b9l24VM9AXcR/24WvG2jR+Jnah
D/OHoz/v6b7Mi62c5DEEHsJE3XKFLapNxBtLExBvwtxPDBbQohHq6Y11cRL3kNxm
+O7N4qzpQJTDWXd0nki8G02nS0rohSru//LN22eTh5YdkUOz79/xK+sXUpKftCro
wZypkcHtgpv6zSUZmdaGBvpf7ZRQXeQzPAsmDa/I1rEUoGXM3u6iEgt6/pceh0I6
HPynP0ErAxSNCjr7w1R2IzAJPeaGqDiRcI/KAvkeVUW7IqmM/I/4QmQ1mALcJ+mk
bf6ZxzHTIz6Hy74DyxPNSU4v5zN8Bqxv/1B0MTGqg8vU3RVRKUzcY6Rv1T0mF4GD
RQ4JvVNSD295zqh3qYT+jJuSfIZ/aBZzvGobE41uX0yWdoEiqVkXnkVUnYYPuBx5
M/9iHdgFlrl4/2b+BL6a8EOaXL66HBwd7jtiBHPvUt+nlKJUhvmSQwybsJZUubcq
hFq4Ar/y/TFO+REJTvz5MZNU83QylJx3YvvCkx2J0pW/6I6R8ywMMGoeI63sEI0o
L2k2f4Jz6mfDoN+hx7Mb0SFjp9VY/x63ZgdY6pcsSPZ3dqM3sDnmZbmOoPSSQVHi
qnMLjUVPPUzqIHNCCm3YLBTiKymiqu3m/IYYetLry6WRDeMmywtygyG+do5OoC+g
dSBTgRvD4dNYEcTsuyiD/R46z2DxapWWFAe7ywydreAlINUlkTGASeJuBQQxX8xQ
wa5nYT1LKH/EHp7E4MsiDraUp1EuiAdY1yPW0RmxXE0OZw8W3ovU0/zKKixAh7O3
vPV/EA197fkbpBF+iKEhmgQ/LovyKAN2rRXjMim+87M0It8yydj1JQJvEub8wYmp
3OWQuIFAkcbDEsQYTL4MgkehkygDYF2oA+0zx/cqEsNrcPIuT/B/+XK9F5vX26xv
0DZ2tfQS8BWcnodhMRUKGZZ5q3pAGVsO4uzYSgYxFIp7gDL6Ba4X8o66MV+iMHf6
xyD32uX08PznylZZph6ryqLZZWyUmIXtuh4Tz8/EsuIYbOSXBrCEhj2N+KxkWLpG
HpTtqEj24HZlh6Q/z1oK0zxUPnW4y8eKGJmb6Lj69QO/KV7vfgijWULpFMCL+2FD
oXszw7qBHS2G+5W4u/4Y32XkbD8P0T9QPd/ef2h5XlwUk+nZqj4fOxPBcWFiW6ly
DTNp1FrB2e3atWRndsvTFd6ib5/V0ncEF1ACBvPMwoylozupWo6k2xoUWnRyE+yY
KiubBIMu/IaZg0ZVCA9eAuNQf78EhYcWPnW35LVpVK3QKpP+7E/8H9DB8lZq/jQD
ze6Mt9sZA+QtJlcP96oQcyYqQmio1jOf8qg2cq/ojRAgfqzDJ9IE2qfTAQLLMJz0
xjp+WQjMzD8HX3u5+nt0gHE7mOdL7GHftCvQ0ICkZP8rCs0XegbYwZMSEI8s1Lh5
2TW1lVHNfWlztye/O3YXmcRgHHcNlmv/76p8tvvkQ6YW0FfI6ORT82uzJ7/T4R+T
RKKI4AMdOCvpI5XENeETrWl4QiOggk6PtTRhCR0zkpJhkrKIpHy3557fz5LAcOYk
+XAauTTDU/EkaEtEf+3QZT3b7kHRWPRznEBMxaK7FvFOPhpsN/4fyyo4QiPXgX8C
FsKfeFmoRES4Af/X7HQzlZ5YzU1Wzsw1Ch4QsJzKVoiH5/RNL9VT4Dg3+xcOgRr4
zjO80u0UrJUDBb4kwwcx3eh+j+Rc6bypCE/FA5dkAffYHmUDPJMcKB0jOxEnNUW2
bCJpzGkGbakU7vGyMrt+RT7l7xab+25+hdpQmWKH/ZgBLAD8jAnw0kuOjTk1G15K
hyC56kdXgYGs0+jXk4S0dw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gzllWmuzuqtRfjC/5yJ6uWB4ahZCCqofsyeQs99+MsNtJqF2Iil/AHFFNeiaZBHd
8tHTHFGAPKQOD77jaZIExvtuQwUZShGPuyqHGgGpXwVa2OhJd+3Xv/lz/9hAIyRS
yYp2zbbfd/D/4x029es3/L9qWrqyXXk1ZrNR6Q6/CP/0Ji8lIgf+ACl+oovOwOOP
o51k634TtFrQ7o3OhL2xG0UjZv6ngo8y13fH36MilgcjD7S3E3GmHNums29m4WHY
qzoAu9gCgn5mEOxMPrKUe8x3qU4TIInQ/G1m0ZTYYMhUaPB+AAvoc4JiooSrz5xs
gqFZuHEYGh6FGqtzXsKVVA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2624 )
`pragma protect data_block
f1lSL2ax77cTb+hCsEuCg+ydzSqs2/b3sfFZzMHMf+k0Xv9/GHKzWT21mT2NqJLl
fK4Y4uvEyluZsoxWXM/FSLOkErgB3Honn0WlvMhJYyM9rPrVLk8uk0sALn/mo72Q
gYI+9HolgrSj1aDWIYy8oUPRSNfiLdlpkd1swWnyPEYIjGwCSI4MR/a+f7ESRvrm
syCdLEY+mP14lHYEz4NNUFK0vcMSG5N5n9eMxyyNa57R+u8dq1QQKGGha8cXR/ce
GCP8tgwvav8gXHGjBiEK291XOG9JrnR5T+nqB5drrOJLBDNgcD1nAaEizplc3sx5
X66cZmJaRUtRe5j1ejaQnDiUFBuSAwNqERxYFSPQl5VcAAFqqkF8zrRzkzKsFrf3
KLka8fl78fBWl4s0CruJ078Zmcv8DN2EfmmZecn92jMPWpjNqD/zoSH4pb/fTdj+
OkcvXY4X1jX42pjES87dOzpYKyC6fMff7k/5tan6KzFq5aTgsGB0tOi0xnjS8hal
+jctRsJ1BVocipOkUxRik3XpTUv+iwrJDn+gnESWhBZVzmEd10KfX2dAOtbL4Sin
R3uyhCRnyGNS12meduoJrZ1ILsYmCkwjR7p4fJ7Yt5V3kXhxd4khM01zZw35ZUrH
E+b4inNLbYVdd6oqkw4A5jQPCqX5OCGHOJ8v8kDUDO+VFMPN7s0L/gyYF1X5eRTI
vYiopUyl0z7Kd1Q/p085HUHE8Zb0ZvI87P1dUcxfdtO0qR7zSCEX4BY9ijto89Kq
tmqPfHGlz7C4fTC0BtwoRSDEuFMGP3M4WFTsrDaD976zKFWLhrX9duVlo1zZixNa
EwxzpPPRtjgS+UtQ1AjPwHYgUzCTXEG3Ejf7O2NAeAcauCWC1vMwqLiL2o8y/S4d
IfpcHOHKe+zY3UFaOI6btOp+z+2Gm+bixOUYtVbr/BrscF2oWPrYlAVrAYz4BlLW
KpMSmiq49W5yQlW65/Rc1A+mkItluRt7h6bJWj9bBdA3dh6oyuRvSgEjen+20sB1
zzYloaFxFoAne9IIFBAJWx0GHlwfLHqfJoFmcExIJGQDG00PSCDeLTJWOAFDnc31
ilvDuh0R8sYgusfDbwiwOlGezSrMjvqm8PCmzbey0lxhKxO359gW2oynVmBux6uR
hgXBgA8TAAkl78ZmSXms1XM8MoKHdmTS+Q7nWBQuF6VTXj/fnGbze2GAMcyqecGL
/mtr0JJEhxHC8BHM2NuTtDboaZuJxe9CC2412uEP3RON0YfXUShCAHHQWDRrejfS
gErqu/bOXyNbdqc6qhYZ8Wlg5f/rtP9etNkMVWGFgvZJTZVOmrQMbsR1L900Txri
Dp7r/qJG9lNl5hJITK0kmgunldUOM/IE7cVi5YaAUN1XyvVFaTJi9UC0MhH8IqPK
rNPeZwR3RWA9ztJLH7UGqsU99Sp5v/UknTAZpQW0ZrGyiVwYpYGMn4ImSzveFSNr
AeQTkw6gmtJJJ316IRZJa/z9WBxm3wZtlxKN1NGVidqSnU4ZPb3Zn2yQG7ufcLNk
HdNN/Gw+JznAr0SRx+agnNXnoaCYprKfVQ+eNATlIgHMiVjTniBoQx9idAvORj1R
uLixSL8NLD353aD7YBOibd8hgF/jS0ITBK1fhNb29Vlp6V+ArBNlvuHULxw4yr3p
cT1YfN5bLySOWD9CVFs2Q4gx5S4n4OCz2fniZ1fAz/mvpf5F+xetvYHMwVTJKPxt
szGN8TYLArI4VgrMC4YJfn6MldmiLb6B54yhKQ6xdTARANAPw9w9zfoxvHfVyom4
N/uhvR9nR+cXRcB12CiH9FP8GVJC7Q4QEI6D9+asK6SJy1HM52eOo6nbSao5jafJ
6Zj00XKl83nFYwHkAuaqpe73FbLcA7v7MxjUECMRgOXueioVpiUY+yKttKIecH2z
w7lnbD5eO+8vtPDyZTY78rl/h+mI6/TtbbofEPAWCX9grWpc+JV9c/YV/Mce+65g
mqOc1LjSlV6bFlHNf8gZXZTjv7R6JUtRnFq2lH9nbTD1RbXXCX0NODhQhox83E/Q
XuWGojYS4nkk6kPSk9dMtIiGzxnurf7WAQpXzr8cabuPS6OTW15GcCTJqJv6pHTM
NIXdgSr5VhKpS5QIbx1qEjFPM+cni7gmM/e3ku9S1wJGLvHGH/HAKXFoIJ56WQfK
ejKJH8M3j7twUb4Fb95k/HLCoHYAwVZDNAWIC3raShQMm+3THVWnkL1UAM5fyJst
IDHjYidey7mfgaODIbzefg+PSIwPsrAfBBrEsqT+Tam9bQIDd0EihHuszNvGZe/7
tKWdLzkxzsm0RYfXhQ7fP1TVcga3kKd3kRULPJwVZhTgfRQ2nJyGaWGEOE+al6HN
4cOtxcFm9zVLCffVLOWbqVgC0ZHo010QydMYJrlJ07+XYc67RfQh1hGPC4fTB2tL
Cb9ZO+4y+oqJA8CptyBXpQsAm3LAU/SAGEK5iRc3LO4b0FbqqCKy6pgVtDXPLD4A
UhYHgL5aQ6TITcJ1JBSdBRAaZFudNFVSBSKv7+jzcpGhcmCSy7LeQ/RQRabc8slS
sRPTDl9JcoizA3G5kgtIjH/6ISBkW6aYHuOjlgRQbRAx0IEJElzgz7iYOQ4Loq5T
4pnXSruGwfhD7lXqpvliPY3Yn7Nb8vXoUmnvdsEG0tVkdtfIJunxyMRved5xATh+
ornxQCT9lc1ZRogGJKvjC+EXXNraaEC2Cr5M530xZd3LONkce/biB/WDgaybmGSo
ojj+OliEWh5nsycPawoVSdvJtGK+DD8Jz5lnjXYrSbtlnFaIDtciKeUVnCCs+Dph
Ewmc7/V2HMkTgYPREZWlYJhIuR93kTuGpTMFUDH+1XMjLnTEU3pSl79tPvkG2lYj
Utqmm5Hyb4Z1ekXHhoJnM1idaYdyglOKnqhY4bsHj81dRvuXnh0O2XiycAZQUA/k
85VNy519gT11LVLgyeNszQLCRjwHXWHwWir7qAONBPD2vPTfp6ITRcEIqP218uuv
PstqgidFaOsEL8wcXPdBmNW/LfFkNrkWqiiLP6QjPpvdhueEFOo/MUGMgKc7fTW2
FZK9o9iPYVDO21SH2yJ5Mz2zVzvQC0TwGwuhQrDf5Cna6rFoviMCIpHgDEE9JlM0
AcD1UkC6L3gEV9T7vn65+FXCG5VC66yI/Y1Kf1wLE26wgy1hyIpwwSP6PMTKime8
9FgBjS4ifEWkpjfDHJM8XLfK6rIMFiBfRJmIwA9DWr0VPlg5qsH1I7XwQD9vAirf
7jlJYrU6eEjiiDzr6NOioZLYjR/AI1yw+gAisHjWrKIPwzHFC4j75BpmwBhXO8d0
qsUMhKfGAxLfL97WWE2w401DCp/CyPLYbEFnADCHMAhw4Ar4FvVBspb3nP++8Hfp
upquZ4NRIUcMJEgo01mwWm2dutHwnGc+S44oCDmKcjNqvAJ1buo+1ZqcbHH+lodx
DSD9fR1GXrfkgC3Z2SZjjf2s77kpqFVOC6JoBlMV/7I=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jeLPa6gNOE49JUIRyzl311R0Y4/eGMIkwxKOaj7yeugyJRfdze+jSL/027cNpea3
wa55W8jH40/kXr6CPrcG5Lw3eE5YGcY6ddDsCG9snjOjOriAoMoquFNJbxSTO42i
IzcOhQWvttSa1wGzWQIqZjAyewd8/ueLSQjvxKbnlgIPHvdNkRVndLJeMRVNTULZ
UR+Gln9vSvJOqUVvf+q53yzL2OitRek9vPFN5p9nlKztb2qaqn+atbe4tZn98s/z
HYqkWWFHbIkekt9WS88qDN9U40LoZEvaKeDRqovq6zGQ4i5qFAmluO9tkQ8y5gwZ
SFwE/buNsz/P3602GkPyqA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17824 )
`pragma protect data_block
2fzUhf1ocfyNhUqH4/ov6+XQ50H93zjMXEKAIgXS2ZRjVRQXkX+w83aiGwZoQMLH
g+dslf5pJzwzoueBBOulmsoX4kAgg7K+kmHEC8md6GXDTSotiQAyddkd3dYOOjJb
37GaM3U4yY+q6bBdD5hfe9/M1nSMM0Emq+WCRBu0SgWSpZ3T/lET4JI+EexWttGa
OfIS4FPDDOmSZzfbCQWuZLrXE0Bou3dw7HXeHLvF2EjjPKKqD7HrtJNJYvXzCDA8
MCHFuUX29z8MSa6u8mAfnow67kMOvg4gIZQ+cu96Buu/U1R3z3upWtqCjLIFCnsV
6WL549ZA9uzKJN+kX8ZFqQzeN72sbm6N7MkKUGBet0OgtjJ/A6JrCmCXpXZBIs6D
lJ7T+mrT5jYEpWHk67CO49SHglOn9iuGA2sYTmS7WGGUF+YzdsYMn04k0M6p0jQi
6yXTym9XTLWvL4vlXzAUmL8StZEFXOvfTh2YQs4/rNI+ZCira65cLgtznyyNLqOS
JHIwqdQxOFJDy+ioyKnYKDqTHdjt4Zq7cngzgQuuFLoS39JRIWwR/Lf1z2qgip0n
KYFq1nCz0sdO2QjfneZLsGR+HFqVqyLbDGG8x6ihKug8shozjAiLWgy2alTyQ1/6
dggg3aF/EEmeNE8i+7aeHpgHiAQW33Kf32s6X629piYQDAsCb0RReS92E3ccK9Zr
XySphc8nv1/nEn3dirG+j+Ga/zd9Jb78824QsE54QJHLwJmzHbOnhsmr3HgscNvy
ipHgeS77MrBycb9Q3s9yfHZkeeUUuxUWtdTScy1Q91tUHbeZ2clsCQgLM0BCX3m9
QvS9WIYjKWR8Nlpe9HKKlRiStTfkdW2LXKqirIONFiKkqvo+Ba6aAnAwskxc3ItD
GznXC222RI2B+/gAOL/mjT6p4cMTtJiLnAzzRsoB/AY1j2sMZHQSJuq7vANJMT23
1iKvmZOZsi3SrdMTl+wSzQt5gpOflCGXs4m8EywfS50QwK+kuqo4ZVHeqm21eKF3
B8F07bEnDrRFnQN9oJd1hyPOp5poub0acXOvgPYaSqjkbcFB9Sstw56+CfNWEVVY
OUV1c6MtfePRn/kqzbqsgctMKLtOc2waGQDJDN5x3Nrl5IX2UyIlPt+zo8vhmhrl
N63YxAsBbe4dej1fj0ygdZKfFgyXtT0puUKaIexgt8LnC10liklSqND/aGz5LYaU
s9JjYNBq8ihbmra+wnlsQRDZavRwMo4b0MHg8fQWfiGbVOSwjfmpmNtfTLpiTef/
4eYVowXIfNpu/TLU+vJOm+2jkmkcP66HYfwUprFAjgWt/lyqtrM7DPjwUqsmpVah
Y7mmW/N9fYZ3H3yFmm7GdoUQwXQJ+YfJImzMLGa74lNLuHqpNyEXmgIqmGfmCeUf
XEENLRHcg7HEWD8ajBI9WUW1weTufHKVyeKW9tLRfxIroyvikmMcK69eyZ1zW1bQ
sVtEAp04stWr/Jlm1mKM6TpALrcy2lw2b34JTKxHl8JdnmJS/xm6ZanXwR7bgR16
Y1Wkg/scdYjbs1/Rbv+w+d+PVCKx948kxZCPDugHGhk4V/xJdrLcWk7GUF0Hbc2h
jIN3hqZn1L2RMB5SrGhhmoHtt1j38F530s7DJx/MnRbCAzKSX36/rctUr7/S2jKy
DvL04zVV1S/T5EaJ1Ojgflr1flBD1D6MDsC9TS/Pt+yr7kTPW3Lb8cozS52K8BNz
QnaQTWUC8fNR56NQKFA1JfXt4JJLZEYdVD9onDcED1hWb+CyBMlG2wXHwWd25Gid
ah+/0d+UBKAEzf5a7llWJbGk9496zM0+ijX2KcIpUbEQJ0RPUAEPHOolPqK9/eIk
9uxW2/SnxTjZ0d94JUMkqIUIYRtpIQnQPnyq1DLyaCXMnVs9WpyMinwB8j6ErNLj
iiewXl4hLQJAH8s4T2TtYUroBq5pwSXeI4zZt7/K5wKLN/zj4A6Uf7scNL84f0u1
mngbN8JlvmuPPG6gEvEW1WrVR8s4b3RQrniLFIybmbrDkwmJmusBszPA0pXlfN2P
t1nVKn85I9g+kje4XAX75XcSXtFjdRYQLxQ8wWGG+Ys8nkmiKGMP+Mpq+e1Mvc1O
Lscuci17I/xAOUJTfkzdFPEKjLklO75bj6hxAvhHQ2ZsZRVENYA7SJcskWABL0qZ
AwqcATp0vzlKf0j5hQmf03vHbZ4OolYTS22aURYKFyWTbM0HbRkABRcP4t8zWD/+
vptPRexFxnULvMoewCkZccYbN50s9cGPZen9VdfzCy278VdokqFiGqpPB943nQ7O
5LDufmWOUQyBJi2+hjzLDEWh+8beYeB/sZtenrljZ9RtLCYneDcDZ5QgdYag5c9p
0EuBRQb0KhhEFioZM4BST/ilC3MC5YNEXkU1Bt+Mv/AWUkGvTO3ebbxJMQkvTD51
8b/rRmYCkelpDb5iSuGNC5WGv4t6B6A4nuJGzwiqKws8F+MLVrN91t1PCJRvL6J+
H4+7bKbBrz5skvOH1jAWE8eRQ5OzuQiJOt3B3RVSwqxusrTPwmvYmW/xBU280jc2
mOA224qTMPYD3z4+YOmwTs/3S/bNqCjOfANRDOQR7keEiVJj9h90F+1xSkTOccM4
dNHaAIkT3NDJ2m2530xwfrJl7q6iYRJdfg6mAU9mdg1lKDYFmSkgqCs9YcAena/5
oQfa58+LYnLLTZT2kR3EENQWZpHRKF5McN/tCLI6TxrY3kg8PrTPDjoqp1rPxmJS
QodXARMi3L3jvoOav4oxiwa7KMTK1j7fwVWGhRsa0JauGMUdkGKzA0NYjehviviu
RF1dDECrlZTqKl/dwIkvXG80G+J1ZWL6qdqP5mBr+ujkUZMHCerpqpFog3mZLBod
5RfOMw9ojw5MqCptgjv04dsAu0FpOWme95Ds3tWiL8UnyeM4PpDppt8IzWbW7ynM
qx/Dx5aKeAEPMf6MA867QAh6/MUMEKWfJ3UwjPMP6i+qOlwjmYbP8yDeOwlHrpb0
hNW/R0X74XHePaMJ/FMMpHrtg2NKSzltra9HiZyAxNGfsEFEwp0OKVl4YZFf5aEg
XeKXePcZMrfFhNSUgemsXlTYJCFVF7S7fSk3Db6FOzSqGsaqenKmNcCU7pP63M/d
zYzvkZ3ELAQ5/bLnIZ/9Rjb7ewfKEZuxQB6UREcyxiBS5iYgIBAP1UTYa9IMrrm4
nOsCnj0oBxm/4X0IERmW8bAgac+cJZvIXKJC3Ym1l7/W6AugdWR5iF8hZ/nSBVed
2EsvBMgmAuZjG7ZKCkjvf3Kkq/JAe20IL6keZ/A1OOGTtRqK465inr36tgB2grWg
u5i5c++qtQkENmoNOtTBzTZrw7S5Y5DWo9fSniRoPUh+vu1X6N0fMTaJxAC5ft+p
GKYpokI+ieox2RPfWrvrmUnzbtS+svIM1GzBNXWDK9YKBFdrM/SHVGtgxB+KDvg3
h7AZalGcUWeR6FEIVJagon/mErNP3u2rlcUp+GLzR8P66HXz6qd5ZAJeaGLJdsCJ
iuUKKddZCIpYmaw5mj9S3SU9GBTUl0WIvKJfKqmYEMj88vSCTeEtsQwrKKCbDFw+
tgM3SdhuCGk2f+VcH2eMJYwTTtPtTCD18U6S5K3Kw1q73jLyLn07UBt3ofDO4Ool
zy6K9NQXDQ/hiRGE0fgXGOrlMdMosLnZ8lKRCSViPtUnIhvf3I0UVgQfDjMZeYv2
pV2sexJCLaQKA5SM7x46/tco7jTb1OiV7y7KVIdSqUjmQXQre0jeNTOp4vIHoeTn
iGf39xeFExAQBPdDlkES1dPO4djYrok3IXOemCRj9luc7qAFirnNg7Z5HjMFKtBr
r2CNaXp/F+P99ZOps7lTW1fjm8l4jOPb5A4+4dpxU0Y9zQcYm7X95PjCWxHjcCj1
XoOvOd/5MhfFLncL2EV9EzWR1m7udxbfBWUeBX4ev3rgGsLEXMtvCTSf4LGGyc/L
ZOz4W5+u9GIIK+GfwPX0lJXwbCUYq3MKExkHbGNi4AmNbfXVJ5jGhb3sgwwf0FIP
MyNNH352uW+YhQrEycq95nww3cxJrTItk+j3GZTERcxvUIIIDxTqdt1OnvRQtJ9D
uEM9TVrWzsb2515WWx/y6u1e7jgb9LFfm6XZXMk9Ufzf+OS1vQftD3S6q+0GKk+8
mwryO4LxCDDs8zzVONWqNhOYcCNAWTuzTtfRTxFcx4x6BDvPUKoV3zlIJCgurtkV
bH+KSmYP0tIjSb9m3RiH5ohkdMJF37f4EtJLpOtSWTj/js6kQKbuneg6xfZg73Kv
qq1pxnvVcY3elo9eOfXeP4s2EJzez6+Hfg6gjObVz5mC+STjI9sU/tpzXMTk4fQW
Vx6sFLcKJDByQfL4Uj07WqqH6uHRGBp6SDjaJOf0G8qic/G+qedzw+Ite0toqK32
b2nbrc7ZGhV4zkTcmPu7JEnLhNy6mzjRJz9gPQdjktz6OiTp37UYGOUDn2rQFatW
j7KOQKOyDhVCpxNupaxKqhEdbPCAbYtMwIxV8K7GiaAdAyTKSRvE83ysPKiMEOXI
OZAFi/ie/wERPpO3x0yAodgBSYbf9xpwU2f0ZLtHOKC5Nc15PGbFfwp98fhB99Br
uR1ihnpaHS8lvjkmicUsRO9eoPKldKtgaUPZLtjwFwm4tLyIxN76ng+cVtFRJwOI
SfChhOQLHnTwn4RvVMfQnfqcm2fDqpYGVyfXuS7SBFN+dVtzcjYGOd+o2A/MIteh
W7Dn6HPMZjfAUj/DPmskNqSFxzClCfggHaJNRaGKaybulQKtMcd79teC57apSw8Y
9IBLJiZFMHRbrrYyQclC7M7O0G9j2knHoR72O+IxPyLQwHgBFqjOy5BJBIUY8s3i
9WmJbScwtWsK67noqISp6pamNtEf6NFSbI7KH16uFXNvWXrMoMMDfBR3x73yPX2T
ywfGzdOtfe4wl4qlwdkkMIS2FGNMWhtumAJVRhJkTSiST0r39XTjbk6dTPeashAY
qclz6mU2UNTWhKsvB6nwyX35X1jQOxqHO82oKP2xXybjNIFPrvajrG3u3pWs+lEQ
EUJhZPqPqlrN1qX2rcUSlbCM2RDTRw7X8Ni0SotdAwqcCFCDBNr8dBh7oKlQgsaQ
WRQPAX92Ie21KBzFwzjQdQmgDohYDEmAZph+HnJw7u4+DiCY7O6j4Fq3KGqReW94
fenL2nNWQXzAH8Hgg5XnhpIsGjynN5xNVI5V2lUTWAq0NjEtkOk9gdcCWixrTbsb
4odsrU7V9LI/Bp2GkY9FDquhCAWhyQxh8zds6jZi/AWwgotFyjmpkTqEm3Ru8xHZ
meA0loP+QLavw1FEMLzgWTSyDnJRt147EANzLX/r1whAx6CcWD1sJu3yZljbBpDc
AbFEvFM+DkCeQYNNW4+pyaQyQq2zRjr+fWzmDyL/c6BVPyjV6NaumgPVZVSlOoNT
boCRFh/WP67whgE+GODuEswXlxKsIwa8S+wAqA2J3wi0jLdFkqDjKVpigJqewRuY
Z5pz3fYePgj6GL/5Dmp27J6ouYfF9BFbPsoawRqY33FsrlBdlvMsbEkO4Umi+vFi
aw8M+GSXTo2FcarIQ+eO9UHe0QGrxcaFioWAVzhwB8ZS82OM/YhCvOcu8Dw9wEOq
VDAH9rbfVm0WSZs9lNBRD6FZYVp68wFkj+/v2FsL/dNcmB3Xw5VMZqi2UOg5SIJ7
416JXAAH9CYQ5H2jteQl1opGmLCQCFKsOvo6venn4iWBg8BmTPK8q4pUP7VZ7v+I
HhxLQ9MQuAopZb7aYLzBuv67mhKy2YbLtnjTNg3ul3AEDPbuF3aS3O0mcSD4yF7h
XqQWKWFYwHyr9Ua6kxkqhfWxKK2vsbNGndlIrAe92F7f4QAkGWa5awFG9ZbtOg/l
Di9i3yQP7hy9BIMcs2061Ze97niw+D5kfzQqVi8eiDEDS0JrHaBhiXDuYd1EfErM
Zhz2ScFrYbQXwaQoJXB554xfGFdtUk15E0bRy1CyfdyeFY+RTotpSbKXOMvFxnwp
wJark5OUrUM2/mv+uSw98jCYzw64ADidQQHcnAB34jBhuXPUI5DAugV1eh7aVn92
LC3su+u2zyrWLNwFbvQL3z0GiM6yyj7t57luiTijGjt5QOPe3Vil+qxrlxOWMJqO
0BKjTl9hlftfRLGSuZlfaYh0r3/XmnYAfANOqkZgqt7njoK48wEdgxSLU4bxAn9b
pbGE3n0/2cCbyjHWqhh8MuaslqDd6Q/yAjM7EgXeH801s+LglsBLTRylQDrUFEHC
4v7dXoClvke5PN72xNqw46fJyH4qyH6nYrnu5yw3BiW5HLv90qEbnyGPFwlO2gG6
xEwX3HFcqDkb+n//iX2XaftNXFO1Xne1Zuf4WkZuDJdfwEhyApMMRQ7HL+XubWiy
NEPFq+AmfVk2G4e0FRzXDmoH0PBLKzuTRQncff/Cxd2RaXs7IXuO4a5v4XlEiXhu
38cTMRPDrE8VLyJKCx2562Fb+IkKDg2ZpXyjMtePxWeLAxl/T5zzQNjtLpr+1fOV
cq4DDsfspHzZ9i4OeOrXolZkJ912xlnEtZzemmMDwqXROgx8v8SjhUmvPUJUpbBd
qsWeD1wnoHlADm7sgkYp39oNykapCBacOVlu7+w83sSfvUevTRCqyUTOEqtjpeBZ
Hdf3ZpnfV6UccyvC2vgWyHQ14CQS/tOIz7OThWcr0S0d6jZN7aVlhTACHKHrjN0M
BNz9548LFQ6ZYw2v5XrlVuj0oSNMk3KgtQj3UtkDRnEWgTO1L8OD+LTJGVvDAbGi
u7niHZqnxivLzm5dE97wuOJEdFCXKacKfcNNC4Asv8zU5VmwiaRIEv1wX3sTCHuE
sO5t6x4VnbwYoUt57H+Nr1BiL/erf7xvpxmPkgHwPvPvuT9Qy3pZ8QZT7f5WVG1t
xLHAx5nYiF6fkOtsHe3UzVkELya/x0HXih8zWC8lyKQb0Yybjv8du5C3XRJ3P9DV
9jpX/zlOBm+8sjDRLRfsJZAF/WCCC20PrFFR7qr0OchX/rIOiUMIWf2FbCz1rzWv
zzOIdg7u558e7qKlXmkrmisnf+B6mdS6ES0XcyHlLls2anNHYtkjNm8b14aZeEKy
5Jgm2vytSpF+XrKJNGSDwOGog/+Khoft5Ci2fXOphdR4Rn2F7+ZofB5NIvpwoxbF
H7qpuVEzL9jXgwm4GnoV7vG3YcVTqCQEhGwho2OtH3oz0PHX4q7di5z+6/xn2JJo
zCjBSGnXd3GScG/hQoCWz8AyCys1fNOFeFqk3+SE308hcIH1prWf/Dn7dRatxx53
BUIpJSxPwgM2qekdXyMbpEhyFxyiSF4LcDSjhPbk5yXi5+1N+x323p+b9ssJ9wH0
AxoUSpE6tdTQmQ8XSaT8rew7wqpYvQH22SsOCq1Yarrrnid4vYtpNhuYHp2EY4Nd
GERMrEkkYpWN1lLqXzy7Yt6TL1nAexEdt73XuIGR/e3/LdEgLKt5tpa9YheYcvIp
naFUXWMe9OC/7IpA+HjBnadj4dqTUMrcdEyqYSPimGjIwmSfWPQKlYWzmSBRS1xV
cHbSeq+wsl9E9j8Vp1pKxa9MUYEXqIqlu8I62MqY2phcfOUzFcQ++DBv/rBZrFfF
1tUadfK+TdV3jzL/3DINkxldAbeikZWAbdY+n16B1EoMlZP1StnFBdgcpRhocO2O
fKlHFF6lVeU6uIQjdJn1aIABgh0cntcJSw1eYqREceF+qPnlYJ+D+e9eh6rFPZtX
aAkLcOGi548LEyLTx0XoQiKucTlBV7kd/OMk+WjCexdHkZJsOfRC2Q8YaYJw9Mkt
/mpVjzSqE6mPFBvKHCFrtJe25EzArYDYAXAaQESBMmolDIunxuZcC/gKJ4YnowDR
bhFvzHO+fKinzGhTNIe6lUfiubyvpSAcuDi7lPSfX1wNrQCl5n7cJSjJi1Ktc4f7
HpJ4/K7A69GeS7ZRUzpmuC/JUhEblLMBv/SQnMWytivJ9EtmG+kqRy5YEWNQ+3nZ
V1HrrJYfl0wmoRBZJkpjgRX6rwRt4mYH9kHwu+sHqWuKhiLx6mhi/or4GtRaV03Y
TELYqJV2KogbcmE7Vd1oPJapM0BLqXgwHA17UZDUxzX/rT8P0yiDfc46JMDmWh4k
U6A+ChL5DDabLzLKWVBjlQu0xN+qwxJJmGe50jiWiDZGGYhoyjZd/i0b/yQRfGKN
JVdRWdUBsAGGh/LpOWFsIYMbQ6/0SbAgPbPkSl9LrnLsLGXusQjUvqfYMHPUBpNp
znNrEzp9VRO8eamyoHQMk4uVP1BrVVjNSBpTGgc3+l3iFJKEwonyCxcmu0Yi1gaU
7pEHbhtw4Xy4plI+1wZRaVzJQ15PkYdV5mpBtgOv4IBiOn0jNesd/4GSrmrniB0C
19sftiPIM0dAIUtJbHcsih68Pe1H1e+5CAeqFiV7cSk6j9oWTmH685SfyyOoiM86
eDbsKdfncAqHcTtqxm98MNoVyC+Z0jdcjSq1rqEOALchVRiKm8Hw5+PwBJos+83M
82Pxqsct2OWpRMqlkjKkCrfKhFzV30mGWi1C5Smh5vzBUEElgj0f4PQ1nkTwGMgr
y5p1A7SUhrT/CHyE63njR0TTL/oj6Qx27VdG4qBKtDwl0vUx0NQxcznlZxmddoW1
5if6HQFubuEsqGJoMj8aLD+YmQFy0hbNvyCl3v0CMkesJdyyMxn92U2u/EhZeY+N
MHwUTlAgfnZOzA0lSbXqL8BgxbvzF6ddrUmxosMYKEcAuc+m/P9EzFMWXdGqa8j5
eafi7OTPIo8fGYZ/aoavED/rWi1MuhdwQNYBDOtoVDnYnmD3K0BnS/hhFzi+32fE
CIsHyqqvNi+TCWgh6ZcdGNrDRXwkI3ZSIqsqp0SEnrbRy8rxESNCHECMtE5+Zj+A
984oz/L5x3gtO2SQSHQ/SaHtmPna3PwcmW/mm3jEAnKMdi4TGITfhOQ16PwavL3I
UcvHiCE97yWq3o1k1AKUnSjvOSxZgfXlHe98XMIh0ELpY7LyjCqArYt/d7XVK7gn
wzfCFcvFnxmjPn0ZZbEVko42SVnwxkYC6Ji+NmYqlVeIM/kgcryiU7HwstRitpif
zaT0oK4YS1RBwoEwJSUA3ZfSz8XpR83jtq1iKaPeJ7FqjL4GJ353IeoDqgW+RxrK
jFOUEDFa7t8651PVx3Pouc6CLDVdYiuaY4vkGwyzQAydrHednwYdU2EYMJvxRokT
uYuVwrcy7VHtGue5V0qtN0Ek2lBMO6OZhrVIc0jaQnXhdvXg9umYDbe5imk72/eJ
vxWOpkcw9BZWCk6psZCmtcIujPa0bEWxoTsACQq+0rAuIke2ErwX3vABmpLm45vb
P95hxK4nA+YeYICOf7DHSHNchDxPcz0Y1FL3E+xfPPo1/ge2vAR0oJp9VtV8TUIo
KSkkw5XgDvkXUNi/LLhQSgMZbb9ppkFuE9giPr0aI4hrMUeH1lnrgboo3DlQF/ND
NOQIM0Hy5mF1e7KBTKAm2ZoDkiIJe6nVZivOPhTFHwksETGGu3yocNz7PLOgGcEN
ArfzGmKxNSbgdeHu2GaEp/gFaDLtldOFP2oTxYAeXCf8NBEVsfortj7apH0KESKq
61S0o0HF+XqwJmb87dGKuMsHEei0iLD4pQQVePF9JoGj3kfM+EhTkz0pJj1aXVhz
Qb1QqFEtS68V5xPfY1YpaaYBXSgS9IsdKPdBIT1nMcdztC1u3Uo77fqY63lVu5zr
xPXL/sTMWiL81JIzvjT1tFLmrAqd7R0VfOqXaNq9kQyicJA9AbfzeSDrPy/JJVjq
j6Ie+/3TCaOccQh1WJN59HPblFDQ2CH6QP6yZwlc65Se3pzDUIEg9evOSBsiXjP3
gbwnzPhHJ+3SMJy352NNUfEtKnJR/IvHuQoexLMKSbE+NWkLjCCTIu1Ub6dbP8tX
v2HOZHzkTbDFojy9RHH/pw3qKQzCUYvV85SeeJT2cGEn7TlEbVxLTlKy0Urx7S7k
l4MOxSAvmCRtx6LBJ8R/Q1hampuV3LyqEab0lCMYilw8LZ0QVB7vqbb+hHvLwvib
1f+IYdJ7OLjrthFhOLHJ1n2EaEoZVlRp+fe3DfPe0RE328pCRwsoyKCwfMM+DImr
tleSpzualL2wcZOmKPAqvkFLEr5LN1xomUan1AO4sVnjQXIKpilGgEX0/t3CoC0X
xDzqv6yRROcM6vjCfq6UE/tkiD76gXFmXD/CTVUJwsNeus0iNpd0/0/boBcXIrss
Vqr3u62ZzjRtgylU8gAcP6Kqh+dzWDsLMBmbn6XhiDEorZHS3FpTud/13E22zyem
US4gvAUwJh/qpSnrtbOIJYpkAeTIAICyfQEOP33CE1DI/TVVQXYeWBEoT103tiP1
ZtlWzmExuoiSnvtdWJcjgogow3hDMxDdkGkLHas1IWEGVy3wGIl8kwj5lfsH5bUJ
vhVuwIoVeJmuKSdyyGJ8C4SRiajgiQJ5F6RYj4lLt7ywsDhsH4ntv6/qcE2i/ZHx
E/9hW4Ltj7eFKR+ndfBCB93ckB6KIwwb4MHCwg5zQ8Nsdnd6bDBrcwgRqwtVcCLF
oJhRHDYpM/zwk1tzT711YIKA0Z2gLUKTKOh+/aVBg+rEVsLHxaFXECG+mxlN5YOy
3PR74OjZxGjizuhF+UG2bqWZYircOVzhKqoeRKBsHl8hFJGvDjI2n8zifq6zuENC
TeOx0erfqcSIpze7/Xbwt5M8FapNW2jTjbSSWoOaMemyCVb5Horw9q/oWOyabPL1
hDBJ7KyeCQCV5mnnaFXKv8BYgFNxdpftMjU0f3BVAByZKz7+gSScQcnM+AIkj0y9
gd385qDL6h/2VPkcRKuX6EcPCTGZ3ED2th+qWdnJxtiMqSUsRviPL2rHNCIWmpg3
9zQsGMEQ8jrEBHJ8Jquzad2yxwgE+5IoMoUU+UoUOtYRVfDDasDO9pCzDiW8j4J6
92DoNyXIxiCUSjj9zVOp2UxwOua8/SYEJHK6cfZ0/YxTMFsp0/TDd/79/AV9neuO
ylEfMSYkCXoQRWTMjsCQOo7Q1aoY9CxpP54pJcNIsASG0jVUmBXc9EYVqcAZjmmU
t0ttMEUo3EwoUJaxz/6+9DcnUeRduRE//SJapHsnHmfA2ZXaKQG79/8ghfyRhRKs
FcuAWabjEp9kRu7JAwNaoQAUE8w6JhDzQipUWq9zZeWxCsZnXAIddZ7ItcVaDfol
HlnD8CQhVj3CqupVjVqC8tR9t1O7NxMQn3xiy1LhbZm+1CLkKLaYjWL+kJCgFEdi
z/fmTtQu9TC//nlnJ5V3wmIxBKVxRiIALnw+/uAWb7b5gtD4LwDvu/bdvwub+EtP
6dt+hqi987E/JAqCgIggC8TrN9kezE0H9Wm0sR5fHTbclHdPlKcxn0zi8yeyOA6k
tFejKrTjGDNvnmOCuv0YHi8qPfdJft73Kd9Jti/UyRPhuDyjvCEu3Gi08IfNJ9oq
sv9gsaJnEXm6bu8CEfxfBKP490HJNEd2Ah5tH9m2lBhttalAx6YoyaG5tXeZHHBj
PBoxJVGa66hr0TFSLvPtuCHLWF4Q6cmn6fXIMliy6yX5XMbLF5mWbg+iiBXxp7BA
cV2Fj86Sz6d1qs3Av3A07s5hU/2ilnHIhkPMbT/VGnSshFPsRLgBMTykE+xLwpjT
1u0l38Ftsdqr5JuuKdB1LfMFFyZES4xrYcZenEER567sXCCGZSv/M+Hdj+ELK2qz
r0lCigoBppZZZDiGZZSAq/lduGr4MaBoSgikztRymlfkQQBRNEhSREbIJtmXcjtp
X0geYXG1PJYhsNArG2xBcWRVnqqxWPSX8ubi8XNMTnoEwyd2aBML2CeYBysTvQ9d
rxtFBRwUQpg+1sEaRAFP7SIzLbo8nFnKJuTqBPE7VLprY49xtSQUNy1yqAV8P4rT
7XB6KcW0T0M+ValUCJMR7wNUouPz/Bu15uzh5bjIRCBQkjPfxe5Kh/YBplYL93NW
e7Odm9hDgNWdWkFvXEU5lxOp0q1EZPnKr3xuVpSsjduUq1Epi696fPVgDalvYRNQ
hB3blTnnIXN9RL5CzAdcqtYcqAJ5tc6IySS5ymdPnl2kxGjbPE/lbzEusKALAFjO
avtyo2zUc/xY/UTC/5uEuMigiY+6dv6PnabwHIG8Dw1fUTc5FrlXnRIof3ZjryS3
QQ5ZG6ABEhRJ0qF6k4cB0o2ZSILngVnqX3cHjqigUvNY9A2JbAcof4F1Dm9znpmm
L8LTCK8uRR8GT0rf46Yz7ZNM++8oCLIPAxnRqajwD6FOCL+JTj7t8x9TcbiZUz3n
PZgyWsuaOqBH2Yvjj3PgFNRRMws9o5BPDjVL/pvH75J1BzrhlzPzUXE7qMcQGRmY
RQaOvaKLXxCVyz40arAynv+4nN7bWFcUWEuL7XHTd+myFqBz5AC4SVL8xv+ZAqAw
gSHg3qd+raQKoalJAMudpVAgRd4oogdLrtOShrlaEe+Ltm2TyWHSNwBg85lBgcgi
nnnBJQOQnFF2hb+RNMR0MhUvd49SnlnLkUKn2ZoeeWoU12Hi0QnsirODVz19AgM+
6oBJQKHJjLXA4zXR9o2Qk9VToxWcTQeu5UZr2MPbVJFNnkq2WGTUvCde72vIpilr
b91XGklEkBB4bDqc0CcDDCWrfYgZEdzCvnlcyL+X1uFob3UvYEXzssvQRl5j5QBG
Emu0iK5c6zncBXGCME0wlldp7EC5jWDxb8WS4HdcbVzJo54vXs25YAgv7IxnPj4Q
b5zwR15MqKhLdfUl4ambPpZE9X7lHfWhmqzIHUBPeMDwDnYU1ly5uRsYUVAp9ovx
BK912SPjvCifeZiCKI0POKi9qXBF+oxBvvr9KkFjUizXvqzEj7qHElsAM/MKZwq1
CBhmzBW+veMvn3oEkfaOk/E+A1DbtnSsj8qIafTEzLzxTWull/6Nkj544nhDw8Yh
KkxrjGiwbyW3hpi58r/BPrmcHTLZTkbIvU01XlczpVEHR0qQWj8YMPytJ7ZwrF2R
W1szKlV1GQi7GwDOJhvQORRP4xmveIl3cmLtFvyX+fUHEtQA7gbfvnMAX2YBrB6c
6AUsLR0flQhm14inh+ziHeufUsAo5fC1Tgv8veUn3QYd7b53WuQnrEmCGk6gE3mx
5GU1BxCchNys/J/NHi9Ixp3ELVvyxHXSteBnCT218BMmwWMICIDrPGkuNPusFWlq
lZSdqMwzCsQk9l2oqzhnv66F2MvWFs8zR8WhSNJpIExb3XlBbBUQvm2ppf1zyHO3
0xxUkMJWu4PlmvaGhPfQpAhKk1oaxRjxpEiwAtQq6sGUvABEAjVIm4PWqkMRNlp2
1JnDnj3w5I9RqGmEpvaoB2Bii/bQAohmCTAqPDV3YZdFaFfdkVbFfcZh5mxRhjbg
CihVRd6avzn1xyJeE+8zu7fFbfqVdzKANwUr88oqmmg20f9F2uO9ZgHqpM1msDX1
M1vUvxh2XCAiYuBab0zn6atwTpVy2cNZk0JXPkNMO4ESL9pl5j3mNpWHt1XjBuTy
7DGRCH87kVv2klFxXqHGHhdH9auDAw/61WvfrCdqQmbPU5bJvknfLuPlL3KWudXP
+rnsTau5oYWL5HwUhoI4iLtYlN/yqtZOXjbOcvfs3EzD1T2+++661KwVfs/kTEp+
DdSfiue18lue6Ym7Y33/9f8ID76Fq84UnVo7nmo6qtFbAeRVe0SE3rx0mnxJ5NMJ
X95TwOid5fImhQXEvjhzGMsXqa54b+pYl2PSRifdVETQmOHO6tbfBFE3An+ngP0P
N+5/das5GZPW7m0d4XGVMPq3pbj0l26KZu33Uv0mEFBsRi8IDJXjeDwndjkoMxVg
mNC0iqeZt/VQUytEtG813rcilhohDJJ0fr9n4MSWofduMbO0dOHtpPMICmS4fcjC
oAEUDWb7WzY/923kd5o4LKDcgs1aUeYQDPgaXEZCa7Lcers55RkNOqMe1SYpkcir
Jjm+4zbK+/yCvRgHwCxeaRPUPKUESQTy0owHR0ypaiY+FGUGTtQWPvLn8kRCdTOH
AkqjeMVuEj9N5zYKk64BLijwcSfhZVzGDSBy7EPKZiJ8Kd4xd/UvqzMt5Q/slnlE
Vmv1XIvo2jEGlA2g3BSD5PnWvQVPc7umvl2uIhujLz6srYs7+ofmBAQ5u/sRHFP2
J5NLARWD30icUIa/QtYUKP57vbP6+hLMDjcjAxOsvHw9yuhWTS+zmPccMerKwIa2
gj2Akiqhj6t8hDvFc3LJvMUmDhq/P/zIwvgkJBe/LQsf9//aGeBs0rjAknRrVzEl
ObQzL4YVP5TwllA9qhYvoNjRAsfa0OewphWJzmm/VLJsTerQ/1q8zKqeumZfPmk6
JVEPq1jNSXMd7uJyfz5JuVgV7Op/VJgqinTX7Gcn8xiwHHOy0nCnCrFGN2l8R6ek
RExfsn6liFLXasMwnMY8K+gszjpkvhg256LrinMr0beXR2BdHSy9Mx+03rZeH6Pg
eir/d0D8Au7OA+2kPy0D/tvQhSlMHxXJKoFEAx3dY085Hheivw9KojDJHJdQQo7y
/OtszVRuzSSQl5U7xK8m0pMdubEQgys52Gl8vzVVqTZZ7+DyaMO2yYs/5OKU2dp/
fhKhQuv/vKWopnQY7ryquJyoeuOxTWt6ivE0WTxPlvVkpGjMVNBpt6GPZDRmbbpd
XaVs6cF79C7FX5bTRIokxO646Yr/lqflx5p2cj8lbzPl8rhXjrGYGxKZI0YfZVFx
SpfO09ktsec90lyXmg4AZYJw7YdHs1nmxXpOCYfL6Ym65xdX69hwap2PvgtN2TXU
L0aWcso5y1h80BY/LoEyR4AC60Y8dqhMbS3ZUPjMVRaFr1jeJidgLRNyekn6tLta
Y7XYDL6vAEZavOzYFCXpxMNp1/2mIo2ylf5o5zVrXuIhUUc8J+g/rNU6E/LU5Ulc
fHWl2obM+a+ZfXvQwq7y12Yhs3KfWYDpJcW525JFOheru9rESzcRUU3AyplVZebA
maX0Enw8d3n8b73oUH0ZwCBJesqAaej1r3psDBs2Pg5/bPft/N+ipSAWgQpIbYxk
InSc+P2mPuGPmX1Q3kyKH+4P6LYdvro04TG1lejtH8qUqtJ54+4LdOZJ+E6xWpWu
bX4L94+HDSAQl0hCPzGtOtWTw9PoC7g3Rshe/sA5cR3QPrOwoyW3DsJ2g7Tb5Ybk
KUB4j6sC8lCckwQ/+5pMx85cjpNSPeZTMbCKvk0/etO4UlYmisAr82unXIJM5Iuq
wF2idMT6Z5enbHOJxKUCrJLrEL9TOnzswKOGq/5XAzJlRKruFlvRnMDTkirRzAU2
e0/s7iBHJGBSI2+jMMcTieRs4uH27dm+zEvHwvMS/uUY8fnC/0b74z5DtTbn3U1A
kkk26goDgY3rfTz6JUA4cYQNOjK6szHq2jyWWMIC/arBlNZYP2L6wDAjLjFl6Ruk
hJNlnA1VMWBl+ov9uNY0fBS1ELJWdEBx0hF2c6TKk3sbZeuKEWsJZLJEpAjNhi9J
HBNuhQ9BQLVVg1tSZ0Kd5EzNgcTYkNFNuMjeLZLlZT6uo0Qnt8kiD1zmwcG4+3eb
2S1vFy7ueFJ/012mcIimQ6HaFo5Fjb+2Q20lXOvXOeg1ysjrWagkzUYWhEkOpgeV
8coCWBshRq3J3l2aC0k9+6DiHEhbenHzPYHQJZGokBYuIVIDxdtuVA6EusitRjkm
3FAOuo4+M3bgo0HgCAvAe0GuCF/lFWdZTF0WR0OqvxoIBbfW69Sd6jjcJHvdq7Gd
u9cTNNoXNEq80clzK1LCXv4JVwNmCAp3fyUs+payEyRaBQJ/Tj9CAjU27eRLr3lq
9HXHMx4FAI0e6iruT1hT9u1AYaiFyKPZ7snDNht1DnAY90ycPQbVIJ7MHlTPr/5v
N6A9pocE32MhiNT7NHTLsypsv9dKSWIOHRMBSHKKsyNMjcGuZ1RjbPDsR/pFGBI4
PAzkJm/9G9cCDB3maJaX1DwSDV5krYM4v7evJhjO2l2tdrqdqJrsYsTBHVKC9VP2
fzp4R0pBpz3ZxSO1iLceWYLcPUjqD4CN/7m09kKUut4Y4TPLLlhNQNGNa9WNNAJA
PaUxIha966EzJ1m8gW74Qu9/VP+JQq3cFY678wks/YIM/oZDcuoXViQ6XzsyKKM5
+/uXWkHvzTHAj6xJHH0eKFJc3Lck3pqp4e1VymsIsdznhvF2gmVhdNRj8Tsbs10f
PUuhkACrHxJBr6Bbrdje54MfxDN0KcbwZ/I0XVbqjukui98rrt9vNfa62Tv259Xz
YtojbXS8GS2b6gMETDOFWgKxFopDSPI9tHPs0tNQR4W9MowEnubtH00jJ/CJZGMH
UgG+vBPWOD6YU02q98EPVqJ/hCcSekqv/5yCVvpaXg4UslDxGs0XNBcwcv2Yw2Y4
hRHSn53wXcbZVzGH9JIcxlBhqMYDQvAPHyd31p784qgkxNBg/UQBKFezNK0/OH3L
5sUkXRALALscvPqrw4m55hL4miReDFcn85xUvqWApuBRR03VUiqHJ9tMrmQ1EmCt
yNWUrGOtuJYMbGNzsSHnPAEcBBQQotFdgKmwK8CwOBJM56d62Ice+nPePCkzs/NI
rjQr2lnD6vCwLhCMU0x0JG+OFvotMdiTp9kdE2uoMziEc7wDudiUEWMi+lx1og/U
ajxZQa5Vpff0CuWEtBIgEZ0pK8JI02NURLRagb4MxD3inuTAFo1VUCL2IdGDC1/E
BimXG7CsZGLCRCliuk6IWUKNqdmTQzj990mo1Fz+6mEB5MoOMahMVQjNvBTL5yHa
QakghT75C1pa5HOJow8SA1kwKjC6H/I0e/Z2b9nbLzsxWigL7zXdxQkluBCDJ/Sn
bjNH5Pzg6dYNbkPTIUAnAApZZ0hVcvYjLr9cMYZM4Z9V6xKD7WVwJPrbQ/MXVrsR
EQG6CRK17w+e8Daoov8FNWKA8hh8DvzDSj8SKe3k5KF6S5C77I40JyRkBDiFkg4H
rfdNDhyuuEWzdtbKA91U+7VsCBpcU29w7aZJsiu8dPLStk1WVY91I5FQ+nh8F/Hl
fR6nfiPs/OhR0LQrolm4NBNFtgwnDGFOYOxsWOtQM8HtXOkNoKjL0tFueqNkGuPt
VyaanAhO1+a05xjgLDP0b5MgvMzCMaaHV+fbTb+70PnDiKb8moUIauvuVqlO4tCP
uwLs78c0c2U8FLqlPpuFpvEfRtfujHsMbLzXAN+V18VIjW7EY8XbQzn8TmQmE3NK
1Z7+SShamXZueD+mhYnr/DAS4w+ds3k9FqsvqdhBFVQu/8UgqYS5Q8D+hQbJNgLD
CdCTHaayNMn608qIpgCFnjiHYKp8xkJIBs2CieIchGVEKFldjg7EUXEr2brXgrU9
4JPwHZ27Y/DqKN37WP2feD/3sFEN5Xi1ujcQd5Qa0zdON8dZy795FPNeuUsy8n8X
6ExZ/Y///D5pLyQuoFxMIsX1asdZ8jjzZLcHt5Zke+k5ajpTYhNsi5unt8s09SHg
tEt0vQRQ6AopfEYMbsZ9e+x7Jq4OCZJjzat3OPZUpwF61fcAexPwkFWDz+ZT1yGo
etYCsO+s9WhvK4ga3q2Q05kDwtz2VdHvwnythhAV0UCzagejIXKoG0OQPAsD/niv
JT3P3pbft/qL1uvpWr8n6QuSbWkHIk/OFwRJsW7D1q1qn1cFGXF7XyRjK/1aF06Y
T8qlUVs52uYf1KtGN6Tt27ahdBmnbPCXEjCZsq4K2mFu5PNR/6PE/w9lRKKAqOhh
Uy4f1f2mmK0JNKzUZbCfOheYmlBHU5M7n/rID5NPV2wlXeO1oYQR6Q1hvBVK9w1z
Nwe5+F1Zut/+x0dRYtLkbf0DhuE5/X5mZcDyBu3Uo3frD/orZ8K1vS5P8VL6fBSS
IMEJ8IbnBrBJOZcpl9MalNjfMNVXGJgGzyv9APNgpyDFoMfoW+jifLxRBcq7R9xT
DlgJJho97BEVT4UfLtZauJCoGqEXOpKvy7tanU0HoztwsqP3B7VH5YDnvBwZRrBZ
8cXFOFHssjDebos5Rkxav0dscB8SGssDTBL8OHC7mGQtp7rdLbvb/pq4HuBJi4Tv
bUD8Fd5P48IemQgCHoKdUHnC5Kkpk1APbckD9lOShBpRdYqt4GhX28suJzj2bIna
2rQN4h1Bq5/WTjtjnE6UZzM1BecZ7x2UXGR8gMP/92IGyKNxpuPWhGC/LfwBwqU+
u/r0V05i8a6cwrnAIBiclOG5m1+/AEaYl036WO8PCENhf2v6qryQs4qBG1yvvI5u
eMUGyIGpypFX/5i+2mfKMOgPi2w5X3Gqr7sym9mCxsinNmI87PtdIUa3y5kqG09o
luC8TmwEASqiPxaFKs4NnnL0H6vJBG3GQwQQp06I3Fvidvqwe8oDAx968YTzKThU
Kb6EWBwlGzBKXXB/nQIlQ89lj/4Zda0UV2xBxnUCkDWXxM7xAEqvnxorUL7UzPA7
liDBOfx9XaH4lvpIjHeVcoGUVBiCyOFo80Qi+dNAl2tTgHqKOStq83H/tmDNfuWf
93gmqYHitRcekQHhYbhL/bePD9XkwvVmC78QbnsxHekInsX3g2q5yh4CEFKKcF7/
hSa8v2MfUprT46zzovDQopC9ZgAlRsTvgpuw9rPzvZDBkflsqGmWmQoS536VagUk
+k/q8IioLQfx+cyYh/qMMOPmxoNy25v5bBZNqHcBe5ZKXhEr8HGoBE3Sp9SMvGBn
qUs9fPu3FY1fl/lgOUdwMSBcg6Q6QIEafonIRtuKB8V7C0a0zGEdf4h9canaR0aN
VFhCtphO/dySlffgH/f7FsHgq984uXc4m+aRTDy90W71083mpn7q+9qJFJyav8os
XwrJP201L1Tqu+vs5HTzuANMljkRLPv80mvMbbKljwB2hoj1/OGu9qTspVK02CGx
K2FrnNamXAoU0YFDlCojIFYSiIMyOgCKBM5Y4Tgl1vAAlLUCvvKMu2jJPyfSKZ2Y
OgWmyXdPng5EthK/zu68gsE8K1QzFhyb/HJXtfVGkZhU3oHDa+7jP8MoE0OJy/1b
1yzAfFMvW4P8m2ov8nnSpoWHnILW/MghWjZ3K7eNB6jr9n+9P7d3jRjuMxTmCAp7
rrMu6vVINZYuBaCgAyflGOEHPVtzhlXxSgaZME1JgK6Y/tpKUc+gI6tlOn+Pcgzu
B2aStAAjtvqR5+JzK3BV17dhARFhl2H97ZiZiudHAvLy8n7Fw9RBniapojPncWmF
Y1YgC5GgYi0B6hXLLYJps15MNmQAppVICaeoTBxmY8tDLxdKGPmL5SL4bIHMYShg
dewZjVhhOFf4Vfoz05uIn9KKnZwnyB3cwbWMSWUCbvDfpxAh+H6qRkyvwYYRg4Bp
OjInXR47oXPJf3HbHQmGzDl01y1CP75xhglGor90ny4JPDM8jSv8UOd7y/yK2f1x
QKt3Ou2+I6uXO9zqXqKa4MM4d4yrMwsB82dm47ibmS+uDPZ6n83hhliW+W9fizdd
wylxqrA6mWr4H2jiK7jYjL+xWteBI5MJ0nur4GBriZ0tGD+4jqImIinQ4beDLyUm
tICxg8qVcMUaa7akid4RnUx/aXWBUsXNmS8hr2V9hNODX0hPUJSuZiYtyzDNANQU
ki9REg8cITR1vUTBwQTDsN0oPuqOOE6859bFE7VApEi02jcFbrSOXGgSj2jwCb5N
PLh9t1MJtGH8Vqe0ORy+hmkm0cy4vQJuRJ+m8Jszj0ydzqs2fBKGw75sf4JkfR79
dCKBnFUVCQZ5X65NCT5PaSO6AAOwXWv8bbAUPhMgpmrjC9CIAiK4n1165sdEPWih
jYcY5Y68gjHFlOtcck7/KzTiKijv3F7lCaNBf6u7JuGYwZQ8A7sZM8N3jNGvoyPR
0bjKrfvOEiphpqbru6CuJ14wAJ0OjCMbMgAtmyPVpTbvCG6nF7Gwb4Ma4fzlrWC4
VwYLBiu9orZgvEOt9wK4bB0Ha+OEluGaLQC6AusUICZTYV9VlcbjEUbGGL2Gk/E6
IFKDFBOZh6qqgW5UeZR6y45QIRYCVxq7Ify94U16MPf/QiRZ2XOCfD4Y6Nggd1Yr
k+9ajDlkakda+9dDx8cXc2sai9Mr7cMoQLVjjiIe4uolxs0zUTmOhDka7TKjlgcB
32XKeEAklW5Wge3UVZCCkw+tT9DFpNzcV1nvGmy4IYasFv/2heFTYVxAw0sq9QhQ
mde3y8wroQxv8aQaPHynVfVfUI35S7Q1qsYXTxfnuxun46BTGkHcY+vCP1WiHRxQ
v9H0wAGgkvXcTd/IQFXxtD7DhhBa71l4C5/nLCwwULG/L9XZoqvCybSpbpMmUZuE
fH9WwMIgYgJZZ+/4lBFABKxHSm+CYk6u2JHi6jJBioH4EC1/8buY4A38DSMx1prW
kRikeu0y640McNJXpBNRVI5XaC6ryh3sPnD3y+whXHZlfeN/TSi71LvosAO27xMy
h4pF+ozTn9B2GWupfzQhdscRHIF2FthDUz/Lis50PJYnPEXJ+BeEPuJwd3oZHcQP
gjEphu+G8xgaZIP8bluPDf3ztKSg1KkZ5I7D3Yn0e5zYh0b9jGbDkvFc9Uy1UbLz
b1gTlTXAINPy7D7/vi8CKSFpiVqZWU8u8x0yBfJjtlVbHOcPEvnxaXPdaQUbmhfF
yBqKun8OxyrKwW57/Hx+f+UXUiVYtwm0fPP1fO9iGKRTXPV8Zg1zYEpgx1ALpYAu
YwwzCNbHJW0a+LDWT5QfFYnoZIzMG/z5ckdzl8Z7qmbo/kV8KZjo5qDYRZQt9J1o
UC90oqbUFqr2JW2XWJWqZGUXaQKIH5jeI3vi15VK9BPyzySz2vulZSC3q5muwisR
MoWXuERDgcR8xhZeUZ8tAcPl1qfJcEEmM8DbTV8+Mut9zhA/YGvEZ/F2e++utSDZ
oGygApX/x9nJQg9K6QOlAk9E/IsWY0n3Q496DjNODAqS2PlzdkakHhO/HV8rcJEo
BjB84FWEtVvUxCjngx3YZahn2CBigHgM8cC5yN0CuJYDvLPmHyjZzuAk8YxRchx+
+5d5B6xO3vaUkNopU47GKaeroJ3JLQlS9tN8TEN6IXnb1TlVBf4qOn9rwTDiXwS+
zidjmfjQ8xxDmR+q7AjI3dTYXttgR4dUOVYYQSnEY64355NE0FAxK+yiwykwEgxi
5R8zK28wH4VfzpLlCOWaKhYIW/HJ2HsbtTS4wbEFqAyWIul06cB1mpTbEts8mXCj
zkxumYERyS/1xtzLfXSYtElZbiiII7Fi9piRYAkB77DNCqN4j/24WQzmJZmSo2Uf
PwwJh+v3wdJhyUxVwvW/QpBvlwoMzqL5SMjtor9HN6qZy9s+AprQywP6GU8CRtJg
sAeihDiAfFBFQnqo7TiSSpVPWorxDQBy5/NaPYc7LTvYzoBq8s+Ms4kGoJjP9oRY
OsU9vDb6IPvlE9htd64xD0h3G96YR3+fPvXRuvMqsaZ1otxDvH2bpwCPnYkLVQyo
2PWC5zNrKIWMPUhmseP8yx3OMPET2x/fGVCbLU88G9u7StzAm4wETI1ivyEyAGUx
mkT4bmolk2/gsx0XYmjDApxi3nYpb4xbXNJbPPI9LpzX+IE9/7rJq3DMplTpm5xQ
GAN+Cca+6aL0dHrwANcFUvdjmWIdOyhMCZcgNWSQXU09b9C+uOoBTpjJIWVsm2Z3
CZM/ifSM5lzr1WxW1GLUx/gi+h04R1vYZvWLG7OM8P/km0gmMrmgFyN2JsLtCUjh
fzAsT1B1q1pKDeO4OTZvSTZMiZtKeHoaosgBXAdh9wFMuAs2etoxGVtw5a8Js4Oh
YEOE+JVtmrli3JDFlDl0roMysk2B4s7jN30mujA0dVk3/dN/MChnaixXL24dYcch
wb8ST9Lj3KcbpUXLUkfMsG0M/gN1+8r6JsQKKMOzNBxK9mtqiyOlOtTk+wWwBqaz
xwLHZMNrFQAhlV09Z1IwQpoOSm085CGb71658MQnsoUWenggrDNe+Asdz0Ld6g4O
MZvhafJyDHnm3x2lpLafJgiwkUp2JzI36rEObSxikJ/I3Brb7a1kwF7XFayfP4hZ
SZ2FLg/h0XzStU/bBTjvjTDkfStxCL+FFSDewE6C+khvb6CoUsuMcmg5wMvUhIBV
higsjuz2+J6KKvM4mwUbzFN07Jkycl68YLP8LZrqql7Md+q9F9uBaQwQWx96JROF
2URhM3garI2QT9FqOIpEMXnd5bioSiwW+b4gR8KC205hKYIQLlqj9a7GVcgtx/Ef
9ikuO63nL+Zuu9TOgVr4kGkUdJZM6AgjGae90x5OrOjh2XogUBPwlwMpBH9NHA9W
OxgMHOLmg529NSgJ1Bm3OK37v/3NhjZc0S+5XvdE22aadmS1SMLMqVhs78qJ/8mx
D9mjlfv6eCZSLP8JOdcUHS8DejGeFg3aydLYhl4d3x/8axh0KnXBGR4POXHYwyjM
U8C//mMo882Z4X/1DIuucJXI3DNpgbIMUXdonSfnYY0vtntfYQj1A1vWy91WGdVY
mAEYYMG/Gw9bGerfHjRBb17qdnGC/C1RXASxi1dHoiBSNDYohdLT5GEVtywUMzZ7
3L+cn3KxGBLrl2lhTlXQRQjxivS3I2XblNBgUJ6a9uf0676FxDDcxSz++Y248aa6
TD/e4Ths55YzzJombKU5r+fAt0uVj7OOlBkBpBXbYFO2TrRUIm3HOg36FJ0WpvDR
291hMFJqfqdrX+0sOumnevwGSfqZAFxyyFq0pBllEWrG/QgN2BZLr+TITI/UVQTe
EAIZZKbExpcz5Sh0Q9/tTA6Ng16GuJ+dxl0GgTJU0Rpz5tGWfEv0dEkR/0aS5vqw
/1XYyjOIsiwxv0/LWyRwIXV+kfTR0VPbpWb8uls5f1SXs+Q1B+hES52yH5rToZz/
ztddyWksYi72uUejb3S/ebkrGCYw8pjb+iSa4YGq9C1RI8JJ+SFVVteEx30ddRV7
wM7m9tNP2y08V5Oi9UjoNYUrzZvikimZhilH0oF708Ari1HW5tPwzcqZ07fUd7Gz
GfW04M6Zz7d1u2GZWXGOus7VFmb2I8m/0rnYLCDIwNzsNsXSQ5sFca7StC15zXUh
ZzP35X7AQZohGwXNtpnaKiRAia6yXwbm0kweZH/68icq58QYkX6nUPNLygwMlqgE
sVpQJqszXLxZ7sElAC2wdEcWAobztkbaFd1BDiQBe61TcZkDRYltYfizKH1QZ4MY
RI08RyAxwTfTsx0W1mBT/FGQSUr+67YKkd2Kmjl6C8QhozM6KNuYDXcN0VDzcOwJ
CBvqQ+9aynQKzj+Dt4Z4dbfLDuLn0u/YxV0nodSxYIoYCpQsPZT9VBCjGKpkibCR
gKL07wFBColF2z1QSwsxkW/uW6eGPV0U3C7OD5JCxKvEkBK3mXlRT6RZg+4p8FLn
lLampHo90K1X3uW/LLmwtFB+UAyae20nCj5oai96QoXzxkgsQBeXnfPR+FUonNbi
ZA/tyv3wkppV7sE+fZdpuYQkW3sZ5ImDy8R/Js3FZzx+4fQldZQwqbE8cpY8PCX4
BktNs8Oxj7mtZ06KmQ/iqi5jwxEGTToit90/sNYxHyYtPnN7h5/JxM7/USZG/znB
tSWMNZwazokDQTlan3OPmOosLR5GlH8VxD4J+6Fdw23LMviHshyioZZCaXuimLWi
OrwBYq7t1jIFqT88R90czMdsVLdZKIB2eaplhuoUjd7TT7bogSBls3Vi4KZGHD8s
i7x3Oo7Lg3+9ainQUeXEETufMxZx6KExjRGLADqdfh1z6hXkt+rVrs1FYVml2OGu
T0cxjn+y/wO5IYnktzs40g==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
KCDZesYNGq+f8wTMBM6iKoNBrOGwHEkSJgtLyWmdrEiE5E7p8FrfklYHCkes4Qiq
tBxf/TBQZZj7HMuikV8cwQLK7/s4GOfikFX2nByXZXWODl+he8d5TtSWU4iI56l1
0e56Tbm1blS3Ix5SrGWyxmqqrRKOMIFyl8TTyWWa4F8GVTcBLpd5obW5Lh3uKYlI
FY3bK61Q+ZYJ1RoMMV89UclRQeFSFexkMOPh8D/GJQrcZN4KJQgbfr2BQ3PQ4XbV
D7sj+Wl2HeiGFGQa3adAZvFA+kZ8rORVgFpZrcoX7PlLkRigjaOuV7dxO7yqaACE
pijMmgoWyVDDBf4v9oeVLA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
HfoRmq9NeNDy3hikkq0mG4PBiKBobQ67cfAWg8O0YQxlHVWScdhPVbgbnhp7yxuM
zvpRMtny96/e4/zSNS3psXCG1tGIMswO8yfKRNjhYalUTGpGjz77vIVL0yu2Fjsp
8CykpcpHpGJIzr/PGMV+kjHWaD4lCEUeOJPgvbmm+/4QgnKCdwGv0pEZWh3pk080
EWELEsoHPbloTRA6EjemdiS2xqG1K1KnlSKBamvQGyP8XXgvXXNfNiQW3ssDPKOa
JUgc58QUDWigeJ9D6yAYc3bMoLdtUVrezuOY3WLqwZOmLN5jGUWDTULE7qRnLmH2
sNHz3r2DalB8qztbVn2VY/yL0vM7WDhm1/PMAsTy7qm0WdFdCiZmsGcKXnox1wv9
N/n2PXTDNqBTN3U74SWsFJaX8tPUIX9STtythGEYLP15Cz2Bp5fzXlPjq9RHCWVq
2pDacS6DjBLNOCxQZWMQyjCTHa+2UqaiC+ZKj3kOtvevpZEH3QpPV8osLipzh1uW
KceesGdaRcmE3LTDfYvKs/h1ydpS/DfiUuw8T1eit6ie0DhF2QnQLgaQf6UVEcRk
dEoX/Lu4U5Lj0TGZ9NGRom/6ghKgOxxv2yngHKKTPfUwdD+8GBjtQIHPOJJk4ELs
n1CRTMeOmRCocsphY1PD66j0yr/tlLdPYbF+WhsSq9Ws8FlxxC9WaatwZkZznSkK
iT0p4NEOrzi4spAGj+XjoLVbFPUYFIWC33HBHQczvicqqpgGyMHMwlMV1l+ce0mx
jSlshqRL/AXddk6oVO3RObiSYKmb0JtYJLnk2PI/ys+oJWfGqnrXUC5kPMa+moME
MR/ZR6JNp9hUV0SnOdQ6JqpO21lXwIk9wwRG3QEzWXRHkmRjoHgqKJywGchZkqw4
c9KaUNQUbSgBqCUO77MxbzBOqAxj/n1yxw1RaAUg+VpLT4zl+52zWY538fAIYFUZ
aeqFTVpBRlsMvYu9UiR8srWOByW6BluHCc9CQjQEYo1KnXDz6xUVCxC6PDYu9574
WqV9BjbKCksPwSEUIw3n1krgsosT1pPJoMILQgCWK+cnaKhm3xKJTOJJS5/WmE7H
ZZ41m5zDbPrLyQDkwOfWbi9UnmF8AJNmpp9+AFzjOpQ/5uMUDyYTjEOC+w6DfgQg
FM1xdgvDaL1O/zEYtpvU8G++GK04ajLYjrffizcqBxWyrc9C8rhdtKt7ljZuy5fu
i+s1WC9UoUJ5JoeH/18kdXFir3HkL2UB21pbFjW5ttbJUMsEAdqGPacFkm6EJprq
44rAOmPFeeAzfJubUJoMIsRbmIGH0DwHEhye297AAKUuc/Tmx9KjoRJjKA/HzQuw
NdLpbrsWdmT3825FeXEVdhJNQGfztmA0DXxRjmAB5m4x8eIwuQh1riH9u7TH3PQV
EBInwloFFkz/1SKSZUGM4ugBL8R0Q5Pd/+9ouw1W3zBgN1Lvgwj7uowJx9A+UEn0
elVKArKzct3hhf6o6XttZT9Pk6QqaQ7eJYzCTSBnmYK+tXXx1yLRPQXoGDXRfnKo
3wv64jp1XqKbsjP1+O7ufLOtVS3kEBebxJD1Y9A50D8jazHnn+GcVIXezeECOPVX
5wLYJvS+TEBpK9a40uXyIdrwIIZvkdPrEKh5EmIB35O0mdNWa9DTostAhPEGVNrC
2AqFq3rm70wrmbSBW6gXlORRmq3T123egcUkmqbX40sMBIDooABswCpcxEC4/0wi
yp5Cm6TCfeELnxUJ3y5ejemUhVaO2J9xuab9H8xyn5M7RglbOHLqNhSVpKdj6VtV
ZLVkDni84xre9JZ8wA/4yWpwv3LFV7e92+l3aVOxo4IEsGA6d/O8j24pdr+fzhwt
npMTtFk3zA6b9WtGThQFVWAN49hihhA4ObqzfKd67Kect16JZHLh74n/2iokUW8R
WPWPQIdBFopw+d7HlP3LMXpOQD4oLnRZKATmpak9d0KfPun6nJk3pueyNZDfpTQ5
+ANCcwT8ilUFkyaFv9gqVPEEKBS2zGyucbu5ynoMMTQABY50qBm8QvaNY7FzF6hi
/xJTFS7QxYK7tMiXgdmtDyQbZxBGiqO0JhFPUm+f9He0fkwNdNPJkuXriPLOBobo
0MxUUjqJwhp8ZcGoQm9O8uMjCKTmzIz0clEn9c1HeocjLoWEYoZNXHe+ZmJPmXOo
/hozEfX4hST9aBsOEt+9vSRW4UJaiLhKe93e7cw3fpAe7riC55k11rjDpUutdjiP
X+9EK+/BdsuHPWubgHxWQBxApj/lA2wJwIkdjGKxLcwaaIb0oKPZH5IsDHGICiPn
j6DX6LmvcQNdBOq0R2fHvpt4/85OxGgP5Cw67ZeOGF/0vgS+4DkfK98/qXFpmg3P
EDnciTshgnQE9mo33XvtH2FYRBRv9xQZQ2WbKcmxFzFfl+DZH4WRSqp1e1jy7qKN
mSQLRzVqrnq5z3Byzv0cFDwDtx6XDyatVJcElnNLREOPxRwvTA8jqcb6dUsfsl/j
PcEje5Io+r85zMnsxo9k11OakSHFmspaMiDnb4nxRN8m3Vt5lJtO8WvTNHmjEy9m
WmPVNOy8oPqPMBG6OILD106XMiebYI8J0Jl3iXVzMZqinPPfPxGHGVNazqmKvygs
tBTWxDaa0PKuOYSwhkZCe8epwIPYlHaRAyVjwNXZg0QrL05hOtA+SQp2lnpbTUms
IloDKRbvzDqjoIZqNgx+ql9L69aTPk2m1QRqKMVoVLwjiauldklSwPz1cNNQPPg6
7EjD8rU67zTKGrQ003oxh7OQWbpEpBcchqvymA2c1+UqbdDOABWTcLsW35tri/G7
h8wbUh2R9cw2qOVFxNjDSrEB/KQZeIfO3IR9BdtUUh43GdQfOSHru9eSnCJ8W/YT
701/NQybaSJvh+TY0jGPWUYStf7d5OvbMMFEjX3X3O8oERXS9F3jG8UqNCHeGZHe
GA79tbHqelB6/WNxz9VSl8S0L5Uf6MYtF6A2sLAX99KH+h0SDiFZjLy1d2yWqOKa
p85Y8MNMNl+kMlBhIKBoOhaWmSq8ktqiV1bAmJmF8NAILdrGz2XytoAEePFfj61H
VxXW+kuK5CA1f52I6/OQFqDU6wUPeXyg8jQ/5BltiprX/fk0cWEk8+f5T072btVQ
0unP9U6DoU+nljI7CybEQS/l4ym8EtFQKji9YpqE/jAjWQQ/N9yudRxIQakUdReA
jrKOJMuyWpK6v7mBjXEsKOu0mWyu/YFGLfui5TiPJM2SIrieqjHKwrnFVrsN2pPK
0E1lRGm8shssc5M/UeypCfCT17Ror8f1DiF2Z6ESUJ+jpaXCV4UvWfiIzw54OHAj
PkvXlk9FZyvwLxFFabgXOEc6UOP1mh0Gh/mjnJ8zPzj//bFLxF2t15tj/If0cqIQ
vJQJCBJpsmc88JF1kK6YkjN76e7tejSW3Zq+OgDcRb+4O1Uj9haMPtZhwOaFUYup
4i5k88o1GzRm1L4eFSOEvhs2nNLJxrmTb7FhLKB3e5ebJefky4rOjn9r29ndYnsq
ARBoxNBNPeEJmQeQHGyqj83nHqPnngicx+EqdeWsD5WPYKnBQ9ftqLWSoA62wrr0
RuPX1Obvy6TRsK7l4Cet7H0/7LABA+5tID0uSTZAjwrZRzlPKwovMnqQWgr7NT1Y
AV14NNmVqknjVeKkpzLSHYbztRm+N+vSAKTSgKibnLXCJyYgxP8yaK/JhKJdOJZr
Y8cqOhABs1AuBFJBZ03OV+0FkHE6+JQW907QgMIKlHHIdEPsNN9eCdvp4T1iELgZ
5tuIyvBeGlrH/w981EOMUg6dMaK75UMjnpXSdrrmL3icb84vESUAgGWSynhWw2/g
Yl8EbaZijKmkWFFPdiE76juCf4EejC//S9/91nZwPbqRGFi3yJWDEVIqJ9prVHST
XAZc9bnr8tjckh/k4A52Qs0BVxTlYiAxiCYF5GQjGCimjVIWV/afXRDrAbWrScgY
gp+S63qpJQ60ZoPyHo987FBIWtbg2JH+8L3eyZNSeojsUh4JnmoaZsBrt6aX6wij
MlKP/YyNUN84JfyzDIZYM9g4/auZ4WzKQZ+7wyvM+8m+2fE+C0nFr97+bSW+VO82
iCNQQQDz4Uyp2zEHLjB9d86eBTPFHwJgYggPt53ueBKeiHTsaLHNPERHw+NVm0TE
WFfUGyeJ8WLOxLc4mSOafeK0M7LnFY4vLECT1F7zyHS3Mq0J1HidX1+mW1I/VBnU
1EvMwtGCNWmo4BUIEUOvATde6c+TC6Hjrn0Wfyj+oqy5Gxq9AGJNlCIn0P1xlRL8
4hCmRN2RZCQLeT25z+b7GusPxKCHNDqwHZKasV54LOgyrB05EtkmhwHjQcvMhVSQ
mR2WrfXB76Tfa4kG+VlgJI8dvu2x5rzD6IeA/JB764XZnUoYIassGlk5sokXLN5+
lA/ifCnOgIA0vDCidjj9YbvN7KXkfoJF89qKId8HSOK61EBcYW32RT98nYQ3WVv3
ofdlP83Xb/PZmasJygL5plHMq3z83uidxFF9JGgkwzQ9Ah0Z7xevZ/lNsa+RnXe1
hZGzYQ3jOpm9jb45aeuNEMM2fKMvFqc/0p3a+ZH8bbQJlt2c+fXIphQ80055GVJd
iOzvME0H8nQrFsVPnmcJ8+76OvUKIjFprug+Q203DfsAn9xELRiRiB1tuIHGV6Ni
jQS+Gezcaz8anmitT+mIq0dbZ/D7tZhk6INJg5DyEwYdRjAHzJR6BhuPS1PfvqX8
J+EOo1cYLc6pTXhAfMVtfggM0YQAZ7JLLM2NNIiJh2pRjbCcW3T39Y+TVBTJ4jzr
zomRCz0Uy/suWaSL3esnP9AMIZMDVA74Bv6zSpMocN6o9aD5+xZa8Ynz5CKelmUW
JhYWnEK1G5VMXMEm7tFEcbHPcKPhedBYoNv43s6yzPvPaT873HQLdOiKP+mlIE7J
wDW8nqTokGMqJBloTS1G0VbRG12SB19Yta0eUjgSFdHfpuDCadXLSHiMKFZ8gher
Y/s6joFIsZlWOkBQ0Zc8YtIi3xd7GM6n6xs3MuYVO6aqpnKQV4OkJ8nRk/obccAr
4DjJ8BwZ8wlUF1i817fSZMBvtYP+OqJWvUmFfzlEWG4y5wLmOyMTVoIgAroAxLv8
A9jP31vz2niK2dM1F61gIm9A1Faa9hC+jQ/7sGcNpReKD21JCXnOTtGf4Z2kchep
yRnS5knmQammaJpF4eou9Hee5RD/XSv695CR8arKAKgo4xO1/uoIooUvcEvRJJhx
plgp7rhRuEpzOnL24lRoVMDejRmRDPrlDPdq77xMM3QRfF9HSxiQB/gZ4OyWgJti
zduQcqK/bkYBQMoMV5cKm36MkfyWBLUg2V6dxBoRmNhZuBuceveeHcn3NiYOGyfS
RwT9ocwfviSEJckn7VrLHVIOB1bGeiLf9VXhKjtdRyJPObRhQnhNZmbCk/O+NnHy
rSSIvm7utrqz3fgsTxyeXqbC+T5yB3hdRfzUWDGE/S2S8z/wjnMJ7CFjRHAbuwza
GwlFK1Tav/X8bc6Kl2SwXKZgQo4aweMim0OAh12jySaEqPd3Wr3HCeQ/8Bil+wAd
hA2QvdWNCHDyys19n+AtAGdNWmiYxXsviH35/0SaN1L0HEPsFdftiMddCHyBj0Cl
/xDGW/T6d8HH2fj1zgZug4ZmX5TG91lQx/ZTm0Xlq0AdMnAaMqqHQZFqYNsdaqyX
6KZGznYMBZO5SiJjiuxYlXdN6TWC1SuhKPJDneYsWay71VWuv0v3cF8sOw5OaxVs
prHRxGX1d8cNU7o52LsJx1wURvupZyeTh7jhNj6AP2v3ZyyLLC3M3uZvNa0CCxqu
ESgU9xyc3OF3hjDkS1bjn0+yg3W/clF+g01WjgapzqgCYB7hzs9zWF3GXHQBWMfJ
hWfb5h7kb0W3XkPjcgeBUNMYVJa8JY9XCzPTURUXRV0WG+gAsDFePoQ5k9ElHQJD
wRXmv1GHinY1x73/XANM26+JUU4eIHcIbFCGt/sy6CI0cBfPSxWpmSkRIMskiYbw
lClrQND/8mUn6DS1M8UIU6JeXrv7hLqG1JNIC0S0VOq3yx6rxkHESbB/NI75MjKp
0CTeEl6ODWmUgXpdsC9kg3/JE/dgpNCTu58t8++vMqAp5WWpcKmZhHfnsAGvU/zq
h3PRXJY8G8a6oSuKvrwFZOC+i5ROkOoInd+wNoLJ5fk3QkV/zH0/0bkaXofW3kqL
Bo9GZn42BBTG/HusG60vPlo5+jRJD+mclh4lsTA69uJMbalgN5k20q4YprDX2t90
gRRjj9YkBqbkab559ZYO+NeLFshQ0Cl+WWJ7FJItlQReCpU7HNd43m217Py8gaQG
AGDfo1pP1rbXyDAIvt1PcfFa+sC7NendVoy7ndVO6jEdynwTTnoBqKf1ZKj3fNwL
rE15BV5HJkq4h0BJySAvd7SDCvGAWK7yU85Ly2je1gU4QYAYl7HS4mUEfwLBbEVe
sWFmIaEaQ9VE33s4rywYu3SVjgT60AHt9hOZpTy+fXDbiKisaEPymzl6QASK+kms
UMaT+9jn9Qno6D5PZKepTrZdv+rANMVnQr8TIQ62jlTH6OH+6JWyP1s6d9b4Fy5N
/2fh8BasWqx2JucsA6vZIAxErnx5t9nDG1of7HJ+JRTsSPWHUy1FUDfND2gHUaz7
Eyp1idxXrAaj20hTKu72rNlK2v3JLHs/O3BXHaChEDf2DK0zG89bbuwfv3vI4rtU
RoE5rHFkQUDzC5GmTUZ45huYG/FmKVMicRBmVjSAva+aES7Hi5DRQGeFDmbWBuAs
j6lH2QVY5rp6jCvCHzvSFr3haOLj87LHrKHWXNIz3TUOm/lCO6zCS/lJExu0THR0
zBKFhi4i8u2lh4OZJVPBDaR5cYWz70NarHw0W6/H/anxsQx3qoi1v55wwG22vWUE
p9bhOOi0HAHLJwHS6En6xez+sR3tSlveA57x8VGsxJOk2fijPB1ageMS/CBQPXsB
IYym16wWubnLgtDP3TrlRJmS+/8OjaaKfkbFah5Pof83ZVgxmNMHwoVNnGxd+Eda
Ub99YWKkxYC1JGqxR5LMn+2fTv5wZqlTO8DIr2vaI0+vF711hDv3Ku8beioJ9SeT
wwwB3G1yjPAGCfVmt5agrTZDsEkNytgRtCGmPh8877gymnUyarbfE6KlOVNLpcvh
DvPDybW2ajU4dDG46JWmvrziFFOidqdUZx73mq9MjlGxBBjHKSM48LHSUM291GqF
kBFAHLtIAdxUat6+rjRzk25TfFdRsot7rEFlgLyXkw6eGqSUbT89mJGEN7OZRTkt
XuKAz/zrgsqyQMHSclth2Gk+u/k2ccfoB5b49ATTudTdwhvAxY2jHlERBb4mGr24
Gs4UaaqbMCu0BdEqZkHR9uf+mzLzlflyEnLwRMsjWUac2Fp7uqv2SOUlSF8mA7ti
fkaG0jcv0rbLK5jfF48Aq1R6WQIJmMMfEGOehxhQORLUGbOPFCDKYOxulDd7ikwh
cN1+biExD2aXBOnpDjb9W41vyfrP/GGqggCPObAP4bAk0gi46wQnkjzrrlKZlyKQ
QQByBxKtg6XabHcPxAQS3lRsOyQvf2WRwp9JvLzCOP0KHGUhqre9F/hI7YIdIgTf
GEuavpxRKgqECjGoDxKe7aY/Y6EB/T13aOEbJOUrKJhx5baAoImMm478+SsWvuip
LAWM2zskuQNu6WiHNRZQEK6WfW1RIFT/fvukCINnwXluUJdKJu8OHdaFQaBHr6DQ
E37so7StuuN/PPJu50RXB1PJ+L9VjbpMT4snVZFxf9Fj8S8ItqX3ANBCDS9BXIbM
3w9DwYa4B1pV0/3v9IGXc7Fc3NiNuDgffi60RYZ4n3oScZMM4SnKVNcHThN7DUod
9ebDLgY10cxZJjOT/I5KURScrnlIIQXuOq9w/FZGiDp50210bp4O4LnwEoeMDL3s
K5Xk49eBNwo60waCR75W4x/S5MYUBKAbMA2/dvP5cvr7/0mJdoySmuEciP39ml7Z
uVkCeeCCX74gRYFreQLh1Q==
`pragma protect end_protected

//pragma protect end
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
a6Kb4ul54eQfGQHok3PN+YrAD2U6p7rX7rbSrftAdxIRbrTX5hEt880mOiyYNuDX
SGdZitZVco0+8yuqwERROTW42cNjkjRi/bzhRLyS9j0PRkif5WqiRM2kBRvW+YZx
sV2FSRJOyGxlCbFb584lyGhNi4NhRM04qO7CDRAhQ131yuLSB3OXc3RYRvHgJy9y
ryDt5Aa6y4asKqQWVaX/0UZRjzeUKRZn6KD9D83s3DikA5MqZ5SXQ+yolx2d05r4
C+zqnqt1cfM8lZRHclpwj7awFKh2vrLldkBIZoKhtS5bwlg1HzZvI7RY00bVokYp
rex+lB+PcsTJ2cD8zHSoYA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14496 )
`pragma protect data_block
xD4ng+d1Os2UjJRpEmm+v5sFS54xFl+Rz74r3iDFergiAA22ar6iYY3oc7aXWSk6
04os32keEMNVxyKL1QVL34/N2xpKzQB1f7zKYxTwB6QcRlcvVwwdBV96iDz/cfc1
IEAUnLnHEemroNu0wDFb6N1qAIvo/XD92HS2UZxnhdEcqdgqFa6zeE4+sby9znnn
4wuYJlTjIWQnOozZIvqgb5hh9WrcgQMKcNFJ9QAcwhZQfyIIKxWohTvUq/HAHWMA
51zxXkgAWo5e8tRGflEmY+LSZmRoo1ThkUvjd8cLCzIZrwEa+YTCiH0ysd0wpGR3
gH5RWWZqiQ1jmtmuqDl06UOre3eod4TUspGk6mRgjBiVeJJWPKDulvUAtDT/Dzas
fJKIxCbwq8tiC+HomOZabMxVUs/Ii82e2tLAM9OD93EMKtq2Z6TQFR6iFSjazwVE
fqsvqr4QwcnnLqii2BeIH7uBpqowWPbSjKZVDaRIUCenNS3lQ1/cNZt5yncXRiIq
XbiHmXKXFsCTc4QHlGTIpnwrnNwOauyVnyCwT22Rzm1qeJ71Pxp0+XnquTBBsZTG
iBR8sxmeatD1gB88+hwR6zQN5gR3wXOyp91Sk1ohb6MWyIDomH9PPDH6M1XpGZne
ReaH4jIx9dREIZcNDD1F6tARgk+1SAh8I8dML6zt12Re/eEmLWXw9TCpRW4lRzRK
g554ETW0JEZq2Pb1IGgt5zxS+U3EmHl2x5fORT91tNFyXcye4JkCwonKtch3BAG8
pDROXCpr4Rr+yUnVJx5GDuQUjkA2mxGWZq/kRWC4DNr8Qa/LYyZgUXe7Aq8Vvjim
0edxzayHKoHfyzs9MYjvAFxKpF/S7Hk+DOI2UBYJKGIRwAi74nqzR4J49yQATBwt
7H60MtzAenbpRk0E9qE2T7sUnztd247ama1qJFh/LxryAP7jFSHRLOvPkQmsYm0a
bKj7eGcLm3xWO8VvNB5UHibKN/7ZO2LaZ35cDoZo6RGODtSXXgy9fnWsBX/jre+g
5dAWFfcqTA0lTRyk9MYxA22hDEurfCnsR8k4MHAjSMtz6yrxwYM8xCdzR/emRn7F
hPaYW2Z/s+jGguR8zxgzr7E0wb3heAn+WOaV7EoS6azL1sowNz2iRMbrWoSQ9lA/
+GHGNxJaDAWaOHQXlVcXY13lfB14fYd5TfExWR6EpLnDIq4Ed412n+MXs1OfrrB2
Z/tNJJTQfQDjzxeBagPHshgyO+jOb8ZWIocucpq9nZUH8F9+TOORvRO8OVBwTo8a
Wyqe95uOUmhiZqhLjJUu9Lm1SUIlwTFC6c+FJfpxVgYaYmmKbNrIdmnPxEo+WV3x
thradGD1gvkRFfZAagIWyTI+8hmjleo0WcJtptFHvMFs2PJPGbEKgtS6dKky8sTr
0kfICNBhPt5vS1DZBK8NUS+m9USrn5ULQVwsCGoi3n9cMIpZFIv/b6lsHcLHZC+F
XHh1C8vYIswhTYPoDtyL7p1/4Rcm4VGPBAO6Df3qeHjhnZB5IEraFpznddiCO/uz
x0dvuMYjL78K/nPudq3+Jo8fkt3uQA4lwahiCrzHVW0CTfaA0XskwRFnms2kl16Y
VM3NYWRTVnv4awz1cinYNzrsCgWD76xwYd9ILfjmUexOJtPEJC6YGSWv2DYssEZq
5eCVvpS+SDEmuLK7Aj2c4pknFgGCPt9Cv0UN+jgFKBokf2I91z9ikXHhPP5vRnKL
FOaT6ZDxgVSRNbefhvK3HnVGuf9aPxrMYzW/XoqDKft03C6d7DYDz+cZ9NpVXgg9
ddb9rEortnnUxwbp4jTaAmqv8CldOF8CG63QWqsB0NW5ag1sMqKVLGrv3HWlm27t
5LTjSPnlwvYoBPTMHJqELDV5M2lWy3BHsHzfbi0OM58K+j8CLu9upu33Whgt9n7G
mftUmj5vEc9GpNw07xJ4hW91Li7eSKc6XZ73/yteQOW8r5yQ+czybA9jikWlxanG
srd0l2wi/Jlr4B9wWlD+BI85lcKAayNR3iosB2o0vDh5x6GV0iFT/wZxn5WAnjr3
oBzhjj0oSBniOskgPOVpyijwtkUWsfn16Q7dlihuHWvtzaYVBSM1uOAGlScwkgGV
yQG2OydzUdauc0RosGkbu0ciN8JUudDCTznuqK3PB5pcgzqMMtOq38hXImqQ3i9F
J9KVqiDRb0Ld94j1MkOn07h3Y6qHwhKORmQyec6oGa41iR4415q57J+HG7o29UkF
krSNsrmjCutad1dHyLCNfXK8QkwznedyvvSNb04yuHEL+f6744zpwLN60f68NbBe
Vdoz81XLlzd5t5D1qxKbUED6h1gVkaGv4onMXziTT5mGur+vVJXZFw/4wAHaXh/a
Lr7lii2fDZRJspvqUHrDodY50CYNQD8D2ADRn+mK1sY2jmxVcO412ZswUCG9TTqW
laWGUfUaKY0wFl8rICR6WdXYCm+/tj3FiPOXRwEjvpZ90LQWN1ExUuClyLcAzPt8
0CWcKLgjsZhLWWw/TaOEzR/y7pLYm/KRY8L3a9ur2rWLi90I43myfWcxclxfJkOx
fTqsD8yNBV46jtPfC93AgccNqkHtcQoxeB2S/0sKm8W8Cgw+67XWO0tgA3+qidjE
k6qmFlBzgeIUCAtprS+8yGcSXuX2ZQNPZ3uR1eJuc8qUUhXM7hQ0h9KT/GeuG2bj
ysWUJBrByL9JUisP5gTgJ9IQNzgybZhpUgpnjASNDZpTbFPr7iwIJqRA9dAK3Ppb
JP3V6vvk05OixBjWJ03FKGq0Pj3sJyqYE01XBep3oHuEQ7QBjMVmN0/a8sV6cvQB
l3mb1AN3G9lFlse8XPeBbrXdDl86Du33SzODRDEQhNq4hufEiX8aU7+cqSEAwGIi
Ri2Ee7ugoqwGXL+1RObC6wGSXrbL2iLQiFZEy2rbAjyfInaQcShRr9fil4tKWwjt
P/CBEO46zBToV05sPzVEuaoTrpVZPpbtCPZcTb0AtVjAJ1R2fexMsUONREzupa2D
T4Ws2hXdvWria0F0HITqD+UAeo/wCCqgTbrL6Z7zRr7dzriuBi0q25KZpWFjXLhI
LShVhh3Dwe4vG80ZnFFqssc4afzRyf9PwTgRtBrM2vHGeDltqs4uJlVlq9z/QSOJ
oSW6Pp0pCAjZrGmZa1BASFvisXljdH4hDJMJBRxYKLyPrVqIG8WFzCVTc+SVWa6O
Q/iQm5xc2X767IlW4k6bW/DfsSoUu+F93tsyOHkBQCJp7H5SW9ZfeOLUMZpoYAyh
aJIr22gsGGoSXrVyHK1IboYh/XX6xY4Hl6aHZ50gcfGNYdbEUO0JRuOPFNMnZnQv
zVhU+X276cL6XU5jy2C2yQaonihze6jaHIxrOe5qVUCSERyALpbFXL37dnkcVCYv
mC0laNEFQ8gIGlf9qXWuH1Td2IKimwDWRpTSBV1Esbyf3KpimPIWCwF+Sc9qhLkG
h4FZww4M/rAKwAQu244uZaIeDoMK35ToKMeI/C03ni5qEtFtl3eoMQTO1BelNPDc
ni+yQ+6qo7gOg5Duyd/lgvbBIabEp8bc0tml9/80uqBTbPn0YeH9CbkmbFVZt/rj
uYpcNtbxEOWhyd495+X6NZL8K9zutrdtiWgKWJ46KxudrWU5SnRaBwpYbSNn8qP5
i7vHC4ODg26h4wgI9oi+dN9oofcSnwI5xFGH2l7Jsp1OXY0CFeE0agoV7X/XLnci
N/AjbtH+12UXChHzVDJ3XHy6SMDfXRqiSF/6+tKkG4n2zwlV+JuBzVr1R25ErUpN
z1FFBgUN/WQxjmriNooGHmfMcJijG8PMd2DXV5oztUE+JkaqcctLkUlZuuxzK8mV
LoL5/2sfvXOxRdL8pOud8a1NvwQnUeuIKFlr6qfkct0Nigzs4EcXcNYROLl1mUMD
3btpmJFB7h9LmfW+ttMXIVmrRfuq33c5vNeq8GlSr6SR/nBiaXizRiCHvzKXPhAg
Xw8l5DiGKGyJeWWvsYzEu4y3Fu+ctXbLP/6lQ/MDOVnMkddWtNdlmiYEPCS28PVw
DQc8C4dQdFgH4G252PEe9EQOWuaUHZ1Zm3a74xfEDFEx+eJVFfVUGirp9SIXwLzY
QnnVinWBktHh+ihz6j2VxB7XANsg4b6KKE0Exjkl48O1BI66eSNC8DOCP15Vw+3V
CdkZTY0kcOKDb6XrXIUXtQcBmCwcFovBCvFlpEO0AOefSS0Fux+o0y1R4RmtS5PT
hB7AtaTSumW+9aeBhrLf1YlUpBLXM1bxLkSdzX2FmA/UkCDrLQOQfDj6WbHtFI8t
WwFw7jttnuzxr/LoTcG2YE7sjra+EI6HiezkZIeUmQ961dJUx++exXWxfdivuZ0h
rzQRJUrYtUAOeYrdjqSswzE9/AYkAIGglGoZcGRE774/JzzVqFyD7hHOdbl+xdst
YXSp7rOHLjqWhZkYpW9jeLfgS9868ejIvdkM4wVplyBRXrryjBfJlNaQasNPThV6
i/PloJq2lswGCtgVyoCCHvV1Vq8QgmWU/6Q7pmaQjLoXzkNUtQU6CiGq1RchmNcK
/R7a5GiRYJ5muS50p8V/CUpC//lHM3CC0h5hJPsuOvQHoi7R0bbDYqcEgtQQK9B5
FffC2vmPXigW1cG/wAu7V+k07E/IP60sjwJ/LNmYm6JpEKc84OZzgsoVCbI9QDeT
wC008dPQzbrzDE6QhNOh1V3D1dpB0SXna5qcbehtU9Qmpj4vWmhgHgUSqBP0CVwv
3QjdIkh10uo7L1uX8uTkPgnqxxnKvMSPodCegOgiNV8O7YXKQ9JoLMkLE4zPZ/rU
yB59yazfV/dpwgAY8wsJhK/56iJ7B3Qk9P5nnPLo5MtqWzUbfuAY6mg/oUyQQeEW
riS1i7u11kJTu8VnWh73cOaKozJB/q2+OS6k+ZKrkPc19VPt0GVPYOXSdqrnIGnp
OlOa0LrQGhhX6sN1tMCeWQkFLqTs3XyP/YzRHjh6gPR+EuLAoD7GPEB/HnDiUO6I
ilYF4vZNiGOTEFlxqzlxdtCk1ZCBBHvRAupXaQS4UC/6CGu8UvpyKiY/78HQk3de
9+rm3KADlST8gjWXgi3Wv9k8gk8uRx1q3nIQjMOpfOOIPZbWyEh6rPykzp1N2tfe
seO8nVQeEN27PpNBo5zDUn9L1zkOItJftqoe4lB+5G9oBB0qXy3E9n8dCvLm3N8N
8AP2FD273oS4AkKW0aNFcafDaWEVcFfIOeLkfRZd8wGriRLpP2yjYGpSlx6G3Gfk
p9Zxa2CD33IvN/YfOididWP2sVFyDfAWX2NgqZGJ6VusYDkb6mfze+QpcKuR2zVg
bkWt4sfiBXZg4lCdylSaG/9avvi/fwwUdnP1sRfX+I3sK5uog3tWgBmrOqzmIrsJ
hB4zU/qcRLaLLpomFuw88ZEZHjhi+ZUhjTgOC3qa5yb7oYZNDbWB+kGhhg1vcR+D
pJtOWLU/sqKoppXcl7s2/zQbanW8hiK+lomIwBJTB4Dm7HxYxjpO1E++DcLoQ4Zi
UbqkdDdROXtWF/ZLJPknXhBLxS+ZVvD6WLTqib5+cVLQboajqW+hcthzHvLDrF/C
iU/Gy/UF3K3IybEzE84+/0eRKU1/mHq1ssPyOhOIJgTvBw0O1jOs4pwPPVSarjG0
i0377uX+Q34l7bvVyYiRSCweMOri8u2zpqkMUw1csUL+xCtzKGAG1df1gatYwKo+
oudBQCu235Vw7w/II8isqq5ViUM6D45BzRbr1Tj2K732Yr+laHTvzH4AZhBWAC/n
TkUTevm9BGIfbagvs3VltNQx1+A4DV3RTqjO+IzYn1HNBn91fR4zK5ZjoYtYyloz
s/BoqzzXR3KOnZ5cL1+vfh9UV7m41JDvwjs8jY9gdFdTiPzRwe4+0gJkg3WdCRoc
BEdwzHHBABeibSZhKne0+QS3GhjEyv8Z9/LdpoI6U9Fk6xJ/ceLY68nJKwp0eQ3O
h/iEcWax+tZkR0m9Pt8vtTLJkt0IPyQMf1zzDpzfLx4e9qOfu1EEyijkT7Uk6SWZ
nuqYs7xe4hCAQn5n0tyvvoL7T00JVOfS2UvmVUoDCdeczYTFWGPdfOlqNxuKory0
YyC829XJ3BeRNmlKG8/vqGFpE5AwlqMUrilgTQt1vcD98UStFa45ztU3zxwoGjxR
mQq58aISzZbg6whO7o/u4W7jWGMuVo5Fw/thMRnbMzHc6ByamI6BT1I6fXbDiPCm
DluYpk6UnB8D4pPp19mroFFlJL9WiQYBut8A8JZEcETtMcjJ1SRxMiJflfNltYXR
Cx9hjWRKhAaPMPhP4zDOcBw2ELQCXVhA7hBjko8GDnlv1W/MeMdD+XB/O6/v207u
pFfuGwE82mLRnl6cFHrI04hohMSh8vvj7bUNor9QM5TwRtwst+e8UP+D6N4Zj8uL
tVEmSb39XAab3S1SC7GJ7nMi7xPxKNv0NiCtZsUv4QKealr6/l4GfO6LbjUzEARX
XYdxdFl9sJ5YIYCT+FR1tUInMUDMhi5DVykvNjC+ELhFxef/iPpiLaDVL0hm1/jG
RQugRkNMekkR4c+wwSk86iARFN9+7rzxN5s9iJVg1e7wHVF0ErLGV/g7bazLa965
/nJs8XBOaIaMJIN/VV2zuS9dOSXGDCq65MoNAUe/W497wsoJ7ebU5zonNYNK35oG
wGlQ4ldNGVWx+KQRBMSJCZxsQk+Frw1FPXKQi/HsZ9+NM2Cdm1sVn9yS/uBBWwvH
qHWN3D/1WcmP/KjoQGNkfGw44qGy56rbEi99wtgam60QRjQDM0rL07wtD2Rkx3IU
moF7KK9V5x71tQeEsUJq91qf/5vvyOZCtHTpi/mRJSA5Phd5LEBiBfAF2VBKK5wN
axNe7yejFE+0T9Ss0lFe7/vQHFuYE7n4KGndAXpjEo9Q7r1FNQHG25bSFZf3Cyt7
ZHuUo1U6SMUgBVBADNd0H29gRvIKAhZbBmGw9ziS7PVVC+w+Y+cOxbDai1psXyUG
0wYflh6LSWc1PbHGeXFb8hlndYKt8poCSqmIyQIM5vtFT9ztxc0G3DOASxKJSpXw
z4Z4BIaTzD4H7laApQe1KfftLIGtvsiZLGFxph27E6tP4MzC6IsztkcY39p2LlAr
9xqaFGAMccWuhd/9yWtIMQonthYipzp905q9kDeth+F72z/slfPhoT/S5BD7wNiK
iPAcFfB5UXtze0Ygh+nWcNfeZgtG6PBmoriYkaUTWrsTC3aVCyLooGjhkBjSZbGf
VBZCzzeEqFdy9mcxA7iXsT0dFRYRDpurTcIsIkvJ+2+JAMMYibid4fnkycPigMKD
XRQmENjKvva0DNSmZ/1T5CZg8xKL+OA49S0I4mGSTx3VYWXbLG6lZMLolGZhgLjl
bmVBMDIQMf9mtUa8dLdwxoCTgzDSimp8JAOGjP1Qda5xoGq6Ux3cmx9IYD/Z8/B4
IkTNvobGuz5dUk/9gkLRWMZ5LSnbYxMrfpRIs8X64cZDH55LZrS6kS/NeUY5syds
IC0ZPE4RIxqF/2V1vu1pZBiUf1ZkhwLBV9afSt/lFlZsRIAUE9mG3tyG/m4D/xW7
DIHV8+xAZzbeC250iLmDbh29sJeAW5E10kue7X0/xItC2E66uQe7hx/BVhJVGXOw
p+sVestr8MEY3llZ4jPKISHXKsbY8gxTNdHSaMd2OFdwZJVuv2zVwzG3wS7ppaIv
gkfJKWF6UjheMFHZjDHHYuWuKsuRp3f3PHoP2pYfnfpmCx9IzMcK7xnmOqalsCNn
3hWtAfN6OsHcuNf4IZAzThAnfyTV/pr6zmJe9PVtFG69f1UJhDB3yuQZBnWbY4Z1
SywAZv2zePiWRK6B+y+hrFHeTpJ84Hs9aChf26QZwL+ZSJ34sucj4AIMK+Z/W4EC
XBj7tXIIjFkzt+Y2ENTFiIQzS1ho0I5YgJMffRuZj08++MXSD0HU1NaeS0rLjOc0
ZGOvl84C/h2jdRmt7wUpdmzBIjWXXEpjKBWEo8f9g9Md/PFu6FBYcfOZIqV/Xok7
08tiQiBsAzE71MO8ED1DMKjq/ttuh/uLKggTLgxTbU8Pwg9IU1Us5xsbUmT5E1tw
jkjzBFmkAtBDc1VPgkPsc6Q5J3xGr1w218j5JQ3ovaNOfqH/n1FDjRn0IemviIeK
1eklrYsZXn0eo9DRS/FYkFGJzIf78eb+RzoUuvsUG2YBnOMGdygQJZO5qZBlIRIT
pFYIQwQFUWIyzRlyCD3X1y1v+sUWpbjF5OCvf7HaZUbStRgeEFIMqrUDHgTVagDu
3LShN1zdRrFO4MdBdUYDL1c0rszHrKiPC4oyyg2RLgZ8ZV9uVlF9kFlqzBXtMEhR
j4bcE0Io65NPIW5V373dNeE8VhCcbv7tMZ+YUFYHnpjVP2PEMFR8Y9ai7uB36/S7
PYJpbKNNFY5uFsZIEzZCqepa8Y6uxNTaAbC02fZLxZY/38h3vw6mdtHwQltj5tNa
OG97jQBdmbygzKPKhlqUyCIeV5ho3P1ChXNXoFAg9elTcBbnIe/ADsqvc+CuwNfr
jsQPxYfOT23xk+0kccbiJ8awFHMpCj8htyhAgW4L/0IeDief/BHbuyzZ5VjV9ZTB
l0Su26LnIiMMoTP3onuAsHtboxXF8zp+69dmoO92tK7OvdLcrwVfUWi1TkA+3fFQ
IYhb562e77U7GQe6x64YjgDypsV8QCZQteoiOdIxLOFhVifccxRvRHQv/7AeCH1y
qXxk99RpQICoMCeo/RzLgt0JNCgannuDmtEumM5z0w0oOE+MNcsS/Y1kPGMJ28oZ
8swIA62h5+NUM/U6aib/IihjuymvQ2+rib203DpakoJLD0niHMEXqnLVlPNCjMj3
6bZoOj09nV4tkLQMH6RRiQZ00dRqjRasyVpJbNMaCCGJiXpWxTVkKw7u/K+oVB+O
2Kiczu4FybRl53ogMAp4BpmhQl7bb49Qd6Z5aQOKIjuaAoF8Trj84XMeWxgjHtgC
4sbPB+/jce5ZxJOMkZTEBXGeAYUQyh1ADs76ymb1qqbkPyT6CyrfedHaqHH7uWts
l0Vp6yVYY1gxqALwkywqVO5e3zN9lSDJ/Jheh3LTg3PKdxrAWWzhyA0JIcb6q3UX
ga1h8T72wqauNPbtDvUP5Fzg2YMTwrDBWEZ2y2F/HVeCrtYyJ7ftpNDOIPlmgzVn
hu7wg+CobS1mHMB19nERjSrLzpFvrqVRququEhwspQxemkgvdJW8bZXpGNwqDcx7
AIVLYSs3m9cuJ1oyceQ+wr4H7U9mvnu00CRp6aavJk+BSl/hmjLMZjv9mCmYY1Cs
qMaIFh8DWfDyzwxSE5KgUu08U7XiBHSc0ZpI+Xxbe29WlyTlrtLMRWdEriSSOUBs
etkz4ZiZZGX8UPZKO1BuLcjS6b2doFk+iv6LMKiUtKeElcog4+g/w3Z9EuXcXv65
KgkvRFo8A33V7jbK+IivUDskb6v2AigmE40YBAjD066dxF8NTflvJeLfOa6wZhXU
0kpQSi/4S0DpZlshHXbXT32xrph7JNwsSCjkaXOaN9T1078C5Y8DMfcKYHW92Zfs
WqC+1OrsHYZUO9gLTkJSAx2S6kgdNDf2UMsI5N05qNfvpUfewHqRjrTipOY+gBm1
1MiZq4EMRzS3JPBUMnyQBvumcHYVw8ftIXFor7gcdjZRiti5ywCmFqJsxDGvOa69
mfF7oRo7WIcZaHGLPDyL6lKhNWQ0YSdzLyK1vDqU3UWVenFjGuXZx8XR50IZV7N5
/MYLgO4r6BBInC9AMRhNbL/mW4H4aobNvnvp1ou6/z8H4GIZnR9txGVnhHsOTkwo
yx0vgDWq37j8pxiLv+OYpcvmvhGVibaGL1eTTfB3D2IavV6rA8rChABCd3Y+xsO6
s/woTh58QUYEFts6aXAMiSosBFUdjtzYCOECjHkj34zO7FpuLWLSVOrqo6WqIW3U
KVS2dsffW2I0IZKyNQb+czl+C/evxTmjEO+tYnvWvtDFvV/eKVYJUCbMPud/pDv4
JU3DTEIfDL4m/rtoCuLLHzpvSikEGE33tgg9nbe8DKYpkVXTLvY18k9ImL47gH5P
dYlxKnq9ekrqL0sKG6Opjvey2lFdp8aEkVlLHxMNeNTcWhItph5HOKILO42tZHgT
E2bXBWuNFWllX3XCv6lsBGt3eKE95PLKrUQXxPxIsRRKxbI8gKldkgqiQeR+H3XG
bu3z9niLnx417DWCnHQcLSyZ1ynTe0K4yJb7dsy7dV8DU7dwsRsSPrOz8dtUyrhr
/dqWiSDHSrwPibP+NZwCAiF3ukBWeezMxQ+n1NgizjezAe0Qzky2NMOznncsUCFW
3WCljwrlWL+yMGwIkN+bcZc8bFziVHmcX0KuzvmLoYDw6edBqKKR2adlCMqqtn0g
FuMI+Zh8XR4T4bh3Q+z/iAm9oiaeu+ig56WJeG8KsZIysjPwdszoj1FyJO6NiXHX
RZPv6dEdg8I145OWHiBWHhKVxfF9U/6k08izaW6l+fyuBiU1mkzmcPpqUdhIO5nI
ljzpQElzS40SGbEs+PTEGnpmZa9qxrcrOWCKr9w3n9pdwcadZ3xIhrL7fwFJJAEj
Ldbrxof5OlSBCUS0u1JEQ7BYu/Fiugb7/kuoi800dFLxTU6rzQggVOOfQYQyxdpd
uF+/MqZ7pkmSyQP/K0lzRJ+wEypVBTqbYWQh8p4Jgod0ZmuYic0d62VWm/IGd5KS
8tZRtC8baiZ1CwC/xcV1M2bbQadIontb0XsiKYszZ+jKpJ1oGFpaXsyGYe/HjJYM
U1nKmNKekFQsv0KPpX0Ftenm5pFllnGodIWkzuJJM86OIEVuxX0x8M3/tWcO0hyH
iv9qS6mgpLnn5b+vjqwwi8IQuuO8nBIcvzbkGcCnvWkcEiePDY+FlXrh8FhckuEy
iHGofQdxIZq9yPBTTb6bmbgOdWAcOXtj9SK+M/wkFtziddDkOk5sW6AWT5c+NbIp
yDJ0hyRF6vz3FQ/1kmII11uXVk06yjc6HKlPCK1JWFMG8+fcv6kHLr/FJydcsYiO
W0XT0b4w8jD8B6lLvBAZRCZ8CS413Sh/Iywm5j3fnMj9NnPJ8gyakw/q0R3nLmw6
FY1VrctS2QGL6wfkeqbFnQ1yPHmQaVmFE6qmEq/sC5liO+1IGo6L+473cZfSwnGv
eOSy/A3Sh4gyDec2xYkTdOK5w658/CVLU0Womko5O3D2TB1TR8BySXxktAmywBM5
WXDkbwwHqssRF9FDhXjPPIZ6CYgz8T+I6NkK1coLANZSZu2nhVgomkgcxdpukWe4
BiMWLQyK6Qdyg/kekgZnew07/Av6gIJX2tb7BpxuzfTnLHkwmkzZ916o3mW1sake
Ck8zDAoe/pA8gwm6FI3/9ENoBLnUjS7z1DCZgVewRjwWo0PmTzgb/FOtY+zbqOoo
I96dF5jiBP5xYO0sjHB6ybgGxc0rPevcwOPDJo2pt70cIiNZ6nZB+X4AKYSJAT25
d15+DgelFlAvSZAkcwdmZIvSHWAx37unwqK6j6ju+ahgTmEo7wQnZO7JLOOJvxTT
9ELwe/9RtxpqazjRf1/cHg7dISv9Iu0aCNWyESjzdpBJHZVpEXO5a4jNXUqCdqKr
PFU02TGT6/rFyqC0isnuELHeJrqpdPCiNB76W/kKxLY9nMGj21QXWasf0X2crgo0
hdvgthNdhk02YzZxMyLfsCAAXbKOEYmzna3jJo4HPWcwuo/wXumHnMLbnt500iIi
Fon5ztb9xjfSXM4Bgp2VPlIZ6XR3tMPwaR7s0zOmx4UCeDLXk47kasOJ2PHXXhX5
esCCfl+TqppvQrhqgp4dwf47PLWBnYKlC+/7XZBQzmCSdciUrsVi3ErYWnKXGhTh
0oR6c36ihP/qXwODuNe1EDZBsUJpILYDCDfknoQILgLFKuvJrvczwmQLK74G5R6h
uet77nDJzSC//fP575QCv4ZVoNEHl1ohoIgZQpmcYfZJgMCvYK53pABSRTWgR8Kb
2ukDaYlj2nxiaaWzCIxdqeWw8YMNjB7y5IiVvMOvmTnkuaFcP1QIGMRaI/XTMeY3
vKvlG772Wi5V3rNUCotdn2BnjHnSqXj3MMDErmbMrKY98YzvWL8LVKHR2NGfAtiL
X6tR0WtI/ePOtKoyBHsHRiW7WO31hU4GWsM5igSSeNoL17a+gItJjs78dPER1kBz
T+8gVzg67r+Aqxvu5OpsWiqmnG03hbLHXlX5MTZoSm7db31T494CkhlRKV5HW+WU
7BFfiM74NMaXPHoynPh5SHwTy0bOPCoI8XLV7dvtDSa0Uky8sbXxdTi97xSo9YVO
Q1vi1cPvHL+VssYFPryKwWKZIs49o8mUr0ldJN216Pf7ryYFsalIg/YbbXAgpXRf
dtUqtmO3k6UnpYQa7u0+3lP9Fb+naRqCwl9USmV7tvR0H841KobGDReypmeN19g6
Em5K+hh7JkNhm27/CQF0BfAVTO5pCumFvLER9HKvP4ujAXhrPuzI66b9uORGpRjv
tHBtIzz6gqKTyGoH/ChFcqQnfwAOjyAKyBCbPxPuw26MJQe0ZHOi3jrc1BfajuEl
HrycvIhByD6Zs6m8k5S4Clp+7B4kcRAVG0zsYx5MrL7MjldTbnIuLl1Yy1sXg8p4
Xz/mQOzztmQA75dbtZXWPFJhvwDxpcXc9BAXn9eRVVOuBBuU+M4vyoti5fxuANIa
+Od5lCEn7SWyA3pLlXZH2dki7OOrvoHFDS4XZptqsQDTdoawOzb54HR8lUBfixpz
9hNkplj2f3CEat5TP2tiZUZ3G8NyZfzorAtJB+o4KEJ0xEQ6suiETtVs42BA9so0
CueN+Yay/RdzwjetrXHHFjjNXBgQotAx62iPOhQTvNhjrzdqpTyPxkaKi91FLpdv
RQpZd2C/U/8/3EVGxwqdX+KfmqUgfpgflkEay78Xk7K0ngOAErl/77O+N3a+eRrQ
yqIRB/0hA5w3g/EZOM4qiFqQbawP6wMRCJYPffaYfgY/7jOz/EguW7BcF3YgElyc
ytd6gUSi/srx1IGTuQf1Uy+JPofIxuTHtZAp63fIH4r0i8D5SSwTY40adFacGvcO
6sP1tFK8oUpO6loFyQDg2WASa71sYmUUaGz44CUzZ6cS0lI/sCjX55I4YvO1c0WB
K3NVbnTP9dHDwhdNdoGPt+UQ/SoZWNPT1c4QEu8Hh4byCZ9uvC+kRNP6u74O59pg
A9GS9VqGIhIHI6nQjGYMyRfz0OhmxwW6QipSJFtULHI499RyvKAycx39VBfcQzKB
j6KHcYMYe7eU2/9HlGxLOH4cIoaGHuRBiIYmYz9scEM04c+KM2hEvAOLh1kRlMFl
V+FznJ0GGoJgBNGx3/fcmpGWgUEV83Y4S0AvjGquWOfx789nYacISs8049AT6NEP
xAibJUG+c5I3uCmvxG7MsnaA598iNBLK0XxVAVLXQuX9+pd5bZ9bvf/8JVPQ3Nxl
To1lS1sjpV7njsENXAvZv+HuFl57Y0sGwfRYHoeq3mw9/ZuTSeTFTVOdwifxmSBk
D2JMrwrX7DJyIxSGRxcPHAOAIRFz+1XEJqjsKErymQjz662+n57FlmdciZSs/0vg
d4XT0SjU9LeyoHQQ4UumeeisPaefFeEYmkjPeWcoEr9BKHQckBHRNEobaO+XuLhV
M+AOAQ2VEX/x7u+I0ZmxwfjjoI3W8Qf8rGLuhU8PnqyxdWTkJapV8/agDVezC6S6
hd9fOW1SYZvoPwIiIZNgE2muDrLBYT1ewNT7H24zaSJwFc94XeC5UMbH46+jWSvy
GX2bVNyToDd1qLxa3y+z2tU1S+PO6uZgM/r7TBuLbGCHVSjA2ZPAcPlk5Z374csO
ze/6ohu7j2kNwQq8YwYOW1jxB15ZS1FeBpCDiqm4+Js2naMjxWAszztat8oZdF8Y
pCV+mrcU3R/hPIAdvb9llqE4270GVcCfUyRCkx6vC1ajJXaJCOW2uYgA34r6OFqA
5/BKNCaC8YZF/wZNykFGFXEpaRM6Bf+ITDNx2RqLU/HGt/CUu2HFOaI3oXp9ATeC
ReT2ip55cI0WoWW3qWtSGszF7O2KdpnYvtM9lxHsX+Vqk+UDLXXbiUnLwIhP26UT
A40YiH2NLT3TsZFjokw5Rx+u2trVHGU73eToS9IJQwOuit8QSg7Pvp9rJnEe5Tu7
Z0nIJ634pWBO7HWLU705MzGwSRXFuQKwrCaTJUZZZ3JmbPk26R4NNMq9oUixSBUO
MGb5K2s0fSuGvuWALgqqPYnkhjeQO6vtQPyfm6A1KhOffQFUS73Nk9yAboWsxFCg
kr6tz+n3pxYbiIXg+Zov2A3v2CZKy64YHIwLENfwUhjCqINoSxHaF9yNkBx7w6Ml
lWG9jCqxv5qXFASqXMmwCOzhManfYH9irt9koJqaoo2bvx7ewHKdk3BggyitHkdz
5NGDon7nXe4gP5UDwwua379eORZ1laFQu4dIM4ZpAFZjNpNjXBHrtkxhkw+hwGKm
nxJ2j8gA1E4/h4zOScOZMYNYo8CmnkBN/Ra01c/7ejcgWgzGdXftNnUPpeyt001F
WPUcFYkmnUOtVXB+Qun0AXViT7N3XvnvOsbZIQkg0eEiJqVSGxlC3sz6QoL+ppK+
iY50kfJDsGcPcpteKM4zubYqMTR3jh3Fl4Z1wdvJcRN4jUov1DZ0yE1fYiNYylfI
l1OHiVpf4XYN7Hahli07sCxpki/uwTJOPJaNgezn/P2oMuF+9V5egnQf0kGoKVNc
jIWNg4zqikrv9lZ5bB1jEHWIfnIiiHVMiReWLZVe0O/x5dU8gkBaS9k01czghM2j
+SOEcTnkY69KichuWdd2O+wv1+kI2XmGl7hm4kMDP+Mr8v8o7frG+v7YKFHipnNH
LIANgamMWsQfUhFQqS0VAxhhAi6fE16r6u4hRayILKK2MuMmkhVn7YlAt8xAATj6
N3Dae4x2gOcDLAE83rPjJaPjh+19FBoQo7bJq3W5kjDLzpJWO3gImbC5E0prgVqt
B2uGvXZkH39J8i82L1nGwrjzmhMfgkn0NCG3/4WHza1neBt1KGtAAT3L2qcPApTs
9x8BpCUaaH2QNNzDZ52iRfqM3K/3o1v/eG61WoCblbuxlzJUdQ1xhjeX22QxgRP4
chIqqOrT8MKPuC3AcAwa3g6IDlAFb7XGp2tV+3kBSuOf8F6snpCB4RVPzX9WTorZ
QDhqnolHoNnepM7QdFLNphIM0kWEgqZbI+4h1hZCFZSsyIorKNC9G39lPrPp7mJq
LhOUSBQTK0dxNy6kpfkYkBq/pPwLW5aScbxLQ34EbqHX0TYV7OoG+bqcquOeTaNQ
Hv9mVEb5o5fPvdZ2vFiD6+mMHt7QYMrBN0nAhelETYd/CimRunhDKKxhzLgkdRsc
Vi1Tjt6bQwA/MxakpggUhUJCaXDTRmafRVCT0o8cwjfbRvahPPjrdhmhAkdf3n6M
tLpGCfke/3DCMFKh/TmNE26hvp9ORLe3crPh6Y0ziOApurPv345UXdScaPI5Ew/h
aKipkWEFuAKgMn4HNUXDFv7+OH1rXoX338bfsCTrhXsWJVpu5ukVOcJbS1YFExFT
JzOzjqWQU9yB5ueqe0dTZuWW8tQVt6d1LBqxhfzb6GZUaMDkV35UwI0RmxZNvAHz
gmqyTjwZlmI4utXYU9Zfs62odGHwhBMQkzIhuDlbmIBx+QbH20kAAdTMKrXvHGBj
th/l/2aqqgPu+tKw4GKavh+FIlT/JgAsPvoEh7Ks7cAXSa2fdLgQ6g/4H4FDZylP
tOLO8ToLBiLRvoS8u1GkoiAZt7xlPparQo9txFMrrcAsxg5b3ydWkM/CjP8HPNGF
munSG+HG5Cy3d6JnOUR8Et9Lo7uB25zQK0bBQ0wj0d/d9S8Tt8T3tI5dnfTTpxWq
Ef8pblQCAuf4jHZy9UXgA+Wrjvqau+58iDLCMJbCXEQu5gJ13JB5n81zMi2Ss4d/
f91vKLbtNvCpjF6jYc2FRlPt4sfgUnQfe/3hXt7SndQwdxhE9l4nLBSy2el3D0MY
k5DNkKbeN2Y7qi9FEqqV7fumFO3pFZda6pioGdpIpa25terxH/maFqz9nmmY/z4j
CwCIJ5p2wMLb/ba4toOdCy9jejxxLnGxqmY55Rd0myjHRy2l6PuL/fdeWzI02wIB
L6vWg6VCLGJALHzDxybIrmeDQQZahmpruC4DnKdIm5hCV00s1WypSMlQZfUBw+9L
VSunyQO+5od8OSQnMOOmggqZsNzCGmUXL9rGoPIsGmWn/Vq4DEtmNejkcL7qJNiJ
JurPyZrxA30nFpyUrAlDaevFW1zZgVebo/zCJj4nBg7DQrx8Uo7W7BoqTa7D+h8X
bfEY2/3qimT2paTR63VCwszyHHzb5adeRlJIifBsBTy9NUvUC/Rg1N7BKoTyUI/f
tGAjSlmv2EiS6yX20VLE2GH7/pfF4Q3Cw7fXpiS8aD0OpbBHRQbG4AlhXD9x8Gav
H+HcU2g+hJFjt7683nLaqJDSd3acFiJrRRmxTrkV9GpVTP0xtNZx9sM47O3rI1QI
AE6eHYnri3CtYQLF3N3iJoP8/gqjj3J8/2Z14LRq4MXLEHVssO7XvHuHoE6GHK4u
T+KJd2pYuJnEyqeA6GIxxq8VHvFog4Bl6SkxISmnzLEfhgRbKMzcXQuJE8JaJ9/Y
+7/6i1BAC+i8/2nBzTQ81T5qefDJmVl79EEMX+wJK8b//mUHyefaFz9s/a0aHQR1
CDCVSqnp7tZEOSc60f0H4oUbpj/y+ZwDSnF7HAyIzdGJG6StaahXqxtyGVgU60ZA
/dE7+ElsJRG7VQHV6pPlvHttHyya1SPRYziOKP7K5B6X9JZOgakIaEqAFbiNx2vJ
nNdP5R9VxljkZbZl3Ui6MnN8r/K+rDGOau17pvwlDWMsA5clRtSqyBN5yHcFi6B0
6CniZPv2uzW4G3tW/RukiVTuMiaDaphbbMaFEsGH9fRG2IRRoulH4bMmDoQwFVt3
rYKp2GQDoqTXZAriEC0dDiOOGvxh/xOGNkpRGXIf8wYUebp6YR49Ty8pYImGBQck
92Mg5oTyicttQJLcnb/QEemzuf4TSYBUVxF7Bm5btirSMT73HzStdn/5vuE1B9Fg
b9N47V5Eij6ftuEcSbdRaeFBij2Mw3RyT3GVQrGfffJs9EnNQck3IcyUDRwVMYv4
cOCDNXwyP+0RZjUvnCtHt49UWvZBbEtbZcRMukogUQX0KIKANqdupz6orkfO6k/v
zKymevEuFWsyTBuZ7BCEuAJ3X3Te0obuDNgMCwjJIDbfMVydMiZWa7DSBPKDHp/J
rVydjqx8h62n1sDpxQ1ocH6PjFMK5pFGTzATLy0OGVBKqXwV5gPXumdb8NijHioz
zwgKj1XSR4sC2zyxsd5Fn1bTnnlkijZxIrz02E0gRGSGVJxJ0eAl4QF5GPIBI73y
JHXhBVTI51fDyUb0IOs9vGfn3Kbm7WKNJiwqAR4eCkqQC0UkAWDaA19SkTUnk08u
Tnyrbtbq3EKDrsiwooTKK1El2hO1dQXvdHEMLISAW/vIqyvFzHOUaofvhP/fcXsv
WPP+CnS5nV+EHB2PYC8qqluO1fprEHZo1uDAp7DsN07hxFca6jBVRqDuamDCgaHv
xQQeEoDOK3ghs1GyseTZM9HKj9d/IMNY+V622xaktUDPuO3zbqznWQAEhpXYYJ1q
wSGJpe/uqOm2+ofdyCHqOcSzoEVLC+u3Yl6gwjH2REXBmj/w+WLuMM0tR6a3O1LW
CWi/HIL72AyOXwOEbeMB40qiB/qNOgbIvV+4nXL1J6GiQF9AjqqG0fjrPq3aYYu/
nO6mMWnhmTVo8Jf883osy8cXQitQdGdrdEqTSId4u+JTyBqOXVF9MksSTijSCFGz
s51vyAcSH+1GQlCW2oL9VvLBAIDFp8eVk4InU4iW6tM11XKS/1k8ZhJxs/g3FF2o
pWBh0jL2Du8L3fwZSax12k/eOb30WUD4ofDcxNUdg7BY7HchegPcmXT2ISFYdwWM
eQA5XlUmRipMi6hitt6VQpEHutPfn8xMpFOJr0KAApwzN8Wm8Hye0FyfV8LcGtTZ
PA+NZfpQknceiJGAKuXpQDV9/efK615si0raC/QD0fCsy0p6iyFqA6s0Zw7sL3/M
gEKFl9CMPgpAlB+HF3nB8EeZq3i3mhn8tK/rcaq6otf/uX4Sb7bRO2pX5uNSobjC
ktUtVuq5ovPkaU73KgyhNRzkqweYdq13LYY7yyDxTWdURi9zWVK9YM0V2RU/OXM1
WayYlwHDb6aobTeuKwwrHCn9nq4zlfmcwLjcE65x2CCVAB+2vFSYNI5dAQrCG8lO
jfxuAuhe3AtJRskuFOhjVZrz0Gm5E7riSjNunwjCRv3CGON2mYGwg6POGf8d7GL3
H7L5h+J2JnBjJ/tym77fPcGT2suwvJUY1B0tRzr+/Hboq6N5UN+K8ML7IJkxFyXt
lfoBfdGCOqBH+9b/YIZMxJmaHh3z8zi5lQeDX1N7ZjGQvIqhYkI/nXuE2jlM+9ZM
LUuEJs3psBS2koDxgLIaF/uSyCJmaPlRFEa5HWbX5Zq4uSXjZ1ZWCv15hB6rvG91
C7NX7lDi/VBfwP9983dWWo17rqhYUg0c/lzCEur5CkxyrDRHwzo6yT5nUEWpAcf8
C8BV0JzOtlSnNdk3UA1fwcoLuYzULaf6AwYqUi7l9st8g9kMLRGeS5bDJ6OwK1KN
+oF0Mbv5tkzVbsFqvyRKI93XOoGbX8bHPIxKgx/+BWq6FYaIMar09+1jJWrlnShb
47ZUKoojcYmZ2Xdve6GnFWjPGaT2qervNIxNFnPJ6UC0gt250rd2OAcHKO8E+7gT
noMViekQIWW4CUjfLeoJTYGmqjYcbcaxPude5GfllKKQs64OMGpMB599cgtyuPZp
gzn+Y9JMvvjs5qXyvn/aIKcYOOsSheEVKE83EK1wBMMZAXtaPiYAxFl9bpkTVJbS
vPoSxPwzifOLD6CLsBgGmVQweQ1YDzsDSy1kcYtbmutXMAHH6jbsUKGzJsh+fpQz
ke9VTaf+rhg5MiZ6+HtUktjMXo2TG4YCkqdwAUlylxnkwO6h6WgIutaty9OQc6hj
9aLWThw1V6FKUFLEdeE30xaqwV63BTXw4+VvNAydS8pCtReX0jCx6OTTIO67QiAP
cqsom+JFR7MiTXpT8Mp0a51CrcLumHUyndujOwABSS5oE5pQQ10Db6zGDh2efeNF
6ZMzgW8hixvAjyjmi/GrpBDB+PtHKOs1UdvVjcVFiWpJP9Kk4cdqLN3IRejWIghw
IWlbvNivjcjF3o3zkL8lWwWWILkZtl22EeaGNN+odhbyCAZng+Yn8RHsDTan45OY
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
CdHQtyLgQAkb6YTOE5TjC3Vj042n+sq2aBkdlaFkpD1hVi5TfXsKYi+lmqui9jzO
GquTzAbiniY+Aq+UujFPPNHNl/HAkbD5RusOQVSZXWvW3ZJMxhRcAMPgGWpMgaMi
ivFhvM/QlUIaxZbRzE+Hyk33Xx6sAW4cQimninliqgmlEROAGxzZxm19yKhwUsOL
hhpkNvyUwP5USPfyUMoegkmXhc/ltz9pdT7xZoZ3Px22v/sVOcgdCxYKpCWNCE+i
BCluexUryvNXXLBHdnWnDS6tAngF8irr76DdcYup3aiXgP4OYXXbbe+EFF3F5i21
gmOLyd0ANCB62T2IwtA2Yw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8688 )
`pragma protect data_block
y30kKVp7TIZVXGzBR0hU/PaMAVFor8gK5tbHWZcvXdV6RFQ+KfON4uNpBDX+7YAz
LyRNDIPAhTuSSJbAMQ9fQLuY80Xr0WWdF9uqDCSl/tK+MLwujo9wnFzpf5phoRM9
U5rWkgQKC4PGovqDkEGOzY2kaRxNlYAboyGkgPNlwWRcA6R0z9eypo3Uivwof7SX
9jaaoLgX4fudpvOgcx5tPSPyyoGFAgqn1oEuTs1cJsSqKZKSgUe0WGr5XcOc2Yhl
PiYZh5F7SNtCPnl7nL89emNpWoVcGlyPFU1jZ/QzfhLksXfBkDlh5pIuxMg2yp/D
Setiyj/AeSeQkTLvuZH+K93fRFmqP7853Bg1rchrnkrI01UlmxAq7tqWrsTCeLmQ
RjtH8OpCrV0ujKOzRxlJrpM6CnJ7Hg2Pqc1HxbnuQPKz3TcJv+aMzJiVuMfVLoo5
t41hOsUJvZNYcuPVouVFg1KS0rnvCwtgoB6muMjFIfYQva1W8DFUvex0Ik1JhV/k
X483jegU0CDCnE/Pit/vFO7lVv6dG5MvlwKLx6l8zt9EAJTURQW7j2hSA9YLTNQK
CfEjtoi2/qkHWFjkNL/5abtlXhrBlgGQUSVTE7cHJlepmOlNRTrF8RvZTrtdnbC/
1diUTyeLARbmZhPlTCSWe6j5Ki5ccOhHNfNn9vivqybHRJ4LxYDhQFXrPz6/PNTH
ZoAdXc4fmnDo68MUCbAcpxeJh05J8mP6H8Xf7Dq1CDvCaC4N10bR7n7NGKXGE9CC
/fuD2LUB6G7R/3S8q7L8CbjOJbSctcGfsxxhOzQg0NI3S7bX0nawAGOf3cxpQE45
1EEVWJcUYNPqSkPLMC7AW2MCi0OsLUf6u8FB00hqd2u5cgIRuksZjPiVMGe9b9Nn
0Kb/wKZzUwRFI0LnRzfweroVI5YmLuwSCre6w9JEQKVNSCT7jb3kLs7YHNzAuZB/
9Gok8FILTtKmRqt8yWM6l5zoFSEUoyPFc+q62mOXDrlr9Amx2lOlni6SModCTYop
62g9AFlbkCXxybEJq+977sHob+WxwDFOPFL3Xb7qj6BQN7hzLRh38WMeYS4M6OnV
XBqiNL0byE0IrX32OEZbm7Fyk3TDGczLMBfSVUlYXpCG+QWFBSDdL2160D7cZPrm
kLKx/xonQdABYBmr6vqZf2paPdjVmZ5ETqDuJNh1i4+HS1e8pm7e/etOS7RH8JgL
1EyA+LdzrNy1Ki0ThjpZ3l7eaeJl7Vz666gPo0v7RRhXo8wDWZNJn5X5u15GwAHS
mQKAv9OoJmamJ6A1a5O+x5glxBcqsTqKLpTPLRUx9452MgmlPui28QzvYNhUWY2K
GUNs97NrnMcQylhBiGbhOZT08L9Prhx6vESFpFdaah6H8VxI/3t1dclPnRh9ZCQj
P8IGf+Io76EAF4sueJmWafhHwhirPeJtnU7bglH9LrYyqtH2p2u0ORqvpQEuRWcg
8TKJf0dAR6QDmF1Mu/2t1BTtN3T/kk1tu8kdsF+DB3EvfSoZtXDbFWavxOSPyIbz
Ba4VIeQsCacRVNbzVN1Vc4rPSMEIYmp/ocUQffa5Y8Mehl681iw1tVVpMYgide43
wLw3AnsbWXKbXTQYfbvbVt6AcRDDQJ8MLcJtJbD3ECzocFEXl0VCEv2HPqaxs0H7
+YQiN1czRC8BFFebZSnkVTJ7Rm/4ErHQ7gMp2BiqY4rGtsqEVqlN5PV36MXvl3ws
UJDRpnGm+L05/7OjGvUeDh9YrTRarul5VmSBx5cin1VvxNa1IiVQPWeg7iG80q3o
KZq7Kf2QIbDjf/U/gJZqTZi50Wno4d0ivm9KHFU5AZLC+pmpOT37rIOmpYFtYPKJ
y5jDrDvHREZDg3NkV4Q41Uru4or45OVRvDLA0q4TKJQ2gjPokoX7jEho6BPa2fsi
CsT1c/Q34MVDOGnBAXW0biQLZQ2X5MTw+qFnHZ68oscfg8f9uStwKJUn9UXpGwNl
+wCExhGjVtjv2SJ9iiRDu0CspREPU85l48H4s6PSOL73FXJfuXTr52BunxaE7Ktr
3QGQc2as7oKHiU9Yi1ECM2UJESd05NDJ8zrRqndJdrBbxBTspJ3PQhbrOIOigYjS
eegnDjS7NHjrF7RCYMkfmWIJyD1QmObPkicyQ3gDC70jLvUG7AN0GT7kA+m+4cWW
tpamUKdrkQY2e/aW14OBZ5j5jhff7ciFmYJaG8nohDEZQDYgiNWKdkV3obJkLGSH
6S4PgAxPbl8wZ2LnBOJ64oePo/sScnohKqfHNT/DV9BtUgotSF5AYfKnV2/bZgZo
Q82Rgy8+t6UIvf4FotVtimHIaCfBtP3AeYMfAkRTjS45e3T3G21x1KesQlR/p2kv
gPrih8+p+fWhOMgKp/5yx7pDs0zb2NXe2CAj7btIvPEZLn0+E8ovsNIO+1DiNwpT
ogMYcxLFbC/SrxWt7W4hr6dA7gCFx2kroaokRVAHOQwU3F6FfbouxzDzt34+0XZb
nyysCqVuSyeSb2ASjdkb96Pjq56tiR/3ULEiQS+jvqGjqfwyR5wJjUweXup8XuU7
IRm6cmRkzOyNtFtPWiF/o6gqa1NVEai47uBDarpxsd6NkrD+BDjy2hpimSkpuvwU
t+ODT5W05uN4glRU+YgttA4Ud5nl69uhl9C0RBt9NLT4cP94e5eXs48qwW8u3r5I
8+Ola5iIYaCrmtKFO2MLS6DRL7z8PMAfOMmq+We5EkuKjT77dj9REvuhek9wJ5U9
sGnQBLjahL8D+Jbgytfz9dzQ3eEpKymls9ewzQk0FhbR6+Axf3a2RaNkXkByJkih
oNuGtFHJKZ6XY71w2eYzUSm3z9NzUhglbU7qrPmOxiGylGMB0pgMyeqNevp5EFsc
47Y13vtFUIdRH86cRly4dd7njg5KYFrt3SBbR5ncmUbnwJTi7dwSwmzpliCewNQ/
aDVGP4YEj3fN4w2aTg4VabtP1HU0Jpiqh54DiNCYw94w+JFf0/XHYKdBFIyjhoZK
UoESezxQuXyy96b8Wo+dAc+nTeeROnIMnMxffJFutAB799lP0KfrahFVqme6vhQ7
yFPj/C0BpXx0od9Y9HF19THig44A1yl4/A3Exezqk5UgFPTkasSlsmBFaB5sOM50
8DEylk+Zc3QkVicOnJ+jNq2NY/rP6i7/fJp9cygE85aJMIKof24LOgWsM25tKttq
hG3ddaGMZeYfN/Jz4Z0YMUMwizWP+Sjz6gA+v2DNAjiW2HJHzxoav85PQJSoQDHl
eTRgbj8hlWsGjHTxckWIaT8wE686JEwLw/tVTUBJ97GCa0lQtS29MbCGko2mdav3
5P/F2pILXiQcM/wvFfAgG7iBSkD3zDZrNA3yu9xlZJwQA1GFPOMi7mz28p1X1jt7
kuzWW+j8Xkt8WhHDOXb7s0Q4C/XsO/RimSmJKGFxFKP06S73ypRSV6E01t5ZGvok
ZxUY86MHNFBWC38MlDARKUSWLefGGOEqmhNmT6i//un692MyrKjxHMLisyVWVHcP
nmfJuAqOuSQCKiQFIywpz0Gw7Fq6jxJZq0E+NdsQ4QAvE1yBTVO3B/hA6WXpybiB
AFnTK/LNVTMifARgztx74jDaQGwN7iFH2EalBPVsmAs5Z4vUzSNCngHXXqNVUZ2Y
C3b6QNEUrQHHInTpJGSEa9DUq5nSreh397jbnE52QtpUXQSeGHCX4gmuIYth5lZZ
Fjm12d1t0G1w8C4A7y37pWzH27RoY/nTCK630mLMWtx1Iq2wbAzHxnX9okTixYaE
8Rbg7yXg/QHCIDOrqtq1PJ3AXtn76wI43+oLX9TZBxRwian+7EBeGh3iwjiLqfep
1gGX79//8pqWXZYuCsUTPaySHzEUs7us7Dz/HDkumDtzgTm+JHZhtTs73v3urwHq
4XZQRcwlY2wTDJbQn48gJCQA1hTMwLJEixXWn7Mh3BxQblYnSVR9OkDXOCuItlY7
8lMgK2NswkJYGHxX3CjaZBizBZqO4cI4KSGhN52V/cWKviE7Q+7XVrojucErFokn
aRRmxvb6GM1OU0r/Aflw876CBaC+JVr2EQE9m3mrRitt8PhiuBJgwp2Cj5qGKBcP
SF0bAd0REFJw/t95+D3fZh2gW/QXLDgz10lLgOLtu904r0K8OYkwr2o51DsTQ48R
oCUFVtid7DOwvbPio6m0GAn4l/s0N9AhtAWQDKGDOpILuxHlDlrIAThFXCavp0b1
KByDIb4AI/yCTls5pyv9fFEH/xtuDZaoJ7l5FVgYMxGaM6FkxBnPuSvkAfRxhHua
dpRErf9cD6aI7I0ElLwL1CXh0ub2l8VDYsPGFxUSLW9wm1NeBMSgtW9oklyVLuqb
qB1jFSe1cQCb9MQZZyYHm35RdSO4F4LDOiGX7BZPVobMi2SgHLyIxoHG5piD1y8Y
iGl5CuBJJzUl95aA4T9QazmwW8lAOAFhSMwklqfqfwkB5qauzFcJE0Vw6ZzkD78y
1P1fGcr8oPZZOcV5MIdFRjk+3zhNXWngT2bNuPJjzCTlKX5LEg6r8MB59a3FUaHI
YzW2bm8IsMTSdMC1CytsLIBbNnFDtPi1SfHEwgXWgECVDLnGyEGjXLD0zhoQv+G/
Dlg7oV6kt4p9DArgUBC103IA7PhG98zaWx9ksjlXVJbZfi0KLave7qVfHRzM5+xe
KKvzZtW5rZPPRt0F+mMg+w9rOGdfb4eoQVvLAHSpSUofgr9+nJPixIuLP9IpVEBA
u/hjC7JUaE5MR43V6hGaCObWsQzfkKyZKPAxHP8sI079aJbMyXXpuEOtgtj6F1Kb
NBpXCrOr3mTCCPJOcrY7cLGKFzrMaZh1++Bnw1wCggR+/1Rzz2X9eXqj/LD6J0GO
MFI189c+PxjrnUYujWfq0JNtVVLGMGs3xxO3w+fmy22v8gGl59SyXXAQ+1TV+iqc
47lPzfdg+Ru2jngqLJByBX7BhL9LLDk0ae4eFWXgi+80Fhpzcc90Qfs4Q4JzcAe3
cto9LVRAPcYws4m1ZCcMERNUucTOWgLXrFbMa86bwvZZctRbK83ecsyNI1P3IsRi
Yvl66U5UIc46RyYNCPAIPu7vbtBR3+UqESAox/6GCYba1euNEHedI/U406hYF+no
C7Xj3b3LF04d3lMvpzpeEOaxahW/eTsbsAQqOYDtX3+ypNsvD1f/u0dI/F1xLNMw
dXbnDHF/DtpvFPT6kbooFpS51GAyWhXAxKNkZHetDZs1Pa0STJWvXpc1yfxFTwDK
deGQPAoCqM3qNVhKrETsq8VVymjniesSIuotaakDX8Vew287m1fpTUyNkqlykSAU
E3TI9hOrSAPS9+T2DrFp7IhkIUficSTTrVU3Mm4CmYypw0WZwreOEhctRjcpYXe3
M0v8NppAKtK81HQfJivvRMug8B1RdC/9c+x8ZCM/ZOnLnT2ySMEAFfGN6mF0N8Kv
hABueoj/Z/VVFBJr/Y+d2j1GER9rCo1L3Cd0IFmTvMi0vDQiS+Ex4QpQ9tjO2d6D
2qggXidlMiEsnFJhWZNj0ry4TPoyoi2/PWjQqmQHiB9q2gkNKVuXXbQQrd/+kmsX
movYoBp5G5QHS+OjxbvjOKKhPcXyoZ5j3Gt1OTTBlA18MHvBhZEqiDfXMC4krlxb
YxhY56k+d/oRjJAIOAVV3Zm/uUwvrLkGsiwdb8QZwNcWsmcCIZT8JKcUwwlBiJoN
rRuf5XuGXtBH0mZd4hKG5IgKXtlB9yUk+I1DSO6E0XI3fmg7XpkYiND/b4GAXY+i
OaiBwasAZ/rz6JrbpFUNxCoOULd9f8GALPzAl1ddTmdRtHbTZVwlmSqjmLwrz+qE
m4ergTn2surVcYbZSBWK58mVSG1QxeaHQQ8Tc/HUSSUa98MjfGj82nuDuJ7i/2Wj
DKUyxm9B1O7Q8Rax4MWgyT/GeLdw5P+cLzQOHGQ3ou6fLfc6ToIdGZkNSvjcwCEa
R+3TE+IeZuaXR2ksVmRApgUpaPXyziDaQ8gpU4MszveXrafUz+tMjBAXbm0X+9cu
ZWmbuzYQhzdunAX9XnWlRm5AQ+/kx6JTmnK0s9cKcx78g8i+zTm9ovB3ZxtIfdXv
1tp/TsJ6YTqP8il2PBrVZL8WJnAMs3hJFUEWXy4u0X/jOB9YdZjNVQpF9QDPnR36
yBcRn6JMlGaYTmc+3ayVLd80NvGldyFz4lCw2yyGHtE1UeeQUBHJtcqstGe4bbHG
rKmcO6XC4/97xQnzBazqwWFrREfqLSt0nC4jNtYHIMTjZXIR739C0MW2imfHirRi
mXsAVKtamYihYSmQxdMxnDqe0b2ibWBBsJH5FiZW4AXo/35Dta+2rTXVwoqOk4wf
RdBikMwbEab1hIyp/J4kcF84GpilrlegsbXoUkrrUSVxLDDY6i5GHEmbMYEdRoSe
0JlbXF4PvUzjW46niP8BMo1qM50PlPB+UqnOlN6sKy8/IoUvQQap43oDOqJdBAV6
0n9npCJewJbjkiTaOfxS4IktB+iJ2QC76F2HEn22OImzue0w4z/7fAzPYt6aekpR
n53yVPxy3NUR54S+iNMOoswakA+mr8KDE+E2lHHXpUmwMdbzH2YkdLgOEPt2HY+W
WtZpyDPbQdTLxuNsrkVc2q76g9JK5TB5BvNfrzhWjkzaeid2XeC+zClSS9MdurQx
kXIo+kGcCjXjdUlU3wRxQwksE69GcIrhcntUgHq51ZmMPzyBo54OhW9+OfyeSl4V
0eluHtFGKW8O5wG0pY5I2+L4Z2nojtGYVW+9aGxASXz9GDwrp+PwlOMz0zQTj1Kl
GKYQCcNLOPHm84yZpEgsMES/wU5BWp5xwJOqnSk8RrmtlYG0TtU4VNYJHPLrENMM
7AHSz7fA5fNY/PinmSEcR+kwXQ9BmHixFxARk9bKEWfnFVO6cUd+f7A2QPcQiSPM
co28KR9DEYhhKHJNEOjBwaBrPvUDHBjG2oLegb6zM9N0qGJdbzPzmKXJ9JEL4We+
amSwS6/Jei3g+0ZzwYO2TUC1Sq36oglytajHD5TauRaCdd4LkDltDGX+XoBuRliR
dv4WHEmJoy28W+v3rmcNXtLw44Qm78x4pIganYaLsmnbrtbFMsZfBxNRVNdjun8S
l27GotsdMxJrBOmON/eftggg1Sg/bNDZfARWFbW3rOBlCZqvtrCety/hxnieJsDJ
rr0Vi2om+wB0G5icCOAm79OqemIG6AclvBwVh9MTP8wEANRLCXjp+2Zh/GQqYSv2
9CTNk4OWNxqO9IdCU4uqVyw9wcs/VcywfxJSQDxMTkMVpEaZMoVehBG8uiWDhSMJ
RHUlHEIMxaPF661TGxmszSr83yxP32oM/S5xLYId90j8kuYssp6HfM4FFErF7szf
Cb5b4ycB+lAIAq2pRk7NXERxj7dCg94p3XGTUa/PVjD0lhEiBEfyTBrg9NN5NDTb
7CHIVO2w55yZnK1RJtK6hpfCOeScKC+4TG8g8aE22Rcz7YFY5KyS4ioUix+fe17y
oWXChFfPpGy2CFIltJkyaODKyhJt+b77LNHIH3UQ3ekVzforToOBuBVZZwN/fEdI
Tszi8Yd5u6SoWKzsB7nxuGmGjlEBNijdaj+l7zm13uB67Eu80AzPQC1As+Ini4h/
gpwoJuK6oY8qelAMG8Vber/UDZjCeqpnwuJTM02RriUrdwFMutgJwwvQSEaWwtRP
4nKTRts7R7SFRK6KgDxl84SarNeuy8Ai8DX9l2pi1a8e/QZF8RuSIJTf607/H4fU
EbVxLX5kDkmOVC2gOl1xjM+MHYM1nIxvyRAdhNUWZOPO+FdSvyKbDcUwHBfl3IPE
h5b2U8wVWjJ1AJvKyHIbxKglSwA7dju5gE7KGb/QknvUpaNfqT+KzKqgbjO1xsWN
2y2HKn1xD7K06nGFnmzTtkuMNasC43Txm6bULFwhA6dVBXmneIkGl1/PBvyntcGe
1GHK4L2O8A7Knrro3f9yhA5UTuWhVH28iPv09o8aoJaje2lb/mKjKei8TA4vpetb
N5eEUKQDTJqUCzTHV/Os0QDbrRGvwczFYn4YSF0AHiV6wliKhb/Gb9QsrKeyFiTb
7/wk3CcvQfyEl3ZaYdC/zJUiMeBVhgm6tE/Z+zQu8VDCiehD5FHYAchHgWcQhCp9
imWYI6qd/4ztHgft/RFxcB3meQUn2od5TbJQHioj5HNE4YVRgrbWfHJhasYmcxqW
UvCSCmq3WfekBoaXeX/ZKY/q2GjLP1KrtfzlwLLsKVced/PruVZrXcX3A1JizMl1
7AuZPAcvpMUEUOv/bwuvJXWRXynh4HFDQ/nMN4q8bfNarPeT+UDwn27DlrylD9PX
F/bGdpmsUHAknv7GnHd4NNyIPft+Bp1OxIXbnLcCbnJai4qNRoMWofKba6OvJUaZ
PsMDYDLtjlRmbAfG0bcUlCClVrm3GpnblhgsAte7S72BvVOl8xNUJYRezCZ5+5FK
OANKTX5hp5qe3ZvBQ0XnaRMqvRhL6OpTbe2snJZjIHzw/haVxL8zUPrUVHuyxCd2
MJvQ+ZRkdYctbNVie25l+dHMbBLpfbMd2gMdTwop0lodwscCxT7ILaAWpt89mz/f
D3HbAbokSbks4ODKdC4eBVImkIgc7AvQeVFY17o/VMaTujGs0g+teJzmA6Qqd13Y
AxYpAzo+r2k22fzz1ckb3KxhXSKDsCC4IzVuhsOmBPWqeX/ZhRPpbPZAGGFi3nQt
86qzSnNR5HTtZkHD5aGS+CeOfd8MxwIxnnqF+jobUx/xi3Y6kLleAqU5yWSEyjS5
H0gIcDN3U7QocJj55KR2mEQt9wdYQSy6Nr/pGFyzVwb0umEq2yOdlv5eHZr0Z3Em
bB+VVzbeHq8TxqH0+LVocAsj38vBgKqGUynt9a9TVGvKhh0IdCjO2wbofvcaN0UB
FRMSTpc07Jq59ZdnoibTCdxLhNAb6nZrcm6ny3wJEAuOLYEnvzW7fBEiyJqINR+u
Gd1oy2MuX1jpDbluYwi/1SkfcWemlb12JQYCtZmG5lzKkSRMae756yMgfnkPnyBH
nw8NrZgFyv4FpGnHVzjxYy6IKj5b5TNgIc9717Oe8v9JuShM+TuvDghWRPQ0YVbh
+hkr+cxR++AXvdtn27/+tU77u7CkZxGC6mLL/xXbPas1Bc5SyoPcmpXoMJnzndSQ
u91MwzTleVqC8hy9UO3ieiCAVES0wQiATd6vDHPTqOjHwGX+6pB4Y2uNSoX0Lfyv
DVrxHGI1pmJg3RpmozFn8Wg6w/wfExCTrPR/51eXnW3JqA2u8UNuQMi8VSuPrLUX
0rbxvWvTgseHq/1ZFUOzmA9mpu5LKMl873W5xVowl22sk3Oq0uO1UW/LFhZ4IsKg
7KfLbxFEYiCOhxcDYtH1RX/+bE6NWJVaeElxgxuMfUOMJWVJ435Ymmwu2FzXO45F
VVV97weZ2WxnWoYrw2k5uXdBjWpNOakwuZ4u8fHv2CheqJmx5SZuXcC//9H5CeBV
YNmCI+kJdm3q7Nz2ksqKE6HHL2JICau/r0MUlAju7CQlWSThXRwEjcir7nPs+/JH
d07Lnf5K3gKTQ5sr/jBzsrOIqmM1bpGD4w0n2UudpJBm6uDO+pAtrRktTr2HMcuo
TZmUb+J8asN3NtaLRGEpRQuBa4g9NUjRtnfwSAtKAiOGLbMMklzDsfQrOe7MI7BH
Yx+BwER6xaDUP1EeSgWJtAyDVg6PV1tprJ8MDsBWJUVlFex0LPNoLKhmZKdukJqw
GUJdEYmTEQjwjUqBeSC1/e+pVB0bZHTAfOq0V9aP+gADaN9LzTr3bXg1K5a91Smy
RrujG1kRFwOCcaXQ7ugZ/Rq2i5FZvabzbjyO6EJwRQvDdRndQmliOlBNaN6gOMcf
zI55vREWQzmxTSNbgVBnlqRQw8wls0FD/PAXdLPe8TtZz7OWqfEtB6ErC+44cp++
pAcz+prAG3a9FW7wf85nX3p7km9VXIlgCeXCTyuSYyYKfapyPfiTREVpSSLyrhhS
FE6rRPNbkzKkTGflHXOshlInf9t7Bc8oMEEFdIQjEW6SdTEPq2NDjY3NhmYnU23J
yaxbhaAOFN+f1N1B6zJGlrnnLSoV/bZzxMRhInDjxf1IRdORhT4UlVOXn9ZSBd8y
9EVHbunuKpmbKvRdGgK90ysMlshHHAA/mKbrH1vyHNKNZ44pY+Lvkdeb6BcvHkU7
hvzSKNpo84M3e0ogN6WPEZMXNAjLaJChSe8+tvgin7DPpZwqYB6C2EBC89hirldc
2WPl7bbvOFtCDrjTA9fIJ2hc5czh7BIK9bUloLFHcTBak3nh59xIw7DN6Pif6iak
gdqsEaCvPSbg5IPb//D8Mk9n8N8m3ipap0mq5HftORhclgoe6CHg4dAFLqTYzfRN
s5ZHdKlr7f3swjg8MThNXOphenZDs/7F8Ob9g2tLE6kGbB9d4bq9rE3vD9W7ClxC
zePKVo7PZixKPG6liLx9zyU36g0HgLM3IUv2Ib15BzU2pdtcSUfQWfExxS9iq8Tg
86IyY5qCRrcOV3GjtZM+8EhiDelyds4GcMheeoY2vjq1MDhaGvcw8Ts0phkTGvyr
u/Ib+1tXzae1pOlCaJDJ9gdJBxSEvjVYU4sTvTKZD/GYwFf9eyLnrpZ+mxoCxJot
Pg7LPCI8TSVcQ+olx/khucCdUI7mjIDP0XqfQ7phbJ683ueFWNr38MTEUR6fnnJS
b8KRO1w9y9CuDb0XTdNl3L1AiLjD7AQijJlV4xLqJbMzsTgSVw/1xPsru/lXRxlt
zUgf+t2H+v4QLLuZM6Nlf1ZuMYYJ4GXxqn9RgA/juF96HrjPWacIaT10VFSPFRXI
F1mSXPBtHsieuFbKsj3C2t+wN1+kfdu+x0oA+R/6A6f18Y5OcTAFO1mJdzaaNx1m
HGF1svb5924u0Wmq3yTSfFFcJDZR48q4DyySIfGBPt1nLQUHOPVDQjDk1bhLDNpy
Lu244j9aghZAPJjDc1mVIC9BHAnaLRr7TFh5VC+unZj7feTgnhoV3NdwShW6Epcu
TRCGg+RVokE+ipNA5T+esm+eHtwYarhM5ZXv29O/xteQYDFASnOPqDl2B94cnwZQ
2pWuvnLq6NZJDzmHSZ+tLO5KmuSnaqqsU2p7E+Vf5cXWsk2cJ2WErmPcV+Tg/874
WepFTlz7FaiyWnQ98i0eOH1VC7TvrJnd+VU/F6xTMXm4PnLcnzNCTcVYWtRoOHMo
26rqdoCFu1kpGIh3ZIhx15UpVKSwPyI8KYMJlbhM3Pjpn3djA+s/CmZS/PRBW8ik
gZ05QGzbSNnYmnJh9CjRvJ4KNKMflwA1Q1/b6gyHiDk4q4AI3XZmOFLTlQwFVRvQ
Sjep2FjYKKSiPwomyZcBsShfRZ0jeCZQEaD6svdoo3d5RWtemk8/iysuqMfL6lTa
Tr4m0ikCifVweJ4kaoTMXV55bkeAfISSByFbylUr/9XOYrlyjXpFVXiiGvre1CbD
ka71+YTmXXs5FUzvamtb6B85BTr0EslSvSDA7g5AjnWyawpViXEZWkXW3Xr57wpl
dluV7QYLsoxgBRzWP7hE8JtvPZZkOq4EphYVGwdZ1FeDs8oGFJSme7QwV7UsRHxP
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SCcIxQvJpcWt/HGie0+vmnbwqjUZFhIUHmTolEuf1oXiRsV99Fn4wBvHQj/wcc64
0BlfXanqLo7FySgr7FvTiZfHxs5cCMXuLesxJhTY+w16PVVYIDMxsvrASOhB79XP
F0Qb/mauC04THtrsTwY9cEBuIY4pBESxTvrF2EkUMraoAU/srWQFdhPPizwzZ204
NHU8OKxtFA4ufUF14h18gBcDokG+0DuwTDaa5zDyrtY2YdWZYUQOt/UQstdtzM+X
RI5+XumaDhs9NUgLyfAp3xijXmEbhD5Khuo9ZhfOF/MrpreWH8KJr79KUXLEMhbO
pUQcX1fWrMnoUWXBBxWkaw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
9/0WKI+pb2uV5iQJA/KpNCTLL4J7xf3rtI+4ThEUPcq8nQRmXPbXQOtlooAQ4tiX
zZA5GoxVdz54aPjkwQCo2HjtZYkUBEwOu3o3+pI2jMcK8hBCFdjQUXTlTmwa6fRB
1Y/gDQxwLqz0JSTW/pmx6Gx4PM2v5pp3aRkoscQzU773neQbgtujRTYJa0QvGe06
OsyDqEp08T0mCXhxr7LhpWUDog/3QfT/m3U0fX9qrqoHfm1LfeQivLmQb8wsNv2R
7igrJglEaz1/lqAx+v9QBlZWVKUKTxcghmGRB+I8E/Nkt6lRgURVAySvZEu6W0h/
Ds/i3LQ12R5vH2RFvjBFFVEtlw3xI2V88gRN0p3N6AkuTrCSxMZhiPyOt+7tTlui
R4u4f7hvoS+G9xSfH4nGmnIjnmxxoU37+DFC106Iwl2oWnzyWqrRPDa0OX0vjXRR
NvmPNkfaQoTbhXDq/nROVxpxEC005Gj6W7MqwPHOzdo0S3gR9L3+sL1hR7LEVx2b
DoMa8hoQhewDQ15eViRjFesgT3kGYooKb6YakLzZ6q+eMkhNzoCgauZ8TueOhmFF
0Dy08OZAIlRXHcuH3UzWeWjb+qM1ufnIrHeCfZC3VBhh2EkSf7i4B2fB1f4XdUaf
BhUt9DOHz+tzmtNUiluiC4Z/Ia0ycMx3jOEI7f0uGflCbbZUTWJRssT5kzsSyMey
HBOzqOWi1qthg6PVrnAztUhUzi/BQNGIVV/qpRIMfo16Wi+HJ0nYvsY/LTb3Stru
zERIu/CQ7u1fwNdjaLTLDpAC7kiUQ+YAz94+Rb8cQq4jgxZTc8ftxRYiDdt+ss8I
2xgEsDXufRWXdY84K3zE8qDOX9HFw8t56xSftjnvaCTJBmRoAjk0jSUwZDscQH2f
a3TkqRlUeUK8wiOq8Ttw51+Bf88Vahq2aRtlR3/7m8qvt2zSt8mIjt1wryqDzlDz
23cHvcsv8xH/2+dfkaPfugbwT5Z2YMoL+XAneUu1r0Bj1QrPbT4NACbI8UHbimQW
5dNOIe8RN++FHAHyO50MuO1JRMcy96H89RmebCx20pgskzmWOsXQ/VDO7e3VPSPl
+WNWbil09lloD10K5Ul2sft5OmRALT7Q/dyXPIDQT/sDsTlGWvhJn1fb/Wd0FnOX
o7WGUNtBUG3cSoII02pVoNcrcJE5L0l+AxuBkxQJiSsZmOToXuC45yOQ0n/VgQEp
pYSKpfp5UwVZaBFdBPNoIL3bZ29dBtLbxFt4AJPiJv07bV+nlVkiild4ocESxUzr
GByTvN17MoKxoHOLrW2xUrM61ZDF0YyEfTQOlehUXVsERVVc+vuttuQEtzyRyQdP
dfez+iMDEcDQp72Zr2fdeZVE29RIVuTbxLgfI/wOI7wClmVWDy9B75x1IUGSeJbY
dt5xPKU8dVQhps3fYPa7q9IoMYl1JtAsfPsgwie4WdbeGGNFBUDaWz9+3ulLljxQ
CY//QpPWInIRAtMhhNs9Wo7l7o+az1mXMjaf1Z0ln8uxgl3xPkugjHsekGJkSxWA
KNk/qqjjHy3jVU6oq3MzSQawKR6E+O0e9idd8Wm2VKxod/RrIRu156V2Vji4oKsH
srEzlOjL2REPSH0xh5yLWTDXlDKLzApx1ilEVkLGJaH9e0///MEpPXUzh/wixgl1
f8ES+mAhIzP320RsPIp/Ir9Xvs4yiq51guL8+LTa1Tn6Zt/p8ndKyZVbjN+u/RQ9
cetXSP+4+mxJiXAFhFbkd7zBKiOlvQTwRzuCr/4MtrnEVgrxqUklGKWZN8u4xxxa
wTgOrKE2sIO7TP8/t0gFC3lKVdRc1VU4dE9BMnTqw7pAB3lDDybdMHfl1dp/JRI8
ZQ6vwvg4APp1+RTlFCM2qvtoUl4cW/cE0eOCi7bENcJ2cRmxiKpnqwUaemArIUpI
K44mrLzcwkp9v5igSKnThE8IV8/xdTCoKP/UXUhdS8MEM3J9aRYZiSubdAR6aPC3
niQ+xUgUwXT5JeErnw+iZNm1l20iyl6EZkl81YxgOBnh3+9ljRFQ2mBDSREBnsZh
1ubbR0vRD994H4JO7yK2QuGidMopi2wQdhD6yC/6lVZtjzFyMhClwXqtafcDOeco
6XgnmhLTOksWhFszH9gy0sK2exPn6qh97dp4iLzfsUcAJNPZ7WOd/tFVobNpMD8S
h8CQJuqXyWpiyUicrrHqBYdc6/lnUMDUrUJzw/YY0E2Nx+NByiuvy+vMYa3D4SxU
ZJ4BMcibMcs/KWmU8BubajoULTCTW9pj0+AFtqKkzBVDnvDK4j26LIzD5/kd0pD8
+jvDHC6ISfq/tkqwP0h0LsVox225UAnv9dMI80JDddDHri9LLFa6AIDEPhJ4f/X1
sdQiLywTE4D5Lgr4U8QmIbNwHdxyZPlRtVJ778Cs29Lxk4a+sphghZkymtxgB12R
vfJ1PJPQSr13WwBzniUTk39th7pabdZx6BZITePC3DZMgeQ7rNV3IEC8gAU4dtCm
DwI6A6TvLxANf+xnVfDN8nlx0UNN0oc1ZOJMkmoaz+IXvlJyHvc8y+156w+knflg
EYv+hktc1jMX11hJf3yHMKUfSwv7PpHll5DSW20ULOht/xOfM3zVF/H1DgmLuxDd
7ePTLehPagzJniPRXrE476QDv7lrlfXRoqg4sKpRvWeR0Yzk6qoOu5OgRdmhn4N7
5/MMGz5j9EMxY0fKApPa1eYC83NNOO9F47ZbWmiaYcOnxIAUeY7oeFiwa1DjV3Rf
JRE+og3+xk59y/qWQkWu1W5JPjeH9WY0/a3KqZPHJf7YA0dUgszovGm6b29khQGS
t8pyxRolsruww39IqedVHmr/kciPf8Yd1l6pNySs8gqCAr3dXFeYhaFh1Cwn1/vf
VN1vI2HL3NjWsT2Msb0iyMjXsDUi3l2yhTPSTG/1YykcdmEXx9BIbZRWkO1Y3gSa
HMwdlqABbdfH0ItAKOrnnUWnvdZ67mYkiLOb63VIOs5c5mcT3yxqxxVq1iWp0VDy
aypd7SA5I3pSv6M9Scyc73xWcS8b/+g47pJDrSekqgvTUg5dcPA4xAq+5b9EyUdI
Rmx8ARf50w4OlB1h1/g1MNTxPxSuMGroUbcmqegbP2oqM1nWSmHTpZthfO+oLoG2
T4T+U1TrtmDpHvw29nuKauPyKFjAaZGlsinlnJDIE7OE/xQJeS6n6hk+c/AE7Lal
9fylsxxr5qxBQsj1eZIiwYbZ+uVsEQsXCkzuxhE6XCUCJMXNjBzwdp2s5EZ3+RNh
+QyFtu5dcShAZQrDafHi39U9t/ShzLjSfb5vD0zGpaNOOiNtBjvl0U2qDqyVkG1w
pOEmfebKE0hFPASex2q4E6qGxlXs3An5oaHvjc+8b+sGXKFwRcJqOZWVK6tddVIi
NqyIr7HOCD+xCXT6oWZDZ3tY1mswtmiyrwYWziZvvBztyhx1Xz72/RMxLYfzOf5g
7TFjemI1QSWqL3mE0elvqbqkGgTFmvYhNnLqAmhmDhkwmutaORUM/HJl8N9a/he6
48UbSyMiGz/8UIBmMJFlMVk72L1ETO/VlSwctXF1pM73OYZEDVq64174xcQSE2tL
l3KNoN39nn74y/a9O4MwVuRR2mvWfrR0S0CwGYJ4DAHYVPwZB465bOwKnRk2i8eJ
WVrMJMcmg7m0qU/5tl9qOpAik29jpxnDi4NRTBiXVloYrKsXePwaETNoRInxCyri
7FYf/4EGSCfm0X8Atd0ux6x+Gw27ZKk+Z/qwzN3DH+XPg7vvovYomtHdMvQSXHbM
1FuOFfP+G0WJKaC3dkvrga9D/a+mZjCyWAOGg9RFo2ptVxVmcwamaFH1lfh5YkVx
A89q1+sJ8dX0MHXx2yFUI7ZNwSptsHDgmyNj1I135dUppe0pR+2anhP6wMYh7/Dj
chNbje+e3/xeT5x/A0tCWF+KmaB9aU5V9vchLwC+ao9S6ufB+W90ILTAzscDcwf6
aRYlQECfIOCN6dDjatj3vrRvxdtcpI+5/a4da3HtkfImEnulTc4Fb19el+tl5R3W
4Mnn5/Qo2UcXtvgAvAchSRcZfWIrAHV1s4ibUsQ8ecwPDG6C55HjbXLPlyOXXxig
oz7G0WlvM15ZhFA0eyvhDDJ4uWFxTEFmLHJuyfxnd0sRcZz4XZq1nSIF9qlm5HE+
pPtWagbtqguKxwfLjMwe6vbhJwuSnE6YhdgBtpDHIDefH9UhYLgqBZIaqI1fe5Ew
wl0vuIsN5bus3lE4H7PJ+/Rk9TBo3OO3KTfBli+jXIlUwx7WMm7y1KMQb11OAjYt
byMOweTX3TAtS7lzy+nsJ59JFsP0zWEKTUaNTaIUvC0u9TDOX8Lw/GiP3nrsw59j
Y6L5zsnFc3AtbeZ4PdJEYL7YnzxxEvRUGpp0H6GdfDO4d5XN6TD7+dT8hctj6hDJ
6r7HMydQF5X0Miwt007AC8HOumHZa7+9wh3MGluByGhkM1bm9cbgc07xER9LIwMn
qgama7/z0bvrSsku4S89lbcFuAMxhhOXs6zv7613mtZveVsxj0rjnXRY1emWEzs+
ymXT1EKzCcKfCM16K4QY1hGJxPX5GTss6tRBV9Hnkba1KWRGtrpW6CtucLQdknZ4
x0Z3pwlGB0VgQXt6Z+4vN1Rm5uDh7rBXOzxx0Kd13cgurx97rEUJwtmYf+FUNlmh
1lID7xt20I10VgxJB5CBlrbLEAwaJtgWoteS/NvtYyD7h1OBSsb4h2pxke1oR+ta
kII4abzQaXnaUne763Zf8lDNWsPvJYvx4/yZNOwdXk2k1wY0f1TgKr+P4Bxe8s14
boukBMB2u+2uul/ctgJ7k09euMUfb+0nhab4C2e5gktC+ke2AIIz+ZCHNl5Dggmq
+XIGNXxQC/+drqTwuGzFd/hrw+Glv/YS1njJebpzxY/YJ+Q0oUAZr963Rn0m5RrB
8fronfdMJOBpYeCWhR6OoFfast0ZEiOUl0exID3GvdUprafS0hCRG4EYDX//xr5p
k1jc98cSlr98x5tsuyXRtdVpx4SOVUZGQ51IMz62bFub+zAWcGmlDzKUb05gTP0X
wU5hu8ELwICzTSJftrgsNKgdroGxW988Cq08Yglm4PnNYEoGoHGlxhAWeIh0iB3J
snHTvI16ueCdB4Z7SGe0KiQBAeT1buoR1M9la3714zs=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RUx9WaFvhMDCKLEXcfOCsBF1/0DOepx5oy3Bz/dLLNcPxmc9eI5KJFF9+9FXsQml
qqZWH7nBw99lIiH6IVjFRucF5mu1KOIl13NWLg4EFL+3JkA7VPv9gmA32jApJWlJ
lsIG6o8PnEk8mkq+VqRm+SjjbCJm4pjzVAnmx/FbVXhIvfJ3cjsKZFPUitoqcITI
ObXyxlphK9kZ9IEl+eHGeekgoHyPcxqrzrZcSqhQKmcvKaq2OEu2aB1PGVypi4IG
SHH+Ji7yOKW5U34rkSB4iXveR/G23uk5+ohZpAbROYuox6O1fD9zRnwFf0ntpkks
aChuTcDDpZa6W/IgtI0O3w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8288 )
`pragma protect data_block
QX1aNwUFVKluWYbmurfzT8O96R7nkYCY6oraimUFYsStejDKc3JbdrU9lvNgywmv
uV9z281EWfEV5Xi04Wf7Zk7j9p3ykrsoWZBxX1C+w0W9tcz2yR/C5nPKbFpyIZPo
sjBx1Ob7bZAP43QkU/kmussXWOlOSRP5T069CSOZy5OR+2ILVZGltsiFqUtyWYsI
tSadZIj4W7yKSrpGtUeIndbN9lJNL4W1ybmwaZUc7bplZ9/QkF94F2fj3tX7UbtD
nFKs2pL6bpfN8cX2d+5aGjqzbvuAqgrobCtFFtihzw7KlEDshO4x/uk90oKoYBw/
nXHV8wjKGk+PUEvasQECVtAM1l5EMsQKC7rTMDRl3AAp2OyJT3CRMEZaTov7FNqW
wfh6J5/13751Z8PD/FlS3HADpIqHCd0V+FV9NbDeUcMKW4sRl0d16vCkoZcCZcCI
vYSNhNzFYxL87/myoMFyyw24uMT0hRiIPplubmwiS+HQ18s/LcLFfA//kwH7qPAY
rfKbY+z1CxYPBSi81p6qwTzs9lrSAhGYG6KXhTCTVR352NgpwEi0xBUMhqiAfrNh
LQjyl+OPR0MJY6jH8XxYe79ESbU3KAjq0tRrxsgpRfcluglVJrLbc8uRp43e+P+B
qd/C7poqww2R7BxMR8jF+VvLv0Ysh/fzhWBIqh1Cb1SmGPHLA79kYdw2WW+ifffU
vv+vLITa9S3Ydji9/gWNzHgbr3B0Al1E3sk6DeFmSVs36b9kb0ZY9jqmBp01+8xM
oyjtdQX1QFNlA4cM5Hc00IB4Edum9Ft+GaFS/SDzWJ4CSSBF+n1r7rbgBd2NPNDE
M/GBFVhknTZLQajuqUSetpvwXmXrDdtol8zt3PQS8JatssdI/cM4h7KAGZLY3xfo
FRJsBGalT7J2lgI6206nSoJg44/sshtwvv6xLLf7d3HlZw6/zef01nUb3Q0NEGWO
n/lVv+DSg4BQFi0PHp+Kxt+X8pjrtnKZEyMvWKhqaD+ZQneztmPFwHov5LFeTNuD
p+/GOW1fQQxV1iF5eAA0JnxQxCyckFl4AL3r/lZN0d1XaAK/+lz6ISoYRnsDIJzN
1z0oZ3S0RecG/4TJNdRi6Mvwd1CorCZ7vpzwAMU+KStvLrKpP+o6+5wZYtDaMEBN
TocBt9SpRrJ/NHY5dg/G3IemDtDfIukg+hXUVipdIY61d/ma7cHglrz6Vo1rdXvK
WHxQ/yBa/S45koKLP1/+12f4MkG2AwYqTuBmlZSmE5i8sNhe1rFFzwqwB43VQQoL
aPVnHDCd7+Qi8B1L5hPyWFGZTH/sjAayeN1zTKp++/xLsIEPM3QjWjWL/NTnP2hJ
CuoY5UmwnIJdpg80Emi1ztvotmNcT6Nv/yBaz+pi7g1t43SLunvOXN014GvJ0elp
J/6OtQOLl2ShbpUExll1GpBEyzPWYN5vQbGG13g4mQwXXjbKG9+WWpwe4k7rNCnM
IoWpO6G1zJd9ybOrLHEdXTV7uKZk+ufkJZPrVvdkbIZ9sqU5wT5o6hXrfQS4AumP
Cc86uF7EU3MfMOoKfJqi22F43lGzuR/33HJHYuETaiUj/FfXQ4KkpvzSkEeJCSB5
4RUVeW/mGmOJZQnfhoNZ93e7RQ+jzf95W8xB4afTK8qf5e4yJrpWhpaX0aj0LpUC
SC/6r22eMxCwqVu0ZAdfcG9Z+yJEbqUirRdW1mYuFGJAE0IBKKLe9tDP8MKpnZJC
4tiI+cIWcz83f8Y3m8cPEHA/KA11Ct06Od5Kzc/Jt4vvNqCJbJmAnMrA/90JxWEt
FiOr7VC5jNyMLvaARJ1pSXR3dMQcqkbQje9IqEJgm2xYFn4VC03Qewul4AOXLits
Nd13gd1QL5CIFtcv5AW4FBa1PBFUKhQ11DaYmzn69bdyu+7Ug4iJFDkiLOlRsj5C
H9fRMAYL8McCc44eh1FtGOPMmrl2dLvXwQi3AXYVdkfdZbFLLv1Pe18gb3bJNMSw
vhAvBDw1fJcve7KZZT23iJrf0ooVrOuH9d+T2nOIa+f6d0peqBU0ZgLSnh8ORiE9
svhzr5vaXQ3XJiZ7oB/YS3D/mDh9UOTmjrIiLQoaNsLXKzOT2THPQF15sKxSZuXB
G5gu3kIBXTaIo2SIcxTNCI2Q6gsJp+iF1N1Iea4PeylrEga0i1gLp78w1m5XcTH9
7pKpi2H2VToCsuuS6lvr+HcAJ0QQvDj8LDuqvVNYip3ZfJs1OsQe6FUxIsITA6LG
mIO2ikElpOCE0YpxNg6gBR7K8XaUVckAtVpqif1eAWoq6hItfK4kk8XXbjZ64O/m
dJoGUrdkz886XumRUp62YJp5m8sg6Q3qKpRVkNjyTnWfnEPtkqA9h2fWoeLT1bYq
LnUUi/H5vKBPx/Sg5dMLOYE4Yoc4s0/ohIyb3IdvhDKvAyPSI6LPOVsgNvYNhlqq
VuZA2AgqlImpqltiJrkHVWWy8KDOiQvUJDTP1aPssnKbM8STO5BHEoWeWfPnOIJw
WsfeFyLO5KM2HEVqjWNA9Kx3LyOvcO4J4UigQdWsOF3a5RlmUcYF7g88ozvMTcU+
b4lI2GkKwxZnalj4gUUKJDV/hRnP3chypcNgBBb08tfQwytRs9jUKKRht8rw+WvG
5RJ60BbUomf6u02Du/x/+AnnhFD5EWp3xvJUHKyj0y9imtWcFB5vHDCApnipAhfH
+M0bVn8hTvcQE/K+P5qRE7uPpUggp/1wliCkbr4dgnx2Q/3B7/y6jruaZtLG7mrk
YTJwWAjiDUH5yZpFSI78mEiNvz6wk5k9IEWv5BWrL+bhJo1sA5WOWGP+R4sSJKVw
oQoEBQqOngurtM5tdY4jNm380xw3SAU9ZoaZfefcDeR5Q6mrVd2yFNxkHTlaM2mc
oXqNtBci0QUz5pVU+ikU2OewrOxKDwy+y+TNZwQXGz/7Voh5Ym4Fqe36pIkKlRTJ
jqpLD539jyv2rj7WBmkNaiQFfhGEIc7oDLzmFamXBd+q545SPQ2xKNS37rfmr4MW
XsesJ3WQpZeH9CXjH0zCz4BhQIM9dX+XDlzh8bk6z3n+0VHtpDzpkGVE1Gq/YN5w
2rDZFzpev20U/3LXQlr25dMGWNc2fZNmi9dmTwX9Kt48lhnOmpxscMH7uIPz+ZgN
YWT4XtmPt7SMug2Ehyu4oAy7ghOUMuWRbAjyy/d63jAQrhJ+SRN4zcjYc+CoG8xM
TgDPZuO2vBtFqSxsbMQU6bbUjqgEpShJkluQO8Ix/mkWtyief7KkFvFHPJHLl8HK
mtN5GBYGVkruTGVSRu4h30ed4QEMwpFLBFvsZXvhvxKsUI0tZ1BJqUAJTgLTFINL
NLihVdMUgb++NCVyhY/3FRhSFnZBWdxj3nlF2ibv2/sPEvPrGxmaO2waZ4o/o2vq
weZlvfcIkh06CfRsMyxKYZp2LTtUeo4vNx9M5BEEjg7e6ioT6symy/fQXTf43gzN
azQPfIXcPzs+0GllB0q9U8NVCV75xtziRkOkso5gI4We3tzv4UoPY0Iu751y9jKY
MljueTg/yfhsXj7bpDXrcm7OAp6PHBr8lOoqNVX+nZ1J7WGIKNYN9KGcnxadq2Cn
NCvs9RWeDQx9/+zqgt4BlYxfXLvmOTLrMZjT2yY6GIc+DteNnk92G4vGMbn1Yvu7
Fpj9AWZMhPZ0UbYjK2O0SxwBtbDxa4xVYu37RJZHWjFpMWcQIUn/qplPrVKlWcxl
j2L6ooYLnwi15w8fHci5hKNK/LHGKFD4rb7WGp+L2N1fXj9YoMNaGR/0kY0dcIsP
JtiyOzA/NdB15eBIfSTKhZNQMmhmSzG2AftTKg6nn2NO/nsaXExG3DbGwZLs1T2Y
FhLn7sjhrpX+Sd/5lXvBFg/9WZZttvTA65Y4V11lc+XTLqmW1n/bE0+DKVWP/fYN
h8YuLt4dUboptJ+RdgimIN4jKx8JgQqDIbMcRjgM7rkjqL1x/OCFdgHKjB4qIxXR
o2Td7rYx0zASEElMiRSqF/chMgL0H2QWXlNrZ7P5/XCMqXlWaFM6O4EpDmpcfNf8
6qllSJlXRqCPx//ZVmmgpRG7F9a0+B9w8b+8EgTrcMyz70vYtjpcWuUI+VZGTL1L
P7g5+uinUT00aN2/pCdGrEOD3nT7njSFzOJ/hU1QhCOB2zp6RC7rdYx+T4OElUVj
i6J5sxuCoOxGnKU0vS2WHSki/vVuSDzOwnHWHbwyg2mKGwN5UQhM+AEnTm22rV8Y
J2064W67oJvonAUkDqhNFEwCuNFhdhn7xE/5NbhMQ0rIrm1mzn1G1xrBcSJ2c5eS
1e+f/yW3pCdgDmmG6Sjl5o//nFtHOUxMiNdrNiTQR6ci/psybTDUsqX76PojDKSc
lDWLqtUtqpIkjuSRgAjxTTwe2o7yRElRVGMhodqlzjsFqV6XwoqpKyzLHrCn8lqI
1ReJWpnu0HXdZVrKAgBVkPVzH7UUHwHwywfTQSZz+MQMTjOPN7BVVw7d0+6V2Sin
ESWYio86Fv+GVNsmeUlCjmMVh8klxCeWI4h3KNmpRTzvol8emmmb+9fkv/l02GUX
byPhGpxVgSmdL6+d5hkv1jsR2jcG74CbTKAKpHggUesFkjenMfOm5OHxzRN8AhEl
dARHscG28+2GrCc6ZxA+RZMu+X/OXgQiJFhaDqXOoxEn1ARgvLIPtpLg3zfH48Ng
2uDkcSdj56fG9/miRdn5MwRJwOmgE6jU1oOP+/vtYocN3IDyjeXX7bluT91ozUgh
GihOE5GrDO7GDIdJPd+OXLS0v1GoCp4LaWIUSpPk084lTRX8zw1HIc/VKvVrLmN6
KSD9aGK68kmo+ekKTi7TPkDT2+ySqfaT9sF3pQNP7rsda7BgZeZ+tyzkjZb5S7ig
Kpt5jNIHPCpKbIcFnOw4UQtlnCFSd/swy/fO7KS5BWn9P8V/FoFqSSZJqABLAOEw
AO07XJmXnBE+dQak0c+5P5GXxK+3F5N6mxGcpX4WZj08eupZgc0K2+6IUTHP+yWs
lKsCXvS5MwD1m2pCpfba8f6EXd5nv6czB1kStVMGxgVMxtKA0kmukX8Xg/eFc3IO
jmA6mY0bGLq7loh1oLNBFOCttGDcEfqXwE45SDdVZGSqtNjuz/ciU/FDRnU+tURH
leyjqWNMOs66nap8juqZpYl+SyZKSvTdsDgKARmQOAL4LT14pQ/I3ITw5Wnr15UH
ak48KSt7JjMdkuaLYx+CAQDRXAaPsSvoShhVGpCCVbvOAg4p1l6W1b2Hqnnjh3GY
X9cgJSdURTWz1SGbWrSIWITNigw+qrsafGDIxuPdKK70i51ecRph9DtodK6jQ+o+
qtBypPIwb6bckqCSd6wCaubQna2Kt89SP+y6XnbyE2C9uBTZtY8QFMUTzPa2e+Fz
ZVdQvsxj7Qfl7owxnWFUK6lvcczSXTpIDXDPRVl/irI4v920pIC4ZuxQNxI1VDQM
VL8b+oQzjYX+PGVg9zZO21VfL8qhlQXwVRblmTWrID49Gv+K2pjUraMZ11s0ST4T
6OnZHzt8hruJkfpTxeNH9oql8yJajWL6UZqiHJfDfwvWz4IfNboo2V05Tzu3/CSW
dGRYTddVdQQiBivLL7H5hUfuYNj7KLPAW2XIoKM5PMeCpV+t7PfLHv1on7wmDdqR
M5XcvDyXtkpj6a3BP4b4K73d4wGRIV4S2JKXriKJpJOr83gyAICPIS/UZaeb/1JW
mBMK0br4/SKqpaoM1BVGEESPfjjES32v7pKJYkPlPPWesimS1lsFj7cvNyHbBWKM
eGOAniwn39gDPDJ8z+qoxtb/xU0OBDfZ/qg7NyAK1th9Ppy7fysSfUBKqp8oMdNX
Jb6AqdUPKGAk18HnsALJUZd3dvdl5zI+ZfueHTBdhvZwTuG/usprKKRawy31RZwz
hEBL5AZQHvfhvjnAjAWrcsDHp1FfL6is8ERFriWpYuxBmEh1y2nqOw1NgejaqFnh
3F56YhagSM5P02Ft6ynY5IYD0lzDTBf84i0iAefer51iMF+ov/DoWxOstZwykG5Z
B9UdrT4mKMNQewk+TCdEFltazw/FHPGaTxcrOqEnVJpo1GAQOHrrVPpTVL0Xqbi6
3iImJoIm2gW1vgOLGXdzFL9TImF8Q3jiRA853mcTqUWP5DhDndPVsbu56qOcG058
pTWmey4oSrgbME5qlTZtzBlPqVeV/ISG0TwFrrtbQwhVBrNmMcNiwAKNdjR0RjfN
J63/e/DAvw8mVkOiK6rCvERKiJ+5kOr+RItA49Sn3Inflr9IQ9dtxjsD3dOPFESi
yDnrPds1uG/JeMQUrU/RNI/kLJVD8pQA3l6gXOIV+yg9Kt+OAD2dx+hXDQil+GWR
IFxQKGrVMFDA+3mA1YgP22B8FLGfhwRDbPQBTXMexuL9TvaSHxs+4+hT0g5bsEii
rTtJMy9J2I8GULxIzsfkgVORPFPRqD17JNGfQcSiBnhsYG4+E85K7OAA2tlflD12
gURTIn+xN/HqKapPho5NXaBJGgxgXTD8T/XzAN9AoIvbOuK9eMvqJb2PtuxFnKls
S60TyG7aUpM+6JjCBj2cnmlhb+9b/Fxt8769zSAv0A7q11gnIza1wWr2MnJhnliq
Z7EjN/Wxv+ZyhSMMcf7YVAVHDto6UPBseKZPS8W8hywL8Joe8O9Olb7yNdRLDEp7
Yz88n/RrYfZyNvyjvyvI+YdVbxTBQeESBfIsqhjpDOhkGiXsQI7dO582T9MVz9dD
u8TEENdJ34gPypMCTSH2dyyPZhH3yGaGLahHnkaEKMrtc5M94CESE9PcSd314dhB
qpS/AWvVXSyPGUkmryQrcn3lxIDae5wWJlBBmS2Q9Anx8QTRb+bMLlDNYaJrdLwe
Cpy+bKz9IlvFprb7HHxIy7i2YNbcKiaJUxl4f73ifbv75qdhfKE0vcQNajq9MCDE
gHo7eg0nPC/DVDcdtULGXidwIDDtUyNDK2qFJpKEpatLuVOFGG0SncZrDtA4myiu
Bluk8sz6kD34amlktBOZqfCMzroqU0wvv5d3dNm52o61TSlZ5MPulGRzrC2eRcky
gR4ihhT1mjgImGrVhhThbnQAZusaeqrf+HiJDuxsnb1KbYAZ/qjScFhKuXfqyBIE
TLR6UHWJLW5f1MSjfaORLLZs6GTRJ3nk3IPZC/Dl2Qtt9WYaxJGHClXXB1+Mzgp/
obAfjctXR17/NG1Oj0u3w5d7LYhm6YLqjDDW3xApm0suTSmZS/C/Teb3F/SA9HUf
JTDb1WvQIA510uvM5y0mXTC4kwhseMr/wxJfVNBedF2hlbp7jCA2TYAoEXvLPMG0
QXrBK6Un90AatfCnJzOWrYc5tAvAvGv8JsNHLIsEREw2Jr4ONLtvzPX9802NnPBT
tMyhctL0YvKgDzz6cdx7pfoOCahGjNcqeE/qgn+ScwoPkauQBBnS8Qk/2M8+llMC
kXdjTGW4z7L8PC7b+4hYM6j35xWZaZXLyUkY9xtnqSpjp1xfSP0iWh/AmDhFiyXg
TNQ/pG3ZmFxwADEW4OmAu/EOWDQcOv0Bss5Dmf8V+5diElFBVAnMgSItR/F8j6wO
S34562NZLx9paAOfurMxlRyzH7whMvM5evuDgJxmfl+8JRWcLd9+D+PtSQn2MHoB
7tg/QWJH3prVUnf2KviBu3D5mfwXOaqtQ0XLjyVM7xDDU7Czf0A8PNZbVe50WXJv
c3YlyySPXt9acGggs0C1YYsfdWU+8weby+SxFK0d4Z7GrsJBwCUgOMDdvBRmKSni
f4Mts0E8hNFxbvEzUJ+noMjBxcdWnbO3WIt0HY1DF+//w1yf0+MM1APhUQI/fvjH
q8djaAwmnODt+neRudJqGrtXAMDY8psQnYyVyuGHVWy9yiqLyFcIsQx/w1A0aYwS
OMSUsqR+pgC22/UH20v5tr20MuwX2P+kF8DYHWn1xpBfW1RX+ElDKWTSP5Ah6jnp
8C0ioFNs+2M4fMbQUSUtYu6k71dfOFSe17qN+Ecs4pjIL8Gy5oNSMkoU7tD+GNMD
qRGiSBy5WxOEcchIkZs4WPbdfyeNomfeO9GH/sg3LB7OClvziVfqRb8X6zzpH6iR
ucoG8SwufmeJnk1NNWOwLSopoBwFUHsLLyJAzmQnqXz1xilG4efz8P0ezmPd1BJf
9eLzsXjLKRc9f0Rh8FXTsyVVTCo+9qaRVqJ8ac8D7dtbgEzwF7HUUoMiCe+hNj8m
4Jaot/VJLMdar5zu58CYQLwjUxf2uU+iLR6yWzRdgrWM17A1m+G6TJcWHANQGmoT
nUPPxbjCCSiwWfy9dOx62qrKsQ736aqn7wavhTgUB04H3LAxt83zneCCCXZrh168
FEDhhyVlPCBrG/aNqfb68VLmU8lJDLKiWudp4Bj8VsBWt47dwvn55TvraC2EsBnC
VFdCk2t+pAmoO84aHjaLGrQhR385s1YU19HW/QoyRJaIctATOm3Ej8ekSbghSbaW
jzioJI831rTXJ7tTUfuWZG8PFbFMIVWUU/28X6MsrfeB5BD3xZtYWeJJrZkWyyU6
65KJlSEvpa2G8vLBmvLDxjWbFSD3Rx+3bQfrkGODqIxnzNEYCLt1LNZCvfd5UPyb
q0Fgq7mdl+ue2P2DaB6Si5U5z2OPv+TmgmP54qfJr7yxbmW6VI4+XPyU2XMf9nJe
JESWm2CI/uhwRan3d4cdCehz8Z66pKrtPIC/bCFu9BHFPWXsZYXndtl/4Y0LMNdG
Fw1nY8R2lyp0KGXFb1kUdcz89Il4SC5lbNfCKTMcPvLRwbv5Z4e3TYPYG+/7eemw
PmPjPV5LT1ccgo6+bIyYRSmUyiPcA+EdaFqAPRSAuwuQ9utIk+uwv61acYN4j+75
defNnlq8gideGTedSRrGhxR9FPkdDirNfC0t00l/I7neZ3tyl16SvPhH1fWrkyzr
y//T7UCgP5XdGQY8P4qcAHk5w/9z+rs/IBE+Wz9aBDwM7jmJ12Zw+tweiiJz8hAV
jwcb/88hQchw/AlqFkr7F5WVRar1OnQLoSKSBtrG7o52WMtvYdvvtwEGsu/F1ypI
GXgia20zF7g+rWJqlzrPqjtJcaoSX9KmrRdR+GzF3se3JR4Nsxd1nxppao5wDkhV
MPdFgQUkpqxUqhVipfLKPM1GqFJl4d32wh+AaqFQmQJiUt7iB6arBqWGIBMrEvVP
IxPZemnoxL2YLCGX0qYgwZcFy8o91kzcPhblY8k5mUz/44sQz6bEeK9einWlRpZ0
gRphsjQHKMJ0SHCx6h/adr0Sxocu/NLQRVK7h5flP1AWcHEMyYV/Y5gSu9NYItQ6
r/AK+6dgEtinoKefA7wwO5I+yU+2Ge2L2b5XJwW7AAZGBcXG0EPMj7CvcNyEGjft
c7JlxVRlaPgBhXWE13Ei1AWBv/h9LTlzx5S8F+qnpMkPQN7dE8/Sz+RrRD8yEYcc
OpOHDidwBQpEHnV42hzqUwaMWemQO06xn3C85g86HpeLOzS9fPUxsBQu4zZGMDRd
Wwm5Ua6z5gk9GZwPkaeXqj1ZufYS1qCTtaWcIorjFYtE+myDBxGmY1BtdFAgd7pd
wDqwJa6gtZ/T6huz1u+bJp7JkwQ3eeiYngsaihKn4CvbGfRL4gqIkDFwmi9S8Imv
oE4YjEARwD75Pq1X1J+HB9oF3o1Gr8WlNZRpSlatRUgfyAIY74os/nivCY/W2jUY
69sFIaD/9tNzkrdof/C8ZWwPcqKMwVQ+9R/EqPQpHkG+XisxTM0quLrB1+ySQKBh
toBe/PcXCQjR2q0pmd/LcAj+U1XCGZQUxmW+oQZVJnTE1/VnAdN71qEbh5YNQUvz
4SqudtZmvDNdpAmucH1xiGSmwF/WiiANAly3CGhVXhCbgn9XNjiv82xH6BmNuXjh
uge5HpxXLNDUIK0Ef1AFlNOuKbamGY5ScJQgz1aIdp7EG5KSO0MzR/s7CHrTrPNi
in4OwHm05IiBoerUqCP7sSTFJ1AvJU5LBrrKClqo50stCcixRGUJdBn/LlR8H1fu
Ewio4hXq0jKZrhduCqsKUDMgu8ChnejhyjWMfQXbdUv1xyPpEbKnvb4Fc0o34uSw
gMFpfmI3tnUwAGZYp2ZC7VsnxkaVhG6OCei7UEdkq/o02BKcYHqGDd50wN4Yw4Ey
vF1WREyGPkCOoCTOmsGOKygmeHGLnDnD8nft/nV2+CV7GEQxVXFIngMOAccoA+EN
WMOsfBfV40p/GqqufcUzxRPKOWuABX7VvSLmDj2zNw4oWuJv98HSOya6ljn5I9GW
ptVi8htL0AvZUH9GezX9ZSzoU21pfZpxdHuYxuV06B0ZToBPN/b7SjGMaTTeYj+B
BrlZAkIEsZNZ6ArUm/4GfCZxsfEjTpJhJVZqOTwxa9ErtV8KlDgs9sbwvzOXBfXF
qnN0RkbiZZQa9tfgQif37p9C5WNZvwyUeExvDWxKLc8w5d/6uNK+s/ZAFoHfU1ta
+p2LGJl3FsjjBjZt+5FNpUhNyjaKgc9UHpkMuagV8yq8n5YKKg0btcYI1Z4BrDik
6xKcgeMHcg/XB3QXmKGJ9lzHUH4iLrLB+e7bmwi+zT4hbhp1IoyKpkA7NxRciZlG
kvjq/pAaanIM110tG6pocdvU5YpMz8kaBf4qq0zs/Rb8UuYiQeO9NUc5yEy8sl39
2kkqOkHJNYTIqWeDBmJDfQxDFDd5fgnLHdBjrf517wcCPNwtLCTCq9JfsUkF1Hg6
4V3L38lNW8zgTVq1Dyhqmcv9G3FSmFiLuLAYH899iFzJ/Q4ERxSYPKWso18cGLFV
Z6v/4d0eFcP+z5dlrmvFk+BLg0HY4ovpAwXBOFPwfc2EK9M7zrqkeuG78gyV1g16
OKnH8C/PRGGWAdgRvXoRUsQiOgujVes5MzLmnLKf0SsAcIbdr+GyE2y6Y0/mFxdd
GPCH2IboGRekXwcKAMdWzvQ9aAsaBKBo4C1qvpzBJHGYGQTcHE9s1WcmCYHpDjgI
+n7s75nK1xOAlNsZzVbeZuqDgH2ay491vncgUgtAntAVXk4RlTEWBNRJOcn9azdr
vqlLDNnbOeDKtvwHgfuYZRrBV5+MjNrqA3izoakYMKU=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Ds5O8KWRr2uezuHrZKf7IdX5mqcnv6sQimYn7Cua80ZtrK8LTimGidEb/8mhOOGm
97PvwevJQcba9AkWHkvV4tVe+PZrlEWl6FY8Xkso26ve58jVNr97xupK4jcKfyp6
M85a9qe2GWCnNNsy1QL4nb3d4d1hDw44pwgqOUOjHwSDI1mDoDrC7M0WIYefddXm
UBO7DxOMOYy1QcXx/skoxqXNuSpg/uuvFeGDD+vX0cTvsVpP7bnh+3Bbl79o3yy4
OO+wsFYQzomN/n3oSq+ac0Q460NNbcAdfNctMr/jvC1xK8vS+P9F9eWT8lrCJ3nm
akrdsRMTD170+dNIqkBHPQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 12192 )
`pragma protect data_block
YPZaceAjX8MJe3omiow0Noqi0o0ca31kgFNKw3ybh/JbooPq6NQm+KDywe77oelT
cdrOQv4psc15sCwdnzpwpoEiHL7y1Cquli/VoGem0q5TUufQxlqrGW/8PXwUmAiv
5mG4V1D8hrO/Mtsn2h28ImXMDl4WqsYSEtuZsgAhpc2xemztedmQIKkF8N4tz/9f
u7ot9+afF57fxK+IvTqpaRE5CzAwGSU6NXXsI7LfKv99xgCtwWiWktC45pUEuSlE
oGWY21gvTruCs4nIPdkBPHpTrRgMUBPZkkXRGDX4npWPKndhLu4ramyh1jWHZvYo
nDqpP1xsQJ+h1adPOHn9zHfS7ca5BDyW2HemQSF+2w57oXOuwr31UyweltiEUzJo
brUTGiwS3eLoesPPfHqHx86V6p4pkCJh4NfxOly2wklHFl892ZlrBxWR88JVA/ut
XT8yg9IpsqszL5a+7gbFN2biqOZOk+2hlHj0kyoRdkxf+d4GpXv0LeVItJuB9ip3
zaJ9l4PgVhJIDy4P89KZqpo0cyyMSIXAYRNItuy3T8WDtPt0lnBk2APNYxvn6Ou7
sGOJJa/zH7je0UkfSsbmAYPof/7oLRXWHbM488oRhKuibssOPrALTj5PeBgSqiEL
KO3lf8AU+bPH7GNXZdBNFS8M0bhyuccACqWljEPJ7nu2FJ4WoFIPZgrj4iv2R6ZR
C9JqWXfmvRFeqcZsXxI7/yQexuGTVgEbwQfPZVC32E69k8Ed5ymin4XwLiZtd6yA
TA2KXjqVcw7BpnJ3elE2FNRxuoTaKYRHiX6ulVTdEbCJffDY5rPhdVR2ruAUhn/2
vRaNFe0EiDZpVgp5V2+DJB5qW7xGB2y4DEkUC09AjcVLE1sDK2PEUiaXG9uQqYqt
hI1E0KgKbP0u8jGgQoA7MVd4+vktEsAQQSIQJeRXkYMKY5PS/teF1RbkAUT8Q/0W
7PLTf2XteGahyBzWU8W8CvE644++4o2uW6ZMK37gIF80s33Jo/wxZwP0tqXjAJ9m
iWICvLB0LIiPPpMIoCX06BQnQKj8sd7BRR8oGqG2sVR9eE7M/E99YASQN6fegNhS
uNSucM1eVIbmXkCCfRJ9NHFvFAZbWkIMyCYEje6V5u7tr24nSW6w+PrNWSFmm5vN
VUoFv50md/bfX21dsYocyAry8uQ+5ZjO0MIBh7c+AQkxDgE+mM2q1GdbBnOAJm+/
1qpNd8gUqqfjjmfayFrqI2R3HIozyh+dH+Hj3C1DWmck5niG/oi8WhgBI+WuqBP9
Cp9o6wKGfySD8ac04jjdNv3TQtSsNXZhAK0brUzL8Un6wRLb8dCAoDAzbVraqKZH
xaxGzhWA5KIxqzslAISPx5WdYsrtSfA0xC2vd59xxyiBKCa+pTirwfEfNLJvtNqC
4gtrS+VWtdm2eADz0/Fzg3W1/f3TD7m16XY9LwcOCTDJf9d/iLoIwJHshjvWiOzY
PRnarkW1EAszQOBc+oKl4fiimwHuL0gg9KdMrM9XAbAztnRthS2u1HebvsC/RnV3
vtLmC8EhpJXCjUu91jgMMbSEdS84KaZ07wVT2jUtiOr6P1HgGpXUCLapeFd7gJiW
b2ulJ/RAqtRZicGAIR5T9VoEBBrZUISGYmeuDMKFauJqGvBbCGVyDH29I6tlkSwh
Bfz4eHJBnNK2Gr+AqqTyehWk0a13Sz96X/WBSlQ95o6BczLDpEf5jBuQsExl5k51
XcKCQeqOsp8fvlq4FsIPh8ttunNRiVxthLZEt22R5Q2rmzvCTtgxPtk7H6eBncvn
8Hc7DkcyBoxdMEp0EYOPvf58foVlxM2QAQb64LhBou2qHQCC7usWDZhexpEuDTm3
avht+Bh4+W+zGJYmzfPWRkkGba/3Maqh3+1v5YnYwBaIsFgQ8AUG6NNQ2JN1yszX
hqjuRPHSwy7E11C6QTDviUeFiXSjp4TXKkJt3GfCN27GUel0KVUwmTQ0cOVze5BE
0BuoJgJKbb92NSiQsICjsTSf+gIFS3Cbd07x3yS3DcyLfY70cdR7gpeWSyVqJwFs
zD1v6cj6CmhI4d2pIlap0R1LUordpRGgX2jz5RomRSdyV1R8h6B7FHqcnbIMMAAN
NUw4/dlb4XIL7iXpSMYrQrkRBapJuwrdSj+pmzdj6HtcB9aKpjpglkk+fSgd1ZNk
Dp/T/+Ts40/+rGjdTg5/+CEKECOnw5CZZLcm67djXK4JdPjSTp4q1toE93W+kwg2
WMxbiFbrpFwvfgris/Wu5bvOFJGCal4lCf17h9MF4HtQiZWfgjoWZVKfdBdXnlVf
a+iFbY4EBBlVClnrmUZyMEyA01qy/YGcYyK5VFIfDFLPilPXDa89D0RZVhVljePT
8UGRH+r9S3SurdvfsVtuNC7tw9xsYId2sXClew9A+8mJYmJWRcpY6A7xXpN7Lp/J
WqfRakAVLE/wOWP3DriU0jqNQnyeDTqWcuh71quK95eiKdIzRAmKp1qbdzvR4pC1
S4TkkL7Wmejgb3uJM46CseRPR8MgUeGucOT2/4RwBBvAdCkGhYs4beHtk0wUkdHS
MSwU3TEQXL+idoFikufNlBHQeVilU4odMTASnslYtLu/M85XCzAiEweVaxpz5ux2
V90fOFiwFUPy6Jq2Vc/4cHQD2y9Q/NPISBUoL3Cw6p59oWdcQgl71ACnOWwqQGa/
ax/bXYTv3HJEkCN/fGFLO3lKCsobCBGr5osp53i5vSBUQ10CZvDnD6fAWeZSls3S
9jST7R1SJG/ctKr1JNWgq6wU0gW3wv7TGACfK1pyr8P9GWN6z2LVdXDUH7tYChaS
Lb53xh/fucXlSlmmrx9OPJZlLvZnNwSBsfVXrZ/xnParZJ14PorJAwRaLuPkTUvy
fQEF/U7U/A6XvYtlO9l9uPpSTG9Ouf4JQ6CT99tWHJyxJVJBp9TFugUyFJuzsFvb
jFYsXAOnx7RsUbzVbw9KIXPFmycM7Rnf4rytg69Y5wXvCHuIiKy/YTHndz7q3dSQ
xRLPc8nDKHmejt3vAfz9HmHlgE0mHiAq/Ntc9HS+WPgiwlTJyrpxhQoz4+0PF35M
XVMmnBe7QX8g/61GW5JERASLDaS8Q0RP4nKHFhtB8Rx8p2vbUhHoOhk1Zj5BU9Cx
fcg80hD99ff25uIRt9j1AvLU9TLv6LYUgGoc60s1txt2xM4szdskPZrP34hIp8Uc
+IK+VYdlAbVSks/BwAtDvd5742RN+C0JzAcIPqYZIkJg3B5S2SRp+YvLhs5UMQ6j
TU+lun5OmXNa0CfhDUR7c0LSiGlViSAYfeeuHfLXpYUC4++7jnDTd1VRAPElUmCU
eZ4xtz8WRBjLhos4fXywiy1LEpj9DI/qanDJHyyiLFmrKwXSd7gJmQ0RU4qkvotN
rol8P0NjQfOLwPlO16XTj+YOxqkXh25mePFYP9BVybXixxcjS4WFr/O6wr3H8W04
nLKpv3WeESFcuVMHORGfdVnd5l4Ki6fvCL06esl1EOrs/AnXJlacNzyOZ1wp1QR7
4gegMZ0zaOUmk7SBKgL4Tatc1OSgurLG9D7N6Zdr128VNS1m9UfUOD8CwvkS+NSo
d/M6/1l3H9SZn1zxo5LIZusrkvsctVoPz3fV41RiArb68iT/G+YsoDBjHjhBJxq/
q+NDb1ymYs8pOvpXzQgSy8ZOmK+DNZMh6/arWqImdovnKuMGGmOBXElTgHZ2TAVA
4EYHUxgRHuop9YEQMqh9ySME+KVgRFyn314+qg67nW8BNuDubKkxGB+ZhljcS1ik
mfyIs2biTbDzljTAHK5lgs7YI19W9UfYT4/DscxJ9xA1yUh7wSMRmeusCh5KYaFE
+Ruul7UwS4FN1MvJuOK0tp0rvJ2AOwF5XHnI7plZD12/2r3b01JLbASTW37sc47m
SVJUwlcI8ICLq5zAWpu6MJYmmu+n2N5LE2B6v9Nz8AMaVytLiduhCVgo7wChTe50
L1LGTkkgIUsz6JYlCpymtmgqQsnvKR7lA8ETsP7FnfBtFieW4HzhXWDumON3jV/2
SzTSEYAx+fmYscpu9f7nbV2xscHFu4bp/0fHOoYxLOBWlCBlrbW0cnSS35v7IPkg
62hTcIRVoYtGRHqBmSULZNrvBlrle+pLzyj+uNDBpJ0peRsz+hvE12aZHrnwvzBZ
SqHHpG7LTTjuSeCATm3tY9j+uEQSNji2jU0P2ycPDrhHhI12MAAibddHoCK5kR86
1TfmoT4Ls3EiHw4bJyYV2h0FAURuFkTZmFqRVW+g6GeQKcCGaNIFmYovlE2sxE2z
5d27OYBP+KODeUpTE2Z374NaY3s1reYhTXPmV4+1X89RtYzo3FiYYbe0H9JhrSI5
VFQiWWYHokhqaSph+TwHDd7RkBvrVHxYWyn1bcHekOsBp1iSNmm5aaNbnBQoEAqW
7OpeIvSgJzsloGKUh41puisALVryzJ6DC9kDeaETtP+YZXODDwKCNB4jOGN5Axz8
EBRClS0KEJ+wa4p/O2fwQFs5o1FWpTGb8tsgxZefvXrMMI3NUgujQBnpkr8EHZ2e
xGdqTdKhlnTlx90HZ6OtVC5ctmfGOSCyG8y4gVGROFnLFC8LnRQZaWCMzKeWf0mN
IW37WLyAI/ww2oPQI6Xc+Hx8nM6dU1glE3V4h7kumEDFabWcVoANluhdzjVwmgHC
sF4xC4+ljS6AStDG+OIkETNqOGdlNa07ZX6IU3WYpCnmadc7kqzbExa7xBdhXgH0
VXb9qdXLVG3ZeOKP179boDxeg619RRgMEPHge35OXzGwwrQErjNX6yEkHt5gq3HY
MX6yvDcjzwbsW41YO1cqU0rvYSblEyXj0QAXBoju4K9KEkBoOaG6XXfr1Er6E6C4
jiqDld9Q1cMnnvT6TWhitAwcvIey0DgtebyG9F4/9JqpULxWnuX+kn9uzikwBxq6
wz7AK+dxs8vuNMGhqFevqHG8LmzhWG1HRT1gYAAKlOGe1eCxg2pDjr+oJXz7Tixy
sPwV+uWr3fVb3YN21HcLLTvtWxb62Ch6fDK7KdrUzVZK9g3tShg0uolEZ0Wr1z6/
d4MMiLaufX2Zlog1ZjwbTR7qKWmYQvjF4mquEgY6JlRAxYagUBRTbfNp6cNMOkdW
+CKnO1qaOrHbHBIEJ/gNSQ8SF/CoMDrPZXr9yphnIduza6gkDZQVvhsKRMKXzsX+
kbXHBisLGVTTxI/9FsxBnMZA9DWzmhjMyyY8v4AReveJv0x6+tCoVGL+Pidc97N7
gD1oCsLTe2jzJX1wq5ba3kFBxVzlqmZ6mXZSUUg4anvTncZhS0qYbQqwrODs3R9p
CT7llekkNfDeDv0wvPTWP4rWdobnY1hqVbpUP6329yF7eTUU4BQVHdTUXoRYs4Q4
WTEeY75aZ19KOt1OhidoI+os/H1MehZhh0m3Jz6aUuqq2UR76+1lzZZsFxY35Yl4
BZRdn/lKGQo5r/9WASGfoTGZgPbGwn0vuYmUDHSGTJ3gAkQswff6mHJtYhGWWBFE
2MNq61qqlziYEnJmHa8yZuJTc4kiUrZV8q5MxUxeyi3a/9yl89hx/EKHstn9VsSL
3ZbuKTwEypK6PX3ff2me/OhCDiKpTA/hUox+6i+2Jah2pBR9t0UqtR8RPx95mEde
eJCgUmPF3YGF2mM+jji9oiaDWuD2wud4nyCgutttEOJV+sFnII6gLMxh9MuugOXn
nw52ZL2XHMLGH2ekr4vxvjVUyM7MCsbGtcv6jjLAOQ/MgcVpnlkHbda4KHcIjIwo
/s0V0zehEO0LJOWqorGWhFL/Qw4EHBuglR/OSWCkQ+3LBDSZhvLrRPFviWMpjXz/
yGzT19MylECML6HuM+WC0Q3uw740V7W4PyjY/xAKgjgz1PAa6BwGUKJMdyfO8Af1
WDBzRTgNFeilusJesOBMDfpiImvsnRJQvcfbQcXLV5ZPv/0BfnnkurD3v3TU7DEo
IcBheLC2nBHNLY3Yf9qZyRuhzc/a1drh91UDhW9Q+TykbeVFMcNDxe5Y+sbEBS1C
W/hoDpeeaUAaOtwXtLsmxfuhb+lnkh8Oq273XLInLc235bQ/p4oMqVRSgN91AOMp
kXmBWDFjxXf1st+ij9GJuT3KBR54+XSnb+0Os+yacBsu4ievLJnrrupg9CTWtd1j
4eAqcsinYeYH3YntM1MR3+OskU/pyYZYp38NzXIWY1UUB4pBxWFy52U+YO5Dobaq
0sBB7Glpyi4AOf6vY540Atq3BCIr2AWt4RayNU01Bp0twQOOIGtNH0hANPDxojzu
7nowMUdpkd71O1k/J8PYF4kcU9m9b7jb+JnoB+srDEKwzcDAUa93UFCCL8DKy6vL
L5CVd7jPs9TmKEdh0yqB8ebtZNj1WkEomTIruKOfyF7ay5Z9qvh68LQd0eGFfjPR
ybBLo90yWvbOpgnBfUPe5UEy3z9aygAjK0/Ylw/MbHwoijYy6dDat9Ydn5Ilg0zC
/AJNUr8sqBFQSP0SyAptBtMQsNv/4gEmZZkzHkfEyUHH0tWEG3Ne97HnBatLrru7
AET8SdWxoGWVLFAlVbKuD2kOXOCw1jnevNhdzZLVftkUD9Ychdei0jpqYQLCwBrz
jMen1ukuGQNwrDADJi7ETQNHaxBZL5Q/iuDHlx8X220aHz22qQRrKVXH6gZNMNPn
2As30NDjvDgG3Jp0McyL7RUtY6ZGGvS2qzBPTEVMfLkJiHOZf2CUykwjtciVVEDj
IRga5Q3shrshd1ngfJqj88Q3vXyK4ItgyzSS+J4QVK2/4Zwxm4vzUWIZjAyYljxQ
+yqGV7PPrHvoJe9BTx90veB1rocNr0ONaezgnJSLHwNEiwIvE3I6byuqVyxz+jGA
dFzvnp3UYjetmtpxq9kVDrFnRN6+whYy8qIkFkhYx55YON+MEQZpTahRBL51rzGt
PnWnzSlXqNungd9CSfOaWZpHF4Mbe6i3LGSz65JoRHF6+pqsGRwBQBgxpQF8arjK
z8NSRZZ0lfG4frop9KU42640mwk6MBTX9jz1WroPEIhPGdYcjs7r700UIlSxFk4O
BxAUaFwvh4lA2MDs58Cxu77jVQypyITjD8C3xFqhwrNc5pi2WoK5P2x7cUcWJDkQ
ejrwkoe1rdGeORgYZX59KuNOVvtNh3r3VlHJnIjldRnvTz40GbUK90gLhQwac7EK
FZkwOgPKRHZMTmltFR7PfRaH90eSEANjqKrjSTFQCrJR78IWW19N7+stOq2W1Ggu
L0fVyX1U+3Hh3UJ21uoInItPZ0U6XQ2Jp2PMP9boif8gIrGPALJt0yX2awDigIYL
oGCPkQlco+6pGhsGOS2QXTdJGTG1pVhiMT7NXSmwF4Jtd2ZVTi1Uq92IapH1LQTb
iWY8mKH2j0tlDegss3Vq9fv7Xdq8NgPpPq5SZPH0JYh/oX4ENynqbZSWyU6JvyGM
OZtZv2EPpMd83Gl+nUumcw1G93vPZhhVTem+dFsn3HcynDqHm866gX1VH8MFYiXR
2ee/bKL2w5TdEy1fiuQ7ymFu+4rQt0CRcI/xPKDvhJVj8EpuFBBaXq2qYCUKMLPB
02bV7Eqs8BBW+GMRPGhasTd0mO0OpufBjYFjz0s8HHo5E0hyHuQu3zaoiOdiMf1Y
HSCW2ua55KHjFGyqc8ZlcZTgSsbxX3skCksu6NC8EAXElgTtBdJ4IYsAtJudFp8V
30Ezks7DkOuN1yF6h9OR37IAaI8PYASepjQgXBt9LLLwW6CtJAsOBwYbtt96+NXH
v8QA6LsDApHouG2LLYTrQMZa+P/Ju1YwlUFt5xsaAZyZ7p8+qBVz45YuqlVf2VHQ
zi5nz8ZuGA+rGOi0fzZbJvgZOfE1pJhYCbt7VaSvksecbS4GrLUMp8WdOhQkrVxK
vGzmobbkqIHFEkfoKZ43Wkk8i8sFswLVlfHTkTyOEUlN7dKqkzUQA9In2GLN+FW1
ZCu/0SUEgNtH1KZPDnG5yhTeXOHUoLVxzxjwU22DWicUhxTIaLPa0l1UM/oEQo9T
kWwzq3Zz4taZntwPFlWTXRirKIju6NTXvhjbvSZZN1TZbDJ90vYiRKS4R9EhM+rj
Zq3MzljiB11K86e/vzQVZMf4XrjUePNjFZ90PDUcm3ExOqkwfl6MpKzi0vBrgL8Q
wpCIcYjtl6WBGjp9vv2BKhtK6Zb+hwONT+c5Z0NiJNvJwc9EUf1oEw4GdDXWqG2K
ue4f/dchhfsl5b751sXSe7abGo4G7tfLBkbfXTe5AV7hTLAGbwOxcJgTD8nX5+lM
yKfdHLoyMteprkMP4D25gge1EisZM283FgYTFFz4W+EFZIBz+pq9P9VThp0VDElO
P3Be0xTspsleQuXivesKSnFg2eXawRMSV3ZzDiv6XKOVyF48/spfBG+APdYZPxkC
NuHB88q6K/JHPcw9UlOVdqdcClEqkHrMzCU5rjQs4eL3szJhIpoVikr0oHchGJ7Z
GpjZMwllhftqsliYWFy+DUpHkmsdh35ssCmZleDrNBzJmsIGWRZKC/3E1q1arMU6
Bfj1Jtg8s2bN7aS9eqxnTUbJYNAHmLOOw0ZlaaP528CX3HRJP33wPmAcm1JgiKDl
gfJ/oaLkbx0+8aPHDp0qP2eGQgOmQNyEbHUUr5RfSB5kawyLrsI5fnbribAdtK1x
2RBUDrqfHLJkohH1ntT3pc7enMh0AEeusPuMcm2RFihEA6HzV8YUR463+9czn0jl
xoOzvV50l6bFuQpgEvuZ39+UfRjPzVTrQ29dMox+yKBZdP+KlOP+CBW+xzuDXGzw
QMbrEy2JQ3o6WeseJSIXvUg6jOyCGS3YiapXx/bzBjgWMY3m5Oyd+RknvEWUqnDk
RDYS8iMEsQDrHZkvx2dxiEKxg7y/l0/vaovVIulKUk3hyOS/k9rMyn5QRgzqReTX
DwLpi8og2wf/pxfr6zMlSGOHg46ZruT4/HYYSYpD/Lja97Ll+ovNzPcMxAydFANb
IV36Mgjh2+qdxdHaGJHvswJ1zl5fLM41EeRlpBDXoDKxigrwf26Iu7c+VwkFKCx0
xI5pG9aECcSznGd1WLB+fiZqvmC5bOlFolXhLnUZokAsG+Kht7y9NhZG65exEgR/
sjKophrsqHZVLX8KrGE2Sa4skxZqC0DbG099xWDeV/BqwgZKVYx52OvnoRH+lKxo
OexNsoGFI6jLe+0id8XSymyaOyYSgEao595uOZYQTTmRtw4bpHpFFljn4HGUlMaU
J9RIU0avuKeCMEBEVOnsdd7eSnSF6yaWQvsJpCTxqEycrDLZipfcr+OSk8xwyfgh
9u5EfD2cXqWNazY02PSh2xJeZDkvXYGnn13/bhxedGx/IHJImX9QjEkn5BsleW6a
J6NeRFTbcnLso99ea977EHY0G7124BtymJzYd+tfMk2Cg3UojexSuQaGAHQ3tora
h5vKLwVl6gpPszabfRVve8z+8wkxrCkAyUF2BbamCwcfsgmk9/iLQBrdGy+632N6
QgGiCYzr+xI2s3u5g02LyP+W0Gkf99oexidreCkLKQObttGiCYD/tbnpm0uhkng0
fHv5VR0LvFyJl3cVevqrqittChyDLHevssAm1jvkL/j8Xn7aOy9ihDTYPwaU9N2D
5PHW8uSZSx6r1ayr4BX+wtHYV7A9B17YGNWbzOv/NaTaqWm2zpZ+Z4J3cszQz4X+
QyeVZVkqz5TR8UH51EdLPnLR7XphgSI9dL4bKBi3eHOzykH3JJ7UaaYmJAXPtF+0
Q0NCZ9PNOXBtyDJDUh2C9S4aSIj1LBqc1bNuvW1UB7W1220jM8fnyS5ApBqAy4kD
QeT/U5IlWubQ699ZYaSLEKgmzJATRhmqgVLZl+4FG1Y7dVopa050F0e5y0vKxoPb
ZrMP3vSBsVYE1FvHXvmp67Z4muRi1wRgBoXIlriK9lPpKCjGdd3o/qBHwfp4Tx9z
VnIlbg08xJZQs+H98B0KtsAVMHoaxNPRFF1yOFc0feYraFjBK0XyaBp3D9bFT6sD
19KL5NVZ17rFY5SyBBRtCOhWWpDQOgEN4QCXEb47ypGoC3MjA9RVuWNCIZs1cuuT
JcpuLIhSTIp1/hzH4VIQkeAkWYmyOtH/ATTE8Mnxe7NLhFvxwHrM18CBraEiXXDQ
KuH/s0ryIlyLo3vAqHKgdCSPQrJW5Vvnkpr40AyC8cOctpEhTnCBmBi0GF5x8G4P
Fbk0xjTvACTaGB42GH5v0z9iDwezo2Tl6Vvgf0J7ZN2rKv8j87qesxPY63030QeU
H3AxsV94SBncbE/A0BAiUoVHVXbHepwIx0qwgQOYNWrVU+H9hoF1UtE6Xo6MhUKn
DTxqMiB9jfmraECQsLYS44AuqoB73z8cyIc5LJK/tk8rT+366yMxdsiSOwsht2pt
v38lx+J2tv9k6sjC6V0qCk0pNpqvmTqw2A0y2wwtAJnRJ6GYNulyg9TF58SbmxvN
wUzNbN1Xk6aF8+Rsmo++QFLt3pOpKjQ+eS++GZ5P59Zl1PkuXpv9C7OqcE+sjgbj
/g5MkpxVvntXIjkhC0V5vsF8FEM5ETBNfnDVWNqknpI9y4r7m8W1waxPf0CtD5v7
/m/lZrFK03LzUdURd4hcVz7X1mUTC/3KxGEtz83boVV6WfMU+yalJHO1PjMPQU7O
yvkvInnip4nJrMdan+RNSqdxfa5Lk+t91L5y7JnjS4gLbnip5Bz72150f54WloOk
XZeqM93MBJq8wbHaMrLhhZAUjQ9SXZ+H0XSU8iXAiaZzhzwABF6F+1yhwuS0BELH
b/DqyGXs+QH5dww0rIXHn3V92NzMionpAxbNrTC2vHb2DsbLnCyaproa8XO76Rnm
nSfcpiqMjGtrxrb4DuiJsh2Fc6O2vDWRSA1LZjaEIUArtbl1+1mtkR+9YI/QGopT
p42yEfov5cUmtU8x3H3Uu4eOE97vh9fsQXupsGmjKVn7Mul6sDXa1N1/kb/liQm3
Xyd7Zig/kxyu89Ezwh5E9spTYBb3jQfa7jtaB8TOQfMfKUVRoD3prlQSxqkr8Jtv
kjcQ0rOwEvZCMqqDVdO/J1Q4rASFSMRkWJ26P9S1xDlx+UNyPcW4KKehD4pMAlai
Mw1EN/8tzHyC5lVszr+7P5xscdt9wgmEtdi7f1vIJW9em8mf98zWLGSYCUitNRA4
jBT9iHPZOsamGmaLgjzsd5O+oNGrekPvrjuo+v7r/p+GkAK5hB9RB7IeA+X8faAV
UsdWFSHGsJtP62iLnBUjtOMQThUXpWIml7FUg3DewuzRRjgR1RzhubOIESq2RETl
BXtJYnR5thigIlDxunqEOUPB+eAUDQI3sdjZwDgY0y29AJ+xb4/gbYJ/Xyks5G/T
jjsB4LOmdDNxjY3LZhDWn1x++Xu3JFoSWQTFuHbKLB8RzKoA1k6PRpuugEE3j97D
h3U/KfkdqwZ/2kwfNTuFmpZQ3/9WBBSHMwwjmYqwh7eTKBn/HI4yYzeseMm9FZQM
QC//OB9+47VCge0TWsJF5b4XtkUNTe7NbHrcNagpsE/gdUOnveIhPgHCd3ggriMH
d9syrpjNhg8Ssu4SygajgFviaN5SkhxoPcqKsKov/s/ujFtBLhz07padrMf0RhJM
MAMWczu1LHXapOhsSfzirzlErB2ti7abqXI5wkZ2bW2dqC9IAVAI4Z9Mhuqgv0dO
k+1K1oG8+jGdGQYq9tXh2MtV2eFiqM4WDq8D0fl5XvUfkuxtLa8HjbmOlSMQe2jB
mxA1vp/rfP0KbtYCVKukGrTBPy3xDs1W7M8FlpG1hJcalQZXSxKeKA3ocICWvpDD
DfyuCN7+TQH1ZXf0h0JgeMjlcTVJ9zNkbizt/aCgPcsm4P4keWnUDKNDQZCI946G
XVNFTUjHy251xryAE5Ee/z6aBLNJrpfDSs7pcSSD4V4t/CTOhfg64yv5vF+9DYJt
YVMZ7hAf8ll6j/gwbUXmNm1fKf5a3gy6Vin8l1Lb9zFvRdvAUzhmxOOBS/2GFJaN
DTbU8gTdbQgD5F5E1ZoRDCAO9zmeqczrpaaK6TCyWMk5iRZ+kXuCKaWn+95i+3MC
vAu7JHN9zfJuho7+Ng2S/1TaSRV6LE2pqw8+MX7o0p747+SD8/aBXDJejQeAAx/y
GKAj7Q0xVPCf3N8BeUBOzoEFVOoIBbNPoMM/DqU8WlfE1CQU1F9oGkvWMD3GmELt
spnhJK1WCDHHd2E8OMePpaY+kfWf21uf/yI0whNKSveK9dojaYn5eMnp2zXuclFk
p97gHa7q2tnm6KAykxIPQIPeIq3KCrVMzsNEHFhTMXZenY6wATGS+6M/xa3cH5i3
M1PB3dyGnCC3bFF8s/0FkFDBln5ZaeIvZW6vfUrqyYXm/tXYV4trf7aHrEm/sztq
hDqBChUNt8pAcJk6TrF6ZyWKOG+ZGgTtHWILjvpKb0MdHYLnsHXYD+l/pCH/hv5T
cg6GNrQSHRU7wC9G4ooW9lYzlRlw6MDQ3QOo2cfq1plgADmHvsaAF29XCUGdut/i
as7RDhwC2L3es4oQyzJQXTCsU4PTRWc1vKFA/2hS0FPdQobUKqxvCpyPUcl/FG4Y
6HnBXwRltjOnG7ifs6gOeyp6vwi2eojYJss/bmVu1HJEHJcv7ifog9/R5L7TdXqi
sZlf5SS9RKL3fSLBwHICML0Z4neXvVT6mgD0Yo/AXovI9KcCK/h3Kyr3ed1pbl7s
XlvVv8uEWgNFV+S0f8NHKnGkktWL48/FPtFzmuHUSddPMNoNFMKp68ojFcquaC4+
Z9EKfteJXXeym1rm0FYxEiGMNB+rA2ZEEAqhmdpc+a2RrNDYiwZSD48wMgz8ZIgY
d4LD5C/6fX8KF5BvCTtDF09dA/+8UIB/Hp+4EvHs9iZ15PGlhy56dy6rkuftK5LS
WdPm12EPBYqZGPqsoZHiig7w5hCEh3UYmCO9ajvOr5bdTyphHPlhhTeaNcQquSFZ
KBCAIvtisTTg70C1Gp4krbCLwI0yCC+CjccYNVE5VLgLJ0Yvx6gluPvbVKwLlJ+8
9yMidon2/HEXMnlqUh9iMLw9A3FNqfMhPQHzK4OcMlO8NXJDLQR3CQN7JgOHyezK
4PbiYAZPCB+CQ/wC7+MlMpSAzHBoBqyqDUVtt9AzSrCyvmrUHdqYgQ23VThgNotl
FITWYo3+tN+mOcw/q0b6W8lM+VQHTe25fiHFWdbLM2z4ndzPvqiUACZGj6hW0yE7
WxURTjBjLQL+M8MnC28h21GxIzUbto594jgWOQMna38W/A22zvhPZhnC0okX+cYO
uPqWecjL5ftiDh9xxi6CHntWli8UBORrIwV0SJWQ6AdiI2ZunDzzUAGUNBkcFh4R
jAhdqzBAhmaEq0UHsP6MQ6Zh+sAxE881laimxtSNJdDlUvuDDoE1TlZutnwSU/rK
jpS6NRkfbWmpPqNDW9WHA2MR0CnnuT1lmelhiDPnf922qQRw2nl/CAzOBbopA3kh
fXjriKUfTjL/Lgt/UrXbSg7oYSoOjPeRI023FMFhnmAdrm386Z4D6PqSM1Iy1vPF
pH4AmBWrz5g1s5vS974yGLN+UnGtyOpQRJLpOfVUBTvdcGnLdZ48HUcPQRje9Ih0
2LnHYfvtKDCWwT8foUnXCWvdzLqBbJRw5o5dVIh0CQed5KQFTvXuX04UUyfRAhQ/
YiWPlVr/AGnOsqVALrDaE+2DWfkzYAoh1wQ0IK02dGCjsq+LhZZ0jk3KuLjlWeA3
QwPSImKfEO8wJnKu+ZyG/rN9TtusmnUKm1McdWhXGddOrbeBiIAOIoITiQlTdHPU
fFa12gFa5Uhp2WTYb5Q7e2GfQTo/Ush6Bjuz0YKeMoD714knQyunwkxSNPW0gwwy
1kB0UDeEChiJDNhehW5OHSg3xsG13Gap+KNpHIKKkCB2VQa1jK+ySAcUnDKsLLh0
rteTZNZc/Y0F4RY6/ZKFr/+CLS0x0Q4GR14+uDdFwjBaLeKl8VVYSDXQDBKbju24
FdcMPsaoZKeELmhZrgZ61xFuf4RH9URtsqibiFq68WY64e91p/f3WFNfritp6vEZ
+jjDMeEMXgHMnUaj5AcTG98YhqN8TsKTY2f9Qgc3IgkqfuG4uIae2yUEA+V0G8br
qOaTrb+r9sI9gfyHfHVRaTFvtS/je1h1xPhJtGCTgFewwDYxKxWwb4R8Mwfpm07u
sKu51MyTvaTdFVmp+tutl09f/k7lcu+N+Z3/nXzwA5MPLBpVrbJFyE4BKngG+eXv
AP15P74S9WalWfDWpbGo+UMdp8204w13LYO44VcsbNz4k/TksvCbBje7mB3ZdOwn
/blA+Twuf/+ddEg7N7JfDTkKtGd4FqXHQBlew0vNCNHKkOohq160QQyvfAmG8V3Q
WRiI9AO02yDE/0K+DMj9DARS8F5wXucnzbg8yku63h+WQil0R4sHgEQhKqV5OGdK
rqGoAWyQRp19JMujsC3vBQ8WXDJTQejTVj1pYwtsng2ip47lJBpkdXJSzOHYtBSd
9clEDjo5pV2euGYCCsOr1dDbBHxDR18W7uD9cy9bmNuGyE7DgPX6zGgmMsiHbA1a
U647yqXS5yJVyD1UAH4FllgxPKGMFgUgrQwjoR2BzDR7poo/qaLnEmXDeo8FUvtm
vJZ0TSZkqLB/nxssC+rhWbmmZKmdTfAbTswcVPnsreBhGAVvqdCsF3/X0ZrbZIl5
XVasbfUjnLaP19aoD60DEEaJW5SuQjo3H/1/Q9z/4gOhSsdSJr1gCa1m8bNErY9B
7GHQmy96IbV/YtO0NOuIX3RuJ/n65lQzpAQIOc31CP0BMahdIfc0y/GiTNzrMfx6
PGaqi07u+L0hZDnwjIlFU4uC1CxOaM/96EU/Zzy4ZDmsl3JsVxkiohghSHGkbVdW
YClABKmZMwtZEZPFOotDbg+b3mYRixrQMNuLa5XeveAIvPO5wlxKAARZHpKYYSwC
/Rdd4UnK5JAEZuk5BzNkxw9JydW2tn9DyB7zWfdzO25qGaZsrqHnyToHGIO3Th3S
l8ZE9PmbTP6yqNh1fpem8FRORisndivEFl/JE7RifPtH1V7jB/shDpguJ5FH9Q5t
2Eu3gUsao9cfdlSGIPi7GUH6OYg3YDhKjlhNXnyeFJFZ36DUMZTN8jCXTGSd/LEy
yxT2m1I8ARwX98g1K1Oaz5NIFMa2D5RSrBHDcKwb21mrv0ulqFTJCQ8ZYJU2xDJ2
Uy53757kFUkPjisWRi8au+F55ufxFhXr0Yri4TPVxgr3kc2o65g5NV6a/rBNKWlp
6RsvXx9R7gLikKopO6GG/3t+d4nW9w/unFiqqbGXaZbqpCA20dnlahmTakxR3O3E
NIc2CnwtrsO0NqFAWnYG3/gbiAV5sczKvWc+nyOAKCRPFU3MUt3z9D4ujtjFucqn
kTplHoKwbHvTNWBVSJ+e+0Yt9UQTF/ljnYwWL4pnq/NwJxZD3w6y9aCV7OjoaIy0
b/iFx7dPxQB6kLmSrc/H9jjD7Tpi1YLA0WWuKsHfkXNDWRKJUKdF1kUozyKLht7X
LehYLzbTox5snZuMoJgY8FU4IQmJDbEIvpbPiWrCaXHOFiptPZiFja3AB+w9F49u
ni6LjuvJpanyEuzhyBwrjyQOuY4g+k7/mNaZnlVN1hzc2yvFLMoUqw3YZDKPARBe
5nNDarTKb7GnzCEEchlf3cPk2IHTwUij6zoW1tSJIb3EMRfB1ppZoNvXoBOUaDmW
krbeFHxJz4iPkFxWw64V/EfP2tLMKXhvg8Ts69W+ESvWsQcGstMW3ZfxeHcIWFNc
VgipBOx+UYx3Nvdat1bCD8PEpUoJoJfbiWfEpaQLNc0DMgzhDYdL3g4SbMuTSh4I
zsyfAxkI5weB7FC4q9K0efCmgNYdQMSuspDqbZBmKbyJIiZfwNODZaBbYiessjuX
yoICW5bjB+mCjnZMFnnbHuPuyaV8fMaUVRRhXxX1Q6P36ql9zIwXgnK//SrnOk9k
uF9bwHpyrYT6TrP9ZIkfCdjSidINM3AzeOecqfJcWuTaDguSBjaJrxbKBpsORTtj
AI9/QRjKcjLbb4WErhVb9F2EQwQMl699MFeQYAL+RwWAEjqvCuEdg4thmNiD2Kz6
3F6BNZe5F6yryVhkH9Sr51GyNR5vlkmL9EiEfxuUex5pCBf0b9fPP/3liJiHfw31
4ojUNMksenDEeYdK0WhsMoA4iYgeROQUDVZUYus1qPBGvCMB/O6XNXpgTwD7zWML
NYio4RVkAWHWGLz9Ss9SxS6ihdwy9Gg36JgB3mMGHuO1h+WszHr+a/4fK4OgbZHa
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JjE9MI4vsYUWwSSBfbuM2cP+7eaMq5BAIkNRAfty5Wab2HZzLw7M3vUHP6CEKH7K
2c/4BfqCPIU+H76dnujZg2ZkVTGQn9pfDjWnEYjr3uS7WjTNCiQ2V+pmxWO/0H+h
66W4FnnJVMXXG75exWMqFVzAizjc/RQvLb4N7dZpNW4EjzkwHyTrZ8c5zSBqv6A4
vmppOXshS9N1+mgB+W+6TcK/CzsP8qGrf9PMsRb8tMdX9x++xLCKsEGnJQtmQF6z
U7ZKuLjQjIbDG50wQ5visAnpMA8jrfi1yydyGiFN+yEJ7NYfA6dgVTelyxdFi7+u
2tjvgi9OxMljjddy5b5q2Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2720 )
`pragma protect data_block
OyOCvJs5evRaiAi6WVZrTLy8jKttGiUYEuq2Z8yM4CGK0UmvrOb0GdcR28Y3x/pp
T8bVwPxu+Veh/n9+ieVJo9e+9XG0D+Q39L3iQRWAhRRzox9egTSNWgQVX+WH3iCd
1W8DEe8xjZQG7f+ZI/z7E8CNWdihfBgSi7ixNkYvFyzIB00PDk2F4KFGNjiPlkSq
yqoJWq/nAuCpIkhJNQLZ7PcNGygW9dEkUKfh80B9mztRay1XHhJ4p657T6dhSVMC
7YVqTZpdebZSMTjRe9BOBEURJKFApGrX9df/XljTVQv6nrHF2Awea23zDeu8Hond
M2lBZYZzzg1mYohBShb9unR7d5oPBj2x1v+8hhZrbZIeYO6U5n5wfMFW9kstIvGi
IWbpa+0DkJu2uFdc6/KniVkErQ3e8CpGp6IMiKLK8Dw23/foo+ZlYiyq/L1N2j3T
RkG6qId50ccap3wIklD0xYDdUTZMmyE8/xfajktgC57bQIpiIyI08/3OYtk6vY6h
KqUXWWtPl0FbBxIN03Dd2ZA6bfU/KtRsBiJ/khlz2llBBFqcjOn0TMOZMYAxKeS3
vf5qB9ss9V2+vBy7P7+MizY81Kz7JQmNUuLYIrrGq3x54Fo8/YVKgosONa+JPg+B
qkUkRiaD87F0Tl2HMzSOLPsjLzpEWWtDQx+kb7CZhzLh556mFPB7IzimXiPJnaOn
eP7aavfjKs/gBF6VveWw1F7/Dzgr6r6BCeti3wNlCQ5zKStRdBwnxAoh5MoT5pJp
x6VXY9fmerepL/VgWXXihEHE1i4L56OKMwMGPexQgjM+cvVJ1qfA5wahUjmCL/KL
PIBTKCp7A1V3zBGETH8X5SVFNMSWYJD+cfqiB7D6fHe3jjFoH6P5dYTD8/CmoAsq
RPaNnnGk8F0/RRgE8VO8gB9Gcj0Npqv7lfPyTpehygu1dRGFa2a3luojFq+88+vB
dPpV49GJlxgLFTSWJL4l2pAqIbJY+hG9ZcFv+BpmTRJ2NdEOokNx+Cc3Lo514Isq
aNSaa6tzqrcfrlHmedG/iIhhS4lJeunRnjwhLT+CQd6QEn5LW+I5p0xLMjyrQj73
pfQ10caDbErIcK/JG0wEB33/BQ6/ot+3xeEsKKNCVrj/R3qGTxxqTOFbMZ1EPXEa
u/bfeiFtMtbfLes5t7fSYHPJLiY9Cs5PBBQnx+0p/4fOG4qIDNx/2TsG09gvZU+p
gIzS7o9DZUd2KDZw5k1T1GPmsbZPWjVpN2FgB96NfwioOepzQqRHboW20p+KLPha
MXEwMwJVLP49dHV8ibjC8sY66Qh+1OlCHpYxc64gVrlCugmcN1leaf3C8CnjacPq
4l6X69eBhr7xlPRjr0sXR5LqLVJx3IsbWZ/BRTKQZq1Ndv3bdyysJACtLHBQsw/o
81PlnFrTDJkfhhZA36JZ6i3nB65hgxm9WVa3ej3f1YJP4aNjWSCvnhpbEVoYC444
DwKg0D8QfhHcc1DbnIkok/qBOINg1nJF/q60hvXkYyaJeTxp27S06Agt4RtJQ4lz
Cbdyee+56+Dfa2gtFLzZtlrwQgBK8BuWMgQVTihtHHPXFJtbrQ/JcB0ESc/G5sTo
u9eoBppUMHCC58s2a9rHvXZwtoZhHCsj0cIWAJOXq7ZE6mw+8ojpFMGLPn3dHEY5
Yte7sylEATJbiI2UoyQYBdOZYb97iLxqgZ9onu7oAI4tAmkZIAa8Q/3R6JNv3RXy
O5ikOvTMEq573oLWpxQdpogAcSJkmIsy0Avixwm237uAGLoo3v5oTfHViviuqepH
Knbw2jxeLsxxoPw3GsS9h89SNUNB8EUA1OMiNIVaohpS3oGe2cZCoPgXdOvQ7weh
WgQLLgnLnfqz/5GDd6b99l2o8wYsQUbV0jmyQqdVIcpHlG/urSCPpMpPh0uVgRyl
0TV83aMwwM1HHT4Qxr+UVJNJzwoKgZDz0aCIY0SLYnQncPMhLkbA9XSuF44s6Hz/
pZsSfnh5aFqP5/HrSOUkUxBvJ3ppFMk/mhCBQ+Sc44ryKaP9M66lgBTM+r0Z21Uz
5TMbI47nQ0iImsT0IQijovrQeOKdDmpV84n9j3iWnZUc8z3xAnuXDUOmP0DMAQ2v
4bTLe6ovgUDDPjeMi3I7REtbc0nIiQfhnUMF15LK55UBfv+JE1n1bn4vJW0a8Le+
TgiLx9/Uw6Vz8L91a7vvL1XH+GkoL5NDp4h3mrRJTWPrnrH49UuE/dMwlCEN05yQ
3v9P4asg7VkT/gW9SyanGT0jw5T+QhEaH2YnFNhSKqOrDgEXF4nxu8NgsfAfShFV
u/omsKGpAhU7sMOchrzu/R/Xq51vOF3GF6NJvzoLs6aHms5OR3HUnpxxU0XHsfb9
cCvURXgG1/kaoOtd/MeMP/wlcOLuEoNIBsvKTlbioHxpDXchL5Va+cchzSgNUBlx
oBri+xdV4KhqfMynOku9JqzouL2PfuvfmXBWVtKeomBkz6VQSrxMRLAr0E6K9POU
ZXrG25kKzOGytskEPCmu/+kDjIt7cQeLqoB5shdY2Uot8AqlKUyjSl/JcUudhiMy
T+lJYnBq8+6M4aFIvEODLjBct2nr1K1xxso0JextKxgoNETPsZwbBy13FwryLLrd
MAin7t3AgfEZsKG1O0idnoStM0d0TFAt29ehJlZ13slfxAP1kN7JhFuhdz7fFWWL
KQtgjL+tTybOJA9vEBBNqO4vcrmN/Dtaxum3V7YO1iuT8l/tMJ5qqJRlIfJJji+u
zKbe6G/NazGf8ks5wI3NAHkIDhSfD//e0G+Rsv/UiHXYJp6dIWCLnrHqQfCDZBiz
wuGjAannzz89gENoZrzhd+b1rm+hcRPayECDZRmARAjGqYJzihWi6chlzm2DnxWY
YVdtQcDgpKtCXRJW4ovOW8Lg6lp9CJfYp3Xsao634a5rWkxYPSptid0Q8sYQ4U10
CLWGSEHueh+ag7F/yWlyBvc0dcJrNGVOEraDQAgODSlFJ5X7lGTKxRg8eBXYPeri
JS9eLDgfW6HBaoLPbtJQBaiSb0RPF7qzGy+2GAU3X8tEoV7ie5gv5mxQ7hrFyqrr
L26X3xoXiKMyaJU2PpLeBX7i9HRmcJs6a6O0miNdQTf2yvjvMXz6nX2GoqH45UWD
p+WZfakJLv51t1IyN7HtUlE6YssxJW4K0WarPjo7ON94TYb6ViFYu5S1lXp07NqF
mUEUYf7tSxAkOajZu7ugLQQv64ySb1MqSem9Nuz6sbEgL79fzYWfMFUnqm7utn7y
t66kCuCxpBS1Hfaobsefn9puK8+Dpx1HyrTUQria19n9QhMLSlQ6BWjkVg6cEjzm
k8cgUWQSoSSLRt3F7yD4n0/uSe8VsTChU1M2/FKcWkWLKmRAW2Bgz0gN5/2adF9q
uZRbT8zmaQuetw8Xw8KEpVGWFxeocLGPCQb4we8MjhG/mU5N+Gnc7XzDcueAWWli
XYw4IFTbTSN4/xCqVlVUNRM+LTvoUTlFLaCP9OAkBuIov7DEo2KHRxmmUvQWva0y
kpwl1y0Y3JLQTARE/kTl4BgWZUa6FHT6YP6tLzn/HuZ4iFM8hQpKWkJZPa+EwdLJ
2WVY37M1LV9eQv7mitVRgpqmHj9qOtJI40JPSw/3COs=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
K/HKiUY2rJJilj9SyLza4IaN+sPnfbrBw3+o8j2OCQPtSOb051gH6L52NYMxZufd
YaFdfVsiBM5T/94WUQVdkgRzqBRWXqSyhhSFCgGnQkAnzbxgc5yIFOUnGnER2rtq
vKXNu1otesRUIYDhwzWI3/ifcWbmxyxVF+lJR/nm/QkM1+ukHfjRuGO+x8Ry8Bo3
0j/Qf7XULv7P7KYZBTECuTPlzyCGrqM6uMhYPizaL2ZDY8yC5taqW3scDlWyGKc1
1vu41qLGq+DiX9joc9uBfNb+3FFgmRaAfrkxmZfZo7Rl2FN0hBA4oTaxpcxOMCNn
IfLhgbjE7jelTzwj1Mtiag==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8256 )
`pragma protect data_block
CLMOx/0i6RdjiPtsqCvh23SC9woraq9ocaK14hoiEptqdMSh6NxKGK28zUDehatD
xsaImffxlswiSNNjNCQhCd91Y32nQ2NO5NJdfmeTecdPAhXQVHm+lfqRMVN6fatf
320pFSYN29Q6JK6b9FDdoDI7Vq/d7BBDRPeIAuwWXqXiFG5lsCj5tSpr68Z1NG6r
FWvkHnsHrssKC7C0srqU3t+34kaoc8Wa5ZONTFlzfumah5REW0laiUlChHMnlXWL
RJhCAieo2o/olPFtaRs9kKQoTMz9TmI1eaxnD8oT5lgM4juOg0hsYHc/m+HUApm2
v5/Xpez394jzhFztf9Gko47U1l8niP5zDFW5JOKcInpQyEj1IKv0w8OatekVGycq
k0/UtjUcEU7e+UxTGN8PQ1twxxtQukody5lyQdgCg8res9hzfQ7BeArJK3YTMyj+
ZXjGX9k/7yrqyRikZ+e6bZiSAyoexsDrXhJSX9UB2tSt/FaI09KmT7GzWjdircEc
bIJNpAUPhH2OWvmmLPc+QnqN+5tXJW78UitH3WPCHWryK4dIFwQAvS9iq+m9KVyi
cDbTtZEjeRTo7Fp80IRifzpjjXCxiMTOlX4U/lcLiKy3C5FLjrPlQfGs804aMytA
3PqQtxfRUCu2P7W5r7+d3ikq9KQ2kSJwIiVPv268VJd+LLPPx2gV1ob3+yxF+ABv
ODgG9XdYPc8tuVPvnXrHfqkSOQd8jDIJ0eoxf9fPkrOqPutaZgeB3yz0dE92b3wi
RLCcaYffWu2Hy+3azbSBobI2F9BmQnuypbInKm1NfOJN/mx/HuMEce4ZnDGKu87K
bcrmRYBw3q1LU25x3ExDiUAvsM9S5Gsd2GLSaa5C8g9rnDTvPi1AGoqDqhp1+fJJ
Zq6AivnaggfeAGhrP2BXsURrjuGfgm85cRznK87SYcGP6Gc7gQrRCbVjBCa8Pzil
soYf6eAyeTMt3oZbtAJUYAPKNKNTXhCBsLj3t/pXrBaF4mJMDl8QMElqOPKSSdQq
uciVjCfAz4AiUH2B+cI5/47nDoE5BIdfFkEJm30fGjany0luhJuAtUadu1fzvBze
UYFLF1G1WUSjxrN+PSTlNPfQJPDi6RedfmCsmClGLLA//R3byD8Oo/ppx2jof7Ox
HcWhxFLAb26xv4vn5EhDlhYOnG5zDwmDmtoxvzkT1UX0UgWcqLci/8OyOEwGQtpU
MHnyvFQY0A2M7RcQxgak8KaJsCvRdzGJgUi55Hv5cvvhzPN3Kb14v7sPiBj6q8Ig
UOdHFzJgxJXwjkBSwj9MBS+f2MuQ17zYqZE6zhVVrnSX7hn1SRo3iYl7CMuwIpOX
oifvPFz9T3RDQ4cqcTWv/pHRKzqOT8kv9begLWpIxKXItHouqO2rxMTRtG+wnCc7
25sGxDRwVSijZ/l/17jJFbL+1Bcs3pnbXuvM0KdSWIi3FILlMQxb4SlBS+1/7CY3
LqS95yLHTmERauGvJZZNEA/RCxVL3BfZViAd+uWbc1t1v+SYKJRsGOzN6e2IRFTN
x6ndGsSdy9TP6I7IuC6lFhCyR++oFfawKD15+d8JFfZc1/VHHasGtXZ+iAFGvBXU
3FxCUQfw+ZcZlAWapHKhmOfFsEIbe84IeNnploj8KxwjsV+y9A3RF+7+6/U5om/y
kRUY4ZYhAojAprsh6K3TZ36ev0sLoFYxjXWKIYVpir1i/atISlc71KlirnesYjBy
E9F579hj/qzbCLltZRHeBsZyxai7pO1VhS5OoRH0z7NzQvsU2B2livqOtjz4V/Vp
vmkLAgXl+fUusSQmqaaqPyY9XSMYLRGNyWZrzn3wTbZsXTIk/G3Dh0JkI5UgMhAZ
Wrou2p61wGdVxQQI+5AhpmhLtybKiXXDoa8kd71GWEs7tKiGq7Ms8pyk1lf+BUhf
btpI3/zSJsS7ckqFN8kT/PyzU8VnQ9V4cIg493Xk11ybGFf5wLRLU3bLOX9TdnsV
IB7rKwmCZfh4C8KMDY8YCwfFxj7rKrUvQMqfJSntJ5d8COIpS4mm5v+VrClmnZHG
uepPMYCU6rOkoyTASzrRYI5i+EjPccEoxmI7jFS8JMqfYysvcf1kBdyEndJTR4/f
AQOog5qy8AYHMI8vAUqMNEHNcNM6uhQjHOGRvRU6tTKSNc3dIHQcDhWW0aL9FuYI
/yLfv6LrShfBPthFm5HA0ZUa4G9fNBF64TkldbsOEs4WwcFoB/7mucVOiXa14Na8
xYILleiN7fKCUeaoh6AdHCV3nY+whBB9NSIh9pBQHu/FlGiBvuuQxhFLJEfJswg6
xFpAd3KUyhYD1O3s2CoCiZq2Kb+jPA9qO5gGsWmsmDzo72edQLkDsrbjtywAQ1AI
zERiRIdn5t6dpmgRuXLKgFtJJ+ea2B9gG3eu8DGUYt7upGwBqlFcnGzM990SNA2W
VJo3NqcT3Sex/RtAoqMsCkDQg5af6I1EkMdMBbwobKBLh3L3QWlqmZiWZp4HjgUc
b8+bL7RHEV1B07DRdcg+JxKIYDOfeklbg7xQLkChhXM6lJ59YQMmNn7Zhf9xxf49
dGF8D3cKgQ2xVo2PGyN2jsfO3CGAZVOjJqoVX5kMVCevkqoAsUxxrfoI35WTiDf3
A1pmDWU+HH1HHpXgdWxae9yleY69o4SkgL5OGub+7Zn3PI5NGSNXWK5lzHIEN99e
0e9xVQy8gkknhsPy5NAKPgN9OgcriiubRyyrL1/yT02PhzkmdgGzy2bs3tMhf7Dy
v2Nt/DDd/hVkwNuAsBbGgMCm31VNvKy46pfH1KGqRoijp3PP6xCrkNAvHHkNjmW9
TtNc+mQLvLq2vr4fiZWG3rFsUiu/k+8VHpoJFWiwlELGY13HhRV9xJh006D0vVcz
LDis4HDza2WZ1MMGn1q/CMglnGrUsYIyqgPh/bBf5xvH40GYloWIzGVS5juHgc84
2cS2O8u+YLhR0/5PZCRfhfrhp3cd2yd7JBxYGZxr8lUOMAy6qyCQZLKZJGZrE6lb
UTF8kfVNQW1vH/quWTx59uNco4uFb9JeEGedQ+4eVOS7xzOOLXE+ih+6tnWK0lzd
6882LWqZ+e1yTBDVNlN8bjZfcpDPVg57s/nX+wVCjR/6ELhveNIDz4f523pf2eAl
5jrsbps1qO9mKvAQytdANMiI6EqyVVVX54nwgPJcyLftQ8KzpIrImJV/Yk4oEpFO
5RoS6a1b8uPckbbsg2mFoGvHktwbE1/i0WLiUfvcVhNyIWS/vmenizd4ztFMLCh9
thHLK0GOffbPfeFQy33PUkUPV555gpoGTcn6new4nP6d7OvAPkOttvVsE0g4wGqK
t8biUdNRYjRr7dUysDa6cIGmlVIovADkBVZukjJ8TCiNiRF/drTJ1wTzIpyUjWPG
ttnMeD0ZK+45lL4vARN8jxj2sCvLDzDeANK2iT1ReuMSmsqOF/F/vsI/N/3eD/a6
kyFYW1/2lB9sc/CFywhCg06+Xs6Ntp1I6YfTgyEtFMYrl7rTSZCTm/dsdgeYpNFJ
+mvY6ADoeQu44mqp9VXfOyUFO4S1uEYPWb7Gs+GF2D6hLxK4GN35wRasHDydoaWS
PxQbVCdNda0QQsTpzo1XctdaVb5D4IrfZqHkaQVYBuS+xexSVuK4ZGmKJtuaV5km
qbObnsnT4k5H9BRtkQYWds6YkjNDHbWjTqVkSk0jxegOVrq8k2r/XRMEfBaX8EfZ
DALsfXk7VpFHgnd6uXIxQSn0GOAPh81xacTbBxbw1XIiypaNPCXPOo5Qea/AfP05
O893wS6ECeaZRyx6CrcELbuM1btFsTSZCmD4oWqiLIUCy6P996uBZkkDF1lomDjl
y66CjCF7Cg6AzdAonQ1zV8Jvm2lpW6LkphAX6f2VuRBRjI/vREmJn+aH2b9KVe9W
KWyEogDtY9zVIlul3DoI8gr4M0lkf+fljWieHFeJ2V1PngLl9soMmuTcfM/bnoFn
99GKMBfLk5CxZddLpirgfX3X0CmYdjoEBo2hj1Wzhxzuhn3sZt/OsKq6Jv1IxZvj
Fjjc515ux+e5ae8jV8o6XD2BgzCs38A1RL3KblZy60ZyxDRdxh8hMU/eJOUxlrgW
4Ez7y18VcW/q/M4Ub7+ZyHVxdmGGLDzFpO9csuJhimi+xjKU/8wwCl9mMO5hlAfu
hJTV2gafo7m/qwCecBWxwgjTF0tEuFoYuTXPwNs1sqhAL8dESbbH2vxvv4lb6xcF
hyXnMYgqeQAxtAvndygIk/HhXOUhpo3o1SB/5uJWimea0T1YzTcj8h+SfcxDvAmu
UtTmKt1VD4x04HmVu8zzt+0CrilaO60tZuMyzOgXfDbzOozu9lA/3xpmMKGs1HGU
XeNi1xDV8p5biQ51Cp8F39yv4qWxbs+LOonXZ8iOHFNGqLfVmjns/Ubc6pYPhcby
0RYl7obY5+nmH1LYBgrKVj8toasp6P+Hhkjuh4MrF5tH+tJ2XFrfQ5isZxLDecrV
CoesyxqJ/6b9wzkOAcSbma7VM2pa9vyZYgWIqyJ6rYINt19rhWvZNeoLZFaX09am
v/Aef+gDhC0lbxj7C6JJo/WZBQEVLuNH4wuKRzcdHVGqjMbXcOecK94PwGfwEJbV
rTYbPPlf6W56qh3iGVHt4BafKo4a4NhLBhGJZH9U2ETFEDVlP/hSBQFKDLBaKcKv
0ekYpjALWod/Uv/IwcWhkoioARKEaCQro3EBAJZfmPeakRXpTRBYN2vBWBMS6Shh
scnYddVjMmDgZuNE+5iMkDw3WQhApBsur9lI3IMvD41X2zqST+x5oGsrdTKugQcZ
5p8qpXrqLZrQpnxJ8xJqgoZ/Ok23GBBv1HOdOBjf2M1jQhmJ2ZV8O09/H2MZEIno
2QKCbk3i0cMXr+m13KyCZTUSoN8lkZ6nmU0KNnrgIxTFx0HFCWJtnJg+hkxaLoqa
EqTOIKa/DaBJMcKWns2EXnleTyY7iZMC3ECUp9+YXLrl1RVqomoJpi4hC1NTKtv8
sRkP/V0ifWTLzFuoyjy2EyzoolbHi+2n/MsfUNoRYmJkziuSrKJFO6BEracVTYmF
kYPEPaE4qin8/naJGK6n8Q6j0hM2fhOqSCRdXkK6x4MEJ/G2Sg8GJE+AnnK7HfKY
gNcDYtn4dqZmnRH5ARPw1VMamPQSBnI6Pf5s/9knnlI0ga4uwwgq4umCNAMVabls
Y7I2uStartzpErE1N6quDECuScuSpFDh5LPKQPxisTbJ655YMMY4YiZ7TVpmy+GD
LV8pyiAx04jOP4aFyPPrBAdU7dhG6GJqXZW31ffZcPIatrykl8kQH5nIR0JylVNl
GWcK8xNZX7qPfWsDsoTNMCcIOG9ZqxUF/HqNjnep+SwOcRtifa10Kq++WKiV1mFs
UZ24YYIPpegJ0wT+Q5v+4TLQ7UXaLNqCpX77JikI7BKRXIdpxUlvdlC/gnboCzhb
nskgIeVyTQi10VMpcOSV61FuP/8O4ZlTWBDWq0dExPmKl+xDBUeJdBY12vVUSx8i
I9z20SQ/hBTphUiseorq4NL0Av0gWjHJULJFebcVu4YY7Po1F7HLHujcColjXfmr
Rm6Hyk8qNpRgVJHh2+3XfimJVawR1SgpJ3Rrl15zbhRHU2Z1QyTLOpfZtc49yi76
3Nq+rZMMVt8251L0fLMcBLtt80m802Mi2YIJnV45E/j887zcrMVB6jbfGgkK+cIV
Lv4zL191zOb0GMsKrNaQnxlqB+SkQjzXLsERJtVnFo4Rg4yXIozU+aSzo+FSos3b
1dyLinJOkSzm7AEUXAjTPLJg5LC9LlapEadlZlrxTx0uLDIy1USUJ3FtOKQcAsGy
rQ8dMXSBLn2s1mD/xvhrodTqZdNKo9WGOL33dnQYHDdxJ2YDL24+6HnAhQeb6t0V
WSIupc+cUeROnOchVnHN/2JrYoilZERIyfNLFpy09k6qtBH1Q332q8h9jK+DhJP+
i+ItxAamRIIN47OCuBurU0LBxXGwJyHxhd8zvn8n6foMzCSpyzL8Q6qvWje6QoQN
B/eSZprPjCsrRsmEzZJcbxGJkBIexnL4tdGRGUGW0cUOdWoASf1vVtHe23tND72U
Chv3c85AqvWTlh7sQwpTIfEu2k9H+ya/9BAk4q2JUWVTWVWYpYNHTWJON9RWpPFD
HF14uPuECDqFB4TUDjMCq+MyFH20v7KpG5j0QoRVaXJcTrDewO438LXPX4D1LNP8
0J8kH6X3YPjLKyBxbTPGTAny6YtcZWt9KRzUOHWnlPeQzb1AWyuqbpn9WGORbfQN
KUhvWkMBqqiSpXVd8j21KEjhVFW1qxIEgu/dpYpHCN8zY0wgf75EJ5BFKbCXCKFF
PiVlb5SEi3EeXvWrFAaWblvQ0JxpSJaKQgqsXCCh0uTB9Sr9awq+i/lmBOM63m5H
3LiTriR9CVV9ALo4EZlHk+TI8Fy9Wg0ffFDAmDgLaa+ck2dkD8ZQkVXw76xHB93w
awCuo64jGjGQAlPSdZhuFew2QeSAl5AVBBxcRMIgnojAbtjMRzHdaSKZ5pIRvvA9
CQ3RgBAgBkvpjMNraoNrA+7Y1YsUl3BXdNeKRykK1LAk6r6/tICLLjf4MwPrbwyc
ayC+zGcg++MkdpLe8xEZt+8QjE0CBAdZB+/JI9wojSgXLOJs2RWBUyNKV/oXAK4a
1UpJywr20rKt/H9wYbVe9TsivhlC5wRaJePi1F6DsjPTECGWWIttIl6V7MtEBOhf
pzRr0amUae8bp/4z5rhWyZAjy85N6skI9DmuQHx6P5fQ3YU8n5rUDG3O0fnoF4nc
i4LmQwAL1PiDqTG/LhQnaxBCGY9vYepRkaSs/Z5A5RhVNbzOmOoGbLo0Pq8bPIxR
K+SV+TIO2kfsxRmWH8wYYzajzrmp11QC/T5dp2oh+NPCUDY/w6GsbSG1hh5lmgWd
65a5QQM//8GYXmkeUrhuXj6LttkSrX/65H2DVs2bSqbwKFabvisvioFRy+HnKkZ4
velODGI6wsnJXi6U1qhr6URdbDC2ap9J0ou0Ip5tyXTYPmk2HfVvi0K4z2OSyaMx
HgcReHszoaqaDmDuzkCbveQmbWEpSVJxOtHMY61vGOt4qQajn1SvYdbe2SB3L+Dy
2qIi9zZuqLx87/ar2JdPbrInVthWmjA6uvIj53Ej4bQVwO9UDf9fT7eMUKY3C6Ts
A9bjTAlv0WL/kPq5f84VS6JHLI/3aPMuUCgGJbLtn/Vm3lSCQj3VFimLuR29cTis
5471npBCANORhGpnQINXOKdYsHclG1XJIF758yHfec5xHfkmAi4PZwJ3UGbJ+wZf
yyPxDAuPDsYG89dBPKLRySVCX+SirS8hJfPymRDAtVhtCAvSSmKQ5pANSPvnRABP
vadjkfq8wtTF58+dRuxXCnJd/1JcqpUdG88SwcO34WSiSLoRMAYKYYwnK451A3v1
MQTcakJSNLYPRObPZ0cTiaDEoItGlkkEi0+hzOYYpmSP6qw1LVIuNQoDGYqG1E2m
7RQSlzwY/EZq4fBUKQnuxq2MD126oPlGwHSRm6RYBf9KTSX9KOhzVPHgdG0RMAv8
UrBovFLdg1qqHvaNDIgFK3c8mr8GGAnEyG5z/YGhIZwtPRLhYvWNZWXANJfckpnh
GHkbt4MrhXkZxaygIPO5ga7jBcxFfYl44iHXuVJqPQJpGFVYaeGuFeymmFG/q8B6
mDBFq7ZrzKz10KL/x7xO6witYr8v+W75ges8oyFbQLtXn3cl7x6w+FPjqGLHtC7q
cZl9BntboIGDsHxtNWbTZbvl4ubUka2cw/2Jr07cpZB6qlrkoc+ANlFY7XKQG/zM
o7KS7ypRF1ZV0guKYuTfpEbUCAnh8Zn6S/0H2Qoc6wJ/VtNs74pk57yPI5ORtbbT
bbF6qbQ1PeOZVlYvZd8HkUbN5bJuM14Zgj1AO/SMdmHjlRHlSh/SBJN38GNP45NU
09icejmwaULtDLTyl5XAOW/HTkf73qCgmDK9R+Ma+hO+OJvaWdL2c5c4MLIx7RrR
AjxoP3PEK23ode640VovfPVYqWaasGr9eVmUO6IfuFqEhj0wMYkqfBPj1eypN3PD
eKvc2suIfLFi90uGo2McbHbKNa9PtjfX+YqlAHy4Xz3wXoVzCZWIyIA4hY2yyTdj
Sb6Zigwbom58oEqqJJYNcsopYuw3VgA5ELzMtu2eoWxihYnHaEcBmOKYiUmwYogE
p/DqiVWX7GULYb3i1GAZ3wWwCEAuyvemjYVxNZ95wrjuO/+iT+9zc8hlaaKLfzsr
MMG5BIZXA5VJgLdZuYdk50PI41GcYDgTpMK4dGep996liW5OrW33BOHwZgpgbR1S
fb2yMJXY0dDJf3p97TNvbGFWC0f+gY5AW3xw/98kABASDeYTSnfz7+dP4fngwzvb
J6TYsz6nznb5Cm4H3kdlxDD9QWMJplYhoHVEO9iE5zydtqmK3R8bo0A/GzqgME/d
nx0DMOIhCR+FztpIVCCsA/7txESQZObfsJXG+lAgBpbx7LbGq5bKTsFavy0Qaz03
eQKXfpFRUttMzquJzBdVcImX9Glo25zSaELg3RC2KT3FP/qt6FLa/yWLYu76HKvZ
K3aarodm1aiRWIHBRvma28kz0MRU7iIZCL0qh3mvGVUcu2Nlaf01/k9qIgA1s0a1
A3/vsajoNFIzSpfGthbwY5EB1g9uAz4+seU7RKt6NeNhlmXvi1h5GIPfzUeErFG5
CxOP8VDHtJYSrHb634sAh8DsOF07EoCMZhVeEAd5uHhzDpBH/SI7r/ikikJD5bQ1
PCTD5+bV+zC7RehxVUGMpZLusET8yRkm0VYZNlh1eq54BfZEsLvTfihbi/6WuSGK
QmY6So8iRTJ3LGlvvgS+r5biazHkAFmhvKmd/WbhAGfvs/zd+IY+3h2WitQI9X8B
Je8zDwbdj+KIVsYlFLajmPomNz1E4bfDRmwRvcdehqrbvOyoMD/J44Z5FgyYNE01
ICyRxYwdpKY+jkPIOWCR0e5wHTQcuCWcWi4ADNooijv/x5sGSGcy0NuipIe18xPW
D0a44QMQtzHmoVnqxQvfsaeRqWppO5UBtGGJdYZqtUJj7LKDLMbfX9d78tesfA/a
htr745xuBcxaHlJGcaP0BJRMr+UR8uBg1tZWiEDUhmaxMsK8wvyhC8cmcpSJDwtF
jJ/6v0x5PChmfsVi2ogicg947klNqYfIo1Rm4j9BQ92F9y53MTQGZAvWICv5hDrq
mHx9mxhqdikeXaKq8PEdyoNsERIgiEVM3E7tYsiCz4ONl8pvUXhiC/+1/ywzik0/
MCf8HU6NMcf2LmnZNJCHQE9xCbr6RNnhCZ1ygqLakBARno0ZVux67z5EVGxLwTW6
jeJgqaImA62+Ow63pMcZLjQBpHkIGkiJZgq9tz/cNWQm2wq7zqkiqdWDbs/CDGAh
XpzGcbQiUSVSNEpqs+oYr6DP9QpL8KuWFDufWEmJg/rlYjZYxk5dnhjJkLw0zYFL
Rxx/G+2Y4v8EfyEDNFvsMr0f2/gHSWeZXv0dO3msd3DamUhPXekqUQ+r0C+bCvLx
V3uhSiG+iYShfudLhPnpEVd36vSqQPz+fkpH2PdYmwQNuVGOR4bJrNsZRUxoVyXD
awVTRQODJ4KKc1d/pY7UNYzRPQy4/HFxz7rTOxSnXtrV8HY1e3iR/WkjgjLp3xRp
Y5wO9ZI8Zftm1QnON25bREUIEvPUd+RZVymZypjARcE4HhqrZrF1LCqD/pqGq33u
pxhS7dRoWFeyjYooD6tmhzARgQb52hWS9yeAIaOX9jVcEgukEkomZSNLNF2Ud76w
EUMi3/dyCavbGJrAH7aB9liQ9+PY0Jz/CwW/6hk88+AvO0eV/XOUmiIwdJDiYHZo
+BRJrdEdqv54Y25TxwnFeNrhjHURwwwKRadnoYNnHH/9pKZpq5HSdgg/U7OJuctw
vw50YDmw1s/kLe0WbcWYJ8nwvKgP0Hv/BG6lVevJIEDrMs6LQ/x5XTUAVupMyLxk
kWhTpbutoyy0VbWDgAb1TTgl+H62bi5a5t9fIhnBcPUN6CbWRo8HtUXrb/gs6MmD
cua2ey/+kY1HFmHeceaYDXAew13Nt5uzm5RnqVDPKYqv6lA0lFBTD5Zmdj/MGzzT
q6DqfInMZ1Hqc9kg/zRAcpwcInqSeEpRxSG3+GJVTUlLIL7dU84mj3ACpxkSCgg0
niKjuQkowZIshV56rAPIBTVc360MSRfnFTiD7gjoC6fZhNhg1234uQWUPzwzN7FB
wy58vDzH5k3lMTaFyi3SYsMeB2qATGOAhMDXtGTmB6eRSETNMO3P5x2MEft2aZ0H
QhVzRLd7hbM3QKtUaYytkjrc2WP52PSuYrWT/MJLLf3N0UXSCYg4sx2DrHZmV83h
xRNb6zk/R5cuzdpOE44Q+K0de4x1OD7klBel8zfTshzx7zos/hZSqCl5RLt/EZiE
fL27oU57/loySViCRtS1FV3GgAd7GDziK2Rgb2Hf4uJynUvWWDwgGU3elS2zIp2L
djqGnI/DaNeRMvE+rct+Yh2FBS0+lcrOXF6QfMxO93CG2aJSmdz8GtaY2X6vTlxE
ob4/N1ZzNSQ5AKCnGwC9SlPIZOO1hmLPABK3UuLU84DQlKB64yV06Qn+w9HpALal
YWSuNqF5Ipx6P0khTHm3Ob6GV8DAH/wr3vHPXqfMgBVk0njqB4yjARVuFemFh32a
pVpdBxiwiReIObCLqsdFqD6qXV9ty5fDJ9Pmo2dSvU3XAuSxCsNSpFvAELlfnMyy
ENRBa7eSyarDxNnz7dVS0zAys6W44RXaEvuslL6psIN1Su95qlIftnWE43J++ia3
hkTjgCNhI2/SfV1NrrQnKFQ1HFpSD5yOXgFt6flerB3647y2COk71N64mnwjoRB5
9uq0SwJU+g+uRmj3AUilhkNUSrqDEnhBDtn9nyH/8MwniQhbJoZac/nE8TEgfsPG
E81QDKdrUst5fxlVTpUi+JkKQ8w/KPYokMDs6GsbaxMG3naF7zdYWIPh40brz/JV
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Uh/As6yCv2pRaUyr+r4ZBS+8uvitRCSaNyD9BNUjeWbuDEy5ZtLx+/1+mdmoc6bV
7mWpr2y3LCVYbv/WI4vhCsJVeR23h9UjNpiz4Xg8aewW0Bs+NTXTK4eZM5K++Fml
dYOkmTy9KHx9fhVMtdxHRaqhVrLge621Bi+Gs60FrgJvVGBXluSOZFThMSENf26L
VbZEAx7pDqPGO2/RS+qWcnVTdenBFO9u3qDyfGJKz6y4z2v0hoRC3ZUu5EOv5vP9
4Ynm/SfEtB+6zFtmQU15mVanpYpqtWpjjNUzBzM1eIZsQERionTi64v7dpbxvqpn
bGYvh/Zw+jY9tI9FNISLeQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2672 )
`pragma protect data_block
QVE7UAFJ76WqjadnfZp5TF2kYoo3FAxw8uL/ACyBT4Cd2GPU4yEMPuyWbxAQ4qGP
aVPc/hfQe5tvf0MBK2vTsz2sz1zel9xazsv3PFfeg7CYjr7HKtZo7SClhcyYlF/H
fmXjDH/KIcF3LszcsV56xB+2L/1jQzZEz7oVzHGjO55NSDigq1BAze1skTV8aZHI
Egbbrm0pKYp8xW8QroxmFDJNtz0vD2rYl75Q3ycuBAyeB7tk+QDjxi3CSJunn+Um
PIMz/uuoEPBgj5iNs/NABIOrovLz2ztrr3neOqw8X4lvCKMpD9O4dCwILWL8RQm7
qeDQNNwEkx8S90LJblFE6potRmLSQziyj0xCary7XIAMkaCEjCuphXAD/SK4ybHY
KYf58XlP+CaEuGeFWRuDWA4nW+LaTGm4NZkIuGf0Xo9dd336SJ7Ky6RXB8p7fvvj
nkY7SQMke39wAQqqOkoD9h4H9eq+LWh6f8++3Si4k6l8UgVrJDqUOu+qoW4yg5Pa
wlHC4fuQu0+JYQI/eJbV2i9cvcq6AvcIBtgkR8YBsDNQBH/Iv/MdMdfcZfNIx6f1
/xxOdVcLayCo4VVxB+Qu5Am9fhckxAAO9PgPSWU8PEY628GBgJ4hwG1btULAaXm7
LB4qCuQOc2/guKEG/ItIHE0n2DtyjAXnzcW2/mIty2R0k3lP2wPHCU/6nerd9qNa
WcajQiTfAn+S0yy2OBfRbDZoRx+xYdXjJiOVNjtOy5s5ZfZXtMlJsUynVS+P/pZI
94xb1wFerKklXjK2hiwCGKh8lxI8XKfQ0vtuuiMQDBtNayIpZHCeaeiS5Yv8X0Q9
9eBrpEg8beW1S6Ne7uUsrL0KXj9hNzL33ZRf0ahgMdPIFcO8+pH/If8YHT2C5l84
/m3/nzTKA0QD3qLxfhr6b4jlmVMR6lC7VqkcHyD3Aw/1fRbMelz5X69BC+jl3zvo
RWskmI8pLTr0L0w7ZW+E95XziT/66nb6WxV+DH/qIGkj307bupi5KzovD1sQqtu1
WxMuuRwF2muBntVQp+jQXM14Q4VacP6/xcjwMkwlt11N+IFzLYZawk8aU/hfY0Df
kEkAIA1sYvK2bSB/0FZZc5HPGdKvY+RlddLd10+VqBHa+nAmxGris8lWrurl/aax
aE+DOlFKbks2to24Kz8aXZ5pFGzByH0w8pVLdc8Q9W9H9lYiUfHwn5gho8nViRDO
7EtggCu7Zyurg4Y3O23+IPZLJAzfFjPp5quTCWP4WT2uqX2yV4xNt0uCN167uCoy
jNRLsSmK6KBahy913l8d+qRwNJ/gCnjs08kOsb5UfhamsblLWUU+gwOTlbbJufAY
wLDD4S90LY3dfTZisr4l4YVX+DNgsJzIadENN44StFzoS3DzxBPTR8o3QDXwHBd1
A8T6NIs5FEWCAzidRfCiTW6SOubGONRATSyokpmdMfnNUmA5qVUM8ZSj/dBj1jwm
twr3A3geOjCt/Do6EP+yhbtyvyyyUDt0ttKL68T148k5UNd8wJ7ECNTPYJNqJ5RB
0cvNcygu/Fh5T7brI+UZFgjbXc9xQOO13uv9By+FO03CLnoBwc5pU1xXfnp/DAaA
EpICJqbzwO4e/bYI8SkUonkx+ebz6OKDRqnzW4Wz0M6uYxigYJYiAE9pHYdH4ChN
vLoPW6u3VArA3/D93sk9dGE0ncoUbjHMgoDvDdZd4eWPOXuHq9GUhMkWinO9PErs
HwQLDNKkcAsI383nopG8QGUh3waa9Cxtks3zlQqftXDzsEXummZh8g05ZEmyqc7c
QN6aNFKsu99iuzw5K7FafCahK9h4dhMfq9MxT/EHxP62kCCZ7uJtwlg8/wpUNfmy
3vuA2tkRps2Ehm6kbINj+TqxUHNtR1jkuJ8gc+gV8IPrjYxrJuZkgxx9OsPWisBf
VEHJU9Vc4l6S9kb0ECMsNQz/WQs6IqwLxWCjA/JCmH7z3HWrx1+Ht7c1QA7TqMNu
3xhagSTxvni+j4yXq4ntbnKyJoTtJzfJrdKB9rMvRkKvDCRLTssC7OtfLCInB7T/
XeDZyDeFczbUl2hv1Gk0EZAXymxtLRygjZws/g7LNE02GOkzvhIuuUs6OOG11c13
oqL7iaBu/hflH80HaXUC2Xh6yD8G4Z89/ftYoTwoqrT1XPyaZNhkbe4wwhWq88xu
kYuRyOdtzeQa6+DWo7pNtKN7g1dD0zWe3a7/EN7tv9tEoUoleI7poVH0j1rCcAkP
JjUl9AewN3q56Or7gU5LrmHdyT6VLM9xqwG8jU0FTddtOI7tJRZpW7eiCUgJUNqK
RiwFEA6MK7+xr3LUhJjUXJbNYx9wwFmXDxptBiu0DiQhAGcWCM4StQeZsUELaijM
eRQzeuye13usgekeUMyxWygrA3j2sMUpVUifSKWxXYVCjvtgt9nbLYmnbk/7SAym
MNG8GDcOG4IWoQyiW5ML8RJ5lZ2XIkIPkFTFabzZr0VVFwlyNOZ7IZIujJkFLSx4
M45p9Fg1uiinQLZ3i7KbJcPcMQmJLACnjNwjlQrilt+hpA4Sif8CXewPgb2pBEwG
QeKY8ejWlaFlvWP+wRo8NBKeo+IzFVeI702Todj1gUvWAOxlFylePAucd9aweIxo
9Iw/TtTbotmlWcjdhoAroDKC1Wf2VDb88ihcmepCSBex/dq06mvOrJLxS/ctT/cm
tzQB12+de2eUWDgupfih3FGvmmyENhuG5hAa0Y6YbgVvf0DTM6pivEE9NhpsToDN
VV7hxAVepHTsXz74SDAEPj1bttPdIAiaYMh9lfCH52CPxhzgeqq312b/V0tbeZTz
EByOWVqBRneRoZPmuOWWYOkSgYkC7erpeDI/5Zt35E9JQchyNDz5JRPUtF0RTRkW
XBCTiJZV5rsaNTPWAWhYC+6ZGnJKAG9W4oswBeJocU4eLB1jf/hhlxtGNzBgffXJ
kHFV367WKGtjOSxxfdsC2cSsCi+NuFHqG+PThGzflIq1C8qqYgu6bw3srVCLHCu6
ULRbwqYqbwachbzejaGtrqknLDkEup52siv8gikgH869eV0IwpIMDbUkTk+MS9d/
x48bCLcoButJZCg1eKY0ncVw74prxeRWoNGCMFrsCd+neZBd2Hj0+zIFPQSfZX+f
tIkduUdjw/N8tL1EJ+7EG2OuNHmlSiKfUvrlcuNNjRAmeVwsVwdUx2umcpC3otId
m4Be7pZ+TgC8yTxlcrP15N4xD/f+JEIEpBuUGWKhJpUUttQedntFJGsaRgv8YzWc
W+T/FOec2lCirOnGmwZn9k0I4zT6J0GpRHqZnksquhpqTyv8iLbG9hdlkgEPo0Y9
gghrJt8IBGftlYAytBbJbiWJCHivP6FwZUi66prdo6D4ctJo2IC2gXfNGytjAsnW
BZ4i7hXT9P5o2yUZfgGvCTceW6l28wx8YSITHRZ6yxtcmn1e4SqCFiUCR8rEPhr4
97s+WZVDQGja7PdWpVp7NefqNfAA7bFZpSXobq6K07/8CtCj0eXAsSUtgruHDP8s
9IA8ozeqdOIHkQgImybTPVFQ00orNiZc64A1NqcJWL8=
`pragma protect end_protected

//pragma protect end
