//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2024 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = tinyml_accelerator_int
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Fri May  3 16:50:37 2024
// ***************************************************************************************

`define IP_UUID _6369abc29ec94a5fb8cea8b396f4b8e4e7fd21c4
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)

`include "defines.v"

module tinyml_accelerator_beta #(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 6,
    parameter                       ADD_MODE                        = `ADD_MODE,
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,
    parameter                       MUL_MODE                        = `MUL_MODE,
    parameter                       FC_MODE                         = `FC_MODE,
    parameter                       LR_MODE                         = `LR_MODE,
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    //Convolution & Depthwise Convolution OP Parameter          
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,        
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,        
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,        
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    //FC OP Parameter         
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,  
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE      
)
(
//Global Signals
input                           clk,
input                           rstn,
//Custom Instruction
//--Command Interface
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
//--Response Interface
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
//DMA Master AXI4 Bus Interface
input                           m_axi_clk,
input                           m_axi_rstn,
//DMA Master AXI4 Write Bus Interface
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
//DMA Master AXI4 Read Bus Interface
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);

`IP_MODULE_NAME(tinyml_accelerator_int) #(
    .AXI_DW                          (AXI_DW),
    .OP_CNT                          (OP_CNT),
    .ADD_MODE                        (ADD_MODE),
    .MIN_MAX_MODE                    (MIN_MAX_MODE),
    .MUL_MODE                        (MUL_MODE),
    .FC_MODE                         (FC_MODE),
    .LR_MODE                         (LR_MODE),
    .TINYML_CACHE                    (TINYML_CACHE),
    .CACHE_DEPTH                     (CACHE_DEPTH),
    .CONV_DEPTHW_MODE                (CONV_DEPTHW_MODE),
    .CONV_DEPTHW_LITE_PARALLEL       (CONV_DEPTHW_LITE_PARALLEL),
    .CONV_DEPTHW_LITE_AW             (CONV_DEPTHW_LITE_AW),
    .CONV_DEPTHW_STD_IN_PARALLEL     (CONV_DEPTHW_STD_IN_PARALLEL),
    .CONV_DEPTHW_STD_OUT_PARALLEL    (CONV_DEPTHW_STD_OUT_PARALLEL),
    .CONV_DEPTHW_STD_OUT_CH_FIFO_A   (CONV_DEPTHW_STD_OUT_CH_FIFO_A),
    .CONV_DEPTHW_STD_FILTER_FIFO_A   (CONV_DEPTHW_STD_FILTER_FIFO_A),
    .CONV_DEPTHW_STD_CNT_DTH         (CONV_DEPTHW_STD_CNT_DTH),
    .FC_MAX_IN_NODE                  (FC_MAX_IN_NODE),
    .FC_MAX_OUT_NODE                 (FC_MAX_OUT_NODE)
) u_tinyml_accelerator_int (
    .clk(clk),
    .rstn(rstn),
    .cmd_valid(cmd_valid),
    .cmd_function_id(cmd_function_id),
    .cmd_inputs_0(cmd_inputs_0),
    .cmd_inputs_1(cmd_inputs_1),
    .cmd_ready(cmd_ready),
    .cmd_int(cmd_int),
    .rsp_valid(rsp_valid),
    .rsp_outputs_0(rsp_outputs_0),
    .rsp_ready(rsp_ready),
    .m_axi_clk(m_axi_clk),
    .m_axi_rstn(m_axi_rstn),
    .m_axi_awvalid(m_axi_awvalid),
    .m_axi_awaddr(m_axi_awaddr),
    .m_axi_awlen(m_axi_awlen),
    .m_axi_awsize(m_axi_awsize),
    .m_axi_awburst(m_axi_awburst),
    .m_axi_awprot(m_axi_awprot),
    .m_axi_awlock(m_axi_awlock),
    .m_axi_awcache(m_axi_awcache),
    .m_axi_awready(m_axi_awready),
    .m_axi_wdata(m_axi_wdata),
    .m_axi_wstrb(m_axi_wstrb),
    .m_axi_wlast(m_axi_wlast),
    .m_axi_wvalid(m_axi_wvalid),
    .m_axi_wready(m_axi_wready),
    .m_axi_bresp(m_axi_bresp),
    .m_axi_bvalid(m_axi_bvalid),
    .m_axi_bready(m_axi_bready),
    .m_axi_arvalid(m_axi_arvalid),
    .m_axi_araddr(m_axi_araddr),
    .m_axi_arlen(m_axi_arlen),
    .m_axi_arsize(m_axi_arsize),
    .m_axi_arburst(m_axi_arburst),
    .m_axi_arprot(m_axi_arprot),
    .m_axi_arlock(m_axi_arlock),
    .m_axi_arcache(m_axi_arcache),
    .m_axi_arready(m_axi_arready),
    .m_axi_rvalid(m_axi_rvalid),
    .m_axi_rdata(m_axi_rdata),
    .m_axi_rlast(m_axi_rlast),
    .m_axi_rresp(m_axi_rresp),
    .m_axi_rready(m_axi_rready)
);
endmodule

`include "defines.v"
`timescale 1 ns / 1 ns
module `IP_MODULE_NAME(tinyml_accelerator_int)#(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 6,
    parameter                       ADD_MODE                        = `ADD_MODE,          
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,      
    parameter                       MUL_MODE                        = `MUL_MODE,         
    parameter                       FC_MODE                         = `FC_MODE,           
    parameter                       LR_MODE                         = `LR_MODE,           
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE
)
(
input                           clk,
input                           rstn,
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
input                           m_axi_clk,
input                           m_axi_rstn,
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UAPD1Zi0Aa9wTVw2r7BxbbC4XIqKjKlX4pUtQMw/qTOkypIg9goPUS37cPIITfdn
KJcl2RrhzmtzYjfmBDnAFQY3sD0c5QJOJ9zK2X16AO/s14aseljcPGBpirklAvRr
h+ru4Y+TB7PhWRAjmbKYd0hy451CPYgRp10WIm027y7i1NPS7aQGPS7tK5Bll0V4
4eP6oV32mnWpAve64xhpOBEdD0yYuebp/FbRZQdN2ih5T8LLhK+Oi9G0mLsJx6Se
3or7G+vnJvoCviosP3qxgvGxqpWr8qwu81T2MUvzAqauaNuFpdris6S7vcs+X6g7
hfHBzxWxzWkS1QvfHyelOA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 56832 )
`pragma protect data_block
jS2N2si8YyBh3rSe2s696QiDgfX/XlNqV7xwKAAoq8sndQz6q0RN+5PvvbByzgWQ
+oSltKlZULR5qyzBwEMZHKhaKkikYJHQZzHy4/XYjFEZBUaXJ6r83w1ZmY9mE04m
nDOq7B1qVxn/oweTFUu+ZSX8rJqL7wLJz86w2ZHTkPCCKGb3oiqno1tjlYzaP6Hk
26Ihl7k9xwkhK6tvURRpZntSWP+W4neIhsvvKhX7271N0vxQut1ry5tViK4WSsL4
0hY9NwKL4BPjjYlswyz3YMK5D46JwTNctpcFoCUV0/9UOFsWDaIeoBCcsVkP3m9B
QPSmxa94ltaEK5vrnbqxDP5NOspoqg7FJ+HGBDUzAdNNKDzLbWC0wB32z7jMi4ce
74JhGYGuKwhJu6ptAPVOmrgqD+pvz/f3SoCiEC/wBU+76o8dBUUZmT6j8kP+SoKW
4CBalnxcqpp1GKpbrXQSc0cAy7dsIzqkilHxZybOucIgg0JpeKBsCngFTnQcX1/K
yp2WCXE0fZz0VJXKb+wkeLtZtXhSKyecSLvvuMuAAJZvkr101tNhgOadgeOCLHh3
fU3+wCV8NgThRt0s04Eaiy4k4smranBvgmgKehPRAWo3GpvBLcytcfBO1ICJzt/J
rfl1EWmERdpleU3oG4DpWoh4lT5XtEnXTTgeFfvJ5tq3V6bgzy/cS8Drw6N7BosI
3ViKvoUibkmnJ48oGsAUnPAbZ1OAysbIMneSvajQu+vI6DDTy4hso8eHjpOwyHDw
xSeFmDinJLYjkbYLvnngbOI6nf+WMara9eJ44GhqG5i7RSZ27DdDLQKiyaUkw6tb
nuQTH0GxWTlrBTdGtfJ6TVp66oXCyX0gJHffyKBm6vO5EPqG4HzCAc3mDs//QsIa
pKGOl8qLZ5Mc1iyQt9GhbPVaNKTWRWUecwMDAhMnQTuUmru2bJTky+H0qo6He4jy
6+xFzfLVAB4laOsKK3PUl+FtRdDmOp5KIO82a3IhMbw2ufkHYfBzJjavAVrXPrcU
tL+y39ccU4p/Zg6euDgN9GwT5+wlDEgz3zVm1qSGYashH3TNBzPdb4JgEQiBlvxZ
wm3Vt+9G1sowPuGaWYfwAzdy3lRvzL1C9gYTHgPD0ovZ6tIoqwFIYW2vkpIfLOyV
CT/8GDmF43BkPf3u3Y0gHTgT8zZ2U+Vmi72n8JVoThEA6Bf+/ji5z/U7hUEAn0dT
i3Zi7nnjAhTj0gSDzEW4v25wQ3WYMSMqq2LbSkxMF3UZhBQ7OPW1YKkJsuMTLEDq
5rEaE8XfsTMNmFnrLtJXoSqiKSqmg4K2zpC0fJGxy8XjqhiAhYHdM4QUhqkhaHLf
T44HCpcAxLQ/IO+u7oUydBpL5Be9DqDcJJvuIULB0cS/V+dF2t2iwOWLcHJA7qDO
/KE40S3Cpj3uGv33jyhWNaetvoj0F5DWhYvzg2Ie5xW6R6i6Y1qxHI+hNr/0RNav
bwv6oIdg8eulHgG3f7PDDJE+AvV1cow4dKVOYj9t8gQrCNi8yyB6kfqDyBb3mb8M
CpRfr+xvpssXdjNdK6nNUWHvNonIHSAfEH7OVzdLsNKvt7WaGocA8mSZbNCuGwJ2
/p3V8/8mxlexURTEkWThxRoGR7o1//qJkoeCS4lY/2TpK6sT/VOwo/JMyX5KLzum
KZtIySfFYC4fljpfs1rE3HtM6arWB8LXkP1byLYGKrr9fq7aTkVGclvuFTPJk7rw
ZPq0/ajmjVJOi4XrGdbQdqRqmFNtQExb4fo9pLiL2ZNkVPpJl8o9yjJbGeyImccs
GSftWrLcTqMQY2fuBThZnEo4u/k1fFey8Eu0EScND87pudGnVj/MZpj8IH/k5Ibn
o2hFdg0KKnnpfmrdbXkCtg7MAUcHqnti5l4YK8jBsSM2GNDgdl0F3s0kh83WSC66
CrxoqGOWQXO1agbBVf1iee/K/z9Euh0nYvTRnEHkLLElw9t8PExiwIOiI4faPGb7
B9jdzk0AvOq6ufAFxA+2HMfBj6eediWfXLXBsNpJCrYWhGEpiATeWR5MGW6fr5IY
kubH/qNvfapWYvi1SEc/5WPPyq4TKuPH9jV5BC9tNzGn6TY3N9W53rfPbacDzNvC
7+cQ0istACwcproeeGeRCSS8s3wyjkJGelaz5zzhoiCir6ONVk1ZDXLciTx7q+zD
x3MwW6e1/9LVc73Z7oEDuqoYaEdFw9CVJ6xAoz3nMio9xJvhjaYV1Q34bC0aiDbz
VLez+w5VlVr3OcuD7IixxS5R/A0jD0PwwHGdMhfppIVxhdmS/FLzNmhKORdqH1kF
SRWaU8Fq1vXbAUUhnCgTS6cx155pEqkIJwtc+mzIJHMyo0yEe1ZENbpgUKkUwLlK
voGbQYHBsREp+RswFbq0seurNOY7t64LhDgw3y3DacnXh3zS1j9KDsP0OlEG/0A/
3gtpIVQWhlX/UK9GOTdq96OrdUn7rPKETIY93K2SZBrv+DUPkSqeO0NylSy1DCcM
xFaks7dUTWgu7eIu0M6w8bOV4cj0KGK5Qvno70bd7vuayOWXOnECDb92jqveE0Pi
zMlrrgjarcx3/3EAPq8eKHPp/9uVlUXn9kzph6kryMW87z+39CECPWzy4L/teHFP
3O2fKot2bcgGwfYAiPJOS/M4YSRQlY60KHpGmYixdv2flqnKBuSgnOVeMvjstjC9
NMlKrr2/brnUjlKOFpRpg32s0RQqaKJHwqstw9K7gIMS7trSFsnFwXII0enZY5dI
p5UL8SrE1o4ef/NpP8ThcJBV8oF0/h6aBzqjmK116wgC5U+cXK0+BzucJ4MvgRvf
gR7+pCPM1ZGAipnYesMhYr0kWeEponJphcV1GPlk7jg3DnhxT3s5H3KHLKR6XH6e
dynW2ofTUUJdmACR5er9/tiBY4v2Tp6fMjCArD0TAAVCd6hwQ3MKRJ3BzZcWy/uA
Y7oU3bq2D7GUPf2NlL2LKnFlH/oP0AlGB/K8wSyow/Q3KBze6/HLxCYCIdm4wqtx
81v/RDwaCCMoGocRxa+WBSPE05IXDLLGXBlrWz80Q6aIC43cxaV9uVWC7kz7te+j
/2oAhHNxSJUIsBMMtW1SjSuBoqsHCvElM9drd2pPiNrlBd/TMPJH3WCApgpe6tY7
fkIAVTGUSznMZ3jp1Z3Vyd46e+KBaanY204R+pCt+1qf3lVmMs8mAFTQZL5QtMFh
H9xvXUTP80Kmak02TFLKeYjiftvMzqB9kIYl44bW08Fysy2O41o1BjdZoE1PpS1y
V8Q6fD2H27OX4soWjRkbM9EWEGhaB5m1azeSrGB0KjHwAQ+hmQQ3RviRc18rWmE5
BpKfJFlGx+rZznuBhqk4kKM1TFjffUFWgfhFHBJwQfHSKSLEOuF/l2SJ9U/ACmnz
5fJbHpYwL+Dd/lCScvQlt8UoR6Xu9PAsyYAmoO++BQi5bvIKv11O5DlA4udoxkzm
/+eouu7rCADChuT0XqHo0Fen++qlU3irfJKW/rxlmrhm2BQGHxQa/y8ohmt18mHW
uvwpqFfHVDO5qoT4XUA3tURzaf1pJKq9d8heI9gHRqOwE4yEjvFdZuKclvgpmDRJ
pekIMqD5qcz2WZmnVniC2wC7U0fw0YFLXe4kFRlcXKUXq8RJOMxFH8iOMHEwHGVq
VqyfEyEOVcHKl9G905pJy/dtbWcugpuHc+uDc6eUqE0AKF3mqy8FWezOAcwFcZGa
6tr2A6tVY0mOoPXThLPwHX+dg22TWP7G77KHf3ll77SMGdKG0Ja3JEWLS+RHHNR2
T21gxe6l/2NTh13ri7jgc5VJDNlLmFtelM/OF3mPFOaX0gOerJcGbkCWBFO0+dJc
m6doTYPtafRDIVCPXFShSUgnx5AVrpmChgVlBQ4yTMXRwUOGyfCD4QpaJh6u5bDA
XiBMoqv0pSGp97R54qnYDhvYAnf+H6zOMu3hiBgysGYJ63pk1JCfx0INqChYlR5S
jzr36U9kA5L6ZEcSWhxUqi8rqh6nRSHQOpIOoJeNl8Lj7noe95ViM8ROOWkv1JVe
VZRXCX1jBqJjO3eV3pZdWfqzMfjL8AkU7orsBaODcTC+rzPxgiim3eDIeiBuV64X
xzHF+DpSv0H5venPk2dHuV8tLynqe+lnA4mD/1xLEN96s0Bc/rNjhBYLUsfAOm6n
XoTmoXoZWRzrXBq2J1fpL2UwW/QQfMzB+BwzgbNoTwDvH0Rlgf7DMZnfIpRqHvHY
YEyzE8d3NGhsy+YfXPQ5if3FZwzSzQEk9c7hss05lK/MdliueN0D7F1LgjEdk9KD
QBIi9JqEFwOPEMOmlSXXm/2C723+Tm/uwrtKIeYW9ccxZ8AG+ClP6m/qnQkoGfiE
rEbhLJtv+8HGRavr7Y/8K0f+Dg2tWuRnFo2PzTGXTUex9qhZAw0fzNG50G2hdeq/
3sclys7XoY0P4HmRpng0z4BXCa1xhECnjqLahKNcDGFeqnXAYd5Rs2vtqbC+mQ+t
0WwvlhXSIIU9f7RVHcgz1Dlr/PBGOv+P/9y7IdQD2n6F1igH3/H6J9wVbgT9aq4c
9xp0aOk+pjN4tFxqkmHo0U1hQ2NPwxrWLniBaxFBKWje+UxLbgZvqIJZSIQ7KtpB
88FwzBQWFDqziCU+LIyVsXSxtSgRMle8gNfhoLjWqCvblvx28rHh1SD6aGJzfYZG
RhiNmhlpgAC3yXaRHOsOntixhXM9kGn3uYInYAeCrD70eacc7e0HICbiSzNAGuGX
2xjdPjYrKE04U13ocKTqbIK7HUi+sZf8PCguE0rcjH1X3rCo6TcJhaJST3n7tT65
UwqpoG7cY+QIDyl4Q7JhmQMyohuqvBtUOhxe/qNI1eSRUw2vFgl4Ois793NN6H00
NmErtnymI0PyleXFwDSkT/YZIFu59INCOvDLjwVW05LzKwzVW0OozOnbczcSL9uT
6VeACMi6TYpQB8UPsyyn5g5rfi1XqJ06GTIVcycHUEkbQMEYqvLnw2dVBrViTNLG
xqx9NsLuqkKuR0oCIlbMNDnJVexqZKh8kfJqSr+XtzBsM247KYPbTbDYi/DWge98
T4Hp+28D6otqTcta1zzgtWIqzrCmWRILAawFYjunZsm3DxWDwaIzF5aSs3IxuPaT
/1jLCCVpPtkvSIE1v9WhIyTTEuyKCALF8HgZPGfGKjOK7uUovSOMJyULos4fkyXe
RVJAeEfkmdFw5wqCt6+SOLrwQRT9TdTS0g0CXIDHWW0wDeU5xiGf8QulzthwTKs/
54CWB4uK12HbyKFmKzPKd0rEUpoxxAFjJw5Yqn6IhZ07r23geoU6twceTOZJNJUh
OgWV8A9Li/wfvFltTxSlunlyFUTNC1o31k5OteQ534Y5d67/ar4iIKMvXq31qRB0
HGw5Dep3+KG9cWcKORhOkqOCb9N1eTSzmfhPmXhrM3POmqZ2izUCQHrZsqAGOYCI
Wgpmi+x3h20ap2JLVJBjWyoSg2dJQFIyW0t57dmxW0SVbGvlA4mzbnXinOGJsUO5
qwOz1WRWeV4fVTtsdThPY5GtpiF0uwRoozr4zQuKeuE7Cu22IcKGC4sRjOyaTlbd
7IIFDsvJwPN8pIvntHiJL2Jy6YBhzsHk2RQrZWk2c8GUzFwtKkmoJxQqBkZC8UMF
1vznAGNf9BtqmA/nG74egKiidZf90S/rbUt/eq5l0dXVBrpagw0KUMWmTRFdglvl
GGNWU2onHZtUpJYd/AcquARzv8GWVUQTPgVHTCyuiAHuEFdPLdtU0F8Rp33gxPPF
Sst03aQOBF/oLy1X2D7KRixOahhVv0wzu6IbnsB63y3G+OMzGo/o5Ks5vRrak8tc
T+Ud7/2Jv8n5NpCbNL+ZpSQxcJyZrnnPVp9YvG9TYYZwHRzk4JQnpyV+mIflDlkF
933HBVxNWejSSu0HHlctUzgGWqaTXAIxYq2exVaO96W+82HiRiwmuFfl3HvWzRrE
UUAhCLtmJrPRQB1eiTDiNJS4Yx4O38+LGPLJPSasx6mfXVSgfXlqBTM/QpsZR41p
jBtHpAUJWOzsrGCLMKIC3PehnsreXwbb1o7MvDq5LI1zT3GLMID1cv9hmDJNh4C3
4Yk4Xu485bP8OEC/0Vy435OVUni0v4A6TxUN2poJL8RdtOX8sNrI4uPHgQbNP31b
VsvNYB8WeC5+WW/CZ7nKcB/svXpJLC2bV4HqI3AOEH4lBTXCYwZdtIR3f62FfXRF
Hc49p2sO2bs+2JIbWFke/KKuiKSGVypaNTLoEQBNnXJ2B2PkiaX8JSbfGIscOFw0
jHBBbM/gbXrZaVTo33gu4JJHXV54u22MpFTKsAzl0AFQwObxFVloyJ5CqPn/RymI
9/zIeL4Awj3yS+xA8t68ShAARsiiioTAvAO9GVTnt7yLKRMkUb5R01/KDePmBLM9
93M43p9fSlDB5YwBfFC3S/3ilZ9IVUUaozSpPZnQScOn60GyyYGdjNczFbNoc+kI
elw4E3dA6qtsm+8MH+M0/2n+ZTm2KvpF2fJFLLBqfsY1AFnXDDjVzYGg5MbF9L9e
bgLuRUsD0cuW3lSzGeRtQwkHetsFa9lz5Oe6elle/cq1qqU8gWwGrt/Cpn42msqE
h/tRo7OtNwwkWe2C0aaJkh8jb4cpGWmmwnzycnzDM8DLgrzDCcAliOGcaV1LDzum
9mYfxivXCEyL+lJdYWPqE8M+/4FgXLNo3YpkuKqNXkxviChJMRNs4KRo1IFcYK7T
GT0Knhd9WG/75jKqyr+xP2HsJ0tKesmAcXvQFwVhn+uliH8kLMHBlMV5t/ONJVOw
eBTcQgGgyTPxUlHGqTzfEr6YGXHemuhHhQIozeepEaKILZEeX7ObApsBny2h6cXY
XuPT2HK5uT0syeV0cFFWRPiJpTa/V0Rx/xCT05R1jW8W+DJ2ssfztgKNhyrfCx+F
n4mQilTeVpDtLWjYqduewyLMI/LW788yPs3/bWx/RxB18qPVnY9srgFkq4IVYira
APOfVNhv3UEtGJ9zK97ZGjaHP5Iqr67tXB8Jiesrccu7IM5a8EJ4hFmcc/TYGzrm
7ef8kegRl60g/TfBuNX/dOESgGgAgTSBTrL3torp7+S+VTrFKp5yXWRSDr+zDuV2
aia7B0CneBsuu996RP6LjXPpMsaR7f2sVAaLd0WHm3yBdQ1cTPsfelJaCmnuEEeY
wFYpPnnItpXtnR5Jr3we8EvwDVY8LPMy0xEXsm8uLZhsuWcKFceDTqVRwZP3iCLo
zQXqVhhHJ7zG4ZVM4RVlQkK0/N06Pbq2VnYsjVlVRRxLOGWPq7BpFIGAZBQVLtOe
tdcqQaYxC0GSrZ253lT1otExOBf5J3Zq3bMhIWP+XAHvm7ARnIpCOkgS/+SiSmVV
a8hyrzaek3JnF6PibsO/dd3qGUNccxSma8ih+nbK65Tra79QuSROdu0tQp0xBzH4
f5COlN6MHMihqdR5ej9ki/6T7aSeI0FjV39M8KVcYtIo9m4D4+ZvrnnhFAmp63dK
H2kah9zC4ps8llMvCIemAAiaWAEgXN716VGkoIt8SChR+JWHwHWUwAIbwDPA/Jpv
zKcaZzpLGZXlVMwAc7K6ITeMDsILj/ItUg1ndPo9AKwOChphfEQDiZEba7Gc6s+K
5j1tAFLO+DsK2tsjjR1nVfXnEl/k96pCJRJkHm7UT8nU5whs+laxbFoLuN5VvNrw
WWig8Ifz8lXmbG1cbN9DQEw5790qrAXUwXr5UV1wKtr3wJr2/C038Ui1UGfHyPaS
4Um5IpTyzs35ODvB9sbouGIXB1EfCUJ/CnLRC5eWI0nhjmSo8bIUkyfVcNYemfAX
NQKOHeQOOAxdyZs63DgVt84o1IffRMqgWOngsGrL86o4GBiu94tyQgkwaw6ay4bj
WT39mgJxfoalxuXZ4+lhdepJ/hQlSlp/JFlKEgpo3lID6Wm03FCmyhjTc46r6Yx+
ZXSVmo0iSrUTmNDgr6Fs0Uap6wNw/Aldsz8bYrM/ZJYddVkmIeBDVm2nB+DFgipC
JF7roI62BD6rz8YMRq2m72jBlitJNj0T2sEHh9hBpLFIxGiv+4siNIHUPlMhEkEL
EBnfxwUk336LkNTqIqh0QTQ1iVYBk6ur9+y3NYvTvY00aNfGy3Ly60vEbs3C/uOv
KMdCc1vtFrHPYCdrEkWiZl9HzE5y6iMqGIGsIExkyC/wp5+3uVQVAox7YXy/crIj
B/SnoRmcqMYrSQSKgHM9DNHyLNZ09KE8hd5n3mtvqyi4XoJXH6XSxs+Yl94DkPp7
BeCcWSP7FMxrIQ6BTWJMohnt5GwSB4kWJaX3/PnqMi9QtEETLhLrQhXmYnfR/nFe
UFwQw9XHPESLu4cwNjRbHpnK/3LLugWgY/sPQbGNwPUQf2IwXgdrE3kly6F7C4nv
teshCGQWPfQuAePUIfCgFeRShmkc4VwweOEmul+d8NezUazmxQ0FjstZjZWepspR
leEnvixBUy7ahGAbLf7MZFQgPj51hfl34Wna4Ody4zIqiyl3WOpFJKLsNYhPXLQp
TmwM5riMVfVIh2JhVJMcbGUm0P1pa4iR9SsAfYvFltnF+v2dtFvqP83ahGSHgWs7
wDFcBPvD0ErHVkpl1pHzJX9CcTNA5w6PukEO6dBGeRZm3slGivHmWV39KTBuBegP
n9cJ+boo7U6Vvn5+Z8pBsUfwinAFyyL7jHMzNVSbNwVn1fdacWdjFi/hQiact1tb
rqktsBmqEv6k++RkHbDgW/hbB1K2jLW8wNJeSwrdIWw8VjVf5eIXrpCcgmJb+Dsz
qcVvFf7xMgjaZe3lBEXXlKpF7IQpcgw450ztKccUikRMyFlFcu1o5GhWKeMLbjYP
sdBAfNdOLYCZMuff6/p5t19iLZrXqlYvySO+LD8CN6LQ2rLj9/BlZcsqvTzxgd0F
enyJ/nQK6eqSXGyWrXZnnp2RSxew4Sz/Xcc+g2A67mggJdqCIk0qPf4dvDllYmYB
IVBiDB0K8kG5YmbBB9WYpVkxt5h+XJF0REp3UYqS4iu/3EnCP+n1cbmHw/VRiaeW
+enMuf+EjuYJ1r39CuBHMusjrN8u12VwMgSgVAV+MBLTUuc/+Fg4V/5sWMl6jh9V
/HqWlS3wgOqMbuoeMJH2V7/K/BqWyzK99LAvrAQJJWzJpSPnn4g4tq8LWlaXvM5z
I63de2HjK1cZmB57CPt2G4nnws2z8hbjKe8CDFX+3BFt0usyJGQDH88emcpNhXxH
ezJMqFeGSlOu/PXMmq8ww6vfSxS1ZPlcSQRvXtunsksR+dj8qyuqy5pw103I3irv
203PMQnRaIM/uusPhUotPekdUGCI3HB+bmRjGrfimTW2+t0DRc4v4xsp7KIDpIMI
ah7UKeQ40n94Pao3qie+oyA+2vLoMc2rjSe+byLfy0+85+e2FptqS+TGXXzlK0fh
XaqCTFjM3ZLyvsVVvCdfcNyFQsIaarXB45lmn7o9A/x36Pde18S9t/lTPSBBbIcl
4mOXhTaCRhxEJINxadROWTWO6UmpYbgGiXrNEvW70C/eQa8l3OSaPIW8kWHGL7v1
WZ5xtsKAN/MR1EdrDTA8+lLR0p54LpJcIMZNxAWjTvC3pL7B8Ny+sJ+xwEExmOMK
Y6PBH9EVbLpApGKWWvU0HrRF2UErwkF/8fA2ygxayuCcoBbduHpW36CMoNbXj2ze
FY8GgsXSGiRKX5W9g6ku38F9RzNr77W91owiZiHs4VFur8hYRymmsZsLN9tQyJs4
A4B7CWgQP2Ex9StifUdvSDMs9lkbqvFKF7JM8MPEXvW/ow4OhvduFmD9mL/CWFrL
h9ocXN2Ol0SoDFV/sOnIz9p+xH4c/0H33BYM+mIblJHVbL7vB3mOcf4y6ypAtY6q
8ETrL+L+P4IiI1kuy5vYIL/yZahQxyuVyCJdVaDL7pNGMZhey3kP+/1Uj9inidm0
YdhQNxUu2S3d2LYFRzpZ0zPOAYAxBwAanBvv4WcUEemtcgIicxYNdPJtLbbFi+Nt
BA9S0cKBPgJzkLOZebhZFS2WZvXicObvYdA11OBZu7Eq9QjAjx32AD6a828+S6vy
kltoofGaUA8aIlipHzC5ID/F6T4pQDtuk5ZNKHgZeZkxQbtVzII5UWHyinI15f7R
AdU1ZHc3pXkRdG0SjgcWrk6mhVWKseU0zQvfuxFv1u+jGORdeW8wRA7zMtRRlj27
mwh0C24/8geTOwa6tfSx7cTSmEJ1LbRT98ojN+1XYgUegRKXnGn3E6B3UR2nLFfM
x5dxUmcbJuf0IpGBaQIQw2tgdyY62XEC5t7waWwZjSH4fyMMIolVBUUTZ/MM1e67
ZYUL5OTRmX3FZyrNvuD5yD26sFISShS/osEtePItJDnNr+dGn7mje+0nLKxMP7DG
FVkHx2C9Bw7julaLoPD3CaSEGHTt4AgyifAycjTv9PTdwuyKVyiMsEVQZeSlh3Ly
doBGo87fSAebTuPTJC1g3uoKLKtbnaP0wR72gfJ0NTb3wD+quW5nqSqK3oVWp2Iq
li0OOcbKb2+7uhseeTxGh5mhC/xNGBYX7tKV8O0XscBU8RHXha4M+YEKzgN/Hele
EhTOOlGyTPNaU9JYXUW8p/tmSMIpzBMDjN/v1+3cMrx9lNM92b3NWX1ZjJ0tno4C
N1Dsi0uCXOgqMPuIjgVrSMAU3gSpDjZI+IJgeGPXdd96+D94pkrk2+OCG4o70Qon
DBLQ+gq1WNVQ3AbWDnRFTw4ryy0BN/8rj2cUVx5Ntdp7q79DowPEsc0jY53UQ+kw
1QUEESUfleaK4nQ8NwpZIbpKcc4M3F0RQl6S6LF1AOM3SyRPipmIZD3VFuRCSz2T
uGJKqbx+bH3czDD47yXjiO16QLx8N4Occ5im7V6T/YRMaoSML9/Q16Zjad1GEkzZ
A3Rob+o4aSVpLsjfKy8KbGWyAdVkn2+J3UyTe9fzJL8/AMn611q+IVdoNVZaOweG
ZELXgcLIwYVSuGOefGl32EIIgHgBWi8Cn8pa8b0FOTIUUec/x3i6IUQU5WxNYbJV
26bAFRDvduHjxzTogXOcoU27f6WY738PfqJ8e2KnLBj9dUrmkNaDqhiKDVx52AVW
4ECE2EgStrJsIerwTb58TbcrrgYrCcZ1aymARqI5vXwD5F8p1otCAsIKnJ++aohJ
CrpXQy/kcbFq04UcnLmgj5B0pgVHrbFvCA53RAoy71z9TCmyYP9aYghjI0veFJUW
Cmxi6+gN/UOyLN6tFmHUWn/mNOzrA/ToxopDoFlMaxXszqSRUiX54F/jNpeHeY/2
mn7+9UZ3E/i4HCustJHnO9F9d4zLfTs/MK0VXz7ArWpoS4EwLAuM/3pNb+ut79Yh
aIXtUDyi4771xi/TsO35qLp3MZRROEN83MdPz4FTvyW1SI7fhOmt8h5AXWWXqfoH
1CIHlg0i4MW0pJiOTPovSHKCxrpL7WAL5GJPXsSKQW16DZ6zLM7Bad8WB8s+DKhh
2xtzKYuX1z7ijWHqhxMZfmu05C5Jm5OpTZ35G7gWDLKuh/zrjCNuy8d0GDL0rxVP
Pgf0FgFhh8VxFMRh5fsilCY+2H7TZsLUSFlWG8d670fukhylx7HLS2mvkOYlAC6y
mBWl8HuUCAJwKfJNCUXzkj+xVL0BokqiNF02G7uQqBschptyaUK8uDaHNkVvHsTT
uZBzdbP5qUHOmQMmq6PayMYzzaArWD6u8RJi6klfyhozxOa7XgwzUikyqKHcYBCa
OyAC0q4NRIYw7PRA16iMGSO5Th6zviqO/kFT/jGd9vM99oyYMCgWXMtw8Qn/ht9D
HuP3/AMvo43+xfhe848SA+VwSgz06HFUsLNPyZWuS1DOBD48atBHcQfZMcZB2tMU
Sncd1RRblJ58ecFvLIC3fuOZIwcv7QemMyD7V8xI7Tq7MlZ46eFODgHDhF9qpDc8
9l4yTRGMKPNd3QZpruQHEelHII68OXOZMq5o7dUwBBL2xwPeGa466Gc2Npd5WShk
hpWZ15YiWh7MkbP7lrmQx23Z9GlIwSQtP60zCCL0fRmgTracrA+41V+VjYLnGhcd
1ANmdN8GBU924v3vSNskJdyaqfxKadG1OzMjBGjiZo02t03blihaKYyq44diZ+1p
5ad2CwmK1WCJZu4Fqzg2WhijPO0hV9iJFV/2P5+jIKs2An3+GtvmpvOPV1rDl8Em
fyL12Z9Cz0dFeZTo5lbkO7gpKaHC0f9yLwKccDdxitBLZwUKj6w2e5D42Z2uydyX
PvTuhUcQ4d7PDe66esDb3qXkhciPg2oawBJ0TdFLLHXr2xi44MW2rzBYjsdRwfaH
7ZJ9grFAfEYzJoAYsGD98v+VSKul88NuCHcAWBCgbicOmMV3OEx7VHzWZUIb3q2T
T8ocMJ/yvDUkyPRIxJAbwy2EqA/EQpNDM+xwQ3h5TQP5e+QkCpYAlMFD0S0vRwJk
TCBvn84ZdY8BQW5K6UmbnKg2GOwFTAv1xJW5Z1BIC1cL01nk/ae15Hba+Btg+WT7
xiKSr5/wwK94GdBGoengQ0znR9NY7K1LEbCKZR7gL6SMJeTWj++eaSiUTAqAAH5h
lRzIWYHKqYhcp2/LnzClqgUdESLueZ7A8s2cv8Eb/m+5q2alsfAH1/0uDFR0ielj
4jy3kCbuBM2cSrqMo/6vxehZ0ktPrjApiJUfN2rpX0Pc4UB1iyiNUVIUEIFVGpzq
bkn0rPDOU2A3Yj0o3DkbrXGMKgFxsEphShzJJoo2h+gGCfXkUk6fROiysXbnwn0d
QFvsmIZBCcRWDt/wmbHCX4YE0adE88O7j7m4C9HUtpnzRNLqC6N/OFNBkeYCuhIA
FmS/3owdj3vCmeufwpHo3PvEVvC/c6USURB3WCLQ9yeZPBb+qn0D0HCHqmH3z95j
YyPVLBDsUk40tFdWbM6Lsf2QIfhnIciCxHpAVO8DMU2exYNfKwZ42md5bS6Qfeop
lXPrYg50jcQJMZLa2XitLOYv6Rw8aW3Fd6XXcJbvq6BsFZjRGsvfSgCUb52Q6vHu
IY3XelpnP5shYz4Uk5hsgQ/SPIm+p3D1VmwFVCNvaqDVqXX7gwcTExzmJPIgKTVL
ukX5y0k0/gs263zV1XaZ+QFmCDrzj1W81l6Ko2UxXTFYeF2lJL/Zr9twnbNBPwmV
9xQsbmIh2PE7wyLtYbaTzAZbEAixmbPP8FMZAejTZdvVR/ICUAqvqu8S/d8dK3Mg
kmmQqwg2EHEnU9rFYtRSUGmnvjyUcVMC9sdum9N2k/3wx9PQ27LsHo2tuzMOpC6u
OYlrP+7z4RVfDXTi48SAYej2ucbjyx64fa/1flPC2PKPQ2eRO2hvuOna5Cu4fvNA
DZSGtSjROnEJMmEewBNJNtazDcWOEOHNc/SZQm084pyF/ih720hwECudxMKrn55E
idzPcY4OeURjYiRn/k2XKan4OgisAaJZPZJgTb4Wy8McZ/ii3loT9W1YMMN+Slw3
M4jkBDXyhF+HxGf12dWywlW4yb6Qi0dxy6Mvrp7OaafKp0gdvaApCNzDzSzebVYX
oGi3y5sKHPfPlvgx+VpGOGgPBes/1iVm0Yt9NfiPxifSfko0jy0zK3pVX7xSRWx2
qVRpaOq924lKCNLhhu3vFODOMJ0p7R4OCvEAf77HE3AE+gyszihUTTyYc4KCJxS7
99gHHmQ4YsTz7WAiF3VDwH8qKVlB6V+ZCi/9GCqMQCPsFvd340HZfyzdwkeviMW9
bkdZnRpXXLGSQkZJK4ciKmjgktwhzNIy8ZMJn8jWvGejGQFF0Ft65aTg7D48LfzC
94DAn94cH69xPo0XQJvepglFNMnBYEhyF/hmuG9tFrRVBDv270F9Fu2wh7mRqS5u
kRx2+9MADzl3PJTzF2Eevozynn47YcFICaGFO5lHI6QxRZLTfgGYM08qelX6jEmC
xY7pStvshYiKNaCV5Uxq5oL2HN7Malb0uJ04KbxwnaUuTqQd5MY7iIAkLsDFAbTv
j8/yfJyiBXNuAnnXZyH/11NGfjtMh3qBdXqqB6vz0YVgezSoGYf6o6ZzdzFugqpb
AH2muGhP1yIhfPci90VLOplBPHgckTrdpVJySt8FKV7m3PDncJZZL+iFtGdpPnqf
nJS3n1HecNR2a/HiYRTv8B9ZINSrfco5dsAyZ8F1z/CinKVod+v5VIDKKvFGItYA
5BaOFhVauzSY7GyYsUdvSLfRu3j61BGIo29ipJaaczLjRtxO1F7FRAccIv9lGyrI
kdQaHjVHGCpXyZojbieLnOWeJvCyeHMA1d2kqWIjItzQnrJ4J6bmj9yXow/YkDYl
0FW8ncGCaf7yc5No1pHQUmu34gDqg1v3jf0brSAeAgna0KKprWwqgT01vX+hCQIg
TnW5zQvRhS8EZoVNDj9/jKz1FmjASFxnKypzItfWPCvsn+qtEU+fGFyf2zrHydY1
bHReMciCjK4aSftmlTnUpNVOrH8JG1azcvSz2SjSfHU3HX8usNoIr9CeeHvQnTNY
FJB7h21FI8O3IYpeI42Et3zTL/bWuq4gt/yXgXKXZhhGRI6KVbuReCSd3pGMDTIi
56c5xyXbis7gjm2WPoUXbmLDVwyp6DRv3lB1PkbIe1mOAwAUDD9+8A+cqkSs6SC6
t3LnHqV5Ffarj5KIUML+eCvNH+Zl0keMjxrigPGlkFbiS/ElYpSJ+aVPJzEU5V9K
whp3CWgHRuVdQj+kszTWid9aLwEfvbVI/NNCDBR1EnWy19ligGc4VNs9BaLNSKPu
Hium6xAR00/QGAKGowD32jJT1QB/15pntBcsh0o3MI5D+FklI6f7UV0b5SguU3ay
CvAc2S4JEuCTxp7RP1JXSgQQkrsO3Uv7eLnxP73X1GSnYaDW4rI9iaQhqpkkN7lC
USZkujwG1gItaVQYZcusCIyEYesqZ2fWZDH6YClPF5DmNQD2Lx7EXaPEu9RwxBmr
ZVM8FjrhexyQxIH7qABXRPhJcX5d6e1FIChlsey7i2Tw5i0zIf20Sc8asnzh8x/O
oWbrSpAa4xBofyWQliDZRAxRxkdtudtqr1ha35VtNZayHki9e6MJutwZiLRyTqcI
mfh6+hYxO9jzfSvECU2dgD7HerxWtwbiwHo5Fb7PGzxiDS5zOmSerGaJ+d6fA6lv
7G1E1hQrJQBdvQugEiD/pF0rYtlWwZwzUvStB0I7NdJcNrjgClBph+s/d2lOXFqt
8kGjR3uwhly9wo9M4qsWGoUqtxiT/u9HoKpkBTX2fJoo4jysgO71NLIYXG5dyITf
U87Oom26gVeP6G+DmeVNNF0xQj5FopQNT+tQO55T2L73G7p8ovYQYyONPuUE+qBN
jRLelGT6RT3YgUTpdj2Gp2Po9MCKnG76khVKULCSssRAND4CF+yFMn1JBuiD3CGZ
N5ke74ZAy3YFoKHiQutab8E5vCXastA2qq/njUvzV/zgu3wgpU99JpqUTNleBacM
Val8PScfZ5E293b1+5H+iBEEVGKV9YFLhzblEmh2p2GnSIJDxVL0ZtsdODqQLf2Z
wRCLW0ge+2K9lnhf0BJDOl8BqFkWhiGp9WVuMJ8PSHsQdePSXn782aPnJhXL6HGB
E4cboRYrWUcOPooI6bnZbppQnAOkuUhwC6urY1dCXYJCJ307IK0EZnlTmczi0GJy
eZeP9YKvWJ28nlRiX8K+QGY/obQxpLirSJdwMpTbGNAFloI8PyRTJ2Gq1ckzBOJc
t63ktnh+cGgBarq5i3yJ0IoATqupc6tbht2L1V58iTVUIOEQIHGmjq5Kk2nK8TFy
iECfXmqzF1Ul4esQVqWSZv3buGY7c/D0aFvBw4NVexsjC+cSKyXvQYmJKjx+xP9i
MXrsKqrf/AU3FjsXNDMOP+Dwb6hECGve1QZGKf9KRs+tIUkeWnPcGe2TJDABbb5N
n+CcMDP8UPaiK2RrLJe/0zdrmur7dApSTBVjHuXd2gePaJSCBWOsAmiYqnUCeoN3
7bju80+3WL/ElhL+GEPq786ytHMy/yOR1DWJj0Z3lM4oR7uN184yQWQIKUF959XP
6Zr8gWti8LYSqmXdHaOFb3sI0NDHUQs/Hi1QNeeKGzlCMFRcQ/VmmTJPZqJJAB2J
KXKX67rYuNx/sZtefvIR0evOmzlP/Lg9RmDA6j+iXVk/8pfJ3rzEERW97288l0xy
bLPdGo/ku6OXpMKc3iSOLavbxz4MSbKSEMzY5l0d0Z0hpxIgfJmqduHQHmBz4W4a
iyyAbF2zJDsWO5QYJm4oRIM67wtYm+VZWkwxqCJwuOmnsj61Y4FYGdA0KAbuD3tA
W/s8c0qekF2vwNZaN/eBiqzDcC7b/nbsDyuuVFWUucPvHZ45WOuGXzYLJFEtIWil
eDwg52/t88z+pVYUaJSqkqtoro/8VaiuztkAICQmQyRZIk8oUtNdqRl9UA5fzFou
MfomJDQQ/wx9uChP8rMKpDRcOIsxd1dne67n3Ec/68zrt4JCMglFESlseqZ0WdRS
V94w1Wzo8YWz61uysQFOJ36wN2zWMCDULnyapBzEuOSWK1BoA8oEjJVPHwzzs3py
nKAVoeSjwkxuT97uQ/B5txNZP/rmla1/R0zKMewlCnFJBrK5iBFuWWgp0B2GstA4
MwkRHhd/QA+/NFRiPb9Kn4FR8MCjt55VubYqW88a9GZj3QwI8e7U6dLLXSadBztg
up4we0+N2tK4e49IYWmdAlqOA/4tVS1qAB2glJdkCvuv1JdkFjTU1BGvIfzLaPvG
dMJD1EGyhgotBwELnxbmKBUkIzTw41xL0oIxG6yCwbfXQUz2k9ZcxCu/UeIRFtUB
GSwrhazB8M+sXlGTspfx4mTOCze2eIL2PIqBFMRiEr5TCf6r38bRU+7cV3j7vj7/
+/UIQ4ZBb1UDoTNMTAuwLEx/gQXXmeMqdBf34eFNbc5uy3jEQcETYzDYr8SwSu6F
bRKyDjxQOdG7zJlxfeNr62o2vryv6HBgisiVxvipCvCXqF3eobHtnYUjmYWvNaYk
n4V2YjAsMz2gLCCBcLN2pKv/Irw4Q4JWC4W9A8OpWg7y3yC16dlvYG17/GKugL6L
76kE6bSYGbWAnKisj35NfuChpHZNcu7rII3dQVYgksEdwWbjN1kgKUriIg7rfyrO
sbvZouRFSmyaObSzb/3HoqrygPwf1Ji/R3qAt9iWujSB+bMa8EyHOHZ6x6eX59d6
hML7f2zRsh9tTqwJnojGT+na4pOcurjEXbc90537QHH2nDm061Ik33IVj5g5+r90
uwkI0IeX7BAgCQRAZ0kA8CF1M31WqV8DvyDtN3BDDzDss89tBe81xd6PWVDTyVtk
1iHwar9qAs926PSd6Pcj7KGiJSL77zdbqiEHESp2uzG9l6v+h5lyr6MlWH6odm6N
Nr8vSj5670/OXiBjo3WOpj/0j7aBqyrcimizZXTN/ADuCJE5RJPuCL4LFrd1ngsC
RWj4SWsSB4xMXIRD0mbwC2vCPZHNw2QpE13Xo74ii8S3itkW2qtraBi/cSDZUwl3
O35J7JWnq9j5FxSwO2KYw637GWAq3ie38ez+fMuqJYGetqYnkhE5FewiWsO1ofox
Iob9uH+KsraEEUa/le0Y0rLEvw/Z+W/afnNUQiGJbOPnYZqEvCM+l4Lwephp5O46
NtHIQ3YjSAiBMXv/Y4D1iTXIkL7bJPmIcIwkQolNlJ0ZVJv8xB6r0oX1r7IQQt+z
xHXTecs1DFjCPXensxrVGuDOq0DSiZhw66yDFTaPtWzEMUaEO1uCLeknTClHZLQ5
K6bcDmCzTVEw24FpaJ31mBesF4KGK4sflZ8nC3S5IZhmT2eIme/npm7lDSRPUwt0
jAX1W95+goUeiGKkTOhNWxpJJBV9NrzCTcTieEGHjrhbW9MeIf8b8hIEMNjF1jaU
lPt87qHwcF2rBIFgL9YhR8bEcHGFBMS9n5PI5bwhe7masa/Oqas2OFH8Yaw+bkGc
5CRDe+Yl/klZUQlJRnQEFENj03TdVtbMFJYVsazqy142lJGbPAMBsneq889KS0Lk
5KH/0H8Nu1U4P1g/jaEoIdc5D/0LP8AnNaENdYsKCF8Y/lycicXH+RlXUz3K9sBH
uJU6cCumPb3ZiXhSPOSywsBouyz6NleN0NlgToL2ZSE8ErL5qASndiHnZRy1l0kI
qq3cGTJHS4RF3DaVCD8LwyHu6SUdNze8tkwvDktoX0Qu2BPtNlNpC1t5/iftUmLt
+O6Narmya5VItvl91PoisxlUM7jGJ1zcSHzKvnT2PPnYz5YeS98/YSb4WSEkDb7y
w19gwyaKfSESFqzHpgxQj+85n4ckvYR9ll9cXJimv2wR8WHpAWOMAyUA+gnyvk3N
ibE7MDhzUSmA0/KJyNvdtIWsMjRQEbrMZZ8thc3TUbFQybl4I24fZjp5YWKXzvHz
jjVkpfRC5kFHaNFBXws9YujT6jjTVdqasPL7J5czx+rk9LNCXVCk1z9dzHvrU/Uo
38qzD9F18BSoDbbi6q/8Du2h/yf6krobYN8vhcpKHM34/QzrKWiGTxj+ZZvEAXp2
rA/+GclgtbDEQIPUrAcpk3w8Z5Q1JlfUBXHAnY2exIyig9w8Y3pdjT3+hPsJeFpg
4vtG7fb0dHq/h/JFxsCyPyU7l8abb1Umez6OSN/ODNhQRUM2jSk4GLjrO39r2pLY
JB1rgw06SVwebSW6YOofGmvJrSZ+jySXbZ3A+5hiBvbqugstbRyYXdtTouyZH96z
eQVlgAHNue5uhdrPwYsr05BUMdAuoghT7VbVY/qxkVMFYiV5VWy2awAOkgABiJ7J
e4bFURIGaJddqqmiYlZK8B8fNc1kBARH4fTVJMstj9tsuOcFxqjEmxssFHNENhoV
yqetfJzKXzimVT7ZA56J3sExDB8S2ZNeCEqLM8EClr0ZZ13sxH+MTkUezsDkaxAY
QhSf7sDdpbg43RgXcPipcBeKhsDM63PjwzkCQc6FcsXXDLnbd6/V63IJbK3IN0kR
NkQYL0jfwvWGlUiSIENilabFq1v6CRsbxJT5B/VE4NnVhnHOuCqk2gJt5wXS4zlk
Bcc6+DXwVjEzafoaWw2BhWpjqp/Am47DPyPJJqRFDB/gpIPDpe/p3zaDO1E7RfBd
YgEAmzhOv/NDWTzlxC5xMpDU6BS1Ey8at73b6NHWgaHq+pr3L3Ee7qwNl+SJ9b1L
2Fa2L5vK2/gKRIex85xkRklvTMCma0klfnC9o102VUUFU7Ry3LFBzFKXtnGKII4+
lF/hAQ7yCPWe/u/2NpHSb8g+t8upPKzhBkXfrFGM7elrbinc0ASUEppYh+weSLRk
fMpeKGkE6hjUstRrfE5clEk+MuBnlyluBBnmQJZBR6AQ+hWu8/otDdPFoB3bsOKv
T48dF2Q/THPV4eo2hpk6xI33wpicoWMw+t3R7Wapux76dN+vOlt5bn15ff0EzU0Q
9Xzz5zZKQwYZR+/20yOBrYz9QrqTwaV8EFKx6X9EFvFL7kGa6xZNRoJBftO4QAJu
KXliJbyDPxiQ1ysX33V6Fd8RiE4U/8Gg/4ChVqGsPqPAVhYSOk5XLwux6d0+9m7M
YXs1M3kzKEJCW8vvPg8ivKf6ttMiRVefRoUgzOnNCnVnA97lean9/zsYbmsdoQwz
LCIaYgkP1G3ijDLgrBI8Ojl/VVFLSLS46qGOiOc792BNim+XNMJTvXwyo2xmJbHG
OkrASMzF/4T6Z7MtKYoXEj8JDaWLr4HEOTI2bhkwsLE9CuML7VzjiDy+y75s3Ezk
Q3WFM/1n6vOopH1I8cGlwegVx2sswAtu+mMbkE6Uc5H+aWKWqhkMr1NmZRtbDvHm
rFWbuv2niujU4WKEeydQDIRFSKAWnQSoefJ9JsPhnZuj3uvn1f0rfnVpoAjm9SgX
KAuFcjeJZJg9mnOp4G2yvvqGFU4xfLXImuv44qsU+b/oxI3ZkSspW8KgsVRDMtZ9
nH6A37KcUisOrwPj1uiNlQ9xeaTGjms+7ZbmNevZw8BBqHxNCih3zZk2dBJ7nQCD
itDBE6A99oikUBN4LFanJSsieYkmwdQTO97AaTUzf8LsiMp5k3MdiAiUIZpNMELT
BIgR/HU8Pz+Gd0xdU0QLEfbC1Mzs99FSGTnb8FOtneJE5C7W4/uX1tVJJP0Dp9b+
oid4LwZjF+8bLW/gLSd1fUCSOQz23AcT5ccqPdUNf09ljjpP8G6vuS4nAmqQ/+YW
tJFeKFK0HtMH10G8UI5YDmJT80tsNwLijr8offk+z03hWC0b6IT6swty1JbA8Sdi
m+qGEObdj3nLCbKzGkSJVrMCNx1zt7/YiIHELCKd/7oa5b44427PqLFT3ubRzqZr
H57BErjcM0IvqvyKc6e86UrFsoVHXxRmlC1IcckmAiySLnN76G2G8rbgwVEIQqUs
mPXC6Pjm1ijaj8Ac+mqRvfV+932gTKbZN9OFfhrbJ/rkVZgCoG5k0UlHBdeafska
Pu0VO2ifumbTsLUVszCiR9gGXF+eSodWi8+B/7Fy8VSU6RMcAsaI7h8FknSl6u13
/bxl/a6mFgZwYjGN4GaUjdTQch0rqy2M601c/jFK1bzMtdhXB2N2LgjhhLmc04d+
f7a1ZU/RMUhK49i+3vFiNLJ8G1guzhO2sdPfOzyhEj664SnGblvCM7daqgfTdgko
9mx/xMzzGrmnI6oSA3NFAJB6N8NQedxxEwV87ywKNH8CUwc1l9SI3LNPxTHa7rp5
3e0lpHgZG0QK1R9nn9yPLAbc6/Zyx1TUH1ZRAqEqkBZ5tbfj+0gNdsbdJ/Ralr/v
WIZcfJhwmh68kWTXeysgNF4kjM4sejGGQeyQZChMnp4WeQvjar3LK3b/emhWvtCc
UaZnpMUl85KZXmT336vWkkc30imAI9lngaBWEC3+BWmnI0rt3mDinjUVk4EcDXzx
5wi5OA+FLJ1sMT6o8S7FfhEADXdje79kdTbpcS5s/lqk5cNBB05LTtdaPcrG1uIy
gFnbJuHAAgYbS1kfztcnhNFrqcBfI0J3QBnES4fwDzAFIUrmxQhlrbdsunaUQk1Y
26vMS+mFePVSzWMdna6P43XFgbMHndONSwu+GRi4P15gyFhr6KmtrxOluwC3SoLB
shRnx7n46IjXnQw5m28IGjGOaG/521f14UirRIPOgrLkHfhsN/+uwKm28eMlmuvZ
p45/aUQYifre3kFgwm/s10wA75e9e5+2arCnyUDLDJryUqKLXVkZhvG77Vz1bpmW
r9rCpSBbIDUKBWIY0U1bSpAtfTsq2dB2YE8Hejew6cYBHMha8P23tHXHSAt/x13T
VTagQuEcYRgzhO3XWdQLFii21j/6ZYZnKaWEdzg1A+TnfbA9I3sBLeciOgiI45fM
ECNbVM5cvT99stj6Ko/ODxYjvV3MHAoHaRjwiHNAKlkbfHb3in4V+BMQ7TPwrAtO
y5ZxspG3xb671FwdSP870Kl4wcoB08xwFoetK+yRReexM+TUjMSXW9sRgtKaWS+d
NUCTZ+KodRDdVMja60rKqSpZog6hkPfuhiXa9G5IwP4LwDKrdL7aW+9+JNtYeUDC
ytBbujSi2lmvHGaNK8d5hbBLm1MiauVF+RxxEUKY1+k3K4qa82CAG4BaykNlgem/
SeqB0h0+/smG2T0q1w7SK7PuymG+nnLeJzE+VEWw5zgRj3Z6yoiU4HO3sqFuMua0
5/GrGz+QI4AT9jmMW2XMXM9ym1+q7LUR8bTqbUDA12RBKKVyb3+XTS33j55Z1D2r
izx+kdFhkbjBJOVN/w1EtCfc/j8Us/j5nSXWoa+2Uc6n4qUQyNcy+k4QkddNDE98
27X2S10ABDChuUsF6BP1RbaeVfowd2kou68GkTfXlN23PWt9Fdi0p4qMHgaOoKNf
umdeoXQ3MYfTEIRLWavLQEr1Ekpm8+T0hwooOqG82kJUy7LmRqMM3Wh8nYJyHxu1
etchOqPa/KcdnmzctIaJvSU/MvtDSLuMGoysgKg1iAdK0/XR3mlaPM732BWit/Fo
sQBOUpXgXHKwKZ2gmzgGKfNGhJkhsSTCZEq2eMbpeNj1aYbvNtTfaqE6c+hNrQdm
OltqDbPGN4xCTHL1ArTZlCtHJNB6U2XdGApM9MsFjvDGsjtkTaaF3CGiBA67ELLc
K4D4zjWHuf5cuKUz6rkclxiiM1SgwCl9XfNpCcpJASJZogMUzZyOa1eEPIxgMh2T
AfXLU8vX1S2dqUNRosvXhSNJjZYiz+kEvwwJUgrjcvSYVEcf7CcPQoJKTd08EYf/
O7F369oF21uYmx3dN2lXVNWRu5PjUxB+q4pav1LoU5CI8QnH9/vErf9+a8ATC/pj
flPgh8OQpjnpWi5pj083K9IZWESFb6/nNkl+Nfpd1JoqClvc8lzh1ATqT07or12R
GNz6U5OO6fD9zDxqgZWqlj9C85Aji4UudmEe+QEBjI/LlsB42obd5oB11oRex+em
jqctf16JSC4Lv/XLvsPsaEo5B9Ibwhiq9KqTBuwDpPCRzh4F3RAZiYPfuHgystkG
64bit0lXPwjHVu6ovG5mM1pReQAF2xBsAPVrKSlmeeZvnumygoTpoTWcHIxTtEMX
kaQZkNaQ9PBdYv9DRq5cUfF24VD7Ouj3xcQyDwZS6VwG+z7XCt3kel0Wbubn5jNg
yKdABn2uj0gDuxOzMYz2hEJRSEKcb44JKnNL7fARH6WqO9GGBKGzvuBP24iOcU/5
DWJkvLfQ7+NIOCH9mGaYRlfOGyEG8izwMhVjbyXD6EFuoi/zJGsYK+Q82LZSdnDu
kmw40BUYAjAwm06XZWoxnDN6XyVXmkRqOmhxX2XD/k4C049YX5Rd4RHIZo5pRgrC
/HmQxBRaAfAentIpgptc3ofEjFtiLr17lghRYinDi/UmqhJD+Q2kSEmUoB7RnosO
9u9Kako3Ukg6109QYRmo1cBfbJZ7TzH0csD3ASzjlsg2JXK02Vm57qfJTNidft+2
TqgreT20lpMkYTKIlHwjmAq//uAU5KUY5fKxX/ae/W2D6eZTvZA8xp9mbW7mpUgH
JCZ7cKfyHsVeKFKa+Em/9RHSFYi3+kxqOpaC90hF/hCRxXaW5XMg2wrQY1sKWqtc
VPhwhyVxuXvjOz2Zv8Wk3aeyviJD6sgQ3D5MI/dy7dUFGelsZvsNo4YwUZl1p6U2
y/MIfqqLlVDvMwk2zK7Ku8SWdB5JigY/NDy5kxCZLXNxpAIhP0/juyXVHWzrkYI6
N5KF8s6RII6Z2JWUBCSdDJpV5YPsofTT7ppgA2jNjvQ6ahZVaaBmDuLc5YQZj5VB
SSKP+uGwQCq3htwjkT1vGEaUeaj6o82x/VvLQUeo+GLEeQ1b9K/+LeLLOs1NmdNk
56ZL8oqyu5T07uDN9KxMRnTBMxBvCIttFCQfGzMq38QWSiPMUMiiuq6mLbrNLhzh
7bFTENgj3HFxTNlH9Xfh011qKx3WEMNSkhP3qvPwlI3AEcNrndG8banQ8QyxXO6Z
C5ZlHwybNt9DklXPeF7S5k/fFrPg1C97NB2EphPthvxWWzw9NWAy8dER2rd7E8yD
cinqCNsydW00+nakbMyyreMjqhhW0zMmx5mJo/9B4R25XXNLJtT6HoiCNhK49poP
kIjXK2HC358U+ZVQ3HVwK8hCLpaKfsa23+c1s5W5PSnlu9wrVZugvbu4yHvXyhFC
TbHye6rHZDCL47J51LHqAFIWurmi43yOZsS++IJrCfRSVJaaA89oTAHphoFcjGqC
udu+w6nFQHXgeRlDFyBOoKtIuyVYsQbk3kEr7ua1lcX2P2LqNM6oEcmJLNCvOfZg
Sye29Jk89sKbX8jFKKRVQzsHD+WnkH+GPWZoyjNvDz4KocGpKTVUHUzpc6ZlYUtm
BNCeRxWxFlo1C+/Tpp0C3/u0jHovxzYk2VyCw8YBnhcAodm9mXzJyxMu3YzzMN94
9Y47pOV0or/sCXKLxvYciMoe/ZpObrSLGiO3lEYwifJHlqeTVJyHM09XexGdU8ya
nO4cIjB5dBmznc3zLfiRWrKJjLaWS0/DeZmRVuHYiSw24si1ureaylCMAKFKTrGW
eVYv6pdQayy6cy4b7RiZCI8NPlhaguzI7hP0JyBwBe6FSxlqiCHDkViiQwS3afTf
pO2AaQm4WyxMiPnuiKcF3161mSmUGAopyj6Hm8wdd28nVHW4ulZ2XVQX4D/WV9F2
SveX/qdkgUnAsVu+GRkJSpEpdqdIjSl7fiCiXAOh7JSoBPOYQgpvcZ7euhvWnuln
UuM3Yl0UF1/HqCdSGRQm3w4UHKkBJlfiXkmwfwaUoDy2jG7sxNha5zxfGjaoTLP/
ykxiuRbXW2ExoswYil2Fm25BdLnwVnnAvI6O05PZig/SOC9fgRLaFVylpkcUrO/K
S+h4BJx+5P36HRpSAGcE6/AV29qHVYHyqQQw+lQyt0F/29Lo0od3UUPs0krk8biX
RG+4cdilc0HZQcRucgJu/gvkbD9ALj5gewY2kfJ8+JiFgXAZa4n9U4cfPgOWpgeM
gg6CA+1dYkOJPI2zBnrDjbjd0LyHgw65VfMCC5cN3RYJy25AjphFu4YLzn8qC+ap
g0dzkDULJKzoLG2AAZFtCyigTyzEAjB3pXR5iBbFz+aUOv6/R9Y1ztpQ7lD9h7zz
6+bw6KTfr3lFJDvFrj9jkDF3OlWbcAdSEsVs7QxdxKgktNnfGhk5fmGNhjgPBlXV
hxuNr1cXmjpPs+KSvH209vxC2q8lhl2FwLN76T1UmsfYOeHHeUKWcJpN6eYeKGlN
8rP84g0EThQquTsQN9cx73yGj6QEF3lBEA0NLU22g8z86kcDeOQcQRtyeUSTnIgB
2n28MgsSwkM3+yysEBMuOmDbcrkEDBnDv2cx+2w+B/cAwiSrtsIlnCcT2wylnPTA
VHW8YnQE2BP22myAEN4GToPmYRsV3X/B8ws8YqCsQltD9SKTDPvtDhEHGoykzzd0
WMSixwbB//+KJiOLrJhPgDtJ14R1SMPwWwqRshhkFfKNG2NX9VM+1dvyuROPeOio
1qtxMvhiGfiLaKaSXneVk2LbzsItA2WKQgd9XoYKLcfVoOLmFjg/KhvlNRkrxr8L
npUDPe03nSgxogU8GCv6b2bZdY9YrCK96+2euIQCXs/ADROhHuK57oRrlef0Tb4V
tDhh9WdwbR0yYHaQ7OR9boIPn0QQte+NN+G9Nd9MsK0qITzxpJOD0OXeanLsHiVA
MGyTurTKTA9Dn4OJarEZWuJJmSxtUgNbzIxKtOPgb69htIH+RX0p6wN/QcTPVPw3
BI3Suuj6zobFnPeMAWO2eaLa9npDXv1KNTuPNsMozQT9VSHolY11VEiipFD6FNhq
cNN+h7ejQ4llTzqH6v/XC2O6aOwWJrg8gWIGX/l1O05tjAGVQMakxPcKbfoibM5Y
QBUCK5R5p2aeCFdvVj0csKqG8RNDql+o3eXXHXF/zrdA3Tj4+fAIgVON6WNCh2JZ
J8fl6GKTgtLkObVdm2bA/IZCodsKjxs9MejuCBxxfr+2zANeqfPXLV1wucB1h40+
948Nc/uRKjEsX5kcXHjVVlIeLhZFa9iPjV+nFcfcy2PNFOMML9oKSgUZqSyxSo8I
fYyNqn2iDCJYr9uwgTIGUGlUxJ8y+Fy1zNt4CjB4rV4zFgfqHLNXfbV3Ny4wDcqT
/PvMYaAogE5k/k0NaybZ6xeLdIY8aofbIC99Kv1k4JNiipH2jc7k7j5GFzkkKfoe
CRIDELDcgtG8Ru/peridxcokU6s0Ui8F7EwdnXUoHUnCO2O42Hp9R0JS6sH8f5a8
j/7Qs3KLvFlH3RFofoKFGD0IFLiWktMH/0MRIZEiLF1dpbTDRJ6hlKE5ZIv9sqp9
ncRJh8Wtfgz6r6U2t8Y9+Rl9gNcp0BUFtOwKIkaEMjFtbRYzY/N68Ve/8T3sLHw/
HraX3JzsF//QBCBWRjXfFv3MkiQMSW7eoYWCs2wZF4nrnf/eb9mLXlak36xicRbS
PDEXHexVYfy0boV/fvURqMUbCkt2Zo0kqWAL9XUmYv2RzLtSFyy+Zqy18kVUBRBh
OUMqE5fHZ386ue9pufwZVC1oT4Calj6+gRJT1XNHtWgbOfZD/65c1vxI9J5d0TL6
7IVISXscFEOpgGon7KAQAocgfrfKKs8Z3u8MSK4WpIRNKVzD8GefvLZZATuGDZ2A
x8PHcaLWdJCW/SQiJd6i9lMOOY9q4Ki3EaOsXiemcDYupzAYSz/Y5hinna7K4sZS
YlcdwQ7pTKE2K0AIZZCcPwDdmjLvOpHzrxKxgL3EnhXn9eSPoxzhgKZ2Aqcj/bSo
B6Cd0ke5omgjsOp4BDWXdCWNTovXyILXfc3eNVxEOQZXff+YkjXXyvLn4+cRUi+q
GbMrkSQ1mhtgHXkfQhAwj7eu7sukNmq0SVhOU4amau9E5SZNFFehhvMBGSP3/rR5
KvF8WMEgS0YHlYpfReStO2+Dt6+snufVwWEQ6yilFDtX+VGQPGUesoUKNMEy+Xic
DEDKudohLC1UjnG33PwSaE0Gs1Dyf9bRxKZ8Rr3EKDDt+o6OpZYY172TpNkKnUB3
P4Q5J2Paa1S04gF8vy6HoNE5j3I5Jf70UpiaGV06DMRX03GB7/MOCbOmj8Olwgog
PddtMgjRRom/sNHC8Lr1Oa6DPM4CRbrVKcMzHMTbEjDu7cgVngLjOR8X2IqCIkI2
cFye5txeyhlw9fFIyOTRdKsRU2W2ZpDIVqjXxr9isBrfOOmyebv6nxVqfEv/Vy1e
0wGZy8jA9uo2h3+JBbuoS0LuLN5G/HZg3kDYpq+2OQ/8srkMxwwTG5R4ihZcTIuN
7uKXwGA+Eg3mjSbQD2fWbkZ9yT2x2VwhdNO6lemmA+v8vrp68jay4pxNgBBXh4bp
9VYvf5tJVV04C9abb9G1pX9SMwhXeclbTTrH2aV1eg2EQP0EuReJjNNAMOwioEuc
KradGFsfzRMSQSh8tTZi+GEDMDwj3EmIoMEz6ynIovd0uejee9AsvR3KrnlhU4Fj
TgmycZIVakuRH8U96zZ6nBH0c9e/WL84bL79GiyUeJZYpj6BA1Zp0A8kJi6SPES0
xIKp5F0bwe2iCabNm8h+wNEkqQYi+bbFGORveYPFlzHfVQkpFBH874c7ga24v/8s
HWmdXFpKDCRj/yjcegdxxpNXNc+J+RobS8+OFR2k+SanmhSmv37nAvSGer8zNqhe
AbxDv8Zt6MGKlFBKWAdEiy9lTDVt1Lua1WcWXkGItMCmTLv/KzkzPDfkbIdfbQ5j
BsW0IcJ9OJO1DaKT5F4kBvj8wK+ivfJnOROeVturEtZnxwcAZOt43uy6j5+L+oFH
qXJ0KTzP4nYIUcc3em+n9my76ptr6wKakQdhh2Oq5lasyBBGcD/gAQhHpbvnA4NV
KBjrXWKTzDBzar2o+Td8tz6TMU7QI2jG+AbhKClCdub0LvHuGePmVY2QfkB7nqEW
/7A141UYtglR5t/2xemQIy9pFTzUCNEt66xL/q60mlxN5rfwuSr59CJcTJkD+2LF
IdOOWhH+XECvh2M2SKc+Q+XEyCbE4bwlBurBLcL+4CYWNhLf7RguwWAb0m8TMg3g
R9UZx+n80whWamZYvBZm/E2x5jvPMUxwQh7EBR012Y9YmIOpnBiDa1JoB7rpxJ1S
BUGlBLnKOvXtp873dGx8KrOVcjH1oBkRYJ5UwRpKZ6WrUnzl0bL1S/7YAhwSsUCT
jNvzgnswOdSIXrK4yS0qS2xYooyE0Gi4X8wYX/A2MUcEVoJkjHSTpFld9jwRHEZ0
owqqOTwdMaFPgIHJQvp5nRIhfmEV38/c+jDfGdlLcrVulqfQTEXcwEO7Nb/Q9MFN
1u3lB/86jhVT0E3YKDKYvczYbua8HXIrSndrxknxCvC0Fbk8AdNHSLP5m/LdkSPu
u8flOFNKN9LvOn0HfeQMeCi7m9dnt5RcLksQ+UDWUJiXvxVwIQJbG3/jlEbCMRII
OXAYgdHTKnV37SrH7TWB5JZsF/x5hgZiyqsrSClbxLiNlhzIgulEmyxRnwz/bOLW
8L1f+A3w7NgU4PguA6jI1iyN6MGOEg7YPM7ApPp/KcXJ9wLScuNyzdtw7LNV81yv
4OjgpngMutw+Arev2RGzG2yRJWOeJd1kA17pW7YcOLLQLyyNY9RyT8EpFtgnyLmg
Zs4nQOpfdjh0DrQIKizRN5HbTTAg+R1nP9od8oA5nkAZUbCaCaIen0GbskzLwYJN
9JhlTant1VbX9xLKYPeoPFIkYygxKbBid/xj37y3JYuW5EAHd9xWueXZRqJSiTkI
hFa6oe6kpCWEsjZVSlJ6q7q7EiSLSHZmrCDVGP6bobNDQ8PSC2WRCAINmgB6u4bz
TplZcuSeTF868XSd4FCsyjlLV6cm7ePCWpTGrVdTKIRPCWejLpezfFFsXQVNJjrd
GX+pGexwRnxBqIxB9/zMJEjPJ58ab8X+6KmEVswHY/osMYngu1HNtk/QNAwlmy6C
CSV+sDzSoyXmgascQkkDw8JKi6tqfxHSEf3SashVzujDR0BT0d4a6ArUd81EBcxx
hRceOeRt62NXxJCF9wEdAlkRJCIF1pGRV1AydHoazEAgTKQR1sWDePAfauzaxEaP
rpAZngqoscjSrZ9jAJhpN4kuaPuIH9+lNqEytbXHk8AI+CPkAWt1x0dQlE8Vb0Pt
FEHCogqCQmq8QoqkPj76bYzzDs78nWmH4gLmgvBspo6yTqA2VmJS0K3Pjv57/MNg
WhJDPfwnLdMwsvIyZURFlsZOiUM1NSYd/CLy27APBVuHv6LwADAXCedau1kejxNM
bqvzRaWDYDAiG1KE9js23opJ1ajE5WlG0ipeir+yObfS90xfn2amxb58EJIw1s8l
uOzwc2EZRQw+mbgW9N3ATJjy1JLsuOBUsdh38vL26q/pbzE0bFxgq85zuRnDA4tQ
VMaY3XXbXjg1Paj7GibUi6ubOauxIjKr6rOkuUFmpE1OF6+LJ4We2GWN15Tr5RQe
e6pjOUTkQdafmB/p6FrEbR3H2/GhFMYgpDEPLjpY/aoxQeLhno/fkUEHOKE3a6/l
5HSeQvDdgItqbF39uOTbHQZAS1kn30SW4Dyq2SJpU/O4bfC6ynk1aRxWilHnLJNP
jVXo/WMcJCJkqr/3omRyDi1L2u3ijUFf5iw9ekOd6Vyf7MRVoLxwtUPZJHmiX0EH
9dP3d7irOS2TuMoJW6poCMyfwGKajNsFh8SqbGmpIRmcXbr1A291x2Xox5bDOmCs
T/y/Z+CYtBOT0YlpxwgL8qHprlOuO+7QoWuAAyEx0TV6/9G6OYgcnXXsRTWmscGN
NmYddf7ZVLhlGmIEN/G9rh1Ib3ID1pelglBfoQCXAAJJx9qZ72koUHhnpBwp4EZ6
YwRA3NVB1dVst4iVw7h8jHw5DUoUZ7j06qCHQnMnDrKs3A3eyTysEbMa+fW/X8/4
F+8/dT0/wE5Ij5MjtfwLsT/XmHrLJGCfFeguPfX+yLMdJFXXJUSF7Risy4GAZ8Hw
hkOql8Fy4RYb8HPpectKzk32rSTdkIr8JQxSAo/VhdzE1oO7q9F+TiMja8ymi4Po
zsFFIqrcSlfSKUo9u8pc2G90M+Hc+7RN/+uBDY9V4XTse+lBBvIqFj4Aj9lzoP4+
vQhSwVqNQ8m7wNW+9M0Y6KcWCaWcFW/aIGTmf6Eyll1XvYyRNg5Zakp97i0RTt0Z
Zl+znXZNLf2E3Oi9C4Z0bHtm9GLAwbg3bDEh7W1c5XkmB1RsveIZo6cj76kWEyua
hSsouEW1f2ZhYjL2WN/FHC5hUno2LHR5HsetqvIIF6JdY+W7XUXxDs++TzVf2c0Q
AAKQRbHCK8CUCUApAJQhikFbjx7S3ZNa6P5f6LLB8xqf29nbNQVwGrKaGnGHdUPc
P0evEa16bGUqfn8qKctSmCP1bLWw+fGOfQikkDFxT28zeugukWRg4RFu0KyfJ8/M
Q14Q/C8KYTTG6QAfFfdGPwDv0IbQ6xq6w/aybEn6SWgCcxKtGDkaSv78XaKeglS0
wx0oGMqoHeTRwU+2yJAe5dYSYBpsiPIZrGMIv4XhRF6LDsporsjSgUEWRu8LiURf
PGeX8gsD7c/1Yz9L4clTcIv9hLW9YB+KK2KPObgLrMN+iEbg4NK6inLYoOOrCpD5
4iVhqxduRraD1u4edvPstc+XlUCXOB8z1i/qGP2/TdufcqcN/5muq4PmcTJ93Y8l
QR9TEHDgCDOR67aN0CEjdygWyFlhbo7vmttbfq3uuNLS3X3UDOy6uzsEuvaIip2J
1ume6RYdEkpXfumLkqzSMq+hJsQgXjPJ1hLwspZo4hE4CzJeD+YlzBrwn6n+/rlh
FPkglInCjxpmRmN22KnNB7z5D49SP8XxQg2dNurwNFBQhOH5syaUGuI6VJnlkRiO
ZUhLGqDMi4478aEMLT8HRGi5NNS2s6qzg7tzcjG9w2JGaIC8dB/R4q4L+z3obyAz
VwNSbPEBZ70cHYfDRcQiEg8zSzi3iuzqPy1DoaehHDqGLkQszt+1BI12tptXiiYY
d8tuzlgHaFJmjOakyqfh1G+cqCY9LfcP9+WoLwwAHe5BZZdPeAMpOMxIRmBgYMSk
O0DrF0x7VdKX+9KHFhXgmnnCGpLiKHVpVoOZqQBxhMBAp3vafHmKnrVeSBDMPNI1
EkphGIsSilXxRH0+jNAvqW35iVyT66aysoDL2SwQa1bIfsjodUUIua2bL2ywDfxT
eQFboCeRvBY8wwxpAjzE6mY0ZjN+4KXeoQ5iH4nyNYJPEJuvVGVOYaWhwi69F9Nu
jtm0eG7fKiEamA6lAnjHGnA6ye7DKMnIRC6zAf1WFY0zdw1OoukxaZA5rMSzoHMV
+bZnHZ1gN4nYzye4v0R8oVY510HpwIEChCJDyEABdG5Ib5uFjwPgd7cxTUhH72yN
R3VwB06rd+lW6OilA7eDc38Xp0agffm+00DVMBgK5lN701KyEzyIakKsOh5BtqZ/
HK4pKigww+IXIQntrnVlDQaPYEHH5863BQ0fUclSFE74zP+rJ9L8WJ0//rqSLBs9
urpnhtJQOFC+UlPsq4/qiFlSRPve97XhaqucLPpT38Xjx0Xrki5kxfnhppUXbsrn
iCtCBTLy6nwPxQEBTe9VKg1ZLY1d538cufx7fwUubTY5q6URvUXtEiWbfpimF7uw
Tkjtv3fSnPv9xsXAsN+YSntwe07I2EU+4pP82iJQCF5jPUSplI/vNtrwMC3MXwjF
oWEr8W0a1hPDX2tSsgoxzFHMr5LuvFermFABdYXgKTCRArsX7h+v5k65t2qakAdV
HPZINlYBg7etLQqIiWxcJ77gRc1tTs4TRurTYKI8S7C8TzPkXAL+yq5vBTe+Mi8B
Rm11u47dbVnzKMyUj1WegxYcXU2gJXV5dzn1lg4sA3F9L39MmAIB2yMSjj2SAhW+
N+TuK1QTaQbCYap71hXbC66TtZFzmE6K4lNM/hRRBRcFPdt5YtO3phYe9UtFWItA
Qi6jCisI5d4dkjnFjxRjsydU56Orhi3CuLLvlFKzFuVoNDX7YllsM5/XgwbU4tIm
fT/h71GidRn9iq1ViPTjWWhVUoVgotD7Un5wlZf5N74YM0W+Xe96HYULH86bxlNr
Yxlr2GvERCCj+Bp2Ae4ch3BdqDXXq7rJo9UIsEOomlsXb4ooYrkc0Ftdvan2SY+B
WO++kTNxHMpjFvmgkGH31P8H0Ed+utnYgr1E8hNR0JhxDpIxB0Q2oxC8e9xWOF8h
rwHZp69Jg4usDJ0HI494x17JkyLDUmSu7Hfn7I+sHUdrM9MnfVlm0QyiC81/nctR
lmk6QXO86EJuVtL/w96oDStiU4bESq+Mn1diDoffgjmgD1DhfoUJBL3rcFyNVV0p
TfugsVqvGNtJ0eGEwGnZIWpzGp2rwqR3aEVip8mkxDgnZCg4HwYQLNfY1INMItD2
Ps/ugmMtqiUIBZT/4/za9UciOk58sN5rP5nUk6xyRe5mDNIK5gw9aB0/hq0qIFlj
rToVtgvWANeMW+vLieZhrpdfQgo2+jtg3Bi7iK7FArwWPZ7Na7eWxKastVF5i4K1
3PTkoCc8weHIBdQqAlEu0rLpie74NCAQCYykBFI5VfThTDnbQgpeTUKkbhew4onK
MRLxOAzc+nbMHdmPHEsqsv4YxggGPm6J+nZ57JYWSoZAnSBDGNZYNxYyJJ1F19Ay
06lWgqXSeogLYMT+o/DmYN/dgDsmAOhTAUqeYMkkHyz1wve6aPsaYGfKN01yTpae
32GXvQkatHI9opsNbpeAKkY9tcnQHevUB3eSPQQgmBD1AN2iPwMjnkgU66wRhEQD
DD5B/ujk5jPNFkw5s3MLlXTjSBvadqHI3HITM85KvLaYsuLiwM1p+UcaWjAF1ZxE
dh3gv4Zq2aTgqInAWKcuv/lhaQgahd3I40pZ//IuKlf6HLiUSLOS8dyUnQjzsDFk
IrP/vMRDF8P0af/LNY7G6BlRQz6CML3zo9Tc9nTvwFdwx/U8ojJu0oSX3yUCK2xn
QBVX1XAnmpb1J7k3XyEpfvN0IpROmlCMPiyZYthaPWSUrnYog/lLS+Qr97Du9z6s
omPe1u9wJ8wuqdzSgvW+CKH9x1H8ghaQlchUWnm630hIyZ8w2t4QmAB8uRzNbcLd
trCVcO+Yyk1+GO87OJEUFyfy3KAO6oI692/hrbySMsSl3iG37czgZKHkAG/qEoAr
KJRs+yc/u8ayqjfT4QC7TyxjU7+fPipwz28lQlOMkouSoNngEftOfqtyavzXUNXy
fopTltXwVYc45vYmMqe2xE8yz7Ov8SoevahOlS4510W5DzgZAwR4rdC3E+oDWF2t
NWSJUER+Y9bH6EVKy0qfq8U/vrCJq2b33hlUO7XaT+ZmNilt4/DND5WfbQfm2dkP
bfMQgOCajwoxcbqmGVzPAds+v9a/puioCerHY106r8feeR25M8JALNpbPUpCVXCE
opO5u0Yu4GO/9/wFVG7mO+A9KoxEUuCJiDk1A5JfQ02PoMieHesPiCVASAeSi8PX
akmPg6UsJCGiJ1UtwqbNDylcZnttgfUUYEMOwauUIkK2XSN+4ThkCHt18SgnhgFQ
dA9LKcNs1mvHsF+Ck8vvvDkUzRvDQsGxTduOqxwQfLWCDTExuqzhkEQ2SzKbba8i
2u6F/BZINXeImSpdjliY6Vl2wP27cJOt99aENF4+8+VjNRkvHUApDtoNnNOeWj0Y
kjjiZWqoZ/jvz81KnMKxs4GJnpgOUH0KETdtWau3pce9l+wSb0ZH240qoznZTdL2
yknJyul1VZMGE8HrDpcJeyddz5mgTG7aeijE4NZKui6r1YbLgGMahcNVXYRZx5w3
otLCAU8YWJU8YYw/57zqOxkCS+iSEpma1LnzoMikdl7E/s8lu1YT2zUHT+BwtfjM
cmZhUI/GgLKLmtkhVIEGEiDVo16rE5uY5g2TWVZOWsfhVJCOwL86PHjA5XJLDUL+
Okus+8xKFTJgY4LRjM/0jVFQxDYmdEM/oEId8l8JhegT+ZtlmcC+YveIvLEIPtjH
ULrQs2YA2azQfdR8hyKOJSB6N004PnKHgUT5T4hZTRIEzKGO/IxxJaHlCcw+p3ub
LW5U2SWJGsn0bCZ85QA0cTvKXBl3/bYCY4zHor/nLTH+dnFs2kAlILCNJNfqf4v6
qmqWjP7kFOtCXtbc/Nxy1b9zPjM7GRWRk3/uP8pG2wm1+FWnpplifsKPZxzZP/iU
ZMwIshwywRwn8q+lGW/tbmFkWBipoKDSOSR1XDt9UFcyUmOTYYIH+2SWfYXh05Yv
QNvvQfMx0WUdmAvMMjzhF7cvNzZ6GN2zKV8kPfYSecxvGts65LVwZ6F0QU56a4gU
1ZUr38CVCgnAqKtAUvofsvTSdwtWO16facH4KSSofk7rWFKm8PV1hsIJM3cUo+xX
jNUVASAaq474unIAirQug3Lod4hraTmlRNbB91dL6ZGQ+DgtCGfrqEYgXb7Tl1Zk
RUDSFDtPbgJ2y5Cf0cwy5KPw4fbUeYq69Mk9tXM1lVcAkjX6qqj93aam1h7KYDkD
D/aq799FTlF2z0HRhI8IYIrm2H/TDqYodhFTNDsGuZAcoJpBhveh7Bf/ONVIZ2Ch
SWEhg4etocjZTl99ADsAVsIxJnaSmJxnKEzGeWbu45L4TPD1uDLwRdOuhdgWg45g
FKmNyTDOwo/bnqx907lQtm/comuNvu05eY7+Qzh6NqQj5icMf1c4owB1cS/To+ih
XhyVwgiutnEa4oVbrQ8Jcs+c7XJuZ6yDOPxZWbKGl3PxJJX9uyol8xR3TwFuHlER
YBLg3lB6p0igDTgAF1wmK4zU5esSbe7lvZBklSzaQZ1yNk4rd9ZgJ47GUvTTSju1
yEtkmVlfh+/+Qw9W6JHo4QBCbpTPfKNt2+o/f4J+7SMnYLkescLUkin9nA0eqZrG
WJ2Xs6Razzj9/PbA+VRPsd59LcPuRYjeBqOpgMcfVJeR/hURpAcqfEsuiTSmd2U5
qbqDf5DXJJHp38P/fnwp1udWf7bYjuJ0GJik0LN36jm1QslDL/T0eMeqUkPPh6sX
ycomsTVky/R+fCSIEKwSqZTuCRTKK0VG/ZdB5HR1xmFvQHiXkKplDQtf3/iEChVY
tFlpGJ2YjXf9D0ESG3TwZxmQhaEDw/dmKkrpODf8zDqCLwFwCudzpWhsOFsI3mti
khHaYC+hoZCKWfJaX2hhQAHz6vJCIYrJkOdBcEXTkF41fItR3zm8oyyZrR4TaObU
QLZ2uFJGo1uI2A4WMyzUBQVbZeVqjdFDkBY1mTyl4d9M80NpkeYdn8hMXZ0zderY
Myrh9/v/cL2qNxzf9+K2jjsKg+ucVDRFppr3b9DeiGRCmvt1ZwkuPkQjanuTo8t6
Cl1RXkVi2SGR3d490YmzXKRg/nD9rtya+1iYthAvHKQhbx3eLzmE9MSRTM3zZB4C
x9D2NtKVXw5+G2qXkZL8KISIq0F6/8zZpqgV3Po1RMAxR7XcMhyYb88byjidyAD6
wOGGNS0JgnI7iNUedNInrdYowwLl/889Vb2PbFt2HLBkHeIEgbrUY8rvuw80csxH
v6P60zbveLtTbpXobkZamCULv+T+k+Cc0lGFqE5oOKZtYTOGsi0Fw1xJtk0dt+f5
PlJCEZCekNunF+M+jpOsINADM+QoJfnZv2+2gHSeuUf6zDTfW1te3E1YHYWkx33t
mOX3XB5NxPWZ+48+XTDnY1qwckTrzg9N7URWIT3giBUTkJZgAhvio8yjD4MEO8zh
lc3WM5LbVSthkDsDPtJAno6jG1F1VXlMojKtg5ewqi42EoAnmFB2FeAXWlqIyW5O
XztuSMGh2eOa82UIth5T6Aj8bzNN6KiCdCnqy1aq8ncuLCesMQKP9QkQ/Efale6y
Hs2lOKpE0r0lueNt6Ksg34CrxRsvTHSWJ/XjvCSQZKhSp1Za1vwXBatWh+aay7yY
aOUApSBaa89NeVsl/DuITTLxV8GCRtnZMsIGUNMRuLOA7TqK1L2qaneeJrJw7Dkr
QIo962Itrm5gHTucLXe4K5OJ0fJxZrfyFiA48/Bh9PL9uoZdvo0rUqISncZJ08rn
zTORUhFHg5nrnhtOVT9/8z8wUtl99V7mHerHUrNjoxQRv8yaA0CBCGaHy+Hh8c9I
xRpawrfoTAqIxO064JZVrlmCVwU5WrmU9Xug7CIgusOmFIS96TqrlOz6c7pGkRLC
Bfv4HUz7ypaecNivz5N1pqvkY2uWkstoHuhdz4F4ufxmSsDnUDOnAfoJAWm8xFxZ
kib8z8GFaiTVZlr8xeyozMzkkCz9LERGXJiP3rByepWAk71FqtYElzYYaf6XR96k
fTi7fmcYDzXgc20C+rsIT5sPBgZuWMewR4ANGKjAKiBZLUMwJK+9sYh80Nx2EWDA
y5KpL18WkhJPqKhgyyn93Y87j0foUPp60+3r7ZZvH6hAg7HxcvPWsYxP0yj93dtd
7Z2c1apUkWt0rfBlTiJ9kP+rK6WP5yjnANLWOOufezfMwV4FgVBhYD0StFE064o/
7B1e4okV0qhKZ55gMfw9FbvsBQ4NmpS1WtiNE1vhJTuZMA93zh7Q9lK+LYqdiizj
9zay48ne+ob81rTz0g+lVTIoi+SvIMglLtYh5+k6hKLvh7AorjKjLpeOhCygiWrQ
wSzju9/r3cBCsd5rmwteEUzDUF1rZEAPdLVvUT4XmP0MzH1JaloUyDH2ky9hOGJL
YPerOCAT0yW7F9FFiVExsahFTtC+7X8N5i4/ogPG3BMYr14Z+9ffm/7TKbglIJGu
6Si06I7Asu/PyqIuRzaZwa88/1Iia+41k+FHQZoGDxsa9NIOp06iN66RJTaDS0Mf
3gtr8/y1QUOEXydH846AuRpM6CS/xYUsZcDMk3j0/QlbgUkIi6sPdr/AdLCjmqN/
pQ2innrupOfSTWTxP/ZqAcPl1KTKqjETYa8y5gktUzdrYfjbnlgKrlTweNjhAiRe
LG3Z4EJJXYAfJYdY7WmtJ8Tjvyg+Uq9/VYg6XVjFHXDo4oVZVfHtKNb8tyTVA9FQ
ALc87+7SA8PSKi97LCnMc05Ort/0yFUM9vyR9isZmbnTyQsoB2S9+X36Be7uffwG
kQaNa7pbK1E9QVAyyZ6ro/+vxP8Ui+qHYBQZFzB+tmsnxrJi95USaeVdiTGCxksD
V+C28yFiKUSjVhxsbXrAKJZbxmjez1r3k+9KR/0/r4rKHKAYXfeHiOU8JmySzggg
tQ8Gyd1DZ0kGdIgwybY9LiVgY5+UZI6QiJNR4YzsKUolXigQQPO2xBPvb3stQdTM
UURs5tJxbQnz/Ttnf6DQDxNTij541t3HJZMZas7Ig86dbq4g3+9yFU6faUVyBeQi
iE91CM/Rd/nwTw09PJuw4Y0AQQcFIx6i0GTAe1IoDDOzuobQRJwRpTtgFb2ASgr8
Cp6ReVr9rRjurlMcpqNDaXdKm9NFm5TZtm8mTCzDWFFRiYTfaAKYiLMy90kKJ333
jw178PPs/ENTaMwl7qQ98YECFzXg9+fUck3mDfJCU788yT5Lggm2GaFdVJTzaumN
3yyt6GOEfgWWEEEFecohldXD5CnL25WQ1yphGUh7wj8B7v8vLxX1o1rLqbVazzUi
POC7IzXvqe8OJirH1uRv549tMMK1oC2gD07YvMWqUfBrY5QIv8oHYs84clKceZEV
spZM6RPcp711l40YPar+rJIJkMqC2GXmC7K9wsKjoqyOo5T6AIqqfsNIHvlqt+mU
32oMJHWw4w93E++my9hxa9Zh4uV3ZiTx+cyH7qZksA4nCygLJClX+G2YSNJWeyl2
RrURb8xxQXSMYVWvQZRalps6BvF6WcomNPuCxAzWBswVmqHfhI/PXZ2+sDH7EGZA
9enSBSEZ9RoIUHnzC04NHtn74BrcSuoCY9nyDz5ibbd3/tDCNrkBl1ss1f4OVlsz
PW8XoDY1oCwaxN9mfp2K1ZqEVD9UK99FhiXtL99n3yf0Zm0eZI1tv7nW8dqnIyWi
9p1qkqGzrg/rBnrSICrqXqaY0+hv7MOOk3xTtFG17sDhWqHPCab9/aeD5HU3oUDU
hCa8RJr8KucBihJu3Ts0PIYtWib7ClO9Eutm5AVI1ep0hbcd1tG2Q3p3LRGTfNPi
AL5KGsvLcvclnmPipdb+M9wYx3P4J2bYu5KcDdm+NeUlXTeypdsp0jc5req0qliG
TQaQgnrwZBqOmzTR7sc+X38zNF4NzDUn5wjDNI8d/lomSonQyxR8XQSRFb0KT4/4
yNuu4S8B8bCYCHNkynwsqH6DFDvMMwnWP1wflr5lhPOZja+XBjpd+8VLdnnn2+My
PMpKmHfobws8sOE/XXXYzOGAj9A/Y/cCj6NxiStTD5MM4Zsirajl+O26TdflzHre
qjIvRcCN58C0iMDRJ7T+OAn7K0ye1ZCOHl6EdEadl/vv8hB551b+WyodEqWs2xXO
SjtOzjz0DjinQi7sQDAh2dwCCjcGiKJa7na5+dnu4AJRRrUxdwHV41m4QuqLfDjT
nsAvWB4Vqetwif4aMTeYxsxc6DDBwFDr2bg23rhI5J3SIw/jsSVA6PpQiw6C+jXF
AOeKlrWP6NZpgohcyPRElhJy1jSFgOINbic+w7zPxe/nvU3A6v+qLE19mGuXDFgZ
Jgcd8bLxpFy0zG/dEBDBBvC9CRRJ7B5SZ1VwhiGfH9CFNE3XIU00t5xo32scXder
xfXgXuXamKGdBroafrR6pJdCPF9a0vSTK9fOllpfo/Zs6TwQ8t1ecrCDhmkaek5+
3nIv3Y1o02wJIpIiGOy4hZ06DMpHfMVIxJBxZ04nQfbNaqyIAHATzlIao1671td6
tvgceiJMYxX/tpofZxXECVPKFEeTc7dY4duJ6fXhS1JfM7PrUAPwcAHzvWWSMFto
zTGEszalnl1nbAvRS+sSRxOMMeAKP75EZ8kjZt1cY2yQkkwa+y6KzKTFeNR940t7
zmVTsP5xg7cNURDyPjdVclo7qiArQOAcleIkhrjsSTWU62ufJCqCaO57LZ0dBqmZ
CsWA8KFU+3qpJzR1KcBorSitnl4M3gNx5HwDz8uVkPYmTe7k4e8acJpyLdXis+nk
/RnUWfHmjKpnMf1Pd8riimBCSNYYnJH5nEnh4iSdSuA+53eXaxZgMUbawQYvgONv
CSbmp5hAk33j1hMuyKkhVviStsos4uAN1PTotIezAcFERKznLoySLDFJ/iTrv11F
0fK6rZ+XG/RbJKXyqDUVgtUEgkq4C6fuPfoAgtpSfIThWZZ9tvlBMnNx/NB7xINq
L41/pxnS3JJueT9MyxAz3XYzEZmSfH0vB9wT8VHZ/zOmjnoZH1VmZdQoR/uWS25W
NQERkZlFkBl7o1AwC/aOC/CLmOy1AdI4Iu3yCm8yuR3HXGY385BAp0wVQ7Qcvtog
c1oBi9PSXljK966Bo3wJkw29wOgWjhaxSjv7Bdl0rLdLhhhje54mAwxOgXAQW+Ja
mNNuNw13HgEqLLtsyPpgW6mC8L/4v+wQaH2dETFDp8QGI7lbQHbWf6lhWz5zRQL0
+6nYKWUA7VVzyvU27FZ3qEuawPEza243+HT709ypS5DNQWwdfGfGme7red2JJ17g
i7WEF42N/rknAKZ970JDOltuqfF1kUtfOxNNUrwCZdi2XtEGqKLmune8rXB48F8A
gt9Ovqu7GdHpOyzG5nu7vyXrBFRtRMLmMZx1nsoCGVVorZr/yIhA7FnBvgV6uK8B
+Wz97WWA/4IC9j7i7JujYUUy2DSAdaHhRwJ3o6cRfMxUIGVMcirSsI3LFxWw7eVs
QlxOi17NGjkEN1NtYrYtCWRLz18oKDltlXarcz4HbnFF77nmLoFSUMXBBKCtwjhs
6mNeOtCYQzztGpcYQAvvXj9n7rvYhUzSO+RdFgYq9x7FxbItH5+IbcCl9JUYuokf
664HJmMxM07HsI/wxDjfw6t/J1Udd/HEDVzBgXrJgP7mL2E3lnwprodQetMqnUft
BpeiP32k9V3nKw/3l18NbUtiMUcIBrRt/c54TVClkE0jk3lJ16EH07T9Ry2cG8Pc
/IlHWFznl7p3v/hAM6JKqAJqVUyxeX3hMFNn1vdxutVJr3CNWLzk5AeiGakt0mlz
R/IiHiuh4f0/HIErJ4gtszGZtURkxulpAVRATK//qa4g63ydGfEEeUf//DCA9Kg1
bB+8cp2J8z5QiTwiY7d6xF8I6SHhzgkCFK860XbLW9A3chyzSmRDGFcQqFygfWyp
ygCHd0g1dqTJ3XEN2d9Py1q6H626FhP6KayAuWEY5vHKY0QzpQT5Uxd0xw49DLjp
GUJz1D/I+VHX+Xg+ujke9fowO/wZlH6EoW/SnGyVtFTJEouwfGp4yZpu6R3WBFZf
ezUtluic0IGO1YPXXu5gFphtjaghsaP0xyduHZRhIYbo/hOp9nKH0Xr5V+59q62P
RWwEJuix5rqQ6sV0IGgyVGFCP+r3NooKRqTlm7JeQXpAsBUfcKPanB4lRUWD9qnw
+eTD/IP46+hyZ1LhFJCO0I4opSwtFfTkqUiV0gB/SMqW8bNbdoNyUF+orAd6JYtW
LKEa52OS/MB7apbeoKVcl9HDC8SC5yzVoN2Q5dRSMohFEOv8rdmHxC/rNuXxlaTj
AUeZibQy0cJGfTnXClWP9DJdDhgPAIPQS0OnOOnCjwv4P0A79J0NIEmYWqWFOBSx
Hol4EDeAwD97y+1zMaX+4vdpzrXcr9LZxg3kNhyEbZVmNWmV4jBLUfMoaN6AXgou
Z9DsvpJIYLrXC/mNN5ygtnGtwhHD7D1cJPAGrewytIy+HUDCCHJ/NZJjTALZe3xD
vQWM4PhxhonWiCdKZG08BEwWiO8mJBTyjULR0dK6pal4rj5+2qNwsZF4amhWB2cW
bs4bn2VfuHwRT5nYKoTM9frVp70bcprwbzn0pyBiaWPmIVflEXDNKTDxroMzX9F7
bQgJr2ho2PNKGFBI86V6++2Wjr+QitdW2SYwF5btI2Abw96Ir3TAU+S8FuXtLQl7
jCbyMNYga92t84VWTUrVFwIPO5TCv2RY0fgwor+bCDlTKE7PkGHUO7so+0XRSsUn
2Dm/hLM93XEp5vXnFWqn9534lEuLBwDsxClJQrVjiJEXn47mdgoF428bs8APiaff
cmOvi4trbc98yBWmczznI4MdVQ0AbUOQjhXOgjkrB+afZ5CU5tySE1tdLiwf9a2o
eVg/upYOrN3iUJvZVjoCZ2ijFMOYyd/xzvzD2niC0dfqfS+pQ29SYH5Ez0IokdUA
Lud0uXJV3hB6QceAfhm2D08F5XGRJtw7nHMwZXYaQQGHGKeRnv6+Op83SHjmySHa
l8VGwyjdesv8IUi4xrVkwoWsvcP5hBIBA9od/88WrjffASxzW+nFqoFKNiBlAKmF
6FPb3bdB6T8qKF/8SkZ6kCQTpSe0vUMHFUtMzE8YY6tpu0dwlgCMZfPWFm2R7gIy
x7LyENE7vRZF2H3YdhKkcc0+95/KSlOvaD70/HlPTE7cOJMaQWw7n6K/WIqDRRmL
NFURSpq4Y378N0apOEJm5e/LBZKHx0ReMRMrneU7SGC9j4T/VrYOM4jj/cglz8mW
0IWhZUVXsQVYPuXF2195c4Q20jm/6KYEGH8bVEVbedVysIDTPE5FaWQ9QtnJ/MjB
iifq3iwmDjoM5BOou/jLOgpb2zII8jniE/98v66C8tGNgFCUcd5v2T0KukBdsf8y
Hng6kdo+DGqSlJ1JInVfYuJqFrRWg0eYlQAofXUh42WGbbuw6l3o8gfC1VDsJS5f
oI8KgEy/xvoj8Dt+6rzu8MvP8Xs2GAtwN5fqFTv2+KOA9Bxv5/j9KNfaXnR4l4CZ
aoBFkc6+khNjOesMnL5WiwPiS9GwDbBp2SelAI3T62frYRxnx2KGY/yAdIsg76Hb
hIU3U3uTgS8M25hRiqhH0PscfKFUjNoZWmhqQfFFoKd08dnBwWluiZk7BgD+iiS8
kchQh89A9RSJWLXnB7Ke8cSG2IdZ8UXusuZS2GkW3xvN7nrkRgUqYoMqO0QKF2dk
ng8kmSDKOEw6HlfWKCZINMKtj9Dncx3cWIUxKGUCAopkl+9p+kc2e0XcgIRKAl16
z6UBj5DFDs5CYFnkiEp7/tN8XkoQ9P1xONMNLBkAVeUSeMYiZLKT2SHV3Y3VmV0y
x/jbMVhPo1JNI9QQdIYoACdgpLpaWNDDy3de39+ADZrM4j7oKtSNNxbXwDAu1whn
WWzwEI0RHjsLwLiXWbOXQ/7BXBOekwimlgWhFNPuBTFjK0bX1UmrmCSqygVoyrUI
lwbKD/4eOnuwQqmAVGo2BEd0cP/v8wNk0ha6DNrg6IN2n6GYQro/ZQ7X0mJK6gAI
AeL1NCCLGS4zmidzKsi4YKtTQHZe1lD18Jvp5tjc3T1Fs3twz+ylnzJhhFhO60l3
f+ehmkXeU702da2tfWFDbvNwNSr/tat2rRObg0EZj5aBUKEDTBykPIt0fUR7SsaS
aDKTQkUJmMlce+a0iwJyu4fVjZtHNGx4UdzO9iqVfGlGIcTnalHgCkRlgm13ZOeB
AX0i9fFs9EHT0zuLfEtRALd7dg7QQaFh10JvDy5eDEa7QE72jx51LyQJDc2dSeWa
pwjeMg3dDRh4TmhhiMH6yLo2gmdXppMMW4LdlmAwQsGr0Ozv58FZWEAfqAftuLxI
kUvZLloMNHd6CF9abwjPW/NLm5P/ePEFS5ZlRjtviK6euOV9c4iDpSOHIxJsWeW9
xDQ6f1h+yzcmF6U1a3IoRZu20kx8cpFDEmuDIq1XVbt9nQs1maZY9FG8aGwzNiK4
aSYjF6ygXLOd4GqE5VO1mgLA4KfYxbl9ReKrOy0bZzNZHBSWI2Uwd9YDCndtFEqu
+A8mM2PkvrS/yMnWpcoEYyUKZ7klUbpqnZ8dCcKHl5tsmu72S1rLANlRxZaYT85B
lfdQUha+1oWip9TGJ5tgp0ufu7Fd8ZH5n5YVSw9bJ+x8S4MzkL4OY/h6C8ynJT3u
+hUoNKcYKgGAgq4ma4rKuE8lLTwpgMQiU4a1GVzCzDmp1qcxxaPugcP+lvF1an5J
AUT2i3ZT/IfQ/uGSEsF9GDTdD2pNjkW8BkK+9uJXR1kCowN9En1TxUl4mK+roNWx
btZTm8GU3q3zepFK1UQwfd0JaFW9JQK8xaLRzVYhW1v8ie0/+BgvjOtAMAGbgisl
AO3UOFt/D6o6M9Fzs+Tws+uk/rQsglAzIzTeicWAfIRLHHNB4+6lyfHH+a0YAOJf
RUUcaXPF0UtCJluV/WakfhMKNwKyzwOaQ2nbZ2KrqGh68CAXqZx3J46JHZBIoabt
fGR/DM5xAWxP/QrXayyy2q0O6P3Oi5pqvqgxc7p+KSQNPHJMSxb8JQN7ynBeLCuZ
Ah+yO3PjWZN4q15hdA9hJP2dL57/2JZmZCdK2WDQfF/D5BSBhk0oNjBQ3THza/54
LlWnf8Az7da4fJsQPfJan4aW6hXUTwC8oGUMAY48i1aQSu1oYKvL8CaN8eWNDXf1
p5HexG8aDXCovOGFHTb95O+CtllrxzgyKTMdqQyHFp/z9UTfzujsUt4w5dJD6KLM
W5N1XmTB+uqqevR4c4iUvUKibihvPeJfmNH/VtqR14Ew2wfjhWosfVLAnVH37ACe
pJvmWGZsknEkyxKWcL9TKey7dRyQeYSjOPHAOKG5uzIvr3EhiOFcf9f2Lc9kXrJO
al/mpb8E8q87J/+gvDG7A+02sEEBSrRoORr8gVBIQGOahywZhaz4fxcwqe+AaM0o
P/gpzMFSnunsEK5QxjuiG/H8By+A3jSZQan/0z1pi93LYQTIVKoJVzLapKQKN3rG
Qtjrt4dr3fDyKmnHhnSovHIiywksarrl7KjU8tt3626MltCCd7iQSEl8KqlSPWRO
kJ0Le8I1Jwc+18Uycbb+pmy/kxZJ+99n69J8G1fIIng4WoeXiqZArpkQ1/YvObt0
P/O9wC+NSJh6OGHts29L/4+LEISi0KXd8XuthdcUKt6994tVbM2rxO4ArS6fvnuN
wBTcy8VYZ3QIamL+oeyd1HSBsEmjRHJk97ai3Uz1j4WduVN4YV+Mrwc1GfIgBz8o
nmF7RUEckVsLV2UKkqIs54P6b6hFRLUv6rvN04YDFKJDVJ8PeiL0NZLBwWiGZj0P
sb0rhX6XCTXBcP3dnRPN4S/eulPcN+90q2KgAhVKom4EWuYOz5caa8IOiRe6ptDZ
SWPJfyukwfeoqHNJ9lyMD0JTrlcYis1MVRmjMLJ3I+0jbiBh04L1mpH2XOw5swLe
8YWsyGzLYYqYoD2+8sbjKlZXTePyfYrVIFhkUvP9aV4APDM689smnSGZrCbowla5
2iZmqDoV+2WYrgQusrR5zr+USidvZs+VVZgSUcMnf1yKjYZz56FUhZNVw6fZxjXf
g6V1v6PjO4J7bBTnm1w/BtZWr6jzqsxS8JYxDO3zPQxLshKj0tkTPdOBP+RoaNsb
ECwITBcgCRO2t6mnjJzgq+LnvmPCD3SU4hHtfL/czHZMwskaFKuiiy9PXThMgX01
ulNGmM1cVmcHc1gqAr4oRRpQSJsIf0y8KgrDDpmW9bh9jUNEyxaG6QqQrxTrk/WQ
yso8x33y4HIoDdgq2BC8FYCvQD/HpvZekBn7MIqOVmyGmKW4YWLcDScAe57Paoeu
8RjGIZFAJNMzTlPjRKU+TAFFGi/FT0Xa98B3Vnj/E5JA0Udv3gF4X32XVtsszZtc
miAtp+0zOV0h/Mp+3LsccuXLzfjrLn1BQKbhKr4Tdfz+qbpdLvQ0hwdXGadpNzsi
tTbbib8DdGyLd/fA5C8iMsgTi+km+Wk6kqZ/x1MMKNOqBcIGtSJ1wGplZO24ud7y
YqcD7OJNDrAVH7TfCen1u7sm8tzULj10pRINhrM4hcbjUPDzNqmmKTE8M8st3fic
/ssTdeBDu3J+5EaQbTJ1K7rw9GW/EE+bDhIklnVmWboZ2elA0GQqSUnYTYqfpjDJ
22MU8Fh4mgE/s+hdPzTGwlFR6thws92SsSSITHAVFYrOG5+sVyaym8WbpZkad0+l
nMsBhTClaVkJAwalEQ0Se69dSAgXqVIMisIr0YA91fFxHgbMBlud+/ZUptB3LcyP
UzR9xUeEDqg6SynhSVer3FObCb2CPruVZ+nf7NasBDQLBDgHpcZJeLvtMwaI2Ddi
CmVCVfQwg8nZxVcNSOnWIhNW9IFbmG098JoQsJRjwtYBAkakuUOw2ACK/bRlDkax
UzlSba+MrS0LhSp1LhIQR4f10hCWEAn9JW++SLmZGXbwmQIdgD+VHp56uAdnLZgm
JkZ/hQG4WQ/oeVRJapYY75+Azx1YQYyOtbyURmZYIpSvCima5JzqYyxuEipXsmt/
YSZWYmFeKJRgsO7o0l5Um1yBogUkTX0l98Zs2A9qX+9jPNdF5JCacI0d/Y+4LaIz
GKlG8nRlaqlByU+KZ+RDIUJtKlqKWD3VgyUjtsgs3LQVcR8SFCUvF/H8+DeB6d7o
rr9ZJE6MT9ypHCi9TNuxUcZ67Jxvetia2+IXiAC3GAgawRTgaSPS8nEHLIGzXNyT
rFpqSpSm34uFFnRKS/cMrj0SF4bmJvxEHRLP4ExbzPLkb09aEvaojChi4OOqZduB
OPK/z7fBJJ9ZZz4ZVL/m/9ERoNM0hBkeTNm+A3NEcq3IWyGC7pDFctrppBpW4S4g
fihObf20ba3v4juo6ULmGesNG9HLkZAmhYBfQCaKux/Mbh50aNXr+d+UPJcTqY+M
7hrmEz56sd367jzofgqX9W6qoOjy9lYwcD5YlmeNEVAQOvYLgUejbpJV+k5yMjTq
EN9TmhWNKeeAcAhx13ozDh6DvlxlA/iwO9+mAjy4tqVLsfS09gWl8HoN/4rsSCcO
DqCU+GPWrIkm5mcdh9Mt9W54ajOpnRU58XmdSQFU0NZt5+XDhYPircZYflJilEvR
9+o/2+ERJvCSs/yTCsWq5LejieBxxs+6txq0Mo5rjEhnsu/+iOu0LTsCX5elVCkn
42LIuVs0UGbQ0OGoJCnjyZhjwgAh0p6GUeoCAfCJgOnZvWf80WEwqBtilqXfoJgN
JaTAiVzEsEQ0b/UXSheI/Jb5YbJ9KjUyPTD1ol5iCwr03uwQ7Gj1WHUKwHT+RV05
csB0Rcjf0hheaa6gUH4sg0y4YiulV9O0H9rwDuzfkyHpUTomoq39vXTpG/cOhHAA
7dmz/5M4RC9a7eNevZpkARTi/qc1I8yC8wlYNhBoOTicXx9vbAmPoY1izoYO+q02
0AmvG+wG2un+zxPlUEf4wgJONAmGPu100Unyx08D74n9BlxETW2d7elWIISJEM+T
Zcx0uz1Lhfxle0/Bbax9rOYqR7gmif1rnqHlVbUykTjS5MmNndGOY7TGf5P3u7NE
JlvIbxwHOzt6jRGE5KgXvEhYfJtpi2OWJIZuzIslS+O/qUFHEVbVTF+pr1gbPfZ2
xMn8/iAp/N3/w+uJPdHl9qrYiC/2v6JWR4N34z3n2bbOZeC5AbXO1E8aRuQKH8U/
YYM6+BMxG7xoiDzxtfrUsB+7e4PT6PU1h3Yy2P+OHJoJKqSoUG3SWhPFrt5MlhMt
IVIQK5A0BvwwHDDCOc1cI7zBoQj0ckKdVFsiP9CvQogIzOxpXF02YdpFrARkmmPa
598tiYS/NXMsPw1KIDopMZt/7RUpDOfShdnVMm1D8VAHVbCJGaHSPr0QoTqgIBCi
1s8fH03LrmVS/wSw/EcO3R7eL1ZkHHXVqEQXDsh4Y79g5cM/G0siLVGc9fpRzwcg
RQs2u7nAxQN68BZlk8q/qgp0EAJ0SoyEvBSt4OQpNL6DgxUr5IOiNj8GqFS48eCL
4mjSoQYhJIHX3oGXZA07aDXf6VeVlKTcVfxJ3vtxbp6ueqOz+D0UD34MA8sYyd12
u141RK8c/01UyIjhdwqnWHNqf62yzhTHK7nklPuzz0HS3eYwpZusLnXlhWpCpkPP
icnM26sgKCD9NoF6iLvvuMNGkRHepZ/7gmV8TpEfYSQwysMJXHH0kdn+YcvdYXNB
+b1HSGxBrvDpxhzPkHjBLEuYcyOWtVMw9c6ZEZCX3nexJSfTD4uZ/uyGkSI6bcHo
k3WJe0x5spOx+HYieGEb03RFGS4DU6T2qnpdk8bMrmyd+1ayZNTHHoTpPxoGuNiC
Zpf6DtXUMfLGE4Knnw93tlCtg9aMOXTjgP2fUyUShiRvF+fXLrrbFYX+HJhSug0u
FbXxpbgYr8WbEtsL6+qDvxVRUILsFFZicOVugi9lD07tAnXmgbljISLdFQB2G/o/
n8FJ9j0HIhaNqCzZgREIJswwEO9QZPr1C1USsKeJAWuR4moPoE1UBPCc5V9ZVPBT
lpQF7lKwvnbl+eiY1vPJFFy2cqr5eiQJXhNbNRqCrYzEu5tOrLszjJ2A/pyvEcEb
PHNGpWrUU30K1HU4OHzVhIN7I5cOGFv3TgKM9YSbQvskzr2V/6lhk874CyDvXd8w
+kyj4vZjC4v2p+IpMsODTWDFnhkECbsNsZQaqXYPD1RT5s02+ZQlh3E9N2T/SYRV
ia/Q4FQR4s9eUfc3SPQzcN65BeCwxfO9dEzmsK8+c1k3FhxxVnCD+q5Pr04YIZ5a
B4jYdMxNHmWIUXRc8mAMQzGTaeK4P8KFcH3pojCRxJL+LPtwr64Q2Ffg4VqLDv6Z
0+URkB1godUFhXjU+RISEs2YngcIPQDD4czf61p0zVbO8f3kIBx92UmpkqOJgUvM
rHeLiX+quLCsAy80wincnUf+aWecqu1IfMzxjQOxhMYQYPjZuRKPt4b2QB+Cwmqh
kEjicGlLEoDlqLiwStqpmcNE/gTQHeuJpnvV/Uv8CwuGHjpvpQotQs5dZEnr8Du4
YvVm9OmDYn6EBuEtlnzWBefnlhNV5JDuE6oDNA4MA3el7e2z4+acZHSLfJQc3dsE
IWWKxETfZN7a93YJRVuzDs9k9Bj7cEkaq1hJdoYCYnJik/jnhaWDi90cklsm4EqT
FcipxT1xzFkcuVIAQMq0ep2eNgWqKsF34hX1MHmPOKXXCOoz8fLo3g+zwuqhB4UI
m8efbY83ni2tYFCafVVvkJ4Nwexi+yyU9arCqIffkLuBvqvhblAcnPiDoMPubrCt
80fy0LG0M4myP1jenV2kBe5q9kVDEhTmNHTZtBaPw7AvVh6lTPg2yTItfMnmo4aM
wyGWeozL7LMFlgANdi2nQZL2+OSfBwlhrwhfybzESBZX+i9w+/oDXQGgbl0393l7
i7LNPDoTvDq6Bbh7+USUC3DtNLm4tz7Zhx5aBY2ITC2Lu1tqH//PO5/4um43Lsak
ibPVYuBrjGBHbPHpAexNAK3Zu/9PX6SER9kgBUrdJel219iQgFVB9cmvUitPYZKj
YeRsVZE3b+V96ThM07mLj/cpr3RUdsbSyFhpMMAzEgyMAc1yz5+0r004zlSl6iom
mO3I9YlAT/bc7Sxnv8bFAlKBbBzjtWpGU5tLWANL1T8tR/M11sp7KsqoPj+76owE
cu4OXAdi/umq2eajre4g7WFu88hzARIPIiSFd9S737KaD7bCYL7X1Vsuim9SqViZ
vNMq04Q4GNwKecEWC4huLTc6GYBPc5TDFxJixp4uOzv0PNZ1aBb+jRuKaXk3XSlZ
cPUlroclaH25zPvIQdIjuN3+hwKKEyleUHMRyV7eWGUHDi15ltk6frzvUoFwxptp
AiG3HqspULIpzGu1azcEDcT1G36g4wzKVava89HJeCZjFFMa3KeFxrlJcM2KUwHu
j9H96AxHdf4oLFNdDHWYs5MnevmEMKoBA5LT0ApjlCG9jMGNzTRQpqzjCwVS2UC2
kchwDMjSGsc0e0lOkBs7LiROqQNCDW28dkvL1TIN8VN0DjDtKGNu3qXFb1cwYXSn
LSAjbhjW3pyU6cp2umEixSFkGhFq+YAlq5BAHKCm51hZoCVM3pNHJFbWQUct9MKD
ncp51HGuPuXEH3kAhi2NKI+/SqQkw3Fksf9JpYq8pbDjZTnIgaJ8yaiR2TvDlhGY
yzwQxLLpeCNn9BEYrgdS1/9Kdpg5c8JLSz+K+HkS6I7RZAQuhNVXHW+d4P3bZJ3J
zTEGuaSl2U2nZ8geHgrv/exQPsFdCk+ICwix5eUTd0VNPqi5ZL4cRmXM3Ip28Gdi
iQVAMWeJp9SYkNMAJ5F/zJqLh1vsjtAzZX8uQd3QNxLbuhFQmEAHDXXrOiVOfXXz
KU4cvw/4UYn4yV+64ZhphGT9PZgRpb4bBpaQumf3Fp/mf2PhTU4FOCVmEUX3i2En
77Fqdc5h4rr0K/fbF4JP4djCruK5o7DL8MQE89ao1ndSup+wEMsKEd1DVZ11b0LV
G1ic7UVo1WihyoNoMpyor27A0TsiVoC9AB0D12ViT4h2jC4t2W8CTLjfDbDI5g+d
ZD2Aw+W85BGPajfWoV/+ypQFvF13XkjmB1ZGk1kMzkmEaBovRHzmAuec1pFXnjcj
BqyuFstIs/MdktS6Ze4pXFQ3nl+tNKeNuygPWxRAv7l16AF8nRGtDO26teq/Rsxu
7r8Naq7Pap5XFgm3USnfuhVDpt3bOy4erCiyji/zyM3u/2BNzrN9+vVaKSQFLpDz
zJZf9NKfUWwir5Cz0qovd1EUrlFzRjNmNDuFUDmZID/nUwIrno055/iJduDghGr7
7/N/WmA4hBvOe0h2/vW7PBCiz7S5gNmJs62ouvi98Ll8DzrCtSd8FivbPSnUAnmR
0zSC31UNK0cXNOGlGKgGke+oxlyXhY31PTNt7OelRwu801r4HKxXqve3fiPuli9K
cqL7TN6G9/gH74xIKlYcNrTpSr+f+xlm/dKhBaN7jqOUD+PT7GUVn+za+CHVj6ud
egcm/chJspwMqXCVPmnB0xHO9KfCRyH9dUs9KOlyJvs4IsdQzO+DVTeJULGxlr+I
+vg/QuqJuLCTo4yVT02XHPERv20SWcxmvCvuDhp2xLofeh3WAPGNvkTNhF2iPAFo
DYiX1BpkfD0deU0U1nXxNi+Bj8RlL3ncVYLf9cMJsP4O7eOrP3kfBXxV/tHa6n3U
1IWqAiOCBsL9/Y3BTPEVpsd0hdU9ld48NYauCEUqGD5W5o9bt9Cr9in8IlfJV48t
UCvMCxHudjxxCpOzeEdv4himfSFcQsPCkYJyY+NMfcKFLpCcFYF4X7p9xak0kgF9
hBBRqF6vDR6WS+/n0XDZ3+9kpP4EqFGWw2GJaxjN7hWbNIURRT5A3ktyjkJ26KN7
qX1dhNliBEtnV0JjRMRUnIH4GqGaFJn0wh2sOlatVfOwGfmVMgS9M4UF9QG+ksKp
aKaUsEa6FNNIZ2bWexOFb2s6fGLZErZaKhnNdUVD3O+pg/Dh0fn1w2Ty8J8GGGsG
Nb6AArtzAqHPUUx9TyhBWqrPtfq6iYOxUj9qLDQxDWPsAIkEsURtvTd9Yiv1/bQu
57mOJylLQ6gS2hI3kEQ0H4jO5B1GElTem7wG+x0mtSRkaHdERfmByOXLIIbNSJhd
MAE5lkLPgCa+T/BEqXiAb1g/E7m4kuZjKq8KcelHin4EFQaCoTH7RXOwRjSLx3Ku
25Meew9LuU0aTkeJeV/C6MCvbKfEpgY2KsF0O/snzscBNPK9K8igGt0EIifeUbvL
8RRaECzOkRmT+33n35IpYx0Fwu1siGCXD1Wso/jiLAt3+XUM4hR/PxDRHikxf+G+
LyFtawWI56xXRfBso+2hHwJTDPthXaQjV9VIfFQVm0twFlP9Lp4J6Q1CIyaKsNqO
Ww2ic2JepgKkjfNBwGTK8PJAEMyga1Lalsou/3llvEFxpF7iFthm0DPMZUKB3yZd
43EX7kzRKVoQg4HP7w0SFyec1xh8vf5ssyfL7nXuD1R4sL3XOG5Z8jb0Tpf00rAi
ZNBxUz254qOd6bLuoZKZi+Kn8+XU/VJsVH2kXz8hoPtkt/REjoxgPXyFtQls+GMc
PTKMb23uxRIuVRYxiLjyxXDl2UDQGGH1iKRhnesV11skQ5ULkJfRCz4XowTe1m9d
2asi1QHYC/28696KBF65eyYorpnavAa6rhljb9SGfTPs0GCALb+9I6nj+x7cI+o+
9A0Y6BoxIzY7f0kHDmoCBGkq0tgJz9O+/mxDoh3zK99oWYH0h+0HF8l62c2KiN3Y
DY/vWZX+2mn3AguCXUcOR1Dnz31B7kipWHNDE+bwr4QM7G+Tg3xoNRFMl65NojUX
AGFlN3+kjjbYh2HGt7wtFODJTBIqFWomCKyV5ZSkp55nd7S0ybx4ZRDnBYuDJXvk
HFjCiGG2Ci0nzV8lJYpBGcSKDg/OjyxfrVwVNwOw3GsDJYNFxRz6Qe9VvxmyD7sx
FiXxy6IWWm3Xao8+jWlgASnepIkSRgaGj5i96Ka/8RA6UePPRJUOogk09909Nlw/
nSKMHqwe4bkEeZOxLAAe33NCIm9cKGEycp9zEBPk+eeRZl17xrnz+wFm2OFRA+l6
+UPX37Cc1z72o77BO4/L8enmglXRuiQpkp6DBuY3Cngd3aXBYLW00M8Vl+DG76hj
ccZLGF0sAmXfZzDHUEgyXKVXgdOQNrnfP4c5zHJ1QqruPg992SM3FI76SQvAqGxZ
3OV0mOJUyGlG4Z6niomh3jA6JuFx4idKgCi2Q1/cFygly89X0TpnrMth3VYV8tOw
U9C5yDd6aklXZpHyJ3TrY7NdXXdA5ATjI1/HGoaDg9vdtbuu+lQzoiEiEK7NJKEa
OyRPa4fh/icqa395Nb9IhAiGZDTHyAHRTv5uD33IdCrBI0YZ6aFXBQ1mV1BMeDEo
fH2OquAm4cSXmQw40YAjQkWNtXRBz42mRZ44sEk29pQsbM44qqqgFyvNgjCcGAWW
JdHhr6b1yPg634V8yfVd55/CkGXp2c5/WV//ABa6ITAp0IgFfv+XOjPu/21cdH+7
8urr61SEKlK/0E4HpBmwfrGJRytUddbfMh9B2Bw+XI8B3UbyZFVXFyWb50yMhbCa
eBlpgsAQ54/Tk6PYAAu8v8Np6jFfHkBkxALyTDoA1sukGczq5xBvrDlOd9bw5728
Fi5qz7TT603dH91+OA8/rp1lcfa+/6/SS/hx+0mlxN81hpsBFMfltfWh3gstxeOU
ERLITQe4pu7vFBVqOXee2zV6w1lkSDs66XREimhYmwAoEvOReaHwFKHMGKyy7pJ9
D4t/HhiwOggDZhaGq2YH9rX6SHEbqBwlv1/ilQ3LI8j0cWnLTqmDlrAOmoLojHHm
okv32gMqPlQk7bLJuIZI7rLpo9mrgwiCD974QmfqeDDt7Q9P6A+390I133Evw7Ub
RjU2zBGu/BnmcS8Iuz6VY1Oy1Ao6RsDQmskvq68fhUUG+uUAeSrgymam/PbOZPi3
JtxWi6V/ucYM4c4pWiyjeI0x4ToMEHxLmprol668NNHzaLyIlIHTKOiqEQb+zasA
PEqHQ59LTL+jidmEpNYmcbTh3+ZUPH3CRPpxvGk6B2lVWY8ZyqK3qPien1mCD+OU
LF0dTDoE7wM2cxL9ipbAQPCFU81MnHfXDV2eMQB+iVPpOZOiMcLB2wFWc4nn9viV
tGNfXA8WIOIkg+q8gkxl6HnGEJ7TVoVC+Ipw/Dq6mQ0wSxe4y3+S0c6qyENLzD+F
pfgyldldJO/ZlwIyxtJH4dKgc+l5VJQmwbdVRIG6hOtYCbeYbEDh77fTsZ8KUmld
9NM+MJBzROt1Q5S3Eh8KxKtmQX2VHn0CvlWLu5+OHR7qw8WSm5TEh1Aq8iwN1gf1
Mslq6p3rCDP6wxeFZk9nh3hTOmS69DHKUMoxFVOQGxuSwH6M+Swnz4bSRPDkvRFh
YBzJezy8nk3BDvupbuOQ1d7pEpDtL/kLILxdCJkj8tyGkdgFYWSh9vqnOzkHlQ24
xLyauYUzKG+d8Zpm55aZtbRMSy2VzxDvTJltjmI1u9cV4i0mgOiU4AH7ngAmVF1v
IGmTH0/dk8RGMNhVlWoXxHVIBZltFuYq8gL8iphpnug6A3TKRC+2EXClVeQCRH9k
GR3rZ0q+Ej8WAT3muIoATYbEWIToUYo8NULCRvOCRT+2kjGTD/COoY+IruA9djwg
8XUATeNvm8eWzIrPU6fXTBrYziJ48v/oVPmEikpFE4yW6Qjg3O0BmhkWD2eSGoVe
uWSdVAEQFJGXpw/IpLpqyOdlHnn7xEsFzcQzW/WozYSwTAhiY27pSSTKFkHkWIxp
xWIIC/TkwCPlEhWhFON58qPAV9YItNP3uotMo4yx7/wsKIBVEzLxdh5zNn+BdQU/
/o+0UquwzuPqOeek9B70BhY6nS5HQTaPE9bk9VrzEm6ry7QX4hDf0iB9Y8hICQhj
uDM7GO1LbLBMX3wGulI6Ze9gQB9I2SjKLj9BTC0MRKfvRFv2+CaG3Sa7oU1Rzq7j
12gXH9JUQZQ/jo8Ftl6JrpGhzyfPBNy4JsjbvINSKitoQSoSL4MbLVEa7lg/WEaK
DVGOZIQAMlpeq1yVKaUblq6SwNXlUbW1ItMcL8I8W/OHsokbHhGZU6JltgeC0rCR
PU9XJXx4TW2/Koyt3F9YFwkkXG796gEaDWht5iAyAuWdzoeqSTh7RulnwMbLk031
lQbTJd2uXljh0K0x0xVYEkLsket1yxuyhjf6MbFDMLe6ml08QCJr5hUZ6lNvXezW
6W8mjcrqjcvEWBZBMVZezGHAlqZEeajbju0Jsa1d1/EUjPAzOd5d+X+xYFkQChfF
2xmTXzyZh0AKrehweuxh19S83RrBH3j0sFlZlrT2/i6YFZBnbNAbJ7NOLRp5KdAz
I0rakBRh4VLsvCrpWqYnSadofJmYMyNReTk39cbtWXpd0xlKahvC+Rq1asX4K/Js
ldnFG6psFdgPB2Dq07RKfuDzIYV+0gQ0QXLAEkRPimQfCmhFLFdZAOgmRH9esQ4E
13trGfgtYducHGRcDEq0+SDv2xlVVKnf2ZXXbGLkgT8lAVeN32165eykXnGmED+F
NkQRmrnPh+SEhuRD8Ppyh0MRHCysFyP4sQzjr3cuBttRBChtJ7y4iMbECgCliDjl
BvKaetQpZqTSUBnDq69oXvilh3spSOtLclnMO0h4Xngu6xkilXEHelg+QnnIr6WF
RQJNWjwhEsR0Mwv11Vd8gTxsiA3ZkpD9Rga/Gm++KRLq3GGbs26WU16+9hwaA9iy
qD6Sfevoag4c9HBghcne4zsc4Ea/VeFIMOEupAALxSiQB0qxhLPHili4PYbMIdsC
8T4mIOjA0cbrJ7HbVoo20odmxKg4LLIsyP6aSyc4ppmu1ouMJ+RjgZUlTjN+K5re
kR3FjwWE4dQoDWXISAZW5ku4Xu4yKN3cUURYpAm63jRog0irtCM0CxeueXpVHBpy
P5YkaEiQ2zY9YWAfI1j67HhE6qh1W1fjQ/PqaGJv7CkX3F9CMrfKA0yVi40wPtjw
laHEm29nyWUudZgyC89OszdjEBsuSaRm4F+7Y9mKealuD33d/wcNwVCcMRDqjwr+
ZPGJdTASKDLPaLa3/8UW1MHAKdOh2pAsmtyqCX4BzDXETSWwEdqmmHisI2HapCtc
R1flCY73dFtXmkwTxC/SAijzmfcGXk+zMR2GOnwxfWntUCAbcbSSlQ3AguM5r805
EYSE8rb8Y74G0imM3VEv00DPAOU3lUJKjO21EOL944uV7wXTAj5I5HzQwqb+3r6X
wPaSFNmEXQ4jAOEhvdA0RcDRcoAIOKe42cJRK9aEjm3mlgd4hkcK/GjC9QhC/8rt
CGpRdZQlppd6o8TjGCqbtm3/RrKqQsJ5K5GAqi8kVsxXnupEOAMmsJHLgNrjQyT4
b8EEhJDaKmACKtgo5iDrAwO1J11+pglrB1nXoIMHxswelZ0DW6ajndwuh71J3cUj
gEs5O0d81p5O+WSqyzQiTnBdyKrQMYP6DscBSkZRcdTnuVl9E4G0AHfLRbxnj50T
xW4QXYtYteizNM4Kp7pHGBJX4Z6mKmnbAkjOco6EmwzSK1fe6doUd1qBUVb2asSh
XTiGwElw0E9CkpoZh2u6fum6kc8qUXwfgp2M4bqQK/uZ9A8Msaz6TiZTnWb087Cz
t4hdAwLK3CckoL0B2Y0gBVIQqKINFaYfvKlsPjZg/1Q+20Lwlime/3JfFQMuhCyC
aAPufNSxGMmmEJKHvzyghWJWBtKaSgVC672+RaMw/KJbu1Ddh0SJIiF1rjvdBYPS
wELFdtWpX2S6HIvvT7VbDBnWtjIEzLIRmtYAPaWirSo43C7Wu7VECOQit9WUaNl/
Q3Ca7pGaEXFzVZkipK1I+dzb94No2qBCyMeMNtBw9qZodJW5mFQcswEBXC0ipgFW
UEpjJuGl2bhO47OTcdsRd06otK7D09nCmjaEg3hyHPGLswwWDWEy3t31gzpPSZF0
u/lhet7tGr4eYU4qPtkoaxMStH2I4f4SUOLjrjoT4b0BHy8QK4m0gqf9o+WRZa8F
4QeCG7MH7kgSxCmsNyhfpzUo8NOFfiXeR7p6wRF7TufbrvZxWespjiJGXyxRnqXY
+PfCHbdHgslZn33uLhv12XNftqnp+QrQ27HgDkHE/4A1vxFSJ7lJ5QPHCLxSOrFq
OVH/WG9HP5zhZOWJJX1hhOYZkmEuZQa2sprB6Vq6gZud9Wyf9/JkuFdg2r5X1iCU
oIAbl5mS5W4j98Rj9vgfL/Jgcnpw8dkoHoEei50Ftrnhz5KOsHs+QCdmKQe/cvp6
ZEi0tc/yvzfcrN38z7lQI+wwc98ozdMLX5+VVuNDPJsDYd7pmLH9YtDy0w3AaRB+
rfR3OURys77nbAQqngdqwhnHKyVNQySAi0pg541XNlsvKNWFyKPv5O3ahnLr1Svp
8Gue1EwDwYraIwuMjNS0OdpSNbPCLX8O6u/IBn0MWIf2Mb7ZEDgOC8Jq9X1vCVrV
PGycS4QRGyUFknEeJSnfvAwGHaeLeedkqYJgYvNxjQMTAq0GUaxoY06T15BsItKc
KVm+2mzKmD6uQbjhArHLd1Q+rfIcOG8hlVPRjj1xiC4hp55AlrNNsuzXWkOS8DxI
Fl22T0S7qUcU82zdAYfwgfvtwwDTZcZnEckTQHkJSdzm4M+zWkTisEVNQF5IkqhQ
S499clYrb1MvE56a8PiJaG9GZS9a3EcljCTsc2EN6qoWMam2dfnfUhhV01TQSfuP
ve1vmdnX09MKEMMyLXACbaipG4jyzvUCgHDF/Z2HHwUFhihVFlD/FXcm809a+Vhp
bz5uxJNECeEw+5mh2tqkNFaQdJC7l73NCTpzws+nOjLOt/p3jveUYBfkylrDyrR1
JQidkGPL+nnUDYB/mb2YZ44/ERHF29PWaCJbJ07hsFXMOP9b9XGuvgLck7Sx4I6K
Sz3Y9R2NH3tjzVuD96kwKYogEfqTEf+onPsOg/stcx7ESMd/PwkunmOWD1eThS0B
JlHpDjUspOLY2eoStHE/flEKnaW8Wzx7NjtvjzwPWNxOZezMI9YHVd7JfV44sfg2
a155QoSyz6tLUjsJbGZNInnACgwxRaIVZs5EExwLMjz5n5C9hRbwz/yuFwwsI802
oyrpVOJI0VjzLtaMmQy6nYE1Pm4g3Vph+GSHaxqppd8fEuiUkKWEDwZTNcNomMHI
hLFQ8mq+51oYoOE2O5OZL4hk+nylL18JbP4tmSkED4vcjXT5IhyfCFKB61lJscqx
N95d6lXpEZGGMcGHFGMmturMZ4dYSY+nBTSDWaB/ODKtG9rQgqI54/YcZWaZ2MON
vOw2Wj50Fpfh55dO3b40m4zFcNkIoRt5nMEJ1GvMsFQexEZs9WImL6dnE6yDGpV2
Li9yMDV8QJFBkME/C3AVQfT2RoWliadnxeW1useiaxe2k9zQ9TCukWJnz7ZUjFP8
Q82rSuN/TIP8aTEpFvJak8QKV5W3YmKdeFQaxRihMkALQKV0Df3l3SWLbsUbHJHN
P61RCRbU419sUwa/ZTnJjjum4Fk0h/BTfzVRgClaPGLrYDYQ7SB2NDs78Ft41ezu
j4yKOXIucZ1ihySqlCNrK0nYAzAPOlSZBMmCnRY+fcGqvYH/9gtoxxsS19FeiAyc
6NxvIODUdE6uQ0UOP7PGQKLCOJwmvqMpPYICa8ogXhZz1wAsMfAioTgVqHbjZt9x
sNHefYizkIaqflizM1kr1nMySETEbclgSpgh+Jw/40spvHDvRAmKd38D0lDOuZQr
tFBFRPJZ10CdQNJg77a+3yknxZ4o53um8ps3uPzynaJ9+9hTuQfQgJbgHO/wEXhK
fOSVorksNvZ1t9B17ha/E64GivFoP8rtelUDPHWMQLtTHiJLDGh0GsWl4ukBUeIr
3lBpYMIipYFBmOlkYnc/EQ+TDgDdv/D8waL4ctMR+/pjBtKRju0JJ+a8YLpQitkx
nZfXik5y7zUCozAxYYsUFs8pwIldu4dCxd5HsTK/brO7YhRO9rMqUQVpZ9hVUMBp
AgGuXH8de6QhEgnTxHTy6xCatFjJiOQDSH4mwCzRo6mc+r9CeimPz7Nc+1IjY+a6
aUANNekukqPuVwEarba8iGa2zEKKYvEYGQTJrX5iWBhntER1lWSnSDZKmlfKbo9q
m/F+8IZi/IiKJd2Ggj0mCH9sYY3lGA03M5d++PFAGD1eroSUTPQHnkJoKQErWI7a
Ue3VDBViApt0lmMT/fQx6WU1To5Br0WGVJuGsfyS7XnflWZ8EcXXkuAB8iqT88N9
3DPokwAgNdyPNM/HB7gASMJ/+ZTY3J0TwHNs7dt1JP2f2cpB1gm1kXcD1aMS495f
Nlqe4OCKJIebY70fmGdQ5K1k5DjAkIZ1F9w4PiRFjVebFT+FhrbMP3rHVHa91U/7
pdT6mWwX2WyX9KocQjfPpIegZcgft8K39/MTNsLrIR7/55AROKdx0e9L5QlUxzfh
v42v+/cy1T8G3S/d9dIpTt3gupJHbEd61srnSOFXWJCbfiWKS/pmE3gOa0Q3mXNa
CSwBjN4ud60/AURftKXHX4ePH57ZhlBmeHmhcFTPM5jW7KkitX5wXcd6OCMGcL0z
/+dZ5SkTl9o1AQBz5QpPHIk2x+gdAGrx8T7qeeqwFgK/AgJgjbUR9aXnAFAXNVZO
zqUc8o/mb2bik6/r454Iob53ZgJgjRMahdd4jQHB2h5uA84SZyf8AGHe5U3sAKBs
16vAAAiJtfsHTq8rCBRfytTRyAAAbk9bmdjxJvss3BHZa3vCjhK12WDsUX+/KSSh
NTcpvhAS5VIREzfCbmGYYr/NZYFS2V7JChWWqs3W397Ich5g1lcu+zwZp+2eIutN
lxkkIPkr2+LL1jscjYwegJGP3VNdozr7WjSfUkd+s5LG9/35r+d0POtT+Fy1U3jE
3HJGtmLY/L9+IpMX8yH61wUHNDreUm6WZ7BvhBBbDTpLcFZhzilaQb6RltNsJ9ZR
XlSPPBzVY15j5w6BK86mrZrwQ81WarSY2LZFNBbdq+JDDlCqxAyXpXLndTn4lMOb
V23Eae0LqZ9iCvjPlN+5/7V0K1wVhkXKF3ahz+TxFm9TDimeRjqoiTpo+xLwe8IM
0FEjdercexu/JrYyD1Yd8/v8BYY7mm/TzlQA0YMWpg4mP/FPanisvHZdgZBzXnuM
+SkrcgEjsjDHXRv9d3lBlj4b9ZRMoPlAbxpgNtT8gcJV28EHzxKl8RwEIlON1sZA
R0usD3SSs0r7lE4oqrjDkjS9LZrnoj4+JTQSpdMqszkDxx5F2hxBV/hUx63BRcej
NmlF/X5Ctyt/cqbTBVYkQTtwF47HP8VIqXWe1zTb60RM4fNEyMuqGqA2o4xD7PF5
ZLN0T/QPNlWP+aWQuTjwbnQx6No95osJ2qVJPKFXHY7rYnbT0hWmGYIyfCpBeB7W
pKY8Zfkdye6pPYhM7Q8w+J6xBAmiEv3tFszVFdoV5mWN59GdVivjpWtKi6VEAOqd
LcS2MpDfiAAjvhRzU47ia00YtgpD1U6K9sNzZULMju4w5z2I+owl/NB4LagLfpVJ
aB61brvgq3sg9CsniYhPhgQVofIBSFgW0LfEkufBfyW+OCWsCAUjG1jEbipMbTzO
k/CmEUKMAnpLyr2nsPe2ILse9L/q1UL35WKeaMNsZ6UqE0gkQTJDDfFNVs4tkgts
q6tO4cKiLqqgXMor5K4CceLcXDIHYb0S/2dgFk+EwM1XaPw78FQ0QkJGTf6Sg9BB
uYwsa0T+F5qc+F3vJiRr5tyE8+fM3Xz4fXmVcaahEBT4OObGNFkNIMLx9tArBN1Z
25PZNMTKc94ek228y4Dhj4M/6LVtBvbQKbS4Pv5rGAO2fH4qDs3uvHMO6d12k4/T
/Vpfm5ZXdw8s3YhbqdFMXzZc3+v7Pkiby5aGWZpNzn4MynkIV6uEAtEBk1sG0l6i
4w1LWzEj/F7DHZn4Wfh9fdAeimLUVhSF7QHKskrTWFg47sxvua98JUuWikHqGJzM
2L6rmCR8Y1sO1kqzUw/u2jfUjLTlly0cbDc+fYpWRyxBP/yWzYxDLcpr8K7miH/7
FYhQVGAkZA4WP/vW1vlZ7Vt5YpLjJto6rHUYyJKNppJMHm8aQ1jae69GQM4ljr2h
OJaSw6BK7+mzZGVGp+VEO5kuNo9xmYS2BTtJa4mdB+TYaPhhJ5U9M3O2eTwO7nKz
JKYLPtISsWrTKvo0qkGZ3+usd0PuKnYYfJzba+/V95WUBdraPzae/8cvFd8kD3yW
xh7+VK78l7OODTabF/vIQr7u6HX0tUFDkvjk9taIz+2GSmslfC1FwX1rTlS0suf6
EnD5P6MfLy2YkjKBDQREV0ScGL3oHZ6f6LIJ24omy6fjbRgKdsTOhBnmCja7740D
CvSIt/tDqV2FmGaunXMhEUHe6H7o6bjqYSkkeF+B/oPoz6APxioez5/z8jA3FcKp
f8V8f4Uv0LWnkSgRw9XaoubkDMu3CTAmwxwwihCgEe46ji5ywJ2jMPV3zfqeYRej
Qc9V/iGdtWVE8FiKPOaWdRb01yTby/A/BJeauQ/3w1wl7EsuHT5Aezu+6qMM7zzL
3RoJGyguKrwQjR1WNV3NVMWTdcbiZnNtMbSToJB53ZhqAJ5YCsaTlOyrBcdAvPP4
qBcA68hdJOSGVrXnLPgvQE3cg1pXSAkh/GDUouDi+eQ3EFbOzO/TR7JpeYlHsnBB
GmV6ftaQ8VS4Q0AQIrdP+IEDtL8WfrjkS9AYmM1KVlxeSsdfjl6gWx5T5NR6zgCW
GCbvfR2qkQSDvebN8XQrCknePQ42gHs4LUfILU96+8qOKIOefyX1yF+XcAYS7h1g
JsvYvbUbgQ6dgSDPpcsi07WMb+DL066H8GlnOprNXIn0DCOssDm7Q11asOgJ/Col
VC9kYFlX6G0TvR2UWeavPjTKDlWE+8rzTYvdxyM9X2sTP20vhb6lJ/YLYabDtHEy
yHxW0RQ7r1IN/VQuZdKoDmp9tIMJJCCGuE9w1CkKmEL5ROc9oosixiJ1qBMrbrc7
7BoLahIUN6qZ5Jay+8pMZOeH3ZrK7YXXSsGE82vBoE9uDFK1C2r5KSdIaWBpprYx
4ja7mRKIdeLIpu9ZOfmKZiRUu8IKJUwAi2UrttAieWUw8atocPhIflE+ciYlpP7p
zn5dU3dNfUfv7Ok97OxP+mF1vI4bWOqt3bTWq0iB7KJemjf2YjjpV7w71Ph1UtaN
CDybQ8soTnRdHPKcNjJTMqlI+nkyGYyK7eyyjPp7mjhqpXGANo4EW0F2W/USnxQ7
UfsE0NVcY3o2tDdBmgXWeZR7IecKGB/0pv11gcsCOQxJ6RBrY0v/DSNMQi5N2LSR
KjJgbkYsHo443Yg5kFoev6L65GfIuavpY47yvr36aTYjZ5O2XPes9Qvzo8VEVuZV
5riTKvSq3Tb/9a7Yj76D4vDOaLRt76I6qoFBZl52hiP5oIPigDTEKSulBPnLXFcX
ssAveZ89pp8tncKkkoOIwQDb2QZQlTuO8xpBCfnI2elNKMFiYd3YClAMOSioCduc
SeBTSJkqjA98aPbi3mVR/tqY0rZndOiE/4fYgxBBa3n2F1yeM9vNTCH/K9qq/V5l
np/VoWqWYwBYbvpVyVgPv4QVeS/1444CnybQeXEBFUVslAZ1PKR/maS5jK3qaCKK
a5wKi4Dt0tdZlpQrMXCjiArj1Jn1lt48y9aDXrW/sGkc+Ku23df/tN+/T2CiSb7O
mhgmoTtenM0R94IGMd+tm6Gr/iwpRu8VD0ar3p9i4aQiD37eVPibtaJz8NU8DxDj
vJsGBYuaDx0jwDrL6/9LC0qGu1Eqd6geNqMn94JgGEOipId4gdX1NQVx3c9ij8rI
wWuEGisGGcR9/u3L/BSvG8EDawF/DQlNX50kjPNCDN8s682/myPPI5fizNVwmEiT
K/YomGvzGQ4mjzk24vEnqgXjGg2gY+m9pETAEkMwPdO04K6rgaM5eP7oLuunDuKd
XLncuBYrxBiqf6b01bc/xRE7YoVAdy7JnX6vcd7S5B0PAayUjlL5ib5q0oRlGm1i
tTHZMBKz+cP4DiwXuSMGmPEQZoBrId/YsTVcGDIjagZJZh4pMUrS69PuN0llNXjw
DR14og+t8Cgj4YgGJbpRS2K35ksjHn534sekW5G3wBgcxs5CgynkwBA/T+xSFBYV
1Dh0T6haRfDHQmgf/MESAFzD/HdQWTQrYs0Al++7QHxazdn4DShstyfCMNhhGjM6
EiRIvjnfkegF3zulCZQhn5wgzSneLu7zAH1pTfeTQFXNRzZAWVETLqeMB5xEqZD1
Oi0uBLUO1RMGQ7gK5DTWdPCfltO6J0NlDtLu3HEOeGgA9Agh4wNCy5jtLTsQS8wD
97j4ZWbwUhLPGzGFu4iKELqBW2EuK2JkbmyTFUfhWAfglya14odgPKxFGby5zEXr
LZb+sL+m9YY0GF5WPEwHBmLC7xGih6xk2VEcoS+bffcQyb/5H0u/QFsTBpBKGOaU
MArJCZnQ8Pt9WG2cpImPNcOjVv0T1+pev/ecFVw1XuyfnTghv3yD/kpC79BNy72o
vWIFs7eXLSFKTsfr6GWDBK8cwS/5ecsXoziHLccH0cSDch+8ydimyokUkNV3be0y
Fw5ZtQG2u+FUAA6b2yE2oGGA76LF/0V8GXfdITU74YjrlNkzhdmBMLRiI7bR8jeS
3/0rG4W3VH5HUU8h1fdzL8sInHxevamKFlIVLXxJJs/ILw5+lzKQdyNoA8svDWwU
NAcYgNDx40tafzCPPANKRaQHUXWVbRw7ciiKBZFDm57hoIGyVxctO8Az7dzD1yGz
Z6o+zcgg0CBVS/fiISTlHkM8YtvVHdrNPAKRLShQVwkWKzCf1ealwhhtuZ1YnjH9
WCJZ4DCebmnJKohoRRS83enGQtC6giNBzC2g65guxyQV5rHUhGZ4Z1eRdIJFoxWZ
S2Luuz2u/2pbn1+dZw2cmIO5VLbaNR7PAjc76scWXpGMp5PVZxXXxfh5tLQ2XFwz
hfQL5+o2v+t9sMwEcOwclE4ZCUeVv1vaaTiTFhbnsKfHcVvF1Lcn5B+yCvowJQ2o
xcqKLZsLoNdB3qTZ2ZmJ0WXyZaWcQwju8eE/Sp4KPfXUxSXqJhxgvk9NE5bPvKiC
7vP0LZgYg9iHC14r9t3w1z56j0dxxu3Jtl4jRPtmS0MFUF/AoZDTM2cCFizYckma
OugGQKm1iPwcf+Tn7fWUjMJCvQDIFFYFGUHBj59ntY4dd/8av2QMNt8um5zff6Cz
gbTVIL2/mfodk0EnFn9vwgsaRocUOPmoP/uX6aKRSvDbYv/77F02WNtyfZVtYMvD
vJtVmlX11amM/JoOPQzmcMXOZNF/9+MHbnDqedbjlBCv6pD4khRRQAm+RyFzze85
J0a6oyrRJtp0VVurl9baBse9MARBnreVBmYt8T4cW1FIkOr/byf22bAA4kGZJcrP
GCdI0NPnCggM/3tClJTSe4xJzQXHJVi7I/Ub2+f85bkLGBZoMISWTrhlzoF26BsC
NUI+6FFmv6YZsd7et8Vxyf2eE8sWgCHVavCDRSYQcC+pcsvZ3UxNRbclxeY4NLEm
VlJo7KWEv0BxfnS9P5miVSBBv4uns9lkfOVcyNKz7U3YSppgh4o7kw0hxVffLjiC
qAuskJ/C51OTvBo5MpeA1rExUyP8TVuTFiWT5i8i5pzXqwsu84CQ0wjse9cEwYzV
0Go7/I9gLpDO3gdYQVkTh+N2zMu8H6xQ3qz2yv61PDsDIKwyVr5U6aQZGsTO9v6x
9E9aN5hHipBDShQDS+ye/XHUfkR3+51I5OxGCvOokbmJjNivJV76nPP1TO8BDDuu
6ErTV/MIEWXxJ/8kOU+WtKfSIFFOFhGQCBG+iwh4wJlWRXP7VX+A7Wgo3boeEk6I
zVWABtNBPZdBDg50MnYhdZiU2Apijuq50smmmP3mS67wKMmc9JYcpmhRkTtX3zV1
j8Zq+V+NPzHdVLamHs0QW1wNLmW3VsSwzpH61Jzw/gWnCLwl8oDYxGXQ83CYI+aM
K18EAhfFT4eS4hnnNk1mMgzo9JFUtA2JzIDm4tD/JOf/k/yrJCjGzbzuSCWmcL1O
y9oxJZoXVN15vcRz4Vlhb5AqBVKpBiXrzbF8h3JBwi7rsAUN5rdk/s6jMK4e8ELy
mB1Btwqv0U2pM+T/urg/t+Z5fjwRuoej2yr8yB08S/3bZHGNCLE8YHJWd6ZGNq4W
7LNLj/XPq8dqUBPy8TaV73OnIAufflK1eP3zQZI3VgkAtF/AHHWpU4okilzCh2ri
HWgdKoFRcn4/0Ki08Cs+S8svCMJDc71vMmduN4lHTpLnfEwe5jU8cS6VRy/uHq5i
0YmSXwh31SrDvz8RilhZEBenoLK4Gc2/iX/U0e/IFTFkndy6WwsoruhKkhSjYcmQ
9o6z3tjY6Fi+iexHth1jEgR10TvapqxPEOIFAjfhIohfylBEM0iNlUsqtSi+8BPx
xAHnYpIYOn38qBkQDtj0A22Cza6i1B6bR8exIPyvHHVwynuJddF8NmvUOfdBKS+q
fIDbA+Eg5rs/ETxPfBomfvZhxLFPuEGx1hY+knhqiPSa5/4OzEuaeMENtWhcQ8M5
FgJpOqrVXW5J/j/nelFVpznlS89QK02rMZ6IBwdDjGxhRw5CkfVp0usjZv1nmFWs
FMl7QyqNukmHXzwAhjVj6kwN0T+gC49eNv16gcAmx+FcnS31g7S0Nwyt2FQpO8by
K+3ivjzbEEDc5vmMlfd/ANehOFAOjtzSHTvtcE3Q9B7X51f5hLZkwWZcEEeSP5il
xBfrwXBb+8KJe2jF5g9s1rrAmlHcCFN3Gx8rOOMH59eWufE864o5/L2k8WwCAARW
j9QyjOGeC6FjBfP2oxSZD1A8klAwp8u2gp9fb9MeD+6K8yQ9vCfwPBwSIWO+IOcb
aNcys8kWPDqBChg1AJTsYJcZ9inTcYvJvw25p2t6QLgtl5itT+LKm+1rR+P3gstQ
Os0C+istGFHv8jUMgI+HbDOoL/UWR/oUAS6wr8EjdYq3SINveN2FvP46DPChQ4hx
r4NiJYeep+g27na8mj+UclYviKFLEzxCAU785sb3SRvFw9D8TXFvoteZWb3TIptI
3QZNJWPiAXDLCNBynuxvgTzO8TB4B7IO+sYGTzKmU3BaKikueAVDXey39fgqqziR
z75et0wV2MR0aUXcs6Z2s9hr+wxDbBRa2jbn3DsnRtTDSZVdQlx7qSpmEzp9HJLe
K6bO43sF2mH6gyzv+jFHtIWNsImGMzhnjHErdaovPKusLIoVmwC3EmAAEdFtTcuo
7OXPhqIfFq+29L4cCHaOEF8FAGm40rpuD4NHuWfSPksicdBM/3EikF26ieFbmH38
wNlt0JuojoWxqZhOKH8f0F4csrdlIzFUSqOub+KZioGH0NEjPSSBYjJ6QWCKaXR/
DwBG7rgbJWksYaLvE9VOFBuzjGvD7DSeueRcRNqZcWLiozhdadpXWnucfdaQ/TC2
L6zFdSWskQS3aZcqf2A+oCjTPJhJ0cB+ZcT7g6MfR3qWUi2bMRVB1pqcV4qfBI9I
akMH/li4HT7jnZ2PTQWLupaffCI7ue92Y6PLO/ZYG51gMH4c5vXg7mSJ95iCIwHO
tvuagYFg9DH3o0+bbx0mHyw2Mf1eg3DWn72Tcjv2tFirBJXjYIF2Sb/kzuRirTON
GnYoKWSaW3Ph7/wuIr0d5D8p9GpXEHYQ3FeFQPzLhlN0tJZZaUZK9Bpb1lHlQglK
xP3nDDi0Sidk8m8BbpY9pbVdS5tTC5Y3UYCNlRxyRy2bE76ly5raj9+uxvqYN3BT
1gEHcbaOQdZJ8Ik9GX+/oZboSZXNy9TDS5U3/wnwtiJWxn/ky3Yz+2lJspDvpoVg
30U+1GqhQmZK36N6kdMX7eaF1B4PWhQPsC09SZQ1/rQlRFzzxrtGpdPwzEzqyVLM
B5XXa/VsUeRrN89xJmkZw/4Amj7QpdMLQOFqS42UnkLR1v3ig7mzkDT5HXNZ1/OV
T8Vsb499d/3NGMq0ust+7KEli7efx/dF0MsTaGmAAnmxEttbBQKRwQ40mRcC28ZR
uBnyGkk+AIP5gOqxiH//rKXi85haQKBuaAkqrwiygN3QUyktzAEB30mHN2Di3F1E
PTbFXacts1oF2BFOEqYaQupvQlyGbby2novYCHp/MkChurc2QX438HFofIhELEjE
s4BVoXguAU8nRSAVs3Uvd0pv6eBlSFnj1OPmPMnOLNNia8EwBY9GCrOPCpEcJmgI
2fgS084kC8tk0uou5dqkueM3guEt6iO6gSCUQ3qUOLonKhELX8idr+T4UXgS4g/H
Z97a1jWwkmQJVl/kLJFbYGRdGmLfUHHCtVnUjc9RSDVmnRjJUzZ10Q77glff8PK0
9Q3bvIKcGhSGgKT518QY/Ryiy9AmQgXFPOjrEvGkiNncND2D0XI2861F8rLDVXUR
wO+q9m5x5ZgcYuD/7sOUGzBDJuqmxym8IP6rIl9s2r4AGed/WV2Ri1ZcJ2j+DkHk
YAfvafxGNE9Cxnww2xC51KRgpU/xX9Th5EKJy17QZ/D3xMvEaN32EoHQnksYALvo
iDby8WN/GBROFhaVyWb8iOLyeqINDD4hv70ZazSDphAgOBnOl5Z06c5+Q9p5lvQG
ZN7eUblIWTTNcNYVAS9Ju51I/WrIXG2xRuk0hrmIKT5NSLgvKsUZ9jHvCUr5HGpc
XQgucxho7a2FnXOnSDDUNrk9wBdS8F94mmeoUS7SnnPV9kuChFGMfhw+/7XeH6Hb
VkU2+xgr9l3VNPK0uvcdY5826w/1N7mlxNVLVP2uvO7MIdTaNFXyomLiV1ZxK+OI
setXlmpXY88MivitLfttVBfqY3b1amNzqZtolOzdZmanwe/LHuV3QVCJbSDANtVZ
6HG5ow3Fb8x37w6Jk47nRRYDFpZW3YnTrc4H3YyH2arjG6jUAaLMQABhbAaw72yE
GdlVHnQLiC/zXTRoRTlqcbWboQKY67B0g57SUHAgufHoyoyPp4bKDXhpWdMA9hdg
p83zGKeXwtBQcQIUQhBT3AtST9e0gm98guZoN5TouhrO18J4swBzYVfbrGAauNpT
0kdxKZCK09+YkMb4j244ZPlk6dOk66X3RFFuhs06h8jjD1Qj9Nhx4O6YXtHSAr69
snONQ4+5Mp1Ew56bkA/AevaV0eG4ndGO1FTYoxULMYt+xMdyGYxjrIcuJhswGY8Y
XEqett1Q6IKIV4GrPBa3pDpyNJfRMRe6tLa3ZODiq8YR0eJOMc6hajari91HDKw7
LRZI8Go9nYl4+N/AuYnwaZH/yzsYtybxI2I9/L7+2NLTAXRTBQ/wPywCuaf3s13d
hpSHNg47rrevjztykIuMi/Kb5oX+DHaNiq3gRCnmcZg0wRhKoZ8Ssdxn8zl1M/iy
K4aPglmSdEo+g/W9jdLhXsT/gUa9oJG/lxGl/OtKiphXRfQ7OlvdY5EPUX3rTB26
PdsgqhKDw2UQJJmYnAKpShG2o4yHglBdF2C7Gjc4rpSLlYa7EfSbmQ+KsTu5CBnM
4396Tz/oCOA2xunyJVymsavRBNZt04VSUZnT1Sjvpo9ubZam8eeA6PrRXQwD5G28
px/Jb/sxI2AcYnCW+FJ1HILnpyYi47Iw0VyIUqrBOOSRezvyCkGpgnSjTX0mMYWZ
hJRbXB2ldnDbOn2bhKyuStUr2Kjkf0PszepWa/EsHp2EC95+P4DswXNewM3/MZtm
RkofTyP2Es/gNKAq2SO/gsVfBgjL2JCqkT69+OwM0G12oX+iotJa+KrMamwr5JbZ
CVST7BNM7z0eChoOfDwqfFjpdxYpen2z8y7nFVZDh+RWnaI6S7P8z8wImoDONTYh
k/mUTmr2NzD03CxLMsw1GSv2sjrd6rMTHgboCHoAZo6FXgh5KW3xzlQx45cVAQZp
cGByDq5ElBWI2re+GtBu8gvlFYUmQQAxYkO+hDSWfTk7coHUoPwkWpQRGfk4F1Xv
LtrwASk49F+HqIpmCzBQP0TYT7mkNV05c/f2NZPJuLuOmXrxwu+ic7uJSw1/45ZJ
l8bGEm4uSiSpx6G3KX4MBXhXzZKZKlgAcW3V0RGo1nxyYYJoFt7NAkwIsWQgfBWL
O0PeGgFHIS1Jw/hCVwZ0YIb10EVT0iLeEHcADHm7MUhDIOQcEOTswVM1RB/IZgp2
FV73H2ilccL0ax0Ijs8kmf84UrSMIrahgIFzAjTaO0QvJpgCzwFbG/NT2Jb1wjMm
GOzkexuuHc49lckrBJaon3rP7cJv5Dukg49IMsGuPka2SMNmIwx2XqAmgs/1A9iR
xsdE5105iFVKD+V3R2Z1icz9pSua5kuKos4IUo1EB5UnefpEIgGfZp+ICMRaYgmN
+2sPlWxOXI918IwSdEEa97XTuOL5UFci7F/ezr6cBIfOw3eKK41pNTFXnc6ZPizz
OWdRkrRzC5aPyyQoiV1A39tbJNSpQV9fxyXcik5zDN7pqoh5DsepihHteCmSQcGA
YDHvRsSIRBv78dKZJoZjblvBGl7Ooiz2vB6vlInOmAPCm4tKLSGsdT6AHRNK4Lr1
oUuEHCsAxDtrb9LP/Czwgg8KnGv2xTPR/HGGNKmf8stnlpbgBGeHGyfa23ZEQi1B
54sBifDSwD/f6j9W+mOrdMBqHSo/JWD7a0ua9CM+mLQ88uNjsn3ElD/G0d3wrW42
GVQwkHlX8uJSLips+ijs8gtY2O5la1ecT/aIW2rwVaEjdJ8KsC1AxsV+aJWNGou2
L9wNhgspFSsmX9iD7Qhvjy4bYNkk08BdI4EwgJ2mu78rANEBkn+uZRhZcOlebqrV
BLRDmj8KX5OXvfRdOK/xrsCVdBc2WFh46hNvWwkb9ZrcwoXW2uZTbZ9RS7+n1r7d
Om3IQOdXTiZBbMSMft1zO76JXsO/3Z5V9QdRgdg7WrZMjfgP3f5Z52FzzC86SqsA
3rlf6lTK+/13q3mDPLfL7Cuk2zzOqb/7vwuN2xwTnAaptH4fU9J9vsEwKy8hXxVX
e4XbBI97MEN4TPmYNBTXrcmCm03MmnPQdi/G1na6+OvtmEIdau1dkX10N/NioD5J
OUf+hxJ4olPj92Od09VHkIvV/J6c5BxGgqkrFDxyRTwx0F/1I1OayUoiq8tSQ0jf
TwGLhA2dscUzgPJzFzkqPXLMLZBVB2ohxyq+iRAitcDwVbfl2u+gZegd7quGxNzY
hKtuhEK1hlHLZgvcYP91KzkKX4o/Xq64aDTGalmPY2xOJbs63+FCn5+Uyp6w33Up
CI7LC+w9n0qfES/mYkEgEv5En8EDOeZBnJM3eS3ZcRLQUcC0Iiqs/T+EUNE9wgkA
10EJWFCtb9GeEbIHqC7vM+gGYNSvgM2tbXvKmoYeFtM6vnN8ZNosqjFaCvPqPVL/
lYfEeJkZW6ZYVxMSx62MeiYljAwIs/i99fdWwXYe8yny5BBRIjaLO9xkuuGtgUKu
fFr9HK+QQe7a9y88hYGWDIZpJLXHjoLVW9yJlSAzn8Do/7fhGCbOTPw+/8Bcss3A
7ra7WKfcBC/cywedFxQ0AFWIgHIAJ4Ln4iYezB+xVdduHZxbmfBtPZk7Qn5uDKcw
sihdc8IMDhM5kJ4/jcJW7P31G5bp7QU6iRO17AeQjr25B/XQwZEGK1A+Xhw8eFqc
YnfXKhymak8tf4Tn/+jkrwmBYyhoGMUmgDi+vu577bDxQJJWoP47fn6pKNxIve7v
RQi+3ds9cRMS8u9UyYvY/kymCO17FJ3F5nri43GtL9pVYu+kitNOJY1KG/IvAgNx
OZzRenjyka+uStpCU7gRPWTR8FVvm7cW54gHiIeVXPc4evg6gyCfaZRfsSSypxto
+h1+HhT+se/cLo5P44U/wuxol+ucQS/J1Xau/WDIsuhmZ7dbmFwf4odY8BoRLmEP
oqEQPZXERPamcO/9CoIwh10jY23hzhbTJ9PXFH+fv+8uapZ0XWGpNEJXOxqrNlOC
3CjdMUNXOizQqQwtGQcnBQfgLSkEL8BmXaR0mKn6BN86NzLt4oqgtLgD2623lxuY
llm3weodmGEJWXTTWFqR7n7mYp48S7nRGFXno9Mjr1H4DN6GIs4dxOXzS48QSRjY
G5cWw90TIAL4+4c4wOn/0Kl85djerPbqVkvB/je8AC404BOJxDKv+LxB3Cpka7Io
yaT5qznAPjelwg6lnTob/0arBHp9hggDxdOI//0HkcP3ZyFtRD3fMnmj8EKHTvq0
QTc9N9/g2BCR38R+lPmrUjGSAvObGx6UvBVJiLWvVDQfo7snBK7L+w4x66qO3Kpr
B36LnCCZ5IJLAKjSZqhgAQinD4X4zyEDwTgO9c5tu7FAaoaOKU66lrAvfNt8kwWk
499sTOa9nbYuyVfT3b2U84y9h6Phta3pcO9Qi5DLWuCRhDDx5wsLFwwRy9pleUzf
9aM6Hhn5TKGTtB6jlez1vcfsR0B5lKUlQgqhoJO/kM8S+K+Iu4C4FXxs0QEN3uLT
Rnvw0dA2UrI6L6Z82WUNlXXwGkgjUsok14JqvbPwelQm4zrlJlGKSAe/9xHhMQ/c
gJTmFF2An5L3Twrt1dy93yEIpmZjN8LIQ6fXq3b4TSnmRHtMCgogKkiflQ+bG6fU
oY1xFSY04tzTAmo/dERnw5ylmQtq2OND6h8RosewY76VaT8ueDxBiWVAVUzbhEbn
yCWp3cOj92SfyYYRkYOfx7qOJVRSZtpLh+8tZKLrvJrYHohdCHXx2zqKUx0FFyFa
RO6vCu1lPcssX3lmLyFSZegWcYWP2iMNequ0wkgz4MWiE8m9IYh+KborE33Kkn5W
IYapSNtISbncFpVb4U61a4hWKRkAw7c+ijQy3ztFVlcegMtlTILvjVlmYUxGEIEL
4zCPD5B0bvtjlyDsIO/TzrVW7X08vEl9r3Dj6ph5oEhhcUqtEQowkCn9XuJYET6s
Xd7rK1Rgcb9OwzzpXHTy6Nd/vBxx3ReKH4BJ+wpWZIo8DcbrNI/oZhC291YmB1MK
fLk6i98gstuyF52TTYt25T5DzoSktxQXXvwhe+EcbMhSm+a2YrCBSl1yCSXJFkF4
j3mcWZcQViT8t9f+YN4Sl3OUI0V4HusEUUX+Ew8vI0Ak7w+I8MnabA37MStNdMT4
twU/S1qzH87c8/F0ttAcHpNqlF+DA7gdSMxgWhdmVaUAk4T2ZxgMUhoa9wCw4fvW
aOunu3o75hs1DDlT3wv34iTxT0CzNf946SNf0cSSNHckUhyOEOj8ex2Y9suzJOs+
rF2en1sc1B6j3wKbLhoIEKIcxubfm2aWx7a/IVbhBvHkcEuqrjjggxrFc1chirED
GEwyTZsEdVw/w6jBoxn36Wfot0z78qc18rg9ryaSFnjhLRgekn1OZbEJAsOAPyGi
Upxa0CT/DAl4oMzi9OGZPELpVGB7mt2HLicW4s+tDs1N8odfE6tpTx+3XAs0m8fZ
F2TgyficaQ7w/n9JrUsDi74WqAX9K6LNaBCrBQk4ysMySDxeUaRBY31Ik+3fOBw1
5s8CHfDFZoInbbmE4Lk4assF6KnUHLMBrjkNuCBZKAy7AELCmwkzaITmmRXiODLp
O7mRU+zBWdVn73YBuv41YeCrrQjI9Wxb+C3pX2gvWK/MO333rVUmunYcortbLegD
iojEptLl46PI5FYtQ4oT8iPeTz364tTMTcGmwfKDyYGsNf0dLr1it2XarmOrDqgq
N3nbn2cN46urWOsFZCfH+s0612KWirB9uWwTBmpjk9XE109GNyyiPhCEMrXz7VFX
9+uF8xi5a/JpkNmiHDmrPCmfrJIPfNjGxYFKK08VzIJ+3o9H7uCMzqmBULHKBWVT
3KZ1IGekIHzqczN6oNNw5L6XjF32C2Ke4fkFBZeardbHBj0+KXfgTMnwZw7X3gB3
JvjXL6kWxh8jwNPnLGZeYxLTcOl+rNVqqjmqoWQHOvtFH5+tqy+HUO05C0DXMLvv
GbwUaCKK+FCuFfJ8O6man0bKh3pCZRkbzKxmPkNG+zOmFFVlTmfJq/Z0h/7zOXrB
uYkF1SHLItDmit/4k63JvUqiXAY3+Kl8ua8caB3JFOaK4uSMdoFUv5qXC1cXQZbL
1ea9I8YTYS+Y1dAhgkR7CrDTmhvhgWP1gdZsidzma4Bjn5PRmmIPFP/XuW5HIf+3
qE1e5YGxWH/cqL5W+YM7jdnjGpghZLrmADD7bAT+IkbmuVOiVCSIV3asv8dm8KsM
SuZfvhLyr78yP8P2j2r0TzueXZnMErB15FVLFl6RoDx1tE69xdUqdvbqGKERR0tm
PMKvQZg6y+g5QLNJa6ojlilD9dyTLNS571wH7GEURmmjhNFVwTWd/4zf/o/E1sVJ
6C43+ipFHa2NZKvtDIvIQvDxr/CLC7wdDHIk913fLQEXRsXjobrPCbpioOgrn8eZ
Le4AbgVPYV6ckUahzFYC5ZCu3NOn5W6eiEMlL+JK0UgCm9iHEIYL21BtRpKSXnYY
9zppvn/e+ErZJkJ95jRjCHZ84kfFYHfLVq6GyzHMegK/wQIyOtY73dfVgNYcNyg0
82I35WDGsqI4TAFqst1FM81r64gO+q2+DnctC9hvNC7MXGg0HzL9qlXYNyiSj3u1
bnCmITvzqJ9L2WHMIcan/om+IK7QjLBEakkujzlKdZmzYUEPrUgVsfMu032xjb1e
g70ioAxR+M7tfn6fVePprthrC7FPDWZCQ6h5t1HOldBGBThkmlN/Yk9ugEUViZgi
yK9jOxvr4z2qeGOIyKxCGE8HQWGA25HiHNN8V7SY3K84Yh2o9MHyV3AiNa1SG1gk
xhkdGL3BQfb+IIbumR3PHqHGw+tXQF4ywqQLOIV37+NZCMwuoCY+dc/2cHomfhwK
f2P0d/Li05WT07rcRE7lmmOFJxh/nTQ/aWiY0Tl+yn6LvpJMpijf4l+JQFKd2uUL
BK8plgD9el/lfxmlLR6jKdOm+Zi6wQSBMgT19f3F8QwmypbzTaYZ02mQp2+kSHlK
NBqqK8JuVAUrryTWIOzm2GyKRuzeinli4F73F/6b3nZdHy/ElPmjcREmB0MXw1T+
jY5SPIMbNZsaAFVqQUZkR3UM448g747Ijq/9AgUGD6Lohy1oaM8jj8ItZ7zlCAVO
yN6d9d4k0i6v50XqpIC8AOq4TJ7fyrfXnzxYceutnVKkqufraJnoI60MIWsECnmr
xbw06svmkYRKKdzaLg6+LLEFq/0Hxc4+1zBtGZ+hD9lPqx+V+Qct6cpcd2z+o7bG
nVO18DEuwiZlHl5gbW8voVwnkpPghd5hs4PRu0ILHXj6FdLxrxqjk2YnkEpN4NS+
IKbiMXLKfh7MPecvo6Ugq5KoVsc6NalmM97pI/a541Sd2ZntXFDsoC38wiYrnMD7
/SOfPXUr+iXTbRp+7GyNSoxsDmSmPZu6G5vkKapdTwgMxTJ62gfdrjECafqh2WGA
/AsEZ1tmidGXhXBdG3O861rn4cBp/zCPncGzmbWAXggEHF/HsjZ3wK+RhVBUMk2E
+OpNTKc5daXZAPo4hEWoAvwqie7bWvfXMO2cpWAF77BzrpFZ2pMNQJvlqBd7HOaX
2/Xrh9pddcyUeJPkygalUZTbCbbasgEJoEBynUVSX7sHKi1YJtsxZC37iWDnChTi
zO+JDavbzWvDIph+H/CcDOQXq4zScDPsBJ3qVdzfu1w1XKHaNMxhphO6t0GZiujU
7f60nEdJND03hf8WJmxE9fgG8Gx/NkGA488RtP22YGefYxtbFY/CIDJOMpTatJlt
/cv18YMxtzYKWA3GBiA380Svkn3Yve7KqdtahWj/KVNuyKhYqZBhEihEhalfVrvg
Ng1h4MoW3mXB/dmyv8sghACsPigRUzRHCskH/KNPZX3UNJZE/GEtI0fKA5mGCG4w
Q/8JwtHvLy5wf0jsNhq9TRhCWtmKhz8Hgn2UgI/BT/sEaV00bQzlaKzw3ti/WWxi
45/DvTyVK7r0/7dQfsLpvUB7KQ96AZdRT0gdLAeegBpp8SqfuPnAevqegoKz4Cen
IuOiJ4neN0eUyNaQZ7UG71lWlFgLDKvXznXo/XnJoRWXDukJ6ERoICIim567XDH3
1sALd2hRv/mDTzW/jzgzlkkBrTccJoEG8j5yi50dBdz2pZrRRuOKg2krhBfo92Zp
WnvHydDKybNpq7mimW/Gr/alEuC3ehqB5d5yN85XmnAECTjOCnVWwKlbPM5SM64b
1RAWIsAH5Caqv5LRsUnmFXdoRJKUtmFA3Pv5Q3/mhTI4xXTjv4NRlEvoT6lqYMQY
m4EiTPFb8AtBgz5n0GncmMKVXprfqXyl7YmBvnXg70rpIq9HU8g2c75PvUppuSCU
jxqcGo6q1x/QMwde8JuMPYmELVxzPsqZHGFbFKQo7YKA4APOo7KsyMAyr8sv7Scd
3mLT6ns+e0Jx5l1pZWCFqXH94BUC2TR8QrUXVYDDJF0aUvXfFIehuDPVnnBt0a3a
8+QHv8jX/gSg9qyeDTaveixQt1eOY7vw0wqaSwnbHThSlGaghjkHXBYOD79uMzUs
Gkems9Itr5ZKqXeeIvS+R9YGZVKp+h8syxfIqrfsdXD/6oKb5U8Jps0tY511+q31
2Ika9poI+GUWFbVfpcuMb3SKZQR3BO5bHJJ25OQZEXQlWywGsvJo1Py6R1D9NtwY
2h6YErzCpeoRx+xXZv1zIanvU+PZnwL8025BCMqBM4sLvRUvrfI16c56EIEGkjU+
dodCgoKtNTQXoYSsLcXF/lLbhXxUq9lIc+snGRxPeyQwWW0K7vBwfCB/5H9eZHcF
kLN1bWe1vLDBPdtKQbkf9o0cOeNR7LGDwg2SlVdbraIbZv7wMYQSgucUynV2ZU+1
dFgAaiV7wsd35RHBnL+/9iPDufMD67JRtU3JMj8jEEPxE3Dh5uInPfYfmOQ0S/Pr
6fHJVpMjMUB7DsfoJdSCe47LBfqaRd+vk3izPdpbAJiCPFNySz5iYFgDU4Vh8RHi
KaIfTE7crlWu7kDkx7jS0qddsprn6mFcjG6Ht9sBjkqlSHVYrvskubphYFJH5AZ8
pOPwgCaNqitwciK/wUVW+OuUJ5R+sRJi+UR6Mkq6aWIQUaWVB97/PrzWZayJ5uA+
OZs8wXnnYoFYsJrWlKOk5VtBmPMlVWJHsRn9U6um0P8z5MiK+Aur4Jg9zk4dlz+0
dHDSxBk+gnEo5c4iBJD1Ntx/NluDNpH83eR0KtKnKbmSAibZBpndBtLpwMdP8jww
5OeGH6XV5rcWDNOInP3g4bqIh0jN0sR3Si0vZUnCX20PDKaNBTD/spynJtUTSbYT
pd2iXrETYINGUZYnL9jSH5HVt4XWe0+97Yg3bADIXx/ODLhjcLRipDwWezga8Jxq
Rce8+3IWaQVHzQZbdzf33Y2j9whrQd2PQaIUyIt/Z4tbWLGd4lFCHZQXWfgnAuoQ
VS83KmTNdtSgGx4K3wd3/DsHWbigl/H3HF9CQ3MPm1TuqOmvXp/OYvqP+DUCQDin
baJJ8wGHeClARTh/YC+h09uU1l+lYPfi5rStecwG423xiO+LpO2lcphyxNhYYfYw
TKnDQxP62tqP3GOxD76JNsIlNTtEFa8W9plv/COuNLIaIFyTz/fh10u0BywoET2T
TTl7kaoFuWdroSv9hKXb9Nr5/ohgCTRK7O8xgJiJvBFrHiI75e1wyRFH9NBuEf51
jgVO0nrGQcESWAnE1zwBXUwi5Exbso8rtASjcVzxo81tzZmtbJZFdv9e4Swfc0Pr
UuE3eYMmuelIl43zZJk4jgCH/oEpK/ouEPlXbWaNvnm4aavgW3kY42Zx1yvWsFLH
adn2onR+PG38Uh0PRFmJvi4vOxsILS+7ZxC1aJw5g0Budctc4VV39bnThdkHsYob
uj92HSkyEbthBhl/ODJbdGD0wOWCOC3mK7jS9DRvS5cafeHQPZa/Y1mZg81gaT30
115m7oKtCig/2m1TdL+67X0U0IEPrhIogjEsYP/OY9uma8RAs/xcFQax8VhND7Jb
LEWb7ljRaqIDj/OI9SdV6dCYFKFOGNsTJo6Le3/d9HlQ0yC/F1mPlPIEQWNoHAWq
C8Kyu+/ESCyw8W5+wSM0tRfNLhnxGO4F9BjflYw2qHjYVUU6OUvFPTuuyO5XlDKY
fwjO5PDC2GMiUTI66UH1e0aPhejauQYxNXUOAjW5LOGh1S18BrWayr9FOPVVH2Jr
dn7K5xonhC7CvgH4lSRicAPZPtWdrBiYTC70JDheTaF0gd6sopCzS7OTiN0Fd6ib
UoCPMsKX3lYUsmB71mNkvGztCGPAQICfLWZxbmctDDIAkkU4WAkFT+bFdAPO5uHw
m9gL/kllN7zJ3qZbJRBSWo74MPdT2SUS8wOhkOysrYgZIc+BKFVWKVm3i9pqA0wA
CEAI54jSFBdCaQGelDVs7k/XuV3gNvhRfGdv6zINqDp9Lk1Dz+uaNrb0poRBnseF
rvnOJGzMGwBNmPDbivTBg04Sye/DXiJ+UWCM74kJNJCRMD7oulnbazl40epQvE3s
jbQHlO99fuTT1b22PBL6H053nNfxIsWp15Gy+Rs+bOXWU04uXrT8f29xxnLrYTRr
/tzsFZdtcItXY2NIU91QD2PBhKwT94BMALcsieQer55nSLc+ovinWz6L5BqF6IiY
PILEIKN+id+HkfsR1sZJ0/QMMsdh6wW2k2VT+SXCpaQxEswyFVdE5JKixZF7xhZo
ifV5u9sVvpcaoYylR1OYLUn3fCvBdlTi1+BoUuhOt8hCJLRD0FFAjT9pxjLP2QH3
9SvI9BER99IhIXarBT8b+exG0oR+qju9KAP6ha3PtMkaHK47RC2ozcS2dihzKB6E
e8aX6Z/Bo71bfvGnaxcuh8rjBQg16WTccApEG4Oc+akFJoASR7Htf08sBj4KHuis
VLGeGfnXav1d3jnLdTvegPoFItwAd/kRffr0sVQp4eBKqMK5b4PMybQWsO2bwzqT
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Qf9fszyZbsBmcg+2V1wXzxj1UER73Dirl4jynI0s7lUscj8XUpblhJrji4Sxh8x7
rM5ML1c694SrpMQB3hEdt1QugYlhP1zQ/uMy5CGfhN39gCQzKok3X4O68lPhk6OA
cCO/dh+n7c4wi95kYxB7/qmBeVIJG9IFQHRydVLe4t/84Qn659M9dXRqJkbNP1Ig
HvJnGdGbU7uiNylqvbs+97RZto+icAhtJy/3ROemdZa7Gsl7S36o061fno8cnI5J
Gmh8xh4Lb0crIgNDlIdpz3rM9PHg53c2Vj/qCIJFZhZ0QJMCTqn81baJmnepQyuM
+6Hg7V66xUs0MB+zkDc1EA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1200 )
`pragma protect data_block
sN4gvOVnacD7dN2gCgTuqsDopbtlQ6tmSjrGigm4MzOddoVmnof9mHY+S28Re1Pa
zhVecm7M4LBK+5G/KKw6dW0pQu9e//XEgZZaGc1ZfYrvuIbsyOI1gzJwBzZop+wp
POj2OrQZPGR52Tz9ZdfjQ50EY7ODYiiDKNlygcq3sdfmRNMYb82BXP4F8L5hE7y2
1pvG2BIhh84yeGaBZcOymmwAO2KG3w4s36/gjJdPzmxIXnR2nWj/hqd/dfB3yO15
ASXnpzt9xbKPlEZJ+ZhgB9L6PHvjOaBBHa92R38m5DwLSxcGF2pqRpkA/d1TWzd0
F7ylPgsZrjVHkN+tdBDDCjrzbpN+VIPwPwytZ5Wk5IVscqFIwnggSob5RGxQqffS
Y8d/2BulxV+EZn/FPqPdWpPrG8j58SGS1kln1hspn4w1HbMb4zOYZXQajN8DE5pB
fGRfDme4hLhNTNOcpV2nwgaIhKGBZk3vlXpFGXF/TDSCaD/aRACPSwYva3tuPCm4
xYtzCyJDB9D16qTYD4wikt+GWQhSouKJWZsvWqj1jm6Xm/I+b/Cr6yacQF7R8Wyl
Ts1hMZe+xoXcAr/mhSPXXJh87UT6u62Kr1dOlyMqU93yG7IMDVNmu4UGcQtr56ZW
Ih6ZJNMdel0HN8Uws1kE1r4EWKGRb2EXr15HpgpItknIYr+bim5QE0uVgyJtA46N
WZ5xIyNcej1nTfzPAAfcDoZndUHvKxgzRV+oaWm8ZaCZSZijcs1sxUWwKqmTn+O9
UXu4+Vq2BnfY6xqLszKC4aGMjHhJcJBZdXCWmeknaKQa4B/s6aotfTCzCv8+1+aM
56W711BST7cOz2TR7qko5xqjJPYKBigy/8Wh2YmpAhKIhxC4va+3VsHDX9B1nN3x
kyLrX4ZokkKknFGDzTRDeFmKvKhkNOX35WJQKYxvy4tqjlZ1Sp1/3hF2kDG4uOpW
tBH/gPj/+AayVe7QQqPB5vkziGxjXowFjFlpKHZyq/ed3lLENd68uiPXTua9hj7S
/jrCumruBsNnQIIHybHl90Xo4dcJpNdckFHwzNYDS8pYohRXOyRyo+ZO1LJ7nThW
Py8JTIcT7A6tcKpbR/9DTY2Jw4vQs/yTzcTisgDu0tz31CFX5OOWgPzMDDu1dZic
ekAKntYJT44T36lUYb+AGWxao/iyoDP7dD4pYlDi7xeScMUMvX5I/EyJTwzHqd98
xtnGpNXAJRCRg5fpeIrRxl/zJvGYR9H+5+xXNFdxijFDTrcuxx+VNqPpW+Gh6zQQ
7U/gkLkuFxNUn7hDQjs78T6u1UE6Lba+MLf8sImsGZb4g2jhcbLOfTQ6bH5rhMfH
zN7oaCvIqotthccrO4p+0KH/q9QPAcaFLH4dQKdrxRv3k9ekb2HjV3T1g0LVjAaX
MkCOf9rfjFWE1Ts9ypXNOt0HP6mUJaGCZVsZD3asvQkV+Tq6nHlDCMt5C5adS2gR
w8DaG1ckm4kJunxA7ST1L18sIMMJJci2DLi7219xC1oFeMZLGRB2Tu26rD2dm9hS
g1MCbja/KGW6FH/G+chWc6QHkRtgS+muv5+rjVW9kGqqWQSfLKmiUXgJVqFhFeQs
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ilcRGFh9VNXGrWAzxPpBP0wzelZgyon6K5rgjc/DPSSLq3rNwoxJ2xfRg9e8+069
ongFgOjDM59K3l0EZ7ja9GsM7UOARD8XuqYFIztCNQbx9jGxs7/V2DR99GkBJPR7
RKG8jP0mThZm4jE/NrobMigCvTt/GUXsqoKM4oXC94qxO3KiWEv9G5Cgssg056eM
/s8/Uul9mQDSuOlYnZPkkk+rJhGYQW3xtuapMTB1tQ4cYQG2oVm5exNbyliwrOwK
+E2Ygyz5StsOXCvzYGRCUwVqcax8fHWOUT/IumyyjiZ0uXfayCDrycvguIV5xP2l
svYNTeSejd3uRq28F1sztA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4672 )
`pragma protect data_block
GIB05k+383bwn+klFjFsJUv7FEmpCZQAr3wd98EkgAYxwLgPj5S4RaxcvTuuc6MG
h1zPk/A/afQ1TKlSVPpEMHk3hy/Mh7pXh3+4BWvsmchXv5ZkjE0bz2Bz4ZxLxpi7
77Dc4MdpMHzsVy8VM6ep6pxvYKKAyKD1F8hai9kJxkpkhv61H9foXdF+1Db4OFAW
Q9T6IaIMQH+3olXMvFVy44ypa1EwDBJiucGYH21UjwgYJknt5i02PZGmum/EuDSW
G4IxiDlhi+3tLSoouh8kQvJXbzSX2o39R867vx6Q/jF+5FTgDhM6Amd45c/1keoG
I1spOkMCyQjQYIZYEJgxiWKQv37WxV+FGiidCjCslq9yGZ5gEvvyRRFy813WKjUX
aFKse2jd70fBwu04aOV6N6EkPXB6byLy9e+RNEreHxchm2gBtPrIvlSJqKQRQ52o
0ned2P4mcXcl1N57k9/H4epJ+Js1pFwfWiDpsUoW2Kbd1LbZqS8RHlGtV4Qk/q2U
qBsYEzw2w84LRlVHf/BKdUdHcAU5p9FvG+zxxPwKgqtqPyV/LUBDbOpomPNE6IeD
LhHn5WGFAc0qE1ht59iBzMrnuaE8lyvnv7wZ9NAAR365UkuHhA79f5vAAuL/2tYk
cwZYuTmHD+jJV7bUQkX9V/9ftgZnsLMHLKCSfVwIuoh+mGfGjZCCtwLibBme6ZWk
PCcyhbd28Mk/XNMxY0Ud8GSiqLlBj2iQcZbXjn5JLIossnssi4SSmMIHqbgEVBPZ
ULQDZhHJ1/8L5ISEFEnbaBjSnDgb1o2F+OeAPepOhcVEaBrIX/SRs+u5ijYFhhUH
cmCajfI4ioLPmqjFLgj6PNDWMvz25pzIGMUMjdK/g7QHqCQCJjldOW4VIySnztE1
MG64qzpnOcotBTWirjHgwImov5AWoFtRF/ObfRmYOrc1AqkBB77Xwl2DPteRMn1P
hkg2ofM97FxgSmUsuRtobmirrMcdiMX9AH1yUelpE8WQgNoAYWraZ7/PnIwy9gk3
NQmWUYAwLRtHd0gWtmxibI8aXlaCsfCHVF43hdW6Ak7hikHPocPye6HnEU6caLx2
JZyePH/YnvvQrSdeWWtAXLoI3IoSMB83/1RVtwykOPaOUC7Uck1zHZ5a9VdR10uM
jgki3bxlKbGnIHDvkLP6wwgWkC76rfFMejDAOJme4qcWAXyMgsoVfuO/smE1G6xO
1LHnmT2/EThAdLTkK3STFEB9JNNf4rVmsNrW1f7HAKB06dvjuthygEKGhId92H2I
xTcV0JaCJdhPhOj0djNMbzIWKLwkD/p0du2PTi+Gz+MZPEZm1ZFsg6ICy9JEfpMW
L3nNiW3uU9EHsPt3FrBmxR8eLTR1BtB8Rb2JLAxLFqG9Z3lwoywKI7vuoV73hdOk
iVHbd7JwrkVcW5xSrnACm7LPd7N3DR8cLtMLG3KwqtVOdtAOn+9W4rH3vnea6eV6
uo+CHYgo7S0NeV6y4ikB/L2jwOlyvXstoZlcS1NSHJg/WFuzIcQokIWVecIwCvOj
wlmCOTVTC5r5FBCL1r1tkjlrLGOOJNyigtCdwmXYAoXt9jFxG6YtQJoF6AdE0wI6
F0OdLyW+44fH/iAX1TdpKMXJ32S+LGEbV8QnO3p2imfrQLQx8+77pKOZVniGbXjt
9WyWk/vVhK3f9fvR76NhfL8SDvzyeIti9DmX/nRv/dpBoB0zlu1ebYGzCd/P3Qor
568KwxwBYKmb9YNw9+Toyz2J27es0rDeN6v0q+rbzet2LwHiyGmaH34UHznwJl41
OdvLjE2Ax8M7V4yK5sCmP0LUjKU/ek90YuA/WzjuvNT7GD6C4C9J5LWKS7qpmxqL
NYXHL8K/uOOYoeeX94EXKamVBBXRZpksC5iwBcolFrONdVh0KlcHarHpz4RSrWLH
UnHxCyuLxX+YhR31mQG9ejbc+mgA8qTQBM4pA1rTJTNPlP5cxP2DL8dviratxw78
0C2Ty2nuvo964+nHI0OiLIC+b99HcAPOten/gN/fRNFogAbkVKd6D0q1gnULoVhf
v3v46qfA293k2zsWBx9JDHLsdlx8rJknexIhGicmrUDpXqM3tyKHXxPTpvb4VDGe
BOLmBnEqC8e4ewZ/akLxfvj3HzwGyaE/x+f6fC8oDWox1x2NVhBaWCmqUsGZ3Nbo
eFXuJbuDbhNSeUS4f7a0KFGTWBoi9OrfuiRo/qg+HL4TxKEQ/8PvMp3OHzkNziHd
bO0MYktY0cYFkuNxwcDYiszibkr7eQGLUrhX3gA8s+MFx08ZaZKQSGw6Ft55FGW2
y2WGC+1s8Mv93vhMWc6yUDOKZ5V/A/zDP8YSPMJOhsr1XCW/KEWJjTpDh9zRulWK
CYTZBZMcJIlqiMK469atAAjezvNfi0REDQeLShv9XuGtri/tTCVv2g1t4gAWvvP1
rN/Ac+23zHkCl4eRAfQDfujHYiiRXopTa5n0KT9a/y7W9F3FeDeCGHURZdK7AWZE
6x5DjoxdIAHT78AJwZ5P4ab+1wDYA3VVPg+piUpec34+CTV1p+tnsEAZIKZ9ob/J
H2r6NbvUwxy10u5/s+WqDLNpZcCMQpcYJpHhLmE+rxbDGGtIbTbYgReHVAsdKRT/
pc/m6WA0QKqInhv8a/mESqz+ygFEzY9niLTI638chOEZ9yyiAG/ty6EBHr6lI4gw
FrnuaicEUAFjRlVEXXi4wPplivDtNON8ZTRKi9maBxI/91C1hZ252jahA2hqt1f2
6dbmTHPmwlBFqNw7dBc4uUfgKJhej0WginAuJ7DidBO7zKYKOs738Qfi4czkizK/
DKRInXxIqLGDsxiz6dH5uD7SH4wTjmdlSonmf+LwKL8ZO+cTvZCyt45CZzq8A4+/
6Xzt1f0k3spFS1NnEdVlNdkMitlKueUbcKoqRUNjJyEQkRqMVWEll3jJQfVej1Px
ARw9qWniBYjdaJmCz4i2YvDgyU3DrMB5mVctIGEexpAqK0fYlRO5IocTlJ2+gLGC
xHX4WYnxo7gz8QgeYuwqWHdd7AeIEKzaPw+ukCBpVegeGz7sTMVL43v3OMalRu9/
Ur/o0WjMO78jAiHq6INeg4CDBATaoVQ8VQgy4mgOkIgTpi2Fynf21tc+akYrq5cM
nok2H+5sgCUMtO1QTTDiNyX37TnbzGSJpHaEFgOvxDPmM461NbvyfcVfi/tw11N5
uWr2ZigKnFTg0UD1s8x9pe4DcdehzU/gTG00/r2omwO/XRBIohIRF8+wXEw8qVTJ
xvoBRal9EtFU0C2LlTr+2fM61L+dcOFiNaCpkdP8lsx3rbDvRZPu6/g+hKxeg3z+
+muoTZcT4yJnk52o0QkCRUqAXDPE7Rkw1UwcJotQmUr9dAfl1hYiRdR5Q4qxq36q
dc7NVBnL9SezC0Jae+HDCtQlgp0T02fMWzpIEOZEI9ygKo5jRvQ1mOcg1E/g4N+F
QOy+9EvFuHpvQv4jE7AzjgJ45DsTVR4V+H7s9F8w5TcROHsspKPFOAXIcirv1NG5
XXvABg4kfZbSvFqWviQ6goc/YJ1cwejAwlaLuPKHQiKQJYT/pf9lfBroX4U9Kc0h
335ESkNA6Zwr0OQCuDYO4zNsNLG4i7HRZ2tX+tvDxDykvgFAbZOmu2pw1iggDWzG
pNpGq05rFgmoWT3297OdMYWBr4S+Hw3zgmnPaNC0YFX40YGlT2YMIlhl+YY6daSA
Lea/dVzt+uw6Lj1QPSM51joj8D8+ASuQdgtPpicscq0Ddg2HBIIrTNDbxiAWvsoE
qa2NLOwzzaIRo0G8yxY8kLvXp/MHBaBTi3Apm8DqJOJUMEFasa+1/VGq82rRm0c6
7bfLPz+0qjZGeC74f+TEkNixGxR9k+9zRHSpd7LmoV7ID5JIJbZ5UMVdSN+rHZUm
/nsmHdblhXfZtR958EyW7BiuV63sDOqxF24/vKUe8FEjIx0tnfzRFeIA8jTGFNI0
bvBTcyZ9DCrUzbiJT+f7JqEAUDbsigaBKGKW2bvfYp9QyRsP4sDxmO/5ZCBS2Mwa
uhy/WwMvZMu5ZfYPy5gpdPrV9Qvz3rfNbe6hEXMJzV+UwIFhMKw8mVRljTK1fMnA
H2sx4gtEJorntJBun+Bmg5EKlb3O1CTdrEi+9T/qRKYMYrIztwyM821MGf0s3VaG
jbGYCDk8EpKhPKCHDTaHnH4KYJPbjLYBdatUOL9KC57djG69aSeG0YnkE8iNBDq6
OIzY1DHa3ruYPqOUmCAUuznTrjeEmeL5wJSNTfU1Ri7qNQzfHBJsJZDAVDfn7nAl
lY+j0Lfgzliq67YDiiFn512yTl28EcY0GeHJS2Ku1vKxJnhpzsj5zOOQNxpxjYtz
o/3w5HCgJof/5Sy1pnlrV9b7SLfSIMPK8X0rUCIGVqkJV932tpDtvrhWUi0ui/Nr
EJS2QM111PcmsRh2ddNDYG9IoKJ9qsMeqMHStsV8eUbIRRz7kM6FcPIA3cfTHlSb
EUwNEnpgj7ROz0u7eRd8boPMahnGOwgIAhGFHT7Db79epMWs4sN/oo4KvYUnRYSy
qQ0AK/rNyS0nBqGEQx/dUlRQFgdcUCAalYjbD54fbfx0H73e9eng5KIuPIauJKiW
cPJCdYYRMDEX3dhIMsxlRWYEcxDulXu1hFE4GViwwRko3jr/tmHszPVXMjkRoc0+
3+McV6bldv1fiQhgJtpVplxuyxZQ+nx29BRQzQ3Nn9Ylks/E9YRVagU7k05qqGIM
VpkK/rhE1p4OOAG5VNpd7VqDRkHPusZLTK/OSYFCyykw/uQGN38GrXzxBo7oP1L5
vVjmx60f1dCTt0INLbRamgtKF27OmIWskqQVm/jOBWUNuD/tFBXVeRECN+iXDtJY
3m3xzgb5SZgrGoxu785poguB+rPBLngsuL1AJ5E5MAquj5SkMq8nH0Cs3hCXjV+H
961XwZHDyKdZKFccS1S9RgRLKshA5C8WI2iIQ9duXskJVyAtcDlQ0Ryd4F06Iaxj
Z3eFaqoZ4DxpFShDKq+/wXmvuPx/ymqZmj2d5Jerg908tuzDKTohjqnwYXXab3PN
EpCZQaNPGynurPgoTvKoskMghPjWLZOefPIkXs26GlWj+BVvb8c9zOnP5JHZSUIm
RMqtpzd618a7X0ZvxXk1+y769PCj25X4IoCxPspfnc07liN9fgngDBgyakkM3tBd
EdJPuqEXeAJh+kBB4HwUJCZMXy5fyxBScos0Q5sXn8oa2Jc9QhjHDhGO6LrUVV7T
iRXiPfX15KMxqHHnFllKgWjOzKqLgc1iRRMfCP9dx4tI+LckkNUoUBw9rwQdBOeF
8j9lA7Nsl8/NPllL6VwQH0rNvOX9HJNOjncdtJ43O9rnRj0Di/1SWyz4+Fjcoiyn
MXWcg7hoMwIrbGm6IAOcJUIzFiETLl7S1yFYuOy38uNtUxEOQt8n3ZIWXad6ezFJ
+mcjbQlWQtHaGsguYAo75yIKO2pwL0VtHP8DxCKgCR2k3j+AR+88qPrqnUuWgMY7
cpTds8NtZfXpF2HrnYTqp1VFpzdld5+o1uhAvpF5gWvEGMXuf2FUB1/pmqSANHsw
rjkwJ0N23IA1vRjyJKizZlLWsrGtN6/OcxY8BXHimf/NHudJBpiNSzdq66zBmru9
cBTdqnsOnYrkEyOLD8FYOQrjOxaBhvM+5mo2TDIfyUXuXlxQARlScG2SLwpt2uDw
nsBwt/wtdeWXwKzo6ETaFwQqFk4rw9hu7Fk3CphEu0hTUjyb6DmnDbU+KjJZgJZZ
Bf5URm20jQDYwmUwS3WnVumBnDP/p7ax11VWfGLkoNk+7M9VzUutaWx5vYn2Q4CY
fyYVgwpOvGC8OkXcvLPf2eHZIOpAiFEcZGbZXkvtQyKU39ctQuYMVO3GBhPytA/Z
/Jy1EyMuZkNaehgPR2Z94TGYwqxtPjTjRhtROXED2ZK6PDRiV0pDBW2f8wACVdDq
CleylFWL/5jFNWA5sVVeqb6plNzZSo1GGEU82QYEG7Hyd+EsSiMuPOnpHeRa+tST
rU9Oe80oFvSw0/BENTqNt6X1jN4aFuhDmQDEeJZIBDsBofXc7Zf+wYULM3YrAiH4
GYIqDxIi3W/VTBzbqemv/mvJer2KopnY9XAEQJgdVF4vnGW6o9EHDoAFacoHCOrI
5JdYcQ0zBaKT3ONK533daZYDhmafX4bvsqfeH1+D3IoojlArCRBtdD0SK3e3vlDv
MwZnBfvMzof2mLXI/OCz8w==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
izvgvDzAcpiuRRxaxdRKN+adMm16posiYX6l1yab2fTfBOCQnTjJdEzNPeh0heYT
qtTGS6Edk7iDsbUSend0MKapaljRW9I52hwZv8yFuc2VisI2DNFtboZDPgV1l1Ns
eSiGELAmxs6DCIlNUrCcJrsfLiFQCP8w5Z3MXseUty49sHL0wra4M5FCZ+0f85N0
p5yibcd80LO6Nff9oT7aP9DS3fbDJhJ0jhufPMMKLlSEQU80iu3H0ZdPWMJs3Pp1
NeoahxcGTxbxA4JzooVQqZlKtJGcwj2xbHLCRR65k4+gHM1LwIh2/IWT0+dCJCig
M6e+d3qoXwVVgdviDX625w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9344 )
`pragma protect data_block
SUZwxv5a7DHM57W8MgiyCbhbcIZm/E/JYKxrINfAF7IsuTSLo+MrCBvMkDqjdDg3
MzT/Pfsn7PtewbcTV+037PtcGfDOWJWhgq7LHNB7X4HoQeSt33Ae6hyp2jclKz1d
g0BXVYMLgd9RXaJiKQ9Gzt4kJ8E8i9wLf2zUv7MZrQib4FAVCQiPDtTJECbggpEw
rpzI4mhDg4/QuuJzy3e7v8WaROW8+nU4qO8azTte+05ugugSjPbjX9x5kRJak5bm
1ISQPmHWf2BFcQ7dxByLfwtL3SQbsfW20rlWjghWPGdKvnA+4FCpHKX7Ay2ZFf8A
qK5WGarJwkT/B6iI9NCsTkIYYp5BRDdJxgMjXl6b7cVs0qx6pEmxHyuqFFh2wuM6
j5E3oqZRh611tXwcxoBLAY/7CHCwezA14H9+VnenZ7Z8r7f1B+Cu/WcOQkLtAUOD
vejyejmdSJIDaBoNStZWAS5S+E1FiosvRthOMO+hvpeKRVJb/LlwUn+6LpYWP3bn
V1//T54ZdOpxi1bMVZbki8F/dnXBg6QkLoDiYSLCr4MK67aG9EsZW8GZ/hv8/u1U
u90TTkrBFYvUumbOGRCJCT02JdhuhI3yN9+EAt3LDKygXSPmVvdfkegF20IzgMNz
E5OzElb2JnsLMIIGccS8PXXtzIxbnkxxA9OaHiUH2dW3rmjsfuT9cWnvOyGHZrtS
hjq+hnhtkUekXYSq+kO3sKWmojJjxx6BdJOBkXsB6Nglh6TQM/BSyt5mE02OavbE
ps8wN7k8BSxdvt8MkcoMxVbqUOj0isgzyeAfyEqjq1Grq4X/UN7zTNhrRNIurwXi
4vdbg2vu8hkNP62plUAZ0wCHSQMJkS3uilGevRKxJsf45Kd1e/IR3dGTj7QbIAYH
ZmG6Cq5PzTwn8wEjn1eU9FrzmQhqzSeJEmXxZDsjuHui6462pJmLzrV7fD1owOvq
lwH75PCTdlSoHJjeF47BHR1fKn9VPoB8zsRlnKDSnOVvP9o/8ioLGUzFo2N9fkXO
hGGgyTc4FUK7nzINvd9qraIhGFwgSQARCeiEpFV8dchdZoOVPpKLw6js8vNNXHWg
RfR6HhCfnJWNFV1gAJaRKSn88c5WJilGzcrm43f060xvFyUeOq68kH9O8iHQuQAH
53ZYtEnZiYpLyxo3wD/SPi2EkHgsekVNgcbuWTzXatg/+kdcRobhaUT10K50MIam
+th3VfLJM58KoEREeb7Lhi74ii9SQf/OyCyzW+kWCyExvsX0UddhUOnOsCXSVuHB
1NaslfKv6ePo54PnSST435uuWbBDTaubo1+DePP9nnvbEmKR7DV0Nrn9iIj9Ghcz
h9BsohDu3DT2aV03Hjji2QuZFm3WSEd71L/uHvucxvwR3VzExuq5IKAgeaNtAmbY
d3BO79NfUIHNdMDrLxrN84xsQphWt9qQZS9jIGxlNGesaQoSG2iVG4sP35Zuxk6D
0sgQmgpNRCm0brqSJF36HKk5KarF2aETHtm+56LyDWrwy4jbvsxf78jSQzWSNzvZ
/pGenq5Q5ibhGEhRrIKqnMuN0Fv6Zgnj9oEdThGmjL5QR4VRlP71U/xheXFK9iE5
2gLt+F8kLsCky+V+tl7FfW0cQ719mFvgHIP2AEgdyjP5Tdz7I53YSG95rVhUvocP
T5ClHQDiyvuWoEPEjQrShe64dv/lh1twPA/Cj2zqwtSLljlRxFrCdjyZsAZKMHq4
s8qDSQ6uhU4+OplxtHfWwbTzHAhSvyYci6mzOfHxK99bsRUuwxUpS6wxaQOnFcia
XioE6eOI5awZPc4o/9Nngwqj8nLwaLh/+k6361L/DfiYn5S2lpXZZ77+3QMsR/LH
moth1dzVG0TUG+CCfs1XYK95uBV+j/oIVh3aj8Z5L8SkYqvpwtOFbJhOaZosVK0p
G172K0fuMRvYJ4fuzUAKpStnXnjnr4SZTKQ2iAqT/URnbKIxeO2ZU6IUCmDCFl3X
jteD9Sml0KFis37g89ZAsOfDZW3+bbfSuAZdiZBlW+6arjx8rIV/KuRS2NIm40As
Txh0BDMBDQWAgiOm3LKG7jeB//3Czqkzt/MxvYVbW9rPMVV7aj9SXBs1iLC3b6DM
aojSGTNYA3I03PRpFndHADaYEz8gPKic4rlKK1VSDVIuT4zs63NYh56Hs2/cEIqZ
ufjSlN1I0S0XPuDVscn+jaUOTHwHPLOYGjWX3ofoCFqdWHynsQ5wdkoxhBUyAxC1
/6mjpYkLBNrxAXuuJZ1eBi5QXH0D+KA+aaSkBkbyJySrntut64VSzbJu2yIHGbQ9
VIs57Vj8HUhhrtv1T+mRLYGm+YlfNqqTNbL8aDf5/E1U9tw2rqq+o+Impk2c2OlE
34SvYjhpkKRxhwyvL5agOf4IsgEyYZlJhdEfpeMpivLEhlH+ZVIcM8ymlhbWCxUa
UDsQXng5GsPYhJcMhkQSghzdAmrimKU+F29vVPBzi4N3aOAYijJEGPzIrTz+vA+A
fB9L5X3yWHWltojbKZY11F+9WDkDuVbwA7u5soGaMvsO/7mwFohjtIqOSGaRwu75
pdCSltvuzX8wzZ4/PQrO1jF7U2sUWgMj0BXJKig9Jtn+C8g6BMc77hjLGDOF2D1w
cvMA3NtB+z33yKccozW3tUsHtHVq5x+vYEA1MDMh1mCxl86ZnswUL/jcOtqvm+vW
r6G5DVQEE2/vH8p86BqhHjDBbw2Ja7Ad43NZFBOQDE4RiOZWYdow+wqeNqSEvFcZ
dMc0sf6zdaWbpegOrh7bN1ou2u4kFUMD8oxKuqLe8SVTYwDzYNvEZAQEKWR/YH4k
mv8e0/mZa/ZxF/GcqrD8SBTeRYy7gSAfs679YZZZiJ729ihlHI1Tn3RLFXeNrLDK
4cIBU2amsPhZBpwCcAYve2Hbpxz6F98ZRmzwWBgtNPQmpxk2z4BJfkh+N48cIeDl
ItJtDo9oE3zmuHwX0p6s0D+yTXvh70TOwNO7/OlXacxjYdejkR28fgxvG0I7hQ+o
qJqG8wwlaJwMKDJV57tDgrgo7pM30WN3StD5vOU4hIcMeuAww3pOjfdOoW9ZBXjV
yjQJsT4Ro/A5K2K58DP33xdybZXRiftN3tK5rIvQ04D4WVdqBo41+YXXfZURcFiD
9bIn73A3Ks7HAgdXx2AqlmgAqhA7LFA37/QKRehbXF+VMR6bAkKC5K6w11vaLpOa
DYTRjKeUEBFa7/ErDpsgscFoascLwmdwe3pwob+FEplNWpgfZuPYxGEmKkr5h+Vk
1Zjt8tT6sPUoZ+hUmcICx74w1jPvvez0mJNpzNQravoOQWfk/hmoC2cT5LQAZQ8N
AxHL5s1awCfPswdMl9jvTOXVIoT/JU4LkHtGXF86C8CSzJtUofM6TxbXKFR6P2ON
OgOpN6rkeNsvzKyPunKQOxUoeNGdUGwdDn2nE8644evDiaA0q0ry0g8vS6veMcs1
9AFc6h37C+8BN6b04GglDipRfO3HTMKVwSkNcx/dCoPH05oxP206nnDjC4zitwSJ
WiXeW4WXCYMIGM6t+8SkMvTp7Iy5E9faY5QJ1Sqh2AQRuhKcFucTbw2Q2Ygk3cQG
zRvPzIcy+FDsj02+flMryYpPz0bEg8xECudn2Ph4TKsci9xkl759zrTVqaAqEsqQ
eJGhih/Jz0Jlya+4gYDZ3mcBJz+MTp9xIbKXb+wPKc+PiXeClHWXfGO1cG4eWFl5
3kW8b7r+iN2aHUgiaF3dhDbRKUgcfBZ+NML/Cn9dcyLUjHxAz2qpy7qCXae0zQY5
SECSGGDm7uFs3gxf85KTPbgmzpT9twLCEgSOpdy/sUr4H8gzmDymwUH2tkaCCBpi
S/iq7Wt/KtuHWWZ3/p5vLR3fio590aVz/TQrp2tu379qZwLcEezkV4lM8MzhF5ay
mALQdx3Cb1p0zd6jJGVzAB1L7T2xBp+6nG1JgMcq2inpULhqFvH//KR4ypg+Px+b
s7C92PIrbQ3W2UnH9Llg6YXr9CiQ86UHBKmFFs0PYSL3jIHuY11EdA/eHLIJ5MEm
7tnFst76sCZQSj/N1+pCe2Sel6d8qtirQyoq5Nr5r636I/r9cKMmTje/kiKf2WsJ
S8mv4uPWbI2JeFcMHNswRV9PjpNDfeyB4L0j/UMh5023pHa9US5CfzwMBMlmWbYa
2teEk/xNzNA9W/dT1dJL53Slw6hdpGa7izK8UCKSE5IadcxFRtjj/X7hoOeLlhem
jsHcrlF3vqzrxR7lMRYztUCCj/9v4NYdka3t2IplRMHdUiaZMlCXJMcmqmT4JDvW
+rTjhZA8rdZPVF7N3ih1iGNlWbR7lhaicBm3UTRRfHuJ1KY83hi9ysai1ScMb6ut
Dv804nHxMh14MBXWW8EWnGZGmcNrA99XRoDMnT92dEHtJuWX29m9o2aLktWHG0/d
T6n6MRcIJ33m2Uew15PJwH5dw4avR7rrP0KUMeiz2YsODhQimEHgP/qZfI5sbMoi
xcTD9Q2CntmuiN3JgUAop/9f7CjyBiO9eHrdriHLW78bd8O4fGbJ3216C1tb4l6j
1Tdw32mSrj5kvgybNXKZezQ5UPQpc08BLbGN7y5f04qQsToj1yRApbCzGXgyK1eu
hMzw3bUg56gBYV7o5HFbz8Lzeqrf+olMI6+Tw3Dng2NfiUnXEyN+TzxxGyIoOFnd
yvOAdqS21wq1miwGQkgM6VOEBCfUO3Q8U7gMktpwlAilqgkiGAqYwqQKFyVQKwBG
J1yMyQk0uNH0JkdCp+86rTCyvSXVYG66aPKZ45UznCCVDI/27ZBWsJUAib1D9Ksk
jQORDNWT+8iz2AgXkg2lIoiYRKGWZyaS2h+D6ybpQ6SZmWY3Z4tKvvgVDPoHLYNb
QPN8tV5aGXkiGBve+nz4tkkXT6XUkKD/Dihs4XV0IJk5E5hebqTpmZBgZrxw824M
a/dddpofheQ+Fw+YedD1HiUOCjCdCC1uIGAFG25O5Dbys5CwS8uWezn0AcG13H+y
HJqMjw36Og6UyFnaUbkZIiyN0qFO5IKNnXjgomeFJXzve8YLKy3cuSAlI/abq+s1
GyLZ5WDcmUnm1LMyPTPW5QZa/TDVEscOzbBborgK6fAORaXQTRgKVSFNV7JPE45A
QNDpxB9IxFEkYqL8YKCnj78mwcvDmjnzpjzmATpz2S+WDHd7WLPj6Vi3brWf6FbQ
B1xM/Qdu0Tz/3pXGAEXleajTkmuxdQWIQ3RqRurIBr8FK5/nKN/YvYbq/bryClcl
okQKK0184WqQQAEkGyi6DLVNbP5mc9beBCuY9eGTIyaKRqQt+9sLv/WN/INXWg8n
r82oqEwLtTALI4KBD9DC3aKnSo0Vh43qnESV66M0wMHrbxX61biCcEDxF20x7wxm
3xwLvdcbKBwiNcioZ/r9YoOSnxRDS4EdtIkDSRXeKKpUpSttpJhqHxpwIf7INPRz
i7dfiOrBUiH38Y49VTYSip9rR9DqLxZS0jiBve4NnVfB0R6jJQPYLKisDGgdsBpC
uqvHbk8BOlRxVZSbbuppBPP9qDPtIAswTWuUOa6BD5foEDh4/+kq8yfKnoeVZFqM
hlPBgUTGsdFhRIrfOzxgSZBaj0Vug7SMhkT8RvjXS2z1noOzpBohYxrDNQ3fRARr
Ee3EtItThSujN0atqDpCHxfQNKXS0CVpj86p66AWd/X3OCShubPRYefFH6D7vFdf
JvESw2MeSfZOgCJhHPXMwSJ0XjE3MBReiBXlj8XnWJJGdW6v203yzcT2nJlC5JBL
8aILef6Vxr1Ti5rv39hfvTTWplhmiStKMqz17aTSbAdjaEHUL7pixWfyLXNBVp1q
a4+QUotofYSazh27E5yyVSchn0r6NwZad0RwDicqp2DGslaYYvT3BOENB3ML9Cnh
byDvL5gLxAQoaEMdOs8c/lxOMJzgi2wgxNJitWntkuZqExThyTS3B4PRXvunudDs
O4v0CJvROUfhrx3YmTRvnIpyRFBK9qUmUKPZTkLbHm2cbPaMnRkE+W2bQbQVMH6S
qAAYpENUVInC+F4bHOnKq6aAyrOlMXQCwWcYLQBufVYe7zGs8hA7QKrEmuyZH9pe
kpjBtTYcBgKYDjpu0iAJS/JClHKmFmmjNyIwARO60ykpLt88moarwIMFpSTKDPqh
Ap44GbwKTmWGsXL13fVjxQZjafsfNae2o5S3qKGbwB0bbgDMo2W917XlxrYZkSUY
hiKBJlqlEnxYfVrOwDVVY/0uqNBZWqQBg8EJchM8tGZbRXJuXks9+Ik/bvjqtp31
OnAREHBimbmaIOjwQfPNU2MdL8QGbOdvqLHHaAuYkAIsPP+s2JJQ7OMve0fMt0a/
acfuv2BR4phuO1hXNQhJnWhbnOniOnqnm3s4fIldzyX0TDXJ9zVDRUsAXf0xHatU
2LdGyXdxlTTFBnG2TCbsEoTNysT1+hIEsuiKk7DW+z1tqJCK63NZ9O+SdmYmb1mn
Jm9F0ja5CEz/KQ46Nd86kv09Ptzw8/EmX/BQlEGzcFp34tC7OdtXm2iF6OyjkLq0
AVUreMsShP+s1iCgFPOBAxtnmC0uLJc+vQryT9wh6n6UCwpIpK8SbiXvnAHkxrrc
C/lnCU1DN+wgPmJFYubZM8ANlwKHMlcFzB5vPgmJvc6RLYvcMEQ7AWGszgWlkshm
ZGUW1pb0SqLHsKWautgoq/9QwWbYAujV7hHHU6kUN9i1H4hl9Y8UM7GkmMEAb8+e
4/0qFucop6WPV0c+z4iLdr/i4RxKSoDUfg2QPcLLhowMMas5VmviEDNRYIfUvhAg
QwQ4Scw+yS2FQJ6OEtah5dBQR+HMBm3KIvQBWWkeeCYKcak3xGxUSf/ZoDbAhSd2
g2x9+aVfY1pv9l5bKWeUSSViFjG2bz53qP+Mgjxbg3g9991OX2YTnn+u1mopxio9
mLfz0Ght8q8gzMLCJJpLNdaXmx+mgnUKKiJ/Qe6KiGzgD9exQrWvH+Bo6AtWP2oe
obzz3u47e44SBVBK4nIHWm3vT0cwIMUHY6NVBuxeKAuwLPd5CFeBGASSO93A9nBy
HB1CzRISAxZPEsYaJkigXgWuTSI3yDYCkQFUs+UNhDHDHItYvva/qck6R7I6tjKM
yjJNOmfgazE4KIfQqFIH5Jv+hqAE/6FRylWJtnCjr6op+Wbo8ebN+17V4ghBp727
qtR27KdKU4YcLsSKCCnLu36rfUifU+WN6hSUE9T7CdsOz/L5PwHLJz9e+UEJzyu4
B2+nT8rUG4QdXkHXC+WrcWFtheb0MkM+2jChRr3QisOKhqBNuGPDGQoROLw+IEC+
ramQfu4sXh5UhwLL2nzIlNc2YoRtjJghtAhk9dLL6g+vZ7bQiSABucfHKR+0HrG3
C6KqM/0s7/JJ6gVjTK9lLQAQUhv/9TQeAxLYyglYMZc7gAJQYPTtgVDH/NhC8GXu
mhKPQprZWraWVGQpyJ0+EU+RMBBgmHYaWSCzTCnRVsO4j/9fgxTSlxA80VZNk0hd
qq6j/huHaS3g6LCLktGm/7M3XsE82jgRL7v3VVoOjpShjASakz2WVc/Zh9h9d7R7
aUQZj59iHmhpqrbVhRdlS2vzWVfm5Xzubi10AlZh8NAM+kek7oPeH0aO0CBjngX6
pevXRL3n9EzJjZlrYMmweQ9fFjhhBfmcQt0avxWDQN56YeoxHpACui+xsKYpqj9f
dgMid90KppwPRIJrqI3a14inaKNJof1L6HKjI/2CjfIqc0QVSFJgfBDdyTOEnetG
32wQdE9byDL6aRkqSDmIKfUqB85CK/9Ow3k6J3fO/fgzR5QocekDJZLOiHlZIXZD
5xi3Tr8xwZM8gAq7oy+LMobHZHeMv/mayA25jsqZiCCiMoQcUXOUJ0Lsgy9sOK2f
IQuKGSdNzViCrhsiolbaR2sTh4yiZ1fs1yZBrT5k289B6Rjt2OY39+92hspnTmbY
/Qp33DGIr77EcML4MnUkSkNmEj1SSlEEfGZuwdzwR8bzCEi8QHs1pY1cREGr21CE
Es6xAOjBWsXSb0yumXear3D/iz/nbBILL9446EtzVhva3lzNVI+hWxHmx0nC4yR1
SYeov71Zbp3JErFRAgiZX2niEgz+LH98L4DGwIIDjmtObItu0Z8P5DDjMtE16f1e
aMLVy22BZST97I156m929coabxQCuAL5Kk6SfkBRGTm3yXy4A55VVNMCONnaaW7W
U+tThsLetzYMIMYy/iL+I5H3SkViDuM9Bwjh1IABV6vVEpEaVLpApcP1ryi975bO
vbzFmVNWd/HMumhB+W5kWW9MLjj2h9LEU5k2SJuaGgBLws1lEhsiR0N5Z2+LPRaS
AMmTzYgUugPqFNWkXeUPWDeH3BqgNVJbFEeuIqf0xD8FvFPE4gu3A0rX6qALisYf
bEeixiBEIxaZ1pHk5CfHMQVII3T5hqZ46buJvl8TfYeDd/srpTvBRbtDpvlel+7h
3HeMiScyNYBhHFz29f5tqFWlQTovJJUAZloUunNkw1ycw0FxgEGidh4fjUs9BzZh
FvHDIGQYHIOXXx1vrNDw78yeBFIVib6bRPy6GdpvinyfP0vG1Px9lS6dV8944Ovw
GHNSPwaCEc7wUZQOqXXArvzqblqDR9qKg2hLuXVo3sMwSz2WVm4DC1gFQQMAUCf4
hr52QVPvoK1mP64syH20zw7GPioJJXY840Fu0kOoZZ3HeEJbeNZhHibi4plxO1+9
Oz8WFlsRhxX9FDa0SAhOhyJHHs1eXq7oF4yVTh59T7FBO7TxFN7UsPGy/0dbOxdd
RNCFp5BRzrwsixZlYHvEGrq0tO1JhvGu3OpezLtpmnyiM0rarl+7QFgxnADpL1mr
Op3ef1zcH8/nTQIidwoPXMHCsXvhcDUCik3fN7puJZgI4Wpfbk+qMnyIYAvNoT13
tB7PSZl5ItuiP/xwuJj+WmelAq5ib+29E6W/GNKSddBAKSsZeivB45M4ZxXBP4IK
dOwDIIjsmsnQU5jXWR7SSVwFYIBBYPkLVlD3/juRQiCBYoU0ju4/KbdfvleMw9Fg
WdBLgCKBbH+7vPFhAugzP6RyliG4s2T4Db2PApCriPP0eu9FRWVYdc1IGBC9qeXR
pq0ya1CY1cf74qSWgNuiuDnZgUynZnRs7Own/NcK1SURFUs5mcSJa5skFEcdXFPx
CIAfpWDGiWcCBcsZkHMhOm1PxDqlPr9MyV0/HM0BdFeeLJEEXHnltQee1wDuFUA3
xYtl4SxPlHdze8p4hFiriAmfIVhsWe7+AZ2JsL9yb/3z0aZMUw4ishNu8qWZsVRl
haCnr/Pe3hmo1oXHu9ZmFN4Mfbak6Fyox6YQaLEW3i/zeKumKfe+4h4+yNIwXDPD
KwQCxWc0BQc44WbvzghyR5mWsvY66TTU7kQy6UiELg6RuvPefZ9sXX7r3ylI3ppm
uNo8H3efKchzyoCjpg8Q1gpsH8QlpQGH/cBUsA9eOs8qVoviH4eJ+48oUSxGhLFE
dTwBggCNJoT51jEFc+gM9GOD3BMlvO+LGEhiuyKdEbCnlDgJz67aEKsZOvwnntQ5
OgmttVovHb3yXVymW2Zzj5qrc6UZOpxaprCI9hj3woGJ71kBZW4eKmi6uh6pXZUs
n+NfOGs3n9PX1fJZMO+jKS7HkvDy1KZvyNBGmg8vmd4EjqlN5WknlMAKh0qIO+hK
6ks1lFptZImBgbPS6bx6u8EV5VTuKnj8LgjDjaXM6TTkfacqB8Jh1V/EwKUoKy8s
0W7bYCdF1saKcXJygafsftPytdbpum8H+1D49CqT/xk1OV4ZKmc4ZVs/1NiSMl0R
DWRhE3l5xMYxqebd7qxpBVLyI4PKK3TJhnNF0xnlpbq7D6LTZrU9kUsVkzVvuof6
FuUHFurtbt4Hvtb4ln2RR6Tn6HCK/D1y9nq80B2F8RUsqvw2oqKx/VX5cVyqFOvD
j5cVhcTy8fiKQmAsBiaTB2/zPo83Z1OZx7dgxTdS2yszLOs/BkPvCZ8aRhkfak95
ItrSzSY38Aw0MW2876C9z4PToDMgjeEhA+vQ293Ub1EBVhcG5vw2D8UQfdDhTWDA
VVMIV/sTXCQjmQSmgLxsDl7/37iojVSOFALo8uFamleM81I3OEjJ920bGRefQl7Q
pTC0CL5AEkljkFrQpZX9ku8s0J5y7FogYUs9IUg+L7ubRdYg/Kw9y7lrzj61OlTR
DD+oouBnj4JK+/cm5g6ouZVJR3UsZlaq7eRL/s0qTnx0eugFEF26ptHfHnppWVY1
Ak/Lyx//xuamiKMBiJBsVXiVt77So0MP74Gj5/21jqwFNXUnBhOUwH/GbPnajafm
5CDgXmUbDrLTXm1d2qWR8DMKofU7FXa/7HgQ0Jd0pYdsOVMOQ6T9NtDCb8pWcRpA
b2f8qunbj5v2Vs3HZzyBB+yA/I4VpeFu1SFXhxwmJoHyDHiGGmeu6bmnXhVeT02H
zvDcMHf5+ZLKwTeUrNhI+4ujzAWq30QQkOnJ1l/t31R8rHP7U1rDgfMwjMcmPddv
YasCWxm6w1BqJKmyKWvXBB9Njo1TQ0hD50JoxeDiRb4mODjQsPmZmpJyfauVKA0U
KAbyGU0qXTh6sTRSh3NgJFsGC29so3robqM7p9C+PhSlhVvGWeICkLLboBmP/5gw
Iu5oBY0/jcY7Z+zwep7SSb8UQX5EmLBxiR9QqSXzxtekf8wrwnr0w5nyMwGHQud0
7NhAo6SbnHr2GayhiCVQs0HYnId9m4IYlZ38vzG5rNHE+92QCfxzPgb0AwrIx0hh
beFF1QzyvhL+TwQ7L1Z5JgG03J1nodGtbcsi+cd39E+C7zVdMPJPFnCOgiKKPEfT
n4Y86PYlKYumYSgQpwHPdG3ZyrjfeXhIcbRIR+OT6lfvd8Y3WaZ7FDOrWCJjksFh
0QKR5kn5yq7phheneRRfePOzfcBlE7evsHPMu5PtrYEBrPgZJ30lHFWDaOKv8kqv
UeLVtxvOHO3X5mZx8zFjMIPLDMdRN+TGal/qwM63sgNMvAWJwGewmpzJXyOXC5Rj
T++584qeXREfI4L5a7To6UpAwhiZJ8f/cUTRt91zUgIfLHc6uo+q0/UfQWcl4oaG
2feFbUgh2AoKnhZwi4Y0CeQprN7VXcUZ3SlxwfsdOYz8Yj3SQvLRwM9JratimTDN
x+Kf5Rolt6LJORI9kz6nZ+tndobJdcLPOz/h6qEnyp9AP4SQcF3WWluyqQq2ZVrj
+U4ZvWuUb/EqmkbR++C4uaUH18oP9HYvJrLSOlZmVaWim28XOHJvQyontQgEamHV
w3hG+dglc63uOMqND6SOy2h6RL0wRNGG8NNctAtumjUKgOwVhbMe/7O4kgqTP73E
Ivi3rBRnZ39cJPTaRvzHDm3FJYLxt4IjHQmSGWQ6+b8xKzYg0qSJDI/l86j48yM+
hrGdCe6KRb+bGZmdkfMDqboXk22NZOqDB6ZjfdDwWv39938ufKfKOWhupLoyVbDQ
udRda6v+axwpB0YpqigV+sWQSPaemtixXU8W9O0hfq/wS08P2krOwjkzgXE2rjfs
/bTpWlP5L6GTiDGwA/1lhE+1s0wcFPN2kRRBP3JLD6ermVkPq9GrbQkmb1ivoAQx
Vu+xpdNzimDM1FiHCSew8iDTV/YK7AWS/fvpd8UahA16QdA12H40zACT/v2JA34B
NMeCOltgrU+YWRNO6P/gnA3hfF8dPUYauOvqwRgK5KVfLc8VX/AvCejqP0oMphWA
aW+4STOmoJDongL+XSP1uQKYHcF4pKp8Pj3kILOgP+i4HKwkjqVMt2iU0I7/0JtW
TAG4vIIfF8BzrRMpR8CjEoe66J2w9R/G7N1PmuqJfGHnR9C2sECe6KpUkEtL9DZS
NWh7xn5ovnerKwtn+8Z8pm5ZCwtnuE3k1d9bIGBVIA4BMKoUbjjX8o9crspJCOM1
PJ+U1EDUMMVfIgkU7tvqbXYrle+wB4mNFXoXecP/haw+BcSuLFFTJeJKIy+BwqTj
aqnZsxPPDL8zKXliTvLo54f0RMgmdP1lfvIJh1Q8mj67cXwi3OUGuEK+YRyzjavl
j4Be7Ri83d7RbtL/ulkP473hkNJ5yPcbmDDIlDGK4d61Avm6Q6MMXYuOdldhICU8
q7eHxBupwn8Ic4aR64khpxZ0HVhofjgqCm9lv5Hld5yP/42nc4nMZ9Vpn4gYpd0f
yteeUwByDX9dgc9cJC6XOAk2vjt+fyAqkarovkEyuR9TbQ62EYHuxQKkJbDuF+Y0
TCqkjljcycvipDdZPltlXbsV/rFGjPAg7KAl7FyBIVah22NLfkUb47fEwr/aEOwf
1HPwtjmKSO8cqp5EMobC2ZVYdm/R8iGS/d+pEIUliUJic8CIIYxpsT3X839g/bCh
m4semd4z3J6mELuu60lHbTGW5uFSixFpnE7SsIBcpz8FcBEDBQTtXzXTiJE5RPO5
d4ONmcix7sHqiHbE5DCqnY/yMpLHqAI8AZ9/DEvh1hw=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dODUcaR1nETuspj/gZCjSOS/sq4C1jc5HEGdJk+0u09u0eZ6ZRfMlnQ+qf6lt+uo
wVa5UKwSA51Ajfrdy5ry+arlzHezbzceaED0vqhxR6Y7e0MXnzISpkSzO9aqyuwd
nkcM2S9PGFHDHH3gnIMcv6t+1xRweRxw6+uJmUe6tQzHIXumt5fVMWhF6JlvDx28
yTTGBp0VUbC1dVAA4MXMpYpWf1VyW/GEztSYllWe3ZzXre6ZhAs1QztljJ65vAzq
rAnNJx47Of0e0qbtdM+VshXt1a1fTg0XpGSG3Eu3hrMBytFgh+QJ3D7PzgAO735Q
j4AOem+hqjylELzPYqCdaQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
0qequHUEW6B1Yx0+ewJgMCORN3EtIbTYbQ66NhSb1Goj7hOCeYnUyprWnthpkCha
pR46k7mRNJ7L0FZOGWSl0g+o7sImqc3HtGml4y7gCccnfboVmYjba+Zg9BvTbtmh
ij352qAB7E3Fh+JuFaNS184Px0jP+uLDmPrpTAGNLqJCDJfVTAfMQ9jyeKQnpsYY
EAPHJvsL1uNvD9Iu3Gdpi/XEqC1DQdMuqSl353ypg0ibusFEIEZ466p1Rwv85TQt
VMRjEmFwPfCPTcGdtq0kfXZCANqEa2VtfVk93pB1vdCoC7A8Lt6J7jQCk9X3WTFH
TWEXcloyv+5pPVAu8dwGfFBt5sJis1fj+gR24QE0NvXFr/bGmXPE8NP3yuIxX5i2
uyQ/UPh9QZqnFXpGcSXRDRIdnUBiiU9+FyqYfDc7tj9rsx4F+g/MZL3KLRrAN3jm
V0H268pjB1j/nK3kAzWqYtlpVWqP8uq6QKPtvYGaoirlW/ZY9xeUGV92c8swgQ08
eyLUxslPaw3HCgH+yNwbMMkY0AVIAz6DyUgyCBNcbjK8ANoA65HMbg/hf8sXN+O1
1DHmphz8MFzXRj2rcd9aycobWNEVzzZtW7kOSOBJXS2mvnRvRuQs212uITmuQcvf
DNNU/sg8YordzKVx6wwRzKnwlLrKXR9tK+mR/sne07X+TwzmRLauezPBlnuZIlsp
l5Td2WZJh0MApsE9J/DArmyMapXsL9yP17wReVi+zCfb6WgwoKZzDsA3Amz7I2vp
QvfWlzZ6qK/d2wNurtlKTTa19Js9yX2KTma0GNO5RdGyeABeYjwtyZx+4G7yHwSs
m5COsytj+p+lwlTnFCEwuZ9PcFpde52FoujOTS3m3ld91QhRIQEsQN65w/4oyK9o
IfHUaQtuwDercaiE5x7HKG210IOyuzhjPuHXFjkD36DQxadgS8Y6mEvhSxeMOSQn
fADIlq0DIVNOtrnYITuI8B9Bu0X/ZSOxdxpiMyjOZV9AHEW/Zb7m/Uyk+kxw/9TH
0lTrEh3ZP4E9GFheYHd53Dna7kz0ZndLilWuEzojyUUXH0g/VAf/nMIXAb7Wv3ne
QB0Gq8xndODBZnPllsxGgR4WAsNwaGkfN7SVKwfRP/iDJryrRSsw2X1ITPRHlUQc
A+UdwoTZq6ePtzRAFhAu4ncfsi6UHc0NDna8x9oh0MxHuixf1uuE0OvXW7F5+bmS
9uKHn7llQB9ZIlPQFUx4DdcKxcq+36FMJvPeCAa8mFokkOsOaTbTOIFxKauqqwr7
5R6NZXL7pqdL2faceQmhB+4UH35Va9dROcbThjocyDjaBxmk9MTlV15xU8Mi/e+b
r9cY9d5PCJTjh8JMQEnM9hOYLoNav9cWY2+TyJAMwYlVQPiHANvzAKu7via2swja
+1jx5eUl40IObzUyL5E7FWM7MFg/+BVnMl2ZSQJgLIaGzt25Pjebex7/fRMOpm+5
lR9K2JB8uPYQcixNTjxaysfJgsxG2QQq9Q+avsBGQGphM3FFWHd1dtFAa37Zvz7E
p4rK6EaMYPdXtHrguI38KLBYajFuAXD4Au0g9+T7J6AcvhnUeWi/UrPEoDQuajOi
b7IQXAWxYg74QextCm3GK60vUo9nH5nPmRKR3s4sEvHyubkih1tG9BnbJZN+bpjC
GqmkP9495Pwi2omvyR0PGTgt1FvpXFOvEJ9aXy+flWABRN66CQaOWr0KqakAaesf
kxmgFFMT1Zp8TVv5i4BiGNZIpm/YrxWrkHAgEu4FZ/NGj9z7vvFLfOryHuQoHDIu
GC7JGLrxbhfUW/si/5WW5RrHc13AOEWZwblVSrY5fcn8dSYizqcRbWnOuTgGTb3z
KP9EW1pprlpqyL4BHJAHfGFC+E4R7w0dsiCqMpiLsuFtbnR3hIIFjiOGB2SZCL2k
IWyNzR/nbrk6bHj99mkqmxQhguNm1dC7Fv+vtj+xPuEIlTOhE4NGnYFaKKGwQdbr
7WCoHJwQrq6efT4pgMVtEL01pKJcfA/Ii3R87DkPSnJtQRzmV9ma5Aep3aCKBzKz
2nl5PQ9oSRjqWjpgEUru+fM0Obm+zApP6Ptxout41sehoPJAIr9Y0NtYOuYAxngY
UuV5/pjfqC4nK7n9jrnh+A+LOko4OMe1Zq4ugLShegkJTFtvzbW5eHhFPdwOB4W0
TQoSm1KaLTHhgFAQoUZ+oJTmFGjX17x+f0Lmn93vulcRDpm1Hkcowx8jokzh0s0q
4L0I39fAe8BeNCHZi7U4aEg4uX4flxweT/wIKj1S2kg81ZL3sZ0m1dTe0O9BgO5B
0ruS+SKj0Xx7ymm972HIAlB4670xVfV1nrCJdcgsIOjpJ5u8qjqqOCn7yvjWtexx
ddll3kb83KVJe2ftUcpAwf1sZ9Hz7aJv5y878rR3wJUZzDYghZL9QNJr/o60OQxj
oMb3O6HjL1LRRq7Qd04S8CFkBsmESwcIUYU+XFUCxFHri3flSgUEIuSdXK3jkEvu
5cnExuck+HBlbbNLQ1Rzq96KOmZMznZr9Gcsj/mV46t9bh3o44KStRMUS+liR4eo
eAgkZBpD18mByEDTm3/w3/ZR3qOoynTvl91msH7lKE3RErmnTI42fyjpNaqNl985
lR7YrkwD09cZA88YgRk4J18P02lTY5OCPtfxIEOz1lq234SsCZeAIiufCqu7VizD
re2d7lNqM67UmEndWHa1gWkDZny7TLMshGtlpny9cTxcCCo7VV2uUZGcLJw4ljyp
GxIQfowrNMvu3KpmHXmKUbhGaIzgFiLLWO7FrteZjFwUhaaCtW6QCyhU04arHX2/
Elg9bYKRp5jko22npAgEoxKvPThlJirRQT8hO+lcVDN3dxeEI1K7Pmlda63CmK25
8IqR11KeT71j/L2QJToxGTSrKu2QqIVLs/mLY84iNDzbM3gF1fWwhH9iFY7CCgNU
dnTgNsVfOUxzVZ7nyT6GW1rubsfAStQsaMcJpOMQchLv/E3E+gfc3V69MF5Qxfi5
LTvCQnadYOigLn30QJKiwTT5pghaNUqNsjXY/99A7mKqQ7TtGqv81QZwZUP6qNaz
xoUaIYsNmVOY+z3FLKmUrVGg8UxYSO24pJa8o5+eNvsAJXxf8VDk9EHVx5Y3pima
x+Op3IQO3XOOjW2QjLWwK88bHv0Pvk6KNXIMhkkxC3FtVeq5HFkL/BNRBlLMBFEs
ZGuQ91zwyVESlqMrXh1U4kIOD8GLG72fM3snyACSRSEkL/gaUqOk13pl/oxeHp5T
AWYyMagj9aUlJIve8KftpNQxvUSajsnKvhw4JoysNpsfH7rbXpHAdFyn7yOvr+fC
29emn08RZhZociAK70Ou5EysTBWIQxRlaatLxHoQkkiDaoeBIXGUAhcAUHoDD6sH
4sSPeyvc5/YKVxksX0r59TyLPQmaR3VgOFI3jlWDglQ8vyaC/s2J5OJBNJWdagi4
2vfXWr7CUsfpNE5BRoYFN9HXdKKkbevDxeLmfNXoMHQBFAelbWMy5+GeXNPsQx9x
Mw0b3jxg0EbmcUQ2Cx5Iv1UE0L4szSGksE86tO52oas0WHu6GtkTk7a/3NyZzmT7
OmPC+UZLYYfolpYFLWSy6Cy0Bm2675Q3NfWZHoYPjN9Dh8dly/C7wKY4l2wI8F5D
ZKKBBliBAYLoZit5Ueh4MEJg8PPZ1a/EXkqohur+eQ4v+3xEkTcc6HRsdv6dQzzk
65+LA2BGiYzfIeZ7luKUP4Z/mc7bYnPuPYPHT+FkC0xVD69DMrSXqEXb4dm0n6rz
SaCSaD4dWRtOfh23jG5N/VwF3/DXCk0kERFPfar1See0t3/KE9WSpArB/UCgUCF2
g9VtHkLeqHqbHYnNQMJoBtMeRG9geRms573MyEdW/vDEXqOAbKCRm7ewNGn1DmM0
Exgq0QanG5c1kjDMIbpookCFYekEBrsadukvX32QajNrLKPOq+O8KywuG6PLjYcb
vGQmtqw/RUm47eOX1LryU4KokcXkx6GpG0MW8I31rBhpHOKtU6oTspmwdoHIErSO
Hwi6wcmi0oQ79/f9AqV7TqoVc0LFkhxHcjutARoLBP+OjyBCWusnMRgUSFmDtqQ9
1nsfqK8r2gL68q4SHi+bLGGOX3qCVR//lxmTnqtCWA+Esee7kvKXD8xFuu4LUqMa
Y9qYvBiGEgVVb4gx4g06fcWXrH4xGRDpUItmMT/GjvRVLYlQD/0XrezlVnHqJlhY
RT+hEfSv1h/VW9ssTU49/DnigRQsS2A4enh/Te/q8CGhmkmqiPVp/04lUTYuIdvW
tlIhfIevaHrKmuWGpYnYyrFwfGxR0b1YIImy/2hiqNDty4puaBKrF2PMy/Q8NNP5
HVti+PA73ne7bxIXNxKxOebmvS9zphOyxU7Xpzox8Tvo6ocqXUmYzmqpDdQbi1Rz
hmuuhAInJ6itWs6uAiKLXoiEcrb8W2N7e5s8Z6c7w+PCmwHscfLAdRf15eu6f5eH
oIfLhHDcuc330taw3TPvXRf5CWkbZ9eD7k2rXGZrE62eHlbfrRfzya0+WWeHEITV
ud3Lh66voTJBZdbGqK7IKWVYUdiqjdQyvo/NvrjUemg8jGoVHatSddCsiI8zv/Kl
7rOrWAds0pUMy/Gzgp0baTS+5MSBHMxROxvjFW20cLWaTA9mfmnB4c1QflPqOHDc
92BfIDjqu9ms45zbxc9qDVzDhwdE4741RZSjBvpe3S4NtcvV82v2X65oFK014a7x
XAXZmqWFAYw4768uD1hoPOHmmzG+z117hrvvwLhTtvnBvpX2UBTbDUj4I1YgwPCp
qVx7lfxRdIG3c0AhsVBiP+2wFE0+WwSvUkdxv0B2bNsXwyFTC2nT+L9dkinlZsPu
4VEjETf8bXu1dKiBcX1xByZGRiWWy5WvDvYgJ8l09IYoTB5hr6A69/cnoxxuM6ki
R5odyAb3rx/sgehcWiKbqHeGmkgejRFFGVNDo8sRK1sXA6RYb2Z5pYiLqElJDaXt
mNWadz8Qpci9YbtpNOFDBp+AuRgBKaFg/Ow/Nes0AaAlr8+5tDk4yXnbdDSkjePG
H8aH2TNRTd7xMyYI4KuBbWkv4odwSKjbwt29q1TQi8ViSOAsQpp/IYJjvTzxr+4f
M4P6apr3UbbZ8eJERW8AXfOuy9iWedPQ8OeQ+yE0XyhzXGKnALXpQMcpQQF5mDoQ
YZB81Dvi1uFg0n/ERQjciCLlxiM+IQGewN9VInX4ipMTmxa0xAUT8jEJq/XCFmB3
iWEDZoKVnisTB1PpNE25uieq8bdyHTK19nl7UOalyDWrpYnfATxai6iZTPIdmaFW
I6lDoOow3ZggFg+Z77ytJ8g9kWZJ/gS735xt43YxEC47gFBbkx7rTv7BSjgOjW5E
RjmJXBzw6fBrg8ywdYdDkPnYyauwB8sLXJH/ZBB8kNkVup60s4/X9si64CPX6jUd
+NzFQXpyHG2ocXYROERqcnse+tqC+kdTBhh9CqGdzPzmkmCo/M5nvStXVY6h8EBK
f7zuckzgGBlXRoqnQQltLzRXa5mTlTAstO+k+WJk08nhhiwPHY/NvAwNXCoVtUb7
gGSWu9JRc4cHM1MlDKiymRapo6QQBgGMy/v7H4dhoZjncDEy9+DwoFZj4rsbU4pE
w7Y5fWphDwwfR0EBoTwgvMWIuyxBiUr8tPqA8vSBaPhWJyMhLVYLWskCGfowqbYz
RA8WqRx6n7MEF8WeJ8gZDApCleEUZDNekLYpcGMzQhxEUvAqvW+BNfoZj+cJap5+
MDAGji5YF+vl7lmuH/6MlLMpL2p7F1zXalmJB+MbXaBrU6fRTkLx1Ms7EmgtQK9I
kS3v6bXpoxv0Wnc9sAnFUThIPrOkFl4+t5+6ftG/AyOW0c2ToUo55R5GJ1iVA8fq
HHutZA6faNUKjEccieLDUeSBDwK3LH+buoErOOxMER7QpG9zbhSStsuYgcYtC3CS
Qjm5NJI2s3TEa9pgiYypM26l/HgjT4/3TgxTkvMVCFdOs6YY7E5ywd86NVxcabXE
xpjGa91xIkPvLkohZyhAnnvkWYx5eh4ChRXKKygVQxX1DQSYLNS+XposCktZgcPI
cALxgszbPt161CQEpM4s+k+b64cQp1GofQUXB6Cr/W73uk0ZRil3YXsAVUMficyD
ApG9SqKLtSk4MS4RKl679/pwV7P6zP2h9Qk0CvEEcLQ3VJvvpe4jFlP7I7e1XYu8
Zy5mcWp5pdbn3nEDlmy0B39Km/+iHCaQl6gXrfIHqT9xdPejUdLKNOvwARqYdEWg
dDc4czWxTpSbXyxFoBlNUsGMGWyym1KYpDO6i1kcyrS4d/YrNjQPupMSWzGcGjjv
/7cWAy6KttGtFv4xHWISkCVTCODsnt8M9oPWGAT1aglv6x3y/TKc6xmmfotiZlIz
bKuYdpZOGZ192D8QZhTrJkbC9lHaVHP+3jqeRfMFN5/UWWFE0d9ggijKQS2TtuNV
RdqalmDaePs/cpu5T/CBWajeCFgGaOU5mJ82DTUea7qVZ/1yX5zxDjQ+jUFlFvz+
bxoQ32aGwWY33nE32zr+tlAzMMORoFp0bpOdLGovxScgUlRPabKrqgqI57o1NLBi
5wanQsoNQGyJfbUlR15ROivh2ju069WFRjUMC5Ay1UM6RCiQ37YEbaqw91P0iASH
fethd92lNWk464Mb1MoAJ3rDulkQT9ckFxZsc7baphNHsXjKQ8bYngS4UVJqRxsf
IQVEWfDZljw2OvpjdAWyLvOQ9k4SrYORyS088IASE9klujyeRHMAtwT3RWIfS/Am
wyrlXLLp2Jwq7WxSMUB+BZICyTXD674bS7oskpjWubu2vhM+9Zhlcrt66AKrZ1Fa
pP2etopS4Yfcm95KEDg3vkqoR+lf7fNSPIF1DAi+Oyyu/t22ldFNdSdB76U1nCJd
zVoLDHknfLZCl4+gE1a5uixjRf9G+aP+UhdgS2HuyFQLAncSu4XsCdCSxUe6OOgG
waOPCDcReB4UPGLiLvk/EqYgeZSGvTsupr0lWrFZi4geiCZrnTabrHg3gQ2T2ZuE
CUNIpHavVEjNnnp0gDQPem8wUiFZHY2XxFj59REFIRjMyUgmQxCCWVkAjnI7XVnT
QvlpONdSdLTRBM742+Eccx2OsaHgWVi5pW0fvcOYIJYHbsrBnYpm2xpGcWM7UTcO
NdjMeQSlVZSpKpSRLwFo9aCXH3U/6+Lc56jQNLNN1MIKCLZZuj2NcF6pEf9YAzvw
fNXkknzmsd7C0bqQAbCNRXlFCKCinWawDucEWbf5XzgXxmnQuZ9XcIrrOvgRZX+y
MU7kEwlyioCL0j9m/Mdl1QLEZ0rcLh7yGNOlgy71eD5hY83LhfNiZFnvthqybBV+
Nlzkss9qycQWjEHYo0FtwcZbA1uJLA79r92uC0XFTje94+PBGzk6g4AJ0lREk9Vs
pVDnJYls2QfJSOinOqTv/XUaJcaPgDZkBf8JA8/lXR8bPVmSz68yt4BSwWGBjeCI
JaT3PbpEE6dI8hZ1MfuVt8gA6muka4VPFEasYpIHdkEfSAMl7INz8ukYXOAm1u1e
HW7ktNxxzSrNwJIOnh4BgkU7ltjF4zEznabj0ISzgSsGoPiC5h6rO5nZDHEkSLsN
4XD+uSX5pLnFyMTkUsLII7xwSDiP1wr8WomjOw18YSSLwr5ID57Jv0d1+zzSBvmz
XvRFZDFalw8yxfUCsNDVyV1AaMPEKkpvJ2TeFMdaq3deJUvZ2J8gO79OR2VhJUUV
TTbQYS/uvUt/xejW3g83qoi8IXsD2ISHC8rc4S3EAAQQlWC7kjT+y/uvWkoeSars
if+/KypWW8/0zr9dUKS9V5HEkZ3JjkM723O6/2ooAj4GEK9feQWydr7fG46z1PAt
BbqkRRXkuWU/TA8oPQrsme9qyp8PIl4xm+xB78hkZod5lW9q/1eSc/J6uJotD7sq
m4GcslJz4bB1X0M2ObBmjf1DZDfYRQZ397uXZ0Yt0Y3Nho6VykinUp9Coz7W/086
skS/NfsBn65Eka2tAqOfhjTGRNexW8d2XO4p+2qGJISNR0E5QnrtYfMiQWsAt9GY
n5rGE3hGitfxF3zTGzUvc/YbU2wY8aFrl1AoLYvsR9q63A66itTyRPsjFTfGXJTl
u6gA/HPvGepNRTdgtnioZfQejR/BOrD5HL7XB4X2q2AKXo4PkwiX2aqt89pKwm1Q
HYjp2yYEQ5INHUuwJkAhtcE68IH5ZNnU1CTOHYAnbXUm6SjuuIGiPst6ZXorE0it
Rwvmh5Y+R1H62GlTwRrK5g4u7auL2vPe4YVwAl/F9yhn5CHbTjAhtrgv5AvZ38Wo
ZA7FWvfDCsdxMTcDbVpcIpBTuKCBdXkJPQgRve81NOKflpHdN6fKzdollpe7QQJ+
bqWzI8MR0CrC7fMX88P2to9nXI4W57jFoVFDI5g/EBbRdi9kubSmtigJXKH9j7uH
pCR6c0vx42WNG6gaa1K/2qwxYF03JnRwC2c1g/gdrBbfuMYXuGqIXAEPCLFumyuN
IDW5Qp+bg+QXzNkf6YyVaYym4qQp2dexFcgM7q4kRwcazI0uq+iVNPcqfPrMYKxg
7hfm1kII437CEFNVkXXyHTWWCvwudL75DjWTzrqExt+LdQx3+rtONgu9e7tdqqSW
upACQFAra/sdVBxxqrWaQ1/OGM/IOuLp+VlNDKIuYyea8NKdiMmtWwUXvFzi8YFf
bbXafgaUDgz9D89+9JWAjf7mCvyF6QWZSFl6L43WpnyYx2mqUm1hLrdOjXbPrezO
83fGuUeTyWY0Y95d2Ek05cIwOTP7zOfD5G/olKXXTbAAbLIgYUG/m0D0pojsSS2x
dIqzSp3ZFowaeYrdWW/MNgzglrpfcAjTe7zr1rG+JaDbsiyUxPBvJ4LI6bBmBh8Q
biHT2dDpwejhgif8weo/lVMsNH+648wJECFg0x9GfWrdgaBzUhnc3a9u+7te6C2g
Ay9w99zfPNdX+cOhkXzHOt75T++WNSzCfzSjK0dBqDierGjgwghOWr2cDpet8Ic2
N2eJh7YrvESp08PzbYN+/qFiUbZGfELH4hN7GIiQ5lUuSSZ8OMmv2djkAc9ttG/S
NF+GTGsTtuaFCoA1JaDcoWdIIWNjk6CYzK7sFxaFaMdich/5/q40idEzntLS+tI3
xhLQibBclpZHWipAiuFBlA6/iAof9MeeewlgpZwROJI0aJZCaBLhey2Yo/YVtEjg
PbZNlT4ZXLS6YyShWcCdhOFv6Ylzk0iUAnoXhEZ6T2RK2GWXBaCzKNclHITcDPXZ
FI37JoWQV8wUi0HK1uTwK69/HK3g86+VXsCgMIMYJ3/3Lzel8Jb3vmmoMauY8auv
yyoJuaNOY3fV6LEvP+YsMUWOe5EAtRGKdhEzL0WmmWAOwteE/lhkUlKZhseI9t0y
ncVGciI2fgM9qrL8ypT4dlDzf/ythH9OVfB8j+NwT4UQ4+UnM2lxasdlXuYGnWEw
7gxphWmYOhHi6dUV0z5u4eZwPf+4a0FR+ZHWQsX7qK26dhDE09BwqImpYSiCoRrV
pAkR1UoglOaWBADS2TIqy5DaCZJa0ilO8uch9RUkBRnAOd9BnIs0HtB9ghh8AXD2
MEQIyiDjxr5jE9hxqJ0bNrtXSjAw+MQfQoYTQ0w1g9raZcc/aO0vMnL7ZdZS65rW
PJVJyqH+kAZqb2LIrrefuPDgL4xdPZ+xECn005gT9pwBs8SEVKp+9ECCQwTXhXCY
bZMsfT8IO0TJARQAt/VBeknZlphEF5YDDC5f6D0UWxNOPjpHaAsoH2a2po2tE4xu
U1CfhwgRRyslbtoDPJWhfTfQi2a/ItXkepF71zEuv+na1Z0ioJAr/EC0AP4SUK7P
YuEf3NXKAGp+sd/jH4rv/mMKxdQjpXoJmEXbpMKMv37Zb0kkKUPmcak2zgCVotGg
LGjCAYjHYa1D7Wc9tBNNcEHLwh2jYjGxHEEZlF/MJ/fZCt2P6Xokr3tGffeGTMPr
wsjT2tQkfbqood2m9FEwqzZKlb+AjBDqoZTLUKZ1ll8tov6QBIlrHahm0j9IC/F4
AlVq8Wg6lQ2jg1lllE+dc9UBEJVk7O7L3YCLtHtEtiEsP99a43V/EI9nreobxfPk
zN9E+vwjo8xokIAQZ6gPwRBNEc9xUVrDKqfH+emtVrWivnrkrhKpMnTwquo2DYIP
4A5GCBEQaGBlVQwUN51U0GrjwpEvIZU0s+x/wtAyC3ecJu759AedVVYag33soKr7
L/6a+qkoz7uXEJQb9rS7DsReGlDGgceDnQ2beP/pNpV7alE+eNX82qf47Ss7zuZi
45R3LO139TfZvtNdQ8Zpw2P6B+3zQlGwLrbCb1GxvohfQzUt3e4Jq1Rc4BzZZCqV
xENQTa+Iu994LR6534Ps//5RQr7F9rkP0PXjykTWU3W2jOY0gZ/0/+AwTZLKNkmd
rR6Ku0SOppnc8pu1aMrpYvAvIjvi8WeUTFn0/xK9Xgy4A13iTmKBs8d48+Xg9KhN
eHQsWW+e4P4PBHJGJ4QUAng8dSt6c4wxLaAm4ymLoykVwSk/n+rYb6z33Pm2+NGl
vU2/xPU/yTEp78UsLS51LfLEsgX+LZtXq4oAcThEJmGNnR2Sa5p9Shiym1XFSO6v
84oJ1lco60gxGiDJNAqRlXB3ErqWmsWizyz4hHwreyRf8CytJENJefuomWaDnN/m
YARpSqGgbgOe5syiKF2yLDgEVB5vvNzxNrUC+D84sCmYVBLR1Y4uTH3CWsdoWv2w
cs2YcrY0ni0FlKeHE3XjbkiwGvs1cRJ5r8SbCUOFb5qZ89FoDXghMs6aQGgdbcwx
Vye/30PdRao0fysZGQdwEGM6/GVMLadLWDPAK5SszOFO6m+Rtnn6UaSFdQG4E2aO
N38rsQ55bOxzjTZ4tCZVHbeQXbhXnnQvwRxWnnHfeWnZjX3c7U3eK5bv4WsDkBO3
5ivaUGHMUDrax6W+DtSlu/H43Gafhz7HM3JDhTBmZ0Q8ZTL2MuK5N3GqbNqy9dsN
FUALltzDADSCwOdrHywMCCLNMaoeZHnbzBN1wp5feAGezQyc08kvrdxZDgudbmYs
tIgADrtjUqCRJGu02b4cCp8aeRc3lzze/RXGLYra9yARyxgQXzr7f+xh6sVtOXsY
eYFAxBNOXqJsGvHZSeOHOQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
eBKLpC0GRlOSkrTltFFy+M9jUoSN6TH7wxaic8yEBr0oYJG3OiDeRE1VO/GlN4oA
kz16aILtsIwy48rWxK0ItKfip5HXK9RGzCs+JE3djy49kJpPFDeYjo5WZ7E4/N/9
gr36amcGIQ5yFKsF9kIpLvHiGhRnnqrONK7CBsR4ckb1mWA3AWIcV77gK+9hBpYf
DST4AhN5dWnxULQ0syjpX+d0E3XUQTLuYBcd06XweXjWft4ORsIha3SORwnVHB+J
HC6J6HryOTXPrtBo9jI3B1fmU+5hagrp3cB2lLFdHHu7yOblsxMqglM/Q8zkg3+u
ZJO3uVKhjho3ITO6tiorEw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11952 )
`pragma protect data_block
f/WJ+2efYl+DjgCrWqNGmv8qyiMYkADErXOfpk7FDIPMujKLo+rlZHnb4QWq0UjB
vdYtPk3+H98+CA4izSipuZIaHNy37ZIU5ozsdwC9nXMlSAQ59ZdS2yumQpND050y
G4T8MYOyXKl6V+LY1fthpGJ15vAOVCxoZeWQ4zOGIYuK68nZd1f5tYrsvdIuXIt7
ngtxOvwg0Hm8w2fjitKVHDAzt3ksK3Cq+tX+tFpSBmfkNCCSEiAciQ4zeA3YJKDU
nIkJXuPirtp1AD+tis9oPrgiY8w7/kDg+L0e0O7CFpb3J9YgTmtUQPgfDntdq+zQ
MgevrBM94ZskwWfTCsXY9loHC/My7jOhG2p/DN0ChL6C4FuBdxAioqxVZkfxrYwC
dhvO83rx5gB6hIjQRya4SE+L4pb8eH4uAuc3xFRFGsJcmGVkYeDtSs1OCMdBq7Ha
+8sZXkPVsQUDl3Sf3rDu1/Bn+bmm9McsDiqTIFAQ7Twk+LjPs9fy5Tenv+JALwB7
a/Kh1w1LqRfAwRiIRH5464ORdQ1eaZsnTzqzaxiw+IgcAYFFLYeWWWfAONLr2u+4
Bt8vdFnWQvDQ2nrShKgViwF8W9SAt5tMmr5emUdlHne9RCTu+88z93dCt2bmS8TK
FwpY3LW9rZ8QdfWI0DkWriRfYqcNcXw96X2csRPfOV4Wr6rjJK+/4PHjXxIScZqD
LX6VDZcFZwVOIot1raft/1Vzv5AzdCwLq+IyatasbXnYi8nsD6tpqXRYIUskqr6F
4qOAXd1VqofJGmUbQxHB8gxeEeW6o3DIJng6PpGPIHmRDDjA72giypOOX58ch4so
xWmUm9VyZdgN0QcMAQS17Q833x6X7nVraDjoIg6Ljq4NMCSSLCQeMwYiIigvWAyP
u7z2eG6NQAMoYKytKasLRfhiRQpNNcCaxMC8TSYrglh5fbLTTucGrHh/nZ86xp+6
GAPT+Tdtwc3XwQXoAW4nA71K3FXj0c/5VwT7FV7UGlrffiNT5Y9nNvXLTMqrCd0b
rxczcXLtMwYbgacWxGTGuMmj1erL1t8e+o1L9H9xaswDbEtSitv9nLme7hLmOPfu
xkKKhYXFhLfBNXAX4jaP4pYEySJedZY36dEXv5JMeFqM2DtsDZmku6VG2Rks69Q+
CDkD9xzqIgqlTZslb96eEkigtK+u9zGwa1OwiBXwXfR/9E+xdEpsLWW4AsAHNkhr
8/rEEUvUYysgTNGG161SIXW5Vi3SasS4W+XbutN4LyuZiSCajkFhleZtvOYkA1T+
n1k8KL2mwuLwR3SmjEnkNsnHWjuwviHqaRWXZafxkHEwlRHcziSeei7ORzBY9kac
6JR2QXnzcqtshVdgIjcZhKfpsuxQ8ITW5REjv21X06L/vGcIh85qT1kMy2elYGSe
6fnfvHf+x+przr7iiY3LkHWc7RMrcSSgFGu8t+8jcyhjrng7yUgKgbbqKvhdO6x4
0tKK1pL4pPxdVQOT8B7IX3P6lwJ1pMBFooIannJeEjUAdstgu8y1lxMMCgu1x9i9
PjmGAA3rJup0a6I+fdl85lmdVF1KvMyQOmw2gQE4vHY9aJWRGQSxJhcaDJaE2n4Y
VM+wqZyidJ4ULQcZ/evQfJiu2SyfjQB5NmBGurplqapau7fiwTkKl3GW0qtt+J4Z
mFYvx+Uw0KhG6GFkw9SO5ZnlGTt6xpPkGN2pZdk8TGHVucswTEami3mKIO+pbxnt
vBOyX6vNAy3XZRwdFZlBKXvEnWHFVnV9tfpk8q1Gm50OAU6JuZoQm96YbD2EaYZV
jV+832fI4dBjXD8h1xoK3XLXP7U5Ocd9oAkw+fpYgoY6a/qMb92W/0MDzBiETVsK
DlG6wz4lS5Y1NB4L1YazJNbuAFf8dMIlBnuAqcJ0uu0YrjQt0am1HTOgPGPRRLAw
af3FncHIfU9dqrEcVa1nuGf8kQnTzIMA0dR071M+8xgF9Qf/NDyuDvL297FAdQaz
db28uSWRdSEhvcuUCppYnv9W3tKQl3J5i1fRTa5xx+pluYoqOFi7zsfISOGNx07O
3BZlJkTqvXNMySQG+9fz1Kg1uFW3JYn/fJJExQL8WwdSVvaNqp4+PIlS4Ek9mgvd
NfKint7kWvoFMG0pi9GrpcdKLjSHPe01wuWvxn7M+t4NPr5yv+rDEUZ9lbyIvx2d
eo6k5/NWD9Wj5NclxPzQCmKlSoJLCFIu1dHdh+GA/niFTV0AEkAiCLWBPRtQgAsN
ATgS1x0kxxyzyxz+2Ug4lwfNwzgin3o29vF4JD2DwmultOKygHCCleOzsnV5BBka
D+Cbmmm00Qau3EM57uJCBYstS+jlPnBbY4YF6XYqqf4dOPlYqQbvYIhTeM83EXC5
oDTgq5do/hdqyRJhgNsyfPKFPp4XHqmcPowHcJ1qZ3Bi8jfi5e6lr61iDTiP44d/
K8lNz6oKXlEdmEPiXbj1mRS2PzS1hogHNGyfAK/+uw13AgoRIZiMalWhd3ekUDns
tZOuUMJyGO0abacCdTLW6znL6CXrxRw6YZNlAfVzWbU8QtpGzJYGBcn1P3LWtE2/
hDt/MnQJ/Ls2HOuDuGBaqY6K7LSZYw/fRMq/WnF4DxUf9K0CJYs4Y6nt4t6ydyoP
HlbM5ggE15sLDD8rZ/OHb3vq8MPtzJFeuhUkgsIVk4/z2ogDv7GhHBs32hHcJAgj
9iwAXl4OYstkFpjAZcfOyf0usAOFPq1TlSEOvh9ll3odLlVTJMXWF8IfxPCKy0rE
BvgzQHEixyYckb2dXW/fq8h6tYwpuWZC6EqXFyz3VfkaJo2ZdFnF8VKlICOVo9R2
ocjwE2BJi4/pxzATHP5F5k73gNidwiGiGomWWkA631HkN7UJsOcyRb3IHpkD9QPP
owrM6CQ6HUon1vN/+xF2R41Ni0DTclBNVMywg/g8Efu7kNqafscTRxJEuQxI4yyu
YtBKVTyYM2LAS/Yw3ePfz3YerhFUi4oINOqkanhyc8WYeSy3Ypl/EJaXPL1yrGOF
T+wiOYoF2hMLBHuePMHakzDiFWLwAaGyd8i2xviErR49YlQQmdkQx2YwtTgPFSv0
c/w9HPKmP03PsiFERhrs+wDxml4wOXRW/R2SZjFwh+bVm5EtOwG3rIXWO2x5LIrT
GaxGR2IgjK5zIw/d27Dwfr9HrYEErmf96ZaplHXXoFCYp1lZ/zQvC8T22KnjJqlG
f4Yo8twD3V9lxnNr0qPGQu8FeaZW5wi67nFF1o59j/ImsxdNHc+rptWb1SFXUdpv
qMg21CBKARH6bhfUe/46CRkiIvLvbk5y0bv5gr5h9IKv4Omwn7lh2yA61EKCl4rb
3VZopBnHEHdqt2uYyG7PQWEsH8/+YfxH3WNoNa/Oj4g/b/Ydmgx53WngDKbEHOBy
PBmp77A+fHlPLT6nJKbWSxJus9FT58lkcScMBfaGrttfV3ykzNcfAI3Pn7856OFV
1+H6tWLfrqQKUFoQuwcfiCyZsycSdP204DNH+GkU1bKh9sx7oMWlanS+D6TyRLSe
+jpVA0jeREhZFzklb+JhjwR+tSE2WakIyYiwokPQ2uoB2Mz9i8Fx1n8u9CgIut0c
JiW1ck3fYEbDiz+Qk0+K5srNbH34wBTmczgI/qjAyAp+pqoQvyInhIwJjzDOGeU/
LsEQ3OnAEbuRSf36/yo376jumhjsUG4Pdy6qJR6GCBs6pt8iUdBcZNoUMYGq+B1f
GOXEvWYNCesR4U6c/4h3fSvhLq+5FUXpjZTvxhEwlYBeG08C9bzvDKu+UWZliLVd
TvoeLhbrs2ClwnY1qSG40BRvfGg1DVhQziLgXHzQ7PQZM/rtMlxalypI0PnJMASv
tIAmT0WSv9/vTbN5bKwGj+6j2i7DtrFa5kJ7bhzrQP6YkIfEpy6QrlXf89Rof2+I
aX3S/+EV5TfwSxyOc8WJ7NvYgaU7nX+/c0XlSofqW8X5qjgct2nm2mTrvvqaRBr1
kywZdF09afh35KL0min9URRbS6RvpqioT/22XjoSv6dWZJry3aMHFTiHJylh1e4N
zS6wDY3w75ALeXbAaYhk7o291vXrssfgcQ/Tr537b1RYtQuhxhcoDxQwvGvCanl1
mv0HBVJxs9mvGSIk8TOVzsw5P/2ONIUaSh0TQZS0wXQFLDPOrKrYDX/vM1o+NmbA
ZV7B8A87a0Ute0SLNZtTiss111gM2yiJq/K2NtNtg8L4rkF8tN0ZllvQTcIoH7kL
CFcC9wEOSYTIRI60CBXEl237XIb39RyEf+sbqrYReEDwC1DYA6aP/ivmXU2e4I/I
ek5VZ9pB02LwgPQ5JaUdSKf+O3fGXFB6caWQQx/fTN/gkQDUWynMcXoocezcUF0I
+CRTtuUFl/xlWgysUfrCg+tn2ISJQsErU3IxkpNSuSgAGouYxq2VPz4r3prb8y9r
fYQ9gDX8aVBqFle3auMGtZ+XlULLHHluPIGyTVmK3wGdxvWqKzP+7M5I6LB1hYhI
2UrB5oLEhfBfLFh5Aavd2OY/4Fykjx+z21y+/kQsUDvjH06YmF2u5R9r/YoMIYKW
tLcJgPvE4vj3VB7X9L7lZsu4Y/gi+VD8KvUUwwoTiOnO6BcVlzcBctEUYGvQZwxl
0AjRJ6BqJs3VZO76VkCf6e+OAcq5nHwqWMVlqcPWd2dysIAB3klmyl/kerwfb2QO
8fNcn0WHZthgrVVMB6s5og/wxRuFN/LvsDk48NAp23HRRBJykv8C5l+a2fei4roJ
MoF7yZxRukBc8izZu0XtCLbAjsyd527+XjesBZ2b3AxNBlTCuGSjFm1IPanY8rU3
wG6BHfTsAvVtA8XlCfbhdn1O+NLaBbrVtY6S9cME1W6HjtW+GjZGEYfxBJFTrpWg
RxIcynVCMH3qoOw42VOYoNqXOazWDye/v2rBAYZyHCZ4HD3qWQBx5wGg1Vmlv1c9
zk5zEaAiqeGXv3LEWfcRy1ghZmTzf1FenLPmvQ5LfS4NO4SPIJ/6TPgOkHsOy6as
4vF+apVGNszmrkPSH6qkrP9K/YxhIqvOeFWboBc60IdFCrWFQMgOg3a+eUFDLzhh
hkBM7O5+ttxbp3hFm4HLdrZivVURBN4/38ZhSq/trlHn3dFhbPmaIErvfy3zL4z4
u3olF53rnPHTYK+BeFYF4OcFIS0uq4oj3zoX4FWs8+lKp7MI7itrRenAHHjfpK7i
l2yNqRZZpAPV9qeuii7Z18kF/pbXvoLgBT2lG6IJ1Ch+ogt1+m33Wr+02KWc3dW7
l+hMiwSPXGL8NlPR2a9vOWleldpms3aSaZLCaggOjm0Mpj/qJ3ZMexY17MKm1Woa
W1pm7FbDM9Rrx5cZLgVzKtrmawx4VdYn8DVeAbhGIpl7IVzVEPtRhpdTkmUC0iIE
SrDnJ/4nPdj4Uvogd0fFk+oldWPhs1KieqrGZpbd4GfLGWw3lRwGkPixGDlmEhPc
q3nM59JNph82Yp5DAEAOZNkh+teu/jcfVcbvZUBobg9Y7CStvpqFJ1V4SPftTuzn
pN+ShvJmSCjLotngmfQ0qDD9iTT6Ckuz5mvPQXELkWcNwAIVTqvt+gmUW8iiwrcN
86QSObPX3p6+SJSGmLUYfwtrqVMbF0zAUkyD8URdJN9CLqkiiNIlL/YkIHa9nEUR
A0JACX9h01JG71VKhhcOLRQ652A/stnFVkq9hOlmEin8Oz1VWYY5SUIgdyFBM1Su
fD27BpryFJS/jLf2jSweUTlxWPt8vDydsAn2vv21Sd7w/REKi1Fp5yiL02jP2UGw
Xh0O0RwfXd5YN1GSGrzQ9A0uIV2/O+JpfrlgRY5a6mOHHQtk9fkQMQXphiOoUcPs
j2atUAumyUpepTOH9nSeK67V90ZeD1dvaSDF20/R7Gg/pnnM43zctQundVfNJZpf
tUSaM2ee7tnFUE5r2T5hAvTG4/9YemMjRKTsfBXnfFXxXnlw1096mCfEjLT8+ff0
j5veIMrs0QZiftm7sp/XqPvm0LVVWasa9B8VvxdTHQ8awNxe5FrwQnNiIPo8nLEa
dE27rBdQ3ysu9sgWqDv6ytICOEljhj3uhuK+sY27org4lEkZcdSQmONoMc19irYx
mUtUPieu4OF5YHTSSBDR8oWYifmQW09N6n9GaMyQxxY6F6o9EcjwMFoxdYYWtAr0
TElhvY19Bx3XM0m8OVwDYTNd+HUDeCQHaDM4ZLTgpSNuvO1iPTlPVVagpk4MyuSm
Utta0nH2v63nJgnL1Eej8SshVf7f0cgyqSjlfnXMaryWHeFS5gRK7GzhGSKLR8Fp
FFrwRhKzzaLkHaClT86MgCWTn3yhF0LKK7HWYI11skXk2jgTY8AjYs23W7MZuofl
FwDB2OP28UdDzQaPMVKQ2+CMNBPkk/MThaahR5N6JTjZhavEnb9wemlmY9/ELVUg
Wz76erUi1dvQbCK3Jl7gh2JYrdKouqsI45f7HxuyRngNPvKwdao1tj/Rrluk4Nob
kyajxI0+elMJQcZfczjStpcWt10qa9PuCN7uxomdrQQxFgFKc4bphXBHAoz74Pvv
86CozjieFRHsAYRk+M74+zFPJm3Bc/uudc0IfYv8DcUWyJLIw/fiL9DhGZFeh1EU
hD1VsWOh+yfTu4hS8KmD0Amohu1Wqk0rw0GQPM1yM43HgujuV/xzAV+pT4CXILIq
FNac+OVm+eYby+wgrPWrTw8g5YTumrFGrKFpK1EF3utwklfj5y74WRbnQ/HYjMdo
IzR3HRGJ3rLwfrVvLpZjLZbHARCFnGVWvcBLZ+ySVRt3twlrIuB5l59obUY00Y0V
5dkE3T0+o35/tWig2R6KEpui76VCRkuIcY46PJAxnNAqvWoDcYVoj/wbRw5D+CGH
xmiEsll0I+dA0/xECJGKH7sJ8yRI7AddKD6r2pft5wMhriUNuVv3A1wf9sFkrVvd
6Ry8k7sKkzqzfJialGM3spnUaElOHl4E0kav2K/RJdb70vUROIoKjJ6DVH08eR5S
I1pAfpbIsCgdyT8cCJAIT0TWhP7kkdlo6DdDJYCaOEqGN0DCfgAR+++H55qBWL1u
vbFOLWzFNeNgm+1mQDzouK+31JliMvoYnJ3fJdX/AdwIXZdGofl1Gm3ma/UAQBPa
PImfbJjKvzkVGaDFPEexM8beK+hlMcmXD3eCC3KWRqfN87+2bPHkwLSyEVdoKjMA
edSZ4pp/uP3MFnyDX+UaBxhreJjrPhFQdgT44VKlARSUOI54eLG4z1dyWTc8VtTB
bHMl9nQtkpDLWYZyFZ/PoWKW4PGkFE3UjzVLS2OLqa1P2aQxW/mOZWmhEcdpMnL9
MrTuVi1p2zMLlc29p1dZRhldbLtZFESk3QKP2kPtD+qhskJKq/+w0s0ZyquuXGtl
xSczPLAWZBHBOlAJRbyHTL/pQRpdRh2dAZH5S4FUghyBp3XpnVTsRA3iVXo/saD7
cwRQRROVICdeISI/lyLjJKQqDMielqjp3grrB2IF2pT2BSI9xNzr9Jj5es/1vksJ
ORepFzVjnPYSneiPvB/NGhtuwSA5UJ1WpZ6OxWFEGCGRhgBG07f1I9ggkyViePij
FdppzwseXYtljMRDubEf/d8k4yckVmeBq5ftH4rRkMM+r/yiw6e5BlbPBFZJjFeH
vUf420p+qUm/aIC/hGstYB6p1Om/4T2uNyN+CJ2BCAM4CliTmau0ucWmpZxmdQNV
dxLnEjgCdDt+crCKY6Pqukh6anr86W/0ELUWcrLPDvxW8uw+/QbGau0hM3st4is6
XxkmHDNNnKQEQHppEjgzwLxx9KKuoBpxbzaNZYxVzH4IaC5YbMbeKqUNGmQVFDvN
IwNLNC2zwPKj97IouJ47hlVaHa9ZW2YsCGeZ2xbb+RSQGDT0c2WhYi6hlKyfvd+8
QBKf5AHY8m4qGc4+SjSK/jlrVInczSusKHFTJu/DKdJ8cw9I1cISWiDkkUssRZcU
El+BKemhtL6tz4LIoOJSrM5KCJ+PROCOPf4P5AVRX1smlfEa7MZ8r4L/LWfaK6T0
Vu67ibb+2a9o/Kzdg+1LGPT/hJBp2whJYg1yJWp8SDJttbkxo3X+J2zJZOaoFsSo
K5m7DOXS2P9KydmPI0Bi8G//u9Qcq22ODdNGGEeEXHQQpibQQD/RcrIsD+YD6KcL
MYecLhW2Fbe9oji5x3rMTMgsHVELvJSB7CCy4tyfk4g3zZPQaBf5hrA1c+w0psQH
GbS6zKxtDsiDwMIOxyiyKo+IRdaldXBYvy5n3jjafC88Tqdv7jiUuGlZ42/UftJF
6xc/f1IUWQpK2zFLic0G+licnpJpYc5g9JAPFgUlPhrA6j2BLSHqPcskVRFfetLp
3rimm0999iuNwNPOiSk74M13Ncb9jslYJqh/RhWiFNkMKkywPIdAwXkc2rvKomG3
afFKPTWmOOINyiD2OFMQjkU3oXf5ePskoUr4mk7O742k7vx0jbbJI9M91p6Aq3Vz
kVERnvzhu7aFU+4pegGmyB50uNULf1YaFnNpJEti28npx0afB51guBHAgDmLBXnU
/BZ9LAiz9i3QsoNDs+UJPBRPR1JsLlcCQS+0E5FOj4rlGDsnKRGaeoNBswlhNjmO
DUfdpQ3RJ877ijlXg8EHOHCKeFhmtekObL6Rx2CX6JPg+cHB/hyufsjH7eheyRxv
Hc3aPE7bO9rgBGE35O/jkxA5kWVNNASM+BWvthxGRRqdVvNNb1mmk43ggxpL+yDu
TCCoLf06FAJKS8BH6HYAQdiczl3zvgU51RVVUvn46+gDVE9PcSpivhuofak1k9Yy
Cp8yEiA7anFVyPOB8KqAFDWaEzrBJlksLWqagUi3BxXShzQXcul3ERMd109HCtZa
pqrx4r7LF4jn/qmnFkChYKY5jgFQOa/0SVXQUXRR59A3FRdNoZbQhTspD6G+8ykj
jV7QKOoAIXtl5cZEez2lHEOALG+U5TlHv2kPK8RqDppCvtK64MnLswXUCLqgPTx3
jQSvJcqkyY0bZujg4TY92NKZQtNfwqQE3AB5EDPCdpQ0LYrETIreftEdBrsXypH9
7jywM1usW2/Nw5FT1mbBrHq6oSd+1mgvm+/KsfcK3x0jpITBnCtbir10KYdx9nOB
eeddujkSjvEuPLE41DjpggOazWBdVbK4jIAlajolEnZMSJtA08EbuRcQU/GGc1Nf
Ef1lv1Rr3Y7s7ZNVM0zn30CJitUnUdFYRkjE33m7i+UlI4GT8AbNCmL0CijQBTpW
jAglx7nQMLBhuMe3RYnWfvAb9nM30BI2qdAoEiEUiUouKqftUXMelsp84ele/n5E
SByvidhNxcgTRnpbkB15rZ0meTemQIXwtYiknFuvMmdh5dUg3/Q+3Ifv1UxcgdNH
jQqLSrj3QX3f+pwM9mnGmRMg+w64ACO7pvb+aGt6TjCYITu/z4KB0NG9mg4YKMCD
3igl46DIO7GhnClhRCXFKi9Moez/pZgsqsCeD7i5gFU1sQOAn4BNxgzWvgm1sH9V
EBpVK58+jnT2DWZhTipFGbsELXijTbW26iJBRpwb4ZI742UOmbWvlA9u4/YoXaeO
Z3Z6JoEhr9QD4oop4amfd4YUGfnEv39tLHrbAqIjNWMsLetTrExlYRpo76zfQ+lS
NAUvzS7HOAJa2aGBmQkaV6aAQc6+/dSPO4iJzHuHl3eUljuTIG93d8akGsH0V+RO
FPVPxn4lTRaQjvbS1DaiZhDR6FZTnxPiWZkMHxRH3Q9BFQeKFQpGU4HG6P9mI5b/
69xTNw2pcGczifOCupA7kbKgOJULoffhLKPJ00BIXZsvfoJwT359kPgCOaR0Aw2q
dM/kO3R/Ia6cYK4dYP+dRHLiVgKJWPj2tYIUCTNFEjHzF9qjsJ3iZEMpa7okjqy7
Cn2tUk30HR4Npp4VSCXWc+dsN17s75xINX8ZlpkmQXoKYjxg1fQrqlKHEGHcfHHG
LbMK67Qn2zKzckhupxvVBlgHE7rLzdbyt/EPcsGe/DK38KI7wRdYTO4bfjxI4jz2
Uyc0nG818ab1j50/RelCAe3x+hNmI11ovxJFbQEh7hSPLWjitYKqgqStZcTFdUak
Ak2+/NnHaTxORix9W+7X9bNCrprbNecRFXVx97a4fXjcCw9DKx7gtbo63TniTqVw
31R+t5q0u2XSvaxfQ/6pEtS49Pkt1hPUiRI/GYJvHZngYuPLheBgT8JSFz+yuuyd
pw6zkDdQHlq2qYounDVJtfgvjNkheOhcerLUxurk6aqPaWXcjuhP2eS1T0OljHls
tzlL/uyGmuoIW+LBmMz0WnMo89vyZ1Yp9JrPUav9AvM4xFiv4kZXt51bThY7WWsc
rqTixXAw2vBVSaJeZ3UsRFdHlZM1mJejwL94TIMtYgEHbnwMVgiWNQOKky6aXjEM
NfpZoRaiLY3pbV7eZogURmHjcdVweIzlkjSEkVdcRAlqLCWCqQQtHrR/1bYMJ0us
MsMI1AimaD+E1i6CrYFn+mx/knnotKiceE7jQ/hozsdFUZktDNICW4Hne9sQqjKt
p/Gf9X89CViinh8FYR2gIITwxxdyriEafoO1OScDKdTx5w5MGF2Jn7sJl7uQMe7b
Ts4QeheANB+cl5SvCxDxs+TXm5r6Xm2JNEOPpFIqqzXPxZyC1B8qonqYlL1PWTOb
6avaCetlTv4r57OEJmye+0lxHduT6mS7CWKdjkQ5Hy6aYVBfY+m2yazWP0IWaKvL
/BhdGsCAvr7wa0XaF97GBQ6mVGzsLjUr52/sv2c2ONrxnH+EQFJGMeYgdTqzmBAF
QWTZH35mrnZxALZtrxH4+GFJFgOOmc8tOBXND1lYH99/uwKc7Ru2KHlXgaIrLtOo
Z8JaRIsXj75QY6osyF9ybuc7Le8QYHuAPIKYiWoRpZKw571A3SY1iLYhkwD4agEW
CPwBqQ6wX18CCep7VhXnagVGYsJR0Z9Po9o2J+vtKur9D0dTz3nmyhTisiv/g79Z
R8QHpAJrkK1eo13CNp88dq68lXXGK8kuQdRYtKEzCsDkMEeCcWw5CUxAaU6UB1n7
/rt3N5QYEoOZYoDJtPfF6wE/gf/V0EU1AHkbSGF0LtLnO8DLArmAbW8y1iFVCQDP
ZdUgOzf+X0InxSJWMX0VqhlrFuT7jN3sySatPgHQK5SdKGC+0tseuWlvOgB24iRe
OHALrfKMkuyC951VmXVOv0w3aRRR5rL4qydpwWuK+xCX9rK6kjSoZNpNU83cUMHx
nTUJOKP6TasZohaHIkxJ004MGj+OTTWgGPnVbvL5Vv4BrfRzdjLVYDzGfdq4nBnw
JlVxBtKZBa/UsycS9AE4K3Nx7JWn3fboVItzznTY9scNyCJwjV7V3/eSjP3E4aZn
9WOAyOa4glri2xK0wDYzyKk74/Iouw+5tr8mSoj0wxYiENFz0ZKZl8LEaDF4zCO/
I0lDIwPoaotCHt0Mp3EIAxr1MPSZNf01F/qsxy8KEGISFo63IwP8JfF05QLxwwC1
6obhB4GHgiN1UJJf13MMBmm0bI88dPYy2w+cYnPjaLW2pcGHFjSGdBgdqxUCWcsS
NJsR6xua90e16CBUL7RiMPWUzc2Ev4HWbjs5PFxfO1Rf3e8dcyxctMiGoyJ8hUlM
eCtu0xC7BO0EnLIzZeenbsEnsB3JCkFhCUOzBQ0svHVin3jU05CShXsU115JtzfV
PgZ2NECj2KQjsQsU7ZuWxyMUwpUpSSYqKqzjPGjy/ZKpgFiG1lWgLjg+akbzEBAu
mN66+sUuScQf04VlegCM6jHYrKWCrxowPIQN5pyiH3x5/Q9BM0AZkQIR/p7whFGc
Rs5bwe6dkPN5xoGA/tS3js/XAklA9t5g9q4hs4TOVobBN1hfdml49ktE0DxbpD+F
RWzcO4lby4/hrqXJuqYhfr+OIti5tqEhIsxTcHRCwQB++AwfO5tWv/pMlPYdt6P5
Y+cUK3ZGtR5e2RcsYWICOx4YIYg4uVFueoSnSBWhDvColycoab1A2byS9TPUL+8o
3V05fl5fpDJAHSygukTAYerJbFgNprdda+TdpXMgeWcs1lMy7EH7LdB9d7jfCeLV
PZ/mnvKBoPAt6321yFTlon13o+GpRYc93JrWn2XCSrRGe7eyTRrCA9SCFRw4CHFr
jNLv3/lirDfPMzpVupA1IbDj7KnjAfPknjn92EOEM8vxnOSVf73h6QN31Sai1tqr
Pxyl+XFpx4Sygxd1CD0rQ3L5NHW1hvj8trPsjTmfFv1FaNqW8SgR5I91ntnnbaEB
TavgvONNIfDga8gIat/TDzq5Q/wyeoZzPm0WwjEO/uhV3erOygb41LYOqL/2nFgh
JlhvC/0mfHYrhWGWATPAAGsTekfm4Nele2uvupFP2Xh8GXPHIcj1EywDHAEkgnOQ
gdj7FZBOc9kT4rQ2iltLLnf07ApGLHA5H2PUnkxeV8WPXsc+Zi8FRm1m3zsb24Np
eNPbQjNVZFMNbBj7ouNL9UejmEL0BccQaKH8CAeHwbcJ0LXd2hczgBDAc1UFxbrj
tn70ef2kP7vuo3Wdqezdyip1H9EoZOFJo5pcUDjfUPAsucQ33MtOZ2OgIM57qIM4
lJ9/z8ic94CYD2Dcd4dmIJdhmnVsyW183E5LvIP19SVVk6GHB/rRZEOlW0ahFQzT
57Cx12X7nrRTgiroOP1jvilTiezS58iYXE5kceo4OcSHAwZfU5xTFZ+6xyRyS2Sg
pM4Ss3EGzOgx69oSHqoBo8qaqPUm78Qk2tfK6qXJbV4h55zvSQf+CdDUmv0gnOcc
T5sQG6R4o7X3262K3QbWmspCtRuqpIDkNYN8mpRXkN7OYlo5GxIOcJ8sZ2nUmk6J
smEhGAHiJBMGuNLxUfFMPOo6OtgV+EKEudLx+g7RzjZYknbYsHaEqyrC0IxM50SQ
PazQodHS++r4+Lx06Nlx6yxJ/yZzMlWse9w4BTLKPvs2p3DspDgfrHNXGRsUt1av
bB7JZc8Lw8Mp0XNC/KRHJ+DilJXYgzrnvwA/tQSHLfh570M+2FI+klft5HVA9xNY
IgCRLgNc1iL6YnPSk/GDdgyOyKfI3VzSVVY/jeVCaD3hIz5XEtt3a/MGMC98+hbN
FGjOdPzNjU7znRqrJU9eHWdnm8qdmA9FunP9ghqdz0MRTcX/Xcm9Oq6tH2JvprY1
I9N2QvGW/MgW/N55PRHH21QNgOSXQDtPwYvFDYRA0ZwS7hGW1aaTC4vC9wZz8dpP
R+D/6jAlbsKkT9j/WSUH4Mc6BVklimnyw2lTO16FheJIIXKefxYG5V9pO5gZhHH1
k+ac9Em4wjGelsf+IHiWcNFqg5xYqIivwaAwjdcjRbFZkjSQmdv+b+LxpWBSI0Sj
g8uJNhc28B3w1SZu+dgVqB8xm//Y055Tg3yhP+2ef2ai9igG8v4FuMo3WFyfXacV
RWcW9nE1QIeuGeGf/9casyR08DZQhbFabZ+av/sLADOBGtwvPAeTWJ/9DpyfJx/m
sMYmmvFiQLz79tNJEBdmD4JpM527rEGiQWP5Z1NeOk/6+02P4BS9EBVgKcvDorZL
wfN2dALK45zpgayynpAM87ug8Qdw573rlNMHxbm2LvB5i09tyNLiqgaDKSWk7l5j
V9MdgTm0yP7ATcF/24ARXgFY77eeUhhyKY6/nxT/Q+NKEpYdCEFtzi4uQ7KjAbKk
Ua4kPCMmHGtn5XBzQDfiTMfmOG8AKnEi3jVXElBrrw8+umi0NOsfxZqlw5Drzyub
dfSAnUuh1NBYtCE7yyCF5Z53xzTjig8Oack8BAqMrIlTBQOSU463j6kelSYnBIq2
iWRwLG2STAyZRXkXcuFyifN7hIfpCsUFoV/DukE/6qvfEwHPMuvDUWsK7j4Ulfg9
zJIrbcevjLwrGUXOLzMkVUj/vg8WPvaEzBSG84EG+XC7qa6r750SX+tmfCxPYu0u
MvjhX3iIfff3h/vf4UUenqHOewzMfqyniefuzY+qd2l4KMLQ1ajFMN1pcc4ZjnFt
Cq+9CqDiMU5A9iX/HUMq6j3hXOHcnFJY8JDWe9YJYbugc6658tEByXisiuzv7LxG
IlRiieC+uwZMYwxmEsVt91704k3bEHZWFYJt7UxraCHCzOHu5yAWiIzgTMKC8S0V
sYRu7wDnkkr5ECir7iYGF7qDrAbjTMWOumcNhmgyskR+BR69eZX4Hev3HKQrpjcl
HstshhAYs6iVzJgFosgN6nHwUawEh5xRTJidSDYUxcqtVBKgjoRckmQsfsaCUegq
RHzJJ3MtdIMA2DIUZV4HfE+bDbAA4AMdz3gqk4fri0H8syPerrazbCEBmacqDgiM
NnPA583LZpM0cEO8pOASRoDPycKBpdr8bGZFme+twRZEfKI0p6V1VEhFSE2j24tn
0W/kejqmR/IfvMBqF6Elb0kSY7/kB7z8CXTsaZrVaolxCPDS7sphMZS7N6xHyoKn
3zrlXb8G0zfsTtyeqCn1TbjNJobUIL4tKjrZuM2k1G35fGOfGeOXXNC01aucTKby
q0Q0a+5q6qIrIemiOwT9m7qpzkpr0f9gnfOcK7nrNQQ7WPtYACQJ4kMYqnWY2zea
9CFrSyIVJgbGjxKeu7BF6gQSwORSeLzZVpgxoC4TwwfLM8IkGwQ3GejEx2RRy8dG
p8opfg+aHg93IifAZdjhmQP4wm7FzVmzIQNDyXhjUH13saS/8nUN3UCmauvrzygo
NuGygf3nloEtouc69QQeJhUj01lV6PxEnpsR9U8xMXDwRP6XQmav2U9idxbCmBj2
d72V/uD74qQjU/pywLg3L1OFZDcO5b892S0EUjhMnRNPlk4AayrZTTBp+ZQ1ZAWw
CWhsg9scZ2UL6ySWmVVhAwQ0yju+FlOgrAlV2OD5zXvaPJ7mENhxG/aUB89smUwo
3g6zqSTA7frz5F7S7iHSlXRrA7lcix+jyhs9qBwsM1EmRb/Q8pmByGAQSSI5KcFv
HZGcXONOiWA2j1048Jk/YjmPpHJo34SENe9fXHr6bCnpkPtS+tdiYwkCvSrr3y5q
Dt9y0DrqQ8gdKIGZGZ8AxxnREVzYwg002iEd7M4vEKUwd4sDuCRd1NsaWkH5zZE1
jOoGZDiSuHpqN6ShDrbqp7Ne1a/FRmD31iHASoASe5XRQnW1jjSM2ubUcmUU3ISj
XMg71bekwOPcsezCWjWRlxTNdnV+8hRcKWj0MrRKEcj1Z6f/rbaPLGpsNXWSwxJp
9ErQQlKHFzUtk5x8PrpuJLXcUzuYbfue+Y0rb0JqStSgpNJMTXzYrcbU00rSRynM
oQqK4whksl8m7A6rPGb2Foaxq1yMo3uPXU0WlQ38HJXQyKKMMySNFZ6l/no0WT4l
RfrCKFIS7dZQGiTvsloGDPvSnWzupWPu9zxjFxTJRYF8V2aTAeRtVIagkYfmstx4
3vJGqesxsYCunCRjrxRiC0gkJmbPlJsXocGLVcaEfV4uPoMgX/IyKetzSpHgnE/6
1lBNjXUadZdIAUopkfye1ayv4+BNJ7yEQcz1pBZ7MhAZALW91/5QL41zq3Thzvrh
xyUnSxngZOF2Icgm1KBPfUq7QJHKArdDCbWvoU9YFWZaGzx4UbX2rnfG2hMC4rQj
dObxU8O6l3ZAMhzjhNFHBBMUxFh+/rY2pn+49Qpi7e/pj/7IaDw6HIAt2Ua8KA00
4Ti3IAyE5LgD8lfFl9AkU85pHYARqKIcQGocFYQqt+d5jvUXvcf7WBfJl0DHmezg
13X1Ii1tkswNW6F0qxQNedWFmB0O05qH2WiFXKa4JcVO8sFqd71QdEdfQCjkN5HO
DqCtXIRAibylgIEv5G2K8yYoaCU6W1wHDS71P6EdnvfUwE2KZuXO+vmeg+oIzGev
t/An2pwF7EM0KRh/rHB/joipodQQRkrpdMsiDO40mjms6W8bFdSbRc/ftMcp/Xhn
2vKL/2P78TZnlc7Ty+PFOyXprs6iOcVGpNY2Qmtw5i7ZCQSzTTUnhalZpbinelea
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UToQoyi+a+SREAKDmGafqW8vC+cdH3YzGeO541dsB+5Nn4DpuV1BDZoiv4g7aKVY
dAmizuerzG98Om4krxIyduqcikgYO7cv1tXmWqAKRZy5l5myuWllL9nQAvhATnJO
V3KTfxY3owCAOkbBIvOCsR2q+rxG8lCY9nQ1P/x1Qv+U0Jq+QNUza6mQN/7zTdwH
LrA6ryvSHtQFdktbJgQ5g/wIeSb0FwNH2B4JZ5wFYklHCepbMmRoP7nP9LMtBSoY
CJFtXOvJzi2o12u3HBsEla5hfeKSlZ9qzUDPhsFs/nYJecVev2c9iRYCfTtYqxaj
e/n3kXtXMpawa2L6HVfMcw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17376 )
`pragma protect data_block
VGv+sjLDioRk6Q3PciWvM5xPkNv0VUyzYo7p7gVDgu/zktlb5sB76HtRjDsrVuJP
SAzbRBNjWbzTyiG0flM+97U08Yi9w7V9EMLG1hHyBv/EGqyicidEwAvYiS/5PyEg
x6dbmvb5633nU+K61IczvIZnEywNuZoqZPa2D6DrxST3npD1gCZg7YrPn+Lq1fdZ
edrkBmE11VEaibjjEx+SYaJpyq/pO4nGGbrkdUAjPdt5AnsYv29xCER01eXSrfUj
ElbW4N6+SOQ/JCleMLye2Vo5FX1SDxYb7xLS2Z/gkT7ywHL2ZewQ6Z9a2+XDfj1D
idzzV/qLVWvoXtsg/7rm9r3rdhtDrzlbgrWXkyJvan7mveeJsSugxDzHg9Bt1QPg
g/zM3MO4xL6ksJpRwAyGpn+XFHKR9qEb9eIeKMHOPhRuY5wRj8T8WShMaYJNJudB
8ThqlTIdcor1S2FMlk58KEqhnPtBl+2GUWAhaOcXZSxUZoY269Z9lM5FA5okHLHs
BzS5NghBB6580gPGCIFWPB1bFo29P8D/5ZY9t5Xq/EgSSolQHPTYg073Qn/Lv0Iw
PZXAVxSJx5qacx4GAD7/rLkNyaazcU0RTiGQHYG+kUmp3hPVBJMDPc6PGLt5EDIW
/VtGqYIFUhI25qochAXi0/9mCDf7bKsO5MRuc/9UK+6ulN/R0VRlvea8e7B8OZXU
ybvCrWu0cqHhTIJu2z+Qs1ho0lb+VbFwC7WjEhuuNBPdpMBIOfuESMGORmEuOI/5
iS6jbtIK7Af5U0YE+Y86mMFqvhtPEunKe/N/ZJdcfamvl6rcLyZQ+NLn1Qg6TlaG
//GEWy8E+yfNyRb+xfDQxjzlORKd69+QoyNHNensyW4QFd8gdJCfidjKSVIuRvSK
W4VoVl0Hvtxlp4bCtRzbkFEahiMsIIlPJQxgDqXfeAVtAAvHeEsXeXwI8Luqu137
5sQZjdbVvFEhFiNPlc9Il6RV0wYvepyTN78JdGxdSTclcRJbZ/R+QA0NjVNQjmWp
DKDJtAb/1UuV5+Jsdpk/mGBJT2g7YMogX+0OXBpBROrU/S8GcDEOPJm4vTA5vyc6
wGf6iDBPksOE7PPQBANlrQqM7NbQGvQUwjWds6olw9ffNuRJMEH0WE6lDtCOjEnf
E1AQaMiFDH/4VkYY92gDWyHluuJ7BAfq7JFi7XC4UQqyqDFFF8JCKJoCRFdT2Sub
eYHvLVY9ClP/YFz65tqwckiabuR9xSn7rtsD5qY8Xk5DHjsoG5YWBNpY+A7K7YTN
l6gk2IflwtkNBUUC4WD+aNiUrnY1fbRxQzBIWf40y7f9o+xKUk7OGiGIr6QYAYj9
wMNsgHUdIO2NB4hhWKXLbHY5GVFPHSIy0Xz53KlII69Ib0Vzk/x5phOItw+4VROG
4+R6+xuzIchgtjbaFm47sqdGotAh9zUAd51ar9Et5n3hOOrLL3qky89Iy0o0mjuZ
E0RR9+b1/h3DCuqlQJT7N+oVvyEy8gHp/p6QgVfQdCbVrAcRkd7TrcRAJLDlQysQ
rFV3t6eaUq6wa9XIUIDILb62WSPd9qjW3gPcbHl8Uzsx3abC0QEMVqGPYqppKh7/
dRLgWU1I6WooImksaVdgYYPGC51o2vWxvk39l5Bw9wM/i2Ek5tL92pnjISZHm4Hs
Yz5gUHMLa1Ncs++XBdMmzQVP/2sxTW5MBYVcgUTG1T7ndBI20StGcdRyftkPgrNU
om6UaZ5H6oAGsurKQGZfQuzBcFwGC42a8t9zokMWJM2/1vVVef0AQHNr1G9IpYBV
uWX6KH2zN+wbdPu7mQ+0ANuy/CKVmh3nJF4A5lFQioHkQZ5r992n5Svg0DnzgAYW
2mMbz8BULqZfGdgpnsD9f8cZ9Sb+drGoexemIvfe0Qd3dzra+L7aMD9G4pNs9RYd
LNhsF8AyFw5x5reequwks+KZJ1QoCYj7NLQvmfE3nPiCySHWBXiDjH+lAorDZw6j
kbpjmotLVKErF4S81skrXxDJMwSxFcWIq2cNhnHujYjIoRX4FZW5gfm+IcZAOy7Z
LxwMSD2B+8cy5iJ5FDRLnopYXkwcNQJJ4M5pvldie0yZBZQUQSeOKp4rb+AHxns5
QIZzIbuzwRsvw9yk2hql26/YNQHWjAJZ9OBRLMnFI3Bg7oA/OFE5Mbb8WS+0GeSM
Wl9az3aRbh43Tgt1S1Lkk7g/cYrZbc4xjIS4krgtcs0JufETbTxfL1G6lb4VEDVk
BkXhK/qn+QInvblUhaa0WFQd+yUTdWMMHRbNfYVQ3Kya79b8esfMG13wN/uGtb1N
8dNVhmlfn8GoeTYYgIV+RD576wBo4zbOk1ML6RHuK9AdQghzOztJuKOwF/DzAKf2
yOL8f2G6/MbfvUEGzWuitAqdg4nn9xriEWNG7moD0WcCnnjIZ+qKnl3DI0JCavFc
UYlEe7OJJdkCSD458mlGnVGKTieTE4iEmOvmMmh9SPFhs6wF02tM7Frpz5SXeluH
AWpQRTRXc7CKKf85/tLVYBPNQOnEcABcD2WfRP935xbk18O8kb7QX0CA7DikMneG
Z5HPKCRpWgLK90LJ8Fo0uKfzO6TYXeB43Eomt1ZEsGz1lulg8/tyf4KIL0ddiy1Z
yY5cWk5V2ecF1TI/WrUlWmmzxCygl/9LgiyJG2EjY7zUposu0llWYYQZhKenYigM
ru0s6WJfClYHf7RtsAbfUlgq2pjRsJ+cQCCZ88bdwc36v1/QUlQ+pRKtfu3SNs+9
tEfAWdNvdkHBVJ/yXS6wEqbOQ+97Icc7Up3KDkommaRg3oiWS/iftaddsob7//iL
lH+s1sD4S7cQEjUJBg8a+S27pjXZiLzqh6d2tCTbJuJ/AEm+jBJIX3fK96JvE0pv
TvoSoHqv9JBSwE59/UX9/68NJJliUpkBVZpXjHO3FtUgJAcNfodvHsyhN+JFQ7LV
kxVM4nzWGuZSwPT1ycDGYH68DzWTsxY89VOTn4c4q+4V6Ad3KZ5mujxHwQnGQa63
iawpXVOEep/dORkTBvjgDKFJpTLqdog/m7gAh8cvuIN9nCETKOm3rfODa3v4H+Xj
IO701j2PgRLW7yShusmbPsDplbIFmUrPiBlGC0YXDGLxQ+oaAaSkKybIRZniUvk8
yU2vFXFjx9K+U8kvQwEAocoIbQbW+/PlvhObWeRSupqSk/EMUFXHXRGOXMrs5X0q
ZBFQ53Tzw/knmibiyRrmGvP0H41F0yoV+3PZojAAj1znwgZ3saHsGvBzTidE12fK
FPoHEnDUg6HQ560WNm7ns5OclL/RzZK5YPP1Ob/PIYR7dZDy9W/t1U9QNZlhSWTP
W67ZmhQfQa0k4EICmaGeGcZDpA8Wt1ST0l+ToMY5KorWKNLplaMgpYtMxwv16d84
KGWBPwLIPhCONve0vYChsvrDqL+5A+VKAljQyz4aX9Yvr0yEp+aPL4/J2w7sDAyz
eGud9eo2gG2EftLKjWU0cORpuL+OdlMrt0uebxzMfkc5Wyso5fBn3g5lOXawy783
D9YBPMCMM5dawoVHnf9lUYbl9061/ySNt3sCQar8cmC5gxu17UatNKDFhZuAD00u
u/kizQ9qzO3ShJhgvKse8F4zXkYRDqCEvxAzXq1IYma+knGAjKJHHAf4ToJHoDZF
DR57J/VxiHzyn0gyLD8c204qi51A2wF50zcScr2aPaJjrr22XBLuzEslA6ZLVp+A
SF4f/S+9HAOgd7dqQftjILa4bX4REBOJlqnuhccDv6A3+ShZqGCLwYh/RNIouC90
Kvl6uBzbQOQwZ+NGHoMt9oL36iCSYa+AdqFBVwV5ApiE6ZkoWErV7XI7EObPHTdf
6rIrdNd4uoT85enK1Dw05rc8MG/yhamJJLX8SjxqkelUoRhGEK//Wj46Dhge6jmD
atvtm3xu+EuxW1y55U47uUQkVyQsnBWZJJgVPiNpxR+1MY62chieEsgSx6XUGIqJ
jGKEGb//V91GNOMpBYyE7bMI2iC/RPMF/JmYiQMZa+GVRTQIQIZRohEM/69zOkUq
H3mWg0BcooAjihB+d2K6N7679ifarnCcf430gXcK2KcpOicfKjDpvjHkzFI/cFdE
w3YqgwpJFJ5upyUkDMegMjI+TQoX2PENpKo7jdQ2yvloxGuX0UYsDc1aqZVf+8yB
SpGD3DrpUDaAQPD5MzNs4RHsASYrwDAwMy0gnyCfcTZ3bFPumBXed25yVZnqAXP1
P8xq6jE2ht+3wayry1AB4XJEAyPiG5ptSPFWR1A7bOl1FypemZbKWFuXchSgYkA8
VIM3hjgfzuB80TZ1HqNAAekWDT0XKC5smNzgCtO1esa0JzZUz1n8af1LPN0XCMOG
hVtY9DfdLsnQeOH/iS6+L4siZuBz7KirT13zS0PYnuyho0j49sg9eitlEcMvxA/P
hwCAtvKUrygcsCBmvN0+uaM354bfFCbK5+KzYT7I4zU6iUaLFarVCRJ9UnHg8OEp
JrbQI0+LNpl5zB6u0BALm26xZ036lS+9asupbuoS4mnieWWC+t3wJctHVS/5WC70
17PLGM8Ry54aPvJfsTCmVbqItaEo+KVim7vCwfjVZuUb6XbuSdiZVyQxwcS+YUr2
5ivGH386T5DywITTlk9g12a+xb8Nk5yBfTZQYcaJQ7TzDRwocWU4Xcu9DBLi12L2
pucpjAevZxOmnL1Ss1ZcdKDS04PExGjnU7JuifLH4n7ROJ/+sDPPrEtt7nG9UOuh
kT6a8wuZ27IjmIz2mlaJxPvkPAb2IOtEngbZbtx1NWqbdMwqsFY621v+kLbiPoI1
TojpD1f/djjrVt17PXe+WSq0M5TcL1N1eVq2PKXAbOYfNmn72taREh7Wz3Pu5Gzj
a4TB8Rdt4r4t23tDCbCnK3mjd7va5TBVxgYSQBmIlfM5AV7lwiI42cKGoT8jKoEd
d2o1UGWiJ0647W/Rx9NVF0ZnVK275ADhKoTLcKWDFF0C1xc9gQorYZVvA65AeVPh
6S/ls8JnieovrnBWCLhTFcZeyTYuszr1UhcO4nUU86g+CYJq9pyoEhicOCIHruo+
QDCdc1NDU6RHo9wdQF3NaQjJYS4i7iIcaDoZ4bTH/+1IELqHj2xJ8uhrv0FCCrZK
3zAQnf8FiIssM5SYAkev8cM6W7mWD+iVWlJ7KMm/aMnIKPLlbrERo4JcKWeuAdGl
LUk35riVyCkeWPIapkEBObRfxkgpzY2jwExr5/hae6zp+o4voQHOWua7UGT3Bd6M
VQ6T9mQ0fCCKZzAgSc7+C3WTndbamf1IsmlR4rsUCPwCoVJaYQcuBVoRdreDHpWy
vp1q8jjk6CC30xS/q4LZqaz2D+1117mounG7NeXnSf+A5ENrYJaE8OBqDMo/3UQj
0ehcRHciGmzH5bDWbH4KJXtdvkF9TbWbndacS9v5BysndHqZLTWehFyHgYoCnvo4
4wCqbQsC/caAX9v8hRlOEjWjHsjyz5fzpZMiipA7MJSOagjaO8p4yl/D3MVat+gD
lEGP+5C8OsVITe1fR7dp0mwvtxCCc3RFV89yvG7vZGRWdEJFEj7s0Sl4xpdC6mLq
y+D4rmUFySk5zZWCMJ5CKTei1eUd3WnaLNItOOmL91MoHoaXJ7BDIABC9HwAS782
3WtvxQse+5GN0M7/ahrlbExn/hthJm1Asfz1XXaCW2SdMjdiMY/Vh6BxY2je77jH
loKA3Y/OJN8GasqKivwy5RH7qr7lM1Cjc3ravjaD+bgIzErg+lPFuRt23cqBn8ua
LKUev1ukb0a3jd8IvvBMXvcveRQDjtiobMUembYT/tVPivAgCzmLlv7Spr02wevR
9qFRFbWpPAibvbJwyb/FBd3Oi1EYRTbqxKpq+dZkqULaYjFJx3PdcectFMJ1L59T
jfgcl9VW+ay4s1TQyRX/+w16ienJKeEqV0AhW+bLgTcNzAWLSvOwvvvqv+XPCAmO
S9K3uJzby/3Q2k8cCwl+/zLDLsLc/0I/Jfli2cJPt5tCPUlQa7vNn9WfeQRpUXGV
oXNb3ToZqgnoIZnG+3fxT41CvwaMnbHXdY5rwvrvuJu3FWjL8ZQ6zJbaMcVdetUw
+n5qXSa+lUGwflFtTsS0gDW5M8znA6+7oaEaCWf29ZaGMfXXyekurQtux1XaTX57
WU894EVGNQE5I+035jw69QF/sAg9bI/Qa3a0/12xKRSTx2etJQAhVWu3dVZVT+ZG
vBkw0GsURU4lHD3q83rXsoEFQBgTatMeqXM/Brur2c8ixDyoULCLiA+YcG+XuQNY
m5Sgh9JhJXuCMIKXebarLurHpqas6JLhPB64AcjZnyc61uleXp3phvo+kiRm6ung
MHMDBEeuDufimdkiYxhjJthtXH4xhB6KoBFaE0sNZmXZDdm6FUlW96mEYYOwzjNp
XvW96ncM2noBJo2Cn53fD5hWF1o/mGw/4qLBr7vKgsLTc7BCt1U0NllUyHNu8NXK
2YE2KEy/VpGtDvLJMbBPSESy7RFWLkqV+NPpFYiCPFOtEHwpqc42z6bhqPNFSj46
9PmJTnKqOq7DJ4KZwcf/ysRsRApeK3SGIV81FWvbd3Zw9GMIksl/6I2ZDZyMY52e
qYETTyUjP0gFsVqMGCLKykvaE+uDfK6TXtx1bK1Fq9vOtNGBOy4vu2F1cXTEEV8j
ZpSi5dEhMdnMBjR7DPM1KvBLkNFKmpeIpvyn9xEXw3oXdIjAfAFCgqvZHRrpqWyv
5jPfZT3hqqHf+V+Zg8WwibW12OmtBg7GyZBUEpW/T+Rl149VEkUGULrRnRJhMIrd
2r+5p3qgP4qJQobTLJJDTzW12wCgVG34M2oRBrVgmgI3pjt/JDKXSitgpdxQO9xi
JU2dDUJHI5RSwGp7b/6kuiGVf82S9O2V22wq9f+NcPC/mcEoD/0gs/s+TaXZczI+
tYdkrswVC8rfd4+ZsLKkIyGQDQWQi7keIJ8Pd7IN82zjTrPLenpMLRD85UqDyigO
WhoQ125d5ZS6vJGCp7GQ/JZ+xRfMf0i1VDAs2l3u9Gdg2tg+I4m7R8MTURbcU918
bSJPZtZVRDm7VaDXdvhdwwyu9/NER5UouRpS7Y/QSxTFD009B3+kcwklzkwP32sV
u974O0rwc0ztQMEwkq6JYnZK3/LUuBHjYTEK/SvN1F7x8oHHAazyh9U4fQv4Zgwj
GZzOh+2A5M7mvjjORZk5+GPYJXrba7ULxSZFUDBcekRS0cwseuBsB5P3zhBu1dX5
9BDGESHSJmODaWTnBMxmLlqszC/hrTelWqfupdY+YmhbdPGGAyk6XKt7+r+spgqc
Irv/GHlGktRYPI6QydY/1iF3SFXTVGsyHAFiEmpqxnYDmpH9DwpIzMLeyQ1FZIUi
ZwV0CH74WGlQJTvimkT/w+C5iBBTxkXw7FLeTJtx2Ymmdo6MTDvuXfAjD4Q5LFzb
Awmx2ydMoB8Rp/H+6uMTUf3EHUt4SW764Coad2FdqT0n7jE6Q2BAutGgBPwuQ95n
3xRj5tUsMSAN7DE8rWp1s92yzwV1btgg3Rm7gljQX7BUFvSZHuQ7VLfumaHPuT9W
MvHxzoxPeLCzFGti8o9YvT4YzS1WMpKVv8350hPwW0Mteg46fsfPuNwqR0cfl141
hG79YVAg868Ztgretdw2WGE2y7JmpIE+Ks5g/wS6NBj76uLraAa7/Z3gkBPpv7oe
07NcgTaXS18uXUDE/oPaHNaKN/5r1X0SFSDv1CoJ4rqx9dGZ8eBeZIwGubmlX0FJ
7Z9+d/qm4SSPZsHUIOxVONkVmjtNJ4faK3RF7ezUrP2V+TCpQzaWilrUMrxAarbl
wSeMrYmRT2NtvbhO9lhXL9NEZBxClO69zeTNt+m7yvIEFXLHwrCEAtDA403odnak
sl41icRPRhHG0aytxIp4juUcnBCWBolPpESCdrut8zLcWeYjyS0RZJgL9KbdhjVF
zq7fTt6I5t+IF5sNV82nCzK6DCcaM330CFOGEkS4puT9+35TACT46lwtjzOc4GlU
ovNzQilvlTJ7gZ2EuDquwDmePDUHHLP2EGXm9rMIrvAbFfojhJKITsESacLS1x+o
Cx9jnZBoxmSUFzUEDF4s3eyKubk4IejerYWxhKrr3HGdrBYnsqiqgb7md7jhOMs7
Szy6xmAOro07y/sbyBnn8MSlgUXDI5IqUKUQYV2P6PWFw2p9wGhvciVQoXqzdGbI
1MZejeHpu3Puz6cdzmBg/6Wnl8LCucqFtBg0dDXW+CBFzcwuL4Hh4OMSdWuJMOF9
lc/Z1vSjIbn3s0F9NgVO+jJ18t4yaXCRNA794sR/jdppcScvozSZDSq0NGYqZLsx
eagsNsXjGpvGNzHLab5KEMTjuhDnlxkpabnE7+bUvGZZ9r/rQaTl8WixfUUX9QPu
ySR2aqCEsVir+Wmx5TvETCj6QmJmgt/HHsyQFKWf9DtwSTJkH7/BOxgzbaPvsAK0
6Y91clzeQHzrLybPyO62Cl+3SWZi/9hCptAyTHcbISvyCSDcQqP/GIQ37N94PU2H
8u3zMzuO2pw7ohUSkYV3oqQMAZiGHAD32aNPlKA96goAgCnCuSm5QWUyiaoJt1hW
g806MDfc1H7rfJScwhDbA7RZt3A3u59KUxvD1A+ppfw1ezT1eZK1j8+SRbFd2/FH
HkxN74kCakadnLjOFNTxXk+LgsUv1oWgERRzxsaWajAI6vzze53j3nWLLz8LWvej
y4Ow8MJw0T2CLLhUfZuhq1ZisIAO+vx5IUXgOMg2C0BR9LzXCfuROFUCvAkgUtFd
8fAtuArXBuJJE1CCIONL1hBo82gKb+rMfqWkS4CvK1Kuf2dQmc3QhVIQiSEe+dF8
ESC1ilFF/xwIgkCHN0etHetHYIzo8inUp2WL9ezGMWpoGa9hlvFbhkXpmVkg6mLn
/OOsJ6c5No19PudMvNrDy8L3egQPriDubuHaW1h6gY8ZX/872JWeHzqrUp4Q1Oxs
DHS3OmdrILc7w7QLfZyRMuC+d53D3xpCnrXY2SSKJvU5grgs/O1sOzxpi07aTLt2
yLLVcV1GvBXO9d81QCRJgB4WOvwT8pJdCfLBiYVj+/9SRX+8LO4+NV5AiNByokyo
dHgwiiC9pjX3/WDTm8REK1hH/epk0XlYSnM5ebNtjPoSAFatkguJemWMEjCymrNc
rDKyAChdPEUztKKkRQ0W/jgi6Yj2O5+3sa5frDPxF2ctT1UfGdGBx9SHNEpFzWoK
SgtjHKiOXLP8IPGD0NJbCuMVozbEXmaPAkn1aoPvj1U0KNM6XFct6Iw4at9Fis8z
i4c2QuiEzWGRkHK2h4qFMpgUdjd1HP3Uz4hfi02v9aO0Xi/VGhTIagUdfbhIp9Ju
qSfXVxVgGBqwOuFnm/p5CwSJYoEtBme4+nav0opnJIIn970IG2nbG9Hiyot648Pp
cp0crvV1No/F16zkB1YmF8u6y7tZbfWYP6R2mLgr0V3RxIauV7+yMRiyWZIk5d0D
6utErW7wj/3P+cZX6Vnr5IZJAwgcMAZB34SkY3nduYkKjteYYcaqNbbAT+VI7bqb
3vsvVfxK13fVvrDApqUbmB6oU4SITEIBjpSQ4YmZ/vPNKYy4BDy/r5B50SL3bD6s
AI/3prce+ExXzaqD15Da7jEOXBxZZ++togDm/Lm7GwQXqccH3n7JedxiWOPTozUy
6NcGanhcPac0e/ksyF1Rt1l4ixJBXtoJ3cZDVKwNGkeQ2DQ7mL4J1cgHKuUI9OtL
6uar+JiDgvUS8xJkWZj4zPaIsmPYuC5m81eNAeLpfU5DtnfJYtQwjTp/rAlrsEsa
VS5kfVzvAwo91Jzy9U6hWghymuf3MYYv+dmgTjGbCa/jP5mFqeAjqnZiAy3Bflzk
mUCC9PvdYjxQTA7psH5ZytcmE57fErXG8yZep28zdt1GCiZjx4JIiFjQTg+YZK1i
iqpUXqVANBFIT7aSprS4a07a7QJxMIibjqHWrg5hKOfC3R91g4gi5S7gbOiZWnpQ
jAX/qZZnQjawGwdKVPXTnNYD8wPMpHLxo23OYvm/KoWi5cXJ4ZeuMOQMcOPTE6IQ
2QbQGIyKRtzarYVmMNlG2EKzcLiFqiXK5fAYQ3dbj9In6lJ4fD5CWiAOTANYOZAo
ltk1lMQodyxViX+xxLG4q/4DSAqKNWFeR1uESrZ29d9h9Cqs7Fps5eA1FapdgkDL
4cB/NSU8a0h35V97oqQsmsgQOpjFWPzLhGOzKcnqnmSP6NvGRCpmwwJ+i0LiZaNS
/NE1XLfu6fMY/MOVVUvvBEPuIbuzQHNzHDfOIZ/VOIbCTJmYCYSRsQbTCjY+0kE0
57tDDb5lt8YaDC/I+QVavevnjD86I1JyFd1n07NWHlRSKlJ1a3D0kcuh2rJGyZiU
SQO4pW/R6nmoU/VR4O9ClBGptjmgxWbHkboOZDFcI2siRd38hRzDHeDviH6eiNjC
+uaE4if8+p5iS6qqAlqd2UOg0TWBkrPPd+JDe6QwTcTpa8KhPmZQ4WAGFWpVoVTB
NKl77GvbK/MXXbwpi6B2mbwHDRWSXapZcHk/scMseWrtZ9/T+5RlpLwNIvdrFZSX
kjPVj5HtQP1JxIyIKVEScHU3WazBipX7CeabH9pJduJHyv23ns5WafgTJYwSMVrC
swkqF3V6zrzhuS0YGOOgtGd+p6N05TtvGa/cocw2mbiy0mgYvds3X0/wRYeyAcqG
tcrUq3Di9I3T61Y98qNkxEpK1d0S7x9eQTUwSxRUpXPPSUibpK6R7bIG5KAhyhxd
n37wi5rOgopr8mVMMuj9S8v63T4zY5sH2/68Fel6xIBxojBVhXlDFA/8iitSS+qA
1q7SUSe4uGIcZvT4ZZXogXgU5YhzseA06lR910OCitZHqlo3+ZaxK9K7MkQKuM7s
5yKcFwiOCgYnbgK2WgfcIpKHsQKnOv8MVUZ5yKWbEgHMLPxBDxkmzMuZZNZQ9Srm
mwRduVspdbPNpcLsKYrGl/kCwVD6BrDu/CwrvbQRF17QfYmmETrurl6x7sNSrd/r
u4SV5tIk5PcBk3rlSmxVCSZUMHkJGR2B4ZWufaxNnsyviSWD31A6E2ufDzy+3CDo
2p6CCy7niWEmQ0nQcunhzquPHunqY187CguE6a62KshSAWynymjTzrm6+QCRXqL4
TDC7nvYdMe+EpQHKum7n4dhFNRc+QL9eUWm0W/lmuFfBH589KQeYfesN/O+TPPeD
jSvdzoIwsOhRjaDXSOayCrjxRRuS1OyIowidGRTJammpOaiKLOVTWieGkeyDoksL
aIo4RUODqolsI0n0m6kOh4+lFf6B5oWvS+0/fAtw4dRGSffKRFUH8fuqECj8B/4t
WbxqBZgxz2QnWYMfsD60iMz6H3hj+OOXcuAjjUao6wF3KkpMAXFKv7VoyhVcuWHK
pUHTWA2YO8LwK/F4MDEJ90l7qDdTAS17aB5wI2SBA2xzFXUc3wSjoIIv0LugQu/Z
XL2RhsJmACU045gdGT2XsLDjqMsVwQyyUnzrFhJrtR0yFf5fh/UhNCbbZpWONiuj
CHkQKn2jU9ATGOXBzxxsZQnoHj2hbd9xOAitROjcUUlhs6y5ntaosWiPRA7ADDiQ
vzbdTBMQ48E5Gx6c7kUaCn6DDWCrultijdh3Pl/v1IFdn6rUmaGzymzIUhGB7gXA
Y64z4HZ9dHsLV8yIPf1uYTWCD4LDETMB9hWx55uFCZuEv1jwAPgUhkQu3nIQGeun
N5q2hHDjBXrlSP8Xel2xbKwwLJIcJwKnMnlevR4HOmhg56reK9ig3iAnFc0iiD3A
WjhQuB4RAcuNfSnldRVZgXnHU0er2XPV8+TjaciQmYvBZjJdkemLr4PAIcBoJ2Ft
2NnpsGgqR1zqc6Usn1xJhig+RaK9Orb7UWcHIjT1zJQol4Z1CZzuFDtxYFdoL/Pr
IptZokg9aBz61zCQ2xCe1Edz5vO5JhNHINU+FZXoetmgeVR/sxEag08cx4Tq2e64
Y26E72ZUCbp+B1LZ7iDF6psj4bIr7687sT5m6MSaij1+XZzw9NEtL9lcIy836VVa
pnp4+D3+XrbHMez9PdTzyB9hLR9QEncR2ypSThsWyauylWKowvRCxOrbVAFX3WRV
T0+Qhw6pVsxzPD0NjKmXXYmlg6CXQMuIY0DRlvgoX6ggXs+Ok2ZTISTrQ/cn9XGe
7n7hpetf+2rUV6YWmzXaBbqEiQheAf+82HUUG3wiagsIjOAYUEg21/Zxpy7m0B6K
3yqESvVQtBhpHxexxn1yKX6S8n2mqVdcTe1cDKb9AvwKn8++XCnqzqoXOzYtjU6r
iWIqJM+bDTRrvfMzzTxhmSl1sv97UcSeL3i1TxRvc3z090Exijf6QsSRoMWY89fC
ZlcqBj6bTyMK7Qqpc3gHQ89HH1iSVQ3GFLrY28gBwSK/q6pwlOH2wV+xFKFW4W8h
Ov+IeViu8fDgIcwreN3chUbJ+t0DUQeb1kXUFcNFXNiWlBA52oUxKJiU7FD7Lz7l
X8JfJ/q8fTFSpsvBC0ZKMaIPs8kb+kFoG5uB0q0ycLrpv9exhm5nsfQ0gTDOJLFh
cuxGE+8KK3/wi9UB0YgSvbEv21IFZIGe8E8Q822wL2JnpZSCRsC1f7iDV8hv6CBt
+3GQP5ovzNMyn7StAdn5OkiHU+rSxcbNhZxdlZdxj37UKIclrt6KmGe/E94qq8W7
ioj9rO/Os6KZh6z3ZngUc+/SQyRWPMpzrVyH4U/WpArM3j1Ff4eWy7WotJCZ+8r9
NpTwAeVNDOy88PIut0Lcw+Byyh0GEDng54UW6pUcSdNgVjRDRQxi2+RosRcMys2l
J6P8nfUK38hFw+ooippnkoyxYxRvnsp1oKXpdy3t4GuPJYQ9MYN1Qcz1u2hq/G11
s5Aj4W8L8C38n1tO5crYrbRkFIPbBVY/v3ijMtXUCN+/bNVU3+cDyFSAsU8rQEpo
Y8x5ts/nbwIzlSsY4urqKS6uX2bjDiO9INe4Io4zvGLuaW+qRaYNE6UlJiiBxGy6
rY/OgzwTS+fTADM7XzExHdgoR/tx0M410g5fBrBuM+DFdCZevQb0VyuNXYZn/T8N
C8OdOwMrV43N9nF3XWIuqysQCO7F8rU5cvWR3sGTAqeM+UcvF/HAy9eFecSQVBo2
QpvOwH20FhQsodMbDZ/QGiNuAi6QrDpsTQUNUV3LYosF0AcH6d5R7so3PYIDWOCY
Kcmod3S0hG5c/y4TfaQlg9P8G+b/eQvYBYIJl81NBkYzsUzv2s+piN0bGFQFFeIo
Ro30xXNy4veyfUGLddkqGUCZ362Tmb5Pxqo1tAf0WLoSROJKJXTwO4k7Qmmw8PaK
kWycgBOa+BTFXeDO/XWysds9gRixKrFFefp3S3QADT581iZ2FT+AOz5kq6TVnBl2
SIh2HPYfGVM7ICoxRhiilnzfjEpR/03PrMM6HdzCmHcyGKL51ZmAFUc4XUYThW1Y
5zNTMFP90H4noi7mxxoNclG/yO/JUgfYhhKNWxna6pV5DYk5jdFBt2P4NB4KuZ0m
N2iOMU6d8NaetKc+KmUrhELznk3e4liDr207/FGaN0xevhaOWlJJYOk2CTNUVq1v
e6CTBUxnPN2uVjoIpuM0h6XeyhknRXnec5vTks7up8FMGKuE9TnWBYOZTdHS2wgT
k98gQWbbnMBoKl9K/YLMNJKDrpHtjd1Ycv5W9C1Wg5NU4VgwzVSTvqcLt9F4RsU9
BbWCla7inatjEeXD2sIrPJ/Qy7zbZHytprsXYaJ4Hvto/H8j11UkzblUOMKhzM8g
DUrKul9BK0I8TYCyNz47n4I7s32d1dpancx7wErtE0+qkArHyaaHe4WBni/X5u5O
clLhnR+iUD7SnyI9F9t4jrIYTbLvr0J+6g1dzeuYCBbY/iccWqoDQHCee9yfQIfO
w98PWysyAT5EnvNzxyPCyG41+N0KYhrh94VCs8X8t5M93D/dHV42Pma18ZPBtYVq
bp1Z81ZUwvvgyUbqm/Xy9VH4CCprci3/kuoXyszywnpTEeOJpB26BvsyeGSy11IH
geZBdZLxl0jHHAb4jAhha4BW/bQpOcwHqss9lXzkR4MQ7RhO1QX5Q8tpYC3L1dZj
YSWEUv0VOccxnDa56PcV76CQiOHkn8abRuTGKI2mieLdoiDJunIOGR2qfYDxFDFw
gk5/Hvs3P07QrQlz0lqjmsx7GVsMA7uua6LlfdHRCSuBbtKmSPuSCx6GzdMOndC2
jwDX/IRqgNJsJg33BxT0l2/Mqn82Yp6trWKgH3Pt9buTgscwAeN1LJSqHg43Vmgx
5Qz4dH8LRSE4Te1bfjNHygrw8FYStc7fX8PlCuxzc8yEeWm0Ccu6kqRT6Q7jxaZh
5QZCuZVxHPGVBBK24LU1rYOlVI5J4Xq6w1kKJ/lHe+wRaWd/kn0UW/iibl80UXcA
6MauvigIVOc4WnX1mpHBQAre6FjV50RctP+MKESxWzK+b820GJs+eGQRrPQ0ilWI
XhAO2RWz5NerIbS0yDQhyG0Ll9tU5gD43HrC8P/nr+hFYtHtvdJyfvmtyAGUfS5D
gXcB1lbEpqOIpgwT0jEmXDyYPLBQkg5kG0ckuaZ77qKjy4AjkH5S26IaPNuiD8/E
RwLkNAM/QMfejRjuZ5NfG5bZj2+k5M7ojusziUXQeK7BzahAl7h2qTUh3Rz7OYsS
DEke+5RSzMG0g39D0higCT+oFAUN6q04Nu9eIKlSUvChzibMyZDQvgFiXOYnshHm
ycJ9/v3ZuhnPdKcegsigGZJCH/0yZRETsvnC6oDGh7g0OAUxjKgnXhOG2mf0rBJT
XQmZ/4NNedtTNK5bgTh2AZCm0/P/oRLC9PdznsQNjoEeskqzSWNysftA7ojcR/hb
cyTQ/u7HziULsevcxIw5YDY/h007vixSV3e+Gv2YTDDxrlxouS+qzUuzr9Zvcqjv
KpnvmTkQ8wgXS46X2VR84iPl9Wd7RtYxUsPEpItd5529RSys8oehXilS7o/KwAH/
Ak59X+vHkOBoI5ygadQFIUns1I01mwPs6XzKDSe//BwJuS6as8H+iR5aqyc9ilCZ
IiQOvsom7Dg1pN4S0iKJl/vG8xgoAM06Y8Lt4PH0eW9raa1yjrx/vH9CKl1lDuoL
DKgN83fWWOVqkCWFeIg2huppLyax7BGG7CKNSUSXK5u7hDh/CLnfCMCHa0CZCk7A
qsA10xgoSag9FNgrjK5K/xB1OmBNy9eJ90JnrmGVzjpUadzLyz1ne9XIL2oRlOoy
WuqIAzvbikSFyLAkoV5xficpw4YFC+0IgUV0SK2QzcX77HqKpKfy/9uATnxeNlS3
tuS8d5YZWI4x9GQgCLOVQeoJmcEJUuCwUe1CD/dGnEpLBlNcA06wVDY9pfL53wGn
BHEbTbDo2f5E4cw50/qXfN1ZUQC3TfzcfC6i/BoI6F1SYlny4LQJIzwu2JM1pVMd
KiFV3fK+wGbLPVgR4xc3M8o/41LxpmIVWjy8KqIuR38rN/Fj8+AUQniPD2TQmzAp
NZ8pZaQdlZXyADMLkljPJV8Lu/RKoeYG6rjAd5yCXLtwzA1yq9s2PkifhwvWCNJn
qtzFUNn4UXOHQ1k1m6oCwPutZgu9aLm6TQKKgLYvpPcGHgVMKbLN527BIWytaoIi
+SkInqaDXg90kNC5BvShwfvm7XIEujrvq+WI7jy3o2HSP1K5NhAEapDNPv0oJZoC
oY5/LBPdu/Myh2XgtrjDo1HT0aujaeK1LzJ/xgMAvj6fpoZ+HdD7typMqnthkDKK
bBK1OhX9AeRXtLr99hyL2xPA3q+W8WHg5NCGJq711g4IkVa8mQKwWVPasDHH20ZZ
wyFIoVpFHRyBDkIfmfW9KSBFGkbRDno4PvLYZwmCPXBdkIf5oSmGQ6hgvVl6921B
W9ydrpViDvli/ICcvtKl4FzmPO5xh5Rg0aNM3HhWMHvEqBh9BP0ixuEZHh1xfDD9
plJBDTZiM485xco56FOPXFSGeg+1Xh4RyQinF97eVZXXTITjodDUwbpvVJYyirDX
dkEUJi1su71VyKNMZkyDrDRDu9ltxoiphu9wDFXP/5YFtwmnBt9wPZKc6RPQEQjx
YEnqslb7HaSOLuKqMms2rDrpGe7WvtQoXjrvnVjsHelpYkdNDF1N4k4cQ7leeZg9
yWlz0omM8uxWDGRtIWrzmiIwZqVj1iNCCM1FL+mYmlerzyBUk7hgnQOHmtdVm3Tv
9LJ/1IzluJuuYZ7ossvBZfRw+5d85CfKx5n20XNzCakx6fl+8Jp8oT/Ss/bel/zy
ESnvvmii7xaRSrpuCD85SJULLDqKkV7ydy1GH8lBupXcvYUNm/N2uPS37vjYm/yD
p5B8aCczEhfuaBroDRKXBjXBDqWXALmkx59I3gw//3blVv6J/OSd1G80WvFG3qA6
yGubbrf32d8Nqx4IQaR7gsGBhZm/yLu4+KfVY0K5WVzHrIWRcmnHzGjigq2snKfW
+C5n9o9rn3iTZeO1kCM2bKPGReKtMLLxacrtL9b+AkefkHF6N+lty3wIsS12dJ3K
5GNZSQldLDGnmzaQlI0UxHvCrnGPFlrKTv2P0BKezl7haJ2qobCw/lOltTvOBJge
yZQpYPisOKf3KWAc2El1Ypgc17qodgAFxjZqyJP8z7KJm2oAJ7ki51ic70OAxe7q
FPtOPjnV9zw5po7TAG0qfp18GRGd43j9lqnAZBvIgJlJDtf/xxnW3hpdsNTpQYcb
6acLh5SSYR/eoybx4t3U80hJD6r523WyeVeQjbyeR8CV3u3+DWl3ChRVAcOUQIUl
/xbKNpFmND3L9YRA5yoMuWd8qT1KGAyhxchgWTbmS5PnPP8BUBWhOlLRxPgVm6tT
uCu0wJ5mPboQy20Glf0BoQrMj1J3wSVnXzYCpAd+tCsL29CVvwLW5qxQ5Wxu8atU
VrcuMgCLgsvggKNV3vwg5mI6wWr3aCTdmlSmURv8gHhpLPvrn7Cl7Oak+G94UXKg
ENiJb49Q4GuACzLc5Qw6vf0gjxdLJFzrqTfJK0/qX3nd2TVzPTnDB98mUduwPnbl
8xYpKw/9Hl27IH0cjpudi82D4dyYr5SJ1mkZRjI7Sg8s525b+TTGsxTz5W8gpnIs
Q5yzKPVnw11+gj3pE9fklpfeH+sA7ujT9fw8Qgbb6hLPCkoz1xyS2i/ly05V+en7
HX+bt8/cHWmvBIsrGrzWgDk1SIdLeJZn/PpLdibtJSd3UeDLegNrdNQJ1zKhe8Ym
X/WigRhgmTCBS0IEQHoD2McdfRW0YiZBNCliTxIV/O1q7E3xS7byr+URSRZh97fv
n/tfJFo3jQWyxNwsANamANw++n0utkWwuNzYhAC3SEURh1ltm9n05IW0WZish2pC
H2scB3hsJXnFuWEsnTtG/17saL5EVN85vN2jDGxtrUIseX9oco6r6zpTXRSfumyN
fle+vPv+afg0FK8XlN2V/f+G6aTUgFOMRsSjqLjVqP+51goMSJcD41dF3B73hdTi
6ZBHHU4aXXetNoKKbTma2+QVa12LDlflYiH6Sqsi3FcvXCDqPexq1stgHDKrBwTn
s3cjq5I9HSjVGlgJTHD2mtr5Svn3pvDuoArjqqtVhdTzura741X+AFIJJ6YHRjWr
VxMi5MQeS13qIwMGD0e+BGAMlcNubueK+rcGBkly6cX0HWMMva47GHtCIwSlPsT8
OAqjm7Zsud6H+hTCDtdne1MWfKzHIVxMuQudLCKVHT2U6JAEj3R17KkRSbGY8UQJ
/ssHthmZaIs9maGvo0LA4Ql1gH9frokC5J8cKIlmJOR6eN+mPLLvIX0oL+scxG0W
xZ3F/Buhh4VCKRmGRXEZDYua+sUy/luLpaMUdlJMhUIwlQPBCyxfjfMmx8KEnrEf
2b7eONbc+yHB6/t6PRpsye1LwEMQdtOy5fuLPaWuZUgOnwV58EznAL3rxb064F/h
9wSnDMKBahrMs45k0HlhG9F8VmmrVjehR7xAbJLVHQHTKHjF35u7hMYPIPNdmbou
/ckIA0M8KFEL+2TMpqmVjIuPTBwVodNC5MSc38dmNi9UO1UADCf65ewFjR2td6cO
GfGmiT40q/81woEaS5TPKlzLeUk3UndKdILgyDxqIxLIWEFiz6bq55g0NlWrJc7N
S+KGz/9XLFKfupUut3pOvo/kD8B50EkFjmleceHrzJGdZUGu9ZFNT38ObWj44fVy
sKTzrxAsUXp+AT7AbzKcGrrMCKzz6hhMBy3VlZnpZPqIIFl9sU/yQeKRKRc/5VaL
BTmiYyMc15QkfAe0KIgxJNVDR6jkrl3W7UJ3dp0bHdMMlOtTdzH/5Ks2y8na/laI
TfjMnKFRl8mKZTeZFQFoDOb83tuoTijF+dmQdDH9vGfq3/qnLFdkMR8e6KhGrXjL
+etor6OsRdYx1cuZt6Ox+vFDbALNmnb2LMiItlBxX9tVT6329B6tYe5engtYO4RR
9pm/vziFwGdfEuHvM0PqVhb3tF/zSA7d2eF3mH7avQHeL0fAe8dJ/I9m+Ktfv3N+
kByIsV377Dt4OTZ4Z8YBQlRTXW8eeq39doiaIXZQjWkKu2ka3DmbfvWEh9IvTj3i
zwYMbO+aLomn/ABpPkzTrhltxK9QiED87vcpP8u+2KxC7IUNcWOMX5/9AeKX3pd6
ekzcTWaseoUYZHTOQmad4onnkKk4jFNrWt5TmuqN5wNYFqdjrqlP0scrJCdSa6sC
wvDVDfyt4GqHrumf7p2WCNcL3Tmfa70us1yG9v3aEWCpSvqaX5gOu0/ndYkRtbQd
WAEgV5yPDTftI2KQE9Ou693fiAB8nRqipgfyV1p/AoH8WPKtsI6Ko5zYTIB32rZK
eVSnoyhp/BBcMXp0GjezLpzALp0ToZKjhgZKFtDU9XwnMhg835t6XYKi7x1PexRE
3xMG33n7zxNZj6mRoLSSqm5M80X4FVytpQ9slhXCgCPVNJpYdXi9GCik62bqJNXZ
Gk2Jl1fNc1EkteunehBm/arGqz+4AlqHGnNgd1BmkE2oefcHHCVEVaU0kebDfCqf
tBQSia+xOnNUZJhfdmshhhgDo4lQVAUb4cmoCUWdSG4Q06wnfhW+7yYY76lqaehJ
KMKl8sgIp5Vihzggj1S35lbsPK04cj4FkFatZmpI/FlJqorYLlxxUxX+xS73gHPj
iNVaSnSg1MiX+35f5yOsOMpPadmZ9HPhEcj4gbAKt/2jTg2vUMD3RhSXIAecVCR1
C0wZJkIEWvSJWMbFrbc3lBMy3cjph2Pi0eK2gfUIpko+fNn+BS+hbMHXiUCLbMVT
m3rz6m6mRJUjqlBSms3QPbPVTibRuPlw7ohMyJ62f8ta8EJqPW6cm3jBL5tfXIxV
fZUd+ONVORxrWODtQvkOqUv07FpSvknIOVuLS/lMwH0gnWrZ5ioQ/BYtRnhDGX5z
Viu5cAfzYKVXNy5nrsnpzVLZSyZNHj/Hsp4uQ3AUNlU1i/T6pBB+/PZ0JO/c2xE0
H1qrqceJJxqC/lStM4cVyEcqRBgHLFjxvccvwAkhsn7nt/TRRg9Dpnp/m9k8FQVZ
o/419bV9PHRutO+c/dkvhwxivA110ePeeTR6BT3NiPx89uCnL1jENNpudZWrx7jt
n48q9GjcATwnZoBa9OLCwnpYj8zOmxXH/S1iKb/OJX+9Ee0hJqUsCJgPpBwy3n77
B7AdSrIypmEENmGD5GMcckmGwl0dfqKZ7zfpWdRqzaWguF890gCVOiQujBs9/btd
xTAh2ukG4ByF29A74kw963LQZnSP/j9Ub7blAbRJYrI5DSYiPOVo14IQ+wpz17Nl
Ps/g6JwC2JSCXYNvEmZlAJZR+rSXBhE4IJjsrkevs9p1qucAcUU2ZpvKViLrepAL
jXFpWVazX6MZR+a/BolZsDH7pvbEoXq3/6Lx1Agyxsly9UtELdhBvoj3EdoSiVt6
X2Ls/+IQuYzYXgZ+MMRygdvls9zHfyOmGPQAZtZY05HOCTddiVGs1BkfKEqqpVTv
wH39i72NBbC4k9BRPIgrkPQJgMHhaCSltMzQg34LQ6sLk4pp2fZ5ib9l39Hfn4w7
/gC0JdckoB2XpFOkU122oDd9F09yIsOHmfcg8b7+PO7j7fW1yypBMfjJMb3RiOih
G7R7Iua83eNPIq12jrWHT6DXoMjbuNolDYTTTiUqqyGXzD4tcGCjHKK5d7xd+4bK
2pOWmgnG6HifxxYU7tp5ErE3sUIwraiozujx7cJpCCYPXC1Us+wzm/DkFJUE1diO
oaxQ+x9AdyW+5kgl15/IBxOOUrP4kKjIBJWYk973iZsiUiqR0tslXfRVdti7MQmF
QgXNJ7qduhNdRmwammEwoUlSLooD/VgYS/CWt9O/2moNhKjg/LfqssKXZsV+rY4O
eXySDYgWXLdz6h0qLuF98m1pbjt8zmz1jWwu3AcaIuXk2VB4Fwho0iORXEVCnSJj
MEB1AcZmdHQuhL15HHQG+8TPSpghw4KYxCR/W0cbiFgppkr99Ovj39rWHRcbbffk
PuAViNa2MPNdo8CdUeJANQWRqxeo4qL+/HV/WcmYOJRLoWoRj38IOAv211vMF0VH
jgqQI3ZfDw/mXKtDzCjN1eQ4jM9TfdnwKZVVUjwakOXt5ro32qxQUjRlqxc7S13n
fvTEfbcl7IZUl2hIrNkbrtpsW2cVAU9bwuWVY5+JS+ovGsuqB+dq6kknMoGYNUa8
ufBtUbrQCr2V0wfxx/oqRLi9+ZtVFTvHrOxHjsQkRTfSLsx6yBmamPj9vO3ULWBK
hSxWhJbq1Gn8xmY0stbDFhD68gtBmlWruvRgArVbLVWAc8w8e9Z6eCAOv1/HLCqe
nqBUjz1jedqHY2p1nIjjF0PC7LDTm5jzPOons72GDuGrrDMs3JiFv/tiNv2ICnpD
uS+UV/KpLhySBnYBFZ0UK8dteX9o5Mt4VLLPVcyRUO90rTH+Y/sKtGDXhc4n+r75
b9FDrPn4ev2sZt3ccOmRgdtmHdmO9o+RwRFbqjXP8XP3nCAn72UxrV5i1wdyM4TY
YCYbmARqqxX2pSvuq3hOY68rpqj+dPm+Uydq35O7xg9nUGAnMprbxnTD8OhFQ8iO
kBCe97vgEeqAppgaUomkX3l/WATxoF37cvI/oJ8CanTKBHIzzSquIyob/e3T7jEg
pR44Ic2Gx8q5asbwq3DZ8onXXY1PtmGClfEKm6xs6c3qsKS9QqvbkWSz3nivUtQk
w1btCEGFoCqOtIlhy5jwwMdceSzKcHX5/xi8RcLtsq+eKfyuRzGIcR4uOE8fbXbM
3jZQBj/IT6s8bBXaecgGITI5ETJsFnyco9AYdmPST0VKz1qFfLoQ5+Uv44FSxvgQ
lZazVpb0ghfBf3z+Jyxuju1y5imhuvc9HM1h3QV1mEmO5XTYM2lGQJ7ZOtHGlwuJ
Yy6UYNeYF84tUtBAYd1Vmrvm1j3SWrKKg7Y36w5SbF9lvyMN4PHg2hS0SGzq/mTP
Poc4tAUB3QKCG6JKiuIXzBrd8svIuJ/GDInRe8ELzIeKcaO97AE+qu3MJVcHPKIt
Lcsp6CJHbKE8vQ/76J/nEQ58Fr2q4UZW1ljI2f9Sa81hMD1SUXRh0wA8afimvFLp
40yZEmYSi4N3CDtprJtcSHPy6slyecE6UzpBkCbG/lS82AntsD12JkiR+ZOG6FVX
4gXzAvWYYoUg45ZR3NCIRn9w6UKVuSbhrHJy+jM5MXpX+hN92Ln3jb5/D+fE6mJ6
P/m+mXqXhRdwgNSKa/cCyVwwM6i0ptos7hdg3zCpgOsmZRPNMDe3a0ZAp51QnBVh
5tUG1o6f2ipkjjwmrFlnreqz0256bhEjtXbArG0NsCETi9NGrcKvprMrDfNShijg
5bwwXJyGwIugNUG6qs6ikVccDKKS2MJNtuDQKsoWLshilW6v4fl8nQgr3EF9aOpy
bvOxrCHnP462CAEht9pa85j0UUHEzMenMdEd4/KsDM7kfH4LKSpqsxniL+p9bf1m
Lx0PQPRszuEdQPdRww5/kMNr45jgu7vnmjTzA7aVcOahL6sWjkxRUc18Q6rOaTr6
tE8mWhcHlPqY71y0PaqGSbV2IyKS2e4ZQQ0Ei+ioQaM5UwUqf4eID/eIB9RMvoFP
cdm2I4VYgpwhSMJVsI6bMuO/YfjrU1+MMgCmPEBMV4lz7UOV4EJVzmR9XCS+rn4N
kQHiZlyNJ7mk3XMK/J+TZ/diecBBGt9ucsgxdZYbuBu7EHtnzoYReWNs/UqGropw
sgfJ0LANGTYyWpHXkuDZiYDDe9fOj7r1zgnZRcaLir2l6M0LjC1M+P1K4hATFzKD
vHlLYEUdLiDI6OD3wMscaqL8/T814oUO37ydXq9a8LbOnFIiJjv1lrGd5xXiydLL
7kiRUjnK/6Sem/f03+KvSG3NSaxgmG1tc/M8rtXlhvC5DSIEzf4TxcWRXjbPmENp
YtGZYpHim4evWOsKl/j8A5gWT/1e84+4pv/QFWFKjJcvuJ5u5DNYnTzZTb9sPL97
4MzHQhmyjyaIOjycl6kDyx2V5ml5Dlb/y+Ggls8vLH6wK3+vO7kPt1f/fCtPBXrS
EhWDsZctZAOOTA6/XgvsSmEr45RtiG8T+1bR6HHyBWo9qD4XKmKbm4nTHZ5z+5Jr
7bjgXjTgwhPpTJG15Zek6pS04eZqG80/oKC+BTU5FnTeAFuZLQXdMUb7VpOFOARK
k/7vmzWPvhipndUNXBJ4Sc/KfpDZVAo7YIHtc9aHdU8Gw6lhWp5SqqKAJvdvTXmg
dcxzTsLsbjxCHiFDvlN8YLxwoXYXV5v+8REHshxWbV9emIJaEM1YQ+DSqzrIna8R
ReisxD0q5VgP8LjyoTm5I9zzXWNIeEaRdv5OV82Kef1WyhadKzOHNw5GLvpzdfKS
gaxPUQimQDMxLLbsOVg6xyh7qs8Zwedq2LUqySD0KvUL19k6n0po0JcJhriUIyad
NvAWtAcsII2SCxlv5drIs1A4eD+9v1Mt416l8J+NHvNL71pBbuEZlMZg4OwdQbfk
ZkpqBl32saWjqQBIdY5N4nwOZ9wkKkVnvyiXzbT3/wF7tW6Tywe4na8V0rPW7QN9
5dE1JGdvOKgRwMCWrqqdcnepnsPsu50htwAudE67BIitC2JUDbY9bqsdGtFnEzJB
1dGlP3kTPVsXRpJd6owLOhEPdPEJO2U3KWlCnKfazk2UBoLVyJ10W4626MQihYOt
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LajFc2UWMOFGohP7/uBJVAMj+1ovnw4pfRb0q1D6Ttsnc93x0G3eTvQhECCtvyEY
VC4fKsZxaBRj+Ydl3tO3cGBAf+skd8anafM6UpVjYmrnDIHkVaTaf/GhUZf/ej9X
AEBSDuLcd5908OO6DkSJL+SU1oiaZttVO4gtXQ1JVZFDToLJD04oymJSCyK6vm+B
t600npiKBpZjt+IfSdUHCOchuPksOkgUT5jGb4Ico2LHbRrNUNAr/N4xy9YQs1Je
w0/lHaFKFZO3+uy4KNj3ZGsf3R4L3+5A4e8i4A2u+GpTVqNRIzg3ITYTEvMPVGBP
xr9ckDjJe1QUledt3kBCVQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1248 )
`pragma protect data_block
oQ17dRVMO3lK9tni2ojCHl96Ckj+MmF4vqVAiwGIO+0SzfKwn0z+onZ4L58Nwg2d
y9UclW10bP7RAq4941ll0SfQnkjfYlGzG7NyqsEZgoBOP+cD2+gw6l8XC2WrzI/9
zRXDQExXEUOHxWJe1uY87/ydtYdO5toi+QqEBRjKs+PWc5MF+OlEwaO5y2dzyGqD
Nnmdy3OwsBCSgymF1XaQQuVleYKQq2C85eKiZSy6CcYrGfIzFZaHlQceqEuDnQlf
BNGLb48ha8tRtGVBzZSbaSxPx2C1iyILCmQeZem1em0iKw/kL6qmNHQTZT8j7c7t
icp5ZXg+4WU4pCl8TLIMMnpOO8JYjTjRBpQdM1Jj046zER7aVxQhElhFbwATfmMX
BjHbiXi3LyMtPZo+gV1QWnjor+FWGlMKSqiiJWXoxNkzU/0BFdnM6Gwmjoy/nEYa
zUxs5fgWmp1gcSLIlv5Nnvl7TYujtVJEac6G6pFMtPypSmseg64Y+NvUiyGmm3zc
1jqT63oHJg9hfx8luCKcqsIa2RyoUMPq2BdR7p9PrroXySTLpVohMzAfxHsOPZXb
XCb0lK1ZkdTtA7zb28h7CwIhijnLAbPzSRaI034nGZ8AfV3Zoy4R9selqn5/OEjr
S5WmCE/N2wSHiXnbMk5uMDn02mJHJLLg4htnTCqc8TwEBjbgJFqiZ7R/D6qBZjtT
4B8hVd1YlBwSuseO4McME3RkjDUJH5di8wVe8SdbWoyIWshuE3rKRqvUjMh3Rez2
meMpJLLBGt6AXHoaI4HjUVix7LzwY024eJM39IP1zV3spQPIENx8Yyj5/KWV4Nry
1vtMAveH5gluNH13DZAs8t2RsSyHBhtUZg6TiGbKQPjydG33UHa1y+3SzFke34Ft
1ZX6PnloBUllmmHRVvvg8YiVX++MGt3WLPwNWY6KebZ67KTyd9cqgJ2SY4KrL18t
Cvu+EQXriNbX9U/VLE3jKY/2Cr/KVott2nlf/MaSOA1P7NzFUrL3WvmD5KcDP5JI
QozZoKe/o1nbgAyCuuunX+zFQEckWR6LjwcKiJdRJTZkm/9KYYczvQullevdc+pO
unl3SDpWWhJ2WocGDhEon+AZo+vujGjzU+dj98ShLF8Ra3H9eljNeFvvPAgo5jGm
okQc8aftkvE7uZ8ltrBMowt8AHo1yhxHWoAdSK81vhj+7pk2e0VN3NX1K+qHuX8F
JqC4J4ybQ9SfC/wiMd2W/G8sp3Nshy7D8HdwzfyABiq/1oZLMvgrGhy82qrbhdtC
v6tB/UZqJvdocrd2GZd+Iovevmg2IT7i88ESZea3LQtLYkYuLVye7gsgcOergdBM
x8J+fvdv0MYETnc4yjkm+hWevmocQIzV0Oyp7b7RhmANWz24tO53+oknoJ0Uhonp
w8xooNRtPFdRsHDRKc+SGksxPvAStXpEnIVztTuIiC+3CHEwLNz1osxjNk+nTjX5
afGxqEtLasLx7i4KWNQtvTmv47uO3Mc/MnsRagB+42aonxmJ/przkkdPcghO/Tt9
2aGT+fDeTINzSbD3L3zAndOjYtXgcrsvIVZowGiaLVpaPSjIYRBGjINovGGLi8Kx
YziowHaEwG44DnJeRD9+/bVJnXe7Xjz37ax0RP1AH9OFAyiwJ97nyMHggz2ZcaYj
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jcMfHFLglvTXNh0/ZgjJuAatgQoSknmAvNZM5U+q9N2GQzQZ7n0UVbHtjdLGFcuO
ltnQG2XDjafkQe6TCBA2HLJt9Bw2VXbIWmPcxYbHdzgmD7GQxVhVZHc7v28BaKFB
MDWUSw3Hqx8uHdqoImQspMYxuRPs2ytf3MonIXbAZ/vv2fU4lqzq669nnAwtSVMj
VfMkziwqCoKHx6uPKSfVs0K5DokolS+47aJL/ztOtb5UPVd4UhY54kAnVGbiyd8d
dCX+1s9GpGV7omEd6nBQHolvWSCLV8gn7kTTQ1tqXRh8adQ9s+O62vMBZKIE32Q+
fp5bEJpFC/QHAvRyP7ub+Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6672 )
`pragma protect data_block
SM91JsddV+1p+NuT4NPRJehVVZwaNy94LAFgJF6Py1Fknjvsui4trNosKJzpP2Iz
VL8Vvy0Zx7U/A6hUK5tpFMy5ePA43ZKWzzLLGKiGsrVAkFZeTsU0q6jKO3LjHD3W
P3pIR+kVjEEZehm31/mQD9mBtroAbEjRIOISoCMMcCVCmyPuEDncfSSHJY3AYYc/
mrx1ezCELL4bw1RRRBPHDQGRT8XGGeV9OpYJCbc87uBBf/jx7rN9uAjaFJ0nUZpB
P54uGXL/UNdB/8y9lqRyWyBqJoeKTJ+z2opHLNqVCCWPw1+MKxtzZGWQ8fQT+pEJ
Mp1KpFfXZsQvMhTxirTRpXvPi5oOjPeuEGiuZ7tLp5KNLgTS8WJcDLHjswGgYeYg
JXuV+p99XbXfh7/GsVBKdaxBIwqztHxwkynU6sd20WDcJsuvd2X0kbIktIrMrE5V
rh+IcMLFq9a9EXm0fRZwZw79StT/ak+9chM3YA/k2u1Tf6L57+eccdcI2JKJu+R/
p4Y6E8VN6kzKxUylW+hAcIn24cWSWgptNCnQYDfQWSqyeNKjHMeFkaZpAqRngK8+
4sLcozvyKQJJXjOsqV3kDysTh0rpDIkSW05Mw2M6gmxFeNvUSp91zl4jL1b46eVi
MCgJOAyjv4IGRgb/Sv/s+aCsHDBhrmYg9v+0JjtZys22f8JFREPcS6S4WZYGD5Cp
4wjR3ln4vU5Sxi7vLDRmVusOr9/enTtx5kAptAIqxkSjg6Pi1UR9+J3UEYGuetX2
Bcq8cH6yLv0oNcz2MZCGLmWTyRHg/rSmUR4YJOjHlLGDMWsaSJeLhr5M1mSQzvWu
PWlaC0eJ6/IBc5hUPavVZZnlM4tUPZE4vWtvdshZZOy7A+sCPio1+0MCrRyV+ogm
ZbSysWPeIJZ8lWMEnZiC3hi5hN9yZ3Z9832ET5n2S1BK2Lf27hQ2YBNqC1reil04
MvnhDyHreu6YllFULMhf+70h1ZjcQK0S4V/8EY79DKiz/8IbepjUO+AXHGxm90m+
A5Xlq2yBceS6duZ3PGxAIYy4D94297TeWoEHahpEbO69jbdmWsD8vmOcLmbB8NUr
FRCBOkc1C6EyL5r89QA17O+/ZxSN2+kE1rgcwJ/yjIooP2rnBGnx+IIdo9lmbehN
H5/L4DO42lPP773Whgk49wymu3f7nxVfCXm/YmsLxdgXby6izEHoiM36UfgZf4QN
gcr4ieMMuom8YeL0UMhT5ZJXeu3fe1/254N8GB+PPDGsuSIWVAFT3rLQfaJOhtqC
HhhnkmaD0+hOePAdx+eGpL+n7EtkpOq7xvelOJ6wbsBro3tTnWGV8+iTWF1VlkpR
axAVOtshVMS2fKinxaoHmO4t0NNIF7DaiU1IXMLStRGlsIQJA23zaUdx5jvYTpRX
Hez/8tkGEIei+QOm39NgeCHodGoR5ZOCsyv51vhQ+ewvbMGKPVqZmcZUO//xnIz+
Nj4yRDrpyWWjlObaM5dGs3h8dG+ltOPNGZHDr/wqufJNUdHfNFE2jP6gyc+Qg1u4
kRH2vqwQdwg8DZh9g0cPt3OZI5007nRGtc7viYlAkjTrYFH9tKx9MZmFLiBUhLDM
RTUE2Yjy3UYOuDzFTfQFQqTD/fep0DQmCm9e8hdZpW9t7xuE9oYDI2sesBuol8+Y
pnA85V09TFktalhEz3Pu1KDQQUX0oNhNTjmPd8IITDxQqnj4KfJf/KCfxa/WK596
owmMcLv6aoGyXfGCGW5TeHqKnG5oL91RXi5qzajKd4em3sLExljwXft3E5bIrLuv
atpIvXtvf6B2hi1Ffs/kJUcGODgewobqxiiONtglDp0l6QQ+RIo9+8SmJ+75hCkW
LXCiBSea0zcw3/BmDzA+AuGiM7fB5rlUQHRge0na/A/336ZOJxYPx7H+DWvuEugj
t8Qu2U9grgsouTSqAud9iCkllzK2KrvjIFVkrm7lkaKg5aam4dWcfRiBK5x5POI9
7fZqIxwfwjLLYNPBOHV/75o7k1MaQo5UR+/6NGqOAa9zkBB4O73nbjag7f0bxhIU
iMG+mXELUARh5+Nn5jYPU3lEoCwQl4EmR8cgDC9iTUBf90gTeo0IxKWRUvjzznKI
rNnXAYmHR89hc1ExdW9/HbXiY+aEzfvYICjN7IsNkz1F/kFJcOQ5mmXnLQ3n6gRO
H3g78imwh6m340kbY9gbCYNwJH71QKHKjbhfgGGMJcGHJ6N8FKTH5wfvWCpSDE40
UxJKqINrqtItQ3jZgbTseH0hrtNmyCRvgRK1ZUrOz/zDz3A4VzKbFo9/uwjzA/5T
wkcI0i5R+upV228aZWl3wewa7fQSyqfPfuB+EHpZWuAZspibhYEPZe5ksGsFvnmG
qxTn8JgGaKKE3+OJQRRwp1Qy+7QKwopgFDClnQ63fxHi4/Gi1FkHHVQRF3gf68ev
4FJvWv7t/Z7097tQL1CdQrBDxqw0crJwqQAl9JvMFYQBEo2JpEI5jljCtDTEETex
NCAJUDZdMDPzZAZIplSKqCXFy7/zFFThMuP1W/Bqa+Syp9z6NCqTVWwl02J/Om2w
MkSGowLJ6whaca4LxOiAG1zPNCnE2a/iy118aMrUbbCIK/eQKx2TEG2dTJHpKjiB
gq6aK/cEdksSLgJk+mzWtFiRatg7a0Wa3APLJnxLcoDJzUttge46/bV1t1gkT7cQ
jjvo1s3Ey/Qo1cbjJbAtQ/bRgrD1OSOcNW2D4G5Dzr06GKgM79SE4RukcMjckL6k
X+ALx0Jc/BSkY12AlNeXSLyMIuZInzhe82zlRXiFrKZ9qHJJe2DAWDFhJV+EcZWd
HIyIr+ev5xj5JcyuoXsEmjcEE8Pav3js840RQgrIk6n0srNEUvLa49aLiuWBjyOc
FI63qo8JMIdZZijsmFMlyZM1QIEnSlf7TuDi3zd8nRy9vkeLqNYUI59Oek+BuFSF
2h/Yip7qaemvlyIhgVmVknltG7AeMafZ1/YcALac9NDGE/08Zkj+X4K7OJKj6fS2
x5T9pnURy0TsTwZxFPi+OI4a8jrJkTmngchI+5KWK2pwHf07rAvoQHFAZO11Udlq
uIV80OnHejRZK4xPwZN5KoMctdshv0/dAfxjPPLnOe+j/Qg50HHaSCLZlG7IGRta
NY3mrME2jiphAP/PNuvWAAfuVXptYh5NfTJ/qc6/993CyZm3vXoEyoMUArMGd2WT
/6gaZVNdn+t9CPrQ/NM00BNQWiyX3pIg/ghL1h4LLVqcIoh8AmagZ+1bGb7N4RoY
afGz/tvtrfxrgtgxDuC3s8lcrMGnRSg+BX4fYx6pUQ2JbAa+9CRSPjZbLXMUlFMR
uQk/1NTfvwE+g859DMz//qsenPrcEAYmCW4LKiBCQYZMf0z58n5h4xrTWYpwjQo2
JXchJ25we0nSuMqI4NQWtqUUnDhqNgK4cahxCIIVuIdrJrVqy7DlcWSkfk6fPpHS
FVXeDtL1DIRgVR8q1d47tDTqqt6qFvMW3SMLVbegwIqxiNusO2O1PIultedlBb4B
5PpEn8hiRZPDfjAVxj9FrlAZAQenMDY+bbD3uFSUn5pSrXRXlHbsGuGz7OZ7972j
ju5YXGkq7KyazE0/9OaS6h1NUdIkI245Smkohk9hcwualS2nhPluyJE9poiwhkXV
B6ydbP1HM4Q6ORaLeKvEz7XJ3Yl928+UtrOmFrc4dLWl/QpCjAhHD7p0wLmchS0g
FbZ38LdFvwVUEJQgIiDsU0LvLrmuC4ccLY5QXsUtFuXSfSCF+GYn5J1mS3sZ10cH
anorCb1DL8KPTAgmoh97xOFnls/pOXBDcUCc2gnZQ5uIDio/IPivKW3hKfSJxdXP
eIsEZzVuBdHXWi/lLwCJbc9DzBO4YkZFhkKxR/oNSRqsBGqRLAOPs388NNwBnf5r
J6rly1KU88tSdHcSWww8zR6arro/clPUosToDv5d5IzUEQ/JtzGnk4vQqPokPLCe
hhM38KG8pO82ybTxfJlXLZ1gNhO0zVkiSujRsgwwlZqYlfgl7KVQp1CHfy6EJ4Nh
sGaWgY+fZDx/K0k+Y/N1DpRuzgaUcaxAxT/ZpJCqq/PBiLuQyfSC7KN6yz0p7xLL
zeGHYGlz+MAEkqMUDd0IgpZUgvM+YNUNZv3p9HbyOQjxX9C+a/0yOfibnPVRbmY1
MTIWgnP+w19KwjzIv08olfAro/VKOj8QNkirXkaw9/ha6rPTRp6+p16JdIHeFVRl
MkvEKHI4ybfF+qQrAzWUumYMBNUaXBGKiEhNK6zGoB4abZvtDj401l8SJb8MP6FH
4qfUqL48VZ3pBezrXtA/OLgUD8QnHzY0ptkne8A6rNEiWLJZ9cTlZAY9YuzhknjS
BxyOFaR+hUs705zug780R6qkxYorBC5A3FOO0T9e4fujSSRRLpz93377pMul26c3
K8hAamWt096inl66VNhC3Kb2aTP8ps49Q3LUjaEKlMaCnthDZMpUESSMVzrtrlMY
jWyZU1YgV1JWVCZGa5I0N5I/bQmv6BRcD1crrCCrgZg6wQMLNlTqx5WOOTu4IGXp
gY2wCyPgXHjZAiJ/n4Fu1ZKgvuSHLSn88aoHpXa60r4PT5Hd8sDw6J3Aen9m20p+
odkA+5G+jgubNgsYUmHaLNrR4nn5LhzFrUyUZ3lAwt1fyADz1+XzwbkrfvjT3uw5
aUZw1ccAIKLpHlJlDB4qAHLJm8TZ8qpMttOkPovYTDOgmu1ep1CR0+hgadfm3xku
FbjvO/3Ep1RZEg7/59MoCUbIAGjMhj8cAQd9iR0e3eQlqmMUzqodreHUioembjEP
Lu2JD28d9KGwUWU2ngB4vZoJEj3geyj/XpB12PfZniz9DcDo928RCCC2EyXXPRJD
dl+uUwHYZsj4aFHhvJjgHpSLnoR32R/KwAoRNRduGTBWX4VCzTDPvu2rscS8uKpS
XQ2GUxUFjJiAUdlyQaQDcVfH6GjuPMjqqYcFjqVv2WLPZCgw8wian8kJrO3KxnoN
MjG1xJGv599IPvdxTeKYl0iVUrrkOSw2FzwocS0PNo+dKO0T6IgqYglp26FlOYCI
jN6UDIrbH29Ijlw7XvcA5wrnzPeWJhkmiI2O2GqW7lNWy8W25R8cfPzgjvJSXrXh
A65APHM1PTYwBboyBUtyVYgWu/MPP5moo1db20M6or+oKDLYeAIxBrKUMl3CyeQv
9K4kHRHK5Z2GpeleTt4nekzivPkQFg8OZrBJ08lE8mVVgCQ70hc5DmyOG63KXGt/
/bMJOtvX7BA30dDqicmHiOqy4n9Kg0+DkCjVWsWcwvFnYS2QzwoSQUjxIL/f/YFP
3kQJOXAOmdMI+aQV8oCDjFAFQknvxZjd0q/Ytx+Alt5t8zQiGJG36VZrTYcshKmU
fL5H2uzficDkjKRQqTjsR9jhfjqpbCx5DmJSfNyOPtVVW0X/eCZk5LnM8SiqYXCV
fXBBCLsvM09BN5SXm67CyFu2/tDNexFbSDLSJHc//1unVjZf7RkeJJ8lQSPyq9fq
6A4TLs/XwAnhmVMQNPIqUYl1GHDuZG3A2+wDainc5CiErRm3MXf5iYXAtiCjJlZb
kv0AhF7c6iRbuFl3cheSeEviuncPhYHGZ8s7q+gUMIYqKNf20fDDtzSzOrhPTlwJ
wR67OOrGNOphlS5j8+vpEGUhl/6SALWo8d7hDyIKArcHQSe2BfWZjv7lEZLiFaSs
DkiFHgsB4Cf6aAGjIFhDn/OI4iW40GmWlU9h5j9DX9L3isg1cI8EM4yj8/TDvC54
PXblC04h7pLgAOofe4AsbJQ+NBIYatJlcK/pW44SRllgY44GLziSGwDrMacDjv+c
rRUHxs4jJEQw1/gVxQ4A+oTfxsqd4CMEzuVByFpAvxolskjMJIfTF7F3BrBJY63J
v3ebLyZpb1IAMhvT7rj/nOIgsN8ucY3Kk4iPjkftdtDM5RiRwiUx0RmqbroXv0cP
2vZUnkwA+7pes1j6mH8cugpYk5zWRGnNMQdX+JLqIe+JGvFCai0tZ3N/dmC6VNL/
3aQQx/nEfy2e7xv0pQIcT0hjr0FbFthIdEvu+3TaMGK/T1tNycbLxoH5lmsERgXz
oFs+DzHwKAR0lY3M3e+B22XiKn03lt94WEmE5tARrKMOf18svKOGKMFrpzdtY5Yj
VaSg3PK9WOn44Sir39t4gSL3RaPf73SiukS0Blf+gDlvylqznZga0CCHPg0EnLfk
g9+QXj6z98kCZw1yo7RVagmPT3N7yq+hyw4hNAJ8+z/QMzuIjLKcx6E73AQXD21Y
oYNwBX5Tk+FnyLtDu7xgSy1+dxJyMpLRrGOO+7aZTLr0V9dRN2rNxjaA07jo5yEV
QTfFmcCW++QbgrLoTfOqP55rAoZsD+QGBbl6/ZLzDRab8qcaB8ZGvPn8lys/upCW
bG/0c7HPqHrvp5ZLriDfwzIiLNfRys4wMIvpYSsZG9DdcQLPLfcnd6zC6ZTi+/F+
J5vEzTr+2cGy1KDBqdn3+BuioQG+4ESbWbQp+KWECmaG0DNQr0Wd/P5w+dof5omT
84aWCDTvfbuNSEl1kzAvpqbJvfnwCzqVT43pUIEohtqBHAmLog80644Fs87QofGR
N1WUAuakY/HPfl1Wj//Ax9gZ2LmCugRRiEQ7xDOZv5Z3iHnMBGWLOgbb8ENBa0BN
3ndzSjHMkODyF1Z2sZrOiP9pDhxnIx6RVgVFTZ30cYIHhKTb1rrTBdc4i0H549KE
fCP9BUL7rDTZq6tIyVI4wgTw1zHrb8kAT8hwPnw7rqPehl3Qbwl3pZmPg/XKIj50
1wXVdixwE3mg7OXemCskmeKrYQOxFfkNbQelfpPbPTvsCrM+stGdzAeo+f5Li60v
kOQWH0Xo8pyKSP++lLG/9nymj1i2JabQEvaZiVIDP1A2S2oV+5S9qPAEEJK12Zpt
joETcVtt2XXbRXopGZ0VSuyvhWGmgp0c2pctLsuVr0mXpInHN4J47+aN31HiO0qj
2XPHM6SnoODFq/QGSHZJSIytdmGafeUiGUv35gLrinGhjnPKZIrclg9vMlTcWW3p
EXnf2vtQIYoq4BqbLwbViCzWSK7l68+aFDPP97h6O5D8PsE0CKMvo5EzT3zhv8zd
URVMZw7QWnlQNDMRE3T4pfVK5IDKxXaJcmjfw+nVwUkYrEmlP4uAln5Ei5XBpVPR
ReSC1WSllF1SwOwvK3vutKL5KXrsY/HUvAHgppcgOQ4UgzOxwiIen4JxxtgWS+yz
qbfrv3N7KiV1nWklNQuXlA+qNYRL81WXBrca6yRTo+21n3BxhGZ/5zO/v+1OMFst
VqXRMb6VKY2xQ4S8cWIWRZYuxfVKZRCAaxNvE50rSRrWIHNTvOigybU5CKk90lUg
xAMQJHgGCBkLyJsfrcy0Go8b9YK9nt/fvym+Dv1zseegCCure7N+uvEcoL4Jp30S
jZt9HOycGvTSSzFQ2SQz8peElT9Erecq+bJAUqQyehBn30h2H7N5DD+OuZWUSWwX
VIT3N4zxbgANEvauceZ8CnjCCDv9C1kZvp6qbhmyeJhObh7j8j/PmASRkQOzxEkj
sofPEVhu/a85N2xC2CCxUH9lDrFTYbMZKPnuQq3qH4HojRnWcD93l7ExTMCGC06R
7yOc+l9uqor4kX7bj684Kv2OooiLTjDxR0aSL7gwQubHmgHUj7jTq2x3GOR9CmYA
ZLh0Qzde10JY8V6mkCukOlb2zvnDH7dSLgL40ryZI4nQ9+vL7+vNKAnSSd1HrFKO
vybpkwc4lfQ09aldJFn8KJyxEn7cAfzkBXZO3Vv96tP/6/etjrD8iQBrWjHBA6XH
g9NiqHyRTkxX2K11I7GASPMc/0J9xvF+DNJ1AJT+sdkkzcgLWCDivr+JnGZ4t+z6
g+9i4x+2UtF/onGexVQvlylOGzBdCVo7bT+VdKSx1nFMEvRhTDMK75w/sHg7rQHs
rPSIThOmuC0Mc1Dlsw7sTvzZ3CXaFSUYl7a4Q37Pk+AtSRiQHoerRjcA2Gd/gAvO
xOGAFT58Z5m7jWXuBIaeCKj8N4mJw0unB66JZez99wFN7YBVzJ7SPIxGpiL27Pwd
2Blw2g85zpGzhiTCxLcuHXEIQ1HY2psD0KfoAeS0GBnc1UlqAmtXTr40+FWFYGvC
taWLiQj4uKdYpinGTr6Ot+tXEHUyCHe4NuCl3+aQG0DhFP0K1dsPFRUs/r9z3fgG
6N3stINfQhXtyHsXYyBBHWou11A0DfypKQU4fmavAEQcFe6s/YaJ0U7aCJGD3tMT
Lz5nHMdjcAgahIK0+kDfhG11KuoocV/N6qaGrytDUCh5Ghl1oAHwfQt8k4EwAZI0
yop5RLZYBnt4MblK7y+MN/TLtL2vh6lz74Mpi5qkVaRnJNGO4WHHpUosHq8Ksfln
/Y9y+Jr9PhuhU1Zi0b7fHbuPAlDMfahCSbe7V3ycHduO+stlpv3o0IUBy2zZl00D
yUjc6t4/YwUYWC1A8OhYa8ExA8/6RZmOwHqyMKxZIb6XP7Tt3Vd3KsL8FtmLLfNP
ZpkcFbWloGtOU9u6JDu7279PkVSEW2p6GyM7SdSuCqdh1jDofbRK3rq7awioPQso
zsTm7q2gMKSU4nfAwk6qUD6V9GENjqwJdfue8xjfu5HBQwwjDBYU3WidWQGeLDyQ
pGP34NcR1tJx8mek8VHNX7fN23Nogi+Uy8DRGT2vmqXCcKiNNrkRRbA0T946gWcE
yX+lNRk5gKtbf6oSKMUORV07znHOXeQKJ9r7k4qk/bugr2BNXhLr/rryiZYVuLl7
hxfy+f4nxRNDYSjoWCqSE4um7EZFTGIdUN3yVPFschcemJD7m/yo1mpgHYFDz4kC
mG7UBKpSQMyQsowjUT7vg2J++g1xRhRu1y5FgiqBocMsVpamIoEzD87ornw7w6kC
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
YXpCsWvvhLEpBM/R8wJT5SRua4Epb6GpRgYvGvqOAWVftaQwhtZ9GrTyWFOH4euV
R0lNy09YplEX3l/b8gc47XqhfG6MW9SB7yhNzNbPxNYdzEe500Hx5Ywm1TgFPDU8
hSnLAwsaBMzKWgwWINUc/isqmuLEJkkpp2nuc92eopFvANeAfKgh2WedLT+FasE2
ez27WqlOdrqQZYddypFLm5GSl31z/winDFUAw8vS55uNkEJu7+1v79IeGs69fpyQ
pID6WQerzAnl4EF4b7qs7o5ZBx9wU2MsglpTlAvBoefZNbPPrHbzgi/SNbSpYpS1
rSjCdKwWNkcsvxz3h0AECQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9680 )
`pragma protect data_block
b5y4LiXxAWTFxEvLjzfkOra6BmYveXcsWLXNHC5/VUAJunVd05XAqmNRces/n1Fk
+1shPQG3rScuRSamQdeXuUlmzCHwabCu4fzo+1dkr2bfC9zFDPxC4KJVVBm4Nsx8
fgPdUkC+KVwij2QZit6poFCzNsy0u+iVKc9W9dyQ/U5BTzgXn7aNz6DXypOparcq
FzoAPYeuVfvD4WrorEz9chuKxeHF28JAscEEQEGzrqCsUAz/ve1w6tG5KKatGjEn
H0lMwug9ht1rQwjECvn2XkCThmyX/m8o/UQrTsz9uHYL8UctIZiO6Spkze8y9pnD
wj7kBeSFYxKodyuFeyLN4c5HxuKXBPmSbpZzIRkpV7nguiPeMIudGA7DUWeJWZ3R
g1oLJn+0M0JI9hXve20U1eNNxAzD+bxbMu8HfZjACJ9Gvb4+SEStdlqAI4SkVG+u
sC2P1X7IMz+j0LakAQS//lXOoR7QGiMGKqgLXxpmzxj0eT5zE4rXQeO3/Dti4DBe
lqKodutGd6oXV/Jm0Yy1S10xdkmglys+eUhGZTgglzodQ1fTp8tP1D0l2SRxAZuI
0pHWAFhcFE/lky/LBtpmlZJdfRQH+8V+tRDnoc1+vKygwx0gxLORqKDcRJYrinB0
CsNoGouJmP8AZEkCKS/B0zSWVBZccubjhgbs5cTQWjMY/UT5C6k8uKOnpkKzRk5T
AxGhKj8R0GnVBv/Dp8Naef+SgW8r9Kcu+ITHek2hhEjxe08nTctVDOXvSA5IwEGC
QZzRCYc62c3vQ+qOjg/5kfnCPONtx19MRUpWORc2I+ZJNbaNpmUBBZgH31vlX+9j
XtOIdXLtj4A06vj9eR8h/ymxeIe+MOLpHFVTgZIFaCQE3cQCiH4e1pWKL2ZHcqhf
InOjWYnLSSjcZFfOgLYn6Q2MSeNcYw9YJjguXWhE1KBm/8Y8/C7YIqJ6sKoAciwC
0UDBsw4kADxfJvuKoPXZXUyce5et7ao8gMu6ZvEOTWFfsP4Ng9RFRO3GskRrpvac
AWJr6+Th0heLen0OL/5QxGJZvra6EvEgyUN1FqENOO0lr7sLghozyQCQuIqAf8Q9
yCHAZt+gnHGRV/brq4d94qa0yofuLej1LTR/6gxlsGwaVtMf3ZeG+cjeI2tPurAi
zL2j2I41fTFx9X/UkGX3y3WswA3VtP628mtAwO/FrbTt4MHwL+PvHnl+HJ+xXN9l
lMwXT4ro7h32sGqIVtIR1iocotkNs3NuwdC/VBGHcqxHYCwSsYT/tgl0OAdo1jMg
n9E970h8RHFlOji1i4kCQ6XcvwncmJE5WogdobgChfc/DzHZYeZQs4QLjZwWnIlG
KSq0aSTtPf3W9QJDGWvCx0V8UE8GApvEqwta+7ASpfcIxs845lkV0QbOmDiHg5On
E00uXHxg4Pwy6r6JYEnk5faz5k2XnybWiYMZC+q71V/cGm4rn+0bsmqGXqkVNoJS
WIlYGSKHLFGZwO4l9g/Jofc8ncK32kLbZ46XX1WH5lBBPb80plg/xnNgSMN/NHWe
+ygJuU8uHdmylsqYFjpZZxWXmkuMJ0wdfRbSfSLyqTgrQW2+d7CIjK2ccDt3k89D
Gq1d3NdOkepnLbzOjRLTCnkt79wMpn31KYUNKAeYza7x3BPZ86QPJtKVs+KGX0zp
/AdlmRtwhrjR6M8nRRASntFdpF5+YTJlh2bvpIW5HVvEWw39OtljDzC6WdIfk7KI
tt5M6vp8McFM+qrkWClRCqmfoYklmCR4HwgXheoUmBy/LS/4N6N0O1jVjxDWHILg
DPtL46CmKmYnhaZMGWtgZEplQvLPbjNLrfVgoS02/5/cFTRv/94YB4fPBgjpnLI8
NS2fgMlbpAaleKuDbouoYtFr1gkEIFIL7fYP6TSqXQuw3T9yjraiZjQsnhEXAivK
NFWwhik6dznm7+gM44q+hjyCCPXQru9C8qGTNycnPE/LacHtrZqry7sr5gS4wisj
m76uKTDoBSPQ+S7Ngnh/Q3uKw6kS6VQePywO3E8qkXxChF9kyuBOChi7AmO+Dy8p
ipqoMp/weQxcaCgKmr0byV1thHN96dQoqcg48zdng4oPmdMr7+E6c59R9x8gVtNf
rvAt/Naq9UnnKZQlgtKcnQ/040pkFIE1jB6IJkQ73gLJizkptaZ7q+Yg1T/BPvNb
zYVvHa7gnv+35yEmJ03tTPuFd70Yh7hywNdc+L+P4G4KN1wcHvK42QJMZq/z5jOP
8BI4wJf1fGVGNq6hTjxsClMCcFZp3aOeRh9xanNqblLWzj9kYX82tg4Du3ULyaWK
M/gurqAbsQQM+RWVwuC0yIRyhUDC2EcYcitLyrpxu4zxmUtF3xuUuxBQrcL0egX8
lLHNzvh5QTiszmYNzt8GvdE87oK4MOMI8fIU6xQoZJcpnqKDYWTnZWCmCqmFGUne
Hu4ukqjB5w/LEyFsuiErRT4KDWxdWckxCtqmX/eAAtwussHVIgLbNOYVlZ17HGmL
sugVEEDS2rxh7dJUlVB2u8H3Bk+EvYAdGmv1w1n0WsbeIXsORN4pYpE+K+hZrlYQ
XzZkbX4EgyVAhoOh7ziNFWXhxPyBleSl2q1LftvQ5r+CPpiJSFyCEQwUyj6l8yAA
OvT3XBe+vP8GdbSXm6enuiiyQtrHK4FyG7B7OlaG2fiyASTshDdMEbv6sNNJ4OqP
I4uU4gm2H+yI1z2MzIrYrS1kxjSPp0cWY4AgW3WedlJaJKKarzgoQzkoOCVnaBRr
QAVHqVIASzoCJg7WRKKiIDzoh6TVAI3JzI/WO4frestPMpS0bQXDIEfJQWkKhVJ3
+xZQ/noXaXgsHGhWG0+GJXGdPSmJrJZuEHYJEAyLcLfdc1F9/CXHYJpAuRxbc732
3L2CQzwZ1lspLiG8EoUu5cjuUqxlRiQt20iLm72WeMlDblqjeN7JaC0bzRYnlwHr
eAmnDkJnNJWfbaFzNxBSgszQTiEpJc2nuf73dhIO/UxE5qazmMes9aRN+jXJ4bYS
dcCd8tqJcRR++Rd4zbg3hiBkO1zElVGey9bNwMiR8dRyybPBKcPffP49AF23UXXH
Ps17dKja5I6C78xRSyDPRihgCovYe2ylpwYkFwiIdMm8ppb5oNjRPtwuc6q7H1fa
gmJiNJy2WirEituRibrzAmcGgRoMuSjhWdCVcKc9g/pYRtrgrTMc+l3W6PtoKGux
DHKgx4KIjqJGU2fjFi13Ina7vh49hIJ/xT2+O5AELU9vS1JEqMGGf/gSP9tRTDol
/WeujI4XbehTOeDZ/iobv2x8B9EOWOnQOnuAEI5tgpbiaVRrbQimo/N5GaUmKQm1
M7fb5UJIZDHt4LMci7Z02VabCw5WCH14Lwv+lZwLYMxOFR2WHBbtMjXNnZVu5bjP
f/eNX3ZmLbnVM0U92nfijbsLGj5Vk3EAtNnOnNLX33brYDscHk1eRNWa38FLsgTj
1Dulq6PF0o8Yt7SPEv8jt7ighkOiHKM+qcBm11M2Rxl1jiRjLzdIJS35xpifxlfr
SIeVXYyWDLXAYilNMDIsfCXFvdjLEmWRnQyJIO6b5Sdj3RSsadhgeIi4UX1PwkQQ
RoGBqSCMu23hNiawzN/HfAhVd5xZQwzRyKbtIfRiMtkVL1KzF4PZG01+t6d9f6qY
afJH4opvHQ0Xcc4s5dwjFnd08xEJLycI1oyahpSPIoWZwgoGR7CryC6OIH7MrpS7
Y7g0+F0MCZEIupHIy0NRlJxDhWVUYJvdmdIS6M4TKElZq3bAVxNoYuyE0b+Pxp/2
sEz8o1smKwBDTIzPCEc3ZjgsLU+ER67TBcZzAQzpElqU/M8waGzubU5C1VVkuNt2
srXFk2hglyEhKim/fbpdQsCsn7xr5jzhZC4GpZeqco166putsZf8o06BzxReNjSE
fol2eTnI5C5ErVGRkz3TuS93owxcVQjaHQ1LprmZwXLvoDK/gAI+xM5VQqspTzeG
DFUWsO6aIWWv/DgfUe8FtYe7ujcGlMKr0XvfqNkny6lGpisqKovKy7PP2GKK8Hyl
idyGRVhOjD0kGig+LeGJcLQgAuEWZi7BScC+fBOHTKN+Yn+Jgx79hko5ztcCn6Wx
kBEoi0cJcXq4eYvwbyKj2EVPp+bC0PO3ZyeXvxqQ95ErFbYt0m/CQqh8PBfyaGkN
PqUTNeupWbA0jO++gZo6LZcF9x87x48vVm16vwKc+wFWYnsNcjbhm1os24AkxieM
7x5R2DN7daGMLRGOKHnHNrpgzdde89NAgtAkefSFmFdy/tSJFqGj3xos96WRfJjt
PO6dZTWqo4wBEfpt1UipD6PMcRkfQ09EM40jGebJxug69ZcXakcbN/kd2KwGBpGK
dUDQzNhSGLzJ+iSs48y8GLerUxvyRjsGDlnRJUrlLWSAacmjD6PnXr6/LKDI9MT2
8N/LQ3VjZhCjDnX/bbnKEwVlXHQ2B4FKZZVLIOBO7NHSu27TIjWZEKT0z9mgAF21
oMmAYiOeuu7Nb8ycKV+WlvwH81YMrCji005u5PZu6IA9WrfhDzLnxZzJlUedkIWI
8UAxCCAUXuLITfYwVPeyIuXIMaZf26szm6MgzgIV+1jnSCrF/MAV65VLS0fJVg4t
7Dyj1WTZND95eL4iO6TydBJmTak9mqw5pC4ypyZlFsA7+YlTiewhRwQm/gYi20bu
Y0+Offu4cxTaLRjBV7yiD6OBYp2PuBBrsAAWRs0of2lZA/pPDOFWCR6rMZy8Zn8R
Za4REc4/7HJ+R2B5Dg8cKKB/C5suRO2jHmSwNWG3D8BylZ8xclOgapar5RxctbnG
IsogSr+h8LLhSpTkhkgZekHuMk4MbuxJnrr3xTC6w1yCUU/OhMDe7VzS0Wx6BFfs
hfTlT9ra+QioROkNMeY0EU5sjq+MM2v+Zr2Lbqnb+z+E8PgLx+ke3y4uyXOikhUZ
+uRzYwTsUyzecysVf/OQW70s+zLCqgywEMOP/2vuntisH47hKl3tfBGsa3xQ9o5K
qxDh62o7kPFA7KdqXwW1fIpVPocKx+21ofKHjBsGhJqVNLrTmJsAu65swtShc5VG
B4h+AkxeBg/Jp+oATbpymCiBKt+8FD5dGPFLMexhZPE5oTINX0xgZLSgfGrRgBMt
duCbFEyCrRud1jYrxIB1gssziEYaNMUO3fCT4Fq1zzGOnzzoPLRJXhbdqPUkaDwG
i9VcdGrKAbESaz2qEvQrbwX8ap+FeTq6reXSUdtoeGSH21lT64+tQRTDTf20fzTu
KMPuym+qSpf4KFMy2p8WzVzCq8q9Y5t+DB2Y7U8s8KZ1ZNH6RSWlUWAnNxnzX3Xk
mGP+3ta6qyktcMihPTXufT7Y0xfBq9eCqhXoMsWsw4j5wfbtkU2eaFOO6zSFSADY
GRqB2tb4ibgakYjT08Wxw2fjVXlspcUrz4zctqdxBtWTMe9N6+Ui3z5RCVLuq2Mz
rjOk6OfeZ6hV8W9+fPdDPSs6znM98U88h1ZvP+ZRWgcULs6/4q5WblYlCD++1gNt
t0Os1jRH1KvgWKSwpCUge80C8ckUuU3871dDu+tBxYw6K2TImI7EDDOTnlV+IBj8
7+M5MG+UbPZ7El1EEahjIwBvJoMIGA+MzBrpaaDsOoXtt7uurB27XyGLtbCz/9+P
145wYI3firNyv+M3mdahhabSh4jnDGnI1ZfP2pYGnDjNQJhQFrkuI0B37t7bdgDr
ZE2uw+XWIyO+zcrg4Yrs+G6JfaT3/zih+/nMYjHo1C25+8sSAV6D4HMrpMtoYxUT
L8LOrhVeNi8Fz4nq/lPB2fOKJ2nhkzkW8qXE4mkqPSRfF/DPc2Tt+edRkSAUCoyB
vIGQKHQSzt2xTaFf+xNSXS9g0D3+GFiyQCGKGfPFE87Jq57xkFAvEIImgqyWaSF+
fKhxSL075XPnQbjivBpWECPCt2cVt6zxZCjI49pjQjs/PXMhMFnBnVnAp8mNEP3L
xww3qLP0daL5D2k/rX5LCUI9SfrswehP/FsHKa/t/dRt3m8nXotL8UXiubu9HtH3
FhwDkgRBGdwGin0p//h0zLQPv2s9ytc9N4nadpCQAQGMtF3qFBx7jNUefzcVpvcI
RyeuVJ0CsPx3ATS1JzFI/4DF6dyQQH7GYYbEPr5xiMfa8DCzttrA/7tsIgFkdV7l
QMCVJOMWA/WwnA3q0BG+eWsikJ4qODqUJspt56gr46OXsxtZhZNKnZDPu5rzpLNP
1VAQcYYcEzxXsjBr2D6C4HCc2/VrI0JYDAcHeha139qbwb58T9Gbpy66hjWQEt/G
03zLZMrf5rBOwo7RT0LlwfVkX8kMa3HlKjfLkFxlrbR7uvWb5ozU02g6mn1OYwP4
OjMfuVaGP6irf6IQWQzCQxmcjazmSwCIBlZq6sRO95+AsPKqlIYpYAUAD3+dxu1O
3cTQf5aVsjNZzU/c4jwK/fGEd7jiQGXVmAl2pZgm1wvz2UjThbzP7UStv7Aak0dd
Yd+DNXFWB3c9a1k/ZdX8h7v5M2nuNnjg1CJq7Z8Yg9bDiIiEqINpphxy07UyI5o3
cGYHiSLBZ4a9IJr6b+k261JItJ4W4uud6sHWcP8/pyRIFgL1mW66yNl8W1ixKzqg
gGhXubu62GyDVLGEeMblYBqpNpBJsz5kTEa6nyBX0VOMpC/GyVlebRX4JArx+Dhq
a8rHfcB1HYoRdk02ltouYHGR1WuYTk3RxyFcyig3+9E4dsXqMCqTRhsU5tNP3Dn6
73lrim0FKe7JhUjwmvn10gGLN9uMq2IPC6ilj/z1qmVHxupClm14SeV0Se62ragw
fPMqGWBhBWY1gHZ85h1Cv1rQx4L0wtMA4fo3Rc/lq3EldC4+1IlLXip365s8uLZv
ePIH6oT/iM8UalzHjQjhbuJgyQN4EUjdiYjjATlyOwbQ36jhXb8Hh43jhC3cgEdm
U/YHJp8dUA0/ijtj2yGKEeaSyYWe3Jj6PrwENg7kXGX3NNe7dSEVWF9IuuZz1mAy
Fjn+NX/hQfQ47en7RvGdfmSL2vr2qFQyCTnhTmgZR4e+K+gKAY8CHB96aZYAJWEx
jmVN8e+37t03TQhdtyuOUtQ92JyCtWffm4Jsjgy6rbafX3cgyA6D0fAdj8fPHyxB
HXCsw8/UUL4+lBGjyMjzuB/SUjFYTuLMsdasaxy5LZS5L+x8JNU3uYoWb1e7SNhJ
9ZuPa/D4HvGO7iCKWYbSYWgHFZYSimXvVy+h5c4OohIiDntOzqQzCCL69Z3/EHvH
3KoiApxyZp9ul4mAgnlGmfo+E5W0Z5FH6EhHQAUwNNvCI+/Rjm7SAf71XpvJeBdQ
uS6AOCe4iVt2+JTGDwM3CiAbevJZ8Cf9FkG82mBUTdAvh7qooc6ctqYXG5pfJ8FB
A9XJ8HUKwo3HbXX3/a/Dp5o4DPpLKRF21TTa/YcddI6gtTzlt1nCdDCSh3pCXsPf
mYQfFV4qHVhPmiyZS2wOeokxM6x999ahhqJ+GKASiUpTtBgIL6xWMcGAYDivoM7x
//1ej3r01NZmX3QKIG2Uy6hfwBOOd+vFwC6R9o1l5Kq0oIgMCWbtf6iprDjb20+V
ZfCz8AEdjg9cyjzaz1BugCr2tEnD8J875WEt+VXZ4Z5n0f2+OzqWOnalOM1RFpuT
FX25GMiBUVsqt+SyhL+B0Hp2JmOjToEA7OrwgTrfQ8XkqOxSj8GuiNUOkXRfh/ef
TNYlX/etf8Uqk+Kdl7vuLl3OPo4xjGHEtTgSfjTVlBX0nNk5ZtGX+EOY5c2UlsWL
dGGt1HbXEbsCnZe+5ba7QHgG0OOx0fWq5daP7ANKiIJy7b7w034k/DKhn/KXF2Tp
sU6wlpph2jojL3Deud/mf94Rvq9h1dGEjyfXK9neSBF5LGDLLao9S4N58yCShsdV
5jDwZ8d/mSsvt6EUwm8zhGpl33jcsg193qO7qGl26WePXWWzS/XO/FFLAUrLy9R0
A/v7Okh8BXYRhNiLKU7VRCsOpkuWxa4Xxwp7HiDxHOAGQMB8yaWxfyX7ffZKfOtT
Mq5YQNjGRJtUBt+SpJIkoWraKeTFWHOTFEKsYj6vXkXIzCBw5MbS8a+IQ002kFWv
j80TycVTP5YXrDLQqM533bdix9neEWOHnjaANxRz1Soe6W0mtFSkgaFuYI6VSZwv
V6EaVDjFxLIohl19i5lwzztfVLOTxSvacXdN5D8w5ww5Ik9T6qwYrrePVujDJFWB
axOrxJug4VLs1cSrQX+hxprTdT5NCRuz5ptGWSborUrEjOSS9Odpa8Us+EnzHc1/
MEeoTlMRigRs2hDhg86Np+su3McQiSSRqfFFrlKHa2iZIiYL8OASQHKk/EaPVw5C
BiC+Yr0JsWWAAn9OUqzISy4QMnGZgB7DjRQL+eVSCcDjF4Plf0hqxDkSWGKDIngo
mkTlIw7sSBzYgYxA27LIHIjncgudUpraosPk77WhrNpOx/17+5METhyT2ScA0Ex9
IKaUQKm9tCL4v4hi1tPK9+yhJZHk1O1LqGu6owsU2ror4xk4wJLyicLm96ZLV4/x
ONnFEG16LSYPrToEtNm5D5NgStrDr1TYgxbTsLbPsvqtcDIpnEySCmirfK7oaIDS
gwmBftnjybbJvi+yushEh//SVlVVuL3f1ohxBItNny6e0dJi9NpFA2AzvaIUGC5C
LGBnKCQPZWhLh2k06GfMmDVQUq2gx71LrkQRUh8cGQH8WPieEMVa+oSTiF4Q1BtB
ugPAJxrdUxrP6AWoU2dZwI9B3jDlLTmuE6g5NE28WKuwqndSOPdA41yL70YFq1aH
jco/1EZoU41D2C9M9/+c07tJTTZjlVL5xElS0wE2Dsr2qepWipVMoh0/8oVxqYYS
k2LR7WQy4vhOlxxPLMDuBEmOZuZOgqrvrIFeuxeArsEPb/AidRpexXj7tfipovWP
3Vt04NIIevDlNCPFYU8QPs6DdQKADU5sIGYCF3CAgRK1X9u2V+BH5QSa5xdmZxmo
uxYXc5IiQZbuUbmb41eZA0mu5C6YW6CifShguPZnhu+YLloK34st1bQP7kFoeG5D
ee14ywYToYGdJMbY4Kv/s5PGj7kJbku9thrvoirIW8yh7lELr79FOYJFgA4whV2y
tqxwzqyahCRmiF4jeDxhFak2NqYQ60i7o+1Y0tAAoF20xNUXfbTmr7DvSVkp/h5/
XdMyvsTwv+5OaKDKaCrGLqfTgzl90E0Uztj0jjrJHh9AiBjMUDXrKaPfZECK0cZE
rG0TJ+FuXYFPkMRVtfiVaAB0WPBgpLr+GvrQVpI0Z4Ztzb0a06e9tMszGYwflIzo
FrwO4YQbZ7MY5BfqF8DqpJsKTDpzLPmTARImJUt6U2UcwV7EsGob26WPDzQAA3lP
mUZQp8coyREyIQwHetFAfFn4LXLktobePlTHPn+90dU7h+872FH3SyvnUp0b2+hL
kM/1QdsixmhiI+27CPWvJYrhiDMeITm0LD4jcOyUdTZFcHso3sa551afgxDJ7oG1
bCbsNrC6mmGUB5rysBPa6D49mbrWPjawVgNQh7viHYf9bdaILCf4HnZCAXe8fDmP
fUW2GGIp9llENZGdDtYGCF/C07VON2aw7K2ZdilHTEqResNllTpvzXYBv2tFFUbp
7IZFZwnaWdEVAp5NhVs6Z7nrbH1cELX1uFIxIOMYnIQHz3HlXkS0ReGz6PuZzHm5
x+9zaIvlPzQUPxhHDVAg3UTohQj6m5yQ3O0i5CgMSQKPRSAV3F0XDf4MaFuNDf/n
zvdAhMYvX3cNbUDnrJnlpBSD1gEKLx1KXHj7yzlK/iTV2QGwB0L6WtuzO9znFo1N
jFqalFznkytYLF9bXtsrxza9lSRFdtkArSIhXTsp1jUYbbB1HXhxeksi7p7bxCgO
68FFVsngfa3em1HrBGQTJjAskgAsKfhrzTjL80uQn2NepRpdmbuZwVFOjrLVKqVX
GUXVnbZFVZ1FTu9eHak+A9Dy7vOyrSB0XV+XY17IegcJp2gvfzbRM0Vv2JZtF/6v
2OaKutKWcwKNZDBJCSUt/Axa20PYi4qE03S987uYYpDBgqGSdZrtQ3YkAXrZMEG7
KxLGxDATZjwbmFzqOdnJMRHQ0SY4KX688mBbEd132C4MIyzicgz+3CrpdcVc9MTu
J6/y/Jguk6KVGKA0Pb7eMu3fVMvy8cAKClqdOleUBBa8OdNzKIrUmP6YIj6pRDpE
+243acBa3U1InN2zfkLM0xhv7XmuXN/mbizls5f3qfo+mmS0+vYPMZN93dUGAfbK
MV3mbCLWnzfaY71aYtCA0ikX7tpE3jpfkh+2PxhSdW6cqABLwtKCQ819uG0Czx4y
+Yr/d+LjXVS7pgEzSczwB7fddohArHEks926VsfzUrRDd4uy6oUjNVrlmE5IBL27
UBPVkOjV0CpCsHFdecmGjDH9xMVer8H0ZsMpxRbq4l4d0UKLurtRgM0sH+QqHIof
2FaYert6mtKF+gZg3SUAB1xCIShTHe/QdJdNnz34P+R2l0gsGfl8NMSKnB5k7BaF
zLLSDqhj/WzYyEEyIs+62X0JBHowZN/l+tnDFc78OPPLF0NfFCNPCTjp9VRKFqIy
fmUNG6EOgSf7FZeKFAprATd1nUXF0b4njjqDmHdNjvGiJam/jLFUVd92N9ECBT2T
EUTdnHeCPgKTXKtZRUocFYe8T6UVYzfyQsc9Gu0bwj+d860Nb0nRmmjJRBObMMcY
05/VTS/OjNU752pB+W+L9KzFqbrz62LEkaE/WgutwU8Ebwr9x63UM4AswsZjI65s
mu4lsRH45LzyF0d69Ov5xJj8XhiwjY2DifODNToXDFtKXPm6gJJF7TfVCy29ECzS
cgxAVq3pr0v3Nby6IVOdZRKEa/2KCLvOJBIglRW8u4T9QPdxfL3F3njW9dKUtUsy
U+w0az/VpMEbD+JxC1wMR9TX/ZV3Q4ptmvT9w59QU77cegk47TFAnFqqiZFV4Vel
lXxBgi4eeXYNi1Hfn56/f63S+Prjpp9LutAFu9gt3ElSE8U6AGwVm4hLXL4d7hxU
GnfWXVfe8hVnlgsWxjRzfMaUKr1vRgXsPVJDc3Iu+E9U6qMSMJqTBl4Gy2gzMF2e
/fKCIXH7kzkk/B42h6WhL7BHo9EM2SVjyWi6TnmcdOMWf9Axqop0PvPvwqcl/JEz
ymHM3WEpFloikNPgpbHHGrtfm9ajwTgHN87XqhwC/QEXPTgKlINcqboO1faFEQKZ
ms4+NC8S2CLK4Gs5jkkGDM99cgVfKa+4iIQ66wmyJKq2z6qdIciOJgdMhA1dxpD5
626VCml68pvSJjGyGa6cEeA3hK8q2GzF3OYTwXjOf6IyDmM3GfL7fpwZiJteA7oC
KY71V5MOrHf92GpcUHZldvuNH8N6wMPF0xai8fVCsInszNVK1Z/hkUbcwaTgoO5O
yEEUmq2fH0XXea/4ywApXPlLEo2tYcBk+RMXGqb+LOK6s5Y3p4yDX1XYAyjMMh9f
Gv+Vr3FQZbfG5SPNgigUA+i9Xyu5SQeIh6Bt9nYa0gg+WE8oPG4MGUfjrLJqeXr3
vl/tQVsOnUZAw/0P61fs7+RnBB0Pam1indB0CWBATC9Xu3SLtEVacv1bwHDuh/nz
eMfdHXNK3/8T42tO8idoLGYarAvIdEVXKFn/fqB5KKUTj8sse0v/5MtYLRhZw+sA
BsaU55w0c3tTTImTsFk3a6VIbji3Dys2AvbL/e5wHJ0ESlkMrZYAmsGiO5HOdpbR
lEop5OTimRb2Sbiv016/2hImkHPambo8T1dfdwEseCdQSGzkSwoWkCfmP3p6hwsM
OSW/QI/L5mCnZjiglr0Gi648gkJpM2g6uWc6qgcWyTyerIg0otuJTZHiVG1nZrJr
BStQvR4k5N22g5U3Bimq5ao+zClV2oVzIALLts1GBaXMkWhmAVfGLnMhlfmEIOEW
xt32BSDAOC1K4G/vw1Gu+nM7Mzuv1HWwJr0Dya7XjYhJ5kRFaUo/wwJZ5on2Dvjb
Ds1z0oM1ZnyBwsmkqrQtMB+KGq/VgRnvh3xPlb3PDAeQ4w/YUaKHQbo+TOQL+3Cp
FonNcJzsep7Un6CafvHztJFrxtI3liL3t9URhPjhSwGYnGPx4LZzLcxHPioHttI2
ec8wrye/MLzfiMGPeIfvBw8jj00X00ftTMrc3D3Z8V5PfHkkYZZCTSlLM2ourm99
ArbBJuk0lYshgQe2YWkRXrFDBDygc2rCpt/XV6JS930wqxplKL2K5FURy+q77VLB
Gfa+bru1x5xYGCYmc3798cfWkyZ+BnmWxOkoSEryp3cadTlT0j4iobR0BUtgEtx4
7sITe1qTKi5JvzErs69/GFPnTuTDwX9+zEe2kZpksf7RhAgDpUFiH+NXMbofwRBB
iUoVsCRnPp0OsufE7c0P/Ls9mwHrj/bzPtn8Ztly7J8ffLAb3sahOr1ixKGAIine
F7nmiZD1and5tw4DFyCkeqMYsdWvImFOZ7Mm22ptkMMgGNXzGZjdlFwO3fZ2N+9S
aZFamnvab2XjGMSOTbHf64vfsvGWSPXuhteM1S38bdFq/I8qJKVTt0oVcD0x2cJO
pLWHslc5IwE0PDlfI6bqbZqg8vShOf2S7ZqJBkDijmn32zhdk8ONrZMmlVG6CTm9
M88p5VaAuH2SNaPsiK1P9d9tdMOWJyJLOI6tIn6gzLVpJtkk9d6tpAEKaLDGZg8L
dI/7yh5YVH7tqZ6Xb15oJHBHuEYD2AJo0XLstAvljKsOMronXS/2XH5oBSRxVqKf
wR5mx7DzgLdrvqis98yfgzJC7DJ2mE1yDAHT/vRRP/bWi/wE2a6BeUiOZ6J/FtRN
8ifq22qtSOwT3LuVr12KjMXPCiC7qtxCCiLN1M5pnXKsdPFqIQc/vCrwvExe+6Mb
P3ml7kAVJP8gj6eFmbXniy7YKMoYkznXJ0VagZZnmg8=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
T4uea9GeqBqE5zAx6f982OAIqcBoKvg0G7MbefqKJjNWp40tFZdjrkcgFuSdb7Oj
1OXJr+4b7FGi9TPiglrSbJYtwL9c2ERguT/BqJRHtuPiJM6tIKt8eMlS+Pcxii0A
uD3yXTR6nJy19qadRE/bWHh0S9q5WQ/z820yRUrU9JCqtjBiTzUsX241kc4p2x8D
iRaiHdQDbZnNeq09+vqB3pGqYLRI5WDWTW6OBhF+Bx5POne7lBgLwVyzxTOJy/8U
mMoSK/N/7WMRx7i3rsT/u5QOWs/CQtQmfPaQeDv8LEhmNugar3z/b+fxoFYOFluC
WlnAjIUdjMv8ytBj0GHFEg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7184 )
`pragma protect data_block
zJU3kxlzvE8EnALmY+1SSupkaw8jkBYjKzfWpagmAruDKVl5oW2Itn/2LjTtqzIa
POuG/kRLi3YT5Iy8DXmrJjsj/XH52e8eOdTWjLsJdOn25qJ6jR8vK/ONuN1gUd9V
jRAChlyb+nxJtXM3gZ1kLzGN3kiEsAQ+aOd9lM2KNsIn+/8CJaMKO+xjFqb5iC7T
KcvHdWpzWUEYWTQx71HBBMKjvQnFrRigCPkOpy7NgDKm0lYZieXwirH9HwUG+whU
rFMxBuUz9qN1HT8hUEIlmmXcYyfrFjolAT6tOyfKuGmr29JvgvyMSK1WJpxU955T
hm5zQmJxykxcoPF9DHF3MTtK1cE7QdT7rSj2NA1Lp6/co/esDOFgs2CUEe3gETls
FrM0nn6MUdztM+xKfzxjan854oiuBmBdRWnshUAMfQeySpV3RSJCow8IkSf3SHfP
SJfZqhC0opFFBXmUi63ovQCuEd4zushlgIGfM4cYKE9nq1418F/GHMHglUZuzJeA
RPpr/xTQZA2Pxzc0ZymMvjQ+ISiPg5dQQ58axRDICLRNkIvtP8LcIXiyg/VDB5/r
+uYM/yCxTkGYCjL0jts6shyNKzPQfdJMCB7AmkMpNUodip8qwjLHOtwtmr2ex09N
AwVJNSZ+vgBCYRzFBz5K/XAIzuvMCNqnKHSpmHv4uSzXsN5CRfQH/sl8MiwvJ+FI
IMhOMUJgXskE090EmVaIGGYCI/BjiXKVFJOyaYldMrl3lbHwcbNuUeZv6ixZgH9m
dr/p5KqyD+CSTw3+vKiREZGu+deJtp00rt0400bQpVHqLKb82MYarvmgyT3LviZK
nLOKO3EupkQ+TUJjqUo8RFgCRHwJHEE8t2/4CmlOGpRSq13Lp7R/rr740Lw2cO2Q
9EIViSoksH7oQFL2cgdctFf5F8LhHJQdQ+lDVcFPvskuvnPLn6Ic+jdETEmb5Qzq
6/5ZVpGUGDCLW0NNHIdyGXTH0o+vXzdGVMgW9dAZsN701FVxoYcN833yENAZfdMn
QZN4nx9t3aFN0M3HnfY3ws4Tz3g6k/HrR7TcqnTHZIz3i+uYToGz2RjkZco0OORy
Dk4xduJyfmqHcgSVqojISuIRehspM7Kow2zWz9w38+/Jd4q5xy1qw+2vUbZKLDKP
4PiNukz98ZKFrJIwYhL0AoN+FVp8EcUsqRV8gbQzEb4ZC6wqAjfs+PL/VEGLDnbH
7kU3kgX7eMD8sHkWL5R2yT+MDmjNDE9i8WUI6gL+ZNfGYxfPXwLxn7M4si5dEePe
qYR3vAXqNDWo6zwiSMuxMZMOCUe1NYtTnVMGv+CVjwXtAQw2I5OVvKbEUp2kdR8c
ZFdSe2Lt9vypXgCEfcd5I8HkFUm7Dht64O61PsXSA7w4JDkwir8/6qY9y7dFVnWW
zxBhqtpg0HivswnxqbeGJ/BUQDdTdqYa4KfgBf3iEc+Nn8pHsC1oCnc7mtMcGVx4
in+QyT4JQnADCmoOo41J6EnU3lKGjw2IHOWfd6vu0mzJiGXkZ/OIc8drcnA2xAqE
deFaLztGyks0436kojENy2mHQPw8hZ2nuN6QcjoDa60vwCbSffawjfuO2L+0tvfx
jZytGFdj6P12XOmLAZ3AGJz9DKYmyybUld22AjLCzNaEU/w2p0pMALQk9bOD3Ye2
g/NKWNhX8ed6aAd0Hp058qnOl79W0N0I+GkxpNaOCaZphYh9nFXotEoj43SEJzsA
a7JArAbYxo4z3IukuqS/7pomJMRnev1jpR4jHg4bY6slp0ILbgqNsPADYjwkKby7
Lt000orWE8zYPqZMxegn7Tb2hSqa5vZs9j3S7URXkd2J/eKAWQY+JsT7DX97nmgG
cPEdR3FhxY2vHE9ViuC3lZx0IdBFi7ofWxObB6CDPEn1wb2JmNnfSeibnzwyD9eO
Un9+TWnrXPoI74LXRmkZcCAL0FuxtoJo78oEx7uSKP2tcmQWEfpMB4v+e8CaZEpc
l+7PGG4naNwjQCaaXwgOnCAAEKP+zRumy0WjGAt4w5OH088UrPiRgDSbWps62wmd
UshmdPm7/miGzYnWbnNtCeSuST94+fwBL64D8EpikCL9x2FQcEcKMYrmOyH+gm/o
PDRppNu/0WMB3/tg1jqYqgwh2HKaxshslx7vYtgj0ApsdqEs2Y1qLXtihV9mrDCc
sTN1g0r5KJ2f1cgpuBWap6nmflg7B/keVHDZxcX2utTbQvvE2FGEJq3CkKLW/w3W
CRXJJfNmiSX/C2zcIzsLlProCBfn3NRiSgLF9ZaUSkzZs8LRrEl3cVwUVGS6LsaI
nyQSjIN9R+CYxu93htIbnVh22Yt5hNEJUfwS3CPEUdtkIL+Or16oo4Z3729NVLx0
s9wB3hVH4FfZzdsB0/Z7ZSTFHk97f12T3qCOD1kfHyrZ5ob9mya9wsjEk8g+rfwZ
np5iM9jO5mJZvwdAx1kfHZjR0lD/sQy9rTYv0Ox+/yJps0OSIwZ4wn/6/qmmrw3J
paAN4LBJ+DnQhQfcuvBjbv2E0MF/gRGWDNA5gnCOmtm3SFdAMoSspOQcgPh3Bee/
5ZLOMkUd4538nKGtdo+HQ6cJZ04m2kWlBQGwhMwaDvOV1YvswWMQlYMxbecYHksY
GlEcEyxRcqDT1yLW303+4eb4ZpwxTOtHkV/FuQ+amtAwbFcOpx6JHpX4JX/yJocv
41+Y9J0k/gqY67PUdS86LQAcEVvtecROq3KIIpGqBBBt3UmAZs5fZZdhUWrO5MQA
qRbNNzLjgHw20Wv7KorwGrslt3S7H/20KjpqFCkiksA4b6PsaB08w52Aah100tft
RcvMH2dpcLRMm/ZMLqy9w+eDO62GDE8wJCtOJ+uoS5N7IjK0+aU+pcenklJJxQYl
gWXmFzanHV56rNwzSmlldBPXYbOH+YF0KZ17MByTaTVEvRZh50da/3j/Hz+6KHry
h7aEX8ln3uTLFCmMtallvBA+JDPfGmYspD2Wb1NOVeCLW2SmMlr5+mBeVEmSC4S+
IHr/13jABKenaAV+JQKmcJfEe20j5wGdXIas+nPiFjwYULyn6LLMLylu+ITY9odb
+G5wvIBAxur441JGjHzTjP+F26dLSrUh8GkYugSU8Lq8kgZdYjOcPiGVlAa/ihtT
rMeO3Wb5XSK27ZnosTeS0YQNr6ky1NLsxPT4OvU5MHkOoLuYAN2vnqExb3U2/844
fuoFtrzN80BezEvNXZlZl0ECiEvd3uxaOKOdSOVAW7zueL5jcFfiAoeBb2hWfWRK
VPkFzxUrmVWRAtZRJLDYtGwgZNAeZ/WZBFpuqncG+IVgNaUlYL4we1brzoxndK70
RLsD0KEXrwuPfxo2Juno/vzfpQM5hARA5cWaZ/UCsXXXCM696zpjcOD4M6E/nalP
N7i+hRq7VsfVHlgZ9eA7bqKwru/5yJDW4l1tUr7rxHkXmzoCIaov4F2cqfFgNUsS
8MNrw2GKwDcmS4CoAjQSATnAtEgJvzdMqawIqQOVcgszLrwTjJ85CNEiE11Z6eXs
IXspxpJLtv0CSbS+nPIdFGoeZvjEvrd2SuLrzOyICaFCIvndVBANbIqxfT+YndW2
ChndDHHPExabiXfzRdzK6fxgg/7xvLwMcR0L3t7VsW9VnVALgFPgQdWIobjG2d3Z
yidxl7uSg2MB/CNRHjKSmBe8MDpFteS82K36LVkHApbW7JxldTcZxCZ9e0vBuTyx
duTXx4YDil8j8j+218d46iyRSMr1lUu34wyZoOIOLfiyyXxY8JDPJ7To4QNg3nH1
oY0eKlgPHwerIgdAs6ChYZGKfx0UR5/LUk91Bk2SahVPdxVXzQW87U7DikYhtZqP
l8ZukabjMx1qLTPz9GE9uVQBeiYhN/PAwzkprAJyGavQZvE8qZeGKH7ybesCwNvA
Mt9pK5svbFAhUmzEKTNuDmLM3ae/+1nMWtjvOoijK2ZferYxs4xTPVeP1uJ8sIiZ
dDCN9duxoiMrZO0CU5J7/etwqyd+Th+jqUn7GhvvkeKAmFxAzCbPfOns5UGX20yv
wReHMdg4nUfV+g0eb0+wMn/u7PDcaak/QMaNylzaZ2Xa4Y9rZy+/qX1LmVoLP0jv
yXahsbBMRKrECXVMNhOKY3R4OoyjSoRUPdpnF+/iyiu3kQv7hkbBenppFEJtQDV8
Lh7g1ATrfK8OUu58EVcwFvoNvmMdgBdLyL/l4FQfHrRQoYaLQ5HYnEJNNalysa6M
jJvjzZlYPigtCwlwj3r9l3zpHTb2VrWVzUuNDEBGaQCHe9LSEpbMcjtcQ4tTzbXu
hTawd6tcn8kUO7BWYGaAqX300xjy5zysRQlt3ffp5H/rQdQFQk2trpc7oZeauryW
N/nH2mh1r0RXpZiJhTQ+yTpsUqoPNt4QjBwo/tEvdrjmshWsNEFV0fKPyLaTKJT7
atdWUhcRT8zC4qpLLEQGumnW3CZ3pxSJ/2VoLzA43IF0kYPxq1fd6ACEppUQfzOc
tSzO9RGDyF+slczjOhuLLaaiG7HVfE/byDrUKAQyxtbld5fw1hjbQyxi7xKX9OR3
mKOjYQuwTGgBk9pBA834ABWTfdvXiFqd6OqWstpgcS9aC48+JxJxus0FouUAgUdD
M8ZNHh99ZlB8/MzPPrcBFQEi8+ZAsaf2gp1RKO/X1aVXv1PWSHUNLtmbdKxZRYgW
FEl2CpODYMPxJul1AeXu51drPHBy28FXFSkUC68pugdm4Daieq7jSDQr661KbKk6
3M3+34sJv2KWBJqacS3+e6BTdlfNnJ6ar3v+kKyyBQ28J9PAlVrtCaTkPmm7FEYG
l/zchrd4yD9RwnDwHtL0QjlDUcCSjIMOYPREQAaTU6CzbvHBpniV8ZGooF/3OYzV
+Ca2G+ssjb1ArErc5Bt1SunHd26nNy7sFwx6qJmzy5gWTBd5YVAn12giIfvtBJrM
GWeKtbaIb1UW1NrHOTVk8R96RuKzPKRsWDCYmmzy65SoaX6dNZhhgeuASdr9k3SX
5H0h2uBycGBxV0egOiv1Q1DH8/O6hlmLUZvvM7ZnEeUQ9pbAal61RyKrjKXILz/7
5WtmEbP2cD219fFwzt1s7XvlpkWHPlFuFdE1QkMgyBffCZ8gvPUle3Hsa0C420FP
+42OzBuOeCrLiawYcewyaEs1THNF0BeKN3/pNTIu3gHai/cQpCHsyQQ7C0rLFEPi
cByOgKbbCaEh2W79p+BKcVrEeZwbYaBj3EJCIrMsP4kHNbd4tnDik4+ZGxPdUzhR
LXgYHuzMO/0QBMktzuZR1aSnne+yFt7XLcQBiz0GS2UWkXzWq6su5uvUGnWnQ/gz
J5HzsfZzdcRiA3/9ChKbOinLCx+WoP1MKZbpfBUTgT+PU6OWW89P1sdiucgfBeKj
q9Xa2nHz6ALAAG7Kiqv5/6NP1n6WgO8QhqGE8spW/rtaDqJcTwqEfyzXpCSN9f5/
9b6nSnIgx8rLzwbo0/NHF0wjwScKN3eJf1lG+d6y8SWju2OTSSvW4Yi/tJXsj4Bz
Fwwp7QqLg3CG94ATwDdPXkn1rztk0dBV9JNT/La2fuq9NxrwmxfygatvjJ3RvDyz
m78ivJzhamvQc9p31uGK8f18/8ife47AJS7oflVkumRi7LcmQUAHDzitkZX9ofZE
tKS85ASOHOHQyn0IgVRXw06LXHeR2Wt1ogAi1KFbJ/xd2vNQjqYKJyE/QeOb70K8
jiFN0xlm9QtHDb3wG3Ywd3SXKIyQ5dqYTPeA5mIP9FSN9l0WDIW5u2viAXBuJWsE
YPyTfmU9yOs0pHnrDS5O9P+2x1W7GubzFSVRF2a4c+gY1HDGAh32hoADzWb+zc2K
ISGbIkoOMuoEqsvFTSa9a2B3PKHWtCniA9kO4eGOMAusLJ701RVBicvTgvFVN9tP
vo3MEy6o3AtIn1CLUSirlcmxkH1oXfeJK51GRkewl4koBcfEWQeq7RBOdS1qpslz
40aDM7vKPdVUjP78sWYbllvIr/VxyNVsIHDyTQlY1PX7033WLmMvqn+jppNT3Aec
X/D51a2BUabhUwokUNQfNqAPEPIRue8/cH1FcK+3UQHqM+eTW8ftkMSXTKngl5Xw
Gz7aB+Mw39EFnBWeXhtQd7kJ4/g7fMFBZu+ysmCYQe2Q4P7uiwDARKm+Zy52yayD
5Yz8W3JBjeyy1OtZCXp/V0wOSMwgI+60a9RAldbft/ogGH8ROw5JuzbDStRyHfZM
zed014SnUVvL3OVcum2xxvMvienkjl4ZcJmOd9jZFlwBn77isXx/Bqd7Uoj5fVyR
02WvEN6jnjvr4UWA6Fu9jS4MfeQ1Woft2TReqHvwsUvLnridB7ZHL2MpXhRQ+iYd
GKMcCrqLPdOBiaF9JhTfQR4SoDHmszeemSnrjiv4fVxA0QNHvT4vpEthonwswQqA
cp4IQKHxrLx7yxH+jDgMq8Rs53cGL+ri7uBoHP/InUxJKvP5m2/bq9Foz0gVJbiP
TtZ2JOvdpSzkTUe2ftz74sc9ukiBabLwgT48FGcARWAsJ+PfSTwK05AFB9+sLyJb
nDjySKbeAOqCv02fORVV5dr+sVUAacaUcUHAmwm2Nt6OGsKaGl+S0c2I7RhnzAKE
dKi2Eao7zqQz/YHUQKDm4fiHJr6UW6C9jO2rzgm2XiH0MHfWdhXudE65fLRah4Cd
dj6amQ3gVhqu5mZVSiDd9VcdLTfYD+E5k5E90/m0yXUjJdGIfDzqJjZV3Yh7C0Mm
GqYo6aFcs45kX15HUjTxK3iYOwIltjKRIWQdi6JzJUSv8E+wye1mP0T0uzdMPowA
PaEepKvJF/uay9UXufeJLbH6i97rhy+5LtRZMweIECo/6tbkzWETxlN9QHaC9uBN
hMFQwqYiLGBxI3CxoRkvUhYHijDeNtA28wxW6fuHBa27/0ugnj9arHVmiMgwrBE7
UOXzreeBUJj4t0mvf1zen29AaKClpodGhHr70F3Vp2PIbwuNfhvJDT08uoTGp4aW
22m8pau2Ig+vyTTrBpB85rPUI75AxDXOeY4lTwJLiGPJWKb8jE8gCEpwsJp8J7CX
HmmDh7RcjoyY//p8du5ZvqrivLlYrtjKSeu/eRl7bhOzfDkg+fc81pGYVmf2x26Z
vyVwpYNkl0jLyw30tx/blF9tAB4BD8vIDh8l7uFVOL7YjpOzxOWEKVbjQMyUA5oT
MPoc33n/U//FNxLw5WAXhC65DcjX6Dt1snTtMzvfRatkGzmi2tbWcn17urLooNnX
cTUfhcyUSOB28nQcW3PXab/rZRumodTGOST9TdkR5TAdRfENa8AnUxlrTvVhvlei
KdD2Fs6T9LD/wvgNgmwe5X+2SbAY757oZ+YZ/+sXDumxKYGBWlfMIro2l0copghG
XNdbZOF6bQj19rOUnLYz6J3jbJ1tE4DYMrts+bmX803Y/aR44KG3mtxSpCNnbHCf
fJtB8hIUaFdsAZf+F9O+5LQYNxkmeGBIriu1WZIjqclwFsoPnOQMZ8UTwWgKWaO5
mAWXmqge0feU+RRfYALl6BHT014jLZYRg0uHC7N37n/okzSngfctbg5UqTyYSpn1
J1X2NIJhi6KvV8AhjCzthhsAnilrbOaoMGsFaU3RJ83s2cK130l51Rq6CHfo1usR
S3FcvodXLM2RNTLNqauhhwxocym8Q/CDix5+xrie5Cgpwjv+VA6OQQD5/StcW9xT
wu/YXxpNw2mnQ/x7abdpVVnrOWPNQjMCc49zdRmgh9F2tIbqf0cpadN2eeT+MsDs
UTQLOaU0FWnOpMWtMevbHoLA6jF376jClcbPA30hcHMHfEGMzr5mFcMt+mQkK+u+
H5qQejoi4mMriHWTUYagsoRGjuh7Zj6H0MqV2yODNEIBOedVv/NtXyPSjzPPnpQ1
sQbknSnOgKnwoNnck48vdxs5Rp9LNTfYf9pnpTes66ykra3x/frVhZd4/TdClT0N
jI8QhbBHnhfjNR0J+BO5wQV/PCYP1ebsZIPQoTQ/4oiUFtXkiCgVBsttJ7CgSUmJ
1Cf+DwyRsVcd3i2ETxUwyI9e2aTvRCz2Zb5NZci9u/u26c3kHLN4U1iNKnPd6eap
5byHXTtaC7p/6WebqEo75MQeH1F8XHVIGGglCpuKF/yP20RRrsrsT8rB/fOy1U3t
RAHIKYBSIozslLsvSybe5HGbp7+Z8DVIroncPNdQX7rDWB+JOV+5YjuzO9c9IQWj
O1y1q99cCsYkYyMp2RGqqSUPoRMOJZ1+GF730ZXbYZ06sPhEFUbsxWfH1894Hdk1
eY64Ve9ZQA8aUWqmlSwj4cVMZykDWwfFZfiLDZ0+Qilitpn6424XlxhSB2CdQXyH
KOQ6TtPngcarJtLkqX56A1Po8SiXT30gjSNTJNC9HSU1ir8wfYyrxhz1xFxX9wgD
8QO2iTUBVkh+XuRW9Y6RrHxZr38W8p4qNT5So1dR97IOdJXfDOuBuV0+EPzLQz+f
xgnEFStFrer5d3b5nBxVfCelfDJFx0kVz/TGOzHj4HOl89af6oki5WWPVw1bncsB
RZ0yxuaW0tpQ6SScuN01RemZVK9gSVP6rdRnbIir/iWp+12freBmr1ubYZGZ7Sja
WBxTgoNoN6v7cpdh9YCOXM2849WxMrkL2K5gcP5pqRKvvmzdQDdPe4H8e1DhP/Nk
iXm4L1/1TPPSvekX+jbKalwZ03MwJFoZmGjcrpM1ejMAHqjxFG8oR5FBV7ZHptAe
ohiCRIZbpDxMkv/c80AkUhjIy3y8tKreyjUAd1ZRKiBI2+jyXqAdmGQ9NEWhNQ/5
bZye/tUQSf7gGoRpFAOjfb7ORap57xBtGbOCojxKo+eV8uMU0U7CGkyPZo2uVDdl
Pgxxb9ZM3WO7cmNJyjusWpALln2ClJkzU0Z/qsUpZl9w5IHqUVXGkn86JQFS8x4Y
jKCR8nEhQWFiwt6XOn6UUF4lTMHK4WjBM02F+C0Bs/t1b1qIh7gR0F0szxJPtHz8
YHmVTGqtYRYcr6/2Ylf/cmKSbwCJ5DVuT09mSCwLyhotA7ur+wThwLs0GqeFrfYm
DFXRPo7IxJUMzQWX1jCn/MQV3PfJbggLGGPgKZJKOftDIU8VzM2maaJBMbYAEf74
7GBGY/vehP+5eDFhfXE9gCs24HxH5KUnL2hIHhJfo0ebcOHKUTP+LJ0KqL5SVYPg
rPtuvx6Yp8cXFNqFrNUDqghuv3NtsMVb3bjPRhYZzGCpaFs/ueKU0NsEyzRDX8VD
/OE36UmfIsAKGMMP/ZsHJZOjh8+bdHEY/Nh+AQJA0RWe0BpX+gd3XMImGXMeINuA
sWcWHdvdn3F0lqCE9omGdD4yFWgrbGHVTemIe6407U1RZXpI3r1lH1fO88LE/1jF
VfcBtbYnna+vy/l0Caz7SM1+Z+oclYGiDhI0i17Bowv1XlSx20qqAkaxxN34cHx3
wIqvMA24Zxzd9VHG+tQKhbRztA9cix5Ybit3d1hIk/XQ7ie4CceUELvYLMSb9NhN
YGEh9h7V5MCvMVaNQC/mlAGc721gUCDHBtVHk3hML+YKiq4jPWxiNMPoA7mINYXS
gBMGRFUXuVIL51i0aGm/lGZYeI5smbZ5Y5NwHgmQ6+U=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Ora39Sd80IDNrQeN9rCdLiDvYVbXVu2B4qK2jOR+0LvkcsMDr6VBgeTpGyp1VZzM
MND0skzRGh1Z9Bfma4cTiahFTaLJgVT2TOKEVFla8R9uOGMKcOyh3QFbS8obHYzA
8mqp3i03rM7EM8xD5bB7Rs8K49Lfc4o0sg7J7tv9lwAdhrgVhCo2FvQFSRvRbIuJ
BYp9oQn0w/309irz4PMFHwM6u0+TaQY3EGTYxUvrL6ofGPCbBaDOsRxsV39ZWEfM
c0d8JOgfR9TqJ4H8g8Tm4Ck9OEInYrqeN9eolRhlAzv1vt/sLNO3gN7F/TEWnYzF
twdHLj1DDDuKCtsqfRPnRg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 21744 )
`pragma protect data_block
49pf/aQ1GxF6wTbRc1XwyK5sBSQBn9f0PNCrkHLal7jf/z8Z2XQs0yDAWkxXb2Zz
+S2AvmP/aYSSF/7r0IupgEpWqZ5fiG6WXR1ozD4nmGLlUi/DWHZ90kkC866e8BJ7
3DD/yu3PdU/aBFVFaozFvCUBZB/copyG7wHCLfF14rnipeXuHR18u76LSGOqnqXU
F7bfGVxyqFqw/Rv8Unv3NgGOwb9nNRAZjVZY3GQZqf2WJOz2PCoop7qGiLqi91SL
0Na+w54ytfwhCNF7jpn+c1xeIHBSnmuAKMFOvNK+DYl6kzdGgNyHeCca+pidn7Q0
nixDG3JLXCAHX99/8US3KKdvMOlB5R3KYpUiZorHK27nFo2Y/dYIrpfSFnal+4Vy
ZC0xuRUa5wsIkqRsZ9OawQevjHv6cA3HsaOd7/EDU52nCJpM7BibseRCqZp0BmuV
NkbqTY1xmcCjoo9bcjZNMnVlqWE8JNCThkxhtIySuvaKU3ynH/jF0QBTbyJKVUse
Bx6CLzevWvB8vQLNUKKZeec8CfYKh0XudYIOxJl/KiEUvdDvQ8zkJmL4cifpNJwN
Kjlo8grkbSrw1pp4+qJ8YDI8SJIdWzUVmwDaTr2cIcx3cFXFxbR/GdTBmlONRH/J
FY4OeYd8GMQzL8395h2hg6ECuzoADd4tVdHsgS9lzy7QkBvuMcroDFbmkKCs3aTt
6tt3/MhuhgZf19Sd8rWvaIg46wR8mkFuOZPN3XlTO0E4kBv0ifWKeOHjY8qKmp0g
/yyYR7rMlOyLkY7Lq+lWLzHkCCHTM6aWojISCawYEnLyWLUQw0Hi0m4+olDjIxli
r/K6jLg+AgmSWekge2LvBpcc66Vu9qzUSAhcNn8BicQF+znkTdELFZ+JRzlOnLs4
frB19+C6i2DlHqW9YYXTjPDb2nILzSg1/MjX1sRYv7CM8bTMQZMd0X4V93Sz2gj4
rSiJS8iytaa0Mlj8sTwLMKQq9waegsMXyqJcP5c4oRJveP5bpReU/aN2z1g2xntl
fxiqmGDpEaDkSs6LQMNbMnNxWESMkBuedqEWFuBzm7q/sfMwq6SjOlK07jGJEIxJ
/SG+3pe2EEAz+ej5zi3AL0ibAG+BJmg0WJ7bG/Lb1PYFCBRt3yJBfi/pqJJKzdRl
fLan9O74fjX0FILhAP3/b1OG3pfEuz8KyWr9QnE2BnXgkplYmlWZ+wLEJSndEi8X
MaIUo+fTvk9DOahE0fUaB5VEI/6JKGi8tJUrRI9YRNjP76A9eeQO0nf5PUTIc74P
j6lP47pzfQJFntCCQzF256iVEprdwSarz0GUrWMxHu/CHAqrOm/srtSsSGm+N0CX
gGMhHW5wfpXBL92auPm7MHI0dIcg2KA2viWhAS0SuI0FJWSG5qCOTj1jDDQgggqm
jDZChYLLFl/6XWu1W3L+Xx/+hV3AubhC9y20Al6XmhCT+q0J6BKPkIwebQg24F9H
3cAtZSdg6BN0DQeTHMFWZSfdT00prJk0A8Zo8+zDKnMDIsG72kjC3aCwZBmeQZKr
wSRiEhbcJPACraWkkBGHbWFM903RaXuvZEYcjzoq7LjPRMG/mLz8mpa5AkrfQG/G
QP2NKGgU6UYjb0E1ZzIgh8UeuUM4Ve/NDUfr3NVb4A/MYv1Tu/l7YSmyqeh4q7LH
ZS2Vxz/4nixEFIWpfLtmxPvv1xuONDVS4r9EYaf6dG0XzlWySrKuDYKP/77LGbD7
biBGTChDMpAtYybw1L08xdmgqFYrx88d4nIzDZSVByXkXPbzrwr1J9v+kHRW5S3S
suT4t0akoV3Yg4XaUTSSJSX99jTHQdPgQfVs2V53SJ9joydiCYPEnH/HBbFPEzu3
jJCnIJOH+gtpgfQyoi7i0dujrnK8Ov+I7X7PkNO+YnBdHjAY96aAli/hNXZ07qJr
CWJUuwYhnU0mtd/+TcUPaM/Z/y9oClk98pI7oBonl0cvTUtI58+ja5PaLHp/UCJH
etXxr5N2hF3veYVPngkntGX2fX4/k7udvGxmmNe7qNU2HDl9ENvEK5HpYnYVs+kM
gvowqsQj1Lj124FEjmHC3aYkcA0f4h/LEOG92nPzHK98CP4FpWxPyDVIHjqxN0Eg
OCb344uDkb7Ka34rloQRPEuEYaw/Na5YFN6u70S22yTjA1HV35q++qYuWCiVQ7Hw
w2J1fKaL46sGsKPgLcDFjYv3gtsIwjsTQTDBmRCW/VYOsB7lXNOWbuVuWraGw2Uk
U8TAt8OgQNRr5Pa/dqSupWhsXPMZ0SCYHFD6PA2aPCsd2sUESQ0eCTK0JqKnp3YQ
RfwdD3a/QCPfPJaVo6bF91stafMtNZ1cGpIfpWopZKCAFqmHs2N61QB0tobSCrNY
S//OP5xvk/hfRVLOI3a9u72Fi9yiVwbBhObfwUkuk7U2J/Y4alITuP68cyF/g/5h
g0ViGYe0/FCI3WKYSpWiFppoqm+XFqfbBhZOGPAVv4EKmfr6efoy9N0uw2ER3Lik
RgXMUcpTdirzA/RW8exW0hh4zGqrlo8+B5CZBE45PEoQq7HG1xJr5eLA35N4j9JR
TEroSehF1hvvlA0WAZ+qgJKuu/L62XLV+H/RSe4DijkKBfH/xmPiFVW9T6UHILPk
1A7gk5ahldyr6ez709h/0qgnMB/B/bwqIsph64fLP5mNdNHBlD1yGtp6SouakPd3
T2anLfYXSCFTrIqdp7xEFaoMhPvzPHYyD1S6r8TvarJizxwuFVYShdAG5nR2LvIM
xpeX/DuJGqFp25GIXodLnjuKzkrt+McppOExkB62mi4h27QJ8YViPRCWvUYQzkRF
5v4nUGidSQR492iD/T+2j02aeAyMCPLwJ4lpHVxA4bUijgDaMKFX/wW1BUNOTiQH
IFI8PQ3rvXdWxwrRKBg/g2Z34HoP7XS5JixA+7DNO2NK1mETwBTIllvqGl9mfQiS
nfuupA5l+wy2UUYASnIKqNzR5W/YhWeNLsii5KWgOipS08lWQA3rC/6z/D1jLoJe
xgDG1wpE+11bi17ckubMAllGYqIKW6fOAPj+Vnrb6QLfGioR5FTj7m4BoGE1UpHO
U80dsujSV8ORUUnDSjuCs60rbF4VvqRdKk3Dk24zznvQ0khtWARg283+PNQVxgCx
5LfElFueDpAKI/6u5UtvOa4aFDcfucvRqahDY3fZmpTRfagKykLrB9pyyuOCoJi0
+uQ71u9D2/vwKsb+/N3E+wY4w9L26pM0+5ZKxX3EkN/Y2QZ/RVydVTvmN6JLh1S1
yKqGMKhBXjl0s7zMPYArU2NFfJ9fSfbiGV80vniUKEZOibupsz02bzAP8ZTFiF3p
ZmjHwB88gnGanCyXREAw4H89JkWBvHWMQqQvBY7Q+fexuc8palu3hPwGEFO56dyG
RnEzzZi7UBdE3uZxSnPuDoEfhP/ng9Kz7/QqJsVV0LFngrlBkh1FOUuIVmsFZSna
rAR0ywZGTBxhfuSb3QsJsVvLv6yXSxySIjHuqcUcSFC0m/NJWj20pgRfM+nY759h
soCKyJRlGKhHtLLdFODl0blHEHA3+NVhXVGsfSeFTCdMLHZtqrtx1UpERGuXuuH8
Ctf3b+9RcTiOnklytDdzytnox98nLUjzp/16yczWshifm/v1eP5vDuYryrYy6und
sHVFjFN5f9juW0UuMOEpGLmznZ8JF+7omJY+3y9FrFaFl46fv69eoNmHSEYXCu57
bsYsXD2cXzKA5swCRLcRrvF1D3cKD6IxGEFDzSxSoLBkymIRR21AXorisraTb423
SPZCSHpOYrNw4OfBsp2ysFit96CubSLXZzNeakg9McAoetd7DWT/wnyPHBIcAcNa
jFyOqrndOzQCFcMyteHqJpz4kLaRnJG2v0FHfe/u2Gv5WShxbrKiO41hx5+sFfw1
rcPQF6Q0nPNIUY3rAxaib/5AtccoQu3tyzqjE/iqkq1xfVDb12yn7+5l/7jbS7cn
EwbAFDHpcQkYfrWUIHdESvYAxdqGlJtOnABxP3bvj5gC+Nm8WY3Acct4IEf0g1C5
ugeIqj8hmZHKulAuCml46MBjJooaAO0iqVTpdHMJLaErmOhHc8kL76dSJ/BL527a
3JVN5Tf3lW3b9MZJ+ZygYcgozzZQZxtfG58XdWhmf7zNmiBG6B4PMAI3QZlEUAoX
9g9bwxtKCqN5xPMwNiKHClFQS3mw+bZBmAr7B7loe8EIg19IY+wQMm36dwsiL2hI
UVq14FIPBSbR3YJdL1rCnI8fEJ875vzi2qRfMyzl/qibmymwNaCHq7EZj6BrTnen
Uqd58hiLQB2QCO6ogtnBW7tyrq6TO4ZVEiVDXlkNbn0mWpM+3O9nIKp5oEBKEF9M
FH58iSjvzoFhlTGSUOSCfWqZUfQLjurT4za1Z5lwqJYznK8FXHZWpGk+khylxcS9
vEE0QpsyHYp3CYE3Jo+VPtwEp8BcoNrGLbnHyHk7Gmjvsq6QjoffVTat1jpUxpNI
X3dfE7b/rFFyCfs6/49RelWDMYXjDGFrvGUckUZM5pz47pzY/oeU3BaiKV5xEIp8
w6pWwNzsyCaCl88I9t2t6V9UpNDU/ONQIN7HjNm2Upze/gRue8FdLqHgy24fnu7U
r3F8/4VI14i4wTcdDjlp+LcEQKqfbYd+lrY4xeMi31YoDawD/gr/1unZY2TJJUdp
ah/eL5nluev3kIksdlyAPi/QcWPpP0T+94khzPNDGW+H6bgsZEpSGu/6xRFyMLOt
yPdaERA8NAxxBwE87tyLClXzPm0WT8hLw1B/keZFt37JFiDcy96UjSk4z1qsHX3v
4cc7DCp2ZEx7y9ZWahzwgagvcmQgjYUWh6OJ+hx9XCoZQcsq0J6O94Eln7t37spy
Q9f0hKfH+WwwD+zWLonP8DZzD1trgl39h2i0fCcEfJgtP+/ojiz3MfT8BMPY/d+l
W07cFb2akaZrzwDGH33Xfiw8TxvU9RbptftDMQNaLflgMto2POWKWDJKgSub5eJB
oTHLCqyCbaT0rYbnQtzK2uSiXPnZqAjeRgS1ZkT0R75b9ltDNJSDp4AGSEWTmqUW
5i+VDXVHyh5YGh2GRc2BGzOzqDmyGOm9LjeEuvEbZYKDXlSA737iXkVPYfOJumwR
vsYHYqLZTEl6e+EyEMfSsj16INSzWdzHI5uyg6eV5YBr/jcKL0EqLYHy+IN6bDn8
M+RinzrhlnI+pFLjf4ISVtCbbFTZ8uuXEY5PpmKkJwHS/22POYLKLLWhf+Muuo4C
9YugVrFm2Nm1DThQyUAmMPs4P/kiyaGYnO/1HpIoyQQlX6QclAJJMO9To/9IK0ae
S4XkPEe77B5wIaumo1uQS/YqkhAs4bzhzPFp4bA8unREqFJflycnd2I6OXK3MkMV
P2rAenWXXJ1LK4HfbB2Pzoc/csvyijqlUeOdLC7YqW1r5l5xcumC5H3Qwot2V4eG
UJhxmYMnPnZvjaaPrrRaHDyd2fcrHeUdYMURpgc50zcpoN0t5ef3huuu+5DPHE75
wz5JciQ8fJfVHomGdHKnvt5p3i9pG8zMv7QTxp43kc1PRWNnB232HzkOnpeVJGUj
cjc114/qZbtIXuQbopvwyZChGjn1ACuAcuFoZo/r+TeqbUblPHoj0noPRynJqfn1
bhEQbMbInRA+mcnMugPNl9FaAwXMf5q+fQ01p+zk9KI8OhGu4VlcaFPRoxxLRlYx
DlYPw0rrmueYrb5Lfp2kPUVqzKpGwx3Pqv9Skj9qk8peo2+1BZZ/8E3haKy56uZe
wqGTjl1YQgO+Fu1dDpqp8zyHejBEuLQk8QfeHjGrsKMxZJWlrVx9IRvsRuIhUePs
jAFZFpwDtq0zCKjTOm4dXbr+jm2WtHx+VY9lSO6EoINrCC0AvQ4wdRHGNud8N0tK
AIpBFeelVt2cUC70PmGa/2xIq0QFOwv9a0l7KnoEYlgat5UM03dUz9vy/CweYhhR
FFJ6RzqdI9oBFTOsWHx8179lf/0SlgsJymOZ2rYkWc1MisyZ8YK+LpS+E4x997Z3
xHXm/wXcEjk5nE/gsCc+EKAap3i613JC+6c7VbRNMEiwF2FUh5rmOsxwFnQ3Tdgr
Z/361+vodHRO8l0c6Fuipe23ME0d65r1sXCertEoPKQ88atllmvH7ty7y55rC33f
2WBHByWNQrENBKyq4cSk0XjNnVvUAOeDEuMdI9N2Aho0WWdGkVuAiGatFiJnUi3m
0IltWlPcir2jb2irBqvsS8F0paTeOCayARcDNQW6pWAxbMwTMAdncC3Z3pPN1Kxv
PttwzrxBj87K1tF3p4CjcNPhooU8u8VG64cg0Hi4ikMgXVSvQnSXTLpG/jAaY24J
setHewcbYJWQz2Old2YhGO3lo1Pa7dwm9eH2LTlrpB35tEvifQJ7buK/r4t5h2yy
KR3ewSJB63jT/zhmU8eN46wTpQRFEDcyyCtqQ/f5WUXknRhtzENxM0gGCU6YDcRy
3erRBj7hhJ0FVQbh3zGtW0bLYCBOlDYZx4/wzszHy3Jp55eO+R0KxVktSJ5eHZt5
9CV9+U9nNo4x7j9TO6SCkxXHbkpNpKvOQPEX2koNWkbdKM+ALyWVoBymHBzX9xII
xjvxL5zy0vbpHDhcbaCLUaN+eirWlENxSdk51dWGXePITlF5IGU5Lxd9ns0z45PB
vNsomuijnrN7GnF1dcb3VVMUKgGzdkUpfVzwxpMLCE6NuZBO5egPGl3+Fhd/WKCw
AYUUgqXqYw8vBAUOq0NTgT5O2a3VCtXJ4x/jdlD57J4codID3rYwyDCf1WAY3qkQ
bi80PCLjOhaNdUA3MMoFAM2lUg1m2RznmpqK48MOYIya0uXPItMWeDTP/gbW0yz3
1Sdu9nMs5FeT3refs4Xg/mXBMT5N01Q2xV2iV+P8iZPigAlDjdVivMoaouclWdDy
SdZlzl5ljwZ5YBCHPwCeKyf2VQMwf2i3q2Q2QtaNm37mBq+bbzHvlLMSaIkPsN2H
u9qhRqWoapXZR4xS+LkhXu+jAQuHTJhrsCWoU3HQKL137osH4K7scPNNwZgnGj80
YV9V/WuoD0DZYHfg9f4umIXhFd4lDv/0XhMRE2hPF3/cNJNFgwDGt4z5AZ0JdKJj
3R6aB5hpF0TvVEZLZ35rBeM6UJmb0IA09HzBIOERFi8nFVFyqFi6JFLPTa8IXk3C
98RBZrt+s3+jh61Upf4RYJyZlFXKsSJfTvDgdeCEAO4OG8WpjjIxVQMlWniW2ROX
7kHSEBYAMK10u/X6jywLuS1ft8grFMF2h/zLIhUTIFZOPOBjoNUOmwQsvvO0FshD
eMJBzdPGv8tujldxTf+ttAHYaUyy3lCZSETfEMCWg11+2DQN4hDHm+Gf+mhEOGHg
5DUHN1lZUu3dyvA8XTpcfTG/afEsH6aJuLKm2Mu/J7Pws7PYvD5rWJHYdHg4Nj3u
3mCYFFwg79gji5ijhTCodoFsGeVmBhj/P9Qettm5iVfQWdDd3w5An/2vBDyWxMBy
4J6a3DbZ79NMAnEag05mpjwU5Xe4Dlh105/LBhDG8AE+Zwm80NWtZn4C8gz/j1wC
j18K4caGxGYZ6oa0kBKwRR4p44OZIExmnt86HVag5wBGraoIevDdBwlDsMW2wWzu
AYOd4+ZwQ45clmI80dqkA9upW22e+lYxw2Cp26HasUX9Gg1rrIHxu7bYPZlLYbBO
oNJAJjYFaQvaiMCCG46UfWZ0ze3mPvJe1ELUVYdIk9Cl/jn/mpOGUMMNsMUSyaNO
fv42ijmo9aO3XKTUYSpHt/mMBdGssOJJWK+EhtxWGKhcSCjPAt98PgKKNrI53i/v
yFIKqhEU0d50cLooR7XBvPIuFcvd6uTaH0wnoyiphC1F4RVuKTEQtwuY3n6ACb58
uFyntaR7dim3zq2UKE+uKOa/rgTmHn0K7z8zoQJmIwg8aQI6GG0Jm3LZP8i+ZzXH
JMl6zedaBFrJ2HzWbrxYFtiU+bwOqCfvVJZzT1nv2Rh7OmtFkR80eRhPlexvLMKe
OUHaNCi4LYhEdRcDAu4p9WI2Bp6Qfyv2XF/EmJqTGDi4N4OrgoKRYBKeC9zMYmSf
unWVhK6pD7Nx40bTVEl9783DQnBPzQ5z0H1j9ktGtLt36lq25R5FVEafjh/8e5kH
OGLqG0oWKeYCwKUBDJ1tQYaXc2yPuqkrFKKqUifPFgJXq/FaDnIVPMbvihbNVjrs
hmFeqEFrbCe4PuI7c2mqhtT6TWukzfyhQElQV73xDXdADy75CN7e/B1h7nIWTQ8Z
8bg2jdIAcUmgoaHuRDCsOuOQCoU6+ikcmqoZYjJqU4TSG1x+SQwHiKH/ei3eDmav
Kpy3/DBreWkrDzmccG57k+j+KWAcuT5DKHPlyN3wGRZYOnOI6nzB4MEDckquA5IW
ECQzwwRJLmuEjiIEYzyoEYbHFeZhEp5R/tAurOUdRC6NTdZxM9sPZ4dEA3R9GaJb
OAzx6Yu8e1WFeOoeYr69gemQJefWDNYTGJrNxDlfSi3SXxsalLPiCkMBBo6ATkqE
A1Fi3oxFqN+a2uL4uWET46iUAYHQmhApl6rf/6N6hIC1Mg4hQHp9xeJW7Lf9jt+u
gTpbqnpK8a8jI3QYeWCeQiJr0b6QldHOxlfXsbqpWplljY1UgcgCr4XBdAccriuq
c5HFV6HudIGLWiMfaSDLQI8MB7CJuYxP2B+Sjazt1eGJ5wroyPvdlkdwJQueC2/j
KbGPra1juY+Zq5sXh8etVBBXBpD1UExRxxxUa4LfNCK1vat1x599BjqeTYqXusFL
APENv7BDgFhh36gXqFqYnprsxavhUkEaLdQiNGqPtuljcRi+x15EsNSnSmFQXqwP
3OqMeH2fgB2wjFSCgLji6ahJ/+H0zy2wyQighSYLKd0lHImQy22sBpwrQVUv2hp0
BNaEqfQR8KRSVQK8ZtIfBSQlHZ7CfSBPT+DcUTpJhXvQ/W8i/CCE19/xNWJqbLEq
r86LoK0eV2hEe0OjStbornM3Oaeg8992k9ZPnXgP1oL+RGmbDCa+MonJRuVpXK1q
B3YccND/4Qdsyr3q0qorcGduV5+J/SNOGphrZXqflQw8NNhMe8404eJ6nGZczP1H
n+mrc0UI0Sv59mT4szR7X1bFLNGIIlW/0kqVUqdw/4/DWlYAi+jkXhF2Sygacs27
8BkYAFuiIVkbIJJGG4CVNU80AheZdx78dPpESG/cb4CBqtHSgExluepznabhsVXW
43FShAeWFXPfI2tSPTJcutRloEZpOoELRbbOsTPKdz3fFbDr/M0t3whDT1Ajs8qX
JSihUgMZk/xs6w/awpW10KR9L3w77OElWZq8Il3Voy7q8e3a3PjYRROoBUU4FXiv
a2i9HD0ASAPtF2KYUyN82yVD2mnsUkz7OPR2i6JMtjDhy01gqsaSi2HI/dTzXUpn
O2uVoVRNw9/sDH/SVEFkEXq4nKBPfYeQOD9Epdv+Z2JmnDFd11vDSJRCxfdcyddT
+928cwAeIT/O/jI3HLpScpYuzjaUu7VkdKyTazcStEx+pd7I91akXGRbvFMtw8Ok
+Dbfz4dysiqYkWBDjJdZBA5JQuY4rLmMgvv/grDfK/dykJAH6wJ47wt4C6a52lKu
wOGQqlipiq4of8mEU4n1hF4Nu/uVgu5w8emN9WPysCn0m47+WHEPtbpPRoVjqYOd
cRce2crrlBNjQ6T7NT8jcqhXZLvPB8wzKXWYRLkTDnSb9sTuKGutxptnVIGKCKn0
c6Tfqb40FbDfZ30Ebfx2Z/J2IwG/fzqXnglW81m77Gk2p4j4DhlmOHwLwxVA6nYj
CajnrT4y8MmxYm2j+l7JVvZh4oYPgt2c1V4z6et08qUCuxdQX6D8M86rX4ju9+PD
2RN06TyEYVO/vZM7cLp5rgcKZvLetDmpvRBIexjX7n6+28UwMW092ZHyI79Fcott
GftLjfiLEi/fa8eAN3Q0+pYT51w2CJfO1dmI9BEN6w9yYkpS8fJ2tIag4HvPG4MW
6E4OFwvkM/dI1b6rSXGnGOsFJeZh70CW5CPDOg23bFa/vCLsLgYcoT/lrTjAHOnO
g3GY3F23O4hmOUh/xJ8J6jNyKXVMZglxVwUVjWV4PKt369T/YeHdjNphKHDvwDWu
sbWcErmNPisK766VLGrXUQq+Z0+9Y3T2tHVwoaBEiv95wBblGNV7spgEW+sHQG+l
5eKg26pnotGLJFfcwcROj7ArPiEAP2lzuZC1vbo+C5P/Wzqxm3q9QU9naGzyZvnF
pN+ZkgQVuHBCXgpnZ1GEnPrAATT2MLD8tvFrcaC3mfSULV0rhulHppqP0tRlq5Xo
wXhBmtyS2n9maeYtfi3WGmhDr70u3F1+Imgpq7GLt7nemRDd6J9LVcvLRZCyOU5W
RfrYczghhxkPG+tI0XGmZD1LTuVHa3dwwDAgE/7WimsYHbuhewImNw4OdV8fB3Bb
+frVpOabNTjrCueFyEpS9HDQp/qjgT3vb4AfpERw5XFLam1v4adkyyPtUXkDNfWI
dcOuUsVYaVwCZKtLJyQzAI01vg075irLkp0n8D7g4n8ux73G0iAtLdFfbPZxm8qI
sRlillJj+kKtKt1vWNPLCBSt+aC9n+XjuTbfYSO/4SvaP4WIgpvzFRIi4ZNLNJmU
FqGScQ+8widETPgdlg2y+uaXLfjZlcVJXJFLvU0PaM9NOfGs0KWJ+YzQ9olvHw23
qkk88aJy4fcZs7R9kUgxz7SBvD+C8jTtAkYkufhSPdIPDygg0LyFN4aOf+Q5tba5
Z5qJFj2YlbrztjM147fJtJLt/3DpllAQfikRkveZO2BgZIfDBoQWG67Tw3Ff8Hjx
d4YjCErX6YaDttA7wbdK+LwP0zIIVznkj1xcwDMdipYSNj692VEOdrnfRMWjN+bS
cZQmRlcQ1//nCdv+6XL6VDUmfup+OQQPqQgo/kg6ibf/EmOYJi4US40esib2wMij
Sw4tGlqoT8dpn2S5ytRXkSfg44YbkevCjeBzmRjSKG/dMFtTxPPgCaDW0z+YpqXC
KR8fKQsUPYmONFYrILFfjePipaWy+Oid9c9Ig8+cpLBCFk2EBr+3kkUeR9WG8bJQ
vNVFK+LhwMX1gF6GL5I2dNhVoWKE6KePC5vYjvsJRLW4Z8SQsYaZaSSfS6XBRNDC
vPPQMtitsKCdaINTlvBLQLwvNIyWvDY8zY3ZKef9dwy2ezoGSaeOkAUqcTbrFLrY
60cTpBfFhFR/AKay/3E23SXjsTa7KOPEpQFw6YDKW5Lgxcd4wErL9MsYnhKGQPWh
z5EBMAPk6+4kn9Z2/2cTDETKkBjh1FDZg2fzCNYhlBvm44CUH2DEEsQ1oDFGcx/W
9ELjX4mP13LNVQU+TMAoCu1qVKJxAeXo7YNFsidJVUB2e0TvUixAbshXiMzDybxX
fOtKLaBjIyjMRJiqFcouSA4cy7Ov7f8+rwgRAs+KoshZ+ED6FpffrDr0T8cvA/8m
U1Dh5O7JXrbi9zDOqoq9R50GnR9FZUItDsWL3ORd+QwkxXHeFjUDyp7WKDWDyLL7
W2DORgnJAhXIEBN4rzFcX/dzvuPobsW4mMtiHysVqioG/LC9d7ApPmHnwKwS5Ke0
kk0LasCr43KYoGmdsOxFftGAceNs9GfAK3mZ+6ydwb3zqyyP0ZqGHX9FqpWpbhGi
i6W+ipVLbU6IRyDBgGMfKq7o3TY0tLn+fJOeNAmHtaGHs+Fhp83YdKdQsYffPkrL
KZKLuX4liu0Q646EMPjBDV/z+JrQ23oJyDx6G7STDi+JFTqV7jy4fgzdhk/sTmi3
FgyPesDqKTHtozMeiarSiMKlciDsp9S3v8ssUK/Xed0aesZD0Or/vz8RYLIwO+ho
T26LlrSgneLIwKRwb3mqHbKdFwfHqyJo+H8i4NEhHRxeqqkkz5KgP9RqwU9DTpJc
BynOdou+2OPjD80KAczOIhxYNw/7iJCr3qf4acO4lDxpk9E1DBgqOipnZdK8e73L
ixLvnT3oCnusF8Jk++YcSx1ChDit361SStXujTIgkvamoIta5tgoQMovSWTiJ9//
jKDFru4SBvGyUQQ+CLWqXTYcC/KH3lAxsShgK7O81rl90wPMb8GxyRG4QiFYmcMH
C5TfqxKAHauMCn9xcWMq5JVigr7TXgZRphM43UKVxYbwTmwU/x+V+LU0mMK0UiLS
9M7Z5gjJU0A92amzV6luT8BNcM3bKniiNVC7QaKXjxvIsdc2/ZorsInAtM6tqlwF
HvuOn03TTOrUo7MNoBs/2jnCJ2JKqtZoCQWnBXSJ7mN+4SVQgWSC69JJtWe4AMgk
6iSO0Xj8iSJk92F+HBEm3Xt8AHtboLxeeKeBLJog75wd1bx8rqT+ySg/SloUAp6J
OXBcRjBK2kQYpqqQxy2XoAWGeeUn+05EUq+HpZFh0UzLRl67+ghCnD6395h7EcU9
aQZEDjjD0B6vaIkRPRBAPSy8slRtKXsDQKSY8pxc8XTmNxziRbbCYLr1xh6pXMcE
+oDwBOHQNgHYE4GRdIAWftpeFwggL5BdgoewZxaXe+Dza+Povit93zwgap46llWi
c+XAYHvJfPmtWSJOSS168iG3u6k5QbvF4AOWE3x7aoeL6j1UrJQ1KGviQlejkXN1
Jhli+x+n1QvkdDT8yrZV6Ix7OM9iT5rzwIyUex4RBlfgvPxvnzbIXumNYagKQzPV
BUO1NBXJsduxaZR83Jh5ZWoPrKOHAmrpSDmjFqge5AO93F8QeBjbqMBou1Pki35o
IcvkU4Url2xY6Gx8YoOxpN97L4e9BPFQwpxx3+in4/alC8kzqxbMb4AsELquph+n
1HnZ46zg5Hqyk2IxxKhFB1WgZqsgjdWlAL4Rz7Y092gYVlJeoII9YpGH8f7hT7ot
YK5xEaGeLTAqy/zzEkDwzV07qlUnwM7LAjawosoBEF6y4O1zkkWQMhqJ0D8ElswT
2p2YKx9KO6vShEmo3r0aCh1HFOP82+b2juyQ1olHkyhHvA2n/qnzCxhSrCirJ4ci
n8UJyvZHkG4HKdUCZ3/NOTenSeFrcaqSCT1MlGaRwzQcrh/5doGEJOHzbF3Besvp
JC9UvrslLar4WAFv2BfHkkvwmUoyCTp99/VmzPYMEIT2M4lWwAoz6RmR4mcnv019
U7/mBiVT/7lck1FQ5Wdlx2e7Pb5xKCsZeaOv/NP+tOg+7cmv1F/XsL1pQqCLGMAN
I8+MlKEBJShDoel6UFXVpxAQoQf94oHLlTkh8lL0fLyEcn+zCRt7YQlWL8UkqnmO
2xIn91sVZlN1vZQv3ndruhv9Q4X8rlQZXNYr7ft66KF2WNN16kRibT8naW85/2Rq
fyAMBx+LtxbUCX/Clx5oCZZOnvNCTYYhn0RuhiAmgYtf+G1dBtKcRk6YOLW7MJCW
CaGnxPEydAMad8hnzf0FHb+w4fPWmYkCLVJDKSwqMOeJ3yaa1wBFE50XFxuDAq5t
PlIPsDwLaPqqJkW8KshKQ6y2jaglFIOCB+f38d/X8USYK3KsIaBcDfbdJnIllLOs
F7z7tKpqmdX/wVwRgrewQONfhKqo7WCvsSVV5Tvjmserw4MY35e8EkXIdYIgp4Ry
ESueg528+mr7Jd5+rGBDEuTgX/ECJD7h9jKVc/n7oRZ06Uq28+kEo55weVSGqg4X
Eh2DCGrpSJrnMiFovWT3sHosxsY/aN/mAnEZ4jQNJGB5u86BdjBP8Mv8VAaUmEya
EXTQcz6Qet2HGMnnsgp7yA9RwViRO3oGrsWEPn7gL+DZEBTKI4IOP+rqcj+BjhhX
+g4VqRwXtlpLgCmtV462oC46/3LcUgf+rwJJLIyYyFk6c8eFqsRe8vjIdbkrbsx0
FyznXgVhnD20Vofn/0qYstWWQb0XKRahB8rIxkjmg4f0f8PwKLWbSEqBIHzi9/sC
pV4K2yXVbHflVpRBkr0c6BlGCH7x4F6QZtrxqPNw2wqHBSfn9RVzi19frMdupBuB
SeU7wHc2HU0WE8mO/6aJhYiAsO0ZmEa+WrN93VBoERLXldbfcg6T97BM+De01bY6
RQU+jc5Krbe1o7nj0fHV9pGH2rfLJBaE8V+jH1AGuLMk5VZqbuctFfD+c0jCUpyR
ktCPbd6+VjhkO2YlpBaTpTFGSAzece+oSNX1662y15MxF+txf0XS2ZagY5KBM5v7
x/wJMUqR+l0Y2YbS1Vm//4njZQQB5JWCmIrZ4KkYM0r47EhfGgciX8IrqCX1gggN
HMV5Dsx32lsb3xLypkslcG/cMzoqZw1OOGfxl9FCgmqgBC3k1kcIUWawYU3VyxB0
wGqlEjxzi2O+FD0WalddNHzeY020t12msh20qJkbNOVJ1gOduBESH0oP6zmbhJ0Q
JxxCnPNo3PAqTkPtehKgrXg5H/yC7ISYRXCOjc8t4G2yyxTvT0v/0IAnsX6JVN00
eO9ENe1A7xKW94BqBpDbcFMF5EZyrwMrZrhcjFi/IH/7eRuM1LZo0hpTRlD29Q2D
8sjGB7UISzqkIUk6bEA1CJ007Wf2aDWsiO6idgeDBHXLoYcEjF1TGzU499+GB4ps
5Ek7s5rqA054oVaqpKI26CP4IFRxkoATRHjFsmXk3PQEp4qHotje0IGeXIO8umg+
JKK/LTpDBud1FkS4gMrHUoTQzZUGmmzaH9yIZRPiZCccCnR/VzdsufU+qBXCaAVf
Af4KiMLNKJpdTLepJygfKLM98L12zYH+dn/42HzaU5o2p224W8OTSsFGi2lEFzeE
3RHQL/DdIcaeeHp7BJxZIT9LKfWmcKqdUnoWJ4aCUOZ4S0b2mIsjaCclFG3GJFG5
DiNGdcP0EL3vKgwBjmqMuLkJFwXFibiJH/hRes/RrJPnK2WAMs7941uLl/1Lp30l
qhTtQfw27J31NZ18Qwffnm3iP6unQk3wV3bGFCxMTkoDoFntaS+TctRenWeOy2uY
Jv90pomv62gnHpb+Pnq4ggbxyt1G+guJLuSWrv1o/+NR3bfF5i1IHT6xhpf8BYVz
MQPEA1k7/koBxU7YigDckM4MAeZVhgdwuXks77/yvkhQz7ZilLV+4Ssy0WUq/beb
erY8PIxcdqmIUgckTYFTBtUOY3suD6/XKZRejovt1ukFlWJ349ZD59MunlFk+PVz
EQdxX5sHBy3Y8X8efnDhjsINsX+r9hdOb/yEi/8UIh+9JEttroquzcohv+c7MkAR
lR+nT9FPlbMxWHFNBLKwEgtjoNEveL8VQBBiEMKZAq/+VjijHVrhBjtdoirBeayM
g0JKSE04Gh8BShaFM4DVCxeGMsX+o4U6XX9AcHVIsgS1oI5OE8c5WjXBw3IkZ3Qc
pkpZTJOtAjY4MpXmZx++1ImankTh2wk+JpZ6B3ypotJXxbStUwC2aG4bbM2NHunA
fgW25JaIvDhdGmW/rf6WAJIpKiGGGLNzxbyjPl2b8Ynx2CsbbPuc9aTKhmvwfDmd
jf0N5qEDwPx4/oIfEHtD3aOS6LLKyDTVwnzHqiHgQ5qrjX7gvABPzUIZJTwPaZzk
e0iUPOiGIepo4KCCFdJisAXyT2zVy7EV9aJGYxa1D+kDuVv6N8aqpgRUkcEABvTt
Fdr+0ph1chlc5DZKK1HbBIj0fZKwC3FZumDwrwIFgZWlS9OhdJGxO0k0bpPjppKS
C4AARispgsCulEKgVltSmv7l93iohZmuSYGauBK/j8dkxGupCCu43xOJo0s1fJqL
fP3u8Px8ZDDcF/L6o1qB7EinV6F/nV1f8NKL4tQcKwGU/OgJDOmEr00c8nF1BSg+
YmqHACVKiLPpX6w0rjOdLb6M7jqs4GTwZojx+byphXUBPCUGdsrAf/ABcnSz25N+
v0Fn3il5vJozeUGpEgwn8chmHzlOS5/DMXuJyXCcxmOMK7gE2Da+UUU8Wq1gXuaA
NRBLPYeomYYTACJbNxBpq5ayoSkH8OALb/WSkVebwn1+DkuYI9LbSx4TULVg2AFs
lh5p7efIeWhByb9/LFpW3b8MO8c9yq+Sc5gXfjhI39qB51XzBGn4qSTVOlu5AhTf
k5Hiz73O8Kt1aB//JdZ9UcwmZqCuPTgeAT+G+fTrvhtgj/qJFuHfXAMfmkk2Ca2B
b8PX8BWFPxdMievR059YSL3osL2MwGBy+GbGjk41SGrOZv8MPzh+pEIQbAbBXofs
ivofNsaEV5d/MmU4VTCrMGZn8Uar7kx6NZHoi7bVNJ3jjyfEA9F8fkpsni+wBicl
Et6CzC491d0X0G4tvFozpMz8/i0OeSPQIOYkGRnyqoMhr2HAwKvvS8Si+F57wQpA
NaAd+o4kvLAy3Olp1HmMItILP879XW20zQXO9daqCK6gncBtb57fCX5Co/Y3cisO
OztuBoU0gK02nqVQPi+OU8KaUeMApewRJCOcJiC65Oeaud3MmkSR+TTC2DQAPeof
F7nXTfxVfFJWeeQs5XHlgtO8cJUD9rqozcg6h7ZQWQOfMPqVJnMoaJq1TNzEozT8
shoH0e1dAS4DOZ+FVvI+mAGTxQs279Pf+A9U6Jn58qgjlq3cEd6lW+H6jrQY4T7i
KaXxIRLmVs2WPjP+RcDueUZtkPpD0ZaMzOteCh/9ID3BoVyULOcVY5jiFa4v7Xat
MIfWaja2f/6TAf1XZJPQ07s2kpLq6BYM5Q21sa/+KK0BVLIxLFztby79ka/aOx5z
Z6g317/kHvSJM1tM9lveZoyutgVxsVBJRkrEkhiiy7Ax01w84kTsVYCx9ZF4ZbBB
ps91FiaLBQlGLElhVTqgpS6FX7C2Sw5TqInEUaVcN4DxGzYAAA/DS6KExchm18LB
/6ZU4bIVsPC+N+NhHQVpUqn1+jZ3S4wm1udAMQd3XpkFFIZKPq4nFeJh2SME5Db3
5jITHrpsbgUeodFsXMPzkkvzkivnPPs+N5JWQlHMIb8yQ50WVRjIw/Qud53HviCd
eflu/buTyJ2LP3bGzsCY36iOWJN4zx+lrl5c/NYfceG8ImLqL/RYVT2SXVyMzqgl
ncbwy/7XupAq9Lu+lNo7bXsW9XaQJSqk2buKt1rgHBwgMnmTGrOcsI1TA9+8gD6t
Jr6aNe3rGouAjLXLlKNh3XAWN8WvOimZ7AG7Wt5h71O2zDlWTCZeZ71CwYwfxGD1
nEPzdOqCDxpeUuyojlM2CljNLTiJTvkZ/0qBSz+8aNdkrR4FaVR/6rLbvTypLRlP
ZMJcMfYT4GkYzW2zOBgUvSe13vN1azFVww810Skj2HKWTIdptjJRQy+5gdkFcB7/
ZLsA78gJF2Y9RoTNbQFtCkBu0sbEdVbh5rZc7vfVA28v6k6mzcLyry+ncoUZvRKn
OjbHhvC9+g4tj2zRg0eF6q3uTayO8R1eaof/JcuQWtjET+svXnN6aIHjW2PjFmS5
3CWQ7ZtMPHFJMBQkT8NKD8bKKrNWjQVhmfrkCgiVM70s9mXW3bv3PKPKYS5oZpCG
uj8T6nLNaU+zHeCVmZYCYleQ9iyHQzAk5ZSYQieBL8vUzLe1+iEu2q2kSvUkbHOB
7XoNXMXTqoeDzFtIzbxmxwE3i3WfisEDn/0lmrvZ3xTDbYqF/UTEWfq4eEHCnUS8
aVpiFcx64dwFSSiawS/yWUcLIYLqBBA6HPmY86871JFdJuZ5MhnfswrOhtHxntSD
DKgIWBYVbBqpSZgHhBjQZWpJnBWQVUMyop3jc3rm2wGfXGTDW/2WPonuAn+brKtY
70C6a3L+JiZO8rd7d2yJtW9eo+ItU3IHNwQb3bqdUyFRYXJfPOb1YnxZ3RjWaRNH
mziiC2K0ayfgrx3DNL2obzLN9Gu93yhtTQtSpLnCpkRbyaDzUyaBtyKE9pxWGxlY
qeCvJq0KblsUwyqpMednn9ROmEvJYWR9HpU5h/Z7f8WVcoVHq0LLu8mYhZXb+01P
JhygBcN5ZsBQ9xhxl5My6IqIu3Etn8yjpBXpTQn35vTn+rKg921eeflTauaogTs0
PSpCRYF0pOqGMHs/xIjcVQawP4Vy9JRGWcztaF9Wn3Y9jC5NVa4E0stUPLDI3NvC
0y7yCIh2FUM05I/vsza+xz/uWan0wJ239gCpQ3ffCp9hS1/9bkRhP5vF6eCm8Qc+
lQ6O3esMNBwCVtCFZP40EIwYWXS7sJjbe6/BKUDDvyya43aidRc6YrN5CWA3ioCB
ZvcjUsOoeewsQCegW7uBlp12C3QzjX6pixH3MPVQrtTFT3goB3yLK9C65UDSosCi
uNffzo6hjG8CQHkqpIS4KUL9iZbqAdmVX5G8gtq+n/UjyYWztgMC8IUV8B7Yjipa
YIU4Bmb/eGYtSZHExj5H3IwML3odllE1m5NoZuRms1MQCb/6A3TqrC0PKG67uLTN
p5y/YIYqi7N3AnOgLnfCpyKxF24oYA+FzB/v/0yjlgYKIJHxQZdPe4XAUh62HWYH
ALLZyLJyW5YTISQ74QBwRDANd0ajS9W4rrzVAcL/OZIe3IF4OqdEgp89gFJunhDI
UEbWe1WpkrVej58qy3hfFbkLlMLbq5xAbxr19vGpZXjyVV2tiesoZ4V8MiKWbDlJ
aU6AN48Q7XDy3I+46rNiaYEWuRUStzV6GcC63+nZlYDCXKTIRc2A2N0/UEbv8IOs
OzN06IyrV3rfhe0yWebntY6k8Z/rSEKc9G/uQT57WLsFIxgyMcyHyuuiAFcihFEj
PJD9UmnrZ1/bl0ibcGS5IBLHlMVCX2t7mruXJHyjyX3tmDabcgQxJ1XZqJXWk67X
nQakjVgBypioUs6xLIt39A/4h/MXpgdCeTMEQcIQO9w8xbK6aEiBqVFtTDnyPqLe
+0B+1f1f6PdyTdcDKgzNuojA9ngYURaKLTkFOgASHkoxzmYBb9YA+rsbwbTii5Md
sOHvPTMHZU3tIklLWH65ejNX/4Quglmig4lPJt5FJD7MUDkk7qfdLmb4v3ySvpLf
3Mh8YHYP3Fydt9BYrADuyPrC5IqSIbbiuw0SEYkIHVAIAaLHr/EJoaKZgwbBvM3f
pi7ahHEMAtfjZ+54r29THXM7vjFKDDxfgD63CJewGdRr2I3uNcucf3rl3uTOQJoi
aFc/CGrghUhQDi7lXLr7iAJqaVncLPuJsVp2b7tymYyL6Y8w7/LH4CrP+5GhpoBA
RiZm0jGJszCAoODv2Gi8rCR4mnAb8a+bqxKIjyXcapOsl5CqlVQN7Dk26EMoxqZo
hkijI2oVxY2Y/Pes6kSZ3zQcAPWNNjxdSow2S+zzQkDIPrgd6lwDYOz91HMkFr9n
TtnoHy9M1B3ci3OkRl3tsl3bHEcJ5OcQQUhcmxa3Akud1uM6FBO7LUU1QeMmnXZp
hKGj5nXLn+Yp3ZzQdhVDp+rxZAkGrIC9llBmRQchl8ge1EHI6iyJ9lAjCdMfwQzP
KwNCHzJLDhG+r29DE3rbvu2Bthmdx3hJWvQplP3bwKJyb2vWQa/NlGHADTh5MVtD
arfghuP7E9cIw41vIBeMWVdpM73N1nXAgZiw6ABsLvosNs+AZPa1/iZQ+ho11CbK
mFyzMT5uceHsd7QM9zkiSW4aobrpQa7TS21pyEULR+TUg3lVVFcys0+9kLfMybTX
RKUfsttAi1w5b7oPv+7vYEgnbx1xQlIMp1k76IgrtFgXUHGWALzbqCNsHlD4UxQC
CNSAv/W9qSk+PARrgyEtYFdzXAayn42YVIFiFshTITZ2BEQ1Rw9d1OMJyA0j06BO
IMYsz4k+RBx/0G7nIvxVQUE4w2jeH5KH4LhWHycEiHElIzMlGuoOddSGg/FkP43w
Z9NbKHVZ2jS+j17ja8OPNJzMPLcTmXfKj8/nlbthsiK6YV8tuBcc93e9dpPy0nrI
s4oX4C+5e54CWKpT7B9EFC16cqke5CGri+hmZXA20IrrVkWhL2AK+VjdhBk0+eqC
Lc2ALSqv6+aLY7ODP4bnMn9NMzcvCUHFtYKIuGrTYRI4+3Fx8BCPcl4h2zJSIAxQ
rLonZom8KSFfbK91Q0v+SNN7XtUrFoSz1Jjrl6xkJtNH4Ufw4iqwIDoHFCpjzDRc
vkXZU/IF+kaC74+zVb42zlssPOHVet66mQsuLUtcmkjARw1x3dneDoTaf1paJ2Yk
Dv5l2F4/HMVMO5S4MLijRdCF3zYN9GpvXLS7egttLrHkyxH9Hs1qCbfsGm4wDRul
KcKZkEpA5CZrG5uM4vONw4EeTpdMhVOYdNw7KQE/eaAlGgFpT+kiDYw4f5+hY/Il
udEMiNO7me0BhZ0tkC1T8C4q/Hu35lElIAQcpYk0odMJZVYtvFgnbCyYlkfqBXyK
nlyYqMangEx3tgu7Iymxw4Hw1l4jF1I9xru8nYdWQciq6cq7F2LcpIzj4bCbMPws
Q+qEGAqIDvQ3ea3tlON/UANVKkJ0Q9J80yOmzNAZlBn1Haf/t/qREN8PMJSRX+dh
HTSSY1T2kxh/O984gpzy19Zs7fF3qjltZ1VEMtrJLyYJWErFUE0LfF8odFRVFhr8
hvra98183Otcz978TNbVkWOMDEMxLCof++aywokA4OON9s+Vo+NPR0Q+vX9X5wkq
T1MhiD+eTcwKlf/GI1TR96HXiW7WQP7odKIlkRso5ac/O+8smOv/aHNYwuDUwmRl
rjCGhKs5wALYxWfczCiGTcdgCYzLE3A8BtkupJvfMBMzJBS/nPLeg9saQhBRUoTX
JFVwEXTMCf4B854T7eTOAsUNUl8ymqASsE08LFIwaFB6g9vAGt+0EeBxvc67wRbH
t74ig8ow0yv7FMtQiEDKnEZx5NOfzy7psBf/s0BuHTziu/pVL+EtXcNA3hZ5w/cZ
Gheuywmfmv8LEz6cxuJUY/9Gj5RtA8ZkIzzWcXEDlFacHV5ql5y6dBxgHfR45YV6
HEnG8aEbv/P2Jz+SPDiNESEOUgebO0v6W5/ZdmVZE65IcyoCeLoCaVDOKYO5Y53N
gub0dJv765vX7nxcw6GpU/Q2X7HA1+8KFeu8PhanLB29sQhb0+SA5LVCxUqTieP3
O8//bkzM2G61t64g74izG/3P+BUThFzHBt7nfNmYaORc7YIJPrBG7IN+yznFGS3B
YIbJAOpz0THG24JvOU1Rq4MpOV+M9UCqsnmMB+9ruxhDaY1mpkpDuTQ+qjcB9iol
ZPblf4arwB48VM10DxBUU2VxoEEj0uNfqvYk3p8MU/GduEWSqj0lcgTQmXOKlDZw
l3iLJdo14WoEHGsXCtAc/60Lav6OYp27O6rLbg+2P/UPZM9jtl1q9rmtiKYwsAtz
9W8MFSENXWCoJyzLH+XFw98XiUR63fA4jQJX7GmHzXk3iD7ut9xPRmvHZgq4WcXV
qZ7kkJbCBokfITQx+X01v2n9+NuDew3klh3ZpOVCUObjMI3u+BF/teKQYTgMtdjW
w9u+pygC/RklhmUYXAgQdO2timTE8cYHpMGpzyUGZm5jbMeqzyWwrMxgWbb7R3fH
rTRETxUBvevVXPtKb2vk1/pbkTW0KDKkUbhRFaMipU4StHGt3F7lSUhso1ZfOW8U
qsaiabMrB3KqjfoRuPh/sta5R/NCtUGPJdTrh8VdqsJ1cvBeS47t8DMsm+wIy96m
gIZNJE4EXizYqu4L9Kw+DVJfZ/maUUYb68dwFWhpq9fBZBpV++Qm6EJ1iqoCTdGy
V+ui4Ued0kqkYwCULE1RM1sw3QJT69yPu3ffox9Fzi+HTjN4e4l4e7yjnD/TD1ns
DZgu++bNAVJshPPUin42yhU07kHBUbOGLq/D7bicmkSYwimD5sVi0ep+6WR5ahxw
HoP3xI2tw/1fGg5KDpxwqzwxGH1o7CSNG4wiVfn0fMtvtxicK8XQeTQNWfz3soOO
CP4szlmp4z/txoYFvqssPzST1M1RLMY9HSIyPAnc+Bq/TDX5hldTDVOqcpAqUuxz
PMOLPNo9MQ8SU181oFFojKIIBhhFE9kICSCgxQ+G246HY5oABI7ZPIhFI0bxn0ZX
Gcu34LgmtiselD1g3Ub7qvMYLeEjV/f8cmdyLb07a2tmYroEsVanVRckalEYjj3K
jMji0H0PiqRaalfK6iY0LqrbiRWUckHF43G9h+ZuSqY+QGM/hdlng94Zn5IzXpYv
IKJMF05WOz8n3gCkZRkRGalm/kckapk+K5+08cSSdgy6ugBxMMwt2tjPQZ9jjOwV
go6tPMAlveRi6yJlTAnlfA4AXKgOct/SP5fSGFFMYCbkUOCcexdFTehBEMIqRaWn
PWYVO1cwfoIeD2J6GutLwBjfFjgljTDdNz0f7HgVEO8dWr/0w1i7JvkJKvTnR9d9
18AuMk+PtWv8HFfH/cw83OoWE18EM6Uhs4Ac/Wz1q1PuaRUB5oPfSOAojNRb4hRc
2Qu2dEMAiMDwwNyFflBilMSF0GpU3s00YIeuNE5UEgd+NVgiMsG7xD4+Yv8jwWXR
TgAM+kZHPUjsMydBNv9Tdb8ldQqxR3sRy7RnhspFUCu6GT8+MDK43Y0iajCo8bVu
3p1LskTLOfTZqBKC1LmX13/BrYvT2taSAtffkdk3rSygj89zZJLFDPdqXxgSA9e+
wajbONXof/Ks62tVlAdtqK+EMXkQOh1Q4g9r9octIiA364+SgL1yXi4a0tkJ1esc
2fgP0OyWTB/hCioVyQhWmDwRHt8NJ7CtU2GwyJjyVS9hhq1F73f8SJt5i42tcUiB
ad4/eepETOSxqgqlQZUqMmUzYeGRLNZPYcjpzSfAz/uZRExt6ZB6kZzCLZFLFg3B
RD5i8UQhlNrbZvheINfbrmuA0E54gen0oYMuk7K+dzlSbolZunpZ7OUYK8epor/U
aY8tZWuUsNkqms75u/mF+fcngCHRiTZbY2qtLKyhtI2v9WNyQMviaolaDXKJJNLF
acqZZW8I1/vjqc9zknEX+GnMyKFWP65xnxHcyI68Pc5v7+QUxOiYtNBsNgLafQsP
SahE5iXYTcbsLFeFArLpTtYXzyZTjxDu4ERbSWtASz4UC3ZzfVAbqUzJgApDRu1k
Sv5VaOnYibH39q3tr+nab4AoLoqPQUcMbkR82xvC+DmOZh7kS1KFwZ77AIqALIIE
9ZaGtMjHG3+HWeHuXGDIJ02jWRYyW0dYvCzAIOX8OhL0PGhy1j/FUH6Yk6HrUejU
xTEr6jaY6DJ7r2dpeKUcbeu/IK+p6AN7KNX8M6lyCk/5X1rSeoVeryvy0v2/8ngL
hYTqF+CPB3vp6jVQBbwUIHwdIHFmA1KEtUNDqCrbnaptJ/uwPQxs5TSTZxQFJEmV
HgWnOmj7UD9pdH9LsBOLCsmOHGCGMGho00Wg2S0sgSlKLVytGM0ubjiC8DTYb/xy
DmAySHimp63a0DYZe3ET7o1f0ulBBnjP238ZO0lhdyZGuVBmPC5FtvUGEFDYazTg
5KqZXacC40Bbz/oQS4AvDDRiw4rq0VvLwcyQdLKRSuKtuuAblrRDh2hzgCour3rI
IGGPYuClLO5O+skO79rcP+cLMpqG61+37hSwnqTy8zDiXDpn/XbuV6qXoLfKryrU
4fOdzpcKnVw5ncVLKS4WYC+SS1KmqexPkoJDkUf484KDQeScgXE/DzWbssF6eh0I
HhUmQSIMydC0ZFi5cGVKbOtgw2ntjMm3Z0CJL8r8kUkZeKp6fz6QSq6Wz1cxzydB
cbZRGgKX1kg8xjX2cZWdEtUu88WRTJgnsY4XTRwqYaZSN6gZ5MOkuxtFbL0SpGDz
1MTF1cZsixkJzZdGeWA71VaMx2Ft4kj4r45DueNwrfO+L4LIljFOCYQRqEwwNpHe
xxapnhuG2lRU6CnALXcoeT+CZoUXUuAjlG1oZQYV32dM9I4oqt6mSQxdk9yhrD1O
Pr1QmIn8sDh14XZCmP6YOvHc4wRIoZrGSVydAxlKCnQ2Lm1ZFfSgmIb+rFlhdNt0
5cvdJdPhQVnCDGMW+PFuGYXfcupAbP2DQE90njx+EV2TE/knT0r0JiSMrkRP0JIn
ayw6dAgs6U7XtrbtrULoil0VAOBHR9dOi3cXquPpM+/WemE41JtwkbvECVDxXmLy
j8NpNPizFsPAXNJzlaogivlk/+LmmNDZ794O4NnjG7DRXjRwbhXh0cOfMA9apJG/
zWQi8q+hvb+SmnvJccuxUCUgSv85lUSfa7KYdO7+ThppIQrnkH88qkbZvfYZ3GI+
IDbZt2ZuR7ICvBdoWyc9g9Mca4+tckkUdcb0HsbtdSl8hqOImAIWY2XZMGiZNe6Q
FZGVHD65iy3C7B5RnNxC2cqR/RWxJxx+vzarjQ8zo4WMs7+pyk8LHgdDK+ING38E
M2KU6h3mLUMLywJijjdG2el9qxwI4Pvdpxpphyjnokhus2I3sxeI3od1SSeb868f
0P4IFHuuBt1tgGp0uB/f+36WKWPSQQ7avUJoSF4uEPZ8gGM/+ygEfAwTIWcvMQwD
MitFx8VyRvPUWNJ9W6Lnsn3BJIKHrAsasj2dowBVNE0CkuKQp/258nAe8dzkR1nJ
E5uol+anyL51XuVp6THZ6zyXj/LL0lWklArJQNrN+OOQHjJkikUhPYt1uphig8Od
M4Tk5je6i6VRtNHo86yzYfocIO+TzxNY23eAZ/a2xKf6tO5cUjLij+xdu6OFDEwJ
1MAIMNUIwILcHPMzDB+P0je0tXaLLgBp7HHKzdMT6KrDhcHGz2GL0VVm2foEKiHm
6pJ+jPWV4DwNiA8YZVG4fBnGkRehNtdBM/ek2Qtj+vOGxlOifTLihJYdZBanBgAM
p6LKzJ2PnE5Gf6PGldKZFtkig52ZQA218h3zNPg9SiCBOtYBpBpRnwu+x4v6Qvi3
nU2nUnnZYsOVBiEzgfWum/1WSAYEGpsMTra80c3zrRIyC2CN/Ka7jtBqWfEhmoW7
ekvD0YlTzi0XZ6LYDZhPrQGyinaazuLxER6iV5eoHoSXw7hnFcs3bnqFLpvYTkgh
lvx2dUIo8u0+WaXIREGIQydVpcP6C+VhY5z+PPbE5n44SApsZP4ylJF+A375XK2e
xrfc4XX9lLEXkBH8MF1FHrmOdBxudnzDO095lE207RLX//0q2ts60IaIoxhBuAvU
GUxEiUEKqEGXyzPkVbPWBdKDHbHp4fOJuO7ivfkutU1uu6xnubPQyacIhH+tl8nd
k+qYzIr09GKRS77s+Zwp5QBxG4HhScX2Bt0xJsBIkbZ8N+z4csoFvOfYxzjl+s5M
NOkb08r/2DmOEKWxg/cZw5RACPfeiRM9YW48frtv03to9qBFGhXf6meJs57zoKBi
Z+7iYpsMMNsT9elUKf2zhEYZbLONy+RkJTZdqwb5KMA91wFyB5kiCHeZEFnynV+Z
hXXI6MRvYI5O1Nd3MFN6BtqxPrOQPJMaxeg/YFbnHReHSQB0iJefGvgySUqIhRQP
LQjEHIwnLgZ2eSbZJF4SZjjodirZvN+hxt7nvaSzx45BGcGefdCHdXpDuW+TKBjX
0jQll4NGiUMGRCiY6SqrfqIDg+p6D2p5u/H8xrtWyKz6ZtsDJwuR2T3y+PETMASn
0/gfv6Ks7S2nYyFWKybuLLALRVBtwnTisGAh5OXrFrB3mQ562Vi+UeGMzgBYEZt/
nXvgL+QZMMOah8sAcAJRpH9wRTTQ4xsgMq1Ig5CBW6qaVWyB5H+Deum8+ReJrzK/
/+qilryenMZ/0+1EJ2lDjfhakvIpBicSlPRuCU3NSXHQrocEv/XOtQ0SveVzsx+N
5mUhgiVn4LDmnQf1Ydio4g+N7/GJKMoimojqcLsC3vN9isJKm+DPk4C5vQGFR2hs
23mxVRi1loi00aLQUaMLpQFAmqfSpQcGmUxeB7Px6i34LdIM27je1Z7E/Pn6wHZc
ZKJ5TDApBcaQE0rLnJAppULi3+uta726crptzUePrj1gtOefSVuGAVdF5/leItRS
48AtrWXxBTmGXOU/f3qtKW8/OBAhGMvHRc9Wc8GACwcq3zfoMs27xMCYzAFgO5AH
BahgSZbBQKBbhmBhrZTz9mSse7vFxptPFKHGRoBeQ0bFI+K3I189X8flnX/qkrot
veH6/yxlrgg8ftYau6ubsS/YArLPcc0znsB5VxjwmcvVEMy1FZilvPpFlIBdrGKg
SeRci43N5j1cqrmosZda7h6XbKKh3WgX8mwVXIwqWaV6+LbKNwoaw503DNuwiEi6
7ETPTWBTamr8gJs7sTEX8E1d4vbSH2dM9rSGbCukyQ39Yi0Of/zLfbVv3FRLVs3A
hNkLaeLMspHAZR2AyG6p6b3hCInQlVrk9zMZL6p7epRv1gjTGpp/HaBdCWL0DNKG
zQIXRMErFu1yFNLhbauSBXCNCCz1vBAI33wcyVUYy5uYG7pAiGbyEctqPWSj5HLz
zKeATWhSCwFJVQZyTzCrZVbRBwsbN0htQY2owwY38N4SFif+4erFFbfy3cm0fqVn
KKbhA7EurSpHh/G2GEelnXRt6KCThXVixOWKDZyA1n8ecGlVCdozeVXk9xmktwEe
1N+VzPkuRTuy1hL0UHVVf+DczwRLSSjD5vCoJJfntXIanvcmlcuJzIAP3hjg0IVg
9H+WR9Y7YhBscNabC3pwiYuZxgjfIkzzS9RnGDITe8LWb/jHINYRmJ5HZdx6ngF8
61SbAgA/evYp7VxOyTwB8J3dvp5yPEb8yruJrGA6AX84QZfo8zaxp81/B8cvKpDo
7VLJ2hWk+Ut+G8GbMt/3IC0y54DmWm3huBfrd3qg/u5syHHtKTBuPEUr5gP2owfx
Qb1qWUp9q40PCDuby23pB1lw0IxR8s0iJ0KoAIFfnNs7iAgzf/KYsJ6Ci5rIjH7f
Oyd7/t6K4+xgZQapLhmSrbP1awIgzQOAFdrgQe2wWHDJaVvY48oZX2XQy8h7Eemh
5B1CRY5UkbhFKfNYBHJMPdIB1Eyh5i1Puv+s6bMvHONaXU3zJdHY7rh5t5RQuJje
I1EB2FJA8tQVXywjp014a/o4A4e09n29aSEfMGkKlvJuJ9DnSr7r29QwNADVudxJ
QE5J3h1OzK8X7MDxAqERv77jLZWD/jE9lMsKTtfu5CFvisd/gYxhNYuGMwY7GRKV
fS16+iG9tLS1MWVZxX/AuhVQ4/oRlRto9M9y8ax39oRfzdmNa9ZW4HY+dz1LEn8e
BkmhPTDXg4QbEmmcP8V5gASFgsJn0GPaxGc1/psHD7VTWcKJ6YYbXY4595ET2Dzy
DUGs/0WKPWg4gR3LemyvyFYDQc10omPK4Hyccpc3XJ6Vg5tVyjqzis7yIrDWgkiS
xof2coXMuhaXnvvvkh+T1xRPD1mwoSYj+1Zj85/5aSlW6CoV27OUwB9d6bFjedwn
/uIwNzW4wPQotEYyIMcNALr799JTNBkc48lRd8Asfm9+ykKmOZzaaKvX+m2on5lN
rT/MtJLJ5q0fURFJSvPzUy0nrepwURO3arwcdAcYtVl5GGpXejC6KxNVvS2YA+UC
ZFY/GZxlNOAB9py5UwrjfOVqLleXVLciVGifLaVXVqa2E1PAKQf/ThsgvvBM0stu
KMKjo08R/nX3bEP5FXwHqVL0kNsIDoPSPJ4V6VH2M3fY9K2faKhwkq6IhPvHdrY0
agMry38f59SqERTC0PZpHweKyh0aZrNgkDEoO3+pLiZeXcyJqZUHHu1li93s1BPt
eCN0D0BQaA+q8b/lowWnKnzvCIoohvBcjkZEzqSP5WLiGlAQ4qI2fmIrDC+x5P4h
Fv/zFsaB3GajNzm4iDL6yU1Tx6av5qjk+XIbFEfptlrT2wc6KKyILYuvTZNk0pHQ
KQF0A0L6BDq8ehob76eysWpBEDVFIFzJUCa4W6+andsAizIZiPTAmAsq3KzpCod7
DjAGELzAs7N9k7Ariw0uZOoCl4J92j6xGFfOS24C/CV4kDSoxpPnPQHIc9ZCLX35
rwER7fIdQgOiig14B1OH4W0tppKn3HEyzPNyPLWRL0o8vnDKH7B+oJXUhhykommy
6qDw/Wa1++36fO+lcSztKSSEubTgltqQZAmkfLyL56y4SJnt6UKlKqjFqsKqqvlx
UsV+oRxa6Q/qWPlKE7blwlQw4Xy/FfPXMKVnVqvswjnMoRaNTMHSqXQyswyKWxB6
2KzxW/vFatrmCmpi2I8yM1wvxAM1NlgA9T/EHTUnU7YJmo7JTjU2w+GsOTFlNX1C
XKhvTUq3lhtLY7n46rv57cf76uuOumeHt0Yq28VzR+XvjMAVR27A28c53YyrRaga
Ha0OViiJfFqD08+3FFrEjKFmVVDOP5lMcX61dg7ONe1zcGS3DbYxZiV2oIX4Nq4K
D90JViaI2W92xfH1XZLyKpqIWBOwk1SILKrmECbB2vWv1MhsXIM37RmJyU/dcvWq
B/d+38RCy70IQuBs0+fCpvSkyhvub9tYcHaJ9+m8yNvF4BA/HrI/MvFI8r+m7DAV
DEREKk3E64qBcsW6dTEOBdRxtiaR7oAaSp4sRDWxvuRVNFcrnLwNWqQ1JQnQo0b4
8xXeiP9q9Wb9VrxtoHvyUJOWImDr/DGH1G/QipD/VWtU/shSUTO6/h8n1xw9lgsx
ye5PNZ6Lj6/BUIqZenyk7tKxsrbb/kbhbSJy9AuU8FNUfvXV6c/velsPOqaYAHCG
jWHJ4bXjGtMrrMHvmHZupjpsLU+yp5j5lkZOIMjcIafWFPtFoBrsrPPZnVc3nm/c
rgcocENaa02OSBlzAR3L+sF0vcBDnDzSVWv8l/w4bmWUD5Wy2I/8C6KcxjR6UqTX
3u4Oz4hp+p5VIBva9TodCO1EzosmGNKb/bTxUkqO1hcpim1LjIuFxw7BMiMfS7EZ
RBDmNjrbUu7Anb2x/In14DKnU9YwPiHVFyG5Q//X8gcO45mIE9QUz8xieUwPAj6K
ET02LJ4Qyfa3axHryQFIQmB0QGCxxTcHOkbYAuA6LKlPZcVG9D64ZIMebY92n3UT
1dgYvFHOA364mF7aHLFQkebO449BbV7dh1pG8fqfv7Mt9GLW4QEcjB0uha2b8IZJ
Vvn1QSTtbd9ofGWRJMuSjz54ayMUHJBeQhENqcTpQmJdpg9Fz6EY3rV1EFn7okVH
gGYcTaIarJD2Iz6MJzXAn7l+oIG1o5PUbH9qbxNBhFl3cm/fTOpLoy9w6n5jVO6W
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HRSnxCJMiWVXzp5nskq3M0WPO+LenHoLgtc1sUYvUe/TiovLv7sTS1sFN8C+PQGA
HTYt5jAa4rbx420Bp4vsOVaQKOOLgH4+UTgiY+puv/GFXdygC85jQ+oEXV/Mclj7
lTukqYct7zMAYMNk7z6mP5jPqHHrFCIpMz92Nl2Fue3Lz3P+ZZt83yI7VOm7Xyi3
ya2VxG/SIoNjRqPZHIabybk7uhzsw2iddFLTYF9hYy5GfdkAJmToZsqMyEiaBwrZ
zW8wPei8xGMhHwLXtPQM45uXDYrlkYG9/wgFJlJrwM69vjs6QP08akbtH28cowO4
bsoTJu6bmipSkEK9fzoNTw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14016 )
`pragma protect data_block
vrOw29Y876etu30Y4G6DAsdA8pCcHUWL+pQJu1CKi5/BGC6WTE8EXMiCyCEBZDVc
lSw9VUtVxGfbxsMwznCcYHGQd6GZ1ta1dcxQbbeZwhbt9adIbJrMDu71z3derbD9
KhDheDsL3B1Rj8Nbi4WjshsTFGRkiJNNAZi5B9GwXbiA1Xr+88tSNeI7TtR1EGY9
dLP8aD+UWv+lwrSB0Ye1jkfIyhjsp3WvQZMaLjbP4EsvhYTjaIwArtkg7Ai173MK
s0fpnLJzMlq5dzScU1H54bEfCU5113Vt+tDjm7wTNtsobLia6APeh9mmSOHX2E+E
8xt4MqN0zaCTIxdOPMl4/cSuSumzt8Pct72wG6P+IeSFGn/QBwD+k/JTOK3GsFku
0DEKUMzU6DjawIgya8F2qaVnd6RLGvhhOb40dCCiZRJzDLEFEqWevrLmO7pT7FHG
XgrK07mCgN99vR/4BzzzeylXbK6y7TVrXtsP2huSZ8a6ZYREKgLfq8LFaC2dq/Ch
7yu1pmrUFO6VDkFpWBbDPTP9yIaherTbGHrn/XYQ1cBKSfVF0Qvyz7N0VZGHrnTS
quYf6aIhN+GLvjKSWf71Wip0RiyOBgWwlKJuxynR63zEas94uulDKHvGSFsW+Pt3
pYs5xmsa+jUUcH/IyPjzCfjfO4gB3hdr2Rw/YjM1pik1GG6pRzRhkOEH+RztChGF
vbnqWenYt3f3lEIFfinCWu9BpVAWcAJZnYNUxluf/BvSa1qXRqV2WYSnKpNIkDaB
gphlO9lJn9xvrN8nQ1vSjQMrpyKf3y6Ns68JI6pPuAOYFKOJP209m5XDgUu6ZTR4
VR4xbrpJOLebsqGPtXIuehRpagewuY1YerVjYGhDw4Er1s3k/gSmNnOS6wKeAMWg
AP24T4eFm1LcHdDGeusVBMEgFm3Pb3nSz9yLdDuPPh+P252UpTOoCpa53YT52dU1
CtnPwp1pNci0sBnqoJx3LX1LTP8D62pYAICkfboNC9HrRLJCUsvclN1U1vuy6HID
NkJTHO4whI3xxlhIp2n15UlKzqpU9NK+h4HWIYEEKKjzzPWSQh/McJgknDbMcuwl
+nMeB9MJS2oPUZ9SkYHl0jpJEgATcML3cc80vkY+TrqjtUj17sReFv656un6gxuq
Kamv6Uk/8h2tKUeJsyiihFyjLkUjhebIC/ygKPYJCX6iQ56EAiq1eAStVYsvhUOT
wkTG5cVshFUMVmjeFQcl7pzq2wrY7Cc0nfnxPBRgd3Y/U11GhzJhQY83wWbfKVxz
TGSZwAghX36iY8GAAEJgpNLb4wBrBHM8yZllo1JukxxZ0mgO3iJVBXRvRjbNY5uW
AJKqu8DNIIYwtB2ggosSf5FKftP0UBOosjSni/oBn0PDi9uSCyT4O/mRhCcHjcPi
PnZytm3eTBSDeuCCgNoNz/NmcbzgSb1EjFge4VbTLa9Amaz/ELfQBn79MtQ4cXyM
yL/BmKJzeDgwqyf78u22NND6ZjFN8YzUw+79cbQ5CYVypMcnAfzZy8oS/oOVoRxx
VvTkHe/o6VqG2jESn1JfM6JQ85YYDXmbC/qmBXuviZvnheNvE7Uw26j4hUsNOjPk
lFE7Y0bWlVjq6s8kWebeDDtn7JCBvq4p6i7i9Z+Lc+Y8ZS/3JPaEXFxZ61xNOP/J
l0zzA4OJMDiECMfXFTRHMCetGVDZwEyQ7NpoW6vN3LNnUJXXwmqQIqQUkxWiNHuN
vAGzXL+mQwUb7fkjtHkE7W8Q6Vie3EC9j5PMi7eqUt+IJj8ZTomd3hxNj4YDc3Cx
LqzTFUxCRCZXOtNCy7Vdt+yuzxJNz7+GZAmhAf3wtt6wHS0Xl0Y7d4MdsuKC8ER4
YJmGkGSS6VdWiKoXie3XDRf49Wd6Qx8VOem0zxW9VANEB1RqYBmIKTn9P3K2SLm5
QPxxkI3tK6FlTqwW9JG/AphKmdFm5QOI9gwgJO2anDFNm2Hye/N64eO0EWu8lE8u
fw2iC5xF4sFX9MvanGaIf3pP9tBl7VW839l/H+YO21/aMp8f1t3sHifU4ea/gmtB
1xvLZNb/RjjaZ+j5q+mVxcCnQoazhNSac0xTrBfplSy5+cL8I8CC/IdZHt/Hg8bR
JDCGLs88CV5Ug/1PIS4wODcq2DxT3o3lenO3/CA8sziClX0Xtq7qowp5H2uKNW6S
r63tvGmJTQuTFacw/qTrMcuVnomfvUbWiMslikg3NxkDWN2ZYf0Fazn49bHXBDot
uAQXZgsmbZdf8fNNmVwviOcIeMp6+CHG7QoHY8f+AHC0VWXiFgwmYgOOGWi5EIEb
ZtACimf8DCFy5XoFpxkHbGkc/PqIwOzHDGD7KlvMUVBesr7+X+EuyemQWSH8G1OK
LoPbLIjdTVMd2liyyKDNQHhCjK81k5HS9B5RXhgVBeYCMfrhpOTF8I5TL5V+GbOv
gB3J7f4zi3cUD/kZZedOmxgcfXPjxTpUqo3JC4dVlyRBPRyE7vI9hozy7XPxBea+
rUMRiNibXgqLnE9wYzCEPbZPNFwnyw2rg/9kRa6lH/jt9AWiHBpWGOmcZoKvvsIW
IRPtuXd04R2TZbq7BgEzr19ZBM5bwgqVhI0RKPxULOTq5YF2wGb9EvEyU/AyiciG
2Tumuqg59WVo86PkoT0Dv3JYCdiPkdkB/oJjliT1M8ob+jqa08bDbWn4tSxOQu4z
vBPj7wbVd1K5TSvT7XnKMe3SaeqjeHGD9hNqeJhB4sIJCNx2UGpOHyMuYrcTJuCv
FxSiQVJh1R8WwuWlEYLsJ6IQ7fLnO1uabFDY1EtbsHjfe5I95WN5ioNZAppPCCf+
/16Q8UGOerHCeqvxonhR3QC5+FKU8twcCbTe7WdR4xnfLnsS/Wd+kLoRT3qnPUbK
0yoF9C2vNqc5uRxuio03qXTizkBg9DctVkeUwYlxIYxtlmKWktDsf2CJLGssAoyZ
wXZnR4hgcclf3zS8zOV3c+Rqlhpumbt4VAMOnuMOvj/xiiiqPWJ9lmwCSqNVIFFE
6KVmXIcj7e6a/JMwFbRxDw72U03fCu5cm2GXeXpmMA29hss8uxNR9QPPz9C6lW3y
YC01pX9Gch0UJaaN+Ewf0qirEp6naXHudJ0+2wlA/rqoSmq2Vm0kdNHesxTlUubj
RqUXSGDyi3a8tMvuNP7XtLGg6SPfcQXZRNuft0HTRjyrTGbK3Th+cI/Jg2yDmNRU
gfAOTQLYS8vqqXEYR9EjnJN8SR9+Fsj8Qr6BgZSReuBOGDWmaUvzwQE9KgCfR7j4
Qpe9Ea/H8eIl25srWDZsZJgfUqdG1/F57LNMhP2gmhBJGA79+qB3LKsVu+Uihc+G
lVnXYDbWZnOmi+C38pUROW5mKrUi6vZH3XDkoXi1vAqwnGmYQ2ND+GK37wHkY530
QA+p8ex/RJRc2HehXB7P6WKfvFF0dvKH8zL77V8/G7PuRsCkrs5h6ZKChj9ZZx0y
RgUpiLe9A/R+42eu6JrxET3i49dGcNP4x1y35Pv/KeQcABrw/zwo3EwmwIdZn91e
K9cllHcMR+j+ldkCMwu7dEsna83Bhojo9JzzXrh6Nb5q0zA9WLjmG5SSHvcvQ2Mh
wLeTgY3FyBhrvxz9s/lLYq8+TqnCdR9n/FUp1nHX5mLyqC+Yh40qzizRFddj4cmB
APZTvkUsWpUZbAcJPpGdtAW3jMI7i9aC5FuKUlkzBCo5vBgMFAFUz5SuVFL3omGL
Ry7O7wh2p/orbtUqUSfEHVjTcylC8yoqabDs1LbTwWV4qAjb53GzzQyl5EU7Q18o
s3Os6OlpYVk0CIwRz4qHd73bxDT4ulCtl5lHBv0uqFMaeJQdX0+Raj9JdaLRwLTS
bFu1zAnafgQMAApY2wyKJeNhojLfNxKprn+m37o4xhSjKtxBc4Qhm28we9eg4flW
Jd+MmZf4v0qUdfbFrc/dqHQi9D/eAtnbfSJlhhqfDqpBRmexYLPzZUagcvgJhTHe
5HZx19avfHhcFGPJmy6kymnXbquKsmJQK38NOup4af8sra6EYchWtQkIr/p3Xsj5
cC444VKBCK5WtiGQqeOgqhx/y3z8mBpbqLhQn1txC3V0whsARjug7n9cADESLYLL
dXIvEIMH4jl95dayIJcFpzpEGHCLihvKJbHDBDsQRzZLOih/Zw1vqbYe9lMEKxuL
eAXOWjEldqqe22UdTxgix2a7C51Hs/19l0k0EO+hXuvO6O4uLogn83PsCtKFeyvY
2TVAw5sR0uHDD43tqENlSj/O5PRkdzoJDAZekLxq6ERp8C2S9mzpze1uvagWeTU4
3dsazsgfADQgn9l+YlwoWtsQOwvYwOvIo39kjTacOoOniRHMIzpX4nrUDKMGTRYq
qgwbdIfqi32cS3Zh9tshu3iBrAtbv1il1pmaE19WbxCbAPJS5n7hRCX6rXf1cFxD
qV87BWcntLywuifIuptIIlW0j93lw7xGSPwQLl0XbhFvqeX2BilVU4W9sKuujkBL
/ZlqKDA1jz7e9FyeLyNf6AujX08+AQdehDyGUIoLI3QK+6tHWqBcF93prL5eWWQI
xvsCKwmo3f795lSOCzucohcIPnAzbBv9qWahMIV9GlBaVFSFdc2jIB0fU4dwgVTE
jUNva6DD1jVNq2hneqbgXu03dbJ9HbHbKD9BtTdRAdQnPgA9/VrH/w77cf6u0CDn
lA6RsLsTYJC/esFiA+iAyu/6pvl17Kzl5vGca05CwlA72a8L3lLNfI9HAtFmGFMp
ZCy+tmUAQV0Tp0kdmeyjq2byQXoN3phtWYn5h8oTLMOlCGSOcTzXLDwJO5g0CBx+
N/XZfQ+eOJDI5viUInMqVGIgWbQUbH9u4JdusSip49K/B7Jn3Zt9RU+KbgXNO96g
XcS8mDYhKRklhscHw+ePORuVksQBNeiCsxYUSYJYe3FTPMB8E6Hb+F9vm6umlg2V
8BAqgmpq32WmCuk0Sy2YuY3u0UtC4aR6CWwZaZG9o7NueHRe046rbdr99r/Iikq6
RVWKthvc7bqisEW8SPhN4DvZo0GwKvDjqF07o3ImCo1zfoCWKvZ/FK8CHCaOD8AB
YR3BG+PqBAR1Fl4uQpdaCHISHyR1hTIljfuRkukDdZ4POpHS0TuH3/FWYd3r6oWz
XyvR1+Yzl0dHDtQwKZ2mpH5H/V8FWKNBdFG1kAefmM8i/CvuMMBiBWH6nDyGkJx7
Ss/zfnAi5JyXrB2Qgr/bn12Hrt9iW0aa+u7kFv7X27dT1V5g/sxkvU2LVp5rfkD8
SiQFzaOWlvy0bOO4+ih4i0PPDZTL/IBUdVPod2KSRmx4qTHGx7ex86WIZnIVHLoO
Zc6qWNn13iCK1U6ubnuTnNPt5Mg9yVfgmhrfPdcm/cSO/xai74bvFpqJB567I0fL
IkIePz4SOJE81Kc7/6sPURA9DlPHx4Wq3LdSQ2zrKccvVYbMkXY40I3a1ujana8I
b+FuUadGATX+hDqtykJFhOxgSyXxanhVtXaz8bO6avwcZJZE/kIDYu0QuVOAwAxn
ree9esStzIiH2J2l/eNPE/DziU7nfuFr73jS/fbfkRVPoFNMrd/0Dl6DT/BzioCv
kQyeATa/YTmTfGl54MP7dD3lWCFqHbiCL+5A/N4Ne6k1Hi3YUNKqemB4xwKb3kbC
940TKMGJj6nqtVvjChfT4pP5G5H5PIFhX4NLjFn0ZMtCmk2LGYjLZzWSqbLtOLDy
VHYj2abeb5Qh8icKu+RZuj1uVYal5jLgeUQthFVW9IdtvjnUpzIOe9unCs6Czlil
oijIC6GgnTm5WU46Se7oX9Wa4Y5ogPUg6sAZcXaZF/oDt1rzVZQWB+XonYZHFZGH
w9rLUskHclu/GVhsvBueUfJrBvLA3AGnNOO/q/otMMplc9Waaf+PJjrypRCFlxN3
UdG/Tb3AuY2IhnMPHSYUj9EwPs/BH0wW/WcbnMnoeku6HE+xOVstO5iK/Tk90rxY
CgbLLsF0siqbop2Xkf51qwj151G0WPuHZkoXo2EbbKMrcXVbnxmXSQZ5yOuikWo2
KCx1haNLL1j3XnaXxLtKCLNiSy9FyNJHCw+ZWxM1EQzj/wxOg21em39VoQ9MfxTl
UWAarKGvquAknfN77AhkuaS6WcZ4gOIQwR1Qo44IURJIka5yBkRVQqlcxXOX+gFx
B3JCphARZ3GrSDbPtew5hcwszegmGNJagW7qhJMWBzWj83bNGz34aZEgY4Yy0xv8
bY10kvANd0nhTZX7SOVgByXEUJtIdKloPovZkEbALbInPm59Ri/MYh2hx2+XfCUz
r0nxF6hBshdF33u76eE5ZxYeenkESpYqXiopVfEX5fEdMM3Z5SDmnZpvISs/qdkZ
XbM7x6d7iRsx50wHOc+6Fdp9llOIborrT88ZR6N8jltnptkFhnpoeroZoz7Xi+8m
ztomqRACZ1rgdyKxVegqfPH96YdlR6p0MW2Gmk1BOMKCad44zfmyrMdAo3ZCSHoi
4TJLVO0VbWOaHQDL48PzjzeN5EehxP7MNSKFLq8gTFBwozITr3F7d7+zF+FtX64u
cS1VCcBxDBt+/CU+8ETD2UaH0JfRHBOfJT6+0bx2mB9QKVAAyD5A3AwHcf8ZfDBz
gdqxdDwSKRidTjIT2FWQ32J5XM/inn9zpUldgybPzzgc5D9S9Bv5n94RsragMgd4
LL7cYfXnyfTngh0LemGx5KaEb6gaqsnQ2YyfKwApM9zlEfnAX1IVQcm/9Q8yggKe
vvI84zwGemNYnq4FuPpe/QtNXSIBbNC+QA+6BaOfRkdoV2feLzf81qpewopS0TnT
mlqUZD8a/eVBfRaxe0SCZZOZk+g7ya5hDySBxNsypcI2GNPTPGzg+UIPSv41Nhj5
hakpbGwUnYpzJc1UPO0BHkTycTjeV/OamL+ANc271Rp3M1mOk7YZA+LQ7+t6rqpb
0yLlykA0WrGsYy89v2aWgfDTyysdoCAOdaLt1T8k+GqEutO0qgiscNS1rar2MuaD
LWe2OAkFV90e3sojALUHRP2mATC7otckCmnbUkhgbbLcUnaom5spEsZjg0/UeU9q
KzODNo/BRxAmVNEsSYI7/iPKyIp2/ueuGKTMwBmJpsKw0ZUUbKnBYxrQS+YeBVv6
MmNoTiQvOkF3OzBZWYkFK/0vzVroD5nrIsoh4TQdNTd6sWyjC5ZKKOURFFTdokph
Z1NuN8t5xhLnDFaJ2Zoc6quBGNQu3+evdnGea5/p0OpGVgqY1f5Dc3aTd7AeVEub
o61FvpyMH3Ht+Wz5fzbCLS2m9kSmDKPCvirU2e3wP56P01etFEMUSRNDVjJxURBP
nWQHqmTVhDlDqF9IPenTO61/o287rt7KqC82nFFni6+PlnmNwumzwwKKLBg8ud/T
IaOHKeSbhIvpWcPMgeNaQpy4z+y1yuGhLpSF1ijNY10gkblTcLjKPtjyYNEDLtwk
f7ldsCV1LkwSVBzdmAHLZQm6AfRcFqOhXnBnuipgKTKWoxPO+GaL+gXUW+bZa4ko
FY2fXkGnuQDVpawrHTsR6VgFHymSOhkNBSy0MGYa26hp+13wzG27W0Acsx/vqz9b
ZHtQwMrvt1zgTSV56K82h8zaU4fp+97QjLnihZyOmoYEuBHFJ1q40oyNtBQ/t7b/
p/N1Pyz/L5ACxBtezjg07xbU+rNCOc9JpnvrJOKV3mV5pCTkMZ4u3g6f4BAdlcTB
fJgLnRFBRdS4domyDvGL0LPvt5iIp4TAuJBpvTABtuGRiRgCxVnO3V5i/HsniSLq
0t+pNsOPAsDKPin+SwJRV4a0bmV3xWM30FpM8QKBOQ+R4AV2ugj/779FBvVtURfh
nLwgwIxacBkDTw7LWaT4yP5+7QdBf/Ah+pplEbl7zmOhcHdnPcEUXEMg38/Ksk/2
INuUzZw7j6Zs7ucio4mpD0mO8x+M7HZYq7ypwbmIFP/533cwIbg1Mydg8RKaomZ+
3fGxiUtO1Wjtyxu1Mcc5BLw72ag+mS4FsloCATdmEt1VYKOcbKmjOfhpkpmL0FK6
/Ft474daBFyEUZ+uw+9zwKFxCWHarQ/jLUJGgiflDjCxbwJO4i7kV8Mblk40J/Xq
v+icZS1dNbL3JNL9+IbO3AFmbhOM4CmBJe11oZIwflv0CucHu1OnuaHUvAahYUE0
eP9LW5LomZFJrMfz1HBh55iOvnUrkkIWDiJeR5tpi8LChj9KbOMUadmiizy+wLFP
UAj+qkgAGpY/SJM7CR2sEWGWwxfQa1MJUwIBfyXw3PTJ3bTcZWmfrLijDplMxSIW
f+UjTsIr5P5ZIyrMj6DT446fOh6oGme9jNw7DtgNkUakYGC6dFJS8QpRdjhQNT3B
Gf0zN0SGEdAuPbdk5jmyIEsn8HsDgVRWC2PuxdPAc394wpbha7bVh7y9rV/vOW4g
0ydLofMjrQTRqRqBzqIqy+wM4z+l6uRv9kgbtifotY6Y/QdVcLK2gMZGznR744TY
FooCo2ydR/HPyBqV1MSOhke3tfawJTWlxJZDRhZCa9247l7eyNkRmIidP+a4amtn
gJsgCVfGkCGQWdENNyna/Z9hf0PT91qOV5zeEQaaTV6dmKtb3SBG+r+DcLXWJksG
9+ExVngNnxXzPs+VK0Gp6Py5VoXwI2hmC8Gs/5QgOdu79v0o1h0/RRD8zfNGmkEP
dfhC21SgtreGtAzrb1dsD5bXRcf83QKrVG8GCjiuXJUoAf3tTLrO56NUp8up7nu+
OjaMYlte564NFuJzYBH+kybtNOYvYMXpycdvNa3JI6cDVHeDWZ3Bb5VuUZ5lT91/
UZyAaz00S77CrTT2QzJd9K62ieR5bKNyILtoWUz+pu91o1rSNiuDdTQjA+VkYH0o
ityER6zFW8JZp3zsLOCnofx1kStQVoxoN3+DIpGU0sX6QRCF+h9gu0j286YSNbrH
F/i6wB7dlBxyH8gAm3c5VTYjWezEcNN6mg5UTCax8J1aFY4M62mUjBDpylzkMP0q
2GjDyHao/iM9yiiYVu7dlc6kefDB7wmims0mBgozM1CDBkvGE/qQqQrerePIihD1
bA/Yq4BDaUDsbCQfTC9FDrUCKlJjdppIIkPH48IjQXXwbGm9lNNwME/GmcHWlFuU
MPZR2s2N7mY4sqMuXBcnnZ+2KRV7gfAzGr7oWGBNNuBKjIurebkOHd+pxdkbflKY
KtXurdlesSouW/dlMSmbsNTC6IeLOjtW/p1baLW1ud+fAqJb4rUWdZW+Z4+j6urr
33/utXttpdcI3iVWjXHgG+KJOKCPFd6U4mrCVO1nFdaY/zJLai0he/z+r067tRU9
vFm0XHzR6o+5lAzpQSfte/wdQ5IzOpyqTJjz5qFVuxBMIl/aIL4pe1Z3Qtz1D31g
S4lpN2p3l6Xg6jOkgdF8Ae5qqnN/6D9Oit0GnIVLqcMN7t93q+7jhPGTqgTmktSb
4QsTI40glaqbAceXYGYiyRpKKXW1AXbh/TBkgfVsBO3juanCLsL1uFeiPqA/brgx
xQuDNDy5sBEpjRWILYITIjW+rcjOSHrH0RKPwOnNuo4qGW3owZ8hWRtUTLlMYqOf
dC8xmeonw60vx8g4pNbdjePuY5K9yfdzXHp84Kq2pNSF9TuEwMNviwlSGdaUMAHb
LVDieiHgTz75JOEhV2cZb7aM4HZScZNwSjduPhAKcGlUp1mrZCOxVUddETe4Tbsp
chjFqT/WfvHFhtdfZayWMr90+pFMu1VpXxxCRM6cNuI2dU5wAVsmEFaRtknSAHHb
MUX8aQJbxyPCCTwYRExhCzJ2HgP7rluWymEfxoaqHZ4OehJId7/vBTynMvCzX9Jo
R2mAQkDjssoYS2yqhD4HdefBagD85dKbbNDw2cwdAybYUfEzSXqK1PJOdbESRVj8
Uq4XgqOSDKQvc8dFzuproRQDYq0B6EHOBpMcKWbaWR4wyZt2Xk9rthY6YnmQj+yi
vEv5MkgfyP8GFo9ecp3iEuHiI8LND1i2ZcxRMqwqNt1l1d79Q1iXm8CaMoSf9jR8
J2fJb+IupL3xMpnV9f9ckFN90TRgQxoshBlzBBiF7IYUTy7juV/BjTx3N9xqkQyT
r5DI3va29iPqqyX2HPLslLjN/+H2ZMh6wA9Lsp3T9IXLNWZJXg2Z+KpFxQQxPvYX
nTeIlEy7HfSBOUsKdRQyNQObSQ4iEPzF6gaOlY4Dcu68MqjfzQk1P7dKJU8sU+Gp
v2aWVZpYAU1UVopp8C95WMzRA+K8Ab6jQLOsMWc8MuwljfpiTr5eR4UGQN8ytbUL
ATmsSIb7dSoQqy6Q3b7+gbSLtndjD4eQjzvSJYygdJq00o9c2zJLiy8FbalDtKo7
+QzooSVj0HRWIxkgvZ3RIX98lPKLP7/Mdkh9p0lUwB645FNgAYnINKCzoY6ozvtE
cTMzbl2jQNb8dbSzXUUnDpu28j13dUlPBpy3dRWzIu8YubBS9O9OEG/++zNToN7E
+u9oVvasPvBSv+gfOs+PONJcT6WrzADgyec2g9yrDSkS+Xq1/ilkBQxF3LPS7hBY
/gfPmPLMiAb9Mit22ba0rXlQ+J+82KXeboyXHqwIugytKdjZtFs3HhhNlyfEHq5d
nf69c/u6n19i01QSo0CQ5FbfRhGpDBcJiu1rjzNR+EGodNU4D8QCQCO7toSkb8PR
94KOITHC79dcHJqeT7tN35Zcyl2mirC1MLGKJwTNAuG7DzujuFKi/BGwhGVHPhkO
YaDPkaxBT7cUM1petmuI4Owmn0TqanDUWXv15XbYCJRKVeMrINWs+T+9aT95GAq8
UoYoeBAIrBh9czJIfaKdS+vnURFQ6pfa5lt8saj4LfWFqKx6gZDy7w7jygoyehra
4MjbRJzDqVRGvIJJAAOkyMwlJdSbfosfmE1ULN2OhtBwDysGulbiU+XX3eIPdPqz
pO8qLY1kU21QGD+ycO+KNcQBdxWyUCVA8DoV2h0K1fHVSv6Ix4kRfEvmKI+Qw1O4
8vaWfmJ78y+WxXmYaRX8BzotLok1Utb0LZpsQIlB0JB/7gPzbSxMFo3QLIYISFrW
y8+bBJcALkkxo7F8iFq63lPtJGXATHYtj/HP9gAa/hGMSR/wEe55M7wyfIIUUdew
AWzXzMGAIoMt5l+c5jPGEtbAgO1DzWKC8KDk4Kp/1yllJ0jpVUdkh5aRtsYqwPUT
rcbWkJxeTYbe76sxDWO8OOB+i/sTfOtdM9rmEMdAYwoX7pzbOhIlbCmXSRQ4CUqR
XOtNNFmLfvRsSd0vAxU7cqBltCApkKr9HgDzBe7151jarb1e0cn84zNhvc10gukU
64MHNVZa7Yui314AhAwzfhUfL/fB4ERLaOwBfiIpjM8OyNzRjsSgjKbNJ6eC/s/X
IJCawTziVQGrsyVXZAxEylHOp4xMZvcjqwg4RpPirCc2yFtvUmMFnXmd7N08SKeW
tfNw/OPw01HNid4LsQcTpPr4ikMrC4tYfWy8M/KWAxz24ppvz3xq34c5CN+qxJI4
1iTJY52s3xs0M8tThyA1OIGTeMHnkeTBsO7fva+VUdhxiVk8SFeHbJ7ONJWxTbyk
FAteKbA5qPCidS41kqzuAIQ+Hjv1oUqhySSP5O68F4zMoH6buMH9Rmg8fc7RkyFD
5cBjk0r5wKlJe5hA72AkowXun3KK5aNRgqqXfyK3qbEmjlU9CQO2XV4ZPIeqZYak
No3wSntd2g6Afe3mzw175m5juFXqZQCT6eQvDUbwliAyC/Zp6n1iclJjOxBtpzuq
/WJq4QccxTZD+tsbOTYEkLF/bb00Bd+KoCzc/GFLBA8xiXKsQAPUYA1RwIOUc657
UtStjBWckLuCSczHIUHiqXYUcHBNmWDwyZyTFcOrRwvoSQv7dEIx77+A2+L3WFqJ
QdHV36kzhNMk7tyFIn7T4CPpL814ufLO0cJcr7w9N2HfUxPZPJjHF3i3F8ahhEjn
wDY4Y2DXf3RaYVYaTEWwyNxPsqzHOv6U3MXyCHbCyOsG93GWTYULCZ0ffQlsAlZg
ZMxAuEnplHXF5cimlNwGKOBc6l9RNAHFMiAcRylnX/3el69o1XJbAA6jDfyXsN2h
SftMG1NcE+o/uVdZ/HxuekDwGMNIyf6Tqm/j41W4O1U2e3T78Hil7A1qahKDK6iN
e7yj9abSONJceis6wkixAa6ycAfFjVG6/gyLC56JcFRs5s1YhsMy25Eyt5XXxUDq
xJ3WqYolKURduhhY9gIqhULoEIsYQV3K9OP+sWK0P6r3ayOJE/QomfSrsKNctMwZ
rspoAP+XQZlvSRD6oBdUGvY8AowFXcMit68RAXc4DzaCCqiU8mQjPOiwpZYNACk3
1LgbC1LkAE6JkCIMTKqAG3g0Q+FY5ZbiDvCEoAUbbtKeSTQZtImLbatHggANR60s
TLk3Kepzl2n4BHkCADDbx61BeCOFIBpLwvdDUoHbj4vy8zam5dLfy2UIZG0cVi0O
rOGJ0C8yOaGCBJLgVDpJE743xHTwaZcQ/hdKd/mvX/jbbXlcWz/8MI+nY/CF8Oym
78F0gl24qUBnM8kwhGEsai0N0ZgmwWlqM92H+Bpb3mTILMEJqVd8A5XQdA/igKAL
z0CGpIgLl/8EknDp9gt6tVKzCNnPD7ISSN3RURrTv+NWMcrBlykp5n8tc3KZwiH1
Resw8mTwwZwhXlxP3J3FpId8uH97OmuQ6OtIYAw73MDTSKjbOvIux+f+IGo0/qA0
BHtW+gRAOFDpaJS2f8NLnRUW45Ui9Q+43W6VOZt44v4qjFDWyuc0Eczlz6NEOpyk
97gJdguCSW0AtmgfnqS6BqNFMkjMm/Gl5/ry5P7CdVeZP4rGCUoLi/4Zk0DkgYm/
opylNVHTMhArWIAUH0fwV0rMu1+3SlmA/Kspp/rfbU1Xyzu5uquK5B+L0A582WEs
YR2uqTrOCiTDYwhv3A72/9nhz05t4MRdNa9jVJZ2RZKxuJmRXo7aI6/60uRlyQSZ
yNm9mjPDnvX/Fz0Drbq5XdQOuzppuSj89OOKKOzgZfnvgWthxgU4/XEkMr4VCm7h
pSIKBl/OHalKL2wsDgFDWeKEFtL48i5Ln7IiaUSjdAWxgjCBQEpQYNPa9FM7KnKr
iyyzVrmOwX7sPY/SzLmYTDZpQd/Hvz9Hwa7LwfZV7zEqSBBSVsYlpkEapE9mQN58
u345HoBXq0ZT+WXVTZZFcQ7WGPZbHZba2bZyeCoplf/KHI2V6lwPTuS1v/36/5DW
L4YxEQ7Jipvfdo8GTWLx98wjvIODpS8ojiRg03KpybbOUmXCx/bUU09p4d/ffPEv
NYUChwXsE/zru9AaK6noRwR3dYz9xu4OFinxqoeNM0o+yBrpWsRXbQ4R/zgf2w3P
2o6reVrvopmboue6P3VZ0EeeDjAaA1kFgDhoWJTNVY9uD7Wq7HdjYF3QylIOUHkT
UlC6kKY3nrYridGNADwMWSk3noohgV3GMLJkclL8BHlEYJyRJh+Yi5UxWX+iq/vp
NVMLgiKpvicnsnkrT25w9yd6MQZXWoD1QWrXGjtr4pn1AG+i0mDsVtiLNu22DIyc
hma82GDMLWpIQ4Slcj+Kouf6BCOEGnMf/s9wZj9e8+0gVS+p4tQ3u3uMkIRF2QNw
ecSiyu1NJciXI0UQj7azdHCUagxp99NiHqUMH1JklmOpXTsueFn6Y4oelX0u2daz
tqLZMqa6Ot7rvl/1DqW0kUdkiHD9GVNG7UG/qAvTZ2WpVsDvErK1WUp2rCcrI2jh
te4F97T3s+ppjyYgTmzKtNMYT8Urv5mzUkRjNSja3gaBoUgmfV4StV3r2VioLXj1
AsFpcFiRH47Pro2MmHPuyuCji8qYuqNzVtfkJnN9hdUXHYZMLF9eh0saCNEaOALO
vk83hxt4JTQHvSXrWf/mjbfVrJP9in4gB1JNMR8T/xtqUHEtjIvwezSw/ZEnRjXE
Yvz5jgh8/ghEcYDuxrOtRqxezzHuB+pHegrYxHPLd8emHJnxJTeWsEd/rUj9hADG
LulfV1LwfHzEWeHKMi3j5rh/S7OrHSlhykfR1REv3IxOAtP/zSzpyMGdTdbBRl6p
JDGmVro/vXqpSax9R4pV8HimFMgAP1WZglyPbAPQnk/PE/hQWl1mKXhwWEsa7F1+
udw37psSwH0mwdM7sFFUm3a7xpXd9AEHxKTyvcloMLEHPk1zlbpXI2j4LmG+I7M2
0HgQmV6W/f6bADgB2uFl06XU3+BlxrdkAEd+DEmmacVwz3xgr2dpKqngXFCyiIgz
f/UPmsMb0LLJKfM5V5RurhmAxExRzYNWdVFEYfViL8WBPaEsVqHiY9VcmwyDRHm9
CDmd3b6oeJ3QRSTAqxpAgxMbjBXXANbC8hGEfPY0MGVbNNpDfo1D0DvmskAsR0Fb
+uxdBNOTz4W4ePM6pufSX/cmOLLp5QewwNSWErilZFH24erhgVujuaQT9yAkRrW1
nz+sLBoql8gDce60zwlfwd3ezwVP8QeQtLW0xQGP2jX02teNnvpn6Ic/gjvi7M4+
YBDzBC5TsVIpoSU0I1xykXeinVy8MdKGzFI0hK0Bf1/pfdo0pk57wa5QklmA+Hso
n0NoRN1A4dCFs0QOZRpBB8nfp+LJnPxT39SMT8qAOYweZE6PHqcGp/+FRxXDY2Vf
XKAUTgAs4aEbwLy+HVMI+wHGAOv/D1jcTxitYyU9+Yw9E1RcwMQ0rZKlK9l46p1p
F8k0i/9uz0E7e0jw0FfbRBFQK6bYAPrbss1CQStuUaVGZVvXISLnyimgwVynDOlh
0xWr/wdlpJmy7WM/tebpj7h6J4DKBHt+RSd+pr0R1VSHAJCjV7z3VFx4SRjFue9z
Idz1nFygo+f3EfOLliQJ1V0enILqXXIqmsA2iNRjMWW5JG1TBIteaUQptBdM3Qw+
2v9A2ticzKwfIFSVjWSD+pNxQQTb5qUhv0it2mgCc7Y9nY+5Q19ls7U2Ih1IIKlz
PfaxJt7j/VKowV/HoXtDuxeAMmLwApGMpkOFLyxnGsyoVp8kJFZSyHoUlQbyrED0
WC9jsENE5rX1NYvbctJq9M4zJJ16VH7yH24LYji7MyoI66yHpOuT/Pv4N8u9ZwrK
bXxYsPdKZgHVl3+K+EcL5C98akUy8nIAf22j9g6TOLPboQ6+mHOoHOX39BljV8vQ
rlMuaQg9baHO+JGKeJrpEdeLQQ1lUA1pRzZ8v0VObC7I4TUazl8y4z6o//S5R2TG
LC0kcOpVHxbJaUTy76x5qIyk1DZUj7dHZG7QzzygvaJD63cRKWw7vXPPQrtGFSOc
huT9G9YqL/aj+5FqrFpNqAq4AgQYZRdELzmudf7yamWyjuhhiYAKkJWeAnJHWjOp
d0qQY+wzRyz/PzJPvaO/ek0aM69pgP7U0Rf5ygeLx1SUc1B2JZ68Y2SPnBuFWeCa
fdtrWcDFwicvLEid4EzqrrRKYpeivkBxyiXNMA+54KIaPSjcYN/+lFeXTMmzYUfC
Tza0XCyVzh28uJNNIFgLKo9xPgDuxrYPI2KOrNy2+hyRqdDlQ5ixvL155oh8uPjn
z5aIIdPyyjVZnm4AeGtPH2g9BVcIaZ7WWb6gyZgMVePz4JJJtTUBQKMPq44YJNIJ
sTHqQ3ejc3fyrNz+dP2jPHPUgM9IDSYUU+1ngcQDhE/+hjX6qg014kUUr9ysCu2s
4JTDwmxkROmEAutDpkzxQHqm/x5CrKp70mZQBvNI1WvFTW3KGTMXDVjBBVcE0dri
SLsTeW+agjikUHCZ05D7rfA3km6gQLnI1+c5hT57xFk31p3Z87GhrK9NY87nc8x4
xj/CJtFQDMDoDkbdusAT20fsufE3ny3+RscgEfU73X7tP4dTrMA7ZTnRy0ySB5Jo
SUMiTeujKX2phs0fVMs5E0ja6631tWTPxcYNQCYnndRsNZlxnEEr0hFKvfgAi2fu
1lSPBljgr6Sy3d1npVyy8GDIlU4x7pwfKjjLEcJ3lh+BPVwehtKUYv3BLB/NBlag
9TuULv9dwJsDIY8ZOPjW+SNkjdyboDUeEXtIa/a9xs4/NUNQrMQ+WUje6zqTvOC9
v2TUEL2AQXXODkr0Q4dklDeBaNdjmiZUt05dH8ckjpB/DHRUwbxtBOsK9B+XKtjM
jTWxLvuxbw9vXHvMTaAkqyauUWCE8Fy6OdTOzhm7sMTgNmSV4Z8EHgR+34O6NKWz
lpC0xufW8pprLU4UId+n6FXvpROLP3hAJ6Dxx9pL3VJHVdsRXNZLLcn/+mQabfBD
shRod6vPnVFPMxrH0GM43ENWMA4yxXhmsBtL5rK8VNr9Ljv8pxgWERdsPvj5voA3
uY+TRD0h2sC5Q90d8RMwCPreBpV22WKOb7u3v5lvTzA5rMHWHoliIIrFzX8aUdeq
tCpIl66mDY0W2wo+cxiuKANI6QxoXel51pKoVGshcjAP3lUq/ZX5pK6JOtEw5jrf
kOTyTbtbCp0HQ7FR1S/WBBGl9S9pvIuYjrCgmxgx09PpWM/IC6LhnIqF3Uxf4l20
MDxVC2ADq0t03A5ptSYlhrfUjHV0E21zQF6mZONnOPUAtOqpHQft/8wcpI4ioAM7
J8zM7iYHl/6CE6YraZd9HgrRQTURVRlMviHGAJoYpiS2NNswHgMwmsRnOUth8R5D
YrqMa7PGR0xuLGGfjcz8V4xc4QdlnhSHSnl8JNxDcO1ltKAhC/SowExT1knZ448N
07UEexQeLiEoFZUBRbxsLTTQY3u6Bycz8xmVsdJsu04Lj6Ufgden72jHAHt3Y5Wi
0j7NVwhBlqR2LFj3/LUhMp+3FjQj6TIA0RLit/o/57+HlmsxeThhBzQUvpSgECWS
X3r8WPDbbwbNC/i7HwcDWA4dt95P4AxhELW2DLk+ayLVgn9pVUDuypR5bq8l5989
MzsTVAcKtsmZLsnqkElSg8wRCyhChTaM/XQqZQdYa5AFPBceqfqUtPgVOMhK912s
tA7ixRjY3Zs+itXk8Xzws3zeKag9QnYG3GVbf0mSkxFKR1VTvpbv5Ul/x5ok5fJM
m6xiw+dIpJff8eZvtThuUGG0+R9FTNgfIJiH92ADfwCRH+qnRJtH/CO6/EySEdD2
M4NNBY66YLLCcJOABcGInt3m4bYKUavuUwM3YUXeG0ezfRuC5vopQtAZQLtsBSRN
7l9ypzQolqXcZQZ/bbTBfacEXKcSS2VtHQXr3RHpB5sneI852wz/8+50/pAKF10L
pfhDGZ4cJXtBpC/8iJZ39NXDy0C4i8QapIlofusg0FSlZqvvlfwmLKUc7ZfNGzxe
6kNkeo51vhT+EJvbWs5ghI14MnXefm8Qkg1ecKMrcg77/gPhcibh8ui8Trgf3G7e
gbU6yGtQxCRlcGJqO9TEdnkkWQbE7Xy8FKLTjLmXDv7v6AoUzFTr0z65qwDBT8uZ
9TdXJLmO4Z2C4EQ/SVeb1K2NUdKi/XfdqQuvcP4ErzhmE3jRyCwcxSxaRGOVaotR
Y4c6Ns3H2tskpV3YsyNkBREuCF0ydWAPEmjArwI7I86CZQvA2A5LLPG4GuOatCF7
sxSXxGBz5uXOC56Ca9ZaLmOiGe/e5bkIAUHnndNvvUYUAJRC+r0tye7bclAtqXM+
Xt1GfQzFvL8FkCiiOnV7eD1L9Mbt3KsWrYnJipIJx9qzm4X2QeYqiu/bxJtI6Wy+
SDkHoyVruJerD6yP89FGDNgWi6nVpMwjFf4+Ykv7blg9s+CrqiwnoxyprhNrlJ4Y
DMOpTLbWCp49+/ADwOLjP6y13W0dmNY9pG94CA/vJJjfyPm+al/MEoJsH5xfsC0k
JYfBhktgo+/lkb+fIZ32Ny4Mhqd5GOuap6qhAhfNd+UwmoVA6j9ey33USeF3gFc2
Cym5HAE9erloao35nvMftoN2nC+C8CY6Ec54KXnFYng46u1lJ6wjtCSe291e8+SX
PvbEfjz9hoS6dJO/6Z23GlYrgLvaL3SJ6v+Ql5CibdVnGHf44nZEka6wd+MXvlmO
9CNjDOfx1eIKLbTvfRidebUUQFy9oqRh6MvEVgIlKWvIM5HgwLf84kHukskpsey6
Ywfi+QoqCSLVQHL7Lfh5plb/baseN4MRdWlJUxvytKohzlCGEqCu5UMfzzgQfIJv
NLht7MroFLfEr/rLgbek5NiNJgynnUmcJlsErosJX7jvieSV6+nleRREdBhy6jpR
Lea+3TyKBkqXNWNoBHT8ZFCG7DMwgSePv/BPPpfeHfqyDbveIGjGyn4gl2UezhOG
yIulhX8cJWezpeA0lWcNi2GAK9enrAmgglb8UfaijqZKFghYGJJvebYLFiIsYk+Y
pCK2SutbaV3QZuyhxNyVL4AxKpM1OceqJvuQ5FWy3CImuugEQUDRTv8blnf8ujfY
19PHkFAS1Ex4O26imc404jQO3K6eraIxtxxUTzFmuS0OxdfN3gbw0T7gV678Efzl
RhOelRWXdrqUQ1Po67Q7r5Gd5FbDMB0I03IH36nBATnGlXfauVhLNYXWXi5GXdyZ
Tv3M0w/UJa7i9hUgoBjE7700AMj5CT1eotPMQw2bEBNv0FMu8AbqFTJ2Qmb/hXmT
2hP0GQvhOJLKRwcXxRr2vrYuNgCw2ATSNTV5UHEEJwLDIAPqoBUCBW1uoaphsiA9
9SnaCqlbei9fGuwvB/yLQAYYIwM35P8MqG+l1QmnUf5PSyvlBeAd1xCzAg768Mfe
mSZ2mNlrBRAj0UwbtLnqwiEQcpGcs7MOfOv12HGw7WMxFdkGkTp3E6iDx1+yP47C
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
MbGsyjKKCW8JUuNHurJXdhvD7/6FyKLOLu/5A8kb5cjpmC9bh+9uRZm51qKmRB1A
ktZw9izBR0yhDqH2CGdvNyU0+yL+K8eeI6Wcn8WxDYMN2mB37NiZX8R1EuTHpn+T
u+lCX+aCD4besyS7OnF5Bg/teJGIGjvxb50TQowN/0hNkXJVWs+TsStLoKT7q954
5p1Vb76igc6OOLnK69D4FtAy/68srhiPkZT7BpCEAHEbrfGH9l4tj0GTowrBX+2x
Wed7/x7LIPTUyF6/rreMyF/mWmvJV6QHSVgdC5s3k9eZISSNxRFN2MHB1yDkqNcZ
MWNEj+9QHqge55ZBwgOUpA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9584 )
`pragma protect data_block
UN+4ts7e1klQpHiv03rCkuk0ef6+sNRrhSgmtiO1BKLQqZzW7K4X1AU2FeYOGQoA
NmMDgUQB0lWNkLk6fjiGqKzIE2JhtJS3MedHdeamQQR9715zatdaCC9eWyheDLdc
2NKtnVAtgUDuIxR5Fe0qo3u4J05Ecst5itTzI+sLY3y30pf69mKskENXtXJ9Mmp2
S8e7ct3due/TFoYkRnTV56T9Sal6uy83iwkQJe2pdPebbhkhVvQ4WKDHQPxJDORz
bxAgliR9yBIoU+j8PjxPbRo64mQcVwfy1Coee8qrEZs6x1j0egJMBlwrAna3ezh1
fXY2be0J9zONJ2hQ3mdgT6FKJpvvXd084hH5CmpwS2qo0CVzr/s5nbNwQZEVIB54
ndHOrAICntzzzW0UJDkkuvDboO3VNHRqdRrfxMpsKvkHpv69CFBVn55OhkUlVANo
zEzujjGaISlGSRFgB+c9oEBAQ2Nl6XCtlv3uDj/fZetS2J7XUhTgyQs4cabbC89A
tZNUvrqvH0U4v+T8fUnDFrw1vDGDT7PIJW09OzpgMynIETQJXzJvP76VSyvQoqnT
ACRHIRBpwqvC761o8IXaj5elPI1r9CucejeAU18NRwUsLbuUfzMgJA511D6cTjGf
R1gxw6eA1F/aVA0xrfKkS/PK1MNh77tNZbnunC1LRAsQP5uXtqMYeDOJ7qnvL/Hb
JZiieDWkudi/TXFknACOzeNRQk8HGUbpKyYGCEp5lWY4c+v9c38YvvWsAClD8jIo
7NO1AgDlZBU7qtfORPmHOJXDRn0uHFF/+nCpq48lEeAiuQpJZMf+vENxgILwu7mI
nw5kxkeCwmrSWIpdltpIutVKlIiYzYp0LPxyKgeza0Y7rr7Uf6UuwW2VGBmySjWt
YOYIdxFSbqAZjad5UXhDoZe4r20spd+3hHrPo24HvUXNVyVNc2Lor244LLgNCpzv
DG95Tf/yVddm7dITPNzi0WKubAG9uJSlzuXssTZ6PiDt/mjjyZLGUH8RemLpz6dK
tUlr6qvZghCdBzg64zDSdaTr3wsQ4DQt3q7NDqLTBBpY3UfaIGZl20Z7o1zqz4gL
dqFNkyc06lsmHrM1+r2cnvD1k/U1fz/rjAOTwr401HOWNBxyKrqq4KWCf3wLYsWC
U34JLQxi58Ki5/pR9cqyLikg4LUjfXoAq2Mghr+aYqaUjU2aykSNvA1yXp6QY0Zd
Pipb2RJe1iYx2VV7IhVhp6DAnm1TjJY/KlfN98+Qq6QfVtuhEnlJICPz6Fhd1zHl
mKP/rRqajVt+wbxaqubUKsqYUynU67rJQz3fpgMs7eXuIh36fbDuKxuwh43FZZTk
JIpC1jkcCycO0A7btGpPrZmCIz67XhkCPb5XnQ51YOHc3giXZHg+xuOms+8GIZsG
dKFpGw5QM30DZcVeJH9MjiknvzpFdEIQqgohPBWozfODlwqDk49ZQZH/FM1YgdOa
AOi3lxUOEP2WJWVMzoS2R4snfRFZZQ1ThZfhFFaMYIx5P1RxH/WeIqMpmW8SyV+a
sNLtc2BblV8ATXxhLAJpgW3RByvxCvcUzLSQAWglA+kijLb50LdrvwgWgyRNkTg2
uTMkvmDXJAenPsQxY7S4CjaEaF9+Ox9CTDHpEnKCXD5dAhEYhGsAnYWI8HGSPZQA
uZn+buAd6in4azxitQj1zGMN110OEUdbxobavJOrizMmBBPl8pBi/UWDxJ4R+miN
0tT3eHbaErm5O/3cPlYr3FXhb/OzrT0EI4H/QuaX71takBoju3+VdCsmoUPk5TW2
Y1ciLjFHApGFKnJd1lIPixQbNfvCiRKvYKFQaQKLXHtUONpXPIGEblcKbFZuHWGL
BZKi/SjK3ym9uFEaNsnEGqoMKHg0kxsgE/MO0OqaW8kvnMS/eYLHdh+MUteJU1G2
nXOcGxAaeLMySWkkdTmyBKxW4cw5BsiaX1esdgGT2ZibooWReBFphVkb28kZr5FD
2RVHW5Qg3ANSCAJpX7ebVVb+LYVFXqeUlD8CSkdhYkq4/M/2xgZ9pFWz3HL5zqJw
eV6OB1y+CGQq1iYY/1r7M2I7VLPyhUO78Q4umGz4oHK3fW+TRIHXogwOpRdif/6h
E9/gkgIfb/Vn8Kd8sDD+ZskmsKJNZNgDWT6AS4Qa5o4M7fptjIc/7B75WLHOCamo
BUyc8UcZbwv/+J/ZLeII2couh0umXelG+RLpwF4+ccYO7RgltAqP9JnqXGn6G1ZO
FQaQ9KhumsPnlfLdpU+M9BBI8T8eZZO0us0+yJQDOV2rtT7x1enqUUXIEAIHB1Qo
jZ6SeZiNBYdwCNIVdWv+46MrBvRXXtLFhZUhjSSHOzCuCaC8aJWGezrWKiSms8xw
KEsf7bS7m3XuryDVneGVPBaSJfdZeV82nHpbOlBGlu2rq6eogjac2MzMRHQ2TC6e
LFXyId1p0S3kPltob9d10ik5UAEblG0uCT4kbGDY7vvT0e/1cNMA1p+mNodrKUQj
KinfpkvuJM1aApOhH1t4RzGvjy/iilRm4D8LP57ucEMWh690AGAI9GB9MQhvPJxe
/yz/VUneNCtm+xIHi9LQNK5jJ7KRj5gjOx9/w9KxhKIKPzqMyFTBXQjlOx8BcTY6
3NHTk6GWWAv4sptGPUuhkfRabUWbIG+0eTynye+go8mIJpAGW59eYRkMcW2qA8Xh
ti3k6V1PWDwxVaheUFv/sBVKlIHoKJGBgScmziz0mR7N4chePfV8rTXRoOF2XcI+
lA//BQUy3WSTZcMDixeUr7fnV52QlfOyu6YXeREwKY1j1k77c8n7KezChi1CSXkX
IDoL1t8orfc65G6Ei6Gp0ZGaBFnOXPugOal+OMVsIImDXvlWQglK2Tpy5+JI5NT1
xTrMujqWzzd9HUyKIyqxk4Qf4RSnOdXEAiLRNnthO3ow2rnXuSpVzNFSgngmJuwk
e7IlfjPMXctHb0WY7adcznS90EeaOFdSQTpHMpYc7dDehHstRAUcSxxp7Yc1me/o
Cg6msyHtWaUu8XR/PwQP6a4Lsj1oVLXrLEKyiJOzC8PtoDLdaqG+5r6fxbU3Qwyt
2chq+8v6GWI7XG2NiY8UkuZ0Kuf7iHbDUJXXk6zpde8QQG7Se/5TtvY0hwwuuGwY
VCjVYbGHJSYA7IujYZN5EiKPzVWD//I537eZ6wIyGoczlk7eFu5MVlT2DeZp++U1
8FjMU2voe6rJjmRvAc6U9+45LTot9raROO16L3xAlO6R7iVvqDQRRIr7wtfOl3Te
IAAaKYUejgC+UgRJjw601Oo0k8rpokSZnJucOFQYmKMZmf19d6PbYDFiV8jr4fDf
L93HMNKDc3S8iCr/GQBWpQSclgnoIWDpXqjEPRBeTfEH0JmY5YQS7w9Jybz0n4TH
4o+IfMjU7E+lzXUvtP/kD8KfbIUSavwVzUfcp7DbdVQsfqOfXGeF/49JM9MIXKHq
aPXl7Sq4lsJ7Y+cYRidNRpbWDWZku8CYYq4zRSOW+x/wrPJmCaXG659yd6TW0Plg
b/zG9VXNwYd0eVuaRaRTdi5uXjFScszWoIYQgjmFxppZJ2NyKYJkMn6l7RpvzZSI
oXEnFsXICASETcVdfXNzrxsOZHt8tiw6OygB33E5EGab/0faEzon2DykQ8P7UdTt
uLQp+o/BfkKQnNpswNu9m9KpBqoTYhZ2ePZV304XfkHpLQhgnFflj5kEWq5TUtam
JuJstCFRND4qQqtvtX71Il8N6QzFcTM+gdKK7Aba0/cMlQvtMMROxa12kS2EBKtr
N6/KeuvLLGjs3zZWkRj1O49eALta3ZPX1owonmUjtsNARI+wl+21qDYVoo2knTJI
1KLs+pqhXHt6bHEl+gl7E8Acc26C5wMPVEHHWcfHbXBbPkeo8HP4iWntFvTFskB5
koY6R/elXjiOgfqeAK5b+mAVd1IaWqx/Gk74ZpU5eaqaiNDso48S7d2pvPBDCUik
XgL8qxw2bdGYnArlodPiZOYUNksqV+vShFZz2pwRyr2z0D5yColH1GPCy5xDOtuM
g12KpcLDRKk0uPOPAD0Q2eoIWjxKay9QoSPn1I3cVtq9eqlIp4dGrXUpXKZ8Z03H
kma1Wstavl342w8glFf+vhAIdHOQaT2tyWMqZuZvpPGrS3V7NeDMj/9QTw6ytyPv
SVEMVbZybT26+SZVIxpyX5VSTvSd5WN1CsyJUp4ojVEAqJXncNAgSimakAiWsJbo
E4z34tczloXNuPEp0z1f9zbGCaCyneAONwv+Kt+8Cpf3EsZKR3CwAABpGj/cVaSO
2SFMeK+yFt1KeU3JfdT3r7FJHqahlG5l2LCVH78RhrseUR4E/KiR65HTvDf7HLub
rE9XAsk2gPVca12Msr2gLS+8gF2qYIHXYicr7N/CDuS3gv7Q2fxuDVr5+FHd9B+2
i7Kyc45+oHsFH0gLJ7ZCnWqKjb8sRJBsPv3tcTNpA4Loj0sw91njv2/D9v7KJB4q
kT4xz1OeFXqjwCJxejkzz7HOaV4CgecZxcsetR5hYuOsNx+xcTNSMIsLQmF7Oa/b
vV/rnvzmsRrDKlL+8IheJV4x8BZLOOiSSgKmegcUlmR3a+wQzw9+K4lXOGgeaaxh
L5RDllPkPH5iI0+MFUhSFN7m/bkzd6mRbOswY3UpUn32xO4irwU8NOCDw3+7wrOl
wlFa26V6q8UKtkTL+bbnUpBsqxAYoThMgspMBq2P9oyTxS+wirR7Hgocd98XTYJj
p//OhmNpFMuegfSoMP4M2/gstUddlmGamBHfN5+tGGK0S0ID/GLuzOi+KFCtLIE7
MgbeukLqoPUMOZirlSxYUrsvSYOUmd6rJ4aFluCJP3iwmJkWoDYEy3rqWwWsL2ny
oxW0iBJB0u+m9jeIn/wC7NG9GLjiusB1SZBHDBi8v0A2Qr99PLzjDktiWnXVXFBq
eMCdIoGtnDKacXcU1kHCxQQrSeOV5wmQ9FbHTktXxSvqJ+EOR3zcVZ3TiemnXySu
n1UhCPdScAsYlde1JT9o4GNt3qfPtlVxS/AOGNPpPOQnOK53uZbTrHJIXUlWDNPX
dUwqTYvIPygCz1ZkiD2oO20Vn1iZ3l2VHRyYo8ruwasVr7Y0IU3zxeHZWd9RIRmC
gYGabmQg/RAtURNBU2xURNaIJl/SJUA98qmh+6ihCkcVQCmjpSM3BJgBWQNLYHZz
FuB9oQvsZskubXfez1Qntrg6HpVSEdjOKEQpmBmBuKRHG+PfcPEPnZJDLgC/wMxB
ytAXQfnpq79lhhGS9ZVvpB7ETNtEHXpqgfgt81805OOE9XYyXio6CPFPqiROjr2M
9OkHjLUwASYowFZci49C3LOjFoK5dyqneZ04fTITpKocp33K59skN/alhONI59Vx
XnM3xCd3wPXMpeuxZ6t4AEHrscYGC/hAyzW0UB10j21F3yTyjaaQocwaMyCslGoh
x46ni1NZScLDogm+AN+KVRL+VU7AIMR5dSsfqIorCq+KuCWemQaA0vVyCBDF3ThS
aIx+/7LfW6AyqsB7CdSupFkYLiaSs1AzxOpgvuAp9Kz01MYeYF5MHa96a//hTTjE
/MK1h4j4KxPyICAq0rAuI2W6w1C6UhtZqKm9MFs/Mec0nBMr0/Re98LmKv+XNsJs
duiQAU8DKNhpbV+GWygVaCeCBl4zX9Hamcba4H3RNtI4+bFtVU5mYjSiD4uiMRG9
w8rQNtQZdKHU7jngzw4lUgwSj7SJQYEYzE8hCekPP0aeBSN3SShW4nM7ZI65/zGc
oyzGgupVHhxS2j/2zjdF33cfcwPDpe9uM9XYqxt3PYgsPhWEEC5kC5+ns2krWxYL
izxLw5hcyKd+lwGP5mI66D8Dsp3BIFhTHMI85Hh53U9iFDJEKN75Dg+mYSriV9Mc
n0khvghrXai7Ln2o0pURY1VrktyUGpn91VrdvLWmaU1ajo0hUl2bH3beWdBkOmvP
fR9LWE9rzW0btSVQuWbBrXfLD315wAS5o4SZ8f2Q648xSnR9N1Nt31ZDl3OH9/pR
T28faCR1RQEU+fqVDLLZzAmTMhXPl57ydiaA8VwE2scQIV/B5RrwUSLGAxp+9G7+
n/S9Nd9WmnNkyI7xprOR/9NoHrhSCkfK171frkf9Z2E8o6LBFw8xL7Y0Qi4wSj+5
BGSfaQ0t9nJl9VCZdYr5okmucCS/149AVWVagvWi4pHVKLtH4wy2RJo4xOlxuAGD
ONt3ZPeh1a0c1X8+AXmh5HFn4Ibkeap3qkCfxmiKzTn60nWGT/BazYvcdkzs6IWQ
NiV1duVLcuyfAezlFv+SBxeSyV3w82Ecnyxhf1kP+NL1A9xkn1TWHS5R1kCFABSB
4DowUaSklKMfLXxvXTKsYdUpJuQjWgeLaFbXyAhSvmji3XRqRhY66Bq8CrtRw3AU
qTok6i6kBAyKRuouCMYTX4Q8MxnpJzAgdPdHNfyMy1BlipZDqWNuxa4Mn4zVb+Lc
H0Oxbp/uX7q38cMl0aQqT5ZTmZr7Owd+2Viuh6XIOAoOqTeL1I1dngI+/Kp5489D
PT/aYbqJJJ00KXhRXrWua95VbNUp7/PUYIENHlKCcHDW7DpTE5faHzSAGV2VssQC
ywmz+yMIlPKVJ77aepDkRJzec9qbQz3dlgiOkckBSnHhop3lyiONw3nQXtV7Wm9H
uzYvku/q7CbXZtJdkNSPHr5jv5vPMBhemOjQNmoD7XfPnWzmkEoUHx0g1YSassOI
uOM7hy5IZfboq4dnplH/SW1UrzxTkV3G9+iZr9AQHoIQHhPbfGPw8ezC9qrJjJj4
SnxTYEX5+dsHZEnjrwdn0D3ZaPjFyQn+ExMIOgO8KDOAeKVTbdS19majmrl8rlI/
w8FXAUQxv2vf9us0b0sSJsguVtbFGdVxXYjV7WpBhajzH3RmWlYnsQwpfUOI63o7
VhIdi4UYxQ+dYROho94EsNBW2lMqlI6XrD03Ysv1NRL4iEwJtZ8dL/GMbusqMKje
KlTwND5bEoj6twnq3tnTzUX/ATIHT2lHuUSYNFXbtm3WvbDnr21srxOTBCCyIw+P
US7kkiY2x8J8BiixEdxNvtmytj57JEhv/9X69y8H7KHe1KYXuw+oKXriItCcAxtM
ScQ20RGE8mjCIYseV5hi/ASTsdDO5BGUXonB9Ts5y9qib8U3+DOK2+2agiJzRgIg
/o0C+YOrCrAfGz8fzFgSTEfxAHTQcyFgvh6Knb7/DqqQIWzZ782g9kN3DVy6B7K9
oMbjglEGRylHMa+xWJ01+dc+F10vi+ZW6h40qo9NEqkVfPACTWjicxkQMneeOO81
etUs0k1NqA7iL1zI59QYqQksq2o4Q3fZLI2wxgHrgZ4aYZxfSzzsTg5LwCaWvqI8
/xQymIL1O7ZcI/MTttU5X3q6RM8oZjcrf9Nd5lD39f0250aJhG3HfTkvXWpYKO5M
6zG57LX7Zuw5vZBPYLM4rmYHgLdKQHAt7zyGQ8vg4n8qEyjejnlr3IesfAhiRyBl
6ucQXc2IF80OknvqvPVlhreT3k36M2Ub/tiMXjdroklCgYCz6YPGu9FL1DjlrKkk
duvBhrTFgp7V+DJ+mCObwjMW5hJTB51K+StYoalS0KHZqgEqect+GfvaChaGseAt
8SFyMSy1YzHAWetd7i+evFGt6vzJHQoHcfOpGqlcaakxc9hyae2KFQYbTLfj5FYz
vThBObRU5t69Lhtis+yRQannS+vV8ApkXMtieXbKJJ8d2Ryl7J0BijqypKt0wXhF
2FvGHdfeEe3bWgYuEAy98+bvkBlvPLDTRpET+TF2/LN13JFZVb4wI+xsd/S0PNlc
6woQHkIZ/LgxJ2fEi+ID6NJzidP7Y+LXZ5423hY1HBJdsCu3cY1E2mbbNrkHIrSn
PYMJB3ovNua2Ds8Gfj1hKWRYyOqPT5A+ViNlCpDVODTzjgGfagY9ohqZ+cHiHIxm
eLICl8io/9gh4FkK/Fk6TceRJoR+gjYi84j+ACHaf3ZQi5Z3qhtjlo3KQTqvr+/C
eW/qq/Q7XwJVHXgda9huiVhJcBGiDqO4/EaQnuLsXL9qXK/X43TE5+kFUrsutWfZ
Jxxi51kC6wmX7JGMsavdPU7mDPS+B4mDOcblQGxWHcgjpFydjrxe85yxPDmrsDQB
JHWDjf1R/P2YYuAMLWYBWGj/jvW3pZhVX3lWeHQw3mHqK3tP1U68Dy+xhgxLWb7S
G8OchNhJzz4DgMRd+UuS7MlJMDDNB5glBBqvAlyv/rN338TdCAJ+5xjf8K4xdvsC
PshU0OMpwlZ58bGEPFLjTXexK3lgjBPhQ7gaUTpJQeV2a+0m1u1RubmKYDhEOMro
h4DmyZz9THxEKw6n/u2Q34XItFo9Giix65XlTFbx8L/NjQk5RR5DHEGkHKLitA1C
homEBdk6vxDLH0rUqUnXHniNttOccS5sdowgVq2h88S/k5UFhhd3n08qBoRmMcsK
r1tW+qctWc5v+cHZE9mG1J1Fa941VP55bIcONuJKi0AV0tWM7FxOiu/jNaRKVkQa
pzMdj0nsGwcERkRfOlhdiGPC471SAn0FydyFsExyAcwik+hJFpNYwT3BYUEIe1E6
49FRQfUkPFlz1AKhias+wspUaZgOG16Q4lphrbAr7DcyHJ4mNDT9CbFluZ7fGJMk
VffQLnTNOvo9S24Kcr3Eex2CcXx8p03pSGFmAyuuXNjRlic0pRl0VIFU3kPdvPQG
IRY3/ozJpOupCS7gnz+XsPCEK09uWyL36FLz6mlFKbm5sVIWCdtlTiV7MheKX/HL
ncgmuA11gR3TQZUxGAu63c0zwrPHQlIjqQVF3eVTjmRgTOC1dJoE3xYUmpXZdkGz
jYoyBUmz5UAeK+1xPzHJnRc216W+QA8/gXNMwgaMIAP/WQYzh9pUbouXlybBaMFh
uTyoEsMznEmX8XCuEOU+v9IN8+uDmv/A4Mm1zh0wn4YkeFuhUbNDHiX8eM9Xoub6
GlsaIku8QYWgaxLZjrnPDOh0SyJLWbs5OWatbHo7nwigwM0la3K1jHX3+9VcbDIX
Mtqa/hCSPLH1Wxxs5xM7VXbXvnNufjlUu125sQFJ4ue5xIVJ1x+elQzVC8L5FZNB
cJaYlH5VaObXX8Ejpj/h0Xuwbo9K3Ldc1wx29FQjroddPOt74HLo6XfvFmKizOBG
OF2V+qe1vLFgcvO/d83ZTdjFiLD3RE8JU9qcJFLDF+Jm7mbVLT7r+UdApHxUs8T7
sWDzLLeiceH1XD8yCuUb2Qev2coXBxc27TTA73JoRufnpnNBngArfO32+Znhbmz4
zeMIhW93j0Cbp5bECG/9eiA6kN4FnQlprzQtokgsbLuzAOnD5tS5OzpvIeLUAT96
VIZXrwXbErGsZ6AUd0DBBkmr9lUMncmkNkd7PNZuP5jMo6VBcYCbbxEvMo5DtBUE
W0WUzAhKTmA9tQMWf3QSUyqbmmBazoJzCX3vZVSrP1rvPG02TCQZRDWU1/RPynlU
xlFh5BZgrvjFt2j41jzXekdpjMLbIFoIH/13H+/xDGmBU1krXeDAagJ5T7M22/IL
gGWmg/IaTjb30rvadXOnlfXACosDl4GnyRTmDDX2Oa+HVNqx6OslvZ2HJ839IizS
YdJFgCF97szAgC7kU8V13C4FV6N768igiQR5V/h+QepUzdD4zFHnJMzUWQ0m9HCt
0k7oSKM1kyPUCGI6Io69c8fZOylNPeOSLO5eX6Q2YbHwJDOC5E7PP7M9X8e6F1+Z
tgCYwMLMbGOTBvyafuZ7gSt0feBrFj5RGS+KLc5QAW06t9nIlbG5aZ3xRv7c9+Fy
CHUCD6+eBkW7mZUnxUEVQnIJyVmLR68uchFgwbjvAdSrK87OUazXGDJBs9L9HC6C
cnFhG8Y8YSEjJJvT2FXiUOHFfE3bvGdLxWqsaQaPX6IUkRWIwxs7/gh0l4CE8L9Q
9zZTeq5VE+LazdNzYmHrxqq9cwihYELOS9CdJ4uy9h/o0VTYrBmnzjfepX8DfQPX
WbZ6kgqAN5hI2BWYiporSStyRxSydt+Wx2A+Dv0J3VnmmtopcmfMZpL3N1jws+ha
WWNq6kTvQm7Ya/l1YftDm0BbUBzZdu/kVIsxdtFmGXTtYHEuvymxmwcyx8dUdjIj
8Q3/4eucF1n7isgG9+5aTAW2H9BTYOsGW7Rl8Audz/+c2FfL5Z9Cn91H8irTPmD/
IgSWcDPqvx2j5u+icJv9CRRHpkrlTv4dgOY7GT4WLsAAzV+VaGNMsKpkW4RQEjG2
dal3G5c+OgIWB7U9up7SRHPSVPMrqB3CYyJ5rA4NFq2f2sNpwLmoiJvjg16rNluh
lXi3tbY87am1gCAZaTZK3hz/dmv+WyTNzgBzFKq8Q4MDh3kPK0f0Vx72Ro6TRJPA
HirRGv660ltN+Rwq4KUTnPyGLDrvJLDYO2/JyEUHL+tYV9JHL+iP/wKF3M/g8V57
8Vmhel6nLGZ9V366G9OMIkMe0zvAfXLQiP23DLwUcjJwvHJmWbXyqueqjWal5JE6
I2xCHRM1ySzZD7Yj9g8F9pR4OgFec5jQRXghArq2hD1NA8W8f4OjWVQnZh5Iy/mb
zwkEpY6KgUshstYKCq998WmX7g8Id7j6/rjN2euBs+/pyvzHrF1/O56lUAfrAhHM
igiefHy0zeUyXUR6fGnLu7RscDZJF/6F8nvtm6qJFlqQg9Zqsc/IMojshfFkMxC6
9c0Wo+0iCJ1ziUhpjt27KhPT3o8PCrAFLKi6Z+qz5GkpNpCQxhZc34rEYTzcR73r
WSVSfeWSKa3I9hPg6ctM3vJkiMNZlBcvp7fYwmVXDVjL+QqgOi3O4bA9gtxvtJai
TEL9Om4PtpY9dHrpK16IUEkLjTjq/vtV0188jsI8yll82WRd+HP7/YYEIT6INn0B
HNN/tkzLt5L/B6uNnVccFQQd3JzzEb9dfwrVDS9ZxzQjj9EJ1XGWMOZET+CFL20V
QpoQnAUM5kJnC2vRNarp4ohXMBKQJb23KIE/Bbg/rmYlK9H4oksbpmFG6+qwzzct
tOqh0j3vZYB7ry58bIXvZ99NQ+ZWG2FO7bU7Si0VCJQ2kDtuyh4WmbUxq9rW+P76
AREuh+Pil04EKTHoFf9Tfur1xvTNBXmwGjOD6YlJ1T3NIn6pBvsVpzF8nHbumWS1
8NfvrAkFdVnngfzXm6xy0gAuiCyYmn69QS7XWHFrnLt4sqC1aM4z72f8HB7DPpKy
/uGf8fLO5O/F051pcn72mZSbR099/R4H9m0+FNzGOra+TgQyl+QMLgQwMhSAiJP8
8KzONBoN1znuL1+IuTSmlY8YSrTkoHExD4Ugt1HqBjGRl/QxywCUqRg21WMlMDM0
V8GJCjLwnzgPKN+3/QQJGWexXNW0fen+fA75oBDUNR7YnR3l16bdrrQdmQtwM7Ho
FFU9DUFPiYNhxu8h3t1WIwV7+tTRE2l8rvalFBgraDcsGjqauF7SG12+1yUwX2ON
IGZS82fcGL7cKGw37TZbr+190sjY+ROiEUBrzLHEyG8MZxfT8IfvXn/VvDCgi1jp
uoSXD35/IbhrsKsxwtskjwS9g1ZyUfXXNVdrTt5N7hOIDTKsv6a43niRU7IdmMvC
tZsY702cr2I1NnauUtARQ656t1WGk5YMj1TwX+Y35csxg+ak3h5p4t+t9akWwmiS
3xHSFDm0UxrbWk0LcGXI2N71YVLhTuSSzuVfAYuBY7k68KSN/IYYZIDd9B9QZQuL
bd3EIq4xIprj7Y3WGnfxeX3E9fEPA5C7gR1k16j189zK7g8nY6B3ArtZsqJgmc4g
ZPV9YsFkkZ7DbDGvp7j+oR2PoFfHVYZ2YQ4Zv4KUx3ZYEDSY09mITcvpD/t7GEUG
pyFUrKjYoxsjwrHxMpEaj8o0gS9QXtr9gRjrB/CUcPJbg9QtiGXuf8XSPf/rhzZi
+bmvg/8EOjV3esYsSHkMpSr6FxyppbcElkXepI9pgmkBNDKJiVeT/iKW9Ov0C5cF
16H9YA2zbU8Xf0PHdyJjtO277JK9qTeMbX5XnGYEqLs0gDOa4nrwb3ipEKWDrm0t
/L9E32pBq8DMld9Mqv7w3oZlKAKWtmz0D+u9bJQJW0ZpzwF2Qfvd6N5NAc+MNk4M
Y9pI0Tdd/0tNuZy4IYhutRObop1yxnC0KXX59W1B2dgRi1gtI2hSiSufpFeganen
1eh6wC+poW3srWZKsahW8mPM7RxU3+ytFvy9U5nrvG2mmdYD+anuiEMToevPPL52
CatUBhYkjbeghHqySjQICKFizZaJZeujbodnl6N7UbTXFXiPB2iryUoy95hX3vzn
ISO0v9txOIB05WansumWPHwYcgVJISOhn+NsB8UOFPv5htLTzw7crPN/sOMPdy4V
XJfnisRpULqmwacKaQY+gzrxeUAUw/89t0zEkDbTSuTU7S7Og94w+Jk7KO0hcNXB
sGUy+736636AeVfWDHngzrqXZTd3pGIAcgtJY1UwN8rzhBgVXNKFE2954xSEFveL
fB/gVa6stBWTPPbuEfi7P16wNRVP2iGf52hxL+k5AcfORa8Rox9ICUK4AkS8rN5B
LsPNmUfJn1+lI0JUMiETc1oeGyHe/6W86Tn7r2OBDOPEH0gxkbhItPWVhTEkXDue
W/os3MKgPanHWO2SC6zwJ5AvEPwFuBjnJLfZzUSBK/7K4H/Wq8Abe9FM8zjIRcBd
W/oPDg73xyqG/HewD7A5TI7kzhpRJmL6w5ELYbaFLi9DIymar3fNjqMwZopLgn4k
g8sLdZp2aWIV0RhBoLZTMgcim0rhKf4fBRc3d4lqLj4=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
c4vqA6zK4P6FyBGZ0ye6IB/rKwL6vT9dCGYXz+lNu2opJpb/OFEMmf9TiynOxc2N
5PvXjpbVckCEj6nRKfZF2+7H6rO+h/huAfypv1oBgYdAI3XKfe/hyn4EpwEA42nQ
XMLUaK03+nDc7RIYriTwNyewTenrS5AHoOmwItzrwAxJ0pRSrqhRp1SK88qX1oZ8
8zslAFOigV+4DqmG++FBMFzaNv/R9PWBJ5EdpmYX5Br0VMLDJ3tZo08+F8u3O+WZ
VYveVy+qO3G01DYzktnVvGtQYfX4F3MXAsLmrJvTnpp9K5Uwrm4unQ22C1CzW5/7
x9FAO+zYZufOHy0jL+v7LQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8672 )
`pragma protect data_block
En7662FODKwpUg//1PL0du03ARXRDOc6dvOrn9/0WxPA/adAZKz2iIorzBtN62zC
r56HkyNDVPN/CvfIi8GD1rSWDBQtQlC8L0MQPoughYegrZpZ/W6FcXeYv2sxtAg9
hwovDx1GIzHqDO+fBjEJnCuOOEbME0NMD9JgUPhegbrSupX7wpn1mc5rPhEHeOVB
GB5zNlKEsjBz5PKhQCn0Nfy3bdG7Xy+bPoIZ9IJFyPWSHlH8eQxjhU1EFbaB8RxJ
LB4/5u+oXBbBPRLgOpHdGNm4pJHxqh+ooVT20r1XpjXgy/rA4E3BwY1R7Kguik6B
LfRRcMlhz/2Ok6lmGnqtMiIsFJMrle5nCUbhFLWVP6kYbcX6yIfb7VN2vORYdL6p
2rh+uGdd9Jiq1zg/EtXMHyphE7wtxNM/jqQ2YqGf4DqT3nw4/SFPBtznaKL7Y+04
nTeYM7g4KqxkR4kv9XXeXYenmzH4p079wIOTR2QvWHkAQ4f0q6MyCo1Sa+BZPvbF
Oxt/0fR1u9+0r8CwEe5wzj0XwybA29ZVEheLQu6TjPg9gJWBhGE6+tRmoq4K3CuQ
Qb77OPxheTHIY4sFTu+LWwuG1dyWU5VYOohFVVYARiBhqnJ009KWcmTBKq52oV0j
ZteA7WsFXZKDpT3gvxW+2UR1P+nrSNw2m/idmELmsvKAtbCc1jdX5buGz5OQQ6vF
3cQ5qRgqylCxI2OUYUpYP3K20QBL2tZ4dr9HhilZau8f8D9aAr59zKQ9kIlHPaK0
0BqhBVEsMWBVFoo9FHxCka+lngcTWqjlxy178oX+BUXtS+rWyjuMBhqbQDIw0MsA
+aGkP0kgBvYf2I7UaY5PS1gL9MDOGZOiSSqHDgErFC/FCDyC7PeknCspobX/jPZ0
SyMWl7e6LC/pX9Y62cTnvlLBsIdOMBscSBUAXIBzsHS1a41gzLHfVhqOCoBCqYSZ
3A0muai763CxeZL8GgIYxCYORvpl8j4w0rztB2hXVAMtavTeAtU5ne0/+huiR8AR
aP133tz1n0AP4sVOTMyOjJvINGxTUDf1RbysENRkG11zO0eljt11Hfhl4HUyxEn6
bGacjBc+pMzrYpCbs+LIWLewmGc0NJOfJnt3grRthZ3OPkxnt3RLZ60jzI+3u7U6
BBNIoTRL06DQUjyW0OOpsgjCqOYhStKLHsE/aq1yZG1ZqFR3SP5IXjvuChJJjpAF
aH2JUzPh4d2t+h3jMuwq8tHKy6veZzBeGKogIPbMkxL3JiRSRWF+zXjHarrSOU5d
6jirLYXVmXRtvzVsR8dHhK7YtbR9bRg1aMA1iax9l45xkklNgDh+3P7UlBCCm5kC
favclLl+IpBHyFPob9AgnbqSHEqz8Ve+awuk/72nTJLrkg38sHXl7u5Cu/CQh3I/
HO9lPsDKzPW5va/Uklj6I69zjzhEZ8iXuAeULcNWxcOChsHLMwtH8bxoysG/5xjI
arXSWi4Fb7FgnaMQhYTyXpN5KQQi8V1EFQVkQt7UANSb5Qj31U4lvEfFA3lPWGcW
7kuJegJL8ryXS0KVICc2CFMwlvMy+v6U32FSVv49lodzSMbaiOKaR77Xw8gK0+8c
ZHEFrvT92zpHOtwcZUZv33dlcSlYs/thnHIlU6zmNLiJEDKAiMS93T+qbni1DXny
KaDqy5BSd18rnERow7/PsBSZfjalf58neDNSdOCXzYz80trmm5hpsPPemvTCqpUN
0lZGdKPoCcIFHHbwnheZ9VYZvNlnT8H4+9W2bDSmIpKfGTDJn31WhTTv3ke06XaD
LyoVDZaPFlbNxjETqU3poBMIBbmHGl+b73faf+JTG+BieqhRqBQ4SMMA2qIjmmc3
3z7xUstZPp2oDORu0nS6eS3SXzU9srzOEAey2bgZdcZlkQt1Dxorr4DAT0MvV+2h
V9orDI8W8iln0WA+NvcPmzZ1T750ZzWhVhsDzTk7iCw+uePT+pKllC3d8xqigZqC
Tq4CtPY6bh7THyc/cSAAvSebx+YQkxrmvgUYTlqPtAq9eDRypm35QUxSXPrAH4O2
xVVwOsiPLNjn9oJacgzLt+9s1RQDEMBxPJtuC7l6718Sw4VeQ0OOyIsXxmMJXxk8
eHdi7nrP6h6hrHFxOiDU1tz4c0CTcqeloOxc/C7Nd0wFg39ZzgiuaPCCMUx4ORMj
ATm7jic44c87Cv+qP2OEr1nQzA31smIjXsbu9nwqTc7mdjqzrc4qBfiolwgVSzqK
cz4eKomyp8VOlLmmbBdTcHcl5hJh9+KtqSo6xX9F99YfDk4DJsKdfAhXpUWmkR94
DrEAXy6wOMKFLvsQfz48yHsU/IhKCfIWLWEG5nE9mIYMw6912IkUvUy0xH0SPXlw
bV3VUusGq0lvoB9odN1wJrcHq0R3B2Q1mUyZfkLBLUzd/S+moSvbqT6kAlazmQKQ
GcURQPCb1BvYipj92dU/vk1/3tz+BsTSr1yWeUg2G1CfRNX2fd6q4w4tpc6go7wD
0vmhvmcjGbOe7C22VbO2DXUQvB8FyGMYljCibUIEJYpZIfa2plfmLAwPcmKpgyAS
EcdazfcNrO6tkl92hFfjye0iUk11/udZp5aqDcres6Ty9wvl6oo4cqXmt1N/Tvjv
ogblsMO4UqPCRw75M6DbHU8yVC0arp7wWARmIhtsdnoNFcM4gaVWkHwSGJEKiQqx
JbUMo13ThxvytgvUeIhLGkZj1txTMSvFE+FPcMlpGF+tMQHIGHkAxfV9QB2t957C
JXdcN61X90fSmfif3cfQXrRUsRQjoBKsUgMTptRIbCPeqKdvDpNkwbICV7qCdyT5
o/xviW6iReInCfC+gmYZK70fUH794iziNmSe0LdY75B8+B7b9xXsaLShTiIcFA6g
L65TCIprweUAW/GJuVBTU3Vg/JH/Cj1CoLHUfd5IRf6G5AzTMgNEPDNt4Vziwxrl
CoCka2C6YutrLCOlJirNDfF5bDFuw/t9DcwDHLBZp2/Sbw6WbFr/USU+jZRwT5a3
oDIpxb6UqESE+0h0HlFKSszOcBqLgmSvcGRlkK+aXFlGC02jEo3kmSV6Z3hhpHyH
7nzsm+TQnxyODOehCpM0Ge7GDbq+VjU6gdhh71+rx/wRsBfjJ4siNxKwSXtXUT0i
9AnUFf1qs80fq5UU+N2FCTaEojJUvd0Z5JNhiPsGAWDweqItHhK4qYW/ry94K685
ECZYJp+uqzczHgY1hAlh9vBcwQE7f9rJ/80JwHw7qtt5B00Twhnz8yUeqmisuoRG
0kQanduCyHSJpjSn2/+eDUib9oLyfJRD/AZXR7LI8Doh+N0cq+6zKOCsDldzEdDn
zB5cI1ctKhv/YSCcw3ZZ5/v+jvSXt3BY5WCVQK0GzqfsIK1yvi5PuuywaSH/gg8+
tqimUVR73hgc3n2qIeFIGCZAbueDGOFfCe+uakAqBIQnIo+2uKpPfIk43E/SSr11
qZ5R4yXpWbge9j1SooognZ3uS+SBijUWiyX8dTZzUCNw0RlUvXrszDTMGoAIEoEa
lf0aws5EoJs/SbaPpcXSDZqAgpAxB4ujdzTBQWwks1n+Bev00mIqReYchiP8SBcx
GS6KBzXPhILErDa6CSZUcBZQTBFdpAOwUy25vPkvFIlG+oC9DrJBczcAF6WDukyI
1foHI7pmkqAqceXM9m0yKQsGlDW9DIBBkDyMMR5VB2q0zN9g3jnQmq4zPdkGGjbK
PoFMRcygCl3TFDQpSAdiOzyA4IzeOdxbL3pMEbyLVlH/ZkL6BBvpLWuJy7Q3B4UK
L5v64piDJ8OKeWrg0e59O5FIRBEYm/Rkn8RSlhu1vHXd3a7YwV30+iX9Mf/if3Eg
VF2DO46ieP7HK3TEI5wj1EcATTvCB5QoyhtF0tmnB0VyDJctkrF18SqSQ6qf0Pdc
vQm9yuD2fLl7gDMxu6cUa3oG7s4EPYbQlXaOSsMeTlZxFrI5OlMS4akJanL1ejZB
0HaQS8D3Xsx/Elolx6d9VQa7NONtSTTcqx5/wZATsgLT2TjR1FfT3WQFuui1NP/D
gZJXpaDm3BwoN5N3mYx0v5kRqxeTe691Oogj+8s3rx4smtpVHFQwG7fuG54b8xj3
qhKP6GKhgWdQy14VOOQeCcBIFAUaKxvzoX2354f2c0hobdv/sOnJvHNkjt0fJ5hl
Gmi0woQYp1cq2QQFZbaJIlL4uDcA46VDttQuElFWwNoaEetKxSZZ/kWwnK9BPFBM
ZQUuUI2ZBDAfNvhG/FlQZ3W/gv2MMQIOywfNwcyEDKd8Sl9gfBn3aLw4iWLDx3R7
9KD3/qia67p8kBVXb+fSVoH1lzZzrOtXjUthB5eGfs3JoMw2ezJkZUjY77C5P25B
Wc5MIUU3NmkYMHUXEXTNG7IVYfUFpDPweVn1/QwrDOn9fQr/kRgltUSwbNkHJVoD
5NQ/JY4CqLbAbAqaNyLD9JfH22Evur/fxJ5qgUPA2UBS6LxnwH6MOg61ZlpVj911
+GWM2mKT0Pvq9BfcC5IQdQljR/YYZzayRK1CUUEG/5PsGcRsovP18+xi5iWkuN7G
occS1Jiy9NzCoux1JhIMBcBZ7nl1Jw42hnyFS8YAXaY1ceyrixAGShAnSj+h2USW
89RfUrfh+f9TSATxuI5jCREgZaovUmW7j9YtDwO8MEs6K42q049aE6pLV1v1p3G2
Vqn5iAHx2e6rLYTshpB+VdDHMSISkFUkTduhQ13w9p3yxYHcDFwOWmtFtgA0nbwc
mR6QwAwOj2adKjuzCVvDEtiehEiEAnJU7EvUcguB5ASHuiB3QsnEONPAxqiNguJI
pD4/fdw4Cn4FnBaRzbVUf8UYPlxMAj6BzSTMQ2NAEtUfMs2nokgUHcHBX0Eq97tz
lvPdBBdmp8CFGNAG+uDNBpku4Lmrj2q4e2TAB7MIM+Tnw1tJLDbwX2o8iRp/DO0h
nOSQVb64JHYgN3z0TbD7SBPLoXrSgCMUMB4eSbLqIzCyyBWhQ1p6I4aApbZoYEjT
8kOVE3dXSaPXfSmbR3wgyxeVqtyQNbezZVqcalxyOyLrV7h2lPWqfSFRpzAazuiN
/SPcYFAaSiYNxqCjqBzox3yzkzBbvyuVEV9lzXhtXGmciD1On6XgGm6PG5yX1oBU
M8ZA+u3UOcYJVFE6jT8xWIAjz9tVPQnN+8TPqf9TXBPsruoYRwmfI2nN90VqyIIM
XUtGDC+MBPHFwhb0QAiYx+m7nECoRyX80GYeXnIKgHIazK2LCCVlPLsvGBoYsE11
26th9JCKJVaU5/zPekDFNP2V8KBR/XEngzaj5Fx7o5LxCFKaAMdRzguRLitcRhe2
8Jf/ZfnnUiL8kPMdeSlFXbXiyZtUT2vwusvim5VJpZSc+iYICIzRK9wh2Ximz1NS
9llQpuHe1bFI1p3/KfHJtUNIzRJbXzZHrNgZk7h6/W906ClAtG2lh/ouEjbKg87Y
9ZG2s6VR3KtGwzAelkK4lckUVojsvDE9njZOhCxHqoNb+ZmeVhQrTSGx3WLWW771
VMeLi0Ke1hSYqzO0qV8nL+ahnjSqcEDBRhybvEng2O9I70fC4KK5LS3fG46nj5Ck
LavHFunLA7IZBzlwv/S3a1DXq/MCOvYgB+oOUdkCJgL8IcSL65539GEHy8LK3efp
AIrx72sO0Xxcj/CuqB1oA/R+B/jXrUO9S7dRZ1oSRJdbCpJINnqsvNjf6v799Aao
+bgknyudg3IOMKo2BVDxc0eFYc5FNioBvDDpILIX+9fPXG2oLn1b9zQpXVDvWiFd
5KPq0s5BBX4Rv/nrAB38XF38pZjgO7/c59kwoqYT7fjteQVuqjSJ0QWMlVNJ7qeh
QALnzSa0Zi8TpCFGOa0jiufOTsRcyaiAGpZ+MFPTIc0vIqubXR9DmpMRa0vDLQ6P
mR7XOyHSsRRqK5LTC2vB1duYFWmpW6jkl4RIo44nAx/w9QfmH4u0GZoeSc9Q7ByE
4VAk4kZr8VYi5jY0u2BfaXHFS759xFUjgfor4qp7XNIIjnIPOYgFo0x86oBp323l
hR8EIbtdo5I+mKc3uXz/aMWebKUcgmDZ5QVGLL1EMd0QhwIuenL+lFMauYiEuPNS
kb0E68JrG2c/0ewzt3CS+fxhf13brqinkE+fyP+wTbxi+jl+lXPStjmrUV/9YDvS
6R4UdBAo4y+XecG9iZy86ar7pc7Qi7EuN90u/C77o8R9rdnz1EuyuHrmNCNVNU9v
e0r4o3kxThwZGermG+Vlzon3S90inbEgAY40GOsRTCgkNYd11q7f6BNBGkYjJkea
jCCOG2raFS4Mxz2G1FmDeJVIJ8OKqp2sZtiZbkq/pybrTJFevuQloMiawR8ptXSF
QW5M0KKv6KE3rBfPS2lOe2OO8fBH5Q4f9y3Dq/sWf9as0oCqAt0BvlLApWsFLCOp
X0BSo1fhh4+As1MrUUkckwJWszO1Avh9gIm0Km5/PUxM29V5c68X+pdKbfkF6alp
XjmKXsiAcEjLTQPaKM73S9A/YAEh9+kbmrJ7+mwAmwAtmMTPXqi8D+G127o1Ninx
Q1GdxWy8kHpqawrmqu9OLrRtuxXAFLDIklG3CO0xGHWtL3LC79Nw+vuiQI8disye
HyjeFgXS9dTyC01Ce6rdibZB4SsOh0Yi8ATPyIuFxHYllBcTa47rv2aXmwUnKo8Y
9EiNsELQOp1FdqP+jjdlaRshOBzyaj7f/qVm3Go4JYpHVJC+5niJ1kqq0BOIK3/0
zfpSKRGBmIYcjvfIiFo5eK42TQoTWCnChXAS6KUSts1/hfD2SXJwIjDRJmSImlnG
SGTdMAQVP8+C9xjNoxL9QXVB3ux72sYTw5U4aN59wYvriip+VWC5+PqHt7ZoQx4l
6zXms51JWBi4xy/4En/kpe3s0/6FSnp9UxwG+r/Sg1oFBodXL6UfcOORACE2jyP9
axAKyrXxqCy5wazJURFHFyjMMo2uEC/tK95llPNyiaOOpSIuw7PutGHpm6+lUpJk
w1MqdEOAlOlXkDkdUZaGyHZwUf2W/exVhwm/6xf9aYpOYIaNRSRsBeSlaVYPEQNg
gZ2wMVOY+KWjCgJnUuaYIUUdXxPQziJLnd6IGRf9Vb9JZNuu4jcW+TxEfMQshAny
dtW15QfO5kZt1CHTvtngJOZbDkgrqHPx1eSBtTFUDrfwTWHq4tT6GXXuIGU+qQyQ
jLaG9rUgiy2CmzBTxREIcCnatPRS+welHojIojD1Ka3gpfpU5LEM6bJxL3JGfsw3
jCcHIXPo0WGrLsbeZY/QgA0WElWzXoWdjkSiJZViVlq9UbexOWymbiwASgycT5qa
5ABScd8Kz1AxooqUSEs2awxveRBDxyLmNKRkPahlxJ35WmVQPJsBq45dPaPDgR8Z
GIm6oaV+tpq8ptcLMY3VlKyoCzhS0/V/BBHjqoaL2rvj5szloTJmmt4+bTVzaVHA
tHoi563Leq0cOOXVpq4f7zBBda5cVXOKRGiHGbxGWj4q6pK+nnvQVOIFJ2GB/W6d
4HpquZ4a5zr0/3kkNzzTbNWMEDiKqpK2tO2uMAuEISeF1tA14W+jFUS4tewz3gMu
mIdCxrzk94etCalM/h6A742wuG+LJrkZ600sOIsKjE0Wen/Mp2h5m9sPjUwKp5fs
Q6b4U/LFkUOXopP6GPH+MDHU6WOWJhtK0X49TcD1T7AbVNlhCXm+8nLLC+5Kp6xp
h9Dvl60kmeMhghxbVjMkm615lEofBZeH8Ota5hG2V1vqjTExz1OMsKrzvO9jA44x
EbKW6cfu3nH7ahJhrF76xBXZ1WQN0Snwo6Omt6puUbHkxbV/dCVE6Embe6B85avz
A5JSQPBMfD9mI84gSRInJWKFkyXJCJFJPhmiqsS4mq4sYVgy+4nM+ucKTFkvhdVh
PonlGIGSS4Q89kDhsdFJU16z1xa9HGwqO6U0BGeGUU2j0jENgj2x+Iu6FT93M/hM
UYxypkFO83sMxttBec7cc5URb/AR6jtjWZA4iP07EpxUsSO8KZVxf/5uAlG91nlZ
4C+lb1ao5NVuW3EcuRRcc/VIjuNS2C5Jg5A+xSZwiVrRMoFNfuPpy6UyMjGown+W
nsadKL2/BUVz9h5fu2z7J2GpNpsE8YFdDJcFY+Y4Ks/cqbeHUwEOs599fIuCQK2+
1rsp8WWaDmScy4rYq0U1ttSjrW2m1K2ETfdwAB87rWffrzW4Ocs2KRSnVNOXnrN7
yDNxy1oPxB0oxC/H2JFDUY64BRdEN+b3w4mRQrCAd+rIR4zxtvZZ01jIJqtAhfHo
/fc+ZOXqlwBGqocQ8/RfU7wMSJYQbJroQ4ILuUGf9hJ5PBcK9GWCuN6EJuKStZj9
YW3denSVsI6WBmKRbsYHQzuxKIkWCzjUJ2GeVZrCyQpJkQk2KSAZw9mklJRMRmXQ
BS/GCPI7DKKZHpTrW31X+3bFcbxhuCBwCwUtP77DiH05t+qrPANRmNTWR4jmuGmJ
9Bm4wGgW+dUKJ9aHaTtlCb9ymrmd5roKIf07Hc1vrJEy62avKG5PtP/JPagrsMra
4ZN0e6tiTqqG8b57kqiiFMAIl8gZXukeSjzVAeSvDFssBsdbN/j/wGk8k+07oNMM
o9lENQnwPXgOHiuKbMQwlyKB/IkFrDtoNGFPDB0LoOYelQw6kwjgqkV+YAP+vLi6
wSNm9EV/ixX6Cg1Ac6fEz5yRtjZZlDZC9aiADnbBECo5TD/MNUA/TKC+mXKIZelf
5zuGvNODUYeYwQa6QF4V/ypRMYUVyhM9FJgCXVEsUZ3+ff/Jc/GdPiF5fAsgtwnM
vqW0uA1uzQQKMETvPTY9F0RPUeTtDa960Xsbq2JJ4INevfSK2b+RQVM4tgxIvLVl
0ScS7BL43nH1gnrfKbRW6tCJ4a1bo/7SPaN5BDdx/NiF69wiGUZ3ytA5OTqpkzvC
PUQDicAAKZdHK7qfa7guinAxIquD0ehjS9pp7/X0grozEc9JfvkymPW/a7LQsiil
p9strdrKLS0m6gp1Z1eJGkdDMsbR9Z5Z2luSLZsSO8LBhkWxHZzZ+Y9a+b29dnLB
7OAAEqIao/4bAIgDVRaSrU6rVffdOX1M6A2e/W2GwAgJzuDFbaS0uMPMVxVyvh6Z
Tqw+/QQomx6rsG8gR2qNRKQc/0OmKSmZ/oHAkKyB+ikuQ30yTkX5B2rcHCnvFBMv
7GP98rpGmkDnSHjQoJNksgOOMNIZFTcf/Na6+WY/M6JLHMelDB591XPV2nG+gBQ3
FMOENblcsvpaq+fLKWI3JPJfoYvVYBzn6cfbV4s0CTozvYuTTBBGuO1UWB6I/IF9
Se0RkKbt0QW07JzfXvniN7GupzmZvHoGKkdfPul/hQcn7e5hppzgvSgFK3hiD3cR
NssIYI3HQ+IgXm3w6JxXuaSMyOBVFhj4o9WE4Ttovhnlwb+LAmOS+G+FK33APyi8
kJkOzVPCDBEf6bBCoPoLIJXSGCwYARwD3IJA5bMpC3cgyIXwhK9ePrNrsDXTA28j
6bgRNri2yONk36PsWPJ9pj6+IAFqRlSAjrCWovAoXesIJWHPDD9lM8ycTCunn7jR
39ORj0mcBaJuNYitaVY4oU7XghMDt6i/wiNiV92TkE8ha3euDdYt6iw5JaTJfVQA
S8pXQqCSMVPclobF+xE+KbNntceBiImJ0XVv1ezId+sWvMcWaUVo1fJ+9jfxSSYW
nD/icXWAydZgdsWIZea8PYBEcyKge8wVG6f/NNMlpS8FHLj2zOqloLWxTgtCldet
uWR1bwdG+YYWPb3mGmLJ2n4HC+oYwHTBitwtp3MRAg90gmg8Wo6BrmVdmk6txfCL
FD0RmlT0dSuJR7m90ONO/hvZ1srKyWzT/nHZIrzh1aBiorz5Gbib1D3QAnLBmhRu
2feStukXcWmVrioWqsXQwHaiNrA2NGz/X2mVVNtuXzQbA6lumQ4DpWPzYqg6Tp7z
1vfHGDxtAZGStaRv9YuMuJ/2ZVl/Lz3t3dcLG6ndjZNoglKL/RXETrdIjVHodgWs
yY4VIjVMSpdhkM8a197cZiDv3LOa2TFTBFve0hyOs5tmwWTbbD3oT+2j85biJW9i
5lFw3AXyTGLmgYLfba6ZlGKjEaEHnrt2+OabByypyvJkrSuNLqtpBM9+FDK7HQq9
gEFekFGLC9imrgwcEYaznUW4nafkxmdjAbvaQ4KQLiRzeICvm+RRj58mszRbNfhZ
+J8v+mw5vJgugFCPVUEFXI1x/2H152RkQxyCa2BwKhaWzl5izeMai8WkmCY91LyL
8Tx2SM58oiqq5Ung49REzkeZaniqhs0SaiMdU8/aeoQ4OeSxzNTpPcYA8xJRTWEZ
1jmxKJHBU+dhwHQ16sj1SVX32uIhpzWVIXQa3WoAly9x1BOyYqTpezqRbRse+OjP
QmvVCsp9jbuZaL5IyN8kyjGZp33Tx+snO6Oh2Dkngs3hJLerZtNZldEOCw1lhh7Z
p2fcMdGKETkjkYRqSAEjN0JQ/Fk93rd9xSStU0PhvDKbapd8FlDu5feTIVIr84LQ
I5gEDOe5JPrOlg9D2DdnaLL6+dcZ39fwoQhA5vUXDwX9pn5Q8ykFlShIAmPH2C/r
KZwS5QTciOPA842GNSxn429WyGs/hQrSsvg+dY6bFysJZFJfEnptNOy3daxcunq0
N5hd+H+1Zt8nfiqkak48jRgZsc5cgMMir52acv3jbtMfGTfoKyYa1K4/ZdVxu11f
J5uju5/Bg34AqbB8CXsKqo+ZK7KfuMNFODQUnpfA7EkG9issbTjobWBoFtDi+Zj0
Olh4Of27qwhdV+6YbXiS7VwCz/LnSp3X4jZeBTmmqD+W/dNrucNJQ921r9TUKAYr
+Bw7hzNKS84cFd3EuyWViTDkPe2tX52c+uIBZbI3UDOWfrQN1iRdiawZsjQjO+Dd
aoyG0PdNalEWiSZiozW2N4qnq9BFvTNOoMVCZ/qmz9a8Iy7Z/cS39kK3wlOAy4Qg
mnt0/NRTGYIsxNH7l/yp+spDXAc2j/7006S2qOY7uOhZA6Asvf7lkSLsRzNFXUAQ
ZvBW6km5s4TstJZ6qiUsjW9QzFy8l6tjVa29fd5H22/rs3i7bj35GL/arfOQSu4x
OabApVMbqKA01WiDTTVnW1Ui1Co922xa4s2EbdFUH82J29qPi4J0ksnto27u3nhr
BGixhsEvYF0ZCWyeRqN7hA57JNT7ggolNlZLBX32qgic2KqyifZ2pDfJU9Ds2cWD
LIw9q8b5eVAHxkLHe3uUkxrs2s8OU85mnbG2fv9w9p9YndTStAG7tgMCQ2AvQJ+h
qHxQKeN8a338ZKWIP+7J5fAZun6Jis77sTXcm6sHYHHFwKhFIHwx72bd34Nu7NvC
VInzOE7wBE56WgvJvP8jinrE9ZNmCCI83dk9C9NxbMbVMmNOj9APLclWzEPLhFKJ
pJbQ7A63LXVUgco9RLCbLXE7CrO99lbtbpErVE5y/FUUbkckDfsR+9QppjoB1YBh
lsDLXbuhazjMm25R8lQI2LqTKixJpEh3WOEaWYYJ7mfZgbdoBiDGxRUJBCnhbGlB
bo42TSz97yo6b3KyNJxKnYS8+d+bKBjBn0XBdmhMQgw=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EBpTJ9JJFdT2w69Mk53YW+mlp3vHLVSKHTe/1pFDrcKJicNQS0ycQGs5a4DR+9lJ
YHw3tFlV3Gll1tUgKwSmTxuKeZq/qMhCxDuV2WEI69+y/07lLu7M1n5UXj8uiQWQ
exmYdnMy13CCnabytgepB9FPhcRXS6nHbEBE9W1j4zkGsr4xc/Ch31O5SIaKFtQB
5EKN2L7WM2fbqKxEf6wgisaj4ET/xCrFyunIR/hhqWjqfJdEDALsTtuj7U4lq0MQ
v7VgEvjdAgeOvR+M617LDo5Qzv9J4G+If/HuDlJ3QFzOtUqgBEkhgjgck+dZNIlE
DX2Mzw9vZuLUPrS8LvDwgg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8032 )
`pragma protect data_block
fng6nrdrJjb4iGmVc/KLGqvOmhd7NC/3SdLEycpsQ5uPFRUrTJuIeDRlXD9qJOme
tlAGTdNEJ8SnZ6/JtOuwCYD8+XddoikHwvzr85/Bcan5j3HiUj5yNf7NtRuT4kVx
P8wGx51hxOUTILmB4YIQ7obexRRWGfk4wFvVZp0VNyINhFmtBlksGyIYuc9XSOVU
yIHweNr6ZPKT4u+7A7sEj1lLIe/LAS1/yhLpUJoGTYXDL+MRKg4VPc5Qc+uee5Fx
QzWGCBADR6RPnYl8GwQbzS8fsT743NSdaqZxtpqllQwaIKA/VeZB172EXLi6hiTR
SGB2+yC2J1vQhuRDG0BCPzLv/xDcdNA7HQwwkMYwlr39m5z+hV7rb5qf0gzHg4m+
CNJFeK5MSvewhgPJlXi952fzheNRqtlTPH7IivqM9XpssvIUOHgw1rIUIQnsqKFU
edjcyEJ4eK5UBtwL85vlPtP671fkoYZGbsLpsTl8VhwHMNbqbY8yvsXw+eXwJhYc
TXJDWJQGWtfTx2FDRmCI8RlxMyJkYGvEaZq5Qkoa0km8dz0FDWDnyKwh1Ecdk1iG
Hs0JRWaPv/noKrFS3LqRXKcQ8e4ptW2ND/g24w5wuqNNLbcQOK+qLLEh55VF8dtQ
Xm0TFfMQqbMC6fcG4luGoSDV4FDmxhxUam86wzvFcUK04cqRFmOCqxUbTOJCv0hC
W5/yXInaMHlo90QKNeW2dqpYf6neL62j68L1cshMhT4mUvfXOVJyrKNx9oYnSKyt
5ooHGaxfMWF8ppu0ek9tyFFMN/YIe2y0nKPbYd9i8VqCgTR6fRvQO8b9Ceq4p7dt
RodwU3uw4DOweoOn0aQhFeZ+JuldYI8TUSTgoMaMvZcmnCSiWJUzksW+2NNDa2pm
V0BJxBBmWkV0jd82ilN6sYZXCy56OowNUlnJHJ3Sa6sKTrd83ovlAotjsMoGHxeK
p845GYrw4iVPVXGoUbJUIXcEuZQnRYUZ4RTQroH+chC+rCj9wuiG9xzAlZKStXfo
IAF9ZEm9BxSHOtg3hWcH3cr+lxRLKCw5e3PvVD7B/vE6Ql+ZjULwzIT5bBgyUmy5
6oorQFtYW7Gpmbv8YExDFLRBDWc3s1IdFFJG40/sjZuEpL26RJ1ywNi+oP2Svry3
KnRLJxMfeUWZ59PdiKO+swR68AjwMdP8P8N+FOLlN3gfm0opBNDra/HyjXDcr/Ea
BVRztBEW9vQm29U87WUnXdjyUcdV/rem3/wEstCGPpyAtSgEZyGfEu9TeOYZB33b
sVnz1QFih9aPYlzmg79WFiCMXEJ7riS3Qrpg8182K37xVNLeqqO2kss+5uFSDB7i
biwFLFSrgnuvyFIhvcZ5SBAxoMM9lUtVpoM0Tg52QzMnFlM7fiIzodgrKBo5rPxw
50zAQRdGPogB574odm0xwJZb8jjb2oboAl0zFFUuhH2MBdhuXFbbJftzZARZfjc5
Mseux3syXHxbt63PtGpWLnNdKBmDySmS6s2iws7t8aYXW2PAIt0Nkmqqq7pgQNkN
X1j/yJlZgBAiWo2FMQR4cu0spbfsCwZPL4ot0UKO2WqJunb3d9DfXd7Q419/PuuV
0hFU+GCFeZ8R/IZ5N1j8zkzPKaUX62WSlFAyvmyQgsTwfU0qN76VwoTkxLxrnvbB
99ooAzdlE1oS/SBcwReju++fcr/BrlBmkr0F/rtqhS4wo3RD7SsXNih+mL53qKox
FRjrfSjrF7Yhej64RBQKxKDSlh3EKgoLERRvO2W61nWz5Vp2vUP1uTPM8MVEg5CG
j7UZNqfn9HdmT+3XrWT30JBK4QcZyxK+V5ciZzUa0fC1W7CrF0IXwN/alN2HHgfQ
Vdr318RITfsc44+LDaqLmc5LPi27ynQyTauG1AEt1RBrZklxbK08hM3Qf3CK7x2z
LXYDTnNf+1ZPiUL4PRhEkUsBNe/JZfHqgSRo9CXDE6kcnQHICmSz0L9yObUTsCTV
DwHHz0DfT3khJvvX7TL1jDjlZhKrcRLveMGKCVS5kZB2nMfUYuSm8hBfNnNXVohS
GL85XWkaWN2mNgJ4ZhlmsuVCe7x03w1v+AQ+57oEh3A8GN8IICXEagse3p7ntI2y
pcs+h4JI60POWiIJjL/PqpVxh39t3t+Xgb+L50V04WR6LD3SxikwFkwcS8b9qSzv
wtvUX29VLm1TxpivLGiPETcmrF1RekWG3OLSXDXlbWmet6ecCHzGrZNlHOwkIRhD
UQVawu4j+IOfmGNZuih9poJjl1bBZPMpwzcUCmIo9DPyuw9B04r4fbmj8lVYMhOl
KfFJmx4z5f8rl9KZoONYZeIIrKIPFgYHQBLXUoS2hyBvLIBlEk8qvihnKp+4V3W0
d+0onEzoz/+NJdoXERnNuXcrjPUuB8DzZ5ba056Yc4ybUA+6a+aZncUX3TLI0fnk
FHskMaXTzmoDkJfk70gM/P9HNRHeWnGZQ7fwUCOGvg9GdPw3aF3a0jz3zwb5SnvE
0/0YF21FrR8dLn+d888G/cvIGiW9AAV4YawJSGFzARIPg8MkARjzYzUG/wi1G0hQ
QkNZdTn3DXYH9ZbwAuZ+459iID9Qu8HBfI2Ds4euMNMnbNRlAOqB7TwT18IPdjvF
jMEkyw6fL8covaQJNSQApkdfFynhIqiWt8ilu4O7XfNibqz/nQOoAifEk1IdYzIL
gTX2Mdy7zgjCmDVsxoeXY70Ass89d3N1BnS3JHGd2pl7Law+KOJ/2YS54wws3huR
vUeQIl3c4m5Ul7u+Yei83qNKzhQ1Uz0mUybOXJ4moIIOa8/tikpqRPYF1iNPDNMG
uSmtGV1b2b8y6p6H4aJ/7Fy+Tk3KM5E4u+Lg6gnWCBnPGuvh+TLDPukSvIkbNY2v
J+fJpG9QKVqAnyzdOcYAC4cXmdaYbKhamfhD1iy2Ew9gQoUDfb6nsh9shkmCJHGP
f0ehonqcI+IcK0lYHOm13q7viamtJTMNGhCfRmJ1JyKAR51VdCB6RROJikrQVxkj
zXcAX3iNvzdyIiSosmbOeykACYW45905uoFmcgqwIUbDhF+oGhiUlo6rKIoL9nMX
4dmSu+Ql2jF3JshPTdQASdSjMFjBA2bvcJ12ZasfDuz9s1qGhhV9fwcFUj7ZD7at
ssj+wwGBZHTfoc1+Z2szJdAszsUG+M9fpqXGRvApzieGhoNnq+FuaUPcaH6512aW
Sgq5yO8MukKKEBCt4+REQTXTptmcEC9oqnpB6t20YF41mZPNdk/Rs/n//nzY3ONv
60NNV2MEqJ0qVQYja0lg6rawxLoU5wxbBOrTcyPswbg0+z3bdQYu9PB46+XeKpgt
KK1KsXpXN6qpdHEII+NffBvvwhGGfW9Z6F5C9qzvVhjTd8mTwiF2GII+90Uzs0FS
I7tagZgh0ZpLXBR5uJrjaL1CdxmBtA7Bpjq0aU0p0McuCGe3RlUzUooDCEcAtMvp
LLY+M+EEjywTK9Rh/poqV+L9D360HcJSiaUFm9lBAheA4NhBZdQ/StE1/8/3Hxwa
EMF4kqYDW0OcgsBE0PiYxa32Uf4ejX1xkqY5UrF98LWfGQojIDUzKMCQefO2+tCK
kC3nrS6SEwGsrGk3s4zXqw1/sqSGkaEypd+BEZVDn7U7xJMh4DlAh2dt1oILbqPW
EOjgdJzcxk+n2VkC3AkRpQ5DxKX2RB/h5MG9MLdaYiE35d3xuyawL5JkObOQhc26
gRdbZh3AMBTsSZorE9v9XdSUJ/gWltehp5dg2Gx31lsWfbAr0oAoULqCuqEz2e5e
mkmogy8J2K6p23UrqB2zevNbhBs2t2iY+H/xVorZnKOiPMBE4b92VZ9pIjGWKIPJ
zdjNpWVL/mIv2jQPXzj4iFY3lEpeeRofsOGNQpCmlmjL9WEA5ZZtIu1ST4csheh8
T4vw1s44+QM8aEOD5H/4IajxCuPbgbTOU5RO7ID1JRmSbRIflkyH/84Vjctzkdcb
IWvuRwi4cvNaachJjsnhFi/NutMncDqEwLwj6cyWahp3zvL7mOC6BFr6gEwfXxWx
co5JuaPftJCjuSPjt2dVtfX+oCZn8ViSNvnHSaWtY6AzQztG/LYydqaTwUnMlFE0
QppEYULCavtjNmK67YRpdPh3qWWrB6q+rwI5NsO3Fes3cDY427iLQZZXoX1zQR4I
BLiOCVbMvaAHQKhK1Byc20kScjXIXpnOymMYmMcBqPUOLrLQThnNxUrBdOikUHyB
KSFoKwVSYJCEx4XVF4msVJTMC2LCqLni2DUQwiI+q47599rW3q6iWc0XX4niYuCl
/REyq2yrF4k6T4bTlqCW3FagGhlOa8hfWGt6Txu17P+MwjfailtD325owAGVBxE/
mADFPiZGxkd1sQQyzfTqNALdrgKt2BfHJY/STtUATSledJYA0SCKTu3amZBp9w92
6XwdlhiFLs/IMghLaOmi0eaMxPIQEwBCqXFlRpZlmVN18IV+iSNSCQ+WPQFZ1JGo
c3xF5Vh7IiBjeflvPhcGoav6YecjwAODE30iXBmo2W+/o4TI+Hq5pekO3A5zTovO
GkUTfAesIhDYoIQqR+/Epdbd8d0/dFNOyM3COAZHDaHop4fIpTq0IhgY59b/KTS5
gRUlejRcUc7wp8DA3aj6Z3AHlmxni4EI+YKV87d2fkY9vLKekZ/cXY9kJhmA0c4o
EKLmx2BpA3utQFRyyj7QjyIgl7yjso79aZ6ovLjJXrpZbIWrGHG304ZDuTuz5up7
Y3N7sLtOFqGIZ6H73XduY9I44JSg1pR3rbxVK6NFNgUyh1N4Mf+MI75D/PqaDTVN
1FC944SUmLRzun/O+AkeMoaY0+JEOWD0bSuxE8vaJDC99DK7ienbh64dORQISBdy
DGpZOk0I6hldubYg/CFuO0XHEKVpiQ5w0LE68zdpbJ1vhQVYyb/1poS04oh4if/U
WpiOnbgC+Zg5oFvC4Ow+PaQ+Hzsss1qUzXtIf5WB6CbK05RtqUdeShYvXUNYZC64
GmC93WpGGmBeexvlunyYr66OAL0nKE8MuhdV2ofGaFNDzUTBI9odCDsUa4wwelCW
+1ISAJxGqelQyJCNpLeKul3Pf8fZxtlQGMFIR7g/6PfTzggo7lFftago9JWDtv+w
a6qic9O35fB3oR5SqE90z+zfUQGFx6Ch4oGjB9jzjUdclQss1HIG0D4SCPjBokIh
fEre4rxpdfiwiqvtlnTu51wo8OC/lrsRoXg09TWq7sizjXPZZtMopRV2aa/USz8l
4nIDMKK7Cilv19CCcnwBDG6Xeg8rTbX2prVVW6tg6S3Ue+5/Q8kIzS1xndI86Dk/
GVc49EtHH+brUBQBfUKGpY/dumCOBQjK6k87b/u603OPUTZkMC6Hof153FVXJ3DT
VHVyJwDYHISJ5w9eylkwdMZ7PtMxxvtCYNQiO1IpDTtnCcYgp/z2xPAuHtNmekxr
DKaUKGVczvBRQ5r8t7ltrbtIaqwJwLNYX0k1kmPW2pxRMCK5eDzTkWIHP7Kw+q5F
WDSHmVrUdtT1hCcx8gykgWiSqpyhu/Bj57JVeKbuX72+opakhupq1fQpQCkLEyjT
QH4uDTTcez9kZRP3L5J0eE+/czOaRIGEAz569rcXXMAOLvyQd8SKRDUZYflw8xGk
jlOQxASn8Oi7uLwsev1ffcARm60Hn8bVdTQAhoK3pnmCfF3j64+Prq+ObGZ745DQ
BF1uSGR37RU1bzr1cPUqZiZkvtF/5WHYL0y0vdfb/l0ZfelvNzfttQcnOUGShkHz
ORlBkha6l2Enb5BQ7q5o55Ab15JOsmiKCAAmMuw5ChW9JfaV6o+KVOmKSyoGojhK
4ZQKIn0UgJzgpdp6bmRoUMNeXks1D7kDjtMmrw+oUZ44zdIzAJiIiqmb16OjKzXu
rc/BsgVD+0AAHXfVsK+JwrNg+Hd7ySZDjC5q/9UTU6IP3j22nagvt0gRTjMMPXKo
2NNoU+UougH74dF/fczPCRNbzkL9ytTnCL2S8RXElWM0KbebBGIYKV93Ph0RR6mi
xMEPmvqRsgUF9SrFpMN8ESK/LyBiNE3HVGx6vc2Fm7/TASJtfarQq2++H0CvHRxT
gdwGtI7lvJazPGU6hUH/bce2BqiHlC4j13wTMq5WfWvxzKiGL1yIRGh9hGTzzMYT
V5do+6HtRqGz690dk4YUwiy+6uKvS/rtSHqzwyrS156FeVK5/jSIsQBR2GQ36aeR
7/kyhQzM6UFtAAjqDZyejdR+suOP2OI+uFpsggCFbTITxL0I6qzY6bVpZl65k5Ev
xcgzven/SgfW/gSGDJjK3WBoig81mKMWKHG/VpsnlS+NMeEJ47SB/lQxkl/9KMNM
IGHoe3ITiUtY/MN5dWZTsDPu2AqA4C7OsZ8klPllU1TF9bIiZ0nA46PpgZteLk5n
z384Kf8biKbR+nvMNXkY8Lya4V0BYTUIetFGQ5tmp3BJ8PFgtJH67P/R+xrgfUAC
nQAkr0QtECgie/sSm1BaXUAgwIfdJ6meDSxnzdpx+FM3+UNqzmHi4/eEVZW6fzw2
wkiVUVomPq7zbLJ5HYFCVakZMnTEn7VkEduqSk0nkZKJ/XrmndxpmCbHwaHKopNZ
/7Q0l5hK5dM2iaAdSRC1SfOGk2Nud8bxruXwxa0GyYT2VmrrcoVdQYk7U5HdgqD5
kKOSti/evhlzTR3Vy+WSfv8iZJ1Ca+AcdgI46cU68rm8JkfUNtns+XvEUyajOMlK
sZyg9XyqF2pBlnuxcACvj6Rpo07dYMKO55pWF5B0N0TftQb/BQw4XMPWSq3yBqs5
bX1QAeT5ZjWn3z+JloafEtdIjXB7RNLDGAvfyLIm+1sgg34DOzQYGF2YlOAbguwe
P3SC0AZOkiJmuRLF+BriRYs7ptblGrDVq4f18i6MarztTyXJhyRdK4Pgfus2QTt9
PX4vBbO6Ooi/TIlftXqa9Zu4W0/KBioR3SaGJSNJvdSU4uClHBAyRgCrOsyzghID
PVNzReUwxx2W3ZprB/GzulMEUnEgiPg9llR1akxdXwoLSsgWucb36qjbcy9CQcdM
K1CMFf4Dz7s9YZnDA/xj5Lj7Ry5LeQ6KB9cA7hiBkf6yZszdB98Vrm/L6t4sbQ5S
hd1GnNwFWcJSBmu7UIPFitguezhEktsm5EJq4uCkqgJWHT6WboU4MG6pafhysvTF
nfV/D7aMpf5OGKcmXerqRMagPaqex+bZ6vOtsl8dhnIZFFiaj9RZdgsFcz9/nkT9
fLIXAbL9O4G8AY+URBplZH4rEiUVd4lrKqbLI5wvZSOKaGH3zm903x2XCJ/f0QhO
0UuiTapMOWMnxPAqpF+XZ0XiK1I9Q2fBJt9C8yAr3vAijnLOapqhgd92Zdzjc0LV
ubVTdMe2i79TPQHbIYXx+Ebq/wKkrAIVUPfUppkos+ol0/spqS3/ZDjRxo8LURge
3TUKo9FTuMu67hNcpbSJSt5Tnk98VRYGyY9vFBZbL0BKC7kw8xHUGwREYhJ7RISF
4Syk7JsR6s/pEB3kWIHHVTXpPxl0dNwSQGoa2I/X+HSzjvrV43GL/4uXI5YLHMDM
9YzfOGUpBKkk7NcTXacnPZ6ewDTqEUGLxeLhv4XkSXcq5OuMJLzONpF+5ga/vc9M
0FbGgGxgsmas/kl5mF2ZdL9Fh2znuYdNDuhJm4JI/4DK1UYegdUU7k+/+RmkcsJZ
ji5m6XI79ApAyPtxblHRjvk2ffs6yNL1fsv4u1E1+83+ifGnkAuxTyzErcd/Du3L
ez39F6/mLX8sEOv6Nkt/eXp7rIZacN3HOKYLBRPRnTQwj1vCugLWbPwzInhEwPWH
178vKcHzLDP3DR1cwsgaowlOfKcmDp8mOX43OP/lsmhWFXTS4uHYoDYKkPLSB7a2
o80qTKJK6c1bRqhda82wObDj2i0iRruhvpnR7kXZAle7PJ/X5UKHZOAyigt0ZHFX
mEyFqTNMqcRdkak4/SigbmrF6Rega9bVjDXn0LWzZMvuRR5ky5MWnlq3DpFty6PA
P1mQHkf4UPmRGdqJ3RI2rdbHD3nptlDqU2UZzYJIlZaSdRvX3TCcE6wvfcOOCQR0
nN4OToLu1loquNccj2rMzMkrVBGEp2rY/6bpB5muAz6mmKS+BWbr9jdpDbJ/xOfw
8Z7pJyTwCa0vgm+uJ37D52c5Js2j3J/5Ls6gp2cvCxe6kW9EkpCeItdJ2MtNidUA
7cJWNupYHMQEHCcW3FLhNQ9P35rejDShM09N9BAkcuUS0FQbyut/nhwPamCd0quj
MPx7fdo6J/Ast1+csJrT3w+ms8UWUDcll3pwg7ehY/QUvLEnzWVfOOuKsZf1tl8v
AGFATvd5s8EcMV5tbFdPknSi7eLOju3crUUxUMr5q0h3hk0/WemUknttX56ORrP9
hMmS9JXbihhaI4mc737tksmLox05qXXvQYUb0Hjqvz+1gK0zR3pcO0gbI+mGfL5p
snHoeZMBGkFbr+QFoeThE64SmJLoqH8g/0FJu0iGCGaZBXnWWU0OzBogeOlJ56No
EbG1dOmKIEb7B6ud0oM6Fs9Kwja+ndn9M+w8G4KX/G2JUcLXdTeYnk3LA7m+9BJU
P4yMKHv9fnvA1zQf5Z9xPPO/hJH0nC+BCB6BmssJjXEeM/4UR7HIX3fk0UyDUyLz
DB0whrEyWkGMl+70+QSGBr2Y4aUc/0QacsevxmjAkdPvbLhrq3EMrrGMMEszTheS
lZcLgcBxTnbS9kgT6MGH4qAkoNjJu1vL/zSUvnnmd9pzl41hE2yICj6Sz35Y3QUl
RNbGFIN6FzP0kNV7e5J4kz2mumN9+xUGibUaaWGOhQXN/kIUcDYQMr1p7/Isgfm8
g25Qip3Oej7kY8bcm7XTIDkMKve3T367PfZpUL7CqVMfiSThF3/M2gGlKMU9bOeN
bNrixXVQnemITT75gOcd5BNFLOwiGybbXJpNdnRv36Ynu82jUWqJsF0gsRJ7nR+V
gwJfiixvdyQG98Drot+osVAruVw3QG8GAevCwgeyXrJNGpV3M+0+Oi4opfFVwSPZ
KUkihq2G8nzFIUFEtikzB8tGOuxq2gkR+jANUCASDuLUXZUj7n2VpHmMS2rohtR/
dGnYqR5NwhrLB9iG5o5WaXup867IbfbMCBTnONaIlLof0R2X+Zkpm45s/zQUJfqG
OP6yyzOV91479Qsz50bTaDKL2shUVOiyhu802DhzOesu+iE2U4BmN0+h9HEydUG7
foCswnYK5pL2qFBr4pDnbTwOod+dS7ifSwBG1W3dzRqGVf/IGv4uM7acD+B4KVeQ
JN49PT6UYm0MfshZVT5/fPnEkljdEdB8O1XaukZ8ELwANc7ZeWfVpEtODpdgwbxw
bDSitdxcSIfndeM8X9WINSq6apJjBRXdtOBprCsuYsF7KIAWtk0gd3l40fNlw1ro
ZIxdvBqLV824L1fRI76OmvEmZG7YnEBiI4bgfYZL7ZnTFxIDHkcNrXGT5uoXJGIf
dCLYMiiz1NY76oUD6MF0Y2FDjbYKzDN1z4e9/MPcUbIBdqBalmPxtE5A729pfi4+
t16Q1CZ2HwxkMRmSbb4VYWSFSrfIUf2ShPjoZbwQ69RZlJ4fqh/LSHhvrJbLcer2
HLrUu0a1h7khnAVc/lgmSP/SWydhnC7pbCdoRK20pOc9b1C79Z9g0yWEnZMkDZDc
J+WeGDoS/hhkxE/yJv0krUpdmI0SzkgG5DQ3liqst3Y3icGGU4wW5Mp+QIO6IsCX
Og5JoRlGBi5VUDX35XQn2OftqiEXa9s4buYeD7AzXKGC3VcdCuLep2TeT9uTsAaD
NL+9gQ1wiIYy1e0/CFdkqFdvfUYv1Vg6mThBOzoh5twErbnAalKY15GqAKdzkJQB
H50WUvqwZU+cStOmACJJZhbZ5yw8yaOhy9rU3UH7dr/XPff0cTVrgIXJEYfjAz8+
o4Q2B79xGHXNgesE+UUPZxoxyX606dYtrV75uq30YRgdHu4cILKeZegMFfPup+hM
L+ioqvmUH66yPRTsS0JiCB9BhXQ0Fg7f6wYAun9QMVgFlKbQvTFHlnAX8W8TADyU
KrSRlA4b2fyYpwcVC6IX9yIJTPzyezUuqTtSBIRfvihaB4zC3MjY1IZ2bIY7HnM7
nNe1H7QFwPztcmronwOnZRjb6/e93+BGOsCt5hq0KiOKaZHiQvz/hdaUIRXZRxFZ
khC2rRh98GftUjlewjZ+Op7c4KhsKTzlOzDk0sYT++4S0HHOh7iRANlOKG+vF/xG
eM3NN8AGjCgx3oXoRmiVCBGvHR0gyi7PyMF2tYwNNkKLxz3RRJ8P+b/3banqhYJp
C+JGlF9t2dgND9a1sihjS31bIBu9mTBh5nYesehH8Cj15V4CylKqXBcbhZOVB0v7
nSRxqFJoK0gg/uWo1DCD6+IVC5A4xz0eK+fXx0VjQMU+QsN47pVNdGs/fBitgGsp
BazBxvGfXCHnYx1fBwlkRbX1qwuQvcB+BmFr2at7PBzjZBgLgyVTi87qKUmHowZE
caAheoLNrLs5HA3rqodjntDyJvAXIyhpXrUCeOQ7/ybfJbU2opsffEvDgnvPQa5j
rgUXslsXRQ9sCjidSyFkVwnzQ7mjf0sPlJ3K5oPwWNbP6gg8z7h9o6RwLXBSQDnU
13tnGVEITm18S0o3c4UBwCMb7Y8dikb4sqNdr/twC4J4DrnPAe/Q9XjTaKG2GlcB
TJeDWfXGlgsHjFUwUiBMsA==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BI7GNbFSS7QSwNRCIEfEzLpNiR3SPphLwNo/C/xKhU+2nEeyT3CBzuyCvW02Oq58
NINJCezlW2aRFAy7vSac9fkxfqvVkAn1QMv5sZT+Y5ym0MCzSIiCV4VPko7FiOwE
GUxzAIcBth3+X+YfhKexDcCSPthk7Uf8eYjTj3X0dCpq7mElt2szqQsIulbbePTA
irr0w+hO3RGRBsWHnnUUhqU6ylSnS9d8XzsAO40NyQMiPLuB43Gattgo3CEnsfzb
hbtOAsDzGGn8ajWeGGxlmWV8vUsrY46O3WCoMMIIPWQc0LXMthbW7d1Vsrk6ssvI
a16g8j4ilTLt9lwGplClSw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 19760 )
`pragma protect data_block
pLMZC9VnQcNnH4NeAHoQ08+LjCM+TTim31lBR+W6XHKhdvYjm1OvuMVYOFzWeIfC
XQa4o2+cJjsyJMSrTNmsE5VL68FblrsnWDTz2oLUX5cZjVwsIxdVU9JlB3YvA/J8
0cJvVxn4RwsXURLOrHR8ZFR3AeWPDyFkIkFdtfFaYL2pngUBzLoe8WaYRIZBmASq
fBALGkC6T8QCYVedtFo/q/VgB+k3M4jf7QNuFOEF3s5SmkwMxsVHXEkaCY8G+dKJ
e+2OMM5Tvy76lN+eitkmdwgGnctF2FBhtuefECB4BDA3xgKwMz6TtoQkoxjYqwCm
2aN8ZS6N+ta+f9hgFVzlCOuWHisgJiSIBLGoJzDmhUEzFAsYJAkxZ94O10YGfqqB
gsDER+m/TNzSjmrhiH3epNpPr1JA6Q89DNi35waA481aW+x2o3lgu8e0bo4XW5uX
gwnjeUwAKHHKodgGgcpDE/+g3og/VSKgYP2wgnZcqSu2dzzyPWtQh4LIu6ZUXQZ/
6fx78opgOEwycFAu67zmF9giXwGZ9o5HHrSMyVrpDKqA3vI17bqB/bZFmBqj6AF/
JGZnx3PK0tYvQEd/CnibX4v/HXP9je8RxG7OTBryrG6C/4ogoy1KaPyhWlZVNuj+
z2M4WS9j8amD1QS+nGGXHkfLXyQSfE7fxHH0mwAok3PXyMDq39BeYCZ6Neu7FqCh
ziiWkLX2HhLPQbVQ6stCyQGSGCFvomGSBGkRkshy+OddjJtvkzCsygceXInTVyBl
6o5idjJtMMaZuuuSKBc5ZdkI2aLsASNAM0FGH0FEILHb8AnkZKTFEu9KE84VNpjt
DetOhc8xJg91aPOaNcM0+vEGS9oC2/zp9UnqMjxiv/CKT+0bAFY67ic0v4o7SR/s
bQFdk9wSucW3TJ7GUglKTbSDAhmPTP5HNveD0H0Xw3oBpTs5mASSPEd8fxc10S0m
b8rL8jolUn7dOwMggBf4Nqsc15Da8B/geoVKkfefgSpWLKO37ouoniS2DhT7pEt2
XN1BjvrGbgbsdPRk3M9iUrHmmYMxPfz/pEugt23H/Ut7Km5FFuIAF0LivgliddKC
TGyxUdIU1qGVAXEghm/QK1BPoMWsBhSmDNgH3aYk6PJsIuzyrmkXeluOOPxFne02
Mgd9+Ewlp05EfoRwU3ndGD/hWs94hxp9x+XQ8R21OAnZrxsdBunTU3SdUGqqn7NR
32w8+c2H/0nb6u59qMKHDueiF4B8LM1Mxru9qEA9Ojzp7b9iF4SGzeCXqV9x5z/Z
9Z+dG10rViZgwVcHvVHqTuA8F70wZuhrm5c3lTWMgKOoygppFloZp6Errz3+/tPC
pC2+pL0O1PW9aLJPCqH0B3LQ05gyjul9j2c3O4Fn8jK+BuTXdsy+EpYcKd7m2o0s
S+ao8OZgxUVc1SS59BjYdcmxPRJoHfltvqYG51arZuqvFbUJ326WSwxUthuxzrAK
+fJXyCNxPwVsuj9d5Hn4BImclZfffgEK33Yd4/G3ocGENfbVsdcXa2CkgUArRMzM
Zn8z2VlWga2hUI2yQKI+HV8b9wQ9/0KA/CgNo+kg4Du2nRrtHFHWpzXlHyGUloLU
LjTCdZONJ1JfCflLO7a4UPgS/RJ1ix/gPzdQRHqWZXHVCJhXTeFpZ0TIWYz9gGLK
m38tpUmU+MvghWufunNPRLhLooWD9Wsi1G4hxj2/6hpoPlmZLx83tBKaoOvhrxyS
fSgAyGakdeqm5jc5MHjfCDzwl1u3JVJqH05bs1xmDTY73+Vv3RksPlpFUfsfqpUB
kduIXn6kHTIJ2ZwZGPWeRQXFO6T0Of4Lxc8nbSozXO7hOq1UrtqzIFBbT7uezXIJ
E/Lxhb3+FYXsIwCEJtDbM5yUmDTeRpaQ97mqUbDxqPYMpYmsbokpWHKGZrKViEwS
PNBHtACMaDGL4jb24weXLVMA325W2krfQQGBBLHjS/aHSG+bjKaAq+MXWy+N9bBj
l3nNJ1Wx1AGQrUaXohnlLKMSahjxnX9mGHaDwTEedHMcsOiS8524cg0QDFU+QkoZ
SQYbI1jBTDzr4CnH1NCzf/rN+Z15QH0JvgwRjXUZjv61JiyFJVctJX7rbEPpHbW9
YKVXkZDm5F3SG+gpdK3zARp2DhzYsREgMe2OJTzN0QRv5qhrbALip9u0IL/hIFiy
5J1QUseUgaOzC4MJJP+0xIYyuwoGqaqpvb/IaQR8YABKVsdlTySw5rmCqr8/CVFM
Puh72dyjzaUabXRxkANa/Z4HHxmKdieVMSh5D6kQ5na4gGd2KmYWokrhdtg/c/ux
9cxah9wNClORyjVQBwTK1tG3fzvi8CxmBHnRzH9AiiD2z92xkZvJh1gl9aXAqyxx
EAylrS5+ttFtVF5awH7w5x5NArx0mqo9MIkx6Q5bN5Z5a0763zUX01hXtSgkWujb
xzKLcNO6HHzkdd7jclkA4aabTxxAKvMv8liGAoCfKMzm1kcigmHuF3VfqwVZrBq0
TkttmtqWuOMgTJOne8FsrK2sS7lopqiPErStnrg7lUCfwTFkUG71+gipFSeXg6eS
lQ2pL8kFI4xpvy/vaHaXrGYczD8btVaBRYRFEu7gGzcU4VXheBF/eAD/SkATwM5d
om0jP6Sfu1HULmi08fe8chfC/0mqhIpGbiruYBOUsHMIgiU457Ai03portjZpXVD
4SptpLsd67X8sNG89GU76qY5uM1IhYFF28YH8oBtyorsdMwKT0PN9LTVJwBHRe2J
8Ru0NXNqev7/nxoTGcOIolvl0KK1Dp5D41V7mxbbk1OsI2WkSeO/lnWqIzlzdg4O
Z/4O34k4Ma/yZsFBjUBreZJDlOIPgjNGvS/THp2LD2XcSNBwje6LNNRypk79fGKK
xMNYcRU7R1BLgBb/Jql6U+OlR57hrFZdyxQLUCiWFblii3ldavHlj4z+7sgVfYka
2otbixCA5a7JU/WUtqfa0aBAp/gWn75fKM/WhYFGpzDBvZp/4tOXa28bCw5nlBF9
Rhabs823LahmJBinjEJSu+RThDwRxyP7IoMFBT68jO0kIVN77VM2/cr3+gnFEiZU
7/0ytTsEuyBqJP1dwNmi+6Mqm/7qRw0VxEHh+YYX87quAOYTFiRKcXHGNScsti19
Kgf7QsLgDM3+GPcrkIf0z+Z1AvJjAwnB0DAeS7dSmWexSdypJHLpJDtiy/Tp9Fon
mvXZqKHTV1AO0y3MDieAvBA9ixZVrYESHzy3B3Megu3Bpj3RSu+T3Xj4491debGE
jQpFVRXhuRH1k0MzLQJ6jLH3Xphfr+z1j8zhkPeoFaNL02QpdXHxlxoH7sTTBxYH
/kq5oP62CMSOCqBX8nSzV4GYPqMJ1RVoLKJdD0THO48yCN2tt2dE0fHTXj4b27wr
FhLgEu50SiHLD+KFM6MRJUKjhi9ZmgpoteFjyEb6/TNr7gJt3o+JnZVOs1kp/izN
akbLML1Hsx83C8uh0vCX9Gzsqfrfgeg+seIwNtuRHGj6A3tBeTOhQXxXeoEOD+q+
tFqFlwbxw4Qzh3Y70QZWC5pXIuHC/uTbYpGF5ejwWtrtyqr2/GYhxNOjn4okJ1Vf
EbLy/bKnoGjeXRpfB+SLUK3DY9VTTpk30U0X70653H/vlGaDsKLkSs7aQQL9x7d5
fwKEBNlj4+Bsgh+SxmPgYJ/r6svqczLWMU4hxvZ6QII+EiLFCAAH2ts4uUPnquz5
EhJxOf8GaCu9I10LvNVYN7oRALD4ywdxcrBDkv6QYNftbbJadqjtHBKr/W4fnIul
np5oL1hg2p+KgpgGLqBAr7Kaj9wor5RlM3BeWN0bt/usUHTseGLwa7PQzYvWUo00
lhm93UqYjBU2Z4QBmq6VmV4AkuuuieJat5hELYSkpruITns0qfcYidaxtFnSCViz
G4bWWVwjT58i+EI3YAp/zqqGwyx7OvGbpsPSwXTlfSmy2VyejgAXEsWCAORqjkhX
/E7etqnB34QgCVgdCzz71eaLkUPQeqRUZ3jST72ZRcXHgOY2I44iXqZ0x0Suue76
TgrMmVRth0nv5Uzg/neuLvxH23uv3molUf3MhkfXBvSdXzNLyzEpA1gd/Y8T3XCz
dF3IgCJNjiQ1aBk9A4dasvYWt5UK/E6TD0ediUono3G1cSjz6kIANsbZfd8OpDor
B94IdYqWLq1MF/JLu8P+UY1Aum7+LiZioMcaIAkbo6ojUzPqxJ4uJZ0Ydo28qaYJ
RWj4TJSojbPW4jzNw6LGGZL4RRxNYoOoIKitGwB6YdPmH7F2iM5oR6Dc0nSj+53K
V9Vp9wWwFdT3r6YtO69WBSi6Oa97O7QyFDYpWVT7vSy6OC27i52ncNWgtF0DVcBk
NWpEcnKz21TuF1HoG96R4Y/WpzNUZYHAgiRm7NYCFssfIPoWwEdJXLGH6R+Qd3Uc
0qnZ1N1bUoIgUjwMiuSJvc3380WiFKkFlmP5uBpldOlYEFZtOkHMleRBXRiBip8a
4nIzJ9pMPT2csuTL6lYxG0QA/6tunBNYwKp5Gx36K5pP7lYKGvKlpQInIB8eoKZg
4ZDq6mnBDaU6A++sJlzBPI3nAivRGV58nQVxGrlr4/E1gz51HrUVVoHfqEWd2Ufg
iKkhIy1vm6UsQw8w+gYbEf+jSYxGmNKizITUIdikqyYjgcb4XXBWnYkz3b9o8O32
B6/kNvGNquhTAwOaLHyeS/zox3V47GEU7gvbHfm2YdlxY8/oYiePHFjjQxJM3Htn
vaw5Sez1c8vPjdbT9t8Gujhq6cF9L73iRqEgsU+FFgB1Igb2pP2DCU99yYPdW7Zs
o87mGpvKHkj8WJ2KfJ0uMUplTe6A5gVBUnMItvANpkirkXOBZf7w/zv+KIsV3T9S
PrSVfqjy3etdXgDX/68F+x2BauXi5oyPsUrwRmPmntOvZh3X7JvHGmfcGQLSl67W
/WuuQH71+YlCxDjB+eUubyV4BEq9JRM/IRp46tBEH/aEHLvKtUx2vJYY9zgVetKl
i6nQLIGQAWF9nmUuiISZ8tOTZZOD76H6FhCdhtfXbWyI1/qDIX3sZ2SWnJlp8Q5b
VLzYPTOzUmon6zJ3Vq3uU93rJesZ4np3WwFuLh3cP2D72uFRNDDQN4OVkTFFwaI+
W7DzepYuzk5GPGvQIDTbXfzMcKeoWaPQr6uu0eoG+KsrhUOKwj++ZOS2Xw7jbGLD
TyQNlqEaGMhS0x48qqHwWO4jBx/jJlr6D6BrgsgixbPlHh3CkQOCfUnDEehxw/Sq
mBnL0EV/P1kq139LDx7BQltTCogXJUnL93cPzoKTtXrIQADFtRkg+KKwyEpQ1Bl9
SmawhTdwNZGYpGuWpJgqMm2I70CjpwkCFemtfeveLoGjmtBzwE44h+fd2Jm//aO7
tWSqGyR8SaXA/h7pxeCoyu0KKr8yEfcPIo5YKS21t/MQW/o4im0CZiaO/ZUaXIOL
3Yu06EELz3Qq41MM2dnjZDS+N47NHLwe9XuRNVZTwmYaIL0jTUXmHOS+c65qXXxg
/8kCLDH+jtB0eEgDWc7gbsFdJVNEK8i64jFWh6TFcCaueES6MZKM57lRbLCx7pYS
cR7KxPWnd611dt9IyfLabNEWrNIi8ZLUlDBHi0gNwzFZBpFEI3H0xwv5GQInxLW3
C+GyzcXpakebSkDwLay4MwAVkDjPffoplFZxIiUq1bgZfQh4anuO9IWEIO+0rRGx
vOnUtD4p9y9bDoKCCk6MC6DOdRn9X0xd7iHCUFq4/MITmE74qL4BIVsRqvIS/THF
8G0QDKKw18ofWJwsY3deNBb6ONCvvHB4moN1SB0diZinVFEwHTjTNMkiy3kEyV12
2l0gvFLAm44YwRe6O/Ls/AxAx25KLwveSgoJ/39VnLqw0Y0bjlKwzzjnU6MKcBTc
t+eMsRl61wPFT/i8Ii9QN7FEHgGw/NOCPDI0P4PiBCFpY1O4Fuejnu6DQ1GWhS2h
GpyGXIDdFlCQHMq/4NnxrVzda42Rcge+/dP2ZrusxkQBFo/rqDhKP6E1H5OGtFzg
Z5V8pv+8GnCBOpwlJE0zvJcLfo2rX0Krg0f63M8R94p+JaJVRWmecUfpSm3qxaW7
Uvuiufk8gkKu72ktcnHzx8LG7KYtbOhEKuMeUUmRHHebwZbNB+eDzFRVg66xxiZQ
CCKs0AlI/rl0d/OVK07StWGWFbnFwtEj1kNyBbXTVvGjSnEJ2lYWXuvF6srIiOUz
W6qf+ZxXIrR/dNUh1UOxONKE/kH90JszzBAObvmPqx7jLELu/roZK/nK05AANhb9
VrItdvkjcHEbmucHhYUr7Eil7CrvoX6EhibsY952lInVlakEpTF1Vu8iU0tzaW/O
EPdRJ6xgkJTCJZw2K6xv58BgDWJ55pYRbjio/LT7s3ETLmhek277gGBGs2jN5FtB
B/ivDPknne9NZ3AuMdRAjXZk7VwDmvjp8VsRuvNrXK+Db52bda94K3mc7GPqvZZE
uiujGBDzrx8Ge330S2gPei55d1/iTZ2RaqPYQOuWarcZWf8SquJEGsOGDIcWgDOV
h39kYdiLII4b++M/2g2d3QUU6WfNXIgf+4qR61Fx+ElwCH6Z8xFyZedS+eRhCRdh
1aJ7pP8z7GyU+zzWfUHBuwhVLNDlAz8OyU0lv3ZIEB8MEHN8uc7q7+CUrz4i8tWs
+7NXrsxsDU0sZjlT7fZd+LRQgkTONHcWsH4B4MA90ZL/LOAVLrs5wzbkRlG/cztC
PXwYyAR17TwYwHloqfkDRbngqgOXtv6nREhoWrGEJ1r7WS6bTey0EdD5AzkZK9Ql
+Oz04btvW1C4Vp0ymZA9/Z2y/IZwztQzDLTAWPpOju9uRppkM9oY1g44IXAKHL2P
eDVmLhYDAG5RBml4lDwlrEiVHHRPTgfzsIk9NdMvEcWzezpSzl//skC3As1zqn14
DFywTtD3gVOKHwb7dkeGszJNTOUl/ghagbUnzlOzwB8HzJQlrDR6PJ1VT/Kw+u5o
aexpRz/LqJHzPFEKQYwQhn+umDZ4mJZ2CQv/iG0CwdFsDcbAIUPbE6xlpd1GhleK
AvtA5ToebrL+apx57xHRjJnb0oLpQk/NmAPZMlICTdAJDWy5pOXtxMpXKjQbGLni
6n104TPq3v/Dnb6YVTef+2sveVUf0EqYPmBt6GiFlRPbW+kMFkg+80dvlWC6fKHy
rv3AY6I1HbANDOT2mw3tOodZbcUEn6hNe5aZz8TbpR9wCqJjMTt/Lgn/nSHnZfsK
EaqcFeDgqzlantMyzHdx/A4hdIS0YTOTn8C0+WKe5xWlPgQ5MR9CfBFTX0y4jyCO
dXZ1k/gDWoSPXwhIYOiWcKFHp3M5j/hPjtO7vL/SUlN+DMjNSl7+NqZ/wnpjltND
VhUsqHCITUvTPNxvVVZfF2tazghguuVT10DAbzMbYqrYZdHE6HpXy82mjGfaXClx
kxidSkjZSt+IKBwvnDQByZC5aJ999qOCmk2CGhXkweiKo4BiZuo0GzEOIl/CDTqh
i+sgeQAASzAoA4TU7Z88tA8NlmTepyWF/23rKLR3mTeWGan/k3Hu8jFgoSyI8vK2
sagLR2YKyapx/BZEjMaxHQ71Za4KNQUSrysnHsIY8SCGabpI5bBgxfIE1xw/Ygmd
IEn/Pz2MRwYQduv2J1WLP2j1aYCNVYYQq49fk0aZLXEjakObQsk2jWUZRd+z8prk
XmJfU6Ox+qmmDh8v+uZWTx9yB4vJVk0qwCYyoceucEojG/e3jrUDFqYn7x4S9tLD
FpCvc0m92KMtY5y6AKYe5CF6KMkknI0U2Xt449yh4CpC2DD74OiRUl4WpYkGKFbU
FAtnLNR3mWJttcgxngp8blr2xF+ZwB78YPcox4kMGezRO+DoW7oV/D+5J6Fx31Np
H7JXPnp+HnLy+z74mCQ6nD4HMw2upHVJ58KWE4lJpFAanLtF7mEas1sxYRT5kJ1E
upvrImFSG8MMSKbNA29NF0OqjjZFd1kXC8dtUa25+hI7M52/MWwcbwEOzc4nhpJx
EiTcpq0MU1xhbXXv12r8JM2ziPGrEZ4uHFrINhSWtu2S0kjK2+os3MQhNVHUOlcg
y69B7Bvtex0svnDnCWdtuahtLDcxpxxs5SkkzTOIgbbZ1VxL99uc5lyL2mkHI4ls
6o24lgzISmiaOxw94aij5G+dz0OSd6nFsE8UCrXiayHTFQ3WLYPub2sfB9l737Jb
iNvIKu3abyr++BFe6mFq9uVmi27mqrUbP+lDbPGybXnlb2e9wum+Ux3V4lUhu3LD
2s0xmaS9iIgG9eUkMrXwthqvXpPZN7PBqM2U0NJmh05Ue2OGZz5d8Bk608B4HzvG
54UEABWfy/vQqBJEJKhxH9RftWWjET1qqqDkOXc6tOhbva7apxnooD3lkZsqHNZM
Rx7T0MrF//8BFE/KdcX04/sNZ4p5GphHmim2kHAUQT1aTz39sPPshg4fpUY7bjFR
5dI20KJGtfqe6CTNkoLXX3PT3PJ23S+lNXXInoJgAcFFzSES6RUOldUt96hUmU+O
ERkiZy69nL7hpnZQQ2s7e9qCw8Fkt8IlBwQPD0oUB3Kb2pJWjArw3DzbeJLNUE5U
3RV0oUjs/XPuFVejTmX6bboAArwlV5IKYprGLZzIbhArMqeT478E+iZ+gia3iVwR
zi1C0624XcZmsBmGuiOrXRwk9HkDaAlFu20r3jXZpG7YoaTsq6m0Lu0J/tQDuyYe
6+QPt35S6ZzV8YdHiaqFBLaunAAONp10bjjvlxEQgkdoxSFzGAWdhZuW4Ujgmf4+
RjPdRg16I+dMcIPH3fz7zzAWpkrgIa+GA5MflCKRh4w+AMguGHwYlkOtviGsNLrQ
308a8v7xRBeTdto3LHUD+C2y0UhHt1RodJG2aDCqug61qKM0EJ8eLNYXnYLI5gCJ
y59kAwnB5opxB0Xfgb+NGhb1LVE5W1rWAuYDBjxFs9PK+mmTGJqnx5BCzc0zD/4D
vRB8XxeTdd+WFTwPMvzhE9dddwv5n158P0HjnP1LmRfCDft6No1/l2Pm4vMw09ld
3NNv1ukpgTeoQUiZyFZLV3PY6fsWBKQgQK605uwZkhFNZPVC6qhehPKFrbBpJfB8
1uNLkwFhGNp9HvhIi5wqTF1nDJ0wrW3UzPOxjuhaANKznnMpm5XJZY2BxLuR5JMY
ZkrFbkbyEixlW6I9KZcuT26NlD1X0KMG31wN7tVfZ7OMD0ejMgL9S6XR5SQqZj4u
LBvNg3ociWFgmHxCEtf8UN0zJmBcXC2hrp4WlEeIna4EZNQCU2qmlFSDbjMbzXW1
AGdPceGwb57ZySTA/tE05lHkn6ZJER0pgzax5YTq8m5RWFL9whJ3LWZTBqk+T1mI
vVepJY8DDHLL+6NV1N0wMoVh1bvvp7hJnKqwLyerIK82tygvwInpmJ/+ScoG4+B3
twN+PG5v867FqTOuKruPVwy//fExyMH+M9W7InCZTsaylhhB5UM0qiN5DD0a0Khn
H9uWOHG5esJaQoahH+qkjIkaaqp64irXOocJuo/Cdoj/hZ976VwoPDrW4lL3mfpj
favv5o+8IbNY7feqbCqrFLa2sJlTTV1nfl96CAffeiRom5HpM1SbBUe1qGuy/yVJ
aSEMdHT7m0f0xas/65miDxExWYF6XP09csM2yTjvTz1UsXrewcFVBZWVZzZTmBRx
QvSSZAouxDFYj20WkaoQvKjGyAtHu8kdeGaASxzkM6YM8gGvVop1lXzheBBqP6xy
DAVXkM2gZcOuOI/zz00vaiguRb4Hfrol3z7fy0X0kyUYs9nwsvMBuXE8jtjEFAke
q9KcRtBvC5uPwBaP4NyWipK2ePE9lEsgA5lLCP3pPy7IN74H7gcxBvtbiNG4N61p
HIPUDtb6TQ0hVOml7AjcfVHe9DCeCwYsAOndR2b7Tf5I2nvCpSnYVSkp8eBcznzR
ZPgf8fDHXTRIbyNGiaeHxo1vYe2Sa70h5QtZATLOmo7zb826xl+fxR10twLJ635t
E6nfHKwKwx6M1+iElJhs6nIXwcRF/C+jSMYgR59j5/nX596ZcjvGFJcScFqmUx/K
Q0AY2yTBJuVpu9o2MPHYMQc48toZ4oRY6UoWo8fUdlWU6JoGTUYVFRxP4R4j0gvx
kYYxo60qVvHbpRn2CF0FfjpBGUkxwT68GgsJriaEcjE3vl0IbCv6nAcQQLkGX2Hk
PQme23EQSBMv1rtOnm+bZ1Vn1vPmjsVFbpm8dBazensnIzwUyU/9kPWPDtO02o7Y
lTKQK0F5qRqrBZ3QGlQFSIJGmf+QR2ClamGkIHVIKMfzbFsM94381nV1klbS8I2e
Nu8FPRY/7X7FKI8+jWyJaGDlwF9kozkd7+ZCHotzM95YZskcNLp+nuZfxpNiJZ5w
flco45PDI0TlKKoWeZS3qX+W7u2WyKqM1/PncWMeHhFsNcZdjHDZJP+ZHQ+wPl5C
RjVtAIvza94V1OEQGxqHROyOh0b7WkVhRdAV9VBzi8AgBHZEBZlQc+K7uCtKHW+k
DXTauLCqNLdVqapeZi6pv6POi4QJxRDXm9DqHZ3yXnbr53FMNYMpC5hJ8Sou5DhI
+bC+QsabFjPh8VSU6ZP2DWhuz9xNziQksGZkkBMqoJ+hVrDrnOGKuMj3bGAoQLH2
a9Ww2BmRX/VM/7ZlSWQFwrMhy8C7SYQFBBarkbS+R/QFYOD36JtMzVHUKA58gDXC
ryjif/SlH7aQYQIZHTytF3u+HRPyNr2fhUceaay0Ec+eI0cd9eVHEXXS3iBRssru
3fyVy/h1/siP+FTXrSUdbaxA7Wtm1xr8D7uEom+08mKQ+AKapg5UC7B928ZwBT/x
58bgUM55LATvOsC2d2rubURe2nK8WsJi2sy+N/z+i/+UDd+DSbPux3+4/r2MDqPa
Y8JLtEXCBSILYlvVNgga+qqpp69HNSjOO9qp6i5dYT2l//K4wvV0j9NtpvtQ03yh
65rMIN8azERIb3A5tv41dLx3HByuGB4szsWb//3Dx2V5ZpygwuRqqZ+Rpb/6U9qh
Je08aF4Cj+MdQQwBO6dk0c51+0Reg8Tbgljc373yoQMca7Sm/j3e0uofURBGBoVL
IwLhOPXf007ypgu6EgUsMgN+34e+6spr9F0kqp+h/jP3N+BflXSXXqADMel/+yEb
mmEXgrj4lOwC4j+jtQ7wuIDqGtSjHEtM6Td7gFCCXR3oar1lJERNjRIlX4EmPPC0
r7dJ9pPZCJB2nUGhMp2LFWDH1G2hi3kDABeF05QU9U6apkXJPuo1Qqw/dsP1WyxF
nUt9BYqsICHHmUORtSGY8rFjUgu/A9OKUDeomioYuK1dX4TpghJqnqk5JGZA6DCm
HzlCXH3hcmk56iXg8/J7kArllWC9PnfGvvv40v1rXF13p3WWXYJI6/BvIp34iKtC
hSD0B4YWOtYfeZDLHbS6IfxA17OrT0XlttebZd9jwVtIm9rghpDbfviIaJn3SLcK
GbDmKFoJ6N+uTFjuslEFd6tiRzitO8DY4cQDNtoGHiInPHwTSsb02hQpmqr8TreU
OjT1GQc6O8YyHfrDmFV6ss+P2Fk8kSpQIoYx9jUxA+C0ojOxbOoyupNqp3DhHm2Q
4V3Ze24GoqG9inmGhGn0VUm//fTj2XtkNbmO+Ft7IvMvSrfuOPU+kR1e7YkNJE69
MOWjGKAhHjepyG04kV4ltyKc6AmsulXrr/+gmdv6SGGCq61JZrEF4ckdEQfv7Jh6
8m2JamZfXAuk9WGMUblw13tMbrF22W1Ise29IJnERwIn9CMb8xj4HYuB0f0LSiCU
KBjT0oDr5ahY2X6t1sng6c8fzKSqKaSWNcG0ckB6R2W6yE8yY1aTt27GUK9UNCNR
FXP7U+W8ge98YABFH5MN0MJkRemK1LKA+NLHpvTQipVv9YQlQlJV4ixMunU6SfEC
CP0bbHjS/PYefYrB0sGj2UXwkk0SzV5Er9/qf4GT7VBWEMDS2SA88yP5h7+33b6S
k6FvVvH7oJJctzESVA/nIePKwY6Fg90TV35JGLnmxACbM+/vcwTA/3kG9K+sh40S
54OK4wGJ2OQGMkkWeVJAD73qXfQaAlMiyxQdbkvykz/3p9wygPOifzI4yv94o9aB
VF8cWvACUJB9Tya7tmbWgXU+Kod2qdsXaRiuUo+DjI13jkJGPV6SdeyLT/CNwHij
QVj6FlM/Aln4dIeKMzyCVnLidO3UmxyZ1pVf74VZeSTK1utXT40DUrruLHYhpMb3
CGPrrcVut82ndH+Jx9dtINU3CGvZxRibTMd+JeQXdrAnpMI4h6DIS4XaCqWmxosn
Q0EJaimBxvuVg8qUKpsZwmJKfI4LzrNw4emiwnTc0vYlJVt4SFrBPi9wZeM5AeDG
fgV1Jimu0ZYSUQ0MHylN3o7nFa+zHoV5xiFVwU2DgFpTopv+Ww+GGPqRWCA/J2Ri
ey0pROE4cLwoHqd/dxs8nF0/dHRL/AxHxfvcdfZSJhRDQrAiI7PAk6NsuqriX0p9
WfPTYxtcHtZlYno5tHXpUIOb2xqK64ZX0zjuO1QDt7LR9RnSezTFUGwe3iLnJ91j
vjcqsKRCOZaOoOu8OhgInO9odl+kXV7uCSc8SFroY+VJ+DtidL2koN1lWWmmF4VT
HIpDURvvI6sS/EOyq/zFHoY/niUnRFcxv2NvKTF3a94GTGjXhkVPIOs9GcpgTVdE
S/CKwqkw1itxqBVMGqeu4gnHrJSxm5O0G14XGTdFabB36zSrkZP8B+BmeVCjOOTu
tJX/q0Y5i0YEcB9XnRHgc6TgKq04XHTFgYsPwDlN8lhFOqy9Z2s1wJHjH8epj4Ly
2crW/cjfiD4V1dCb0eIE8CjN5/wfYySapJb/o9EkrB3h4lWx3zoLu/2YEBnV3uvH
YUnPEp7CZFOixCNf1LToKQP/b2Jo7/cYIQ3HW9x11K/ddEYQEZawMiZlR9lL5Gzj
mD+3DRHNlO4Mw2hcpl8fsecmcY9URBI4/pvLxzclanFOidI0nu2T3txEnPcAm57E
WLqcde5bE1QWfO/DxuPwsMG8ZJZYxu4W5J2BXpNxecFoPtSTEC86Qh4xPXZh9qO3
sJdFadAnu+1W3K8RhUsxzk7U5PZAsP6KvsnFip1dr5ZwQ+7jZ5vXQDBZoHJNu8rR
xjzRCI5vcltJnnJdcF0ErQfluKuJhyFg7KpG+1kM8DxP9jaT1lZ2oHmVeMn8kbbc
3lFBBRUqCGTUm+lseMqdQbgTIWWwhmLHvHf7XDCwelogULm9EjkkYNHSI4ISnt2K
kgNuf/3lK0VlDn7JUHmhVrwS2fqX3VaL2soTcU4fJmAZxZ4CoRix153aVsGSFJMe
uxlbJy3gDCFKIpbO2euHssJq2d54fV5Nu4RW6KHka4I1moQND1lq10a+4IQeo28y
DXUGahjIq3t7vEC8aPYv5lzkcrvuwehyOqJzxS2MYeXwpVfugxm92aPaBrQLs0fZ
g/A++i/BjsB47dlcntOxuUtYqiIAJRUW/NebfPmXS3zpwdmHE7tOZ6VOQKfOqVG8
GHqdSMnUoMkSbOWxwbC36+mAlYTqraDIepRrw6Ry95OoIS//p/734r3zuaYTNwte
t1ZWKXB2xbQX7ThVUcP7LKVcuJPPj8fi6iNuiAmV+NQIGE3bKuEROfwC8/Gcnlfe
VHa/JD2n5n5tSmP122g4GaeRLzuc2TbaQb8ozZYT6RMpjvliDWCKeejXf19KvOdf
PZbywKEB5PI72bEwz4kh6WhL9Zrfihn8/wQLC9K/b4+zhrjqCKU2np0v4loO5OeQ
tzrej71cLbPjo7GjPqXLp9SJeaTRhelO5wpqyWDPBxeO3iShTN6ftabdZgqwyKiQ
3vuRzRNTc8GvVuEK7TxBYZqL1Ied5M+ERcxhBw+NIu8ZJ51OGQysPVCjhK0820Ri
FJnGuos2Zw9BSTJzFBqY911v2f8GTi8XlRYMnFsBSm3LJXSH1WH9N3gdDJZEjuv/
XrWUywJ2g/VDDQViP9IAan+1vZCmUa0OSnRrOr10f1rV456CEka5oqTLJuDct8tH
zB7FesNk9V/xEuQvhRlYbqTB6TR/tPOUTztRWSe/ar5x9s6xfCMSW1Enwq/JIj6x
OWDe/gYJvlhWdeUypPNyB+C4MfgzGIfebj4m9vOOGghw2O0E/myAHAI/cvrDTW/h
NVhZQZHBn/c8izNAvZceTp6s6klCdXmv5pYus9rUzsXfOYmHRQmwMvZmFoPOt1PB
C4kQvIButfqjnU8ZPJc46yFatfmwUH7+7ce8r7J49mUQmxdxOAnoJzEKqvgBJvbK
EBiSPFtLe1g2urNwbj4AWw7c7ggXjOb4xl4N2rj3AkZ9ZS83cH7nzViizLP90J0m
45K9/vbOhZZjfJR2fRFM+lRV0MJ7FyTRMkfcDfiVojXwOKIU+dq1tXDkdJJn7V9h
mWuUMT2wNkeNHyaqfh9fom+NchCm3j4zrB5sQTfLXHAK/ptV9O2QfPAB46JSHagC
QaRQ63f/qa+12BSKzov9t5nrnSvLWYRopeuwGoBdnN/BshV8A+zNdvvAAfFsYDv8
c37rS9CBFJbgttBIw6L/D/AIJN/4xLOSqBhBHuWglr5ipPYmfXLCLMzsbxwL66TG
c4OShWHB1Zi5Qecp242OLsJc9hGLWAK7JLNWoSnGroGqKS4TeVIL4VH+Ze6M48LJ
kvRfM0OLIQyEj6f9kwvKwwWxQjARMwdl9GJm00+2bk+nV7K6i5yBxASbytS/vxTJ
uAaEqyZkPqGHqxvfmzg1Ken7Nyi42fBzlpxSvJkkv4/WoClopbfngphtxwZtyHPp
BJZb+w1RaqPGPx3zsv+x9CD7N88IAOlOnUgz6CKJs9dV9wDG5Wieue6BXx5+onzK
gPTinDKmM9dpzJ1WtoMwTQs67C/7L+cLAg95U58j/WLN4aZ2dZa1/Z9GipYP8BRX
8lmWtHsykZbBkBD7WJrvWB/ZL+3/y12q1Jso3erPYVJbbHD30P0W9ayHi1lqNs8y
u5UGe282mg8O4fXzW+4pz+MWIBrQW1dahZJz9mibfUVYWS6MqHxiIeXRfGbtGG3c
a4EXffgBtiICHEIjO5P3yOpNTmbZxSxUEBHtHw1PrSOXC6oBi+F9A5fRDbcneRE5
cfjOqOVo9NrXdI04oI8eLWW8nCWmgND+jnqDQNs9NZblodMHijVomW4ZxI62YgIf
sB4dSa1pHyvQafK3xk9bGXJwPYKAm4BsDUAWqWW872P3CTKbEkVKW+mKo5+I5uke
xX9ASVv+kYBRV9dcWNJOONQ7ixZiRd5ntzYNxksxMmD33B8Qxy9S66g4y8PUaQV1
WbLSsx5VrE6RevQBqyS97dIxpy4tS8LQJZp2BgtMz3ZzfuOdwRnQCeHhgvP/P6rE
5ldIr1qW9/ztpYA+LeCYLzQ+cqmNEoHJImxY0ozdlmvHg6pkNYwke7JDWCXOJiqG
J6pp7gfb33UC71uuMRgDMwOIflUXKpONfD+WnBo4L3Nd2Hr3V9Q3U1Heskbg6Rpc
uZha25SHUdf708p/w2wKKFzpaTi7c/toEUieZu1fa6/C3bvieWgohWO/Z7+9goCZ
olkhPCie+0+a0jEbxHnXDAtqu24Cr+Pzt7mivgaG/aiM2HaqAM+5zPD+2F8ohwx3
wNy0PsCJGDMPAUrG2hO0Az6i9t5slIHvf52Tc3lFLefcroYOX/YqTYX7h5u2qG8K
uviSt6XrJ/b9ZwiGPjCBVLD+UIYyvvZjlMEd61kiLFuO80PZl9Cj3mWzYVsVmHeO
pdj93RePiirZ7E0yI4CWKbdAkHD7kd8JvuEIwbhebatkQ7rlNbSTdQbaPq9gwvFs
PoH4peneyRGCEqXfLnP+DSmf0QolSw65nt3KYlrcsCdY/x1ZE/xe5hm0Lc7LUAoh
KRF+1rmhCUu7HERzwmHsR0a7h7BlU9OrN44/8VIpRLdq6tP5AArnG4nOmhFkRGVc
SOUlUe4iBed25WAEzbU1MlnRIGpoJP/Kxnzzhj0WQ1z/ffbicTfA5vGJYmW0MBtU
q9LJmWlLsqtyzMPwZqRMVB4gEikgwOppWt4tbkbNk8XGD+W2WyPgZ1HadCWa4UFS
lQx0ivjJ8ss3dHDPrtrnqAqXdrrsQ9GP+ErZiVoyEu1H4a7xLL3n70qjraJRGjir
zfr1+qJknJ4VOTY1vK8P9oDTdZzWcttidJvaXAzJRXU4xhuJ4zxXKfHnFxuNV/T0
uKvZdHsX8Wlj40rWHbfDZ06SuldtWJN6XUMCbc1OpcwHKwopdUGPeSG5wZkCoZ5c
Hz/yk1RGnoRKXQ2Ohg4R11AmVHlTCjk7mVzdAHFq0n8ck3OoGRIX3NIRva89l/Xw
s/rAxuKyEToNmD3AQuTPsbXJfNDQdw7HMGhu07lMU4SV5VP9UY+y9LjGR8K3EeXi
GvOmhobpRE7gsZARvc3Wer5Mx7UwszexJDYwNtqpkJ+o7mlruWKEHG1boFdWDdGR
bKHG0w1I6D5zwjm/sXV2rGy9ixniaRDuCB2TYAvian0Nn4VTNWSBOeOv0idXffoK
vd9wmzo6vzy2ZNRhJRaHSf2kjkujNrZdCLqGWiyQrCQVYCEUP6OedErJ1pn0LBMR
+LCwXEiFwJq5ajdGfPccVCc6+o+4IEVwpj+azModd+EDa3fa+m2OoAzjhxuS30Rs
Y5MwOnxN64aBy4TzY/nqo+7CNbgq2oeCEI10HiX+aDcfQZInGHqwps4N16Ugt74E
YMbIljE6Vq7UREuJcPu8BfIXLNyMX4vQCCeyqaoOAHBEFqkKSWe1cNVnQ/Efdh0r
mezmASrQeF3thD85JJ4BUPO2RFGRyAWEGrfyUb25wdq3GH2GJLZYsenpexQJVa74
As/avBE8wwx88yWWixbze2/0VlluTbDOafKWbr1pwpjWIO5BBUTRKVMB4IaOhqT2
rPIlE7ptNvaKxHflV3Z0jZOFmOVwR8vD170QVoC97TWW+5qijpmm5KVsljS83gF7
2HSfJoDyeMg2W+Y8WBYis3i3kn2AtbWQD+8GjqRh0GXynOiXHJYV2XkVZB4I6Z3w
sS45d5DCMaNWbNSwRdLEQYLXhbg0txS/jIS3Ui41ntNSJGJtp546yZDM/4Q2F03u
gXe/YaHcZTSxANo+IyPGCFy9VDV62rmKr43EqQekdlz4GkayZhHmliy2W+b6mOdh
VtsVWaRxNxsaqD7A8Lwvk14qjYFbNZxzMitSbTa9jwSjwIlX6Ed33wZsYwEF95B5
VxvQpYRbuTxFNoZFNEmVJXO0Amthya9Z6ziMiLINNbR1xi2smx/Gclkl6fmc5fVn
DVHEuFeSRJ51JX8qivrlMd4DdP2Xzru++aFZ7sBgiXgjwhVT2UHxSHF18IjmRST/
oEonf0Q8oZqXszvmvtR2SLGF8x2bq5hwlvSeK9PREqLz7RlZAkbEKnNmUc9yzRFD
9nvcmMqa4H42cN8O9BFVeKnVbaOMqv0o+5XO2OL+mGPY4jLzesCZjrDv3OGV3Szv
CoxiIQlXsjQ1EE6ZgySOr30AZSpIkVd0QpKH1z5C/36lpKe/ReyAM0D5W8kqGgFf
7vD7ygHJ1CM1A4FmV90PmDX8FhB8pXlo9FHIgm2iWfPl5myixf6u6RCyLEitKzCr
FJGXPzrQUWfPfbGKodUZxfNsuKvawVy3pXqKE5xIgIu6Vyfba9Ql2U6KzSXf0dj2
EgIqzkKvDIthxIBEME8i8i+9yP/0hEna7htF55edf+N/GZsfdjHLWsCKaqbwa1+3
BZAPgW5OC1iddlXiQzaT8GTZCn1XIBw5yPYhVIbnnhV/Fp5FQKcVnXHImHTWRCYd
hgkkChe67Z4I+4Oka8OI/ysoqtBJmNNyDLqCfcnFeIQMFrljC2nc7j8YBGVeUrwb
WLz0rFQvaluoLisvqOcNcij8v3pnQ7B6nOm7Xtt9a6pWs79QFlJ3OhaxdNVT01g+
/hrUuG006lzBuyssoPfCBpwqWuVTmH/S/INU29ixbfkmeWSkc4LOwK/1wuq8PxD4
029nTZIf/k2Oz07Yk9NagePH3KbUNuNXV5RHW63+rXqYJm9hoavci8WPy+1yhnum
Pzia+JI4bPiiEy0CVRI2swfqjTEMukytkw1MUHhGNbVavnlPbOd6AXMcPX/mBOjZ
NZaYyrA5BVzKrqUjQbXfMJkRgfirrlQYLKRKSJDpbTWabzrA7lCHw+uRBeWPAHcb
oH16j5dmbHBk4k7PCcgmhCVDjQA5r+rH6kIOzCElQOkYK6lj+n+3C4qDSwkptRPG
FM9AwT9rtrhun8xSRuAFnIL9ZhEYtF7HGtmdHIf/taAPltX9hUZ8lX82jl2YLfc4
Cp1nSJM90Eo1mS6ALs/bciEs4DtKZqYIcTF7HACi0OZKTliZkeNHWxIMlAOYtyeO
0ngKcvIVFnqhuqBADc1Gr+rdj+s8NJRSw9OQEe5gmvEUEFeB46+wsWbJ9Lma84Ww
h0uJZqc9TZg4+Eo1m87F99BDASSh8MRT7z2+fN4wT9ACIrPPMjnFJ+ZqWX9fj0MN
LPulgsEeglB6jxJi5Qsya6G4FEg5a6zO0Ky/3YDh5jxUOwR9qcXBp8D/MBiRKDBW
+wHiOsXFBossKQ1dE+8Dl7JTZP6x3GePxHU1djnwKmY0htxwgIDe7zpOov5VirAB
tKx1CDZxwsa1lecwAYejey/YjNBUyKEBVzvoAnJVo+yDA/4OPrn3laxFvUK60PFL
gbP+2i8p2XnLeUu9zIsc0n+MNh3SDY42DJzlqv6gWS6PqPKSsSa11wz/7bU19FUs
DfgL/iB88kgRQUGiYS9OqMgYobH1VbplXw1sk4JLFNDpM2hTyjWraYIGMic4zfO4
ufiqGOS8iofK0zYLI+BOCQio5gmPtUvfLYD6SVe38SuUJcZTAXIxb9JdWuCsgrTQ
8VJy3PVTJK7H5XYWLEfnjPPWIiyQN5Cn3dhO9LhSwadD8aaoN/3OsLP0us/gvl4l
XVOHdOmAPKQMhIK7jFJgjx4h67O3OW/bgxH2JV3DjVvviBgKDmd6ypCHny6Mpbji
kP0v1JrC38QKo+Jw/wl8TG+fnu0rsFEm7k9uXpW0YkyKozlEt2dyC3k4U0axLWH9
0H5DQ2lLo6pO0oHVbzBO5k4xAztbeHsycZZxnZOvgv6jQJFWqJ1KyL2JvlPyHJRi
1tdw4Bw61bgIB5pjGb1NRtrGnDalay7QXAA7t+I94ac5q2GN24eSkHVb7fD4XxBj
0MtXPePsN6EZdivRGv2SxhEwLrAJ99TLt0gxzD6EZKMA2h1d2r6xZwCoQZmZtRFD
cA1AIl2fH/igIaWDPd7GAWc5Xl2KS2dhLnX/yw+rzTT+FQenWDng4VnLkigkSELR
I2570NJqXBA6v6H93ZfqMDPUpXeDPGAYdJIEIe2S++OSdn7JoHnsLZVayHgEgmvY
l90/JrQ/N6ExJ7TQd+jhKT8vb9I/V7kd8fe4tjAhJ0ta7+QdcnVtL4JuBm99q6Ma
ndsFpjo4JHI4TUoMjrMeLr6AOcg5X+QSIEbGs5JYKyW3TeFeQStLi3qnaZbhdsqt
goFKQ9H29RB8YAB6oCTT+wpqHhgiJ7O8EoVszJq5Lr9GNAIMhqnAtsUnh+treG0k
azS0EQrTzeFdea4GqAKVTZmUP1LrZLDXz+m+AzUODJAn1FKngbRlXv3LBMIALkq8
aKCBVGqoRkk2Hr2cmO2UugY1j46NKL90h9SimoWRtVa8ZTgSvbqVK/Uq+LpyoRnh
TN5IpTscqnwtA/t8U87D87iKr2ifneHY0YcYd33tinyM/qxVG4rC0UHqE9Cria01
pL2QDGuxW3olkNRNWSsxSTsMp2uJmo1pHy7K/e6fouT7nPoSTpVHsgLnYDDKKDEX
ElkU+UPL3CqqQZpn7kWGa2+jYdFBs9L1XtzQT5fhDxlwugpChmo7d3+LdoH3oxXv
Ivgrd5knyvV95AeQGPXYdq2cPaEX/Y9YMTbscGKx931tNmw+/5O7zjtXJ+jI2mry
SbVW6tjHYcn7BGd5GGUl7UUb9ODyMfKfDNp2sYJzvV2R8wD+Vq6QmiBF7S8jkGPM
tAkm59EznlS+NRItSP9B5tO+QX3UWQRDfWQzx28XrYN/+W3AwH2G2u+IAautGVew
GP6i5j5cWquMHKFnwpBYHy9PasbqPCJ/S6qBNPrPQaEFHbroJZvWMecXwHvPqx3u
5Jjho/ou8fq665YOTC4ki4BYZUC6wOdkUa9VGQpbL/uWH76Dv96r8DCUGvoNsqZO
EF0SOvz2xZA23ylgihgAJSaZG57ju2rnxOTMni8ewzQ0yNB2BI1sMC8Ao5Rl3Gzb
O67swamSoVZidKJ2v2OeDjykNkdRO/x5wkTi6zYhr248WJk+3d6ejQLk+vuN9kP4
o1nymKALTMfp38F+y+OCGAqwQc6ij4oGvMaNO0FXsuuOV7uxoBKyGLVhSKkZgGUS
+L5QGXkDlsuDey/mNGFpDwLpM4SJOtufE+lfTvysYPD8SorbDNr0tehkElwquB4r
TQ6BC9Yy9vItwx1Sk5YroN/QW2epJlpQu3HWxZ/sZoPYDWYW3kDXaIfrjlSKm57l
0Ul6dd+UyhoFny+H+Gr+uGdj3+AONKK5V8OBwIgCsrWhYUC/k1eHRy4Ls6YR2ldu
2jcl8t/BN3f9qB0kyy0Ar00ADK7o4rCbMx0w29RGObfMQ44hKacvB/8HvwuiQe51
E4O65WO8VTd18Z7Ai9aaYtGGQG7dGZUy2uYSf4GXLkjjpNzoLvFfjJjaZQtn3S8I
lN1UfbOa0TOm45m8EclhbEnarh2wX1e76bkyHQUjzdnyE6KxtvsGlp92PYlphN8b
wAcvG4eGodiuXzZAhPou1hA5vtIPsfAJfrIfsve+NPnYEc5x4L+6lTt5nrto+lzT
18rEUJh6XYKoohTkzBXDaiO5aqWrZ8JiFPtFJcUchOnz79gnt/yOwCffdV3AavS1
hJUsNszMuIxa2NStad6OSnzAtpG0UMDs1MDw8RqozdSGfE3xwnItk9x9gewCvTlO
LF54CWGBBi7201mctXuKjsZz//U3qEcUN2ByBjg/MhXVTJePsDNw37ZqMedkmnS2
rfbydFpyu37zOysZf3Mz/cFUhP8Z5N3jklGaGbnvvbRlcbnE9p8P5v7M9IDtYk6m
s+4QAojIw4NLbP0ke2fjYp9Pkf1FJloX+E5ksd/InnRjAhsACmpsH4Y1x2ntGHnH
R6T7fvsAAFt3Yz79o2T31o1uXBoj8ZsoNRXgQ8WMXY7Ka4mUzTHx5mBgTTEC4X7w
tFkw3/RMFsSC0piZPSIquWgSOFys1NfHqIW2Zvn1LOK3cavamUlD6IvTz/afcZfG
/SGjIbL6ZeN3+4rr367raPmeXIGQwfbrHv7zJntIODMGlaXySJerDCNUveEo1jGZ
DMOk6BdJ9yoqVlu0xjLcncTnlMA/ucjQlwjI76UasHk2aJZz/inYIZ399POJoUJC
eR++0WQ1qKMrrhvdQ83JN69Xzm/PUPYc1UFH/fU9RGkXz+y/6UudBT9YjBQ/q5Jk
giBIxyRgKtUrj/bv4pRG6ak+gLciuyl8wLetR10JXZ28tzweSYQYQXBqDWaWXIEQ
fGYPrXtU3x2FmpPfVCW+tKh84Dnbjq7k8iVpkEAEl5K4B4bfYi6RaoZgnoBx14bY
1VZObFkGEltiq0KOkPDvmP0ZaEumJ2A8erlXMHXQJWsVALFgjFlzmonaygOUDlXu
XSFK1HYssnkChfAuakCT0iGXa1t0MTzqv+R198i4HUals+Ic68kVIsGi/rIjqjZP
MPCfLMMqLqRQPKnLiHoQVdXKwu0SlSJFXHoECXGrDsatWi+cdDUcaWTkO+hhPFlY
42XPJFr7sqZO/59RHy61wxzJK1NXTLsgehZXOwthlZ6E7oAwCG1UTeFqky1vZrJq
xQExTd/W8V56X/3G6SCcxfbH3BPISQzUdX2XBdJibcBqZjT1bz69KNnum4551Nul
NTbDolVSIu2h43quRmFZTRRdjhH5zNDC5siN36SYn15xiOLPQqdzx5W9qWz22lKb
NKHq5SNpcD7+NjTaET5YlyfZFn+mQHpw5WytsS1ADtf30tv4+m9Lq0WEiE0+8Q5R
9sdmIcIjVDW0CBtk6AvWExeVoQbz00mO5ZcWDoc3Cf+VDUp+qyQNNcxzycjQSi5+
/YQvWgXu2/zz3cT+0JykXbotA6oCaP83/4UDhwoaSWcdXBQZ6927PGojVtoY3Ef4
HvUba27w/RtNg7i7uP/dwhnPA2nfXzH1XAqeoxs7/pV2WCDaUMNtA1VfQtvr+bf7
fNXsUmD/IYOgmZes5oWPNID55aFuoUZfmOZ2FLctam4CSxkV1cUtl+GGQiZ4cCD1
Kx2Oqr3v/51a7m7Eo3qvVbZX7mlC+iijA8ebo2qti4erokxk2cySdiZGcsjy6UOX
NDmCN48EEeGh3NrSGKng3ZwVV3pxPI9y8iB2BEV30C3H+IJDxl1yAkmS/k09UDiY
q9dSEIai64NSYYK46klN18+xPpCnqgzdKEjcS6KsfS3lSefvluuHPb1emT6lK1EY
oQ243sfuIVZqftBMgVgRzq9+NI6IWMin+qgvKdVfjfanq2KRgnHKT4aF5l1UUt4f
F5DEexeVBY6UfijzZ33agJEYCZSvWmhKTa6oeaVW6QXh8lWbXtoKdikw3Q6uSdaO
nNvNmMObUmI60KSU84nsDuIOS6M2HVgb3X1uL8XZ9G9lth4jkcY0MqyU54SzLAk4
IjHrSv7ubLHBxO16TT9+BCCVzCeyx8lof/viUzvowpDVPro3eGpBX8fvPwUW1DMs
B8EXAdnuGlV1T7xxStsTrcRC1urfERxMn+WIQdRuB0vlVV+UmsZnnBvAoGLaU8zU
OLu/0NTp7GkNnN7u5/CyXzmQ3h0nFWsV0VCooe3+YJmyeGxrCf6lgNLeKz+OyP7e
mIYr7tQ0qy8EMPDLADR91EbE56nRoovAcQLpI7iaAsIXapNwESXH/5oJZgDajDK+
5meH/paPYxsLLkzGxu0MEzUo95OHRbHEnwsuJwGLpqyMwAiwzTbVecnV1rakGE1o
x9MuVCjiwrOpkw/P6ZaKz9kOmOML3AHY4nnY57VpIdlafhBNEWRnRXgcQO7Lo0/4
0QddUtvmfiyUb2r8Bpo5p2FvXL2U3pglV015tM30Yr7vad1NKPCkRt3PdqHPq463
E2bv+cv8lcX//In/dqrtqBZwW1KoF73RXo7+RvnH76fgrQdH6PgWh3QsD9aSI3ud
ht9OB16OOBJBJPEEPPMeiqXBtbCys9bskV7CN8EbW0sReZETuI/s03wwWNM/K7an
7HUm09Um+7FMCX6vW1Yot5ppbBGI3uoM3FPANNKDuQfPmSsX20hjMUtfQ+4FeZlw
yGoSkociumVLhoB2e8fuMeV3z7Rvq1hb+xu89ZTQMSiL85NSI9Q1WFJQ2UUK0uCv
tBmHnkr8QOoPxp70nJhLpfbsRDGCZGuB1ZE23KXBALhw9yOlzHCFC2/JAFvmnJIk
niJe8YWvTIn2pezemLFUnTI4ImPcC7xFXCTX4cmK7rHY7YOv3z23RUueavPvjXND
3TbHmyDMXaoCopcXb2Pb7Y0dARCK3pRPknaPXV2v1qHD9Yik1jHaiYg4fN8LF3au
VDKhX49hlRGMMjPD7LokrO/LyzHACgEOWt7CIdkHJJpQIp8ZoIDEg+G8KiyB8aYW
ASyqptVm6NHTKFqmDqnMSUHcBvAq8cJkVdCynHN6Jdsznc66RaxODEQkqMaKzZk0
cgGGGXYBW22LGaWcgeq7rbuUtyl2+SRsajJI+UQ4ATFlKNJO68SBjQs+8Hu1702f
f3cjk7TaDeFhQFYCKhsi0qzUmCGCn2cq7fLbMnE/SYT0H9VM8t+eRvEgrJk6B/NK
SDeH+v7UF8HRKvAnHQdhOVgCY59KUU0txUrCZf2yl64k/suNEjLCvsMOexqgf1ji
AomtXpKNvNLP9dJSztGu9BQxwPcbLSMn+Xqo/iAUVzd6G0wvtX0XqGTp4y9TEqKg
F5hQB0XsZqMt7zsSxxoaaT1l1o7Vtw0JpO772CLYYpYiDfUIivqBcadFv68GRGJx
8ele5tKpauTQFKVqr/P3kfTbupY5dZC2P6UH1kykATb6DnXPrBw/o8aF+y3IgH9Z
D4taB5WiaWsXGdTCo9JqYekIXDXRCwEREUUan6OpmVWiOfGZkivHYNSliwT1Y+T0
FFayUcL+CTQsTpLvn/H4S19vvsS12VOIQbRHmsz1i6eK7QTVMsJoqTMsI6cWjz76
kmee3FpFYftlcBx44IebTRISXbDT1RO3Jhsy9Lg8OzTRjuU2G+ESswh/thqctpLn
t+iYOTszuaiRZOC8jLOpdeH9rOLjMOo+ZC78X4UCDwIdI/E8VCgZppIoX6OHVygW
KcNn5sicPNftOTQINTC0wtBEIpJV54mu6p0RL3pDlkTJcPv2N8F5Su/E73GWh0Cl
SwY9TyaWc0enHFdGuPwT67SWu9ImudWbpeuPApAzma05hLbzp8/HF79lYGAix/iV
UUTYQi4OT9Fd0A637X69QmcjjZ4ii3QRvc7S2E0KM0aEhlFj4AW6qf67LXviCSP3
hp0aKfQIYMgEJ0fNIZ/di0Dl6grJv1K26z2CBm6WmoEQF2h8KzquEGEhpxfuLuf8
Hh1caWWFq2QoMdft5i4ERZF29zKoWgv4F6CeRfApbtcGoH/xE/DU4BhWychQImtl
lHiQH6bMznmmz8WtIoJzWT69IScc7ad1dMORNPIbFpK33fjRKVT5Zks6B/21wPoT
ULdNOhwZ9CnhOSx+i2CCjXUB9O4vqiYzhw+Snp4cuxhs12ZI1YyH911jwGp5CnbC
akCaYGFUYbI1EOEcpe7eZ62IpeL0dfQ+vK6hT20n/MLEBRfWeRC5Y1hG3/s6uWSR
mEkdK1rEUOdNRhVkpValu4EJ7AX3qBGh1jvog++OSsjzrVsZJDIp5eAoPYgXXSuP
q4EH81QGWVQu4O7LemLgjr6rCBjMX+8noNcwI/U70M1YnNCWqPPGdOHTIGGN62N9
w6l+xPP7YRCKqWCKpRMJvsnZuQG6fgHKgYSGuyr+y8suG6LV/u5hq95LD8wcVTcH
jy38KfLaG6DqNXogdkVWLnqHaz+U5qYR3Rs+dzL4A0c3EPszhFGiBav/nKXFXXzj
+Nk1NLElYUtZvq3hUQifSdTzUO2FfmOaDG/tKrHPFv8jACcVzXxx3IHFfeKZI1y1
oFEyxeXCBY1mNJLVGwvuO63zUw09dyBGRvACrQ5s+aJK7hhD0/dQmoWFg58MuwKE
BWZpvqO41joXpmENdKufCIirAg5m89LLlr+gv/YD6aG1CfPNsdtO3f7saLRNUxHu
fY+2a/Jd3e4hgbMlTwxsZprIf4OQ5idLzm9q+0BkNAm6+LFLeJWxBdz26kncjeYQ
ibMS3veJ0hU9g36scubXvsopfuo0gLXYI3CevCb0QwScONv8gzObpvYcxehTfKb/
/IKlkGePGllAcoEVV28uux2Wm1ahK39/qGm/1X2rqQytlJ0F+Kums2A6SYE5WEDq
9i5L3POVqZcgLKvJn3s67C+wutfIn0rdEdOapi6QR6egl1wOJ0vsLHcmTfH236Ju
TMkRfuxaOoHOKXEaQGHqUKNCP/goOrPJlxUtSRSWgvap4Yrvhh09dqrB/GMWEwBp
PtnFtFtxLUYwP0D62UcBQ4TfPQcwZOI1drl4+5WfJQ1XT5UFz0FBdf3ESa+8nFpa
GIosbjhZadyZ8YGqV0bLJ2KmCFiwh6ihpRhrGMiWaMDnraDhYjo1R/19HpA9sc/B
nPjihD+iutCp111Qr0lIDso49bvKpn+Lh7hj+Hsgbxfuis9Ot/uZDAmXuXBJ+DsA
/0op0ncsaeu34tM5DqtQbzMFu+MMm/mybx9oyGJQOpyAqU1MeYTEDXhZgkDEV8oc
QM0d/OYQcyJIbnm8HJZih/kcTZHtbK4piSZ9Sb/VRKUXBEm3Lr+ift/Pu4PI7erd
AiX//xWTOQ3Too8C4qNKNmPDbTj1UI6RJ/hLd9+JVMziLSwAw/k7XhXbiVSyBsqJ
p+WT3BMb/z2SyRJhbobzwwLHEBmtZ99sTQwVMRIB4f5zW5ZTV+/oRCnPEVsOI54Q
8PXeg1qPjXmqSzvXmKCizT7pWmLhNPkWjzdclVGpMcRDatHChSvWixeM2vXzy1C5
/fVPxCEWxjrjNpMgoJxmNN1IfQXkzrJREyRP7/DNbDR1//qh8b9VrLA7qZZsdkbT
M/xzMNFToITdxEZySil+c6uQE24LQvovRXiWyYJzrF/cSUt52eaCckwgY/Gq3oQ7
fEO/aZdFQH4LziLcAVq1MTM1HDW2HYr7j3LSbb5RNWQ=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dY+B8wkvlyHzHAcf50xA7+ZwfwKLisksekLkTUtOcGbqbMekKzSPN3nAtFIE73nq
7qX+MS40ZuYZ7VyYH3FDh9VtJuUOTFToPH10z5HgWNqdLp53mM/oTAv67FZeBSZj
RKQ/963GAhRdaSCFpoCM6liizOoIk59aAzhduvvYnMIAvTe75tI+9msvR1NWum3D
xQuZ5st98A5R8lsDFnbRpiQzr0xtJ5/sP0HEVxEwGwCyZWuPFJPCXoNk+fqo/Riq
wWG4gO9Wniv2WgfPwfLB9eyQBeacaSbavvtxiwLwbLPlfQersSmBgZN1l1fr+xIT
jBp+85a70RlaQTBNTHIxaA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17360 )
`pragma protect data_block
jfit4u2wovGtSRsTZFQJPCi4/fgOwdJObJDAZFW2y1ZahwYOJv8pK3Wk/YNIID5K
miXFq3SUl4xdLcdxduer1P69jtYT7uW/+O/cpx7LqQLJvcKWFHPZd3HG1Yzef2na
cPkqgj+0g56ZwymXRXY8vjYbgEpgElk7vTZ2Ivu8QurXFERq4TdsZhaVZZvZ8gnh
F+zNeCwbbkygTDvnp85/VxiJ+CVNq1e4QckRutGAckdHEWlziF3YsWTl3EDnOVDC
CLwHhEI/OYtZa1o8biECOzB3UEC5rQL3xp/vKmmts8tQBDwwLQjkeIcZ53Q/l0ec
5CW8kAvcFO6Zd21UPiMzuEEyAf2K+ocG5b/eACHZBhb9NtsGjaj4USwKFzBc6hJs
25cVQxSA1euOsk1s2SC6NGJR8VoecVG5oK5GsZhLmgRLnJHyQKXbyhnQrKFg2Rsw
yMGlW3PLSfWESRbz1YRLaaBBDQJNNYMsdX7G1j7ibIWhKaoPKa76/SXKM/EHH8+h
qksCqE4SIIRNXDmBmkTCJTVwjsOvywJbycH/J/hGc8xc6oKWi1eR1NYD4ugQBvTA
SCUe/xnksNSxXypVLwSafzjzIZ0CKrzQq9TUYnzw/IXT9CccbcNjm0Ygb39Kjoms
JKDpdcwBNT9dePqiZTGLSLTmE5vIk+aJJLXCg3G9kP/TeTma4/nt2pHzXwVVVvhU
5ax9wS0auTaT8YY3xY3uLdOHlg0g0gVXca4mShL4tGssM+B9UKtrU6kztcpxsSFU
8hoF1BCmFVK/o1hPXJhXld72bz1lmElRuXI/KuUr6JyK6HBzDUqbYFHRnnz2AnL+
dYGCA33yjzWAf72PNXRkh8FVQAriR7Bf+ymBTYMSYZI0d89Hr6LeyPVRUmvbuo7j
JT39r0lW8uAuJIQ7dk29KLo1Xei6V/xnPGGTEduBPM9vEPqnUS6/VvETz/lfUZrg
cpxBxwzTwufMZB8BLSQ7qGTZZrQWJVGv3Z3PQ9Bv1QZoyAgVHE6MNjnHjU17BoTw
M1hqaSQhtOX8PwR8PLA3AKxDttxdIrlOnHM3SeMx9rIlMA9LK1QHIcuyreIhfPk0
Inoa7mA/VLUVztlLKRoo812jXyDubGerLcFONIIq01g5nG+ZrXzhblNPHxwHiZVT
K8fLk4BviEwkGaITfv3m0VpCqG+ZRpfIuYMT0Ln3ST5uzYlPoJNgzcU7z20trg83
lzNBbdjKf/JIrPx8hjrexOjEC9DzFGC1HpJj1Bxf0LF27j0QG28u0k3tzQGc/xjD
pq7nY/zE50DYaaANZYU8BCMjnWRnNCdoQZIAoOZ2V6aPC4ZwrIMNRvFVDq3wMMHC
V2tAfGm9nwsOjwkt5YSsaXI41F7IW3tYQtEQ/3zozvrAp9V4bcqKapKfoDcJH4hu
Gz0hS+GMrH7Uw4nxm8lCDsqb0GgKRjaqF31t5dwU+qArOb/2btRZf1zwz2/C1b62
IYglWVRlWmKOYYMR2JsJQoJic2fP82UbT0yC7U58hWmYzICDsmv3PTgs1m7+Gvkj
sn7Dk+zrWGUriMhGOpItQzHFOxCSz9LU6Ouo1NpDPu/K5fOSik3rRoa8A/nZ1w+3
+SLhzUzbgInZ79Dw3gr01+X9Y910bDQCx65BX8LTcfYB0DO+QyB6XqGH4hbWu2zp
TAY2WNN5Efc6cX7ZDbeR5BL5zaNyUlfurYJ+so2Zaeyk9AxTMwQJleITqDlLAExt
UAOAprWZ5JPH6AOGDiIFL67XC/BW+aB5IUkxROv14Tb8tXRSmBALjsJZ+ijI/7te
Udft2GZNZ9ARoZOy6tGhVct81x6RvTSOZ+C+9QUWWwpy1lz1RxyF/MsdYScTC67X
IHP4St2FY/6B8JlSG5CxrM8nXw0bkHda+onuQhGkNw1rDOXa1fwAda4LqczbUr2/
65GD7b3iSCY3NL5AMv27fYDbvht/zuJSb9XULd4kpxhj1rc8K2loWZUH5Kc7vu8f
KC/CqLZYpqC3fRNI44DYvU2xLXmgI7RY0TH6jq+ecnv7xikKcr/eNs/ZQItF9hEx
ZJyQlYB7hnvQTWWP2j2IueQMB61N/zxOrENXv8/2DGdzeHgOXkKC7lj3tVj6RJpm
XGypj1fHrV9Ac8LXpJN/t1vkuYvZBGHdo/+Xin1/5jV7c/F1rUK9BIi8vgk4wNJj
gccBEuBjOPxN5BjC3eMK4EcUcj00yLd0J9+7IRbz1hf9lsKq8MP+ISLZedR5Spnt
L1tN48KQh8VlOEZfliGgtQDY7cbcLJuFyBfFvp75JaHftby6OJ5uBjBfMzNEq57z
WSmx/My1o98jdkPtK6mnY2O/AQRYXJvI3z79tP2ePWIVD6TdMhLdxdFe+WZehAgV
3U72uM5l4Y54riMO4tFkvdZNuFlqxP2YvKhks5f8wQ2lQKOAGhPvPsfUXHVgKkT6
on01tSSSTmbYY+BOGTMteOulCnOTzM1MHy15uZbRIFW9b9qlP4iFR7H3wjTHz2Fd
t667Vto3PbiZKTVW+gEbz+jQu3Ep/zKInawWWukLDMeyTQtYTlx+DdWb87FdO4jq
zXaGDBCiuvhUJdIGg6R7HbnJzJCGjdClwQR++urLMpVrtIN3/GeZzQ6CXI8+LzG9
LFOWIhVHzDfOjoo9rAzVPhN+LvnAptBTh7xmpaP/6KA9dKvwto6EvVBdFOwlU93e
SNRQDrCEkVyNZMP2+lXpruY577HM6foQhZu/9bLh/d97Et4m+ac6ok8Tm8TDXz2D
fk5QIiRTVXVElnNI6YX6LWvq5DFfUEkEBDEafIIbdbonsckmZtNfbgkc2Qj2Yl7w
eTXv84bvU7l9QxTrYTkeCH++gIYI0kLUip20wwzmnEblcX6jqNLFA4Ay6glZTvio
4uhCtt7EtKxMpcffZamZtZP6yqmoTMEsor4DPy0nCydETH9LTu4eSaS0ICtb0zc9
MPwCHwZc94oqzx1pXFgPKwjbQm7VKXl0tJPtbAjWlAyc2rIFUURANsM0vZA5ctU+
cY2IjpVvwkyuonnK8wr9NywI58wrpc7y0UPufbY8R2xQTffiFTMMj3bCHGvpBFRF
aUTKFH116fPs9XcNQREOsnS6HlStqlXWEkygEQM1zlL/m/4kQ1kFaKw56QtIJXrP
fqCRfzuVSnTTCiYY09eZbSLD0vB+oHro6sU7PKop3jl2SMrbAIK6di30YUkY6MTz
CepHDN7/qj9MwEZHuCvtzr1XwG/bVnj9Rpsl4xONtnfRsfhKll+ZweOd42nXrkfN
o24Kk+SSL2J7SbrSB/tBHSnYq1KXCSKP1F90/ooGy4kV4Jwz7Y0Fu46ksXlsTtXP
Ocrs0SAfh+mgurnxHalo4lPMu8CPK/UReD49DPwzyReVAXgQ/yi07VvKipNTUNX4
rG490j/KkfyGpGUfOkAr8bZW1k6mk7tsLi2IzfDjXkn5kSAih+/b4wKPJcJf5E/J
8Ij7NFPGb5f4BgpIL6oGkElN67+HzQEtXmHI3o1nhFmObhb+1P+HY0GL+tscYRsq
Yt3JZvzWk7+UYsyK3/MOOuQQCK1X6fsUQM7xX0JcyO7nR0/zclsglz5S18tE4eC8
mdxQy33fiHqJoQm/v3F4erFqJZWKWI8xhHv2mkLN4GA9S4gZRgMWciQnVAIsC+FM
vhJ4mJHNuJHrwUIL36nrecheto7UQ7ExD60Nbmn1rGAY3vY9AHxMGtaJ82vrHezK
9kfwtxKmUvh0f0fGDngRl1Z0PN8ZcwuAWkOxhmmBJYEYNCosz82w9rNlrs3ZZgRz
PUlqF+nQtSqBI/SuPx/rvBzLuTlOUe+2l6mMmn/4bXawNgcms7xn4tMc0BptD1wT
rd2ZJZz/iBEA72aMyXj5YRH3Gg/ubaJXWe1KcP0KCppJ5kOJeFGbIYyu3XrmsMdj
vRhGkLP/ZhFrd6sB7Io88iYl4tm6fsWznLqwRK9YbP8QgEWphgtgaTrIlaa47ril
Co421pes8H1Sd/3g4KZNnPRzd/qF1SyJk1+UTZGkwuuohrPlKu1ETKW9LxWxgLDV
rjou6SU/I5nbIgbJlxmEiaLXnIFz1gZCzX5ruBQiYyOhgBpKZ+sX09LA4YAjF970
6Q50JzDb9YzuQtLwEaP6VI4vhg6Hlvb2cPVajDccC//aNufjF2H2NNaxVwqoD5Fy
0LxNF+DHFhmEZ5czAXoYXPJ+yCA/eGbTG2/yS8u3b9QuilfBBkGLvQT94G6HrL1L
4AeMe0bcs17AqIKLXXTmDWvYollnTNRNeh0oDeCxdQCVyq+1TrH9LwVmHAsH+OQT
TmczbDi4zdT+EnT/x7xWbpdQS1KIjyEXkqF0y3+u+MQ39Aiueeg43f+VU+NgCtbW
EVHfiSWKNQOLVDsEj2ClbBLhXEWG/OLpGJtL8WP1lOQPp7H82gNWHfz8c6iIOqy9
HMfJ5iBa00Qam50A3eOKMhwk2blmzuesrvKk6m6E0gQkP8bcIHuQZfTlHqAF3RSv
8oboPsh1BAdSovpji79gkh1g89jtk1JnnWRlrW7NN+ZZ6mC/Ti9bnyHC7tR77VoO
SoaXQNXMmsZ15pKw4mx6EHGalAX1mJqc9twNMD9YMR7tdUlXZ2QMRjA2UhE/ooTn
bUnG7G/v82qHB4nTCXmErf/i0Jgv8e8RWjq/Hw1HxjX6CjCR0QJQSDgggV+hZ5DT
Dy3HR+V9xfG+DxIF1eXGaNUTMKNmk8xQ34xuaJvAUi+QmwpJZWgV6c4ZH8BqtQ4a
jckrvU9ILbThE4HblwZ9fFu2Mc1hXTfCVOSuk94n4zIm4xQJ7Yhp1fCrRWFn8KMo
6oygnQ0pGWN2RDSGlWOeXtL3V0wzMXE9qAtlrHaej8s2/LCNoxg+YNqqNtLBaHcp
PF8995x3NndNb68hiL0WjIVe1CPyBMWhpU6JafRmj3jmvWaNx+Ie0G5BM43JGDE9
yOQD+9Yhy0Ob8MKSd+AolX2NoaLiBxC/FBoXINp+ruxJqZFVwMcX3AyAlkR7fHlG
qfaiTsRgxL7yFb5VCYnO7txBVaw+6Hf11mkEfOrwGdrsXZjwzcnVu3dddS2iGLni
joKpIZaCa2apdbN+jiDBPv7vjLdNf2TNXswJICHAwrW3q1TxTnaV22/a0egAAOXS
0psbKpR9uSoQ17hut7mODc588TlJAHXx1BSQqjgClZwHOAWRy20mPPm3F3nYU6hU
7TC+izni7jdFbLKAnbNwELR35OA+Xq55xHZdCF7ERmthOgoxn0SMH6MS5cW6GRLl
sO6KyLSo/Hv5z7qzeyjCdGUwDrPO6iyf2UOliawiXSsTZSmEnMhPRt/olQN2rk1f
O2HwQ1wVxPXIcIoaR6xEy2Bb7Rq16tK+kycIeAoMKTqqmfgf5P7VEX2aLYOXlpGS
dnS/B+04R5Y/qH9O75sURVLAYgGJo44wXCWz2HN7ggllIcM/vrPmDGceLb5Hlb/b
kM6InJhLtLy8E5BS71zZMS6ThAsVwgGbPKnzDEl6VmH5Mr4LMr3WTkKwqSA5j33X
aysww5UiTxVUEo6RiJDr70rBkqGL12dk5UKIYGKF4peBJXVn7aX8+2nPH8b7Olxe
cCW+3mSnDdPFbx8IXuuTEjgwGUy15nMXdiPMEMe97Hds9b/02xxgsnGkyEhAXnhi
7rS5e0OOFtDHAQPp9DMjmpi7fJiYkKfAUN32BkaYCkqYeDo6LHPVQt85MWu5/+n5
Za4mDGkJb53vr6slZpyH3be3JQd9fLmvP/8xSCnOX9N9kSypuSUVUvaxJHBJK76/
aDruC5A8qfS+By695lVRY07CgCamRbVTxv4qDfbzWF0zbIsZIsOlgWTd7UWm2QlU
ozKk2janEIndv39WuQP/8iVZE/nwmVmZP0ZKWCoovvbyg7avA3Ajqn8+Kw2Yavy4
Th/tENrYTPtUu6xU853XkZBTGm+1E+rxMmBRHXtNHstVAtw3ig2+K9wQ4YBg4um6
jVyQy2HDap+Z27jhnmQ8luVbaA149Z4xKANggTa1cpZBL6aaNbXJAMpwdh8GXuk0
sKqvo4m7dCGlf0yI/plEYL0zpUUhcb6TG32H7CkpQbf8PlpNv1WT/59TNR3YwyAh
aHvmVSVs1p7+6xpX3y6iXn6b97STqjX0d46FUfHMU+G4O8kiDpk8UyafgXuahlTx
Kp2UuFGFnVXfhXYEhVGG+eAbwmGYeoYiAF5kfCrE1JaEgsj5CrFJ6aqXRd37sHXa
YFlPEuMbo2XONwnUReJdnkwZ+5IviliMc+7XaKS1ZyuesAbjj8GpzYiEri68rZE7
ws3R1P+KyIVvYVujDfAiLlCbOKjz6A6MZ/OsUuQGaMoEs848To2hkIs6Xg+Oi6sK
CZi2U5Z4mEvWSIIfIBQip+NJVLV5n20mFYYXud1exak4og6IleIIhgatHvmzvnm0
iBJQOykyyfntsv3tu3R5iMlkyWCQGs/zr4AqEwKakJW/sULFr1d5ca4lzov5HkY0
DWVEPIpzEziVTbOLUmQSxGzxGH4HnddYTpHwp6Wpycl9C8f5qC7vXrl3moWjIOqD
NG9UbhxWNcLUEegmX9UWB6FPkHzVcqkKcOmBmwK1TQ1PD5bxnz7v1Ozvgyo/PMtt
gQLytAZRclTm0eJ/coHarHs0riiyiELUuEGnvd2zrloB8JKv0ghGaTLpyRiF7gt0
/1e0GZLX6FtMPKhtYkLMgFlHz0pT5/2JP128SnEiO2pvP4n5QLtltg89T6EHA/p9
v3oA5zKW2TIp57BJk/loIN3eTuF4eN1kWoP6+rJ901hq6wjgsMoRQ1AP5KpMZLY/
eRWSHHfe+KSm6WAcBFkkD//buqTqzjoKeK32/ljKkMmyezb7WeBH4xusP7wYifEf
2RefW6PMzuIa6i3i5e90SC4AeTnFcQ+zNq87G2wbW418b/5TWSnd50k8sUL/K/R9
vJ+inq9evXOdKWgwTuHctqwNuJxD00lwjZb/mntDgjJBXEg4Qz8xj7LCe2EGh8Bo
8fWYlu70mH9uVoc5netBOYGdwOV71vBscg3WxU5AQfadnLH5f139wCzLd5YP4ETv
snsKOlavBUE2aivoQMt8QGQHkMPNC2QhTL52ijWS6E7Y7CeGhGwbVxda7ENpz+B4
rrZQh0WofjV5QI5sh7oeq3H7XKS15js/ALawCnaR0pSfvHwZaZglnTD1pMWqbD7f
DRpX+6mPBVdQPo8lG2djxW4xROPuk5iEN+qqRfWS86ALfe5Q7aR6f80EruS0pTJl
HSF29k+4YikUTFV+Irn4AJCnncFqCDzCNAznUONkkHDaz3iokwYEr0cdJRb/z+1m
lhIQ8D5pbvjrPy+3BVuI0scbXn/Ms/MOR2kAscgfmv1jKZuAHI8HOVuz/XECR3dJ
cH8xDwJKp+wSHo7xRcIFYP51UD89YMfo0JdCXJbNpdwmTcJHZ+wNX3afLt4X3DpY
fYdrtuUAjJ95Hy/TEG/2PmVJGxnmIawFUBj7UxT0y48zE0aQ3c9YooC2l0yezkgG
CDrdVVRduTUobX2lTwIk+PTNaBbhVapnYte4WyyDvdAqmY3Z/q3bVvGXX4dD6QqH
WFXKksdGpx6MHkHELQE5IOSMqs1m79LqzqfLLsEl853KEHDneqblrci5efifae8w
2uex8BV0Sf72Sn21TGimM0MgFpCcyNJo4jpAu6jQzyFmowueO0du2sAFB5ID1L4X
SdcYt68kXzDZ+k/VyX0cjzmSfk0fA/K2jKcqNEVlu0vkN1OgxsMLPOmV1oj57EHJ
TpQNbNw6dwVbtO5bBtltO97DXWmdSdJ7cI5vJ3DHYRG1kFMm09GPrEphXOzTozK1
qtZZgnL1OxFh90LsIGsIZiEHcwLE57QWqKSbuTTEPtOXNx56K4rN//76F1RWDjXp
kV55+F3SRfzhF/MWIXS/jqQYe9vR3NQVOap3N8qvtmGthLFQiZ6Htl2JkksZEbu6
SnW1jHlrqUo5fVermxD3DabdpANylUTk9dCqjKk17cSAXuHer8ML8cYgPYoN4Nbn
EDPejIOxl/7M4dNGf0wtoxI0x2fDm9oq2Hv5vdHYM/T8nqRHj5A7/jqNx3xqIVh/
Z8RotxpaTcmQ39pT4YYkV1uljAhE2W0Q7zlilx5Em0ut7OTu+qrMNFKLQpCQoAWh
pBM0dSkvRLJ6C6r3CzcBOtrUBYWFLX+7nsn7zHhwqJYce9YQD6zZsunSChG66Lqi
c/Ki+NLJRkijH+ZuNnITZsIPIkwvetG2cIq4//WU0xbh7yGsaPH+gdY3J467i2A+
XHe7CKw3Cf2GySvvsWazohe5V8tFJEg4SoGmPf1eS6s/J7uj/Uv8CSVusWLCttG6
8S/UnXeXUBLSJHVZxoBp2wcR5ATO8e0PtVsSXnN1tUImL28b2XTnlq960IteBx6Z
ixNqTqHBAUH7BSfxk5/I7tKXZNuJ4d4UrUTRkZEC+cQC5mCj/0xAyHl/ECqJfyCa
1blH9aZaJuviA1gyLRaN2pSEL010IAg0Lc7lhZM78qU1ZpQ/zkIVsSBVjbIyNVPS
ykkcZxi2ApK8ErAtrVL/w6Dz4tY9vEGwCQ1yJlV07bd0SpvMMVli6tmdrY0y1mp6
WQ00oEQ9N783zXSvZkBLR+Xk/U8LNQMs3/nv9IStL035IcUBIkRGG3+PfDLhQb7T
8SQEQdjB7sD97DnsREl0Y5pDJUHkVInwn/0wW2yudS/6K4vrxxJEUgO0HjsEJGV4
rd47U7IzZgKDtoLpw0IE+NUdQUT9tZsR8PeO4lbZeFz9NWcAqm0OTQjhlHELMfNx
PTBjOpOvJuTFONXin36nzkhJvGglhkQhM50bVw6hDueAbZRGM9rQ8gI9VktkVR6c
IHWFbrRoiEQfWuTRL8zFPWtRLrwDVibO22iNR57VFs7MLiasOz7W/gSOyBH7kPMi
w1qTpyn16bgtnRztcewlu9SPg7vxTbOVc+5oV1lbxsQy7sCvI0atgZWWqf5RWWXO
R9hDZeaRi4g5v8Vk44S4VEREqnq7Ltpd3AwLAn+VJOfOqSV4EWthxh5kuP6AJ54J
DL0qm+WBZmqCZekf3MpUOrsivd/VAzNHiyCO8j9IubqMkNjeKUKVIKxque4exfH7
SkbzmzKw5USCaB3oVBUMmJiS4AeThl+XZR6laHuN+eoe4fvJJ9ISJeUixiwpzvUy
iL2EtTVVJUEN3QY2aEFKSzkJOoHTRB2/l3y1Msvse20FDw/SdwIybDF2xnWF5rhz
DLuwVJWD3G0BkvTWJfH++zbmudB8M0XLsaLqu9ITaMgSyU7SbF+B96S1kiHzOy/c
xO/8CIxY98tcIGKvF9ZglNQnbnPUt+r/AY39Se+3LLubHkcroJl2HVa91cO6BJZd
BF7A0+gEx7GXqIbyXTiQRr8Q7XcRcxV6dx5p4VOC35pUINW/ABb3sJOUV9ed7yOY
hNg75g2/BFNskI33/7THBLTlZd2wiS4nC2hIEFpsk67Xplt8O0kJ9SSRaYeuueI0
xmJ266lJVq86m2Tl6xL+wcg26+X2D75saNLlpICUuzmj87IJ+ZJwi8KeMso1K1zx
rwpfutEAbQXMbByVluAUL+7dFmiEjUtrE2L0AxqkQbKfG01s2K9kvfwi8zVHSgXO
RPlbUL79cCWTL7VMEzVkYCPTcirzEXl8ZlVnBqMBokvVemDsow7UpYbO6zfBP6OO
ZHlIIymFMNhwOPIvPkUHESy+rVmnSf5pz4ZBbXyvzFUnMsGgFuxeyIqo+FoFyEvp
phJHnD8jrpUxMg+KXcXxL7qKJ7I0TrvnykpysXH+ujzdSY8KoCzF0B1SGcGhgVSv
L/nf2Xy4uGl7G8XLBu5cDTTEFJcHGCn0RdtOn5ftwZ+Xzx1ZOoUrVwLBpzm0ilKo
+dmy8vA59REr0xnRF5Bymr7V34srgLLWEGlc+CPtfqI3eq3mSDuGqyhXGa0eAY3f
6kkvmS5EDmrEWOqB+m4HUBOQxHLx86V5hZBBLcE0O3juKU+Y15cMBGHFo8uu18Ec
hawtJkbar/AJl+udhIyaxRX+mIBOOsRCuf4aURyAqeXoteQyaLkssL7RgHDRcnnp
d9x6/Lt6WwlGBlsgkqVl0+y2iMRrS6Q7fC4T8f1EIDUXKamBYfHZn7dTssyDIoNy
4tyfRO1Gvu/wrKR6ug6kovNzDWFtskv2MCJl8GdTENzHzygC5j4KNJcetxnXxzTV
AZZYBUI5l8RLbbM4vNYoTb9PTeriIAOSIJquJ7yUNCO8wsPaoSqFd2MDNEu6qpsi
6IOxBy8i+ZqVYYnfZigR2yVT7FiB4V/rPXuvaGVA1SlfEbqp9ckngyVoOMiiopFx
22Ut/bzcveOppPcBcgkJVhGx0knFoYtGFUSHBb8HNl0kEPsoW8EFbWQpqSX8tGuz
i1lmMexu3EAo4J63I79EryUqFDWSaV4A4s3sMGltJe2NmIbPcg25yuI0mRWKidko
NcrQzX0Cjp3pPedj93YtOtdy+vgKMCnuBRiLVsY7rgVtsZCAzoREV7sOw/tfoOJa
xXQpXbH4hae8+kWSr2D4DyoQ66ifxsJqApJV6zckqk4RJNK31Ev9VMEEsZS7spUg
CaLQrE10H99NyJNcjOMDUHMwS44ZSp9RgAKGNUYUkT7oG23YZ1asl4HyBfCelOsx
sxBEaWhfWi5fFT+zFbFX1JUsycixwhVR90pq94ZCoWHcaub4F5qtd7RV6ij3ylBW
scB5qdjGi5yRj5JZPMkMoVL17m09QcYoYIzh8Dsa5CFQyQ5cAB39tFevimVCj86J
l1edKvEZWjsN5wFaN2Cw/CXcz1WOAeZRU22mTs+xHozRgtyFiLA7Pl6kkSIaUGxy
i1BvDHAhnInwTH+simI+yc0XnAd3C8XLT8MeUWyZampWrUc1GGlpdrVTsbzCi15d
Jg43Iub1QTys1pSn1xNFvHMQW/2ci8TLG8WwHQiqKzttK9vtWtNPcpFkiA3VYp/V
SGV5jPzVcaVy6rrtlJdrAYW7zI93EATRvhhqwmoREU6snAN2bg+5vb34yWMBC5xH
wCjBC7XQTmIZytSzRIaK1rI17fLOKC9sFbv4TAyGu52CnzLWf6Zu59rQ1geLuclj
HNe5FTj25vBbhDaGr6kQJfH83EFQ+cjM1JszXQFh82rc1Ied8Zl2NCdTyaNchky5
U+dK8NKJLUq9z1OtxGAsw34NtZG0V8qCqm2105kLeqq0cFtxM2CZV+6dIWlkpxJf
ECMxMMINZGf/TxPYLxNtRrSJjb2Mh/xzyswBU1BLrCU0fqVenvm0p6ub2+qnEIpm
pWPsGBex77Wy/qoOmLo7X5BZuZqTPOLl3REIUFnQHBQgZXYrh11Fv2z8FJQMa4An
GPhQuUbEQ6mj3pqaozlvD1jI+79MY7nJTkngbJ8d8Mf3hVURPS774dFVAvRZGl3E
ztDPJYQ5D97MI8TBX86b/Yj98DTIL5zxA3NWmg+N0ijCSpEECtm4Hx9S9chmojpx
im2zz7ZCIygUOkL4oOmuwhuKJg8ureG5fWh6kmUBGhifXa4GBO4R8DFl3GA+RUFo
1noJCga5B1NxB2umjDQKwfUb1iQ2rJV7wO8lzzmiLq5iv/2s6lXAJ5XLKDVs5onn
qQk+k81Q7g3W3obvw/9QHxK6QTJ+30C0DgrG2fGvYGDTHM3cax7QdjT87G7uczEF
LOFhw/ZxWgKrqepQhw+wQw6J2rZ/mbot0Y5lNayg40phesGwlY936nhPORTPyw8a
DMMrOxFmQ90U1kHRtdxcW4SjpAs+W1Gq6+jEp1MRDl2L2petRFlBbBZRVtCOUdqQ
1a+lQTbKasyykawqwTq9Pp5feVq4RGTPlwr/3yIXbUnehzOf4t4TfziDi5mI+hzc
jW6vySp0jMWsfQZUoDy5FnzUksDBLZ3qZ0rS3LHSr6w+WWRtXHliGSCRfsYrrcTG
KlxHMQinCyHTU7J9DjLFryu1nhAfG0GahxkJPkuitXYfjTDdXiksqa/AqxdWNqlO
yQ2ZgMZe8IXgCGwWKOyTIYZStwiP8GX1eWqb8VE6aY26CXm8KuC83zK/Kk+iN1US
MeMZ4qLf/RIQwMw6CwJhdU4ot3PXMcqBDHQ9D8L51KoD7W2W1jwzZtWH+Zl0UgVY
7JzHCSmeNk01xnNF0O2vqqafwr9NePzZeJl3Ya0gIQQHthtC7KSggXb7j6Xb+qzo
6DOIq2xz8d9aWSSGNUwn34LKxic/66997Jn8HYCczS9ytpFoLlZZkb1AnkGWRZKS
eSw+8+eWgdxqFzdn5MS90Mn0pQG90HQEmmS+8Te0spxuVHXBKW9ssY6tnIwvu5Nw
kvDebscd1FSYZ6z5jS79axH13keg/Na1ho23loT842fdwPLxyyShWHeDTBft2T3D
T/2nww2rlN5y2310dLQ0TAGm9zcZ4AEwemooWl9qmJnyf6KYaa4hhyVgcRM9HMWB
Wr7G/sNIaFyfzmY+jhgOFjjcZ08g41FJgxtYDAJV5Vkmdt23iQTF3zokgF1X3Wmf
AEzG2tImcd2oJZyPdW9Q5f8d99vwFQn9AYgLUpQpltIe1KoYL9q/19u9fWsLkWiQ
gJUfarqwJFozJtOCg5fCVfoKckeS20RDmAOaoqlvVmHnOOu7yuLjbX1YgWAYJ+I4
+1ANrvkGPZl67oDKtQaL99mgp0zWQ/8AVlxf/qA9F4UNJ+Saq/5bPI1ne8ES2I9k
iXs8MP9m6TKqvGGLM/FVs4uvKoL3hU4r1Q6thyJmq/a+06rYNGWIfWqP93dJr7Ib
QRYo3qBtL1TvQQjtHNCLlzjUQr7dcThoFDp6UNGN1dDSAxrXJnKC5it8DxmtdBws
U2Q1pHdp3lZbWu08wgG/xH85bFz5NOtwx7J6ALiFtkIdkJkZyre3twO2c27YsbEa
ewhbAXYJUKuy/bwQ0IjgBoU0z/gQqISzDW5OjCZuPI21myA0lQjpzeD8BX3teRtA
K+E0eCnGU4DiTtZiRbw1kg6AE/1Ljdh77X77KRY+IP9reql/WzyXY+Cyhz3dxSJf
TL0tkqgxu3++B5wd0sCVUgFU2oMdaLOL8bWjyVlVFj/1A/+znJNUzrUrdTg7usBl
iV5Yr0wD5KcEh5a/8Mvxo1mBKfc8kEcpBtTsraYK+32HKI4OrMT8vQBKaVdIliVj
CBeVH+ALgu0/NfqZ5JPXJySoSdjdVcEbLi7iBIYAhtrTxS6HiuQTySAMmMpNFVTc
Wq6/wFHvuazXn6vkKoxTf6u5APs6ebk4V/WMAJTaGzupHHDEigg1m3uUZTxcLFvu
guXb5mJpEqehTVT39ESqm76l/d3FqiCCwAl3j5HRXhSHrTEb5pyMQLTU6IVdEtq1
XJUAzOCBs72uKnpYar4VuVf2JENW3+TQ6SyP/bK6FHRB0XUjN6yl7b3TuyHTD6WI
fTZ5smt9YDhWRuUYKO6Z1bU+q0emyUFSVij7iRNBp9u/nnNRbs5UewEJ0OKZHPKR
4aqMaOpaO3GmGBFsOGWXgpGSM2uIndZ3Y+CBdyiwFnImom6DHNZ9WYBuOQ8xuQyA
xPzFEV/iLsx7IFk0wMuevTZoM+qJh7Khxy/a+284m2CFSa3Vq9cQRplEigcmLDFj
BQvcuu3bSODMK3XTCmW0yeHBFI2UO/Oha5u+wgNa/DPR0GcqmSydbB+MrI2XrmwM
H6W6RIkdPL5xFdY+3kXgXUNhecDFXGv0ttx8Z8w9rR+/+ZWSFdGi/oDg6+Fbb/Ev
5CXu+aRUUiC6YgzHkkRtesKm9qX/58FQWw2FB3Abwsjq2Dw2E1i+Cqx3cXFtvSHl
Y9SKaSvq5Hcc4t/D4OM+sZIhFh6Tp+/2reGtpG5f0EFJmaUToMF+S4seU7tRv4Am
uOFeaY9gTKpibFv9Qm+6cD0EgpoEp/ZooZ+xvk9Qwuh1Al5pjOpZuBCsh61fbY+K
11vxMM3jLdEaW24nJDUrqhtRxNasuGjyQWXXN6m09G0IvscApu32YeZqh2cYZyhT
jthK6pQUNG9jU8LbEk06MHXoIGn+vDXSwg3/H78i4Kb0F6o9Veu8qeolx/8iRJ7R
GxcMz5i38t1E+DtkZ/gy7nlUOdrAomLUKbAHbrBu4IC4JGldwAa6pkXA8Zh3h2T7
dD9jJlb/jlc3c3lGYW9X7silhLEW5pkrwJuQUWnpZk7qoX/yVBQaEh0+nzFz9Q4O
tqCdwj0pb1ji53yEM2l93/RiEpEPG99PEt3GSWx2EFTgYfrzxqrJfazTKmIWaALV
+QIr0MQSk0awEpiLozgQ6HBANuhW+DDDYO46IX47AJiOr1S6plvfcrUCcH9yc1f8
FVzc/yPbsB4wt2rtktmimESvEXUUbRvVzePDYNUoeagQejt5ORF3GACpgNYFmcjh
CJmh5cUncb2hIOFPEBSCg1Ae2Gn4fRD2KtUwyFywXjuRyI+M2johKa//HxOEr/1V
FMY23T7mPqKhbTjG7hZnWNP0yyb8N9agi4xF1pZOgPSqz4e6M47vKFwO47HqOJrz
Dh/DwAiZqLU7nsdnYZn9x7j08hQzJurBOh9h/GMBT1TVUeXpJH7VxAIdxJ/Ez+GV
so5Q/n9dVgmE62MASuhMni6zmnSKv3h7bLIHU/9L4GcW+AX2v2AGc3+FCdhNEbsU
X5jmVNQwLfkEuOFBCggPaYYlKJag2/NoApBFSTPtpieIIaiXLWLQ2mIZPi0nm3gw
9P4NksJSkMMGAE2/VoPC5nsSaZ8D6BBO5uWCqsoUyTjH11W1OfwdGHMhPCoNnifC
hD5gnaKjjTsS8j6LsRMH+9LkrQo8lRWGjMglpHSpAHW93kBVq3NZplp9lzNTAwKp
3g1pv+isz8VblQ0AfDUlgq5yrJddSsrtUkuQ0X/tWGmjZAnS1f+cnkwWuMd/C6TX
71vYXJ/CZ+uq+o+UJyIpyaO6GZ3AWQ0vitujD1NfAro1ZlG5UzxFeALJQjvzaiN1
O+MMFYQ0W+GN7W6qeQFAqQXPzERRrSZ3Yyx80GqHvy4cNm66RW3CQ+YSoTiuTCh3
GT7Aj1dw0ionkgCYYmf9Eg6ZzDSKzUAJqYnt7r5zJU8oMtVOev0fpAgV9ng5dc4Q
q93CGY7WKXNfPQa1J51nD1tE+ZBgtkOFkrVi6iEOyX9Orxp3Ppu9H+6Z9oZrMAD0
vjNa0w8Qm2acCv57jGietYG1eSrnDprak+DXvSag4b2l7e16256ikWFYJrdhDbst
XxGnGJWeCi5NK7ZiPKX3Sr+Z44sw4CSno6KnlLtdFz+crfRm+ihQkgkHFNxQ6sKG
5uKWJwkuUdylzNqLVVkA2BuS2fgpW/lw0M5kSOPpmmrvmIWnl2WZn1LTozhkf4CY
rMXzk9/qDqVziIEo6upV2mQQvNsuWsxZCRX/31RiZDv7bguS0iiI32z5RKiv+asu
yFatO8aI0K0p3qtUL3bWzHPXSWRUFeY/s9TSH4khNVpwq7tkGZfudrURj7eavn2K
Fm36jAjknZL32PsFn3mgYuirl3z1tDjBo6VDHnvsuoLESqkvyrClX8vxr7pEdPI2
gZ2KTSqLrDLG5aEfbUhz0zr/p2yhb19tqoRFONQFhZMCFHPTLhSHWaAbd1VgXcMV
+/rCUylYELfeT1mafbutmFFK2RVotKD143wC51B6EfGRVl7pOIXdXQ60cGDQz1MC
j9SvOlM207w31wD51jMTgppQCJhSmKvMYCpMb/e9qSPi9ajO6SfBzz6SuJgDUyON
FQFo7/XuRjuEwVnpnpmQ50Y2ar2RSWJ37HPp5lAbVKPwELLyWkA0BiJ6XeQqmoAX
IJXHKJyMlmCiNFzFAy4MzVwQMZmXxhQ6OsBlW/EkFA/I5IyrnKgp16Sg7McP31uQ
kJ1nklbA76ZVQBIeyO4t5JzhjpwVZT5A4dfe3HqKNMYWem4wczWViACpS8OXuRxX
93titYp/XTcXTPtc86GEs20MbJZrBvVC9U9k46KN2nrRcH5zWxPgqsMEYcMEKpp4
7tFgd8uT9lMMnbITbseuzs8aZk3+dyYG1wf9Ofu3EFGtELlNBqhkDlBMnlX9m6VN
ECxzSoqyOt9T4k1FO/iBsjWZIknXTQSUr81TTeb3w4u8Hv5W5RNMmBo4g1kI0fS3
/ZogLQ+sVoPbKrUEJx5jCGO39IaFaVq1SPm8FhFgR4yX4Fte+msGp6XJZXmHXMRB
pazYpMyMlpzhUAUcVG+rJmPZJ09ZsFF/89JtmcwAPTstgmuQo21TNIsXjl2/4n+e
BFohStq9q5uZk9l9pNiSoAEc2RuV1KSdotyqWtk0GXIgJWmP6IMho7o0UNjfdPm+
rXAUYcb6+TQpt7ZIP5S8dCA0uoSdGCeMsnJ7o1K0tygoEJJo7XqpVFFpwuiR55b8
6V+RixBIYbdpcmgqSixeqJUL4oO81/CKqzvHwOdaDrRgaK5aNVibloffUUUlrx35
IfUo36BE2PBZFY1nCyP7yD7egaNJq0wy0VH3fHuT61G129mWS9vQ2odhizBgn4IC
UvsPcVy8OrLy1zX1Hg7yQn33kk9YIDVHznF4+8ZEF8LsKqskXKEbh0FT8ch+lojz
Pm4TLj/PmA960iC17lwEX6kI+17XpSMEC74uCIotoJXdLPq5OSUUBOWzW5DLE06i
X7qmwN2jqaeC5WKex9lRvuv8jxBmVKZ4zBOvVzPMB5kIqHvq0Rgo2HhoUPAkVzy3
D52DWP8jNxgXyiA2iY54VFZTKSEu+ZHkjKebWbc+hOn99ZaHpjMqFPE0412IME4w
jY8sAniEJwKJUuJPf+K8bKxBt2lLyjoX0tAsfmYwKz1PmvSpfun61HjbCkvLlcwW
yketqTwrEgsP+MAdfNj5kRnOBaJqSsONV685vrlEIapM4zIo5428bVLhhJCS6fEG
4UWpyIp5Xb6Y3MLnQV3U9AFtoym4pvP9S74uA+TLA5cvvMfLqNhnhujpcglSPzDh
zlzlKg0GN3/ouO1UfmKmolwt82mvxrCv4izgOVdP43lm7MaMs1vMEcyfg2LiiDDM
Dwds11QvRhs6A4au0VCdEkVIZ3eioetIO568bqIG6KQgcpHg1mp/DEXk+PZFXSLz
XOh+g3pSOd3ogLtzzZpOd5IgMufN6Vs9WPLHYu3hl7VRGz/Fs6FsMk4XXwzoC3IJ
xziti0wtCY6rqteOv1+awEUY0zvzqtfeGS5wRLR8hjcGzcSNpmttTBCAgnnp1pnZ
AKCU7uDnrrv1qKfkcQG1C7dzjmYcg7KBqobkRjQmUK7KXlEeAD2Zft+XLjzLmX8d
XpimWpiClWuEhDcRVg6R4BSs6G3l2ykU/8Q3iovizXOiRHgXYslA+7BXRIQWi/ju
v3pT4q21L32KJj/Sy3ApxyjtRpY6aS712ls5hUlS9EdpG/naljntH94Uu3BXxgY+
P94yzchKAj190MkkrvH8Tq2wwswtgL8NYrMPtdHA8RSjg8DOy0jWgBlVRecRWRTw
1xuR4Ckt82IVgzOwVSdPhqsTWr2rnycYR/qhrI1+wKGTMlwe+3M4yPhjet3yOOOI
4eLZHi57/RqAZP/JOuVeH6cGZxz0RABvrZdhp5cLArYJgVD/pdO/p284/iAFUk8d
LCPl7yAsRvzzNPoWTSslJEV3lTdLo4pZLNWNgo8zxiscZJaaeWVMJ8M8aqL7GSGc
J7uN2o1+Y6q2o/MagZET1lAlkcx0K8yKzk4azis0sHfLqA7N20Vy40DL4dLw4M4g
8QLcqH0Z3WXlONHr/a9QnC8aUp8WkipK/RS8zIf8GbYvcmoRZDe1eqmghiOCawqW
zzkrnCFbIisJnu/dDeGGa4tZ8xdj3vzdaQMW24EX4DRUDCYUgAwAnJ0GTtKJNFMe
9X4LNrXlh3gI4PRiG6kVvN6kzFbNWZWFhP559SDqahthtDnMQSxl/S9dC+3+EtXl
A30xUwwt/jKULISGkaBo4zk/YuFxqCiqPJsPU+ZNwP+EbQxrRXmxql+9ITsxqxZC
LKK8JJKT08Tpx4yqDWwqmug1qu78YylcZ0CiJlU3D3sf2Rb5mg+Y4ASgU+Pnz1TA
g+9j/WuviKrH9d973s1sqaxg4XEPfnSGOZ8ty/sbG13HK6uEe2ITtrH8ig6Ql0lg
as+EvOj5mcmnDytvA1Sgm4SBzXBJLaZZV/KwVf2esWFM/EHWDZH3Ett2HuToDDSO
3r1u6+0ky2t3LcepcAeMLxIhrI9fV4WJLAWuTx8dqBGKA/pFfvcfaQokE3I0hWif
vEMDX/km5//KBIOkapNUlzy4QtVndqWUth7ettf9FePItBa7LNcpdkD6n2jcfdtc
V1HLaJjo0L3jZWjzB9k2zzxFbU3QEe3UVkwOGRFxhOUcKad5fJpXPXhQnR7DMB4g
GUwOg6oBvS0Ny6r37JUYKo2xb9FLobwp8feqWvEYQADKZ/KGAQPoE/89OkaslWwC
AdduCr9JSP4TNZ5cRzqzgauS+3vObPQ1ifXTEzQi8wGD+rxn2KIzwe07fMwJOhIb
S6EWGxgk+KpFfRNBMoRzJTnngRIyMGBK01HP+hV+YTro0H/TrwJaQGfeTbHHXagl
9YHJSRXhIvqFx2PUXJQo3p7TGdSPaBO035iesdGEVtskPFJ0bYJm8v5nR8k+bfRV
FcITBSST8yWkPR5U1RW+TjkLM8dQAWTJhrEgklJK3X2lK6msd6QTjWSTMCeXNJq5
qM8xFr9QCpxZO/Scm49uLjFcCaOyjtnUcIX7jwNhHz7mmrOmh3ZzIuNm4ZaLgsK7
laSyjCV2uhzJTX0YoMUu7IbO0W0JkrdHuhGKrm2zwB/QMzhaquwDf65CmeNext9O
FWaLtbmx+Ju/FGUeE00yB87XtLHbtyB77hh/Gyoa1y84K75ta4j4v74udJeaBCd4
TBwx97mAqhfqM+jKeYI3o1hxsp9wugOIxxsSZKAljAea4PVN/Thf1+61SToZu3Ig
CSZ5bRjks7Qoc/y8ndHFjlHT5ASF7G3cD7uUbuRtFy2mpJpfwJOvSMYXo7SQ42mE
RiQBrQpF13p0oclhNEZL1o8MHE1l1+U20ATzK7r8z7745SV2BJkXXjfyZaU01LU2
LC/c7nJYlOuEfmGy2fyqhy85vYxxgusFivMrC8IqElima42ut8lwsdHEWVhvvBbp
0Z/AVNBhJJgNr9vX2RXOYzBPykwvR6kg+jxuIBGOLd94HM6nzHfL5DOZU4t/j0jM
hJ+G4IkJ7NkXZ2SpSdEi6CKx93vJ6RY7rJpJvAg5JL0HTvtRKUvxustdNY7OlpHt
1kPOM8fufmB5Nsfnq+PK0SQxEqlqJrRlyvR7tu4YMGnKY82tXPU5BF4v/qL/hEu3
IJyG60GfmlvfszjRK9hQGL0S9dLM+46nhHGPCosHyp5tpKSqAv0e7qah6pFfhWVD
h+s8j23JXnQwOJib9c6zDmDymo3w7VeM2JdqNh3ZL+Wh5LFDRvSGbTMYQ6EKNvz6
Gzm372lC+Wn3drgrubkzDOZEsKR1cu0H4l9aQHpgulIju+4gRaTVNurPlV/z503N
qsskOUzf+UPLhITNBM99gUHPJc4gAlkqWU2HNL7XinBLkqifwJBTU7tawbM/vos5
Vrr/OxmDvSwvRyDQbHUrZaITSsBmJcSzKPxhBSIcY35p++1I2XBPczsUMiCx7bfW
OiIfXU6FQv8EjUDGuTlxq789b9TufsIGBK737/FGHZPQmKq0hodkHi2Pu705R9md
AXP8cKqWwiPPu+7CSiM8Xy4UW3GrU00xhNbeSp33zVzTJONR+BdEPeR5GYVZgFwb
wOfSdtdIUPmFW6Nhh9d2dJhyTPSnznATKjwGoDD9ArC5Za/5F55NXivg8G3TUd3D
Izj1GgvVT96EQTUhQaEkhCKAF8D9KTmYi+57uB1HwLZW3XETr1Jumn4HbyYYbUSI
GU/HyvI9OPrupsB2ZkBSE6VOCXmZU5GMazbGgnDoomRHdwcNyc9zXlBEjOIt8c5g
jkOWx4D/V7tYf8rgygtVEHoHLoOvHtuDx2EtCYNdL0eTWRGnK11Jsmj/1w65+Bfb
NRpamGxgH7EQ4xqKr9RTb7IgTcM9Kk/4UHyz5k59KJBx9JSNP9sRyWK5Azj43I/3
5u7LIfZiF5wanKJtrRXx7ENsnXMi3m6n3WuEOMcXpB/h/unBBoxAQ/cY0iYK4nPv
ksCwYKl+IgXRKMbTaUDCofdBQn9y8A3IAevXrCJ3jpX9Bq8ZCPPmMaxXkKXPX1vC
P5PPXHK42/EvbuDCEWCTVHF/xvGHmvQ6A/z2nY2FQtMUEJN3WXzbLxQNQfKV/dbq
DQREoSF7l/kkMhyZ+kGRwv8dHIwOr2HRxwrtFLsabu2YMRiJS1YhJOIkNB3P/JHO
zSjrADhhQGg6TK6Jka1owO3aPJ18y4VvP/GHxLFrFLe3wjWdniCg4lh6qVt8UVMl
BGNR5OveIAsOd93dEDvmGw0opukfkkqbXIbzbpfXlFXsTekPSwkmn1fTtODERsRk
2TaZmtrRIlgJIdIBEJ/Fue3+aq5QH1uEFww5StXWGHorcl0DzfsHFj6dXywDjAzC
ZF/QkyT55WaLBVuJVaf62pGJj2fkzRhIKEtxukEi1gqU3nSjZpyZUwrleAEZMRW7
sJ24KQxYXhOugQrypfMCkkJs3+OoF5I07pY1Xicjv8/YRuGmXmfFxDp+EsEDG7MV
+oMVHQGUZjwzklqP/m+vl10/KLPNepBqPt+uLAd5U2zQgK8PxIEMWe6b4dET5cMa
YGuDUWHlVzNxCfDFUgybaNLwHbT4E3sYcyXS/lLbNBpu/UjDHTbc/OEbiJdvenx2
ejP1CcGKJUfxkGQrw967E52tQwH6XODEqSirCZdJaB9sYDqnLOh63q5dbkM85j9M
FFPyJRz7f5aQSzZdEMS3jl/Z44l8cBfUQ3KibHJqDx9uQEE9qgvkMr9Q4CtZZq7V
R+rvxdd0AEpRJTAFdirVmPP+ZndrmeVvyKjGsB7vkHb7IA1Xoc/Wht/Xygt3hO3m
/6jA8+bNxhPwGYGfLGzyCtZW+jT37v6pQiulxXuYh3k+zdvWP09mUqwmmuy6CQc4
LD/ggjYyzvNRfIYyabD7i2FTNuPsBqvg0sjOQQLErHZcgjgVeK08sGgjbBAKa6dZ
3m+83GnTvHjMjgKg1dk7n5XYoePuVtNhjAYJ1l7lJkjFrNwmik+9qDX9ZDgna2Rt
eIjbHEJCZzsJGuwDA/+YMzayH0UMDfWI9zYjiDHERAQUiitqtmmdJeSZgDUV2iPV
3Eb4UF1KL/hMg4slNh9qY11OtzmpZeBCH9+5dA2fMkE5jK0+MFUAveIzwnYadaHS
bE0SxHBrVM6XetdWjvMUsvEWCJnymPuK78yaZot/Xg5IEfv53QUBoUpvM3oRezj3
vHp17YaecvtO+f5jqzBwu/iXwz/oacBlh23vcV1zcd3zgbm5XmEGfIqThidQ6Cuj
E18pigfRsI20bM96MAVqxZgktmUpz/zxhGS9Sp6KdZTocfoKdIeZfignhYmZzbEx
iib+OeQZr+ZL2PzXzexnzlZsZ0ggt7xOSs87PiDgYPMO2eUKsfeReVf36qtb4k3B
fyAE1N0AyMZpEPxFwJpKDXG2/lrhGbhJVSU5zfuIxNKk9Cj1PUw+100AWOM4jPoa
TQueMJwnITbH/2bKvnVTrkB6RLYg0W8qy3QvMxsGSDPuBR5DvPUEHd3IBPh0aGFx
muDd4kcemA4Dp+wTv4yv4Xa1xPoP5z78rq3uSzBDyLRUEIBpMPVvkBcZ7bSWts8z
JeQiFSZYX1ZalbnkGWJeiiUvWxpSA6Q0Q4gv5/Gu7a2ezEzHQ3W9lpTDHtFlrZ0y
CgpViB1jVo+nXLJaD+KosIGwlNLYQvxg/tJWpLwc6HrsepQBpzW9SFWkU6d4aq1j
T0AyDGr92VXxDu2eUwtmIy9I1TsqeXNgMSXqQ7G7ytsGwpJapHMFusP5/h0yjjac
SbavGta5Vhfvh1Yv12fLzZ8jOB6KcXXt7gT6YHEz1yQJ6/wnQHYGi1s0RCfjV2so
Y4bFFjLcDZU5YBXQi1aunpYFcY2yL81/Td+v/8Ymj1t+OsYP5veS+1VBqzWzzPei
tdCl0vIw2M8eW1+T924/070Fi2pXShnyhHpiv8JDRa4YsvF6PX9NLRBYBIMhrAQi
1FVllBnOaaYEhlkn0Axht7lCVSVA9NR8sL+1WC9/opGUghTwUmrvwdHPGZ6L/5p5
MVbq74rzLGfUG+7QI8Dh/AI5cE4yzOD07uARf/jJN9qHfbj2Y+VmOYSmTF286qg0
56s+3N05jz/6A7i3EgPUy/IUvWZ3EdkQmJUhkX7uULwQoyK2XUAFss7xjg+6bvzh
u4a1FhSGDv0dyGHyqMRPZUIRWrz12ujPFgiDTSE1g0kxw//VUtKe+Kkx+2BkvY3r
QxKZDX82UVx/7WLcv6b95idku1yT0P3+wMXFIwfElRSMTB/rCiFIFzieRThslHGU
wzZkMxwp5DBbZxMr5nHdWw+XQW/FszIIKw1WPgBitxUz8Jnfh+2mrAAkFjO96PoA
7Y6+YHTNDmjPfQoVaVGKSxUcCw4b66v+rSvJtpP2VxUip1OKOX2rK2LNVRghPAlj
PHo0AQSWBfXsK8Nwc4PLI3sn2WeLOlg45Inq/+BI+qRcewyOWR/8ZYpQeM9buj/D
X/NIroDA06nfn0lfI7rde8ZB9/ncoiMdz2KcpA1QA8r9BNZuJzhDmNM9ZpSaA92c
9AgReupTTc2KToUjqhpfB+2MeK9KkYDKdcBN/M5RDnUPZZ4GHZ/oVVgYe5TkgdSg
2wW/PC+KeQmHRMTWY3//rEGB/vj8nF2X3h3AY1tHzA6dy0MevzISoyyYXBCm5/C9
SKNUjWZ6Q0QoIQFHK+LoTGo4w4p0akHAllhfVhNqarxV/nOdSttS8g4tNsMlUf0x
/l4VMYAPKom4Z1X52KZCQLv2z/OdrI2A4qRlIxl0vYRP41BRXiu7rq+X+7EmJQ+q
1+yiN1rElBPwC8DtI1Xxl1BhJHHtRIvt8nqjWVWAw7pFATaWH2gZQLXB2+VS1Btm
2CovNVsgN9k/Nj/3GnBIdL2FfmJh3anO+ugXQVv4DRezaEX0K2docD0AeaJeOYTS
/8jDwg+UOBJAsrzesLNpZyb/43q6gAhQ4aektw4G7UffBxJXiIPrnIkO4NQ5l7rs
ZvocFFmwb9OkmU0lgKj7MZj7nH29vaQfrmfdi4V2lqc=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TnAl2DexAcT6xrwDzAldu0dX9HH1RQYn+hKz3K/a/4fmIeCGZnxoJ5liienvxrm9
blczhCCnCYnav8adl9QgRaf0lV8eFlg3rkrsdnHrr3ozKdtKeNj4CgvCVLVKcGD1
QB/pDRIUlB3d9FJQx1guQhgB52XiiOLwG0JStERebw9urY7HIVjtxzWpqIh2agHv
e+gqFlYYY7s1LqEOx99dnTryxIpyxJ13V67DvLYjN8oaG3BW/YE59uS0hX6djbLL
PlklIl/HwLyeV+JIBOzm1lvuhItnI6AatOmHF5z19yos9s8WN5/7wzSXK806DTs0
T5ndrbEGRmTkFf9LbcltLg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22144 )
`pragma protect data_block
bCcJkFh/lY5qdjB1lCapnxdRnw3m1WOI4hrLVofVFSaiuoKmfeKsbcGMp3ndUl0o
DasaKGVuFKXac5+IgLUokGJbRkmWSdXfvcRc9FS+lzOIdTuX0MyI8jhmXWLvilhL
wBbc/Q/vHD8rcQyfPmdVfOMaGV8zA52kmaJF2OyE3Im/Qu9TdELYEM6b1KnOn+zS
+hN+W5TXysf61zfvXJ15+GpqvpofigEl0DfgK9w2a5uIxM7f9m4Mu1qvpYKBWyV/
GeSuf8fWbmNr4vr8cetTE0eXWP6zA6utGi0CkoGHLqmwsRNRwHt7bz30+f9kjaBM
nDJ5C8LWJR9UazVg2N9mqLa3PrnHVcoxfwSOkx15Bb7JKdpEJxqGH+QYk2MxWkQz
hYZsR+VVURiTW8usj0FwR7klt/GoXCaHGAr5VnMVzXpD8eFL7XMbZiZLuKns6ag1
+xrTdGUaWfEtCKZVRZT0n13iQO+TPgPsjsirFuu+V8puUtzDfZ+b2rC/NtOkbaN9
/uy02FGYEFZfxgK9GKRLxG7OyaEo3YIDf5CHgKx4MNS+pg98Y05YRV/aXq7JVYQE
/p/9PEwK01WvsE5DBVu54JG5qI85Lr5NrUK79QqhBbS7F2/WS6LZ0uhegNmgidwK
2/qj906ZmcRxU9LHL8iiRL23vK8ZnXvziDCkfFRr4Mz+zAzHuwfVKa7extnuYjt3
6Z8z2MvALF92pZsB/nrQLr5kdxI3CHNKNr8/0lS0mmyLTGpFFOCt4yxbroMPVon8
W5G1jD6+SjgsIXg4pl1/2OL070SGGhRf6du6BJqaAgOm0OcSdvvHT3r7wYwcCP1Y
9mSARl7CgEGplYwe6JWqn9QZ38OUHtEQTycsxgowpPEdWKogABDadbHOajfT1y51
DLMSVg6HT+nbosz8LHRFyIE/fRgApIszlbPWIwX2XtX6CYA8YSzYwM5pd6PVHOCd
N8kHzU/PrlRxvTHSB+mueoip0srhE4ueabPsLAO9KHLWHuwEEIJr2pOt7DtBVR+I
W70oYkFETYZyR9HPULZu+gXaFR0S1xNMg7ENnJRW1Y0WOwBe6UReJ7zOzqbrSsOp
Y+2GPpaI0Ul0eWcePoyrM6xzCGTJ0gwZrgNxCpbHWtxex261e1LJGR+iNJa9LhyI
nsTj2fkLHHaGvpj7P6NBG+Zrt+dSyNVLZRkolRJ1cI1eK1LgbqNuufMkbQffnQXS
72HcsExFw+fVrYwoMLjf7VH0hYQALmYexwTmDyW24CgpxiE62W60cds83HdFvogf
fDGqOuKwLgI6GZXsBsvwx4CseZU3k+rc70xoA/DtwB2XltjWanZNdVTGVhWmg8Wx
goGDbGRmHQCdcneKy/ZBGfQLqdgAWrwAUv4szTiN/AUmUPlgvFWjpXVbLEoQaa3z
UkeTH0CLTzlHuGE4oGZBrwgn1RU+j0OEibMZXl1cTezTuLUJfn5CcVOYvkheNaF5
0ESyp47JjbfbwbxdnDysPO6X7r5K4PULGmn9KiQ47kNHT54Mth4WoeGFF4Dg5kle
w+Zntub1xgy7IJ9vivE1lFy5ci4H3XozjEgNvoori+6Le529M/MadTvhRZQhsSp8
dC/ieHyaQ1XwFtXyikVxCBpYXsqkd8R1vhhtlsSRbOUF21PEieRxaISQZ2cXcHzc
+zM0/dbC4jyryUK3mzb8BsoZTGTvi0srkIO5RzS6oY7AzVxt+MjCZGfGDcDbo4m6
z1Wh31ft+ykSrvqTMCZNNTid/x94Jbf5qNeZ9xZgm4kTCXFlyvmWBXWBs20BpY+Y
v2YzjYRrsLVk1k6MTcx1GB6xJ4bqxDMfNe5ZIJiLaQjTPXq8JbwF61JZOVsiStfk
atVL6sFK+Kk/9+OfAxbe++0eoEtlmeeU/AoxEFGFcUJpc3ot/oxrA0hVtKPb2n77
HhGAJD4fd7j6URzgm7MFtg2cUPRlBtgjI/XVSsZ65anjyXssE6AW+SSR8Xcb7Off
x3AjYoC/20ifx5Y+eNSIuYuufBC3bpDD/A3bR+3eUP8DPYXbrvX/2fkXKfJIKi1G
m+8hl0IIoTtBKCUMlz4S8FfqgAajO7S7DJKZ2vtAm3tUSiBbZJvkjH3u3g+7Wu3T
TzdQzuWAzrFn/7BCdrpOqIGOBKIFhnTtb+uOANgElNA9c7pMEQ10Wer6WX9FPoyU
P5JTCCnmaa4k4FYFMZ5JSRHTkGpGZydW6VLGmmapMe/JXPuUCjBIRP44sId8Ymyq
nw/fB+UULukO50zfz2dUYKrotzImGbiWIPUHOqM8syPlsIOrtAQsRpQBwWxFh6vd
j/EvUnN+0pQq+u6AgZri3vb2pJXzn918/x3OQh3I6g+p/cYFr4Sjrk0IfqIVmyyK
IzrjWPkXQEpvbZEsuT++R73cyHhT/uMy51hIDeJ3MVXzgKrC/WhZ3JaLlfXkPQS9
IqyaHI8WNWWaM1X+niyFBQH0V9ooJGps3TylV1ajibKVCnKb3PlJt8zhy4urd1w8
5By9G0OV2jotensbefeUcFc0gZq+eJUoHAB+senJQ3NUWdEDfw0PZq4HL6tyZUhT
4rVBuhzIoAokhMbzuauqbWV+bPjpBtp5uODHIbsRxr9EQQQJiQM8ErRLQl6S2Ux5
77xFGh746iYG4CrMiXDDVALsgJuZUC0yCAnSqvSkJj5sWebjN0+N2zVZvy8yEio2
m8uc27bcdWlMxW5cR5XXKhAT2XdVrgcYZa9Ib04rqR1vuZsw1//nOTJo/qWNN0JN
2BzL/bFqd5uOj9g/UD3dlaICwygItmP7z3YFZUxjioUbEso1aNIZGRVf/VhQiASD
vVdAa2FP8hPJeRaJ48/0jPGr3igSYze5ibbwJ6PDM9cq8x0JwPzM4f2VwDRejR3M
iiXXGzV8Buhth0sKajvfGXH69A1EKSPkzS+GQwMw8JpvoDz3hVocafSCFAmwiqXa
Mrxws047teSvGNr7/vvmEo9bf6cyoID7RYMPF48OXypB3UuePKClq2GNMUy6LP/X
jtozFQTnMhzMByluRo8YNzHzX5CgsGHTKd5nAZNJ9JHduNoIpBP9FuEQqURAGhnd
tJDnpYETv3Nr50LEU5uglrv9pr93OpvMx9Lnl2N225YHgiyrsf/YFC/3gsAJTTy4
b+2Jnx49sBd9oadC131XimASK3RMMI9qUvIsRTAVR4xkWDX26bY2ZreXQOO6pP8x
yJq46388Ce9pAd86ASX9b6QmkrTsrtRFSMcBPsyXOwHjMLo0NlpX9UDb5aDFakMs
lnnxJbizSsWhWt5tzn8EFfAxBHHR0E5Krk//aqnAtDzABE3LREiIbacqm4F98Sqr
NWb4RuUHZsIhdr0Z1eFOVjTfAl2nEMm6qgIDeoSAv1sxv2NwHTLc7AB5IHheEyqX
eF8Uv7m6zqDcWqBvRGmFoyd1XFwb8Gq8PAQa6EPHrIXzW/nU/TrAxXJDrIKJxfUA
//Vx59oWk9evaeieoGyF6tDoDp8DLGD6uEOR7q1iw4hmZG/SDX4Q8iPPhjn4v5GW
WFmEIah2AbRRXtleEGRPINjjaAgjbeIFdsE0W7atEqXBJusw3p4GK8LhU02SiuOJ
HEFtkGj9j40yahfc5F5HH/KsgtQttkRDeye0h21XKWZh+LbiTdV9zaaLFpXunWic
P3UqMEZEtXt601yw3VMhw6Cd/krTzJwC278fOOQb9borkt0gygLnn0pUHP/7Lclt
UIe3dMjBIoXbYvnQAjZUp9wF/EK+gyFybhzAQtC9e35MeXQbRbTmV1erHIYAENzI
9nQobgZy3ZKf1/sKGwPu2AGCfqE+3SkF+uPDJ/ogaSodKDa+vC3fRI2abT4ZXdhc
zp/Ol2pHx7/E4LqO4/EjKkAyqlgUWNiihxIGxK3yY/5gLgr5T4mDgbOoS8X/tv7h
APclQgrLtMstC6+dKmYKQnlZjMcwThiXDRTfRtn3i8uyQyC5WleoE1Nz5VRb9v4N
i7EYksZycO7GPGKSrjeLEEaCDjVNGUsKJ0CPY7HhGNC1WFe59RIBb8oRjp0fOPsJ
tEkn2qCivuoZUMmaU0ELlEubIXd5WhLLBW68RlrajpFm/l+0lym95vrluEIkiLkw
NqpmbnMnWjBmmor5NKhQwO+zXPk/CH25RC93K5YLFzQfIcfzExzWivSTJ+aH1AtN
WkZJepUR1mXFCCYwh6MI6iGh2TjYFwzWElEXxZbHqCTDFAWBjhiw3iyLwSSCOiYz
k6JZRs3GFcGZEp5/q6EMEt9Hw8G/Cewncfsuz4fsWUsd57EAMXAJT9pMdBUyg28z
hvZ2AEI43NnhbUZ8+fFSQmMVGKRWjyhB89VfaJVE5xucdkAp1kSmwGklCp1tHzO2
QlBp9szolOTz5dv6+KG2ZptVzOmALef7nN2qWloY8YMvYjhDNZ6M45A4a+yqcYXH
qJv0xhJMVnJBj5ApClt3eXRv9TMm/QgOYgo7kGnM7ZAIO19zfA/MfsOluNiK8Cjy
2ReQ8DZ27yDIlT0ZSrh5JdtkDwzQKgUZElP/2AygzTlaun66gG39rT2lune3flO1
lDe/VZnzmsSZPx542f9QIuTR/D/9XcPn+PgCS+96NduAzSIblmORsm9Wc+FTGM+2
Wo9B8n+MQVfzbQrf2GyRKNkk6/NyZMOjdsoTTwtylBIf303/5U69A/alGHl/UnPv
B3X1P29PrXGLPy+oUsT+9yQwxQ/MyaA0+NdBEGq8N5fnvWobOKSWkmPC32ox4yjG
tEqmL/OZjXKCOHrER4NUSSMMl+Z/sp54OKRk8rexZnY+/C0svOtgzbid1YvfELvV
IF4dpeq4eZMtI28A6vcHW0SMCni/J/IL4xExHe+Ss22COGtshaBhIj9l74n8AyZi
ia6guTrBp4ailFr01va6fDmciG1qto2scRd0TQTtKZKnySIKnJAx01x96hcYB4ng
AvCDs4bXBUrg+jaXvMTriydQrfcDaaPqH/vUy0cwh+NwwZPA5eJG0ecz17OWqh4G
trDQLLvZczSptEKWc+LW5kmW12dHZtP1Hb18dwQ99KK9RebsqwWTB9MrY+F8UCzd
clvbkDuckcpMhvwbxBTCfcr/oj8pqRqmHT5KXiC25QvugyIRTPxeCEtZetmGQikI
XhLZloYIzcQKM+RT++Atu5TQ0KWEbRZkuuidEA4+1ZcqBBB0ApdNhwDGdOdbAGr0
wLr9im+bBuhjQkHjQU1EFoWAHTImA3ccmmDQM/tDZrmtonidiobZIPgq8reLeMEJ
hBMlZS4Rg+drpTG0B3+QZUYIxZ71ZwmFtWU/AAjGbJNjwVVi8kugifWw3xnNZzQa
TyKaVixpjk5NQojvbS/Dk7AgbHK3zp9PpMpd4a9fPgbzsYc2SSbDHit/Yax4U2rE
GG1CCrtxM0IVBLeJzlX8Ms45qhGhox89rybqlrfDN9MO+prC8x1P71FUfLSL92FP
+MTyZSeDLBhx8Ym8Rtzf1dgFZxXT68UrmqIXiPdGUfyVFgUv/K4oRdnG32z/3ydm
eZSlDNkXtBGg1dMLVRar3v7ruH1oDQAQIxuSa4s6SNXubegj8T6UcnV7bk9fTOee
9EPD27wH7Yf+9FJh4te01OslCTzrxgaDDBFJoTdPjKOlTUwi/ekkr9aBy2ihb/PH
VAnScS57SFNybbPVaeuKhr8KY4q7sC+X3BXJNACS5uC/f96zqdK2ThnpxPq/dcOt
DDVowXqUNPsJr/k59/wC3/XFPF9CbGDJ9gZfRXcKwpBhgN4Y6eZ7O1MtEdz1wT3j
YamDeIHDHHDXg22NLA/OVRnPahcSBdZd/2oiCrncRadQMbeqDnzSBFN/fiXLTWGI
gUZoO1k6BgQyLao8SPuDGP535JMEVUvJ0L6tR7KO0YdafCo7Ja/UnLQwVuRiYHeH
kPj4a7MICduF3d+L8iSogNWr+ixUA0nKSOQgivIeqWc7Cjrw5UdpJzmT1OAYKW3X
I3pHWY6vnfJP4GMg3UVJ9m65M2GzAekY5e84102nLQTZJP5mkzhLmnEFfOROJ1gI
1c65Lta6VhL9YJ5ivPI+l8nRINPeSe51v49QK30ZSGnySWrQEbApfM7WonEA8Ps+
yWqmvn2eHvzSQJoRg8KpuKzC+Y6tHOxbn4bst4FS2gB+4Of1XEIbLvugc85ZnUep
hSD9XIvoPPltoqLvI+9EjtDAUT2M17WX8kXHqIy1lPei8iZ8J4Azi3pPzAAlCQnc
iW8VqnUQbePhnqOjSnEDXBnK+eo2VfjYJedzIJBzqf11MA5/WBcpmC9Mv1QrP7oa
WXXWjfC1G+3oWwRJPxT2qocsTbaMvuWNksBCeURjsUaF9AYgD7z6JamWCvvE/lOw
f4XtmQ8bk+Sqde4tSTE7Kcz5z2I/5mCelro5bIzSMN0vbLc2EY0ZZZyy6gfjGroR
qx4ny/ZmGZgNNXbDKt2rk+VU14ikLBBoMP6LlrsA+00KlZwc8qCLQGPUju0zRZRF
wDpJHJUROjlzIoqs9d3qqmv97TIYOhnCf277VtScIUB1n2C07Io/MNNuHrkbyJvG
d+bysL3ysvfVgfYg05HRZcCE0PGhlZOpvZb/YYQcFCZWyPrxTAkGGAuYHeb1gRwF
pJhj4d+lJypt0Q24qMmrJvBn5FpYy/q8Z+4rL/c5GAXVC1y884GpBSE2/8N0eyWS
E5ZdxKc9trGBbXvp+Hfrr7HZIk6AINzxw9N6uRRQaJNKZkCRL6Qpo0uXDuPjclVf
ZTUACalePgp61+eUm/ab6ffQQN2167ASeIT9c7kBZuvrLWI8r3ahJYLApsCK92ez
c64GwPPyH9TA585l/dZfwfiB/0OLakIquq4UhpE8AVV1PwrwfPkXqBpflCLK3NfR
QDWZEpPFY1/l2M7v2OtJVguSFH6EgmP97AUZUbVhDVeJ4faaPWQY8/x5WGIiKu39
gTc9b8dPS3U+rd/XXCMl2+hX7SkChmx5gjSVm1ocFE29dQ3Hy6UGUAwbwQfYHwzR
nrlEby7eQ8G00jcAQlsNaV6d9g4sSSUWd8E+rfjf0S1+DdHkI39KYfjP130c+BsU
s01G/DDd40n1kaMCXKSLHc2BzeQ+vhW7pICEYbq1n0Xw88a+hSGmq6S0yDGo6I2S
yD0g/nCSeosG6p9XHpTfw/QXkvnrvrWOEOfp/jseCN3Jt/ZDaKa8iBAjS+Xvt6mu
v+dji3s2qNoXrpR/mJkYXjcYC9OdQXf7MYYgFkVROKlpPAyN7bN2WeoLvC3umTu0
uFVbDw+uLC4EvxW/eKm9TH2pScX/PQk/m1Hf2bzOf3uzh5LQ86Op52ghqDeU5SfD
rprrGcCdAz+zCwY+gHJ6SrNoDribQpJSlTcBR4fM0Ub51tawefZ1FKWawFRplxVf
rEYu4dBvXJzrdC4DH6CtCQKjUQFEybCb9s2de8k7JcFaXvCXQYyQKAHaqqEgMIfq
k0QXStGeyf1qALZ8A2am2pO2yWImO4c4CRDK2tZOI9x5lyjsB/9YZlkjuXzWAXXa
LLsnUuQ/9z1Z66CKHEY9bDmNt/xdG7dvHMU+lJeI26HSd9yaqKK/BIY8RniBrbRG
mQ8lqzFp27nYxeMCIy1BUOlQI+ldGolJSY2vQSrl62WtAfTfdbwbnDx23TFA0CW5
/mE/1wAYa5Gm06pTVtXxVQ3RuXkwy9Ksh3Mou2P9/I24pFENe4tMlt+1npdSM/Ch
yfOmrSuDGecV2xc7CdUhCanxLmkqEX4pRWqpmqwN2gj8Y7YyV/zFBIZUkF1OVn6B
i2QvbjBYd1JvcUrtQ8BRE7XISmCX/wJio3GolDhh9fNNeuBY0vSFeu3y/qXkBCr9
1QdYoxEoRiQ37EQbRG19XvKz+WqxvJewObyAE96xHqNWZuJNAfR0die4sBKBXdM9
F1lDOT9P3vU8UWjlNht99QNyghmiA3sJ3R8Yvf+dzFMOhu4bV9h5+E2HJ39wMCgN
/6y5ym65HpqIdxLcbHqyeqOc0t+GoN/OY1/nsqiME8xxHI9AlLLeVi4DW0LfGTpC
rdkijqHiWiaXvbYt+G1eAkiHTT3oko+s/B4GujnDqlT1Vmj3Vg+TJzBGNG6ZmS0F
REPSrkv2rlopji7PKVSRHTnfnolEPyRTX9y2t9XnnLyX4j2X94aJFJKtWfmr2aQA
1NyI2fzv3Pq4VuCyvqx/0yIKB5znngQGsBVJ0mXP5QsFw1kuNkL86e0h1K/WW7Xd
/E8q2iCyZWI7QeUqVnygqNO4v2sNpG/mP3pyi9VWbZbOHgc3ZmtsiYXiCZhD/zEp
MINntCW2h0zMT+5GDBmMwjGVNmZP0LEialTiAh0EivLFOZjdizdXDtesr8zCZG+q
BaZAgXWGT48+JG97mSvcZvpAlmvP0ONN2ntyz4GtnaBrfLozc6KEibUuxsmxeOaN
wFd2qW3/S26uJEKO+1+IfhNHMZWxVxZPpByH6li9uu2UBEvCs2cGkVFARq57hPVx
JU2hHxSg/HYEnrHBhKHhs2fvkcjIYr9dVC+xrnvHZmhdX6chG63DE00csSG97r86
QxVw+tZWW971AUNVaRAO1c8pBraNFhA3aVg2cGYRp+dRHgKjINH2rgA2Ap401Ets
y6cg3dSDs7qqXllUXLUzzhXkLYUkuU4K1IuF8m1I/u/hT9UEskfMeu5moTRlz2ft
lN7toNODfcSSEigm7uKK5o/x0BBBHUN4ysq9BTUsdjiZ19DTxtjSVco/x29sIAuo
U5NnFv7U9ipgDxDfd4bbfdME3cpZ9GzLxe15EfwepGHImMYtcNW+LuLWqnVIZpZz
lXRHWAOYEveyT8kRfuJQoo5LlXmLXDB2UNPbFLvVuLryEK9ObHCyV/pPC7qzSk6x
WEW/gT8iCiYSJzehzL7IgKkTo6KKjeQ7Xd2PTAn4T691mi4VxS6Q11zX3RcMplG6
87xG83HeEcLyMC5ApnA4+EnDDi8iBvG1ppVzxdeMRqD5mn7QAwtwINJ0F4grtj6p
s3suGYyeEsiLtAxfUEM4rbW52EzP8BpjezPI1xTHPFvR9MMFrLe2XjnjptgS/6ZH
YDvg9JB+05lhmerMaXhxyLiEu45OEQI1NdoZkuiERixY9xYnglQG21tEjCWMl2+E
/HCxAUToXr/DylrxfzwlIYnL+qyqLTQ0WU+Uj5bzlUsdPfHJCVk2naA3OTrCOALw
jtjLRNd6Ioha2lMFOqLaR+N/lo12uYLeDZLcT2CKsRIx0lGtXP8z97anCBBfLwzu
EmOYaEOaQleejahrL/VhQyCPYA6S+nmROEvCRQcSRD2Al0n2qQ3qPE+mJhzLPZ9B
INuHS9Nq7ktARmOBv8fcSyR93U9LMSR+omRbvPrAtiXXs2C2PymYOlnYogDjyJWa
tFEeif/n805VJHvP/aUT4/pdmPQO6aQnhOAsF2fZ/DDtVdRphOsaCD8ZjCU663vO
TGpYXifRdB7rv82PMCzzLmDmb607GyuWWvtitP5nnwQ3LIF2689wrxoiXuQiOFHm
9EcQ5+BW5fGxapdNdmLtlC2P1NRX1wdaZXDy6IY5IdhdeUeIZeuqJZkVocCJtq1O
nVdcVMT2t5rRn9VOn2JcXoAp57L2DolFRjMG10T1CTytqi/96iMgGFXTci9zNBAE
DoVRh9JSnWsfP+GMn4oGcR4fqYwqT34CuToBAiW0Ae+2lC2aDinpT3X1qJob8B+r
z4zGIZdEKHZT83ZWPKZOHhVPR4HxiP/jC0lY13FkG0y8V55WkkGKK/G141jqUhsa
EbPu/GHuCdEQ6xTtj+PNBl7GK0Fiz2WKk3GJumO2i8BORKCooQXpuA0ANkKKvJQZ
2zIS4oU4t2mTRjcuDq0iCQmOiCOK6ffQ97pVbfXmJC5DgQSM8YSf1MumMVZur1Wt
LcHt0bU84Dz4plD+SXJ/CC4JHb1y8zE3uceVNUN49ZM7Uqo7l8A2B9GyKHnYGSvp
6OiD76yk4HlHgeiztc7XFDP/2qf2janAayibgQFVuv5xxeQNNvuRsBumlYemAikc
G5EGXcrVpjctZQkPzRc3Y+FkyAJJdVrfoM55m6P6gVxnIuNoUG1MrfNzenuV7XFU
OmHdfYifMLqkomwlcay4h4i+UgyQMYx3aSHNNvXIJY4hYVpIGBuO9QYSrhMDp4l/
7bv+dij4Pbl1cDEaaPaXqHtY8qPhSOouH+dhJ65BoEy4UPR7C3lCggH0HvDrzrLt
Maz13vexcnCRDPXu2itZz9jz8rml0cvAcjcDN3GjnKAetQ73Eld+vRKyI8D4lWMc
M2lgq89+Ngf0PNGI41wCpy+g0V8+kOFVfkUEcZNs1/X2zVhsGrNwOjHdQnaxC58j
NgplgBE17dqhs6EplDEOdyAe/QLB1z3g7YMAkStYx+O5gMIhiWq36/CtXqypiJtP
HZKpIGdaacJ5tVflWK9sqquqXAE26IGEODWo1HRLsDwZOl0Gfj2U9Lzk5O5g7NSb
307aIhK2YdzC9n7WHKfmXq3Y8aJ7qL9eX7R/LfpVIisDh2Lfasc/ThVdb7ytx1nQ
7AMSHsx3JRn+dHEwXg3yy6qAaFbbM1uCoFMK1FXDhhJnpsIvhbxyJ2lfNn5kobAo
cUeHxFmpHAtekvqbT+aTtlCi3kQ4zVWbKm3iL2r79TJm17P+6tv/+UEV24pIpDTw
lmB33ObE9LQ7K8dVz6m6hoKDAZ8PKS4gbHWzPImb00NdGJNto9T3K7Fh0+kogTeh
uKN+dP0YZ0BgAPlBSCw5Toly9ncW3EVTYK6Y3TUIs/s+IU23Eb6QvTDwhG+5mGcY
1GLaaF8w2bEP7d17u7VS2p3+afc11cfeHwBb1Opu9CDPgcKnTBfRKxSGE+m4Csoh
mDdm7Ta3If8O0srsBIXScuQX/WPqlGz+5tPvzTW3GsaPtqqV6H635AU6pB3pk/un
aMXzq+5sGSzrS7LYJx9ibdMNDg8nQi8Mk1KMpQ4CuHMGhbLz6hu9c58rnAV2l9P9
jkLDBsxS09gDStUwoHAWnSXDMeZko52Po/dRhI8nZzaq2Bf7WmLdafritbdRdNNP
XiRC36cb7WBkVotgLw+2wyrdzNm4xjPYowE3u47BrTk+hH2ZaWSI7iolXzNza8iJ
YdkuqVCfUjzEV3cbSjmPZvv3XxhCoA8ROIEvneYuos6RKU8LaRdp/poM18/Krnxk
pGo0i8Aqhw0eFfoJtnCnoYR3FgcChcEWPR3xXzC+s/wnXqxiEee9v6UwFhVScl5N
MqkN0BQw3/8Q8N81XQ6G6uYyl82HYC/GsIBnch+qndT/yrSOXuFoczLKsXAQ6zuB
ANphnJGKzhy4QfMyoTkLCcWDIL3/R3/t9xNM6clPhV29zpVxtZZCknG02twIxbXV
k4Mlb+WrIot0O/5Jknbxu4P3YgniXTfZVN5ZAjKvuYial7tHUaipiw3A+IQ2bZ81
zfZoRqr6aGsEVUA44BCvVKBOl6TAEVYJtb3TH2B/SsvCHcbFOlMHtZ0Q7pMzzs9o
PM1uUlQbbGN/ptO9prruzx4EcmKQJQTOE2OBrMwwiaEsQWPQ4Qhzm2pOmEUGDKMd
Xxwe7yl1MT3gdVRndIYRoylsv6g0AzlAcyGvcftT3TA7KlB0oWShKBt4Kh0R/DGF
Uxe9hXL0tziZvK3pH0Vr2rUdWYRsZxfK7B7ZAHyj+UQZ/j6fTJDR3YAzM0s3tfWI
lc8GFFDHic6ERyfchZMBbW1weuX5fnPmpkwJf0ZDa8OSTggg2zrjcR4O+7FBDXKH
6r+8Veb1FQwNdNMIsqUZtcMHzPYMHhAhLgqV2gfv+ieVALOF2TdbSgkiuiX0X3fX
dm3siyi2KzGwpmnznBcuhE46VS43UQDJxU/k6++6hZ8DdgcWbpxzJT8xfnSVE59y
zwPvpHqPTEQIiZlayF7Lt2yXp20x5cSST/TqzvXvJJ29tJWH9MRNqDNv3UrWI/tC
Pd2KWrv7MtrBXt4QsTlRphF8ObpqJnZr6I8n0zoXduMjQJOOLvOz/V0HE50FpFlA
35mgSccM5feR0+PV/WB172QDf/DDEFvN4GNH4pclhLnJftvp5T1DjjWZudLBvijb
AJkWdZh/ichcOjLrrCLNakjo7lXkUykjFcG4DZcG57u+2jAQWuEInCZ+TthN+8EF
YoKgGSNd6fxC+VKVlx6AzgUK3EB0MYOi5vq4UOjb58ZLJddSmpZLW0npQ5FzV2cX
H0FWBqEHtAswSDDF7K40yLQ0IVAXVeYK/DGRTu8BpvJpRv3r+Np2J7BXlNQGjrby
Yvk/l8IsN+GIacZnfbzm2EYQcRnt5qsGJnNj6Kgf4fJC/4dHo5xurLLzXaK7YyKi
iKm6RRtrgqPHmhmonGG2JKadFx3PQLHTZlQ7W8d6KT4EzlMYfJiodTaDuxNndiEv
TD5oNVa/EDvoEkKuiXYu4s+vq+pnO37pBTV9mreAiUPsickEXy5J3Cs9sgvqMFE/
zxhsqnMFbjkHQQ60g+UK85OZNpwfAiQftVLjcN6/32fXjs7ZBBAjw0jTB3vJVRsy
DhahPoAa4z7868/tXwFGrjasmDCtQV2tTmBVpEtq7JXhGYvBEquQWLQygg4nT2xj
wrdnkqjHOvbFdwnAqjux68E2Yu/qJ8Man7Vfu1875bYOX/qpHqlq5AHnWX2+X7vc
ukxup28T7UNl0fvjWdWijz6V1uRc9QHINssk7J4GXFs3acC0dnN7YgjBlUIbZfwV
OnxUvUGa5RPcrl1UpEvSLR3Z9RdxgXnhaV8XWQzPBLdSMcSJ8tAooX5OjEvwbm6w
KX/fRr+QO8/LzUpdZELoDhK/B9JIEXIWR8WERvy8UOho453wDuuEMkWtH06QnHiW
D+Aq7/JcmM3/4YPQy/trnkVeDNvs8PP0/9BoGKTtmsgciWEOAASpfuZ/TN7ymdIi
GS9K1OEYEWZ7IvkmgnDWwVFhpNTAMpasVvWXPJaLCx87FAGcup4ovI3UfNXosIcV
UHhCBM3OHdvs37ayt1MotVuH0dJ+z/86TB8SC5/J92uncjNsG+k9G3MubU35YRK+
x2JNPTBPwAxwOlDaZqnCtE1OWOhqG6Cf/OFcqlAEil4ONmmaiYTv93YcYWL1kUgV
CLq/KvudX+Uf72gkxIvJw8h0YEfq++7g11BKiwP2oo518oacXbHI5iP4+uGY9Oce
0RZ2CUX2Pf/NJkHhZv68nnqtibXHZmvqGNBpd7seRFMHWFa6zAzl0K9sjyWXbqsf
8AEPBBtrcs77ck+GgCU1ZQaR/i0mjsVJizrVqOtzO0SguZ484+DXdalIKniKkw2B
m4v3D6zZ3hvizO0uCVrvMTLP07ZewGuaBlP6ZktyeCCzmQibzo/hLqb4ck/VZN6l
Irueo1j393tE0NIu6erOAgilDnhczATpxOJvH41fNFp9JayD9Oup2U9Ie/HY0odn
+M4oeamATkmTemPFXIfXT7utMl86zfZhFxjs40yR/tlO4vWqNmy1Bt1GWPusZ9uF
RrZcRIUbXO/gVoMEIXKzKUrmrQHzsJKUEeSKLbNwMExVFHHiBOiL0tKBbpaN1kci
7BFfgq0V6f+3aaGP2h/IBBObvb7BAjNG6AFGT7lgGfnNk1IbPIuVeLkAIFQCHal6
/dr2W6aAPxq1gW3Q3SWzhRN4vTVSqCbCMbol/63pRbwS2LaxTJx/Or2QBUg4XET7
+PdLDw0mkaK8EhhegMfzO6cpdg8Kokyg+vQiyecIxQs8tfthhtPCXdF/gt4ECvKH
5zKIjaG9SjZyb2XuwuXiT1sfcHggx8ZDRo/FrFPmoCJ/7YhSvqD/p0N+X4zNYLFG
PsSJsFfKM8XmwBTIRfGwZHzoEhRBCfg/lUrOx2woHHsVWei94cImWUSZRVQCIt1e
vYX9oOy3d+S5eqS94BjQCZSUB5wXIf/R7HqDdlkNHx0yPGyqoZQiK4WdUxOH8F5/
IFhJF8/EDfGtemtmFK+kqWAYYYnanuwZbdA75r/jaPo3PT6q64uZpR33ZWwKa7W4
PBDAQFdrfPglOzoTHDHwhjNJQhJMELHbEXWbfK3Xp3XiVbPoq/L/gGJ4lDUbg7+I
vuQZxPkiE8CUUBE/SJi0R0sEzN/hti8UAN1Yw3Q4nMMNm321G9PiMu/8GbY4P6h4
wIpBjPvzv8EwSu8FQJbp3zs+BrbmrhpwNLY7T5cYHcZ7ZD+aqCmbsq5ZLAAyi7Hl
GC5yL1979neHfy2hizS3A5iUgukQaNpOepZHR9HJATn3ztcQFt10LaNH4Kf97h2W
eSyPjHvI/dyz0k/jo4XBf5/uMpIMzwKSf3Xl/Xkvqd5/2VRQNWelJePj1K4Ev9cX
js9j9fiFbZdee7xLenun9Ki/X2FQRH2J2fgwnMQbyKvixevHb+BxRuH4qP+g3uBN
4xnACM+bsXH4xbqPqjVZyb8RXBauoX4sYhbhVvlvVZg7WIN+CiaySm0RR6vRgnG2
mVFfwmVeia/Qje1eLUbr5apmnHPKDnqniexKbihvOj3Lf0hV70XLc4OeIge7Z3zr
imogjDOQzAN9spxzIDfxUWV0OSdv8bPqfr5t4VlzWVDlk7a9j/HtpYd4A3TrO6zT
7NBxUJIzhNcBeIpDZiKNPyWGXANI6tW2XhCGjPuiQemNaftIgigVWCENDnQ3eVOF
WWWpXwbKk5Z++KffWJgP3OlAv6D8Gbd/xqhou2Iwl6d0CtVFNNlDeDDqML8ilcuR
EypnbI8yhhW9mb7p8hyDh07XmtC+gtZg93mRqrQF6L+cAXuValpSimilpIi0YLk/
4HnOqawgxjXKjtM2L9wMiZod9UBctKcPLm5aIpXmE/KzdVcRDAVxGOPy4tFGLZk1
QQPOTvbuJGWyZQP4LuPk2ghk3kMsgLDcJ/8fV/muPX8OnM27mMd4CykorLi/euBX
ye1d4a2oxi9gwWFT5q+mOPwg/IsnlXJy/f9C7+babcKvne4g/k8dNJid2AumnnfF
EyZtqW/U2yC8DPmsMoKso0cb5Bmw1B/lbBZ+zZQefahtbgj4S0Dd709p7wpSHl+F
MsaglD0cUq69EjMgcACeupXx8Q5my1opFQbk8BmCaTU12c+oiKrNbUE9ZAOdlNSI
18w1izHGr89UeS1Gl7e5ojTaN9W6vdOUxGyjv+epH8KLy0OjbGxf5HX5KbnV8LjW
M0GCObTKScEZhe7xRgvNTcI7I239MWP6fjdp2B3+D9IRY72xUEZ2LNXfpOrXxAbk
vkY0SNTAsR8G4T8Hf02bHLVkHHkuQIVcQkjgv0z627zXOUYioW3781zMmrECJes+
Ag219hmOulgp5vrCra9PJifVVULNvcQxGw4kxAD7roPDeLm6GR33I0XIiJ+0LJSK
8xyI1oaZS5mEdGwPz4OeHANS2r3edJb43T6mERmuQ0NUGICefEDs8fOV0ZBS/KzV
Udw5PFpI1TYH1vgbwuKkdQJNmAtP3oR5IDka2V6jZOaaOUt5ekcRNU6mOUGeusSD
vtepUE+QnZfqLB0DPjYysQ64604MOdBcZ1sFF9MMY/mtaoHSF2VSqns8wA27eV1K
nXQHUsAG8g8VPQc0zOrhimf1ilxQ2PM+SonPCocX3ar9M/bnSsytnrBDT4h5u1Qa
25LBk0wfHdpj0LlZMuWb5J6pObVjAL5/gBW1kpK09agFA83EkP4ACTcBCmtacqwn
ZXI6b2j0guAtfqpvMoLUxXtg/7mBcm+vRnDv/me1X85G5gXXW15s5uU8RKCMYmNz
N7pJ0lk5yf+LmPgZVnZU524LCCdbiOCD456ypGn1M9xSpORns0AxSkCCJUzi9obA
2CIE1kTwLOx7KnFD/K5p4YecAl0TEEX1kz6wzRk9znJQdHvKVRd236bFtZ8juF9H
VbkKI3HniW50GzksBSJJ56ZMnir1Xjeu4I4/oSDHNxgZqC1ST2sq8KZpgsaa96J2
aN0uHCi5STRcn1zZQot3JURlmt6WPBq4mmsbxWCWuZKqeFzQWm8PYyY/R/E3kiHB
MPv1OO5syxUkpUFLs0YqNR9K1hveuw9xEPg7CiZW6uhxJDTYdbqJx3RYPNZntYCJ
ztkQsuv8zag9AdRUxROnb3HF/mbhNsTsLPX+6cqM3EnJP9JtjSO8iPkLhQ1Y4dPa
QkSf8a5Nrh+cBI0ECypI+skZBjOvqS8p5vdlxRN9v5XxMgZqX7avPbjes3BK8IBN
c7KOpbDXgCsBqk88DQQm3BrWjcb9kXVg7UACoK7TjEgXNo3GvsEbkZXZ4j8WpxzH
XLCz7SZt38SJSxc8YnkwPhiAcMLx795GWXWtXBU4J0x9YEx4ed6b3wPVWhJgOTwo
C6+3t7NUAk5sEKTTeF1QG3VomMGsYCMe69GRI25nhqujsHk3Qlael2Dg3tCvIJCH
Mc4OGJwWWfpEBfZcLruy/yo6rpcr7TLBw+2R86OYQ2OZ8rDmeXmSW7HeED4+/1eZ
MoBnCb4IPrbfsxoIXbGRxxjFDvIXeHV3WNSuMk5t+eAttxXW8IsmVCwrWYisd7+a
O2wM3TcE2whVI0idiOMlus64+Yhxmny19JuciCLG+CyXisrA1nGaursTfpU9qzjf
n88kBeC6T5PRvz/hK98wTsfCLMgnT1Wb25rNhCQaqmb7DKc5nrBNDlWK4sXiK2hD
ZSir4mzFUzuji024RQuZ7Ff6wTs6ob6nS+cCksgNTosEMu+2RQur3LODo5hIytju
fTt9U/wiSltf/GEFSDZWkqTThcpq9PKOIFdxt9w1OXQeHJ9zBpOgLga7HbFMRB18
EVTMVZKzW08mXsMa/061DYhRPhXCYc0lT+Xd00t3kS6YUuLdg0T3NHwgaWm7rvEI
O5f4DNrtNqHwPGynmzPkXJhGzGCzfr9YMfHHsicda3Z34Shs+2QpSGyhe+Nc+d+k
vIAeltaNtYjTrnyXhyLr04cPKKGZMqrGJdY49LJafbritiYIbghhDwQ62q0NOp+B
vuRtmlSFklG45mueB6YHdzYROOWkLrejCT/cHirVJAE/IttaUA8euiPNM7wdhTsd
bKElrcY690ipHMQ3YaBJJ97T/H27+Krd0W7MWDF9uYhKe2bQKPgP3r7fAYIXFwjo
bTR54JGcilTP0A/kEdhunMk9qjZZkkGXDsLRpJVUYyRbiMQHhGXwJVlsGn05KNsP
pEk77Hr6Kq4hfHmhfmElk5yQPRhE70D8ERXnTVL/XtjSSTtXxwHxL9/hoIKbyN/6
oIXFhh2FEqp3r7HOGTIbZWVEEiK7p7XivAdRlEnvanNEOzDj15k5Cntn4jFJxWB/
6wJFRRi5u/sXFOVnIbPcpwqDQ5kTotuYIjz0/77BV3CBkm+gw/eD1MsAEhGwvtEu
SINN9TTE0cAOPnsPKda53mA8bF/JjOrO7Vi/pLNrdxpF8ce5I6uTASMyFeDyrPe3
2xQzVzpDTRLf9UpK/djC9O/+eE+HWmJVJbSNhZkfw16DR0U8Vw1acKYjwD2KHFnm
kLaw5pWGDs7qPeYGJGVKJEnQkU2eQrMS5Wa+MA4KKm+rk8UIdeNsXxF2Knj7LnJc
luje19l/7hX/0QWtnCIV4/1IzT6kEWMNXJNDyPyPIj8uGbmomxhHTjukOrC1mTil
stcXj+bTaAvKNCib4zqBqZWDjzCpkL/b+k7LZhdQx430sxvOy02EtGf52hMmkMPo
48ZP+mZw9FxnuEmg8twa5Epj+4MZPF6xDmBKVFLdyOAgxMRrXJMXBQIkTPyCQePC
MznP9Jk10l+s2NLGi2LK42u1DM7KWGzlXncMbClifu9HOZMco7gDZREOmNudOL6o
+itNWfx86HzlLfoPqmDt3T3LlNokl7xQb6jbEwO89U8HuIAmvDEhR/Xv80s7dUua
/76lx8OvhrPs6jwjJfXrQaPPU43KgkhLR2zvJpzCG8WNsiWS6J33G46rUp02FDh1
ovUSVNpj3ZUs1WogmGkz1BBDtsp3crrecr/tGUbZALoF7SBqhpoDODhrhoeygXUV
edumdHvJ8Vn8tCsop4WYoY/NqhL1NBXMbqth0yvJmY4hub4/GDHqzSxHFf7Ci0YI
vf0s+ipdgLWKzCI+GA+tbxfuYV8o9b388qYTK1rRjdI2TmLXqf++NHgARhFF3dod
JYJD7t+21TeW0GK4qp2iD5IR6neVktlIu2/wXNqbLHn/lfyDR/rn9NrPaYD4GpU7
oli7wSSvytQGNa0S2TctaYm2bK7QD1N6COPHFe0dLUdjG3HaY0XTUMyNcikFRPnX
inOWMSnZKrW5e8zblFRSEHhzjeppphp2z7omxCfVdvGIqz0497NSILUjUXhCSuba
cu0FidgNjYEfxksdwH4/KvKrUOUKBZej24eN65zSq156A+AagD1MztGjxF7KnZ0Z
Zt4dft9UP+TvM013BLPa8C54Ihig5eNo7KcE9S3emEEh0z4rrNVoI5M2BUzBNP6g
47VJQhVdA1codCuEXXNqA+iOKQglV0uAfZShQe8UcvDv0+A9VQ/FWP3PWusAFXZK
w8KPQ3xcjcqfFac85WXFIBiW25vGhcGHaByIphKgg8lRlrgSOYMfvokfyBRr9EWM
eeoCai1UCr9CYzaJq/YYwJJoA4Mxdmzh2dtEsr6tNrswgpLZ4ks65Y8M5TUl3hM9
O/LxjmHOj90JMwU38Uzl3xHnxwp0yPqKZhsHDpkAqgE0mt0kDaWK23ekIn8XqGvU
E5jxvjieXoVWDsHecjB3rAROP7HehS9taC1FT0rmjy7nuXmq1Hg49uVgTzv87cf9
3cFHZu6OLQd0Np0Fd10rL/P2IlD8bKMQPe5glzX5UeHXGaZMu8QDqjHGUbZBMAiv
aD0sNBP2qGnCl/N8pQsffqLlaPtKNE64UNkDrU0t0Z63Kbn7+ddGGHzCRObikYvS
9Eb2Eagk53QRMlE6L6MHFoD+H9Z0b3KawvWEqTV9irC3YBgICscozdOkLfzl/Hyn
cl969lP3J5t4T7ZELt9vMgSYFU7Ji82w78aHL9Pb7hdZKaj1nAyYLNs0mRUl/Bln
vqUkEVZqYAvt7o1Veax0R1NLofgqt1/BE9sz/JetZxvBXpJ/Sg41HcZcSm1TUCdl
ieyqUpF0dnRSOQOJ6qha1g5lscEb7H3Uz2ef+tBLiyWdMfMr9uYwBL6klRtVGSzj
i408MWipdYvF6dmU5XdSspvw7SMLnUEFqiuBJmdWAYRma0+N6yhSkXafqgS7NLWi
hTGdWn406KLgwH8Na9qyl21xWiSf7jVdSHqTcKnPqq9B2ov0peryrqz9CFp/tKwa
CiKup3WFM7O6gmiGRdBkEXVe7fHrie9M2fSLqRlDiP0V+fdVE9Ir39b39pru9Yde
KEVOygzBZE4crOlLPIt+L3FufJM9rtDXobxQzmlokiBciV0CnlcayRfj0be+BfBQ
bSVXzi9ZGcS5dVaIfsJqHDijXfE54ibgJ+8ekzVAg7aGtieHwid4UBjzVTuD08Ly
8PdkVdcYYqszX6W9sgPjbgJCLuU9jYPp42zXBVatRtVnyRU0CQORu+AosuPbRKww
S7xdFKjByeERCHkFVTkRDmNkUak3LxfP2Tr7FORdMWlqkOvxJnsnK+0k8XQwqOh9
wPqXrDshOaBswW2OeRAmu+mI+YQpFEtOBc6eb2UxLMEcgTYWAPS8q6zx8YmS3kOU
El6EwDmk8arblE+wb1fJPcTS+bFLtX3Svl0m5HimoDck5AvHM374eFBGIAseWI/q
Tqj6YmmQNxb/yLSMIBBeC3aVyeEoRxh/jVPhGIVQO2CN1i2fbjLlh+XuEtzpBvYa
0K0GtlVPoG3Fgrp9dtpbJ+ymwZkZu1Ze4+g/rkUUBPrKcU69WhIfHWUFGGdjHAxh
LyvHdMVi1idxWfAJBVI+hly1ks4JZQM3LmeT8l/wMWrs+EVV8qTT18Bx1UjeiCCm
uKj89WT+Xs2dp1RKVhD5hmuYmsaI1cEbqe0tIfOkZIyO3WOsoNN/+sy4MNhZkpNI
haSz7f+wHKHhDUP6sanGYobTp6GUaMkM9vj/5c6p4dUm3f4NAa4cE/vaR4LVCVFH
wZnvpXFmvA/1dhKfp5DcXmBUqEN9IJ+J15v09N+DQ9Y3pwuO7d5E8jdezGUYEb06
LoAdZTOV3Wu7PwQZeOyds3mtZTICZqn8RaHokfgotayfOwCzwuOjA5c/BZQ1eL+q
8w367vAJEMdrAz68e418OdEKOEMCBtVbBdBDd3gqyEknVjdqzul8ZLL1jKssOPI5
RiVb9oa70yawLXGE3qT/vw3ypPW2FnTHqWRvq+O1QaNtG3MgBrhTdxOAsrlpXine
BkUFVqt/YBQt7fZtBN1UAA20ai1cOt2JcGAsdZThQITLoGFt9EBgRjU3jUwnhuXs
6Mt0jCVx1xgA6U8rz8ycax9+R2Jro3ByV+1H6CXH4seK5zEu/4QQ4GiMdTfkqjFl
Pf9zoiyZ6vpzuSSRFlrlMXX3ug69wW3YHf2UfnGTWaHM1HX3J4iJvdhS+XKeSp25
d8vOtk8zsGGHeJWpMisz5bYTs7ZtqUpgCn5jbBQszF+fcAKC0B6mGMuo5N4IJev7
bXviwhUc6xrDs06UZO0TOckM0D8SynQdgNQnZi6ecv0cOZPKbnSYPXBUGdYVug9a
UxwB4rHwfkMSh4rbaJBCN5RV20AOnIVrGYo9Ip8Fame5xX5L/wcBaCxv0268HpR/
3U92L5/ZZkd8l3LC5Eh3xvUH3v8XwFIltiMa0osqOBMuzs+SU+IrkiQn+JQoxud7
TMD3cn9rF8F9rpglkTLRYX/OBuLPeHERP3nOwAxgG29iBcc4lGtAaocaFuPJMk3G
YL16IjNktDbrMR1/0JICLVdX3PkEFPdpBlkSDaMC9fNomC0s/1gCPw1ogihyohGl
l5tDdVDNHG00dm7Bk9gjVXStbVn4ezkewvuFc2K1HqAXTVfd0vrhUbj72RUDiEZW
9MofWKq9iYgw76cVd9MszTzEJEZTnhEpeRTKbU5sX5gE7dEw9OFMl+YmI/dF67T0
5uKMVCycb6BhZW976ujoFTqOZViLsU9pUYIheHQPHMIoIndzHpdDxyxT3KY88MX3
uRy5/Pw1M4HTxpDk3JIiLZ94QPnJsvzzRVhyEfDkCt1oh2T6d72olp0eJcS0Ltgq
n7SNHIc+1ec3HBr/kosHhWodA7qI4v0eUBFmPBod7gQVCO9rqhO09+ZOEBJbmaVt
n71r2nkZNsJuUUHtq0H6+BoiGn8LK620/YI+Lv+RqplhdUa1K+hlFSmY21ubgASL
gzyJAE1451viU4srRqkV5O6uAjD3Y3OTGkoVWth26v9D7XTnGJFEsi/PImxYX6Vi
wjSJh6yt1Ku9NRg6xrJUh77AFJfOaYPa0KY/8nv+LixgnSZyVUVGXO0NQQYVeDz/
j+OCtkDYS132gWdTnJxOh7XBki8OtZGf0yGNdIfImmUARIDmrHXQfv4xrFM0IzMH
cd2ORNjAE080I+c383bxsLADDW9gUesLC4wyboA2qhnb+o2V+SpMcciPtVE8/PAX
1vY0F42JbEfsLrQRlpSz1hSBPOD8rW3kVz/m1IT+m/K+EjwXCl9M3RdymTDToF+8
3Z2kXfvda94JycTWPLegpCURLo5UkE0/DT7ytl17K5Svq8le5aDfs2i6Tdmj+YOw
sH11MknaYfTHt+iJ6tXNaZRGZItY3VlMwbyC0hCSREi5Kjg972yJrJgah0pOO01V
Ypj60zmSD8xC+yZT5FivTBuEqaeamOg4hFT3ZuPvuHofakcA/Sx9jSP7t19eF+Yv
JpIK6TAWBW99ch/d2UF7+xx+WKppPWlEVvb0BBYTDBzdIGpBDPnDLgFU3/VBsGta
Wm8qRSkFY1UrNkJpEpf6QUuPSCMh1tFQ9k8ubdqJwSYwPkdBdSE1Rd7vC9/SxeU3
YdQ4o1BUVXCFJX6kn5XppGWgED31lw0t+zfy37pCnPvWz+sOEIS9OSBF5GPYQuoi
f7ipwjdrNIlNqlsViIWzvR6rCuxGU2GWqZSHsdSRzuJ/w1GtL0kBNgaGa3xq4hAW
PsjeLbHuSq+UO4hAgwt9D99ivCEE1IH2FikpAAAzAYXR8bDt/w+SrsvZ6P8XadBo
ZQBTvm3m9Bku9sF7ngk4C/PXD+S5HmmAu2UMVZFrniiThgSAfxDuI7N8DUGqT5c4
vYtTZK65rlQIW7ArkVd0Ii5xfXpJqS1HU3VJYLuSlH5cz54yPplEWHuc8DL6QoK6
8mw+sKW48Bg/7uGatI2QYy964TUGE2JT0GN27rwDuPq/8hR5cIXbVZ0/zfaRTman
38uMiFvXkVYNFyeK3NwWpGLSn3fRLCq9PydW9Nkkis07De9e0/4WRnpGMPef34hw
nuKhqkWc4LyYSlehm0mE9V9jiKzSaD0sD4OZleceGjL4JfabLU+tOwuqgLua9OUv
p9x6GioZ4vhkdQ3y6sFsM/tJ0XzNw14WHXtCaTFDsuRaI++qvr3KUiZTsiNOtaWo
7fog+pkv8ME9y4q/uU4Ezgckb5KWRh9jyuVmqFwCBKs5Uba/wsFWmxNe/S/Gumtb
Aw0ttg6JvZNGSWntiqAD3EMJrRs9Z7CE3sVnQ2/455GjJt7xXvUIT+KfPnkzshno
RKUqmPnXjYrQSJ9W7f561niywa8Hzn/048eCTT0z7TMBDFS4SEMsC1E1BzO4Ea77
MboZFs46miMYYQhW6/upLaVpMb6G8ZZJFxjqqz3QqtvxJi08BjRKO1aLMi+ciRP1
6O+JdV3N+CYkfeZYeJXzF6jiqAIxYeUJzSsN7iCWwBQUOmRCXK3zDkvJuRAl9A8c
WolnpF44KQFONzeUwNnoVroKm2JnAApm6N/WzvmFeIyNdZSXm/dCiwi8dFzQ0DAK
G3iP+rfkIJM3jaP/7seSooRczwRn4Ap44kR4Lg8tZimEPUTqBoh0yzh7xzmXiL6H
EH4S7nE2mqjlerxEPFOY7SJmstUtbQXSswqZsiy60dr25u3YiS8U1Jb+jpK1PjT6
We79oLp3Cf/5fJBclqdrMhHgeXgmhMh2g7Ki93E+EMwT0wSmnq6KZQDU/ydBXqPT
kPMlawKHJSQvN3dCareIUgVmS1IPxxAj5ZKt2B4gT36/d/VrxeLQdGIW7gt/PGtz
fHJjaXi4haY6gh8ga9vQFh2kR7IajTD8Ly+p74ZeE0F3a9clrvDRChj7aOtMe+Uj
7drG22vA6dc2UTDY9EK+ZygFGmYeG9uQlnixJCSR0AMNq/I7oG43E4/N+0wWbMZx
Qt17sy3cJ4iguvUfY1VU9ZwcqFtkJbmsZX4BKXMwCTpcG3jifw9TGoG6LQc3E8dM
PEGnM+fcqSN3wJG4Me5GgiWJLMB1bJY1OSVzAzRlCyHXYYoL+JO5/v3jljqNKztG
mzOpYZtFoCWQiLvEfsS30/kEfpXMF+gsNm2zAMgAlBvSjq63POArXG2OVTAQLWi4
8+3iPP1TlC1ALtDCmqXPSxUmtP8EBncg8IVqBpl3zSkEpDHKf49UsiHlNLz1htip
ia4enOIZetXPcYb2vM2kQSPzkUt1i2O2W/MCFUg2D/659rV5ld45PQtldwC6AF8N
1a3nauproOBH02U9kRHE+0yUKTu813gL+t0a2zAXgmV0jvkiRgiKgirN87PX0hco
iy77EkzlmmUkX4xN7t884w70+aeWbV/8sxF7IhJ7mSNl7BcQp/YuI47MZIvoQg6w
ipIXFoaC3hoyrXXDR/qz9311/LcxYiZkyg+ngvvawxoSDxAZU32E1CgsNmD3GUPC
Ngxez230GH3rIzGJ8S6Wp8D/yjyl48uHuPcYWMar1XZM0Za4rxF4edKNTFM72hFn
iTcVM9M8aAX2pS0drB14RRqo07V7fLfsk4h4J5eqJvxS0NoEEa4vOBzgQYZHRniL
cKFIDj1/vtZFTBAdN6Njd42OiANrsYwDv/fiL1HKJsfr6KJQWyHbKjPD6RSm8xmM
TBt+mLPUbpWciz5bf1UZi831dU3ZknvdOcRvlRGs+UNR1KgIE9WDwXVYXOGQ4Ilc
Ii9ObcNRQ0wljLePWFUEhnt+pS/DYeol2adhMb69J719FHi2L9zgmslXI3KY+hob
arIzgEcuwKvAk/Jd3A717OSQ07P5xo7C6ra27/n9Y6/FMEWIxjfcweUzhFCw/A88
Ro6S8RmqpwtIJ5oj4lrc1nwAfW00LM1Vh1j0u6gPbAcAs+sHL9dzh3QjhAcUsrQU
THJ9itrOT54wgGBlXTEOEQeW9dLUWNKbx7CVs9JyTYRDMmWGlijvs/xvZMqELLmI
gqYG+hCBbxbShaLPVQgmqkVrcVKl87GfKdzwO0gaBIPmcsUE7upVB3kQjKYjLILM
tBVX8+LxIh+3bzayL0GHDJXjLxl906O7xgt9Wg/scjw3rv6m1ErtVTK3sPJfszkD
Bz+CXMoKmapVkBgWgl8cr1cSGtdWGFKotRQbEv9+RKhq+jOdHA2cQ7qfBjNYTDjL
Uc5N33A+eK6p47sTn5x40VGF1fuIO6VLr1qTNAm/N0hUf0U7u3Rsu0ldw8k6Y+B2
8NuFI9yfNGxmd2RWEtVwSuKRgaAzcNT02Xm9Ibog8oUGa5VCe2VxNFk2kSuMHjD+
8nU2akNeXrB03BINDJ53HojETC7Ddlh8YEJtJ6pptrFb920mK1YewAdk+n4NRfiN
m0LCq16pGg8Q0j2gxU0HNNjJiW/bmSWJDIZmCFV1Mo5Akxw5WLtLlOErd0bbtV8V
RSsbxCcPsZesz8mvF0BMN7nxhCHpKqKpbldnZ9BcNDnWd5UXg3v6CSI2k4vGrQLv
1+XI99u77ktYPtoBCJq4aHGO6kh2JA9OhXgMnTEa5zKDsJUfC8bSHrYCbwKzkeGy
UNbQ7vjSQrjNPv/MxbNL9BOOtkQvfFewV0wGlOcysG1yd/coPw5eDEjQotVf7PfZ
t4Fgpm4oYle+R6kyB4+cjQwWY2qLe0qB4XdpOfpzeePNR2SbAf/fwQ9qcBQjeJXw
CtTF39wlt7WJjpLj5S8yI2fx0ra88evjfHbIEJgkehjHBuDHfq4rTDeZv9MElAw7
pT0QFy3Ji01HuF9Tn3eV3lu3jjEJRvIXWNWwRL0ZIfWj9PqT/+RS2HRWh8nwQEuD
hyyGEa2Cbzg+lfQFIBjygQmfj+bteyLwn7ZpueWyejkfvzGAByUhLVVBadxkIwed
o60POK8xsfIyIBAOXnKjDAHmgsKNt5DhShzFraeDoXF2Vo7MacTPwwl2i9FoT45z
27NWnxfe5ilfr6O/CU2SXyLWxWdIIecTWdfI0sQ9WGQDRltZ8CacVe4yn2n+2C/E
fbQAiPeCaZr1I7c8Ecf0jUHT4yAJ7atYcL+c8AGnbd//50xgChka/NQQ2o1b/TWb
8rl/ffw3yGH+AZe+2GkN8tvXLOvlpFl6I0CE+t/Szea+wpckdQ/ftMrSpqqimnIZ
xen7uNHHULGjr+z385hsNdAd4feZ6VW5tR01D7yJz64Qe19zVTxDInVXI/mXBRtF
3cmHyxcVTkevPrI/2JBo4YWkc6yikGL+9Sh3yQ6qk24J+bfMUlbjUfrhx6lvrIvz
Sk+FyIE1QRLKUuGv3ElGgvqhKLjO1ieugOBpBnPRxHugTt6OkHBh2ogBsetPhjWq
yHGqv9VR9L8azmpZqcJDEvLgFbcDIJrt4tqf16+8MQr+cxp/xgFNS1y1WGnFy4ls
Seg0TLd2MDF8VrG+yO+/R+crPjXAXMqp3CwZAdlrHCzr7iAjnV/IUSJyCl9R8zFS
VnOd6hRz4ViW8XY7zipBDkuGRgZ3GCg1CgM3cYSH4yXRayWFsv0oMaM3jWeplS6/
mnqDkP262gtC1MedpmXALDK5xpfOl9ZqZmDIU2obw1dpq/vqMKGbJ+WYNtDtnfr6
7huzZ6ZHmf2IDHwb/x6qElyu7T1KBI9BogXLKNgk0C+i0YUXRTvLKgDCBV/VM4Z3
Rc68MmElDD0A/XTcc+fnv3lNbnhZYFzrgkIX003H6YxtI1AnlVo4R79koKRLwifc
acExZTyYdNMYJlT+4NgKtIo131tS/IvYvlvZ5Gl3Jgs8c42fCZlsAxQUobgcZxnp
IsSVe1xxY6g9K1vvnnyj15QSoKsKma4LPlS2oN+yMlA7EMmuWVni/zhtMIVSSyVy
gjtvYCLQBAZoktPburoRUaaDj8JgUcIds0WeVfLwei9tAOKIh70kRqCzDAzhVZF8
88NyFHqt1w2+SSeyjYQG9bg8o/5l/UikVcujzxth7xqBtWFq9Q8Qn1mX0AgrABEP
+iYUdP9wiNhvzTVSIAKe4DHwJ4KzInk6VmjqISdNMj0OwqS8QarGXTB+J+OFBkkb
iQonB2SPgYL1V7+AICQ5RfICSnscefBr0eYQWkbqnB1VxOEimUGr+XXshbkYEHnE
A7tcwvpGeueS8kaLwH+9YPph/TvQ78tmNtk2w3opoG+ke1A+bF/Oc6bl/iB2Vy3B
eReRWU9EXBEW3iOE/qvzWassO2xtUx3wo6C42aVuoYbIynSSOsq0YbrKYGxOo6r8
wjl13aB1XGMdGkDZanq8T0mEl+9p7pf7ZoDNW3HaitR7iDQbPvtd8ODl2QkNf1Lf
ypU5nSMuaKnW2TyAiMgi73RdqoFDWTkTyFVf5te/JbdxDMF8jHGUaIJsIPiNqy2N
AUe08hoX+gGPkltgv0wLX1A9aEUsm23GmUAyU1mtZwpzQk58wuIAlLUDlJQKEGhj
6XtL+nwRkEPLgIlMsQOKlpuY4OuTB5YtWNsC0slDH1rDg+nczwWfkJftbc9EqnVP
9zbW1F4LjVHpUqZaL/aiGQGnxayElWyiFPMq8NVj7uWQOwEfnvF6AkyEHLSPMOhA
eFjAYuPGKuQfPfqWuOS24S2XXyoVgpkpg8YNYmK1BF3CtbKU4dM+QrGiR4L8IPdX
OXgWdNK1zkFx8h1L0ZCllBkL7c8iQvH0camiZMvA0AVU3fyJ8SeOdKJ7jSgfaWc+
oxtCRMJjCYg79mUYjjhOpr37Y3lOiL9p04PlH6hnZ3ugms300mhmtDtXNOx4/Poh
t/NWiqt24hJ0xJIkh7QSUDvpSoxYg56i8Q56+uCFYgSSC0CHt/bYc3qzzlIvLUAf
mukzAvYSD4yFTQG2sUc2bgjDTvNrBz//ke5rMFP9A5SomebA0xZE7l+EJOZu9Kr3
m36887uYytV0cxjdSehzJWbFI4k61yiJlPHAF/xKRGV/47M+BMsFXYpjOZ3CMRb8
TQqAy/O0bFxTIDp8ZvFd661IbHcGvagTe3AfOc4jmdclW2q5Ra60wkLR+wWfwQBa
0W3IA+O1+3ema3Dii48ROUQEdmVPc6s5Ta7ZQYeqNGqEEaDLp8108DNFHFwCKBko
ypw8pg6jA9fqC79daWdCMndgY9efBViyYWeJQOe1SSFtOy60xSL1uRLX2Ty5i6Zb
vJ1tJPbHJ89UezCRuXuBnSUnzqq9RvbKNXqrYBycM8NWjwuL8XSns2zTOo+7PPi0
FRHjuh/3BUOfXAzsjo/VPs7QBZarzWDecrSyEtcu3L+tdRM8TcR5Uh3Uz2gZb7HN
TL4b5ot5fbt2QqnNIUWkt3fFrJmK0nJuMz4xdjBbGfhfTEoLOltJ4jTCm9jLLkqd
3zKGq1Euf22YOq9uFbYNB4Cr/94epTM+FIyYxrD+VXz3x8ioTfTRmtgvWA6Dfbz4
n/m/qVt/QIAURQXwaUduAR/iZsAxB78/745k+oNohgtgOg8TW6rJVQ4tsNc7w+j1
1tBsYH2f9Yo2qZ4EsOwrhJUXDGlm4LdHjMgcxaYYMJvIVQC9AxJrjd56t7P4ugPz
eCro5J4/PrVDwV3WjQdY5wYhW2qoHdtXx+S7R96Nhvd0Oy9lRixX2aNTfHHQeS0U
Xg+0VLcpW+QWPvOtmyPrYyPOTci2cVPYtsQaph3atkmjdWABs8Y+kvaPxVMdl1c/
Dl1BjQ4eSoUmYWyfGCVEKMhquCWBz5ODWpgWi0zUTYzTlLnsBP48Rh7qC9n4WLla
f9i9VW3HZ/4edZd19pwOnNViHnsJPYFu1E0tyw5HcyehD79iuK1rZSZHdSyLdNqG
rYpnSF6hyi2buatInllLbfCuUhmaS1/tUtZqdghXtVs7ND1Ez8NgYRtxxoRbb8f1
Q9fezP5BqjYxpMbmTpb0oQZRJjpWTXFpA5AWU1oA+HkVTlV/N6rJ61nGFqlI5i/B
JDpx3DiGc7zOkWq677SWq6adhkDwIImQTrfZGsMqJIbfOKOUlW7qnzrui6md0Iyz
mC3HGA3o/dg3Yvjs3pjoUZ2rUTgmSE5JLC1MwwBpvUxSOp7c6G4ej3hFdpQTbTec
RV2/YvrLVt5bzVt4vVeW+WYTJDr+HKXw55BnMrmruG+n4pjAJ09IcvjD+9uDsZf3
wf0i/l85SKR28UbdYoX5zZpa07wckHtqN3s94o0U4iva/Kj6Z6z34EHgnn+hwsUa
On3TTLQ3g09nH9WDameDXyG2siODkZBkriSxwpiN1PBabGAXxji/u7N16vJT0tbw
cfToZjr/o/NnHEwgt8WRRyScp/ySx5S3y12EF1kILXcJxp0ZBT6eSIK/1/p/PuNt
hdj2yLoY1ZPBJFwO+hGUScAHuGwms6SbGf5n0zAoQfM2PijBJiwuX1Nn010UViNE
ilaIOD9kFtLU3RSjL7zw+bCBLKUWMHNUq3GQ2IuEIVdGXZLkL+t1rMqySe9jr4XZ
AKPobqbmkUqT1vwcGJOrKvS28GIb/0n5ngoHXvHvQveaNCoEE0dz4rhbD9uTjH6C
uKd6oLqA5Mp7j5TaU5ns+QrcafYmqXNxuzek2hvzgJAY7a9qKJ19KvXPGK48QdXb
6oqV4yZnftxGodIWCw5RvBMU18bUf2TkDk9281URQwg60XoRB4SUHdHNWCdE5PPU
RTQgmp6dFqZin9/jCEim5D34CID/P68V7cp2U67hIHwg3Lsmm3mW4mSdN2Go31fq
zyqj4MxYj8MT0M2c0UWm0WzGSVOK4Jr+1Y/dsOAKhfFsibREXRFug5p1LkKafKY4
Wso+rF6gO46+tAESS6rIGgR/O3djnvNf7uXYJIRpO9Wm7Z/FnzWDFHVbs/nSnsyF
7H52PDLdemtuF/vN/w9wxE0ds5QmLerqmYIaOT1jyekty2wM0W1VVAIiNPEx+j4l
zv2Rxv6W/Q0JM57Q+KOI9BBAUuKu+tW3i5ihhu+YaGlCBfU0taKiEZt6NXkRXX5y
hxL4uWrL1S8wNAnSN81Ub1L7uTSmjslXCeruyVkrk39pHMgAFoGjq3E0X9Pyqavi
bMcQ42y317ASJ0gemaJDuwKEZUS9fjazQ3D2rf4TDkx6KMmply/ficXhD49UxFHO
Aq2ILr0pkm40lkKWCcAJlz1HpYwmhBkgyrPyU4S58NcdV5Y7VQNXsDsn0EsjiKNR
7eE4omKP226Ge9mw0wzvjnQCh8xX/G6XxOzG2hk8fK6PnpWs0PIp3HYcO3HLHLm6
0bwJYso4JUYuTyXNTwZ0terdmMF7spEfE79z2uI1+BwOhC05M5cMq+ar/SIpmSJa
I8uUoEK9KVdHH4EdzIhReRVGw8P6eC6dVsnzF5uRQz3LZVltvE+P8KSu9asO+ehC
ez2AkIpHV3wBszUj2lenZQ==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HgKYOU4gaRPjXUSIvLkYgUf1sraIwDMcckqLjc8PHujM/Jj9J3RLZsriTEO+R4Mi
A6F422iB6ukaGHOH87d+GTXXKgSRUDsxJ7DRQVBoB6CXh1ocj5BKdJBEk3WhSr+S
lI/OAryUbKfLkRbrw8mYndwVzr2T7Il/4DnLuQkd1sGhryVwec11NzWFqAlbxIUA
0nX1vFipii+QAyTzUHsQu07lP5Dv5TFEeJCGd//n3rDIyQyKh+CXKSarIuLDyjwj
Tjnul1vuPdFnebdZB/Jr60bcwm53D1579Mvu1fN3uGZd5fVDpcNIKLre1S3bGdBp
XJqijFVcpKHYqb7eKgm1Pw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2016 )
`pragma protect data_block
z/bl6AhSN8oXMVzuyi7jE9R6XCg4yK+m19gQN13454dqDK4ecVZebbZcozlKpHPC
KpG2jbKdTY5gzUAcrKYRlI/VyQ50nOLxr6ocX965mQyN7HVGnS0+gPx+ckFXvVrW
xs/rSmGfmpmUWAhGDN/J0BjpsrT7RPhgYqOgoM+SyZgVS+0nhJ6XABRlyb5hpz28
Ksn5v9VgESp5W3tbJt7DR2lNiAo2cUKYIRqTIkNY8ovp6VqlYCmS1VoXJkbKt1Ga
2W+eensmWsWj8hQ1ocAc3d3Xls/luHsE84iVZRikxGsrjIWQds/uTgd0rM4FH7m1
vpJsMlRlb/w9y0OQWB8n65gUAkABJYNhU6Go313Xoh8HWJ8zSyaFxVRZOoD4+UUx
EFnvn/PDJ84rkGeX0PYTub0oOH6k0SbJLATirmlzFCTh0rfBNbVGlbJBH99LKfC/
s6pAGIW/rYDb9yFj6Qv4Gf3R3PCxXjooKYtTKkEg+7fJNtn+Oz7QypdXs8roIMm4
j2XGUByMhXJrQ8wlv0RlsKf3DJa737yCP4r/t/g7/usGXHX2ttTj/gIP9hfMUw6E
YYTh4riobDOK3hIcfd0TB3WC17n9STLEMupGNS+CjsDCnbYYSicAuKsszrw/pwU1
wx9/lALOd8bjY0sqo0lQHPbeUKqASGlYqv2i85QQJQq1FjdKNPtHbib9hw0tC9Ev
uV3D0x/7OW/eQLNhYhUEBom8PNR7p9uGFOFLcXmbaL/AW/dKuk3LzhWmw5peEtt5
8QiktPfaOYazIRzE4wV6BfsfKcWx9k0etzNl8rLfpN89H5rxjeOvx1yX9rojU8I9
cW2RFQmOvB0GJxf2EXuN9ou1/N1J1Ki80QH0MNz0VvtrBfFWD+7UvZfStTAXvhTn
yIbizQpKzl+agcOyjCH+CPoNLygH+OC1MA3Il7Bd9VsY5Jd0ZT48akie6YyuVbB7
agDUDzAAVMqBSWmmV1dO5rL8bixTHRDr3SBrEser2QkDPm7Dgja71mSx6WmPJa9l
UYz9IQ2rd3xA2WaT7uwaq5sSSZOhNiDr+Gco0OTCLvBIVChyX8edVxAify4i/Ewq
0bHLiWSD4hcl3tQMYazCTVMYBOqignFm0lZQlzbSzFcZvyBb7Hn36c8rqUIkgwR9
4eRBl6azgAHUVrvS/BgqX3ZHNvJLOEYVB8uqJd4EBLYLr0qr0cNpxRi2cHHu8ARe
cPYo+omYWSh6P1irOMt/m5tG7Idv4zHFJ/J9JM9Dsp82wLFPtZ3R4mIATJM2gqF8
MU4y0g3Qll4Eb8doVlK6Mm6FNQ4at5xpM5Ke4WVXzNR3Opp1wn8p53YX6SwVIRgL
KZ4gSSiBdGui9jU9NU3wk5k5UebIUEbcf9194lWUDG/ARZwbkQJRvtHuKCMJHa5K
aDmK7CBCtoZLF6fpUFk5mKjDxgpF7r1DtfZi/SlSuk+M0Sc0lVeHSNowGlS13D59
X/RlZCprmFv2mc7u+xDkFuBxtKFRAf2u3n3Cox3bwSQKZCpaBUNZX6VdhgvGbZK7
T48jm05KcZVRi3W6KQAX0aWYmJxdOiLHIy4/2dIhisw/ZhWXS7HtI5jXp/QrT/DH
ZoSn40kWtMJ4FvZ9s/O7lNRKVnKlPJTp98fIsrX0i5BpwoRQ1ruzpELP6PR11aQQ
U32x6X/JtZznHATZMHriymh/YvAICJkbOUwPZddNV2F3ba4wO+DYj5MC2Zcl6Xa/
GmdLQQpGJBpXlubuKO1YOOoU8IayDFKkptvXljauOuO0HHBbNhyThBQpsJ/UeTDK
7ftYdOyDEYZ7rUjFaI0sW2lwiQ5DUVI7Uv7Q4I5bQKLEe3FLg+iJey1eZNnQczDW
I0NGe92bLD2zzZXa0OpQsKA2rmEqfmRn+A1+0DUy/3kmOvR+c/AlAzfOM0uPnMJY
HG0vJIKutmZR685rWFsKiSXeZCpmtHTLe9yOsxJMVcicZYjaVuSaef/qwlNbxcNr
ySIohVlDGUV9GaJcrAz9crna9MQd2kAaLdezGP0eIxol0N5rzdf+LBTXB6OIQs+H
fxSjSTwNQmfbiqP+J/D6pbR27sUTpjfLP8DVOtapu4K3/Wyki8RMxq14CyRwza05
bWUYVCNm+LuRSVdu4JF4Mgx0VcTMa/mWx1jQ94XhD5Yfhr0a9rf6tULWpXtca1Gh
hP+UoTjchGkN/A2Knm+kqZuiK0X8xMlw+Rk3ytmf47D9Ti7NVJVabkW6sprsJwTO
lX01OHTpmtJfGvDHSvtog9D39F8vvPhVORte3U1bY4XWIbONBFXa62bFaBRnaJ8T
Wx6OP21WDPUJeZI3MFc/jvZUDCUdEH5zfCC3TFwbh8C9MJg/jiyyfW0QbIGQvWgK
MLpTGKOtiJoc9clePp5/apZ8kRebCKlPSXp8Esx4Dinu5E6RdzQpjulDgJ55XGS3
cTtWXluvUEomcvnXlW5GEFWns7TtG3szIcrpkEnn/Ye3K7qsUim+SyqxSoohu0Yy
CBCUfUkdStHzSu+dSlfma1UDeBMylN35GPTrHDApLlCR1y+n71sQQeqcyenbt8AJ
sK+Nc+d23jOHZeGA3B3VyH7cFahOm704BZmqbHKyUPAYwaXgXDu98nUhc35umwNt
Nq6V2bQjR/6QGMJeMo8GjGn6JY//oIhDOo+/aTPtqaR7B1iQKEC3fj9fIzKGOjLc
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
IOkIEipAcYu3JQEV0/sieb1CIvnRlX3a9JO96qOxc6kDIMRLXvb/jQgsYI+KPxpM
K89naN6kHkdsyPFKIn/VV2Pjn5wztcNPphpiJJZERsbh33kveUf5WTKuhxoNM6G2
f/x49ZD8qTUjezsicrqOzy2m6ua0ETn+YkF5QmjQqMDgyuuJYcwQzGQgYKqbS7PY
xy0WY926Zsb2img+aLOKLor8AUzqNyNZ6j+3dkIecri+4sYCoS+lNIA175qxJhhR
I00F5ok5pyXP5FbWuYw3aJsN7t/7SqpR6NmnxHld8nRSfOYwABICnTPkcUXjUmlp
i4QEBNAZdUPWKdXuJ4jQyQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10976 )
`pragma protect data_block
BScf9kOaMyvFES/zE4hvMv+xlq5NU8sff5by3KAr++U7K340AP3WbRTAuirnnakP
hbPyQAP+Lv8D2y5axr5b03mNfI02BnZNyBedCWvAtQOgyISfUGP09rq+PLSR0lqD
EvjdQVNS+RPMqhRNdGJXN5h2S2DjfAJZtwxpbrq0PaoIeeUi5W6ZMinnSdtcYRxG
riKxhRAiKeKBc5Q90ByVc9e+c/7S02RIMK/FBcU3bzoqS+EURSfdBJ6jQ16waWXz
fkHx9RebDO43qYwDOy/3sT1W33JrX4aZOgtO1box3mRY3WEw21fSS3EAgUM/6JvK
eOtiS08Bo+tZXVP83u+M7rZGOtLjlk8Yi0y9X5FQs5Wf+oxVU+MmbQZd7ihJOXQw
pJ8ghRyQpO5OlpGDWD5SOjZRVn6qlVB7tB5Hbds+P5mvJDPnh4JE66u182pign2u
uHyIZS7MiCj24HFIHsxVw0LgTB9EmFrDIjEooSbZPjmj6wgVlCc+jCZHrWioFS/d
1vtMexJMkf/bAaLZLFj00NoIiicGZ4Oix0kaUvRw14v1YyDpse4LobdI1ilxBCrg
h8H1PzSWXrFJzjirHSHAHbUJfh3WjrAtjo0/7i2mQKBw9F+T5Syd4QTTbOypfYFH
Rdh6hUkLEeAYH3wP4Czep5SrPK2RI0ixBidiwqwYtI5ZQ/bWc+3hMkTkNtb7lw+B
AKp1z3/AnxMNLYWSD5UtQQWFOGpnGvoIb3yzlRSwziII+8n7Yx1u8YdxACruFgJP
J88WBOgh9Qg2RrdBMqIaDqA8GPxs+LkKrugz+6gR7qanDR88YNuDSkSyYDVD6Qbq
HQKuTItzLS6foDkl3IQn62kJp1lFHaGS0hhbmHhhDQ7VoRwU+38Y+7iUmAJyqYVc
Q+4TKp5J1JK4tHbGgW2nmChMOs59kQd3G9Z2lWUWE62nwb5U4r4R4KERftwioezr
dS9O1MelURmP3R+EPmiGVJSY5+fTwaKFPMEYpyEO/wFTiGQtVEmF9dcGMsAFHdBX
NFFI7gTZLvulhcJHeobbKA2wr9K0+fdY6L0JAHzAyYjI0J41Ou7IKf+YSgT5Mh9q
JSpHia5HRuHmteTaLdpIdcONWceAbsTwGMetEzXRvTXcKJ6vhcHat7JYoxqLE97z
KK8LD0m3xu1pFOqPF2/e6WA97t46LdzAnyRNoZ7x2/UfkmsFyj6KmeJySukiJhWE
zg5EBU7YCpFkbJvhnr2zplRFFmZpB7RgwZVIiu7hQ556k5lm/Qjvs8IcRTH7qJ61
LLtCtYe3Y9G6EJ0GepSfreKvLZrscvFpv0U8TfWjIfFHVpEUjpUkuR46gNY0zwS+
DAcbpFwoSkR+76Xtds6n/o2WZ9fGftPZzZQFqOHm8Zy68idc4AS330dKg92PiBtu
KRzlbg9OxrVjmRLJ5i9JB9RP9wT6e/zZluJ8LFI9HnSZro410ItDoRPc1GQoJ6bE
HqPpItaeNfp7AEvDN9EEp2rfWwRG5uIdtnj8zeU3OaU28wxT7aH0Ku7pp5nv1Qjz
tXc5Jy+JA5MR8RFSuCao+UHC9R857M7bvwrdzawXxL+tQFS37HWBd9aYd9ggv/Bg
ZQX2BC3xo9DoT/A3wah/zhlj24UOOdwOmL391gvJC6GTn+iI/WDyT14i/0GLf352
xh0g6u0LngTeQAjkrhouZmsZeSEtEKCcTchYALmdsfzPxhXVd0sl0NYdVDX3ow20
PPLNRIA4dUxPEwU5Ln3dOl21sIUZ8KcFWWY2j1Vz2MQmEe/hvf3qcM2/xvOSASHW
ibBtPJTzWmAwbmYepyrkc6DhUpFkkivYViIf86gYpw9y81oLI+vE7tqKwh+1l/U3
p8YcLFtCN5N9Bre4uBQ6XfojqNdlV2lcV9/bXlGvKT3ptflsnozya3aAkSQ4TnkQ
gn9IDZ7DNoX4HaZxWPgjeq7jNrU3j0rOTwEAMt76TTj9oJNhDKuE3AknkAUUxG0o
M0P4mOGv+JdsIkXil5MKP6PA6BpaNlXxGq5TV6D7Xxyzq/7znjMLznezoD3scTOB
7fq6Ba4w+mndyL08Mn5Ea22GQVc6tK/4qYH6Seq0d1DQAxSLJaBEvpKlJKCymHLm
p0nEd3iXhFFoQ8IDlG/GQvtRPGsQbp3VvPkKrJ9M2VI/dC9UzlqlFo6UGrmy86TS
bSv7d8sgnH22+xHbGKXYRP7JU0E+LtPIrkcwp1AYR39leqsKuJbbw3XpY0CgeRkI
3fo4y4TCX75ncOT4Al2ikG1Z9+GBQFZKWO5vqefne7B3igwlWjgfCFcmGTyEVi+n
S1I7hgchLBJlOT5IrxY+HZtsRpSwo6ZGoVj2cxuarlcgXZAx3TtCqaCliVa7+T0Q
POJwd2+tC0OcWsG506pBlNDrtBBO6B4NHg4piiOq0ruheeNPBEH8ynl/BMYDwR84
BomVU+0SJhw9c+dfUbAd8kqbbV9FHlAtybpqjSWUW8Nrrdt1oeq9w+s0DH4krW4w
1sGDmQeaiF1qZiZG/PnPqqLkod1WJK7Sbr1KzFvmt51PWdWy24rV+IF3u0Gv3sFf
RVqw+v4HpSK5/bG9GX8Cpv7ldYKdYIcRd9N7RdujjFgBs0W9cVi6pZN08MJfx6FX
GxtcrDCuK2CLPgTceOZJ54L5F0QhbsIk0zKl3cRZCzhnG3AIgpV2hcXxYYC7deTL
nqx9sAe5LQU3pqRGYpCpl3Q9g2nTSc4aIEEz/yg5OZyTcMrldC+LajsTt1TKAICB
vylyYvLARDsOU2f5ZH/Jmpa7L4KoMzlkjrfwc9yDKMTXYWGUCg2nC3rMK7WGy+w+
+zjOuvXLaDTswCYITTidZahH6yCYUenOcMbajCdMzyEmtqOCDvYzEXHnkWUuP0lC
ExHPuLhJJEJzaO19UPtWosIu9U0zTaEceasvua5kObNTAPCUJfcstmLngatkrrb+
9fdbbq4F6vWQ07py/Ck2O5XvfIfrce3Bpoe5pKNxUhLgSrPEwFwoXvez1NVV3S3/
aupLZrT/NWeRXj3yKgpiq83J13yEFQQHXF10lcB2+BCkjZytA5nf5PmW8i7IqidM
MeAXkDXu6euM3kju3GzJD2sUI1JvNkuE6hVwW2e1BJ4BEotg3oR6tRZqnwZYX6fh
JNBOs6uTHNu7by2NX6+nl1Fr0TbxJwl+pm/HLYFr/NRZ2FVcuACAOVRcC1tjmGpL
mBjr89A5w+7Sx7RDIPWLqc/Hsg5la97AXj1YN0LajLoPVH/KZBbZGwZAocBHrnme
ijAaHXHrLfMw5U3zDsl0Z9Tc01qa0X513XHeX7eiZXwVEBiUG3swiOYsCc8615HS
+NhYUkM048L+kpkLxVkgK8379sXmRILiLBSbLJBuNcGIV6Y4n3u4m5PBW6E/eIP8
SCEqyzRgJRm42BijenWdbaYBs2Piadxne8hO1pA03JQUr7LKxV1rfXjAh7XSwKu+
4Bxpjho11WFveEaU1OyXadGoZ55pa4ex71fwLe8Hc3vL/4WZIB4b3ZT6l5D4tb8M
HC3OXC0SyRG96Zx3nTjRFT0kT3IpWSm1ui5/QT/OJuTbGGa3LfoDrQTrt53RufUw
QrZxElk7C69V+EteQQV5xc+K1WpT90wOZKK2ea8remKJPmp9NGKlmK92D1yYrfic
zxeHxny5B+h6XlmV1IWsZmuUXD9klEhtO/bNQy5/Q0LWQLTf+anmOCowclMl9EBL
oGqqO13aUDDY+8hErCA7lyeeP+TpHJs2gkHgCnfG6uzY96jStiDhiQk+lXS15fFP
rFyx+a+atAwtvPTrJ2tVqswq5BC5xyVfmVN4vNmeCHgSc0rDyZbJTy0e+iul5+Ls
ntKys79PgmyAsoa/oTBDfTRC2ZbKdhUZTLH6a8DvG0gOllc+BpZMINXXyF6HKfaN
GZzwX22IwiUmobRp082uXaPCPKNkl71LVXzoiEODLwK27w9PHdVOyrR1w/9STTQZ
ragUHqIvGMoy6I4+TdXoPd/O1S/owoOflmEmmPuo2mdeQJiOku/GBXNL2nxUQhJO
6nv6EbuAQ8Jc5g5bmOcmiMgz5dmKm5IpL/VKXluyBgneC4koJlrBDVYUOec16SEu
0m5gNXDnU2N4Iat3mHHVScPLB1OsVtepjulqS9c4XkVtcMPhfq2FYU72jMmuwfZk
RI7WBDTzUh+3eShSofdjGa8TTEL/GLgPll1xcAErtVu+t7HmgishsCd1ETD1l5XN
2YHt+OqCj2xkzAx1nTAWxxloUn/c5f4SMAQ1mtb26Bz7pi/aDa1CVDgU42goYL7B
NOyRsTDboOsBz/Qp8gh3ZmkVUyRk5hpZ+095WoUpPQ+My/pytJDYsrklcpWnIdnV
jeb7t7AyKLi7AxF/hxudAzQLFlRpI7zlR/QgdtSzlp5MHmD+5IeQBRoyF5kMmuQ4
aqFrdsykKcDrl9oFZl74xUFGeO0IwdZoDfroSNzPcJwbwj/2z3cwn+2tWDmI8eC4
ws13q6IWw/OBOLRCGB0qRxXMlQ4H1jyyL8KJaFc9DzbRUazM1HAb94Doau3PABll
5iYNYiPIg51LGZEIymIv3QEB+CY5BC8rmRp/nYstnb01XokFG68DHKdnFefcXeFI
NX3SG8YTSOeq3ESZVnS+5AWFQLnJH6PfbmaMmxR80RW432naFS/uRKGz3Wl1pjSg
QnNmRyUEnfQKrZJLWxyLXoi1WHDuvwXmEyGS58S7XWbCBb1PneArxQjf9qAiko7D
hnK93u5BA2osYVOishhTColq4OLWvJ3ogkx1l7TDTeL9KvtVKzarcVHl4PrIJ9lu
Q4Tulgs4WYoEFxwcKYSrv3fgZyVy1j2Hhmo7A6W61DI7aRBS6F9hCwUFIS0volX/
oxsA2LrwtXN6ne1HD3w9k4RrVPSFkYSwF4vBc94TY1PPdwhVWrQ0SAj7dFOo1je7
2wGBAiaKJMdmQ5i8qBr3QG5I3xuHT5dQFacsmNkCD/4KG3K4h3BMt6m1zzKt8otu
WmSkJUDEp+2nCaR0uBtIKQQrEN4LTQDjLySP6g4jQN7OJgGJPSILP1sPo1SM0hpb
FmFTr5b35L9DIMOkISIt1KkWGlmz/S0h1zY4jnmq5Uq9dJ+G0FPaXJBKPn5x67tt
RHER9m7fz3dCpaTtlwaCG7sVlVEJVdy9FM8r+X9F+GFHPkNOPdbU8Hq7aoWVC5zX
GwJ541id8qjIfiTCwUm5M1XDShsLcatDyMtPTHY7A7YLKMPHZqv01cimvwXyhQbU
/4sADGO2Tq9ARoP2NwcBUdwP1BBQNJCb7yXU0yPy1weGBcmSjA9c9tO2n1H7HMff
Gj1fxldAZRIk8hfrrGNcNeImg8FaIcIObqkuufvYqP/qrmD6FLUUYxNjs5N62HbK
K1bbC4QBYJnX6igTyI13xVLCNI7Ug3E+gcK1VdbusbdP5Jpa+si+yB6uZnXd0vQ0
ZzO4PIc7onQOkQiLlJWtFCUZBmQLuEOeEyMxElOpsAfb7czhK0S83vEimzGQOOpf
5hJf1GwX+fT45BHNKSdnDgp2+cDDSpjvkzWDH3Z9F5A+KHCm75BAPUAJRzsEu0H4
QaBd46k4rdxD/IDkkQjs2n2wje0rIW8kfqE3rMiTUwY8AkTwZlTCbNbTaO6Ecu5h
oEFUh5E/kOLSmcvAthl0r2KTCDEs8SaA12ZjGZZKCXsqXBlG0N2gEdcJFyInTdwE
Oq0SfC/w6fUpuJP1HQojQtKqMR6lvBEweoVBms7JrqQKg5JKhCodRGL+B94jU5l3
kvE28d9wO0HGm0JKOR4G6nlohwCADJaYXrhcwOJ/8HiageNIdfa0GdpqgR99P7Fi
JSSdl8RSnMRSGnXQp6fKGNQmnFu5IKW8yUtLJk9mQnPuPVBmVrSdA7mlbDy2rHfD
3/M0Nboy1ovE9RvW3OI+gN/TixbcFCoC0Sra278DhBNZAjW1KWZdiyrntgPL1SQ/
Vp7d97SYRPGQ/rcMlZs70y+OuPbXVZ1b5kCAMDMedoDK/rJ5hHf1zwcmK7ki9k/q
wkh9FOSWu2FuaIN6C9jNnCj9HdZIWXb5fOUIkYfxop8r98Eie31DzZRCqnuVnhz9
DxazWJg3Wir/y1fDjCmVZ4QQGGG4v50agUa6MDd8sjaKxnmUOwmPdizpja2FfFh5
7jwnnpit9oHVVAfGiNuTUlS2M71A4TGjed6gk0pRbYla4FX7zTvkvQs92hvw3AkC
j8z/DeHbQgivYL8vxl5Jk5kWIDMEhj7D7plrwE+nW3XKjWb0tNPPobLMvo7pNPHo
jjCmwPMDojlWPu/VqLWnomg5MWwBX+73Pxb5h7P12XoMT8Q7xggclHYx+Z4/CMJt
MrKx/nuUZPIv+Surf5sMmtkpYxvXyRC2ytpl1HBb3q9wvO4ZRHL3nwELvEmHOvtp
0SMUp/BqGWgOA7g8RrIDjfKucn6H1FY3b6c+56Gq9w1bxh2jlMVCOleqDwmHXYMG
rzAbP8VW8nhcQQ6jBxDzaHmjrWa+UFt46T+k7PcikrWA2cWLu9RGDlM6dq+dnl2t
NCbeOc3YcxwVTFUKcBVx6ng93/gU7wJ5bWmgwQLuZyiRODxtigpx/+/HkgHUco0R
hSx3mrpFzTc7Dc0bvFgyk01tCAwddIW7nE6h5GtTx2VNv+/JanW0zKtNz11DpByT
b8AzUkBwHBS0H1/BcYjk2xnyUre4C+k4UkyPJn9XJ7lba781ynXxoJ3/XbHxsVAr
1ZmQWfvf/74NBMQ01njwHJmXhZ5I/kT4LeJHhFOA671qWT93PbH0AZjrvtiZ7YrV
govy/izyQqaTCNgN0LXdU8FObY4qVK3SeFRruMqX1xVSsjFp3dV0SbmWo/MNTBqf
Yqjwge3QN0Ppvr63UpayB2YlpHRX6T7clCbYNBs5IOlkDQ7WDPR5Qv1bBaVquwQg
loRMhQfX+1GozUIGBPepQvwCvkz6A6cyU6o9tbNyT+1msxq3fUEYzkmtA5cnLFHg
u5AL2cs4FRv/OW9xzJzt//x6Z4cz6mIJlQ93iJwwUXDShIYCLV0u3X1sVYJ26K5U
7eJmIRZW/F8QTSgNKUwR+kheCRjhmBLscTQXsF8YFwVFJ3zsAYQG5tmKoWp8Z0uJ
uYG2E03QiIO4a47UcIjp2xRFBqlXqWuSuPPTFi5hmvGnpd/bYSQqCrBoUg/Hhyqc
p7NHLnxmOpQ34wjrbGNI8ccf3Iz4cJGY0K+kgLQEvrK8dvXib7MrtiByslfKH19B
zgW/AvQuCZeIbB9tXK6ucn/EEYif1Bap30H4St9WjrzlKVO/wzsOLID25m6sKiaL
sR5Sim57hbTDRZTF7EYbExTBF95iF9BvPFHkmeRzGavuUqa9DazjTJJAgVlEl36N
cl5bKTNb78akdbuVjHs4ZQvA7Wr/YXvGQnJ8QU0tr2f8noFvw1V2vubfsZac5DZM
6kDvCAp5J6Xw7wgksh9xJgwnkY1fCOl7AZ2buabh80NcR+WNxdGbRZqrWEDxyUNf
7yPzFYFWxE+FS66mvJDiLy/scJuUjTojQ87xJlHo74WKrfCxxkPVd1jLtyCdbDmS
drkKmWiEeEQb5v/n3jTH7f2zMuPLMvCC2R1BYZU9UkV9wjU2aGSLY7fHXhjLYfit
I4xv9tCQbft8Dk12Pbnbv6pHQwPWeCFwamn9LGc6gMCWE36Y/VVIPRnhGK3zFrKt
wogK6iJS+5t6Z7C9kXQMuuKWHlaBVDJ91DMUhL0cq/STQLyxPb5EgWX/2hEnKWMs
qDUlb/XuiaPixuTKokZxROvmKSdP1TkA3/+wRK2kBFZ7hBa5SLZDYY396hOYHrO7
PmxmO+e+TrOcmk8RK/aZGGEAP76udMaFi9IOGEcLrhcmdmXr84lLErCt+382LJja
UE6q2IJiVBSeQ1e2l+HPHI7r4SlUp4c9w4JK2gx4+2C1uawyTVoPXXSNOmSleBk/
7byLaDvjzuTpmVjuTch5KHPu1K3XOSqzGUpioE+GERKof2In2xurN/nIxeEP2pHS
Lhv4h5PxjRQrDQEHyIy9wJtid+nAax3xp2aRhb2TuYbeujcqZIeHBCY5keq0LHUr
Pxs4zrSQoDgrCn+Vn3fjzGA840CZzp09VA4qSdTUU8yURN2IABA+MrB37VyVRdMS
2uFrPaKw0KGZytt/0G7TDnYNyPvRyHEoJjhOGax0klNaXTQCETa5vS6ZOphs3ELA
2Vn8YTa83ovddrRjo39xRR+h0YPQuVrQhc5sX7+NsifFNRd+RigBVXM27AdFF2Ie
EojNtp0onU3ikl5uV5eGq4G0jGEiViANEUunbKtUFocLLy7zsjfgtlvTlBZ6Wb81
/Tq9vcm9iyNoqixI3WM4ga0Xf2rhMSXNu6aAmf1Bws+dx8/KhlCDhlOSM5YtyKaD
9hwiqMWjcj3eKLMMhme2Dn1Mzqx3QzndyIAoX+oOarpiaHuqVklUvcpTpf3suH/Q
VXM67RiK7pQ7EeFeOjWNNen6pVWIVq20nobp7Hu+ntXH08g5kK7vU/V97hC73dI6
V19ji5aotDJ5sB86fmMD4KXCegLauzzOdPA/dXW2WjH1tn7pJ435qhbAfe2SPDo+
vtjL2OhI7hVFTUUp9MotT0IcwVueR7XVBbjuGcezz63T80755GGbAIm8Trr2ReFW
N8h3jcn5ypjLz7Wpqj7VWBAbSlik00IfiYgEJtT3+OuK3w/iwNtTdIyHRjXyaU9p
jPp0GwqfyiEpI3JkgYXDrl4zTGd8we5NCKXw0zTXD2akat8x71tP2iCQxWkf8Hfs
DdOoebo8DXDOgwe35Ve+rxhVznF2+XmAJzM68rtIQUkSa0zpbJijAgIRb+PzZyqq
S8K6GdwyPqwQLnn0Ry/JTbNFyk+Gm4ThKoJGOBWM8SXQ6jgG94WJf0zBoUKqFb0k
ZowZheZG95xyRwlfRkDblLrodtFjc/rsTAXzjw/Q8NWA4EfKv/83nSE6mUTNxy47
PbT8QgwfNBC+CPXhS68JrbptGrB+IngrarQv9aa/re498RbjddoMck0ZMc7yHw6w
oXv1a2aCCry7CWGIRxhWeHqXQ4VUitgzCEZBkBVzWnIeASh49MqZdd/YSyHV//wv
RKJl+Eb/D0G3ge+pNWUisdpHuuoZjeNtBGcAjB/LTkoX4Yj+SMJ2bUYbbvv8fH6S
tl0OWkwYjeGy7FiCjLjW5+9a/b1bZZ9B9wcJ6tghVoqvNJdLh2Ex/6DmCb2U6cvc
i5jQS32bxD6QGRD3KiBoqmyESAQai92kkIKoVWuy+IHty1Q2Ch7HDs8HhDObC6ok
vluC/YcXshuvVn+awfXRKv7abrZJBHaEJCAybrZ4y7H+vq7c9rpD5iuKrxQYiuVz
f4Gg7kb10HhrZPrMxwx4lCFGtjPu2SxZ4b7YNKWWYCuccKcfcbgmj9boKglQs3c9
ThrG2LDzUERH2qcYFAFXiAao48PjApDsm3fWhAuNF2jhBLeeGjZ77qhPGpJlxrEv
trTxf/xtCIuPADiW15Id0G2h8jeMEWAr5dq0zjg9jYh95CXHi0kzOHhjNYl2hoJv
Ex0Lyp1BhA2UtxWsbHpcO4lowdcxDmickznUGJCBO8zZoG6DXCU9PSd7hFF6Knl3
CZzk9QSqd01pWAal5gI/nMYqIf82GMTn71cIn8jei5x5hC5TJjvtHecqatRggCeS
wYH3HlaPUVyL6IshQBizKWnmW6wxiLz5shJHknT4ee7jXgK8PkcQ8RDq0P4Mx9p+
NK+SEkpt6SIF/2Of3Tle5Q6tndy+mpUYH6sVGOTjbKM3FUq/d3mkAIcHMhiATuCw
fVVBp9J79jaVkNLG0U4nz+7pfkAy+REwj4FuKHcelYft+zqIN7ZdE2vgFImohBG1
EtRp+DeUyQz9GuvJ4RsfuRXHeMnLIKuJyJjSEjBOGuBIRQw/ARQafoL6fQtDkVO3
5Htz2mi09BgiFh/QhVr2F7pZcRf7TddPXmg45JJS7C14fQl6Cae451Xf+joFGOte
13P5U2RKD2ncOxvSo52psicWZ2y8RAcnkqJGSu8mmc+atgZeLF1LhqwVlgaXjOxs
9f9zNymc9NytZkZRtSBvYAIOf0nfpJXpwgmWyRf7EGZwM9nf1LYKoEbRS8VQmHZd
LwaEFSr+svaMThioI86e/wikuRORGkUQlRnN7mu4CW/rpE+uNAY7MxEOV1VC8onc
bLJyIbj/Oh2RG8O8MmNoF+i4jfSsn9vvfuCYIj/qwZHDmuGg3nv9WyNyfAfM83PB
U9y4iXB+vevuwttaTxPX5YUIIHJMHryObQ1QAI2iD+Drc1cXq64QXdBd+tlU72sn
tKTRuY0yDtYzr7+Q/Xi4QpSm1dAFI0lwSaaZORxikFiHKM6dUEYgS9lg5fgSTW6K
h/UB6ESitX1L2VFFHu/IgfNPlFC3P+ZoCEWSuulNNnTf6Y7t5bx9bKsnOAVo9DkY
xkE0wRu20nOwnxiopIZvGi9BJe0b2mZ0hfUnmndccnHDfhSXXyinofgDpaNgiZff
uQEt9lZrCPjWC3NtJxDxPjyKhUhzfJQdPJePNq72etRyiJp+fsFfd/oCq+Aw8VOr
qEIkFW4zLarTwnpx+g5D81V+6ikz3cJvX7AspuPXIkF/FHVWEvuzH2Tb/Jz4Visx
fR98odqZOFw8uV7Q7tPB+Q48Z3fpbG/thLajGm7qdZ6U9HJ7H5Zj/O/6hF8f2Frx
L9wWMCGva1DoRk2jnCZKcvV8Z4SibRQOZZQ1a4Cy7CJAajMkQzcfyn1pG2Ba/eTe
CwnuTZvFNJ1jQ+tIGw8qTOjvXtlFRFy7tYvOs0v9t2neErnW3oN3TUSd3NhEFwtx
kW8yXZOB52hPZHq7TuysCZhvDlSfRLn71VeyvgLsIm8rhdcdx1AJ+A+RhR9BYWce
Zfa0DvWWMiW0DBrwqqmiSt84dFq9bvkkq8k2xH0OI6sID5B4GaFBFvfBrVyJ0mp4
tCgeXrPIk8evMo7me3wj7Dln4PX9MB8j8UlBgArWwbuaeRtzmTC0+X+1kt1RniYO
uyKKSWx9m7AYWnowIsC/pfDCN4gz/6Fu4xefgf61wpYzXOgUMQop5tiqCa62gxjg
gPl2eP6er0EalPti5lX3mQiMK8Cjpsfnnda72/tLGNqQbcrS4Hpda9ZpLzNTDPm1
WBpgACltSX6HoNRo+nZY6wCrJIkIFW/LM52CbqWiCIwMn4QymBtcmSMqUfhpcyHq
wlIhjWWGi0bbHzYWojTW1OARHzvtNrTixgEluOWQdUBE2V3YwznAMdDpz0nTtOPq
qWHx9VIIt5+6IQeXZv/oLfpNtVP7o6XVKlNAOaqg801k1tUbEA7zZ1ZF6Boobq9g
yDYzZFwPRmQH6P6nRgbzsfASCNAWYjjqnwYXY350P6ZiQ0qwki9xcBK+O3GOMRXS
Pxn2mTD015WnJOjZb2zgfyIKTxGH1aE0dnKS6mSxQhTL1UXG2CH1a/N6UtqjPMmM
x/S5LOCy0tv9YPvY/LP7/7IaUtz7ttGZU3lvQBx4+h8GoxYnpZbzZ0CzpPnMu2vr
82cDhUaBUsdJGucdvAbcIP+ZYtFe5yoBzbRF9r/CEPggNe+TeNvOyXrYC/VCuUHe
p2lwWRi2kRAN1vB0KN35GhvoJTutwUJN7glknfHBiDHnX78lFQO/qDdEdQYM+OfH
yqryB4Dos6BkSePjXd6pVp+3BxngVQKXq1SIu5t3S/n9mTCf2kuZZkngdkLfGIU2
Ie0IJrbAgEflXbpMCSB7U67oR45PKLDQofWn/YN5O/CBjkD3uN/GDR9xyyvnqxdn
mrls/tJX41dtpsmyMLHN1DpJW1obXPhlL8ywNXRrfDGB42tz0cEC/F65KOELZfxE
TR3aeKJXqiDG7IdVWGQPnr1tWjiKNGONXya3xGO+XMZAyyxKNX4p1PKVIxRt+VgC
fs8TKBvo0Vu84iQaf5bz2emFAtbowA6OzlOlGzv9WbMygjbeTdlXvA9ABLDUU32X
uvgnPIYFqwJ5vDGYdC7ph4rShKlxQpSIInS9wtymkfEVeIAO/8+OrykFXGQbMt/e
8Vim0Wc0YkAeFuPsfwrbgNIUYvRcre37P30fiFxFZR6RM7mlqv/jRT5G5OYjBHt7
TF9AOyQGaZgT/fNEdAZQngJwNSYavzlyHJfZZunMyIAE8tEz6zI5tJv6CUP703r1
5d5u1dkP/tfuHwO1qNwf9c18VebFyFTcz0pDMkTsgSNVnl41PpCg97aZn001h28j
PgKheDrDGs/F0Bjm2Y/S9LkgS9wPGAltMj5ffg1OioYSSx4H2eq/aJfopPWn06PT
e2bnFnHRge1+FrqBQ+BSfPPYPW50rEOvx59qL6nj6la8PRIvCt5h1yNa16ndC+QP
LzVerQqBwmlpCvWpI3tSlJQ4N/fIbyagTVwbK4WalwJ2WAL2sI24OHHcePhaZPYP
Y65rE3YGrGoapXUjwL/J6SsaZROk0KmijJb7agjRmfahe4VTXpmDrluHPBaA0+op
F1MX7lX4WMNgvKhwNaAqsLzwwTES//+Gq+Ar8lCOK/F3hkfXYFM4XIz2M5DkJ8PG
sFu3KIq5SL7Ep7sCNqix7CvN8KO84dOPsqB5JPsoF2o+fb2ZLV7nI8xPn7AICnsE
sfeSsZ8IDIfSqDH4+x8OlG0vJM0oLvMjygGV08WWBS+JhQu7QrmXxUE2LIh5uazs
aNT940UCQowb9PRZL6+PmbYzgCjklYMB7qyRMeTxO18cXoEzLUReUdMEFJbhP11w
MbSkwUrss+1EvlLrKQnZGYfbyueHL44jNWM4yKUTXW9ujKAjwl5NueFoCX4QrfwQ
+hoNHdSbwMMb3xi6MhWO63RqRsrvqSla+scAGWgd2NWt2CYFLGVob9kGT9BQKFLU
9fo1vt8jetpgcQe1OcGIGMIFieXmpM0IiuIIoh7anM47hv9D4v14AslrO9RGfRPi
tTQ/9Yo8zdrX0JTfNTVxJcE/1iUwkkvAGkozzQ4sOAKDDfzk3dls2zH1NaqmJ2cc
iy7gyz2WZhb8blBQ+M24yPmMuc1gLnLCHAML/pzFYikxrpcteerkSvAh02otlQm6
Yt9X7xRixnlSTJCRq9Ma1kyZ5fzmg2F1iWgBqpBkUdJetXzQZOoOXjTKUo3egEdC
K+6aBTdermKxUkqPzstBEzXNa+thyfxL4puQ9+OInngpz0p42q7/AjKKZ3Garxux
IQ3qp8VuCpliGx+E/3HxL7xdz9Uwr/+3Z1KmIzUAwQG8mYqyot4EpSSpSassGPBu
HySxVQpm6hArxORcpuqGxknL4xed62BTFAr42nqjV1AmBH2BF5u2PEM6yNmh+/Et
+gl/EBMlgbUy1zncF3qkRY8KnClAVtZ30pOWNcvbyeExNkt59lltTuBVYTFuzfJk
sKIFTtv8A+Ys2Jo7uaNPqCDVzy7FbeiINBjZ0LSAKPMJ2FYfDGJa+G24HvK19lrd
nd6l9xa/OGOAI1BoVy0U/r882UeUmhgED5L/SzXR3jv7qLRETLhqChv2J7f4Heiw
XvMy74lZExDaaehFE93LZKAGqiNnozpoypMaJOJa2b9T66MnLbbWajTEQrU1bMzZ
KJyWKdi6pcQBR1Z1C7/SRdQY0RjrGyoW0x6WGKWaOJq5SO8yY+oVaktwK2YrL81o
YhC93vLNDclBFXSEPok8JMaMKz1nwVdxH89wbG9MQRe9VS/j9IiEkJu7Tgoz3uIO
MnHC/GWMoSS9LtFB52sxRhd2jnNHFArsfMjgia7LBaexw03ziGY34Tsce/u2ltC7
GUY9vtwmtow/S1KW0DwVQG3z/UKApQ3lBVOkuh3zqkZtDi058BETrHVNFTSaYBga
gMDbvrg5uCgPwp68PNWMc3F4MgW8JlgIbH6f8GOX4Pexx4jojkItVaAXHW1CP/lJ
sE+VG3p1OynvWYvrJcJqqEtWnzeT2BWS6xSZxJ9NwY25un6CZJpv36LFQMobFe1Z
JjaE3Ei1JR3ug3dFYLy6PkgH4GoeJMJjgieQnHe2JJg3pSKL6V3v4wjplfY1RB/H
xU+gsTdl1yKmOGdkBeSSpUK0PHDp1QKYxqH4DUwGk9pLBoL3s/SWyYmziabmFJBd
VqP4Sm6fGTTfZzts2x/eM78NgkWUwD8zA51Bdk3R+K/pNewewl+h+v4dfTG5U+mf
BuwzfUSy/YgMNQIVgsY5mhtCTL3JneqdgYYyzwNXH/AVdORT42pU29hK080U1ByI
DjLSSypFBkhb9VaKoEcjIATLzhTyUc3GGufoBlSEQyBaU6woanKM4tL2K0n6VDJH
92R6XeZ3iuZ/vFqnyD8Klt/dHnxd1Cm1teQIgTqBLbqBw+ySkUAhicJ/E1UuOQiA
JoDQMNXWwpOfWNLlGlgBKsJ0Hsll5wuQcI+CvxMYDLg3SBJtRQzYqJurcvnELE1Z
mD5LzWpnm4zrqRz13u6tLOoMH3lOtOuy7R8TBnk6i01nuiRSUT7UcQvbz3I8OTCo
HmHb7+c/403Yk4uD3NVGGKME4KCvS4f0+LEAb4d19diyq07elf94tQaTS3V0GgFZ
yxPsxw/muqms90qV2JJQLh5cVlLR/ik0mp9Btb8NRmIVFuvctbi7Baxrxmqd5px5
7hIsKKdUjsPwQtHAKqW4t3uKglzKJVkUS4B4im+ZfFA=
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
oAPkM2KHNJlb87fFFmzvgNzk4By1DN7tGS/fw9UJAujePmav2APGBok1mHg50ql4
9aYkZWup4j5yQS3kwno7v5YgDvIJcKIIv/nJ+QychCqU6jq4HMmmahfMLfvmgKDk
ae9WCeHXijjq+vbqfcofN3E077KurX6hxYOxeGyXD966TwqSlpyob58ElBpJwGg/
FnmAXU6R36ASnTpLNvfx4LwZ7xMW2WEAiTzwubClhqiUURxdsD4qFPo2ePTL97dj
hr4kC4FAEL2UbUa90X+xvaODR14pqBFCx/8pS7CU2keM4YXb/i5owXskEU3yhDKo
CF3ER+h5zQRKUhodqtS9Jw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5040 )
`pragma protect data_block
JMwW49Uq0Fc6uFcczmt+o/stPdkr+f0/aKOspZV+HFpD+q/jzdcgHVeKwh1A9/LP
NjKF7OSa6fcu7mD8h/Ci1Cukivkwi6mdr26hiasiNkeizduFXhlcX7P9kcpuWoTt
liApD0PGfvkJPAcTMZ8Q++3cjgO1tkMdHaEIhcn4phcO1M+yTcRYCdNmfkBk/xlP
ZHF1Pj3/tNjGEINl9WTk+Xc6BsPrFckBwuF7b2ndnFUKoZqoh8yPGoX2c7kHUBh7
TJWtVB7Zrnp+djLaL01sfrGa/xgICLTDIT9SQrIIJrSmO1SgNJ3DRydOtEx2guz2
2jjad2OYI2wh60B3W1CaiXMUYl+PyiRsdFwtjlBA9KI14Pw6hcv+6nPMt0TBJGBl
aLMToG1x9sWgvN7P75W6gp60VMcraEeBbfm6bpSXJ1rvD2UZ+aVwQJHPzXLdCxmz
QbBkR4gyxIE6lmtBBmYOR864qWEYzrcqExZ6eO90AFxNOYYth0Oj9ea/Rzu3CBmA
4xujW/XDl4vdvhB1ldK4ZL6RuA1SbFeFwMkHNsK+a2b6QlJoMbynerFMkn6GwJR2
lUdoozj0o32jTp61Z0NV+WMP6zJfEUlgWyoIxN2NxwIX0neo6DMdpMRVeCRz2uIZ
x9CISOdxValGUM2QPeZvD8Hsh98tTfsf+SXKU8YnSGPtZNjQEc7kDmBKRYMKUT7A
qtZeOhRsBt1b5WwXp6mIKIM7hoXqH2oxfCF9GoA9r0exKb1GC+aMW5w7o9WV6y5/
bw+VVbgkn1O1E8gJc9Zmc3rZl9Mp7dpggBNS2rDbwiD6AaHvIZ562cgezssMLtuU
iPgqf3OHyO62faoETNfhq03kCDIQ6tQ6Cer6wS2/Q7NX8kKyV7LTiv+lEnZL//B+
PkYZUV/YixGY5BxboogQBsGTnqu7jreLWOPxNn2ZFKjvEMKEKevfB5A1O8xgv7fT
pOXFhLf2fN7plMI1VemBP/zJFrnGdk/rOWQ/ha6NO5vDnIkQyWk0uKwFmbRDwIzq
acOLuyxvr5iYo1733ehL1z9lVSXQC3fS6Rwev9sJwjNXc/5nCMZ5ehOwfOHDm6R9
VJU1isMYJp6fxHMUpXRZ9r869XrsGwwlkvYkl9dqZhxVuVhdU7vnFCIA2ISdckDY
2Etw8rMQgQ+8JueSsl9RxY5kzd8I66dSd6GOD1TRvmYkX+KThe787GYcSUq5WlSj
uDZyz8dvujBql2kswwy5CCOm2ykKwgLdTiy6reqizZaENyc/zAjQr+R/TFBIllMt
zGWN9GVaNzcXECuSiiO+TsvVyeVLO1BZvO34WE4RaUocKzLTfXgDllegRWQAllXF
sLhgIRgCbph8ShB3jezMIsn8KOfeU0UV2VvVC0DRDBWD0fgYdHoknNAoh3+w5ceY
2tM/1wLKd6fIfoN2/WHgpcSYKZ1urCLIUlVBANJ0SECeuOxg43Sul9gvVSZ9FuP0
i7QQZ+7xYUheMDOWiJBHsJRPfYEKNWLbbPIGDABgnYOyrd1U0VrhWVD2mUYCkjh6
C/TIC66fIoWCMt7y+6jATVsd9sfhvbi/k7BX0oNHTN+eaFopIcobJxYkzvygkM/2
Vb7mDi0fs8vaymqbT8Yb4CW3MJDEbbdUgcsqsh4863Gadn0oSnfqBrPZnHutwTM+
mtYve/490xOn04gWG/NkaTKjLaS+3R3/qX+npQ1ThrNO0Ud2ftVeM6gBfKrlmBaZ
dDFU4MZUeUKuqalr/c0gEl12c/kr2i8XYqGaffIc9CjjAODT+CbnE/oX7mCb0Ccg
FO3Q801TtXjSfUvNpUbf9Qb3RElkK6dxWSZLA0K0y9MaHWK6QXfL8+6x5KukSby7
1qkgNz6GnxiEsLXLOLw9M2kBuzZdYk+UdRthXfc8qPbTuEU0eLCFrSjyn3hGq4fN
ICIT8qyFanwW7PMA0wagSKFrFd3YjbdjVoVP+guKarnDqpUCLkfCjjQaevqoRAGw
HfKPFGjr5Cduk9bQ2i9Ded35w+DtGw5ZgMJHy3QeHwsE4KFws4BXf5STtbR8bjv7
8dvYFqF3/RbM0gCQo2BE9pHjToHPFva7hfVi/6rxUNQy5mWwKd29trlD8t30n+7k
1yg3aDua3EL6dfyonptA0NA+lI2bUu4xo1eX2rOQAHd5KzORQKwCKRG8T4Lh4EC2
bMwN7/RXRhvXBUz+n3MRaQR3eeRkomvHj3C4uM8VrELiS9mYTetndApnqjlk/fqQ
94BFeBfP6hQ5jZeewo3OtEL3R9Zc9zglnlt4BJG8hCLyk+jwlqRlIwCYO12UTTZe
wjys2nT5gv71J/lNtEfX7BPBQb5bN42KCFZGt7jntWKsuATdNHz6JG62jYcOtzwR
mRiHIQx8yLPwQkbvOht8iUimknwHgFAGfyzL8nOZzO3zPalb0WxDG5NO9i0DCT1h
iWVZ2k+tp5MiPbMHp6p+KFfkO36OpTPX1yPsdQ67HQ+Jljca4gqLwFNzPkP/1vWF
+EnAqbDzuv23c1mQCO7tSjKXo+UeomCwuMz0qi5txAJp6SRX/j+LU8MfqxltpUdI
ONfjgur7d0C5tDo8kN9YQgyhubYlyWE1gJxzNgrwHfh6VjnfcgLA7KTdQSuzXhVY
1R0eFgX+ZXtJAeBftFcQtp2M664tP6ArgjaVHlINJBXgDWe1Ccinz6y9toI+ZbWu
tXVH8rF7E1w7gFXLGt5635rH4PO7JP0+2lgvESfT4G/tF3eqjP62nFCNcg1cV6t/
AKHH+K5DnKHKW3Ka9g7H1WoYPrVTHyzGKtWvhzFE4sQNh++WBMTq/jl/laniyFqu
FNHdeHQUYoJWtyeh6KxyIJTD5PtaNRtewsSNhwscukBSUdHPzkU5WXSj6lYsWNp2
N6Mr/JOYZjeTloZB2zS6Ig0UA/0w3yzB5KXONyzGS4feNFiaDcFi+u44RID8ZD6V
j8S+/3FjXovf4IlY2S7OR9Iq2/MIHLYm6GATfOYpV4vZa+rb7bx6Xf4VnCHi8aUo
KiaodzXKL33r7FAxDi4SGP1uAlwxC8b/BlIsoDxqfMzLfty0uPE4KI0ztPpcXYw4
Y81RdXrQ99d2SA9Dq0z57LU0JDBzpGSKdYWXLyTD+raLTYrqynHHJlBa+Y2PRTL9
Zw4jaFg4epGeSA1QXz8gYu+19893mRLxrCTJVfLZyF1BSxSsqkYQT0oZTlBErMdu
PRpRKbBJatfFDROYuQ/E4D2ERiy3OaI/VhxTrBGgcIkk7CTu3xeZ80HOd9Occq1I
+s8i6FaheACTe4GiNmQ6naXf/PkoCEFa/6CpvtAN+KcfiBtrumXuKkL3IYdGqmbq
CTnr1T+YSlySqx1sqhJcQwZijpRy+DkJM9+Iykoxmp1G6Z37a6w7CAEkBp7MXh6P
bmHC8J+C73hdNLtpJzJim3M4E7EWm90AjYXaNVuWpyeOUifuXkdVCsQo0FYY2Hp8
ICf4rVtkmmm9eEoIrMIvdnVwzxAk1+4baIcZF/wy3sWoxb1jTB0BHfZ/EVcyov2d
mQb9j1Wc/uJPQAXpiYOI/sY7mc2ps63wBunWU0LoZUenN9A7xibN4cN7k0fzgbca
EWontGYyn24pvoZA5rBtvU+ZJMtqshY/HRi7X2HlKK3BWVqZMdrBwhgUtnBAf4ww
T7XAPxPUIgZEHxw9VCyEYOjxFZd4vHBK/OocDC2TTMxDW8umZd+aTJ3gS0cgEAQS
Aqr6yBqciVOWKYajoSyOhmdKS+yCeNXpqYLcRHq2U/wIBZtbXwNmpZoCUvCLwXRx
YQnP4jbYvbfgMIxpx+GG/Y+WNNEi41vITcx7wpD5qBgARRKJSmVqRMdYjcJiLc1A
GCutFE62bNdHs2eea1AWpEWomLqdXxsRf6ecynhXWAUJi46akk821cUf1wbViJpr
nVBKDrAMslUL4BfC6nkvT/sQwMfgaXNCo7nyemkzYgkDCH4ZVvf02j5wakL6pyDm
UUuQybdZoepRG9VzY3h8z+1llroaHVt8x0KnBghSeCFXIhF1XQmgNrV7KkJAx+wr
OQYMyImjO+EeRrqLsMsHnNFvy0px9eISTrrAlp1FGZcFu2P4YhQNmAq088hXOgzp
NC3nA8vJl/Ki7EKru8pX2NWDyya84Ft9SAnwjC6GhCP8Eetxvm0d0lvE387KIGWw
XE9BhC6FNb0fJu30woUWaZJ7i0z3Rmvc79ztytbHvCPG7iSUk6B8B0SUvDb4wzyT
z8vEEYBmW0E9BHh1O4XCxMiG8uptb1puZyUKd6IHyuHT53kSjWz2N0PrB19q0t01
oWdONmXXFJgW9DYJRJdmh7FDPuLRCnav2KcaQtSU8wjJqLxHADLUCI7GLvWZXWAb
Qv/d2jAZtY8JmXI/JcRGhPVICggSAY+NeBdiqLNT4VRp3NKhx7HwiuQnBXjl9d0l
cctG5NWvxrdMSzd52bL17KncNjF2t0g5USMLAFtzrq2ErQBdgQG18vZp9WFMV+9d
+J3xnjCfswIDe+9JqvrDcAwngmXODqDgQGZ18Unx75rg8nLT1XZzS1aS8CEVDhRv
ETgvL8dNaoKOM0fop8sCSfblQ9sZinMf28th4TYqPjIgToaiQIOWKMa2+fX6brFM
OJlmwT9UzqEbUm1D62MtVixbbe8+Vz29ArzMS/dSmxu0AKleL7DmQAQFkZxkiGFt
GGZVkjkoNgVxEaFOtzUAKEeEiGt3WwpvGcoK7g/kw/e4Jf83UM0OvC72gBmu17k8
cIW3AX12lT2G7OgEsoTToVYnrGWPQyxZvgNq1NGePchhVBqtctYdCeRX94VJEuIj
pBeBtOo249bPn2yMyqL26Qg2ZTDE1yZ+f5XxCWtG+Lq2nB7CdRg+HoYhEFa2nXEc
uNr+9pmPOXI/lkPsLGMg0W83OGKIUQxqnz2zJFAzFSAQQEnoPGT2kuS1cddDr3sf
lfrRTQc4sFigAmnDTd87iVc00ecmFhTdVvUyMD6e8leuoxnrK0Uok0Z7kaE7NsWD
kqB2qQjzAlVjg1l+dyDXtAxq6vGBRuvBPPTm3nHCngkFejN1/Ysy7+WcdUJ29ncg
okQJgeyDvSvmkRTTBY+25zRRTlO6bHoruaouwpR4Nx9wf5gDFmZwaesi1bIhYQQo
Z8FntEbDMf6Yf1/ilbUEkgHbU5oqN9ACZ5N4RvJlHEr+Z+wQLBOSgof44kfrOSev
/bsMG6tgOpHuT9VIoMypPREuAQ6xR9LiCqO08FnQHnazgHbWLpBH2NHwpMO+VWVH
dcVgHPSNgJA8rTjKC/jn4JWN/Mk8G1X3Iq+FOxIzzJFiVxBeOfIRHJii29xgsDmu
1yXB6Wk+hzJMNWiyGZJnJ4CEtmvCNx2HS68NnSIFeT+ednbSNLF2t9wqBynIOVHc
9EuUJ2rGVnZP2hLhBQpkvyRWZo99Edx3YvXJwtEIvaOqSr+F9cFfHb9SVZGewFjX
gbZyOV7hVWwZlxGgsWuOGbRnNDNUNERtfW3FGVpgaxt5bmIUHYK2HSnXGkXXGhsE
1dZxL7h/EaQyrr5UaFgS2Gz7mKYKhVqhtQsmW7ZqGF4OfK3Bt2s4m8R/Q078hTDL
Nhj4SzfsFpo48eco9lpDcJ1uRPP4YZ+IiyTRa+ywN4vhUqhfWNTNBhOHM322NkWq
SgyU1CUHlaBtuZivlyKRxWEBhl6NMEQbLw1WPfQ5OXzYlp97+sg1zwctUR6vvaQ8
bEqGOU4VII/oo9rnd+ehg5TN28wFdk96Uy7m6nfV1At1JXDEIjSPbV44/BOCUGaj
tDrw8wFAtP5yBn74k6g9QUBeXvmOXUlNEU8EV18QU4NTSugVrEBsDGIF+vI/wFnj
Rg5tdTIiNFjNxtu1s+OsaepM/AoSol+TKhhIzzyMORDku4wtFExE/cUAdQAjytQz
hRtPAP1iVTZoZ+u/WZh9QQkWl4nGEN8C5kUVpRjt//xxcv8iwCEFjWB8++6SUkPy
01LSRw1mWRn+sCBl+GuYRuvSPI9DGfYigSYhvOtfMqrP8hRqwRVvLta8u0vhjn70
VYcErK0oeIq0Eav3VIKIRu2MupSHVoXK0rn8VYNlqekQs6KmDA1fOB6Er4KlqQ5/
i3LMlr57W2lyetXZ+xecfusl21Fty+xjAj5FEhBuV3egXb8GXrRfpS72KxOznNzJ
qDdQ+H/n0t+C+mtGqTvfu/KYsWg2DkTMlFR244WoyX0t8hvNe+H/w0fekiuj6CLN
G6MouzsO5D4ninYhRc858iu+d1Y2sn3hX+7mNIi2AEzyOIOtDIta1hq04EQnqzOf
zErCkm7lH0JVSG/nRdkhIalA0mVTNMKQYWYnKQjNK4ekNGq/Rv22HJdlXR+R6/9W
FslJ6F8fROEEQ8IE6bdEGqZrGbCMniznCfq9ZhIxAjZI1G3XRFsY8J/VQs99pyTV
DS1q6+UTMQVblsyM090nF9OPlxLqSQ6o/5mdpi6+YCoVM2gkvLKk0+F9VkOKEIrH
C9lo2BWReXElUsW4wssD3HdjqWPRsLd640dbbavucOg5U5IGvpQR6Sf90Q+JJKBV
pfz1vcCbdq3GnlMpL2CFv9WiWmzuOEovXxNb28B614tHLa4ep2+BNOBraDa44UtC
vnDtGAswb/dHF1I4LdLji8POQG8hqXP1HMnS9eC+ub+7GsVsc3P6ovqNgjZFJJUP
p97VdVNoIsZX9v7pd/VQJpOXvMys45O3AxzjoqfHbOd/SkppTixGwYnokrGZh+RR
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
MB0G3Yzb1/1Px0LlOSdUiew52Q3l+zclKyvkS/IqjhytkiepEHjHi1gCUsyDgXF7
ivGodueh3qopKn4//gnf9GItwEIbxePbK3bgBJIleD6arvrgLLDxfXDOExpd0oQb
dc88AAnceVZEG9cbJYVMWUhl2DqHECi4c0p9do/DaBKf2PXMdz2I6FQC1F/Gdsme
hJXqqRJXP8y3v7bu2jmoT5EBle0o4P90CimRrnd2i/Pbb0EOxn4RSZQbNsNNBN4K
wfooCLHTRNwy52xH8JyaGnii1Xx4irwTGR0hyeDzvd2/8pKMR8R/bxmL1n9r2+F9
4jhZ0IFWB1tYFLzUJONZsg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2624 )
`pragma protect data_block
nlkE+0/Yk/HcBEWumm/MdWWXuJs4ezsTYId0d0a+fwKkjOABwrHIcXjVfwwiXBxZ
wEFyuoqyOxpOvQgvM/ip09jf7uSZOFnWhyG0eOqDbVu9UYpLatBQrDek7EktpDhg
73ogMeFMQ/69E0UIgYl+tSBvh/v0mSIRObIZD/ILXX1uY5++0FrQ5PNTHZR6UjPt
jknjihvviprLPtiTiscmEW4QxZ8OdV5uFmgQHjm2puRiaRiAX6ZVSx+Ya44Hlpsj
5c5KgartuXWgI1xtanvYjdcNY0oc95j98jg7YwhqueSOJvQUofnXjjlVE0IHaYBR
19G/TL+73W8XZ+V5DqthDY/dKzhaaq8jFP1WD4jCoYSNLfd6ivRLJGnoRxuK8ePS
zWo9UVpJuSpU8d1d5CK3nJSx0lcBbQ1qqr86WQmRfFN2VZ5YXe092TgrkhKqAGEx
rdnIRoeyfLE3WFOmzNeKBIjfH1SGCPjwxBJKxCjwL6BeAeChsMdACZ75duHndMgc
0gT6q10LzBbt777Yw5YNgscO2zyxVmH0SkTlzbimVGGb/kWI+hZ4uQfhVew+2T1J
fYqhV23Jpq1r1VV/Z8f04hWpfY0Jk3Mbai+Gkva+Gjx9cakP4sqV4+4qUbgJ5sa2
N3Ls+LUGV1rArKOppbN1mbtJ8EAQiaK1xPXw2fSpwuP2ydN+HsRvXtyZ7y4iasOy
5doPW2JF8rZhafgHLpDQGy0tIllhE8eCiOGvjr4njzZcc3HtILKEM1A815BWit8B
FZfQA2Zu6mAAYFumCJUkqTWwNH03JQoVmKZueAG8GREPFd77jWrLAkGNp4f0QLT7
Q0odFNYRWhWQWwmhVa204iUH80bRpyNr+aWP6Y927viRl0DmL1UrVuTh0kIgvo+A
oGmqYzvW5QWQm7Cpbxund5Lfmgpnuzm2WDe3dKFINOzFM5t1DtyBf4JyAlMWSKdL
ZPLaaa0Z0w6MhiYygamlyHHLIAmRfbpPLw6fTZYbUViCRfLm5Pxt1CJb9QBBKYDx
etbsI4Zwwz/8iPyN5FpKchN+og1irCST/xljmg5mPNLcvguHANMpHOkWiRAUBMVi
puZRXoqP32E3mK2Z8GpnE4vxMbANXGvcOy56/N03+auvSP554y4nzUH1K5P+/ich
LzkVdRO/WbfVgPjJ25zlzrYVVOBIDeTITIwxcbDNyZZXPKF+ZAT+Crpb5Ni1tB7b
zYodutJSqR5qKpnM314ky5QKk1wXQ8ZlpMWPLZIvdSozg7l7yylCFGyGqbo01ooR
5A+lQ9bCQSqQ/YUJPIbvgenFilpl8AnHD0j9FzygRvbWAB7uvr4McN8u2ftANdPH
YVv12LV9ELre0kUXDpjd66D1vjRYbrD2L0wYj13M5ijxc1WfW/2hnE76gM1hDt8Y
NcjH5vM4zaOjxfgXbTGQoGANun26Ip9W9Bnr+TeTBwXhGjmlpe8pSE1SbzvqDfWQ
6SEU79TaKHO5AJ6hx0XO0flTlxiyvK5wUx0izcZOlFT6TrsHA5+UMuU7BzdsCbXq
sBbUrTNo6WJATgpqEs7/gIIpn0nqzkyzqZQmKhpKjwQQug/jiGM5KXAvqmJeeV1i
E9LNtEiAveFZCGFR6cGffiDqZH9XMls8ynWcoCtuy6jHLMwMt25vv3wXg7Pf+psO
0Tb3stX4Z1eY0eyyWuucOif2DcItuARSTRQqdR8fuVl+lz535YgF/609wAYF8xrH
Fw3TUFyqcIyiwgxgl1zjKKUXq4pn6jen/km63iVW/s7wypFzZNCY2AmEUP5dn39w
SjxZ4K3B28fMfw9vAWERZGjvTBX8IC60JUQhc1/tCpvsdzrWm/fD1d/x0c1VhnBg
PntoqA1TBchspwCTaG1KDPm8/fPVxCr69LgreKYUYcuBTKtDJI7IXZIobg2bT5kq
JOTL7uJrWQswrgMrCUqH8w9N8QEMG89l1VoEOFbhpX38VkjWjwgc035RDo+3FLa0
+kiW5NsPVicntmsi0koszgtwcAt0+Tw8PtGoGUzOums0WUTOEzuMf+0LSYCLHFJj
xRmFkp6b2erYL1d0nSzgNSGn86v99bnXnz6c6ZfZ/zCEiZvdRVRTQ70FBvf61BVy
YCcHjX7u3jRyjiXJhtWr7UQj/RVFesk6/n47x9FlBWj0d8tipWQ3nu2bXZ1D/8PW
qbklCMgMyh/CyvT+dyMDKHeE78FqsJ2Om/+E6yiwrgZbwYp+4Ijf2NvAfrJt4/v0
pyVKnrxJ0ptPuQTg3j7Z+x4BcE0pVbpRXAIVM1vJ+55nbCppJJpBGItjH6P0XvGY
wjrtCmjRH+an83uhTYLCCog69XvmVHkw+7UtJ2oR0cYkIL0yxagJUr2TVtKd/zGM
SxVqTBxfCuwOPCtytVjZNl8KP4Fn5TIrHUBAN838/KDtS/VbYIRlhXUBEcE/vakP
VoxjocpqTLx1YEQREZvqSlJqL4YyVGHgtDlpLALgiRKKOk/Ipfgn7Gy6P9l+63td
StfuUdDPl235uS8+PalbQFdyT1VqQL21s6kZcCmaF50wHdsYT4nSZKH2vwcvxs1w
pPYMVAt70HaiPh0sMbG/YKj1wLfujfWCDrY8B8KRtIEwMOIDBd38iBPKoo1AC4s5
mZePBMDLagHgYr/3GAsSqpGqH+i2ZHQ9JYgpNy3IYnYsJBXBy0IBij6E1c/qx50K
FtH2m0bquYeCpl/C+wTaZe+pEJezXb6G1mEv1YlyLq2pkCFSQ8MWGsqWTk5b5OHW
Vx4g13ID4wOC1PxePwXlldVhw/Z0CPOK2EncwLXV5LZ4sfELtTY0crnjq3Oc1gx8
kYVgN3y8LXhUs9xXQxgvEl3wEpviMHaksDJ5GmjJw8M5ZEQpTCiXUIWK4Q2EbBhz
kuLlGzLMolv3DvCTTbZVnxMS1XZ0Y3enkrn2C7XWnmBeY51629JPrzMi09j11MlG
b38LVFufp1Mq7kW7CgVnmRn32DWdDCJvRpYNWmhqCh6DMUS3y8wRJnU/Lx1P4KsU
KbDWOX21UM+3u1ZNd+eVuQw+KGxPHi4HExSg/ahKYGNKM+eW5X8K4JYglCFiWF1i
e+uScOO0hXlJCoI/cJ9u/GQFquLYZhubHoRyiUH1h5xypjyGIG/QcxnlCE5K1cBF
iWQ6BjYD2fD6MpW55oknOYf1COZQoHvyIMl3Ev6PxDQ5Q9WV6vbgerQ+fCjuK+X1
PKsr34Z0zD/ZKG8h39EVohvGNsrc58KBf+rnTwBxhH0EP24wg8UsrPoePNI+Vop3
MiErOw5Q4CZJn4oqc5OcIDKUNVx+mDmSmiVqHdHPh+wHaIee7i2xDBCnFkbEP711
0CNqMWpznVAzpsqjIvJuq8PabkL66yfUpYBBToYjjOIMxSoEt9l8NRXKtW1ikGNS
FUnaDFmuidxO1rSqY5WFMhTodFSueRASqn9UtzkkHpvS8ZShOMm8Ho7xDwpUVuTD
kBbaXOd9I5w40co7qly3vIQfrYcXGmgrXw4VsQwT5eI=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LGJ6iBQ80N47vdxM0RQ5lP7Uyw5k71jMXBe8ROQQ42WHfiYVc+LuiEeFr3aMsdDR
imEH1OL97I2HOQpDZEL3ciyi95YPxDjeJeUR24LEJHyYZaA9ReLnbiiki5N4D9IH
CGPjLycTaztfTkkAydGfEAR5FH3Ln3e+0NSLjRqkC+wT5lqNzLKUnJYwA8JtA/VD
Z3rPVDr5WOo8Bm2enNUYbYyawAp2aC7K/Sppe9dYLTzI55Zmd+Cbgn7hUaGyWz/M
U14nz72zWJL+JUx3fmqCdYyZixHyvOf/Z3LQfHqqnHRbYl1GkAcs3GrClKFtSm9/
CCX1b1DjF6pXo9KPFLOHBg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 784 )
`pragma protect data_block
+p0YjQhFP+GS6Ed4JanumJTyKxx2Fcz2QvT3GRi4XHwuwppq1lF+BE3ahp+Mkw66
OMpjHD4njtsq4zMoTyqZvSLTcXlJUysqV2VPEm3bliwRHYqmHyoJ/BWui0AJBfPv
71xVb2ReOZkl4AkZUiSdExEiL9A0/HD7/Rdd2eSlNkjs0eXzB1OYnwTK6A2kjC5V
c73C5cmdJKGIciikZHAlPmdJ013Dg+Kkg+I0ig72TE1KsjIoDJYMuGGOwJOsUDgN
U1jUqTsH5vBooK1450qBcoEnY3ifWS/+89WAMIRTmbAbuxoNChEei8BqsLtrQvT3
1JTCPpPZSVR+HYTAcZ8eAxN4of7XHpzW+b5wLqKKQZ4kNqR15rEqHUwJLOaHvIAE
x6uEOUm7qlghIIKGxaqbtAWWOmgko64zXkMV/Jt5eMlK1K088pThsMh2gR3C9dXo
is44ThFLy3YQx7ld/0ceqRxkruwrvqGQ/+/4ovgo16MJhmmDz6JVpr73bCipTZHq
auuA5lcBTI9tRjwEDUUta1jX+AfVfoeGJIxsn7TGV7RQYRlU34r3+ras4ZCkOlzD
q2fP/nXoDARI+Pk0RCo6cg4yGCLLcsQOTJ29JiXZbmRCyqq9kw03d13VCVZEKyuG
B7Q2ukEKgFhv8w/VWGlOJ8OFbluvDQzZstmGkPf7T1alo0He9chpkMecARbNJHWZ
pIyypoCDDuJbqobL2h6BYWlxx1pifBGheKAmMNBvk/RrvGIimeK4I62YcCV/ZbaR
idPm9ASLLdDZS6j+11k67VnLLIK9pPfzzrp+Om9QkiVVS5Uy2Oz7L7bwX9AQKL4J
eO3dWgLLlajKJ7aY27JvNmY/UgfMYYmuB6dMgDWe4ng4o8XcA0OOkHN7vR0PdtOY
hbSmzu4ar67W8gu8FDrJNiZC9zDUmjqY1VkIVCKkYuibkh3E+RhbFYHzyiLhlfiZ
ij5BtxkOuHuy4f/AurG7JihVaI+RZug7Ym3t1xpv4qdZFesUFZv6L/7T/WTtsRym
newv/laW2akPKwoOHeBolA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cxGtwFn7oVkIKiir4xZU1AI9p5vSB9OUZSDF0uoDr8HoIWy2G9AhaTkhFVXHlxME
u7TEb3LWH/oa1qtX7ER1TtFW9G7x1VNCwtXINOGs0mpCZlBVNu29UwZqUMgrZM+V
ZOKzZsF8hAbRdo4U1V6/o+RsqFaXTMGQHKhgEjvFMqJyn/RA+KXydu5Ip5ZqOiLW
20VDnPCKj8D81soq1SmB95Tujdc0H+Ks1mQ2gqfcNArYADSqld5Vde92S0ICyKcC
aagQa+XRPOez5cySzn3l742p2hJwAI5KB97SNMfT/U6yQxecNCwjMkK9yXelfuoW
kFCts2Ps/bH0UWSWq5hiQg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
1lRTvs1URAQxSvTZwBBU2iWBkR7NxdAw2AVGR1MfKm1iJgyHh5AVR2LVHqlL7/0c
foDw0hc1z/G9Fe9A8M+fdEUEUoz355TZMiy2I48deg2YsI5YtV3i5XzpGlRRZEaK
i/zTFODz/V08pfi/mOaxf3tD4s+SgZFFeTAdSavvWgTm1OCb3FVgW0synszr6p0z
LYiWcjf/8aJWlb3XymgoL4FRUJymjEM/Nsw/pxh0XW4G7qeZLGicD9QG5tILBrjT
03RXSmimB1tsKqs3x7usLlu7v23Lks0hoY3ch+O3D6xedolua8SmZjwHS19xLVbo
l7olWgxoQF6kDQE3jQk6YODgf4Jz+1/4bXAAMaP3Tkm7xxngIdQhf6MKA9Vm7j4N
iddYkRUMVRwB9LWMNfocW1oVbiH0Flwyu1BOVx8aUvMNa2BBuV7O1+ShTNpW8wUv
ZuXUaODFDbU4wFgldB2qDP9mkIrTZl11VwQ9uHV4C64F8AcfLPhL+JsySiVK9vy9
DGA/NUEXhKgdwcHrY6bfd3qsM97Im/i4sj8RmLPGeDc46tlRE8QV+2394pMgVLjB
pfKekCQf7E7BDA5bHeTJAyJCH8e4PchGIJM6p/aLR2Wd1NaRmnBoqmogk+XN5y80
CUnRVxnkGdSv2CejHH7PjyXkbNZsFsHE/HLh/jELWKh/ms97TBQWNpailnZCeakQ
JSsKPPFy1e1hpYFAE8TwdV+Lb1O5NM2kQGoVemXoG49fz3Prq7MzCsMrcS54mbXW
77G1+dbtvydT16+WtlS7sFzTOLx25txLf1mvt5FnGCJZth7CgpawP27znuBRMayW
8qlQO1NNQimMZ4DR8LqFptFKi5HrRBX1fWECToRQfqkQeKIiq8cSJdutYyYMMr87
C/8+LLFbiSNAN2Ozs7fXIPDmpMQG5Tlqezuja3XYaU8=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gEJH1bfgZCgqQN4SMWM8uNunDSZjHZ/xIAxRhjhL9/yMWbXL+1QxX0qg8TqTaaxG
goTskZ64xEX2DCH7NywnT+BXz9BaFLMqEcBITDzTH1cWC7HGH0MwfoDkvgvFGi5s
/5r3o88kzbJXcDiQY3tSs7OwkotRWDhkVVsbxIAC1w+sUSafmHGm/f1Q+pATDL6+
TQ3h0rctHYWIIW8V9HgmaC3eupH/Y/wGhPCyJX4ybdgJlBpDwPBFLDEI7ByPSvVq
QqIwLRIO6FAW7Z5qwK9eOiy26D01sipJyObEmKT+TIeRUw0NoUGhAMgP4d9wu8kN
QAMO5Dz2z3g5mKxzsqc4yA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1792 )
`pragma protect data_block
Vt5xLUgpOY0zRHmH/B56kBdatz6InSnXm4mN43RwmsJM06Z2W78t/na0xq+OpVz7
0U9GFbfPHtGQEw3nx0gkjdkBTiyQFz4HPeaCwcV5sDphJEq1jOKLT1hzm+QvqaeO
Fo5eI7GR/pIIi9rMs2faGtfKzwuN4RuHauQpbzxwzmF1GVQRhzL03cFmEockEskK
DCUubZuaTH3vpQqdLAyn3SQGH4zQ+7+f+wxr7gct9JzV2o4hT6/mxuZ27LQHYgnG
15NL0kR/PEncOHOCeEt2zxyiMD2LwAyhnLgSfAlmoMm4NzMZDdgDX1ySY9J86G13
bDDFoo4BaYoBVPBYi3XkAVL2Dlo+F3jIcSJw3dMr1Dw4aKjivWcbbl7lddRmXU8J
mWuUEtcqz0M9SbXeAc2g5ye7l4BuqNw5GNY05BT8TlLXJ4TeVuyHAMrPuX6EvbhQ
VGA0xPOBLImCA4nhlZ9DELi0Idq0Yxqnup2v19T9Wk9cxHTuIT+MPlUNa/iuGekG
q3htR4Ctdcig3ndb3ZjVPPv9hpmKS68io/9wCJIhriNYDuhGvycea0ntsnJ8KU6A
s8aDRoIRjUJrNJATDKTX3EmB1lTyrQG39DdbXDcebLoJz566Lhtmv9dkOQGEq+x5
ZvvvyNoqCImNB+qrRg5Vvb7vCPeU3o3Raf7qM7FDlBuVC2xMYOzAxgWAd340dbXL
CiKMfCRI7n/iGiZYyJ6hvcTVU2OR9PUc1gzZ8E2+LLuRwzIdejGskXpj9X2FJISF
Gnn6HmALYFE8rsXz+UclCwo2ACpa+Q4pYy3TBINMUNF2mhmD+eAe4BTGJi0+Kbim
onw/0AxEDYJD1+6daGPLSIXoWKG+Vle76VkRXlSEHr4Zm908U79EfScAkHcvnS/j
eLJ6b9cZj6jk9bvWKamPnFsnoeJwzwR3Xjn7Ln1+XGvQYugXwYhW8gET9UL73Yoc
EnwBqLjuaLOTApoJSZHp9bqvsbeiCB8TbHy+wqj/KD+i8aHRpbP6GcmTvEnysy7l
Cf1Rc+lWbNPEyb3Sud+eEQ/HkITCaJFQ0vpFI4/DWgD3dNsiB+X9RE1IW438ysI/
jSYN3QOk37MPH6CEVGs+AenV/ROIzxF8uAGMQRccbdTukhTmL41PjAPwzHz77uF9
MwznRAlrmc9pMS6Eezi0AGssfIoTmQbGn7GtRloeSPmlt9phxO84gXUqZmrvEjz8
nYcxZ7Rmzx/B8XjmEV2F+3J54zNaPuTw+H7lC47LRwtcrEk2oOlIjP3sYP1VfLPM
qPgIrrVjl4S/7RyAs7ZMqsHVx3IbEA05oq7mTUaJoN9vZXB/hWU/Q8yEVOJVr+HO
ZYFnBeAphWj+cKcDqnmfwa3W1Ab0/7Ru+j2j91QI0tkO1yCyQ3XUfVk16NXXoRRx
fejrANvUQA5oYHQXikb0wl49n1q47vjqNgGMbpVpia7LNgZ3pJqr3NX2OuBC6NCH
lMmVkRKsL4qvDncbLcqmzVD4S9k994vxDXjy5aszMuhaeVh95l3S8Vsh8yE40pUy
xTOLC6NKr8cTn0paxSps1b0iyVxKfsQyXCPa2ZnWWe3vcwsRWTeo/dy/mb9U6Qt1
8rMLt3k9SQ+0vc1HPNQ9THNZEhZNUVnzXC59ZbSpGIM84y2fR6NdwljvO0vBuxyM
MpS/v3ip3uQDBLE2yQMzZKDrA3zD2oLbRc//ai7Imd51svElwI1A+6S0gzkBjnuM
l1AeKRCBRAPrM42fT35c2mI8tQHalAPCGj7NQVaaQ70ZLcwr/yVl4GXUbfbBr41X
AjvN7NRVg1GOxNPNLqzyhVombEklmO3gHPx0d5wtfdXfHSqFZL++dwVwwpvZ1cOz
t0h+vhjL4yBYTscdYoRz+Wmm0BM7JWkZiIkprV/iYrLWanOJozkh39K53btADehJ
kGrqkmKoVT3tzfDw9sJMnrzm64NiUnxYyjkJvvJ2IucIxDLrFTK75c7+h7kTVRXn
pu4xE/ulfpRGuF6QDFGSwlNG2WD44K0GgIV4jppJhb7YiuClyUN4OsN658gU1Caz
JvHxGUtvOVIc7f3EUm1xyEpu23ht1DIj7XgGN+3T2ECoPMpK4mHoyf97nIMDC0Nw
0hGMr9odOWyozpss5vzAGq3XNq37NzyMWVsXjphypQIAP3jhHrhw8hzfwttM7dEk
voVk6o+hzyVgR+SG9rVvJTqmlJg7Ac97rwduuR8JO/cWZ9H6q4iDXl9j+kVZ18La
crKw1GFNkxb8s61cOJdLohKHfGfxChzKFdsf+VLwSOJgV36m2RRC5JIhzvNTyqwA
/T5urkLRn3+XpLxJdASpfKc2oeqgf41JL6dDcOC2yDNKR3P+dIc1u0Q1KylmekYs
PBMQLuDVahiSUyW/EwATsA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nT/evmSZNC4SzAEE6oa5dffpg2F9IJ0pnxrNNeNcL4Zl9a4Q7EKLH+Xd6suPEEdw
PKTyecEQDl2IExIng+m398xJetdCeMY0sTLt4WvCxssfAYHLhzLWaegoowEWqFcR
/MvhjPDfVqmCLBl7JU0OE9WD33FSywb9QtU72Zuzly0+TyztsQYgjdF1eS7hCwbT
T+KqenLmXQ+KzaxK54aE2k0xFfHlb1Qo0HYrJef5JBy7QU4YQkUemDbieZu+lNe9
EYB6vP52S1k5gFoc9/Q0LcxGtMJLEvI4wHqKvxRnP1pucwaGZ6Vl2PXZlTUacjk4
0b7eUr6kn4BGnxRqqPzPpg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 38464 )
`pragma protect data_block
66L/AvmzA2tdP2WOCUYy0OduUGX7Sk0AqBcIHSsHJYAK9dZLEUEnWfFIooHlglPv
yQwS8+zeRD2YC3hgA/iwIzTPoJgyxFUM3zPTOQ1883DnyRFYM3gHPigQl4S/Uj8q
XfiktEZqjIp83FoZbm/QWr+wV6wO/KWtb8aDqAU/Y3nivGkGHH4EByMEu7HruxUf
w+g4Yhnp40bIskjjDN+x8u2V6+mcBAWcSjv4zhlxpxoEF30GBJZiluhMM9mDcZeF
OWI7e/UDIx7FMr8NBtKNWfFvoZc4USYvZn1jqir2PAZkc4KRdhkdOILmutIauHkD
DWyVm+DB82ttA3VDNLM0SyuRTMvpHCO1lPTHJ3+biR8Up7fUR9MzLf5jbYKqkd0E
G7PIwivdeklzEg6TYMtmmUF2nXYGYYIR/FcBTELZdi6XXC4FZaPzTs9JrZysRm7I
rV2FQTyR5vdUziKVI0waF4hcmKSCqhlpvQ5iin4NwdR6pCilkF/rKue/AN8WB2T3
87NqORZouvBSUJnT9nyeTQZFwZRitlhOm7KKhMPaM07F+aDXpYL+0Q9QuNVHeY/a
zD6+W7f/vPYW0ThUJL1zZWGIH9X+kdm5j6yp64HZo9+sskLIls18zjfyiinkQ2e0
X0jxyI2krYJWa14+0LK60o+sGGXoxWW26Fj1LnGZ2XTgX7zCeXMDG3Yccm4ARqcZ
ym05Eub5LF4JY7zBwk8e7upUX8dVt4R/Xo6lu8b50M3fNJRtiB2jdP8obmAQo8lH
TaimQoXJzQSgaB+lYcOqSClPqBndorVbdGbwYLmjp8lpaUejrdDHacibBiQFyvaX
C1r5jY8N2ChHJHD6z56Ix/UrnOavmKXYmJAu1PahcRIVZGdeZeSgE228wm3/vWBb
xBwjebM+6K6pJ2PYjCYMtArjnyK8J/sCPSJVML5Gt2N83+nmRfoINcl/PxtNzAa5
tjgfQRMe6/xYPoi3tU2tiwgBdNSPJKlHUTPCvrSYUZFRwFsOBcUGoVK3yRoS/TY8
1srbIao9tB4PJ5OKzG54Xh56iDVy678gaTm3ua6O0FOOz1at9sqPPDrEkjeg9lNc
9pS21brknTRxOM6LK4/J8Lzf/qCjI8qCgoPpm/nP7N9qTcOH3OhfzbL+sy9+Q5rb
amlA3Vp+r3CHqSSbtnkJXKUr5xXZVxI6Y8g9QH/ZH3x2h2BOSopN2/ijyAaNyPZf
Jv3kd35cyHv437he92TmLJm7NWvmOiV6/A9LGYSgN6OaDwyNfnX68F3XuSSIFvI3
P+4N2mgSCDENj7I/f4jfEiesRURUS8e/BaFB42QGJedtJABCUY4mM/1JZOyLZFkL
mF78AIqdnxiKvN7e0VLLUgvG7soZVmZihg5LJGw3AmrMOVNkAYox7jSiXw8TlZsZ
bBpeiikIs/2MbcF/cRT/BLHgBWHp+7BWlJwWVtHEMLvjtn5gtUvG3fiSdhoLvhlE
HIujN2rWSMrfId6Y9JI/cAy0H/o/F+Yux3vxDgfUUKmxMD77kyEeekudigP4H+V9
ljH+r2/4xc2QqcohMTJmub8eUcyzMn40Z1RIvUh63cx0Ueqy7X15GLf9C4JYLLd1
bD/IKaDZTIEZoyuK/a1/P5MO1M5sWVxa/zkIzw+KNyL7hApN8iRJAHOLwOhbYmfL
qAqB0YFNeNPfSe1NsuwMsJGO7w40mVyZbMdx5aPukqVkDxuDefn7Io9S9Oo70FUT
L0OVONy6joz6kbRY6z0mM47nuI/656VJlE6ISbG8YXmDx8Mw0Wcww6TXo9GiRFVK
PTdnunkin8jqdmEugILdRz55F/rq9UhAJKZouFfDbuahIpB0O1s2kSEEsMRVzhXR
3jmD0pE5GuXPJI0qcpRa/osJJPegouF2peVp4v3TG2LRI3YL5FVEArO+TcxZN1FA
mnLGcgUXPB8n7HGQUVD1DBCSUEm6TRSRchCDgnJNq4I7GyxYw5Xn/AtGWxiXQ+0k
i7ay995t7jcUWpUxhBzgu1zZLmr6lnqXwRYNsw7McBlihufuPuF0BXmF/DC509hW
nTE8qjxQGRg26+fWM3bLh6D5j/DadgSPHmLclXPHFcaKnRDzqnmctBgYgadNswEk
L6OSX0wqj+CPQQQPnADXNPO+T5M8KLH1khGYuov3Euj4zVD8w+mDU1qxunsCgYuW
sDrMQHrzOWyyIpwH0grWsh5kVdwaRDviU4OXWDcDT7lf+7jw2/QvUsmGsZU7CfBj
og/s7ueGGjuFW1QEqOSdFdSlJTI0hTLBGgTYXOprpDlE2J3elxozGHYoxMTpI7hy
3+D0CRTpLqo1AJwZXI+e1GSCcjPvVYGTlTuXxz6WAAIxw2uWREOOjGdDhAQyA0Ce
2Qp5dWdGKHrbEnLvW5pWZK70nLiqJdCjAfYaH39yIgGQtzru7fAIKDIaSwzvprRg
WgywY8hztuETLzcpo8weK1yh151oBOz9sZT3xIHkJGijhb7ZCjxpl1I9bUZX9gHb
8H0T2PP8QaNazLRfyYDHS6VlCalIRE3uao9Sa7dztEI1td0uDeP7aPBqBzxOJM4L
5uKbqufYeOwTRrn8ycWvDw6AwQvxaseLkrnAhWuLD64dgIbHSA9WMzTJD0TJLssF
pgEXczK1l3TxRDS2eSOv3Cz2KOobRcb30V426Zskc5l4GY96p60+rE7twfBD7iJK
rIb8013slHsBNdGKlnxMUV0pgwS5DFzzfFhAbNmlAZ+o6I+ZlBDNIwS8pZfqkCFS
VQF0NdxAd/6TDkNL3Pj9kpWQg1N1zKbsI9rPknnGa4bnb8dT/x9wQcFo9kzLHwnA
9DuxGM2jJ9oyy74u4AIyV88XSXC3YYfDcAbMWaUkXw1PoCw6EaNQJLK0H58P5oX1
wRTsyCiqEZT21nFJ4pExass2xeizgkut6MqSzQ9qF7c5oWxaOrcitHQ0fBW7s6vu
UoYTBWYuEKtgBR9eghOun1CdUW+QloTcCA3+Eo50zZcbw5etPCaWgMmGMcxZrIZs
snjDGTeuaGFLAcnMntKRSKhvUzEIB2qWJ+WGgcldthB0Wmq8baoEGJdU/FNi+btr
Pd/7w/J9n2kbPvAafNwhF/6IVIa/9qN9bVfPNwpEvfK6K6NzPvTPO+fIr2aoi7ku
UHy8N4jmhbBtp07oMpXKdWQBbJqt19muvU1Oi1gd+13hkNpL+uv9dPnj9oGcAhdk
CeD4CQcsO2QweiRpTDOsnTb663S2e7+uq3qDQWebMh2fa2FMJYXftuQOVHPxenPJ
pJqKa/TDX/UGjGwD6t8XupUsfXUoX+q4lIRJ4EBmCboD3IjusViellt9+Ti55gY3
d0WefvgYOOVMNslyCstRZJ5mgkziiHgRlLvMmvSj3UtsE3j+Dm24CgXU6iBvcX1g
NpxF3+l0huSOOPO4GsSroq4FniL59Aey2ICcdce5kJlSoPXyXKoazj3VHLAuXO3N
5ml27rf1+0+dnX6g7ZIrhVeGiy3cfmpNNipCYPBGiaEvfXAiF1GUenUDV3GZ4i2x
a+ARUjIMLATZ5cannwPVIz5G+4C6YVZuiKyMrwNbN+94evFvEHbJAe56X+pS1pl9
aGyQB4lJ5+7xGbm6jivdHcSjwuqCfA7yZ1Q+CB7w8X0Qg+QLg9EHtieMQW/EhWHw
UhiHB8p+U7BZBV6/KVh44VY0LVy2JkKUFYBUOvsR5oQsuOU8onaq9PnSP1BLsBnc
NEqSOEgvDsnxc1wtYBcwttpxqbOuKGNAMiWyH5pweLf3mGSJCDeq/JgZsc6OI2pT
Sj308c3o5XO5GhteS6POhDbqSU88ccUfaF4wpJ43qWpraAlBvoYabc9mwfOFwPTO
ztkNSgwnzS7kKSMpLyGn6sVTx7MRXmg73IIJCalCbFrE9eP5Wm+D/PGTQPwNQ1cO
PpWq3kLCqhJKFi1yYreFGl2h6qM5uTyWZRFDyWhKXwSthucNaHq/ABTqqHYyEbsh
2wsfb3DTaRzqsZVbR8+5TKwzR+XPEw4nxKDz7vbL4xoJf0RN4N3JWGBf8JArRsvp
TVPpIh/4ob6+BFagfhm1aCkE+6v0M7kw1KD3Kn9Qqjo4tjAsvQwklGyj1DfUZlEp
TeTuq5+Gf+0go/fdQY+bok3oCtSV8lnbhVWlOokz8OOcqiMZuaUHw5WDFIaCVQD0
dnE/Z3daeAX/d8fdzZdwT+xYQpR9gjZKw4jajyL5/toyMAOfx+e/AA/t/Lx4bOcv
dLMOUV7DCO6FGOm7QGivQKisWowm4UZjoUoOl36nLE/o90ugPwhuV9kvEUarY1LF
gXfoHJsI18j06ZNEcn5RJlWs25VGh26hsV68sPCvoDIVLRtsS/tDM4pV7EvB4WUG
zlV9CN8hpmU1lqOz0om+LoOLrpDi20xzaYp23t9Tt43KT2uVNZzkq2d2+++g0tor
P39PJE3MNTWCTnuBVS8V9Vp5R1qa0k4K4nCEcZm6VtqZOSBg1bck7+dLlnbk3llC
Mt5XXRbf9izx6kldQ/SHwpwEEnILoFzKXCgQjlhPVVLavooPevlOI2O3saYfQGDY
UWcT+TetsOX1eOFW9fbWqwwZZ6H2xzhdnewiaOMW+aTmIFuhpA/TCAd4JB6y5W1x
3RmbFrsgg4w1iaZdPRUhOmdcLuAZhV1akllyTtkaNJG0RAp6vQ3B9xX9ww8YOIdC
Ryuvqz4G/uXln7ZdK3IR1WJBwq/QixRHl3XUjrtUuqXW0i3Gnb/U72onn8GtFV3B
OuJYcoBn1AhsQlFHC8Hh1Zlmtyx3UwcyNvlyvSu91fDc3x7lvEKIOLA1n8Gdr5FQ
9+/IcuoLaJXxAT81cXc6GxCgZ3iR1aK+8GPdtG+onB7izEBthq3TVHLMYC/5oBku
FkFKBhJ5lsMkW/0EtdFvBd0j6W70C2tC0DNxTrbcUDWm0T9L2bYFB4aaUHAaLFpm
CYF0KHV7jLFmX+U5l1iWBXLK15UhrTHl5Uh23FFiQEs/G/0vog75S8Dgk1DRxvum
rMierDh0y5slhmsinNNPmnIc5aNrFB11xqGPOaJhXEv2ZC+Fb0F6AcHffVpqAOcV
W3Hyj08FfJ4dsC6UiF9NFqA0CVk11682MHuLWfroQ+IKLAVWo97DWIa53IfE2KCZ
KgZFOjqU7U+IwPuvSfe1ylm0mD6zoy+hj64Df4QLGAIw6sDR6Y+oSjT9pBX2sJES
ez//1sYtAKAGqG+LNpqaz3CMPIx44NCHj/RdekCx5+ogbEe6aiDIpxJiALTjlbmR
h75L1UlmH/58ltIv7wbPiDleJcTt1tDbehnpRpB2N/y6hW4VUnjtUGwWFR+keQMy
+49JbMq9eKY4aJHJFdoOh3JSKVA6cMVPBfa8yhM3A8EfTP/natya3gb2vMd01mcH
3E1QGjvan+tV4ZuZkltmNI/0aulOowEC+iRUumoIskivRoNGSabiKIEfdl9WqgEG
XKDbyST95kJ4bXth7TVbRE15uyE/HtucwYbhhrdQXGph4h3UFcQHrj3czmSZtQIo
X88heETouCHs0l5WtL2BiIjmqli1abK5MOq6EbiQcGX+OytR/7bf7IuWkSK+RWn0
hMPOdPYr6nEi7AiiUMe082CarsTkgGtiSdyGJcKkjj5Vqbjw5TiXNsUnv1LjqE5D
NM6IW6mnKkOsEpYzP4UIanicBdJBztswRAJ1zlAVkMZ0vpC4Gl2t88S4MlEear8z
qhayji2BjKQOeENzzlYkZnyiR8HR2Wm5TQvTll1O2kfkspcEPUnJSOeQfZWW+xGm
hCmu8hweth0JCnVmEqPibWfBrr7VmP47/7mSXWEGszqPQXNGGeaPLKjooE5rDacA
suXO7OYjgQtuM4Kg9tnCHX2q8e5Skj4BHRmLUkiUyiUZF/roMoQIf1VZ2wyCDVUQ
nkggj0ViLIPetIn0g9suEvj0uLoz+zW5NIy++9pI4SdPSCAmHAjFFdclCUJp76TL
z74lqkrc0bzm8AzqR1aIxoyAONPlkIZpK8SgaKYjX607hFzzJ9R86l6N7ro5u6br
8NSSTiAeoaKfsPtZImcoMIpPpQOnfxEjiF+KHeu9NgBVUbyYCGdUXEihrxOC2b+G
XqfeyskhEA9jVKJypIbOW7YvL54vm4qwBXxFzca35HVIxgjPaSR9WuU6AF58XC8c
RylyhU2/jj+QbZVVlb8DMkZ0gTt4Oi0tA9EbkEOrhI6YvV3UDdtwY7u5yWHu9335
yKTjaXfeE41NGeoDIzBnCStUfqmwcAmfpaJov4MlJaExJOxAm2TrrtZfNjVf/xM2
bzJbJiq7WWLp37N1Bl6miS6J4XNiUgvLxhodzTQ4ut7crkE6jWXNh7Q5ClWaLBs9
UYhUbYiKs/kXhviOsYL1fU2FZPkUcT0hiu/YjO1rcRBUPCUKPTB4lVSGb0AR4d6w
+2wI6AXMe7sAQppyt/SgyZdh9IVFyO2SDNaXzVrIULpWNO5NlKHkpqgDzNS+J5e+
R1zlrE/iMyDjlfiVijxfGpLqhcmKnOkjwq+ssVZQCeDGZMD16CtTNeFSvcpYksyo
lCBCB+TpNkn6akVYTPbv+9kFZh0umHadqFgIUnGI/QQBJqKCaAaqPCtMhfVD76Ma
H9f0GZ9NHb1+VOIpjN6iWtyyXvGfSUMdl1rH1GnLnYlMde6QvnJgvOgxfwpTf7ui
9EU2wZ3lStLYU5Xl1bOKLUviI0b4wm5FbLKBAXgkA5l1D4K0Ye9RkHYEG0WPN8ED
ymCoN9u0ljWzPLQrrO20YVv3/q2tbbhEktljJGj7jJYISHTsPwnfAbV2j4R51+23
si8Iy8a61b5VKH3E/hFEm5px9zGods7L1ZJCpjZqojTj3kmKhQvvhg36uRzeW/hs
x/JO7HjkzE8nT+Xh+vfVVUCJh2jNAGDUbdzJdnZzHnjs8IKOSo31zlTvHXYxR/VY
oMrM5Z5em6n9tIzxoC6F0jwb7D7s85A9uJ2LhM6NCsbCJ38hUoVP2Hf9dicvVsJ+
nWDvfzIpSWvgAewXSetXMv/HfhqInS3elctP4mSCTI+Fd++phoi7dlZG2ITis1ho
kgnWbSc6cdljebSV3bTlVVgZzy2wfXqxYmyAiwA0kGy7oZoQzKbtLkQkmhNezbJr
RLxYUAWAXOLrF912jhaidb8hbBTijmFKfaF8JliMqL5SNAoPfjNRpFuXGsaLkuq3
t0BUkiFqPtW32+uMp0+mPMgUP+rdTqwXylkcI/snTFD8CPOfsrqfHAfXo7uoZlfU
9vKrnnWo0455eyB4erPuO/SDHw/+dqTThxjNx+FhU784qTMtVMRYTFreJ9N1E4t7
zwy+aCIeOhdYD9Qaomru6KJizRVkC/AeD3UZbSJWfmxI0tvrdoh+wTMpOx6hxL7Z
l4wnr54lVxwQRGoZkHca+Cgg6qBZf5Z1OH5nuIHrWzNJM0BBB+PkF30jqyhG/opj
ocIyOGh36e56agaralgH196EjA7NI8C0llOu9SBwgQJCHkHIhpASvkf0/B5i3akL
oJU+RgjUehS+Cbvwj7sepBRqPCNN0TXpTX27Bpfx/XXXJcauc0FmJF+UJKLjeVCC
BN5JeZvdxRdXaIFBjkP/ASAHUI/CDTMVFwRisX/8TcyBybB24497xXEEdGlSe9PT
ivmBzNvPxfIqVg9Ihf9gQFi9JRlDI/bX9qEHYxbWQuSbwB9KHYWLtzrpFBB7gNUB
SjUVu1kSOS9WMMJuOn1jUABZGqXzs9hxGxO4gvMdxbTb/YE+RgtiMpiHS/8n5rAE
wW8YOPQP2vu0BrN+5WfcdhbzXuKDrWk5B//XcGeEmWe6VL8iWvCeZmlNN+91MJ6F
EX3InRqoz4Vfvkcy7c15HPHooWTUIbnn/S5nOXAOc1EO82xAFboQWKyeIRLPLK5K
lk9R9lRQ+v9KtYw+EybQNnGJkCy53siTwf2JP6jOb54uYu7QbUXrUyHL/+IaijbK
KAOGhx9N2CBLndBh21WpO/sPWFmC+uJR5JWV3m2ETz6g+gd7gn+PNdgYaZzwT+qr
9utFC0WmLYBBrcz7vLnC1/3k1JOnTa5ifDmycrM2kAibdOoaqad1t8tSnrIAJS1p
K9/BrXB0/+pWzz0t4QOo0c5UXueQJi2Nv0sT1bbJ/toLaxa2Q1/j6DwbGLBp+rby
Jr3GipAK7fwSb5K05OqlGumzq8Vwu/OUeY3gEi6KfUsn7ozVlmyp+X/iYZhFMWaT
lIHyBvOJ0B3QCmZMB2fyQVMXn644mzykNH7IAKLTH8VSOEsp0UcQ+mAjyC9Frmfg
obve7acOgJdTuTftYQGSremsmEe5Jl5vjt2Rl71LZAvGQArDHHJsYUlbq7VplvDJ
k8oGPaesTtU0sr91xHiZ4M3rA1xVxGrDbauG7BFoO2sWZ78FYSiJU7ngSnLn/sdj
QFtL99IMWk7prBE+ONK5/PBtTC1E7dJ4EtCVEt+KF5utL6Xq1CUxgJaFzXs9Sn3A
xTI6Ij5+JSDRo5QeZJRIpU6BlAHKpA2nFIR3mK6kdb1ebbJJYuqSrdnYjP2VljP5
OkH/Nd8JP032GqKiC76ogxKsRbu/htdlmVLQPrO0LxNKi5hwnJWTxcL4VzYQbN8t
u3rRGSa2qOkN36vCAWHq4V+EumVeOya+0U+68D3QE0eB6Elcq/cgtWDYqZDZinqy
9fCXAtRtYB0eZuWZqwfPOghPyoCM3PDJktiA01ns3s+5G52Y1tpav1gyAZ657TLZ
P6h0md7188kd30qY1JUPvzv3L6Z1fHBvRhjRoczafh+ofGjFQLiGO6ua0OzOgYhi
ulUzNrVmpUCsn4DmbSUD3rWTswI2LR4wC7mXXGxl+cpJy9peLwXxTgTO0GxgxoCv
vRUF68WULgRUL9ZtLpgZuuBxo7b09TUtTjw8uZ9XhmYS1OFD6bcP8/oC0/OIdh80
byaqeFpsbXzQweoqsfU4rhWMWmL7NnVC28YCEZq10UqWBkYvqI5B/SflI9fwC4eK
/kr7b3lTww3Itu+MeMKFzIabsT0Cb4HHtuP2LYfyNzyF3qMpa1h+KLkGWh3GHId/
dOhIQVaa8Nvrv0+g2899OTWYtAGRH/ZngD8I3h39NNf0Oa2n2HTXfnSgoNbrougB
/zdOXKCg5pt95O3xj7ZR++KazrlLNr3oR3qfrkCXAVzYDodL9RwGMnG7NNSPG1hh
euH4OtHXJLAsOa8YJfUPNVZ757MiiBiQJNQAuVvm8lgFpNSz/3nYEM9FZy1otLw6
bZWZlVCcRJMJktr2ZHze0lbrtWteVEWu+4DJ/F4j8FRiKjNEp2Fl2xn0vpup/c4d
RicnhU2O79gomdtn9kPhg/SZWUcQMSoR4AR7WSm26NArG13L4X+IYELr85hkTOPD
XWocZJyfyP4cMocgmtr6QFKMWg9vwtKFJphNiBRu8hjzGazrX7FiZTPLEqObqUo1
te6HDGtQrE7COWbG0xdhIK1GOYFbX/V9R1/ZxEFGMj6sjSOdgA/TSwC66Elh6MPR
rMkKJ8j8aqkVVxasZeyspApJJ2QNjgSWt2/N//FSOvO5enGEtewsQBLV36DICMPJ
vO/kRehBe1RmxWGHAKgdRtl9UIKHq8YoJvDTbnolKmKhuHnQ+MTE+gWrEKCBIFiO
EIRRfv6pv4R96WQiRfpEb6ga667d39wkVxCPl90UwTKAIUr318P6wiZj11CHoBwr
BviL/ElcZ3UO8+lgnL5+1/FL+D6of1W17gwMHFyV5O/bbR0HxYaNXVfLumJzAWq5
Z2+Ni6vQ2kXOOQlUfbMnu7vXPSkjxsVCG04SY0OIa1kpFXPODmVyUjHWg2jrb0Hn
DS4d2bwNH1s1K3hLiqqmztQ8BsEkVnny86ldsQ7HNTCGNKND95h0mGxy00b5xRf4
ECoIEa6MP0X18KE9mODRqTP+8gjBCFXa03zan5IzZSP/zNeA3xd4hz+SMX+vFymx
Cz5mNTPEoiFag9jsHLA+gcX1buCqkke71J0kLeeMlGXxa3sy7UN4MzhJS0DPsSlG
2QvotrBVn02ePWLexh91CPTvIX9ZCabHajCxobzIESpwmYC9EiMSWi8VUexsJLi4
HNeZ4jyWTYXeVdiCH2muzxMVb/5/j6QKcBVSosXdybM36Lqr21gkwI0hrhwF+VrN
ffXR/xtADqhTk6YCNykiDG9YEusOdIxpDeC6sZYFORDxQZQKx/QaiCFhy8gk7miZ
d703EjMEMO+ONhjR4kNrweEoauisdmBgmf52MUBpujsLffiy7RnsOzguts6vZjyt
OF7XLI4BMgjrNGR96uKBEabx9WxL8vBmURrXjAdSZ0cRSca3crAnn9iwkRMnR72W
JFQOXP7UG7kxi2OhTBnyJCLZgQkmTdWmE+l0zUttDskL67FZRSjSe6ayuucN9zNx
4GtNd/WCQ0M8p745tCLKZSulmgc13N2T/PBhCljvSPVTQAUr4WqMx0FWDTLeDL6m
1DMWNpNO24oLNqyZGKmR/Erc5hB4XX/wDCqbcwqnV3D2ScSSxBtUWusG4z4lZn2P
ge4MgxhFuxalzirwDukEIEq7S0aqv0RvAqq3OjtuEseOtbDRelnirh8+a4nx5BVH
9r7b9pcL7zd/gN0EIIuahAGR525OjmleNQkmg7kj2AuQcWHDAqUmftujR7a1xRKX
TmRFaS719gShlUHPu73iv22RZB7Yuf5EKL9c/riqa+kyj4b6HD51MnfiEDVWCDCD
wxiCjZRo1HP/U8Vd8syL+VlBoiHX6PTurAwNnho0wXE9MMz1IHtLOOj5iWtZyE+8
WNMk7UJSZkStB2HSqssteQsfO8FTWYZyKpNGHVN/9izvmqbErX4kgbcslg+9j4Nw
YRVRZvPuNV3hZLys3ibv/I7yPUnMPCOUpAyhvNB9St4HqKo+hTX3NQuBB/qIaeaG
pqjO6MCTMZvIzq5nPV+/Y8zTuH4esa+QW4+jm9VAQBvGeGvLboKJJiRXpjq4Acw5
xqRp8J9FVMDjLTnz+vxwzueD9/Y8ZUcCdrbQfG4HG5YTd8N1BIyz3H0prYo29Mle
Ii+2zPvd9lmHhPwUKfr5hD8mHwmnaO464zoi9KOQeJWsdvxBei1IfN4h2IIyalcK
U6M7RF1EL4eMmycDtU85iVeh1Sgn3Ajt4qf7PmWLHNmuo2Z8oChyF06SZYgqt7RZ
SyVqgwNicf+IzkS2ifwpcHMlIfWEzFqFJPAO9+XnFIsALq0EdRwS4/B8qXEPaCb9
e7GzN7l3ZBkHzABNwXj1w2RLOT2kL8pWK35xXX9TU8kVnQBRGqjYdUZ92z77fVlT
0KYdDU4f1f2QSk9cG9Ja2By6wqgKGsL4YJMYMMfHL3oLAfILb0o2sbA6IOGRoYz5
zDRVdLHJPHJGBupFVAbIAmvCheCWeLPjyswXlAbofMLCqSB8Vbokq+dkKO697m7P
BRCR9ix9sN1l46i+MUC4JLwRgjMx+7TEQx9mZtUQ82s3nDDTgxSnipQeeD+jcfiE
+oerTkS2dA9g7d8pctDRXfKiy+dnxFC6arF7s021RadblRkkzz39yPlzzGhh+y+D
fDEOx4nDmTx/jYNlGM+nExgseElSixwvRPi561cdYHejIzJaJtt2ib6MzkdTYYle
ADeEvuvT+C68hRMziSCIakxEGiaCU7M6U88uC/clZ9n3qqI1xA+v1a711p37fOOm
/EZxksWrGIlLZZMwKgfnCxsAJLZdbbtI6vzaPCqmMyqI8DxacYRiwfnKq519o4VV
7OuYekvOyJ5y7G7suFFpNx87lRsrtFKeywsyDypdyEe8BcSdVa83L6KysUUiqrp+
K9lKSRf8y0KMN2C4KsSBVwt0+xnKBLENlROTYMvBuVtgMUmAC697h4A2tX2CRCcW
clGuLedmfmJ6ySFQ0l3xEyyHJAY8Yu+bo25ou1WKTzbpg/H7yFykIaBBqwIt0jDP
hXm9bZk1nPQA2Z9zUUT/hsI1WbOvVY9/E3y5UPNbvIukbve6WzlfOnCS43Dl5qb9
0kMq3Hps5BdXbbrfGDH5Af0yiOupQpXvmWNoQbPjv+Om/IF8IjjP+C1dlu9W86x7
v2GyFWTz1/JprDEwmVdn2R5r933IRR7IZSzH8fY0AUGtmwIv38RbB9YJhCAqgLk8
v6nPl9RqmvY5TRCl2nICYDfUHf0K2/E11Kui2UFBRROdoc3UoJzokqm9qJsXkm7t
EH+Bn14ZW4wjAtpIeZ53Fmvqh1PDJQa5JIplYKfL1ialo4ytynH13FE3HfG9jkri
LFdz/FfcDOCK2LoHag1uT6e93Cs7dRAl+kdnYMgDDSbk9n3KkImej7YsyWBRByj5
BzKuiMs4uOktW7ZLP8K99AuwL5qMHKpJQ+QrhGW3g5mylZdqnnloGL6wchkNShA8
vWYExrMBr65fv3jh0vlO7H9oEDUYmO7ArZgrInzUwnN38pjlVkfxPh6tKXv4RJ0e
vhZ9i7ZPTGHPqd0MsTbHpPrmTOULSHFhLcTM9+aNLILWSbLiqh/wQl6MW2WUSLBl
vGlBIiHtmoy4tipdGSq+2b3kb1iiW4/QO06E4T3sWwLrFCBo64+cQ5vklbRVJ8J4
MspYDbm+qfm+kgXsTCV5KEBUWJXHuz7AIYfCeLmO2NKE9dxZhjdcuArExresLXuI
jwPhEHwQhhW4mpS/V0/QKWQWfP5dJqbpK4Ls+d72bAD9hu59p8j3FAO6cF5YtJng
1oRuhAh22/XUBao+o4kFMtd4+bkBSIrCTLWtiBFmt9t6WkoaCN/tYpkvcQ/efLjs
4OkFrlC8ONwtY4Cm6mogKqMz5EYsbDZyPj/wN+zhLU6WV7XdFlSpf7UpDspQbTn1
od0UeVKxut7sVIpWouf+d3rlpjnJ9yqb6EEhARNepozAfkWSJpKtQny+pRqjc43A
8PMFNWn4P/ZhDqN9DmWbXIdRbPpcWHfiZ7Vn9lk1+sOvfbCm91nM5otAmFEoBunI
6YtLmSG/PJay0rBqeiL89m0vb6X6Q/uid0S6csmqII/j9LSU00Dp/FuaC22hmaTZ
6juRVpWPNpOb1LZkhDeTleFeyYjAuZnClrxIj+W322RLap4kgaI0A12EK9zGI1MB
IerzKhyFh42CY+5o7x0eXr/eOHMHYf2MbltT210EU8ftPjr63cfUR4WFDwYN1Dwa
XnU04FHNaU/E/OZlEPOpOkkf3eoxcsH1kLHV+2dpmFxgcFukFdsDeyok8W9b3ZzM
VkJEl+NLWVFHSGjVf5MQ/K3fnF6BVt/51nlEwEuU7KPpIz774+5lFK4Qb/IB8JAr
TZYk5bxssRdnmJP0DK3HKR9SfjNd451DG+pOl4ipEwk9482WY3O/BGwsM1P9DULU
ZUGJXKPgPd3eZ1z11jS+yCucP6LcagEvXeej6tBnBwC+u0OcvLrM7A3UCoVQEuHW
6Duv5/r6kGnc2LSlfuWZL2gjcK//1CyqGhFt1V88U1BK1JsxFuw/bmnEdFglFFvY
x3VMoyWYJe8WnADJTC3KvusCRQGjKxoNDK5o6OYfUSjYQw4fzk5XWNiMPXwkxRfx
EU8bggQL1/ulMdZObB1fL4Y6BrpKC5xOukSgTEDiOZe+ssQCyYqa6EWWIlMnO4c6
P/uVjauGxxDO7Cgh8FViAEHTJOWLxUKBYk29FxQoyNJ6RJVaohClIbwqiAQTRlAH
5jXpp2RkZuYJ8mhmOXPQ3S7iQ/dnFTaTLHt9dWtdrzVN0dK8yU58ICSWEGPoowrX
bjF3SUnRjEGrhuzjIg0WWXDVGxUCFi6n5Tg7DSvd4YZ/s7/5UCM9i+UbIW3+aVQN
JZ8i42w1q5NXvLl/9urVr7c4op1uAqZvHz1PB19cLG0G/y6Y3XkyDz0Enow26ebs
gtEPkwB2Lb32Sly6CV2ZsiEo3SgC8c1NbzfeZhds/XzTKaQaRf3/EU3nw3GerZ0P
x734FeVRUsfZ+MoIoDG1EOoF27hgdflAZCs+LTWz3ZpH1gsxgikwhb9tEsfJkqO3
ptgrRtXykeVrE+BqY6HceTQbBif/7JtnlQiSo5AvH8iNYUTK3ONBFwI78iwutJAU
IaOMXsDRDGhnzZZVlscDZ18DhINU8/qS54IfMv07EVdQGqOriewtONJntVqemGYT
yjoQ9mK3KSQ9FhB6HmljX46T4Z2aQa83hqTM7dUryacXSm+jxwHg/ciGjTEUtdtu
qxXpW6Um19dpmyIWPR6uzZ8udRIBQCKEBuDnWybMb3d6JR1Nzp8SJzHNuDK2FyqO
y+BXzMPJ0urVDPpAARja18xr5R8SHJZyNDC8tVU0+scbaIPgWQ74O0AqHFV0HP6i
CCp6pnYB0MaxcHlRIp8a518BKv2qJvO4VvO0o8SyjtCCCGoLIfgQmleibKdoo8qV
3WjadY/1MefngFGhiGMLOEy/kMmN66ARFVk1zhu2CILV1MEliPGMwI1G4wlw+XVm
Mb/r3nhBQ3bBGxSXU4zUT8FelCqIfSvV2P9gliwLaFt1hL46c56QrTsip7NdV7CA
byoPZjn+bzRA7E9MuAZtLlu48inbhZG4TlO72E82LV//zV3OPDMROjnbYEnmKxu0
TlUaAgOeF2DfrCutcy3J4wa/Th8wGKj/DkrMxESJpPFYCWAs5t5/oAArSXuA5bQ7
FCrsmG3O+kmTqkPpKYM9bOOwCjHmEJaVg8s+wqNUDUvJsixUfdJF9JsYDJZ+mERD
rggOSl9ECqu04PRx6pGzwaCMpnIo5MuMkhM1UeqfXHr7PHwZnnU1wUvfcQhjWSWi
vd4dMT2C+COAR1hbth4ZiPVWxX8qwh8/dHmWMeL8hOFoZ0XWBDGeV+7hIaGkOw0z
d/dSH/sfInhdDfxb5WY+NSWAfJ/luzn5mAybqRYjiY6ijHVxlFfc0/632qUpaL30
yrACrQjdY5/njyIzT2i40gvmL3WuZnBxKEjRT7ZuZBDMI4yYBESNQWnCbFw/jbay
raeKUam0kAHdm76IAaMdUnV4dw0CygHvucS27buf6wxAJtIRo4ylByhzdut+YXH0
FIxNrPi+8J8Q1OJwD4k4/Kb9E70fnqHNK9PPZUN5XADO4bzemayHZF4g2IaWGmeP
pjMKi+gwhLCG8jlaE6mNa14LGJWZsJ3htZvBLrNUHLD+ufDJ6Eau3MPhO3zf4rr3
6pDwN5cosap3WQKr/doSwe4TQTQgeLUUM1svlDGYwz5lsHZH+vY0+q6a7oE/m5mj
vxxIdbA8hBiIMHTdnxHuJLfTcyEzAAsc21IHNngZAIfGcSWH1iEblNzQ/htus6gs
13PEfwoBWk329XydV8ARQLDtu+SXVM3FM6TXBMIL8od0UqJm2QbzLPIyzDJqZu4u
A2BhUO56XV8jYfPYxu1oaLkXs2LPgE9Fdl7xbiuirBIQcTduTD9h4D4dMTfVWH4a
FXxtT5PUSWVmPJTd6A7xr0QYPUj8hd5kAFNKp3/WAVpkSWRw4mmKeRWVGDf92QRc
mbLuemzYQ2Yz10VnGisBmWVj9bBvNI1qnaXNmom3HGKXylP/uUMxjLaFDO3mVhks
n0zoxcP8MNLeN2Evj8wUPWLcGWb1xRL+30JmQNUe8sytBXnBxofhXZVSEmerwrNy
K1UBt0spHFdiZ65pN7CYROA/BxXKD+iW30FAhZdC8eQ47CHy3KZKgSsHBI7BWKbQ
jSlee+2iD46pwKIcm0Os08w7w6NhOi9p0OVgZPTsoS2lm40qbwtbFr+4DKeeNVaR
k7r3cAiiNM9UvlTY6FK54uhGOSp7c+qy6k1MVu5EcbBEteXT40Ka1JZlLCpDPO+5
IyjzG8pZzuF8R6RTDK3HE5Ww7Pht4XmH+j+hMKKssGL+mS4Pa02vIIv05xJckklj
09gpFyvtPoz4uyyRv8Z7vPS7QzOYFozIMSfQASvx+RCqDGTnRrrms53EYQeqAJAl
agpuFpMkJzmErFpbMwn6Pj7Z3LKFOPNZX9EnUduGRmdFTXO1u24uCh+cLX/mAeAU
Wwp8owNW69OIesWu0B4Gg/riOJ3rbNs5/+mbR08YYtUPMTCmTPP4AXRQhtFhc9dx
iMf19Ep8a33S5+MqBB89BA5ECcQaj/LOgbOFOsUTnhqgellH5h1fpqcEyMoG8Pe1
udgI+tFJwr0npNwDgVxpIEpdix4mUF3rAtM3hJhjv3BYpK6IoaWQaHIafA03GGEQ
k4uVuK2OfbLoanWly34vkDy3Pyq1Ne0uLruYtrCojwAm7BKv4X9XEAzYoeU5UcxA
iLz0pwV2OC8nSsIlqg/fp/5mkrAeefZQoLxJxQuQthFnI0c0rOtaAsuL9APl+jb3
t+kYrwJQKOozTzeHl9rDbeFkLTAu5Gey2Ll8elJN5hUXjOuf8f3GKFhcyakrD7Cg
rMbuULdxD6qLHcS6Wj9K71eLnXqkGJa/QJvS69tiZovmirjG/ybCZEqJRIKy+Sw+
W4mwSPAcMh1BKEl/ViERyITelQzs7KDC7uTdgYvs/bVeniycr8bMrvTmrjCgdQh3
EPmaAYij2KLEYb20lteZKWij28U1Bi+grQf4EJoUjxG2KotMiH6ZHcCfW3SYjj6S
yjzIL5GTnWcbYtNYiJ350t1PxZuVoOe6RTpZi6gnPWA0OaMDBR3R+6k85szOVw12
Mw6qZ7JDWtwMwong/EGrsZV9bjPUpepN63NkMzLgxiXR/eMwQm6jP0M9leYEiuJE
+7FUJUZieBDDOOtiR9Un7Plrj5h89uEFowLIEYhDeBhUSbygyCN/rqcbAvpbv8Ec
S5571IcTe27ORJ39ek08M0fFdqid0aAM/CTO5GqYJVnITbvwqC9zmEvnpaMqblAh
5cHjuHsc6cVNkbJcMxK2tt3xJf94PY/Ed/0kUsvPZxpY6IzTmMssX7FMUUwNfFNi
2aGk0Djvam6mcp2PZ91O8QF19NakAima/ehryibJ1sCReVqSrCzo4ADVfPEh48cn
MRjRasjLQerKOx+RaWLpxLp9LVaJs0oIxtfuNHpIQOmLh6Qz701SwuJUb8xO7I+1
oY0j0oDE+VhoRo2DpkH/3Tn3hAw9An4lfGluK+BH7916WIQfA/hIHVK4QIQ+P3vT
YpvLVDhgKGcgHKxGgQUfDlPjyObuklwVHMSoHP9oaykwRfR9HbCi1+trTA+WevQZ
s/IVjVPzEMabBw4OUXO54r2f6VzC5CdUgEqn09rwYI2xS9XVEppMsYrDYTLp1jAE
IliFft0ksvJ9a8FfwTyJvPkiIhvznehkk0Q3CwDNx1fXHmsHqa3eZ3Ph64UliGEH
QHClCE6kYKTokO3aD2SGt6fbpFahMxx32dcs65LCXml8fJzrnkRaTmOguwO4hAU5
N39ovJi3vNd2+6+B3TZqFe1APERemaWm4Gz8VCZJn0DDC4MnpJh7inD7Fd7465Kw
9Jzp5NzQqnZqDaJgiTAwgfn7cpJekaev/O+rkoRWjelsk3CKTcEmkLiGNVWYVtHJ
HplU26EMR7/rWqXKiidDFIVHTScQORHnu3319mOpa8jRl8Obt+G9HFHVqD4N+vTW
i3/5gwfjOHz1zjyBVdv7NM8oFjVuNX2VLZosoBgfKSwjVHeOy0t+uOyHyD7zjHcd
ppomJtmmjSSyXi4kzfiFECzt9xdTXsey2pV7tbXBMErwhBKDhU0QO2HiD9je7+nq
vbDAnKrqhA0xBnSlJHuFOF21H3Sbp2cpWCKD3it9jom7eSN9svHB+V6gsYfOc4s6
RbOfd0svhNexYcrver2AA7ybMKWleKFJx8pemDH/vw9SmgYibi8VEEJ719yO7Sbk
4dwyT5rsQcuAUAnz+Z2kzkd96TP/WEMCL7ywTaRKxK3SUh6q/MMPaqIhr7E6zXpZ
ZiwoaEjw5AkkfZngGAvi9WdFZ+Dro26UA/xygMm2MKtp+DZwFvHYNNLu7aFCC3mI
f2bF+Km7H3SBJg/8V09i2VcafiESVgI4N3wdks7GBVIKVgLHTe6pKDMvfmZHcTjD
lCqTyE+iy9qpan0wWmyCvLFuo13X3sc8vAKysEmlcw3+j9DEPsiN9xXmUb3+32zA
RKbG1JWAmV7q2vRTuClm6rD+1WzFgGp2iZ+8EZtNEEGtPsQwUPKA8DM2sX4IZJhl
ylpvy9UzlkV1J/6dIF9p9cgx5k3W3MOtSrZNjKwblmjS0DOjKZlboxu/dUUABycy
D/mUeyr4ZWQzGUQuECoaxvHr7XS5FC3ovbkyT+1T9JMatSn+EWBz6YZGOcn2JNil
lADbaBblkrA1ARnvOweMWzSOQqPcfky3RalNGFCd8490P7sIVkjKnniXmTUwr6cS
3Q6BqbK5PMl3xRyvNA3zzQtbWJKqthS8puxMSEhg5kx3nzm60H2BY/1VDO9HcuM/
4ac0GQcrcCtCXF7INtfeI5RYaXl2j0tJJZMJ7ln0f+1pRnViC4usOVgCpJFvj1Po
dUF901CrfvRg5HvBkbqCiGREYAUymNxXq6log6hrFV2wA3P1GdWibNoBWmIEWDLb
2JwhP0mdZ8RQMLXbFlfYEGIaDz5BKr52YdpDtxFbkt6/T32jvsQYL6VybPBANXmU
HeVc/36JtZ+PjK/vZAgToHo8eYfwqgjrhSXj8pLsVoZ923L4CGmEoJliX4zQNSzl
JoDkQ9hCQ4rBtNCwV6xycLlPB1YSWSAIDaP5K5ikuejsE228Z+xpvOORIYZC/YOB
Xzt43eI04Dtleog7B2pTtYgUhhxTxiGbJJPB8dA+LCFZ08NbLhXw8uc5KShiqsSd
th4j6anZkEjDfzyHHYqGTzzR9QX6JefWd/K8H30pachRnu3zrKaGRU6EWeVnW1Zf
yk0kxJuRFJKKOdQEBa3VBntX4NV0aS6tL/zlJwS+e/dFChpl7coKpu3oNCfyr+cI
e4ExBkhlicpAsM4dDcLLSYxFWwtkV1h83fJAPr8Vyoo8C/C6xghjQGjk4vm1tgZa
GTElNUKU+yAmBpgvEELHADt5WcosDD5ceaEB/yBbBcnikP1AwiNuFvOkpDKsdDZT
UXG6BiBXUs3AIwiimEdz3Iiaqmj9aAigxcLh9o+oVw5eJHqnM1Pqh7MZItRY4CUD
mSmNuyteETW1IMKyISX9BDz37uQ+cODQVPpQv2LP6NCO4vouW8x7vBHw2P6DUBNr
wpM2UNNHIdyDBhYPHWcbiXBepVtcwRS0T04Ru6kMrnILqaAcEJanIriL1DQegKID
3b2jwWbARixTlZWT0wcbyVezPPNEC/UZs0maVgoljzwD24qWcdJzVHZ6rNREGn5H
bUcE9PqyCPSYV8ZUwhJW5scE10UvwiCsnW7kJYN/IKAbYalrZrIgr7d5MkVefq7b
9c1FjKqnSPm6oA+zuKwqAqiOrt04mLVQF6zHl7XL9EjfGi52Ot8B5Bp46EIj10sP
eu8g5g36EcJ42J8Gyi4g8kuV1gnS55JqFZBR7Kvwdg87EqyvHmXKOwZ/z/8paf+R
ylGUUILPy7/kmVWxQR4+tzRo0ZB9An4qx1gl//NmNEhzWYrmb6uF9hEYqISWi0pO
Yri+Bv7tF2L2IxtwGoybde8B+G0Gg4wzjQrHK/aY/SF87JZ6sa9q7Zbv/ucThWIB
TnXTIIotwRorfTDO8Ks9gL/J+ewkMe4RNbNFCX2y5VemadXnCNBZOh8/GPuzz9Od
1Qcm7NIyUA6zUPSQyTaHcXhOV3F2th2/0/R/j8zCX5q1FQqWgrtFH+GXm2M+jYvf
0oatdXba15TmpzH3Tz862m6IF/O1hfHskVFw7qcPd414Qf4FqNJyx2Ndsnnf+1fD
m875DiMe/DuBeU9qXiW4J9y2WslfkDKnJ0DYq7idGwVBrI5MsD1XtoVTPpKRmB1/
+NUj5etuUDDEiK5JamkrSoU/ENuYvapLf9RXBM5ZpNukh8xEEYa0aT0HI81Lqdxs
MVPidi5c5CgQKx1RIJaFy4qrOrgDHJqFZe/BR9CW74xE8KMmvnmiqbc6pIpeYflo
ZeuwSjBy8icFUD5WtBKVwza3/pPKQlrniKaokx1Sz3D+rjklekRy6efwKqlTwhut
6CIwLwt7HzrQIN1DVmMNkhJgHiORQAxXDOzS3PvjcoI3MJHPbI5h+CHUYT09BX5W
NRUKwgqjLQU1u3gDM3N5DMN1aGyqYoPAlTyNUA0o2RdyG1RwDo2ofOO6+EMlOXXd
ipu6X6hnDfOUG+7LqBvNQeTp1zECto6cuDW9su8DG4ye4oRVZ8tKrzHEIQXmqPgm
RqRoROpRwQvNWUBiRVMLST7cBQF4kEgUVJBTZUlOaLg85Ao7x11hXR58awqzPL05
uz/fxjlvAT181O/8d1yvhKamah8UkDKwIrcnvuDbUvLwhrMY6950L02LbdQ27bs9
t83UWhIx1WoVfbavGbUeXMNZH9sI4lsj9Z3qoTgrJ3yL/N6efPNeT8KkM1xmKYpc
IgEviocSc9KL53z+fdMiNwW/4DpGzxbLE9U8ZpxXDOCbEtzkJcxvXXj0vnslJIhg
AGEKGLtNmGQxxUW53rIv/8uQqkhiAqkdSCkhY63AwUa8MBOi6SQSSU+ZpmmstHU1
bQvUlYt4KqnKd8G++tpFZFrYa4bwim0NDXfcctKKcSjUheY/0rx2rkCwfhfLJNjJ
HQEs8288k17SFrydLrMfrE27/IgvKvmiuwiWZv/2QgKhUdzVhMSq53lBkVeNeC+w
Ozlu8g/outYm7uRgpgn4ZF4Y5GZEqPI2H0HUOFvWnSrY/tEIy4on8A8A0qFL44CI
JgZxZbpAxFl5OcRMcdG8jOJPAREqoj6raUNGii81fwIyyvhvuBAj+XdROefQBhkh
v3J57nzfHSJKKgsMckFv4YnPkhqEaJOYwCwISRNcYEuYfeOSUt0wJGbim8UXZ5nk
Q7xcrG8am1iPipDMfMtLB1fUp7QV9gapOfa7DDDeHGYu22qfwu7f7UOHCg7BB+HU
8W3D7E14aISue9Vz6ocPd43W37N3n5pode8cET/UEgn1kTjErcBiNFk+fmsfbpC/
laVOjrTa3DMZXiEoNVj3Ryy7+IZHxG0Gmt4YLTYk/S3otsiLmslcx9TKYeRWWtF8
bO6nPe7GIwdKmP/Qyr4b1IPkG2t4Zlc3UtvxEm10yR+ZorhMOzSDRbN86raz2DEL
2tgqqOfvILX0dBanBEgItzNrVUMuBE3+Dy9q67bbz1YvOau/XQMRAbVAG7AAxCJV
4YZKXrJ83b2KHDWBmPoIcYMujYE8/fdV+qJncUOP6S16TO5zO2VZJbuagOkKDo6/
zdWMV/XUsimxML2xAfrWFvLgDDrovAL7GbB9ZQxL04Oq7Y4RIPwuTmoAx+1gAkoL
nrahEMwG6a/hfKFU03XcqMighvR5YxgqolBbeMfGBRtOX+vbMqScDhXQYC7dZAqi
1otl2SLNSsmzGHfYOVHYdfx37JCS1W4TKtZn5UtnrEood1qaLnqQ4Ni0OLKBL+0q
VToo8q02zy62Vs7kUrHgQYLQgl0YnY3HJ1Uu9IOsK4yLWQZj/jbHiszXEbPAK3HB
hPd4CmDbtWxvPov8KeTS4lLpCX/1/sftAz6izvUFgqSAyKNKN24yhzLfM3VgmV+f
cWl17SNnov6+B3Xr08smACTakOSL+blAH1s08T1jK45CmQB5UMGZcCevRGPD/8jd
RX2uMiZacWYo/N1XtJXsBWrE/muqcGksmh9eiRINMGRdGJ8hxRAhKTJuZ6hzpnLi
2Bgg6oFmzSuDMg2edZKKszDyC3ru/fX7X4jSLNBWn3BueXNZFBW98ZH3KqY/rO4K
RDDLtpGbP0YKORfrJ2MGl+o5NjkZyofnX2n5YmPTkTOnjNyfBvhkYRenujm0WPfL
71BqnYDu84h7K9FyJFUiF2sJ+ydT1srV9Amf23Ibf6OFfE1hPH8/PhiG9dqzDzoO
uzWxGRjKC2XU4LL4swxZ8wzRfHJoKlv/ExhLLVa8SyGt5qAJejX9rD5ItS+wq6IZ
m4Dt7meZxGI7edLeiCfNu8WATvgv5lZhr3h1GhQ1yWpUDoH5vhzFRyJ4afuuLySE
gnpJwd3RRYkOgAwCQCQUnxaq7hA/Vd0ptC0QvDGKQNvkab4dej5veJ6jVzrSL2Cc
W+0ooEu6gCLMALWYkcXd8+ti2X1YGTeX3XBdzJ2PzMyZVpmFKmabWbj4pa8RmNrQ
isVHk2eIZvIMII9QWmqii9euP9guWqNAizVuhEIZTnoaS9n7FW322l4nU56UdxAP
MT1AkpOTgdcw4yaa1HG+SDVEn7snGwgOc1YrHHnaax3eBSXr1jq7m7rYtpmFYpu1
T2YGH4pOIzktRdGWPkI2seUbC7aL/H1db24YrySHv4eAgBJdQZTtD1QDF/tTubai
H2pXPrDdFb4IvXMoJGJKfIiE3eX087qDgAUZoy1OxnBkujIpycbGBdR+b2KdKXDj
hT7FOHHuHRttl/rr9aicyqHMOz+c7rZx4FFqRmE1yNWn4cqF5A8RoeqwPVYasGX6
fgEzksQRpoFhbE2XiLU0YmJToxiCQYdTo4qntmx5D4dIr+7xnVGvGHlkxx09rD4U
InBqJyo4Ju6QoU7SMpLyR6j8SIVR/9fEumtS+fbfFt9xbkbSPOvfpDo2n1FouSvN
O64kK8KgIbfGh/P5R+K3q7VFUIacvDpWIbXBk1A3WXD7Dt5gGJR5CzrIdLvX7TDj
DqtFU0777eMPsEuT0RqmZI4qr/yBMbwAFk404SWDEWTCqZUOs4+6zMfLPcZGwWIK
CtDfb3eevrFQLrqHjNnXpb0C5/Lge2VDvmGK5RHD5rJMbm+sijMXPNyX8OX5AHQH
DeiqS8nsbqJ70AZk0bpqlRhGtb+keIaFUoVE2lTZmvzTRVbUwtDsYLHFgXbq9/Hu
iKoaz8OEqaCLFYJKrtqHhJLWDXkL54zfFoId2Asp0AcR/FAeRTRMZ/ZhMNBqm3Ko
bq1EXpzJbdvTaClkT0MSJcHuCrpEgjQpxQqN7VQSqLyfHp89czPAFhkiqh2Q/xQQ
E68ITJlgaNijoq+zRK6VnXmSPXCzw1U6jEoQS233/CbV92KOBWtuhoKfz3mh/PS2
RyWmEmqCOOCewhf7IJ/uYPgE7T/BmBbPF+h7QpoRBhvhAqcdPYVlu1nooiSOzBvn
+jiewooiLy/2d/jCgd7w7qgao5zfUurHLhxu/28Udcof8MmUGN3MOVU5DzXNBJfT
m1h66IfbPKVim69M66eucHVp0yzKXljjzM3m4jatFRlYdvZYWaiiUW+EMlNq6SJ8
LEGX9E+JZNESzMKrDoKq/bVXB8PjznjBLXAZZygbcy9EWmquvISaZwjFqRe58oWh
2co5BNwwJpsosjdu0nwIF/DDeKM8Wnbawf+VRZYHbjWGziHSxZQCg5bjcQLTCpJd
ghGoIoI8jlQoFCfOxAhiB/pFa00pTjjkYoLThEXTzj3DZsfmvdNfX9SYvNueVMhb
eiKq0NnbaO2WjKmLmvJrQvWNHUbOCDYC5nVbO/btwGB85iCuhESrRjGKBhu7gLil
jheWuCTUs6C9ijvOkc1dADQU1xXLwuLp/ALM6XsTZkq00n8UggP+H7saZXqP1mbP
2pfhB1QVthYiH5zLtjms6jAzLga02RuoyOaCdYL9dJBYcPpyYYZuqeZWsAgW2CRa
xCD0WswL+4z+1XGXmuCEbIE6x7eL/nG0OCvX+FIXOV36YS8JEhMdJPKWvWUpWtqp
C6rHnaDMBKYnm6xNt576WJcC3DhhxGO1Xh1X2HhfUZGP+qLfxPDQv3xVEO68ucBU
g0UziQOuWt1B8BDNfPX8AUK8zNx3Uu6pqPvePBrXTOXakl3xPST56FvSIhgdd20l
+1LigXah+tD/is00QTbK6botpMfj1cIwYMSc8YOF3MjlZIIy03YQXIi+NepcIrTH
OfbEb7RYl2ih1burXZ66UiAHnNj2KAr33dQfwkopmsMhqG7YKKzRCkWfEbCQa/Dz
q5MY6FhJohFvgiLTY2Qrh3Wu3/vENVBZZTImDz80W6aZ+JvmU89fW4byvtevnt4v
jUXpuKFdT0PP8h2q/cyWhwxul3LfO9G5JHqpD/tshoAmqEb4CaUlApPgnHlmkPub
FIN03v3V9cfhec8rWpuzvVNhyV3G1PaS127xQBDG0cLtZgvy8VCk32HoHcmTvkx/
9Y/gOE58dI5XC92pSEMZ9vEqFeoCwMgaBufkIHk/1b7AJZC3fChDfgmKKP3ZOkP8
vzOJdKtLM0Iw0ZcpUElr5aKUDlr3D95IeQVLnqYEus7sXKT2EeQCxX0UFqV1gkS7
Wq9ZHylpKwUn+2HpLWpfmsePecv/aW4T/Nsazh9x4wWLF9bvDMS/Yg+o98t8Td68
4LiqRIJUh5vKQ3burF5I9qxeHET81pBhMHkkwk68tXmzCrySvSU3hW2qbUO8eZx3
PMrkn3Aa+4EpSmo8ZN3UYam+0Swle4mZZ8y1QF7icPC6YOXg04TZu9DziSHxOXP/
/WNwirwERK40SGvhRdeOstiEh/WvDfMw7Qs9PP+9qqcYy9tzoxjB6E/eJ24eGNxA
+Z1erOSdWBfqR/f+AS8kr0Rnv5UUmcxzQC5TvgWwUBIWrgDo+iPSj8bAxltjGMN8
tnmLce7Jbc62Q1N7mz2wWUSwesDkCbSwfJ7vqlw/a2O8mOKW3E11t1BPN1S7Q0JL
TmfZyH7BLhE6136SJaOxkRgLy25ptEf9VDcb6KVpcegwmcpE1bIWdvucXiq5mTPl
SnmCBzwmbfIft79ov6NexyBZ0L+fITl6139tBAadxZ+NQHq1xdNre+As/9fBa7MJ
OA8/JU9b7bQMbB7S8sqqTemR+RRD9juBI8Yz1NGkZljSmOXTNc/NFnYpsO9rJvMw
SvyFlH0wA3PMrGN5vJNTJCyy0LXTeyU0TiO0bgxFFIXST55DaO6F8w8MBCSsawhW
TTGWcMbilo4RdfU7gXWdKk3/Gec7+Mvt2E9a4aFxOBalHnNvFuunFE0QEU2rC0WC
XKnxuHP1QtWeN50tjHEQzUZVeWz5nL2GAtc8GsXsq+47vpxMAj6rgDWkcv4eaz5p
uuBslmh/lY0tU2DddWTAss691QVPPkbPaCvWLSewSg6/9+y3oIoEEd1AIqMJCNd7
ZMN8/naR3Omm//ACbX/jcB8D1kbx2y9ck44LBblpC/eo7jp4rbC6yShHVn0KhcG/
g3+5qir6L1G3ZCrwoWGui3MKBRsS+Nrgwf7UDWP0293VYtNrd7MO8XD+oyd3bfTn
PJYJsdX0GcPOpNJO/oMAiCrnQIyBhGdC+3+p1Obn4PTMDXSqhhXAmKp+GcT5y5Dk
Hg+8AR50CzcGyNAo4z0X4t7VkPQ0Cw8Sh84JGbLcNw1PIWYzx71kB9Yl/bg1RfKv
ai8WNcwgDYjQ4iO6gTKAW0OYItHuGeA4XYagCsV60dzq0RSuJ1np37l1TGjO6hnq
0x1DYt4wQOUjf+i3NYnVQNTFwqPU7EEAUwjxt+mLTAi6cWlCdVj6IZNm6W+JkTgp
qNFXeEWHyyV1HRE9duNMHK7bykqN5If1Mk1a9NUTphHbJ4+hfQt7nwE9B+XTSPNW
us7O+XnksMYFfo8Xie47nJV4p4vIkid/hWDFQKXPNacR+U+LUHxFJDWhGFFxCrc7
aqPol3TY+Wt8n+kHhPgpdJQin4YYdbx+pFl4PK9gmylG5nvdOg3xD9uWdvMR6QDR
+qBs38h6VOSxN/vdWbaiEYP/dmh2mnaW3zDZQFq0hlc8XAGiykcPQ5kY/lz1VEjI
fLfoo+6q3luQjjY9u3VEODNZsZfrmIwQh/it4gxPjW57WbK6/7Y2y2FUnolDtDc2
mvB85s9OyqXXYlapQzw7nUTe4W7F79hB2cw9Wb/BxinawS2M5n9KiU/UnskB69aK
bYs+O15P00lLFUnSv+3J3qLH0WZdOWGVrML/9HzrZ6UaTxGR4fjFBUrQ6mplMMPR
CHpV3nEZZKsLdV9hnSFa24DFcHiFLO+S+QrWK2N+WMd6yn4dUZ+mPY6EOnLF7PH6
olHfMJG5urP1BB20cCQge3KIeItfV8c/EvTJ79Avg8RlsYe7IbPDZ5IyoFshQuPY
MgKuIUPEszFauMdYiLpLvvMA7b8tSrFGL6m/TbTEZZbtX96uC7IlM4rIKCXlXKsi
6mHXO6BbvWeaxKdAk5MXJn5fmX9JhqMQEFRXWLFy3AXe4o6Jvy756m/pNeqJv3F8
X4CyWpAzBGGKQFbQtKxZBC9ksGAMoIccG73jD/2yLlsmTmA7bv8dJ2rplfpL+uge
SNHMjrkIVFR/d6QBqYuFewBf/5M4aeKGbMRocha3qCCIXrULH0I7xRm+PRV72bO/
rPDT2L9ZeJ3euTea7R2ZtNe9XKBbPD4lhbDgvCbry/fDiRe+nuegCVJ0C6iQgUxQ
56iGZTc/Q40ZdEC9aeRlfzkXrrKxgK01fHNrl+nxnqzLCYQfa7N3C14kaWSH/oFS
AFerVJiKAt9Km2bZCrjnAZ+Dk8mSn2O2vzTxcZiQtr56M8RKw24or38YAeSs76uP
ZAesVTxYkKxACGx+ufGQyTgRoUK03D6n+3Gmbod1e1yfQtcFIxSM1RUHD+/+z/s6
o/JojqQp5c9uanmJViIHZM4uC34aiBccYsd8eYGHh2Fr9FMpYX5i9wcDmqRD5SP1
5UopcGPR6UAdsQgx24pppTZotjhz1HZjw/8enEGET672xenBqQh6FxC3I2lLzgL+
Tbcg5BN/jeXl2G+i7I6WUAGjhB1jJ5ipJaghQhaLA4afzy+2CeuHICVnORQ6lPQY
UhdOF5rjs0BLsm9UdTaX5kBkX7PZto94bCuVGxdyhmMMNWSByz8fxIRsfjcC0lXR
WYWWmgoRMzgG6nsdYH80Vcn+cMiqss4+F2PVIFZI7uQ8iJwZlYv95G77lWrwdvx/
ByuAkObF3vyeuxQmc2jT7KZuKPy1jZ6IioWAMzsKphe2OG/FyBBp2TsgVIbOrWE9
+2S3rmS5ZeRsIlcBrZGDW4Edww53gqn4WH4mnw7UmE2587/lkm1b4WX+AFBQXvRF
deu+GOlZ2bcnsMtFbgwsXWWTOIsNyA0Z9Kn5i75gmT1sp+R4HP20VllU7XAEwL2h
6zE+gDP1SmhPTGLA1ClzSILgCIk+6jCqabX9xgtTPib55jxN3HUctCO8Vadguv3S
Ay/NF7cIRwNRHI47NUuugb7zNYNaBGE0/xIulIWsR4ixO/yJgnOB41bPeNupKTxg
DWbasN60Se2Aln+kQrDMLY9WN8Z5AtijYXUDvFUoEhx4aXU5UyCUh5nYdJbXLY5V
Gk9iUv9hmblziiuF/QTUICXIHmYbIpwLtyRVaxEXMAeEsA1+kMgnUuCwBwUalkOp
TUvRxqnR3xsE+IPdxLR9imD0MFp1SbnSNth7ppvrwzAcGQGWGdnTvVCx36FZ3ZYx
ZSBXwBJTTdulLMsVUfEcosXFbX1fQi4zn07uFvdOehhuN7Mwcn7k1TsNS/5hfUqc
uQlg4WSh3asXBPVSW1GyEnO99nTiQrG3gixb253jB39njvXt4jGJQESUZI7GX1zr
aap+w3Q2PK5PJecCy5oaeZLS1rB+dBcHsrAFKmnaBm4zNXvHzTdvf0ZM1U7X7A73
iTXqDLkvdiy0QWFDRfV31USoeyIHUT4F7Jw591OcM6X5d7eBwxvaJ/LZi/wweJbv
wbAHv0WIwIoWh3J2DQ2+pbB85uT5pUVTJW2LGzOyJKCxw2gZ6BleBQKaikeIyV1e
PGwZC1zhgJomS1wAW5mSDMzF6udnYrQAmk35e9IK1xG8GmeVFmUDyQP8WF1JGLU/
IokM8iJoXkIOLTVa3yd1wRqXrOVfoIKSyQUryCeRQf4bsyZyP7teRmrYyPahFg1I
b82B2pLJZrXkRsX6TXVyJUJXaJAbGFlhblhCJrpVlhjnHpJVB7Cw/9JgeZI0DgAJ
g2XneKEEhw+qAYvRLV8Hfuz0eAPjq+M3PYHruzUmRaIegvm7NRYprK4WX0iEvO60
b3kGJ7u1XIzjop6NAthyI06GhIJFHJuNDJ21uzRTbW13jhLC2HX0Op/zWctQKAR4
C/FnQACsjAObOdm7ZJtrVSBScF3JEHoSg8TIzsBZrT5feqX4L5c6q6b9WTaANZpY
GvbxJkWVBESPyauzR/PvvYiFnj4gXdYuTzJuyhS3DYixXtStyRUXO3XtECCjBkUO
EVPnI8AyG7AkzWBnP8pD2B8w1KTDZ/Sd7tcDZwXkX5SObqO0eHOdQI8/y/cjzm38
XOOeXtom8UpJdJ/YGazrAJoyYW4f8X/P8iX69iKfYuWxhOuOnobwFnzL4Sh7NHRJ
mTuIe1zkSt2IiMUZAc6lPMRzGVGpcxUlBM+veebw+0VPkh3ENauZx9/gLjRAfQZT
cHITte1RY2EkERVnDmyKUVDC8I8ozfZgeKaebZheTyE9G7bp1+3tLbqZshPQsnA5
SLOb7IQxD0N8KxYkEpvFguQFFNd2FdfIgDuvdTxb0AAVUbU/wNYaqzUks5d4NhG5
TOwv1hq7N/ZmQe/lrt1vYRTE0ZUHi/ANBwo/QXzCyiHmz63xbq9C9UEJUWTdUEwO
wJm2I/zzkF047eQd3X21qXrulwBUyMOjzOtdARsxyG3KNOtPuL1cT5yDtVaQzcLb
dOTsR96rmc+gbOgVe2LsyNrIVdZ4BA0Hl+KdE5vSP2CfKUeWM5B9ZTngwh0MLCmB
z2qGskMSsmydLvRxJlsL3aNLUG4JLJ0iJ6CyBU1rbp+3JxFnmRIPeq00gh5SafOl
prHhJQbvQlBi1UL6T7Lzf/5/d1OsrrBtR1ezRUxNNV2fP79Zdg6AjjBRjLAYZkw4
cjQu+NtkS5ctBHyEfFxOWsBmNvFAGSYXTC+qc/hr+8XiRaQVtH8cRtyttRArhHJ9
5O1zfKzwpNk9yj79bDlTwLNqgyM+5cqf0DlAaMsDgfF79T4nQiQrPCAJMk3DHSLY
UbgGLfRfbRwVc1FBMldRcB/wYs0vnr/avMvp1gQj/3kuHHzzPciy6cNQMF4St4gr
ZYJ4ZgMBwb0tBQOiKMmgsLNcKQQ9nHzb3F65qiGzAjI4E3jMGASDdt86ax7lT7Lb
aaZ3lrY4ZcIO2qG7FsLS10ijl03oiDLEf/NzH/+dUBOZhcuHVybql55mnwvbPOnA
POcrlYIyXksCRtA8660Deomr345ochB1mIgvs/gq0YBg4r95T3koC/m7+EiB4gzN
fYSsowy29BFdDs87AvXbs0icRwaU9X6QfJKwnuoPsXyACYIR4hp9u3V+wtGZvK/E
C92LOZJxys93Ru15RefT6HuPLZYx4JJNNlBlzq6UuFiA32ME6b/bnJ0vZyeFAtM7
1K4NUyp1N8C1663qeGjktSmEf1joud/k1JvNdLNlaMcK/pX1ECshAZwI1zMamy8q
4IqIn6hZj+NtzWZuGM8ul6MjP6Hu9ECbVk7P6A3MIa8Qfbfshu34BOlk28bo5GkK
2jL1Cfsvc33CqtPZP6qtI0WiTfR+wuYoCUVPhS21oUw7IptPF/0F8ihwmP6C/wUX
9p2VHgeznyZd6JCRZ8LsBWr18FqAk5w1yma/Igc+VSK/DevJSgt/iYPDgB4BA/N/
MYKb2V97pEgSictyBnZ8bZEPdei7V1tWXN2eLLItfPbPggYULyuyLUbk/n4+qUEZ
nY6Dtj4PGPo6Y8UuNnCS88SF3kg/mT8NvQ0eFSD5fZbqApDVAUpPd8pN6sEKn9bn
dswuuqJR0xnAc119aPzobmsrDGu2KV2y+xou4frWhthXTNaKK4Dab+2sHiesCcGf
8oA8PgPFZCHmsd3/IV68uzW+humrSaWNnBWSzlyQkyO4RKrP4mnht4j+UjV4tEPr
uqwGiEMPsHIAgCe5G1N7E2kZiTowVW/xgvlwuoEZp8winRBZxLSj96yKtLUt5qlt
5l50MOQpF5fs/sbrxWZ5+E4QvJuYrGVbjSty2h8Oc34QxQXHIzY+wHnTkibTKgc8
De1wNm5zZRsT7N5muazE+UJDhm0L0yy0CF7Am4KBPMAeIM8kf4fO+XBRfC6Wb3iR
6pkxVOD+MA2PWGTsv8KyAuvcWLFsqRmprT2beKoCc5xoy9mpGpDMt/zW+3DTLTCt
7rdu/dK2COf8KgSzT9N+2G+VfEdtUcHhHWkLjr7ok2jyb7zj3NT6OiqzjnpqIJCS
V5DEueMbQthVjNaJB3ZnE7Ila8b6JfJz2bU2GW3rg09P9DQKcv7xV1O4QvnPl8Jt
HwYD5cn3jU/aAZvjUcJYN9Jc6EyIniPpPODCRCumpzuswX1GNd9QQLWBtIbJHCIh
CkOybsMPxw847jFDz8xUXKGXgCZ8GujPXur6eYruvlFgmgWQGYUN6BmvEP+9Jcep
ZIDmKKaIK9BzM5Wj2mbX4HlcwoJ4y/zxZfZLzggux40CNz948HvKT5ziZ0badE2n
Zr1FARpBq/a2skefpF90mVbEV/SSUUb6XliZUFDHef7YEhTJ0M58LovWfzYd0jpS
eVv39sa4+WApCDv+tZU1vd3fvD3rVsXA5yj/PoaH71PozTKoYZN7lQxPEpWAwBWf
Gh+Uo++ymLZioNhJSqxKAo9sF9yqW8UDAvQhTd/wcMl8TVYdvWuwWIdYiW4xDz+o
iPfVDZ6igyOKtxoCn6Ztp72IXiR7BuydFMcw1/0UVSNYfB23pY7KUaMW5p+8a9n+
7paLuGqr5tR3P175I8jz8fBEWv6OqwAhaWX5pWoGZFUEgSSF5R6WaIt6qviuqlfK
UmNfi8AlRv40J0AvPmNKhWDoFH0GSmL7h2mNYR68FbcRYmKYxpKJeBt8FHpsl7HW
VTnlO9AMkwTOuhM54H/diXdHbW29+AaN6UEUUFlQIcBMAgjFzZfvdkS6RpRFR36B
gN3EdQNeZMf/MPy3BQkSDWicyh3WCStGOkkmQovnxS11fRYG5r61IMf3a5hYU5yy
xFLtL55srIGWQWgm99IUm1n1y+cCoeL/TuO21GRfcxl0n8sXkb1H8shwYdP56fGl
v7a63GGcg5PvT6g8w7AJ0o6gT0scItbvG1k5nR/OLppn+P8HNakIBvU2v0mczkft
cT6C/TbCSdQn8k7n+u3JdEEtH85pN5hrGyY6L6fA2mofmflOPSL/QIcIP5t4+v3r
U5MHPoQU8ZG4MVZMOTlh3kFq6xXfa9OiVibr02q1t0psS7Sv9tzaNbicNGWCKqIW
Oic49H1sqhQ16WBoZcOlqT9b20Dc+mCJm0mL8Gzo0APFg0BOvo5xGE3Nsla5pNfp
+u/DUo2YimSHv94/1xcg08kR83OUFdbwszjF8hlGtzF8+djrBA0NXFqsIUIN/vgB
KGvrN7DNRdcmxKDG064iA/lNeXWhfoFrfmhiia5dptV2HPpKzHm4a0aanONJVJV2
K56wLLrtvxWrpY8znXWKdZlsqurbibI04nN67onyTA6fnDk3ksz09CRkvovlXAyv
D4plsbjbQ5lb+VaHe7xSwAF6j2L3OoF5ampTsGStMlNykv+GC+tyXrXBVY91K8WO
N1e+hCVK6DSvZ4k4Rg90t/UYp4uj/OJjP7IsyhraBn8SEZBCQk5eg7yfq+UKGUm/
FohaFYS5XWl42ptqy8kfUDLjOCsEs55E+2mkvyzx1a5opiZYgQ/5QmKKF6u9cvTj
QOnxfWMJ/CJmCyzT7ZaqIBOrvs5P7qIJggEOg0ZU9JGs0P7W/1hc6FcAfUkflCw7
efsPRSaggNsfjFvpBHIg1u3jTIzrcagJITN62oLTX/98BODKSqL01BbVDmXhyVVh
4jBjOQTazoKbWDj5X6exG1UAYlsSq3TZzMlUgv6OHRuKY2L9CZd559vuaHH0dRDL
4l5mx9i39I5W+ZlkJPOEdGyw3v6yN5XrJy0C0Xnym5a/tkCKwbZLkIBhfOJ+Yo7J
PvxRjliFdQOMFiDtXS8EnB8PpDxUDBtGm3tJ5EmTPIDxAh2jV2H+pL6iP56pdxv8
1hdKsDlhKug+t1j2AjJVCNBhFbcBCNy2ks5lz5rsAF5cT7lLIPTea0rhT7V3ZkaG
CGl7Jghiwzx/OAkR3ssadBTHrgGV9gHi/enOtrsvKio1LGmph3lrgh40n1fOgA8J
XsTesenHULymeMxQwNmJID2ZdNBA31M7DeQD5V8jOinfWv9TJDi0RYVrKLaXhaqt
6DiYVkHbZkmyfH3zcaKyi+/3/w8YH5Z17ml16ZdWGrukJ4E+H/nPWdlKtv6IW6XM
jW8rQGAvVo4kl45ckqTLYS+EUUC/rcvaSsAs6P6hUp6jCp/7GM7FxOR4M1K9QVja
g3c4jUIn3PSlzCLK8LFOgmntYwLa6qXsif9DtRJtOHG+Op+Zs9Q9I4v8vX51+aEU
NQdCQ/QjRKmtKRTNGq0X315oLcvijqU8Wx9Z8QG4KmqIZKBhvCx3OQJiLc0tz6tg
zKJlbpaQ2dI8omdVCDyRnQLp1IYuffCYXsTXC6oqQk31UpP3Vpi/4wM2Czy1G0Gx
UVDYmRS6Sc6TA91hC14A1NQ89byFStfAMRzeZ3vmpqddrGMCjxXbe9gXWfWGxtWX
Y7PMnf38seiiwYLjtZOfoRUrj6SAbVqhSCpE62C5szASEAawPxQfmU7NxGS3qFHV
1LOSie2sVaXP11yl4Uz+IjUne24ZfH3YpOlac+Z8NBmsPup84WVX/eYixpgB0rag
T34nWoCGvfh4mTZsDgVkqZ6YY9TmSXQRQBJzYWa3+5x0o2C5ETTA5Oj3mciqXoCS
9KC5+xYeVEt2SrlzinaSaLRBSvNLJCGewlGyxUXndJkwj/5lV4i/eY5m8sf8FtCP
icB9U7KHZApUMADtOMJAKsD52tAuHhZvP8d2n1H548CCkHy/gjMqAuMss++4aLY9
1Tnm+WypiBNF6Luf7hYv7iL/HGU+NiH7mJU1KB5rBWX4uaf0kFDFhaN/FMxcsc0c
1Ziq/8Cg+Y3lGo04mtTA7f1mS7mTFjuN1P63ug7S5LP9N97VzIDhZp1fMidx0qWp
gcefc8d6LwWNc4kJJ/p6dgnP1fpDhGQTWYuh1fBdZALvd/wR137Tl5Csylf/Bfv4
F3jSBEBi9CWAS4v8co+O9x+j9zEb6gNtbe0d62pJTNiJIu0ddjcozOfRebeuPGsz
VS0smO9R8dLCmSeDMGQhMyH7lBU77BLiCzOHy+eUvikv3N4Y60WvJ6G1jtIQViKV
e7ENMYiXucaz3npwhDIkE4NZ1FzLdPn+ELGBT55gBg1x3KMaa52NJ2sF8xY/dENe
J6p6ucwYXDBt3sOYcnvasRroWbb2cTnuVsCPfZiTeY2T32Jg1MO0xC5wIwUrgJxw
vhnzVr9qbpce0nfTubsioKxtak/UQVpK4hnTothjnVHZ9lndauqe9J15QfdCQKbO
5PXFlD147MMCPVOg4NdzpelVT+0lcZu9y8i5hXzY38dTHVasgVaG5lHAvRpnaAHE
5KubOvl+e3DT6aSQjNIqvzyNjFaXZRLZI5i10W9+JkCzGNHPZPdn+XRDSAHwB+T5
EQZtd6srCoA8xxbwo8ZeLUnBXCSlv0RzI/RRw3uXd5493TI0xepSEYmyrbXfhNSB
aWkRgFkMhMjZGPCcAuFezSopUsAP59GNPkm5to8RPGyWjRWAA4tSC3i6noreg2bH
uFTLtBkYmH+Y0qyV3E5S02kSnYcenURrlW59+ZW5oF6AH06EGgh+XZvoETn+6G9K
UG7MEdYMNVhyBgnYcgsMxTSCf6+MXg7ZZgykkeGGO5v7Bj+y/ErMdk9mm++B0bCX
SWhZa5MIM303umIq78bihX1p5TjJLtCEQuKCnnyc/b7H3IeVj2kwRfQram5X74qa
JVK6bW9h/J06qfN5qKNZyfFgetlg7PsD9ia62tNqXgvLdi6hY4vQwXGb7Ag4tBGq
RY8r01UW/dI8UqzH+OoYsk56VCnPuf4kqRfyhCCwH18kodp6RS8edBWxNgwXJHgE
uIfi1SFmhZG5f5LsjIQpUkpEpe951qrhr9BEqugJfzTo+7/V/bzs3oysR5rVNH8G
hhlNB8Se3F+FAi9BWoFJmfFddllSr8BIIRF4bJOx9nK4hL6bWraIklT/kXFK+9DX
YGvG/KFgpfubyk5VR03RTE4WlJ+wljJZD2PymbOyeZk07VG49Hi1lKVq3AkEMCFK
vL6lKdgNTwq2D6HbEkHSSRj56lz3ngVpyxcDD8iuloW3BiAeH6Mh261R5izS0VyX
fi1NgZZBa/9+QvlRcOLm6e6QZznmBY1UUkH/sKyEMlpd9IaXdPiVp2HD71fe18eP
3Nfo+5sDPBR7Q4GuucZ05icvNWtt7xZZV2nL5MSRNaAqTNa+xUu4b74dbI0IFRWv
mnUDQF01OgvP6y4ib3feRGupL1MsKIt90noHxtpdfNPPRx80U4Rt9u+NPK6g78iZ
o/12MaeeshObopGxuz86iSqo5idwsZUoDIx2JXZoDMImpF9om3CSQOEowsxr1yTD
idlbs35NtTp5EnOdsvpZikirVKhdNAPaziJlBM0dCqbW77HRnXC4I5GKrE6a8udE
NI/Bdfp2hx5eZbAU6jomC8BiQ+8tc7jnAybKPqn38nSZsnkAL78/iqd4v0lGuwjE
LujPwVcfP39BP9CJn4LX7KSaSR7eodlbU6ckeuFDrS7kvWwr18Pxx54Rxgx5h4i9
nPdeDPqvU303kpEu1PjqapTHKbCJ9vUo0NevEGALaIKnUyx579rHyhkZdnMF9poa
JL0nKbb+GI/Ld1YGC5IHxU8TQ+N/tF+AiTA5zr78PCLHa+HE9w+ZM7dlsPIAK7ye
4BgTYjLlQCrSnhh2BJ43utgTd7cR9xjuSevePvMqI8j2ZfxQ0oTvI4SY7oonD/4L
HqbsCPpdRnxdH6z+UpbRdAYIvWv/MRk4SrR45DyqLO4Yd+xroYjyV+u1r4+3kZ0q
kzpGqUvPogstT5SjC4Ipo90Knc7609PHyp6UT01qnKyfnsSVuLHLGqJzGmT6ubLa
gm/vBbw4WWn8TzZuN4juaD1TE6Spk0qJxjWxkMNw0Ajrhb/ToLpIZrNabNrBHgrm
Q67aaVTwQCmrKIDkjdQZK9CFGfJ/A0RZ8mL5HporhvCSy0u3Ad2+JwPVEJH7eoTW
usabxZ4jB5wrydYnqWYdw3H7dq3Ws3OL7Jehq/O+J3PhX0wrvWwLP3iDjo6ijPnS
oV2rmPhrKq7xGCKXB77g4Wp5OEXAgMZJ3EdaupGEb787C/cLxaaJ6J27Aiv43X78
MJEjrIXClJXSLpZj/YXQw9kP7yyJ9x6k9ggPnvsw80y30+IvBiloIQJu5ExzciHo
PYlm6Y70irKmKEEXybJW2owx2jVmxYYbUI9tDeZAJ+lR60xllBLokSdAxAGx6LiQ
LgTceWYg95oO4t8or7EQBShWqJS2+FGM30ztJeajqG4tft1wtDNbdOkBaOU68+6L
wSUqckzVNEqMfRRMtCO2PfLCmGo7OsG8tYIzJN0J10/UDY+R4k1L0KMllIYmwORy
3WzYDEEyMnNVGR5FdHUg4fRKlU/ov+ozDl6i31Y5Wfrmbn+th5IFMGjyuoN6cnLg
TzF/w1vln9Z++Cl3CG7uE8ZEtBycbeV18aXZ/quK+/GhqoimS5lole9poYD44Q5c
GItsj39RPhn9O5Kpd1t+czLB4i0asFyXYMB/HmrS9B6JurMf6QG7nz+RJKQ7cRcP
tbZRLtDgZ2n3DDwOd1YoRKrwWoHEG9aot0at5vbN7JnC/OTzkyM2XsAG1FhVBruJ
+EziuHXOP17R9EeecNoKy4VeR8+gdWL8UwaFmy9JrxAbBr9UIMwr7kebEoSJTJAu
iXsmBdWm0+fKDCYH3d08AuSQx6QByCctW6LsG+B1wsF66gQAeKE9tdOQQjdy4Fwb
COBl+dky5dF61wDh+FSxQRsl27rrHeo3lUwkxI5QJv4z8jRAwwzp4eCgrFAQ+qOw
jw0mHI/pTwida3ZAbj9lj+YWL5/oSfxV43f656f4Mu/Vv26bpgBMjmpNiZo6/jfS
IsjzPwebShJuX5vfwC0T5ROlozR4J1su19y66/sS/9QswhdHWKNdFhbHjN2WBwNv
BgUmo6hN0JZLA1V7KsXe+rlRqsBLKmCQ1qCLoQwfFLL8LS61qmBIsWUCTYvU5Gfm
ICEKwhQia2ofC8PhWGY7gPv5B0F0udX2AKJQ2pzzxYjWFX28TmlfO0C17sQPqWmX
o20ujYrD4o8WzyhVOHTNKDtbBVMnk/L8MmxGD1222BKtbNUSbZ9HU9LGEV5AIVQY
oT8SPY5xg1HbC+v3og71nKZ/t81YsGjXEAUBIxquPxgI+YQ7njnKW2EGpWaB3ooM
lRelJpIvRSjqY/0SCHCMPa5ngXzh7Xjy6QE39vitUcWKCZ52yIRfBCQNFA2rzKVh
YKbNSFqikklW/NunawKIER2DKUA/qHcefYQcNzEVNkDhvyqnHedFa7GRvJ6B+wlF
uOOBh1vrW8Bgvyh29PMouzb1mNOLihAQTwjNBtD5HBQ2ivGXQhue8DYnkk+bXXPl
aQ0nyg5fs1NOVm2U4nIXPmgT2FHZU+oZaz+yX3HdKZn9yJnvEK/H221qYjSCQJyw
s7+NW2PxeAD8UL3INDpI53+E3u54N7bx8LojfA+7gLZLdV7YdQt4Gxrx5dlLejkc
Q0TTlmvQ2xmSJCiJ0FZr4PG3ADcSnM1hxO5nDWtCD97JMyoJqCXvhmF3wG9rPZku
PNumjO3wBa7wDsvGs78AN9uivCe1yVsiV1N+UnJyIWmwLrvH1pkhhozDRt1A60oh
eKl/8P0zm4t5TLpb12Y2BMcU6rv4jDodS6zTD9/DEikmQqm1EwlERTVEPmPEUmeL
A4kyID0jfLoTa3cvh9cS3g4MZkUIOj4lS9U7faxbVmc/RaTu0o0DT+yiy+JPsBEk
0EgwRfSVdK7ds0ozjZdyZ8WofeAS+QYfDR6qfcjuMnRBGO4Q8ymYpeApgkUWHRwZ
VyVcVOM037mkQRrrBcdY33S2y1Etvw0VcP0mL05t1xhUVAwXnVxF29N5uw1/pIri
l0L1PLtAi+H0nRJZsHZomoJj1Ix8D/6u0Gf6LbB6HuCJTjLSRd182yJ14DBziJJF
0WrqlWIdnPHRRlmNQdjJVRUL/+ORAtPzW89mmeX90h+te10LxNSzgizHtz1rBhnK
Njs0NGCfKoEOGWW89cJQJuG2MELEcqkhoM8tKAsp7YMJyrRPwqLRmICv2kPn1QTd
pbfOZqJOCYBiJqnDqTE557g71Bcw/+fzw/W06/Ohic17QD956m26kp2BP+7E3QMs
8YZr+D8dS3jfSLm82radtjJqsVlQSbPhdjlql7y6nhJNsMDS3mLIeJxCY6YjlP/f
iuhxZCOQKBAh+tkFINU33GEdFicA8Sj/NW0H4MN/KgbdO8li92dyAvZxljGYKmyy
wTLjo7nuxgjefLUHFbXbgEpOVQIeTULC4fryqQdcLhNXQD8TIZnnxN4aZ3vDvyMm
QgHpa3OfEqGvxWZeQWQXdPLQc2/NZ0KPDGdh/2SdFrQpHivnjqpJ7dJ2cwQOt0FR
3YblS3AnS/jhFHA2bU2frAuK+e9by1devSDA6vCPwZryVrevvlCJrJNr0io6o5pO
R1Si9KXrMj4JV4UqqXaXQgeZZq/QyJ5R5mKHAhEgyAn3ndKKgsjOX/gr0AchEmKF
V0Bgm6iz5ZRzCFjih56pA9NEXrGxsZyF0jtLAaI4Tn4WgD316epbjVAw1UX3zrjq
7sk2pE0g/WA6P+FtRr2dN5J0r6w++xLwBKupwIKI/GvIFx53D6O7nQNziBITYRC8
gmNpq2taQzFVqDGZkllJqM/5RIRXUlCTaNTOO9Tmjkr/BGdZT0ML3xlvHmEiClqG
Tv9H6K9eeTfgmtWoS2XliLRv2gVcKyenbQsZjZaDko39l1W1tR2iu1GHcdChjLx0
cEuxAY6pRt2YUoV4AVD4R4eTJ2KVb0moqIv4qpzjkSs8NyUDAPEODXqS24rV8pho
NlpIKoRgUjk1ry/ywOpaoK0hQ7xteHZuFtOs5gi9ZHiVukgoLJCMCaDYN+qzr3D0
rgP8U2xN8LkG6kNLq9uEWJ4bc8RLcuZi08RJjyCXmq47JUfRFkbefJ8sP/LyYRnH
VaVs9Rx82TmtyIuUXJdHEgInEIt/BaGj+pcS7/bycWMBP73r+FBzLPKIat214BYg
gPAYUgQ0f66h3N8fA3rS5hQ0RI65dFqVpk65wYvOcQYR4TfFeDYZZIyaQRXQEtp5
X+TsxFo4ZhggVchqB5RKHGkzWulV6yN9lWg2Gh+GdI+Gv4n1wgkmMKLzIH5+iYkB
lsolI4NsjpbW2Udj5V6kgf+hHzhwSe/FD9908l0/BkqPgeX/kzusxDv78gS6LZsU
cjRNP1hXIE37o12dmAnNpcK+sSJZYKR0BMC2hUCFCs+dfZbG8J8AXi/Ofi+11SzV
/lSbkjn1IkUFLomauzeTg8wl6gJn3rx4cMm0MLJ0OPLz4HahiX1MLOdxmBlNHmy2
XJqGD7zdO3UbEZ7JGRf4m76MyM6YSM+8KY71a+XBdt4dhsusUSarUVKoIWs+d3tb
gzFDwRvimoBgEam1Qe2j64ZMl7oBbQfGqfdlO02dTTpbfjWZMQIQL92iVyi8EQhD
kg40kkyjE5g696wZWj9Bb3xNQOG9HQUmlgpNEbk5TTtiUwiRIuPOK5558n0SXRBP
lLCJRc/dhKXEeOt7rz2cbpG/UvTj+E/N5dA3azLENxr02nu0MeGmOXikmfla6AaU
6Y8gxFDoNSHH81GeGfvjfeTDN2M5dJwkcs01QFjXIT9ydnGi+kmlXVH28nbvL9W8
hEf4FMEy+ZRSD7vB44EdT+hnhRJF+vOgbcHdSoWN7dGJkOop7FuzAnavh+DlHxJR
ku26Rt/EhtHKq2iag2ntMcjSHoiU/TLAVY/AweSP1WE0WSoFEVF2g2mnrHpYzOuj
JPchlRvAQus0qt3yVm9D0Wob/9/st4M/XJA2zL3Tn2ktszA11F4eM6F57jrFYM2s
rTZ8ApaLznxK2zACbl6toITjJlMskzlChYKJOHX5n45ofqcoq5Eg4nCtY89r0Ci0
lrqOd0LeYG4HT9wkLj/DoeFO/DgW8bRhaGilheBSKppNcILfFSmngba8vbRR/Own
yfRNT4uvTKH5OYvsDXRMSmiQqIAzKRWKs3bmBu1Yu5CRwCQkZegiOFBfZ9w5Fpeh
i/0tumaZ737UrsSXsPfe3+dCQQKXQi13TKG4wbK8aXDz69ewStpeCPuyFw3bF4LJ
gO3kT5SjGMzK7BKgYK9C/cMCR7jvhdINrULjohkx6+5RKDasIn9BPrRT0Pd+e6s6
v90y1F91Ey15tc1UR69FjYGhArzn3lkbbXRKJ74Yrwlf9X/dzRSTj2kNZc66O9xK
721DuD63nefYR0Zwg56cqpRID0BUzM5oNTnsG9wNOyuctvX62Ie7hDKb0waP360c
wy/HjhQDUBEXJajWXBaztC88KYeyXgtSmhj38g4TIw5u1Or2LqjAYumYoPQAhLf1
TP7DuPbipfzhv0XqN0KmZ9o9tUQWPZIvp760i6LX8+cGbhWserj66aKRuigndIKX
uosWZ9zkUvH717iKGAgfBL3jtXscUnh7J+NraBlv2mtDmHyhOD/sZ4RNXQZeh4uS
vr731IjhsaaX5gcuL/NBl+5ZfMjpfXKBwJD8rTaQ0O50YbRH7xUSNpURbP/UNVBE
LGfWU64OT3FojuPdlDsCPPvcOEV8f6mQa8rVdSZ++ArrsXE3RYi51bv7A3O/FUAW
bmmr3E3ugoos1z7np7SmuxL7nM671Ni+VcSb/ty9bqt4BoqvnpJt7Vrqpc5+JbkX
0xHAOYt9RtitsKLkzy2k+ayqgeN+9rfTt66om5BBuWPTN05+38jeAXD5J6R4EBBE
YFTrf9NBkWAeL2lyzK1of1ifD3oX9Njbk4lTa6Pk4F03jgzzlXvUeqIqAb42EzOI
ANYILQRZHNCv9iUdm2SQAAaNPC6gX8dS1IQqP2XXiXuJHw7lcXWbtTKKVMJPRI+6
WztXcFCgZQTfYNH4lbJHIqfuxSG7TEcPXEWexK99jnlQY0oJotNPLrHHYCemwH4T
bcsV8QiFZJwXLoeL7A0ypYVo6tzRe8NcWRv0Xq5QlDAW6povGwJ/wf8CabVL4E8x
oBu09NOvzQP6vZPE2/dahkRZX6FmV4jc0AhyGnZ8H5JJQnGTGwMb9jyD4DLXYhcV
twQN1ylXa8zfRlhkAEgtoOcouoxK0OFGizFS+Do1lcTRcCTI2aFMkhLRut9FkUTf
vSQj5aGE2z8gDUWLTyRYA4LxC0JlW2b3+mV0xOaCjB/keU+MnR2TkUAer3YL9Dpa
jEARl3xbd3LQ3/VgWgiJfp2HzLELODAPdjceMYm0u7Eu1NIExuwqHkbsTWa9VpBL
u3Ju0+H8c9ju2eUXpzzOLNQsx8n8h6r6ZOYOAa5/Qbyp0X3XmULmb3CHLD6En2z5
gNzt3SeGdZc46GqdG5JILztc9w2Kh5+nGJnse15kj7wjc7YwY1HAnQsoB5iZOyzw
w7bOoz8YS0BjiJ/G8ozLXWFc7M6yE+MbeV5UqPBxunAMOLcLk2HysfVQugwKgf0h
2XP+9QBe8trigY9QDEBtp2ifc+N90z+25yFXZw3HqLAWZHSyXhodOSQ8GmAySUSH
q3UmET4nX5FOa726ZqmrQHV+GYpWqtCLHwS0X+GjyFfyza9aKAkkIVleY1WRq60O
Il1/7mdPnY5uQhfU4ytHsv7tXfTo6GXmn/74ge6VPJ6CQ15n96Bgmn93mukxXQJQ
fkOirJ0LvcxgKXFa45nQ8Wd4AurjUQMzrsL8FaaybJBZ0jFBOU8G8rFC+vIYGUo/
V6bNhZ6CxGkGTTQ91sT/X76QSmIpqQ2ZRFOI3cVEvLUCojIAvDesrIAd5hSTcKHO
g3eM7jfB8YRpt/awFkANa+RUotL0eDkVtefHjWveqIuOVrKNXDqUlsY+Ei0idDVX
FRDhXID0tUTLuniA86tBwgMief45ju+09JnxdOmenJGxaCuZqt0FjNgURC3rvMg/
xaSOBzRNlUmh7bP4Bmo4XPewiHAzpqfe6+FXENqv4zVeeq1jE76x+h/OqylRSSIj
1Ln/SVBwMs66wRXgjNjyvbAcqo3TBNvoVWfM2ghEbQCz8Ds9C0o1nV/bMCfqA4MD
4NuBS3vtAUz7ceL0dCsbW+WSkSNfCnA8NVGDG1uubmkcdFhvnjbgk0S6DieqiOVi
uPTvdBnC2kjA8GSeXNZNbsgDSp1YirNlS/exRpUjkE/QEIWGXjkzBhEzHAMf9tq6
9kWeSRMtdKkib7PK+2hbpXLW19aCvuYdsnHS7HM8ArriN0DzcMiiuuzUiPfMU9wJ
Y6+SRjgXLLaYr660NyCqA7qKrSfCzheeCDNKSGS1KLy4NuPL84PcaZI0WA62vGMS
6gUl5DSnqTKkkweyxL0cMnzoPOggzflESL6QP58mlvR7Ye9+LJmP0w1jN2tcPiEQ
UyA4U/meliwL2oWgVR8pl252LwFbY93WW4BVjSvEIj+2L+I3sf3mwhUwpY3u8Hvx
sp4G5jq377NEpG4HkmTXDeWNiMqgvQKvdlPYUcnLNHR3ASpNrGMYZ5ziai3fP5Y0
H64BXKVHQLBZrsNsDqhjU5g7Mr+YL2lfPxbqYWKt7yxDKZ0I2dFa6BEjpQp8eNqa
G15YswikKtc5GfW37AR3k4RSQPciNdxY/avzPnzRLJFYyB9noXn4Gr3eU27I46Ew
XwBnebDWucLa3ucCPJarw4Bfs/EIaXV1R/Og97Inr6jsKbC1Iy1JqVcZMtkOXJR0
FCUw2wN9nfxTxzjg5CTrzwbkJgnEdQn5H/JebxjqCL11pkH8nim2yCYkVeN4Q2SO
IMqyU6AOqz0mXeJEV94gZ8zB3CgH5nHYUeIvywvYLWmbYSRz99U8VWHgJEPNUqyw
QIYGN6soGVssU9IfEu/xJa9hg06X3MEG3oWo+9zBdU/n+j5XDZ3GPJ2CsQCqmfTN
stYwpRyBjq0qWIBEIm9ASm39STS3goKzbLEkD4/SE12oSyjLC3G50UqdP2eDlS0t
UNJWeZCmDUmD+/DABQEZNOBqA8d0zxbUSv9AqGoK4Va99AdWRcKomdD5QL7CQVk4
rFTemt6bbJvmYYxyqp+4lH5N8WI20QLmBxJkYP/12eJZxtZTp4pm2TJw/vOmA+hD
CuaOa23aTN9hJBQ22B3E9fRsZJkMJ/vdPK/V4Y4OM92VzMKxqxHfHhcauUy4Iq/4
lcjX72NdeWKVUxtbB5/Nuv6ac0mFgdl/QkSP5N/0mNNspnpn7ppFZsWDivSG73D9
aFqkUxzTNLltBfN46E8l5pG9sGNoZk4A80wAPk8XY2bGEHl1y4QS3Gh1cpFEEMp6
7wSy0Q4SvQX4r1bwXinGQrG9n+gSmz4wUnN+7vcrGJjqb5LIS5XeXYXMg/xkvJJs
s+O9XGzFvCCpy3GkhJI7SxuhIg2O4AHLi0J5NOYYVD0Kb1GsEJQGxb1gjVJop2Pi
k2aPr3Ol4juICd3karmkYlZIoZEBI7nbgCazcOXcChKrgm98yVGo0QmdycFcVOXi
i5sMlHuK6rMOl2T0fhK8EEUkNXP56aacpVWuHXIxjcLNdtUquiwaRST+sEZed9Up
HtlN4c5VKlrc4k28G9aUCr7QDGl0QG7dAszrdCP+wr522tq+BzxP/FjtsbjtX+1m
UAwlOhXVI8t4IYAp25mVdDjjaUHsJacLPck1JTDqeru+9nntS4Ym+1ghIH2IN4/l
rAgUdoWsZhXasBLLQKo1eiEp3avfJ1TpxrCeB/ANWow5XNr/8fizoqLwfwbELorN
2h88Y2CUxd9ol38DKnIq1RZf+IKHDV0utrpR058F1iy5jIvysn3hL/IGYv7cSfwu
xXI/UJ/8ZZWEfewUhXWxA7+4BLmU48WE3/GERVeUZVkUesTGIepoG7gABdrVwDRQ
iMFjaQcGbym1+120jDFpzsqyiXP6T/QFU26ddSJAjtl4wR3nrwGf/LrNCax3Ugwi
iukhvcFanxsVBMPix+1wdrkEtUfYKAWPa2sgMDnzS+2bI1Pg+v06DscWEk5dpN8p
EX7rXK1CaFoFHztdEdvEWk4fj8xuV9i2yZXvnF8AmNzhHLLC0YbA1Gw+KzT7+vw4
5/Ol24sRAtGZ+HaoTjTa3CN5UibJFXAh9d8NW3k82e1HMs83fm8VVsJ0K2RKwGdJ
4nRLSzFb3g9BGleTA1vVR2QKXafrzsI+L+kpgGXC4imjMGlSrHkxPd/oL5jLuwFB
DR0o2zOtNo4VQnAAXNLwTkdwgA+llc9Um6GNR1YaEizUHD96ONEDi+ZiVmw0z9xO
QYp+Vi3LbqIvlUv2pIi6EDRz4XfIRQaDGExIY3e+QDLPUrcVWVazssW0DcKF5mAT
mE0b++69TnshIMxIqiC874XvRE+Q0BnTZwNQaWzewXWYn9iWhLmxtGHPMHE6b9zx
+ZEkrVY5RHSpf1xBQjwdcf1klEWkdK7NMGj0VLSuXdD6nY2xwS0E0n6YD1C3ZTgl
6nQ0n6APHFQLqzeLufhClPQRQxBCqE8gFHaUdoj9OabJ4KNpWXM/LY64JhjCTxZP
+t1VpTSepZoMrYx2IdL3cgsTSIF9mnT5KhdN0ZZilVtyU/5iqVzAqTP4nB4OtYD2
1uebfISEjHP+ZI4cFhnXi/gxuqxWxcv1ivxOl39+bE4SH3HOqEbbq96IIlB9Tqb2
NzpEL1IMlNw2jEbWbkC3m6uqxeFmYW7cdiEQj2euaVheR3PcDU6DWkK5v8UbtU6n
cuBtUMKcomMahB0FELQ/IWYixAdL+V/ZiY/qjuPtyzWaxkXUWT0bcESHUjCGOFM5
9UIAAwyL4GWhAC4iKpeWjO2neBT5z2iO3GDBtaCtEnCNciidnnEidH+FnTqHfStl
m7XMP0oeGAoE99n9xJnovckd+DYOlfrbeZnoTKc0G41PTvOoR/9M69gRDzECrHFA
6z+QCM3lR6AW+IAPGfia7vKiRZ8Meb1RFOYvbaf192EQzmcLvqXSGLXzbO1XsjVH
i9i8z+rryiTGa4i+t/s2fDzjaZtQE+4tRuZ6846YwDrnEnkV2HOIxOBw9PjbMEGB
Eb6ZuC8OUT5dcbltnf07VE1f7OkO8SGVcqG6Z+a+siK24Nm8xO8M3SaO6BigayUb
o85D4P08FfGa+2TtFkgDB3tiTWC6dfCMfb2UxuN7xQX1yFsvLG30v9RszDxfV4tk
UqT7DeWc9iRqz8kT56erZMdpdNmruQ8wGUq5nczxfoYH/Vtq+eTrTAVhRQDoX/zN
z458tTVTb5KHbo7aEsQHa2etKVuhHXkrXJhraPnYiZ6iIvcYU6yq3c35wII7WrJz
rZ/oVGMJoDmSLUY2OpE7ROsmNNHevUgRBhWyWuqMNHc+R5d11cScYXncLypNi4M9
HRcE3spJ8gXnDmPs3n741dDDjFyhQRixBWSKmDaT/s/CBo++cXkYu5lE6DWnjskt
Ne1eEct2e//e0rqmTHkwkPLqIaVsCzx1sHakuwSp/dbK1FWPJzyvvG6pJxycbfxB
IuGd+Di+uxbyhgt0So1cGSGIWKSkgeZEF1rqo+Vkjvr/GqV0WoI42HAxlfuKSQAL
tzBWmjjaCIt5AJlzVc51XWpVY79G/oU6RG9Wjst+WSs9HKYhZcZTWaa/L/MTV3iX
QI/qKDLQpuKcq/NbC4DcbjUBCnWxC1FXOc0SeKDhpcLakvj8eKgBW/K0eFEUZbV2
JyW8KtNWuMmzBxTplE9g2wOSboYIb9snFIxyrFkuseFYB+TtAwbwyXaacxCq+3lV
vhihkEX+N+rDAVdtPdjeua2KC+NGgaMFChPsLt8qEnLHRb0Cak6Q/acfmpkPVTjY
h3JBHwSkHJcxsvWfeuChe0eZcl9FZQHCUNBpcBy4RCZo6PSRH4b/G4relJs2YlHc
dQmHfGLMnJAJB/4kdHmKjxHp+AlFODcWDno2dRifX8IeL0I5GCcQ8zQD94qEu0rr
sSKNr4/hnRVuguzqUrw27+vBzCnQWxz4lHj2EZ7hLPcjIXkvYHF3C2Ii3Gbd4Zhj
p0anpjKUJaM6NJWTBG16B2r9fZ/ovIR6CzYMIz1nnvhCLaWl9moq3KOAv+DJYpKo
TbkChRrv8t8m54VaRIezKez0cPARvl7hltXhXOVzU1PWkc2jIiU1LGOs2UUgkDkU
pjHgrcKDMW6Ms9Mv/Vub9a+PBQfFugSQfWKrEuBqQc2xlX94dCZlfZKsBFx2sYmV
fDp95HwF8JQTSVTHI6IN8VRzOzhmx/UXFDTu3Tw+7/+tbJFSiEJmKHwd8PUV5cgW
7YoWjLe1o4V5R74sLq+3YMSfhkNdraQ/ykQddX1itkrT4VxuN8HRljhpS3H++NOX
jnFAbQ2FgAQoqRhgyUv3FomlVhb+kpxAhvOnEWanX5pQO8BE08I+2ihD9BxWN/J4
rnRkyU1QuY2EJztSDIiRi5kXeqZJlU0yN93Y6bW2mTGMTNYIFTG3YDHlv+ShJH6r
xtFkrxpKc5oeMywcGAoVmP17gnViolppK1TMhQ2P4kCTn5MAXgmAHBvTYD0HzSAY
bog9m533Chpyq9u3C9wWSdxHz2k8pvc58JM7QeXLk41l/J1oDatt6rlSSJMtuYJD
7ljad05jYcnEwYFKldUORsfUobTqSctVfDA0JDCpl9Y93eDx6gD0FfnY6pytPp4T
SIFX9BI4vB/COTJtO/jUUxwEZpN5JWJI6JVWGUETW+14GO3opkWhOv0iuJbfUHtX
izlaB/EYou+x0taAgHCKM5SeFeH+r3dVkFHrrIrwip2zy8CeY8D/be7yr32g2Wlg
o/E8PYsbRK0OtJQjd9NmGfSP4s7tz33k96xNpAVNtHsdCGxThER8/04k/jiRpC25
1NjVf3ZjdKaOLTQ+XArh/7m4SiXkkeZppybq8mH/JsYlMx6kk/DKOtBjcZJusUBo
DWdGJLo+zsArNb5FhvxjP7FeGfwClEBdF65nY03rnNDFvJCQhqbTsDDwOvM6RCLY
FT1cOtwTeWDfuCd0aJPpbxMNJEGRdoGKxJLdhO389R4BsvINorFTxva/w52epfSC
+vDJKJPCcmCrVm9hhDqhrYD23WnePmj4hsfeIKdN4FS1NAe/munyw2dORGVYKaMv
YDGirPkDXxik3aLNU/RFcIsHZHggVrwBtBoV5DQ2qTcLNojU7Aw5Rn627Ka2bd0E
BgTIvn7v5GMCPtFRorlTWiRf21MmD532BuyP6X9DaxP0/wccc/DijQ0sXamvXJKZ
cy+gRPetJ/dd3aj9cQ/gJ9a+3iUb1aofMjuSM9amui1aKoUBrJsB2SH/kPpt0IpS
8mtiffHWdvuxxwFjA8pB6HAjQ15+bIIbkoCPSDl+p2+6Au6zAs5kOwibRDtcHNlr
uxL6eH875LDYBC6z1GzhTOd3/zA/oVJIJyzLqEWaNmr/dc3n6+o0Pf0nTT4IGojW
gIsu+5MfxCAR5+Wwe19iY48VuUL5QHn+dTZvWqz/pMeaBPDLkLiQdXpgCplvotGh
NNuqidoKqmGyyeJLZePqF1bF2Sn0tdm1Rjiz5UCL+iGGYF6NBtMev3BvxbkXPyIH
xf+ij9gz4gQTtcejnr8+WZeuI9WTLjniRfzpan6KKVdND8CrcYxo+y972yL+RYab
NQ6stUEDZf9Wd1FHlFLUtUtgXf2k1mBDoP7uacG0fojDMFEPUwX57PNM14Nrcyt7
OJOQMOOfM+kbpdmfdnpOeqvrE5UtXidxD60go05k4wOC0PjagUS8eFoYB876yjHl
VT6ksyOUlQwFFfjPyJN5L7eVI4jj6UCCbMrkLwC5iVdlw9NzvuDAzN3Dwy9LuD1d
Oc5i+ytHszg4KOGDHjN68azMvoD7WrbEYw26maXHCXO4s1t/Dea6F+ZielaoOK3m
Xop5kwdvgM4CSqmok9iPzHOe+CNqM/e0eYZTltJ9dp+oSHwy5afW18Ch3cOhp+2M
qzo+j3JjINBw2DOkATkvW3wSoqwX095lUw0ip5iSyJMFbuzbyZgLUeetNotn2NnK
Vy+U7LvBk3Lg9uW57DQIOAe1yDDh1I5HJn13/rHcXibpxe2vET5mnKrAVOHV/M3W
UDjFpjo5MRk43EPi1Liokmr6OdP87MsIdG1AeGP3mtIyLqbMdvXxu5T1CcqEabJK
NdEn6sl51lmU3rsuGshcp0MplUYaZb73Iq+pzUOOdwE2epBX3kX27HM8Ae2seI/w
Q4R69jI9LUbYZZtHtapkXFfzkTB0bMnZeBkdlAONcHHt371fq/Zh1UTWpiW7iLNK
MemZj08SfDE9i/jPvjvg2AtsgaAc47azByJUfEcEL/mYiruqgTOxhWCs9Ny7eODW
ck/NfidtogrPCvo442Vj1g+SpLMnmbgP8hneJQw4jLJK3lDBT7OvePFuF5KJB5vo
pE/tG6fpHuOPmQesuGaJm8JrrQNTIczBXvBNl9OoSncAS2JpG3Pgb1yBVKAPGki+
/w5Ucf3Xx8edB06VYYOLWYj/peepjqo11o3h1SK8VWqkBH28zE4I6eFiZDvs0P5j
sl40JrgI0caVLUmswnZZNGnhKIC5ZpLWPXd35dJm+26Ta0qErEG3EK/9tfQDIEwo
GWP1IMtlL27N9wq7fvceIrHUOuLoy7smOAfZ8uE7aTppZFwPrYh6CKNPkjurdMvj
4D2DP+ls6PLRoBk6P2c1t8SZunC6F1zJdgLiNGV0U9eDn/3Bi4agmh83Ht+9gDq2
WIN3oqsKMs2TtDvqHDhpXhJJTpVuFoBxijvugrvWQZGOK824I23vbCLSASy5yzyk
4zkehgdCLiao6DAJMLp+b8dvjR6CgXDQ346Mvu6aQRb9bvg5sftYruF3c78+CSm8
MIA4rNndvlcqUIsZ4/xL8L80Yslyd/BhkemXAasQLRfFRsYjbkDxyMzZNafBtk4e
qk/1PjSKjd9m9zqYEnl7ynq19bsZfbtZGy/aWDaajGiXcg5wqsSMh1nCCzq+doZC
7BXeZDTxna0yKZjRk76kdNbUhco60Z8dcyBtBTS2bXo3qVrq5tra8lqc67zHseKq
umMDmtGu7JB3zB0tCiJptc7dKb2l/k+lwZlWLvCovk5tnzvJ9RhYtHNo+pZyfD0C
4rEzfVEW5XkZSYRbo9ySuVINAgXNmDDvNqT/jJAuUswnjPpcY6EFtyRHRvWmXSZG
8d3L79Xn8VICIXYdR1TqQ+7KOZNgFzVkYM1JJFq+aPyDf1lSBN8bdim1rr1QjYtB
jkvKmRmqWf+ytJDXWpVy5GWIYB68xqMcI9nkEY1cu8lRNUbwkEgErDqCq1hWUhbs
nVjx1K/M7TN0M/XoqPUAE+TdJQcOy0s1qegq4Qk7PID1UQbhI6mlPcTd9kxBLNM+
Uq15ZgvyT42+QMOMEutczjTld3YvUKi3F11/95V+jDDUKl8FjTd5mcxFUehqbv1h
5Z49i7dfuTNI7xWCi2S50/wYTdxOyvE+8zjO/3I784TDbZbtXJTzXGXY6SW71/Tz
plVEBtw3NnkL5Dch37iDHoRnBcktHcnnrbmWEuVSXsLNpRtfxsD2aAkUeH/LOJCj
5Xy645oB/kSnP6HkliO8Sjbo3C1dDvcR6lkA0GT1X4ELxGLbqI82woi4/lCn9lEO
xQ6RQOw448ooN+v9XG8ef9448XB4QMxEqv1oeF6cIOJm0NE4Ng2PBnk7vGrY/Dq3
llAJqHu2IzCMwNyLjFnAJxA18lG+AS0mZ/0WCCuGtTXKZTV9CBrielNUvsS5pfSn
8yuUL/KbVS9nDJG4paSmM5JUogDfPxVLW9O0elp25xS7nEweXgqme2B2y/3OArW7
0+JUkC9K2mkx08qazmUahE4D2p5zjaXOmVPWCBIab2sM9r+vkOV420IhRO0adXMo
8iGb8tAnpqLnY863zt8vNL24Uj6um79KXDEX/3gvt5a5xtGqwCBD2v5VzAupHage
fEnD80SyGzlL0+Asjb3CxpLCjKyXhzvVqZ9ckm9cr37kpWj9NQv/8P9AnxvyBFFe
iCI25qFJwccTBBQrBzd3aOAsM2+TTaIe0wL92ZrTiZ8282cp2gnweakJ8sKt7dcS
wjTsaQNgdhM8oDuL++Ho5XuzNFgS7KwGj/+O903Ypk6yvMzZ278KFP3FjaOIFPgr
1zmekuhYMPfmlD28eSTiWfIkTwkoQUpUM9ewmCV/fk87mHmmPaFxYeOoiVBAIv/C
ggjrsxbKwTsOJOaP2og+I+Ej1LbGJRdLdb/Y9EqLjwjCSg9aRxDzC221aiDqgcaQ
aPW5gZoS2S1yGCC85a/xTLHGYPcPJm6+IfnugO0c7edbNLkgLHRHH4zbsCOjlX2O
D0DiMebgtbF3lHvikklBQqJryY5w6/Y9LLAVjI4UBD0f9c+Iq/Fufd9MlbORlMxP
LAsQIw0egO1FD1G6g2P1ttrhlC77RcLfOJ17q6Ty+aMk7eVPFpDhQAX6J7Zbwcvn
vLd4+s4xi50LM4wgjQYS03qQ054GuiZWU76IYWIxStObtNdq4nioc/ZRtZ3OwU5y
uX0Kkffwu9OOBVPksciUlfofYDs9kJ9RkjrvycE59zUUXZAaO0AbE+Pjry/JZTXy
ySOAANlzS3AcsFe2jsT1undfHDMT+iaKaU3ZLHG1djVKUsBsvxq/VdFHnw24laFM
bscQQwYeeImev4aVIXOuDu340cqmWmx9iP1aVwou55pGD04W3CvRS+iQfyqoYK77
A0Qg0uroSJyulGSkZqIjPVF8OM0Y1LRo5NMc6nLmSpTusK7Ffk24T0Cdrvu8HlwR
62Q/XmPlw8XI6Pu6OgYwDudu0AmYQWLOzcLOU9x9nsvQT4FrleJuxd8qkA54FcRC
aibzbZ1aXtoSnFBH8KkW2qYNEmLgAL174k9J2EqyzdD0pM4H8hv0WoBCSf4zBCaQ
JCrauope0A7WJMOeFHPhAIDIpbaSvdbwIEImUmL7Vwe1KJeEENFv1v6q12VTuQsK
IiALzRe7TiQbm8HBtBIHmvuBaievt5er06Z+l0gDpJydCvLevKa4IspBfJLeYYiZ
Ogyi4+GouFnaju/+FpB7btOSkwEZHMTcITV0WvCsH5FgkU7W5lgDzcLELxovyJs3
w3G2oN3HhIc3Raqiz7p4PXLBSdY0hLifX1ImY+1QroTYgDbow9Lxum+j1PEFN0vw
0VCql7kcnCMn2sYUgD7vhmUno195Xu6JWANaU9ANJZ3eyUUnW0k+HwkWFr7kC7er
MYBV7FHhrx18xRi4vx+9ZPhKMkUf7NHtbPxv8edj7uL5tbvcP60dkKhVtm3dctRz
p0OkAj9/piWpiNH77qs6KAEPQAY25tJ5Q0Yb9ZEQxWaJzV50tOgTNRQeWXRAANMJ
ViXWWkhmu/4lzYJlBcz8IC2To4+RvRzKNKN6xqlf8OmSBx1yvFgVCP+CTDC3Gp6m
ogQJKhJ2zQ5xKDeSMhVdvmBlyc1Ig2Q/7J8NaepQUucE83pKfUaoJzx/6iADI2RX
TYQSgcpD8dJ8VyWY3AOA+iWYwIY+TL0j62OLN7vCGdNB4TUvJWogcbksKMbzNHdE
znAUcLkID5qSX7xTNmjSk+alk4o3maRmtiftO3Yoj+K5w5IwblUSykXQpQwGfhwx
EqbugLE9OAwTco8V5zzKV9VIq09su7Fl+Qc/+lRbi1CGazPUypX8G+79BgpETHfZ
dE8nQbm06vAgs3IVqkluZ+rUF/9hPW0E0C7mSvRtI6zUOTiWCeA/mZ0NmiGtCm2H
JJ/3pYPJpQUVK0xu6B12riVdAZl8HLjK5HCKSWwoPeMEQPpaTh7baK2xIJ5xXzOD
fSIj09X4qFt4IenlC7CotIQlDBG9qzN4KT9WVXmmvc7Hn9+XSvQkrfpwOsYfoZK7
5FUgGqlg3RU3wuxAJMIzo1s1fSJiA4n7BXqufEXl478JEwq4mlaoIu7F0yXzyA3A
1D+OhetaQXYeMqYuEE1A1/MkILDH1ZVeKdKpIuF+TQIzAPUIC29N0EvdReVquADy
6RvbNszrFPSd+HtZk48mVmRTbwqizPTrl85rpPj5zxJeaftCP5SssyHXDruAUKpd
Uknf4lMEEW42Y0Q/0fecRdzl0W1wtwjXAtA7ve3P+qYA2KUGQfYTh988XtwzN/cN
tbUvZ88lP3yTNtEzSdRZMPxrEK/qgbSTDKmiJnHQymRfhDm/Lk+gJGIgDL6nrYII
hQnnkQaHzUTG3e1J6fBRJD4VacILkeuAjjWByRAEX0sb//CRJ7x5AgAlIAYGuIUf
/7RhKIWaFuLJEXZvDjV56NGEg4hYGelDqFnvjZ3HCIf2g71TiOSjrSDSTnwl1say
B43TtHCBEDdshvf4ry70NQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
k4+hPwwozLkIkWfTPkFKeJMtJg38RmkrcxiC9qYP8vRTRP5v6CK+1HyVB3RA+UDx
bAzgTT+aQYp5SJwv0PNrc/fg8Owzr8yyRnsUfp+Zfwq9PLi8cmO/Vqd1oMs3/t0x
BBwDdVmMIfp7Y6EQLlNAZCMKEbfFrItPTiQdFOxTqOkLuAYJxujiH3MjpP6/YpMT
ijifWm73/kB+6jvcUdHpCN7rIskvNLatIZiNpbNoyJH3obPsPWESc7ZVWjFXsgaZ
4lGpJmdzLOs6hnS7gkWkGE4n+YqaoYMn0tHV3U2cI4pRtFDX8G0U63pfrPLxcNq7
WGh1eL0TgmKN1NXe9WgIqg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2864 )
`pragma protect data_block
iMmfwX83e6h6WJ/xzeN4jFhvRnUAlh3b2g5HF9Fr4f6zQxM325PNxyNsF1Mejtgp
9VjUg6M97HmRmMxNpA/o3tLc3M9N90zBeHxrqpb4XdTeggxfj+Um0HdcUKuYKdNJ
PVz5GxEfh1TMDUPO6HmJk3mexkfaF/2U91BQCTPIMrVoGPQMiQYGwI8x+nQEurH9
QQIbwrtHndwXt1SSWhuVD29OaAkecoX1gE+Mgrt8htu7pOtTFgKlUKyrxIzrN6hD
bERNk3wDt8tDlXdYDrcJIpa02SZG6eXkNgD3IfDGQZKyq4qVr1yBS5yNGEy8lhh1
V01D4EDtIl1vaNtJZ0qdZwXvISa6QMc+PM4uSx1kXvcutTBvax+4ImoJExnc/uC0
xPmSgEMRW9WubXbKv+3SMsXW2qYCGM5NqspOlMabEtRskoAQVdGOSR+LH0Q6qoax
EtTQj0Mr9QDAXCvYvCqD8WWFNVJ5Ytc+Fm4rZWF7ALlxz55WBDOg/Z1tW2D5dXor
Vb27kDxgz+PbYD7e4wwxp0z5krWeNGhcBtJsjxSZVABS0NAR2l9EACJT9djrXxJX
ElWvL9Mg1XI7hov7I647pDrx7Ze88/MNwMQx44Blzwqbgqzm0/fxat+h1/TF0TvT
dcHRZyAilkk2Kkk+V852Q3FJjTq8ncmQKdajX5pmq1l6sbgbDX2+RwxVDlyN6Txz
LNEBhjgTVsAoDaA06bM9EQvSWbUbmMqvDJaAR3/TYSy9/Clh1y6tfbCBmlRftswK
pnzXaNfjkHC+KgaZm1bJe227HQk++Gq4WskxzbpuYzjKSKyaXOvVwzM1QZbPUA4U
1F2sfL1akll0j7t9/mpOhFKeYTEKKIRW/gmQnWp7CwB4g2AHCpx/xapUNFP5gUDn
0v7462NE379QOPlE8AWeN55yRPvtU5Xcet2v09e05C3Myu7Up7JULI4/SsS0qqvg
SeWB+G9Ob1Sz7ck8f5j3/NrLJ4JDfCB4fLIKfTdGR9glE6BHPxspxpRa1nMB0Kou
Hi9FI/bBCiHDdwIwjljyQ7XOYC2J0/T2UPFPYXTSf++YNCJWvc0dIV48tVk2GFwE
GmikllM9fZ5ol62QOxUcbjKTWyD1pSHOaealjYOgPTcv1z2uB8JvyfWMcE19TSmI
e12Cuq4nxcPTAhPBlAGQbmgNa+qmnj/0PNI8sV6u95w1hxEkfjWNKF9LUnPynXh9
J8s05MzB3wfC+WVeNMc1NK8SGtOmbbaTKu3ICQYtuMI4AMeFNZJrbVyr9vjLc7xA
lq2cevJuwDRuSM3qsfOY3akpgqevv5gnsHAJn23FVOXyxPtNLs1F4uesDUckL4r3
QKFcyYc/QvToBl+0glTguoO4nF5AJu14dzLOtzGPyxxl2a7GyGF1pLLTu7b+j36Q
x/t3CdIkracrUe6JKkVen0yBpgMKWBfWjMgtxHG/DhlBs5a8BD3+Uq46AlwIQ9zF
Ws3B9+Y5xsfT6MyYQA366VQAMD7b9zzdtny7+XDLojS4EzmFnC7y2riHUBrel8/0
duKT64FvzZ4W1EE/ot0wGrQEgY+2rfogUfnnH3bAX6bp/Tn7f2O4HkhtbMvmnX9U
6Wydd7GQpYpt15cKvhXG9bhZppGYJ6SH/vS/CPyisFl1QFkPrORgFtDGqZ7gMhFp
2vegl2l+5PThwYYA6wjqDiiFf2zJE9XaknThowT1d37NVHDw54p0mW/Q0CtuZwrt
rwQ9S9HOk4Z5iwf0xe2r22EIzpbCyDJJU2hrMJRTBmbCrMLNPYGwDAhe0VArZ63d
bxdZVzFn3Qzz2icnWp9S+CnZ4nLui+SPaBX2ZbHhX0ctRO55Lg07dRtbtDh6mLKr
bxdGiMLwgoUSpTGAHApJbiyjPnTO1/bNLQNA0vVdJYWMJJ/LEN27eBlKJEm/79TH
iKCYQoYMjJ9V7NJAd2IUW+ZmoZofVhiTXtO0S+s6g9diz8nEzxkJTPpImF0du4Kx
r9Xm1f9Y5HB8QGUz478Sari+ugODzbfAhz6iz2Udw3bhpmqLWaCpf+dnUK29LgCD
LQDPvumQdYv8vbYwnq0bzv7SQgcod1FZLyteEbL+8AKDBp3jn7ye0fQT0KhnpKfn
/YRN3cyQlcE0g77tdREcIquycy8SZMNceot4DZHrBZB/WYHZni5sKQsaiJW+iiNU
SwOkEY6EYD4Ji/ulKOldQT9fMRhQuDRHSiXju6AElIUyZ+RI8P2pv8XT5WHcfOvC
LNSGzBj4hFA7893QAE3MjARaprzAx7cKtV9Yq4yfByTSOla8aN5OTRrV/ihfRgyX
khH+mpUtXSQZfDRn7aYTzsge1uWh68YqkyW2e7qRNAeRSHKkCKINDnU0XGlCUrHi
ZEgknA98r2ZQvSNUXrDSSWb1jExG0fUafqM8tSKAZAgxRyiD/IBYtpUIbMU+5yud
Z/zhD4tJwHuIq0RA/z9h2GG6c+3xJLfjoDQyFFSCietsrRGyE6dkFwedKnuMrcW9
2kQ/+PPfsZJYt0YD2Ml9bIPocuuQsyKU/pAX7aLqQlDPqqyxWvUzHDdqIKxBqX7R
MkghNm0HhKsqrFKHfLFzXDzOawQEmgd6ql54xsplnwvhHlva6fEtg67zGhdLTHCQ
bqq3ZZ/RApRtM9Kc/NWRD7wd1a/0s/ouY8yYLzbcXh95e+L239Db3l/oDX/rbBNP
/G0DNgHBICNQ8iBu1k9mmLhlblgt1xGDLqrbIGEXY/FhkBcou8FZHqEWYCp68NP/
o+AH9QOJ1SM0H8vaoIcvk8VehA/mULwTw8VE/LE3rUf86f/wjarDQ5XXEdnzb/GS
+/gODhB09lrC5Lo/vVTkSPp5llWCXVw+ka92Hv+wk8c40xagQTQwQqHEs2mDq5N8
dTVFB4hq0c81OmxrQiHfQxeJE9hnsAoAWkcRq+0PKCYeZK6+m404u5CkgmSGJtjF
7NVGGGfc5Z+u58N8uAANyATTtSBGhDuxld5BuAJwcN3lQyavgoxoiJqpZrYsThia
fQQInsAiUPh/C8saVAy75tsLi1HrqFNzg/lgL8q+1O9eml4ie95j0U+o2FSPAWto
FmkUSD1Ca/b2vT2+eCcf3s7RpZCwhWcFw+Czpf+TedZ0ZKbvtCYuvrXcrYVD5U97
BaB4WvP1ngoLvIioZShMqOwRu8NSkqdFwvj3HlHSqbc/hY61FQr9Rku5KR0yVrTf
R17eHIbYXGRu9vkxMyWdci6C1zD39PDamTR6j8ZI+25bUV82oYqVIMHHQ+YV05Cs
OJqdx0rV8A6fE6nbB88fSRqK63W+7Jio+xPo//O1Hq/75qTmQwy+NfQJCUYqEwSZ
OFlnp+vBkPmtiyAz7VGzTxLM+modsZ7+dpsq7aMIPJhsqoW3w/QyYUuqMbZiv9oS
3KBAjfMuJ1DEChf+9jrcNrDzNipf/XjyDrtjjirrAj7DXTrjopl6BILLlS+v2lEa
viD/XVzfIgMZNvLL6KrSvE4z0Tq1kEZwJQQqeERXEu91+9hMiQIN91Cga4tnRRk8
qyUifYXi266VgkYLlb6zn8Phe//J5rTxR1UIw97Vp/b1U+Hf+0Paxe5b1DWJBMWH
SZu9hwiBrJv8sfx2WlvkcUr02j5p+kQDibwm1tqS5sw/PzH0PUCepJFIOr0vYgzg
K8CFrX2EYNes7WtRFl9WcNo4hH62QLIafl4+Bc0/wjJdYyrIqk5cqQblnm50uZzl
eWJH7UPIlvpCWLULC44OdbPwQJdsaPfh0TYX/dQn8T+RT2ZCcitUwSRQWiLEYLhf
0ejrdp2hPH5EEEAp+DsnaflRCHg4P64XLfQK83C0erw=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RNNODAuiU1LsZvtcR2Akkt5C+ygPCMmyWcYEUtB2I4VMk0/LqZExeA6oCWxqjQjv
2areY3VDAGOyM10nLQcQ/yvq52CpaiCwJWsTp00Y6X3g+xw1lwv8ZoL0CxC2I2ck
IbqLLPJMk+acdAhSCoerWu7KX8ubAU+ccizaCaJFXgtNDH3MnjCvBIxpBCoFI3Z2
zV68w/j5vS6Rjr+jxAWP0MnLezTDYtaRxSo5qqJdwNersEmZpYszC8iLCwqn7SC9
n/o5td+Ww/mp0jOGB4QnERiZNcaVeTsAIBAEUEJ5IlV5vvHqwedGO/Tvh5zzIHJA
TKod2ZgTzhwThbXTMBy/Cw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8704 )
`pragma protect data_block
fVFAIdwG6x75uqIs4pu2teuoKN5zDGwsXEQb+pIITqGkUeuFj0JR31E2PN+e4pv+
bG3UTp2RB9t/5ToYjM/btei9lPse4/zZaIELrq6a+pGEKOyf+3wtFLIcJY5fbN9o
4Q++PV+mg47gj8pFQ5jv/ZYNw6WJX0HfEYHFo0ZM98JwFo38frLm55GWLP47UyaU
DqX48GVB8bPIB2ETKrIbY1ooNL68fGQ/mb8LWy90/d+BlxyvpUOMPBOED7ikSjtq
/EKqbHOWAazwHGHQnPVF7o3d7d/vxZCeZ1Db5Os1PNmZXrOJKek5o1tqxpmDY9WQ
lGvufBhBXdAwx4QHXxwjIugmNag7WxXq3Cd844faIvwPoUMfwSeaNDqOlMxloxHc
o+NxQ7u05/DDBtM5pN/7LuKbAajlrPr8bBFMHWglDuX9yXWyiU1kvsHtNrRXOxFG
6UPcJ5BgVqAhEIYiTSun4UF7wdZq+DodFqS/861AMbhCYNAIPtwTwXVew7FtcEJW
g+cu0VAWNFFSIWSL7quOtVFFNBmo9fCtzUf0sP5lQ0/cTMUO8ohPkikeEdYi88Lh
CSol3cVbIurK4Uh6jowN1bIUPX738ta+Y5hFQK9iCLxuoWFBiKowWjHk5PFk2wpK
0p7BnHvvQLFZxtKU+9WYAcJa+ku3yOptSLG7spLKIF89CPtDG7EjcLlVL/J0KjgN
Jw9JvtDqoKqcnp1odX0KOl7244V2QiI4PXvGo67gQJ7yRhMOyUAgQt2lOjHdklVR
vRbcOkfdBSPXeFEQQXLl8ZebCz6VdtAHCwWZ4C2Tasc0rVh8hS8NeUaF2e3kIdqp
1zen5ThVaEg53xGIKrSz7VmH10Nq8Mftvqo6F4mxCkss86H2E22hpFin4mVEjCRv
On9XaKcb1gQSeB3+opEVAF/uRRZOFT+yydg9p1w50nUzbzF1e1CYVyj0ujzeBRxg
vdY90NzVZvn/O1ZyLzACIviqjbyrfMvvYAtKsxmFi8wMLp4iPbXGwRagQ3Iy+wBj
VSJAXLOJlnwb7sZLejW+crSWH3MpDWO6XHtdGIFFxKqMa/VhLQKOsfhaqIMUvEJS
llOlYMsihyRordl3Rv1tvNXitkJ2so23ZRiLbtFYBV2UKFv5XBYDV/l9UDcNt3rJ
qljrGY1xEcKNDfID9YjrlCeZvqUwHjiRQkyJ7VLtPE1LFI1StOkRGONC9/sioCCk
I0haMhE+Hht5THkSwH2g22iLfk0bKlNj4QzZfG8bOLYum7LjoDSE3KhChPubN9Ta
DPJG2aWz+tMI3uLYTYO2jK8w3K4+L0WUZjw0AWln8FQtL9OpPSPmO6hyfkw58cB5
8T4ml53+Ue9AmDnEkh8+zPmpJi5LpIQ+SHMNpYeLLJLvTXmOFse4r5AbtM88JsVh
kPC/QFvOMd0d+YumPCDmloBcXUgpi80eI04BJBruOPXgT9MwORLtG51mCdA3N/rQ
DrSarMnkjf2gCNi6aI2MQuffTBnzL+4O2tjdc/5AUzZ4VfMppr7zZANwTGdVr7a/
iubQQoPg+/O8CfUuE+6mrYBjeRxJumNj14x/BpJTBA4VXtBuV978rOi4cQGCM9VO
9SV3MYqlfCYN9EKL9PNt5QKLPHZNaCh51Q3UVjBqTjJ12ew3xDkrARQYunxXXzGl
HGT1F7U4LjWLFdvp18L/9Uc25cQw/f0xUo+wD90BqiWaJDgjGeGGthr47xaPUMUv
UDL8uep67AxRET6PJzdqQ+4Ps1thTQlF/MswMGaX2+KjEOgUUuFlEhNBXbwfiD6R
t1WT0wtX52v7oG5XVV/PuwHVgtPVD3/uwMJILjArVxC7bcuErKJzjUQ+tmxgCOsv
+wQFTSXEUNVnXHO+bfZUvfaDVJn2HaDduIdVf8+x40wePp+LwGW7nBkGRcNGkufl
fpQITQDeU/WBFSN1RO86468CyGTwTpA1QBmOsePavaz3ByMeP2EzIzJX2hdo38Bu
yq9aEE7rizHxfU8Tp0FeaaMxUW9+0fJs2fuO6L8HVsZz30pGpwzRPfZpCPyYhI4T
G8HPFAqZNJn8AWrJsNbMflcljKxmiopSRtQt3juu+XhpH60gdqzZuzO7PlwQtBdi
MqRskIUokvz6Ed3NriQB9Wk6YUFPl9yFRE/q/ARnWpx47YlGUgAoGGo6XXHw+lhf
lGnen55c2OaDAHPn/dxdlsI4xVI1wdftLCCu/nyqMbhWWjSCqDFUW3YftxrQxtFM
WdZ+5ikbkFX2/zLFTgLPoX2J1NcHEOFJth34j91WYEhrxF4GtYTaYRg5IYO0hvyn
p5X+b2ErZbjvq4lk9j4CTCn3qRXvVTCMe5Oi3T3iUSwU4yZvyujyGN2VKEcHOFMF
mQ1wkvSKLPD4eOxidCvNzPtpxLSPM/l9gXRoggFuuBVGACbZ3d9OmHl0Gx30NE8z
guFkIZO5P27vdIU217LGZ3UrUpAejLG84VAra51tbYHE1nkmB0Ou7Ibx/5/e/1Y/
RVUaBe7HMFrVQ7IEwe+4AMfRLu/DStjnVhfQnZbRLRMo8Npx9P6Ky4LCo1vvjuka
jPl/2DXkdWvTcTru2eSjEho8ps44SrQqXOaUf9U6HvXl/sYqzeIz3sBvF3/Z8R1j
RcJMaWmPkZ9Ylce/Lj7cB7tOZ76N8xqO5Ul/1MCokRxyha+Y/ZoLq+eUE7wu0pAA
zXJDUNXbppKWbsIatcbbNxxmLsWPXOAWAZDcCJktrRcMCCIPlf4wET275/nzzB7m
NGAF1ISCZrQYwZruur3AAqpLwcSc3ShxsLZTyD33qWI81kd9EpHy/2T5RBLUjfx1
+4b6FhqGk3nvzlF1AB06i4QoETpegDQPTi1DUGYSKZme2jQpyY8aurBm+cWAkE09
q7pQU+wgPMJSFdwMlYB0rVkc9DhSz/cME1v7IffygzNona3Ck07CFYTywq+z7WI4
Ssf/SHa+EEWSpw2NU7JsEjtuhKHEFG3aD8u/EIbQiVXJgomkd2M5wQJwG82ZRBol
khutUbSuJzZI+uHwo4vrKDQQgWa4kjUpDIFsysExY4+i0g4EviK8v9uujiVjUHZp
t7fhLB9jHB1YAuCcDVduAlXoJ/4ngJMo3wIqtOuMA7zADRm60aD1PYkEeBCPuFxz
hNAEq7an8ZUvnZid7YA0rW6xjJVIBfqk4ON/YAgiQHXtnal4BmSaF6s/yu9hZt4j
Cb23GBKGrrH/gbZerXWAPjALHDgZrmZQ4wNC9o8PaRCX459cvoL6IsxX96MzT2M4
sbqHiMjlddIUav3Mc3wCvu6oO3CIbQWi37F/e3WzDPWxBFe2lpEuE3cEQBfiCrGe
k1MWCJEtBaEAvJV1TIfTrni/VFVmGRj+4EjaRjbBDlgwb5TEvjJgnf18dyaHVjgq
Dg5kB50+8UC3vdj8si3MXbR3RoSNSzBYowBl5PfsTrXhisfjrlqjn+Y62A4VFb5S
vD8F/zwe1fTTbrNnlwEVHxqfGD2R/MxIO7+kQ0U4DxZvctzzKPVTvN2afmwVZ3f8
uQUbpAQevRd3arvVd2JjObHXrU5obKroYJ+ww6ZWwHRBVCj2AC5MsbpdAuSOO3IG
1hzewLZwbr1VSBKC/y5eBBwLc4OgzKGoEgUraO1dUJvSpyHy5H9bvR9Jjlgxw4Mp
HdVqF7vtvPMNpUNIBvGWm5oxvXEoEssKCVtYBMUrv3dyjW/1PxXK/VO927oa6slj
x9velKNOPd5GU5ISQAB5h/9+5YE621EGu31FB2IQuZJngpykmn679yRfLBuLL3jX
4UdFEyKxBYZakEYnLYcD9GdZUKrwFO+LeXVExWn+PcMGSw4KpUTak9/KnULy2j58
bDoreD1rtRYpHoKqbwCuiCaWHv3Eg5VD3O19goyagqJJxjpU+YA+mkXe/63QNUvh
+YXxmMnvXKhxneFD39+yaVfe0RM7FJqOpVdrbEPrhUVc2yQ8iE659g4flSPMBVK3
Ntm6iQT0xnJkhdaI2cCpytUT6ufMwxraQi6HCgmjkuq78K9X+iSpcFbfe7RUy0JI
SgjhOBzydQhT5gxXfi43RJ++5e+X1HHUPcVYhv/lZEAqLyxCdW+R1yL/kONugR+M
7dUUkYjk/VF6fg/kGq7FRSkjYwIllI6h2DMaWcr1M/w4rvBZWAbydd3zl40tt3GN
BrnXXtgEGjtrtmnEvrSToiGlqLRWrc6ceCw+hqGxsSSospqDjlP+D4O5DZcOz7dS
Ul2y2Sl3HnkOAjFWy5wh04b7wYwFEsI9Ea73+hnknFBxiCKkmdlpEJ8yz0+hjWdy
XNrukBqydFI2in+a/+jJfnIqNRpUIp6NIQvLetVnnxmKn3LOjqbxlGiTVoax1NyR
CACLRITG58Ta0JkRERFJUsPpGnHaHs1ANhEegQsB961yHTdOEHfQQnKBH2zoKOq6
h+hYMFugzBsuH6R0RdI3pRuZWB6SGtzmZtSQHUHHG/YWW0la/E9SJ3bdJJwAXFw/
9DTdgfO2LiQHy5CfW1UB/L94X4AdjW2fghVx0gPjm1jVuxxLC+r1zDT/D1owliC2
6mBrNw0CwI3EMoMSsiM5Kj8CO0YNXu5AlZSmimQjvl1ZF+VkumPBb8r79F+zEVNo
sojlsI2aiJAm678Fr2xArhWU/jqUZEY6Qeu+/WxnEvfr8gbA/Iyhj7My12h94EPV
l9aNut1EHfjCe3miGOx9zILefVScVCDwSMGDj8wnZV84pcISS+a/YovOjPEtxAPA
qUDL3CGORD4iQxNliobd50QpOnD6tMbgLCWQvXQnPmQ43/TEimBV7bE/t5/W4xtn
gkvOOgByTlBeWObCm+ss8W4H3h1KIFX7HBuMf8PvWaP3DiPsUFRV5/gHbVnxQ92Q
ItP+IAbXB4jrm0LjSldXjp4QDvpxEKnZSkmuZFwk/hcsmw1oe8k5J98qicXbSRbO
/uBP4oIQoccT2/JPBXqr5hnU/4hQe/jEt9cLlawz29UgVOJtHTe/ub7xTyR99HmT
zqtPqTQY4bYhu3ldFuX/44jTPhTeaHq0XU5reOKoyyOoTZFAn+te0G8MIMkrL5RY
BD/bdJ+c1IE/fMPaEmlzvHnst+uEILJjzCwxO8kxq/qUf36KQ8pHxFB/4o4VeHj4
+IqIK6mjshcTpOtiMiyeQLNd0iBk8aCgHtv6l4Y78iwFBklmaQ8cQ/XPn15XSEEr
Ed4UQKl32ALXjGzc8UD5NhIk89zYxzsoOScS8UUPjeNoaVWtJLM4TKdUMAFdp72T
TUuStyE3RDGGq7J2IbI/b9DWYF8Ak1fbbxVtnBdSOFVpbFJ2GAKni+TtIFFaH/L7
6VUwFudj/celCp146jinTjDUxRjD6qaQe+nvIO5cEgJiLBecmYdv9+g3K9uQmt80
X2BMLitiyiv+4Nuxwh06guEkfYQbZhACMSuALNuHjPRS3QPIwvj9+ivHnqai++AT
x8EJAclvRlflwEkOwT9MXuGrV2Mo2zdBJCvl2xU7VJN8YbdgcuosEQQvDWU5cf/r
Ta+QfIPgcippy6stQPn1TogFL3D+iOtGEzx3sufbgykXdr+pCHn9+qq0qS3o4eNy
c3JibtC3xIysBBjfVclZ6a4B/6t+xt8441LdXIh5Puqm7CGoGz/FuveSNkDfDj/1
KC8uT0txVyJ4hOn8Mu/U+Uu/abOhPGJ4bgBCzHOrH19BmoQkhJ5k2WEYI6iO1oN8
4KdW7EdFJlIo8fFPhPXt6HbI0iMqENRhuu8yC3fDywmsPAmGA6lUqC6vXVK8+5Hj
NxVKc/jwu2MmXP22kbp+/OZLGNYhICzDOUGaRrOq9zAx9MF0SWrLYkaFwMZe9rAU
/nR56eTVRTGNm8v7Ks6vO2vczEcijpxc9jF9Dl5DbKWnD8HW9OX/fT/un/puf34z
n4VSk25ZnMQ/4Mafk1u+JznsAnRlpWGGQqr3RBEoSfucgpIkBcb1poRasH95/4og
2YQJpgvlb63CUCATl4kVz2pbmrKBpdjKgtz2/hnUNxUESfg4OPU9WB5GpAonzT+h
EQrV+39KwhObdWcO1SG4G1fyvKmrEQUFfAvXd30Z42J3CxmXfzNlGsteGRFEMEui
PrdLYKECuiCPbdfNOZSYBPRxFGQpSqYnXQH93G77s7Qgr7OjuEcdkAC41jb4YdkY
+KldJ7+ldKifMPjrHEUWJjwivNmh8/EhGmq3zH8yDNyRzmQzGHCJ3DlV+m08S3ZS
WqY4EM6HKZl4/zWz0QJSCF9PjD7v8dD9uVy8kqYyWvMXCZUFv9znAS+GO9gDmPFW
Fw+QdOE7S2UGh42KHCrLvq0L+IJuhhqEWzz5dofSO7ix+iXFoglY4QfjXvUZELLK
06alPUoPts43p1eRwT7HCLNCTr4EFNbMLyyK9XrgVPtQ9fFn53HJtru6FGt/bEnq
1YVEPB6T3MU9LzOjJbbHKCI+tCxkE5Mcvg0yxnAA5UORuMCqQOdueHznyrj7Z21G
3U6lZvM8fsTHRO2kzTRoP2PKZlbENp5tl7GwuJZ6bVQPHMtmj/XBkHL1pE4ld35X
XjJKe2IQc6yaEjKKpLjDfPfJlA8aQBXH2vtmJyn0ooowyRbg67jY+4c8EgUooh5V
ORAUCI71LudOCc0xmXnrmszHXCRl2aI2SpOom+ALj0giRwTkZBslQBUc/UjqdFkB
LzRKoLgHQ1NjAJFMt6L+iqxZnDRyaU9iYcQhg6fWrM89aEdlk74E2JWgOuNMHKb6
bz8Ew4RMkXehrzOWleZboBR+d5muGzHLn4JhzEDUqAoQnz5oAS56ot+fOUaQT6nK
L/7+CpoTZFrZHpN1coOKDETD8CeU4ow2ziE3Xra2OULSw3hf8eUXaqiHha7AV4Z5
rWxFc4y0XUuM7elqD9kSJ+bhYiz20MvqNvduwKD6g6mfOXI9o/0xRcn5DfHWezxW
Ml5/OW0TzYBW8FT+kHzrlRFpLOFz9tOpGbk6Gwf5mLyw4F+PF2bSxcjqVd5NFdAd
sUtIN0C3/rk7flvNzYVxKXsjWsI3Cjq2LyonSXLtofmqJwk8RfY0XJm9P5fSGEUL
ly+OpFDf5sSXe+tN5bE3mZz/lmwfeM8D1Qo9Q4I8P6fuRjvUCFwvOXIGSrSElrCo
QDpHubQ7218/gQTjj1ig1/AL6M7kCFJGQH/bwV/3lNzuNlHmB5LqOQTaXbfK79tH
4Mn5un8i/fzytsdl4yju+US/c6OdZ1jCDnQJamaQ82dAy3+eHnTeip/kXnoiRFGl
kzszWRCCfeZX6ALPJAFAbM3OhZ7k6nK/PkPK8GjhOyDedM7vO9dVG57jdPTnupz4
2ELctkgEhWkuhdUk1YVzjDeqjJVh2t1UxGufcqt2GjBM7QPwxUhfaOGk+ORWeINd
BtxNJun7vHrgsw3oC165TLG3M168LfXj6ifGA2AEop+0vO/YUN3rWwh/z3AlH2f9
NNyA/vY/YW+I9UXD34Doch1i85wfkrCmftD8kU/tahi0TKsP+3PnF0f8ilhpPylU
cUb/EizU1otQ8iw8x0Jwf0BFvPtghY8ryjtIceY0W9i8HJybthzU2HnW5NHbDuQr
icXSxUROcrcLj3m/oSAV38SyuFmCHKG6OrpTP4lhzo0LuN2agjxKbOBjFM4oVwNG
SdpPPga6O9v5oppvQWNQizX63Gpg22dR/9ZOAk1m/ZQj2TM6ARVob1ZU5CNPDV/t
3YRuNcCtNJWCGGE/EkqLRKbpMtGYAlzcbCYcgfpTPZFLvjjQGplERxF7HhpXFJvB
PlpP9UzErm4hOKsmF23rFcCwG+arvRxwW3zbSfx8LSA1aAwU0pQRHdwNaww5dinA
ZhtmUhaiioGPxFydObC2rOVhjKkSv/eLG4nvwuoWor+dznuDtnSNMpXBWgM4eWsI
Y4vaseVfHTIW+wNP2EU5xA5/pKCAlfl4SezjiBlnR3K2Moz2TOvxBSCVcgMy369P
M1MBp/90hBFFA8Anq/QqQVkeDAJpZEya9r9xrBo+vlIdwF0Llc12Tn8hWLv8uQxB
s90oCt6aOKXT53FNmrV7i5oB+pS8+noIq1yPZjBJrR2Dtr7Eozdi3aER7T+fTxBI
1n3AwBJQxM1+yr/7OmoGAnd1aGoAYCoZKhJ7VcLsqQu6sDgnCXMY1PqfZpNfO3MC
35hQAe7HoIIRMOnkvIGriGmBI3GIARj/e86MePgL8ttlAnE4toC0JgTHuKH+oB2O
JMIHzjicfN2wdzJUnX9La3lxzW2MLZW63WXaLpdCwUW6H2eiIO86EICHKu1MAum5
K/atRlAYZ7Yp7hZy2SteOdEpMe4Vrn7dzVEofI8fA4hHa+fE1QAb7KG+/8sF8Tjd
+FnNzbMcHf5KQNSbHQ/zj3iI4bP8nFSelueaEBXSzeJ4vOnGlGyjX4P7UH2kb/bY
TSQoCHIsVR6/bgCkxPj8he/duhFvMxv32d3/6ahxbLLJ60zmR6mBePeZkILT6ohW
s7+Qx4mcUFqT0WbYn+q/UAXM6Mz6dulHZDGJ/jAhPj/Gri0jdj2yY3GNHNBbI8Ml
kA1ai/IkiDsBsOUE+D+qeD7bFrZVPrXCrH/Oy58Pka/DIKW61wO7GtAiGqNtgUoy
u8Z+6nkElBU8iFi1zisqDCxm2nJcfbQhr6Bej0Lw6gD2rMmx6+BYBsEpmyJIR+PZ
9PeRsFycdN539KOavLk0TC3//RmlxBgzOFEnLOGqoxL9xtBQqSjACn3zi1NyoEEl
s0TF5RlLCMM9BrxhRdwhFoZljNvyjRkKGlvHQlI6rrqwcZCLQ6izz2UrJnDGTKKr
3wH2drCer5JId01wuA9EtDWKvfLoqAoFkaokKrwmLLghgoyAAL8Ld8tCJQ0SJ33t
VIChnGQVKnhignNPeLV/pKSQl5lMgnqrfHxGblcfeMZG7BZNwbtTHqxwrHyS92xN
DoOLyNpYBxrWD1QH20ILI0FDkQrvtP2o0zedIYjGdalO5fuD+WfROSWJG0cgkGQJ
+EBAKRrtJyOwTuO265gLNdKq1IO9T8SJXALZN+f3mrOPnK06VH2Aoa7JNIrKffIM
eSP1x74TP26DkYP1hcg3+K8cRuDVO5AlUO01jb45afGAzZTCk91NV0iDpRL6cNOe
+RQepDfaqE7cASQ74A2g0rBKI4IfosY8+iTuZY3NnnJal4A3SjVvutib26vbg50b
Xbd+iq4e29T3ANXGot7ns76kjOfJwOCpOiZmDmGDMcHQjr9rOeI/zb9zOuZ+K3C6
iSHobvF3hoLAIoJiUhblKhYslZ+Hp92Q7O156Qe3Cqt8aftw43G/MYgk99VGjqLk
H14ewKVwnQdRzZMdPfbPMBNqPqpI/xKCZSv6epc1IHjCLPQIUJs1K8fzYkXlvXjB
rIcErwiIdPFdWK8wUXXavyLdTI78IZOKVa5skUNJkLi+QEeYIKBlW3DMQefHMlvt
2vXw5qAj6+MG0FXFvsOX0hgiBtQGyEgktYOUY7T135X+oEOI3GYvt1UAGecDSgFe
ID2B8QCAJzlNSOF/Myy/MCHBBVDVaD9Yr+gtPewZHJRG30jfWFK0VHcf+RrQGmOY
YrQ3MEuGlv2PNNDa2aTgXdnOdKJl15ELvIXkAyQD8u+nIZtPSfJUrBorhypYOOGs
0dbcv2HxSdrPFtWVqXeInIO2BUdMYkpJ+bh9b07caPqkfmAxrdvCiAuyYPlxAN/y
75RCqNMN8qkHFRoAyTzL+HCINRaY4z3xh7MbNcoToX0sf6Nv5uFVycb6jit1INno
MfRE+INIXaFKAA1LUVI6KVnLRon6O4gWEu/t5ZfUckRgHSXjsjVg/yK8g9RFPath
IEY5EiAb2cYUXW39B3TpVg0so22KHtUESrwqpkJGTmebqw3mPizrF10wZmmePH4y
k5jNp3ZmQvZnsQbHFB68BYBb1lhqK0JK5IgPCrlNRTjBGccwmPV/IUXzW8A4HoxT
NhXhgLm1a1w48lbY1sh92/X/hAMTAIMjEPQtWg9g/WWKw+B7Dyr6g89SOFfI9j9K
HmAg9KxZxSKz+PrUwQ/G+lFu86mfImEEg5ZFl43J+cIJOql1HiqJRjUO6H1ABEyx
FFjgqnR1HQYOPVVgRzBkYAx+euNtqWOeqJ4sEyyMTgFaim1elx3oqe2X6dQSk7E7
JMPL51E26MvbPqXptVmP/CYNZNGIoEAaUUTPoZVJvMDeP6E/XW1HaK6TjjFoLkLl
r2Xbo0/Q4WOMmeudc4+lUshKMIT4lN/+Bp4kbyb7tCAik3JyAoMbgoLPYTZSmVCk
vWjWduZa3ZWow26TchldwrNoN1kB64y3jn/+JjLvgy8j/7Olet1uS3cSfXxi/WJf
hXgri5y+T4JPO/eiR6nmLkeENPwDra9ItVFj7joBlx9ri+p0dj4D1jWEDrw087pz
3rWsFfX8w06I5zZAWWnTysPfKhVH97WNGptyVP+TBu4tAOueQYGfalwPgu+V1OES
qQlcx3iYcewSvAPGL89OT+LailSkSJIc1GcYCZaYkkJ7T8eUdwL3tkJBPMedrLxa
gvXPcP2UcAe6mnw0Tk7fx/me1Qeu1Vjce7NtAsbx5oGtsBSLIUIAJbAHTVY/VO3j
XuaiKZScGzX3msmJHJ5EwaphiHbgqZuwovtl/daAINMOfIlr38nCujkqwOCyJPqg
S6cE8aXQ4O9A/0GzxyrNLB9BppfSkRfY6NS6Ilio3Zjeyr8w+gkCJ090QXTSK7sC
O/WDYIRWj+q/Q9VNDMuB6Jl0Ziq9QxA/1FNR452kIobP1Ms4PXLfT97kUsMcbH15
dlGQIv8HbIPTKWnTAsyc4xclHyz8TVskgJFlJxuHeXGtmYrVjuUVM0XUdiex/WQm
4Qes0fBvtU4WFxwzhiTTCbH/cv1nRD01mAHQAe6khvPzg49bTiD5iLHR+Mk0qGZT
blP6nqxT2XrolYzUCkp7DLvYK5Gj2l23rz8rmgxgt1AhcwPseHpWbU1DrEzYdtyq
mZzIeyJfe2OUZkt7STHlBUNBRlUj7snj0jbn2imLFjWYzD5xlR0OMv52ZDBKXvJ6
mjaY7R8biHE9sfbk8SFCYXFyejCjYA6qIL3YuOzSbRwJeniv77LQPfEA8ZfC4GgO
rj6ix8xKKr3hvi/j9UWionYnu+jT7OrBnJOtmA2+Ht8I+sHOHS9FwQDr7I3EPYkl
nUQBY6c7gj4ctSix2vzW4K4nT1ULY1eIYboac47rH+CGontPGbsItjDpGSLtNZZj
9hawWgd31vd9dAjJSeiGdHkJ7d8MkVMZikkIq/3hbJvUO3n80TiPgyBkbxHbOZfp
KiCjiwdP0B0j52vuy7Sa+oideVRRJa6LGziVh39lT8JMX4E5mCocJTv5IgDkoh8h
Oe0tW24SBKIWlKY4W4yAwzbTNUt6QmeH64207/9Na7T4AyzxbxAoIXla/7N6UaFQ
zkb1OSrJqljNCOOCLaXOuPfkPXlrEyJtQjzTVTQrRDJcSet/oj/Rlr3Oom/bmpok
ughGld0ozuaaMGuwF6+nYg1I29+NT4xM19nh1GqG0w+zc1zphy87+IDjN33ycLih
k93By39dpYwOol6adv5zN5Z4czJUkCvKgCbjzAThg1esQm33zCIibIDB1NCKZzzm
a98u9KUhJ/oQsifyYtchew==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
mieWCq3D9fwjcsp1ImT3gbXsbTbDT4PQ+EDd3YpmCXzYl/kGh7tOsoQqatuZ5Akq
uDl+be8MQBY9cDXGwZmqqGkCxuaqzPtO1kqpFN//E+GajiFaDnoR6OLnjkN28n5g
cCMz4RehVnom6k7bgWrcfVoaXd/szzYlXaf1vic921E9kW07gQ0Sr+yE1W1+bug7
1jwLd2+YhAV3bc9QQB3XX7al7uLjcOP5WeReDJtv5jZUXYImbmWxZOLWSsLGJYiz
k+v8fEUH6Y/AhJQpxKnKBoM1MegfC7PItSt5jEDv6FoCMnznjqufEpQbHOmPtVnS
/MF0TDosPhmQo5CcMWxiVw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8400 )
`pragma protect data_block
KNdY4gw9tOBTxE/7PoDhA5wxZI4oba34iFv0RfJaeIAjB3/wuFvKUrJcqRK+zi6H
quzWu4G/d4n6UJdqi/v9PFERMgCA47/dDQCIGFYpoFC5Id6xpXTyHgCeVFeBt8s8
LK4E8RhHYDfBNOo1lqYApivIMkVbDgNZe9MRkq7i0IPPkpMrNzLT2zgS+Ai8JV9k
7NOKKm0532nDu9JkztbHHx9bLOMA7gHpwq9kr1UWjcRrd3L5tsT/AjRpiT66Updr
96721BleobCkzOGSJfjqUK2VPxyl8HRf6+RXOOgQB/hlkt5S8uSEYAj+MmBMyKBY
BO44cr5DBTiAkl64knQ79GTzkr2C5BjmoVRMtdI/+ATIjGGCz+vHZuU2rXW7kh7H
uaVC2dG8kHbETwNeyqflpzSeKKkqmq31JJbDRWG4dKJ8oqIbRWflWwuE2ztvxbVg
cOjaksOZ4T7yzMfZEWHJH9kpH6NoCfEn3/FZ8ltSEo0CLYws3Im9BN1JbZr3DJVc
75HpMJfXH/LGvWFIvfdfGd1gg5ujOXrQwg9RIgs3MabisjrXW7piaV35daecxFVS
xw9HOInaakpKrm/gIvaGXmsNqC0T3ejd54EFyrtMkvf6BYuWB2mHeavt8glJRkh/
cDxFgKZNvzby3h5QNF+jEjJpM7qWh9U+Y33i5LZBhvt9Ztu6LUZcNcfGiLcZaJGr
Uej1ksqNpBlQE7J1Eq+x9ZR3Qnb+r2/PXHshlkfwunqnPqvN6WFOGzXao/WkPfRR
NcdKH+mtXY8DW/HcBncY13H2zSMZIo6W38cygmrlM60mDCZu23+n4n2pURTLHPCl
g+a0wEX7YwOoAOihC688EjidMCUZSgf1VLB8AtsoRQLh7fDA9WSujNW0IWiCVw6k
r/gRF1n2HuXSKiaSJkyWJdL1w0UtHZ65cxPuYPphm0IAWvm/bMHUglNUHmPfWcFu
Ira3pyal+QxjK53qI2IEq5eywZjpwv5V+eLbiDjQi+hUN43DSnmo08a7Id9xpUss
EbgVw5NrszCJz1r/2XOL0YOxdup1b8JbmiDWJ+iYlnpwnJJn8oD7t5ukgzz1Ka1b
OrdD6DbWfKIkb0XYYUZuRUU/41latOgd7igUq5mHL4os9Yy4+1j35tJyEX/25OA9
LG74s8Q1zyu9aIPFneCecqRRfWbZ+8G2FjFXTIcZEsnRkPFJjUoCoI40dSzgL45v
RCLOCRd1kLZe/wfjSRXgrjvG3swxhCIGW9DVJOgCdvmWMbPydk6TehGugs0H6z40
25xVWWhzwi7aVngg+dBdUJfb1rbKejp9/dkMEaD2CpuhQKwUqRpC9AorehDGuYVo
CVIt9jZNMnBXkqLxYcESneecXnRoYDbuyBDkTDzdcphNY15foI0mOB5ST3u+vbjd
smkKYdWTJP5mLGmrVqy4v44wO8bxJIVKwm2SRRa6qrHqWpw5QjU2KqYRVReqP32c
IwWuvywSA1kObVobYi2d9b3ZiijFLN0B5hPqnE0bda5ZAyqX4Adp54eSLOMiQThZ
RBOAjSkrzW0ERsAeuSiZpF9xI44/ISUgAAQJ2k9nYhBVDsqqBWKymLqJ2QhHoR90
/K8vTVYFDPkPHvUBEoC65tOBSzI9gsXR9o2ywmRYH1aDmxOz6N5fIB2oTPxtDVax
aaRAmrOffqVOLk8IUOiDS7X2dKhYahk8KexbrzW8QvI9vqocVkU7h9IKQdg4oSaz
8XISr8K5Wlw3XY8g74f6D7jbz+mZUqU0z1V7fnFXjDt/p+NVoVlL5p+7JuSHZP+e
rhO+nLBZxiq15Iiy4N5Xlrbapf66Ytg0/v+8/obCqItm/ZWcT41nMVntyznlqih9
R2Gg7GqskGVVlzS0691/NNjCCou7eGdRWGYAn6hEAa+wCDXJSxwcxxdgYcI8hlWY
wznFpT1cBUkncd+w+Sx6rwhiMYRVnPYWnXz9j8TZqh5UP3EHWq12WYXY5ht0zVyA
v/OTmClIxr/2g1VC+uhs/9+EeFba8/mLb+4l1Rg5AoCIO7uMjfK+D5ufJy/Zmun+
AHoNsGcS8VvAasg7xPwo2NR2Ig4TBW0a4s60bgmmpMD7p5No0rqQMWhzlw+2PGwL
t/56jliRE4O+uxLa9rkJQ+dNEKtr1iqTSvLomSLuES8mE286OdrHpZN0+AGqVgZ6
9DI9psN56Vs6T6LqesR0GMZNJM1fPCnY8rkFHdlL84JmSOQuePOxrvN4XU+AVlVr
zcthWal4FqAsev2bvgqRAVjdfcC0/dnRWFVUW/26Hr6ZNkEp9zTdi9Zo6Q4jGZw6
RYV3hQdvQtd27FU5y74cxtupW6O8JfGn+thVdzEEURDiVxqfzpOkcbkaByQT4Nq3
LnGsiNdqnv/XNQdAbkkjhYkQQYsDSoTeTdUiBKXj7h+n0hYJtqN2X2rZHT6bRQOB
pVHcqHzR6f2w4q5HWqjLAhoYVE7RN+xF5Srx3BniwdQvf7VLc0G/8nBl09GezXcN
msaMLGkZsZHvcnkdl02KUprqv+05vCMfB8jCcFMn2AaoDT70JauBo0KWgBLZNvU8
KbHkAvuQerOGsdyoh6MolILtgAE3124smB98m6xKdk0udZYvGy3qf1yrCtC6mllh
pWzSmGb1DXHV70Cn+B4CZ7qVCJ2c6K0z2nTQKxH2rYlvMI0bF/X1MQCYr3VSzZCN
KF8hRC7H5bJl+hTy0UZvw5OdB6Whbrt+iSZ7uvwfmOpOiH/djUMFQrChJR3hhryk
m20Wh5ud5LIT9umQqGp69jP/xLxpwbde6LuXwq6sP8vbXmxSUe5RqzYjgxhmMxXp
bWwsKhFME8j3oXAwtr1vQsBaRaxJ2J15mJ2Bjoc1N/rak7DFwWLsAzZiJDtWcDOn
iKTaRh6wcFMJwPwXPZS/49QhydKkosHVg8RFpeijh14Ee7XqfkSuofnhapVvoAOB
G+GzZrn1Uvw/g2IRE1cmg04MaxOUSee8/JkAUhft4uf0GfDylOnERVkRL69EIz8l
4OTkK7mok3BXh7g4HMOnpodwcomE2RZVWlMqpS0+0onM1xHDBvr1UG+wkjLUcLFX
/TE1G1Fsajqr5Nq89NnAG+MYC+U8+SBdjFoJEVb4Iif/wUTOtgxOAWkTn8a4KMmx
rry0OAfvi5LE4x0hCDZNm5hrQ2UxQGdmZak9NYA7VpT5OAUG1iAyU+qzsqxxWfq7
Q1z859xuXzt+XPHp0yyoqu7s8x4ls8LNq6oLKch/LaXfIDnAnQOVdFxkOB4ZROaX
b7TKWY9Wsul8r02+InByjWnLxg39yK5fssfOhpCfWnsqxjGrUjPLwBp99SYK0A3d
FX9OYTTplcL223L/nn8abmEyW5LCey4XqHabSTKvGG0GZ+80HkWO9sesAV+hvGb6
T6aK5KwqDj9R7mi8iM6Ix1FmnrDEnwOAUG477w6P8hsZPxwO0DurJa7CnFsu2efv
PmQQnnOdj5l6kkg/AhBR/0FARbPfIHNERvPwQMoejDP8GWGnCOGRL4o5RnKxrtnd
EUldZ4o38b1ttADfbSUumrVIx3yGbyRCXRX88VbBicGc829er6VgclJtNjqZYp0x
4K7oBF1tktb10M30oHokU979hE497n3W+gIKFnBoQ9zqr5xShGeatoypMofZwDRb
OHIg0QKlzb5y4f1DFBqnWhb/DMM2d5JWAGVgKfEz8ISxGBkz6q9Syu9ZU63UWrP+
rlwqrfNA79FMxLPuTnZ5O8MIBhQVanFmeZdw8Vp0YLpEi6NZ5e6nWr2o611Es4h/
NRmCeh6rItJR9bvrJ099rQMXmAkYNTypRpG3ZCPM+2RI1tUNpohZdd1TB3R5x+ju
OOj+Wotedw/3hJ/YqR5Fv8M/h/GTQn0ywT0lUApqFxEEH4lrai4lmARaGWv/A7G4
NvSOerdURyyNUPfnmjlYM3tpCvzyKPb/JAD7+v5aE3Dil+RG4bEWmnfSecCWtHIC
mL2yt4n0w1zExSSjUOePyGKQgU8LwfyCc8CnQVnV5GW5PtX0ji7kq6/M941VF03f
rc6qpKkZeEJScZrOzCkrc5tuEhCpTEc1Y3RLIrL128jAvt+hBf93JaaYtTTEtXNr
qYeLcS6Glk/ED0AH4YMH488+4iFfFR706svXHC5Wz1HWCCKaVLMHoZ7yALlWELk8
wEHu9fnUIoqLol8FEb5Dnzef907XNp4LgbKI83gk4afZKUSPY24xZH0nURnxVnYm
b5nLHL+eIuc01AiPtIUkdPYPlJLiYV/XTwI2XT7pm4aGK41h7h9rzyXwoySU3n7d
frbdL+EUlpi9tHMyRj2fh0b4IFI/X/BJbE+A3rsA5vIBCJuzdjnUy1MsX0ePeWuy
SXK/6DxAmPe+Ke1OLN0WNarDpUPoiHJXE6QQw5MNdH7xfOYBq8+PSvNEfthDMLqw
wLpe9Ru5WcSYwEF29JuYy0dnprPRHknwjuitfjBN3v9sr0CxJKns8BGaAlTW8dzE
zeNqAkgwyWK/J1MhcD5dhfoQ9qQfP825I4QG6rh5XLbBOStjan+fN+D3X5mByCB0
i8VYhc/yRTJ4fir0pD8JLxkT0QHjugDcgjX/sKxplPeFymDWSuoXkIvZjkRqGBfV
kUTTfYKvVzkH7Qg0tqP61Ve4Dbds3ris3L0poT1AtnQPSCQLWXFTgI/XJ7e7zTba
PW1Y7A+mIPXdjTluiiA0EXSC/7jh8HCM9o/4Ps/gCPbpoeIZyDDQXHKJDQE7+HEU
b7V/eyeClrV/vIvEwOonVhg7n1a2/ktJt2db08GPBzjzmeQEtu5Ar9GakmbiJaAA
qFLJYtrFnHRapYdpctU6TrJUfEATrAUlWqxa+A5UM/UNobSkw/5BKfISng/y3c55
41UafQt6mC/pEYwh5vVe+jOVu1ng4+wFgcR8bW6Uk0rb4nrob2M+XzljvwCfYX3v
CaWrf/c7Hp0SG5PDHUL740VXP8nd5SNgcM8Fg+2DqdQGiu2naM7v7dU2x7RYr4zu
Bgfoc3v4703uTzOKXxepIBrddIYeWbP36eDU1nAf6bdmhdpE5ePcW7bVhimk/L72
mZrXcTesTwRKeUaqtgjZUxuw6aDxfbcjujg1WvO8mzsaw57DIc+i8aN5S+gpyAwi
7GeoMzqHp+1LrliH+ntf6LHjUyRqktuHrFfuOxPLqJcnDb6FK6EGkb1fk0RV2MaI
yTx3NIPJ6NHeHX3NvuqdtpBkOF1+a+FZzX5lcVcd/zHGAx+pW3bsjFqmS9BXnkr8
cJ6lI2FZ635HuUls9zh6e9YZcr9/tAaI+1YBDo0ymvRLvMAZlCca2V+7E+oJn/s+
h3nux9+THsSXIHWvyY0BJPYzM3QJtqJK5uCJ+K4AyvY8rs//IVe3mdhcdjqVJXgA
qstMF+EI2OsK3ckidzVm3295kT+RWQ+KRDZjQ8SOxJiv366+On72swOQJqU5roKa
kHsL/ZL2y5RiCVch0VZR0l/RkJhp2Lf4vI7z2D7BX9jRP0W6RNTheR8qiiBCUvJO
UKSRBnr8bpOLZvH/jbS8gFU0bGYj1fm6NwyU9py4u3FHeHVM/rtl7s9kVVKCDgvM
XHLs345KqUNT5Afbec9i+2ca8fW3iJPKlj8BxzUWS6sLjReMX4ne/mozK2wVXh3Z
O43VawfQ1QbkbHWcBGtJIXi9OqWqL35PAw8sCGdgerMj+YcRR5qKcLYFFH+Kmv/9
D6pZk1N4Mk2O9M0Qdw8Hbrx5BIUrG6BV4JZfaAl7BnzbJCZvxoEsFa8dKrEM2WXt
foJDXJ6L8vwdBKE6qYw9qpfL9ZTdbdaEcr84sf0ytAUx/OfFhFaKhHg9Fn2MEdnv
dqsCEYPygq4cf4CkIhUFGuNs9g7BHyRe8XZfM0MWzfcecO/pHKOhNi05/17Vf3l/
hdJh1IaTfb/LOf2nCEGTqwWYEinw61vpTdvB+3PQ880PkIf5DvPL56OFZZlzUeMW
G2YwRLNYZ7giNgAkPAHJ8RrteVYuMFtGIPAe4rQ2SU+/w0/xWvJE/XyZ6BXnuRXg
Vd+LN7GvGx80CVq7eqrLz5K62nviuxasSl+7k9X/RJXkzIK+6cEhhwPlxSS/PiQo
DdB48eY9sLVwa+uL8nprXetL/fOy5aZmOfKIn20X85e+QxurUHGRwv4O8gM1IqC/
RCPphcymgaL0MvTQh2rUMGh0v6/YIpDxfBi0VNTrBseV2R6frJvIq9L3qQnYjslR
gZeJhJwmtyeReozTWbQhglGaoLkjVQUTrvwPiQ8EozYNosnzNLfbC7zIeQz5eDFz
dh34xjCf9ALjOMwVfZCGy/IeYsIZ6JPY/vggTeYUp8pzXjJObWfCN+sjeoEU3xKu
UZRuSpF6htmMHWi1s6q0EYc3sgEAfgXhoPe7JKzuYF4o7ApEiiIHlrWqZjcunFW7
YMQwWIIUOBRoMFV7CF9oF2O1pl81J/nNh+g2z6dy0JgvxklC+RVc6VfBBJhFtbpA
rkyI5RGigtLbgfQqK4nbFKK7R4Bm+lt+6BV9EiGP+u0//66ORHEIpcP+bPDUNCm5
Gq10J8rj8Pt3PjXm9f38HWZhfT6vtOL6xg+7coZfmhv9XGGsKVM3UHSHIZyWZsYs
WrG/3t1Wp5MDEKruQNAY2mbHs+tgN0efyChMGNMd0WWNnbURWoNyO1yn3rhVcb76
KXUA4yUHZz3IX16I5lh/lsODludNoM0tfjmX4QCIWyBaRC7jBGPtbnfUEUhd7MKv
vkgXKBjBuTvZ6R67O2GSOr4UDXeveDHaVg/M1TowGEYdtBw/be7CQ8hD4JWOkzgm
Iobwuk9ccTbi824WrJtshDtdHHA2Una6UBOKSVHdGH89gNmKbPBFAvcBqse4VUtw
KDUTOa8Y9LtLLSi6RaqxnH6OqnHNFqqx7Vue8+hUIapqffhe240can6NrbPbpdDc
b56lqVnBoBH50jeionbzPICbuVGRxxqpORPsJYlAlWYBUsgxIHG7BivjhJO1eeCZ
oD+gS3mMYBHCgEkIQsdUo734tYOduCMWJK2kKAVkNC9N+UAJ2/J7W2HinGJ1tzNq
8/Wv28l5z1jES8vYMyXIWX60RgP9NYNpzXJaH8HMLpodhkJukl93GY4/re9Pntpg
7eie7H2Z8AAsYTR4LiJpCAyCV8mrZaFfou2cLpz1lqtCxSUu7yv0ahYH/3WbRmiN
dmtRNW5HAs4SDdWYWTXboG7OYzLpRjAaf7VldoxXhMWHl5i80pfIg6nG2LIY9Smu
lAbyaxkflGIK/6z2D12PIVi+zKnnK/eh7sckEgdO5H5NpIEe3NDsWfpWur1K3VDH
gFG414ahhr6BMlKnlXvCcc0tn9BDv7arR1USwbSXXgBVn8sLwSz9MSYiMEx2augM
Q+bA6mFmu59et9otUnCGcZKEKDjvTgiPLRzKEgNxcUW1+ddHasoShoFvH90ljE7F
38a/FXZNvOh0xmvIJi0pqm6A9yaivJt8pdFoV5Vy/rOxfuM5y3Tj+jja2C9KJRkg
ndXjYhIY7ILwvDo7HNbz3LKlSnFOWAADarYhNza/61mLhUq6pa6yNUUOonaMnyvI
9OPaQLgKV9sRh8D/Hv0vzUsuJEUXO1+i2KBqehr0yrDD5kYvQXi23CRn8SfN+w3Z
95DWdjUD83G3mnBiAvmYTfOOcVjz2PA0HXd3OCHHBMX3NPRYO/YNplZeZTtJ5fCG
hmCEa0KDJw6RgzPE+9nV9BECun0QksdbwKNTOBf9f0vJdsRbAOjRWQSMPCBDIh8b
PQLi+fkyTfgzvGU/9RwzNW78kziKcGbIzEOj8IH0DwZQV5zW1sR4HtByeT/ySdQl
clBb8JFl1nNqRleBKCWH1TcM3Y3FkGtmDiJjrf/PGD2LR+HDO1ACwFn13uwFxo1M
bQGHrR99xr2oGbFEQh+fx2krHLaM5UCUeWAVhDCKfyQfz2SJpB3m/+FOXaA1+PEF
WelcjU8LMHb5Pyv+EugTCiCYO8J3lntxwFCjz1VFJeiEjAA89bySMct8AA7fmtXx
uU/5ijuCfi35tr9Yt7+g9O3eT6N/YDSj1tUMOuMjJ4O0nxR39830SIGsJb9flRrS
o8tSbXsuQvN/HssH9fyTJ5nhpbA0E1Tv+tSVvlrEYuYjMbkow+88KINrhoHfBuyh
QBtQK61cj9uwcIw/oh7OpIoK9wNhZwWfZWuW+iBoahGoL8D67IkNDrCCrV141rCj
olRdId1N5tH02Gt3uRj3HS6sWbzAM25V3CoJNk8tBKj5fmHT93oN2Zs8TnHvWllD
EMrh9a/IUoa2S7ViSfn8TmdFOJr8uZlwMpxa4MbHJS2OwG+SHoH66/OKaPPF9BX5
b9jzYshqinXoUVoSuUKmvfaMKxDLAmpimiCPHdXp7AtxRZxtcl6TnV/gTgufBVRx
/Irx0zpc7K0g1XumyN4QNJAeM75q2bd14zCVfamvdDexbxm3mXYA3qHzv0qqsSW7
Fb8X0T5edHYvi4pPfZoL30IkBkiwLDaWrWyunNPGU+oiEOY49iYClkcrPjr9x0yY
81ZiWlyV92Q527rVkRL52lR4P1dlAEGVva9TwIqZKd6fmay2EEi64BFsJ+bNhZXD
eVTv2e9jbEgz7yB1wztJ35hhAB//aJjQUk3g/8I1ANXU+3aXBt9e1NcGrmObQEjN
OMu8wKSLxipulumPGjxVeLRmuQlDfUpMwdG9Cjl83RzmL9cKM6mcICSbaKwLcTj+
XQtoMqjgcLzyLz0+7DnZmoWDk0GrImXiTaKt/HOinYfino5ZmJ9oy78FtqwxAwNR
dTPz+oR2i6pAz18bot3a4Xo6H2fz4Xf7Bd+hj3dkGc9GHegxjdogNtBdZrO1WvtO
AqvvfexLYA37WW2kRuNIEmKrQWETfEtjVVc+RMFh68Mqn9gxbdV7dWpvmJcok9CL
GG8KWnnnunY9Zki+GFdlfsqzskkgjt4dm98QpeabYB5rCEdSjZI7v6ka1NcpGGUG
PQANyOno6o/bIf3t04PwARwfp2hmn1KBwU0xas4GGkNNeYiAwkWA/8kRaQJ7Vg17
FjMC/9eqlnarAW11z2l5UrE/Q4xUfKbXM4PWFMiAy1p0MBTLyHgqFaI3ADShBo07
lLHUuMCk5wxVduQOZN8GXPQ34fni7l9YX3KKQkQ67kPvG4MeC3tME6q0EPkTRqo9
3iOm56DXtn6iD0Mw7SvcGV5aNWMgYcauY2AHrA/oMl9v10MP0y3BbMBFc1VhqWFp
tX380SiXyjrzs95QqMg6ChL+3yEzwIMLQIht9ZlO7vi8YferKdeneNu4guJ317yO
cLLzoGb3B2Cpgu66mt0CQuzlHtp3uAwrJNFgm692qQIKVUD9VE/MC5KIFPEm2yF4
x6adqYkn0tU5JT/8eBM/tw4nWGmqjsyfYHGatmmlMrsCVDSC/iJWWe88xRXQtnNa
YJ/OFOlIZOrtU6dxRP/TdI00FfJ344cB12SIJbWPaIScYhQzsOcLBCbT9p0hWWPJ
5vMLkSMCYYHwReCPS+zAnEF9nppq3Dt+VoVhh1v4IfMV/ZuSDuxI5Ydb9HMtWa97
PSkgA3f08d0lYgdcXW6NdBva7dwqqmi0v29U1Q4m5mgV1rbvYPbjku3+LuHgHSrh
CZjCeDlreS4E6OBZrrlFtigfVwEZTHqtKQM3UTLGavwKQdJB+Ml7PiXUXTNkc88y
7T/nXCxgUa1ZozLbfK3K22HvtPlieFVnUwYyZmo4Xk1J3EyIw6pACvsYPbM+52Lm
/PWboUi2SxtLzWiW1lmwtQmuBGS42rcyGG9Vf/OKAePKXJPAZIsAGlOaeoxqs2Ar
dd+euaIPbfngm4MRMN06t1CL5RD5fjfhzEPrPA6/R55JGSVCtdfPCUC6zLKyPNMd
OgLuetKgQXjyYv72S7345OelSXi0G8iDyngLVHQtHszQnQ9qORq4GTvDmjd5Zeb3
VAO4fPUIVqSPpZ2SAZh592rAC5LkngvyBLJQtB+52A926egsL27pcND6XqDXROk3
cVRfSbRTjfqREJdrPfTmIN4vzC8EAn8sWEaC8r0HfLB2UN+fAkK8zfbmXXdm68we
o/rdqOB+KMyiFmPwuOhATyj7T7uPAh8abvrrAZpeaHbu825aQohDuwlfMGO4bc8k
eiBpN/EuDDdSUQjtY9+F7A2Qiyh6ieiVa40Q1QMbSf30WYlqBe0ShaXkVT2HH1iD
o6crDYT0EFZBiEnxqhgHeK6R6ALcvV7G4DNg2LUl7zyMq14wUDTLzHV/Zhw6Mkz9
tzJ173pEaBQbLhEsMZsaygw4+8R9G+fNWDzypzEtmijAaVYlaDOM7q4G/2685M+j
OJyIx/n0fBwo1ekGudNQoRcJAyGoCr58mr4xh/aGLkRxzbLGaQlC3mu4OiaM8Sl/
A5AVeNuguOY8Yc5t7Nn4LOdp4T/ldv4DCerp76UorLiaNV+tyl6oNdotF8LRZvRP
rfz++coK02ctcN4VeTXvXxzXzCDCdOqLQ7kVIv2qOvTrH/0jD1TO/pBeIINDMBaj
2gNk0SlKVSQnJRDB1xoIvVUtOZCPzf2qvo/XcJvqt+Xj18JyFSe3yWM1Ygryd0kk
NOkW+8vQUfLqJNMByEUm54XxnpBAq2r6Mj9ugyBpwc2ivanM2fTeKGeMZOjHV+3+
5n6dCvTLlmafNI9lqVrFIkCsoLqtvgZQuVYrJl3wovgIl9eQaSy2FGaCi0Tr+DgU
NbTrAhnlGO3kfA9XW/lB6H5AMMKte5/lp529iHdhr7DijNtgixRg+7Ta9Y90LovK
u4QmzdCo2ZFsPaWYrk1tV+q1r1834YzLVSnESQCaMCzk3+UfOsEkBqCeNt/O3zvd
2JuX3bCZ55ds2gPhtZqPlzQ+bpMFKZIEJNXXkQMfN1EixRXjVMA8uWoW4QBb1QEz
zln5NQgMCQ8XlmnvrfKNub17bOrDRKjFGvR/w6fpH0OOZBlOdne8x2w1zyL6VRpx
7EzNrYBrARDTN1g8s/O+qo4tBbto588NZH1sKKyHz21MZeQaAvBQL/xG9Xv3SNhh
Uy76EHPaFnnxc2h8DTXrT8xW2AxT6pBJSSgMUQ2q06la+Dyf14tyNA/fL5Fb4ek/
QeGPGS7tEOvX8ZwRp7Np2WcVw4E8I3TpqjetXG0AQD4HTEmO+bST3fhqAgqqhNdK
ODObTe+rc7+bN4H0JtCRNDxaE9qQMzqJEThRQESWD3DcbuIHDW/WlaKIFCSYYcRl
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dHR3I1QqLXcoIr0HRL1/4Ri8vJJlgs6/Y/areH3kxjZ4gt8IGd/W8kKPdyHN6s72
PB3XbCyEBaIDZ7G/uMv8+6pkmXq6pdHHc0QaZrxgfQtrRlZoqyID0E56fE6ww5SO
+Pw2L6vXqh3ytz0Afd0MRsLSqhsTRJi7WyjJubJ1JRZxhqMRLPV0rVtCvIAiM6Nm
RC3lnxRwKb3dHCi0SYKs/ArPu4aKxoHBxHUbKh21HYq134GjaoLtRfB4F7Pm4tLy
Z8MPeil4cPcoZb9hBhOKRiw4CsNmvyG2GEqBjKGgpcHQO6X8x3QfbbRDvIrODJJn
Kc47RhYJTx5v9TfjZ7eTcQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9456 )
`pragma protect data_block
KzyvhXJpT9qkd7OJH/IjKYNy1IqDr2in4sxuTS/fj63yOdcWcoAQXkI1DevOtp9y
9LS/JyYN/4jFqjE6b1oXyP1QuKqncuTwnCCAVG/DdhD7cQzrz6zztUdvAK7YuHNW
bx3AqekXjNMVtApW2GYqye/1dzHw81bNFJZc5WppsfT7msQlaBV2lVR1Sf9JvhA+
7qafH3ZZ1OgevJASAwZcKrripj6mTg5jEF4oV3zsTz41etvTY0hyuvazT4QL6RlS
UGQDkKshRUGRpR/EE8TlP5UiNpimQ0kBOaNICp42eqONCtj8UktUeNbHYSkE+UB8
dMoml0N9jJ6GwDtkG55rZxVrn1bSdpjdhNeC5Kcz04yZrwAs82MHtAryn7z4EEi6
buqjf4tGzes4mQO30RM4AfgOAHlyrNB1E/F2J43QTXdMZ640JJQjygwWQPxzjMoW
j8Dv36iBj/7V5ckF9KJsUf8BkxBzfydNVBzZfsAIcllSz6UDv9PSDiXwwD5bU0BY
iDfbqL0hqNYCdUWJjriD5Bl3VInxVFLvOcVcwsEFItgnJmcnsjF9JS9LVfP8ME1c
4/vrjGiOVvtHK+HNZFHos+Uzt8lBHhykhXWVBUstyXVig4uvdUBeypcBpVCFtiy1
jral0ZEuqu7yiTzQodfKzkaNn+AX+btDhTJALAcg33CH69I/0wxY3tlWhfduP05Y
B/IzxNmnJkOf7Wn+Nqku+Jw3ngh+bK7FaRPIzZbLzDT4rxLn01wSTutGLRrCAkrC
MbC7XvCKkoUAY8WqEOU8mVe6eAyfKRfjjA52wrvnj4iNAH4y1pNZ67Ok8Jm18HVM
bGpw9Efp5luoij4zOW+4o3P0VLYgn0Xf+d/48LocZE8lx+nUR/xiscBRJ7r43NEY
uRBFp2auPB2eh0E3ZrjZrAaI24zPtAOsYIGDJ23IwiUjvStS/jAS97gP71d0wzSE
FQgQWRqOdM2PrdmJbT8y1zajAHrtvpAb6TTpTEjzJxm+j3QBMLAy0mN/KzDpXv2g
tBbN9OkIcDDGDLrhxxjl3le5rDOoJEJ3z0rt9Xh5Il+XrMlhtVZseuCS+k3XLDuS
yBBYRSFKCMft+kKuc5u7ymA9k4VEWezTniQDbrEyEloYkudkOegBXTFZHUao3fQz
TMiAQ0RSE004rkXOnWqN6z9u7Oo87d4llfPA3MgG906of6Rw+n5OM011WzmEAINH
540HuwZ1HBVVdWnidgg+RqIKMmtV5luWztbUdM2J9bYo0Nn1g02Tvs8PtrXsE2Vf
gEpYg1U62kOH1uBZCBkEuGiASZDlxW+zpwNYh6IMnWS/wJHGOxf8Lh5Ta6bXYO75
f/1O1r6H/F/nv8SVzwm1pyajiFzmwz1I3ebBdFMGWDF99Hp4YHJHIeage4D3rAe6
KgVV4rRy60Eo4dWVtM4FOoXunCDoRy/cKQMwlEaxt/4cD94H/l2KZlKyRZTes4z/
8E9JHwE1fGvi2fQe4jd0lSJKEc+jhN+BM1Ec2xRm7ETS3T5MymTAaqDZJjU/VmoT
MpigSiu/bO+EFA9tXfgBEwLKruYADH0CSplMgJu+IUrfiisd9vG+Y0gqaxm2F9tD
z8Wunq+tfryr6B0KmrVLpX32CJP1P5tmz/nOy6h3u6GQkvdQFMkXr3FzRriAGwKd
Q/dYp/zqTq1Q1PZM6xKxQcG60lK2jWurKU7P4xy3OWwlEgtpCIpWBnUMa/Fw4Ibr
Me0Hg6u1Dk0oqbkUb1MCjg+n+TVnTkfxVjAbNqY2/qonra4n0tPO9sJpnuLQrd+U
XLyBu3ctJd7PnbWO0wVR305+sBsK16m+cEMw6F9ET4i7ehCJLGTQiWYkVLCgnnIB
ZOKc8dBI7sETrxxLlMtPGtpa61ecPYYPiD4i9sBWNuMiQYOL2dRrkaByB1KZZiWc
YVG+qmEfC4qis0XLs/pj/RgpQF0vrE5fsZBk7FTQ2o6/ERPa+I+APd3jTTEYV7y0
zhnCq3/SMxiQAvA2sGL7jiAXQ6mits09k3OnQVO4Qu8/U8epfZd0WBoespwy8Dg8
vRqr6V34AAHm83kC+KIhY8jyg3Mcca6wiis/sELGhwWeb/JMQ9e0rKbiz4qwNoid
Pj/fUZdAJtHhpiwXKSQ0esdxxBY08R3uSmUVVLHhuhRfquAPKdP8/Zq7mQE5LVdX
fKT05IPQ5fMUWevsA9dcUWdpGhg3OdQTmVT9VbAMUDhLEQs7Ojc3v66v67q96anC
nmv9+9ApTXExyfmqijdeJyJhMwFv9N37LillzSA1f2EM/8AcEc59R1MDP91gNI68
xhsMW/pI7/u6cE9u5DvKSZ8Ztypz20gcWG9EXQx7NWmt2PHNE1OXstm9hzAEHiIQ
DfWM1hl5e+72NxoDztbg/lzCQx2aJHAnKj3tBqNigX/DfKJ3ymQ2mR7IJgfRi+gl
r6w7V5Gg60sJcCLYCUkbr6t5gcVECQ/C2Sy+Q+IN+Kymv+1UubhYehjEuqNL5gtj
Dnm2ISdEstP80xo2j/fav/TA55zopJcH3cDrN4zSAVAMnmpDYipQ3ljJPJT6uo8u
QI/hFa1usiHv8Q4w+RlOjNpDk1o8jMQMGafuCdd7e5cgSV4w0bTZeaH2utr4exjY
X9mgkEZSBH+Gi2Gb2lRUuRJnSgE/xhI43T7zTV1qbwX1kjJLmsZpKt2LnAJ0aNJC
w8hKDrb5hpxI9fKBHZ6mlKi3Hzo+EDDNyAE6WTrWW68JfZf6spFPFOKW7Bms6xSI
nzcUJL32tO7c9PNGI7Lz4SULtKQ675bHX4xoZ5w2s7HO3BG5S6PTdd4S3We/kwEI
jjixtcjq+EdM7HgbPd35PAH8oU6cOOx7T/j4RhgwvQtmwDHOtOWwW5k3mErtYmir
6GGhj2zXzsC6aEpOrZ01R+mrQ64JgQ+9AXM1D3Nl/S1GMj9TOdusvWeEO1sRlVjn
OXprJi9yoVTWsY/D7fBqz55SSUid218h/mmNjWnwoEvB3zESjZHq29JeysMpmIc4
itbE85QuFFcJrQnuoyi/Bq15/gqQ10F2KPNhrnQoXsPy2LBJhKIKALvm9qLsIIK3
TeyYnplPlKezrvZM4R6dizzDbD7w5N9s+Ttoie3WRIfhhrwJI7smdzjaDZBHTvyB
ULkaAtKch/MhcR9r+4ogX2nRNIDwXg5j7V4wxE5DmKqU6nkl3DDbva36abzRCzod
k3l/SeYuUKrbZEW14f/KR2qFqQX+S4TryntXKaMbJ0XEgdLifYD4ZOnd2j4+mU4v
fuYOCoZ8UzdM89d8xL01AkHCuhgWcoNiu7EgXkToGLxdJw3lWaUWkkVdAl22mj4S
eY8V4tM/OM/9jOFgSlN2R4agHsss+2hwmDhelcqJ5RUWd0JRy9E2jUecpjnD+y/A
viRLP8HFYlfjpgnRnq2YLvrVZEXnaQtFtsYhsU1lg09x1hDnrXeWISRL8x4AP+s8
XLTQmxCVXZedPfbQASNX+ydgHwj5jTR7oofBRyUjn+pYv6QwIbvdIehsbLcEdaEM
CKBrBjjhGGjWeqIQE01Gm9CC3/rMVluPXL+zkS0LZGK1HzGuJfgsf5XEjGquXKS/
hei6sw9uICMo/tGEdz+/BUHZfPEaPwwiVrgqEfILfbb0SwaKAo55WKc+KkYWyTlh
pgDPj8UrTyTvMQz8RzDC43E08GaqJExwd5kTR/pE76DSSUt8tnF2iTwBO6Lxi7x+
ZbrNGjlMnwaPk57FfUugl6TsTFx2P7X4/2QEJcEfRYj71bsP3JM8O5kpHQAyJi2b
KzwoYe2dPFUoO9HVT8GYn630QOwxcmmD4QIWabqezRMfZoCJGYhsa0yP9D/JsGpj
GPiEX78mOKnNljcwHqLEsoqEb3nhowxJ5pZGh2KC8Vl7YKelUWqaqJ1I1ysBwQv+
+kMV+xBws0VKqoJu7R6C0wFu+9UYN2Jve1LTyAY+xkWCTK412GwUh6SjSbOajOTX
0mu7et+Es2q/IGoIvWyaPPtFf24AY8tiGhe6t/6xhIcONvr2rMpyqZ4Fv/BMQwym
PKekfrnyLSjaFlfCqRZL9aloktLUrcC+zK5pqd8ghDF1bGbOLa1xLHsCEyeRqdlv
KV/tlh5Vh0DWxX/OjEeQTyWmDfWuvLBPNun2tAxy9CK7r2SrEFpV77SRWY1dt5Zi
+p+hSyaGlTaPv3cfFP0XthX2gCZrwBQzK4NAVhDOwtBP192RVJLiCLpZNENN1qSv
oJdv1CgmNmzHb1cVD85xi96LbQF9PfisPTMHAk3XWmZ/y9CtyDu+S51FGpL13G6u
kEuFMwY6cHT5rSt4KKwixkQm+49rogCmEXaadVc5txCCk77uDhL7hnB3zKg0W5GJ
wFWTT4Gwwi3uRWoVkRr+dPhSIkC2SOCxJjflhQvfmgr8bxk8GIZRF/P2W3R1useV
yb80FLvmZ4VTbOfDjXgq8AXapuB15tED6Bhss9wyl8dTLb61twK9NbB7ERv7E0Pw
6yktcFAhRn6YFOeGZMIMWmO3hL+SQRWQUFf95x0KEvmBHfoJJRdiSs3qEffH5vog
5gepOLN16qMqQT+ZGXU3lUXreC6ts4rTMbO3PbMVX2A14ThwoRxk/Wryc3okMvRD
4hybtduo9AMh851IIqXNVukpZ9jZwSBRwhKFjUhve2llEpQu1pYTqVkm1pL8eX4W
s3KjabwYI86sfVo6iM1oqLic9IQbdDWgtOw7LJIQld/0c1q3+s4Zi9aEMUxb35yV
qh3MnvKkDjDdGE0mMYS3b4xuE1E7G9clBDg9u1rpHZ8VJcNJOE9eE9QG7q3evRZY
PvLdZlxJXnT+x/d/ARFe+wxydEI4WbqoPd0bvamJb66+cglWV/pC8agPvBe5lxc9
ZK3TWWPQUu+23Pp1tFP0PTH5kRbvaapL9BRnI1cymOd8CVD6AfyrZsduIgdgeyhi
naEa9kwkcSfcfmGmDQZr+2IpQq5rxVj68WJCO3eAFB73hL9zs5taO472GxdVCHL5
kYVgZGmbKeSJIqzU4PsQMhftZz8bwHrv1UpIIrGqUsabBMAMmYHLiqfzPjt4b0U4
K/mJDLa+MrUJJZBsLAuu9mIlO5z6DlsZYJMPOwyu3724SKvqdkjRNKY2ToN+e+6M
Uqg1H0FeOGIYv0zNAVmZcdinYRVmJLXTG6L+zKVjfDzVr8N5tdyXI8QXVZea0CbY
QKm7/PVhVoQKJ6j+5GzyS5N+DfxOyxZVETcs/DWwXBaFOIPdYLTfISSNxPpJxk+T
04MFbsRsl5+KEhVm7ouqNXByVhkNktjkCqoLMqmDMIZNRZd7IjbnvkHleCMltvDR
W+4QtQUpb/4A4wU71WweE6fuztdvrnqeqi9sibK11zLjCIx9FPBtRKKavc+o6SSE
SIIuB26eHflMjl9vH0fTnf5nw89gWAQsh3l2FTkT2Y07FanyQFKNLli9GTqqNn9u
smbckpVHZaVKJEh1kYLfIG5xWb1qOOvD4DyQL3IM+nX7iurLye7eyOvm1tVVmsbR
LrNhHYNa6HIH0buBLahzZVdVnipj9pPdvLG1UsXsHKv6Vb78Y2yYWfwkKy0WfrTr
e2ib8rmihNStY3D4ApeZPpobzfwQCTtwpJzuYFRpx/3LZJ5iGNTlrrAQmJNud9SW
kXwt9rvFnli/HEdJIcFj73obRNC+2PTCVOoiRUO+HhamfP7iJsL8WEl4XeOTkMqW
Hto+9Go5NY12fmKZl9WxfB4VZlhdOJO2ZabK3XDrhIYAB/lvkA8uKYoIDVFgZWb8
drGhm+qZ56Rds0JzihcgEF2jiIYftwHBHuvHV+wmmnDQFqVxOxg/yHZtWQ73D5ob
zm8rWH9DwBg3225zwYmixpF+uYssXJx4Rhr2WM/v+j+TEozZnEqtuf7iXA/ywZ6L
2N7Y4i2KHjy9uiq9QpyCuW1Fss/MSqjiGfd1kAa8n/tDMf/KKYzmkLTVsbpQb0tO
VXhbZh8QAQmIYdW6r+C7MjzHwZzU3EjaR4GiNU43h4h6i/O8yGKSaDE7oowPIAb8
CFIRCcdQ+F/palBvnWo6v0gCbdgkDsgV9hMzSmYdkHZ65RfnadP8NMlETvQjQ256
fHAS1JSoohbQAplpMULi5oc/h4qbXJRuWoOkcMApRUh7FFcqOfllPPGZL/RtVvvJ
OZ+5kapFGr1LANIMZmcIh4QD5ij6cOt2YCBfyi5vd4FihyVP2JGV+qdgVR1STZup
2t56ttsbFtzhBzcvNaw3nBnB5bjgVqSZe2XIUHKm8rwf7CTzmP/CVZ4jvZstZMGC
9kGPcYvxPZlcvMGPFv7P4/DM3MpU3PCQYO/z3Yx12KNwIUr9c8Bf1BtqZbA1p4Jj
eYL2KIajqB7zfDBunMKB8bdNzy6ufk2FBwsr1CAIiyjIFjNvNS6tetdxKyD8TvjS
SISrfdW6Agvv8OnxvXoB+JBlPVXkZr0VLnjvN1qLHQlHKKYX7kGxMsr0aEZocEsb
3VoOwtihYRpcOdFrvnNOOK4n14i292g0dyWfErToWL3mkHBY3u+bYQPc/apUixwR
xA2LnLv7zVtN9miD/Kz7PtdeDPnf3vOD4FYsC5PHxBF85tiY+RryC/P47f1c77qU
CtATM9nUZAay3f3tqhqSR/P0qiMn1rrzWxISXW6NFCtHlRjsQUhl3MVhyhPGOygn
R7HlGPew9KRCJTTnuHjB7sjFO1KTJn3UkI0txwwWxR+d57fWtANeShPXuiwesbiF
RjSc8EA2ZoHXeZtV8jPTu3RdWbn5AYBOCm8TOs76Gl2rJ2LIykDEqHlSPDdyQvLw
zDKTnRJELteSs0Z4EizJcyQPOtCa0UMc97cVhjLCIFOXIYR83zLwjkvQzf1GYhCt
5u/IYSuPog4igHx0GaeO+dwAnAvLoKk2MCn/9ZiRX5m3TX4NJWdVoZ6O8Os2WD13
7KY9ZwAp0XlRX+amPIQt/658AECqHtRtxZ1Rut5xq2lTDBqHEr1XxNLHy9iW8YOa
z4+pg6AoPWRZizCJexxUqb18SdNMpzeov7ZaTX1p8vmeHmnEEaHXSOX2W/ov9V/B
uPH+9crRYON33Zk6Nw1MIzKL/mIHVspqfq23nkAcdvDTx9KuTZx9Q6a5IEnfHGVN
g6bBxX4FlXE5WLUykUn0XUQXagznms/OMa5FboQdgtD/kOPuCSDRrMm2F+eiZ9LH
D+wnuxXrF//8Ys4cGvoFBPUkTvXFaTPC+0tbX9WI78apQVnIf3mF2Bv6bW6mevbu
Ti38eeUxb0BhjaGX8D8hmvpILoC9pXuFcFsz5tpDaObJhvboH0G4nYtqzpDaGVwg
fyjU6zyNZq5XzguT00KSZFQnNwi90lafrd9nAUVD+OrbqjV1s7XE6M9jtlW9L3nc
eOoP43I74BF79LOTzQwevbzeOeWzcGf1Jrl8K3x6jo0tnpOefdnVHvexpKBstxZ0
CCoNonif9zbOVuaRbJHpqOFAKooRxMHdP2B4d7mLZNL+rWAiG3REW6hMKKX6PSoK
IaB2c0AJhZo0MntSIC1mtK6i6AVnGTGnXwMYSSuW2vbeVC1ZdxVOop6dddGfwwm0
W22K3iUYjEEB1SlNZhuRxH50EvjN0nw98v65ItXa9Xl/0Er1zAOyKduNv/f664GG
tHXOQJsj0C5c8K36OrHgHhxITzrXJOXkkHYXKv/jJExmeqVDkcFxcJ97m/8cjPyC
rUSNXKDBLQioEgi3tNPgmgEMvhDLzzRUCIEhg6eY3U8IT5/ud/xQOjAaOgLXb2HO
6DYUjhsFG+AeRGrvZmzXP7HfVFJuhSaJTvldAvkSTOSlCt085fgFDVl3eEP67eyi
J0bBFIeVabfo12Hb0FLRjWT1NeNXhzZCX02D2aCwhBnQ7Lf5N5fGllVYlEyD6E64
FFx7tjjEbDo9hPOkb9YRNZR6RLnhz4mt07SXFC+hmOIsXqMGnYOvsB+4r1gZ5bR/
YWltYnhHrIPJJN2fRtTpMZjZgAdC3cA8L4AIa/1iWWjQOHzPDt1o9c2BStpvC35X
KJl0/1q2yzKM4POuYWpV5IN9sCJB2DW0WTK5xBIeokYyzPdGChWKzBW+LcfMj/i7
ppA2+XeUcX7Z4c6FB6TESFuQ/7UIP1fFsS2mTtIJUlAD1O0AlF7fGNdbFZMhb1Wc
cP6SF3kx7MktFLMJ8rBvJ1Uu1zCkgr3iUrXzP5j3vgdedMrwZFNXJaQ0nwC+RuqH
/Incnp/noaJ5LR/nT6kPXae9FOZ8lFNrf8y8yuW3XT8gnaJrXsotulLeFMbhQe+u
8+KxdshujHBru2MoVhG5GdIK5Wr6uZ1Iv0ZtkVqTAZGIAdCjh8R+aqCdsFJgA7Pe
FJ/Gx34WhemWAjV4z0IA8tafPcZrvHCT4/v37JPT+66m7vB4Xn6adsE/AGy+VKHB
+2wTjQZPKpyNG/rfZQZx6Foo8lE3K6BHTqPjdw2h7Gkju2By6YUqIc1G+YHbzENv
6M0dG9D15Rczcf4NRkk58NHpTYiFy9PlhJwfczxje5MZJcthhPoidvJurW6xC6aD
AQCtert0tGuMdmiND3NN4MAuRfaT9LaKttu3sjZ+ufIpwjSAMkZL3PQb/xQc1T6c
F5qUqB0VZalOwXc+U1RasUtUh+ElQ3m7gFoi5q1B8IS/rNrfMu4y8vWFL15zPnpT
xWj8rvFtI0K0B3Ua+5HLrrs+2qJ9bQVcaYsVSpRbzjNZu0nWihGrhqjPDQZf9bZ3
eivYCq9gq/W2+ft/HNlxzoNv1ydRKnuYB/LFOo379VY2EvgKXFvcTxOPoUWMeOUM
/4hUQ6NrsJqzOKMSpEipSg4fJAAP30as0u7DpjPr4CxuHbqesguYboc0cTJJSBKu
GQBuWt3Cx2WLmZfxLDL1HiHWD6BnG8exeiMFHqdbvI+xb7OgNKRK4UEKdYXXF6KZ
rSnKAaoiQytgn/akovvHsGhjdFViNBN7papWMToi33cfCwzLWa5QcwPhsR8o4DHY
5I3FFXKn0fG7fpVLVJg+zRbeDMl2Ff7OqmO7+QIPVAP72OO2J2J48/4o3rB+v+MA
bv4PuSiI47okxZevvyCxBM7dFTPA778Iy5c2R/a30gha8is8t/QR9+Pv+f5ouOB/
0GVko/lz+nfhDZ1sL+AOJbV4lpIyYrdbrgPcEGjBvDmuuLx4Sa+2S0A0i+oLB31H
yvloUqB5G5haqnKgaGbTjdaKHXOdeMGc2YO0p4HSP1HUzOJBoT0umVBPeN+VYGgD
k/0+0PN02WiIZ20+Tidv7ca89ADvqDRoN0QWk+HLhNLQsZaXNGo/1rKDAHiz7I68
n8tcj17dGStI92ZBXyw5icNEs+fkVMyGmDhM46fEOXVe3i3yYHODZXGyWhZz1zo2
h5i2TYaUb84Y63IwnMT1IkGJBm734MVabOeFyOJ3xDhXO+HN9m4sOMW2s8KWEDMj
wrn1DGEQ2b/rDh6+NTv7e3tqtqnxyIT43C1UoUTbSakk3BDyoQdHC8lyfGhuLfAK
NoBCSjENaxkSX5A0zn3g4iOH2q26NxG7TMwTJJERYzUE3yqrkhsl5G8u1C+0CVVt
qtRcvR7VJ7Twy24tbKaPiZScfOX3XCnkuZVUPxEii0XgsQbilSC9D6yS6Jo+8UIG
T2GiRckcPy9buqiVUQA7h1T2jzMLvBctNfD6mGAiDqkwaLZla7heVPv+CTscE5Qs
vkqdggVK/z2qJtIKdY/V/y2O5q0edoz1Bq5kirAoJ33T6sboL+bVRo4P8Rik4FaE
zETo4HYNBDg6YIBS5kDRamtGmiayBMGVWi+VTJr+QeD99aGQkwa8nrSAjUTFiOlI
kDGvDYC3cTDQETIDmIpq2EGtZh0GyxsLrpza55L0SSrWrT4Iqp/+9sQwCTQIqF7U
p3pxecpLQY2HAOQi2Dq/n6gX3SSn56s7Y86eR05cJ33znXCtFTHfr+8lciKYPn7z
bm2JT15qN1K/mcDKoRG7ZtnTZC+y3wYt9YvHZ69gOavisCdRzLpGB6qa+f84pZLl
6+TdWrSxT39zoF1/ZxPi8Fvs1aNuW7BQyy5cgWj6G4wXrcLeeMm/QkXxRe5VxIxU
hfdm1YSf5X2x2hjIhCQEyUPSaDX1Ia5K9fb7JfDzNrIRqRp1b4GA7K+WTlNQJaJ8
4quKbeJYoSUzJ3jROOetQn1h07r+wMdnYOohW5rgxdyA30a8VokuQ25S03fm002t
R7/fOZgicxHCYGhwmzfNZ1cWv5CQhCPTV7QtW7wskFbgzsN4WAg2TMiI/I8FGEgy
vd071xMG5Y08BO8zC3T3mBkEfs+C4Npe8RVNz/whPcw327NZtYZ2UEGexO0I6Qos
RV8JX2q6Kq76ChDghhS1E76/dPRDfN0s5ZOyLYV+UlrfnoBvh2S1NTWbdb//VnRD
uj5xEriyitH71lMJvUF+wjeKabiU/e0MN953irwSwWzNKSwnI76xLKOxnfArKFXb
rS+6Fg/t07dr3E4yF+q6QINZn9Q0MGppw7oaRqGABMnMx8RZ3Z3XmYbzwJLWl7ak
Ih6xaIilr3iJQ4rBmr/GuJv4QbL0UjdDBZnTZQHXO1TP91WJfE0nWVaOaWSDsOFj
yOaEvjtk1wdBx23h0KsD7Rn4FKTU8UuiW6dKQRu7xukY9qwY1eKrMILPZforKO/X
cAMFjlwm0r9ybpqwVMBWjC5dTTiqfJhoS6pWdgBcsvuJ9SpGZ2db1LkhlhO3UXFM
yMHvAooV5aLMC9N9SKJojH9M/FG3x6z3PDEZ30t/CVYjNwcGm9SjMUrg5hzjxjYM
pv5erpZTy5BXhBEtAVHU3hM3PSo0SXwa1UPcKJB9hFYatyFTzVqrBsTv9kA5WaHn
8aILAVNhYe7hsMtGBRClBEZ4fR7QgdZLG8OOAT5US+bwk+MgVZ+BwXEnK4KaS9Rj
KOlUwljgMUzBkih1v+6XLibBO1LN8QHhZGBu4E26JHZUix/ia7hBc8iwti23v9S/
/lIsLES4kHgPWzBDGcJ8pN0Ph5JU9f2uZrLbVgkLfM8tYnXdhvb+p7Xgvk6IiFpq
9VsxFXRUAdQjYMPgiSTukQKCXL1bIngie0Csi6aQfiB91gxsDKGEU9LfNS/2vqQv
VMrRQNeJVKElGmdk8bnQGWzGlxOBM7oznF4IHwt8Sqe7GvdryNJRDwWB9Q+RtWmm
Ae40RUOZ+3xpdz0C5HFIqXXQ+P3n9OcRHBgLFt8+lktaW/W48cRonicROmhdXif3
HwLDjNtmNZSWwfs/9urq6jAqsww2AN6b+geI/6iFkyYZeX+qNATAbXRgBi1YxJ0u
qFombhhvJ2EzUCs8SJH0PIsxmvzHgmbWYhIMAyLfYl5xoJoMEM5DljaVSbNjk7a7
/eQjTLHyldbET6lMfSgh19AsKu9ml3Zn5rLFgx8zK7VOUc5ebMyvc1PPfer9lD7r
HhF9UK0svMmaJSbme0bTBUoAuz4B/IPVcEO0xx58bkOgr8Z/btIYznaiaq4M1Gpl
qhfsGbOU/5ea7SvFc7GX5pG6drTnNVFDnUhKyeJ3V1xMOY/4tidH05pmfihMR/Zv
/UfkO/8VPoe6yxgX5lfXqPWuCp5t/AEOTjZsjhFadoibu1tu+jSBfQ2RqV419m2J
/KJOrYRraP6827ETvIp76Iz+vj6d3fc7V5U6MluQ8g7F3J9uTqoG+kYeVmJKtSRA
DBNk1TvVOiBFlw7JPBpI9iuAanQ2waTiknVZHAS4J2KQ46aHwIbB+Y798d8YspTI
Rt2cH4eIsyIs2Luqq9iSNYaDDRD3BTeoHG1TVaFlvyhmY+z7Lp4iq1qbUHxZ+HGe
uh7ptqGTxUAdbfNYm2kFVL2kaXTuLReH26DPYFm4DUbzglZ7qcZ5y8BFSX8zIkVk
2jLpwnJaXNvHel1/UpNvWWcwXEE8dUJLYcbdGq+ubAkPgVIvSJkq+/4RdXRqXxRl
qhja3Wqos9kdD4umG/0gjiSIcWzMkMGVM4HGQ6t7JGrI3yct02uuUndJqCfAnOE5
33H1HPUZHlaUrepaTTUmvjBX6XnvUWMBjLvaXfZrpThzVoUHL4lAKqvZ+HvdIc9+
fzD7zoG0e0v20qxvlgbA82ZK7HuPCI3Z1u7WQYgTut4CH8aG2ofxb+rWDWlqxx6N
dRrLoQGXUk6wWVGvOHO4bV9GKslBDtaPz4Bqr92xo9dHBYUmjtIvmAUX26BwvlRn
DYO9CVtwHnUlw2MWH8IjaiEIekVnqQHxdKDHrQXZTF98EA3md5dGbe5JpQOf8Cmm
Vzqw+4HuaMi/ccK1ATM/NTffx1Lxu7LEy+KH/xOydA/tt/kJ5ucOUhs4biQbO5kT
qBL7QYtXKQf7AKCS5GxQeNQyunZkcA7MV6DE3teJAa+cNLSdLAO071O3OgeIZzf6
LEg8wIES7psFzKqUStXg96iT+dlRsfHN1gu0GcF5LGMvtsBVfKFiq5WR5mh91DWP
7C1pZ7lTkNiiLI7GBt0NZtgzO5HTZ5QxyAMgQH1NKWXozc5AaZlCO9PP8kJ2Nh+O
9dYtXFrP2rBGVOF/HeD9AmVTyExq5RXeMHV3HQUF7A4/O3hVRREj2PvSUi9kTEcs
EeA+/NNjGp0XOlX7t9jTH40jCgnwvYq9Kj/09i0qOuRpfarq7S+aYUpDVruQTzsY
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
mhUWCfXVUzYdjOIwwGTRAB1+XjGKNK5EhNXevqED26VXJdpOEHysbezsR3pLnT91
OxJnfvT0T8oqim9UTIUdtHRHo7Q+bHRVqeLfgnjCdRFglpITC9s3XpLRgxoa9++K
AdNWsdTgxmotPmi6SIN2Gn/elAoQir7H29ukSxGSPSO9rh99kImGtOVmqeDTN1bp
84wMX9Mu0mSqUt1ydxFzCIZBFQvgpBouXbjhEsGVeO1SFWbCLJBkwqWAH/pZjO9P
8TiCMUd63wJB3wg345CpUcg0hPpTAVz5GXDPLzByTR/gTfU8D+atJj86Vbln161O
DOGmOO8zLLWQOg9alI40mA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
sz6EKsJjYUVnDkXxqtPjY6xjUyI/1nHAVLzzuxMYnt8ta64QnfeM3bubXiRiCqU6
QOjab37HFi1BbbvC2IBuYFCIz1tkUts66ZaSFXTc+u7oO6XmnM/BQ2VySrQ1Ig+/
QsaXud9xj00X4jjVQXMk0gmSD3QuTHbaZcts9E4LNpSld9ZelGC2vtoPCgMQTbbT
0tC7Byjp66Nqs7BbX8ZCoTBkbE6B35jIdRElgM9MkkcEnwqIj7KDu75FD6sgdqpH
lWxZph9+ycJHQNiYmcselIoHdj/bPGw83ZOaDGW+W4fdZLoSSUOo3DV/8bzEUllM
AerdsL2DMqpq8WGYexFgW/ycZ0JuMaFAvJeG44AcOf7xw360bP4Y1gmudvD7xc0U
JS/5F17+im/SjJgAGWQc2ATJnJLf4kYivY+0vZAxUQOgY0IBFKBerk4s9vbCGHWh
KriWZfqWAD1+F3dr3Ko+by7hJdXyzWwslsrwE26SIXZbafNOCXvgag/ZAXMkdvGc
b1TL9w0XYCXjcdPFe+DCHkkjOd8PxPMhna1lqAKBP4514acDisPeBlcdOC7msPnL
oas6Ugg8g3nBrkPG4CyCov4q/Gf/J2FoNbRM6YROeS9t/r2/Yxk3NVaIroBd+M1N
wNooJq+nyRR75lo2PVuOYzTxlLVp/c4N/cwNrUnZgnCfTwXt6G1GM2KjTFjCXoXd
gXCWInX427tkXlZLyFN/R2t1be0aJqzJCB4GT/5YtZFMfi1qhDW4CDhgeghQx60/
h+4+h8dQfNRd2GGJjWVqh2pODDKh1p6ezyoInqVKX6SsC5MQ+3TECVTgyvPkdvAe
wYSpQUN5UJmGvvtC0vXhb9zyLOiKSHiDY2MTVygxG1gOmHafH2fQ7Lz8mtRDv5C5
vnDuwY0F8VeMOOsYEXgIb2LpWrA24vL7D/r2IK1QWXLNl7i9yq+YZi8UiW6+gM1O
W6sCv0xgMkDJxuXSbTD46yogH5OiCCkcaBTpUzoWcI5PEmUeBVjp8nhwg8pG+v77
JJm2QWj2x82PqG3A2rqDmmnJZ9a8F4m+QYtpFk+en0/Xp2Wc//2sEpbjx6/2Ch3f
POkyEigfo7/P1B28O17Meu9gl1ZGN0hC5/snyyOhL/IOWajAjiRis3uqR/Afbkne
MKiiEeZDTa9kDrHronAMW6b5nk7CVSt2tmBX3W0RX0icQyIRjhQjEAMz7Wx+xN1I
3C6/L1MBAntzJFOJAgjdsUAEZ67zLDcSpKzUh5TsLuZSdpoRNWX5d6Z2lYwRU/oG
k1d1bD5QgxlxkzISlN0nP2BkFOOP/8VokjTjc2epadO3kUM0HSHK75cnNuc0DmYL
Zzz/NTW7tsSZzb0/V/2f9nab7wYKapduPb7kInnsk0Ffp0lXRdPJleVlRhkyw1Gq
MlAfnQTTtOR8qghF1Sw95BTddsBmZzm6Q/r4nybyeQ84a0flM2VXWoMT00wYBpa3
U//NmcNL+5k+th0V8VFuuj7K4NpC2eS9TGQ+MCvy9RoE1ewx63nRophkvKJo6aGC
GoNfIYD653znEQONtfTAc9ePRn4JEh+jD9rjh9/IkCg05AoISjmTIX5uCCQ0q5o+
8syhFVudRKsPMtsxZy5qF8WjY9/zhIFP/kkfVYOmJY78rNBA4K1h/XNYJ0KKR5py
jJBM1n5vKbnP2vztK0uDEYaPgCvN9oOmytSbMUJMgSm4SKkhyZxfAWUGXhRvxNy/
bfXm2UYcsDa3UNyKrQ0w22pEkdPfGrKEvktKW4lkK78+S/et0E0FXbTPRUpX0lE0
VdUVn7o4eiUEUMD4PvKJuzfcwSanz744E+2Oso2ywT7Yw67koS3C42HVQ8k6qgqm
z73smyzTDpIKLSbF3qmMYIz+PSsVYo9D+EtscRnES9qphq9WJnhdjhXVfVxy3tvy
t4nAW1LTgviusGHFOQwB8s0/V9UcmKWFJ4QXTu29EbBHR7QFT/rT6+1vM8o66Hos
y8gM8Bei2tKqie/nwKngtgJNgetyMWON0zEVRj7gCNn3axuJpVz+hL/zYqnauscv
03ZxYcjmbN05PF4GCgZOv58c3GqmuqQJ9AiAVBnJKx0I7w57hdr/HGoT6LwyUDkU
NOO2j8vWuJDfuHKUXzVziSv4Y/jZ/erqlClyZEaMEa8ytcevZkVachOwHociUrzi
iNQqOb6jivHfRU6S44aGNS/dbXz4eSGGcQO1bbTtTPUT5fnlWxGP64E3PihSDZmm
iu/OpGVikWDjMdloEUp137QXEOOQTHIXvCUN1W5PGp2B/mlxawXbKLD58+y3F05P
i7RVJnXoKeJmNgDEzS1do+IX1IaNA6PAV8rBPvnAaFQsktEVd42T+WHF+Fzn1gA9
5SKieo0ixBRsodi/zHEewtwy8hP8Ftm3AGu0twmhrvO685q4kpYBWZLedZvFm9LP
veTMxRK9jbWpO7VfPBMhhj6SHPO6pSusxQqdfuBCy0XuYawnlyM6I/o66J1FjzoD
38EVCwm3q8Uv1hXiHg/uxyVrqr2JPcNw4qNJ06nMA9hi3EzkP4IqvE09jiSc0l56
K4C/PhqNaHWedM90m3FdEeg6ta9Lqc4ekZSZToCvJmCDDN6sLhuzPJHLv9n3Agcl
CcYkmxnGPbco6ZAfCGFa1FDO/zbnbxgA8fSpQN/L5I5wnhC6iADrGSyLP3AmqCjf
kgmtCr5OVu6WV0/p7AlxHj8IJ0+poZ1780TyG7nh0TS/64WZ/Kh0k7PbiT/Pms7z
mm1wP2eisG76uVujnmNJZq4VS0BdnDAoz5cyQJxy+HDIUjmaxOBlU6fm9Fzfuw89
m0WrSKF96CdgimL9IbFCD3ZX+Vb5AmNNorYuApvirZl8G0voRHz7grgxqSW5fpHF
IvOolFJCuwoTGpqTMW7o+fUYc3AEQRYQym6jRXsMFd1/mGPi0IDz5wJp5+e3ade9
2eVHiJgt4eWFWHZRwpyUQ40fmxz/QzrVO1I/gSbnSwDJnEzRqhq+0zdsyotHcBve
L5U18p7+hdoWWXTmW49mm4E5tGFCZSUOFFMazE5aN1LXVAW+eazRmDZcc0iW5zD+
gx+LGUAqzeZsddBaZBavLxaObFnd0EdglgGxYLlcOf/2ZnJEq1qmuo8rUpY5GKcA
6EMfpNKSwX69atlu78WkoxvwJxa3QcJv/tRnUNzUcQFvYdmzQ6nNw2zujX/GLapY
FoDDBmb6tIhzUgLrYkUS72QNEXmAPLhsnD3xbwrHP7d811Dx332tqGapVhoW5W1u
QS72A5lXQetBssJTfXC3KcYSDGqKTZ9oyQS1ghBYMXnRR0EcL71z9+o5cEq3LBDy
3YSygTb50BKTClFW7GuY8XwuAn9qpvdGfOHaUDe41BvV+e00jpuIKY/vdj2Ot4sV
+jhGUgYn+yVklg97vUiPwGDM9kAJ/f7w6uqjjsH3aOYSYgHF4xfuH3ytUSFZa8HQ
P1dvIfvUIJrCylggD81HNOOzHdWuviSahHRG1wsCOTgbnwpBJMJn9OuFxJOW67NR
ZdI3CV6AbPlqaLg32lHeSTxok3LSPx+YJ+SwWvt6l96Nk4Yv2diPmn8xFE2kZiFG
8vOkpwslnQ4qEsdjh/m7ANFKTjaK8Lt9zM6hoWNBvlBj/mvWqUCeZlsSUVx0ZrXW
07sosJbPsB0vxarKL8TW6jRWm2iGh1KxVXSPf+bs6arH6L3hiubYO6oJzuZn/yr1
oORNv4ZxRNRmCTyOr/7OB6wkGgeJ1GtK4ByoIAsvkORYCweshRoyv0R2811rfkt2
Fs0NXjH684y1wFJnA1SVb1rHqO4HPltXWqlk+gfm20U7dhGRoBE+dZjwpO/EU3R9
pL0/AOfFJcGcdOA4baaaYUAHJaQk1hTHUNOV5qm/A35TAEJ07ANIdpZmqIgSiySE
a5bjzo8/Vg7Q78QzCNaMAkrsQeFLXNsvV79Dg6184LZNNpElZpiN9hhNQaY+tsGe
tVGnti09CGlctyg+LWJ4DqpXeJXVkuO+maSuXQFgL9rnKNnDw8wlDnxNhVluLSwQ
qVLthvHWpeO+bxCSpmCRWZyJtW7M9lDq5pfSH0HeiRtCw4dMu94bTXNtgTudGf6G
DCd4GvzOTezTwcvDnFVWjF5O0eL1Nbg6kJW3WXBMVFfIj12DKVVWaMWl8NBkaOn4
216zR097U/sGzEwswI1TUZCaysOmu7OR5kIQfomv9iQYsGAdPKCf1KToKopsgK6I
kdCaWX/Tq3ht8cPxYZjbRj/vCC+1MdNj2zNhgC2dP2RRURujwddTydEoHraoGSV7
vuJvlk7W2PZxtgzn8fnz/JU0+3l367pl1ypp33NXGvnBHJwdWnHqIL2Wl1kzNKZQ
j4xUAjJuZUQ/Tze3P9UD5HHKJvHlCxM6xQDGvwzxE+vwiudbg7DU6A4PbYTsxXxk
dHa4SAa1DBbjhWgVc0qck0eZCMjQgu50s/FGR05qiSHQ/4RRr3+VjeFfxlOuRCOh
+ZkazjbV1biL6VyFZcbeMjJSfJKnx8dkU+go8j+sPkDAK8rp84MrN7ABBz6zLFaD
ily5aIsocCVtR62WmhC2SR/1umSL7d14PHkscwyr3VX5yEdU22PjeH1s01T2AHZb
XnMW+8HJ+cncXmITTO19AViU8jynbHza+ad3WCj4yrDGF7EfbourdSc+6V2bZvoR
An+JhaSeozm8a50yMtmO6hIHHABBwTeXwq7C5rhdbRz9Wa3eiPAe/oZ/bS7oF9/E
//Y+e3vXbHVPnqcEoLVFru6aSW7n3qJSjZFFvaNDDUpzwlWSMqIvqSEEyo1i1foi
B/9Gy0b9AgQPoU069qI1LjyWG0V2LwLM+lONmK2ISvQomOfngkvVdrrf8VVsivzw
az7V6nwUtv/kOPNKkHzk54f1ae34zx3JdBjCcgMC5kJ6wAvfde2E6fcrhtospxkL
kLJ81RMDYPZ25qK9hoR/NjWHwTIFjklCXv1xRxRBDUF8cXMXcpmLY6T03ktLzLsn
uZFs7QodRxDISHvogDUUd09DKY1UfWZsgNUaOu1kj+4035Bj0aKJXyC7jGjoTHRS
n38LPMh5C1j8gHJHe0U0LtU89IhDoSiDy2DT9c0cvTi6BLsIEKcNNzfAC4i1Dwqi
f2ipdopXbdB6e9+NWD8LTZ26st2H6FXU3tsBouZa31FU/TMuycCAw3uU4kUN09vk
awrssfIhkHFenj5wLFAIaVudRb/rtUa8s8WH1zaUemHClpDz/YidTC9izP++9dGC
cmTkk9X2YjXzTPm8AiD6La8n7NnsV7EhdWiy8vv2se116zsRDCJsNYUcEN9pO2Uv
JxBXXlE6MLEJ89xzb61S9Mn0vxgNeY9Lbx5jW0axxQXo9oJqoMggUqdLHxAMw5Bb
KdWDIfu1mB6MTzvVP41XmQ48O8eWkAPDNQLZbs3QCtDduvDlb/+0H6+F27Fm4gNh
jOLFVR5dfrv+z4Y4HGdu51yBfvElda+D7gWs6koPprr84nLNIYOJi6yPpeO24LlM
KONXwG3kh1ohkmqhlLWla60kXPYUmxl1UXLOis7jr6t5WdEW8mPYR9MuQL4jOTMz
XLznLC7+QxmntQr4jUte+UXSN58PxuRUocO95f5SvOhY+bHYFMsKzwRk8UVwQYS3
Pgz/pKc+a+UaYvqaMC+3G5KzajRW6rHj6PnSEQcHEv48LD+310Wavzk7W9pvKCOI
2PRUZYqiBBC14C6TSr6UpdxkLLPFtXWP3s+y5p03GH8TKY6gK/gSI63g9kFPA1N6
IT4PcefmO+eaNF7TWz6shU5Oh1LU3zg+0aYajbqBykJA0fpOnLcrhTas3DL2fNen
YGehIKxSbhIVwwh4HKSI8jfX7nwdyNrgspRaJBZNkkW/lB2V5VJ7EYB2/ZgX9MoG
8GWUkGohomKb+FkSvmUU19kwjI3Si3gSYEY7JinOHJQ/G7nlrvFha1uOC7fmTCso
ryptxU0lwQugdfHX34a86Ce0hdOfmPjNXR+Vfdn2lgkSGE+LAcGZEXznivvhjWP8
kXyIQRYpIHFcl6quknSAN6be+rquIBNwJ1gvir8Rae2m3GPtkwtE/+J2cb7yXZVL
HPEIBSOdJe5jGJjJliiFGLHZvO4In1dXhYTRXkjdveXWawRO5sQGq5C5T4/wTxGA
iS6J27dTqSuEdl9osGAKMa11S95TZ4BnGpcCjjzxemCZjIL/THh7D8JuvFBJFyiU
JX0pie98WyV0ZTJBrrTBqTI95QXPwjnMJBwA6a7fbsq9agY4NRGcLrKpAuvRYK3W
hPt08nN4iMhYURrBQntojoZxFEJFlOgVMti56wQepsmZSyCoq1nKHzqvk2L4fIsN
DvW+CuVoUKrrZzuFOfegeA9oijfHDp9JeF8ooYKEDyWR4WAk1j0h7SNbNFCyFLQm
urVMXzfbSsQ/iRGN9TphucqSzsipuH8szPWe+OsZzqFRvTjm6uiUIBCpc+3oOUyD
aBCalrZQ0lOTz3OQ5RjoKaynjowTtW88JmBFv5BJvBEyFOR9P7nZ7kChpyJwnqBq
5EmrK2t6ddFaptz90hdLo2vmnK/Uk0a5ppApJWsdyotsm9SQonbT7hS13ynCEgsc
eYms8rNn2pz6jI/MqNGtx8W+2Vhge7apSfWIyQ8GOCwH393N0xMhU9KKfBrZdPv3
mKSglmUXl/ce4k7P4agTloWFgd55qNwyA+n7B15txYpBSzugXNe0hQwQV4I1wGZj
e8d/ugWtMhT4XPIciWfgGX7VF5wtdhX40P/OOwOI11umJyh8tM6uavqxt1RyPAiv
9bXgP6Ohxh6cWPZgMXXTb+pwDiQTmIQkJ5Eic17JKmrvbexx8CvuTBy6PR3k/4Vt
jKoslVQKw6+O7H15tH/e/adYgbmB4bJVI0pIHQZdGqT/fQ+2xfHrjKgBM3JA7q+J
/y7f32cETKjBxq45Erxb8Nr1g8hPcO89hWxbBfobEiuTJ2fOUn2pqWReC7kWAyva
YXOU2GymX+QO8GNrYjUTSmzIhcMj5rD2N0WYRUVn3dPhci1t2kLYjwejTfTtiJMi
yc2WrfDOAEj8OABSBu0u2tCKDRQB+p9ImdHXb1Bbt3pf8ZJkerWR9bZHxLsWo5U8
xcVNjOQOxIndgOBLKvefZ14Ol/JxkwWneEgZkHGAXisEcODvahlX2CN4maeFnyeN
xLnDtNw1WpO55DhDbJrPC1Y5RS4ketzRC5uckcVKcM/lpRFK1Cmzp4fQNUHZF0Ra
3t5vtiJWO6YV/QnMKmwfwyvtMyOMdKjRVSs2Y4a1YWgyyyUSsmPUcG+RWIlhAcqK
Iq3jIfd6cOTwSQ2OJHRa29OhObT5NPN2cxExXhCzwdHePRXYvlouL8ssPMUcMJTb
1b96X0gZHcGUJyalziK+fCrET10Vye/QCCjGV96AiFO9W/dG5Y0X7bgx1Ab8kSGl
in72wNelfOoBN8hE1s+lovlLerp/4wqx0exRvhEhqYNdeCLj2ZEfU917PCXsGHyl
tXGMI9IleORMzUM4m5ifbszZrLhTtf4SA8+Jq7YDhEbEdU1nEpibvwW4JCjWESti
UNDpiTQ4Kc2IbJ577eTAbmnhTELGnGc72S8Rhn4Kx0pnQYFR/xAb+QnQbWGvOmuR
QhPi5jDNmN0c3/cEJIQyQUyExnuEAqGaBdvGbJJ6XSJq8rMeKS6S3gxBRLepO+h2
Sh746thbev3jRDFy2D2Go2wDlwLAmKspVsM13NbIwhv0buu58jxX5lgiVhdFOw+5
sZPoL4JddPHJNSqJpIxEhcVn6NZG8dy8Dloe9EqO+6Fcy2VSaSCNuYOSDAjxIBMw
w0vgU5ssYA/JUZCbVqSN2lmGPjYajCigIeFEBkAzYTxwF8c2VNWV9o6zI88zx0HA
hqeSlwhc7i6kfmYzd2TPCc3OweRV9mzNH+4jXcck8ATJUofRFSwIxuMjO7xkiDtt
NZx+JJmFKTZLxXQWag/gAkKZF2MHlFqqmYqtwdI4GZOSbJwUgWOrX1NhGV629xbo
M+39J1tFiyCXPobWmueA3fRyLuCYrSDJCIhcYb3C3Jj3uUz1PTwfXynvwxvsMFtO
Hal51VtQ1CuxhxiGUc4QY4VKXslaYZkK1sMuqG3rXiXgQzr5ygDzloo37z9Fpzxt
26NDtH+PTa2w3tbn0zyqe0Gzu4ytvfZ8AC0wb2n+fmz4t7RVSdR8ecEtyUlLgNHB
upKhHrsFLhxfMAV2foqkYLPermd0hpsfo8ZIwGKPQD3uf4IIwtvTt2fSuN68Z7ps
iR5NgcZ5pI8CQxkd3wVYUskYUYirJ/6szqNc/SQy3SaJFkj/l9dAXlP62gcXD1Z6
ZrIwCq7zQ/j3kG57IaVVzXXL1IYnLwjUC77zznYzsf7J+7J7Q1YyJUnni+4JDSml
NsTCu+zGFNS/Wpn2wjgggALn/HIK4JCStxzhgpQms+ICGcVFIuFdrttBelh1OwDb
tmYUBZuY//UyToVns6f09dU6xp4vdgBhyFWQBEqjnykw3qL9xf+tHbszLz/jXbzy
uniKbgsII1u9PFMQtY8VJQx2TQlShQwzP3D+Svx6Xh7yMzrB/lOLWHZtIBGmq4NS
WnLBbn2owtIfsVAXeRMu0q0S+zjnXnVkl8oehmusMnqI+Fn61VDTLD7yjDcVcmAL
EDUrre1FeMlnEOUpuJGmOXWS8ZpCN3kKlNRFu0iFF8MDmEiaq5eAhEX9VIWYNVhB
9U/f42QlXm/dAPqCTqO4AhofeLDXBW/fXR2YUzZEFk2ldetSWu6QVZVwKT4Pz3Gw
Tb69PEb4AUUQRNJ/0c+F49AkAvqywN2hF6xYsZHp1UEW4k5D0i+9M3LEuJ7lJeoQ
QlqOm4ME51Bg+9NWuI6ztaYzq+FxZnf390/qB4MFtbxv85E4ZCIjYLII1KT+tpiX
v0mrqSLYyfLxQU/+IaUtoQNyON73nYnXQcEJeBV9GMBxHxlFZTmxt70ZteUQlDwd
y0khQFrwPBAHBqrNR310L7f9NZt6C3ZZE6D1muWOoqF2NTgXwAbwVNZROgO2Fr1W
6s7KUVcXGxFxG4Lud16WmL2wfBl9dP8/phQPblJcZoE+C8Gv79DiBoqdHga3KxJF
06MO764Bi/ysXUpYZjopVX/rFIQSV2KWl8EWlai2AYUB91TByGsybSm/dhzQC/lS
WJvD1MF3kV9oQjuCcSeMs7HqjgQWyGR5sP2Oj0EG5WfRp6ri9k4TcIt77UKkxRWH
pYhzt69ZgJSLXI6YeQCiHUPXjRuX51sJ4QELR1gE0H/EwBvobGrJKb4rdWV0z9QJ
BhkBqU1hIJTuY4n3DPRNbQhgUwijlLiUr39zVhqu1155Nl9lfrGl6Zb7o/uF8WS0
FXO8stRRIZM0HLgEAWuWylckZhQj/oW/Me+Cc/Kzly/yJTZ01Dcp6wgHutl1WmeI
/mkTTCC3RgIEaSdtYnmPThlMy1OG3e4Il0VRwr95DuDLoT+aMW7lnFdEsmd08uVQ
cB+M2Fgg9er2S68TkiDVsbUd375EEi4uW05NlwbActhhVHxkP2uwhahYPZ+FvzUF
2SpFXIQTLj+AXgi9/2o7WF+o+tzzAyRrWE0GQIozzm9zC6JHOFSZ5MMkGGPp6eD5
LPFPZ9Bv2Y+ItDz/z70ZlSqV6YpIzjd3kZl3Ww01YcA4LV3oShqKA17x122Q6fLV
2zI7C6lax3IbYe0DxDYyFs2lF2K7Kzhdex5YLfk41u1RT0JykkwE/XBrCKx/WD+b
e57iQlctJkwGfZ0VNpx2d/9PG2+QTEpQLQBOmJ0mWPUZKWl6sChY5Sx9CyCFakEV
PuS4eMvoCZF7TJfv3LtqD7N1gOjSewk6GzIjt3hqlNZvvrUVBiusJrUMmTNYQ+7q
6mwB8LO64+tflUvOVRflXWz0R7GUEQj1DXyHRIwkoIZNSWyUQzpg4WQxrJ/+rcms
pQKmAO0R2AD+Ed1Z4qCJ4xlLRR1xeIBtP9M62/Hm/wD9GaI1UkK2r4JJ/LOyXFXl
hPpTHMK4qqNJv+xZj0wXhdi7zTx7fm0vjcoGSpRsd77KeNfnUl5Rvw0L+Je8PKZb
gK+wvVqVOTVuWjqR2qj+XNXHtX/iAsnyjqmZ+bJrdEGdedtjio5kOhkCnYYU0d8C
B4vjn04JMM7PXeahE3MuyworAfXQ8xb6MC1SVONhvcryRO8XJNsdqS1xtx0hKYwd
yhaGcUPQqPgwsq0lUknhy7wlcvuIMdQgDnXFGif48Iw/SmWMG1SQNGDDk+RhV9ot
Di6oCS/kk5SLMjQyLctz0RxfUnZ/7gdIAOCiKMlLLlgarMyQSz+f6McZIP9GOlV2
f8+KCpu22/8vIL5eL06ToT8THRRpac6yZnIX6lkLjZx0Wt+pjSFFZaIzcTCJeYaC
65A474VztH8Wp6D9WQDjRts3Y98A2pz/arf17wcQf/QvKZiNRDOnMaKtUF1wUurN
Nvi/U4JENsxyeUyUE5KfikclkwFHklrfxFLHb+hjp4tA3DSfbL5B4zBSFZWjW9/8
uofgI7YCVIUcKv4YaU4h3ykhj2pv0yaP8eFTq6zw3Gt0OVHPcy0ce1/2J6BwUSf0
DM2Q4iZWivuQiQZbV0B7RFRrPYLRrIa2pM2S8wXEgmoobzdobAEGoT52b1vWsZQg
jbq2PKCJr+LxxxpQE7o2ohi3jOsxwAz79AwWez7NOIdVYXOLhc2+g0cFu5jMEaro
PPVU1bzjNHt40GVB7zEUwXEii5Gi35F3bKLy+Mx6/DFSynZ/Urdh7hotzGN0bbTc
+gZEg8Ukj+MbRC/EhvS00j4MhLj91hw8yH49eh98lrVXnTcutGm7oDtLjK+mtbs3
KxZQ4zEGxQL26Mrrd6EiWoXUzgmbtH3cdIQA8NlYjgn8lO6BS93QG5O8Pngv6Npg
CdlJB0oVbfgg301QCzdIRuLKF47jdD8j2GAY6fTag7C4vEZCXC7yBuNJMNHW5L0P
AZpSA2stdwdckO5yxLyj+UjiTMk/vaHtE0J5jIHeRUPZ8YzoMAWMByhB3CoAvGjp
lXzs0bHo8OmG20jnn2rGxtXD/HSMlQwPRdTDpVMbdb+/kF7HrXkZu0M3v1lLLP2a
HDnPx7HxH9FPYOJ25g0A7Tr8oktEFS0325RZozZrS+KiLU/36beNeYNNmiQmcLY7
Pjb3lA+ceyvCLxx3VN4C2K+5tD2yyybqhTw40eJdJYrQe1uRzGRcvbCcaNXi6gKc
eqPipT4YdPlESxGRtHe3gA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
W4xIcLAGBD8bUOrVS+fXcTQTkyhnk+f/lg2XBAAEMa/kcMvBTKBkgxUnojFBuMQY
tJ65EITvYXYG19nMV4GBFv1dvuyjmvQMDT69OaDuxdjqQVMeNBi2JmaIBD9AbNoz
vpWK8FaA3zo4+aLBpXZyBcZAlV6MW00Fsc8UjrwTGIoVkeiDjbOckQqZMdsGJx6J
Xn2/yAtivucTOAKH1nY+wy8XbA0nnuyfnD0mE62jcowC6SPqvGvsr2adVJB4ZFbK
2LSIHASjsa064ZlkmzQhUsi14vLkr/DWq/jMBqGueuTPskVh/VGsgJdVZ6566+Hy
tuXTdfICa3ocZAW/JRaZ1A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 27200 )
`pragma protect data_block
TxiUe4/dyiXajnyiV35eaw/MzDKOkbLktd6TmdC6I2tefwnF88WdTJyoL1gfY0Lw
H5imyVCQexAIm11FeFVie1s8A+cHgKpHkl5yA6wrUOqm1rz35ojvwPlYEJ2GNqhC
jf7q7EuxBLpJ+i85uuMOsWhDCljTR+GDlImdSjf5RFsk5q8QwRZXivUiNHZwsvPt
2AJ5iCwarOCuXm5rTy3wxwJTonrUPhUWia7D/ZrOE4RJIND5v4wENcnfq7e1Q2RF
gqBzDKCfhrdUnMd//YZGBgNiAKz7eIQ6hBMKtBHPAb99cK/30S9dDmXSb13P/7Wh
8m/QY4rZkNT10WO49qd75pS7GkygKrM0p28426m2mgKPncxy+9acZ4Gf/Xw4zdZR
lvCynzNhHBvQge2YaMQpC1kl4/LXixijqtwWHn3c2xa8qF32wKQRYYfNRtGjcwVp
MNVwz1Dmv1WJFgS2ZIQAvJZicyXIBmKKyolEuvtuu3b+95pB52XoGMdGXDA8zgHV
9EopCHNjpYN3oQ2OoUPCmGy9DL1wrItSgSh0onZ0UZ40seKSghQC2O7LdJkyXF4E
Bkb+hs+QhxUT7Abmp+QOuyheabBGEXbBaklNiF9G0SWGHEQH/w2T+8fq0ZlZsDoV
y0V8TLIlUHq2n+J2X7kMmgStzLm99ryy+6Pwekhwe/R73aTnl/6bv5Yv4YPWh0vL
d7sfdkZBPCJIeuyDfp9uOZf6RAinnloZf5v3gV0LrnYKKWEiDiaE6c5eLHqLfmiB
k4SwT3Rqql/IAMvKLdU4YUH/jUzByr3W3/QMA0pnbBBik9i+w+J+lv22nvEo3wer
zw9xSBjsf8bn4PqoA+65W3xSmOJ0ISv6Avw76Pex6hoGs1EP1pTy1Jt8JVK5MwCx
32DDutcRjCvpxV/I1egIXdcZt9nvXJoH99Y2lKMkSSAVUAOAnknUscm0V4MMVc0V
rO+hGtZYADL3L9cCHOd7lhIAuqHr+Int5p/bu81Y6hIwRR5rs5huYGwbS1AXaHfx
PiHsro9Ozjy8WJ/T+CaUV/kGTXZbgadrRSmnSfxQGi3lU14LMCcneOuNbrNRLeIU
pu8qXGS1K1Q4KiIh4kDfaCb1MFMqV+H3nRSsKhMnRNmzaAMu+/ibWsTJRHXmr3cW
pkh8V6e6wHLhOCqFUbmVAqvmOZ6nUs/FyRlfhMuXrVJTX+A+lumPMqiZzll300GK
DbeAE5/F42GusydEXVf0soBKFG+7w0BdIVNIQxCyRExTLTnnMijCmCq2AjAkaVVN
qYHxSLIriRur4eEvGPTiTXB5NxfqH8lcBOJrFnOO4NzNCIrxD6wRY9LlGmotEqrZ
wgfJZbIZa8/mRTQhx49ROSIyl6OS4MqULJD+54IKuQLYR0Zz7eNgoQJNC2PP9mOa
BkOTkS1I1nbzTYpUzKjHFLsCKEFEZ6Bs6MQv3KA4tqA4SIXE+eLMBCJSRP9nyNJQ
1mCwJoMAgYdBo+N5nWejOMkt4DGWeOzAxvVtwvY4rP2Qzjdo2hiilmZOfU+xadrK
S1CAonDP6mwWxVcZ6bQ3QlrGJHJacPi8GtXFXlVCcSPAOfBpQz8Up3rDYnp+CDK6
tPInmCnAMZPjSqxLgwy0w2UcgY38iCbcPUPorgvhNwCq9hEooxJR+Uf53qquechs
GYe1nXwXOaubswZ7refbjmR3IHVu88hYgsw8vNbrQ9MO7lEYQx4tMkKSusk8vwig
w8Nkq1inyUD5kdRvat8WHNERPTbDG6GtLgH2PA8p3xGc+xTMHOh/M2XU0+QtZTkr
8f2trWSCj+FwKzDtuzin+B8K0t/LMwn8USf0ZT9MrwSe2yyhbLsv6v0o/UqXtqDz
mjyXqYfUr5fLGHDh5PU0lADePoMviQjSX4QLIEFXIUJ6joqLEkQo+9iu/cZJI6Jc
tR+O69q0tp7O8hDgNetIicZ+HTFJalgSAUw58Ezak5RDvLdgmAR70ZMIP4mpCsXT
sI7xSbo1YuFvc51fUXEOhMShKcSC10Sxuu3GbUzlXJc3XBJJh/zxpe6QZpWtY4jQ
MsIA6qlAEfequ4uo6Os5f8zS379Sqg6FAv0eQiNU5tLpvlFRNZjjIEf1T/gIll4f
6U7zH/Vmh8r7LkZVeGf6ql4p1LU84blLXNArctgKoMvMQ/LhHe4rmGetglWW11Wd
4FrRi8MnEUjIW/TXlC4mwJ4gCGFfS3Jr6QSx+RPoBt/nvj1M/5hlQoeqMjlwLPzf
qzulUPUbh7rI+5DEkSXHgA3hhbZvEUlNiyLmOPDZBVWhxcuqY6VwQhJw/6us5wY/
c7yNCB3yCW8SrxoPXEPj37b8gPqTLrHV0+95/eZ84+qLang7n1uLINQAhZ8/PakK
hGz2nAu5BYEWe8TLyS2GOGngAApZF1zQHrwEXHqcJRrxksv424thkqqWUWZdQ5Po
Q/QU/SZVBPtrvLn2FiOtwaKGYW43EUKxLwCfD8W/RsmwVDxeQZc54yVwrSuIKwNO
suhYzfJwZwX7Dnja507jUF0DUJypnyUwiQo38+jhTuuAMNJvB30D1nr8M/Fjzeut
sxCHfrQpWttwaRo2T1mawvtmdBfeMRvvdDN7VFRtYrYL8pbkMlY0XVKcSk9hFVHa
GRKJe06H6zYa1/Qu5a+Z0O1zYu43EEc5pjXhjno59dOMVDHsCHaQ6c4VQHs53Z3L
ZYEE7oyWJ4ByvGG9Qc+mnPfcAo4k+fNAMPN1Lx+LMe+rWYL4/i97MdkXSsyj2M+G
KR0y1jOORPDmPrNRz0BfuM4Ej3iNgIE0g+T1xxKyZ0SantKar4uCzMpqM27uZIWZ
HbKS54PIJ0DpmKDuBbAkI3arSuacM5jnBIIGKhR3QWOZLwPV1urjeF1E3kEVe9g/
AIV4+8KvbDWEBFORSoYi4OcS+cmvej/D6m3ZmLyxzOiWVJ+HYDANwB4U2u7Yumq7
4wPuJNmDxPWM35ieabXGGZTu9FVCHy95sbBL8jttD/rGZpeCJkbwabsUrq0MkL9X
Uml0fNvW4yazlKFI8HBtoxZBfBwwxEl9Y1wiL66BEQ71uoOzjJJ7xbF86pc8Jrss
KaXFt0wHAEQvv6SdAjA/hPNW9139IfUWP2OdtgoOXuCWT52M4qFBBLCQ2VRx4Ti3
MUwsRz9NFVlVMmgMMOu270XtErHEVnMzFU+4pR6p3vrEMz0Oi2FmM0NtRnEV6mLO
3ICaIanRNkV3UOv/q8+uQaLnwho13qqVgcGLoByqigk2I7WrQHh8GPeXUJk6Bc17
34zJJpWxrpOeH4TNmzf3pKumfsGz8jrepx12apEVikHpTuPVq6ZVvN18eQUoa4cD
YZq7WugjcXhf1dyorYSSmDVAFzBWaoAL72rknolX5EgPBpnCoWf76sHwTtN2xdwO
hgZF/3tH3PMko5Ys8bVfk1HiaNWPiEHEadVC8V6TDbd6qA0Gx9/ywfYx8IF1kENg
On0UMwobaa7vl7abjE9vz4gMV1Eb80sQlgIChG56KBzSXsQccwvEqnll9uFBk4AR
k3WP/+B2d6NCYurkJzIRksvEvAfsjxJ8GBTdxJW/xVIzmyEABy4HDlluTuF+zbpX
OoHHgUkZ1sG6k+9j7iShCwxW9+b7JHGpEg37fMwvrS0dyv+00Rkoi92ZlzvN1eon
Oyo0IIjWeS1P5Kvf+FecYen6DJxNYBHrwxnntTaui9q86lu1gDBGUcLyYA2itXip
feMI00ajnQQq8TbTgOY5jdqQeoKC853ACS2EXqpENihpMCJJ/Sg7qSR2Dg9yP/8R
XxVeysjq3wmbXv2IeVcVSVfDNc1JUSYlsn6GNit+0gN2BPNao0ZBPTqXuAeeKWzP
TJFPfOYqOXD4J7I+MYvqotBHLgLlQmR7QQfimRgWe2B+Qiyt/tcl0sl5Wk0NKTtP
yep56wgj0R7qqYLtIt8IaWkWO2ts4/XtXSGLBx40tpGcb48LaE1UMjQe4mEL7k3V
ECNvU+w99YwKK94RShyRbNaQ+wqpn0wuP0RWLzW6cJuj0BI9L2HToNrbVmW2ydfF
NgAnrWsWMoszxEWAYuxlfGcLQaN2zf15eNl3w0R2ZMhaGG0izpsy2xmiZj7fYxtC
5JwJSRiGuWJJ0WSG70O759WnpPGb9PNzAGVMpoIIMTzF2fLH7Oxm41bnukUwwoto
vXA7so+9LOFHjCqCYsPvexEAghzgLGDDL8BHDqVvxEpVf3pgGS0lGt1YhA5zg1vt
6OnA0diudH6npzIx4FMa3V+Gb0vh3wIargbi+mDpeyD0DiuipA0taKagOZXvDDQ8
VfUBBYrBvZRFHxEAt0WsZ3/zEtcYSBkzQurKhJlajqkX/cWMK2py1s/kY6uaRoBZ
fYmxeDgblqRIzy9RFuhaiRha9APDGrM3liQk613af3VKaSwXjwGXCW2rBJdEsFFZ
T9vI+fkmEMrUWOhMu9C1+5EJxrk/XgKX9QuXiq5laukcxx9VT6nPHLj6a+Wc7JOq
PiQnwOeEfu3Y+xW3CaSiV2Cb32yANMGgDkmDJqFQKAf3asOsAkOz+Qcd2GCYXoe/
VPmqvI2F7vB7iiar5lMLMW8qd5BPoAztypc6NvBoZcghNoZJh7Rho+2hDpEwcTxj
qukKI+7tw/Gin+jWXPPCoQ4IdM8Z55JmqV+aj/2rqtTT5fNR+eSzu+dcDBlceocG
H6HKJgeVs5g/oJtrOIjvT/zV07tkxv7lnGxI2RZDbGbtzFWGrWb0hJ2Uo6RWA0wq
0B9GmUTBk2AjZBy9pQHw8SbObzIH1oTeoyaATbF9vlq95TX4vq/Sbl2SE7hBHSKV
RQXRP+1QOizQkwpd1nTz29kyzcXge+FUyx9C9Csol0Vg0iGYjy1joDef3BASdLbi
DCMTlNrYJMRDTIGsQpje0kGW7RKUADuB8e0ri6pJeURDprBxdrVlSR0xSI+hXMjM
Hzt+WDsXIdOeI3mCE4xx1nt7PfEQl2znZrYm9zK5z8IhwdzhDb+6OEbPXQk48R1l
mvbQdYgGJlz/5lv5heQy2y7MYrW+Fus7vnV/Tx/MiS3cPTIkDiSaVn60OLcbnL3b
Ti9effehChLqAirLxCcNI4jHP2WY+2J/xTxiOhsoZaxvkq5onKnZi4hMrnVuBMcM
HCocLJKI79y6wucOpGHoIeKzefOO0h9mg5Mja9RfMkwFHqXu92StZ6KUZBRzj5yL
0HlCw1bh2uWufIh0TJtrJKB4WCY2tVOGva3lWuwb0IVErrYeTr/bWz98Qi6tiKlx
CDNT+/6ecn7qi6FatIgHuAgkdBh/KD2GuL0kWD8S0kDGcMai3t1orwO0rnl/Hlbq
b8qUXmCPFE0g6yZGy+ff7ZuDpXXa9Q7ZQ984FiWrkdobitH5DqTGZV2S1U8bUgHh
sgpnj0/FpKISMnirbT9coBCbftZKAl5xsHHoQTQv/oeGfbyjKtFV5LRu4bsRo9Fm
YpClR5qT4zLUSp+zDdQxR9CcqEXl3TgC+R/0W1eThYQoGC5ZN7gAVy5udSqy37M0
1FBuYSFfyL9nnFoT61NSYxGB/CHxwz+BQtsv4kDhQYLQ8ejIuWXRZiBPIsb/GJxP
CrUlIFTUXJsEVtSF3SNErxB8rG+9MLtH5U4cXFzbbRVzzoki2G9Hna57kaXx80jc
L2SWVDHg2+KnLJkbXODDZfZlHsNGiMDYuzlIgAgQ2pPzehdOvNV4fnqtHadMNWKj
1kNNNn8roXAyP0DNB4zGuFJpaWBsbzngPnLnLANPklmr7D7bU31GeDk2TotkCJ3D
3pgKU4A/5xmVDBnFqAc41dcy+X8oy3GXZqMuZSjl7qcRLcRhRpvqxaBcmd6Slwqb
ibbc3X7lTS3PGzC+L5OI+lh8PY2IDgZs027RrBrQRwANDUqfl9SMnrSN51FyLBEE
gM5B+mwI6hpPu/+K4in0NT2BJflKD7NeAymr0fJAyn0Y0u/WiRSXszsbQ1STr7AX
z1TSKQswI6neKEuZfxxOFSAOba4z2BnhXNxQGksIvQ3FZFCYRdHAK7o6s7QHLSHu
cwPYP1DS5BtPug7GPkMb6vj/xs90/3ZDeIOOBV+PhQ7tKlzz4/IAiU4+MPClLCCs
WfQrmmGI0+xiNyD4gdFMOE61BDiVtE4gobC7GMSeoA0/xr1m8pLEYrDfbEqioHba
C4iMyLNhaT/boVoQcvdr7SkuysKkbZRA8+36G8Y/KuIteXl2sxjU8NhPegN6ps+0
8aqfjTw9JAnKz8c9SwPhKGK2R/0JDxD8semowaRYOXF0Xm8J5GNSu63tyEO8SD5Z
T8TuoDsiBrXdwWTMfmln5D762H9bWVTqyp+8yokCM6hFfvr72NMw+y/wrYK7n4cB
TlmfBUfEsY8xMO7d74qkvnANDaq3F1env/ulc26M08QxyGzRREVF7M/uI3yWyvai
Ywo0kxoz60AkebCoqwZ1mSfgkgmNkJqFITfbY6zRWYUZkQeRlu3NkXq40l69mSdo
bltHKsw+nqcKJTz2KP4pJcRziLKSL+HWlxBClt3Kd7bepDpOTh4RUA7DSotY9Zt3
YqIYKB4KZFRPt5p3hFsNJfQGgvz8EklmRFmeR5FlOmZKL7zN6zGC70+H2GnunFYU
j7aSCtJnmwLQnzVfciarTnhngIiyyQvxdB5f/ByItDO3QTr/N6Ug5ciREnQcNIWz
zwCtF41+8npn2Ul58Xq5ZjbSvlSzcv7teGS00enKxMe24Cbtau8dk94Yve+yuk6l
xgwZBJVISk9FPUOaz4H7+N6pDioVQK6h4SSBwWPIjEAU42/P5DYIVfKrw8VCJdiB
elDiXZ8g9u7gHyQ723sdnrTA9NhYWHMo6xkn12oVM6TJITOtAkeSBQW10og5dnjK
xEUeUe+W1qSy8q5mM/6grT/B3DK6n4VbOrh5Nd1x3C/Tkdx4MwRY+4AIJGq646jr
6jZL59T9wkN2u/BbZ5LEzcSyjCrWZLrm7+/RABHqlBa0UL0lNjs/u7sH6mY2VVOJ
YphAiIaWCiEoyxQFf+nG6dNwOu4WF5g2WTKyle3jcKRD4pF4T01TRZagHyGlnUcV
p2DlQ8tTSDlpP3oIb6V/nwYHJHdv/cQSZowyXQaDsIOMhfxW/xnpRXRd8GCVcTqf
yIrG6PAJYGFLvyIEETYUQpBx3oKwBYV0TX8B5YMYUQ0Ceq/bIqs1HO4IhmFCeWr7
95VIkMsCkOWqdod0aTPEbC4QQe0y5ORy48ek7B+Qi+z9IV33esgblkVgqdN19G8c
/BAV4H6qKXcUR/ncMpSa6fcpa5duZOgDrzuwNOlZj+JpmtP+PWqjvaa11vwm+JjU
6neQQeaAOXpBFi2xsXE9E3qGnbiksFzyB06xEnsQ3C9+ApvuN4D3L/x8vNPrQrOZ
HVRPaVEbDH431U+8TG2xV9bCNxmZNEKH1YYTyWauNtXGheDJJBAXZxeDkQUoUZRL
qMyGlpLJRm6KiR2OKyQRdOf3mbwGPs/XFEoE0RV0ESHdXyCnJEzzmg30BscR6mtX
MZHxfFu4+tJgSnl66p70U5sbifuJyJcihwWdsVMyMgxXKIZJqQp+P7n4hmWvcsTC
1gj/xPs06kWEGB4vJeW43QUd3x4XRPPLInfaDt0igZGjtKJ1YBnl/B8I/ybzUvSX
ZEJm+NWKJXbSXb6i4L8ZdO35gp81/b2DDbZavR/2UCEBNNhl7vKkKXQXDdLqRJtL
30VjUrinwHGrVkwxdZGOzOiEQWdfjV1t+lEJ++7aZil2F0AjRVd1A2aPJKrEprzl
zKE+NvVmdAxwSLf8dlGev0ZEMLCiG+B8NpohNotfnojh3Bj8tvYXZw64J+OZnVi1
NVXPmHG6lITKEfk/FgMzL9BikPXCU2wgwu2IFaXcRJB8uwlB4rZbrKzax3iAmYi2
ccVywnBaCc9gQ69PfCqClrTKxJzCALwbbXbsOwE2O0mKXmosCOkXZ/eBx8Z9i1DD
qU5jtJsgIT9I2QqXNKDUntrceIrwYJOnU/U+c3IQww9g4zF77Bk2RdaIMCDhOyzi
ne9wZ9duex8ZA2hkel50OuagcrQK6Zl40vLz/k6/SOle7fmHqmZkXIt6CTp2rWql
1slXaYXQ6c6WfaGS0WCxFR9LW42BrtwRxKoF02dnsB28j0NtsAcSBUEV8egefsFv
160GevLAwMgoxQeQEYVAg2Omg0BqVkgEC0k8YDzeDnH+cGkHsL9EA44inYIAZouL
UTVsYk7lt9GZEdlk8SxRp6/Rjg5UsyEd4jsPSBvuPrZvS4kTlC/TjMKDjwUQLfZS
cMZkK1FYQ8IRcGL10gFdknYutu1b05h/kMiSZHDk2xcr88cF7uiazMYRH+w9NXK1
MmYbNl8p3xtPkDIk2NWAS4qB3SwA6GCMUQVW5B2QEZt7bLrCbGEU9PtaRV+Gh9Nk
Z3IEpO4NfgBnsCJ8+HLJ60h5jxJrfeOhzVHUWNCrliO6rkXAxD9MtWlmWWZu78PB
Xk0lTrGVQRce8py4BKXzwVrhYb0r5u5twN3if/LLeYByY6NDOpVWdsNBTwgwHiNB
L62sYmxKOWbgflxaQHKoViE1Y3ysejpiCqC0W9adybf3PJv+Hk0KLxdaOtVhI/Yi
W/2S4Uc2IfkEmectdNMiDtUU7ddJ9WBXKemf0BgrNflaXs/DUWIpwoYT8xR6wfVs
FOHs1FMl8M/bLMP4DMWgJcCiWROEWsW2a8QRGd7859C+9zh+tSB88DJP6wR9H+6m
g7fQtv0qmBC8XBodxbyFxw32hlItYNs8hVxS+8ahJXHYVLcDx9UTtxGzImG4V5r/
rFSkM4TfEcdJBJvCtK3g8J+KSrMDQY5pD4vxkJmphPv+V6LSt2Q9AaEE7wFMit6i
gyt4epKKiAwbvhfBN3q6c4TpYQhlmw4LBBhP7facqeYKHxgo9XmRFCC5zbms4JPJ
vLUvuoTwXyrdiHlkF1Ce61213VKTAFg06NAx5z5fmulWhPe8ZTfAv2USNKFEXc/E
h7uZpv67GOvquryMXvryZAuJNLZWMm1U21esuc7ezbKLYzgPYcHql+mcHG6gyI9K
wHB+K97FekfXVS8fHJueqotXVY0FnfV+7s3H22JZuPkxYtWO/p2h/R/1vkqEDO3/
tUvqJl1dV9Z85HTiHThnn+9jMYkvDD4J8xn6HrA+0fS+jJ35EW+5LSAYX4yAbOgV
WolBwCLctmNsME0hLyyUzgtgfArJuuCJKM1pi1xALrrG48JGecfQpoO/YhmzX5nQ
A75dYKl/zxGvguigRC5G4LOWUg6N+gunkzSMUhRdmdDK99b3F5tBpxxm0Pnz/0GG
vNy1vQLRgcPGcPC7X5JEjpfvfzCfBN54liqQQ5bB9ywGSRYu4cw1/9kJQEH29MzZ
j50lkggdYMiE7u74/VNQeqPxdKlyZpvuD5ErgI5bAoUKc+VuWD1M1BjAZnp+AiXW
vpa2bGD1EXpFFAyfsAk681r1MS7+AUm1jvt67TzHDAr74IHtRejOUaLvBVWb1vlx
ewMVJpMlh26OsJgjWnJBb5ZdIrUOFtvsmTp7KQy+25mQwaJLrytAfSpZjrpX89nj
htT9qkOUOtAfkLUtcDe2nZiYLeE1fOl3MrVQvNqgU5IYVZg5l7HF7z3ITh3NAHu1
4+jqBQ6iOqQ0rSSMcqHggD2IEZt0/Wp66Xto1IHFK8rzAJx7q7LAGJ9NWnl3Xm+e
pSLBs9KfEPt58kg7G/kz/opY95u2fWpHHMHDAbOsO4IgUzUuMs5gPOfcIQuN0Aem
WOMfkytt0A+/AaNYxtczZRMWRDu9C90qDuOXRBAGe/nT7L8S2m1RZ6brlNXCbtqj
wfGppCu4t6FdCHFMeOFP6OLE/KX32x9HV0Tg+mlYGihea90U7Ho07E6WI1j6uUx2
BQrdUd0DbG/Cn3nepPpzvgWmTfLd5nlUvzCuroXcBI2S3TOO0px7epLPP9iNFTS/
eMtOXKtyHtrUBcmY2RF7EZov2JJxcaljLWtlbwCwcrKyVQELOVni5UBJdPInuUod
M08+wvqI0JE6SMCRNZa7JqzRrdNC3+tn/OX/gwarbonIxYejIQGGzCXwrn3P+oEE
xGdVtuo+/buoUPblavRs9cXFCZ4BrfK98IofaRlEfWBXmGw2ElYvRXiBxm+mtP8J
08XyuYS4ZBV5n1cf1mdfKTeIB8l9nOGqP4Bx+Reu0ZpLoJsH0e2IyGkfVswvbLAN
t1L8wR8O48AS9ku4yKNSiHQsshkzw00gYlVb52SkejAvpcpUUY+xGWovLpQ0MjXg
jfCA29p1FfLj2CI7KsmvA3O3NWNLg0Ifa9y/wjwqMnox9VKpwVcfSJIYCp4Smmnu
THFprpzIm100JYM/zhSe4pnWrmTW/jCd1nR19vBJKQVN5H9aj00H2GkoYwAgB5Qo
TyxK/zeyQUySiP8fZMNq6GOt0wJQ/HJ71Movbx4Mv+ST5AitySGhWlZ2FV/5h9OC
bdaGSfR9bgJU7vfNgOXedpGugLqffatWbtFeV16GwtTBaIJc6h3wRIUCcwqMJirt
NrYkr96XkotJ4sWJ9KuBpcorLQ7KTg0j6yTHjtIlHe2fuGa0Z0ckW2YwLpHPXAIg
EU0Ut2Gg/+Rbfs9K/GwnOwSZs30/e91BJADVSRR3446BICjUvxX+Elmju42GxqAv
8MBeCw5zfjElQh6kde9h7IdVQvQpTvFBf7advKhN33VaSN4Kt/klQY3ftKD+KWVR
M0Ty7q6NV2iwQumLmlHnV+q0Xvx4TSnaEgL5AfzgtQogVSfaMnD05JUqKlhqlKw7
Uz8QpMScCeyW/41E+QXmfEBNSVC+uJalA1ArnhtqHmvujqgsXnWci6Gx2OZ1onuO
5ckVYHf/3Q7S2zresGBN9gylTuPDUF2yCA/uJ4UAAc8sQrLvqfVzgRbj+ziC3Az6
g+PZmn5zpOcSHF/lL52uTFIymh8PF9NXGNXJjIbE+H38mlS55l2xesa0KWBS1xLc
d0IA8Cdp7EBZYhl2GWiUw71VthTnsPVjRVr25SsibLhdxJQDi1UXV/1961vqjuKJ
5GuB2+KmLvZPhCZ+iuuIG23xjHKmG+wacWj5dSdDuau+67KkSSOj6AuivPxmW6tu
2XP+BM5lVob/pwUX/TLSlFvMhjo2F3tbS8vFu/HZQRekL5m/wWPMCV1/Vi6hmbpL
77rAiqoTpUnpxMSLFFL42nFrwF75S6g0yczkyrGR4mKtm5/MAjLaULa8F/uZQRmD
EeEE+k61gPQv4+yBaVtY/ui5drlxm8ctAAXh1coV2eBneBKmZ4zqd1NDdaWVnRyB
uPhByHLlosj/RbfxZXUMqW92bciVEbY8DfVYGxodlAK8wsJsOmUSTTrGcNwH+XXm
Sl4R41wwlXO6FOEkkFlKSaAYqafZoHNkYQ9YXUe4pZfegs8NbC1pOuj0sIz/SQ2e
iKSaCoF0gPvWBHGrwYZUBf7B5jtY5p0n5rrja2dIvd21MJ6V0Kng4niw4KMOJGRK
Tz0FQag7H49nZw/ENFL0wFGVFkDzkmEfiY9xhPWGaQtwuu4bFrBarkLRyy5b5K3F
hZjDB3P20gQhIhiIaQqy0tUX/O2UQRylyCPfPcmlna3Zyxi3yxOWoABUFTY1FESv
MVLHtimIjY/3IzsT7qaoFeqRpCxf3zgEnyqkhh2h7sylsnTUsnqDMzwO07Clrcbz
TrCxp/qWefRoCqheQZcFoL1CfLcdStf4PIis8tHt+Z7rVztTGZnMP9A3MnxZQjPe
ern/2KsoxyX68/yVb6valsP3F6kDdPvcRFCJD9Vw81HMRfl5yhiDWUgSgBhgklhf
1X3JiCOxYeAs9NmBjnyYEA4tTpHEueqbZQ86bhaOWquINe+I0YI6197MYWcMWFcI
/NhgFfNWMV+VDnXxO9tGO3LHjNKXQg25QQEGp0eUhl1pHIU9ySMvgAvXWUQnJm76
vgvhuiaerTFpKwIu6Qt7audpHLIVlWzboemqH14s/GDPlSXohLsJuigdvSXba/+m
E80B/1zUMpq1spv5T7BHx2FKWJ1WlV/bKUDYSdB2iv8czKjkjuaae7GO9OCk9Afj
HSzVYrJXVz2mZaWIhlQE4a6drNNQlMTPaKIQaOaLg6f2fPiLaif83r//dvOWu/9b
mbzqa7l3b0j7L2cl7TjKn4iCgQi1HgEgLEYrgXuI5QSklRvpS0tJ2g4GgOwgRBUf
ZdHef7m4UqOS+An0yCEHPoEJt5vjjtfoTn1TWVyTAPcHJXXwmSzobJ399f7PVEcl
TU4scrvglZGuFPxKLta7D7pPQx3WRhwbzK0j+cAm38oJLKVcwiR8Yk6gkfN2gkVE
Vrj/DO6l9Wd/B/+4/pWz3NUSNCpkD/5u1GmTKxcbqXspNmcT2kO42hazqXeXEbjK
9H9W0MRoEZbNcUQsLly+K08ld5b4gkdrZqxa99LDs4JDoIXCBJJRxG4pcqEklCzu
6QUqWB3NKYoO8giUVAZbGPdNEf3j5zdhYwA3XmS/1zNukYakkCgftj443L0wNic6
JKK6rsPO0pLdJKBT4vRIbyTAAFyiI90cKzilZtwA2huF0JVPLKq5IWcuXuPclbPm
hhwj4fxlpkwhjP4tHVUipcYVrYQmxkxoZ3tAcnB7/7iqxHPrhfMXL+T2pROWvb82
lo6LiYVCZ+1ZfAdntWIHF7OU7bOvqhOK4eDhB2t0KooisFR3NEKPtldK/7mY2tjM
Homv68iH0EQn2JSQ2MJlpvk/Z2c2wU8bBGAJmraXO3K1LsiAbP0jZb5bXQh5KETo
xzpSszan2fBnfRQ/OYF5c9atjF9W36c74i5u6Uc+eo79SoP4zPp67Qq8uRtsE3G1
WkzM4P40zn9OCPVHoltduHGvRwkGG55VCCqzTbL3GUsCtuVBlK6wtLbDRgKZhWaj
0ZyF0SgySVtffoyLVp7rUmze8L248NaQh8I4weeAHuZY+QQLVuVzUshPQ01svRQ9
UnfMa5t+s26ZziyRdgecUWhtEcETBvhuAohnbu8MMh+hSZBiUxK2kt+awZ7SXupo
OqOwJr/Qk8jwpqNddeY7pN92bMJu8Ub7QCBHKGmKXQ7EuHa/tHwFmStmpgM8asPt
6EvvsL87rLV4qz/xld+8l4PMdHYb3zpDMdkDXNYoOM0U+JjZ8EPJjBakrZWThl0C
K+7MKagEmHcM4djV1GohugLWO3QdDTGVfa+ZKXO6azZ71vYKTMmb/6jelVLY44Kb
RhSU/wWlB+8E2XmXnoo5sRtaF4YUlPPcYsxYnkuQq4OSFYhCMM0Pk1HVouJqKqUv
sLw/IfTwMxoX0nYAgJKw8qldfbog/SHKKzQUsRlnuYzLKS5SjkLGusaG5AIrjbWH
MmakzNxPRLgGyY00AlZGFCvepEnWJ6X9i3TNhgnQ3kmmxLjsEKXMFgvSiTqLkcoE
/LoQ6XQgwNwtS1p+vl+4BQCWZw9O6CBRwsDV83U4Smk/xUIoD4ugbNKmxB0nL4Bz
vL7wMQeMHZmCi75JvvMPj4QbTwHF10ZrYa8B3nQbB8MzddCF+7Kyg8BPwOSlAza2
8ElSm5h997eLzq8sFC/s+KZwUS0Ujs5Rex7oT1mgK6O/MHFaW7fO6vdjtLkEPm+w
5rOc2z7XvHk/ZDam9g3mn2viyOlErdERDo39rfLLu9LUdf6HHCWE9iXuSnG+MGxf
ubolKaYmWb/DDk3KLy6/CUdPT7znn01E9X/ey7OI8CWoDD0xsKGtJq7pz/ipdXoi
RJ4lOr2VlHSftliu05gllC/tlpKOadQqsj5brut3S6xMXkU84eQivNtHUhe9F06c
x0S4b7kp+beMP6OCkYdnPTQf2wWigdS8d6L8M0XwEA1z307y6jBP1ifYn0RN/jGz
4paWp6JGKO+DvjSu14YwmLs2XiVb3SP41Xr96PXwmIElCdXi6mIJM2cCOg2u/rSw
Qh8doIssYLNRB7SDje303who/F3R4r1dVhgqgWExHVmnAUT8moUnrqdehxGflkFK
QoZY8tP5VFjwaBMijOFfO9i4NQJwxin2JfeVqE+M9AxzlayoZqrNkferNqKno6i9
iexD5ElAgD7ktndYnlLZa64Eti94opOIkCk29Q3TQjCKPRnIJx7P8D9nz1RJXoI9
BYRQr4HAKT1h4pwitWhx6t7xujOyPrjpsNgEYMaQxHUW6fByik1mqsaCvLpyaRYx
0V1/XVPpu14+Qj1xDMBiGiD0byTn66EXAqg8SXBd0sfMRtnuppnciKsIgnrhW91R
awyOUo30pEGaXTW1DYO2qtPiaZiy86rMSwD0k3qlg9vA2oDtf4fWRKkZMALWXNR/
svGOf/PCzhoZgNaPUuuARH80Bnp7ca30WT7RysfYTLeJrdKE+gBo/cTt91zP5Cw8
zFQosg9jmnR7Xudw96dlxLoOOmneG/3cdLEHjAKT6GQ2liQSzdmWTW42FlFk8hOM
+kupwgzKP4rDaam6WaUitAHpOHGRwO4Bkeurbb20sscmrX3Iulo0JwUE0ejLnK8j
WFwhNZ0gZEx8Vvgd6xqkxqNhHkOsePN8CskPT0V4MeJM6Ib2mjyK05xXOZTWp1G0
37FzbVK6Uhh5G49QxQ1cG/PdvDdkzkrBGl6d7m+/4koKzwRK9isu+ImVER22iDn4
SYADwRhqqAx11hvBEesPLs2PIJFKl5377bGvB62gS3WOhHVHBb2QTkf3eb/GN+3u
E+7ueCiUL2Yj7pBxC8yhjQgOZCz3YC5AkTejcNnBQayGR2FhVTsO2aDodpRxkUVu
12vshLypoHMRyvCW4XnIbZ7fmdkyuuKtRr1xI46ofb2j+2lo8FZ+1wNY+wR7gWfn
pUgQPEndzTKxyRqxAsW3PjpxBg8uP1LASgwplcK60lVcVkGvhCQ2+P0xC+SZ1bCp
Twi7TIrSL4Q7fzIXYm/byrAJZSCqT6RwfuCxcAK+g+ehGz/PqSyD1Fwhf2xBp7xh
k6HvKZQdOVRnujiJo95tBqxnVjQaABS38pxBKl2bZxh9fPLlry49IG6W317JWWMh
ZX8j1lg2yfAZsxgsoGWC4YZW0A0xa2IgxLlBXv7r7FnY26+84zbSFCzRHHRrnfTo
M76UYyfu87ncPW09Txr/Hh7K9EtZd2LBlqBKAwGZ1SXYsK8/c2d2tJrJbqgER17i
8PcYEp6/wb+wWySDQGa4KO3dCanpeEudAjfRY4fqdbwh9IJzEXVjeTElUjIhJoZ9
Lbrcm4XpAw3lb6X/tRUYSnbtO2yYnGGJSpPLAHLqNdRgGxOrn6cnih3BMO/WTA78
VYsP2+9iaslGy50PymzFrJ3YiH69mp6+5UeVJkrkW6oSkJ1lMXOsyFT/XFtlwEB2
HmjMSbvTCa6J04BFRUaTjtfO1a58EMNSgHrso8LgJ2OITSPJlR4R1m/P7cVs+zFx
Le47bGwmTPLxENnTMuoIFPCBJJx4Xn+4lDndFkPQ4ryCfA7PHThr5Abd6gwglFPz
QeuNHvxeQfwPWB5US1PG4msuolnxIXOJmbpm51z30vuAWp4qPEGBLYWvAWlEBRgh
EZjQr6sSvmGqSUNtuN9PZAvKEF0kopW2oxdeOFhhoV5QT1q8hEX3I4FiTPqUK4nr
SZvQFH55ZHdIqFBU5M72mZY1XSigPDVLslz/7mdgu9UvjRwaqFbXC4yjj7d8AnC4
AMjPd79kBJZOk8bttHozQjtHcNByVPgIeCWaCCNQt2BZcGotn+3Q8StEI+y21mFl
FNMoigCO+wbrLJABNPSKLrGIuSWyDadjZ3zf8ZuVHNyPEoJrtEiLEcU6kqeUDj8u
ZqcxOjXExPUSCpBAAR18BlaqjRmUMCH5P+5AJDbw4AMeXuEtk0q1gil8+0yH1kZa
/3+EEE6ym6Bku+e58ydUvE7dg6GNGzu2x+hkG0xBH6NLyHkrunR+qDu5ddyLnELO
7AzJ0RsyrCQBQAQeR497auTHM1epNdil2wrGZ880pOI2VfFcBidNKwWr6lB6W4fi
mVpKHGw4sq52XyeNv8U5000V1dJEVcO0b1pIoBPzh+mXPWWs/5V8Pb3js2AHyVmn
KIXO3vluZLygGGcgn1JEchjOGrll6PEAMIveaRDRKr1NuqVAWWB2YLXX7KLF1OIn
pmVbTg+vsc8sPhJHuJKqDaRSabQjxKZx++jyETS5MofHMCRWwik3pmIF2gqzk6Fs
8XAixF/kbISSQQUjWpt1UruvWvOL7cU7mcePNhH2I++RUSUFwhl++sZfMNIQhXNj
DvBSkfDc4/VHGG965lMQVeFFYmZxktm+Jt4Lr0T0B54N2fX45rCvt0YmZoHo8Slj
nLqyVpwHSkgFMa21NrO/7ydTUGqf3kaYmhgDd9cjhj5pQB1hupeJDQvcovDPWfTm
Rv5KDV58qGWRmuRvLCnj+drXX8iVrko6E36KxqFhyVdi5JLsa+/ioxnikjEzGCIE
EmdBf0+zSy8qrEdqLmJzzhw+AGEq+gwSZptiusspCb4cTL9reGUVy0oDRqilrgTr
Ab5nf7MPrrbvztkrm1GkctSpUaDMAFQaZNKFcTaCkOCg6Ykszqz9g4PrKw+jAXwt
6WxxPiDhLXDn6Y9eIR4oX8X8aPb71FowzUrpMQ1qrVHWcvM132ZUl9J1WKwFki+x
Nhm9shnhQBsjJuLppW5O52k4IAQY2/E4iErBLmlLcNx1d+tNunE278OrhvFbQYDx
Z4TFEXe9AUxOjQAiNFx28wQRZDKhNsCpGumuxlnJQzVRxSw0A1sAWE16cAoMHjlP
1tM2HFUVyNIgtXwY0pUIXAOc2pt/+qT/wpK9YdCsEuV9kItbGxp52b82zluIwXHI
fKK8ZeTT2n4cBbIVnQzGmboOJQFg7WV9Oa6TO1ozCl203H2vwF62+sSPyysX5GKX
Ok2ve0RB8Tj6lGfG0BCem2hoiCy3xeg1bsita9va+IqM24NJa+PwcDXtNfhiYlva
Tsxd9rLTTHO+8uoHRgZVf/YjTD1Cn4Gy980o+k+pA+y7el3qCQ2N3blPh4VV90cL
Rnd3jJ3RZc59mmeUvqtsPG0TewO+HWZWV4r2KJDT1kb8Vp7tKS1Kgg4oP3ee+h4V
UIiyoI5AZihEVfpmgHrS9gfkmdB9uhZnmHWYOVT3H74hN55+DA1z5+5RRXnwQwT7
xEuIXY7FrcgScSYHZnPbC4xKgknx4hG7qPvpu4mQ0QHCfl9jueN0krWOTrC6OG+/
Qpm/VzGbCobEkTqmesqlU2Cle0L22yNLYsaqLW4Omqu2C3MUE+FMl82f28Bppdlz
RURKIaqkrPf/EJZtFXaXVWspOD2RNAWQlOjjWlVPUQ04v+si8+C+kwYrv82W5Uss
i3jmO7y6zQNItd5V7h+1FhZu/qxqhNdDUz7oGzLodWMLhNAUzCcvvHHrRxoSkf+H
6/Jt77vy57g6Y6WiPcCZjuhnWcScATP6XiLPw4UkXFFKvq/mqYEQVXz3jsd2Llli
L4+HDEGMKYC2YpLoNiCAe2ROME2uZahb+bQcotM4U/Jid86ogfBGPy84d1wde8ZS
FXTeeqeSHwRhMeqlwgwcM8epxSqNA++10OHUPGmc7117g5c70cbUUbBUqntoHmka
RnraFtSe0B9r4duB+qtSn4faNEr3aqUjwNtBJZSOJaTD9yxy7QFcHLL6UtQ3G4m8
DKSPmkCbWaYFpp+vxlDfUdPrhJmCMFd8i3cxpWGlIR3//MuqtsYYWiIhbsLWwQYf
8BK6nhwh6Avfj60f0EzYMCDz2s3Ve20yJZGZM5lVYrSsWcoaOTJWTWn3CaGKYkHB
iYNhEmEnH5fqnu6AESjAIx2w6VS3vYMctDAFgtO+J1nzd7rgzSwkT2AVOGc8jD1f
mvJ5pcBYBxrtUGH3OAHdTlzAOYKNqgzzshvY2VRq/gg54+7tzI8BLuHQaHhhXbDH
ZgzJlL1DAwq9A9fF085sAEeMex379reGNrMqr/E70rD9E7d/ZDonFQSUWtF5zYr6
UN0YAqxKkCrnjB1BOx+FujPLpJQ0VdDkhdBod0FZl2mAAFQO/fvAeX4gMnAXOhUy
e/FKZ71nURvXHNAJ1GiedQdjKO6cjqs3dB+OJiWOZ8GdgOhCXpI8Ko9oZGFwuNiw
xDBQkGjwBaAznjz7fuL0l9uUAqvYm8j9f8h8DByMvkTL6KJFfUKhHie3RpNsbPLW
LKQi0AFVc9JbeI0HK50yQobSAtqjZ3q40zjiE3TOS2pS8RPNeYrhLSm7S1EVKiBC
LpkX4f0xsvzzgtDSZQsEbAXsLe+v74frKhLdSZyesdb194HKHA8/bPpUKE8FAuSd
V/vN+Pb+SifU2MgZ8nSmVyAdHya0OBe0s8GNbjabRjpvf4snBTkjnZxKcwgJHkLw
bbWK1bCGkdHRuSeqTFnkTT7C6MO3JnUJjMJid0iVcvLBvg/M3Bb80lW508Cmfktx
KHE6ifzN/oA3a11slPP7SHC0k7T5yf+WN+vtoGJ7F4rDCaxVnFkCq1e/C38Tgx4x
cmNbkhorRa82a2HSenDNexnB35++CgjXIDBXYVfn6OzJnmI1lxYTrqDQHrBVBSN/
oOLhAhTC9TBfeasgvsDTMhv0+RMFjvEtMyVCjIDPU3vPFFUSXaW86OtKVVSjI2HL
Fo+h5u8cudDsFcMA0we7fd6IPrN8Qsa7Dz2ztPaERhamfv85cq2HWgVfIKqjclYw
vVqZAxruyDFp9naOpeKy1VtRzaOpufa6UBRzg2wUf2iGyLkeeqTSfO5170MqGCsO
VCtc+w5IllfaV0Hy0DaBuOQP0djsZKPAzYOTv4+roFFsqICMtNoDY1DCzVPYUsoh
EffCL0zdYoeCzsllI0UiFk9i6SBGZAf0H2KCSaCi32zyiBshqXDfgRuvnGDvMXFL
liX7s7EdQOIi+uVnUBMQrt0x3Kr2bm7xPoZpRz7B6J5WK7d5ovqP9ivZVV5hpTD6
v4YyY8ZlBHs1DoQ3tk/jLsPz0CsVYXFFttrb/cFWlGFkdy7jVYaB0o+NXaHgo1lN
S5hIRoghsIBbRCpy5rM3rrxhtMWfAdSeLC00dAl1yf9V2ju1c6cUEtRB9N4rLZlM
nvtFPppkC5u+NnEBLILHpjqwkUEe44M9s+capZpOPFIWYukoy4KMfCrotWgBeonx
7xOFCYDTn5AnVKym9CCbyX7fJElVnmoN8dKmVgXukbWt/9sJXN1fuJDkXJCtj57w
hMUXxPIVwttwGOvZXGCNswUmIumv8D3IbTbb7hqMozdxBMBKgtvwpfOXTWRDFGVL
q1iJxKFg3iAXhN5MAWsON0fR3Mplj0qPbteZyIsIfu20WQpR+sFwRUa+7D4+1PwO
aXDXYP981FNAXKwv8ZtvMHzbxCNfrURUV1LR9RTn6EFTG1EjG+0IiNjo+PLrawga
tYnPc5/ecVeD/RKKATYT9GFsiHKJu3ZvwGIs5NlMLhFrN1aXr5BDEcGOiRzGppU3
iYEgjDk205sEfVbOI0GJbYEksIBHwOf0O27UWFGO8vDonsL578z/VZsl9Lp50e5J
OXaP0HRUBy3spLL+vuCDfGtmP/6lPLGJucxDrqwVFx+z9bvOKu52Gp/fjxv+MQVs
lGCCNhN/fHR9OC3dNMjSa9odm7Tg/h7aeIhLqOS/nWTwq7lwLqgsxzFYspFX0DWV
8o0KchrnJ9Akn4Fr8YXTtBcjFPo4XSFNq0qDtL0S8mx5vGq1lh4+BlHq7cQKhjjP
VODv23bs53E6wOtUvcBF51JPuTbPtp/GJ5OiAyb0uDdGCEj6Ppx/fYt8MsnGXgi8
ER/EBF7vybMzb9FCGImmoXj0xJ7h6nj5i4BzgitnOefMIKKPe9dgTUTokPgciYMp
1+LAtDeFd9p6d1GIRg6xCnYxu10ebjYHLwTyzU+gk2r8GJv8oVQHAfHYm6S9PNie
5+RPwCiPJVh3sN9nb2RIRe7XLzGC8FTHo9ulM33Z8JHaPcsaaSj3WQ3RxumKaBI7
jRNDcyhYLypFUEmkff5TmAYYGD8uiGq1sjMenM72jDDzfwnpWMmMJppqv9yshF3y
rfnM4hcAa2GIAO5PvD0VTg0e1xzNRNxWOsviyDPfyhRiFL9Ll9KLcpaPfuHQm5OK
pBmOl6M794v5tOSyhjAn3N/TqryW2zs+sk4+GQOrREUzXkc+t7wHHF2vEuyPgTIm
QOhVp/SIr0KOa7NduVEcJivEHlTfx8/B655xJRu5wNUGibf/j++ofukWg9y8ktpg
9glC3Nke+tEIePzWBPFjm3oNnxFUiVnoKl6dLnfFLvEvV+GSxSg90dRDSCBlatII
3OeTnvscVloyAK1fDb7nXClW/fEK4kcuS02RJzxrRqypII7mG0p5OMdabLInXwxO
j96Si+vwP+GXNWvDK7zaJhL3v0VE2FFQln2WtiRc6JIh4znH8gExqNoaSzkVDsjQ
g/il4ZRmKJKFFcWpcfn1HgoTYI+YMLo6oGL2aG3FU05jOm2Z3EuP9XDCy73LtJ7g
ADf60f+d0+Z/huFz1/cdqvhg8rXi64iyAhUZgL7SmozJokeHo4Ilf4LClC6oZZnW
n8a2bXU8dUhioLlkGVUXWyKhtzDNOMERZR0Dlmop7yjwd4xX/A3J5cJE5MDVN3za
2tZlFFqN5z6NcAaR1z+K91mq9tR9omNQHiMsgN+4OVmm5KMEDB4TZEJg6Ex539Lu
7zLhBs1hYHABiUdg8ImhIxWlIgFjI2ME1Y6lvkLQWwO6OCL2ezYGYw5Wn+Yogc8o
6x8RMNFw/WOtGlvQZ2jSxZK6RTHhB/3qEJnWqOkh3lS/f6qu1JF7jGNR6qGLM8YI
PfqLCaoZ9pPOHCziPDk5Gg6pP5vc+w85RyE1zyT8j6PcTRE1X+WWCaHzniFG4Jzu
pJcIsHT7OtzxYdEmm84Jvt+9eRdfPz2lSU23uclZgyEHtJjDn28xl8l9/Xlixlq9
4DXPrBiE5aUMoQ/z/NhXEeqQemat3Juoh91hjCTm1T3utoCU1u8rk+XdiNsne3Eg
AElTUL9pjT99/eif/QFuhArTFZurdn+PP/QV5s0RjdqT29Viz3sZxR5qSmnJdlBb
j5j1hzH3iT0KqRurn3DlnEJcQRbmewrIb9mR6XDmAf5ZBnQ1s8C4gNpj3alfe/Qr
jDip7r/NO+8P3O/EWiaqbYNKIlgijSOkwFHiNIyUs8FWum9D/w99e8+4bbim0KMe
9JH44GW6zkMJFqz9lSx4FaYcvNRPqIk1pHCponAyohtHCTz/tZPEa7h8xiqy67iI
NeUu1aWAV3+735RJ5DL4D4n7rb5hibT8WVCCq4XjtESNQ6RclAzGOAPDXRniE7Kq
YYZ3cyaDSQ5oeR0dkTGN8RzKYnU0O/XeuTv7Y3xD2fMpcNgrZzYjh9ryA9XvlTVG
IA0JA4FSq0TTCBxb4omSG6rAq+ccm2mE5TA6JVESTAwvRA1edNSKlzVf650TdhSW
+H6gyqIB3txZCJT35bzYWkl7WJ6uHQcMocOM3G+B+fzrJgI64VASF/3haH/5wBJk
2zOYxE7rhga5UvtrDpU4laGiR3p1u+k2CkmqnbnhTtiB01RRJ4ITo5mSIJQg6WZL
xEcCDK2es7Bw+FrIXDz/PcVST4ynEe0c8MPTpw2mYEvEJsEUyy+5e1baeKhVuUDg
BJ1esI8TqJE8wF6ymfFgNnMrJTWDnCFLIR5pTsiW+opjLHvaTkUsOSAXySfRvAlh
ppDFkQTmkZvWI8IV5Azi9OyvQs6K0AJZF5RjAuxCZWFxNtVACf5PGtO9k8HqUfHh
a1MwEC571/KnO0XMegwpNOppg0lmu3Kreyr777p4KXhmnj04/KoA2swesn0HV1uN
dilJ/h87txnq0Oq+KIZP09v9UiYaz+5AuHT7xwITNLf16WjTgSATV3LAKaBkQDhi
V1/B0vNnapl+oUkJkP9b8VsxOUu8sYF0xlb9K6354tZGojrGD5+5fWRcOg4EsQpU
tXWyGVyTKiW8bMEGHesALYzVC4+rRKaMbscihX/KTV30OQBERpOj+YfI8R/Nzh4w
SS9PKdJ2GzUGYEDT+aQW/DyydFoMUL1TT/hdpT6HQSDFjGVkCd0vWZDW61lzaICy
zhvGJeXsTC2aO1SBzGw8hvffXUFo+3Lt1SRjbfCxC3crhlbP1WrQOs4Z6NaKijKf
hyzH4xdB+f4dq//c5lO7LbuOCQb7cqqYTh3XH9xysyxEGPbLK+9wq0VEoqr7uYI5
3yLO6Y2PgrKYNfNUivUARR8hjMTBtvFeTPxcj0V6dkzppMJJcBGfrnvik4j6S7k0
cWrsE/R5FNPSiNnyLREXuS5pb6sWpASI519gpAYOlZHI68bNpmIt7/T/Zt1LepMz
2CDt/5aITJpoc3g6fM4UnqrdFeYwktZH8pCv5QjQu3Xqm/4JPvGY7rVyvOByDum+
AFg0Gbp5V/zE7TiOZph2bGCPGFobeQ0ycH2ykzQD0a26Ai35duiTgHdwocIJCikE
XW8Ttt6z9ZrKXus7+S3N5LT5iWNRpSZyPQHyQx+j/n/oLtieAuJbPZn0giwZYSrv
GuJjU7usguy6nK1NXkadg8mtPyNiikgHabvmYyN5lRl6kPvj4RfQJGXobjZ+IaMA
WN9KEIH/FNkgObVK/qrDsg4y+my/uOxk6YLFh1RiO2MrFrs9MLYtmhz3YYyTw05I
vApwC04PGPqFVEPdkb5aLRVTChrCMq7vX4jg2Z5G9iAcWGpgmMVWcR55hHBSxvDA
w2GXyw6IMSHWrXKmKt35U+iZ8HfkzOHJZiBeowFrWEIl1p6OuWgky9ILB2bPUth3
1hfSww2xmMG7PjkCAkKIJKfLYjv8NaXLwIhBiSfoTgtZMSJlJdOGeeFvKlR/IqIy
vlHr3QCJQcsXZ7FTCjiywq8Q4W9BovRhcfZfIoWqHlttyz8QptuO9Vc2JLyxAzdb
EpzU+h6a3X5MGW8ohJrUoN35hwab+BLknPpDagbvaT8RJuWExtcli0fMNSfjPshn
wET5rmP3pXwQAoWARnhvsjOn9bO6OqtO9C6fbHdfdis8Z4RIif7DKVVpCF6yJI2c
Lh8wrOc8zaRzfM4yV2CCvS/MLfKYSQLrl/pFTQxJavi7x35xTAz5LKYnH45pwqnp
l2k7P/tnLWgUCXjwlkczBsyt9c+BtqW2NwoSSLf04tw2ivIv5FpGUpXAzToHxGkx
JtZ5yXObcOFkeIrRly2cgIUwEUYez4TvZKzHpciFqSaQHbSupPR0yM0Ump1wBwgf
RVr64h5BDr79cQWQPt6Y0Asz9+oEHWFzFp/rMk1xLusEFnOnE4FSCWzp1IMWGffX
GlWZB4NxtHiieqQuDywa7+MFVBowfGtcGwQadPO8l3CsH1cxOGfheY4SWPRJmi5l
gR7vPosOFKB4Lk2ckCgTYThrux/kSq19tpiZqUd7QlVMMciCNOtYKDK/zbhszzP9
BxdwmEASgT7u46uLiHYFVwRzcA/B9XcwqxsCrDOV28jQ4sS/M84WSAXeZet4OEP4
PyaQAlHwS7hu5vSNANUVFGAGjGNsvh3jwORBE8Gbgm4yF2TJwxRq+M5VRIGMLUTN
K/x1FYMYLzifF49uthosuhWUBGaLC5X2TItODDiTZbhFyXtEr+7JGSXB/IVVgzKq
3kUXlyfZPkPV5WvqiToKP8eQrTT7ICv+HpCcx6H5A/bOVjYaJyIJN6u4X1tp0HKV
II5Rp6oGg7/I/raHU/0n59V4C6FikNoWS557lRyDSUsFZwPOIPd+Ziwheh2QfOTp
onIumDhDkzcQ0oDUS4yBPRQyDkciHM+ZEgWhkOgf1mbWCVtPZNRkdIuBdvPqcqMI
h8/iHuUE8/pGAN7EpxTWIuzlf2a502BD+HxYeeWeKuqvrsJYjtw35bCSpsZdCAHO
OxaNvW9BQuWLsH7qN3QFk7qJkOhqRwbonRm7yYItsKmGLECdR9I/MChJ1q4FQAwR
lVJH92RRI2dGhe+5eNtI7s+EpXVj+QvovxBNmf+svF3BPmgFtiQzH3Ru9lWghsIp
cZwwbKmun+uVqZSsuH7hB8eRvTDvJrTDv9M3UXB4SGlhaW7EhH7GU17mFwQGflS0
7RxuVhQNFxmiWWVGkAO6Xm7I9xLpmerxle1cn6aD+AIFGtBDSrqIU85XVHe+OKGE
sSHkloSFeu9VaIor59W4ZkbVk0j2iAQUtK3WYmQzblcVuF+Zc2XYHJNp5KFxuI4U
DItBxeA0DyGR6vQxXVON4XlAZqOC45G7sbpR0E+BPaNdmurShGJnWNIyN7/k1X+e
kIPZQLSJeK331YkL0SIvoMjFg/nSx1Qz02QW6WmmJWna5xLHUGSd2jh8KZeXRBzA
DL6wtIZel2asP64ZFZSdp/msv/LYuLiJvcers8LlM9TZWCu09f/dtOBms9V+8Mob
DmbjMjCIigAzJfymPwa8H2OrsGyGgO9EHHq/L6z3DwZciknMSV+Dls3pwq7Sw2aC
SYf3F3TFo5BBit2rHGWUTsKP2i9teyMdcwbjDEYWFVKaZIpOP3/21tLfX5bQ+p61
vWykd6TQ7JaeQRsmhlptQzbHAH6FlACUWb/LQoTKtuh20+n893q/9moaKguZmJSx
GOk1ZgEkQdnGysKpw4ZYpM+LHCDCdoccKvC5/nIPW+tf4PZzfvDacB2xONN22jRQ
yVAtdeZchTe5zgRAU/Io4yGh0z5OY1T/ZO/lHXMEqNYH/BPDj+zJTxDYOyKRG93X
UnFtvaTIhd/BK30K9FCyLIbviRvlyQ/+xVANaSaImvFrDcK0EQgAEr+yzvNJJl/Q
4xQYzfSyLvkcWNbGsOY7hsZtEv0vNCkOk9FLBXQb0uozBaMFVG5om+FvVh0N1CpF
IRjpXZHoiEtonL+TPtyxT1Y2g2XYKdNtqwhiixwz/qu7Vd1MUl9sk3q/dxT3Rsq9
bxMmAVtoV6iyWhqsKzSNu3eEskbK8LRV7f5L6hZjInf28vG9rYc/qG5NsH6+0Pov
rzP5dG87LbfGfo3qkdVaVsWCl54NaDZ015qWQPwmD2qYGiALx1lVzS6lOPFy7soK
lqWqpjXvleXA+XXbfD6oza+Iw0JraY2oJ/EPy6h8i+StHRvLfew9pt9dFaxP9p97
Ktv+b3f6UfTypE2YUq0in2PVSWxPljpl6D8aX67KFYgiUnlGwJKCDsC35DtVCXJ5
/5VZ8+GhwUtXKTXnF6OQ5yc4nN2Wgn0B0+/gNSNpocBVI5Hv+Mq8iw/9wKt7qb+6
9N2ok2vhPTZvk+l8mzSDXjavlpRYoEqX3Bd3XUdiPvVJP0KxIBoki148vdG3l4v9
roNeUUoJqurrV/dhjLpsFQkFP2wiQC3hbCNL0vznuekRjfPhG8YLdx3XrHgnH6T+
pXgncWF19vJ8NjAxaZVXISfqMBsW6C6eJkBCeuXnZioR1EOGI43FirRAetXmvhF0
ndM4Vn8xQbkHo6B9iHIDzeXU+NRe9vBfTMwpx2dMTc11Usb4X72wvVq0z60ECJWc
B+TUW7JJ2wrBea5wtH3pl+HVaoOkEfiiDtkiNeivHFC1+zzT0j9aKMtH+Te1L0O1
xz++2ap+lKRV8yNJSFf6+5AH7ZRlDVPudOnPrhOrgaSWCtv8+GuPmAuoGARW4D18
pEgpS7h+AmGLMLPcPvzX6iONPZnzdko3ihwyJWKioWcH6+CrUEEy9m6JVS6n1LaL
qySOKFY4iuWHGd/LY496GTdU+AoYu23pdponvMMq7dr4SVLGyB8TQ+TrqQNyrtMu
/HcWeOnEGXXwoHbk8D68+eHdmkeeRGdmxiqS/wFpntDYaTBqWUFR6iz+uaNAc8Uo
1f9YJ09vdp3znpbg6usS1R7LsQtAfp2r3hcQ69gGUH1Yv74Vp1nI7M4o3NYnx7cx
xFAEZD00IptdjuWfg71X2zD74S7YDFMv1+Lw2bToqzy0HBBmRadimBtUa4O/M7nq
f73XV66Qp8CIDWDclaWXGuEMk+5YcmAqfDI+20cOSiwv5ZwFGuMRUd+04YDfrz4a
woMYLxW1Jmi1x6WLMbFe1mph3WI141aZmlUkWb0d2sXAF8DiwTDdTUNMePL59Mxp
0tTEhHZNiPLdQ7sFj7eAv5cPdDviaotNac7JPWEUxoLP6soNBunc9jxt37ZVKCKm
nJH5aIjnJ3C/qBby4I0focHOEFo0t2A8zpIf8m9HOKb5fDnLiYbgsopnnSQvJdD6
KwERPu8zt0toFhsGAxeVe9qTVaDqEHh7aFS633+9ut9ydY0G+cc1cJPT3VQEVjby
FS5FCSXvZEscbsh9VQESB+5P7iqUrRQF1FlNyfwwXJimBp+HrSIGGnF24L0D19gZ
I+EwlpZZsoN1W35riJkJ/ttLOW6j9jBHWz0Hg625O9pWQIIp0kWFhjECmjMJG8yL
S+y6ZO2dJuCVswZ9E2AktdgNDi8UbJHZ8KTfwQLcCTKKzryCBeLKN54pbhuSE0cZ
XDR/s8+8OlAwaM4S9mVQ+BjDDwnNHa9yDPVefCN/RkgaFuWGGWeYzujRo3A/IniU
Ig4y6/Tk57eYcE8OxJOdOad5RIiiGYlsOiXG3E8U5XUKX4dpu7eaVkN0QzKvEHCo
wpseu2fAAMKAT/aVMn/Qb4dqb19qc/uTZXbrtLfmX8DhKfe9gItJfzMpQQa8rTXi
0CXYnl05zNGAY2k65c48TKKyDxEJo0DmuWoY+TZdVvPgl1qf4YKCMtymc2kHWVyJ
763GuA/kY7NT6qvaRdijLipZFiXHKPEmHVcTlHy0S9dSGjBVD8pJ+w1R3oMNKxYU
yVhuULi8NS4jInp78KUt0/nnnUoPLUoiselvRPG0XsLuKdHVlWOR2Zaq4NTaZmbF
0dVHDsIkE8q5C8Tlhk+UZdgEYCADW64m6tN9OZK7dYOlrvJODhyUB9ULgsCBNd0N
lT+7ZOfDkSfWiijZRKQvsUSrdmFM1JCNBpDOsq0V0kTe9CoGaW3dpoqaHVJMWfs4
Ywy7wYHWjkXunUEpKsYyG6vHBDCJ7nuV+u6bfxiTno4O/jlkn5SN21RvA4prUx+J
5OoUGG3ZFFxza2AzWoX11XK5tcNqR9b8XJtoFwHrrBtdIt4noLmD3vR9WVypSQA1
LPy7Yn9cQg2i2Ci8Vr0hktj3m4rS3z1l1YeqPShAIDTjxopb6bt8umKZ008Yc9jb
moba4rKQjcOigMvJuO0YWRLC4wg3boFlq4ZA0Y+wvFRiivtn10fA/pJfz1/QQIG4
8O3aRckkJfHW9MuCFY+QSlXZHPo/hGAluI8OVdOY5J4wkp2jdLGgNuENsm37oP19
hYHYzdMIipccaYEKQTp/O22GGFPTNFtL3DPhgnEOO2T7Yn+Yz1PZlsaDw1tuUFCT
QkwjKAFK0ZQkkv3Kv2eGiCr9QwJSi1Gp8VSPo/LXQTwO6KRsFV7uiV/IMtPfIMVS
+3bjrWXdfdW+KQ6ZkMTHW88FnhxPJMc62boa+vZKTDaSNVDFIo2AoAQWftOD68bi
50uPR99I1qBqJnQGsnnyJlb0tmG49jdZKPC41hbtvoFMq50IRdcpwa26T0FNFkbH
8DBIM6sLPJRYf2nOFiBtXwDrbWqU3RQUHxySmdW+ta3F6AFPrpAdbovdQCrrSE8D
mhhoiwuE9TryXwKf6ojE3cbM8KKa0krhkDsl99IUrYT/4ZHjkRwj09vItnjHuGn2
wuUibG4Y7cshrXlqvFvSPnBO8qpU2jdj8Nh9dJMX7UEvEbE4JU6Y5cCinwxsaiRa
WwwwP2wTl2hF+VY3GZiWpWF0YhRoyaiCrm+Q+X6PAf6EUrXWp1qYoL/rIoNOJSgc
MTcLeo49uaQsOqxiwMHSdnbbx31YsGeCvcclev7C7mh1fEHu6P/IDiPCN+4YhRWF
/7WDCN1HcdSDycsaLSXC9d76Mdkg0q8/QqfENNqjmeCUTZZFCumHNFutGgrWEVFj
D5L66F5OLFpoNecwR2niBzJ/AOhTKdj0l7SrXEWIKkbSYtkbT5SL9sngKxnEs8Iu
np+ANShucYS5YB3/m+wp8nOoREu9lSCIGirhvy7HRG3fMZTBles9/d02+iG+xqCg
1pfHGBIZNeQV/jP1VfYpY/Hk9rUaOYmGgzA2KWl2/xfYZqDte3a+DE/MYgo6qzVp
eOl3NPpc8o9wjpWbSm3V+Zam00am/59xiwn9eRsIT1NHwYe60KcMiRzdqU6OQA1A
9UhvlRWX5X4+WkcYYgXLat5V6ZxrvBCClEYgh/P4hHVMSh5E5yvg/Amo7UsCRlai
70C+YV9Te3eIp78SMnNPAXaEDsIpmYxMId/iFT5ZkG6EbYl2loFvTex+D2pQUCIp
VgV4vqkykRii8bXUk3nes7C5P+ECUigxkccx6tyue8dAZO38dXMXN/TL7k74QtlB
eUidvWUzF92bihoS5FR+UTy1E2VVpshdFJ9bnLXBpQaL+udwK1JA4i+B/t9Xu8q6
51zk0/tpQFZ2paAQ+1pbbyPBdRxQfAJ04pr4rjqM2OrsC7WtiBCZqCctzapG6CYa
9CTg1W1St0/ucswGyU/40X31FjciweE8kVr7MB1We8SygtAJY/uj3yHZVJ70Q2Tv
kSNqVkm15Qa0SQWgOxAfue3jhKaxams8AwkZVmHxc+bO1PXp7fCdAl05RmG/9c7H
4v0EsFDwFOXnzxXaQ2V8PpSwTZUqYZxCfZ3SfBXYeBvPXffH3wxrrGpFMrGitTeL
A1Mhu9U7OWidTShim8qr70Hg3ez/8Cgz5kuEA97n1OFzyTkGCt+icV0lyaZDeoqc
42yIS9OTS/PdQpGgLrRKSCsd/nzNlhC5Hc/JtBlEZMG13oVdcrnUj4Fev0AHLgVB
egB7v+tATmhCUWVR659oXdCb1GUm3X7D26LRlXYUhRRO+69gA6I3DO0dDxQ7D8ul
NhIO/TtnqWyLCvkjlO/7jRsgqKV+1gsJuAs2N3jWokIck6HD8UH0mpseBvmpkSVM
YX/FMf9yBvRt+q+A9H76JsO65rpCUQBkzTWDauUCDpWb9A0eewH4QVeo9v7/NpRN
EN4lKHyQR4MwU51RA4wM95HALWW3CiEtYmFQ0Mp0wKjwxKqOwODeP794BiSa9eHD
3Lik7fLOSyQr0QqZ+vMOfakTjlNNfqM6KVWPnos6Q3x0f1To528CSd4Aygn2iwqn
4z4WnENog9GV0x3lcE/ZfhD71TsPnfWsK01fSDlp0pDuQPPlJYNagADVKilZkJnx
H4cuKbAh7jzgh2vP3lxtPU+aUyxPIeI/77fMRXBAYc6amaMeXN4zhoEMRFUfSPla
rctyPp4VUiDnyPsWV0bzuZRUcx/oZE0g+zN+WLMry7WgFYX+ZAoLrftEq+2WYU3O
2iD8hmJDh8p8uYCkOGXUPgsiF15vONmFMefV9dZ71pj/s0iMdYRU/Fu1u8RQ/4UQ
61ZrbtOkECoWbeH7+eua5qTxiX1+MLaxRHnSHIAewjMlYX5xYEoRGh/pr1Yh2iDG
jNU9EzDGp149zQtlHheeJPxzpb5tT4iJzbkBfSPlEJNGzdvDRkew673jU3+kVoTu
pFBM+4aPtOPNeZTpc9NtVqL7oq5QHb7ygnXeN9h1NoGNs0TkN4z9WWCQRTd1DYME
O0rCirSyYOtwW4cweLiWj1yap88c6+pkbCkhJ025MpNk2IrVn1fYoTxPHy2bU1bS
aH1TzHxquay/7lpkzDWW2jtAugBYobu6GlqtADB74KkS4FBbmSHjmSdHwlVyrsd7
Kao6nS9tBUXSWDF2wJmQ3jnH/iKPaD+CGnU7ofgSeklBr8Yhn6KeAfBXi6EKrGKZ
ARKqod6IU+/YAsIvYecUWEh/vpkgrgQB5qywnN1hyvOoMkYK+PChSrUtLTwFNOca
x25cTfT5RjstaTTgOqZlz/kXfkC4yQhobgx/Xt5aM5QfduispjyBixLqyxhVYnGL
eOig553OqJxtD5s2zmzdBjySFwfwFZGbFLXkI2DmFoZaSiALZU3zaHx3VCs7o7Eb
gHFi9nKXmdtlPw/fgsHLRbMVUow57ECuRVqsKWPrBpvVMsNvS0Fpto4270ZColfI
mZvBlI4fG9F3fdx8D2KcXI1mpbNhlcc3MCghJ5mLtZyQGR6VQlPt1MGGDr/TY8Lp
8DzIp4zSBFqcjTyRqc3lRTJw4fH/wbErHxiqwK1lrRSxQCzwxLkOUGS/dcOHt5bl
S/zaO2gXnzuzJCQv4f/4mAY2IRdknWnGqobmYMQrMgX7/WGKW6XzOGKI2kD6spuJ
g9nkJ2VYQ3RdxHWp4YCwFCKOT61ZlOY8oMA5d5Z4/amxI/x26YSD1AxLHUYJCjvH
WhebYaMM/WunFlhhF7BCRZ3ZY+Bm2JDIO6ob/wWVSxv25mb2YqECWdN4uM/EsG/F
TPuGbnuaSNvvnTB7m73wqRzX5YtNqWh7QZ4UjT+Ng3g19a6/ViZvT0+bAQkI4Wgu
EWghqlvmtreLX+wWWcZrnu2a+1ttd+YOCEohdcA8+eHYo7Xeg4G780Sce7qSj0Oi
3fL5nLxz/jDJ+eTYc6ZE5alB7t3C1Ugozgasoi/UnjeMU7hPuNhf6zmQCpmIeOa5
bWGKgGjhO5TT59os34Ipqra5YgYYFWlSGSk2CbTqu5mg1dGhqQwk5Qi2O/Esw0dt
Ef9mlcSrSVfgMbbc4/SAhnSYTP0V5RfDmpskya/jW4hGX9EIUvgIztrYkaohLye/
ph8FXu1SwQfNj/i4DA/mpT8tx5Z+sllhdee0UHkVdw/MjnDXZWrTWXvP8NBkQpD7
48W62FLTCaWcO0IOdchyiNAMEoLG65feBG6b6IAhnatm+Uh+f4VNzLnTV4Mc0/KN
8qwdFwuI6PcdC8M0kmtPBn0jMewSEv9d6w+g7fp5qgAnA1JKt8f6Bt2UFv5OlgEe
kgnpWZL7XwEFM4tJb80ezGf1nD9dZBktOf5o1G8WyIgqB1VY9c3uobEalNWqbs3O
eZBIsznvgIOtdSVfxxrWnaAS3RJQbJhkvKgJRg2WTC84FvPR2k5on8okzYVWFew9
PV3OOHdZCxLmttAkEZec5ZqPLr3L4RKzqQqvU96XILlD+9T6GAWYo2Cs3OSkwvzv
L9xVVw7NpSLNtrrtAj470Sw9ffXZxErlMu1GhcXq/P1M7sXRHIxP7/OFTJG2eFo3
Q08YgWScJgwQ/1lzvkUbSTbp+2DzXAOMlCpell7vDW9gscI+jM2jEo6hDutu+zb4
p2v2zNoiMN35Q0uu0fY4TMeQ6j1QEBXp49q5hwBFH0Ai2nrl17N+oDr+OFiZfG4a
2i+ZWpisBfWimdOcgVe9TXLVvnWmqY6Os5dDLM30zQh9/s2iFMTH50WOd0M1Ksxe
3l6yGGx6E1O1IPaE2gIcMa7FE99IzswKt4xj+guywZpZGIOduz4zk6tbw18H2WXM
PDvzNejvD7E4aqHV10loSJ9IGvIA6PlfbGYhtkoFIGTXsjJZxSvZLeJ4Fvyel4yO
45KOi4rMHNon4KymxLtEJ1xpbcCn8i59AhllmjNDGFT9A0wW4binfTtMPityR02U
QWnIHHMS8tTNaf4XCBFrsB2lxv449GjU0+Yohz4WVP51KPHGLN1olTV6IrQh7dlh
h0TYC8j6Sh/0kMs6COoQqMJmUsNHb8FkX4DQGwDUqmd9pQcECl+a9uh4d4KW/9PY
b1rwF2wWLNb6Sbv4Q6vnQe7TJMIL9DTP4hWiHfDUAyJoNr2y0lENcIMU8EOOh2MS
+cwUDNycoCOaLqRXCdVs9P+QWYHc+8t+bVuUgEKO1N3tiPbYdWkMOz24KRSsVumQ
drZviSknX42g5kbWrrDlJkg+7dh405SwsJzSBC32A04HhR3suRI1vVdltva6QQVR
TxjViS7tqKmEOscrsOF3y8mBmMvZJaf0LUwIYbABbIxPFW243m7xyFxlucrx9XRz
dVA3vsd+CK1fztp6+hGHG80euqVOgaIFPK0XiN9VLWHt8Km4baGd7vMKs94hOgDD
oJus22eWyfudeT5mz8iSEnK+rl6OtaYYziJbojRgP+FpVXFmFyrREkVnJrS3FEp2
Jnk4K1mNsBMaUc6uoIMw7Ru6gZ/Qcf7hPd4b/DatO3kLiqILQ2aq3jjTqSoVIB7b
aWgAup0NKpYhjlMlRwjMN33ta1C38NAITLy1M3MlaWTnyZ8p5JvpeRqiZbt0QsNe
xTKclPrW8bXMQfhCNWFqNQlRa9Eqz50tMAlfGoMmc6oXWUdIL9COSZv2iRl3F0Ou
z/cOmTwHph7gJSCm6gIO/STAV24A7gRKLaAuSlw4iqK3ymoxCnfSqVrQrTtsMtY0
5VTmQfLRT7q2Q50vDMqh2QN1WV1sgLyNzNxuuqn0qx845E0kMAcmBbmXrg0n4jmX
jqY3leJJEsz8uN1fLJvBRBLWgLdJ7a619B6AiKoseDfx6NJho+phxUpm8hxJd9z1
B7U7G5WMrXm+Lw8sT0cmT/xbhkkORwd4UsVEeOv0BL46Hrq6tYq7SdS8zymlPd0Z
GoT3TfETy1NBOZlrt84q/Uz47OQYjlxQeDyyW4TVwJlH4c6ZC6dWrA/UTGkKAwQ1
Obgg4flewTKHbNGqjufupVvftE87HjcDlYIysnhXkbyex/dOwMitWG7iIte0Zgc/
gFYoNWJYQwWka+C/1iJAvveSXDh0oBeQTN8a6+DYM6KCT92iiPTwOvvkzKi3dXJx
yadYjj7ho59HBrNQb41uosShVy1N7FWDlb52EQKDsJXvlII+upHxjuVjiXB4gD4b
McoE+ksrVE2RtrhCWQu7ZcZiAj8JILOFgILU98Z8HF4MN+ILPsMVp9bxG+iGpRQR
VR1yNpjIoiNm1S/t/IVyRM7XbkiMp2ec4tQLVcwWgx7wjsG3ztvz896AARWisCIc
AZ5EvwFy49XyYyNw3DtWGiTZWi0zxYA7r3GemcVd2Bf6zWLJEwKoI5ljknFl7BXY
2DtD5WE/N14YS+nP5tdSy0/DYIbyXvxrkVZA6tJoGEVchsMHZzJopby9ryr36g6f
zvNaNgF/sb+WxdQ5gYld3AcRu+3ari9/ItfVIqV4PimaORm6gUvzs3ptpESCIKNI
nGyEV/a1CWWztho/KOFmQayFBthAd2XEAGVPM3a3U7+8QsAr86Uqlyx/WIDbev+h
FEPF9OJgweF9prF73BJWgShA1beNF/2aoMdQwwKGpPF6+z2c7O+quNM7d08SPBAT
Hx5arPoUGFB0tw3MuL7yp68uLURug/CM7FlilAj4W1fAP+lBn19zI0FO5GpS4Wgu
Zj5Mn8/EVD3fYiAsezbiTHZgRvDO6jFNGIVF1kBfjHw9BRQdMlWSVcGneT7wd1xD
7iDHj0b1LADDh+SQgU8voYeB6Tp8nC26vhE084j70iuQwh2Tz0zSskZcjCtwl4IU
ufvVAgdbcBq1uDG2WwcucLqD8vVfkjo9/ytrzqXRkFEiy1C3w+k9XJXZ/0PueYWl
j0lo8UYvQ03/DhTJJ0Gltxt0hqj0md9eLNH7UapprM4LFPbBC35uU0DbY7W9v2P7
70tyYA97vylu/RPlCeYOKxaQpySqxJNUa8TgssqevMggPQU7z7sqRci+DfqcZM6i
3KpVHHLZmGqeghVldO4SSaicBRwFpHFx6C9z76KV2oD6EhEMyVeBaMNa/xZtzk4W
N8YIwGxn68USMSu/OBnvYyE7tzviNkwD6B9p4mwK49dDula2/kJcNJ9tanhgoWj2
514PKVV5yRvnVhVYjshI0jjbhpFQ9VT6XQM0wZBTfIUTdie2LAO25bSlJu/OjRgP
c3IrfwCMGZobQmkllrriu3TqQpP3xnqkaBBc/TnJDZMhQP8ttRvyj/t9Iwbv0FdI
hgncTg6sOdfJOLkrggExhMX0FN3i3m4sIvrvb0O/7ankhAgbi+uvBdv1e5sejdK+
J5+QQg2iMRGtqOAfz9vwX/dugcsueT/vOI/b0eSjjRAw3fy+GDNng0vn8tvfid/a
rIv96LOuXJw5/ZINMnunIaCNHbt6ZznQIYOEVQTo3hWZE1S7RMXMkjeGMfQue5Z9
f2sDayqqM2OjcEApPd8E+HmpjDTq0UgaLIjDNxnK4oujkQ/St6K5SsKQzOnZf1yx
whuCoZfGK0wju3gqyQ+rQv8aRmKgQie2uep9nhk9lbBxII4EcSmKNmytF3bSSF4S
S72JaPY7S1mhgmMfaWeis479tmdrDjELmCu1YKdxVapK2+pMmTM49CHH/4N41jw/
7JlFfc4qk3YnfrGQ4PQF/TDqjbc09iWADGPUZILaByAaZIs77P7mTsKvPOH+hwsb
/axOM2X21JBHWdVTMzNTrZnAbYWjLVMMC8pmvOx8gVHgIO8elskGrxxUo2oFjAOa
ayrvnVRZmTc0BtV+YYksJsicNmzamyh2tCdMl+dHZQ3jRpyw4z+6bACGd08NLrc2
n4XidO+b214lbuDIZF0uBZlHj1Bq/e2C819rAlg0BDlObxYs9gJSAOCT1xs5I6p8
CkM1WnbuIDU+Kn6T8j8Ye3Nd9HqKcrlyoq+r78dBdklcLYs/RFxexvf/LtCeVcms
8LwYuN05hLi8uKyw/UGS641QMqvcMtg2s4G5ADAZUZLqOSiTu+AtgopIYWUabx3t
K1r9MS3EMspazrTCpWlRwDtTI2f+j8bVFRS6UfPfVow/CtRyONClPUYIX5S8AAfg
e3UG6mKTeEA8lWc3lVE4tLpXhkCZ3ljLElh/geIOmqbmQMlwZjs2qgJ9i54e7Yv3
uz5h9qViO9Q5/xKRF1xlPlcWJIlwJTqT9u90d9lq93duIOaMmYWJmzx4zJfARnw4
3MBm3dkNoREd9o0PixUS1xWxcsro1WycYDHcmgjVVefK4Re+QXwAf54oV9JK58zq
OQR3mhAi1XZ7J4q+C316kmTXSMR3UTJMWFcHfZ1H929EX6cdMlPJ4P3ro2TZQKn1
go0JUe1HRrsP7hE92lB0x0QS+Ta6Ukn2dE+52DJuHdmS47QkYHPPb2e1Su/cxGZv
V/HOnVZrLGIOrg6E/jdlrM12JIr2Ss2yYcH0TDr6KrNX8WHuYHmAsz4SFVLw/cf3
2oZI4hDGLr7EwHcbB0/FZ+01vG/XtiFTixVjP/TOriulO/BQh7kbHI8bnHtADrAD
m0sLb+k7kWdINzHNEBqJdH0OQaxR442GwBvc5u5+vvXPo9mf+BzzpxIeQK3U6jxn
opXKgsHk+JEcYVoaZ8yteHfvaYYGbT0xSjb072Oq8YQUoKAA/zyLjgpdaAmelz4L
NOnJ3EF4GQzNZO67xNMMFyz4Sd2tGmpxDcx/gSoTwwON9MkesMM3Cg/heujpYVeW
WVe5AZXYaOyb/A/aR1bWljQSAUOD19Ghe1xVASftimwCfNdZ2zuAyZKtORyo+7Bk
TYxCLcPlc1kIbyJ4HY3pbkSy9H1O72/84nrVpoiP0wf9P9dsYjcXJ8bVauJxu29V
Dmh3ZlXkFBdZqGrn5FuNjCeJ0NEybaB7giG+rDCdnK805A8+CRsP099+/Cz9jdsl
2PrZ5in9lzBqzjAexakDEPNSRSgVRSCine89x5qOsvg7GcIhxoMEcnv5dRFUfDr1
qELgqzj9HU2qQrmXWtLtu81ETYhiVC/AvZ/zaskalIATdo+E/jL07LB8xOp6eL3c
X0ZyHYT1VdyS0YRrSJGXpQK9z1/C7ZjtwNgpOCyHYYO7y/zSq86ouyDgkYqFEOzf
WcRQzwmY90wI8P7ufrCHmMBOlqOjMd3K9ueLz/RGvdtRW5yM1wL7B0dO4zSA6jGP
rzbsJhVmNrO8melUSZh0LGLNFAtxqI9DG7wFXiqNDBCYx+lYPrV4aOFKHuvQk7nl
hNnlZix20Sgt81y9LDpgXQ+DfUokQpqA1ElGPCpedK7B1JvYpLUjhDQvd8dR18TR
iR6xSduiQ00wwP0yH5kC8ordmhuZxftdGUMwkX2S1WOUyB9v0h6CQXON4ulnxLNf
FuWExsOUC35obORd6ObS/Tn5dRKbtBy8PiTW/UHKMfyC7WL8i2BMGcHcC3CFol2X
RH8XDFdqWKFA4L6xdI3xTIbQWwafmJYu6DVjJMV4pPb5qb/uKnb3ewmyAlRd5H31
+mvXemBM8QPmT6dpI/yCysyqPnrNGiUrqO2CbFCuMRoXixVBIq4ilkHHU2N7HkRj
eusq+LAiv0wCUvhxz5UaLDZlkaLDtUe7/lgptlJcZRlioSWNcvg2ioy0WSrhCx+q
YTWsee8jH35UmvI+Rmmq/9JkYowRe9RuzDquS2s4J3bCMrrG5O5EZsXzaD/0Uecp
XW6dbi9c6m/uw/0t/0bcJL6o8u7ARcesHacicYLJ10q/AWxhSih+4/mbHyHwNqUn
9ZNOrzXDVCT4z8DmLSMQk2kAiCAIobpxZKMz+amuCrI=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
KumWNg8HpDobrFdOtRHSAXwCIfKfo/yTH4VvbSyBRxTDsp+zLYfICpi3EbHnz4ts
62g+v7aeb9OlwYNRQNY5seyZ46GDByXjru5hjS2Wz0V+qXN2nYtKOjBuPDT25wYq
0qcpF4jGPjLMdxdb+yOuilmHAP8jXcfPm08R6+Onfw26aSJghi6SIre7uBxXq2/o
U56SFdhHzcmwkS4QwtDSPUS3aSz9vJnB0oe+23MG391M/nZYwqDsYoRMCobJCkoJ
GruOIwPRp5TKLuIT0t9cY3lZQRsDLCPwQiBBXR+/Nug1Tm+gCHJDNqYeC3Z5Qvaf
cVZbCS/oXu4jKwXbY4i/Lw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9232 )
`pragma protect data_block
iDCs+EEGQD/t4Lrug74YWrWZCWv3mS7lB8Hg2dhcXIiYM/uj8cHt0UedlDD7Hb4g
8npzJ37/2cm0RP9gxOAk3tXfLO/tz5Zx5dliz8yrDpnyVNdPkhEUtKKRxvP/XNo9
oZl7lmQZ3WqtzXl3fH08VYnZU3RBsRj4/Ns+Qhs7dE53uAW+Q+KhqI7BLHNBQABo
EmV7p0bvJG/LEk7fUqBpdaWz15DA2T6+ldd2dtrTDOlZOsaS/OUvi1uebFXs8bC7
I5RGzvDABHjP2jmSX6dZpEgnrUHnD4ZsUOv3PpDblYVXbklkQzPr67wOKJAR9vDl
XM2q1J1yCt0wiFj66jaEbB0TTf7jbT7VxKtunsgSKzsDi++TpsVxWhtZwGZAGsgN
KU56QBPR8YBBdynHUcsQIh37lP6h8/CNC+MKQYwPjaBWOZ+XzUVmWHKmb75etsmx
0Rm/JEL+2EDVZqtzaE+fUR1lBE85Mqlr8Iy/bs093SHZfAIhJ9k82gSwUDV3glRc
GO6qez5hQRvgNKlNu3li4H//AXEVLKvsDWMVOHVHSVh9cB5LbX61jvpa4dPPmEVN
GVAcQMs3BCyHuv1i1wRsnroK4pYO6krYWkuG7ISDMMw+tcCLgZEuS5ctGVCaDyb2
EFfuyFNO+iY9OCrIbFxaLLCqkPcbwpfrh2cfiK0tIudYF3YoTyrPsSXG63/aTUmb
TpLi/VMlzKAenXsNJ18SoTIKdFVMLvRtKmfeB5al3ZNsP9ib2nBQBb93HjOsjspe
Y1AjwXMox26gqyHfnV520X/UXwmXM85Zh/Qh30qM+N8e5lcqpGyiMiDp58D1dBZT
fSLyinaSw92b3xssFQNxL/7pEt9tyLj6RBHbYLyqC7ZDQSr5CearXcMsdZFtLI3N
Z3eah8zom6AiTGQnEX15iLssecxBRYH1qdVyQfdTX1+KStxsWdtxqDU5vFgkTH3W
ls6URePWmgA7YmX36CbLVPEBlEpNpWKhaYLfbpo1vPMq/o9VPbL7+vGLziUUTA1M
Tj9FM4aDMTieQYfc3ELSyP5VfjgP664pUZGnlnczkjongn2Gt/IzR7uzsBdbc/s8
oDOFqNDTQHqfRrzEebvRvpROSkbxJoxJ3AvBNPwTjBIdMJMySw+V52bsysUu9QZn
DKx8Ukd0v2jYjhHxrUEuK3JewPVniDXtuo/iB+5UBsXN9UQkeM2+XGka77bZaCeH
NGCmxb1IMDBBHli5HTQ7P7cvdQN2DbInTxfFoiCFGblngIveMboXp6CWY5QYbpYy
TiFTFRsaWWj+w36siaAoMpZiX9IQ7xNZgGmF1FAHZ5qnLmySDCQvq8r0S9hW0zQn
V+Bs3oXCt6ju7CTM/Q+sWkVLj+PB+0YcXBlYGG+hWynRAiFT+JY6Spuj8iSEPNEx
vkWu7j7jo7P3HQ2dPvHQsW4acEUDXfmmXwqSOCOWJFkqgMdOIkVMJ41DPMjOw7Ak
FzOkJ99tn1/PAXvbEGcusX1ZmhRv+0BiLPT+MjE9U2wbm+86G/wuhpe2smHTvqT9
ajOPARFTAZmdNyHWdvkSjuY0B3qBIYAJzRNi4UGqJs+snKYZY6B4O8RJtP3kSEPA
OA9uRt9cJJ66ln/JCGy49n9FnaGexDSkUSIT9/DvM+VzT/7GFh9wGN0+nF8HH6zN
8yx15L2JsHij7Oj+EpobNU/yjflgz1nkOkEURu0G4e48HPeLvJm1hbh1ZcF5RoP0
BeTpAmz+gxNoa0pFVDEjnfOLq+e10YMmEBK5gg/Mvb2Vqr8CNDYO9kkY7rfLjhYd
W54+BHQwhrgKMR6kP9Jj6kCNqyGwm7UlFII09acZAj5U7HFntD0BN19FxX8eFxsr
cm3PcedO4lp5oxnpi6ej+q6Vula168oDCnGkA4oAA0YH5rov4PmRI9ATgTosd367
02/iDiWcGJahVanTOqx4K74mWbVQf7xmGr27XSlmUqnDvBhmcZEbie24Tcqe9KQk
4/QYkQzj/7wzAQloZpc1NsIPQ+99S7UQrw2Q0HM7Zc130VCFz68VYpPMWXPvjbE8
hncQ8oZWHTTrOVlXJ5YWIIW3rDKxhEo412nTcG781FofQInj+w4lBO6mvuqYdjjt
YVxXxUm0HVfdkCieSQSw/YKdaDZnxoGNVjtURCEPqpLl/ROd/HzPHC3dgAXfoCQD
mHdQ4lAVjdE0l9RkvMOrgCEPFYcioOssUQLoRuJX3eYdvLkapefUcLwJHe8Vwe7L
RHPHLAaWBfV9jgsuV48Yoqfy3hKEBhZvqpPhdv7p4MXhTMctkX4RNrRJs64gNaFE
FtyhvW8FxL2/pBkbjEEorqOYTou6EKwKPF1y6wf51ElvsqOnARGZXjNQQOXMukc4
KexHjLIZW4iiLV2ShmVamT1NXqSqI18eAQnkqvfacif/c/hA654ZLLx54MdXIEzo
PMCkFX/TIJ282p5rZO0g1eTxnGFX89pnZVWn1LuVEf7hXw3fUJp7EP/Q9+clE3V0
WtogwKhdY+RcbnNc4bK4PRBFxHe2lM1sCQGehkkpQlEP1gp38dC0gNaMF9zzeUQE
fyl6RzfAxgrUFWdXFiIroKLvqilnAA5DUpxwmKa3sVdpry9pwi144aMcM+RUJ1qG
I5Fz701XlmtbiYs8sRCoP4hL9/+RgPT8fy+7eFp7NRihtH+Fl4Z9IRvrwbXW4SvR
W/r/V/DTA+0GxK6g504jNCQwKWoiCJdAHmQHzr9goi1RDCRYvDpM+rJcQzYuxFTY
ONCpIf65j3w+vOuTJbGZSh5lfbZy38ZtIyNzZMx36NECMoeV65ADGB1vnKH2FMUW
sm1lUrc6KHqFkyR3QrZaI2hMg84zotpTBTdE4Ayu7W0GGPsFDSp6petrwZoH6QLs
Mt5gJu13PfIIoAmXRFIDLaGO8UMPBK7Jlx3ia60JaOoIihRnKERtRLPFG+ozwYLn
B2HESoHsYguh/zWL+f/0xoiPAYqSYJXdP3PnXib3sm6wEeBprU9/tmVW7pSjRVc2
BGFj5H22rbnPP+Qb+ajnb2wLnxsYoqdYpp0vzksM13nwE6ZVvlsLKMMHHy0us4DW
bDd+2P34u5qjR85IfVKFT8V5aMKZQQJFGQPJ2W7y+tI7O6iLLR7Zn6y7oxLXDyG6
YTotBVmUqpiPqpVpjqIU8wUnWXSg993VuOZhn8isBFdPUknXnIk/DwMP1LVcRGRM
yFxYSSjwXZ9F3BgbKGVHmGyyS/erwRKP/7RiFhYcZSlJ7Z1xmnmTGGqizVz24rNf
ZoPAPC5gjXay6p3XFOYiYitjboGtjgkbaVZo3JYOT71+ZArEWWqC6W368StM9ZST
73uyD1Gszj5W4V7eczY02oRE/aterEj5qN2PEK63cseriFJpTjoAUFXrK1XJeJKH
mlnRe5Ih13SLn6aA22NGLgT4AU07Hv49MA1u3Aiwzi/TcTw/m2fxRQIRpMdQtmRC
1ZpuTjXdQ/EspOsgFJZw+S3P4bqNMZ64lcDhEwlKjTsrkKFYDArwbMaiix5Pzow4
b5rn5B9AAuk7MmelfxQq4zzfb1VPfbSNOfdehSJRdGW+ZkJS9Pf+7p0u71+jmZyi
jHublJf4UfHI6bJ77z1+6DcsdmNBPRV/+io1EZnnzj6eY+WlbvM7z2PRtTNZENgP
7U7lo4rSEJmt/qv4JTL7MSx9gCjGMUZ+xSDHj69q5z/cHgIhMfLyVEqHsQgdqqkI
REYi3qgo3QAvHuM64sZXWsEjduNjeSOouegUAxsi4sLbJzFm7MpgW0bJs6TuYNCd
rp5mXLn9RvAUlJ7zocMLAunnBUI0BWRfRSjg4OEfW4uk9vy+3xJZ8Bh2OldvV4Ba
j3YmKjEOCzvOxK41xoYvcde6NcgnxJqlJ6r9hVo/xlhdHmBcbA37XubMlUlomgB0
NQQDsrG0pFGU12+3Xu3tQoN3u2S1SPrSFNJ57gqhnOTbisZar0ZPotvFby78p5F3
Xwon9pEuSpc/G7twRYqaBcGZX+GvZEPzmWltdWVMerhmkR/KV1vt+UuLnZERAE08
NkgubIx8WzSyWJxFtQSK3NvwrzPChVRiQd8xGHfaQ80Pzb4T6ChmsggDDvQWdfC4
iMi0MfkQK8PMXij693GnqRTDW6UsjosnyU9mF/OQGBxahrZChhr6IOD7fecryDGj
WQyKDhRTYyemqwptPxnVX/g2ngdXp2OUeow/d+1DtR1zQJOf+DWZTZ/X8PHd2+Zp
6xNmsQsBLHP41WtE6g9Xwd/beQAm2Y/t7Ok5dbqAj72s7OYfUczNisBdVpdzpLwc
UyF49iakmSZbezt1k8diaz5o85BWbcwPpzarQXHn+GSVDOczJXo3jzE1/sCf+dxo
99mnh9xz0Mq+yFlmMReujYjGiVnCarYwN+H10RX+klorUIBi6yXA92huVgEY1DcH
aGXupoc6ZLQT11aLF/qD7zxFbTrzJbsv8w84smetoJwprGNYJOfEm6XLno5gWDqV
jmYzBxB7SNhvzcEoajarVBmYxuPhgZ7ClF5UcsrM5tzd5uTUcINcCy/oDJ5TWW0k
g91WLFNBGxqQ7KkIvrx1Z8vIpFR/9FEQD9v9eMryFSUB+h0U8rSybVQhcPNgsmlW
NR4TqrLJ/J4sk7kcn8q9Ij46txkL1ZM+9XSgnO5Uvzzwf1VNpeNxS/9OlTPhH2Gs
KGDISiaJTbXCWkLMCs0AOp47Ou7XFDxl1q53UBceelgRSCw5njQSiAWkpzxyKnIn
v07dyYf73RQkyk6TlYa6yEmIFpxO8zKlL6I30vNPn1oTKiOPRWEAy7EGPldpFj09
pIHgWzTbCQwLZ2B/C9dzkkybRwK76mjasb+dNjTNAuC66RoV4TE8sUuV0vfeTvtN
YWKrXoQOWJi1dNVqADPiQ72kTZIphAE7Q5oo+nOmTUHYEZ1x7CIJYpbMkBQa9KrL
9XPQeNVADIQ7icksC+UoWg7tDGYlgFyvrT9VefRTqtkWk9h2uarUfq4mXJvMKBwS
tgMvkfk3V5QNWWxbFV2V8g1ne5XWaTOPOhr8VspYk81PPxok2inxuCQfts+xZ8xI
Z/C1PmKjeHSEC/UOQmezALpQstdQbenPvD3aV/0FteOny8JdWGWw0OOEoi/JJ5No
UMA0yIRHuHndLNhmf7lYnJ0zkJpA9/UbOOODrw5+KuJijhTYgvSXgWblDNEXEfm2
RX8PAYYjYDu2tVC/yMiamIP1gvD54AchAncFYQPLDqsSt7HJJhHQKsOGGqKBt7C7
nKm9zOFO1sTXTN8NypA06Bdup5MUPonhySt4yzgPglnwN7lyAtaXRRpFS7XSzl5x
X83iG3B9+DA/h3vzTO/yJrmqhidC2g3LJo4+sWtdNZhBMGijTTRiXCpK3ie4sRoL
KkEcvFgpowWL4Lj6ikdVXVJFpK0jYrHjE/T125JmDGnF9x3W0hCzGPEnTpzm5ChA
8TJMJurpqgbK5UIm92Qs0gAtILayVpuJP/HQ8y7E9mXLhFAfXv87PhvZAcDy63Pd
bVlBV68VoTB+nObjqTi0spUsNhYmzJfc9HrR17QZPL+7OaEyyIZkATP3kP9OM1QM
0bUvb9kOGLXm1NxhsLsoTg9ti4ssRubSjOiTLeUM6OgG2PL8bMf0i4dNBeDvD7/G
VB9DwhVJ191O3/zRi8OXININxPbN9mRfaQtZtN7XNVnV+wo38O0U6LIC7J+bbAFT
A54vwIdRmV5VXBUqtmzSAe3vGegMvlXHclaLJ51XkS0xEFm0Sq/pKyZcxXKs+HyC
1q6Sz8w+rHsQ8oQuq2uVijJqOIvLpY3VnUx9+KG0Sz2AVY1wOR3jhgbivuOrCKDu
rQUssPtP3SAWNzGbabHGEX/xhewiicY3pG3FjYSihHuFKZit6hfbnh8nMFvd5UQo
jOZ/MTiL7R3Ux1SLx+vR3UQLw/x4dJRiOf8iBJ25+4vdHGppywjIoc06PmjJ49zf
WR6tplw1i5UXuIIvNOa2BUJTc2YbmigHrDxGAGTZ6HZr8TlWG5jXkqnq/ukN3fx+
l3P7sEDCBeCxHPApPCi7xHQA0Ngl8qcsjX/bo0EttUgv89HjtsLLz9jVkQsRPRe+
Xn6m7epeWrOV/wJTQVz3tGRZJ17ut6FGVzkShQzavSKTfF3pQFAnLxaK0qPpRGn2
QOMK99n6H5EB8sC3lEu2TR7QUvfS4gkyyBx9IByG7d8TeOM0btZJWRbU0dJo7sno
GJ+7WQoqlXq8REGVGKKrARvqg64ttZngQ/OBw+TJhWYCEKOgO3fFXmWCJ+DqE8Dt
5iGlz9STDqj/gN/gu++wdU5tX8xHLflmS4FOyb3TK20EG5Kl5/WqhRXpFqWvt+FC
3XzV/9aGf9tHGnRTIvKEQ7vQ8uEuzvydnriLo40aEOUIQm3FkHte+XS+whjVn/uK
VxQnOIhan0Owzq2Se8gCiPi2XUqHEg4gH1dPYdZwkkXnQlx3zQfHT4ALFhl53omB
8KI1aJ1ivlJfvEXy3f1s1jnYJ9QlRxxPP+/Dp2dmk905j3BCd0ZAg50zCH0vOW43
sjlh+xut5FMYeMmzqAyNF7UAOA82V6BjbG+UR+Vn3Gtuj3qYIcscb80ha3/LaAze
i0Wf7/harxnue5IY+QCmnw5ZCMeyKFzGJhunUOwPhHMXFX/LnqDXAEV1EbqDc1xE
msBWkJLakLVnhL97FbJwiLMJqDjWL6CMIVECGBgovl93AigUzMqEFv4U5y984ePQ
6c2a1S6jN1UxhHuyZeElk3bsYTEMmsAFcWW8thf+pJoeEBOsQK62SqyrdAIXsLvx
O7UpngjQcxjcWxEWrFO9T+6j68aUeYpDl9pP4se9GR8kXpPUG7wOztVFLJ4KgmsI
BxHkRVYXiRy+uvhyYQ81b+FN2pXo4d9kuFlkknIE0+5e5QwtAt1x32dkn/UFM2bI
PiqpK4d4BfAkN5v/ePjL8Tig4RJVmWlVvli3HhpArsrivkfD6vKzEIt69YO85NwX
Avr7iNoYeUvXyddOTI0y/ddJq8JUQHM9BhVygEx25rvcQft3meIs9txuwiEZoh6x
4xqQ/73yI4+IVzFXqTkEZ+uj5ge7eMYmZwwXK+gaPpq/btsezHswzzhKQNh58OJu
Qt3yv2LYclIF3lm0hPNwo8xH4Nyo5wl2O8BkXlxNE9pPgtYudyKYZzVQfvmAkO8w
hxSvn83VF53ZjPAWPb6ud5N6TVvHuBozG5EBVNYcQDzdKREYfvHlLB8YCSMIIIzt
9AsvU4/FR5WPxwAYi9HF4lgXiksmFNKaKZLJUbfZYTP8sMtSKPCK64djnS2hltWP
+9w7hahhspysLGCltVZPyQ4boWCnxNi0S1PTsLVOH5g583epMPYRwZAdHeWQrGqU
spN70Vc8RKiy9v3j8A0ySqC0SYE27Nz3NOhYXeB8x0AyMkiV0w9pGrREvK3Sla/9
QAL2O/Elj2Fnx4iwVONS1wIZR5gWsnTa+/x/pAgH3eacnMs3FR9mX/+ExKDHtq3u
snRQvyoZAjEx+ykkFx88EPmAmjtLF42WpIoDYyyrEKw/OWnq4BSV4Aga2olopBWq
UC8NyAtX43jGosJtlS6rfm601LKKL6gc5i6MvFro0QKL+eLqYOFBD9cip+oLpOQO
cDY8JJSdJApxtKLAN7Dlhe+2Rx3t8j9XyoXhaphnIMc+CzLWHP3X96F/nfq5JhcF
bhSdAYN9y52/t7f2yfl+ZEjKgUJFHDVfpNApzZ3V0YGRVYgZmNC4QlAdwsmdQVLr
dyAhP7FXMbjSUcAgtTxIEOE93oMCpJYcJXKh1/qua/JsJVoKVRZRAMnesTezxU4I
DwfrFP8bAThAZD5Exakjnansxqy7Rqc3K5p7MeL8T5bA154bbQ8vp1TM3jiDW8BS
HrGhaC6AFRU3DisoCZQAHipoPhD9utOwecyDI57bCbj7U5aq+GPx9kiGpqOKYTAi
ii+0bo4HES1SeZpk0Gq5udvCq8Qgm7dIE7biZDnHTurfdUR1ictIcCkdf8onM6wW
rhP0n+CrFrGavu5HzYngX0SfML+AKmDwOE/XfE9onhdvLvAUd3dTP0N2O/2tx0GZ
Zfz0rbEvx3vxOWwoj/vdl5pU2Xlc6qtKEo2UCPWvYC7ex9URdEnSwzEK73X88RHF
iMextPchMJYBsA19vQCSc4em3zqb61Jco3Sx3t2Wv5XmKsi/2I84/Ta8TsJKPoj3
qkvbCAKR8701l208Fj8/ppanT/Jl6uMDVaSTH3CS62gYFvLcnj8dls4G7sIDUOdD
quSo9fH7Pc/9aehzkNSeJWOMO1bS2xHh/CnuqU2GP8eFJrLNISHjBQZScWuMlzIR
jYRMJRPA9K3srsJ0SaASa8MWPBwrBkoLq4NVn2Bh9ChumVzVKrzLhFraek20SZPR
vaz9aukyGzMrbdJaGfuRaV3kBJqNjOuCshjm1Ua4qYGlKNyBxWMypywegkPBOOkI
UwqvKr63ZkT4gPuFZ18pQgGyNHDfB/QvtdsXMR1nRoc8YoJT7Rfy/1HgQlqG7+QM
7j9UcbXVOcZkGVu7x/plCOK57URmkGB4yRTZqwspyDUJb0/TJURpgMVh4C/bSvAS
fmkOYWWP+pryeaBbXJPfMpm3aJWVfPqKaLuA5okM82ZVRuDMgV26eJbYWPlb3Oi/
f6nmpJswBHgYUMy2jdAUB+Jn4aUTGD6xX3hC2t9EjGl3lBHYIkSdXH6riXH0zu0O
9RJ7ZmArDQbozed7Jxj6F0W7W5mJIEWMchBE3furk7KbIoehpxBGcNSnYp3PDa08
EiXYICJT57JA4Me/NG9+3XJV4YYYzEPMqwVHvcZph5vyRYox3R05Ir3JI534jWU+
v8nc2MWTCYHXpuo+EU5mX0dRCh2bYepZIsiayjJnLCU3tFEuYdJT5gDsEzQj93Xp
7gR9FaIDfk7xd/NgjCw6pDXK2M18yJ0d5STJUKFBz74wrQwOOKkD00SYpGvnFvwF
joGxUxSpEd1KKqoMXWxUuq5q0sU5kk6qx0Vn6r63v4SMt6/Nb0Lk6u4/3ElAYHwA
NDJ3/Qqcp721CtK/pa6ULGH8xwtf0jqgR0JorhAA9QMqGIcFObaO2VOlOCXi4ZGE
7LZwfSAlm0gWfNbKVspccMaalM5NoWzbjEjyqFFNRWH4eNmysVa0e/I76Ad06zOC
l+WHXFMlNQusxzjCe+YCSpSkben/cnw7QTyDAz8Jr1/NEuP77dcyubpN3JJk8X4F
lSfM0Smhf6qpPpMMl4c6Pi9L9mHOCIopDiHa5B3QBAx3c16HXzcpWm7Jq/yMRmO/
4rPsvd9c/+PIl+6jkJIoS+wmJGXsjaXOCm52TjAfpcUKu8WPcxE8UAgrphGKhw0w
mMLOWSBiZI20+BlPHIfWrY8msoex/8QwR3VnT1XcyXuHLgh9h5/Ijs9eUMDxBkVj
usJsjd1gzqb4GnnmoDQYDkibjcfUYw4QHDjDsuTieAexnCiuYT24fsiBwc2QM7cV
Du9CzlpSGZA8ZGuHz7JqFpC0I87aU3+gnabdN63shpUIICnVUfrYKda5xIAEp2WF
SvMwaTB16B6qqszJ05qSByLysrTfJHljs4+qEh6kiYJCLBvtRvyuUOfw5Htfe5AD
S4T3q8FpM/xRvsrul/l5upBhy/i8CELDE7uqJJ+E7n1Zf5yiKY4Qm93D7YVbA9f2
5mIpYnFNgKE/c66MMu23AyYWXRzjYnFk+6/EoxFR7QVXIkRjqZbwKUReNMxErQqE
6yz8qEDCumaN8APEGEwZkwld7IHAFaWiguRV0cA6gsEzwKYxwvDqTw7IXRqrlDxV
67rEG3py7cGc627wnJvzPImahqmwAbm/kBc/ccBL3Gmn/93lmlsr/UUOfO+XVABv
CXovdkDt6d4nMoWWE7hL7oEuw8XlaGyrUWMagkwrgKWZFVRYPxDOFRrqYGSQ72gT
Xd80qpumHaZR8kq9Am2Hs5WTf7iz1SFb+BNNAvkjMEC4zYfHpt2VQdy40DD+DLe3
QyVF1LwQF/EWaCVkq9bp2v/0pcT3hxKB38yN5sal92cF2jsXUvx6lpmKywtc81O2
FKadtCqGfNwePfYE9mPO98d8ii5PcDwXsBZ33EMGsgoXXIaSb514Z48Q0DUu+f09
n0NrqQEI0IDpr0WF2JOPJhJm+rqnawlNYORKHCFZmMZWfULUEeYTArrUj/kInEP2
yB59/JSiq8DEkz0tKaHxC62Y2UaIzc0Ij9CxRkXxExNbZhVarGwa4rEybZBZHHx4
f9MAS+jvoyfLLZ1snTjeP9NrdX65lKdwuGqAefVzKHZGEBmnEg8GHd0DxZhQZHBu
9eX4kqAuPWJooTv6maUnBRbjSbwkAAaxXmhMfvV60awNfMqtMe9gvAURlme/3xN1
UBZ17uiQK3SOoKXZFQiperdk35H3mzTErkbMfNauq5AYU3XZRQidN4/FAghPKPWE
Cd0Y9WT1M6yu02edLuGMl5SvB+y5dzk+Ntbhl32sGtLpP6grCTyElEDChv/OKXET
t+mwh7BOLS5SX6pG/mhV8ZH7K5vBpjf1xQ25k+OyYFXecJ40a0vahAK8lUFaL4u7
wtD791jNNA5g9kSgxtwFQcg4543wb/soS5Wg8UebzuDZa2f9j+dA6CnOZxe7TPZ5
nH6IsOzdq/QAXykqwwOOw91m9/vLLTX+atvnuqln1QaKjys4fk9xpnCXUX7Gwf7b
2RdPnR19TrIjwPUFV+6QA6kTQ68j1L0AJzbdNkdOkWRvpO4Ey173KRcYlaEtv4uf
QYBotIz+O0Z6sQkvbg4+wGg6vNKKv2xaAQ9Mmeu5vRDlxgKrm+mCYHEEz5XDvlod
1HcIRlZkPMy+o7s0TOB6lKY12rWc4mGjJrKzn89jYC+czxbh38km+smaDK2HDGhW
PQkXazwSaMhulLthzlK7M8+N9OBWYN3I8BciqzQy3ZKhIVOWzx/eNJJW7LZjfITy
YZbCQKgtSSwcu85+9as/juT++werMzNOrXU/6vjHxqyPYdZtQ+sjrfSHXjlduGv/
Wqvwv8oQgntzPDFz/tg2UYdamDXFbro7D40KWK4W48WeBGuv1OVL3yXSd54i/DbY
Iap5SNTqgBGPdOplmscwzHvZA2sQk8bVymBOCb9HnQdsi6AWECCotkClk90DSkll
yBdWkLTXD81g4OLUgSStB56Pm7kz1pYF3Bafo5pTIcGTPDHTRJhZbFhnZuxr2Sfy
gyuSQ4ziXgxymJ9EewSdPM7vv3gh4WNaU0PMMPIAqRGrUd7ElYWxFk1p2rMkEpJ0
xYVZlZOCnCEXZ1XS5yiqMX3oo6m+ugzgkq/bs8DJQLt+1+abbmkK8bEAI61Pj/Ql
7SB3RDz3qmh4xP+mN5Z0y6vGwrL0BO65XUJYZ6nWDpK0pJHLnPI18Ptp+SnW01uH
/p4syYSBZCYe5NKCRo9kwmPTj31i2gFkQLOXYjALrAmfYe8RUweMKTkq7KWOuUCX
ZW7mOcMS4yhTzeGsMy1I4jMFVKoVQdXy4ggRVgmlZDu+UH9NjooVWJSTuEiqV1MN
35zL0G2kqzcd+FT6H/Kx7MlDWumdo83P6/EAdsYwMFI3CTEtyGSMHFe6k5Jxp/eY
j8bHquzSupgyFggvNqRhfmLJQAdG2camYGynodBCFgiEfk9xUUFxG5UVGwTSzKxc
g6jiIs23ADPoEL7ZLb+JLdUI8A23J0+KY+KW0JOAOWVkcAAIAQxKKnWllkf7GFeM
QeJFXWab5u0d5Snv+cMJVmeEHzwiLH/uQxd2bLiqV0dG4WqdapZsWFA5+Eog9VIe
XCeeF7Pj2h1cjrS7Xpbm68Vm0gRA7doFZKD7nfGCIuaX60Yn48TQE4xpUCV6/Ro+
C2ksUP0542RoLKDLK4gf02J6KpXxdAQlzCYuBcgGRVbsv+4n+vP/UpDZhtl5Tr8h
4zeoYUZOGveWMqSBM6VJMLMLctVLmXEx4Pxh9VeBK5edYc9EEPMimzQ2IY723mJz
TSgmS5HovN+r/HMSugbVyt7Vq1gYJrfki1hEOsmI7s92p7E1GhU9EO/HGFZDtGds
l1+dCGhoG0nOEA+Qd7iED6nqPQIhJrJ5U36vtuUpD8l9pGQsXOwIF0zmSVbzmslI
UwyqFnesIcc+kbhhd3J1/BVcmHY1ATo2VqehxXtKwpfRKXxX2AOg28juW1ZXy8kJ
YEv9IrP7n5NVxBQzKUc76htxDGQzJsyrRQIJKvS4J8z2235UHS7O6CBtCPDLS/F0
VGCen0ZE7Nc3lI9NpZWGL/hN5LIwNBNq9vpjmKdqef4iPyebfMcfWmU80D5ECnx1
kyKx6wSlb80Ir3G//DgOLA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Y8a03G+M+DQsxdn5qbcGRKWzanmJN93ooL37a/xhLj5zEpy1hai4eG29j2PzQIOo
ScEdAKxMaYxZkaqiSe1iuw8tPFTeQxDoFJF8SIiBmPyKaAs6sXOtxs670MVnYU7q
sZ/5KHYpLczSH4/pQqW/wUjVoTWe+v1rfLBEzq4Z+JG0/tIBoD0FcYpRJTGnH7KO
PSp6fgg6ltSEAzmRo+2TzaEn/SF2KtwFefOZJ/qPXBYzQMzhvkk8ehxY0HsT4AL1
du+IiaTDsebBCAgAvy3GKGJIWfBCwttZEhu2mUzKcmpToqcjokx/+Ksnsg/xtN8A
b/uGm6de0kOHBEXbxCajfQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14768 )
`pragma protect data_block
K+Fn3T6fKpnWTHUihgyfLIKTtlja/S07jT7X4r5RhKpEsA9J4vR5zZ/eT6aUQ7bb
3aqhgM8F/H4EtFYrpX7fDQMgpiqzZRTQPHWLWtk/cl6uy6cr/5aa6Y5IrhZLAYiL
HCXuq5uL/6Dir+m4FuqhHHEgh6spYVJyWLrGIhu9D7ATuln0ynQvidhMv0jGG79x
A4OXomgydjaa9mC54sFjbBRn79WS0Z6aQduF4iqzml/yDYFTU4j3Lc4SvZeDl+5g
q9HlJyKjjHgs2RN+vVxYJ5oR9rwCzfE+ux3s4x35EY+gYmii+Yb/XANW8WttlbTE
7mLzJiCnRX5cd9DG0kksZYJDjXQk/gB9wwxMiy21q1i8Es1n6+7YSxLys/CAb0Hq
0WEjfqplzRJbqYC/rqpsE2fqmuTfYEutV88QFkcSd0eSbK5FYcutHzKqPzfpUWzI
gAmwghOH+be6LMkxNvYh777s1Bm6TWPkG+ZpahsJCS6VDZH46UrStA5UlXuH3y+x
zNY96VdNPBveovqw2tcLdIiPbfABPWEVNV+MCTGeVQeTCmTbp4w0vHlQNspBcyTp
jKfhCCiLOFiD5Kr1JAnV/FAMf9d7MtZtXgD5GJ17zM0mgexcJ8NJ22B/NCkexRoW
P+DrEnR6hzHQO/o0Ebgiu66E7DRyif2DDa47QsUmehfh0uYy0gkzhaGhaNlvftSH
2tis8P4H49X+a7NPKqBqj5dRHVuFwB0SoL2AVk80BN4Vp+wyQgAGXgQsHQGg2oZy
N1CvMJyC+ZDxWNMWcOe9s5nYsgoHpDtaazCq3Xe1EIw45PFIcIoBC1T796HWYc7g
G8GvSSePOA47eQraIvs/VaZfeazBdlreVjGw5FWr88FQdGfs//cFgt/7AAWHI4ru
fb0pjuIhXaFcldR1ClJzjn20/y2cDJtsMWHFy2Aym5+POgxSwyLIdrWteOZmJL84
quzRU99AS0p7tvs72jqXtVJ97MaZfmt2nQHve9rT1sd1cZLUsqQk6SQ43CwWuG5+
3h4hlaIA2wbxHX4euz1B7GbnPp6QIwx6KvTd/lDwVPsJMTKY3MN5mOIC7nXTBKBr
cxWMItBu8KSUcoADwUlz1qAOd91SLZXfrv2fPvoYfhQNyDoQEnqf4tNOYKGl5lS4
xjcNzjHzBGXwadHHtiqUTN7Ye95rXNCzsoKB9tPEHpiLbqRShrfTV4lWxUlxNo77
6k2iRA8P/Hs7vw0TDP9bBTQuRYDaNO7mbxCrD1iMiEjs+FwD7lJPSCWGs3mNN5u6
Zs44Pd+95oDTS1UyFERAfFUPicAwca2CffwJte9chZp0LvdxIiI0vRelB2T8wK6J
dTMj6H02J7vWMy/Eox2RvwQhF77Hs9xGJa6T3fQrU7MgMXjSyVHJsi4Hl2uCQj+h
pTtPU/eJdS7eaIxefOYaNycyMcQ1bALpvyivdn4fb2hAIl/3J097mY36+yIGb2nh
VnTiaOmJTTxwmOkYiJPjVcvsWbyUtZp6zAIThdnWiOZs1KBM0McnrNG1O0UFtSO4
kN4xs7+Dj05XUW4UyEvJWpQ9n7Rz8s/NLHnCElgD3NrC1blf8uy5+Vx4pevLZezP
JZmD/DqnrPxSaqGZE6xldSL5RKI2tR9prUDdoEXKDYKpyM7RgUNOLPX/yKWtOQ6g
zxe0mkViWIet23uxTQjfFd4+cG/Hxwn01ozNWxvQmVTk+2dpkpY6CR6fnkAyfeSO
PyBQ1n9fJ4tVgLn61cIcjhVtlUPwiL0gHnZ4BUdNTu3HfL70W7XRBi+F22CrAcYa
d048vN+89ORFEDPDFDUF9IPPOVzc2Ts3IoDJe3CfmwBpCib+SD2ZVM+NCEPOv3ot
8pZPwm4W+qGReMXg9mLUtsAFxxCd1FqCjq6uhJiNl9fMtwu7jUOM4tM00sP0TfLJ
0l2lsQdXGMZpUQnsjgrevDwbQWhA4DK581VZqUKXVbKJCNTKWoe6u0PCDmkxyQ1y
oAFU645lzj4TRCu/3HOTWXhX/NzJtK7JM7pi+HWsKptzlPZHiJhv5bUDfMdsGkf9
YtXBpePo7qFXktzd2Vid50XpMivJ+WLbUblgDaEPcHQnpA78SCicyidjO4Y55MXF
4JIDotrIj8sExRFEaHp2N6h1nCRp535yKOHU2YIkuoKnZrplNIRvjd3VTJ3+OH0r
wjcwnwdAYCfYtbgz5MO4Y1+vVO0philpQGPGcsQcy9ZV9b55N7Ue0AjIV36UgfMm
r3xqIOHecpTLmeacwq54xRk4cLrD6ME5mZ9BOg8rRto3LoV9xN2xex5agKbclWwL
iyGcDRFN0ybN+DoLKglx4mJqYgj04en0Hgx7s2FheeQqBY+vTzkMEBPkE0I1uoLv
VCvqXljCC3QM0Y9eSWY09A5NwO2RHMFHH7XRdQIxNEFZzYrdXZ2WnmpMOIAt3DsN
9SVEhieCoAZOCKqACgavqoisfzHXTzvCzBQm406Q1acTPhQ3nXqYa6uEOt2BmtEr
NVZVOD1rSq3O0zGlzmXuhlhtUVtKsxmRyDV4Q33uMUt2CxDYvLdJkwZ6G6UBFogm
mQOzYnYBiUuTg7sK8vVRaDpUMaYLltMkgmjjREKbOUjIUGLEFoLu30kC0HljbV+6
5NfuZ6JkH5s5VbnoDY/dipRdfGvSjuqgk2laq98BUYs3F8GwDivA/2Gr0FZLVfVa
/wUVAMyz454yWcwjSr5AP5avz2brEiH32ZvoBLMx9t/m38nNkTHAwKoVMEYmjVgK
z3f01NZggtkNaA96cdtaCCOFd/rvvBWI6fHOZindwWsirA9sAp8XXizSSF8oH8UQ
N2eOyWLmM/h1UcmtQs3kn393A8z25hlMV6sePiKSLJkzA+kbVZiRONI0ax7MRzQ8
rsmZiOx2O1J4vXGumTBLOa+fEbBjJhx5PdOQs8UKSETOoeNV7b1Ks2rWfZGpQfi5
Z3a2M4foiPb6TMFHHmFwQ5/IwEyBD3Ywb/RGlUxJZk80YCesVbRDcKgbWwefzcuD
9KsDE1+rJrGFtaUpP2e73ov8FdbN9CsLmJoF2o5rWGn+APeFhTMLqrHxVG07uOo3
b7tdPr7ODKLNit8dCk6RMKTmJe+eVInmh3+w/kt7mMs6ITumS3NHmznPz7h0Aii0
U4wxY3KD81FO9Q3DucbP+uPqHHEepJKlvgE0HuiLTC5GBAB310tk55pwogd5ib8E
7YaZDAPC3hbgGAZtqtINN61ob34DvQrmxDOuxwGbgDzYGOVjOsPjHcUu7RynxFhE
xxVYHtXPVxT+tEa/74ye20kJ/v25O1dkbZ3RnofkjkiBKDLR9C4VdtEOGBvAIY0h
XlzG0ih/Pu0Tcag1r8fheSvfg8qzY29741YlnHuC0DTYjkYNhTeirFM/+Z1fAfGr
PFAq0aUgdUZv8SPngLftP1rtbl/HpxryB6EKErS+4k+ncufZZbbhsTz7iMf0Be7l
O4SZ0SbjldxWK7yXCMpGoPrD+4UUt4fRUtE0ov6mGGOt+nSy7oiPXwsj0WmzLMiz
vS5VgNELzdnjh5JeQ/Qqoc2xFloxX5arfbX7QEmVbpO/9HocIOJL5IQ/CSWaJCA6
FiDHxbhZFuF96DiMubttppzJKe0ZnD23gW5voTw64Lc99sRSv9sTQsDNLdRBeKow
WK7yY/d8PVD4W7JLvw4U7O/mtjU6EXbdDJNzuejv93t5RnCsWxYR938+UDms6Z8S
UfYUR/mHzwvdcRuV9pQ5PKX9oH+2A2x6oqUl6kzDIOcMEQD54SXRB6OStfnNATj+
oG5fXmWMHHGWr8NDh4+yAmng/jJwluwaRcOzpyUL5BvCCqnZxxn2+wVRLORFN9We
tubNKLP+Za65k0OmBPh8/zjp1+5+ppWbrQeMSxQ7dctLwKiUtdCigz/Fs1p5YIC3
JokCSV/keNF7QiI0ZoellHqMMwX2i5UJ6V7uH1N9vo90IcrY/+CcH/OMjdp5dxzx
GkRpHlpJ56J6NvAfulGoXijnRlc+oM3Lx4CrVpR2Ppe5QKHOM00hAcxlU54aNIjO
63WAokQjNU8IkcmxzlirtghzgprAj84z5afsl2LZtYK/Djib6GWBKl43nYaJ3sGI
PwPNlZoE2FbSe1czexp1iwB7MCiTDD9N00lSqzJ6ccHkZ4/l1oO15uOVz5N1jb7L
bZJdJlx9fuvIq8C85lPiTBs29+3N68VVGKr+328W90eHuwxFxCQ6/PC9aBboCyaU
3zf6LIH4wTxFLbjGBVdrnyC7DFDsCGXqmeqDAayB1cAcKap7KjiWoHVmaLh6+uPE
di/P3L2vJOdNkyCOJPL/Xyq5HmtKoFhvgw4d9iELMWknfsa3j4V05w7Ysd/MJ3lH
O9LiQnO89sfgBDE23NHXsFnslWeFuxZF81vII2eVjsC2E4tCl/twCrFFY5ueJY3r
8dA8TDdqIvExxDUYAizIfYBjYIBoD0gcs2GVClnVTYfMub/UgXIkk3KJdzbZCMmN
1hwtH5qRAOzZtIx93QfNiD/064YPK7MvwizpuDmg6TxCaPhoPkNTVrmN9wYieFN+
UOjVeXAWHQl7Bxzra5Y/Sf96NuzZZJEdPvtVw0/4NbGkZid7XFRNeFKsqyngD53J
qRFvj/0HKmw/VbD5tSVeGHq0mBkgGkmgqgIU3s/gM4YzOdq5FhEszazaNYfg0f9I
zcujtXWcisz5eqH4o7A42ZP0TkEz+uMIfxZekwUbPb5Zv2npvDuivgboAoL3BQu4
g24rS0/9DOxJymDoKJGNF9ejsDd9LJuhwy/DNODYa+DNBlBZtc8yZPYxPjh527JK
05+7k0LbuApNUvOKGH22/KslXzu347e4O3YhS/ZCQmHCdSK2mshJIEgZ0Eu3zCVD
LjOC4eZV8L68afZ8kbjquMmeU6OxUdUvYjcOX8K062fSC77oU4uCzQpoBA/VYGPg
/COr6G2LCD/MMvIvVWAMhI2IZeNZiPlWhWOxN8S82QLJscXGttzEvdYGSIDrz6Xh
vquTBpbNHqDsT4rLnw3M84mxoRbXl0QUG4O3LVzRMD1vNqlmoiTFknZ5CtZQd5al
26N7eRGa7772mX6BBP09EXQN3nU8dhzP0NUdn9frkkkzubunLUwcSdHqxhOCBQnk
aBtch2NZrhAQoxeIiGzPP+I6Ru8aho+xOcM55LW5u2Kon/j6An/0Ztv54CCgJy+6
sWHue0VmOzsVPX4GZMPKuH13C00Q0xYFvnXj+w+DgkoZAqoqt5vdxLdelFBGSX/w
f9vKg32LU1TYTpCH4NFeni4dhn/F4lJbalClbKn/FuP8s/8Hht4yTOiovm+wEV/m
CW6r8L5pd8NlIWCrKglI3/xPBnI0+h71hJyWMlw2wE+OQE/6E1/XzkrkIOEb0E/z
qXrXA7xd1FlmUKMevXQaBJDsxQ6weI9L30TZfDC0EiqfZSSy2avEjOuPt3oGfOPM
V0cUFn3nOOr1LNfjil+NQk0pDAo6fBEQ0FBIyEsPw+QjOmJ+Zw+13ZqeVIbDXNVm
SSlot/aGxFNt8sP+w7wMyDS8UJPMQ9gk3MmaERJU0SN/kC2U8xWZu7dXv+P0r96D
rcWesLQ/HX2NaoiXkoDLjIRXpXNpoprxkz3VHqKnVoxfb4qpexgU1fhdXDIopbTk
/ym7fNns3V88yH85mQ7jC6wD+Ehqal/uR3ISjv2ImIVBGLcxuoldhCil3LQeKDqS
ex5/eurc241/MHslv++NvxnS3lhRoQeK2NW7wI34qgNKRggjUp1yN1DiaiVnVMNv
l5BrhlDjylmwumxqDsHSa6/jhkdEmTDLc5lTvuqwi40zRL8/xWtYJzP4xuytenT8
Sms8i34zWBKNvAUCwD/yKqo1qQrvfOKpnCe7/4tm2MlReujgC4/nTPEE+ZinciH5
+8NvxDeoM59Gpky3pMIHcaBGR78PQL+SBcGdRoTthV0JRx8dBpdNJSz7+eVKVRuI
yO4AIMxJ4k8ng1uchzL7xobsLljfCIGW6V1ZN53TC9YAz6ZJzE948nflmsmjj51U
1IRpKbYtmgTdXkXunfJcv81bojpFbPIo6NCFSC6UwRNeqNyONrkb9T3gKCMVpXmo
OFR8/Rsx+5Fmzh8HzMQiVNWHe5bzYOoWAQWevbzxQQZJa6/i8UnL9UD31LbnySay
FAHhv7Onpq+andofLnEOLFfHiR47Mr64H9KK5b1i0u3Bre5/UMz4GE/037MU/H97
l9wmR79wbE3Nv8lhIMmZMGvQOb0JsJsC2kqALK3UqsTaAitfBuoHXVZ0qXSUmIF6
2EfAi3v3WGnMkDlqKlNwga4PX9LaQl9GThOErfF55yBt2KwhRsC/dcKU2rlKf4un
J5y1jCFx29IspIvk0JhxjWunf7FJxh5Moi3Gu28g0Mc2eKCOewxGb8la22hfoWgs
j5x2vNFHSG+/gL51iU3NusDOkFEOgV+eukI6S7BOMnLiVoJFV9x54ZgH/ffl7Rie
NnS5zxCTVCqrP6Q2yYsifUUvbgbwTCxRbEsEs/txoxaEvRK8TH/nLZaUK0rH7Dbw
Pj2vHu95G1nvTnHSUYVQI1w7ot4X+CKsUWD+SAVvnxGop2nBFYOFUOZUBUP0Erxs
u0G45Xmvm2V43OZtLyFmjdraonMJKp4XGdULBP3Tq9qIzNI2Yb6+6hFdOeC7WOFz
JQK7tJTTpw/G1SbWuOa1QUQp2YklwgqH+BBjWkF7BPvipXZoGtAsa0cCNA0V+hLI
f0M66d/4wZ9jajxGBpz21sVdLkI4081ELaDK/90dWxBNucB/BNmdq1MVSEw51HNe
BQrZbXHbNZsk30CFLpKX2AGkelkvUbaM754A3plgtqGQgrysRKKTFxnll7TAMYaa
q8L/bgC4H2oJcUSzCGrJbf51Fbyfv29UnejjL7Im+p9HTATFuUoxtWLAGjPNddci
mhwqchaf2mEg1IFYGRF8QVQBFE8G0093kdEDfCNnAiQNlbrEiyQF6VWp+qrO+msP
bybNaYUu0K6MgNgTSTL5Kw8S6EodEviJ/0i8g2DwAP4oCQ/UtwyJIsPEEDKa2suU
4EuQk97fBwE+jYHWSjtHrtj54p/RGEQ+M7wpa2ueWHq3Zk/fSvRzJJCj+P0eay8i
YnRsu44Y8j9SO2Jd8ccx5+pYjfuZBcP22PW+ak3a2l2BAFTJyBKWlMWtgo4ZRIN1
RgWWyX2bBbYrOHwkScJ/L3YKGChBt7jN2qRbJYdFXimh4jBf6yX9B68jhSF4IB+8
XhANgezZxqWGmb2+TEyix7l2WjJaqh5Q5H4Ud9Y4X4QeCZ+SK9/YhDlAn7En2jWV
UpjoZQkAyWpr+Z1GvOpioAMAaLV4Dv9UauQftgF69ODx10WWajjQsLrsvETIp9jm
dYjJ2Y3d5ej2ugi0Uk06JciOoiJOHvmU61Aj5M76iqgDEecpR41beeBXtl+rweNV
dv2u/CQOwLvOotzIwa2OWuUprrisu/IGh70T5Ts4G8I5p+B6VQs6JrMwsKRCxYuc
ownn01KKlWHSceYgpb/RW8+hrP9f2V3R9/5hWsj8xD+vlmI66oSNwz64qnmTZXQm
XDU5muggI4D8m7Fl8DktJVDJDn1LxlBTGBLiGtgZcnEcGFUYHXpPl6tkVaCujlaI
m2pmPM6x7HNNepR/hCdv10pe747yDoUA7pkyFmdSJJE6c+uEwxB9v+EvNFS6p4D7
43B9cp3+7OUWeHqOL3K6u4iLeyHFGY43uuux3cBDGPIESNICw2dnPXXywP9yGFx2
a26XmnvF5nBrJsetpnvUzNLz44V97GtZ50Yb5p43UjoiNHgThpmtevU3Ad9loXYu
YE3HD0mmosjIBKvE4OZniFud1jtTtj1v1FC31H1lln1bEMUI/riD9VxVdZ8dshpi
Wxsaq94pQFimhczb0LfVP4mIX1o2R6m5/Fw9rOX0o/lEKSfzpRM+rXwplXDLUxzC
1YSEY6aoJIzB0QecTG7wumr5Ec3/UFWJN4oBtSkDMXCc9KxdXjoxWqVyam7nmsGf
FTx2rFKoTsZknFkWouB4aKoAD5Vp2iWTZOAHiVcGGEx7oD8qltVbJ1E/gcun0Pss
3ok5qV6NTbGvgjbZDruslJO2nr68J2Z5a36Nx+l0oLSYdQVx1pllnrG75IqHvU8K
LWfaOZ6hRuPIO1i9ijcgrsi/PlfCkcWhUYIPOGrce+M8KK0O9w9QPoYBTfL16GCU
gJZYIfbsPDfNnxgqMr1w54yoVTlg8Bci8Pq0+5w6iVDMaJ0SpbRnOEgsrMXJ4fAb
u/UgHZDRqMTeVxYewpwQpchq2dSepebgb1ghqa+HtMYWp0OYzbkMfGVY6jC460uk
jjFTvwRU4wApgibuynIXfkW4Y781vDL9YeXc2QXtlAJjRq7GJi8EA78iqbBIVfbW
fk2T737vES1i4jU7BwScgCs66GDzm6fW37bIH9Wjm31OJfi2iFv6RmHlJf8y37Ni
ia+pRcxFjncPvwAYaMGVo8lBHL5U1QNnC8LcOR+OIaV2aSfxKkaWvJkvKamIVu2/
YV8e+TqDnZP5Vv2wixZhYQpdzDCvJXk1JkIHwB4nXOgfIXTvwqiro+d5E1inpMp/
2M8uErlMVpmgb7kQHt5sL9BHOMtQ2FkHgNjOV7O85JFzXNKzedVcgp1QETLcFXbs
/jpW8f6de51+VEbgcdV056K8Fx2sPrZ1IkDNEPU1/RdoEkVKtLMm05F8fc2fDBzD
ijHC4GGM9mgnXeZILQkx/xUkoIASmRnpiz8rmd5KBlOIDMAYcbEYqM4sz+orc5TH
gUdMz8xjgr07uG2632zsixp7174FZmz/MZ6dBBfu8hcekDxAqVpVLGB0FOfjIl87
ITJ/tXr2zBvPfHy1qnTr5p5PuSaDGpHM7tKKzYyN4ic3g6CcwwH081Ndf1+D7Zyt
fTkcY6RioCytTXCFETRhrJRXw1KxXuSXtlOMSWfqarywczBR6Aiy8ZhPnuM/+5jb
Zi1YZlvGTi6meDiEiq7ev5+nae7NVdCxRIFvce6ygFei9pMvFvrIrJmZ0EKaCGgp
5g7jfLOlIU8N8bCiERTMr/LFV1vmw4vjLhNaLbRYZE40m/ZBYTY7yB6S5u7bzzbS
CUE5YO2fjAGEsxvywOeC4aWyiMBMUDqXgXglZHAELXe0WZzO952/OzpQzw150uQS
WTO88IX00kKO/SA5WJ24TFnKypParylcMgYd4EE1ZkmIXTNwmKeo9P6IYJ/TTc2z
XQXQy/xP8p0Q8c8v7mZlITgMgU+D+obgHSzlX3gdIKKAjNaU/Re/2v6Lq25Tkn03
7DseRnag4XgWRAnVXG+ObNZtoXYklwouRmnTtpL6SikyleKocHFvkmQ4AbI6WxrK
NnOazYHaN3jNQtHxyrlXvFm7m/OGIpDX4d6KQhGmexxDRKiQvYUSHBELLfInbUke
/jmMC6KJFWvZNe+x+EJ5ooSFzagdG4Sr95C8qULOMFQRJgjt6zOWqqa9vhuzM17G
jTKFBk1e5V/VvKGcUFQppy3xS6syyg4pMyi+0UFRYrau5nvx4fZVE0oSr05PgD40
/D/nyMRZJX637L46yYJ6yJrpUGtm5TcnVXFW/3MFqEO8RZ49bF8lQt8zcuoJn+h2
x96+/tesNwGjMcyqC1Mv0qnWC2DZx9J59L/jFosOODexQGr3DYlflcvCpc4RGv2W
mif4ypuRBzp0DFBDaG2h06o/KZWEmaiuop+NXooV/doeQ7p0kiKNoZm7GVrQk3Sg
2mWj9gv12TwiE8r5GtOiTm16VM62N1YGo+mCd+c1fgva9FDytMr9LkRSNVAnEA+/
pBCjwvihIe5FPyYomi2Bz9raAiV7CYuTYr4r2RtDuRuhxTGyN8xcIjBc1YcF3PBR
IvwKCWobvkambRnPnhEcRJdXTIx4APSLEauoEqk2qpQX/jBnTAjonylJSVo3RdC7
v2FguTfu4SM7b1R25Y7QeJDf63gd/bHaKNRstrm8UPoy+E/v7DE/mu7+6iBCVSid
x4rTTplrM4YdYfdd55nwcTsiKNPjzsdraRaiRMKNuFLu0OVj38iA59D/kXTRXkik
TWg4W7eqT3075NP1GlKtS9hKPeV4bE+I33ktK5x573vv8eN7ZiX2XZdIQ+OEnSzA
SsjiI3ZmidkoeNGvtgfzXj3Av1x4QzmKWInmU94nMd0SYrWrGs45SNMZEa48WtFx
W+lA+B0sfiwBeHKih42bKIWIC2tEDGNCggs2jl/Q/UaGB7lMtzYeEMRR86cN5WyT
i7Aqmd2w32hoMZ1atWGEEkvrepOnVGw29Njup5XX/RF+dQfEbvqxC0M9IfnCorC8
+E/sUQD1CCOl34u1Zj94uXpxmNc6QhArRJvAhh235sjpC2wXjIzGeS2Mi/VcC49M
i8JK0gMy99LJq7B48hc2kPqRNSvgPsWOwV/rUKDfQc3ZDsViZf/Dlu438JdfRI/h
8RiDTg7HKjSWVm2vqCW/c/Mk4MnUxOOo/IgTv9s+KQ+jHJLcLfSKnU5SFGu3DeC0
4fUGYVEz0P+xTsqBlq9NF/ktsr7SJFHmf7pX/O9dO9x7LxcRbMFeLodDhjh7Jz3z
DluqaHKLEL8gfWEMctCVbLH2bhzCIufPEN41R2a4P4DFUrd9x0suIqZ8f5hbOZoe
C+pjZ5XvDrA1hSBDFkpuQsLNNLGPYcEK0Y88SNV6+5t4hw/hSSCxA9Ua5FkBYXcO
bOOqLQ2SLMTMtv9HjfsHVnFurOf61pP/X64XvrP5eR7E71ksl3HvNIrjJXma7wUY
Q6t+fM3/mwrhnSU022Zkz7R3Z6wC4axwIjzCFsWNBaB8QPAhkBwTwFaiVrFSlud6
xr0Ezc5Clar4IefDP7sbGdH4z/9FiXP0AH7CVkVnDRSXdsaIIadrhTUEIQV22F1x
EJSSOQXxqoyKyFPGygE0O1RzDGrX6UVz23ngXwQF7u+xPduUMAwSQ5Y9Hfet2nGb
wdtFqvp2QKY/AmjdyuEUM3uXkHb7z+eO9SCbp8AohHiUIe6PtdwoslkQGEhZZfx+
U5wojkDLyzDPe9aJXPslqgc8ej14MqwBs3iwDbUaDh4sHifBCDTixpIQgCcaOZnq
ptqA1YSKOF0BEd4eiOsksA2KaiP1H1or/wZI54Dv1eae+D12PXSl4d4NgQM+v1V7
q0vRlcB1xXqVycpvIt2WeBqFhveuD0wrsQZ4cQkoxRyiJ4e4sA6HJf/Ps3diqz5j
c5MuZNni4WJAnwEqrJalc+H8K8ckELspdgxZuTeXkvXM+dJE69Ujl1WvXnWlT07d
dRKpt/MYW5cpFLcxg1eJatZvCBo4wcXOwpC3hBBs3oy7o/E8Jnx5dnwwMgM4dg2W
cgyAMHRIbHHRiBfnXyTv8vgvlf6zZ5tvjvKBhK44iBXLntYofxblwgtR0K9npuNX
2JemYQPAJhKOpGNLaOql+ovi6UHAigO64ivR4Ip8o0mDQvIBsq1cfUh3zjkk48vX
5Xqym5jnUd10J3BlUDlcPIURu9oOrxSJ2/rgjZ7NQo79UUFmJ2Jl1GL+9kQuyca1
zphzkCXq3mRXJm8MoYjIaXXTLN2wz14uKRGRoen3XMcNiiFEwSgCQe+XuRpH0ORz
QWaZrn8qk3DlDAiN/kwXgev3Htzg3hiyBzCIHxFXbVB7s/KZC/kZcJ0txSgFrwgT
uvF7PiVgm/HLoZ5K6VRVyPu5JdH0YByD2wnQhnIH+Kg1ZndHGYNIbNpY6DlR5/zp
X6tMP/nJIVC3gP4v2Iy50V2gmVeLT8MCashZkHcE+2rP306UbRje2VS3l7z2il23
eYQZCYED0AINR/49kPRc38rb1Y3ydAmlw2RV8qKIVgdSCz69N8tm68HIuua3AGOu
jTkiJN1tMsi7Oq4R7jVPAiK3m51TMApU4fVF2/BdQgFVe4jYWt8ecvxK8+1mUvpE
hAxpFOgA+4pvJbF1Xpzt1N8WhfXIt7STrbYg9+W993Tup2QbPu9ixJqapfOSartL
aCpOUvCSDPN191i2eWj1DtihY+kTlTtauZvp9OWzkfFdCd+xu+mBKvMjwhkgpSwG
bqyr/EIy6pQ+E6KXh776/T9ou2at0TUIxr05u+YlI8ZvrLjJxzjaD2b3bYecciKt
W9j8ft/ykMaFKBR1GbYF+TLgL3Xm/iPrUg2n59nX7e0//gjhHJmeig46hy4lqRVj
hlbaBxj45jSUT8lyHhF7SvGQfrTD4vD6yonn9C3eOuXUFodwaSj8jDnSBu3p/QY4
zv/ahkhDrNNiHHgNahHN+9z9F3OqGjAZwrF+gW0VGv5LZ24DBKHLlr/u2t4uT6c1
ftACFFrVSeuJsNnrhhA92yXzKJctR/ccHc/yOy3NsyIO9FvOprgdY9ylWDLV+3cB
v8HD7ZK8ufDYC9YkmpYqSfEvbxWzZmhLjAmZfMw+ws3xiuY45ih7xGM6MzkIErJ/
Zc4fAO8zntrrEaOSF8BLua1VYXSgOTrJsP5QZ7WlH4NWBfVHNnEr8X3Vl+s0Gbfi
DyyfqB4FWk1wi4pvLUj1MK+QY0xmZ4Z2eZGvUFUiR3i8jw92eR7AXYr7pRxxelrL
FNw7yQI39O7FmT/NsGMfC1twh2VX6G0i14S9dFw8yC9A65XpsoUjWLHxLCvP9NW1
ruYmutQDX51zl2HFOHPAp50oMAYap3jRiCpigJoJ+3SJkTfEP3TN7Jv+3PTweiAO
5cFH8+X8RfKKSK55sVcmTiTUEeYTjEEi/gEIs9VNzYxMcvIHznUYi1CqydpwwOeW
52Yhh5myGrNNbssFHfYYSdhQBoO761YtYFeucay3prETdj6zjo+KUpc+ZDAtxvMR
qji52qab+aQem/FAzpycW++wPLv7hehp5036ukvsniDnG6AgSBZUYbl5EOvq4J6d
M90fL36qncF4Vin0Q9GvdWTeeUiwdFlM7JnBkeRe5rtt2jOZGD8bxZ6Ua1l3M92F
CtypyijdD6cjWAwN3OW20slUk7cy4FvE2PE6ItcGtVhUwXWrb5UJlqswaw5mXkWC
9h1tJv/Uag0TYte2Pls7UDtVw3IakQQqYdKDEMtHESco7/ITm9tIcevEE3KkspS2
Y7pFUEPgqbKByUAF6wrEqDa85TjB2YOKdG1qiFq5+gJpXxQttR5tS2HgZZAUni6+
uWkT85Hu4JTKV6XRIeIfw1u/C75KQHwJHmhyoGLvx0ywp7+chuhPzwrjAMls8D1h
0k8h3+2RF0kI7T3Mf6sAdcC/CFiU/FqPMzbWJfWBHAmbBdxMnb7B7cBck4Tsr8rQ
xlxKdMvKOfYMFLkdUPDN5nMQLH6X86QEIhLctKv8YckQSh76cz5SZNDg+vJXBdXq
sHVqXuU+/zWQXkv1XLXI7Y+Up4jDDU1cEc/Jf1+3fLIYiypDmGKWDb0znE2C4r5I
3V9pR7SSq0ThAQn0RiqN7E3O8H7oHBD8SUqCohoQq+i2bLls4u2SpTT3Kojig0nr
N4CtDi7aAAIEFS540aO476zf6uRmYSOKYzwgxBkvE/NfIPAgLEK+sNYWtVGF0iwH
ieS/qYeOCpRy+eSOyS/6sIiWjmtTL0tp7yNQRZ89z9XH6uxROs1lmdTGi/jqTOcH
hkWEDpE7PP6dpdbOrycyFHl7iAHbHYasRMjAasDT0QTLkovl03vI82z8mYaftkXT
W8jLbUNkC9EQZxiTFIMEQi0UNbw5RRDMFDgir0ybnq5ElfPSzhiQwtwjNBvJ2P9B
yL9cr5LxYqZ9ODLZlxwR1x/l2YpoWzOJP9ydOH7CtdANi1tjrjAw/87rIjqVVmFf
jbQ55ZKzoT5mE8hf5K2RevRNb/XCQaMgWHfSfsT0optV0r6BloQSnJRKfRnkmptr
VGnr1PnThtq+s/8Fhvu9pL2LkqpDVnFdH8vwmBOtj3CMc/OenvB94IIQI2Ct09OY
KdYRU1NE0WwyXXjTwItGbGhIDnUDJG36nVXdWyM5Pz+hiEhS1we7KnBP0rU0cOaf
FGx2puUeFEMHk7mxuV9L3D03Acz7/aIfGAEPElVhvAPNhO4Mi+YjLHNayaDvu/7y
gErtXFWLxkejgoukDKxAyYCbH8wB+pCdXK9zQDXysIKk2/euD/GPDc1iRHzoXI8t
Ose7RfirEo2zYNMJobdFVrfMPSbgVQhQq64cs+GHhZWSTaud4UGRqaoy7V1aF90t
wa714yBIRWjjcpyKwQ5lmDzSXe61/2DzK8RsebGc8pyJFJi0XbJPv1SdU+9uPFSX
rhB5kJe/RKCrFeMoGSL/CE3ABv7gZoDpwgQBdS2wjmiuFGUbNtjcpN7w2sXtQxic
GFp1HT1eu35wvDyYAE+z62R2yinDK/jDZcxi1qPiqK2nTRHJ3CVJO2ntEiD+z63V
VDsh6YMJiZdJuIE1PtEQkfteRSA7GJisXy3QioKEZHMIQCEFnBXgES0QqVWY7I+f
WHIY+moSqh9pigESroem5lLx2/0RLqcLrIY5bUaj7TZE2EfSG4y9rKYeqxy+0wJn
DgWb2UBpQxHeVwCZ/41iTHO7B6bv2yHLz9UXtn82Pss9yu7htt7J0CT3Jgodofld
VXroQw3pDp0jIZCBSNxbfbHuH7fgJRQPET4fu40S5/JuAUasEJEweHVoT/Npwx31
mWzauqes5Wczug0/Wf7oU1hImJ9hM8kyT2ah53qdj+jqWWaqW/JNwSAkmJXr1fzG
ib3EyZVokbKtgoX2gTQhFp5lcWfZuXQoTLOEstgt8u4TFJQHHXZpkZ8PmAh46UZN
JjFa9FFcx80xD4XDRjnnBlQlpArEL1gYevSQ4K/GEqr2gQyBqHnyW0+e4VYaFc4q
5WQ6tae4OvT5VA4ca/bJHGQLDelc/ItHo062P3rYNIeSsPSBHeaSqCvvz5YTGzxr
kq+VMZWXHoglEUHznYv9fUT8wa7edMrVfzcMEXnazyqw24y9cyR5RjtAxDEyydvg
Pwzc0pdXfIHNCytT+A1XAPjIOE8qSCdk6lP6ek43aIwfUmWhh2aLF9uuPdwYlAfK
UHXAFCjRff7eKZ0owReYpl2bfihZGhwogiGq58rR+xPzU4uxC6VHz2DUbsA1j178
Tpm+jxwOP0hp+BHiWEPaIHYoIFg8dNR2mKmpGiYtBMlskdQkt8Eo9l/+gWRXlgIN
D1GYhEkyAvq1eQOhkWWG5DEomCbq/T7FaKdqmsP+zi57Iw/7vrgEAszpaiXTV4p0
nsCD8keIoh/ORhua8znc49yOyZwdeaCDCcLTgm/rX1NEUipykuC0ad5JH+7wmgaI
vHhrL7x5D8NVNHpp7tDwNfv7PIze8ZnwcSq24bg74d9nSpcNQ/cpSisepN1eX7AP
9MGfNOkslhZztkyPYvSwE+6Cr3jiRWlpAuAzEoBjM26nx8Dbq6njvee6QD3AjPdm
Ybv1r1uPbCP7N8JCwJyxZ9Fzz40dWLMErv61j/Z0ofNaUvhdHa6sI2H0LLD2SHpf
Zk9I3KRB96deKRuYclABds8FiIuViUl/tldNmtwaNATBra2iIXML17950hoPxp9Z
5A7ydu5xNuqZ5O16frzAyrtetuF4ReC4rv1JIfn2u6lMrmNrZPPswN6yFj+i8VaJ
oSRaflBKpCfCaDUdV6Kups0G7zzK57wTZqaToCXB6cBEzYtSCd7dVtsNncgKC7Ug
Y7UKJObtdiW7lnwsWX0p2BW7ZP6gJhCRhIwajSZ+ymsNzhxoN00DWFaJBHp5ziNe
yMPpuWsZceEikuHeIlCdZt/1nPrwstmo/PxtiFgmRPD+rWqjGHKN7ETbzSuXvx41
eH3Uo9UftT2RhKb/jcYflDTZvthIdA7tqSJzCKzjJD2TMEDLg2qr1uCWPd8Rne+3
tui4Oqg1kQCLnsG3Bk+wok60mxk57WON5oA7godoek+wvkGsMamc+f6oVgVpWv7+
66L0VedMuw9YVj3prtNHORi1cp5TluJz0Y/9CHBcUGqjihDUMDfoiBEnOAyQeF+L
Qf0hR7iBihNQyUDPWUqvhEuzcI/1OJAWtxmg49eV4ZDCAI1CR1EoKVdooc0EYRx2
wAmrFq0QFDuRKT3HMuj1xUhZHE4Mr5ljQtHaeSnyOTMqIW8v3BQ55PkV2u0Mqid+
J6f69JImAzhijO6m3XtyV09t37EQWovq7lvaTjvVmsCYyB3OD/yaTKAFrOYl0RkV
VX7OrtJUmRBmD9eyJlvMlDIUgCMQf5hSD2wVNXGx4it1I1XoWm+9Yf/F9qI1TOdB
91Gm2Z3wtZ+JXwXV6ap2w7Lb5EOsJvIVmHQUE3GDGPWh+uKJd0rfPJPmttDiYkXZ
YylNwxlyB32wD3dhAT9xwOUUQs90MH72MsX6fhpAaGRMTb/gkuCAwR4SbSa6o3Yu
GgGHdoorHq899OK9dM/9LIaTiHLgFggwmeHefom4we/6b3AI5BhYZcH7stkOVveO
RytDgGOtYhVihnNNgRhjuNtf80JDAVd/A4XadllmMXknQox54kwteqe2pg8pMQuA
PQpv2Iudf20i/CnQ/rQkU1pFUo9Ny8W6V5FhkxhjIgQdSO5KidNSx6AxecyD2bJE
aWEr9nq+C9avkenXmP3cAi34WHFXI18vpDoI2emB70urQnISf/CgOj8FuSsGAKwh
l4HvzNnNadEkUclyrMgiGuTEiNzniQlqOUFouOj8dMHatiMlg43WDYIofHP5GJ6h
Qdr4Kuvq7Borms+p5PuWqyk1KqAXoEoN6rIhNLSXWBEaf1tGH/vVOD4srREqRB+8
CyZFnld0k41ETk01yoniVECOqqqqkNg+Mi3+2uVoNxZQTCqjWRehme0awzpf+1uK
lTJjXx0I/cmTz+UEQHI6XTWDIv7F7NOceorH3gcC7t+xb1i0I7Dn/b2oq0eCL8Y1
ualgzt0Yjrb0dRyBc6ccRsuzxelV7uODQCQwjuXL2b9JaLX05nDBFz+0Q9BripDj
awEE8mZqffJshTjBjlufWv5eG2SenGEjvxmoLBWiAHuxP52giXUILsWk7uNgzeG4
4c1qNI/i7zxX3gh2pOAspIWth3pp7SoGHS89RU/di7rKDKGyQng85Zpv4uFFVBnV
fVfE+gGuO3/J3qjZgLc46NZySeZR9N9U5JmoYSCER22lrisBjC9J5fYh5LmuUk1L
53e7dtlDC3W6n48HgIYcU7mGMdAx475/7lJ5oNFJK0lzqzt5sQrdGqBIFqODqK2W
NDHYyr3WpZGzbPfA2AthiFMElws7j1qR+Z+4Y5imNgPEtxA2CA+tMam6UoDal2fp
Uh1UYSOivirxToUJ/jowTl0ADeG01Ujx2YQjhbGetfWSJOGj7sulvIMrgfrc1VLz
i/IXGUqCk8BlqaUtXXNgj8/7jkPwr97gCSgd3kt2PmbCNU5/meo1hjRvxztF2GGx
bBXRZK2WQyhxSRrbxH9Kh/UJ5xO87ZYV19sa7fnOJmkPLUGhyzQkmjjE5OUNJXSa
erqlTU9b6ONbW8yEN7iM6hDUoMdWWNEGfUk8b7sPOeCBF3AEfkXaJ3EPrOc9p7Ty
T57DOM9qk9zH9QvVJmEJJ3eBuYg/06kjwa4S4nn4ZwIi2e3UY/+awGjGhz/UwB5r
+iWZ1aEMQlPH2DpVAl16EP/h1NkBsY03wYpGNA5zNA8NTBFqZzgjQT/IuY7q0DhD
f0vhXeTH8xgcOXz17+jVQjuFO3kXO5CzRcsP49fUIf+Ex/14lXntwVFBvwr2A+1x
HqjcwZxdcnBvfzvIrmyA2Zicc3TjWQ/KjD0ZXAsJm3ilUOB09yZ2tmE/FdKmH6qX
OcmJyHdAOqaFhZtnE7IF7xkOTA6AUQmhYCqq4wntMalZHsFUebHHmHV1cv94/GWE
FtyJQruByTQa4xf4WtGkG5ZD5vLxrpY9Y8+55eCfquzsSTyg0upZhN/nYtQr6s/L
wk8bKMf3OXCHRuCaaGQiEOXJFewIjPadBDyTagrBQ1qxo1B8XXLvn5roQv+Qh4aM
Iq3LTmfI+cNMJXpDHHpvTIz7S9BI+r2FctvJmLr6F3NHcJSyyqPqqhrJH92thEXG
EfkBeYB0UcaOAaUo8QBcx/KCS8D+Hj0qj28RwGnewNA+HIfaDbwLHVgUGKaWsMd7
kma1dYusEI4O6ixxnYO0iM/7Fs9bDWQjdZ8FPBAF4jRukOhJnTwMSfi3vr9G0m8Q
7uxHuX0QTA3vGjTglkek0e08Eg12aL5bprlJhlfXknHXH3eY+wM7E6hukzEVXjzW
rcfLlgimAsT5d6Uio6Q8EsRwlfKC28JA8gcZXKYvkBUbAOnSvlWW3udwmjtDkurp
gEolmrwhNRpi7b/aZmcoJkry0PJDY6PHSs2Lf2zXG4dtUpdA3KeRbOb6+msIZ54y
Y7a2Lvzl6jRKDlcLMcZQOS1xxRKD/4XN+jeRctL7rLpFjg9IMmiMXQizAYIqUkkY
NlNBoLe5e9pyZlH4o2GlSgSXeelH1eU7VgY246ZJAx3La9iGPM0VUbQFiPfvSO9B
L+eDa+tvYtRGQEiken+33iZV2ENAjoDV+HoBNxTBFatTTpuPcg+G2SZIOagsoISa
yCs8TrPZZ55EYIDJkkifuMhhi6oXnV/xRIyouuKl0LvIobuBHUThZOh0y2cWkEnJ
7XoLbpbm/LmntMXHWzaWIbnqwA/+D0qG3BMXc6YzesljMcTlrCUp1goIsVtym1TF
3t19eG4vpf5shIWmXVAGHrSDEfM2n6cyCHANjupnGnMxsm0HFKZmX2YOmhCg4xFu
y3GaDdDX+K/weWqsD/SXyHaoi3U9Ef2E+X7wdufLLpMP/Gv0J3pXZHOFei4w6f+3
2sQwRxKIda2hGyJzsXJ6eWI7QipRVvog8LiylD3h93Ur2YhGkWCcPWtJ7D8HdKNb
6lc7fbF7RC8IX7HV6M6NnSKtDve4WaN6JErK5FjpVwOKSKClABNEjryoFdSKAwBZ
cF1Y8EICWsd022IUREzgQtXTcEsYK455RylmjUGAoS/l/SD+h8AitZPQg9bqfXzu
yPBxXRAVz4GMytTo7gROtDl17YL6yWwVC6phvK7PiigZcfEtalB67VVyp8loJ6n4
V2pPzb/Ie64SNZ21me9l3LPjYPfoG0yTcZxwitkuuAL/3feraHOscaVU49rOAnkP
PTdxOWFDe6v0CGwy9DiBorUULFoGDt9p6JaCS6mtXi5B/fN4MQwfEGFUgzhKfJnk
BCkoShxjvREASBH2U2Z0o+hju536uvfTOCoq/GHLrGub/ZB40X2JWXNU3Y5kRMUh
R5c6fpPvdUpYfmwmaNSU8dqTmAn8WTSfdy+qPrezWFxB/Ta+C1Qj3Ew0swyjmxMK
pY6SetYvIQTOh4LhNAE/he92J652A4Se/IJ76EkaS8TuohxlWM4C4Qgdjs8rh2bI
wJljLLpiu8rKKna2fA3r5gySABmUOItLG8qim/XE8XJyChb172x0Mn25ujUemgDQ
1jODwT0JL0CMReb+8QSIanJgmTVfHmku6blAErbWMTYhwX5lYXIkCrTgPQkraq90
RIe2Rl4FPBQvzWTf8oLnPg89B64pQH//67txU7r7Rw01J7X+PVD92LVJUNgHaExF
OhgE02IDjFJBgOouWC6bGW53dReeoo4RxrLxEB7KOhsXGDOAXoSJVyMCBrPFoAc8
EQ+0CC9zfplVn/dnfjZw75pI+WEkeEt+PsvX+9xDY35kPh+CUQBN2P04FZ4dOtkX
FLqOkdvQsJ3koDNYAhc85bfc2hdTi6hCpq0YxcnSdhI=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
S8yXTVYSoQL/3zYuwgbWjaiItkNX5TIy4fE6fksi7yEuh0rfcehE0hForaHSOzmJ
U7mhjPOumcUUJORmR0XTBk615tQSGiKFeYv8L28vZpCgiMTV2MT3NcFFV6GY50aF
OSlIDQgKIogW2tFMM3W3XuNhyQbbXViuvYz9YY8HTz+9ltGsA3wHlF8Xbl9lYg7e
xUQs7MYf6em0EQ+oUnJPoBQuYIWF7RhsI7/Lk6F+iWsKzunttXIL1TZzvLmi2x1K
nhhDMVTCpxf6bFOb08UkNC5W5lGFHYYKzsKWo2Rlp4lYfrWclvmi4tlueYQx07mF
IO3x30RPtnmS6w33RLPQAA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22512 )
`pragma protect data_block
t7Vzx1+lno16yktNlWYimD/1LhIx+FxavxlEmhk74SfQtfmSDF1je/MravrNUi9S
AGtmq0IFe0Yf1dYDCxDNS9cB8aRz/lqiN0BqIj9s2cQ7plYlWMEhAiQtVemXJpmX
wST4xb1vk0MhooNHYhz55LAKHouGjFzXRRhgeweGor5QwN4QD0UYk6/NDoLSpe7C
UZFtPsh21+WFm72quC7ZkVpGjg8xByY61McIHms7QyK97LC26pgYk35EIVzz/wIe
rUJvg2rtWV42Ptyq5o6EKULMynQJgtas1Qw73GVdiI77kBWxCAuQR7woo/JzeoP6
Zuta+kOCNybeVFMUUaP31W0xCMS773f4mc4ABE5wah9mX04POY8R47TGShSNgNpe
pljvqfn4pDywrC0AeAiEhxk+CKVHgCOt+cBcPalVzJ7miP8ae+79E5w6oMkjqa3W
gaUc7Qwijh+ejeG3RGKkAeQvo+NiMu7gXTl1BsPKPc8iH8l1mmnbROM1DyIbt6gM
aAJsj25TqxHNbdkWX92a89dNkIMhmyTmJbCnbl0mxOrm0ap+C4inOPlEsoT9Pir2
vR761yDTTkIQYwosMQTBsM8ZoTDHa2IeAKL1kmgiNa7/OZr/H3j2BwqBBo426sWh
gLdL6JroDocdpAIQGqlVVNuflpc8pOR2d7nNGYplP5RQBbWvZ3Vc1JU12IsqMbiT
cdBKTfpWaK3tUUtT8vm4QR3BIYar+DoJKA9f/GWSggbIrbSJGLyG/GYA99suMbOf
4hd2MYBDL1TaGoLOxEM8Z5Yp13wtIlBHBh0SOU351fXa32zPMJWlq5TYnz5PcOHn
56l21/r4X3R0+v1tZOFeXtlUMigvBd1DGJEUXwM9eHZzb4ZvD0aMJQo5YQE0u25s
pnkSVINV5ynYEe1dR4CnSBrepKWuAt3gTkUd9blZm2rJZQX6lNoxHAFbyVloPtS8
n9oXRl634L8uyZBR6tffe6G6Y+Waz3J2ZK/ypjwggjF2h6Zk8H9TCPiUgJJ+M4x2
i8Gp8wezgU4qn7/vm/jXBchoaTPye6/DkyGjudMpZe9UB6R5zIdfQRPrBKBUvJ7h
QmLXvnYugKCbH3N64VV6Gf05Qn7LbNaYfPRPczr7fs+sXFRAsPKFwU0mxTZKp2S1
5LZDZUSyIQ0z90waZRzCDTf/NHce3ifwkJw7gJdqzT78yttdZNvG2/VE5s3ppbAi
UEZzo/FPajzT7rO8fcpVMCvJ6aYKP/Q9sLcR29fNykFAliG6BMBiTCufXagXgjii
uksxSKtxfK7HHcdsB1r5ip5/RrmSyCnWo8kWOladguCyEa1NQb9omA15xIh7OlCB
Q+nPhd/HI7plesUkali1GACnMi67mQHJGMvgf5hY8yduDxgqGcidrxp0YI/cwYdS
h5KBMmOBhQhyPv4A2J9V/dNMnzRbiytGBerHzgARyde0WXvSaObL6e2IPi4ao81m
TsEjOqC9AfbsDLSt1gSB2zQkbJFJH5s1N7cAG5/98Lul4Fzu5lvY40kv3fVPXgJg
GzWA/89HuvyipOQbgPKjT33heAxanc8whXpxh6cE4q9HT/xYiglLu0pfwfhR0YHM
qcutBzj678CJk0LIbOYLCx8GPBhL9ys/CzjWzMbhBc+ovQ0x9bZrUVikfJ8Z7v10
sFrI8dYhuI3LDK9k27SPJB+8WU5bd7mfOClgBN7CNWI/54eNDh4cxxfWwCNfrnNx
x9LQAIm2Rdgcg66mJKuHNzHjQAMOUEeNW0Yi6gvUBZs2dK2XDDTUFyYgmRKRh7rR
bwloW8XBVwt5rUYNZAg0RQc3sf4ZAeP0G4PmRIkFp38r2o+aHUKhtNM4QvQrRv5c
ApKRGpslej2WoEBQgmW8UTZlyKOE4YbqSZJBwvzWenUO2M2lObFrG99DzWbcOlF2
13J0zP/lfOfJMb/RZij3BhNp1AeACtLIPkibzrwLCQH0cBLsnptB9rFvVJqJgkTu
zxBaVvor/I26o+QhVtxB80M21gjunPa2UkQb7EgH+F/ctH0MmD+lRislU7ja3++g
GL4AObsjW0hNY9PL197ggfGWgIh47I6WfQC0GowXccErxA0MjJwOX/YvB+7WthpE
vHvc0X8gtbbkzW0LdShqYJB/53qxE/avxzfkjTM3D9gao9j/S+Kmfn3/VDgpF0au
QlAD3vTNcdH7f903wbdNzcyvsgDL61tRnXS2vBu9ZeuM3SDjpyRjJagvDBZHolpA
8K77b8fk83UrqhE0ArY9WGmjhW4Hj40Fg3tGPJnAHGWOHKdm20uH+7ZSpomVej8l
GL2vtLauOK8mks10ZzHBk3zsm/jp6pRD6fc9+/ltB3tXmODxVWYNJUjvfYaXa6Ir
xRkMeOdnXAZCERF9Q2Sau++3Sj5nRCLPw+QRdE8elH7UefHCHGHZ0kOb2JvzoyHp
IrKWU6ZfEAPyQFnINAsLREQoRKYcAF2ZHtubGHSGPJm3GLrd+648L1HAETg+Snf3
KL8wZrWqBxSo6lq/0PBAQTcTl6BqkmpWKLADKXyttOb8cWqZXj8URxaGqClxl2y0
n48qIUsC8x+a0SOi4mIZxgRqnSxFA+hFASONeKhc3LC//PIOP+5P9RTJVQZSWRwg
ojgsbHG9zp2lyfhItePpf6Ia2a5y2aanO3AchPWddTwsuIdrqriW/NRG1a5Aj6gq
BecMWwzadMu0mTHL22NWIyIrgc0SXGXnVYtvY0WkbdN0Y4+ifycvYshssLOCIzCB
9ZrAk/gYS8B28/E+9sPd+6gIjo6Nd1c5Tr7ah01nv+3ZJj+/vtTRM28VJVJ2+6zR
yPXMFYx8rj7xoyQvQrvjjeoTspOE4acNczqthoKu/5h0EKfwAmDDX/amjjfNWgPd
GXhHONkDYPdCZ5IbGa4Mu5nXXZjUbC+qEaF6KR7+4XTfeEEwqSWeOO5pk8xYrVaq
eXLWzTwTSKpvxIP4x53dzRCCALXf9GFOI9yeFCy4paUg7ptTieGyzYu7ZdZZ4vLH
yjBs052tIKJXhJ0dKL/rah00RcemQ6L8ASN9CallDOHYApP98gZ+6Ia08p6nlP/z
rZ9Jj+OsT0OcsVKqu/aBMaw3ZQnBrsiwD95faE6OGCEsIGd9SBPPEzXdcr3/gKIi
Jgh1yCazkeitMeQ1LkgJtyCWd3ZzQwh1k3Z2pFfvrDah7qtsvoCabbySY6iXpywy
ArFL0L1yESJMhwqEyZxDE241+6wlmpXHHp5r9m68ZxJBUwCcyo07d4FyuDrLe0ku
zRMv1iCxmL5mQG30gvuR1uDhhhx8M8FFCYgSdebwe3UmzuwzWHAh41dPWOOQHEYV
7gDRd4irqL8pHjDgvZE0S6mPGccPsZqA4jcBYbCut9UEWRfuh5kd7BUqUjIx1uoM
5Osmm1iGsnrWJSytGMame3ds/yrlHFbZl8ut71uwM+afH2xhO1hiyMAeQWjKwY58
eOPkJ8e34m5GSjT/8Gw8GfjOyPDHB49uga7GQwec61TohFEI8HJvnI1sUwl2jKPb
hGvrZl1RQVBjdc6zfm1f0Drxb1rOiDgbBOzhKsV/HEhSzAcPzfXr8wcfi+bi2wG8
rhP91OA9kSU4OzB1YZZsrfG0IF+q70yTvl58EC5RmajohfTyZFRU+RcWKy7yr4Jh
MhTKAE3Gy0Wh9nQ1NO9cJrWT40vVRS93/GcSnKffwIQS/wSflywAmzYhfl08/Yef
jpbQ8gu3BQyreRz9skVH4WBqn2GiXmLQS9R/AFKvz+Lso20YwIQk9KwUUWhx/jk8
kPo7RGjkLBFkM/EWWqjhNKnLZuPReLCXtCzGd/BoWwYPUYxmZs9fd23rWVJroPJY
wJN2WEsg75uXIMKoN+4ZUZjgoA4VXmuUH1dc2yDgxY/0LU/kzB/aobhvdKpeeh3H
Jea/gqIbAJe44hfifFzOnmRkmrfm8r/owWJxZkX70Gt45otY4+O8ZOc3Yjz5ZYGp
JjD58bnNwJDJ/vgjUgU4D0oCU+KHgnFQ9kBsR4SzFz7W+36AmYaXydR0xDXdYeAM
IXxuRwATqsrlJXDd8uGtBqGjQ3v4JY/A4qwnK47trKr5F1HNGpbhRkzjFQYVv9Iq
RJPnR+Nfb30i43qqY0i9hBDbIArZmd8MOiAUuJKm6yyUUDmrSZVrDDvk+WATG/p0
dZ7lqzFU+Uk0h9f9p+av9ennK5gTgwthH1jto40CadpwMh7dJj6cYtcktgQHPVVk
zMd6xTT3PqiiZ6cZKTmzg1t9ZL4e00QRFaYAbDCdQU6GydcvWVm7fuNl51BbJiBN
05XGpZtbbIvc8RpqniIfh6yZENHCZYLBuh0VE4tHtOI5Trl/w0652rbE8SjJtX8e
b5dX++owaFQYMYB8000ZpId7Z2Dg+omiGxaTwETKcDQbjk3ToGd3WkKVRfHeXbLH
apq3aL+Gd1e7WA5oTMMMAOucC3wRU3urqmOHDACPdhIPv6NSzx1YYfLgh80vIVvp
NeHJ2PA/8I7GU2Y2BJ1LuwLKHDFp/vizJlzsxd5eMv3x8cRu/KRMehy0O0676mt8
2cXUykqwpVeezgXf+/rBelnc6l3lDXJCqb0sXGQ2aus/pADxQ3R8HxbNgn2A8O7C
2TOAFjznvBx+RB0bNagT8K9WEIrN/vcx3+0FpLDqmTwGjLyw/oFVIITJTvjpBwO8
NIYHtUp3IMJwBQGQ43luC+wuzL9TKTYjuSY1J+/87/PV51CF5pHQ9EFZTL+rTGn8
L3yOoYjJcn8f0O2QWlPcXJqrUM9UJpaQoVb06DswTDQHiNzpTpr6OmzAv1HaKwDg
ieCwV8ZtdORl0oDHmdO9cdyvzGhnyY+3Ltyw3z9s9ZIBGRVeQZ2LhdxaSvH+P37A
Fv3CblA/KkY3EROqSdt4ePg4XE2EwmVc8uNaYWELM6HPgjh+RsdHRHIfGiLAzKhJ
pgHGfJCECXQtXaIjxIUQlUq+XIURg0O1eiHitJRJkqevG6wJlja1oDHR3nbY/pZ0
TCskHcQIWl14I4P7co0VnXdjxtA5dzUGpyIR5ucCFFyx20A5kV4ow4KfSUWOOrln
nDfbYVcb4MAs9hYeGr2YyLHkMAJ7jMByqRDr7AXtsASJ5Wk4wHyNGqmQRUYNsMEX
swAl30zQnjC3IqYZHdCM4ilo5akfUX1ki/5mpoQNo3gnEUkUQC10qbuIaibOwUhX
+g8bsw5gGeAH/FYyMWGjzrGBPOIulxaF69HHYFXHvHWDTYW2NEP+o8BQPpbzdH6h
WJsQCzOt0Mh7kV3zxCn0bni5ZGyX4JffqpMNXj17piMgJ/juWiRYG5V3pMR5eBQ9
+h/xSLWLqPbX0dx2FSnSPahOlrRT266Ioz1lM+TYog8SD9/wVyGThQmTBay0zZyk
RV7RKzOyzi/xvySL3Z//qG1WySE/nzEtVrr/dZvF27isVPSpBsKkuTC6p4+QDRPb
no4B4add6hk0CcncBaqqpphzd49ghiZZ5Y4rDLi1u539kU/yZi2XhCk+XfL8d4Tq
1iDtB4/BqhAJhL0rOJq/60HCVBddA0kQEPdN4bBAPrxGSE5CXy6vc72pgAMGAB4L
/yRYBMHcH8ylnZpmw2hjg4KiGyLRgR7uQT/U6X6jlb4tUn7N3Z8jnqt2uYGYhk9M
rZOZN/3JNrt2/7dIdzZz6gVEtYAs/4Wjv5QiFI7bsB2bMXMO+Y9sPxSGApV0U0H1
Rofjnlbl/9x6hsDvrGGGGW4bJonVqHw0Xj+Qu7mDa/KlNI4FqJ9mc/3soqc0MoIv
wEWgdVt9LvdE8Z/v9y4mfDaXONWFApg4KkRVE925Y5bD87w6VMtrQR/gNtRYq3y/
sjWqlPAfCJp/bIivCXcoo5oMbcLB/KegOenH5qXSnGnQ0qaxcmuNQG6ZY0/lp6Qe
rOK5c5XkdljlGM5Q1f8a4TN2qHAWkSQywKOlLrnQoCBR+xcY0PpuZW7nIf7HRQcD
ahOhpmAsnUhLTu0GIWj1VciidvRR4cg57twnbbEyCKwa+Cl9tkIuosD1BfzY0SGp
GqCahJUiwhbZNG+bVdU33pfaPia9cVnHd+t/UiOs4EG7rdidcO2JCncOqMHd0n8E
w2cW1UO86tMYYI5CuNHQ1Hf3ESCrM0QX36s3KKmn19eMlPh+72Dltmiv24o2znXF
9eT1JRDZ4TUNLlysjZ0eG3UkPKupsC2Otnwg4eU8YVqTAdSr3g8PYzQDdK5TrF3D
gQGdJwnPEmVzXqD+X9GsnZoIWmsPIcPK1E6Ger+PXbTnEgMVCJa205wmkLNGT8Wj
VjkeWo0m5p+QvF8RbiDRrMLK6ACrMsGo8lLeWviiwgPbjXoOO/1hMrwOkDOoxpZ5
8EsmAg7uyvA8L6Tqevi76OCA3f6/Oz3S1XOlxEvCR5zWQpjJreSTLZQiE+BYWWBP
Ic6gmPDOQLPYO0tzOi9hbSzrTzcWGc9r+GNghaKo9lKcFMRx2M5hNglgJX/3wRN7
8baWtuV2PsxE1W6euCJhB7AzBjvjvIlQXS2L/2MvCKKsrm/bnuwjEQHCuTy5HLow
vtNjXneTOZPcdMw/AcTdENu5Qbeix8pzUklIIel5tLzvFlo/takRUEiGXl9RxucV
ZwfS9UkJXc+xvmMxuPIkOayOJfIDjOosqPcqBto5t8BEHXdP5ijcKM3iX0zr1own
/Pqe9PWzc33JKq2KddWPt371LE/7M3NzLl5gYgOoKLdmib51gfGz/zW/w3Kd0Y+8
gHeOyA2HOoRYYCumMP9KyrYQvMRguRS88enDwmYhsiJHLe8VessO4lFsfbapiXm/
pVZ89qMCzRMTdKfx5T64+YmBQAEkYIuR8SApvxbZa96j5rXqh+AAirH28IPYGozt
C+ELaeFSsfsWPnwv9/pNTfV3gT2HRLjTxkqmqkmUhF07gaFkzFokFGZk1P7paOLP
rqmMGPgr2Lw0+Y0H/csfPUrV/pr+tugrbQTNSBrDzjH6pl6p3qG/BA6Omw/qAKYc
iSgZ+brH9L9S7+57J4ZbiTltHk4miFT88vueXIfIH1pRuNIQb5pCdRlPjhiUlBMm
4T8o+eST4ncYBPigcJU46d+rAp8+fx5Mivgp5Xyn61BFh6ObNGiouDEUv5zm3GX9
kn+OiP7xKOOceyjiV9JkIC5mxpAtrgJ7BS7lV3Aqt3icekSyUutMvSI0/b28P5oT
cUdHUVgOManYGcZ6cHDTMnoToItCILeKJssGUv1EYo9ccA0b15qIPrI+JzSlpxVU
vl9D2n78Z8iCAI139xLqBh87zL/kYnTNh2F2t2jOQK0bdtV+w6h9m74d0VIrHjS/
GfaTazXfFkKOa4MvhibNm1iU1WI4hcGjGjGm0MQNlVQZiGk8DUJ1gMbJINFzWtfa
Nf8U7bP1HA2KmkYSSS/PRiK6n/Z8ItKkkEcc4FNndoypx43rrSrdznB85UBsObk5
sk8HNk7Xzsz7F5s1UAHlVJOntIW6BzOcBAcZL1vYvcCSmWadGSVHn7fcT0Ps0aly
QAzSjkK6AuU8+31eeQtLAUn1fF0kvu/8iI1zvpTDy68UFkMMFqbRscp3+tS97+tM
hkvV6eZTgPIMxRluztlUzykg9otv/9kJUWtwV1dwK9RdOWGmx2tsK2Otux9RCUMl
wSgGoHZWDBpKB9wRLAts9ErNJEcx1yqkygKb95gK3h7ULe7y8l1M51+Aup0Zv8vj
23cHRDz8pKCBmj+jniAU8S1dj+s2d8FMXOWeg1fFZCGaoVJL/3x5fnwib0v7OdJf
NXh0dngOH/SEJxG/Ql40BH24OVJmp2jaNdt8VNi8a5O7sTQK+UbCa4+d4yP7UKyB
0VVXh2cUMphjXiCQbW+/M7sYu0bIUX+92cYCCmb0S+lNeWsYiaXA2x7zktYPjvOB
ivC+sqWu3pLxMElr1UZlnBKpB4YjJ+nGcyFJIgDb9qpJ4kXYTUDt+E+ffXSMyVgn
fKHVxPfcs/XuLO5sVCUFmeJT1q/NE0jN7XaVseNjgNY92WEwgwPhTpDtVNSSKHR1
28m5nAAx6TxxkCfGCzugyYxuORTv1TVLjcbtYaqhVTdt3wf9ZJi8XWs/HCfF1BA7
HlwRvIY1Dz3hk0CKT5AhMVMS13d1+TEnU4oFcWe8sno+MTbpBPvqzcMRcmh3xrGj
VHQFIO4SccEXixfGCbxx2J082YOJke2fYDOOZAT3KpfM5Rx0ZcOM3csLn/kk2HoC
OcmhXPQ7OiH1Iazxxe17tFbth71mzJJRgbgojQTa5EJgRTXnJDLKpLp2rASJboOi
a4IFd7Pu4FYLLVRsz2flhh86a3lNwpPZB9AnMvYjGmBWTQJDlRn4xKXEl7kzUA6F
saUXmfkhYX4BpDdKvdP/cK9jgtQMCAl5xqLnblahDHu/9E/mZqNyqCL4cFsh4YCq
pRmYrC28qUw/BSwlAzQZHk+iCdGCKW19RBo7rIy/l8KSNkp8AvzL2Wauh/o02Ijy
vCCM/n3vtw+yAjGxj0MVzklTbABq+nZbi0NcaWiEeGZNIUczMd7Qv73w57pbg3lV
K18oPnjVG4qwqAO2kQFvFW4Aq4WztQBnjKQ9V7+lw3H2rjcf9E33TPjMCo5HH1gI
biSVgLc7F5UB2VZ2YF8E0ejQLbxdzUYI4/d8dz6WEt1ZGChbo9/Cwi/7A5SzNRmx
jQddfIfZjSQbXcWQcP4/EfDhyGutpZpSb0YIceJy7IBvv/x7gn0dzWBATTXK0ZJI
kAD8iHukGAK543mYLLejKE4P8hHUFkwemwoLYJJWerGT0SZzBbEPoBpRFye9MX57
z3lt1oGtknAUuEh5Q+zjtCbxDtCBJIq410ItghiV1+iwgXgYbVNSa1G9YDcuvrQ9
v06aYYWwNWk6baIx8ReoCNiZw5F1tjnDphtKo2Ad5VN26nIQaGn+ugFxHeou0TSr
xuqrS+oLwuKDXCUxeKCQZGnyhBlsLLD3ZtrTMDy+HO2Xb7KqEfycJAAm25Xh0spz
8lBxHHnbKr6PjNm30lUwnkWD/IjebGNjgbi1KmsoRawEpK5jegrLr/ZDRg+NL4Ez
NKs7k+wGAOv3YdvHsJdQeeo01tdTM1E9WZ2kbAxuEnQeDRl4NRw2Sl1rB68RDYwK
Wbus2SBdJK4hh6ZlRaWbtHJ8LMM4olqyoCIRx6ciVdNcvMdM+sieA0IyW1+/m6lz
2WZwAcDgiEGd/4nlNuIQmveYwEPMYAWpHGZR8/lA/4o2et+L1o43x+/G/zMRit4b
5inbQqrQcdocx9DB5YUWJK1SnU5RZCmnSj8k9yQki7DJKrU21U2CMnqY2GW2D9ZO
iDbKeK46eCMwQPFdgrAfZ+NOCCoo3bbDoJeqioNfbNSYGAgrOXPvQXoJszakbO/E
M86ShfoXUkB0EepHAOc1q4EGOt84pluT4+AvsC8OY+SfWORW75SzpJxpEAnqOAUe
QVJQD6W3bNGoo/btweM0Pod2Xv9wpAJyXXldR4MMu41gqZAts0L+Y4znsjpQWPDz
H5dkAqDGZBbCWcSRO4xuOgkuCgtU2shZLkV8DC7DepQsyDzazfbETyY8GvClh6n5
6vmL39I5ArNBYA3118G8ac8XBlQD3kT53sMzqk4qRIMczlMCWZiNR0RMjA4jLVnm
LrGv/bk9/D0/iCGbuVkNetsCS4UWgPKwYDLNlIGHtArw5FY96tx/izPHR6uZrPBL
SFmefSyU7IJhs2gvWx18OQFIyvI9Jr0UtyMk/ZZCJZDJZ/IYBTZG6JdfKi+d80wy
wxlQksUHH69x5suLNECtWdI4oZil5aZ+jxn6DAT5znyTvK0hZ8n8+9GXqGLReWqD
Ucb2w5eGkn6jJTpiuhoc04+en9xszAnnwdhaRY2sqtrVn+1S5NOqqAMkf7/SwnLp
I/ovadpeCaMv4VLjmypJ1J3ULsQFCBEEAl+t9i5LkzQzvXRDOqYYiLlhqwxzNaGn
R53uSoSMEVq2aqF3nKxG2m5Fd1EYw+nYp6S0dZweOtilFIUSvqoyeQqzDO37vwMg
U7JGI7Xouzcf07WEL+P1M5zAEi1s0/HfMSeBKxSTSueWPXbgHMq+OBjiNujnEBFh
nSuRFpM/kDZZGYJVUF2E4eumjyw4HP62AVX4QNND+5zvOSd+T15Pbm0e54PVogX9
n6Rwqb+i9ZlOtZ0UUv6B4lMuAzUyMtw3m++iUmJhbIbQngazodJFbj+nmcL7ZFmG
O4jUJq4GF3kNrbIZxD3iArWYP+ZcZB/622CfbwK3/EVWtfsqjwLaEA4pj8ePkodO
n5wHWvSOkXcdXLIAawVNRMMP873o3TYEVkvmNhJlO3Ptvalu/lu5BydRq7jp61Pn
0uy5zYf/oRIfj7rZGGog0s7tgUx0lI7uTizN3+3cplOs7HRJlXjnO/MewyYz5JDk
8GEufN99kivFa95axSLD/hEcGhAOh3NbXUjyxVcQu5uy/KJ5tOQRB/o0H9SZoMjm
YxKHl4Jj5KVD7GZxzZIxkIEmHXAy6IWE4kBruX73klKTtudGFbdZrC1U5aWkbvNG
L0WykMkdUkgVb/mhUT1DSc/iBo3ApQ/PiI9CKpvUMgdUOH3c6qVDFyzQtcwnAyx/
gX5jwj8JpcWV61zC+h6vtlqWrD8oEXPgwNOT79N3eGUJlwBnZFHqn8nrFly1fRsI
flTPm95N9uILIaVOf1I35fL+AhtRO0odg88iwYJVR+PVUcz0Udg3gDgdU2+zPa67
hCQshqAfX2v2mtkwGdncI7rOh2fIrtI+xkIHr5LgEU1yjYVENxzZcK2BB5uFvaKA
RzMyrHSjEJJlhj8uEYWomyjtkaG/2qHhAwBy8N2BAy40yq1tHR1QERB/A6CENlSK
RJ4rD47gg1MMDlUlr67seCkGSsXtw8Xcws5zS2s3gyGEnACt8FsJsBrnX7jHhJSy
BS+C96kizX40JoF+rSJGkfyCtcw7uos3QCPpDc+/AuGiQbYTkGWWDB6LpYI279+8
T1WmarbETxt090Rr773RiW+2S/gzfPgQmhxjsBEkCLgazmvyld6ukyoW67jAkGqI
vKn/btxFBUd/OEHJktoLykOB4mQQ0BucXs+oXrmoeZxhGaNnVcSZFCGnNBCWFhh0
RMnZogwnNm05oI0su6ScIi1c3I1ChH7OiJNYm3aFEWfZQ/f1zbG7az9JZyoImpGh
J9muZOr29vcELtzf1BA449e9DYCzw7Ng0ydxCXzrztHXZ2+dlGNWCJriTSykeGQS
+oDv4jU/2lVlGrUrud41FB3INuxDBZsO6uG9YcNxkSu8bfEpHXGXW/0UzfUjFZKk
isZApDlDW1yd+SLm6Ejvnf2cwR4gQm18SP569/kQMiInSy+ILdLEHY9QHa6ch4Gz
7iFhksjQtA30YHYDyTF9H9H5OJavJNP/tf700NdxGwaE/W1fMLNAQEt1Xi1jAfGw
3VE4PcQkwKYMRHejh+kV3chUA2LB0X/+yOc04tfpUr3XPIEmrGjckbxrj/wCt66R
ZVajJfJQ5chMaf8ZWGsiFbr48y999e5GS1LH1rWdCqN6ku4TGx+D2SjoK2vWGbgc
sKJvTGXnLD49wOs11n0PqBeH7GppkJbUiDZwdnfUrohuaBifcMkNU8WnjVq5Azhw
WCWpNgjf+1po+xKZzxRhOn+JHqK2+chTrJmLIpVhf5WgLz4yv2Q1sKt4efgyEc9r
GUXIm14x8bWEGidkiRUJpT+VWu8BNsTmBDJ5gNz48J98amOrI8DUrMtDVegJx1mX
Za5JFPQ+5b+0zCRQPrYPcyFTsaQ+WrH4AONOCskb3sshYQRLYnlNzSUpFNBz7iEj
QhwPrmTaDLgTcD6QZTgwS8n4Oy19K261wWxFAF1dK0kzdOZ1fLX6EAl9wNxrf2FI
W7AI05TtpOWaFYa5ymYzaCNkXChpcoX0dcnSE8ZUG++gSGV+69Hp6bA2xdWKWcFx
Zo8dpVG15dPU6NP9RBdmujdJ3tVmKkSWiO5ewFSgrJuX+2CHjwfXZx2RepeX2qP+
+Xfjf8f02Co0bFplO8kpdOJCFsylsbAnHsvE6DNRTnIYhKk7TKSfwV/9oVEWTYzO
Xoz/7KRkj2UGjycoGFuRlsczZosFikkExvbXIZATxBJ53jJT7r/z8CAVPF44DIpL
0iT9oyDdf/Toza/EEPZbj8wbDE2AcdeydGcgEmH45+rvqZLJG9qpr06wRcPSs36+
np+u6m/NTCBNMlrfPZu9THYE+9HILd4dBpBfWpZRz8ZHicG5BOJ8Z5jCQjYTvRv/
nrOGHbLkrPAlKXipIm2U00dUcZqwX6bCfMkqOwe/0t56MhGQ1tLv5mhsfvI8S1gb
KxqcP7BdRXLNwBd0HYwWW5j/kUAHF/aS50MlKoNZ28/ziOkmByE/f5u7ucS2Dwib
F8ZUOQ07or1K5fIF/ayiPKdfMzgQBOm6vXOBdKFHyBzAdE+Zkx3NR23klxjGGHsc
DDLzJcLTcRM6agYEbQgQ8YDCArfyWx1QBrsuDvo2sjKCRJNUoUE14J+m61GIUZqp
50FNA4yChHrRBLuONQNBFaZbZ1I8rhtxfvgSpaNQi4Os2VmgY/JoUuKa+4lQ3Ju2
kFUxp5C1lswqBnFO4f8ArnD13V34zJpd4V8TsTUyJECruZK7ovw6LLW6rKMqVGsK
7kD9CKsToChwffN9xBrRnfMNu8J48JQdPw/mQ5QyqfNi0wjg4pif/rO+NBrBcA3J
wze3L7L2NgngLpqCkoBvmsK2ByHHu6mdsID2fVGQgpeCC6JEdY5bcMU/47GuqiAT
gNXtaNoGOi51sjiBomJuF0124bsR7UXL2gcbKSu5CgY2NML6TQl5iaARw7zbdW8Q
MAhpnAw3FdKetfGwm5vHKmau4mlSLndBMeAfZ3wqfLx2ngSWsQfYylhvd2+kIYYw
aoBDC20goRMzmTPb3XkFrchD+MLVOFKm6HJBRoHggoDBt3V7gLoh94k9rOzRYw4X
1ieXrPAOZB/C+WMxiMqUlUIJ1g8ZYgpCR4cre+OHsfdJWhD2VcxqXllA1RR+1VJl
oSTjW2jzt1wVnI25SIklWJM6+Ob+8v8FWevHAn2PaRhqRUwuxdjnnHCZ8r3pAbW8
2BcPd3rnObF/rg3Ywvmzcs2sXq2Updb7ubgiMzGT+6v90/oLCVY98mHxW65ou+Qf
EdAoHy4LjdpV4LougbipO6/jmYvhOZn8Ro9JSRwgsl3aYuQnZmhBzx5/5rvAYRSW
13evNvCOaCMqwIdFReXliHNqteaWEd+opX4yV2lJB6F9J7oPR4bymb1O1GRMCgyo
lowvRmJwHg9GYQu+y1ebJnmsg4GXr0ukg2ACdSCKxndW+kDQkKZUyzcWivxVZDNA
8IUNSrGM1td9cg0cTsVxQX3PL8+d4nWQFdbt05sLoRcyPoym03IzBoo1i+pU2dh3
H+he5vstU2yl0z4AIFsRBDpMKWZHxMQrdvygv5I0gDdhQpNKQHSlellk3lBEmozz
KaQLHycgSvliAjAeonY6mvYWV5zOywt/S+1jDniv8Pg+1dU1jH7228pJnQ01GdZN
Rozc6okXvVG1Uk9y+dkv7s8cBsGKuhIIbVQPbQt2pAa/9Tc4eOrYcBKK7moGJrT5
TcQRJPs8WGZjZpYXAnq8sV1lAybEiGfEbChHXhv8TEhBb4ZCLwDB4sQzU3m+OPvW
SGMVk+irAjwed1wAClfyWlAUbRzm7UrQrc5YCzd/NRxyqV8XTRpQ/co5pe/OScEr
5huhfJAndEjLEOfIylalvWwwEspR/xIprDJPT3CGX29ezdcnnCTu9MxdbXBNwR0s
207GInQYe6ewJAntlfxh5R40nPMJfOThgzCi3FZGTyaFwHuM8NJly+5xHHTdZiKX
/exEytxMEJ12YopR6WnrdYO1STTsgm31rP0wBwZEwMFDlGn7V+/AREcuLuA+nRhn
1Bi9nRrsa7kSICs4Zh8vouKqcAhrMEGDqohDFdYMzwwWGv3pckeOaogWSmyPAzyv
PNxMc5doZMQclwfYTMVh1wdV1Ls+jw+DqZlUYyZ5G8e01MFuVsGHWr1mnDwHz296
1W53FBwhxWcAqnPSNuaSL81ktwx7jikIzm4ixL0yw+5UU7JjPebA1fZRc01sZ++Z
U7XQZLqC1kQVe/vL147dcvzmDlCCZtue1KUBygnwz7lwZ/RdHF9Nf92n+CcKBEfn
wcfpWd4G4sdwtVIWdehBxojvjUsem2NyeP8QtDFvIcXwv1tj3CFQ1IRXyCO9F9ob
K94EtSZnD/TQe+3r0WM67nyQdoXlho0TQCKQFY+LcgB8gWwgEgh3IlmQhN18BOFg
2nPNDgpwXdD6N1xQ5yV469lDGOSEiBtqsYlYPJ++FSL27YMCY8op5/uR3LMhtPKX
57J1fCueienOLl3NA/pdUB5ljVwQZzn1vu10pmviz1tiNGbfqYRao1pXnELhA4Ta
E2uLfNNXYYixmEcvgJSM6asyFbeKhdjxlzS201DYf0vFmyr+KgaN5896ZzXrIM5f
+qDBCEYw1Wg0uljTnnkZF2cl1qSwyzqNhXi2jRbmIiRTAv0q/54bIsgOERnJghCe
7EepnDXGPFEjMA9vRclAzEnEcM973UeUaA+Vc9wmUm7IDjpoG+2xMs6FEJJAWWg9
fxEKLR+tg/m2tX6IQYZl76wUjVSHgzShSqwkrAy4TLNVh3CDs8WzhpQe+f4hWm2b
Wya7g9+H4EsNvYKi3hNIFsfcpAOpR4sijUfPUyxuz4Hsjk9NhGv/dmB0XaMy91Pb
ENn6IDO4VqTj5Ke6/citihwdmdMCtAuFQsGsVXpSx1jss/g/QcIAxGT/NIRUWeB4
cVJIyFPHVk/M3UpuHJSqeNItd3PRehr/QKxRDwFaosbV8Dh3u7T9jP+nT8nPlI2/
BcxgIJHhU8SP3oSh4vFNkI4D9Yx6t+orbatCyOqJv3wW+BjUEJ8Aax0poVLvMcOH
G8TH86XCF+EF1gNW++KThRxCOvxhnU14gNPTrQuBdQePeOWZKrjr9qaID+ncJJcA
0bXO1+PK/yS2v2lYPhMDin++1ZXmo01DaPQt2n1IhaY0DTaMlvHlVOPcYYfwHeXd
nocIMRD0E0kHVXN2i+Eu4Gduefa+S//xf/ZNt0kKWzEAyhZnjn5AeM8uMPRQho+a
XEjD0EvpR/PNSlaYdia3QIjx2P4P8sOu5yfO3A4dCc3qMZGH50Cri+2ig+pnlyKp
Nmw2mMcS9QDTj5dN4xrBCaF5QjipCUbkTuFdwpw68tFe49X0RynoMCVuLi5SgBmW
ixIYJhYKoig6k0tdzkrHXxrRj4ayWlf7emqln7q2gkvel4IR0D/CCGyc8usXOsVx
ZMRx2I9c8yy9puSNaQDX7Ry4Tw+5zmexsKzYjXtBmXEa8r/jCrsVl/xO3Zem9C1y
fDnOzona6NbJi3zM4aboMYQp7Na1aVhOIzcyJSLTmoiqt5JtUBkTAvWpUXL0r3N4
2pLO2W5xiK0clhJOTl9L7k6bxJLg5qqY8Xo7L3yCbqzjRUv1h84F9aES25f6degI
AWsr4pqvQ2FYFlx+FpgNR83KolS27zTmumog9etetRmAqOFk0pF9DPoRZHCdugZT
Ri/1KP2x2vNI6CAWf0sozN1iN09UA6ddSK9UYsWuZHRiDdN1A/RSlTi5RgdBlJ7t
3eBv9LzukorvBNcbj52ZsKdbzDLZcIf4A7pmOqHltxhLLhNveSeguDaDvFG9P9zR
sEzKtUVF0JFPyxRdLC57TmtF79ERNd5Fl1hWRrN/xPBQYLyiOnPpSbaS01EdMxsh
wDB2dTxlnt3KMKVghRVberzbVOjVGbMITXWHZ42APHKhk8aH86P6qyet//1o4tHC
v+2rhJ9DRfGMz65nzYKqts14Iqeoj3N8g+sts7cse1WqNDNA4Inq6oXEM++oElxY
lsiWYBf/D21OwHBu6cYmADFC51nHWrCQZBctKBk4eO1FJVVX0lJkMmysvjB5LcMz
BDGWsEKdaL3OZmtXScriinL2CVeFYgTx2gXzvcavtpsEqygngAJnOiiLyV9ciMhG
wjgfaWa5DzyJIllmsyYsM1ciKSLXC2ysArZMHu6DQnhEUkckmEw0ji5+SepTQ7Qk
IkXQlKO3g3wiXflwSJGku0+vhko5zgUbebftPft53zQLrjD+L28clxaOc+ji1g8B
g+3xFFeUW9skgu+5kH9tOiQ0kK+HnjNTgZnqHQVnFyoSH80nus1W161lPEomIl9Z
D5ShHgD14A/mxoO+z5WkeOsW5wm5TTzesj7gm5wlSSpNKhSPzpNK4Mwt7jLxuXA8
7XFUsbwzxvcwj+n4hMB7vqOKYs5o1JGJa52TRpJvFxIJN9DxEKlM+jVNdPfSod6F
EVoLGMtvn6Kxl4hWW06Wn/zOZ78TqOaSSF/uJU0gEqbguLPQPsohnRb2jeIGCgWx
F4lxkiLDzPdaVSDuNEIuaMlX3wwE6hh+cy8UNGf+2sA8DGrqERSClVZm0QUA/1aG
RcylCHCwgmTc83LbZZSITYYfeIlRZHnjzQkluBlM1N7rtbqUraTGb26cnPtBrJxq
k4vOu29qVtvCT5fwcA2WOkHV3EfaP3opUeWP9vkgSvvlwfoRajpw/mhYSq79HlFN
zWMMQWWGKRQYbp91ZHM2iddxAjOUVaf2jyL85kXD3tRc0LmiPqfB4r6Wl9pl6rEs
Yl4mIgra0DnMczzWiSl6qWjDZjIli9BXtw5Vu0G4cy+DVARNWH5c9sIQ6zk/V46G
oQ8D8B64iHi82noAoGAW83NLBaq2VeMrzsb+Id4Q04LwM1zmd9VJRAObgJojX0TM
Fqt5zSZ+aPZuKcjdlDIcYni5vQO80mX0br0p2Q1q2yojAx2ylSWvMS0aJJp9w1Xt
NVedqVlVAYT5dR04oFKbjElQrDk2hPQgtn4NnwIw/YekServjik+c9RqD7BBKM0n
6OkA3rnIOqjDOCzeAwWmMxxOlriNxCj1zGUBE/w7olWMYNwoW5/tSJoUtA3yzxP5
hoyBb6+8kY0Oybgmfu+Dh5OSwn2Gyiqn3NkjJHiTePss8LOUQ9pxumJ9pt7zoVZ3
9gVYP4DXWyu0SEB/88oR0ufFA4O1bR+hmdCPInu363R3mcUZp2v4i3mrOng7McOH
6ZnD5/aCo34l820+5rqpukWezn7h44EdOpcwqcJ+PLmRRbqVrMS4PNTgYi/BJcA4
L4ru/yZNR8Cz6oIcwzdWiDqHKEdu9Zi45UUl/Ybon+ZG4y3UjmR053PX3J6UUoxQ
bnampUKi3Q25KaGQSUHWLUtdFRCxOkfhcZlchySuKgEbyKXPRsln3D5UijLQXval
/sKq9RK1uHwj7gFD4KUaUD6w69tPGZgt3g2lAKvGsMFKHLiuhTwZ2qEIwOVz3tcR
aKoK/R4TnPD2dOD8ll61hhGr2lzLfDgTbiOZlUUR0J96/Z3RZQNY3Jmpx6p+y666
KDxiwfzAgTTm0y8WoHX6j6ZaQRr0kxHeqIad9QdH8hkhh8yFSISBT0j0zn4eyYNb
lm4xyQnh4lBQ1ff/HeI3FlKx1Kj8K50pweauMPYCsLKiEGH2/+s4iTMS/choelBx
VuE7IRPQZWR9pAYEFgFgPTZqodjTdDYunsawhGeXDD8SDTgZwdA+KlUDKPC2IHUd
jA7NGxmnuKIhe/6l/Jqc180hMaXHSj3w+P2dwPV2webTUkfXW2qz/czfC8b57e8B
DttaLadTflixJOb9dDGiNZfPZaAqL5hA4qUcPOQKGeGDQpFRD8PAWaEQ+5I2z9uA
jEUI+kkNdweJT2iDZDpm+07z8xkSDkMKcDdkconzKa8pbhwbKPW4rpiUxoqVbEnG
vv8x8KdFrSURv37L4tTt9X56UbLOWS/BznoWQIg80Wl4psdm5xwIMI/qqm7VMqpo
Ly0/f5cPuCmiod+k9q/lapqFn2xRcjhKqSyUKgzGhQtvTrz8D2asxOv76SnwsNKO
W2zazKg64Y6/wwFhbNpMRbO3X2gZts9g/SPAEsbQoqUHF6SJgNhokYMIwLbUmXNO
XuTaCjDc5HzRlWOUEssPI1IwUainvRdzTMYxQpR34uPJgQF8ISQl5Pw0mZjP6Uoy
GKk3h+nwnd7SIDsCMpWvpbzasmpoVQEYZRQZZW6atPW1Muu19JQAMjcCyQDZxGxr
TW4Wo8/AoHzrqje342OWvCSAK4xSeu0kyC9TkGmj/Pdc4NsmRiHCpNvr/CnfFnH9
jPnGXE973xvxIfEXwY3G0kpf6QRxSCt69Zv6MoYepVabWoER1fLJITxiCI345KIP
jbWWhSB7DetguUiTpoAIo3+Yhnu2d8IDLCeMIcozm1qf8//2c+WLmwWZuydGSaLM
BBKSClp6UW0z9Z+l71nGbQxyto3Tvt5xjfqul37DnOLQ3+cmRwQgPSygApKATRH4
gvisKjYB2SQa3ZDHdoxGnQx+oN74juJ/KA2B1JjXAM3sKp47DEipuUJQsDhXjVNo
mVMXvo8Ivb8DElw9SdeNfESvJNjT5rQ9HdHF3GhRaRM2FnKHX/6C1jaPkxkhHlKP
hzzSE/xpA3SGkBDJftU5Ort4gj4rgwSJhV65Y21MCf9L/P8aQLXTCO/zjw0ot+sV
bfS52DorQuv0WVZE9dAmUyLZrLOMqMDAaL5yhZWzZj+JWJxfaWOWX2cPUrGvPn/a
iBmwgtOBuSm+h93or5ssc2iWxWovndl2vpMIq5vCmjGizNBQ6EJdAQI0l/C4c6Tc
LPkfZP/AWBZqxJ6se9k2Ho41JrdBdSUsxE42v4FsvSIL/BOMaxTEKB7lb2pKPl0d
ln+/5d/GBJaX+U9rRdIbvRY+oQsf3tphfrivc2rGnI+dRSQJWWUB7mbflBWIa/Yz
cuiW50O+bK0TTjWBFVhE+VM4/V0S59FCPPRFuVCpD4Mkha6j8e/BJc+Wn2BrsWjc
Gp1wb91F5n1PBd10MqjXOYEbRsbivCgNQ4WmGOyMYCnA9MH8enKMMXHYd/dByvSN
59zmd/e4jCCTeT7BSQdExUyZvAjAJKYAvoPZLu717a/J/9BWnxNTg02zdCW4MEW1
8+WKuL+ZCLrS1R6IPTcS/irF9nK9YfgdDBiRkmwGzM5+Rh8HKCJsdmdHUajp+z/b
v8RNXGq1V68G86DGD5tr43f39mPUeZno9Kd2IsH9p5cuuaWIaXh20jaiNyGsNtED
qDjiLxeLG37rOEZcu2tOyc9PuI3IPtRF0CZvfkNRlolmY7piztulYP/iTwaTqUYw
f+8HNiMJQadU8I8GpUC4wGN6zHa6EONIrCjxc2Q0xw9GITJps0z+erbAHSbwm+zY
mjje5e4R/pICNxdcQARC5cB8y3FSZ4u4x4sTpUXHfj//ZmiEy4+5T2/cByr6tG+Q
8psDdrH7vPWSbX8cS99mElCAcAnZYiVLoq/FVJ3XnFSyOJbDiN6bqzHBRI+grixY
eICfokSoRauqNtMhbZRMBAbLqLGVNGET8mYvWr5n0k/VaFrj5oeHn6bGUfNaBUL/
QGLq7wxQbSWKZcMP2kS5MGqt0AmU5uK7913CfU6AiuwoRlDm1H0+VVfrlClWj8c2
xaQ9bAIEKWEMnjPAIKKfnQqJ+59p6kkvGSTejOCtYhyZOWKw96Aw8WJoDf/546Hc
xRVe82DoRDcQaMDvStlIAutUA+BtWrzFH8wpV2VoxO+ch3DpTlzRe+9LJOkqbGp3
ndRkN5Bsz1pnk9X8XlbDMo7AVuKl7RR7Tcr2yz9uzrXMjF3Peo+WNyIrgDQ88FyK
5VctfXjmb9C1QvfODvitAGzpg31oOixi5ubLAxi6vD2cuXGWLDZHUo8uqnRb4+CC
EMxpMNrvunQK4OWpmsIuflJqL3SAN0gjdcdEhe9VEjbwubqJpFndbui3LaGNTRhE
F9fQJXToh0xNvjbMynQiEidTRYFun3VBpnR7zXXMy8wWkQkjKB+RxdD+lX44riI/
FO9wCdIPtrywf4CPvdYOO3/V5p41elbRA/h/jOEwgKjLeNzr9ii8n06sMDBqdlXX
I0sP2CldWf6X47Yt5r30ktY6hQF0DPzGKcAF5ZPSHBqVbqEyDR0eu2A0U4A6/hAt
L5keIz0cb9SyJ0/Sj8pwu7vlBxPIaEHYScfFN50TDOqfwTGjzRpVyL1wq7cSSHdb
rA70aWa6QGQEO73hmv/Ll8PhLgj28sgDeoRYsen2u/zMJGU1FdVrYNqHbqLdtB/l
nJ0mlMOKcBspSSwnWdl/2h7QNrkH9QQv/iASIGKfmdbXPvYmcdWk2YTOOo8v31nG
cyTNecczD4v/g0S6QNfMmPoOvvMcoHfSuPgpOfPtDyM1jEm5Tc4b5J7hAjkFusHd
JNNKmcpT7/e1ast3UWpKofjYG+/IhT2G8w6YM1Vnkpn6tZ983qf7wNXfO64ZwuP1
0p3xkQEw2a1rRv5uzXRVH943/sSZb2A9i+9Ay1S9Ebp4/R09K82Nfsf1xUqQqe3w
GGvlwHA1gaA9pb6H/9FF9MO0qmPBBSCPth3oVh3Rl7OunW776mupNsWfXmxROdMz
84SLhaMGIYRISkf7mcNs9JSCRrY/KxIOMs8xw95vxV1DAJ5hqfvLcvd7cu31xxXs
K4ecr6Z7aPJGrwDFav+KmiRhqlV9g5hLKWbFBhn787Zuzs+Hpx0UoiteLWgtqAv+
M+Y/P1OPo+mTsYJFtqTdtbUpYvr8mG32I1K1gOoQJ9KH3UDb/3W3ktbYo/tlJuPb
hPmgNTBWTdDDAwJcRjZGnoClwg6l3VCo1kDtd/AQhTzmlzMZxnGQbWfdDZFOoaPJ
tPU5hZh+ebEeXHsyazKMVI8nnis15o86HZG4Bt7GpSsz0ISEuNKj8Khrhq4hmSWK
+j5qK0QMZIgS7kA66poYcOUWRKaAllwgLGb1ieAo3jv1duXs3FM32W3u7WoCN05K
AMiXW9TrA/BrWyDPXpRUtLndHgrylOud1lo9k7TQEpm+as9dAkfZAIueJAyNKxpd
DD0PUTTHDBwwbnrteJluRsvcqbCIsuysQUSLaf0YF0UVoQSyUhrBL3ZxpNRvZXmI
iVJBAarDe9ShHlcCdRx08sRdZ0rWmBNQHd1Ph9VQj/1zUb+cof76/CTkkijGx/fu
FIsXwy2Bru16p1wpF9MP+lnYlbAajBeC7LNiWv4miE9MvhYbnUbqDK2V2rPBsGMq
jNX0Tty5JCqlxi/RM58Mb7z9Jq8gcfcXX3yalgZBfHU4ivdm6qoy6k1E3r7G8SmN
+jeO3praBA6k++P0+ffodKUbYXmuUgXGq7kefgw0/vpp7bIPGQCOn5XJsYDm78+B
te/LzAP/a5Gn0np1SQEpVcx3LAtmqe1PJXMCvx/4YdFyNOPLML0ztmSMWAknpImc
B+R/9+KqLNLPtIerpjlgivxAtnqbMPlcbLXBtVa0cnzPLjzXlDLTPDvYr/0pzeUY
0X/r/oeBOSL7bnU5OYk82C2dQCbdIZDYyKGSRJimYhF8Ul4RTL2JbmSqUs+amgqx
yZlQhXAOqllmIw/bM0HMvWIucU4tyVttkoXyBB4yt2Wbp+2iCWMzReuEIrdj/BAS
eKADdN4zce/ignJcfHD19w71L/gAxrZMYZ2vEsEUSKUzxCz8FvwdkTW3Rppe91v2
uznfmhPizoj+F7EDXhxrxtaPyNuBZwSM/2K8PNPCyFGrNDquE35ZVaJ4Fd5l9JeV
W3W/armG6azzi11MsQGryiAoxiD9UCnHyctieRKxv/bxV+bSMivVIFE48qmwhCmb
hB8d96IsCKWnzuEQZcRjQYgXNzAS/sj+JnPjLVfHVpr4YwpctmSONVsaX6KUuaD9
lOfONj27LYi/hZUCGa0J0gj1aRxr0RUwNvP6zacz5la3y/Qk36vvP2+YZp7Z/Svp
GY9RKTy6+mWdV25H7xBl87wvCIgjPq/t2ZPG0x444nLgemIXaSc+rejYLq6/YCyy
VURxUUs++JcPxCKWyznSxlkDPeeQHw4QMypt9yWvjd3PBOnoHVzplckng85RKciu
xT8RZz9N/iYaKlP6cZ2eNOG7RNrlynhVRenUZScdVtvI3/CTX9GiQ+TpCLnTZ8qH
CAAvE6gS0mpM834d4Z/BYrXiIr096qy8rvefiPpk/aXsD9k4dy+PcH1DHl/bdJFa
jKrKc2L02anMsdJbp0ZlvUDry01yThfzCi5vr/R5lu+TdZwtP9HIglEMPZ1s+uJ2
RjkgffI/cP9esaIKIeWfG9qCE0ILnj7nRjo6CKoGFsuxfJiKkeaXaQvPR5xaHvUk
VW9hzYIKMJr334b8FEXIFymr3Lk8FEWaMRMtitDt7XhdPc2ktPu8Z24uk80kSj+A
3ykWJ42o+Pg/gZZx+IIF2f8DbltJex6H99jluUfeIAGsHHnJXwe7qvbQ7OtUilhX
gIzMCZxkVCbvbXUPaHDqQxflANQR0vDGdFFV6gJngczv3Y35xvsLiK7Z27OUmDE2
2bxkBUeF5qze1b3aoY46v5D+NdCpnwd/+IT6bUTe+OqpxFt+bOdtxSMy9VMhAoQj
KPFIABWDG3s7UvMHQHj8UZU2A7DjgDjFsY2WX/EgjNEu/4pxA9u7dBAPITw1QYuu
VBTOp/+QgC624cBZ2iYzVfPoJT84JFb8E2e793SNt7fQqNc+Eq9iKxxKTCe+JPK1
aQsEAOezkCi9QHANOPjWyFZ05mlXyLk3vSsQwOaA4owlPjfJfj/AAVkq/x7PN02E
u1qYn4R2qmHXb+vQZSvjKp7uu1lor7Q2HldtXwG28HUg52nBChgEHEbKKCRjm+ZU
BByUhl+mDlozo+hndICs+DBGjuNsT/66R3/DM/tSQ16b/FjmbBTvSXkBpVcs4O8n
FPyQH7InhXh202L/RZ5DObRpkOqj5o7QBuaiGijKtjQTRveseVfgomN19u3oYUj5
xkuWTIiEsV8ecKJninKDj5nOqV+reNdMPoCWuJZPui1SdSdScMq+lI33BLu9tWuV
55SCO36tB5tFpsZCMjQsQmL3tJHWZimWH5Noo29BCXOaWVXR4PIRN4rzva61PkOs
jdn/FSu91pO8rNrAB3TIAErb2BC0vWL65WEQ42X7QdZgBWBW0BHw0F8vL5zmDmtK
8vVmVnSRoPFY7oqZeZ1tIt63IU5zUCihKOt479pK0qRVpudFmZItZ4Kinw8dod4o
aEtxONpP+wYFlHljHtwDwk7DjnKG/VQHJiX6SbSfjoBACFsUQaRTUXvyGDTFiJAG
BPIyC3v//Rd5RL5CTVzdmRyHBnK5BgQQxFGkNdAHRvfSi3hSKLxIzTLfVxsocdKX
+PAENeHguVmPvumfYmsTlTI2hzjRmsEjBOAnoPbCEAbR27oGt92D70E/2m+3U6/r
FcGIHMgX7m8DMSasYgjl7WGZP4U2vq9J2ll4TNj0j2PSL3QXyCTx5Z5HIcNBv+wG
LAPBiNUwsnYQqHRvGZXUzkn8vVPYfB9lc5dnW6goSjnTiQKcuCX6rlZu7a0U8BXE
Anujk2ewh/20wBK9tj5etqj5oGCOIQZEnBRK8xUjSs9cQvXRQbg1vfBSFAK6qNda
2ZscTF0+S2UB2ZkVDyvrYtN7EQnKg8NsK8k5z4O+SG59yp3ydulz3lxOY2ROIbRq
OQAln2+JmkMuxgUITThfl0gZgzdUuDjp8jKAZAsHXEJCECpAkFFJ2pxK88Cv5nN/
a204ZCEVKi/Q3o8WUs9NrZ5gArRQsQKp2x2fRGYgSmPsrMUmDSsuZIuEP5V7H44N
3YhbtuB6m4LM9HAqzqwmuWHJ36lkHj1ezKWpVT7O+MuLD/5OljsdYLyq2AfcvuLu
6lTDDEjCnbEiK4qvEVH5dU2MqjYPRJMuVzoHKBxdIxaJpZQkX4tLSxJ5Nvfc0M2F
/Pobi7FoygfQkIN+5UbwHqnIoFPrjuci1Gt9o313Z6Mjo1Rt5ZFTSo6PSjIVyarf
GnI/l9YiYTT1hWuoN3r6hxrcGoDW1g+wz2KNLHVP+xQB+RDf9rRiLRvY8b7U76q1
nHu3Nf91HpLYKNcBQp+frO14H6Lw6HY013sORFjEbksu4UFY8m0beupDU3BZluBj
xhf1fSqdxNn6dAyDB4p9GLS0ZOQS1AsNA3lH/b5oPYuL44H/vgfpVNlNk9N+Pn2W
mbtFvZaYgKQpABGTwlk5Ti6tbAiE9M1RbqwFyCHTVmiurCFzm/1MqOdLook9t3w1
Ncv0ccbVLsXLLLcSRRX9svY48GjW0wNX1MohdkWAhTS19HTnfc4+nyftHvsdTVuQ
/F9XUCi9WuvVGqx1sY3NMw678xOZA/oHiCQ6nMwGzgeqUQN8ufCBhwMVc5Q44Tut
HuVKdkxVtOmyVTpNFiprrP0RtVCH1CcFc2sgTDX5qRwNdLUAIlLfHBDfxWpSIBEI
KRue7VWhVpiSgORzQgOkKkrZHRLvSi9azT3KWmUwBABXtbTxVWZqjY8PZVIBpRDX
6txGXbPJWQ2mJTc6GXQZW6JwseYawN4DnA0DkOW/SqAGdIGqnaM4aHsapZ2wQrYe
cbFllyo3+2bGw2+TOWuIBqAHMu+sAn0nvdNNzo9QKilB6hKVyp9FUl3oqZixvxXw
4VSzqvQxi7YwZ60YgIWgh1mv75ap8yFjpXHr8ojwZIWqHfFnyEwdECMtYWj7Tyrm
VNTs0sKK+7EfoeZA4ybenA2uGQLAVRMxagGz4D5fhLomBrJTLOVDV8RGV7lXmajp
Z1seT4PMfN06qtt65q1jUOSyMlx1eZhKRUeNlaDGfRsZjR8QybgbwJgX/zuNIZ91
R2ytrXrkSSkAfZQsgv8O9zv/oeXAJZIf+rMjuwjU0oCHWg0hwHua/HBY1tKLmSol
o4SfPbLnMWH5hTE9YuGPUYsCYettg3feibsk4+4xy3tu6bY3Yxv1ZGTx1ccG1ErQ
1WKMqnLgGaxRk9id3s+EzXKh/0z3P9ltOaEWQLM0oOObddL2ph4oCvOw/za57xPP
+cNJ8ds0j+AfDdPtK569Ucu7Mbgd0aUqOK5AW6PoHcdQtGKGz0gQRPnj+qX0v7vP
tvSYQ4Va9MLWVqpYhPlNUT9v4Ta8ltwGQTGUdCQJRN9bdEbF8JjJxZw5qie0IjOR
XPwEaMxfdRMHtt0JOt/OElo3TKfRzgCWONJXFVV8iSXp5aEAju1OJ+oNcZ/YN9XJ
64l0aF/NRUPVRa65nwAfMM+eix33r4DkdJWJk2549YV1IoMp1K8e+X2M5JdqC6w6
jRSeMAYyonYtSs0O1TcqrufAi3sPIQT0JWuMGfcKP/YcyybIydUACOXyzVr23WtP
StIwjhd7tIuiI+aYvs5bBDTLFvgtqgAKIkOx2YJDFLQSYhj1mnxvE40joWbikyTG
GHMxjNkGEYbi4kWK9+4MtcNq7EnwGP1KbFrtHAknZX70qKi1aTOZXDMlpyiWbjvo
zSJk9hI+o5ABsOVGgCIX/1uYnsc4WDQwjFX46w70+dnVvKO5P031s9fmoPt/onvD
dfy8AR2rrkPavLSLGH0i4R1stH7kOab4NfVLMpGksrFE+hygm5xzBwrcRavgBnpx
l1QdLdyWw207pX1IFOi+0SpDlnQSg8b1DB17pCk3+s0pfcEO2pFZg2rmYISfyMJO
md6L1N75oJC62wlF9hqKX5Vyn/sFg2utrgSfjBTECwM6eDTlwkNcTIOga09diO6L
sowYWuErgUfIuK55+b/knTkFP2w0F4tq7u/kZ6zFMK+ZX4IAGfeysbFXJ6gEkeyC
NFhDtQ3yG/9Rfk2EwylUFvvpWCA5cn0wsYeSkgRYNfYfvxLymaOwzGlDCqrSja1J
ef+vLSxjVqWGA/xpA4tSupzgdkz3mZjnw9dlXzGFE9aw3yaiu9+engOm8odTZTBb
K+qwdsViawMUWLhhK71d15yMHuBOSXkHv+FkRjUzAdMLLQ+AWHzT5zOr8YV8dOrB
z9n7lZU2bGCF+hGmKNbps+QRTS2Ld246TnxWD+23GneoD6QNQU+2M/UIHPa3cD1b
CpWlvT/TrEhFLpUsCA04FwsQSOvrSR2OZwUBSpm+1jWViGL7jxqkhzTdqyq/ymMZ
uIhYPCBH3reDtlzw43r39ECkjQvv4OH5lAq6yVg1oM36HNx1/1rq9JEv3pr2u0cg
4/xfePBY30uIjoWn7h4VCXheWaAUaPJ9Z+23ujjmWzdABmQMsAxIKC/3ABn8XK0D
RNFNi/Hsvif/MXxpb0nGkNbq5A6UcPazuTuDxbptl4pZm8sXk5BY+8xoE8kjEZcY
KtKOG9h3by1KQ2fsfvx/s9mT5snnRjLL4SuUTu6gPJIhwGBXVFCtNPaAkOnEXdBW
YljUL0/7lpq5jX+irvz0TmhKRWW13JGQ2ghTBwqMcORsrE17KBGv/ZyK/eICx7j8
a6z29nna+cD/M1yhDDms6DBIFSGDTkDTWbALZYfcZhtIddSDRpN0B/Pywhj8qaW6
PZcBwNstuUuU/giXTVG7Tcqe7aMFQP6e5X0zx4L3U9q0XnPtbW4mlXopBLYEWyoB
JUhwXL75Cjr9zJ3SnzEvHY3g+Jchknm77/1qs0k1VFk7sfBp6pqpJq6Eo72D9+pO
E9RAkyGcS6IpPDp5b4nBCnH44eIZkHGJ1zO2XZ9MkLKJzVTwfkOWqMcPJW8/enoQ
CAbiGsxTWlxmcNmhXUhM4/NPq/ewIqAWnfnXrYorq+Yd+4SBXcrn06S2EhDNs38o
oIC+IQ2pOQdvJ1WOFDLQxBaGE9fPmYtRRDBhtKgIsPP5elHdgeh0tyOOpnrUKP4c
xkXdvUDV3tqG8N1BtmgXRO76+15Sz6wRPt4im8PFXXU07+cAZF23KvnK0LHciLDI
n0Hhfz4RBSO2bWjGScqoVYONHcnRZd40qMUwXduvJNNEwwh7cGyPEtSk6vPaC07p
KJU19vYuNQoTxyhyJJyZ2WuS/mPAxEVABi323kfeiiM8J38jKZIUpc43UEdXvRjp
iAY139zE3Xt2qGgjXZ0lmvszoM4PRFd5D4SIKer1EwxzKdeQmpCHYfrd/ZRAjhaO
RsNH/ZBX2ceA4bE51tllpYl4AfI9C6Z6l17wCo9D8w1OgUS1kqOtw7Hz97Wlrph/
8mb9AVmBHAT8V/wp2RqouwUQFpRqkKdc4C+7ejL6csRjSpR+05qA73cdvHDrdJVc
t/xoCisf4Hf2WunPQ/bTpGKkXJPGxU3OLpCKYnHVafZ1W+G7CXo9M3gtYKFIzRQf
5Tb/4E45cASu6kb4nqgvqkmWQY1kEBrKmsFEWTOzT8tntILFT2jlX4ErnvoENyBy
ueanlZEa8T8kxcjDxMQU5B4but8qi+C8F3Tibpz2bTM4aAWMCx2rLtuD+SzygW8j
3aqpKbqOHFzSuL5IJOA+Yojfr8kWby1JRIg03J1U52vPxgDE+rNOFAOccjNZ7tg6
zQcO9FyoGgpCbKEkCTYDGMvNlN3S4/jThKCB8XWDOuKyF3zNK1CRaMWRMyxWcr5h
i8WPCl5NX7diND3ffYStDcRxsUYyEVcQRvlKY6X7KBV9u5ln8bcVAcV4mFwvLwED
xKIQgTIoYYGlq1pIa4YCKUgcx6FcWtTyzOWQnAb+uN3/r7TU3XKSfGdRIJ3+qnCV
Q9z6MJkZ9QZ81fhFwY5ogWSocIeKltPz3VXLsNjBFJj1wRGD3Ogg5xOykCZXfRbx
e1lmoAgbkUl2uKdEpXBuNxZIbKCbEwTZP/CcEerGqwcYl/6OsW1quPwp91TLlwBW
MlP19SfYWFiY4B9WsIwVJXq6i2IxHC4vuVQnP0XuYeuuJb03Fw6rDF/3I8hlLHXe
/tdA6XsiG5rUJr+w0Cq4IU24dcMLchQbA8V8zykByk4wux7cIDkxhTRTP7/TVtEa
o8t8ooMv2zmz5lixsOiVM3RDf9AN+04NLMVdI/hO8Q/KmScrUfry7evyHVidWMLQ
aWKxl6rDdg3N8KKQvKIGE69Errm/vefeE7gTcbATqbFW60ehck+LBr9WnVvJ6AIs
mRYO7v3yM7VaTnCbT3itI2KCCcmSig5mdJqR/5wM+/51lZjxt/1UbEGHrag8+Xdo
mXl+8IYQpHg/aAXaQxJS2y/3hvxeSVEPYo2f5cs9GYbHASzGqLaG4RlKctIIOWQf
ERVWr6h+c33g4aZWXszEmaASiQm3+TP0G6Et6fetVxbuRERSai5Vu41+nZbod1D0
TziqLixbiEnD0WbWiVDYuprpy2Gb56o+Zc6j4EEeSI51NwJCD3+tb5POmd/LAqET
o/dNcrY+DN2n3kpno7g9ml1L2LYf4OhmLZJUXchE8Bm8HZwLuJE0kEEEXjo6dEL9
Eo/484qZGuImFKDaONbzWgW67uBMHDwVIZpvzawZu3cntT40u49rUsADedmvXt1l
2iDW0EXhE2GkdwN02VXrxy3yzg9kLHNde2pzGCeCTjZofISJSyU4te6wofrpUGLI
UsMl7/0HXbWBispiOZ75zK88gSoQgFnwwH/q7DlOkZFOY0vCyAm8h0yhLgRUte4x
PaSkPHW2BGWHxVXrGImomFJybt/++9MVyyd2Y/K03KjOf+NXWWw5Y/mLI+8Yrp0z
r4u86baaJjwtzolxapoS1O74Zd9KcJjFnbOqX2ENGR4Ht8b3auUQ+kYzqMhFWGyS
ODAsETEn3loW/C57lhCDZfYeZ5wc1jDjLoYaSyoEO37498AMrV53G5GLhAx1IsHK
t6eNZbc1ZTNttgPnF/4r6FMcALImmnaOnLZt1/WB6vkPwHDlZjyeh/1/4cW+8uzO
KVaCbjlgQfK0AY+QY/daDOjdAXHlfX1/NI6c5jdf+8xhlJmq7r8jEJGBW48my2W1
uWv38XN8AXf9dFleFwmjFKh5/D+dIWnmcnsL17ZwISZx7ut1tMU3I2kfiN3GTo++
2AzZ3hTzR+eCkqE7Ix/xFgG4UJR8Ugl+rjmf/IQAnqlXEQSK+vI2/OMrHaxzfbLZ
Kww91WPYagexwUInzFuuLScES1SEiyQ+ZA+fUEb++i/gfKszdTJet2M+p7f0OooD
nz+6X5RwDucBNF4jIfJjcKfvZsWiKfVbmVWgOACYDznLsj/rAt1XicLlV4ROzIN0
XmxS5fH3Th+ryVP3LY7hBhI4tW2kzWtZkyh6kr9++39ZV1MlPXdT411RKGVDp3Rs
DuAx+Mc9KWS8KCqWmyuJr6WwGK10bye/YYJ3HOO7K6H39X51rBhtkvVITyDHRcGg
ojxpdVGYPvVy9uV8fLmzddIRtuWwRUy3vRyyYBy74XzTf8y2NEVDhgmhFFNT7mI8
e/x0aPyTMAt6nKPEKmYvb67rU4eSIc1GE8AwIECKbcj6hKUnPCWm+7Ta2G2r8wF2
+bMbY27vSEwc1XukzsB7LGh17VkxVfwdliQRNt7z42Tcq/zCYjUjtrrwxWbSmFfR
4eygiGd27U/qyBS4VD45IjSJwhNX2nHmej8DE4NbACqMpd2GGYdHzy7XEzgPxb0E
pF1QjCrx39Ntb6fWy7kmJh5d64mrUMkpiONzoYoLSETERibjRvcKHjXaNLI3rsqN
TT79spUeEWjTXAMdlqx3cjVlbDu39xBky0skzOuEBRbv73RE1hf9OOd1RwO6vyiE
ECPHnO+YNJ3wFFE8zXqntfl32aFFox64IGwQl2sP+j8mSqoXud58Q/YeTUXf/+4C
HEFGqFHhnC3mFMU2tbDxKbSKNpYU3XMu9wCrzs5SAl4pMFzDAzIQKWLdiIAG6z9o
24cC3M1MOUT873zbBhvUlQuYesCfHSkeBvvmaUJPHK7Fyuweorj6Ms7bpu8Ak0kG
7Tus///JhacLDbPiZ7dth6pzGJsktw8ins/2jP81tM+vz3trRziHtt6mikyQMHB4
x8fUnQdBQDdloQVmwhB2QTLWuc6JZ5vEJOk9X+faK8kVP7GTyhif46jujoPk7N+6
O4iZKbJvLl94iQIn9iHmfkwAjllnDmGB3mITXEsKxDEZVbI1DDP/JucuHC0W6FHu
VbAz51OTqjAvb/LqksY4ACOWi4wS4gmFmfoHd/5pZwV92e0MritaJh59hxQ8hSYt
v5PztI6ZIfSVtzDSl3HvrEBwFsfZ3MPXZ2maVWZaM3/Pdq6SqYhdaNetEM3Ow1oU
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
DFjG3HCDoGcflUs/wVlndelckFVug4LU4+vpxel84cDYe3UWqg1mXmVFh/GkzSQl
mMKuwrsMxB7PqDXhCEsifNfpyZ2Hid2MKOXDDj7c7tBiN1IEbXbMI440L8HYITFg
p3rdwlxu8tKzZG06FNvXbaXQLnWs+oXDsQKQC6g7hhFH1pN02YKvNgskWLiTNsp0
q93/Pu765+8rIz2dzW0Cb5ogEt6wx05dgZCYuhnU4JPWP/2Gza5XXAC1WQPr6n8W
blC5Oc+Vj0lkRaKkI6NrxCkPCBrvfL2GWbvSV1eYzqNNj1SqF/yzTZw2r/tEXGy/
4cxlBuOoBvTXU6xpYPHnaA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6496 )
`pragma protect data_block
2+chGmEFZ7mn1aU2aM8oQStXG50qy8D+7D+qcmRwHP5yBi2CT9SdUggGl3F/lFKT
BFCNVyNX38YI8qq3tZjwvhAv2//gxnxnRa4ZKQOtnsDN/j5RxtOTGHCinHsimwxK
Blz6DvbOHhGQNarc6l7TaSwYRaNTFNhUEAgIYM9nQTr1JdJJaGdaR0nIJhULOJDU
hved5np3x1FzhikPIxPCEAXlg0VLxv7Gl8vAC/zQVQ0Fwwuyj1vIbm1j63bY2kdi
hjRA8x5qE1rXC37v7uaPuZ75f0Vyr2msg90xcz07ZcfsxPVfTNutSTX7HkeQ7CkB
HjUfvmAYFpqhZSQOZUGtGu51P312QNAc6Q8DzuhY2ACEdmpz1tw6YJcwl+vmH8zN
YzhMjUBGTXRy3oT5eJhIhgsqK9PYmctfb/Yq9Qs/prsocKj39Qc6qeEVIxugkknW
PIiFX/gZPmwbTICJ4I2IWjQ/ioBDodMcE/XBKL/koTXHfopKrbLNCRLYqXpcA2eH
5RxjVaFj+6RgLGVC0lSh8ep+uC4WP2oB9rePvA0UbsKGrrrl/VEqorQvyRSNn9Fz
pt4QOEcVmuDAcFUfs23dPDD/TLfrGzc96U61LhGAq1skpXLSfeR4dKUfshjPrAJi
xZE/pQ0xKl6iiMuCxLmmZ9A0tbv+iTLpZtxb9Eep8NiXdyMZsuAju6T3j8ydpTXr
D2TJ42C3X3gZoh2Pe3CxmPfngX9E+T/ZB9kWvBvx+yQWbe6FNg0SygcZnkl/MNgY
6BDXaAvuf2okU2XdncSQJYNZV83U9NLTSBDaetEpRxjRWoMMbNKnkvupK7DX9HO2
wI6Ie6teTiDvZSeFmeLDLEcj43ITAKNYKouc7dWQsWswPPHEohJl6LfKYi/Eua3I
HiMadNW+HuhMKuW0ye8LYGklbBnFe+4rvZZUJp/mJSzGs8QKGTPvE61kZreHLo/4
a4I6PcmysqDtgCy/nSSbynCj+uFoNr7GFVCrqVi+B27gr8XG1y6iESZfTjcpvM6U
rFfputwqngr3OsTsxjZnJ/srK+H8uq9TNKDYsSxDMw6VbKwXbbML694JfUytzS66
zBLl+4t7hATkRJ2M9AgqM2i2mDYdgXqGkiNNskLeIkCk169NP2b5tWu3/A1OImX3
mcbHdSrIiZisFdiI31gUyuotZJjoyNv6gVLWN9BVxuiHoZkoVzAmIg+/R37CXNU9
VS3F/FcoC0g9WkTGnvS1KlXBBZilpMAOV6exFVDfbXqNB+oOUtvgG6uPDExOAGBx
C57TiFbQvPriOG3WSukadKq7J1SvodUpTB7C5OkVnH3Znol+mZoAVu/rh7cmXuTp
gSC+CqrRq0V8hJU8CG4STds3fnGYNitzRzDng56YN0ULu083Sng4YRyNbggr2uZu
JB+SXhi4NaMndQo41x9aWsjX3Wo3egbeF6339wuLDqiQOT0MDYRWEvBhqG9Ur/sW
xILYgPlTKuFO067Vd6HupeGtPCfH+IYdeYjzUYhf1tB+CDa/dUlFQw4Fne5vdESf
wEyhvJwXOANkfqRpjEgf7ex+xPka4n9BznHByr0edQqJ+SVPHlEMSbI+P9/1oCPG
QxHNrKr/Vg2OBso7FZb9CGOU11E08IZ52zoHVnkdeoD3F0VG1G3QqkxDHKuIxAs+
ZiUbomf6K0gYJyVcGJ6sP4LwRDqfrzTGxiWSq300jVtmH+eOcqDmttJOKkwNP38H
ZwqSaKjCAg3vf/y0BJr2zGbYeVUAxfsMADjLb1vOOiFeu5PmM0KBwFnSfL7wtQst
VeTXBbSf2C+k7XT6vz566osrMnuSR8yaXHP0T2BIUJJukA/yWzUKqFsv8bSJ4e3X
Y5dA9ynI2NgzoT9dzWi9dXzLCpw3nA1prfvI4ROkOOtXquWhBjUJkiSBS/dlJS5e
He3JJLLmu7fnEDCL37FVTSAHuhm7zcMlZgJAaJEKVfmtKePD5qOXzLd7zgpVyPdW
+izIIOo9ncJygMaUz+CZJXD92afxWp6e6DbknSL5SfAswVvKNcSIs1PRQwJ7TA2J
vqn5qOnJAeNj+PuWZ2ZVw9gRF/5uga1FLU6iQkXPRJ/IDBsbT7AqxW48S0MF7FkS
/gDMTo/RijdF19nSN9CoOVp9ItlRVT60CFJSpR0fTmQYfBsTdafZ/4XgQOJ7SRPB
1r7vPPELtP5k0qSVmJGQ5rULnmqkogREpRkxZcinzzJp4fpcI3K27VrooxUoGcwh
+cmw9C4I1MFUQwxHD/LNw0tlK60gkC5iAMC3UT0k04Eqmd5jo38DqSsxNnzdDUJz
Gx3nOxV+cdD8x7cX4ghBA1RrzAEIQBFYQcJBs8cPoHDJxiUyxfkPGzhATKdtEEYY
mvxvxMzKVOEW3ExPhY8jJBTas6yoAZ4ShXGuF/S2ouy30KX58DMBWPpXpZ4IKOUL
0PS3Tm5ePXjSG6JjVQ4MazfEBm5eBqq0cHv8+83zxU/fX/GU70G4ZRC5oUr19TYA
p0anuUHoOlh49k5ADJK1UVj+yaOBPtnOBYAberGXalIxp9lXKfTkaiqo2ThEnORc
YiuXnKqk5ALK95tCefoh7awqLoFo5YJpKMvYbF6xAt/8jIOfiItfKfloniPfn69A
meUriitjBRW4Hzq3ppZ5oAS5Caj4QraxywC1tLN7+ZxQdG7rdFOqfyRaaW+RcxEj
hVVXU1QjKaClReaI05nNag3bE1z5ChmXBW7BiWYACjBJzbIuCaFxojevGGcRRnAV
f34XHL5SwEZKInuKA1qY4+nV6GRnpkduq2WOUhHKw+zjEJSAhEtTQIWpG3bCHs3D
Z7G0wgjy0S1xxaCYkgS4FJLe8mlklqjqb0hc4Tdh3hh54TvRDRx9gCvFKw1q+NdJ
JsgWzDbgbLnreoFl3/H0vJyTicE9+dm2ChvZ4xpOt4KIPMJWkhVHKKgSrBbwb8N7
NCOsXDFGktHg9u3JNBuLS1OHGvmLXVptUS/jGwCHifNPA5zBf/eE3OJ1gR3RLYwk
T3/lQXoFYPvH4GI/3aCXIl1Nk9LCvXS04rLRkYBElLOBrSb2Ab4WOSZ2Y0KCgoJj
Msr862FD8qZkhO2NcxTXXA6EV6zDHnY39PP2dKv2XAno/rBLiT4b9mvfvMV0rJTs
zWjIbYTWMY4xPI2/RC7lbhTCfLD4e8XZvFc6adkT2uQrSiaDn/gb2lqmCTOXCbHU
QTiiNSqDwkbOcvVUbmNVUee3UwMUsrlUOqm0VbYCKMU5wAPL0ROR0QSqG0S6U68N
s1hWNeh9z/DYMJdTmJdSILzwCI8+vvhhndNqkAGzSSuXIe8PdIBBhng5XCiqzX8p
hzJTCVRzOT1dHnihgdePIpf17UaNCoE1HqJUYRfsurvGyCSZHm8HtDhvFdlbWSrt
M78n+Yd8RtNPb1yv8J4hFw1VZMAz6A7ZX5VBF2kKNQ7rzNvLz5A31CEHnW4OhZWO
LMfne1nNMaeLCbG7rq836ebni8F+ipogS7/13+bGUXwocg3EjT4Sk/Z2PGyvkQFG
jSr5yWqjMFwPmFr/KjMqPT/31Yg+Keez7bGUrrBbFII+wxpVEdfDUz9O3KY4VpDj
scIojls1lGYj8du/MoS8kC2W/eXIBO45fBnF/aPcrqDZz2k2aXTw5TCUFSiv3z2C
P8CZqCXFBQQ07/QUdbe+qmejzChztJbSjqjdiyAeApJKwOvNnn9eh3XKNHxSIccX
G3XMps+leFR9mkxRH6JZXyXZvI8VWm1Hq7Bday0wa/uihY36ABSJ7QX5mg3tO/R4
rf8JYDHTr2ZTYf790FBTTB3KMwN9N9n4hHxn2KVL3PC4Ybqc7aqzCgT65UbSyVnu
Ah4uz+KC1YIsAiWjNWWfOe/WAwobOv9x3mp+T4OLBBcXrBHBTD4ymyL3rHiNAE31
Cg7cSEQ0immJ36vWC1rn6PdXZcdSVcTCgdEx16XA+AJo8AD1kyJOqG48O5xg26dZ
Zkcs08W2EoxhGKvNKsYStPtswoJyVOdD/bTLqF+DkRevtGYLULcF9/Y+9V4ksJiN
VRVcqImTOlMf/bb6C6OcONAYjJZanelMFNCp3cUrUIYf3KWASvy4vRiCc/5wSvlR
i7DeoJAbkmgMLdil+kjsj46+sIwVdjqtjqfWNPCuEjQzXHN5kmZpLTPCgOORXorr
n1PbMeTJfjZ94KiZfdFz2cEXcwfWv5vvoeBDDFj4vkHBdHF9qC/0Ifq4zs1jhUJB
tAU2utY1BLwHKepWmMSMSU/cVO2jfoIz3gU584usvrjX3LEf9VZhe3qN+8tvK6se
rELSAauwqwfSZULi7/DkaM8BFqt/tbA/sJqeSuEbslbu6o5os2m2E7c6kRbIohjY
EVZSdmiDjUGUJvS8YeO1dBuIXDh36A46C+T8Ivlqr6YaAkLD9cRZIwGlDAeTkwDG
aNT2Od7RWJgW1dfX3uQvhvBXlrgtC4Jj8YoCbJ4B5BGba2xXCh4JuISKdugik5LH
NJqXTCT0EIzzjagxniyhqVjTYOxj6n4r1tVzn/aoYtL/s7u/pZGzsLO5wkVKQjNU
JCK+FLYojSVMtI2eaJ0HigEoHM5NkZ9pH+jjynPRUwDv4e8sbUtGhlhF4gDUkiWW
8kqtkFkWq5s8uZkHSSj8xNgwWzwW8STqqMx4mjsqkVPw170y51pLggKNSW0j2snu
tgCiqvSgTWJT4YzaZnqkOmiIPAl5dC0KBLCQQyTsfBwzD+jDKXfE+VFWVKrJALIc
2aBWxoEoH8ZWy8thrSDJzVl12p/XRKi+cSIHogcsUYlJcVxGah8Ca1KCA1aGBXOd
LMwCf1O2OETI/7UfzqnHr9/BCENF8t7owkUrh1UiAwhpI8z3XaaifsEYl3Oco3Bt
TTisLZJ3JR2KmX4ZcOB/OdeXoaQ10oP+IdPP53c4esSQeuXaG2d4u1uvUa/8GxuV
qH8SZf/lCawYyPr6zmRdyNBSAa1IuEIifVjX3IFFAH5vVaj6RRvafOmtAtYn6ybO
vhPfKRft2S5TCBVa2yFBTUex2BMYTw76rJSRyjhfWuflGkY/Zjo8Xay/Pv+HudBE
EZxPmo7Nmu2xrABaj+g5Sf2JNWJUw9VBdbKa1/dXP4uvhPnZnB7H2TaPPcYigsA1
2ymCRuiapjRmt6FDPBDEqbhXnBbuZarHCSL18Gteo5JA8ToU8H+vRVOcMRAWSxNb
xFYHsruP/QOIt5x0z4Yfg19tWaqkl3Deb7UxiyVrunrDLd2A/m1g5NeAteCGVlXL
5xbScduBvEdG41Je56RUtmV4Y7/PgZayHirJtVxkR2h8NwmienOu6lVHOuQHceWI
p1PtrrbapWGgpV2m1W1d2Aex287AzekEHvsLGPli3gh70uyUrXPzF6JmeWxunl/b
lgybbqisURJsCBeWLSPA54m0re8S0gijQiOtEv/WWbokscKrYez5ECQjGdkkdfj+
d95lTqmpOZMFYtenEs1PUmdhaVNGmrN2RXFGam6ErDm9XWPR42AsLXCpJ2kShBct
CoCsfu0Fly24ZQ63V+hTMOMgItMW2MXO8wMztUwFj06NjohoyrrOJttTADze5ltN
mJIVSdSWV/BjjcheVzO10PeplTghQlYk4x8ikKNNjI8brko7ZtIWItNjDIXK+3PS
cr8Q5GT5mdHN4AJDnnLcddvU9zv/vDkER/TSMNQQeByTr54wh8EtTG//UJ0UHQh9
tn3L/fyKcO6fwEaTAMcyXq0yiK9zPz0b7tCNpNcfhXQnu1+2SJIdaH16tUJgejGh
t8XZ7HlTLo+nNXfXH4VA9e69G9+/v8jVcLV5iaS4hmBMEPsZ6JMoQbpAt0cfuI0N
iVWbqxQMoFKQVkHnMw0hzPYIQvSVp1S//zcqEumr7f3LeQAoVV1bUW+I3D9iuHsw
/sd4V4oJsuOVSNj8ynkDam4Mv4sqCNUxZ1OKXrZZjOA04E1z3LAnzPOrGhJjno2V
t6Ca4fqlX1r476DQKEIemcXMj4apDOy3mgmAdM1koA8ZP+HUXl1+Te1Wqa60zzM0
NpLOCb+rLkvp5emckbVOvpzAL/DmLWxhN50dPLqsbHYKZjKQLRSlCXnj9fL4fp3/
BXMnfiDDBE3xBnggp63k/vyNWgAGViRXEWN5nuHqvHg/dMA1MjGXEQ7TnLWPyCl8
1kRjXSzMNllKJ/YuqeOHW7U7rkhrcK8UHdx0FO06WtSGPSaZCen0IEFK/xvC5ujT
7kGU2wyXn5iA2mM3fN0mQExWQurBBlDv55VcxIFnoSv3NMGXGZQhumolCHCMrfPW
XNKZyfObdwKqbE94karcpGwe758rlRzjzRFU7f5VWPCNAGNVYC/TYNvJAilyu9gi
iWt8pKNZWW92kQMusi1LYt8uo6GBdDXgLikNUmqK5xANqhFt6L91ArsQPWuzn5gi
8IRLRDtV9IM18Mhwwd/tEHvSx3Kk7mWDqimFOohetXuW4U4Mu0/dXA3/1t/JvmCP
7r4GcL58pcKpBs9mz7PcVZh4ABIzrpEZAR9b2CqemE3HUITs7gnAwIAjd+SYIhz0
ohHQN5bX7FSub4Z7C6lO4lCmdTlmF8kxBkVK2tJCMb1V2Ggc4JGjQyRc3pUL0sg6
22B4/eeblrIwvR+sBM5UH7+LNWDhpeR5W6qKe2nsth6QI2ODXv7xkpQcEY5jPDZ1
Ev9ZOmF8yPXjTvRdNSs/qd36n7pidFe+iHenOrfdBRx0Hgp2r++d2Z+rYSZP4MPk
LvSXNdfFId1l1w1ACTWKbWgUCq318YDIihs+xbUu0TkmgOAG70w+YnaiI79eCrWy
LB2fB/c4+zEjRBVSrWDePnRAGTof5nj8uam7u5EfDN6Zf24dWza+fNhDg4GMXFfD
1DoZ2Hss1wlvcMBGBjJbqdmHVNslvRoLDFjqWoPbJnQFc+gRcL0YNLBdojbJYGRn
sxqSg22KYe/StCeJneo3pwBvpe19i4bKWICQqwKwMlhUo0X2hz+rdiXKbq0VJ4j+
NGzrYX+oFQfPHUcm6szoGqDTvaJf9ed26hxl/r3s4a1jdvvFp2eRDdCm7fxVBiut
2xRS6D/30xPe86A6SyE+YsmaGyUMLtSxwVGeuwznw67vjNrdfaMMeprwdnxYSwNa
cTAQNVpHAgA2OOzhYsJ5E5g6dgzjrH1sug3p0xDqZik2wOdecdk7YKbhCNRn9QjC
645Jt+yrq2QkSVcOj6VoJqBl/rHSiPmXXmiIuFSCObczyedy6RxWvCL9qFcxgfoF
et8mtse/1BW9U5DQg06+O572luN/go6vrkadGO1B3u+3pBGuLYTPkemnMhFgyS1g
1QxBMThx1taXGAuh5djcmM8Emi8DJjF3FsgiF84XHM5MtG2lJKqBXej0SVsH3uTA
1GVDo+Ce5glj5HURnrx8BZH+Zkb1A+YzH7lSfhFtTEs3WKqWNDDeSLhjO6M5RuFW
ffpR7bSxfjxe4pjSz4D8pqntd+UeLupe9z+kWJhHnRENRt+PEhd1DjBjs8gSzgTL
76G6F+6n7GMt0NjkjOkjklWQv7InQTHVyhfnpi1pcyTNqLyL+RGUQyuhLkX/ViRN
z7Afh4fZYxS4GNHXaQSTu4YYltZAAkHnT3gnvGH1CqDKP6TOqbF/BynjtKCKS200
/VSIjuaxZpzlIu/O6tpC6ew6x4YTIReGDaeY7IfJBr3HZ5gf5z9/OdsTKz1UZ9NI
N3kN2dUHctMMiN6YzYa41pSOGDJ5rYl/es1hfZkqHXn21ifxKFEm3t/YsXHxiw/5
dYhfhx+RK/qm6DxQQGAnhOoScLCj3Ke/XLUy7EhpAKDGDziPTKrAPXRlD/s4u9VD
A8mZUExIOMampOkooj+TBV/e3ziYYCZ1iE4cZcdU2n840gLC7ZPZLghFttaHNBaH
yI6Q6Ys57efvlxt2VGxdHm1JRo1H9FW5T7WcZwlq+Xn/JmGIdYhdtB9QOCSU2zSa
/xptiRDNjOJmN+hzV7oFFJNT7SWUcohgeoULsTYWwfnLk+xWEQ47Qt0tMG/m+doV
30+pXgIatX9vaNzdBBOgVROThfpCvHCj+jUMSLutDp5idoYDnBTl2iQM0mtg6vxV
khJ+jpl9UqBJtDhiJZiCCc4XkIqEsm7UvziBkMEMFzryDmp/KR+zzVB6JJcGhKBd
aga1W/scpeFH0VgoiLR95OqlplR5QrZ1np/pwQlWAG7hLmtk5pOZGFz0KjuW4byZ
c7sUwEFohxzRZKQ6RPoO7ZmCjJ8LEIZzqwZRanmZPVAYLAscBvVTDQjhuIJQuEy4
AW0gaeWUuS4tPEAKrUv/Ftts1DcMcTsxM9lmr1onX1IOLawWBTxDGpMOgulhAXKI
nP4Zom9ASPn5dD8r4gZ161HsDqRvuriWdAx43z0pDe0nX62418bhEdzCqDYU9ZWI
LFonzRXHm09gXrnMzG5tGFqBzWF5McXXHzPEkDh3yTR7yJgzJJ6YRw39hza9Q4Ty
we83vUe6lb/OrhDBnBOE1u4jn/SPtJVqJwC/6AXO8uVDqPxZqe2HZZBOZJ5UMimk
/qIgH3lU/9kaijFFV+2uPgbHCRYd3/S+WJ824KBcpaogAPTOLQ9G5XdL3KyxVu+6
O7tAc4Crrv6N8wuv8zqzxmMHEY6rrCVzdc68RB173NkpfnjLmF6XkyBdFs3InUvo
FT33zpUEvi9yevMwJ+otiw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
aqn0cA6KossU7EB7lxZBaqvfDYb/9OOPCe4xbve3s3TyzFkBWVgwAdxLVrgtHqXn
IbeMJA5nFrO1eAjEeUYSgjsOUKBFPSZYOWhN4pIPCVxN5bwX/5bn5Noa1LUWyJOF
lR2ooZqkntBMq0FI0WvvWmHAOM/jlyLOc3MC5qVHi+eiludkNAc1esEVOXhOkVA6
/vIbwHgx/7vQk/66CIj+j7nCtAT3B7xSsuf+xxkWEsged3TqpVQO0MkdzmMP24zH
Fsd+PyaArBTVhy9pSiPxOi8AMjqXvTI8RAM0DKkpjonV9Ny0hIZ8nIsNzyYvgrdT
EdPMj/5dSCJ+lN5iBwt2Ag==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 23728 )
`pragma protect data_block
+3zG/WT46y1sodERSOl6Zv/i+lnnN4ccsXliMJ35A/5zXrhVcy7On/AVySbMo0wp
9Kqxz0oesQvI7Ir4Ft+0MY8s/VmnXTqbYmzUfd5V+fegGE659lDzCZj1LBgFGhMq
daohd2lNzoNHkOgMQU4/gRZIWjmT0nWIzfnfDdCDgWmDi/OVC/0nze15Guegrt38
1xM5UWAsya6nkSdynll7qm2/9dWmycsMPg4sBp1vMEw4xEJHjvyOg6piy92Z3oIf
ZZN4+cILbqo5n4eJwAlCJ/qibr3gGQq899o9HKbfrDkKlyHO49ADeBn5gCBwvHk6
o3qz5ZpkyXZ7c6xr3fuA9qy10IYQ0J8b/JXdDVISBchR+6WGd9o7x23+mJ6evzvW
Y3uCa8WQOdK82hq6riMirSiARxHleu9e9BkNr+fxbq+jZsJbZYAt81N6xoecBnlL
doS8VtLz5QtcHL63HYn45cgGaO5GZF/5Jl41eOFoNmuahT18Eqky6z8nOp4nNO7V
GDigJEcdjFIzDok8ZG5jlu0A7tByZERUNaJJH27pqOfPAUaIGXZKpmQI4WV1p5Xc
SHrS43QMTNVAYqq4rAtk0yu6qqmZHunHDLWBKCE21NYi8nzQ55VE9qDNSotjFPBC
QFFpFpas5Sok5b8+sNVE03sY9x8xlkLL4+4SbOg5Xii0Z7ir66l1E72r47pVTOCE
AWV36m0IWtBsxI92ov5NmBzRcZFb9fCY+NpbVpJEnM6Gze/eZ1Kv0dZ1za2Z2uCW
Yuktk64sRiodHMwoJTXRdk42ijrI4UQfp6ymZLiDLPo+TqXR8t8z5POgLse5BnfG
fX+A2isFhaBIhl0EPDVS3MDpUBx9jY/RbBCGjgbl+AMrVvqz8D12VDmq+XUhwwIG
1h1lvX/u38sWow2jBhEwWKGfBLbgyTCFBNTzCBFWUyw+i+xUwwfM11g07a3aGC74
fc6OJjwZb1qlutKQTypBoysEpOacDvGahBTkBeXTkQJMCw0R7alf3rounVrlhm58
Woy4lazOWK1FPDPFBqWkuoqchiM/jw7xVtQ7ZKwMGMGaRbYkC3F5Xg+NEbtBzzPJ
ccp3eKWP48gF78nMj1/puuPmlj9n8fq/5jkTCSmhX+tVIJ+NTZ9BbuFehV0crMkt
YsAoRt61TnnGKGU1tpVn39ajqykSBokkkM8pUDVs901QN4/vQVZtJcnsosXig7yn
b5ki5pJtOvuuctV6c7R8+K8Cc/dwr5HA0zkKqizcPW6R3bQ2Sk/1tzS7A4Rw/QTN
RMU3hlNJ0JaJynJWG25th3UIVjGfrcdk7wcr0mvsHkO/XrASDqPnpoOKb/uOQqRA
o8gqvZZfihIVY5YooCcr4bIwI2zgNrT+PHqSc8R4Mc6rQq+UGL0bMJ6gapOLMrUu
zjJi8Mycr9mj82lCgbuFdXXD5dI31sGPidsqZmyxQc/gf1EzAw2i7kIMWDGsP+/k
+T4xiUL9ZOeewfhYeqEVMy5ILN1cXuZ1ScCrLvCdhMDeKo4gIQzQybVHct7KwYFY
3kWtqRf4t9Xj/rM03+1AMDSxfUxdGSHh+EqSmVp5ssCmTVzJx18bxfbyPhwaJLiz
5S6D7xVGn8FF8rnttBN2dyFooAsFLSo3n0o5oTkJLpLHeLllS9liLrVtXqKHXjeC
azaLxblwgEgCNrSSQIAZrFvzn7zy+cVwk9ngc96pNxKA4x5fU2WFcvh+vVzQzR4k
0HsCE25se3E6Ua8q54p54xF7vXAxu2XHEc1jyH047gPERcg4LmffaQGvD0q9Vahc
8+7hau1mCp5g/BKysqbQ5JPjsV5qfwC98aLqGHUkXbo5echaCStfYQIz75f0RLYo
QbhczdJ38fwjJFZVPe3U4gNVGDRiQy9mPJKmnC7N4tdcSOEsR2A2QqqH/hAxYao+
oov4L9qzi6dH5DNMwgfSquKgX2tbLBd174cok1Wbcd6Gi2Wn1ebpgxeMPEphO71A
9s/vEMNmFowmtaKe5RVHaeyAvC5uUBbYLCuxSLtDoQwlDJ49JUBXO7UFGiczo0/L
4swAqeBJCFisBY+xVj1pe6XlbHJDfNEVJqlFkeB0nEgxSFtDxiiwS1BvMs7H2x1w
FiSQQC8rNXpcaRGfu6v88vEcKYO6JbEAhiICkaM7sTH++PiGdR3OegZVji/2a0aD
Ss7/lgoMjfSd2Wc5pILUudee3nMPbimpzWknJElltZcVWQSAov48S+kks2YgFSaj
mZdeJ+vGGvLUOVoZgD1dWX8EpPyf1n6o/gVBpUX4d3PCHrdMgklIdGUpNFNFOUmx
yL8rB6zxjshpUIJy+NLLMdUaFPq85LzbAg2UNLAtCp2ETkLwmvppewCzXCbjcBes
yFWtdGySOSeuX1xp9Ak4eULBeC7vulYvnetMUxuajLXFE6HjGFUGeCQvFP97wVqi
Z5BidXLiVU2Uvrc7/eOgp8FEgf2U9HFZWiFrW1qkbE7u5NO9ttCCoMZbdBjcVvYm
yQDHYVKHNqOMIloWBqAYtQZD1NcWRVbxEezzvVsv5PFpE+UP1JC/ApQJOkio9gsW
YvS/yPJmcSm3kVgYXvhTDE7p9j07rxpi3svDsMBadGsRvUSQNSK2/iFaD7oWp3Zm
yOy+ENVGG/+qdNCnW/EIGngElCHu/iyfnYa+D5SoSh8FdqFjBq8i4+Y6fGMYg4Rq
5SBCyE7XWgDj5CCzaqCu6cQjf8M5XCUKb9Dd3y7Ed9yYErwCA+ts+EG/jWY57U8I
QkIi3CiWQTJdNZNkxg+C+4+Py1Djv+KvvnazL/chFZHJ9k2p6XYvQMJoGHz3c2L9
LqYHTv78qv4OhOvIZhwwn9hr15vEjtUOdhZJS/yK7+bbymXmWewvF5rt/lkrFzdS
6YNbACOP4z4oGhVYoSarf9z3H5HVPo+Jh/BdU3KB9cmQ1SV6FGFZi72H1DVXtcNG
caXHVnLqA2M82EIJFnZ1knjFrzBLPBEoqS1QnDUYNqNl8QcpNp/Z1CxRGoGUeAW6
Zpynoft+W8jpHBOMh0pFIZD15T9QmR2iWTKKBBRmoSRMzmqNnLKbRvIZ5kD/AyOG
T9C747VAw+BJGjpXD+8stsaJp5Qz765m1t336H5Y6rqKBif+7kEA3/MoKfq9TKRC
LipF54YqwDEph70ycDVMab9ixKNOnpmuDQSSHU57NXb6ZV+8fUCpLYvV+Xto2g19
453OZsJcjByK2K9j+ANWesjr5dU1H5By5qHfMdP7+WG4Jh6DqJHGNu7J+qLES4jZ
OfUj/vi+EpD6f56pConaR8ADAdIrXw0/q8C00qyXgbt7Wp7gI2lCNX2ksMctJzP9
PPYeKK5CM9reKn+1YHVRBT1ajlAD4YFBG08kuOLBmx22o6CtRR5Fs8s95lfsq8NW
FlJkHROEOgnq4Iyk5w05MCR/rzn2eEKi7gP7aC0Ddg1tju6hkagNKYkdB5hKuUUR
l6SSLbZQBoATiQbfl/uzx52Wdkfv735M5o9T5DOZIpR0eadk+EpxJ37CUS2074xz
oJ6J6+xUW457AoQOmLhFda2Ehkhrcw78KOnsahQU8uyO3/vACJC9uzL040y4ZnD4
fGZ4OeftCaeCGUv44tMqTz5VHcd7QcujTi2sGEjVU+0F3IGR72YIEEP0Xs75MnQ4
3HxKWodb4Uo3xCnOuwCAKZbiYrCWjmsbyUYv8sx3KMc8vJR856aI6BVxozNffw+0
4IY1m+W4yTy4rRn3qH3o7ESVda5J+ajxA5f+Hyevee4HZ4LkNZPGM9D4nIl+woi6
H7I4P7Hnd9xdWFyktcN+For3KiQmvfpkY31J0DTMu1t16OAO6hnO5JyY+afVSMvj
KBQSz94Zf4dsPxaLHLdYBReK4XiMLUsPrQczhV0hgtoPMn/lg/n5qBK/o5KMc47o
GfwZyC5cexZQJsa9qnL/2f+6PqIyDQ0l98YtY+jc0I7weLGQ/AlcduMfEjhs3LW/
yMzsYZvGrsAl3fNzjN/9hzm489euxZgKJtEX626CPdkK9rVuA4gYmnbElClQKG78
Jm9cDg66Xz2mhYveuQ0yvwDgtcihhS2JU8fheANB4EF92VCygntVQtvvelHYZNwS
1SaXj2DVw+E7bkruFqS3Cw8cfsT/kvZHCKbvVTbbH6wWMrciU+IF5DGUgPjeheVW
w0yjGU1aVbY+MgG9KrnJenn9Sm98jPxzig9uXbUNHkc7sodukkir2XSz2xd4SW8H
pJvtMTq9DN4eeB3nwFPjUozQ5IUMaUBGwLKzj8sbv+fAa9MwBj83iqOd8CKgFRES
1XtCOe/XfVdjM+vAu9OLlhFHJDh61GnPqM5hVjHu7ejOCAbjIfNV1jC7cw2lL4VV
JZ8jTXzy/PCiNNE2sOxS4/7yDH7GwLq9PxFQ9TfxBbA8yL4QSHtIvueViopclB6v
lDno//6cM2dvSi9/ZmjE4rb6tzyETBnZjfYB8COnghhugDbljoOybseiE0OPR+RQ
Kg12K7mHXK/xI+Rq847P2Z22zE2LUWLXAS1TFJopNECh0JZFX57Fo6XS8jybv3Zk
H3MqwkaoqKDK+T9qr/2HFAbjwAb//ouPm04tQnrZBM8FW1ekkOejidi7QPDP11ox
+zP+/yxJ6uHnk2bOlpIq2zjGjPnSrwNn8sc4dvhwZUSHwSaDsh9vi/oU/cjC6sqD
gxY/XENb5gwsZ1amYfZNb342YmIE45s+ZTBKMAcE2/nuYhyoE9Y9rmDbhXhLhseI
hH2Vo4F2ebGvyrLVoHpDWcvVawpaVMXutPvSkYUbyStGEFwcR0ePgln8FOmLjopf
rXe06U8DhKyXhwBUxKT2RRyWkF6o2z0HJohjk6l0I2Ybxu4N1phB1cD4kvE2MPNL
i8JCIe9YTmmHrdNmutQPtRCGWXaAk76wivh7zF3qfYim684QPtWblSiiuOdZ77+x
jsQ25Djc2qimjUAXASqcea2jry/BN9ExsJnw2IHuNj847d2sJtkfBAmlGuuGKwH0
z0hSFkhBDFoekgPhj2qhh184AND3afnoSQvd5ChKCLOARxaTnVnE2LAPSsnYvQYt
LGlvLVtzr7YaH6Ub9P5VmHzK9hyOC2TqslgaeN3IKYRiXDOWCWqObbWcMUaJpDNs
iXWlZoU4DNtH3KDMUdq0GWx02POM59C1F/d4/hk/G0MQbZVQWBgLn/IrL4k27E0j
oVA/5Vt7xX+dgaC8XMMjlcfV97VFdmxDvISgJXBGdrrnu3W5o5ubEb75M//fvH0q
vvxWzI+ACCZXzrTyxnE05FYEyT4giBtjCRqaC/9otEHyjL5S1r4SaMz4bhs8VuSc
GapCLzZk6fOyTOG87v71lwkq1Ifx7sT9qFKS0AZ8ZI71S159QyfeoxFvEdGPRZCy
RIfaxEPiIRSDAFNranxppNiA7/IQiMy9UUajsP5hi3O5GITO7XDynaRnbSD0WclE
d6YPezqcxLKIWpij6vilhzi2gU98FaQnqdQm0liS+nL3yFBJ+0wv8jKPzVRu0mWy
3iIavzgiL9BRwU+i9T0M/8Q01OJQ2gEGaM1ue7bSKqHU6p9Qy3i00kxZeTL7Dcwo
6p9a2vZxUqkcl7TN+lAKnxVMYC4CiC4MtPj9uDoSnzcMMLghLNm7Qe10MkCR4LYZ
13RRxzwd/kqvLhztPd2luOW4BmE+77bjTk0MDf1kOyQhkEAQVam6UsA4l0TXAdAW
QalOgDK5FFQovj9F4wuDZMfsMn6qW8urUVl+3h7FNmzz2FwZ/mzd2R0q+xm7HZQ5
I6WpmUVl4fBj9KaWLXWtbRHyoo24S7NS6XFutZbph3BGa0lawG6GMbuQgY9nSRet
XH+Zb7uOO00Zlt7uNoEv7K+XhtUv0/IGU2IlI6mEwoIOQsd4k3596lG+Mts8lKhU
/lQ1bKUJ093/BqP0v+/bam9SAymhqBLSCBz++e5FRwBBoh1FZtJoCqoCOXWqFfUg
FQ4p3P6G3vxszPaNyPKl8YcPw26VB1wYLYUWI3p4+9aKYrazPwhphTtWjaCAUU13
In/8Y3ny/U9iyjH+0ZSXzWqR6tYTI6yMI43rd+T6uQQb6icCwje7y67D9ZgcPAhc
Y00WWoNo1mVNH6Z6ltyZcQltj465V1q15/qCP/jrK7xNAULJuljVBpcemR259H3+
AmW4s3sVgJ90wcHuzmcrM0r3IH7mbmw6E2KD8YDJGddS4BEtaKfQ7xRt63KFZldC
OhozsYzSc7SikHlLO1Oy17BabD39qKjtF3+9/HZtwrl7HceKOe2D/1sAomrkTHRS
DTrVGCrTcEOZwVmqMl99HR2T5SYcTPGfz2dS1Od/HTACOH+auE5bQ6s93miX6qa6
EoBlTCVeb1SKCtDpoxHWJ8MO5E66qydN5gRFoG9KXFaM/V1QLKqcHMBAFdw/w5aa
AsO5LW7Rh55chsy+Bk805YFInwakcEHoIOYNInXsvliGij/OoVUAU7vf7O2smS9F
Ds2LBpdw47ruF4owLmg2/WNBnX7fTuVs/jE32fegJbY87PHmCv/n11oHoKkNlvHa
mMXtXOzj69RnldmAZpSERB8hjxZgyaMs6o+XXnGeIy9EL8VArc5BHDl/BkBfpp5u
i1Kc14SPkKGnSwigJlpSPyKwBKWL1g772tjRmjW4zvd5MGQqxt8td+6/dS8k5y9s
+oFjXn5hVti1l2Pag2NNEY0GxJJqf5Nr8yELC9IqopBNKLGP+8DMIw5vn6rpD8Wf
bvfqM4zKOFuK66Ru+TK1EkLt1mjsYcFpt3ymaBU2Gfgg+60XyPsbxi7IJH2nIS16
ldg8qvxai69EbrfPqVl/Zd1rH1eLWTOetfspscRKWpGKETXdu4EZoHK4v9dYZ9MA
c3tUkjqVOmrVQKL965+uUEv3uMHFwGhUT25GKIeD58rlJs9Joxjj0E/v2gR7Cnda
De0g6cTGD7073eZdRizlgo6IPi51kbxEp7TxMs18K0cRdp8+FmURJjqKaVi2Xh/8
CyPF4LbBLlspDHOEn3xQI6oZ0UUwnD3SgFcXs4uHnL+BFSzgyx1TI6nHAM6w7d/v
oZlnMjuIH8haVGP+Pnzq9r5uNLJOHUvAeNtaY2Y6Gb5yLtNjY5qGWrxNF3L/tFXq
/cuLxUOGpO2S3II08NqSWsnJPZV8MSuSX747Q32QdeSgqT/wOqvMFZJnIrngjTyu
QqDfc9hw11m1HsDJab5CLWAd/k5Sc10GPDu481INABAnwlOTQ41ALn1k02ELJ5/r
w9pV3owIC+suk9wjIP2TqADsrgR2WS5yXufDHYkKpaqNNKbPe2ARbEShYnAqKhzr
Z2MNQeRLbAg+hx6mpFl23ZSxs4abr8Ues40t6x/JxXScg/6cJDGzog2zNWhGuGal
yZDkDc+PkpkiyKsasmSZ//HgimD3BvuZV27Ijaf6xRWDQjWwJYDz5oc0wnZasEl4
rHQ+Oj5fuCmAYOv8H/QCzMn2CSZblxcVjWQ39HaC9x6XEGiq9RoVLHreLzyovwbj
MQIfy6WOGhPc0bvKJYkgngk7jVMdpF5Ro6hoki+pvnabHaQF+Oc/I8UgmPv07U/b
bBgr/1WrVw4PdeonWwyZ3u8xZcrkk6wOl2PcuH4UkiE4o/q9bjU/4IY6YwtQJVXH
Z6yvx9jplA8lh9lu2acj3kyZmGYx7hUt+Jn0jKV/ESBJyS0at3EeoHSHoscx4WtS
OtSXS7aPoPhgUmuSMxfHy1RHPf/5SJ6etSB0h8bBFdZyTy9oXO6j04lNOixh0/bI
3wzUQRHPbTcuC8OQIrIPHgBQ6MtcnBxe2zwc3wsbRDY/s+hB6p1t8Xt/2Kx9Gwan
sYdHztB3Ob4ASLjIImq2Cc3U9qFd9G64Gg3fkN8crs4mkJdJI4CYoBTcKVaG5OLE
8Zj41USNNDFrAJJY5bwwUM6omJChnS8UvKzzjy/vOaf8YTr+Bew1vn07RVVk6Nhe
QIQOYbm5VyB4sU+etj86MgXZiOj/rFbbTfps0CsI2NOScCBcJox0m65zTsX0ew6o
zhuC1f+ro/A+k3FPNQK+PUUi7NhNzsvoYD5e8ssg0+YUkge7oWxELCeE/yqiYYxx
09aAQqT9IAHLHsbu3LZYStrDMbzcCqEBxSohfweTQw8E22XOG8QeBYAzkulMP5lc
41+ey3sU1uz/EFS8tloQASfzi/Rcfn39+vGSLTF4Q/swTLAsabAkqoALRbKvnR9H
RWNq9+iWk02olgjnTtZitGUMUr+cbRz16UNNrbZx8yWlIvmgzUJ+2YYUzWeRr966
XkirRLh39vt25ROxPncIoN9xa9Hpz8j8aEnZ2ZP5iDt52FGDjYlc5Nau+dHT/wn7
EXXzJIcO4KXwibaMBVXiL08DeeLVVbh20LM+i/A9Y9vGEvexwnvZfxEmxVTGgxcP
Ri1sA6orF6OPsyAq+CDPb2OnThk8vT1D17hnZ61qN+DmyzG7N9fJqOoHTIgQ8wE8
Xej2tKdy23Ard38nQgEmLpTcBQeoKwQSrRSpOpVPqkyr1MD2Z7eMh6SgDlefpI7m
UqK+p+wIvc0nTm64svLeWYgiww0B1ZdjrCJ+oLLaRItbJW8jCbTem+oMyWdnk49b
L0HBz5134zHHkQLFoXhhoE+ZmYncNt/W5jUDx2d2cEBMVlP43orCc6clG/pehPF7
oSPoHMbxxYn7KWWEMKIXzyZRAdEjm6MTTcoapcTLDeUqE3h58l4X4fWdrr96poO8
9jEGNaduxTJbIkV80IRlrfOAri/dpfGLOTDdHZ0XJlzuQtGtv6i3sBXLmbt5taGF
1FdOMkGH45sEsIldZQOf5/2f0y7qrznKmm5opw9ERQX10c9bcdz8WdzArQ+MuDpC
+wxW/lYDq1XRfxTuF5dELALdc1QkcsKDCFTSpiDhYAhr66rVDuPfHsiSfXvaO+El
sEkAt++WQ1t3tS4WMlGLCl+5jbL4bJbXMx5kA00M8s0SJS2X2UKSshCt0TAXIILf
AF0bG4LI674CPV3Zwl0PjVTXIVH6mgxvCHLwMNRSQh7qewDoMBaQogr7OBOnJfcy
30S1b7t5etQMRwIIyaziaXwpadCF+m+SiQDbDSH7cRYBPeeV6ZgeUpgS7hxzIpD5
RqINnsPgqOgk1osVvyQeTUNr8K5AFyoJ76OLfXXDGqDx6D84f9YiKjYCKLYVUY5i
oXIuhLyyyWNVFxdDrPozMgwtMEEbrXX9obVnhTrvrAXLXvl33JoL281uP0ZjGhi1
kq6hlTSPht1Tf7V8DJaFuV+1BMIeYpT3ELvmSCtGpSF7cmT17XtJ8ddp0R8x0bkW
/YMpUpE0wQTD673nuAr0uQyWfV4Ylrxv0H7vCgKvlnJOQo+iUcceUYZNPNgz95EA
Eta6IC2lweWUvBNphE7jfXAPQCZ/4pyOLcdTe81VKzi5JimX3bHg/7/TQpyavZ6m
wggaSibRvBUfrkbjm7Gr1740HCy8qiYNFHNvZUvQIKT6Gk0iv0bBTEyFdlha7xoP
XHnCGgfCgq5DdOmZhur05IDZxUp5po0dXrbpFm1jNijMefrg3PioVBgz18WnU/HJ
9WEkZZEo7jrnae2LnGRgd/NzhekHGWyCUZwj03bvRuT15MuEU+0QEURutEBUdXTf
UMJt5hPNXRGFCPlr22JAFuzxAgiwK4Dg60LlodMYx4hvkMs9fTVgduTquhDYH+Vu
MXga1hG0a0OzCtC33NZc4jFC9Lh735mnKDcjIZjcvC2uGI2oMXS+Jtx12L01m2FT
tZ1pBB7fcod/TQgz8wf95xiAzBAfVWHGz7ruckm2Q/W9ASeZceJ14vFufKk6mDFP
GEXx0Usip0U/0cRxte3Czr79SV25eDwMRRQJknB9jKQYSE2ogQOI1Gei81fx74nZ
vTwHB6NmFsLj/rmPekN+GBScKSiMxg5Y2lUZCd07iCU8vn/nyYTRY78bh8fERh7m
FkSL8MQoKpce556b/zJIfFZces5tzz9SfOWsKmIZ+7jWga44sg6efWuBeY8O5w/u
aoT95YpimciNArogYXqxk56PKY8r75T8clk3ITgEs4uwbv21XGB7ea5aTuuaajPO
J26AmFfOk9bOZ7fAkX936mP+R2GL1OXJi6QH0Hb+Us8UejagAwdMdpasyGbulslv
dBXEhtcR0OUGZMs/0lI5GIqdiQLWzOjlQZvcbHGfkIe2OYFHdLCeVLIqYQIjn09d
MIfYSRmRGKevq1MnHx130jvBR0OgHdmDGubzsYDNnhU2PyGgzujAeKMC60aedjdY
M9tAJo+4qgdKFwZuwmlou9us32a+dzZMdRp4xniiT5rpJ4ixHxlngQglxEBKsg5c
//NFhgNZTKUbBGuOZs5a4rCfe+7j+AmGvBZIK+D/MwOAEUtnCxVBCrya6i9jXelv
YRzSIm3uSSVVp1+Ej7gRmu0GxGwzMjoN8nb29SBYsb5e1x0Wq2Q4R9TuWJCNJbb7
RXg69nzcdUYYsQSRSvcKft7yxSwI6t4RBLBQkup07GsKoL6uQxRrXgD56Ajq+2nx
XK7RTfTAmtXmVaHrecNHt+Bh4UhTpxi6yxbWHokUKC3oL74cpbLs4U8Ssf9/kYHu
ohCQzEIfJugt/jn1/zfFCBRxAAY7Kgz/Z9vl4S05iP6NuGidMd7/CcCiE7oCGyGh
Cz7s4e295kdRvoMNNHP0/xhYyd0HqvWSltRPYE2of8mJxksdOO8UFGS1mWTB/hc4
19uidvWYbzkItonh6hmhFRBCJdmF5QGJPjYQ9cJ6dGGx+ee7+57zGaWTzlGg+gaO
jhJf2yI0JxTj5FX+wOW65o5D2ipshm1WM2+FwnaB+PF1akkpAg7SZtcZ17Kt9NFX
+5hMzgdsnUFyXsBtRlqy9mbZxdWQlMOOyCsU+UrweLFA7eWj1l34cOsLiXCx0zdd
+Nv24TxotjQVP/gcXt/Z9YOaN2GJnRmbOJTeNln4RrTkDMb4lF6s6yKSrspw9cMF
kNCI80l7UnN7+CobOak8ZE8VksUMHcgdU/2h9Kp7M23Xf5KOOWZHezhlXklMo581
cOcu9D2ooxY1yP0gvXi6yXkStpMXI9LFXzxWmpyquHs6guh24y9+R7SjwR/97fMH
HMd7H8RXL/MLhVCTlZ7VD0rJ01P6l8xX05rk9iuekybaWb2zIwCG85ZSdA9IwvSQ
iMcG8yZz4ZDQsevbdkMypvc1tIKb7uP1cD3yqXpu9ZFYyzbZLoVoTwo9PKBBWGub
/1zg6hotfFELgdYD7sbHEIeDu2u7U6bnI6yZEY/Lpmp8fI6YsOZsnrTk9afrc/mk
OtmIQWWhmJfAkUZS876kP1aCYLBTJtjLof35CcaNXqKyBubW3WoAlN6+IsN8CKmq
REEOfxNjjPhhc3WRo6WwEVMtysMtwhCRnysxB29obu9yrvXcWnxstjJfsTiTX6RS
PPlyzFP3C/oIZ9Y1dnhSDEqTAaK5dZSkztz3kI2Be2/X6ICWfX1ljWC8oR7j0PFe
DVXcpUDbl5+Mev0BTWmL/ZWyW2+gTuBA9pKm39qIezWZjWHwdqLeCUfdn8w8+wZJ
vpEpm7eDu5ghYJP3mKVELC9AEUSvBM9BMi86BaJYYXt96NreaCTOoIoXzzH9HzBP
6kHJG0aVRuoJ+ldQEyGLEkKp7ZKe2uWdADWW6SdEJPqiq9CgJCNb9g5sl9Yf3YCs
4NhYTVXO0Bqb4Kn0QEA4wp89qXU09G3Hzp3p5VYV+gGC8BZAGvSSwd1lxYelkGHN
XPN7hRYeoh9B0Klh0CKJCKKTrE2xxeHMOPF9UMGN4V2zZTDldDvWFWjXatuaJD8r
rxO1nZphoBkyS39vHuSYWqR9jinQTfyhZSu9ibuOqIB2RzDhOTB85OENKNO0wxpT
xje+JvsOoQKGDqBROQBqTHiEI//i1Q3XBkfy7VKQSw7koVb3WJSqhMlQOo8Jcc9H
ksizKW0B0HqPgpx6DPI+OMIhRSOkNA40bcp7rp7trN4T+oVWnX696ywK2ppzCMaJ
NA3LjdEPIEynWNvNBdHeECm8KL+HqZp1l7mVnmal/GepE9mhdQqYh9eKwNBWGKDg
e64CDXvsl21HjdV4nDTodoR2xFDBQfZO1cTdmCiAiIpMvVMBPKMmbhJHN3/XLyb3
mKKoucvAUsd/9rcyMOCcKXOowo4Z91QQ41pyt5HbOTjyeVzonrqe9FFJklp2aOyc
C6CDUkv6YDMkTJO3In/ZhFLYH9nulx2EmuIVokM20TLECsh6Xt5ijoQNzluhhT2t
5+8168wrIsJ9ymoe82vQ4GZfYbLhhf8ns58b05X0M3NzZ6j5DUgvdfCSz5OQ3Zs5
/grLzvTl3q0ynCNkdWfCtTSgQPKoIuVE9j9LHbtM+Liq620Jd0BlTMrK9DNMrI2M
qPv48eQaQdFnDB9QfU1vjhHpP1/hOcMOIxpiVNQRJYp/b+r7M7pyREUqtvJTapnm
kAq7Wn9aiFQTriKJsfWpmqvvTZiN4NXeS0D9Iltzai15zhduFia8p7dQkgMmf6OT
xVwKHJqIAKRy+rBvc7jNN0K2nGqzMThMOz1b0u3RoRRqTg71Yku6exxGj+x5cgIs
0UebSbIj591T0366hUuQGaMcE+3mxd0KeeIe4Lm4MJRZN1DIl2iLE3iX2K3u3vUm
h0AdaHp+WIOiMhmJBCoMY3GO2MZdMZdbxrl7usMxfU45tCjEAW/toz9bSU1t7WgH
IbiydNbqNt5lG7fUhcPdOV77stL+fcUV4YcAYxY+WzGB1vup7xcrMM7wdVV4v/Dq
fqYhwKxGD94nFog1d55NHNOaoSkHTOV6JOyt0E2X4LAwdTpgYAr+k3OMXpmMxidU
o77kLeitUPDv4qRkl/ViLOOHI7JsT5MeX5K4HOAw6+L18pZgP2kRGOa8ptjACw0u
69YYsFrqghBQOD7y7OGNn1u7oUI85lJ00/7BYfm1eUUiAA3QThxAL2Sj7/nj1LQw
9Gf5sqwkPud7K77bpnLAa4TrK5uOdRcX4cefQyUGBjQHcflTjEie/XBmXzoamIla
Fn4PSpaDGKzkjMwmI0jCgUVOGUqndEdZ26qyRPfFJIuoFkU9822hKRzTmEiu/ZL8
nW52Rjsqln83fR0FESM4+6Se41QQzu1+UAgUGnih6UNfoaOntHqw27oCbgF0hXtw
gx5l3Cxe0uQb4tCn/a0stWNHI0JM5tbkdLCF6KFscIv5vyzn09O42yJKkI22jQ+Y
wtZvVYGltaSnth0Tj2W0IR1M4/NhSiyuMVnEpUW1gTNeL1M5SHrz4X6c1QtQ8tpv
cBxoX3DlvE+eLx55/mOgOjPJrBzomPGdOcDyTfpQvWoZWAg/0YDcWFj2WilbYCiR
lQbG/6SvsUhvITTaXXoijkr3dx66k4nYVMcsM4xjodAR26Y1PjrVxpMz2kCsMQt1
zedPIBdz9I1mLxLRJ0/8EPBl3AEtywQH0ausaECmrdQSA1phoOnaFU1qeAN2gjY+
BkGPs60rFdwOYCyvN0LF0RniWE6nK9X6vX3OgrQyav2ORDq6VqTS7fUuWKxyPiGK
0iVskmsyvffRIkWgEhQaptGvJRJ7pnSuBw0sxXOUO5NHYVdzHXk9XLtHDg7KRCnd
Pl/kb5tgjunco2RRIGIdnjlnRe+RwGHml4MQFppHwxkYW2t+e1wG4OuaAgABrKmO
4XMbA85hXEuBmBznXVgWRLEOognx7b+kYBMI0REuTroeLuAJero2ZmOu26D9VVo8
mHTsdgC5OfeUcPIJOZ3jZtzxNs4Y+mqs/qTDdB7I4yuDpQJj6isflvAp4tmF8jGY
nVUMlKmEVV/UGcR096zDkZDB8cFmH9MAol2CoIHKCr1cwVMyW7aSAFEFW2Vmamib
oA3xhHNwVPaQ+oU9Yk+8F+5D/5N/M9cqtdgDClFCMkl50VwgLZr3MgKTMDpewy/x
v1ca4GLk7m+cR1+/qao00Dxj8IFhGLneF+TezyJAloVVTZVkNmJRYyRTKRUx44xG
3ipEkS9wRMYM4iteXhlalnPbn6VyLTLcE57XccoiTFIycwdse65gn2VF7OSeSS69
rBeZyw5+9wiwre4TrKz/8b9VpNEVp2jSYtw4WE4Vi7ahlGFVr8KvUy7863J5Dd/h
lBV3q7NNfLFzC9cOA50p27cIMUMPLst+hOI/XHGxntYy8cHL5VA3IOlN82lDALkP
BTO95TXLUOPsFfNZSp3NTtPedT1XpIJsv9IClDGrHC3TltT8k4tQ3qz3DykF1qyB
MUOZGuZAgEagP6oAOBu0gnHo3pVKQvJ47UbBD94Jnd2QVG/DLx+rr3JnPEmtbyyB
sDsA0IpUbBXBK044JwYhfatq1vSYBaZ8klYrOsNOR/37DdfaBFZS0sem8QfiriYO
vHVLIWhOInpJYD0tpPlhjqNnFe1vfUujFXg7k8fHMKjiFpv3zS/VR3xK1Wf5Rna0
bULD0Op6hQUIvPKKrrAJ/yyrIT/x/5Ot/GHaiEYR049ygPcMgd0xqlJgXD/e3d2C
A9UYQaufuZbeAVmLAg9rgV8unJ/WPyGdsGhk4eMZRH1UkM5jnKNFnt1QZD3tRJMk
NrYTfeKy10QGpMdkIHlTF13SDVNJpNKFekaCof601anFvAkP1Ws6PRPa8lIRVljs
lBSgrBz0CpG7Kezv0VG+mrn5apDzHGr0Z+TDbFKT1JUmDW8EGJY9YgaWEsCDUnXg
V1oRrORJE2JYLMR8/qnrYfSB+JljpOxvWLefDk4XwV6yeDTTSFSH7C0cgNCam+vW
rMOcJ8XV0/EJrdHowTQjUGeCkPAxkymMWpVwVaqxC/BJTTCvmw8v+HyUkB+IEdDe
Rafe/L9HssCOsvX3fAvsSnuzs6nt+4cmrT5rVd2yJWjmdC01nk7zZYaekUQHfP5K
i+m5GcTEDl73CWwt6PBTPUcORfmM3BreDPOlgXR0w+5o4tqIXMIgVjGV7RCgSceo
TnYdgPUvbsATfL8Cz0COXzF66NQ3g93wKXNqu0tOvmc9wo6TeZTWqLDt6OFw5Yna
5yIsWU5wXqIiVW0cMhEMcwpO7mw5J/5l9RvLiMbZavWw1OkZo0wzr6K943T3bkNs
hSQ+Zb4VYkgCiKGxyDibWq1hhZk28fHYxQw1hnbWH0ewNBlw6KKxCZuT6oz9dFvh
MJ4FhTVZ2OSHoQ1LZNGdGSpUCMnLUAidXsLsLoMUPKJqKEQokMZrwIv7EpMXQVFV
nvyeXe7KvmX5TZj3s/HWt/LCTbqmKX+IcYDVwrKOYAIPWK2iHK+cyGJNCblglXXu
FJQ7A68suOQ4kDVFgw3fjbbotXl9ZZgvQbA5XcXdQ3H1IUg6WufLAgnOc3/iwZoz
KvjhIlj8CZr8ej+/0thvBXchdDu/2E9nwHMWv/CEszKrT+dqkFD3HRYWD35qcurV
VsC1/guzc87zW4O1GTvvVmidPlsaytuGllZNu8FAcKTMCoxO1kb7pqHaAkG9VjF7
YFOEBPwVQeYoKsJyFydHLNR4WSgXP6nJIf4yFlUs+/GKlsbwF/fvLn4G3CVmTLkZ
B8kNMGHkcN6f/4rZ5Zx3Cio4gqCh/cp+hWNrWDr6N6uRUiAxteMERv9SleF/Klqj
Un1k/KW4lxM0/TdeMWQyYjJYD3zHGDb7FtbqkDRZjoKwHqrvmDv2B+FiNhfhquvn
5dXn8uqeFIrarfll64k4b2AaNqR7Q6ONVXsfoTjne1tPJMZaW5bspBwbt/1xlgqL
ce7QGSSyxmLQmCdeCsh5OfFFnpQgcistOi5aQifjuLQTwJ3LVfx0b5HHWTKMFmqp
ChSSVbttmL6Lxgvs8ZFcXgm/5Ib0+lhmKXKPy8Nl6+d8TpUYpevQICV4iMjYdbl7
D/Frz+GI/0yd0Jn9mhaePh3hb2GZD7LWZaRCmNbJM5Xcwos74HsnVu4jutofGuw9
FC78UiqFk7l9lwY3Q9tuhkNdRFZPWaZ/xPbN5jCvmUZ7zU/qSlYYzsB7TggV044q
asg8gqpYEJ7WMbpYEkumh/pMB+wj8Ok58G//YL9sescmDOton2LPuBNI1Q2KQiPe
fop27ubMO9mt7Ey9J0OuRvMMhwPvKUVceOJHE7MTujQ4BdgUHWp0tXjkpWgW6rxw
N8cGmcuzvsKAgrtv+JIBDvLZF14dzxSmnKe0uayCgizrzJbg2oRYy78AVlsH/8xB
fJW1TB04QXS9F6Yeg3elh8RMgmMQollx2LFXjAlS8QqhQ1pPr+la6jK2ivbywAin
8frAFKVUBZxyQEIhe6OEJ4RUckXCsZEHzQEPfsyxotyqnflBNIhVTmNXrh56Wo2B
IEK9EL3QPMWJ51LK7QMvCaqNymy3UHtRE01EqQig2vDr1sLoNebZSqiTXOFtyTFh
AjxDkMbY+ZneMROtjYXs5VQXhQFLr0k1/IKeV3xaUkfxI88TTJz7Aea9f8HmHNxV
CIImrT0GYjM6hzAHeSe1vqJI8rWV/XF58K/ZUdZ7rrAF3MzNB4CPj7YUC0NQ3Hcq
ESp3GP46PHTqhAbdr8/GObF2sR3Q7Njz9z6HU6c2mAI+sa/HEJlOPpJijLN7lRWk
joA6SJKTzQr4/zd1gFjfcR0IQvKaLeIqUukL2z/TMDWZOGovsJKbqAYnszpaijbl
0tUCGgXCtGoZcl+XGxTlZVzQx4po3PxuVTCaanlSXB70C7ocTh+pMSwmYiVv6EYD
Bl1q4I00zqKl0iA0+jVTD+KnaRk5WLFqpb/3m9dujra6LprVKUXM+I1Fm1bfo1AB
AHJiUlWyBnKFHoAMavET5js11sRzKO7iXhQjjfMIuaOmqpjOq195aamWvGoiZbn0
reRdXuJNdhDwwp4MF3X/b+mYkRXRuoJX5WZkW0v5ixk8lI1JvjWeZbURJ2UzUKVL
rOLUaq7W9Z2nYRmXDT1p4JE6cw7Nzb1FU1X+QIJtaV0bP8CURPAJGc9oLLl9TLtf
e3M3QiLJFnBSIH6jlWSWId8/iSRT9rN0iMxoebw+52/8QRBusjJpc+r0p75WdqmO
qYa+D0/MXFh1jAQTOX2s0UBtNKDbwUms8rDvEexSmaXPJD8WvS3RH1EuiAZMBPyU
953RbJvYRQV9JwTlX7TM5i1BYBugx3Op3v6OJxcmjCubWpYGBBFx7zK1+qr5rFDp
RdkkLa0h2FC2MvHk6kbvKuBH920yPXzII/wpJ0oVCepfox2tjIJVihzGV/5EErMf
qhKDlwAx/CyAmUZwMJ8qVopAjTKUD0XFYOV8RL0TGFguZ1CC7IgM3QpdcWyCT+Vj
8ZNkm6OL9SkD7AMAbsZ55D0NBrXY7Ygk8xNM6tk67+h/1jFCciKAOxZrCTtYetL/
e7aBKeCSTNqgLfqUS1f/FFliBNqUbGVZWW6oVy67v86LcAOjakQrk45puR+/sbIC
8X0m7ZrOVmDh3wrV1vKnKR7A97a+cq3a5OH1+K9G0aTA+3Exv/riw+4ZliisDJ3+
3tpeudseWO5TblBlmGBKfQrW6TK7PgEv06jhNqyLdrrU20iGyuAgNl84TtCB5F1v
95ZXQwId/qSn+Fabdohu7jE8DQSLfJM4zYRaO7ffJ+YGbC8bH8H2m3GDN5FAHfbq
AYa/3wDpqOT+1H3Ttd9at8kE3uPeXGk3rcin7Y3/zOSuWSse4i8IqocUKpdqvYgC
TvSzdWSJbAFFCpfvR5vHqKEtux+H1nIWDZqu3hEnlzUAyhJbBiLGMMDvPs4oz+tf
jJzzPWoxLVyyhe0qjy3Qzwx7jY38AnTnVt3lwFDyMfOEMfbm+3VPn0Eb8n59IaVO
bVRGF9nXhnyQPMONhp0sZLFf1aHWbGypMgN8oRLknfVzmt56vGCtssOvgql65D+e
BD6QqIuhtHjQHjmgq0Uz/UHySMBvOiY6Thbfd62EW0s2+3mQlxoHCA4FTfiflAUk
g2xad1Bstm3kw3/wFRhIkcG5V9piDSkF5nfj6e6UvPeC9ld6rnk7mFIYsWzyvr8k
WeJcJnhIbUmS9IyAuI8HV2jn1Y/aophVdVpQi4kTDIAnaqx7n0W3aoa89zF8B0Cp
g6Ws92euhZ4KQ5300jFvDyUQ2lz/LsgFORy6B+JC6sS+UvXIgXoNcJiGGgQbYpGa
cMu3ZqyokCwQNDHQnVXH7GNNWRj9fbAAkb5t/ejJ7vBlt3XDtTVO1iLwv5fR3ndL
WzPgPMVyoFd/VlpxcMdoIhR+mITtOBKhtbjf2WqHuOCRV/J9CMjK2bjRvmBxv9ji
SXTOIezpNm5d+AHcxeVVt1RX/OxqRfQa1ebgbArnhWB9TGb7hnZa848i8D4ht+fE
rxsOjW1QVxuBGK4RhQrOSdGHcEarbZctnErPK7ZyOcD1ggEF/C91gznGpqq71JJF
BXYXDr0lEgbsjxiYtlmdPN1RjR2IAJgiJYNuvDbN0pti18kiLOOqK34WLwSb1Ver
Ql3JMPTBvN3YdLilCrIsqrpnvUOaQlrfxNf2LBwnIGmp+0yKNfdt1wA8tEO62gOQ
um9U9TO+nFydqLPWXElI5iGV5TYLKSF1x6GErs86uw138zxQVyZmDMU7t4ghjj9C
X1kP05ff/AON31XLMIOKdcOs56XWgVpTldxSqf90Lx6G7nminoJMMSkKLWd2pD1E
IK+0uKg+D48z0GpalRYsHSVlZEzJz2PwT9KbLv8tjOxlf0n+mmUtNyy7TqQvsfGG
5lqmjkziyqQWjKk2Qy/EJw3bkmJYuDaRnxgTAv5SWMENWaDmxcJi1mW6GFtNfLnu
0HGq7i4W4agKKkO3FXYSKbrRBQCFSeW5Cr/HaWhLMVVAGPTSkzmfbAEZIABY+A5t
8W6ZngNRu8//4yDPhWa9GE4hJEBRhlg1WOkoRn8yJUOwzsrHnNQVspUuErXO97F1
uko97RPtAVDTKs/TBwktLwvKW6YOthOtmK2hdDFsJfslGVSjRKRVob1BLg9nv2W0
FEb0d/9lklzHyJsq44luq6enO2HzoZmKb4ZdYIK5/4YK2rTpPWFcrlH98KaKBfCc
BpR3GwZk2tsytU80AHy4WSek40ozQ/8+VXiWyiitRkAwiI/j9R1IFoyaLilvlAJU
DSJ/r7KFmAIZGhM1AiCLm4ZjbdgyN3MpTDD7kLk7/1lYEGp6PNXK1+th+Oq1nc6A
fCfkc93+Kcmw19XeA5iq8iSgjfC+wWXkR34CaXpxejIYq5Kl3kxJQbsP4nz/mzKh
dbI2sh3mlQSEiT/+wlr/AJ34v5uZs5Rgj3zS1u+GOijeP10cM+ZpOSf8FBvEFsMS
eTFy3KZNRD1mhwyNgBt6xX9W8vY/lMbqARFCtlGA1IxXhHMfkQQ2cuBNOk5rLO89
u2snxAUKCnfTJBRgRtgeTKe3ei5ASK/b9xkiu7W5jyoE8BC3SEfgYSmKzrfz5ieE
yXIVUEaSYAxwBTe5k9OaIjhoCRrm7hZdLoX3HAJAWhrs5kLjzaIR4aja30XtCuEB
LXFvX3I6yaIRDQ7JNApSvcc2mTIMyQEBMadY6jr/fsJRiFDEvw14EY3euzSC6TeE
6a9OM6ZdcQAT8y1Hy492miAUL2A7ZMnJEJS5o+gYmAFZkhplfWZ63TefYLiiubf3
yRa4aFWTi+eJ1KqvuYfLBHPEjforE+VJzMoUDvfuF6P8pS8xaPqzUnFL8YhICYJo
lc2t6T7OUYpbvvAk7l5BPUupm6FNEbKqJWRePjGU/tvRT2opnTwigTPRJUwDN16y
ba3PxWIgAngZK/QkfIoI25aCIoPVu6GV62xVOkGPtnyOrbrPsZ2Hlv/XRowhQ1gH
t7rddH9dMAYor/aNHM/qqfyKKk+Hb53Q2rr7pwNHw6wNtpoi8YpSmLxVJyCM23i0
KZ+Zp/iNQZF/8X2UNhLM4JJPw+Ov3u3o4VFqW8dYrFIaMUqucAESxF64I3bWsYr0
JZ3NTXCh3q6EE1CKv58Bykp4MGywnd7jlYNkNIQSxeENkb91/ruRC83YUIpBxUj+
zQg7c16N8efcjrHMry9PvuuP3wjAha8kysnvg5wX3bmmVcgQP5kkzIwVutFbNlX9
E1k8Fm0a7ECYYD4bxzb81wmUllYlWHVICicV0iXsT/VNw4UgDRTfa2F/JWPxSGOX
F5FS9PZMGwNUdhIpI/AJClRHruz2ze5Z14JKiPjl0i2BbKkCX7pB3OG79paVkEAx
9ldQg0Yt3hRCA4tbqXQg92pqZ6GFYhhaxjp/FULWp9xbCH74wZBR3LMsU95mNLJr
CXtLF+RwRuEdgoc5OGvGQszAmaKSDNq6tnKbTOxOUk6TMUMx/CAjBC79XV3X9A8F
8JEkVXU4w3fiu6WP2dWq5h69GxUU4tTt8Saj3pUBhSF71xd6JO2YZJ4NxfRcCAQK
NqdEGamZ/0XAToRQb2EYNbVRT2YYsEfbswTWHIePrbaxcstkZtMR0pTT64DrSEkW
xx7xCNxJp3uLEI9S0N9U/S9ef/mEZQ4EQwHu4UwZWMC2NFO2/sXTA0j2yXIqpVeT
RneFqEB7Nh//APgdm+3BBniRwWJibJWB/TskbgDHXZSSFpal6+l5JYlfp+wEVmZm
RrKCjXPiPTLYoVeRK97/4upsnk5KzLiBDAWXjDqcTrbhmbPC302m3wD9lBq+zcwQ
BTuEmK+UXMgrdPBiWHFUQ4FCz05PeMKUQK0/vOhcnrA9ksCYHcDJArgIDAf9xZp3
VFArV9lbqyP0HtKw45NIZZp2xuItZK7CcJ7VTbISTbSSw8uUpwHLKfVYZdLpAsyj
E9mbdsE4tKFxduAunW01XOSYhjpDppDoGNWOoY3Hsq/tqsAuqjqlBAyWJ0x39Svn
+Ho0n3PCNZVdiKoIDQKHMCQVoq4aP2xmejkRgQu55AjEj0Bem8z8lIjireI5xykc
HPzidHkii+cEVgRcL/O/4x/hlyBzBUIvPEQEL7TJd6LiiVBv/j+1WyVpAiCfr/86
o1dgYWQjneUzZC04+RBX7wJz4azu85MsOtFN5kLeYSlV9a2YRr1BLvzrh3c/9poX
e+umUe2210Wk1LgwIcY6suRPGhV59dmrGukY+Wu7m3s713qVZGB4r6PYjhnwOm7W
TFRU6mYs6oVNQSlEd+RpXnyF/juWxoGa+oEPFM3uw0+f241arIDCruXVOwItt+p5
EUcQjLA4pZp505g/5WClWqnzTpomzuz4fWv6Wziegr1FnZ1brKVmz7j6Dll7Zf3p
RcIrPSOK0TN8zEAjkzVqIZiUMXIE12W+fIuyPwdLqKb9BEivkep2wgPw0ARjhvJE
W58tpQFEIgHqm/tyqdZAT2hA6w3pviQ1epzrv/2WZjeth8bbkWxM4iIssQ7VJCMz
KNaNSYoqeyPIBqTdA1F3LH/p1A19AUs2ve6KWndfWR68j2MRgYFOXZYWdjNdNIKC
Y4bu9lCvkcsC9NIglF+6NPxCJ4EPf3CXbVAqjfjUB3h7NLDOZd3GcDWUllp1D334
5eNdpcWOy4JzS8YSdPHnW99FJu3ShbQjmolGHUdZcm5GFdzAUmaWST0VjN/mrJAD
MXlonFYn08sWuDbnBQa33ebkGYH6UzGQfqNsss0b3EkjBioXFTX8Y5JRn4On6NE5
rng4d6DiVOgohCMR6i4J9U8NpD/h1I8O6wBnATijaLeakwtsVTYS9e455VgQnQq9
ExIeJwDF0o4xk4fAJXnuuuGAj8sTW/ZfErHqmoPETe/Pyomq9YxkWyle9tD4OdpL
i9R3DxazM+DiE3AaR+qUs0qsrywbIx5V5874Qhd5nw9LDASfqx2DsXkiXOMkINey
MoQyp2FFDzo+0TVTSDr7xZ+yzyupMNbCRzSHy0o+yUgQl81j61NvxevREgYQvXjK
A59hDKL03Xc3LwVsmiBRfbluz9cIUaK5JF6Xj3vuB0KF3uwcSkX3ywH38TSkx6+9
JLXEX7ZVPEPDyr0f/T5tVSeh9JV15s59K2LeGDVLrywSP2wb7z681ImGZd6JTkXO
jnhWB6hKZvsdUGTN4t1Vrj0R0AnQ0l+B3S2ianIN/XM3GHZlDQRN/Wb26wSaZd9a
ca4bF2CYQGJBnCsV3tzsYBxUP4nKRnjNJLb2rYjLYUGvuF4+4eeHjtG9dxnvyDI6
v3u/SoebBo9ut/qly027tftkiAyx+6F2lLP4aiT/Pj9It4NcyJB+X49Pp3xmIaQ2
4lXubPgbwOWhLoXrQ+El1Us7+AdeTCmHliIIof9TtZA5XWMgpYPFAK+LrCLLEOrD
qOZDgOtAivCC62VTj1KuZAkRF7bH4gzFuXbnVv58R++6Y85vFEEm3V6AlTOpIB51
wUZJLGZiYCoqWzihPqhTwPEHKsrMhQYY/qTM+3ogVL6aKf0aFtHFHUbP2gyM6RW2
XP7KYJ1aqdxAoJJqaMYlKaMimbCZ1yEic5MEDXSQSAp7q+wkR12m7x6V5+vT6cI9
PmBs4E8BDJpcXW0mt5v7UHWRRFfPcwJWztvfQ9H9tPAvGW522FUY4+87nEpEu8Cf
0A1v+XY12dwPutUvtyMqV0rfiov/tAEy48WUFvHOIxkxf/drB2NscxERfWWtHoUN
3DUdNTqZG9VroUA9xCLdtGoeutXbNCx5Y3hJWEn2Ft/c/BttT3EclqOt5WsBruQq
ei/oFDtilAJOajVE+r9iOm98Anoz025Z2gOo4frc6UEbYDFzAnpSmBWDa4CTJ7En
buV9ymlY6LgN6sGVzL1PRBXsMbLH8+pn/G/9NGa77uFaznZC3pB1sUlk+3lhtYh/
7w/OveZCAXgnuqs581OZZ7B/vk7OPUdZrPAx48wjpnVqE9J6lRPhTMDuxxcezthg
SSImIFUcOpuhN097L4C0EwX3U3xfKqINUX8KctVz2UxumcQiuMrnbdbEfPMPWk9x
n9voOS+mvUwF1sEfJdzIxuByXBLVpzr5QdzsxY7IYcsxyxkW7sIJlCIWxeZsGtwN
eZsMsM2OTGX2uCXUCMz8wVYjoL2d3hzaVkqPycGJp1TEsI7hFN7ihSVB4qBTFWD5
l9kqic6BWlwA4i7Bd2o2FsD/7A8rJd5smQIJh0xLjV+u2Au+iZzjPX+dxLt9r4eB
xFJ6e1fVFn+mnimPDgJENJaFxXryI54VRwGSX1JPTq1HpfkCYsOnr+PWFEwx3eCf
+bBdD22qYO2HXXWv+vKUvjFAXolnpNK1kBesbm1UQFEH8LC7zr3XiEkF7Gfi8ZeZ
rbkArONLq13iF+AXqRA/ggnWW3kR90cHgMnmqRnT3FQRn0oqh7FV1MbHIF66nZii
0L9T0RBJ3IhRx9jUnM/OaQguyMHQCFG/OGSRXoD3/IdEPdqZToD6gdrysgDcjRZO
U4DIExjr5JWJCzIa4SlmZpVJYLZ/wKJaWnofing0GQkxI37/+ad7UKBqKbfhP1pm
W9Ysa54VuWQ0Dl9b5H4ALUjaZ9ZGBU1Fy3j6kDnOLuhkZyNSXzVtL+vVr3ViOv1+
KjTCEoTR8VT01KcXNLgtn9JjceOj64sgbb7r+11QZ1BQwb6amdWVOuuFtJx9GwVo
7zrwH8/VRgZlBs0COK17xV0GMXOjrdoeLawwXKiNtfHsg84jk5RerHL+U8WPVvM4
aq5hw7N9pp2lGSTN0eksjXNZ8HXPZusdz599hYoMCbbhwxa8xhKXpYTUpjaL0Mtz
tFm8/lhItxUu6tl/RTbjCh5niLdffQ0fhG10OQ4tEl4KeF0wdkcK6o1f50EDdU03
gf2aYy3PobVbSIP2iOFvLejAYF40Boj0w2l6NQ7ydP07T6HDMtRZxvOdP8knXegL
6y5wchBcAIDP7MyfMVQLZGA9ue2OTpXxMYhiAyjKjE9VHn5I5bIFxgpehaPGp57T
l6W2c8diGarxTDC9sDQg55s25anpBFofRr/EbOHtvl0pqCr2OMeNujfLzQb0wRFh
Ul3SrAOx/Zm3r8qbd/HxFbXCS9xgsITwHQI9ppiw8aDHY5ha5r8kXkFsNLIJhuEX
FsWhqhQiYPezudVcY6jBcE2q56jChzafIBTUrPRh5T/QgDFb9upQ71obxmWiYN/M
V9pWzeBCr4ihMh1tWzZRyOjGM/lM3erYCm4mfkBUwSYV2A7xYXXSoihxi//NUwkT
GEpe4ymTb2synmb0LhRwNT55l+ysd3MWiGi9eddftfFloMzpKXb0yTLHOLNnjXct
E537pOiSPfitaWeqVZQiPRon3cSUjawG33gl3ygDOpBHU6CIJADeiNQ9qOnPqkwt
4bBRHYQtHCDjuG4mcNTWDmgCr0/tfX+LFgj1ecWutoeiNGAxoOIJ6uaaOWRqHgmG
7AVtoVCTtDcATeb/Q9i4Z6deC8XDzLV8791zQa3KPEVE9FY7l0B4qQ/Y96SiG/Sj
2DqESUwOQ6IXS1kA7p9aq0G3o03oPuIMZ+1pBXoRdWELFX/Zcx8ODnXmlzs0fww+
tH3lt/9FmQoyqQqmqHuHflS17/bZOpIGaZxY1ANf8HWjgKiSdP022gKm+uOUGARN
x1MUUYCa+atIawzY7S+CCJVVo2iIFFy1bwuYCuu1QheWcxLTSAMAVOF6wjnDbo3R
n3fwUpkpFAK15wPT5R37OjDViNHkkHyFu2MxF7UopK4tHgNWPmafSk9lWw1VLHTS
BS+6TF33v6MHJ+PtShj5VZHODiVw+0gNVHukJK2MnwsVFmDyjPEwYrWGqcm2uxrN
hYsxPfhbpcbZCrZMKZeZTW37wgEd0E2QSSipKjCHS7x+IBeoikR5l5VrExFnJQtt
805my/nAEE0hq6Tm/xpCGyujq7iuTDxw6Ul0yUqCmoLWRaUSjax+MHa2zZ1KYosw
yZDzxoYtDmwf8JRZCrk6StkOIsPUen4ppUka2hY7Hz+0wkn51p9Fi3MuhTn2c4Rv
DgoiIIxUnVzkkdS8LTgSryhBB+1mAbC0CFqAEspWOHF3Q2OFQoUYCKMYdc03XGt9
n47W5H8HKo2dZhSJcNli+/P8pQcXg5opL8i0KGA3XzELyShK0NNzi6h8HKDjRepw
gt+eOPdOgx5z18aL427Xil7ppwVmu4hqIgUqZ4vUnfhVYrSS7P75ZrnuueQzLBhr
q1xeemBetYVAJKbR2iZB26A8M2SKd5HQtmj20reaU8nKcgoB8Yu+KkbmvcaT7rcU
I6a0vJdVpvI3YXKRBt46KYui020dABCat/o+9lZV2CEHGszP2YY8Hs5LLN62hOyu
VwvhEeEz/uHaxlkwIIGirhvmf0QsR8ZF5eGYB8NAz5/BpeHAGn9dFSsAcGLzazY2
qVSXHOW2Jc6YMOf6VBeoP9NMZIhc8pyAwbsj6b+WFxOmt06qD6NWIDXTKt28wBCg
sDs8lxlbWY2KVK4QTn/FCWLaFYm4PO2tVzXh+RwcLp9Xuc0y29MtBd7zh/UZj8A2
fJt2RRgOZ3gcZ9Abt4CqpGtw09Cb3Q5qFgrIC3FtihraB2FK45qUF2zkDeCCdUug
dKbu9VrZMgc684QfdxYB/rkx0GHL6ivrs07UpUaShx82gtDiWHWWdfvKkx5P7Meb
Ie4ax1gBUMsVihmhMc1xPJrysNiS4sFR46V3gG9zAy0WqTspGLPAa4HEN9ZHbzen
t8rvDj6JrvRZ0/HLv0dn/LVjg3hfBtIaZXfZOloxIxQjOws1ossrvGt2+87hIet9
tDJhqHxbgM9yqZN6/yNRm53nRji+P4Uu0x4XIsVjT7AmujES76t2d4Yus4QUG/YM
DtmCCXTrs6xlAw5X7h8tzUIjEgn+o68sXkC+ZWi7jWAkD1RZ97ZhJvP9+BqfVDEs
VxrGPYIFrNPUlxo/JN3aLbM7e4s47rHe66ERmwbxU7gqAakd7iPlfL6U42GmqMMl
3LddwEf5QZqWdd6mKWUOndRVwPf1dz7AyYmF99Py90tpgq6iGm9eQgA5p4BdyOpm
QDmIFuXLVkRmXEvgs7lS9euZr8pSCRRmBACa48av6jS6Jznij5QWDw5GHeiszK5Y
oRqMtooKMylqiuLNMcnA72+z8qDIvbOe29Im5+letWMZMhYpJQkUwHxnTiRSNVBc
Urzu2LvCKloSMRT/eHBNWjZsNrxpVuvRu+cpkZ7UyqoYgn9m3tV9lzV+WXSkNSJr
aYlAI8pDwEhncHVEe4acEw6+t3Q6PHZZACD1zxvAzqlBvd+S0FGdl8Z3nOAj10ao
NwQjNoFbkaB6GuCiKUrkoXaepnDZrVwATiOLbJQuo1twLJZNUjSi1SNYXjjiZSlB
tFqiGCnNJGtBhGhTU5yUWP8ZQS7QHhUMuh+FJWl2IKFA6nMGe0VxqykPVG+0X8K2
OJH6Wb1/K4SLSQc0nkMi/9yRJBjGTeKwd8+tiiK6/vW2JnMzjgHWnuWyWQ2Xt1UB
uOqZWGTPrE4TDdZC3/Lw1TastSqv8NksZY/53C6IFWb//v7aRtG4gqOT33McbgP1
FE2rwfFU3fXGcMlPFfvTwTPsIbkZ0jk6WHyjiVfeW3k60AXPDfBPKLWwsd3KWL40
6jC21BxGjasDEUMyU7x6z8JJM1IqYO7rC72rgU3FDdPLBuplgGrOkbwrcMIVAEZf
uOdEF81Km000NGq0INwFiwAWmugfYUTbNuYZXFoGLE/KIpcBLsK0KWBwjSEuthNx
ra1n6BrW1JbiQqDEyOSBdohC2ig+eoa3Sq5isSXrizAlqICQtTWNdtgBZui7ujX2
VJVM/mkye5mKf/aj1iZjBZzkHhchFlIhnJ9SkIWvcgJ/dnlJwdkRtVVdNBB1ltJQ
XuuFxGCDr8kvP7ZG0X143BrByXjdcBPKSKyFvsO311KvD6ACpgO9ssH9CbGrI64N
fehufYx/XifGMRSt39P14kOcs65xS6gMy+FUfCwicUHTX8oDvj8lu0dxw7hu7gbZ
DYAvpB1UwNxE9kT29HpM9osm6SPv17Izd6OACxzCJrtVzLCZ+Iv+KDeo4JErsIri
C3p0oxE1vF8P9FXrDisG8D3WV18MdUNNBL7MtfEpfoTeR2gjlOF6z6rPRikJt7eE
/evbdajYaFy5G9L2q2PwVZCe9aGsCHjmhHuVYYiFD6U4sfal2FUSkE3emxIuMIaJ
Zn44ffVJRTjLPog1jQU90oCqoGj3BU60cTqLlObYjI154rNO24aQYjnNGbNu/KzE
1UlNHdlq+EyEKyky/0EpA6yN2ztDmxaw8x3AU50m1LzYR4ZTp6zkefh6bpro/nKI
arRTT/yXhuWYOCdh1rMrgIYhezcku35eAPVuXi70kxy900ES0MsHqvKJUQUJ8PJ9
SrqvsWVZ+tR3KLt8nfF8i/VkazaJtryKkbV74BF73BiNwO79xrrUJo5/Jqg8Yl3e
QLqdAWuC9PE5FctyrhZUrRDGC7XJlBBwgcISSwVak8kN3ZL8gDh2Y5gaGoJvoOKe
oIwZgt4Ngiwy44Hd9RCpi/MryhbTky1f/vXnVUlpI3CAAOoyspng77BZPe5G5z4T
HkiI1lpf+Da05tXJ/SeDErWS4hjk834DB3u7FzPzIndWxL7yeHuzB0FUGd7DJ1iB
PXeM1Acmd4wxc2QsQLXEWMJYwr0CRsLloVVvgRpk89172y6zDqYNIK2EkfUYfju5
EMFslpbXTMBLhELX9bitFbmkNJtB4GE5UEuViPNWlRqsSzNNxSfTNsUyk4KXe+jD
7dgE5jYMAg+uBOJMHv81yv7V0jJ4IdpI3Z5HjRUhbEpuZHpROHRlXfD6avJ3Ke9p
x/E52ugsqi8nKujMIksLEUiXcFw/CpKs54fKDnhcR3KZJB8/STdIfzxw3lqVFirg
QCQZEdVYTC6h3PhLkOBXzIu9GFETPvv81zxdLeseb9O0lOfya0ETPLmF/T56t3CL
XoM7QPAFWp7fYA+CruSoOOq7lnM38uCVB1086LdVtPtLDsHiHXN3zwUrM5WyEKaH
5ws5fAAToiPMXxYIHO8a1ybHNUi2SSUK5ZlfHRbCwCm9NyCFEpMKJyg8Pw+gKxZC
yFJesAnR8qEVCXatmJttzVyLQV407i2d96RwkEN32VXiUitV4NC1p7s6j1QAXwWC
d6BfmegREpepc8cbrwpiVEPdFOidooRRAzOhOEQVfAwIZb8T9vqwKlZN3bpTvqos
1ut9NkfFGxZ/5Rw7z69yOha61aB15rDLVtjQg0uv63eSOsJUo4R5EzcZLQr1GYI1
pmRYXcN665wHnjWDeMQU3fx3a48aLReZDNHOlT+A2wTWnRQecAYjpcaMwXi0XunV
Yi2ugZOjS7Gpf9qorRzpkUQBGokycRxsf7yIy+YZ7nGSpzOBY+m2wg8dtsKXR8++
v6kDRkPDTXAAVoPoRWgUGjXs1BGgO6x278M/mgNgFNfHXg4hclXd3Tzj7Z6sC4+g
k/H8ZOPNMAG1yxj77ykrSatZBjso2VgsdrzCf7wFb7AGkBmi2pqeMjoCNclO4ONx
fnihfneMPG/YPivg6QkBL+f8KR8alPnZC6dutb6aTAFO0KC9MiKhMwgAufZrKfCa
RSjziQWO/eubxv7SwZT3vn5XdNQfkX1tMPAYm5EpR0WRsol9wV41CErsXTJl6YKP
HvoMxlUfLLX2J7tK27tBQtSnlrs9vGM/2nO496Dp4eG7L8Ee5H123bvnwX8UZ5fW
S5Y4qeE3v2W1edI/8jrc24SMHbtr3IR6bEU336ehlKkBoJuJeHVAQlI1xXDGG/oH
T9jMWNkyb/ToSfcK3Oh6+CRR3rwEaj64VY9Gj1f3DjCgG8/mKDD7Xbc4m7/YAjCo
F7hds5eddmcGR51Lwt0RqNFDRh5Ihevj9DqV5hx9+Gp1iV8Pgcy3ioH56v2j0C/Z
nyTGZDiQVSnuh/xcbCeGe7oYKAUKBjYZTbwOsZjwAHxbk8YFbRK1CHDeg0qJnAiV
cvmOv+Ch4rZ1wE00DavyapFXRI9griOkcvVnfvAzu9kRDV/mPt+5eE2Txu/lBcjX
HwV5D2MBzTkIroKGDZHiaYZMZSfttzFwGCxFtt4Wu1STbmDVIklXAAeWZvLBVKqq
eYaHReq896QolR4yP5ZNVOH+0suD9YuNxdnj0ED5c7iEYnYomNPBwR6ACfgQS9ZW
wkFoWmQls2wPxCJzdh/toLi9cyY92BcQ4uvDKHnqF/Pbch/O9O9dvpwY8g91hTWj
0R3tGxx+jc39XPRAqs3yhgZx69kkFGJ9q5ulEhS91FnknsSr69hjYAQbFtbr7j+9
HSISLdPVLWpJK2FJnxBDmwiJXMb5KJCxAO0pCbf9CymBAViTqY4Emu7PcEPM+C8a
HcDv52iOkgu4GjUWV/+/4pJXo9z4jPAH7kX9agYlJhpe3NjPeIUDR3kA21h73Thy
E2DAwMmuCZprNC1McfYrgbN3Knm/i4tCVhCWiYr0DdhRLoubgIRxowtjPj/L0bVn
hspdHHuehDYzraTWF3oBWKu1KsxZMpjCe3JizGmSN6rvLIcfz7ykpMWmI0HuSX4w
iJ3/Ue8MLqgCctUrO1q22mllzkldBrZnb+mZH4T07oWSo0zQxm7xwBJtMgl+ietB
rT1hszp7y1DnZiX3muJbZwxBpSLP5gLPWsLNHMfjQZ4O2jYLZIiu9ZyU64666v/6
LdDVbWZnfx6GaZuVqYz03ktI0byUaa4XhaPXxcLj5ZFE7SnkggYaND5vemXsRGPl
NoH530kxdlvAatwS/My84dF4h5gVQs89sz9h/1lqaUmvTeMu8ZRdrGiqKjF9EEZ6
bSX7TRzMa+2Ou+3H6/9znsrlPhRoCPDlcM+8WOThXQQVpgNyxaI+2Td3Xk9aUnf2
t/+7hZkBAZwKOuV7bhdYV+nlb8NxbAtgSFiVGRR3bqykvju4qb7TRGI/nVHaXzyJ
LNNgoAnGu09NFtjYQ0VFEvlLeFRRIxlJ84yK+17h9E2F97VJOp+FUBglVbwMeprB
2Q6cMxeWPPHotc+8MacH+lf2qtbsiDH05O3WvBaLseQr/U9wY5zr57x47cmC+nUi
172Yym+RdhJw6NFG1HytI7ydBhBstUac84tw8hvZU/KWTxElOH/S6vBR0hAOjwTm
y8kBITtZhj97M4DNdw1Vn+otAOZtOewi/FIy5mG1MvVsEELAEY/GIBAk7f6c8L5j
7ojTYzlDy2Sah6tgF1CwOL0W7OguFfwdnKblkdCrF89Pig/sdrzrAdrTKbNI1xAz
fObEnOPEAV3w+01Kso7TZpLFJsBLAl4+ohQJin5rrGdYuuprWqSfZBy8q1h/IzU2
emm5jHX2tVrUkVRMXDBgki9VZDOOdqUymBvs/LA4ffVcwr4WIKZyVFn/PvZHsPPM
sCCtLJ1Vk0gQ3+gU9ccpTmt+Bx0Omw5prO3dv0uSRsAKh4a/O3PY2stxfG3EGV2Z
ZrDHA8oxsCbbw3mFqnkitRt6CJ3JnX9nJaj2Q9O6MJ69WxsqA8GDDtKu3r5fEvRN
LYan+1BBo0ANlw9Lh+y0NBS7ggyevmmo79X6SGQfML7HTs4bPhnhDQy4hJxF4HJ4
nAilMC8bnJcr4GwBb9Glgc88jQ7vA/EQRsel9SdOj2fizh0EgA9p5zQahtf91Jw4
5t0SXUHhcZHgClKDtGv1Q3LPhAlZnqsDbS8LCfQP+G/eILNSeuE+OdumoQk1imaj
CXVFf7MZHJKquro7ox7buleMfaSBBPPEYHnut0L7t1ECsBWOE6hbDvwIUy7lvoUc
Rx+Gbum1I9SR6fRavj+LeLKOaNGPBb6B3YNcOa3Cki7HnoDIlcwKzWcXIMBtWTNC
DqRTsjfDrqvM7TXaQ4bngriv1U6OpdZvNCVM3/3M8Z+10KPeuZpKcgvEVTT3xabe
97Odsrwe1keSDv2qDsuF5By1sZEy1lkRFpTwEtlL65Ed/WVpBXmpN2LxG3x2MUSl
cEjHhFFmN5S2GMxYEgyOGpYWn5KkZDW6vs/2wmnYY246LuMH6HVGdW+ne5ER8Ar/
YTpQylQSbOYiEWICMWB/AZoJof5WltNxCrWFKDNtW8sjaq6PiojaNQJir+qVdQbk
a4a7Pu0NvWhOqkAJnbgu7h4TT4PL0vi/+h0lz9yVFTANKoG75yYeZt8SmfIuiF+l
C7u9DrKs22HbLz+mNzv0dZ68aD4haV1ilS7uEJq7qsp2qMikU1hMZIuJWW/KANjO
ntk7jjWo8LayYEctkoVoDw5mK8NyZVQuqUJTcPyO5NJeeZYTz2uy5gtcZeY5/Cnd
D2sAWUorX6N+H0pmehRFVFpS1siEVGwKvaqZVTql89LGz1utBdMfzRE/30L6qCmZ
H7EvBoumiF3byuJ+v/ajWS3L7ikBq7w1pJLYF7eRDgBhNlbogAroApefr0a1PmI2
kZP6QquiwsKsIcxSu3giSVaMyeFBjEMefMukzjmWrfeRUkIu7oSo1iPUzR/Lks84
otG+lfTTE6JKJLfqBWWvAFs2EKaEn9UNLnDDDpyXpFg4u3uWi3Y10+bO5DNFb7cQ
DA50CBP66QeB2aHOEUhImgiqWRDSgxLIfKqqwxxkdAN0ji112w1lGsoPo3QVsl0p
9u2c5N1RlL6VPk/14pR/1yz6DoHq32x8p9iPpuT2NnBWS8cjAU9f9GFIUC01EzTl
LiSgichXdR9fOKZBXsIlv8sR18L8db2NjTTzpdveV0g+/kzBqYD414Go+RzZR3V0
lyQylMpuWD8lTO6fK+UweiWmw21gDiuZYg2aP/Xok8G+nMi4qQGgGOM8l69fuPzy
EzBCRXq403QLU6aMJVQdvh1DAxGN38N5NYnhu8Awm7JJqjC4MRgRdrZRBwc3DnTR
4bYT30M+q8AIJGHc8U7zfA==
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
U4DweS/EANJFIVnOAUKo0Hn8fEh68YoRThMXFgLmJ9MCTQJCaAaIwOmbw+e8r0qC
bVH/JD9CRSlLmWRLpzaJvDphUN4GrnMWaRusaxSyqGlzXsokn6FQF/qIoftUdatm
XTT9yG9cbfRa8124bU+JqwMt4ncNU16qpkT4Fc5ECaQrzwCVEqM288azVGLGWiPg
CTaT13DtUptS5a8SR9isp7CQHDlN6OH1kl3/MJKCfbfvofivZBPvbws2AcUrD92Q
20bmpIb5mgeZR4nlsQzwSg60/BIywPB774MpVCsJQBVb5VU+dRboW7T2p2xI8HuD
VBbYbh7P1hT+f6RbsGCCxw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5104 )
`pragma protect data_block
rr1Wxhv8DxgBtSr7tLTkxNDJQCMt5vXogKKrUomVmmfmFmpPzniUVUtFhIJa8odV
orlGZ4Tom/HZ+9bsMjXRGijHdrtm1VNKxWBMIe+SFfaWZPaMEBaLQRdv4pI9ccoQ
vhj8xOtSpQjyE383wstA8929SC3fZER4/bkjlZn5/pVpDxD+c5/zT6vpIc4z+BTu
4Bsom+8UORSni/qNLJL07735XrErrdCxHVIAZSjaHjvBDpecBLktflGqSndYzIQE
V0FZN6Ap6iUUeCIXbOuvEC23caGhl9NIFN/xub7cJJV+RSYi1Oq9/80tNHvjHhvI
Nt/SncNacd0c8qkzI4ESHM6M5+w6NP64VNR+VaZVmXR1cPf/qCjKkliUsP5Amr5S
CkFhL9Qx33eu9rttawJ6z5NZuEUzOYe4qqqvFv2xdjYq1lzd3F+MtO1TRB/CglOe
2elCcaTddXlAdAATKlUAlTNsOIw+sJvN+nN0fMhNQw0alkQJg7VmyoBrFSiLaMtl
8aT89JcG8l6zs3hICaEpLAHxdMCJmKsV+zR2JUlJ+IxI17J4wVieG6UuEqnkNFlT
S4L79tKSies6UPVh9pNYDQmnfBAo2J4svyNnUV2uKDwggy/cnWYdNmlBORrnI+Cq
KiYpman2gDU/KMUwpTp6GoeqONVg6tCrp7JyWPM6jsWjXJWDtw/rKYlge3iRd1HR
4D2nsK/AO4LSUN3dF8aGS0VMWWMdYlojs6OCs7zWm0sWNBrO5VtvGxPP1OBOQ3IG
VgZmHK76CPvoeJ12aG2oYrYEjfuZ8KBosqSJpezm2WQPJao2w3jgzFjtqluffgUQ
YFjDTzGitbl/FszK65vMDEjQLsIGUveCsjCps3wd+KKXeZ+18BuBN5X0jMHIp4g5
LwgUbU+JCwNLlaJfIo8cmAQP6DgPcJ5MUCOLrYjZIYILnIFpjUu73lnyXo7fNgMP
ydwTUPGlCEOshbOknaf3v0ea5oVdo+xozo6DJQVTknNf0R96lqw9UMqFRfdh2bfS
7TevFfx2mf4brWAMHvZG4p+T5Yv80f2IeViacNFJLmcBI527+MCKuP1dxoRrn1ik
HGahJenvNeXosbl0lpSlPOegchaqFWSbZBD/uqefRwurGG5U8SxOmXFP8iAOaRtv
V1vtIvOOX15LTs/uOk4Yb9q03esMwUdgBoGi4BR7IU3xeCXLXfqH5cjAui+AItt7
hVb8vJK/tpxw8nhNQ9yHf/+9QSHTJkBNkbdy/CFIlS2cgaNIjaxWYtkyETLA9py7
icTEQVV/j8j1ARixbEQxtzprZ5DFlOUiSALzRs4waA8tE2Cf1Ib577zILJpDFiVI
lNNr6uNRtrqntEwjJgQEXaANaHHrv6lIErObs2Hs/LsxwLmF+SKIiazXzdgwqcQY
oIe+1YhUvLBOoDwnOSmh7vlSSrt1D8QrV1qsHHcTHrdI2xmJj5ryxBdf1IOfep70
ivECTHjk403rFWwwWSShLH0H+jPakqmAXzphLexBD8qUiina6/xJJgbStrMVRc01
bx1ecz/RBQXud5mMu/HpvT1cdZS2Y2OI6HiMZL5a2g6Xg6HaXn/YYl2c8C0vFyA4
0M1Yjr2bSoJuUgOjTD5gbEKAdA9GUl4eYRF0/E+jwDbrq7mby1R0E1yqYF9GDrAj
Y7rzFduqGf6FWC0oiUPFShR9UFgx2dMsNkdFJcrPnQ0SUmBCu4B+DeS4iCun5NFA
Y0nKJLYWuMe2wjn1Ee1cmpdpfAoiSVB4OeZdvWxpoRai2/wR7ElBPauL28wA40IF
4bMLXoiXrX+OLxnetIL1zrY/8wFh1Ksw/Qj4h46PCyqSuHJsZLLMEYzNVxWoBsBp
2X6e3bGtxFOVcMpAg1C78fsO29ykd3iMj2z2SBfuWNZCqbvdJKunjzXiz3xdZi0R
CKql+yatq0HTMNy+T+lLK0FayeNUC1pMnrKS+4ntEOVRnEcHQ2wD7t0X1ulrTppw
7kTOSKQQ/JQuv5YdDJW7DskkiLQfh3kD3an/Gm1BJUYBeRzjvWbXR3R9Qnqiv1TZ
jGPVEzMONPwvTgqt0630e+l6ewszZwpAaXWGmGen4mzhQ20eoKxkO0JC9wAtr3Le
3paQT1NEd0Co1YAcWSh0AduA6Vo3tKU7PEVztp2pFTY4KNaP7BtrByPcha1hBn1e
/OSzPBVBNYVA213hUXTx3aZp86ACKLSxClS8ihMMnDfJp+JBtk0Y/xAGOpbPwc8b
wTd2Hp7qV0pGkjOy9Ls33fRZayy1B17RgdkH44deTtyFQ7FLVVvnhDrE7QQS9iJD
1H+RJ/jklivdXpX/X5RZ9o6ZIGVL8WLA2I09DL35acurGv48TDWoBtXly4KP5iHS
XxiHRQVAUmS3WF/q4nbi9zUjKUCwk1xbrs18lnQli3hzlZCfD7U/XTRfXScftvVP
e0GmgGv0/yqop3teX4leLKsPJOYS5izZ2AyH5fPSUwjY65nlRCdTVqAyvqNSgeLq
84MEjxx495DELLIP7Q35q1cLFeK3eEe19OfhZXxUSZFA8PQOCFs5Cx3PtqZnDIHJ
m/SB1we2kDx2yV7ShBPA5/dxfuS1Wa+Dy64duusVw81rYkG0Itx0Vz7Sx/+gLXEm
N53VjNaD6SyLgogbcrQtZfaW3v3k2jS4pCQY0fnYuBC2ld63S92ZvnUZPvTrrhv3
dEYxoZ2uz7Incyb/sxzN9qXOeiYrHADToK6AGWOimLuN82V4yxrJGt1CszrgMhmX
+T4R5tMlFP4U8JJlfRWV9IEAzoKgk7RAMEnfNYBX58V3Sk2DtBw2nWNB96UBQhxn
gPPZBlHWkK39FLPv0dGqWjmG43hm67bCwR8aI/9b8oqVA7p5Vydup/6k3cPV9j/C
W9CyupPo1bhynCK9vDllJlfuLEVAJgWdn6mVMxpj0K4RyNBUAsMHplR9ijvHmHgG
2qXANVeLMMBHQFlSW8v57FZp39nHY3EzyrJ+9lYqs/tKpgXvzP7xTPVqIy9chZs6
Hesg8r8NPQ+YSzrmNBRQEjvts4d0rsfSV02rO+FCuC4aJKBo80DvGcuHLQkU2P/6
jvDe2pL1X/qk3ffNnf0QEl1NjdwZW3m1567Io9VxSygvYTDKwUcfukDmaUGyU0gJ
jQxnILaCn1cnT6rSDoHD2/jAr483XfOpT8qwsT7jWlQNaC+Nn05MuevcA0EFCIN4
d6mc3QlrsuH8lawe38GXq4IAgZ5mmTbUFQ9HP4b2Jd1LlYk8c273vGey6/NdF/T7
/CdTEhdu56pynP54rChnM7L3XDueb7/W/d3bMAtN4uNzzND/4K49crWQFKcmQCvr
3g07Wv6CHttLNHyMyFwwQlMhEVWQtAvz2+rVs7Lv89oapasLy2ozZfzwZKcAxB30
ywmDXrmvt4EVT5UcKFv1lxSflfuaXByEOODkjOkGodA2+4hLmgSNBQK5IXyp5XpQ
aOXQQdqWsbJw/lgmAdgZzTA0h4bzIlDt432azJ90I64imE2z1L+ytC+4sjE+nXEf
0gmpJgb1JwVbj9kR32Zwu/7zvuk8wc1ZKPWjh3yEGL6xeYeP8bp7dtCa+K+ZJJZk
H5Tuc61DHoQ5L1MyIHH17023d4zUxShQuY8IYqui1zLdkZMOFFxIWHq67KPzYXQA
+DN2gX2T3kx5ghk7y1NLL7FIZEPLdytp2I2sq54UZZxmaRcbPrLEjwezzZelZDJw
5NLL9u1T2HBpW2qAGUvXL0aFaUeQRqdd1zFH9vwQ+bhkO7mxFsFiDTq6qG/2L1Md
zlPtSwJXvP4ACeCJIAmk0y02X3h8EGSVyLEVCDefbSDjObJ5vBcqXSO53sGKJnBm
WXbqql2vP13T0AtfuFwn/whm4iv9oWIy38FbCg3mQnw3H4l76aqLqdQ6CMHcJ81D
knPEX/NnUzPzFQP3HKGSQFg6DUm+GqL9ddGOIXelglWCuRC72WfSLauP2VO3IjPD
EXKhYLkmCfyMnhyN74xZNGSBehbxoUOA72w0hxWjZEC7s07ZtMODFPecLv+8Rkdp
V0wf3keO2zY4jWrgTXG58yaaeUtOiq/G8qj4pTiwsS3H35ZQxw105gaB/3+7Uj8g
ILTDFJcXQ9QizTGo45lYBS47oTXfx+cY1pRwm9HDGgabJFopL1smluzJLUvwrPQ4
RnFoMv34fOqimP6pgXtdGErkRh3Tk/PuQRaWXZwURH+b+k7Vy95YUqsrVNCaAKcK
DfVE9fc8TMLQkSolYMYFpPuAMIigXnYcXxR1DqxWMfxI0NHnbcXYkxdusJj2jBqX
24VYdQXIa4ynI94GMInOxieGrOKhB79JN9uznzPyKfb4yx8FDJxBU9rMsCi5aTi/
AErmqCuKXPiiVjTdCAaJr2QqryRiZ1uN/MaqBjARyT+bWwwr++Lx3O3fNg4KPgHe
GP/dgMuwkKoIbL8BYXJ2l2G8AbRiyH2vR55oIqQQTb14a7yW90Pl+Y1oKGtWqoy6
KGhhUh70n18vDhoe4vbY0xZMCGcp11DAQqGUFWX29ElZ5ebVdJxDaxFbTmFlFyeb
kF+YBTdPWvwwSY1aYadyw7eEVP3repLDftL9eRrjDTCpz1sRSq4el/Zt44kBHW29
YTlZyGT5FFu9ZkxuMCz758KOUhhO4Jj0ljRBDcnsiKtmgpb45EIWvQSz6TRlu+xJ
F7MtyuCjt7yTCgeBCMbrsAlNGAsyqZmak/M38QhEBcN7WPniS8wnUh0z6a3vCJrv
MfCDntDk1dX1PGnQ6cD9Xh4yyDabzhmuaOP9Py7AxF0spIWXIsHb5OcgAGsl8e5x
iVtPXRiWCK7cohZSox6zq13+uzGlqJPD35lvOuaf+haq4MBi6LSezXx5E7GTpqh4
iRjREiEMO4NDA0kcH7fs+4hLL4BU2+jSiVkIN8AREsRDT48WSIEZk4ohs8N30ONE
ZqbNu/LA77G9v6UVfTVSrW5WQxoHYc0F4wp5wTsc+Wl4bqKoDCB+m+ouoJsYcT6F
HUGucWdC3ISRzxG3pJ3NC2Clhbm2aGDqw2YI/wB97e5M0AefU2HOlI9RQVSMevhT
rLianqEVlc3iQFUT7Ox1q6IArZa/SOzLG/S7BykUnUGl027v1fkbh6JQpOBT7eQZ
pV9mSQe+gcLx/93Ih4jeTfb153M+yk75fxPOEpi9JOsvXMmHde9Hzwzyx8snrf6B
sikUrVQzc7bP1Xjv5d3IiGxewai0OPTZe/X3IesnvvyVACsNAYsThXx8HjPVfM8y
OgLO3UI/wDrQbzxLFVK3jWu5tGE8jfVWC+2mo2+IEI/kn//sHyOY8amnr7aYcKgX
F6pva30v1Ek+vVA+eZUGSuypZnfd48xM9+4r3x/kFk8bIKkKBZk3BsqPMWLNaQUj
EgeSCaKB7x35sYoda0P7m80J18EMH13Lg02wTSeBzqIJUOorDM4Mwjx0CftHsOXw
5Ygjpc4h9XYjulZ91u2d6OWC2yzt6Nybjs42Riir5/TAI8OWuFOQccU0i3L79lt6
yMC1+cyPBkVXV03q1BFHyOTR0oRwOCBRFtMHIvAav4m+rWkzE+7mSG/6UkX/gYj/
ih7Ws+p1uH8swaM3YdL4jUWj4p3XIccO2F7otuqljsRUD4F6Xg6ZSKPq4UbTyyqG
mBuZsDTBG9E+lh5NKdaWQx8duNS7R72P+14KsVE4FRZmw6ilHiNCllSncOwpfuPT
7AiUIPtALi+VxwaCvqnwkQDEaY1NuZ6bZghh9XpuXVb5M6ziWmKnNJus5/tYiO3/
JnNXAwg76VKI5jpeLAuqRlo717sa2gC7XqX/M8ynWoMl0kba9GkKdBTZ7NAGYLO+
zGcH+99pc061/QB1GBXIxeqsW/hh1mqnGsT7xJKWxddeVQzl4DwZy6nifcbzvhXy
kqtQr4xediz7NEqvlqit5srNs42OCM/vBSd19VTVgF1xfogTGlShXUXj5Y2FRQ1G
T0u+Aac7o8nRKoqcXf2XGTuMPLYaExG+MfO+lvh5L2oszTuWfc3tfAk6hCFQJD/A
A4t9Ma7rmIJwLkms0PANsNVuih2R1tJqoGGgEyt6OLxc9Ed6Wil+6EWVPS7e4wvR
1cwYd+TxnxfRvpCm0Bppe6bru1OTtwfYkH/buVFJBCoIFN5ztQ+PZzqfaB/9/Z4O
XOie1QcdBPn+dBVTFQqfea0ceL+QRSKmk27t7HHR4wNQq8S6wBNENxLUePw/lzy3
yuz5anySXg5OhtuvQZ/2Ib45c25tdXDiu7C4wPkkNWP0zLjiYvq3CbBiXGfkCrWh
WioCWbP9bhvv65NhwvYncUchto7vCpB6CyMlpwaErtdYCotV1EY/epVHT46th14e
B7JOWFn7foe2bSLmbYV0vwWGvjhgAo+MdhjDccaqokxNH2MgJIPjzxCjAFCeeu7x
sdupcrZaAJOXc2wC2v/SsJlJ2BaebOtGEimXDmXk1/Dgq+hyXlgQlPSvxz+moBuI
GLa88o6U0VZbU5+rLwvaGwAch+2csLxej591jsp7ZrlbKjLLL/XGf24Wa9a5uQ9W
TvQ83Dlbv3RV1k2ejSbUsvnvHyp4Kh748m0N7A9BhV0fEi0hI4wRu3TUi+0spWpr
TQkrsxsHph1lkbs+a3QMMHFqgptmmYuQ9XAlKFS4WFqx50nuq6OX623wKcwBQreZ
8RiGDQiuIrcFdQDkpWjQrRkHDMYY/LAFKjOyqQDKZlW0zVmq+Xpx2D3aTI+B1jNu
/DNlzdoqXL3G73HtmYd7pBb8S1eF9DQNTPVJ4ySmW8NHE7l0NKHVkzkxsoba+43p
WnUDerJUt5QpZN02twywIw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GJC7Ikt7Pfo+azT28+TqStu3kM5Ec6WTOUl14mTw+UMY+/O7ozFdRYO2Vm+CrgRn
zJAQDFNHc1VF4nd+oPyX5DqvXU9N+HxLf++vcWwPuXtuKvKeo9XCLLvJk1DivAdo
fi2ceH5WtXWc+HbVUTtDnfQ/sNIzxUMSONcofDMjjrJt1Zbb9528UqBCARqcgmZR
MUGI9WFCVSrtvPbodSQYe8fDgYi600HkhK2C7cTg/3/3riDfRlmbbAuL0uhsLE52
6MGKoOsCrvtexcyFHLsF9KNEcHRfBt3/INS0rhjxLTNCyhpeuLtLZecuMxI+rzoF
z2VstuzxtqfUILvlmJLgSA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2624 )
`pragma protect data_block
MrmupNOsfRTjDCWBUltQV9wThZfCPcNSgN8apF3E1qsemQLzS0gmqkCS3LmCvy2D
FtIYWHn9m72qQJ2ij4uVxj9UYkBU51iGptScGFUM+Nd52w14Bo52b/ZiX+ZPgYaC
QJt/MW0fU5y/5jQKf4qENDLNY4xLGg3NKW+vAzZbuiaEJydTwKWP5MDCSsqIHPMn
zVzBnPVvuJELpppIlU9KoqQIJr6slse9aZAlkyXew0mPGnApZtUzWu2w/hYpQS5K
kTlgp5V7tcZOYOsqGLDjvdroqUfe61Svdv71xKIGb9rsNk6Wz8VJpXsF+1yUUHV9
nH1j2fy0599o/PpSbyllOMx2wF5mge9L6tM1i7QYiCxbu9Z76ulpEYl3Pl5+PRHG
Y+f71MLgGClyvTXaOlcYfOXKlSG4+8iPHoMhI1WQ13cTmP+2PcadEWqmmG5BdJD/
Kuts2Iy4Iyk+foMg9YWlJIexVULOhJ6MDKG59eZYmse9kQT74MbL4Wss8znoKhww
fNoaAlTi4vvL09jwI7hxL8njHn+7C9fno4NCxkI0OlFj+uNt+Bv+uUtLjk6vnEBC
qsFKLdCacb/HWRnxGPWNuiFjdsGsRCLZeBc+SXgNyHOt97/jx/t8VBV3eT+JVl+e
J7bnNvRrtzivAinDfHxWlfToTjdo0nioOCm2ZEENw+3NB9FqdfZRcKiaUL934Nwc
8U5QTG7SUqPoKV5y3GuoeE8R9ncDqmc2WtYrERIEMSj0MfepAFUkkZZsDiahqzbD
I+BAJQSOxR25gpZXU3b89RdF/pJ8Pp9WLhLfiKXlyr4PZjKHqdNeOE4VyJZJWHOb
CVez8TsBG3s7lIuMrNxhuMoI5NRqOfwCBGvAysocN3f/5PtdvokLqZLlVS3rMrU8
MW+d98kTO+2+7ikw2BnH8HFnH6nXUkbd9At8vSNIAVUENMw7GSRew3hMQyY2Fy1Q
j1uwBmE81AlGgb22ciQuAXVrFmEp8jU7no4t0jQr0pYNZSV4BQzIjWXyHWTXB7vo
giORCRP2qL28544vpbrrNQ5poImpsyil8MGom9cgxdRQrx4BBeqWKabVkl0BXykL
Uonfg9p4yXM1BBSLE9RF8b4jlvEoTiQ8lSzymTDMIcmD39vpAYEI6oG1HB4Mo0Du
9q86z4LdSHAkoCtmCRwD6tVXAGGWEstqyyBDzoNNNRA1A/LAsZulCjzxsV9HvfLJ
8NW4020QhGkqo6KB0c6NwSWfjgzumhD1NYI3E3LpHFPi4xLHcurVqoaUu1jlwhaM
DZhVSyih/M330ImD8+Auj5Q8iefuz9xV/TQtgPVd8G+lLeC2+MuMd3INf99qNQx5
dVAhoL7w1pXf2XhULdq3lDi2F5aZGy+gCVoxIp/p8XfGSli+cuqjJyEWT+wDk0y9
8C9jWpZ1UnXetAKiBHwoGkC22dbuZJz/upYB5LuN8nxUFAqkQ+maJ2P2rmHrK17s
xedyA/d2KpOvxgjd5RtLqaDdREAR07TaP8rBvQ74MaZFQP88Qew63+eXm5nwqJYn
Il9lYYQN4Pj+kl6U6D676rE/m6VCHsk/y557BF92Pb2uw7UaNnMPKYh1nyXb/1Uk
gTn6kG3IHqvtkm4teSTe9kSxL3PNi7jMSG1MQlmtZwNSr9BA9+fDA6Fd8K6CVLKd
PDfwT1gExhOHm7osUx9FW3iAewd6JeY7b2wHcaa7uRv6YXQyrNTeGq/yWNQjHkgG
okZWpSM7ALJ4O6bP6nKJ2R6XDRm8RtdcBBdBTcYYDUCiGasOjA6HlsQi6YkOPrxR
62IQ+/IDOVouYpB6LHV1V2PfLB+eb327hpKIDyiOVCODAd3irFDiTxoIR9yZQ+4r
UTbUh2O8HxPJSgUgiA5U3v24qfJrhce0YHHcV8bZQJVPYlZZn656hrZ0r0V0PbNk
2oOsB+ZvP95HCVjnPG2VgItonqvSoT2KOus729XOwD41G6LMRQGEPHeyaC9lDNJo
hbBBArhsgQv7ILCrUXjiWSUlVucO+RCD339BPzoB+Tg9tHtpjfVDjwGzFHZ0gTgZ
xGZFKub1vK0z48nzSfeZ2LmSSZJ43JCZi/is2lNzhZ6JNUtlxJRgpHRiJ16gyzci
EYiihDiyigrt5APZcq4vszSOq0+9vH596Wma486FXTekx2Ykmm9LpuixbmtbEHZ3
mTggV5I+PCquBW+3kiCvQLZIlcRdW5QAcYNvYNNvwieHrg1khbVGD/83YQaO0rNp
ezuj+4rOlXMKtxq2jnYKx6mErpv8Ob/tUor+lfhoceHmSrbXJnzK0TEqsSN+9Jkj
HNalx0Ahg5MZenRyF95X+SdC6YJ4i9NaNOGZ0EC+QbT+Gv7ZsqisQgR1Jaj9taYv
JDaoLzcFed+ZPBRAeVixhEzymK4ZyWDqqxGBjUedb7J9F3jVY6Egra89l9cfQh4i
swLZrIgDKpKelFy7PIqU7i6y/eF6Dt9v4a0Yx9YDSapJVPVwj7C84MDHFgz51oUT
up2IVmvbnO26rmVEcWzefxqm24aWTWsARPd5RYvxM9Ugzq5cWuMvfQPuMrZ1mSlO
B9ZAXCFt1Du0HGx2xlJ7cT7xpyHOsjoDeHC3pefk0rhR/NFJmPREA6hOGV0cMP2h
XS5BJncAm3TNhbKeVzpVhRfXLx/9t/GQhbE6S6Qrjpj2idiWyUbjFmfOPy6X0/LU
fbbz7HSi3yRIre+hLqFH63DS3KPp4wW3nHex0iplTQOdQ+/zcSfIzsbdWsPWsYVW
/5EsVZ7CA5YkgWLqb5h3R8LkeOxlAMu3PoAwvIIaqCl4wRWkh6g4kNQQH8uOCtnO
k9lSu/O8/ZeAJKlpvjf6FOZ9TZminhvM32uV2Zs2BM9Bxcj7+64FluvUc7ygwkz/
+wlZmhFjbCjpMpj+rEbVdphcuvDsIdlS68WIIILowbCwNaQ76Zt5SXYBdOdBsj/A
u/Q9AV20LvFDxlJxG4qQbKjzC2Dl1b060TXpxNn03nM3orvIr5J9n7rW5Fp1gKUw
b0MHSfoVb/ayuMFxBpMQWBQ6ZsEwsMpyHh9cslfcoln0wXrDABa+v87rOQVOlqGI
27syhx6SAtWYepUAogQcU3opFhH/LWnZKT+TLGxD1AqR7BWcHG/i3DHMA7UyL4xM
Y0kJ4xSTK/xqqm21PUj/TX03aQLzwhkbYNsyaYbOPKDrgu2RHDQJKp5KuLEuhdvq
bEa7nCF4IoV4LQIrq88z9fuNeQTSbJnn8IC8npF4ThhSdZhuAWhCK2fzW0+hjNC6
vfaY/hm531San8RSEZzhpTMU01i4GKjfbe52oMu4t6dz67Qui+P4hZmRorPbmIgX
LoFUAmQRF1lMHJMqoKYx3eNg+sn91wb5fwhkttEzCbSwrsrV/YMtCos6evxVYySq
Ki+630QkC87q51KUE6HaHjQQKvosxPRkLPxlYo2Nb5FUayHnftmLN9EmdRzWJAoF
8RKRBIWCgakwU0hqozP9MOSmV3dRd1AcAG48Aa2lHg0=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Sm0jjN+I3VT3DuOcGmh35FTdHo5cEGlgLcRh12zHoez9KAoZc4C4IRizsALrjHBy
hgM2xLJP2LU8G42rhf0eKTUMB87UEH7+cXR1jVciWYLZXIbKg1oyeZmixH7xyT0V
E2hCnwAcmJIBfHBQHlFYW8aojXEst8fNmgPKah5TDR3p21Hzu+GUThFHvxPDrl/p
JBcC2n664nDPCeK/woR+Z1kf4PcFm3sD8VxZOmWqrosUeTCMffUsp4iewseRJ90b
d/lQjwSzbn/FR571TkPaG1cooewa477ca8DdGScYqhisjoZ3Cilh4mTjOwTYYUjO
1O0OXqpvhsxFkPlJCKOl0A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17952 )
`pragma protect data_block
sdKbXbzMR8TkfDXOCACSbD6KrpIhyqVfb3O5Li8pqGa1H2cUPQlLyxdYmMC7P6ef
LrWRgF5IFOIr5tQ9RINJXaJBk6MZBww2zZ16QPvYdkFu1brBJqNINz8GmfaaFAaQ
NIKXa6nQ4nUoOP468y8/V0jHodQX6m65jKE00U/9Mr+uSUGoYffQlEkZLzR83IlW
Z7gJk6BY+r4pgWdKfF6WLBYTHZCUDUoAV/f9OrEA8o79E+6k/iyaOUV5KTHpXctk
lXTbsLuT07BPtp4dxRV6vJd6hnRot0gkJG9U0AHL3CTrdzhvP5SiDsoWyfV2/XAG
IRutAS1XWiTPcvdSbUvYQZ9sQji7J9dyPPeYLoN9KwFcAY2RJadoSClB1fXwcTYu
/K7QolLZhSOnZpweTvgvvD3jfP/XVtgovAKV34COuOtC3oJtKR1As/eb4MjE5l98
rGpD4woOkiQr3zg+zAdo7HcOOycbmzMvMPzfvYBY4uBuVcIwTdBbdUIy6xTiFI+a
Rl2TG7foBuRUXwl4bSVqe6/TCUm6BO55M4FOTq+3HJZu63a7NH8W9+liVDmaTqD1
ydKO7uuKME+UYFkJ3RsPft3yOuryTE4VV2t742H8tjEKbAQKhKBBy8OFVrTwy1LT
jBiZrFcEfV/Ce0Z0tH1PHyG6MtKd8eRr51nV7DrEV8D8eYsuRg6ptwksQOijWuA6
e6N8lIyzSyQ44toL3GAEoCzvzHbW47PrC3s7D5w10lxrfYI/3TS49Ow/YEM/RJo7
TeKQplqY0dzybClO6Ir/dTJ3UgC4Cu13UUvKuvHvPTPtQbzVurCufiSvbSrjpW6K
8iyIZ04sLhcwSGMWUaY8BUeZ48RXyG4Ua2S0I4LiIJxGHdtqWYA2Nheo3aKy/T9K
vN8/32HRmJn62f8L+g/lgcnA+ZoHO2JmPBwoHs2pfJn+c/msai8sbAKqWWNhXTn/
9LeeeUqRTO2ubetva4kQQT6fiiWqxiDI6RBeLkA+VQQqBhYf9/yn7aTk/LPaYbT6
Mo4y07AMdaG032oclJFcItflNE4bIeJOGYNKDQc7s7ld2eoyBlIO4uaRZtKrVA9l
ntlGhCPhK5sBX2PWKth6l7ORf4qeehrNUd8YQnhlrkC8z+hl6w7XK/EQPPT9gyep
ecikpskoAgbH1guKw5tbpRJPSvvSG9AJBJm/1Xp3C61Zqr7Qlvk6VLcso6s8uzGt
VghE/QrUmVAyeupWE2jWkiQeTCTN1WfaO/kEhTmssHrVKyPY1wjyGJacLiq/3uFk
U3Wh0Oa3Dw0UZs/eVdJVkFMN46zlChlGH0aR6ilhZvrojdOWG1e4SAAcFu7my6nT
tG2hCuT2jArhOJZ5fIRk67Yg04VDuJP1WN8J9FumrteJm6GwMgEjmYkvlNQpXmeT
3G2GRT8r1LzWxcFP3RBsGkD0K+Ni3YyK+eR8xF/aTpKEJy6QEd+LBSV95EZ6jcpi
XtQ9EhMX0jI0SizAm8gcMCbOb5SD094Y9BNcwUpwZUMaLgo4TPjMhrJ+4dfOe1V8
DJ5weY1feg9O1QFwxE550vfeGM4gJsIJPS2jXdH4H1cjtLfvb6vel7jowvuihG98
rhcWf9FiujhJlmfb9JTQ9RpvL/vqa0Gg4TSeicek3Kx+v7DYEXIFliLoXUHgCNvv
rG4UiNyDlGQPvSbtX/N/idt0OJ2vP87hKB4TxVtrETIgwDSTiA1OQ5Ij5eaTwYvL
cFYp0lVEn9IB6/dyHuL+gbM8squid43UM6cymWLNFU9ObQMc+UFV4VHGyJz+Kzjk
tbFY3pnXgqfdN2V6YsQZaZ6mNAEaAprmeLRCkUbnT9FdI75ofxyeNr3KjMNvwvkB
TQDC6YE3Pwkh10awdr6Am12mYJy4VY2M87iDqkdR+kO5108FXI5EEnol7yiBetUC
7kxOwbJvnC4a3iZCA8YXRFAGgLW6fODUrK3TSvdmYtLmcz36kieeOfDMKX5BjJQY
nZFvGkjnKQ4gaREd48FD/OJBspR4RdCPsmNLU+9Iz5ybTgsshcib/nfmR+K3QHr1
eXjVO8tgiuqQ8GrHDNULmO9mcGzmhzy87KT7Vg3j6tl3mUtHDzQjAxX6uVnripuq
vTllp0nxrjqQ9pKIxmhKBzu4yVNmWMzXGYoCazcD7Bijb5AhULuP0uxRQ1tiNT+M
3+kLrCEv+LjkuBGLWWe85YrVIAuvnEpJjllvBDxIJ+6epc4veIR/pg9lFotBZ619
dLOtuZfbegvLASDpkzrL4yRDDe2YJeAscFaNeAF1QN3Vi/9Cbmq5kGx48bUeN0A3
XiSNQmsO9jhW+769FiItjSTGXDctwGuxw6ro4NF1BHmHNyAoyi5HURugbRXnAbEu
hua3lhwWaUWaABpe4DUg4htgrFJeowzGHdduO/jmfrzaclZ0miS9O1gxyEN6RCqd
1R/DIqOjpzICWEjBje/tdM5sU5tD4REACthBxoguUa+ihW/bw5bjEO+LQrenwYaP
sqUthy2964sYuTbRX3mE8gceeqwtsvxBfU2c/NMfkIeTA3JAmUKue6FmxybFcF2v
5z97XZEfGIUM3UVMOjzjXTjsev7is2pgkvpS/eIPA0tkJdOYTjsg49OXjqlxK2HW
4Abddl/1KJd9ntRvSu3wPXIweGLvlxmjJ6Wj/dpcW2JMS62Ra4DKjuNZWkxqFZVY
NC7by6PWicjUL0VbDptwdvzgpn6wWX1gkyO9CKKkuHg908H7RSuArzvkeZI802O5
0wx6Q65hfkWa2NhDFO4aLwUABZ0afa1Hq/1V/6ukN3GNmgveI7dRel+PMrF428Fy
HpP0jQhyPar4FPv0gm7LuX5QLRT3y8AUsyKmH5+35u82iZhISUFvn3D9xI7apjO8
5GDRV7jPWTx1fzRy17SW/Mb/ygq58ibnsPFfdzB/AOgiaCJIFtNxsahE1blE4bvL
4EDqwKnyuetk+kvCXRJBwuODcQ7glfpN2EzIgxOH5/5ci8dia/Bbktdkz0bLwk5F
YvIhGzzj/g7l0KE8dVyzFdQQFr/tcuVcLf+DTpAk1NKXCw54UMUanvjbDjqQ9Hmc
Fvj7plN42h5fIsJ2vWz1Kg0M0WtpRkoYHb5/wn1kt3DDX5RyGXmz/kq49nE2NDWw
/0ieA3VfCN8JqGTkyX+M9BHiXHzrqAa2zW0cYc6xlzUrL4GbecUZO4IgZeA2G7p/
0ujeq9BuH2Wj/npoW3Ou57IMC8mdnee0ts1XyJCNCbKaGdQbd7AeWvajG2mC0vru
mdTDQ5qqdQoLkIpRNOnd6hPU1lW3ZMSwpiPnMLLDjV9diNX8PiDEBASMp/JHc+Y8
/UgxGN85r2tCjbVfmA8FBSfYenbeSF9mykWfzsYu6H9H5o7icSDVjsiQ/+y/hVeO
e6p6vp0NwWcEe71SxWHCTr9ToRx25cPnU1V4oM7wumTp8As0MICw8NWqOvsAOEsZ
ddsbEvYgfCiWsJyyC0TuYdMHxXQLWMnM2UOhx8ZkXTVG/X1zqu+f9Pux1gDQ00zg
ypPC4U9mKBR8edmFgmkWK5NCdtdQp3pxjPBb+jUAuc5yNl7bIjzL3CWE3irdjCu3
0fHqLSmjZz6e5V0XEJqoJBvo2Dy6BthMlSZ2wHGfHTwQqK6W1g9ESddiuLCl/JNS
uuXdkLVk9UULXHcgId+afTT+GSNXzjLSxW5QzI921Cg5HDM/N578BssXGRjDh+wF
blHqQq7581y6cgrYn9MFIJdqrzvWwRZg2htcWPX0GSjIjSLV1TWzXI5i0NbJdlm0
mOT8qWj3s345VkRmbVOeXxNyqgG7/HfDLOzxUmFXTR1IY+1kkvvv5O3HUuGQobxh
bJsFNz1RdT1VP4ToWevMtu8e+wWttmwUOh5wAgoNOv+YAZEAWrOkyRJoa5le7bqB
tzzguEkD56sfAYGhweIZ5JFL+eYDDLu8RB5Gt9Rly3Yp7reFc3QBfXsQHkdCTx5B
+701zQW9r6zVQY3LJAXO87gmpxRQj7vLJkaGdzdLQ4NyYUzGDQqR81dqNRinlMfX
cdlkhASMfylBhsGtkacbEGxVAfMRh8sa+6Undko0C+7C+t9trNhBoCh/sqMot1/q
EZuI6TkzlFnKg6KuOhOumSImRrWRvISvKBw/wI6xURygT22KB+KxHqVw9zgNKIq0
TIUps0htpsaIXcHwuIMY7P1/k6DTm3yBge7/o0Y0JBaa/p9vXtwOKlYmeMk1lnsS
WdgBxwCp+i6uA0/XVZcam4bdImS8lGXu+/hgHUzPg5D0DUXUVPgcmjjKgJ13Lkqz
VMDphdpNVdIQ5tu3jnNMRZ/JUDFwfgo20HY1aw/y5DUSN64PAaEW5STJMRhGWp85
rv9RyszuRmpGo24zkAUGcMAhsuIBYYDfvqu9K8DGuHxUqhPdTK2kjsmc4TXQ4sZy
iYG0AQrZsElc7wQR3Q02ejaeRunbolBW/VpWh2Ii1UhsCunuEepJsAyK4tCkg5yO
1EdXZJFsSCXchSjM/hyZG2VHJA6uhZREl4Nrmc7X2B++yxKXZMeY6Y+k/opFc6YE
o9NnZNDccQxg6Fws1YeuIV/DfUXdZYp7nqCJevtN+oSxSt+AvZDQpJ+yRNJ/NU2s
+I4pJnZVvJ0fDK8ThuFmWWz2qSSZ0F4LCoYtQMdfe/cRZRiF+LLkRNzoPhg8WaVm
loD9CQwdBDVknKbcWrn9/eJfVYdRD3AcHuHXE8mNT0YO5ZIOnH1KA5LNlMnjn2QB
Q9VTQoS9jOpSFlupcTyRiN8EeI3hosW5bi2pCC4LDm/0mYVGvQsXtgB8O1rgSkEF
DHF6vG39tcxBQJuDhezd5qTIUrSbdVJbAggd+e63oS/CcAt9v6odDDQD+m4/zVJp
+HJmeOb1/2+V6x9Wg6u6a5AYHsP9t1HXSAgh4lDSDSxg75F6K3DO8POBnSnx2BiI
crDPZf3C8JU55etsDgDyQ3cf3AgUlekrYwI9iiIOEw5+5p5noXqO4dYz7V9BasGx
iNOvVjQ0wEnQwBU/bi3F+gfdn07GWgqyZFr7R7xA3W5xUHhtv4niPyuZCt2Y1aTF
EHTMLzvDqnAbEZ12Q5w0zG7IgG8xGgwQpcsQU0fdWfFqdOt/F6LCOfH7EXTjWVwg
rVusSdbZ/Ria/mGSaZCejQM/GVfLnrAUIcKiXc1+piu3ocol/5nGbBsC4ok437Kw
3pSKVCZMa0KnZoJCKqHP7VV+FMV6sw5HhxNjoxdQLGw4NOilkLlqy1a8SNS58c1g
mpdYp/7mSxFFcu+OJ6Iae6z7pYev/Ss8mPymAsahlQxa58em7viP6hpPzZYrJpPJ
789MfghCJWRdSaX/ksqicjo03yDWGshD0hOX8DOO8mIS+d2xyCcRmwMLNhKAdyGI
zwwJKi+hFCB3ZEFqk6rOQiuMZjGTTBPd+9lSAcevoMOe5vRgqaijO/I/F2IcnU/t
tDjbhy/ZxXJBQK1u01ZzvipadThSqtdxS4iOM9b8XCHTmD0C+bgUax7fV4ZWLJVj
YvFT/czjj0xZi2kAp6OgeSO6BtTn4xDFNDBq1+TJxmFt+/+rSmTufdJNtiTepdYy
yqEbHO0YRPLADUFcrZie+hfGS2z4F+IEHtXNSTwLowdpEQ32c2u3rFJPgt/eRIrt
xtszeJNrydWqzMPzW0aeFpRjSf/2Y5g2aom6wflSgglZO5Rs6fmG5WUwN8PERJi9
SqCkbFiSf2K3lGJpXiwh3zwFevB9dyShbnlGHRV+4TjHJWGR3pUmOesHiLRTChRU
8o+QUPwqY81Gg+Pmn0/vv73ZHSScMIYJTD2mwJHNMFCj62mhRzTwBPk5EkQHSD+8
PRX+vPTwiTzC4pFBIgYLWghCsUZ1og1vd3bCsEtG2rkAeb2UqqIN7sm/Br5INjIY
W1l3FXGE1qPRnCEPU2Dl6YBLzUmViwFxOkhbpCv+8AoGg/Nh+UpkCYXyeyA1QgNM
pCP9Ld0ubo2haxithlD4fi+FHqHJZdbtLXEM1BLVFI3PP710rXPjaIZuzDVWNLzA
rCgIvTUmQzFIZoj/vEwgeIQ13pHD3gzT1oDQvHuG/N07HGxW/ydBc4LckmH9DIwo
tFUiHm9rnF5t+hh0z50Ptqoxk+u1bliWlCiFjbkZFxr08B3Fev8hEnJxRKKPUoev
fNB/w/4A4bhXciJ1pHZ8pEFc1czPS1ILM1ZXj20Uifn0V6hpFwHycOGPoqxtCgAP
CIpYgJPdm5A3u3+NS46KDJ43ORLT+rvrrNgKC4nNlPC1nkGfPNyIMv6lp4O0brwp
T1CNAcLSklZkrhMDxNjznmHOMMwNWDN6/A7lp93Sw/+cL/VXrbf/fcpag59Srw7u
a7p+8GYrZcBvFDty0eSSJiWDfAe3lcmcDf/xCk6b2NYOS6On8FddnQrYQwOjMT5Q
qrtgsme/eATANwRKHSjsGQ4jUl2Wla90G8fgaEjWoWQJV+Ty1iQSkz9QyivyceNq
xjMabMAK69Q/EtxgfYuwlE+6l1Mq5Qm4ZFKXX52Ngpgk694VKKxCMPDR+oV9HokZ
l0SXmURd5LQGzd2eNwjaN3qkWMwo9smCGcAMUFGIHi05fRbSVTCqSVy+cHOGD0AT
QV/BJLnyGDV7ebniHOEg4hFmowBpLXjbCObDkVRQlIsR5X4zHy60R3MjeIwySrLN
emJbOeyGIy8WRR3Ka9k/XMHewawYIympkOzwc3E4sSpY3gzADuazu2rOiS0/P+s+
0/4BMhWLFzQtzlrRHLLcNlHDg5kJSHWaucOWZlTSKqqD/Cwg14m/4K7ntAvYXkdM
FhA7reeJ0nDLuUP60SNnH5tRteCo5xD9hrNn5dOmZMCAO/R/CQJRQginkq5jt6YS
fnSUT/u3Xhuav0xsUMw79TYs/NLNSRl2YT9R/h8hWLbDPqROK8tuigr1TkAyGZ0u
RFx674N2m+F1DD1/orxV/73lFgIH++JXyQgcwmE8r0cKSJUJcnYALZsGNC1lLzdb
sFadDozJYRXwKjHWLHiIp5jWPMkrrWicm9haQovtwzuVwHo0wRM1uf61Vn/u1Uex
7Zeb2Z8x+uxKydiGdu2+8rWAIssxDvUr3aeRI+3dtI1E6EgSb969gIwBEGg+83NL
E/XNfU2iFYmHsedVx+vvOZa+1jwwrGul80BDn8nhl14QJPECCiNggceIioL7+4j5
heP3Rpp903wMz66jyqQRtrTSoeWINWTJS1XXeLSduOgtgUrDiaENJ/kgqIm/oKF8
Mo3gsNrTkHaqztLgUaARzz+FIDjlEWfMANNqW6ZWmZeZCPWW7IPKqKiEbQtth/uX
/l17or0jreo76H+UYP/cEVjSP+2k7jbAlHGzk5mveAtH91lLg6OqN66fsXiF036S
xgRxXrU381EDWjF9VY2Lz5/fpZ7oKR1b4Ud/yUXWIiKuM3ujhHCyWHmWrSgEK3eD
kVE+jVQJAKPS6icYTI3Snz0GMaj6FQGOLYYJAO1rPBoHwFqKx69WaQ9mlJEU/oEr
46maffhB8Ck5mdh86NGBGyKhUTxZOT6s+5YBSpheN+URlGJJHWojvBa3aWlTKchl
fAd11tIafvNgiJr3b29ka+YWDKMhNJI6tCr069pfniCxRE8Xl+6u2owKBQoFvjDS
9zAWy4bY74SINGMYLMzNMp/Yy6bBwsrH7oK0HVl02Pb69IldRXn1yfqKi6Le3wnK
BwjVSQTJvLvDf7njyxYUTopvt4IchEz7vDady3/8tGjxeFgy4sL0bhiB1HyAuZXu
uNkC8iqX3oJJ3+ZdMkVtEuvWn7HWc3LNCddQA3BHUDcws7rBHPZUmgpkjF353Crg
1EZZvxV1QBb4XuhZNG51CzORdn1mWJlCYzGiK92A/Ki3Ka9BqFcOiO/E8Y/Lxx0/
jazViCTp7rZyX8oiotiHD6W1lZKPqUqA+oybETPL57wlAeN421nr9UiVNPOt3Tzg
v0XkwHUcE9+5M/4xZ41Qhd3HWW3uRTxu2YvulNl4y88VbzOCg0m+IIcK7GrYZyRo
/8tcYs2XEByAPVtFsh0VwKwPza85qgibtLJvAESS3lwMVXdDKgyaAYSHuBcSEXWG
aoSJjQG+zEscCnVIVk2xG/fnCUKwQAsjZu3hz6/4b1JYiS5/oTo0qF3bQfv8HPXc
n3RTXi49VpxPbCeLSL7I9PaVAPg8IbO41q87LOmJNKIBMv3Nz8DWAI0HYyXbV8Rl
bzG+CLGDlPqurJ84bUFkgAviJoEc0a3twR7lAGjOOclGZwRb0EdeaPPxT8Q4vHyA
2N59vlo9r9r3E4U3YMppOaz1iahEfdG8y8psKj9xv1JH6JiIBXmLVkOVxNFMYBxz
igVtbsu1hLriGJjaOetBNjtKs5B+DG9qr1sXrWFpTHkmN3rq1rGueiPqt/oT6k+t
juCnF0iXkKYRVibkJnbVMgw25rtTqz7i2ZZP6/9kVqDpdlE0NzLZs6bFv5E9uqFL
rVP8VqPS4DZssnlLQeVB3RRM7cSxBrmBJoHUCwuUNnHKemCEA/K2ZL9ArBfVgnT8
PfjbXBhyEX5n/U2S5fhCE4+QmWiterO8w6j2GoehjgrnbgBG+2Hdc0xMCxBvC+OF
HovBmXIZJ1IoMP1YbWy24S8x+DQ1d/e0nom7t76J/N8LVb5ZSjYj+D8PDXGFLFD/
w8Y9otWYILAJDwCUfM1Ol2nq9Czg4NVH+CwRM4gaRogr0bj9akHZ4enU203KNb5i
cCzZ/gByWsv4hHNcjxjJDpx0GltwPrXnDUCjf8Vn9z1T2Adi5eq7L+eIf3eDK0cg
iqqYfTbBUzQrQvSqt/LJoLDv0kV46QLpF6nEf2l/1Gu1mJI5SxvEV1INF/HGV2Co
IhWfnLCehQ62Vi3cHLw45Rn8r/Nof6ufis8+ZE9haD53VsR27OpwT0rIPQQTwEs+
Mghzh5dfICJUQyRldDmSg6puBxBxKXFP9xQwDgkKFNk+qT8dbqm0ZdLbgPJl7PYE
7Re19zaduGbq8+NoN+jnGUi4s6U7lloZUKGN2ULIvO6GZGYhAaR6468R4QbzFbIj
xjVLdGf/iy7CRX4WLsMuCeDM3iI5qV9NwKt7z7Nb+tELOO+wjmnYGO7OdQl2ruaD
E6AVeEgqFSgmvlzsJcpwI2OEBQaFk6dPtNCHG9GcLt/qyt9K10KkowoyFs0sXhlH
qAYpgmI8NZkU9VOUPwW8b8+/CSLN1FpUKmZaaAsZLz265O52G++gxH6e1DBITLIH
gMC21u1Nfs6L5X/K5WI9/G3C0wds+SLiz/zjKluwIawpGo8PispCgeIjxl6SbaSI
iy5eEq9NCnWKnwYdbI3BECWyKMufXbKTOGRXzAEkxJ80CvQrBIqixHPh8FTjZJYp
ZoLUVwSamWiM9zW2WxhYqlRamd5iEnH9fWuNh4gqiCCorHpZ+LJ9RJYdg45/1vU9
yqYL8lDrsvaQi4XReK7cPixc80SdrYNMt9dueY3KLCjOkz+745YUGOeM2FjodcYk
Cw5SVb+NPNsIhLxIuwm7kIwklFc3vdeYPcAa6pab5j5+LOSOOXUCNc2qMijeBEPa
l2y/aKqr5tubjHC9yzg5oDa6dAitCNi/eN55tbEIuSLz/6AhaPAgthbhc3cPY+Da
H4jSllXh9otT0jcTlUWKIOVgYtypws94E9I4tVXbTUjxs1fm2zMa7uTYA6X7BpBt
v8+mjkxT+xrewIwJHGZKNh8DXOTrXeK1XlN3xd1Vwk89UyA7jUrgKgGt3+576b1j
hiZdJIrVeDTodDik2860pMEuzNJa57lB6T/9It+LUpTTwMq+GqFm8J5dtoAWN2UC
n73JS2C34wxnreI9TEJ8NTGG/fLcBeWyd7ytpj+ai9O/oTEPcnoXN9dBJB5eMXfF
03lITf/V86RAoUP4O34ckVav4qAZZivyDA8EezfM7QiNQh3wHvIdizK1OJ5eZJvd
06po142xDLPC6VfNqLGzDM/zq7vesZ3rv3Sax8c8lQrenBIs4KG3ctT2r7g4n4LC
zJ89XmYhqeVXyAWzIrcpSZJ5iEJlBff5qycCsbiW8P0bNAr0zrC+xNBwUU2S0xib
MSfRpwClb0uUN24S3NO5Cr2XWqxZaBo8LUySViakzkjPnLF/SL5Kc3UBDKOpb4xL
o4kxBQoxaCw6l8c7U7jBV3IhdxsRuXR/eidEyyoQVuDUltFKXGJCqp9NHL0uqswE
V6OQpkX6P3pagyBXUJLf9bmsZCjF5KawiRPIK/PEmG+pjPMMqWYIValhjW0MIXXT
u7Sn/SaKCteZFXgc79vFIfGKNW70Oaf7korV7qEeZuQaXPz02t2tQ5BXoZ9Vxw7H
L79AJhLs2dBdUxLnL6egNN7jABv2gwBBZSsDOMYBN9IWoteM6p3Cw74CRqOAjv6W
M5/pXRKI1InvpJIbCLYrmw/M7ReQ97JQFN/nl7IjLiYkBfh1Akrfa1PSdgT0OJIe
wNfUuuw8cEj8fEH0LlROPStZhbiRT/sTZsnQ+gX1fI4+1xoxiW9D9YfCet6vFmP6
Z5SdfwJoA4YEvuwqb8+ccSwuxn1xbVedvnNnI7kaAsOBpoJ8FGucIrRU03c4iCpO
BBSdx9TA9j0hYuyW4fMboROZ7Q+IG5q1RbAIJbwwno3j7JhI0VL0Esj4Wy+6KPOH
KDPS0NZTZOpzbrbyGq5Rv0gPENAbpdQSbuXcGkTmOXf2AY+yyGkyW8a2Ts+P2ayL
O9QVRl5XG7z2tHVowjI48GaZuUOoRlPDyAPI26uXGhnRgE6RvPG9xkU5FdSO79tF
wS9AxtYzsQWkVQszGSKtAyDYnQl0Axd8IxbNISG5zwTAbZOSPpB3iLqNWUPDPxNE
Dxv7Nl7rWddy9gHFIpZ1VAxHw6EbbfGUl9dGZl7b7JLXh9xmNead+UI846xHCVif
D/TWbSxTtSnrXA6TKvBtXc0mmYYcqEWVNqFKi5WRHKGeH8y0nwBjp8IN1cNs8c1R
1Yo1B703F/n6ScqKZXeejPYu5MUqoIRiQbFxfHzLCQqlxtzuzD5NE82t92e0gh8p
cgZ+Co/YY2rMJYzUG2pBjrZY4trA7t8Fy/U20B9NnMd9+JL7BSOAaO5ff7vyfvkU
FpUutB0BxTtd7OtkWpzEPiw4qadMfls7B4AuhvFACaAwS031riFFOt4usq6X3Xop
tf8X8oSXcSmm8+uDXhYJe/3wEgtzO+/G565FCLnmZZzZupl+R9dAm8o7Tdbr02U5
4ELxpMM9wN31jP+DXdmT1yk2VRFnObG1jEl1kPhH7EDcbBYn5qcZsZHf9jO3Asjo
j4fZIP1elx6QbZ6DaMe0c8r60P1tsJ5Nxhnn6CXLtuz0ruSxXDkn4RhtvTFZ4yLf
jF0bWOFHy5VMlIWjW3FhTbZAPuEdn5tRu1BXCdgnCuDQ3Xtl1zzzWOeLEjXMy3SP
dm+Kz2m7fgFQ9s2ko2KAw//Qcfl3V4u6zjANqloJ5YVSoh6iXkJZQeLR1xP5dfi8
zu861Xm+Q0G24iAJZV+kspOjTas1qfB7UOQEo8QYcC5Q0VKeKh8vhINW9O0zwKTb
vaHEZVKDBzq0SIeJezrMsGNnYqnkguP3EHoj3Ye+Fo2PUuQS544YjIheot71TSvi
jst6q7Nt6EcCcdgKY+UiBK+N6JdYISAT+uAXoNvaJOJrITRDqoQbanIfwD+NUMtj
Y9pSZyNgsYgMLIK8WFVPM3hfxgvBEw/Z/rRJGEkHK+W/Gai/PaS9l5KsBnIDn4gF
zkJP38VvE6b8/NMRhJFatmPeHYhwULq6xQ57wKCoGScyZu2fbXPo7/4vklQS4Ss9
WW+B+89UDemgx5NYsZ4/XV+3W45ehKR2bYLpu1wocBmvrfLVYEJdepdxV2d6G2xp
cKcOj4k3bD+HcnE+0geAgZ/JFz2iyi1oTLONrxmKSQjYhe6b+UvDz4z1+0F0czrZ
ygaU1Cd2Dm0sOdW7azZcO8ug+qXM8x1XEEYnCaQ6VOl8JpZSImcFsBej4+PVQWET
PDEAqmSIvK5HD/PpvtJd7YHei9xX1/3VzmNOXsmCmtJH8pAsr2OxDa13jK9CuvTc
Qk5CocdJak936OhcTqVK0L6yodyRYcmrOyxfkdiLjQTgfQEtkxuWIuKkSsr4l9ad
XgHMVbdVX8mqHLR/DaBeQkb4hf9en4jTzObj0hg9UXWYWLu9Klg3icE/ORRtOg6E
3BGjA239Ni3jqn1791lzXuhgLQ91FKbB4+JoV3gtTPzGzi/vJMcDeRslmIaWu/vx
AcVpn31Gv0HEZlyp+8241y98EF/TeIZJ6Vo5sqKwquMCWqfux5IiV8m/mvoPEW19
NX2nrnybvAVW5eKdjqdPPpr1wydyjs+WGlJDSWLcq88stv7UVAreffp/K3NmSPz3
WBt39SIDHUiV+UqiPnjjv4P5YLjLIvz0Z561Of62n8jt7E7IB2cCqMBID5qo7J0v
7pMHwzBCHL3dCWrOhSJ777kws1dSIsKwkF9SAIFmlDQGNzdbsX6jSpHZtf1B9TBY
QZ2Z/aZY9eq2WZ0qF/Un+iJ1RxdcodWAHyEOeWskuiEU6mVeQIAu8Wkj+x0TtDGn
erfwtL5SlOao7Bf5cA79+EVJuMP2n/BaXm40CJZoH18KYd30FfTXVbEDk+UrHzRd
+noUpN/OuecEdVJO4p3nJOOQf5Sso9NQ+GyZjr2ji9IHnSNP9x9e/xdwShfpVRVw
OEAFG00XvGHTjOdcnoRtH3OXjNGa8m42XWqPNGz79h12WK9MEbAz5QmNimc5Q6Jp
XjniF9b93FbZIykjif4cq0ngMDRJ5kBF2/42gbpQc7ZmnnpgI9qjZpdIQk8+RFiD
uEbrNy9b8V3Hv0PHz7rarbNzUIS+eughwHm5BCe77mGtzx1+7jsPiXM+jxcZLlnC
kJJycBx+POw+Z0zrQm/8dJmgnrkcG3DidkluQgWCB58e5bog5KmRpzIkmmmuDZ8+
znejq3DIF0XOL0CVIujmgJNGs2qE2oM1KakJMFaZYfBgAGNFd6sg+Tm8ohqSP6MQ
iE7FQ9Bo2d2pFeovaS4S70m/lRSkYQWje9j6iq3tD7m73ep5O+cxirv4qdhubiEq
rfOGYcLoCWtPkpMX9uYMcu+4ZrDw360AqXrv2yPXvG6WSPH1NP5dTSckNWFLlLJE
RzP0B/IhKbWcKYqGcpEgMi1821pjOeq0gKdnpbBHwwkFIx7fhNJ5dwaoon5pJ+fO
oq0AtuHjedYLO6XBFtRtW8S3o+83c8Fh1gcZ3i3PKmcTE3YcSTBvPlXlFG3xHMMF
U594hSGeMNITG/4WOsu7TgBXK67n4Wq9gLOH1GqSsRG8hjj75AH251xdXHfaGhYH
G5gPvPEgQX/z5icwnTaXN1UM4cOnyDa0czKODIpkHlrPGMWzO0wYet4zJ7S7uuj9
BDcCeq2agh682XEASTfEE0d2vtQUVhfzUZ+03HAVevhe1cYMLOfZZnjAfS85EdiU
2GhSQ+C/AxyKQf+fkLF5jp+6T3WvAcDteDIBp4CwuIdsN+rYdnkW0UW6NHr0k5x9
PLvw2jUrJLriODr8u0nACdD11r/WurbYpyITAXYDDqmUPrSdou/wEcZanVTlwbdA
hBKSyVcpMxuEHSmqPfBMKIYFksNTT6uZsOlZ1k+4/3ys3K2YfBoCOKdCMU02dsGf
ek+j38HV5jP4rzjiLs3tsPdH/vCJjsHm4rdxC2Fz+svSyLz70wKrDDXHBNJPmUto
7S7nq66if2HfVfQQRyjjSHSwTyqu4fhTomb40YpqgWxZa4RtVCbIH8myPecqbefT
uS93hndvfzl/Qp+xyFlS632C9LcpPwTLiN6to4NTyjci0AgQGLEAo8x7g17HKsGT
1k+l8yq6KQV2mMWZy1hqCiKRTsmC2ygrjDcStNEWbBVnUDn+oPRmkBHtxFy8dTdV
AMu7mbvIucHCBOZWJq9KVy1ygsiXpK7MOu7KrpESrzW2Ct9T5zOIDx4i2OdwE/WQ
BPO952rdjlwsxYlhSS/uNmHrUlrcOOZUvb+gKFHp/u9zvReSfZ6NCNyVZmj9jBZd
GmTzvdumv/v7kdsoHee+CR68TAs4C5vCNOOK7m/L25ldgg86UYayzm3EuiuIW+2g
2y80IXvmEu03kpIMmaKf5C4Mz4r71BDZIqMVBYJy59A6xDa7E1xLBuroONwFmCNU
qtP1ntLI0aQtfez/S0dDXyxm27h8ncf4fWyQI5RMQkPsGGwoQ2MXX2tSZeiSMtGj
Z2fHU0c0T52l9DmUSWYdGEbIeXb7IzN/m80PwrN/SiAmsQrrdjo6yRcsxctRckPM
WqazxHPY7Xm5qgZC21IjEk/uKCnoGnxf5VpGKnb+Itn3Hm4/svWxkglqNOMN6Y8f
qPNH6y1vcwTAHbNy4KzJ0K0x9WIgJKygP4H5FLXW6/ASTSHEdkG0oJhiG25go8OM
QyKn6FojZOm6VssqRxuW5t4ZceUZJunmeFsJ7N/Sb81VI9rfyU2WxgwwT5Vr4vNw
m3ahwcPnzqjS4DjXFtamEVcPA0R4XnlUa3uB+9240fm6TaatZYmZMZF+7hfQSwzb
7spd1LgxAKmYBabu27xFW9i1GCd8dpKY+cEzWZfAf+dOc3cwvHCaH2qefTEmBfN1
yl+7VWdIgSTqYxXI3bhfexqXSeSLYu0vmTV5fLLaX/k8pUSzvsBLE5j7hDi4kNzh
8OaC5xtxqvRjXY4wdWUiGAh389LNvY4sAm/iPgTfQvE4cEo1iumRScWOTiA1hBGr
4xCJXC9Haw9sGngj8VC0RylkAPcL9feMfWyhdwP22XROpid2nMwALnaurqTptBep
WKnozwR0IvE9hf1dcO28tWIquNHsF/kavNOlh0tUGOBfY7tbxhD1vMteYEaxGsr+
P6c68O4uWtVDQpCmU/s7gG/zcSuNXMk0Lyu+fnYkj28UhLBmhSszlCaUMB3M33yo
pqlHSbB35UhoXA0jmWNbLkXGwbTaBxEQDh3GXIBKVAaIADTBik7CDQcVOMaCsyOq
o+Iev2sGLCI+vZlWwbjg8rgb+L3lIIob5BMDBrTbQa0FmohkIZu9okn7+SFEtTSn
OU54r1Z9jijr2gBlqAmeLyKs2yj9MBs+fjlHLJ6Hqv/rbVK14TfWmHMCrlZ1OuUg
qfAJbNxp5qi2teTAMUb80ssT/0kzSsLBANsurN1pkk3ZvW3aIdMdulVWkNJ9dtV8
jJ8NLKsrKK/wgcnwsWIIBBI4sjDBsO6vMGOGavc2D8tDc99vRs9R94534s8kQtnb
FgfJ0E1PyW0z1lckO+GCjzHI8nqec74nrgFRTBVlZdZBBAreaDy8FlztFEirwAji
kDqOGbIXp4Fj+mroAAzWqL9S1AUQOkIX6HP9g24OWzqUV7zORfD8C0NM+VzG2QMY
v2mYHYT9QyAY2uJb3QwJ7fDvxc7b9XBl4JeIwk7dQvOiruGiFT6v2FOZhiqwypMP
gTWfrJe/WYFUxTC+SuaN5N9G8YoOa2VviRLffiVBcFbRTy+fc5qVnnbSqtw9LBU7
F/yXKQLeWLFCwE7sXWW0Z9x88Pw9eu6Q8yyXKV/aLRsKkZpqLFn23LjDD+wW3OxV
xpuNw+JjAmGpTu6OwOBkfOoSjT34vFYT6wmFbWX+MMdNZ7O0JDzL6Vl0KO/hoaXG
/w6D4ZAiANJCtffuJmyoS8zuF0yz0kR3EAzwF003KeaACwmkfllcssZcGsqGTJMk
DOqVMu/P6EFuDdP9c4WBFrnUvATM8vc//8Ud/bZyFTp5G+5UtNVx4HZEaWdVxfQ9
TBwt4ZBNM9pVEeeBoCBjHqaH3USXtAdkHzqgUPAVYx/yxs+PCcigmvfWs8gl6Vxm
mlXRubXbimsCn7HJeZwLKSCyMaFTpwxSC2/sqeH8UvYzyoRtLLH9fSLicrp+FMA4
aEscBi3UkWYO9g6xqyV1yNIiv0A68yXCfGKxIdXpDKnMEbVi3xsIAQa3uGHw6Un4
Arx8TaAfGI6B4ngSYRT+ByMBgIj/i20sfJ2nMMOfe1GK/gIv1X6FNr5cOKJ19nHG
GTtD5LjAvZ58Phltzrjx/bPaqr+W5zq1KaKjgrpZs8YZMMV+eAbmkgUrq0xO5VWi
1lKQeZ029/2kn6B8E1b+fARXbYaEnGC5e8zrkKevfPPXxxdz3zu+3rEjQLwITFGQ
PBDfMKy2GbVx2GOoB+kq4ssmLwYCCkYBciMRImursCH0klxdlYFEIO1uQDWAW8hL
athR47nVzrdveGNg0bdPY9g/mi+0SFLiEaDvS1MCi0yuhkecb2+H0dShgfRzJiUO
j/KIu8eD5gBl/Q+W+A1GWsaRIv1qa3qxEAQFb8gtZU96FqVgN+YeCrGZfmZs1Mfl
mNCWLjc1j49tZdeX/26i4afVcYQ+ouTwzjnaKjbYwcf4AGplFSVAnRMbL41kCQt1
q8EHO2FpRbh6OEfRcu5vASYPbC5qbQ0Ah3ff/bMv1xypBFmWsLNn0VPXcsAdOhE4
UXqeJ7imQIPXaF8j9ljwyW+W5s1q6dR2cH/FsFtSXmGZkie1ovaAqvvaMwScmQR6
TwvBnTaHaTYGwliLQKwH1gJNgO9vxUmhv/iqxLwU0rv+X1YCWn0dUd7DGkk9F4Tl
huV/51aA8zHG1vhFCJ6joDk89XDtwlPXaLkR0w9L+uvuQfoSxLhRqgNfXVQxqWAD
XjlFy+rQptdN0MQXf+M9955tmr40Tjw1rv9lkh+nkDtPKfSPkE/+8uhm9AJHy0vE
TLYfoWQb3n1k5f6GY2zsLnIaA2TYJ5SYBjy1eIiFB5bKi/6Ao7jIMZTCAVAVu2xO
RLdDe5J+q5bOuET78kclRmMQbtVKhgGZE6SpFVc9y9+PTRIAUcdV3MfbE2r1akx+
nCS7Mn6wjjcQ25lyaw4wdCBcQRzBlI/idYO6lPHbE9zhkSdCUHfRHs6ZPuTO5C8p
J3t3CfQVmzsr99zNik8LtDgnO8WuM+5RhC/HMaLqktFM7G/d3uLvNa6tBosbMzqL
CkkL57aa4sVcape77hsL3VI73ta2M/cf6r3r4Hr2Ch+T/cR6sNSOKgXj3sEy9lEv
7Ahr97T1kdS2tn7xQ6ARwb63qiF9bfep4KCzhjXFToP323JwceKi8uvFyod+ZZs9
SpqXsSUeOadaWiSNreDaxhVoCWBi3vnP0d1AbzRFcZdIfcSKJslmVjBZhiHWQeL0
0KAQ8s0vZrj3xvGbDo6kS0S3suPLdI8c+mW1FhKN1cwT8+9t25jNTnSHfDx9oCqC
MqRdWXYgN361ShaVy/RTw/NNVqrfEDZoxP/BEJGPeXqiIXBE9AcpWQ99S3K45DG0
SioALLY8OfJytLXgaH8wSoQQRyclPvBBZAOuAkrtJgrWZfDAIu25TYdUeXEnYh+y
q+BLGea0vYVP+iV49ejqNhgWQYW3M1RWxroUuW5tYbK1KThHa+sMxaJbv3ykcTcw
Q+pGScOeGVZ3p0Lih8tb8y0aJ3l5cQAgimFmFcnrMx1HvTgm6mwrQUB/kNO8V9EU
r3yazqFaw277IJ/CPLn6U9VYXXoXIqs7E9Kjk/CWghJYgeCddHo8dv+DbFaVbxdd
N4bjvei6EfkjeQUna0p70Fd97lljpnOAywL+ZJRO+J3pMe/J9hV28+aKbTG3DkWE
yhGcYfs+oFe1/RONn8djNOfGDORTRVTqQ8+1yKHooDKXs+OKU9PDYfloOGNPMFpj
ThaLFxd1sqscYB11oh/o4pg4HkLRu9i1f508OmxcVDXKQKV9fKgJoAK9MXJQoTYc
iVKFzmRtpkyZEYmfQgRx/XkbWQt16DAWiGjkMr6HEEn5byoqMlBAVPW755pb9Mf1
KwDEPL9CNI7YK9D+lZcczN3iRTrkTiefmOkGT5UWVs/cejwpYshB2FUSjjjbMcpi
AZ1mXKQbOsKLR+ao2kfmpRPJtv4TTYxKimF36lUE4mmV1UQkcwogMzaRkgx/r8Mj
iaSG7Jktjf4wDYp2Bev3/I4p00dALqs4RTLxvTyxS3MOCyRMSfzkkNags6k0IGGI
xcLG4G+ZxIpMS8gEa7Wv1m16G3dTzsPY8Kdb1ud2ubbHYum/KN1vGpvsClr+bZID
LGGC7ByJyTmgdp6SHQb+q56dPZp2a45BW6xQJJ3GuGxiKR0JMhHcwmRTGkuchd/u
YncetoyvO9KJ4HxpITGq47Z6IxFAsrbEYFcBvLVz6OYlXx2WdGilkSYiklm85KUF
xmDYw/SfG2J/+ZwPrATJULfw2ZSp0HVycVaNqQw4gZ97TkOx2GekU6jW1IwIZ8kX
FqhdRI4/bLau9jeGLOlxxKozTUHkfYncKU8qifLxzwYkKXn0dBR876pm+2L90lKu
KC32zoQSHu0Kiz16xGxlHdl5p5VeKW8wr3N1bTGZUpy0NbnMwMh11A9ZBKJzHa/k
Rf0PNH+K+ilQT7/0N0lBZ1jPvJ29JWzghiKcoSiF0gr2ZXDwR3iNfkrzmFClY+WI
PKecVbpAUlOjkGireoZ+51T3XFbQjfX8mRyXoiLcje+86OmM4pItxbRE6LgpFJRn
nmCb14712nlbabGUL1mGEc9A8WvikEBHta6AB0d21/UNIlTkN0PYOSlk7W7WwvSP
HijW3KIeMsWPzD90PDwLOn3HvA0WT/I8cQOT/MRYtNX120W85I3z68xmhvfsKhwr
aG4jwpN6snzByPF55WyTzwdCCuvUL4KkaWJTr4N8LS/QLQYD8xwBMaRs6gXvyRyU
TT1flqrQDiYcfTw34Tu3jsPu1Vrxqzhmcq6H2dgpO4K8cTIMz+D2bx6DRmgGrgZE
ciRGrrGaGQquAwIzzsNSKm+CRBdLBvMQ8Kbf3fCQtxKEgxuEYl8PmqFQ3oMLuUKJ
r+gC/C3fLn2xAPDnomLCKk5M+5NvyhfokLeTrt5p3WZxPvrn2T7i4caepCOh1NKE
JnsnglP0O4qkpy06gCcdRMpeFsJBcVEjIVDsyMdJfw4k6a77zr3dCR3+UzDYdh6/
Ec1m6ff2bHBIHwmx53V1+7binVMQj4ajiwq4GgwbPMxaAV6pUyRhPM2+beOXDAdQ
ffNcbYMgi9urDgHZjlZCmH3fB9+gAPsRkrimxhZSV72yGuadSCsC8Zufik2cNGk4
5fjPmVqFRbGiDCYUobZel7fVjppdNvQLPWai5sEYwnAtzwPJOJrv/BaHic7Fu0S7
kqNGv1Z7ibsMgfI3eTYvC1YU7bzq3igg+hsouS6v2FvWNweBu8ICcv2dAvt9DEsD
PcmXjQEw6c+FhEPRZDfauLqKkXyg8LRcZoILVaSh+Onr/aTgafnEag3kaRSfCcFk
cHkWOGumEkX3tCBQemEgzFrkR1xQq3ehf0mi10Fjj4evjkSSYTVSA4cmNJAXXu9U
ZVGqZyB8staoVK6yskZfnjCDVlzCaRm9CdSddmLSdsMrmm+ozVDRIxPpfi+02rfW
pvMMa5Jf2kOHydUNlx9Uxrsjfz6VVtkx4wZzOoBYih1sZGvKX6xZ/P25hRtamQB6
UZZDPeHJy0Utfd3+dFcrBW9RKMef5GFPWxj40K9pB3QDT7GNgRea2Db3fWiCFm/a
8/Cme8jo7lSqp5J6QPrPmo713YUU6rpLdtMFO/6WV/mkzrwM0Ag94eRRWVB7kU05
75/7XJtu0ONcy7iED7GjCw3/Rbtu3OSBhvM8K/loOra8a1Haq6sMCCkr999OJI97
s0zsADITzQPHZ0lIZjmaB4++nlrMtaUgI7B9SNwLN7xyXnH8DW9XlBHGJTMI5EFZ
6LImRzPolRRGeqNiSVXT5Mg6chkWc6h8x2dgPrmjUaOFiImwYuTjQ0JC9s54irYd
by4bQHHXh3dcUlvkP8rcZdudCGGj6o4UEaRX0FRv6B/AWnrWuEYwS7Ud3QKt46Th
wpPStBkWwfTQYsUEfJIeCWOIVZTF3KqW3KBzTPBkoDak/ICH4UJtO5dkA7WRilVp
CIM1vUAgFKt3nEKk8ObJ092qUcNcP3AT6C9Hxj+hbjCzX/6PvkxtiYQhp2RL+rEL
MkrKWLIBIibPAb82mHzR1DFYfuM1Rc/ENH1VggLG/1gTwpfWwMCPCualI/xchaAI
CuCmlP1OMZnB/suh/TjzeI+kHOaTshQOz4by65ZLoTsuzgCD4id2hLAZepb+xkjd
gBw/hupT7dZ+JVDBmrrz8S6kTojDWuaFYfSC/F9REW01kxwN/f8fxzXyA8RpmZnu
sey11biN2Nof0ntYqPULgquzx1cUYudERQru4GLCFfz1Y26LxV69ZMJE5npGmkHZ
VZOjbNwB9cpRxf7ji/tEAtOkf2tGRxjIPvBD109qHQmPaVLIqipBfZLkT+VbUt+n
+CUkVrCxDUCQ2IxoFTXUmXLqTX/UR850YUauHzRAUQ1BBpiA04n+vomftWCvPeu6
RfcefZBUYk6EdQzXZF3Q+Y1IKFh69+0JQjZzNECW2Sn8qZKn0V+5V0/Io8/bNf6S
u6+Fa3DruZ0iJ99Jhe/Deuz55PN4rKTpabJd5iVLYZ2LKYhFF/Cho0yz/LVAZ0Ey
h7qhqGwbz5Uq/2pMTdpC+ibq+CSXX0XeIKlxTrINf/AsRbxIxtNeGrvTIreLsHxg
22nCXKPkMg4+JAfUHc3SuPETgq6D3enVr4T9X45C8FXlvAdRsATOq8NrvY+hhAhE
xs+XdsVNXthv+bi2Ruqef0RozL6TlSqDhxIhQLfJGYjRLHYkr4H/imSg2RWmluUg
MvaDUf039VLSmWlVeEsBBSpxkDGznj9C9/r7yDeamFlJoMwQRFBewIzCSputPATo
Dc19UPrZ88OHtIuF26jEeXq5hvYittPGy/WgMaqSBarymxoIKR8twChWiUGpvZtw
UUzqUWd6dyQFb0U4+26bz43jFFBjUd35JxdxryixYNxBKFEXi2u0Fo1PW8XLoG/b
rA063kDIFEhkgKyTcr+H4XooEO2HkEZDjJqVlIogHyBo/GBlzAnq9spUyg87MYVR
Z5eJCKBhjub2POixknONhi0Kxwy0ntQO5wQNvJMLiqzxNd64JD1pZKJSjqYpJI29
O6N1qncanwDCQeLvBmcsK8vOtUz1j6Tt8T3h/No6VKi79Y/Yd72TgGwod+yqE292
XGH4zeSrzJH3brQzWiz8+ODY86v7CwH3Zzt0iY5lYEDPvZJ/j282FJ5Rs/ZM9+f8
R9qgXodMkYTcGMaiN6JpKYsx/W+Lms0Qo3coVWHO585ars18K1wUTE9bEpw+LVpV
y/57svLxks4LYxuj0Pbavpbw36geZhMCzUsiercFyCnqu0ML6pi3w3hA1OOAkypz
C7fz1B2f7g31UgzvrBmSvg94UrP65NRfgoiQJH3jISJqY3F3r+cDJyomAzL+JToW
/3gd4oJMPqnpGz3yuQTGNDpiIQUDeaWs5yhe6xToHnm/v1Xtv9AmnRvF7xMlTsmA
lGYsclveCFeqyuDmT1RsZ75ji9nqcrofFWQ4z+EWtXT6uKqouAt0AEtQoYDmIw/s
j6Q01q95oX+wErhm8+FritfihUsZuy+KMSpCdBXeki9BiZT/G7MyYrC5NPvmpvGb
JJ3GMUywNTzTGpij9i92gZJMyAFTBn5ELGXDEkPefHGT/oklhLqMOXIOahRfLMdr
ERIyB/cVoPPfjyniQyUSiJB7p8JeHAnBDsPM27MWa8RRGwuWXq5gu9o5p3ya2c2h
X9cLnnBfAPrOwLSZGrMK5T8Pi4rwGemxpuvOsdMDxFfa7EmaqouMyJAO0Dfqx51R
4laSC5xrFVO5xXmOwYcn+h0a01UUdqROH0Lm2rz/gVIwvxQHWN0KXFU8H/+JmjUl
aKS06cwl47Y1nRRLwQd6/RDNtMWo6oo49TwKkBC2BBHzbjFCdZVXtSFBZ9Yg/ZlN
5ds32pvFF61Olmc0gfhUvbTl56K74uDEWAT1x+7zMZGgwdTUPm0o2HNdGL4sHAlA
ByWMJ+2zcWp2Mso/H1Dkd/FdxDvJqlDWheUd4IR7vev3CaIWFJKyu7ZObMq+bs5F
xcoLJPVrhvBQu1h29lQENiATJwf6EtTCVilA+koJwjt862tIyqBTwt2P/saySnY7
9l2kIqrNs77oZF5qKM3QlFX4Y7PHXHIuXFheE3W2qXjcGxK92vUjWcz3dobuEO4Y
9x+IIHWAKP8pEYmmd3lnNUmgC+5PzNXH5vTBuydiwRL58uuU+6XwHHx49T1dlxg1
Kdi64E/rVLEpVdVYkn6yHH9nNhdfT9d7D/4TUJKaRB4VApkSnKEx5qsxKfPr5ROK
vkT7nKEQrYTnv7dRiCM8m62CEljVqkg8j1xyBKPEcyFtKpR047Mj9Ii9WYai/TBX
WlDtRGgrZcmjZJFrDZkvZaFzlIv9bwvixYfvuiKFR8QI9sG1GIWkN4M9MuPOgNPR
mgfv3HbvfcMIJE9xxM0Mm/4eIv+Ne9RBJThbWXmgu3UtRqgSou7+LoBucKusy6Xu
tLNpOTs5+aTrhdNF93Wci7632XSu3V45Tv+Xx1vJo6deNVzggGta/+MsZ3sagLzC
6G6L3c5y49ExV6t+P0X8FmJRbchObXdyoNOiZwvUSbuCwgiAM26K2D7Grc/dIjUZ
n6KSys6Bi9NkEieMwMbaRThu7UgXvywWbUBWyUGoAx3VoeXwWQ0GINT4TTMCcWvR
yiBcI1p+4Xuh8PcScZtTCnvsPJ8q6898srs/HODzqp348iQiUHdLjuZQXkFtIYzY
Rk3jdjsTrfJ2ItWyxVtwha5RKgHaLjp/gYZaSlJkr7EresJJyRbWuEosRXMturpE
z/W5RBTQAVbj/6bgRBuKyQZCIJgmdLopYZlJofQaBbzfzYa8Zm9pDqsJWltkINFy
L8CUTdo4FgDtH5AeZPJaFk6inTcwb+n9Q1Tyx/xm7Ma6DImFz0R2LOsG00P/VO8q
s5LjaXII2zedvfJOnhHse67ATFLbUjrNlvcj4v/kLfPrAXYmctEQ/SNxjndEgQ7g
Rcnz+f2PJO/zJ25qSn7IJnCpe0KoP7DruiPrqxmkoLXJsusKqCoY/SUwIFnpQ8hr
KJEhYD1BwTPc71exGkM/BxIaNOjTXZhUjO80GxHFXljWXH63JnMBRVCZYE0OtJg5
lgiiKvzOqHs9Rftrsts2Qh9zaGos1x229NdP5cOTaljrXFkG+MkplSCR3bS+tKzK
JpUOWJ9PpqumqKRyowtiFY1VqZKT5myck6VqM+vfMqZrVPQkl7HLLwXdEhFIscz9
SLC2sJaGYS6UhXtfeHImWWC4xjy+oWOhIOkHKIMO890JgY1ILTbZ/SPVlONhdeGH
79TbNHzlK+qsBMU51YxnE6fa+wcFIrQHLCedoGb/R1qCrfSXarLMll5PmTcsfjUK
a9/67YklLggzBtgefb0Jxit/mwWM281aEEfJgh7coDBREXhGJiTwo6OQcfruwL1q
3GC4wxJhog4Yv07W7TcYqwOdTwuTwoWHCkYfzFfKhzW331FsAAY4pT6maZcXU1xe
Z8VgKmSC14eR1c4xMaKivifx4hGRsKNlTLp3wOV4lwdLvx5lgKo99S9/UweQF3Ex
49rO03RbCy05qgPDVBs36/JsvQTa8D5s+s8g+UfNMBXAW4SEHS+5tiqUjBhxlIlZ
CcumeIwyc0NS5a1wqwJ9C1hKL5FiokXJaz9mMzmbMunTTEXSadjXE0MlX+iHgwe4
j95lAi945EkkpcThjiAbsvdPW1wV+I3BMSv1bnBle/70Kv2+VzwDPOImLyzmyAZd
5cLYfXiUEl2bGy04nPTeCpn1qRoAnfK1QFs5VY/BHeuVXyfcXb5pTlGJoWmwhC9O
B1mKN2GeHfWRnF2HD0nEnwVr7Ebxt5T7Q5N8rlHIL0oFm5v9Ts9C1/ttTZ5TVNt1
Fll6uZZmFmqUxFTF0M+7PbtTxbgSTc+AmWbUkJr6OqDW4rmNtPshLj53+wz3NkXT
ckKDa4+9QxAxIwYUSDrS6oFPHAtZd+3rLd0fdHFQ2RSGEWTHiWnUPCJF2zGaQOJk
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
MViLbSNfznox0ifZuXXT9O8lZ36fp09XnMsWGnctjaZRuqY5k/fq/t/VGu8eMaJ+
Zj0Xwn8Lt4DbHZpxJqTW6DID5ha1tYZmGlFaknjNhA+ShnnLFV71yuSDaMdiO5eu
1mC75P0TQ+hB67oeRX8buFztaTnuRlxvPnwb04UhzgzFODEOW0iqOgajx4KUnKGz
LnqKRdK5MPwJt+X3QomDh3k55b0My8OfruHajrtW1jmDc+nXQ6zOY3c4qmavvj+I
p4BSMhK+byQsa5HRj/3Mn2KtUVMzO+q0rvj7OBq2zUdaJ5xFGxUoZCIfSME8zh+K
KatPH/XqDw2QBxN1z69JUQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10416 )
`pragma protect data_block
zJywOcNCYCPXebFMcTeAwzIfh9xuZPXO3AFUymz9F6jm9of0Mfvv72Zlg4PSucfI
2usb+4vZv+30haqF28UfETHzdC0x5YzprNBZYTGjXrKee9Bx2SXndyjjFKv9e8jm
vBppAqtB1OkQ3ERg+J8r+YCnpyFT2xtxwDPsiBwSjBRiv3A8G+Q6iG7vSoGbfynE
S+173Q25lEHMTx7TtEup5SnHIyTtKoCi2/+r+sgyzRTlZPjutL6V1+V6+oJI7dxv
vzDdfdcek/P3aI/hNZJwH0Fhrz3vkmcJWXDF9rKN+C+PXIuqCko7R/2xwbnAam7N
GT2si9ciWUPbAxQr91yOc8sJSehH2YRQ44hHDPODWsp42FOSACeezdUHnE15jJ4N
wkrLP6cFenKrGX/wK1DTn5tpnbwGsZK87l/t5Ftv79hcLgIX0hyVkEHxJH4fLj67
Iwk0HnY2C4gnxY/iE53HGmnUcTYgG04V2mF0nF0qLehwjV5QNJ49wfFBcpPSYuHh
CvNFMxEc6OKeXJfmXfkWn7CqsfLt2z/YCpIrsx3XXh3bTmBHmO57Z/rhXSXiX4wz
i/cka/XFV7L+ZaaIDjdr/HJA4jro8kXa+C20Nhd2njHy+GJ9EGi3zHNQkmw6sw/U
j2mFzIsg5r7D6FWbXnQVLKG2UMVa1MbbSqLp1pq4tY4agJfmPnfcsrkCnd7OXgbQ
+25ksNaH2oiv3xONK/pMyMTbMAldbsC5ZziCsk4/PGQRxqQ/k3vZSwkhISnvgKw5
nus/QNr2Y74Nn2DcNtVmtZRziY75VMc3yPhJfI6Q3q5Cgtb3evabJX+alxT/5vbV
GCZy5r6VJA0oJmU5pUoeplfX4VB14ZZSs/ycOazaVRUq8AQS4OE3kAAT6lJkZ4me
0dJOAmsI0CLIRx1hrugUhYBIuDJLaYeiT1t/el2GH9tlPG2lfgX3YPjncmnXzAuH
UGqSapyGFHAX7j2VdZlz0efZPOaYl3kajxMVgUM9qBB0E0OTotBSPjYiEDEd8OxN
fK4hv65BFNXIgCreXNyetL0/2Iwe9NvGYAXYO+2M/I7JctljiF0Awdfi5tUH31ut
IvHNcllTR7ATuTN6fM1PO9EnY3tWlHwlHsH83Whwx/2VQ36tkYTjZu/GL/ne/xx1
Qg8v2jD8qcImuKTEONdTS0S2ShVbLadkXbakGZKea0S48/Oabioy/jXAJPNWvMTh
Wk35K4wZ3M5aaNJMBNarrjOxEy2Ms4gxSn+S0hDMj8rPGGnZHnWQqdXp2Bs3Yoae
yO9nnMkzXLS0kf61mxeXZeNRNLQUkXD0YQ7yfYUiyny1fuFqW5jghUgUzzOJko/V
71hM80BcSfov0lwVOkYdU5mLiPJ1cAGuRkhL+BGY3A7ngQUOSztfu/CAWiRBziqw
PX/iR9I5rCZofYYnLkVvuCRcB/0blrtylrGLYvjYFR1T8CrIoelOhMH4ieC8I0et
grogzkDOh4sVJwN57UeO2qv0ga/207eZUdSlh46V8WgR9PyKFkpcew5Fyz9lvnFL
NU5Gti9krDHIhS9vFvIKZBaiFSy9nBxgN5ky3juL9PsPC9zI37p2yF00lDLspFmy
oXsQi98odV9PRdVCZuGond9Ok55kxpvhqaMW1OQwpMPn+Te0lOoZyKWy9jPH76j1
7ElD/IQuEtwOgPbEbrK7IOP7jwQ+4N9do3K5hOCWLulQGLZA7jHppkeOtdNb2NiO
TaSYhRV01YQp1wzPRNM/5rL7sreuZqcE+gjGRvGMQR65oBtzpWrUdFgOZ6N08nSp
e8fdzpz0ohsq3KUMKDjfSzEI0tOj9Pw1LYOrjOLa5YYJNFx24wwhDRMS7HQw2iFZ
mQDzYu+WYbw7/8uD8MZMX70l8qFQbyfS2jtYnAeUf4gJSMt6ezsts3kz9CvNsCmQ
kxAlaqEc7kDFnuU9e76YiGY2YKKBtG5QIg/srsiJ8CdmyF+oniJKZzjKc8uY4Jq1
rIw9rgHdOoWhgzIh64O0/ES0mMJTgonzUAbTv3WO4HG8ARGgnuc4gHyOQMNixL8c
WOtokRXwwnQi9R/ot0ei2VxnP3hFVvS0SWlB7zvFjSGxq381hiWsf/9vyH+ujlAW
vI5ydW9oP607tJO8z7UP+IvB7ECZRufdBMSBCYPiBzXm+lh524We3WCHh45ASl0Z
8Pe+OZ/1xl9SJg4fg06h4dZMCiq50to6UsLiY9VCnRbfcI3LaS/6vtH8S6K/OfVn
MLHRg0I7qSIe7STd6cBr7iJAXwcrX7eRvTb5rt5PsLnBJVNdI4va0apvPqePgK/M
e0gEBTGYEm6KHiBTW927oH6szWdc2p+2Ivv4Vq6jXtdhBgOVEE3T/TiXnO+Gyp8j
Y9RC6rcPUqCsZc+PlSZbwvvAOq17jICHnrxbpvjZlDSak1qrmg0wdN/DRX8ixQi1
QMuguNwDPdW2ZnuomFKLFgYSdnNGWy7qXDOEH+iYeuVn3AEkO1v8wmhEmuzoO+iY
LeRWuuDJGzFUAtZAh6yc0fKT+k1Itg6gs7dINrQm7uuRA9lB1cfboddA10Fsq9rV
0xjh7UpJm+SRns40M5YDohwFWMLt76N2evaH0ltQSdyzrtmt4YU8WpcOfbeT/rPa
RMyziUHM33DXyF7ejxV/fqrHU6+JqZZROfxUogbtWkMeE6zCoJum7KN4S84YYcpf
uhf6SPDq8vtR3qEDqSlsP2aY8Frew7LMImeqPj8XPlLMQRemd8J5XE9D2hN9V5oH
S3mr+Y+qwcy7uZ17tOtNtwCNm0jx3mSeJozq/OFvc5ZdAIMlm8Up1IrhY+h+G3DH
tdMP/oFIm9H/937r2t6fmZ9jnXzdJN9vNWCp+fAH9D3Z3OXfcW7D0M8oflRY/FO3
c2stx5p29xOe4aOLrZr7LlgQwjDJ3KWs/XfnJR8hl5PLvBYn3z+p0XvLB9WrdSjA
BkXGHkBdPtUMEDPJKjZpx3q2tjj/S97vwJS2Xis2amKiDj/2JpyvtkXqy6A7fuJt
pJ+BgNWJWKLY7B9NdKUy/9DnDDiFPzpUTTClDpFwHDwL+7+R/eZSf/j7Ti8zYMR8
apI4ghun1o1vUXbojTGXfB6d8x1NB46AklxKa4jOtzKiXgHj7vtN9ONkbODnbGW+
EzHUZHhHBRH8tX8jDBzK/2Xh1haWafvwDNxTzmoc/QAyiQ06wX0sqbwM3fpOr89h
wwNQZAVRIxmpXuGuzmqm8WnhUTqJQecMy3urjw1i58AIb6rgCbI94qft35mlqUTD
A+xUNsM12hagfW+FO6S8iuRSSV0zgKF+NM+78wCOmj8oAUy6XjPTKicNS01MakAJ
Bl4Hl71N/H5dHzdYdKVISdS/M9kEkouM8p3p1YBb3CfbBYCPtw1HEDj6s6xPIcB5
oZ540MuIcqw+5RPVQwTRmiauwbBtc9ZPTCoE+0/v1PuBi2JpqXIyVcv7jCv5W7iU
lmdqyobofDdCVVWkKvPur7H5XKQ6pjgBLwZHwW+wWXfI/0n3mQBHKIfQoAzcQ1WW
wAHuU1kvfhHvyyGkMf1XFPz/xNTO/oSYwusRf/1ra7S6lTSYdYSq4o/uU0oYHesP
ksjL6UvMd3F32OaGHlSH+hv0HJi5+Flt6+KvQaIAs7doCz5p2qFJCoMsy/IYpH2p
87v5VzM/AcofR57zENP7CQ4iHHAErhK/xeN3UsRtqI2tarz4Zts+V6MuVQTUBIhs
cCiHtyWgT3DDO51iz8bnIZfk3Mr8YWykE+KJ36rykeD+8AYA3KZmP3800xYZ+jpc
8HTXw85+xR//2eiCrD8kJ4H0DPK55tN6HQpRMq1cvHCNm8bF0T1jxUqbdgTBHEvT
/uvyrT0VM/aXKlluJNQAfdZ3l5ynw6Df55gbaL+ccAKTjw6Io3bdJkjYt92x8FuM
m1eK84JBCNpRvOU6ogCKEhfNBQZqdpnto2Imh722r5M8s4+e88L4NiTJ/tbMPaKq
0sMved6BmWfNWSoAkbuk96zMcanIlIxBuHEHohLaitlANeoDoCH6Mo9/Psga15pg
qTxdxhWBsIIlHV6yiy2BHjbTTkae1I17vOy/5ursMdmd/nSv8r9tk+cyaAg1UmGf
sKKGabo+86ubklzo/9h/AGbtSjYE8OLR9ABXLmE7tAqFqQqn1jxA2y88ysHiq7WW
b9T9ixNWJQGeGBv1sQ3fHDEA1BZGymE+hzQXYsHxNRvKyT7CarupmUXot0QUpW03
NXBi/XIPvS3nFisNrmnYSQvVAXwj5YGb6FazwDNnndGBQj7sPYg/ZmZ5b52i5A0r
DRGF68AXSoYBR9wtn67LKbgj+OaEzjjVfBh6G3ZTFZz3EjtKyMk1AKEIE220XCdt
EVSp+5ktA5GHW1VHtTLLQf1AadyWFQ/xxoIqgTvj6Tz3UGD1O16QpXnem0EfXXvy
10nfyO1z0ew5IA8kt6nSKCp8HpGXHjCBAPkDdhGN4y+gKcnD6sLoQPAeiC3VJRis
nLTKDItgcZ4AwUHBKLgr6zdFtJDUltsxN4rL5HOxozRfdW02z7DWbXVxPI/nt8UW
iUUjDORIEgrRpd5QXLT8liVZ6+xfCoZkaDHJHQvhJwj7fw9y9Oc7aKrjwjw6yzPa
eK3TrKQDgRIpmmeo0J/oz/o51vcli7G56gSoVVI4JbNRTnEAyrOIWEn0WTIFUdLP
4Cti0h1Iyio7v7iXXrDbOmBnjq0M/tChCNSzsu+RYts6qT/oS4LQAaE7ovkdUhJX
kWxlQ/UbnxCTRvlivVYdtzaWfva41VRI6cUKDm3DstoSXINkXslP070hmW6h8fQY
0pyYRUkcPUjUq0oRIrwS3EguQ3zSDuddd4II92qUapLhxl02MYYSfQxixUV3L0xw
RS0gUQTbHeIHqVApvmyBwWUGXKqw82tnf9kjGqRfHFeBTxi0tooWWBUHGwcEYcZY
94fgrZU7ty/f6f3ZBPKHFoE60p3kJ1js24EWB1aTift2X96TPZf04E/ja/x9+9yI
yK1NPLkq7UsXVkhyK0hwg6roET773m4/Sn2uRUK+Izn5HpuJQaJRGdvAUyHcnN16
2arpix03Fz8tfZDBW04GLS81rmCgm2Hc7g3vFKk4ttRBt+LBib57B8V/xXzjM3vC
960hqS7OpMAcJ1RHRpNFUgnwurC168vQ1IW0YXXOl0iFzv/a7fYoDDvFvZDoRrmR
1Zcqpm8K0VgOTnvm9+Tz6u2Cb7CQLLOHJ2iyviCKuP1ho+xmxp+m4w/os+0P5IPm
mFUfWZB2v1Afe14PPt8d4jW6f2tLEjcaQWAy5KUUUEvPKYww8uATDA3knCSscxgd
krDQaehJhlqIUkJLbQDBZde70Roe3dl9uiVU5PwtTc3ER/NaQROHaC9EFOS0PDF3
ZxrNuwPmvOmPhySYhzpUdPzFWOK84Gs1CXOkms/ZyhtyNP+uKvoCPCW1zS8wBY5J
EqH2XJNe9WtZt9+3RmY+6Gu9V7ehfHbWd+mEpP0Svud1WFYxblUqsuFcajZrEHQG
uBrh2/VpslhZZnEPkldIMjm7j7DVvpirxYznJgPnq75vXF1iBr9kYb09qQZZXDZy
eDWTuyCi0IZY9y33ySAEmUjx7lStxplefBjtjNw3MBf7QKjt+ALaQl2BYcl3INXL
KgMwExJM4aVZhcjlkjtPRnVKK9gpt7iVKShx0K4KoJTAV4n/djTwdrVnpTxjf4ua
bOvULIKcES04OfG78qMnO37He1j5eiq4UQ2ERE5rn292ExjgMMrKNM7XWrPPSBSi
PiNuHmFKpQHIzTxkJiKpOj/6RzBUM3KKHNIdm8/c3kj9nkVTCSKO8CycPyh73PL7
xdQfAYJYZfym18wdgLc4uSLZzsz+MZ53pim1qSYqENJkd66PdsnAs3sqCPuiLeaq
eNTLHY/YrEEw5kGDcX6ryl9YgZXtZW7LIGIWkWzhEX+DFvD0nUcBibv3GeIAsSnl
7QlF2Qgc1nEfMdte3TvIqbXnZgWH93DFhetqSyWN25m5Mh2cQfKjZR1wnKwkAnCX
po2QiDDBAz2vPxgkX8wyt3rOAhwB1LjG8sY4Y0SSHOes5W+7b8I+EHqhSHApyaHG
ZLH3UGMGvrEzxqRZeMAMaC/ZrKCoeumUKv72JZyBbN63Rk8b3Vy4pFBLl998qmW9
zLQLuaWsX6j3Hw5sMek2IwogwdFyABa2s+CvTTq0seNaTFvVpBEYmsYIZZ3lapp6
JNtGbIs3iPAiuRkURdplyeGx1YPKErYk/4qJG3AypP9sWuAYpKbvgwnbymZ2djdq
up4DCT7hnGR/GA8+M14E3TwhTRttbZYP3GkBXGWRVrxGcKc8YlAbYkrPz2WMtPME
p27kcDk6Ll38t33x82aSRY/QM3+F2gn/UfwF9iVUnCYVRH4OM9oQ41DLPtAA15zp
rRISAG6OuJcNo/n0k0XCzdsQllAxkczYvre3Beaq8sD6ytr7w2uuCFyzOvjRZR81
EYqVs/gsfKMQKDm7fcgGIzD+aSc/lhx+VmXOnxEW2dbYz/+EGPqyRQYKiykvibXw
7ck9DAZysNHO/Ifwr7OIQ7ukwdQEs2Ik0CyiBvnoCvUusRCyuLHcRkXuP9TPO7rM
f8bSVgNMi2dVJaRE2iZ/xoJ2n0qYwiMgnBvxyEFmXwlGU472ofybeUQBJMVKOb+z
KJWF817pW7IWmOS5l2H2tNMtvXXsKqNBdzDTcvrMS8j6Juf7IkJkTVxcKj6Qz4Ux
3mM5wtbNvZZs9UChDqYFALR30apt4etgmt11f4xPaoqkyW+1H4dH+fjNtHNGkHwI
2GRU7Ua7GxnEfOZ0rNspT+j3IoQbybkuTP4q9aPvFW1X+BsD28ZcUttkfiDmmqSX
Zfui9hETK7s5P7DqNYH3Csd4urxXraPL5VrAXJBwcF6snVnSXGO6cbgV2cno7yhz
q3uepUeAqmUU27SWo1IVmIWhpONSmkYnBpKI9JLFRwqlbS8dHstGQzsbRJA+Jos5
71EYGsUEWEisSccRCgdETrAC6W347OxAma8nHOszt/wiOuT4PgBU8bsc25rVxvZ1
ky5vzGw9uJk2xRgifguZOLt/U+9jgRBgUnN4RC4qtPoGYYry5kYhULd1oyjJlO4f
ewGiRU0Ekl6SX+Adcm5GQ6XDTt6yg5Il1LUES+NC1rNAUgWJQv2Q/eaVDmo+Y0Kk
rOf88WXkywx3JWGk3geaRB7aqbzYHLTVlUNQpWpHN44XnPL1P3Z7l+qSVQfrW2El
TBswhlavdW+W+YZTpA4AjyX9OPbevZzzf0mOy7MnJGfhhdTmY5AEXGD7FKE9jauE
IF2bTwmEI47PueIS8i5EzB+lbBpoK2OEdZ3w0uLOQH49jQgm2ZnX6w2G/5vr0wqA
edWtXNk8h+onzadVzHP7UXl8xpiW/7LsrHjYlEHwFdDzN5PwlxfsxlmW62MXaqXK
q4k2PNIgWLkKV57l75dWa52TloKJou2Kh707CfhkBKqQFMTta0TSIA2JlQ7dh/ut
nJNJn+H4+dqyZb8fzOKGrz4EkNZIUB8TOrrNYPtWeGh3EwbzF26uOH6e+2dknd0n
qc/cNZI058I/B8I7DPgYvqycRylbfp9EemO6Kw/lxnrNMWKFv0p3jNjEke7dT2f0
Rpw84dKZOO8If/JptuIN9Ypa6ytKbM+tL6K5G4TvC7Bogstk9PGCBUN0OiZT3ABb
A7184X/f5wDwAVjnrledSsfvTUulGb5dI+pz21Dr4l+WXVKqCnZy4z4sYI+enlRL
lUdWq2MzuJ1zpIGKbjLUyxd+MaLNJ80ZqE35DOh0iyHo5T+p66RXBpUcPkTz3rMF
iXGAuRAYHwf3tA1E7QTDyK5pPx+bArjtgHAQ8EU8ywRJ5KMjP5Kc7+z6vmNQwWNK
hAXoh1earep3pZESuoyO2SFXpamsk1m9V5sl24CClnGc+M1MSR4fpn2AIcS1OeZr
0w8v6Ce/59N+FCauDTBcUofF256rGmRQCz0CwkyfeFjlywEVqFZfpAlZDHTQfMOJ
4itUTErCVMGGzqQXBsptcnc2e4If32BsEuy6TVjfOGAUmsz+O8rH8W2ZAXxmh8+M
2Aa7jH1Ycnd+wa5nXn0D7IVKp5amxNu2BWiXtBKpuRHRNICl2L83qPsCjhaPsQsn
8UM5VogJsJAfBdhUE3yI7rYxoDX0apzCGAUn6cFGBbFQENiLFVq9EqVLrVt+ZRt+
2Ye8QOb4Y4JX5N5KSCC2LKT7PvWExu4CSGY1LU/9LLUSXEU993lratPx5SSdQtCV
UTjAtZFvy3zUSvYw7ifS8A1YzAuWVB/r4M3hwAXk+kraXRqSU/aVnflFZVTZUMIp
Pk1m4HhSXKtIZDRCvRUAlNssfx+r+ukGD+/sdcdl9VmT6f9RCNz3wRlYl5V5mfsq
HQSLs7sQLV84TsIGw3k1FBXCO6O4BQAysXCASnaZCjPjRBqQjpcwHa9w1aUHQnhx
o6KCzF/ih2ZAZgJ07o9s7hKYw+obJ6RNFzbyKoPadar+CAshpi9oNw125Jv0fIFi
yVqBLHUB3LOdlbUQlXpx0XgodQnQE2wfC97O7i5go4EVAaOka9Ux/leRdDf4WAVg
u/n5vYVxyVUeLWdNB5hDoIzVVPm7n06OAiJ7EDevj/YaTnQ4C8sGjyXwXQSaGbBn
Ncn0vZvXGi8ZQbFip9eVnWzvEXB4nFwsHqB7yC7RRIFgIzQXPsTUtyaslJshwj/n
wWRjiojeqrZPCRFWf3U2frOXp0qvQe628MpeqL2KfogVTNozGH9BE45wPgCdagAb
DHitWslz++mfaSWiLaMyamUHoTy9zEwB8zLDfkRZ/UkaKoS7MpRRHcJcS1u5LJpO
nLXV1AMQkeM/BL1Y12OR5Cc6Mfyl9guyyBxkQnuo2/6XbW6+g0Yk5yAisv4ncRWM
xTPHXyXCtC/tSwmYvWnCMZZ5tIjesx4PVdkmiYiSyyZz1FChibIhXmV4LXuKdaBf
6RsKDRTyRCTr6Uax19bnumO+xC3cd06mC8DpcB8N7ECV59Vkl4s+uLli8dJKhZyQ
eOkz+Ky0+pKpBl1zKmbdaIJw7NyGlrlvL0FxQXkPvrribGMjkkMPLWGwB6RvWZLg
BHQcP/Dq06cGrX3JjB6FbgQcUEWeBJggn/r8XLtgRpVYJaGcUxnaKUwkNY4PJeOv
OlvtSSPKpdX14ggVrz4rKLPLkm1Ut+wWf6FILeC+yLl2A4CjG01mN1fdEhYnQnyr
aq0GIkM6Q4LPww/OSnYorkHccIFBXTFsxnK9O1o8sy2fx+p2fW0JzgJTK6/OdNIZ
VlpPD5kxzjkG+oJA7T+U0PzoUumy4LYjApxaY0M0ZsQ2WRQr4krfrlwfZFjS4gf8
l5Ql4KdBFUZJs8llsCnKvf89jg89V2XXkJD3/kZrSz+BEEt1I/71DGWfL/cGMyvT
QQwZ8T5RoB9zGELLofGddG6UNzpjNaECuOxoUtfoTpXCdLwuYfGF3Uay63PA5CFD
P4YW1Y6sg077QJgRV7wNBL0Nd/trGjA52h+Af1bnE+SpDrp6GnU4ccoeNQ2TFz6R
y17qwjZRmKCkjgVbUYMGNV5Ja44ZLpNwTEujocP6QUsODgSqvTHVP1OxAyt8zPGw
dzmNL1UmcWgL2uSONZFIyNgMO4dDZiEtDjkjbHHwBQBIyDGK0bpexGUdxinR4w5H
CxVRDoaZUfPY3LgDB7B5bmFzex4me0/Pod434QZCkNG1RnDws+SbunZI1L36UG0y
P69FDIBbkhSFILd7Em7EtyTFXUWSukH62j3gN9o4x+Qmh61Ua4fobEyDJhMJmXH1
a2YMTOAXFlg1PFpBIXNEQp4EgZwF3KCuYszj48nWmVvK9ajzGUqfBFu9KYO/xOtd
djaM4YwxGKDc+/D/sPJqvxgDRV220Sr0rVb+iBbK7vyq6sFWXGB9zx7td7tRphPR
SWLTU1TQGa2BuVSsZbiZW/55DJxSIUYwZYlYg3nGCG6D3M5Abkh6CRkRbwZRQDdb
iUOJKghjniaLnFwSiqSU+w/hLm9AftfdjKYSr23Tt2dM36nxem2NheW6pIGa8L16
v4QWZfrOhrsO7lmf2rEAOSjSk/q9xdbiyCtjscSfP/BjqU2RahHEsjHSEVYMusfK
O/2dZ7kunhURMAD5D0ypBe+c7kS4Vh17s4m/Ah/SN8w3mYk1KsHhrS1K7UjHjUXb
wkM9p8PTNDdQxORy9j9vEqrMwHjXvlbRMmLcN3dZd5nipTRjgcFsrwywaTSW+p8B
THydActuCpyBskGnSgUbQY8fvPYGUJmJfb8fHezRvS+tC6x0QuGNUFPw6hg2u769
enWanbV3rrTsZcUmnAoMCpbvRTCd0/B27fvy1Y3+/WndzBnWV81qaOMx58plvdTG
A3x5u7MQ1sKyIw/usFUCx1kKVvwsOuOQWse6+lWd/BRMo0wtuxobepQU0K41YRz0
wjQtDrPbtMS82JtqFK1vn5UQjZNWsrvA9GCuCDUbA3dFBZ7RFP8YSDYTjl0w+l4y
1ni/LmviG2YgsV/Vm7XikdYt5+N+MaFex4iP+Tfs/bnzuIETYYIm/0T0IDkSbcHb
omg6uZlQs9ehQPP0DmJTjnmCL2Lnn+7sZxmM8Q7+9rfl9cdV0RefYlBRziWo2p+0
kw2XG1CBta7yQMkMnmPb2LvRauH9bIR8CHHFyQ98CXgvANM2dCZSiuiJEtsZ4ru1
axt8em94JJn38mgDIcNDAvPZmRhs4TtLeL20C+dtpJtcXXk30fkzuVdAIhnUQJfQ
+zuRRLHeVF+lJBt3HKJtb3nCqVxU72mbGCDwVFMKiuqV9WIZcbGp9UuyuWdAdwJ/
PF3Zs0ci42LWetHBoDmi+A2PeXhDZ0f9RDhAWXXA+jSSW+9+mKo/oi8eMX//zYTW
zbaw0GnFM0AgPufJmyOoA/sXxHmIJzpYylTq8wNrHmNGgwqJr8cotv/Eoo+VJU73
UqDhOolBgXQEXOYFtnRXatQHMcSBzrzYYO30gYdnqmNrlHxu3I1vyBt4ZiZnl9UO
XAiv1F99oin0Nh9BFw+SvOAWWMwuxN1PJJHS9vfKT4d7DyX5QUytOPWx10MXbInx
UGP6pzs/YvLU2eofT5xR8zC4HLyLOrC6bKWNWp5GYY2aSK6rpU27zBwcRePOap54
ON2hQK8nMcThW34iwQ3p30ymeu8wrsV6Fqb0/dqaT0rE/7Hf/yf+2A2GVDJLJjhs
V8PLB6tGN2z3eXUorszDAS3Pn8hhyEkYJbbEpN1wv0se3A6/3SEEadQnPtuBsVCY
GzJJhZOHIV15GMJELApTh9rWs9eDDEf1xiBhKmp50moX/rmCy3fj7uaOYbmRifeG
CCoZ2v5UZyyiwO/YMDh1kWqYAPySuM7cRZ/Vz3gUZK/B+OcaIB6OXG5FKXiSM4UT
CpTPABH2GclARGug/6RQho73iPdJvCFvHQpYDFFmOVK3p3mVWV9fiP5eKH3Wudqx
TMRCQbTPi/HigL1k8Jzz19kmHl7O22ktk773rDUuB1JPQ7Baot+GRhIyCMp+0vhH
zv1rGcWXb8OJoKauKrLMddjOOtz0aScYVgKTxKwdbEpAJ29q5wi0DnkUBoVcGDMV
JvfaxtbKZ95MHO70xbsESei5PpFoGgFeD9plOBLLgmtgtHYKsxQChc5SnBhcNlhQ
+c+jZoKrZROkZdYSBBuLHfipwMzR9IQA4PmYw9QdL/B7IC+k5XyMhOBBDDt2Bl0O
pCM7XmaCPE2LmEJ2+qxI7909F7KDkk1FZ3S3mXBX4chahhNMVmB8zEYJ0HgC0Q6d
pQ/2809rgbWCYxTXRx6DTbakk66QEONn4DJku7ZZdCWKBACSOoVUnTiFSKQxJ4dl
XWuJPLXhdG09ga1kxOVIJzaN27TSVwAiCqXmEjtSus8sC+62ILJRSj5dXDT3sZ+7
S8Qp0NTPR5bpvCxztWm56SGf6XwjP6x+cm3hJVp8squcpBsG0/s8fvmXxU+1mR9e
48pSZ8r1QY5FddKc5PQxRiTrZRrB8VmXpKKLuUyQhi/TgQAvAHengUEeaC+OjY4Q
+HLy/C26Cs/Q1BmHx2JaccBaXhSEBE7CyJpdpsXLTJjm8iQQjocb+UUKU33pBdRm
MVNb0VFlQXnHitvLv/NtWtHvXO0rEjMuhasEuM29KT4dXnZa5FQNfUo44/VaWtsZ
x+VH0UtFxBP2mCj0r+scURyWGZWOzr2fwc1FoBm80XmR9/yOXlr8Bn4h372PZ4GD
G7ZNHDcDJIvYEOwaeeo+6arZgpRU40DZFXzxV+JdwPTm5d1Q6ts0XOIgmx31ohyX
xQRiWs7OcDO1uux9k8P+ChWmC7XFnmavvRRgsUEJdfatEl1P3qjQMFJCh5Ddg2vW
Rohbbb1vGENeZ3i9Fcj6womuZMlsaKI9hz5fSkhVjSISAOJX8Bw0TcD6PymwUIYa
fz72JbMBE289TN2jMcB2yePzLHzsXelfhpjqyO4I5pWCmD/QsXhwAA4cPfuhj0cX
TWERu/sJWJUkCifFXmx/NRjacotb4oQyD50JjD8SmgJ2YYU4g/+5Lc9JrG2fXHIR
gL7YZzNUAspgFhnwEAmna+Lwt53f3g/36tbHXaKIGDAbCQzcCauIaWeVWYr9QsLY
gLrFnSJ64PyYpRwhA87X+hUs4x19uffZtQfMFbAhPC36FTAk8Nu/nr5fP/M6VmOR
bHx0J7lVBmhIH7iYEEOHvfi4dIGLwLuuwHxt1C6P5GIYh413lqeI7fkoaXnRhODp
G9u8aN8QXKJ9R7ctY4beGj6z78oUTE4vduwqVey/weuRRo4uhnGvPyMvU0lC5LS7
Dt2rVYfCytyRqDEmiufOBCCEefuk5kW45BIW2rmKuNowLE08y1vBT+Sgw36yOVFO
tFAJlivisbDw+BRIc2t9w1XBzq7hnPys8yv59oA5eKmx6LCHr6WOSOVt1wPxD7kv
wy14gvJNn3BVxmdSAoCE0FwDfktpWPKQxfW1VUYE9BJEKi9yUcCWCuYci6Iccrg/
loOU6dsvXnGl1PMkClGgPv+Xd5DxKxe6m463QZ/W3/POoKgEksgI46AhuBnBJ5ol
/qd9flPBAUX04z0soSJMbyoV7AWmvGTVnr4V+7qIGBH/IL8L/daa7mAwKgADFjc8
g1+j7LmcbwVYAUSPYpki6FHdbZWIalTeBbJVAV4K9TvRs7MTIM50e6oKJpK3r9cN
GVKApkzw9UXoMqmQN6AYPZB+64/RF9vcwbLJo+Jgt452gEd7jkivnUkfINN0doPy
xYXs42TzePp5JVAnoEtrpfkuMbn/OneqZB8il4aVMIpAxtnikpN6ercw9JBuPMlx
A9a3IkVfUV2SzJ1mLiPtBj78KoiSbbLiFJEtZp6Cs4Cd3ugSVc+17+OR9DT0v09T
bTiYEuGGbBERSHmbKvGmfxQeSFhf+dLcYq5i3bUtJb6JnemvdhtCKd/cS9v6joRl
dr+Yo2xQ5s/9Rcx+P6/SHi8kuV1BfVGdmHWygpZlZt49i4c7vp/ebml2FegUjEv8
j5Caet4s5WovY+BgNDFFJYYOiBrSLjLxxRsjfdFQsrrqjl5OGn74DhZdNpAsChnP
1IbPmmyyRFEyXS45ocgYMLpFq30/9X4MmOSMd88ze5vF9SIjWswTFMtl4t/haquK
S4KtGuD0JkFMPuJLTkF9y6Ly+sFO8XHYr5s7hQL7QSYWByeVQEDj64wt0NAfACMi
A92aCoVSmPWXwI7+NpeUjFbg/Xclx+R+ITmRhh+u+vyFCaAwntF2ZaDu+wH7beAY
KUICuneS27z77vizkd5BA5dTVEcpDwRitI+K8XYChevA2XrsX388iN6rl0ig0YYw
GbBHm0EQ8hzhjQlN6++12EXj2pH53K1Qw98SOR/aLsoErsKHhr7u+YjvLpm1vcJk
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NX9eK/fcpJPx250CwLkrh0HgOYgUdsMsQTmSHK5884Nk5hXw7giXppSgf3xGNp4r
/SdRjRqBqkLK9ieVS7tSIjIS9kC7xgLsOT8J6V/zvR7LKm3vbht5Lp5H52Op8mGw
zaxA5+dDO2XvNvpfdlR5bOUWA+YCJOP4Ilxcb7rN3AJpspGZsVDzFP28cDlPm8QU
RHdTuDl6jSXx3ewFEWsqxnzWNvMSb0ZlXcPCybslTuLwlqUVJAfV3rtB3+elnZK7
6TYNJeaNoqEgjiV7dC7ll9jejzoEnCsPXaRMgUujdUxqMRTrIUIRCpwdzozgcZYa
ec6W4knvQSMiz96MPqZq1A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
FLfeYuICU3yLVgpEZYAG2A+ZttX7sF059WXHL+Ue1Ar+U6SAZ3kE9wVBrXH+VDeM
2Ctvza7Nt9U00dVgv+G/9Gbwy4spXM8sCCmFnmcuLLNvREeJY4u3KmQ7Xb2wip0r
BZYlJgJ0QvNf+ezdVWw/pKvKXZ6qxUDv2hk2IMJG0cYOIXHNpu2Ba3v8pmkQCHBC
kUA8EQhBbRU696lnw8kHBAFvTibyUJe2TjZWE6ENjqLk3lIScCEjKoDwsUpT8Qbu
cG32weCnlU7ptWHLi3+zMaYbeqfh0BQqMkmJD6Hy5nHXnZt494Tq/Ej8EwjVCmZx
m4sG2hT0rZKbooFBKx9phGhuIign48JOB1hqzK/N2xNL1aiI96aPY0Gtqz8KWDVb
JrcAc0x+ULGONxiMBdbX19FmjKFxLbOJnP5v04m+ZV71zcvYMjXZumKD67JLNFEh
3KAu/6Ib3CFBHQOpj+kOwLAvYCCijQAvsqTVVQ4bLCJQBosNlFXFzcY95AbSX2Tz
bXkdxYDwjI9AIV27R05hb+b6elEDyqBMG7+nc40pkpkZ3SA2Muc2h6uu4KIdekLE
aMx/i6FzNa/L3U2z7IRBI0H8a5XyviVXK6sHiVnFlP347mElJDvfuC6PVHzdsSTg
u3ceu1MyzWebypaYdwU5JWmWSU4Al62j/hlyyu93qBQbPGpfdi9Dkhr6qLn8zBt3
j8b65kSK3s9sJGFnN2DzTSNyvHN5Bo+8I6C9OYnd+6zOK3qXX33L5CFOoMKt3el/
QlKlGFdMbiiu0zMADDtqVjBvUcge1cWKa+evH/MwU+O3oN84ofxQ9/04AE2/qOL0
NRNt1zdCIk0dtzPW7KFyU4fC2xiozGV9sGR22r5CPFgECXLS/btHAePiOydXTJuJ
LiPofDpkaWy+NI8GeYZP9Yi4lGlt5aHlGzxqzO4SYqUs6T2UqDF7+Dg8BzrPhU+i
nCPJhOv+bq6cd5+WCMnDa2VXDVYGhCcNcgZsIpbJJdoE3X7XZSKzjvxfI4V2kLN3
APZ9xjIDBrfngV9sq5Gv1zevGKVVL4aZNcl9MDnGYqKoY0Fxg1FkGGmBRV+K2H2I
xw6P1oJE2aGHaFhRe5lLm/3a4SkFlVESrxzTA/tep1b6tA3WyxGcgdzWTh/0CYw6
Q91aeXNZgLBVeW/kFz+w4wpL+qvEtNejgbQfRTy7Ok2NudYCfd9RgnQCT1ib+Nt4
9WUdnfzHHZVxQRRzoPLMZ4FFkfhW/tRXGEiPgMHBArRougI2qv2O+Oo7CYd2p4je
whsxi/oLlIXFs3TJvp7lc/ezMKi1GOQrsm1GyvhVGrP691tv6wqy5hBO9Is2RQOS
XUjZ/OsoUgOJaPUxCUWgax4pdXMcfxyFpQIM9SoqAdsLvYz2aSWXS3UF9LLxENgJ
y6nxDpnRHP51ZaAg5/6zdIcwtNhjKadcAhXMDr1Dp/EUqq4+Gcs0Bg/6jUE+Or/8
+lIouwRD7cn7cb2bbEIvzQJaBMrn02Qz7Q4WaVZWuW/kgdX75FjxKcpVUfmQUxsX
qo9oe0S80cFiFlMTQX+rMhPB1ApA+7eFqo9hy8TwDz5tmMxKwJyQYtEGxQB1CenC
8SYb1DJixtn9DQN5pSbHQeHm0Rt0Y0+L1JwpB7L7c9h5//ng6SbeiPRkjSD6qGf8
XIayG5GeqJnVE/jUXrfQ6wWGx50/9ivQL8DHBELd3pZbtLsKRGUeMweaVa/XjKGD
NbdsRFJ5a5h4d01qsHdNnEHZ2IBN9ZfPabsnskL/nECl6lvkjP7Xbz7vz+1ElF/m
z7jPX7oGGcgNIk/l/nfTl1l4RgcnSzFQy2Iqh8edebqI80SYvVa2iXzP94WF0ZeH
GgsLEEZuaCXO4WcTGWhuDDQIKzQTiBsPUhtcYsjT1+5NDjXsHdU/D8qFkKFonglR
rvwnQG1mS8CbR3vL7uM6qQILHrOr8ntJmU5fioRF9iatbNyBIzsIf+byuZVcKPB+
9c8odEqLmG7H0iA+DXkEe3j/+DrOXsSenErbOpspHUExy517RHz9AqbO4HBrSWHK
HfHoMRbpvG5ermunZoEieQ4PSV1M6mAe0pumO94w69IEmi8rxeEikjmNdA8XPcyQ
YuG48HkbGrNzESKG4dsX9Q5xxB8vFnliKvYAWwOUeWnUrdYJe/9SIP3/avVlnxGY
zF/5aPHKfSaxNqPpAOF6PtCv+EdFLJaH0oNKXV/XHU/M6OyOjuRC0J6sOjgj57KA
iI/Gkp5gLMi7nR4Pm/PUHdrOkWwYh24PrRdKU/tprN8et1b9hgJ6+z2UUIpnDGdD
cc9H30lKOWq0NbHf8cBRQcrVq/e26P0vDaxgfrZvbdPUBHyuaQAvTU6/QvsKH+Ys
bSbwBnlhfa248kW2naoerAFETPuk2tLE+vdGHKojYHVo+s7s+63CU+8/YalLyBgK
U/hzhsAWUiPjGHL8uFPAlOtfBLPhnvpA8+iTug036wXsiifvWqJoLG8Ko7iodIwq
lwEpt6AFl/M5TBSGYAaH+X6q2IKPeQmvwnOvSOKyLV9kjed8QyB0mPqr8+sMTDpW
ttJ6nelNN52x+V2s3lHOjUobSkbf879w3zQDnaene0gIkEd5s9y5c01kNnQHJpT/
9DVdH3/8RH+ef16rAyt4033yhOiOYclzzMmvZeuzDJnP0ZPb3FzpSQM/NZ+PiYeH
f+6j7RVeN+21gcw9EjnEr7+oOxacJxp230mqbyJsrK8SMq/KYjw1MrQeWK0ZHp3X
VBJdt1DrgGZ4211qV4IUMx7OBui9kJJy1APhYMFxabOkHoAMYqSmEQkHkkHC1jBc
cqxE3UJPxeq2SAoWWAWxPRy7AIIxOjysXmsN1f7WTZO8km2Mde6NPr7ACTnAE0Wg
WaVw2tteLwaB5+PL/FpXifSvmfrNObwEsuKp29D6M0mmAouyUpkFbS03vVpo36vr
SwOwY8JWMrPPDPlvzgGNY7u3etTR6Xo7v0FI+pgf+INYQ1LWYtiZVo/hs0YvejFM
iT4OLNt5ia9iUvY68pvu/WgkVSJniWtgq8yhNzTZ6rHITf53dBBDYfWofv1GuBKX
RL+hoMnt7XCwLMR6g6EU48w4FVvIbP0r19IVA1Rtp5NveX4MW56lQhT0ncziHCHy
n+02Q3d6faykrF1S8kK5Ne3KTEpFfNJxMMiEDR7ZJTnNnZi93NoK7TsTGIpvy2Vy
st6suveBdN4+QfoiNy4C3Oahf0YmIFkRpDEgs9k32Sp/12BaKZ3FQHhwjKxfZtqM
A+bRJYVSJtyphT/+t7iA/8IWIQMrKO+cZINe1Deo48pR3/MfphjbncrKkQyMl2Yw
mlkXk+Rb2pMQzxMKJ/IHruCrv8NGTKlIBXYhwqeAFzfw9xGQ6YqFghoEvofaf/Ws
mxjO5x6wF1wyV+QUml7x5SIX/b6PCSDQp+agVCYTsG2vm9FxlJwZ6YJxZZiiyP82
GFkgDdF587FszrXPtEe2+L1QG95mES6Ozb4NaUmW+koK7VHrvLYBJB7kXmIfZ2aa
1ehai05gT1wcb5HLxDDkTucZzjtEA+FO4dBIyKJaEik5lWg2yzMO5JkGpkHWp/gy
89mCFtwIfMpG768tKLK9XDedUK9gYtXmHLIcnaCtRyrYEAMG3Axa9XNpP1lIu3EP
PFSUWYjCiQ3YQG1X2pJXLKCgmgjiurN/toPyJlNkxRH1oAcCRsPjdEirtYpYMoSm
LF+oDUABtsSbiuwp2EqwXN9G+QLNd4QkxSKDRFibuqh7C0D5JYDKXtcbRlhCjsu+
2gf7BLv294ARU112HpculhlK1yTj4GOJy9yntkfpfuNuPIypGSOZ5s4hb98lGRz3
NzzSmT8VeKYadAOytY56kIAzyr/TfHmK4hPHiW6fQtEmfRknKuHUejRpSzTBRH63
jgBuS02Lq1u/mwmGrzP6eAGnnQhfKCc44S5sNOtEXmOQzs96McDTNpNlBTB/4VhB
ZHyQh/vBl8Um5Orvu9YQpRxV50+49kGLgdTl5wRrJGfoxRLQWadfhb7z7hGmqXMo
M6a6fj6AptUswCpxT+FitoahaY4/qR3cHuv2unoHR+ILE9P97+cBZyOI6rI8iIzf
JWEa7kAJx865rRJUsp+LfbDAwOHrgAQPjaIYIb6iLl1lqul4+L6wEFhg1dY65M5Z
7mEm+Oq+KpyeeMbQtNqM7RRvJ/g64PUOF5XyL+J0Olnczb+DalyARV0GkrHJXdh7
aFopXLR/sJgR27pTOoJZYqQOB0rRAHm2iZPxlDOxWlzANDxRRSCylSqhUs8RG0JY
+WulQ4hVYmxmJeYp9Lrxdi5W++fklSwPh1kDP2Bdfkk0EYXHO9dnB2vX1MGX8G93
Hxc4FTlOCGBouHw9x/ru2DtRgP6GB68Px7CXE7/3qhmZoVP5sA85VwnQknCSRlN3
7n0xShC7wKoXmKiWqVTWiLPbASuh+77en0yz+V88BrCqZT2AYiX5kKsMHZhqbxo0
mUNy5o/qMcIAnTjy3kdHBk6nQ2bPfzwjjUwtKGQeQM6rb3KRCd/D6982WExLfk3S
zzV6dvNPeDMrysmDp53+v+s+Rm5/9Han+cwPnI40WxLadf+0Gb1Ou0fCnE7AIqpr
ZM0BPwfxRYi9tz1YwCpE2BOCpvnmmJ85WMh62hA4tfH8T6j2Qp6y4JF3HupI3jXi
55D/X1HztZXksx+tWOK8K6VPE4H6tDe49JYGZ8i8LDyo7vCum/jLZyaFgENcAkAa
/9wqCkaSOZTcsJjfAi7PlyE3g07ufiVZmaOnUZfGSYRZcHjg/vNWLXjIGtgW+b4d
TG3gN9lROtteg3z2hntogQDJ2ZTt3sk4sKsiY+QciNVhZHfPOwNozQ+OzyUkce5e
zEumffIobJkx2DQIwACLBESRrMUfZV/FfioLrtXLgh5IGPqLwallG1/ziOfhprKK
J0jUnZbkxbnq2oDaGEaHoNrZHSkmY4pv0jzO4/M5PV4rUxu7KWvHrwMZmZNFcmu4
daN19DDpz+w+5S4XSBfX/FhhiP3kssM2WAYktm3HeGEIdWlYF8a6s3PEg3Il5u5y
+GAPueuuohHtECnMMpQjlxEzLLi8YW9qdRWvna8ycW/Lhzc3I48Qb/lO3Jfo1P2q
A5L/WaJCRV6PAoUnxBVPFT2JJ0mF3XIW1y5JtSN3RYwYObzDolcnLaN6hzu5Y6Oa
nCMtRl3vEsdruLx2t1rauJk8ufFJCDNgHg7q6+cCiPk9pHmV+xcfUTVTe9eI2u4d
2twIs3GZWZo2dmV/A81MjVfS88axYj+d5rBYR3VSHuqOEu1fgeDkRAkeihGpW2sH
ijyD1KoXBROdHkr2khznVW35eBKEr6wf3XCH6qB29kjNhszVa6YiYbCO37pWqths
33Yn1HtxPYasWJMxMMTP8Xdu1rSRze9CPgPsSCwM71NUyBOHYzIxaHkWRSEVxP/J
33d8SHkWQPPpKmBErQMgp+beAGBiZ3m5Z1C/RT4n0merOg+/UouUfvw3CU1Glzhm
DkqpH9mNF/qUZcYa1Ze+P0ZWWWsp3p4eM1ra6IafNxAUaYpPTUaR0k738w4Ce0pn
xgcQzWuKo6KbFBl12Ggf6cymSoeo8amPvk33nY5ozp9aZ9dqZz1WZUPOXRUJEuw4
GnQ7mRLoqucU2eI5pZj3+45rh39tJ3L4Z/oweHSIDfe2eAUcClKLm8GmdMwnTqJC
qI6ZTubt63iMwCJmY9K2lH3/xBVMthiS4uOgWoLhzogfAzQoTjzVox3tByEHuqiB
5Cb5stzgzmUw927iZzaYcH1bkAve8YSYcR9whmqmnzQfoHfhphVxy7tQmSUtwGqC
Atj9pvVH107E4QuOwZPxkRjClC495Otnc970FYzaIIO6/TeOUnMvS3qtWPAm+zrQ
qLB+js5cmy2vASq9+0xQli6oM1ug9ECoGO+Ep5Wd1NcaFpeqiiTLx2ngEfdTxfux
aeoyOyn8Ft5qCWwZ58IaCZF9xK0mBxBrI9pp90xMdDELI0kriy++VNKh2N1bwh2T
SelRNhyI4m7z8SPuQNAzEHX4gV4wuIqP5Um41q6/Uwv6zt7YZBPJg93EaatP46eK
mNJBIJzv7Hc17V9tmXbj2yc+9t4EPcTBZfSA7QCcvRtf7953mpEkdjIKl8JxK5Bm
Sup330UgYR7h5q0sZj4ztkT8rSdNyty+kV61cw1gLMl2xPt/mZbJ+zOux/9wfe1F
NVSHgbXiw0MlEHHeti35IAN0uudh5nxZUmui571PH+46+O5rc+tHUeDPWEh31m0C
FF2WQnoepUQX6/HKG2EWKZkYrtPumTklOjcQhRNqe2OO2/NrbQj18WF0PW4Z7juk
IXrrw4KO3q3dg70GIq9CP7XQ/4cbAN09BY+ACsD1n0fpcSvmiHdDyZSlOu3oz4JA
CiyUMmoH51AmPugDr52xZYdqlIzdimuLShFM5a9hPpYiFqdU6WO0wxsRMOnEwtgL
xlrnmntVBmspcuO/y4aU+0OaiR2D6pYobvE/TutwDupKcv4sbMbSh/VLqeTqibRo
f5IJCAzD7PKf6pyNI7Tf+aAUguz6jKN8ZL4ZPlRnh65QF7fb70T6LIjfRTpl6kYu
eNuGe0rGpo3jfvmZiC+HQZrheTKjNesr/5eq/RqMBLT83igEUSXIpWhAkKkta7Vq
qg9hlZCFpzvs0T9dJ+7HyQxcZ0ykWBli/wzDd5cjn3XCPUlFrzpIB1Z5Eh2DfHsy
SKVrrht1gkJEUn24U0cBOixnUWkdjxbmtsTbtIwLq/Nn9BfnpSKY/mt3cMplG5Az
xIJOQCgZFMWPxM+CIKnaEER/YWGxSfZp5QzDTS50G8pJZTzaG+8YgPe6d2jvPo/M
RnrATXArrG0qxzivhxQIRJrk76yUiixi9p+SwZ453RmC9CS0tb5WBi8Zb8Gbj4So
svr3ER9DZ3tYbAgXZEQg4x9pWEkYuoXNeRXnY/6dXFh0Vm1qntSwypiRwDbWYz/d
mLTY22CrJ+44vsLOKxJNKDy9w7UeJD8zvO22Gm/pvi6iAgKxeQZuAwL0aIIvhh2O
1ueaCMSVewM8ruz4CzArbXDAKQfmf4nD4wDzS4zsCFJ3aQci7v264fp1ZY8sK3uC
nETgUpGsCFJA4Zf6Gv3xcAZI+jGiqRiC2IBzzorcV/bpp4gvmjolhP5VgPs8w6os
UenfseAvnMUw5eQtA82Qma7lKmaVZ/t/tphsd6Y30clVfwnuIVQ47hMwuzlVso76
k/xVUPv9wyN+CFkG/8x+Yojb3i/xrwy08mjuLI6GmQZRe9aF9aZhvh2zsc+kSVA7
s0C+1K1dFkaZ49MwOcQOVrrkxIFezB7hogtOIVEIwG7q2v3xJJo9CcDdBSqsko3c
lFUN4KrHGJ6v7d8Dk9PnqkFHqRJQP/l+dbGU7+W70n/4GuwS/+4fecMwmvjtGt+D
A10nnVrWbqVYkjuCIs7mQlJDHRcwT6F/zLu+aVJblZVNHt11DPBe9sdJosoBh/ih
I+RKBNaOuzea5DQnsv/qqd3rOM3lH+VwSqQ4MrbiscB962vjqvB55y53VnrYITQ0
VQYhT1RSLIeTkX5ChKywDYP/BuDIP2OGc6sPkiEmjY3JpqBIh4/4b/opgakjF7hq
aIj/myh0lSXTNa1PWCNMkFiP0dIOjvGpHZlJvbgnFKsMaRn6xCm3h5yWeH4+vr0y
cGQEY6V9z60kE9otabTAzi+rqNG3jepFjZ6V5O6V3GvdWv+36BHZTc5bOuAss4qv
YIRZcXy8zAZ5kH45ygDuDXzBGKCAabW3LrGoAtXiJ5S0bEZMmyk2ja6U5Cacn+0h
r+HF1Y2mFnPawG8RZGCA92XerN1ZDNN425DD59JWdrd60xeFcJYGNa//P+w83KVf
6xVEAJ/lfCF5a88K5GkdocYIoK5l0WEFze2uRP0umR2waDiut2j7puQFlYjG2hLN
aGmzvuSBYNgwE8ylsSz8rNLYYTPhbeVTiFQyyOFLlM5CGZEQ2YZTLL+TAZpEJcML
Tm0lc5jvraHhpWo/czjRcg==
`pragma protect end_protected

//pragma protect end
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
d7vWpuGYn9oM9nvFNwSL/Nvn2eFEL0AUMjgpeI+NrTYrFc8Vx7vMxaODnr6OBqmv
/2JDyBxgZZ+VoBSnn+0rZySq1eGC9vwnfYvGsbc5SmQOTEscR2VkzeznL9PC2fzW
QugX5HrpAzvl/2Dt0d4A45nBg6L2ULxS1XCAi7uyEpFKSj+qkYXAYy0yKZBKDQMQ
YnFGr+HAyCjj0hnCTVtHVOThqnFTbZ6NMSItXhj5YdG8sV+5yEwM83vGuNyUCXKE
fJKJVKEAS5kZwMaZ5Rh9Tw9GN38C7eEQ/Clk2H3AW7Ost/fGtMv1GFz/W2ZSsMdO
RpZtk7FQInKN88xWDlDITg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14480 )
`pragma protect data_block
q7NJGEBukQJnuPTznIZt8ZazhcVcfKd45PZDWfVQezVuoPA72Z6JY7Ps2g7X1l8d
Ah11TnslNV+xdKdWmi4KOSbZmCtx8dV6u4U9S30CpRd1RwZ+MOiTHqIihlSrVpEj
8BsxphLp45m5HtD4gstUDAQipzP1dZ7+bvkZmMICPSSL+lLKXXPQh6jH2TlDUopi
KfZZo9aVELNIAXoq9BhVej0WYIyq4xeS7yfbw1512kbAjvhidJtzlq47rJgq/Fgb
6Pim1AUvIC2teGrVupfY/M259iPB7Tp7I1upebCRq/pVyTN6mfaXfd4S555w/JlZ
oOVHqFEVSvs9xPnV6l5bw+CgrO2UuaaC6QkSOnwoydZ+Tmy9EKXw5bmyMEWzXefY
TK2KqJB4F1LHmKpqevN7qf5kwTbhWPoG9HgsPyA/RyDi9C5ERuz+VsFFirOZJIsn
KO0a5/QkdR+jHDvj6hXgNMS+hFfIiE1++YKDK3K11ZiDz8IH9ufzte6Offa2sEym
44DVQHbmp/miUACXTKy5FL0ph1F5F394cOQouTcbWIOVxQnyHHUhWj8HEVl7T7Je
olisszEOCkMHc7LdQAssQuf8E0BLpotQ5OkPUgeOntMWNI43T0aFSr5tzfV1piSa
xw54WiKBgwhkI0v72VboNNiyxJrCwkIxTFCBjicf36NTY21v/QVveCvHGrzo941x
sO+Yzo287AfDZdEC5lICX/NE6jdGhsKoOI2NtePKGaS6N2EAionxhyyZvtvmXdtJ
yjhVGeJzVkfGnOGZzofd81dlhPLFJ8/0C88V4NfDh2iH72hVEwP6cxhMpj58PK7H
IyI42fhkxWqYh4WWqRU7dKTgl+DrJtAM1bhunxz7f/CIfR6qnZM9gzqACyE6NV4A
kerCo9w2k4RjsNmo3kWnNSwQ/zlT5yqRhbdFBXjdB8kA2KUlkHP7b9jSYwkX/8yS
vAgC64pCYrqMIjRAnSI4rAAeWJNdOtP2hrP+ngvB8dSDD075ekkpZbScAYbuEstv
54Fn/Jcz7V9fESHDsJVQiPmdm9qLmM3Iz1ZdUQrPWd/y0LgSgL3HMPKYWqRLejFt
3evmq4znM3yeuqOtyvpw9zJjL0BajsrhHalPUn3PlgShVpX5KVeHOSm+v1J112oA
L0orjOf2GbN7hBnHKL086RTikdEq+Kxh3xzyB2f+EtlzrApR8TgXctvKdqyw+WC3
uPgJ4NnJf97pTg1S3/QUvuMAWO4rneIG7ecFVHBfabby1h6aksPJCD+OwhzrQLC1
uP7A7tKP4c9is5OscC8z+stkFrtNUkaGhQjzveLrbZfOs/P68nYr6uL5kcOjUSQB
gP3NIsH9wx48lP5D272ox0NT+Oq8DHBYh7YUh5/7u826BwUfdwmSpCvRoz+mhkXt
J/jCJfIt4HWzMa6zvJ9UF4PrqdJf6qOCJIbmb5L7J7aSNgv3cPRYs+34B7aBGY63
o1gM7mJmdTU0Om9RHvlopZRh/2J+FEI92Bl4315rWnSnO+N2UfteKCM16bx0/gaM
1emfouQ8aEu13dnoZ53zC1z7fLRBN90CaPOcVIkfyyIJ02gCQ7o++JOcST8pUuhN
xgu01UHrWfpNMB+rRtneKtXFjZqqEmiRoM/ZFfrxQFe4PUWyQgXi+Rod1q1IJN60
ko4m8arkXU1JsG6vHpOJvwWOs/x/YyCcOCVojxIgA5X/6m34nPe+po58vxeWQ+0e
vrMBD0qSxRuHMC3tfBmOnb9URYrrYTz+1K8zHa0n9nty9vDwS6QVegovckf96uo9
uSvgzuQ4qTAh9jIU616imS8d+aWXLNHilau7JcflXToREfyAHVU5iYKSbMDc99gW
iD+C/pQ1W1XW6p/mNDhbRxv0RChZdQ0vWjUn0/NEaE1U7cl8EJtbn0mq/qGvbGlo
HCvclGzigUpAmHnieu+vzxLYa5PpTKnZf++6XOM6QQZLal3Ww7lDW1R53IEcGlme
IFADoAq0qMPiwjPNZZZvGRhzLcIsM0g/IMWSglKz0DfAkM0EGuq4gapNyJA/VpUc
Zu8BmAInOXuoLGrUfoo5Pi3QHX63CkyqPiAH9frt4JpoNqoD983kemAggOEUT7cw
vfXIKU2GD5mw07Evmn6y3drsOd36IC377mDK8WDaCs1qZftcgaolcCCOfF8UvS0X
drw5dCFRjR3PDlQ5bPJY5k8YRm85fzVHHdO8vc9TS/M6zPtC3oeEgAffZC0SViTj
D7XDDwfmipuT3BZ/mOoUZGXDSMasreutdJHhi2N1fczEKoFKxPrnhJpVRN8+Cqwn
zX9wrqrn2ndStG8WE9qkydBdgnD1atIGie474nhb4nvIcPdqzL7TSbmn6VZn5k2f
UMJepqwAsbSpEahb47w0XqQ2CvuxHagwJzDqXvnWZWUbmechZXT3v/2dEpwO6jni
evab1waPATWyER9Yn10bqIrcH0VQgtr0VYQFaVgm0roAymz7QZWHXym7pPNj7QvV
xo4EZAEJP414fSqidZYgCPHTfzJELIUHgYhbdEPuxHUB/YvFDsQScpqVim+hQZjm
c2Vvslox2lcEDtw6Uq5GbduTsurY6+LYKOIp+Z9Oy/FIY6Yb016meTU0BUuqgTPW
Hn2U081Qbi7ZUNXuTREDbMa1aeQ3oxobBnRr0aOniqhMA9rxPk+95OlwxZYouMAY
WOd9nak1OU1YnHvGjm3mKbuO4qMypkXZmElbvn18647T7LwgaG8PJdjMkJ9AfWDv
Rest1uVkmnI63vBmeYYXKxBujcuHLt1KE97ra+eWRlFNru5x0dTldC3p0if7OQ3B
AzUiNOyKyQaoJljcuYq30tP3VZHs5YFlKLdb3CFb6rQ1G9Zn0a8MN/J6x4oNbMSw
5ZcRyZEitxpaLwOMIMuD92VggeU5ol4n6aJZZGZwDsrfYiV1MfHnd2audEyzrUb9
o9mdsXI0e/f7nk/GYHexPwydT4iVubKsjxrD7UNhNz8KojKz4LVUrxrT+zvI0oMS
MZ1Po9Gy3WkZiivxIGyxbTY6NvhBUkhgWd/ecTsuOp+VdmMmvYd+klhSNkdL4tQb
iKQ2M4dV1jorynTib1KpSe9lYtk/LYjrgLG3fstOo3SeILtCr6ruQvlTTR3WBmrY
IAGe98SfG3LztQkB9JciiiVDMD8jtLYgzudz9nToVqyPq5eSdFkN6x0HXypQLCjw
R+oCxN5AU1ISEeYeBhMn5eaqXSAG5Mp5DFXo/922u2ghGzyE0CHEwlVgFArfZk41
psFaR2p26uW5MN6nsDKEcY8DQgWGYZRO3hFqfSw5plSXBgl9Q4ktOVKw3Rkz+/bz
dJtnCyyuUYzUlxDBpuwKQu+y4USQGFAaW6V/C/8uJ+BMPt8clvcS/N7uxPuRwC5Q
sIHYOAH8JN7ZG4qybAJ65JddlLAfnW7nD8ZQx3vQlfERsSKM58SONyyFxmuyROYZ
NyVTFgT9CrShm/kckkcFY9NKbK3TAbZOCWcXAOeCYGtJiRcjk3TzeBE1k3p6XiMs
Le3liE8xIIBqQ2G/0jRuK3Bw2LkOvBGD/vT1jOfb/MC7P6T4khiP3tqp54FHqJMn
vFEKnAQ3uCIFMSSsu9c+H4DL63lwgYnSLJY9iHsXaVufFChHBcHL17MAaXNnyRqV
h111A1D1CNqZq07n3uO8IFbqxDx1Uwn+K/U2qRoxt0QO1ozyUTnkpL2GxHVWucMW
/01yPWp+TtazNdS6MKafsHgn6WHjmN0oD8mccUf8jtVWI+6NYbZpQzrGEk0YzWLy
3kBuU0lodPoZ4XywQ6jjSwqgAjPEhU968gjTo4TOJEluT+k4sROmzpSqGtyBYszs
leyUBrNVpEsDJsLSZMu5+kd34gsUQvqsDlVe39U+5NkL9RadaHUaubOEl3l3gtxs
+ikEHP04pjfEmHJeSDJPd361jYLLecogRjPFqFFBXHb1rleAm2C7TSVbhFsBPcx9
APxl2j9elQNGWv8WjtWduID9YXVYkBut6t/b7UqIImoNoqHUxb8mUId4yW0PABtV
O+EG3Pc1PcD8OcHy5upd2b6kipgXXzXR9jaKyh3+2jy7q75mPvn/9g/dGBFHh0vg
fWeptoLX9pCkSTeaWN5hgrz9kx7Jt4ln2HwZL8AyDjPzc4mlKFBhud6o9PnsnMlo
D9zds0tiJsGwH/d2TZQfqOl/tazFbb5YcWNrT7HD3l0lJ4zQ+SWdWpanvS0T6oAB
BHFabI7vTOkri2/k4+lh+YeuRcPlTQwtG2kzYyd6CKrN1VB6qnnBprLZSGK/S72l
x/5edHyCgh+zVUQLA/T/ywVm+p/oog9frOac67RdaUTRH6Gz1IcSddRaf4A0q497
nSapZ8x2yWU3Tj1RJHtos1mgMoU2p2HTfXiVi6xgV7Bcmkk18MurecT7JnArf53b
momTTdlHosqq10T+NehoRd33CacuysPRpxM0D0qHM+cm3xeINclDjC8a0pWQH4AP
Iyhj6zArdYmjMXdaHlOFz6YZ2wvXsINm1budvISD7/OPEafH2/TWCBtPb2tyO9cN
AxL9mECimWNmnubEHcZY8QGymeGGHhudtQBqS6noApnuazQrD7/L2YaJYZZo5HuX
p9Lwhf32pnGr1foq9QFobJgXo6bfrYecrhxH1oX1OhuovPhMiEUAR8qmkNdGsOGV
iU9hNZp5CEHGdVp2fFWzlfW76qmtKimT10EfbPzS+/CukJ28rzi6nVm7lsUXMjQR
mCTqoQZLswc9z6nmtGrPCZSsnE/RAcU7OGPJ3OIYgMN0o3lkfSHXgxYhYjifl+Dy
HLWh7BbNS5jsjE4yff/HMvQIFJLvgsIbQWeJjQ7O7GbnZlcgUQh01WvNBeT1Ksb8
N0Fsqvy4O+4fxMFKgNwamGJHkwxfK1NwWlc18ZmpwB6949oGs8Ldb+qMKaRGTN6O
YUxAv7lM7zmffTaCkiSxvIub+ErOXlXJOp3NUDv7kDQdMfdCKpT8ytsBdp5039zm
IFBJKslwBEl6WSvU7L7VMPJOHpscXF/FriOHw8JoH07shv5FmUUKhd+GhLAjQ6rR
OvVdbDsYYDvhnefg4Ay0Qxhht51Hprlvqyuv0fjoMDKgwLn6ANtSwAvfE4JRY7Yu
Pa0O4OzcI8iuN3Pd0ml+R22rqY5W9zl5Ynyh2YuIGCapv+UP1Y6XB5s2Nmw9G2sc
7Zph0cLEFN9FN88QR5V1Kdkc/uv3Ku6RBpbUPJw64nv3c4gl5ETCC58rL5aHi8o2
vuhCow1nBA0T/YpYRWMoPpN7EkOqlnJzxeWPOmf6fPlu/7WuuwP/O5JOwhkm8ADZ
crE+7ehOGrClseY+pgcfG6z77VZRxMB9jXgXXacTdb8PDtAvPsOoR2RziKg20WcQ
tMcWidGmpiTdWahy7ojpdkoMNEhmAcRSrqQzH9B4sTMxYU4NlmAuknAQ6YkVEG0D
jmwRWcFLFA/OehitIEhiWZeHb1ZjdiNQeBt8hQJQAAX4w6AXgMHZ7uhwpOXBsyHV
RwC2oeVLilIwx+5p9g6d11SEfOkalDZj0dLjakpXGs8u0OoM1a3EMggGVjEPqPGx
XF52G5Rm3CQpqcVx6pPV1lMw9NzhZdQZxLXPGLRBYKngWqlVHe+C0mMJq0HgLup7
AALIRD+clZH6IIY1gGVrfgJcEhc0DSVPSZLBLcMr++7CM5Q9AB7wwA+g+iw8XeNs
z7XUkVAb3QeCOdKR4uWpreQuIKowiYylLPgubzwXhZFv9A5I6M8jcIyFFf1NC1lI
kmCQuFL0PefC54K3kpOyc1FysyOhgk1pBq9tVhUkB08eKHvZ3ZB3GSKgxfwjmciW
T6X9H/72Rtdt1H9IGECVROtyopMko7/SgRCOMcnQiGaEBw7CwG9s9TLMn4U7MiCb
MjH7TTlcF9/KzMe6QvMgwDBg54XdLYIegjPZC9vCFWvNL0fts+uYungDWlqyRBZM
vJOgwVaIhc0J7eMnasbc3mk32ZelIkruro0zFImHhWoDn6dkxd2DPH4ndzaHkTnJ
bhHBitAi1qq8JPCZChEG9C+J2MLUdeBFbb0qyIdl/rWhKgK4BUqDlTLc2B0g050I
u8JTXzt378Uf7SebugeV0w1HW7asUyDGQtR3XsE3Q2LfINnFZataBLOsRr2DRUC9
28XwrQfFzU41/vmIfS6Fo+Cz47yyNua2vhQhY3AQ30XFx5yq18yiYNOPrH3flMhi
0PpoYSQc86IF+206CsXWmTc7ISsQ3G9Uku7HcKdGgY7xCdFqjU7ao7cnC/Gjv7/i
TcW8za3MKNVnABawWbf3gkqoZsXrrCC54ORsZrAV8Ew2DKf++JJJcgyli4zqiCMK
wYcVdleMncmP7ST/YuVc30QR5jRomHLnWXuHtFxABXE0HH4ysChHK1q2xndRm/9V
eQ5chWZ8p5fslOEWGT+Q4tu5L9hpZQkg0aRpSSioyxRyaq5LomTjbmLoQfkdHxUz
VpGq8iQ2gQReXAoi6w4Nm/9Fq/Xn2L1bq1O5sD0JGwODi/QOdBHuapiu+E2gFua0
2h2lc3jg/6bfkVBTi+yq2YBMGjH7StWoJu4Pu0OxjtYIcEAbN74JXrGMhNXqT5u2
2rVsQ8tPsdfP2up3Pkbli640OVXNOsikkWqa4p8HVttUzHhdn45JhQRZqbfpSbZg
ouD1Cya8NttdxKjdHBDpaBgJYe0DtMGXZQ+DGOmOBmLpx2aJBNAdkIkTp7LLyk04
Trj4BncDfVQFQVXDT3QiCC+fFtbijDIJpKGr1dWWw+8Q0pDAQT5E0ftIEU2Zv27L
3gj1XJMnqT/OhZejzjl7OmyiP804GGqBRzKYbDVyoAn4NvkotHYZj+HoFnFQR0EN
2xPylvnPxTVKXII+dF571kt/JMCi7kdG+box5r4+Y6vSg8ArCO+yjQbayrirVJIr
oSRtDHG94k60pT/cQZ/AGAjdwpMwEu259xsmo0rcxtrW+xeeK62kKCSchNx/LjFW
DsIUXhWFqfgqSYwteJUHZ2FNpTX6qakUhuYwPVYb8t4VQH7pZNU4YkFUml47reSh
4nCJ/6Sac3U7SuO0iKpr1xtjcaHBKt3cBSyP8aNNVl8bDhnd6imbMx3tH1psZuVV
rzAEG2UboVMcYEtcA7JJpcQtvgK3wplOLhQA3R099rNDI/u6EJnVxMNJ3YXK4jWP
QdSRxiPqr6TKtLr79GtZcM7qb4ocRUe0TLCzCikxUjmciJBYChccotM9PgAG5/e4
m9D1/ar456S/A61w4Z6gfANPihps/Y0v1nkeEwuaZSc0dSwSjNo9Nup2Cs8sPj7f
nxlsumPGJZTabhvOxtUdgvvj+w2f322uzRfnpF6bUN6ee8MUQzQRijUcfC4/WS2x
/VzNV82aPQ6wYz5x5/gyY/MHJpQD1YYo36yW1dUQrbI76jjvE5VwvMsduqRPVuEJ
yk4+ft3RwWUHy8GAAyhP9a11cEBxU2E7wPoB2ciwWBQh4AvY3vqEeeQ/xAZ93/CH
vFiffn52+zlOOWixLqTyQ87Sidb1W7nA9/tc4ywUT0S4btv1ppbJ/IEIqAYuknhM
iZS9i4NV2OF0OhMhGQMVgSrYerhxA8L3IyRYCUXt5QIt1TPc2qHHiMaFJrFIsEnb
qnXCiU401u/Xl4t7YIDJDshgTLtb/lF44qYSApFakHGgxFrNmpKQHOf5TnRP7EZJ
LmCSW5EqEPv8EkbKXWvUvjqEsRQWlESkG8jsqa9+zc2YF43CHzAqW84BYDr8WltV
OYZfoETR1tnh08aZWRD/7ardOQ9I8Hj4Yt5XWnbdeI3j6O04JyHO+0vGiHq+4Rmq
jwg4SSR2FJR0RsNw7Z2JRhr+yCK9wstuyHmob18oU+j69KV/vKMeQIBSKbsbng03
q+zd+q4WR2fijV0/PXXs2c+AQsy76mIF0juitTv6+fSQHWHBdZZ8mVUpV4N85LBl
ydeC9KVZODkgAO9sHTlqJE8/lNGjUpUQ7e3wAHEaTVaZ0d9tg0xinMwjqDezAw1G
owdWJcGW2VymdXNzTwk1lSEAp38dwXrGlOJBODpZQZjQ7CzRsZFe7YofiK60P7P4
+o7qBtcJwGCmHbeldtDRA6QSxqrjfKOAhux35vCQnSTMS9/Ch4HUCUxvTgwEMko7
4M1bd02i88+Wl8AP00/soM2OA+oW1qU2p76X2PBsR7Ie4/Yp18UXvywb+p8kL1pA
y+mdk7b0eC89+2BvlcEAkRXyJctRU7GNAChenb8/xn65i+uBcN3XBzGXI5NaP5zB
8gAZJ1byq0YNOD3UigwbrO+EalmQ0i2v4ikMpCw3f1NmbQZqh7V1MirnW4t1gxwz
Dy22VTPqBnxWvwbNMxVQENwzO0LgHleNIrGLP2HKZzhUdyzNXbwzz1Ut7Tp0scKU
XoZkvz42U5bKKiiDzLESIDOp5CgaAbTo9LUDDbhVQEDH/xhfZ8gGnHWLalpkjOT5
thlzwn/grdow4UIwjUehqyYCp4kSVLeV8rL4MXo4U17+tL5qlaTPd2PcrplHDHrz
BYexYCxDF4jM9U0AQqrQbjNWDEFFLC2yZNUBc76OJZnUyOXcSh6d655ILK4aFxHL
sZyUGfYpFq36yclqP6VPrp1ELU6q+7MjvRaNJgezOMrdXuiOl3rIMzvnjepibG1U
pgg80d+9lZ6r90culOftgKfcSQwa05Qhk9TN6eAnt8xONblnwnLq8W1xiTp3qz+x
94bFOPAgJOY2NdWLZ0R9r7QiBTxDPcSLuBYNJGiYvIR7sEobcZSRxwFg4/lrzLRf
Dk+cgYdDcz1gYE5eYy3pXJ1UkSC3lLuz3KPglClgbO9Zh1TYFNEEUm0JVAczI4fL
D6iJ2e0I8PxvTeQPxOdEDIH9+TeD/XdTkZxaKZYcit5228+J5dz0eDE+E7U4z6aK
mrgZNIw4q2YLU+qo8aIAL7hqpEfosxK0qGw071MiHBSI1kzoscF6gSt7bdq3DIpf
/3oA/S7p1lBukIEUZFUQe0x2vpMmSYm5PrDxrqDG+yF6r8auz198rRhe94IiGzSF
uiweI+nlitE7IVc7oZP7TMnrYeGiaWdnrBuatZEkdyuQKEgvSnoAjp5IyDwZeqtw
V+QCGGR7HGOxTqDUAds/HYWdq5onUfNnp41ReFD+EBilhtz+BP4itLhi4S6qesPh
kIEpCX6hg0FiBCi1ytgALSATLITtirsS8wdV2CIK/W0fWQHWWM0jIrxzgUqv5190
oJFI0g3z9u8FAIpJwjo9c+dBxfSkfQ5j7UPe/AdAkHBVE7wimCX6Nk5ViZ0x2U1j
xXixGoDHuQwBZ79beSj4pSsrS6G6qaOIhJUMyxB0N4yaN6xW3DiWHzksgbn9MF21
H7OqcnthNJXuxz+CxHxq9enoAC3AHjr5732ClhGCIvWziAKmNRiVeyEXaACniHOm
QeFtjbDGU8sy3GdrcNXqMHQzjbW8DqIySCVlhBq8VFW6ybujDNSn0yPeB9ERUFcJ
hLtsBJcG5J+ewAz9HaNI2Ornp5Q2DhXsfVkVttYFn7wIz002ORQ16M37pfrzebCc
ulzweLgcAYU2fdm6vBstgp04T2RGfJO3d8o+DDOUR5M7Vq5j/ayCwkG4UCiBig0Z
Wk6n2Up9IbBSzE9hXMV5UT8ov1S4vDmzFIu0ORW5Cr/f/BOlhin01I3JcHNXiPmh
/P3TKklrMhSvyxSSPEhTjAoMLZ76B+yoVzQjfuju+r5zLF+1DVYUoOx8mmQc1rEh
tlZ5dkB3M3bdMXvrXZYbJx2P+Fua+ZpXAwk6lmkmtsDGO4rtuptEhmzHAqQr+sIG
2OuKW92XzDS2XeAagWRLRnbbIg4ebhwDXlVM9V5FZs5VVLH7yPJrklTCqHPlpdKg
ysNXCcm432Fzi0IpXh03jmQLZ59Qn3Y/GFHQFH/lzHdQguqN7FSzLyDbfDe+lKM8
4MmltWb91NZFm3PE3LFNj6uFuld69ooKnbBBe0qHgWYatiVFAyM2bkqx5lN3MJ8h
c+Klx2Qn/TDuI/KLWv0R/McEqWmx4vNJziDqWvrRA0cK20RFpPorMuMzYer7Rf3K
XFpeVBbVz4KQP1PJsPU2cZ+vtWNGQUSrs24EYe3XF0FGpEdaeGaTRdkNR6Hh739k
IX63GhH0jYwvhMM/cfIqawssiYq60jMyKKdUdGf71PiaHZRNIChtbf4sj3xqwPgF
QmJJMLYZmD2l33WDGGJSLHvU7gY+BldhxSzZDn5S9Y6VtsKDqblRZLSgzUovsvL/
mBLEMh/rDtFi7OY+n4hxdoKfsOA+o1SZmdkusZHbPzbhqccNSag42J05CFniOOgO
5gMOcizIsoslHK3IZhLYyKfV09VrqUvei9j4ElTpX/Yas4kKAl2YNBc2bEVttBoW
gCqhqvGEzcDs0nGdeiTplxUaHnzJZVLTVcU1/ozTgm4lexKZ709hu4ux9U9JJBJF
hRoaqL60IKrtAqTTZR2XCer65lEjWH0djz80p75JIo/W09ol2Kk8s6GGXNXjo20I
C9HkZdP1c9fHmCM3uyMt3u0zDNfdJoATe4EFcArLFb+TOgH5CCYgwVWOxVzIskJi
2NrjnIEtHvRTVjj6ORE8sJVv2Pu/4CuPA4MxE/lwaZ8AJEN570pyqkU9fP04FTVi
vkqlxG+ynGKBBlSzgrijJ9yT1sotoIO0PFoEPB34kA45C4TZWzm/GtxYp25nldov
fzWVowNey/ECvKoJhSkwBDAkzAYDO6lz4f/gKWPy7U0MXmluxtZ6w4o/CCOhj5Dg
+GBZIdG9DUjPz8fuLdtEX+NofQlIuYVV2BsaEoc7CjZCjlSbXjIh7TbqaI2zGyhK
/pKRbTwo7x/DRPKGHfhuFWuUgQsn4fYnWmO5i/59YKQxP+lYMwDSzcIKI+zPqDdz
OSblqZZoE2HO8JLHLM11A5fdAsKIKYx6HHPL75U0jbzDVYE+DRnbCRTCptDMOQbK
9fmOyJ22OkmVpmmDQaEigFAUxM/2OtGcUFE1H50j1zvJVH+iBTiedaHiBH1xa/6f
Nhxt7l+bb4d8FrqhS7zrlRLhawbb/vXcMQ35HTrlxWr6wSffaf4c7MWiQ51o9ang
Jrxjx4FpNsjPxrmL50tlxZa7DMROJE5DsHVVQ4CWjH9aS27GUI8QB2bv70XcqxjD
wnAliYdKqapG5tbbHTEzwlQ97UX9btkITkk4Bad3ZrsDWMAfR4uUo9wChF1XdNDk
ipMguByXPAGzrui8sVo794595yF5wQqMcnuIdqcHYY/BE/WhxsARE2AFpw3F0cB2
02SmwU4o0ysE80jnl8ZDKDQS20goLg/Yza5A3x2vzoTAf0Br0oCryz3c67gIVgHj
RMDWuNGAtDt4D3DMq6oruf2FH9VhsXyg6PWRDhr8L6YcIKbhuV90id90ulUMebOU
0BT19hozhNpPXWJQ1HkVO3qp2c60n0pRXSVDdl1AaaDPLObqjMqiWaUYQDV0lIUI
QHf1mJEFJyBQ9H1C4bG1hmWQ2ATTs7/MapXbiEpxUWSxqQ2+gwPnsTRvpE9V1wxS
4V7uFo7T7mZxtlwCaXRPTrnY5sBZJXEh71tzq1AOtseEhwfTstwKISRJUvY7bHls
efz7w2oZIOWwNTdiP27o9K+g79lqnxtFzgS18z7mxOctmHNtL2s3KXgmDWMTOfib
PW9J76m8ei1buV5MPIQJiU8HoqugOHTSmJiI/LhaauWBokjOjnE5Rwy67xxenn4N
IRoRRHOkXqTE1PtVBIs9OzZMwR89uPFTUiDCQcEhJGoJKdjErsbrGnSJz5LwztFd
nVLvsmLXuWCIAlT17ROV4mRqChwxnqJzDZaIGm/eofJ8W1+bcVpeocWsjklfrG7R
ysROGWSgyE4f24oQbPoUNykWqLXh+cOB/RHvgwz87tOwkJRcCYzR+ymT+kGWYBIp
O5bAV3+Qh7C/lsulIN4wvKevdI/sHFg4VYNCjmS1gPewrJCaDwkRBif6iznEaXU+
BWdC73Si/jNatTDvXTqDpAshNg5TER/ae13sPyMMGHiqYMEnfPgW6knfJhdB3Fsk
7b3P4DugjsRGGj9MyVg2hXRifaW4DlH1oC+C9JkZrcBJiyPW+jT+ey4kLllnSvto
XQgEk4AsAp0nDJyBa6HL/fWEMz+Tf3K0O0reiQ5uvtuTq2TTloifWtL1rv8MrfTT
j40i5jxhKQm2W9END6QAcYYng0ZXBiJcCtb/SOCK9ddLnphqrEk5qvpPVfkisluz
1FEMaSuR1sdHrYuo1j+YvVmHlT1sYOuxNRZdVR8HEybVmPeC8xtYBRnGldkqpLiY
IiBjLTw2pNV7u4Lq/hbf8JyDP6S3tLynrCiaurhrHVYRse+kRrol9qQ+hVSWlLM8
9HCpI1D2WTMGEJMcu0kNGl5iHcz/q8ytgqRjxTPsMaNWdqJkNprSYiZLRn7mP4rf
+5g7UbL8C21VFh9O7xrvmx+SpkqBxxgsqCecS/cl5/pPuDeHQaY6cd5lBxfVdTyw
9MEO2LNDhOYvEc5qPPw8lkXnfTlE4hSAhQNqFYhsBzoNbVw5R8lEER3ONpQOBF1J
v/BpBW9STvV5j49l28XbLNxjiVB8Vvr6LxehpLfNotzy35YFF7lefo/aDKAJYn5V
NUKaEavjPwPnnNb+F+p/XneK3OvlvLGP97Y6JPOLxMfi28IKax95igBuuntN8BWQ
fKCh5Iswz5hZmiftdAXfkIrzqtzZQImMPRLt3WzRcDSl46LsxL8ds1fTY3Fur5aL
H+9IjMs+yZpPS+TlM126gC7cDyD+I2XmxScLtHtbUiEV+PGAVyCI/YPYWyu3GjLy
2+AL7iXg79kY0+8nORd1vAtxrMD1WTNEZn3tSEw5qb9ZHs6T8q4iIS0OBmFXulKm
Qr4E3Vge0FXWurmFSEnH0krhYzUXoHBnR+PWIbs33LAlBVXny+IIjzI59rYQhugA
6J4Zpp8AN9a+PkwAWXphBi+7renuk2kgySmv+zfSygEAW0+ftoObb3HsLX3WLADe
K08caAOhuvrgtisS3/Tqz3kbguSCOh9fp9l0cA6Qey0PUj2uzs0PaZp07xlbELMU
vSjIhkCJazvePAz013KGZSMnr1oaK1eKprZ5IZINn8X8Ja/SNKwXT/tE8lbBwpZe
zurZFMmlCt4gd0gDWtYtBQGbAlM438Gf4+wS3DNti4cs9AphUD0feaEaMTD9LtZL
NZ4+KhndKajHhMJeSCOUmZBHMbWowQT7OKeFKVMHG79clIov8U40r1dMFswu+GKy
sQeOfy5CfmnkDnenIGvCwZ76AJk2Rn50n14TqRuucGkhmHYP1wk+fBYBLpIuHKUo
BVq3Z1A469J5ZeB7NhAGWwNeTGy6aABW9gpVWLyZrc2lsQ0GV0W+OIK2sJOeHNYE
ZV90hAbPyXvchwdew1sWDL/M6NUSB82Pvd5Pgq9AehIwFbDYNr9uJI9AihsNHdog
6bbtQhkGGsV6gF3pVO/WeJ40oIJqGPNsN0+nuacBb9aJ7TigioV9F4DMet5LRx4y
whqixBrIcs9lJdZx4qDcdwWgN5OEcdd1fCWgbUmwnjAOa5phwUexSQBK1w96USL1
1JSo+ti/aOqowTa106uuSFBtlKau4Bv0ugcHjpG0Z7iU6rXcnVdVAxlpOGS4Sz6O
8mJ2cdNT26h2WXMmIMgWUrSRZJCghrbDpgoPnpuxkZ1lktg0mCgICaBpuRLS4R4t
6uqE6KYK+GPK3IFWZ/L2qqMGOftxyaeNn9VagWvftyVUoxRg7VZYCHwxv6kKFtZ2
vnSBPglL03G3OGy5D2yzDs0ec4YmjeWoUo9p6BoitdCwyYLSR0WeDuwJUoHwDaKi
3MoGZyAEJA5JwBDoEEVIKFuZp3bw+Rxa5smiZ2YdVVfBGp4cQmsSPvvl3zpHoPqG
8edkwdYLwuA+Z/PwU/A/hlHASZiC918IlizbXl2nAYQzRinG08kf+97tCM0Klgrm
RwHVPO2ivXgvg56mMWmjnWMu8Zb825Q2MuiTMbqIPhDvmAZLJS7q1L61uOPS9PKm
aXU9X3g4jNyBsILcZWJQVPkEAL3cw1buILOwIaGONlWN+hRqYAmbwwz6DM2GAS7z
lZsZuI63QSc8gtbrY24NrxidFVs/xJH/lCwz8D/8gGBQSo5z+/iyOJpGePW7Gh53
0c+IP+LWWeUKs27McsMCJJXIJhOvGpcoe8bGwkj4WyaF0zitHNA+sldn140iFzmN
V0NQb/IiQ3G100sx0pu1H/ddkYKdYTNXzLqRThom6T9+dSG75IsCLm/1Hl420O3X
oIwPs4hYcFoBIYUu7uAAq8c7Q2I0ycpofrl/1zpq4aSpY51Wmx0r64phztezJZyz
05m/aCvMdze9pkbhFAIoK0aeL7wqt5/47u9lbnpeeRO8h0+VePTlC/aCsjL0obZM
72w/2c/+oVJhuZUb+p9hTRzthoMZndwCOE9KaXau8nBzlr1R2ijh1ZWqR9+BO8hU
S1BaPDce+73YHS09wiNInYDk0UPiR7T/X/CqHldE3ep5fT9pL2bYognYs2xEq56I
km7p21KFegWxa+DjaHt5dJ/OjQZEuVc0pG0jHPq1ceGqQDZa+OgOEkda0PvJQu4v
7ajuUHOc9sa4VZQyitk/RNUYMrjXjuQ40iNvTtkKWSkjFl0S0asKbRolUPyfK2FC
hdbrhhTJSrTOC9DWxQt/rvraCnj8ryjTlB/T+sdTeBBYdf9J+A0rjrCNNRjdXqRa
pIlNrdagrrctPCkaD7cxPhbW5pTe0sK4aMsSD14S4RQu3PkmWg9DO0aBjCLK482E
t+8FBZQh3Id0TkgZBvYNApRw+z5OAV+l+qiXLW0kztPN4vZOI54Tpj74TpbORMw7
At+IK3ftJd+5iLmJkxax2blSQGkIKu5b/8ryst/diktmWbO0AkefMfVIEE4IPIQs
wUw02RSCB0F3rq/XMOxtHFHSjTu3neE5v+oazAYxte3QgIosvzp+cQs8LM734F11
rD87XlOyBmfFynocyVOfZnA4Q6Jqexg3jZmMJiamM3CJ+fuG2TfDmJBjjw27zTML
MoSjmXCz8fep5RcDoflYTCWDD8MZZyj34qfihTqDVLUQAlWSUiCaKNmHLQ8hNiWZ
4+Ba5GdZ33mr9nbLw8whU61l9+8tsrb8w/F2DRMjH6MUzdvVeLFtHNxqk39sKCOD
CwdgIMRYOe/52xFRzqWj6lSSBjjNnm1SsFr4yTe6tHHqvyAb/GHY7STh52RyicEz
bkeSfyg+rhToU80j7IAyJBgaCODG1f3silxHz+OT5p+qm/uYSau2dG/RxSKiC/3E
vpIzO41PueK2dJzpQ8XKmVBB8OMBm9ZgHzYvKK+JCtBEZWjTN4ZHwyBEGkrZl4SV
aDwXUiYv3UL9hzK2ecjdZEsLVIEQ0Ha0PuJNs1CWMagvaOBiA7TSe7TGNjWhz5C7
BG6SA1D9UHBXLggCLHFvjiTYQSAolaBrxnzBElkWKFIOUQ5ZjPbsjwKnI/fAttGU
K+Q8DOSMQtZEtTMzjCVfQnp5FTSSrD7bX7WnWeETiAXWkrwKxCG0ZAf8FIOLH8SC
h7jzwUxpJNxi0C1LJt/dRo2Xh9/1nfetVHdgukXNq/wuHAiyzCX+nxWHMEvDs2pp
6fR9NAQFPNFdRY/wxeeh/3a12xyOnff+xcRzX1evXIESxxLqDtztOizUCyQdILSY
kklv9PSgphSpQNyPCog7E0eExBdkkan2UCqIhBOK4cnqqbEapnEBO/owuxQXE4ay
hbru4cah2jK2vLjFrQGj3XGqG4+sfX3tMzvAOep8c10RB9p6jTvMc48t8X7PnZ78
38eudrZc1aJq+VrjC3Wozk9g3W8fu5ltRpD7s3zCLHxh56U86ID6iAUxHR0NKlLk
DqrbhxIj0eD3Y/FzbSUA8vXD7kNbAlOeYIRtP2+lQDbIoCcpBuvph24tvtkMYj6o
h1lkEu1FuuQgbyBg0KSJoKm1kRvKAkceoRJZbdtlSrMyTLrJJUlSxUjblBxATCk0
nn67f30Bk5k74lAVJ/+0U827co1kTyOgyo6O4EnB2TQfKLGSuCSwqSH/7edX01AN
VOKtS9d9BsgJ4SczWIkB6jySUKfpuZybwkRCytcBrsjD7XxYe8UaO/JDdo+T5iHY
ZGSHUrO3bNH35ZKex4Ua/6kpjUWMRjsxJX0ag48HF9334PMkP3nUwSf3Qfg+uLeu
niK/a+0HGD5Y89Hg+errR8rXlOFF2jOlEm8UY1N+PQlFtoF6Fv+ly2Xty3M1Pz5L
np7oyXSqzG3ODPDoMybLhZrQqfSBYwFQYCEdLPwTinzZt240ITc6vyfwDXJ/LBkd
0FPo1KH0W9M41got6Z2l162ZlMcCnJczjN/hQzsFsBMTJEbtnZ+0CdpoAvp7xWA+
gr6jkaiBXLi+9+Y3OaL/VRtVKeFagpZJJ5oKB+qzsOm0HTuq6VV/c3Rmz+G9i7/b
MS3zVL/09VJAiWhIcFy3uv/CHIa9Mou9/J+biOX1KBcXBLWMVQNCXM7q679LWyJb
jbk4Ijdcvp7gw2J/N8PmhACgWnq3iqCMzyUttE19jVZ0zpLrhTmkkypzHSfJjqxm
XcboW4Og7xt3ejCQEmg2WZgQT06LYjBy+/fbcWz51pCA8Tmw9em5fewLc4lSuGm3
oeB0P5MU1ReZpDfdb1YUFPqCudPC8O/SU6BuZFuzrtQAgp16mmKNlgoB2IvbxZl7
8zNSIQxB5akdXeX6sLS25PubFOT5Hol8kvgFKAZ4lsAxAwFiUFJn0QBSgoMOIVn8
LW650lKvbqT3UZJRwnIIyY60R89p6L+/j8ghhtTiDOk+cJ/W1eYZ1iFePvlPcAvf
fwGVQYdlZ4ht9jnSfvq6QdZ5tjvI/7RErcSOf/OUiahoHkUv6rxVPRvARyuQQE9K
pvGEYCHFlMKWIJcUzVo3D+ykqXqHWIw9xgAfrsp3O/khub+DyMOwSs3+Xg+8dubc
KfTMs8cwEuSJJRXkWS3uhtJPUzxjrmZiXLoNRQ3pEIJMTQyvBNdZy3Vb9JY6fJ9r
//fWjEPRkAgPWDZcAAhyGEAF8lP19JPbHFsLIXRkbrgmqq3vNZU0ShL0VKcsnb3+
UMC4rHbrQ2bga0r+KpqLxWHFo394EuzhCAWwKEMz7tDdqNFsgqZbQm2St+7+50fs
u5bO+ucjiO/zY/hJAiovVJOiDrfaW0mhxe5OAL/tyL7l5Q/vbNuAfVxB1j1KcfaJ
wEt04g4TXXN3s3Hm9TG17mu6jpz9tGkYQe97qnnraJVYAh3obDqriGXuAV90tRhQ
jgfXUbCmQtKXR1BZ01hRMyM8skJhlDCkM62ThbXkYRcuuUb/AhbiBEIGgdpB4q9j
STokD1dsTO3MuriWa8P2SikyY6uq7KIoaGwvbb1n679IA3F+Lj+6B2Rb7QuQjIig
C8LrQrqXScAqG83YXjfhpsQCXI6HdZNpz4OONczu6N/iSJLFT1sGazYR+EShyom1
pNJGMFIOkW8+2Meso27ouaJOuUEWi4jChvH5b5WLPrVmN/PWolrpjdTg+z+dowlo
2o2y2FSceIIMWhFVBqYeMkCjEsao578aTdQwzhE+B8YFiWZckU1OBmgALVbW5BTr
O3PdUlEBz3qoIec+6GjdA+utddS/aGp4Z6rB67XYdy5Dj1jyLehTkhuD32b8GVLR
bK8KTaloxH4aUfIZ2D+K6tssoEaqCrYuM8QBvtCvMLiPEAXqUwoTQvyVCXbbzo+t
0QxSX5uqbMJWOFUaaHrQOGQFio37C8vAU6FfqRnkhkaCue+xq+CckegTEWzC1qsz
r3pdpe528YjpL3J0XOf/L8IBpPSHmJUTAi1S/DZGTJ3DILh6GONGged/Or42KM7R
kSf1BKyNDB9/12RmOSVIz2VkETPijHPTZvOqoJrze/8ERMabA6n/m2RZbnuXHJqA
e+FnLr/keybSfIL3h+rvVsX8cJ4V9nTszlU0+ji9OCdOz8yjTOdWoFIbsZUS7C4/
armxckwtthpa8fAIEars1+lPzEbPOxODE2aoKHD4SNxcSeGubwX8qftn6AjSg7wu
HyWNS9S1UkBjHMwqPrSzJph+kiG7FA3Ozz3twQ3j+pMP4tRQOGr0t54MhPZ3r0bE
Tmh99mFlXSA/aftUX0riyYGq/icuTj2iayLQlinc1mMVBYIdTqVVOYmtO9E0J62J
KvVNJrYkjJYslqrSecrqXDlWV+iOKvqL6nPivvSpnmbVTNdy59IdkYH003ESTx78
40vYpnTuqPEvL0B7hbMz4MGjzeVElICUROZMWjpPu4PURcw+34n8nPonlv9O6KY5
tePraJC3+BpiGfd141N+oud0M8AarestPV6lqxDogdN5kzzez0+4hSYvE55CWByx
6tey5bKYT0FZrqfQICtM8+xachS/pKsqZn2z5ppLvIZw57X7576GmqlLrefrZFma
G5iHFlPHT9NnUDULOwVYD3DiLnpfTS+ixUyK7dCT/XP5eoI8BQzJuRHJRW3ojimU
mxKPgdzmdMWz73O6ri85TzN7dbldDji1EWeuV4GbKUnx7AXQF0AJXU26A0rzKHx3
WURbpwy/MQz/9V1dDGd6tc7ubid2XA+PI5zvf7ukzn3jtDLdlvDuYeoXxpCeHcoO
db6ivoPZ3Mq2YbVoZzRDDVpaF6o2BiZb0d12WVT77SUmkeR+gsM5Zk74A1J4uych
UWegbeBv3ujk9+du1HHt4a6zbr9/Kk6cPmn3HcBwrJ6y96SMp8V2m8thM8QU95H9
qcYI6e7wqIEe1tmoksasuQg+AoCU0bwpaJ6NwdZMNVROvVsS8G+3kox2ms13XKcm
Zo5ZwAaJX7/uXE4vfv0h5CpNHxzDe2z4ifHn4x1cnXr2nwnNXj/MukiwxF9/N/VR
Ic742HLf+5FfKxhOFJLyIFDQIXz9brS53BjFZ2z4MgrHp0wpmgD8mirUGmSzm7g9
upQpzqKkFpWoUWWGg+y6YOcc2wWWwDYmZUj2Tz5K1b2FUuKvndqmTF6N5EmummB1
m4rMvArK9ioqBrzqU/Vlulooe2fLR5r0F+lu7VzYSydzgU2MTGMSvNP/VbLWK6+W
RBYJm7JlTXbbZ0eX2ckgcwm8fCyCekocIfD456G6MoV2B7n/dHnST9BCQflKOX/4
0zaK+ZjTn7V32EIVD4DVtPNuQWSNaSyQ52W9x6lgEmSmnNkPtLjdjlEajVmsAvDi
1MMPM0ygfwvXczqhBKXKupo9Md6sw7H5ZVBIDiOp9QWCorJZLUp64qgLyox9pzFc
lDkcyd1SFL3sH9UK7MA9NbpkFA6Ob1pAUewIeh3QzIk=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
H/eJ5Un5Ur08Ecxa+wuI53b78sfCE5X4AG7oIFIt1RbPlEQQG4frkeztV4FdBsPW
cjXw4Op3qAebgjJIz8gQsJ19WYBE2QC8j/+nGlFs2c/abKYiuORxKctoxDH9QHNh
sEVq8EtLsHJO/rmP4dziQxp3hwHie/E3wS3rw+lxLFv9J4JNVWdndhCjhTawklWM
Px42GMKqSbyDxDr2wgDFg1U9PPoCEtosVHutO4HioTIsuLSIaKAV1HqNdjCCKBSF
NYULnbmmDX1A7uG9BClompPPuyizZ3BXM75MuDTfx1Vlzp1+h3DIygXu8o5bHynO
0jjzaq3kSUftR9wtn/O40A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7632 )
`pragma protect data_block
eR7Sxgmx8bdADFR1G8o6kWcqo4OKIT9/6c5i7BNO/oR9u4TNXJupl2PxJTSYEHR/
ItZ2E82rGmBA/9MG30BvRcx8op10275Ny3jmos16YFx7CJd4gHCJBIwwMxeo8CJX
+JHI/Q9AI0cVlOdqaPdMZ2rQ2pYfI6hkd2m4sbYcYj5XB/6qUDC+NR58qjZUIv2b
kF/opNLAQVlfoJ1rxnjR3eaGGuvizYvKAVhBO542Hyx/gsLkLO5Rzx3yFAhKGIar
NMDHH3TxQKC57BK1JCx0rE7FtSjxiLRf/84lngr0bpUyjDukSnI8gJX3SrP+4xd7
maKVuKLqOaHtCEPbrKyU/s4eCq2LE83CmyLbPxCZOVUn2kNf2TndX6ipnYGV3eMW
L3h1zP43DWCN7qQYbGdvjK6+VNmu/r10NQYeNYsgi0VydWfap/PNwtIhJvGgAKjn
xZUh/vKi3oaAxw64DLw8Tal12ynVCkpDu+wLTRfPbHYASxhIcFY8B7ioftrRgRqr
ewRqOLy9hrBWwLIV+cIVoLn+kYGimGiUGfWa0HrHCNZO2EVUlTXuBPdKlRg5g3Ly
Unt9rHr/z1FG9aomi6046H6r0i0/tkd88P4Z3Z54WC+r8jHCLSY88G5/c3eO5EYe
hD7nrCk4jSW3aR3gb9rqypq8yO3WnE9kqolf20dnjduh/2hrGzJaWVMi7Y3XM4ER
juPWhZZGWv8yVzcobz3C5/Bf0yHw1oaoU/150SClubSXfnM+5k4X+5DE8KNB1RZT
bEbqvXLIVsQBaeljpPhzqV8pKe4EVdpkgObGWEEl2hYFeAiSMZ9/Q8tWQUhCG4/Q
C9aS88u52DBSN21zhqxFVYSVpCq9olnC6ZEVwgzvV4Czi+O/2YMi4AW78/52ZLFW
yxVVpN1WK5wAcAeCOygbQuNxzcVx50Y2j+VU/jTs3UTCcL+fRHdX6KdXWVHOUmAW
lBfSzzgNHT4poi05gyH83hfFY/qb5CWBMGrFWQ8erk1p8SguP+afeNmKa6Zx99W0
SHjogbdZTD6eVnba1uEmuZeCwCNalGU1aGvcbeW50e8PQ5ZKaGNzQSbLDtaQEepb
lX+k0IaE36jTgF/vf+Q7v4j6bnpBDbmuX/CAAbTfHmKeZ8lZ9B3z0Wm0XD0jegX5
8pXdrV5Ip97zM25V+ryQo+U3cG1774/XLipl0sgbHmP/s4LSe4MyRWoLAhE9KPJf
R1LTxbvAjn673hRLV2doiQB+9EwsQ2JKLqmaq2X6SY51F7AR7oybvvi0o3NrAvcW
ozd7qxNmPiTtHsJSohpDTQ0gYwIV5wUpd85zkfhzOeuKHUVLS2MWJPGKVBqoSUzh
9mCMgpttCpym58unh3OptgCZFJBQg29gEPR7iHkC4TxTuPrOso4hCXEeYMq0g7ME
8BAstoYfkNARdJJ9HwxtbCahvFJMcZorOdmw/+u2N7CGG+ef4dJrD73b/nrcbTGZ
x2XBanivx+zyLgnNgeD5S5c7D3tQQNJNa5nUTqVb6MTNqX85M4vee4tr83xld1kq
ns/RfQUCvp6rGeZQ/ChgNI3oEboCK8eixwAfyAzIHD1l4o+6aZwdFmSNkRGXlqbW
/Hy4mr6pYvnSlfbDqZBu7Jl7in1KNOpZKzs3xHrH9NlgupfKZo2h05I984GXz2AS
UxBxDkqyeHo8e6rwUVoUxiFc99Y7obICCMn+44Oeda3pNbBJo6SAo/37X3PlzRCn
QnE68Dc2JiEsAQVVaUV9cBvodL7BEW4d07Ed1U+OHgkbm3kx27ULdDej3eKKvVjV
M97G36gScM9iVdy3aLl8eKqFxIW4xJrNPZ0HF7BhdD6vBrxOwewlj+LE+Avx6tym
k4cvQXrqKmXGdazBShAuW/7U8s411eXkHCbJ64tOc7kmyS8fIZuqY9RH1xMDxwJS
Z0HV5GPz8aQxlxjH8S/7A5Z0jFeSj9O9/F1W18AeJ1i+SizCqaX60RlIAvTKYY4S
qQjnzmOpNxDrUVapdsPkLFBY0Esfo8k9bpVJPwMQIt1NCVn+gHoNruNQ1DI/GYhP
FXV50sOxRrH7his4VhV6Tjc2rC3T+qgtZFR1qlsbw7+0BhD6GFUhXQdmj/IvKOUI
6mERMkn8UF+CU9J4VI4kZzWVGTvmRc82Fjj144oTAzBmzPqj6ox1FqOa37cNWQw8
VV6GXSdXPtHLRCkY46RaWIOCQpBdsV5is5Tj8WqfSKkP6QhxLvK/dNPO08L4BZtk
uzMxXOzH9hv7yxoirHOkncU00dyu6lK/KINqCypFHZidgZ8T/cTpqwjdpqoMNs/A
qO/OS3TA1HjmH9HUfwtA41OLdIG0f7Va+IEUNQRAxzuVS7+k38j0WenmHPOaRArf
6S0KWGv+VwA5jHZf1+C3gKFNxd9iTTmqpisrbmtCWCa9Ht/yTfWywWnWbhCr8QaD
GRjSWALrhNJN+8dQgTmkXmQl7S4mD6dcoAURAa/70lPdpEbQgwWeZ1LnVonbPIe9
tWNnlmopV2A6m1bjMZYNNov3nhzaZ5jX5PACRWZdKLiCxyYiEW4PHRJs4vzL0WCh
s4Qi0Qf2eShCIsugxIJcjTHE0kjGrcE3q+ysO5rMwjY5IFfzOjEkwolk4ucRJ50m
0f6ObjFzWO6oBK9JcDyotesv7+OSD047VaJhC1CBevJVt+niQj0tTJq3qgXbUS1K
1Rw6V3+m3yLCA9msilH2Q+uXADI2T0f+Rodox5MRW1TAKuIsgdvUaYWmv3BBth6Z
VGeLI24/Me2Bs0c7Bf5hZqzAmurEoD+gGSFh1WKQU0jyPpm7ei5NvXru93VOPh8S
fTT0XNgpWbQ0U5XaxYd0wuT6Tuhpyraaiip2ZB7M19Xyw1ihe8cSd//zU+SZY8o6
PMcqioQ62UA52H36ltCSq7edT3ovKzSygVxbE1JyIuNmTZKN6djx9S4/ShYbp6+3
Y3wBdbw1IFBybuLIv3oPr/tqiLEtRDDD4Qiy4ekConYYYBq4lcZQ+X5Whm+BdKjt
Lx1+oSx5PZne2ndeIul4s77pCmhiMUx4br/Qqnx4I00GQyRTgB4V46ScXCROFj/x
FXlyoeLKR310JDjoietRXYPRsn0S06d897V+xSUjDo3BZEVr6cpADRTlGbIsDOPr
i7+VVBHGYmSWJSTRAyhGobwMSn6sbuuUGoAssNo+AvU5oxmJ9BrCngTX2g0rRIFa
xmTW8rzX08Mz9rCs73Jf6l7Bds1kBGMr+QgtNDOWc1Jidxu2XiW6zNS8gtqH6tiI
X1FYgmCuaNkOm0OgU2DtRjLdGe+IZoqZ61aKtu4jnTs/bSDS2PM2yzgYXr/+bx0L
Gg/h450KRg1dq1I9vnwQo7JvvzwyTvvVVdAo0NtXdddOdz8qTDKZIr1JBNhit0Tc
FFqogYe36U/iQ/+QfUBGTie8AZ1lGTK7ol+kc2gF6wXSBlYNOl1tbRLK5l7/T5MS
0wIYxZmBwrCBybufqQ5rXHJreJGdCJqy13Tqeh8oCOi45kDqhjE8O0lFdW5C7W9v
1ro5578a5NoaUOrynMIAB0hYubYhcJJ4PH2iK9p6019B9LePRKKG+3yU7DnlWN5M
tBgHbT6Xz6zjTi/G+i2Rvt6FEIMfE7QualD/BDdmk6cR2zb6YPj976eM56f9CKwh
kd3vcGeoJITkR9rfl7d06zzS3HqERC9+3OqapguhGPsUm0Tna96KdmfbGtueH5Pq
xDVjWN15q9iQLw81JHqDNiFsfxq1+AiMEgyG5wU6nDOsH+UdlRyqUAONy2R2WDMy
bv1pIsDHYwsNINpeC9WxD3Gd9UsBPI6KXxVQ92USfsxB87O2HvTK7HGS1CveGmJ4
XGNgUfVH+BI17g4BoA1vuNw/ddtX7jP6J2wzdPynnQQtWzUyQzYlS/5NmsVfJBi6
9bjkI22xfVRVg3EVEZ9fd0+IQeIl/pGtDJPo1TPtIG9WIuWSYlwMaW6neMfJdkSz
D9Mdc2mV0xssmA+3nH7uOsICZh/r9gZq9oMcALFxw4i3wP7c7AtEt0VDOVAWVygP
ctQki7BhealHqdIFja1s5XO9HOhN/7eFnSaGOTikjJM+YveDxDTenLjIMS9W6eCO
HHnmEDnfMj43ocdEbuMLcIV9MCm1BVu9XDg9yh7OYvBT0KLmP1DAKnSwWEqQ32J7
JWT3AwdNo/bJvFd9vDEhssue+Vsw1EQJZur+0N2JxVYbOU4PfcdivzpzMJiRale6
w2+i/Viip3BEMW8aEZyQwZBk9BX/9O2FKFXiVvPXsIZXc7lx0knhzF6qe0DqCCsJ
pI8404WgVECbs/EXW7ISeKWp04f+ZPSLvAmf5un3pcVrx/hNnqoRsK5gQBhmm6pL
mpXvFocB/lEl7Dk4RhMMQfNjVNP5VpV66Fo6x0sN6LZB7ePrVzxSmLkInnTkLSL0
ovkmJQgKq+gLu9Hiuwr1qrc28hZELaqxkfaSFU/VWBVopsn6c1pJkymol5vhgrE8
/Pm9AO8jgbhFNZjVdu3K+ZJLPC5YRvLj3IvAzKPPO+cf4FmwbUaIpdKqr1W65AN5
Y8Ra07Z/1kWDvtE4WNtJOM4/CkTNKE8974PgLrHRFxtB2wPYkspwtOZQ3UASfH/n
sYRCj8biTsG42tR8U+YfL0XeJgpI5BCtwYCJ4ioXlaTfz8smb+l7c5gIBRbPpj7Z
bTnrVynbmfEsx028AutpO0eKbFRPKn3qTWOQU48zZwetj36b10x+35NTr5lwLSsi
rEu/JHfO3aoetcpBT597epzRS2OdvJH2aTF0R7B77oS/FpDx4W95nkpCiMgJqDhG
T/xkGRXuyL/KjqjUcYUR9F8YZHbkYvlC4NQiVi8D1JXAAV27mQR6CqNbkQ02fbJx
kfiRrGUj1GDNye1lk1gPND4qInnyy9t9ydGvz1QFlgiO5/4QRE844PP96fzhb+xf
8Qskm3WdpjMxAgcKaiHyhbt0FMF/AyGlEMFjSIxUwrBrvqpHL9cEvpQFDLHaGyis
srFnGQy98tiYh0Kk/aeL7PID84vi04wl70s//ez+JS7xSF7kqyYYaTFRgF9vyj80
PC8EV2IrXdh3Q2tBjGVpt0FXYgxKfqUSN67EwgJyvaOT+oNauOqraU/ZT2X8w4Ux
078N32mrv5xUAavlIPe+3LRjxzWY0AbuWcu2czGX973JmRacGJ1rvE9de9py6lA0
4IrSHyF+dcSILXg6lA/ARwy7VaGqCF1UGaZ/ZWfIxtLPK2gkYu5GqpDbCVljvGi2
hJ/UXDhNZKyJck0vQ7E4foFKN/VMl0sg+9hYJfe9ntnm8CUSnIItcGAyYjK2hRPk
FTCcsF61OlYiEsZ/pbCER4cIgG+UkYsUpVwxccDI6KncKILMCocXVVVuVrxzm7bg
Su7NNzBz7iUiuxDbv7c6P/AIdxDhrXUpl+/kh5JA7KAWaOIRRIWGj4qcOROjMtr4
u1808alcSmsxmS9+U1rbrJQr6MeY0tKXNOmch4HiZCHrY0QwCCSXHjQxiC6rAHzS
VTE573wJ80OuqGDeZa0bkD8BozFrDh9kDEfzl964H5iFyUE2knqTAdES3QRCC5fe
5svJFwh+De6CHcxy5Fd1rOpViMSRq3Ozx3KzrmFWpjTfLs0bqpyN4tF/wwdq2SxX
vJXfT+kCoElXpgN/6QIxQTC952ytka2sU7T8GTnkCLu14spC+uiJlh2SSmPX4z/A
IEh78VRpmyhzslwyoooEuyB22gNi80WEvkq1dYk5p2RV9yLmJWGbT0SjC/IYHF49
x8jvz3Y7H7AQJNUEEO+YkUUWsCkXqp1Hg66yUcaYXRhsWN4EbQS5pCyjorz/i2OV
Szf/8X6vN8k30KvzqPT0x+Y12cb6pjTKJGbxEiZDbQHpP9eS2Mx6TV1CqPNd7Qai
Ew0tFC7NKdlz+p6Li/XfYmNr1DoH37V9pUk0aYh6rUWyIWu75Vw87FTMopsg3W7U
i8/T9KUZr3wO41+NeYrndTksFizuKtNmg+WXT4XfA22xLZ6Ncl4ZoMNcmuClQwyI
CzlcuVhZCW87gMKYSiHDrgzcoBqX9qMTps9sJUjScC90DWcc5U/64XzWXHqqcbii
Vo3QWMbFuUHgtiMCr7PeDevR5CBrGGprRdJ+kAENN0NPjh+bZKEOeMpQlelxu0PY
9ElXVibojh47jLgqyQMyHLmAWThSxPGdJ8R3ZZ6KNASN1UirbDL5CWKslDUkkp2D
6os4ZzhYCvPhUxcdWS8NvuIMWivAMQeGLalFRu5Znyqp2a82KoH6bybQsEHxbmhD
Wn72iXLHnEXDEGeck2ODzRiPPFFFVGf74l2iw+RkkZIyUjT7Nc3aKaYupg4bvgkf
dNBmILUyTbR7VFCiSbxEpEgrBwzHnVWQArAU0A71Hdfi/LgCwtI6DLDMCPOYIpBi
acDJtEb9VPrvaEddfwfIRU0SREMkzlrTAEH87gVQr+fEcv3cc5OEUbZxMLmNIwJc
pBpPfUyj6elTBW2sPiziGPcPqOs447qoXdXtbqfTW9h0vMrOhGzAa43G1wT6NxNg
1uoV9bP22RRui3idzLWe/VMO5yj1KEx+97xZaQa4RgFoP0DP+OtSBe5vEsNfgfM3
fjw7xbB8/t4HH9rwRqJGrKId9c2yldsqhGtR5qwNDVY3lIJuidSB6EXPVNL2Vjmm
ThSHy0vkGOUmqiZro4SlJcYGmfdmJrXAevHe7V8BcCcQX+MO6fz5r87LBDeAgS1e
7q5DWEw0z3U5MU2GEKtEOMj9C95GIPMoz9MOCMiHWQHYrLYSoUpODAe8PoqXofBC
U6+L7kPwLpdvv1q3ukx4MKCDIHxbHXUM3qs+88cQAfKpq4opgHch3nXdab5gyZh0
+gsc5adOEFLtweMBg2QI9tKKrbIPi84K5l31tHveQLuuGvNKT2JQ/3yU7AzYcUmV
xkIDAJXFHEU4724ioPV9VT2do2efhAe7wlABKdOnUK+vLYXE7Ve9zccZ6rGlBLJo
5ctr0i2nObB21KQ+l6j+N4ZXN3lEEN/KNudSil4mpPqSBKqw1gfyVNgNzHkxWdwv
H2iFqoebUVEMYF7sak6GjOuR/fugnkrP7/E+dJish+cQIE9G8YqTuSBmDik6LXGT
1iRnjvP9ttq9ef6oCwH0ae0oWXfx/jS0g2IIwY91jipdV69R33gYl7CjSf8E2uS8
kbDNxlFxwFcXiInZndL/fPcF8QBEzSnLKGJ1ybJ82WtsH0z4j6msNrXOJ+Q+Blg5
SIBH0sw0Xo71BLq2DgRL0lq0ycWu0K42EiUaPYm5aBmx5OcjO0Ta3V4D1UgrBP5u
3qFUtR8eHVs7E6pglVXmjEGDj7cqdLCETVCB7yIMxHSR5liXFy0lDbxMD0jiddT2
2T3Dp273mjcVFT23yxZisHSQ5B8f/HgJFV8jpkw5ZivfUx8ZyWle3H/5Pdl2SNtK
9d/YWaorcE/XAsDBn5e9fswjREulzOdJHYwQ8U5LOPIfUmG83OcV/NjW4Q14ZqDd
4P0hBhe9pQNRR15S4A5ZZ6ZvxscpnOaCSzC5iav2SHL1qXmSVaxaobihIoSIr0rF
vyTZyeaz2ut73AgRwI5JglbOAeTSmJS1zApDjdn02QI4R4D9Zc5vDi2+yE0oVGmf
PxyZ6BE2CUkL2O5WFQHCSo420+j90gkDNpmXZu7USCWxhbYc2EOnsPIUjK4AUGvX
f9TW0MqN817CjzHeeDrPX3TAJ7bqUASrOb5b7Q6oYMTGDdD1JVs8QUOn/GQkK+lS
YZYlAiT4LTURxMwS87NZgoxenV8RuYta4ZlA/U7lz50l/2+WiQH9yjfl9sFevTN4
mE3Si52e7cbNsaRQzERAd543nshSmxLGOVWHPNs9P1G3Y9rJjuVMRAQUpLpgw3a+
VJyO7SveQ7Lttc81va38iva9tXT5xxfwARcE//+8/SPpznNFIRCrlEzNIZ22zpvp
C5a2QsnfAqeeeYC6zvwz0nvLaRfaejgCWbD+IGxaXOsKFdynCOKxrHYcz1CctFp3
5bghid8rDElv5So1aava2Q5CKkl3bhS+nC/sS/uFXKmvu6T/Myigr7p2RR6IC6Kr
ZAdP601Grsk0gFfvtz7uOAJ0v3CyXffq1HdMVwg6lKNxevSUAtzKarlazP4BOXlq
LIdKOrp50kCwBJA2kewHvPyliNrTBKNwfuF5sNK71/KUcxohkRFRerJeR8NaZw3U
iIh9RTZsUj2IEEkYWJ4rIQiaUXUD9ELETugwyZuqV9/Lx07N5alr6gUcXgVq9Sxg
ODRBYUsKNwFlxratujjXRI078DMv5aD8MbV60N2a5hmYdYsC00PmxoWpb5DhW2sH
tgoWM2jeopIs/F7794fKdKloRhPjJmq5fJZeinrXSVITREXQ5VkM0ebqM5EjSXLg
sRu/SuBSI59Bc1vpaVpGNtgy/qMitzm1ZHiYJ2OcxVdTh8oZ+zhMTK29LslOeTzf
nrwdBFjW3hOeihtaEF5v0po20e03VnCJEUHgyYC1q1wBWBTSe9O47DqMoe26sc2V
SAkckBhLuEn2pzz6mI8CQXrErpWssy3S1cVupVwkcte/7VFVuSs3rOHtdd4VQVD3
7/cRgLQBJNEHlRSOB5K1U/gIny7CXy4QZ5Apk6zfOgs7UuJY5y6fw7WstgrHRHd5
fLoaUrfB/qT7W2+7Dmir3mOlWxURoo7/QcYPQMieBsPAGt7NEAsWk4DlbV7YtW8L
hw4I2VL5IR14XwbO3r+phyrQMbtAxUCdFvLBxvHzSvNYcxdRc2368/OwROw6o0tR
1Q8+U8vKYubiuTP8uGXIbzLfKqUti/8MLlAPObAcwQzlM40WouYaiLyiTCvmxDOL
dVdQi5Q0Ap0JZ9FJUyoHV/Wo6BuEbXdlkcJBjl9YaweZgBI08fT8U8umJRxP62Xb
bFQLuptb3/MbRdE52rfoDfUYAvT08f7fwlvUB0Lbpfdz8uuy6hZAjx33lo6AaAS9
y9Jq+V8qOYzaDggctHFE/C0dHc7N1nJ8sMnaZbIWtIfv73qB5Oqr8Kbf4ebQNBBx
v4IZ/QDL8iIuOKy/XynpD1CJ45E8TBzHld+oKZcOSFA07IkWBS/kjTF7ghmVWr2P
S/gm7FaX6THRF+e6QAP1PuTtEOraCqHy7iX9edHXhlrbjofztauBdIxrEgz0VSs/
O9PA9r/Ui2p+7p/E3C+5zduLZsmlv+xvfWFgQsoFwA1AXYgBZXqOJ6yFZla0Oi3J
jXlLR9BWFnNhUBXlW6KzTB35ta3r0rWgq2ybOeKu997zoov+6gNS/q6aj4UrYzwd
cdESJtvMHv6LFzhjNtt/1bEEVcDBbPOGaCZPTpR39VxASZqr0fhxwpIMue25yzKQ
1dMqGPl0b3r4fNYlYfa6yyymkXE4Ncd77Lfoe9eOnFKGtd5uS4U1nNcgACh2Ejw6
EOf4L5ABd9zu9TpkBIjBgs4e9fp9LqNrYv5n7LwCPaJFvbnj1jIUE90dJK8U4VMr
cQ+K08WtJmnN61UYA0XfyYy+q8uIW7AWxhf+5q2GsIvRj1kO4RErRKidmJIORQSl
gIqsNA6JkbL4esjwNBpd64oc28pIw8AJM9HsQk8GOa+uBTV0Cl1SiJWfWVDUj9i3
6LMi/DVKA6ka63NTKRQ4crNJ+CgqPbvNcZm2dQmQXxEkQavc88RIQlwXDElnz6wL
YJgmBXKLqZqN9VZfPR19+HKvAHx1+PQZmZfYUug3rFfYBdNPYf7sSFavoQLJVhjR
DW2ZzVrzYwDo/OtTAxwhYIw+Jc1eaA37qtjlmXkDm118vvPDxSP0jW67yWxxjJmu
1WX93AwzufexbVREJaEvy49cjh4AtJzeZFBb7ZXHudXshHxmdkh7YyNmMN1BQEvz
qTvv/pdtn0Dqrk1tShlvRQeobNlTBMNzdCWKcXS/aeBo2ir0zbI0KwObDPjE+82f
MGJNRy/V49t5ADgZDg6JF3xrPYGnamkiGz+oLpnbq5xs/00DA9GkfoPW+FUknCaZ
+kFCpcNx0idI9y17mKpC6tNhVIhQ4qio8zfzMqH/enQZBKVy7UEKlnFKrkueg3xo
VAfce3vbBxEr3wyiduNAMKEGfKEW07t1ho3099vY+vxFiu/b/vDU1x92ZhKxk+rZ
TTJXZPTcp84WXqcgHyky8eCMxYSVkfWOyZ+WFbCDnsPg4Ria+rYy1MiLhZJWzBVw
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
guI5KdUq9VFCpZc9kXtw1Uw30PFRENV0Qgdmsn1vro5XuTumedviCk1DkeEx6Yx7
1XrtNGU6Lw3tAHm/s/xWYELzBkdVlwxG6qH8icpBvkJ0RqslYwG2Y6jtxvEUpCHN
8elsPLcjO6VwByAdjehUpxw60MrYIcN6WEkgT7DJ/3XrNjWK3d1XKJgxh/SYRgKC
94REZOWXNlFknRJl+gAt4CfM6BnTsJ3e43D954RmUd8Nbr6P/Igu5OhgcKLAuSIO
dxDpqzDCj/VmK3ghP5uUKCblZiSmjdsqU2pXZm/oJcB3uUzgHs0rmTc5A+/qQmFs
o+g2wyojE+N+5cROGDLcdg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4768 )
`pragma protect data_block
RY+ZvQxIdXG9sHCd8h2S5mJedcy0S/4XwTe7xYIpRdE6KgJ4uUNqDv6x5aQseJ5i
TvPEG3Z9iX3P0NqMNDeeVhUivYx3G5+i5R1tr3VxUAoz0irRPSqoTtYiZ60u6UyX
4Kb75v+0t5NUkWeXJffdHBMQwwkvGZAR28rNi1M0D2SiFTLUp7uugREIXJmjcM9w
l8T+qIux+DmjsnMeTgvFVBd6g3e7TKQZv39MSAd60RFBV62jGRIMJM8eqE+K2nRb
VG6IQVr/PykODFtns3JKeiFaoxAxMoEfCuWLBoMNyOyVoxdb+LmEVcm+wo8eXcEo
l9bzX6fxVhavpk5+kKqFf/QQopw/QZfW9X1+JFHK/3M5b6umESt7FF3WxnBihoyA
euzqkIUWGaqk9E9QgTWYZ98UNfqLzXmg2UJPAhHDjQigbofrG/l21x0keTUXZCat
rSxK2d3ru4SPFXqSbKd23rdeNKF3SjhxG2Ct0fVREJPDpg/teBEhZz9O1tUdUeM5
Gwed2M3QcblaIEqrTZOiYmFI807k8HRjs2hANedVm8puhaTG6t17VhD5lGT84VIb
U/Cy9A4V8+cV/YgbRUs52OVJDW7ASFNosBnBJWJHo8x1i5B6m6OYUnBl/ZqkSB8z
HrR9SdVvzmxHC+GH7PQj01Qwrlu5U5KcoXwAquzJQGRo6BeTs+TbhU8KcCu6TZ0x
qgGcqXOp4+XbtOtFQUUWBDr12SQ/a+8rBF/u5oRwF3tPm4/UKMlzNQ/VbP/4oAXr
KiNDD4KwLXkYQtl191vFvOvF+Yyty52t9ge3tfhE1fa7+m7XmBltX/WLXztss/4f
/J1VdAZcXFRbq60m4llXdozc4GLuV9fUNrbsil3f8zd8u3vD0O2O5dq81Z4IqBnq
2y4ytOIBbzJDfJnSbCzk7dCusdH7vOhLuIvn0fOwphfc+HF1PGhoHVQgy2f+J/8M
+KLL+yCEGg1QgBghUJaHRQebPMG8oNdLg+3FZhnCmh3JJDY6J9yPiD1OuS4IrsI3
mZkpf7l+dsihp6y+8XduzkEuRrEuDvi2befMLtLNkj9cGVWT/+HSPGS3Wb9+ajcl
dN7TTeiyhmxRRvSREUZSrdErkFlYroXUd6QiKOBJnNlrfT5jgYmnkwblY2/z+WR+
15aIzZBo51rV9jbUvbv0F/Jufa/HpWGnDsgulExQ6OiOvxfWBmfQwhg5ADXc2QCC
jliySWL+2wtWuzYHiI/W1m8FllDIUQ8Uu1N6K2Wxp75cjFznUCNbRzv92QOv3r4L
yp8+rAiDJKiXf5HERHPh+sNArGiATdTibgMdvzCcl9zCedyb2vZo1LmMMW5uu+7q
a80C8aYyXQyXg/G2sxncz1ZADtVEp/PNnkgasqP8xX+ljpYEncagC85eGslDD7YV
LcljH2y3QES/uhg6hO7+4ceSQbPaXRP858uc6MNbhqx1jnaLRSnlHeVBRtS2WBvs
B7s6LqqueZZ/Sxtp0/4N14iWtVPlbfPLfW/4vPIyxOlmEujzbVEeDsjgJUb2C7/u
zWdLOhsdpa2f+WQMUyiDLo2yWFnL1cCtWnpxJfSTnwvotU2Ii+WvFmQr7x7Vr6fY
jNgq7A9xx3qwVsVvg5k/CINQ4hwMAg8LZBSsbf6wsaZXlYQZDrrup4YhwThi8JBG
chE8HqQiX1N4bQdFFYkj9x4i35cO8QdWIQkyEaHXUC1tKIqe4akOOYpcXusl2gEg
xjj9SGqew/gu6ujdabr11LSq1H5wwNb1+YaLiZIHZ6aevM5lRs1yDgglgRrfi6kq
mjG26oucluRUWKOJzlK74CujIy0miq6ZnyixzQmUVFt0wjOFVVdgyk1jaNxc3Ng7
Jldmvij/bvG7P2McqBBn1yedzw26xjCeLXOB5CHn4UMiVWxq/m0kmEPO5ziOBqLp
4sH3IqnHdC3eo5e+o2WywD8IcR/m2K9D2jrs5ovZm7BRu6qc+Naz8c+Vv1nD8FW0
zR6Rfgw4epGYlc7Ni6lBHcVYPJlpAS2UxUcb2t468ZozdKe0DLmuQZDlNkvf1OHz
b+jU1LuztR/rGfSztlIah0wIf2RF6b1LYyDxyRzcvwUArtUeJSHyxXQdP1BzMId3
Xndu92fV/5pFyW2kOyQ5siYg4Hven8pk7OI0QqvllfV7ECDQKTv0PyT3vaWQ6LmT
z+NAeqQKsWBIRj84j+xNVLjDGAQyiRl4Kh86c/NRUzaon9fd1e6dDk9PuttMXsEG
I1LiNQcy9fD8Lor1+aqsfMy9WMa6Rlz47xBCFeIAh/CF8Qry7BUB1zgSO4/UCB8Q
xJtkcvMCAlSxJ7u+JRvedhXM+80sIah3RaFO3poIJb3EEt6gfGMQlA897t9qj5dw
nI3BisR4YCEYO4QL+2eZMdMF9qdnPYkETu+wSszPn5EmuaLdyS/CtyBP9UCmulzD
ABeE4y/rNWTheGREyd1hKQhgZE4YuDORmLpbBCEK8w5RL/0tx3Yd7HoajpB57G2w
6D8D+tEv+Guzf0MNlgdycA1wX8tTgaKOBKJPX7DUItQsFhl3nwhi70i+I1GJr1F5
CAu0TCwOosKcHnun3Aj2Sx9uBl2B/2FB8m5ccdSES/02sH7vjLAa+FIE/yEZfwvP
gO3H9YfcGAi2j2HwE12N0BdbpP++cf2WUksZFbArAe39EQKRNvzL7lvS25yYRgGG
2RjUIXzxubFwVtUX4jnXfahZMCZuHAoBDvaigcUYBLBrzAYgMEFcR5iRKUujmP1m
KEipb/SerXpCSLppcm3yYhEnAt1nZmgwfw3vgTeL3tbvQQEn3Cg5nMN7OEPjX/2F
QdrYDdkksLeWZI0zi/QnpFsJCaKWLfBDX6//r6z/OrOiW26ax9QuFRX4Sb/iMjFf
2u+U1rOJsddalWBEKhfRG6PUiQU1nmvZUPALimN2sJB0Z+8pKqkiDKc8y4G0Gu5n
q9+TwKugrFLfL7YZpa0OZDrzEmFMSbKCHRRn0MFFu/YaOKH8Bt7p3bTbkWAbPYeR
nl/QJzqzcf6NEzZiN2v8QoIIjaX7LigFSyM9Mfv3LYtV4Y0tM5sEfljd2WIZqc1n
YKsqMPBjf3/qJ6pW9RrzaLUcyWY5KC9dCIrRIV8yQgzGk2kfkFsDaJnPtAwuzGIC
9FlJmDm2cLmXz+T3gmWMLwxfG6O8Soo1p8Bhy6KlqtWiQehdK/6Z4CGsNCC5Bfxf
PR2S7/TW9CKnzIdW7QSLzypmd09u76DyVqVoBfQddAEE06PLE8gvTWMG2272U6D4
NnlJzi2aNMoSZPVgKulz4/qWQbR/eKZ7xxosawioBbRJSkPJoFQjYbThxkAuTeX5
yn5j4XSGYmwQmwECxWlQhavYfIdv7XlAIbUVkxeUiDB91j8dppokUeCFMr7EaqIP
/aP8AVh5CEROcpuMQIVxXD1ja5XsC1QC9ca2jlKTLZhMIvqfjFQ4k1h8QDjFsvs8
o/ZCLlFkeTwVJqht7KUtgiSkNTV90GWW8KVcHyWkJroCywKUA1Yva/4QjFnskLta
oZR8x/tpeZksZFMGorYbaMgJ6T4lJfTJjgOLgDxOtvcZmqfojjS9Di2Ph4ScW35d
3jq50k7y9QglDnEk9E9Ypk0GS/XVftorhmcGCOjLtsV7FfTEs2ecf0HcJKfVMzyq
yo5GThEOD6bHtpPeWn0j3bCHmSD7VyjcWgd5HnACKDLXUYqx/M7tCwkckkzAOT+F
o+4kPlnNGfW27XFteyUz171wGAXWmEP07zxfgX/grRQ0yQVhoO1MluWEb7ti7CQm
PNuCPEHH6kc+F/+JTHMXC1dmJhcoGOk/bQei8bH7BM7KJAicej8kIzhjOqaGwEv6
+gv3JoYqUlYzX6cAgL6WQBSiEO7d78gjnJlNE7beIBmYmmkMT6cNQ7OhaoAIApg9
iCPTCPf8/7xRxh448oraUgJm4YFYmwZBWiylENg86/c2bJULIFOkezTkmcR9gz8J
oqWuVi8wsa6DT2geWovr50LctlnHBEYF3b3/pwAqJ+c/9pmeKM1HZ9lE5kYEtTNl
nH0ew0floYMznJq3sS8G7OKReNWWezrfLFLT9k37os9jZUMkzcElX+ewfPlBr/8e
VK7CCAICFFuM3mm/eGQftB/5RBM7ZrcCkxFFid2/r4dzmHFuj8zuUvb4u5/wSsa/
vsunMb8hApwB1jqNCmv+C7Vktp29YqO13rx7Q9JBTpg0WX3kGsMb78EpQdonPWzx
VIZtW004jFDKZPNxlCrBjY/3OIaAYqjcufMKnTASgLLUfYEG24qWICJPKpBgM+rV
6eh0FIMvXMO6k+/hh8tILl7tiE/hyr4SEvXRLJ0Y63Wc/CccNayHbKxRqxr0lHIE
k5vfTVsp7Hg2jaEt5+UlW2v4SVQTKBf7w+ot8gVsbQWXbHEl38sG0Mvh+FiE8dch
2yZ7LiUoztvfpLq5mPe/aErZVqvAQ1lc9jw60Us5DLeMcK8fDYjkTsOhFGErh9/0
g8+cUpfjpiuGMjN728x8oFYkn8wbxoeQlslwB3wIKIN2xs93CkAhsNlJloicSp2D
tovE4fz5NXV+r2fsRxEWaD1VZU3koMxtNaASHxcWKmWjgsF/jzBcOolkwFyjbKLP
g42CAXUvtocTPUZoXGqa2DEnGOK8f0eEcbsXdWzSicU6Wze78DLllrLAll0yiqbJ
3ElFbPdkIhoYz23X9NHTmMC0e5pZkA/pAIzMLQxUGu2tcdsNrghqUKOmV6kEjmMm
TLPBvSIK5DGOXmO9dLTTYHvrRN8AXqBB3T0TCR027RKRhDsBalAb/S6Waotb3jkX
W4g0/ozqG5PTpMuqnyfG/Z9NYg1Ap7vMjLfAxWG6B8E0lU5ERTXbPFiAkaZ+ALky
j1GR5ve4aNP3DMZMJ65TTI/lLrU/BiQiTM3ymihBo14n8Ae8OGtWIg4u1gZXNMan
igxrwezCGxienjM4INFnpqr2rJY22ZBaN+G3noISuOr1t/rzFkXh18/MWibrwNNR
hrGVN0QQCICKLyVyx8cXPG4VccrFC7s3Vt/AbPLDCSBOeXxE/vZatF73nF/SwuD4
eMEKegcLrvWBT0iTrRDlEz3eDIhmfPcKr9EQCwURq8h0iveeG5PBd4TUq7pn8Pqf
BIl1G+X2MxnBjpH/4dpCzSArnmiSG+51SiHWMztEZE2Q5fAjCDT9ZrF8dR0kuv08
bXe3Itc1MmcPKF32yKfOjkV1gqHBPE1RWjBJrCY4y1nkFYt+W6MLUbwRWJwfHS0n
bw/F6O1uMd1c15X6+svYV77sFtcjTHp5jbNDlSzkcUlSPkpS7OLuDkUFvxUlCKtZ
Q2ZfOUX6mMYw7oAFENS75q7j7lTODaiIaJAuyXKaR0p0NfNLHsA7kjBhYfUgDwZF
0cpOfFrO3xEM5PoQiHEe1qdun2xBrofqhQRHnbGVWZ5midLstm+W0mNXIEIm7Ed8
LX1mo30fsJSsHRneff1Sru5g4+0hwFP2Bi4YzQu/yb6wb6MbDqzmCG7wBRSQAdik
FUhIsqt3zDLXieJAOHxYsqdWIEy1wMOaKZV6ihWxiEbNApicywXtJ2FnxQ+kIcru
SJzmw3bAcFM7ppjUY12Wdb68B7Gurm9Cc1C9OY0rIk9WxcQBHwnrCP9RsRaR9Enl
yOxU9fz2AFz3u9EbSX13DUSV+Z6Rv+HOikpps4IeMcxr0Nq/df2EI8pro7QSjU0Z
Ist/cNtCJKzQ1ayYID9H4AMYq0iUramDERWcLJqd/1jkqqSVzowCNZ95abYxSjJE
NEIKnKpGPQf2L7euH9JvyO+j4aKi8Z+TMSuToW5cPYyUPNv7iwflZQpoWG8zt4yX
it2V8MWtlbze2HjvjAkl5WAxcKidxG/Edqz5GCieYTJnhutV+d+pDlo595rgb1KW
gbI7KyFFPOYk9KnDJt255lD6pJTCxRpps+EpyiZwpwz+NKSgS3ZKciXogg9gDD9g
mZAYVNq8qtmAWU74zkhmpUdMcOzJgqeSzwgXF1S+3ArJ7lvX/EnS6jwAtfs6DEdT
P85EpMYp0yXCWoXLV6Q+XYLDAe4ozR/DWsbibjdmkErAxflNGkbO77p9MYTLAG+I
cjLEpyo4vQGnOEndHT40nQCxYBWBaFLzSAi0SErMP0TWnzi1Cyep3tekqYhOKl/s
2jJWCaH2TshHrEMC2dRiPciPYnsPgq5l2Fjvu3WGeMnDRXhiQKWAVwNNRDNRwPmR
VX/dtVzsMs3PGVAK8fmDBTnWyHwORr+FmP9OunEEJqFCsy8txR2Q3Oq4K9Kwj5CY
DFO52mr9URvypBCoNo6BUAMUCihMK51G51uPoCouONW4KgYbEcOmZYLNCH2WItyM
/dP7wflge6856xG99Pf8bg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jWB6dZW6ajyjUvFhpXknGWdKwGqRa3lWQ8OwWW3d20DBU7I5eEi5JtqU9hRh9sR4
MkTKUjxc93IbFGrW8J19lRUZHNwD8OblLRtCaD8NVJbvqcbHGKB3BI01g6Jfd84k
MPf3e8numSl9X29ETyt3nE5jjcYUVsovp/CdejTujjAYMP57An5aA/YacNerlmgM
K6fC8JHQQZc3HuCnBt21+SCd/aFLbFv+4gdnfiiHaL6FPzsApuo3GnyKidehlStJ
LzHhQZZoi3qS+A/sTMDKcXT8Hp+3rBT4vvnWgY1KKw+m/3GmKU70u3vbNIVkf7e3
Y9QRtxo+hd/ZGq1c69cngg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8720 )
`pragma protect data_block
PYDvmDGGM/JDBATL5/N2jZweHmYst8txInVneSGCzQ8f5zdOKxl+kRUus+WffhhU
aY4dApYC/eBzYuwcJazkbz09BuOIlQRM4cymII24LRE4VVb6d2JUqul2XSRBiq77
7jTJ2H8j9FErhe0t33DzhbJjsgi+GalbiEMXc5RHD7YA811Nen1nnkJD1UslqUo7
nCBoXQJ5Y3CwfQ/l/n6/4he96WrzPmjjG4HC2AzNsE8rxLOkipbm6Gr2H/QNCNp9
uXbN3VBO+HDHfABzj9zfojdePDG1Mz8mbJM6QvzNXC0xE/4pXJ9p8HNiYmS/OaaB
kWXf04eI3lYB9VLcZo8yNxfclZ6ZStAVWUpXUQIYPfs36ziT2dvORElCOzxeXoSB
fl5YguYBrZtsDbZa4mUtmNc1hkQJNYj85OVtyYl6uHJ2VFBfVLcHoU4jYm8qbxSh
86g0M3XDuWMh7ZthjAx1RCkcEYdDbQS4S73TRIycpoZyFRm9wuuMCU4rDk4UraZi
SR12CYYbqDd9OIIw/tYbxku8m8OCXkodwVheGV76Narw+ev91LJETdu+W5tZdj7X
zYAzewZjFZx9ZICpieTCmObzltMNiTFRmnaMKY0+HPnzZh5QnqtFvun6R8vEAbnK
3QF+bcQFOkjNwEShZCY90yeIoIGlcUCY4RaJs64ibf0w3tUoAS2CJVP3c/vxvSt+
tAVTrYd1hw0YTnHuOhIYoC+95XQVslDCPiurhTIKhkkmYHrZLkRHDL1oflu1m+/C
7TnC4UvvHAjvrVhqvPbIHK/5cdLHfGq2ROKuIDfVSlsleIkJSQKwqZEzrgLWuyva
/bIPFVV1UT8W6AB2txCcK5v9H1MooPAAv3/Kf7c0tQRWroIrw5E7dR3e9dedldzZ
6F2F78ykj1g1PgxsZAQaJmv6Ebn3q9JOjkcj3sHDx9M+W/uh5y9iSMYQlUtH2jRe
yNk20riRsXvd0VR4HpT1UjSFpFXrNBuyo53dLiS48X3dL1cyakJuUHwm6GEOxM6E
XUj19PNrqMc4bQIt2nGaP4jMQukDjwY6Yy6mHvhVLpxYe7O6sgfgZwszj5b53pRh
9GX2PkzOr0r41QB24wPFCcPAuI3PoDoGEEss9K4CDt0QbBYxfIM5nMF+NiY/As9a
65HTesACWav6B4/n4QwTno6IcnbBc7tZTdsQieMaTHES2g/eR+4wQO8j5x1lFT6q
l608Id2qEQ2YURAp47EhtWiO4jjBFaJq8L1uiWd9EkrDGRSLePrsoY9oFNma3+DP
6kpumDMYFTph3xyxK4bhOvd9MNV09blPU+LOEXnn4ZgTgdzT7K/HsFAmaHN8DK73
UC0xw8DEzijWI1NPw3IYTyn3Zt4WnzHp9pKKMA924kg87+UYrXFae9Zbcp1MyzEX
Hy6prKfWlCzngDKtifvCOl9ypU4JNoGwwZDRVPwFAUZSlFxhLClNp4VdC5f8HsyK
3RW8TIhZ47WN2aU33yD5afI4QoVbY7BsEBrAjwowRMVVySBmtXV6SJ/8KlD+F38Y
xdYLFk66MxG6AtuhFRPehGeUyagM+zNBaxnFsw3iFiUofWINALhwMm6y8o3GZR4N
Yn01LuTp43OzStVV3+qypFS8nmA3Rb3J65e94IFspGAA4f88kYG0iJUgcVRPztrb
PLOMIwlKFwLs/e41OdY3l8gjrQu+ODjj3QzLHB5p1sZKyK40YZifeJIGZFsyj95H
PosTemp0eMmasIPbo80A5XLODYvK/Y4PfWM039ifYvpixNB/7gFIs25n4mIX13ac
+IApL18dpRrZY89ujo9aNdFICAqjj54OBz4tXF0aeKBYK4czYVQjWhmE7OM6xuXX
T+xfXwufmpui8E8tIS02nc0M9HrUk+/DPg5hEJpjSYhkPJsQhfs+Kf2Efo3SRFX/
EU1aoVLlxDdaH2b+1yhQojytjTXpABr/36VdN36fz0wUTDAEyGCUvSm2rBEkb813
5TuHBUFx2OehsdqCmYHWXKizUGX9b6uRKVZ8C2cuCdA7vhFHOY73YFixprXTCNmF
FzKRQEF7JrJ1Xbaut+80OrhvqrXiDkdt0Wy0oDwXkLBF7H5sTTugE+qE6hLLVtU5
1aF9AMvvgrINd1f4Eila+NfxFfK8vO1leAF462tRnIYSVv8FafdzK6J37Czf2qCq
FNQ0bVh6oD/IeXnDpN5crqbsoOKzqYXh5ZGVqlYn23mNH+FUTM8k5NLg6qkMvRLr
E2ozvalPF/t4umDtPe3ERdSWHOxyTPSTzA+LqpmQo61+lp2EtkQcub766bxge1nF
mg5CHxTuXR4ZSTNzQ/mWRTUxLwPzheX6SivK6eP8ZD97sY4IEDIzYpsv2jnEjsy5
/ObtM34Dxtb9aSR0UGs9cHavePJIODSkcEN9O1GvZKyhGl0Tp13PBmP60Ok6DD4i
NTknUcoXHoc9AvKf6ubjqabvv9dF+M0FUzFCK/SobfAAARFJtFd7iq55rwvaHhWs
YcztOjwRODNvAWvzMAlpeBv312r/k2sTG6gQOrQtlFAIc0x0kJ/JgncrCntyraNj
9hEa4Zc6j4t3lGAZVyd9r3J5Rcl0XYUVQxsT556gVlSQu3ORNk4lT+Z/jQAVkcvR
g9cHS3FC2r56G7dUIdOMFuWldwMmbzOjxlYXCNBKb0FXgYeqncLDh8md+yAn4Df1
dIjdJFEqeZvj9YDg6VNdhIxUfKwQbBFJ/W5cjY6W24stkbr8hFPFWA5bM57K0Omc
0n3lIvG7cX4M9p8crcGCNEmaLy5jA5zdyV9Wz8eE3Ixk9WQeRA42KynZ2i3USdAW
AzGbW2SUD1PCylfAgOEeMY5DtLXgJ5wJe25EGYNwLD82WEsSfxy3MQBAWb0FzyRa
KbTct/RYtJ6vFLognuhAlyp3S31l8giKsTcyDWYEms6V0YrGW4EEGSxNavrXyvee
98UMD/ZUoQDzeQTQcRnhz4DCp9+awS61cN70JroO7etgtO7X36saQbiJ59ukoHny
i3riMU7D8e2C6vEQ7M6CKcx8L9wTQGkGy1JJUlMXrHg+tzzCTn29aOuHA8Uw1XeF
bVfGOF9SOYve8b5V51SN/YeEcWCNAiAU+w9qjiPBGbh4ExqhsKQygZotMnPJlLZq
wVYd4SJfMPBKyJImLkuCwP2FnnI/I9BtIjHIQGgpwUB+s6EYYsikVa3CY8FPY6BW
ft37m6zN4Nd8Kku/++HD78jxKz71EA6FyNgYFd/UN8vtp0WiiafFzcork1BRAko/
liEaJUAULlDcA3w8Zz5O97iZU2zlwL/8dN759RM6s+O56AJLEn/VFUZ1fjam+AcK
9APKxad4Gg13UuNeF4E2PnitABiJW7+VbMJ5cyR69dAOrwyqlCYXOonbdxuVpEVE
H4Bf6zru7GbMGg7xt2mX41ot40XMElmz1f7XYxLoge7RwX2TNMiVMvho0G5gFlxo
QXIeQuseW5rTtwoStjqHMVVkE5282oOw52K2BvnaojE583QA3YwSM/i0tZi2IDYB
nPF0H2QfwkUEQPL/P25hFC8JM0Age36A/gGwx2bZBwPZgkYyQVXhR1Pkr5EBVw+m
EYUTl+dCp+tCK6aqF5iGSa//wc3TVmyD2LvP9kt2aFlS+Q4mGk89+2QmTYQ5RwJG
1zR3pWQT4sEY3wyICd66pTAKujzxPAYngKdtsjYhnmDzZ6vGEpbVr3YaiZGIyKAh
TCYE5Fky7bns49orP/UxSouzQUIq1LQ+0i5MMFDlRUcyNY2DJgBanMfWA8SokUYC
7DSIXV158yXpjsmG1zQDH4bUGsGwwjAgxrVCDcmM6rFCu0OGIMJv/gOmkfMv2AHc
fn3WNdqyGxaE8a8pbfnwKOjlLzSRs9tkeTnhRZR89A+Ul6dMUPG/HPclazbelvBS
HXOUAtRHRElRlVyPXIb3oHasp3aGJS824A/L7UUe2MjQVcAVpXbagR3qaE82YAkh
i4uwpW+HZgZMpoKi20FUgkuZ81d7drsTlTTBRXBSF0Vlz0IuJ4sq9kVyqGc1W5vO
MKF2F2gcsiNMq53zet4YSM3rTpgT5J5dMVXg+cQkSjoLxanOb+tNjFyXGrENO86I
uOlXDLiUuIEIf8ppZ9t91v+yIY0JCJ84DnM+WCjh2p6jR0q4jNDwPN7DtZjq0fmp
eFf1eEg4Xd98lrL0qeXQ22aQbUCbJgJEa4XyHi5m63tJlwO9y2A4J2cBCcfn6PoJ
hEhZOJUf1GG6rV01lCpokS/TNs3YniolKAweW++y+RugtS51zTJuslxjRcT75+Fx
O1CuowWSGu0XntyIpDn6JLFj9o3XQqe9ONFESrXaxirhgR4PvH1xpG5cLzx3XNdS
+qiGDxJ1spRiuRleYflJ/C+/oWi0hPDQ0MPKSUn5rX1F/SG5sub5hRxe1VlcuqCF
mF8Nwx0XDt2X117c8Zr1VioLrE+hDtCiQxhN1/pt9Q5rFoVI4f1ohduot0w9d6SU
kUJDQbN4m21PCSxJ6qQLUGFFKc2KkwDipyG4fWfPhgWl4mz9HMtHkCnkIEt0403V
ZrC8fP+6wmPA7UjRGAAB9ynCksie8Bx9TfS5gjN0RTnHWXBeefVgk5GJcIeB1+G6
ua0PeP7m/pbC+XgYsBgj0OH+ZP3279pKS05RlQxh4XC9NjFFtbzBgujU8cSVYiAF
NvgG2DAXKf/GqD8B38JelsQ7MRR2/uBjTAFCREm6DpXusrRdwTvD3SOR9dL3LZwC
Z1XvDeFUQra8Z5grNlPCUvswlrznfyCGI4XB1GBGpNX1ORFgIAq3WVsM0RQjMzGa
Qz5plqkt3Oc1W+IBjPbdN6AC+LAQ0pAnsB6UoWBbTdRMoAJ3Ft0nNoBVeo4YrFD/
li6JFXymFVJShfD00f9jALrpZC4gvAANxd0wRSFDTWjLIZA2CGFEe9yHEmxKkH7i
qp0IBvqtEx1yZtD/B0qD+nUw4KhtbhBzmdUxYyYwC5tsXbYPYnjK/OrK2gppgXMI
pmZfVtxMZVppKrrY75eB2dgfkaU36j+3kX8WUOGb2zjWqunJyzXqGRbdMQr1YZAY
wgEp2pLLAKIbECFe0GlrZwxPcem7mMtCiXrpPvdXrUzpbzTFT53ZYPj6tkAxJcVi
3zdRRuCJWrkT9iP1qbpYUOQzOFqlt7Ee7AHb2h3FxxwNZRM836yVoF/cqtSHFmWf
CteZPrryECpzhkgDMMwz2zEy3sXII07afpP6hpkmmk8RG3YgTYW3AR8O6INlvyvd
c/5igUIBj/KSGJYPzWJKayyPtbIM5vepJY6AEHsT1Kb2V3+IxLljpe4UEmsUO+TV
d42J2aZqkpS9U/ueZkAXLxG1xLuzmoS5aUKhipL/fp82wzXRrcrq+qDpnBlUzT3W
rk85E5Uw+6pCrDkg1CnEPCPUAo4QIXfuy9UgIZI5vLcxmwmMM7k9aZcQcNBAeMS5
SNSD3CBMydByZXWC1dIwjROQO11fsEXz75LjuEPY7UFSHczJ+cvCgb4AyU/G9Cc8
9GBZPFKsD14iOBOzcXl7Xitcc4CXLft7NW9teq4ROjAF5rHoJRO4B2yPclj30eg6
MMrR8QN6rRcNtMwIS8hiHdvq0/YTlFsCixcwmCLkvnmDWG97shdZgoSRsyCN6h5T
kuvnwEuMitQbpS+USJUeznKk6fsj3O9WZCeNfPJYW3ey1MRBxaAXa886wKlMi33w
yHltfvNEi9n36GiyE7lPFjRvnRGM/QOhuPLI3VzOyeOPTppLzzaEXintMUaWV3+a
z4iV8aXUcHGbQlCK/kSDBXCkWGJ8u0AWTeyrRthPKLgCbAqRrZL6qldzZs8Naofx
xhuokjQZ0/mu6hANM3SD+b01pmHvx5nV6rUPdi5FoO1hqrc2QOJi22IpbFDx0zg0
dlAdjC3eaZBnePsSWQRmVrvFEngo6q++eIxgXQW2Hu/Yi1IEhOSQGAnxV9I/My4N
DoBGQRZHXOVUCLMIvu9RoPipDjSU1O9GhBdbep7lyUD8pSq2KxB1eMtz/SyPt8HF
kgejX9ERAaMVjdMtg4mU9GR36XelDjU1LlOqJv1Ey0NV7WhERrJMxJhItNT0vxwt
ezv/f02c4i+mCpXrRFivizzCA/DNa484ApZcvippAkmFU2TiUZCy8L9EZs1kryza
RbKsHzvqO9Hob+JzwDU80K8Viz4JaiqgzB9G/G/GiPJ5pF+27ftQgd5YMNID9576
bWLFYZ/WBAXxLKJNrHkFvW1RscDGr6QWhADeBxUBCOAkAXFRdu2CH3vdZhjk6KXh
NlS4Vz9ulQC4LCMvJEA/fv3oPLBSkZUWiq84LVS1qdGhlsRekwj0XBuWEdFdhv+V
IfQCBYoJhusIgf6mj8/q88bXLsDNzWYWdPmaiI/GwzPlgWadnow0pXnKpFlMT1BK
n0yKoq3B7jKsJYfmzP6CwOjr5toCB+PaImNa0eoHfPojoauQJog1jbjBq8aJ7+0j
m1nJNgRrFOUecUk3oLSnceLLbsHwprbaSKzhr5pFhRZDYfU59SjpGL1HnKY2mbL2
JADPjMpOsl3inYmEnIhZOtMOspC439j7V5SWsSQBYZJDg7VKjL1eYfNITmpNfF4w
BDETQj0lhjiMl087QBQje0o6BSytVgZDdcTO816xKisz4MGd4e7QFwtcHgq+Yu3j
PQDiDhbBo7+MdA+mt4ENKP02iJH0vfMqBWKKlsiM63wP9DTV82GcQsziwHWUYwZx
9KGSmXJSK+DiDQuC3rAAXR0/Qaa/FvkVh57oB6tX8Ia33sBkfkcDUpbmkfiJT/8F
b9y/1ReDhkZR+2jAg9hRv9+a80xfFgs/s1q4Dp7s8znWN6uAU+etFUgl/D3Sb1de
5HHfbDjORYPav81mKE7t5UANR1mumKp/V8xQ1BisrIRS2nZfaTyj3wOwbYglyCs2
oRdfyZj+IxCRjL5n3zMn+9l8qziAXI/SsyaWjAmleVDwmdBhoJXLx9mfpGl4SlsJ
1On0o3ZvL1ri/UmBoyPFjP8bOKI5ZwoIA8KhVONbImR109/9Yd5AZWcBrCOziFU0
tHB9GYJS+jcJ3gZPEMCuvQHWBaKyapPavrsge6rNVrhDneasScje7EZ94OgKEGON
1gLT0vM50xj0TCIB+Kk/XCDJ7fu1/FMIdiWI7gk4lduIFpfHhHj7G2pV5q003ocW
w7zq3+1Hrx7vz3gH0/LSetGDO7LP8V3dI18B1KznLOpEwjo3e7eQm3Ok8xCWRmaf
6u+ngDzIIiN1xLDZAp6PK478n6MFhdsy3gSy7S0Yh4yjjU7OWUW2S5F1E8mzRtuG
yKj+fwY83jjg+MoC3XNJsOkUsbwlOgFPyJeUkw70aOiT8ZjlacL2C5eEgvKKWDcp
pu0FuE5mLN2qs7YSz2Tm7uZDqVaThZNCXo/mx4hY4SeUW+umgnZk+z9Ooag/ORC2
icPLJiLwaFHlbftF10lx6hA/r29meK8h8Ei4l+Jm475DoogmgVvuqfkKjivERBrG
zS1INHn5zF3C42nvHei3Iu42phxL7K4NMZA1EuqN97r18DyQAmBKgX/FF+cK1rm7
aNS257b640yKiMI4/FzfsCScl6HVe56Woz2YkBxnY56ozP73PcJQ7xxCA2wNYFJt
MKsqCwS2PO9w/qfFtrkP6++gvZQ/HiSfIpZf0i4iNS+WCrV1xRF0o1VkKlj3esAz
gApJFOi2mKGuUHS3+OeEKu3jVYdljyTtHaa/LdrgDVGWWACTapYEmCMaqyol66Sa
n4Sv0gvQm94r6m32nOqO5PqgkgSgHd8xDkqIX7tPImVwov020cZyRxmvYC7sn0LL
gygKPgoi+T6oNOqG96+hpGDRP8t56Bk9VaAMqvSv7pmqBEOXisOTnjUNbhBJqmMt
+M/rD9xq8p2Fc0J9ImD4WkH24umY6IeE56d1ioP1SygxIA7caPasEmalQ+Fn58zI
bv9TT3sYoVTLun/wovQnfUNzUb7a4n289EUjt6qkZS+uWIkCCgjpuzcN+ntmEL3E
OjzW2i4ZvWox2qQdV0v5KJgFrt9/cpOhDSZbiV3MX2np479Kqg4AKmWzOpTKE1jF
XaKIOrIOXPPXHhBmYAF+XcRw4VEJcOJ5e99C8v1/bfx4M4RFUGkx9ArEoZpgfu1u
FNSOVMYtBQQdfUevJ9sO3D3tDSdDO5MBquP/+NZhyYYdbiEZvJ/TfeCk2VgeBESa
r11jadrdi1wnZipRRTUulZlg9UMyapMptdaF8SU5O8DQ2DL/QVE7UC2PT7Cs/qma
XlM/XOs+nsyrAgJobOsWJAFXL9Elsqxdd+8+GLffWnNzSo6VSKFD2IJ1IpRh80po
uhONGXbClZznA7jVwYeGh06KFWTj5Ib6SCWNyYEy18v7vkk8EeU9HQoaI1WCqs7d
yHe44QBCVa+w6dHh8ExI+XLN22SDWxpA0F+A1Y9nGtv4CAmkqL3UAkgGC5nJkTar
UMNy6YVXC+udhA2iA3H5aXOkzvmq/ee7KgCZCOhuqEyKhj0e2ovWOIGH8cyIoT/K
fbkLUdfcLR34svqBhxTQ7u+o0lWtrT1ga++95q0jXX8lY6B/jWowU/IO5HoBQ/Hj
GdXDQtVwnga2WL+J0FZZ7fw3AUYPL/5I+FGDCjOX5qcUR8rQozqOzy05rBN6nljT
g7gmAhueMkf1qomhwHnqTG3UdbpQCZ48vT8hrHG3qX1Pt/lz8ESHF+LIptD1BgeI
g5apY8y/7KwC4ZdkJ3CkDRltbn8Af2H3yyk8p7PfrnH2eWShn8OgMej8O9LLA990
RG45aNzpiapTPHMsDGG92qdpItba4hYKr7x4WrN95AJwbqypMshnjDR/TKW//eRS
ReHASEubKgszJwhB3dVF2C9h2o0o3puJV3bXgKX6LhgeggvSBV9Mq/QSIdHq4Ze0
JJgnwXaBBkUDKEeMSZqILNo+G0t6lAqM3lSkA5ja/p4EhcZytpdP0indq0d3QsZL
zRCjIMeo1lrvknFxhkPyp90rSzuGcUpqgUL8Z7keO7EuO9iz5uht2bRZpCxotse6
YX4+9tPmI1HwkuVZJLmlBC/sEtn6AWYlCtYCfAtDbPM0MCpEBZ4ONoiZWGRXoTCJ
YID7kzycwDwDn8Yju2mo3LXnQGiibWmjwo+1VxkBYAp01YiBOOl6V5XLveluagdK
bH5xCOjM4LnSiKQZqSw8uD0r4vuHTDN/FQXhkR2qJpY5KQtqLCDoquj9TR2YiHxu
ECkpOIEYqmeRBCccZmPSGV6NjVigtZxeYtj0SJPmczlTD2R/k6ty1Q/T100ZW8rU
J4aQ1G4ACHyr1zIsXBGP8GIeJzNRDDHDl3iCA5mqYSCLtbfV1C4+K3dJ+GCcp6a3
UrvgiMXt3z/s/UusZENJ5GqXi9bZl/cni33RewDYBxMkvATMSv6iFdFDNIhtVjNI
dkGY2wtPWKS0KUy+IbXtKDLLaToG9KKLkojspUxVFoMnC+5pFemkP3/hAmOioQxl
3ctqAXWBBknWbyRV0KiIUZ3XLZ9ciymaZ2mjRYL4hDeHUvW+5ZwrRhbicDeimRGW
jz4kgicT591LyaxI0Jjl7iuZsMjoDzjLwKZkfskRI8rfbTMaXVQdRPWaBUKIyPWO
ROG6zjhpertdQHZ0HC+VfcEFAPeQBRwFACP63W3aXSdwpLyYvyCP0JB+gnCG+nK7
i8wHD/JZT5f+N4abIf2mu1IacSJ2MINEdiJOZDNDo7s2o3Rh48zHK8evExx30E3J
2Ag0QpZQcqPRQ8ye3JqCCB04UprP4OBC5HnPuDwsbsYHmFHVKRN7LWTzpO6pEV8d
65a27v6+yNidu2KXPY70CFyDxeWuROJi5rgqhP9JPRgIrMjpelMEcu0bmlO8QjrZ
/HXssPGH9t1azMWOZg+lv4c8SbzqxRGcODP+qxq1AncM2r4QcVSj4hTru5UAFYNI
ji4+GICLfkQF2k5zJBgqdE3endcPvZM6co19VUjaMtnr9ZpUvuvbSA37FFf2q73i
OcM6vKEvUDVrzy24T+LF9PGXHs24Uj6qI49J7a+kkGWZiUDYhgPLiBWq26Y+pZ1U
EgN+Cyvnm3t+tgPrNA70AYZMefZ2+/Ce+CBUarH5TieYvs94Fj0/Kd+CONPKeeWK
t1O5z0oNhdSxfaW3yiynUnHu7x/ZAUCTBD/AyCRXCI9T5y7nQQECwOcaYxDyFgTJ
Nw+CnBoR4fEOleT7Inl4r74+zh6g6Hkavsi/ZIF9jtl7CdrjXvKd7lMtSZHrjTon
PkMdmXqSq851kOK3CAbl7BC/7Iiajdhjvt7RGrFf6TWpL/vh6hqNeuuqT+g50Noj
ZCXUPN6k4C2ukfpp3qjbTSElH99Sh0dT44nwX1sp6bFFdQJo2+GUqVIc9Ouw5mU8
jkO2DT27ZGrDV/1afBeTg1L6kaNZDEeUr78VUExf0ElOCT3uPWf1KeaFj6s6MWjK
zLPPhor/JjdYLYYpbSQDl/OoSRgZ5zzmxl7kQj1O3nrB97Dsr0aRwLCOQ+hJje06
ooYbVyuzkxbfdmHGtDv02rj/Mcg76/6n6u3fpTNas9r2l00jxoW6He5Ahb9TpqLi
wV8Z8MMsQ6nM97HIRL55zkbIRIP3ODM+zyoa3k1e09yghz3h81it1heUemiMTNw6
onRKCZ7RPfNWv80p6GF3WI5g7w60hYU08//v+M+N14mpyhi0Bx8+Co6C11AjDp6i
jxj8X7M4VASF5x7xXK5k+5d3lQdA3n8WJzTYMyF9K2H3EG0LW4TYT0d6ftaO/Q2D
8n1rGWdSVhUREjfVsxGAupt3JsUvz5p1N6/0Pkj6e8FJ8lcV8sZJLhua6EUXEHqL
Gcpyq2MAEZu20s9IBeZ0kPQUCxH1oka5X3VMA++9eVsxYuSF/vbN2A1hnz7GeaWr
eiRGEOiBZ+y+3zP7jD9CXXd+XkFhIgI/n6zW2Eef8CfWcZ/I/9cSZsLbxelmAzyv
oMIpOMNN41QRiD7ovbvsgHc2/kT0panRKeWfniM9Up6NEoyaKoy2bxTuE3uT9pF0
qNu4wmhTB0+mqY41hlKRmroRwBlVe5Z14UGw/6eNPFYND6mXmmp0B0fq8ykFTFer
FJHYK79Vf9UPsLh6vJw6OXqeVpK3bQ8VtVbyW9fyZVnLdROQlmMthyKqIIUZbTo0
QEpe8z3NSCCc+ji/DUe9TkYXYE3Mg8tZkj82H7pk+h5UNJ5Nh2d1NRPEmUlp8bVw
/JHfSv4xRpwW+FsOARMRcvz6uiLGDHmug/m+4E/tqCZ04mt/thZPqQFYqej31hgB
BIt4TT8pdc4BhsPAd1j0Pzmth2Wixoyrv/2zqy4o3T/nbg31lXBlXpOF7vvxMJmU
qaLAnU30UnERZc81V+yskL0FpAyyLTa8tvG5ZCdsW9PuNKHaWF9u5OtLoDWLxb8+
ykkz39eyJKt5thgD2lKTxC0Zv8TUy+QtjPD5dZN1CgRmImryfeNX3Uk92HXWz7Yd
+BGLNdQPRzJSxzwPT7tPU7C5M731s6gCzhRRcNDHOJTKtfDleP5ptv+MxbQWZ4PR
z+ZWx5U/xqh1pMCdjNowAqLJkMn+wqiNA3Ll+I4EtSDgEjZwhW7YJXSdV26TFE4W
zpNCcLDJ8iMeTQUT8TJwr5XtZWm08RiEiv1mjKJqP/4=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GA0w8QJfUFkCwAuNC14A2OPnVDdQqvL/rHtQYxwCgAQRm3/8lM1oJVxDLmAXC0rt
YpuB5M96UBLPpTDNzkcz0YSxAabcZ/RH79shYN1j04cW8/2eeece+GRKOgeAz4a/
p/0gvIfFKe/EYZwVlQaYdRUzUwZwGDvlUck1axwUnXEj39DmBeY5tBbxmdXqoFKv
/oZDA7sPc/1VZCKQpX+VnqGfhp2qY/AeRFscI56RlbXGUrZGgWmplq03+qIYGVww
icHZNSPEmiw2Zxfi08BMWwHDzxhuPLu0VYxwr2un8ZTmEFKLgY3gxO+n/Ms0Bx28
eKrkU+jxcznZKZTofliFGg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4336 )
`pragma protect data_block
Wan+JTOmavfR6vfVY7/HHgmTd59vBzl0IHk/SNctx45gGq+IGYVu3RcrSfOh2KL6
H8ytdqqXG9b11FJpg1Fudm7jwD7nnhJBHh+2Hcg2cjw2BYy5LIb9PPg5wtG2NKCQ
jk1/ONE1S53+gpgyquL/QUsFYT9ACBAZsgzw1+o9zAl6Q1kEGLOK4OnpIV5uafu7
phIyMkG0gVA4QibHbyYA+ymRslbPWujenDldweIk0E2q2amLYta/ljQHJKVcJMHm
OdsUWgrtO0f8VSaeTx+J1gKkMN1yvWsx6BRd+8y1q9rsbtMNJD+ETGaXQ0D4MR88
rnUqNbLNMvY8kfI0YJFfPgtfcTeKT7hSpZzTC6bkRXAyeqCqsq4VCesR8KvS/x1I
03U7N2NLjPtYH5UQuoSOqtSfdTw88uZj8mbigGZufHALJUOsOMZ6rl/+X4raS+Iy
+fPg0y4JFsRqXBtybwDm6J99n6iCpuR5d0rR/wcucVy0no10XfIwDv8QEi6Hgvj9
ey57fyodWZRD66TcF4V3kPNFN8+MXE4bRlmOEuMToWNsn6b7b1qN9lUmA6TgKAPX
nIWh7QV4UB5WGNOxe444oBlBwpBtnheQIsjCKd2z89VukCtFZ4Y7/bk+QpEGO88W
KpqBKwUW7B+xNYI0Kk9HTmzWYH4G+rLgScnJzevqCWP+h2qetEgCjvH4Sf7BSY3T
pMLY1juLds0LgsWuV7IQ77mSPZl7bYUpZLJj6CdO61ww7noPuLH68VHz33en9POl
4FiwQtxJDzqx/WMN1xgbHeXKYXUplFNdWP235P1p2VJ8M2wGf3BHQgYGbhQ1AWHN
DjQpHe7vKFn5DKOahOqTeOtVsgpITGgRJLQhbdWjtyRdJ+V34guE4Muqs2bf40j+
dQfmRFSoAhKlR4h+td7lfTCoj2O8k2y+pqE9i4Cul+wB18x4Gtj4hjK+CDWtJjj3
WZMBE7s8GHIvLr0rtRkH6s0/hlqdlIJzGkte0eeWDmQ47s9EpPKwZqaT/1eFrlle
x5FYw4bX7lBjUlPVolUUCHxfsaN6fPejqe/7g7KBoZ2Hn3NIoOoFDPWDILupRLVT
pI/jLKIplcTBsrAuB7GrXloEeCC9m+bvKQnAXHSNCjX91EYMSy+7VhR3xdIg4COU
ruFjAoBNw06RARgThluNu953myxrNJLyEJo9JC61GeoUNoQFgEPEHoZnWBgQ7x2C
9nDxP6jOyZtRnnagU7f/oLK6ACRDVDaq/JU+csbEH92H67feSA+p+1L44fkwmxAp
idRsg6glxGqbUIbLnl3lkbmAdF8w2UtkEnWuEoM7p5gw11YsG+m9scuDdzt3xggs
5F2JyAcvrlC8SaE3xZoHGlDImgZ1eqlEpJcBXIHEuEKgwLH39c/ohKFjhwFZ1UiO
CoOOa1Ce9Hi8H/kMFLLYVNiTyE9Vx/ZERSQzj7pxwE503xbZReMOMLym/n9kShQ+
Q3kDnCvQstRFcWludVZ0Srp3LlDupmF+pxaJNbAGcpFpx3lv5byAdG8TvIPY7xvo
2wWo2Yben5OjCZjyanzifI8qNdVvBtd2T+gzwWGB70BXyflgkzFwIzyhDjTsa+KH
pw1W8KZ1SuP7fwb2tpuf0ZKGAvyyYSt1IK9wzjpsXrJ/E+8ljSiTsls6rfmQa6/Z
p1ITG9TAfe9rOpeYi37H5DGPeKxoLMPVclmlrEKMcoDR/Qe9r5R3y2nu/fmHIfXx
vfMdW+vBso134Z39Sg3LaoInfdNsVpCrNU3dKKlEOVy7Zm216Y0f3u1ul541RF9Y
MtlJVMzFUx03q6IZnmukH4mdZWYs8jSfqDIM6F0podyk8VjH0hIiD2q0Vvyp4rSg
zt+wQswgQAhYNZuaZ4N29TBDYcDRQgqe2YOK50B/HwKlklWRtzBtGpFG7C2c+yqG
jS+sev3+5LqrM5ojpk1nBQY/n4/Dfp21Z0dh6OlgMbYA+e7qsuoAuwTOOn6oK0de
t8EtULrQRV0UNG4MkRkBVbHtO/HCme/EJT561BQY80zWfvXtnzkGtSiD7Kbsnj3d
Nr64Oz1dYktMhq4c8D3sJyotN5f0IQrQ6iVPrXny1yFyGRW2Qgfehulx8Gyz4cNJ
1nlbGZd2rlZWNHDYqmEKlvAP1gJwr8tJLNscK6I+zMxH/j363IOW93Y+E50fPWag
iEZ5hAU2EFyykr1Yut7Dw+2Qp25qTWtin8bguW12a+aYbshiiUebxdnFcqTO5VCV
VHCwD5ffJz3G9R0YgVPARzkkgqT+VT8DEL6/M91eDB4cT+kNfjnyRGMs6G3hC3Wf
pjsjaAfNdo92sTivf7vMNmtZks+6sUyky1D2f7mCTxGur4bX+1FLLjRRp4Y/O/zo
XWG/nFR4jX29ZCS+bbVDIc7p3QlmH1OXnhpjGNO4EZbnqiDyMKuJ9gvb+DbRVprO
jBVU1JOds0lbmejPDPodSn5lkvdpah5KQy7GW47tbitZrylPlNXSxMlpFpUonOYg
4ErF7Nv+lKvxA6Lyzedh9SaUIY1pHYGIj/2FuJOAqMNhNva+blZ0Hm/mvoW5bS46
eajpACGXDwA+pDC3dy4NAjDNyAWILODiaLRJ4RFL2VYT3WzJVPvZwaSPoP+rO7y6
QcA9Xcw8lyRc/VUtqJ+WfJkk9b+iI4Mde94KE7en3nskpLtubhyX+NrqEyyRpKwo
mx5gZTzUszV4wsy/wz69J/LvQq/vOO+a3iHi57bs2wJSZnkl4X3hvFl73N6y0jFk
PznApDSMRWpRFcVnTp/pecFf7pYVA+4xVmjEhWkRjTytX0emGYLQpbvHZm7QTf9p
FGGNtzif1pcWyVpcYM1C0fJmtXD+cJy0Bn1y9ObGKEcRpwQxvdBH8i1FTts3qMTP
WYxcj8PKsVwmwbKmZzZ7n34+Dcpa2eds73sIKNc+jrAEiAhUkLXDsQj0Vh1AZtvn
yhxO6Sf7lYywx2r6HVdauulrt3gmQqulTQyPH/+1I8amsZguk82m/GZyV/diZMyY
OgByr7DkSmq7sj1gHptMrFueiRf3qhSEsts/yQg2mcZexrYKylHkyvS1qAXdMGkV
eHTrYhNicWpjnzJmzo7mKCw4srYMdJZZerF3aVJht4s6n81TrsGZw0nOAlc5F45e
wcy6ideUCvInvruCny+0rMtzAyQE632i3EPhvbdxcYPhDO56RQU+xwGNQarDevy4
1c7y8etws+NgxD6udju8Eyoj7OxpvovQFhPK8gm908VmHi0MSxqHShuVmJeGncQ3
ZmIovAD1WiZT7BXLOoi/gFGqLkKAnRuABNHnhzGzHxch8OxJS2UJWm4QfQntAnKj
jCA/uLgmninUwOPd6QXpucsU5UK3kja8MkA4NANbjcfQpqQa4UnyJxBR/5L4zNN5
ZRnocbeW+tVvpvCTOsAxfTyVZV8iF99xG3T3O6K9ZTG65jOvpMf6ged1H4J1HvA4
XKZhYGanM8UDaFy3K/7TteZOjXg//0c7Z9piVBemdNt6JDMhckYOM4JoadWc+g3z
cElVVRVKcksLz4af9o3L6oBA7+uzZk/Ib2B6d0ZsgwfEqzVDcoGLZ01T4kBSuiXT
BBqle9W+gmVrkvopmdWtNrOpt9AvyrLaqMGxHlY9/1PGfoN6JUu9v12Puybb5+ND
2rLHRu713/aQrtUsos14TiZx3hrPZxS/5QwtVpjOtZMxR53uTqix/Wqaer+uMVQl
cFWspaYBrB836tTwTdPBgfXKlMA7TCmd/wpTgxHZWeX3O0rSQFb5hegkXUupXRLB
f7HQxhYPVHv+lwjBtmshkgAE+YWB3s+OirxaoGaOHaqMsNQFpfes3TLD1xO1SMEn
tYjthwAzh+r6V4C2GbWlW9OAUXC4xlVYQxm/cbpSfgTupHbDhJGoNMs7XXuYZ8IH
b+OXZ0z6i0qh4+W+k2bKTvH/xqhhJcrG3/qYHCXM4WXAYRbWjldWj97zMiM9qu9g
mSEfZM/O57p9qrBc8XssYauj/Ae1r4fL1GAhcroUnJiKkNyBDZvJ5N9QRVER6tOY
HwwXlPvhkyEv7XNzWF5aeyeNgm4MWKfKi6yn38zpApXVwI85KYfHS8+ZVgQAChDd
Ugk6EfOf8RDLYHdfu6LpO5odPhHss3EQd78Ew5tXJkD8qphdhuriekqR3FBio0WJ
sBFo/okWGYJF6eSSyauo/UaKtFB8E59e+n+5hpodPLYO9JGCG24jnD554LJSINY5
xdKlgUD6rnCxol6XXgQcMlJRN6Uq0pEc+abD48uIeViNpdLr0lHRvxhbNB6to/4k
lexKtlKexuvuTVudlAFVA8bik8G8ukJYPvLHa24fglMYEv8EvhVBf6hGRpjgKFlX
SVL7TM0erKbTTaZTWifk4j5wOmyuSWe4GCPz0x1p/KRv+usJlRTxhIzV50UygsKA
QX+ATv2ly/teO9n481H7XLHXvp+MnpZD2/ASbZGy0pmyMonZfex62YZS2xXhjHmB
Ifi8O0Uv667g+dvDnkb2ncxnwrI7eDf5l37TPWHAAoBL1lsJT68CXli5CzLH1Yjb
wOP8VjYneEvNTyzSnt5snoc7ezuBPAeWwWuj94btMydTXx6Chm9fEfUeUWqqWYvV
cB4fvvJt16fZ0osWPH5lR1P8Lev6VTAL3S8r3dqc55yMMvdB5jL2VN2inREAeQrC
+R4qsetlgzr6DnQrXTrF7l9bPfGgSjVGKuxZ9kIGJBvXgFhiojEB9phySMb07Fws
ROuXrOqN0gss2l5YHa1qqWZRIOnPMmbhBww8kDzfO4hQ3dh5fW/VcjXQ1R8KEGSm
ksRIz7eoRHbMOtqs0wJFM5+EQEE6l6yPWQBO+ZxfnzeqJekW43PH7Mb5JGnTeBlu
C5DyOqvcuu7/DQosHL5DBpFCV4bHhaZgTMq8WHTuPyepM/0+5MCoB/ZRGK5KSosV
ig9y3fpD4yq2K57uIrOXQY0ZXLqe9fs5AFX7A1p0elDQLm0LV9imIQDab4+WlT99
cIZ+a/Rs3AUPYPPP/qzFoykXWcvwsLyan3xaoPtrdxgaCC+TzRcmPHLHa4mNLT6A
zBNubXQ2Fp29csKEo6QveNrxsYX3JMWTf7ArhuZea9u288K9vxG2BJ/fBHE80m1B
B+naxaqUHuZuBhvvKSh0BOmqfT/ms0QqeNVHeVL6TTKsMyMLstZCq/+N/Z77qp6D
v/CS+eyNcJ1BWmOWUQYEfJJqfzBl8jLg/j4I54yZCV+uhfNeGW9sHDNjjpU7aG8B
jE+apK9Myq7LiZC869qDVjbq2fzcslk7eI6uf2AQ8sz4I2p2BSWaNkx4nxandJvJ
Cm2nUvTdTGMaEjvgsIcTx4dUzO3+YeIZNU+w5uuULL3LGqFWrRoCvj8fPFzGBq+9
8DbeEFDznCBNsB6NCpIy1bkAvq+PvpfejOog2fY/KisiNArL/f9IZrAlsccNbpCA
knmOL6bXop2tdNKNB+lr8KG8aezXIaser8Nla0DCrN2BfNty6HllD5+Pqu9TM9fR
jSJKO3YxJMarupa2yZNsZF2ekRK9hCsOsqCPD8JPQJjU62ItwiFP7X2iYGrJVlYF
a5ywxzr1DSqcy/Ii6GijFk5BZ9UYzkRoMIR6KpuhdhuS1V5nwQ7eiMtop6EVgf6m
rKsJY1JbijNkZBe3pEqU6fK5SBE7hBZTFcWSPSRXz+rjGxR6MExnqC9ZL3vG7IN2
8Mue+Tqp+Y9s5yhgUm1w0dx2K/klnJBxCDYYY77MSCokofYT1IebspJKFe17s2ZZ
MuNwmVNQJlCZ2FuHsXUMVQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
L+OB6r+6msaKXwsC2vBIb6daCuW6ru0Axog67EMGEXJgwyD50E1ck8jDwoveAY+l
IE5wS739QYfl+Kiz38WdR3XIGcb7ocqULZgufIK+hvOs7936Eq+oJm2SySYYKNI6
I8WdHQ1EsPaIU2q8qDyZSgi1RWhnNkWGvUs0r4KFh9yrcW4OaW9Q0fGVDY4M+yDe
rM6mvVLlFW2rUuZY9r+yJ7s39NiPpFVRRwuysw1uGb7RU+Z5T6cKhWzGFc9lCpZF
lL8aClN2W6QwN4s7YBycR7mpoaTzQS2BfBIrzmX5VbOKy7cqczTdN2uBf0QDcu+z
njjRvhacwfhgLVnt1LhFvw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6560 )
`pragma protect data_block
syhF5sSEU2PBQuF3SSRw+EB4UsGzF1kDHAA9tgQ3zXSnS8dBLSSpit0tD64VsAWb
WC8A2C/0ChJUVOzfRGdrgKRvMYs0kzM1jNFcgL1rBxwKS5GrnLvDw6mj5+jsBwur
iw673NHXLQNGqeQ+iC5fLXPrb0c+uQ6ksEPMDxq+9B6WR5X5skIulP4igqZnwsq7
6IhLTWvUMGTK9TVgTd9ertQ88atxvAdrgqytv7z6VojZEqGb+bfYky16Xm4QITs1
UxuQoqI08i4T3Hk/8T5jSbkqd2p0hMSbiPLMM5Se6KZxqDnNIGJFIFf+WaKKEL+w
6bwPgXQNiP5WnspjzIrFjdYdkMCfvvmfQyopB7HKi3qhfYfUSpYgZ1E5u1X6/Rip
KKj6XL80tx6V1Pmow4UPoYEUD20NW7UeOQTW/bZQrivCJaxvPcj+9v00WTjxrM0b
DlgdA6hTzVPWwRZBRRAxe3TA6vr6dcUMbmANPVKkeUOKb0gs8aKexAYSh4l9Gmiw
5gSd7fa/wd18LSuxYK7OgzBKqlH4gWRmuRMPWpIEwbVdO7WhMoqQ23zqfV0umkee
6LSUV0ZJ6ThHJfaMdH67M+DqZReBxftveGjHo2xwT2v/SGsMw1VJnSEjPSkAuBcx
4lydI+p+Okn52qrw+/vDeIZ0lJCuuDyrrmszYGCwD1nV/zNix+4q3yax2vkuBg9X
TaVY9N6ymLKocl/vWfynGFmMY8SOfX3E4cocj5PWBjhHme3MyPHTByu1lS5w7rIl
C8yfGGruXPVtVNWOM7UT4XkV4qqJ7s1Ftrga6YXUy5U1YuqaTFd2sG0wgFoTlLeQ
uAe0fNT2Su8zSK+5PTRQ+PATozAkgz4zdmsp7QSQ6d0ZJf6g66EQPWZL5LfBRIVp
v0NKkjtpeyitKhLKbkrMXB6Wf6wu3YthNZnzuAFNXnQfzQvBeg3m08JtICPzWPv+
J/IDwjWJHfYmT5ErLhLDBcBSrBPHXOJ/CFYiQdmBB9WRjBcM4a15F3gSbZryURSG
As/JibsV3szfpYYBtbldXANKOf899J3BDg0oLVDiCvooN0XQXRfkWlb9BJnorhV7
u0hpOVmCQbPqQKUCW4j3O4eU80TPQCghRRHDfQ/4cgXzldlKtXXSHoEFEf3nwLIr
GvGnLbLMDT3oiwiLssgVSryrh5ks+2GiLwKIFnamESUnjho/Cu2Qu7cOBcqL30Jp
4qxakFgLYH3QsE0Zw6YwKzaEr9A3byyBUTo0IdRcKsCZm0GdPa9KUS/39FKXL/aq
aG1+++EkG0+hFjWzJshY3+bFh6CclIN693DtljnLNv9eC2qDyTGPvyhJvUcRIa/4
1wfoU1ci0181nVo15AI8rS2gcCLQ0Xg9W9QhLSzNsuCzYqlyhIbXgrwX5NLXID5E
SEuGrHXcjpRiquiivYI4E1FcWvhDka66Z1uxowHZpEyhlYItrRFOlXjEs+6fcMvG
z6TRxzFwUNAgvUGk7SyHedQ2qxefbml+UKoF2o5kTQlffRjyP940upPdyHFBgOX8
FbVgXQpy43zhss5NI0XShEY2SB9S0CnLuaAKOuoMYzFcO3ZIYqAVxZ3UBLQvdvzr
cv81qgAAbJPOksRDqs+p74qVRksPw86DuTkK7gMVhWcPxP/8iFdztcy32f6+IYZI
UppKWpCJSIafIlLR3o+JEpbmSXpaWm95Q/6/tBNpH4EFcrjr9MST8hpIAW9XNFrt
yDP/TO8fB5LIBWrhlbaHod4T9zzUE/Mcamt8Wwc4HB4tI4S/8Vz97wFHz06oNlwI
zcJWLw1Ko/lwK2XNd6dF9l04QGKzi+ST59sBo0+Cp64JhLHftrbIGZTTra2UhLBr
1oEl8e62w2q7cOSidOc8NUGQC00GKrviLF0TAXF60If7TcpmuMZ+r60IRT0yC8RS
shUtvy1tV3tJcKypJivt1VkLs2HES6z+OAe1KYvvCcWPIGvlATbT4rrieXTKETKY
fz67nCJsBRSoBvjHNZZDFcrl2lbPC2b0i/K0lWa3TDqKlzPZn3cjbK6ybjT6Tugc
p1z4qsvF3120xmjlEY8QkXDm/msFiWcIHeKnB2RheIPiYEX0/xcqr8W8BG4R7ZU/
YX8f8N9oUm98lEeYTe7RYsqiZRA2rKaSS+ufEFUtKlF/3z4sAKtE47Qn/z7FqcGr
I2rSNclcP11X1YjhMh/mu5a5HNjOMiwGr5D8GMwIET5JmarUZbfVFRloBRgpSDlU
gwOFAvUifcmGXkNu50Y+EBCJ2uao1Rk0Kdsbn2tdKyym0djO3ugU6gFpeE54PskM
yid6RtcVj85qTPiyLXYTLhUhIi9Y0i8nXaIPsyJpHDfvwE2aNU9xwsygnulq7lFY
fNLd1XlN8t/C/7sEZS2COdKGROSGihB7Vdf7OZsuhfiG/b+RGQz9AgUbjS83TIkw
lJu9VLoyfcQAfrYpY2XChxPgcXWi38OJHANfy9zNSbxbfA6NLnatgk0z5nzplgR3
jSvp6f0BxJT26EmCthhLOCm0ERUr/wH2NvBdOOfa/CRk9B7jZm1Wtn6uSCQQuzoG
ufMjezESXjgwBu/km+QOp35YedtCTDXhBqh/jR1V047/I64cYGIyWGMeehgMeXfp
HS42X68eoLUDCBGBpDPBxtzyJBzLG4m8ixtrOnBjnha16sddseCKSy9EiyGF7RTb
Bx1U3tkUd4UsSwqhJEGEEqby8qQrxHUvXL3QppXHWtrN8wuBJZG5IFye9TcdZhNl
aY53BP2kgoUbXO+oqmqmwl3bxRJTvJPMvaGOSLX3vgapapAEZgHcFwgcHFMPT2/t
yLyfD7smLWf0uyob+6NEqUCxoibbkE38v/+g29vaLutnE7qi4CPnCPAkjkz/LmVg
PW81hxPOuhJ3K/qdUMAu2a/auMC5xe6RYglDXmJyR144t6ZIRh4GnPY79CCggF2b
17biIkWObbFgwrJ2kWdfEuS7mar8L2ugxp8JIjSKnVJCS3NzA1SgzufLAZqTL1Kk
vuPocGz9ke+TFWIF6JuSKoynTjpxdF+sx3pHGR6XMYeYHqvrmiTSXgRGoV/+qJ4o
Wl79OYrEp1gCJZoPO4mPYJn4zQPYcV2uICTPHiPnrEptM7szjUs1hX+dz/CEz0A2
Ru1v6KT2HdiBOXI4OjxatBNPulIRCWjHQy22wgrZuZjBhHKiwkE0ZZY2JkH6ZXlu
cFLpg9bJCo2NkeJxYt13LuVZ4NZa2ToKlinIPoT9P6RQBgzcBeahbXNr/luATT54
Vt/hemLga2uzT19gy8w2WfIggAKWiQH/rYn8YAVI0zk0KRAU2jCD2clqJSBYC/Sn
lJtK2Vtb2/TSOinPm8nLN3rhQ+ABQ1b86zyrEPXewRoy/v3WrQZQQH2+eu9F6NHu
92R9xZ5iBScm8uBhNuCvfAlJNExDNLADpJSLYAUdOs+gylnH0S820bRUQywyNvY7
cQFmYVJ/V9UGOtfzlJmTJINWpfLTM/DEdi9GY0FOWaIBKP8bxEDQRk3mv/Ul6ewo
AfsB4POosY9TjGl4ZYsEd1QWBgnhIPMN/EGIEu38JRt2JWkQmwAW9LwPFek4sJOT
uGrRx6qOvlZGUCdv/fXI6q8KHjtXcSiKbHHQf0Dexn2xgNJ/3R1NzIfzwTBXgrX7
wIGCjJCCv5stwNgQnwOKWGKjMZQaiRTpwBOwLzQjSqFK2925LyeFSP3wkyZ12WCP
wGwRcE9XjQCq/+XqUmUYVSgHyNCD+CgcTX6ndkBuohBxZ6GnsrWNNvBXkyGuOtzP
r6A/39bvT0yNuBgq84sNBxtrMKZY6n3ZP+gxjVHfNhe7onHJ7sWLPC2Csc4nAtlq
wfrGiIs8cGZnhRtfEkWYNmh0gdzqG2zYhsR75hv3vC7HZQU5BQvHfIFPbiWGerOa
Bg5zrw9mNrBHShdUECheczNK+Zzew3p9QU5N8fW3CXAe0+emIRbIdeWlGlsajMdN
kqH9f3sxvopGemacoDaPsciFrTDI0l53yaIkOOCrcWunhAYb+0tjkhDv0pFtYlTo
7hYtr+prfyVZzVyWR2wdmKHkTv51AbgcMBl8Qf78wMco/bBPZNzhlBwn1hBUsAG0
vKvo7fmduVbZHPBFqv90uNbp/dH1laVhcKR0uDxeUmFN20py5UnebueHxqjA2Pnt
lLxv1X15xUy/AUiSs789fMVSKhuuYY2V8dlTpvtXtZcNsoa0RqUeabCQ7ECvOXFj
KczmJTNF3HItZTlheOtJlikt06qqk//YCMVuoqpb/vByCFR7BOfv0lIOZqleCBnr
Ec8bciqomXqe0WZKF0FYlU1fTLGexTRGeAg5G0sGX5ukc8A0X+RNisExtl4eFoK7
PX/+aPCLu1n0IH7KrBe5vDEH6yvNonN+r5En6ms4Q26bNtMcuA/Q9bhIibuk8Q79
qMsrh3j1i8IZ0TEtkIIuw1z2AatlaxFuCcOrSWABKs9JWLfrjACca/kV79xlkpLL
ISlRAEufo+gOMX1/ApeaXHoPPYa2oX+AFrp1HG3j4YYGqtb4ws54UqrmjMVEKobj
3PYMkP8ymq25pEYQIdZHntks+E7BFQifq0mCIiSST2cTqZ7ujyQWQQ2KYVsKxoaK
FL+t4dX+92GVCPDr4shzQSeQEHmF5djwhZC1zBocHPdQGRAiihw8yhMnyLHZmgNX
Ni5/N2N5S+/wFBBudRAdN86ldC7vuRywv8w4yZXbbhLUVvb8sAuMa0mSpkXLsWwe
tdfiLEhXphemSsG8quEz2g6UPs75f6g7lJ12w7RSoovxEizdH4i+/337D4DOam15
IsxuUhOJpntyO6iWbl5zAS/zDLWX1gdFLWmr7z3hIVIQbT6/6wZIG5ZK/mpzICac
8d5KAD2m+Zn2ibqhWnI3zdglvuqKc7GVmqQC/i4epudy89aSmfred9bLSa2tkZmY
l07TssadBKCpxB2kQkqAiIOKRFQn0VxrrDs0s3nCWpF6CG9LbRq19iSiQoROuFJV
a4szVuWCwgnpVHVLhKZaeMNK5SWzQjJHnoGVlu64WOENMEnRzbN0tZIMjMt7g28Y
jNoGMq7oVfYtBF6wemb6bSGAmhjWxW/niUGViXyERhT2ad2JEp4ZXfUGwgsLKIk6
Uxto5GCEHzLgLPSEOZVKMxVEzP7Gtwx4RIm51+XgBZBUU2fom5qh3w/Mn6eiwcH7
+TghYpfar4DG2IBTSdKHHf85flTtLhsR4OQcURKmsDDGJFGoLaVo8JA/Mg2zdXmr
oN8l7UeBEtflfvrUaIkMnTXsdz+FOevRTT3neURQxfJH0e2nhGO6uvq7ZVnJ9P6q
mKOcaVBxonERmzmo/EsYoJUSRjtSV0H76Y16fmn1XTB8T+JV7e+p7t57JsmXVmxs
wDSRXWDxDRZQ4o5Z9CA+A5gj5DQkmIPQMpU6KgscTB2iT2sGfHeqJrrVa3C7cECC
R9Jt0H4VmIioMF9RUYeu5FP0c2rXiz6YvJgt4tq3XKuFPqyQWo9HsMB3sHnGSGIH
7pvtt+d/eMLsh2Ajd1Ky9/DiByKSNx4z/n5Ids91TDKb5DOmpzyluCH37mCnHSVK
m6/q/oiWOaEMKc7Pz6u+tHxaEsX9qi/lZvFRGXZ/et4PBGyqgS/QCEjn/6syTbUg
OVYyiAMaB0+xmoDZAeqqStl1Pdzl8Zpg8dPjOWlbHKNtA65pdvzmpqCTfgDuC6BE
KjkkPRSiYPjpZJh6t+ifrhnSFebVRpFvFwYkx2JaP4AaS87leFdMv6ymfk2prjXz
7qD70qwXrouGpTemPOMEB8xnnhxOO5dVJ+YRvlk5FzIzigpfK4cGuH5vlZ8kAwkS
v1zUQHoW6b5g0lo+Gq5jv9BybNCmeIv6CCWomdIG0jVkfpgCqauUyVFlV4vijMnQ
5JCxCtZoO0zEd3B4HzftSumta9qBQpLnXFYP4MtKc7tSEhpwjy5T99/YZWaYPo+b
h1mHbbIBkRxduBqAbYALNmXuckmhJXK/vbbXFK/67v6YFP7lmJ8jc4/UduObWYb8
7LZEDFifRVJnw9CNESE9qUB1/Uxupc0o34g9Hbh6Ajy3YnVCEytiMekr2iBP+ptk
GAzdB51w59h6dqur59o+23jMLWOFiIhZOFR5AOy+f/YO0avrFLWFhjwQf+0uXva+
yYxGplmtg9YyWVcf2ow6DoNKef1xY42uske+65BxQhVz9HkhyqT4h25AngfEDvP6
OwGYu6xzKky+C4ZuQK81o1v/7IMQX1XiAfzcivblrhlYoHYvJnCPpLMoB4VVM4Bc
8t7AsGiFXorJ5LOMsnUo77aRatibbn+nwBJ5P6UnnYe6OATwpivZ5jVdi+0j8xKo
3b+6xArNO4tmFLmi0/zn6IyweEY6oUEvo5JZ8pTgxNa5caZ/PFSyCDBMPQ5JUuM3
j3L7hRkGGuu24XWpiT7rqfOvZPmvnQ19XdvE4bqZ5ptkPFBCtLKQqjWZnC/0+kta
dGo3tA7gU8Bz6rMoszMIOXEwdJxNgaKJnKwapTWal91PEBjullNmaK0a+3GB0vxl
cAz5lzbtZB/Yr6aGMw3buJuLFThYRR7NQS6Ife19lVdSku3Ena3D8fkhOiLRwseW
A7ilyY3ucRBfadAjHH2g6kw1NncUWSfudurybYg0AHzrAS65KB9biX5rjpsAOCIc
tWsKl9lqBCBcoBd0T0JLQfR4WRsISMOYOR5MbQWIgvacvMNy85vMGI/PhgGU++N8
wczWAueBXd7kJjAEeECEgkvPY6Rk+CV1ih5dLLqX+r5hOlRe2WQQaxEoQqZ5twja
RuOzCRmlD8NXNOQiSvzFiwZmbV78yaqmD0iInnx+ngagdcvR7QqWULgqzS4yUwa3
GdPsi+XmqnDVIZt/zdluae5khk5a/YW5wfoLNdG5jnfPhdF9bjQkpNFhAEuNC8rR
d/L/6rvuDS7exgEH0gokvPNqTpOO1aewF3PtdfNdHKo1h2kzjo+Hp9fAX6QPvAc8
mB/HefBQuygLFX47Ump4mmWfqL0bcFD9VHw3Cz5X/O4OjN6s9BYIJ3rU7/3CcYCO
CrsSE/7lNcJqMLnDJLZdYppsE4tzJPGBUl1+d2WRPGLAQ8ugPt4Q+sMPQ3V86KkW
OIOQM+wplH+FGkSbUFXDP6bJ5/Fz3Z3QcEF/xGFts7ACEBLgUSuVhk0MAiNvi6Of
tShOD9u+qNHkrTYOhjfHsFjha3zPoZ7lTLskixiyB0HPpLlfxS9rJWRvIn/xuxON
Z2S29ZRITS7gJMwkHA37zF+yYZApr/GnfXlA14culnqn34whkuWGxRHgPBXuu+yM
zxlqMQlEN8IktRsSh1NWQHe9qGx9aNbFR00siWNgW3M9dOk4h5XN82/LyWLli1iT
8J+CuBjSLU2OL8S1gih3nq8g7D6BvPN/uqdXPAvyNvgj79F69zn6Fk0w4OsoAGDp
2ghVBXR6BxMGyNRTSobnC+JKbhw8qgWXGdGerj6veMwXdvcQGBB6wGOCIEpFj7I1
BY6+f/kkX4qsF/TQ5xtXYPeC2xd+Ohl3wZLMfot61C8Ilw+zTTzSMmt1oa6aHfSA
Ggh+BtUwi/5vT4wKmN6oHQXEUDr5nhgKF0Vtj7Pv3hRq2hV1SNCwVO6nF+pD+IWu
AFEKASLexmn7JOPZAZFt7ooEkPAjPfp+WRbaR1aprOoWExSACkUIM4aW0y1Tl+vz
+QKrxWEAY9Q12MdY8tiPU+ptRQaBvQPxMjiYT04tc2+tiY6Wcyk1eErJPRMXJfor
EQ2aGPH5pXm1gSY0TIRwcy+CCVAuFExbjA01u8Ta3uyXq5zqY/5L0S16Hlt3uITW
7OnMj3L/0MS97CKutWwf6dWisS/5x/WlDuR/7j6UofPv/s3LbSFSyKbN3Km1Blzj
1szOANayHpU5nZg7TtaGqn/HctG3pHUten+7qHXoo1rGJivOXTi6Y6TKx0Yf/4BK
Vyku9lFxHAGuc0mibKXDBlGQi9xR0MJwgPuS46hraGT5TmdDR+QZYy8cjo3kukSF
TD+cZWK0vBerG+PVPwSzxeEH5DZEioidOJJahc55hd635jtiv0gwtRTkXvSHWzBn
QEqWtQlv06InVdl+O13CcsGY60guc4dwMijKQmFJ3gtdTfHtKhiLv6cC7f+kd8v3
5QZ4F8ExsNotxQioE3fbrbzTehr8QQyrm54RaP0LvmiYHPf3PxTEmB08iy3wT5uK
oz4Hv4/HzomiudpA9Ac84cFIz+TLPOuM1QYJpmg2hE7B6Gv9c7n7SDzG5IsspGDY
Oq/XdDQop2OMh208UbnlsRuyioahGcTRZrhBWqbxudAhqy1ZKvwgtvLTVGHiC7kf
m/j/WS2wC2oAKwckMUV4OIV9brUudYM0xEkI+5mGhTNQGcTsDdEiWUe9D1TZVIKB
EytK9UBGvCOIPKWL+lUyN8oNnZCl7mFrjSIvatG3RanFrmca7fWwfuY4lDysfJHP
phr76K9EIkzAVBjLSq4vPgLgXQgL7ldWHi0ZGa2KCXYW42EVydisvlkCSnDYAGUb
TA4G9tQHbVmDhYwUZkoQF2ApzFmkg77oldcwsoHEw1L/77UsDvATLm4tEDEMyuIA
i39L2Df2Of/kCuS8OxJbIBxzU2hlsKWeLokrv/5cpJjSbPINOiuATXsSoBpU+tSU
j6RGI4Q9Otbn/vOYrNO0TVCKXHVQb/4/3itP3U0XfobmReDY2hFZ0rVPHCAwdyJZ
v03Gz3ag66GG/8D+M09ok9b6Tdv+CICEe+UYYdF43lg=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HRwvKvP0Iyw8inu8XypzN0PB/j+Xy11wXJhDeEME2VxdUwgNj00A8Owen8yGmjs0
FBL0GE6MAMCkiAJOWBc+HleWjieTaelek9n2x2kssNp3i0KZLrGVMjBeFsMlDSKc
jQ8k/7WXRy4MPmRjYx7dr426tOKtgZyHkUH9Iqa5dRnjANYNagyTzpI0bfmhjvni
d7Uc4btjFJFTcaISLZV+l0ujALktSjgy1Ipac+rg1YoXjQM7NTpT8HjizY4Lhbcm
WyjREXXPa9F8iYToYO/rYOSOog5MiGY7EXubVJJ2oLTmNpHynaZg/BitEZczYaWM
nQvmI21PlUiMtzDsQv8n8A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8928 )
`pragma protect data_block
cDqNIyWdRbaFn3VqLvREZwNH6EDDLXpkSgYp7lrmpvCWJeck+JBEkyf4s5TkX+n3
Yp4V4AaVIZ65lHI7gOgUIsrLlAcpcYOxzbU2lviejIoEwmm/PaDsUjuoMW19MBUn
An4hHptj9DzsqoY7FlNZqIIzoRY4NaJ1w1kXIcz3jb1iRly/sbGkuF1jkj87b7pg
VRquyaRzXmjo77vVbHDlBZZUImgJ1NoMzm/HxKBjIUNAQLRyL2gG6pKpFwxFr0Dh
zKtnXwDF+SzprXdmfD1oqJRnl0pxChapRJJKAqu4Nmad57R5M/MyLV14/OpdNTQ1
v/c9tj3rPWWuHk1CTD61edZTR0w29Kmb98fV3fMRbkO1H5y28yOKEzXNI1c1/SK1
N9j49xPM7FDF9fwT4TYPKD+EGFm04mdchuDbx5e+v2+FjiRxIu4RrKgm9+jYgMPi
LSYo6VbukJ5okvGN69wYdBQnl5OPeWggCNvQUBZroPX7XuA6iEB3vKrVbznlbX75
6QiVm0eamXk/33u2/TSvVIsSLZHK9PSfbvuoUfoxab8WyQ9yHlunoEZQ+Z6GBRwR
aQoLLQlffH3QTePd7X6iT1gxmguC5VUGYezYTYg1ryfNZn1LQxnw9KRnL3+f/g5c
gQ516KwGYlGHlTkQ33v3AKNWQtdcEsaQ+eHW9H2rSiDahQapKo2DE89NYruxGtgh
psAcvKRvBiqtAkdQOlH/JuEI5LY0yfU72N28ZqIn68hUFWkvdxFQqWmf0tINeyRq
srtqFe6D6KHUXbKpQuymL9NGOUFGyuDW31kvIxDu0ovHJaFeNC9Tu4tT6UcyVy2a
Z/p0BBJ0OcIcwGH2ReLQvQV1o1UdQxtRud2EZHFLcJ+JUE++2ks9QTg2olt4J2W1
vGQrivlDrooc0rfWTnAdMhtQz7YH7F9fR1R8tLTC4IwAYsACIV4DQI0xRycKs97q
4AZgc9xVAyGdUkYY3YnaB4hJ4FkhHQqu2PY85AWlXjR/hiYdCSi5B5Bhg3nfYJPE
CA10aVB+wYx9pTA+AVODT5sO7Z/k7RZHLQ/qP5R+8a0H57OAn+cvBQHD1Y6gVXPE
S7rNtKPPjI7gjh8JpfmgcjoK62QFL6ligLQN2mF1NVN0vIqgI1uDnOYFccSMNgSj
QO38cjnumGxXSKVHHiRV3/OsjqgCuZwUThvNx5FJZcoctt6IdnhGHKSgX06Nzmj6
nHrDqKx9DKrdhGVv+KBLCo40FDSzPZAsgd4XB9M4dF2CrX6npLKTzdzEl0oW3ok5
ovJ9ChG58eNbHcKIqpu7pEnn8Wu2PQDhOPYzT3XekocKVaGFE7xMNU93swdbZ7JM
ux0r3repbyeSmyidbzwtdywSGw9rEyG/Tant+IMHI/aZRAX/0sdLlwaE4fJtLi70
5aLB1UWk1RvEdU8rn3f+hQXbvMbUKuGTGJU0ob698YPZZMCWPCu4PRFG6hST8zGB
MaKjdPEFBczHst5st56PNIE+ueslmLA4M7wZwO9T1IkRtj0Bnz+Sr833A/gztGqp
5TvkQfkV1SrfzvDM4lNlW+4vwSqeGOydF/JbyQ+Q3VK/61r+w1wQD6zFN7Ldrave
NJqeOZp77371cgcDkpDctZo9DP9i0kodqCxFBEYZtxgmaYq2kpG3skzs3V03xfx7
k9SVvib63NaomHM4xhSlPqmqOgy96jvyOINq7eVfw3WcooJ6No6Kn9EdgGKMnaxT
h70AEi7/wjbY7OMWxXZ+XGS4ElUcGGinemx5Gq0ue46T+DMOquTUg4iby+9A69ut
qa2QEqXAjCfnd1wScq4x/7/nNYcQweUr+FTrsBVKrpxp9LkqGVd9Upm+uJcZ8TiD
lDJL/S3hb4Ybvzk4KFCArshxFk2dZPY/eUowJFGjiFa4oEOuF2Zvp3C9Bn4o1g+q
EZFCylZF9VySo6c1Epjyq1RX4amvRaN7Mt3zkysspHEDYz0ndfelp+Sjq8a7DHb0
oM9UNEYfWySBWA/oPdZLLKY7UeSD9SQ4jKPqkl3v0ZUgqrwN3bGNvMtHBlHS3mLe
BFLlCITYcZeZzZ4UWxU9JNhMjMmsKPzOr+pdfn9fdZlrytnPtZZgckdqcUkJrqLl
pVY5WuxgumBoXFuerDHi9R8WykguYpjgwr/gNerG8KiFILEt6wFhEwtG7QVa80ao
nm74affYi/Vs3IGjPY+o4JUXwTjBTMJN9WI61oB69n2t5GI1nOw1Gk+mIBTiIiWC
tcyylnfyqV5cJCF41xw+yeGPIHdnCTRUsuJZ/vH6E9q7NLdXskx599KkpuY9j7Bm
mB40xQeNj1P8Oic6nyM6P22tmHXT2v06lGrgWbWyreMyf8s54mW9q8Mpvoq8ptsB
inOCZ6Ch9nqacCT45g2RafIEMGWXeM0N3Bk6k6C+nggsxnVmOlaghqLnresf/g3O
fMYxV7DyhBTPcxZJ2aRmsOzhnVTf3AUaw0csqBxnOzdCqM7FOXdLFjIKLNrQzwiE
j1MsdBdpKGIStTkptKgOCvIUn/RXWq64oj2jcJT2KBml/woLiEVUYNs1WTnQ8m8V
hxV6aAbUdod4tc+f2F6a22tKH85Hmmxzd4zWJA1u7xh50QI+wwVw2H/ua+sccZug
DyUs50UBTwcde0f2h6u2mCz/u7YPZY/Mg70ggk67lmyPjLofMhQQ8V3rmSJKv59h
aSLvZJlG+bLCsMOyVlwLwLRXQDflIldCQ7j/8VqDFQMfVvE4VtEAgy4OeV1NQah6
9uwKvnKXgC9g5ZQT62Mxim/f+F2lpLRbkCuNUEOUCutSgMF49N/tQCVesmjDkDGz
lXsPYYTGNMsZj9nr6zbNxszj0SV+dyi2BZa0/40IhPNK8KEYLTqQG7FpzYgjFmLh
6//pYJjOqqgYHNj0Or4AIJ5Wsh2CtROjiv1T1UmdolimSKXcCi/EJM4Hy6jZzxuE
UMVDb+/hIB5aQZOBL1LzkHHpeGp9DE9fuxZ7T3IwKtXeVZQ8dUFH6GZc22DJ2cjw
/6oZGKadu1tyrZGagrgXCuQUNGjieTHxFJEmT8xvU12o6xz9CJ2AC3mtFniVW6jK
EB2Cf48AxVnUsgeHY1rgTn7JM6djRQB8YDwuIkSlXvfE7U149a8jHTlqTkaRV5Kf
JZwHSQgz4x2AKvgKCm4HPgnVLfEUAtW2jSQv+r4O2toeOL1nw01l2bNnQO/iIHdc
mKcJlYGXwzaYEsvKMGEGw/ykY1dVpaVgw40UPpDCMKvyLxbhRCVME+mvon2yz8td
3WJVbbBrjTUAgNTkLC3qh2ZeSehSSpuqtjCdlSW6mzuOUmmCEIT5DjD+RqK+KFdo
pPDSW5dVO/+bfGLvSYUWCj5A2vJfOLixeVMn0ujjwuLp56PwzGzF7Lp5ruVkneZ+
ZoXL7s9YjYVgv7WmGYEtDb3ha85dqq2SyvOWxAe1r9coftnhzWxPzcbnJjqcv90B
M2/2+143ytpcz4o7P6RTLSCkJgy+if+RklrpATIuZlGpub6Gh3I8rc657A9fm8yj
h18sW4BJdJMRgmRr5fF116vZh6TgsQYIS0E+5gSzPMv/6bKbzP5rlCWYF9nFQm8V
HRcHmDAgdElRUa9zwbOSENPdH+ay1Goa2Nm97AF/Rd76OUK9NnIcNr78HKp1qU4R
27suoN8QzhHYni3ClI+5EmGupAgY/VP6NE+9G/lb1zueEfeVwft0n81ytwRYlRfJ
iEs1oJcxDOurbXaZ8JPSvzq+UVRXSaXI6G0jGMO+DJ+Irj7C6OfdZ0BrBmBkkJhi
LyeqcUaNZvxeoK5lEfQ5Ez18MOZJjV0OpApg8Xin0wiy8ZF0cBcgLeETvPLttTTu
oeAi5+JQPw5nfujmZeZdNVt2GgShWhba2EP8WnXREfGc2STyTRwvqIkwOnrCxeFJ
1led3Lsil+Kb1baWQFEodduR5SCXtLUwMorrDtncDT0qXSKWb8YCy0LKKuppIjET
52Y+Z6l6q6P5YymPDwKAOb/yleq5kHNzyI9pLtgmaLB+txm7Ruh9Kb/Cq4/0ziUU
eVQemmiUjrgt90QqYSvYL1LTpQVkB9NFheBb7U0w9bfVmILznd/NVKp2usQ0qA5R
YwBvY6e9cKBmWJqlkP+8FCPajYLlwTVB7PzW+BXZE1+LzTKQaIMomK8O9jiT0aaL
UamYvE4V1qudeZdSDBpTsoMwpN7J2HlCUYRlnWCCz0UfBaWAVg/tbcj7QNYHT7Du
qxSrZ1RjHMwW1X+LSxVXZ8cWmGFOcPWMrYRa7bd4yXlZ2jHQMmfcvVV5WbUHEbc0
eUpNn+cZkIg3/J41+iKRf5hHEtaD5JpGUtgePwY+nR7hNnRWNy/FasFRKG+CgbWW
Dh17JCTN0AfYKaoIFOtMm3ME6wa9NtSWweLZqxBZ466lc8HWWuE72vjoIeDJzXfd
phouRPdKdqdGlwix+zqhKbZBVA6SZSHrQuVT3wGKKCDAD7+eJY4iNKPBv75l0fzA
7rcILpuy+uStg4r90i/Rtnd2LPJ5C53gQotfXozRlRBGuzycxRIECyX19pbl3iTz
YpwC46A9CKqYGpTxYkLgxTXimp7nF1Fo//6BFNaHbbjSijIyxkfy6aP0zqjNzI1+
CXs/sd0/W41fKOCNo3QYmkvTwBocrGofVXg2c+7BEk7OqyFvswhWemW7ApMagkUP
SECepg79LuHiZJoK4aJ+24nr9UsOWyY8u7F4cfg2aPcr860E6RGuL2d49F3KWW8g
/yY8RQSKJwosFB7HvilCtiCXYWfY6sn3OYFmgzkqm7ze08FiW8GwTuZWSQo0N+CJ
k04RhvozgLHchGtdJp3ZNt9PVvFJNAPZGVA9Pk0OcY+DhbRQh3qXG0vWB5ERHFsS
npRIEMjwnRJZYaS3OROvM4WUaWIwBYxNTc7S+TGj/Q8E+7nt/7Is8ytpm4GK18Ty
YGLaN5ThaQb3jCXoc1MGazN/AXB3uKiQr0wWkXgJTy1CcMaWk86GxmBNEOiTuHEU
udQEwxvEeMtNrs0NGKxAsNyB3dbAmHhT3fFgIpJYJQdCL8b7GM3fy2scFZraz4Ub
aiv4Bi8SX1FbKz7PgSSmAe7M+RUQhlB9u99M6KEUVNTF7OmkBhuqPeFoiJuseqh5
In4D2l2fLARYCFwiCXretYYsYcenamRT/7ZEqNoIWQUO8a+Vhmc7JS0y/H6jO/xk
NN7RqStpkqDXMQ4a1obvoa0fRT6Yi6IbjVWg4P44SiIG+Jpi5kuHDoyMLcd/u+tW
Imz7c5+qWtOaJz87YMh1E1B868Iz4HMa3H3Aepur20/i/3SpS+9eOErE4e1M84VL
MzBCFap3YVvHINk+UiM4gdmk61O/aNVM7LkUKcNag7Dn+iYd4aWCe2m8de/YL9HF
OtbEGyhOWNzU6/+JdMAxgL0KdKGPYHoEhx/wk/YjEXrBsUgXVdRYduVRmLX8P+AD
ebjPG5S/OhAp4Orowi05u4T+4pDnBC1Zv1+uP5yTFv+InuGwyucY5Q2r+C6NONhk
t2XLMPLCv+rO9G8wVwGrWkdrlxfCgRyzzkW0H7K1i7bWdnHMAgQBgny8y/6Wt+ea
rGxRtcfLakGltm3mARKKUdFDzSvKxzA8qtvg5CVc6hIHQi4kIkEGbeLRMzuE7ysM
dDER6ug41IoTwOTWLGqbYVxSDSQwGdSBIcprXA/Z0sSpMCQNFOwbjKjFK7ier5Y2
QuDq6MHV9S2qg2PdHN6lz2KQIAKPpF9HjeUDpbP5Fe4lG3TJ2UsGG08jmvXpUs/a
gfW1E3DvBb4+6f7dGDrYJf/rHBVoBHueyLH8WugrcuDVnyosBNyI7NgXQpDyJ1xd
yQEogy9oMD3rTXulxDQ4f7oLdS7DRuwtHy5i/7bxsy68fjQBy9bcDBgP/roki+Qz
2UDTs2SKO+T/uT0IPTxeEUMAva1h0el1GUSdnInswjz0e4jSHSKw38G3xfP9Rb8K
9MzR1uSCzJI/D5HRZ3MiMpsA6lkINZJGJHQcQR02DeCLBoFKL+stXTPp6Qlxv0C2
62EeFPHk7r++uI/Iz3bv93agoMPg+4z65wQhEHP+Czu4+8EtSdw3tfiJhY7xGh5N
+HUyJVdGaRcfUoIufvbsvW2GpePGMPqrgv6NpNoCr8bp4EX9k6OM8POH1+gcyQrt
GEVnih7L9irUn/3g2uVZqw8XPQGqi0xm9TUcXoeqkB6eVBIJLV9xyIbPPAEZHO3S
VjXKMzQEgYkjA6zmrOOqrXP2naPztMJZvQ/6zaI1/AXknNI5Wbabc2ohUiaDZkMQ
EiVs+jN2PIW/luEyOUsduruFYUnwiyA8nfWdsyFa0fBgLjm6u1yM/+HrTKwdZBVi
lKZiQlY5FOQRfKjw/g1yPkT3uy6AP3b7qp1mY3gJ81UDPUvdH4Umrxa2YKhdrACh
GiLj/f1A8OD+Ubjnd/Byku/20a0zqx9CmzFDPMvthDEE/Zph5xff6L0Gv+jxuiWO
c8Kn/7d7z97OMY5YYHMGMDvEUWR3bFi3P18jZzz4hmcGpIWjCzU9Uj+sYYW8J2fz
z/nJmCJeESmJ01cQ7iyXizwN1/EdA6UFStaCRUUE3dwE7g2uDjp39XfPMm1wLt/Z
4tR1MWHvzLMsX7D3wsh9wzjd197kmXG9dcv+v6nicQWieR4ErW/SZtMc26xVokt1
SfFfQ5OgGrW1FzNRTxuysWWinoTTONT02bPsJTiZgCuRx6GEY3b3e7N4SoYcnr4R
0RiYEnFhGLJdnU+LM4tfmgpc0fJ8TyuvLq7NUMLzFhJzdVUdvbsyPfIcFgkLnekE
8M8lLWD7wtj3WW9v0SnxcRWguIy54cjDUf24/50glGncofz0MbSDrkM9v/vSFEYa
ikImTK/C9n0YUG2F55BKEdAIAdUv7sUha9beWn74xyGxnP2oE7ZbMGkWvXv83xdT
kWFFmZQm+ouAu2tuUMQqbwvNz825sBA21ff9uywDTz4myV23vC/l7ANb26rQQXhj
C2AGqXqLLsnCK9kAcwx5HLMijFxRp73sIwoNSWxHDhijcn6PzC9JfrV4M7jR/6CI
HgVoOsbbhHuPAfyNluGcBv3clse7tVAbH1V3cmOSx8UEf2w2sBs1ptuVW0Z42Ah2
QCN5mqY4VuZF5rE2QmHYq1BRT7Yav5PuTBQgdYZ9LDcqsTWVgLzVwbUYonlMJrUI
rUsJw+SgWFemL78OWlPBWpGPffaeV4/j0vBK08XsJVeFWI1jxQ3kkiWySpvZa79P
6mSEX8esSdv1QXINSuvv/NdAicHOTa4wejIIkAqMwq8VM9Th8Wk/p5cE0EI/h7BK
14z/QCPPbouPn1pwU2y8c8f44iFn1EUYlgD8PFWM0d3PPui2AyUmawVWx7LpoTLQ
ROFHN3jgBQ5302RZ61/iI2Y9lB10k5BEwmYBjbBMvSpSDS1T8XHU50B50Ch3G60y
4iWnQTGREtxgg0Vb5RYah99ZzxrGj4F77ALYiSV/4d4By+ttjCvtTaKbFQOXD6Xk
9/6Kjx1NIgD0mTbhHSic86YROsM+MofaahrfxrgKx9Xrba/IpcHaY18Kh9fGjLqn
WG3+ejosuSDtJHU3LkuKaQsQ1YAz/QGS/WS/rlFMa0HTggBn68J5dJAaIPADvKt2
a3xyHnGbBGJdfyfb9VeTcyDA9CE7KVNZxKM9YYHdSXvXXdsxwdram5JzNXT9J366
wFgPEISIBa7ak0DSdMGoYDTSxK7d62agwgFmVHaLTy5LVpd48Lyl8rcX2PvSkI79
AAyWoDqIEjje/5lMk9/gIHcTEx25jAVBpODQPfX9onsIvREraT/J6IQFj9xfjzHP
T57LYA+L3dxgC//4z0GUZ54IR27hFNZlhp+d+IiaOBvHRXwOUwRDLu5i2la3nCtp
l+/nEJJKaQ7TkUNIyBr9KZUVtk+wnJOnlGQLnPswq0jYkUu+sV5N9gEK9N+L/Np7
RLdzlYEUmT1ncnUk+QYkPStUICEm1Z3VbkHcGOMgc/jrY9Xlk0guTFTt77PFb9Tt
BymgpNPKlCWTd/ljmBJ3jgM9YXnQsYrPGvVHMkyrmuxLFg7N+P9hugFjJm5jjRxr
eP+Mhiiw9h2Zm8bJdmn5nTaVOKaWdA/FLPM1dT9L2GKiN4Dm6cWQ16J79RcXry1S
IYCqAGnVjLZtgegPQbIJyFqDK7p3744tYaq7yikkBPfzOcX147Qu2VFCUxKDlCpa
YW5U8zO5e/maBkXwXaVz4tSK8oq1IBJip3upQ/db4fp/OkrxEpBkByie3SMV8arz
iBEGukYrJG3UG0VWqLGQG6PbRj2bHBxtA8mv0Fv/212aomhBufVHCNeXm4tiO+3A
K+P8hxwrk+2+3YRWtZs2DroEUdgmSW1gro0Bs5yGa7k5VQafBKfCYZPC9/R0H7TW
ehwh/Q9Obss6F4xiCVgkhDSpmDSgUtOdrJSThlwutHiznOQfSkhrEI7NS8vEq+TG
q6EBvSK1d2GSyx3vAQIBWrx4K1N2CTsf/dD39r+s+egHlbqg0n0gUPW4q9JLk+6L
8kZvQFgK4H3ZUfnC1pQ9PJT2zHJVvTZLFROSpD4Mhl8Mwu5Skoqav3SCyR7h5Pr2
GKs/JQbJ+dsFR1YUyC2/aVD0+RgbQsYRq89rzuAmUEfAo50yV4plMKkuzB7FYGWT
ycn9xwaAsXCwFzs1CHC5hjakW6pLQcjr6bft1vTz5/v2yE8mAjUFT/3Ts/9tIYcu
ib2LrvSQVn2pPFmF6wtNlfJdnvCrq7jH0rmEynau0JWyRvrj8zqaZXUhgOry7tiD
lVD512vWrFgg/JGyee/ZYgAgYtGtGT4pBoaVHBhO4kA01XyQGG4/kseFiNbA95dd
WecGAvchq+x5C3HslUUDXlcCnaP7t0x9Ua7KsPeC1Ts+bXIqYNP6GQlt5ByDo1Os
m3ALWwwnQIb+i9Ndv8JwJgJWwpWwWR5OY98uJP1FgeURXHNUIs4vVGFaF1KvVoQO
kGCTDWdjrI+bCyRkkU5e4B0QCemEdpC8A4op4tkkuOAaO7FrEsW2ot4092gDc7u1
QE2ilpOLSO1RFZ4ltWjlHDf76RJytg7WnRueCmIlz72bbhw/UNQm6Psw4KpHrR9o
KPLk/o82WHdnGpi0sgABLHja39o8/5EwUgxFQmli2RHtAWOF1KgdO+nyegco3ZG3
kwJH5kGVYz+QuCID2+iHUInM+yLVhdHFPKdHWDKlFS6hxih0tyqJO/9opZkXADhz
NTYgVgc2f/cb9zHCc81oUvoYfdpBgN8GkJ4raQPJeqZ5WGCDVvDtS2M1XgzNycxf
zCGdXsBMnuNhLq7kXvjtK5pT5n3gz5r/vjE3JUZYSYKB1d3je0TVjZt9/YcBBfRg
8aAEso4pW8gSsxYjYOwY8xCu0QG6xQGmzNh1oVe8QomcHe5LUiItU7Egar+o/ueB
F4nhdXgC4e7bWWZV9LWZCWl9qLzByAoWXknM7K8sl/UCrWhMFiakCsUgC6vCevtN
xegZokUZSmuXqpOw+cnYFUy5aN7CWumZrTt2Fryem30WQPMTMwqYeaF5PC6Qnwk7
0KAae3nM3niP5h4O/MuoDcsNhMoKtWWttxQh8cCZrKjsk67sf/T2UcSinm92byjA
GtrCRGt3VNPrYAvKzR7Omq+xs2s9Ibn3ycNf4Gi7p8gywYNFggFJSlU7EZZV4ZJC
mF/HS5auqUHEoerkx16X7g9coVGiT9ZLEBUzlJPZ4Gb+KAfv1nOOVYnTQqkeAvh9
TFwCKcFC10ady2ZwCEwVpPbUkXGAx2uOFatfATmUFiUdXtDrwy1ODwTrKl/bE3+9
kajpODMM/gCqutls1TZcL59mhc1dhdGTof3IejQhbcIm34AJ0Kzz/T6dwBRIw8ci
ybSVm3v9KlSUnU2CMibD59xPftVTobc/+7xzOWPKBqhuhwtD4qULkSqcjIGRqKP2
wbuZMaZ7m2aQcX9xmNewFI28p9Wut59Keq3BR3c026IdEwXu7tDbGrStmhP33ayZ
sBLnAYmjjzN5rz5/qXdA3P+EoF7tZkMWdCuXqx2gPN3jCKwAyqOTfrpB68L2VHnW
KrCfRGTob2LITq34/vfSxJVabPQ4xOBucGgfo84GQ0jhTjdWfOqtImQZL9EcJ0eK
1FJcgqKuczF1+TczoEXRWjhjV43LsXRekx1p3VpHqcyIuS/BozYqidZVVKRzmXrl
SdPzvwCMzaJYirwvlIPwBInMYLYEi9NPQPPl0SKYlIP3lKjkDYkKuSJiC5gFINJT
EsUvPPcdRP2yTye5k+iwMlWIdS7SVUyM67zCs8r41WZaJZ7audpC6+f6iBaX/QOA
A9MGrGFtUq1TCfvz52vW1D+QGbjeefaDZtkq+y337c8qRacnC5iOI7PZhAph04qB
Gk/O+N765pLH9ls/ldVw6Qpn0XZ8Ht4TAAgS+2AFLd5WAznvGKvh8a/HJk7xWmi/
j9PTtJ9iJT+Ki/ng/Cp1wSPCEZtWYdg3VMsCPBkrGJ3lBRaduYb48tDgDytKtgD7
H0ivZ6RinK2Lt8hsQlAAiHJXODA8ysJe7igpPtbRD9N5syloXu9IuVtnJm/wl4Dn
zQcYQbSeCYcNtFBxL+3OI1zmbgTWlifCN90WBOeXyxW3lLzVY61mPnBFOnPSNvNF
xIcI3AjpsOje4wz/DZk2HiQgJ8CUxSFUKpzrJlTSlxHalrC7LwwkOKwp5FyItSTn
UycaWKa+4JMq1DulWh+CTIR4Tf8JftT7lsQCTXZQApSOXy78k1udDhkdV3ZrGbmd
kYjn3wBKTmbxx0NF/4YeqKhZ+13kivkK1As9Srd/jr7l87QQoTSAeJlhTHx5Dh8J
1I4XTESgJlSQFpRvBjmK0IzsFhX+0RlPUTz4Y8TlMutoylOAHGvJa1nBCQU6x+Fi
8Yn3u0wURTRicpq1UPzr7IMwbPCUY/cLDJ98E0h5eqd+6Nf9KmSH0/eQTpjpOLd/
a2AHDKaNSr3CBdsWsmtsTY9OlZiHDQFOq2oAdunWt/p7tPKLa5m/ol0NY4u53BPB
r+7++J9T/yGmGgZvxcBXwDDwLK1wxAKMqgFxyGqoqa92W2hKL6MKjaaP6I6ISgeB
bOK0SsZR+y1KlWP30pSRn3vsOutNup4EWnQxsoivy9VPzhZ8kmcursumK/To0fxU
W3vb+uQd8W633NTqqIrxEXcwhVzA9QAZaqYL/MD3zbmYhAN2BsCr3xpnTJXEDgwn
ThkCC8Y8EhFbSGmjhvH9hTCpabKaMmI9PU5k8KMtS8L4AUKGq+7D8h6JowQB5x/o
lGKijxvn0cFbckeYdeDGFEe0CvwTurkDmTcvxtxQhGVhLohonJyNphuhIYi6ki7G
szuD7bqb7PJ8kXr2Yj0RhsMDXfP4bMmH/r418absoYOoxKZscdhMgrc5HAvzNUNN
tnDgRiklPqZQMvujE797Q4ybAtj7P87IwbNjzq7efsRoFIpxDWgv+70bygD7g6gT
uCTBduq3buoXTLXRD9JfvqiSWCf3K2OospJ+uYJUVwt6O5C2YyggYtcwbb3uWSBi
toXfbYTJ0Rpj2OB6S7+8xdKugQs1cXZYGG6TG51Q8Tgfm6+3Kk0YXlLzzQjIvuf3
1IkAg4dEzuAI2/q+bk+wzHEURFZIUw6Z65Y6HZNOOGvSuTQZ9Pou+B1WhNqR7egM
cEnI8PvJMhb7u0i6vtGMmdEUsbsr4QDDjqlBrog44UiB2G/tLiFdiQpnDQg+Pn0S
NC/VEydKITmot0/UjHWyumj77gkC0GZDrDRbi3RHPji9LDLXEQUVgfh50FIH9RTH
OijsMeOKpUcwB0jm+FUHulcbmbI7QuQLVwML6bIbkbGoKOH3bfGMKVg/dfZKFqos
W6MtJVavkwtWek9NfQsebhL2JETqXf62lLdrm2ifagGUCx4TNz7E5ZKaRz8FMmbD
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EZziChaigivdHdpctRsvO5+WHxKOFlIBE9Vbe45LrAfkHEBp84Y4KQdOPUz029HH
8c7OLPuRdz0ZTZVLREIQv/lKEiyAXnFfuh16tuvELE7DsIyF/+7g79G/OsXxG8VK
rSmk3sll+1vbAwCI9Xavc9pU7VF6gzY8dzjY0mWpf8OusBH58s0DJH+VcvRwpfUv
JyS6Bq63VVxGUG407lcPa6rK+UmeFIzbYrfhYlt8z7fz2bMegjXOYxFQmO9+oCjr
CdCm3GM5XHetRD0t0SqUgO+qGB7QtqFp9ubqDvQv1QcrlQxeeLgWxM/K+PqVTLuP
0GIjlRKoyEcE48Rs8Vktnw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2912 )
`pragma protect data_block
KKxSEX3RZ6zoCEO+Cm9ZReOkDOezWZWkMMHGaqA3OjwTErpTX565yZzBoUE6tJ59
ZMN9k5gKsJEignfd11ynBIbp4NaQCykYPjgxzDeZJGz94lmA/+PGqNONNZE6TNOV
ErwhgtA0QW69Hz+qBzrgQ/LigVEK9mOCSMlEchACwGQSW2YZJzROFFcjzrRCs3Rw
u3XJ8pEAxSE4SRb01OSkhyRXJ0uKOASahfPxCxm+dsuPlg8nDEA1Z/40ZXGhwt3H
dq5y+0+C9cFLRWFZOmHtYtN+iuBu5MqxNrzuqWsvhGR/aqh4zaZqsEDvDwzXEQNQ
DqpaqmEIx9qzuviKX1RgrcIe2YQV9lJp6ElP31BFquUj7Z+utCWD5RSQJybzDrTj
lBvMAweoTMAVzOnbbNBHPWx8JJxWjiHxLxxea3SXlZhGTcIkmU5jgXQ9hDiLlMnk
VamMxmXJvWw4ekVH+b3tqWOqpHf43wiIe4aDAG9exkgvRaaO4BJNNdcaMl+jwznO
/vuww31I4jHV145F/WP710gR0Go10dT8LfmlQCweddHCZ697/QdyZA8eDo0L1tRv
DOb2gR4k7UqmzkIa78uDNR4tQMgZdK4I5Icnd2W5TTZP6++DPT/DjuqldPdEeetO
gIzjf5dYuPrJOefpHhLjhUB9ixSGchs8qMJSEu5KDO1VtRNcET9M8KwtmjzN9dE3
43c8ihuxF13AGScT8zz1djUI7DAya1X6lRHzWIksWFrxOrbmBWhIXbozk2sS0ayy
0QNq7jdmeH4OcuQUVNDeEOpxsFP04tW/V7+XzpxnynD4A8/6+QYx/hpfH88ldGCn
leQB9BCAe2OnIqCojopQsesHbu3N/VB9CkFF4iSe88b8Pku0vmBUJJGhqtAoWW1G
4DLTIk8NTWNm20moElZ2VQbuXDG3j8j23gEVlgArnbRHDggOZxJ2JQSaP69vR6YW
pr0WNCPMj2PafxhHKTJwsbbhU3vBva8yRTI55B1LNw+le9y7WoBarnR6U5D2U+v2
Mv4yfOolTswxvIhx7QCXN3kFp9z3+DdPwcIJDmSBL3xlt6yaoQ6ulKfwu9GHFfVW
SKr3cJhCTEuDTmrB6Qkod8c+OcKN33OUX9tt94M/3nG9sjFcwucHf8DG3sgf6OWX
dBp7as/v1UMtplBy7tsCQybcrIHAR7anmhVjPN4LbpSlAnLVtRsnrLwf/w8tH0oR
19BhwaqZkJZdeO6dRfO0kp4KXDu6jqM9btHmMgfnF2JxrUiYsRxqLMIPwU8iBInU
1zFfum6mFq+vQ2tUeTEvs357znlhKjVpoFIuqghLJZrBU/5bj58U8rtrAxPhY1gc
lXBOSBhWTwnKuavkHc36DtuwgOb+DTsvOs4X7DrBE3CqNEm9FSXe7vR3CJSCbKEo
wemFEq+3x2iDrf3OHWwQwjIy1tUxtDGRgqzNJvg8FZ6D3OjrtJyqo4ef1pEdG5RJ
WqyplUmKJEdRUAMLpm0uY4kXZiTPsBoMgnTmhZSWpYXMWLC7JsHoq/ixvUrL49ds
laLV1H2/OtNUXj2HDCPoW6tzns4pSi4APrp6wgLBYN0bD0bmqxBZ/ak6CMVoVqii
mWNQKGgfozrU3Y5je2I5QRqkY65nVWiDDB4YsggTuzq2Dx1ENgYWU7G0RDdE1HUy
qfSdOhRH5/Vxvq5va7DzBWMYllFkKlShSTX9OaMychTAailxOFumXDwdDvaXF1VA
3yMSIwC/9ClxgLBORpgzWj66jfGs6I9G6H17oBq1K8mJyhANp5Fi33NJ7SMudSNY
yFKa0DCuo61xaZwej6NrDpRzrk6ugO1tkn1BXWfGCXyLMCjBkGVHJNaxLm1EhOQI
9/V8HPJj6+NlcpM+1L2j/Cu21LVs7cGc6xG4lsOvFeG67/rrgOO+U3w+9Vjwk4iC
7tLHAdOSrgHIHYNjMp9lWuhZBUJDVKtyojqCYBMPXV3SSRyfrdIaljJSd3PMxg72
gAA4F9AqULd2cYbnpPN8mQw4gqFKhM7UYhcXY454FW8zPgYuzCWOsejkp5pjWOJd
RZqJy+MZb5T0p+7dXIAXGnQVBxxZ5C7+pRujnUNkfpV4USYyPp+DOhe36JxfuMt3
VAAYXYhQfE5xPpmEUnRd74nDPZjta2CD8c3o0jLc2ArZa+hs0HCM8fVIDfQ0kewl
8c4ThhfuAG+GhpxIjq4VrsAUP5P1l/vGwpffV88D1KcVPoSPIUHP6Hv2YY44eSNV
pQ1laxOPIbDjEyu4YGFtkCbw5D/yOCc/BUrxmYq1A9QvT8JBSXgX7AyiVyFUu50v
AXpRZVe9iGCfYmBInZtfaH9ahSx8zQqwiWehbQUKSTOCCvXeA3cUClLlCEypyNQu
eRnWGPoIXhBzBbWyipoXwYZazbKGRpjoqwVvdVLQw7LuIP0prnuq6NKrWCvmp14v
vdTN1gxWjanzGoSRm221rsxghcruD02u9aZ8a1LycJvLSH5tlYpUSUMZrLmC3ZGj
etAalVoXPTMk+R7ADLU4g6lnYsNu2CXrSV2VICIQGDcGOoOm4xtWx264oUILFWOC
jJoyZmH5hnc8Z3v9jlPt577U4cRcZhtS2L79wtIu2eOhY4H+yyr+AAt0aznfXtAH
Gm9CPmdFPVwckqLwXVPt3vKAg+YpvS0RFzFpuzwJQQiX1ONGuoyxowVvvctJI6Ef
kqa8Zqs/zjIthdNGUqOq1lvJx/ieAaNKy9ZcTsfPXVpLCgB8balfSoeJkCNnDNvG
rGB1gYZQuQj3LrQLJOCWwc8VrHQT5XYxNhfy4rZ4jVWOKP/85XFpmpIgO707nJZu
ZKJQ6cdl7rYfJ99Q7eRTc6uh55HswnYrWG7rKXrj1yJaUcLZNb2wlcejqyAF/7r8
Sb3LNlSM4vAhbT6wOb5COM+CXqslOkM/iap7n8zxsARQRuQHyzBAf3ksQH31Dit3
kk+/I46C+ndV0RMLU+Bdby9r7avtB0lpxeqJ/vtKb/IdhzqubWTP9Ll4EM23mKwo
AzhNAQ23ootNO3WtGXyKkwpcvgreT6qOPD3SirnHcvNkBVK4/ydcXW1hrPEqFz8Q
4FSfsTUEKjiXjwxq9/Iih6Es0X2HSl9/kaaJd8S6KsJcKjKQUuat60SimzPbf+XR
aAu8TPoca7JDpDgYerlNkwdiUf/UI9JRsgqXfCFUbFtwb2eFrT8lFOZK+e2XlHaS
w2AebBqeijJGHlF9upSPWv+yRZeNoyHjpdBfVuRTDZgROBv++FCAx0vBFpkPNE2E
XmeMTrXA378cBEknvs82J9FPOV9ZlnxY85oAH82a9oaYHTVmLDXpo9L96xyFsuRS
aADiTBrBEg579VlLXOpPRJEowYe2Qfy+WhLEhXeENg2/aOq40J2mwrz2XAV/5tDm
iWe4KLDjaKt/9C0enS+5Ge941pQxGygDEoPUKgBpc0hleULDXE2bz9eL7n5kOAgA
EF1DMakMQATgvMoVVFmLAqML+f7nJ4Ozugva9uqAFLBPTXjgoLC7xmZRmnlI1wBw
LI3BYm7TESFGb71QvRvpWPSzYijRNrP+V29h+buVZAWSin0ADfiQfbpm8Xw/Rauh
VYMBmuOcjI75o8JAVE/VaMUZMjFnwWiQnY54CPWCEQxiQTyjJgcIUKWUmRz4CxN3
+U9ePL6Q4PTvbBlKwLhpE6ocEJWohsqlBw63EDK/z1DzZzr1T2VQkbCscEFQzi+E
9wmlspakDrvHezAr9ZrJgZWOKzYcYCYyO5CgPMVPGIY/mIVWBj0vA4YHxPOus72B
WzoS8xMXsKx/44ZR+89+3ujChUoekApNQAF3AKga1pBTogwKiJPo1EzrJNSNLKDH
69QcfdoB9kU+PF3Wp+upbdiHJi4pBVUQLjg7rtrXpKE=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
iY4gumT3F1MUpMW4GZ/BYWLhwXxZ/uCiMtWRt+jYR0fBB34cDExKvQMuKO/CgwC5
4o6NN99hFloRg663YopG6wKlbULiacaaaLogo909/2Fx9z0V1VipWTzplzBwUokd
UX4yhmG1+s3OuGLg9S01B0iClJKyoxBQHu2TBx6iOr2mGKx0OvBiSWliQfgJE9ra
BB3BrG450gltL6J23MW4cwDdhtYEO/FSkVA8SUvhtw1bW3PSshX28DOT6/Jl0vFU
mTapZ0yc1owDnTG6fV12aVgbI8wMvuGDqmKJtNE4V9iI/zR7+IFLFSWglQ7HDcOg
3+lwuODL0eVgzJD9H5kJvQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8016 )
`pragma protect data_block
/KxKXfMgga8sJBJ5oFce0C6tRJ86LMaSWpw4dLQkXC2TngxiOdGgCqlwOfEdQ11i
CBlFutDTohjG9AkrIQmu3VlzZ8U32yMslWm+2s3CIaysMvDYrHjCxpp0DP+oxMK2
EeUnOuzTTxPUiutDwr0CsBYcXCNCAIlc6yK8m22SoCXT5vn0Ba7ucd2SwRwgGRMq
gZUdgzhV6Th3VEz0CVkC372v35pz/DmhB5s3pHrGPuJPK0xa/oUIgVJ0NF98JUm1
+JdDy6qhzwIgBkDIkvv4MotZs4lcwrOV6tCjHJyeIy0phXB94vwGTMXhQc8mQ2nU
N1rPLckoMWcnlUE/azkA2wigF1hRjMllispBSDJQ5XE2reVxJI2rWv4DMMo+undt
+R1EngLhyPnu0Du5T3uRewl11pBE1mFrtSdMH/vRUj5/lDYtn9krF3IRAF1SWdnL
ESmyvbk6UNgN0Abm9w4GX040pZVgHSkoDeBzVR31tk1XQv5aP/nUncHTX9drWXVZ
V6vgDi/NKzAJdPQJ1IbQgYdgTOXZSTYQU/R31QApZf3oF6tkhFQtoMAk24Ypm9cw
kxIzJ3goNot94Qj3jkCgDZzPPfQf8bQWar5+P4vBTMAR+cmjUdjffYj3MXnM8b8v
HprXV9XacydqDZWdHRAxUmt/eae04bEfcmlKW4YEd5Q89TANsrP3vBtnGU46BlEB
IPZPxi1RrwW/953EA2q2TXxxbUAWfwgrXxO436tgpMAKb5qxb45EjNQPBhdl9Mxu
JLBDo03jmR8LLKAAEldJKRAbHsp0A0dLEQO8o0sjvbitEc2GFV4KWYJKUh7YZxtA
RkXZTek5umeYlUHp+Eh0LSgYWaF+edMhrIvWbCY5eEs8MooZL14rZPSUj05lE8HB
BVBimrn2RPwKKo1dOmBOs/snHPlf0EbpwxtfxFG4/wpue392i15Gg8hHezltm1LI
4WcAH2uIfT4JHy3C9DO90MMyZmbWNPwhZkDYzwBGp4V6Y7383QaKNUbF6ZPxBTKB
UtLDvn8Lq7XuUh3iv6TswFZxVZdYQv08ymI5uvE5o/ncr7aLclEZO49gTrQ4p/pY
EQujIp9hQDMOkWYxgJ+yJCQSKLSOQpXq26sljXeRuM3pUNbx3UJFRpieBfNxZgib
2N+I3icUARaMtqoW3c721pT3IqQ00hqYOjJltUk8lRt6CwPBhmwbqUdKbFa9CZaz
sgcBAjFPUAiFreZ2EvIYB29ocAnKlSyggHZCSv7GZab/VGKbRg1VI8kCdTWRNx24
C9pVfQDiL9hzYz21JTtBeT2m46Fc4GBII6Z6jndlgKtP4EPf3/ejCM8B6o9P0ynG
z1L0jPMJ0qFAHtzpZfd1xJSUVYVBAHJ0T09sSa4Lr2FYSWac66J+0bt0uAyynVgn
MOpHdbZd3WW/NL5Oc4Gc5Uo8RUoM8+tPOD3aAnmNfz6FspanKiX9Z+gXNEP9ls1Q
HUW4AWcTkBNH/IASMTbWiZ/qCvGbA97PxFscUqfWfBmIckTWs6EP9ZN/Nyqp29WO
L9o4OAaZ9dAC5gFuCDasmWabLDnH4gRSHQq/hb0levm5A50vhfzRRO+hjmA8qJMK
CNHqAID1jL/1fMOlXVCWWFq5Hv3buHZy3CGb4w+KBZkEln6TQx2NHpHT542AFZuE
8jAh8ydDYfQWzXYSyDLWbMfs0DVDkPsPtVvGsUU9g5cs0vUvpYlkQqMJF4WDmYU6
nsBy4l8wRf2mHvOt1AJUShcTfpimPwmJoR4NPRAuunfoWhiFHCVuNkHMDg4dMPOS
0uduHcEZU3exWg/bXyjuF2FLr30D5tBGMZKWvs8DtKjpfNMJel/LuPPJEMfbtxO1
MvHRIDUeC8G7hqMG5kjZGp9o5xwelDZ5DVs99L0M2o5W6C9Q3EmNelU34jD87zgt
CUWNG4w7wOy/FJrlBqKGmH9QU/tEBQwdBZtMfuRtBsev5bW1528oJ6suI5CWn/eH
Sq2rEvLqaTHuKDimGgIAf+WxSLxDS6RtBh5GAi+bPbFeedtPJe+BHHHnN/rB5VqR
r7yjl2SqhUmqYjVv4icifD7RctPoaVMT/05gQI6bmr+W+0xM8yT2b+Z+gMVEb0Cu
50km5cL9fo+5PFDfwzqoXSHV6hu1OZlCn9fOpU9GhMKt1HmWyC3I19Noy/0w9ipV
MvZAOUtTHjc6CpeM9GilbbsL/wvwIjjyGmHw+sBqBJR6KEQBY/UVxsCLGmCbG3oJ
SWLVEjBTPxBpHRuRPB47USfzU/gv6+SOcIifx/os+hh0Z7Z3Y3y95hoA91b/NQI2
+62xAnsgpHMPl7gOxXV2RDPtvYVCkKmQyD4sA+DljyN5PqsPWF3HuUQa4hOa6lSh
AjIO6qh1pcgBn315raUhdRWNgeSrpS7vFiBTkYf8R/ydItYCFeDl5i6iRAL0KMBJ
Vksl/+NhxdBTqQpWIERNa++rxwOSx0ymOfcHi6m8xQyShclIQVxitDPNx7cFGzT/
dcTbi5sHTDbI0st/OOqYFZHTkSxBFZBEZfirxVcY/PgK6FFwsKXXlDvI+aNtOK5F
OAVCGRW2Mu4STZY7NsGF/FTSUmikutC3wj611Iq8gtkpyS1h/jNxQZozYLW+vXzk
/5xS4kvHgff5ldnH5c8YHUKBZIvjsFjtkJcLao+ZfTNrwl8kavmFW/rbInHme+R2
VD2Jawaqx+K2TlK1/R7zFQ3zW7DzGz0jNMHzeQxh9Z69Xw/6ueg8cv5OvrtI6+Vl
eXvcSoohRQ62MvJyxbOwkbhAlsukkkAUE+e1Bm+SALsV3uznRN6PBUXeP3Dd5d2U
ONiS7MVIlE/59nFxm6OrJrL1uSrIuf82WxuCO3m4Z5bSIAThMCcZRU2HYRaHbOVp
y4TFrxNYnSlqbQ02qIemj1SYeswHGL4//O86KrwY+aiqeDI9+DmhqHPh+P+zeCR9
/AKtK4pGjr4Bez3WRIN9ZcRvFNPZ+yi5/YfNmHdfnGQYEMnTptnnAryOo7yMRDJd
F482nxKHlAzGcmjUnMkpY8ukS/5bgXF+yDrMoJkxZ5eVb3fAsGgEhdNtfvVOysFj
O9oMlBhON9ZJIulLBwUlfqUaTcSEhRL+z+DyuMS0Ueo4gIm2bPAj6goVhGpaCdud
SxVDlyCsYO4unvG14nYvBRURhxY4z0toibMODPI2Rjh4JqjsCDjhHy3DmRprb886
zzjmJCIsrC7Y/iELzDZPxUbsW+g8wANgAtvg/ArtlAei2QVI226uy+nT7+UIRmt/
vBgEvdA0XDv1D2Z1BJCNJWSXcVeLmafyZtkMJG2aOB5D0LsGIq3kwmYy1k/Zwxs9
3VGFnQxegatMo22oSdpdGaUIUTrpPYNmP4+1FQ7eO4Km2lU0mfJdcgrcTWRiEay2
BORaDG0ZyrXgRMKyHpU0du0zxQp0D9cUKNra0iBUd9zaCLZJ1K1WL7evNx++1R5Q
r3GhkmnhO4zG0p+hfE+fJsIr/C3WgSjDWq3tf3a3RvghenirhywX4UaozMDwWuhu
+25pIWYo0am0Zk12rw0y458WZfil56BWrDVcxrVpqKMdZCUGfziKSm+DDph0oph9
p3Nbn536KvOKDqJzRcbzKKE+OoaSmsivKvqkLXdMy+kMfhpfAqGVz/yRxlAoTivz
cTWkuA2ZmqYwLWd6AxIKKHuxrsiR+xPq41DO2A18MaeHRV75SM6BryXkorS8k1w4
pVI4wvACccEaOFMlGHVKZ/Aq5ohaD+dMD63RZnLx31iyaNMkRlgnXZAmfhDukY5r
f21fJbljsBobIQIFYtn1ro3OqVwIgWD4LtrrfPUUnG4jSlIYqBEi1kvGZxaJ8R0p
ljPj1qjrC4NtgX6FMTALQHSUwYadrGqQvZp91NZqBZ4vfWxB99aV7OCi1i1TGe3w
0A3bE3zez1pfim5AERqxepmJb+3J3ay9NIYL/Kc1zOxYl2hYjk3+yxuG8ji4Eq6b
zXVbb9eGj/t3mKTU7WR1HqcGZM8Kkf8eCWnEx+TVM7NS0wbGPqGHK6rw/c98ZRA4
f5blWvyPSXod2xEaWhaehXiIWsXdtC79elk6kaoc7TRu8+cAWHE31ZBtsF1krSHz
FPAWENSpaT20TBWyBw1Z3fwi9pg9EBfKAWo5Dk9Md1nL296Te2sMC9OqtANF27lC
zKuKib0kDaXk3ojrCiX7IDz2VzJsVHaj2eg4NbLrYeidP+KXrvgo1oFnhi96S+SS
M2OAXu5ZD09xZAokGg/B6TxsWvcobCMSXkoWDygpq6tpCc8hfEYcyQaVHns8oaXI
ClSttP4HzcmHXPoPEuiWEUKA8eSWKwqMPjw3Ad/AacQCKUvCqCllS6lj0QRdKrXL
2/cnBWuCza1zwOmNfMf2t4I9P6GYzIhcTDzZltz3swUgJXcsUS6tCFK2lc2RZtB6
7RUNs2YSDhMj6nIJTV/LtVaWV+VXMz9MNhe4hRnAX639AAHOp29knXJ35/omGVFA
bA3VNEZ9pJHw+sPpRk7zZTsoHNDxQEQcfHVU9fkwMRvug1ILkSC4xa18+dNkUpQ2
75l7Q/AoK/1QGDdDpRsLsaxZak0FQxssGctCEo8xq3PtCauOwIwJd/v8vhDNKsHz
rMbjZqLNlpSaDzVy82E0EPFmhz6Ghn04XP385ruBeysiUgHHHHDCpW3iTU7kHROr
VYEtBNAA905uI+v31zCOqOkGjWZx9zKGz56empFqdVRfFbHQGjUv3/GIY0d+oskG
vB/UatzF/scT7HJBLItWHmc8SWzTsy0nfhF/VlNURPrIDIpovjosiJqgQ4ct8REP
bPAyGQgGtrGR69ZtOBSaT1tOxjrTJhioivv9idUyX/QstlixIcOcyUT2gO2OhH2X
8FeL8Npap+Eenz3jcIN8udmbBrBJFmM2gZc8jWoT8ag+H8sbhm8m/ZnAH+K1HEDr
AeE/8eDs1ykWFMQ4hAMsUlPJfxO1+hFM/tSlfI2HEv2jzTy+R7aCmhH0bE7HuMno
YpMYgDswFPfpptu13nxZG75rpHJ9OoV/TVAXPVhUBoTd+Z9SV1K8iIUf6+LXdIM0
vqClKm2tBndweewqhT49gfEJxRCQitnfJ5/OEzGFG2WsTJWH3WaCjKaeGCTaDhXC
SDmq8/7Gm7vPsXpWM8dzyBBa/D4VBYXOyuL38DJYIU0LnrPSDlhbV0IW8/ZGuoRT
EC9G6fil7+QyHpzmZnq9wBlKZ8jEoX1GXHr1O0g9GTJ0IV2ZRWZ3FgbjGhXpCj91
bEHJ5fNnexccpsEnJNRB9wnFOi0/hTO1BXZ2Qo+po4YZp0t0JrRvFPiprasvZ2EJ
UxbGCJ3LLU6bGq2mNi6au3kXMz2lD0jSnF7wf5SG3kf6Du/LejYwNn3HzBeu9tl4
YVv5kslnBaXiZbSfukM2gF1bkP1Y6UJSEHhYnRKsvn8VThkUAUm8AzlvR/bp96gO
3v/TQonqZtmlNNBMoDCcn3Jr+sl1gSdPNC3mZYPrzpSjgNCjNBX2948zcIo6zysy
L/0R5ugl87JuYRHeQyIXsnzJ5vDB769KzKvwak9x06EXGyrpzj0+zph+Czwx+Ovp
zyFhY7BKYmHgR1WGUyJTABfK3yRJe9msks7l/h3jCQPLb21a05fHPpLzryr9JRm8
zlwyJv2bIm6dMw8wSg7I8TQz580ZVabj2ypxs2XY4T1kCcwZy//XliBYksyCA4i2
6RfcXn9UGo+nN6MSshx/xFbNjBSbYJiRzV1uPZX//kaTnlv6KI9R3D5pXNijmYG9
s50gHl+ZMRlHrbnOJcXgRjQePuVrYf5aKWhAk76qX0VzjRmb8pg4trKVQQ4xp3tA
XIv4vgazgUngTFbD+e1JchxdPLR/kobxfh9v6Vi+P3fWu7D5SMhUmCY2nPPkffHt
qepCt2A5VhhExShcv07rs9tds8JMFjUk41ynjXfUNR6xqW8Tq8uqqVkKyJKjSwHC
InMEI5JIgcUwek+TOqMMZM5VdO9/a8X5hQERZ+Sg1CvuPnQ2Zzo8LkZ5qTm4afP8
NpVGce88anaDWvOaKT0LHmuLj/TchJ84tyriBK888Td+6MhWO8CD/bmMV4YPtP8r
5tRHQeIEDW1MQXsLhx5aCbzqcxzv7xQsRqC3pMwn2yyXSMGUVAI3WO/bvR3usV+V
Mdl6cBxk5Q1OHkdTO4vIhuHd04qEo+3+CtYlZuHZMl/azDfTWTC9PbVBb3HlDsiY
sQQFAzp8S/n1DWclRLrS2B5qnrAYvWTHg+rvKzyLoFDd5nAXnIRe91uSNLcS8vuY
gyF7XCJ2CLeUtNJvRuU+SEVKbdNhk8RY6xcRZlhPpTw2pNoOaDtN5NPfscDgg9RZ
XArrABywDID1RfmIC2H/SkyWddhhwTJ1U30Smai8vW6jhHPXBUWIFwgrwsLaMZkH
3xBgPKjYxDYvNLlyrZDmw7FV0rwR4AKIz0D9ngZlsxhjeBT4PKCfiJ1zDcBszVnP
NvrkzOOHoyJgJHg3zh+9wNI0apquCF4FkixK01K/eMQjBHcylzCtnirxURBzcaR5
BtTrHUvhZqfIMl9nEsMDZT8fVWHBsjpTGw5RuwiLEFEjVvhDEtbLQmWMdbxCuSoV
L/wJtJus+azCTSc8p3XUp5Z8e/ZRDAGc3Y9hQ2UtLozZLQ5Y5svltPJIkChDcrbK
Jic5KXxy/vKWZMXyQXW9IEM+vXyMnbh2VEbgjgUU/9xWL8EbZ1AT8rwRbX7dIaKz
11htgo2FMrDpDp5iFZ3aqHiG7TKb6enKiGeCE/uu6w5WYvbyxabj1j0sfthVlhDO
vCbRybYHdGIXKKe8+YvIjOq9BTDtayGkTXB1WZw5h+yejWXIF35MI0YaEIBMRYDE
bTj57fCOTwVXMHGt+OVSxX7XTMi8+xOg45MgUm9Tu2I4h9gT/jPgp8rJRtdUQnHE
WvPcjSkZG7uGkP8g6wgoYF6WbRlZNwFro56Hy+42ZiBNehXlsJOSZxteGt9iu499
P+U+nl17NKCtYno2rVf0QIKlcXqK2c+AQUokjzF3fyz7+AfPvI1ancjovVWQnOGx
ebK7GSsfpvYxnvQTSqRcRwyBwbij6nkUQniZHws0YgKPnPRg7Zmjnf/lPH3EgdgZ
uvIpPC12+1yAtyPb6VMYW2rbA4JdOFStC58w46QQ5Gcc0+fZLeHxat5wxFYJQSCd
C1PfLxuUrUiR7pKQos3bv+5auNfSztZMeUkNgi/EqOcm5c//1EcuwOVprlXMDy6P
Dq04wjbPwHX0n/DS8IXIX1PBV0+Tneh1wiKdYP1O3mCKxP3gIj1RZkqauFdj1edg
reTmAoHjBmY24j4qmaJ+gSdt0d36jmWReEbqRIlkmDRPIr0lXoF6k4qxkkimfxLm
JwOS0bUNK1ZmX3bgotJnrV4l64UWtxyxmH+R2m+RkrGDHV5rwn+ZjP1MfYpsrEqt
QYnfN6C0F2ocN82+G2c6+YlGJoxfnO0e/KhPHRUCvxnFpoIZZXiioHrFwCbh1qcv
EnWhhtTH5/v5grzqGbgC3oHMnC/jxGwbbp7/ToUIJp2WinZCXoVDsCl80OibLIXh
rEUaZiEmTTe/zOtpKOMaIKFOa7X/CrLYLmWgD47Vsjld6e7WqATvGAaVQ2igjFCO
v4GLlF7rzMG8BAjRHbnIMSSbZBPy2w5iRn8/sAhEs0SG7xXmZ/cbI1Ka9cL0Ikqm
qcLMimi2+ibYTnmtvGSXs971mTf4BYlolu6yyG6y0VHk7JgtvUwGyiGZWfXN2z9h
kJOcXqmJqrEfeiutMfiNNHiwOaMUKZH89K/bD0WuEtzhDZh2h2vd7r+bj5B6cyY0
fm26yk4QxkmZmjkvXVGQPU7pnycPEkYpT+8/HuiVzhN+wglzg7ajhtScwlWbUB96
dPOJmO8WWin7Fg4pX+kz9P3gMlFXLmAFGkszQQ0RSJpOPTpKvYUJwZkBvreoGoY0
ulLiEcp9FeQtURDoFd7H89GW8NHuocNu1I1lH3/tc7n9MgoQ6Z5bSYLfbQewq2Nn
7SFyZVYoowrF46A7bkv2AbjLE9WgofUrzgEdKtsRNX1+Yy3cTgMhNJ5Z5Ve0+6sO
IN1Budn7ItbrnQtLnWk2SDqmmwWm3CT2nlJP1mhDgBoiATC2KxHmJ3ugyB/f1A+v
Bgo4voklzZ9XpK6PM+IJOnd3Obdx+gW6ThnacBTzhCBNRf4R+6J+8v6rmhszOfrF
THxekTHlFiwaDcEzveMEjbrVJP22piU+2X5P56vHmurZN8PiCbEPxV10+3U2ObY1
8J891GMUx6aqA6XBHKpoOylL6AYoMBgV2PO6lFXWdsyGaMiykER4oPnJewusF75l
gs3mYsonA47AsCyR/azVTuB2EyN/6QqNp1EcIwxy5CP5abILLWmgAOrIc2lYFfoR
YyzslOzyvCrZBa+xvfr5LbQCK/8GEJL+fJmZ07//CfhrGQ6af2JHVh9/9yk067yQ
oBgmTmxEZxHXpe4i/UqR7fe910Ku6WhrS3lTyye/7BjO0LrOkZRwqTP9mHmfUpJL
BLPAr77DlP1ghXV07xGh/IFQHDmUu2c0Aq71wrjZWMcxYBm0h1+KhYkWIjjFFD0t
M8V+2mHNgTyytU15xvGX/nfyV20pDAtevFppFSCsx04vqrymsgSmuHGTyLSIYCn4
iblsAaZIQpTuVucNxTDG/20rLLeMCPqMYvn+UD96dxurOow9IjPIy6eZc2sWCDAr
OXwwzWnoq5tu1TBlSLuNdvKXoEH6CBwlepjTO2ufvYKg9zfp48hPzML32NjjJ4B3
6XNDl3lIB/RLyZ4fNXLSYTKLI3qTyqO/qr/giUzLEzsaqGsoVf23kUVS5PxcwJ61
LA9jH3gwTCr/U2SG8j4R5e7048860/KLFViRFKwchYVodkYq8qAWg+huAcvD6gaP
EiIHRA1n1wrIR2Otbx04mSg+2NZ9vdrPcS/40yjHwkRV0oz7VtQb3VYK4+K7H05g
v8mwHkJRruZ+Siq3ODZznrA02H+kTfq1FImboPjpPI0NlmuDgXbw/SAhPCo1LSFD
IV9H8JVD7wexlb9w3QKZelwNCimUQ0CyRYpEbJONLYAn/HuTDYVFR83NDwAmmXlH
KGN0XFyUywhQZX/IMgbqxSt+IrkykyLYoUMiu9UsorbnduTQKt9L0I2c1g0Pkqzt
JV9wY/4LX82i4s60DDFzRi7OJU1lpb1yLmLtnOG9K6+cO3P/ijdYuXqo9BqOn3DE
URdeEXB3eub6YWi9OSXvzwDG0qwfR69T0KJZ3TMfdNg5N8V1oTFr7+7PLgvE+t29
/N53DwNOAz+tjAgd7cBMtJyYY/vb21fwMoYE6JKvaQL6lxXjZPbrO0sFBbHtpLAl
EahC3NAIDVmcAJTVNsbvKuxL8/mw9+VZQqSKH/Re0XNWTBuu8rDg9HeidyqPXna7
8l06r0W0hhW8o5PezPIwb3GhYfA+yVHQeGFH1nhAj6K8Mjj+RRF4Jd6IRfg8VnbN
b5m+7WC00E02y9pVfFcFpNXFXb2dtgQB/MeJlfSsdYIQ19Uu3GxjFzHzkeYA36KE
H85lCPfKTk73hlkvaX148TuybEILuLLxYppka3oxBmk1sUbsPQjxp4BcKVp1ARPE
he+Zp3l2ZnvaYyN1gMVdWPEJAr3xRvD60r/N11saB3X9hAtCUgG36oe1djxFy1Gz
szE6NcJZsB9/skChKi+OF+jfe3jcMndULExZcZchErkoOKzMdZbczGsmS/FVamh8
xVrC1UU3jUKn0z49Su/1eFdJs6TrbqbWuK3A5yPi2NcJRt9McQl8Pv/I2Q80581y
EK2z+ueSwOQn6he8O40g60+wEptIV2hHp1QIkAckMEXOoZGWRuKLQCkZZCbGrSuN
Bn7LEFMa5uETgAZkmvu8MjpmAbCikqmCqMrx7hhxkrPcfsivxBUr0PUGq/4fErlJ
nG8eVSdb4kLdw3nvqRaUmL+mbgvenbJ+vjb+Pwlt6Ai6EwNbAnQ2IUxYPT/wrR8e
xw5G/WMRV7grDVRrMrfs+xX1RR71W/gHpdhn2UVaVaZlGe4rqWu/JHVxNxkpcyg1
5vVT/ZRVP3JdKM9BktwOwgrPhtmg3OgFVQDw1vxbQyVk60xO7spMqxoxNuhV/NJB
7EC0f/kAxzFT68rmLjEMUCP20qz+Knjtqrpbm3Yn/OMkRG1QHUMR3XeOQKl8fwzR
JXiR5xYVPIQlaDJmcN1sN+pDX+gK6HgYY86tmqbc5pdfj6+j0w5nzVzDiHNe5ML9
ZDQXsgDQx6K4TZ2Lh0ErWvNQyeAZYGThBn0BtS9qv9MWrmp0ag+UDsZBwuuocUiA
QABFHG7U+j8vWX5Vz/zJi6+yrEbJekRFrX2Wt3h7Ics49zx5mZd3lqTzBggS14mS
8bnjxprgLSciQ1M7cwC6rfUDO2aLUdIxW7OKv/eWGeh5+QuHzOzjcf+yeBBJypl/
i/f9dCBckY+/CcsvnL8wg7gtSMRnX8gvZCteTMcKnTPJsaEb4mdfOPqM38VcIAE5
bdy9eedYcnhLcbH+es0OOQBVTH0PPTDi7/GmIIZG+rZhMSK/wcZ6XVHXXSnz+R0q
CHTtGHwvYg99lALN4igmMP7lLZT+adgUiSzLJaMqxzPwtN4J6ZyT/wpO77z1IPL1
mCk+cYNVicylI0kQOzooGIELKY48l5G0Fb8laSOExf8tesOZfLohzw6IhzC0wzeq
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
AlkHi0WxFp0KDehe7ofN1u8vvf/+tkCCObhBgX4rlbAWI2YKGMZr9L1MIe9zRSEh
U0eht9pEqSOlgVekd56EMitXi9L2PA03WqTB3JE/hQHgIfWo5144kI82SlcflZZH
0srahMja7jc5CnXNEdf9VClDXJUi6kJBH3cqP0e8lTpuucOgWWZ3zazRmtONmYNi
CNhjd7WOQMH5/tn4zScF7w0LquH4iOfnR9qbRUPze3oF5EUzWoysi8GKWvy1D6k0
/phk2Yh+Hy0H9jR49KmyqFzVByyPNbFqA4vv9q+lS3UhpUT5FUmCQVrQZ2w4QJIH
/iaOMu2LGr7MWl53LLcepA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5392 )
`pragma protect data_block
/cw1MoPbLytNslL2TkMaHjKU/xg5AYpBvMKZCvrKt8fKzys1TmSUdBoycvKFKtqv
d9/27q8i1p9EF9dzYJpDL+PMHHIlb1N/drHMGv0gimcf5Q01+ZvNgpViXBr4I8Vc
O6aG5j9rqp04bZ+d1iItCbGPZFP3Mdlc+nxEkZY0kw5P4/HrhwcDzKkskCHfKEAI
3E69MdTutxRMQQDdAExzUpuhLNuVOWdYZ9cV79sUIYkW7s1cb+jTVvTsYrLJo/zK
iHo1w6Er6u68Pk4Uo5u0KtzTDn5tFVskDJwhMRS9U4p5ORAx2hFzWVtJhLoxa+9G
+Fo7r5VxyPc1HL2jKKHyI9wz0+myKgVnsvWj98AvY38ly3rSFuPITtz+JA/jzlsY
dbx1PbiWyMDDmqMrZktWFKQ4k1ADafV/N3FanfOkYD5G8o3fO9Ri4U1PLvwkg/W+
syb17xths/g1iFSl1z13fwpkErjNu1xch7DVyWEqqMQfnJjVIRboXWPTOXLxuqjd
qVvnhvB5aRd+n3+IVcwov839femoiAFxI1vbjhngg4QWjs3GSAkWHM7YK138quyF
vZZUAYCnxZCX0loqa1ovYbr2rmQAkW+pp6bsbch3GMWsXPLlVqvgFezKzva5j/zC
2uLz/cEH3x0zu0W5vqvxH0/AGuFr7k94+J0dkMUtMSwaHOHEP4IBj/qLmSQSJfbh
7G3F471Gh+ia9OETBNz/DoCmLAjEHOuaO72bVfwvIR/4HIabtXKjyFJCe+yyVQKv
SMP03Pnb85ZXwZ480Yqx9NRHB0h73EGeU/+6EYUJz2O3WJJ6xH9ODbiCcPHiJhXi
UGlC4RSSd00Cdcom7bMm1RRne4OaYD7UzMAJnOfbrDR/JHp5CXRUmiI3P+bVuBas
hROdTlC7RgnQjrzuWZmuefCmp2gnR3lrxH7yUzHvU1J4QzlVVt+SEBCMVkMJXox1
2Q16k/2MNifVaICR2AybKEyG93K4iqHG4nyzNkFHhqLyzy0rOYhAjF3nhtpdmOwA
bsnZi5HwVkF6pcK/iNjYTBPMB/ZNW5i9hY2jRZpKDBSHSykhGxifDfPbVzEcwHB0
5EwPdYnc8V1jg9BsHq56Ahcv86Ty7nNTHOPKOGYRNKPZG6RgzxvuOGhYZvsDiHpD
FKh/XrRC4ELmb+enk6GEXwKxnoVQHL8vyqAVEncGYp3vH8iKp3383JU96lgcFwpy
yrC8+BQ//e4Fl9aYB6s6AeaFXRBIAN8B5GT55pRgIvG7MI2mtJ4/NvoNnnIL71G4
CGlqZuWUFwO0Fl5q96kl6LeaNb5mWirssYRpfhxe1LhhHe3zmdJNiG5vth7h1zsC
qua9R2VJ7HX1OCX8YwJ31MSbOFWLODOTLUodY0puYA78szfHAHy990xOHt3Y9PML
qb2BFTiRrN37HTjA+vKkL4jawEN7F8jYOL1l3H4HXrIt9pac3BufDOm600bJeIor
Ihu+VoUIIVm94C4duvi2Idp7KPGqFc+64AhMEujbstQCFpdocQ4kvRJAKk0lfKoX
CbPttO9+/OxKvJZ41bCBc6PolQfCF8+5PIBqTkyyEfuB8w9sP+Tk/HGzZ8Zc3Arw
potf3FucAl6dX46G1B6XPmDvy2dcik0z6C54yTdXjanvEfB+h7ob+2pE6g3GImP9
6/d/otT0ruKD/bkNdMni27MFLb2bA+Z4o+ugv8IsjCTYmikPHz/wK6mhDct5Ww/A
eFszkjxZIQ8QXxJFVRDIZy48lY5q0SIASdQItwTc3Cil+dcW3nMvd57GwkHZUiZQ
O/zv5seid1nsowhuHoK6R89W+7etQgP5UPwDNEqG0rV+dcggK618sJXMI3sgYLLo
Sq+DrWQUXeNPXgsj05I/POhXBKv+XtPB6TiCwJ57/S+PiShejwGDhuSEYv56hhvJ
UdML5h3JFCV8shbO2IBFdCWZ6opm7gZiF1SFeXAW3/BprmEEB2grWGE1KBng7tlM
9Z1pXoBtUJGAR9u0hyKeZNcDihwicHBn4tHVF9jUEvGEnc3TU3Fm5mwwKdCdST2V
cknqPi/ACIUQW7CS9rTIoOycoxl4Ox7jqbntaQ3hOzCUTcrA03mlhFSmT8nPjxO+
uG76BBtsN+09rw4D9f5w8Qat2rUqpde2zd1k66teuwi10lkImmywJBmOjY26HTQ7
t+SOhSeX41D7HvreRKb++nesVf+Sec0l0MDB8CYN8ETB9Ti52RVyKpMMto/wIUe/
CkDNz4l/Y72TwYNvJkH4R5KOeho20cu7/tBHrRmumMaq9X8wckkYwAQKS3s8XnNr
qG5TBpmUeRXssWmrT/SUueZ/q27JqkTfoSkLkb0gBZlsi9Oq3iE7hEP2e6bGxyZ+
/gcBJKqtB6/KYwLBK6DCB1OiMjsprrID7hYpQWmS1oeyVjWuKSahy1v84GJGhyOm
Ne16Z5LNWmmMvfBLCgaHIwhdDtucOr9qmtdD0Ef49nAOgFLWwjIQPDfKVSIxMC5r
4mptRDIebi3YjD96Sr7GJ59pP/LTEvBi59VNtkOp1VLg8Fw3FIZ1UgWN21TBq0uX
nmmeJLj1cjGEOJuLslyjOHHkX00/bTlr3kZ31s165GsiCIAk+UDh2md2scHsgcdy
YgUu9LgART3SiHWWH4Px+eRLBIOBcr9qWq2C2wT05vuRxgWdVBe0eYRxhb2nNv3M
sRvhDDFIbc3ZU0qPl7pRYJDYSKVcbL8j0YL8PvYuhYYoaknNvEjbauhRnAGT0MSE
hv7BTAv/qQYWiAJX3YApfCNyQt2Ict9n2QcjtWpXaNmXWUHiHKkePFsVpl9SWpBt
AVC4Xdy7BEnvTZDZ1U3Hyq3Y58LTBydaCpCdJVOC2bmcr8h39Bi9kZERRnBnXxTB
0UeP3h+IDZoRcPOvQZWMknwnFNRK27FfQdv5fe5bQf/sZ7BA9CW61tnwbNNpmmUF
NlTjJy59Bu2n0/4gx4t/PC0suKjCPxyQXfnwhslerQz06japvZg5pVX4LuvTOfzO
bInabmkX9i1M+0yugIGu6do5ZDmx5u8YfRW33LPlAKcOTIQSail3gu7TfNqtgT3G
pV8YnTqcF7IJ8HyHjxYaN/wrPQNk61X130scKqCN3l+n9cPouOLYA6V3ojqRohUG
I4HWqzDccvVIPrwScU0/Qb1N+KYzcfSZxSScBxUXRkGCSvllkv51fkx6J3NMWMZH
3+JorNshYxjn/N+k5X8H58A1ZNdx3LBgLC3iQyAn1Gq8jwp6lWqzRcBNBEur0OUe
p7nCqiFDEEf9AdTwft1cTzRd+GqnRDSYqyShrzKx4k+BMK6fDfZg3gGz8xeRg4tY
bkfuaX78tfIwBxPDkLHfypYU4DL13gkCrfkk1F0I06/h6l6y24AL58B0awVBFhTv
Upb/tofcHQ1c1ugp8rokdYWcO0ebw1IpGgSgjMFHOwRjCbqpcK0qNdlts+LfqCB5
JYsDBwQODwd9R0AYzNwdlyPbOqyfk43kU8umpcpyv5n9Bn6CCMxEBejDswFzvr/x
XeGxn4hC+JWbkJIPSsm7U2/ZMYejbpspdA/tNKV+ncoENkQm6b3N5A2SvkHGMyI1
ZGPplymmkLIshmabpZs2rw1s1HAzxAn5tLBJLi9rWJb5oGk8l9lJS9/V9qDSL56g
XzppSM75S701iFAL3w5AQnop0ICt/ToHBhxJVx0DyfVE3votqrW6nc5EICWNMKkV
8/+Ms1Gc3sL4SFdAOx9QonFcv1A4pi2y5m8+hbg1/rgnha54ZirxTgFctkWJWi4x
MX76xXrZIYm5H4q2O40m5/4W5pHp++TXRp28xPRyvDfUrS/P4lAnUNi44LtXoD7B
H2BrFwmcQ0qdPZrbM9UlM/daynOBtrVyTl5STSlAsoGdKhOrTn39lO7Px5fzVWFL
QuFP4TnBouKOha7lDbbgez5Hs/EkH2NAdhsES7+BeiQW8GL5yVs95cvj5Ke98mBC
sw6DMHV/ITurxJiIo3uV83AlgWn7go3piqmIIALVXtEiUBdXnoU7Q5OWg+DGPTDV
+a1lD8t7dze5WCA6JpIoipqQ8dcJL+cYEcVuKpvGOPDhEK9nShBiEJ86rGogAhuE
4u+Um/Sdkdrv5fWQRPop3mrYNcW1H2dQN5xGwEdv64WzcoDcWHIpSBa/tAXTzJw3
efndS3DFxuoJXH1yFYl+o1Nksbye8Y+Axk00Dbsp5JABm0cUrwVvWB5VeRKwQvqD
Qug6LSDHoUhjBqq5iN4CgfwgXr6fThsPvrmGAhw0thmOfDPIDi0ZYiJrre0s/u1N
fD1aCujnyiCrGKRD5gE6wNMYjEwDeB8WpQLNIrEa73qSnR2bBr+mHalO9mtBJedq
7IjaPT+3S8+Cjt6UlYILaFWevRRNBucH8aGSvWr7HLK9RGUcjhbO7DCuaEANmEr3
adYq7h4XplKfK5aMzYkoTSCTgqMerzoQVnnFIGeNg1NiV+RNI1O08vk4O1O+MN5H
EijNmMUWqfaHdiy1l6bXs/mClCdoR/LjkmuqsLsC2wRM9S21QIRcfUd6jcE1Yne5
XTonEJQRouBj9NUpuWEelM4lXdzDFGG8U7rlriu2c0zPteTjX8NZJZXT/XaltkMW
LD/bS0P2Z5qYHfkFgDpvkfMvy0rVYizbhiEN/ywjTlLQC1mEVGWAjCo6CInxfLM4
RPLU/iVIgKZc+CTwcsAZl7Lmx2Hxyjy+JS1ZMYSl3wJumgz5ZAkiEdrQFnQVrF8F
kLZDvMJAUWUcTLWVx3hdlxfqsJm21t6CZ/Np5HkC5HT6YSbe93oEm8Xj88YDZEMG
jAWiKo1kC7S/dfKHWycHO3C71YNv2M0hE55eifvRabTR0K2VGDlYCPtgFJ6dzdvO
cu7vTJd4mVkgI3dQIzD2sfz5Acn+2gHsGYbPDLJ4CQmKiEwy4JsPZXMGQY4s0w7E
j4DA/bBYLwsLbcSnlqblnl+W8Arlbs64XlszlnwA84uC/CzA6rF5ZVwggadE99Kt
cDZ+juGOYqZuzhY43nhjiTZewTG+swEFJnkvdxWudasjxyQwH9vsoHB1JTEe1JAR
0GmdDK5Kepe6UX/4NqX9GW59YgzBVNxX5GMZdGnsMwBT8kGLgfqwAmiqp9qzeVOc
bD3qo+BwwRqdsEjBTLAmlXETTLKqtRWDdomomsgXTxwMi3v3iBh/nYLFOkO1aAzY
/sGqFLnhVT3ZD8rDPfxgIyR/qvN5hh5AxsuOam7XIb606pyg9v8b4O/cy5hByp4E
+wS+/PobBWRRcbX9F9I7dCwjclF36yES6ANZYSOqttVVJps2R1Puvvzzbfg9FVtS
gtvFYgRPYJOl0FlLi59/BL+pkiHjn4NEzQTSOKoXGVjIhLEz68Ti8JOxKaKYMxLC
6uZcnikC/NVzLhHb2CG8vQJTcj3lYiakeNUC0jQxzk7mJVftt5p9DtnJvsp6i24U
3PqM25ynfQwca/Ruxvi1jMT8E/qiEX0Erk/0Dh7ZIyBMUxsKsia4v1ch2GULO1oI
MulDiM/MAORPCssZ4pvzM6NFhTcDjKe1rXABd564N9Mro10s70/iiotWr5S806V3
qDsI8VQztSAHfXmn12+ffyKF3uZ3VWbilRo9v1FMy5NCcoC7GXR9qqiXxpbrcXFB
jK8pvrE2cWvfVtdPnwfeMxcj1eWQxz2vYqGo1eXrXgGwV5ZSuO2OIBkJcxE3GqgZ
v/MN6p5r9hy+lA52o3kwVWR8IkVPAFEG8wGexj91MM447Hg51s/S6bXPYI2VqhTM
3QfqIqMKHV1suOZmdG60XKJME1K9igsAjKIjJ3KGm7wIvhy3izEUrwO1wKLt01JE
dYYh4acaZ9J5hNba1unJ73plT9FdxkAsMZc0i6INGJeeWJ7/AiT5rXT7FaxN24OX
a8cA99gseTDEltPOvJIDPU2LN2OkBXm9uUUDMnp+0I0vGgCAbk+deLY6ZwRQ8lz3
jR1imkQIfYcE55g6x4ytoI/HXk5OQbb8I7NtmRnp17mJmbzv0QedJ9EJAFyV5SlF
Ddp6+pv9ZjqLL5csZLmFTiObCagsgdri3qyGH8BmmdSgsGHHpYSa0VOuqfDOKC8a
16y5aqAzZGA+PMunr6X/BXJ19QKN8JrR7kDgRCqqggW0nBWrnHuF88HdKua/B5e6
mBAjwH0Fb2++pbFHC13DGBm/s+8XFCbJa3kD83S5R2B0Y6YY1eHNKiR9EZlH4x0l
8y0qTwfxS5C4trdejggsDlJVBXOjlrpdABmsV1zk9pY7J7Ge6SnqN4wxv3viOdLM
kaWyiHAf5oEBmosb91hXVGP9LFcbubGyAZAns9CEJAxexTPj0O2fK3zzt3sG890U
fPL3/nzYxuJVEiFskZwDUgQyvYbQRT3t3eYmTY6YOGFCTUCXsj/HDn8Dv7s3Jcg1
9hrZg+6t2hwz9kInwIRDhAt4/V7JKKq62enaZdKHbXqN/QFM/2NSfp7prZ2C1WXQ
f60jyl64kAe7/B0UQvrxnalH6RCwsaD3AgejWfFgCEv70gqqtyQ+8zFWvx9BUhTK
TcQosGljyfarDh99K4n/yj45C2M271+ojgwN0kOnx736gGZ1ESy0xBjr/e40fgCW
tWUroslHvgblYE+8gAoggyABHCWGPjHXES+VTyCT2wcqDUS9nqDDqodNFl8zZSI9
Mb0M8q5eieCvOqsVEXwBYC4ZVfY4rYT+VZz5WDoOlbW3QtzvLdFI0yhx+/bgRfBL
0O3Jh/HgDE03M0Rb0YFmSzGd4APWQbyRqRn4qhJEW7cefZMCiM+9+819DvMGrzoM
wRk2pt0sCzQWAAT8IoZGV2X/plIbfhmddNx4esdZfwyLCcaPA+yP6rdZYhgBdhVN
Yeu7N+Yx1UaUT2VmPieWhEqq9P7sclJoahlAdEVoBnBVWcU/7wc4fPcohAiXYUxg
xpAlWnNcUNaZv4V3aDVBnOTnssSE94eRYQex7TWd+iAYV7LticMk1kgaRcce+Qtg
BdiXlSNGpvw5SvYp7HXr++REvDKzqDSSi0uCjdbkVlmO8O0BqYAi5Gbk2+bH42H8
AmueuF6GWvvdg0jhpbei155wKwh1J6asmQM11i3X0ks/95f/63KEvuY75c1qyz2s
SPknlSqqCeEBTvhsULj5rtw91Pt05A7l8NKirix7+95wXzo5+B8JSI0G6aUjPuK9
eD5UvdtSs0ClHCyv8M+pcw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
U7PYkLBFroPgRS7g3jEdiHbVrifx0riVWhJ0GYR+nrvW9/X1MW4iyOa8fRfUizyz
3lnEDw4LzLJPW/3a2qj52R2FZplmCUAh4kyliNFLLYRlamTzXM9OU9B7pDyBNzy7
njWNwUpcmXAVLLDmdSI0BiAEwNjCRRlKQrT2C79Q2zqK2dyEExEqywcbaKgOaadF
9/KFS01cOwoLQdEpk1XsOl/CmiVJdguw0LYCAHjrfW28GVb5cf7zkzQGPtieY3/I
CWkArGCli+9cHTs8nBkHt2pD6JEs+1JN/L+YxzXcA13L1MwNO1YMQ1uy8ooq3M6t
P8LMNeQJZ9wX3xsCDbjVvw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8864 )
`pragma protect data_block
W2juK0b0X6YIB6KIM5X2RRw6siQD6GNFd/+3orbLi8oOVTzSAZa0R3s6RHXFvCu/
m5s+NazDExTuW0RdAhMp305hxYQ9oXRz37XcdxfxBwNz1hO68k1GCyWvOGGWNODM
rvJwO+znB/qy2kbCV4UgjkcN7Nxv3zd0mSG8ATf1GpvGTW9jGehGDgCoZ/kCzUs+
XY38NR5p16iUT4PhrY56X6na49IAPzNAFS5TCbg4CI3TlCShngS8neWCyhYv9Hzy
JbBSb2mTo/J6dSYZrFE1Afo1/cMn2IgS8DBxxMEfp/Cc3ROMUCY2pdiFrv6sGl3f
U3IqzFwjdLTtvXeMsVJnNdg9L057vjw+3dHpXJSmw8CfSmDaeFUj0awfVnGAjExO
rBD/ND6kddbwKH8AsRhyxwTur3I5DeZ7vUd7nUzzX5Tv7MbiVcRblzrYsTK14FGK
Ml345+xwhp/IMCtJHArDuXlc48MeAcBnVrIxj2i9eoc0JezqsquJUNrtTB4eBvLy
ppDmgj42aGT89MmGUKqPNyZHcPxy891JmIkFxZZZ1AsMDzpXTsYx2yZq4hA2+oNQ
XewlsQn+MRF7yByDeEGdzgWIfpnUvHdi1YO2GYAQPBPy0sNWHi7GSdDK0YjWwhkp
222ag1CHKSBg/WaGBQ0eP/1QSsGplwlsttLTUNcILMKY8kMoxjHrEsu5CSNhUoZ/
TtTPjBGoe98S1w1UanXlqga/hv0Q7dFldXqbdeActWfGsG1x09yoNdJ4y49kwhCi
s88Dm57h0/3/jJpJAOo99GpF2v45YBCVFs6/YIb0IZCwa51f7ok127aLQ181eEvU
lUPq1ZPF2hMjCWzktbsvWUwONuOsmQjHBRIXPXdcj03i/6UtKfblBA+QdvEZBg0r
8Noh/RUxIDPDN0uF+8JnNN/Zi/Ss327aYRR6LpJFs7GtXnhcnnEgauYD9JuoqBvn
oN7flHX5RPMyJUSuIllBu/kBySTmVGMa5XMjICuOoh8hdg3kkaJgZYymlo8KNgy3
Mah12g9sTWiJh4HvYrtUgOZ5bEj+d+nx51GZ7pNep5vtKRdZcsKhBsaO5+EnruNv
GvPW02DpVblt30wMoTgPf6bd/I/Z53KlYOHROQfz3FqXLOWiFTuvfJFbwyuvoYJR
6m6LHE45pCtcXULka2zzzD8ioxPP5ONAgNbiWDwDpF7Kubkz5ZEej8IELxSgFNsW
qhkL9GCAlsowHCW5c2i8k8zLl43vVEe8MmLTly+QnLkELxAY+9Nur/Yt9TihXm2X
S9fTmWZt2vSUY5UZ6o7300Z4HrOFDqujYn7GolnAHIYld+bfqVAT2MNN5apGSoGg
cJevhCVD+Plmakk1z3dER/2Cl2xaStm8gMnFNuAwf6kJ0+qfJd+DwsKhpczkwXsF
kfAEtWHX6cYD5yu+C4VBaPiSQVlZwahFhOS8JkpOGS2h8LSIymgoQPX0xK5IyKuA
lqrpRnu8ydJIz5MVDaeQh33FrKnse0vJf46LFHI6CrKZDKUiPB/IUy43f5URXPbr
/rb1XM8IM/n5v4HtQB+7o0PoWqwsFoFncQD81V+96/6Lh5fFxrq0bJi6x2c4YF5f
vSpLlRFYIwlcQeJMIjX4l5X806MdTdEIm8MONjJOd+mMcMwPW8+kGV/wSB4HEy8T
rtyZ0lI7riU4Nc22xaoRB8Pszmz35U+9WNN0SfT+poRj7p767fYk9Zqd4lIxIxq3
vUJE4DuDp2bXpiY9EXnmzSvWNn50go9XA9Ou4hp6iEkMAxWdQzmkNQ+0OlZoPL0r
KRMYwgTomr0uIFESLiGuEQAYn0IvFeojCGyhNR5KVMlN36rbCYHCGqFQRyZZ8/n0
X1AV+PvfotKdts5LkR5T6x2K22+mN97Ot1b9ssgSM40EdCjHxe25gVsnIoxBpQoO
tmxjzG2TZOsRVl4sTw9FgvBkozpw8d64g91MmJNWp8q7BuvaxayFX4vQUDch5h6m
um3IU18r1FcE/zQVFzIH7esn5q+n/WH85faFukoYRAOu7oq5Ftwv/ypljSQ1U33B
L4OeOoyv6Uq/3TVR4zZQRu17e2Jy4HaGHFiSV+lr+7hBOFUeH4vDvTe7GYg0fuCr
8Mugpu44cJOOXEX8Ks/ltlVP3YI95eCd98DX5PNV1YQPJWvsRPLARPuYl4moe/Ax
ZC2jbZU+6+o44S5gTZPmUiKlGvj/68DHzcqkaMN3sVQU/JRH+nUjxoDoyI1KPCM3
hSVEQWRAdIJFzzQvhYDGkoAaRj2SkGy1m+DKs+yHpf8F1s1aYxDNAx/kTM3s4uJV
sLunhZZ0Sm2ISLDysspi2IGSP0TAvkuCaH/DRzvzD0JYiNnwRnAOtJBY3zdx5UyE
fs4AEhn4xA2A2g3zUMImEMb9gm5o2lE/cXK2/Otkx33DSK8mfKbFlgF5I28CyhTB
nVHD3gKfzF2YPEJiN8bxKhhSJGPDx4tLL6UviV+97v9zyZMw5m28GHu/04mWPk8D
gLpL4FHdsCjNge2+Mtrgydfgx/0i1KxPkpbOj+mCPS894bmoUyjs/pi1NDLyceYe
OoBpecLnQTvCEPEguX8f1G+jl3uTJc2CzU1EFGZs1xS6PtkXPSG9OSlp+gzLawrk
PcEyd0QXBSVYikPtXTVyB70rO99QWP5H8ne6ccW74Y1Jo1E0wrFf9oBpka8pjQQv
emrYwH+aQsstjZ98tLvk7xAmAH35WPbRk04161xtiqVdmTxXCrICUH++KoDhGOym
PtcqGrYO+WRf/9ZZkwz9TSBIllAiIxr8YCo2wq49oazvlg1yjActsekMRYMu11zo
gqMHcpV52d8oOk236B33zj8yps7IrD2qsWS6leB9Hs/NuflFwkH3ZkeLPhJDA03m
+Koth1ZvrIXQ0MtQwOFHY1QgbTMkTxMx9CQwkDObt5PNUC4pvKfEQvAHMtUossJD
YiogLryC18Umn3soL2wzKP5IHEZnoETx/IqBpOFtz3kHq7vLK05UbskItaojZJls
fYQ9htaOD4WQcZtPhJG2s/ODzTzVoHvvSqVQs0Lyz0rwYBzOi3KB4xlqLmdlzkSV
m+oOaQvnc8HVgid6cBbarFiQpoAzHJ5Z6K3XhAd/LMRqLtCN1LdpDaTw8B60DMD8
f/Uz9OhBPKdQgr8SKbKBc7WWxaw7k5nxJN1WQ25xv8M4+sGZMz4PzgzE1AM/rMpo
i7hsqLNPKwEouFTX8lRZ/ct7ODkfHv23uGRDII4gSMY2RddHS9oCaf4jtIl9DQrb
ssseGw1DFfiqHnD8dcAMbQz5LvwZuotGcsh4cLqKKLP8G6cFs+RoLOtd4CjHFCLv
LSe4F7xFssfJX9/d5sHscire+HxB5UxzK18CDowj6fS5EsRFXR9N83nrx25yvoWd
lZvkRzi0Dp1qo8NYlg4YBvra0+G3ssQoeQlvf1V/CDq/VHslsVo1cMvzgVU8T0DJ
FqmBDbBTA8d47Gqkr5ap1J/AqUtuP2wu/ZjNrIFLQFg51Emx8deltemHpvrJ0ZrJ
AKVTeIBCItwiyeZwN5bVxsFsz2Yo7pICC1XpyyiFDBm5NCMrswm6DuSfMSZXWdBH
UImHVuRUy9/seK9FCnOM4em8nTfUtVlpkaZa0tRG72EoQZDtPDtTrWYbMqIR8cgX
nDzcVu2DZJaEfccrI5oDFDQV+JN1AdvPmnPknRYLvqcdOx3w2h9O0RGP+lEb3x5N
bk+WvazlT65llUUrQ42vsXpsn1tKu8j/e+ytjLhWHo4spcm9cvlZpIRnHMTnaV9n
ZJXrKKSXP5lccn/QbQBO8I6cil84vptwTyEwxpbJfjfF/iUZCrYQXC4LE1R0k8Ls
KczKZK58KWwShn4REioIosFm423tC9y9Pl4Zi7PLB/Uz1UAlkoinXm/IITx4csFd
0iwrhpoQIK+Yzpcwv0Etxrx2IrfCNGAEfJkIO5S40YJbEa3obyw2OJgMMcomldp+
YQdEN2mo0SnBl5KFqyf3YNk4Wc+Mx9ehnY5yBGOkamLmw5EnVJCSzr7sJYP4hfJt
kD5Oz+oIFHe/SOhTEPfxma4q1nPdemLHNjvHWVi+MUjMy3Er+L59V1yal/pctBBv
bHvVjGK1CGlkhE2yLzVRtzy06yxzOjihs1qpnzR/48uik81HWEL2stPE+MmzKWiv
1P3KrYKG4xrd+FwRLp1x86dYYe9eICNCFwxcyMlHbAMtEWOV/+j2GIx3GRjjFH4f
XLI2uyDWmmH+jSF1DEENwB+r8gdZyEZCwCcShxMTZpASITMnkgjjcAew7Jang/SN
PyssAgm+j12ESe2V0UtdeEEWpFP/vEPGHPFbgvuEct8izbcZi9qGQcEyqJvG/O3B
51EZhunVuOg1vcvnF9QT47MrWzDgg3ZkXvBuvC/69r8sVP1YVDKlhD4POzKFfFQ7
H18FyADzPUEiz7zCKwDCOkKnNVyrRpmpzB4AxdA/M30rQln007UQWIVqFDz14yYk
4ljQEFulR/M29EPicaPbaKGKGQeYHjUhPBJhO44nZCKXzBTofMqSP9iopI/YEDrG
H0Ybd4iYsURV2juaChPE918oTmoAurc/ZaLX76PgjBeM9okBbnpK/kNOmUVMZAN0
q3WV6cOtltnzyDe1PNZZBotJQIiOClcb/R5JJeFKK8h9OMhnH/kWsiifjcD5e4Hl
0yBZr/LQZo/LsBjsggmwQhcP1JoT4X9lwQxhUzguwS2QZHiMRSirtAHosI/339X6
FbbhQapMln5nzs4kO0YoWQZNN5A1hikRcIpyyd+74B3R9bKfsjAet4kbO2xEvLjj
eCgALJXXnN+AhQ7aNbnNPmx+gKmzT+4pwoeq/iOFouRSxuqw4DD2iwr9u0PVTxIp
sx1wYML/EDxZmsVfHzRGGkznx3HPrSRkXNQ2sd0O05rvASV6mCJsrJLGJDrOBiQz
PnLX/FmU7A6xe6gPtXeT1RYW2tXCkbwMtUNIx92dBMsssDjeYTfeAF3XlxkKHVi0
F5GlD0ocOh5F3O3vp7FtU4gfAMyxiZj9aB9YaSAIY2X8L/4GtrkbA8oIcsAdCtvh
H+nh4EkrPP8ju4ZqCUK1q3QdeKXkrvYgkD/AZfvaGY3OT6RJMmE+DM2JN3H60DaT
MujFRDMYgq++oGT6lJ5RyaG7NTlbzom/Gbm8B85aZVYzgM1HAa1YCCKlGkhXO6LE
dA/00UPtTRee4f2yqtSxHZp5nfv1FNo17546hIZ4wk0j8u+JfZCWKvi4FtbS1FrE
bGqxIbohsc2gJzIYXqshVOJIxy18/DwSqrWzPjH6RHq5qCMwP6zv5qSjUK74/VZF
JYTePczM2zzawrpPgPVhoWYKqL5dDid6hVCNCzvCkOM72jsWqeHab5txZEZ1qAbn
wBbQrixWNaErWlFU5O0ldczlYBxcOfIFd8+I13QmVvgqW7vxNKOzAUlJ35bcsshh
tFcb3veHtauUuvA/7nGnqhzSi9I0T+paXhIFf6NJTV/Zw2NU7mXjZWCkF4YOmx2G
46LBf+5Ax7FqRBYc40HkX5F17seKD/Xeg+ydacIpUNQeDqbn+T/8BrBXEzgjqPc/
pukWWOsy14no4oHBG05YdtedVvw3lYaqEYe8r9SBXVc1IOGMTchT4h9lr0A75bf3
+t/h4V4xB4AJNKjpKJ3DHnUPYqBIntCEnpojgsY7q7YI1WY+SmGsQkDfGtyN27a1
sVgpxblnxaNJ/y8dmAToyytTk9WfV5z7W5XWUMYSPXxbN0aC6BJKqq3NemGOTAS3
uKs+rCzWAhfB599FwkYIrtrA3M4IApvRJduj/PTbhGiuO1XsUBwDgPvaw5pYMfID
NRNUYL+dbMBqQy2zGot4Q99xe1cAMLrBDIKxhXkM2PJTsDBf8WdJhDCjjUA00XBa
4eMFJ4vrimk0ShBm7pHSIbjEQPg0ke0FZKRePmpAsLMNPLOqaLrJ7ilB6LXDmFK4
BjQm6ctxrx1EEa4f9saRQbmtgJEw9xTRTiYxypxGYmFSfVMLT4SYUnGV1gQVk0QR
HKl/4l7JM91OJZZ/Z2Pt8N+peG1Z+1JelLm0i+aIq/F7m+mcxZ4T+azgUBDQe7OQ
gEFLCD42y5yL57572PCX20Ocs7H4H//QBccuNmo4ZVJWE2WySJqDk7dmd+e+kkQo
lJz1WiW/QZPCSeJBCKR3IsvS2kdhyaA6wO4JMnyIp23al2gapZUC6tv8VTnecG3k
4qAaMq6AqU5l/PingGxSDIO652h/cCRafR7HCu6wUDGcTRH1Q5WdrGsSWd31tGmg
D2t3lLkJOCKYruXyoxhjLRht95tBklTmE7cilEw4Zjfa0FuVdbv8uxLRiPoMrK/J
iZwe4A/SBFksoG4BnsbmTGaI4D3J4NoGcKbtoN6uDRB33XbHwqhyTr/Yg7wywCCB
q/SshdPoK5c/EyJ2YorFah0ep+RnHs/6pvEk0CHrpQ0nXNkX7ROMHyb3UcDCNHcU
9o5/i+1i3bRJwacee0Biuqu8TvZOIVlUvQWG1ndz56G5w18iM5dQV6dXthefZsgS
D9MErCgnfZ6+1cXQw4l3uUR7VUa+/x19AnZFkEwgQKbCPzA9RPb5TiORR8viTFPn
apZTueBGvCw3m8JFyBuENxRiPWlqE9AYW/CE9qldqKbSSdPdgz4pVIbTwovbNF0d
umHjUUGb6pJTHkfAAeoiZecTXwyhvxGjlaEISJKlR9fwnq38+INIf0ZoZhb4FpWZ
0WWq5HS1RDqmD3yyp84V95lwq5WNNLMRj1bMWAioHbWG4NvSMDLMq2KKeQd/OPe3
iRT3IvQ9OLumzr2ijxshTRRZS0EAyguXdBv8LiTqyWgQixAq3jxovvJ/ClokhZZ3
KX597h6T1JdGLpZArlrKevzU6hIcWbHUj1x6vTRFeIeHV10uNN/69MUvPo9atjwS
p/bn0iLrxCPIbAg/EiXDKxfYw4NfNYMaLXaWlBVxUY5DwJXyFbBWzZFeuR2jCtP6
YIsckaxLrGIM17h0TC+Ycn8MdUwR8qA093nl3y0ytj3Jb9iBNxMQqFLuHbQ9leQU
lmamBfF5Ap557sI2pMCRJvDQTqTxkv75IsbthGP4l7lXroTTeshzhbe5xdBkE9TP
y39Iauz0s2Av1TBU6zafCSeJNpO3V0BcWR63lWAu3TaEJQyUQ6hMs+RPztE0S/xD
01+I7rgNlCiUQDIGdNZJJj3cOqQwFzDDapTHANCU2sJO5nndc70Ptw+v8nsKcMwh
zUT2156QSgejBczRYmmtj8lnPlz7UQTpHa04GQ/+MhmE6g3Y2DZANydn4DJx0Zbf
KBNEryF26whq45tCNA6i5YHXTx0uUEk97eFCeCOJ6BuR9Tz9YZykd1bPmpR1kXAl
4Tncelr4p8WyjMxFB05IHoGOA4dBmvABL5mL7Q5ZrzSMHEXpgVJehLij5agPNfcU
/YOKFfTxV3AGbAa3cpgfIFRKrxN2P4RdHEC3krrDGaUV3+dhcI2U7luXlWeWP6da
8B2Xun9ftNRvIj7C21sc61YFvH52zY4BnCCptB3M7nSyUSUXxDTNX6VOv7yyBlGt
kzte8Jx6E8DEQ54rLOckipBLZwX+LJ9+oNIwm0zIphuWTwyRomTXBOVIWSWSrizK
hzGY4jnppNAgyHzqOffDeUPHdg/9dr3LN2stchVEA+sIJ3BVMQhxc8HIv0WdSl3B
hxg7O/r/PEtLXmtRwzZnTmYD9dAoecQbIO3ovoG2yBD+l0HAQtCcfFFipmBL17aa
4Uq6F/eCqaTQNDbmIWNmlKw4RMuMVuuU4YvDxhwhAqC0XTv5S4cRTCXq+CSmqeI/
s4UdlVpo+d8OvHVtwg1NojnT5g6OuDvXYdLnii7n7vsVOdBMzoCUttJmVupDqRyM
11GOpevsFo6n64PeQqTjiXi1jJ6upjTFnP935Ec9LAHLci+sGVrMrcH6pwUfgLK2
YPPq05tn3JovAAAhS+q156NOi3Y3UTW4e8nPkUoG7TpiFCywsxzEZvknGZS3iji2
o7AU+6Bk4CENEZqP4RgG6UlO+MV3kocSqATlFAr+e0918gP+gjzYT5x+1fwzoq3c
/MnS5DYm5HN4q+ilXOMmVpH/GdjSsgzxxU4KAMm4sYWW3WOnOKT/nj7IiOJ+oP2n
G5xNVDNEy6plOKyt5WNrE6GzwEsaooLVODFxTABM9tEtOOAWYS/0fQrRo1o1KyPb
mBUQKJvepgUtz/ocQ62OLazOLbsyV/8XMT7hJWoeu88ZUyItjx+F7o4pFEj1+ZhY
djWysc2cA83O24aYSpPzRQRydUJQs5ZYazuALicpj0ZjF9MZUw5p74BjGBuV5cXK
FX67ZgWzjTRpU+S6Y5BAPa94BKmPCjWOWy7rx0C6VmwqRuAG/HrojQUq9TKXkPPk
4mt5zyRL8M2jEkvdoZ0fSVuGDlgrql5YBGidbHifbZZEQYaIVed3mLvXGZ/Nxe5o
LzmSrpnP3ImGkkSOw/KJLveO/TSqJ7B0ndc8Dwl5FGO+TOV7JEl4g/86mMmuC7sq
1KQaaeFkelI11ngkofUiTXB1McpWXdgqtij3cWIuQ3MKNCvw8AGnGwFZL+rAN9+7
fiQDt3Govo7kgF5Y+jbC0EBW+bUODL0UUg8HB7dgEvMaFPMesjz+VnSDQqBQVL5e
0RmEjP3HYoZzzYzYo3fTJDvy1Eazoru0FPkuzGkCJd76oyzpEVen9F3oQyjMpRns
Zeow9W0DvAWFbUgX0K4MmJ+/I/hP/s6LVuTLaT06iORaHMllWu0XzNn4Fn60y8YD
1zoauB9SLrXHUTI31IlIkJgNKxrOHCZHk3T0e52v6vBbZLnWOWoc7a/uY/2MJS9r
iYxgaaZJAuGyVrg78eXdpPQkQWJoB7rIcRxTH1hja4SSMqmM/kSNvwFl7DQLEC9P
odMdBjQH9uoX0IwTnG1pZVF53624lPxBDjW/6ZgDMiETyzoYM+KF0EQIKdzQJegp
fnygG0D2PMQo4hUcN40SZN4i9U0HJq6Azf/2Ulnrh/eQ6H024UmamZmmGNh4tZjF
LZY9V4x9idJ3J0khJk92wY87+SAVm6SFSc2j/4gsvIxdZ3onZd6IucMATIhyIvJ1
AOAZqIX7VZgOsTkA/QngRHgd1bBZlbeYup+m1doywQ3j1rIMA7JNMs1smn6T7vBS
V5zdOG8cdztdUsRTjFnvqRxGO7eQ3LCLNzAqJV3/MFzV5qGhGgMx5nJZc7u55gUM
8mt24odfyDZdYHyAQ2Ee+a+HAgrJ7kRynArGAWkkZqXhZuEY7KIHyRWcCNm12Q9V
wVYwDUm3T5QmFBONPu431jlyhmyernms5AuKNY1ajwknsidff9bU1qcWrzOJSUjO
+e0hqlRhF/xekjf+8CDNVM4b3pRSc9O6ni7oIt5d6n23AEm8/Y6ouW8W3jiWINhu
0He8IGH57u6OI6ga9lCHpOsU9gHHpYmdYE1Nzx89iuT/ICPcBQHyjCYuxvtb8u7l
HGT1mN6uXBEZY6IG7JPlYAIanQfl8VJJ9U6WbSsVDfkqg9o0dgaGyB6ryc6ADWQv
Mi7GlaJ/dK3hSgXltWYpuA42xeH/BtVlFEvVdKiYKVbqwFSGbI8zKSRCIW8/xbI1
gBfOByAgVRmFTlGrqzXUZcZciC6sbXD6y7Z8ynQN0CfNg8PIelkUqB1pVi3HJsvy
uuXLwuMewXa2fWOa0K24al/+k4kOSIyaHpUODOAw8IKdnbzBIPbhjyZ09Sm7HGZW
CEl8aSHW0UxxkXiZvACoZqC0Jya01Jr+msjyLizR6CcHNiUArbaQDT3FOwq9MstO
rFnpMclqN/oIkH0zySXfC/eQmOZett10efUpHnuiGEnoHLhNQAc2ggwv4q5zGaLA
rGIodB506AIfFohp4zMBK9jVXYbylnr5eABltGhhBpw19su6Iw7f21Q0ShcStQmi
ETWTBLQDirkVU26usf9ngCdn//mpbpnT8YULp0/1JVYz7OpmiBQPG25DmFNPxWby
DVWFSWBw2WWWWI6WJoRNd9c6JGMNPdDmZDQra3Vif309w4IaUIBnoov+eZa9h1jo
33neCTi4Xw2a2z1omQpORPhH4zlq2aX2TM4XQFoOHHGPwWJGtO8Cp7Etlh7tKMwl
WlutZGgob7y5oidtuWo8r1hKK9hqBWydL9W9MSZMI2exem1zdooejxR2JZOHyNtu
KhiAnQ9mGwqngl5JtwMVMvwO8xe/oKIsXeeF06SAOY6S+r0xP85D4f7jCEUZvWOV
/wc3HSUJkcRsYMcqKHWMaVwDATayRkLUk0HRPOt7mwWfaOPrFDj/486XQEdMT+TH
AjG/1kYvAILpdyOxHsmeltLKrEP39zQvZF2IpoaUCgNEktJFc6dWasVfRUjPn7Jf
sodKiQDtj/+e5dgwaKHxQB+5gltIkhTnhj8eD6h5rJJ92DqA8e4ADFC3QNIs15ew
BfRtn9Zw6hLD/ITvhnMH7sLfOtWV/c/wTs1A36rwuUQM2cEaEX4aieqCqXyEuOKn
U+A+XOFfFM2N0qwFBiwc7ufs7HNEOoSCb/9YtIR9oWiO88xMMMzxPKUIux3X/hM8
NnnRnonLQNmwnEGN1nBdq4TUf+d9XhgIf3RAgUexeX3OpJWyHG5Bwqb79dkArwRO
gx3RYUzqFwJceIkaro/jgbZR86iGiHt3kAqIeJcLNdms1mXOjcfCCdm/UHZHlKEx
IWa7S6IknsVwKOo21FiewKvAPzBKd+u5LczwUVqCHZGQqKqCNmNzOYRkjRUXPjGG
lc7vtOCLJDk7Csuzvvi595MMhdO+wJTG3dWTyqDxWI4BAg65ouHjX/eBcL0ZtQac
eMAImkUje/bK/FOaik7YXOZCnL1KOML1xwRHssXJr6nXEhJsYOTEw9y6zIBlGm74
6JJpOUGN7oKSFcqHDDjVJCHg/BXjDwYguRhhPYCkEC+6FW70K0afn5nbhdDmWdwL
W686A+V27MZIyx6qOBKal1g5ly+jgSPCnkvKgJ/ROrc+8dTI5SPN4sBibSx32j6T
0tjZy//ieRiy/N8tfm2YN7QIx7ORdPk+c4z+lQFeFe91/nyCMK7g2yfFaQAbBDoa
BhpdUNA3Th16Aj7stS1YDSwcG9K1WSiKCmGeHj/8Lhr3PRa4ISZgSJOiUNwZHxaf
TwvwZjAv+sOtzSQCzshSbnYxuj2hUlrCMq/s3u1xzIg/uLwtEAgrLXtaNuUa83t/
87+eh7Bu1V0nyIBGFvQJfdZNN2O/5vYNuqB0NseMW5W5rCWjhrfea8F4n7/xmRuc
kXV5TE98wlg96krLukqvAsQDoKFNF0B3M5cbo76H7jsuJm0GP3W9vFHsfMSMeqa1
nQD7CsoISRV8MhzP+ZxFzS1li48un1/UkpkqZgM1HQ2dtTvVxr2d0lcE6cIeBP1y
qmSE7Zx907TqHbfOwwGEMzl2J/TuNZ9sd+5WPyhzWNdbns/VpwV1+epNO/w/8W7a
6SLTi8FhaA1UuewNDql6FfZBaV4yjgX7SBB8j8OCkJxtvYjEuBSiXfLkDGPOwebH
VoZOHCLQN183i/FyyWgG3sEXqpJ5VAF54QhnE2R4q6ucFwk2BUwlg2ZO3L2HSsvi
VvqiewboisD7b0u/ca1WOosYt7JkiwIkazBUfcZs0pCDVCaz3ey6tNPVzwy47vSD
i9Q8KWvRiq4bY8sW+qyDlea3STp4xGGajTbMAHQoh6fxwmilAY2SAU8fPsRQXlXo
/GXqspY1NKgseokCF9C99wsmsaqhSzWmYTjqH8nl4v17X7OmlYS/5gvItcPcUR1o
SSvoGOPUH4EMmtEJzzyeqrPVf3yKP/uI1lflkjJLej8=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
OiT2dQb4Uy/gEdqLMC8CNqlBJV0KUNAMS0S3akDLWjzWwgpbPMAu0ohnbS/no7R/
zVzjGshZzllMwVv5CVEgR7vk10gyZFhDNyo9eaEgAI9/3YDHMnaF7J19dm1dRkU4
AgETyH3eMKzFNTWJ7pswRrj3XPIA+Vzv7Sr2/YzcArTSEb4KTD4QNKknh9fsJTwn
PUC19jwL2HqqHU/YQ0j7sC3XmhN6EX5Z2e3+iIXC9fx6JbKZzsTQOWqXKQxkUFAD
HakyLs1uEB26ZWhUaB+H7U09XlMv3a8xVJyGH2gNcxzusUr6F5EX6MKiDAUdpFiO
EUukHV9hH3L3Kj8uW2xwiQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6272 )
`pragma protect data_block
6ekKNtJj6LYtfU241tblmTBY7o9zRxMc6StHbvq8muSNt3Dle3UF7FpYktUorwJP
xi2XkdYcciIByQ25BFOhB2vODFe3Z5wG+D3Zv9KElE/aU9mTJMDfd+4kgaQOKOQo
+LfkxPaDqu/Lx093dHiD2XgRWe36dwX2e7nyrbEGOklIo9/EsQmu8oPII3mDb5Rv
BujPCgd/HssNi2thL6L/VEU7VgQzxtBq42NLpoMPoL7joS+4kQgxlILIvhpft8Cp
glgur6aVTWk8zsQ4sBuTCQu1bCsI5BlgP9FTcVvIye79R4Pd+lT0DxQ1cU9qI4zM
cOs7FGS0jmLM9KySoK4QsUgCMHElY1CeSlzpacyjSTLRPkgHfB3byN3Z+uAwg0rd
hG7eLLinx3PXz7f1Cy+sdvNYOayzmPp1lYCmcMegb2zZjs60+VcO6ouwSjae+C5M
C4MbVy97JqQ6TttTkHVknnLVuz5nHFR4mA9q/d2zclz3Ea1gdXj5zY8x+WvwPaGT
cSYd3HATEpxeg/vZAuxkabS9YD1Z1dv0YhGqcfoAbRBLHKrSMe3iKxHzefmMytIu
pIG7uiu/cAb9LKHuO7RIUV1cAXC5VzXfnKX2QaXieK4YtuceynzSz1DH4S8gAZfc
GslYsg0DuG+lm7ZEhjKWrzEc3SKOLPssc9CdUrN3ZQF1dr+m5wy0r7UWBzoJHmlM
acMQrusOIJwDpPfEZu4Iw8yccFEuWLleY7PVuW+w25rM69BP7gE6983GiRpPO13T
Bzsdk/S8hFl7xRGfZgKsXl7G/IIPdGjb1r0FY4dqD0HjJEtAH1wqNEHvjFU8j4rX
JUVoe19RT5/zETDzksqHEUwkF7I9kWN86PS/MTeirPB2joSUphPn3LeCrtoMfPRU
MK5Ow76hdwKQeLq/ALbHRTlW1eTI7T3W2FaUabN8TpXZSZXbC9blaQxdLJOx0y01
eYOeSRWerTVFcip+1dwl46yaD8gSP39/Y1+b7XDd3nhc9JBIAZfcKd6pbX2gkWUD
7eht8tKcYdDgzrILjhD3bYtxwWZcZV7B/kXlPgENWTCiNMR4oVI3cNOOAuU2hJha
PmI9phjiVn2C8MobVifVmT/RDRLG9XHqS6UiErnWolClaM4F8H1bL9lKja/+SLGu
SWq74tQMf5TbesDH5erR9IL+VVM+fOw9DlUHWm7j6NdJcW5HIKyWI21xrtuDryHK
1m3fkTqb8p0S2xxcNdwwZlLyFiUql3LPij9hd7nhebPgUGTNoQWnKUYy5vlyeP43
9yMFJp9FRBqWxly7qpGcLJSz842zxdGfUh6obwEGNFIkn8lXCHldlQSTNVk4yLNo
cLB4bymk7Bn5mctb3mhHc3y03it5+GSqkwBYiViXw48EyjRwtPN6Fnd0S7ubiAlI
09P+P+RejaV8IbFyQjJyRDCkXI5ATPqhZsdMLkXK5pLRcV/C+LAEYBt2tKBZzvQL
faetDHOnsjfCWPyzMS3w8iJx4CnRaYFc77dKD8J4+KH04F0yiw5IL75CNb8XCMxQ
viXqXHRh6DXwLdNbzOAE+3+jDEZKN83iTX8OlOoT5FxJ2Qxoggud0yVvN8byYFiO
4Sby37ljCJ+X9ApEURdOZ0Ga4FxqpG7KIGm6XvBUdB7ZNuVipgs7dOvdngr6eFgB
dxsMF1S79ITF14c0LNOdFoOI64PQxFFoco3Dn3pK/mdT5yePl6ebT7/INBy3Zykv
ohBkIbqO3aA2t4xLQoTn1daaL01mQy03p91Cy6+5/yC4NKKwLRvF6qZtWuVQ2evQ
OKZb7sl3eSp9zWmVXeY3Cq90uszQhU+1cj3nOp7Gxo9pdxJDU+pNcSHhnDWQr4WN
gW9+n0ch24mETUBMRbg5smibalCmhekuZb6xFF43+/ywOBaH58qI2eyHvcDSs5HY
QnpxEJU38pZWuKg+swGAb4NJPtL97DF3PhdzmUrQxkQebcQCkMP161//dco4GC9e
FhoNZBB3D/4dus9LAkpXtZAPK+bu4+U8ryWn3QV5K+UdWsgb9RqW/BGvPm6pZgLm
CvFokl8rQd4VzFcPN3qbrCZSl2tnBrYc/j+sHRKdAopMeMV5o23jBN0bytX+KCh5
TRQMSPkVeeJ6VsAkWkielsw0pNBd2A0cQ5JFLf+13yrYvk9aZ863x23/f+5qPZyF
3ZIiYytUumhzk4iR+8aTfybrYYwgDjy9x9jG5Uso+SGjvKQUIr52S4nCefnUsDrR
2+ojVxjgVuEkp2xeOqCrNBIMBIPgMMQnF8DjQoDDIgMKFwV5gO+1r7E5TQhSRPKO
i9f1oIig6Tlf7WrAVfnIe+xEPCJ1YLshaoTNG30QPNFgv577rOOXHg/35+DMw+ab
KAlToioogw9879kHP5SFy/wjQR6Nc833l5BUiIGAp0ovqLitaugH/O+yEB7U6sNg
oZwqbN/qLWGVlTCBnPemwVkcN5HOkzFOWodsEHqpJNF3QWGLHbWqLDjaXlWbyUoR
w7u50MO19di/U7k/zpAqk1Tm4GA/ZAPf5ojdUUeqeKKGoPqHSt8ido3KW1Jtbbmd
W67VPjkNq6g9QDxomhLHLKhu+89atCmAlPvUwXKZEa8JWTtzf2hrfMOHXkjc4YET
ldZs8gi/vI4+rLRu6ssdVse2RHQIYVhGjh/FMN35uVWS3U4MbsM8+5UVxnUC53Eb
fmjepQ9mVdv74Fug/lmgXVzAbVX2A64Q9peGW5tnXB7rD/7Ov6ACWsZDbvwtGMBp
kzHhjtNYBEfKuln0ijsZWukPSm1/xwneIlYYlo3fYOGWxntHYaTk1MU/FJJRi2du
IeHRB4B3OBRPTjgCnxWCtJQALkGfsmxbWk9FjA+CxqqMLTHoqNLgcAXrAg0PliLC
pUf8NfkLF34wcoRONXUazN40z9oqynlZmH5TusA1r6Lhqf0DsDeqvawcoXO0zVYZ
2WpysPSXmzJgNKW/g3vk3UgYX4nxfyqi0PsweybGc82TlBKp6wpy/24SS3CTNXHf
/ztfCHQrC0mkUMYD2Ujz8YLJdJ9sQ5p43WSRIVQoTwYK6ezAsGN/9OEY/d1IUiAd
guBc7iX0ELD2I8B+XYA4Lq0YZmBHOt4pKAOM7av5usHAOkuufvRrwcnC+RA87ss3
wtDvjUVgcL73AWCjifqeD5Yhpvu0b3hnWY+bKpowlRIU8at77BWb/g6cerexAdJz
sr5jT8LisVGn8ZO7rryYjJw0JOCoz82jZ5ld1Xx5zU2H0tCIWl/Y14RbLVDTnUhM
zq3Oi32ZaSJ+t3psjNjnGUtnr3RXez+kFSZz9gZ7iCUKPfruUAC4j527yNAdPQAF
ZdEFJ7eBcp2IQHDBHUYzu+qeq5AZDlUkXCvuI5qXtzJWAIPeiv/5kL9V8cVg/HBk
rOqdUrPUcw/+by0+F2HKPm6Z+9tBSrPQNhOnO4M4ChmMumIWNnpwFxG80qapbbFb
kbQaWhp6KFBhU6dZjoc4Y1B+N0aPLNrfvjiwNiMO0D1z9E1R5VHKUPdJe5HNcCcd
FUDhvoZm+azNSFNXcGenyI1SRRFxIErG+GKRUkfbjymTU3RswGWi/uAsN306LrRo
HfUPT2dpFCEuV5LuCduVJycIz7M4VMmS3D1MuVP7uIaeYOgQ/ei/Q4VfE4JX5DXD
lz4ARo8DAsA3kyT+ZBjnS3kPpmySvfE5R60mnQW5sIFrKW7HjOpmW5JvNpJpGLcB
Z8dc0NSr9e+cICKZsBqq/ooGGyiZjjLfjnicbObs02LjJXB6+JdoJT9aYYD7E6mr
nT47HECFlA/B77Xi2KlJRM5E8r6hrYFzyNh7dxUMpXujGuqFEEQmfZvTiPg6C+DZ
roMlirv/jIXGYYy896CDkDRrZZhSKE282+9GRFgiNao37bWL6IQGr8RUKKzEFxNL
/lYO8q/ozG+DgnoBQDY6HgO5U4dqflFzQEjHaDAgUGPtOPbCAa4xWcMpcMkYYBSZ
J09yTvlRIQrcGFe6agDMGZd2PXjWaZXwye3Ojc7pvj12KiCcelFik2HkTPG15Un+
eIRolhwEBVHE2sV8VDhCd1nYWzi8nRm1rhirdSMXvHfzv/Ug05Xspt+ZCzBBsHoZ
8DG2xMXPIzEG1CHKYBnRZm/zrHVaEEa5CJrPuBOkc1PQpnnAt7/1XsJ6rQvzc9kN
+56aLo7f1fIKa/YmX43RD7gxKDvzZJfkbWhqZP9Y+NzpRNapftz3/neBODqdGp6H
TDxfA3YADzj2ld1ddUcvvpjfKeIf0x6TkD1VcD72LGBYON6gg+dAPM5hTP+7zG4+
R6VmUowybnndduqRn5GCir4HycCwJKbUEI7ti0MYrjuxIjTu1riXHMsHlSaMJaWL
xII9e3hOz+1DLa4va9xK32MOT3uReFqYBLuuAATW7pshuRtnaAm/WQgCqZN2ndye
A/g4+kh49WYtPYsLep6gg3SfD6vi4++fvLuWWqEN6/RfZ96oY3ZQ9XQezPz9Qocs
Sb/+0Ke8Chn0j7FwEL7NpG7vhF4qn0U7VuKTsuEz0QsKWs6ufrgmjkLsj504aPd0
IwPEe9b3iDlB/jkxvgEHIe+1LsddXVbcVrTPWF4VK5pFA8+ruv8WpIZqHTuV6Kp9
N8wz8xZaTUa6mdfMoQ/LXdVdGMMLsRj1i8W99vF7OCwEPBKK9YaR+S0X3ZJTHSRg
qoH1XInFnu6/1r8pR/ImIku3iAit/CkaL+HQhjyhgmef0GOr4m7lvy9kPLqWGsLq
EpTl17TAqK6BvHM0DTjHfZfQEHz5royCXCOh5den8FqW2LwEWLqyIi5L6zBTG7gf
cOdsbUBhWIL635Ku/vIGTXG4jkIqnU8bzvid1CIcSUtGyd5bhELgWYfI3XUS6vTY
FnKDMU124x9pzGkkCtNWHpK5aHJJt+OD9Uu/gzKA6FppdGFQkBaHe7YEyQg4erFo
zAcTMN6IrCNzt7eYbRApVz2cgjUjzlq8lymzJPgXYyqICl0daOSuWVrS4675g2Bn
IWW+Upyze4zPvSNkMvBzznGKdrJ90Nhe3LYVMH+63MmviqrAxk/3FKD34WtR6lFH
MHZUOeYhNgV8vR5uQ6RRgB9hpsAC+PP3f0dcOrywxXUEF0pf7fO2eZ9ER33AEbHr
2hPVwIOoY1WlDea82IkNEvyWK1B6zVvjsFuO1xTrhk2YfsK1FiR7zhRgmmpttbd1
/ZqwFZi344hcDAWggevU8sDi/jl7l7j5rgOJLpe+eOvG1G2Nz3jmrQHNqzQDrkWV
+zX/G1KoXPOOgOY0tfpKPnc1Tn/HYQkkY8l/7bxr+hWLtbPEc9M2c3UdDmBA5Gem
lRPufCof5Ow32RzTlMOTVktkHC+KJUEErySmXgCJR8DdfcmcVr2SX0YZGjNzhswk
sU2CwnA08tE6jd/NQ6aURw2gDNcRnxzYa1nO8VPDwPiroKuS+gNXcMZIJxoG21iy
bLTneluBCbeKZaOceRT8cnjov8i8TApg5rSrtIOiUngYxpdsbbRKFwckPt8fn1AN
aFR6hP6mJ+9xPD/tv/i94AD05p1VRAZJ8yj3IXkUzk7X2gKAgIxS9h9oJvyBRqaD
ajzwex+nlT0R/mPacFFbxATTeRlq8LWjKZIv3AKqke+GsqpQFWhBV7WXTq9lz1yX
7/Z817YnPRyz+g4sTiRKBHzbLJapvmn1WiUHErlYWX2VQFmlSFmwu+px4Ose3RUT
HZOeIJF1owiiQDZ3a4ZokH21hvsTvEE75hZOd/uyYJAnbS6PYbVCzY8W+uzbR37G
pJHuKz1SIKzdXT26cnOfU29PgqyNbcIY//yrT6tztGqHWhc25zBPC7NgclfT1q63
TV63vbluzgkwHP/dTpSZJOiibOcV0lMr9AZRaHjbICvzWBvuNpvV+DH/CUqeDxqn
UoO73bl18GJzL97DW++Ya9CGy34V4e8FoGeNi4qrBUJFi17KP7UI/P7wsPwvaEtp
7YNw0Mi0WBe671nLSsx97OwPWFJ/ZOhact3Dpf2TW7mzWeihwO1jirgqDhgmRVJN
1ADLlDHzZn60/KnJOqIka2x3AWq+A2tAVnnUHlLv552IFUXgUmIc3PShr/TcbVp9
YmIYjzyDh2jFd6t+yUvIeJ4BkV1rFv9ASQmzzRMSVyJ5Nshi8V4P5s77JPWY+N9P
PvONq51kQSuRxMvO0lqMuXZTFElh+Yi0QCOMPtFq6N6F+Cx8JsQUOTIncfumaoU4
59NlEz+dlTjRZHx/nDHu3H8Qatci8Yc+aEqkdGYuWai3mzSA4Gc1U9GB3LhwdROw
IP2MtXzh+WYSlsTI6ZZmkBDZGGCUjClXQqXn8jL/pcp8h0GKrMNjgZ2jc3kNH0VP
dCWGDD0k9yzhWItC4JPJczvBlmmd6SduVu4dXU3bTNFXI+4oH3n3+PZZZmghyPsV
E5kwrIL4DPv2U04+8/31l9ugNK4sFUJWOdOQ6O8/vC/iltq8X2yeAmZUMx/Pmx6S
wSuuhLBSXzEHdzJo2Wz8z3Y2ZSnQLZjaAJU3lYeOWW/Y71Tgmfsdd9d1X5OVSYFY
/ouvwNdqfXBY4ihydSFcjxHb1SGNdNjNpBvYWZNPn5R4FtRhPh14sT2T9Pv4sXZn
UNM+pXb+cd0YkNwHVOBvOJHFfWU3DoHy20swLbN7bHyOzOyuM38xtyg1btVnjrNW
f/JqBSm98rALkTsHiM6vGsueLchPd5SCObVpB++vwZeWYqNxezg5qRXV9M/ENgPW
jjx046UqXF0pGSLSM4NHwdtZDhWQqldXE72JCzyex8wNFOjIHooc6lEFl2wWGFbS
N1DtP2MF8Hc2EENwpjKJOautfBMys1ji94ZQzUr3cmN9v58hQ/DPIOkLVQlN+PCB
52NXJGPu70ifeFVduRkwdqRaSXB1LMwfaaLRe4SON8VnRlSFKKe5Bf1hBdBBa7/B
z6bUgLgyCBvZhV6jSXTxx0iMvmRXRRRY/0adY1DRrB1xI3yB7VWJkXN44EF1wfih
eyC9+mhBokcjbUuxjLubtDXvMAwqaWbw5Q1gwc08JcHgtjdJp305Uq5UxpWLJXt6
mg6CAzw63R3x93fX/Y5BCQ+VIDX7d2Eu/Bgw8GRptYMJRQxsfbadgVTWXQtAgefD
KTWThW7zq7PYi57PgeX+VbuzN4gMoKpZgR0LaBDBIkk7+C3b0VoVRZ9Fr1X63Kds
UUAwmGMk2yxtuNnkJhRUlno59ME4CQL67LD+GZIrol3mhmTK+f42l2F337gSrgKA
r2/2bxkHSAwfTQ836Sdw/kR8Uw3oa43QwlF7xs8pxsjfoSyGTFfvrvfllelqJw6d
5qHtXqzGS3dU69byck83FMp9s8RXFzKkKu8Cf+HkWsGX1UOkNPAv7I4yCAm6wzS5
/BK8kTL99OHGpcdFR+SvUJtTqpVMt7nlU/IQUUe9+hHZD2QQJSoSd1AzE4fDrKZH
zZwDAjMGut+QZCA0z/i2QhYmaoJgub+TDDCA/n9hL9kQcarxQQFlMibdSuupwUUY
1p3lshR28BT/vktJBDn54MlV5+6fAL2M9Qx4H9su0hTELP/APMHMUcdjNkRww44e
mH+Wr0L/QRjcHi+QRP+uhA19M+64Sqh3MvrwKWnrTUPfdv7Ai0+dIHIrDLd+CgCm
g65DqUBEBOYMcvlOx8k4U4KTLDu7O3XGjAA8OMm0DUxa5YwP036+oysWdHf60j7r
Lp79B5PfiFjP+xmE7a3yy1xXpiNst1OaHHxnFRUE4oK5QGuIHmo1+5Z9zi3OoaHZ
ekPojVRYW4MWE32Y87VspFZZRMzyGaM0ZZqf11cP+vGyHu9ucTAXOkO/poOdnI20
RCBMmDnpJejJADmoLzQYpmv+uv1u/rOstwXA+/UKLbcsWoK99UKyf1FYNIm6iNwZ
mSezV8UPOtEdkqNhd9EkbI00NJdT+tbNYIctzXCODVNa6Pgd8Kl/UeHtMHrC+lKi
FtvvDCdJwIL5k0pYOmbCer+ELHY5uD/euvgaQZnVgBVK86+7OLKA82VL+ua5Nf4e
HCFQiveeLZ173EoE5BHqOSVmSVt7SqI+ErVR/4ExET6n0u/EM2OjouENfzXuE2zc
IN3L0g6NgMDRe35/DdEyGF/poWIN4cBVeT1VtCH3AzamvipDR/2ARWR7CVoI8xjp
s83dV042TyFBt9XLeVAfxiqQ3UR/wkRIXv1yfbRbIk1kYNw9VXUqlATmT3mxiQhh
2u3xAi9OBvIA78fpHgn4FQw4pXj+idAdjtyIHOhBNjgK8G1Kdjvn5beXZiP/Wllf
8MNPtCZwdQup5HV1mDCExgle3BRaWLsPFgHYA3n36Z0/zx8OdjwfPM1pPTnpmvOb
ESokQReieUyy8TCmRXF1Fsg4XN9Zjj5wtaZYYDA7yno=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Gl6v2DgxXnZl9eb8DrAVo5uuVSLeXggrTanHLhJlxfbs8E94IyIfvcRjODGoz/rg
n2j8Gpdul0uwFSDHJRC2VGdGU6qhgG/ffX5GRHgzYMBBq6dktH6Wi6J5kDnIxsys
ht4vi6uFYOsAZW1PiGua777VWTixnsQPsN4Ctql/pPPGpKRenm79ICjNiWoogsEn
cZtbHAn+4UOSxlDz/JdIzSY4F8EKQNyS1vDjGPhKBy4JxPXYy005O0XeymAqLuRq
488oNTRET4mt/mvfKX/mzNkfzGa7PICbLJ6Vj5pHrfpjNgfz2C0zesLzFExLShSd
G/MORZ9kDIIcwAIO8IUOvg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5424 )
`pragma protect data_block
vTYTUARxAhzbYAgX96sZzGNP4FOjaFGVafhfhVdBwPLwArfGV5MOcfAR4d8FCQ+l
2VtBqU+25x0KD7OH/xGY68/qNUoczWyV6Wu4q114MILOJ0FaA6E90pBM3q2aRLhs
gNoZgA4+Veal3J3PgBw7lk4S2cQyLFc9cf2XCPgB1MNqyc9tDS9NQkgBuCTUFtNr
ySg2rOR2e5X5/JSdln8HbrNz/I4BTXlzyqgHqxNhdz+Cu8YlZFDfn6tPn/dYoRyH
iRWee7Gp5wxv8cB3N6Ao3PPluXwj6e3dfbKGc8AfL36ofuaVFv/b4bEd+1WuIpEX
53bz5ksbe5B0MnCbm1hai5BKVIfi4zKdvJ5BDblEcMQNovS1V9MUU15v1Q469lw3
d0n+k/YXNKi+QYcFLKN/pGcVpl6rD7VeURnhfUPU+zYungxiSM27ynJOXe9PDSRj
gipVmxZbc9FZfOeNviZ/uylek58OYO8QerYzpAp/sjFSEVsG3UVhVMzQNtCFGCTS
OMygf4zUpsBbaBkfraQFCfsOK2yxw1pRKslQFNgxDFuFsSZmeTdkQJz1LOV4hGy7
cVxhuJ2ezBO1/BAHJhpgQiuWPeJDGtxBaV2DbsM1LmRKQhZ6c1A3fzl89fU4Qwr6
dHh1ZvfPAQjEDd/uXKkET8T+7+gUk766/GXiSiblirsbnm9sDNhKb6WUw7qST6CP
WTMW9uvOmK2bVSHDBciHQ22nw3vNck9TMTmKKdP+QodCA1ehwmX/lyu/aGzebPDl
kflwlEYk7ikPYUXKTwZAYwB/cRq6hS1l4KskKF/D2aMOCtKEBwh9N3USIQJg+cVL
ZsqI6kHdcDwArHxVSd87EGbF20bnXRTjF2e3i41eFWCdahpeOs9Mvorbebws/Yd6
FbpJzq808QTgzjbRAdxIbvFSoPSSBVYvzav0YFM8f12+mqf2hiqebph1G2fMybIe
3OxRAO6z5JYcUd9ntGjy2saHR86FbZWPEc7634/Qydthoj3bltJvE1tEFl5gn2/U
B1uUZCBdfczti9Xp0LsDfeO9/IGN/Q2KKvpc5sH7vGDtrmgzbBJ6zfWaE1d+XbWy
hK+S4y3EZJx4vdW9rQk9NEI4Pvc621uQDaQjt84RfyrLsmO16xfJ3Zovn2LohxpV
K8k/faZnbxOkB13lgW4GGqxKgaMP+3HyoiqcGPWId5WQoqskgTJq9eobyfq8lPNz
nU8u90vmQYEBTg8SmVEDOJhfUSHGUpfc9vqZJEkxzSaQkC1MURnb5K4k6BhXH7x0
HBoQck/V9bybds15eZ4dZqXNNjRiyT6e8ZPZ7tGgLwM+zyCzw+imL/yHmADTTPL+
Ht9VXkfSAhZpdyM1vz3WAABf7iJEqyZl8Zb9sDGZg4fBzAcNW2Sh6cmK22lSUzir
soz5JCRB8p5ips2GUKexXJiOSNFYu9xAbxZAgBMw+A/4lDWWe4GlqdDY7gQ9qwj+
sR6+50EBwIs7ibHDAK6QhRZnvoDT4Y0WetAq+absLxbF+EaEZum4E34+MTSag+dE
+b+7WbPySIn3XSnzOK/JkTuPGuQ1pRX/FvOG9PV9d8ra35SGJ+6ahFR7Shhj+eBi
h0mYkDge/l1Ixze1Zkww2ozFsY2MyW7//iJFDLwCIzBYuEVgKYzmI/ODDRyaxk0b
3y9mdWFWOtN2DaCyCmqataHtPAAPtoEizjqy3Md3AQ9CpPMz7ceLHA5zHwry04fB
GCsPeQnbnFUjG10jbNPtX4LKZ1IQ1SeVnKFQvU+6pM+jcG8H1jzqTHrfoO/UvlhB
MRNn+DODxvYlI695S28YliW8uDcN/8Z8fTBZE9gb03m1ivbPvPA0Xr/u1pyazjAq
kX2bgDH29Ko5AnvtoaEDdzKGAppj4O2L2Iu27GdWtmIA0hlQljGb+bOphbsQm23E
tWmiKllgkvsPsqBLwIHEb34yO+U97xsTThTOdCoR+QWV/aGBUIfOZPCj9vQJrP0P
NeIyzgGlomaW7+KP+fQW9mv7ZqpCiPiaZ80t8UtCz92zfMqGPBB8d8sus4tjs6Dh
ebhQVQD6vI1Lp8D8cKuyk/dFaWchAbxJ5MPnrH0uyv8zIqFLJsmloeQWwtyf4i+t
xIYwhdlsSznZYOqU0OaLFw5z5zkR92gHvOfXZfqO4Q/6+CIFhjD8lEommSUa4Ra3
Bnfh/6eC9NATo48PF9bnxusZABHeAbH6t3JpIdrmj7xe14lSAB7mppNnRMrSjRQg
TJe83mJXpA1lSqnJwB6Yam0MMlchHi1H/fQMh9/bwWth4xdZzYNKs81Zx0W5m3p8
7OEKdYD6Jzc1I5fI3u5CanFG29ZSCpJF1oGMAlTSWuEghZuTZk/6hYiMHEbleg8I
yHjRKmQ8VkDZ79TTqihSTs/9EJrgelX3sy9J0WkndJPM2GqHUo+OJtVFVmr78Mey
kPzsKGN754xvAjiuSKBRFUxBraIOHbXTkCPkpAHbJ3ltjgScq+ewP9zLv1Gf39UP
X68FZGibT1g7nkU0WFqlz2d0UFXQ8FRwVe6GlRI3ngTkomRi4/1Li67NHcA6IF3q
TyZ+8l9OsUByNM2PiGXKdpCRAl0MpTyuggCkppNaUFA488DdZybHMKk/npP1bAKl
IOhBFNzMq/n4+O5AH2+RxmyhnBncHfPmaO2JKHx7paBVpUlr0C9ow9vKOPYrSct1
FfP7ZSanKRX1q8y0twv8byHarynbohd14231lcvSNwizzrOBPu4VMbQlNdvpmZ3D
dxiion0WXSGKJrTL+mndAmJ5gASnjrS4tlArzkNuE1AkQrxw5E2LWw32EfiBEoA2
ef6/+58IGnrM7x/eWb4A9K6XRKCM8kjhq2NAPqcuayTWGhQYVJkbjyVbyHeizoF1
EFQ6H2CdHceMDek71HhLfoxNRKnfmxQ4WWmdHDYsoEEK9920OLusK+6bV49BETUv
JU9vptu4TtSFvj58U1yM+e9QaXV0wpRsgb5+z9gXuz8mSE3TonkAK5an4c4Xqmer
nrFblqEDp/jTWU6PtCDbDH22pxt7GYYT+I2JDNJCoF/wrgHB8lGXHC8L/K3VfX/F
Acb7u4olmE4jipAbrZhmoAApoX/vxkwtZWyPhB1Xf9oVaf3pHmfTbiLZ75N4E/SK
EixljQ3EfPmVoDQsnLwlnFcC6m6TSEp1eyJa43GjcvLdid5/yTMYJwWFDh8FANO6
swSw2oEcJQGy+Y8FYAadME7+BriMikRdHzou1ADvH915a3DaWb+KMfxFa5itp9yh
dXnqWjKf8nsMXEy5c4X+SOA6rbPA/2Ce1vKxY/4ytZ6ZV5CVIWSOPmF+6jipNM/N
Cmr9Tf6ryK1rDE6yJIWjqMTGX2PzR7GoAUrLlkDXlpn3HAKwmi4njIb+0+RwZIte
xclnM+MuJDFLhKNBjDGqF8aYWfuFDxdvOoWO7xRs5Jrp9tGxLxneQnwhF6K2vLT/
4wPCABTcSloelFTbPcQQiBd+kP8qECEsk62ZF86EMIpQlVJlRExGdRVqz/dY8JMK
Is4yNVPEZ5Ro10vmjV8mHCWcXNTxNtOeF+cZ9gGiMYtX78iW/axx97XE1Fa7qT6S
BX9HqyaY7xVPFhzyvvzgXIXNrEA+tzyw5Th0hgkHWXUxxSJQxVMdE5pJzVbDY7Ha
E3pE+AR9xDbLjssbgcuOa1PoUq1+KNCraGrs3Yg+HYoPs3HQO/RP0ud8wJT0N9k9
l1XxWhcyQChjLA/9i5gJ7jizXWnsRC1FJz7tj2CvVmmx7wXmq6GJferZimLaJWM5
GLrJ+simOOrfdmjJWZAt3EV6540ZiTnC3MtOaaGJuHBXKrjoHPemsFTOnP4/escx
1SCNqB5y2kDOxmGTM3xpVp2L5F0klaLXVdj0i4jUrKI1jmcMm5md2JYKsaf87CDX
R7nuM2XmE0a/QeeNlFTx1q9E/xj1j5HRx2JR/x5eKV5HR4wAil+Mswjb++H2sm8M
3dSIUx5e6WydmbAx4ItMd7HVdnTn13+Uz+BBtFwsDNhSAnrzhd6RvO6cxsQtgKcG
U68A2eqZ4RDdV3Rz2izGpHC4RSvNPhEFXVX3x5Xw5VUdvzDpJWbUCf0R9x1l1Ozj
N/aI9eWClDnOxmESemo3tdq/IGrIwrgZ+ZFIt4SyyZSAN2QLYW1GEQ3FPmeXPGoZ
gQc72OGjlD2gVXroTOtziGiOKc3pjPXfACveg3VSwG71rKd1wLWi+fVu8M3uiJeV
x64MeDQ+SCoGc/PnEULqbxRAD14P/wGzqwy4lRhL/jJjU80nBqiM3hUPZTxMx5pF
tQX0YT6dVzjK7+bRuMe3llI67B2hqULjg1i+tWPwzt81CG45ioC6uGFlWE5BDn9z
wJTlj+bDDrgMLiu2Lh293wlG/KZ+DVnhm+a1l+jPYdtZi14AseNc/VnYy+/IZ16j
gcgcIzLfEUGqVENbA6U3aHhaXF/KlPlataemCgHsAMaQ8DED8ifAVPeS6Xzr+Bna
IfLw1viyCdLRAQRfOegMssvSbYlaG2OzUEJVmTehvLFlbnihmqFhMdx9rMlgYrLl
LeEF1t7ivx6Zrt21h4GmDteygvyLw+Acn92NfKf2RDf4YTXrS0Ag5sxDONKOw+tn
cNLWK8aTbILs0mAWJZmieG/LR7aa/1aVlEnFHWgdxuUGH7wesOlVhsnxZF3l7JRe
CeHa1JCGRHwJ8c2yDIANgjSIuLMdX2xAVUcZEnTVfXhpQ6llQVBakA5VdP8Qegxg
EyUXu4KfRVLwQz+gDWSsIO5RLKqNqdt1Y0m1O6ShTzuyeot3HzZInb30cGWUsjlE
UytzaOvJ7vBlG6kHJCfvTJX1pFQI74GZ2UYYnZg4m0WvS+Cv05K7iYsbuL3SPG3V
/OIWZ73f9dc0tVRimDs5ImCxH0+LEV7tbkavjsft7N9SwETWnAY1/UBc7bfejkW2
3m67FqMUbcvyiIISD7gypFVeRu3rjuxuhuOxl3vKqj6wJ24ThH9Y/oMqVBrAlmea
Diw2Ln0C/1F66YBGTpwj7jLQqUJb+NnnzOM5rrlhIYW43akLnQh4IscGOBcOArSW
yYypW/i65NfqnxVH4oLxAeXX080+wJmfY9ln82GIzAOBwqAGko3vhDMQzifXhoTY
dyzxFASUCaNaCR5EbO3nLmeGHoy/JiSPVAh+FViQLS2BQ06f/bUNV/dZ063GcTrt
iyysLg2pzaIZ4M+1C6FM+1IrMj1Nedf7cRzJ5RnK1LXB7QVAdXpM+1h9aktvkOMK
6VvDr9OH57TcSCFJMLxLoPoUsjr2wj3Q7Y6DO2oUQUV2PWB427NJKDBDAwXyg1nS
ArQ0M4KVxgO9N9trHT8U1k3wifRGiM1TmB5cqCxe9HW5wV4PfqwFIUTniUWyQrBc
13R/HJRIE0mt2hkhhzAMa1WUWzfY9mVjmvx991sYHGhjPzRrdYYXp9u7ja8bHPyQ
fnubby9uPBM6T558lfW21AlRbLj5eSqiXaMD1QP6j8dhaZhEs2SLyc6glvlscqzn
uYfG/a3P+WmA46rtWPuJk3X1fI+PTEI/DTS/9v/Qt+H/fdOz5NmsEj714JyZFgml
1SVthztrL1PCGEadkzu0su7XNgL/kVLXSZU1SMXZSpevDWg4yHkiGhWj4hj0ZdNd
wSYkK7jNlMh2EWrO25pqP5YkgcgaTvsO31284X4VbOW6+2HFwZwT13NkT0e0qPIt
p637PHJjxaNNRKLG5Lf4yphQCVa0Ryk9hhzwm6qGRFFTWgyDy1uVns6ig6SXr/9F
Z9Nw+L8FKVeT+qnL5ms1UqMeWGkAQEfm/Iwuvvx9GOPDgUYNJOFrJfYkc0CikgeV
uqg4TAluHk3p1GM1a1AuAxzUXDHSuAgLG7AQZi8MPy2M/Z9rMholRZx4/F0+pMrM
7ulpPEkWd23K0NfuO+oy3AW5Kw5+JkipZqUvKwGQJcyodRErOqnAm6kYIwG07fJq
oqdqmgnNprfm3XzJ79SmXqMmhrxZXq2HMiLwk4/eb3AzIWIdGfSmZnXJrauk9+9F
/Vkfc37cb02UfhMu44oSsEEQIMm9nSYPT6DJknM9LzR5CHPPE87bSkgBz4FYPx0r
Y+J9KTtMFubMaCfNUwlZbgJzSS7zlhLD3lnAiSotFr9d9eD5Ai9USDknzAo4pAb9
+cJazoEJaU7kFLaNcxGwwCFxEAs0Lcd8i44fLRQFLtnUryKIKgPmop6dzCN9Z51I
2s3li13O/S2Tg3FTHvJ3Hu7cS6YAhGSEyhNR3i9Fa52FafmwHc7W6vNb4LuRrReM
PV8TTv7jnAQQ44nmazOq1oh8dNVHVAWjDfgv7lzrIThbRonYW1JctucYmclCMu7z
gY6RvHRzT+rbJFd6+a7TRMlg94ILEgj7Uy03aTpNp1VQ1uhYKV4Uwv811THYoq/l
9WdSwFuQGj9IM8ago9cgwY8szK+oEEfdAP+/d6yRkdewaJkRtSfy/q3mjthjFVNX
8DJU4akHUEo5m9/HVgXdat+sme5toAp3uVF7BI3OZ1u3AT1H6b7BVILFWb3R6noN
QhujKpQL2x4NiuDO8+pljiaHOcpKJhLA/znw+edVEuN5wKoZdQK1Q4brFhr5IZmU
FwMJIjJ2c16ujoNP6tMnIMWJ7T/CYyur91mfpR182Np7ItzDRHB7DSoJU2iucf2n
jW+L2oORCIzJyx0TKF+z+I+Sx/vqQ4FDFj4578+Om7cQtKJd00TILXUJkp0OZBYf
4T97PHDwufZ+2ADSOXdstTcFiPtb1ln9bnbllFVqUJP2PoQeizKJYSPRFM9qKWR7
BSqOuaolOV3idKfMa5yTm7nFfFTZHtokoHTKIrctIS7e/loW9LkB/qCficzVIBOx
4fHMQvFa+R6tDu0JcjiRB+IQTJ2f4CAl999wyjc80eKPCi8M+EcwYNDymxpZ626M
iTjXF+bOTdIPy5iFBI6LboDieO0OXbQ5ng6Up1A3NLPyCfZME/YxZ25Gs/8yTGfo
Fnn5540sBIg+CC5OfkZaKzUJS2yZwscH2GRX5r+9A96M8HFVTmKwSch3YrLiH9sX
h1i+NY+sU+mYwPZV9ox5j6w5Gqt6b6s3NIhXfFgz4FDqZCpb1Y6Y5hZDNxYA+co5
+yIUTgr3Zn35d3PywlekiJVvNnfyJRiIrZrvrVa2VdmWiIYXFzzWajiqzsTvK27v
tQYo5gO4RrWJXHGUpeCiHINjDertPv3ImdodcekmPKc8kd0Gx5G31YAJY8G2TDHZ
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Nn2LPg5xYOw7mWC1SD2qFanii+cCIXqazHspnjsuEgFULZ1aPxN2xi0n6Hu+7LVN
s+SRJQ1Zdh6Xtv0Yh68vI4Hwo0A0wKfXZoOYU9b2EtSjtdb+9TnIlXg1zP1idzrY
hktUPo5JX2q4kediXr3MRMamKwY8QH0idgVHlXu3PBmWjddfvyGf8aAUNtc1V882
1GiHqYzr4M3SN795MBi0oFk13E3oEAj/F4Wbj/v+PXOMqcTrEgUyRdzangDjc38k
+SnAqwY8HuawoWLVOmKNqWV089/0gMSPtpH3F0W0wwwLUfSi4oqF+FjP4tyHUuwf
jq2OsfY9iEtNjeqThP+1iw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5664 )
`pragma protect data_block
o5KWN15TLe2WrJc4HxRjtkrTvox4rwmsIfjstCQRHg05B9/nTLIPvkOM0xStC2GY
WVXnI1v2gf9/k3CrAIjtHYTt/jhQpYvknio0AaDNJCesbPFJJSPIiGMfwQOtaoAj
wxOZYEi72K+X13C/uEMCXDTVPXp3VP/L105XR8mKTbGlLWGFRlPntus+uiK3Y0GH
NtDyRftwuzyYm4lZ/MFBzgMTjY36K/vzVyjqwS/p/7vksnbO9jE0nYUSRYYODWr7
LyQq0VTVdt5QwYbyAhhmaEuj/dJX43LveY06o7SfeLOwcHtqTjdZ39OiIVk6ze7n
aFyl2tVJoa3Fp/l+yyCezoSC8+Y5aYzIFC/xoxJqUhulfejSzvJ++ZtFlg1LRYwq
56D3NS6dMITiLsmksZPZdh/AfvbY37Z1FBfXwjQ/NnrGqGJxbx4KdCNTGY9urpB1
NVuzr1ZEEtD619Cgf5rGAhxj9UdqQW1bJeulj6FpvcYQ8HGl6aIjcfrFbGix/9ay
6YJZEBBH8b601TsdInGQby13iCedmmvbmWOBg1jpAv95QFUdUMcjlA+MwvoA8ZE9
rkxsRnL7PVlH+TKx29WWapsWIzD+ZIzYmMhgmRXOxmpA3GRf/F7irhale+6AM+Ds
aOJ4y1N5FQlLZG1A4knZzjVtYD7MlTRry/nkkObC4ubH/jWQ/6+BQAGaf+jgt4IW
3oFHEuRnszav2NvPMLx10VsYtuyk28ALJwyAZitvBV7Yv2OjCq0pVUBIwMtfNvs1
nAZf9bvCiFxc09j+ZcmkHs7itZgbmnJYxRBW4QLbeIev4fZ2yitXmPwdhB1tCd/E
Wg/FuLQ01dp+Wqs1hR6jqdNCINuFiW5Y7qmWJpX38rqeO3y9qIhr0+sclLXGaeIp
iRCyJRW87rsW2tZ7hutwb7tp03cpUZSa+Wcz4RIdQ9bpVWk5I602mj1QR3pHBgNF
moXVv6Nk4LSgnwnEPVTHDYTp6s4XRfKMZkd4ITzZ+kBmxuBvIlJIFbxYHzRar7Xe
9sPJgGlWJy1w8IJH1av1lxVJzaqRDIoCH9KDl6PKHEqF5ec/8+MLxH3eO8kl7/B4
Criu4I4yH2Pv6R6zHkOzFol0lL5WAtxtzPxZypXP3hYS+nfWXg2qaXaMXwWNNrvr
lwBy9k/7q1KHXfmgVB2BQv39quMVbeLoJ/mzjGcebNItIvG29WYopoRamX6uhhv6
xnl/HpbRXN0tEFFIjjMusqA8JFhdt3axjzpkNXcGar6oynHvkIfqNfHI1l2iO9Ym
eWAJe7wOCGMsdEDQYSWq5yQ8XzFunyrBn+o+WkKnxuCykqBKoXB4bMEGpFilHflE
zMDUxxfKZ8pHHbvgrC4tlgUagM2wqq2O3TmexocaDfDmM+bMZCIT0sLcCitSmFhZ
iPq7q/wvgsNF3dVD7b+sOjA7WvIeVucQkqJB4NphdStNXx/wPGQ5J0AIJVeNgPiw
HZTc7C6N1vyEwZAmiZ5mZGwPWWVQksoGxMKIG/iTpxqxEYHkvrqZeutmT5q/B5zg
GQsaDaN2qN1Q2OhZTLZJmckXaOGKeRltg2XS84dJ3Y5SmTo+30dyigoHAXwIoESo
KIT0sPdVschBl+SfAdKstztJhnspfRCpWZ6QrNGgKeOUP3sCuZV9Yi1qkOspub9v
2rLvnO0gqTfikgEkmouqoDP3HbKTVRn4O7ny1KZ66j1Rh2JYo2/jC+73VOs9uzD3
09mChIrk7fTjh/x+9ARkyGHjeOV4FSkftrh3H62sDcTxCN00TjhkPtzS0/V4PbX7
/IwQ+uzWUlPBa9lJ1TC/nKNtLT804b+wIcydMChoRkQd4IRQm5Ejz2WU6J1Zj0YH
p9hgFm8PWyLoCEKG82Ztr+0gVT55xrcLEdL7uUONZuWbemDH2nUneKVQjRSMX2un
GhXrS+VURPYKvqT8Y0Pp0NOJfeS6sFn+39FDPHFmOmFaxc72qoQARgTi4qke0DkP
wpNtx97N6yeN1Cn7Hk+BsnP3j8C5qwAVXlpTlhhgjqAFk8AlRUXlcSJHIZQX3mZe
22nu+O/cWEftIuXAUXQUPeGyqzrE01FEg4n9fLRu6huJwYZJzdOtaVS93vAfRaaW
wg/8H3cTbpiYmL9s9gIz+imNQMAteqrGsYmqfj6ApbP5LSTHcoQH0jA1IRevSHYr
JjWXnuo1abhmZF9bGFz9wPfqQj5x3Qy4PyzQrpvx+o2XK5Ngygu/rHJ5Cqqu57Ks
CZgkJ+9S1KTknAj33LjZK2xvBYZ0U2FGRWiGgucWb6Wx9DlHKL436xk0WCUhoYEi
4fRV0dvIcv8fIVLuI7WonUzTTYzuOuBmrBuHBHmITbUN03QGQjB+c50SG9Fir4wS
fkj6H6UDSUp+V8Ihd6qOlQXwIx0gH7jHZCjR2fIAoFqfzcMph9/1fVflqs3irk+a
M+drxTFRIMlREPPXZzHnpcBSz3/X4W9hwBBg+cl8kck2moco1rIbnoDpJkPVuI6X
sZC1DrXaEeQvbQwOvN3w09encxcSuzCqh60frV9pvcJFaJPn3ytjOQlQm1o9pni8
CZWIfHePR0vlHrfKRt/JzIBmY6avPl8EUAdr/pojHc1RToj6hpjxG/9/OtDL4VYt
tYoncjokrKgfDII/D3XkTPLaug7MaNltdO8v2FQUXa8dgrqv9YkJitfv71LSFBeS
bBcKA6R4F3fSiKIIkpi+kRB+abtxqgQ9i3FrHqT4lgtlFJscJJVTikuD9FFRHITC
aTyKs2eoaHKCi/LWWMlydbt34WCxCbDGDzryqleyiAX/7QnsL3J/rbFnat4EB4AB
IinRMPn/OLLaYffQL0hXOH8ZqyqfK3+TqTHnYmrpOauRUatwXOFJyHuga0ahacEh
saAMxFZvWneh0VIPkWdQEbtHprQYlD8tnKBMm7JnHo0boJhq9xvSQ9hiXUdYNumr
ULYkHj8I57g9ShYqANyK2Jc2VnIYAelBXfGEizaaFa9BFSwbqe+UkEg9KzlfkS0Y
FDQlcNOIV5vuRrD0QTzddrs360V2omPyQgr5yhvOHGnulMpBF9GMjd/wfdCFyIBU
ccOd/0wXGr3adCgSRsizRvuOPpYVKrNre7v5O/IqKPUEW35vd1PxkQ37Cx0MW0jP
b/lHMM3LATIZOh4rhjGnZ+Hrm/v3yPEedr6KC60mw7Sv/fVFh81m+OtGmKpk3zEp
LNaolDebp8Qd1T14GF7kMNPfLG7nHWv7TBNw0qmb1QZzBEKEvdpfwHeqyoqnJABO
GSDRq/+qPXvP+GL/oEaBojZVsKOKZnhdc+4O15krczyOBaVoxkcXfCbu49zUeipP
cQDdwTQtQIS4ZtFWWr+gwJOhPVPUDnW/Dc4vPB1zeTrfphacujTH7CqJCXxQVnvb
n5ZUX6tRwE4vyBuxCBWqY69zUWWFGUVaVLyNo/SHsxJ/fy4dQuxIq3gLUtKMDRUy
vC9xV7EsRms5N0b5RHW87l5ywUqXxdHtKVxMFrlEYJToCPhO+vfRhBNZizJDTqIR
prm0KUlWoC75LMoZm5GBx45rW8aYqTn8ylPg4YuQWWBSPLlO4aSNFL+DlnJbGgoh
pBb0yTD489Vv390dGPFGrfK+2xr2o9whS96vLQYPYgyJ1yNlm+wpby1T1rSlDh5w
+AFP+Peqtyo+hgfpgHqxa6uf3mScV6uCinPypz509AmRuCbHsmgXy2pzFzbzq2+n
1t7SidlIuh6qoh30W3wrmJaws5vSz60RFcCHyAKhI+nXTvKIr+THlB7GLk4tmRJ7
3O7TUcPxA3vJe/SQ2uNeWcERW5g597yJL1cMbXGTo45jtQDkREby5TFI0THX9ch7
2aB0jmOzOvMac/k2QXQdAaZRQ2VJbUVsZ7dt8IVnuJ6rpLKdtlRH06f/n61ilGxP
GshLHyAmGwQ26W7Kl2P8lZzqVdXI1UQxUaEspVHeU6UDvaK9S1Lkt9zfjZkRzclj
gsN0FkaoIOuGZzH3yJyIAjvBMFr6EW65IVlZxZaDrk7dQ3zNSjGe+KPlLddCKIQd
Ww7a5LnkmM8i+/pSTWXpLS6rJtQ7bnUowDq4njmw9pIxHfJYV0OPgOnLOc+X2lYf
nxEhcGGL/2z4KHqppPpE+s/pDKiz6/zt6qvLkp4q7ihEDq7tYErm+oL9nPu1LfLs
ritoSj5Xm4mRX857T59yHXMnQdy/h36THIBA5BSczgw8zj5YdwPr8G7SNkhWlcSa
2GIxcL5QkwBvDQ5TV++qqvONpM8VtDWwC4CVJArxZNM4Oy2KsCmxsm/WRxMTK5bQ
WRDeO6KwvuGEIciQfIKihx14WhfxML64/KzI7HQEPSAFdFVNPTcDTZV4j+4yeeOS
EhUtGbj0bldlIvvRRlbLWJhHhf/KvKG9oZH87g5ZXn+hrSmN7BkRveicm5H++2QL
nLdTHBIBWLlc7mcx2Gfw6k0NbEs8iWJJxUF674Wbji9wUUOjBx07fBVhkm1ZmYe7
kTr/w/fHI9oIlH1M3xaY0xtC2E6rQWOTNhFav20bSwr+Dl2j2Ukn+/gk1W448rMP
XQzut7qWI7bNM5Niq5xTc0rx77yIjpmdOpLHdmtbDzWSNmnCZHw1jyMdsyaiPSzT
y8p7k1pY/12NryEOytkCOaDSOXt/MCetA1yA0MO8rrHGhdyLW5b0OXRCayP87Fdh
9sCxx3SMYDunshdCq/hXTsf9LfcUTTVIQscvGjlJhqIu6RgpgHW2H2eLPA4fRkGa
1WlUZM5yb9nBzmzqyetmCxZgfZ8fXmo8XR1D6wgc2Y0HeEqmq340BUd4Hi5z8TJm
SV8tZleZQvrJvj0GKo7wiH3el2y/peMA3G+kZU3VL1Qx2XRCdIbcqPcBDEyRydEL
9/Tx8TYolq6GMPG5UzJIu/g4uA1kqZhZtOJuccwXUQMvusP0y1Kw/iv0FNAWTVqp
gxw0yIxflKuOrnLMZw7iyOCca8YYLwcFg/D0GIqJOGTD/NnyN/hFYIP1cbRojKqE
m//HqXwGCBlmXeBpWKEaSUj8Sj74mr8W5gYYQNe7zIqcIT9faoWaoD6yvcm4fskF
/LalIfVRKdjcGzLH4p9kegr8I8Ce362jQGIXvD4UtTc5WINWZ2jrtALYPbj4VR8z
91q0eiJ5maFOnA+FvOraWbqib6MhgRT83aA6cF9FNbuM/Tm2KwZ9NT5VJJ4BVKU4
XOb872YVBpCaykdf5b1g1AfKU0SMLvHKr2sITSgFDvAqXHW0/Bg7OV1zqWYp7V9b
MtU9j97AMbxc005HsU/eTV1IVIL4w9ssT9iIw1ITqoZo3h8lFWIrGDr4hJcofXMG
MsK3nBYGfRYXsM+iUOvDp8h0csHiDMrIC239teUghDQCJwBQZCgBMtavJZZpB0Vr
KbzHan0lQFHa6HrnfmpkxxCffXMeun8R3VdqfpZEgjCXny3GrQSTYVXCa/Z4llwc
4gGRmzV7lroP04O1SNXDOrioACEn2nSeqI6jKC3HTystCYOy1+L9O6PeewCiPvja
dZFRZW5W37idf9ZO+XE+T4dkToET/0L4MV5GRH4112I8KUCZPCf0fgwdXuyzDVvJ
9K13+o3700VkJqzvnqh/ZV39sSGQxoO9exKRu6oFYxipNSShV9A3kqL8Sm4p8Qb3
ZuOJGNlvnV8O+3ja6pPgMCdvU4jJ9fqTjQhgmO5G6NC2vU+CzfkSpP3qm954VTCI
qj8r6SbYwg6JGEhjObw1CljPzpaYzZsiWROJFJYbTy9Xp6E/bc4YWisMoGZB1jHb
tTK2dCq+LzZwkp6fiyhscg4RFJ+063FZSrXx1wfzTEOV6mlRT5e0REHXpsHkZaIg
T/x7N461gxf4ck6DibJY+V5FAwUIya+/w/fvlLIsW0ThVQKPGeoXzR/iVFCgsp3O
Zk5/CIThWBYGBf6aIOZ3MYMvtPYFeX80+ueoCEiV07h9zdiZpTGDh0Oqsvr8CBiG
ogJLvlH7lSlp2Yg/FWu0EBo3WKDtXcN0NEX6t7k6iwhrOv8o0sDBK1KYh2ooS21B
sIH3lRaiE7rU0AX/ipuerl31E0ImTNJ+IXAJGK8S4DC/97ZcXqvYocFa0znrp7wp
1O/bosM3hOwzOrwfnO+RV+/h5dF77A83dukPwqS0BjY5HzeLOw+BJoGjznkXrIsa
CSzVtRfB7I6O7lBHuxL2qKUBTxZK5uu3LLoC7HOQhcuF2dWoa6YX9CFdjZrV42jr
mA6qpyStygZCVGL2p6zMrL8J0OJtzAk4YKKU1yS06Ca010wnQ7kA0bQ60PDud2ay
uVWZ+OmPISpiBtYmY9qZBoxEqCR0sbbE9AhpatGtqEGKUX8vQAfJilE6NY3nRqF4
cfloyS7xIusEGpJE+D7DKSX34pVxEjL8hgWespL9e/23yZBxTQvCJSpghMqc7G+G
COTqiNlg3Hge21DwNZyT974ixj2IPqw5VqfE/P2Gt4v978UJFcdQ4XAiVfyZPksD
dhh91ueDGJEkeX53/HECq8rCjghk9CO1ilXTfE+zFkUhhU+K18/8ir1G0vWGO6W1
kIzPWC3Jd3bqRXBHkdFrKjPszju0LiUAKyPQLR9meqTYYCvDzeTe0q0jqB9B5YSx
+3K1ZgBUFkQ1Dn4aVTbZjoi+Kp9fI9xwzuJ8C0JtrHNV0duwZXACOp3J+cxwGPBg
ATXMMtVeIAH5FqRl7yyOUdSh+HYkBzg7DDF6c+zS3fz/b7fM2MEZyWJmy1O8CS0/
8Vd+FJE8kUWZtDVKOGF3qVJY9MClN4Hw3Clgb2Qze/kppGtW8isHe7RYTcXdopt2
oQ0LrQB6RFc8v20928DAlmzM/xOJk1dBsSXa91qTR300ohpyavJLeHRJp7EMnkeZ
2EFd1xklmu5SP3g/Wf5RovOpVXgfIcHA6GfpJoa2ZBC4eM1GDD4dwZpmQapRG5Ba
g5WXGtS7q93Z8zJ9V52s3ytPiom8OBbyNYCI7IQUr4TAzm0b2UAPZIruJFqk3IQg
fdibPui4EUe9qS2BxRxKsMI7pgV6GpmNDIPsWkooKfQoJXmQbnsQE5pGRe1XbqdU
I0V8vK44qe6g8aIIYkPhs7yO5eE3JwuOcT5sxWSY2zv2c23jAMwoLr7D/Pt3+wj/
nvhcJe2xHyASjeYKoHm0pwN2IaKJ48c+GqOlSj0h3Aj+RuvQTOrpVL5LUDHg8K+R
FgFRZlGip4O6Hv8zC74lFKIOwV6bk15TQgpWir0AcgEIJIxwZFuz3mgm0y1otvnD
44iclUR/EPxDKXdPyw+hduARTZg3h5Vy0D6xu9oYaEO/lT2xBvgbWngHd54WbdNx
pOcTW5Xs3hXbo/3seKCXCtf4fwHhiUo0L7U0xkOMQ24xSFFwIbgC9PCLh7U3fRU3
PJudr7sh7lehEoKus1jRQeWQfZvSz6DAHhcvP+kh8LCO0kvHVPZhbFqJfxgvTRoG
0CooQ3dGMHOq195FOVzqMEroo4Te7oeeQDKSpKEnE4kEx+QigQQACO/K84jXdgna
Pw0LYYkhlTBR7Bdsq00oHvWajQQOQu+Qr8L+mBw/7u1DxjOk8fYxVDwEJnZAG1wk
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
f/Arw2Hor1HeYNVJNj5zUW/I64UnRb2mSBG/V5RyEUCuO+4FP5OyAz+dklP4ODon
yxYEZeVivtV23svApSwNqBNjanUJQo8MaUVp2g4ycH4ZgSyQ3re+H4aJa5iiryRu
rGDRT5tkwmVMKTzgaxfaXfK4yKS0cAWlkZNbYj5GhvOxi+pfVz4xBQamshWRIZOE
iLS10fNQtIwi1xKGtuFy7vRxFqVKOOSVT3XUjKMIk1auPFooHOR612fylKc73t0Z
cdnE6JJzBbSXQyS1ISsQMis0fonnmh+ay51Ggi5cOU+fyczdpQToQRRQW27Mg+YT
Du85tZ6WiS972ufqDC5kRg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4720 )
`pragma protect data_block
1KUjYZ1TD7DaAC6b7ajrIu77MLODRzJt8oUogqUgtlxbV1ODIdIRXwDnJKh2bETh
FfiU/5L9mCK3t6S9W2WmhBzRWV4i23+l8QK5GxgRL/JOK3vYNC4XMXcDfmxZRUhD
zYJGzUL/gjGgS77eYgw0faY14NtUUetqSRFXjdKX86RLSbUdDWmTtZ0pXSq6iB8d
ufCKsEq4LYtcVD5kzH1yrwfUl1TK/05BYKNmMdARQoROCUK0VySr4LZXtLv4ynS/
HpR11iGZufDUasd7Gf96d/f7XhFa48v/NEFAD8V+yTy802jBLdlDGZGTC8Ho9pHP
9gFkkDiGq04VqSko9CvDb19NkTMyzX/BmIPp+meCVUOpTt+9M0QCkxNsHlGHDs5O
hJpKgGG7l9/2YnePI36aXl7EqMTrKaimkKzJHGQRXab2RCGFRZNr31kO/3ZhIgrh
mbI86PC8FsLOHAA5LwBZnvK9F71ttWL5U8GtGUew7d9L5y3AUuteU4Bc1tJDxLyZ
VDwVWRxstlOGMqvxg6GYwRTYIUXVa9eq6qGbNEd/LBsf9y1j1706PZcN01/EQ6bB
0eneHQNbuvZ+FaOsq9TiY6zXFT5/n9BLDC3RyHsZfRCwBmgi2QwpkEKAgdBI2kcl
kOWF4m5zvxSvyXT5PFr/fzqzAA+Yld1bdZJuEggo1VxvrBONYeryLdl1+VpJ0AtI
i9mMpFfQCcC1Q9KE1f9PlOorCo278VXJ+o54aTGa6zigodbizLFSPMiVznNbJsls
tzrbPI4w1tmV2ynCbyJDlqfpW2TsrEzNy+0v88bfAaEL1IBcQWastkc6514Mch63
IN0h/MJgiEhxaGB+fv/HTALTdfDPPCk1MvetIndtx522pAj9EWQ7bKL0JBhbsQtb
Jv80U5Lok4DIeqEDHynhmm+wvI3xssVoK8JVd7hVQanN9hCf8uaL6EE20wvhpUxv
X8YeYMMYpgS+HZLemp/lcPtk4n/rhVNzNC+/OW3lrVnA15mQkDxt+nTy6+OWQzu+
XNL/NUAGl5nd7V9RKK2ytJcYPAjcoUpB38ky93ytkE9Gr7XXO9w5D+FijYKpM8Ck
r++gktrlf9VQGnl1NrU+xX1NzB/8hj8OVGcBkR+YgTMeQBNXvKNXCW3ACej6/rd+
CTVmhcv76ROs+1y9eT0WBs83dqavNmmo0zP4/pG6NhmR1yMpe8QXj37W39Qpi60C
u5moUx/aRqH5HAL5cM7LfqrLABkCmjAJh0szQMTYTOVBaDTghXAgYLnM4gdXbxPp
aBYkIljUWVZt7jJecausIBB8Cktn4ObkR0MNQxILq9m6qtYxK/M9yTUJ1lPjDO8O
BxmHnx6+lyP4r4WatFtXNLRx7ZjWEDI72AFnGv6V9OAuzW0Cbs3e0PSYC3U1A4CX
h3+sXfqs1dK97z4cw0Y0ugIkDWT7HUqGZgukTNzmNT9aukeOlNMTUb/Z0xVuS4jA
+0EyD/l9WDMYADT/9L0HrYz5ZgINTMPqYpWHmMLYZvg8gWVO9O93hskzuPAW8/Xp
2zm0cOseqCLA76z3VmBaVpg4DvzGLGZkBM7TnztQcKiuIyJ/wHj7rPYBg9ka2FsY
BaZqXbrEhufFlt4MkyUU/nBl5/3qj4kMVuQuWYnVBflmkNXL/ugpROXEMl0hiFmr
duB5MXFNaQgKMeNl73nTrTpccyzBeL29zdYei8mwbBdmlcdqIKbDQQzg8dubmPX9
9SqaJ9T9FEv8bgUTGgyxkRIHVvK2po6o+Tif9Ez0bGC9s/jNTL/LNM2NQcjlcOVu
BCajeA2CP+CsM3cMgAJQTH6vsTUGAgmx8+qMgiF/HCFBYPMwRswW4dyveylSSEDI
WHippmiSWnS/SRDqnPF5GxWAmhQ6WPAoJT6KF/V6kL+BUYgFH84d5zJ0nRYi7QKw
K3O3U68eAMJI+2nBQvsHmL16VRADeDwiKFNEAt2hzzB8cVQJCZTVjmjtbOIkvjK1
AJL/dxuOljFfgbDlFUkgZTBPrmFgfM0OHNC9363MgXRz7qjVXZZuuYkzK8yQa298
2ed2dCGPEoW9bDabXMK0DQT4i2i/RCdI3i55TKOCWpJtb5GO/G6V9TAPNTK+BgLz
Yi2hYzDCuve4FpsgAeGfZtJN6x+9yNhJNe/MC+ROYZzcNz3riRTCgOVSyxPit7Mq
IE504dScyhFO3AG1Q3grgp2+1pWrpRQQeSgY3VYMpJ2i5WR/ZrfMILEj6h1XRxBc
4dm8cjF6WTWMOs4BjqbYQboHxCTOkHn17NBOrgA1PykJ7LZy3v9wTDsj1RzNy3EE
P7D7analuItwDSvxV64cQsiHjlgd/87xngoi+JSeKyHa8ZFKIYQ3pKji7074jQa6
n8Zf2osfYmLCIJmox+vRkCv/wdWIHkruCFCS0+LQV9nq5OF9GfF7gpLN7ihsyrll
+GlsHCdCqQEky6fHupJ2c0YVpGVeDeBLhKWUGVnqLED6F3Dg/cABabREWMPOuQcM
5OEqdt4FbexiMqbTA+XZDmbug5ci05AWxDE6Xcq7rnCRQnKlW6cNssoc9QAyOd8I
2QH0rJSh7Tk2PYF3pCpyk52el9caN56mN9VBIOoWMBrCybhmglKP+qa7cEhvUxbV
yv8Sn2B2Pdp7WcZiIB7cQ2G/gq/zJm2uu79fUPmbRnBNhq/vLBrIiB3XkSSPMUje
jC3Kl/xDhEWOELArvYzzkgFWkVAl54xkf2URVcCR5awhcCp+pSX5Y7jRGBCWOoTS
MLBXtagPvoPFQ4r7boiVWpPVZW5jkYY8PexsBCHKWp8KUpfQEFGDb9carsQ4wYin
1KyHR8qBJzd70sPBtdY8zGC35YzqqX11iPGv4PdKmd9eTziK45igRV5mrtAPrVJT
ZOIAc8K0anSU8edml4AeuUgAXbrDatujfOPzMg+Wcx2RnmUm6Vfl8zCpFVIWHsKq
vH2/6HPeqJ+3xzHIBkif5ngPOCjXFGyBVlx3EbwY7TzIl7KlkgNUtV2+kiju7VEX
JPKNqN+ajDUo/9OkSWHWulpDc7GcbCPhsUeiNh7acIU+N1l6yOfztOyjK3PW7b98
fcmXsEmvBSnH7+oXJ6QNHBTROoiSq3Ai/EC/4PyjpUKecNg0Azh83rqMhSAQARQp
Oz4OiLp3cyxwTLA3dt4gg25ghc9yLwbdnZN5GPXv7svanWd+biO4qGChfAIydZK7
9z3+i/x9c/3+YT1wah+dPDZTF+YrjN6E55ULMbUkjAAkj524DRTr1oSL3KfBmkzO
69yXqoLRP2dG7jlh7bLCSo8A4K6IDe0+SIGkSMqaT2lM7hqgkkdaqILYxBweSc7N
JZ8+SyKaIekUsgZoIjAiSassaz7WH3pR5HooAU25DYroAM5eyA7haM6/7ghvwIRk
rTxY7VsX4PkFr89xfSlTxpn+s+flgG7rrifi/cV9OZ8vaXx0nbyuLLuwnXG/9qWl
vLywvVZlvfNCQQBsEZ/fmV0sUwxB/DFrOvTYpfmcAt8FKV+3CwGn/wBDjlWpjlej
QEJaG+pLk985oLIL2y4z029WJzitULxLqDxgddZy6adKKqno0Iq+vhnxmkUzlaWH
34vuFud4yurnIllNb8+Ljl40qPxx6gurINcF7974fJqp+4E79SNo9t3NAhM3c+9J
cGCqg8TiX0w8+/V0x7R+KREeoOkWjtd0RUp2AbAbCG5yxEGoty1O/+PnvwC1t/58
rbsjDBvXvvUkq8htqIH0rX1GM29f+2Cr18tyePd7vdHFH3jahv910N7OV4HGKCPI
8Vhiq2irJSCCu090DjkYApQZs/DSzZvaXG+2t9Y6tKcKh3POWvGlKAVuYn3eJm/y
wPkhZ5eqLmIJNW3wAlIPeW3trM3/KMHZpHpm8pwlaazEMEd/a3NJVsMUKH2dUidb
qNrfMocGp2lAFo7jZgJ/5WYTstGto7OdEcmOFrG/BAwXjw3KkJNNLN/rKlmWveic
6GS+nrz6L16+FiZhkb4/44w4sGqfT8Y/6C/XnrZWfW157xVpNl/ZGjqhJlJPnWYb
wErL9QpqGE1OEFkEHeSNdzyGC2jHnxUleAvkjsfjcDb1bTYBnrAvLN+J2SCBkgxV
VApuVA/3jspjc4DzCyXzZqs7+erZ7XXoifj1eY/z3uiqbQ81QgeWeU8KO54eNoEN
S1Xry9bCsgMr5gfyB8gIEtvBHMyHCdwYqfzMhbrIJzhi5Sl4Z/puESA63r3ChpwI
OVIVCwf9/mMf47KkcULB7k3X3pVOBlkb/aDumJnCbwQ/vh1V8Y0FWSMKUnFhZmhB
ZD7FllVGTaMzd1bbgfsLGKGGB+/3RRPvwwKPwoo9P+m5BNog6Psx1m/V8lK2PyWA
EKi7BV/Pfijs78KcvMfo2SfgSf5eM//EyOmN0g18TzEMqP2bxTjm1TR8wH6DQr+M
nhpcs84/P+wAcwXXMQelfBdYLs0WBAwtkCvlp+lK14Hr8/dSK/i5EQ1ZXNroWm1z
QM+BkVbxEtqRJaj4me/snittKNzpsuWOqqS7mNYXJSBd6oCMEOXFneocxOHJ0fSX
M5z0j29Ob3KZQczsR3Vj7nC1onkyxY3RHv4+w6y45U9McHoZtXKwQ4JZkErA15JH
1GuTb00/1chLy1kYKpc2ByQhgGUaYNV0Nq0PfLUV/0wd2XM4IQq2YvdLmZB4AzEE
4N3IKH243Glc0Re5C50UAXmnuqn41RlhS+dXJXm4UO8Zy7ph9G/J6OQAodjT59Ai
viEySNCE4fez1DxSDHLi5/rul2y0jyffjGfdYFa5o1qIrdlFJK64x9sgrBayI8HM
i/quhkftYOy13JTMVLkyF4MbCyRiv9u66YtBnqDTuV+nRDBlJ5ykgAALIa282QBN
G4r5l9kVwsLWxbbFeIyFuzeFxf8owjvmTW0mvssSKPoFGWN7reMhVCQAuLabDB84
aEUFseF/KFWozezjNZMyGP/MVPJ0bZ3+CkNtIWDqFZ2eSQ0GNzmR6qt/zPmy8UmY
8Ugii+0euNidjPAdFgAzD3s1VgMShk+s0LaXqmAJcL8Z1tDf7R8E3LkwzkpiBoBd
CZsm5OeMkVSouslmvICIfcMc7Nb1icvmJB+/FGfbO6vf5OWlCqnRJo5eSaS7CNAS
zhmDDC5iVXY0uBDyNBHyAbx98/sEaKM0h0oeUW1ocIMo43w9XNqXBYY+sG5d3Y6O
1UwWJ4tZ44x4Z4rBI1OKvZRL3RVV2q254o/RcmvSVTASAYw2oOuXnYj/rMX+TqsV
DOWmzvRUfEKZUVXGYlSl7JDYr0Bj4S3qi+7YewumL92bfyho6bVyWlGNJaOd2u7h
Lv8VukOCHz1awZdP737RlwVBO6TTzh0gjEBPJrxhk8edTmnpu5jycQ6VWnilgViN
med+w7fNwbkTx0j5yb9852dsC6FPklBlvcHleobZP387/lp8oR3Qf2J6z79fA8kD
JLMaWCnlrlSviPhXVapQ1QYsy6HvUkME+9xJlin8CPFp46R0drvBdW6q87ksNJtk
FLUkpdJxii1asd7oSUZSKaaPV9Awuim9Xy3UtV9guS/Xihp/4CA5XdnVxcgcGS5U
9+Z97AwWCXRoD73P0ZMjFIv862tCvyzIwi+gzZA2Hdz6WA17AGLjXrZBHo7tWXYn
ycc8wAhNWNMZMZvEMmfAZ2eJCMYFzd6wzFXZV5trDHNfi/oQXZuBJHB0jfbq6/ud
eUl87j53ZRE8cA79fbKLKvD4CmlfLwFblIv8/9/E9at29CTkzYLVYKodZqHOKm/6
FG2+/SiL3Kj74Zo+97fKcsOOtPay6rTIRz7UK8XhwLg/SjwyB7FNcK9ll7Hkj5+M
rglDSPMlosQ1ekh/9LSH9dpVGJGhbqZqcwIY8+NWaZUTtmX7mcg+b325DXkogNtD
WeIfIOmaI67srZCeNYCMLSMaeHrEYOOqzsz/S/S0qoxIbVWKECh/Y+JhkduxIOP5
yVWyN4v8lAgw2xmBbn89cqsvkxsh783IvZamqM3tWUUBJWoTw0GoMlxVyKCb3j0T
ccvThdkA6URqakGnf2nUeaqgEevzCATZrTEiyWmdZn2mwhaL9+KOJufY8umtXdHS
MIeiQuyAHpgML6uxu8ksHbZtSKN4XOJCcf2A1JvbzXoY/0XwWD/fb1/Vd/0/H0/9
fegJ3O64vz9/eihpxh1LQE4dvwELkR/KCvgPiETpjG9EJa4B5N6kQ8awjDg0jiz4
sp5+VInxcWqBkV9NuSyAWeR88bYGQ+E3Tm923dx3/Z9otQbCZEEJcIUymFG4AGTK
q1ZRI++ki7TwYY/AXeACwg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WJp5SQfe7+vOhL7eAAh7bCLYOueEbZmRsYZiNl95iSvC+MkiDemk3CwI6BUBej+5
ofw5UJOMqAID6OsAu46QdZOCZlZyKYk9+KGc7EVTtG4rXbDctyIuBkvdzLMramih
MXTKpXnqVEOQvybXWw+td21P8LEDvXgnQ5mCLJFJzpicQz8F8oB8oYLD084IfYXd
zNp69znYqlMkKUV2DzAA05Z7urKbOWoBpBj8CuDNOgz0s8ErNctm1iH8BWbCxyXF
LMNQlSC3zfWZUwetJ16t7cVRt7bJzehRnqRtQ8rohz3R320WIvbdkYWY5q00VMSM
WVwF//b8Q/MENxkyKVvTOA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4288 )
`pragma protect data_block
YMIVKpm2vsWNhV0Xh7xHSQLKxovIpifDaZI8oxuC32Hbxx5PA6BdJxZJf5M3tJJ2
lp1ilPPsVwDjK1UdLcJkAKWnmhKhZyDAKQcchCm8m8oUIBiiQ40KkqiQM1qDT7Ge
Fa9ssD34iugmJP/ygEjdFMiUNxzxb5Kl7JjhTcaT4Z/9GIYWUtDL2rYFDFdxFBA3
v/3a11uhlLLtsxdrZdit4C8tgZeqdLaId8EznKCofvnbaFzeAeCWbMXdrPGBcQrN
APuyb47MGtlKpuOAyZXokpUzp8Obxo4tM2bzZq1m59PsHlv9YdcZ2eVTqePNH5fI
XI4jgz0GjfZeanOVTFStkI46+cygSyzOo00CSkvrp/8OhfemLEofyMU4+OGLcoUr
bNMn6HyBpFMUoVydatF4t2yOTcyHPAf59b+r+m4hNkEHHE7W08chu7uHpTnbX6Rm
JPBFnNSZLCtZfBrDTubmPfQuXslC/mS51sxsTmYhMBV63be6L9zSIgRK6PTkBMSC
FWBJyOZH5G1GjEtbHzgcW+Vq3O9UWoU0UhArvoHQorQUYAYJ+ZbesOLOYrkEgjzi
Cbb+R0HNI7yJ1paTQcZ5gmcPvRSTlhSxpfazpsrBPMztt9Augj4rWFRjmu0GJHD7
8uA3JFrYXtnDk6TWc+J1pWfJkeS39cTYCIBALRAXIzQjjkOlh2ly64cniVil2Qbm
rawN94Rz+NgsT69nUhsrGtpRSG9//I7K7+RTIYIJLe0FAKtNvWxjU+L6ADSYw+Wn
hJq5UxR+fq63HNWVWpzO22pgrMKzOJVlR4vQvwcSxbT5JOk3PnTyGx064jJSxCF7
PLgPdD+njFcKuf2e7Z86d5cC56SvrdR18qXUhQNgbAPlAolNCoXoEHkT5cr1nsXz
vpjhXyxfrxvnhAAa0r1m2okQqpR92A645izbK7iLadEyRKGprDotTEk7qsnSOU46
8xWQ4ZqnjvWbx/Cbp9LDKaWEHMwisji79aWAOaA/XdaZYavefZP+qoY7n5fbEPAR
GXSYJ4rf43z6ydAMDGWjAIpy5ci5rP6pxVLlO+49IAEIzaaJo4HXOUK+fDdOwcgj
UAR4a+ufKmCmJ+4iZkyKDJjX8OF5mv+kTd9zvyud92s0eW5pXKSyWLDTRmL/ho1p
10C/jW2VdVSjXDtxow3XSFgVJYBB4muCZfnOx14qTHKpLq6iCDhCSxWV4JRuMEh1
xbRHKU1h2Ceh+j4siuxJPFM9H1MP4gcazC6WJd90MOq6QGAwaKpcCBGbmpCZKuRw
n3cg4YVjIQc+Uv5HmEbzBM2RBQWLxGtJ9Qz+MrBUfq0lNxmC9H1Abnaiwi6K/csZ
15Jfmo+TbJY3TvI5AeWqmbuODRTFpnHEHU7dm17YejNGfbwA4xP3NMVvvcB0TnHj
UdG1MQvx8GZMN4Mu8zAds5wqIrcVyznJryGUmD62s+2TLa1YDbGRA54XOF9NFHc3
G6jJ52rigLmIZezsoO/W+n9jWf8xym2lHuzPKTgmAXSORLMoHYh92yf0c+sgpf+g
ovbvyxrLUM9cbJ6zP9ioTD2DwIPuhCBbst/iLjyQWZta4AJS2RqURzhfuxTZJHRW
tuVZ1fM1qwBf0CPTcHW/Z3FpzrPmdkvq1gEkk9btnQa7bctMbuz3v+nTPp/8xkrb
tqx0Vg0pmPJFREI2u5b20bnh64tw5SfAozgZAIEOhSoghLKHohZuK0NMbmqkN1q7
lFy4pfksrhZfhHVBggZap8UYVKPjYmMntAmKrrSzPvxsoSkGhF9dtH0MtdrXYuap
RaAT/x6D3W/5jcrpXgIOfi6lCmA0EWU7vEfjEEd3dP5RUDpG/V1plYLFchxq6KIT
jrbysgBp54JM+sIzzsKUO3bEhSIEGAoWxln7bPJps3XA7kyflSyjmzJYvVE0t7mI
CQaCb3aY9/wIpmOildKCUnhnSnlP4vKrztWqXpL+xy/IP7HLcOMX5QeYobv8YO1J
4TOCnT0YtTosRLOPRZKHjep8ealIJs+Iu9OfdKQFJtPVMshd1N45neb9jOu8L7FS
RnYYcsYmEqIZt44mXFt1KLhH43Xm/Oi0NTB8a7Z/iklMSGvDO+I+LlcZBHRYNYVN
WHd4sL8yWWVZYv08AZnDiPUsLSpZbW747ZpBpbGCLAOfeUmiPPOkgh0G0JOmAq4x
esPwHM0fv/Qko2a3+SGyWDQSTXEzFsB6BP2sbMUG745972hXxUugzpDxjsA5tPBz
6kVgS6UMJzd7BiLicYN8TkTwWrLHL8gWkH9ynYWsc7aM+fSxIzAnUSW8Yt91Mjq7
LI2gWuIXOjgAgHQnFTglxZTHfUmW7K3lm5kvdNugAR2ImpxPdRAW4NPaa8Ah+NLq
qsumc+v6WM3YWDz2nI9nWe3Dz1NoU95M4nGACEUEqkfFoWbYKUOfcZwq82xScFOr
M1thvRAYD94Y1fLJqPW5YaB53EzGiiX5IkDKEhtJaSqmMqllFkh62a7QCFsAJLJR
BQds93unnMpNc6zrEk1OpGZX29usP/48GrqpQEyV7bg2q0I3mqX0DhIe34fwdM0i
VFV8VCZFyy1CHdRqgzunwF7a9CwBlO8WMUWh6+cFUvQRqZk/vp6D9mNl6ASOvbDt
rfslT5r3yagdj2FrIzCCWErXUpG1Y9YU1gAKK1xUgfGLMXns+0amEt41BqtD/8TH
P6s8H/7JR0C5UBQoiDQLrvBGexMFdSNhWcar/kmaQ3BhAA/Ml8fGQMyck5WMTTzg
NG78GKGz8uHCdqGNlq/V7w2Ehdts76kiier0uDafUJ1O3ny0wzOuUuCMvMNFqyCP
+sCfPUksaKCLWWPpdDPciLg5kiw6PkPU+bt8D5vEJFw/JRE4HqVbvDmKYSOeadwb
Z/M+HlFbdKgjo/HW4tRRN0CAQogVpFMuI+I1XbLhD46H6Qt9CB8vcL2NurRMBZUU
tYBRqe1Lbj494cr7D58uHrHHYm/5+ighPVo9p7gQu3i8yRLyOVS/J1PEfQ/HeuqX
BnNyN3D3XUErOoE75ywGn7lAYZcBfxSpmU4/3gKa0tghPmat+4JPtZxoGR2XgPgV
ZnbHcK3LeSAZf+sHhS5S7EggeKbSnR0LA/cQqqdn+k87iBh4usoJA0WJC1XFqOnz
xHyhvaITQ0LDOj5fLUBPXHA5E+00GU+B2/0K5GdzBQjL9MgS1viut78gf2u7chyN
ASuY6cgkTLqoGeV8pC/XKgYOAbOq8e9nMZFCTPFiKnOGPNrA+ewQSBlDcBrN0OZb
xq1RC7+EDCKRixSy2mrl6SbwzO8YQ/UGrfiw7ifd2RAqNRS/ITUsbS/QiD4iR9xJ
HHrCSGcTOedw0imdS+kQuKXcsUid+la2PL2UEOp9aXabNRIVfC7s7P8xRd8RKdSD
ZVpgtIi041r71MM4dZgCBrrPI2R5Xd2VS+ALuKBfxkVvUA+qo3J6AncbX7zvc9WU
XvTeIvI+Uwzb76PPRUfvGfxTgLqxxH6/PLPQoW02SjY2rix7ffUSCPcimJLAMP9w
0FLhk6VHjpGgXvkrwBXPdSJIfVzkhiJNHWBvtQqaE0i98jTDkLQFaL5frJEMQdoH
WnjPP9NZct5mRZZvfpaPL5ibFkZUbMM/IikTjetevYYSeNZsDikcPO7RXZge+M6h
09MtpHXUaNWgN4EXr+r88E8s7vnXL5uCtjR2s8eBPDT3Z+VBfY51Ynp/eGC7JP4p
gVjLoiVMJY7EzAjiU5PjBVrhkvbOwt54N08rG7Ozs2GkCFWsSUI5HedOOOknwc4o
qaqOxx0UVB7KhdZIPXK/HxqUFxKwMh5funumPxlj5b8Ov/o3zIavQMRqd7xeNmiM
F2JxuBDzcnqKf7FpCMYGtj0ujTovzdBhHp0CjWgQexa372bX8P0AshTVsG6p/9k7
h44MR1wUOibQ0tYCE4EWtN/C7w7oXhqktE5z5ByRPWOIJWmh2EMWacqWu9nVnwWz
Vg5YgR6Y4oqDM+uzODiqrnLlv2d+KUjQHs6XlVr6gzgGtJSMdK7Lf26qlE5V79q8
WxOXcYuaTuhCZrQUZXSD5Z8bIYciQ+yuSQTNoAToUXxjh2bg7f/DFRUG2eaehj1N
RS9jabSCSBmdLx1FDScP0o73+0RnkZ6M4j7Yc8lOI5V4yV3DFLczBy2w2Ze6N0Vs
PCf+tGGZwDlxGzDuNnVgAS9inTfGalQ8JXu3+R0QPVEvnkdXnXxoaaykx8JgZObA
bL7PBUJPKaHnjYvJkySV8XWbTIdW0DNlb0p+nL0C45HlAt5jNVgQaCUUal4DQCgj
A5Alsr4EqfBaKII4MIgA1wvTWmd8ngDVS+iQVxjUjjTz9O7fsmU18j/ZDlbjXijm
NxybTfzZG6cEHoRadfkQIsfzM8Pokl1AnT/j50aOj1oSZVLDfq8k1qyAqdSspAAr
qjbO4C7UpxoOadqce2NvkegM/fXViTXKvE/J5QujnTkbcQRBzXKDWIcJagzaxWiB
1yU15wvpmu4pvH2C3kHCRb2Sc4L1d3wr5D9G7mgm5FkEJ45gDQ2wY5P1/68+2slO
W44A9zIT9Bq3TQV+yegYuHP12DLM3Meo6u0nHhH1X8Jt9BQVteZRHkR9FcZ1frPw
bmuYNSwbT7O/U27XxfIguRYQXjRxS/5BiIiOtH5g/jceqEPA9kjz2Ikw9MpXmOsK
kJNfaC8mooYvnXBzAvO+aSrzpddj42MMzxRrBZ8sG9kh94O8Q77Ql5smny9e7In7
o42snvInEkgyli6YQeB5ZenuX1PBQ9H01vRc5v9D07n+FHvYJyG0+cmhFjIjEkIO
zUtIr8vGCP6shbq4wxEqPDLl3OL7vcoeBm/gqQlhu6gR67FD9N1iflOnOGFOm8RN
mHWdLwaPtf5CMbkJ91T/L1/V0XF4NLuaIWXXqfZu5yDWOsxQfs90fWNwzlxo7SjY
5sbOd6etg9H6rhAi0LfGLMKzG3ApEoo3+Mu7zCWQYYGSbLg1PLD2nLoXotHOUQW2
FZJtqOPuVaLZFzuHESBp5HHogplIlvBdfDTU78+vmrtiJXiOoH4rPV3M9qrE/V3P
Dg+IUvb3Z2g2dk41eZLoyWmiuzJvHLUVRsch7KeixvDgjPZzwPgoxZSUTs0bR2jW
oiB6QANTebyNnQQ+/BDj/w1Z6zYXJkP6AtrP/cSJ0P9pHoRD24pW//TXNCIA4gL/
+06eQ4F5tvjJewECe0i6nxEr8IYhbv9azap3bQeTFw+aHwCckYXACswyv8reL/DR
XLh7ybT+rLGXETgmALj6DTLNi4Vbf9pKKsnlwDmf9Rvib+30SW2BClS819nawUCz
BDWpeGTIaQyb2ocgRFqUdDICHC4MY7DtkhFcXBr1eLZO2RwSBSglFpf4McM1zRfo
PJT58GP2XFPzJDVdUtEn7TU3kdWva960kdf9flucMhmPaKffJLH4oadssgUYQLyx
GvnO4w4rXC0egnZJM6SgWe2toq5reflhgkMcEtGMnka2Z1kv661/GXP1ffIfQwi5
BmQiSGxYoWLm7BbDQyl3B7zugE2CPiv4YbX2kMsc9objh8uhx+2n66furXxBNhBP
phbqOH0Di2qztm6mYLB+5m7MjuMq1h0XwFa7B4LXf+4C34FRQnx05coMKMcbZ970
OaJcvz3FnpPONoinjbHHTqNIjn1vBOhMRrBJmLPqIPpi0kAzxewe+Q16GDXysofp
Nra3U2QixsuE3QGsXI3UjQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
MaZofawTk9++MWMLnPzqMS+oF2gt3qouGhPthVn2z2YqBT0sW41KYSlSUGikbQ4H
mtCNZZVOdafSEprS2USXkcn8z0jSoI8ANoQ/hdMgrZ1IbHfy3ZCv4dCssv1VVEk/
Wn9pIACY6jCFtxvoxZbD6T+ahT6ty2UO7GTHWLXfOdhBmfwktH1cydm6pqqsaqXb
syaWxbGHKZQk+tEGAhVYxVMuhrCtPh+TH0Uw35nE7ILT7cyoOnLRjylkx4dlUBP8
sM2YI6fTPisrS7ncW35+b3BBf4LRKloDn5fyq3/SJ6iCOHb+qDZKYTGHjWSh9Qrv
a0MwyRgbYYzAZZ7q5leAAQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
TCVRyHJfRAEf+QwHaj7KGbXXX1DCYu4tREJxh7u1A7/hNojOiqfC6cXm3Pv7rIYD
3v/RgqY95CX5CQPYyLi6WM86yYmw7aaIz1eUqVOa65JeehiEXwf8qN8+tiY2eMwt
9OxmExect4ixDPViNKd1UKmq/hJa/wC9Zzg496ar7qEeXiv1/ylex1kZ1W7sU2Lx
hk8qZBe4bj+PPc4EZSRhCuVC/tbO2eP3eCnpogEVcjCHkGtglZl10elgXSwrt35U
EQvkvQ75T7z1TVjgHj8EF/jFBH+OGPIoh9zeFEEbI5Lrras6MiZAqWUUl8yEbxfL
5/yqKRWGCAtPCp8+FZbz6YXr3dNcsynj01p+C1K5w5c3pmET0zdn1a5BxvaFNBf6
HUKEsB0QW97QkyrlLLW2iXEJVxh+5CZWwBoG/A2O6+BFMFFLUmdJb4Uvjiafrzdx
zM+9e/x2wVmnE4IkRm7PwpMQzWYSNca4Zu2FT5TyBZhONcfvFMV97dugkWcoVaOU
zvmcLJwGtt3PhW1QTHQ7qbuaB/Btolfrk9CIryxdLEsg20Ny8L+KP2QykjLZEKls
pjlLWHU0THerCmJzM1XFtQzbv5xJ2bofYHqTJl43tNgZczj+LX593vn6ol5Esgiy
v3qLIF3lnWywCeTgTvtG078GxRQu/ANfKXZfrHACsAm3wbjGSPY1LM/pgIdRGxax
SMnXCXRMrZpDLyuh1FPJBa1lUexGUJ9riGO8mQPWr/2KYkR4sn3qVtnxtKMLL3p1
I7m+VQlHB6pMNc0gcgqE0nX2uIwv7nOM9O+raCo4HzUp5iLPv1joyiRvuNsLcbEV
yucnJ8ZKo+mF9P1FSy8LGR0xlzEFkEwbU+vfaQbKEBgIU5rBN4/A6jil+WX94nSm
VaGqbrCBun1XybcIAW6H36aJXDxV56EkySqPtTbjkmVB5KPX/NUdRlqiwCd7r7WD
Xkfiwd5pMSWIPp7NX3d7dphS0Ro5FYu9La2qhHWf8CYrJ09aV5F5oQmtsmNsIHXE
6U7QrrIMr8jJ9o52Tm4ENcnQn0RxvkeYMVtlJ3rc/JaQFKITCEdxTgxmQWmKFqeO
n9lHIOAj5nrrVVXotftyLm584oUl61xQLVhrvDLlu//2S34j+vf13TSobNLGyK8W
RazZ4rmZ18laGmQBeEEq63bzgGg2hzDh3aSUDZ207i/ADa04+/GPbEhFDbfpzn4s
wdYJlbwPWQdKlMlNf7tzbzV+4abWbbyiGPzAVSztcKcMznFb4sPAPXbN/Zg9OZ3n
2DPHeVF3ApNpu90IcK4G04nx6V1WkEINL0NhU6r4sBpgBqOaCWWTJJWGKyvkoIpk
jCxgSM+wh4gvDdpa1es75+8Pnm41OGmFXK7fLqRkFHJ8WbQjNUtiWbDorD/u5F3E
NGA/pjxOkOT0nC8CCdMKYc4Se7HmLVSyNjyj9r40+qEB+aoqWg/LGgTuEqUwNTKW
7RBu8a0yUdiaeM6D77TqgUO86+//8rgUnA1Ho1LN9T1w8a9sLZZfcy0brjLGF70T
Z5zrCSxFbMsUVFB1NZEZHNrsu74mGS0INGfl22FpLVejr03+ZBMr1SGzDPzDOBmh
7Kdx0/FTVPv/Wklv8/wUWoPhu2kc8+s+WsVT3VW9IKlLyZFRTecxFYceeyBIEBVJ
FXzFDa/VgxnjVB18XTvhcDc7pvrfqJWNNwCm4Si1hThYJit3DJUl4iEhX2vZW9P1
8wbPG3nRrYk2mULSlFPR+gD0ida9ysQvWbOpYr6+dOC/uhFUXD6jxLYJ40Tzzxm9
Y2fC38rPo2kzb5H49P/N11x9DZHsSBrVYJKGKuUVfD+RerYlcsdw3P2SdFi29hd9
ct7AZZ0L++YGfl9IuHyXZ8lhd2p0cp7ZgvZjVr2sOQeR1wi+6RGDjG63ny8G1txK
i1dX1JEUC2aQE0w4XSN+iHsbagVUb0xTQDNFopeC/z3CPjHL8ikym+3SrwTeQ5Nt
nyF/LVi8ryROyYly3DU7AtCOibXWMF/VkeoaWfsxuyRbeRlxvrR59/uoYcxxrKzW
BhXZGdsHVmbLRbdzbg8MpqEH7Gp6vzjVCDu24PzMBNPQVUDqC0v90R+ycTZZ778N
5ZfDC/bR9yLGeBPGW90c53AWKx9OV9kvbea/wkZpYU84wdpRtdwBYsmIZfAS6F9c
6Yojb/509NQJh+y+nGnjaszhQCcUsH/eCPkcy0JKjS3/x8r5Oa4g4065/5PaB657
uMHLcVNwYkikcgbIbjGQC6XfGUdkDqQzg/+8W7G7OkQyqDWV08Depa9beWkB8Ab9
LBZi8ga6TzIVQr77+OduKlhbBAwARetkaW5unHy90a51oP+tBh+JaFi+cZGlvRwo
MCtBwDn0zCZ+8hkTKpoFhuBJT9X0KU3qRTmpF00KoDDgdMXGUBMvExwTz4TUuEa1
UhzmUOzFFLMpQhAqwXyD9VTfF44hWT63Mi6GTlRs3uiqSk30P2jhahYd2WA81B6i
DfU9IEX460MdutT2UON094+PyP5w0VRWL6lhjQ/ZSh/PzF5Cal/3IXNA15cmJt9i
wabWxjG2rZvm5yNcWhNnIJdyBPerl0q63gCJVJP5OIV4m+rFVBpCxoMBu9xKIR0L
Pkq40H/dO0wjHheCHaE9tc68q81n+j6MEBzJ6DbCsieaysZ12PpHTB4ungKguw6g
qWZ+Ufbkj8VoD+ycxCtUjqs/7d+Hd727EuJVus5/hYsPdRX6qcz/w2KKm3t8cKXx
ZoVqMlEWpiBT43uYywscJpTEvkym5Y0ftiw++3lNg1sxYG6wmeUUKUTJsm/WARJa
l49Tsvli0HwGSrxYF3BUGvP4C5+Eoyy74EM1GJIXAtfdQxTJbT8GdDuItUQ6DhXV
V2U5rAWVxY1HVMC/GXiDQpTiWsc8xQZKH1jo0QxWSQssJmKFD8on1M+DdB5TzJ7I
xf3LYZxDnVjPJXKwAe8p2lAEhMGPnRXyLFP9NMASEStSdJKPOGClcnnO7KUz96MW
d2+GinuZyapfgnAEQJ4cEAAUcxGm6FR7mEVxdXkwdoxoq/iRPGl41g7cQjk3lN6h
y0qVO3c8HjbHWD9CBgV32FzTWUpmAu5FOoMMDgrWhfjJFXEzlgmrTZyV2qdwxoxl
uD645KQp/HFPkDNOKn3JieJkFvhjt5kpcmKVwtGzMieAKxwreKbh9AolTgZ8L+0v
N4/98ELZn3di8lAYaNrLWh2uc5Tu5ReI7wwGGiiZssIGr8jDaBVT8OscvK/4gorj
0vRx+bGjwrr0m2Z4OLtr0Yb6iwsvGMEvVS58s4y+WSVkTU1iHkMl7vadP44GOpU7
iN5QKrlRlwFKVqQ/OIJuhadGZtMKDnIKOwJkt5ClHejIkLK3DIEDCFVt8g3qN4cx
RYxJh7d/m8LFp2kviG+tBsrX06QMN/CiKsmh9GpxIUA6QAagYtXV6gmiXn0/XQA5
tPQzoe9CN/4wuXjIxxs6EfdsC3BxwkeAACrrNPBEjhzBu4d3TZQLtPGnVett+sa5
lk+KTU6REoNLP8JMUA3IDqFXBcpJgZqD6BUFyEBQmLxNndx5ye2QOXvXbyCZfHGJ
yCLwU+Znloir9DXc1yyJlFUcg/hZUYCwLnpPivYklqyAbASQAH0zIn4ZwuVTrRz0
HLQ8l+iq42M4CY3INT9PPbHzoN1UZC9QBjrqjcbuJqd61kFzA3nuZ7/gSn2kmCbg
LpfncT1c4j8qnaMGFnAzteayV4Kg+b+mau1CAMqDv+Zrt6DmR8sAn2+0sxBW4yi3
AXGm4oiY65bFrAQMyswSkUxl12tYMT985EtRyItzpZYSQlx/YOgRyVVOmQ+8yuIr
59K0Cez5K4qRzzrM2xZ0sv7obcXIixl8xkcbL13a/eh0gMhnqcomm+9xEMcYgfRk
moZwabasen5kzhwIreWaw/Z/sCnmIQYZ++MdPNM+s7eHNVS5Gn5Uf7/2qI3fGaW1
tDAqQnvM/Vglxr/ACQILONnHPKyNkRx7QJGpVh3gsWtc7RfxY3yuZdYTSQ9Hq2kl
KTIl8D02ZJSR8Zo5/ykyG/n/ncOPu2/KLl6AmkRAA/Rv7AZDL99s+98IE060DIz7
UDv4V7fg/P+PG2XZxof8ug+zeT+p4ZTgrAkPa7HuKfUMdymrP2NdpMvMu+tPzA8J
OKCZPDXyiAobzDcfd9GJ5fzelUFfE+vjAjtcB8AspN1Pa1+wH8BrAWA3T8A8KVPq
CvLlfIHkHRJDCR35Bui1qAza7RPXOHJmttCR4FCba6OfVhsgrnBHBTplwydR5i/a
7hdR/OT4ibCWhSytdTYLHutj0Q01QkVccBi1Nnks0Xevy6qDRRbagzmY6fQ+JP+R
Q3hDiWvJqM8iNTGfBDszUGzDFaz/Tvy5NQP6Wlwu32IvjTbW47WyOGgGfOxg2qjW
FcjZ7PHSDIFKFef878rqifMWO2YQCUVH8CypaJtHspozLJpEMPhqTVyAD2HOhmvH
SQpQwPQc/LqmOkJxZUifpUWwgNdv0k3JMt9XqWTO2uI8iLXZODV8CMQqQrlbI4AD
3ywBl/wKbuG7z0ZKxWgFiGLPcEyE0KCSqSHaKpy5Uy9OL+MwmDwkyGHgt1o6JPyH
I15oQKNEtbIrd7mcr4vCjI4xbXjTvHMUoV++0mKrBL3yWGDCRG/KSrs9Gb7L/wLt
jUAVWfv0bZAWagh/18+XDFiVNQDdQZ3RvdOx7InYGIBwfTjYDmQeASQylzm560ro
BqvHKdtClUmqEkjVF2DUe0f2Fslh4YCLBlAkFWmUr5Fdx06FKroUnQCLgYiDjCP0
8I78gpDFNH0CJ+HFXBGhLdJFWE98e2FBDwVU51YrB/mx6jjY649jJn8URrkPs4fE
Wg8J01m2hIdoIpt85tEmaPPWgcBOoVVbe9kAKJ7c07LtcEGjoqFpr7zlw3SmJ/b1
/DSUww9DaOdJAKRGChN6DQcnUkiIVCVLy40s6nUfscLuntGhQW2yVl9P19mm67ZO
HrJUwixKexJLFGudcH/oI8E9siadvSaksUIKtAcLFhnRtUO4VutGtGbfd7cHI4U4
RdfomSlihF8bR4zQNbbn1oxxY/F0L99zNZB2NOzkqajTn4Bb9zE1kvA9zf3bKbql
GGn/7gz4MGPaVrW+G/r1Vcy4atuu35DPyV1clhwQXYY=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
J8mB6bBEmEZ9ho85W4fpp08n/zUgjr+RQt9aAHcbM+GiKI4ntZkx0Lxpb4ZFeHB9
uosWr5y2rmpuq+s3378ZRQdar7H0zepQ0f8zSQKN8k0wBL8j6r2AECYMvB+dI628
+XmQ6/fzOs0sNMrocqh+SyycjPkf0uOxBwN4yJ8tuP+Eego0gs1tX+V3ABBlzQTr
JxUSp13C+coUB88P/MNj0kcWC6oqiqiTyZGoVOIf2U59KIJ0eXjmN3NSJIoik7I6
P3wjs1sd57psVtWUKLxSoW1ahb6kyX22xZwnGhP2pnuiGpM0U2ZE0eK2cQnyoCoF
t7T0ikN1pGv7rtJXCXOc0A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6880 )
`pragma protect data_block
5QZlETDo9zqxuklSG/ZNOvyFWYu7EERjmdRihcq5yKG5EumlTtG0pKT5IuxG88uw
oAruikyNehEp5vbzdOiuCPrcSiOOSz//hHX7MRaD0ndR1tjoFdGol1K2vK1hlY9M
QYYGD0EWpnD58h36Be0kd09hGYYcM73ZZ2/4S7b6ar7M+43lSSeXPpnRbp/aB7MP
CMA/9YUa9KB/VnbeQqbX+mE9Mh0Z9l53q7bRhJdsfI5QZdFWalLcJ6UrRXF9eRjB
9/ws981Xc/S7I8PhNlwEa/22MmZhEGS+yX1ejFTPe3ns3cMvcFsvWpk448A/N0/L
wLBYGrDsniAFHB7uzfcoC9g42juPRd5haE/Ed7zaBRLKqhLKK9JUD7kdvxFYFgzL
P0gC2njdE+osfCkCZuoVpKx/oTA4ozL/s2/VMofERZqyxb+xGBQlHjJz5THlCn4t
k02dYsdsRFMzoeRbv4uug0phNT/LJZYSnAfNkw1dx16WmxvRmKaKnKyj7dVRs003
vce3N3HCBcQHPSYuDulJHtfjxoZ/tDg+C443LEMWKNAySNNmWfJ4kqgSM9YWXUHS
/t0v5Lmp/EpUJeyRbcWUUpTbvPEprYzFFvzwLA9Axu/6ncn2JAp7Hw3CAVjCW3R5
pC/YfeTN6vZ7iYkxla8RhZttkHrRBHnWtjADuU3lHyFCbwHslktuDFG1vjjL4Ehp
8sFTw399Q5SdU5KDE137HKQEVPgPRKLSJ0YaSh0iiodUYDPcU+o3By91qDCnZkNw
yK+Om2UtY31YuVs0H5HLLb3sTQsvAdByMb43FF285tYw1hlR9KiL0XdFXgnfV7/b
L3EIgrKbZSL8qQI4GrxMmCrKBsj6gUW5Em2+Gu4tBRb9kK6bNMGr2FGMMcXwAtbd
xP+82tgPqAb5WW5Og5DUH5rhyLxDz6IP4Qz7zJY3LNiVpsmGU5gfIca4Vw5CRCLo
9xO5lk8TxFLjuIf2KUBhO8CgJZmoyq4wXHF9fmsdh9+hbSUE+7ApsBGa0GBYIguI
fwWYT0SR2fGd6S71jBSQa5WQyGGESoYL6OPbcu5ueif4gTn14F95ERa87n02Op8P
CnZo89AaHKFqvGUmPFfFE8QKK+l0r3O0HDHWkfxFZ/x6/+ryReGHA8bJJei2bF85
qgM0nwRrOJyU9LVrJ9LtbxAbk4wrc0QA9gOfYoS7kZ+c42Kw3GPvO82pMQQ0EHC2
vE4DMvJBeWkYSpusCFSkN+u/Mzn6XWqeo9WifTWblnFP89C8G8PeNODmE0bnbpaR
ija/M0cVHI6ewSUMtILj9ip9Ux1dycFyB1arPsyfsGRIZVxBggy+AODff5/W00cm
a196wPPdVO0pVxIC1k4QB3IghAfD7Qw7GkXoZQWBstT+VZyse8admQPw/IqWxJvI
+X2aNYdEOCv/4D1UJB1x9uaVMFT5H6fD5gJOS/JsfzAPZF2ejxQw32k3pfSQbkke
odo4sep4eSNy1LvFPtgC9h77S1uoN0sO4hp/9o3aekB20vWdjDxu4SIZ/ATVQbez
CVy8vL6LY1/1HJGStojMgSwgFMneqmGhWOWfgDRE6lo1W4p6cSJTsKMz7as5Wgun
si9cBCmPbx/fV4NK2upzt/rtzcJbRMK37cbhLAXWDxyKnw5wr7Gi5tRr8O4G98nI
WoNY70DW6f2kdWrojirTQqXQe4usRISAdThL/5mbIpixFd1COBOVTlRph8MXVvEt
OpYA08vL6MJ8q1EjB4PKwWv3Nts8JT1tI3qCdR4i89+ELFKizeh6aOuPX0j9Vl+J
ZEU6NVscrQdGB944GMA3CztKkimqRHFQbSjRqJhr5bc6RaH/nQ+Wd7IT5sbddk8g
zjCwtCwzbi6iI4dZesADqo6R1DDuRlBE/Uvj8HYxrwtgvtTAfD22AWvOFT3qjdlL
9QwdwxEjtGMVRPrGGhxiP7IGBGNff2kZ2bZFxGPzPf4KSyDc/JPZ/LP74ZQDhVeR
MnP1itA5kcXCPkGiBYs+2t53HaCdsU/zGELr+HKnsVeRN+RDtzPJ2nF6zyaUqWW2
oeltUK8XIiBjQZ5XPh5ACOw59rafpOU+fSNUuLbyDgpxBRHw4/fz/5sIRwcPyify
86jeA0kty75IyR/mjd8mgKiN4V3ouKYhCpFKPYnLRA1zXyyYHUH65uR3tc7Qzi8v
7YiUs7qMttdXCrh3TrBVCC4VMnbLtcC4YJRRju/EnwTPnoo19QQ+4vl/CLRg5huZ
oWMOe7UhJ0ek6bjZHxYTsy8FVOtWJl6+BoYioWMiagq7dhPf85AOkosG9ZfdssSt
wbIyZSX+7eJbVHXPvGa5QSpks6r9cIKtu7h9kqRGtdNYMGyTtTaE2kxarDg3rsrQ
O02kZ1bwBG5XkCWDK5nZjavo3/LFRpSJa4/eOSokLLitJJhve/IqG1bXhTYaKIQJ
gKyKFJSFCSsyvCJOGe5yv0gOuim7HgX5emafAr2J8+O3bxj8Gy+9WjI6n70qeAqj
s9Y+ZDoviZnuq66tVkKo0ddDkv2qgsI80GVAox0lSdgs4epwLjimJIDy/mL4NrPN
q6YhUpkTdl2wlEq7OU7MKAqsGD2BPxyR9o9EMQIT2Pe9m0yWsINnu8qqJcTHIlW8
aIDdEYOS+lZKXWhtvmnR2u7vMdcvap6SpAwcAXedfQyyddoIhzAJwkl5KyDQBi4N
72MzMBQV6nZp4NlusD093+p9HCv/RdNR7T56C6X0h7feNQXuV2lWuau9F44bsESY
bTm5GZ3w04L/tvnmHg4eBIDWXyd/9XWp0TN1q0VNwo1HPWvcgsFLWzwXcEhUX4l9
W+2O1T4pcbu4WSVhYegAJ47d6QbQRT7YQPMYncnsyVsyd2/6Cf0/fKDcK21BOQ2Q
3IUxMIpJBBtxMvdQ5t8lmM0o9hJWJ0PjVXPSh5tXmurS7roZjpeKrcssYLvWAKOS
HJylRJESxAwKDXqRK3nvhnSBzxyJzCmSLaxTMCrQVPOhh7/FVLrChdtizwf6OD3e
v0CNYfluPjTEOMU2t3kYxCgujWnxcPcBmS+fDzBan6QbWLQKyMNeHILsTSELValQ
DzK7tWV1WDZ56mi9cXUqv1Pa81cN+fi4xmVINXrxdQ4E1LMZND3aDxDVtctEIrGF
SSyGt/5kHzy1zf3qgbrTMgOdGjITb4TkueZ0IlkhgNX9hAWuGZsiNG9QXGPAqnBe
tSBercO3N+gAFz/gd4Bt/HdOCUeoWRDLiSKKaRkeENb1bRLwU+rAIDvYtAJv2CXR
4mRUM5L38oKT2sf1rp7GsQ0i2L4k9gFjTaWYdwoCfou1xmC+eGG7rXG5WeLBGjWA
te8HWGf/cWEImQF10uxYPBgIBJdwP67b6hmd+x4Q4+w0UZA6SZRxUW0BlS8IglGc
VkFv8sDtiCtcQFWcbIaEea0L1Ymdktb0f+erFiXo6Om3S3mhneflkQubpVLrplQL
fiCXKzNeXCruj4qzz9LeyfapDgmhCQCphF7FlJfskkp33HaNj73g0psZ4EmQ5KKC
KgRN95EA4hgj7u1DgLuCFOei4NMwXv8vBdvOtvGH19VyTKh4c/iOXGn1ztagnlZk
7Olrke8Mq6f9t7OBvNVjp+IvwsFW0KN1bmvW6CBaDmfwrl7M68LqEYZD08V9hp7w
EdBeLzD8IlSn6kRDM9YGHVv3K+QkF+RVveskM6xUaLj76PsacjjxUPzvlkXvtUFB
j6/p55+O4yuyS8ScTEzhOE4usbX/QZFE1vrbYGHMNOrlkp8VqTPOGTiQzykUjVxt
s6kzJ3dhyyz8C0zSRtiWhQXszhXfPzYAum8Hoxrbm/O0KZMEJJ0sq6GqoC1FB8p/
lGLcGNjpLov5Utk+mpYMbmtBe+TJ3TnUTi78N/Ud5nUAVMb02sGmKMmlUpNoJjs/
NW506WE+gF81sn+4JQmcJIhOcpLIxUJYtEdpIai2+gEHAGFYbmgl/1pvqFxC/7ML
uBLRbhXgWu/ar5UqWbi0UGWCX7gSUJbYNjr06XGZYrKEYVEWofteYrfkybFcTqFg
8v9qGUDYbiMloF99omilp8E+XYAiLGXbMNyR/1ZPHNlmO7XvNahbwS42hYDyCSJl
4sRODtUAMROuyDWrSLGETtdgsAzT1e5sMuUNdocEE06yIEmZyp2yhlBgm++Xh1VR
j2edDziFBfWc2PM8436JQVxcas4X4FVDNXb5goK/qpwc1x7IUFcgHMoFTARuYfxN
kYqoGVcPl1NTdVXsag2dloI/21YqUkpyLbNZysE9sYLc5mV9nFGSKCcCK9dRnQEp
88M/dGqYPCRl8HksC5JjNDhtTCz7iFb4uCr0K3ohQ7vo2dWS+sii14SaWhpQTkBx
KLm4+wJDryBB30UGDECTd59Kqjvn0lBylse56W6CGkLozR4Yx2s5Wfhl4depc/7k
KYzaO7SwXNegaVsgmwofYByVSAO7nteqGPfqa3GFz2LAbzb6wjrKlf43Te12c9hR
bOt3evyGWarPINVvy7wvslm7xjh0wQ+r9FZUGwwB7831PSDfWX2JwqpG+5kyJo1C
XJ9F0YcDnUdjcp1y9plyeH3XPJRCRYEYyvch7SAbk99OyrzxvrW0mWAvETzv08lQ
rE1ef0yx0vfFSZPUk8yNHNLK+eMfSNapp5bzCkap1khmLPy5XCXNjpdIyxmqosjJ
Bx0l34so+oj/XLOR+xc/IeTm3L+P8/M5zahwJREKp9YfhMnKQtUMP/M5gYu8Qlee
nnDJN/uvPNo6TSkFkgKKp20/ZK9rSx8gDlMLzKmACjNWTl+RFwFx2y62/iSpIsVh
4AOlIOIwVck4LPRlgNjwO1YSMUSwOU4BNeu4owvG/RBLyXJSMBpSUnDtRbON9a/M
Xh+Nc8AO4CbVLDD2cBcCj14ddLKuGHmei5JcuTcA/NxAX2MmqJ6BESAMfbMytKAu
pVsA+o7X6uX4kXbwp8hpf0KpEYHOYRVyRdHro1tytZoTcv4u0bn70+clUmqudOdz
AQEXfECJmCXZxY90KiDBkmIkCD90/itJP80CUJuWALtWepIpqaiimulIh1G3RXYX
ZwrZGdeZ4/HOLw0wmEJjldNqUrojGX7XvA0T5Y8Oubhe/blrMcopNg2edRDbXPki
MUn3CDQndLwATUV8/fYfQPDFMIJ7LOxSsJMF2mKjYFENrpMvC67r3eFHZDfOLq/4
V74om3weqypTfXPJ35xZJsB2cJqLQWc2eL4w4qsfiGy310btAgP3PfBSKVtzQtCC
h5+iFHzDVueOWw1Bf4RX8RHwjpwEMRFINrj2zXueDRxBPQxcbC6Gp5adEMDzltNJ
TgP+8e71GzGJnTxMwBsi/MqjQFl3IBTEauQ9tbyFEIFR/rtylrZ1Fh+pLLYFD/Mc
pJ1NC8yiU5jBSV3+lj34wUD9XKfutFfXA4d1q2mGEh545f0Wp3DpGp2YgjfER3D4
QKhgiIdqBPdjEd2pYgxolOCFbwTWu1oLcZTo75wMNDHtXsQXGq7VwkPTFonHg4wA
DZ/DLRn5DoFC/eZuCA25QmGwlD0e51MXhf2DVKaNoSZksZbYOKH3rE8yyJqpa3y4
75wyXfDudloLoz3//QcP7sleyvbYLfQIMcmldg3SezqRXL4OcDqxn3AHfHKFzvXC
B3G9sUxozPOGCMaNHKv/o20CsNedjxZrCnDiHLj2ekUcVt9d90a097WZD3bbMe1V
tJtOqxiNeT2GlgOl6epOqUdD7/QJQWyif9oadlG0PdcQ9qQcZyJvPW9nM5fcS+Ba
ClE9nZ30T/GIWF1TCpOiE2KPbXIhAvMD8oabs09NhUhqSVmn38igF3HiKHZrzci1
fhctYYesZIuTbjg10TO1xqJBaJudfoD+cYAXaJqPRyofgsPEM3sElHwsX4SvOBSd
iVIgjEUaoxiJ3w3NiZAxeXNRcW6gJulW8WAG5wIC9oInivxDcTWrGBiYWAHzC0KD
5Gyx1IxD/FDpkqXRvnXp3ymp6CQ2DKHj6HKWDRKap0zwgdeHgfKgKmHqPM1tHAsO
wZXlUxyMmzN1FRyqpEViL+q07IJlhcH0JbVGP3v+N+HkMFvci92KX5D3QPpOsQ5x
tpii3RX7unOsKtiAYdFgzAgMbuVF0GLmxudgEtq0F65zki3MySrq9jZfDNvEPM9J
MZ6+6HyG4eafiuIZFufjpWUHd/UPef/cs58m198equM0VTqrBkHt+kL7Ca5f4I4j
Z8kPyuwDn786uYRnaAAsyVb8pRudpB1PdHBRkYxeYB8SkpcvAeBbnzJJXP/fdeq5
BdKdww5marwSDz85umtTQSdTpqa6hXRjLrUJdiuG5GFuBQ3wqcn3/r1cfcoQHr7G
My4rEILJA5TTUYZ9ZzdhsoVMXw9GpqO7Sm+JoVgyVffMWzu8hD2dGnDPOQRMfliX
Dn28wFDZOwTkhSPAVRenunsPVGXe+q2ZvgiiW3epxim8d2ITVRuyMRSeM8puXa3t
32XK6JA7ri+4n/Vywvoo6Oi5rf4mSmpYfBa0TjrDSTmLqhLbpBKdWEVy8p1WgNXa
L43WeAkdz1X5U6jEJro/6EJy4nfZo24nhoC7gmbczgFEjmCH9opLSp6n3PLABQa6
9K0B52grY29ci/1xev7YdLdP1Zw8EECU7ltreZbER15vWmc2/Rjs6QtkeHUKHdA5
ELePQe4fIrArnjo+LGXgugZPDW4HUQ4c6yO++0cKKYLuG5PZOvljcQ0jFFZ1dCq4
dzjmLavgAi1uEvPcWZQ7eF7svvNyVR3GSKgAO+y1Jww5jSSTa40s/5QHbOhYfUib
ph+RjMUhcLoMSM3ZH0lpTJiBL8aFfbs7nXpAPGtPSMGHrzTt+o/JZyn3veb018Lw
0jh6pq3/ZTdBOfehoHklix+ipP6ZGh33e8ocU3kvoHeM8FlcBtdBrRqXndE0NH2A
qP1jwbN5rrkL38rJ3h78vTNzfIg1yMXcfrD5ZqvuwCc20yep3oyrD5Wlngfxp1uq
Q6IhmDUScIuDuoO/hTFnV/M4J49a446sIJmhZMaW34421f+y4CRUdzzTZDOGCaMh
szLfqeC+LBuPFT90TIhg0ZP5LGOAt2q65mjW6WeeCpxbzSVB9PB5Cd90hIgFP2at
fDITGTXZhUKsYgiiDZb909ZY6KnmG7XQQ9f7PA/wJZ3su93UnIWsLI804X3qpfh/
bphQY2gFqXxbkQTpIkPskXbLFqzU17SKEN18IAY9FeyFqq73FkxNByZNzqiScc//
hmSoGXZOY8dBuKPVkTc6H+/hOfuJkMFWGvN/1D7zWhNCjmLYxyounu1omL0Kiord
xWobxVLz7j4K63ykjdiUccfzvxpZn4OT8YhxjMU9HssvjgbdCq2wpRYNFEysF5HI
b1GH77HwoSSLBjkyB1C9VTLQoR5dHUDRGtFo+fb9PT6iBOzzX/QD80+OXogbkwW7
sjcIeAW858R8KAxtAMGV2VncFgsTQ/LfHIK9GvSe0BcjPnyYdmOrTWdcxkdmz8Eb
n0Z4KYI3zkXPkj1vVe0bbuEUH/5OisJD15zUekp8cIN1ZQzeC3Lz6V+10I2PyWp8
OEKxTwIxqK/j+hlJ8kvDg/C1lDIyIFwG3Ba76ho/DhT5MBPWXtShigFbeV8JdgOK
YyJowJoQgvk/KGwkV+fgmnVssm7Q52OWZPhA2RYohWG5v0RZwGCQA77NgYEmVD1U
36kU40veGZltVVc2ColHkduxgigt/BJeyYsFnY1hCSq8LmfXdA041l3IpzYqW7Ki
xRTBLTPA9jey+y1V+SFIgquGU65FZWsBWYR2i/NRw11m9r6MhcVc/KkSlNTJvJKS
tv/UaW1w3v3XjjMy15YUNHNBW36j10QybbiD0vW4e5hlpJG9jGcEau6fbbI1v5Zk
GH1CJL561yawgbk91SZKZ9prHKI6blT8vGpKs3xd0HXMHrbGorZukW1mXI5jc7ZK
9iuvgPIab6xbc0wCYAR2MlNDY8WoVyuO2Plwk7OopM8FBjT1vP06rOk7KPJz2CfT
TS8JN979oI0BUOgIA0LJLblscL8d7dJm3xHlp97Jo6rXr5TX9HvVWQxnYnGX1k2m
8wqJ/9CaUOWwHm/Pe4jK5qxP9SAgP+q7qdnECY90+evtk89Gsd/B1vS9Pk4xDvld
2tAbik+Ec/zHoHJTSI7QBdpIt68DAKCYEGkv0/bBPMCAlZE5bs+Y3tPfvE7/YI4+
/28hZipUCTING/3TVh9ueRX+MtMmTd0Pl1RioTJT4uTxDNdNCApSVUylE1FCf/X3
jtAxyQS+T/wGFqLQhElDbX+8N95T5iHTCU45NhD90neo4ZTwQGdcx5FKu1axfGri
h4w8KB2cQmglbFkemyasCpp1ifbPMvg/pTKEuaRIpvec2IJgn8tjEpf+clpfOHvv
ch5EA/NjlHVbVlOo6GU0lurXlqmP5hGD0vUXZQoExVbHfMNg3FViev7bvrGreE5v
2+f1kW4hiNTaFwXbKtTmsSqCdNssmCCdSFYpeOzs2Hl+7EnHm5bZLmuros2zodSD
kurMezfmMbytiP2ETIvw8VsHQsPfcQ+hOPADFcb+lZ9Nt8jAnjJTLtzoS7ZfnHdc
aDAY7u4wBHUuU1TNtbjri0Ec428v9QLBYloNe46cJLySiaX+/7bTBb4PT6JjsZdh
BvllF7z4PYJJoWINMCkRzdS6QETAyjnPOH7jwdhQc5m29ys3sku+Al6P6SyYcHXe
kXFfkuXohmUMpB9wtCGGXM50td3YUiOcGytaGBjz+Q89qO/ywNm7du+IZivrJ/E1
pI+Nkt0LByBYVBpd2A+DoRQXLveYkMCFgsrCZUbONwRW+yBmK+nVxKOWMXsPVL1D
4LnvuJ6W2rxfEaUAhx8RxHPQiUjCpKccSHrIR9lN8QAn9mPLFWQT6vfZOwquBl1i
ZsfEHk8glPQvxrjQ5y2VFTgy8QSVU3EWorFNt564CLewDRcKMg5WSVCJ4ExEiYxY
+g5wRdZ9VXcL4Vx4O1R2tE8wJiBgLCuwgcg21mJj3j4i/q08Fm4+t2UD4kAosGDf
/TE+CA5GRxkC39nh4qiD2YVijTElVSJIhx9pJJaZk8eL6+8zpQlKqllt0JwlDnLW
HYOTaXJtYKnvK4AZnIkRj/xKgaYmmIKPwPrdjAoeFQyjYQ78V7vw7QTFibpRMwHr
LqcRnjWX/4LpEIJFEvgACQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WRb6vIrIeMH0rcgQco8e5Gkf6THu9UFJWNJgZg3aOKOUXdSDRRmJ/+UdAat6JZi/
Wz84F8/+pdacgV4jIl9erDeESK3/Aib7o9AcljG4K5Z/prUpTikiL8i6tTQb1UGM
4ks+xWUvRtbn205qIDjuA1lMsiGmUwCjqk4wfa3J+fkdJk4BBHGzANy5eOW/fkMx
usaFgyGiUku1mamJcebfRUnNVpx+u+FsKIB3P05CN8jmWtiNdP25bUvTxpT88QyC
haLNIeK6yj87Q9BOfPwFLrU2uAszgAegghPdp8eIxOegNc/12KeeNepyjv1IDyWn
b83K8dIbhibhvmEH+OJdUA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4880 )
`pragma protect data_block
3EEpoGJ339mUz7L9jjU/WtH0DZOx6NoigAaWm+GKLBAdqAW26YRovMVAQ7fnTud4
fJpWgXi9NbJaKaEphsVo5boKdVh9ogw/iVPMwt8bt46b1zUQ8eOlbRHAfB+VVPol
mKEwh2xrMzqs+0ncrIVZUqRWvymfc0xEuy1Hda9658f7Bt5eUX6rprGqL8K0TVAK
lYYsQumJ0MmdiUobWfSmC/2tdMgZxK2xMryqojy3r8woAXCarwk/Qy31KgqwXbOH
1tV2CCPbWuJ52Q86/s4kGE03VQFaZeU6xeuvte0JUvK8fe98xjX7SZk3/4aRZ1+Q
4EvM9KTgzphZbYM409yA8fyT94inw8PbltC32t+HVEv642+esORyjyxw7u89QNMi
E9Whri7f8vWF8FQZ2x6GLjZGs03z5XjDYX2hfrKXg9e/g88uq70exJZYz9FRd/68
V0bJp+n7H4vKPUP8dc02H2RQl6A+WXv5QbENIHW/qExytItoRIxQXi+mWAHV7dNS
1YPmNyLwQRE8RZFNB18NQDXg9gPt2OqNyDZRCiR+QdO+BYw5dmsoZdTpw412ib+u
UTfgnJ3Fo7dT2Z4Qeq9QcfS4FDRJUEXH86Z23Jzm/nPvZyC1QvWhGeayEF3Zr6z6
bIGI3m8u0HN+sNliqfCzIhZ9vsi+AbT/nWV12lLaMm2XFkeoSBw5E2GbfRdxBk4R
/OrNwRnhJlESekbwMHuwsz4hbwPZpa4/W/4o+GrHyhePWgVJUdbxjnax4/LMYp95
fzBVDRecdsDyvtRW2h7k1ETw1Jc80KrzTObGJAY485HDQ0FsxNKKK5LlJLDBIwB8
+He0I3qVE6p/Qd6loF/3HOaV/C4U2E5+GkNlSjZ7ox2VXiYuta2G/OZeUI1lIcXz
Zvbd8lEl04RvTJ4tqc/BXNi/osO6xscriEDmickYorjre8GRmyaTmCCNo9mhfEwd
Y1MqMZj/1IleyrRJBj6dM/H5TBIL/2jHrZB+jNR2MUaLFf96FcgxyqPKXgPUXepD
FROiNlWSi20RTmgE342Jbc/LXifOZAbqFCG+8drolWZCSRyS6iYrm9abWC3WIzJ7
CbHpKnt/sas+MyJPzMLafmANHaNTmhrJvtiLJ/7aYwU9n7jD+/jdEHdJNAhJWSKL
OZ0rra8DLOvEYT0j1vPCDJlYhzFnZ29aA4iwT9yb/bYDidHBwc/h8lCv94JBosqb
RgWlfs8sqJ5zaTKTuaW7gqqQ6h38T3CxBBgFa+yNTs+KttdMqT13p1Y2CTCs5UHN
kUteW7XUDx9azbco19u955yezO08trG2wzZMe40blmCHQMTW+PZkbvsaQ6aV872m
Pa+Z5uPdaftVIqMDDoRnFEm/dUh3GutrMymjvyvGoCkUQ9BPSrHFirQWO94r4jtD
wHzKsyXVV4GaS8fIn02Jg+3B8NwSqZcmzZ/ydoEulks+/sXwhhYJsZNrdI/rszg4
841eyRhpba6aWza68kVAqvud26sDGiQ8FcNS3Jr3mQNoDcrs8viSXPYEAHDKrtoh
FIXaLwIocZxMVQBQDlCcCxFI0CvdqhRyCio/tOLJda+74fTgGfpaVB4YRttueD9c
JHV+KcmS9PDDkR3DuSrPShHNyQNA9RlgtNiOStRplDRKveggO87J3NC9cohylU7c
8PK+M34qf8Mn9TZpsu5R4dP3cj+bT3hrQ30HXSujuhq5p01ka0ptyrw2CVMGlhnW
9Nx3YW7v24wfjt3g9ZDJ5k6N1anB4EGOC2wj++lav9bW+VJNxi+Je63KWuT0MjUm
cvZkX+pGEubIS72hWQcoT1V7YQZ/zrukCKnNOcuizGngJmg6vDtIjlROWFd4GXOf
U/Za1FUZVtS4ylxRECgfHW4e82xqpAvhy9Mk/pMKgSEFbgJUDTMWsxplSDwSpcoV
tYKxhHLK85imIHjqIj2ADYV4v84da99sB/UZTTZDMLDE1o/N/1lVH7kq7ihteGfF
dk7FuIObhVzEiysB/04bp3SpFsrE4srSGcgtOenYWyy1rEqkW/Fc9G4ZmZ9u4uJm
VXXtsc1Rb7t9PUGRwPjiQKFBoS4VKUPeiFGfqdBDWs6lWfD7kZhManE6M7h/h2wB
8i8CC47xW5SakRquwCIwSqTpoMsrWS3vrOlh2aDuCYZ82UcYD+EO7rqMT5E+aq3/
RsZ4RzaxZCv7XCUkDxumdQv7uDJP06mS9ZSLg4t7ess080d6jAeDrtD9PpQe8Wgm
8vOok6E/1nGULPx1QaAhnSsHUpKeOyjHdXQdL8tJMcB9eEGxMtPylr56fAUjZn0b
R9drSirRd0nNN76RV01VVOb/5Gd6EcrfTcqLOGt/kMEZlxHCa+LWA+Bim2sad3Lk
MnNGUun+8RVxild84KP3E04gPWtrKTZTpBLd0j1vh7rKlcR6CWsU7Q0b+AZDXXc6
633YDVkGYLIesRKLZaet2k5O9+CU3M/hTJlSQOXLZoxBGKY4Ub7vEdhepCVKAoB5
k7mtMR1k0okp/QzFG+PmGkAiNhgq27oiGB22O5luPONpD8uV8gnNtBEzPv25SKxJ
zQXxJnN1tUp6wbEq1CAmg7aRJuOkXPrrdXNNecc9Rj8Q3JT3dP355t5pO+hsBalz
EMyPV7Qcmmg5zBadkj538Iab6gZcS+yPOZ3wVLczltRd6rveESwIzrRbAfqf+apC
YuwlJ/AkgqWmvEjTx+H9WkrRNI5HC5L5AVfAMqqss7PJQPRcYyHS86ZHKVnKK431
51C6jFe0WPSQzfja5MG2nt7ubIKdnx+RyBn5LMV6dF8kr3Ut8hTWlb4qnm4eA+2E
Lh2rUKmshSMX4YXEaLsSlZq3JjJMrGmlwizc7mFpdRUCMuoqEftSiOoEXiQEjZS8
UbEdl9UFfwLZnnvOvVNDj7fcyJEQMN8iptWVQKESluGB0xQHvd/T1TmsF0x15WSO
reC9YC1w/gsNt6+PHHzqJwKpkNke6d74IuBYOFjeuTVvHdZ/7h/Wf3HhgYwkMMc/
J4OL94I0RbkzacWL/Rm3oIc+MUfSF8Gl2KS8fiJJq400//XXhgKfTny27VCFUyiO
VZhSdMKl5zcC1ewKIpriQz/9T2tEYGrCgAa5rIV68SMSHB9AmLd/C93u1mRYcqe5
YSoG0ABwjyiW4LlgfxdKQzWZGvljarIF8AKlL1NBKVaybQzzprZccRkEp7GCSlbX
LMEgHQtrpRJTLOzhOZkxhLjKuXRuZLL0t/TUznDpCUo0ubYiYS81+3hhoiRLWdTc
kTYXwcz8Z0SljL3phLV67jTybBAXX1AVUKBrN0mE8s57KffoebNbUNjBvQO6TjuT
M0s3XmLc6BaHCjzK2nRmlC1PTHhuQni/vJadVJlWURUSqvM2FOOaNZiTUM8t4V2m
w+8CxEK0EBOGLtPrxw8DvQ6hO1Nm3u4mSM+0NflcxtITvTVtbR2XYDMsxI8A9NSJ
8QHqUbi/Th/N/iBJDe7GSmJ2BhL3nysZpidpJYnFXXy+CY4K8qysFjoAjn6+y7qt
zpgnB9jGGl3gxBzU4HysJISTlyvl5K752JPV77mByk4SXj2WqFLja7G0Ki5uJ1Vd
Y76akKm+1Nczxd8DkiE92cgZlWY8B69hNXGizfqfwTdVnQZb87L+a78EKNn4PKhC
VaBOV7T67Ne53YUsC3DDPBfaBrC6QMz7qIKImpa3AAHurELsQ9McH57KDUHj0/eZ
BfQlxKGXpjTLh4URp9Kms0lmRB21jjCGRZ781CQAYAJ3PQtntvQXLeMpoAwkpJeq
P5Dm9K6M51yzIkPUfVT1ePxtw5wO/WyTaZR0BdMA3UK25wDq4nStS77+bLc7RuLx
fzDn395qYDO0H6gZpA55VuaNQl7ECcSu4UdbnyQp7wnbrR3qLkmFvHP42GlvK3LW
2mevs/1uuvdXNSPM7NqQKXi+KZZ1rX4eB+0aC8FRggxxlweNqFkGKacn2QOLEKwu
PRlP7mIh96W13Tx4TI6jN3z+taaDlaDbqnCnfrKnEnIduz+Q2IRPsZxf5IjrIeGh
jn3kD6OxnQCTM42vIFD6mj4/khIc+Ti6XBBx+yLlOuHlPCb5jm6W7gl6+GBhoWuv
Zcd/q9wcXqrJumKfKNq6SOh2V4XxnPRwSjAcSrm/h0MKf0nLeeqazlQhV+Jf4Jva
z/xsBgU7fraqSh7E0cxwArOru1h9agxxcD4NlY8dm+18uEvhVr113/RlsC67/b9U
+8P5n2yM0ShpXeqE7lef5ZfUqmurpyu7xtzaVTT3R+y9dOU6FI/ncunm/M+SrqTF
6dX/KxztQZATlCoAVHgfeuOODeFVHlLA4f9da7lnUJYQwPWzSO7zlPKI7cPMZ9qF
k2sZF36SZnLTozuUglNc9jU+AFJSJAzSqbVpM1IS3/5QvNhxsY3oqwUx4ZaVk/AF
9qiSo8E5zk4qIn/JCaYI4PLKJgWm2gBY2KSx4+BKJA+By05fB35/BsXhjHB7J5Zv
sSUNmbcrfOqf7VXuS4lnBszFUtVp6C0A6PUxn+Yri9vujoOClabnl6sRnEOz0awD
gfriyEg5nFXj8O1/zzsVofIK0kSo2PyTg76C3NpDYV1an3WoCPFs9tnW0jwPYqrs
r5VJZDrthOJljQvl3UPFkpS5gl3LDLmJXU688bz1d21+a/As+REeJzC2NkcKeQPx
jPCvM0sOWQp7BKKTbhTo3AOy0laBgw1NDCql3QXYifbp/V+GqsJzLbGeF8SIi+st
G96sc5ihxu+vcSfom+M9TU4IlwRuhbffVhPUsPk7jczNhP0X5HzNRJ+g1JFmemcd
SabtmGLgma5xH9dB/A9O1yuAhEgTPVfArhDBhEOhp6U3QCEi0oxtoqQIEtUXSUdu
jM5EnuS29uPEF8DIWIOgpZZsnGF3C6EAB5mrAmbEexkAk75nUoHVk3gfbmdmVgBq
uaU1UUMh1t7jYTsBhoOkVxMWuvJDL8eB2kVp35Avp7AgdEOCCBynj5eeXzj4gW8n
Rz1xrhta8QOy6t2naTKkQdjwvQ90/7hJBiKG2vEON5iAPg2CpOzS6c1oBd5sXc0p
2O/MkIRtJu92Ug2pn/lkRJ44hytx1cjVFYvP58kTybBM13U02Y4IRvX3kY+QJP+P
UCwWG0UWO0Ei/KmgBDoMrhyvx8mJZhUzXjVYcIEM3CdeQuoEQHyMQmFR/FZrbpVS
kBi7s/pK1qU/8vdS/TbvBS970JCwQ+IS6oe9WrIvlbIWv6EiaP8Ai/FVF0r97xcN
br86995Wig1flftns+4zHADzboQL0ItcKFM9SGhlmVOPXHsDPZS5mJad5z10yv7R
gVZz5lzIYEvi6MgpkLja0bkE39Mo71cvzxIAvvkrD2XX1Ea9eeywG1NXTMjUx+1f
4eRzQqpULy3GcE926C5gf8ygSf/nmzYBmx1V92Jsk4ZcH1xpRKNl2HglIuZDYx6M
pYQV4g57OBQeM2z8sHegFjStbVeVh0Bntr9xKlqw5qrjj/yICuVvxBfwJxk6XGh4
05qjhWWmGhygZ3aiST3z5OY5ZLQZnM696uDYqErGcDUnDsd7Z+GjHoO9vo1p4JZP
mXXoBC0PCcqXSKb3r7wtyGLx/G+Hl2nQU0AR0haT1+ytq2Ys3QdL1j0ao8JuORBX
Eu5Bo8maA9QzkxckgJKksBDgySgryj//avaOiP8RjrG6IfzVOdHQ0cXeEGTrMeLE
JqtkWd0dMIspueFW9LvWd6xaDiA/X0rM81lauzkS3aYkDjiE4JK7gCQ/oER9wYeb
soFYyygPWrUAwjzKHZ2kl5Ejivgs0sWvm5279i495bwHUYDwb6mCygwnxEgMy0DC
aMpqP4FTk9GRa9UjLeUi2G65r28rSR6x7mHbZ0frodt44CrUQE19kdze+gDjFUNR
8GNKimLsTLr9BYedPp4/aTAgV9AMh3Q0dzl4m+aP5NmMCDtZ4viI21p5Jq23k4qT
+lEPDAybIcfoSvKTM6NdzR9Jn+B9t7vNPAbnQ9uTX4iXwOedgy2phH2ySWrfBWlJ
r8h4yd1oU+L4LAfCkVh2dZEAoQj9PEg4VA+qZVILhWXF1mxfHMC7z48mHVNR2EiG
kMPZg251Qz4W4yXzELLcXIduQq/aCLDv4W7GbQRQd6w1yplR7kjmYKY/j9xm9ORz
9Q2drfFn8Fmw1Wr9YLpnsOcxgkKhcRnuJuM7jjkC5uDBBok0gkwILgzb0UlUrZk3
or+4UbsCMZF+B2Gkjnt1vUpz9OJrsuwnO1xWXOCuJ9I07fkvOCqOr3i1y+yBmXeR
0MFCNhMafD0O21ACMIJ3Nr4mR5QQ4p8YVDtWxOwPIbExpggF5phc/L8T9+0gHvDU
Q0I9YeTX0Pd8U0Pyoa+Ux574DaegCVBpsPFOcMdFlHjE6q3WagNGlbZkkuM5ZZy6
truPK9U94rS9Tuar6UJwnOs/RwgZ1O84S/KWG3sZuA7zPNoLXP0U6+EusuAKEaar
ARrykc0kBowKcJbV2iNpV0fMFZQCTeySbHOLMjKZMXI=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VqH7R+SeIxY56oXhyE/WKHArC/GviY3FKz5Ne7V/RQH3bgysVzKUU32KIqbt49Ha
6TH/LrBAKdVyQ5X6XTpnWf8aJoSZosAnQn1KSaAHi3xOS1ub3HqbHbY/8Rq7VA6x
vniZX7emKTupxYuNkvUhIbbIDaFgSzHBWXareOSrjqKkyHhIyvLT/l+KUHKYoYMr
Pe8LDFWriRu2+GJ7WvjLQdnSQ4y2Ds3cc97cF9qxraJbpH4aQbCrE6vJ9FPhU15a
L5yVNcZp8CDkgfT+ImJXJxjF+q1HBgaIpnVBzY2etQyWPv3ekOyi7lA+F4aM2nZq
yhTXJu861fhAYLrkmDc7XQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8992 )
`pragma protect data_block
h3RivJWc8d0vQASbIa0PHyw2ZS0TOEBqZyZKzHqLitLvbMMCHcnSpMamH9bq02l4
Rkx0N0NqtDzO6enhuf8T0Pm+fiXnAo9c+u77K9lCvmZ40SVVuifSwSTvsynTKKxt
cO3bjJ/Le0DEG9J4j62FHDOBTkfAYd7PC7/u7Wm6z1WZx2I8BI1kKEOBOVIFhEh0
IKguKM2K7wnyJTZdggXa7SZd+Cm44CHZHAcTvtDH6yb02sgMtG8A6ARPWh1/SEef
zKAn1YIh5YGdQCnM8GitkGxT+k1xNaMXbacSbyFpwE3/1WRVkjypu1yqRjfFRCAx
YAHXGNQjVvczfi+t7gRf+btCo/mOS8JQDsmXASqxXQ6SSx0p4f21ClpCO+rV8KeF
njuCMlGEZfMl63NmmAUbtNFwBtGzs/BWdRZ0qP7RAnQdc/D/wwZQ4EjGJRvu3tFg
beREX4ckj23cvkgTybr6GZIKmTu+Quk1ws4pV/sjvU6gPTIBlD+FE6SqCfp/R2mg
ZGCRtvNvKFN3CC8qwoHErY3Eq0geBAWk9ZF/9IPpKfsn0+WHFwc4Rf6icLUPJp8o
bNBTYqOsWdA2z0sXEumhDE8yuWP4AsbGWqGicTV8MS/aayKlxwEYa5G0GbxYi22e
5AceJlPxa28+EyqKBoH8ZXPlvYZ/oTCpxWROQj7xnLd8+fwaSx7htGnf1Ioorjzs
9H+jOJ+UwSC/tROWIE212oYaVVON0Qq4k2rnjp+X7ZJb0v/jDFaW+2wndqzUvrE1
BmyVf9luSkNVTOF08wand8vsFhTBO+OyN5d1xbmLrmYSw0UN3znmrorhtJYWzf/E
qmu2jAXk3I0WR334Rnp62zYVe17i+8FWTXZMo2h3gYh+UaB5aejhKTBJB6yATL1i
Rxgy3EWKkEHik/pTMSXJrGzF6Kfi7vOX+9vqzqvHO8fAB+ZHiRQ6zs5sctE5v3zf
n8WJDrrEhLZvrGE9SQaknq3/KpJ3wR0Sf2ce6WOc3t7OJE+vOLdczzbsb7LQdIqG
xYQv3ivbt+GQeLAoDQsmhs0GlgAJ7kGm+4KHkUq1IsKva00v1BrfwaoF+y2VKujU
RSiiWzbSnzeSpdLySFNp6aM9+mzdmT9Szr9Waos6nnvJ5X4H/jO7kvNSo1C7Dsh+
Y5Z1E+cztcOA0+M6h7kTYTfW1dhid95RuXnshZI4xRCqzUl0M36nOQl2E8vftRyK
S7ndfi02Y2gU+L4AH+j8S+1NqGmV/3fWbPVbQ8OSVxFEsE8hvz93qnJi+nxuHlg9
2usXqlb2RnHb92qa8mCmdTdl9u5T/jRw17zEfcBQd+L6jVZt8WDceb0Z7FZufKv8
hYH6xrm5sHabq+/xMeBK0RGoN/CQaLhjXETkK2RcRyxTsQIIes073x8C4nKSL6N7
OjxBCMoRaMp8mzmxHHdMhYTS/UYp/eyxn02ywxuxqWzkNKL58pbG/Kq5nLdALGeu
6LA1RM0gcAFGV3D6h5iOxFMRhlOxqMtz98Pvu2qcgZ/MZD8PSp6H/FlZjVItS/6/
JJS6xeyWLS4KW+TNi6nB0z9TrVsXsJusVfF0p97TJ5wo+L9ROG2O/0OJUvwd11LE
T9ZC+K5+fUpKOyNJ+VMHhuberp8LQxAajVXJl7p0MYUi7ZQMv7UYnagxeYMmDddr
5f7ONjzsyKGFrAMhz9FfPtlEw4RzSPAjeAp0xghTv57B8ntSOrCVBzpET9HxFTXO
IueSf8AXw1bNzvaqCtOqE6bNEC4gm9OxRTuvMiN+jCPhpF/kz6wPlk1r2CGbMU9G
qedQurfDh3CsRL8zbOePuOhUauhaVA6UTdxGdlDtmFlEsDAwDMZOm+krLbZ5rmDJ
eMggGrkFplAfEDOua0eHihbyqhWKprRaPqUPev4iWRMO4LQKykAs6Bo4qdeGo4y+
s/+zSppkYFPJBNF5xJDAZ2r5WoQEhjlWkN6sfmtwiGh9e/eMJGuWsC9nfANSiCDc
VHtu0QqmouyCIo2bOud/NOYAlLvZdFvLs8iVc7c+DIHRJv+B42CYOqRz7a8wCBGU
MvSeLDX7KFN6CDfgkUys57L/Jf8aDkDbHKZiOGmWwSyHYx79ic0HoZDb3TmWhwyS
V63oNz0Bz4cRZIqPVfDTeaaNvtYo1ZVCEbjkX1NaKYVpe26UB7LqZh2Et7ub06jr
nRHlzkK0o5cQ6xZFrdybsFbGzTL79J+v5SfVyEr+J/VU1RNdk8YqZII6AAzSHcMO
xV9besNetk4n/17BybTVQ2wFQwaYUbb5LJRF6EqFkvGoFhwa5wyeo4KadgFnJ7uX
+5xS0jApD5qgxnmSsDMnBNNjYYGmcfDS+bM3fKSoaGdbi+sD6dKdJOELlwR/paia
7g7sRdpDgwW6FOgwVBEtd3NmFBx+LJe9OytelLJAgzc3Mn1BSMKo4SHMgrPiqLOD
nJZx4o9KZgHB2U39tge9GItqPAXUwsD1mh+dEfMlmOxT9MFEPeMCbj3IVAOXhrPe
+jIg4kBGDJ6rYmprLPvWX6CAzQA722b3GaGrDjE8nUzvY9qSoMhrukR55ToLHgbp
JtzlvRWcBu/nVdEQoowQGwkkb9/EwgSAoxpC1vAQZ7cOOxmTrYjdBbz3FM0IYrof
cZCsBjaYK6J+lEl6sPRp6vbH1AoU//DOrONDAqmcpbljscVkxCGYUoj3nYUpxhVL
l57ieLRmKARtooToT/HADR5q5bHGWpMHGFiDqooIjKBgyCavWc3p6wCjCdNfSl4b
NironhFAIb6SicwvvbKYTxa2BB60w/cfuPc3frs/cLPR+ctI7Z28sjmRGhwgDB5r
cSYjV1Dowu/L3nu7CBevWODxfuXBulBB3WDbFQWi1iN2StVLUUlNNcp70kMBamly
Fg78VNF8sj3r5hF9+BQU69lcMHGX5YPOkCXqT5KlW1JF+R2Te3cTSyjoCnS0xhjA
7IpyIgso+u2z55BbWG0G3w2KX1wXED+kPNfLDEJw6+UYAPlz2KwmFObtPBeebn2W
ka61MYpJ7zKaTkWUueqBxOHQdVmZfbIDLTTIH6/XTr4iCISyIGdz51FNBzDrjyUK
2agMPf7+HimfTfWOU5jJsWSAj317WI3DNNHywXS6wAYx0DGQgjTnS/EUTjfDtQLd
PWxAryDOfRVzwcUYitsmVXJ9EvD/vhlQWx1yXekMNz0cJ/T4nW8Jav0vdNUt7DN2
stuOLMq5k4iQU26hzKcpVpzHQAqR3UuUZJwopaJv/QSAggnQ00Zw4FsVLo5WcjMt
d06ZBS+lA050idmc5lELuGQTv6VuLdW4nvsL8jMUocYbNtO2D/OcFBom8GjybU4W
+gN5iPGIwRNIgzVgSs8PBBYWSBW8k7x8hRyBJyUY+sojtPHtWdu045cEiZgF/pU3
UcQ+oEmyepeAb/k/AvhVB05HPEKDjnPjYz2As09vfSpqRAhmdvYmzUzV+77e2ouj
dhZGqSRgKgjbTdFpPeD5juWK1/Hy0H1uyWoqhLkisxlnt+1XzqnLdOXLUPPOrzal
QOdf/1BO36duSEQioImOWx22Ck0CiWrx3nYfzlQt6fK8p2vDjRWvyUIZVl2e8QcJ
9nAGuVdgUCxh9WGBAbg1Y1bO2th73/0RKnS7fA9KJiaoAQWtMRfARfV/vT5Qu9L0
tLVRWL9Kbz/0gOv86LdKNMJ0kUbmsvvUpgh8XxUNGI3CBGy4c56bfq4W2bdLEh8o
Os6mINlEK9pJftoDXc7VqQq6gT98ccOKTP5WzjkeEHKxVqTR4xuJHHe+xGPnQ1CA
v2BtbSWdVohJlfQrq2+DLz2eKs16Aed42m8UFRXzOXUpRd2FPpNV7FL0JyVSU2hw
2UflVn7lHXariVIQffPWBL2IqXuixN8K86FXjcyssb6kikJkVAcdBmcdhb4SUQLG
zMZauFR83FxnDRR11wf4OlHzbwOSlwlgzwBc6Puo7R51FNzDT4DCRqTarfJB7sDp
7VvvE16HmwJX9Hpw7VtmBX5pgZ5HnxrWaFkhvBQE/CyBKWSXgS0yoaufeg9KV8rz
72gFxbfX1iSdyvyKfFNjV+sbk5Q6v6rTG9qjt1gsYOrC/rJCDAABO6zjsp19T+qY
hp5xpVp+ovDzt7YHcHyh+OdYMGa+O+tGhxihJnLdBKk+9q14DgvmVAAqqW7sv8tZ
LVUjtrkF7loWRYC3/TTjYJRouUm+oX6VWX/aHPjLD1ww/28Vo1T9YRFRhGmmRU88
uFYXjEOhbHm1cqXD6tzweKR7Y9iDJbTLaTaJAWb7iJ2TNeXxBWerfDwzZhnubSI3
hiZIATWo4UzD7i0jIvruwHu1X25EtSIUvtaQvd8wLkc3qQj7GYvj781uIFy2MF3w
d3axpNerGILx6biQrhqbpMGUA4iYm6ZsaTbIygWoF2KdhojW8UH5yh8V49u9gqRn
XJg57MVLkhnJ+Vf2dg+7FujG4cwAg27q4Y4qEmp3SuFJ09QjH3fvbBYDF3vMQNS2
WhzdMeVmH5vxxroH8PWnABxkDsMRPgwIWuunTeS/sqWg0zo6+Vp+Gw0+4NilSbXo
PVNhT3E55wAq67NVMDwTWOrQ/Uv0rn/zNJiWSNTyVqvofTjNni59CKmYk2Xqd7sE
bpuMQjhDkhpi6SXpGPBKaoggKnw8Atqbi8/j0nYr0/ADkguG4Qil5uoK6J+7A8Mq
g3yvq28qO8YM2wpTZBzaVlvn48F6Eg4OeiU1w6LJceX4vrRgmuvHHBHSz5p3k9mb
ccVxnKxBVQxlgITQUfzO8aCNxEj2mn22ATVF5ycoz9Zk+OR2EgV5HTWx8U4BcoG6
lLr/RLNvuYzTNIycmPLslklQRzkw0UeoqKmVLTOIYYONWMhZQosLx5K+Gj5/5AhT
wGgsr7RsoCR1flYUFVZm96Wxs5Eq4YNTsiCiF3RyfxC9MTSrnXSJdxmIMfIdQSFs
gDPAeAVW4PyEoEo15AVCEY0obl72X9J+Zy40kFcWWuOt9qaSyrUMaO2/OcXYfPwH
saBuAcn+T0M+Kdo/jZEqZT26NYUQlwxgSiMrSgmrI15IczaxGJJLMjWq10Breur4
LNLOdUIv6tGf+bp0qRIAiYq5dvuMidoTaS6+FhdT56ZadlmJCmp21DVrPiAKJ0wI
BgXoSe/W2sFqE0JT2mLk1LCPVxRlCHdb0zIGbTHtaLfmCObLFcpco0NLmK0CquhJ
GONPU3Lo5nDxChNV0yIXRLHJ1v2SdUntX/91ZL9IU8T5KuyaZ78e/xNu1NOovsOZ
a0mPvRIYRazdJ3ioRjCLskJINyrimob8VaEao+qfMGUBt9rafGKAeLI8LAPBBgbI
CTlLE/6Q2fZFyvTykxQ5uNZq2x5S5jpzDgNzvEmT9PMf4S1I8OmiGBaCWXDybq0Z
E8YTnil+UDX3j+x1O7FdvoTEs07XKYXwHte0gvgaxzxfjI1DVW/ON4fTuBpLK+JA
CZFNbMMPxxvI3amot3poeP4kxqM2WU9omKjeP5ggRsQ4k8yXMybS7IRgXMYWBgJK
0PNNpStLe4pUMn9xQIomP6NhzelusVuf7yWdauIj8PZc6T7bZzAQj/Ig6b22wmD9
jaUZ/KYrs+tbl0rgITBDt+klrBbT/kyhS1sEdZZ+78Da2xxqbt6JP8KQZSXt7uB8
/sfElfg4WRZddWjDL254qT+pguggsNGq+eZCe5zymY7anheCu+UTBbszjrpAK5OI
BXxotoREnJJ2j3zibRPmh0ZegVzEvlw8BE8+4JXHdLS+rjG9k472Knw17PYtGrt1
/TuGkpEZnCUai6RjKpNfxeQ9ZF7y097HRuaeaI3qk2XXHwYKNh+P0xXfwHYZX5eA
N2Sh/pyWlYNP68L0wW7lsNjTu42V38uuO7xscr6gCLooOKe1CSPhIJklM48FuYAS
+zpWcFt9zsX5cGG/RtQh2w3SQAYUkf5lr1C459K/NqgvJFG73I1ZHzPqVjrwBnTt
jJvMsaPj2TfgW0lWY6z5+PhKtVSTf69Gi5kGHyu+MNLct28AUPXDPvK0Y259nJWv
P/C+dLkcZJXqRUAsUwWVr05oqmMjV2u7BSZr5vdH08lcDFqvbImJDhhol44I3kYt
YHFZmxzTnxb4EYfrOxxKzw5azSDqZqo/14lrExsNUiRaqlwj9gHED3frVxasXg1i
22w59o8x8beCMuBzzjkjuSKyZ/P7Jzywwa0bXU5p/IH+jylKoYCJVGO5M2SxoTHk
X1ZuGhJlnAG27Ct4/NoZ+NKrXZaxFoJvt39fP5jcyU4Icjtt2rfR7Lgtl0A/zmcq
P+qqCjS9szvoBvCu41BsPbIZVqW8tRzxxm3SuJtdixNyZlKeW83PhT9DKDS3auNW
b1SvSWcAfkXD+1lRutpZ4BGeDysVFbSq04iSIoKZGVuEVA2QzMdreq5qfdBwu73T
9m+aNg9Ayr/UQKDsMXTmgEYCHE8LPF7P4IegCAhcSTaW/O8Yr4YLEdapHejy5ys2
aRRQaxpKDT0sb2gNIasuH5jS58hqxfWEQDSys9mJ4e5I1aRayevZkoLN4qdVD9D3
awNJqUA+EyLq88HdrSvSGE677u083pMOlM+53FwJtuPx0a+V1JuZwiuE0nSfXz56
I8SwwYlvpIswUiW+U3yl1YHMmdYWqqv4VuhHmRMGIvMlHgt48zEk4apTh3eWUIkq
0Rn1fvId8e9sumeDqB/5t/6Mq43UGTrRaM7A3QjbeZaUE7XjEYyjXC1plM5fwwi0
cfeb/sUm+hyxDXB9pHEHQOCC9W/UHSN+2Dsy3uqlX+a47MpQIsNeWpmHcMAuZ+YT
PX4YMxtv8NnKLgOCIb51DPYerYXZep+Gd15ktjoFL1GygXgBo9jCBrWBFTkcOpyI
jS6fliTFiNk4H0qPtcFdsEKitaeTzOIoD5Bih6qBsJzy5pdy6CgatIkKZCTZDfYI
xW7BDn0h/2SmUmwVoMrtz7Y0fbtItyY1bluO5wn9zy5+Mnnq+X4ObtFZsqdJyKts
q9Oy3/TKJRfsAFfonpLMVtFm3ZOYjcNHJfsxzcCVaZgm4akyRVSoMrllM0sETE5K
jOJMsWNLKtZFeLVagQxX6kAK2oCPY16N3xHgE8xuyyc66H07b7tqIO597FLOaA5h
2gEpFuD/QoZ5+RmugxVcSxmh9n9DyukV4bOVMoAAp5lTDVWsQb5ki+HqwbtBilGg
TD1IXkUxuiXhxEN4+a5FXYom2Wb7JAB5qZpN01KyfuId9p76MvLcJUu+b0hdcVDS
3PB5dJKAcGTZVXV8JH2B0K16dI0zq8LWlJU5u3GS0rP2rvbh19hWPGvZ5FRD3qT5
D/+4gUtVXE3/k1QpwNcpUE4gIbBKpyFIzBwSKwtNEHIiA/UVLAOKQwLFAFnjNkEP
am+6tS28CejjzjGuPzp5oyjXHURPfozJjKkMaK1pkwxrwO2XE07Ruy9JFZb2HXau
rUA+H8tXQeT50NFtYgx7gzIg/warBz2C+kgxz3BcRfhuW3Gfrz+z+aWo4HDqJlob
N75gsBEIwDiq8FKLmUlvOACxncNiPRhrkQCIZA9weC95J7wR6k+2c/QKLVyRlgmg
uX+q5WkgK53PnKzhFYeDwVR4XM8SxxMUSbqNK4KDmI7C3U7TKl97ZqLftWOm/vL4
WYgEoPrNAQ84Q2kZY59j3wZjfBROqpw3UOCGAlhNGGgquXCZ1TreRZkTE6at24yt
bikDsDaObI4XD/CP/qjdbiOP4k6n8J9I70nFHfytT/I+JI0PttTQvACDGq7OgUch
GoIdYVxUqy7yXxtLRPYs7bbVRI0gB6Fjohvg10bKdh5EA3+/pu50ac/+TGF1WCF+
Nyt/+dipObrniGFj9eowsv11i8W3haXoruZJMK25SPp+eFypkAhAt1ZNlpN2k0nH
UOcCuCk7mR/o4fzZal2r2Re6OK8L39CJXuC0C9JKcJe1P9cJ0oEgap99eLA18t5w
Xom7Gnlf3Sc5cTX6yz7BKY552IFvI7y5SMV+xkmln/5m2Sac617UzmGucbZEicDp
SYyA7ZR0hnMA7G1fGBJYOj7i9GJqLcKt2AEG41XepvE8FBZ+FTflKOB9VbH+RBcw
iTGZWInqi+SzjQTSeukftX1+gNvdL3LBucUgsRcYmGmqgXChwWSOKpLCwMG8eJuH
NgmeIx5Vh1Do53PMWis/yqh/9TjTA434zi82COBTjlMWd4E4ykYvCQYw1XJ6moeY
ghESWYDrOnMEdc0Yv5cR3+0jiz2q3XalR5h7pjz9uskIo6KqojEH5RJrZFONp+Eb
KWNcsYT60hb3vw4SEck3TQnaSdted91oIAq3rRuO/Pj/P1WjYvCEVm6YYtl3yOI+
KGEClJNjgmysTuxJmKoX8P9fPAX6GAZmVWQ9NML6skIXSoLrvCXlaG9NeRbUFNo7
irJ1DfpfvDhIMyf6ZZIzm15Xfv7ttHJc7jKeYUyhEXtb0mszlNvt2W3V3C+DsRCj
q1CEe5sLAlcIMw4doVKFtf+o+t3re9n3nnkUkJeecyGckMPgaxYQAPvUoPithUsP
o8srRG3unsnchyb6lbVi5jy924ochGheYmntiF7Bx9KPvh5xSrQKnveN0nR04FZg
Gxkraa0kNinXRY5BZk5hv89o9v/ZoQV97gSWZKUQO7MA1PUV+LPoNn76eFP8QSF0
K2zvGdbf4XJkuC0kMTBLrXgdMiI+Q2XNrDpDwZzQFy2XCBEO8dyfWUrDgmPSFRrP
CMWYJahfix80Ke8WbFYB1JkgzxftMymljt63MwuaZvB7UtEO2KfGBk0ur+6IynTv
X4qioKGUcSc07L54Q4ga2OPkBIolUokq4WnobaZVJnO6docs86NouIiQSsX5bcwD
joyq2fmum2KtMxrmYMm8h2FAH1+Shu7L3E1mB3LfFgKr1PR+IwM7HnasH0lSC0DN
hVSjDkpNQUuPwQ7jOTIRQrNby1i+Ic0upSE2nkGFJAQF5mXrCdCzLN6y4BhuaErC
DQr5CTk+/MQwHghCSc0gZLCC/wgxV8gcxeaEGTuPDaQIH/b8U4TE4p8KpccgI5sN
IjM/REtendlDSzvZWHMDjk6c9qWO2ltphTLU5VOWZq8FiZsAQr+Q7c5AjvB5uc8O
JZrs57PjKHOjPcqhhIpNxJzwG7vzDz5hLCzhzxxlHHYWlPVEcOJin5Jxv0KxDlnO
FWn9d5R+zND4VvMo2lkPKZJFPkWo0zgMsGOzaV3FaXu+XXY3OksykswvSzEjieWI
wLk+uFomIdgcTdaGoDJmaspwRpzQZDKqGoevpga+ls9SCoGIB0IuSxpsaRzo64w7
EeTUMnnODAKhzQLU8G8bJk6tIbEHAKT//6gukhq0m7g7nyJhc5o8omzanW1QmjeI
ct4X0Yfvpz4J7FANbe/fXRkUHQICBEoheg7r8m51yLEB4cC6/9/qhgQZNBTA0TMu
dwDKv0yWjjd26MNR2HcboXiFhmUuxH0sLnwsDg2MQn9eUF0fXCJE5eKHSamnYSrU
zMbj9kN4zzCxwkxonR9bmripieEjfssISRYzjs4oosDHF56NBA8DnzqpPmt4/E0b
L/s+FlH0YTbo6Y1ja4fQHK5/fQFwA5nk1bP/gm3TxDQLZWHAuJ8x7yLOJ5QRXqgW
syXvmoV/maQRFAcirFHWrYqsl8WOSsJ9/kjHLWsO0gTMLUAw9uVuupi0bX1eU2bB
YT8tbnnh3ljHiZHxBE/LNyJcqXV6itCjXS1tK+50RorR/QzNzlq4uctKuFvOlYlP
HAiZxBxxM3KT3sGOadgvO+1uGCZ7H7mvG0eWXm8WOwRIuXsNpdtKukmsHNLcNMag
ibAfrsgf7RXLHM9ZDoWN+A4AH+g5L4GnfXWVtY2MHInU6+fAVkrD4tZmhGlaqNiC
srG17tLmDIPcUHquyKldX5SiI+gOeE0ZHCidYGGXXxWAn0MR5JnToZzNKv33pUSw
e6ib/mq1n02w6yEMzsZayG3wGjzuqEJ0s2LNnyW5p/aKCEnLw8sensGiwTNLv/vY
v66wXbkJYaPkZuFdxP7Ai2gGUongi+nTmbD+M1VJnhLtTqwX/ofR6/8l8wQlL8Ld
FsERdLPlZK3pwb5cCJ8Bo7X1uSBc8iw8B1vwpRfsTRvD/jD9eXfZJq9hBY/Fd8Xw
rbPAg+Axm2wkDO4oSZjXXogRdV/wD3rLklBMPcBvqTF58OjEAbAUIz8LSlBelZHi
vrBetUeCtx7W1aXrGADqQl9AyUU9hOYsRNzzUdcZuQ9itzCc9VHzlNshGOE4Zv18
nRJkHfFaOW8phrJYv5ujjauWchuOdaif6oHmU9Cb/29KK60s0NILXOm+XHX2FAAz
1/qxqlKNLLvUe6iH/7pyqb5Lu9K5Y08nGcrYq4p6EDeX/PJz3rVJYve9lMPvlerU
EK2gg9qoGo8n3etAzWxa7MT9sbmwKfOmZFa8lPqPedldS8mcm6Q8DqSL1HpvgBA1
z5Rh9OKVYb1ZeQQLbqR9MEVgxqmsTZXIG0w5L1rO8syB0FogjIlNIyd2TQKOVqxf
+0boSG2szyS9fkG3qNAxotyNWb9tBoQ5B8e2t4k5uL1PRF1KlY/uFSEG4hNMdkyF
bCU5WGcsAZ3fGoyM0eg6j7KzRma8WIxHNjTbnKpUNe5GMz6hIPl873hUgxZ3y6Xz
R1FKaiVHYAI4w2/1yDYPBR28txWQKL+ZODfMsHnywF55KmCwtlIsv3RmWarcLCeW
lZAF6KADhKHk7s+aR+3Ec9TSK5pqNxjFq3NF9uBczBdlfx/djBKtTKCqtQ+h1EqQ
XsNhVDjoPcdSPwb9ozjq3LecJxtv+D0vmYqdQA0YqFnOHr9mctv3B6T8YYIX+Neo
wymlvBU7uCwXRoul31O9hxwSs/ivixGPZ4/HgTqpzMD/BMNDAhsmDDPR7yFekypq
JHv5EIy/V/G1LpNc78w7XbK8lEFAwPfr7ljARZV6Jc5CDoeqUzI74zmJmoym30vI
0+pK7CCQg6fZGXhXxZa60ryCX4DNrm0RJd+ouH/pgOQU+pEbRAvo6pXa4zcugJfw
cc5TIPQc9M98m+Ra6rltZILt2lms84dGOOqYlyw39Z6m6yrqww8irrCABO2kvHjh
rlDJ08wJl/dlUf6zuZR2/yHYCrgUI7k/hHlkAzd6mTBGxOj/7KsgmGIYWs0K2XJ2
zjrgd3lx8A5GIld8z+NbsawxH7JkYGn/h6avZ7MQ5fOgskqmgl6CTPaY+0Kzb9i0
j5TPCYUfO4Tk4L66hWlTesIaeurlW2qMoRPgDICiKcR4FlWwOWO+ifH0eoddzFt8
/so0f5NRWxtWEy/LOTljj3sYEvpDRqrcG0RezUNTpuOeDYcKq9YlHzq9K0kZAfKy
cWAa1Dau5Y3ao4DtjbC7gB2lO6xom+UqhGFjPA9+lFJHgM84KDDGfaZZHJR79VfQ
hv6AbEzevHVg5mutTRmv7jPgZgCT2PqlR+bLfoMJ/o0JO3fPU2AHTz3zEz3kmf9g
8hi84AUvyfnBdEjq1sUOOj5KiPcOZBSVIGUsIPhE+rww12PLOYNxgMurj9Swdxhe
8v/WyvLLrszY9zyaoaiwFayjSA0Y3npSPQ7bJ3nVrUg9x2HCxq6uQJSa7b+nQa/x
DDEr3BtG+ocVgQ48pdLzKPT8ukzTTpHLGoduaJNxmYpUQ+YucntmkUI2gknLRrth
+vQpyKo/qTB+zFcpOWWJbZHpEnDt2KwSWDBKCmSEVP62ITITPFJ9ochU3BB7mS4G
rLq+OOFqSidHwx0TJzRXy2YT+C5qnf3Yg7w2oP37bxuE1ispNsOxlr2qq8BP95gH
3zrrjcc3GOV4OgPc4bEHcs83/+KwHzjKi55iLJnVVUpYNBvl5JypwdECKVv7DRl5
pJXw/mjOf9OPKhfdaYxdVf0UgoCU88A/d0l2w7QnMUHwW46hc6fqKTfkh1gcNBM8
YHT0Mr2DUL95xpkKpnUSOkUCnzd7i+cFBIjo8jFHLzYwgj0QbDf6QiKp6Rb9xngd
7iwzo+ng6U9vh7vRBg9aOg==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GDu25vFp3dBiYVdCKqTRWyLeRxI0JSQukAaVw4Nz3wNgF2xUNlxiwEHXLW9kQy+w
PUAlUud+qQ9K0ukb2cuWBr2inUBr6Y+3eNvK+cTFn0zz/Rkix0NPU4pd/VGGEnHQ
Ytq2QZX3K5fm3SvNCTfSUW82sItW1Ywif89g4pEIxTiILMoOkIQp+KWPA2pQ2+EK
mjdJJzbru3QWSpOtmd3NKQr5RdTLLMwrq1nUIFPAzQ/JNz/98jxjStQi8FcBwVI9
ngIBLihLpfOmvuUzarfVMP7b0UIIPmyCeFt1PehcjYzUHlmaLWtzKiE01PkmJU/L
UVY3ZrweVBGH1taTTjKi7w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
T1rVeabNOqK3YONG81PxC6rROJ+NgZWC7+Yab2vPoR0aBEwuY0Zo5yIVbMPaewrH
eROofksE3DcN6TUsLDI7XCVYariCTvFgpnUYtLnj004RMALmN5Zb8IpUKohO/RRf
lKgb+UruDDdSfTQoZksARjLs/M63e+zel3KoykAQOkQQVmYfuzEp19uUfwkKDKsS
WROgluoDPFR2eB85W/ia22g39R5fOjnUkzsNqzrVEUNEMnT1CM/ydwMFVfLjNiSu
X/eCRSXI6FNm45SS/GGp42fILL6Og18H19ihbTipIgzcy3Jteo7ZsSdOIOFSKsIY
/yqkeXq5gUTXCaqYCoQnDbjOHXcLeUUpk45fWQ4KFg4uKz80CqnA7HtV96KutC2Z
v2iFBjWPOJ684h5Tz5BdI3X4ll2FUql3fzCUzMsCI69BbodgzyM8QpKqQGmhEZ0B
W0E+faqmneAe9PbQ+Ubg8qBSXM2jqO8sk+rXDx4O8MROahQxumWpmR9Qvi+A5BYl
jlOgVuBfMETVN0gqseWRnReDQIhM8ntRiQHcIUVxbrnpNSJjUDzArie3dhkijRKP
H77N6ICzI+qqvHql6OdoJVgCbiNcZa1Zb6f6hdoEadeASwN4+MIqrwaQhRnYq0be
bEpU+UZ4zbCykFO5r9XrzMhUhItk7qNb3Bh2/EGdVDtI1jchWU9r1cCMHHLNFuzZ
BQ90i8NdVva32ogyYYHIJGwbwYaMrs3kNDwyj8p4KDCgdVbgQxA21RZMv0iRoCNf
fD8Eh4F4TuftAJvEDwQzMikhnJCrVbRR74pMHFwY59LWa4X29fNOTR4K5foapT5e
tAtxMJAfWPYx9Fj3KoFHIq8Ez6l68W9X2rvgSrBIwKBPChkwWWsw5qMAD1veODaE
KEkBZruBApjWGYMTLM0a5/a9i1iy4/NH5Zq9ZaBC6kZs0NFzi2Jpd3QElj0o2nVI
w+j+XxAJLEWKiUO8gPPVrZ7spWT15YvZh2RjTlRrWKuHDmMQ9s41hkHelOow7Q32
E5gOkKaXO6BC+HUVdui9JudN5d08vvsoAQzrw+CP9e9Q+RM+ksnfbcQk2GNWPwjj
EGyKF4XNQpQlCzAMZyXWNK9DdV8OaaUG9aberEIede1C2ikx90SZpa7GzkZkovzV
Fsp/x43DhTEiz31dni+txYwIbt+O57HQ0f0ezhR93GszM7pFoZ6NFxbbF0deA7bV
lqxoml37m8RaBEwtfaAbD7epGvJiaqRcqelDx9Ey8JKaGwS7G8rZiEjNFfAFpOcZ
6jnJ6AQfz9Ab9XYPvc1CTJQUdNvZegXlgzrjA6DSogvcYRMIe2B9BtnSWv2gglb4
K8x7Whypr8ZNU+0jJchLkiji3/7fraEaxJ8mFx4oBppfDeIFWlHc4hqKtlGzHTDE
oxAW4S1dGY6JuESHWR79u1eCrY3A3opDZoIqEKz9XvrjvxQTeFRfc0DAgs8TevQ0
IGsQ2v+C5ydsYBqlx9kJdzBpcGTSVemz3Eg4QLp9GWgudwUOSqCdtPawXRl8Ml60
/S1BXBbA8l+HI/ArA+kfDdt6KXL4p3ES8IllNY0H6U3tUrs0jh9nCsBUMekkUMO0
FBSbUSeCexH4f5JD4jxsJsYQOVV0PaQpmsDEruDMDXw35OYJrZaQTmGCzv7dw8P4
duxQPuVlooVVDWxLnZBvkHGTVkUYvpsVwxN6JWwl0iJ4ATG6XTSJCSU1pP0dxsma
WA+uJQpUVuBam0vv9K9Zw29+8hq0mBlhcU31UoRgKQp42yS9Ro0OMvk1tiotBtL4
gCQxgHt3SuqZv81VmxmklZMUq0j2in39PmzpA3hArfHFcH6r+uO5Kh07IJDIxCyZ
Is69tA83zn0C1LqX4TY8OGFK7PiunXY89+IMdS3HOxe4zqP51Xtc/g2M5YIoE1am
0hy4WkxcXAjwaI6ykvcJtgZzxOhY2FiSX7hZzXlXDinFjzNCHhPYrFAEWNSyEWfF
WlUFJ7R8su8W+6QwmT/GJQT/0LB87bcJNeXpiNz2Ega06TAXszevjjDD9MLic+2X
vyU1ZnwlFPNBxLOX5GcDGtNiqA6w0nBI9cFdaEdOHiIWK/UxQs9kAccuCmiIwB/Z
pXw11NDgA8Tax/TNlxQZ/6WYGI9mmXixFy/wKFMiaIGuh6X2qhy1Ul4Vx8n4WcfS
Ora2rHvTllleSYF5YoussA3Qq6TufZXk9Om0b68o+pTo7jE/EM4HE6qRpjq0/XaV
WxmGjiVqm59XCPodBOD3vKMbpe8DABg4Yd3RmXTb3Se6Bft71XXenLEb0l+k21QX
rfQUXv/YWkC4itSty4oOFiAvLnLY8YsGUVA9uzo9a8SzYCKw8LRZTwuelekGKqiR
w27TCfu/3Dl2St68AA6SwU7h3BFm/mOncvalt6Phk+KC73Lbrm3NEKfouXomuhVt
4NpKp08whTqtkHzCjctM2aozFoFNIRLLb1djmLx7gDS5HK79fukxRnXuN73gyrQI
XRzGxmbjoCqPRXgXyiDnmuW8T5yP9uCzjxEOLsa3U0vBk1vBGCN1QLsv1G+5Zp8b
SBcGnGjXIxPP8eU7bw9K0J80alt/D9k1n6IjdUMjT5FcJOl+QKAs3aQFTtarKQyF
aDm3tHGfeB73xmLO7BzbF5Ic0t+6FfqCyWV4NehUfMileqsc/H9ztuUwJlrJtadO
oItcYjtV7/+8wEC/oc7pUoUwqdXv7msqqXHJITWAiP0tvUSradtgi2eK5zqbYy9A
g59VXQr/TjR8EfKWgqSzL5LTFW8nPxL7QTZ2wDZgOqHr+NY7vh4QVWT+OsO5rxFX
deUKXTeEVHmwOCcOf085Aj6zzEdtIDzp1+kl5chyRJymFlA3lYU70kYUHbxIiYRd
4iALQWsJ8Ig3ephYl1dyMk/dmpfIHt+ui7brJNTAch4Z8dSh7Mg6cWr7quGYmng+
1py/az/qZXUCvzdx6ceJ/wRVx6ZnckKtJJeE4LkkRe68GjF2W+VUgbtPu+qskH4u
nQPLAaufRninSBnokUEFR125o5bgE5L+NBjnmhD8OGBGcgKjCBI5GpCLtDQtfKRJ
ertKWnQXXN6VJxCWeg2FxTyl9/WDhqze536XFd2lPqWGtWwUyA9beKrGZcQpIZxH
I6u0h0QRqulNnwEZul2EMiBX2iyCs1natsjE1BUqg49BZGkRi6pFh2Rwg3BTY5oN
PxKVKpNj+bwdNwgrIRxps6R4cl2k2v7tgOp9DdvC1HZQVuJLpc2gWr/EOnZ8XTwm
YpZW+bZggkV0sEg7GXJhbBTIl94It4hkeNurwoEaiaZkmdlbfSZqozINe7BHBEjs
iVyZCw/MpS2MhgBnLqM4ATdPqYVfP2Bd5nh8b/jjb18/fj0b0ILl85gdPjbKYYch
ej2Fritd8KePQ1dPdYFQbtlBSZa2+NQdPEK7lik9vA3YHHjhJ14h2rVpV6zJpsRJ
Eb/1Y6ceZ4DdG90jCS6FjvTiVLelOqrkYDcdB7IZy3AfjNY9ODDZu8IbYCwW5Oxc
obdwIU+BB+PQLqMT/LYMiMPI+qdCohEK93PJs5pjEFHGoOTHK52pFb2Meh7D4QNa
ppCn70YxsOSOno8pAmiM9kY6iUUO0tqMmfgNcJ0WnXzTXVFjqbx8obeOid+ryKlP
jf9blo1AHEABE2a/wK3raJ2Qp9Qyzkut5HeH+QxXcdeqxSUFaJOo+QyiIThmN6V3
O74UV/u9mNNvVyTnOqIQm6sqz1msrqKRPt9lESR77zoP3QUsoV64y05Dxg1tdUzg
qy17kHTGu9V3fY58UzOVuvh15hPQbrdCmQ0tcE9jo+FgXv7RGDWqfkpemUhakIuX
/dSOomA+agcywkx4nW/QeRQWPwAynJeeKzKvOV/tLeecFo7Plp9wKTJhMc+zUCBl
s4iny6ruyuJBIo1Zg9hSQx+0aHnvXQrZwQ56vcDaA3BxLnB08O1c+6jDg96g+paj
ADpcuMhFMbLQMdalWeknRB981THBmqUz97TSLYKe6r/AYh4Ap8NQe3q+lJFZgX/R
KAXl5RKKaRmaFI2llKH4geiYm4DhUxGlU5NhAPoxja+3uOwQo3nj3XGOYhiz0g0y
Y6tCeagAZD5hV1bEYuLprckbWrWduLuXQIrV3PsrG3lBpJ7azxWiAqaCz/SGjpGf
38RzbMh/cfrb0nJ06f1mX0c/sTd+4Nn+nPt5vIpv//NziDTpywEj5SsjPjYZUBMX
1JKqqYwiJpi+EnMMRQXC5xyOlg1WMwmFqUkkLBjt/Za7pL7xCsG54nuwf77WdJXf
0Cg3oO1ss/v3F90qJ3x/mZ+MwFziaE/L9sPi+/5CpCLM0QfyaXFezZZU58MKHGUD
KKWQyMMYJvwEKhfH8deJGNgeczlnS0VYaThWwWJjsjXtNV6XlI6nmX8KqBV8SWfB
CDIdZ9GZMGSPmWDNl6DRY5YW2nmTjufjOMN3iGjMqT01EXYlycq8F+bl4tHf9Re1
7iCit4YT0hnUm1tgU0I5E8fCRwhgdqoUkfd/O/WKWjtmrJHvO0p1v5EZ+Hj4QJsj
De5xluagD+svoooKvvRS/WvRk4o/6tNkO3pgem+W1Hr6NF8EcQzWhF7PmFWhkbHI
Bk/d6/KdqepjKhovzMped8mbf+lqrGeyJYCkTa6yC9KcOq2kBpWwCttXSMmp9ZOv
Tu+j7Zx+ap8P5ovJLpKj+fs+mTghSHjIII9h1XpYRgo5QBwyGHQLA8ixhfaSHxSQ
y3ef6/mAPXT8XntymzwS/Fl/HGu45QmzKle+Qd5s1d9dOijrOxprViuiHaxiqP+H
kjErfdlYX7jo01KlBuBYAFy1TklJTO4zIMfmUn7AQhtMUsmDx+1avlD2rvrP0k+I
Vm6UiK/AXF1dRA1Osvoa4Tjlk71lq7hqvKh7VuuuYwYZV96RsBYnjeAtJ/sjSfAZ
m575CbBUGDrsG7knvvCcZ5FDhqlkEWFr9T7UmQ6KR9UY/qNf605xbhV/DftctTY8
dDIcnO1AelN15XcKXQ7W0pTBWYIhelatgIKPKWoYQtj8q17zKtICRvbP+Vt6Qwly
/Ai39HNgP6rDX2qLHNye3x3SBw56AKJyBLUPswoQ1zc0itLdNsGJ40ggTQ6kxNo8
FG+JuN+q15YZN6GcNTnzilL8lMFXUxNyCWIxpczzYCE=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WFegiNLewzfD//YR8tMnuTmdg2CLUp0ZLO3341t663J4W51/8sBpdPwteFEQU3Y4
Z/DFATcAzkk6mh+ReuozhQGvvJorlnstAnpU+N0s1tM6PbvNRy2PijV33al1EwIC
gT784MepBV7gbcpaWkJlUa3N6Av4exBGFcGzv/XKML4pYlVG4zYpRVj0sVKAMoep
a9UkCKnKpo0A1EqwAhYp6u9F+9V3Xpa4esOa2GvzCFCufa7O+3XxI194WSsyNNug
Uw4ckQW578qsexouLInNF1AQIRdIZn8eTXy/3KPByrrXadqx4xDcM1NgHVpkO4Lt
CyChj4h4N679v8DYFDPKng==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
jd66vtGKZkGkfgDUTVKQJXINlMFD03VxjQHyXgtt8vfS6Qa+LPFhXS/2rKLUUOvz
Ax/B1zjWmeWOX4/jnlksiOdlnIKGpsmAWussxzzpWJrAdQJJxavAmjbrMH+flIGF
BKOMr3xTajh7wztvBa3v80alFwvSBjg0qRIjIyx1U8ZoBKYFfv1WK63+kslnUTxA
u6oVTnkx5BlbqEuRYV/kofjFnxZ+CyhGmcn2UH+OpjnjsyRr4MnMEr2EqoTJTZbS
/mgiz4PYVmxfCaBfrY/1ccbUsAkT0jdEkjvAfRl/owmFghZ1lvDweKdFfNqZSi8v
LpLfoR4bLeMKQkxRhKvEvroui+fxF6rqCsJbagcNn9gQ8fbw8+g5BaDQhubnK6Zo
ireJ6PSisliJ+h4DW0tRomrw6KtU/pDxnDTPIKGl6yzRxL8WZ+nRY2X+Vwz1SNgg
wWJd/z0DsVfHR9NVcgaSfoq3sKOiXAzfv+qk5tur6HjcjxVe2Ci1KpGgOa6HEeRJ
5WIBXtuidwdQDH+RAnU+jXCKrx3fbhMW0mT6NNqRH7kL1eYSLXHrwvZQCRkerzQu
MvTcMuo9litE/fWMtDSnXQgJV9FN+lprwd+lSunI5NhzppfKXWg7v5AqH+hQLuhy
qH+N4ymTo7od7hZZwHkE/A+6LTG7PrOwQGR+8lqPWYRyZho/0/mcL3t1IJONRO6X
T9CHmv54KIppY3+isk1uUts9sPH0mjby8vl0bX/rnmEfk9EcaEcs5lk8Vz9P83Qz
aFRfqKSyU7nFEgv45xTWZ0/e/pq2Z5pRwpHQqjsxx5jPoBaBjZSK/6FY23Y56AzL
7zs1ZqmyMjKKKd6HHB7eoTVXwBytnGb/HlR9IYbWiP9R/MbQ587J2Y/bBl8A9lCj
wT+K4F+AxsinUw4d0P/2plv4OGnUSl4z2wKTdIGkjt3iI81MisdI+9G/iwp1fFOz
Mh1K0RB0RGbYjxfWuZk1Spckp3GR7pCOzuRalimh/REMC1PDZt0fvuWSE9RfbOcQ
3sqQO61H830+Bno1PEyVt1YPk/tXVaydyVZ2LFP/2QaHOnS4AKljjVM42tRdfx7S
smMKUexOENb7KLO3WancR5mmLvXRf+dGr5lgCMep7TTN+PYMVDZWXyylLIZ4NpSx
LQytaGIDtDmBsr6TPDj40sM47LWNJgxg1F7WGWCCwJ5BPh30n0JRn6i4/NXeyBFt
6aE/1gmkOQiyMUHBOKyuNF6zIQC1/R6CFGPCjxTdkKCCIpdWfLeuxp1AO6N/QVuo
ExY+lJ0aa2IhzqLFh9xOn7wuxRVo7GzvdYOy0ukLbyPrTFQu0oKNJ1sYw2vNW/9c
SFNVn2mBIxxyiXpZkXjV2JWImYu2drzbSqbCSaGbYLRpQsus9ifpExWSo2CDcSka
HM3k1wM0Jfbmrkv8Dh/1rucR06pXyQeX1xXcaNsenwk5WaVZ+DllHjWVU6+gBYZc
M10i11yuuhUdn+xyaW1V67e0F3gUCEKCz3Cb81O6YLEJfvXWwNgm4KEKsnV/kyE5
Rm8xvm5SxS2cjKHcCDHqPr6Za2wQ6/8/c0fsFGqsL/3hM04hv14aAVRrPto13ecW
8nxJZ4UKYnSTFsqPgmSr/NCpKq69/wdeTfaYctOXlDtEllowagdNkONIzUyM1T09
eLm9L641Uqz81+kBHa4eo1n4/2S17/PAnxsQszSpnPmkpIJMagCNNqMSzQckCpJn
SqnE0J5I2/oAxqGSbaogjTHrKjSNOl8/PMos1Ynr/GSrOR9qwgX3b4pbER1BfxtF
kCL9C3BquB9gTfxNHtPKupGj+9XNaTpb/sjxFKgxrscP7fPZGvireMV+Kl6WLNfQ
nkGC9JcmkBvF9HYb4IBeDbMPZqE6mAZkVOolcPeCSFVA8uvqeFM+84SRs4C+9jrb
eOgvO/M3hD9OjKlHr1j5ie5ggLbhooxrdAE38NVYmZPVNqqaK+csdViJwEln/XDa
1oy8bkmLSS2HAhvaAE3Cxm4CfhtdldjoIapLa3mSl+J8ODHDpRMyrq9cWjKsHH5A
+BXWEzwpm+9Cg4JWlhGB04GzYSJvnyRklDZR6wtRGEAQfqZBeLqCQreZA7g7azDH
uW3TrS9Ha4QWgccND2fTm24XajCUFlxTBBx4WtPFT/Eqgc9TVxIx50QzIGNWFTCQ
P+/OHgM3w7SG+r0qJRmMIDOEBIIwyplbDAsoP7SiHWMQneXpBihi3oYzuluNb5T7
fOB+H/zMNACP6+/KdCuo6Gw3eOZN2/y/vemS86LBBS8Jf9kKHOHtUHWnsAvcs9eb
rSJpXL0E3DEiB5t/gy6Q7TlamL5TdZV083Nt0WcBzEgAGo0SnzJ8bb+r/WWMe/+1
47F4chBBvTStM6wZ7cnQkyjUnMXt+oguoS34WF3/0fmiInAkuvBHuEaRpKNGoRFH
tEbsYg0qm2L/o4IfKi+a36S0C6LCpLjtbxDgufDxxmjtNUBVLAW71CmFTiAzDMjq
QxphInL+qRACLAaKER7a370umHozlbOp2gLqAiZCzZnnb7lmoSZjqrTWsULU1gK1
0XDvIrXTrxpogEblwZpZbNh9oADGf+w0dNwtVJYhRgTQOaYuUV4pqJUR9J7XfW3L
SusiZE7RkihXTs5vd2y/XBWd89WM2fT5R4DBQWnf8Z7J03z0uhbiC0i9qKBMgHZN
ksIk6aBARFxdLFvUdxpC0ZLYVJ5PWUB30aI14XJy96p2a+gCYCQdxaHSTSeh8Zwb
IoyE8Mry96Ka4KouBXiQJOiOkIdeCxPDuhGUg4x4I3ISJ4OuRU8wPPYNEyEX/P84
ShIQlN5GPk9emvtHM3fjNBKJMT+R8XuUqc6xA32HxfV1XGXMPr7AU6a9bjFoJM2/
OJ2aBoRtWX1tqmVChcgV1cDWJ0XdvtkwXA+rIsAOzJ3UcybmKw5ey6SCxe9lNslB
lCQ1eMYD8/4Frq7HRTGk91Hbw9Xk1RGk8jziN+HLfJn4SahY/7MRYz25/CNpjYj7
c2oYoaxQcgczZfJzG+ZRjQy0BX/oVRMPepA3uGy0/oRoD+ibw/iW8eGvGwt63lxB
ecoNw071myCapFYF+cj9WtLGza01QVTuT4vBqb8u8noF3j/L8L91OKNOsjFtFpjo
VRVwXXReXncHYC0yKN2Ok4wVnKB+pERktpBssA+3/2PI+jAsZAA0A/OotwQ8dggu
wNnjKRTutR7VsoedC6gBxypNiNeB2LOpSZd8dXoBSzCr+r9fxO7Vo1Lj+Wo0Q629
Km2LKgSQlrxm66GusekhWP0b0pJ3vjFJBPoBYdxA6HXjcYXhF/07yp2TTVCFcZSG
ALhhm0TejKzeeXhglEPUQmA6YM9qx3edX4iFmO7iNhzih7hxQzP/y2hQe6dW3xdV
bcHktNH+iH9y8kwemFNUqZIdQ7idln408FFpnWZHSppRvHXvCCFQ5lmboKcNPb/B
77UqvzRn9ABG63II1D3aRo1eRRTGjsJ3fgLpFmLUkHKAkv066Xq7WZM1H/YB58dn
C87LQsR9+k48IwBC4wE5HIvxSKxnFv4tUbrgUkH5gDV2rrx0Ph+zyU7+4I5nNmxd
lMLkl3mrHXGdMfpGnec99PPQt6gkPxFuq43Rz3Pv1GvnRPcy4ZLczomMckTLdDXO
zcVnY21vF/rej5uZoSRSrC/3iTSlE5YnPnIpn4/tyQY8VbQBuu89THRW20kcmE+q
eNl8tQqAlOcV/gVn+xX2TbbV5Z5em+7cqHIaU8SHNvBiK/ROcwa9kZ/jrZspDyr8
zEx2Gp8nPVW4SF7te6jZVfwG0eCnzpfi+nHQCEuKd4eLuW7k/1FNMcf082E4DcBd
T1WDuL6Nwl2P4Yw1OuqAKYWWoNcT5grt+hxeJ+RIR7HiIzUZDb6GFYn6Ds61zicb
WrvC7pPja66+eI+1v6JzAmqbCkApkB8Wc27R4U/BZWlCdLqW1z4YvLZBYVCM8mVt
YUgLy+j3TlF9VREXYgzdkdzYaRiuh2J6CIblFgFmXEReB0s8/ISxzkNVU6wjmVby
xboVIuAtf0rPtSr+B85jPrUVUh3IHeu6Be5v6NVVrJNnZVq9OnkuXHBoSOR0a1Ni
QZzSBBU8fxRniuRYg8qoWQf5qoJR7GZ6B9dj3ITzb41sXpLL20zwvZFozzP8vDpw
TK3APTzqkbO2n7nzXWwW784+oKGYSogtT9ypNh77J8WrCVGIrghKBG/m9Rm7I3NS
G1xe0PRmJdWPJxxxccX6BGWSlMc2T0EHBbTEUXkEymn7Iye1AGgFZq0TkeXEoSRf
x0dPaBmkvpl1/hWbTKfTTn2EtfZQ9+tRlNvZ6U1lu6zUTK00wrvmvdVzYGPuD0Vj
8QZgZQs2jVq3slIcubJma62RWxefnBhfThGfMjfzpJ/YZXJugw76Txj4wAycprgK
vjvYfgc+EEo/TBLIlv7/Ozdx50HdBQ5O8csl6DuHGu+lJueBhumqswVDrLXNIatA
89VkP1K4ZgODE1fsWmL/nnn/TedT7y8/r8ucERlSOPmHiAr6zEYzFk2wRpgRkF0g
EcMcE72cRIcDf1YU/SjPq5vW7r8yzy4qqMF1Q1LD+Eu2KZ4bcsajtk8OlwcE5/FB
l44RFXl6y22s4YajahuvInxqAwlGL78Cg7hzOsTm+dyqit31nsde9MaGufERNCik
FdY1UH3zOIDjWYs4NN8S6UMNrMTnDW2U1Ov3Zt0RJRItnkTfsfcW68a6o+t7TRMh
FkBt7AJIgLOzns2O3ju0708zqnD/EqZq2kREy+xNF2jp56vbnBlttXUFN18S67ld
EMiZPliUV5k5HtTHRk6R9P93PQzkgmTO+0Fiv+k4YZBwOxIgJQx1pB2PxxYaBmT5
4t1+5f8iQxl4Zed9YAiuuYpDUEGqjAOi285KpcL0vLftgJR3BqURhWbTUjpUgse3
5ne2MpHW1X2W7mYBaLif7ZuMw8Zs0lfYwPfgchJFBacYiPL6VD8YqA8FlHPg9IoG
zl2zojHJ/x72whMjyD8tPWalzepL7PIfH25lbsLLVojB/Ix93ql+MRpgOPcwBy8Y
rzy5FWroMui36Fyn+OAKs6JFgKPhNh9OLcsAUvBipRqDTit8UyVQsMePe3lt9YAF
JdiSJB2y6rbJZk8vLWQkRMeKQGT5/ZUP3Wc2G9fuJpE7wmtRpF1FJVOEel6tf5YZ
3m7a8GPkBb3eepEqXTmJqsHg4L83+pPZBYtKBv0vIMkYdH+lVqxYAlz0eVM7QSPc
h8G+xug2BTdassn0ZOleQ62lXK33ZCLC4np3Q7qONzK+bKHIEOj+mqxq9HXw4/Tn
mkSXUS61zLLbm6ivKInEYcmXhG+LDqnxQbs/TfHcDVpCb+6yMie6pmCB52U41KhG
OxvnZSse3NMurhE0Eef4wtKWBZ3uIYxZKNTXUwHnoLrXBAsH0bX8QddgwL4fY7cO
NqWH7DvHrjoZMem1VKa+8jUKjepjCraXRl3Jc3/lg+f8QI9nhu45cuQWhxiDpTB5
TBYp6fZ1T7i2fhHkGXqwvsQP7ylK5XEJL4VCvwzLt9T/pU/+JbZYvNGkasD4pi3X
RVNFDlglfD3hQkTY5m7HB5cnohvVL8QC1adcckgZvZJVxj+5w9m8gNNIYiJHgFU4
Apmx+XnuAun8Tp4Xak6Ok1bC7Hms9FcU1K+sod6eIX4e9DJkbjjBskVoxW9z1ZXw
bIgLthokZCsvWLMXepscbOAV2Ek8DAIaEL3ICKlR2sM6++NFVhVxDfXt3A2RdhMx
JJsvugzve5R1lEzDLYWJVMEqdVWDVvLqWTCGmcXL8JZXhNYx6TmodHruW09XbbqK
vQ25LiTNQHb/Nclh3FpEbTYLoZCRB1CofNMLcTkCMwaDsnYq24LetuG9jx5N7zth
y4t9j7+rcgWUb4ItqViiTboR8Q3ES2K7R98kWiBy3+pQ2NelswMRs+/qV4tLSYTH
MNOFCmMaNL5wGsQdBX54MsCfhjNy9ygX1a6knorSSRtDmk9GQXCHr/+5IcrVUxyl
/WWPwzs37VD2baYXo0hNqJWPbzOGWpJvFrj5P5oqV6lk1m1FxrULSzLWfJbEwpV4
xWxOzcqwWY8eklG9Uhuqat/R30EaJlw6PwlrahL7V5lTCBMDFekPjutBOGANyFnC
3+HHJr0ybehkPPZF0/e1xD48Sp+dYLGbtMo6ylE1+ItsInqIX9hqN9/YZPDt6/5H
MHT/IqqeRj8mUKTYkerkahzB0lk8omOhh7eW98dK+U+DnvTV2q0dg4h5P+EirSth
xfSJV2G2cTE7sigMCbdRQP7IkUk5e0qSfChafUo46qEbe3uG+yaBWrmxNQfLhxel
W+ZC1s20+zbZW2YRLmtTUGDb3lOb2uwM8XqfpTjo2aCJq6TwFOA+7xyG39mGDCzy
3OwH+5qB6xodTnkycSkvyTD7Erhz0NrbK7m12ZZTbfGWRXEXwAHth+fK+KIPI5W7
x5UtESyCdrr77ZI2qjI6+dY+Nay9kPJDe3NEVljdOhpPsi32eMuVjmRx/UXgepuA
1n//XGFGYhFTiSYmO/Ls74C9GyJzt0nMshWyvEAAyWPxLPqejz0/WNvbcnyd3nlh
DkxTLxNy7Sh4+WjXotF9m+gRgXTtrpbbYNOA+TROTjkEqJIEQIIAcx4uNHHqUXGR
1R3ARHjuiJ4PGqi1n8MGQXK2CJrQkUw70Yk7EJm5n56nNQqNVgPIFonTmFc5hVPT
EpwDeF0gR+E+f96ZSzUibXy4R8NDoo1Afw1VWUhRirduZVRukZEmvebZZVH+JR7p
+xKc+Yvjp7oHeSlBVIyfiBzhLWAtEFt8nDz3KI5yhRqIEaEereOc92VFqcTE/wMB
Eltv4WfIajY4oNIMJvazv6i24P4aoZd2idoxxgzDnASuw+qhFbUUu2wVpDwZzPMU
yNnLpLQHcx2cWZqMWP7TqRE+hff8oKw3EUS4B1UCtKiTvcfuELQixxXk6iN2I0fS
RngJEJWPlkwqmNLZJYyyk0QRdD3x4dvgHZT1bJHRFOf2FOTA16kfzFxsurgwbz72
RfPiw62iO+NlnRLGg8QFwshaRvro3EjF3QmyaGDuxaearhZWb9pL8wrEl3RBPTyg
fdUFaqAt02axGzGMZSdVjfc2cdu7IMRBBjAjS2r+gRpb0MvMlMWAGj/8Evr22/p+
P3UlP7OoSI33HoyD3FZKpfJlJ6aVyoc7CurJjSPqvPYVOn97C2fngEDGfINXjz0n
zVoB9hwCRXQiEKDmFbL8L8RnOvAIV0bmkFPX2GjODxyVC8TgFOQ16+669pcQG2tn
isF4Xj1TnqTj/kew2IIdIUF1OrGSriJXEkI6RIa/Rwi7kWjSNrgmacSTZk/USzW/
mrn40vbzNTFNMsX3EFgD8seWGp66X9gBHkTy/E6lKuCHnTlWAgTQ52yCAoeU1GKC
Qr2V6hUiC6eLG3uXOtmhhi5QmRhaSdZt0kqvWKxYJgPXuvTZ/SV5Yp3ATSk7B0h9
3hryZwVvy82mrYGe87UqTB6BykpsHQTaXaxUO7W7TviwqITqWK0RlF+3f7wLmU8+
jE0Zp8qCmyjFkC6VV2M43JIY6Zgbp4RKysJAW2WmQrhm2CJ4deD3bhowZC6IG+mD
47hwnvjvAaBsYTBoThD4KQaoQjdJYf8Km+1f0B5ZBcqUA4SP8Hpisrl7l2pfZ8IL
XW3XAKE/RRpRaAslErLV6JNIFQLFgTckutyheKp2YPe1C9W16DzCIltpN9SfeWeq
Yi+7NTGcW952EX4PfE0zL8JjZ5k2fMH4vjORGtCBS283FZFs5YT280hhfT/+JlZ0
JSn/MhuFkRY67qf8r/+eDr0NawxUhLps8DQki8EF3VZoD3+ZniCurP1t3hkWdPN2
6khCOvqKXOo8u4+yhZQHN6Qxm1EnOOdCux+hEcxFwGENe1A0CnZgwwHqQE9Ew1Su
mcQkLTpd6UG37IrMGRCb12GAndkJBwD/XZq6pPvAYlik56jeKt0JE1Zo1Ej3oASV
sbc0TsDZFb0SrhL1NZSAKp5Akp3fGA41UoPiLqwiinTWHatQ9MTPLOqqT3KHNKpP
H4cmivpM6Ij5fhfh4gE4vF/ss06YCEhT5FRFfCUqecu2+P0UBqGNqtjKwmX9sgTB
LnPXApqMxlOSZRGGRwhtXNE4lHYF+b1NHUR01RKJd0r2cm11gdiYuoHY/FiEeQbT
lkl5ICASBBikijBll2N4657bmd9ptTF24fwBiSuHWYzpXjQwNq/AK0whq8rimkmi
McuzTjzNIfS0wcBEwHH3h9VysmQRP5wYyxhCz+tx+gZjqJHNGd5rLzXyySocxPN8
8uNX8rJOg5kannXpauV5Gra5JAiTub/JoVMijj594K+6DJZBQBs/G8WL72RUAvzU
PQGDlojEK4UbasiGXZun+N3zwOFzzlVQUKP8mZXAY6kXkTN9Q3CeWNNLQ0GGSkYi
bcmX0k2sLL5IkkMUtEAl7kDcZxE5CSRKMG+OyZ5AgVNt5WoR+6uuUhHTmlptc7iw
IzieBK7CDC3/Ie2tc9KauaXWLJ3Lcr81oVmKZB6T7cQXPesQUveg7T8ehf5wGSaY
fQXLJS5wpKyvN/eI1EAtFgH5leWCbMRPLdkXAqhPj5j7YyIRS0D93Uxae7/U9UMz
9mmDeiBRW7bsCzBPxm7hueP4GNFDopTCttXwxnbaZAKytNTguFEk3uRARw4GHjIq
DIkoRQomO1g9nc+LMN7j5C1Pe6qKFKuaR1TMnp714OHtl3ZTxtJ5v3N2KstnpOdB
zSWPPbmO8Bj0nf6QBkOyZQIa67aYXY/oq1YEHMzrW/l8yD4DsLCu40OTdbpEAKeu
LT5HbU0Z7UGf/m5weNR2BVWvfdVLPdGxTH9GiDUQKm96RMENtfCBLLc0dRN5vp7J
8u9km7lOm4TVJh+CreqEwGZCas0s81mqekim97UVwwXlPU5fvIC7s6rL4EKGqmRD
37WMMdfE75wK4wrR1Pj3SdlWRxLYGDtTuKoskJfxU87G5CPKrF+GISEXcf2MYsgW
wi4ME03MOwBKP/hza3gxx60/q1NYN46W+Nz8PQj1VSrej1PNrTsw5FAQU6a05rvA
a83irZk7ITv56Mwi0ssEUQsnMvzkK1dq0WWesXu5Rge2nxXwjt3AXEmLdE2xeim4
v60X5OEXUXqMw238Zbj/h0IyMHY3bi5+7sjIzXAvdMxU6LxhR9U4FgwuwiJ8ffoU
VFLmItY2RKo4Tg0EE6PuZPG8FgdjN1sEsQ/4qq4eyOuljqC607emm62rV8cPYUxq
NFSVTLH2PMn+bcb/081QzC/jhzpiGm2+wRRh2dk86t04FPHedIvtaqPNqPq0QZed
YCDzGtns2koMwCG1AsGoZ/+uzNRZj57XNaLjrf75hlHUeU+qpiSKk5fx3A7+eaMz
l8fzBswQrJkvWnMTuxUnVfyaLuuu6sYyY4JWc7RIW7utb0UABrbjtkkxdXWc3FRL
8O3qfXZD8dKhxFlmIB7MDhBs17X053CvRadOxwfD2nuB1e9psRf1OYo+Du0yboEA
AzslQqKguEfqmnpSYqnVA2schPPuYEfGmR+plRKeDszV+MFel8INCz7Maiweg7xf
pz+8FDO1w1gRtyxy+kwZMlTW59craHMsYsBpnah1nCXD9zS2i3mRvHHKixKhqSPq
U6uvr3XmfNZScNoT7Xv3gy9ZUD7lLc3gzrqIn2LgN+Hz3Ds/Kw+iWWlsBplMyfbx
A6ArmXe+TVJ71bbQV1nJr6hsAfZhsfgOSdvTQIfOMPlQHJtC3URyeqrFlnM5ejI1
WbuUzSFo6fcea6zWHTSzxcYhbgdsqQ4GZlqIVcaygN/PYs8W32Ykwt8c3xXN7t92
CnSJZizBbByEd9gx+f0tIzkzsy7/cC3XeEtwK5ehtkPFxuS0NHOloqOgcCWKaNHk
4sVUtEe2AsmC4um3EUIrePMpEyNTRHi284EKzaC0jkJuXmh9wfmVG5Ww/dICJuzF
JiqdA2FZkV2PZWAsPwQkmFyfl8RQ6QHRQMlUm+ScorN4tmK1RA/2EIr/4unEkQnn
8I/ORzA58Tsh9he7sG6I1ITRg2fMImn8xsnRwrPaZ/nvhyDrMWzbWW1SLCEeGAqO
aJxI1xxfERVEHPU/pSH89043d+zm+3+hc4CqQokwNrXxOO8dpzShLudWwYZ8mLOi
VUM/A9q7TliOEyaU6xQzgNoD8A7vPC+5z9DjUqgiGHSTi0oqLrASSUUlZcQ3qz2/
WdyNetb/GovMdNM3IiqC1Mfw6SGPh1CoFX8LKg6B9ab5XHR3m6ZlDNdbEQqETInp
b7IuGRUjy1beA8FJbmLgHXN43NfoX3Ll7uFTwcPeVdXGRhjoES+RaC+0AD26vOm2
lPPVLvp5Xl2sovFZrU8nSvxnaeecShdFaetIrfSz9F66c3LMJCUmHwGN95Zz+aL+
G/OJrgDvDUNwACeH9dEy6yXUUnUMirm146aM6JHr85V19yk3dsXQXP07aqkeB/IT
6ioia7nDVOlv6BUJSFlYNGZCuh7Ch1fHFpdbCxFQ2t4amyJMmij5Nfro8LX705ni
hd4F8mx9LBb4hoDEo621VsX+hy3G5zES7AYB46WMQdYfIfXwgbFn1nZsAAjw77PO
I5wleUt9GyuQlbMo+hn7km3Xq/7rTUFMLhyG226r0zQtjkP0v0CZWNiRb7cxiazB
inaogHy6QvQP95+yQNzhipB/rZPHvYVa1xVthqZeIDD+0WN6kcV3MWoRttoxdHs4
Ln+hYNr/SoVYaR80X8wtDxp7BxR0vInYNaAr4Gnm3mRirSt6/NDXx3yOgwx7hVrq
TpgICVqBp5zgsGJW8Oa3IN8VvMQuQjEb4CrqdhoKnCgitHKp/V7Y96pATYFesoMy
CV4zdJDU5dj3NE91QfCFHPJ3sjyS7uW5WtguNvK3v2evSpR7Ox6mcZnU4hG1z3ce
nPYTps7mMzIJeagB1+i8wdPWQyVgBWm2L7vn7HDE/5MYScDI28YrqUnBIH+Tt5Dc
ENr2zJcnH4okoY8yYO8qmF6MGs2Q9jsqlqEWJeqovFFFbZZWVJdu3arxGM9HM6aH
5RJC2MbRpiu2/TKxlGmsWdE9Mc/XDhmX5DPmGjsmw99xPxjZrzXm70252SYZreSd
g+xmRvyWM+N9RDtK9Hw8Xw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Vl4fHut4yYEbCUoRSGeWlxSaIbqGITd/K6W2sIiXDHoiWQtVvLTZfLVLHXQitdC6
8vQlLfVt3MYLWrgahLjJsgOBbVvowxcPWss8j85Xez+IOU77vSmdTWvxW2U5uiN+
uZZE0JyYDruuKxMC22TV/VHO7XPxwpgYXPiANbC36KSoabmKBH2TsKTzjeOKq8bv
xn4H6iyBVN/IQe7KcHruOXfdkIzTbWFLfmSSiZD4l2NYjAOARyiLa28kpih7g2ds
DoFVCCPjaEOhMIp/YK8mzzTW/O09OMS/3UyzCOsL7fJavKpb+mgX54JsqHA3/DRU
tYe6hLE+elmKiqHCwl/o5A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10640 )
`pragma protect data_block
BKZDVvFV8a9vM9sGUB63bqhfjl4xXl/sch/c87ZB3gHuME5O4RqxyeV9a9BVHETf
589wbGZIS4vXZouE7ZSCwiVr1ss7oCiJWY8qLBjX/ks1WH/C9dgIl0XQFd6OHvY5
pFeJ6zmfYOa0SguH53GCTwnpinSycCrwXgRZokXcZVHPNbumszio7Z1hn4z56RZx
0Gu6U4XnIyQXnI+YFOroxGRT+B5dMhJjohAgE257WNARGgjAl3YWqXyASZwl2xUB
IDYuy/ydbufGOnnwVOIVhFrah7A2DPptbcNPMOSph2QTivHkD8x1jwP0Y6S9MK1L
xGfUEmPRFgVEjbNCBDqURMlTi8unuME8QrWjOOFi6v0WC9xxpwTVjHq5L4Tj3pEr
tUrNqTrJwQnVLMXTCfouKFQAJaza275wp0k0iVgOh4yHzNGKLo8yMB+wFbRCaMzH
SePBcbaaHd1oIQEBfVLlL47P7HFzZWLGTkfi9iAMo+5pRdY9enL/qV72W3JpAwXV
lqhVZ6rgRdwAv1Gt9s9Hz+4EG+MmyMpJ3lseIsuvAFTOCPxwLBue7cSjoOyIgZ4n
Zb0RjFJqJiQkBBSLNXkupuOkp1iHbfLisiKCwknsX0Lyj1n5fwpkmRPAflorGQkT
2L3rTV+7OAeOVaxKphEHqfQ7qFMgauEnRPB2rNrl1heLfMnuz8aze4yUAebAn2Yy
jmwWOtmieym5ZXt5BDaoADrQtY2HL6I8havgKGZ69w0Cl6TM7SMtPLIF2geOBsj5
jCYhIJNO7bsaSEDvxQ2K6ea8F1RlUuCGkIh/0p/DkfmF+zq15EbwqgdWmPwmhaO2
9vd2n+vItP1UOwDFtfR9V/POa4v8oODuJlM2qDWLySOOK8WmXVknK9qjn7AaIKr9
4ss4QJnkSgam0o9v9QWn4ARMTiJ/z7HHKG8MPcPhl/qcoBctP51acndOexCqvVhP
9i1TdF7udQJ0dlo5UliPcLLt0QDpfuehgKES23legkBEq3vJ/LS4JgaQjNQKo6lF
0VCNE+wErr+tVMojsWFd039zcRgXtSHLt0LTQjiV0xNTOk4kYwBgDseB8mhfOyK8
J70N5bvV4IrjMKE1CzXHFQT1PD9tn+HDlnGBMcAZ8lswIRFazCOkjMLpMYric5QB
UOpCqOSzQfvtB20BS4PhMnZM1P7S9POUDPkG0XTP56jjbI7WmKlFJASzjPaFyIwS
cSfXuiZWne1kRrsdCVIkOLoReEHJIVGeN/ddhFyJ5zzUXih6vOyuV9Wv/8tXsSGl
ercNg+fD48K0Chs3Vl8UqM/NaFGz5CXhED99pYisOPTW2r2m93SuX2G/H+GaJKQW
uTAUWB4NmOUqrKTDsxRjGpmhi2UMAnj4KDAMGVpYCV5w93TfST8f6wJfSgHyMNyh
DEcNEb5vEM+FDc3r6YP/ik6ncatde2qedbcI+KzpO85fd4Ri0ozITNw1eKDmXbau
8tiRn6pKwef+IcC2sZFsjLZDbF8i3wnECIRETDn4s0Pofa7ITLW2VG2IIiOERVvL
ddZbhXXVlrBYcmgzPTDU5Ew0HEHSwKgzD5A9Qy8ZEH/56YImW7VNza4evdiln8z7
wNvJBaazkVbD5ICWiEEW+efb6QMrdDUgYnviDckwv++XkeK8KSd1AjXIfxcpMPuu
mSc4ishBPA7RnXeEiJkaHp8poj6WTbGlA4p3QuoJlsQzNqgngaceY2mPbhHqonM9
cNxaGDeZxw+QsLz+PVkOI0tM78FSl/jnVnueaRcK0s8svl7S/erovOUQ8e5oHfad
H/ExHqiqFUrXrnqQJ1yDyocIMMuGFpajH3DUiz/yHdQT8IW4oxNH67Vma6fKXWA1
vRm9FTI42g2BfCUIMWF/PT3ZjeV+i4avO5Ae9McuceDl9GEcr6V3X2ere8nmV1IL
yEV6T/l6ioLrA7FtimNQYQijSZ1FegYXjFLTPXGiIx35tcO/q2M6q6mEvPz6QDSF
7ynurniPuM3zPGgccZ9897niHveUgPk3ku1FuUQZz6XgFfvwoxwgFwDBcJiSmMn1
Cv5MfVzxaXhE1ydAw3AhNSGAmk789hLJrisStFwYKVCnlKy7HhliPW3nNFyZc41r
7P9aP1dpXqyo7QqVNMtbbw8rwwtT/f9LEYD+7Wm4HSLk9gKyPKu3252RJ/wwMfar
xz9KDCVD1m3ymHoswZ0cAmM1y8GfXGs2jXch4gwQ3EWFRNpDzkNUTSZfQ5zLaJgb
i0m+bnUX4aHAN3to7mAuGSgwmAZjObcpu+zoQC0NyhgAs+H5GFtIOHk9JvkfqwVK
YMjDUG/yIcCW0awpoJXhmUqzH3ApXR+1cWJe2FHpvsmaV5l/eGJyHy2GrAq6H+Ym
CdSxhBFdO6goPHNYeOq7iMPblKX+wjQz448IrTE7wuJhZTA0rNvtiaOnykYA+tL5
Od9C13y7tQBPdnNXdKtuwSoU7vtFVm/i2XC1kKherokudI2IrCWYuvvUvy+sWSPK
Sefe+EUtKND8bchfMHuFlTQenydgWW+aeg4ngAJlf4YUFEVkP0mpNfgWC1l+Gi9A
XZ/oZ1KiwAycpbdLeQVsgNJPsskEiTTWsnkJz+c0Wtpp5QJfVSPyrpd0rMJMvPRY
r4qDbifQEntLZMLiSBMyE1D40SoJsdUtBpIhD7679lLqSMB1UhG2rKeV6DI6xWGe
xGpFPoaMH7HNdpjr6dOoPPmwF5mTX0FYM77T454lVg+rEZS5cBqMX4sFLmtfWURI
UqsdOnDNNrm+NTYJ12hUlIQLSngoe/CQlUOOJ2ajgmBWuGEsAJXqG7E2IJciBNoZ
qvj3UzACMZxPMvWAFzSb2seXwsgBy/oTMkI4pAzoKKe/3f2b1XS4079hj8wdZTnx
rmJgD4afL7ATEHZw42H11i9KNiErDQ+bCnvSys/2NY4f4CBEybq2Eh8ikja7vzuM
57o3cymf7KWVGZ8f7aCLbOtGkSanmkdmqa42lwgxmich5HY/i9U7mtK0ewdOmXnO
GaURbSNonJ+HDcodgI9KsSKNWHa/gTeddh8YYPZ8W1gJVeDUgdRNwom0beITj/yG
v0kIPrtumILsnWSs6NIocJaM/A/Lf9dSKhqidyxJKypeLj638cN6ev2mgcaxTuXi
v2szOL4B31yg1qL9nK4pPVL6YVCcGzZIDKiwcYOeotrS2AWtWdtVfFW+2kl/Q6U1
8umdWdnshF1ppiAnnoRSHcS1din4XJWzy3mxEsxLNzla4cO69tX079GTmo0E1Pvb
AjaOlqldHzl4EYHX+VCuLq1peWxoctSjT1ayZ4IqL0SFsv/dtDoqB+FJXdxecPvQ
Sr4uiJfGe3ImQg6P8KuD78UxdAOT3ulPj8cEIE3Qp6pEj5hpWK1LZvbAlJXmgA2C
YQf+f4w85WEprCvHH1i/p4qUBMT0CyrQJA4H4ceHIcSp4Nn9+nkP2xheR76B3XB6
aeYbDzraUIBPbNBW7aHl0J6EwmUdg8olrvbP8IIZ65iAFPp0/HoqzmXPQSotYfnv
AfuIBgRrvpBfNmeauH6X58ZYWWFCRIT4/AZWk37FvCjA5slTapiLENtVm3qaDmP+
2mNo9p/7O4FfvGu9VugfkB28+A46rlsWJl4GAD0TkZcqqcT4Ghsro6Zbv4fhVUEp
wYMDS1jSFJ2Qz2xZY7z46GqDLKqfoLPud2BeDkQnIrmwAR/AtQkRckt7vKitMSyP
7NRCGzC2QVT0g7c+OBvLOnVt+nyZK0JmaHiaeyqa2bODfBi8mpQR9RPyrya25Lw4
rIa5KE+6Xs6NudEpuLQ8AI3IzetBjtVsl2RgPQPBX5kuG6S7HDLXODeUmxipd3Ml
ooJXjPi0k1WTnnh6Y1KXfDcJ6F5eu/8H9Us+gd0OYfopBDtxuSm6Vy6NG0KKLp0E
+Jpuxbcpj/n489ApMTtKVUJkZV6Yr8FDf8U8NRGn8yv46uhdkUF5Wm6prXkQvqqn
uXQBhS/YaBTDy+fyaFNlYKZ637P1TwCH4m9NiogfqyMxjApnqi8/VOA2mOuIBgTE
kfF+WmhVHK/3oLMrkltEF6UdlsehYN5jST6AL2HBefgkkxtQWtagxDZWMjvRV8WL
1FJC9dubfG7s1y961ICqeNb6nYfssPlqX6Z38P8PXgw3JO2MJPrXr9Ghwz6Dvlzf
ylyG/qGxZ2ANjPhEThMlSmvSQ3Yl3MG5rFfjYdV4NPTHKOY2U6I8MLTaSb81sPrd
LJANRxY6KtJ/Ma5olDSiUmm9mMWqlhdwJpaBbt/ISFPz18katLnKZAh17zk8wCUK
evS/cSrtYCYZWmUecinqkCyebx8M5bQej1S+U1Wq+3tq8x7NSnqDjt9McwRhV3Xd
/lZAp0SmhRvaQrCS4iALPKYlqDLIxNgLSZV71kacnyOnCPJBpFQojwqjR3xQb4lj
5j/zrudk7Zu8Q9YlLLY0OH09HPfT9aQ8+Rwki66qabxj3BgxkuVwEw4nHgizxair
XytLowBbbPirqviodCx1cLqiDZgfCCkVv9RX9P4jgfEjGHDFtbCOchWludZhQP0f
Q4yIWpfTRPgbPlTuPp2lzUIT7BkOuNWXUk5b2zuC9jVhvyYu1zo1p6LWFjwNq/el
ebcL2G8maWEO8Ad9/O84RrN8ngDmbwRDK7CJmCrW7msthOyfMv2y/zDg5fzzo2vJ
byj61YcFCVm4AmrXXjkz99DAL91pQq5qR2uy8x+YISZWdqCh5MgHmGKvJp19x2BF
roVGlIJNMI0rAVYnqQTLYvomUZxJ54VaTU0gbfJc65suoytaqSozEXK1vJPGchPh
3MUEkA2MeRwNuwcCJiPaVwXRO3rh/jkAPvtUsXirtkkMmB2lZd6oIVkxAphrfoNw
BWNTDYAZTrBF2WDass1uMKhAqdGU1khyK/LPSfQFMz7XG7sRhsGCU9lCM1nko7rN
R4ATX0kcrTABdFatqAZMVASh14P7MHoYUiRzDckaxi11015b0GoOn1+4R6PWFa+s
gfJaaupOpBK53b+Klspos/5bKQhU6nu0kMXTnuROl35ZM7z75rkm+PT/I0OuERp0
O59Cv6t9xDzESeOgrgPiDypC0y/xNXRt3ZweQ+wkMuutskDfU+PsupWexs0/SD3C
iVmKTd8RySrEEpCaQsTmfgyN5cM4pDV+/nxQWKmDjdU2QUTbiFxU7ICJPL91OKc9
WBG2gEkzcuem9h647R2ODOQQoqV3OOzRVL8vzw6q2GWN+WXZSNHxwHikfTCV/P7r
/hz5VPoc9RTrrCV8z8MNCG7/To/ZOKC8kBWOq0BxMiVNYdHXEM/qT20fGB0fA+Vs
CF6FGXhM8V3kJpnJ9K9RCWFpuHNRCT4LVmH+sH9M25p5jybm9hzg2bAj9KSHikHV
89zSYzWNK1C05dNFfVOhF3s+U6hMAWLemKvGHciiq3qBFXNquJiMd/ndabfB7FH7
j+C5Y4YRNea/Bcd/kSj4jl7Ma4TGdqpQZ1yDOtBp8xXVZyjppKiP71Bj/UrqqnqY
hFa25g46utID3WmKBV/si5S5a/9hv7EuQva0LQyb0/KBEtFRQrNpv8x+I7qOZSrW
bxZL2Dx3rBrX2tkNo7C+WzfNPdUMefrThWWi9gGhSdQU8nQGIPLhFSQ/hvgBBWIV
0XYO22ix5jV+Rrx2BrLWeum9P+F1YCOS83nQ7AnLGwct5adg1OhoZfK3bS4GxVze
DvGhbDMz+HW1OWPyXfuOhwEOVRxibDpijqTNr4iL1UFSCp7mblDlgmVfMZroj+v6
0WiuQBkaYpCaOHThZmWzNH4vg4mgwIjJok1gF6pAaH6tPL7lcxU0cY//ihfDP1YM
WO3dTtZnjaZlFIi4Txt8hy0T6ppV/WSz8earF9XGd2RHwwE3jNCBQNokF7vEVxxx
87TSqsQEjSH3Ur71k7e8uvKiYkjOtJyARdtecG/qqcOWEjYXWILfggKMKAgkqANw
kdkTJWCpzSzTfXi2Ce+wpHDW4dmnrtnrFWwfUtyKDBRY3iUwdnqwu3OmKgSE11n8
tGPk10oY+RDAUGZekGLZBoPX/D2X6S1AMDQRONeEvffRpajxMuvzadFwmqRgK5FK
5wE/DnW6zIPP4FRXY2T/5T28DPAEpuVcVTsgdFlor+rl4cZj2FwB03NdjwQ23sQe
CGhs40l3jPhnwVul/zP77b9FpXvyg1kteWCjzujNvD81yywojsYOAgAIawzMgJxJ
QhE2OE7PHVC/Vywwp99Ku2nKDyp5cEbcU3YV9EiWl1qLCCOll9Wzqaga+us2JGBu
hKary/wAvpCp99WCgi28q1KzgWr3qgYNR8Vs5SIs37lrDeIX3rWd8EitYTTt9zfs
pbDOdK/PH0D8h1HHfQWpr3xatsFTDN0221UkHbYI+GPf4tmcvBjlQ/pzaLuIOcfu
n78tlN4Iobdxi2FBpbX/c4CfZxN2HHla31FWz0C7FwtIvn1T2CgKn3Ta5mR9lbx6
fRJpsCF9jqu+v9BL0hMOQkB/FUHIGtF+6pBV5m8mzlQuTBmHTCrKIeRbybPaBS6+
1V9/vdWKBPYlSkpbscxeZH3gryAHsaaW1IliNgD8m7AZlc/UMBTHaz1xt+3wrxoS
Vyuu5uozbYbgKDt1oQh78ZyiXPcjcEKawtsdyGCa8dHYCKIk97IRWIvE1zDL8Y0T
08QCIWvvIOP1fKuuVj97171WRngqaAF3wQ5kLZnt9C28UVzxnGeatpt454ashyx1
KrODDgdNpQGxdW0ddLnE2eCv45oODz4czetGw05uaYQoV/TgETE4IgIJA02rYq13
msButlyBr9fy8MTG2Rz4O1S9jatdZ1puunFe4Ot1+lG93kvgzCTk7CPuaBYzfRBG
N81POTqE+yzS9ZIyV0bYQsID0+8MWFi1I6a0D+1ZeUJ/fzuGcWf9JJvP64VFTNVL
MkOmQ/oSyEp/JyTZwtgffUMl7ynFwIkXuSBFsaPVMsv/i16PjnJT4w1PRpN6pzxb
Qz3QDOHXYhltkFcgzPuEKBMfEdhlK5Vzrb8ATardIGGAWeEAnXosjRKwlwnZGNR2
JPSMfMyoTL+spvIgG+miJqOd0bIqhqUrR9Ux0zh8W6REjp89nbuUFdVAbCdevoyO
qDqtW+SH9syjIinHuQ/mQ3hoJNMarzNC2rwRIvV4XgIn9M0jtX/kwr93o+UFDZu4
o5NfegnoRd2gYWnVqpiNd7Ig/N5Wz5b1GCJTRk1yIZoehDb5GW42VslS65SIgaNa
wlDfCf/E0NF+EWrd2LtKQ0miPn8GjyWJ0V43SLBJx5adrhDJoUl3NRkEXrXV/dMe
Lt3GTSV8ZRpY7SszjzPZhmQvGkcC4708hyFt8fscfetQyFjeBx/O9ltxg1QmN/o4
PIp3Br3JKMmBO8dWz6uOTGkBA9Bm1hBVaHWMtyJ2YpKQeG7QArtfBrRkRZFvuYAN
NZku0RkbLOGPr8kmpaLxKXCQAGrFGgv+KKpciWJhMnEbMqcszmlFwScwZ8bJtdIm
t81azMI6PG4bs1qouKr6b5KpHZP6Esymy3EwwJYgVIJZLyqVDAhw7tnwf31eOgtv
CXRyHoQw4RkykFqSXkISA7PkMEB7noivyHm559lJHu8swO432HIMQ0dgfVuqZb0c
DqT67sEeOCw7KnbDcFv5+J+vUwm/Ne8H9UHVTDdgXJ4UBcb4QuIXApP4MXVmYNsO
3GnjYxUXUIRuU9HG6IeNbEhJfHcrpOMFtz31Br4nIdTYWzvhxGYjIArdIwMIMspq
kMU8caizOcyxFPxkLmpkei4EX5frnEfTRREPqjZ4bIzntlCZ+/6luLKPK81LJYo8
c4OGHkG6ZE9aHg/ejZKksLNB/O1lmU1GI2pcRlRHydbZb7WSbpfoP8q+pwVCga6S
PYGvw67lrIjdbrMpNtAhp2z4hWIrmSttTYp73POgmaaB9+LGh6JxRXA+0ZAOx7Mi
+C5SaIGveFOJINk8h4EL7lEbEKqy35pKOqN3IaRdG3+9dj/d+DRJIRvcPLQcJjpk
xrnB4ZrTdTUqH74UI+VIHuMMWPudVWyNlfcWuQEEWaQix/2+qrQiGU6qSK/KdJgY
SRkA8NyjFlt9WyCRGkes2g4sb2YgSdCQYMrjf0HWirHSt9k6qfMBkNHhEKCqZfZn
4r1XjULQEp5Ob2pW21NQTWktR3P9wCscyATDTCDGHiF2jkgCpPsuKpdBmAzqFnEA
Nlt7WXi4mS8yYDdyvh62I030BohANEwOw6sEOVRWF01pki/0mGCofYYdl/pmUnit
051EklcWR5kxN4CggKfkv6AP4f6mhbVNWl6ue+8mfjqp4ORuKc2U9aW13avyi4fr
AQ4aN7rB07+8Xcr3K9MDoZ6YMCIOUnO7iA17nDdE0sRFzQea14A7E6xUoewrGB0f
QyH48cFHnaL432G9rgefm9QS97BldtmILohl7FtdQLT7/HJWdTQOj30UanM/MYz6
34mGv9UNC0lpBjdrJsMvHn45sH6voZnPU6SPmzJKvn1Xxmt0EMH8tbOtr7yoFWE7
gQX4i7yU28nlpsvB3bVRJkjdLGEd15oVE20eUa1n2ievm6TDdXIqS8Xtabro/K/K
eXGQyQrlyyIFwGl5iXfU+iK/mSsgA13GZHqe5G2xrxgIW4Jl9PePW9dPEDMyJH/L
MGkftNMW17dx8a9STnxKm4uoQAulHAzG0JBpZAXHqel3UjAMdz4pTUJ6Yk7fXfNR
cTFL53pEpw1B9Nnvu0S7WAToCneFJdG0lQLyg5mrNzv3voIT1nFaqagaOKEHORez
5Vsz0ihFnueNymlAYL7ISPijon8O/iUoSr6h+Sf0WNkdYoUVoidznDOzDpPoATcn
3ZOO33w9+IYI5UEe7wGVMn1BcblheKuvC3mRGpKZasxXrUv1DUffPS7EvU+TpShf
sWW67tk9oXT28fLl1RmuASICBeYPQnjN/BALVhQ60KmNAK3pKNsRP2ZzEF390U/R
Ax4h2a4j8AJ0FYkRTEV22opxmJKvQ1GqNjAkSVPsWPavS3RMD2TUKDcHjcCa0/FQ
wzP5hDNEtgD9ySgZVn2u8GP5DzWxgYAsl59lUqYX0XUaHH+XPv0cixaZTfX329wU
13jMcWj8sLItMa8NebNyxHfqCdEbOApVyHDRTCQ0RLOWw4Bfc2BfvSpNAgIXlPz1
b2seq6ALrxEsSyCnCuI08F+W4xUyW6cOZggg249KtA4DNh1wRHVNFhvFL3um/oaW
I3YsRxJy+YkEiLUyfQN2la/dazHzgn0kwM6I/PR8wDZsz/3N2DE1vGwQIBcQYwr6
8pVvHaAwKa5F5uSxdRMDCN+f6LPs16FCvRnCdIpAqbNtz5uhx/9Eo8rmqko7cD46
ya8jSlIFmI/YDssL0db15xiFrJXpIYbm6Yxfe/NRmgP6lN/gaSy2CfeMhJ9cvEO8
Grr8+WlBncBMNdjp54TRBFWTZibN4XJNF7yz313ojxhmo6eWfqP4vgX43Fn6Vup3
godpMBYiqwGoGJEOKhhzST60WgEXnHMcQWT4QFW22AE8e+uPsqnN46uDVh3Bc1f2
odln7vUNASn4vS25Rgipwn2JK0UKKoVHO3p/L0QZJIiwD2L92E42F1ItqUNn51CT
GKl0bU+oJscbH9OQ2KJk6HyCtNpCBqqgErItNFCLHSUY8YAfmvNoxyAGMtVPeyZj
BXjFISb1sugHyd25Fuq6O9FalDus82HBgzVUVpgB9q7qDn3Z+PcUc7lY24WYOpdo
ISzoU25spmfh7HqrqUvftwT6otQ68tMIiwMDW6ZQcuextIj4ltI4/IVpxqDzdb7t
B4rIF34k6hexNpk1hDuluCN2UaT/KpMPs85zZGBPzkiml8OLOX6oyIMuxtWFvFds
ZRYzKdRsFDyaVeEmVUqh2RNG5BACsGVnxxBneVgJeavn5YJvsEVo+VzLsvK7brmF
ZoWevuN69V0WV3gwINRqEhyMizGfOBB2XCEQ12OoaJpDXzPxwTisN8Lev7XiPam+
BduY/seW5/beuuos/VXXg3maxdailjZhgibEr1nZLYenpm04tTNZvVgZhToED3HI
Tgs7ioBvfKQDWQGpU7fH8RParvnt8LHKbt78fMb8yXHTFltbmkbj8uXS1e6Z8V7D
ZW1mBRQbvhDUyCF8W/QYr+UEbB0q2Qomk/AzJhgA4J4UP76aZKajk3CBqbUEvsSl
nBKj4ZHHV2MHR+kk0aa+Wh5mUhEckSsFgmxH2soyrL38hdCjlE1FlBTN+ht5w/0k
pW3DD09p2Iw14qx/hicAdMo1IekEefmyEV/e2aQf6lkWUIm9SOj06ubrG5WKufDJ
OmsbeyVWPgpFz5vj/L7OfpyPAG42UQQv72tRKKBseMAZQt5vzI4Iu8Sts3rv512P
j0fyeDL5taZuQZyzOPZkM2p7fswbkI767Kge570wVzhOxh9NWuXaDkckJHPk4Pyx
hpvDYnvS1xwVds3Szf9E6/+Al0En9zcaAJTEVWR3F8zDTh9RCw/zl1623VjoyIcZ
6vJvSbCJ+j/KptKqZf5OhbdoKtIqxO0pb6R9yN/vX3AB045Tk7HhsysPOD2c5SQE
DiiT7r7A1v9NStacrZFiTNeNOVWRyNY0lDhvdsbx6ZkeRSriuz7E4rusXUnLuFQs
9ptT9n60GR9eJS9DtJyawr8UwafvgrzRQFiSu4RaceAh/DI6SSRnFs/lqoFWFplQ
bvAql1h/ioye2oBiSiC8sKja+uWjbfXyUUrudyz9KEUcMWafzzDCtlrhXbesE4KM
vTtWDsTPtxG91mKPSpU/W35JgESlOC99Lzc86oOisU74ztcmQhfzNwZTp6ZtBr8Y
aM5JnxRzrYKB5P22C7I51J8PgLDg5ySIYPa65Ip5eBhCS58L1KOV3bnjdhteZQzL
y0fZoUSrAYFxEzPN/CY2whJmc/1UmodmhCKpFEPrwzhZX8lSBDPhs3GmzHugWwiL
aXRGSzwHq/F72wk7LLxqdQFSLR/LeI9Lfd8NOLMtvfmvv/Nzxxx7IASjI37sRvfz
m1O7M0JiVpnjoTVsSu5HVioXrn4VsPVT8iGYqXJeiL14tMr48Q//Hcfw21ftwdtO
0mUqE7DwMVOVX5PieHYlv9NGoX9nQORCGrLjfS16+GZFgGQm9hu0oovGO9pxi5FA
YkoC7ie7tasbvVIBrGCbo+YSdEPZ/KJz2GfRzdMJ3y50nFpvDuHb8bTLAj0orgSg
ay7VHDNTZQSjv25F+kaCsCZj7aVTaVht/IMI1d/DOvSRfNeNY2rZldJf6Gvdyd56
e20LubBhOdxUy9fkkP87abPzqnxLSWVJM8UIPi5KmdCss0fhFTqMyd02OvuZvIJA
N3+r80zJYTufo/QCPlN9d26x9ukRdcxwr0k/QBfo11PBMtdm9RiUwUS2M+w1y87A
Yv4z2BPbhht5YSsFz1k9omveGlZEOpjKww+znZ4M/EZOJzfSIprTJU+hpQyF4djp
+zkOLHfNvBOerf8Q0XF51TBgXDESrobxM76+g+LTmWOH7E2USWmBCn95xc+Z+0XK
+j9JLsZdrZTXpCqLhxfAzai9W/BG94/3WWpsDSnmTbY9CiLbk+FhIFu6i6O3O4Ks
cfvvOALvu4E5ArB/aeV6Rsyvb/XwmBcYGa8k5P2fkweZsxttHpJ9MynotRQaq1gQ
ndh4zVvtwLOPk4s9/Z4LZfDhVUTXhfye6sKleFRUyIIHRt00oUZcOlTWz3LDPfJR
F6xzr6qLSzaDRouCZV1lpiymKrobPqXcwxNZhkTu8txP4lAZy7WVdYu2ji/NA6Eo
U7f+7IcHXK9zUSh3r/734NvCqG7y1NScCCIBFMAn/qM983UXLe9yTpVnh8TW20SL
9F//u4ajXvibDnudOam/6uRPhl8xyl/1e6IoHZWcL6MHN15rAkapU+JnVt+z7FuC
x9j1XHCKkuhxTnh799rAX0hMt8w/CfR6IRKepDvCRrbWKMrr0CQ0ltOfgHSN2SlQ
Qdoz6HMW5ujDfYvbFiB8kwVNpAdXfJ0FhI6nfdSQXq1v7jm3vVEsKGteFY7aTBGA
ObWuFiTCtFALiYeTuOcEFOX1I2Uq/wnWV3yb6OpwRP+cEgVS8iVqRVz2eRRvOp5/
obmRGYDsaAYfJlAf81S9jngOg1e2c2Ei4hg3xtLAVPJ7Q3uObiUJpn3Iz8TNV4d4
hUH0W/YiFOMtO998zxrK3KCMvoeslnEcmY9knwQ+d6MBQjXmhL4/KaLELttrkolf
mENk0PQMiq7jwvLih+wJZkC13LXvCOHHyCHnjY2rpOUR/gNctbJZWWhjw/cSTNbp
ym/2Riy0hF5gIt8dVYXYbiGXR7f0eg4gBvLcYEsrmmAlTZwPVLlO2BD3wK3lMk0m
HKd4wz16Ap1vodUUwmm3F/dRv4Tn17sHBPMg6j++9BCvGJFN1GH9SDtw1BDz2IPJ
4xfk/hWygwauWNdVICJTGvQ8quVdA/umnphNVlG7KEDEPjsL1w1O8tHxvP3Muaf/
Vi+L8mK4aLXFNYU41NEeMsW8rSaGdh1pQ786W8VPR670NQ/7Fe1RseCaZAI9tOyp
s0EXgp321Jk5RxZPJhFmix3b1P9W0HR+MuZzpCZaGtryuu8iD0Spff7ppU/Sfb0o
ThbK9PbpFe4oBeP/AbMGlNO3H5nXkEZH03lRlCSJZUsPuj4uQLB/AraI1wnIAStd
sSs3h0+koeuY5S3p7B3C5RMZLNI0UR1IihSXDoYDCR4liiVjFdQtqapiMLlphN48
aFuubsQdzwPevlpt4tDGyi0fMFxQ3fjbDgL0QVYcIVg0n3+0Z241IOQq8QW3dNPb
Mb+o67Rh5jCwl/LR9NvQXpI0f0pnukPBQLO3qcZIou3c2UKS0BdVWaMLCH45PeoX
jVsUtlu/Wnf7vzAcj5ADoJXz27nxBA2gyyFl5CQyPhsj0KOPZL99AANZWQA2nzpb
Ba/Axtkmw4VM8f6PJRP+JUut+U4SNNPQ4Y6sGMZ477oeHhOl1g1jMPXuHVLPvevN
ANgjb+9qR/g8mxYbEBGNHkuulRGomwBP5rvtxsHUJ9nPbU+ePFDqUUDmsu3QDtXx
0Bzse2yhRnDMs7WpQd+f4Erj5VF43N/GL8Dxe3epxYG8Kjnj2HE8nCmdoZuUxOX2
O0s7AbweVBn/SH4Ft2+iIqJ0jReh2XXJRPrdsVXhiu96HHtemgETj09x9zYZif8a
ULlrM9Z/SgHPVQBFuWd1t58E+W1csyQHq0TfSQCjJYRtGm3ecZtu8+JoOXxfn5qq
2ox+0dHmLfW2FO9BvTIzW0U0H5wYqqu3wFeWQDuPaVfWgxPA57DHqO68aOjaTW+a
FIN6VUGSR/oTF7FyVuqWzoJQiaWy1EZ6nkGEq+bDHERgfnTbsK9j9JuBh7TCqjgT
9HR0BjOOw1IYTDTDfAWxcRrfzYzFbRNE2a8bX5svsBIYKU5DdMns+utGuCU+PVS3
BJusyrF8+ajrWXEPUenppeXd6HJAs82qwdy5YsR9W/eUZAGsoo20cUH7KQkMo8mH
Y1G0z/hUpdBFoFTnNAT7HLVRHOf99xBQI4J9VBV307d4RVdbMYZwdRnhQU0atxKH
NHEKzaSHP4HyCjyxRId22So7fnWE+8JqkDx52+y/9jO1Bc5ebZ/fuFXk/y7g+Aic
/Mzd5wjNtSr/IHrcTxRo8ZnTxKxZWsG908sPtMmGhBCs14RepgxF5X0gvkWUjTKp
fncjdRoS3/4IEcy8VWA9S0MZ2U7Sb/xshnL7Rwqy9q5B31ptngy+drjKbajbDzUJ
lueQ87PR3/sMV69z9+GG10rGb8tzv0B49y3UiyLxT2XqTbO1Cytvj/qgHl2C42t3
blRvq9EIXlrWycyZSrjqAhN6tEvWA/pw7mfPODO+oAMK5+E4VzsXhPTetxvhWxos
NGZQpGnf2ia9BdTKJd5OZYe1aDBtOtZnVHsR8Ws2NO2iNjeOxGiO+T5Wb7Hwp5b1
zoiiR91UMOmfYIr165B9RrttcQmtf8+TI+hQVMJrd5d5LkDbEKaSMSUlY9H8EdZK
uy+Ccp14FbBPftHRw0NlKny4j6dKBxOP+gniyKrXpAEerQhrZxvehWbMldOy2pTO
t+S/NP16UX/nMsrPRyA2afAsov0UOU7AmwYUjlCpBBY7lEsHDBXk93Zl4Hdke9cw
F7NQyODpiDsGGBARq/NFCGby0UTsVDzG/HHdC1UnCWs=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cdfvj5SbLXTQLlq7mn0nV+T2QHJpE/G+qUpb+N/I568zqLwU+HFLXjYHgs7k1dsj
RicHhTPujYj3bwi/8GJQKCMdtlcStsEBBoOjLiXEIjej8HgJsDSJHoTwA0DbqrbC
07IaSZ4sZHRq1rO7fpvf5gvphI5+tg5unEf+nvM/P6x92YjakarkbdvidVDNTNn3
LpYL8V+PLOwHT3Q91V2S5QH1IA6eD+1N9tTCesIBLxg1Ssp/nZTlZW4X8cZue7e0
U4u+RumwdZPsm/Lx+3qD2liiq0iMvO30S2YDBqtZKHxzrC0us0xopY9iS7z8yZAp
9Y1yfOH07n8aEY1zSp5cjA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2704 )
`pragma protect data_block
xPy4sk5ty3RicS9O5p0psc5xRZbcSSTQ7Uf1f8Wnapun/F3/ZEb9dxj68S1Kp0cM
UxYNxT4omUwwQ6rqCRlKs6LBVzCQZynBl51YrZd6cAUM+8f1CCnQO8dRaWRp9vJK
Smi6URsXJkgu9Z0cpoELXcti21F4ZKJzw+3C+GrLsBRi0eq8TW1k45pQD+T1MaBE
14jiT/aW4lHNcU/mklvybaaC2AvfM1On5H6A8UGHuNcV+qpGdGW/maTlPej7lJw0
rQDniMxzZNraz9FpCuVOd0v+PePFm6yctqaze4sxNT2a0CBsigK13bDkQbVmYU4L
NnRRSRbxaDprgvU61DI1p1n4yDYq9f+zt+PS7YIzG9QsC3r8jiZYK43Pn1LrSJ1U
6/Tvs7eF8SocqlKp7gqYoh6CwR3lQcoQqCNXKzfTfAyXXOi0yA0ROR9N4vtJTdUa
dFUk1Oyt5rQhCuajy7mApLK2DFL/5kRwYuHGlt1F9K+48phbNZ5FCQuRSVlqMW9S
mXxfl/21lwJqS6LPgFywHCKgRDk2JEZGsfyblSzbE3vbwgf1fcipVffPJn7eYkCU
ewP4Szc+eU0WEW/ufvdfROwPXiJiMM0XeOS6XlCDQruE6gSgUL9mCU6HEEj5bZyj
L/REaAjBno7gX0luJxNAuFbBx6iD6m3WM1IZnKf0OloD01uL8olZESyAsToBgCg6
6kkOINWuU4yexwK1zWRKScI0IpHLtZmo5HqpEcdhJoWPSzi3/ONryfd5q4ahSbZs
492ileOV0nNaFP4XrXjQKwlo3RDiH3+X/POjooAJDw0t5lRDIQiSbrMFdb3Ou8lQ
H4nHGAmPDyygSFVuFqyJgG7fBr0QBHXpxanSoj+i4sUvalLwNsO1eYdQ/eFbVMGD
wI5TPwe/ni9WtOwljz9U6KoGkGL4k47G6Btl+u5CrAix/DBwXD3DllY6tUiBWLyp
bBBOmbkTXRGyb6+XGQBAQqV/s3JdGlifih5hkqcnYbbF93iHt++ZMQ2ZKUkeT0sh
F4BzCfaeFdTrtZ1xOohYpdCeuopBDOWQ1/fVzjxj5P+eibnHCttpFN1eA6Qwvb3o
BL+zgaHtaZWeLY8kss5/qkVK9TK/F52xeMnvOiU80tAv5eaXYCsVLjnAbSitD6Ap
MQ55THBYEjinhu/nRixwNW+dDRKskcjDJVVOb0906AUwsmgTUhWt/o9/4sVgnv5h
BKAhNJ02N8pgUuSs9otcFvGIDHL5zMbMWUh3gPdJYJO3Pfcs/Bp06kKLGaS2CvBN
k30uZomUoOZGAL6EhURZoBU+RoJAq5Vdu6RWAn9BCNiK8niGpDBQLa45nnyXMgl7
24e8N4Wq7A74pe0bCd0cNa9f3C9ynVyVi5L8rwPIfSwqdOk6r6wlI76uANGXOaLo
YAo5CfN7btqxnl4sUCpyyJxJVQvorU8L2Hp5amRTYjSG7Pfjk3RDVN95+lavm9Qc
d3K6MjURiKBkZ6C8Bo05PPq7+DRLlPn7WImIM0euRWSWZcMWc65YoxujFhwYsbkf
hdaLeRRyLUMgzrCrYyjqIvY5kbrZeJo7NKo9KKSDfQ5ZbINH1t1M41hoWES4x1c2
8l9Zv6lbSLng2BXkjYwwLC/cVisZFyzf408VT04e1C3057o5EKhTmEbax6WNXzlz
hPRjZWsArlM/XUKtHUDQieq+q9edPW4qNdWveujJAUYOugtSap4pXton3L00qY2J
fwegSfsv08JMPR3YLb4ciIaZ75UYJJpfJU/xDd+g0tqn2gJ1waIMk4XJu1qXbyDl
pPPBpBpKI8DnRzToJVx805RLNnkJF/i1LzV+ErmaGh234zx7xZ33udSTZBN4kNfC
9odkNCp1XzuJ0clzq3GAYkQZRoC69jdkAIEfgqT/rxO9IOgJ0V7yZJ+yf4G7lP+T
QuICe0h2Fvgc0EqmfyVwNg9L3kPgdtnoJ9Z+qsgzxevY/etXJT2//IW7b/5o5Pby
QevMLYFr4BF95SoFTdVTlGM/tUsRbTSvI6x1dflbDZqyHVtq7O4dtv+9z8JNq54t
KsPh0rYjr6B5KImKsLcG5JyjPPBq2x2L96B9txWYgO23ijUoVhQBJHKaGmXaB7bq
2rs6b4kI/lIh2cm7OcnbZAKI/1y5ZbwkihxOmS+WkITzw0ZMkx1a5lOiltchs+e7
1mY2+ytCcKrmrm1S9G0i3GBNQ9jCEAcrK0G/AMNunuky4TDtETPC6k2ie3jn4pdW
mns40pMTBeAVdlm5+qmJA+o9VQujhgf4fUuJdnJxRPyFBaxtIxy7YH8mOUlgHrQ0
eUdO+Nu4Y28eTpd/49xQxwjk74uKv0UuyhQKB0t/cKoHYOS6LVj1NC/WP/OTpHhJ
nKv2np8820wYIc9lsf1m8y8LQtfOjaouCzWBaTsFCyZabY3XWQlkn/mMq2X2cKuY
K+Q9hSzb9Atc+zn/OCPzXQv3v3DsJAd7i5ZKun6iEgXcmI+dSAvW7CA+rL5fTpH5
xH9MqlZgVLVX5tmUwhMDTUSjXmbgOTJzQxh97HM8GJRv15J/PM7b++Hb1i4qbUmd
Y0QvyRNTEYe/I/Tab3YBalbt4LWU32L1Xzc18GjHB+Y4/R4fKTPqwhGMJQnI8Qcy
5AJBvHcXljlomOhp2ny/Wl6bzS2uBO5D45bmPr4GsrC+HTQ8+SvvI5qwUzZgTKEy
gadHktqqH5580dCOGxO7duSc94qhwP7xtFyKCOndwX9LDp0LfVwqx/+qs31AIF67
/lbjghIh8xtZewWUzJ37WOxfWH7wnG5I31x5/UvyBXkhr5+dMs3xE8ZWFJ6WftSC
fi000ozzcfZFK//6AjaG0yPvx5dSbGUIY4Y1+GRW5BMrn9K5Uu1PEYQrlG9UeLHj
FIRhM50XhTI82FhguGIS+zNjTyKa5z9w58sf123Uihec+m+rElthDTbqyQHiX2by
71sULWg3IbPr9KKrIvORTkOiOJjg3FRGRsiVxiOsQxXQRpGW47p8chZeV+cjXRJp
ksH2sL0HiENuUu+n+KxHPh/Gzo/O+bPib/6PkiAolh72DP7xWzA5LSd7L+jdTGs8
7Z+BYuhvYB6XQ1BicZ3JJBa6xL9TBYDZrjL7JXH/oT0Zwt6ldjwL2RcRi5j+moBJ
MDug5TYMcVHNz7fRI6RV7oqZ2mXBARV9wDHW35rUA3rRActWYdz1XO5mm+n4d+2I
ykcIwSuJdbm7wQjEVUyaU2T/TOqfU0geGRsSoEFnIYf4Qi+MKY0h0AUJPgcXGlow
rntTxn/lGB15s3D2h8c0DatQD3H60k+vwEZPG1vWXLGWeYf3gShApVbd8LH5ihTJ
4VlCMp+m/DwyJsojWexzLlL2gVVyWoP5s62z5vINa3TqO3l69znIkIWWWO6Iovez
jl3+P6/x5GIawPUSfs1Pi6rU52T07LIp9dDnFn3YocFXGVw3o2OsMvfqCESJoYZF
aTY1eWqOxi51i4irvrc7qm7yS9YFcjaOteYtbLJDEP8vGvFumnq0Oqw6hyuKUtqn
91OsVzfjZfqmAcpU5kAQB9RZAzyPuieIMcefvCgEHgUlxPK+MevWzm7HfNciEK7h
ztGxkei7DIdHQjAHKxQ6LQ==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VUQ6Aq1RpZBmWqxH1gV0jjcIS4fwNMALV3gm0bzM2z+DfCnnVxmSXllDXe64/V1P
KxprX6DZGjPXN4NtU3wLIe54vkeHGM6rIGrIzKTBsK2tGil4dLFjcnF1oC8lq8Q+
5jOTKlwTcUTTn2XG2he8n9SwX4Qk/S4PbmlTXdabDpHNnXo2d9bcUUsfKMLGYadZ
2pv/0x8YfdbJ3q6oJRMeDDKzP30uBdqZ/LhU5V+lUVt3VW04yaLGZSdncERweQLj
5nJ12ZdQbegeO849YlX8vYn0B15rVdKz+jzgxwERbYF+km9cTGFPgMpv4fmjFhx/
2aZ0mbWLleKmokfPheXHZg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8048 )
`pragma protect data_block
lrG3eKlJd9wnJSxa0F0skitmwHusYh+FIhZPoSxhscGHDTRSPnN7QXYU+4j53bbx
WTwlOmEveBkmTomzxTGse+s6aaXI+7rUJinhWubNAOd0gmtoalDvKQQD5CjWe0c1
ZemFBS1GalVm+b37Sqx5enWfS1VxNVJSvKkthl8Tqnh7RyffwlSHJ07ardciNYFM
jUD3PadEueDOZkBrRMThJt7bXdkAHlq+Zqmrw4s/wC1UK8b7yOLJiBGR2ozXEjFI
+NvKr3FxojA55lXcI4levzqI83PxQOkKVTBnml3xEv+uySQMH0VWXQsMh87GKw7v
YZ8XWUCQMUymaj6QcTFgtjJCKDnBSs8OPC6iyHxIaBwI969a602E0hIUpIkgPcct
ptrCFkSXJSWLULikHtW3AatFBf5vxzs8qq/RZsSrr9I58JOZkn/RQIhAW05Ib9Uk
Tv4rFLwxDuYjidIFREdA66+ayiGjpabW8KWmjMm3wycnNAMIf4ut8Aojk2oIRRwX
vPXnibVwCGCIIq6vv7g37PlgyaiRc2hKpst2+ibnJEstTYWZec8RAcB6KIrscG/R
UkagdGtmHi9IDOAtYz8tf/QMNg+EP6Tvag3mb8gt4Z7xV9dm8UBaJVe10XZ9l+vo
pJxWSOTr4xELDfcJBhDSAm0L4l/WF51k9hZq5rED3ME/XILqudYNIdPsBU8mpyPz
dgjL6SG4fMMIBPYE71hHzTSUodZGcrm+txuHn+TxyHlwHihGxqn2Q7b41MzeGb8u
U8ydktAjCz1uuw40h4SDVmckgDZLcZdTm1Yb7K1z3FItAIL+Ki3nQr29RwRkvY4S
Ba+abQjgxlCKR4iR53Yb3MajbhRRaVlCcNVHXwT4dUXe2WSzjLnyJ0H48GVkMxQT
VsH72Po8x6I2BYcVaNDzCU1/wxwiRqG0Mgr61u9cpzTX5oPLmsnsihIsoJdQ0B/i
k4JLtjD7PeyjYSShyYgobrFRH3BaJz1Qqwyp/8ZyLDGjGeqR3Kq3QVNvUpuPMaYZ
Q2IP8rnOzN6RoU755/56vCpZTe8VuXX0JDOygB0dqO8m/XjyTa/lS2J+k/7QsTw1
7s/J90JJTA9dmBzt4Hx7sLzjUvXYkn65s8/mVQFpNBvmuD3eZghm5pGkfMSrfJ8P
TBfff6MchNi0RqmcTp7vUBOcR00x99VHGyVyqGm56hqJmdMhaXvhDixGWoh7PkB1
DlNz2+axIxPWRfrvU6L1XG3Ng1+u2uSANtzHMydS3/z43Cw2oG7UoIHS4mwTu/K5
V4X2DV32Wve5uij7aaevQyrtkyNXxJCX40lIRh+rLrTXZHADaDgwxFkwpw+ir24v
I532FUNWvSg9mnHsLZUH6VY8cIQMLySmnrlbndCCjT6W68brXXGO9V03TG9SybZ+
hrrbrk+VjJ+xqcR0XnBpt6DV/55pvvlGVM9N3hmtHEhwuVq/+AMZ08ymJPh2v131
cBpFayxY5hmIXU7AoUbR3R5wqf3uoK4GuTKCQ2G1iI4yIZiyDcYa0PDvjNViJMZH
bCN+ye5XWEZJ3FJemOraV5U54ap1YtkTG9lxKwMf3nSiMvipFxXN4LDYpKYUF+Mo
/DZjLl1R+X5BATEyh+PGlEfUccam4op9fCnfI0LgYZX31JzgHzePsx/RbnIzfOj3
S07eYhkr8A+w3f7Cu0YbcZTkyXAytg+QMYUpEH3O4VyhzYKJ7iThHZb4zR3CfLEz
nrhfACcjT7Di6XVjsLsfYg84GbA7vdN0naqvpBjs4aaBND7GHGRVynvr2iUEc+nC
MfeO3PFyrJSZAr3+VS06Cp34Qekh7kFZlDw47OOHTWzn2WF/V3jw8xElnnbCkqmN
bxoy+bb4Lz19/R3WTRE2ZLkvw3Dj/A6KMf3jpL7z8jHMeCxivikGgsaOZd6Ch88i
qddNY89wxtJQcnicGdeDb4uOpjxAQTBazEn3BPedMbSzuXMoWkWFRI+Odwcx49r5
eRdw/5Vus1SRyCYvRh9tYJSQMLhAGe8AkmQpDVwAy0rF0pR1p/3nqVPhCbV7Ts1b
QeNgIGjMuVRzbzd+GQm4JcsmYDEsOUtj3GXeFjLChclvMUt8SIed/xKAWfmGOiK7
mSovkCL88d1VbEz8M0XTLHPdLfiww5ZXmdtvFMC80CoBaZ/BDrAe3Ux+8Y7O0UNV
ECeZCxqkSZKOAe3oivH1icxma2vGti19Z7timcB8WzTI2cNxkmKPV4D7v528C9TX
H1hCV6ZEMI77rX2OayGbRDDj+E6woHxb3SlH7144kemfGDQevkYX9aH5u+mm/bU6
0JwAieJc/xlDbebWpJaHZX8yegKAvHK+E0Bm6AQtXOEtimU8ILhyhMFwT462PPa/
5i2jjLGpiArqoR4zog0fBB5LfcuFcBJksnW8G84lo4npNBpMgRZ6RzaIITPKvPTH
CtiNGbKjIJS+9lH/Lu+RjEIm84wwU94d7pnHGxqr1lQG0dWxpyUZQdCJfyO8TX/O
ZZhs8kedjcMh5KySYxY7Hz16+TxU7CUQMDtMHvy+GJ4TWjtbrrFkvNE4ujUiHhoQ
JPeDSNlnJfMa5Ch9BIxOhCmYjyZLCGnJ7oU6CSyW7qgy1kwrogTc/z2PfaYsSttO
h+cqH65FI9xfpATncJTb7uhHChUFmYgVWt5+DDGY7ioV8HidEmLsNMYfKm28VUsv
F2tWNaYD6dhF8DchMvCaVU6PzB7NBFFZV0vqwk1G7aWtwTINBDEuDD4AdsbQnwJQ
Y5vXHsBHtvMM2hyi0DLH2jtzueqfUllLB+pO/VEltUocyFzAdvomGLU4fZ9NlqU0
i46vlEeMmKki4CS8RPQkEIWeaS2kChnx24afsDNU4vkcYiHBWvvwE+jt07VtxedC
FTIWljXWsFUdoBBu018B/ykiLJVAGxFGbTXdTSD+WqzJQQDSrKzSterPsvKXijbH
f1DakOtP8BjOSyWpuDXY/8z8dm/Iqpg2r6IowHT2hiZaRlePPB/n8Xtit7NUx7MK
MC/fJ+nIZArT921kILr9vO2luO6M3MW3HbBjM00+UhCCBQDkC+LZ2b8DExMkwDtK
q2surmKHaYHaCw4GsG2JgjreY38tz6Wegy8RmxSnMcaas/2LT9QCGUab2kFBGV89
xHAt1l1avfDEbutYU2gy/Kp9wtB4RnDOg7ooQdPc+cg5f0opacHzOW/n/5gcz9lJ
jVHjez+aJzLG0foVYkB+oTg6ptr/zNzoxvhvbsIZYVImZ559SiYgdboY31pIqowH
8bq8WhAGout1cPiubAUZb76oaou8QH1lLebqDFBOtaSqFUL3dibTv2guYY5Mdmyk
eRObe4MrNM3EPo68O5tJmNNF48m8MHy4mBH6i5XtcMJyASDAkV+4CjFA5i8z+1Xa
OAgwArbbW2Pc32YJrIbb9CxsU9ughEAnWkjwIpU0Z5p+Q5hCbwqjkqTJbN5yfkvL
qcsN0qiCVWdFWzj0Pk1hbr+6LMA+kkRBwSx5GGmFfxNVLOB6Sgth3Ts0JZoU84yk
mIrGCW20+aodB2kRCYDcQ0ZbkCJRnHv4rnqlkHP704wDyJX88cBJc1TDme9GpMIW
DpTT83ILEYtqicoL8gASUEQuj7UmMY2wGLtjIowzD+3wPsJn1YNVs1n8COW9szSk
hfWJnehq+IeODKLN3J9/XivaYmCxIaG3ACewexqNXkGuoOATcg84RtK/R+0+ylqW
2XkN2BPSpH9xdh3XcLMUvOK9sUMzMvgFyth0et4Cd7Rqm1+P5E5drehJ2QVO4sc4
W7BZN+PgEsbj1ao1stoaFi5ZplnaXrIIYTHoHQs46WXClOm9mcoOIXitLRrBavBj
guDwVMsnwFsgyaowHZj856szEkW46n3lykX7O2mQhxL6DV4kcTah/An/HiTnrEWw
tbGgDxDuQ8GmhY52hgMF6eWs+RPIg6KXfKDeypTgv9CyksNL6Up/HG8VkurFCQPc
f3UDboRoFmDwimFH0F9oxht6c7YKRa1YpahZa6D7bsTVYrCDOwinvWyxvAVkM2qc
H0kIZ+BzWhaiTXD1TKHh+/YGaKePXd2eSXLboGNLdTFtwRIoO4Z7tljJRplq45uC
tlvtfCHW8G1vNvGTpBqb+sdj3d5PstEF7QKxFAtF5G81hx+wwO6TNb1C6KMD4jGI
aDISwMixSaPhOs6myH9vxLwBEGihn3SNctjKEAMDLdaelst2yJmQBRIQWhWW/7Wy
P4jDoAw43WYgT5vMrNatEpeJonO8woDnbV8uxkuMJra+z4565Vwu+OP3v8Naj/zq
Ks3XpBPFkhpcE5bN16DnuD9FN1bhzW/omQBGGS7MLu/ZX9OGq0qq3EYq23uUJJpt
/Swn8wrEQeEJZHFT9E4X6Gn9ckEO7sqw/EYjAfOjpgRsnLm6naxrAsQl+IGSFPZc
JBrFlaFKnP86XA/FNwUxi0VcWGhlDcKkrHq3obJgsgZmYbclyss6mjyIYtQtzqYK
EQsDC7UEe0rPfQVmQgKWdW2BrJ1TXqDa/BUS0uV6CMq5okQhVc7+uW+w3bBpq7Iw
8Ncun3R8MDz1058GcE+HhZerP4NJJPP1bxhG0sj+Q1MRjIiFmkG1Nv8/mt9Zt4wn
oaOJhKfgR8sfRUqEpk0oEunj4Fqh5KVvyF5mzcoftoqAp78rrOopfzRA8lJ8rL+n
iG66OdBdcs0eOWHsQUw7GEZVWNIcvP4C/Bi0AY3PX8kNbyaXkgb6DCaFhqc6j8bE
OSaPDG9C/mioCGeXl6GG+t+Dn8vsgOn0fiKd/xLocnCKOg+RVe/38203UrBz3hlu
q96B8ohhHS4K91uI0nxu2s3Rd2GYSsO0ucRuuvpxComixj9K7lG/CAD2KYJg30PC
diOGRGrSYOpJ38QON2POCw8o/PH1TijS/Aj6kkq4pRuK3KrU0SGeMrIOe4b+BSi4
EWAHy/mAfzOjgRvbdFWeLZyJ9b+FWWB3qQ/l61rtz4vfFlRDmef+w2v/fqHpp26G
mQ9ykzECi0NlOXDT+gM0ed0MAbBLnqIMfcNe/Q6aCJCHA/grIg8uPQiKTHVOSTgx
GiNCKLubi3r78G0BOZOAyfzOie4VMnrQzkhkat+Qgmlq79wK04GbVpyDe2LWmepO
We7xcRZfEuYgwNnH2mpSzD8bSiqbvWO5pZsmm1cunHFmR9jwJjc/2nFTr6Vi3y6x
zv5vAIGXPCM3BHQ7x1yIJ/Sl1Dd43ycbdkxLhQY1KQPbD+cdzo4AcEWJKUB1w4MW
oz1ezdfCtEwV+f6OPyDxS06lNdAcKXSPdPXTZiybNNVdGjf75yaDkId5tcM+cw7k
A0b6FxXwpVn2ocqovTjcYVACfhp7S9W9gB+amSQdVLex8vbwXdRdy8LYwh8X+aqV
+uoVO+keUqLTavlnc0V0JUmelZrYYLZYafPgqAXRMaUJqVfTF+f5TnDyPWWdZSwK
3QoZBv8Rwt+ei8ggLEQ4nPWmHGdRQDosNEEB+b0U4Xieq6r84RvLh87hkYE+KYDl
OfweohDfBnOS3nc891Buy0Jqw8Q7b4trkTgCM/X6GKqEvxJHQXxHoZGxY2KOIwcy
w8vCggykG+qFdxmR+8QDaIAzNCjUYoLIkUR3kHmYqF5UNikuV+uQLEDzL2wTXPy3
dmtHO49WjICJG5oyd3PwwFwarh0k4cE45P9fVJ7xqR+QYko8fFIk+rn+Py70sH9e
JRvTgy/ue5/CVfzTjR5IHXQEnyiFC4Rz3zuUAMjTR1Rw4WvpZ0Ty+en5ihCkLGhd
0QfM75+QPJJ2jcanz6WudX7Bc+LJQUP2CFDyMGighs1Gfg1KzWiCMROlzz63101I
mVspigMNdSBCqMqAB1HF+1Sy3eAZsxHor/YwRxkLtwj5RZIJ7PWZJeiqidLtHG21
HeC3msbTX5+izoMA/pYyKGV1TkBvevFf9Gx9Z9pPbteha2P9YlZlQR62nHfmg5C3
NhbhWbws3fosqQqQwB2Y/EZl2d8i5Zs1kbo8dj8fhv+cqZeCgHXNLAcpVnRqwdTo
bMtU1L/HpdjNFB8m4uGSiFhFFawQJkSe9q3UrgIdVF0cajirSLvQ7jVwlXv1nYsS
SX/NmicROOyT9669krDxJQl9xQvaCfb91MrEF9B+fZnjudk5TGUPoQKD78DXn59b
Iu0JHdgyJppz3LRlC+7iY8M02mt8jhedP0nbyYGa3AWBiVp8/8nTcPz7zk/YdQ+V
n2oZa+eByh9zzxiYLyCz5WoPwiUEe7hSAL+zfnAnQNqZBvxU2rCE2mvW446emwaC
kg92mlGpXhtPmUrk7dpujj4oygNgcqRq33F3EzS/U47ZtQTl4LWj+4VnoIHIHgwl
XIy0PSLydn/A+mg16qBn2ke6nZu0MHHHutfr9Abqsh4HvzZPP1l9LOwkxOLSTBf1
7NFqlytRNriFCAmlobLTTjyVuvZ6y5o7vDpCFxLo1ei4P6FOn0L9qM527Ofazfi6
upAXEbLfIpWuwAvjB2/m3CNcympUldfc0PcY3ZPCBOkrI50rUm1OIylpfOsp8VVi
AyMxrcxHD1dN1g5nP2eUhx7Ls+MvmOGHNUn0isIjES/cW2VScjTtMRdpbgahr3Ry
L3wI2vvu8w08RcQpyW6P+85ScT3dGNYC5DuvsfHcTZd228Jg7dvPIk6+SCRiy516
sG64PuHcpXCHpSCUZOXbjKI4PbZ/nhL6M/rqQbeIXmyiDUUQZqzlSOxOvawoNcUW
QnHk3JALbGh/CUTeoJ0jU6plaFLKt/o6lg+TbZ9uGipYWViux0UAVGlyKVdo73Dl
kKEsfyJBp9k2iq/GVhYVG3p6rv2cYO+Yn53S/7JW1ibIG4WYmHMYazrNjKejVjPy
MXQVCx7raaQHrRof3+NEqyJJP0YUVJIBF8P/ZeWxMXD+hrEToW3IYWi9U3H5ZtBY
skBEbILFnzeyqTbGFan+b6blYBJju1ewzDtKR1UzlDL9O3ExpA3iIpqnBn+tXKI0
e4Ewyx/U2L3pCPK9CxRanEjPqrTlKtbmPkAXb6AzbFyrP0f7ZfDHimI6LgHootVa
A4WbgPGnXQxMsXvrfoQK1+SCS0D08bBcBf4Egdkreg6MWXSr3M+GMepmOjbzTqdt
LjJvk7pRpw61nnFhlp1rJTbIFuYAiD2nRb9n0uEqp2ApC3WTn2bOAVJ44QIJ/rHw
Fz6CzlKb9QEx1mpYxKSn88lnCONQE/xQKI1LeJjzWh3Df5gxgWbB0dzMIHcPSgW7
Npo4wMbTf8bWOMBjwe6ImYRiFYc6Ytd6ilxSv7GX9XNe65rSfBMoX078I2M2RdQ4
oLXJTj8Zl2u2jZB6LIS2JS3oo0Qv7VMzSE2V/aujcjkc0m2m5t0QE+4Zs52zfOSK
T/BltPGfw84AEqeNnPCJMPwIrzcWb0++6Wk7GQ7jh0xzt6MF9YE8YgDZzQJaQgsW
zQ9/vBRXNeFVVqbZ3qlW1t/K/1bao94I0uxnBa7DrsfWmJmb+ZchpiHzeHTD5/D6
UYtCiX/V9thsJwy5jflhLslL7a6tKIlSxRpLICSyZPJ7eZpatcORW+hm6xuY4Any
37XaqUsVyBQHQEcRl4VPOSlNxUwCMJ7U3jQDVSlsUqf+iUERj841jJzWK3x0+Tah
owrc6MNCO1rPskGG7Wvj7LUVCOvm14tNytq1zF0wtdG335WkgVIGRqiGIlFo6nDq
G55Nz+ZuN42Ru8NQdi/DVCeFf9vVwtMxubuY3FwEWJqadb+AQIovF58xVrOlgq3T
u7EaxKEGzuvzdUUL3pF0jfc2ZOPmbY0ezXoVVgdXJJ28nw9noCExcHaKfPTsn43N
Rbuhmm9jqtff0XDFpa+TwXfTw9ksglMI2WfYe6VUKvdDJWhZXCDhDUAqMStIXzPm
j9NPI893NLTSxnvIA/oMbJeD19oNDeXN1fxMeJJjV72IwqftPuG3xlAl/1pdNlgw
X4bh6O7IxJpBRkH8LUQirAUbG8/KvWwyAqCs9WpvCfm8EnPR/3+9+zLit4UeqWTw
tQd65EqC/BnuaKNEbwJe0AsF1M7M1/ZpEq9/kWqIOyjz6B025RMbE862R8wT5BCy
M7yIiFn47o4s1ACzrygZ+6LERfnjKkXjOOugAppzax4uQlR9kQB4c2ELuM0pqZYP
w0KPQvEzdJGEVUyQoIJgnW8BMRodSvqnaM1Afzu58yGvfreGvQ+/DbmbXRBVhaJ5
mwh0qUZthkL0NyWUXsqIAsT8W4Y0pWb90KlPqIC32jo/r9ClNkGYlWtTEhXX9jlA
VqRgAixyFOxslvnZzUShYuBWnd19j9m1+D+AvfEQ558k4AE/Pvj2/BBmnTc9YEhu
LoWQjNkafwx1xEeCifnrYuPRBNrXVPw8ptPiXuEtRkiZgIuTYCP/iF8eq6MOZhpn
uZvxrdxZA0wQsFw1N3AHznT9D6qUjbHh5/Wsg8p6e6Gl1XE+qeszOLoI17QjyKsZ
DxfGccXfZ6ZjXKmtTyBrQWjaNmBFVVvSCQDSUEogxlPLWNLEkOTI1GBhIRYPq+Mz
WBxoarqx4/U4hoHb+CxMJA9Pn0BCgTCj+1w2LRJXPXfeDAmYKQMHZCa9PMv9Ep9W
TYq87uz8yOqVPN8DqOdqg6+IvcymN3g3Tiex6CXcDPo3BR2ZIZ3R4ZrZWjcZWmfI
l7nYfm9O5kelhyDo0A086ldMkdtKoPtJPWLktQRihTPR8/UlsLp0yeJ+fgSdIveJ
Z8theGLTGaIsZcE5UqQw6JT/r5bGx6uGGyjWHANstgMqK5TjuULKd40P17w+sTP+
aeDv2RKfLFdFekG4lb0C38zxhs0s/LS3A4/u2F6wS/a9tndmOLks+CtzbEyihkLn
2aPgACne8KLpPhNnGN69tCfLYG4YV2kihvVHM0AYO+7qxR1iHNnQwmiVZFTJSfaC
DCv6peRvGZ1CSvmSW8/NveZYZPjpBbSvumdFdXSVg+MSthH9RfOG6m5yaQWCeIYY
BnKKMkdOdlzXqKZCRmLVNrPcRv9dQHthwBz5vEp82jTgHsNAs7c+nY6vK4hpXMsz
FYISZimKRdLdgR7phG5Ei0gdP3sEUSGha/jvjm4weOE1vy+64K/h14qK584mixWp
4ZWFa5zxx2FOZPOdwQCzasyf08rX+fKAjo2MqAcniADLJbs6MbCtsGpAzmEf3QRT
eeruVRs084p4SW/dc2fBokaIUdjOixU4KR8LUl4A8Kxl+k8Qn0c4u3MKVwcYSgiK
1yjVd5D0xO+SGNip5YzeGdIgnxe/yfbshPvdpPRnSVqtU0sZ7sfB6Pu3cDGspIMH
N0lZPJd8Z/pWq3j2xzLQZ/v2FPVAcljX+IEGZXASK2P0LSawdogsP65ZSKn/f6rL
lTj4ZHGfCXzwzQEkuBVbwxcoEYc1/PyZCnNoNkPtGnhDAMztm4jFP/abMajNOW1A
zETGUmd5L/xYeVWkG8bdSN5l1jReDFwTsDMhXT1tvi9AMmrL5rqHMRM+L52MnZWM
WKVjknZFqrBXkCLeu1cHuIgr9m4BPlgfG7vnhEu2Z4ob821cw4v7a/lTIIwBVdx0
kNe/RHc4Ao6s+tBwb4sQl8yVTlnkFkfPzjBeC5ti23ty9yjc36Kup7Z0JxUcZEqO
r+BwH3aNn7IrEItQrBAGl1eGH2nOMCjyjkNA/KKaJQzLCmmTsm9mtLTjt7FoEF/o
p8s4bPJ6gCC86XhWkLZzgInaUw78qNPCx5xqWMMaP47A9oTdKH0gut4jbX9FCb+i
yueGESwlD1TY6j8c8ATOEZl/iYj7DbWQhAgGqy8E5JgL1Dt8kZFHvQGZQipJ6IAl
PV4LJ4Qv3qfH38CfEwMsGnoFvVpsHkeZswPllOUu8RXrIHoMKlzJwi1XexHKPi5K
WVcLLKmrr8uHBe374sLqwPbPy2T95s5MwRyvt2tRPANZ24NsQw6RxEyB4TojaVsR
f1bGIPo/fLQrgi1RO7uay33u6vlXKhlNdTJlFlFVVFs/3StUuHaazRcKOupO4COu
7rqN9LD7XHCWO3VkBUzGRIhDCKpINlxFMa6bgw/Bhpnz6s8eDgBfsC0wnFHfsL8P
HSCBHnWqjoP/O9JOLD0dq1nzc2Py/Nh8AUuA4J+c+Gsg467lU++xcxmON7y0Y7/S
4hedOvKs7jzQMrAtdMxGM306I5aPDeqQQ8KqMQwyShuoXUxIL2E74KGyOdmY5l7F
3X6IB5Ml/2ssJE+thX6p2OZT6TF4QvsE6iap8CXMkaF7ac2IqK5U3etmWJMSyKqg
6QUOiXDZUhW3J81/BsnwWBbuP/f0Qk5JlPe4Aa6y2eY4yiigaYZlbjNW6YCDitT7
p/yg6muO7y8+62qTcpzd6I1VScolmpRxUj+ih7GHgQAyXNZlA6z+wkywsJZ+UO1R
fI5/FcHwPfM212P9seAP1w+9LirPEOKQKR/YN7VGCd4lUgawjOZpQWcktHEND529
JbEPpMxGv6Ts2IzKrMdqTaaqYYAkGSGlpMFZLbfvKm5puNywJWLdq5twz+/8IhIR
KQF1UqyesYDVqwpi8KZ3eLrSpd9FZRMxCcIHGM8zB2GdReDE0qAtQeZ4Indk7FSW
3gnca7Y6XvDax+4wxl2r0qFKQPupIo71wtWTVNQ8N8/gMA0mEjVVdNhceLr5I3++
zkI3xqqKTt9l/U1mNVjkMh7i9GSfIo3QAKZhoo9/6nDKaMM/a577gD9LLmJR1nE9
AoYN2bpc+u4wzMlBua79uGusBJBus2hTQ01TeVjq3gc=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
eN4RIYGSJJazrxdxNMcDF+mRjDAaKvThNgCczSHIWGBDAMCVvJhmJf7L64fH2PZV
+by/RYIPm5TF84D9Hb8+tr9dGXQQ+rEh2HTtCwlg1SwNoJxrtr7GyqhsJYc+xnyy
QvOg3TL/nqNFjKWY4IpwjDpn+uaFCyStFR1LgBMFHJpgHgVXdWL86X4CBEQhfik3
SB+Lg/jm32uoIMlDClej6gG3xtjqCDwEeDsamqTz0LtRU7ggE8IBiHyC1fpw7MDP
UPH5dmiFXFUsCK+482ZMfpu7Gg7nwXsegOebEWF7w2qIZVEAdn2zna0ADDuQaqW8
AMbQhfr9xqYjSyoCgjOGdQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5360 )
`pragma protect data_block
XXsECC5Thk7Jx5kkCDDq4JQ95hqFlRaYi34QUgBUshzjW/aprgFOABNUWRle6pBk
uFNqzVKv+0DYejp0msYg+jqrN5OGj3XYeM3J1pHpVzwhWT8VzhpPu17tjGFUJsRL
cgd4Zfmi0NSSkXP+stDNPyAcWSO3FwUjrS2DjJADsB24x3sC4nUii+d+waQhMXLU
AG/bLcWhUlWcVXFsycFfAMu129VLQS4SKx+jW+EoNbJ9CmglBdkLvGgdDNI/qwnu
anJkxHymXVug1qTopZks2MhCJKGLHpoJwrJPxCs5T9sQUybxfRy+Mp+R8au4jsdZ
PpDQ/Yz89iobfpPU39vxId1uFN/bzjEAJqVuGOIA17xlaoaKUWlnSRxgiJeFY77p
ZCJ6cLjG2gJAFB+FhO855FemKjEOxG2m7O8qswHF4b5rPkb2BzS1eGd0QflNHkVb
vKtKHLgbj+KxqJqWugsycvyEd0+0yA/dqwl0enkq++pyZed3+9GBrFgEq9H+/wSy
rj2F/i4U02JaxOQ42Qkwtj+0jWnxSCyJ9ntu9B0dF1ZiIc/s1SmSmkequd8NRAYQ
UCu4mUji7HcEf30TvQByaCWFBmOPno69x3/cxG7AkzU9/31VCCgHHtCjSOb6egV7
gKZsMzMlCILmEEFq0OQFPbukLi75qqyNi/LTOdIw1R7xVd5vbKFzuqhLVBl5IlW4
IU+ZAT0Wsl/NxUoGw9bCOO8ad3Gy3UdQ8Id72L5R1vn3eGJ4Rode5x5Nw2xG+zDS
sP8Va6JKA6BY8exkXjPecyaadXZXjq+dy7GCqIVRQAhXU8VvZaNjl/XPRZLy8nf8
6YzxXL/mL0wsk3oDjMS5tmvsA2/WhuyHCfAYjjgEQ7KcHLbhMrKRJ58otUJXE44X
fM/2FV9iQEp/Bc4KEKq/fk6vffXsEbGqCw86ljLJNzEAJjQC/n1vca5+tn9/dEfw
Hk2J77FxYtqF8rnXS7XmJgWvg3EHdpijg9TyzsB9nPWohvvvD3DXAqxBMtLikJ8Q
i1bkATY9rWcqS0UKuRJ6aKvITerJx3pprnzi28+ZGyY1+btSigFJjDGFpcTPyfRi
LEyeBFUqE3rC+e/l5Csq01vndCB2HgR1uDPEPs8U3lNk5VfE6P7xK1/fJ8wp4u5h
Y1jiJowp9g6dAzcqbqTliwbLAYbPZZjhKNBdgTWlny2kYnCzV8s/s4Fccb64U8li
a61pLZStWdr1IP4jRiSxR+3S0cDEw0C4G7vxg6Yp6Ybx/TogE/rdAOU8mzy4tc7O
YxEKvzMHjUt93gwZj2wm5T68TXOcWJL4FXhfshy9YdyupSOlpHR63ty9TyTbU0hI
ZSD0h5hU04xSzanXwo8+CsNZb7LBMgps7eYuRF9pnBxsx1bWmGwvEFn2I/eGZbms
JrCfnlMLKz5xwO3vVRJfollIU8Kcd08G099a7sY6plKaTZiv96jszWrAGKKXyPNE
rswvGF0jSQU5yJLukADtiSOofyH9JwGg9d33Pl5FVqDZ7mXTAgKwnIGtan6C6so4
N0akOifgrD4y12VT+xgQcEbjnjBcNhNgmnf2WPSP5ibsEzXKlqwuGBL0jBpPqbPP
HkP4OnBRapQyRF/piBQ8M4O9CRCyiBJUiGWUVzSk/5GKLtRO4T9gq6ummXdqt/l/
cLpGdfGjOHgt4EVAt2SD4hidJrJMwINjXJ8lA2eFl857GNCHs7JO/NowQ58pk+HL
Cunmckvm+mUl4NdivwVdbaYry25NPB/3L1jAg+IDGBX5HBSqqywg4j/wbdAS+r3z
8umOe99ERQr4Ay4iJ6w9x04F5YQzBy/Or5ml+dHBs18e1OzagDuuc17Quu4P5GOt
tNfAZ2pvYVJwI3f3xn7bQFlyjM0cEmQwRQZEjN6HbzOexYLKkwajDfufY35B1lTx
PkbrmudN3WIdTx59wxntN9OJd/375sIQgGxIsC46DuesrtRPimFCUUM/RocFhLvn
RcxGZSDHP8feB+nK6w9Fw1SghV87NsT7k9HQ7tgguE3ADJb5eYRO2041yFA3Fa1e
zJkcXFCaset9yS34olad2OwsMtapbmGuywMLcSA0autmZHg7Juua0bpKjEXrXfDC
NcxuAdiP4wd0yQNcYrXFQMKppIpFX7ApLbZYOG//hnXQfC+6BqfMlleNp/fLTzuO
87m9TE6/coMKNFAigepDXxKGWKZwZ9Wzff3Sc8gm7fjJvkg4urlxzJuVEHI60y1N
KfMdW8MymclnCmVAN7zQAk7Wur0ejrz0QoYoe8k2CGGg8dEh6raYa21XjRdxErGR
4OFyN58+LKi00xDaVPTQ7Y3N8ZDgvY37tm/tAD63jBnvPZqfodz/xrurDBXCu5h+
6/Er12Ads4ZzMD34zoosT+brGciDwxqN6xOM/RukZXfO8Hvg6OQJ0JGjwhSpr0nd
oHP0cLDZlMybphpfWSlEHLbm8vbugy4O7RlcNyOQHif775vNy/JyxlV9f/Copemh
ZZauPNTdWxRvywBgh4dFBBWlTOcUSnDc+vXXNKDSW0S8n4wHtC20C9u0C1HxtwvY
9+ff1cOzG7TPht+xXXG+pUSZDUWC4olZIlv65LESfXVydU6GnTM7Qr+hr1St0Am1
tpVXuDhC3kWQOxUZzWFPTkKlbfCiJFmuUV+I0xQZJJ1MDw33IKfKacsiRMM7XMDu
YWBokp8HJPyNACjPcCqsLrtalpm4pVIfqFK7PZqwkQ4u/z3MmEfG0JgZn3E3s+UV
Hdp/PIGnLHrV6hEpk0KXx7h2767nQaweyt3EXSYwYX/MzVd+neePCy02pLYxYlCp
HQebd2gqr62cQ6PRLcdNP5VySE1IRACJNFWn53Mre+6reD5Uwwz6BdblHzk49xwA
0H/ETIr0JYgN+9tnVdYfYses5+4KAFIsuvOwGPWeNhdckCznQJTDWXzCUvRUzfhf
c0DnIcc+L+YE28V7F5pwDf9oj5bH7LYvPKcMymrsXaPCW6ygTykug9vpD4B0sxZa
BeuvzDPxJFqE4+zS4GBm0hAbFeHhR/WnuDTl3AVazLHLrmsk0dc29tV92s4ejZZx
Ti2W1n2a71rr6Y7dW612UzagK3VXpfNn48a6OnCsZvODD6omOCOfkpxN/BryxLQO
B/5wooih6W5Q4cgrKoqeak1r+G8K2lEFPRlC1OIg4evFxv4+trLOfhA6k+1MHhuz
SRvcWZTkOrkwoFhYldlhKAwL/FCSwEPpcncQOz0lvpXqE/TOYCEVMUnfP2lmTU2B
HJ+zK+oWsjDLUjqP1L+RZ4YZHWZqUoUd+vm3COoGzdMKMYYPKxhRBynTIK9GhM5A
3LdL/DnLDlzXile2iEicd37/PCzpB+h/LAch6n2ms0uaP4DdmQPTsvQfRrmy0e6K
/vGtSgVD03MPGLOwCxJ53N76iNK26JdUSbhmwuvma8KQ4rDHeEaylPRwXCj6X3Mv
Hbj4GGOpllq66jx4xiDiy/U8PpVmO5fDV4ry3vw+Yau4lLvSRovUesmg5iKdom3x
8IobIWg7tsDTthxxMN2AcD5IstNanwcouiDSj6UsXd7140Rbngy7Qj8A8sVWrGef
/eTZ/GhCxogWTCRUYjzUsCx1OT1oGJmZ7XZQDO+Zbyuws+aT4Da9ycwjZJcLsgP+
2l54YotbPfzeaR5LJ1oD/YXLCQdHoJMRfj8uduPuuQcNNqVhvf03wK0G1+biDrfi
7vV7mUSGAMwZiWBlf4nWTGVt66zPmF89hLqQwd8Iw0bwsWv95fS6YuwQuKHfIWuA
tZ1jsYu4hU0hVlQnKaylMq2jxS9sIkGmTSggUDYIrU5PSO8JAQAJCWZaoq2wH54O
okS/4mHDGedffDCys7GfW5aLuJy0eLQw0AZC7kuEu2/JWN84o8mcA3NUFnM7CAhL
c7qVRy0JWuVnDJoUTxt8GTU60rkRa3FTWyV4IzwT4Hl/GFggUMJfZ4IKFBIvShoK
yQhz452XDVws2xkcUbSrvdDt+bRPTkJAvs3oysw3uF4KtlAc+tjRBijvrkL0pei0
t4NzaMw2Uz/SuZKpV41CFHUmxQ0wLXUASLbcURhsQxVHY43g7bSF3CItgQ9x9kq3
BP2VicbitHbRjC5EXqG5f8etzuYro1csutsNc6/I1tFt9zc6/IIWgoq/lsbotMli
fvnOvGbZLMD3sj//4jrvogi7DOlGOmkphAWQsKx4XEwMVVQp4WWEnSONN5OwS15/
+5vqoZwkUTe/AKryAahsX7KP8SFva1CHsuUd/NavVcQ5hXJ4Ju9c+PVZw1zXONmq
Ov3SMgUWsUnmaSI1BAwvCepee1ixi4KUO1vrRPPcFJU45qATj4q4UiaxgctdVb3R
qGFKETWN2ZYrl4G8JQznVD3kpQ0fc6S7/HCnsK1KCo6HjOtELO1rz2TRUeytDgeI
HDGIKgpBCc7jn0vwk9qN/yRHYvwrTQoV6huHFCkgTTklHKum5mPRxakjp0ArdUmF
mTjHY5fmmJ6t895pyy9Ya0eCeS9HMr9BnEfh3CUPuQCxc0CvubWpPnHdzLdDETUO
mgUegtZgXvaCpR3XSEfH9oepOvTzixkKOomwyOhdh0n5Z2egx6zLP56kArTP0uc1
3cIK6uFkx7DhY23Mk8hM2snSYC5ZL4YBJbaAQfdc8aIeQws/fY7JdsEHjP5rDkaX
7pGoeeV2P5bYDgRbvO6EVSDPlvU9zSQo6EarZQmaexHDF+0GatMRLiqwAhyWYfID
ql85Pq8t5SS20h/1PMnDG5wI1h5h2pFnc4fJvq5/I6SwFsphltgfElpP8Xm2kHRa
Rr+55VyIpTXL05FdophmZZFlg+mdt3rIfbZmYAXRIgqrqnBq4qSyn6RQlqrppBS6
vUYnU5GvEdp/7uCYGG2oO7e9w6+6dqY2wAmeWhwIPO4a6WSZRbHL9LYNCtstsOOV
LQnMkQteX+NtaLzu7pzoFNNg1eXRmoulVmr/S0U/klxD+mgrMk6YXz+OvZoWG4z5
zDZVMs4//g32nOm+m796tgq+p75ea4Fn8K2yGYQaCC9CGXY8ZqCwJ6RZwn/Pjvs5
CUh9Ewz7fuNO0H8rkfJB+Emion4u/xwlujgaU/wlclzPR3kY6H8EbjD2mdM4xzf3
uH0I18RXVXYzrO4ybuNhdh1pz2/AG0ItqGB9f+bmI9dERwj0Zp/ykIjV/6bdAPwu
SLy4PVrOK4WlZkJGNroia1aH1J/oqtBLw4kVh9hIFtdV6wszTqz3AheZrHaezIfy
WntElMbZOdY2n1IhK+tM01iYrmqi/5aLCyC2KyYaaGmbA4ZSJNUuy+YPb2dESA2B
hvUcpUpRfjYPMSoIIeVpJfNMZtaB6qTSfblk/g5np5uI+4lrYI2MKl4fkVjTTSmQ
fLvuk9cf5Py2jxCmlK3RrpSu/zQ+9Yr/jnK9/hcXm/Ij1T6L1YDo4XW1+w55MWCE
hDmO57bZcR+aRGBYe3yDwR4v6/mHTlc5atLIj/wRhHNlAGYwLWS6XSnbtOF6E+XX
rdGJac6hD9HasNHdxRmSVzqPYq9TR/AC5oZBLzjLNmNfpPt31k92k2KkzA77TB1v
jLp2amOGi+fciBxsg7P27ssmNr1OJkLqSM2j5tXq1EmsfmJMNgjEcZbfZjkcWprW
rnU5Dx7Vh9IcCfCfAu8y9AmjD/itnVOzcylfKrqnPj0ZCqHsJxBlpu944mYZ5nww
8uFNs0YHMdIoXc2tggN4qb0heRwomn6F90YwIPzRTqJgADT+BceiktJG/PDV8lQL
o0XqQdt4yWc549x02LQHzt95n+tP6WLNe4VviXYXuosIxtiarXceEG1URE6xBihL
bwwW5qR8bjhmzIBRTs9qc9I4/zgyzNy5wA63dUFxdpFnuXvkY3RmJXpR4gSEXXkx
Et8YRNdYjVG/mUcHvlS7uB9AizZNtovormcBq5fib7kWX4eqkEEvTdgjT9rnOQCD
5f3+MxgPKfM0UZkiPukVvnnLxnw5WIBdRVMqwjYMfrH1amtR4Jzf02FzkcaQHSTw
djpX4Wr0IrnQZmyR5MHESCyoU7OJsdhDFh3UWFvWYw1jNwT6UPfzRIvL8/rLXgjc
8nWNeMqcO+FAAAhQD3/34paByF96uMWpYHvaV3I/PcGm4VVHf/9pZoee8UBzzv7n
jkC2pWImF0ThjEpCTMLMsbmpgAPMRVUZxDKybjMOAHEIzRT1qdL/Kf3UI8PfIkuW
zJ3EHklGUrfEzr64skfxsHmRzz8p4RaNenRIjFGdplprATM0A/kEvkcjyEI8dZ+6
CtBl6AdOyHX11ad/ll03KRVbRYlWais+NB5iExqqBJ+Oyv5pXmx6pwZGk5U9hHzU
uAdluzkupbyU9O0pL0nWbILhK68jWlEQAZ8HeUIH1+hTPwss51f7s++isF0OfLxV
Nxm9oipiUpE1pgG8j9BUAQOLfRY1bm/A3kbrT3DlRcxSz/rBT05fXEoRRnSPMjjK
FsRdrOKi8l7CsGQn1SOJcmu7lTLjA+1i2jSLUnfoKU75vg/NLgv11XtZ/3Ob5sG5
w2A2FB3O5cWKO+B7dI3ASyeVYPUrmT4VGbEQGX2XWG/fNIGb6Ub2a3PHOY9ULkLf
EdJGQLiJL+FT5hNTKz7JC1X/6dgVeqqiBA3J2InhOBb69V6sz5gFV/q4bQKZrSgF
hj15A5pVW1OpMWv9MI46Pxi57Keio8wvICdVUBSV+cX6Ur1GEGhEmYNrT+p/cObT
W+I4cijA+9usDjZsv4hHwEALV6QjvFbIKxx+wBZ+GVwzBfZZ0E/5shJOgYw9z11w
deLBbm1hd1t0zmWoWvNwNyJprGyhUfDGJjJfHOO02vl9r4qiXhT2h8cLrKVDoGFR
1mJV8i39AuzXAWQ90wouAWLvv6bx057wRC8kkIanuxaEWZAQRkra9koCtPUYs1Gs
ArBpzjVIPtPcgg3Dpxubp1nv4lqqeGjCgPl6O6TcA7WTTN58D7v7YheohV0ES0hd
JLP+bow2lU2WxSV142u1VYy9bnfKE1+Amv7Dp7HrRO/H2oN4ij3ddD8VuS39JFIJ
39zJZR8xMocIZvmp/trVgp/IxeUUzfqMB1W6YIO2Ri+7uzHo7L7r8RMtilJWtLV7
e+T4jfnkswHd1mb8gtvT1dhc40VZqKG7pqyuSmZPK0A=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gr96dDK10Ot7xxUgs5lZWdYkb+FYLlCczH6gZ+cpzV0xA5+b2GmPEW34/NxALLTm
ewcOo4MOlTQ9ek9kvCdmAjHehyCQ/jvPTeRKeh2XKTEBeeJY2yvNM9+88pdQlpXm
pwHh8hcF0iU5AVjOf4IfWWT4faOpkMG+jq822keyNAeKRjS3fzJ+mvCBlDETCduD
LjOWkdPSLjMjEALkRA9HfJ6olCthFFPb9agrEe45OZRlfqiUhkRr9nF5gh2mpAn9
E3HvdMxkTLNBxj5l3/gvWgoXfOHD73qH2lYGO8PvhBSJ4VVQdtlLgW2RtnQcDJXP
9PUWeL8D5fk6QwdpCo21CQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5904 )
`pragma protect data_block
E+noE2zKVrlat+wnnq6S4jYSqj960aBElJK2M7RikTq5vEXGQYQ0rSwu2+OloXi5
SG6P3D2Wmph+R0C8YW8Lx+EmnIEQRXMxGj5ebSo6S4p+DATtntiUdmf2++INnHs7
BlJsPxBg9tujPjJ+5FIlu3/JOyiWc2DJI+amZ9ShdIY7Ll06P1Jaq96n3UHrj4X2
7Kgr4+rjKh9KNyTxkmRpQIP0YyIEck07rNHxduNGFdLS8DK0Pi5hoHQr7RR0VIfY
gzTQAyM2lp3GDTinUrIsOYDFrIFaw38A8ls8wyB0v/gpJH3OCS+vzD01/xJKXQOE
XBAAzZfnYjBGu1LMW1UPX4HzoJhUS0EpJ3bvwXdR61W5XWarpsLITAh9GmH5xMom
rxlC7v+wpvHK9PFojQR1PLWc1fPOQFAe2ScJctC+TvjhDcKXCwslQLCu5/qtWV/T
55FgqurfLcaydSZ4rKwQB2AcFa223ta/NRe45dFDmfDmn/L1W/OFVbtq37amw3Ph
f8n6ebl7jqOIS7H4XHoMfCxzrpS3fO53ulWndeXDgFYvfPHQl3O128tufKkiMMCB
diJOtXbhlZeibJU7oot8vqxXve+QoA2K88TK7Y/nl3FwHDRyE4H9stgtQ6WsmR0e
St+y2Vr4CesMxtcDadtfgUJK+lZvZYWNXlQZ+FRPlD0/x4oxDXB/SXSYLauckxy3
sZ5ao+WyO6cQMdphTMe38vDlReZZgge2lScLcnaqR8SUw94+d/+FlXXOaXTEsWHj
tPlVeyzD76pH058XfAVxNNeeQrnX0sZoO8iFMuv85ynKODjBeaUYRndVl4UyEgpH
6kycTODdUrwgZ5uV40uNFunHaZ9S8ZIcBdXLF8Z3aOXLzMK2+CEQIaW3n2/WQnlp
qPwamQeBFfiUEDOnqhW3uW/uSfKyYA7CaXJgD1yNw+N4OjWHITYo4E/KJ0ufAirp
GQ9VGHflUu1t1FqYMJyT1I7hWLByUskhAVSyCTzyyWKMzZqGjuXI5UASZvjKqqEz
PwLgRZL80+HnBSbR/KBlkCQbafj7PnXTKU4nYE8gQixDbeRPiknR3Xl7YveWsvPY
JayT+/S0NO1+XvkeYWpiLv+HRVSnuNU54RejjqwzT7dBmJOohk9emGU9PVLWSeCf
gX7cAV/paskJDrmSDMsbEYQksOfdZo/Ya5rN68RmQ9Huk2m75AuTbVIE45d1Z3/f
GyWPW3kN8BazqG8Ndfk0OOe5DYyg0D7mjaGNFFLV+5hhWe5tNl+0xSAH+A6miK7K
elut0NspwNckQt6IkClsT/bIvdOI3IoI57GNkoeihjXS6/MX6TFJI2IVIxMac10h
uUUCcxCm6RpIOnFmhAfFlu3L28SvIz7Li+r9s2j370VVlzNWP17pvT39eJAqlnRI
fgzjBhgWuD7s7ao9JGI3sdJUSTAY1PQIQ6Yb6+wiT6AUWKRbjdas2+/KlE13Fu9A
hiSk5LBjIiCCpR1HmXWf39A5VZJjmPGJEKRlzSx8fBqr0hnYorwfUWQSC+9bHHhi
iK8mk0wWlJi8IkCMM8CxoCXXKk8YOLF/7y+v21cliCORfPiMtaArwrdxVTYAdE4K
SOIo/bLul7fK5J+vKqg5Qcfsh4AZVBxWticLiGs49YONkA9sFfWipd4IMaR7J8M0
ov+YPI/KqFHU3duu9LBu3jR+FvrB65xFfirhmigsineeVqFrPPvWWboM86vPRAHf
0DyxcLink82XrurKWkFk4IlDgSkNg593Ji44PboFsKMbitBHR46sc4Toi8KWXzKH
EUrrGvslw5IGOzp9KAK0zNruh80/I9yLeL66esVsfB38qlj8FF96w45xrqnAYtr4
dh4/LPJVTmTNEoDDmjpuVD6TQ15C8/cZhhyLbiKgXI2OXrfdqlYKNBZkJv86fNoL
UOSlAzjiHp0rJk6R5vkbz0ynMl3gcX6nqTutez34rrCBwRYviwxKIGyZs7gyz23x
D7NrOWDzhflc0iv84hVBrSotnP1P6aEbbymzPoPfvo52Bfg6bt/HqYRMZVo+S5cz
zcEawrO9POqtqStoCwXOcxwkYUmg80ylUpFo9nD2SpiwjmLmqyiGwhSBHg0Hg0Zx
wJUxgRpx1byrtk4UZQcO1JaRKrqUAjbqJ5edfG5EOxbAdixnrK2N9WwJr/grkIL+
YLfVDo51L7R3wMOmRWTqORte1hI5rlJyIf9etsom5uEXE/jV4ArJ8g1VT9sMQOhv
SGba/O5NZwZ1l3j1v1KZXptXXOkyklqh+1MmIttviXd+u+7sIuTfNVBAiuKptP6P
OgjcFUNNZXtlvw2E2rqchfLTYgq0hytxWDIAzx5BvlZlN+vVSK2/9qaH03+dEIKj
QrHHPKw6GWYfX75wwsqEgDfLKNd+1jlSTdj5itxlGxNxloOyPrR/aVGp5290UMHA
wssIRAUofK+wzUSiUaRTzZmCYvCxWi4nH6tVYkJ0vjgLAEizzXl3xjbsQp9XKVod
E2CGh97sqw8hX6A/0tXRO25HuBX8KUS8gkh7hFDrWwbW5SJglTJkOqLp++D7D7rd
SPBsogiCEvMJnsgQfGDKuGlKH3VHAvmyU1JYawo6jB1dBTsUKsKP1DSFdKgxW211
sTjKv6I7KjvD7/sWowLLF5uTH9+g7BeIO4Yj7Ap4hH+F1MeHgfEziHc6AEm/eir5
Twr3L+4I/jcksEQLDMvXeb9/Y2Zfyzl3ZS8j9v49dhCyR1sVUKxgt9/awoKhIRMN
gvFVKrPKZ04OpauaIz76DR09C9AHbCuc300O87Udmhl6/AfH81UFwUFnMaqF6ZHp
D/4XvKzyyIaolmRvY/xBuflLxPbuSUnokBpAN/Iw00r1/xzHgvk56STK12rQnhaw
9c781npOTdb/QxzQwogN9g1d09fzu7s6wY5zyu42fG7Y9Zq1wKkj39xpaqlAHp6S
YHZeGO5Grxnv0AobmsJBTc2IePhAJ/bir0ff10/8/FkaYAl1VqTM98UR/7YUGwqQ
ThVlipdhE0V11Qg3skAzPOQtwdo3W/7v7ty8SirFM2yxZDLEysPn4hiTrpMATgq7
DlfWtAR2E/9HlzdhhkUttKAscn0inIczcCYVFF+oYDnrdP3F8ayqPtoBg3VJ8DI6
BdBUZ/jwWLjW6ZDDO4R+W/Gg6pIr0YlZUELWeHuUaxLnnAp2sI8CitirEcup3EZz
SPUtg1KlmLRvFmEvOfdXlamgt6Aw6lTxMLdY6AAK+xLBGmb2jBe5Ig9XyN285DSD
OzVjyn+2jcWdSv8UjXkFgj6EpmuRg5uVbNMkgw51hq35r8DzVTE+kr5dU3m0kV6u
YiyWeI3aGjR0/f05syVWBNKnEdSAgk27SWbFSJmy5B4/g4wVsDioYkP/6OSFm2zk
UQGtsKCV/PSGaHCdSaPq9WhCTUhviyLpGfvGFKUgdnwJVBcpKa71QLOgeVeSozwe
vDXyzXmD8Ar47qcPMsLt/qCNgbuRgDXtJoPApH9l/ebPDdeKMPT1pJ/V1kwQ/YJA
t5SrHeQJZMkbwBhwdr1uOHSX/KoOr5K6iFTrwNCWVjOmRAgSNN4Mm1v7pGLQSuEd
WC74XwjsJ/2hy3czjlM84RFB1A1WQCYrzprV0UuS90+du/GkqKjOJ94cxA7BNrzN
L7O1+7VfRgSpdRghqaFpmMsq16AGJYjGDJmjp61+eMCDncoB6JzRFEmTZDIAgsqv
5ow7nTXc06QJ0owTIbCQ/GG9ZHBgc+trnFar+E0sxyQYcgYi+5oFLKR/eKRDHHBG
KZ/E5+HUWxC+dF/5qY24K+IFc4ae/Zuao/Gn16Kwgc6SveBh1kJit2r2svvY8UZZ
JmCeD+pA+YcI2t1iHNb7o17yRoiDQbMSUqxW7Q4BGYCfhDsQiagq4t5zyCZLVKvv
xa5axtlz/HyCrM+RH96rptuD/z/Z5g8GnhWzcEV7xOul83b0UhZbKQAuK1LGxNRj
fxAONOKGtgG2c3fR3wce3489Oz0cAaRHXDlLImdl5PiuOKZknD7hDvCETKL8cKUH
YJ3aoGo9VH2RlG0h3/EOliZpb31BXe83nybKVs9ufN0O30lc5y51y45eiWZF+Zdq
Q+JBge34fczolbdFGuARvZqcif1/mzNOx/fZNX6V1uHUQ+mj1ddfj/KQ8sdUYUgo
7UNdC2dO4EnWJlRkyNBMPvoE1FG3tyraaq14iRlEAPd/qQzKzqrNalggGUv2MuKT
r2WelDvA7IT/PXjW4Dti9PGhJ3ozXuaqL3i+NAHHF+IzwWpqH+DyFfKR2PwKDZxB
h2C2t95qCWtm/F+OZ+9bMhC1gjY1Bh4tWGeZR+26YVONlPdkujaLJtxUXpKCTxCV
1iiVnd0cjDDCgBW6/ILBsSgZzk89uKdUu3oTTVaaZE1hdH7u8UVn+K3xnlDO+uih
b/QX/RFUvevsrco+2evT3OIULoQN2Hmwyg2U8CXQe1kVSDMFsuObU6Uh8BL8iuio
XYJfS9dKMk5qlMq8fLONDpWSj16AESkTf11BdZQ9D/LG+VYrdWTjz6zUe8QocRDc
yblPL+dzgIQR1Phjq27Fw75QZELX0Cs2metZEKIfMEV+m4/5s+AcqciN2wz8vlTP
22+qNv+WjMc4aK08h88NULFaYxadAoIg9bUay3dVsSbsAL1GDMpRG1BnQJBCz6Ai
o68UIYm0wwg7M9yJAtYew8MFLoA/84TA2CfMxoQMP6TgPIo5i7reb+gnYCAFwDjG
wyqiFJVN0D5nCGqTyjwo1lw+3CdVvqXzjoA9197NV81dWjcRvtV3/IEpe6XuIynG
fl5QB7ioGAazKDWBQWLpkEw9ucV1GGGn8f+SgN/RdpeUlLJfFtfMS9ADRPCK9Hlf
bwF0TdCzT4yBnChDCISYbX/RqWysk39kRNPfCec3TWqYkC0ELZI6aT69xaTq07ej
bmA/KJdl9Nc+KmyYFJFLXwW45U2RLGVS51q7MhrTSDnU+JUJ0W053uLlAKKtkoOT
jKK5914ofetdANG5Y2jvEquzrAS5hvXsfoaQ6Rk86xmpY6+onbIuSoK6XW7Zfwp5
wYujP/vqsTDZjX1l5g5VI+fXrsOIVY6h8GD4Jqei5oafnxgi88aPx+/A4RF4lSFT
wOyZUvK8N6Axe3qIddJeZNqVjX8LIZAEmrm6H3eDf2xuJDMjmvTh4h5hHUbB95Ui
QCo0pwsUEABWEqeKfDjB8DsdjWTOjtGfoTW9rgSvdqS8PEDEbDwmmj0/9Rvv882y
ENADeTAbMfVZEYDvkTV3UflK9/eyMiSiLCPUVTwd8KNw9bucjjqk/SuP1Xgu6PA6
bbdh3s+sMQMnvmuxpiFTJmOOiGRNfpoW8UFeJt32Gf5EIgHGUzG9+/BuoETaphI/
fAOlLehXxdeNicPituMVwcpdkBACpSvTAYLEWyt/p4rH5twcoc4q/NVVodnIOXHl
stuRPoa+CDHMFlXp9u/7HG6TwvnGqtvJJJi19pJyCpWyecYrzyXu1PAGa5eV9ZIt
a1ACr1w9dwy6Ykbp8GbCVaKqBzRTHPF1K7S5VcTbOpXir559fW92eSwgD+cisNni
w5E2/M0Lf1nAHnDO2X6a5BrwsnHkcTbWEE3injiSwbtvpMuqFovLKhrRbkQ4qIqC
PFiL7qV0ark89Xk/KCtNt93zn4QQC/3bzHNug77lwv4QxEf3l8Dkh06NlNyN7GHi
3P+1GBH5zVSfXbOoWphy/+LXP9M8V7oLCwEeQJkIlZW+SauKTlOSfIlbYsHPtxeb
shmBagabOK8uiZHh5uwhha4hlAyZytVR4j0Th3m4icLgAE2I/z9oOvkXxpQ+ECX9
23A7aKTjAzOaZVFIrk7MNnSHuLiK61Pg46gqxSjB9kMbp12KyZHJzdy+sGn4Yl2y
mthGTUvhPbKdhCqMzNnON/dOPyPwb3l4cdO4CBgnR7gVQthvHFJOhlkfTKJDpk8l
g9h+9T3OPKa5Oia4cippz71QIyYjC4xaAXJdTh2IkTYFTDzjJ2GyUk55W2i7C2+V
OgN+jm4Z946Qawa59/BMyIPJrGMXr/W5XKV1I28Ssf4N/3MBHb88kGsq7kFbg2F1
vVfMdNlv3mSjwsJ9IVpKpnOuGjqYGuVNLA/9tvjL64AEw8s/M0lMsryI6XsZvjgm
bAl7WHPJ3ZDjoq/tf9JvjDJ5NWSLNRJ4+EqMvJRTsBf3F2nhQ4B8L0tRorwQaYLn
2T9hWqnihHeHHB33YZCYCRuEnBJpfifgag2mS/W2TkR4dUT4aSOpp3D2Nx/HPqUi
kXlZDphDQEP+KOTgTAvyYI4hqSa+slzgpYYv65A2sS6xEXkq17Co9885Ya32Mr2D
eRwwyhPnc6dun1eSPPUgpRMjkgNpEmwLxdTfG3dtH3T+HI936yV7VmMh6Hob28iW
9yJMO79tesksWJjgBPmTv2HKqxJRvFvMatYF+PZBGcpyCsIo/9Bt7Jkl0peEWEN+
32XeuUnfjA915Vz5Pu3j4Cb0sKNoMUt6tV16+kM74zs4yIq6lzkvyG4WEcLIAOg8
7E8OBxPpXz1kiIv0xBpk+0/n87LEU0JGv4pBztuYw5LiQcvfE+09HzT0T87ikuYV
uWq6lF9R0U5vsBzOrQF+JZpnZTlscG7krERdKccw+QIL+lRLRiVYU4ndsBPv6+fM
+PFfN4Vfq1K1dg79EWEUSuVFqNcw3/qO9QfTG0Tw7k5Mr4eETYZynh0WjTxvmMle
Ae2gjwX+5FVdUSF6ImrxD0afp7PTvG2IoiIv4CBXeSNSCKIYoEi0mgw8akyRCW9/
K/uLuyoLtJZEoi8usVvNrziA21mzKn6wP00UYol3h1s2AUV+SeICSKIZ+U9GWAs8
ufwBmHHG5b4CvS/UgE7vWP5SSglU33c7ZBAkptJCanz3ccjxsECqt4bDNVXfNNT2
vkENpJ5hjRyJ8knN+7Pznuo/raj06eExnKVaU/qgWyOoitBMGqeyk1J8eN8iaSD9
ZdXjZYUA1NJPzNYM2kUD6b3On42pMDxD0yhMkQAciQpThZXhqznTNSavTx0Plyq5
M3vZgBen+KM5Uf3bmOY0L6rBPBMq2OXS4FPUXAIMonijUMxumS6GIl4keyGNu5V3
l72f25Jp1xUY9mU++1zI/LPGyQeuT7gJDaI8gqJTWARJzUZwNiVt2ZCc8xE1RG9v
GUvrTnCJeu+Ci8uzM1HnWQhxL1ksF8Uh9SF4mV9LT1kTXG+qBF2fiKmYgySGXKm9
J8bOFMoWKo3kmWpBqUQPaH5VXm2pSJQVM8ZMo+OUfrO10oWRTwbi+wHmOCAkEsJi
r3Mnzd9TBDolxPuNIBIoXsYcmBc0eiLHuUe+6RCRK0pMN5r4IbwBkHlF1nToehwR
OH2+Dy0rVNpIMcDSZTRM5wzqDX1TPTmMjPypiq8LqwFDwwP877inR1JbU6zkip5W
LG9wr1PIgbRzAjEXxghUl8QwK7YdDJLtC8ZrgLbj6ExlXvE/1EhmcxlyHuJTpStB
FKA7wQ0MAiOFbBZ2ycCObLm8ex8JhdLPKpnWay9+zf3Ci+ozHg2GijRY4VnHUlXs
jC7CGwpDeARXy3jfUQlruB7JJq2O9+LQjqlgUs8gX4sOLCQTUKZ3kIHoJj/hqzSF
9gEWmR1NyluRvfSuzAjIJiXh3ozaIorOX0xXkDGGE5WkO75OoXuDPLSrL79kGgrY
ToeXnT22RcM3yYHQW7EM7hUYN6bpj86ZysSvQMfcyU2+3qVJvLrtG3QWhWDS9Rxm
FZL9KAxRgb0uTM+DFgPY1NGIoQ3XullXwdnwwI6oS8Kapd8Qw3SpXe9Ldqb9yTSC
EZkPoQ+EM2qBavn79aFlQH9VE6eFrZofdRdqQ461S06VunQIYxXXuKD9xWpL1Umc
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
OlJa6uBve1fFeDp4sFTlyctKDuuwNGsKuUBybmPyEU3SyqDscySoST5zZ55iuv39
CYAeTXycoTnAMGAIdN79QMhIRqDGDyVsE7TlXT8IGHdiRKn0rHucJXh1AaudGfek
fGYDcU1I0i5SHpoAu7Sjg3YLeNO+/x5mycnXitWQM8GsiqPBo8X6pXaP9koeitGE
1s/J84T2WlEb3srGIuqtsM9YGp13QggHTpsNs3gOEEKsYgKZN1cPq/hqwkzrqWqS
F6wn91FHhY5YRJqRz7I4ZieURtfxIexeXDMudFLkhssVUqLTi2T/e/qnIXzC0C8k
Sx3rR7rAULOi+ljIQt+Xrg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7648 )
`pragma protect data_block
dajm4oKvsI0Pr8bgbtbrr/Y+ccYYqqPItFYOH2yVOyFqfF+4ddGogWKj/mMj1K8u
hO5cD/o8eda5K6W5tCSO+nWddrMAab+FelUe0yGbHvEjc8C5NGxfRPMIrvm/IuGF
CcT+9CPVpc8GaJHm8GEeimhlhEVSqTEuJfiKLezvV5LvicVqOyoX1kc8EsqVf6Kh
Sh4tvDNGebt0I77kBKXDLVR8r0ltcRFxte0I2vYHWNxbQmwiP31eQXIqgQSb29d7
Zsc/XJrJl1MvgoCkCkchdldhVkOgTGGNwaHtXbhpUlQVVYKfgkJtYGxvXcGfeDWT
jxds6Pk39UTApq8K8Z5sJubxuRYL7l8SgqTNDrp7D3XHwfRgIBkZQSrRcU++Bmx7
FsDcEaNScCOOOqBa5KuknSwrm7yO/ZbOUdJrX0hoMFwz1uW0Dk5sMe9Dgm3CODbR
wCy5l0/E6Q3fdABJ1Ai0/KAypbf7lun9k13D/4b2EBA5jCchAvHFxBRzj3c75dii
CoMX/UmfiwMtdWjzAgWq7Clf8vbkfOGUYRqd7YhbRhIJwQl8CIPube4YzPl4yrC0
altcgYtPzMhsjYthRkdsL6es+mxKm3zENVD/xHFDAKa4/TIP8wUaNhVvf3tnqL/T
gtgVkkyjqJCSfAcX2fuBJdP3xwXqENmeBiskwG+vNChnc9YjUgbpkRUzLGojm67J
NQVXRBfzo8Oc/cK5eznoAFBmsDnJOo9VM1c2LnDkYm4h6ijhOznwNF8KdDSnsOwz
nWZBcGf4NVbXV6zsS/+88j6TqKGpLoRKS8l9cjI9/UUqdYvuL11v0+mQgn3z7OtI
KPG9WdJocU9dAYM87WmSrWAjpXL2mQEP7kLe0/n+TOi8s9G4HkjOh+vZemj04vd6
aJoQb3j89aZs0VxEtT3SYdfbwcNj+TVZcY+44OE3EMm7IvR0yje8dg6o0vPwtmWx
0q8HxtfsLe6P2n4LyMipEqYn24iCtt/nF5KQwFGN4Qdp4A/OGPO+ERb1Fm0ZsBbP
cl7dk5uaGiQ31zprrlq3ncAJPTbB2t4ok9Xvb04rgHKKf6m9NUq2kn9EYAjnX3aQ
uQS/jekN2FdJPqvHxShLlrD8B2jasVq5azTf74IYHfi+I17HMyCeaxZVZvWs9UjT
3JWGAs9utOk43itgiye3f6Uz+6RlfM+E7B0hGr+g9WJcm1LJOK1Kq5t40gkmNpcN
5CUhHupB0MGz5rPCaO/ISwNeP1ou9+t9eDj3US9kSdtnf/gvQfYngXWHExAAHDcp
8cN+J0TuxWYyfzee/+UcB0aU+KhVTJ/ihEM4nkDfUxUDikP9SRmWL8tDmizgqJP0
CA8G50R/DaoQRLa/8Qnmo2nRC++NfkvkBO5qldfRejPJZl6kM8VMaTijgVoOweFF
AYQ2bLciaxX7ViQO8t8udYuY2uYktsA+cSMgYxi14WwBcw3ETzn6Z6kp4BYqyLeJ
86j5gqY4yh9ljBX/KBJI4ndxCWGX9teaQGtY9vdbfIa1BJ7lkkxnK6miA3+WM07V
uOpHCtRbtvKMlfqVSSEm0VPnj2bdkoRJY5V9MQGlX+Ofv8TEFPESmJjFHs1+i4B4
PLvHHkR86AtHQLkC0tvMLzb+8vj4j3ajw29F9BjbpntbQYP+XCV/PlQ0r0TbFdOc
g9Fd4k9CQKJ6YG7eNM0iDmmgPiOGSSCcPRHdGatFIg5dtXyCbJYTr8kVxB2t9ClG
EcuDcwRbGwd3tQOgCyNN8EkHnybbsE53EyzXklOUmavYzwMfQII6vfPbabv1BeZh
0jbCSOEip+aPRJ9iKEOz5jyOD5t0DS9knsnhhT1v3sk4qYreAI3GY+WxOIeLxXXK
Xzx/TbRkjrzQRrC9O0ArUx8kaQqyXD1gnco2ReARCmanCUefEhAZrb8bRZccEe64
2m07Yaqm2S9gYksKrPD2qZiVOHbxwEas81u7UaWTsvKLCtblxOGKHK7iMvehRsKj
bCVxUfr+MMq9TvoBJTBO9wl69/VdHvOJGoKVN+fVqV45r0nykDRPAVwR4+TlxixX
yuaQmr7l5CT0BoLDwVokddNn6Nf+ORiK74MgaxTuFemQxb8DSxDhcQ5cHuWzkUNe
0v7IVMfJeanIzzgs7bZnAQItunr7pnTS8zADryWb6Ok7WNKXlBl38PrTwDkHaDiP
hLOqbKwdTSQHFGCtY1SbboXkojNNsZ2K/lSGNvfOx0FhbzomHf0HZsZI6DyKbinz
NLCRJGXsPva0LF6zIUQioTTdsp4z8VdBmxmkIAewHDRF2BhhkZztoBCXE59gECKx
ZKvi41iFTz2d5GDinDzh1iUOxGWFVCDCnY8Yuur0Gjv27She8j/3Lz3twOL8HMJm
/XTVeNPjeK/CM+Bk5leh1eH0ULtr7dRsWZhYXuQS4F6VEmI1uXC42ye9Cm1umSyD
2oOiNzTSixKXRpP1jvSqZeA3NBpXW9G1UUFi0+ZnOJ+IpcAXm0Q9om7l2k1VmSp5
bs/vxtnP9Hk+z5Hkvkr6yPeVzu5G/4s7GKNC1NDy5KJPxohWXE2v8YQ8bBrMkf1B
N9OMgYeAQkjlxahJq+5WO2ZLqSELJ21ga0oSIG+k92hDNIBtmz/74QR9ADxT3M8L
BHk0Qu64bw/5bOdvzsE7SFSlseawDvlhHnDb6RlDFE3uSOQwGJeOQCFNckYbdf8V
2PV1m7sReTvq0WXTOuaTtJ4rQDYxCI8wLuUom8MKkC0V7JOAzEDufytJU6nC8mv3
nzH6iJHWYz04vREAhBrOysDsIzH76AHCyTCl4V05z/IEeNaYMmeHb/XXy+apa33N
S5rFaWBWzDoqUYLwxCkbXTPOE/kEbNVwQPf4XWK203TIdgcvm5ONCHmGLejEctV5
Fl3VW7ZQNsQJzLofUWOoan0RQ6/NTIuMdMiSQG+QM+0fZlvCVlRPyLU4o+TY1CFp
ysOUWg8KecTs8N5CYBmuDbvHFCBbKPBRrwUtOD6gVAfLWcX89+o6wVC3/81Hzi6l
T0AVbVowp4RDGxj6fKrs8eJC8IscTjqQ7BlEnMTu6sgi/hgS8BccQbW3E1KXilie
7NqU1g3yQ4BbGyKNd2BkgDOtLpZVjU/hmLsnQ/TREzS8uWFdArHC/e8mCMklqD1A
fKCQxYwdDGOHKd9HUMh+J1z7sEa28c1Nmlsi5JD1dmthI/OL9lkMbtr2HCu8ib7V
i+b3KM3GcZwPlfmgKKhz45TCQcUPF2O5d1PEgcMkbg/hIxu/YvfvhVYt4oVt4DRO
OqroZD5sMdgnNPb36jEXhCondPbbP/fIhVEHjLI11UckF3PQuwISYNPC8HC5VMQR
Vnt0gEBAmq/0j7NHoehExZZhe+WUiOjN5AuFbnq1ArMKH/o4rMvTJCGdvLfxnBzg
uCjdeVjp/IqV95XSOdLAYr7xoMv/3lksWpUDt/Qmxk9s3lcOGp505cl+65R9e0//
nAGDDcn9wW6ALzHLl8Je4mhTNiloKcQdkkNY848c/tawBVy/Az/UgsisY9vsec9X
MT1ywk4MF6SnW9ev3BSXkJXdNlFkN8Tf8T9CXb+92OzB2F+FI7d6fgwVzG3WpjcS
fvX+2kd/wTJaUHldpNxL3FU3jXA7VFUzUGs0on+RYkyAyDQD4N7TGCnHIf/2xeWb
yJGNr84+erZjgtR9hjVKTLyrt2Vw/YIq2CXJ2Jeg7eLQmYLJoY21juIqK8VKpByP
pWSLdYVzcYBrcDEqhCIkcwVQkbAaeAk8jUZgS+DAfzw7tpJ3rKm4Irjq8FtBELy3
FAJomjnb+K++yVTnir51s87XflgEoFfthx0aoVlh6Gr/+pSKAyLDRcoh6YXjVJvd
icvjbubwN470OxcwODpv+u7BX70RTnvrFI7A0fB6rG1AcgkGj+F/GYJ2wvm60JxM
4dg4vbCxrZMmlXR6khCU2jcWO05e386MbPMI4QxliHAkBdpm3lLxyxTwYxeEzBFc
QYgGpOAfUV/BnoU3w87MZ7TLhZUurecJmlh3EM0s3aQdyCN78XRuVZ5zwc89jLAn
lxhztI0w5+Tpw81H4qecqxSELq0b2PxOXcWYLbqTPPJ6RjXY8Co9QApBGUWqdyrX
xLZz+ABjlYs9p668KaipD4lZrQBB06lmko5MWJbZPXGk/92LoRBlqEnFzwz9i8VZ
/FRHAu9OETYS2040t3ZGMgH5yur/37RGNH6z1IimrSnjXKMW1TIu/iGief6hVXPP
3HDNxt51uFHI+oY0UcYEdruFccrP1lsn5u+rfQg38BxEy1CbMyZkwizjuhl9oa3X
OUzRGGtWXeU+ZfOnVkp6T4MhK/bgrWupwa6guYtjP3P9Sd8lz+qjKpDm7+FJNe7l
zu3KJaoPtPfjSwb36gziJz0vpojMUHeRJQWv5dohJubYLv6hdtMy6xKJgOQtz9qA
aCMB5eU52MKmfkF8OtxWHJ0objEP9FTrSbvIh7J9nxokhokaerF25gj+mh9cy/xC
Qjlilt797vipBZlmzk45c4jkjOuEbgkYG9Cy6SgkLm5cnhKEjxWvjCLEHtBvEMl1
nGwpJ3U0MNeZefsrzeoJ3by8WwC+yQ3epNY1FBK+S+crYt2CtZlUNcFBCqvcvydv
mqGWedh1L4Qz64v6ouRvnQUNUzYDb++pTUoid/OmQXu7kB0PqTm3ed+wyQGsAe3v
en1ZHPm3zbiMRVjTuQwp1/0k2k3YjTKfFYypxgRHC+yTHMUQbykD0w8TxAAj0kVz
d95mvHJ+BWiJeDGnOUztm25moRNrQLBlWaRdU7SQgA8ERZM6XXtM569bY2RFDrC4
RL+YGSRjCFl4NotBXoLmOtbgNtjl5EMiRJyjb8e52BptxMz2EjZocXrQiYC8GsF1
MPpj9/OjsJhDEwsMCF5FxJ7KFTZxfHBuqRKAZvWtt1cej6d6mK+eHzKb95jHfxD/
3VaNb6R4niTRpZYWwlI3LNFqeanS8bK6Nqvwn2nNF2zWhM/V5S/pdOrn46UIpz8y
ull/dCo+vrC66oy68ORUk+YiKPdv+7gM7/UShcAo5kS50ZFgJDD3i5ziSBg3n8lw
p50wDPjpj/8mpqKxyArgvIUpYUuQelPB9Gqp4bl8QzMpJCE4u3BOvXWl/uWdC55T
6WT7HqCO7H92PivtOG6zXpWsFZ6Kp/z5se0dZfRHQ2llcg3s2SmQAYtt3ywj8ci+
c+E4/1/dLOatCOkM7OQRbln9O6qIShf2c/Sb/VPKuHeF9GpohJoLHDIVqv7YVSGb
kQ8fDZ9ECo6dIuR/Bd1VEH2/7eLPXoIisim4EZonZdUm/TZCqMi8duniqnhf7zNk
VETxX5ABbE+zRnYMy3OR2kU7kl5wR3i9+Zf8wE2QgwmzzLz5HsCEoHVBd/sACv2/
1YLC+W9+f3KMj5hPNqFzpiT2WRFnGWHLH8lVLBQ0RqDYPDr1GhwifkexbaczAP4p
cuR73Qcg+p9wkGoamy5WD3s1+ZKBGbLv4fX58wMcPKaS4uOovfBEJW+MZX3L4T04
h+QhAQu5n6yaeDKFohNs5UgfLfrCiVIzQyJhoygC9yjol4KNgpvvtqeO6OfGqL06
QyUThH7gz+1MzonClF1aWnBlYuhQZBFHIBMcgHTiBOoqgoxcUbCKNL96ZqdXcvrx
GxQ+avM+EPksykTm7AZnNiiC4Q7z2M5UQFAUw/9tPLk9M4zALuWWR164ogSUTiVA
+i7zs9bep6iQC6vs9raLN1WRK7PO0Sf3R1R5Eva5f918Q9pDa24pPF0koc0wO2Lv
kkToMW2sOnbtwO25DPoGU3yPsEoM8JfGkaklaWCAbxdmWbWvkrKpAa5yx2VqiUOk
Aqaq3J8XidTS8PhWTj8B0mlesQtVJLPcNCmP3KDKUzhR3E4MpnbW0lOKqSY/0ajs
vJv+uTKoyIwWo3bXhsLD6nzzCQmBlFMpIRBeEt8A8qzUKwIejGT7kGEl4jEfJiaN
a/kNujNCf5yU6RuGyLCLNbWnSsZr8X8OUBNSQJf538y7Q+EROfqFK4xiBsaJWGIR
U2bKdnHRs8Kyz/dEPEZH0Wm06kXYNx3Fr2CBtSjOm84jmSAdjRxvCBhPk2dnEhXf
35GyvZOa0yCNW/7IJdhlTK1XIaf7kDFakDrtJuVLJpngC8qE0VM59rXaoMxzX2QY
yF2RxMTvUnX3N6GWupI+9nOtsImEoVmr6YE4oaUNQCZ+e17vwy7Zv0vEYk1hmwxG
tDw9rXyE+CoqX+j/Cl5tfUZxAjj8zn7+VPvFdAJkrvIi1K68nWvIjOoS1G1k5qgb
hBoe8XFYEu6TWE9bAPdQGgqUD0+ORoAg1OQavH9Y+xXgrNFzslFzKIWg/BcOe28K
Ax2aSGsWdvwTUgivK4TZFpOfX0tGwWgfMdTSQB/c7Aaka8E2GcMQxc7Mo42qkv9R
WQ0hnGbLhMcURaDIyxd9AISiPz1hgM9FEk6UdSb23ppGnpxWc62zAvldKiZxT07F
c41kyUZJaN5vZ+hU6MY9i9IfYKxzNvVPcBxtTBKXIYxfSvEbgtdpKXJMcZzVRq1C
T7x6BSwuYfnD/38jY+ndLrhrcok3UpWpWCgxOLZtWC82iwfz733LA+TJdOMGKFf8
G9p2+VVNAl8mT9LEBp6Ox+DDYzoUA64uBfMUKZeO4/G0TygbAjEz+OitzELRBNI4
67qpa6nPgG3sgnmS2irjaquFoWz/eQ+SA2kRR77qWPbOb8PX1l+EYPAXvzUivwI5
rc7D9smoROd6YoKY8QQyzuMAL+Nnw52AdB4wR7hbGD7w5qBtQC/c+gppN/DBep96
tpr20wOn8A6odYP1RQ6wruVJ0pk2IJp3hPLNWBl+sLkHmF5QhqXF2AFUsiDm9MkA
Uoh6LwT5fciXDJLOm9AyfTbAGOwQwO+IpyGtZFRMFykVQ2bElgt8OPrhM6g0H0np
6X9o/9czUNiGlzftlKV+PTtm2frPE6W4yoKWh0nthxxtFQq1OzOrvcMmgDZIHQyV
QnTLDViWrJdNZFsolgmnuu+CAR79yvyBXTHJkQlBvHjk5yunAE1Re2e1vQFTcm17
Xcc60b+DcGf/Zn50g0ZPnWOYLYhYxpNG/moa+tsn03C8M3LPVrQjsN/JpSNAy6Rj
whsE4YgcXO/RewaAz66C2xvxYW486KRizQCzMHsMD31bQvmLaHtStEPrmOoej1mS
GeFpYWNVu6g6Iz8SJzvzPcAfY/pZsC7eeOmWM6tjOqxo+Vu5gyB2RkoJQidO9qoH
yOnSHX7ImK3uaxfx0xdVy2tzQ8YTxFvpGpvxz10xXNmOlhh346k2TM6YVcWvfBXe
dgAFj/cp3DeaXl551OqEH0trB8XTTfGBmQbUMN2VHKyJU/MfM0l9cdZAT4mQIW/r
o4vgBI4ctVqmXsBgrzbRZFhHuCSWIAyP12DW2eHe8o0u3KlcKpLXiRXFbarIBu0/
7e6KVS84JeMCeuqvWjcfovbKgHREpWxbhNE3a39uwBVaqHEry/WHdi+HLZ7YUjie
qsAEIarp5wEwkGSMPGNz9xE7fNO1S4cyM7AMQyGFUoIkkxvLmOFxy4DQl09AFvxD
/8byaciCBfOZShMuSsfzkISOWVI6GGD3YY+AjeyYzp0MP2aCL3BAWISScbswGS/o
6qIraEGzZck9ZRwKxq5p5ziioCSvxhM982HbjUFRIjlhW4rTUF+gkjylgNIUFsjF
/A3nkUTjT8gN4n5gvCYBX5hAHWUmabXMew7fYJoF3LgxwLToVmm0YDYm3hDX6ggJ
58Et1rxqQxpf7I4fqsjlji72SghGb36TCaXJXe8FFNVJ2M8JluoFYiOra2dgjkLw
mJEiFDJ85VC5Tz2yeUZjgDRVt1mURi6l0RwvnI80rysolYRU9Gp7S3hxiLrnAWQG
wIkikOhUCQhUuDzNGYhE3J0QeOTdb0x9JqTkFgLiS4L1pmNkwWMqw1BKoPl22G5x
akOCMGrn9ZENNxlApJCo2zVLPQdYT6c/kyX7d1Yp8E+Tzvk5t1VbXDV+6ZxAaR1M
IoyhO5djy2neMMgUjIiS0g3M9u5yCUUTe1qYtgDtBGplYfaT7dPf4IY0GOhb6pw5
HHhHB/XtLg0uDgYOt/XufUhJh6sZGLwTu/NbkWD9qhv7pMw7tro8G9zZxS2pqROs
3/s2YhxPvVsB2bXtQ2JdBUK4yzLFOapaYIwESo/XYHWwK0eCXUQNLjD8UIiYtqRA
Ixg2UJrJNedt0n2MDhn8dqWV1Ib+nDOd7xl3pmATifXjRAKqu9lYzJo/4x35IHNm
pW4dtSKWzbBe6+JVCNfLNz73xlKsDozHlkLxq32L+ouOQaB4bDhz6J082Tesu9B/
/MhM5MapMxF4RreY113ixZ9Ucmcp6iw9QMiYfh2pZZHPzfBi2DA4BEeXwhQpAtKT
GdMd2Kxk7FgQaWXXaVX2d1FHnTDBptLbAEguQqP50rweIwzolvpO0oUrxsrdR0dA
qYYQgCrChMBMCxaNsXnCpWuISZPD4xMUeT/lhCDlJCIijMbWcP9vkP60byc2dQSf
ok2IwAgXG1UHseNpUfihiL1F4oATy5LJF/JVLXEXhqCI+MgOjALQ9qAD6Y3q3fzN
5aoBzIIZSbCc3d6Q1jc4+R8/Ndg7MOY4fB5h6TUMHPN6JZFebMWBuhMZiJTt4lnN
8v94DSlIjzGBvZNJn8yaUFtInfjbG+QivVS0cePL4A/Prt8XC2Aj0uD+2KyV/dvq
NSGtSrww4p2iVIKdmH3gwwLq0xQ4PHyqzIjCEkg23ZZRJKAMUTQKcCzDCgj5jwiM
HK83hHSrKdvEcGD+dHiaMwVIeAUWapN2/pqymBv7TRz1nvA8oit4UrdCQ8S19RcM
eNzvdH1hzmbiBwiQJE5k2PuCdTdaJr1F+yacOAhEat1746/2sPTRGd58W3db8mkH
2gVnFHBV69ZXwfotpTioJjKvX5UkLbJB1SjQuP8WVvzVJJkLC6CN0Wbjss0dPuSM
1gERIP1ArZ5xVuJTtOuGtmd6w43xoxVtHkO7LK0HCpwCLfhm4KU6JRuSQ2KKkfaw
O/SJmM6pR51VfbEKK0dlCXwNUIAR0kaA7oZ0dKmfls2GihM9uLjsMIOK9iVet+Ei
YXjL34OLEHSF/A4aGw/pMiV7FJMSPBGTh/+Z2ABgYIUTi4LgGuQGzylThGQVd7Ct
/z1HbF6/StRuW8KOc/KewK7Wo3zMwR/1TiXUsn2BFB9wKUKTpyF+rlbPM9vXfPTm
Dkuvy3Y98z4zG5S21l4W44MYBzd03XVwMugB9trut7nJG4Hwv3W1nBupYHZajsME
6Hzxja4E/0ohmXUdfyCE/RC3gCXtGRF/CoQaMW8hmT+qDNaZvrm9Grq7zegX0A1z
WFcLClILKAs2jWWPBw1Sy/vO73vw67X/ANl2m1+0Bnt6abD1S+Nnmtty6sWT2BlR
o/GJyyw5tv39Gs71/14SOodFtzEC9M2fFlLD/B2Q/1h1sWjkZdx7dDHVQOctdwgE
LDtHJNv/GtkCt+W/glSk28QjXPNUI/XufFuA5LIMfc9e/XykGGnQuOk+yKhW0OgY
2Voc+0wGJbR+RRGug8PU0RURd9EMVC5ufY7blFYG2eKRtgLztwXBPG6hkAmw+uAS
HXLHulNNE+JLTtmgFModFGVMEeikyQMjul4yX0IAIMGUChi83X9tA8o9bOOKply+
kZTF3FyB+wjDTtTuT81zHPqWRP2epKcJaxY02hrNUfbj87u0i18G/+fpANLlerwL
9/Jw2HliGc3XRH9IZiEgdP9bwyry8hQL4fmcdSBlaKulCcw7lpLTRu8Jj5jn1Nbb
fB+VPmL5zYAFNozGUVnR2XbpONCiBh1mFcehLP2Kezc+MaSL7f/5pIqx7BVjstzp
ppLJDMSHSeBVd7qn6zQ63JQWW1paDYuszURCn7NkNDIwS33vH4gmG895vPdyHbCl
uBqEHw2dj/79l1fO8PxXGh/SE9/XxcKr5VqjlmNaAWUYrYLnPeMJfB7A5I3qmAV+
IxnJFwN6Sn4nqEaGrGUa32x2EhrNdrvCsxVlPFoJanw8cGPzgHPIAu9U0EIYEYkn
aKGxynL7akqP9sZOhoRvWdQ2f0aVcGa4HZIWwSsx6JfdG55X/MVX8zEotdfdhvhh
cWjziqNrRyOK8AtyDXdGl9TNEpnNJZQOh+tDT+W/eDVVwyy+iGuevwi2zFjq19DS
3b5rp8EszhCUz50Zd7m1jA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SqeSgKE6qiNGvHOk9wBu7XxrbNt2C/JwZk2y1nKwvdT3/PMRH/226Ge4V9F2El6O
7iDQrb1dS9GD8XEP1umwg+al55E2CdVW8O/qCUjtnXH00v/kicZylKP5iIImeaKe
4qD1KP3e28YbFoiBeQ+h5kXjxAHmJH/MYZRulW/g5Iv1ppndQTAehMLvfFr9fCUT
RXRjeYkQ+4S5JYZRfb4qmJeKFf9bKu+vFCu50G/lBmxiuI0H1m8TmONR8b2HXHHA
+m4/EwAl6Mf6k9DRwx8NWQvKijSVwlJNrbl5KABpcZN45UkK3Q+e+YYiPphpaFst
e2kfCKy2EJIeX8/sreGgdw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5632 )
`pragma protect data_block
L9ciDfliHHey1kYJRcLgxXQgVE0KZu1vQVPYAfyf/qqoGyFACyHdSEYiBCxDAvJL
4TCBV8mqRzRUxYRJDms6r+fRY92kEVxwGvfEF6L5e2wKiJ2YQIUdUnrvEkDpCWdF
LmGEu/ktpHaHSg9tKA1Dp8nJnsgDr2hKyVFWKRXMzC68JTNHhXDOcI58Zy3j/c3g
4qvhN95zkkxXTEFuloT/wuc9Mkn0fliI5beXTthQGlp64hDrQQ2G3V1QTe1z2NB7
GMjdvRC1/n+Z7UZJ5ceoFzQRf7xQXZk9t9B2vNEpmA2aNtl4gx/NbXx6rkJcBSV0
opUtvK8D+F6BnDe4peV2RsPLKyjC8luofKPl0cGNDVTIGfiRVus4FJUeudlbrhNo
TXfhm9z0s4r7VCPBvYqgBytSrLjIBzvZs+xpwfb06J2vkrYYQdBCqxc3SzCnS3j5
D7jio8yL8LT2mQijD75YgOpbM854LaAvWiviWRd+gAi5uY6ctIUDbEgf/Q3szaHt
/q2KH4ZUQYiwDPSTlK9LAPM8frO87XNWVp8rZ3mORhghmNsgl2HDbCKZWYFPMIEs
NoLIfUQ9utIGrrpNwcvfFZnTG/+PZ1nf0he3mOGtcxgPuBQueTCtfg8dIJ6CugDv
PAL82jaqPSgS8100Zx6V2x/3Kst8ZbXgNUvYtGX4TYdAaONVkY8a9GKpdAf5wWNA
LlBePX+wxQpvbfvdxB7DRW2QHHJ2TzcJl/95cy8NxHz9qU57zrIjltczaI21InGd
23chmKTxBpn1kWRQ9cFurqnDe/UQkChLM2x0fn0cpcuPZsw9KLYHxCFlJ0vHmjpY
mYwuC2P4K40l6bX5xdKNmDnb/V+++zeniZYexHcjfQcK5N3OevyM0uUylKE3t52/
5BPLsBpDfsIucKw9huFFZXl85wJfJnrzV8vFQuMOh8ZOu4rBnggvgf5nGu2jBQXs
jaXAzh4q4q0Bk6jDqtQpEzeW/h0S5G8N8Zol9FujkyNIwQm6YH3Wfg0jsiiW2EO0
VfgbbzF+wtG/HTPVWnS+kNhPYfVlLWfc6mLUPqgdozs4PLtH4MYThiT5hClcOPiS
sTJAWHeqRZkeXnTv30iLMN9vvKBQcY7/1zcrqQgty7YOXHUeMM14eLn8llfpaU45
1tZngtg9diZ4Ugu+ANH9IfZ/goZ2T0SFz3IEr2BeuuKijGpHncfI7A5cshg5dyUw
8wXBvvOf+DFjvu++Zc2MaToB3fyZXgs10YU6Ny9ghOZMP7wiFpm+tHH3PUloa9lZ
24F9WEFL/2DajHvZFvH8crFNxhNxILeDLG5ZBAsbZELdFWTOF3b63ntKglmdAQcM
+HCQ1B2HRuxmJkCQo5Y/9SBJSJTOAfpu+Y/lVHD49Sv7sBuyq0cRvvA/pV5yqSj9
4Pb3H3WzqCY3TvNwvkTViHxAINkIyZm3OSd+AoE/0P9p+uiFPt93R/Dq7OJWcVQs
D/GdfAXvSh4TXJEBdu9l/VdFIWXUWpJPhSqo9ywqX1OnJXg+Nu209nykO51xBfxg
HG4d0gAk9b5jEqm02yfgXXzZYZtTpbXBsvHe9aPP9UHQEPf7QbBwNqyU4OCYUQ/P
VxHtraoD+fL61/6+1HH8CCTK+biNF4V9eYyw0TcaUWe1voMTuSLtdjJX6sEGYU5X
ZMSNqYe6j7vRjNxoFw7QHLpg0FQ/Cp8sMayQJ/gSt9Hmh4wQDSzZTJ/nf+sT1O3Z
T9UZ7glOWetBA2UnEBEQsG5kjEgWTpz14fvFGPIFL4oZeGddsYGQx6ZUVHu8QtzL
z07x9QAhKxAoPhBdfS5zHldMSyujT4ergm9c+OZfF4Ug4CEn9coQkyB6cShW4WG/
o4eevqWeZaojYRqZQdXiBdNaVtFK2E6juRWmdJlQ1n4YTP7zofLL83vwdtaCY15u
/X93nkVJGiUjbtwy12aW6Q97c4XMp5VhsRLcsgPXJbm6PlNTnLVN9t972ECXV2/M
jBpt9afy/FcSUkgolWMJF+LgmC7zceDVr1WW4zbLVqrRxs2WRBfu0BrHdFTiZHq7
jCQLYHLdSETMtyrxzm5u8kf15k29ifkRY3+CAyiyDJdQi1sp4iCUjkwiti9h0wXV
dEgK0sPYRfep4YsqtoHjOCSAsbPt/m0qgXkpyGNEhiFH13onBQ9tJdkFxhgNqzQS
PkByrx5Ua2bRthB8Cc/K44AJfN4OPgyUvvQSZyzo0ufBfaxFVDJcNo8CdIIBfqCs
HhGoARL4eRC/6SR/DACMVaLMhzk5BAjc2U1u1jgW6TMJLbahE4JolIXPLyIBtdps
7vwYCU8srrJPlwmBi8CzLFZ2Nui69jgpjoEcFXV/uEESb3cOMENTeWBmvQk4HKft
u9+hcV6rjgC7vYeYiGGD9O94gcYKYFaobu5SjUQrP6EESedQyZHxS3kVwXCNHefq
ig+mla3GlwW4AxpjHCuJrD/vZ34K8eA5JSrkfagRccppzPhsrQuYIaD4BxIK7wus
j0sSF5zubNnz8MgjU7gStGOdJWMJgc+Y07Ev5HhRLjx5Hm0OEhw1geNdBZUbXiVr
kd5rdGUZ4kPyEdiXZ3L+PD0arIy9euPGsMAjBiO4gcCbpa31+Z4gr5uGe1PifLDJ
rOkZP2qVkvKJzI7WU3YpjzQrxCkNYJp3vME9ZX8U5P0C1BojrF4sZ6yyxlx2Us6x
1jvvM/e1F5J/uc8xzu1A2myuM5eQTbr7xogoafOYX+Q2EaE+GnNEWZK8ecvVDM3I
0ddIh05/TDWQLgIXZ0E2vcSAOySO6zwLvXDa8b4o4Ocnp7gOaPN8H0mrHwlsmqzc
no0YHTEorgkiQgrYEK3fWSWH0Pau94lH050f4C9MIqlocqKYSN9KbLpknPqx0v6Q
zJN9l31FVgi3ekt8TIqakz5Kbu9+L+hxmU/AG5f2YOz6zT22wMG00kHuO3rNHeM9
BmJNBIb+MhJncUIxBZ2hE7t+jEA0ft3bhByp94aBw7CBi8O9T4m29Zrs5EUO1Gh/
/kHawjqdzzsT3EMbsE3h52d+gIXJ3PbE1FfpnVDiGtWFvbEinOIGRKTZFAbFZsXE
kPS66GfP7gvP+kXJ8F4AAwzcnhgqDlkFrKJTa4ucennt6ESmzPaW+W2v8PsP0Bfa
aspb/lamNZUbqtNQ4QgPPFbBChnNagpH8xsbEJ7lCLglg96yjHwnFzEjtWBJmLnW
x+B17iA/e1nyVlMzFpQtCf+VsoD3UZ/CUrt6szeCWPcGxX+N0S9UjhNFt9rQHL42
FTOIR8N6rYcAc/oYDAHpA7+T4QQxsspRowLnLXkpnLxIqfGLC0/8L5lKOQsHNXLx
EsTRsK6pILcRbhgGCA5Y++SQBHoCmRwjCE3IPk9BywRjClICL6pUt7sPx1SXx53i
Mf03RCyR8r3CJQGzleWl4uTNRN4F1eYhHjaZV2wvu1WdPJiHiMTLsbf8XdVJw7Jt
xL8a552pydH0AfE1X8+Sl7EP6UIrlt00C3sbHya5TxKZk7ZvcW3rdQrLVklfMrVX
ntUPSMA2f+5JuDXAx6ir7CHctp2cVdLUWV0+PYGiO3PnJGSjdxkMHAHdutrtNSO6
F83OK3Zxv1pBn3BAj6alU7Lk8ZezR4oPTvT+NVMuN0nsHhnv9ILRauqH82yMIZfO
eRj4UNgf/61hcqWI6+KYvoFUL154MC3c+GUlO/p6T99WtMf3dckY+GNBfM9VMT0h
GGht1mr2EbuqMOpi8lUS7HlW2532NZSNIWEtaenPaqSILFhQ9BQwoj6jeuvk5Scj
nR+/ya2Hnng/nU6Kik++vW0KPVjndsRaWp3h4poJHEB3nc/rCbbf2L9KmLXjc87c
JzGHiu8w05ertSXOHWuP90pzouBE+N6xZq3XXw2EOI35P9mddFYUi0w0/DCMj7QV
7brOrxP3Gty79hsymjQ4hew8gWiWSVxyF+jxk4EwJzUC3wlYSVE3gFi2XdcjGahf
kLpteq68YaUJmeQne6W5XUJwoIJEkMKOd9K7ZMXjBr5q/p0KAsQI9/uYmqlepCb3
qvt7SFkFMAVC3IKjQjMdKlMDnJkfbqc7qRdqXD0dKX3qLlI5+A6wQUcIOKvawOm+
6kBtexFGjRgPFR4BSIBPAZDdgHgiGp12XUZx/2+D56/qYdLNM52nVhb1JNm1DDEB
N9DN6KiXKa7Cfb+ek+Piyp332zOCrnP27maJkXcR4XcdtJ7bETcKPMez7uoOyYe7
sUjup3pSm9dkTMUDdA23A5Z07l1YYQ03zyPBucZlscyGNRmwqQOIMlyOUl+TAo5P
LSlLgRmVJRG11n/BVMmGQBe/CUJhHzDJ5OiFi/rg9gAeuR/BfBOF0EOw8kxIsWof
hcdUnflqC39TMTqJN2Yu7yeNctGBneiuPwY5cOj2gdmpx+Uvvcm+kz2fTfbwnZs5
KRiYYH8Hck1WGNuhUKSR6oigvgsTRg6j0b76rk1lVjHmNOgda56u3YqHp0MwV3U9
XhKkh+Wk3WahJEEgT0aQgJc9CQkG+l7amMCK54jK2D72shW4KCp94QAm2RpR+uFp
jK38wV1NbFura7whOVriwqfO7cJnqv/WZFRaXxWjU2/oF8J4hWokuTp5ECJ6mONq
l2c44pKiNUuftPzvI9Vnyn1V30Qgje6kqLAiSkjBM23h2Y2ToISa5UYjDk593/tI
TE4VjXffwdH4iuRiEazlj0swdX2XDgwWPsPYR9Yuug8TB+Gp502XRBb+S3CaJVjr
izFo6Hs0Kv3svGa2zXW9BNeJXI8ZEWluO/QCPDkUHAuHZ3WV5eVbRii+T/rXymbR
ObptZzMDzlBLNmhwjURgdg3rvGyYNXNwzfD0sTfJKC8F1ouC9U+VMLGtAPQ9f2a6
IoBfzBTL0M/aappxHgKl2DljG/McgtUKC1ltgv5O9xseLW84PuIUHPDJE1cRGY5Z
2pFhPtZYJTa87M4gEEpehoG1Oq0Wc+4mt3qPyHwIXFuqaMe9K28O1Uf+nUAIPdGa
vOB/8vnu/yjuK/+fEwPZ5QERPYAy8ECO94ZFm0FVGTPuvIQ5tID/Nh7QL0EtLdee
uaz8Nv3UJ2xy+n+KBJ47ozd3lkGRn+oG09QuXX15Ex4tfHU0rOXZnUfmbCmIc4GQ
yBItC6/yx4xipKSO6SaA8wRb9RmYLw4O43Yxt5N42DqrxCZCEdv61guZxjddp6bl
jC0kq4APM16VljuuozvfRUMKW41DuqyYBnUoCdqBYtA64rTSabsIGa5ypwg0RQxn
i+7/6GV5t5G4VA9Fs1TPtzQG7TkKT4knbMMIUDf82nlk7mZygzV1I2t13DgT5eEg
pYP6Nvb4gfmFNG6UbgTZ4Bat3fuKck1jAn/cVesQn6AvcqT/U5MD8k1+pXrZGwxy
JOHzrzfEFfAjIxNek+ICYVMbPaJbC2lfspRo9+dm9Clzg2j9KX7T9ZZOhCefzAAr
RDgmcChihgQM8q7BvsCyJGYBGGX1qk96JX1Ebh+VjzHq+BziAVnhZrMYJfUDFp7z
gXNCAmo8O8GTO4F4MAdzq4851xqF68/+wJmoGt5V/G2/JKgYumlrmx5id04iiiGR
M1wfL6DXLBG1rPnT1zAx+ZIaavHUTmWRYm+/O26zqRo8qxS39Dg661jUNpAzXzk3
37i4w8PTyB66GpoQjdDvvqUAirILeU8u6Vqa9R10v/u4Cfl5Sp2b6MsVQb7SwnlS
eWKFCHc6IqVxzgT/kELupzKhE9eFplkE44YshDkCdUE5DD8JuBC04cGJ+SU2lzIk
BQoHC4FIeMMJ3hSlkD/RRr+UbPAgCpqWdjPUY8CEnEAgvYxg2lo4NyMsa5A92kJl
zfdRMXoMtuZREwAphZFiwm30tTi0VFz5OqC3EHt5ejWhty9eoBEuX2BCMZGMZVma
+2BANe4y944b/sCg0JdX4OGjQi6Klb7I1xrDMzaZ5c8k7GLsTJmWuOJRzgCyP1LG
bLNaX/Oh7ueaUpzrHmvqIpLdX8HlYXW6Z4XcmG3I6CFa2PDx/MleKtVd4t5tbTNY
XG6WwPGOWJmRRnR1Iay/ZBxm7cL8/HF692ABpAF3UEeVQ72NKzESnS0bMhd3Oc2f
a10eayUqJfPKr3s5Sj+nH9s4orQNG3a1a1srLBFpzWr/y7t/ZG8G4Idv5oYq5tqd
Jch5ob4B7xvfZj5APIXJMnxSP6wmMvj06XSAnvPd0/Ycu/+fHyyvjjXJALU0YXdY
cUtx6ZkjtQX5Fv7VXpVdJknmMxVtnW8CfQOOvToY0WqRsX2jCDB7jXjd0TF/0i2u
kupqmoCo/dOgSkyO5RO4jr3A06vyovLnVs8EAIdtpUh6ARKq+5HJbzro9dqmIDNa
JS4tQ5OZfPlS3xxMUWS9/BSNMt+BtCZKTojU2ZSRg1DnGWz0SaTHkLo0TP8+mX4+
USSVGXvnEJJDVFhYUdWOPMXrNF9LLjCLVo+KyJEkpzoQYlw+2+rhI8o6G8/Gtm6B
J2CD4NS3yeHNnRCK1bfyfcPopZG3Sr1+SuHjvf1wzYXZfRuxZjOvAFCupzFJ648o
3cHSU9Iy8SPezdK5fZKpxpPU9Mb+4MgK9AJ+11v9O2SvL0e4AxaUTsRE42lDDi9B
NvOtRAWwswAuuu0+ddUBOcaLOZ21D+f6O/5Z7/lYtQQxtNnNQB+1jc0xXrKLJSz3
RVCZhz0zvmX9ODBBx8oJqCvS8lyfN7NGgoWQKSba8tzMkVS29WLxuMU0mxijbfPy
ErZIASirl8LcTFkIt91Q8fS4+rwvC94rD6YeR6KmmtcCczQoQw398gO38Pf9qtbR
wjPinPPIRu7FgFKSEXpV2PEbbQWekHvK87oEHBF95zP55I1qV/8yKK6dlfccGv1W
andWQxyrzYXdzoY23z1Tpkfhc+XoI28JR3H7ZMupW+0PnysN7F0JAuUNUychnK3H
y+nCZ4vydJQDgtRqdk7EpAAeSMFeSQpkXV1t513NFZK7i2BU93l+Dlen7efixYyr
YWCi/Zkk3wpY+xYC5F4l9UO6fH9EOCYH6hktqHzj8fr48LAKpKINgEYu5KcWw+O4
uHf6W9w7fISJTAoA+MVf9RA9AArVa1UswEG1RBSZ47cnJejAJMVzK3/nKDS9r4B3
6dn1DCObcNjkLsgOUgK92AMvp/CXaTTTacdcHWWBYFCHo0iCUg7lgYRo/uuz4XXc
N7w+OV3bglyz4Uq/p5SJ9SQoyCBUJBzhMcz/bpKfq+uExuKnu0+a9E8jBRni+egH
eIZpUzqcZ9Fjq3ep4tr+zp3Z0MWGSRTfkW9k/8gyDXkKrfKe3Evcy8qGYGhH2I55
7B1vsVswmkjrEZ/cSZW+lmpPJy5MQ8VBQENuvIWvtz7sZiEL+c+fTh1GwhpHCbi4
pNUsjeB9vQQgwl2DN6NpkdMDce4kBEyLf288kc8VNX6ZtCczPglejBruhjQoHT6/
Emp3iRXCu+btfEbkJtwIC5PJ4GtfvNs+z1Yn8glIjiPTfBVrtd31omSsBeL+cPZJ
8hZD3uunwt1TutQXC+Brvw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JGwyI82lqjhS73DXAo4f78n9im0jGGDjuyhD3dZmvWIv6mLi2buuH4CLXnj1ugkD
xVsyUfci6Xo2+XwDqicmRkmK5fOSRaKJcuSAJv/zq6OUgMZgvHUS1T/TRxMCWDc8
3Y9b7X+vH7mxX/oVYNvpzx6Br75nL4da36rziXMLZIU0T8BEkY+OQLO0fthXRfqU
pSG5RiQC9gnPErIdXzpP+EujW/e38n3b9zfE/+GNKXVKZBM9oa+DzlY516Z2EAmu
FLpBb6S4YfkdcNEW0uR9p3wjcfOFjL990vpHoJr6nNt2Q7tbvxLf4g/8JkUMexnZ
QS2RrcQ4b5bfTVJO5feuDg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4928 )
`pragma protect data_block
a3EjYEYjNp48FyqEONXFPorZKi66ytn6AAoJVdfgmhFTEkCFfeTbTe8wsQq6O1Dn
tze7xyMvObRdVgKu+eQJwODYdB9Ik2UG8FCysnJSwnWTZk+vWKRD2ZJhDliVVU3b
f95BanLPNInMhwPgsToFwBbCw1c41za2GaULS6xjrkTru1gzGppp1+KQLE8qoatG
N3GgXjIvElVQZ+GbHDj1qdwkFOLi8xM9bzlEY3MuN/MrTifeRaWfmlixEIP3Qq7H
1YYtI5eaKGp1BsARKTW4naRG/ows4g7QY02ZetQ+8qqFyqqK3tiPNdunm2CBoQrh
TlGQGl1H4wct98YzQKjMBYyr8iGhiNY7qCwx2oSKNAQ+jwBrJLK+jxOymG8BA9At
n6wAeNlifgqLwg7P4o+TuP/JzmVQnpTIv/cnbRmrCatMmm70ZR3h+wvu2rBX51HR
0abxYiB7nBaKUrkBC8RqtYslo7Lml2qhpL2mftXWoXH9V5/6XSV6smKJNhEZ8NB2
RxP+582AOokJOowE4NcPbnxn8TBrGTC7GYZdyHWIqIgxc2StxQ/8p9JRMoAUhQ06
YPksy0setGfwRyCngh6pTy00UEtA7HMlUp3uYGlZ5q7TekQS73gr7BltWEj84sbh
DL55RlOfL6t+LrzEJbemjvxy9v8wciARhr7jqEi09BUt5nirgxKCRdCz6ZfDtR5R
uSWM4SJFtE2wYtdHeL008HCSabPqqdRMPS2zw6BsA6d8mppbvvi7cXeQ8+MWfnsn
lAevUdfgo55c7q++CJZiCB+cMaOTVd9z7QB/FTWxB1yNrriITF7T38o7D1PGoim0
JCE/VCLh2KwJhJuDgiESHpbOcDMUmYz9iBfxKLZ05PX+JmhYNyNHWGlxoCkhiPZ3
JBflIWTd8dH3OplMq4N57/jqIzkICLQlwZSofKG41uSzxPKawnwxFZKxW1UavLV7
KGcf1YpDLxzpR5pvSIJlbVk40eHhmweA7FuUM3zv4jI02xXZUXYHGqgIMsXERIqO
HgeorziUgKgn2PL+e0RVgPWwCwooWxyrh7g4FWKASgE9lM2yNJch1sBBoqbHvAg+
9PnsMsTQuEINILE8hz0seQ0l8gbu4txssOLLg9IGanWBL4VdsBiCjj38AqGWkFDb
brFrpUWIm2dIFY1gldBUnti2YhsHb/AeHzrqdxuaH+lu4+I5suLmyDysLSmOC3jD
DC7oVI0KlpIFfzttm5J3cxQlZeCLlX28dmdq9CYoW98ZbRHXZwjIX9ZNoYWGauPj
pKRgWzgGLZVWqZJvaVIfRlJaRygbRfQV95UpSeKsTscrLAsfuucvMW9JmdwaM5X+
Xu1aKDYRymAGDZjYbOfuW/oZIWn63IQdehKYYhdPcPK4xbHFD+J00xGsUpim+dcC
GMuFC69VJqWY5cBMPt4XhlJcXPMvjdvMt+B/bmW7HpmpbRMWYkQYi+kG7axjIfK1
17X46jCeqvGP+igS0yFeXMWdv7Nr3x9bamDPobSDFLu0RZ6pDmqvXLdXgJz5lKO0
N5kIgCUQFr1AWwC1ULRAfRV5J1B20DKqOlQ1UopKdJldCM7GHabtaY8blQFmp+8P
PoO8He6Fxg8z0fE+IZ9G1Uf22oJpqXfuhhoS9uEJtfDuTjIhPmKzkLTJ2y1KcTv0
cXIGS5iEZzzY8MUFd8+EMRb6N7UV7UiHlba47TGJBttf8Z1Uxn8f0sq32bTG1guU
Cjqwds9N0U0YsPONDXGpPoELc/13Yu8l43PrEidKuCfYOHTcLiL765v7KVdDZNFh
fOCdQvItv06md01N8vUUFd9MTOQSdkY/yqHEt12XPuRs+jKNgfo+/HYuQuHd4CpX
FnpBtjjRjx/Edcc/+f53UZQjiK0lRzjqpkKCX4r5P3PEXR0BeUjUQkdTzUNtNxb/
Fist4wCocHfdoMi2dnaYNW8rB1tGHTVGSHuPh9viSGcLkjCDNHqXh4nFyp8C/QgM
68QqFUKrNAd4AXQ3fOutLEDGGmAPJQHuAyYlKabtLy70j32l23KyR/oJ1fIuca1V
zZp/3zHXGTeSLig8QrDFo5YxGzGeGqObYJl2lu+qJ42560cCO+aVDncUvyCXLJ14
JVRObSIKTCdYMzTYzsHGX8aor6RiYzcbypgWMYN1I1JKDEBp2TofBHsoZP1H1FZL
F7C38dLHpwDi32hSZHGxJiAKs5TGOq0CVYYhLA6iPrgplUF+VaDosazFHFeljL6z
DKVPIeWP++55Xvpp2XomqX4QdPccMl4EEy/DuiQ1fOrMoZUN61h9jRL6EIM/swd7
LoK7ZhtGxdNFF3JhaZkeqB6cU4/ubGBXY2Srdn32AlAF4N1lerthJVXuXJ5S/4MM
Hav7D4XpA8KJFG/+mkBmV1yyTnFQck4COwZg2B9czr/0n1WAiVKC15bZCg34GHmG
nhODbar4AXvMf7QbM2C9UheFcqIbK9AcNzi7UvLCeAHqXqqSz7DmQBy1IAppRD+i
nLsvUCCIPC0rdpWeaUipKIKZzTdIPrFN0kKct9PKk9LjombEvMWj4jKrRV7jvqAX
iiCIiAq0u4i69mWB9exUbFi1prPzmHn1o2KRGcsGFB6xVUaMCkZn8I5Oo+YNNy0P
xGuQaL0fpkePcognVb/BDhNeli3jutWwWTU5KHniieYnwfsUHcBQLC6guz+AdBn9
K23+SQ6x7y/O5JbrPGXVKiSbjz1saBcISbEpCsIvdw3o3UPBg62vOnxnMpjir3+7
lQ3wos4jJAaQ+pqomBZKfzgiYHNNT3W0CFuqgotKe66PUxxm+p0eFUrAOiO6VvLo
yqYNcQpwTQ5gtSE2ObnRLBjAxEFg1HGRIh5FlTMT/Yw2wWpZABswCyg3jo6oTut3
39Vr2frleV4A42y4rbYpW8LIqYmVxtqLoBdW2Rp20wx5fe1bUmMMwkcSE8pO6X8K
WDyissj0iWy719G7/Z3twlxFn86HFIuO/JBXinm22+ytSf4zNVPDeOYP5tmu0HcA
NhriGJl+ToMG7Tzj3VJ+YrStv0llhXC6wJi9QNrND/ROxyvq7DCBK2J7GKyxXoi7
dV1bf4hpN+AJB7AdP+adQfBFo7/9VS5JFkYYtN2xrUW7k7XGFkhj0vvhGVTzY9+G
mv20z7R2E8W57jOSqvELk9RKCTffosw+krCZ6J2zgRFOUDGkCZWXuK+XM0V2Kjrj
1mMF800+KV3RzzJrAJD05HQJBScDxslyNQlN7av3vBofdY/qsfD/zJZFzfITM+C8
YRabeKTJU5syEETacOoMfIy2TNGlG15jqzbn7XPA0/E6rdjl5icTtpGMwDR/L/T0
kEq+y4T+oIq+S7XVS4olCkwjeKmdj2opsI4GR5lmwaL2iG/yMsE5KL7IL0S1VrcV
ARpJTahG3Cg8WmrEGl7n3VYDBkLWic7Y+BYOJi0YNSH/6ZnVRzmz5al/A1g1jk3h
1PM9Cj6Mb4MRqgCDVCGEU5yOmd7svnxWtqqGt4ueTpvgSN5yZ/wK416f7sXoEGF1
/WBxrc5CkUhkidTRzLVCr3IIMO6X2btJbra+t1WexT+yVjGC8Q8SK3SEs4q/fdQx
9Ce/NHMamxRLHmmU6+O4v7tz7I5ZuKjHDEqsosHq/DujkntEKVjXA1J8OB5FGIQV
ZRDPyBCrmj5bt0i177lL4HD6tqcC7jzbCtGXv1q2LnzjKZ5Y4pDdjQ5uRPh604ME
W4lS3uv4Sl2kGCpy6/lHEB7rWY5g0DVnMUqqWqt5R+4AOoHe21ppoWllzHrTRcn7
G0ZxmoILl4x8SjWsQRyKAKrNJWoRBMV5UIPMV61q4I7WA//sWZDZlNSSy3nSanhj
sO5f0urPMsgJlZ5rfV/I09KkguULx0TbQmFL4Ut6UzbiNUJyJ/G0K1bimL4Hz8CM
TMsni/OiOZgtRz/TiB620rhcgLnc4b0m2AQJ4AGJ34MC5CMuE2zWMzu2v0VuJNl4
gUiflkqsQDMrAMeBxXK/fLDgjDe/m/4/032pehACPGcPKHjMSPtoswF5BEHPQnQp
ROpx09a697LjUvYLwbnxKV0LHvzQzXTJiqoNTTPdkKxQv8UiLoZQK1XF356FML+H
8BnbfPBPqQlAxULS4MyhLg7orXwMAROeRX1DPBJYjRvClIGHDkFlisdavZ9178IQ
mJPvJBU9CqM87f+JI3bQvlHWL6zRiarhaznmBp6PZj9l544UJ64DptUwhIyRyUp3
ZGXbK2RlpMEvmgunZOrKF2J8bA8gu4FedWYZBFNRzmS6T383GFqiiK7qBYWfvIHQ
A5ioR+O4tH/PBSduYUz0tbY7ViQhSCd2dUtD/JynB3csjgOhUGFS1teIxBShMYC+
fNQcHROEN2CiF5ub0hSJ9IhzZsV7WKQJIj3F31VjOkdHuZeaIZwrR4VrFlyCgGc6
qvuCiQlTRX1L1euMxg5sva0Bsl5lcRDNEROxymo3farlicCzeDndE2ED5sYkatBD
bWcon6DRVU3sXy7c/LhrznyHogZYqcnq+prIBJmjQ8RD+XLpaOuqns6WBbQ4felE
cNvKNpH4L8SB836cWtFeRBWZm4jF7RYTVv0Q/k7UpGvV+8gcrUlfVFx7/+uJOil0
8WYBV4XzA1mTbiG2feeG7ypidPunyI9I4B+zFjpPbiCaeyWpLXpobWHk2lVbqw6H
vt1+Uv7HNxTo6z1fMgnvL7BEkHSB68+De3Rr7VDdTErMcypRYXFDW9JyWhzSuUyp
144oEATsRVMFKS6/ZWCS36MJZWipQFUJHkacayl7WP6IVO4HbduGWjmq+8mU4g0v
jLyGbG8cacqX0GHyRylwEUBflGZ7FXhrqpvpGxT/8klevoVjWOjq1ao2q7RXuprO
FbDhq4j5knTBBO4eEDCE5WxLDOGXetPXz1otr2MPTulkbsiZ3hRutrihlkoqgk2G
UekWadpwBLbtvowc9iVEpdGtHhliiQb0kAnNNrj8TQeYuNO698bcBD1LdLRjZNu3
S3LU7oUiDM360OBSlUQMoLZEJiE1U7QRK39Z95q8swtA8UwMT5SLK8KjT3y79BOC
b4Gp/zhSeTtqOIq9T88mU2jhFcsJUI8AoiUH1CuAmDGMjesxwMdnkOwLghp4Z2rL
BtOH/rvC1trLUFyPdBk6UQzxfQW/jUQ1KPFHnUoD5G+kVDqOcu0Mk5U3PCgyjaHd
bbwL+xj+JVHOTAmYYRy0+EkSAUo2MX5nPdC+Nyj/b1S5WSUh9amXzKcOx6xLaJz6
LzTgDXSnt18Ao8zFhnmZpYJ98zNfC55rXNUMYbNxAz5HIWynr5mloZjYp4nJ6sGE
Iwn2yVnWXONZfiyo1rnaAoHH5SzZk4Gb0XcmC8xxq35N8euDpMI1yY4oRnaQ42jL
pn5up62+WXnVPD/V2hPtRD5dXKicmY0TPLNrWAuJtfWP9V+9WWcR3Crd/0x2U+Ub
9E1nw3JFjXHESLJiGJkoIx1B+3w8OzxNp+SyJf58kfSPT/ue08sxOkj1Ejz/uTBn
DkCcqZf1WtRcqrSwAuaY6Uw1qwMO5mShWNiAnpcmFkbl2REbRXVG3NkTKy6obiOF
I+iGhhzte9F6FU9R/RPIqJUej6N87GDpWhe7eTSPm9OhUmaQq/YoV6OY/u0g5+6T
UHD2vEEAAypq8yA1/ix3YcPsRF+yOppC+qOfmBtKlMXgVgH0+4SXObsdX/uMaC8E
6a+8WCHa2jMPS78+Tsq8L9jFgFkKHizqRlqulVtCcLy8EL/mb035L2sj/dJrfais
p8WczZSbKSZPlFwHmNAzFxbDN18U2N2NPFffk2+Ufj0c8VpWpVQ8lZ1GRltSoArh
JtbZCN7f4vROVzr3MAgKkIdX4Eoln8GyHuabtMGZ2aH19EnGqt/7aN4TMlD2iI3L
0EsrKX5erl/aWD4Rw8jb2NseAWq6oaLKoNzChputZMaLzuGTAf7/tWN3g7FNyfJl
VAZarL+5uJG+ZMe7tLPyZ96YNw9yXnkcZ6FmYuOc/9fbZbhnstA+xJbuom9NNUeT
z8e44fmdgPmna4/UD6aziTe1Jya9XeSmt1t0c9PfDjfrd7PjL4p/lDKMMPLG3eyu
h3r+yarQDKRYn8RUNO3dc53coLAj7wMyowPPbEiKMQJjlaJ7kn5XI+To+cH5cYe6
7pzNsAHx5ZFDC4hBzzMJnO9oRQpMqP2IK1kVJ7Q61qQ7qLjKfrQ2jguXtS+Eyp8H
EM7q7Wx+T5z9r5Hn7w1pPIji5QLND4RFdnIGF4+/cONyAeiWkFGqU+Xl7kOwgIjy
41bT1e27eyXNFQLnNe+lLBDLStDfj+FcjSr5dDeo4+p7ATNGr3LWrlzxj75X3Pll
ex3OaVabpERkDguNKHRjQRt8fnu1MAkT72BzpUF8x6ucqgEddJZ9kkUJ/SKTR3Vd
ZNIoQMud+Obzs7oVwVhjN9TZV7vRQjE9oKhgRNDxbJPbc/EGwm/70zcsXRKUnWns
pVJ1Zl5BOvBFuVF2iV0UuFwAND+JdD3j2N56iqSeflLHcMdZG1Aa+FuWRkIuuSji
8dhfbdm326potxxXp0HKQCNUmVgB8MU126GMNz+70Ag=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bxFskYBbOQXcv3pWFeFRRIeNh1HVRNwc+dHKPSeiCKzoo3kVvg+M8rTKMyiolQ5T
KfRafV18fmgVhEhyXq3HseY9nIYvTeEdNERvWEIQHeu4VApjXcX0IojbcA9eFoTY
L2QLi6b8q8/P/neuqY7ds/YFjBZiJRfoFFcmpszjF+JKn0/GHQ2Aw7aL+g2bJD5+
TCq2m9VbQpF0uxrmW3MSfGi6OeGj45K8qeK0G6PAFWBQQtQS5MBqLKh5SXxWJM0i
5VHJU3WXeSvSENZKww/nO++9SxReWYmQvaULpSHcn6SkEdfrm/VlZfuwe1B9a4JR
FyHm8qohtnKA++AafeDlZQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9792 )
`pragma protect data_block
LJQDPCzqIZAmBk8Wh9COcV4ugAC5kl7r9ajGXO78aX+JzgC+AcbNQp25g2hxs1BY
38eNXTX8NgsvdCkZL5grdVVvq6xgGgi4nvnncMQj1LNRe5WiChyFZ/s4aqOlqWN5
l8d3DTaNI5JDg+wDnvQl6J+tp330HVqxXctrjMxuVE1YPuZwzJCNz4H5Oh3IBMd5
qHv4F+PziXKd/FRnVFSRpEYbVjxS4C2xlYveoMpnN1NoUPKaEEuwXIKaRojcglpT
fhod7U3K4DwnHmIo8mU0J/Y95pt6Suuu+z+6BW5wkcnXlktUa8tW9KQZ+i+FK/w6
x8HWwfZiDrDPS4rIM0NG1TRg0b3oinDf9IbX6yu7YD1ADPPEr1KZy2jqHRD82FWz
12jeNXSZ1X08fGuE9AGOg0k6gL1+fzYvdg8Uw4qaw3O1Qzp8vtIOwbySq6z4ZKS9
SCUwebMLQs9oWZwMUh1Qhu60hP5sU+s+HTOY3d1y/TUspDA/67nLDbTpbFWAf3hp
ZSh4XGzd2td2TzpJm9u36eJYoqzhFtkQwM62CuNPWLCvSdxMOxaMcBna9H/0JEaR
G530zq9OaauFsuhX8xGZ0zYNVETg6ILteIkGwICHyXEYuq5j4qnc3gyKcLQyOK/D
mFiJx6JYp6lkCtOTWRhnP+YD3gxIsilgEF65yN1hxOrI4wKBCZh8voD77GWlspTZ
l60Uc2OrUwCjczWMoMJD7vXmadv2V8cUCd7zyuz/V5VBM1MXzltp4kix9i2IBsFU
CuYopcmRVA7axHEOwwrdk8WkW19w0+RRA60Sn8mIOSrvw9W7pKypkhU2wbgy5gWF
RsuJvIfEqvSNBlKAxmvTNpa+cfq9jt/kbXR2eX2jRrOsUo9zFNkRXr/TP+aqFfvH
WVaNa6P3zRmZQDs1YGD/XlWyUJmxaQVQx9Z3ySQikRJyuLoAzZM5Hs4PfWPPMuBd
W+hdTSn+tumNBwxXD00ZrM/5ghIapJKlNKVA1YtSLwfH6w5+SAL5/aqylz6+YiCh
f+ctqS5EIKFQF1ZEZ1gJbZonHjqe1jznnpaJxx5T+SDu2XvjEHJJevVqVte0oz39
QnjpKb+tenSxosA85oEvJJr+VFWhHnANu17XOhaztwmefjSgIkXHdNjognf0cd77
eoG/rJkAXBn1wkfzTUz/6YDr+RN9+HTH11G/9nOM013MPPeo8t5T+ckjTcJLvqmD
/RXDokD7YHdFq51zfD0nAenNtBHaDyc4za0lOD5H9JUeWCe6fskJZ6nWYywgfrwd
P4E2E6IhWvNcl9ADeJGp3O2wkjcpMs2bkN9qEZvKu0dlgRsIsERXvTq+XZmgrsFv
w1EAfRfiSNqIvdTa01YRg9lMCCwU157Zisp4wHsglgjSM5rLRzONVdaUgFISG8+t
PiZdAMWyN4lhiOMdSWsLwy6TQrB0m/GGgrePtOvU2aeCb3IpfVVNzg0WQi0CpBfL
DNPetwYF64sA7MMOqPQsggrzsJkuD/khynnctLWAtZVOoc9cso97vcnXB1+6a9hB
rhdaGSj2T/Bs4rdDRaDXY3ay7LVmlVB6v5oAozxRwQRXQc96AO4W1pG/azQdR3OI
Ddx+xZH4VMP6pb532ekyYCU6Wu8BUbTQEkIAdCjOyhlkRiCh/MxuYYNx+r0QcK/s
zLKwWc929Z89c8eUIlNqMlPAmx2qHHjckAA5LvVr0QLe2TM1WdDkPPjSqjx4iSBq
latocVWLKhXvFTHChHJaNpkTFlY8Jd8gToJ2NVcRgbEMER12rwaMe2lg7iQbdNpr
icfLJK2KKq7Ixc2t/OEvZ+M/rAlZShJNM0CHxI28s2miBB5tnQH1I6NPbLHlvPpq
PYKN+szer1NPYXeSm4IpEIi3/6ekdVaqOWqtuTo2gtdiDXd5tZz8mE4ov1PkYrV8
aJ1uF3LfKD+ygW9mxln7TZCl1R8BUvvWz1hERDE9clYLfTU+EI6cQTH7dN0weqdn
Guppvflg5qsFxHAt/qGsZHHIBqTeh4/UxlUbaWiBrz9YiGdi2OAuDJlzdxiBpqJA
Nnv7g5qfHepyzONHCJ5MJH11ToV2qXYKM4ayEqS6fTA/JBB/DmC25a4hP6j/gJ6v
DLHO8w5azfUZ3ovt7+PP+5fdD5+OyPNCBmDMjfSnA3cnGUfLr871mgZpSpj8f0ZP
vJ+eNmFlP7//oOH5YFqeyIZqp56fywmKNKZmsqYAOTlWq6sYWHtKfmJRdMW1E63L
7mA19dE7cKxZTUP1xWYqXTir6QCuKKEvZ27XCOT2/K9xP3n3dhmXTRLykxjDPku0
h1lWHOyDkFfOulipCgVVLjuuBIVD2nZ1x5LHjHjkPLc5l4i+bxpdbqGP/JCICenz
p0DaiLayfYHnM8yARKs6+j0dNM9RyuGxG2SVZFxogIW4WwbQLY/rL/qvaKpBdYbq
d9Bx8BK5Y7UomttwJ4qIRAFd7aBLsP1XMVjM8+GM5ejscH3y66wX82PaO/4AoeYu
77DesKQINXvshEhFUHddeOA4cTN6zYEtamUEHz/B2Ynkm8JeaU6+eHTn0wb+a/sA
Bi+LIGm4ecGRqnKWSmME2LCiyU5hpTM3Wr0mNX8zIOj9nRCt1xa+ZkubXwcMqKy5
1WA1V3a5+/QOkulgYWkr/4N7CeiZELKNQC3ODO8m5bL4guz6lFTYWAHOBCCC5OQU
q3Do2iv5XniQptYDZ40JGL9AjY0j3lMjaipWsYtNWmsegmaHJJhytW/hdAN3PejK
fyqYTMZVnmBIlywoH2PGIvUi3S+5kYcdppv1BRZEn9pIi57ZpeN8yaKPoywaGDhX
08gHOg75bbxB1XiAhAoOoVpf1yvg8GkDIMIwva/CCn9qZVy77LKKIkLLWfOHlU8W
ns70kFpAC9vKB6DNYa+NiS4RvD0ytwalZxvDrs7lGDy4R/dcgEC+sQwjNzo+zfLw
cQ0L3sv1E3uLS9KOsjiYi4yMn0Z2Hj/KN5cf2AredIIGqhIXq9zSU6ERP/bl9vqZ
WW/Afh5rk+N7GWE3MRehdZEulZQBG9Ui1KoWyNzBuSunUgqRASeB4B123lKtsmTC
m0RwCHPdfZrYlPyzBn/A+ResGjdQUh/rh6v+u3z4fHNOVhf7cYo62XymXLDXOhq+
CUrYDYaFLETEA8GDUZyqbgWg29bPEI4Jox093O5eLEJmx+eTzLN1XC3erFSGc8G4
XOo0SNjxh8hiJWxp9+otIla70NsDZIouWStuMKVUS4EDlEXcsuK0kHdujrmm5GTU
jVXd7LH4EfKJfOzqFFSuBTGe1egHoHGMuOOIVntPuSyTcb//gMHjosuLRbi+g/bw
wr8OX4che6XadsPp+w+kqMIPHtJI74ZBtBBFMdDFS60FS9uMRbuoPOrzoJdTc/2I
mGO025A2WW0KYH3qzdLOI6OvphIgp4UG7wXydTyRXSxkVM3edIZLgXxQ5HksLeH4
fSp/e23m1m8YfWKmfN+/2YAz8m+7wKpEEbyAjAOnPL0mXtcmt7AUo4IDZpF6tOGT
2XZY++m1tOmxguLZkzbqRKXRdVKNxY6wcUSu5e/jm7Lqg/LvWfcZQRlZ0fUoDDbY
BeTIvJM2Y9nHVR7ZknR6QOjTiEwKASF1FsW/xrDTtQt5lsGZVsDwOuebA4ohtfGZ
gYfm/5sgmzJE+oWWGcBGqmNgngow4+t15fj28CpuoDqJcEabQ7SuTBvOab7kB1NZ
m6akpkL3TBXd1AxN0bYltpSp5u5t6qPOgZDgn+fFjtE+3URXiRNckHRIiT7HM2hV
VVJghPtf46lNKxEE7FgJ06lcWvhjjp/2to7dQ/ckuaeULY7OyI7s3qLtPcywn0/W
LSWGxgThO+LQQBacR2UHIQ9ZBF25p7VZheu/EpZRxNtWB5ny1vzkPEjIbcyq4dw2
gPgv6pBYe2C0Zt7PrDW998bEtp40zbsgWFxaMe7aSbFzxJmMUGJtwko9rOgIvBWd
/nm/UZUoHMQniFVlYASSFHAQaRj5rxKJJvPXrwYwIjv7XZvRUgV+GkdTPpQYPK3Y
xNRQPq5WlKtyxbJdSinPvPoggEjVmFUNRwk0zZOFWMbtpGt/+FVdpLv3yY3bORGz
7GD7HI9Ot4vs9iUu3ltV2G2sU+yLHpl4rIJcq0XY4F4vavXkGiIknKK+1wT6aQyp
B58a8mNFG2XxcExi46RNNJfqanHAEVmeByI+gKWElU51JnWV7+NW11pNOlmZr566
RBAPw7/kJ4C/BEGkYuFeapHzHWMcy4cFTJRLCi+Kcw5anpU+twJSr85GVYoderOE
vv8+NAXNnCEp/LrzZhSdShTuUmw+JGQ413kjYF0uBVI4vV5Ssf+iOEFOsfs3/H6+
HK7e6Mde+itgg8d64MjwZvG2+cB4oHEoCTNVj97EFvY44MhqHlkjSPjsKk1Uycj+
35T/cEeICLC/uQF92OwkjI3a9T1/caX2+Q3X0g9AMKi4K6nB30PRDBPyfc5Z+Y/V
UHHLaQeeREcChNhViGL51QWJT8Zx37Cxo9YW6333LxQmzWbISEX9f8nnL5suCMms
Mj/ov7yLCETAaWH4Mf4r50X3qN7nXWgAAdyGD+aUGjUflsRaheBDsn/18C0j3K0O
cox0QxBP+BkwXGjrMlIVfu7sASGaR8h5+S4bfAyFal6gOnxHhr4wN8K2EfFD3Wy+
vjhyOs6bVL7obfXt1rATy3Q2RCKierNZ/3VQUq2WX8r3pkOfrmvFOskLP4K89PSp
4uoWWVWTIKlfzFxy2F9a0otkCRilGbnW4gwi4voe5FmFhmS6wuNEC0wPhzIw9Bqj
YFu43up7QZDIm/L0R9ntsKhTDKUvfUlprszuJEfjmcW15yJ104EWDFmsQFKG68K+
E1gSVNyxzzpivM36i8Ol1tvao2kEqRDxPrlXZKD3YeBU9tClN5DEAxhCAtO+4TO2
aH62TlFc/w++M95vdT++Jf4moj4RldoQNQ7l6soHHjlgIlDi9TgFSgbInf4LPul/
kQUBmo+YIWgvHFZMzwr8Axt3QxSTVL3UewEt7sUhDpbRdLnS9UKw9IKsgtbhUKJJ
dKx+pWHD0YBecNFROdI15pdrAFLUL6sPjiPdOedBAQLhL3mUgMffPqqQbbgtNbB0
HAqFE44CvPfcMEytGXDa8F3Wj7Sk2OyJQcUz+OV/QvxeaEIrv0CcC35UJTN4hc+W
9UxEI04J896u2fcDIl51QPQ36mAYUYV9wt70WbO23eO85XmJVpRm/J5R3GQC/ihj
a15roM6UPSbXj/IPG56tIvSz2QUe8nzxspa8Wn2tP1pT0wUWbMKIDHP/f7f4ARaD
HKuWsSBuxJurDHEzDzeEF70nUA4DMhMce5V18P7jt3Wz3+slFfqMeUXaSMBy8EhJ
QYuTLOgwh4d1+6/0B9o6He5nTrkVnGlkifjkhCuhy0YX3To76YrjS7s4E+pwUUKS
GiUT1n+RSKIbgeX44KYQ1cQgH39vBX9puZTY627x2CqyuJLj4B9cc+uWR92U2EOW
2bGFz3k0/BOl0KIb/NDMMu+Pm2hvDeBf7By4YzIN93IR75q1aC0vJaRTI8taYWOL
ggh6fhxlD4uOM/FUX5Dkza2I0sfqZgUzLFxZhVd7Q7bWyOXy53TXQoRKWYlOF62t
AgbXjtbBx3RvrwavaeR2pAf0cAyIDfpeYkHcXFpB0qTx2O2p2Hl5XbDrj88bBrKk
tvIbCYMb/IImEOTSF139BQTsQtkiO2uXYGZtwEzCn4bbmDAgpxl/vPcfd2r1i7wA
WAEPRhQfQ5gqvsmlhn+kGUCOXhGLMUcnSBUn0AfhqymEtnXmT+9atoxUUJbaI/2l
9vtKBy6urRBHSehwBbg12PCuaHnfWrRQ2fKXdI7Ls0pY/N/Da+F7nVVrQQKcb1fu
jYhgHlRgJKvt211TDV0tU49IOxkuwhQcxEZN8AQw4EGLvzzpQOenpAPRdzz+H04n
M/aE4RyjTvPM5stmaUTxSXEW7oFhGZYhr5bUFw/OdDjZ9obLltaR5xKCui2Aii1K
IqAqSBiwW/Ang0BM7CeHEzf1yehqnf4y/SiECmusYcb4iyFs4P2S8TnzahRVB4YL
1SeoPja/rXyKwr/N0tZbuv9VffGk9xq2ae687qU4PSTv+uJG6o35NniUM6KCDojs
7gBPBsSpZM/BXEvk/Up1DFTkSkWjje6mvSiSxbqBEXNZ3OgR/cHaAt4Fwi84g+nG
Oq3Xu36ONVL66tLoYdhtTIXapwyw1K/aEz6h9du/mjWTLK5iTDhIcrcJIayasD7O
SWUMXBg2Q3v5ngwhT35HDzHtGVGhyqmkReQef22mXWauPFdzCbaWFh/Vp4g5z4Kq
WagjAUWmG3EoFDdJkUQOKZMQ2jvo/680sNwkZZJrAN6RGoflNdctWd4OeIpTc0bB
3nvv4PCGT3ls2TB3dr7tlIhhytadvK/hlhuwKlaYRalzc2g5N8QPTAB4BqsL3arX
JoaRnt6QPbLh9bZ041cPcym/1/yi2B81/liVrkSvx5isbNkJqiV629z6GXXUZwi/
pTOl4qxPHQLaBTvDNMlWQ3YSGX+P1VxebHRPrdsR+3LcEyH+TTCcC0KA5Tc8t6/i
GVdBYJSmGfsU2lcbn0V/PBzHRsk++FGyKQOZGXO6e9ycsgIFW6jUppbogNXXa3dT
62s7HgjNjfiYG79TrS7WHn0Mo5Dwc3UqmDb64FpC7zwpDA7suedAWpFkOnRh8a+X
JEzTi4bVWWb221GYjRaCP8zZeZOvDrD0Vd0MQxW7yRXeyiTY3nWs41w2rbE758dn
mlxH8wO/UQ5EgSIazNxJUw7Ud+7+78L10TcS6pHn0ZUKTxkJfa9RITkFO952AzFY
0ggePAsFM1sfSm4QVtQqzJSkKqg3YsdxcryPLWpzluaoV0i4EySnp2iFVNSYbXKo
X8BAcWo3STX7BT/JTZP0xtwOMfgCNwgeQeYl+xm4u2VzrYjVQXo2/giMiUu/HB+r
dHNMR/RqdlAbFItl26uS/bPl24fv41JHtyezBEmKVWeuV+d6XEuwMETHGOmvia6i
83i5QV31Hcdfc4+dXBFpRYOsfk7OQKc5xNHJDvyJe0FPTdnGiUioXlZXzhNhOY0Y
S3wcB+ok+zscigB7TI7L+CYHPnp4kI8XW0XEy1nG0uTksybp4IdTBjkIHn5PfpPx
HtDtd1MaAiIcacmB+rsPuKNcPXuTyvi6+/xDYb9NQ8alI/QUqZYRmbnbjiX3oLaV
Gr9QX5vW1/br3h0kp6Hir6K/46DYSwMZVEcBSKx5ydPEOtHVjQPF7+XaPRBwyk2H
mqaNQ6lxlp+nK3QX5/2yxuehJcm9r1gsC4Ym48AkYYC32ZtUmKEOtK2Ugb6HD2jE
FR2mzsyBiqHKyZYZbLv1nvEQOBxdPGMhVIATCCYMgKz43wOccA8Fh2vFJSzs47jk
fMiiUYhSrY1SfKG0QfgVt98XyZP95l0Y8LY6W/Cvnfe0QhkYLVdIgINTa4Xv329Y
bGaOTKP4JkYlpPYnUeY3P9+Okuo+MpJYfcGHCDA2Zym2UA4lOoIeLhlFx3PlctrB
FimZi632oyBgYc63HT+n6xKseZKdRFrJZYYOYzchqo9cttcHuB1dhLMP1JQyx3d8
sOfyne4RRTcBqJ9YNh2cEDz2nhhXnC1c1OaMfiRTZWZKV0m7I+gbVz9oHEU1u+Sn
bdm8Y9UDudjtGWF6lLlHdV1Ue4PiUrr8hq9ZXw0565+CTdrS+kCspLbfevmyrIUI
Dp+tNCz4Gg9oJ6unr7OTO6MJe9S+MvzvGOhhgsO5ZWfWN5/PsOYQqlupF8KVOWR0
0hMB3BR5+l8QErNtyuflm1mpHjgtM0D2N9qbBsLjco4yC4ebjLNQKjtt12CVPvUp
DMOGEFj92Mpad6YcBxfpwZVt0lKcNpRUgeHzUcSBX9ooIFTZITCRofc1WAiihTL+
QcXiPZMG0WbLOsSCrWQ9zAnlBhwEpbMCTKPmZhkDg7r9EjyL8E5N4OZ35UvE9DDs
igTWIBAWCZMOsadGMKD3zN8B2uZ3YPOuZ/Oar7d+foGErCzR7LKNBoSqXcFUy7th
CTh2BOiPYJg1JFdl+Qfl6sqSjZktTotNTXlwIAU8Nv/9o+0k3dj9jQ4+eNZK8wCV
CISrwCWRRJZ8d4qn+A87KcrTWvq6UDHJuBIKx0glUgXKl658s+cXF8pPAu1hak+F
DtWjoyKtrBaWXwNE1T++eNuD+DhaaPDJ6F05OoG/KKuUVG98aGPsEJzvhnalkKQ9
v1o9NmI1VjHHBuKSjGr30bC8M3AogPyiD69+NgRFSGJnTc2lrsehez3CEEuMPVAm
5Q4atFZpDK41E0x+jQxaq/Ns5khuxgivqkEgsBPAHzV4KC0aAW/RvFfR2qxBXzXG
VjNH6nquyOHqujrEo0EBpEXyN/FY/bGOIeqGmcNQSwKARn+ZBw0jQkMQ5l9pMZxP
R3RU5YnoMYYrdo0avfOxZaXwiFgk5qCSE/uyZginmTffDc5ff/wvwKYWdyyJPB6a
8ob2mf9kDbau/2kYF2DkYYtQ2Wu6Le+YjdQwYiFPOhAEIiMlc2g0eEjR9YadKeiz
QpXyKft5zI9G4fTKuVDWwP1AkzGP8G8wDPUzPd8Gqn7ph89vzdYYt0ylpaxeENY3
tJ7aAx2vfDPipZrOSjv60geEkxo+zUG5MEtnrYutW2S/KcbP8beiIM7bvujUZGzC
Aa5S4aiEe1unQrHDfsabxvHwVX4FL2bHyUwOo9g1oYkTm0MaQhQte/FrbUm/AJ6a
Eax6lnw4gGzJKegcNPlG6bHYVrNueYfHJzaV/pFOcN+vQGMGr1Qqg5CRqaery49X
T5EtBvTTL8vSWySg4cHhutU5yej39PNoIdm9izdasqkjPPm9JWhFYZPmyzZKiK63
bog77/XXIyiKlzFAnLfDlfqERgBRA8TO7RypjNbyafVO/HqgM+aR62ZCsBgQaVyy
0FL3HuC97PuEuJ7RzZmYq8aySgyaGIA5OFLLgM51mrpZZsymhNhNIC7M7yvwk4u1
HA8UKm7/bmt+/9EvRowhfdrV+5WwV+F5ottXjzprsCtg7vVV+5AbHmUbucinJcLP
sNcE/EWf/6U/H7i9FGmVuXYQszq1S72JJ80GjC0JTEu+I3kORKbzjujVTnkHpvme
5nmQDx8IhB7PONPmY6ydCRIhsMXDB48dn1UYRAGCs0ymEmV1U+J6gRY4J1UsbqT/
62VRv1nh0t9+6KxsVNO6oIrezrPI2T7YSVbQMHx5sk2G9NrST1IiC4/6NNAs2oSB
1tJTXy7cpFB7kpXSo1ntnDqbnVE2eXMJCuLDeqlGUmMhgCXMjfhKYxt/+npckzjD
GjhIP5A7xTtFPyUJw0E5e+m/xeLE+jQqQkKlySsEs89YrZFRXgS7YvX03ObjYZzc
vjdmZXy/wLU7ipSHp4d1a+dvF+MYr3MsKt7Gbj3FYRyqC4y05UbdD9S0rvF2JkTe
Xbw6PtHRjKMdBXUmdiM2wIvr3BIbQ7nmAp3v1w6TO6sUPtlu1s2nCmJ8zSC/1Lj+
efizOkRD9Q55QFMAb8YwtiSFrEXo8qhTjJ/ppf3VoTIk8DGZiKHJyr0l+0/mRQyU
uHFkhrFDnYZ0oNx6vIxK8s+fldHpWLXEPgAR9t30t/eBNz0ssiSGSeJZ7eRZtxL6
SoqoA/LGkLOBqRMGbdyIIX5Bn3sdkM7LeFboTahOCHpszRV97CYlnk2oiSbf5Ur6
YHqzTakxY4TtS8gvpWrtc4Hs6P0i4zLSxmTlep4o92mJbmBMDsZ3kfkqVCOPebOW
zXbAZfhcZF+kh/2s9nCmbfFxsKqOZYfVUSUKGhGEja6O/7WEzXax1KRnY3awMcyA
a9h8MeZt1A9ARoQju80E/3lu6k7nmlrd/4x0fQZF8sGvFwiN05nnCdcas1dprTRV
E4F2+9ob0xcPOfEJ3clKjgabsFaDCEFSzFconnLM8jIxIYOp/bWPew04nz0pBe88
k4NQoa2OIkPC3QrdxPyTLCj3XyI0FIx0Lns7Vc6bNzRHn09kue933rGrNkO4jHt6
bLnkhcE23oE3W7AC7kUjUYqqQnelAmvT8AlFcxhqHC+LV0QRddJ8C1IQ5lLXZB6d
l8EY0A+K86vTqKDpQQLiNZ2Q6yHnG7y4sTK8kObeSr4q6r1DYtZePC0vi3rdWRpx
heasJ7RL3xQRmta+ctYtYk5CCQKOvS5eiYDE/nnrC5Dftq+tCuXnwNMyWqmxhd4y
sNj3iLrcvK9SKsB6a2/wmWjkosVVLbbbJHaaJrfGaOUL5Ptng7x4ZcJ9MdpwcP7H
99Qu7+WxWG8ckNpREAFECZPulhahzdJKnuiRB+AJjvKDVSGPoQD8nMBear0JLBg/
y8f9ZvVvm1VfcHtcjZDeg6VyytLFzMvP8anXhWH5hcLwB8iZ9+rL8/sBGcJ5a4mb
XcUpnNW3lw8I/vvvVMkVSp1vsTZKMSXyGj7zsRXkX7+UwB/rBHXpQYaBGpdvU4Qm
N4+LNaC651fl5VbetlIKDxlitu6Ra9UAHz4Rhp/3ay1xOb54D2gt3h//ytEKXiGs
0xGyC8T9LgVXIWQ+DN2rmmboPwIA4V4gAAMLZjPQ1cU+ngAbaF2RkkCpJyIHxwh2
rOqQKAfI8YyyreAhb7glF6IJu7ulDaeTG1fngzCavsyghTXEkvyHzx7yYNUW/yKm
C/fjJ5gpic6iJmV0RK9MiYG0ntS9IrN9bARC3CcG5EzddMONtGybdzdm8kU3B4zb
42/FXrNM2+aVsnRAV5g8xp+15ROE8ViiakKPvEAL/a0kne94emhAhO4a+cVtQTU0
Qkr31XlfqUCpfYpYFlJz0qV0nm0Ejk0ckBqA3aTxThc6CZas2/nA8X4I46nw0tQy
mewhhUKbH0UH90sPqz3M+5DtxuYs0VTBf67SDhVU20qJivRYjardMYL5qzwxnYCz
8zhIC2dPNXZZfEWaOiVo9dkgeQYA8LkyEeiEx+VOs8oP5VIbacYhvVFdo3j/VvHo
9Q70WDXyzMAxdMeeDohKCLdR2u2SfK56Zw9iU5qxWDpLzcF+Q1SHwbXwlxk27sX6
4o1IaUEMrf4zlvV0EJHg1p3TNZW1jLXuwkaTM9ASngSt8yCKOognr2gKQi4nx3CJ
1ffcDN79sfeIDJE5E6it6DWsLSFgPXbIKCKOJlYePJl/4iffiUansK0ZzMuufkon
iYr4c1rV3WSGa0XClUCP5SAWQTiR+N483fg5SzNqmfa9ytmzAki6ZS9YCraMTswx
8a9gatBxzIgwersLT2f5uzJMV2d3DQLyWFlJGaBNGU3pUnIywtdHccwDIqIL/gpt
Hd2oTpVoOVch4qLTk2duyv/vIZaE+JrUoqBfBXs/bfpFeaclXxzHtCgQFVeovT5+
wzodGhXF12yur2TYvTbcSq+XSzrbxCSoi1VUFOTMdaVRZu1601u9lx5CCE5335+N
5r1rZzy3WV1NCuR/cL18gEqgcrornHMMbHUN1T62YDeWWQnSh610Sd/ch5LGaVEI
GJCDe4WwugvMGA8OCyev/RXP/HucNv6RMW0fqOX2j/aBglgQgYZxqIPy4JHLEFWR
9oyy9jMzl9oVz9KghWvdMajP3VgHXfx/0fCXWVHbvJhIsvkHKztp8oe2faW6H79J
JCqr3nVZwBKS0HJ73IH9Lsn9FyS6ISJjZ4zzmluaoID0diHU73Wh+P8MK1rrf3JF
UvaNrAfU2c6vb91W12E6RsLEI6L2jjHhoS3jCjXuQsIxNi7THon7oPO2uMokZz83
IVLHfr9c7nLsA2wkF7n070Uwze4Hs+0E3vGgzAt8AQxKtMEg/X/mOlQir1mIPjnE
LQp8S+9Em0pq6BHDYPEwtp0wcETaZ0sV4KeSiv5rwK0AbzuZoyfyM1AXrAe62EBP
6iGNy0Wr2rhSP26V6mEdrwKjvhp9KoAAZVjPW8QgEoi0fRdBWwFMbiYAz5NjCWCJ
D8JhtM3dG6E1RPh6WDakleicgHEjMk4L5NEoEVdZhAb51YNS1lF0alGRMXeKQCxT
1tPnF1BsWDeyXNMjx6wU/EAYqACjJ1AlLNCbonislDRExhOsggoyOG6VemZXQZlT
MMpiX8RslNxRnGk9jCEx85E0RMllSVgkmoo69CaNL+yIPsXdRqErf5xWE8/t5wq4
SWEC9lZHX74PWx9YWEi8KALvbvjtWsZtJGRRE2qp8ikWDysYmnIRLY+N684JWkqM
RXilIouASUGPk0vqffLBHY05ukt2dwMhSLw/kmFSm+kBPY4Luw5/drd1TprSs6y6
RFbA+EToxdj3iT6hyGBkfWJL25KL6OjSyhAz+8fB5EqNRGOrtuSh7oewlE9bgUNa
jx/KNZTMyYCRgRyIHb22mDvwIRJFrkADXMkJikSktt8hiWjNkqpZ/i82rqwLczF3
c1VE9rrjMn4TlpHnqhqXjNNhf5UjAm8M1nAkqmlPOG03kpuJeEu4koP17Uu0fiPZ
gMz4ywSr6rWTDaMNRFC/BJrkawNpNuR97nFMe0QNJ+PHO6EU2/1ceOTZJOBCVdhc
hsmRWd+99GAqiN2+4k85a7qx7CjXkF+IoGRxSqzpExPJ/hlgUVCcT63eYwpy5jQ7
rUim6kqBHW0wJX/NYHdx3livcKN14wcLUgWPMkXz1wC2IhjVxMtd0ycAiXFYcLrg
ribUH7neEh1Tu0hORFtEzHruPcMIPIS0/bii1t8eR7R77N175BtW+YxJZcuunSz+
CB4Fe2ldk28oq3tP2xUDaa4LSVWQ0oGuwt/GP/vSeIRx4/Syicn59sREa7dpbPYh
je4rwwQ9zUmQIQ2xOovKbEsR/L5pPnyo047I7LHd3EU58bzcVEHpzLNrv4QJa97F
WfQ5+znLCs2EHbIRaLoDAELoG4Y/HCXa+jV5pMJNMp6mvUGyoNOD9qsKTgv6hsQ5
37N8ePoUQ/4G57XeSzIidP8ef+0LwOQjmWErsPsK4vqkwEmOaqZ+KhOXyA91y/tn
tAPPFf7o6lSz0GYRsz2fmV5xsDSXCYIAEmzvn6bCe7v131WkAOTi7ZeF+UFc46Wl
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ea5lbaNlv5Tn8BiaXEuMeD6xtUpO17+STLSXwALsd5tIe1hTlJMOiaIVSJeA9i/y
ovWrSpjcMr49a3PoAM8aSARvsGg+/oVN+VBaPyp00Aa8bInp48gWKzO4gAGQe/Bl
jHqW/sY3oimMHZUWNIOCF89MxFkarWiLBYwjMQxWV0GGioy31jQSInH9YLSK3bPx
ydwrzkfP5h/zQ4Z7gcvJbNvxVNqQnIqfcFUrRgofrWZExgVPE2vp/da/A37rfVp5
CQbO+qkbXZYvuSjFQ8uFvuW/UDZhoxc0UXU3Sd3fEI4xg957eHndy/0kHdoUdPTp
DYCky2ES1OcfiNaa3ZBn/w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6256 )
`pragma protect data_block
t0M7Y9PO3iIKAO9pcOQawW2W74A/bEzpAT2wwoNw6MtxbBsIJKeHC9QLSe7GZ9u2
LYgFhy2mH2c6oceAPqZhMrAmPbpX1v0sv+i0fiY48bAg7SbKd9vxj+VYKp+fP1jl
FKojmnawXzUlBdA0Z9zH7Jhh9qS8EqaYH4KTDvm/rI7siEGOqF3qWOQBC9wRzPuV
cwKSM0Q1AtJ/R1F/iG7mmqOYvSyK45b4SGTwZTEJh/3vNQKhST0PlR6Xxgenhvmw
0LzuZCNeN+AzVcHobTzBWcquTXASxn0TWLYSVeJ1vFU/4gSjUVJfguMdlhAJ3QYT
EMHUDaBLL8e3M5+o18Nai8ybvP3SlGzyhUrJfT5OSIshL8Qyjh9ctmf4zo2Zlzbn
d08vbAqTUcTf4ZGO0s6V4vTiUKhwjOPpCsvTr3XI5/YcQHRq5wovYJr0kv4bpcpV
0rwnN5xKd19UaUhxH5xneCH7SY4ZWzXNRk8oa+wMbvwtGklSNq+CgWDjBRUP+2zj
hbRnzpTrSSrH9I9tyNOHZOqVb9pClc19bp4rofpUPZ2Qb0Ne3HYdSpvi4VOEuN3G
K3hyllXrdpXvlGov5i3k+3hQmsQPuW+cVhdHJhn9GedBh9a8nJ5w/r8PTr7jYbui
aterCwdURPv59HZmbbXHr28Xv5O3iVpECa+4Eeo9k0oFK1tWD/9l9yzAKTUnOKvh
B5WuDxu2NnDy3Efxh70ORPDuSvGXe8mLEJDderlAoaTEKMopWSIbFaGbquXVzmrN
474mheW56vWCUuNVrlMc6zXucWS4bRYBLiqN0v4d7YTpHRnzq7maaanyw73RBxQN
buQy9Lsvji6O0Cy2zUcWEH95pPK3gA0gsrMFWnBDN+JR7yn1g4i3unTtjikoxUC5
1aMpNZDKRufWIpbH4siuF+ePKWeZgiN0X0Q8EPKzdKFLtmv5wasjSEsIBts7raVh
L8aj/WH186L9jg3Q4BF4v9DMgezq4lFusfseUfTxaEsUoaQDfi05cVrUWHchhikC
3wUjLwmcDYsbWnswebF+WttgX+7MglDvBQ6UTrKDJT8JlNFrUQGySb1+DJ/QqKpO
Hlneacqt/pDdSveV1dgiH/I8ygot/IPgHRfdzhfNJ/uCpQx6KZ2sUtpbyGqQw0v9
4FX2tpbJdIZBUgvaO6ZEELBm3/AryJXJvXx1I7LI1af+wV8qqeCGOh08ki/zixM3
SYcHcJVv3IPVdQus3FU5tWl9VEjpAOoBU65Ehu07qN+DtsXlq4DPnK/mA+EZgsxf
KaVTMK7Doh+HfwlmXqD13L4O3TvN7hKEurGhROWe+8ilkrIeSpf8NZY3XXsL8UHJ
djU3nV37G17np5QyD3V+7cqU7v+q9aj0KwT3llCU4o5ezZ2rHx4ToIr1tbUyEqO5
cFhzdxzL++7otMqcFO85snhQKp5oQQ01LD9Sc+P0cXzskXA7sJejV6IpWUqefAOo
Ep3NwhH6ryTTdBPbYoUQhUe8ekuuZPx91ze0+V5IuYEU2UU3G15mOkz1aXpjh9X2
Kjp49LCtlzFEh3up8lGsNf8qGTqDfativIy2aKuTQHogNP0oZTthNce3c0u+TFy8
Z8RtsQPEegvSgMkgr+YJf7kCOGfWfRbU2Q+hx53WwWmAFNVu1/BXFugMMqZarwzL
vKI3ktDWsO1ObjDaZHaQiCK8KAGqR74zkp6XDutaxrppEqyxX9403wI+nlGL9aWB
+5h8ot0NK7MAi/796VhbCTQHQwonqjM5s5+790NrFosGj0X9HlgR/BFSOM48iTSc
/71oW/s1cTxeN1lenKXQDUtURzitXJEGj4pq2f4wXR35yDXWFseMWt3MjVFngsyd
JNLeZYMP3ifCE04hIYcfXeLd/yoTp8seqGoym4Pc+HSQLpnTPvm7VwKGuhTeJmIX
xOP6rvDmUKY1Ybw2v6ADZXEQAD7owyptsMDB9f/95sNEJoG43DY1xU37sRbhKBLx
X+ZBNnqBeFetqyYAIImUpIF+vVHDBo6hOlM7BIFiSRmGK4lT7bkVdvTC9cYZjvHa
vUWNpusQE6jxqukPCSv62GhT79uyQGBa3Wts97ukKvU3WONlF4AyAb3/rsizY0Lx
A5c3Ye0spSQL7pwVE2Ql6PgmQklrvzZc2OcxmxOZjiGHnNxrAsOx+1vr+WfBVODp
2LEfi68tKblneCKpXepsDzJX6rMkVXzlJKEWKNEDpvXUv3CUd1O9zvSpvwl+GLqq
MKJVhkaC6z/Ui7ktOR96UqamNqXNVtB/qL3mH8UPzbCeBy7NtM/2KpR1oLhnmk73
966oPazQhrEipVNoU+42IM5aQ9Eyls8Z2vWFbKZyLWh2+7U7q5kYtKFQpvgRmt26
GUKFRQqIls7qVb1zfTwIK+sKh3YbzhepEchedEkR05lsUOWpKcpLbh/JypxKPi8n
6l64om8ieBmNgK8xSjb30YT8GMQxGD2lHaqWUkp+5/iPcCKaMZSMdDC36tvyoBBb
rsRdeEBx/QJa+ZMpenkmbCXT88+aTGQZel7m3uPCY88KMxpGxIwTrBGHljfouywX
1LJM1cn80VHLKxWjwW591vVfPC0J5FCkBhLwy7XwjniECy5hYQK/PPuX/Kz5xJko
Js6mHKAfNjuKU8fA6oiOqHjj/UWveMXcKEjPx9WQk8BJzKMWWZUtrDwcNm/fpmXn
IL9sfJD92nwHxEomE6fkTNpHwZNhVt3NouuWzVxXlCk1am28aNOhbjB6hRrosrPQ
c+yn3mjWTbH3tX1nVCkGezD9BLXCcTBxX0yGgvQnr8LcL1MHMAF35vnumzbuHGET
cFr4oCbeOJfcMUKhd1N6LNyDocGAaaAIbuQ4a223RyFhI1h4HioFD7oNaL9Z90sD
GS8JN+X48x4FLsk/jM+z7w15BNWFQk5LPG6dcgAAxVYvO0w2MlJnNlrAW/Iyyr7H
TceMpow7aPFD7akVP92qeCYgyfYDGQ361pUjgsIouA5ZK0SF4VtZDy97vMDJB8K8
3aqDRXppRsS3Nh/EhjvB+Z+Ru4iz7f1NCtib0m1LYVdytL8VWSuglHx8qIHQfNV5
tHzA8M4N46fql+W1+lHY8SMo/IiuzvSOZo4wGce0pr/DoOgxteF0GFQ73FiZLU6P
ocM6gy0dd08i/L/v+nPBidtl4EC/CwtcUwPfGgm22Pme+Pac+GtVpO3yNmDAxmQd
pZv3STKXTsGgXSTxCeMu7hLUl1UmSVCE91Uovj7aOLOBV/S8REqNkkr+RO7tKpQR
qfQKK3N/eXyMLRc3pte33ov8fNTCZxf6M9xqJgoDNDfT4Plv7YHotKDlpC+9kMYb
Hp9ahjqRBQqoMkO1YEgM3Agn1a+S48E59mc7L3SJPnD994e7DorXw6h+fvsObFJD
KFokFnTkwcNXA6CnN71T7SIvy7AaeXgIHBFpbmqsVm42KpUhQ/pCp80OX4eKaj0h
QZUo0M+vRBla4jlAiUv1+sElqLWdWyFK+M+vyZ98En7wuQxarmrbINVe0o2KGXmw
I897G5/pXT1/kG3ABa3brrMn6rkd3ob/fWlluh+5y18pY/v2g9SFzQwGz3CJFVOG
sB2YOfk8Bet+d1UHwIrT8OZ/6dSOUahk1YlX4Qq7+u8U24nYXANvZXWedwrQiG+v
tJXz9XeSSIhvbnJKeSWVqIy40/XYxdXbAAD9W9BsrvmU9Dop7c/QuMm4W2dGHQzQ
jNMm4B9/yfkvvv3JYCz/IrAqdLQavQ3xBYtGsrc6zf4s25t3On/f8WcGxt241TZs
qcUpxnM3J7xaXjnwTp6Yr/jODcYluCF4V9qBZ1vaYHy0qXkiWM3S8VBkke3GjnQ9
4mzfymPbpqoGaZI+YRbaNch6+wR+OCwNeFg+HMyE6DE5B18VPZj1qojGFwZS29CA
ImWq48IFjByP+BQrLD9qwu8sKkreYzc1b76pCgz4jwPNLj+ASKWM4W0FIyJ+N/sM
d0yn0uAjF+6P7K26DicN1wQmYeJxnDbtVAQwtGVnADCWZRHoXafdJcpm1sOXKRjA
G9rI9jpyR7GYZcSsSVPqTY8F/L/0xA/oOg+U1Z9JbonK/JsGstqi3MZlpRBfXhiE
MeJmtuZg8yHEVj7b+k+QJXk151kGt+f1Xd9kKdW/zzFFMOaR5I7Of/U+3VYFO2fG
yr4L5W9Ob0yaG+iQGrvkf/ZSsFVoY4WfIGclLH0QK7AOeenOOK1YCEsMnZ9cvXsJ
nV/lCkqwhxXknMMxmd2U4Uy2hvGivouLSj2GAEH/Z/HO9FQueBLqRb6633Aeuz7y
MhZDz61AySYqe1wsVt/coTPiEzteNOyXyDuW5eonhEQL228lLaqolq8eSH1L+TJu
fH38RXmp90XCFGl9G9FkcVSLbEi/n23LUmrF8O+YX7ZfIPimpGMGxdXaIJPHVzCJ
cvaAjoa4Uj63sosGAWY37QUnwZknxhrnff9LQfYQxoIyQ+WYC2B9U7XOfQBka+02
Hpqa4VgirXLqQMsCo+xKi99enFUhtl3eN3kTW2x+NgtuxxWf0DpgqTguz/RwS8uY
F5W3JWKBaQyrD0QaDwDFdmynUNoDTx/126t1Q5RbGJ0Y2zdXG/wJfeIx79Uh0tPF
1lIg34TwkR5cqaKP5CsnAOpUVdzoiTaFq5gG5BBNi+iQqBG7hFALJs7AcULKI2hV
lIBlrIAJ/U44wZMFuiGOsUx+AcyndGPN9rtgzplsGIGwEHvpvRCbkPXxi/kBlnJ5
2Fd2d2rM4D/X63hbd1BP7tI+3Qt2ca2FSBhOr3Jsq+0yODnQxGlWge+r3yGnVdwQ
ymAvqn0aylDLpcnfRa9Zso/TpXaGTpDbtF1Ng/E4Zns7Sxr6tet2pcblYEmOZt1c
MskzL/w2SZ4YRsc045ONUIIwUeZr80VAFmeUj7Pjsq1NJRfKhgg7GiEQDbAsXHVu
OLQh/AE3YBG8N8s91ETtdYqa0rf2rtGkXAKfBR0LghBGMlHU8yUmladbvaX2igHN
uN8ZiChO5xASXB3EptBWmqW6DRe1anP9FnT1xFLy1+eWVw7uOy2He0u5LeqbU39j
RZRyxuH0rgTKqhUGoBlouEy7xkhmT4mbZEhHyAopnGEOSRRB8PFYF88dcUecRiiE
XBACWNzxi04MQSMMijdzZ7mOXPCRo2ryUafoH4FxjsWjazRRfyUGVIRkLlnh4H1J
o2ILvCZ/vhDtytmM7p26Qe662vKmnaM2AEKlrUFaTJtkbbOyYPzuUbYuoub3/Hmb
OCdXkERRnx9SoqHlM2OCP5FZY5DMkIAmPFLOw/bTDEkf+nAOMF3FdKtukUO4Mah1
2d34lD6Jrk43NErwNzSJzcIb+o4ifbf+9Ri5rnaFcngJhB1UctjPwiL2PjPn230v
nOzn31qi3oHhqe6qtZb3qm4/M7mmZl8aXH5/MNslVZJuk3qyx0gtwqqtlLmRZSKO
jFPgg7mJXL2SEtq+9PoBB3gOJ95WjsSbNBlodxhU7eFNpZBJ5527ByTvnTQv7DKK
BZgjMYubhXbOKWRd9tkbBuS49j0l6DKLhC0Q/G3bEGrYRRsH9dGyhbafp+wUiNcG
SMdl1j7tmzBk9ttKzcLusdGN97eCctiOCCKoMj7QVEJAvCBclWAmLed8p7hSKRD8
xissPP8DuU7aY3na21Oh1MRHOTK3Q6QuGkx+yPvA+lQmfBZGph1qGrR42aFucBpw
0fn49Jd9JYmzWnnyrI1kRG/z/9kRYTUbTD4IJBJadRCZdGm267+HLsDshlrNSpIU
eaVqn337Be0MtdwyDz/J/x0fYvXv3h0XaNWiLYMi/qXc2PxTRR2SuwiGvm7kiH3I
31ird71kIWFe+x/gVtT9SxgSzrryyXXY8eS3OVRp51MkGqRv0QqZM6kxjF9rMu3U
rm6YE5XDp4AeYDQuKckJuB1QO9xrDGk+otbAMWuYWnB+tYnH4L4ic1RTLeVSND9g
ICDn4XtVDGx8jkmqJmrSwITYaqtPgaaRaZfGFjVN35jZ027N3j/WDni7ZUVisJxF
keJi+zzckH/Z7HZSvJBo47LVrhdGMr3q9VUWp5OhZb0Vk37/4HdVsxUJY4i5sV3k
Mk/jHKnKtmpziJkRyc+J5ICj6z3EA40fD1zb7jvU0r5APydSH2WzBbFrTTr8J6xs
v2S1dY4t2BlQX7FMQ6wKpaIOXWOzMh9raak5gBzFVCJviCrxCsDb1fyAbshnLENw
IIbeoVWGp0MELUA8G3rrlltmxq91SzUoCVW5sbN7uoTSQzObuuBgmjnbPJF2SRa1
5kz2UqTiKaWVpsaN5QO90866H/TbVSrwjy0KnICthpx0a1LSLk1uTvZ1Sr3QRDg7
bP7dZN1WIGDzKygT6LZs2X2w7JxAL6mWGkeSgheQPvltqscuntemNUWezOHtd6Za
9cF7Whhy4ZQJFOnXf5ZD9e5kx7ARLDNwMIThk8fTxtS8lKwYY41SOyNjfY3MvIVH
AQ+AajTLKm9ANhRQepLGruSpP0UGf9y/JwjGh5BC76SdSNMd7pUqnY7rPwy+G4BS
FtyAUn8ignGacSsIAy/EdWazpOaOQNAbEwpbEZx0phpY3REKeBYl+4ZfP5/L3296
IgIBDtgwmMNEtZ+PtIRLAVP7wkTGY5X1OHXnlWKCgBGzMQQInJwj5F6IBwADFw6h
eWC5OyWvbgnbKvgTiRtjRNF4BwPym5VkwQcSTaA5qs3cx6NE3DARSXKTbuTw1xBn
1SEi4GULosKR2Du8NhZ4ULOJuXRYqOUygJrwzRCMTEfnRNHx1GUtL3KFVSFUoXGJ
cPndfH4GrsPSusNxB2MLFVMVoxlmEbKHeQ1xpsFaIFZ9HjoiKUJMuNmgVdgIT4PM
j18laVMXfXrickOd4o77R7dhUjiYBuxOaMjzasuibgKvjYJANbXyToiFt1AownRs
HsuIucKisvxj13NQfA9URa7z2yZ8X8dxHMffnaKlxKFYPho5EcGLgs64wqlcNVWO
u/0l179VIDZhgzW0d80yDcySaHXGAo19F1RWa40KP1dXiz+9ICrBm+8vwSHkIcyo
otVNQyOHb95o9su/f9S0DLfOHRIgs3hGYF3iJbt2IWtE57k4E6TcRhma50sApsg2
JZqEJe5Gtj0YXjQkEhWXEfQqIesiiAhQHQivAOxnc3fD4P8RQT7hHJ3KN7f2fPr+
+kQzXaC0Q/AftAiIV+jqaHmjsW59jTFwjCv6CxQijG/qJWAFMuMz9WPyO1w2pffC
Tu+Whc8NonhngrtjFSLnn6kts3g9mSJaZF9FdfdFnPlZmpueNldbiaPZKUvMxyZS
a5VpITWbqKFlgR3Lin91Eq5XKOhB9O3V4aDU/7KNbemcc8IYmCJdLIDEbevTyBBI
j0S3wEj+ZiAkf1tmiX7aqFYeIXUn6WvHfQ0HvDDEiXfwYY08x67OOsWasfowg7+I
ftlAnKivsgB2MNaJeL5mIlKaPpOnOBC5HXn1yAK1nBUrSc6VGQpo4sZhojGn2XGg
tSFNKpfctcfx7SJctftvhYyqJXo7fRGGj47w2vNHH0jj9mufqAghmrSH4P7lbYU9
uiKvNrgk8x9v1olTGywi67iNpo1Hm6pr6m8A1eQ776EIR6M2818zYvacy124ZNQO
AoefoVlYctsqblyTUF1ug1nWNy/df0/25+57Fn+7rgoRCN99ZwPbeq0F7U/sfB0i
DlEaF0JZAART/fBY4/Rv0VQMI7Tnia6cLgqNKQLEH/djJTpQlp9WlXaJ7R0KC2sa
HUu14KSab/CqG0MRSxp1CFw/0RCT8Fzo1Ne4Epckq91lIsEjlPQh/oUmALa4rDzy
y6SdbPp/Ux2IG/1KBan9K3iNTVE9qWg0qXLD2sqHZmXqR12/+gRvWkEiQ4YUduIX
kmwBRXlCfte1cUCvoujGLrqfw08oyyiWESyMJOw8rWrhkKRyPyTH4WELRVCVH0Ls
Zv5VDhanluo5FjRYMRET+4vtrW6UIExlT/QvuahT+GQdUbmiiHicJx7fW2tVbnMq
krsyyulsYuE913CAgCETztP1Bd43zAt7BTUrJYVvBSkaXjak7WhS4NrJw0rnQZhc
p8d+WA73h/xeL0MpTd23rh0thFFb7Bo/EkkhgxVZHzcIibdQytd6eoaOhOlsM8P5
Z39UwnaRxSjmNnSgxPRjI/U/G332esu6Q+tlj2Q93HY4ory2aVZyIwyo5M9T9tv+
ccKiBXqh6zevVCYjjcXLTTAEEEbOmoHEZKfXAxM3FFT3nDuNXXvfn3rTtrvMZZ6i
gSSpN8IPvgaXxBfc5I9PgFTz8P2ODsN9Iw1Zz5ECe5STAF3lKd6YzQgDAyv3e3k3
MzDm1CW7bMe3ThABjQa6GA==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ULQ51MPouB/XepvTtIkWvgb64Er5dkBZt6mMpaj677GTMlj1OyG3taFWn7Jikzfr
hPG03ML4M4nyzjXP7kto4R3ChPoc3CqpR+7UeBJHxv68kmtJmutJLGaC4Jq0mztH
g4Pgem4Ex+Ysu3YleGoMQmFGqN5Hf7d/Rk6ryK9jOfQaG2bf6xPn0NFZaFhq5NaR
GLzD8OGpA3ZRg9A60ieXn0XhVf+hbkDd2gDYaOvuGReudZxJzxCZLsuVlTMuIt86
Y1JlOHxdIDNYVukFVI+hiRWp4+Jjfom4QuAhnI/rUKjAsSdEw5oGuS+17iZEtZn+
oa46fFDUbE9EOf3rRInNSg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9456 )
`pragma protect data_block
fkIWfJpXKXqwONbkwDVu7FNAn2QuKMr0X6Z5ZtYGrx8cYS1DDaO9Ow6uza3uCWj5
tCkQPUPmBQA1Qlq55aEp8VZz21gfZKNtbZTFkIK5irhCKRPWozk854Fs4s0djfAp
vxlfb4aT1Qafn8RLBxyL0yPRVIeOjMhENFfJ3V/Bi52iCrE4jyhuaUHbTXNEyXR1
Fk8VzWGu0FEMB6VOBy1N6RsrGHh0A1Ms14tzLTq5K4/XUZq5QRrtniVUF0JLyc8D
AhBAuut6mfV6LMdx+Ex3tax5GNCRxVYAsTE2lvjWWy6JPppK/yMlpivSDk4OAd5p
LdAqgevctByXgvS0PqfqQA+qydA6ZBX1xwtP1WiE+8VUcxBfI2t1NDnRFxEKpDFv
JqjIAtfzuVJ45AKV4RVrObA1xAyhhlNYbLFbbODLuf9+lyxADdbRMFonpg31HEEu
yTechmQ5B7dtwDUhIz7/GZJVINTSBTqkPx9s1ycwraTpT/dY8UXZyKG9lBVo+Kif
Lghzm1GN74tsPFwIVbxwgUbMGqdCXWViAJP3FrWEJyvwgjWMR9YC/kZzhWNiuLI+
n/nz5GWNHF2+6obgIKWfPRiPkXP62HC6tU0RUTg+POlNuTo/RZ08aBiRI4ZLZ6zK
QdVLCYOZQrDRuPuuG4qAsL8FJYrc4C/w9vjkHsmqFkdjp7Hh0eyTiGjhF5+H18WO
S9mDIYsM647qaqv7NjQPHFEtgjJrITUhreNLLWNb7D3iw8ltEkCMxYum/6GIf8by
IwFvbS+jPMQJULUMhZYTum7kJ3//tjOq3mkIotCNWPa6+wGJQEgt9/XWIyjmF8Rt
A9et4F32VENxqAWU4/vD7ZWZLGxdqq1EEXtinMD2KN6Yoq5oT1QDKvw48YWCVPXj
yuFFze8SCO+Vixo+9Xw53lqz8Z1zxq0/QK4jqEkVTRoFV4LCDt1pGtWYKcyudWp5
OjBCZrDVfEddvpz4s+gkwwIvuCwglBtp1fWck5OtoEZcjoWz15YGDOgs99IW1W4B
KrT/E0OUJURuyqYAJhioKGTp5dlqyV2pvI2zIg+5ER8ig9i0LkjLsaL2tZQwU+bQ
RRysrDNTl+Votq8Bg0QAfnqacoeQ8TMMtcKyh7pXIC4qefGnjKc7fvbWjLj0jDFx
dnKgQ5kLJ5xLqiyferS8sB7KAuEVWpb7iPsHqlqhncfQb3jR0XrjoFxo2hrloPQm
MRPKl6bmrHlcgWkL4Aj81uk3y/grhGIHvt+m4UU1NZFbf5kEBwd8WbU4IQag2Uwi
wIBB0Dj4oFoOQIAifUTxlb3dMuUUP1Dt7TaWiyL6JkaHTwvOwhB4s1gYCWhKzkG4
1crxUIcdsuKq/RjusXbqB82AMrRW4+G0ID6m6flmVJeLVJXKc3sdA9BSUFnQMD32
vuvzxYdSZeZW9arDmrEbvpY92Dthy6fQ8cmFY01RrMs5uClpZChMGxrlXoT3DU7H
WDVvAv3X3y2lZmTk79c5LBTJoiVyfODsiN6PiFGV3GkrMqlysyIL6K8uuzzK+No5
QZtfeAdvwoJL6IhZm/ZcGZrTXPdpWsLUw6YNGU/2bg3l2no9u3gw6JRXFUHjJ24h
n1mKMidGLbs1wdmqeSyaR49j0TWOrUKyHFPgpGmPrxvl9OxjqrGk2Q/r5Ln/+nuv
VvDrrZQGYtJptqwHJiv7HsZqX+hw58ekORk+m6rNG97qZdL81zxGT4l7MKDo2+8e
TBSdqNv5U9tACwarCiZcKBzE8Sl9lYuStgouGM0sCLVE9Dua6uj5TI70zCKo+m4i
7kR8HaNpg6YcK9fL/3XOakAPCpjSI3ooKKDnfcvMw3ayXuIk8eY90qjSxPUX8vnX
DiXw9LkvngE0HFYNhJKFatIQIoJbtpn7J9lUHu293GbBN3Xdg9b3KcCYv35xAruL
Pajnp3NXih/cmHvicDxobglBYfzwEfsA+672Fd2bcv4Yu6sO82llaV/UcGlx99PP
JgQoTmFdIh//svmpV0T4i7uUsBdNA7h4hTbV+Tq1P1FK+IHoh3S3fuapbwhJys+D
n+5cyqFTcP8UlzIvtPLifaNTlf9jwCwoDXheYfxdx10IwLUpHXQhRFqmvuo944ps
SVo/EGEZ+gidXyjvyWg8vHGD3nVocaVvKBbGYmuoV3lB0zCdmD4Z4XfRRNkq/iBx
r6+s+jS8/uKMj+vVWTkrSVhsS5wJytRwpbHJc5mzU0i0t5+aw5DHD6STb42bZaur
KHg+GlY6GOKNYI3neKyA4cEeqUbBnNtT/Mc8toIwugE4p5AkqpocmbLpjkgYIUhx
Rd7PgxG0dz7+d8hCbOdVppmUGOohZzRFcGyC77CUADFxgrlgn5xPi9iVSO67v3su
CydjFGM4++t/8OhHD6N7V6Ou18+iHfyXxPT+Ffo2vhIq6WS6RNbqc19h5yJiRffA
XVA8H+guSzuoiWv09mfLxGZ7FgJg3gZVeM/4Bmek9V15ToahwNyImEwqFbMUHUur
W9/PK1Jl2w78BQWt50+4kV4Wd6k+WYWCUkMDJIlcRJBmI7vkZBc25kUSdI4RoTwl
FI4p5xnZ6LDodBXLJ8Ln8sDALgiIfKpBjUr13tRMQSZWbgeZ9tTPnOBWgn5EhHnG
QFi96IXs1RPyCbCiL6hrsfgBCTrx1pAqQ6jO4Y1ujFNeeFixvunQ606A9L0hs3wA
Q/s3YH9Veu9vX14Q3b3pzBP8dYQSddUd6FodS7qH0EhtyOSgrcA2diET11AwDUyA
lsV203e5pUKpG2uVT52MkvSKALGP1DIWVSvAxtATXGGhvBSqp4ZwLEJSQaK6vWUd
WZG6ap952BmjzXf+w7SxlLstcZzISRoBKz7Hkv1KdKL43AeOIHRQ9a8oEUOCPvgv
X84eXae9DC2nBCd8aZe/FFlZbBfF3Z+qhKhUs2HQPqu+W4NdH3J4UEQwz9vMswfR
qZSIcTYYNdQSQ8xnZFS2zO+ys/PrlLH7F0VY5KZ+4ZIPwAVGqrcr/2+JXMMptfl+
3GgNWmTTs/Bik3NVxmGFl/zptKE9Wfq/GZ5PLhcO9cMcTV5TAQhkJop1yFDLgxMZ
RB9BfHsrVxn1JMbcqzKQmWDuFRQeMyVa7a0BTtpHfmatUW7tPo5FGjABSqkUZJRp
UqPwFuodU/2O0vWQHZYQaSPnmfDTmRwItpX+RJuZAiH7I9z7a7eSqNA5BhTWWycR
hrTlc5n8IH9jG/C+Dm6Q6tSjauKxwQwc2NnEPUYC/gPnM7IeQAL9rCqaVj+iFhza
dXqyuZJd1ijzcoyhaMFeBKjCZnFuDP2/afuP3Md9WtzU2ktDnDo+wN82pdw3WBrq
0MoGEQnBH2P+j8IqmQZg0a0F8ms69sBe2YVBX3g5+XV9nUSn6LP4pSjU6My8Awpq
Zl7LX6WLEdxNnH5lgMztJSHYFtl5Aiwqer8tA9uVuV0iEG8JlEUHtI8FVQlRZH2o
rBaEONCNaqHo3S6hnH4rhwV7D6X0mIhmGuWbj3K9WYYVGKZDAw/Y0Cr3Q69QKCwy
AGdYH8eZMp+HEXEGpjn3/k8o92Kd6TA7emob4QH4C3AXS8D1Oc3vRqJcn36hjx0W
LkMY1wJQyRX39K4xj19wwJ10lHuxNO/9/p+OPdsecnVylD0bFUSWfTwMWXPCcpLk
47cH+MSf0NMI8SRwJXtkHdnp/FMaGofvryZ50ueEDXwexNTGvlUYBkXrWWmu/cqq
nmL28FLyD8ZyuSR2EyyHTodR6HzXJN4+vNBtM/tvqFcdeLVNpmgE3Xk39SrtZ9MN
4nqF7XXKlMZsMg/itpDxLes9hDmM8QJqsZhTEVexsVzMb25YkpHiB0ZLkKPNzilk
D/+5kZBkEPKcaxEuu/OkokBXg6p3iPSDrgelxjVn83AOm7JcUPl/7IgzqPs3ljOm
B/a2UjO69/xa7OL3wvNeXYV6FJlt+H4k9eyf7tJPhnjnwbVy3TeFJLXKGKKzP6iT
Gv8P2UNgZEEdppJzzm50ySJYURF+qp/t22U4Wf449DXrEuuGC882kogRryyMORuS
a35Il7zFW8YBWc1IMcvOtc93gjJEA9kNbw5htnNpBqTRD9DPeD5FWbzpfImq10ZP
gkvAng0dpQMGTWjWu7fOtkWLu4Ci/6oaWEvFgQwtGZ0RJgaU9IvmFfPQvpPepZKe
lo9DXl1v1UaJRyY53e/RCgAN1q7+i4ilF26utIoKenflgx33KoaS+XeAyYXwA91P
oTKXQnS7I8zPQYxvjou8VdAOASdGsdU7dN1jDV8e+opbGeYL332l30WstHjgoccK
j22x1HpuZK2O3XY9Cl+M3V01A9qbQ8ERC0ugMlAlCOnAasWbmFrVNA8b+JysyyAg
urRTmVDyhj455mrc3dfGjjNiZs+Dwg1aHX7+SdHkL1CExLeNbTuh1cKbDMpflB/Y
W8shc3egtCgotuj1pCHHu1CRlbB8ZzXv4KE3x+u6skYUqBhamU0Dqajf/6fa5Sg8
PR54Am/4+xrHx2yS6qWGVPeNSSAzV+tlgG1KkRCcVdMzEOUvsspw3E39+FKwKVVM
JJKr7Bqr51nMMoe1BDliB9Mw0FwVZuovgOFWRSxyR3kp86pIvDe/YF5x0MdRt+st
uNVkdPQdDTOtxd02LkQPpeXAWlMfht8UO3CLz+Nccf7SEWyWAeA5zAaXLH++ubJA
Ckz6x5TADo4te2PtEWwuUXUTqzvXMoSuE4i/Ympxfe3YpfK9ngxVUIkCNwCsPYB5
JsViVRuQB4ENPxBg1HeR44HizsNdDbKBlT4HYREhCV9r4/WEzhE358PYwiHT1n/C
mrUTIatnIHTVvlmQIyPL6jwcRNGewCUy57ZbytxDQd8eErOPArRtozTru8fb903X
OP75I9ui5aBth6Ll/7YkvWmK39Ozcz0/s0IZmjPxrWdWNZ00c1yiQU+IqrfUZVRQ
p0CnPSa8+n21kN/KY4FnCk0/wEWJJEbtzHLlNUvKqY4GyKxUX+MRp9XbJ7SRpMdI
P0FaJYtr+rNo/h4uaX5GT1LGoSUG4zYTt9K2ivKtVjgRSTivdmbvibf+8JM41Rwe
qsg/+PGKSQNR4tGEvsXva9TNSh3+6L614k9gR+dxEhJc+/wqWs9Fy6GDT+MI+P8a
6YohYI9/PgqHZ4ZFo9unCB6gxU4elWXL2kJvk/bSPTzgssltz1DM5OThPKd3yPhU
tIHEdPfTxD5EyN/oDg0BcatBW7AYPEeIASylVfYbWFkXXRUIrRzZ0xhxRNfzmUMi
uhnU62grYPs6ZaP5Gekgp8GM5+q93TPvfHksGEvKTEHVQASd3cIZdySaFGRoptre
fmgQeCGKutEMfA5WPZW2NzumpwquBMwafswSCJWa1a9qiEdweVdY7FGLh6lTDEQn
LPsw9Mm3KQ7lI1qgrugnjCdgag0rE1sRECtwBl03PjKolRWvHCx9FvTQSPzJiHyo
H0HlmkPyaZ8+Gjh2noWgxIopTo0gh4LOc2CJ36+q43n2AhEgs7m25XQ+Mn6BATp5
+Fl+tbsrO6qcHTifIBu1Ys0wUCWA+blCj3CpPwEJKBgtl2bJbIw3bo3BKJ6CUPJO
7qYmbuV9E3rH+i0WkYya/KwpCKP3E/g3XJgyWbJjbisA/RIoF/9thFMQl0PlprbO
78H9X++mEAH0n6bySGHsEo5Ofx23c8QjiRo6jd1wqiibOH20cKYLz1QLDK8IglUA
TVbnam0CD/79TSVWztXajvsaJM0vHgH2UJVo7G/If6Cf7yybuzh+Lmeb0PybQrpL
Ol8WJeW1JT3rGca5BkofiRHAgIzbPTblYSsoYp1acoBOTUIDHEDYPjgjfjcYpn0V
+AozYS1VfbvrDu+mHyelTMv7UQ1BSkYjgGB06a2qGcoFZnOKKN2y+yc0CFLBlv6c
dKZQVRinkWxZULunX2Bb/w/jOlDslF4xUiRzuLYPu2pDzJ+IouTUeUwvm+IjP9u7
+SEpKu8IEWBmp2WXgPsgHkWQJ3+Y0ABi3qm5DuNY9DJYdyflX3BBPjNu9zlSLYiK
TGQhdCn1iQYZFzgJeXrZ9ctmT3My4CsfoLuOEkEJ+xNJes922E31B3+n5eU7ptwR
AZc6S1AsMO6nAjBkrs8fH8hn37DnVkLk9f2Qc6lFv3ug0e+UU+9QodgmZusC+nZK
J8Us1Yrn30AG2qWM1OrficN6YU0ogvwnGbgeY0eIMJYYYCayxgXeW+IxAQCMW87w
7Q1RYvjIJ7kfVeOWPVildzZaE0nRufmT3oRVg3pIPe+hsevPsLIEdh8tcmGubTF3
ruCW0P1hCGXpGmc6MtdPn03ytKdsfB6HS+uqyqvC7VuktVTAVDH0F4HuZoq/pKx/
aMbiKhukGsTZUsILxTC4bHqZ5zdqV8LC5NWk5kJn/WwcfrjUho+CKQkFT0l7EZPM
bzB8ywzhOcUZtWhVUBKTBgTNZ+UQScS5C5tTMauCbz+mA8iAX/8zw4JqiWWv1B/7
7iG0IYSgT4XoQmfxEUQdDyq4XqclhqulRqpnJrVXrMYNhUR3E8I4asV9ug2koeMN
mFUJz+YkaKt976pAeMZibMAFxvIjwhCOjrAaEcm65WlWK5lY3qCSFRfLR5NnJbKt
DbjsgLs4h8CtN/BVxkedWp/v+cAD1tIuwWhJ2K2Un6tDCMz7DKGFLx05SDfgTuBK
oVmxyBBs56yUj6mDKCzX0UEH3g2uMhRrVfRdVMzK4lJnwvDF6bmEgxJAw6zIft8H
z6kxS4fYuOertfawnxMHBeahPTODKDG32f/yIc2DD0SWSZeVzbeDXgW05mClFPBA
MmeMHEPGlesnUNpil8QJg9HvNSWBfKo7NA/ddUIEnsnoB+R4QKrXhtxMegamG/z4
RzDRAWoRcUe8I+cRNzt4zNPs1aVJZXN0JqXo1U6TaDew5rIZayvXxeSPjJmf3Uie
cTBSCNko16GEDhNn8QU5j8dEFbNB+XwltE32O6HMTQgH4uQTJOBQ1ErD80zRY1rK
qd8dLccGkkHpjCBY9NeTkwN1Gn9qF1l0vSBwxxA/F4D1Fp4K8mS/RWrTlwbUnQoO
gQ4PnPOZ1NowMeH0AxA2oYdoeERmdI9+rOAxnrATychy/omgOULPH4M3oTTw7+5a
3ECUOxd6dqm0ORKAQcMAifB+vWdiV49Iq7qC+8IIKPBbLFFyTnp074ry/Z3g5p+0
iz8NaN4CK8aeoRuWvHmP9DDQeGM+sEjFrVozhE77A2rm3xW+FJtebzmzrvzOd04I
r1shklECjdIw8RLzxbpyM57FrujqqCFX2ijZ02+SGF7JsE/iMSq/CIhYSBUISTFr
suFiCp0U/XM6tBHkLUPUwAsCQZK6wXBPdSoxURiZRkw8zyKlg+fahnccrawzhCkL
CepHBqPO+c6qQKQL0JWWGO3ViPdabyk7ulXAJK/uM11Nbq2EAc5mD4seokSN4k27
I0znBzmD+LQoSgFYggDboyW1bN4JAIlWTNfHBB7kJCcRpSOfKGyiWxjnjFuk2ald
QU4SugG7BtOD3f6cV85sStUeU8UqZ4Br81FiR2Gjaoi9uQ8FWlU3k/z8Ib9gVRN5
NNYAeKyb/SEBbNyJgBu7nZR4b2CmHvdsFUBrjjx+zOtoSo1PHSRt8CqO16Xk2Uf/
12WNm4D2hfW+LQ+Zvs2+mfJgZ9/8L6Ap5Gb6+7wEl0D87cMAO8f+QqRA+kRdOJ1G
kqwdJbHG2h6Gid6Gx72vE0k6OGA79ZLmv+dyiwHu5cduKHLrTsVHpNvK20LRCOrO
BzvCRFZDiPADZQuVr3qy3Ec5+Cd3mCjgo7aYYBgOYzA5ylloKWTMzCRKViEByswF
HreWZKZAOXPrsExewzHAKIHLgLZwqKw6TB5eDbQTLXDbUqdrmH5RG3BxvQfF6zSn
TAgmjMX3b5Ei8viXVyfyFUICvugPS6FQ3ckSH3yZ3eA1NeR0hmHNGC6oliHp81eM
Ye7qRN8D1BWgKvfqZSIEkhYvaUJK4pzdHKXSmaWc3ImMYR39i0DAnhebWg2BWd3Q
JXa5VKZP2fiRtD3RP6T6hStmagdiBwqwx0VbjToPZMr3unvj4eFX97+CCwoIerzY
c2tHrZTT0J/Z5/2NMurui5C3xOu1OEkAIVPANZR9S/cJG9WQNNgfHTJke+7FacIh
nQxXsMZLtjs650/IF4jan6w2Te+YvK+0Db8mOTf9p7f+WME2yfPv4QHB1GghQ4AI
aZzx1hv9FAvlh0ISUAAAXaq9WuSfaYAY14MxFzKKiITOnse9uy5TpZ5+t4bLjEjH
/MQgP3kBxP6+nmHK/tuMlSXL8qisLNm5Bu0Weaz8b4sgoEV7wRclcRS/y9S9RN0g
3se0/MaCSoVP0k1N3pCbNm6h4KiKSxXkn9wqg2i7mf89lULhBuUG+LElTG3RPbAy
zhzG7C+Tf9OGUAokWIWqtEgr72X3tZnoc07+p9lrLByOipvVa1SNZOQG08wLK3U8
G3WG8VCytRPoUk/wiqqlsLFeQPqYZ1urqQ2sXXS4ayugfyfaxkCFtz46JEzXRhhR
fzMkC6gvGVf4XqHcHCfmK17FBPJ/iAtF6NpuwamiVUtivnplI4+pbfYZAEUaDQDK
r+Qz/Bp0Isyk6ynhEm/r9v0ck+Qh1TsCzKDxixmXYuXM3yXO3iEFodCJDs3o4YcZ
mHRe2b+2+KvKfgD483PYbwids6R1VYz9xpjq5x27Jo5s1+W+mJTMaeh/4kV5xTeW
YxhORUINbgk7qzAz4K7MLgnHSvTiL/vs3OQGs5snT68zY76bBRERP40dh53+xto7
dqaMpWv25UBA/AItnCyeB69CEN+H+BH716Be1sBE/JVY6qbbDHme9uOyzFWmM7h0
gt1WVI1zj6jmL9Zv55bjlKNHQix+8qlJxY9WFfysB1JwyEWlU7uUTbUFMVNx/FwD
hstqLwirtmqYGmk0fjten7eQJFQVU4R9rdv3ucysa0JxE6yLkHgnK0hTYHPCfvkG
Q+Bcsy3TouOAco4j+Zv+RAM3okKSlsx27TURFJzYhA8U3emfz26FsyulSi2onHrO
jf+Ml3jGKSx4Zo5YKvbKqe4YtVSBUHbNMpXErOpgccr81hu/BLUubFKM0KkN+hH+
nFvlF52LZy6N6KXWNqxKPklfrDfaDe2H36GEGKVC68KD8egrlS5AgNXllwiKwgyy
+JU6SCc7WvJhaoRGRW9DqbhLjiOVEwHJ2Kh98DQhOEabbOj/DnFA+ygI0T7CUkcT
sseDbOIUtCaoI3lHVv/Y/8hQp6uBfHvYhyqXrrh6EOecvmMPbwQWoG+WMZ/XHTDZ
DgTFqR9bkUTUIcz9eXkN/31zJseliMnp0TNJAav1DvUFE8vmXbvhL/L3cXQKhmFW
5KSVADffn9uJPCj/YsKOy9IpIa4TuwVXa7wO8OVwDxYNQiL528phVx4u9Z7I2enG
aMK7GL+agxIoriW42FS49Z6hAJmh1Hd4RnBYZsbQs5HTE9Rg42Hd0bcc9+ob1BRS
glLTmXCFbkxYaRr+2bCkVgsgHeTPXDVmkaYy193JYFwQRZCdORv6AbQRuz7gLrcU
j0fyterZowwmRfML6WHnzSo53WKMCiBOA6+ydc1Eo53NVeNRuefFAhJz4fWlmEQD
Y551TioW86kEY07wWBVTyax6s+acDl24mXk8iIn1EQH4D175kTT/UbwEB95tMVBK
jGGlp5J8iXdri7/Qj0hPVBbFyv4WWGi5cTmD9hFuJPw8EGUgsgxRAaEQYrXrlRAE
4PfM5zV4aoBuNmZ8IV5npXKhlfhHVdvEiiXs8sRz6U9jiSxIggrDxCfQYct5Wbx9
ErQPln1mdBCOwpaW1XRlqwDayfBu7EGzjpyE9Jzkg7JhpYDqnK9ZDTqa0SK34syD
nvQX3XhUA29tvWDU5cU3oAlOkcP6kBNczAVkgWZXazLMOY5+GYtISLdU8bDVPo7S
j1preBw3cpY3PrgnbSY7teqTnlZziRjJ5RB+3QcReG90egNsfRwlNbWmWATKcXLh
/Flm8GiTF23mYYTyJ3bxXEozO6cIlVn3C4AXIwz32wrBOEzfA2ocUEfPehstwMXT
YEfEZSxmPh1x8zv8lQ+KeXlhrx5gVe7Z5ti/yM0t+mRbwk6mUoxeOzodJ0VAWS49
meuEv9aNicswUc8QnLgcR62Wi4VZAgO/8X5yV77XDLp8dPT1euNp6HMaRbg6bOx/
PQWTfe8MT4d+nybt3i3Y5LyzSn9GVZOJBDKZ7aFejRfaa6W9hlR4U9XavQpLMulO
0PNvX6leJxzJzWOfsfcXykT1UL3CLFPwI5oZCl6aVoJeCLOnxOrBO4TfhGIbaNXX
HhJ5a536s6nuXCfuqvL0yii3l+7rgxemlsymfBkIOoZPC86p9SGdx5tRv003B0Om
5m8aVZ4lwto1NzIykPfI6TI5LcN1zOc6MTXcqhERf1aXwcM+Jd5Du4rEUkKmOM5a
fiNNOiE6Y9NUiADvsY1D53u++KZvjeik1khXrmdXbpUDV0wniD5rP8ry6iQBZgFw
mZ+Pox/1Bd+mtqrRaE6dn2xouk17KfMWcH1DKN1oURNmHfAWNBvlA0swdZUTkpcM
nZ4+95izepe3EUG1RZYR39VKv537rtwl0HThutfLB5liRNxg11nXT8XM8owUyLZz
jOX3P0K8ccDMFk5BuF8kopSQq2cnihaGTxxiHu2NO/T6TqnfP4KviMybVEV1HAhX
sRLEWb5x3Cahs3Gb22NkUZn7aFea1Tre4HF5vpg5Ipgi3d3EMkvaTWpvBQ5o7Vta
5qKW8eK+cazwEpGQESqxx5+9X73g5yhlKtpsYXudkLES8K+7knPje2/aG4g6WMa9
dWTI+xrACyWZTQuB4Hsbi2sSJdZ2Wkogy/hRJw68IJRPb/REgEW5EvKSOOUxDSlz
4E7ivWshTk/us+x9NelO7LRx4rCWv92AxaxqckJbJqKBC0hBQJEmKPL5xNEAaXXE
3R3uXOHcTonLcT6ZKm0I+L9OlAG9nJOhTJvA4wV2Tu85dOEFzvWZNufaT5f8BK3Q
YzwQCbA7+v91IdYepvJDyYSSb+JkPInQfXPgXzwaPeC/w12u33qNCMBQpR4cxjfF
LfhgSo+QmeSuUANrAjnjKHBlxc21vh2gM6JDZfB0qMjdBBndtbs+c1aXS1FhPnec
YrdolvSQuj2B09X1NgwhNxFoSrF5adRFmeWZbcPiNb94f4s2dXM378xtaasj8zHL
nFBXsXMQiTj+tVrG5CuQ6ZNQXry/2yEUQWy301ulQUuWfnT3eqcykQUDKI9Qgsx6
Jb+y4d7RKI65otYd7j8IPxChWxT2jfHYgdL2XkEZhomckKCy729molYyzOnLRAxv
tcr1Z1owYN2y8sIQbUGe39oYd/kA6blIHlIGnYG876CGZ2VX8b04hkDXV8I3CfEj
rLvXpMeAT/7i1dxM0zQSPRU7usd1qGlEDdaiT6RGtOYSO3abWTTEBXMS0McFyQ4a
XWz+WChDva3jbFnxfv0l8C1CVqs55v8BdNHe55y9zolNS1NA8ei8hlmbL24g35dw
ZMUju1rBoY6/1NGkoNcDz/mGHfxZmxY6b+01WoEtXJjPblqaTUS/l2EvCFTkmHfR
av2MJwpFpkXB5ZKyVeUunzFdi//+uKVVgQVXER6QGPKSP3dGs7PVA2dXMeA0mWdi
KdemdwluSmL8x44GyHb2W7QcKyVdDK66niw3OQVAzCqZAaFtWX+gs0cmKOfe36JB
AN5ADSmrw59ljzAjjk6pt1rCd2VolQhcXlpJy8qjB7nVX1Z53rC3EVeI5UXHmpVB
XNrLfIFNwgVTiswppl+r1b1Ue1cVrcSDhHthKbKuKAwMzOUHHiaEHs6GqAMNHy4N
IHLSX5ad059p3iec86yUN1oUKUOLR71wAHQcyNbzDNB+fvGcPJvWBIxFh87/XJSc
O/gMM5E2qU2muYZ2dKFqKHPc4CsTQgTnHVtjQsCJU3QoMq1UBhOBPoZ8/v+5lyzo
k/XrtVH7kLnrqhwOk5hmO5kOloOEI+94YrXAZ2Ulg8XAMOXAFQ6WRV35x7xu8yvg
fBILEOFBG+9hpheYgITyscQ9kSTrCt0CUOBuJQAw+92Tl0a6Fu+kKJl6Vy11AfJe
891Je3erc42oOGs2MpkYzd2GNtWJHAI+HiekYnhCtu10D6lwxWZ6N11yQA4vWtF5
hPKzWSPzuIrRFBu9lTG5Uyq6PvwVOPuXaX+GIPbGNxUS1hx6YVYJtzAzoBUGWxxJ
G5hQ9vE1slKT2IXwE1/7IxhEdSciSp1E5SvRaAqQBonuAw9qLr8oL9+TmHz4J9d/
YroBYc1O8o07koeKmJkh4/uOrJuzzopEWeWO5xvfTL5n4MjS1wclo6B/h38JsWbR
9/1HQlxksLdenWcoEsEKPb8UKxkCl1/2Hc8HABMA+8LUT6XggXrrd03yqsMS1HJi
Fre2cqUV7Yx8lGeG8z/lDnOshjP1vHyqfnSC/+jtvbywJqVyFdEpD6bZU7MuudiQ
qpZ3rJxsUrs4wJ8e6k0P2XvftZioqwAkG7c8b8dNcKeY4k8oI1F84zCyjbOMqfr2
7b+xvoAecwZFKakeYufgaBaGDWOkQBAgUKYbh8cZ4TqYxgT2vf+7UkZR+tBN6Zn2
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
XbFl5qGRNV788/G+wTigFXjnOBhle2VWZyVZs4jTGY+D+xMsmpjVo2uK2cnb4rUL
cql9VrLasZe4UtjnoGjXRubz7kFxnp8oNVA+SF1DaJvB05V2RbzqiAD2NmVoSm3y
anvQtOKghMPuttpR2kBtwOwsQW5ecdukEGewY6lyUAxpohOOWcdLz7UlsXHixBct
n1OJa3sMqHqt3cJl7RAM5gHuNUwOLpvySl2YMFJHpYyGodjeW/jLWFA1GJJBO5Vd
7TgJeBuxjGLQGt43YZPt6L0+gX/O3Xrdq1KzsVc6MpoiHNeJz4GvJmQ3zQy/Bh5j
yV0d/f8/15S9+KFKO2wDTA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2672 )
`pragma protect data_block
iyQkyujt6HSu8oMLseRFbjhkIMkUlI1LBrxMVGzL5lV3MD+Z2Z7tIGXtTvd8huCY
mI+DF6Vr1DCV55wzAkvjn/MJOhThkQhNUSCRI4C675UHWRcqJeCBTBguj4gBZgR4
q/eRYJlAD56/nQ4lskUIKc3ckC7wP8iiZaaeKblv80g5bS0CV/UtADI+Qge4Vt5M
rQb7lLBV3Nn+fqR5DJvzS2xxcabsd7Rw++VBpkrJKaEcwB1aLgttIXmkJiFlc835
8RUNuzMo3J/aSIA6dYUXcLcm3WHk1QXdKf/UgCCfB0L8zKeR/mRLAEvBnv5rzSIp
BXW2ra8KXLUoMqEHypoXpwacbntGXch8PjdiPzHnWoRWKMhP2XZaeau9PprB0kpJ
t+WlereQBJhhV4IiDAWqv8qNoWdRztgqz2bWuEACr5ok4rgsChojHrobnhFbhTvO
7Xjfjx5C1+8EBxFOXJVzCDbdU1Ce1NU59A36nZu/4iPF8D+EL8hEZ2MwSDP4IyMm
c2f4xKUGNCNWMwrp6YdLIemjFWzYFdmosEb5vM2fON8XhSnxy3IOQUofx5JhT7BU
1xvvFsZCOGG09eBy7ma9Zyr3if6QOjk3V47NfYrJwpKO/pWzjpmuFmG/zJskPWSl
ZnSSj/W+h1FdVYBQggViwQt0H315jP4GFy2BPwAgY1Z3JTOOOvzwlrR7+hewH73v
mf04iq/hy/8KOgcSXbCLf1/8LCMQdNoI/iaRJ/ikDVjOQ/ClcDQNcM4zthU99D07
PEEVlTO19+w2WpMA4yW3EMw4eGmhJari3sjRbbkMnT/+uIDOEnM8escPNbl5qT3A
Snms9B1xGQNeBtLbiOWohqUnXg1AhZcgBmVFUNy/m2d2Lud4u0edErFYAWiiWQH9
CgT9LKPCdMrMOB/+VzAl/646XCon8Aj4e1SuoPFuKQ/p6VwSmsxsQVsdJ+BNSEqq
BaZhdHrOKAXOPw3u7p3LviEuUe7PkTm3yYDLbTbXWsiadjHuTmVXlCZW8fXPejtP
hJWXj3tTjarm8nMfO4SEPbp6xRYnH9FgWjGydWrEhBVq3PKwq03z8x1TBQSzql+T
7E/95hufyExVtevu4XW0hcRYMJn6iWx5Lpe41JYAjA+MpTcDJJhmcvz/CNaP5Gjo
P63vC89UaOHMVRvhri8mzKyDbFCIkawc71s21uqWNgkPkSvfSa6KYdNl8lONDGLA
vWVTxXWCgM50YMWPBQhLFhK5zW18e9733eqlE2oDWGIpp4JN+aG0h9ecuFHxsGVp
mC3ldpP+c/yPI/62ILrY+1ubeyWViAX8t8vbkCaAGwqFeAtMsxc+JBMYZH7seEMZ
+l8SqJ86ZFGeMxF9xpPwWTYDnyIjNbqLXT0wLYV3/exCTpW9g7FKoEJpVPlnb5Mg
UBoaFeHHyDt5EQW7RbGwGE7ZL+y3TtGBIX52Fm1PRQAgmHCLJyw5B/kyeVfQRK4l
7Yp8QcuRDHM13tCjIUekVyxb/VbVpso401mIZ7NShybyBOzfEqPB4FClrEhSUdi0
Y7pWLWL25QgTcNUzZKH3a2TCVBazXa45iKbgWObktsvRJjZNAUniYoNrpWzx19Mk
PxP3B3rMM1qaPPVU7MHvG4o/S+V4X4xiQnoveM+afq0Y83LgNcdhQkgKbE3txzqG
8hZrsI0l88ko9Z9jnd1oELwpPOpcySK8ZktGVveGTZ8W7AgjtGMya69t9BzGTJbd
slOR6gYgf0BnV2DnKBcDqlGVytrmN2vnVSOOVm/pkWjUwptH+P0WNkIZ7EslTYgw
P1xUNunf6QMk4yvx2fYWa1IYG9/TbV4zEocWBMBv9l8o5ALz0ovAniYGEUiLZPln
bWApnqBxHuJKZjNofkO+o+riB0PAb0L2XT+GSEBOKHvnczc0lNqgEpWt9RC8OnB9
2vV4P9YXSjZ7DZZs2krmPcmLiZ+gu1gt5cPlMH/j4yIoJDEts/NB5KPwSAjiC0cE
DemQf9kh2cZKhD+qZmpUPH8WMAOAgQR78XLE4yr2j6l8Gfxa0exUKm0pghvOvuTl
bctE6HfvSmBSpOeC7kk29qRa+nrNw4KTV23rR/fcTmZXZYLtiBWinPrT5s7EyQ7X
Cm6vGJA3fIBNJjUFaBcknejcPYJTg0Ads8Bvn8DroIj/ndEqZQtZ3VqEfMlQUv5C
qDdKEOV/DogGQ4bGpoJ/TrfP7YfKQApBekSKxsud+BHWDlU08VZaCBfbKFMRFVby
kQxREF+f1Bq0xEStkCaIyHX+SiZMDUpBmSNX913jDyhfXNEI0a+lq21tgsDbFRcS
xCVTFIU5T4+zTpxZgpl3pxzL7UvdjaJaq/yV5xt9DEcOOoaEtEUe/U3AuaHkzlmk
Kn+6Y5uXYEo0VSd4VLSgRkvZcf9wt2a1wlmOww3KEg/XiDBaZtOSfX8JKpevMHmj
InJNfc3OI84piMI7oMejJ6ElFrhqdxMRIaH5Ro6WXYZy4aYejvlFrvgm06wJw48B
5+2vhQ/fN1oOpjewLZkk47f6vfviTaD1fkSDSO5JBXo4tnxDVZ7WfGgtSh7MZ96d
BXIkcmu1cPlyulciDarYnp2amPbssA6jqVufNQ/8ehvm9QQSEoWXEUoGRdla4WV9
I6PKMrtD5kaJbxv0nQSzTWZUqWTggtpEBoL9DTkxQgm40CSC09gCU/2VTy9k77fA
EietlAPBNogy8iRosY4cBzlYAj5yhfsE8YnEKqqlnefM2B5M/gCRYoePO/3enD1R
K53ToMhwr+nHIY9mthgQ1GibDp/1wVVU0gIsIXlBhQ6h0WojYCSof6CzJy1LNYIX
qePzaWVsrEfv1o1O7vCDJ8lDyXq7axVGocAd1H/8ppH4ijwNVPbNDemNUyNyHNmL
OiPMDED92jJa1swzgofHDqwGx0ZiWWCV6HCMBKrXRIndxKq5V9LVoUd/5tEZFuAV
XSO6bGK7K/QhIdWV6qh2gvoQjk4JUzdy7jn+MIp2+PQQ3EgTIubFXviqfZ5agHZS
JVBJK8txkerenO8yVWdAiIJOeg6ybDcs3X4mjgYi9Clmqy8augOtpMNo7ZaRJFTR
JeWn2Ns/LCTTzJwHKFCaa3o39bGgJ+kpcMvlO5zXOKJtyyKTIXpiqjtJl2e1Qusa
YNra6FSESh3HTE/rHqVHdOHuwpFV+Vg7hPFusfqKzQzc2momnCOuPn3limqifVol
fCeKlpDOlNDZ8PaYpoxvAqtIJ5wIj/U3AuTyWKsLOJXGDiF8roGCUacYEWXW3EyH
c3q3H4z0UyT1guUFOIVAnPN5q2c8uZKoc36s0r0wVD5c8xlwKQkmSF/l4QwdEdb+
O8UdAEu1PNAQIgNJnzuXdNqBMCF++kUy96gny2aLa1nbMfeGIrMooPTtgAtPfji1
SzuMJ2TgwxFA6e4Q7nBR2ORmxniUoN/GxWeXLf271e23oOjcFUe2Sj99/zjbth9g
RQ5zTmNRSnlppAO/qdtuJu9ulwNXUDEGFgD/415N+a/mZG7PrE5u+iBzOnNRMlc9
OtQTFVq3ppc9UhL4qotvCZnWrulCl3zg7CqwAKzIDwc=
`pragma protect end_protected

//pragma protect end
