////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2022 github-efx
// 
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
///////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ns

module slave_coupler#(
    parameter        			    AXI_AW                = 32,
    parameter        			    AXI_DW                = 32,
    parameter        			    CB_DW                 = 64,
    parameter        			    DEPTH                 = 3,
    parameter                       AXI_WR_FIFO_RAM_STYLE = "block_ram"
    
)
(

//Slave AXI4 Bus Interface
//--Global Signals
input                           clk,
input                           rstn,
//--Slave AXI4 Write
input                           s_axi_awvalid,
output  reg                     s_axi_awready,
input           [AXI_AW-1:0]    s_axi_awaddr,
input           [7:0]           s_axi_awlen,
input                           s_axi_wvalid,
output  reg                     s_axi_wready,
input           [AXI_DW-1:0]    s_axi_wdata,
input           [AXI_DW/8-1:0]  s_axi_wstrb,
input                           s_axi_wlast,
output  reg                     s_axi_bvalid,
input                           s_axi_bready,
output  wire    [1:0]           s_axi_bresp,
//--Slave AXI4 Read
input                           s_axi_arvalid,
output  reg                     s_axi_arready,
input           [AXI_AW-1:0]    s_axi_araddr,
input           [7:0]           s_axi_arlen,
output  reg                     s_axi_rvalid,
input                           s_axi_rready,
output  reg     [AXI_DW-1:0]    s_axi_rdata,
output  reg                     s_axi_rlast,
output  wire    [1:0]           s_axi_rresp,

//Master Local Bus Interface
//--Master Local Bus Write/Read Address 
output  wire                    m_lb_arw,
output  wire                    m_lb_avalid,
input                           m_lb_aready,
output  reg     [AXI_AW-1:0]    m_lb_aaddr,
output  reg     [7:0]           m_lb_alen,
//--Master Local Bus Write Data 
output  reg                     m_lb_wvalid,
input                           m_lb_wready,
output  reg     [CB_DW-1:0]     m_lb_wdata,
output  reg     [CB_DW/8-1:0]   m_lb_wstrb,
output  reg                     m_lb_wlast,
//--Master Local Bus Read Data
input                           m_lb_rvalid,
output  reg                     m_lb_rready,
input           [CB_DW-1:0]     m_lb_rdata,
input                           m_lb_rlast

);
//Parameter Define
parameter                       State_idle = 2'd0;
parameter                       State_aw   = 2'd1;
parameter                       State_ar   = 2'd2;
parameter                       State_done = 2'd3;

parameter                       aw_State_idle = 3'd0;
parameter                       aw_State_aw   = 3'd1;
parameter                       aw_State_cmd  = 3'd2;
parameter                       aw_State_data = 3'd3;
parameter                       aw_State_done = 3'd4;

parameter                       ar_State_idle = 3'd0;
parameter                       ar_State_ar   = 3'd1;
parameter                       ar_State_cmd  = 3'd2;
parameter                       ar_State_data = 3'd3;
parameter                       ar_State_done = 3'd4;

localparam  AXI_BURST_DATA_NUM_WTH = $clog2((AXI_DW/8)*256);
localparam  CB_FULL_BURST_DATA_NUM = (CB_DW/8)*256;
localparam  AXI_ADDR_OFFSET_WTH    = $clog2(AXI_DW/8);
localparam  CB_ADDR_OFFSET_WTH     = $clog2(CB_DW/8);

//Register Define
reg     [1:0]                   cur_state;
reg     [1:0]                   next_state;

reg                             aw_busy;
reg                             r_busy;

//Wire Define
wire                            u1_wen;
wire    [AXI_DW-1:0]            u1_wdata;
wire    [AXI_DW/8-1:0]          u1_wstrb;
wire                            u1_wlast;
wire                            u1_almfull;
wire                            u1_ren;
wire    [CB_DW-1:0]             u1_rdata;
wire    [CB_DW/8-1:0]           u1_rstrb;
wire                            u1_rlast;
wire                            u1_empty;

wire                            u2_wen;
wire    [CB_DW-1:0]             u2_wdata;
wire                            u2_wlast;
wire                            u2_almfull;
wire                            u2_ren;

wire    [AXI_DW-1:0]            u2_rdata;
wire                            u2_rlast;
wire                            u2_empty;

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="ipecrypt"
`pragma protect encrypt_agent_info="http://ipencrypter.com Version: 20.0.8"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"

`pragma protect key_keyowner="Efinix Inc."
`pragma protect key_keyname="EFX_K01"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_block
CsnhTznO8x9sc7At8ZuVw4FP/dy/mLnJ9QP5L21jyKWivijmgUzQz4pDQsgubs9/
qh+YdoKppufTD0iT+iCBY9mi7Q3SQfklDTVS4JAfovnd618CuAuvkeRAe+hr1tIz
kOWvI3RbYBRNy+B/baEN9WI7MNsXraaieeWF1lYKHiNEQP9c4oTuNV7o0pm7X5dL
NzUwvSQaQnu9AaIORfotR6cLMLpTk6mID7Dw8rDJckoIi9TKbIiTQP8msW0MPPL3
l81KNYoP7IUPIj3PO9rq1kVmnIyOYWWjTcuU0CjRJFGWiKkAp75NfSnyVIM0nhhJ
P9e5Kuk0CmUqtmyIZ+gkiw==
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_block
NF4H+pcTafFDNfb+3iKgqTH0VhL4HX/QkJbp4HIr9PS+5Swj3AAo90J28hkYU9uA
rIN9V/IdfUdP0wpaAe2CIaHT1Xf+YVe5cWunMyXNM3DwWmI8dsziQJI+B0jUSRjf
CfdXFSD34o8YaXLHQoFpiwbogpt5hmouugqKw9HjLKs=
`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=31840)
`pragma protect data_block
qpNgCNCksrPEltvuIwAWirlvbV94XnpH0JIinMXV6avIqOqgcVhlCvK9tmocIWJ3
AGXtY/5kbnPFmhH+HwgIs2Lkov31Nif8VCtNI+2I8RQuIx46VJ40TB3n6CrX/Bwq
gdyoIQfFGBR8O/+OSIP69DLv6ISPW4LmCOoPXM+WTlasGyPqcqn7jvB7ZqveV/kJ
6gM0Olv7aDoz39vuW/fpD1gxnyxIqqJ1XDJBMKly/Q21SOoY4Q8nN2cDl4yYjWbL
ngaS5c9VKyo+J9SKVhq6YAjAHjwvgowUkeUfKWGT4QjuacMgBAiEycpMM+KV9HH1
gYq/4Uy0Hy53g7ADfIuqHiPMQVQ3PShGoGWkOYcan2WY+sznQve3VsLJsLu45HqN
dOzcS9JYVe5d6yuV93xZyYRWHFI3l8CJHEh45zv80xfcGZqxfC3arEkWIOGbdmsl
YJnulIK7u60Ep58a/K8L7tlM9e4jWPC9IEIWkPEETKePu+0gKx/EFFOhMlAGPyGo
xtXNGwuFJ7nrECdR2ROeuWcaGFkPGzulsnnG4lGERpA60bPwJAEDMRahCKeyVBkE
WUv8gLsaMJkFDOc9c5yPCowqhe2PLT0j0h6sF3N23/EMp7hr7DGtCnzDO56tNEiC
rT2UsRMjGQdzIUw7G9XsUizvpo3xJpMCieBBuNvrVSrCCnGrH90dl4bifiN2sXJW
Ps7GRKh5/4YDxGdw6GnbJolHg6/qLWBOUx2LbpHEIcSqkKqxfbNovnfChcO2OG1A
Zk4O9mYa2xfP2xuM7a01LGBneACxNBAJFfEgJy1sRhxCtit8hCXJ2GWexbyd4nrJ
ao7g8hurW2ardQuG6GagKMOTy/lOK4H2XrFC7on1RQc9I9C7N0iapB1UBkfGdFis
ILWK5n/Mh9Lg4nGbYryv5Jo0UNKZzLu6NUJAFGBerCK9IASV4qLNcCOWeR6et3+/
jSR+pv0JSinozFDrZi+LJAIH8eh5p8hkUb9fzM1YCGi/i+qXblvTefaBrbq5lgfI
QXRU0ozxs8BC44Un95kC5t9a8nmnuVwvp50HPlGCG8RgvCgRWChprGd5FqAQo9PG
9byVSUEj+uwfhLIP1k0hoIxwVxQbI/21X3xCDRZ/hvFKsDGE6Gda9PMahvxpgwHH
IdBq3gPyMk+eywaEgiv4sxvxF3v9CmOZnvt5WrnjakTL/QUrAnbwAEs/bo4AQ57y
rWIkkQFTIVakMQa8eKoYkEbLdolPBHplltw7TSiRy/qKfRrz2kbTT/8OPVw+zfXb
t2RztdwKffXcX73KqrPpWXb8Yge8PJO4XVFYlwkbddJVpWMezZiUhbehspUyT5ep
PD9nuZdpyZZQ5GnhAL7WEmxZmMI9I9qtAY0vpysZ9G4KRVQK5YiZBaBwFmW4G+kj
kJatRveau7q1AXQS0BOW6VCNLjctShgEKM6Qtw4hQ9EgtKa87wwvBKVycTPjfGcD
3Yugtx5Q8IlKLmQ6jU2Qx3KzFn+xB2JRmnAWwQ9pVU932n/c5TueuFIDHp5v9EC4
reUR1/ZnDDTPTZjck2VBZtinxnExD4zVzHGO3T5Oao6SHGo/Jy8vy26d3MLjJh08
6BK3u9zymcQZWVct/Bw6ni4FUFbdyeAv+79Jkdo4MZwVakkMEWs6i7jeOLbsy0K1
tRYNDZYbDHauPMfdCigIrLMYxoWn5pGjF/k2LhMECOeRotTe1w7TUxWaWMRIQUA/
pUVcWQT6cD7m+7kWuWAQR5XDgYAtFllBvBbHyGXxkc1JoTGPdw1Et1uHDUB6gpMM
VIRv5vjN1ZJ4EYQc4TKa3D/FgP6/sJHUkTyjxImm0dabzPTX9VnxsWyCjtZOCQ3Q
RDGG76SsXfs/FFeBj6PD85bm3fX8iTw3vtEc1j9QV/VxcPYgOw/augL82lmyTB2c
CDnaWCFSWBIySRke/zrxANGoPl8y4RZIa9XYJLl4KDEbhgd010lGv+uFo6l7LTg5
s7+/T9T6oGjSujm8EukAIx7N/p7qQOcNN1iYB0FGFWfJIa6Jvvd0Fd6CBd9U9sVP
GqyIKtQ10HIBqpzCFTGBzASePeb/hpWKYUHtPs+z3kU9rxuq/i3xRfKXlAhYpwcB
dNQGC5SSEp1egPoY95IX58pO9gW827nlyg6s4jNDVKB/noxUO8ZXg0euzWFQWV9P
xvPFQy+ebAsoxX6do1ZDgqnzV7r4gy5JNIbFplETHYawwQ6UiFfS52JXzihrGqy7
QQq/9b9oXiCNoMSD/oWOODOZa9Udx6iWnsQTCl1p6V1nYvrQO605FmAR1Aa7JXPn
u38hJD3cJv4hCuUtR3NQNcBaSoDpHzKdhe4B8kJcsEta7iCYVuvVc/iVwQorHsHQ
fTCLSZXN3kTOWy5Y8D4mJoyN7XVaPo5zR74HvNZsjD+faWu+xHdOjIHCWz5uPCK6
7d6qPqJUhzNWehpe1WymwcmlZHnz8mM02E7aYBIyO86foSTrOpJByKk+iNVfgRaR
fg+6sNRgtpod3GodiX9x0p+thtDCfiWHyZiKnnk3aOAQ8LRTT00bGyZvsVsY5Cga
YyD65/LQ5c4vLcHzjVWeBZanZ0Kv22UPpa6+Q7WpLdpjxMzC/51xbSEmVOXHpacH
LXUrMkFqGu16lTTwA2gGFOAbbCM/VhlsUx+NxJ++emoycfxts0YPpYzj5+H538nU
b3p5rsA4yojt4b5xxsCDn0Ft7jy5de9ArEVreacdgMziuAnOL7f7liYAYOKB+Z7+
/68YMJsDBUI54GpiSxLchIlVMUXF8XrtvK1IbBj4nPILUTTMJftTxf0dSiPw0Iqb
kYDzsbyvhtj/aX/5vfdzsqc0dPPdWuBMzLJQUkQ9aHoMS19KubqKs88dP1LpvSxB
JCLwSlVcxDkBanE7c4WFnbgSkLy4j7tg16owhhDDm9MTK4mJw9f1ZHz7p0jRHORV
V61yAM1cd3SenNs0OpsIflmmZRBq5VnnHewtb1SJ7EPt3ipIj2EmwfkYDaELjdTk
pLgynnU54vUJFpJmkzJ+qLBXe3BZ4/ErcraWrtGsg/tp9XwqYlUGU1z8oqklGU4B
cph/CnPwKus8mt0woIEbk6Vi37LL4QVcSgcbkVyG+lAv5RwU4qqBXXSwM+Otux0M
lrhfTI15vmmk/BHAqmkJIAZEsMFaXu5EPSwdMBIenXQby05UO5cgoO22VvpRocmK
lYi7167F/eMjyBzi2U0P7s3OeWCupZEpz1330ctNDOD+GkJglZpdvfWUfwEp+x3S
Mv/G9iSc48mHUhjzWR+sJ4BJHBRMQ1iBghX2DtFVKDWbbTGKKJxA4FUDzMz4g3iZ
oVt2CcF+6w8GgxZHFOjPW4bXrW1a2Gfp8EbqdCIaCzAU7yMKBmfQD78EMTMM/hhg
zfHGirh2MVXwuX5oe9PSw3cLeZM/xi6ju+6SctVXnKnJA9yE8o33cmzplCrnY06i
ksvbsUpr1cHuKvRZRRfa4HLqKh9znO7u1heleX4gp1tcP4mArQAOXY4eoRYARkZM
SpLwALzyA5LxLvLTpGJExrOzwHtZkmou+22WPA89D7Cdas4zQJrB2IttLP5HJZhA
r2wu3fr4ONXr13gECsA/FS+nF8rnS60IhOqwp7SelukX2D1IcqA9z7JW13nRoI9h
CiYk3ChO/4wHaMRMY4ZNU6SYTBDsQ39MDEmG5YFwzlX6mLzMmPInzEHgH5vfVYbh
yFFP0F9N5eAOtgZ+KtAdXJVccJugZKGTXY4p6A4jyPoJGv0LocasKNABmEOE9AbP
Sd1Jvi3ANwft5W0ROjCp1AzXwME7K8eMR5ZWHmZpHr3Glu02fuN3wSaN30DoNJ+a
cPeW+l+mA81BDfZ/cXE8ANyEXTio3ndwD1UAhu/1Th5XpN4WUPtdu+LYTW/n7JdN
htaLkKIE4zqynl72bGR1lsgkbGZFIS5UMG85xa+MKKNvkUPTnMYZndRCq7BFpc/I
f0GA9pd/odw+2Ag7LvLdR8HeQnL3RUbCnvfOBO3+eFJpFDK3liSaoodVwlBeTfMF
BJ1SLSaYHBrbjHzjzl3P25vRHdSYAKsz2bG6b2UUbswzWFkQY06Z6iNXmZdRvhDY
W9N4EjQ/ASFvsDspt2bzVzAXrdmavCpvoZY4MpjbgrsSq/KGLgbU3FJk5MyvEbT9
i6tYbuCmtDjJAMYRVT05VEqICyco7clKOp/qBgTl/2AcyPKo15g5tg6+aUiNCBAX
p/+NeGaVS0A7vUKVOo6XG7OqkLDBj+kpH7TdAITCOJHC5wr9JEBXLkbNLYDAEhGy
d3K/rpZbpyh90VRfdpM4cQ1Xv8KAnxiqRBPy2ZiKklLUWC6TowyKJZ3Zc3wEBHUX
V4MuDLbtcbvf07/paEKIhZzynFEhqUBRkbC1FGhMfTpi/r3F0u0ZO5iAniW3am2o
VIyrEH/zmoljcw/tSAuWQpkjJu0cNKOXouZJU/kuTioHqkLl1jD2mZ8BXHvcqHU4
zClsCZi42rOjC8QEYuxfk722MzBwv0el1DUGyRDD7iXX5qYLxOx9diqQO7Cka/kN
lFb6bHSAkxur3RUYfxZEVx4f/Gf6D4pr4Q8+850H2cMZvBKl8lYf88lkPhbKmEHY
tY45OcnrZ/aVFMrTt4thr3RhvDg2NhqZedtBMtKovG3N3b6OVBVLR3ry1NBuB0c5
5zvhMhG4OyMxqzw2j+G37a8lsr6N6EJMhWS8PhHLlWWiNgnkrgFqeXZjym0Hx6BT
kW+zmoqCUvaSOG7qRwUYkyWtPfUpRUcQs2P75DNamdXAnkiNxNjdZTtsB1LiLOgj
dG/HnEkar2utUg/NqLDlot3mHG3z89sIXIDCRNb35iArYblf83Smm/ouk7lHjVX4
s9h856EBqBafPvSH48oS7XuLlSdwY0iX4WcLgMcMV/pKGoAOffnRjHrcksiK/7MI
XTdlUSu1LjMqd3XdVYV6+u9FYb1nX8ylUh248nX77ntcsSn/wjh+Ew37kcZ2peF4
KI510zGY8YPM4TKzeQhHsZ8S2Dp0tZ4kdbQW5wp8AIy06dzz9khmmDqWooupN0aW
XaGdUcGh29wtNbHRiQgM6mcU+KERrMmcdnyae4sO/kukoJkKUDAOz+kBfUcrZgT/
rUQE8D2pYXzLcb2qgreZN11xTgZfINKWRD3JF4wI+yXs+1PqnEwlFQ6Qfxk0JvSH
2yjq90XEgk1PMO5X3Q23eP6erhnb6abT25oVXAEmCgEeMdoHp/5LugmqrnZAemaJ
SYhbWsWCFtoeGzG/BHAqpmRse3qPSf1e92ls6xwgBuQnwnGQG6fxr5AjspeqD47w
oG6NCR+JpKWlcKGhjkTfsBnbCbLDQQQnycAS1kS1xhgufDf+Bzr2Vi1aIC6y8z+U
3o54A9NKJ8AtgkLw0curFmvoFDGhi42jdGjzs/13b2WqC0sWGltr6rOTU8nkTrqY
y95x0RBaHrQI4L6zWBF4HqRjmZ/bONKtPEqyg5I8en/x3DK4qhFjIl9FCpLwOp+k
ak6UIS0iqmwrkTHUR2ghNup64Nk+lKcSz63ZzOvJz2Iu0OboahFh9dWzenxlUERd
8pQaxCQpeIEGmLWYvQ88mpO2jA1c1kP9FcMdRevaMuUKAOW1Z1Qr9dO1lxN8mikg
boTy35Iql6nuDDk2wRgIlbw117gv/3RqkzlLGV4SOvrZwcGD4JaXE6hlV2bU1vlM
mKDezLYP6CexrTmpvN3led3cFiF/JpBkeJMDG9pMwYMyZQy6eA1mgeCFqgvL7b+q
yg5p1TilZAS/G9wChCLhHX4KFUXH77pBpu9WMEgKxWyW9bTiwcpXkAGW/ScBoeUr
9wQCKQt+7KBsNuM/lB6CDBq75JAuuykCeBYKsMxUZzn8JVECqyGJLz4l/pxD7/hT
KKpHAi9bhxCI3TBC7UdNeWoGn3vuehmXkOc0dg8wVpneIzOu5Qv5HNpBe60+RFj+
5jPmp70Hvw0bMGy5My8ggPxZdMDWSIdrgztI9+2YOLk73JV6IW/ZjInvFOoLGKbc
jnXkKhSWKemgePxiskrf+emIS2cANkpQfxbmY+IFiGxSvwIrSIJ6ODjrcErie5up
rDgm5MUuSq6bEwen/FM+wrzOyoleul3LKKRt8+F3WchVBFkmrj3a0CDvokuUnySp
70rWgwHI8ilbvJBOjMbXD6SScaMcwbn+T+mqS/lYIU32Zaq81vFzCsK+m6C9VtqK
FZa0xlO3ULKxdUAvJ5ypSe8flLIzx1xB04meLqTynPKzjY1BcwQR+qaHk9ea/Hav
WgtfDrK6lkMDAs7egyc7EtyEtL9iwMuckKHIEtwFSpEr5i6F+jgWy7dVzct74oUr
LXwXc0cQQdoMrWlxYI1S4XNJ7GPbLRLXHEiwMCiliCpzGrFmvqgoT9ZsWE3fGNGC
kl2quu75GtcI/HFj+WAh8xgOYc4aCc20OEfLQeQc7uSfBcqgBMUWBQXaEXEZhLnk
ZqOf/R2F30CjO9AGbtCxnISrZ4OaNcHuYVxiCkqvINWqtvFlCM5EhCGjrsNvGQi1
d3+oDckHNfvcGr5n1mzq6Yv2VBT5gS84s34xS++y+EWaC6+Pw5hl//vLEjuqhVhx
jSqPWCc19T5+fa3AG3DZWfA0NcdPA+8ROvru9u0QcqpKfNFJl3Z+ROvujJZGPU4B
SSOWBF1VYvbVHFVFE2ykXhjvnPGdv0hrg/zKtuYeil77N2IGxG0iqCbjko9tz7if
OIlix77wJuwqfZjCgoK51QpMVwnmmYVR256/bG4E7WfeiOJLzloZTagMGT+6T56D
mfh9C1qM4fscKIS1Q7u//QitogGZ7pP481gNNfALxPe9aTtncdGqD2lpf9F30POt
51xtOVFE8dj4AF9kWutHz5ILtFHlqsjqZ+O4vsT5k6GwhP7XC0NUUlE7DH09N/Yk
+6KGTd4A7lu4DfGnYHnrfuzFhIJT1ZmJjTyWpPjsGYR4sJdtCfwWpJnMXC4XbF6A
udiFLsy5tSLlGD7KLNoXXamK7Bih8EhhXlGv0blr7K7deAQucL54K/fsxerSvgWj
snevFNPTJx0hXHU1nB+Svq63ChqfuX/nv/HXSmcKwm8bzJsrq5pE4wBpUL9btxsC
pVBpJ7eogO/xiLsGC1+IQ64U8LUI597q+Y4stWO3ylbjGq2XGrI4Rz90vA87z/8J
2EVls6S+itnRiIwq4PZOD3hIlIqS4BLugY0YFBGwjI63tnbH8toiweUlidR7ODRq
EhUVHE5hvFyOO81ZiuiOKYIy9gaBvgf0rLRaYgviwUhPOwFKd9RtbPfOuSq8YQM6
q7yINK+MGju/cadvEfVjsfO7lCKT7tWYYPncmkM+kN0QK9mPCTnTyntUuqsqGz31
IWIbI5aZwTjRXVY0Nh3DY6HAuf1vooS+4O2mbXAYuHhmP66Br0naF86/NxTCZetY
M4l89ryg19mKonujVF8ccKT+LORyDqF6PKJv3SF1l6rJSJZI8vjT5Rvikb8ODMSo
RNjCtc1tapoDAnti7JxklORoVX6im++lyYJXdGd6qAPdlZZ1uvSZ1dnPzpPMXYfc
UfLQD0ldT90ETiSuV7r97E9wWnpPwvXulvqXOfLGWHExX7/Z/VTkVGHrvV5NXeQ+
J6G+6L/+Ywh1pUCPYKTmRsLAXZrenfOeb4Jn1cDLmZtRDB4RnfHOLScxGKauxy+U
eMs+LEKJbpB+FM9i+EpkPAZp7Hoi7M2PG+W3/Nn6gwzodE6F8ncgPnP3ll2+sTrm
jevI+uVfWLGmFo5hspeZlazNnRskC2FprGy74eV8g6XwboXlxilnv6KgbqZrZQ33
DCI8znkRPKZS3+QhOhKbJcrESkrwwACmqevDLxW8zHdcpawkruPCVykbw929bIBD
Gl8YBR3tvNKIAtsTeXK0E37o7mIDb7ZF2DoESrKqf8qRFaAskjpPukdwzfHEQJOL
FqktQsSaoLlC2w4iCiXNoHjnq/N3Wl2rMtrju5U4OpBKiMGV19t/XfBXTcHQH90H
akyfARxKKhwB4fk9FEm//GAnSo18soAQLRiVNzH9DjYUaz0eGHH3s6dNr6ZjezLj
GRmhSYrtjjpnithMC26k+eotltkFnPIUbAHHjocE8obzdwrmVB094mS+A3wLvoTL
qMpYJCSg6jB/Esr/NwzHoxBDoWAChABFAMfOzy+IR1vKtloGHs0Imlgtp1wZ5JVk
2iHpjZg4WPnKzW1thOUaAx+jF7C8k3Pm6qu7Lb394wQ8GNj71ewTGW7QAUE4h+cw
ByP1UeA9bLS2Aehf7xIL3JASDe4VVq4rhlkvuz7kL8aGg2izU/SsnLEYaMxNOby+
BmT6XGwFD9JZOC7jjgKJlWTI0lH7GB4e/+KOgx6yY7XQViACwIKSXmf6BKbXFf9C
xy2B1xf5apGR1tfJdXos24OBgl8v5p0lDwEhY1zrvkbke9vpIAgp6puH35Ok7EmU
E0hzxsIwemk6dBIKUJG0IC2YjEsczmP8R549wHNjKBJRCMIk24aEkQMw+W8Un0mW
XHN6WORf3HFa49mBHlw98OddCNtsCeAK/J52Z7C9ci+jeBSzlK/zBtnn63VsqIUA
zEb0Aa2TYvn03NBOs6bpIVvAiffAjArmvn1U7bokVnynHuzG2IpSL4mioTQ9qgQ4
LSJwCkSYauYjEczTvf3TakMlClSZIIXQYoRiunFBDpi8vwT7A94+wycb8ibbAM1E
MB1OkDuZZhTByn6vOL4+9zx19jKpAuRBKAe78UjGfjjFOScF7aLUJJBdrykBfHHF
aW7I1fZ6HvM+Ihm14059/WU5OPUzxUbFz4N3t8MEm7BlgyI62RpP8a2E2su4uXiW
3UiJ1rgdMH78ONdjUth/KTrb/f5cAiQH3QuqR7Az4bunIdy2RBChQsbzs0S41mZs
3ZY6I1UbXSVlC2/cP/ON6yGxSc8tgCWKkhbyF+1kNaC4y3gNcUtDs2Au8nnIoc5o
aHOvXZ09Tv5Ha7hA8ocrGI5GRVhqIGwkc1plX2beUeCbL4InXzCTgYy2KrsZVjyo
bHxHGpzwmdVe5Zi/REXMQ6DJNSe3o/UdsXUk5EwCJoieyEaCrnNopM42K68EU5eX
ph2OIq+/JkK5dm7FuPgQPvtNHtlnjjJbx34ZHEbqaNzmg9ypEYvSCozHdmKK1h24
fFsUtHz1jP6+orqyucb0dEhih1b/y6WL2N4RLRxIy2Td/Y6Huhf3TS/B+bvxqIjy
etIj96BBkmDWznOxz5jQ5q5KeQLxyqHbAs4/mZYBVSdPDqatLlcHB7AXtnYC2Q0F
0RfdwQ7KIkq+LV3C6hiJg8FPM3pGDXyzWHHUL6fMs2i9b11ieUbbuVEBVKrYkyZ8
LN4lL+F0/qQHY+zbDfEbutHNRXFcG1dqnh5i1fLZMuzNYzRU1MsRPRo9Nz8GZ7A3
B2yBscnavKJpXrpvlR+PRUqDWZB3TgipPWlnYFi+U5cJIaih7YkAoxc5T09B90vG
nR6ugj3XwAZfu3LSaSyw3bVD8FCqkhO4G41p5Jf15cWIJWDHTyDmt3HRSNCcXUJo
COI6OSU5v+QY9P8HOPTcCNm/wpzXt4sLCVSOdBnCYyoZcEXEdvcf7WJpvKO4IllU
ARtji9AxVAzzHF7VrkDbHtAjjl8AnjVVnG4pXt9KEtokdRnLOYCq3YK9ZD0cW6N0
JY2TrUZ3bqIZLOVuomMmEK4YQU2s3TRHwjTVmI+hmzOFX5bUBbYvWhXIyx73IVJW
egzQdKJQNZHZhNlZyObnH7ahCJNTGp7O6XZL2B6cRdQUlkXBF0+6tWOJCTkBFvo8
FbtVQV6fxJ9XVz1hpQpl35uYuhAlmtKHMZ+ZxTFT5oaI35d4jpI5ZCmCcJu8PMU5
re14S7p2SLWJZX9mSkPg8RZwhBMnlO2UahGj66kGruM8W3qMcc6EUM4k7kqvgTA5
VRkHy6VX5mM2vTObXG6qvLaHYxhFKLqslSI5rk3sLlRXT8vv562dgafBZFurhbFx
ub+DwitLU5AOKT5d219kYWdYSDub6hphfi/bIU8lFKl5+BeldXqiTLm1hkUIAOJ1
QuitKk04KOPGAVnrmnvB3YfIZobKYjI4DRzLa3HE3UsqOvejGO8XS6/e1Ozzo2kI
5acQ3lw4fYQml75qqmIRogOvPdDThQQjsQx25L7iFSHr9MZmLOswbjfCd2Xc7ncf
bVhGmORt0Hh5H/y9c8SQvWu6ZUK3arJKOZFUQ2uYy7XCdXZvO+OPMpiju7DxrQqn
rn7Q3Ott0D2usTvS0qCJeT40eczjNgHNz6pOD1IiN1LClpHOzldNRki/co9azU7b
2C1OatwcDfYQbMZauYTcnW2INjtyGtQMeEcHoT1N/bpqRenw64HWcnielapEJ7TH
FBgcY/qFP9J9oBRN17F4H7B1wR03KgEZiTkr395KW1oGUnV97XiNw/FMMRUacOXP
48Xe1Fwl229oBokU9ZwzclUuTdBuz2ruIUUxSLAG9dgcEaMA2n05NPFDF6vxr/x5
mrJ+ErN8RCt4u/JN0J3Rd0Y5SG1pVpazIjYgLzpB2aIBVbKn5KWNwGBRVKMDNkQd
GdCV65KzbiF5ZikNkNHBwRDkHdRFxjG81oeQ38sfhTOjJ/hoBZnnwHTHAIU8MrtT
G46LD+ieZ8YeN3QbofRcGTSQrTO1vYmTSJR+k/JX4cx7UVOGp56kWvWvT5S/OWGl
dqROuNza7Q1xtSfU5ctRbuqMnDeh2uliB8YYeP24/OTBjouA39BipTea/i66r7nG
ovJhQEsBZ32mhxd/Tk5nkP96heYTMl+RCIZ1lVTP7ghZnD8n0zUZCk+kFOlx9ynJ
PBo0GZtZssmNo5bUW2v1Y32AjhS8raN5HSYlvwwNixFSPFozwmLJC70XqTap0Sub
K0kUyWLMSKlDGpTqiLbKtyR4TYjNeOlfHWBqwMdwcCsr21/tBaOXvnH1x0RnnZ11
KMkyWmv9ZnVpKvD6NBys++DW/nm/dRKOB9yNYdm5bvZtGERLKaOfjAIhpcdOELsl
A4n+CYC6Owutj3Qdzm1vie1XZlpAw1k/br4PNbyJFBvXSa13PYgQRJyprROHBjah
EPWJ0e4rxKCCpJDJprWTs7ecW34DHnA/33rKV2a87a3PhFgmOudgiR32Ii3DqX1/
92MxUEL15mdtBRvSCvdK5migNGET/48dFlTsdMrLc/DwDFGWk82UKsA1YonYzK0W
jaQDKg/tY6KFYGh0O5paGen0Z6nYyBhAzF/TSHBP2UcI1KekWdrPPImj3EYNShqO
8EueV5jr6iUTJtf7ATQxwfkVwUWZ2fAMhufTf8eokCEJ5LHZ8+nNEJ7HcWCmvyip
DPKciniPjPMLzhNy6QP86PSmxBNekj6uoRRmAKczeRJO9hSKVTrzBnMeTKl54SWa
AQhJCvWH5D9MV2PPkZ6U8CAwRulE9295nJC1ZKZuM2hoqrQo4UDMcp9CL2V9EVrQ
ffUu8NkasVKLKC4H0Cwij6VdMTTYVtY9Ug7H/ewiCvTuNRCUll5/s7PqFhlOGdv1
hAnMiIiDieXdiItUAaWhpuQTO/B63pdABU7F1pHIYgYB6S/XULpLafe1QSIQ1AJc
H8K3pAAi18uAAq7ZfwCV93QNeC0niBKgoydSjbpTDXTt40cza+sPt0i+u+nUXoi5
hgbzfoqmft1qXLK7PQzKBGgLyGU6DN3DTkp5lX1qsmbRom1dx9E/WGhinfdjnXrH
xH/tsQ1uiQ2834CvAcNdANy8AZXC2u4xOlcbSpN5N41+MN49+48yW+U62SoC/P6H
XBAklwmCaYKR7xESmXgKe3pCXlVg98F5wL9cetwonBmp4jDvZ0Jj9L/rU/fohok7
iW7ZomGzMmx05pM37rDtbEyJ8B5eQAWGYPHXIdn3x1KzRHcTZ1F76j4/bCz0HwV3
dTkOlvyTmXeRIIhVzo9TJ5HSFpiOon/ki3EtgXt95MwB3mFsvVGmVKWbM4cV1tL7
8kPouiFsXW46EEamn5szA+xQTevuCYxZnbtZxKfdGVFpNwQvLR99AhAboa9upiP5
8/egQ688i/xY9RSzhwf1ziTou800VmhWdFh8FQ/Yj84UNR7i4E5N3zvilCBUU92/
O5IZsvEP+fIo1nRSlNVKn/TGCCS6G1dwG1Db7CkoLM2Whjj3ArDVA+s/+lF8epga
N3f83PD+0Ca7qvkhYhDnMLDI65b77XhNErjiQNyu7zEfgGac63peZ1PAdtKSAJWg
fzS3mQiwRbWLeYWSFWuLhZa3SagmI6LGyAv3TQtNxknO9d+2cZNrsdFcMvBUWf95
AAI4xNFxfmiwaOfaDk/npYK70mteYetDakkKbr2rDl3J5hrqc9tn55IIAIe7OFCF
E3IvT99CDkyo1OmVXRIxW/Izrv67WZkdPpv1Ic96vFyJobNftPbHXJMrCWOoKibc
KAzvu0s4Bn5ooeC+UHuw+ljVgrgLCBbJR6y+Jb1bpbKd1rwSv6nFm+cvmYsvWqiI
r/CY6SAP+DXG9Bzy7XvQ5cnymrBWCfk7L/M94pTQVRjrJMUoEXhr1bISFfymwNNf
hIrUi6HXLyVQ2qs95sxR34y6FR+ek0ObM4Gs39up7U4eJuTxWjx9cxdmI4VLe3wn
ihcYFkt46OqvaVH1oGUGt92R/HbUoiDf0MDTxu61Afc3fhFoniTO2GPGzelhIDyq
dTisww2CQngi4YF3agT7HXX1u/SRFVcmIZpGK7oGoucn9dtkHQBRu8wq97QIc9S8
G0i8WQvqkt3++uKdG84HQ1PYdVn7bLJloQT0Nh1O1qlaGEc5I9bACCPipFwNoiXV
U1aHHvOFsI6dl9KsmopQkplV9QKFIM21ECMIuIpjFd2KVXZIl8tx1g5eH83ih1H2
FFu1dNFSxpY10KdiBQ2NjtYms2S8t5ET3yBM1aFmheudTEtJ6ZZLoUEx/0VY91a+
7ZCwYX+047nGt9HKk7kYdDWQYAHqBjpmIIA3CLCWVFsa+YSZVY8YUFkHKPPXULJ2
cLapTBS2hiLh/HWL6bgxILtmgUmCVfE28H/E1tDhbFwOcstmsoMwCCezAkZQlfEz
WKIXmhdUqzaYOYjACqCuOgS5qoPUSP9PhPgSFgr/rGSYCk3tBsSddpq0WsDKEeLW
Jg7ronDZBg8buHwb3RPKgn21tA9u0URZ/by087bjVQHuj0VmkyHFHp5XKZotcVVZ
xtLldg8UKywIEcW6BuKKeTiLKZ6yXkExME5lSyDiSn0cst++YCI+2FuLQHsMH1oL
obKFzpsvDdqFHUBq/So3hpoV4GGbX4iHaYPV/5aUhS1YB5HM7pR3v8Txmno+46qi
ISHGbNBvn5nCW1Ek1tABtN/fkltiEYUH1DcQPYPEmQMJY+Kq6Mwy5FkFEJWujLAs
s/lZ+pdCDtFo9t+G1GOO5upGATgrTcUekbugZn/BcmdGUhjirrn95JS6dR/djWsf
V3j5dvKrmYRgerPyoAXIyxL88RNopiaIcNforOfZcro6fGWCCFhbA61PJDl1MAZI
U8zi8rTWOl5ycBFIPhAMeieWj4uVeHN9OqV3uRtCDuZLlAs7gs5Z80QAQlhqD8HC
ucjVpkCJgB3xmxXLBXP5nqFkkOKIAeI4Bz5fR1527mZKXvO/ZaUYy6JgvIZ8yZnl
0O7QPr4rogJDQ/6/Zhquj5PfYpTD6/bVW2AI/CSlF+i8nm+n40KSei5HXfNcTe0D
+qUeW3hiGX25M2tgyXJWX0575dq9sYt/3hcBvnqR/CCvmS0aO7GPaEye4435mwnP
c4YvSJ8y49wPldmCnYBix0J1zjFggxKdUmy7mINvhUfzYlGc/GTUBFkJVs+1aPfN
fTUa/CENoWQhpEGDvdtfNjwhLeFwzfGG8HI/prEtNWCM5a2cw13DqNFbZV7E6ZHW
nOM3j+oINSmFsmVsFfUatuMMvI/xEj3A6kghfvfmPyhHOUP8y1RvsSnirTdWx5Yv
IW7BT8PcQoVmq9ZZTHxqpManSbg7t1WpSkgvfg1bT1QJIwstGsMNw9LOqJ/y0c8O
vtr3AhzYaUUoTzdG9dyL1a511xuS7uA2Pfo5MNIwH2f8MdBZcCrwyPS5i59us8Xs
dsx1pghwWQHQBUQZb1nZVwupFkZvH/kgVaNvQwieiWmfBcsU9HoWhN/ofNRkb+7y
UPjqz/zh++XxVopVT2yRxyOD/T4minyV5Xhx5dhyeeeJznSdI0U3XR5zBsnTbYXE
P8Dg5Fw/mh49AYnsVKVFey4K6uWGaNPnVDGLw/mWENbqiJg8PySmOD9VbbDhAner
BTY4i1JePXgTcgFW4bU5YqinackKJfzm+AbX1YtYpiscVDdHZHbV7dw8gpHQbTbI
sVWLbB/qDB766zKoUFpWlsJYlNpxuMTeqkxT+AdlgDcgWcEVYGcYDxiUvHHhfZtm
Ucagcq0cEVKZwTU0fxCv9GF36NIhnCaWp5RIL0JGC4W97DcCKGbRqilCHav6K8uH
U+IpBFqTkv2KblWu6Jwl4wntJ54e8Ti+f0ISb6LVh3N0BRyP0lE0LS7s9lXNASa0
CQS1DxdrBQoleX2V2iMDSHJojwxE2jkBsvo5h8WAXDCz4YFiI6G81iL8TqFu98IO
ZE002MhA8jOjit1Uh6JMGco/m2lm5vuTjcBb9Swje/9lrAuEx6OVJ6BMa6awF5oS
QttaPhFJuVlXufmMy/y3eyInhLU3Og/q8fpkAdeWSXzY8t1j7YexBk2jU4MnZZLk
i8h6CWqAnZwn323UcBUKNzKnrIwwtcbFN/NMjGLwrLHnTuLrP61+sNMbqwpUFX53
MFoJDTL4sukBonWmuxetM0WXuAxjSNqVwuQRWpoH4hX1TpcALgpY2it1MAMD+Z8r
Jw8wsBDWpOI8QPksvt6GPBNZezeMyjQh/EGNx4kVLEpHB4W/zJRxQGX8PYTznDEb
BDBza/+dxWLrkLdIxysvULmZrRlp5v6YbneN5gBlPZYoEvsMvex7H6B/CCQsgp8c
g/UBP/6FGLVb6GjjHI3hUxir9VGVViY3vxWPWtykVxK/4k0AoIUVF62DwBQ2iTvt
RSF6PHrm4a/cxEXH02IAPA8CGxyAv2GbxLPVUn9uhwpVncTC2LBEN0zyU+zDjWS+
E7ASTRI8zeciFHp2hfnKJD5fmffyEKcaW0JOFDKtpijpjBx3cLjZwHv2LFJ4toXE
6KlO3nBJQxKMMyqm/6jK7IK6LEv5EftuVjK2YyBR1qz2eu9HrFwTqcqLiDATAqHx
/1lKgr5+WF7zxcKc8bn5CDvNOJOnqOWHsRaiThpaPUctt6GVYBE1Qjf35xOpamao
8x48nXHmml7twdRUdbweRfMLzKsYhl2WXKdwSQ8Pd3iX9a+5VDv+00kB7Q+comZK
eeMF3f/0pT7K4Jyk3ScexVtxBcDcrF4vyN56xbHIxHorqGxDZt6eap1rFMh7yNXr
QcdnzeUD2V7xcFoFyrorlp3y03/Ocg243wmphJUKmsi+ueLhDDLviXlcPkjcxRa6
m91j/Bz9a42Yk6e0tgotsZG7EFe6WYzDq28P8o7BREvtYkMnbjW9mvLgVp6ieNmU
aWg5Rpr6oBcod5AfYlIrYhORjydKJVMhSCyW7YGNNPAmBpOpnjW/BdfIiWw2kKNF
Wk3sU1hHIPLhd39YLLOAkyvE/38zrenWDZ8VUPSiCU+6h/nR+yZnis9NXeUXJxgn
ml0DFKOVn2AEmN1KrRYTFb4jomZdoTYXUTt/yb+X9y2S/ZStKPU2LL4LnaG+CwU3
oqOrZb6WZrYMSLwe2eWg+izFBJ/gSFuOI0m92efun6QQBrrMDnGnqHpO9K2dSW3W
eb+ErQ6EIo/LFV7SSzI93tlrEfhaHxCMpb7bDLXW5ghdRaOlqdK72IVjGQGOwRkD
PttFXtVBR6b1t15cAN6xArreh8NREXNPBurXYCHQTsRjnhpiiDB/0TihTJwxfhzV
GGHqlghGXyBBnOVgPA/BTmfrggvq/3H/ZfabkqPPy/dwRHOfbPugkbIjoC85pRDX
uzrZxNmTmnZ56LOkBYqCOAl6BJOqw6XLJngbtWjvZiQn0Md+pvNhhijTet1Kx70O
0rI6GeWE2wewEMKlSK0XmEhHVCeQiIYzK40iPk54QOAKxSJ9b0+DlybnCvqmnQH+
mEcVXS4CgGVmVGk642CuLum+PTv2+KE4rICv+rVc4ifjjOzyXh2OvCqxbB2t6UzX
bFDWaRpl2Y8FCxFoP2UaCWVNny43GhlgZWu9eWLYF1xOxd/xi6o4Jzg6XoLT5wif
2I0M9QhoUvwlCrPskvbApmVM1J3/cCGI/x20SdoiQl/9egdc8fWSxDz5xsqMEeWK
aCiB/9YIA/ivh+KJ4DYUdTxodcMJlS9ACOxiY4Y8g4D+YKx80XJgY7JWlmtHUrH3
9xkGiY/WcQzV/SI6IkbDmxYwh1SgEVb+7jFoKHK+iun6YmpVnU7BSEsd7lfng5AP
3to9EJuhxMZPYe8CNN4cp/ulT1l7bw1jEb6pzSMlbMwokRF2jIOQNTK5oI5jxTnj
/bFMiFlohU7gO5HL/D3trELG7HleevG32d4NxX6w5gxAA6PQVpKk2TaauC6dcoiJ
Kh8jBvnhGtPO7PGhkRL4EKe9CU9nNUL9/QOFRv2K+5ja9l4YLfKGpY1WWMtX3jba
g9dEYiiA3tyi/LPiqnrUpDvQU56T7n5ot1CeA/YK1LFeUWr23JFJJBlWxPFq34HP
stNnPvU/y2w3nklgm/qqGiXQBU+SFdk9pH0KQGq821JvF48j2HFuBBTPC0Z0yX7V
X3wVPJ2MC5UNJWVI5ZpyirGKMg5hPm0nBptm/yaHzXEN+3mrr6GkXo3aAp6UyaZM
FeAjkj+zhMmARfMl4rIFz9SetokqO6/659ohdY549Lx+2fDfaT0yh7d4+cbItf4g
myJpHonsOjAPYWlCQIv5rOcHkSvmJlVCRp3VDFSDIZAGOkUVwBUKMRit+YBfhZnC
Ilh4EcGouXIFUlpHgX/1MfuUtPRZ0snihO20WV0oaZRWsEeP3xJM9VNaINt5Aomn
oRYA6uFf5ppHhYYeXlYLpK1t6RqVxaqTfFLJIRtvYutNNWfGr0UUMWkBVmjqKjKR
NWU9z9fcz7NaPSEaViiwUgXOkcJhIP9d/qFGvgH0os8+a6xzT5vKvtA0ePFI7fJN
PfAas5gcmk2Odugx15gSaDfcb2m11hSgyAOZZHKbRTytOwVpl0BZW2YOcJmppvSk
EAeb9kU9SRJwMtfdlHV0lP6RK3rb2yZH0SeSq7tR5/n5RbB4Ymuyftn0KhU+cbJ4
o5ZSGo/XPZR/CA7HoOC4PBPEtlnQ73xIMyqVixJk3XZ8Sm8sLqvKhPmak2hdg34b
rCIT6bCPYj+T9UmJH08/7pOmth7DaAHSyybOX3MJ8wxf7XXNZis0oqygLxKx+iNr
W7nJt0S29Yqx7/Boji7VbZBe6gpA9y6tXpxvds8252Q/9j63nk5GeeAw1F5ew7yx
su/7B5waUlwAf+SGbwtiYTTqgjD/RnFL9oBhEObtGr+8DeflTlkQOYtBdvWYNuem
0T7PqzL2HKBpP1Ecv52f6Ud2gKWmMXlcvhU7fTtbiqopur5/0M9cDmj7ZP8r1AWc
m3EVx8cziHaS5fXprKKUnd0oPoFLDqSgew3pFDf38Hg5DzUub9Ybhjy6CJWvHr03
nNEgTrqCsemd4nNG4QvUuz6wFVuUGKIuBHlWgE1AmBypGj2J9FQStpSETOg2Md08
5MZnMXinE5bwBe+5PmpDJXKDDO36KRnC1CGuLN+eKseOSxh/T0PWr6zB9zAPQek/
qZxRvyhpTplpVBfzgSN7eH1FG2y6oxdaEr3mzqlOzNjpnnk8Z/Se/owazwP9Fwln
ZeJiJrSZ6Ut+ttzAz0CBwGQ2+zlhnsHWdnJO+PeICPjm6mnoHqLJSaVGEICsneDk
fTw/mV+Tf1WIO999bp/ZkDo6U9qzeXQc8CivDJxJlwmFbVDrdPsReYuGDVSPRK1h
QZIFDXgWh2ica1EhxWhjPX9PX0m1e1Kul2jZE2KJfE8wB1havGXfSvuecDKEERlc
cj/5/a6cAzFVfDkFLEIV23r2D5lu3c4bnLZNhXHMTzYId5Zn49FZ9vxVOSyPwHeE
d78tCKhUTqt9EUGfpKJgIVtFa6JqF6IgTRbatLX6rtKZo8KM8W90OZvym610PVTt
azgtOh0m4UX2NUDGAlhhaQyOvP1WpfvlFPOiSS5cDWCXFTbtVbwPwpdTe2lFn590
Q/Mo5ZHoVj3iq8AsUbFYCwr0WyIoDHYIzulm7J1X3GrSgkH5PgNWSoVI3dAScI+k
ktWvDTdAQNLZzJse5z8yieL4i0g5nwcJVpoU6p2+AVcaVJ3+u7015WSr4EEuMv3h
Hxv6fVEtDGwh/3MQb5QKhPEdUvxUnAUX4rjdEty9+npEUzF/QHQfQtu53TDY7OmD
DRdw+KnBVe1szgWdrp60FM64oqPwwMdyaEMxKe3gbXsuJnidkeh5aRva+Ebp/1EA
3z6hWWur2m2m4JGw3nO8HA2ov+9CFHrWgoYrigxJCs0GjYyFLgzkJ3WMhVC87+Nr
43neWopvjRVQW9ZFbfvaEMPLXVMSK2fTp3V6FF5bMOSm9aoMfFETIkkhfmbR97FK
HxKnyWjcRNl9+BjrgQH3pF39QiUSxVAqmCQi/KWiDk7tg2IXYJPg+Z6wFl+SLKNm
Tv7diKw0f56J6a1Ijeei3wbCF91O9+tdmfz/wre2ALrSI45oBa4LYu5+dh5wUNSU
azxpdX+/14ItcCS4+gZEKjmFZdwaR0aMoGtfeQOd/cH8Nl6mDlL00js1TQI0gxyN
D5p/Oy7p+6lZfCoSCVJ65B5Ua7oOXDgP1ocxBL82ETMrRxffiatM2yx3hFjq7+I/
05tLTmgHLq/ZBXwkYTAM1knkk+iQSHPYApMkXwCviktJ7NHk/4lth4qrQHFLD7+V
LTAZB5+iXPKU8uiwSOWYi54mneT/NetPygNBpiN6JHC2epjCid8gr2P60gcvS7uf
qyrCVFq0O6mOyCpb038VC1MDu6y9jN0luRaJ8M2z8aR9Gs0rcZaqeqpWUYeiL5py
0UZjXt8FBNUV2rrygFh8L2LGVczKZaWZZUo5BaRcgsoYw3fAJKOXYyVYYFuDx4Os
L1HHkGOb7FdLPrr2ZuzJwkqaZVF+5IARuM+K7diNN5CLeYmPzyDuxEihO4m0KAZc
8mlTtTEqRUvIxFrVbVmWk9OJ5DQ4cHkG4rmvWZakw+6WOJ7NxzFbeDLKlOr0WRIy
vdhS8ByvhlJoawjLpL/XACRqlRmw9gwiJ/cHDkzfXrTmda5WJr392LFngGh/duCK
hJwIVtG+OowZmjzItsFLpFyXfucIscIkF+dtPwEsBw+o7uN9dEF2Z+GC1xGgoqku
4onTdTwReql3ewcHT7kAdkCvbZkAm+YtgjLmzr5wfKMFYXd7ad4KKUwQdVUI5LYK
K+CTxkQz3VxUebP7mT5FvgDDDYtk37t0cbGFoaM4eUClsuRejjQ1ytHnQ47eh7VI
DikDXvmocESsbLGDuyWYKoJSqHgd+BXgqN/toUyDtkv9xaqA/z62+Qj7zdkMiiHb
wzQmWPFWbaD/4U2gdHJa2O8G4GltutOGJnvGyiRsxzX1tVhDkFO5obczsmyxI373
WE5LlkDXR2WvO8j0OV+9szja8i/e+VYTMpU11QO5GTx1Q2jCO85lDRAHu8v6F1kV
8hiV/5J8lkaHJKERPyQi7GIqCkyEBhY9nDaq1atkQw9wDWpDMj6whXY2e90i5WKM
1nkqONPBg4xs0WoNjoHRWlHnDdfpmQO9KOWAPyEN027WkSHvfX+EmIHadNQkc7nW
JLrPPIaNmPrOdhiok0iOXn/IDnNWfu/WEPBA3OopsxdpxjtEoVayXsuWX7r6tMcI
zV1nO7oW3FDtwrtvvIZYEghKHI+ul7NAcuApYrvim+ISML+ZKoagnj0pAg2r+Emi
Aex0eIIu/gigEpxxocCDaa2FhNrD5rfq7ho/WCyAWsDmN5O1crD/+o4Tj5jyqTUg
ZbXJqjLVN14s+dt99A21LUjw9JM3gkFa/DlnNKmy1XvhPCV6RpUJJYVccTo9DSyL
sGwovSwogajTRFXKq4IRkAOgS3Aj/PQQynZWTrzSX4uh1kUpxuT3odF0eLXm2zfV
rNZzmODGFPkBeBCsH6bdgcDlZ//ywcoWfK1iUwpZ9mowwGMsOigc0TYmMkHyZOUb
dzUuehFeKr0XiJQA/bUCsTIS8qIWj/auyZ71pF9BBZJmAqAM1Po4DWMEaxRwYkDl
e5MO+jFne1gebyzO4PPPbGzNtCisY9GY/XtuZeqrwdouJi36TMPBBfBaLcatxTp7
wW9mm8bC15Gz18w2hSHmh/T85LGtD+xbI/sxRiKZzBhXW6YwR5GXsvXGlZjM8lM3
MZ4enfF6FKuHFXo6Q0eFnN9ryLqoq6Lpcn9l6DiGz4XPeWuMdikQl5qR1eQnGn5I
kH0ZXlof8PqVtuphYr6jpf0MVKZ0kpHvzTGtAinVsHKWOgEAGXxXQzczdyMKhthB
CsvEbS6W2agJAkF8smCXRjL5PUf7PV6UaWutAmrkW8rNYE5n8DYt/53LBPi8j3Nn
I7Yh4TagNqA7DWvOqDBV6qc1/PRMDwEUwx2dF4wK+NNm6hfe8G3AoPvXJUwkHD4G
TSHdToVi/7cyfTsNq8YTIEkIn5SLLh0qY3f/eI5GfunRCCdlketRRC+TCVXeB+T/
wnsXBRfJHD2HpvQaaxcwiow6mgS13GaO058PCyeIlvNMvQheO7jVgnyDDQqrZrP/
yhX4EbI2OVKGlj+9enOyhOKA/G6XVC+NFOajPHREVIdxRa+bJtPegvBipi762aNJ
NPJxvTzy94m8kNgOQlsAUXt0wHfg1S+4yElLn7BIlw9Gg3bLz3UAqxkKhtVMiAQD
xP+odqd3xMAOLBn2L1mOoZTMl21Kw5DKp2jXhZ3ZZLn+06HXtj8+myYKERNgm6uk
bGjBNdV93tOyRzRDwX/gUEsm1aI7ceBdG/mWy7LugwmJhDLBSLkhCEZf8qkGc0S6
RA8HpFJHgv2YjMIvVbTs/P7TMyN6+A2Q6KRmTraqaw0NHlThc002j241KluzyIks
+MrrLgSZMuX2CiamHyhelBy+isJIzVFbcK3zfnQlg5UCbFpL+kQWxd3VkBFMVQDU
FdIdQwVw8Cx7j2MJhulIkZGtLr6aFaK5EnLZCAgGpby/i5bIvJ5jv8NShZIS6zKM
n0+tXHrIKHu2yXotrcL0iu8Tz9YxMTquXWhEBI37OnZHND3aj7FgXmGC47/GEgk+
HLt7istwoBVtxWxC3J5pJS75UG6oJgi6OHaFvHMSlPC2n/pIIjEZxq8hix7w5d9n
BopgAhIXiScHpPz4RvmGHJ3RZTJ00LPuzFoakeec0jXDWBbPBq3SsLYd7NfLeRI7
8Eqe+uWBmhjywNINSALPhoJOITIciVGaP9oyoa5QQJEjOBvKsFn8J4Ex5HdECHdW
rbQrOe6NxfKhRgpJeUiz3ZieH9NzpTmv6Ni1dbuV8woM5cEqVdBLsjlSWGjAGoEB
+I2Hi7MeW2UW5jnadFHpe8w0cs15RlCIC5l22V2U70C9admBeCGizznkAGcNQoXt
xHkyp9SCy1Kta3E6pS5QWV9iRKg6zVNDyN/IB7o5k6VJz3MQE5WP68coLilG1VoL
Y6s3nwJGqRCawluUmEo1W7KoRE8k5Hz+dVFYIXYNiOs3xlS9IlcaQzCPAc0lhp2J
XjQs+rlz3+C6l9oADt393Ovz4CRDIf38ZkOdag3oD4ki1swke791uSVsrsykdU8y
GwoW4iR3a0NWhQMLkVXPdNdtpOnOLvu1uZgkrjkiBghhjV8w6UmzV+N+nrF6CUrX
PXlNw4L06M+TbHid3dtRlDTcZTWHP7i4dfy+I2uqPpVarmVMeQ6NWQPgHeNdubv5
1LiTzJWsspnitSUKu8kig0JDTYbXDMOI1PL8PzjRrxkW74u1K2xKJLtuegKPBePI
HPwZ9DGaFJZGtddxknDwpUf/6PVj+xez8phWqgPSm4Yax/bj+SPBzZWl/KSUumIj
+gWgz2to2Xce6xxwI8DO1H2X2/f14SoxV3lQSKmAT72HAA5DnVofc2X5qUVvQC00
OczanjyMs+xUTMsvOiI0nS+jwMmDICOSThkT59ZEiT4USxrIHTlocPEj1gi+HfDF
flQOcwYXAoZRff++SGZSkavCLaaHQDmmLD/a4v3ZhjFtrI+MM/h0Sd8du77o4E4J
ZaixZAFAMJLf5/Ov+LKVb55a82vy7ZYam8U7XTmelwYYTxdXAPXYmR8SJzDzlnUU
w2cvVtpV6jEpMVqj7ft/1PpBDlAQnumV6n9D6yN1XnjbMKevK3rJR0XbgH6ZciFt
2T2jj885VsNahaJnf3PniRGR/lpxLNoYD/rBCwkgYJm6CGriwP8QQ2r68uA9EnGQ
UTow5JjxaD2SiA/riu/CAihy31DOxvwb8spFJrezAFMUwoCsLAry9HGSZIXYHGgk
3HqpKxKFLjuYh8EsgScpmI9nWHWacRS4dyQ1TBIsVjjte7FPUW7bgwtC/O7xDbzo
ATUSHHkrwmfFEZZVVIUOvwM/6Yc1DbTOKueESXycMLLpHG+o3VMwzS52OEvWAucF
5qEWGs82vbs8P80c/trnqsgTGnz+lfg+cPPJgcvCFgihnQQ11iT8tFakyPAZX+jb
NZviOXxr6bFEHOM2AkFm4UqTWrjIjTs4yIEulW7E1vAVktmy6zvlHBdmcEHXpQ87
b/Gz5KwLMQXekFgqiYcFEC6w4xngxsF+Jabkx0Dg+iz2JIKyDdoMcjKqGkjjlQ1X
a3aQDirDFcn7IaHooslzekvdNO9Hg7UVhWWiQYtytV8q77ajBO3G4ms1ckOWnjRN
HkCklccyjmZjLEtrTV/uZ4Op3O6cTQCfjB9vsrh97VUf9Fw1IcDlV+eyesBcf6V4
yv7nebdwhCfR30T8Dke6NCMfaxHEgrVo5LsRVzF4BeBPIZJpsn+dpSPS62xtoAb2
xlmH0KTh0OWOHr7ZHOuPLs35X6EKUU45EHs5QHyb2bi2+Zrsv/kGHQ/o9rh5+v6V
TopMw3JqKIlTEuyMEQo2jTMG7cAg+FxVsExhxX15/ZZOVIkevuuJtYANkkMSYmTh
GBOAlmO4nHzXUB5RyinUhPsJHwhFHYeP/CCw3YZjH7qJR6tTFKHqz56VDKks/Co3
4otSx5dw43BsByUW5bxsd3TX3Kfgh8v79lWjnlocnhcXwZdx/9rkl1gmTcvy0AL3
oEbGWccrJXg10e8dbVqc+pEESxQbHvkdeW4VLYzMLjpMQpGyakx3fCg8SZgoryfz
jyFOEkF9e2aAixoURdYFwxWXFUZnlUodRXbHCjW2132brqEv++ajoeVaMsz3Sykn
lRnTbuWJezAqC7ulXFzycuVmjiulpXygvry4P+jEM1KwZAJ+VpZjL25yVNR6Y0V2
u2OZTH0XnfboRzLFzg6ZZB8o8wOXUrziFqZAvlN3sPL2F92xldaXwdWHkr8XoJ+F
MAYaSJIUUJ81GFiz7YGMGxhkt8rNGRhc2PT3ccaviFkvNP2ULLvdSYqOQedbJDya
ikWrTOGzEpFpsdFNDRD/4b39YFyyChaoQZAUDnwuwq1TpnbI3s8Fz8NuUj3UCv7T
rXvMGgmpBHxoY7inqXA0YVvZ6XsQd9/0gd+x/B5GuuczH5JaOzOu8WawSjWvwlUP
EvV3V2ut9LGJe6yF9qPywah1ZvsCrKTONymrLFwhlQHcoA1KfU06WCef1QB0k1aw
Wc8Nyf1wfaISArZ6Ggqcni2ZgZk5G7z4MUb9+xfiICFp7XgMkJwkS4WyhnPLPCBK
tXqnUZm2LUiq87a8OtyemfHvY8UgsXw65UZAc0qewdk3G0GDaJkn1XM2bb06OQuE
mOUSNYLXcnBw2NDFwlUdK0SSnwfp+CXcFg+eRdrum1R0bOThAh0+1XDzEgi+11uR
NJrP0KNlVdAs1kuoqVoM1bkeocMMw5CXtOx4mLa4azEOKah7BQLX98RFDksq8WV3
lqgKe3KpnneLQ4aRJfCe6JRMjd/IwVCfhWw1noT9VIDEG2wD5poQZEu/6x2LA8li
bCopnN8xFcdBdNqwrSZOwqr8W4pM/OYAiW02bCFsCVOHF6Pl17niXdszYaMRd0zJ
iB2OjK286XuouLSCQ7yqytVLRBXudrUUJ6/ifKhOQY2CG3GQNpeNmtf1YubkPpmU
scm+lUHh/D9LRWZkxNtLSpFmKRgGpIRIpE6hLizCYG7fsf0lD6FMA9By3FjYvh7t
Ei2RNTmqN3ReXGqpkrUCvQOn92J7jNnBhBGUeYOywZPpmKotgnteCg1UMKauS3xV
B6zLTnp+X7vhZM1zQ/pdXrnlVGQZ+RfirnAOGZndNNGcMX/YlIdPsekuDHPLsbmz
gPx5T6LtpGb2jOjAfvKosWHcqWqo0CRgh80HlBE6dZCfTqHgZIk63UUHTvZv1CLk
p7//JiQjoAyKQEPAk3/R1X+t1qId0MBvswNe0NVlUn40tl9xnXxAib3Ip+rLM3XO
piCU6cCCcf1Njqn7oPH1rjicxhfM7RYYckiiBBuf6HsXvDoc0yfpr5muvLS1lpTD
Wnv/ixnxZ3w5SHDGYg5kgBc1Awl74PX8YNT24d0oAae+2lqXUOaYejt2xCbJ08bW
nlDwElXGI2nnUBKio+MYm8kxIOU+2sr36akpscfIdY2MBQpS0sbOaBIPsPMFvvZv
s1FHAhjFij6j93k32urwDx1UttYEAlu/LjpWoZqdAGdHdcNHtIOJ+sC6EhhyRnZc
Yr7Difqxeut1s/j7VI0w62mGskioL77MtZCo/OSI4IlpFSUyEq0R1tSR/2Ft86Mh
V0tpmSfrVEVOMk6JqTxjzM8G4fNnKCP9yymjEVmPndvH8j1iBPhn9TW+dji4ACwh
Ua+Ikgb45UvClnPqnsADWUkjmaQsnStmC/xPbabw3IePkWivk/w8GLT3iHSlB8bL
UCgQZQDNDYKQ1HGIkb6VmRqh4RaCXwgyrYlHda3gYwN7EZtrMsXfdrxIbx2jB44+
wl+WcJ6SoAfBzr8RC+x1BhA2y9tvEBXZFQs1wZTZhY4w8dvYDFUPeTH8p2fB9jGS
gpJPsrn2dmJFhkGOwen1fMntVT+z8CNCdbrrwy1kteWwRqM4Dl1PJWRSXeignVsa
8uH4C2j+DfM1TYwZpIeRVzWW+IRSQzliLCrGfBbM2a1gBJX7YDAPJpvJzl/psfmB
poSZi9pxWHHfMqW7nyqlRKdJWdboms/u83jfQM4dHSAEQGy0bRz6OdaIboL2KWXS
msE97IW2J/6aTf/g2zW14z2AKpUmCk/sSEzMBN3AP+6GRKFusuZfzMRsvnCqY+Br
pP+Vr+Dj7zQGfoVkwQAlM0cCjjJo5ZLS+gju/oj+I8ipFuNFo2xA9xUgmi0q3hAv
8adJQBve3z1S2hjTxwWBFNEBSuwt0H/rnSQzQfnVjDPZpqDHslypHi3yzYUwoPCv
O4NKMpGsAtVgOBAayT5aZt0lMOkxDj7pZD4+n922euUDteNp6ygofyCkgCe6RW8v
QUVxYHncL7m0wsV23urDrJMLl4E8F3StiJnl9GtsakQJ2TTV/+gAVsHsRhCrehmn
3u57jRUyKnMYzoMZaICe1pgLQzsKv3IQ3MG9GO0WoW/M9T0JOFU37weQupsDmOfU
XU8ksN1UAvCkF2B8+i7WlqB5goGSCpw8sj1aaHZ/C9jyw/1wJJT/zKekajiC3YQh
BoYeUWKaINfcfqoj1RiPsdFGS6mi9vZnJ031uzDGVHUao59NExC/SWigr+BpY4fv
XJFdx4sk7D9mID1V2JLNqwZbAxP1zN4OkLpxPlo9jYMD9g6PaWB86iZZrhQdOGym
/24EF7AZ3kwvhRCswTvlcbVgKUrXW6LWXIF3dLHtCuxQ6+EPShZjIUHCQh4Ru+jJ
JVLDiAUIQmQJz6X4TZHeLi/Fh0QhztwZ93FIFPGRNiYfnHtdm+tvphOZ5KOFiXZr
C0vuvUDHNc40zyp9DeGNUelwVDzKYpR/tXai2pJ6PPI5YRIm0Kvyuhq8dimK7gQ2
gLEsJtRYHfk5piB0xTSzVr2bF5FrvLajd4BFGKpU0y4Uq2u0WXCo4IdmFwylfaUe
e3+kYi/gvyuibt+2Yt/Gk4Q5m192dXFcvuOeSDC3LhPYLZUGndrBo95OdukxQm3+
TzelCb1RdEo6oE9hSsRMvNOe8Rf3vVO6oC9cb3w/BAmhp2vqbWucwtXME28jbVCZ
Z4CA13yUrt0jUoCnG28if1HNL/LcDpbN3Lm08qLM88M+G/fgFWPhyz33EuikXVIu
F5zxGLvBsp0AjLpLinLfFdsWu09q4M+cZ2/w5l2E3wGD/n0ilMiur5l+qzYxaZIS
+iceKtGELdX+PyimnnjwAbG/B4HQImBmZnJckxQURxOwKwlDJ/f6rVwKeyuT9JZv
1oRH3vqw5Y1K8eASXEP+rXI3s77Wgvd4KVw9M+EN5QlZONR7vLKvLCUWfKlK3ee6
8L8TKGrbqa6O1zkxjb4FPoFy1/1CPAX5UThi6x0mNH2mkCFatfj3ceafKwEkXJ32
uYI6XNFbjXtfdw1TxIBpwFZqTUJioEDFC/QZ14Gexai2YeSABGK+BiQzCGcSuB83
gXbS7+e3la1BOlGNcRyOwvRo9/0L0eK2SkyCbz1NAC0soEGdeFyn48Vsefdna5pM
L7KggN9ebJ8JscmiG5E4eVWlITlqR7w2WbZrgUz87SGeL+Tbi/UoLhetJh7d2iya
KMrrA1I3XTAXIJj/C4AMG5tUeO4lOEQp5w8aZU8LADyQLbEcCW4nRrjvWpSiOXtr
CAhL0HGNQI8UlHZy/jSTL4wr6jRCOizwUXmIkSO25DaVtt/m0mmejOH6SSuIMO7D
kES6Z/v9YQ0PMMBD+qBFSWm8iojtS3oNSdHjLjRkcNcoQl5PYubxd0JPdgqDZQEh
8LqaqBvDkZCil8cmg7UxgVpS/ylyBXONCd+cFGEcrwTBeVpl5W5btJEU75+Qo/cz
0/9YD1UBJrolGooO4Gy5B755gRti/P8hCg0piLB1W6KXSIqNv5jciOXXcYsqU8gR
Eborg6tsJUnRdDg53WVq2R66JqzqEh71r7gspnJaTk1muhO8n/k789G2OL+M7Dph
1FnkCYKpiYk/oBXZsyzZ5oN9FosNGRPSV09v03lsF5Fl6SLVebJK6x1CxrChxC8A
y4SyKceKUbgfVWklJtCe502ZTA57ers29F+6oQNyqT1f7m6wvm7zlIlDc8YecqoW
ymmiV1DjP9O4yjeTqG3zyT9bMkkawT7exXQtYkLqqTC7gj0gwn0LnovBKaTFD6tx
rHWbtrnWaqdGS84wChn+NwFNwevZCMS5cMCKZ+V2COvLzzbE1H9LE8NYsQwZ9eSq
9+1MV9nOcOqn+8+9Ptbarkz4hYvXdk38B6syoLDVTrNq92DYwCiG4DLZRHRypiM+
5d9ZXbEehyYu9Os5xvyk62jpOT+kY9NQsJyX2ocmFiFb51d1iJVFxSZll1LaYOIc
uTMtXuz1C8UkokEoSBEuHW40LF/9fRMnY/aZvwFOxpz8xGthY51ohv+Nz7RffJje
b2fVsIV5tp1Wwo4I9WdM8ZqpuBUHNMcltvG0cExwWnl0V1fUDAzoq2GkhAV4HVhW
jo3BRqKKp0l+h4tW9cp1HlPVKeOc9amAy3W8Y4XExliAJjlWLkNKJsQ+BcH6VUR6
Zfgdx/vnd8pHFfzLKOalN1JxgW+GXvEkkc8mO+evOBnDm4xQ0j19j7xnEIc8zCYd
huV//x3rnOYPHulI73gY4Osgkwy9tSgkxfsI0EmHfCOtV/1efv9N7Yg7NDBAmtPQ
vPcGXdUP1RiD9wRgDj7vAQUOybbsxtmeK/2Iz1Qf6wvARwscOEV/be/7FENMk7Oo
LWPpPysWShrLO6WgVkrF5YpWDH6oWMir2m7PTpuJFphdpUrnT5AC3kimcj+9I5cP
V5WNK3HYO7ZAB/RhegzKjLApUhK+f06ArSAz0OMeptHAMINNCNBfjLvpjD0bBdXx
hnIgPE84NG3snBPp2JKkyJmoMNunDaOihNJeD6cb9oFGXRPo8OctheSAA2P7oaod
NDdjr+iS1kvdzpulbE/0sUy65+M7JWViahRHJdzDj7aLLWM1MdRzcgdazLVkK0w0
G7wstEA78SI99lE789xTA3oR07diH26gxk40fzLxt68E7ZouHjAwL2xcko016Il/
MXHpeqRdIqgNyEZEZrbI8mK403SUcjnYtQULBD+mPJMgxsMSAr1Ww+cvWJt4UG74
3p8OVHiSVVUV8vnrOsmr/tzbfpe6zdj7WQuBvsxcLTljQOleu080IitTdZvyO1Bf
HGlopaDCtGVtYNaZ8CwREjjhiyl34vletO1Q8h3ncsRGpRVLPIrHk4AanWEjNn9I
l7ok2E9FRvGyFKz7a5vCuZXsgpM12A0izn6YJZgvP4HnUe2oBWZe2iuVHSV5NdBf
Z2bMqsv47HUjLu6hb/70BawhmFsYXAqgO6d+3u8VepBMSO1Ws1KqxzFyHCqYgyiu
TFSqeB9eFlVJYiE0utE466hBQATspSzZcD8X1dlOiMzOnvigd44vEeeQzUU7X3ZM
/Pnb2TZ0B95X8JGdBQ8I1N+9AoRF6FvuX12kX2Hda1jKD74a4dplUHIc16UnOejl
kKnoxmBEs+69V0vF+oNCZatW+IyUzi6qCqWyLUvSOnXpBeHB63jkOwY3SZiuriVJ
Q9BHWnfIWRVCzFc4682wibVkFl7QD3S6MUVYvBWHsTVfAl5P7Gbe0qE3fpV9tJtQ
j1B/dw29bs9Ofxpj1K2q6H7KgKybzg5P7+XPukTcedIk/Zehzytj9ZZmT2a4btxv
+Z4L4J+zUhSzP0XUxpaDmS9dDYtJRnkQZb9Cg+YPqrgi9EKe9tNHk2YEyZHBpxrf
XJSZOyplFpIaTDA+SGYqfhtFTIFTaDlFt3Q/mMmU7/cedCxhHDk+HzbTipsApkLw
24GeVcv3E4Av+Awvnb8lq9K0L30LDKfuSA+XJ0TM/JmY2Aq12SHN35rNmugoVXZ0
E+qHkSNiZQMrKmcJl/PdnmwomdsjKQlU4D17a3UaMExXB+kNFHQvJKiuyVxYIyvP
V3St1ShqEDRp9/YkkJ2SsYvZ120dRDbGZc1bgFRi513wH2m29PJpn0d+tAoOvYhI
nAydcmMK9Y7N5wEzu1JPKdxHHjSNnHi8Yr2a04r5jkP9Ek5X3q0XL7OpCSbtowbc
HW2aW/dBlDsQ0B200UHh9JJNMoNZAu2K/nCBCKp/urqh8vLIqy5IsM50gMaVarOS
HaSr+aPpGtm920A9A7e3UBtCwIf2gOAOtOt8MCJ7abBi3P5065VrIsPutLI44DfS
cSBWwLdfJjJn+biJgbxkXMVL8C9KfDjFzv9XV3L+jjRrnka3r6bemBT9Zf02ao95
LqQhSxn2cl8Jeyrd8eXpF4A8Xu5THasfeuceQGd2Or/OMFCbjjMScnkxyhN3JBW9
SXqeeKvD+uPwNa3mVDnxm5kLS04F86b0maUhq40nIJTGBstuVws9Lwqb0jIvjjZ2
wvtzT7nJBoySQ6haxnA0zXFR8i4j6YI2W8SMQMvf0L2aiwlvqw8UZCr/zE8CiV2S
VUB3E+Y6ilYkVALbQsMEA4nSctRdfHO7xwSx+GF5LSYsw62u1M3w98pmwYsvn6sf
hO0+LldMnSAOyAxfNXKmSSF2vDo++AcjP5HU+y5x15x14c0Lu/nGZCe35DctA6XK
Sspats6ANlepRckYoPS++AKjS+xMFSbrW9uD2BwICHcxO9FG0wdfI8VO3BaISmDe
ql6nvbFtX5l5anPIGglpXckdk0y+AcrrgkmFvZTfXuEKo89X8PNh54YOg1nBX/N4
EfSgaB++jtVDzEQc91l3pbOe7Y8ubO8s134W0DdG8gHWi8HcFiNRP6X68I5qWO9y
26PuYY8M+v5BkMRk4U9vhx0CcLMTNtt9xeKhEHsMHFhHqkXCFXqedxovcqWbfGJY
8cR0oanl+MdRImY7lJpM++JCERgWIQujBBP8O0CUEPZhRpBn1BwpUk6LjC/Alp23
ZJfFFwnJ+l54Lz6ZHphgrEPeNWWJ/g4IY2PQxxnHMNjpSuDYTDh42gBG6HVfH7at
rS0QHgsO8TfmP8tUQISlKcxgRt31o57SC+ojG7maUekCZbtpOXKBHKv71Y42qt+W
wE/eljGH0FwRShznHMx8l/F70RvuOIp+PWiHhmL/Cl5vxUE/FiqeA8iCgRVU550T
Vr2gsseqGn3bEO/WEVtz5pEj2+kLoHmx1x8TdcD/FYuz0EzIJzJJUhuwmI0BD2H8
hB0qJ2qeLzzafwUHG/yOM1wbnERKDedsT26c8msrXVuIJNaIwLiHgK4hdzIMk2Fk
SCVbRknr5kqln3fea5c05PY/D59RB0ZbmCNhiJUy8saj66l0qgSbCyDlvx6vJrXF
pb4is+Zh1eMwDQDP2hqj6Rtjh1Y9k5pKGihDtg9ulOf23bp7ofRFZAsZksUqtk1D
QKT7cqJf135Pbo6b6CjAryIHZgJEQDweGzLObh4o5znIjbm/FYoVtWlSvTXGeMav
knWlRxAK5Ijabtyx+DnDg/NkC+a/TMqhsk8SoIfEZ10ut3QaMjVztHJHt3epHEEw
pg9Spd68VGsWACyfLhdXiv90VeA/ZmYCUlRhHgNltVOEJGO6BmPHRJhYvR17J95U
dLPgVpGhEkikiC9DxsX+t+wsMbcNHX7cu1Jm405qe4VLmGAU4UQpzXtoocbbMz1d
jzJ3wTY/EepXqOR0CaZAjw5VsgpTmG9xkImCyxVa7Dr55dZSS8FMwPYDKj6eODx8
CsM6j1juHFCyzzkjsu6c6I/javvsZ/oHzN36RVxbWuf2Q7gbNw73FZImKpXVkgGz
CSU9j/du1VU09A4z2QQmocP/Kaelm0uWnbECT4mHZuSMhEOLHmj+hAai2zHskNd0
/Hv7SOLxt+R2UA4qTReU/D2xgz4WMKL+WBRCmwSVCI6BBjTPFeVUILu/nrjVDz4Z
o9PN+DslIcFyecXe81QzDW+oD7yvpSBVQHpogHgkUlEEtdv2uSDo/2mzT9H6dsIN
6kybM9FUomi1/wpya+loEqveLLzBWdbKk78idXFa1x87qH3FX5hDCohWLptNB71D
iPMjbvyTZXeJU6fa8OIPHrhehPSqk0YcqP7iYcwLD1B+n6LUS3zWLwftm3k9gXLo
ReqmhFV8TF775EAHI2F2wuat0aoY0oABqdpHpZBT4qAQZSznEIu6Irnb7mg6CyoS
k8dpliNkEJW6Hgq+MD1sculJT5hgBokEfRjqRl53QMTTPUyOGSprqKqC7WHN2LhL
MVL2GOQpvsVFhPf4Lwg/CQItsKMffpgTGEBymlyjxLtwxWCfuCtPMRHRM6ZoPezY
Hx+LVkGWJ/LCuciyBfXuAfCuv3hGm8aCWS1nZ7/rASLxgS5Ixc8YX/oF6R/UODaT
v1VrO3jCTCSaHNPzGHua1jC2XG/ASzJTApn7mBdic4b7HSZgRZZDVEoOxIJSEkWC
Q/PJMlBWoOBjBL73RZ0tXAH1pVX3y59oQnJgtq5e7i3NPDgcwuBX2SMjTNSpK8mH
hnXpYNM5RQlFgt70zY4PF2vl0oNRflCdrbcvy4f9Fjy3HPxOazat8dPa2p/IWzs3
sGlsP1Xd4+z44S4QaxNBlVtYPcKO0kum1w1Yk4cBJ9YWyBqxqhYx9Xr9HwlSbMcC
lqJ/e5uHtP2hPPyDXzhTeu9/sprusUJ2EFUc9VKjPnT84wEoLOaVoB4Ymmazu+jx
DGCwLUDbzgL22JSRVk8jYz33182JLjOv6Ohm7yONVEi5rJli4JOYz95zarcI8xxB
xTBZKC3UstSl6ybuQ2DEXM8JSR0Hr0MI2q6nc4+IOOue8Wm9O5oy4xYnCvf4nd4o
ZLtvs5q3tfMbygJHPzeusmVx2P6K8o9yfg6VD+Bzpv6xQczhu/sksPJQYI6HXVWq
Zk54WjJMoaZZoexpErjMQDbnm8c+bkR+6mlT994k8F3AuG8HOFFt9+ZMki/0+qiD
IR37ZWc5oz2flOKu+CXR0AmJQ9H6iO+HSni8JHaF3xjDpMg37zLO5RMaLXd5OdYR
+BOHR5ORexK+hTrQNHSVN281LXcN9ioRl4bvI2YlaILH+Atv/jzUR7KYInLHMgPo
IVmLn8wvT48pwSgQGQyfCXwC8MExSbrm+X35aV+r4uVOIiu+Y1+OH9DKEq/XAGE8
i/rwE6wVo9e0FDJlUAJL8LVPa2bwjXoEiEdZAxp4FomLGGwKCeYiwwQONEh60lMP
sqsN8TWoojQlyEclul3xZnXMRcZFKS7fmsqBEdSpsYEVAdLWtTmcEJF9WhrJ8Uqs
bNGWnj/kX8dvwc5k/HxGjY545232sQB286f/YGXWwx0LKzI8uf5YD27H7W7/UfUu
b0/3adTbcWvbU7qiCfH2fdTrZ/NI7tWZ03HPLDxFKXjR6eE/z2tf6m886N+EkyoU
IY93aXdwUSyR8gAW9cvHrH37MhlvhQIToKbPSUMPo/VxQQBx0/xa5dJpDg9Wnh1L
He195QGTKRIz5xUR0El7cvfCTAwfgBq66wTo0uoWGs6A2eAPjFRsZmOkr0e2egxl
zQetYU4Q5UHRsEkzEtOCD3p4UqTAaJgLiWvyezjtN6A1lwO4H0Xi/mJH+lbQF8to
Cxf1Iaqf8301cpC9A0IJhrr392h3QzgZ+hNdKbRSkvSalJHQRBqn3rlpYraVPy0X
dT4XWPKZoaXPb64lQfrpLi6Aji0HwyN7HA8J3oK3EpVGwhEFlvMHaH/rqCqAA3zo
TJU5FQtUtTporaV2N5btfRBM30ii5YgAqoFRFOrrDUUv0E22vniZfMcZvBr4Hodo
juU7zThkJGyM/e1Uh2y8KiDePo9f71eAqnIIlyRkny7LFZyrndVpTLCH6KEXGwTB
Kex1WfJu772nPBEAFwj9VHm/4tn/DBQuy85NRNm9VALd5UXrWrgZCi7z5rG6anue
u554vivy2O7mvb6W5irg7L4ehm3ZXo/qXnr7Ce/1dVhpzn8WgVm9QVC11PLKJnRb
OR0O/Vb5iBug8/GX+IkuNByC7CTl/gp8IS1oXk7cAQuTfN+FCAR9+hhk8+wt5NjF
FM3soauynxA7Mbqob9sFJv2UJomVh+rcT8Yyw6vDkJ4qLEsVvrZJnbXs1QQ6DtJT
z+05Xo79g4sAwSo0v4HUNcS1KLA85wF2nvW7xmWWWu8RBCMdfFjFHvwtZp4mOjRf
MRPU0vTqAK7gleNprJTSaQutNPiLdQ+JALVTSXolLa3FDZckGlKHBKDLJjPs9+wa
4W4z49Tw7aBwwBMSysRk693byM/smbnTS/ihWIJhOY+83MqJh0+ySmhPr+4nuNkS
zUjz/lM3WhlCBWVzs3CWzIrFmskUS9Rf0BsxQFq15MJax+wDOFA0GclM2TiNsIcq
OUndPz4c2tJjxvrOr22ZT9QoyRWWK/IiH1oi99i05g3T6OkqwKZa4Ovuskl5B04M
tfBpMcFMOv3uZmFMi6W3TLDN2gbbbWIUM83rAuw6xPa5RAZTC2emA9eHFpvZ5wdS
I70up9baNsR50u+Ezioljcm5HE0AI3Mk6qetBeYB9ypY5JwbnarNofAomejQwXMZ
efC+3znNJAledDjtA70+XWHcVIgePo34DUwRmrC4R/l3jGi2hyCQ+TtGARnu6oOn
nom1DsIhiVmh2rWTmWiNYeXAiIvlYKVENGnUAj0dSaaJj76drJaWiq35yUWmRd8L
+bHuf4lYOSBO0sm1lZnM2PaTdiEkH/8hYP4MJw2xnuWs3/oX+Sl2EQ125HtRP3mh
ZExuNcS9CrTRk2J2tmdHhAyq7zgwq7UG6kNw6zcdObA+GX6DeKYUwcEECQvwPEri
BZlfmEJg6q11MdixUDJ2rJAd74BtYlC6aptLYNjqLOZMm+/tBlPBQodx0+4kMGEJ
aq5nt/fr1+7yg4z0CAqcOYzPBirHz7XJR1XAad1r43pcVI1EzB1Zg/ozcrc6r8yy
quj25S2ThZncPT+nMdPdeN3Mm+7ISnTOStqoGSZKQfk8V2k15XBPVT+koibUbIdd
ZJxS9BBbBzMuh+zc4GynMEmvIskC4rv3IlSHdyeQsx39ydbKsTaz6QyfINj0AlHY
Z3bFl95elWL/6R8/uCyJYf85bA40tgPK8hIXreQXTAw1HtDAaflVi1IMkosdtOlU
2hMMYJqH6Nz9UW2zbjhbKISSuRvrINbhizyaRjdrQLVCh5kCNbraGmyh4s1ZruO+
Cc1FHkReJ4y7UBDrNfdhhDU8NXL5EiLYNRWls/n+MaGMPvtK42pX4G7QKm6TKk27
drC7GIc+furMYRr/z65BtFMuUEjGLquaT7UopJ6heP2ksWzas4UwJkrLhvyVtHfF
7dW1xV9qGSkqqfg0piEx8wX2JSb+LswCpECL1C6F2CLwGCiaTYJfKBsl61p2uY5J
W8oQPsF5XVPjJ+gAf8vR9Dh+aTUiWJiiYd6AY3k9B3Jbxi4SlNX39F9dZOHg5yXC
IXMV1pYwG7bO5fumesl30speSNBVx1umYBsNeSDnrvGUCidNIuKCbShx9cIt1+8a
mGCK2FDb7pmJ94aUq5ZyrfrvxhPgmyTPy/8YYTYxNEUX4Gou17hXa20u7xeePMtU
jGy9zNqQrYfXeKoch8E9fPjMoASdnVsoz39zmpfSMEAZqbaWtjdLa7QZH3Ft5GqE
EE9roC6HBjO7K508URxwF0qDG8xjMmSAUzZ4m7NaekZ0Avo2K0qvnT1ktov9epYH
d8lnN0l8VQ3Bzf7iMYZRHg/HHCmCKn5qcC0yD+xp4/e39bpA8bnQLLNYggIHYYwp
tshok5VwOjnFzw+FeHLkUJP5nxAtvN6ic2FCbhc3mZfPkIcM/OsMG4Il2UO5dVy1
viwYuW3aYyokbh6nHroNVCvLkIR2kvx5SSe2oiQDXIcurqHnxCbdF16JkjIZz3EA
ykQlupIz81Io1JQkf1+eQGYiXoNR4Z4y7do4t1dR8JObeKhnpPdIXfsQBAnpA5E1
bsD5funbPsoBYv49g+rutk0bejCnlo6DeID5lalUIAIsy4xox5yE+IgA8V6WMaDH
rIfhd/aAzP/hqOO599Oc0z/8yWhM+77v4Dlm3BfHVR5qDwKiX47IfYZm6vb68X3u
NYUg89SZgu4F15AwQUk8yQ9jthieECoXuO/AdFleLq350XxWhHj3KiT8vCfUjiVu
RbRzNlszxtdM4C+qx+MRRiz6oaAc4bch+cfgnAKQACp4doaAMYGlTk5ZLG31Jjsf
oAZzVQZrq6eokNc7DhMo4iZzZvRafEjUdcWoKrgFg2c6fl40ZQExm6+HPxV6Jy2K
g7qbweOZYvIhZWyor+l5wZK0VBW8p3D8zejbQAt+LrS2QPNk8/gBNTaaIv+lGWC5
Ne4gNf/NAuN3KM5NtNQKx1oux0yCyodZWq6i3MJ+LJsW+lOa0IcIat6N1AmsZXpP
MyRkBCDpLRiZyPHDPRhx2A1FLqhZJYVkwY1Sqt/GnBAZhTGc94DrdD0nVxGI/cCw
P1w6T5xH44RLHzQIQ6NE6xSiEVNPFrWrZawj2t5SyNi2Qi5sW3KgaPABbLMMDAKJ
66WUfq89Fk4HEl8qQI5EE5l/zEcXkezszIrDsreYJX3F/UQO8QZpZxKwkwlM+omd
WeUN8UWBFZTAFbWj+hw6t88AZGklK2tpUivGmrqAtilC7miS+q8ac4Fe8seMziRO
eJdmaMCRlFQy2Ag97cpJp69Eq1WiA5PBr50RZM2sbvWMqKVZEizbVE4+ll4TQTHL
5hPfJow9AASDxLStNJ2dJnqBpwq+/BqnbXteyse+HEpUxFOtg+QCq8tvmGLxkAbJ
hT/gS963RnX7LCrVokimu/C2/CMBFVaDvh6kecCh3fwZyDf39VyFGp/enKl4NJSP
3a3VszEvBpujELMDnpFORdw0KuF9EzFGKem8jbDgZhiYHd6XBd2ziEWCYwKFHATf
5JtlQJsvPRx92KoilAWc+gMr3PI//dxcU1bjZCaquv9KH3FnGddvOwSA8Vlp1tDQ
PwC61nETE5A5qBAY/WZ+BrsfBAcRLngMHUx4q/4pmrxloOmHPFWdwq+Bazd87Ho5
YvpxK2+8Zgl5xmyhmiYChD/4y6XXgOClaLHWh965r4mcoQEUBHaOYMcES9cjWKRW
elrxtkktR8dp1oATrGh+JeC0wbG5pvidxhEJOTNa0YGYsIPikokladwZ5gsv8F/d
Mn/v+b978xHaBfynUDc11ihLfQJdmG/BEZWc/cswYJ3puWnU2qSfXpnCdecYR+3w
0gHAfQMBFucs8GiKEVCE+0aT1nvRv3bzWdTxZgQb2E1oSnZVkcxvbn032xtrRxSg
R6W6c1/4QpxDr6gcYdi39kXzSzGQ+xc4rfn++rzwSAHdamSP/xuJFNU2qG8hUjui
GKirI5blVy6TZf60eCo9n2AqB9WaNuzIG5PdJCuSjdeh6C9Fwr9crymvZwOjfAEY
cSo8xp+GKPgABh2JrYNiMYpQnnk8ToG+LnDdrN57pwNTV5S7FR7bsA8X5RSIzaoP
VYzTKTcVBSC2NVwdq1gIfXDBjyFpwek/gknOkQwdykSVoCGFDm7A7RE51oyeQLRU
W9y6osg/e6IQeJxJBcOn7BAIZXC6/MYFFmbpWZ2SKYmDLfO9NBDN/b6y/WbI1I+n
9hcA3okyc8iAgpKqNur1DtbxL+PTK1oWJt3BbC6LgoWQZpG49Mt0GaMaW+bmj5NJ
F2h+aTApPp19n2WFIMGP1C7eZf06ypue+fqNYIj7O0Dk4A8ir4pVVvfWdV7h+gW+
zVpeqrF32kvoawzM9t93aRygvF5ia86Un1YRe72E4RUlMTGbWyD2KeKtiMMjE7tI
z0jcu1gNa1l7xr5Sn9EXvF1Da4ILUlv1pwm8ZOhGRxirUvBIDClfYitLhqO21Q4v
RLEpm/YxDhduPsWHorM9DzcgUkovhObE3JVqQohri1gjU7c8RevZEsecnNA1N/SC
DdFCMZ3XaiUaOojDBkiC5UioFU+mzIaf20pYi28UfL4PR68X7deWvAjcgnoLT8Ef
L+8ObnmcPOD44DL/r/rPyr1TQ9f0ePsxcvGgfebIIRLPH1n1I8ekTpBgWwwsFreI
INFC+DZ29Db8Nu66TX70jCTt1ggevBwL1XfWuVdN1YE2DlKY0MGfFa8FCA2Wy1HL
uaG0nmlxDMPEAse97hjBnOURVxBEbrNkEddOq63zKTOEasGXG79/EfR/GYaq4vRk
2YGM6v7LHVKZq3BK6TokyTb5tNMv9P7iFTDB7DtUxTSo46Y2xxTYFJbwhFi8OFFC
hM0XXwww/r6bevdWx+U0g1LCt3ZIdla7kBGOUIGNTynDVwXehhJTEkIHqNNNyJdi
7l76ukYZbNlTQ+qJw0Oj983c7eMlQ60mnfV6wUO8WYj1Winl/xgW8aQDKDzGkKKl
5svt22I0T9wITNBg5nyX2ViNaVV2mcyEMefux09bC6sxBMPqKSjVked0o4CUu61Y
k/YcWqBPcxXD8wwUUhjn9ikgTGEO5+nMCe2yKRpWenBvLhGJkdT9cxeTiNVhazOf
N9FYQtqeHJmaz6/2xZMEJUDCCXMUIfXr3o4i2hQzxDLustzyojf4DYN+BUg8l/Qp
RWWvwjjSj9nSW1x/+RAELq9A7930XpYC1GqNOH80CjJW6JaHyGfnXj86EUSlgxWV
fmJIG6YTUjpAnjqxOuNnAmB67fllQ2guB/cZurmK6oGXHOWuemuGUSddKzBbjBOF
rGwOxPE9+KX/OmLXbDN0S2ByateyWtCaCKGqNAYHHdhmyLULL6kKNWW1wdkNLrpM
XlJU7zAphNmvqAOM8UInjjJAOweLOecj3/uLUt8vWLfBpoa6BZ6Bk+CpgX/bbo9D
+uW0DN4omGWmgilRKFUgV0pr9CssQzbNXJhZhp917IaXuy6jiN9RbkbBDcFR6KTK
/EqkNdjl3+2dYZiTxXhru4/IWFjk4S886UmxzKQ0cyyBRhH+rcibaHEpTFr5nDiI
aoq9vwanq8+UEmdRn6ckFv50HmpIfbfUi1emynnieH7/Ki7XMMe7C19MzNjPGeKy
RNJm5WE2CbQJkwg70U8Y5zK3v3BIklK8n1duvxoWAi+wWVIW+wrxKZa5GajwXLtJ
KyRDWJAl4z1OO4N1tZk6H15Z8f3NZt2H8QIbQHUQSg628FTMP7EEVsXmZUd4hfX0
tdOvDX53o+GvFokzox4cQNUaPWmMADbTlofz9J55eHEMUXJluqdzKaIyiq0/Q1oJ
PBhCKlnZICVgdqTq/U5mFhfHsXmZe5NOQFrjoXBlyCPSZx66HlPbJw0sIjjXBMnX
pkXoDG0XrrySoC/ST0eDvZCWZfayWX3PlthHS4v+4zw3m8yJhvbAxqdhhjG7gYBv
xcmi9ybhq+u0IwEn2b3vZn4h8tjIId05eE+heFTz+MOrX2A07d+sigyCUsya9t1R
gIk2FPozYffO2oqH3kuXGq78+Jc5mITyxblr4j2lzbER71ByYjhSJco5H5SDy0ol
3XTHS5ULLoKxZ5CV11oaQP6MioPNfRv/KXGcCGVXd35m0rISApXTbI+1RIjpwXt9
+3e5NFo6n7Ch7qWtcL514ymiYO6g3TSgW5S14onXt1d/Pcnq5lgbzz91T25vKYbz
TLY7vlbgEKawnYZZKUVVRa65BP3V+hMMdAGi2Vi82R730dXqQhA9EF6HwD6WWxhE
dlqiNJ0Lgy+6iMNOxsuByQG2bJ+XqQJSywCfjAdIHcjqIHlhwKm1w7sszF2P6V9p
ku/oF0jHVERytIDaq6vYVIITCSXO32sxFj90Bn6sgL9PJMkzJUzYmycH9c8iqVGC
lTbrGrV4sf78m4yBv28YA/zQWNamLamWXG68d1/M7BJ+sYszjrMxRCbTSsP9Rhyl
ZNslHISw1ySs6TlIkbv0bRr+R7KoxWN4Vj+vaiU/Bjd01rahSIBRkh9fAbTKdps/
emduD/L1O5m0gZysCAU+avV3TAnMUt0yXNtLfOydUZpZfi2zQr2TBjz/Jv0sat2L
Pb4V+3SobBQeRge9eEitMfQgRHSIk9f0itO1uRipE9jyB156N7YOlFExIHa1vXTs
W3NOPkPzPhqbeSTruPzF1mjT5RM7cEdRcKl0M28UGWu4qbQZxTODOJ4NOXtGhM1L
sJizxLVnnpaenYgXwzSvBDm9h/4ed/7vsd03O+AcGHdMHY5j1GIgMmk2vYvZr6l/
hcqZUTW0v6sgecPc3igRCf4UncbTV3izWWTdJzttiKqpyTIUMZN2Fpj375vCM0SN
e4CX2+oOt8D2vnB5KGro9GkUJ6qOgJJzol0akK20e/9PXyBJxZp1n6XeNLxDHdDd
nxsWWmvA7EXBefXLxOQUnQg0fUVcSzUkH2iZLAwzuRuv9ILOPExxwlkcmnSIHStT
3YFpns+b9mP0eqg7gF/6Z58+73RcIZelw5PjEIFsRwx1p4Zj1O5GVuOry6GeE18a
9AeC+VIxYLmZNjtbzzP32czEym4hKx42xvxmwRpTvc+CZ2guvG9ofsfaDDya96/m
a7rgCSIa+aJQjaWfQ4fLcjRvRcFDZ2ChzAsxsgmFIUQQLy1KqKWS3jsQi/sU1U7A
Fed0PDF/c7zrKxxblg1nM/lnTVpVLrRy1Iq8vRTr/mAzz62+AAeX2iNetHA5NmNS
79A9A0oI9eU+g8mOC3/VF7uoi4a2a8JbnBc6qoWIALBT0kc4xLGBoHXBgTiL+Ge4
9C3dwDg7Iy5hbIu5Ihl+uxRDtPzTqI9hGdFJh8GSCfL521X6j8MornBQvVULsCEu
zePWnYuWdoLyHPG+SgPr9b55M1ErffnJEvrluSEmk+wO9nLM5FK+i4r077quDmdh
jEkkCd+n82PCSeeyerjFjsm6ZBQDl/0q2MiRTwgSizIkIfeO3WzmLNgLSnEsYomQ
kkcdVgcDC8SKLJiD4sJj7MPlT0TyehlJBoAL8eXmF/dG1bkx4wztPpRpXzisRjIZ
Qejl8UyBwtILt8OhkmU9KmiqF/V1vOYbaByggvtbSEU+OFQxh8h/fFMNT2vdL5XW
lE/wKVrsyc8TeBD0nTh/4XlNZ5bI5gbaROFy/szsUZll/TDPE5rpnA7PhX8UnQJG
y+8rFBaoE5c71JBsi15WZ5ez4f01d+lkMUvGAcH2jrZQ8OdxLqMbrGNgI1EHPY6A
Jg9eb2Ea3LsuIJjHrxdTjZ2Dbgh2FWC+uvie5IkCZkIBWP35muiMpUqtsGGWPQVB
pAOxOl9xHMsBsA813pvhBpi2KpP+G8PeZpYiWTcYUcYq/5vP4aGQPVGqemFfTUXp
ikfBaT81Kvj1UQ205jaWnZudp1BhHYiXj+vta03/TPg3i94Bjhy55HUN5jk6i5pd
UfKDL7ShOX8OsRU6axRuxuAWvJNJP7GlQpSe+C59FN8lEdydw9ONRA6YGp+U/9ku
m6UzwghONSl7FJBNvG18scjjWIfG4ba/Gju7ZUDQ5TwPP6eSySLIlse362RNWH26
YLtkMytr0D0IdDfjd/wYwSvdnR91aZjAF7T/ny/KyKgtUZr45RvkGOKkT8pxHJBT
C+xSg5ENIT+t27N/VbtXz3CDC81orx0P+HpkqwBZ6CD22Ob78KGAqBDnLRG4m4eE
iM1TJc/ON4PKuCuy2mjbM+/xr1lZS4UFxzD3ZLMYAMMI6Mx5sLQtlMRSSY27t8JA
HsVIDgjVlW4V59sREdK9pe3IHLYwknyBQULMNqUzWHCAfg+7B5QtL+0B5Im4o8qX
aBAOr+iSJAT3yzrTzsyBIMEO9RgHgVMW6OSDzgifEMGDzbqEJOyj8uIDQweTpGke
rf1njCbUwCKVMT4PpVndmC1cgdh+5+eZblZ/iOY8sPgXNL6DYjsLeXWZ84RyZ+fT
fr9uHnpebjEArNC2WEH0YHZhkEKTD2NRnaC1hZlRNVmyWQGD31P5wOznFrzC3HUk
mW3r+evfKkXIo9R6FqjkNUYDGMXEeBRMRYThozBDchx6qBc6s776u9z9xEPlfZdg
dtgjEcU5ezJwvn2+ZgFN8w4T860WYK5HUK4100h9hu3MmC8oaSerwHrxVv2zn5SY
vQdacZdz8CQFxNgmeILtyocYrhM0c3SVVYsfuAXgu01Zqq7w8vSAvURhulaHJvD6
wbPbj9QIK3OyB6kAm0bU1XHDtMUwotEp5YEH8y4ia3Y74t4K9IRhloGBJGF/Et61
IHK0FC5WVBlvIsYUhe9Nrag702EnlS28tG5Whxu3W9Jj9Fo3r7noihR95/zkkHgE
YrObQZxmZ0FEfyyi1nENFSTMvP7Dx4DZ5b9Vn9S72cZ5UYUaMY4jEXx7SoMi2+MN
RZPV+Ed/q5hg+6AqSeQ6PuSDFnHNLzcVbdX9QA7vJyg2PDjvZtLcpTEyylPR12fm
sBZW2Ve1Y6GVY/Sp14KOjIicBOkHPrhh2Y31zO5oehkna6Vaz+HkapzDYsfL17j5
ix2rxpnMt8++2ApH8XehZKsx+yp9IA3D9xh0tvpmZABc80m4w+O9Pm9SNP5meZgC
yFFp4X06kQfiWREXg5PhVjp94NIb8jA5FQ8Ax401tKM9T61FaPMwg4g2FxRAFZQO
yeecneeHt2R1vti5wVcYqqj9nn6Wqk2okAZgwcpfj4c3Ke48GiInKnAOTNrFmMRb
ol1x9GhhZbpIZbUJpnLezq5SshE6Pbc+6TnrUmrfx4BDUGvirGnMcfVmEg2KcVm/
JqquPKaNaUNFtH3Ek4GbOqNcIDPI4MEEOr7jGVRYATlspj6ZaLcg6YC3Y1lBonmB
9m5jxGA3ye0zK5ViGQ8wGQFIu4Th2CCij5IIAg00j6ZfzsYm1eSzqUDNNEV3GaTo
NdhV99MkSo+NdZIcp4UISrtm7yRUdZlkp7CgW8buq2HvbqOY9ToYG7qHRBwv6gEJ
Yfd1MncjTbbkfJQ1CtL10eP8vqfRTvMEZWZfqrMRkgNdbupWYacHWlzMMI8BH/WV
W1DdP8f61ynxXc98U6vgFT8q2Ngho0mGk7dHZuW59spdQ4L/7kJSSctyDdfh2T0l
/2osLfifOMg4LpOG1E2v05poTPtXM7tj2s4M1eTwHbnp39xi97zHkgFQesOvGGR8
gwzslS91yTItjKCbm6spjNhp+tJv21tDBjkRI0+X0VNFKGxm/q8oryKjXLQqnL4o
dnekBS/oI0U3h6mI8kJMokmkoRDyKLPyXEo+JYS5jbZwyH/ojouhymvTZ3UKHB1W
xjBn0QUvKP/LPhA6uLCQHHAtSp49lSRgNz17HHw43/vmePBg3hM5U+mE+UtBRFcQ
oS/Bm09yHI+DoeIBpLNSfg==
`pragma protect end_protected
endmodule
