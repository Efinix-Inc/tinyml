//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2023 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = tinyml_accelerator_v2_0
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Tue Feb  7 10:54:40 2023
// ***************************************************************************************
`define IP_UUID _fc770eb8d5cc46df9bede998a24cd569
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)

`include "defines.v"

module tinyml_accelerator #(
    parameter                       AXI_DW                          = 128,
    parameter                       OP_CNT                          = 5,
    parameter                       ADD_MODE                        = `ADD_MODE,          //Only supported "STANDARD" / "LITE".
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,      //Only supported "STANDARD" / "LITE".
    parameter                       MULT_MODE                       = `MULT_MODE,         //Only supported "STANDARD" / "LITE".
    parameter                       FC_MODE                         = `FC_MODE,           //Only supported "STANDARD" / "LITE".
    //Convolution & Depthwise Convolution OP Parameter          
    parameter                       CONV_DEPTH_MODE                 = `CONV_DEPTH_MODE,    //Only supported "STANDARD" / "LITE".    
    parameter                       CONV_DEPTH_LITE_PARALLEL        = `CONV_DEPTH_LITE_PARALLEL,        
    parameter                       CONV_DEPTH_LITE_AW              = `CONV_DEPTH_LITE_AW,        
    parameter                       CONV_DEPTH_STD_IN_PARALLEL      = `CONV_DEPTH_STD_IN_PARALLEL,        
    parameter                       CONV_DEPTH_STD_OUT_PARALLEL     = `CONV_DEPTH_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTH_STD_OUT_CH_FIFO_A    = `CONV_DEPTH_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTH_STD_FILTER_FIFO_A    = `CONV_DEPTH_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTH_STD_CNT_DTH          = `CONV_DEPTH_STD_CNT_DTH,
    //FC OP Parameter         
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,  
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE   
)(
input                           clk,
input                           rstn,
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
input                           m_axi_clk,
input                           m_axi_rstn,
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);
`IP_MODULE_NAME(tinyml_accelerator_v2_0) #(
 .AXI_DW(AXI_DW),
 .OP_CNT(OP_CNT),
 .ADD_MODE(ADD_MODE),          //Only supported "STANDARD" / "LITE".
 .MIN_MAX_MODE(MIN_MAX_MODE),      //Only supported "STANDARD" / "LITE".
 .MULT_MODE(MULT_MODE),         //Only supported "STANDARD" / "LITE".
 .FC_MODE(FC_MODE),           //Only supported "STANDARD" / "LITE".         
 .CONV_DEPTH_MODE(CONV_DEPTH_MODE),    //Only supported "STANDARD" / "LITE".    
 .CONV_DEPTH_LITE_PARALLEL(CONV_DEPTH_LITE_PARALLEL),        
 .CONV_DEPTH_LITE_AW(CONV_DEPTH_LITE_AW),        
 .CONV_DEPTH_STD_IN_PARALLEL(CONV_DEPTH_STD_IN_PARALLEL),        
 .CONV_DEPTH_STD_OUT_PARALLEL(CONV_DEPTH_STD_OUT_PARALLEL),
 .CONV_DEPTH_STD_OUT_CH_FIFO_A(CONV_DEPTH_STD_OUT_CH_FIFO_A),
 .CONV_DEPTH_STD_FILTER_FIFO_A(CONV_DEPTH_STD_FILTER_FIFO_A),
 .CONV_DEPTH_STD_CNT_DTH(CONV_DEPTH_STD_CNT_DTH),
 .FC_MAX_IN_NODE(FC_MAX_IN_NODE),  
 .FC_MAX_OUT_NODE(FC_MAX_OUT_NODE)   
) u_tinyml_accelerator_v2_0 (
.clk(clk),
.rstn(rstn),
.cmd_valid(cmd_valid),
.cmd_function_id(cmd_function_id),
.cmd_inputs_0(cmd_inputs_0),
.cmd_inputs_1(cmd_inputs_1),
.cmd_ready(cmd_ready),
.cmd_int(cmd_int),
.rsp_valid(rsp_valid),
.rsp_outputs_0(rsp_outputs_0),
.rsp_ready(rsp_ready),
.m_axi_clk(m_axi_clk),
.m_axi_rstn(m_axi_rstn),
.m_axi_awvalid(m_axi_awvalid),
.m_axi_awaddr(m_axi_awaddr),
.m_axi_awlen(m_axi_awlen),
.m_axi_awsize(m_axi_awsize),
.m_axi_awburst(m_axi_awburst),
.m_axi_awprot(m_axi_awprot),
.m_axi_awlock(m_axi_awlock),
.m_axi_awcache(m_axi_awcache),
.m_axi_awready(m_axi_awready),
.m_axi_wdata(m_axi_wdata),
.m_axi_wstrb(m_axi_wstrb),
.m_axi_wlast(m_axi_wlast),
.m_axi_wvalid(m_axi_wvalid),
.m_axi_wready(m_axi_wready),
.m_axi_bresp(m_axi_bresp),
.m_axi_bvalid(m_axi_bvalid),
.m_axi_bready(m_axi_bready),
.m_axi_arvalid(m_axi_arvalid),
.m_axi_araddr(m_axi_araddr),
.m_axi_arlen(m_axi_arlen),
.m_axi_arsize(m_axi_arsize),
.m_axi_arburst(m_axi_arburst),
.m_axi_arprot(m_axi_arprot),
.m_axi_arlock(m_axi_arlock),
.m_axi_arcache(m_axi_arcache),
.m_axi_arready(m_axi_arready),
.m_axi_rvalid(m_axi_rvalid),
.m_axi_rdata(m_axi_rdata),
.m_axi_rlast(m_axi_rlast),
.m_axi_rresp(m_axi_rresp),
.m_axi_rready(m_axi_rready)
);
endmodule

//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nrO6ejqDCYTa0ONpO0W7AEJfFo5ZfmzLT5LvANrpYqYFyhoHKIo2P2LLbWPrEU0C
SSKZBcLmFsxBmRH2tk2m6XXCdHa0zkx/lWEiVgWI7dEbvHSTEnm/pngw7gFLVEWE
qalwVbvfwsdbJqH27npi3oi8NEM6B9SwKyy7BIrVOS8mn9X2E6k3fOvSe5rFjNeo
2l0M2TuUFTsDmHkYQ8h1hBkUbU1lGgoMeidlmfAsLw2ZBLtS2tUq00GM763dM/z3
oYSFAiCN7Qe6ag8YUjakMNwO5NS6Zyt5cV0G45RX1arI7lduivREHNmy3KR09YRg
lJ5mbvZ5zj/zNFAno/Pg6A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1200 )
`pragma protect data_block
uMUBKCD0qoa78zj/tW6HzpT/tc2Ulypi2kVVaaNxyXYAmf50H3heXLzog8WRrYGE
Cex74r1odd7Xdqlo90ttuLr7+E62a/w3ahOLJhtVv2D1nMay59SrPAGD853J+w+h
Pho6vQo0JhJ4wj3e+3Wkrx06hT9gkdF6NjH/AO1kmDuMkYgNG8+ORqpunReyrJCn
mvGLfZRk6F+PCpHFwyogG/YXtgnyLIxaL/KppC7YljJiwkYqBH9FPNaqDdOqXSRj
p/nTCdczIBM05pdOjeKpFiq41CX7u7t07yKlBiCCMxaTNdC6AjYShzOYdiB8IFcp
eyQdD5RAWu86UyxQVf7M2fJbcRoa7d9cdRBmCRb89DX+SEubwXdEO/coLhiwiS++
zOOvklpiJot5+KlUNeIjihBByF0S+ApYLi3UDXaee2uTxmXj4IUki5BQTw4dmuR6
eRTjh915Qs8HuKWnMXL5yWCb4WDwdCtNQ++MBbbfrIcdDP9Icshxl2wJ8OgVOWMq
tW9z2A8htHI1qi/6EnB8R+pLZ8m888JKlQ1+FqjI6ImHF6uSLL3ydriLAHZGcsuT
3CFdsp6yT23l/SN89Ovy/4hX66DptmLUWggb5OUOQr6yaTi+Brp7p2sfOtD3b9L9
bebt6Hy0biz+JgxlldxZR1LGMs754mm21fMItB+3suMf7EUEwFTp5jD/qR8WZrcc
6X7IE5qdGwM5Q50W0gj7woBY78G0Yum4BCy4rFkD2PJaImq8bPEFjZUMb6s77fDI
wsMFaeF+Hq5rVQkwHczclxz2N8/GvAXFdeT1cI3lzfufisaPMw0xYTvLEPEpOC84
uH5Gy05TIXYXHtnf30qFhei841VCcxF2HCkh0I4JUuFoqSwx3b+h3Ob7QK4WKYSk
cFUEVIuYQ97oXfXuPBqrfO/dVHA2q570CUO0og3oZIcQawAtYSVMnNKJpv6JI0h2
GSWJpBLQE1l50Pn04RVt0xi2D05kEUjIpJdKkD5pa2EzXHH9UQ2g1u2jgBZ6oVpA
JOUoL2nqLv1UroiPlqFuptiNVsK62HOzn0xVSk4SoAWULEsygpZWQcW+Aj/M5CHU
Gy8FJ7aVvQbXTd0+wZoUNYcGJasHcs/plkOsDmZF8CyKzrDwSdMzSx7taO3h8ad2
ESfY+itNayWiGwry+VwlNgM7RX/AUiB7JJYAUn1TTv8b8cS0RRtX9CCXNIEXVA5m
EhW4d6bxOfm/+VYQptz8fsvHcHWIWeYB+iv6yemwEXCPP01B9t1BVQgzje8ZG6T6
yCPTCI+f9iCg6/l3KEEqxrO+GrVDAZsTpqK7dNpYl3UCocKDOsFYWVPfYy1PTXOR
jGHNipJcIA82bk5oc9Q91DBf0+M1h9cWyjS15JBHC+2N9BKODLRleGoR8dWkPOos
MAxo848vAN42JMuSksYUuLh0BjIU9OUoDf7ABVcUofQzWCdB9Gyom1afNPPhb352
JwdNHsualUX+tOy3hhVHhdMzFkVARS9eZDT2GWbGY+E/o6t6ml0bvZFzGB0VJ3Np
0vAPXLcf+PZJ+ZV1xYNMHzDshbujEkIDFd3pPYjkQrCwZHVOHvZvgal4FSzBFZM4
`pragma protect end_protected

//pragma protect end
`include "defines.v"
`timescale 1 ns / 1 ns
module `IP_MODULE_NAME(tinyml_accelerator_v2_0)#(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 5,
    parameter                       ADD_MODE                        = `ADD_MODE,          
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,      
    parameter                       MULT_MODE                       = `MULT_MODE,         
    parameter                       FC_MODE                         = `FC_MODE,           
    parameter                       CONV_DEPTH_MODE                 = `CONV_DEPTH_MODE,    
    parameter                       CONV_DEPTH_LITE_PARALLEL        = `CONV_DEPTH_LITE_PARALLEL,
    parameter                       CONV_DEPTH_LITE_AW              = `CONV_DEPTH_LITE_AW,
    parameter                       CONV_DEPTH_STD_IN_PARALLEL      = `CONV_DEPTH_STD_IN_PARALLEL,
    parameter                       CONV_DEPTH_STD_OUT_PARALLEL     = `CONV_DEPTH_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTH_STD_OUT_CH_FIFO_A    = `CONV_DEPTH_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTH_STD_FILTER_FIFO_A    = `CONV_DEPTH_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTH_STD_CNT_DTH          = `CONV_DEPTH_STD_CNT_DTH,
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE
)
(
input                           clk,
input                           rstn,
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
input                           m_axi_clk,
input                           m_axi_rstn,
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ntATRqM+901z3+wCx1zlCCMXpq07hUdRpV9fFoiVN1ezANX8O6AC71GS2rFbq/po
E8NoiquteEI1/UCQKva8Hoft7iLkVn20kTVSiGKp2T8QAn1Ye2ZM4E3JMZRHoU6t
HsQXaRpyJTs9vq91xC5a5Z4hhGWkpR8ZKGrN2cyXNEOBRp1zMDzfiIYiqiw2J6UE
dyf59nIzsdmx6p7XKFW9QB3tfG0EXIdJawtY1Jfcnf4Q/4ZPb1op4zR2SHy02e6p
8tvLcFMm0IUs6OEgDu3oTFkeHdlTZxS7s9aFT6ovjuHcfYoGTdgu2JnmfVSDw+cj
UTTv48KDf+ZhXomK6kqkcQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 40336 )
`pragma protect data_block
gtXApY7DZoOCHUyEujyDeYz43tM0mGepb23wAwIZsPnlU7Ga1kJvKpDNKsVzUM5N
0n4eAOYXAgNQvcOdwwjmMV3S1bv4m0YdB3Dfto4LRkK6+f7rcgxjI8W/i7455UX2
YPOs2l+SQuw9JGpqXeHHY3lVwS7tGFdjk731pIVr2zrjB8R6xA5Q0zEYuFLhOU01
xQCv/tv7zyAUhOfyPMZnXDQ9Oc2cSPVCLlQ7vK1pf18WurLUrsaGQremslNzYZwD
2EjF8lWzbC1s1MYl35vE+LTRe1+sU20s6WQ8x1YjdHfty7P/+cKd6ceS6BdKwoJ6
PL1qSRVACZARqspW+izMTrjY/m/gcLf/TcPjPJgfzC62UBq6vo+6MU6oJkIcmorm
UXv3P6za9+AC+eCLUyNFbaZ5AZbiAvcyD4w7LODI0HBpYEmo27L0nFf/OuF0yNPE
cdN9lTY0CFBOh9zxMDuo7BmL3GG6TYgBOZbWOYPnU5MH+DmVlcrSVbnQWNHcDCQo
3yvXImfjx14aHS5+wMaI3noXFoUbiU04j3EcvZndDptYuRRVlA+585qf+NsUfTuo
pdJbjtL5prkvvyR/X9oVXgrcu8Q0FYa3JCZ3PTpTNblzn8JFk7N3RGS95loD0R75
mbwKxDOw6vYTwHI6Z9Jpi9zN/OS4M+3SA1gX3WmOKqJhIXvzo5v6xWN0lZT5ehl1
qDG9kDPj4J2em3T6DD/yY9UOGajHGOZhLJhDBDcT466nXy5F8BDAFbqzqO3x4Dw0
hR0wZQWtiDN82EpqJEqqioe3BoVNN0tb8nn5pZ0jR85k8xwdbGEn2TQ2jnwY/0n+
tzdShblgnJ1jyBfr/6gSgW64H0aVcFL6gaG8HhxNlhdbDmNaEY/kT/ZV2HBl7ZRR
WBp+jVIyKjS0bc2MbsOdr7wv6jNHes8EvL3Z8cS4CWVBE5PrVENT86OivdTWw0ho
Q0yO5k//v0XGJr0bc0HNedGtx2P0QuvTUWxngnVax2lovoU4yv0JM7u3NAJc9bSP
R+2AIs2nPPWGyzKDnO5i1Pv/uWXP7yvafiL+7LAmDsjaTn0k9KtnhAmME4sD3s9X
grbFQNWXuojeT/3JQAOnCHQrWWY/q9rC/ueD8Cm6amhAhEMUWAey0RXIJcmgs1/y
qoQwXKcOH5v1aEd6RZkcxIwuBf5fKroG03DvV/58wcEva/zMvca6VNhMOfvE8m8Z
qTHF0JG79FgJDadPp7KycQDqSgGl0bLwNuG5EuYT5mbJ3bqiDPHmH5Z8BNPPYEqt
+miJIuLD1f2M/fCsTKTequJG/ALxh3K9Ep9UVdvAvH5yIPa6PybOmVAYjJwL4G+p
zqhR9fog8Sbf/2Brr+ZPhoZjg6kjRpYPnPT2AkkiImqoqd6rR2xshqw5Btz8AdYv
qT6AQG9B4bLZbhhBPvm2yzAdRslY9aXpv1jkexJ36PItLNTaUJLTi90d3YrLO5Wn
PSgITVqd14I93zvmTDngBy5MguO20730ahiv3lF8PJuzVU6tbmR1DBFI1fledP4c
9oY5hQa+ApbsZw0QR8Bi4AU+l9yA9+CTplOgReKM/taM5CxIvxtKYHsL7nSXd1Zj
080MLqDUcOuJXMBLK+Q6a8Wa4WJB+k4Tb7rthvPPT+1CDANMZkx2ZAmvyXDk215w
uuMs+sSP631DkVCvQah4A10Y3LYy90Oub1u3qLsB3CvjieBYttdkw8deboaEIqjh
UyF0R9xbmdDkS2omDlN/EP62EYZymaTWPz1cQtkz4WHBUBcxtBajAmZs7wNd4ceQ
RdYjxpJvgERXp7XhGRucR1wtBEZUykF0rQbOphKAcsmtF2gSewYE+6Rja8uZBJf/
6ozRD6hj4UpFWChy/qvL+CDe2U127MAxMIJOkRiefQwL3nFnkPqtL4cc7CUjhLqI
go8xyCD1EvdVoWvT+T6hc1Y62JxGmVGU6iB/PP3BRx4vz8N3ILhG+wbAhExB7y2i
4B6wO7sZCqj/8mmGWBr690u0qZETXUVNlm/vh42BHaadpqvix7XOemA+U+cmF827
MgyTVEb5ciQB6m5o6PV4nH/rgFxZ08ygTW6qu8QVa+xGQJbiyT47dAJP9kW6OQ87
DwEAKVrB21lPvJiwDnvhyJyIMWVYaESlOXloo3C3EcmNXngf/ljPeJJR/VEo0Dja
b3lLwFrWWvHGqmV/4vmoYPQ9FjjHKqk7iPHn3PQT35hJBi4vxeSdE/j+7dT9Eh4R
mh/fNet/dMBuGloglbQBhhYpIjzIJMiQH91BUZQ/s2SdBSnLauctoSLuou4qZ67S
DrDRfPaDFk3Hm6FIfvMl5AbZYrewHUkZ97enDX8+1N5a1iWI8O6X5iNKkSgqJ/cl
dDJQ/gsB4fVJqQpGgb+wHCHhLfBPrHawQnFeP0HVh5WY+hb3F4CCiqeiQ5d4xx1f
2yYDGXL8wWnwtmQFHpBdRWhn33FOjom51naNEpTvY6Ch+ztm2wAwqe0IMqhWY9av
wv/dpCRpXR+lHWNcFBtQOR0k92by4pLm6dxgozGOfa3dEwlg1JyD0tzkLlaM3Nlw
U00EX4OIsRQj4RZwqDYAspsgesIPRt2F5h9S5PuUk2o75xJU+KAxNs/NIEkWh+JR
hwFT6IQd8hBEZkYvcvzf67QYfVa7PzX8gUcMhue5/Hmk12QRjpELoXmfyl96rgPf
B5SZ9zInrVlLpF6XsVDzLe4vKc6UBEhvedpsT+18nErrMajptjdXCVGGW3/5Rxqu
KHiSEIZIbUzON1tDPIgr8dAObWSVmS73f4Uu+GL0BgrSbKicLhF2mnqZ2wP3mmSj
5Q2rxyjWf/mZkPYoTR1wQeSpUik7dn/SW+ZnQ2WJl5OPuA49HiePWojYrSnhqewp
U1n6q6vMc7bYKDNOupeMBByB3w6xLFpkzPGqUhVqzmu2vqL1ybGY0FZzea+LIxnT
JMDVhQTFXafEuQa7kJlSGX/rHeTq8gNEDPuD35FmNjrUyfyDj+kIR2LWgWhu/UvM
EauhTmUQ7pAzvUgkgKd4XGJIryU3gtOrl16nQn0or6az/9r5Y2FRBP78bZiIPu35
NTk6lDiCK5iSy00UxCZNL1d7IUq0pgLUkHfTE23owLYUxI15LO81BI4HUwZ90ioQ
didHug75ywEdYzs3ACPGzYSVrcjJ4P08P8QR2moM6pceI+j2A47gl7pvAOvw+tEE
0g7eCo38iyoOGp05OqMXZ7xUB1GOLFFr2ssm+JB2IWFPdyEN673nWYX8QjFcydWC
RqbvBl1dg4l1KuzzThfdmuGGi3FQLBL6Z2Xt1JKF7InICiMB6GpvGGxqn7B00rPy
sLYL9W4P4ZnkBbuI64/sqA7wSMvgaSdY2UwNdiT4cMSC8h1rkwJKjMt960SXhSUl
TBV/wmzBhvamAbxB5ENoS4RMPUJ+Nge4zAZhHslCHrt42HZKVlv4Jj7Pnysd+eMv
ndydV5o1N8qFxHB4RfsBzy7zrHtoVUuQe6v+ZyEEckniGZkfmCwkfL8IdPt5G/4B
/St3HNERLb3RuQFIMDIhytLARt3nc9U8tnpU0ELTTBRFvxUyW0R3lQ3hy2LDGa+E
QwVHhrK2o7sXo+uIde7dTqNOE7KhU16E+tlW9LhQistq0ullo2qe57XSUCoSWsw7
RKRSydHrWXXzsIsXZTb+yipKftcGLVnJtKss9pry4y5KfoVzvNKwy5wz93pq4dW0
kRsuUOodjaM8MLD9Ti0occyTRlgoTcbVM8EnDCyz22gTxXbzyqnifMlSXHzlYjOh
MGYojhXUvPrRrDpLjI6tLImTzIvcc6ngjd8Ad5RYtApt2mTamQHSDgVU9sCHQqM5
xXzrRwPKwC1B9lD626njJvJQZY1jrUUDhjxOVUcqxmpf8HVERoWQJfSOYJIbpbE1
tl1iN5PWuaj/YtfgVbiej2XHTaVOOrzBaouXovss/Z321NyU4KRlKdv2arbOG+UT
YoUNfxNQYRUtNYuPdoArXLt6hR89tLPX+RD6cfRwRzfaMnz73bQdda/hIqj39KnL
T1mR9mHzulBityw5Z4R++Y6Yfyor0RKbetfaDuiBs8YI8RzGnoS9ugRte2n252zJ
v5l4l4i9qKvRNqVQuQZpKd5BShN19W6we/qvk0jly4n/5lPQDEAPA5GKsOOy8l3H
mUBFqzVywrDVIBhgjKyjXfx8U2EbjOz87F7Bo7wlujOpBlsQqAil8T4eT1e3fjOO
Ta5pwaOvPBSBVoIp3UCUJ+g7ys/WxC6je6XG46zCC6pZ3ojv8TYI7AKG4/VHh76X
GIJqNB9WoOuuQttlbsrFh//BFWjQW8jRQOA5I9eGTyi3WguQVed1iRd75CsyJJJY
zTsTlzXnqheYDU3kP1fPxHQjaN4BbonErSSMOC9PBBkRez7p6Ni0d6U0qPmwL5sY
KW6dEmI0UDLgNparzLr8RyaQcejc3j0HdrRymjeGOIt7sr9CwJr2tlYzz9i13vLs
dyAbxP9nHpmZK5V2aS/McHMMnJlQRcFPuP1MyYKf6zKmOPKIkHe5iBE/0kny9r6h
nhPdPwTs4rHb1+CkiFgMd/ZPaBYAgPugDr7TyySu9eO7F+A0PjyIqmF81ThSo4IM
Jcq4c1w6ye1opYqfqO5KPFi3rbo7XNDBJaAyPKFRfXELOHcKfGAqGnbEphp160t5
GDn/Y7+J2wfcoQH38FKNhheDiGK1pf4w0oteJcQ2ftwjelvWhGanJmqDj0ZlTVNy
iO45oYjTTER6BrxCFGbw2bpeaBSkl8nLcog08Y+Qsrl3cxb2VTPEYr/q2JCaUhvV
sryvykbQJaeszlWUHw/fTLWVszKE3qEvGlaBiEX8pLpm1+omtId58DJiy9TnxwvM
ymW27sr2EYRljQGrK8NLZlivog9rYn05A5cddo3IgTMoeYY6EQ0brBAGAO5Vj5ro
eKwxWyrKWF096hX6T5bZG4FS2tC5oCKc2l0Q4fluLq8p3LmY6Rau3l9TNh9I41Bz
x6UF1+n1+klynPuvt9DnuRvNaHhRuFrVw2J5EQbZIOjA/P5Ye5XKwOTONW5ESEOh
w1PfnHK8GwTJHAFQbV+k1LVTMJvp9+2pjbVgSFcA8pEUus9ZqiQWXo9N4Uz9KYZD
+6swHqKqHZGwLAMgF2L5+2fajNpaCT2nBXHZX1OBTaq0dBeER8hdApJB+o3Rd5V4
Flo31EWbHzuJrjl5bUZqHGdNj30c/i2Xw5YyiHY1d4xuIFZ76Epqu3/PorF1PAy7
Eapb2fH5iwVmr9z78uFaUZItqBRM+JyzZe4H5xqz6iQ276r+QbvdFFyV0x8aLoYD
7DGOJ79YpoV/YKFuzVHcR/KKtVhKDcMCK0Ze+4l7ISlOFNcu2i80prP6vDu+ZIrR
gAeq7818owsgo/QU8zNp033qzb5Pujy2ISkcAR+RU9yeicK2HsoylH2BO6bxTBng
oQo+/rV3V+oH0aGklIXEMiEgR4a+pcbN3HKrbPCcV6v6uynjlde2+fzJDWUoamIk
HFa/yQoPMYKEcDG4O0xFHU9EtRvgNqdf0F5FE4Eg7tpsyQC0Yx/a7x7ru0Zb1PFs
Bo+iUg3hWTwRweQNpVkxLHGy/diScRGNU7pBWtNMsAWAzOT2Wy6McMvkjOVwoRHr
SKKfdqTt9J7RYNJu8PvnpST8d19RQTSKspGjoCrQGY5JeLumXzac9JZ2oWweOLCd
FHr1b2wvnPhRYaSuhVmmzmMFVrUAcOPZsNAXp7/+BfTGpqIyX3+o07jHx8VD0XBi
AKj8wC7NNfozxdUUYmrW0nJbIaSA3OQAjGdoMom3cSC7lvKaXz5/5tqBodtHaIPn
Rsx2xyRUtKxCmSmaMKAE4ThcTDncNdPR8ESIYQk2GFvkhBamRAt4EoWRsoV/5ZhU
w22mmF6gl5aPw6qCKp56hh9veRKI/nNo8NQcbX0dXgNogkZWZcfmiv5OG2I4FaWD
/HFyo5AB/z0JyDe6ZD/2TZyhFLradROO3pq6gXxn3C0ioVUfDh2bSf9FTvJGDadz
XeC3EJBTaVqphT1VX0HxWma3f88bJu+NG14FmBJ2TRDjLmpr1x+lSskocbU/uqv1
/LtRXc8/ESJvPAlzdNXw4YUwpYN0jH1VW4qbWI1824Y6w4FfkcG9km/hBVEXjGGe
4ZB2qyMZJwNlEHgUubJfcrxd/BgAc3N71haotyX+u8ydCv+zwpYuzEvdD/YpVaPw
gHoF3NAAQtD6OJMQb2AkXa5+8lVrLEFKbgn4Ubz8F7UWXLEWBXso7n4FcRRDlXfI
7gb9FJWfJ6Yk+3/C7uELDpI8S3G8+AaZ5MnWmfeJbcR8/e+cRhZmnB/zz9PzdOEM
la3Js0QHgj0uBSO9NTdpcDTT76DE/hO7zurZOPEwm7o3rjJPCiwohZQXX+zgqleL
t66qRM41Dtx8VdAaGlWPR/KptEMTYsg6In5kaii5XIPOce8hNMdkNjTOtMcI66Ja
Wk+P3dEVvDBRAuiAJzv8/D8O3iz5VOyRuFDtRDFJwZYEHwPvTK04E1qGFU0j4vVQ
FhROMcJhPkqXkIGCLESs4G4TycZDYTjjhcBVVsMc4uMTpFzx/15EHTd6UD+R0crf
s0/HbUNXxKPnhypswkVoQOs5aXVZzuGG6VFIUUeLqtGSGUHFnOqXIJ1ye+/thhEZ
adGwrVw1KIiEyGBAMcNGP66I2kC7E1mKKnBFv4s9CwEiHveBvG1OpuAlvVnQGBTk
x2/5E0Xcubtjl2MoINlgKJkQcIoeCsJAnlrkC0OeFa6G3P7AzMM4BC0RJVQVx0MX
vU44ml664iW6jbbdcX5wGo/bAohtgh3Cnicv/PDJ6Y8ZasvPABoG4notdILDnAYC
bAMiYZPu7MO+qDT5+LdJ+fRC2f3774CKVrM6XOASiGyxZbqz+zRPNyjkyTSSSt3L
6qoOi9KA7lHSoUW6tdXGCG68El1GCqpy8k7EuSHRfDWBjvd2fyanZIPUXD9mhq4T
1+HV7vrOfwuQ0LXkQ115wz/ck2H6h341cTUAQdpc47MPnE9kk9lpOczhEOpfysmI
ZHI71r2ePC4VGt8bEsEs39MiLbEdQwbVar9fagrqyxoW0ROdNxHm4vEhGdTonY1t
4G6+UkguHNz1R6NIYQZNQMo4IYBR9bZmVEcSCTBGnbn7tr9K+yRyDNMttWTiKdzq
l2ZRH/4631cvVWrA57NoWwzFkM11L82h3KPfFmWW1mmYi7SMQZI9Hhf4BRfNZHYA
BBMS2Tr/xLXySxhpoHlamEGPKMs0tg6fxIvcFc2LT2aWIq3fg4nbna+TWdUVJiqG
kSBmABUn6PH5qCZth4aBE9D73gTRxk8U/gID3tvYaaE0/k+ctx5MJW0FZHTFxFw1
jhiMNKzsVq86Wz5/m4u9grtvV54DER6idgsR/vc47F2LzHTIQ5uMHIW2jzTdg6Hp
Fnn00CopatYbq8l2jgpeWwvSS7+oHSoxceFPAXf1oROxsAWGuROW2FME8Tj3GWz6
HpFkDhj8yMe4Cd+dffhDETGL3rnP3zoJyZUE1dgnkcZq30Y3lT8tVUtK3vtDAUTD
L0Z0xhvF/uE9gQhXNeNC7VHnqqGYFny7rI35s6fFJHqpRmpig0v0dzxuGywdE/jA
Ed4Nul7hQtQ+NYg3cj32wE/hGNGyYYaG/ai/LI3oowhg7I1u5YtiKswln8rt2wM2
nJZKVw2XSSOeOgDh5YDBGEmpxiipagByFp4okBiJFUaufnoRb+kxRBVKxN6sbJcH
n3aOdwScs0Ypcn9QbSRXY7R7AcUYv2vCDjFZ/Dn5J9IjumhdAwvJhY4jO0OrJqo+
KV8KBRJ3fur3eDk/mZJB16YID6g+urwoEpfaoj+MhyHZauBYYZ/HhgSc/5IKV1oM
63Fx7JsH8UHcOUmVhl4A9EKbsB7xjBtsRLeMINGoq/DJZDUEFp0cZ8JfHwjV50cb
kyY8WmJ/NFAS0gR6X4X19DnoFCjZ3pXwQY5QQzLGaTkiSaLC5S/dvmHtsqA0s+hk
yX2SxUoX10D88zrCgq0OgkoBOmU4jzIWhNQ8QZdSCyZxu0mtnYgjMRQbzKF0/gwt
K9LYBXRdJ6WE2yzTkNCnI9I0bDcGuuxTWMi7i1VMWkBUyym1xz+AK3wmRG8wbBHp
rJqG6lVhyZqRZVIhsrrlutD+WDa+NjO/nLNMePlDny6t+qFiap900cQOR8WPJlJm
p+5MidfZqnaqQVpPppDVejMcHxqrKTAXT8nzA8cBKfln3xgOicFMZl6/hcAkiRgH
/lkK9nLQYcfV73ij00TE3Zl6E/WatIPbyCKlnTFNncW3j3e1SYpsQTrUq6uBv0oj
WBd7PKORBTKBMu1NBiKVYBPcqEa4jyFtM0OYltktyuawAbhKAqOo3eFVHZ5I9JQ9
/C7FHM5JDV5O2QS0NnxG7mwCob2C9JJV4XQKUD+N6XZQM5+s4EW3/vBybo9iTkgg
IP/Fvnsurmifn0XY6gLHjrTWZRAbb62LwQS/2fsawBRmIJNj6923v9cbuhCjc8wR
ndE/MEbgNRQyT6JaLlEBowcmn/boSn5gzjrl3YsmBQJqgvXJrvjZaRIgMxim8OZ1
xWv8FgcUWd5LAUKgVAXmNOED5hP5Og5hf4020/U/Ry0NupQlcWrWI+0ZFb6ZPrfi
eYSgC8TjA/+dV8P3PzekmrlErRv3E1O+f2dOGCyGiv8fHJaWRy6/ALi+yyGFgxym
Bk/yoxscv/oLEU9/Da/xsW0sRbTjqub+jP8P2RjF5aoXLYcLzY2gp7nvKB+5LQN1
M6dWEJYs2YD15rKnjILhCF7r8ZYCiO2QzpgoF9AR/I6y6E3yfAeY/LPT9FAfQW71
0AfB+rHQLjWMe62oWcgbF9E7jGdWiqZW9XwqAoejqk5QWqv/DCdivNykLPocFdyo
2eJ4rxbmIpQjBnk+/5qrLJKO/wUgXZ2xUSOT3FKRLfuT/fe1k7eVRxPM6Z2Ti0GG
oq7SY46jkkviThfp+TOyVsTLFgQjUgLPCoRCFvbkCdTXZL3/wZlHjgmxSc+XTScG
xzqQpFP3374dMPDDctN+5IWK/G1gGmyP8z5n2o5ChIuZIibAUnQKmcCpDkbfsWp0
XLfay0NYp+k2DnJML9wjqZ963kdQrhPRwv8AtYnFVsQ139hFK6P9ATY5DixVPYyR
iz3+y1yoQEa7bRTmkBvS2b5A4gRsyYCLXEy6waUrMvF5mJBoUzfTaFLWQ7q7i3p5
Tc/Pu+Ejr48b7pULOBoEzQtmqWsYkuAGCy44SvpPrzW5LMVSi+idVMtxwwx+TCAI
4D9dlLz4nO6VXlfl7JDw/elN0NQXpUQVYvWhT5CPTp1dwAZw9fArEQdnougXJE4L
2aCEpuZ/ExrLWvzURG8uSoilNipMbNbaNSVeJDn6evBmzpFicVCdKK6/LzwrKd9X
5DUVEao/zIdW/KDfAeJ6SB2vH3y4Wr68l+rw+gwm7sPt/IGqsq+qTwyRwVKoHyWp
PNdS6xaGCZprXw+lIClmcw48ol/g+Iu0waogIAV62lnfWWld69eBtvl6NoSBt/1n
KlJgY/m+siK0JupkLNeCORmKD6gGFaCfnWdPNNABJnWNwQGDS55TkqzRazj8YHis
d3K4sQuhCSX3t5hnX+XtmE+dm3Zg4vUkFnb4tNrzqHXNoAW8MVuqKBuS2FLboFzE
/QqgrpUUCXqJ9pu72y3WTEn6e+ABD0j2jhnfqbZrDjQMHshEwlIMAfZedcqkTyQ2
KxY6OHGtFYl7LlooNmUwq4jKCpM4K9ftWUqVcLATpUEkU2Ve7MK1KBTuZ+DQbBF7
kHyvKlKom9+6dbP3jmrvSsEMMbkMSKDMy89gCJKCop1HU5BKO5QtnPtDLBD96/yB
k0XDZLReLtospB/+lnclH48/YxaVBa1BTpl0opXD+HEC7eXRDdtfhwU8IJWJ+DlN
KNIVCermCtN/VWPU5vM4iYpsFEQXhqmoXLsNjYoLkQosxmO4vfuV1/TBrHWcQnIV
RI/HhzMqg028AOkptfX/eL4jaUAcrIAZVhZtoAv1scuMXD17M4yyocQPlN6FE0bO
eudYzLYfJMnLkUhqdiatItL1IHXBTKc97JoHh/SKTJN8sy7Te6eyS/OijR8jTCAP
sWPCkXwr5kfsLVn8ujWbBSZtcsWWalm3pK+xoA7daH54hD1Y3LK8eQVhDT/KMEO+
2sWS7t9anpEoQlFdW7JnpUUe5gotVfFPwZ1wTI4mUifadNKTFe+jrk4zzmGZ87/+
Uq0wrQKq6tuQx+IM+JcVJ1YaCoeUaT6u9UQ3izSdr5oFc1mb9QWdXyB75jHrnNVn
gRXcL9+V5nvNK2aq215WrC7PRa4bIpNt4IrwvRCI9GLr0VaxADQA6S+QmMs92nnK
p5yrbutKiD0lO9jWas0ciYNFtRDIHBSN+wnqnxYUwHSFvDA7BseuGCC/EsSGMJgP
GJcjgzrUEo30BIP6rpYQNlfvh93Q7kpTL7st1iVXK6ZHiRoQHbErQcG8uh/OHYsN
9zjRVODg7T6YcH6Gzex58EOQyw73fHQNsSK00DddO4/gVNLn4Dw1kJDt9Nau8IsC
itS7hFi3+t75gSLGC3Ear6J3PwZk2hI0eHB+Ky8nWSYPmEkVz6UuU3m3xiqaNuF5
6KL+lGHqAIX1KODX6TYQ8jWT1/wJDQmxShETDXrXd89cd/xRBk14fa/twEQ33Bth
xSuDGr7Dl1km3Sx5KAe6v0u94I2Lq8tlTR6DZxbbUUv1xYDpvOlUwH031Z1KK5eb
VR/vJ1yYJoaL4/1KUGkPmMUL76Ho4Fj9lKE0S8mN43c3BuCioflr8AZRc0hH9YXO
vjvH19IsprY5D2Jp8PSEbKNk4oG4KVQ/PqdJzYPDjtkhQ1sdQ7fSSsm+kMY06x6K
IfC3AcxUZFGFcMqbuENgBhoJdReX8bDbDDFmMJjB++i/q0R5LzgmDPvLjh7DunDQ
AhiaLMt8UjZxqX1cmsfejZ/rIDTnmspIOY9lF13iHgg0DH01ZLg4c1303dO14i7P
Fe4oKvTDnY4dijgg2taPM/tKhR49a+w05cnNQoDVLC4+6SuQDqYl2y6xTaQB82FU
Q2SVXy1PEN7KKUDXK/Ynk66aGaAA7lZVEmaJRDDsR5an7M3ob8vIKMa4TqueXQxV
uoBaGyQqGRm609edIobstDQ2jaW1fXMljQQw2l7Cn6mcklPQ5zhCbp6b0vDMgj1a
s9nDaNCJoO02/SIiIfvTNvZwuCq+PayWAGEpjazpQNbpdQ9/G6F7A9wKXmf91WPT
qAu+MsPHM2KgZ7QMgugR0xB6oOQxbYbkzdXxw9D1gUXOM1b5yAtl67rTC5MS7JPF
HpBt9Rwsz48TBPNBsQigOIcShaxSpD9wsy20M+4PIGFYzXloZ7s6o52PYvsLo5Wr
6WQgCaQZR8yjYq+/ArPTK1kkuSOj8my4knRQVTpXWt0ToFfOc12mbkKDZj/5mBn7
jNmKps4bTGQmq1oIQBdFZf46wuGqt95fn+GoukgsUk14yhwDPfiPl0BegXl55EYb
o/P1esxVq5coWdeS57cVmtVsZkl8wiG/2LvY9vfyoFoqXFNWPNMKFg5PBI2q1Suu
9CTpXgxkgybLK7dlb3wabQaW3BQddX1kz1ZhGRR4UvuklJX2tBJHMolG2K1CtLpJ
T/XNoJpblmE7fHqZJKa9d/YbT4obBDGbdpTOXrQjkdsMJ6/YdSphCgzmbEKiwEIr
noPih4aMDR9SRW62m6s4TDpD/hPdsSK270I95Qya3C1Ht/iRnomS1RMFug6BTHiS
Vft7m8hE4vaLdXisKAW8c3JmmkSj9hG3xsYbcVUXK4WE0ri31/kW7k8n0psxPeOJ
S4jQs5Gow2S48wngckT+VwxW9M0aXQogWUf9KVMx9Ucu+6qXOiaMFYZxg7Jn9eSU
Ts/SeqpP5VBQS05RYPjbZMeB5q1c/hSdI9MOAjlGE3yH0+ZKCkU59GmQdjRXDowY
Kepkt2yEJLrdNwtHkdmkwLwz8tCWHTzJITcOzzUh+PrsvFrCt+kQz7T7QGyOQFF8
4QfN8OCVVhz0SQDXBTl6YqOCme+iSFanGAGmjivQ2GGVzX5v8aQ8b+yXO90Se2aP
zLXofsbZz55nBUbeWb7vjq9RohaBwd2mEIVJzM1TSZH3ruQo/PCkjQWTuq+qG1JH
DMtKxgyJ6lQ55ncF4B+4rUS9IKBTT9iGNjTIeDjYNVEJSPA3EVsURTPbrvDHso18
xUpHW3W9UlySNVOfUu7u0WHpwvfIHzWRAc3IecBHmiGgbLVGyXMmEQeRwQX1kzm7
2bWCR6E6B8kSc6fnahYCzpwyNFiCzE7UPayCq08LnpxANBhe7h5y7IB6weYF8k4W
EFHizqK8zFujx+fdXh+x0Ia0rWQvgUPs0EeqajIi49H3wN+AYRsgKAUV/rS300PZ
XG1pV0t8yBTTQEtIdgC7RBvtfev8CYEIcJdvtdll/M22U45KA2jLTQzSMvp48Q8h
F9IgsVKhff5qIjH6GG5rI5ahPRDXJuL+Ym6PeDQua0rNZrqhYnN0mIQU2auzQkrc
OdLcbpr3hG8tGR/7XRsfRPBw832bd0CBx2RLufyqe465u1BYMH8pFS5j5wbrw6Uk
jU/AARxJOusaYSZxmxiVY2yGoQgqKLm3rdziHOFoCvQ/r2vnvw8TS2U3mHkSiJpi
HKTSJU/HmQ0pJgLxjcgnlpZqwn2B12v+jVocyzxaW+ByFYLwXoctL0tP49132JKg
J1/XYlcmek6dzTGobGxhTU8MSCIF+L5LJc3AxVvkWA01bqeuy0LavFsuf7VnFAvE
O0IFasBwjRMQ9zmeVeUdRn4/rdVoaJxnTlY0MsCtIip3RmO7EeuEVaWriOzjNpJq
j2FLYOIk+n8yYcP+UyYoxFKdGwKAZ9t3j3goZbNS6DkCWIal3i53xCnzxuz8VlbV
B+4qgZKg8TFG9124eGzzwY8hUnR2awjkHX9vVjzfT2fzERQKqdBxpb1+tDwB4J9J
2Q46uIbikeGb/pzoA/VnJB1VjbMQO6kw926LpwdEUpGivoOuoOBwqVMpwQL4Fhfz
6EY/UpKc3xjvW8A+FX0WBS1AmV5dZeOQnydIHBptPxeTakyDpuqbNHvVj+ndPnwl
svRk+E99aW/I0mvIZhUlALUVjmMa65YtPBWxHplMjaJA0oOEiGYCnWXWRje3ZM9y
hDUCPTCh3/hBahuj0ox0lOdoBb4nn7NOEzXsTaJxmvNS/v+Vc/M7vaB7ZnqNXgz9
kn573BL7iN1rZ/Twj2kgY2exLrtjlO9FrQCvqRr0Pph6dRV+CLPv13XW4SMPtfWm
ivHskDnfM6v1dNDlD3zX+ApY9mBmIlbXr+SKL1s3GkcVCOtgw9W175rWPwaBJxvc
cDJuQCr1B/pTyVsXacmoJMo/lKUVj5zZcPkdKAUHqfqa4NB8RNm/rJpXVaTeUdS6
nOSMS2u9Ii4dUQFmcxkkiJCtQQOnh7ni1+avwlF2jP57Fb8ANx68CwiKLbVHgRz+
FTIcaUjG1MmYcL5B2Pl/W14b7HeuyxntswxLtVSx90/cEwxsI86y4yHtukmS2tYl
y8SXmc4OqK+roXOILC4TQCJuRf7lSB1MQW1kkKENWX5fqNAc2vid3XG1YUrVCd5i
5AeU6Et3/am+m4VejVkIn+DJxnacBsuupMbCE6EpU/wmglyJjqTTjhxCZM/rOcTM
3+oSwtcrzr5kb/3IVNuZJ/Rw7H4ZFh6TuvPx6s+lqZuA4v8nxTrEf7eqj4iith3u
YHHPiiwbPVwYtOqpvRvTQ4s+vt6FE61UTb4K0u5ookNcmt3nVpv2nqBHrs1cqP61
2mDuX8LObI72wY2mLreemZSSHJptfA2mWxTXcfGqF2L6PgGGnz8rApfi5kqFW1Wd
qUyCV9FYGhVDgpJX24umSLwcZ91qTxefjdaGXjzmhVd3pyUcsIkAxQis0yGhy5nO
LVpGeOxd5OQfNMKUHQ8wevCIiQMYfDLy4ONSs/DXDC2sWt9SbNLbD6IlDVczIzL7
BxZIj1cSfOyQOGBsQ8svnHhjtlZIAtcoRmEyXHiYkNL++URRkm0Bhd67e7701O31
t3vM3HOKIJ/IZQ6cijwXxNglLgSgq72E7HhVftAEZYcyZ+IhgGkltn9ftXfg4kPO
84m5xh6JEUxkKhCQLrFcYrIVYPzYhx0BRBvoGa/b5uoAq1VVpjYV+Impj0RcmGBd
UhAjo60laEBqnksSOV5r1ymPN65OqVm7gs1spbhTcb3Bh5zmkUMKOTcUR2VD1RYd
im0kBsoLAgcrFO9u91SxPoP4bD51dCnJ6Lv+KvWTYsUbMtHAbBd3QbzYW1i9tqyc
UKsBmqIkI0f7l5/3z2apnGUrTR4WNNTTUFWVKIW2DLwryiRAN/pzRI9i6Ry1nr+T
ouDrbS2ONVnlWHOl9v8u0/WvE/Dezwkpo4g9nty8fjD5MLvvBk1H3SDNFtZYRFMG
hPYhWGa9WGCqT20Kst2AARYAHcZMzTH3SJlxCbLKxXHv3BxvBhICbxcu1igNd2DT
HpEExajSs6o9SZmQGt7izPN7WrkMYq96kNL3g3bxixINlKp4zUrI6A88mXiMRJ79
YQ+SSFI8owIgr9dgZcbHOF2AAT7Z4M3Ivu4bCp4tZ108ZFuKKpKADxupw1WHqvug
UJKy3GJ1EpeLB15BpJLwuhz8mafrsdIK90mgvaxVNrjdzbTCh/fa5Z4a/2vXofQm
mawPqbj6EaYxCHMZqm4boNd2mC2WPAX+CbNKuOhFAWJgVBWEf7S+GhnEsXsO7VBF
1SxkSrkJuTPZBygp9lTRhRc/S2p5KROfXeH7HjP1arLJx355JuxvNtv7JMSvVO3k
HdAA+Rv2FrmZuWtGTO/vvxr9GhQeJa1NRbL3jBwVG39wdcnevv8tFmjoAR9cSS83
w6j67uz+M8ri96AA76tMBvJEoev+sqL21iJujB/iVlAzmwub/4A7MnQJ2xUpoS8p
YA497RRVGFkJG+OiHtp1C6Aoil6tXnDf6fJ1YZSUCcvDOZ1vEEQsbvvSPWPflS31
BAv9SsXTkxk7Lzt92UBIuDvW6OldJKoVrPd1yU+IEtu9F6VZOWR4IWkBrVjAGmck
baEbQeBx1kQImAD6bl37pAK0CMAknu17sDJow5Qj9kGX3oTd3ukS+JURoactWZEz
tuZE/myFbZu73yVMB+ZJ2jMzZSsBXgxsKWqxSv2BF6d7aWKtUENSkAg5suyso9Ml
Mbtgg70pfOvu+k+ORFh644wkQm+kzNvkAycDEGhSf0iN/CGu5Tkk82lPws1MHawJ
TAtIxF8+A7jYx0680DQZbFarnLSYfaGkMs54EmlUML/rzIROd7UNIIT8SalWKvxX
yj90RqS/A1fY/2j+wwXEBhkmCNG57HIdeY0otuMAEWTOSEp/RMvMdCNa/NvPlP6M
zC8IbOtrXXhUJLtvjJiYTK7WI6P4Gooc2uXNiv7VTVpzZ6/Yyq/v3CsfzifIxtwW
LsWo1mRY4ClUQO2MkxMtgq3DdoTexwr7co9/iMhniXEpwLoDYwdQ4PEyQp2ng4ut
STbsmbewrvngLkjxGL2l13W4AyyvTSDkx1e+fUXMexm6mv+T6Muqnb6SbQBMzmH1
tGgZ0CuoBeoSleewi14B62iNfwuWh6aSXzlkNqZ/uSSKdfsnvGheCDKQ3Faw2Xh6
21PDmDpT+e8kTK5OStoJ38EyjqQSYZ2PhYK6FLksVrFzDYhk8GE6Xx9G0gmgs9r7
AEXLn0jNq6TjEC4szHUibddvvWnFlkJzbGmC8I2disR6fGGPuJG1RuUFcvZv5oOD
iAoU9LQA2qMTsLUoxcSZPC4Rs8opxAOkjWVlrEsW1snzC7L3ESeUNPXlnhdY8BFJ
H0IKv+yXlJyhjlprtmGbKLOALX4N3I8tieurPvZd2u8Sx6m3ekiXjqRQ4xZgPcGU
Hib0QeGkDgUCNBQgNxYGg+I8uQ0UPetwxa7cnbedyTzjN9/wNGa2YvJXBWpVw0zG
g7UXzmPy5BbhApa0+zR07CHRKuVgULMv/ksye16wWIa0OKew+O4zMrNaxLgMmOSe
YzuGSn6zf4Lcmc1GBTIPnyvnVJsE/tQXFEAWPDYgiC4jY0XQH8WJuaUVVXHiMj2O
poih6McX3nhopgooFl1AtsWpe9zQr2Sm+6OV4K45sX4xy3AdymSoa495u6DvDvHL
m3liMeLc6EmuWREztBN9QtL8NtL1qNjMjUoc6R7WBPs+UgO/oW0FaRh3aU6fnW7g
8sbv2GOz7FSk8HfPzTYzW7BytlZNnLxYatOzRUqH9NcOeliE77AO2mBxk+dZgHkP
RWZfN+BhR8YTh1HyrKri8vKgM/vhY0+Ulmf6BXAAtlpgvEXrEvgBvYtpAiN2MMhw
wD0d/ik13JsB0ToxzI2+am3HA4s6h4hXuBysT6zrK9jHDFRJcoF/TnqCABSUA6/3
tznflUTbqWZff0LUD4B8W+tYhYIafFQA+r3KQp0wiUeXknIOVZC2wKzof2mpi2yd
BaB1j4omERbFh0lHMI6hY5U2VD57VKZc5U79XqK6McafRwlxM/ZXDagYu9NtgZ3x
7kmbBKkwxhuacVvRHBWs49AXqg+mdQ9a/dAR+EYN9KpsM3hA8bHNP7xAJHJxrQjs
BAp49NclPjNDM10VGHnBYUv+vAN9rFWw+wthAAc+dR0YcExyfE/E8qzARM0tl3if
lQRILJKCZdrGPkhuWoPoYQ7+YSP6ZWyuWVcArry2OVOwKlylcqN2Z7Dw83/nyj6C
/reQCm9p62N+ip9tx4/63zLl2Fgq8kiZUinPNxYhg9xnzKR/Em5ct0yoh4DZBCWN
WAQj6sM2Z7LOYVQYZFyczByLgVBa8GGsjCmr9kKYvwMXAbCowfZXw3y0ygVbesDp
ckUSl4gCJB17wkRSxjxwvWOwimdQH1w+kuRBcdEHtBxnMpoYKF739V5c4wCwsJUq
4jgvRzCydClkrqmqRzV0079oXNs6a2dEwWCuD2tqtVc4llmpfVHHf8BGWisyQ230
xO6cwTePqKdN4e0Fk+ddipfknJI0LqZHxC9z+me86hh+ej/Bla2zAMh4SF+sZMkn
RJygpa7HOBp2Uxi1iQJdG3upDA4onsJRwT1UNQxwRswosxC+1nD4yt0GXOFwQZvR
Qw3CIUfMx21cNQF8OFIQZOHtlhYAfH4SO2yJWkCvjGOc6gu1wzB2UgjuH/vUtYBc
t0kjuJVPmHVfp7McyIfFJQnhlCI2AlBBVvotDKy4ZhgLRaiOH6EhNqRgjKGVcASh
HKayiOguRpCFvWBqnFQgGZQyzWqZVMIILmR8fJy0+3bRz05GhVzcThlfYAvlbM3O
hrguefnJRmUJtbzvDtHZf1xxbpgfDJV5MLJnf3/4OUD8JiR+CcIrHZfiDB0W3TWd
LccgcickGTmNMxuIudUmAEFerG/s4xJdeeTxtbPeNFrVZ8BcRREXsxbGEhruEIxU
BuNPeG2/wGEHIdnlVMokqlj/FTe4BVDm2Z/QJZzDSgEzfCCk/NzkJDMCqpxIeHR0
f72CzQrh0lmITTmmjezPI3iT/m7bH+ZlGwmAJ5JWfM7W8Sx09kNtFdkUkSKYf4cr
FUIm0FHaL7u/Q/3IJXt3OKr0Gf/0gc0s8JwlUpTIPtRDOLrwAn2bl8swJnBD6hbm
+XZCWD4wmUUFDrJp9qxwlTIAp6cXeN5KWjOk0N7k9Wo/rjbweYGhaFt/o2t20NvL
QniU1u1eqU2jSYvnkVuL8mAZFNuQqadt+mF82dbG6/6PW/3W9XrurijaDaFvtm45
iW04h/T1YGu0tOAk9gLfiswLvd92aJgZLvYIlaMA2ElkiKKjsCH/grHHYn83jxSv
SuM9rBHfJ/b5yj/x9ZavN7gp6rsjwppjPY3sBSgAV4PTWl+9ystBZZEKK6MoT63l
jefOMbxNqqJMO6Y3LrssjWpKCe0AZBCzVaklq7VjvfWFivFnwILxAqE0/3s08b6w
EQHLloL0LIX+Yljr5QlmbP4UC+AJfOboyaf5J/JqP0lFDKl58gE5YWIU5DLvNIPb
I4yEMlPl1EtnGd/FeG37QN6U+GZbKAR9RAYNdPUm36iFKpXhuVVr/GiEyT6uRJvZ
SfgPRbXHrAutLyZo1q+rOiwe9ACCnMWipNsoRggs5ornpC1SVyn+OGNbx3Pqpn0L
NC8oxx9V176MMgskGSKjQ3rMrfxKC4+ZSs1iUIpfRPSU2tE+DgnASxIvQLSwffhB
xzXUbw1tttdd93JhI7FpVksfSRVj2PXg/ThZKYGffCfq+lf6pxPmwOJ2YBQjhzjA
TFEyDxqrSl0WsJmk//ffTCv4YgXFf+bsLhu/zBdN5lHc5tg+xPZJmMu4HobPQi4H
fFjrmffhSNwNnmkkje1zNW+KpW50YJ0I62PCeS5ffsf07ZS1abErk++93jK/mZL/
mbI6/9lViwl4H1hr2zyd1AG8pN7GsRvDinnl1uV2l/xJ9NOoG9eEOeYXEWGNr2DH
aep9G/mUrZYjaqkGhcZkMEXG6fxDVh7olV3bLgLYS0GlC4IYft89MWK7uU0Ctrsm
yjkrFK+tj8ob/A8eY8Xfg9zHM9CFd01ucB05CGsyyEWwqJmpM2sRHtKivm22nj96
DhkL6lCJqJMdmRpdlLFGyFoVMiEBtBYtKdvw+sZ9DGaT6akxBT++o2qQoQrhvAy0
Hipr/UscoUlkjX8QeEimKyrFP0WGLyjom8e05tBu/OSOTSRIxVlYC1sqN91Gar30
NPczB+C6n38IA8c4+Aiaz64DzWCa2y2KXrIGQkkdHttoBjwn8WUc3MFwVTF0Lw5n
98rJoOmk4cspHvjvyh1ZmRXxnZzZTvRK6ncrza5g8VljAa9Ai+W6UUYDgsjFS+cw
ZwUcOlGIRFzHGA7PmLzqcjvPYWoPftlaVlPrIp3FPqlB2w4qagZIAAbkkNI6vdlg
Zp+o0G5VyVB1Ng4Q0NiM2ZXsVHBXIIAVzoMJJV6Gh93Z4LtDlbyP/C7KOZVY526d
P8kT5JJYoqPnxN3krWfT6A4YbaCV1NKeMiiZ3+N9cQtT8t72VdFgYzMMXokAhOWi
MJtvWWdckLKUd0t5gqxycZUcxos9PEgABUDSP1k/ok+Xcg4XjTa0N7kZVZgTgYs/
/aib0aIyTjg1kZJ39KgOdYF9YxziF5U8bzYrCkFA1BOizcC3B+tz0I227c3sfBE1
UlKazc3MCL/Vqqn9xzHpbMnKcWbk7pYU0Wg1Kw+Fas+RRKLXl37A/lklk4YlqCqv
wzEdmZ01PbHEotFh9twHjcVL2U/k0OPzJDvWkiqNH3Ieh1vQ8Rf/wF7Kx+JNNVvc
+SiViwWsrktH98uAndNFMa/P4+9kV143jHaOBklYPe4iHzTtTgyHEW3LM2PIWE20
jng31FU8pEbx0rX9YWxwiZUB5skvKq0MTXDJaGs8D96avr0uDon1W+xQhZnTV/Fe
Hb2Ztef7LuGhUT9yXqwcbfgsgsk1bXK57pt248S4/7JTVqpIoNTb4F/Gw/CBQGJ0
t4WrIuH7Ul0DxWKq81u/vtKgfMnOmXjSmtUwQnZmlzX5Xs/1UPN0gMbGTDhu3xVy
I9WoyuXXdazPlBoJGIp04Rvmq+qfLZ/0ZHqSuBwboGfKRynLQh6QHs9mP0FX+ok+
w7gwlpbU/+7CjuwloARn/mbCbIrCyuCCx6URApHx3668F8J9/p/tEjjbMEa7jnSl
n0LMhdszpz5oPoUrZ9rsOtBb9+DuTcUD8AUhe0BdsG7gHtdjkc6sLfkbKaVO1q13
/GlqR/e5a0yp5+URxhgKMB+9c7M8QrpwYnYzBxrS+UNT6Woj97kuy37tkeZPuzkh
4iz2KHzMePNMDADfJ8vH6q7RXlRF0LoY1HGw002KMstARsWm++mf+QyL+lZ4ns3b
QzoVRKrD6etov3WRSiQHQSRUUWXIo4rDfUdGDqvIUufBWildho1E4mbB1Hf/ellE
+SlKv02PaUEtVVRKVDbkYuL12R5zrPIRsgoLIQpeAmggbvNWd8w8Pi0eLKpekvXo
U/L1GTsplKWMsZFv7w8yBFI4JCd/GxGYvDqwAsFgwsN3HAkMi3MjaYA0A8zB3YzW
EnFUF52vpxmCLHYSAKzJrXBFldSEDlX5nbizQy0JPm2i8DayKS+8BmmuOXhgEwbT
WgAsbF4ycqdot3Zwhhll+stg63CLNOD94ahbRHeiPlqo8IX32Thd8altm3fK0Je7
//DydfOUGqCVZLM/YKTlK+yRm8ql4zj/EsaLp54QR266gy5FC/iDydSigIumQa4P
1T04de7dpMKOMUFxhEEH5kxMX/LUD7TlGXXQfS7BYfsUppiS8ozyUZN0YE6s1m5Z
FIAQHmYnA1ToATzkea0Cpa94uYfADHnMPYK8/0GRJ/e/ccmWXYczOBZv80nN07bl
CJUtcLFyCSQaKPHr7hdHWFGFahXEFuwufeiOrN7WbB2ApnfX+a5JqANTL1XUO2fA
HFJaXOYmxuEHu6/YqQhhxGwL8eDClJONSQ3IOUYR5kSm1QSzffUWLQVl1ySQsiAC
9aWCHf5uSlUee+WvUYaXrMwXehRVLMOvPOSHQg/4r9r0ISDscaTy6/2j0FcvIEl9
I4MPCt0vM7mbixZ0CnFlwZRHjjzbowCS+eH1WAPK896IlS7FPR9X5gKXGiPC2xth
puz2PtiCOAJxutet/pkRh/yEbwwcFNhHWyg1Qd5TPWn7HxGxnSLgbNIYzEORiUlw
f4WJQeksv8fA7GLHFUgjG1kalqE8Y8qMA/lAfigsKUwx52Qfd3yNAwhZBeVk46mX
Pzq+BTVRKMlYBtPp1hxOvSBNJleJV4qe63JwmdXh5wnI4JASpS4K3lOx6Lj2qLx+
NIsjodqg+DShCbqkmrSuAjAX13BkrJ5TAO/fGscvaDesrTntrnp/0T8B9JNLRmoq
Q9zW6EyTCGp71Bcu4yQup3AT+nvJojNaXHluwvgZ+R+X/oJfHURkOT/6Ud1P15c6
tLu1aOog/CKUl4u5UUs7ws/0XCaBMldHMKmtx9FD1hkTnu05OHjVFYtxyzey+Lte
JWLSGgIgOLOnEBYAlLyw961bJrVuMjR/SL4uo2Yo+9qDvCwPcqLSQyxHOLzt5ObS
9uYSEZSi11wOrgpv4YOqcL0Ka0Sa+rDUym4rFgzqO4KQkTdfeQKgT/SyAb7HNZjR
TWNdZfu143bbs5tZ7kThWd0eWUJmt0q8efo56Ox3ummL70UtlsLDFV04Rh/sFEJw
enCEzcttU4+N28JDE9w0lG2IEUTeir91xj26hTd8UVe6lR/9ru4obCusKJ3qyHL3
pLCwg5Yr2yT4ofYD8x7F0jhYFUV9JsV4DtaC9lxq3YDTGeDPqZd21qo/m4SxAF4o
ndY2rkbE/0HLpgg6S+UBpEGbS+jHazFS4URnE+z0NqUgwgF4uKgKTJoQsueFRbD3
JMFEQ2fJ73/dMIKqFPksCFg+BeNU/vGrBh+E4U3rpyIc23wQc4wC9DILApzoqsdM
FoMaglyut+W6G+xDFim9uHR4GvqNBbIq8S/QCzMSyabmPJHUKbhchy1SV6yLCU4j
AQEQIeeyaQDtYjaPN7BMAEu2/S4CLAP0DzytkSIwGpvbo7t/nXEfBqPEJf8Pqvha
SeqvE++YIgSmA6QiDUJd5ix4FkJsI3D2TXsKRt7RrbJx6HLzxpOmZHlLOrIEjByn
Ah6xK63YEN7u5DnioomtQsJWTvXf/ptQ8NKu7dpL9/PhgNwm9bt4cQ7nxvokXlJU
0tGYghSuVBKTPA5+wHLOpCztgnY11AHRFdDShrAY1XQKaN4VztUJ839N9JHEx88N
MicVCljDapJxA8op3w66l2WNVvwq1X8VbJX4fjcjGiy/xZgXanGfGm4e1DzV3epr
N9RGk+PS94DHI5oIxbRDG25Eh0j38m9xtG50hLKFjlxIS0LJ29zogAVYtIQG5y8+
Vjsn+O7TRtxhjsJATEdot8DUXsdCWnYbMC7zUeRQopUWT/Zw/ZdLwrkz6Kji2/UB
x1zBs94ok3yszO9tXf4xlYF8Ly/eiYqXV9pIV7V6BG/tmrnwLcJ7CJ9M6KcXE8+f
kZ71Pc4mxRZP8H1+r+Cjs42ftDhLKZkVKOqDqHKftwaf9tqPGdqTa9hS6g5DIlau
Vg32E4kVw1IS2rpY0bXm8XOsB0hZypqe6B5tSMb8+j5bDVBUzWLodJnL4V7ri4Vh
srtoVVzVhLgQ1vkQwRTo2ano2uX75fwzTc1pQwNYqUStbzyzrpNGH1UE+k156+Hs
+3H2CiW31mgwh7C5iE66EdDyLltup8PqKaT7oo5nntwBaklxAe0xMKMWglohosRq
OHigblOylra5m6Z7cWUF763mFAEgJJB+WVnjtDYER3pEpIXMzcc9CgeImfFSbXIQ
HZccfJMa1TsivVvm7ExIS0b2pEbmj67rhIboowIwJsS2/fnZIoytJ3vlnQV7siv8
yRkIzKeFgyv7Py0Ngs7OUIwq6o6DdVNPeggiBm/sqgKEip7WoCIIDMR6Ovk2EKuI
iTeFFhJDPMnY35u5xNSOJP7tehcwOkZAUwq5iVtuJ4g+5RI+Z8E+JAl1GPmzT975
47GSpty4L+sLPpnTcl6MFZRqEqgWGPtJcVsxcFRfp5lCZY4FaCZE5rKVbi919SZ5
nE0frf02Yz7/xdRnMSJWHosN7Pv7VO+odY9vZnb+iOxqO1DHZDI2DYGpyybyoIiP
aFiCOFYBLFAMIjfuPJG6NhK7sbxaNnXZtFlxrjCKbm3gookCvoOa9AvnwZPA/p1g
auI8EsDzZqxRes3vYKRJD6O2Tdigot4eIGBOE/j+jbaQ+pKFc25p3oIFE++O/t7w
qhi6ZbYOgBPxm4pICrwentGFxwEimt7Tcu/VZoDoXNtbhTTuuKw+2036M3XF174D
jIGNm6Tl864x61fIGpdRvMkvuWG3flkm7UkZOhHYN8qfADkiKKKQevX0AH8Y4L1K
jfTwbydS1q4gQ67mjDEZJWLCatNBExk5f9r3qW81owBT49pYjfEAWnfgRg/Cnszq
gBfCc5Y6fd3T1zJQlrTrOYjTEbr6YoqOibWiuOO6il2Qi+cAqLkGXe6wzNNAh4bd
W6eX0ojq0CsaETkc6o0B+t1Rsh09/7XPhH9jevTcxA5dLRvA3RKIr77BKucvjkh4
3gw2bx8k9FNz/h40orHrLJeV/frKP41VWbn1LCTn1gIa7lewpNKwrBIHc27h+rBh
uyrq+sX1lCS2EtGRB77UpbNV3InzRU8q1Y1tqvotJ9zmLQyXKzYJtdOpNy50nSrr
hDWNWs+/+3GULEz0pLOzCqJyJSceclTpdQLRdvsobRlEWFTcPTR8m7TJs9qIvdHu
fiHSSOD7+vMzx9y92o35fKv+MhcWwotVUwfxwkRIZKb2UFOAknd3HRWOno8V8eMx
DWSVCBMMz2g1Yzsx/ASaF63EzxJm1ZMxbZIItY58lhuew/7IUj/Y4OJV3Ko2wT1e
KjQ6WJEmuQZrfbHfYKnFCvWicrCNdNEsAPDTFHwz/bv9g1u+JwYTFtsLEuAdhM8S
0dDYWpni5fXLQnAxAab5g/zq1L+bUH0iLhf1kNLhJ/t57P2T7/vf62bL3L9PP5hH
4In38G+ZL09h7NvTJBh3Sph2iwUsohXovLQFuKXB5krMlj9k1XsmH8t46IArnjw3
7n/i3eM2Hwdvy/bg2u63PKHnvbaNvGMc5AqL2ILTQ8HAsE8ysu6u8mHeQAme135u
8oWfazIJWnIpK6LffkOQOxb2dehX48beBIFWZIN4mkuSH+/KQdBdQoIchvXn37mn
hQ5bpMsNsCxq074rQJSt0HZLqvVdeX5gmjiRqrvWTVjyupir88gHpgbwgn0IHcLN
fUKfIv7ftFTEtwoKzL+ZZ1FACui8XAR1fpHOFjpxCyJFEXEsPTKtjInRId/RgtHO
AI8ao4toY/DzAsjlh8dVPrlHbz0W8aDNkUYFG1gYdm1Os2i1aSwJze4oSU3mbkWF
7/wF6WHphR7MiI2Z2QEmmCzn3OFgfzz+kRYMFQz22bG3fGDJteNfpp3I1bzumBuQ
8vSgd5My56uLruCwrBCTKWi7QlKwzq0yqFgv280aaarEZJlTpLM/TA/lq46VK/m/
v7ktLbObSA7HPPanU94RRPgTh7hVBevnGZ7zi9ZDHa4UKepk7NA7y3cNuw8c7Nfc
AbEfxoerVUZspqTxlMrPscz1Q6J1cauIWvJoUCm1mEU2KYxARicaFxtq1lWiWooR
i/W9h4kR9tFCw17n7JQovi+ejV/obTH8FRGmOoBHYZi51WjWB3pG58/ld2W8A7F8
ImyeKe9gVLWd1w1ACibI7XQ8c3liV2K9OQ/U2JdGXkX2FSDIM7zH2V7y5AtIQRQ/
lFSA1XGgLPJrw7mzB+cDNuanB4BBn+N61z6kgjVdcUZhLRLf6U1cvQ7Q1RKSSmmd
KinkKCWLlJJQKYgxphaYgLZf9BAs9eEahbmW2i2lcEuC5Wr3IqLlhKLHQUPG2KQw
iLD7ZJJGQjzwnIN4oFVzwt0c/5KhfmoYNeNAV4IDd/b2xocTmhj18QDu4VzCaeXI
qAlv9/ZjzoprpoXhmyJVCJNWalmbjInZ3xSAvoC2C44TPaeXjU4qJX+uFphTyGSd
Wq7PApnoCb3KOku8CWKX2It3nrtrjdSA+Ap2j9nHcpr8z7L+4NmqJDpjF1OijlJv
doCtPLg+FLYvBbvjzcxjkzWifpL8WzwRLiQ+2Npo32FyZ/1OfTyT6WFWzRlEVnMO
TW506t8myLT0zuTord+xf+2SD+jcu7vJ5Ro0KTaKUipxUUU0bnJYTYKo6leFgfaB
CU9lrdnWCZi6u8jr3fXP6UHCyyCb5DZrKKZOyhnRV0FeRD/5jF9d38Hp9bccXiqZ
5bupi3dMUyPvQKH6dCQfICxuzW7LncByuzcO6CztKpJq6Gt70+bXRutN9dNn4CEG
6fJgEwSywbuWbZ4VBqa3GOgksdvwCiF8i766SFSn587c13b29XgTzRbkfiYYTy77
FhNwOBSJE4Kl3yPiar10npa6/u9DudTGtAtfqOKzeRPlNcM8qXGyCih3ZLGzSFC/
7jtSOBnVABwp+Txplw8fbKddq3IFDmE6cAG4XmrrZv5NQcbzifw2nEpIy+/pBjSp
enn2fPSqjVcbPSjtnUr8qXFrmrKfH6DQGU7pByA85ij6TYK94yw/mMt/OG2XsrtI
PuULFlgFvxHzMiDfxEg/nJLDjrXhN/xzyrlUi5c18oPO4Flkr0Kgy/Wxxa0/xzWH
LfbkKNuPJqEgRyMhjIVPzPksJQ+SsOhN7XY8vBzn3yrfOj0KN4tYu/ENmMcYOHfX
h4nm459uNWMrWtefEiatZmkI74FihwJumtW/nwzrMn3+Ut7hgxZRoh7sc4oz55tV
GAixcZ5oh129gnT9nT5sC6F93NctJFsZ6fAjP7+Fr8mRFG40DPnZvhG7/OYgSQKo
8FmiMKt/jS3cPn/mVP+aLf7TFxHP736/aKZkG7AMOmfn/G0I1WqW5zTs1F9r/vE8
4cQpb5EVp6oxbmh4eaUeyZCU3hSu5vqHbxK5Jpj9Hk+XACEE+HXIBcV9FZlweDyp
fAOX4/4VFL7gtIJwi62yNnXu4L81zbvNgDw6TrP0VazaAk9qvxY3CSCyOYiygb27
JDM1963tS0E1q7tZ0vZxVYa9pPrqiFjuZW+T4dN3DfVNNEqBCSSV+gOPhV7utrcy
MMTjo1RUPAd5mduoArVm1YL84FqpCK5PJ6ihWzP6urfyLkFahB7XjW8UvOMuHImW
hZZCZCA9Ieu12+vTF/1SaHkPKikz5/jL+c0LF099DppBSgLZmqUKsJEG06haB0Ol
RUz4vEnyzyps+CXeC964s3SSEy7TQ5Np82LtIDExD4EK4WqvH/0bOA8AwVFpdtJi
EDSawsu1UJbXLFJQUhfxQBAWQab3EQlnmyhRAp951fjMvkXsNv+/PFDmMB6aXzkj
17GqPyujyN80lCACL+kre3G116aPy2T/rsN+Log0aT2FvfWI4HZAsWA92RAUc4TG
Pr08IWSo6TSKLvaQ2EeZcNfxufPZr+uHDua/OnSZAy9ewW9daShBVS+uMmc+7vYs
Yocq0e+O1WBCjpLxRJziYYdmMDNZkn79+yWhdLgNYMmye7JHVLSOUg3dt9CmHLqI
HnKxMCtQy8b3NyU6BrHfW7sKURCCY0917uKz9JIrUzc1YHDX6NCP1o9xMPdGKzyH
osqA7yzoeG34MqSb+KrbUE8TDBbq1sR26SZDHBR5ncv9TnPNaksKOGARfktLNNyS
/gECzxxTrI1pzQahg8+2CFRAlkjZtg/YxR6XdGQxMWFxt+qW3b8xyDnuBwZoMgNt
A6BpiM00PkYEXDqsnpXbU9Fn95zUxxgBohYGWvMS/izYBlh3UtWaWd7zanjhjc1x
4qrbJxiaZW0UeM5Q78XPtHlMlfEPiFhrIqE4x76Dt0sz+2qlgKLqu9JqWZ1lXPrZ
goDkpynlZzLHKBlhJ6m7jmOyzfToEmHQwAkyt0jtIJ3vf0efamkcMgcNG0lUzAly
VV/vKMyHpns3kmS7SXKG3zT7kl1ZB3kELXMpE829IlBo9nIsaVd8xteEEg3KeD+p
AXOO6Gosk2cZZUEFhFsFErox8lf9fPMneXJlpEBZ0FUZGuuELmtJ3FmRuVSeshAE
nkrHfp+DNCB3u8SsBJmnCyB/v4guVjkaqR8U7ecLaBVkt1RNwd/PTGm6YiP/lwpP
N0fnsfunDsJY8ZRym5HT1PGmJ1LHSddmZ7Um6iL2eds0s/WDzgjuHKS+n4jowhNm
eKMqt0mueMRTCkAKP9X4BrTOEUM/GBKPD/7jGmg/Ze63imygCvRqgPD7VEdC64BD
68yKI+JP6cPX6NJdLNLvlDxDrmWZHUJA6VAHioJ3k77r65G+0veV3B11HDQhttxV
yduMYbRbw0HfovgdKhcydPoxQ/8cPiB8tVfA/zxuqMhUthWt84BUqH7SpUNNpncf
L+ntLuHgqNYydmHGpKjkygkmnS8PrJZQYQ3ZZRuYAR6msXEGWCoRl5YdS9H67Lwm
WphIkupi2FkLQbuWlCwooNjXilvmOTJM6BMlPkRlKZvAFnszKsi2fkGCO03R8y90
ByV7d5G01GPGJLZX+XimQkWdlfDC7iDO3oN02w8WEVNar9DsK4Dui0ojHHW6B5NB
jGDzoEEKp068I0TGCO82OeR1FCXVKimXV48iIEVAN3orVaI/K6OdHaqcb3xOHy0L
/q7j6fy1fpS2qB0h9xdz938poDFc4bbg5qdMI04N28j7cdfMduh2uZZA1V8IGSNG
s6VNZcC1B891xJ0QDfrDFKhrHBGHO/XyUz7zWMXBk2fCgjl+Yru2KyrdghIXtwQQ
Oa4Lu/2jRWpsCC7ozcU65Twdk842r/6Fc336Tc4s0Nm0dEgo17b4fQPJkrD8cD47
RD1AkZwbcpNaBjQKVnJm9BQLGrnPsM5KehEQpEKJoWOfVTqklXuZjIvnbeLGN3MG
bV9mIBbRofMWc5iB728XTBITTxejtlr1tFumsII0HrAQP2RF7Zr6vcbk7WsbimTA
VphRoEo+fZVtkyNa2iRf5rqYdZyyBod7tn76oaW2V8J5Onpmjw41+yTxjdeMV3Ay
FN0JucoohpcWB/yz6ozp4nXhTiqeEyODY+mCz2I7lV/eQ6T2DdTzT5xqHaG/M4km
6mn6dvcmHEXPCqpjZNZ7iU08Po11qVUST/s02TndxlGnoims6nB0t/oClWPwfJQb
KCO9xJ/f5dXJOdDcyiFbnHrdnS41NnHuy3lhmkjj+0A4eZIQD7gaXpfVUqg6YFNr
amNUWZxd26uGOZXPH6xHYw8HdDCq2mWeNPYd7a/feggxW1YdtiBACwP32LZAb11k
3yznXY7uWx6FunMACofm7PktPgSFgGjduoZ6tJGvsiVYUtG4Ig2T04IySvcX8Num
1aAWEwvJsEUA7AGfUA9j6ihzt2P6lrK1iFy2dKajBB9lcliY5uwEcnWNZQSCIpks
cXYKT48aCiqlIRtrZluQROu705qVClx2YOYPVYEI2MubmXMhii2dqtq6BBQ2q2cB
hHsulfzkELy8CkQtDcpXcatey17avt1ZX1s5xsQDDfqsIlyk1UqZqyLi288cNmoh
baVEX5mKe3V2VliLlq9YJjG5ONqzHEqP8irV/fR5zYldEO7E38xGb59siN+4JsMj
zfa6dj5jj+bUMBolQXaBG5BV9IJzsRJM39qDzovqYTHA/hYeugdoToWZbbA9qJf3
s1lBpNWrnFL6Thrmfrw+P44ap3GcZVUclDo5l+5g2y5s8grZucNqJ5v4qNZGTw7t
ZNtX8JHuiwUBr1uHBSZnH+/R/kgo040Tca0KOF664DIEVkc5jicsaRIUGv2Lvhgd
zI25KxDjZGF4ZAH2VmOrZRR4a1CW4zpDlgpb3d2TZr+hMGEJQkitmz3dhvGKa85m
iDNocKWJHgnm+s6UeE+1YTKoY8QIDSbrhNVRHe8d3eqBZ+kvVkof8cuYtu829ucz
FPrqbSrMCLTXcPEHoe6oV65IcaLoJ+4SZqQQzbngPexUaK8evfnpaD6qEaGFypJj
GwhJeK6el6w1m6l7JjubAgbSm5z3m20jn9GFFF0xKHQlp34NJg4Xn7HfCXNiZffU
8c6uVoNRYUWrQZHY6BIgxY/M6VNGtITF6vvFSlZZqTNuI9VFYXGHjb8TXCTgueyQ
bjsSr97qeDC17YFbvuzFHDlEsjtYu7+wZ6zQoSw1NmLlZKkMm42X5D+4s5nIHm6F
OtUmXqDAEWHi7tQw9YS2tR3qnSBTJCZ+ROLZeLiWt9xH/T0Tt1ltpZ+xvlHFVSEd
bF4eBsB4V/VbONObZ/s60XYapUjGHoEoiUuXIxA2N+s7ySfig+w2uMOjpGIEwnd6
o4caYgxVRBmDXsNYtvcOWwk9wMoQnnnjHWwWZwMTPFK1WoL1UW7dwaLF0cg47CID
yWwyi9/QKgab4Jo0XJbuVag11f+ee702bYLG+OVJsf7PFoMJ6Wq6OfL1mOmNbgjR
jljUM3xXXvGzDuyLYdmCVR8XkPpG5AcuUBW6FBoOTyivTllYpkbugr0uE379O9nQ
i8b4TLw9VkeYwZV50NeUBI3qtxPTQOxRSC7b6S+sw2kozqxKh2mIPSscfEpIgfm9
xJNHTQoIuCXzbd3VBkCTUiUnYuiMatYlX6GgTiSGUkqSGc/Zj9+lpRmlgdm1NpKW
t9HG84mQvMAewBOMrrd+NiG1w2n/rtY5JKAnGnIsPaXv+D97Wy0gSiSPmkITbbka
2udzDTgge09M4Rlrxg/eE7Y3IA5gWp/s1NyOrfwvw14QIMJzQumtYaAYfIw3Jgq1
zDsmtoor3dL1p1iTafYuPclV7W7tAwFvz7ibQFVvO/uYKZqmGyGq6AoOEG0sfnTy
3fShqAnknj+PO8HjKCthMiFHZ2ybOo+AvJKDzTsEp7g/LFOc4mz2Lep5ogVLtAo+
R6m+4yZEsalQwiZxoYraGyOmfHWiQJBQEjv53QYLAepF4+JXOPFa7SfVlzkXXNlG
Xgk32EIn/zr4sRdquoEqxpk8RdipD+RJtEGheJS0/JA5Zy2uNvsQe9OulUb3k1km
ddAAd64n7cri0pO9Z6gn7XdpkvfHTJ/68xmUuJH5LzkUO6AMgXRSLGtYCIXWIKVJ
X+u+VTyvJZqzd/9OPFECrJEDHMHv+9Gr/SRtiOCPTpTkTYOV8oCj3f0iPw6fPBO0
uPv3aHIBa046H/gTgmLjloi2B+KZdOxf3fu3XSUo5cDBUBmiDiMlFzg2ffpxXXrt
kANa+CGwEAeWo1ue0ebJ8YEgl3qiTaunrZvQNhS1+KgfOPuIjYH7xA1KA30yIgxE
jjnudVvOGFMzkLwhKNxjanYSkgfpkc1DUANRnl6N+0pzQ0QyCL6myCvFjCgi9teW
6Wk9zpoZxXQK3iW3A5mVrB/jcWcgj1bxodtNGJMlZTGKNKbAYLqyuHVfeHIOUrXc
EvGDoII/wp7MPx55fbaH5qHRfw3wIzvVT0JuxtXTpIZWVzvyWFIbXCKkDV8uEQmo
47EomkRIk5HfaXSPeXFXW8M+vZEU9nuW81vhD1NgtMC8/IJlWLNSLhzN26Jen54v
hYA9b340J8vl/4hBBY+Pr/to83IwW6HRDy5fvia8pwWRM+Afm2S94T85QojigkhS
5HmsJmfVy76HWDl7vZcGLyTRe2PI68oYm41fHxAQtOwuQhI7330fwFWRrpWWFWFk
ggmX93lMh7X9FKLzZlNexpw4JVPKa6XSxajvf0pRJ4APci1mhnne/KEqgWRbAgRs
wiqjjzoE480KK1/rZWuLtnKvGUuuAb5b+lOiP7toIJMJwGtdnwutjn3nkeeV5+HC
U1jgBKWktcs9okofbvA4CZ4qUkYBroSrcMtfm077qvrnThrsxqyH4nL0TNYslw0M
Iy13wFKk59hDV4x3y9Kn8+BVLitd/nyKT3bKArRCLSTvlT3WmKM1LlCiaXhZ3trl
4iAmDruzIvLAwdcMLC66jTYfGhJAvJE7TwZfgEheUQ2t4sVt8E8ZJwWBWyq7sfKZ
FPt6xW7SN20jLQhj4dMJa5wPfP9qqpq+TZCgcdNwWGL2UpmuGTzZNy0M3gVENGl8
KhZI92/kASdmDAsSGuGwzFiRKvPwsuFY5EThsxclCpMvDlAHZqnX7IrWn2ZS/Msq
iEvhqybezXo8QYGqfBAidtjqtjAjamIO+fI+dt7RG0qkAki/1MRNP1eUniaRr+Pd
uszMXF9GdbRi6KNtyx3tsit+FsRCBH+ykeagJovLOKZzJ7G04iHubXOyFkOubbfs
cXxd8qS+YbmIHX6NeN+Tpxwx70JbcbtUq4WKTEWPOY4pt0HIqX6A0P4H2KJr087Y
h9eZbN+LLPLGZLHLFj1T1Gw3hNqH8JwvR33JMccWPkyNGthK6sqAbkMl8Q0BHuc0
BFgri5+qlrpJK+IIdQr8GFGoaWnfw48ixPkkMZThXwvUYHzRRWUCuqx9JnXAo1zD
2RrVhINDliyDiCB4LwsX5GWUt08cAUHkEzdZmk9ZgZp6xzIw3JGPX6tNAc9uK6DD
GuJTLIy4lAMOvLyN8ROagZkjJg6nlUoIL8v9aKmRdIlZHTZpxJj1EJUwuXirim0d
xujabRvFG5g9QPoWhLgAxRY72JCOKdspXtjtc7pc1GnvDga7+ajcEjW2ZGG0ewwn
BjBDKjGU9gf6lxku/Od26yNJ4EwwNAva5ChBFkkiuRcI3tYTl1L8IqI21bq3ppfB
eQrvI/qoGWixQZNgj6gHBH78TZVsrM/WTdv2+XBG9Pwubemr8MWyC1spXjr0OfFU
uHWIqkwUQLQw+A0ak6W4tKYuXoLpcbDAQQeYvz+KZvkG+tnKrZA4bwQ0RupvdtT4
2Php9ecbbjiYDN5lM36ZrrqojZCdYDnbzkaX4kkXUV0kgxRDn6Et+bdf7Y5XvxeV
PMsxnG7WpajPyTeyX245CT0nGNx0f38ZI5oBXqFzY3mniUYIGafb2/UIxC9+6jJ9
qWqya6InQMxyKxBpupL7TAD+SYwMdGGFrCDRJTW/4Bb+wEFJzmv/8i5hstwKbKhl
RRwxNcWpbNt0HgE6XbApHD+y4g7UmDDWW42yyMFQRhlZC66NUa6Kbw3oLARs7+yV
CaOt3TEfBcoFQo51CmFzuJsZ+O/aQwNPmAG/Rw/zxvmJHc3mxuIAH90xCcDRmv0F
LWJXrJvLHOGnim75rX/SJ3+WFTlqoBvaBsjkZcTJBIDVUowrz1a6qyx2xewzSYSH
f5F3/DvcgL71J+DgaDsk6FVEbsMnPqrlTJ+gtAC1W8TzMpnmVXIQ62gN2KnsgAXP
LnJiqFOvaplVNfwYx/nGSlOJr0mXFAf1fnsXusMqh6n5/sJcSUJkl38cD61lMgfJ
Yumi0aBGkHB0djXL06nNEj4qMGW0Wt8IZwcy5cm2JEh2ETkRdsfFm3wTnZgA/gMU
BEtKwwMF6TKpif5o+AOgTi1aZmZHdFrNGMxw0+lAhor4J3LDcuISe3/iUjKutrHU
Wpo3XRC3+vL7jHE3JvGmbWZ+aENk8PP8wgXChLwDx9ThjPEOct7gBd5c88NPhgFU
4cfgZ88zzfl+xBJ4OQCFhfYST5pCn4N8/ec5s37CZoReXKElN22ruwNwtfrv/h6c
Tngs78npbZYnUZqFTlHGGa0COwZnkjOiKnG5ULMg5dhuATaGWHFLbpknAiW7NJe9
bNjXhZSgznPuXXtikvOVOcCzpAicmaQoYo+vc0oHHKaAgHMfHjeM868k3a9Jxh4v
R/GgFNorW+QNY/Al1AAzyCDcTAnPn1xmLoGV9URo+TB/kV0m110yG2a6h5lT2B3o
b6SG8ANwcI/fSRCB22nLFE5pDs/JsvhDWAXE/K8zOsm3Nrnu0fGGoGR5fnQQdds6
EVa89aUaNrHV84EKz3KZwBRhvMQq1+UdB7wIh3XZzFH/dT+spsLJ/TI01aqsOqPz
nImNVfMvQqt/n9iOs3Sec+xwZH0KdOaXGGc4T7s3SRTPQqK5n9ImKq4kNHpeMKt2
sfmiCfi6Wv1OBtx9TOZKkA/gC0Dg8z+2OMq6UCSBBWrXorU6NydtASd77otTnCfg
V7w8Z7k2h51EI6YBQFFbbNAxQKN5sNTZQQu3a5LYUK2QtBOhl72qtrdX0a9g7DVy
dwdnY8xosZkXVIx8iOEvRYVYLywgjMCWG+QaP99S4i5mrsfm8mwOdUE/fFWGBU3K
yoeubSZgULZhcx90sGi9aIgejb+FIlezFU37tpsRrC8S8f1dEaNTN9Z2aacXmso0
+BQw3M7DvMadCbGXZ8M2Xd+AKkCvmaUZEz7pFtMPocZK0iJ5ukMUUtisSXm2PTmD
d44TSj2Md06I+QjQcurT82Si8nYPr+ZoeYz+nfJiFUMhRsVuWN+/B/mhebVeaD3+
Cs4O3hztKY2EtXaAb+tDJCnbOA8LCyD+Kx5u+l9DNt00+2a64OkhjFa53OxNP2XZ
VZhA4j6gylYqPzJg62iyRlQp14/aWL8k7rKBsTLB3/pbv1b+TGnUTx9AocFrLnvk
y8LTjl2yBEWmeOYD9LyGAcVGmUPbJJLgKlrxdKVG/NSTGhIVUv3Cf5LzxR5a63vD
ftBLBHBZkTLkq7NEqYMFveImgfK8z4IjtoEQzY4kqGTGCCvmKjS+96ZI8Ex0K0d4
iasnsn+MPh0baZhIbBiobAhdJWVn11rELLkJ/91sDuTb8/LON9wyzMUueEKaQG1j
PGwpwpq84rqUdenDfL1NfBqqzRtoGlrg3Y6RvV/SC+vi9x9EbQRFD6I1Xl8R6Sf7
xQ78JS0owpMQ2PZzVWP75kS/qIg0AIoJkAcpxZrfPScjT12LtIjf2ZVY3hQXRpeE
A+/d7NV77+XL2s+Q/4zdwrP1poLgeUnIY+MxhiOr2hixlURMKr4mOrdxh7/jysx9
j5i4KXPhXlrnWllZbyMJwRSdIUVz8wr2XEDfCyU8+b4H2wBvV1kmMfeQr9umvGUu
JUdNTitcq0EK7WUWFjMtCvdOPb8QcLKDIv6aTEM0cIAeMazv2/Fm6VNdz0QlP9eQ
63UD20fetCaiK63A22uWL+M1SyhdYvWJGCElFtqUmzpftGfPAchIrdlL/pKG7u7n
gmOUgabqicCjD284UbTyU79kexe/8ZcV/f3x+Ebq3Nrz4rUBuL+Gobx7NAgtq759
w+mwlNHsSsc8WGyom/SS6CifLTa9OCPzbfPddbX6g1HxrAYsX3gDzsngbGoIEqEw
jjgb4cbRInigzihfvgE9xRPxsTfIud982h4OaExQ80bIUCnhOYCGeU2t/BQjKLLZ
dd16BZkWngY4QtTmNL8XtI7AjPlBdc/Uh1MqOpDhDaJ6n7VnrBrNfTYzkLsnP1hQ
789xhcy+PSk4M/Eus18Q/1pLzqFQj3eOTLQT9wRGuAh7NeqI/dpXYBJAmeqJTnGT
GlEqvu4HfYgZ8WdrV1HGukeCjs9Zc+E/KtAws8WpSs0RQo2RSIe3pKJp/y4jEDvr
KYlhqZF8R92YB2NIqBG+8Jf+k0mD14YzqcsLiMN2X74HLgNdsi1jSU8yTH9eb9p9
J9oO1TXfaU5i/kI7VbOUyJCloVwWW0WpZ8ZBhCARHrWg8XULItLh/B2zdpN4iMAq
hJq9yZ2uPxUUOlkiZtIzJPe8K+THkMVNm9HCP0Ger+21NzTwdBE+FpBpC8KszRTN
71BYeA4iOktcYXrQrsdrUkz5TBFzkM2vHIawXJ3zAh80mERZKMzA6WACoz5HmpH9
Ys6X2S8XB/hRoFaDiVa0fqUAegtn5HGAzTyteaG9SF5q5D+E7AQ5YaOIfesfIo1e
Sum+PlYqQTMhU8AKR6mNqgZbQFqrfo/2RAFikHwAEWQu77R3HudYpJnAb6trOTtZ
a/T7UP8MkpkZ0WMQCHzBiXogN0ltFdmItJD8/k9J+ve2yEOvAkF+sUjMWC4iHram
q2OkyT/4Rs9tumm/2cOGFhdNUob0XfmBwOp7oFoePMd6qRL95yt7zVI27rDnEPsV
ROYYgq2b0F8cYatvNT8G8QQRGFAoyyg1PmpjW+1Wq+WMJJ5C/4Fh3k87dlFjlwJO
VDwI5aW7l0kPVOene2pTYvDkHN0vVfXMlHUh9X4YkrCz3ZiSrxrVzv+FIYKTdYpZ
aMGFJI91DaNUR9IhjjCRvZbVnacsNESYIiabViF9Srg8aE4+QcHRyghdq5NNwr9H
N0VURjGlAW2e0wQjGX6qzsubLOVSpceoTpWTaqkXGF1s5mRa4uv4VZh66FHS3sOp
sc93LfiCsbda7ufys/MLkQ+hna1nOM94gOCRSMD11X2Dc/g3aAaXEi7cBH3DP6t4
BG4nhMMA3/WSumMyJtVEbkuE2a3tmu2NAWfiB4bF/94K4/zw/9VtQltYq1c3wWZc
EeVpExrxxnQQx1t1yN0JEbI0mMBaKoS01UfHqZEkc8haq1Fc58IslMEdGFgkrP+x
OaHixVu31EFN0UrOd4KJR2q4ORCiIpdHDIilOa6ozV420e8gpK9ZkQrpsOmABKWc
QotQKiZrvr5gGHnh0MjGqKQ+CxOebwyoYS6PJL31Wr7Y6Zw2Qsv/qlGgdzOr5IQM
RtCij8uhSa7AoH+wYj9GdUWiAoNobGk4vdprojPmjlFjIE9cCiTSES9VTstx5f1l
YJW9b3gaaDEpdjcAPseSvxqZ1qbC39mCTqceg2OapC9mxXbj0D6GV7THySe4cNd1
6DaJFxAwzZlsx/NKdC8xYFXDa14oCyjpUbW/dD//FAN+oqOWGlkAYd4/6e1ameQw
oBO1cjwxoZKEZDuyLnnJn9SFYSkWHcwLlVdWJC5V6ce0NQEPIOLtPvwg+4nQJAip
tJJAaTd51Ffc0YhbBgYC9zdd8HL5s9BG5IPeeooAr3J67fHgtLWBftI/3hXcO/wU
erblN5L6v6pKV/0LFm3LWHP4Ab2Hs7G81WGwyUpCRvNxe7Pdj82/AP7atV5ucsy4
5OSIlufOPqj49ZuALeGDfjId5mHpMQaMNjriUA8KH75b+/talN64y2LpRymXog/4
ZFHD5AmVQua7TzEUPzuYvybNAlMdS80Tp0I+COGCgxztRYWlJWYl9wIRTD1JZ8TN
a/2uTWXJeB010AM7TCngxIs9wF9h0082kA37jQ9aLm3dJ+VEF7aTHKceEq5ayLZS
NR0ke0clF7rIggHdLyMQBO14M7WQSqgWxHLpf8pbip23nnpo15Omr5hMT73BsVOl
RKr7MP/O5pmTeE9RXzH/tseAfK2E6Vf9IK/OJmGSaJRGkp1tLck6gdm1lWLW4bQO
ALrNJrHLSupgXXUnbKDJYdGqs42D92PNF8hv81jIFb718pE6k+ciayTXnLjx1PgZ
bNfF5UrFMdqga0M73C8GbPk1s57pWjFC9/NwTKvulxABLS8rjB64F5rfB7dpdayl
8hIX8/l0VudknXg247fQgUXZinm6r9GemwlmQNWribKMw//lBHTmHlMqDQ4rebbM
zl14grxlbGjjX/JewihzKkvQcnnLa8FQ3veAQ/eu0aZFBXnVczbVQ/FUl1szfs5n
o6pIDjmiuQ/3W2ftnsY2qjiLyuO2E3rRyWaKmljsK/xadi4QVaSLxsVuzfc8JM1h
EXfKC/2GOLKKQOWrC5R6amh5oYl/KUKR3Lt4If/HFBdZ/TZRfe0pKTQcyIa/sKMJ
eroluVIJrdGqvDrnWj7r59CxVZemJPrL7oJ3oEF/aQQ9waJoWzNsjddPqIZvVTuW
Tlv7cCXcFTeoySK8kySLMEDva7fgDZRcM/Tx0kVsIH2XB2WlUD+WAWZ+uU9g0RNa
P6mhxg5EfFyXc/R31QQYUdu36rsQdIjFzUet2Afsp4EFMDaaAhM2Jubww9GjggDW
VfsCnSBD1dJebzErAro0O+pdpEkEBET1BoM75W7ERjyrvR8S8sCFpL/U1Cj1/XP1
xr1Rpey89h9GE3ck3+xGOowxV9S/TcacFy3w1M31B3JGAEKjTMvmhNZ0eRqjG2k6
NYmGdx/wSd07lhL+DspyDWzlyxOZ85ogoaJInwygJ4z0EHgu3q7oCkygOcUNuvdX
i4LKMYGwM5TU4nikcPcsgcG7wIRyBH9aPWCljpZWcD8Sb82cDY2503NVH8OLnUN3
pvhDNZvxD8N+KwU57hQh8KjCrfzHO25AAe7yNZYGaNzpN+EJUQCmFc9J1NEf2v/n
C9awk/dDhUI/ZwL11RNANVJkzGx9oMhfietslKnIHSzD2iLAXR2hVNWuL7zgPjvA
JyLzda1rvUDoGjHR5ldoKechpAKBq5Y6OX0YMlVxRPclPIEG9MJBJo0ieAu4bv09
neE+WZ9GgL6KOiRAQRJbfdqkLFlSYaJDZcaR0SedwiR6LueeFgEvJTfXPcB8e+s4
0XURDq+aTuw6zE2e3aSyG/b5TibVU7Ml0Y67KICGAyVFkm+oJOYEaGbrpWXrP+l3
EKduRI/Sn9yhY9EbymLFHKmlcWXjvEYwUZ7eaR97QW7px14oeHGss1QyiSuJ+h7h
QihbH+IflVOsG8FKYnfEYlPssOj37OIkeR7J1fulCXyBrlAPQJZOVE+f5yXPDorZ
wpTaJTXcTbeix88bto+s6+GASySC7AyZAKAHGeRc5p7g7vCG9fzMyrYRJ26SBjux
EwTAD7pLcNYLSG1WXPIuHEA7936lhBjA5uapxQTMF8TK0mXUqFXlPBBmxQyiTnEh
d6baWHsnKCnQGUiN8g1n1h6+krQw/A4JM+PinYKOZaoNc1wk6OlixM7vH6PI2vKs
vq5LIVz7qGw3u4ooIedeASmgoR4WMMAjxNIWUsJs3eSbLUGXH7wFe6ycsE/xJ2Fk
LfUX8hrwZhpqrIZOxkpGUSYqOygCWc390Yn/1vhGBc0WVq2Eie/myY6EYVsj+0kd
UxJb+NzKNuTLuxF/KneHYqYfQbXEgfFVnj+o7i7951HrtqQxg18Bjiv0J5dJLmzw
2xiH5apIw5eYT+ETrWQrzU46zLTZcgCTi7E9mgWWuUz6dMN3Wf0NItLlSrxVognh
P/rqBGwnul4hmJ7u9FCBLIsnBKfdDl4fwNLGuLKbH1ulfLk7N31k/If0CFJDnARw
AeVaGZmaHuNP5b1D9PsO8aUfaVaR5areXGhkod80VLN+y6NMX2khrSZwBnOsRf5o
nO+SggvjERiGRR0pCw/aeac2kYJVRmJztiHncYXSRQyGjn/r8+hZpzPNWw35Paj3
19OciixEKmjiGKOYGd3LOX29j83bKJFfagduiL82k6rWPSdiU9fw12a85UJFwIKn
Nd+by/e3jne1vVXpjOziBX51w0KvHQDEs4IvB75LOnAabL3rg9U9WOLhJoF6vkKA
fjm3c5jggxWeH3GT4NjtLDFwKTTIZVJtQlM3cc2cUZOE/EbWkcArlLWMHF14fI/A
dVxE2tf8aSvTFGT4zdFh4L2PR/k5LrY8dEqhRnPLCkLSBo0g9puF02aoucJnKcvw
EgoYhDmNL26+qaW/M0m2IxFhmOAA08+MtLBUyueTjXH9Js2s+K7fEFn1HxvGH5gZ
GmxcXs8iFQkTNUFeS8Zw6ADkcconlPuPT7nHJM3BXVqiY3Atn6I4Fn/6TB6lsIeB
GegCblstmci4164hcQZbb458VxsL2fQfqhqXCSsJOh2cZOMzgijQwXrDahUogZKI
MwM2TkGYblr4fSpczrYw9iWYoePEuCZNQaT6BqzKyD8A4OGBGgw7rNd8FqMDYsHy
05GoU0N5hpcHD/Xpa2FURopnknfqAsz3Z7KU1t85nhu681EBrrSBUCcAKdJPhjuv
krkQZ8JtIM5ayPWkOmYjz+hsvWByb+A1qFRkIluqwjC215w+FDsL21hrTOTMTUtf
+POdUaIwh3bFHT9lLatyRqjBBfBg/2vV0qfEvZ06cMXRSu4oVLQUiEwzecF8t2ea
0JFoxO+3wEoPXZ3JkHjxpWS9Zl9s06Y86YeW2GCFSWAG/4QnPNsDNWqtsU1rfmX0
GFb68nzcA24ev7fusGI56eFb7+gwS1qA9x2e6qgJA5ROcJgdQK+OY4Fa+MoemoqU
7z0grMjloEnBsIOTsa5FPjGqMfEIJMaky0k+x9xtpcuzTNnIHqNfwJ13fnVtfc5z
/vyuEvpB4jO6/xyxyoiGEtxyrM3A/vGYuuOLZzIXqYefWWcwJTrGC/N/gCODxkUo
DZFYDX+fXk++Fm9U/EollGPAuxrdGD3/r6i3GoQlakW776EYDN1gj+VKpPRKZgad
g2LlPA1uOisc5yMc7WG8oN2ja0ZV4brsP7Ye/BosnZOiLEpbsOMwUI3kHitZqBDP
xFohUfcK4r8/pmQat7BpKrYToVn0S6gHqtfvuPUtBImHwTTp0/bswrBBMuGs4OWS
hpDgsjAITC+pE2/w5aV8e4hwLlWAZqFsuSeZHocWsDHa05ersRRcek9Lnj/NOSjd
NENKMcs4lUG9iEOsrT+V1MqCSp40mZjgbXeT3dYGMeSa0vPWNwqaspy0cawY+ztr
eYpFQFHAvWR1AVH6+rBUvyrxe+YoYzNe1bOdn+LqMUPUDmJFeHaX9UJkI9qqG6v4
ZL24KaYHx1MH/G65ZSj/5g672uTM7UFMbbNAf6xOfqp/EKntJzWq9tcnHMa1yH6t
oPwDR1ihQh4nqqal7RSzsd+Z6ZmGaC8ypdV10l3QFwdDT8rrjv6Sd/zT2sbUPz8P
aYuZp2D1yPyKq4u9iNaAY+TsGnd+dm8LTC3X8iMO70Y7l3QlOV/kA+C+I3YooSwz
rDKMdUr+v6MzdcM8Z4E/NrvAsHPxnkL1sAhUYJp3C4Ge4wXeVOCRBqeqV7HvewQn
li/P33Yc2H2Akn19VFzLgC8e3rCwtpVBLeYIRCCmxgRL8D27FFEnaGtfIreS+pIK
FLC1tfO13fGdtsdEUD/18Lf3BZa/T4VCMzZPFgzJrDTUn/jsefkrDuG4X5e2nX55
mba9NUs6COnrJmO/T+9ThlNF1YD+OHt2H26NVERLc7hwSne0zDNbpHIJa23qIMXI
N6TntRMK6WQ+fTt7n4LlyIG84Y7eKuu+6FbBRBu4pfTObo0oqp0Jdl6PawCMMaKw
AUpij2WpZ99CRTSMSwNG+UFufhba51NUWiRHg6hfI1RhdHSZkigOwLm6UFSllILf
Fj1oJbyzQJMKQtu9NoBvbqO/vjZIZlJq9cyGa2ldClG6Eo/sH3dkqZ5YWjviKnRV
Yk+aDErkfxCnJB1njea8i97quP2tH2vuGYaoIaR/aA2n1xFGDS5yFsRN7sQlIMX/
VyftWpSPiEtdp6zTXkaOE2agO1NWs0C5AHQ9G22Z/eeJ8g4wcVYGWZuYd+rQjj6D
IJN4h+2bNm+xRMfpb/IaXLoWGva1b3JjtAfXLPyH7p/a1ylgWP10Pop5jPHKSkzJ
VY4IvBQlMwjlPBJiCgaSXQ5N//0Pkh3oce06jtjIV+gRRcATbZuQVC1BygQ5bwjO
dCQ75w91x20g4lEYG3oGSVlPWGYOpMLwxBiqU3INBKtFR04sEaBZNJXVNdok9uky
/wkMaBk9LRZiIesZRl8E8AexxuOmpFx0lnlg9zC00MuNHuS6qCSq0cKqoK74oTnN
s/2R50FVL71wdNLYOK7lqZ6B2gtCabBiLcrCC2vXXVpZ/VXNtQEYhb3uEQI+7Vsh
24J7FFwk8C9IkSmgTUFhJNL8Jw0zXfPgrW55S6ak9JpVBpOC/zuYLPHcnQe+Pdpz
9TlfuC95BxT+MxJVQxwDIqbl32bIO6+c90jhK4hFxejSGc1B9VFv8pQXIlcXLPkS
LfyUEzpHQ5myFhcegRDqgrC4+V2sqzC8OYVIJ364GmSGrVpNalJzp34skBOVhNwo
aWEWTPE3clburLE0rzBqb61RNhLL7uSwuQ7APkOqNgx7DgyXr1JdCi0i6ND+KTLM
9euWxeItGRP/1HRYOULXKKkxlquD87zNlzkxQIilX3GNjaXsJy5QMGAFyx728s7R
CR44yvpCsobTQh06OeSHLHeizK66uzCzPZmScf5szs/0cX3xfwA397IKWQcprJ+F
MIzjTQpl85YzPhlv2syFna0bo1RwDww1dvOagMQdDI6stEfCg3maBlKqO4/ZwVAx
O6OejHVdoPiocdBEfYkWe+eXlRQ1EHJaEIQ6rVWej8qT1deCLExuVlIKq4zdoN4Q
4fQMl2lQwXkcxEiwDj6Zj6gb8lM0nDrPrjGSLi3gNLGSoBcj4SEMYrhP/lcgzLaP
8BEWp84fUd/NNLuyRmcKPveWJljQltBydn4fbRC+GWdj7o2sAqvmgxndNYEt4Gc/
2n7autby9pJYpkreWTL0shYGkF3PxbI1/6FUaf1wCeFRURL7Ovq2RGdfuB56LAB0
7qkbTDus0NUnMm37Y/BtjfaIRAF/sX9LklUF6UtXavoEm0L0xH9/y1x5yHUGZk7O
Vv0Aj4K+wfYQ5fy1ZbBfmIS+PYxOOe01jyUTNKDUo/UbZHJAof1UWMcF7lzmCCpM
OvbYLyNBWi3DDMutMJuTISKCzBEBiEL1adyOHNcRVt3XkbirzF3n1o2fozhyyiBi
TYPu+iJSoXlGJIiiJ4FFvB/akBfILkwa7F5b2hIZzf/dvFwLmOG/YXFAyhosR34l
nzfRbDNBoHoB7bcfeMBRGYpglmhAwUn/a6KyoYHCKDN/4B8gejpYnoRBwy/m3fq7
vqlnHJa3ZMvG/BAT/sqoxkqsrO/WoFI94Bcyo6inCoB3k3tGKxR2/+/qW7Gr3KzL
WcnnFKcMFPkkUn3dHwNFOFqs6/7RAsD96sKSVM1EWcjBetQNla/OYza+obrQ7D21
M4Hhtn7LhZUyBSqfvld/GDpfj7GHF3/t05HtuITUx6tsgSlNOj5y4oAnGp3C2c/N
Ct5DT7xm/AWywf1EvgpzrPbR/mmbgsKgOX7WSUmKTfG21baiVq9sRShrFXLR3JEP
180Hods1GQfYvRLHgqayTauOHrU3vUYgb4I0wAJSx8dXVhf81th0irKpt6yQ8PN3
7D/h2pHT2/UHvlXIdyWV/lwR37dfvdPL+H5EeQwHm/Qe4pxQ6S1JvjjKdVmDH6E3
ZFRchtk9W3cEjdDeINPdbZU0DTF83s0EPGRvutoOidoJwZKmap6j5hTOt7zqGgpz
Q3sDl31os6QnpNwWQAEVGo7A4v1TZksnteDvV80vJAmGX1WDehmx113s9uGUqacp
J2E4j/60RKtLV4BWbJW7iLtKt/tu70JBoyKXOO8XLewrul5uBdFbjJIN4QduLJOT
MURuDHUOOgf4dbDXgGESyxF3oLz/K/8l98vNYmyZKOMNcaCyPWt8NJqC8uJ8UYtU
mvcRw4vNs6qALxypB77yKCJGZ193rWLhQvHG3S54t22sAbV0cxADuGnJ/c/SGitm
8ncWH6ZeuvItZCL7xMOXbB7qJ6fVQc8h0mTE5JCLWNfdtpm/O9J0mUIWBKDk5b8m
9rgwtXGF/ZsZXMJRp3n866IgN2LtpLhPeKiwQBW0g8QzPj/7+4/CJ7ZPHDPnEIWn
TRmwPCbfOc+csrvdNRUTNpWrgpSIq6fjuOdmGeyAzBItZP7hTxRIlQSIbKwojHEw
ePi9lg+sGPHjWeJTz6/nXH5uwaEekmf7ymZF2P9wxxHu56rFblwciPXgpz7B+QWd
Kzpi5CNO2yCYA8wlq+VQIyHlFrTmaMAc1LK6QwRV7PRNfXrs63+8lgYfX6zxoUoR
NCq3/+yVbwIR0J2tGCppqhMo+rX0F0G8fMFl66boqBj9wOeBggFaUrUrCU0h6W0E
qfP/Su2+znSvQEt/ojbNRSlL/9sXUjjTB5H8PgB2y7CV0W0nyyy6vqEHutOyJHFe
AKlhArfQHn1HqmblRRsIausDAmk15Y/HQ7xMEMJH+tESPuoaWqKGsQuRmWA7mtfG
//XSuoqfljtN8a6eUwYNl0AOi6KQCgekXVpzTjpXokPh9qA+cs9SrUQGdqS8/F5+
cEXtl/eqccMUlaskPggCxmWlCxR4QH7TApfk0qh4VLcS+MMTJpBtjg6rzT3kVEsU
KT0CAdykaHSsz1DrsZLg7zj2h68zqdaruLk50+rTY86sFH/GwsUFdH5MoMrQF8q7
Wavb0o1NVoYZ7W1hq65iP7x9g/h+OnZEOYt6bnxIPYiIeanPOJEY8tGQrH14Aw2f
Wa+j0iIxd9kcuS51YWS99n2AfMmQLcJh8cEyvNgDIihTZLwWEtHh8JSowU45+UgL
GlpQuKPi9hdGR2VVgOKiScDbST235PthN6KMHazxkp6mb6p+Rg0PkDxdfxE40Vi/
viJc+zqo5DdRq0OQSAiOkhUpB2SZntM1nLyN4QmLYNlSszY6z7mVVKOboTZndCbF
GfR2e6Jr2TxzrRstIfe+7u+mT4OIk9OL73vsKx5eXLyxb8XFlYiId9T/A4QzzHHe
RPFtGAodZt+qDCU81MgyBiEt2Oiv3WMhI0aILCOHtK+AhscZGkQWJt+WesZF2q3z
idvDMDHnJ8diwGxbyqyV0TQlU9g10s+Pm3KM1FbAn6yqMF7X2apS6gqDytQNJItj
Kx8yEavVCrla6Tz8zoZ0w/N5irLjtG83xMQU3ht8PZvAWkiw2HcwiLlS5tjJYlBd
yWXB+LkBChQQucnQWKAhejQM0lex38vZ+FN70k9om06CsSmTXqBfHwnY0GPPJw2K
M/vGYOHK0reX1u53+sM96PuwOa3QtOhmajVRcq5KPUxCjNX7gTpS/qOvZz27EeJL
JDp1XBHWu45HCImJ6zYO+7exySwHOOLYKjFjMeQE5zWk6qz1gP17AG2w8XmmzE4e
C0XpktRU7HckfXIX++mU/DV6lLRCwNzzs8caSeYhCSKvgzHQfgFIouBUtJcRBWNs
en3bk8Bf5YvnrM0gavHmEG/ICscqQ/07NL5WO09EF5WwqHWc7iPI/wyqK2C+/ws3
zOHGsFcuayTuxwX3wzXVkPEB1TpVWOejTdf8OZ+3UcyYtlApQu7TxmL3uk4PF2F4
1wRgB8U0Jq76QVVtPHrSCKjjrUsInGmWRHpaFJ1fm8HmQHZBtgOA5vgQ1Tvbvfqm
tzrOjliORZhmIUjdahOpGHfIf30nLJeK2E0b7IXvgXwIdn6TVd/bVVfs/ThBI3r1
rq7Djp8ao+8inltVo417l7yZXR6NgqhaKljeZ2/DBkQK4BfKgoTbDBR2XCjuCDFO
3yme3N6OQsoj0MOkkf4c+7BxPUyYcB3UadVRTW7AIRCjiyeTKzsk74W53iBca269
+kW0X2h3USsDO75GUIz5AoryhW3UdYC1iUt8eei/XDVPeQ5rtBIf0Azbmu7RadQq
dnwk3yZTitK+Wnp18/O7A4L/OB0S5T6sdQhvSI2sKbJHaP6i6UP2rjw5PJEznFhG
cMjuBp2KXo4sS1F1w1PGq9l+bMg+Xv/HnK+/olvKty4rQcegiAVSfzBnJ2UwRgsT
37GhD/JpvDvTMAonVkRqko/Fr2tmYPnKZ9uzyOVHkg/h3QhzvUbId9nyUsrABb0f
/8qOnLYTfWuk8Wb7l+s5yHpPv02Q8nb50CZoP03AYidxPpbId1kvnl22vzE/fdkk
Fy11c1nnTHjUpr++MKKXIzXBazN2z7+pO+Y7cVzhb04eBxoFzWq+idbeY2bhoOds
3yPqvHWhtqrOXwT6dBctic/nG270S92I3Uh3SsJhtkVa+p8vMGkS4Pr6+SU/wwfe
nVZZUPRJKSP0JeqNwGfOvntIzaQ7rI6fH1msewBARDxgLJq2OzyVsaAMcykUeUa+
EAOaD6SZtypE2nSiS/rQb3cA2wCvlSMCraib/riDa0sg2WBmOe8F4AqCsp8YZcmt
y6x/s1aCs1FaRPljhe9oeXNtMgyTCXTN0HayGuaEgtxKXbJPMPlxsBBBRvF5aiY/
+W/1T49ZbBhF+pt1v+T1o3W40xaAUs2T/wk27WFtSbgAYFs+3G33Hnq/VAVVmwA4
TUwqfNoR65yc7ADK+308tNvFXBevp+lYXgM9tukHK12og8fjwfZCPMC85TIpPH8i
AIXMO0fCOpmj6syJR5mb31JmLn+vuzT2js4YjcXovjEBRXcbMYs+0cgkmk9f4ijk
9JA7KzMfhxC37RgNvrRHdguBdOIrUQj1TK2XfP1JvuABY575Irvj2YXtR+FfQLC/
YROoYmMC1z/u+u/9Dam3ZKX4/J+y9eea0hAPagsmxWyp5j6djMu4Kb4LGa0mmEsk
DBHmniTDQ7M3MQ/9VM1lpMk03D1JKhoLhibu5OpMfSYtttVtoKPsNKU6TEz7ZDDd
C95ACfe2eYjlD8d5TfF1So30oXSgPhyqTVp/DBVm6dqEUFTkrdegu0RcRoH38uDO
52MVblfOXqcMnm7PeojpJWd+zFGaK3/q3x0T5k+47bVgreq10rxGyDi62tOCYujf
G5hSDY4+4VnSbvoMUVN7EL7QFo71hEmStOlotTE8J64ibh5uvVAVplrn5IxGX4Zu
yOipSlYcxejLyFkJS7Wxr7McfU9W1m5bZltPnahfTlg+bhdjRLLKfYzRwo66hD2e
ZlqBcrwsHyHMXMGWLSmOFTyN9Iw/VrvirsOs5oUAOe97371ZHa6YxKOgRqx4Azdt
ZFEidNOESizsY2nQvJHWZ4i0DxCn8ueCDTD81L9r6s1ujBaYmP3ZfI9D+2QRDpcV
Yx7LZBcuJWEtV4VfHszjkMThpl6IH/1ErAJeiOORQrMwd9lEr8LcqpatIQ9mZE9Q
q2co9U7dKAU8hPt+S/q/5VTjQWJkN2AeF73A/gJ/DTVfHHSCY3E9YH8F9L0OI8Cm
Giya2xoE6LEoaVazI0G+Z4lApEMzXKWZwJ7cCFyGPPvO+EOsj4bhXWuJBHLQFiL2
bHpK/h+efcuHT6f+9s6TIs3R8K7ONdsyyef/bUXq8vVkCqtNkoIjzWdR6q5pd3JA
J5zCPB8sFb/7LIucV9R0Zvbhpl+mHoemCSYUcN9p9qEFXvRa6c/mzGd/DvWaxgjD
I5vN7ihRx19souB628eg49Z3UwnlKSk/eoMcFGjICvAZN1JoH7axucMCiBi1e9FU
R6AGTWkw92JN5O22zZ8hndStMdCMvC7vO9T1J/s31CeojrQlGOSlgL8yuSHtPqdg
9VoTl0G8uCb9QsDMezRHU3G0tCSKikIovvqpqO50ejCMcUk4t/hK2jDQFkmWVdky
yeJNSHk9Pdkwe4NFEhk1Lx2eCODXEQ/0o0jokMBsW1gKpT3mGFr8H4qntxWZ9jKn
CmC8/Xyc2yW/LQzqLCbkOc7PbGbYR5K1oPG01D7xj67tql/Vv6P+zVzDJJejnRQ/
ejROB8fkce2wrsCPZ2wWVzQCS1w91Zf+BjirtTW1IMUsi/78dDdts1Vp4ACg3kEq
ABku9jMTU+E6qOSlnWHblT1yjigABwoH8qD1VqXnt3jO9UfwsDpakC/Ir1U7ReRu
BdJVs9bMoBDzfUDU1Ou6geCOJBdOSA5QtJN37Z7iE0uBsPYtzUQ1DfnlkCjAwOpP
J6tBBIUENus+YEs/hkhiS9o2NwTunS1ITpDaWXIcYr5xiNPvG5CbZzbO6Op+tsB2
Ifn/8X+G0FWv0e65P8gVNPverivI7q70OwB3ZsZq3HLhuL44l1f807PZfY+9wUTE
xFCJCXrwpJx6KVZ68eYos/BiQ4IyXWV+W1yKBb+eYtJ8VgSywsrv0H2B0W98vMR9
J/WAGURT9vXnUHYINtd9vAvOR4tgzMi8Tm0wITwzuiFss3sWtIfe4pll2K1gzTAg
5tz1MEHdUIWiKYe2fkdW5hP0q6RKjlXZAcLZ8qprL849cbXcBuWw5prEXzngKM3d
b0X35R2lcyMjDz9WjqP+0jOfASf04f7qb96JbYPyLJ901TQ4Zn4lgvbja7/SUlU9
mSPL1uHifMyK1DcGKgbl0rFoorUngjLQ2ftvDfBj3MePWjK492eEcLvQF06Fmq+e
/rQapTicgV9jMdLAYGvLe/Fozhr1yd8bBkk5VqPv7MXaxMp2jRmyZLHE4SEev+Qz
JUf7xuahIy78+ZicNQkfG8jjS/0WhUMOJB4gikUPhUoVtVlgXR8yzJFT1cjla5aD
b9ZtbZenotYFCt7y5wAc5F7L9qi4INMMnepE3GDWE28Qdl+rg+fCe/HqQIubg1vR
6ZPKyCXlKiKUh8bbA00Hljd04qmbTEFqor4yheNhzg2qKhQHJ5V4xdi3gRq218CC
hnGCFBr2GKfqu49m/Y1LFp/QViZ+v99nrsXbOncSJfT+988hOufolqabQWNtvWAy
6u/uhyhoTIXvDFJ6MAcxa35doXmwm7yg1QymBoee63N9OavRVtICVrGxipg/wmzn
A4qCcBV8ppnKGJ+0EoNDgJ1TXJzflROZTUCPripOioCB57xlJqUi8xFgthzFxywL
LW3TYMJciQyJpW3DFXHhNGaos16XUS81NduMn1pSYu2+1ofGb1eHG/SjsTuHAoee
JgqjsbndjDDM+zqfC/kmGM8GJlBzgPDWGIWmxeCHgv4D7JyKO+gNQ8TGqhoaNxLZ
iPxv/7qt7HwcrhgyA0c0lBZ7OhEdHk7uzggFjQuPMEPlYdTQtdqaJyUWWBLjzbtV
rVQJyPlvnUjM38eFqXjA6hPXPGCH11GS9Nef88POQhmPxcZbEbQG+B+oR+8C5jXY
cv1aXcILUdNNUnhV33XRALontJD8yTe/ZCZwoY6aKkXbJRXAlUIJaFO60bEVpw+1
90ylOMJk36sDfTKWuRZs64V64MsNqgEVJFST7qaoNkHyV94EvUMt5PuvFbw0cU+t
NxTRcHo7rlp5vAgvEmZPHk8dYtB+RFSPO9dDn5PIGwIzFNbqlZEdd9pr75oE+zRX
G9FmrgfGlpNjbCx0BQ3Y2p7h0XATHrs5l6ZphyI6lpnBOdhoxl8dptQvIDYOyQfd
sLnbARu//HLUcCaTkK5Io8U6Bk8ZDt7b9nUYQaB+UhTAiG3EyKOc0CRjO1fUhhib
GVzWjdl1ifsiv3wJWYIjjF0ATYrXAp1Bot0CwHB3NsKNzfH4pwoVHwj/w5e1yZUV
HVIVL+tLmKBgUP+/iWh7QjQCXl8IVAMqBsJKg7vsoZV9HDxOcmBT9kxk/r73hDPA
iQu1Eu2wzonD5lUANWaHbEPTUY4vpq3bzhuN1hKpN/jWe6IU90SZ60joj0GDrIwc
qLsHx9U55AMIZw7ikNBAQfP0kfka7h4o48bykOmiQDN+AQrMK1PxqeIfbB49ySK6
7KuD1Wn/m0bSDDpmTIdzsI+5dLUZJ23lN+zv1EXIdh+wtEkleDkpTwSBHYGEnw+j
ZiptYctHckfcyBkh2xlgvnqnj+tc4M7xutbkS9sQbRa4ssACDnOlWDATGijcgOHK
fHvsJjTVA5NAPLzgbdxeF6ltsXOVXDKTuDiOFIHIHhIQuxJ2d3aAboJJ59EBHYrx
tutMqiAFfizknb4JAQ9Rj+ht+esR3LLDpiv8lpTKCL8UxLaBhF/UkyOmRe7ZJrLi
f1+lrxY4LEpirwmAHw9XPDZplEcMLIG5haqSe1Qw/rfuhkldTQRD9+5F3+QFIot+
YD4BnFrHPaAUtGteoXAyAt5GD7HZmAbLY9ihM+DWRyEo6n+TfruyAT8UWK6qB9yV
OsA3TU94Z66mv1hqHT8kdFiyzuJgKXEzXRJwlQXAFEaLTvyJu9l7o0eY+9F003gB
+L6Ar7jVzohIt/kn2X7XcS4bTTLmVnr5oSfiTps/s89hZNc6/gC5udABPBNRYeO5
r/s/yLiIvuSwDiCnrCK4Sfe3Ht7usoDtDpb4f7VHNrAPsV6L+ZoPUcYuVdKBNSmt
e2tfAqZkCrmG/I6gtt80xXzddzPBjWXJ4EBX6w8bXHDPwnToyj+TJ5xmkC8dH2KI
l93lJf7msK9qsxqP+97B2oD+r7C/MmLNabr9qB75CuaItuxK0EbTxDSVo7nGVvF4
/0I/NJGEgrLUykuIvUn2X8wWAV5jmmtMishzBj1Nwnurw+lcfVhdXTyIjs/rclQM
q9a5w0quTYzgP+8CjuPikUgepql3uTFgS6ga2mGwk+D90CkhLibmBUfiWOguRwVP
acWgZ8QryPMlTryNLaMCQ1ZRKHuOP5LnJQae+PmLDsuLZg22f3hFl07pxZdxNFXV
3aO4YX+QyxExKPM3O3gDlh+Fro9EEJPq2K79rCI8RKT8ee/GqgSHK8OQoDCqAvv7
APcebck7WA8Rt6Q8DEARNeD+913oH9BNFDD5G94x8WVhxjtcjvIy04Wi506SZbXQ
hFlggdO7psgpiy6R8ZvfeEO1ZTPptdOZ+BIDmyxZbYQHEefL2Oa3Cl1mhRJF9gYr
ST9gVw+VBA4qQNsVuyecGWbt3Y6y5h+rh62S7VXjna+sd1+8jPZe7fppU6r0H85F
7NSJ4/XYVyITeB8i0wsS6XpyZj8zsQOKVHs3Sys+zDmyxXXgHFHhDTr2xcgdGDPm
1cUTyWPy50zoKvn8YrIiElt06ewbDELrtAl4Tfv13sQUv3HBSTU7xaR3TNjqJwyj
rFNgItGvdZD1HciHlKUsu00SLYu8qvIxhoXlHz4lWKTN8u+XmjJ8no99Z/uCPXkv
2bMh+tAfsTQmmSWqcPy53VgP+E8zPvrCdGRwI52xYYiAwpNk4j/apYSmvOVv4edm
Ex83GVwPwkCrTjFnbz4YbBjl2rqIAN1PbttKq3ViayYM4SiQvs8UJRziPhBCVowx
iXZq0mugi82thq6r/+BngRp+FroQIb6I4756TUOSK2PNaecjR5Wa/wUuykbvkwFo
IZrQ71ONyZNdebP6lUpBHFJud2KYSEOBR4MUqd8wDVxk7AwQ6+Kb2gV6L6QdFYwZ
aI7sQVYZKFvDKFysThUOlHq9krPIJN2jV9FMhRGI8DCkNFTDJG+ImE/gBpPZog5N
o1Y1R43Pr3i2q81/f/HYl6o6OxGV1dcJxt7MpR6UazWNLCt1PiMnU9xlz+7UFG+5
G0UvBB3vTRASyVXiLCXuANkaHkOHOaLsCrW60zh1dzduoW2fDyUrKg6xn1F9AexY
Q8DWtW+s6qpuHhf+IuoGq09JNPWriBhCC8LXTsYi9RYsJ/3uqXFmU1udnfhRtoys
5wh/1cCDHQLCq6xJJmsZfv5teZQXcTbOezVykQFkdlUIAhp3D4XaAFnlY5Dm5mOW
2RJhuKMgoStJQ7h6suSvv1M5wC+zWK87Ijn3I7SRQ4pKv2QuQla/iy1UoIVnRP6P
hzdUnmjONPaGLJ3kRlAYzu3BfrA+Vm8E4YZN+W2nkKG78A6hsOsdespfBdqbx0ry
LaPHqYXk00BPKZ7ybkfJL0sz1l/TiRkvmb5XWTysS9KIHAha1Mju7k+wuYtNo6x/
5PdcKk8d790uOfIeFKoz+2XVVuqrXuTXlRwprL9rDtkKGUpjvd8qRzjSRiWWTct3
AApvrtA4UPnzuj74r/n+EYb83ykR7fM+AmPS5TEVv5pe21lfPJcePZ8/UChi2MZM
0DV8tdzS7KlzrRX1asira+hWYj/SZ/EBZYAx4tb6vC0VJAI/MVeVgIcCKkqj/uP7
fskvqrJJM0NUS3FKxJJPdczxM4mYnWAXVULXtOwfkahnZTqn2+m8AeqNOB727ZsP
o+98k+hgzAMh6jKxXc4zyOLFjxv9C2dPhP+YWwvUIMBn4a9eSzTvwFo0yMDYkIAT
OIMyzGhidz7Nw3l8x2G0s2L7FhjVB38uJHvmbsmlCKTPmh1H5XLfJbhRW/6XyfGr
7XTjXiVTvrf+eN4nHdNr3Uz+I+snkaPv4vgFUSBuI94EEkzWCzt8YDrVqsHCAzap
rB0sk6qnInismVg2kmfRmqPqjB8UptJlakzqM8HJ/54mgowHJJ4Ep/EtzRuNbyKp
oDCCTj9rxV1fhbFTZU7i6qB0f7prH4aYGB57ZOuVFV3Ep5HVm3GcY5ClmFC7jVKE
RnRrZQ0OeGVLnpRIcXLmPZw9nk16qE00bpZOHM1Yc6Ry/sDgHE/SmqN4+/utKoiZ
eaRxnHFXn2yyLprwv5tVKFDEcLweedWnakfIWaojWJaVvc0tEhPG2k/dfXrG1ljU
tCffuW9Zfmd1d/YoO5lrOYIiHbXlgjHmywrPUQ6rwjAMl4uhKCnKqfZvgwaSHsJj
Z/PKT5Hu0/c4YKjlcB9Rq1qVoqEwvwQli7VFecZV+lOhkRqS9OPIu/Ly0JdNAVSh
IlPMqaiIuawinR6TFLxjy5alfgZUnPDQmtqdIapQa52U/Di0N3lpCa71LiJLKIDG
z12g8/XSIyQcE/0GtmFe43TUSh7RuJejcYyaTdoxPv6ol7C8jKhQdDNRx2F10lbH
BnCP/pXU5DiMUWJPX4K2NUbah4NNaZI5PSSrpeekY3YcZHm9sjPvFC83C1it5kOO
mg+5zSCIzndaxMQ874qm1XNVCbfXhBUCblhvdT7xGTtOB5xCOo8EEYr595UKRNKF
eAhi4gPwL04/ZP93HRmWUSXbAk3/MuG5+iQU6A/3yq0eOrgj9zHYJA8CxTTuYq3I
E4/vh5y7rM6hi0rOHa2VCdmzDQhFK7HLZcQo9eSRvl9WmBgUnoGiZyF29EE3qYlz
+JnguQqZOWzb1Foct3Io3AGvkp1lue7ejXhZuJzgx4HvKHyI52PwzVoXHiqUGjgE
0v5tBrmUKlzUK/xzdQ0mu6wxRLvxrxV2ipDHKit6e2njthW5bs+KOhNIPEj8uuP4
lTxJuYCScPZHZT6+RjEBRrLzgu3LCsth6rAt9fG1CBsKw2+wGn+L+c/o+1zcIJ94
2absM9QDvmaAkWiaDPMkpovhC4EjuwJ7n561J2Lrc58p/3KfUVknDT8F0wE+dUFS
T0k9bStn3dZOkoHGGW+0Wy0AAMNimA2E6Ca9m2IAyirJvUIUSX+7+liwQsga28Xd
THDeRZVIzBGdr9VkiAWv2IXyIecQ+ebYBC0qMoECG1uNSmJY0uRW7rOVrdhcdiHM
JzrB6Z6WIhVbuEV0SfD/IbuoYTPo/4qQ7kUJ5eG+HV26wSZmIQ+nKndbs16fChpi
2qCrZ99db+olNVz9mkNX9WFbuuDK7+Bmc5Wd/uF50UZuS4Nz4+9gpmcwcQjNKem8
l6+nMzmbnhbarxXuNzyQ4wA5MD3z2Ndy7NW6JSIGcDgBaKmKQAup+4E89G3qqBEC
wJB6pQmtcLOC6v5EWj9YxeV/woOLHuaxs5khmiDqirZ5MNsM96CEF+Jq2zKk2evN
bM1DW7r3Y6c83ZlgdBA7h1g1p8kqecGGhu8/fpnDayDIW1iA2mmzog4I0D8YcwEL
hZo3enyuFnzKc6Vz751eeMqVPv9mPBfEnO+5xALslaZCz7QingUD4QejF4c6uKY3
9G7Gora6N81p4YL4gzjw9haQ4HeWfQtSdNBM9CMzexRboVSOeYUb+dkJk4YMuSge
diN0F/TeQ+b09C5n/JVRjo0/ikL5aUztnQV/0PWPiuS8UpAUAMfFOxylFBvjJkB7
HfxERBBXZOZHbsYXQqXvbGIEwb/OmxGWRwglnWeWjfC02krQH8t0QFuYRpKQdL//
pXNwjZfSvWvyuBBUdfKiNegjcqSf4ZKylPOaQ75v5nV7j0aEaFruZZyZ5/Xg/U9l
zxtRerodtyU97CTeTJD3WaYIWjydmBHKidripsj66Yt9AV4fsiYUeTs1/NmTqJqI
IUljpghAHlodeqdKv927pFpasQjL97+doSFHi9nlxmqaLwox23h4QVSJWbiqxS9L
RyI2CMr2Yr4OPoFM5Qh7ynkmcAXotHflSoSpGAgCW7xAW0Ube5/Aj/Bc9I8uBaDg
nwCabNoqDxEewBItlRjZ03maO0qPnDabRdC+Xp+gcFdyjD/GPnnWbX3erE1NfTAR
BPSkutUfP5HXVAo0QIMiGqjV0xMLOgdEEUKJW7dLt7sxGISPWFIgBkbxkg4aa1Qh
Iz/PCXoaXHWVHPyN3Pt+T8Nua1q3HTFx14ESRHW1C2grigHcXg0bstpJzAGBdW95
GmIr0sm6Q44z1AeOgMqUFhjpctD2vtRgu9sq8h4X+JxmL4W0PlIhv1eUuntiqqyy
Di6jGAb+NS8ET5VMye5e4bl+2WBgw12N8hGbjiReAFdFYSwrBHd+ovb3j5kjeYg2
Pg1UCP8U6hZcZVLz/Equ2kTB6pi/fCUjU9wg3HTSqgXB+M7gGQOq6Ojz/ivqfVTk
xCF02p/PGHLLI7xONeaThUMhYClCpRp/X/ZYjyXQQCrjvCCHN3NpBtZCPnhbl0oN
yXA3BwktDHRqpW3Lq2wvGcSA/Cxl2lrz8oyMyYHZdL5w4uJOIWXvIO7a9iM8wZkl
gC5Wp6tisaY5TBKU6OHong/crzV+Pr8zNNxY7oqo9X1i6XAB+8VgXV9sza4K4d0C
JTWjZszOVY00zb12G9Y/g658mXI+DGL4XlDz5oq01lG6xEBUCUn5mOgPo1wNGy6P
zdJsW5xyMJeiZsfksjESUkdNEvI0tvCZxRRw8L83/rqef94niErGI+t4UkXANlcA
lPWHG4XXQyLcKl3JdPievX37orRG+sWVK9F+mwXkns6xTYKGXP3TyGyAnEFsUtTw
AxLbcQVmBrjpLlTeUzWTZlUdzMoDJDPTB59cSUSswxlZ06aRkaJZ7EkjD29hs0pT
bkQcMgVqAfCY47/GNIbE48aizOgAkSZHb08bA5aHTYhmD9kZgubfzSPQsMBCsFCx
BY+AEuQEp44nS8KUR03q//kb1K+GsOC9a6rpplIRn4TFTqCH87QN5sZZnJuKV4Sc
2ZFoUkJWpXNuCj6Lmw2+IGHOa/H7UCkJjctedOmlOmgX/TQpagSggII7Y5omHfHk
VzChkmbNDI2PVsbK+CDlBdtB1k2bBiLoW08UtzVq6RPkZdzFtUIlPS3tiZbXHQqR
C8qOo0kYLibRxOQWd1+kHpOKsy0ywiFxor+SYl1xkbwcDu//V0X8Y05PXe0ioAAj
pm/6MKYpu8NjHZ8wUbuNjB4/LFKlWSeCXN92m6gL/S9JPteA3NAPpj2KPgQJ0IEJ
DK1x6DgcgT+jDoVsIuniW0+Buk+M0sfgWZm0jgXEUlBWUSWNF19eDPuAS5QwP5Q3
ndEOGxZq3r2NG7nkTS84WBJrkx89k9QMCVyp7PJoHcNepU6lqBEuPPgZkGmv5Cqa
uZq3WX1Of0vcTdUvheHWts3E9xr4e3M52fmTOU+cFRCnGikNuRYW58upbTvEvFQ2
4dh4++oXqjMNPOmOdJhBV3yado+jDGjjXQB0e1dWojNeFiy2SMhlq7P30R1qSlCO
vOZyCL/IuNJdP98NVhCDbg==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RGmrXSBpGvzQtIlSfFGZyubpD6OD7nkxYErvk5OqY4AbU8T2zk4D8r7bJpao6v+C
c34wCr53xlvX64G5iF5ckAMgA29TlDhpQJxMYfYyhsvOFkDAg9zvSVHcr044itB6
tYeEq2auhSnEv80qpAQ7v+3kFJjSr1vis7RMMDLt+2+JvA9tvqCxkFaj5TBFt83d
J7h26zrRT+NG5O9NsWqzbavQPkwi7jLWjJ/oVw9C8Dbb9ZUldBsURCEU7fnA4I1Z
8teos95eQboqMVXbkfhNNYRohLDs5+/StUmOfglCwJsJxfkAJuFPahoR23HgkbcW
Gt/dLtSrMFk3BsTYV7RC5g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4672 )
`pragma protect data_block
eKiBO5pp1WcNwqLAfpYgm9R+G52oT4Y2QOhCnZFJEFXzqiDaIRqXXFDevmgx9I5R
i+Yww2nzGlLG6YqSaJhul+xXvR9PDacVsWp/DHw+6XLiqI1U7W+IL21FzvzrXvQ9
/mGcXepgr3n9loZfekWavVUogbvnvklkIlfMVr9WqObmXlDZyBAB+VBawVqbrv7Y
49KVQ1800RP3bur6o8PIaXPeidEkzrREymSsDM2QDzKyHE+OaBEzGVsCyVxGkdUf
FVhN7ttcCIs9/c+MGD1gocts3gpQXgV4GyTIejOZtpzgOxbtGBMtcw95BOVOndzg
Wuh/OjZMssXcgJc+FzjT97GzU4NiHXlGr+AgZPRDqzXPZz9Hv/omt1zA7XVWdC3s
sH6aWBtvzRwU72qkUbegY/wgbDUxKiAMAsCbB2Z85kOmxln5Sm/eQn6BAdukkupc
CDdWn6vfPPbnetajn+61MaaOAAdFz19rZ/9UdVcafEoN5dHfELCwmOv3CQ1uqt1U
kW27cVs/vqhc+4GX2xPHRrJMXh+7irZ9uxvHsBLUvPgsP1iv+p81r9TbwKWR0hF/
hqQEYpF1TgUzWI0Ig8MuPDP9aWAYmmYBt0MX6dkInPzp3eSODp+JnUdR7fyV8A0r
BKgmSl99P4xxJ36JyHeG6sML49l8SZR0B8t1cT7ugG/JrrDBsizKTFD/ZyNPShRw
B3skCBWV3htdrSdCINiFnWDyY9B3FeYZpqzW/427LdFpUHhpDmleIjysarPg2BnU
9/5WEHSkfq6K+1kMI9jyNqwYeMtDMTGeS6BkNs+gUSSTyJ8l2nPTELtgk4nB0rjt
kHwknXZv6D7oCBIBN++oU88lI+vphlQKPcUgJS1uuleQ/tRVgfxROhiWYE8jERxY
Z8gBGydv7QOr+y8GvtTkuMntfNy9X86eRJKLAR2qa8Ks8FwFtCqkzmL2R8yRO2hA
mYMcycvVkZvJJu3eui0aT1Tz2cXfmmBo18VQflxlXqmxamNKAy+BpHYi8DNROQr3
Y8Rbmg34ovI5pG7tOTly8gXxqnVBkbxreLnmtf5q6J42idkbmBCgkouYyBq4Ji0o
vS3OZWZqWaiNjz0DcfCYgp4Jz0hiId5KxClov/9CRgxV5PcSFpIM9OjHqTEAy2cr
ZDUBS/W9maGBZzF58qG8XECl5caiOfG1YgXprOR9yWgggEKRrQmS4q53NStoh+fN
Bls7BOgPZw/2LLCtOvtJ2/w6m79y4bbpsY/kqYlpwzSg+69UDvPj1HQ+uaNpZCMq
WbqB5c4F6MhzY5CiwrZ1kaxheLoR5EIC9MBpMFcXqTNdsjWeWxxSkZoQ7u/gBfyC
l+/L04Qa0mN0/ejfKNnB3+pSOEHyZZ4pPQl0MXYbxGcxk4i2r+gDV09B9A2D5LE7
qWc6/0Tnzm7V0cfajO1KEl1LentzxVzVy4ZVv0W69qk4RtR1aAbtbYxJiP6l74Pq
vbJ2/acx47YwA0VCDgPI9H8jGBGAiL+faIghwiHllEeRbnpyV0qXLtJgxZrHT49I
Y974ojTQQoHtbBRD0Wt48Dm80bnclf3Va70f2lWoPYX3nTRQrpDNkC3MWAJN/MFT
/rSE6JKGx4RSNzUZ30CN7BoN+gfaWahUxjhplkfZc4942U4hMsAGTroT2EAnkaun
YYpXxwSig3hf1ZOk1tvRPKVdl4pf2Zl6WwCZfUxPdbei4HbKhL5SWvWc2gKwVSQk
O5Z196tRX5w+zQuznIucKWzHQz4cl/VLXtrXKPFfnq+KJ+EWmRXEccwEr0AC1Uh2
PtjNRcQ+W/DOkhgOtk8h2/+TAPXrfMVB7Jgn8TcwdBHpxptyemFyG91l7TTIlWN8
7GujDgPFUij8jQQIdiZMn6Tt/lc2nsE8x6ZW9lWrN8SpxhWvM7/lLwILRDttzARS
RKm+PbyyIHWiuFgxQnSBmlq6i4zX+f61nY/rxdkDtFXTmemSgq8zlaVfbPWEH+qH
HMSks0liBGnB61SC5MdUh+q075Qbj7c83PwpBn+zAd70cJB+XA35aT8n9q4le3p1
knFkUK2rFMHVAi+SrNIwzrZ+qO4lEr53vTP42Q2bXtCkUypnyY2vykHCh1nTkXvW
RON3C/ILOzJQPonAl1IaeWkDJ8mD8UzGGjNB2f071e5wpq6dGxFmCBqnl7lLxlDU
ozb1hf9icvPEjlRyMtXl+PuVy8WB6VLfzhb4AnNtxxJL5JGxiH6TeqbPBkDGGTUM
DQX6mQTDHRYrB43M1AzvcSijE7yutVzR2456pxvh6rAn2oBKPHwI/EY75ReDotvP
3bTLCvwVoKsFvoGDqZyniRcGGS6lMj2F7hddNkpYhgifibC7olHqb+YvsyQnaTqZ
9iVmPmMq3FfZ+JlTo2sgOHx9V6DJgjK4UZR0C+dmH/dAuTDf0DtjytOgrYRO71Fy
0OzDC3OdtvDsxfJPbhjVOgqsDGH3ntqm5Ckya4jwdNQebS/eWU+jn03gkyfyW+vA
1jGsW8W+LjGv7ACZzQ+zVUIAo1rCiCGkewEUPM1cOcMhmXZeKJ/w/CD5fBEHepDc
VETBhROL4QqZkKy1LWY1UElrjYXO66+ZX1Zeu9R/Z3hlSbCFqWLrSLSsCoCzcs1L
ifKMlYPxMZt1TXPDeqYDbRwmKs7wNbxVizt/PrV3stjWoXcx9kAlsk7DK7ieI6AU
8CPNxIKP9pxv+clYdyxW6a92eutebiMiqFeN0xT8Zd6gGZAXxnB+BlDactEKT3Vh
AbjSsd8JbgXhjjHWy0hxUsYpcd7K8ooq//YhYnlaflqvW/dLTUyb/3PAppeCY/SI
jJTecWOOj9gd2BTzIgH4ZU1zXDLQFnW/YyFkHjzS2dQfyyCwqZh80N/a9l7Cm+gU
Xcw0P3VFbTFG+JB9OuAyT9IhdBOGWhB/1MaUX1DT7drhk3XSWLhh4soU98ZaeObP
aKvp2iGmkKxEnLjwJuDYCWbOGqAZTxmo82iRENnlNHZJNmBP394bBCyIGp6T1h4D
BFan0zb472aryTzfxHe15CQSeffRlZhOG2rQofuCnMS0YGtxAGz22CBGUsjvuaia
HUl5pPHIxz+OoXxaRR382zSbQdcLfBbsk6YmLjxR3NhC4E4H7ueHha056ds6eWTi
LJX9qWqWqMCxtC3dyXdSiTaYKVDBmZZ5B7sjkSRwwJoBD59OMqTqHyjzhliMBWBW
J2r8g3tnV+yyJBVNlqvxGHU+EhNJBwzefNAq1OJXu0LAaMF7qwtgK9wOmY04fZNJ
VimLOasOPJIc+YlDDnXIwKFZAA+G8j2zJB1AT4GJan6iV2q/5jqoEGjQA2Nr8Qem
xyl3I2uvyNpWyYIjnVv8PBjzjbg0dYtzZ61JRtphgZqr5PlMSG5ARzXT6NlH6iVD
nM7F8n3u2qXSQ+dlu7Cri2bsFRSSvhbXpj/KiYcJZx+GOdTpFeSN8y8bDqrXwdAN
2qBlKOwTX6l7G2simEst5xLyS1gHCbie0XOgup8Ld1NQpQOvDWi6Xl/GbkuEkc+9
rDtSMyhhS4nUWgnebg3Hx4uqrSQYvvuBzPa+0Tn/crROnvoEKe/2/E9hDqi7tpYi
Pp2TzGF7y+JRxP76VKf/Ldn/1xcab0vDxfdkKjOKz3NBVT3QT9iu7AtVGYgzCEoV
qFm4eXEU7va4DHprcH8vrtiXkjwIQW6wN2MFS8Sf1dD/NJ5DwzfBqtKYEMwac1B8
Vvmnf15LYiQddphm6O/UXUGigSZoIzG59jhg8mS64ry5oRe0sdWLPvvNrosfbF0i
EA4yPlhRXl39rkN1rf5JpOcRjcMXzs4TA2V8SqdoX2eYBg3x6u3poeMChLhAcSvE
tSyGvnTMrpyxYYTeZJtH45rS6QYjbuaIZvcb9yOXeV7zp8gLGXuFvE6gtBua0uMh
90z9r8FUW+vNeEnI898HeSY/evvXicQ/UHeOnOSkMKDXWWJ5Bmqr90WFSbk54X5g
YqE9HQ71qeAakibXX3CbPZf5dHgMheO4wxsK7g0HYVxlHLm+XkIvAwgOqEaRQtK0
k+OcrvHA3wSRw9jlm9jStHJGup4qCjt8kb50rfxWyhEvTlZoTtaUa3wLAC+znNEf
Gg1C0Nc3dl9TvskNO/DiBXS9DpDSGVuHHVpKuyKkOIlmwVPnhM6RFkY2WPtLHFVi
F01Xp+BrwzgAyzL8fL1qd65DNuQB2zHZq+QBsEadSBMzTmi+A3julCf77faLHvOo
YZ/dcl5b27iYEZ1qjhJQuIRCoH3RHHYZtqt9h1lQ5C49b/mGiZjOlHMYJcxIXh9W
muEwT3wShVfUP0NqSCHIvTKqkHlyG8sZoufNlotz39sMivrmF7tK6CZCuGItPwnd
Edhwg7I1EyhKlbTLAGkUc6zzqaSRP5bOvxrcJgR/fu8SL2osWykOtTeeAaSmu5yW
zD2a7unhRdQBXtWPyMLilbYrZqCtdaBWiKyMEDhs0kqRQXeSFl+XtshezCKOYeZ6
oh3FGoUaoGZ+q5bs84RIXR+SxrzxzxLiNYUfrUkXonrqlc7Pqz6Nn8BCEp9ID+RL
SbRtXYGlkad0l5segA/X8fgMg+CKg7JIJgsljD0Iqp7fyQ22SrQpjC/VS17Plssp
UIS8AHXrGuuNhtGOmLeOvbChi4piccnH7u2Ex3zeyZ4pihQL0sZJhISMej/tIVBQ
fz4V7n6yS2IPc1jvMZsg8A1oKDRvbRP0yc+WswlDVkGiD/xH9kHvLW3Sg24I5A8A
UBOrQG02vZHzjDj1ufsaudGBB2tIJVF08yMv3EOXlq/pLlAv0hL0fQonPr/wHLjq
c0aufmj46elDvDQjHVSe1KAwbbQjiIc4p+iMARYory3cLP8qq5ZDHTBUU2Wqmv6G
yCpDuAx2bQHPvHric9u5AMQ/LvZpPmfo2IVIx6OBgIRiPT5Y4f/Ixm3RbLQR1Yyd
gr/7vBirUUdEfEPvuNRuu66oPIPBGZzrtioXBRyk1lm2MXZ0iFvEfFcdCCqtUrtx
kypRrjOACxlGGOzJ2ykH4y0tcdPwiaJq7YfDZeJmoaNZs4LBVTC8NjISmuUigWwG
LOMnMR5seuW4K3vJZfIea8nzlq6cRFXTN4Q7doKe5ETQsetsI5U4nXjdW+s+/7f0
RG3eXf/MiJ0CezBZIKpzWEQ9GcE+8pLYVwmSEpwVEfyLkpZ5sGiQJTEXLZ7WLUYX
p4w+YWBZV7AHqyf/iTSYC9w2G/yxFjzI5/ndccUZBU7rqfvjt2/HmlxjSF9xOORO
I8DaMiC/LkEYdqeL7BOd328/mX0EtcDsZ+btYQ6zh+nJoyS1SvmEdvr829BciqUU
UI1jkbeZ/aiYSvOHCFvt43kzk+O3vhdxDJpsDOto2heJyMeK4UX2hmsvBrI2uAaH
1VqaDC1TnSoysk/GLMBNA7AyUKarOl2nGi0hSu26gqTo4FfZyoQL3+g8EBHReMRx
LO7RkJOAAvec3hUcYf5PnZPzbcuMqN29YW0dwps+76XL47lXpw4spQ82VmmLwcrJ
AFlI5VR2IozPvd8O3iB1FnfLxvd9u06HUitRpl8M5CHAwuC8QuQ77e+6HHCXfOuQ
xZ+Gwu6NOUAyX/bwN8WadnHTB6g8tZEL82C3m84ajbebfZAKLJwD53bDzrWWg5aA
eM4eqpBg6FhPBVWin/hy5120RvUMenivMKT3/WC/bwLXJ5O1Qo6XDWoxDhDXoSR6
wpRavH9VMEN84xHwwifIVijX2WfsWf/69V1wQ3A8pMQzMwsTlgpRPr/TwasQkDkF
wc5tBSJJxCcVSq+MmVfF13tfqeoKPWg0CbHNQjF177nuv1gTPgs4wICuHt7jqy8h
qTt5AeVKNpJJ0t9mAWLfAnf+c2E3Rc95GKu3WUMi+sAfkGCMb4vk7zwf/Kc1LcHy
RETwzZNRbXBbMrEbQzCGsQ2hLdEFNPTzZPIQio1OUr8HbbFPbY1LB5jGEQQM3S0B
vxOI4au7kQ32IJK8RBWRgsdnR0NhSmP0LCTh69Ay5pqdgmDIwTeCs8dB9H2LFra6
GuQy07L45qGgG1jN6UVXMlaamHk5NUE2nusOMTuxr859W2ZH0ngn0iULLfc6IoOP
JytldBOSw0PpS+qWmYx8R/q7eRj8xNKxs+ZQc78SF87WYCnURrHw8VIuQiNmdmVj
gCUYaS+Jc9olZ4fSS/Gh9krtEQM+PWHLHW3wtIYx9oir7bT157wccLuEaTsFBcia
LfR76n8O9R+CIxXCGBp5qQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
J9gnw4aUsoscInV3O7EPD8AU/ULwKkGKtej8oURuJ7qZeIaiNjxr2/9dwZVWTQ2t
juazs/FDlzeU7+uEaNd9jROGrvKto9aIqzNiZLXvZaX+u42KjqZlE9mwHB9rnVr+
pyRVMo5W5Oru/Rg7uOl97/3TwUs8eFUkLrpz6hE7DfBrA4k5ucRaQSxjWblrYVH7
SBWshX4OFwBf0YhWTScHZ3WH8knxyR2CXqYMwVH323h2FEt3ahjhbKZVqHnCcLoT
J06GjCvoCbr/8/R64dR7hVgA52af+NcDnrJNtDBY0yxlOCGHU6r7Y6vwOpA0gQi/
0tLkMHJ0J4KPgUrtAS7tjA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9344 )
`pragma protect data_block
p0YdwG/RreKn4QuTBJts7nlTnskW/wtlB4hzGJLi+K/PSSPXzimyzeo2/pYpAV4R
3f0lbO1oQOovsXsuykg2wmEaYMpkpoXs7OBZ72Yh2g2dFyqEpwE8QOisenC37MNd
nW5kS0anK9ek1FR8vMzTaOFZsaQROyJEi2vnrc9TEIXr3iim6U+yVnxYYC4Ren+v
IJPQ4URyWgl5eg1MBoXtLh9m/21ZYZBRX1GC9m4hLo1t+UduzPT/1J0Svpx5up5t
Me73KoCFHmRNGpH7AqQBFxsLpsZRXXr3cdG4veq7gwfcQaVqYXvYQNQAlWnxkD0t
ly/gygcoMAM5geNYqpdNJ3pWJTqEW2oMNBvIOTZs8aDI8iOKs7F0iOYU5PJXlosx
NqvPHoAJ2V+JQz7wrRu0iN9tKvBYlxxQPrTowatr1J5Xlj73QEZPDwgkR7fxPhXv
MHDf+fHpJE+KdilhCBWOKPUlXL3Q6QK11SEEtV9ktuPzNrbnQcjnmA4lsQ91wW5p
CL7bQfykX1a6LjVDq3MVLbyEhz5PqbdUmeq1A8RX8hnNcoU/ffK1Vs/aH8sbZ/FN
44cHxrppV7J9DhecuO14zi+0ZQJTdZH7keYiEkVhlNiTOLLrn8TwcJMX4ZzzroEz
pnkRf7SnhUXn7F/jN0aOimS5zsyfbFyiYROm49rhNfJWbI2OaHElnjgoCGdFD4VS
jKP5awtt+LOmdbsvnTAAHC6RJKWTDvI1S8Lct833eNByqq4LbE+qj4b8Z6Eait+s
mY0J94SlOLTjwtfUeSIj0rjg+z3rLqssk5XI9DYjXHtXjRkhrgB+75QIfMITLOGl
ZtVZewNefQIiYG6OqoGnSx8t/fTDw5WAmiEzMtgIZigD/RNtMs2Mdk7QQPZcli0T
9B+na4V2tgn/KzJ+lHW+LW7SVARbHDRcKtDtE4hEF0WMrmWh62mDO8/x+wQalN1G
tCVHsJsOhZ0ER34Ry5qmeM8AFTC6vT5NaZD5w/OMLecbjOIQaRMruT5/Ty4eV5/Z
zqRXU55YHAkn8ESTclhUG8To2CLV9KKJ/TH04rvHu1IBxTaxXTioBDZbPegrGc3z
xW1AyxRkqCWopIu40Hcmv8DL9DFLl1v5UBxGlkMOsyISKyIAb0PPqHwcTPASnEni
qnScRK/Bja/j1cwlLyIMRIPHoUh+GxGjc3umC7r0TkRq9c1X4aPu8MjMuFzI3Q86
MIlkuUD7CnsXtraXPxkOew+g+ZgmDEVoEwlxCt0IODVHpymnjyVt/LV2FIJxJDsD
w5B9EyLeC5jKiT3++jobGePLJ+TWvFyHy2SOJrI5P6tAmOouv+pHBzfvAqBLnPpW
F6glJkvpOpr0rXrx19xd5hLhU7US/WoHLI+DzowmRPIHXryoDrangeH0IN9t5WeW
RuNM01TIht4koeWNcDbo3f96tq4GZLYtXOG2W7jmszAx6QZgh5/9wNd/mtF7JMjP
ECYUvuUJMo5xM3UTrUu1JPKRIHGnpYJAZqwYJwqzH546t9bhPr+CmuNwBTCueSRr
rXuRMZe5TdebPbK1Oem2K37gByTsvBDGQGefkaXA2NaFAVdH9IjZzdTscCz3uMgJ
L6ujJZmQWmQZzts/A6nxQqkmj+f0JXvIZVR9rPXE8LEEBRELjQ5wFMGoP8KxFuuN
pyvEWis0Z5gsrgOZnzoZCxcGcYerLcY6KU8YXJzbxXMdX8Z9dQbcQs2xGRzZZtHc
JUD1UQWgTx7xSoQvGYPZ26WDJGz6/pIl7/NW+5dpT/fl2s7VzQDJO4u29bni+169
Y1oXABacfcuyq3ekJMHRDl9vfAMbVC86RnYIUpNn1phckFbnyoHD7DgL8bxXnGUp
DQ9nes6J00r+N/VpuhcB4JUrTJnT1oky7ZvJMjAzf+JOFuczqTsnkWLj3iJxLGHy
6EMkFAbm4E3BPVO6XXzXsVXSYcTsBTVdoCuP+KYxPJkDbdRD6lpXP1GPTfyXye+2
1Rjl4Rv6e8kBxqQsh1wEnjMm1IhkdnkhUTA1teWo4rHYEOlNa6J+2UXCuBdJEogV
4/6mltm9EMoDF1wcW5MiZjTY2VaE0a4MoTEzqZtpW4RjNHSm8LuXomtaJbftHMQs
PRNMXK8CuI6c5V6mnsj5RgcbOyZF20ja/YourQ66pDR8sa0jI9JOe6oUG3xxk10q
k/87X6Tso5owgLbqqqowR+MjnXZCRWOW6EwunmGk68LB0AA+MmmFPAgoTF2ryvTW
XHDFnqY/xfDIdU4iZOeYPheEAAxGrtB+S5A35KS5PoGw+PAxtut/nEwFKgb69cgR
eVq0aFxVnx6NrHDwNO5x8WJFxOKz+XfXQlhH/2EecHSLPFQR2xQkXIc7/xy6PdxK
HYUTMpFFSqcySeLhkEWLdxJYAlDqY976cGt60RbXF6M80xZo2pGn4+LzUrfr92q2
1TLnppYreHKDqr47bZdNNik6yOcx0l2Bj8bex9wIktT7dmMdQjtKxhA4XI4P7Lwo
R0hpHzTkVaxsARo+vwfhY7wwI72oNpESLU7HN4CFN+O/lryGpj2z7hPW6HVQkDWx
cwFDNFLmvPH4GwmDvDfxoMsUCkfnjj/nmlJQzkdPrH3usBG6lGPUETFC14B5+Tl/
3mG4QeeS+PGgpfl3v326gRIMotBz1lOyWMNaguh+i+wZcI5ZymOZUHL8HVyXDRzP
6pUDOuL3EoQEILw6IOiZ60hhLqaLE7UY0bS9MKLBoLLX/UWqNd18L2G2v0+7VnbZ
Ja1RvhnY5Sl98Vs8Lej3ID2dEFfx0pK90k3JRw4Vm0WHgLyAC2GoGZe46SU7PQLp
xo/fsewnYt5K/0RN+gsLcHzTjNxJElhQ76i4bDzEFJ6m+9KCKTSa+m4jmxTfjhbd
evnC0i0w1Fd23yTdMi+vfcJOfVhPxBIifsXN+lEbGJ17yh66Kngy1657bTihfWWW
x7K8WkM1bg/HvW0paHjQGiRo9uiJ3a7iY9TTG4YDdnkCEw1yOTGYWmjYrJXiE62H
paq4PnMtlN9jRqiN/llIeR9Ac5hTZixRhsaMW9kwIwxAjN8Ue9HwsZDugwq50k5v
/HjFUTxyAltBNmFws2QUaLB7fHo4snKMBVK566RPKXHIlPPj1bwA/8E9peoebMoS
klOt5ru7RoSLeJHd7Qf/9+qBCDVl2+h7qQQNhKVtwo5/v3Kkb6VDls9ieXws9Wlv
a2uQWdslalHgjsvBys+5icbV0JFKZsr29+fdiQWjP87TDSz/OwKinqMvoSDNFH+R
iyemqjnfCpvIQqaZy/RHXTbNdTHsEQoH1A+dZLjDyjmfvhjnmzQolWYXPecgYPR5
PulSp9vWAoFIoZ1jik+WHoveeiBK7WBHo0UnyBARwgNWp4PNMtk3BVlqNk+amY4B
FSGJRmE0TB7Ec9zR6s6J+spghWGq/XUTHz4zH7JtYHSGgDrHtCLauUvC+b/OLmqt
QA6/8PdpND6HLug0PsRgWbJYKcwiKRjYBSgLKOZlnsIjqD9sReqwVSLv//OOKILK
SudpX2pvqe2kCGj/wHAPo3bKc6o/L2jTJmf3GjzAI9HaqDgYnMxplZKa418RLzzd
FzsaCCINm4vssKfVGzYtzkWW9us2z0tD64LBjvoLK3qXp99/G4yg29lH29OL1xGK
QWHbiSNbPb42FYU7SbZuN2G7zdpDPW7AgPr+skGgb0PweWTDKdP/N8tbOLsyJD0u
TPEumy8afPFNTOPqSOWRugfv8420gBXcCbXvDojmdhtd/4PujufI9zB6NoSzxEa3
DWWUrm2ns4krY8cKgAoaBfZATnaZoTRpeTd+PdlTbNBMz20IhaQUWwEQJYJWEoNA
eaR1agy/SzegQdEZhPQ/Lzr+Rg3Q0r5v+pgwkyvy5PcPPeQKThSprxvQe/f+BkXu
3J9xF2zgJ1BbYWhwnxkdDsQMR0ZRwdRA8p5CO5QASnEaANqeEZ9ezb0ZswjBISxd
6O53+WAw5A5RWRNZOMVuEAkev+2NaY/ZglxBB78HXO5m3p2iY+W53FoUcXKaCvTP
WgoXYO/WKhjatg/0hVaL3N3233053QeDCkb95msD+Ht5JbfYucY9ruLyccUyjhcD
if6ksF71JqNSTS8hnEAMV2MArJvT6aVwoG71JebUqP1mWFf7VFLDnjngPjYgicRJ
7j/tiIBjKsGlm+fGQGxGorFzJ05fxf1oOTxRHNbOE6I1Rd4QrclbJHyLyTHUR7e4
ppX7xQR02BTjQWIvm03Tz81dTyfdinqgSIvObmOluOuVbc0IdZ301XhE3gGdqJlY
UHPnsINuQDnAyvqq2gflzl2Fe1ncQMuRy75aFxTSKNSNLL2mNg6rZPnphQ7RRZOA
ia4iGtvIliEEKffJ/t525AQSPK3ZJMtPkBuMVIm3StbamV41kW2hDxMCvXPwK+RF
kSgh1TkdfIORVcYk5UogQS4WQ4Nek81NkB9M5RTqSBbhkJ81cVxfuat2wnoreRD9
IdJN/7dtRLLppHbizQbskL+plR239+ly6+30t3lkUTEZA7hyfgQXwc8qyx7fth8/
SUVZj9ZxrVRhG+THEASCJ70BhgpNk/91SaPFNa5T4VNJzNEhJn+mtjLMVWlD0OMA
88NSeHdf96Udi3j9Z/rJXEOmMrhFiqDurM2UFN9xvL2xzD5Otl5lMZ9RL5vpDYzi
fF1DETN6YQkyKbM5A3QdUElkrs56JFYRmOnHD21FW33iGuoQl8QFE7aAq3RFVu8K
I9OWQfdxnzVFdVf8Ix524MpOjGNtM4m/QUN4M06l2QHC01MzRW0wCjRpzU4rjhk4
aH+hjLFqb8u1L6HvyLlndcH3Fsx6TYwY0u/WRk4++rVYV9O/aP9PhpEAS0FZuaOC
CtXMgo1OxkQOP9iuH83UN8IpsGendEsWLtZg2Z2FiNLGdIBcdWEhITx3PIJAGhPM
oT39mkTled17mCwrvs6FeKTK6acpfEtRyQu1vjqa4+gsZq04aCSm+BN2FfF0ltnT
Qy5PJAKJVA+KTFp032MEQW43AcxyNpGANbrDnCOJ5dgLCxulyKxozTzhHc6tmacH
0Xa+fygswUnYo9M/Pvc2gkgqXzr+Ljd2Xv7K7OAnBUdA12Diu+LeMTM075WiLrPo
errzd8X7nEf3pfhLKxcNNPBSJc4P2X0nuc/SYlyl24ZeA/d7a4VYCtcmpMa6HvOF
wSN1YH5/H6sGbJqe2HmsANj1s11AbbQ9/+MfpzupJVdzEq4VYECnIE84go86ndW8
8s5nu6Xe3+wEjSlrDKmhhQszaobqNlr3QUW37k0SEqKLRgt7BSJ0vNOp7Z7lXiA0
080S6QDhfm7TBjJjhN/Vpbv/Y/YfCl1SrcYC3Ebu4ElfJzpCktJ+PPJw/Lr/YbvO
YP9AW1cSMmulRM7gwREGICyrG/rOLqmVpME5Aazk133UaDx6HExSuoayJDcQ0cB9
JyUK3Efs73lAMPjtmY1vipD4i9dzVjs6jknB8OoWkAnCqcrRUk/QyauhnnyxgHb1
K5EZ+83cJwvkdX+pchk053i1xbP9h+3NM1x8b0OplQ+01U51U0Jn8M8TkUbhoU5p
TvIMgf5f80iLI1LopAuJwijIrQ0RiQuhicrfjKwCMCy3SUWtYjLcSnjSovuk0g1v
lKbtvWzYAedKaxc1hufEFatCBcR7xbCr4ZFA5UJEDRuXt8syY+bfyrFVpk2NVPag
PCRXmcIlAwAHNxKuo5davOqPF8GaeDixql332jJNVf1YQIySuQe32A/OxRfzmfC+
b/6wB5gTckusb7nPhXsfDahjLu0A7T4wr3G++eoMsRmjL/8vCxd4ocECfnb/7Kkg
MGa4NJHAe7509gyXRY+nvwMrlUu7icHjLnpoK59WF0rNqbxlM+OzpCHNomTCVzwx
hvEL/H6xRBOhYRtL75AmArqH+IfjQW5D8zZ8va6qayxFTToO2DYSMN/gtHF5RsjZ
PjClSnGTJRWAB/RRLm6f85GAcZECp402PJzhCa9sKg4EtvBZLdV0KkYqFp2Y+Owr
0K3YtADyHN8BBxJc6NOavMQ+zQ8An6Fj5CxuQkLxGznUczVDLaJEe/IGr4+fPpVC
xUsFeY+okMeIKoWTRjFyLkl8PL2CodOvGEU+GN5m7AGCIgywC9qEY7U+CFBOhz/y
Rv+vDrIyxUJ/zd8DNvZSOXIZt8/9nTvot84eD3ZNdNJcW5ZoZTsWFAnfyBRv+3pY
oJZjBisPiCpW8TcJIm/dedC3Ad8psI1wkAvFcFUq3JiOsqF03WF7VeOsvTjFQ+Sv
NYD0sxVvvbgDvJo0mlwHi3Y+KK8UF3oHhjcb8w3WGSye20sYWGc+HOEwsZ5Ji4cu
n4SlY/ASlHUzey1OhTkZa8MhMSCosXl2Hd5aNjLM/rXffwm1NgzyaGb3o2xZZ+BG
O4ev3GlgeW99KlDCuO8dA1Zv3+9Hg0wiyKUb1Oof7YhN/sQ+k9d4H2JoCtI4cuVD
slzZDt3W6UkXrVcNrq7lbr0829O2iYIYOT7C2qNw1KNZSmkoforOzX9SsnezlPfn
AmUSzsBK8VD9LvXhqO6uMbjnwAB6Mdar3xInN7QMeJvp3GxRM+KuxbuIENPGuu1k
4S5uJ9FD+zzE9Mps3duTNS50wfvhUEAklQdGS6SO2XmkNMY6HOmdX8+SRrkxwTp/
iMjtwmg3l1pTyhGcLfXCQ0wLrYP8fwIYBgSwNUdLbOh+MZyqdQLezp6QY+z3g8vM
QxcvXP4qXC65z0oPTQtB3w374NUbzE1oYsxX0kPMgz/jv16Uno3f6rX41e/Gn0fn
lDm/vHPv6tmMLvTIAtxm+PNNhg8RJAKyVn1uv8SAIv3VRgN7pZ7LBF0QN7A8g073
ix/gZ87Avw6Rq5m7bocBZQeyPyd9spddttIF2W32g+LSXEPoUIgiuCD6W8LHVTlx
Ixa/OhZwwq+f6aYgn8CDQ09bq59B9ZycP66znKAXdIZSKnTj3GdqBY47W0LI2Oit
zKCuLMCH3ikLvhVGdFPiieu1fWgQEuJN67NgQi4hk5jyVgwcjIFdhtDVt48lytKi
gUaZYGLeui4EkPdi626+Gvx7OEHwL4nf1eWh9zqMaNOS9qTTwcQ3SerKA/UsazDg
EN6gwAQivrdyMh0Svr3H8akVT5YcCZeUJWitznyfWnxug6FoBvU9+QSAUUG5kIHy
7y3Zhqd8ZkLT26OsCUjysXc19Q6XGvwd1xcD7FR5MzhWHUvhZbgkGcIm8h6toK5p
XwO4pFJPUzh+YOp366VhR0QO29Jv50nv2yOd8rma4iI7Ih7lcO+u9fk3l5WSPsuV
sIME9exhuxf5kMaqKWHfuGu/4yphlXW8tIX9vGNSkf9D5zkUsStwoC2mEy+Ei/pA
5odYsqkbX9GJjgXF1vJ2md3rUCaX4TVFNLVeAHQzaQ57vx30R3t8I22f2rXNGE44
FYjCmFS6ScJmJIwBDr6RTO0BSSmcW15/M7qKPOZbiVke0XU79O4fp/lC2/zLY1lD
c7ax3l9d4hsFk7fyh0cCekGGbl+oK8wfnB5NrRlxiG46Gdn0lVTidIC2i2hBZyme
SrDdVhGjJIqBT4JAR5n2YNVJJTN2s31+nrh/DKO360mqc1Bvpv7QyYHGnTtC94FM
I9VKL6pEpifBCVC/Y5eEpFW50qISsXNAouCTM5pO5as1ElWV46eLNghJwadtw612
QzlKwNbugwu18jIhDmZ567eoF9GSDNfRU4i3kFJ2WFqoJrzKGEme/4O1ONPusFfh
AcVDCMv1fnMeJWA2SFP07BlmLP7s7Q0WryLgVwAhhG13gwJsTIqsxOYVOZrp6otZ
9beHBNM0E2lOIpLWucGSPiK41HQTBahrLU7lm4WnZHuP2D8QVamR7hdRskHDWuXi
HdGcJbJ0dSbG6PFXf4W5vldhxlbe1TLPIIZV9PRJBtxDbNQVmS43/yH7EImHXYlR
H9sDkXslIc+RY52U9gbm3sGmWErnt14dA8kvchdnpN8pFCsW7SzBkz4/Q2TOmE59
og24wEk9YTcFFx8Fd+4L/tdmbdh0/vfzhVO/DeegWJNiiN2i0BxqhWdtVDcECFHc
nkhAWPtI12jyy4K2Z0QE13Jr1onl2D6Lr7NLVJMhAWj3TD5j4mgEBTnGcApbd/fb
zmMA7ji5XmO7Qvl/wmXPslJ8Nf63XxGr5QHLdjAng8ALKl6i3ATZ9g8TUONZa6CB
0Gb81msIiMzAkyaylOEqA20GXKLeg3F67QaecjzlXpKqvGnm2vMFBZENhP4pUlrl
mDgPPAiAb+Gky8jq/i7uslFpFCgspCgJuLbHbTZYoAmZ1jduX9VuEZydjxCzn8DE
kh/ncA1rOv2CDYe+OdMj2uUjNHQB63egJzPlcTbrpWEN7wcmen3CrZLe1SeOWDBD
7x2QyychpkdLmJ+qCLkjIRno4K/riMJmcEUXQEJEqMTVNany1/dltr2jtMy5pgUs
atCQfdbOFHVZwSrhHXJv0zBOqkC9i24G0sijvDB7M8ptj3r/xLdftkUmoHYvvQTA
qJCdZg6G6xa0M0GoEU2v8azI7feI4jeGBTmzfBT7mLdRFHDyhDrh02MzwXTwL/Nz
vVRf+vNJP7Gydy4ujb5vChm7V+0CL4XjpfXlcSHkIoUdbGnt0gQ8Zq3cTKk29540
SJmNYXMCaXX+09+BfqqatqQuRrcSwlmlSMROSGGRl7JWs9MoXhpr1kb18+xuOKsx
eZU0+iaVXWPSIaXOG52Jd/+muklW4Sxup2+A00Qt0dfqvz9INsNE9nKWgZGsaeNL
IGJc9CeyV0jpP6z2I4d/PNdc/9CvQqc29yFQv+vB4I5k9gKoSKCSANlGoClpkdCF
zyGWgTWCav8VxLa9tN+E4GtQLReNIWb4EsZ5GahKJluMVJcKGz9HZ8nlbydrzW8g
92Zh892pdhPT/lniJjlqpI77RnoWl9glQrxASHw7/cxYfPIYkfLJ2mT1bZjJ822o
u3aV0RCVc/9wKKPt2Rq9ZQowt5opyMIlG4eB2oxdZHlQlsKelnnZmfvyMkFNrypN
AmyBnaaYPYKidnvu0kigtOWdTB9HE/sLALhILXaKNNO5Z7Jv7tx8ie3INZSAB3S/
JXv9sEivFgHEOZYvssZ3NUy4ZKtl68XG/x7gU+ygg9iNDPdMPQDIqj9l4qyN8NQv
J7m0FCzwIfFh3VyCq8802LJbhBAqb8F0q2J96y1xi4U+Rj2qFINwW83GrPQIdu6A
MR2euHtZ+IMRcLbhFMpuNiHGmhcLxCojjrmKTgEIA7FNi9ss+phB62eYWWZW+FyD
s9KgJgaCq8z94XBJfhs8jNsN20eGvHsDmBjj6nwJSowcYEMkoNeZgRoQAD1HzoiP
Dd1Q+qE/nUXueBFH8H/Q6AnFRN0EPkTAwQVbWp22bVy8ANbkw8y+W6QV0t5uYZMX
z4F9Ae0row6WQr5p5GjBJFlZ0Gk25pPXzDvsLMG4zXyXnqudvD8HO6dBPzhT9DEZ
ImlqIgXETyCk7UVCQ12dYcwwnHyh2GEmJ650JUTokPl8K1M/5ZVVRfSQKS38luhZ
QSRfFVExK9X4Cb7nyfnuMzUwzRDrIL0oss8hh4Y8Jd/GtPghVxl1Pt5noDauoUiv
xUHK6Gi9wFoQGpW2OYzJmSWZqEv9FzK9kxgnH0Q2KLpo0rVUUJriZc3Aunkf4Oy4
IvD9biRQPoVcQTuyrOrrcL56yNzGO17fKyZ7zFNdqqEE1ClYq81MMo4+1KTRU+Ht
OEUvIGxsRQU5rMAX1qc5NsqtTzEzl686OBHk220cS7Yx5wJPObGFeL06fHhQFJNy
bO5UXNsFKEs/Wy83qhm8SNs2GjBf69pX8GVOSDHJ2Qu8TjvUNK2q+LCF0nyklPtL
9QZyrufKtr10NtA4Yi87L2cfSo0EEXj0lFFLfKqt7jN8Tnz3Ctz8lqKdYhF+Y5/F
8EHO9mlxqZKI6XkuhGlpBuq8eDAWRTHYZUASStQH1tRRzu4WE1nhfIJt/rsEu+xe
5xixjLkzUmlDioQIdNyHL3CbLZVDkXa3eRk+6HrnbJrVbbAATCCtm0kJrTkZO95u
S9m+PIf2G9FZnfi8DbrbUWgflJgsL0jhQ6jMYLTb96yjqRbXD4em+jzoJRfB4EKA
5tLAecVrW81dC6XS6aXdQx0KJsf8huJGmmeQhSbMXaXwjWIkfBw1uH74mQzS57kQ
m0UmPgDYY5SoYF+b+Q5f6annxaN+9hxFnF1/BpoS/oaD1gkXQFq//9hJviKOET0f
RRtekR8w3ufifjV5TNyDrnQiRNaVanjpEzYDZCQrizz6wHQrW+E5LrQiHO/5oPaH
2bFu5+Y3Ur8m66FFZhJZp8cI9iJyMzcbxreNX5gNqhTgGnqchLJv2aBu6K5wzDra
NlzB/LYAe6KbF3iNAFsx71vEFDMSQ772ya8xEjAtd4hkjzVF3HG6QW/Fx0NKQzV7
6FnC/c5KdPw+485c/r3RhM5FEp7WQkNcB06DCbiD1XRCvGGMhMzAXyTq+jjU91YM
nq1YLkF5NfAS2sv0K9YbuQCaUDX5ZZR+y2+xsT0VXEyBcflqhRySEruFAL09UC7/
jI7jN1VtCsTMy1Sxk+ATS4t/9O46IW+tTdzOOTuRwPiWf8LZLEE8Xzn/BzhATwzH
epnm0/tO2cqMiRUQnUbL8pDxywWAuU9RSgYlMtMvLbKVa6+UE+CtNmu+mncV/sKh
oV9tkxQTymY6M3x3Uh4t1nL5uBtOJiAYaxUUeLj9nrVNsI1n9rqTOvR4i0LEBF5c
ZsaQX/k9/IuLO8BQ9YysAMjz0Xce+yF3Rl/xVv7w/1wzLTmcpVnhSNEmbR6PZvRm
LAzLPuuo7kZ5cNvb7vjuXwZvmthaJU97fPHQcpE7L3pc2bJrw4uQ5lTBdFR0o8f2
x0moYpwf8eFt2eJWgho3m2G//bW3jTHIAjJyK73lu9+qY3EfrCz16F76948DyBf3
sz/rrGVIPOY2HLNwS9Wca4WShnGzd4ZDIFtQlCsEvpPNPYN0mPr21k8gJj8gbwZg
XUUKecAmiu2ZcKqK5BUKozFNqwp9SWbUPRDQnHa0TkV+F8pkvDyoQMxWH/zCUno2
9BNupZNl5IiK4RXcU8AcD4DD/nZEnqlzPC+sS39dxhjTzCCWtvihi2C8YaVFKmRb
TOocKQE0DVp63S2DwqSGZxMNUia+Xs9/BhX8Hti5ex8JFPN1d70sDeH8SqhYVyKM
zH91gwfEuzuSihVm++SkwW4QO8/qCmKQlOP9/4Zv8W5ZLYJ8D5NbnBebpMdfYdOE
nQGtU1asuo/WnhvGp3frgMacBkCvMdkmXQP2fjDmWTIDqZj63EklIg/ObKQWnXki
CXDmbWIdSa31aEIhvgneCUnvv/Z4PH0Z+iT19EeAYFS841Fim6hyt59YElaAzv8F
SW6nPnLjb3RA4Of3OOs8NI3cbFa/apd99ZivRC2jXT2LWoYhcsKU1goLnbwZhH9z
SBMVF6zH8iRBAd+/lat6iG9K7pz6/St76qbv/sOYePTMP1k0050wpqhJeUvYwuQt
Msk3a2CyB8XJ3KuxfLOn/1MPzvpX9jrT9BhAkjEuNuUlzRM9TvZf4w2GJblxfn1V
Oxf+da9qQ26aLCaaKLGUA7Z/ZCb8EJg32Pi5Hd5ykuf+zZ6AThZInSNsArAwhXK6
+s6zuoKJEiJm2PYuIL6hGizop0efr7JVv6D7KWqBNp5wtbMGW5etGaEgKWwCfePk
Mh/o6hQBz+hg6cz9abcbM55AzLvujt9cbBUTXbgjgM23qX0GOTXub039TKgd74p0
J044PLudaO8MtEIPFKJuJSjfAt7s8plgahu/U4GVBqCzb2/wsjQSSuThFiin0SNB
r9OcYZVMfAKks/HZR8tM6WlJy9byMCwRbSu3BxLVEwRAUmFBwo89nMJy6tlVfh/c
FqTGB96JkWGSgjSsMjDxFXVIGAXnMfYIHpKzHfOwEhQVowsvTsV7pP015IRnSH+2
7KC8HqmBXLiFzhKHVGgOvc2LGToyc4eAVqSLyih5jP0tkPy2Lnf5o/Hq6I4yxp0Q
sG7fZE2UikrWeshdmix10QPQmlZ0kVEsdQNN6BML+fyyGPEhwViVDicZMuHed6Wu
4wxUj7BUL4czC8GXQ573aExNKLJduR2RLtUWUBL9V+nUNvq3Ar03QSo9rZxzTw9J
KyaVVU88lVJCUtJXK9lW2XOKkjMdRDM+eLw8CscvJaerTnL8WYt/AKJbOy/cNPtH
xPU+gJShn/z8XB6/i5z5hBPksh31LI/sULLaiEFJzVnZwGBlSMwSQ5lIuAYU96y0
rDDlf8Owp8gz6uoyaT2T8EpTUdrSgC8QXp4mICPUUq6yhOoolTDJy2/6SGfdl6e+
6J/klfUGs2teCP9jShy+U0d3lzkhrnmEIYGdknhaZ2LgdSOF5GmC3hz+lmc/2Naq
RmkKLl2RVBQPDCLICj/h+s+/rfXcYFSt6z3kwd5czFs=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
KB4ksH83clXJb23qUaglabSvcPx4G/oNMuSEbv2yfETOHp5y9NoKWs8vxedBDKFD
gHIopcqFIZDRixgzDbryipcZgO7siLP/+zaclaFDsH0hNSGKYU1pjTi3DB+Exxyq
ckscR2ITBMd8p5P0VwdPNbWp5e1fa4gQ/pge2vIIecHVDVjURnMW6oxNfYTOfFym
AeNZq034N9Wm0zdtAz0okmpOqhElUcjl4u1edCF8z+1HOgG+Cw6IhA1WE9/F9tQ5
4JQQkjCtg53uweSoW2fBoGfm91qxyb8Muk5oRgYhldyFFTHFrxrEE4T1TU54b6Id
hVSBdSjNZbWTyPU4PELZ+Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
d9nDpEWDh1mH7dP7gLGYh3eblhKuul8ys2kY6sO+eJ+GZLkPi3NauyekZjVjIxH8
SDz1nbgPJH46s4D4z5pHjnr1i+PoXs0luo6DlcmZxfCWFQOnBun5vwztZYflggEE
QlTSJYGkWDM28MoZjB0jq0hh8/+03NtNxKR1jOWpHoyzNz6nVioG998piNtWy45E
1SP/4SFv/8qzUDFGi8FF1ZS99/uUur0IybmZohg6mLS4YK5B6TFHQGGmmluSHm1C
hPsAIVu67pvnaCmA7JD/sM+/x9X0pnSROrwajFVPXIGbgpIQkUM3VlIZ4+3QXyvt
AYxGdNkF7hRORYI3+lf9MW0F0WUy+WMR2XDusQi38rywVPf6QCPPuqzGRjcxrD21
sba4ofGkMmeBqdHyNmYoWvVuJ1np0JcmAiK4E8uR2SFLQmecItFbue03HrnFCFPU
pWoGV8wuU2bB0jEm0JnXyD5iPcv/kKeErkEErg1Bpq3YyGqqhirXAvHiMlfNexv7
gQmf2PfRDJ2Y7aNmLmH/ITmrz55OwkO5F7NHsf8p/Fowf+tuHATd4LHbtrBD5/Ug
0zAAToD8TQxyOIgmvLsgE+Clfon5mIjPxd2pYLYxdM16FKmqh9sfGTMvcRz2Rcsz
rUP1LeqrDKlMq8yeqkZ9RBqtrTBFgPlrInvDZScTQz/4BE6jGgeIAbxMy/Thqg4c
Jix6ge/okUz5e44JeTJe1TkT//N2H4PTRQnKEIw0lmLj1qmg+PDaajtQkINHA5kR
gsB1mdHEGhN9Osrfnh4Qgoh+eSOl9Dw9WMeKfA5vnYlrVRejPez3sLqcLYpJhqUC
fA+gduDGOTs/Z+cFZgcdkPIvNyJWOLpmljnAR8ZZa5aKkK06MLZ01zlOopNi/RQ6
0QryyFCuf6xBvLodFqbQ1tjWjrn6KL7VjFhRcI2oSJVOJ3Pd+rBn5t+6bzBDLaCB
WnZk/PpukJ1u/LXyiZyw9NQ5BNjqat8GzeRZUM/UCaHq6T2C56ibRhwq55t74/nk
M9JTiPgIbulglea09zwM9p/gYhaevslCfEFJmD36wnBJu1e55A2rvDjAC06Z/SEp
JXLmDpPqYYK0trOO91ZiCd467rHbnrfockgnvaXPYAIWE+b1JmpDwWvCGwdQ93FB
Zc4SPYoNIlUho9DV/i/EKrfhSYKkqkya5xiH2DmqPlOmrHcEHHMdrsLN/YKG8Ciq
CcbN5I5Clo1gPIr9e0+4w6qPoE4iGTpbx5bqMM5pC3sMNBAOzO7a4PvLtM9YIPpD
qbsu20Bj9y8jAYx4nEnwUkdiotNRm2cCy+e2jhCVSEYBG4DQFEjCTxQRm+cIuwba
ddRraObmoSoR4i0EmpXOm3oNnDuMjW8Mdo6Pan/Fto8yXnSP570jGzDNe64LACHU
uMcgvGufsakgpolvzi0m1HG0nsCEQ3w2dD6mPiK9dmN8nljw3Jb3ht/q5UOdgeJF
3XkW7K3XTplfwc9dSukW6JxHLMl0Zp8fS4Pgx53LujMEOakcRryf2MZv+VFvMEiQ
CA6zydE30f6g3Mh6obLSzgQbarQIbV+WyzrIQ5kTCr2J4qaXT8wwd6w67IZp/QwJ
IG/RK66klq0ntrsUzeac8M9bf+HsfeX5e5+0RRWScM50350vdKUOyTXuL2QWmsNm
gKv+GKVfNKxKgtE8ayy5iQkNNARS2x5ZECAcwicK8GEGX+nG0+hwjd8QolvkhTFH
OwhkbRUHzTxfY9VJe0IuzWwC2vBQTBFbu6kmnSH2sTi0nXqriHra3w7J4hsFUKMw
/bvh40N2QOQaGPCdcDsRObRsZ6JK4LNrayUeIhPKrxn4TcVOYicoOGWbjR0K8JC8
xR+m6yI3olgUswTgldgyjOwn3/Y4TAoaKYnjMQVbGa0nQH6GIfZBheNlI+22Hh3m
yUYFw1P3QUKwYIOMeDQPPexuWyrNWw9ijSWdpV+wwb+aiAjutaDL1CaMShbEO7xs
bbFm3DLbXocPuq3qGg+x2P5IwtlrYa8jDFel/bf4fv3BcMkX2I2xOoOnK9qXmrBq
nNsitrNZd+V2EMv+ig5j89lZYz4dW692OqXRHZbsdFml9AYMNXhS16fOWumMJW4K
Qg/Ew0idxHe9nN8EfNZLVN9Y57j698Rd+h+VRoc3IYejOCR0O+/qa1zYYFefdxjd
jWLH7uJGPx6h9aXNLWEy/WGgRinpBcbQIAZ3Vq1/TxN3uW4YcjnRd9xL8oIqYuWM
OYhdWgv1XPbBv14fJrQbcBXXLXorgPi3hGoRpHPONmvdtWaLOq+iE5/nibODW7hZ
5cOqybB5zmJOZrmh+vAUOKCLw4Jn5KEOngrO9bGFqsV1nzxKKusuZFYgcB6x2I1H
eiRhtZQaYl0464uFJkyo6rcoG162bMk7dZ0lsZi5AwNIgh6wVhpGEU11Gbio2MyI
SdcJitcEuKqHYPSbNhebCgjpbTMvX5SnyCu6tNYICpInlVi7HNnm8Lt3TyyTLL+y
1vg7rFdaqtY2S6QYBhH+zRTsnY6NJ1YZKT9LgKnvNUavd8WRml/z0er9CWUMLl4+
s5RBC7vYHACz1OhnFLCilCPPWXVoyF/JzObQ+Ak0RWpnGWVM+Okk4ZAxpgDThObl
JxOOd6WFlmmAcyJQG+fc4Ix096Mg17J4yRB24eWzVsUwF92ErqMxLSh+boD9lMrV
MFJyAu2QnRsTe/sjvNcb/dnLnwObOtun5Lsft9Bl7mONBsQo0CaYKlZDrem7Ua2n
Bs3O9SeLHXpUt7MAaX+tCbzrO2YLkXq1q0mAWuQLhVBPtOAmj2fb4dPjThcVTIHv
/KBgDr+4JcXT3muwsPFHHJOC5scUx+3aVKUQU8GDbHyx3h9q2UHhPPRsw3U6Ch/l
PCmZwbiD4sFhDkgwcMP1Y7nLryfpDVFilSEKk+L3es2aM6RGZJ2cwV80pVcVy35F
CSw5je/oTktd/TVDwqQO0V6dImOANsVPvqig8msRTYIwWm0sx1tRetp1wkRlP4Qt
puwdbvZw0yLvl2KQUIRZYrmXGzNypsI4MuPb2lT1EjeuSaPBKmzXfgNY4cqXJ3sC
C5ZQ1uU5pxP9NQw8BOsveoAIIy5HpUIWJDGjgz21vUWfDVCjcu1K2dsYjx9yoBD4
A1Hsg+Je6fwczlOmGsDvUxGmeTdVDbUDPcJLkb3StCmSJ+3qOf2N4Z0cLOCU93jj
foSW37w9KNvRKIR9imLSevnFYUhs4YvmiEMAOjg7cQq4ea7ipDsF/omonSEmCAGo
bYs5ZUpi+Z1LeCm6jCdLon5udKmZ1j8bFF2N2T9syC5ByTtNJkrUUfw2jxDHbScl
dGJ5hwEA2e7g0dUSUU38JGDkP0xfsaT05tFeYZVpBmRAnMT2BwMuslGt5LgXOJei
U18+nMEuhwuRI0gAW7+ORCBuf1AAZbX60v0XV1MCYufqIy8IusMYvTkn182bDVd3
RcdluLoEcrm0YsNuGBnttbZXS6xX2r54crenJYHfH6nIBrDZj7XDU8tbRCge6mwy
cZKX76Ig8553ZNI9Ld/OhcgZQCa8omfmrn88/5dkMJygTEHz1WiHWQS4yIcTuWni
sA0SCEMQU9HiFlzPZlm1sZKFobkBoG6vVcKBd3Ryilz2U2ulhClNdOn1YGKalBMj
2uha84wt2+QUdvaIq7KP5//YWdH2zOs5w/LFCUg0oO2tWrL+9pGT3cL3SEORVRyu
Cry3j8+P7RiCf5ANkMuu5xi5kRUg4pOh0IwJB4C+Kzu+jD1E832EuDqR8hat41YI
BKLQlew6BXW58cC8wBpyQKwNTiey7JuqxQJIVf3dPHBQ2A5EcB0tofREsZkbi8Fp
ufT2cSDvZrdKIWy2lSy+ehlXm0zx5+a5ejuC+q8pJnmzccfNROqAJKpvIub+076Z
xl+PRLG+D0zcG05oNbWquyQ+mFWs2X7NyfVaGhQP+Qxp6dYpSMQtfv13w7gObuD2
+loXZwqu6nOrEJziRdHKsONbOnLNwbOWg6MINa3+Ypz+5M0lgoiqhBvIJOFrO69G
whDTm+9I3SPeaOdoG3Kx/luoF9X7ZcFqPxkVu2Z8pgIScQgPzzHaoiC3Ko9vW32t
VBmgneyTccBTUlEtW1iqHZcUmW45I29TEBFe54TN6yjM+AeyZMDyJzzjHkAUuin/
5L5g3Ouhn9FjSBG8y+xXJAKYp2vw6uSsp4L3hTSkhtkJLVrdjLRE/zSjmaB6ZcmA
+PQYNQJ3PG139qUyCgG0QrLsw0MyhrFbBCUQuEK3C8hvqE8O3vo8pgpDfCHe5Qez
FCFnER9mP89fiWxFaBdk9NpGrHbpagkvdSmYE5oXE5kKApr91ipOR42U2rSs5ABz
NvmVDOO2KdxOyg3YI9a1GYswIzeN66TVTebLxWTyciv0DA0XqSXXq9LFlOKcBepC
ljDHsGFPfflyjlzZpMNxOrH2FMBJPLoK73ANiB0Vuq7zMlDt1oY2ObQtCc/Aj6LP
MgQAQvyFXR24+02XFlelUJJIhKQ5iTXRnPlQ2XZeZwIlR4gwXahiUHn2orLvtdZv
aJaMbGG6j0Xcjt+sa2jVLBy2brLZfgTgkaHQJ8vBdcsF691jHO/gIRJLC47bmSsc
hpyzdUBQUlxkdjaoTu3F3heAyhSTTfXtNoRo6sKEX2cU6qN2N/oxoPGc0vUMZ2ua
LSFIquCNqNOe5yiV5g5nJ/pjSfkrFK7PtI8haEXgdb6R3Gk2RAGdnmHh/XNkjxyE
ob+QZEKLS2vBepoNWLIRAHpvfVUckyYHC/9e7sS8Snu7J3csKQRRaqCC/fW/3nlx
SzN+BPWFOpUDJz8oCsTNJn2nWl7fV6AVv2A40Ybohiz3V6OB29A6DnMqbyEEmGDJ
0jayJAsoV8ONn3iGkcyzeWboYZ3nuWQ7UombURkq4aP5twRwbZnBPesv84qBhbxy
GquODYqdPWZaeefc99/3QG9R73uxo/1TIu4bsqW8G2k3o/POB4KH9yKURec3yS20
ckbi2XfgLH32DvOqNepFc7AmkxFB7okWWicZDR6zaxq0GiBTsYxL6ZtmyKTSfalf
X6sy77OhV/FLfpaMlxoOVDcJKGBbSFd8DOMEfmpFqhWFeMWIkVvPAXB9lssjVSqg
VXzC6KGpkS5map2sq0LvQin6ghSoJx0A+UJ5QzmcVswZ4cNmzLwbwY01TFg9NS9Q
6S8lKaITbzYnF5s+YECQKWaBcauQTfFZGrD/8Ie+RxkT51RdEIyIONH4QpUbBXuq
HZLKCZQuElHGQLPfvyGHP4HkaXg8CrBxxPOzKGzyGJrILKSzEF+PJTqNHKkaIsln
qGozLsuDbDE7LrNsIMxOoZH0AFqMGg4+4WrUjf1rf+zVYdOWv3Cvnww13ekxuQrb
mK1cuuKclyKW/NLw0ZXEBJqgQZNH9P7GE2gv7akeyCdZKFVb8jzBI7S0o9z/ei8l
/aYVaDcyuxvbwJwyeGKiOKzse0Ff++aQViHKKVWy6elVlyXG0OcXLgbGKce3UOVs
UWkVrXyphyatJFwCjJCKeMzuExd+JLcsnleZ5t2idWtLqfaq+kaPNfzk744d2bQ7
8V7uS++WDQFQiCLqoRMeXqX5ZvGp/CSb1ujlodKpmJeAKWgagbjUG4+92kv7/IEw
UBdTD5CSz4qWAypmoTFympVUd4FPSkqdJc6/pTtRZXiGDs63ElIMehIO4CGf+F4t
kQkX/Bg9GbnltZKWzzlNer6OBsqBgnHCPHCpzh2dSBlU/c2JNdACK28BTlquoVlE
mER6LuGWJp2GBKMvRVB/jytJsjNSHGvRuSvIZSISitRqx/2LrG+6U4CpKGj893mD
SlWDso6uGC98uV+prtfuJN8TtEfmnQ/b6/kpHHfzDu8IYgAeXMXdFUQR9gDyBMDW
Fwa9mqDMVJ7WVjCJ5JejfstYz5HsGMa037VsaKzA07qmoN2dhANdgWEVmepWEXDw
4ulEhO4n40Dnjp73o//DbfDkoSMd/8eN1/Mnux35HL3d4ST/ipK7YNzU4/wpXAmi
18nsLyPvNlEWf5ZIxLXJNgdDHRDbEEqsq3cMv2WpzDXnOIFZUPnA1snZx0DsHPgs
y4DsfSG2PuNkAFQ5mmMGpnS/o1U3MybGbSLhAk6xSmQD0X+85kbtp7M4aInrHCno
yr9Bwwyhkkf8D2YlCMuDyQ40V8Reb0kVNlU6iHXJ/qeiwCPfmtYfb7d6W/fdd2r1
Tozqnc+WxRcLSvBHAFNXOQp5ZLA7sxepO/eNHpKKkDjMHSeoXrnknaES5o0PpUIQ
MzqiLsHVMoav3aHrzqF7d16NSauTZ9hMANB2MUIsT5Wg5PP/yVBDVCPwi70vti92
lypuorW3v/qCBy7Ega6+NY50G6+XpWi72+vQvXIrzSy90R3u1qAvp95Vy5vymBTK
Qi9uwEZlO///UvDRnoY3JNzC2f7HgA6jJEnVYs+5WAWhjUDudkFGD2fncNeNS8yu
kfDVZnmnMjUICEDg8MzqZHXLcnwxDSWCmghZg7+4ZU5bvNon8baP23B2C3X6ZHOM
njHBXHKHlgaMuEKjoEPfDfPJfmP7beVgq626+Vs1Qt79po1xcYmdo/i8Rg4Tj5Nj
MZrcN5G4L8MZo/VNHelxyxZhZozVtdgfD7wLAmAiqzOHHV/XV6jVRgqFEuzmCnL8
9sQhpMa2mkbXTqnwkpxmm6Yn+0AlglZPjjuvOOS6Mkj0O2Xn+atuF33Q+GZMfdd+
zE7xWZtw2dpzYZFgMijguv25+H3KZ5Y1+8FooGzHRYK1DJSDhLOC4xcF5FQG/tbQ
EW0Jf1omttgS1mxyo9xVJT29fD519ZwvY7E6vGnygyJgGR3NsvFOYkZPNfY5geK9
wB0akvneNJMBX9hdIuDyM3RRtykfrk8WuXam/BxCmIvI0l8fYy7JCqKTV4pFFaAn
cMtlrKgHVCU0Rw4H+U6Xlraa6jfCSYE5V9dxVxcWK+Y92gRnyovwo0XgMRKPnzcr
c0kavFpg7/J4GfpBYCLzywbe1fIRryeEPtDrLSIkvsK8SXnoWfGs/QA7D5Mi48BH
yhT9y+mNihR/ehY/rgdCumZ428EmzOsRlztI7gIJcZ9gFAk+3Xrmhk/Tv18M8XGv
yb9/Lwn0Oy2FSL0ch5rbkc+v5U9j70c1x6UubDArKapaWzEpPmdgUuvrw620NWIe
EExYMxtLgf3Rh1x6o7BEYr8Jo/6ovpK2Ngky0ZRNuw6k2JGf3DDTHzcMoCV1FyQf
8WDsjqJieeW9avLfHdWvjNlmpuLRruRO4lCssSDzAbLX+6tNhDBC/iEc6CHZ9dg7
nOPNqiwJ7u4sSrX80FX8VdOHF3KNzsLJ4OXJIRACWndza92JdInnF4x3DA0Zqr+R
0bWdg6gcOu2QLUj9ohMddGHKBSMM7/05GYfbIjbowoMXkp4SYGtOtdPWz/20Bn8P
BceR+fQ85EDjYgCT1EpJieXxJiUBfhgmFB9Ahzl7zXAkXGzzamwdXP2FMfjLRl8K
Pzt5JHbkvHXXNgwlogEf6a+bNJ96N4H2zg4dwB2XS4yFmMVbA/wpVmXhfUhF9Qxl
t+N0tCSofxpDqqV1Jtnvq4nAKr2G0lmBlk3R+QSH6tF7Mr4rP+VMQXxLPET47re0
+kclajByVu6TUQ9D/GJaueyy4VLrRtAtm7VWb9FLlXseA6Igh7RQYYifnEWr76zM
QkNW/l0G3m8O1HSfbksGPWrvrfXKmKaqrqrnYGvbCYeVhSyt6fxaClP2Gxn4Y8i+
7sP7Vx1mAXZTEm955y53WQ7XngkbTtrZTHoEgkJPHewBVLVdnRJtoG71bw7BIGoT
wQMlyxeKNDzro0wlhBiR1qsbvZ2/zhaDXfGsxdpQQOmRk/TvWgKFZqPN6yVw4a7I
ojxIqKKB/iGqMmhLsBp40ei79OZt7WjVG49XkBV+YarfsJc+B8HfcrJW4pNBY4RJ
KnFZzJimEsjwGo3ZqlE0FccCZaJZeGGnGKuqdusgNSA4r0KaTts85uak1VjNPHxC
rg4ZUtM5E19jWLUeGn93wEV3+kxjxzzUEmSbgGqfKYtNgoUdJgEIL76/lBTtRVvS
4N/dplZBaGFgCWxEqKOVh/nElfuMf2QKYTRP5ztXbhvA2FgeebWU+t811BAGIWYt
2Qu1vW/OYc3shR5+IiMlW0UuUk68QjaFuw1kz9Ri+hdzBhwQVG8ovaRYrpYh6Zcy
V7tqR7u7X//TnYcaqmqQG97ZW3O8+vIHhMoVb54uo1pbyrQpNW5L2EQEYnoH/jq2
8bHML6CBl+UGOKO0oz4m3qudtEgTsSc9/oRp7LOEjLvcV1LlhuqXEKldGRHFY0Vi
Q49DKDyZ08t1DRWvatDQLMuvchIS2hxy7NbUB2VADaCsnZghtiAgPWxwqvddYxR0
6JliOoqqymHuY/vnWRsf64LUMs31NyFpN448BU4FIS3A/2Hm0jUHL5VQkRfDeJOD
fKondOc/xhFx+BbKIrogtrbM32jcisqRi00VjZx5/J52d+rhtd8cse7q4YWimrPf
EbRnxf8uhYAmHG1ju33L6HfAon3nAGve8frknniCYM4KbW9o3okLZCYtJVlJZbCt
IKB/83GBpxtCGm6EoUMThKhEHDkHo1RiOmoR0+l2wbqaDEeGbBsf6fuwfiV7EE6e
2XLcuqv5g164DWdJclQlqty8kGazN5x9zKTbOQrw5pfbBhqlBN3YN3HYTVUhaUt7
rnfZGH+DZGvXlwP//Kv7DtzBgkZwPDQgxalZpJaO/brEPoHrYVU7u8Xs994MxSZV
180gTyJZ/oRU8qApj35YqbXoswximIL4fjmH+F1Brqj1W5Bs6O9gbyGZHJl+eHU5
6m9RGkvmZnb6vEcvQgDCM031qU36gZoRwdvbYDYVWhhEXdGmVqPQG7ocoiYhCJhL
y1nH+ZCmgBfA8VqOf8NS/sc1rEkHftYMmYGx/BiMP5f3h8jdeA4uGQFIAaysm2KA
6Xnf7NXjKe33gyrkxNl7px+VL4TyfuQqeaIBSzYb6YDY4lj1mtMV7dR2ofiDfSdr
bbS2zSytGrD3KhXU65jQET6SsVYs+hQjuWHeVgSa3me3dLVWishqbPR6k72qYWDz
ogEUpT+gFuCTehPEuMyLFJOIZBZ6lyNGwJ1h8a1LV4F7R40CJHHk+W6iuiyAmc46
HYbuJJTJjR/YcjGQmDdG+NItuC54DcYYpYg8A7r+UOOU4GrJEtdEb1iVSPOJug2r
JNac8poLWLFaxBQI32txqX2VHnz3PbFTpe27eKVMiE7Wd3U1HZi4wx+otC7RaV6Y
4N7jkQkK+rODuwjLeAPtI80OFcT5icsJ05JjjUsqSyHBHHKdojNqBV+YUbVqolMq
HxsRjfwYsGhzLicKWyxlsttlR4rw0AqSCYc5ZZn2K1HWiRB9WrsPSHS4yQkR17Sl
MOC/GRFmtKhVP/aHY3hlXki2+JrKy61QtFBw2SBSG2OZ8QZrzlEmIN3arcnu4U+U
NocQCWN6nOoAHecLJhOyQuv3wP1zF28555Qtm+yGy8qc++n9vNs0+5AANoiWKMAm
yAI89ry9NGJRZGConvqdCDD8KDDsQtgLnZ8nutTPEZMQFAOo8LTBYdCpr22O9rDs
Q3S95KtAJJIBewn/BEeI8zfwezE9C/3A3+2PEM1IyjdoVXJtlL8ymwPBk+NXnazX
c1RaKcaxJhR9KX5bm0i5w/RYtoVC4WJ4QjwkSPSvRP5xsIkMk5HLzf61wcTOnhSI
L37D9QOy9+Ve4sGpb3dsFZgchQkGvGw8LLJjkPuP6/OiGFPPP4tM3+LtStdLKx47
UEbZQBsSq7fI4KSA8ZLJVSKu6/Q8nco8L2ma10/lQOeleehZ73fN5alZzvJkbKZB
39EvOe7PnxhW0wOJ4pVR1WC/Qw9iu13Va951+hngCpNqNgaSV6N/kN2dGimmC1Hv
apGzuHp9noIoXZM/l2tuhpOurAMjIv3AlLIecSNNyagMf/fWD9xRh3YfWsEquqsV
NLUy6yU/EHNIcx5qMF6SgYDXzkKaT05kB1s0bYs3AmmshODwlak/i6InADjmdZ6R
WjOq+c5qx8sHlTK9dsLA0J86fkYhaDNiNm8OZKfs+QTFLwS+D0i3fS1Zmh5MZFsu
gq6GAeT569E3CW9aJV8WCLapuEl7XwoWLNp5xmJoKX9mUcPQ3Q69+AbdENvLRJMa
ap+mxFJ03gkNuRlVOOXUbZ38bh9OTQib/FUE6GBB3CcAl9GTwcBVJNOnjTg5SIFW
wbM1RqqlZHHL6OYa/C3KbaT0GUMcy4+P/j5Cr0rMVb+m/J9TkHD3AZKyviDsu/sL
PQsZ63vt43QglH5Ypo19d68ktwUK59VzNXkx/YdCUx0Zg6fJ3yjNIQKwjuQpy/6Y
162nuhexnJLEa5BoG+8UpbST+1NgAqwEo9Zh65uU4w2s+WuFnIGR7EIMoiUyPZ/U
40j0f2lXn++FnRaX0zb7TyoYWVTXuEGxIsLlq4xcKCDcFKzt2FQKE0J/CKzYA9G/
Tut8POASmAXy4dQuWr+RPAwP3+wvKqPPUU9JODfdguwo7/k+BhtDf0MgZOAQR8h/
Utk/NWGC3CW/MVGtSo5q3cniP1qms6ExNhJQZT6TRpHX/8bsK5DORlffF/Fpgv17
3Z0Rq7kleFTFlufxdagTyQEAICM2ImNQfNNxver0QKOqtJ80YF06OswM1FCYQ5FG
psWB+YUzkBnuhBjBlez0w9FZsk6A/hStfkPxnPmF1Kmcb93xqUIzVA1M7V+Lu2VA
0uzNKf36bdnAkq9Fhl7FSeb7VLWcyU6OEUD4z4kGGBd7OwRx7Tof86576e1xLuGw
g60ubfGGs9RwnBUBZc0px9idUWwjs4z1j7wTRv85NCisldOYUtD/oteUPOosfBTg
+z9rxDENFhJM9OXJ6a1OSN1zAD/xfS6eGjGywN7w/rI9B5CVSUQPIwQzG8xODF1R
iturQJbf8By7kCYDITTQA4yNzeKGsHjPJGGZayjg+O+o26Ez16UDGGa+YtUPAGVT
PulBpkHC+WFIUc6k1kgHLveCjCMwN0YzWUJSbOfIeepzq4B6W2py2LMbVzI+JXgz
QI+5PB2V1MXt9pmOrjTOBtaJ/T2olyYrL51xuXFHTg99PJaVztbe+w+56zzz5ddT
kNUFjKVU9m9KjVqKEzkTHQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bvyN09ph9OLb5W8jz2wSPP8AzfZERIsRjKP784d3mCHt407IIVibMY88Ea0HElLJ
FOOZK2I9EgI5l7ALMFYgatJQ71oBd+Fl7PlkQKQWVc96Pfp4FutAhEsujt2kQ8rZ
6CIgkXZKhIoy219rkLb6PtPOYykhuffE06f6C60xLLkoTOGtxdWpUs1R+ddnqUrm
kAwqp/3YgZcx1y3W/XuF8O+OGtRxMTKJJVDxSmHeaN9vKhcLwwLvn+ikTH2xzy6P
9vZuB+7LFCBuIw1dt7Cn6B3APmzVgfn8JEw9Lejo7YYzOIndcysOxyG6fQPL55pN
SWo1E8WB9CuiKQ7603VYqg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11840 )
`pragma protect data_block
ZQDI5KDwEWvzeVZbVja1/0Ot0WB0d+CK0l4AKHSmmS43BIbb9BxMfvO+KSn9jNQB
u9N2Uv+/JrRK93o4X61PTbSXLVC+8xa8e2fSXMsEDKYCUe52grU5zoY/T5+lAOfO
ftaQrci4iRR6qDDipZTkuN90lhAOPFgd/r0uBsI7w+35fdNO6EN+LaRcH59d85fK
GisYCjCQZifI78sHsWoNeRAt1ovFAUJtD+UqvnXHjKR6CMuRILV5FNrykxPRyQ3r
HUjkwArYPi3cLXdLDbwKbtKd8XHEsF2UAZvxs+jn7j06+PbRaictjTiw7ama/mrc
VvvxNoDA1Zeer6PLCLjY9e5efDkz2JBiBe0Uyv9nVnanvhx9Z4ZYg+wp+4tq/ZrK
YHKfEdUVoD5iGMBCviEBfizX/XVZek9+9Fe4W/RyEw6aNYwRACs12Yyt3IrACnar
6M0aRRupS1Sf0xyIcK2JPJJ+6tYWYMTlEC05zN/UP/LReShXneRg2xfNf1ofdlzr
n5bz74Os1VPRovewRUpFp6Jub960z1h16qyTdMOaNtAY4vReuVKIgSwaz0kAgUvX
2UU9Y/Uvsgo81VSabbNd/UKc/6iyNRBWOIskz/4LgUkTCtzuhwchbFUUnCn6KJoY
GMehRuqV4K5rI/uOrHJiHUq4iXMHjaJEYbJPfQde7JXpmECtkoaw+gnUb5vS88aI
iiMYNBC+7ZgZ7dP5SwUtTPj+U8bobv8Ne2WA4CNv2DOAD0cwRFXuxCfgrvthub70
sz7UVA9zx5M9rlOPCxKbcyZ4wxGP6U5qXNa+ldq6hEY+ysKjbfln1/yVHL5xkNwY
r6j/X34pzGJovAjGKjwevcTosUTufq7deWIPXjLXHoWNbeYuKAp/s45GPfsCx3ub
eWBxyER5BOZDiKyV9abN6F9QKtg1oeL2xWIx4h3B0UkQoj41xjLnjmILtE6y9mUp
D6A8/6s9LZ28tJ38tjz99KHiY3gJ1qwtZ5YY3Ilj86q6el24Unn/QM0WO9duJj6o
bW2AeBupNbubCPC3yf8bcx6qqW8OsB1lRRRryDG88XB2xUkfqRnR70RMd4kVshGG
xSBnIMC44hiILVxtII8K1dGmhASkj/TqhqPTdhWUr4lxyNO/4xSAANRL9i+xwR7v
CPrCb9RZq3QYGVBf5AcE4GNGL4y4xTbhznlINo63FlHGXl/c5Qgo1dnTPz8a3gcZ
Gro7Yw+9bvsMJrqOevMm/jjM9qpUukVb/fG8E48riPV1EEkcBnbcxjR5OxPWKpUo
fr+YkbPm1v65LMf9r4ZcZk5SIXS3rY7Foolr1gJ4Gc0/D0ZUnXejZBO5kl7T6+Fl
c2Vkn1Si9fug32y5I/NQAi7g1vwj+G9sfUoDupYOXSQCg3v2pyNMkrDZyYnc7ctL
lhyoHHS2A1iG6FD0VWSqFL18WrD3TC+Up7vzzKc6DKJnmDpxuQqhqH1uNkywMpdh
sxJ//HnCfhcMmHQKkUrrzFpmmFc0ih34ZSTZMfV1Xg+qMR1JcPvdHbQthE8I0Fl+
k+TrzRVpZBHM9CvWZrtTL/V1FfWIhbQmUoGiEzMZxlSDlXFepeeXtgaZeKJwQOXM
QyNLPALpNJGgoSXpxvHUaqHoB2u/U6lGhUNkZL2+zzrSPnwDMBtwarhbUZ87qV2u
Rgd8nL/aaHJC4KutyXtUCiLJ6tCUVi7igBZR17zaMJRu838a2NMG8RMm7pCEbLDe
UnewHet4KAaZv9Ao3SlM0Dw5m5+HTlY+SOFgWaNzNidT91mt04LlQ/tb5F2Zv40c
/i2glGwml4MFoiaGVrt/InHS6qlTKGdE4tu2LOrIBb0YImLAFxiuMysrZZbMfhBw
y5abdO9k+kB0I4LuXc8fcxZcqSP0MdejCeTo5E8rHpzwFWe/DouauHCiFfZYqmTj
mGw6xkoLRMq6D+pkToQuCjEQ9rQ/mibD/2/CVmaJXy3RRbz9BvmZbhx28O1hTy0A
ZYs9acmWyd6Fb9uIdOg0nASqtgRbiqQqZ1OmKkt6eyVvFMIbc2fRIrfTmXyqdug8
W5Ee78JqziF2mm/1r9vnnfo/y4s6bnrNlVyDI9Jz491NTmGvaDcgzy2AxqgkFJq0
48Sdk4q4Vj5CKkIUAV0ngSm1c7CDyprfEpJIe9R9fRyyWf5g6UFUtRosd4O9fLAy
pSy1OcWE7ic0GBvQjCoT9BQUIS8T/KkOu9iDkPu9Db+l2mDLFDRPBPwsrVKHlNHC
Jue+2eYQ9OC7jUbMcGZqZcBy/6ZeH3O7XsKkR0yNbSNfez6MkFp7j3TL7fJ6ffrx
4nxc8zYHPZg0kQj73UZQUtyWCFygisGb9ICTllosRx1EG/mG293h3UT5fCQOQb+Y
fWWEJBpaduyfjWSKjt/wgck2W71Ak80WlV8O0CFoclKjw1wW3YZI48atJ+4kWDdu
Go9HOLr+/2yvQuS5wZmhtbTI8CM2DdVbH5wEk+o1+H5CHT2Kixp+hlrN79jXYZTf
y2Ll4ezUsK2NLRTnzPRDqAPp6OdEB8a448j+w7D/5O8x9kfJzRPu/tLT9mqU/x8M
+86SIo8xQWF6IF+KWuWxrjAr9CFH95acFIki/iMCZfPGxIIP+i8oMbHF9NsXdH+5
DtF46ZIZ7WctjfFfkEiWSQgBr0dP+ORyWytQYV+TBUrzUlmB/QsmScOUpRoU7H35
4clqqNAaQwA1M/oWfJxH71pvIlDEAqIfZ19GDuQSv/9iHG4dInteJusFOejYZadu
e+/QWy0cf/q1L1o1ja3gli4FflJwWT/AgqhGC0IVxF9LSx7B9CWnBcj4GfIU+99X
expXDe2z5Zt/RYMwvy8xUKQYikUfIXhRoOgmbkCpEvDGA9UigAUc9AVRN9j8eMz8
i51n9aDLO0bCHxm9SqhrSuq5GrACIvhvZUk196IWgqXC9JekT87eWapFmaqiET7y
h68VTolYn41rnhcQGHDKE/T4I3X3tS5AblgJRl6139FxlYYcv5WS96hcuF9gbJYm
fdUq79XCoet3/0maKB8y5jMllfJaLX6v5iO3/YfOgG4X7aesdf9e7vq0mSYutdWY
32O5aVlMzPcYiVhkHitoZLdOHBInT9MQM7/F4WP7T3kWP+pk6C4p66j04+cIeYtm
pqz4tzBncnUsd1EvD5+q0BIiZg4F5HJ9ssoqV7Kyjd0JNprg9qkWiRDH638+s/Is
3ZT/Ogug5JOKpL2WRJ4PCw5NvLTJH3MUn4I9VtQqGPw0PRcKujUK3GM0MCFd/dMS
EQ7iaI1+lG+BfsEAMqXQegibnPEjusTp8Ul+J8wIU2vMmu55jl5EizPSB6hdD2vz
5ttWXGeush+5G7PQBHJ+baja3KmiQERnfClbj9bOy0cePBd8P5MXhFpJIO0DYEuM
sEkR0lWML+1oXIDCc11biN6WYw4rHLx6iQt68nbtI9ZNszNjk0CpyB/Y2NWhT2kZ
E6pkTNVmQjwFCd3Z4LTY/rTnfm0WCdFkcdPAitHQ+t+vFlp5RF8A4etxs6dDUl9e
2N0rtQlXKh0rvJ7ts+qUi5GxkWVsgvSZUsqtUMDZQL6+0qZA4FJC/rIC/YFVqH8Q
JVO2JnkFVCWyhheHD/ZLT1Qu5OrJh6kExt4T08A4BYSsSwSgmyfvVBBitmvC3aDU
yDWZ5SDs7kYSGpSxsnQDhdaQFS9ouPj3n1OA4jyVN09lRUHpnCHZK4We0QoG9UN5
cV70T56SPq+Q0ueAneEQj8wVaaOGZuv/1GyGWuXG9QL6NOP+MM+sykKgC/aXdHpQ
NaEg7Ki0SxDu7iMfVq7o4VJtraskEU9ECfJmLZXq4pZvbDI6kt81LlnkMGkPA/1B
ec8MGe3xTQeafJuPVoMgEsnmW9AqArbMTROp9zqJhKc5doBMxqiWtHm0V7gRvmXS
ZjU1ziL5MIjvvyC0mmVJDmmdVV1UJIIDmxAx2eU26oZyGRJ+xCwpQ1IINaAxpzpj
mbLOUTFAqnILO4054ykWiQFzAPKlumuN6NFRX01MSHgcFfcTkoQCuXjj67Hjgkrv
lt/YTJX1INQFoEt9+dhtv2zI4NtHKQVUf0J8UhVngiJ90oAguNP9HFRQ7t94zkDq
I1mVP9EibaibmB6adl78AiR8hOQmPWEltWm/e37mWAlT8u0w4M7sA2LqXZcPkUOX
f7c4USBuNxH/t+vthzQY6JL5Ik8WJMHdRHARprKpJCNGZq0ucn1RaH8ATctmXkPc
3NCgZvcSAmVYmAG2EwFq9o5j8cir9qIjh1+kzbUY928+U4nHeLULd5x0LWxUDr3W
9xr9XoKYZAG5UVmYVMld7uKR9jHu9lSr+TWYiLu4kabAT0Vaay0dGzg99Y9iQZiK
EmkaQNK8DGC75wME1wIhVCxPUayZZyFL6XKOgVuOnARTagu4Fhj4Gtz40/0qchXK
BoarCr18vEo/UDREP2tb5GC2mO/g4XAqt2Jj9BjyCBzvMIy0Nh4EXUS9N4xo0/iS
o3KnSEQS/ohqTcqB9+hBTSuAzJ95ubKdJojr++aE5K47TGW2BehIAMEOVOTANG8w
IeJ1U9lCWPtfiYKSDevM40qOEzFw01j1aRoeKLvnLW4YBEvX6awmEdmlOmzCgcxA
DOX+28dMK00O2satyR68XoAHuQxKtwrLx+DBzox4Yl2aafyB44sZKNh/7cKd2lNR
/hQdAnOY5gTcHCBaz+e8FwHo78+8USVhvPsUfwjba1rDqkSkJiLVPJNkMG2ZmnOk
8MnPUAbhn1gjgHTDd1O64BfMdIfkVqZ1aUTOzNF54jACL3dQN7I0DqGD9F9GJpWo
HOCZz2gDR2il6NG8d7vddvlkmDFSBRxLcL6M0Uz3QcfZfYeVIxWe91cHQU9lq4NY
7bWcDSKwaDx4pxLw4GE/paknEFrlqYQyXT1CZfoD92myjJIyWkfsMlfo9NmW6wsz
Extft+43WeFMI5Vl6WLYKi2QYT/4fD1WKX9QP2cERDDe38xNRddKr3IFcmU/Jw9V
LePgCpv5IBOCA96rt/89HP/0fN0JVOIe4CuC3kzy5HPuQwpvsuQPUtBtVLrrJ0pY
g/FBS7WACReUnI1tn3pT0PwbQYromikc07iXAcMUAc/W47bExTppBanlDQWjdOFb
TvvPyOMFYtMYPlHlbJ7nlv2oAX3is/G51XBGKlFHOIi4zjRmZYtFv8So35AB6TCC
Hi4QuFoHj6tpabl/77jEuE6tl1NnOyF2+3NsPHlJjWNk8Ef5SonrDziop2PkPBTd
J6YAA575htZLSdIHBrKU1oJvVvKlVzOVBlwVsulGecQQlB2p3Vj3mIXauKrE+euC
Cx9q/nqBvJZqiO6zksBeCmWW6Gyg1xIL5+TNyjiqef1Bs3LRF7nsxV8xY5Ng9MO+
k0/XQJvyUR05869FqI56b8oQbgVk/5oO3aUs2LY27Pw4PppahTJLn6dqWJF307C7
d0K9NX0EdInS2ueOG8ddTE+xMbmkIq+WaHp+b6YCe8mKwxBLXYs6mEphrbIKHFv5
f4z9m/AEaJO7sC2mbvIHfsZ6xBH048ry82d8e73TmfAz6Wb/9teSlFigyBucXvD7
xE2BqYpXT8AkC7au/sCHLAm51Yy/GV6Jen8MoRcjkWWhmC0cxFq2Q98V5Wvi6BuP
hgQ6l8vpqTkLq7tggVsE/okn4AwF2sYlLSVrhGBe/C2IMLngyBP/wiD6GbJ8pzSx
Tv3M7an9pBfGmB+9DD9+yO31x9YKaN5KsQ+xG83hpxBIHpGp4sAKD9u2xah+SwIS
6EvPQgt7tnnw9LVqxClJTdzQewfknA/wTn1MAf4UTC4nF+2jSIahZ7FVpg9+9IPs
gLPhEJYDxtThOdtrXdGysWuoYFn3rVP+AT0myJaIpKyDlfJBGFtZLHsBOx3+/FzT
G45IpeLLC82LbBv5EFYAlSHO2xKHd3QJ56GPlIy5NRzR+pWxMTnQ76rozwLR0x4f
Rwp7J8rw3fWd0sbYshnE7apMt+hQgbgduCBSJy3/g5/oqyA1ygWMaugUIXMIS3Y1
x7vmY+2a4OkxNn1g34WM8HZ0QQR6jkmOwOVQcEmXLufSTdznxP9i8IGiDVYy9eny
6oSDbFuVdM1P1414S7R4wl2UI7/9Ld/WnPM5qt5dO/UDrx8FhvdHT8YR1f8VnkUp
JlLpZaqqdq4HTV3WsXl/O6vR2DQ4TTAHew3FZS6mbNQHb3fJzOnpKbwW5ls5bzqx
WDUgVZITDLue+fgBCd7UxlzfyY3hMHSTXMqFM7EElYvdzTTDOLeVXop2mjd5OfoJ
LsubTx52DULVdaOrKfIePfDHypGTWEkt+15+SkYcrRZxku4OIwhXof/d384zauP/
a32RvIooJgzUcPJud1pFV4DPczs+QyCwQPlcqR5ofn1S0mt8rYkXWxzPG6so7Mdn
+J7aJFQoxLF/U2fTkDnO8O+EfpxoHb0dJqJ4pXwqlKTa70Cir8O/ypRxTodMzmJd
xtDOj1xAwtqd0buOmftdYVIsLGmjheGEA0xpYLhA//vwTnPewiBi/hAkHIh0VV0a
ijn3wh9EKZgRiC9Qtws5DYovxUVf+LxvArK5xpeDltd5KQhkSzyzIi6uqi4EDZeC
nQrmP5+Tc7yXIrg5edM4Uc35PnGD8Ztk7yYJe7Kg/a/PpPVCPXaY2eBDRGM6bQ7n
n2H2p9XV7ldEWj3B3dc2VNJ//+nkCUtOsB+niztCCZMOBhqcZDAJ/kXHwt5kMwnV
eSIBmvt0aDZMHcg4cwX5OBCumPQEKp5wnbOaRAVSLeejNKqN1YwyOQvpmzDIZ+BT
Denbtc7Fz+u1yiuhFG+IYDQrgvbtfnXwri/VF0do+pK3Rf2btSril+Y8QgSSD+AF
wCkwi4h7J5J0WfuGbXOYbIQRa963UNiO1c/uCXlHDfH7AstftGPOCDQVwSFlnSAf
CPHCEqJ22NbUo+MMgUoePaa9MLkUAnylbGF0rk5dfEIWEOBys0ol9V90s2GcUEui
S5odSRilgxNaJzve2Dbit9DBU8hlQm7fwG4zemloeDPFx+uTo8+KJUhFqfND9Pwo
BmqBLheZCfVHiI2Jy5t5SD14GODiW7w+D39U1u7LmlDJZhgLcReMsvOqdq5K7+Te
0rtQP8Ye10YYMjiqPViDMtdqkvWlcBupEMx5I0lj93wOxGFQKCePgDjELSyzXzbT
lnZZKd2PfMybeW0+7bbleAo9gic7O0TT6gK79HdSKYzZKyNy/vK79x2YebQ3yBFU
DxGTmFvVBEHzFvdH/AmtzxSOBcxvyM5EKfXuuzGczvV20OIcAL4rC4pCgEFBJqkS
+QhIy5CDIZgDDx5CZg8l2K4xqFcmJWh2ue1JEHmnUsx8USRa22sc1c7fHHYie3ZH
Tfneq87zJPyNrAqV3hsoNorHrUtrcHcuSzYIRYiN2SIHJtsrzh3z804SekUePsc5
Dy4BfzSHyVqsBSnZ3nK9f4QITqSfY/Uof3y+q11Pe+FrZEtVZHi7exXUL4mdf5SG
HzgYF/oE58mYPQDr2z/OW1rTaMofDFDkHAvAPNCpxViwJoontn4Jat467rhXeBkw
Pe/DzRPTFYkxwFgpvOBm7zbgawBIURgDuEqgxyv47MoNz6wScM9clXtTOLfMqKc9
DwNhs2+4xNZR6dhkrDBTEclITVU4CxkPFe3zowK5ircZ35OzeopZGOPMUCpNvyfu
AiTmucyBeS3LWrI8pttBGOk0G4w00i7uq4fkmnlDBpzG2cmN9i4udjc+To5MZUUG
vXiX9NUY5hvtc3zZ2DPqR4iFwdTYwDnM6rsPrpcZiy/+6f8OwqdkuSgJnocXx1O4
+cCQnpw2MGOMhk2eUfqMbwE9qb+TFw0QMRo6Whr0VkUeBIUhl1/CLbl6FszcdvNs
hZFAT4iTptOUZawywtjRkur9QDYbuWC2bKjyaE4cH9E6SSavX4l8WegbJQkd/3Xh
SJZRaR6c/a4C0ju5ISDmfQIo9H89Wgso9dt4DoUMIfhI4oUM9W/p4xxG02EOoA0w
G4pg2gkxr8ljNPdtMfl4TPSTYEPFbK108n9N9oFaKNXr/AsJ/kHOGD6ExT0tVVFC
qNPX2hXe1jmoz2zB7/gidArXOUT+fkwYuIRmn+cr4E9Ssdu79GLEoQvS7tnNI7ol
R9zgqMIDJBRQjrA8FS7o3txaDqUmvWt7ECxa0HPgs/exK6NeCDqGLVDqp3wV549A
Etm/siIpI5tZ4PmKkNfq01woQGADVT/6r8h7SuRAfchEVNNbyixArf2dprwLaXmU
zzSd4RbhD/FkQu9LpkB4IDRYv3H53l/Jq19KwtaPcvLDT+5r38G3ch6zTOTRSDxL
NgTzSUm74JdYGbZ2knnqpS9Q3oCOxIEMzS9P6UVjxTR0pgnQWvEe9KKPWNRONmT2
Q22LsPLIRgeE6wzv6Tcx+K6aB/PmSZRwIHbe4yhhl438CaFeMofkEJ6KemFp5aHD
t88x0zKW6vfdzfz94l+eZw3AFk0EUXvSuRgvgw5vhm+K3PQgzvRmsou7SCvx0e2D
U47KUTOLcKW5IdwovNJ/aalYyWni9vyRPECCRiKf7BnVqyFTt1L0ScdI0TSTXKfE
5CMNEBRBj5YVtKYK9jkh9crzrH786zO5Ane6xU1Awp9kT+Ir9D2zE30tgWn+8ezg
yrVeC8+aY1X4+PNnrSNkpF4MwK02TDpDZvuWYmb1zEAXIavReObWpxSMfTsHekFg
o+O/NgZAWUvg3J7i62fvhMTKuXzskSE6Eq7IJyNyUKSq+XA6SZT8gydNs6Q10FM0
KpdBWFc0HxKSk0WAwpD1m2R5uFU6phSFu66EG9KqwAzJSjI6ILxvJI9TBSwyN1R+
/BMHWCq5Y7UaaN1/QUsa8V2GnlJmI+jmQrGAc+nHQG6gQ6h89zTbBoEFEDo/nEBP
W1rC77QbZgC0EJ0rb2oh5DKK3WMpads9Mt62taPLt+T1Ffg3PYNRyRvJktzsUZlO
gP6L1y62jPs9y4n3OML2Axp8Q7JPMNC2VNCfscJ9JT/scJLUzCFFD6lcasFzxzCC
CkSjqokmJuhN5DtTFhjAUGe9Y92PvNvTSe+wQvtdFacKGqJIHv3htfnOqgcN9tAz
cnUVFPTq++K/xnPLdn6bv89XWuFvMIX3nC4Hud9V7qIx/WuDHlETOgzHk42om9WO
lVxRHs7MJoDv5Zj2mPWdtAtZLStIP90Np0lIwFJdPVPqwQXe5ptkGR45fFP2lED1
dP6tpbeeZzwbOTQMThKNz1GFrd0aoAs4o0BnA13Ac9nJdnN5SzM6F65acIuC2jM7
cFVE2xVjXBv4IpCAAPuhODjEuHj+7IaKax1h1n5g9kG+YCEfotU6p2Bd6L95QF9R
QXGAh1/hEpn5uuliP+oogiB32AH9WaZOtKGdLfZxG+AQQPvSJRNadnDCzKHdvHBb
7Vdi9aVGg+bqzf8BVeHLjd+SYlbNNsc+JYgb7csH+NsjalBuiJ+Fg03DM3ogoTkr
nd3Cl5nakcXz5YoNQFFN/7Ek15FN6IVlb4JGPG+wQMRJYJ1WQw7UrNYzgen5QczY
aur2AAzcUX/bt/zCfWr5jKL4aoxnNoG7TkfBJK8nbt++SM8zS+lMntvClQbWG6Ou
LGee0feYw4uQJRXBsiHH36MaFInlmRH8TrAfZy1eamC8sq/mWR8EaVNc75T4op5B
jHP3sOZ5nuujpRd7U68S+z6Juacx76yQvwmu2qT6Rwk7d0NJjR0OoHx1AVn0+iEm
77cnbnDN5+yVC+4qA0ebTRqNpBN5suGlmjKw8ITQ5NIa6Hbo4+Uy9/v2K4YGweAE
7HunjYFmCYVyGuaOfiYuCDxpBNjUu5ZnJpLu8fVEqXme1EJQPJgA2EuE6qwmfoYO
N+TUJvHVypR1ZwVblEVxlMVD7FEWwofOyd3OtuXWhZ7nxBXbYUU+AO9IAVjkItjn
85ui409/LvG9Qww/8i7Rijeuo+iA8RgdyTRXX4DVpgsNK0oka1rlnMMpRWvzhoqQ
u4lw/Y8gmnlb4Dtw4FpSz0ngxuc/mvea23xyQhOJLO+LLNILLXrpU7cQw8b2VgLo
lGqITun7+ZRnTvJyGwLXg9zq1Bj5OUGo6DP9YTWzLX7gPSvgS3SP+VgOk7UL0kC8
96hqHI7VfjaXxiKsWiVfmGN8YECpkgQ4cb9LWEXiw3K5b9YXMRk211VhlyfwmY0S
bMNKO/vuD43iJf6SmF2ZXBUCiNtxdWcyUC+836ynuRBE3SVTjCByJ/CS0d4jK1GQ
BG/xKnG2JV4/C/0A/Ah3d7IbRL7GvNttNb/MSJXpQjEbQAg8KVzwe10q14i/7Hvs
zhF0/wWEFokPoOnUa8A/nzaq4bfQR1gck1qyluSkrXntAWWgFtOu9zKPdHGdhmnE
e8bkovlChAqDNItsPa2h16awW3wewoDzZzCOhWZuHNKeSjyzXn2ri5Aq5XP6nhc3
0vgRZD1qkiwbfsNWt6XSc/GdtNstmty3yv6d4S6cGpTUHcVKSIb2nZjV9a2SWNij
AMgfj5fJ/ZCOLu/a0tQHvr476cKxD8kS7+1bU+2gb1Ai1NHNv2Ou+ZFhphJ66z5J
rv/9IGB4In6XoU5O9Nbmi+hTTV6hj8oq3RIR/oAnmHJgO/mo/+s91GSeIu7uHRGP
gEs6jd5PF/fwxPG5kDUogDvX/nqQj4B234lKNZ0svsVsKpp5phc944ExmuaHaMaY
qgy5zcqQDVqgAO23+SGGjI83IBTMoUgFgrU5SXTd4avjvLVU/HDo2HraszMq8M9e
czFrmdrw3rXq54GeETcJhYJFPN9rS1Z3+PRlx2CBZ1EmdTlEMthDT98AsYNwRUl1
tyX09OzlCLOGCqWuiVsjgymAobLSjIE5pe4jOF7k8IVzC2JPfHwsGExFCgKVIJWl
VsGXEV9HQ6yXh1W5ed1oVTdp0dXX8gQ21NtmHKMSEKAyZNNtrGoyVRSilA7w3fVg
KQESwFvEtnGrejkXqWpEA0zgnYaX61U+LanVPr5egU4se7Cmqia/NtrN8RNLJIdV
uOdDV2Yh2yVFZHwJb8PpKMbZT7d+u7DnGX40klL07XmVwj8vBo/aihemCQhFNM1U
9YZlkdfUiAuGjtvAvhPrZx0DDrHXKk3YD7J2uzCTm+rYSC6Ys+SsbeOep0OwXAWo
vTAXccijqKJoZXcLmFNlhyNbHV9RF4uhDPEkNaCdniOvvDd5XbiXa8pRbljgU8N0
RM8n8nrl5goV+fah/qf4hsFk6dFRDfO0kXdGNPuIdz/EUwFYeVFY4y/CZQiT9IyN
pFhdOUcoox2GxN3vDfhbGuO0ppTTkAdGgAOpDrac0R5g6Lug8QTi2aMSkAJcCFHY
F7GHvKNP6KsIA5AGQeIdFH0Qlr9v4xkjHRs3mH9JEzdP6cLC9DMozo3FfEht3BEI
6/tmlcKezn3Eos/xjFptlVBdUSBK/fTjEwJmIv3MX+k3Iqz9GM6u56WNFHbvOY65
gmXbv2/DHo+0WzF0fiomL7GfEX1ZXMUJT8ffXcYAxEI+8mAZeJKPNTkH/nrkppXD
vH80KaQvrqgsHtLQd/0VMpndN8IvKm3mzYQhC0QpEzbYnIqr6SZr6tWSDlyCGuAN
/YxmouHXA9LNq9nTFZHDJpNi9BtiTsD6hffnoi2HSo2szizju1BFDVPe/bFzpDkZ
UQyVNxwxtNHqU2UiovsFRYUccH52wWTxM7j0zSZevvHHvCUUEttW2l+YySIAB67h
NJPO4y+Chy2Swz5MnL0RGjILeTqjWBNmg6OLcHxlNH+4sPEUCuJvNi+EvSU/UeEP
D8qyGTLlMRXZRPSNxQs0wUWqjbd78hQdg1u6jy/V/PyXdfpxt3aTLXY/N96p68rU
RoAP6uAnUNVOPF+5G6B4OpZogHPvFEDAKROTKLXFbb43u3KE0lMwg4QueMyoLYLo
zmPCFvLFE5+oB6CUZv0seI5+1VbqC6ki879rjRelNEYvgWkonGTrmYjP1CeTuOv0
jYYDBL1C7CebIX91oSGFPqE91yTReEqUOR7qPmHCk1RBHIfc2AzBQRCI/6bmBQFZ
bz48SOtKKmb/+Qnt0mxzm7ABP4J3NmJk8khbIIvXcE8rhKeFYGMxZ10PpkRvXkTX
a3cwjISwdWJX0Q3huhxrMp1CH6NnsZCu7GVnTn1DIxe8dVC5Tvxss7etAsBnoJcu
Sg+7Y2Y8tP40vDu+DlaVsaI0Y4Oll7eME3tPMewiWV1VqQsQqzfYPEVmHEOnIb3X
cEYFeMGkzBI+Hss4acs4DLg4MAxFC80zZBAiOdCEePf37ALitazSxofaIf+0ABNe
ZZ/aVWIXp3ueQ1xfLwPvlwjnfs/oVIHTKRUfiS1f3p0l7aXK6l/jeKlwg9gH2oZU
uEEqmRy8NVbP0q8WDzl7kNdV+rls2KwBKLT47EI/1rstD8vDVUg+Osby/3XQ+gpk
khz55BVZU+boiu9o1nDgsrqisapRvV3NadxELvojIwMqUyxSCq22TPMB51RUl3f2
l1Tu1yltN/8mUkGBRHEgAj0Yn5sK4QPT913mMcOB5Z5EKzSiMrDi1UV0cNWr/njf
DU9mXnG51kjiVq7xelbM3HDYYNq6XEdl5TIuietGCvFIUANL9mV2xOW+H0IycPcg
4esAyNKCu1UzXSLZ1Jpb28ovYGcLqcsZR5DZuA34TYzzV4pJa8E+6vIBQZqWZR5B
9uUHEXIx5wV6dzGlEPuMPHM7znR8Ajx+yNtbzAHNlB+cIjUPHlVT1bz5N+vPmT4v
EWnVOY8irsjkOSjzTf+DhSza9tWVZ9E+CgW23Zxq2EBVJW+6obMjgfrFSteor822
xq1PhAQOGcXhrKk1WLcU7tNyPaj7Vbvie9pXYzycEn8ZLhFrpmw7Q1zBM5e6xPaE
OgxTNHQ5N2782Nc0CcmdWvRRSSB/2LaYiRR+uKPI61s1tlI7vQ4/Il7bAT+t0GN0
KcRtnwiL+pqFywie27a2I5yr1zFeVmUhybk1/dPcN2Yx9RYCtP5DVjbJh4IAtabc
+7le1XDxErss+Arw0ezDgNGDQZMkqE81aQU8ELBa1NWX5o2cJZ6EBr7ta6V0zO6R
pYWaoJyBk7fjD0qQus2n0P+iOs7a0lZ/IyxyKJ9EaXsp/BVbF2yGNIHaqS8lE9LQ
PP81Q0kmRgtCS8CxdMR7+ZUrx+4qxXQkHRE6U1ngYPeJf+3Dl73tFFJcME+vr5T5
gDmE8a4WnT68dYGeZti26Mn0k4RdGUTcjMF9b16PC6z4RDuR0IQDlDUGrWAg9jjg
lazzdq+pGrdXOKUhAnPY5UygVlnyOqOurRMhla4Zi8en2bG9pAsudABKxKovOW6q
jzzAv30nnTxDr8sqSQt9e+xg7R3r78p4/G3JBaUU8+ohDN1jQIRNNDFk4lyvG7Rp
SvOP9HYTQ54oyfQv9tHHFUTOT0ZHeNFE8qyCvYPg2Q7O+25kd2GVkMRCjgVOhjJW
s5H48VE0qP+1kv6iP42/bf7abZZOuG88AWLbjhF0QNqR+eK+nPasBwt908hjKpog
mMtdt1Kc8aH9H3/E1YjAZ0WneKy/fe1obso+mTANFayCGf9q54UJt34/9TGafpWy
qyg6EwhHGpKUXuT33w+aIwHZn0xjbJP0KUUyOtbd1CmbxvNbNW3bK51bUGbkPfVE
ia9sEEiIUvDbAq8vROi9bCbik5+gpCVp5BaFS2P6QBEWYTk+fsO9q3jLDKU3i4uW
7cbBEauQ/L39DX6MoZ5WfetbbARmL0Bd0gQANIF4UeSjWD2cHK5BvBUkjcqGeXRk
oI5GIwwM8rTNXZkVaxF/8f3QOuKdogyx0YKvnInWHkdhkxVo83W6i1V3aWioCfmC
2N3qK12sYyazlwb1R+dE7xlIjsGfGXanwEZ0FPxJYs/MPGcJaGu86pzen3Qz0hm8
fDVS8xJcCEu3bsfAhLp26OoCfqEpVe7pey7BTDG8i1dnCyQEc+VfVp8KaHLOaNoc
Mo4hFx+L4USD/J2PMNzRRZ4OoBbs97gV4u8jfrCY2C6PIQWQXYGQ6GlWNxTTnkcQ
tIVQ7V+zonq3dwk3oFea7BUMos2Zl8Z9B/Grkt/SP/Pxid95iTIaPw9L7FkUBb2B
t1Yan6JY2pz0XJA5kC9jiaAtREjx3UzeF41K1KvXJE+3/Sunmt5EX7T2WHaYTAQx
KiaDcoJCJxrFFYZEYSH1CPT5yVdBa8xp5CGYXB1ZRB595d9sVLA2H3Rk3gQOBQ74
FAfdAsSgV33DlvNv0F5TfnC08J/2PUpY13toLcZcEau7k/0NdmZ+3dtL9FFTaGqF
5Xg/TDyWc9JAXYpwIxWAjy602mdz/Y8tkXvtehV8m1CDkA9ddgENDXh46La6WEkM
2irmou/JKojHI+Ubs5Mqqv0ELaq89pKdp6zmXAZnGX6Qg4bHVGNRsmUAMjUJp1iB
DrWH+ETRP9rYs5aCbTeTezfKPDgD01YuiDSorpRHjBkhy+tPRxC4fRgmrbB/pfKO
aka8Hb2u3wnnmZuhJFcOv5OCCGi0Y/gcMcIgs+vmOl2Ca/CQToOTNGtfBJGgSj3K
DSFlGEIcsX104nJtzMbfh6LrVyB1gFEL8y3cZinThymKwPs9SQY49zhz5tbPNWzD
EtuO8emZ9is+NKCibp4hiLw/iBf9D7rF9zdMrTn2NuicLikmu7EXy9lYlqK9mDoV
PGFnmXEs+gM/AgnK3DCGhcbTxyMtA/d8y3MChWywjpNcJJMMLWHlSX9Cxv92473F
WSJcT2Aq8MSJdggNIPRl0ZGaQEtlkdTJCcrVzb1wA39ptrnw1i/7zqM5MocuXV9I
x8ZlF9GC49OYQsQaJtMn5RtLv9oacX6GJ5XFaaGiwHk/gs0ICEOmk9TN70saadwc
gx+fgVZGG9rOs7Ia1c8/V02CsApe0txbktbpFJxdMcFCCSGGdNPkw4lxooLTrIrB
peJkVGKV01I6CKQl/Qis1PTWwNvWL6nN2RfBQ+0taZ0S1jzwwrMlRMNEVG9X/gSF
YKBYjDiOYGEsfLWxhsjdYEZhINJU/hbVeJ0f5ZYEjD8CQi44ic97SXnUEebruwXM
wwP8usOdA+5eT/AA0dHMNs1IEEZcNXtRq49y5I7ma2ZUcu8YlYL3B1nY0TY7wb6M
hyRIwDcKUh/Ao5/lnNwp6MCb3J2MOy0on2PyD+/UoiRCIl/Cems0zN4gbFjOC3w6
wmgpn42G5rcn8uJUsRF2W6KvbYxuL0XZpnM/CAs358Jg+gfbP+Mr8Ycd9dFsw+gs
Wo8Fqo1FcjoDtCWE8OfchwHbo82p0kxkACbmBmAy1nwZXPwgsJNtkpdKYX8vwOuv
pn56ooIqOM+OpEBojBYWjop5faQ2JCIw4j2n1r0ol4VGV0l4sTyloD1yl/Ge1zVs
G7LJuHhK6ZqYUuKyTPLbcKOrHIJo5ypaqRQH4f9k7v8Ojw6DCC+uZUGiWg70dQ8R
HayOV2lWVXJ2lhBavDRwAP4EnyrGyxYw0JxbFoOyqJfeCOTOnER4PitpZ8fkSbTA
1valGqygy3G/DniY85KIiCUS69H/Qj/i2gOv5YvEJAiC9kKuhuhvIAqB2iQLbGpj
sHdSPaEQkSuNmqlO6yQwy5+BN+GVqsqsjvVgjSuX+5Yc96mOum2CCyr5F6nh1G+2
jkBFeV/kaCROq2H9OIbda9nrjF3qoooEAJuG3JiOgUYFPQvtJAH7z9nDxVXMlkVb
kGuzbDT2rw3rLA7bzmH3aXh1LXLD1AZDarhAknjHpFPlycUK6S4WSHnsxkXh5x8L
xjLinoLUMBxdseg1q00zTU/X9akCga8KGvyHoBn2d28=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
XoPyulJOiBt3oQrickzgLd8F5WVnOJENFVzis7rDgCs0Rp7xalXa90gG8ZCkSgVZ
aOp9pCtz2Ya5tFnQcfY4BptqmRJF8Cxdc2cz8XgFBPkWpVtxefZMQwZGuqGSUkoK
FESOEDsh5g0MPNTXehg92yoEDpfjUQDWKrlkYexXFaTzRlMscDomHo3R+EIkfbjN
lSG06jT9JPkQ5B5KOFDPBMUQQkJegOAuCF5t5+jl6MEgHJKdwx0cTtiO0S1rbSUw
usTkvssB0LtMQPphonHhyzPrHCvPeyQ0ay6o2DfLE2h9DXcYb0DqerM84hidfxrg
VIsixjZXGcRSnMcL2E/1IQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17376 )
`pragma protect data_block
yAitI6j2I3zEUYP076yCTGv1Orkwz9QmH3MTcjjKcQgZBCfD9lQW2sUR8HGDL27h
k9IoQLgOttqvkEnEaslPKPuSRK1oUHt+H0UVqykw5Spb/nkWVi8SUUMeWSH9rC4L
cVNt/B5w4RxfC5w6bEDWAQByMr/F55J0um5Nibv7ipaBPA4VK7xB4etE/NRL6Par
wQ0dgoQ2agujstsGcyM/GD8hkFdzBam32FoBstOOYwTS2+AK3tiiml5EefGoRfOm
Wl0mwXWMa8uuN4op9yfekNwgH8wRdz/CAm6EKCFeJ6bufa8vae9ZruJJS9NGYbEd
Zyg9HhPJlEEpXGt9TOfoQVAeNsX+DHx6m4lweJkcjj+aDNJMmK9ignxHEsRcsTDR
6oYSAHXKAXc0Wi7cgjjt+zln7MQkkUnoGFAbPLmLcV4JwMC/f46ruXYzWlUf1x1c
1sgDvE70OA/Y+zOjVa5M29S8wuz+OtpAGcERgMS1m1ZXf42/Mee0Z2o07E1ycT60
ms0EGz1LuQGLck0bzdNperAAoWfW0ErY5nDMI+uHtM8+ddY/OIyNeuC2Ax4tgJ/+
t9QXcN1Fk6pn78cCYbK414yqhrRqsScTfTumCt06ZE6JiuEGkKzrQ0I0WTHZmcJ5
eI0MHUcgvNaMXTTg7ikA6TACJBv370IeK5Ts6tYayzCZzr8xcM5JiakA/wb2eaFP
aih+bX0fsN4/JVCI9oz8g9+vCSbYJr8e4p3fbRAH/C0jaNhCIyjHnFTftJ9wECWX
lvXeGO5+SM4qzvO2dpVdjs2bIsMZ7whv4rDlOU3i9frDHKAqgQe5PLaDy/ftSe2u
HluZZLQRQTM6vcQ6T9YC+kae9GYAmGTGufh52/r09hjwPFYyH9zLypFBJwvR01ji
aHIZWRZD+5pwtuJLzZiHgOTkEqsR7WKucXGupZEcX6fKIJWC1FZJ7fv2yjFd9hpS
KssqurRCrT0UO8C/XTHW7fUYi31BOTTP1umJvHyTy0K2LEq7iZRQorhIhBBbZI3z
XRHg5MwsLyyzHF1A7g41h273hFANRuQ4ndXqBF3NyUgK7uEhX9QT1NmJPq7DTx3V
/Cs20ngWhpYZLketnuYj0lUkYozmc/Ea6DNqtn3guswWTGcVvsXCDBEJttoYw+qJ
DhDuGkOfMHqraqsA0Sp3PhKMJ+lG4OTWYZIFh+LvhWt0nyM5bLRV4D6XEFWmB4KM
FjnJB+yDgM+5RITz8oknYkpFHMYrk8KlarlnI2kvP36N20h0jYXyJvi5wG2Tr+wf
Qg3nFLJQB1uQf16YChxC0gdRZngZYRn0UPO/k3E1Q5aOm4pZHcKUGwowOL/1og0G
9puI7BCJy93KX2kEvsO3E/lEwLrS8ogDwPEfVTCvO2UI1Z0I79hbYz07wSpkDWLV
vbhzoR1wuJDgFMnJGMUMs8R1gO8iqFAi7folTC2QJobELVbkmK88op7b5MfKgDK7
tXFVO7YFkquEeoJ+mUS+av/1zash5GnwdoYKSXkbLN6rVoeOFQquBaVIMpThAlJD
pmJA6o3Bmbb5uVkXS/k/yIB1dAclDJs3moZaroGozw+u5ZovezlR3BoUe4L9jQP7
owIiJMO2qC1DbGwkwmR5R/NQ1/7B48IgwOkIxBJdPWC5q20VRgfCPIkoi31fu0l0
p3ubDWxuePKArxHOG2i259PlOmCGKwkKBhjr4KmD4Q8q/ccOFJXYUVyksM0a7oZP
mwUFAwCz7r/Xiw8WzWhhzdlWotlnx2fUXWVhiGJ7hnL8MZv24yxfxGJV8uiSpwrr
Z1ei698Ul6FWdsOoe2oFd7lFgOu7oVHplLLp1TlfjQlQKLXPU5pjV8MFVloCjUVy
dSrUEPaLmTDE6R/TL9n+uPuuT5ECBm70BVUtrttH467T3F/+dHhr2aUYqgQ9Nikk
uLAfK+3lRWmABQUbEGTEgzNAFg/A6JyWwZ6I+PBuKDlz7E3WnklSy7JED0CC1SQ4
k/6YU5kRIAomcR3ffsEOX128vBlMQvREJMT/ehCsmLlda8xLiqFXjZseRBNMnpeY
S9uZ1spD/gTUMIBLfSVVBkdgSbLkT7Vaf/unxgvMdNJJF4kZvsrTWsgoXjYySvsE
V9edD3+jIJYMCaJGVxOIGO9Gdwb8/BS5YraagzQNNcLg+Uzq3S3ixoRATmJGk4aZ
FN6MzIMhtwD0LLqu0m8Qk/B/GYcvTrw4uEpOhlXWfFFIN+V7OenFV+6uOFQO9Ias
6tneaMqegMT65769dU99Gc4Ekpumd+EYGILzhLZqhWSRsFp+kZBtXhyNsnsUXEce
T7GEAxeWUNyh4BEX3riAyjCweg2XufzKCuQweibp16z05Vpd+jpZg5Xmk0+Dzh58
EIpGQNGzDOTpjrgo1di2Yfx7Zkg7pHtgyWRXEMtIvKX40mcUzPx6myaCUofbkkxQ
uq2AHsEWGyeyJqTpURR4xOP7MinpN6nkrHGDZeGvZqfiMRRWIb9g7goR9evYoeYy
8WfyuSuMPWbDMJAos96bMU8Otw3Nm1Ytvssg1HoUOjTFF4E2Vtm7ft+XrnyM1n7q
Sq9RnKuLJ/c8LZ3B2YTU3E+Xfz59rg9Dhf+rc/7Wlg3uTsvKWVEPaPCuQwPqNf/f
5dnNsW92HU+3nwnxNlagAExXgYJPdSQ/mbwJrH8WtlluA7H/jzcgJyOnE8PZPcVS
j/wnEJMCoztAl/+O4fGnVOJ5muPjSwElfBYj6g0qKsiPBXEQJUtVStJez6rOsy5o
ZoMEmIKGCyhINnz35dUBt77H5FBGuHQO+LsiEORhokgid6ZszZGHx9hFRYxQFOIU
kbO5bNkeg62GWi5SutF4KYFnkeQhSnHCxYslPmQoBKsngQNqUl1vgD0bKFQ2YGzw
/8rxeUUj/kCjKkDAeB7OCdI6flcNbU+wn/coMtWOsuA7fN6SKDCBLQpzt+zJTpj0
09F8XYMkwOqZrAXTVapyqDKnSR88d1Y8gVR9SE9mRX9qoVr3ohdS4tLdXIWfYhIp
07FDlqC84vwoz8nwuApsfY2RCdr1JnVmF0FJX8gfScGM8IDL4aP4VyyYRFA7Vjl7
+jFA35YMs973qSUXmwekWpmtqlI4LwJ+PNbyq2g80Si/gUv0/21vG10tdVJl691g
d89e6Kexg2lyx8prhLbSS+1Wffo5iA8ieGueprrUD0U532V0T8ZCh8aFU5P8bu6Y
Qoech16yM4A6fRST8uf/3ZqavhsD0beEUK0VlByXja04K7z1GzAVQG87kYyYvFeD
vLAb6zHj9LdZfoToegowTAyICniqe8DHvmpx0LGNOUuotiInZVItx/+SteshZI0h
+HHaLmGV2Un/iWkL38jEV4jqCiZHPcSjSDYD6IWZdPK0LKqyVmt9d4hVOmoTNSIt
zgovw9n0lCTTYp2Bu7Nj/UBVxQgLmGck+TM85QN5h/jSqLrDF6Px7TWrlwxDC7f1
cjtLxnBSL1j1mNXIODk+m5JPsVHIzgkhhQf6fT2aeem13oz22Kej2Baw/iaFC39z
OfzJF69LxSMsQNILx4bYM7OZ9PkI6x/soqCXqYtPHE9fciQyp7+nuyXvn7LyemJJ
IQO63JtXPHe8mxZFl630Yf/zs/bX1Yy2TIga/murL8JWmUp2GBjzLe6Fayyl3n4d
6C9x13RljlZYZg0sZ+WMe9ejyO02BHV80pM+lONXSR3FvEG2gyShzJ20IGqxp/as
4efWl1e4uc2OYmfyqXSmPEsJt1JVWxpuUSX/eWbcTj/V06lMIjx+zs+dbxiA1ZlB
87Ah/KBdFeQoni8cAmzdSjOa9D7x4f3ihlWMmkqxYtvMOvbUIpR44LN6OZQV12+W
g4JFelFD+5ZfT+lUGp+o6tZROlDI/S68ibE2jSR7ESaj6uMASrvMpPsMr3srY2AY
GsQFHcO8+9SHoMt9JqHQst8ehG70MCsDSuaPWecHGNUP+Rf1VsD0iOBm0bMHI8bO
jyIP1jnAKBWHOT9Zn+N7e6ZxNFl13XGzx3GYRqJhUxIT7n08+KNHLUL4PqqhY04M
NlTSjjFl+SymfLalGyfGsAMkqSkL4n1gB3/RSu3oonOa1DtjUDy1dAZH9DHKH9bG
9wzztmqNYiSPAcJ+yqbq0k2NEEGwSf2McmvB/0JuorNkJIeYKcIXFlNZ/JsMOm1F
Kf0Kc6K5r4n6MNGdHDLzCXrysuDcaSw7lU2YqQF2kPokr3E6eCHE5qFmRDVGhBEf
ittFMixia7KvXmXwlHuqbU/4bxZBtOqgkb00lDBWtZlFPac4RTffB4NGO+3Z1fxX
CoRNIZKlrK3EUMy2DvAjIZW/Nzze2TMxU9Y5LXY1o9GUIEmok4WTrowJh5yYc+AT
whrnQfoh3REvdiA5K1aQcM66gQbgKGQjVOfd9KAiF5Tl1H0leBjuFdqIS9g7onuj
TjicTiMUI5wrRTm4iS2DEF7xaxtYTCQ2OziQMG7IB3C5goLE6I4X4cCwERnpGxJ2
mptkNDCL3udFzKIK/LcApZUjYYZN5p44RhzSpAP97SF1yldgyeXgqZxme6vkkgfA
vVD19+Fb7m009RHW5mSZCSuFpPKLmG8lUzP8ZfsPAZmULm8tTTkKSZozE30uiHgo
h2rs5/y80PyzPFF7dKTRv8BwBNHf2Ci6FwmdR5+yzVhzpad96fw786oRe/o2Z7jJ
uVn1xGQWL4YiKTZZaZz2+T7sem+67+XCyNQfBXv8h1TyT+Mmb3nSeOMp5CwCjCGu
EXJPM9TgbIaD+uhnaZcyieGDRh9SOkkJqED/7yb+H9J+TfgeigsGFDucyJcBzMMu
mz/GQBY05BWaOvP+8OEXLiXTA93nMiKjSGmP1S01C8x8DBTOyUAuSMJdmR1HSEIt
tB4pV8fJnjiyiuhi4l1DhCgrk0k8T+jWS6Gx8Bz495+eaJvPClce/BbfV/KYTKlR
S0/oDamYs49qoS2dg/v7uimw8L+0GVGEOHLUIDDXk51AfJdgqq0J80j7WT3oqYRk
t8I2mV/etldvWlOhhyc5ERWIXRa6zB//Q2HuJicnlGn8Pubf2eoUqVBwPF6wKgI3
OX4RSBvSdUXCUNWr+ZLKeTYA6i6t7aZpcUzaPs9xPAbSpShnL34klN9cKy5p+xxp
57SPgns0xJECbJlNyaWbHCZe9NvPsfRYBYKHLxwxAPB13eimhslWnQVjCuZcM62N
XSTO5WVULyuVPYlhUSnuPmaKSzRduf6MYJ7r8tUe+VGG3LAfJecYPxrKz2Oqr2vh
vZpyjeJObHAaJscUeDjMeSPkEvcz5KBlBNmB46ZxeahAi8ECY7waDr+ogeR1nyE9
ycChtEQ8/38VjTMz8kp8ZILLKgU6uyfuLuRitESYjnV+FqkCYQPES68yxgPvMa+U
uckpRvSh4jDA+9Y59wZ6K4cRqEQQrfXQoMxAOjFmMEJvdubKUz/ewPnDP56jcSOv
7hp5MhdK5C23ruIaIlaHxS/E/5d61Bpz5ghGkKyyDKnkyltRn3LG0V3q6b877WBj
vSjnmbTup8bcjTdCXmV3fSWgB6Lrqz9E/3tjPWZCGjgCJIziVTeBexYdXLyPQX/y
vl6E9XP7Fz8iWaF4amz4UW7Qd4OcI9C0Rxnbv5ezGq3JlJQCmPLcoOL42hIMxWFj
Gz5heq586fNdOmkUEOuPRQjWgI9TeOoehubM5b+d2DJ+NlNBVVkx1LG4CL99RiFL
G2eGmerzJz1Yg+F9n7KyRctPWsd2x5e6/Uli/h5anv3HFx1W7n6Q2ALv/QnY7azV
+WXqsiiBiJEC6gREYpQ0S+kPAUTkFVZwXR76/6nfOdYVmPXBwGZMf0ynq2fYeyDB
LtYTp5eb9dWOJwZJ7m8NFwInXmJb+lqGTpxyQ0ECzICjN9UKVHY60KirJ2w3sXkJ
TAPn6eSxswQkTpqKSNdbw+YIYZmYGwWmi9GX84X8mB5W1KqI2UXUTAKmJ6dzb/wE
Xq4/Is2x2/+JiO7i/14wCE9Yui1KgtDdy24c8NxjS2izte8W1qO2zDRtkDWR1bCo
/Hx88Gbn6UFn3p9w2SA1QrSHJN+t93ll3FbvrT+I8/wS4CgWaWlWhi3UmTqh8J/F
+XjpfYoUOOIBHP7l/3zntEP0dxqeCDL4XDLqESPX4U+8u18bM5jTuF/8wfeqZoQf
BRJS8f0aLN1GTi71Yjjdhok8523GCX55eYKNEkIRir/sg4Trg3j7MXTBCnwQcirf
soXjPm0STmsSp7tzGARKBuBxGyeH814UKlkLjPqZKHZxsN14ydIhjnBfS+55Ddt1
DS7bgps0dt1CmmWWkv582Y4v7wE17+NouzoppUF6Exleu9X+ZLNXeluWMUeOxPuW
GAF3FAMBDckAJP6kt+GxB1zZUUoit4F7LN2QLq58QTB7cV2F9KWYWSTL78GalpiT
7BFcXHTYAjxqK0rMSOR8SRNeKwFs5Ofac4nD5jV9tgDM4i1Uh54M/uU0losIqmIz
p7EsJoQbTsNul5pRQrgyyabRbNIWtRyj5eQQOlOsVcsPg+bThpce5XjbA0kBXAwD
FeUpy/h9IjoOdf82QmTcjVmdWSgjYrDE8b8s/RG6WJ98XK6ueK/WQrpbAO6lApow
TVojW0T7nLMLHSv5m23rfu7JHIJKHszuucYTVff8XEzfmtKjp8WWMZvqWyQhTNdo
/3YlCRnQEd783g0/HzdOHZsUy8S3IfFC4c1RUuwjEfHsER4wmVVpeOzeOeN4DsZA
BSV/zCnzW72I22opp/i4NbXQ9uzkE2odPiXtwPthYa7ShwnedvgRpC9qf8t9+caC
Z9pmKxRUhaXwYmk3WdqUh3cSvPDmeGGzf5eTUEv0dMnHIX3U01Nq2hp8U5uH/FWz
7JCo0gsKYklHbhEC7geWpasfUjV//YUjd0GRIGS5J/8dtn6bwbZ+YIi0l3W9SOJH
xzXTJQBRgtYfHaNhKdJvnjZ5HTfUClo1QTnqK7fc9j8QC2kMDuxlTYFtYipQOGtB
7DURj6k4slK9IOadJwcBfj3EM/akhO0qtuJhAIHnpdtxky4mpdtvrZ60urQM382K
OipihrK3SB2T84ns7kCspTEq9GEiNtW6BF4F76l7IrwGBasBzoLQAS6RW5RY9AAl
KTyWCNk8c9NsVG0DnklWcm8XiQhX5T3lPZut6X6FGxGJxXVT+/rG1cX6q0EC1t81
vfuMfKKF1VReAR3iHSuga9/5gNjb6+BDQD1hXgazTSPq/GTqDg10bVLF4uzRjIxL
ygZEJG3IXu6qACV0eWmk3FUktjCgiW6D9E1V3Dmtu+aYobEHc0Fw6wyT9KW5Z4zS
Gqr5BtV9KQ9SrJrttSylPB1iVcANdkvrpp7RoocdiUnJUPDsKbRTitFDIYmZtP3u
yVhpGJm0FJ7jUIPv0cT/74xEAJN6rkytXUH1UMx0S7AWQWUPiJB9sAkf8knRtVkW
6vomM7Cs8hFglS6s/9dAnKsE20PBDuJb4ykcilvB0LVryO7Wu3bucsvAnBuKjnMi
BUOXaSpyjBN+m66tMLscocNUqXRkyS0m6uzuTK8f51OCxR5VfYPwTZexmHRzbyzV
T6FTSdNEALpkUq/mL0/ArdK0CRTpqnbuuFX7+d2ys0xYYwGKrihDYwNjQOKzU2ez
L50eJ1xlx7rd7c3KpZDAbIk0Ne1ntjZB+MCUtqqcXM5koT9fst8G4YWB7YqWlPw0
OgeIFU3xw/2AA2hdRHtZ0hN8r2JW1x3shLGzb9jLZVdAWOe9apcC6pk7CEvxh+4j
vejd3R1gTkjQsVN7c0rAf6FKw8gu9nOqy2Pb4+58cDLzoy2qTjmd7Dl9P94NxQ3W
6cy7O0a+niDbWBayUxFhNtBUVarMNFgR3JtFO1lzOd7UYVp1oHQJICmkVNrQysNl
60bu11SSn9KEHhjYM8NiDsriGyZ3s16UmVnuCZdj3K6tdNIG25oKmF/1Eq4J8TuG
cEz3SwRkd7Ec0e/ZB8EoFqEc0wSAqrCsVe3CR0WB2uYaTCBNR/ygYxtFD6tR2D9/
MCNUmuZ4ZCUzO0JzcYMukPYygXkbVQd7SYe5KYlw0gLJ25UyTO+VEgIVtLHBEawK
GJz6eoew0ESfMpCGpbnz/o6daeQGmSOZFIStsFslpGdoPYa5aCwzp0P+PjqdrI8d
x8ObdDaGSKNLUm0BsTDKhvAWzskDSNd8Aeew5svt9zgJv6Z6B04uvLO0S9UxE9Os
V+AW2M+vpY1SdgDVE9vjqUBzfpOKokImPcAjY4ERXrnEgDpyjgGgFRJiXdNX1uQ/
PVBvRErYn2bcaLdpmjdVuaJLdRSaI/qgm0HDTMuYFCclsQrpBaMbiVPg8/LH4Fde
bi2EU0AHRPD/rlOJZnyrmXg+9j0TKXgtRDdRd0Wc2Is/MLfhi3AZ9jCoZ7xqkriC
dZuVkoBKvtCTvV52diMQTFqM61scwCV5ntIl+WZsZRO2XdXjRJgJLyFagfWnZqMY
tEKiTYXPSM/KG/FwFqjWM2glCTkJRVjfAN3UYK3TCzzRFWlbVQrz3w2sa8LZw7DI
InsXYLZdbsW4s5lzLFnMpXZwu9hnPy19WV1zJrD4/gpPmNWI3jV3HPBjL9I9/3PM
28JGCJvkcf8F2axLEjKVoHbsmuwT9h2gO7POlcobI58WvDCfjL2NK6cuOT4RyCk5
JyjZ70iiFT693m3tr/T2kiE1JPHkdkl5JQ2dMHWJ6up3rZ7eE15TxcAsdxpc/07U
mSnqCUIPuo3vRQ1WTpUhRV6LcG1moMAajS+Q8hWknpD77L6ijfFizlYfyamJkMW4
0DimQZD9QTd0enJaINVbhN5tKfgmTpwTzSjDnI84T+nN34abzvzW7H/F320+X8ju
auN86w+W93xCHfGEetvqHzR4fRajrrM6VejNcMIRoGX0uMw+wZWceG7jL7hp6Ucu
RBotzSoWZtHVcA2p5k2l3KFxGnswGjwMUpr1NnjnkdfpyEYH3ilwD6uNPzpWGANx
FSvZc11vpI+U5MDN/TnnjxQloOqmukXidGS8kh+8IOruGFy9/qvCmqIvi/tNEEJ4
o0Zkwg962XcZNNSGygP6Ei4sDPH7+2FZaHcsqJ0oiz4WQePGNdUyxz6GW8n+ugwW
nWQe6yYMvGyVVcqdioD7yazMS+NYLm4n9mVYrqVuxZU/LqQNQd5q8Ym8bFKsEXeE
DKoC1mSxV6nnzzL8OQOM9YwFyxv4j9uizXvIYD/JBkjysLzpDBG48bWxe+M9i3x6
8UTyks7Lojn7VjqPFYahldK4tgoj59arzV9aWNPWAyIfUPDl3YcEQEi3dc115DC/
VXuGeqDwfFCVWwg1bkOeDrKaUrnyb0sNVdOy6geFklWyZq9vORsYwWQFGHkbPd6m
YIMek9YeQMuWWYGNy/iFHBCgMXfXr95dQiWUnH0QZ/s9KQlRD+hEXrFFhiCZb8h+
G+Dj8F+pwMh8PJa6H4wabMT4jgxzaZtSq1ND/+SF40luJHs2VYqSXXYjHsR9rnjb
fomk/XkAVqhGMTfFDepL10Z8L4YgkSUMJPWbDKMRxDKqxbM5E4/X7mbJbW2Kk8in
lPOiejMNL+oC8DkdFSnSM5pFsxrGfJRybWBoM+F/duoQkucnxXGhr8+4hScK0gWw
aTxj0p2DeIp1Uk8k1lX6buBN7YfNWyFtQNweqHtFbF+61pVG93A9IYRfURQVFlWE
ADfmPjd0ZIuMtkeFXv6qnCdei8PyXnf1YQF3CX8Nja2nlmXTUf2mnoLxAZLVVpV5
V75N6efdVxGDgsmC+q+ndaiI6dNOaISlTuov2THRHpGiSMGsh5+digOqt3Rkh1Pi
eub3sxmA4eTKDL8ZsmHIjbdEPT0Iu0o6BKQJrbpHeB67Of70VlVdp0/2CnqIgoWe
3HhVbjaSoqmHVaVhX9aTTAR5oH1cOiopRE5tTGSB6idQLkXHZvtHrBBC1yAvfMWg
d1PrykJOc6leARsUminfbCaCwE7elTpA0oPb6tSqiB4ivXWTx3o+eH/VGielh4Wo
c0Ii2URmb5kAftXxqLoKkj7HcG5E3iYMJN5e1eUmhhoQBYNv359BZ9X8hQC7ESpf
gQTxmLBrTB/JjpRXh4StUIcWNrPi+bgMxGcpgtd17ET12pHs6ZRo1UogHTSXfY8V
RAfCfEJCgoepU6DVOIIYvSIQSUBSJRZbUtiGeHC+aqYK/1o/ujdpMSoCjdud/Y0H
uA3F8uF+9S2/FLOu9xXaBmuO0vqDDATmDBKgEoOfmoPozZfVu0KdVJnkxVss39G2
9F1M8MGmBLS5rDVADXsf+Ip1rL+rf35Z585lUoAolm9ZKikBDWoC1im+9gCH/1rD
DG6tWPVWPWfyh32ZfnPH7IL4I8DZWZ4M1N34Ijj6skmOrKpxppeBRDvzGx21VZzf
d0iT+bZloY+HE/cKbyjulf9hKDsb57+Pjptw0bDPDfNK4snO46rKTmqI2o1YuqXE
6fa4Y70pDfG7x3oxsYbkLlHeqiNAPqGIkW//dypmjydiyC2ngyhgRYdVjYZbzmvp
Sqq37gm9mzQ8uLDPGOZT1DWgZxa/90ype6VQl2A5EuhkJdHj/fe6VF8/8LMi15Wr
lsW9QWTYbRzbbyAwe6BgJZmwFsQuGE1BIawhWSS9rMUoyU7og8dHcMPI2UaZLs/B
LH7akkmkAPnVZvpCisLuW/rHEBzVWLMdoiFfheWfjXc3meMCGoK8eNgRp3OlhCdy
Td6b7JowmYprSWooko64q9NlwlGQmiz+vtZHjc6Qi583Fz56OUuUg5jaNS6/ggrL
wV5omFqzdrIqXT/UVoRcXEruyQJqJrPWopBN/myMBOZ0f9FIa24hrciHXB95LWnU
gU5oJn1MrTpkD9laGEW3A7QIq4OX+bJh6GK8ncwiLXkmA2U0D7N7RG9DeudzuSsO
FVskEDRuRW6ROklFoE44ObC4dCN/VDI+t8g3QL+etAqMDRgPOhtewnOV8nU8eKrA
EP56nqjgz19hTGH/X6zbQ4ObLAURZiTu4oeWJYPir5tsRDwxaHBevMvGU/yHVMTZ
yLuasBir7IQKbkL3cauBxED4mhj7nY43LH364/XB/GQiOba5IW+HahDv2sV+7Abb
nM5SSazdNI2pD61i2LHTZAvqofOCOh8jkbSLA1UZZng3sP8yY0QQwAe23vukth1c
BL8ENl2uohQ4g7Vluz3mwW1uF0tIOePZ5MDGfwD0FgNRoWwvloQIAsAUhbNlUb7y
H9xa5OWKkYNjgzVmUtRWB/kxS35j6/Ww3K+My4CKDAOyT9Iw/usWa1W3uGXTnCw0
vH7PyphWj7PV6iKxSQLppRNxqg1uKvbfUO4wyt5dNpoS1MZeKjURjRwpgOZCtRl8
0wgu4KEBJGcmThUCznCD3gT336GxDI10kvcsRsgxzDWU7hb5Kr7WGhUEqXOTtA31
HI/eKXqEJ+uRBkRhvvjmYqNbkfgiGE+dlU3qXFDlWI21zq3xUB0gl6JstGoI3ZF7
4Z9miqw7Tl+Xbu/ieooKefSGUSK2aXqyuvZ69U8R7tlB3bnFcCpKUQPs1jTNOHp3
lo3Dz7tYIL4KsLcx4c3xVdUl5Lf2kemX3sFw7bucHwKxIZJk0jpFn4RGavn+2cwh
cqYmk6o4Hb6dLhnZSqbQdrhHcasVUrAjrx/5zs6R0ty6+GJXTYnRPSWofUwvS4UE
uXqW6vPD+Lnsrqukz+WJVSBt11zEnJAmYqKOtfVg9WBJIdLmPyBmY3N/X//wlavu
/f81G5mxvl6qPkHe2t44T1U1qvKqI75RlkY/WjLse6emBEdErCUEx/03fDmK4VA2
n7K4jGtDD+zwVok6AQmF7CzcYAKfpeMpvJKq/hC554ANu5Y5w4DHje/LrtTp1v3J
rqqHIi6z19vyt/NXXjcFMEpoEhgng3Isy5RA7A7s2JpkB9vgLEH04vKbCFHMyqvO
/JXEIBrNiAaHxrztIBqGHYJQnPYy7bV5HWS/i1SmSf/NUaLwIUvHrL6PF3QszpVs
FOIiYD9RGLP3Kv00ysq/zAMzcel+Fg0Qur0t1/NBUNCCAG3w1cW6SCnyBnrllF4J
sVVZlg/rnIq/mYsFqVW15x2VzizhZFZnSzt4m3irdNK3B5qN2vA85e8hWSw9gHKy
oEriyavYOwwGxe+8TVJiwK4nj5GbY0Qnr2yq8C/OzUGpmLv01DvRh58niUNg9rIY
Hx/xSNs8aPdAU/XZrNZqjHXmtpj96f6jBR7Fzxuk2Y6+hX/NcjgKbYZnfDG3lfpz
1F02wOw4gkNEgofJqSyvSwp1waYnrXgUADbof55LKfauEzoVg/oI/4OzoAqJuFYb
MNcKTX9EZUb5lwRNMtF10XgKlCrThuGKS8EC4kNHicmV4TsQgd3e8ZKpF8ga6IcU
f04EETKz8uRy3eEvZwpMCb7dvZ/gD22iDEwMkKmWRxXYRGrhyrOyfhY4oUMpDIIT
ddCxG//8/wr7w578hNwivwDVJllockbpE9x25csZmXJX32YXhQ+brGH1G38S8mx4
XTVwoL0SymXZ0LEIErvLkdbTznRSoPPNcvJRUCZ5ETMJMnapANhS4IlOUO1+mUX4
EblDRRxIJgScNcuy6ikMr5B9PrA3ptONISBWzlvEYBKOM1fsbbAdHEVgKIerediR
gRGl1plT5wodh4kai09XPkitJCq5naTh3TvOKLuWehX6rjItOIdSb74YttmeecfI
wGgnR5eCVIKmfilvM/n3hJFJfUJ1ZAh/0xuJrhArLlmXpOj9xOMpgTvgn7uGNSY2
qwSfyMg52AbNjXzTHVnTAyDqoa4jBgWtHaumpNiKMrQFzS+IyYMkDYckXtkI+N1j
N/Ff5Ill8SpRhruNzv+RiCqFrAnl8PYT9wR9NwLHy59A8cImGwq0szu5vgkvOsC/
TbYQ5YtD1GPrnMbKwqx38tZ+xdEcA/7HwbEZx59E6pBOADYtFWyiC19bJpm+2bp1
FspNvgpa75tHBhEVz5zqNoEo/uwsQnGwEB+wMH9iXZPVqfuDBNCHPY2QBoY8TVVi
/7g2sYb+EjUD6Pf7QitR5RCbXY5LCqbkXEK8zBy9PS6j/HC/y36Dfi/ij3Fey5C7
AQHTMC2bW5q/aDPvaKLzAb5oKUQN7hajif05QogdGU0dS2Rrla6kY+dPgO0EdBC0
5vAymc4HTEMf4g+v4OnOT7BWAaP0HtO7xGZESUphS1Bj69umerSE7Z2p2PxUtWsU
DBeWj/mmQdk2x7yarGIkKgYgcdXZL4ElMEXO1Ba+4FdamQAD6L13D2T0Uagxpr1e
GTzCTflnzOD434lHIJ2FCuPMvUmRu+zlA/Bfidi0Q+JRj+AYyQ+TRcl3EuhbcIAg
ZIhN09Dkg0dyZnvFADvtxGmLZN5oZrokj1OMiK8xEAqF1/EqQr3J9TI9dgiS4kxW
3NeOPl7sBfTbrxzScUaWPJrH4B1o7UeEKPncRFeepjEbhn7DJxIATt2oiuhcmoHW
vkXnMK7BLwOyvBnr3oCHM7dWJGEzrMmOmgzZKSkWSfp4Phml7pMgbJj4qGjPhOUq
aITfunMaGl+u5m/+N+9GaS/dfR81HBiS11L8U3LXNYVh2MbRNnxUFyT249N00gMc
3FvxYJvoFTNamWH+ukgyJJSv34M/wGiIoYSkHVHF1N/xTloXL81KL3ejiIGsHn3k
DUdNmTgSGvlJxpMdLw12yORthdDUou7wWyCezIo1c6ft1bBkMWZgYwNM/v2eQoCe
n7TPCtSm9tKNWQejvT/l6p/oVDNzdJ/fLnSgzXgGuYZlgXy4QZ9w4ZMuDfQpnJkZ
jEL9KS24UmkQVgdcARMFGLZRWpX0/EQmiydropxAIi47qSW6uziswK8EEodwbgGS
0OCggPmPuyDqXEeaRQ0MdQ0JpyrsZggylu9ew3eq1qZXRJp17Nzse+1VvD66Q5+H
VMhN2fxA17ymj3L5ONGxtvRc1uFOI/54pQOot97OUUGzPsgENOUPFdxEoxKxpqBP
HiVlK1IwivwJDcrFXlkx2nu1aYVrXfoY/34TNAJm+y8ymnqtxPErWozlWVA+hDz5
FGpmif1620DCUkrvsLh9hfOZNhz6MxAwTUPHCV+AbdT4UVB3J2RYV+/wKfy+vD/Z
r2QV5uKXVa0HatcMwSz6sluDFJAkQmvk+d6f7Z/Dgy+rvHoER02rnfVs1bsJK8lD
1CvpLxozfwgOsc2YDwVfiJgJELVTHJCYgwGmK6oWTHEFEzNNImmQZC0KOa2I9+uj
lm5Vl8gqoXOxBR6cEt0gq4DeFWVPbKOaotfojTkAGiJKLkXJUMq/JHba5pCvZK9i
n7DIyBiZI42fFe2lR8GW4opRhzR+GUkgZ9gVcuecvWbIovA10uTDN5TuFqdMplFW
Q+hlMumNEOXSm26u2ZGkmNcjN9nE7seJ5v4k1QR7YxEEPS5lLCr9XXGLCUUJxG+g
7KZsDMxKoi3LrpJ/8/zp34aXnfr/Opx08sTbKJ7V/3lB5J/dqqNh9r/qelSmEVJN
041R8qmNbQ5ft3KXxM9XF+WUcr0/IrK8M2lIJhrRWh0L1oPKfRrWt8fSGKLlrvBi
Rgf1VHRZf6wwmuUobEsTDXdu4+US/xbGtTMl+PGssozCKuRkcOy5syoRfddZA6aw
Vm3fs7QLuiQ8vg+2JeuOV/jleub4P2kD6DRTbBZL4TTgk5llTqXNqgka6/z0HWXs
sArqF2Ej/hCR+kQUhVYVNwBbrWqkZVxx4r6ILxA3kJq7CHH5zx41KOzTt6Mnlb6d
1e6n+Ynqme7Rb9olXn6OiNDsY4qTLte2uNvi9f2tMq4cO8vdkcAGYT9Cs2SCoFQ+
Fvcaoal0qOr6O2s0voTdXpAYRJpOVgoNY+7FKIhhhYVJ8fzTwvpil8iYlJqRoyu3
1a3YSIHeDrwQLKC1jcu5z867ju0xSWUfnv4KEahCsXcFSo2RU4s1BzTtzhxel80e
58yoPeVnkSm+9cH041/qlYUWp9qzPzogEL6l6dfwQ2Z7Ojz3ifnMtChxgOADxQrM
0yT83fg15GzgEts0xA53fam+BGO7Uo1JZMP+cThvz+zr+Q+gCRmekg+SvNWA1uaH
MYi0quI5rj3XS7k7EKJO/jT0xW30JjKG0m+gOnGsegjmTC5ky5tg2zBl7I8Mg8Oc
uoALmOrHzi+HdN1hHJlzxbZcdhYLYBYA944E8/HtHq93S5TRoaGHxoU+Rr16fMZs
SWSiL00oukgTlKJjFbj3arcfBdmeN/qb+f6GFeZcJASG27p7nNcphMSWMIFhXSqQ
K3Yo7GbKu2TlAd/NhKh0ch4GHznx682wnqxjP6SBxZ+r2vbpx0gynP4HfSfjTjVr
4caqL5XeQfDwYtHNoO/NwR5u9jOD/HyvGeIJmxlHnOSeGuzmqd5z9I6Yb7ndqJ+H
HHYtsGoADIQMMwcLVWEqW7fBZ+b1QBaeF4DHpofWkRp+PoDC2kC+yHV4z8XGzdjx
YiK8ZgHlm4K8tI8tgCYk9uHMdmLpcgUV9PwAdm41w1AkTFpK4M+CQo3vfOBSpTfu
e+t4KrstsLWZviht2XtYgBHfSSVf/4l+YzHXLYNDxctJuK6M1b0ysHEZEl+6kiGo
qNGNtxBFY+tgcw5zKJpKL3cK8TAeMfA/4hNgMYSkth0TYCotNRY3TxUDPCfhA2Ws
etuH+sFS4xG2Cuz9c2gdxiQymTI4MotyriLo3g9eafkMNF6oT2aCwjTur0VpcG6y
ezjMhw9xJQWvyyC7zNddheTBjpl6WgXW8Tl7VkrFMav/TlKLXeK7kE8+QPiPYqq4
0cRn7TuN/ptB9idtx0PQ6Zg+52ZHjcA5YbkY+ugS3Uxa74r+VvmzNYYAYL7h/T3K
Rjhsjm23E5UfLYX5RIskRbm/8xKL0QkSd6FLje09eEX/TB4RI69aCrCTzP0bxpQZ
+x8/5dE8TdUfM8oYxSM05ss8yCGmkHedwImrIPonq6x0SeDF7FC/dphud9CKphh+
0RHOQMSWCbtX1KPCR8DkGHSz2ZlkOcBE8XlkX5yoFOVqJUTFq6CNXmM2hH7WVe8S
kjaYbHsTVNw8idqoGN11QLYHAA4D9tRikD66QPs1xtLhnLLrdc1CkNs+dN2cxkTf
LRHtcQPaagUz7cnFH6iSscyUglpqNbQXYz1E7t6vemECa0XPzYTUzHFNUF1NBgno
n372DZ+rIYPCK0UFYFpLMDktWYU94jTUtKTlhuxcqgPMJiH68hlOX+W/ZH7+MStc
WxufIS7JWnxlWNTiKYAa6lG/VPkPm+i5MwaLszpCkvcqxGZqk3cisQ9tMn3koLw/
80QfpWoOF/5a9l0OWrrrMVovHg0GYtNSwsRjakiovnYtjv1kiubLSP0ryD2ubfO1
msIZ6wK1OkBq7sLlEI4EZo6qX//E5qpLihfVLeXehAIAGGIXCvZOJ6P4aBPyqsPp
ShN/FzkSxe4zsPouveMjoIN3UI6zsHH6ZP1IOH3prQ9ebsEMwvhyzhTB5yTlXerD
MJA37sHmss42CS7q2n9kQoFdqZIM6bGUmuxcQIagLlub/IQz7p38KFYB8m5kfLFL
n9EVKP/nvt7T1xyjBbS8FW/nRxjOc3ruDdSZTSNR1r3obqx7s+1bP3BD7dIu1Im0
MuJusy2xAt7Y5vyXuJIOgmcPiSuGodiquJJSaXbU8tliURkwNFj3OXlk7F3Ri5mC
R05MAQYkqjhY/vtaqDGdAc47mR5/RheMOn7ZPKGbjWKWQloQztXXnaj5f7FfNURv
6Fhdu/YhlLL0YXQ3ri2r84yOkde+emeY9uB4x8u9dqiB1mTuYaxV6fKcBhFIVdfR
HyiXpucxHOFbuNmG2jc5hM9FHqPTKv5ICyf8I46+jONkER4lNBrz0myQdwk3AFiG
y8fxZssrNnfSYXDXCKlGlhNWSwSZqbfNuK39pgURZlzLJGTDxRTkqMES6FA8TDdM
w2zwx2LQI98EfjPtQTgOuB3Ck9g3QLQsSdeVlnp/Df6pWLnZNNYAskS4pIA/0g3P
JbPB8ex40v4fWfBcwchN+ckQPr6rVCgDjFA8/OuivH2W7QTcjoW1pYi+c1t7YEei
FNViiD2WiMOiRU66Ey/or4PDto3N75TSe7PXDGZElXAaCVPj4oH51JDT64AoI47N
DwSfkpJwhDK2DgG0AgZT1XPLEFlpg8NSEOAvpuJmTKG/3QoMwSfOeulUBxSKaUbQ
a84M/ycKf7PZKi2JiQ/sX9/Xn6lABgMQOgp8U0lprWLC2ENuu17kVU89idOgR87k
sHAGayvY9cWfIBGYt5wVGS/aGSHOpX8tgZ91dH8/i0N4hzL23m/AD/aRTP6QnZNR
iYh4G6ddMwjqL6OC6gSJDn/JN0Mr7W2VOHRnXcAaAqDRR+Fjvzy4O5AuITOIjF5h
4NgSR6mL8UXmf/Gx7n7el+1MZH11qCGzoCjY5LZOXxrp/Ep5Ywwoc+q75P7sK1Om
+LECUgTyyfDcxGKaSUGD+GvUCpYSZooO9x5mdRnJkwBI+44nqka3wO3dDz0MANQj
1YC1OS6IMS/MGXpvZwIoM9vDRH4vkve+YyxuJ/uEjT3H75T7FAtIA2pr33TAqB8q
bZwgTENQwMUqgpeQVAxW5oVeZ8WEKqgBfnrN3l12QWZzKOJtKFP4b6sV7I9d25CK
f/1h7+S/WFyQePICto5UQSA5JkrNFOdfT1LYc9Svg7zXJH7fg1/2dOIb/JB6v+AW
Utw6xYapicSRpBCNei8MsF+jX3btFVD6XQyYcyZ1hjDiJe3I+B8Iku1GpBnIiuqR
vczj5gYf+7yatzXdbimJSmGgxAAB8EGk0K8qzNbo0m/lY/G68V9h9yGxLWmjfkWx
srwgeR5E5S4Vmgsc20jatajpFYM976007X/j+YYUxTrQ77RHqbQOluraScO+fs14
64VV/3FO1t06vWmxaYMErOhxT90ZZeG5de5E1aScHlT41GUReiQMczSokn1yLlz0
a5SJAz8EHBgKxgzrtH+qEGw2ie1WUzA2FzmxDTx1jLSQAJs7pL0rIe2ToB0iOdBD
+Qf3/tvTYHUMAj3X/k45Eqd7+dA1XIP8ElirYgzIQU/JgVQ+RvCRxhe1TW4rd4E6
H25GarCnWgZ3xJ4I+GyeDEvcOeoXD5ko9qqFJ0EoEJ6BnUlscOY0X9YxxHKCJKuT
/Uo0OjDKmdmS1dJk/l8WGPd7M3xwlrlVkzaDps5QXjzCvokaZ7wbrjmGZnksIYA8
UyArQVLphjLGFk2wP2bTH/F7Zc14A+m5nOubv5FfGODK2YHSnO9WE+P0zTeRbqyl
W12umIgoLoeMqaBdULpNCkepMvK2KfVK+gXgvM0Wsp65VHlvZDFFU9KNFc/szgXi
bCQpFUsHLerpvBEHNbKx+h2ucomyPReyjTwzllKzbJ3Q7Wtfpta87qY6MSx1qY9j
YG1TpmybMdlWDi13Zu11Av8xkDmKHXDxjKGxBHZNizhWQSBGRD1oIEgE8j427l2m
Y8Xx/ex3Nvum8mid/bNPo8G0OCeuD9+4PFmcc/MHv5txtcl7rEWR6PQYNEy9srjW
ISNwfPdQ9Zqqd1LiQGZGtPij3f7UowJisWfHXQWmE57VTT1Ny412ihdGu5qwJSmz
JOVp0UpfVnt3JILLc6qki1nhWs3wct2xd2i3toHh0ifbY814pfY7v9JuCWpZJ+OT
GXI32IZHsEHfhbJrv710B9T/NPCAML2wxh/iXBOazeJGxOSOcvAGxDI2z6AKlSND
BGKvcD5tuKHb6QKZQjlUy9iabJSjsxxfFFuTJA+83A/79dG5yJuQhN5cwfjHeoGU
TOCawT8TJ0Vh2epsD2R8K9fiJPCBC4Lu7+sd0f9/YkiclChBWCwIMBsHtS1fD+ys
RFfW04teDdzRD6WXWIjmjdUfNj/blXZMvxfMSsBQdRbLBwPhq1EAPv4oLbR2pZKZ
bVoAdH/R1E5NYzmHhEDQJD/2XeHeaODJe6KuFXEYt7KieAutBa4BSz62Ntj9IDQd
KL1HxqnHyaAyvZX3ctIndBa77QwuuHJsJEzWhbxe4Ke0Xa8TfcX8aZG1qsdHrEj6
i0KPhKfGrUXy3sBgEgY7eWL8rC4n6+l+6j+ZKKWN3dq+4uKe8VOTIF/R1PBBttTC
xr4nB9hWNPCLADtWIFIodaX4IACKQOHqmP2Y0uncfbQ2Z2Uh6nO/eF8zaMXs5Bj6
QaGCXDLbvdTe74E9cgiHYJ0zwWjOSUwYZxh8/SJpqLsRE40kbDnNvCRZra0RwroG
VXTwQ6JBSiDehs5Qj1LQ+79hZ1qpk9i6RKWhiE9e+FokZ1RPuS2/Tn8+EHvRF8ji
qLOgGtu/wvruU1YB/az4iy8u4kq7Y1ATGaKnglzbwT+SdIlCN6JHuxGiBI7geUW1
XgaEKHsOSf+G+OLYZdNb7xzwj+HwZB9DO7uqEDCpSMcraABCqfistjHeXUjm1qpj
admRfe/GmjqJ1iorFuH1ethJq+iPI2UfYjcMXgtlVliJ2VfmComNsQIed06YS4OY
sq5c5uSsAq5bUry6KKckRGOq3IfHF1jBwucY8mMU5t49noadQjokENQ+N9+6vCAb
ofehLTi3fymjm6vuUcMbM3JM9EmC+y6VfCD9RaJ6kThyTPfl0UOkbvXKvTHUAW6l
67AYPf2I4qlgByFWGiFzb+YncHT/wm2R1jAuAzBP0h6wFTn6rFgHQ+fShI2kG7zQ
l4Rp/Py6aFnyJJAw/1Y48GKKfiA5y6ykp2VM10jtlf7EqEs8ZGwVdirRPXwy6QD+
B7fvcEn6quOUtawZ4hgtSXFTx7Fc+r1U1YRRsexNXlaud8euwzUzVvjZnNxbcLqw
jed+o4na297I6Ovz0+p6AZdokJUy2C8RhF+q8xkR1UyA5H6DoTNHZgqXpBJT+90E
F+LMr1QDf649D3/WSkiobB/jWVgaYBf1qZ/GytVO4nzTmru1MLeSdNkFW1vibeZr
TNplh+DhmUCJS4gxiFtgs5Z8CFqfZmCL55fWerVXzWcqdevxo+ktxNqxaWuKg26A
jK/zQBZRZzhHNz/stb4OdYQXdrdAtByMIcFpg15K923aogXMDI8sHiz1WFEWEtN3
psyN4RpeA6XOGrQ3PabD4UgVGQszotKbU0CMvb43r86P7zy0KJo+MiCJALmreZy2
Q+eFgPSviY842plsRfJuDqCKTlEBWFTU6wuoXWwvP50d7k9kHnH0jlDlBHRcKX+R
zOBt2vgJb+e2IW0NUouxy1yw6LGw5VT2pFrGg9MYPqdxj3027y8aKJoClDM59Ffe
cvRC1U9atIBftyHkfxyqiiSmqic9YNIMliOqOhPyurC1TEiIOttr3qWLgsNbed5h
zICvJFkWtm0hgdlmnHYOyu3mX2ZNyouPmQtfsPl2uZ0bjKjHKdhs1R84cfl+L2aW
rpbhWgq5a5w8lM14yJBsWAUrZcbiq/H1QuJ+BTwZrBtnbYhyFW5eckRuZ3ezperJ
Ia8JkTFFf9rCVwfXJkZWX8NBO7gWjwnokGP5hDHjc74j+YvvIGl/T9TrpATJVJLq
6RCN5ScsLKy7YAtvFAXjFO88GFOeUGYz9lJ4DDKmu9qVLZ97Q9d7Qdx29H5LRXYz
+vaW8koxXry1AO7oxGGTtt9llQmWnhOOwDP0EAVrjFYtP+15r+mSO7N07+emTag1
fDdNsl/kIIYbnXCsTlt/KmlSTvcTcghFJt5ASF5tfrl9VRgPxSpn8N7BhTsUZ2PA
L3nlMyjlE9XqKXzFFm0gIyHDTZTdlz9MmpdbApn6UkyK9Qnq/1xz330BssKLM73o
h1IhofsuQMeai0n02o498GBJHR6ITYlCuaCMmrFfv0sfdYEY7S1OwW5sRmvNkwpG
Polr+mQ5De94wS7aOOkutKdSlHpN1TFVA9r3k6Q+34isQksXCi14eO0l7Jen1u8V
DqxLignUe5xH4Ah6ZdQ0l3j3THI/gdgMB+we79Fq8izLVN5064TH7Lj9Hn9O6Kyh
K8O7Ac7ZM2HcW980uzeKVevxN9qfZ5wNqcBSOLuOntuhBxlSzCIikvfR8VUTasjh
OP34/GqzUGAdV312plqdOK5vZnOFqgXyCwkD04aLh8Hm9SvmziM98Xp7F36FUHKb
zXmXoyff085VT+8qtc7LU32u76AJFKCFopATLT/hSAwO8QtK2pcICcGXnXJdRk/j
/5zvJGLvNByMCi6MYsc0GRRjU29S7jVsyt6ByKcRUO37680tbkmZiufSq1ugtGQ7
VYx84f+++ufOAuQp92R8xf9rWmUXCFX0CGBpz1Y4yKVbMzV3SIGAbUjQvk3KE6nK
QGy+Gv5kRttAzPklncReWw/B9bH+pgnNOV0T8a4c50ta+TvozS72NVrrI1G947J0
LcT2lhd5Dj598jw1ppzJlIjkANlaCtl+/8sSm9OoDHo0crUGo32OHhfebp3uEt0b
WXwH8yzlHayicUstyKGXouUiKdCxLcRCF9bgeTgUJzF0FKjK3ljqTL1Jtmp/8IE2
BlrxKi8AQoOa3mcnmRecuDZFtOCzenWfDptPjT0Lt3bQpp9+0h5MpaDcbfVmCpYv
dZO2O9tPeT5YtL6PrI4D3HnU34bc1IxZ3bBfl0/ZDOdnC+7dYhuKfvX8wlDx/c2t
dWJ20UzTNVvq4XeaIaK3zZiE/oQodu3ThJJuNc4pe+g1MYTsyG2mN2TvdzueusuY
+7zQu1crrdgaMc+6o0uU48EywwKe50aG4Gy9bZbQejqAJ696kof0fRxiM7t2x6lI
6DWFy4Dk6WN9Q2JE/FkNvNNwoXpaUoAeIsftmlqzhHOnWMLqtQzqcqvCQMQPiSII
i8fzWtPuXvVbfIkruzWtopvc01N4Ov2PS8hR2sz/buB0i8rAG2eW0jf5dFrdqwKs
BJiOoDGKlHzU31T3ezX87KBNn6Tv1ojgYSJ0ri6VsC5GZiucQiT3C1HXFoRYyykv
hgc1N6JdGTtl4f8osmVb6rQDuyTW7LUaLUuAbXpRv/0Y798L7UuykKSETNAqYvhp
vngGXE9VRPILhyO34YM288WrQrP+47M/6CuVVUzpjpRIym2N3g/MCTUxJ9WV4SwA
9ma5J4Sb7w+u4BDN25sEOKP/OTZ2EdRfTfTOU8HCnJADGwf6WqOi6o0M4Z45aQE1
aVvwg+38562NBPZCnBhqIf8ptBThBdTvTxAKttXCRTqVxg6cSYLa995FeooFSEa/
eO56uptOiz6LQHO3DqZF15Va7pKq5wxx4/mYOewPPmtFRSnVqx45NYLxBwCr8ypP
7gGjLQdt+/pfqPkEsvadhlaJMiSrY3hOlZu57XPZ27axqq/9d1Bw1Y1rSJtFec6T
ruXSZcX0TjK6KnBuUysNSOw5ILGG1AoeZaP6WnuQh7qo9nuhJ6EZEISG+IC5alaN
HlP2BL5O9thn6FNIy0tqKkUG186IScaUp6OJfzvpBao5mLIVznpTkrWbF7slHUqU
0VihiCMbxDDpYxKsdBQsjoOlCZLpDgIDlwbNZH0BXFBIOmBwvQtkWpsFzE19Oq1g
335SbdXgaKBkoBZi3oHbDctZkESik4rc9KggRz3Hf82cKaCfkyaD109nJOkfil17
S52Yw4KY0NvAuhSg4lozQ0/Aqh88NKk6ZrCWB7Of/PpScVtIYr9O4Tm6nybNXhiS
oA4zT+fPNHy31dEw/w4ViUzWCbxAfywLf+3twDMrOeA+GsxxYKHEQuqFN7p0dCew
RfU+ek1JyX41I+kNt8yF+Xa/H/y7OdLeFC3GLVXdtMLJrvvGzXuOACAKHG8QO6rM
uALsQkEYTBUxooRTmBjAS6uWFcJ27pa+DSYpy/xKej0ZS4Ih+HLA0k5z4a3+eKKc
U28deR5XMqZh/F/4I6TMxa8trEsEt+mCyRxuxdFEcQNvhW0QhwLIHo5zvABH/e3/
jUXIxQUpi/5QA6UBMqyZeVy23Nf/O81s3Olmn2C58IF5g2J6mioEmAiZTHggksL/
sVtnJSZhPQdJ5ENiYyq7LtAdhxjeqL7ZeqrjUQWMdqIalbqdNy1k/T7fnb/0sQ1b
ZsFuQMloQ+mLbslrTI2B3hj5+TNWeEaQCBSHSxhGGEimpWShgPxmGtKZjSOtZd3t
i9ZjpE5J+LulCfgv0WvCKG+0bheF5Wdzajxi/Iv3wYFKnvq788cHGLOGSvAs95IJ
JwaDIqaAmkuOzdv8D0GBkQTfi5eryKj+8JgwN77G/SgLRZmpL1pL9adS7+lkpOuD
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VEG1l3F4geEptZqNoe7u6JRdpeLd/+C+sIvfDe31HCQiL3kp8heYTIjqgziaxFci
r3BdnJzm6rmEjX6IQnsFWYeEOSPdJbBavKp/YN3QLJVfkLT6nbj29hGykwIe5ub9
JxWkE2Va4/6ykHaMTNMBoMMTc11kW1CldFlC71/vSbZpgAVuT6qsafhd7/0zHxHt
MYor1xXUcDu5kL+1Bl/R+9nB35k3P0Ldtw8XLskAO8xEK6sYKdKt8djAKVQjSd9G
kjzuVg5btX6TJG0NuaVxu0EcxOlUgmHO8DaRnhdLq1jB3RPzNUv/08mPyG6+QPz9
CYVzC7deopmdDChZZN70LQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 20400 )
`pragma protect data_block
5cHqyACFEPCYc31ngk9nQv7sjxZIiqY7ZxjLhV17jXWBC/Eddp71NFLdrKnHBvYo
QY1CpkD8Hsu3xdSdLCkY5hx8e8WP34i6Y+SLla++fp3QJsGjSrYqnVqKKHEUazCj
cQjJesmh0n1qtdlPhkc24gQeu2TZVxTQ/kcgo55sWccm1zUcFCEZDJJrcQdzmwuT
ehSpI7Up15AVm65y+jqSeTO5Lk9esW2vdr+r7lNVCLz8LluR5ameSGdjaqMGLMjW
FQPzSWmh/0J8RLyCNEc1WOXb5bKlHYLV/tB/asUB5Z46KBRPEMl2xahGd+k/Qq78
B3o1YBpqVhk8GiTBZZRI4126KrF/BSnye1tEULxqM70eGZtUfVktNDIuAsICduqA
rDnelOHsMGJaBWKpxYzrOHS5JYs1sl2m4SAYNcOTIsBDuHc/3zo2262o2v5h6NPn
kz3+eXSkkMUN1Xo2tDRVcAcHHWpIHoqKlI0wY+SPai8Z53Y3poyr3KI/ijfidz7n
h1KPldYyrHXU+tkAMcJglYs8RSMNsB0OvR4s0+dKM9/6fTdy9iWeitRenhNjkdx8
r4Np6mXGAJ+wXe87GJjTRsk0mMTbzkdNzZJQOZ6q3zR5kGHVMK1Oxd7+KXLdSQ/B
kAzlUc9sNQtiLsKiHqLF8mgr+3gWPZXRWwFtK7zsXHnDl6yys63x/Vwy8vGy8TVq
xB3gVApVSXlyhqP0NqHu50v2HpZ87pge4iVWOmF1o44XiXc+KUYv5PAnBUHRMQn8
wdzyyff2bGIs8LMEey8zqK948dvop+wtoAOrg7kxs7egIEheJpVEd+jUB7rPBhDx
HLY/yu6fE5luwA7gLTI3pNArUV6/FzHjl+LcMTGYMEXg/YNVgr6GxISUCwy9heas
acoOTuXm03ACDXsLBy6+1j3/iLMU5KQG1NFvbrwkj+ZI2SNYMz/y+5L1SeEVlbV1
rCOMPW12BnXspjlvyAB2VgnAnnNpZx0tGvOnaPP7rAnDpfVhJHNGtqN2dwCg3oBJ
QYtGEcqL62qClytod4wuz4ShfVTFAU1fVB5KBfKYOknFkZP9J/rxEj6xjgNgwV69
KN2QenpN/Bkknn/3L/8m/ofXTHsQvLhP7fY0vfdq5HrOqHfy8DLRx5fi3ZzwBb6M
H5V82E/Tc31zvHpLukWS/qju5XHCfFvsfO72KExOUwRIHzq6eC+F1IknZo1RPxLq
QZ86IFNQiqEjSH/LC+qMU/eBKOd5bQ2IIUJaXDX8v4YNfeOzhibxCAmokAcFGmKK
tTjKzBev29g+4AtTr72VgpMJ7O44VoEFEjsNUpGt3Bxi9g0yH8VtllPUczcdko21
Um+zWTnZQazQOElSzEQRmzGVhgEoP7IY4vETJArjGYFUZb4gryMc9FNYb4eINNF3
5WEJhRsHNFZaCZP6IMspA7rYMXDV0+fUfNBgixm2Ef/GRpXkLS7SqUtFPO8fyhd+
GlIYBYK6392oz3Q3c3hvryouI1lX2FFwxbmQs0bGniYeArKR/oAqZqecsFOCyliU
r1l1U/fnLme2xIqrexuIduiuxnfu/2qVI21UCxIP3hTr51i40p1hL2fBasl4RzT1
nv9CZyDZPr3SEpn/rtkw7iAL3eS3i7fwu2dsBYLezWAKeaZOODWgaVodXGJ6ezkM
En2K4JdsOF+bQ9lZJPsIOKphBm2OH5m7Ggirk7dHVfEf3pKB+nY6E8Ff55X3wprl
ouzHz9DIjlVNILGSPBC5TVSde61HtU7VrS5jJRs/ccbSv1K0UMLmK3s4aQM76Fjr
zCoO+/g7s6QPhOBJ4/cIC0RmFPqXTRi86Aq/ThgOVxK6FWDWQmRW5kx5WyHzRyAL
ruBm34N33lQGJXPExSht33avI7fB0dwEPXTaUin0mBnTSJ9hViZBgQssXAsv4skS
g7Ccoyl2e3bFtiECzqY95AO29t/l6Nh+nHlAja0KAJn9m8ThryxYI6nJ+Rxry13d
3+kjjhgFpasZ824W2QgBkidRO7VsAlZuLh/d/cgIgaOMjzIgPCk8+8587GXG6H0K
XGkMaAuEzrJfsV07N3TwpgRl8mnBcQUk8FXN7G5IqCHXG+tP1bXzp+9Nf4egzz84
HJUYTzxHP0/Fm65ygmVxtlNhI4g9UD+lNLF0Pl73AlYfT8NkGjOeGg4z7JMBQo5P
YiPqXSZwCHKAue3aHbUEriQVmcHdFdT7IlvB9vcA+Ht/A8UFrmQy1q8FPLlIpLA0
XfnEVotwIwrVT8i9z0bGVlfGxJMbFfbxqTh8eIxTBQFRvNHdusUSDBSHpR8npL/+
lPTFlAA9++oV8qrhijeDBrDmJkagW7bU3VNMgkgNGhzrXLwN69aZhzO9aO99uu6a
/6+gC2/+3WNdj52uwrw2VcUegp4lC+YTITGcoOdXzcNgsItaB21uFBP/qeMH8gI4
qqbRDI6xEXIWau2XHvkR9df8t3hjV0HoHNuNzGzaJI6B5u6nqO1FuUeLfn8AzS3I
wj0ms+ExUvguStZJQIEAct8zDa+h2Md0F1bMmvPv5U0lcymcog2e89wRhlBwdm/v
UEt7ESmS6A4JN7fryrDswty1UYrazP9/ow6bRYC7YB7sTz/GKc5UnQeYT1gQgwti
4utcrllVuLqTNy+2Zl+BYMzDB/ASsD2YwU1GtsDATHapLV7Nj8uQcY8U1NcITid7
yZsFuKX0pbBR9LFS9Zq+J8dF9FbfsZqZ7H0wKQnjgb3ezO56wiTryMr5gzjch83R
B14niU9E9JrWmTk6gfiNwN8mUYxvST8bGMxgp/fF+bTLtLHDcM/r2XCNyfoOLI1U
cjwVHkO4iQ+EJp0Y16goTTreGFd/EfbxvMdeOf41YqV5a4+eC9iP2eDtzjcCoRrV
MhVIF4szSYWz0bvMNWObOPFR5xIc9uc8gTv17YFg/gYuaNcMhF4jr76BR2767YrX
9/Znn1Wa6bDY5wa9tJoRrgdqQhqt1L10ckel357YZYChOpl5JtzZT+TwBf7Y3TLc
fhM7SQQ36xFN/5+EzTdRyQhQhIb6h81HZS2SIGBKeAR7069CzTdPN3ck0I2P/oDi
X0YVMk6IQgTI64o+4gzOjNX/GirM8jcFcPWtAb+3/cM7Pr2C3hLUDcv3jZDayxNP
odJPg219DD1TvDyOH54V7vLYBFNbDXA4pxMlP31BukO8NhQL17n6bi3UEpcY6ihx
Pu4nspcyY5Ixq/IWx64M6DLEXb4D1Z1xaPG8UemQGiEUEUX+P/vehBTS+GtE+971
+ubuQRBHbpfF63ZNcgLbcDkEcXBK9sIzg9RsSsIwRRpajT7PR7QqyjD3ZAoWLrBv
eKaAvVkXgNirgYegyOedQ9BKwrrzxHsmt+8Xe5vqUM0/s/+S1t08OeDsRq24i3hD
t5xUYXgQEbL/szwdOAJHb4Fmehrr15I6pRifk8tCxDeYdjS3qwnc7hDjAhjY1r7J
mtJ/O1J+zpDsivC8505lZ1EEr+xN+WlUyHf2ySwEA9gXvHKr3DhXS9S1F7ZWxjLU
xYYWfNhISSt1llmTjzeuNBpvXKI0DjGHyoI8WktIjLH/ICb+LBo0hp1Is3TOJZ0j
WFyGi3iYLDsFQms9jbirewqe1HHxX8mV/83J8Jd6iZfs/nJfHnYfyJP0fHeMO5/Y
EMZPICqtnJdgb2XcfqXGj3ZA/JZmtG19RrKtq06DBKdb4a4FFIO7vBt8etp2TReU
my8GKGnQFvUNSYppIyH84WDZOwAc3GcLg9nprShvrpifIUM8k6rAdMZlQkQiUhw8
yiMNIo2zyPQj9NI4c2fGvUs02NR1hovDFauHv7xGBLuIoynOKLZV3XzFD3k/1O1k
9n55UN142wjCrGi0ccPm2M0Uo6F9BEeGbZ8sv/7U1IkeotfNMiRqnaKFsgiMQvpX
Siq7DvmmtBD1Ge/aTX8Z/2j3XgjFumEMofPd2Jz1SCPrIygiSskWEzDrfOTTgboV
yeV7wmI4ah3I/9eHfVrW1AQLsF1LoDlTSi1YCMutyqHSXn5MNPL4eQ+/lMZsvCUW
OU1OrNNx4CGJqWXxIwl8xSTlCben0lFXn4LBLxxcQGG2Q1NMqjJZHx3qLXkr1VlA
cHJkyB+OHGAf9MMpzD1gSLcfc/j9clqNcmv4RieZrj9SUvwP5A3wgTOAByqB4+Jv
t3u8kXY76WtHP5NMX4iRSs+9qO+W30re20vPg7eGwHleNseZZdnpZJdNWDJhY/Mp
yzDLKe5mfiTQSXU5BHEjTx/yrhxBD4K2LnWMmVybT8nuxIqAN1dhpPumrU9ygutq
mpOidAB7uKRDnI5rN05B8PqqkDb1gXOf73P1EH7fWD81eL+sfKvTIDs3aoQnMlN5
zoAB3TDpKv7F39s0vi/CZbpV8TECW2sdHgL+smI/YLj2TIqmAOtZNWhf0Z98g+yC
Z0Qr6mUAsWqf/1/4e598Pt4rizFOTqAHmOJw5+8lYLvp1yni4nZ3+2ld09rGYV6G
rQptOPdCFchQBZrZwEOX6uy0hc5+uAfsmqL3fCNEQcpDCh1X/rQcbjhcMUNK5QkE
Ru3IfORTCZP81ojNIKxxmAETzMCNKcZmW4xLzPzqBEzIemasamViwf6JJhHrHWRS
MONuXtMQwcAj3vRdjtsQkJ1+gGBYoNeqi8t7ex5bBuT+J8qalZVZAdSYhWS4Pmh+
ie1wCGnpg3LZn81Nftejc9iKzxSmTNgemOOH4L+lL9oTfOxM9wUYirp31etwA48d
uWnJX0lKpXn6JhZvXsWYH9ai5F17C6wOenuXr5nKFHcST3DL64046/+T0A2qUUBU
nEZXnW+jGG3+aU1wRBDle3XsVDvWnCdq/oW78M0SsXOwWLG9IyezYlqEXp8PHO7N
PA2n5k23FPMSmOlFL5jbxgo4OBjCCNgTseldV4TmS/xx+BMlLOXdQS6r2OqXKQUb
JdI+xD/IaVQ6QqCMGnLHIIkpLqmm95Q+VkNKhxxdbFxJLqt/0wsvhljONMYoElY5
OG1o3uOYK5cAyYqhsciu21UMn9oDqNmdsESK47S6+CMKQfwVBxvT9a8Cu6UAQvtP
XD0OChQXFQnYDeEjLhkOvjAhSa2r89FeRgv7WGoMN3/kY4RAyNR7cBT2c3PIEfWq
ELhBBQ+GjzNSD0zuYrI7+tYd6G3lzEmWYvckcPAgxepD+0fVkaJW858J7BKxdMkW
sfjfnDh4wuo5rcMbGRcVN8co4W51HF0rd5ELpK7B02hJbXZyCCN4392yrJom+aik
14qaea1zHUp61nVohICu/9jrvrmd3TroMotnUqGiQNvMhjtX/Q0CKCceUTGQC3rE
CEMj0WwJ+zwr7JuoCJ5b3YrQpNRq4rrjl1IjlrU1nkXNcZHB/F3a0qic9/EFOq19
ROkeR60c66BNCYhVAOVlNVnDK0q7tMwPh/JNIKpj/PfIJm7sk3dohtOIZ4i2FZCI
Vn+YmTFN0vlk7LEgzmes0rHc0VNdCa0TvSBfk87tGEhSXVZ9MoETkt7lUF0ZAyJU
QyptQ7Sdr3LKjB8YN/OGMujBv9iniXMf1Z+IgHZSMoM9A9FnEecbAw2VByYn/0i4
+wSsQu+WGjvACcvvBvl/ZiMRRfY7i+tpdLdNcrDFak69iwpk3TC06Jlgc09EcNhd
KO9eKl3ojVEuQ5DXOQLHXuMLQqb2mEGaCebGTPfCuZi99YbwYMSKJZbknqaUYWeQ
10LsKddz9+DlDquWPaiRSO9JwpIllTYYP2M3iHQ+p6bFaPymogYagLW+2xOWuDfp
I70T+GY1HzUoVfiAlMqPRTY25psPKrfciTL+mBPmtsrqVCgtWFx3NFgP1DaPosOH
2bMV73XiNzCe5R27g+OVX8nuhzy6hEWM+FVOUA1bluml0M4J6jwy7lE+DixcnxQv
lL6ST5CAtVMR5SKefkJYjXAZr3UENXIMQ9jysYoc0mqGf7Fk5jeY2SU40rKtjasN
2c/SXMQgAg7oRTDH83XyCYhJDzZ4BApTVMH9nmgGZyF0NLVbrSUEWFAp7CZiu7ye
6vrrANvCrRRjYFDr4cM/4ItvkUKlMpSqFr0M8pMSUyLH3xV3N9R+fbmlutB0qD+P
jbPI+yzPCjFAcLwiFuvmV3khgrtSltoNmuPXDiLp7qqd7ModiiB5dsUv+dbgj1NA
tIIDefEkRdkpGtSIvYS9E8oSBEviAOmmeDBP7ndoX9gz041fuj/WSctzEtT2Sc/1
7lsOooLJfyZkU3KyOVCp1Pel3nfTubPmTRThXxny3//Ddz/fLTOwXtUg6jOxdgJ9
XcdJU9sKCboeiyeGxlhLpTrMzUiGxCkcqUrEbr2wXYfT+ECvrlUyA25mRHABx63L
lb+9DijhyjyrzEJs8iM3jOBR+ECIweT7YTYB1RL0+zoBvpLK5+yHboqLqD6eqf24
FQonRpvyPKBJ7hlWsnoHRI0pqTsP18yYGihkPbxfby7FWMd25mUHpwqHutNqOc8/
LM3qAnLmJMYkoAX4K5ZziqtMXmSsmzvMIFkDx1a4Kz9LiajoPhU+u3ya9E2Zv5nD
gYFUFvpyPWpsXXOa/DRWrF3hz/yeklxApDZhlz1ZZ8vOqQp5VQcp24MtMsKxg2zT
RmxqnNxPcB5SBL021LW0TMeaQ6fifaR7EHLGSfGRJUoo9XW5lg4c5VM6qR06dCjv
xgChQhN1gJrphLXVYu3B8qgGmlmt7T0d/sxn4q5+BE90JyAu4Yyvztaf9eEdHP+v
QPb7V4XITtUiip6WP9U4trKT7bvAJxfCozv6HZytY8nrD3TtFttL3XBeupYovgoK
8NrXgLejcbz0AdssybxnFfCL5Tmsfya0GsHXdqdWIrs4LHgshkYweTd3UxNBjbsK
QOYO62HXrQCtv2j9C2c0LrvieCteXvKSFubHPynKz1mE+SkI9SHz7ItgwrdaUo8d
Pxn90tqQMl3WJ9DwcxHD0T8gTTWvb74m6yoTw7umbEtb+5G54uc4YLc19eiD/Ew2
QNgTrH8PoHRDJzGEj3oOZs0ZxkVs9yoO5JN1op3UWufIak15qMkdPTThq2vxogUB
29mZJrZwDvNIlMqQVPnj9UMwK76XQ8/qaU4b8V/aXI6J6ifrvZ8CUSorwSrZ6WT/
+sIQfnF64UJOejHk2OPzgZmGvPOnSh12v3Pb8hlfV6WXSPxPImI0Ek0xCKOcBw43
ueIKArma2cvhb9abLOCxYwoGRj77v+54Ow0WUK1U4Xo4qmP1AvFZqPQzVD/7fP5I
HStxRElENM6NVLU7nbdsuY1SPZhaqdKhtd3sqxRJOc4J+KGMRK2BGSZT/r09PNzD
nrBHLTeNlZaAEIbfF7Vbyxa+OsV+inIC0WeSgFSPliPeMke3ljJOeMvpGqiG73U2
3xT6SpX56WMkHBgX9XPCtuDM/0DFFUETU91xbzpUarOrtd1mpii/7EJJVa52539J
MlZ6XcJkbNjxQoT/hDUnthcenFqNJF9krfQ6ghwdhl7rW5qDWYXYQO0xlxgPjXoK
hrvwDg1LuOblIVrdatzlh/pKDk4vHUiRQT/D7wf2PEAD6QsUWqxwbLF7KdUB9jPi
+tYAkPXxKxnsBAiJe28b8LZnw2QEFub4tosg4Q0ZCHcNtoWqoKRa4P9qiddhZ3Cg
qhiSDYoA9Y66m02rTvitAdr8JHxyxL4kKQJ5N6qj1rY9S8FchkwjAm4KnVHQt9u+
7JvU7csdBtztEOLHKKYXuTSDUUZ52+DZpxiOt5fS9DWnRLzfeFFr+/ieLoUu5Pfr
Uhr2gm19j/jkuhMvBg1/q0vBI/sYaiw96HL0kGYm4nHH6rHpOFCtcccTT/5i3qOT
p+1BVLV0nGzaccQKkL3mzoGcx//6tcHm/AQJR47z90vsEEE64kUGuDjwzc/TYjn/
e2vhjf1pE2OI2Q8LczVOYineTuWOcxQq1nRydFVl773/Rh5U2cAJZYZqvQdEIkSV
VVMTS1uwtlpGbueTbHy17kfJxYE8uao0CYu+1UZXxv+27BKYgddKyy2zUbdcrt7V
uZZMt7m1VioBHu5OnCo00oZ27i5ujQ3OhyXDLAcbfSH2Y2wnBmK4rZKQikm7YcAs
kGT2KNY+/y+q+hqXgjyUF/BviGWE5ARx59CA93/eQkuz43hjLbWfxXMFO8auJkET
0+mu+GmA6cj6A/DkS65kdpJsCHmSw6cKsNBSFjB/BHOpYsf5J8Aq/1GYq0mxagPm
K9SOdssYoHLRxPbHiFmh1K3W8rQxkxywx2jFkjdwngTavNSm/OdOhaf6eqdi8Pnu
81BNAaGDRFCtextQwVda7IZSuezHoydBz0ZuSJKj3BDj7GjpGWW43NtN+HwnqlrI
B+StuAzqDQ4QBTLlEx9+DZmiowAfiShC/Pz2Awiy96Vvu+/PW+mfzgY0Az4Ha+Ea
IqeyyE8kxcXIgurpm3juCG56hfizriEWm4E7pl2P42WBcCVJIowKMU4DUYppsT9d
fXD1DUGPCcnQ3XRUH+3Lqq/OZRIGz+ctGhCI3JjOlT8RsbeMjWYnCzKf7jPKOnFb
aJRRjIO0MpFvftOjGQqXwdmBZPk/GJtYjeHsmt9fD9YgFaYGGbOYt4Ils0QQh9VT
5v5gGZtF8QyQQmuftLLY3Ejjzsj6t30WVYeQ1fzlrBVaui0XxwL01HC+Q6DEZBAM
TDQnnHRBj8PrvbFu2gkc//B3vWeNQUnr6h4/GSN6FULIldU0b8YmY1Pg2yvbnC+9
Ob/dnjRoDBj+/s2K7+mBs355cN7+bVRlfu6hi2dqShw2cMQWSSnShnQIwkQC2fVp
GbrsB+G2eUiOU8IGEBxILbG+ONY2NtjktN0BwWHoL0HvPBK14xqgLmsILlUvSVKu
Y1Q9UpetvfVcqNOsK171ebk1EaPW+uAOZOZToAMaNyMSvIgrmMVYUxeA2zz46qAk
7IB1yi/p6sqCxh/bsEH8QgIhDsZ7u45KGyMQMAt45OXgRkScVqN8oSEh2Fl0waML
hnWx/AGRj1EykPsfvVuDPoCKD6UKAMaowqPN2YjnXxmfeoyjh5LIiqBt4sxs6tse
P8XGLICu3zR+IIrvEUpQJPvypxraBL1prrF/3Hqz4qhJ0L6PdurWUYs9fIi+Ji4z
xhMjHE5YOEZpKiDD3wjVTsYsFBCIqUJV6eYSNnO4dQUAt4Iz4RNlhuFtbhEdJgFO
joFmYhFLRqevWNr4Xvurp0icg4CITykIiwnpClLvJ+6arhJVCIIGXoJCVw3xYKpJ
jQVe+Jdk0Jcmgh+RDm/gmgoZ7kn17wjYeIPSXAV1yVpZvWzOYJw8yh9scluDqieN
Slk4i82b+t7MOkUIgc7TyntKmRNfYOeIMIvz9dt3GdBGvxIBiBaK2PoUbi3UFdcJ
v7j9DAGpWrzOzTK/jHdvzbYJOCaDoLE/KTdM5qZRUPT2wkCTkLXlN7U1mJd0gxt7
gsXS8tZCWGAQ2YTEwxML2Y5PG0dH8U3FA5eiRxEGPWVNK+lfeHBIfN9vMpiUfjZ6
X4lUuEMLCWz1s6sbF+N+bqD8QWsvABiSRzTO/GHmaNyfhmtauDQNOXUn+HqZ/Nlt
MJG+oQMyFhajyk7NKuo093Wn8faiBHU1p2gpsCo/qTdRsPFNcGwrXn1h4N/4pwXe
NTdZhzH9cv10rBCtii3GbDW5OTvoRYAxP7qdfmudh1yRluXUHLsZJJTMXvBqoZeh
dOLhapeKAbWQQjfpRiO6sXuptK5IXFbZuywTyIbJMYDuzAILDqqg1Ytg6yFbFOxh
atxEXMQWQ/X7Cz+hc+b70TJonmPC/0KXVA+eySVw5g7z14GV0rNhm2ezzNRpCSz8
6NEOKLEDdI0627IvVerayMWRy7p0ix+U8MstqsepxBUBfqAZhYSQYHxCLA8bqrWF
iK2XUEeFvt8FpwTCccL3yCNy0WMRk735+kdrfG9GPOheRLHhSuhi9/w1EJuMB55Z
V86nJPzgDCj+OVs3ptzAajRil7iNx28+7itBvLc+Y/Wh07Hzf65d9mmyHf84GilC
6e45WGHZHttouzF/CwcJazsgtppK+vOgbE6PO/o2xPJ9G2/6N2I8Bn//Dh1O5cqj
UOoa62HlTd2/M+SkUKbkzWsmHVGLPb1MBAI11hLZuOyAObNzKvANYUapTHmmF80C
a+jlMou4C9m3sWOKvKi1dAYJNVlJUCoP76lw7TsU6tlMASF82YCeNvuHrEjJzzk+
meJRAG/P/s3Oqa/IkFWK0Wl2ICrl2vyzs57JMrjVIKdfSKgkGpngcpW8sKq3K6gT
YwBDneaA7dgIr/BIeHgAUHu+R5RhqHzglWNppmvHOCjE5glIQHfrLrKmFAeNJqWf
lzBz5LYqlypnjf25hRiRXZ9t+QUwK847mLKiNwC3TaNI9SyerLH2BnXoH5+KFKr7
myGuIy4QJ3KMh7kXT6t1tG+2yClHadnEBaggCO3VzRngh1g1zlt05eA8kJPGccl4
W7RgEc4kHi1uu6QFabrwx0CRe6BsvsnpsuVZZ3DbBib+KPvyPG3F7sGC9Ob/nt9+
9EFyQvvlg5tDGpbEYIP7DtibZPvXOEq3Kq4Y7VzrZkfVxu5rVejJV1PzZG/Ls95K
yiyw3bwtAUqgUr5YnbJrnXDovC8bVzmIV1xyfuiSWdFKF0aBGROi61oHLKr3Q6GQ
pcqDMEAJNuDtQ7M7GYU8zmXAdnacfRCPKtiIw6QhYVPds/uY5J3mr1iF+0BjlKxB
22C8Ail3fQ7EOku2Up091HtcUqRkJtZHu2MwrL5nSKSKwd0JR+RR5Cm3mJ5c2/mY
DqtdCWnRta5fGMrYoE+8wKMYIslQklxSQo0F/iVGqOqqRqL2/rYbCTkexpmWRxX8
4nb1fzXFaRGQeiOGRXG8US10w7o7aenbkxH23158DWQCl9khr55RIPQQp6+0luxq
8ecHvQma7T+bfC6L3Kmtp7JjJCp7XhUknpmARzfGNpxX7zoHjZcEF9+jAGD3b9Rn
rlI3fZG/t5YinUcJiys5tfDl7WSuBAWTt+IWWxtORqXL2TEq/i/r3oYPEXnh5qFL
u3ZLj3u+0IbkIkBPp7CbxQ+Bav3jp6/m1y44Apt/j3ZL3QVbhqcmub9G6CY84rcE
rZoGPPBjZK9poD15guNbhMLl79m5IzPn5+V0frUYWcZOcL48wGEDLGG0jlTHyFNi
40Psp3b9YykdfCl1SZErfhEge5xk2tgEZmYDaXC7esSv0VW6YAYYPzml+PHlJaQN
BSDKRZQGG7tDGRBk347a+6TAjzNpRLYnTtS9JhL7CqIbiG5xGcPUM/vyWreEi3Qa
dQ/aKGAVQKpt/08xOIZ4uFv+HJVt2GpyDRdTdXHRLbbWbreQFRmu8+L8JGgsF03r
BqWh97uuARZmtfNLFj8VDioT16IToCoKQT1FwQxupVceopqGaz+yTPNmEyLX+1f1
1GtTieYfSCWfRkc6g19Z05JeJXo2LeDgnDtM9qd/TtA7IiSL2jPryEQZc3RgUpDb
CjQYamYxCiaOBxx2QbhrNSESpLyqVat6seDg4v/frTmY6zruxu6Dr/FneYbcsX+g
1WbOMDhR4k8mpDSdeCBMTqyKDzjsbBkBifz180DjRhDo9KDQUWpphz+mUlbGDqgZ
6LhOJbOn+VyTVh2o8sTd0n5/lZTo1yWOlDtBFH7VDNmhBSNYiSCikffHy29+rTyD
CojckVeRj+B06uG36mqCQ+x9N4YFUonf+ufR2+lZSZS9ItaohG6u7r7g9FHEWGeq
01Py0Ksmr0XBpcMpqHfC/nMrCbSJpd3nK6rEQFPAUii5o3/MgEVB1asQ05cGhpqI
V5swbeTefM4k59uwcAVE0ahYeLSpv4nRy03DmOBiL/N05OzRcioniruSMQwu5+WQ
47JOP6zm7nzG3d0P6q/+mpAph3j3fXXcBe1Q/CujrD4B2/P9fxR8woF25u3LdkFC
zAh+75xDjFUw9L+SpniNft98wS13eg/6eINrvRMlhq607fGUn746BrgoopUeproh
JhYEtyeluft/dam/PQNe15nbBHcBOFwYbJx07wwi73JQw7HCa8A1YS9/UAJP3YFV
4G8sxieq5kHwCDP14YMVHvqJD0YSDU1TOHxjDZNFY5Jebak355ceOMTdZ/vFGG9N
M+IIx0OqceiYGIIzF/tmQINJe1ExlVpJn+BKkUK52bSC3gQSzzCN6xy6U8GAAs+b
VufLQzeuGOu7OmEAIQDGLepvLVHAi2CWie2D4YZkQqXV66Z3Aqva3807zA+9PtOJ
H7kyBFq0vDLuQSn+6RWMIU5E5yXPNgVd1e+D+OS3zUT/7XkBP1lZVPjVgc3uyn5v
34rPcDtLWrxQdBpNRyx1GhzNAOndmHfA3glhc9fb/sLvErYDob7RoMpnOi3moVEU
O6yXDJraLqwzVq5rQCzbMuUW3Fu0tbq6E7NH3Yf94VR5cCnn4Hbq5NLx6Gdw4Kde
o2wJzHzIA0v0BulMjJvIeKlj/dWbyTIRqQp4w06uccCEURH/CvI0w5dDijv23Aek
kHApmLb7Jh4SLNkxWIdjUSG7g3XaLjaBWbjX10jrbIpA+kDPFo1meaS34qQo0RrI
tPg+DnnF70a/7b8osc3QD/9i2SFQEL4I1WQULOYcKgK9sQfIOZ2aAKsprhfYbrqY
ehbgdNwA0alUN9fy0sSssx9SNGOROZID6ttbDG3tvO4MGIAmdiwSroLcbRlBfBw0
N6LG3NSSE4shbNa96hvKh4fDLR6c4HLwNDWhK53zCvoLTTPddzDSvRKtR9LlidRj
FiBq8th9MYq4By6YAmhN6gnTQaASsKx7CeJLnVWZWLSRYxRRzlHyWjpQZvRa30ct
NWB6aXf+pu83nruYWPdwFKuvD53M5GAJE2aS8QGgUNF2fZCFS2nw9PPleJD0MyAQ
kSQtgEJGxQz/aJvUfYnzwsefZh6g9yVMnYoZ2f7rz/q0m5LXjTalVchezr7Aicj/
tm8QfQl8zMZ0cv0+ZNvDrEiHPa+Udafi1OHePeQVNCL175ez1/3ZCf7mq2xD6sOF
rZJn4R1RblsNhlWpoGOQiCgh5KbQSa3xhKdr/YUHkzlhliBRJUeNn4IUUJK0BF3r
UyhU0va2eHPr160vnL00gSTZu2bVGZI/nWgIZZP+KlXcMof88ru7r5IaydUxsvR3
tnUqRVOZQAawfzNfTOlbdp9dhNIy0SN1v3DJqlOAMsdU+FLanuPrPRUHzzVuigzD
hCPXIA3YzKbcjoafSEjilYpueFZwx9HLrS7Va3LtmxiNq2ZaHHCw02qbQRgOLx4Q
Qb+Gp6GhX5BMJqWgjVRqqPMC3Orn76JTsg+hM2zLsb28N+M1DqtSfUR3jFsBHHw+
zNiqKNBgZ8nhCAHfvML8B46gDGC/ic0q/upMW/5wbeuuQe8xjv9vJ2fWCYZ6Uhjl
flo3uQbtBOyLAbUR5pdLbNs+mURTrCh5dBj4QGhmDogbDnDX5xlNs1iWF1vV1pG0
rKnq0Vnigc0g6QIfty6LKSKUvIMsbLzCf/SfRo4mlatpcaBCg+2k68Pe9untE9ov
YxmCkZa/KGAyZOtPEhNjsQV7AklrNvj4MqWW7X3mqFZE00BK8O68Z/jK7JMZQq0V
ZjK1TgiZxPvOvnEgsW88EY1qCAkqU6tF0/014v/lDhSaotWa+Ev2I7o2tmK5I9l3
WaUJOVpXJlWymnVH96YpwgvfpgTmK3pJA9Xpc9ZeUWJbPcRVWTCluivb9ahTKiLt
3iMbfNcFDFpvMxM7wUypnIug+UO2gIAsCWTkL0Rzzoc7SvazdJwVbvnDtgOQKwhb
5m6+GC+ZCHkG+paiZfLQg6PSlSU4G/NPvh9cS0E8OWxBnXQ4gGPhxuOppsNC3dVq
Nru9sfGXutQXBfcyk2mNS09gBpTgUbhNCAvvsKXXo7YItCzCZVaiUBPlCGzJcJl0
d58A0JVyDTZu1NPtdFBTiHyeM+nv6f9QDJruMzShQ04GwwZoX3wKunwFKC8DQ5Z9
nm3zjgABYD36+7S8+22+LVZvY+KRDkKyTxgguuWOjYNK0T6h1dYG1eQkO90a1jCK
bb3M9Sjkpf89LurXv/eW2Pxba4XVOl74rO3PWYJ+yc1PN9kgncZVcEVnxm0n+wV4
1463rLuseen1BLPTJBn6yUjHj9c6vcMozHlT+UOF79a/Y2nYaxMDbUgVUvoPjyeT
e4G0w886tGF52gNH8ErCCv2vQC/UmSWDiKUeOY1Zf7QBjzelChzklHddlW35fNp7
kEOPFhED/jD/lg5PC3FVAtEVnG4nOGx9FY2oITTnlvks2NCAci9mwisrEAePKsK0
lwxMi7qIHn5VVBvIwOsDNxAyWTKv1pnGnktVukR4Ub0lsUT41SyrqaskQrO8J7TG
jX7UanLrJ1cxtGodHfBPRkZ1HjSOWzGbv6spUc6Kx3WX0BSEhtlEZYUmRWoASeQt
D3qGbMbIUKfFhvrhBsqxDft/SGzikkdYhgnNP3Mw0XLSLGanAWbEMSp7Fsr8SOJm
+9kq+u49vk36njPQAVnjzocwX1XEgvQL4eZ3IzLiGSIfcqghFxaITBBTtyvTZz6h
/ob/qGa/0XsCPLxY5LN6Zc5ZM61ui6lYVHlH4EkGH1un5H07J0vDx9UueEAsvgAJ
opxQDySmJvvCzQHDGP9SJoDUoOCDNWXA5gcce06d2qDd2rOcKmCH3rA2dGXrzHmJ
gGiJwMusNRUfXiCKtQJQxqTHchfhRNLhk3CGe1xfTgABguA2K24CxDSUBL8ysvYo
LoFTpEhmcK9HE0pdqbtfu3l4S4PPgU9WCutx/3CNVbsiKm2jIxqQMm71yQIF/dTu
OpMzhC6i+QphJS6UK4ohN5Bq5Pmg4cgFVNGPWmbRIPgAvitya0KDcYDEyEAH2fXn
ywxzB2WBK8Wkf53JmmenrA5LaPtshhuNAirTtmXcQ4FCr0VbZH9Q8IFMy1jYShrN
0OeccJtkXqTah0K0H33Dgkzgx6uuYyYCoUFINIlmckqGF1CQMmpFtpAH9zocIZID
8hvbugmDeUdYifuqdVZGWsYIj+T3VOwPoohl0XkTWDa7lilGgJQw7V/ycvcQRiTs
Qc8495jJcnzUcth5MhM5cBPwUsRJ3FA4e5k8gYZWTlQShVTGvU2X2VPX9mRwj0gV
aNnGMS4rUNhSKgleI5JcTtoJszpWkClM4LFPjCGRtYDgIoMOEThxdCuPQdF9fWJ9
r0hbLj6zngQpGfGjeocvFUadomZOC4hLjBhrKeJhk2he855SOA9FCOL4W93Lav1J
OpFOvRncOI2ccvxazBgMGoWhdGTHyqLll50PIjFqTz2l4xmpFgJVgfojZm0Wu5kf
kZIkPLVg0dLmcU+UPJU7gHCqterzeLHFvb4jSrPugKV6GKjxMe3XKgHqVyem4Wkx
j1PI/hZkJ39rXfO3iL2mqNRJiWMOOuGTn0SyLWikeXukeeQg0562Sij/MDgC1/A+
3zOAtS7EJnuads7lvH5+ZXLZdMI489cbPjiyWWcb23ASvb1+jhKPtr/NWBRANJe8
NYCDuvbJXMicf4yH4OKhDEh6j/M5PGyEdXOiJ4w3NalK3shXSKxmf7/gpRZdgQzU
2gBsiVXmSivuZWwfXP74VbSULCVNLUYkZrlG8n4lds6dGL/sljJomA4NjRz9zGZi
JGoHYfkKA6jedFvH4Ze7UCW2BQ5vGue0PsudE90h7nuEINlAta63DUYD9rxlvI2q
xGyOBppfvsSjPBkfRyeQQvvRF+KcJVXfDSfsIAggTJOFkk9fnLriVUHzGRmfoH1F
EWDl9xjShxy42puipyxQsmC+4XgJI0fJPlM2e9u02GZqXiRAvSH5WPOBtdf+VJVq
xFCnykOIaEmY5C709nmwd93bzADbSSDLSAxz13nS07INX7FYBi9+3IJ7ZU/pBO9p
FUuAI2sdKMuGy0C45oOQVHI5Y1vwbikun0dPI7kcVlc2ZwETICGOYkF4N7BQaxmI
7B1qWT3xmnV4EyHg0Z0zMD0vje0dN6mTPwnsRvS41NPVU1p5okRNmKccLazCQrri
0/V9Mb1+VgNTdU/lvyGgwvefw8bo2fnstZ4QPMw+NBIBa8CdABuUjtrsDDawL/8p
oIatrxTQBGqHAtePvjLElkqXZBOGhJu0gkaDBpaTthNyv/jIMoPPEAkQgJ98ZTgM
TwDztnqQ6FZSrKskB4kg944PZO8xPF+dr4uJ64xaV10dRO5Mt1JckgLdD+RenrLT
okadKsSeSkWKAtqnNpVj3Ot3zL7FMDQfOGULhzQPSnEmjTc1mp4yGJZaCK/sYhvc
Q7GZ9uelZCPJ/90rs9O3ErC8yrs2zse7vEKucnW/LLsHf4If+7y5hsAbewzR4OpA
k9x92A/ECG98uzgci2MdwN2jGN0DOxITupCXzev3QBxpTpWLMuQf0xZdEb+G9D/W
CG4dIhwc/4E/0PE6VDAG6PPHpuKp/wffHGMePHrdHgRLcucSUBk92pz+ZCqwDDdw
ZaeS7NWLLoYCe4M1x5MiviJPhKON8n0vpSMZ6AFkqg5a2ymxBHQ+0ZVDkBxw4iZe
OiqetLY4ipvEPIKwuJn6xrF7uTk9/YsgP5dIA1Pp4MRQSi3GMgWsc73REmztQs0E
kc4IHo0u3NJybkwGyZ80rKNblnqw1/xaI7eux3MxVp1na/gAQezY0rkJoug4SXuT
xGmyr3EPgV8DM5yyxb4/HjazfnsatjqYK2AxTTcwGOsNHGPXdBNPEe6fdpMXYKhD
vI9J2vH0MqlMN5oSeoYMEGlzi2JH6mnNg5yy+SVQummJes5gL7sVk7IoXWGAQKyI
AyeTnnUTNR9UJtJX5xSuXBvyfGXjWKxRMnRLpOEZdoaAOhF7YDdxT53i0p0d5GuX
iGV9P2sSTMpS+hlbL/Bd7ZXQsLby+aqIxfpS5e/5FezA9AOGRwcJ5fPHZ3wqmHbi
1c4VmUBw1QhnLaadeOH5aSfdAp+m+wrsO5QTukWxWTxeq/kgmmM1C1L/UOGMF5y+
G8Y5f6euHcztL7AhAp0YDwGxEpwS5u1JSJsMj9QZ4oa74oTbAW44T2eX/qOnquz0
Pqc483rIi8oYtEfmSJZ1ns31LeE0xAWQNkoMoqQQw2cQGFF32DGYMP5YrxG148hf
LRJ7Am7VO/r4bx3jZBEu7GTqjP0vGbB10k6LUim2qs+RS1laq5ZLw+X2WvCP4M5K
8xNXRbJND5xhkQ+33sSDNVc6j3qJ3U+bvMLfw/7GlFe8NcIF1PPvxaFyIfbwVFEp
3kXv30+/EKphiSHtWM9s1IabU5QB9LSydGr8kVS2P85tt5N2J8AIp5yWajf6Gp5q
MzADoe8wFcqiTYyz0Xz27/xCdrWtqQo3Y8yebcdxSKrmxaFDSvkypuDd/4qKjwsC
zKF/Py2KtmVWQSv9JgUcvXjTUNrD2l0nYUpCttzgLMaDEpRb3yOVknwqA+SURGEH
kw4Lbeu7h09uyhyWyadL/tf4w1txsQULpqhyoASAnLKZRKxv5IPukNKWMhF3U/q9
MWdkyoj1RtXHJA3YRqL1QhDzgZf4GJ4R/4tkTnQky2lLGocLioUISeuHVav9A3PY
By2ICuJzpzQo9C4z+dM03bfAoAjz5RDlFie6k3uknl0CAs4PEg5duzSUSjxctrEP
HJzHjCznKhtjui5evI3TYA+xBHydaVdBBD7ZaTKdd43Oj3/Usrri+AcTIAIY0skV
bXGtDGHXtUJ/ESNuhNO7BCBGKy6IneRhN/8c8n8Om93NoQt5JY3W6peeiZKTBUAV
D/snxweTd4cwdm2svP5+RnLX1rMD4tuzzF15ja3+QGdt/0GDxixHRq7ORhVuArcX
r8d8EH1fOEI2NOK9gJ31XOPNaf9P/u+D951X9DYu2ErbhIZW+4OmPZL+arzcogfL
M9Tdg10Ie7l91Sclgmc3hxTfBEuNnY9XSTM9773WceKwYFA734kiBkItAZuRn9Sl
Oopsf0yz7HXhnOJ45jsrQ4yh2cOLUghXIWM40V4DXHBbkYMKD7tdD3PTDbPeTcw3
6ALM1qXfDlmfeFxiarADsebDqZdpVz43ZeNnfUVZunmz0lMcKZdofmjysuwSSJuk
QrdP0MCr9J/J3N8Rz9SndRO8BHTau/Mr4yNCJjVHnyG8+Q97FUqBqL8TQF21i+C/
wrJ7rhs+1+CI+/yeHSe5hVtKB6nMWTVwKmGR/Ia5LTptjtI8WrRu+ScQjK2UebGO
CwiTL4vC7Ua9eIkUuvk0v6fqwaJ+jGAlCHXqCeCQ2uv6UpO2nKAoi8tk2cb93TE3
mOz7mo48exYlpf9HUIsWe/KvUvJGqKc2LvlO19ixCeSziIfeaoQoeGBj2Jlj/9qI
1yhJ4wnky9/8tdcDKAdG6mfchDpMuon5dy9EeKqcH/Pfjvz0D9FjFnWwrZXXEpec
giHyZi57hxiwgYUezq8T4yH+Bj3O6CxboVWBntXv0rWRL5xauhvCbcRTxS/Ugv2d
UbN6ndhSm3HvohvWS4rs7ZQ43zYvglleXsTvQu0X7fR2vvrHsgn20GQc3QZ8GB9/
5d9Wlg8dNR85xFnOSkdm38ctR8NncPC20kNw3YIcEcukAqSZU/wXlE6uJcyhOSVX
fDo7Jx6and69rq8DXHVDD8alS9VD9aGSgP8fXrH3q1oSBg6Oz6EQbePtbiGlcdAu
jDpkEoLVYZc/wO3VW1omPdofk3J1XgJYsLSvpuZWYXkhGfol3lgfGLFvXK8Pm3iD
2s43OjuyvcyUVcSxTd6ftTQ+hgteI5Bz6cTvZabkOLeVvYrALK2JYaJJf/otmcl5
HF4+WFxR5YsJ2mZeXTdVU02dSgjmbzEZI3LiSqHt80Ci5al7f46Pc5LC4BLXK30s
4J3Qi6+YVCIVHXt5S0kLE63jc0t0Va2OSn12JULTVxVJ/b4azuDxD2pGAtQMIj8t
LImBZg5G8fg7pG4IpExJSHHpLLWpacb3pqy9vLRbxXWcuVo4PHnf6vr+kruAQbZD
f7Pq1Id3TsFeFSnFcGg4LB+RRjoD6ah1i0uD6To0BXYdiCYlMRhDi59elYNDi/GR
4Caq+vtQKdM1J1Aj7ToFBkic0i4Uaa4cWBp8IByet776m46ENgFUAO1mNWs/NyCb
j7TMiEgtOPYydcZGF1QFeZkvT0UgMC6mvBvvaELbqeUwKIVrz8zzGrUYlG/k1is0
x6xt/S2wIwD5XFHhwulmNlQdWWgnXyxGKRdYm2vmXxSnUWTDkzzVGv0BdeQxFMLo
VAEUkQ0r6p4wadPh+xeLlWIH2hsjUZFQi8Sl3iFUXkt8+09Lie1Cc2nSBvyM3hu3
PuDpTDw98CHqSr6850+Tuot2kW3Xj21T9Jya0pQDBc8YlV/gwYuePEEDcnb/61YO
inHOPtb6jGv2bAjMH8ZBoR0n1XgNw4azhNAcQPcjCJfDwSMxSi8fa3FMSMJGSI46
pUKkrVYlo9y1E4fKzGXujw9FGf1OF3EK2AXooIc0QJ4UVnLxDJhhPBOJlojE3YU0
aZqAymtk5Sba0BzlQj4/d1IXJXsOMN7gHV8dJB9hNWI0R4BTY/36pdPDaTT9/IYS
kBe4BpTY406VJ6vZdBhdnSM/1/ziwMYyb+QYkRAc5jTjvNFJZxRWuUkRfDK70jsJ
yPNNmNYkKrVUSQONTH4CVtYBYhVyND36Pzmg1r9puvyyu7Kt1s9j1zJEvquv7rcQ
wK5SwZuJaMrSnf8FEsRra7UlY1nSZDf5Ai3AeaTzf+SqPCebqbqHuFqdOQella69
PTekUcVGOt5A5QVujd97ahuwi4FxpjCo1xpxWISZdrjSUWq9XGoJwpg81WPC72pa
Sn/q6fJAIOJ+nt4STB8Y0WKvvDX3cUYQQVyctCccDAgpujSgzfjdKSeJWTxPJBtj
SnF7p+bgPvTZPgdKLhS0zyd73q4QOr0EXsidq22Px4+pTcsK8L0dhv2szScY1WqV
VIUXXAzm5CJs9qfXbPoCDF7HWNXRZfRu9e8cPn5zbrhth0qSUAuAI2jScC7bphdc
A1gVCVpb3KFZbfVsEmEMfsljQUIntM2Zm/A0JIKt2AchWGoFZ6FRS29uTmF47IKU
3ddI1HRYCECe3RhSneN+biZ9LqNbP5ES8eWc59idTMt9WNrPYZ4oEyemivteGnzL
grg+zKlsAU7XtxISOlDKxnQcFxhKpX5XHzKbQ/t0FRJKK01Rd871ImIsMlQg9a24
adODGyLAlhU8iWlsNkagUYyTgnYK/vjPunyxjxAHLd5FHDyyYz9A/cqJ9xMaqSVd
s00Qu/NUZ8tKQO5nqyn2HCKyUxDolwNgSY4A3/Dmv5rmhz/j4qGH71Nwkv50I3Hc
sqUNg/cVea6aVH+jxsrAXkwvj3EGSuPBQo4Aztqjo/iyZd+p+m/NyZ00sB+jx2GJ
T7IqupM+9iB7zEKxLX2NVqUnJqQsfBSR6LbD4O5a2RDN6skn8FpryxQmzJXEBvUC
GB29Y1WJiwnI2/kJDmPTqoPXDrSh5aJXPfznR/xBNrAi2flWCHHGVxjGvAnnKUyK
ACAqB4qYi4pC3IOlzM/4VNtez2YDSnIfhsDsu00Kkc0a0qv+of2opBiaKROJa0Mg
W9iweNzoBb6ibGBsEWUR9Nm82OIrZj3LXRxaOZq8X94t6bWP1z2RYYNf3V2nPyco
tKHVU5/19Ncl1GndOim4wULoKuSI53AbMvKacE8bF2DdLAjcq9pP3RvezsV7A37W
jAbfz2oyXGGzhzH977vojXbPfDr1Z0Z0FgTOKEdWP0I9cjniiouN1FkOU92wS4ne
thKgIl4e2gZx+6D3509uEecx6sPUATO6N4xBvw3abRBTEu/AIXIE+ecD6CEDyrI/
6ltveJQmSvfMoCW/u3zRcpz5s6ZybvbjeyrEfLyO+EnYkklV6+cbwTq+uD/5IhWV
AaV6/YOs8KIWQ3bJ9b+dx6O/1kVA1EBltvVf2BCLKPsKSAxTtW4oys/QjK0+a8TW
yEJUb/W3JZQx/uhheMxC2R/BYgxKQ8xHwB33xOTRWr8vh41xIRxYvBqL0UnfRBYC
Z2oGmQiRcwtOm3gllyLYsyZqd59b+S3Jldl+kJ9xADIZIxk1WASHSltQUa9My/N2
GcNjQFntcH21GlrdZFEgZdj4qn7ir8wlUC8xVaMEkj8W1hnlNXELmztUC5LPGU2O
j5wYOep5IbtaUS38eLozITd1ngYfA2qGu69LWZOOaIxZeRuERQ9F+kpYMke3fJjh
smeyaICsXp9lNv04jINpzYcMkZtmj4yw9IWsZGDy4j14iEjU7VbZyBknPLZHUlTP
Gbr4brGcQ8ucKDIwnDCmQkioU153g8Br9gKehi7WddpWh2Aovw2om397sQ7UW09A
JFE6PAkFqdEPOxAY8F75ss5brefLJiRFmRIIWNVgrVuOy4iQGbrC7rCBB79hXkxM
bIyCZaMRbRTUjlIWU6PMFVR0pxTXb24UrwD49FillqMrQzKtctfSi0w8ZpYAvgTV
ySbPjlbxdkzF+tALygTV4Ocjz3ucC31fuWMsWHID5/ckWC3fqBHwKGpj+U74FP9d
EIAv6yB3lprmpJMZuEn8dm3HklXnUFVMb4ttSZ2SoBR9yUNcsdDvj8i6Ui/qUnXi
APfXRmlExY/doZVuiP6K+fDl863f6mXbjk3BKf8SWErdqVeZkhmn4fVz/smiqQes
XkSaVJ9pYh6DxXdrYR9w+eHCmWUw9ION+7oaldx0JqZZd2kpGpdEAJtt4wSSj6Wa
EAKIb1EcIl22xbIAg86ZGUW1jcFBgZSclFNC2XPhdg1WO3LPNMbx/lGCNNNkQSms
Gtt8NLH6FzCg/JSFKfW+il/tDXU+hRw48HaZkEzwelxT6ObuloJ6zr7idHm/8Vwp
kj2zZ7a41WSQyzGPm84vjQ9Ot9ecdmm9x92R0F1qtharvxTrulmMELkC8XLDWIr3
4+20O33m3bGOBxzxt3hS9vzxcIPo756IzJzBejJ4hp8ihZ96XwXaDSxv8TL3tuqC
V6d9ssJC1MK82hchmZzWTUQpvHMvq/btffPt42ybB+rwwLF0gINXHiTQ+T41A9iL
6B5jOvcdpOB4VKQ6wjTWjBetnuTZGPqw6O0uq1NfjqGCXlUwfWtqtQNbziwaxAz2
6ZyzP5/WYZIL035svEGThqCN/+TBr9jehHjdRjaIrT9P9IzG5aY1avuTU616BWuX
xPb6VK/rfg7bvGq4O26EUYk/6T8WJZlYUgRKZLQ51TchOG+83qdcKSp96v5MGDLW
FajuwTUxIhCjmib/qLiwta8NVaoyQmpjIpKxLs+wBHqQuvPo1v0FNrZq8zR4kW3b
I5Mo9PnmNbJHNO/o+kfsUe8vqbngphSTI2Qtsyh6RBO1Xci4bERnYMKduP9rhpP6
cxQhZpCcOKdSOibwzVazU0EZB8ayX0gD8WpXTtDI+zXQow1rekLi5C4yr5clCMuy
H2UoFLrKjtPfk/Z6zxc9e7ajEhOKZJrTc7MjiwDHnxaqG5GfqdjA+jvEFHXgCof+
iLRFUbY+fHBj4tLVN35r+kV+c8ZORVEOkG1XuAl1degkj5bTDp7PpZLKzQq3aAKK
C2PVoeFJ406s0YvKlWkxyVKg2Ghp9E1MzcvolbayvDpDV/qHiI9b3BCJjy/zGPZt
IWg+HvLdqTnBm8ATS5lA9zCPvfr4a2XcvjWSYjMIdL2PL+0LVUsVLEGL+C9cu0S9
2ixo+0YJrJEwKJJjr4ocZ+OR3Zc1sdQfiV+Fq5HCG7B+J5c+80rzVnoiupxAOhAY
JhBR8UKiTb0ZFx/yZrLztGYFTXJYejg6VepRM8ahs7vLj0Ji6RTGl+9n5iNobdqY
AgVTnq//Ed+r+3EMF8rzJxvCt59Sxy9LlwdmIbFu/JVDqpSA6vAd1tHFFuWlL5xY
JCVQ32PKKCDq5LRkmnZ/zq966nFEFNcRl4jOqyIf41QnQtpMxT0RLWnv5wvK9DEt
3AGd5kNXNw62BWZKDekhgBVYf9ajxezjPwjOzHl/Tr7NZ5DzF9TpKEW+VFxRyxJw
aS602DcsoZBbPhhfitH2ORQ/poQg0IgnYDYuZbkddOQ6xNTY6XHHsyYH3EeiaD6B
HKPw1TWI5iwr14rNBoR6s8qoopFiE3KbJU4a4VjTs56dnd25jH9TuHQ081+PntGh
CTjWpoPjzF/iD4+lIrMQcSx8CMYECghGpISsV4MkE5hdGgakJgSlmYH9ejUPxs+J
2B08FKvHcxo+BKuiE/yDsNzF+n3zrpDt9dTsi16UVFWq4HtDMn3inc5HswNgKYsK
ssK33fmKF7XaqQ5neaqRSHrY6YaVaP43+uOrQqYx65Q0zkqrg0ro6/tNUYwpL15S
Jwx0S1Awew4R86PFRv3v3BQ5uBoKxBRvYsnvWqaFtSUi8cIBFares2D+jvYGNIau
+VcpGoW89PP2BL4/CGnF4jhDGsWyy61AZ7if8xdWMZxeAH9JJw2sjnynszzUjAoU
Ji8ZpWw7BdfiLaNmXSXGhPyI4TxJ0929ngLcPx/JCt4wsL9SLMIvE/Ki45EEqtg/
2b9EEc8v7sRnMRxqKY0QlTWDorSAl6VwyamR6HP6A3PVkS1kMMvkVQ2BKRCzkQuh
k6eRaS+GIIox1YMjb6nJy3TD6kwesMfQfTxdLp7i052cuZsgYFF/SznsWATE0xqe
d2jo1ApIlWk2sPMs4YfNQHE6N58gHUD/zz4uxBeTNYnCawqCH6RpAS41gzVCuDLI
QRpz+ZmAc/xHdoB7YYaNeEj+2e/KKV7ovEwFQMNVklc+qCt9p0ID1uf+P72xGFaX
u8g6+n8wPVRSG5ajouB8mHkQ46dlThxGUxX4pyi7aceXT6ls3lePUY3oF/jUlVdU
xEDaI9+Ui7vTukpinCO8th9WnG5LhUWXH8d2j+oqBV17LEzvwPr3vGA7H6Jz4z8a
uxXFd54kugpYdlJYHl6n4JMjiGTRThWiYsFS9ja+XHDrIa+GJaDVppaUU1P/qagB
6d7LDmuOn7vBjkOFh14hfFrvpVFMTQ+sm7tpW9XJMsBlp0pwvk93yn+5wdSiShqf
GkUTCH/iteTxGb8lo3mm43Thbu1zzSpEUs8nybrensLZya8hAjPlMzkEn51tLDCq
3fVOibTnFrVSqfOGDkT50snFhenAgbFuhizJHMbS7vKt5CiGLc+2fuACjGjnTfqo
GbleKjbqkxQnqVtotwj3ajRcjuN/Lrf83SEOLdnGiIvtvvZ4yxgtBeLunuNk3sBq
DJZn6PlJtoh0k83roSG3toGCZWNCCSeobFxBBJ/BV3Tw2SADdwqe9zxxTSyHbHDt
ZGXQWi0rFdZvAowdEVI25TtOqXyITkqb+/f/Iap90HzXD237Oe3JMbDj7GulAEd4
5s5sVvyMlifOX/hjiDkbA8ozF01RFxzD+bIDki9kjoRzOkypVFiGWykOuvP+R9JM
G8AT7c8iLWf0YwaF509JGuCxX0WTp9Qb4yGeMP8YI+ct8NeFajYKvZ/GF1oy+20a
d1yZxiZnEsmihTPUX2FWyBsS9tpg4znYn3oQjGNxcJ2YWQw1B2KeMEGwv/k3CcTX
U2qlVAmesGDDuT7zyYFF886DcjIMC5nr6OUHQXqAM73nZI/mAcHe+0em8NAwIP5d
jIpRH6LW3i03K1fsqcaTtdamrLNAraX9nc4C6WMKZLVfFnZK7mOHQQvamUHurE1U
SDCAOYszFhVfDFHmt0Inru9wP+Ptk0dI6ad/cvUKlyTBT4NBns5f2Dlef+J9/oRg
FcAQkKeyLNVjm7cSAO+jm1ulNuayu8W/dPLrwqBnyBEHSg0hYpweV0yPoKeNvd5J
wZJruOg7UZk9TFe9j8XDGr9Mi9U49zjLY9GlST/ZgpuIL6eOqO/dgz9fAzxf3qps
msaTMaiOgNjVWRdHYG5a5UVHG6sANEUufgGDx4sXKKJEp4J0JEnpXFagxSguew56
BI69CIi9l2G8Qx9OhzcWFQ2se5S3unNSmI8UAvxa9IAqbCpkYB93LS44T8VWKOhq
H3+i/JHl3lR1CyhbUGnL5KIC/2FDRW2nOZlxdlpmWkA091oH2SYa8t4/BlXPi7AP
1s87n7+dk5AFcwpO1MVne8yY1z340c48L6MvVxNhyZtQOet6yUqk4PgQFgPHQAIJ
+n1EJ8XFSRYu0CjpxPXRzpKnnPXGHfMbhG/rHvSdtv+rvYMh+8gsElMZoaQ18zoe
0YryijExoSySVB6anYqVnVEBk86sCZi6y2ZgseDlYdup+TUFoKZtRdhvwN15v9mH
inMPFgReuIAHXk33JIirn3bj9peBdA8eOW7Oo6jDv0eCsAbNUENR9BeXPDqlV0pG
tqhTQmSvoXP2pHhWUEPzGx43tIeAccR7PYrtsRbyVfjbsehGsTxGnSi/BcIYROM5
QJCNExVH5wN2q8WV9TqTEgF7oM3S8dHh/8Ao/MkoC6sR4QZoBTlIYL8qqYkGCs27
tanzi2uRtUU556CNIb4wIrDeK8t2dTJ52dMabdpFNWpVblpniBiRlGLKJzUCiXjE
rzyu7GeObxGa+OmG7D2q/C5gEG33WU7RqQQzbS2LAxNF/iIxDr4kFkMQjnFrOOYk
a1UG/Scrb2Gx+vz3Cqh1dhkYYUTNhITEXn2nQHIAjN1DOdGlw2Rd6ynGNd+Hbqjm
tTECFiW4ip+hCNA3lB8amMk5c91hNYzhq4BkK+M8mSF/63m8Md/OgOojbhV1Ldwn
EGysmisdiJg9/smkXHoeRfBLf5YGrsw7/yHwXjTy+i9m/dp2/X3SfU6/KEV6ySi2
pikyrPrTPSGPu/8xSnXYvJAjCWRC8vMMy15BDZVurmV/5ujyzVQTnb/qZUDvLG4z
P9tUAjzfizWiik/btAv/0DMAjuHz9f5Aq6xNS/7v5TAs0DvbG0Nsd5wkcxnNfDTu
Dh14MtNr8rBWlhPT+2whdcbF25bYGz2PoYt25On7V30eFe/hb3ni2U/EdxhDSpXt
lTVliyPdG7YcpGB2cXTr4IhM+omYD33KIXyJKsNoIpnPotKKclU5HIusAkw2DN87
fVIZQg47eBW8hOqLTMM4cM3Y8Df0Q/tpdMqpDyUHivudSH5yIl6tlI8dGaXD2nKL
50hnc/CBqCrXPGBmu5tABmbNLiYaswmEJiybJoGi+7DKlRhg9Pvix0Z80i3ilMFu
XCViJ9Ez4ewDySArN6DbDVfMe7IEf8durSigiWt3Lkosr3N2YpWrM0k2j49k31vF
spRK7e9UYccjRSBmAAJb169NmTf9/dg/WvTvQjvLOtirQIuVI/QgY1Z5obc86yzv
D330bbIAaak+xpfRCSAisepj24KkgQKRK3LE5txz+u5KgHL3qN4yWqsUL1SkNiWy
iNs/OY1c2BhAKlMmXCrO8glOI2KEQnFmbgAKKQPeWsuRnLlaPBamiBP0MS5On5x3
rM9hCKiR1IdcN9pjZXc+P16c4tpCUsgd5bgonMIF41RQKDDp2dKO50VuJ7OFo+vT
YNVTCkvYKWNhg/T9/Uf87gqkuYsXOQ4XUxWliD3iq2T5vf8N6VeOzmvs9bhELRLe
RLXK25ifi1+JY57rTeKr5zMBwoUjkSVDnUYo9zb+X3ndwfhGgm5LIbTTYIketzLN
YUul7Yx5Mx3WgwruWKi/9gT3wDJ3q1A2MJBzRVLDCA5AOBpNwDFVQiN8dgZ4V658
KE7IaZQHqKzHZlUCdWrhcay0xW+8oBp5O0H++w/4Fk1D3rNrW34JUknNUBQtu5VE
iw//kPR1zPpTIf3dxYKV7dIvrozu1+DVWRmkIXVynivMSjtFCV0qpmanfumRIS+q
NvPhCK+9+/DnvqGyzLSzP0bxf0a4L2xV9i1LVbyJjR0fGN0tzBkaTI359RwMfE/v
4uhhP2pF2/0t2S/FTJ5vzKoUI/DrxrBshSiDmv15NKnps+SvsKdFKrJS+aYHuOeP
5S41FQ8iu1LP953w0ZWj5L1+ryG5e2ISIvmI/P7R++e3ODzZHIwIGIvVcp0QUCd2
v0pTATLV0leQwtWg7w2b0CbZO1T+31ojTryYprZ9+b1kuptREzFz+Ojeuwi37K5A
KtO0oBOEdARyoJ3TkLJ0BQAH/t/fFOkyizsSzBfhE6gDB73gDHjN9e/l+84ZbkPo
2XxiCvO4Mx2hFG8fXeiUW3sh1VdUXEK80hcWqWcQBlMfPzUjCnwSRd/fobkos09j
ksstcDN7IYXz6sCCm/j+qVhWf9ckTNJ2OZH5oT7IvdAHG7yjmW1iMoI6Z6Nfvv6O
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
O17dZn80apQ0cNYfTxSUeuOoAEzwsR2QodTsWBKlodm8p6SapxXBZXtFrU7HxHs1
CCXBfCCqmtcqgJUvWlJaR+51eABzIOvl30sVUiD6LZYUcWsJPkaHssMpSwfAkGXa
vhRAUEQQu0UtTaG99ttMrdGrZ1yswzs3GRGmYvD/F6OtuqR09L6yC/eFsrL/7O8h
MkyJg4qg7FWeYIZQxV3d9ydCGQioPBDS47hP8e+oSsWYwHJTcIWYvD28DtrAP6ef
WlxJSlSyrSs00kqUmoAsAVwANdDyrdbAue2uN4ZhmQTbEzMyyPtyy0Ni8EU60S1g
MZLnMPlYnYRkrKf6EJ+S+g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 784 )
`pragma protect data_block
bhR/JbuLrPAYKuwbSNoJPUFzek52HVb/fyfcOB2S/6kcjIAjK82tkZiT2xlTgOfB
HkKeN0ZC18i/U2yhGK5jBK7XEGXilO0zqmjt+kVcWuJA3f+BN/ZAj8jIIZwTq1XV
uACLa0g3JjEW0qPQkL3eD2BcuuqC4LC9I3rwRnwhnFj4UpLE1dLqACRaACE/S5pc
C0X1SfwRaCcn/u+9DSX2zH1j41Gha1mY4gOC//9sA+6QNKqkQoBC7wfQEQfce/F4
wGHFG9YQUaaFrgiXYG7SEriweI5vbfGz9Nrvj+MMj2FNllg+MXdaMczbLIhWV7F/
UQAPqH2s7JXNAVQto+PgS4D6tbGXHa5frfTXQjQI0IQmBsGzpmcCBqNtoG2jqXtq
3hUBgtEIbcYobYpB4pAYyUg3mXbGjerejhIY8BCoLVfZR3T1if9kla02kWOJBQ06
Um+efjyHleDdDZ33bbvQRkWEmob1ltAG7N55vBtcuc103ojcQ45JxyJxZei0KSeT
NW+h3Jx3KwfvrT9ZIGMjJkzuF4AyFoTspcRIiOygDoI5JueWDEUiCH1LMgj725Ug
+VOhbjrG0bWXoDufCp8IuNIU924j67Zhj4xYcpGWsu5makj6XF6zz37kmboe9dXT
XKn5aajXmb9VCZYTgQN8fxgIenrTaK24fFwyOg21sqJjpkZ9qK1sbpYOphYEztKH
uahMGNcKbULhpb7p1ghPg+G4hR4xDQdeNbgNRvIFJ8W2j6ORAncKkS632LYvjf3w
JaVa3275tSrFOqbWHmEFEIRX+0Nw//lgMgAAxUcas5VKPISKh8NGDdOyyzudwl7X
bzR6zIBQLCkNEI6GZ+nD9ifKvwZnCkB+44xHD52cJaT+ubUNLUYqTphoj7Mf+NVO
FPnfpImN+9pFmIrI1i3uYshG03awALiVGQTQqMY8TwxIDhUayaPo3f1BGfPRfOJY
OZPvqynnJDgbLA1N6E75JmYC43/iW0XIkBbOlxOshRcORM3ELnY8BeTvW7O7RYBa
evTQBJdwVxyTIVMJAvOGew==
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
aOHw1BsseDz32K1DP1JrIEIJy90ykQ17UA72WhiipJLQ2XjhQhRqv653vzKn27Kr
agdB0oJGVeMoUAT82RN4H5RmimJgSzVWhCrq0raix3I5TzQoPvFwg9c9kGc82P7C
bn54U95A0leXPiKbiGTrV1xiW47bDs94EYPyP3MhIxDes5VcFZPzqOf5CqCo2otx
rH4MkJWhvtBq+jwX38JYCFc+MganxNyiOFBwOf0kdXntDxBCLVOdRUj6IgRiV0mH
gvEi2FxSPaCuZM6oNGm8EcdbNexi/aAH2tMT/yNqQro3Gts1vhRTH8PvtUi5ABbY
9Yj8fJ9zRtU6qdMSPfnHxQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7536 )
`pragma protect data_block
eYpOZyNFMBCmqbPAH21vavzlcMJDFo0DecaOn4AqEF1MnUwLehkvd3p+hmlqsY2D
iyBuQDqiyEdGQ0TMllXSlny+M/8150m70CT5YfUfjYk+h5Ki8hf3bk8re5Du97tx
jw203cfl0WcylfCT/LByMsX8aul3hdrTW/P0iC0QbEmK6eMGPlOQwXHJIXd9qqUa
OlVU2dzhIj3wcCEQONe3Mnq7bBAebAwvQfFDOD3nomNXurmHy7XfCwYqu0CzrRcc
QaRvYP8ksudzRosukux0OP33SyP4awgfy3U/ZBwsx4Ne1lkmiGb31BhcwJLgm1aj
WIMU9kjWt7dZ/kCPvZyx5NKbHZO2dnHLwG1i3hsiXutzpQArFPYS9e3rRgYi1BSv
Y1SOKqgT3ovhvNRY4bBLAAJouAKk/VFE4s7NVcudvq/bCV8caI/dMbvDf46D2uLz
6qeH+klArpnImrAalRPo1T3kj2iW3miPFUZ0LzHorkKZ0mj8eBjQB3HmuGu9DkhJ
K+NXcAjLA8MDBqdjUMqROGCzQaRg4tb+TQphF4WixDKvvkgLl8ptimZ4SABk5Njr
3skFOkGD+H086ktIOQ12g/6LdMY2EvArNbSLBP02FnvnE+Z+UmemN2NNfMw6V7ZX
bWdjFP1QZmf+4J2Hr5JpbmVWYahwzgfeZix3fnju1VL9exoqkgMcRKGdr9JoxciE
YzmxCBtifW65/Kq6NcpscvGV48hgCsbRKI+uplVF5crzJTDcp+ihWdwh8ct7T15c
AppIyCO/v9nLssNjFZLBL44BY37UXrRV/xNlYOwowxhLdpJfPUubdvKodK/oeJul
WiLDxJ0eBcupu086xfVIQasqzs/3/dLtDAUjjYEArW6ibQIGsrH0W+4dC1mnoDmo
s+9L9EHFgpkuNYETyMu7sbo3/w0+gI46jGILHDt10VTvuzO4pVwbh9VrhTtvd90K
G5NOtsEvvDFCqupGj/vyjyNXtwkbWMnKOtCY9IUfgjgBRu1DL/frIoQst5pppnDC
a8Yl4jM0IpvZjKyslA4nlhPzCcRXUW5iuddcmVBcVQoeoAlu3wOCim37nElkl+Mu
OILByG4W9W8r+kEwBN9F0Kx4zJU+6ntELQTm8AgA1txANrNkS1wRt4lSb3HwBj9q
QITmiRDcF+OeGRszl06Jp0bkFL3HFxrqzJU1yqBvdWYPFaZX+6D3pvgm06vdp/1s
9UklPjkfVz7s5xLjT8WQ4tBmZaPTOLSfWopoq5EUd9Wf3xUzmU2WgKnNOfbQnZNq
pjkvVP+M8qxlIC/mKnYFR8CxmNQ2swIddg1UzpaiVWse5gHfH00G9T/UIqN4BQBP
E6JxQydD3o7YaTuO6LlWHgEeVKXnUStC1OKH2jeVKRBzE+S0LLINlkTdh3sZ5++9
w5OqkA+PcXYO4UO/10mBL7YicEsWx325oEKvDQFgVun7pmyOrOHIH6jEaE6ozJbW
TLEcq1y5H1KYW+hMmWVO7gMpwirIzKwv1DK6xhcTCuUiiwEpUr3x7F9XCE7BN19L
EC2AV2OEqDTpYdEMrECsiO33OrjifsrtOpsnjUkqGvSjlm1BcsPvqy6NNW2idvp3
vqHZfmTvgH+h+4xGbcbXObrY9lNeaLZeJZW+Df6Mc5PrkFVg1W5YefiQ9SMlUpSr
WjrGn/uzRZ57LnZE3oVqjUDGQKovvUrlpb6jj9zKek4dpXbCxzLfsrEcC+yVGEML
hrLEO5hcaimrN78Za44YpZWcRsUFRNzjAx4KGewXIeH+gm9Gh8ojSFiQ9o7M/I+P
xoYXIyGPnWRYxJvCaubNgsbjLDd++q4oaU9R0bY6aPheTvd/fMupvjCUc8Dpz+Ae
oXMfu2ajwCN7blnWVElD9P6lgG13iXzU3+/nHiofv66Hk1sm06Vx9BWC4Q7yUOSg
cPzoTC4W++Z9aThs6JdcWDpsPanSr6Y/AHCIFLYbXu5lvOfH8vGwwWNF21/M6z9w
SaauF/I/SrE7KsKGD/l6SiO4LUJnOFfiou7OhKdm5E+aeWdG2qgHm/D/bXG9gPWe
ri2lKulbGOlcyg+MYzb8JQfaWy4ZAf7y+WEa/aPF5k1fUxIzJXhjNNENdMqNPPMt
9GQ/9IH7AKAYZldonu+YI5g0o07zJo0IdZ7g0YcKMIUUX70GbpcvoRzPA71IhS6/
/PnDXDyQq/XQCjfdrobwmcaRwGbJGbqekzSWU45y35zN8dBPAHLianW1FJ/UBymX
tGSxmTZbEbzuB/az7SZxH+uUn2Ehv/q3jnVKtTAaPLRi/3qXBeYCXe9dtvxoiR/o
2/Yk7HbufjWLlYmsUomJyIi+28o4COGWwD1jcjAIl10f3UagfGGSf0oFe3LT9Qmo
EVo9gh7gyyguCkJGYoqESoiQ8CrFEaLbkBf1xeCojJNgz8ev2u/+DFbExcrVvYOb
1ScY5dmbOZRw+f6/x1wip1cZRYOa8vaYFFYwunQRyxCujhdtmTZdJL4qfJ9NZA2F
+hAiMpO9LT7P0gLy325v4d0UPP/HtoSbHMgcPfbEOgdSy8cDYSYTUpcNM8FCKo6b
le88x+VzN98AZ8I0Px93ZZmcOe7KbVBj9v6IEecwGLRBZe659kheKxoR6bMGDQ8A
9PAhvC5oy40T5NnnRbWJPKaIvMby6DoHCYDUvNZLgfI1qAbT/a+5GeHxmn+IodUo
D1S6I914++TyLOyV5dt5ho+/QAv+GfE3J8l2cO/c5We7WbFGerAHVKWes6bC9CEI
iKxZ/VXQkqD9sWbfI1jtnVCb3fuAB77z5S0dI7P+Q7bCpqfMHXXJ6c3k8ke5U34d
er379sfrVM+waylmwiv2Qi4gKMcXkrwNRRu8CqovM7xLkDzXlZitpNT9GYRbN9r3
o901rkg05+F6Z/yLw0h6Togf/Mn1Mr5b2IjJNQT/KT3b7j5DS6cq8L4mSTuhdF4O
TM/IBxrEQjUEYra+HDEIdJIq6ZsKcKGfLTS7rUHKj1mZRldE/l5x3evo4lpYCNsI
/B/6d+R0VCCdrQxDyNzNCvUb1K4jFwfu5COL8J6/EcK8QhAAIdYaWCIOYPw6EDnA
C4B1Ysx64ldgNrsP8XCq6nuhTNlSLWET4UgihG/8fEKRTht/BiGGE9pTo20NStD1
gQYAqaKHeRZ8ydHHrnBI0osoq8QhNiU27tvkPmQTMQ1B7MyxpNQQp0y6gPXjHGoy
r4TvOTxCXjz9WMBlcHQ4V3YBqLdA9SlWJiElpZh/2kVwHOwmOOIZiOGdKZ71jpdP
3fvswJkMf7P6swwpSu99p/3o9dewqqgk/Nt0GfeG12EB4aqSi26GNsUBhJet60RK
3f9NqFPu8MhtCIjZga7IjNhMlh2PSxJaam7vnSyF0tve4plEGhZQUGq48l8pEhJu
r0CdeEk1OwYMohDBDCjdTAy9w5Kw0IAlwibmnxfa2bACIJSKW4ctWju9p5e+FxoM
jSRD8YTDhhW3pTvEUCXExtM4kKGvxMXmjxSYtk8fRJxSDM/TgQpR6AcNO0ZnJgsi
piS9e+tgb35UFuycHGaiOpEyOU6pmqcQQh4bgjQVXABsVz1IVr/bKF5lAA04fGyw
Fkk8SviEgxu/CWCoLUWZMSRFtFcC43FRUFkFrmbe4MNSbB5w35eZDnGZ8ssAIh+Y
jNE5nf4WcqZ4GrQSL0lzW7Sgvz+toAHfk7evwC1b0/iOcLC66ceSnTbyaz2fNC0d
QqDOsp0iHTOVGLoePkRp0pM/UL1371SkGNpSeWhRueMoT1+OZS86VfTNONS39hZc
69tSA1VDn30HLm4AiI3Z4eoUzYZ7swFi1xHOtUVcmAVwyz2nqQuekyrg9P7M7DaR
ADu4of4+GBMavswgzbYuMxms9bvrKK4cqjc5XitfKnwn33WUynio9CL93f2OQBi8
JKQUo547eKWiQ+IsSpy3AJ8U+F4f3VqT6udGDbldMgjXbGz5AGip/zGgcCWlXCxu
zvArn4cPo2giKnAxuANtXGJg+4oXiUb6KwFYjxeAi9cNsLCsm5P0XIl3gc9maYfg
1JBdNZ4U5x+9knwivbORKHs2sYvZPX1O0TBNLwv/GFbY4F3y7f2frzz1e/Q2fQBH
SR8wgOGE4NdP5Xjm1Ve3801gZqy9SxVWnBIuy+n+N8Iy3zKibeuZ8/PzaL0+nNgy
qKdlGN4sMnp3MxIzt0LqyK9tz5GUeL2V+sLS+YuiZDSlAYEwCgXnWNXqd/r1FxFn
ADM/BnTzU6yfi+IBwN4RXzXYC45yoP6lDbaOqalw6Hfqt2wDJ2q0ax0WciW2vIb7
dda/a7jLnojKBTAl5klm0PGgWCynggsG3RNJSGmX1g9FIRlEIznjBt2T8XYC7zXL
IibgtOySJx4vKrut9RYFjeshuPxTgdtqxUmmTz82s9pewyc80ZNQ2nIUgSI1gfZL
d1kPeOPFQoXpYbAcJuG1OqAbVyvWz3OYaIxr4vFYl9JSBiCaEbvTdAUvxHuS9FR3
kLXwN1Sohe5OPEZrSubZYzmQOA+DPR1PVPsjP7dc1RNMvxgWlzfUyLxXZveiARhr
FbfHY7Vca9a0XjBID/UZnnewD7TC25DiVS+w8CUd7stw9ruYgbv5DszwXZdrlTe4
khiiHoLfXwoKu2DGtfnxTuN0MjeohokxV6KJpORrm8pg52Lzr1c+TJtSGFQbwmc2
uRVakwYL5HLU/WU6oD9Z3Ibzyr484KR/giXl8OsgnE4LnhKZ7eZsgZKNFZPr5vMt
N4Lby2wP/7OLWBA9Qkxrz9UTc3mcmpBEpUvv5//jgkngO9BQbKVLz1WM81O/DOeO
V+q1Bj4UuAm0U50l+SivXlZW0AG66w8BfxU+TUq/QdXpkKAE/KJOaQI3OMKPSZQS
V6Oj3IvF1WehuhtDcra3TGuYQ/2i2OFoFXsvkOJHfn3cjq8HEiQEVB+2J1PHO2p2
/+IYO5L40g1vU9OvS+WV2skwsBnDru7QIpbAnimaMdhsUI4ok1bX5zG6y1nkPCp5
JLbVMKdZTGP0UGRQd/rkjMXX886ep6JiOdamFan33Xe8RqrOEa20Nfw2/WMzpLXL
qaa6tsuE8ncJ0Alu4jVQqjTVh+CKYvmEoLyxItWWC9jmQr91zHkskYlqQ6KNi8J7
Bf0MWRITeznn8ry+Bgld5sCq9FSW7zxAoiQUmpakBQzUtMJjvzd4gY2m+DX4Vd5V
ZXlbiu8kDzju3w4+3KAlxa3XFPozHtTVEuM35nUAaUx/FbWYcKy72hnhWjQW3n/g
AKA/xzLk+BMoL4He81Ad/lCXtz1V5giLNxVHT06MwHzdRJiGiwFLexUadUTVM5zk
YBFOBOH04HeTo1AVTdzw8kZcE/p7JY7rNLc/v/E/gh4G/0gb7ATCotTHlMrB1ngg
pOhhYUL9eAWSpfnMWNkxAA/1qoLWd1Fe6NDdGUo3sun0q4TNnyZlN/NhvC6zehGy
TtzGhvWRAVTaXzkA1sfg05194KKOYPTTBH9vXy1kUvyPky2uHHC3/El1wGZrqKU4
5tyEEz18ZNye47kCAlvuFtuCF7XfQkz7xS4DO5Go0YIt5O5FW9DuKNjBAv5hyUoT
1lWMq6KF94s/4C1yhJUp2KhQG0dpa8tNxO3/jHF9Vsbr0dD5lv8ICRdDP0l6xQpZ
iGNiRW3+zsCXJcMmxF7/HOCdyqGhfJS0xCpMZDsEX3LExbXj/RvPEA2a2qbXIyYI
CkzAdHrPOy8V1zuv/VICpfjzA1MKTBuu5a6ezF/AQyFZk1mWrKTFYmvfPXeDKHA1
u+JcgEU9xV32EyQc/rrpKkz38h5NNpgF794mBQE7Xp3SuJbqgInGng5GkldcBSxE
OiGdSILWG5dFZMakdG9gTuE16S/PSeQkqCpOEZ1OcRbQRV7zCbOeyPt8q8yWc0JX
FZwyKgXgOG/sjin3kj0P3/6/d9dNdKu2v6fI1nqvKG8zp8URz5m4jz/pz4n63H4d
o1tca9dVfZ/CDHH0pgv6xecGLXfLA9oEB9oN1GTT18KW+smgbuiiSzw2cF26zPCa
74fXI5MX79IUk2qaKDMUk9r6uq/s51sZqTmaJrZ7rKoGkk2Fd6yKcHXlMpg7ZxRw
ztEDkxjoWewJGHlt/jAoPipX5chyK0Pl5jLj0NMVXZPQ8KFCT2I0V559Axn229HW
ux2wQeSa0RxZcEeZh4KvUi36fKsCa47xU9FJ0aKltZfEl7ECoAbdHiXfUjdUyihg
tCamEcVcjJVxK3NPEOiWAw3Gr9wvD0zPixjKOCk3HJPUXNpl+iqXZqyqLeaxfjCs
ZFSk1fzqIG2Jz3YOgsCphHjHAOQrwZXu0RyAttjc4iwQSGyuYJFdTIAFdRKE29Ed
oCpqteXVTpbkN9pRlSCwbkDM4OvMApyZxLnfJqoGF9H0MCI+OJOTNAql/0pQm1cV
zicW6dRHJNEgwKRl0s65bBfXuBqCEvu+kBLIkpb7aMCv8MvOA8D5a8oq8+gef9oS
DRre9MrXX5CHaP0E3EpR1ovJWjZsPFtjO5eqmNdcCasnj9bA8SxndUAD1ma3nQi4
xaHFxQvTlTzCoBMzzeYl073lb1rLO+mASLCSQeyj+3JfmIPjNwbcfglTPxH2Pd5K
XBdQ9xY93x0KUB+g+spP0FmxBfS05qvx4mkJWM33QjdY9L9npNWqjRqmItVFSHtp
2YDxNfPs9zAg6WYVhQXzO1yKOraXWZYwI/0I5G9iuFozerGAFrpcNgYzu9QkgVUW
5MoegtmNwvjsGgyWYGoCCViKEwIerksN6vDuQ8+3TCXwRaxuNdjbcPU34YT2x2M1
gj+e7BddBK2sTVYBsDzBe3haTBMVheYrbkQJrXMvh84SQEktc3i02BConAcyLKBp
ooccaIxBi0lsQJ0m7lXryjRosDnbgjjjqr+iRWXhknOco5/uoaY5aLxMXoj8dyKI
wDXi+n98vcDM+6xitfUXk07xi/5Ur3GwN/e3V3VmMsi5xh7jVEcfIKxwYpKvkOJB
cWIIJju10oMNxt7PqAyut7RCc2Vh0POW68y4UY/smEqJtnRh00UIVsV1vXDC078q
7pdtf8AOk7nTgKlt2OxFzMXvEpUTO+T5O/kViSKVcI+Y1/smzVQsgyYdkhZjTRND
b3LhAzNAPXMtvnidsBeD+U+ao+YeDG9ITLqYuVbY2v9JC9Lee1ePc4+zpYTC+BLS
0Eya98FFYTwNdQ/arwKLujTnMNw6GtU8A16koSR1dtfcmCaKrGNHu/6ICKMgYu4X
zEiIh0WQvODovITODH96lUBcrgLXKwNQY9HWBxgCJOs08hXd4IiDTmNKW2o7wPpA
jbYtBljjJANMXl+gZ6P3SSeBTKyW95hza59nkOA+Qh+nBgPjQVD2yZgUxfZy5stM
sXlYaZUAIAnD3Xe6cTxAChR4gu6yvCT3lridhBHoE543d4iXq2HxaeYMFCm/wX0X
Nhmq9eWnCC7JvLMmDRSRZEguCh0Lqgy4zFZfGAvtvBwiWciAYVL1fUj6/fhyzjRN
Kl5KuG0s4G0g0TSWSqEmtoS0L1jmAl8bJNCRqmDjSkd7+ECKzMTf3H4rS7ZCkcqL
pwbGMTmJ5BX/A+ZSeMdqDMIMgzK1/xJo5RzKLNl2Gm6fHyGyXDF7NlRV2qVyIMVj
tZO0obZADu0UYeJU2Cwd5Za5davP5h0Ji8IfU8DVq0tdgFbTsiDnsY0nUambFf+M
TY6bKCoZmpXGDNLHdJEbyuf0rnZOWX6KpcqecY8EAm0Cs4pPlHlyeq4yuF9IDdyQ
6HBXJTuFeh/3z59g/s4/F83EsfhlhP0StDUwwcr6zNY+uGJUDWVogq6gfXj/8LiH
Li4LzZrr63P7x7gk1clQYIoDu+qFl2cZOk2sM2Tz1Rw2PH7WcGcD9Cgnif22x6LK
VDUONYz21dELCP2elM3vvJDLbrhc0+DOUJR64il/XGNLNB2sFY1xf/TcqEgFT05N
lww3LPzmaVTq3+eHEszts35K0Yd9gJg65JF639heXj8JihBE7C76eqvwWZW4NJFV
hBXWoP6JtgbuHI7XcLCyvCOI2ILjS/vOngE6tMNaAeH2+YCrbcQ2MYvtASjUiPvd
4f5eCjuL53ZL2URwo2r9v0zU0662M9yTWQFzdVvmhJOdWsEtc+bdlvA2k6ClfpJ6
8af1dAuHPEdjPPgIhcOh4JNpdN+htynWgPTzZR7ye6UZKLgH15wIeQdE50RW1+tO
myKmB+9PWaXzcrOQdLx8rTeRKocj58VB0WsBCycQlltDohXRb86KdpXTGMJIxTTN
Fm/vN0PdHY1VyBIEdy41irQzmF6L2VZEG2eq5jOsNhw6OS6SXPG5fxK5dRiuOZOs
i1DRDdBxuf2iXWEpP6ME+ok6EpCj1pXg96u9DcrdwpXOEoghhTVqHxUyThyeaFSo
dRjbyonjkFnSOvmmA7ueYJl6UdRbzMRw0yYi0fbSTiwqETDZ1npbqL8WMU28MUyQ
Mn92v0swZzU+14R+ko1+NND3eRlftXZpJYM7bR9EKmIN0v0cSEgiMz/Zv1W9yXYP
lP5KtJOpaaOBjqiTAC4d93dCN+mEVcFHdect8KbsWQX+6lBni9pIQzqyTx0L1Xlq
DjEmTxjBic34AuefP7D7FYjc3YUWZDJLjDpOwp3T3hWogEPSf+c6uTyVQGv8xn3Q
Gp4TlQFB6/cFeekMR3Y2EGGwVkIomNHnK/EhS7bn+BwX/M6sJjl/5Yku+XVFiMRT
pYzbznmu1X9XBrS/i0jBfjp41HNg/dFpP3I/Xg7f/xrXD5c+iQq7aX1XMqQTiJJm
9rIDpoZjwD4sTNPVyRby5kkp47DTTuKvnLNkWd4vMJOBt0bwcRoItWk3H8ThVirP
KLliAFKVnYYABTlkUnlO0VwXgvuoowdzum6Xp/N8yHNEipdOMSiLA9LW7nmoMrfV
i3ysfRN0uuw4S3sPvZ0rBfR0OVdAlY1qUTxbubPhH+q55EJguNJzzuT22H8TyOi1
TA/5Fkn+1U31MQFRQDTOIvNhI8uslQ9muGJOAAXO11P1ld/dKOEnKggrg6qra7Yq
jl9sxdBv/xXo2v+LDAI9QeZvI9LOGRol6l+AQmC0eAjOSuYzhxGmaGIjtU8f2W+l
bsZ5OLr5WpWE6E3J3+Hx6VxiIL/2aQb2nwfeLXvX6Si1LcRQ1sCUeUY4/gLinHqx
jwhVygBpuL8w6Me6JlSgDKgwmlSXSMi27kEeVHPOY+1AOoeBBZQJRqpNrvruZnMG
Fjh6Ko+Dl/hg5cLwRTscHUMvX50Q/SJ3r/6LGjt+sej6iLkPevHKP7npT7hJfUyV
lu+UkdnKBShsIM13EjqpPTR4UtHiWefYmGfg/3k6UFXz7l8ZaWQij++36unsLl8E
uQ53y17PMKBjjFsucLDfSxjunZbhA4XLuXDePohHjK9/WnYu25bjTZhQsjefIIv7
WIKc9yxzb6U8aQqPcp6HqSjXrH6Q0iVzxRS6hdVri1iBEFfa0D5ANfmp+jiyGkjY
svZSf7XPQCssrgradmINQOXfNFgwrVMzrsKv4ua1aW0r6Zq84eld6rt3QWSKMD0A
Qm8nA1nsXMke6CilQmnlM6ZNeHUjZ7GZ3ioT9Q4iKsnj9JbtLAzH0St6uARPIyCG
PZNdH1LeM41DWzvBGDX91B7AgbKyIdopfoKfB8bzHbPkrG8k8o9Bhl67q9B2xsha
O8PJgs6W0/9253A0Uy0IrEJsGaXXwGL9nfxcNFCTAo85dM7tZr/JbMKq1Y4CP1p8
h54HvbiXG63qR3m5q/eY1439UZjET4wBVUxg3GUk6NAtkx0fkq6LDgHaYFh4kffr
OcyrAbO0H9TEgBV1IqEWolrzDXTqJBa6gAcceCHMojkRa1e2rqzbXD/urj8dgRa3
TOYI1+9siHkeSrWHapCrcVHsR570MeGHvOHMfYnQ/X9qpkS1/MQTtRkQsfQ8fql+
Zg4PQbvcncWrledjmzPVMeJUNtSTaFwVQjakQf1komgbw8Go2ugEoEqjb/8MgNcf
7XEXohDhV7nXIVYJy8uPKutRbkh5TjZtgUNt5JdCgrrygg1AvESAltS3jvEI21uA
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VzMhWCbNiNWs5sLUTlEVnlFnix466IvcOjZXvsC6qhqgtIXSBZnRpdqIOeDVl2tC
ovGbi993kVVyq7Bm5C2bQxy9+fLxGNwPKAoHcolhSBImtaBRNh+qIsZ+Y8icVpIZ
4fLMHBzzWfDmCkYgVx1CzqzbmVQgy3vzwDMmNklxNPHsU5z4/boXIqiEwXibs8Hn
JLA3QJ6ffs0/3AKyCMxNmeEHiBdVyUSdohBaDmejAL88fBRZ1/Uk9QYtotpBcqnO
zdmXLQ++gkpfG9+/7J2tuKXOzO/PFhR3YYx5DlPTKm/tR5Zp7+tc0Db4mIuoIB37
otMsx4IyAIVZKOVbtGL5DA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9200 )
`pragma protect data_block
LWvHc7KyCLLV4lNFpQuDDUozGS1wKRf7It073QjL1/BZZ86fC5LlvjOOkEpbvRUs
z7TSWrZapYA9QGN/iWA3cVzqikTIe2X+uuPJBJZaXBVCC8Br68odCqBcp47rWrk8
zRtRN9zXqSFcQGxwSWihziXgZ/cJubv0NskgqFTCZPrCkwU38TVtmpXtovOVUc1Y
02knd3hDtbdDA2CUpl/cGYlIuN4gFuPTq2Gg7g9sWe6reJ6ghjJteOB5XZTwFuo7
rkC3ajxJYJPsyly3710YzqdvyRuf3WlMmo3NO3LP4RjtWAwM2mqw8SYOQ/esguTW
UU6mx//0DKSWXvAZrrBWwCs/4fvM4FnKUqvtpF4/M8HtjZMMBtt51ebFNGwfQKDu
PyJ6Tkl0ckYgp4ZLIpdqZNSoBnyn4i8V7/vGV1/CV+V9kkQoavTu1q+VOkAmRSKz
I+YI6P2XY/0Ejlfo3xSt9YU4j3X/gc6vkrvwVbJ5aIIY44n3FZPRLuTKRZutunv2
boCgySVVDjz/CBNs+0hOLw6BTU3+Ee99XBmnVcMLrDzH92BG/W+hLj4NSWMEP0Z8
B4dEmB1qa/glfEZXf2t8Zy+3WHClTB7nK78Qmc6yBKgleAClSBLXSADEev4hB9qS
uvXRj3JaaWP4cxeimx2JrT5+Uj6yFqvO4KhG21MaDp81OpfBN0Fw3+sgjrLO/P/s
GREWZsWDfSynjkuEpULzC4YUp1Q7URryt4UL1ZBYIbaWiJKOceJ175dTdpxhv3dP
y1yTE3O39ac8zQm7FlCZTS25mSW/7XdQBBp9xJrsZIl9AlVfdap24xsuQYzZzzaa
x2Lk90Ng544MTZihw02JuRk6Hj6QE4AnHxqSpWg0C3RDLGpuqhZwlGc1h7rXTEg0
E7DFuKkEbPbtTrnL/iiOuSdpIKO6ZomiJywwAhzYa1mFzsv7rIoMoYIw1xzF6qn2
r9GLBUGWiX3TGntmTH0M8Y3f+sZTJ+ryEbQPXC8HpJ13uRwFXMVS6bqIVzG5Jz4R
AHe4NH22KKV+IJ0JxQzy8GiWMDdTaDpzbyv8A9bl0rfd88MWbM6lvvPz0GiNUuJI
H57OlAUck6AbbC7dskMUCTvEvlgqwLcMiFB1y5nBmFxDgbZOrz9UR9RZtvPNmrLa
IQgtm16mRRWLQMXz4YIWPEjVEaJjaVFQ0md21X7HIR6NK4J2dQkcrnN2GSbzPaf5
2vP9H35juxclWQ3w2MRSp4UCYrHRcZdguXoNIUJQH1kNHWx7hVut4XoeNrQXg0GL
5lKUq2PyEi2Es3tkSifkXiCukcdAIXTM1CE0kSZCCe/wb6xwBXePWSgFZljSfzTO
ulLt2Ia1bhU3LVzK4vvybWsUmeQVfTdrI9QG/gq6GkC/jHYjwDvIeMzjNh3QcY/9
BN2cHUVDzejY4L+oBw/Fcwfo+VfhnBSPptGuRyJHr/3Te3ESQGNSf2og5o0Fog85
k+SsrlgpyQPOzKstVDfRikwPVrVAUr0GdJqv9o27bsFWhWuc0iUnXKbDb8NNJptN
xA8aQ+zEm8j347Y96kpawa7IWhfe2InAv+F40bX6CSe9wv0nAqrUjDDnnJ0U4Kt5
NmNI1yPVEfXLFFF++8aJwLDLwSCWiui/VdcWOlWxUClvdWO0lNXYeQMs1a/Sxvs8
jMLu3cvXNa1xfIGupAlJ1DTgz3rUhe8LceEg6qVlCkLqvxSAjLG5zOKdG4eDRCsE
e/JXsFtGR/yBY5EjG6WWpu6a9ZH4QVByqCky7YDHZ2ix6+1D9nHGNb93p0DTcFx8
3ZEr35ezb0ZkSOBLqpcpXn5UVA/7G6BSV0IOpGd9XVbRFI7ZvTbILaqq29B72Vyh
7qpqEjkl4X8xt+kPGPEeBF8lyYO4FlaFJu9Ykdz3RKl3fg/y4BPnQEkCHa55qm0B
yEOv5xuRFdOISpg4z4ok9gNf4v+kjOYpN+jQrzdedC0w2nsv1ebrrUPUHJmaK5jB
EmTE6Fqd3uoKGgMUkNySVk4bY5MYXannGR3j376p8OoCAy28IujbKcGwaG51icn+
4Ub8lmH4sJ5GBHlhvwtNFQluAFk2SV92Ic/eqm7T/gDyKgeNLeicyc25LBg55zsW
3LR3ANlZNAzIBRic23zgyw4jIR6MRJTgaj0OLWRykpW+ZMl/piuX9sHflaxKbt60
2DlfEkDDXUiIWQ61l6SX+88j93LNJSNeiuabInDuiGFwE+YF9l+LPa60wl8bgPcY
iOmrXEVUUW4fV4Q5j2ywbtJJmk/LfPDOGr+ImF6MYblx2lnQxyToWNRA4y01IstB
cNfAc6FY6Ky0It6/3qCS/zx7VdpnMb2mvZNtZx5jROO7pk2UnZ74PKRJ5blE2xC9
0OJzPUG6xGcncrUh9FlP3xIUsSDz1cIwMkFeD4PUHq7EWDRPhUI8/irw+ZH4PcD6
2dUl98w2Y85S9/3uejve4nUrXozuYrw0wBW5Ss5cfAXS9BYriviUXh++Na+VZOTl
+qLv4wTNVR2FoBGPsV+KirOLgIRG1acV9Y8gJov646myPu3z4uKtCTtRZIbx3cCy
u7Hm6VwUaVj9zdwsABif7t6ANrMYTSKx1x0aoMQZuOszl/Ue9QLkdkkqqLgNFK8R
BdG0npdeN/Rd3cwQSJBjX7wBpvSBt9fA58aaP+QtXjSvx5A4F+xk88YC5HEpRedI
A5jKlFDnkNLoQDdgRlAAhcCu7mQ0gpaJdHkmBTaVtVO5gvxOef5a4a6IvXGS2/CE
x84/UKrj0mIyt9j4RPCe1P4lJ/dCbvlzqzNkPmiUipRSY6c7irDHEsKuAjYg4+Fm
FmmmpMsVrLkGbfoSbkhHU+qjFdmgg8/mYHUBqzUJ/AUvriMw1heEqmts2oJM+4ek
EW8TTTMj3xY5V75yTTJROq4027luYdacRZa0y+JnkMMYxitt3G3fxkuzpzhqYzkZ
sl6cjW0NVS8xeS8EKND4nxI2b+aCJdtALFnY7JO66zHk1VuY5ZHGnx5Gn9CqJ4gR
qceho5xlFZByaGoByLxlJyv0SlLPON758Rco34iQfl1d3RsRzylyj5h6625ti15b
FGBvOzPYJTnGzhckBS+G174L3Noj4FNSeaURhn+1RsIkxY0m//a5eiyWaX/QuTJl
GKk86SDri0vNpjNU6EH9qqmx4RxdhUXtiL0jsIzNa+IeRImAJNK+0D2fzzK0Rg9v
RNW+TKS83cmXx0NASnec9+bMtUoxatrLJ7Jp/Q3/Za5rmXlIZ2xmWJTY9ca1B4FJ
BBgWP+eA0Mp5G31I0k+1qMY2/YZPW8eOXnP7I/HtByh2PFnOj+TjIUu4kGTrRn/B
1D5Jn/aE7yLxGjdq62K3bwl74FQYPRdrABHyFBjfO0r1TriuQ8k9eulyB5woEpl7
joKUQMoubeMkj90egtI2x6KkDPg0S4L5pt5GUG754WPIxrIAi3U2lC40u8D1gVrG
QVbeXcJTgK/yD9mwOAaEN3fHdsjODvDsaprUZHVoo34k05EsS/RzzXBMToymhb2S
R4wo/f1I+6ZZAiIcldb/HtQoZQNn85sZm8D50bW27m1IBpdlwcXzWYpdg5L9AUzS
cVrFQFBDGV0owscIEYRLm58XSPkwZS9Stae2CHiS6KWTtN6d0PJzpKm7ncpsnIcb
C9oCPQC0qwjaUfw/gctCJrGsfY8MWfU2/oiu+OT1003DrscbVRZ1smoA/wh1bqgC
AJOFFmdQpdQjEIibx3hZhWosQesDUwkX+1i/YzkYx7aho8llTqC8yqTCr04Y/JKB
r2exYnggrUCS94UxRyz4PKg06j2JYtIDjXfvW2BWHhr5S0nPTpsgXB7qNDbWojZ5
2h8qge3xbo6FB/GY842u6Y/2AVrAkATEBLIy3/Ma//B/N5a8mGo86XRr4Kfsvusa
KVVbqEMcOWTYXQiPzUk7iHN+VM74iIffYQf7QMHhd171Hj+XtEehURNG6hndUBYZ
tTC+EsJxG5mF2ih1mxcZQnv1USchUEqJIelIoC5jWIpwAzJy/sUvaso2Ww6nfZAk
FJZe2u80iXZFj/CbqzFBP44yLLIptdC/YUFCHrtnRY4ILEbO5wjJEAfm+YNELzfA
GDbnJCNmCQ+HTLL3833iumW0nJw5nme9ISRgu/zM/CSP/I+ueK4SgpI87SwC7lTL
ZBGDuBIjyJt94gqWNLd/unEiTqnVSSQge/gIlw6aj+Q/6UB1c3P6gv6sQMLxLGhz
kieOv+brOvL/s7pz7czuvJ9ow2Raa8ZWElMdZqPNOF/8KHXM15Ig9OmzA3Do2t1M
wiDkIc4kleDMChdgRiOYYGPtqp3v3qqRduH7P1ObmwnKEsBLzgNxKmkekqD2lsjD
W6GNXzTHaTMe+nFeBTK7I+cMbFo1g0VFbPUOorC9w5kzz3p5cSxUYQ5lDNTrZ89M
9LHkwi2Da9odn32w/8uGqKCc0EuL8hGm1p+U3e4xqSavWU+qaQjTY4fEfzblvgzV
0NQB88ravFmMdgDA/nYeyDnG6sQTIBHInpoplWXZodg7v4lDPWkG6r9fy0Fy/LHl
WTMjI/iM+lqZfQqX2DgVPoFIDbsi19tYCAkprvVZrKds9NrmU11wIw1U9jysQfxd
NDTzYqre6XjOAsQZnVx5Mq8vkcOsRcOb7mnTe33nH3ROlxFEa7CcC6anFU/rysjj
79b+q82pwXaz69HKabZNGG3se9nY+asFAic1IO5VA332/lUN9d+hHoxksJoKH8M/
m7NMUg98AHQT+MHO3HUHhJ2FwoIJZR+x+uKi8Nmg1YquS3Vr25BXI/eNQj7q4eqI
xEGlyPhoPO4jygtrm57xdl4JLSj+WA87bclxnWPFMX19VTj3YwB83GfeXNV3MBhO
qDc9emw9mEAyhrdGPnWVzrWApbEtHHJNhsFTuXLN6m6odiDzhcLL/8EfofCkCiHr
P2wqGm1NdY+QoFET220Yjq/7DqVb+8UbZDUQpRsH4gPuR1WSjOKR2/JZAMLC4qH6
lNjoXjTbOeSxeLBRmHGLhg1WDnUfJL35TarfoSqa5Q/w4+VfodmaHjmvY1llI/sG
x8BphINXjT9mQBJtcCErH4PQXGAqxTMDN09uxExjP09pGuvnIH7JmMD0gfQUFXjF
qcxVMj2Jbxc96twFyqNLXuQ40Be8M9eZnobXuCmOZT5e1Mkr1o4kdBpWdeSogvfK
Ynr3XvE2xYaGN6pPJUOzgWajK1SiZKLlQcUVTB+evrF9iplTHY20bsIKDU5oSqad
lAGNZXkEQhlnRrQSKXhlLqicatcqjdMGkySu8Asn62zOZTduwclumVq8vj51IvZo
zKOQjsLUgzOrAPNSg0Q8AfqwNjeSPk2kAxwAzv3Qfw/127CFMYZ3x3bffiPdD49H
pb3DwXkUM8ndX9QkBgrzArZ70IfZ+GIFJ03x6fLT8agSy9FdAUApUGT1oGD6TE/f
fzrjudKqh0VpYWaAkmC+rYYoHUV6L/88MJd88zBaraTElQexCRNGOdRXrbjPR1S0
UODz59UuY7ER07zmP8werueMux2lubdeuE1sgGrYihtieRvLJQ1t+HU8QGeDW3vu
8rXI2Mf+EUWA5376DE393i9g9xhSzu8NFiIhL/fgQ+ozgvBJR/lntt9SNNJ3Sd1N
7bkiXXRFfDcdyzublbRPqT6zkbmd/JktPX52ScHWljngAusEUvVlb4JnrCnZgrT5
im6ztUM4PwuL9lmn1fR59DaEmTcbC7kirIXtJA64NdktG7Ml0y7/poME1otpulw0
4R/j5RXVs2WGDC+FodXliVsfKRxG0u99+QEaM/sq79QXXsDSx/k4yqNfHEl+zs7Y
YfDSUmBlTPiXDyqsk9Hyjzhm2Ike6CcyKlfV1u4hrqjA9hFJWiuQ6Fu9gFzRvWaC
yRt2q01DXrPcPxpDSEGdV38vZOjXr3eo54DdwS58kkllb/Z0sF8qocTLtSoTbI4y
y6jDKFfjeYzKfg21nn7o4IxlpKREBk9nXfpmBzL7JQEfXXtycbYS3CnTuMxOvatv
RPEvwX/LqLj+4yrg69h5W7a8VjTeoqSDf5t4cR2aDCGadDizpBERtWRkGX5z09uV
ePaEw65w6eMDtRtoJEcrDeKvyR8AW6cO61Xg6ao7XDWe22iC7TFTxmByEsuEdUA9
Wx3z3u2uQAq6B+BIdoWddypGelFqmtsK8PljHdenj6ATwh+9raP7tHP3CH4NylW/
xcWXh31K3NI30WPMWFg5VMLVj2FF4yCblhH0uMTRTk1T4r+2Kfddih1lROd7dGV5
g44xGtROHTSXdBeWcmmAg59820ZORoVYUiivi1KPJdy5MIdKw6l3NXml2RmlTSkI
qllghH/FwNWocdmTFzHeIjyno5MpCtvHE0lCt0zceY/aawZmipySHsQNMr6CoEIN
xH1AkAdHGE4btbyllQUcwdmo4zJeTJ8gpSGXxiqQHGEmosjsCtQKE1iHhpiSkkPj
1agTLSA5YqXzQJ75R1gh0i/nboBdOj9+cSOW6wKDh5oXtQ55UbQvDwveb2P4omZT
M4dAx6qWfFPrz+eWAfGMILncSmhu/gvCtIfSK3aAKyis7zbjxZTzrMnTtlKFrlsE
1WjKpEvrYaEcoAkPSHDCSeOWgKrP/hCSRDRQVRQk02775QE1I/jnv87pku6SnXgx
bXfwpkh0n5/v6JqS1ayn+eKwYrlWcsvho+d14N2ggC3Wn7MJrXNs5VUaB6y2Egyz
dZhnPhSLSouwMKijoI6aE25tMd2gx/mWNCBSh0QOM606m1Z/GysYKCG6DP264Zid
xB+gtzks6XMcgX8Z+J2vl+P+vyJa7hasWiYJNMDEr3s0woqHcWrbqE+N6oOmVF30
vKC8QUdSwLQeK3djNymIdT+J/ZmYoP6pM9ut0BoveyVTIxBHIsR8CG6x5en8dWzQ
0R1ryvQlY1GPR0TmnXcQwWUSLhAVkOaB77agkRS4CTPfXh/wuEOVdYSEBh0tBrnV
nnb0Ex/axUTDcChOyiKy4VWIQhdSsOQybrWFly8XWBy/7GyJxQ8gi5gNVgAS5Do/
wq0LDLwGPDEiWUjPNdfFpBlXu80LgHTM1hq6OYSZp/IXnDRpsy+DLDmmEsMclYC2
cG9nHBatVY2lY9WW/TpOnecReRJ2d5KJcHaQdCdwXs7vI4fz0jyBB6YvjaWGLnm9
C539znp3oURvNXClCHnyWk+jBqTG2NJM8mm5YaROu19sFN0HalP3dsgBpwtYHWn7
Jx9raNrV7nzR6dnt2kMQZRAp8pptCUjW3MAs1jBzK3BiNfKPJHNKGy9600IXnASt
hQuKbOaABlMHE4u/jtMXE64GlVpQfeMwcFkFNjh5NNrSURVhk6dNwsWD4BlGQz5l
BsZDp/k4w17dY1vGvWTKZv30HJCfMfRKaegAtgr+7/w2EAhIjIVGZU7kO479fD/L
GSHkYjFBjOI09r2WSb2fctHwrvH0T8OteEBKwpfezcgWCfM1dhdK4rlbrJVL2id4
eCSkNs301Lx+n1N2r7zIV99XbBGwKcniGM+9MrV+Go1OmqBN5goXAvnquC6iwQMq
XdZWRx6w4EQb2lbdJKk2fvxBpWRMJpo8wRAQ7gVszCnmeTA3QIXvdLAgGUZzNO45
rGRETDRfak+Bfy93Qe8XN11ajKsRVz7FRenAJ3qnywF13Db4rdgoFI0aifne9hwG
OesPivHBlatuntwsepg0F5WN2KoKCDTqxGZSTR/jLAnYKXx969xm+kqJdm0fFyZb
ocP+TjWrB6z8SMwhIocOaN5YPLdiW3SFdhpMbefCLxc10YOViqWkft1tLcprdLO7
teNENJU49wFrVm7+KzZkXDBYUlNksGsMQylFwjIvDl+8WY6xUp3PXjVKJZ0RSMJw
8Oo4Tq9VO4zl0qFFUFun+Tdd2Ax49CrQ+mJfmpFtHOLrDeipv7do/pZywrAIJiBd
XZ0fj01Ys7/BrOf/CKnANKY0rjMu/zTXHZKD2aCfjZmWJH8G2MUDKF+QOWdYWfKq
SiV2kuCCcgNuiY1SzkPfETtHYQ5RR0VU1BZcBUDOU5YFfiJwNzpSmAQZdfOVMLnV
2GQSIMFFd5xGSVTXGxhlX70nHUIENBPioWsmaKOm+FdoHxhqgHmwJvO2ZWDtFUXu
EWRJni8YNF4Nb+iCgLQ6Ue4PTpUjbPx6Wz9tb4LwLSBx4qrbujPVLU+SXdhZGsWq
A5pMHC7i97JPNLTcZIkvgBNbeABzVEuaucyP0U6o+raKg2f/Xhj+MAaT5fDU4kvx
Xo1z8RxFnJrqCRjaEG9yFUVcjuFJUea2i8iVI+mM62SxWryRIt+OB+pLN+pwU1Kf
i6AJCkwUJMQOS6VqxezKCnTdIY1Kl/7ECngugd8ADPgcaQpVagFTbDUI6YGLQFz/
EM/l5PVuhEDtFHBHcjFFP0ehVHTQqF6vVpvwKa8QX9aYb9Bof9bVvPyWHnFYVXnQ
WxtkCesDt3yuc5t2sjJAu1yHI87TdwjEaEhGl4J+iYh2E8PgTchr5dIuO9VNd7PM
vPn17Wj3Rpn7o67G6l+XLNEXnM3Y7G4WQB8zKWBRw7pjGgssJno6t5raekqNa0OT
zhrqC5j75EQD/M3D6hXnUJNqwFJ3feiWXVGJN/YQ5SI0xJ2dXiKnSIsiqy8xeLaU
ojo9GZLss62Et6LrqzdRLRPfXfgE9gQYEf/Ooha0szsk/HiqJwvV2Y/vsS/4Cf7v
aLLGJ1Nvq2cbwlHKhEkbpqqnGrk6XCQAONKuEFoH+xIbdZLqlsQTuEjZGnUzyqnD
2X1l0eWfcsFq88mo683W+dS0ip8xL4/0PqZQdxyUTIlzhMV68dWst53wd0euOz8g
8mla8ywBygGRIEFWWHWQT8cqAqsPGCHGQiM0gI9WK3yPseFiwd15kIkQyucWO6fv
DQL8DinlnIbeBO4VyYwVy9r8OF4zq0qI8n573QqjrzkDfnS3p+jhaXCSuWcxesa8
+LtrlqWzanFuvtMsjjG5RL573FWnLxx94mTOcMGXV6VS0TgEu7jTCzXZsUiaubWj
W269jnbIbdRasOOJxqtyeiUijs83E9Pny1/rUW9WXVNOHXCOhH5ZaIb0yuGbEWeA
6ROPTe0PZdlhKTabZDkWtXUWlGueWka8UmiVPFzZVjMjpgsjgpTBfITAktFJ71Mi
MdNMmHO8RfNjHuOUD357s8OdJOUkLL7YgzPoX1VluZxhh/na+tj9mvdK9wlSmCTP
pqieNe0zwQ5frXs80asWZ8S/9N0eUOon4TvdlWIZn5MEbNtJ464mf/y70zlPITuf
pM+kTA9bee0djPYLNT0UZoBAwNmvcrJIEXuNCVhUk1hVbXmvqV1E/d8tbh1sUBZH
ydMS++yLuKGtC2JgUAprvv2GUihfmbOo6DJSfw6xqU6O9FYBTP/tObkghgczMDvu
G9O4XzgC/+D+1zACU+PURO8j946aHC3k+B2Nqt7gpy81BvfrIhi0GCmTw1UF644V
EJ978faKSY+BvM5EtlAo/pm7/BhU1W9qXVWvGtiXlS/PlKJ2T10ctLp6yU4+C79g
3x4W5fu7Eqx2BoDnJWCKXLJQII4DAJfpJvJmFBj3n36Y4oXr17gF42mz9JRwxlpf
nQdnAS8IpMK1fXTfNPZlLN6EtSCGG62R92gVZOnCwgEwZLNuwvKAaIONlqH3/xxz
svuJhTz2qByIlw12wxk+Ip76E4cd00YEseAUm0z3j7ZWOIwNB/m2dkUwez/vHfW4
9tAJyFW9xq3fywxFYsd0X9NSVxI24nMGzzxxoy4rSqFoIfYwsOSgl4PMlN5qshY3
dr+ze0his3TFz8Q0Jq6cmDCLtuJfQwccGqb2TNbZ3RYtR3fyQJYcHpk1i0uhXsaZ
9K9WaZENvCuyzC621kxLydzhk2L5Pp9CjDa4y4urLIV3g36JMEMX/d/x/qWMD/ei
qsjlQNLYN0aaxLIPEzHcRQV5vXnmqHaBvlzz61ouFQ/AQIxLNll9j8cdUpxqvM3a
dO65wFibusqZrk4E+QyOP533XI58WkA2ilFFcvNTolNOEezHWvRo7XDGH2xj9Bl0
sZb0CdywvgTyxKKtgiS7RO6ScfCkFQspHdmTxzbzZQAQwfm4WMvdGs4jJ64qDiHP
k5ccEZByjJkp7temX7NUGZGMnW9zZZmdsMwSx5f3yOmAP2TzmJVRKdlREZQQOkHm
RQvBtUzMIA9Jwjmc68UI4sOyFnLn0VGVvpAv3wjpHdWQczhLH6jKA+op5vQrCtY0
P4+HUD79oSFNZJlSWaWdBfcuWbY39E9y+WRWoXcLCs8TkBCW0C1/Z7EDGF60am6z
4vaTi/dLo2PyYblnOT0/Q0FgDu81ZvnxI2LkuLrXf07geRz4+hpPLS9IFbDUPUOm
Ws2NTYQNDIZ/m1wBxw41rNfU43K1jRnJcp0xNfr2UlOB1JiEpvr0IJ8Azr+YmXxd
iA14JCO3C/Ud0Brsl7WCAVyz1E35F7siUFMC2yUW2AP5yb4Hf06t1tCVNxB6xDI0
+g3216p5nOTK8G4xko00I57T73sO9UIhZi3iyDKFjHDyVEtrXYXgiEYR1URaoXdR
Wun/SRjqoDKVP2KqwCa5dBvK1kvFW41u2VWEiwI9mJPZ9jR0xo1a08ptK4wN61FL
tzsVr2p+lCzZ5iGocHT90s7NedSSuGJ8X9qnjqunzyXwaRLmeFVS5DPNqzBDr0Qv
++NQJzcrsrPazRjgpfXg8+uC4YVO4xQB7oUiIA3TlZi3Wwxt4ZldfnavKHl+10tr
NHdBvTG9oznkr7Wk1tPwu7zpYZBqjXPVv4b5epA6hykrtukv0krE2o8bDxqRb1Ow
nN1RvTFzdVVsoMaRO+FDnTTlZgNY1WjtOkvF0eKaQs3g0R+Uxx4+e9AXPhYuqQgQ
FdrADwNHRPVCU9EOkgrZp3agZF5P1os9bSzp8fE3J1moyYUAPsOJCLEXpo7nP+ib
0sygw++nbhtx0ilAAEOeSzJ/FdV/t9Jq8gZ/YE7t4hlDOglCDDchgqVUSnAsoImP
sLB4snfQ+PhG1FQMSzPndHIu3Wu82IfPElF43ejm6Fmt8rDFkMIzgpw+vuOQrvCX
GCpK5H7OcIkmY84vn9IQztk7+QFpMwZFckN4adgqHh55tPWWk76KMkgKVk1FNoeM
+8vflUlKFsJNgd1AJh6jToIXN1gU2cdj24pwWVpmAfBNB7u/SpfEQMYmF5Wgr9nB
OO7vyuGoQ/Vk4l4YrzC2A+ZAcCdRn3BxLeYmo7ZMhcHrX/4bBoB9vlxv15/T+2Fh
ZdXGmpfZuR+cgMaLRrCfZzf76+LsZC63ij2IE1MkODfn23OPXw1oH/Pii2QXZHxm
ZsQFfRN2dOt8txT4cr03UXOWhWgeDM3BDh8QDmkoUHlpaWnCRbQaPpRFtrAGOWWp
Bv1y3PBabW+jwckHuVZuaof71swqkRIkyWqigpBtZIb9CJ9xQnRlzjq1KzsEsshp
YAnmOft8JpuvJRH6GWdofxh5AzRtr+CCBgQD5HgYYwFYPbfX24/pnprr7WDuVf58
h+MIfA4Fqz1+de64qUoPTV2X8e/ZC3YFlSdtnTIGNSHXNIBTUoM6rtBE5OsdkJo2
Us1lKJaQ50EHaXQvVSd2wjIfO+/cbz91xdXn/6oLN9DEwFgdXmXsOGEDn0BeE23L
tlcxxXbU0n1mi5e7QJIm0SsdBt/wP8VGWvdijw3GQ0BhKA80V1bujyfIyIjsIVRl
DBa4YDs28pkWWpGyNKC3ZKIutJdWeSUNEyz1LcML4Vq+hwkR/1qns8o0VeSIUrOY
61Gjvh5bv+ahs2TvHoaxG24yxc4L5oL3S32ZwpGUnu8GtdOR0e73tWcRApKGrKNH
IiP4l3G7ZfLOPN4L8Y6MHvmPYvqyTmJTJtIGCgEWxPX7tdoaBY6fv114BLtXfM3N
Q6I0GVphnTvMISDLcs9KKnnpgEd/eLheXzs02pEwbTV0OWLdwPOMZB91yHvqTxA4
XR2QgGPaEQiDkCbYxtCE7xafCNvfXEGvykO78ZG0CvZa1uYpqHzc0HzT7k1KC1te
GDZyIyyp6UkTjftVNx9oC5cKQyH+xFjVH8KzTh7Nz3faQn6xmjh4pPeK/aSBeDSB
LVrc/mmG+BWf8zSt46n/mZicZokDZx+H+l2tnY5HlFFYeUeFNLPpg2X0DWVJdqED
xfw+YueD74spiXEL0PjORwzsBjDf8GSSBhVOld0qJSaV8YoVd+Fr/STWZFadYUfH
xfoCnMegqKqeIs7OGQBn7BPhYri2UUhOT3OirNJU45Y=
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
D0qov/DvaMtI4ZmAnYLfBbPznWq5uNtEOELbuQ3YM8dIJFc1JhYS/Fb4U/zlBmtM
rcXTQGtKsYpLY63UksQGChUWRRBFzeuys2HTi7YMdpoB03V/DUgjh9myVk8l4NjT
bINFFR8FK5FSpzH/HN0WMbFwT//Avk59X9EZGKCiOKeHlm9qXs9m+WqRYaV9bzKq
CezQ7NKqiB/JX7gItJyvHhkSAKoPCCvQ9JdKDnyWUhwpjKprj6iIiCmP6v1zqAsQ
JuJLhqLk5r/rIM7rJMvZlgWKyuOhlePWJ0updSGLWXZFovo7sXb7zkvQWeW8sPzl
CcCSPL/weFj7ohDwqXhrAg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 752 )
`pragma protect data_block
KSipNmDMqcfzVUkkKHBhaIiIWQ/Chn2v3nyRrJPUV0RqhnlDFaQHUm2E49aeo0cL
Z0gjil4xjFSFMTy5AHayBjGTO5OR3XaB+TIsTbTQA4oiC5aeOlTisbTYPYH8Iw8U
cGBAlwpajrTzTvKy0Y72fIjurueohi8nU85/OLcGS3UjFpMtJ8P/yfJeSeyiGtr5
qr6a2hKYUJE2JskjgCx/qoNNLmbpg/j103SNITNH7R/cDe90e897G7LUgYc7HT+Y
hNjx8dTay2mulRUECrI89lkHBFJGdmcjIZHtZnzPEDoWpV9CWKalgCViw5Xf1K9Q
TKy0AO9IqhERpylfC8h7kQcfJlx6B30zPePWyWyhBcWFxgT3R+3RJwAIYoFPPbwU
XtbAkO6KzPrmxI9VTCLgy3vcvPqQ3FZvEE1W7905nQ3FTIxrsscl8eJYdX/0PUBn
+6f0YzEPn4vRiAN7UszJKPALpSVKEJdwZS6+dR6eYmxdP3NJstrN53vX2/dlNTiR
aW2tbQ9xE1prX8JPXx7U/vpxP/U2HtNe45JDwcmIveoTiNZNdthdZm45lVD86OBU
EtnAazUrLFYz5/wSCFVzuhR3OWnjz6XufJbz/MK0gxhA1S1Sl2f4S487QWAlApWk
u9r0ewhnbnpq30P60LRshR105LcY3jiGsGhExn54L90VByGuAEaU08o7DedvOXkB
gAy+zs8e4k+DrlBTVkav95olCmoJG4fA0itN31OqITfg/WAS3+5qL+DtA5vc5Kwl
sf5dgreJPMvPeif2bmNiq42SOMb+8BAyvnqqPxudVfQSmcjoOOCwvlTH+jRuUS7c
aMWfsjJiAUmXp+506NjpMaTIKPMoXO0jtuIKPC4UZT8MuAPikvpz4UcF/PgSwo51
J+5j0fFAd2ThZRiFXjETDc8oQnoB980RKHxxVacL8LZszGqXBxn8Vlz9rbkTPhP5
V0HEzuP3em8LfL9UEMmtnLyeezGw1zhFTo/12RJY1sA=
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
iQy01Z+os3SSRRL+pwwNUKKpm/AB5W8XYPWzEQa5bn9VaQf3N+exalmyEKSBibKl
hQf1/kYc0jXG9XiWvPHrejXxU39NETRGeyqU6+9q4ozJLEFwSb5Y4t4QGMIBjnFb
o323YVD2MfNf5HCHz2j8SGoaJUWZmcJScmB36i2AVAA64SbjO/W67a/LmJ1BiQ3w
PYQjncn1oGC3DX8iqqZYhexyeJGvA3zIBDUbEkUX44uVW80P5r5kUBfMo2AowskQ
j7yIiASlBKud0tTV3umctFPtF4u/012kPFwoZ4xgK+UjiA0c/qAUknw25ZIg49DI
3V/4N0Ddh5cotP0reWzcqw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 624 )
`pragma protect data_block
d5zQ9F1e3F313yEB8wTNkpwlOt68zVvOu9NxLAiDaMxA6SA5b53K3m7RCqONRaYf
mUFoXDQto8W2D5qE/uaxb5uf7eON2JvWOWJMf9E6pslfP5XL4sDEpKqM6FNo/Aob
dvurEx6dzkJjTwlV64VlNfoi8Ve4N+c/Q0zcZbBlAVCswcMJDer6K58eCYpuGiXJ
Yu5NUeorwxSHym8bl3d8IKQ1ULDYFk8XQy7X7P2jGZ9roWiLkrB8zBktrxzwTx0U
wQaEBnOBWeJtox+pJ/j1ms4pFS8RCYTDoTeayofkcsugU33EwtP1Oy7oCSwhHIvA
Bf7Sqlh/vva2ZBRb6gUoQkRqwC9A83SLclwAWbxSzLtqPiXM+yyxBvo9L5RsOA3s
sVNf6mCv0pWkofovnO8pgm9Sd8Ax5D+QoWFeRvVsF6K5ikR6vRIZmJBqMGDN5rTV
LuHHGB74Xw1eRzF0fjKOgf4X8yVg2x4uzy8fg1XI5aUiJG3px0d6SchXJLrCgXTf
qnZwdBVWkfvWUPDriEGuo3Eflw6Bs4tHXd71nRTuASTMOYHqwtvMjfD6VUUN2OHS
7kGcn+kNuNHXsNzqpYzH2RDadwriZQ4l3W8y8g8V05046AqTGCr0Pc+yJDi1BtPh
nTRPoR0LfG6If9kW7tK6En++hM++WqCfcVR06+CyZUzIeTKtgEmn6JV8bwwTlX/z
jWlUPQqhUEgyXlEze/19EbltaBakDML/eZZouyaD34LUmE+uIHhaDFDTvkpOuE1R
SOjO6O4zKtWCSxZbC+MlO0lnyiNP1eaNRXVtTfYrmi1f8M/Pt43y6ewnHzOVcXC8
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LJYzhqpgWUDRLT7lO2tk7a+l1BP1IY0wZ6TkKylUIyezqD45dipPrMLpnjkEfODV
q7Rkl4A/yqzBZmdka7s9Vff/bVQ5g345nVLq3qarB/5wQxokx1Tqk4pJqpH5gey4
w4Bnp7So7+KuYJYvCUNx6XGfkI1/r7IJBWla4qI9HIumncMEOCji07N9AEBWJWxk
htXHPUujVvtlXl9GXQaLgl8mO98BJthL4ywtwQgEQe6t7fy2k7a9R71KzPuMbxvp
TGVngOKK4m4GsU/rmEIY3teDVefDlBBhOWIO2EgMedmanWa9BySgs9iIxD5sWAHt
Tp9l7S44lQQH9E3BlwU5vw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2592 )
`pragma protect data_block
nw+A9fNCvKHkweIiDVB6uuHdBn+8sSN2tHOwiNEV9uOzAJDS9cDRCuPVlYUdWFIG
5ewuiYEour3Tw/3IabwfxxbDqspLrxLqV5QFTGkynFBEwNvB7iWgfxdo1iM6d80Y
68B581IvAxT4UUaxRRmlVjf58JZUPyXRQchgRkBJmdlXJMo4cvml9KCi5yyktgE/
HjKuCynW2Q8GuZWMQhdSfbYudse388+8VC5HZZ7Bqv7efWBYJFVZ60I6oaFkbilD
YRvJVpvG8AIrzD7Eq2rY8cm7vmVpLG1gZ4w698LurO6mzj6NoU1waF/slo+W5Ipn
K9UIjlaB3iyYOIgPNPoJ6ib7cXJGpQZadSKVOIeBerVBTqvkYeGs4c3sRykG/WGi
vNHgTK4Evw9QHaPRMUzcLuZJCvtim6A5hRz0OfOno1gVEgvOOPpm6/6uki1ZTXla
vkmBVJQX16i8HdloLx5KeFYIcocmu5+7VjivlLp6ve5muiRDVY7lq+VwR1DKsglc
uLjVp7RXXb2edh/1SLiXAzJQ15fMFArCHRwuA15kxhW1sA7AiPWKTOb40HNCkYXj
2u+HlKnQXR2IxpKOVgRqyaGqZPUUC4+OsFNoqqMZVGvnMqjZ3D/0iUhIbHRIe93P
crZdFm5mEQJobx/PmsY2Y/sdUA4VrinoEBwumboHcRhMqXxqO3qv+Prbk+zoeLUs
a+zqcB90bEq/ruib4LRGpKdurPE36PqknxF2vxmCjdqT+ZVInwWHIpotSGnDCUae
/AZJvb0uWVjFqyRiaumazOP8Camii/Hvofi2YbByNNDeNTR4mJ4styE1LgWm3Di1
FFOVkNRTrwiXLep5Iromad5YQCcPr/eXDAdC0Dnbd+fSE34S8ZeUlDvMdTsXpDyT
Xab7gQ7ReUapy6KBsbOJEahUywrzAQd8BWqSP45LTePI37t4axunWdfkQAFbNpss
DLRyNnNU7L1ZGHFr8DCe1rcPPaeACef5uYbjTw9zioLlJC3Hjmu/CTu30eboDJ1b
/83CaT8+aao/57hi7SA1OZsHihfWQFg3iWOd0QXjiGOqFA4LiDNK/MQzquF71TWw
U0nd7/iY5965jZyt5DytzqxkJUAQLcpUCq/2YbfI4Wgb57Kt2d/8qQZ34j0TRxnN
j3KxhbNXcn9PAILbnXtDyraVB4B10tyaAeTwSaoCsnJdNMKGnyYz5YkglMvNRNwQ
CNO5+e96YshKuGQxypLTjdurlagkzz2cETV18M/P7XBIN6VV5qqaUQt1Ii5MpscV
XBu+cVxRxB1C+LnUtWkCZerLg22MsQJJz9PVHEnMN0pnobBfU9ypfNYSYTbMcWdb
lbq5fV46Lx3Tpni8HZzJo17n4Dol7wYdpT8ssi60K1MuRSyIc1nAUiwkrcmu/OCS
TpLUPbVebJjFRIi+EwIyVnF49gYThRn/AQz78kB6RtjktxkfVz5Pa2KSbEVu6IG5
H6J3+jX05iB3giIcb+vN8wglowVS6ApwgBXiSEQzROt3zufGcQHMpYjqoVpnzOVF
NElAV72+64TTsFWDWdbAQCnzFhpH/olWHWpL0HEGALRmmKym33gJqyiHelKlnI2Q
TTLGwo7GiDFnryzEtM2h+b5X3nBCCPvam5AnuKbRAzBCLygzXzl9x1ZByPXScb64
Z15g6ozaWHpUaekSEtfT6kbRS9EO92LKOq94d6GSxIyNFLEn0gvp+0BWHiBtU0M/
qBAEW5jeqBHPa9LIc+8MaTCtZHoDMW967yigMxVmjBuPnwlNGX1Vxxzdg1hwGJOQ
cjyNLFsfX4DnzFdqicmF9fLliJwdQ+Jqg5XVmrcokI6vzggc3BXetux4/8YRjgw7
xoWUC+BijcTJdEG2ydmR6d9QiuEEpSqevpFd8AN4ERq6znKNWbgAs4YiyhSLm8n2
Dh3PI3gun+X1zP/0lzJGRvl1g+PJ77ICiKpTXbVVwepTy3i/vd0nmg0JwEdZ+bo9
66VWVC2ENhctuJtMABbU9LvJC1dcRILD4Bqcr26sfLyp05Aj1y8uHQJJhI/SYeAn
4FHEx1AMnll7Ifho8dommAJj+zeELWNUJ3bpWk6rIYKz7TouiHAB5A6UO23kkZbP
T8J7gOh2PN/viWTAS8DbDv0ctOzi7sXm/tGia4neL/YYZxUwzmGszfBJ+GR8Ouui
6NOmLmhUUjqxTLdBOvkqfvmcB59BN6Dy0EsQDbQp59rB/o9k+VRH+pPNIF6mdmj1
YH0gUXt+Mo8Ewxk+oHh0HAFOzeed449+avb7mBG+Ii3NWvJl5jByQZ4Q4WUhZwkw
D175HmLMCi7nnAHOzBAENfYf8fnU+9THp8VYYW5SxvLKcWHPNxYgja3jV8sA3Y4+
JvNyZtzKvyzJKyxFn5vePmwLQvTw1KpfR4wyMe3F3kSIlK5bMd1xftPKExZ5a6eo
8FxBNa93KtbCDKiUaXnHUn4YjOWJegDUNjtpU9c6coFzW6mrG7oeyy0PyuVF0Ksz
73hfNVKa6dDsep0RUq6cfGKgklbjMZKGfixooURX6lqeLHfwbVKKwE6B94BrS5CI
LZyw3JNKNx1cC5ugyAKNwgyWqymbAKuTb3Z1a3PlhP0phVzOFmJKs/v93HAsSmnz
tCh5sn0y1ahkOV7iUVc+AfOnEHrADHcTVH1k0s/LyBVYw1AZai7htbK+cHh07/ny
JuUX31qfiWHpyStR0EMNA8M/7Wf0hG0zL8KZPB9cx67DVAGSHA0AaPp4+u9+kanD
kbnnL6XJp2qRH58iNsMrPlMX3DlAYzcfpPbhKRJIGi/Pqv2sTuPf2LvreOQzegtr
NC2yOnphopjyDw15w7e6kQkq00RBxBmgkSXtnyMVcW8CJnC35guanUj2CGbl7dBp
0VVAAgSwO9scWpQx0Vrlo+7N6tVtPBSidv7ecaY3gP2zjx2jx4MkMm7W/jYEk2Vt
UJuOHwCJQZ65oYA5IXzpAr/Rrv9Mh66sRJ1dMvT1kE+bV0I4tXOBSmicdxsextZq
NBvRe81y7/HhMHTZurXB8rdPQTJe4peKluhUcB+NWt5ozRjdMKKRqi6+/TUXGXsm
nHEVqwe4tZkUvsRS7xDaE8cYnMLykuQVB05UudxK7dm41C5Ru/bfI7Aclrb4YgPV
ePRusBhSaUpcX6pNQA4xmfBXCfAKqwIlkEexjAP/BPi+ZIqpFqSHioqnCKSYkWfn
XETniE9ofjV5Ydwrc4qLOGV+1cYqDzd4dXcm6Az5aL74a1fDew3ZpdbogfAuUfQq
ftlRqiWslQf6ZT/V8dzDy7p8r+iF3eXmkvF0cb6UgxsngdZmsZOekGxHDcKW2aFW
fow8nTTDXrFRdxfXq+TsY+iUqvqM+3qY+cjSQqtJ0Pi4q4lGPeU7OS0Zyg0z6BtE
p+B9MK56UiuZLp31P8mHlC9iPFrDgdLIjbW7dzFqjMnkQzOIFBkndAG8gukVYf8W
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UYQgD6BMBs3FymQwlW3gZGuxOnZ8ecCkrvquTd4taT9+NAMEfkT8PjOZveerZNwr
CjHUxnjKGd/1pE5FT9pr4F/r14jO2MEgkxJKvB0yefZZJmZBc5ka3tx9S28spMs4
MvisAK35rpXOKh5A7+9BxGqpC6QuL720uUG+P5IoLMkCblb7nFkHeMEtax0rZ5q4
f36Hx4VEjfzzY4JGOQDkhKSzW5JYtinHPU5f//FKAgbsimWTZvP48bEHPJN0bclf
j31Km8E/x5+R6vyohqeD4P0qct8jm2qtBgVhQR4McorEEkVWJsBM49zN7p2dO6Ln
DnmvvHppjd6jb7ScF8w9WA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8400 )
`pragma protect data_block
zZrMmJ4lG11hjgloV0Ars8dSS/k2FHQXvDW/MiW8RRzUQnwypeUL13oHfEHwcGEp
E+yWCZGyzEMGgxISTlc6GZdhfRjd+kvndgLFBmJe1ZVhgyV8kb1Qky8Pt9POMOKo
JItGxV5sRcP8HI9ezbEayE5Bb/G6B1K1PR8irZy/2JFuGZFULROb3ED7IWwtjHX9
6o5mjvDxHBmIEVGvpd7vQQFhDGxMLUqpjPFDFeKXqzhf92Vlp2ZnwYsKvEshtoog
V+Gricnf1Hl7jAdPDzhOcrSysrHmtC2sokV2Qg/tED2PSBHya5qVehDjx3itl40h
Ofr5I5GqzgswY7pwiQXlARF1wu0yisRf7QRnqNvSozZrN4WiWGCNM0xYOX7hOCJt
MusHv1rUBrCOBaZQqCp1fyCh00FDPNBxB4LouoldGZc/9waRUjH/NwfLTuaU+xk1
9bqYz5K9zLbxd2ImGSoPEbffmuZEthVx2ppp/Kvh9t2wpSNEt8knm5MAmos5KYB/
295Gn6clccsvKBL9/VYaQ5yq6/rrY4O4W0eWTUAppKEU5lKs/IiF7Cn1g7xYC6hE
C1YNaoScLGP0BYbv/vTQDy7RcjmpVyV0Njo26bCPv4veDxd79SXPlHi0yEzt1GW2
udqqlWnoywncL/6dAnn1TpvAcmjqaT4w8RWDP8hqmLA+SwGGhHqGRMnH49iHc+8U
56Brp6lp/+Fci8HNUioFHam1HGHHFpZS54VGDT51hnWGfW5D1e7UYqiuEzj+xJOt
PfFKiEif+NclaDWrdhJAFXiue8alUebHb7CAVaQ31WvvnASAmCr+pbcABos0ZPzi
pKFBqwKknK5bhKD6UeMNVIr76odLdjsyGRw9FAMH4D3AMrQOD3xQxHp3xqCWm8w2
2BNHmvfW1db9Lkb/+Yb9y7G54SpRwSAzE7hfOsrNEU1nXZfXyauSwZyHZ7yug7xt
F2YsTGqfSt3YeriN4jvWrBsZbGu32FBR6B27YOEzZBxmMzytIMj24UjFMKrmLJVi
51i4LT7ob67CdB6x9qn3y9E/4OngJgAG/IuMP4iU/yzbRv+gwJo4Kitiw9t+s7oy
9JBHiUE+q7WophxqQzuKEmpO8bDRT/RHQCEiHb4TvAkevK4jPM4gdMCsp3SveGHn
yDD4uCEymTYp47HUfVE91Jq2tV4XiTw3KWuy1xUARdQ3PlYG11uSgcttJhgx/9/Q
M1uzH1tIHAnZoBAv53XUhsTbtvgEEGd31tV3z0R2yWahRThkX1ajsZxYAPz1MlAw
4L5S9KRq6baegRz9p23Rgu5DPkA0BPunUsoQkWvCx+JUg7EF3yvYecQD6o4UTNFW
Xs2Hs63g4iwonSrGlJhyHSvOIIPmIjOE2Lp8El4p/B5/2kWC+Lou+Arh5znGPepk
3g6DnbduirTDvN0TmcDO72Hrrrp68LVnFKdbUw0vhLEhgiqq4x9Dc3ZPRDDY/wUK
Ucy0zNl8CilLxXPGtluOX0ysOSoz1IsisgviSnDlbRRNJkuRI/IayGQYGoG8Dsw9
xiJ2ESs84VYdZdsEdvIGy2CyIJMBXOdeCNkQtiATQ3NDyuUpGuD9NCL4RnVni+0h
RRC1k15ePUs1ko39FK3N/PwerMDvEFqiYKoRXVTGLmtRwrNvR1NuTxLM2RoLzgr1
z534XIGMVuwQq1HyDxUubr84Kk7mDR/HvotGshmC5ljw2PxfNzRmZTiYIp/59iSv
i2RO2R0OHkGd6nPPw9iW6IY+ugXnQATKCYOuVQqLBk6Rcz/3kOMXB9Fa7yZ/R/Ix
bKDiQpMP4aMPBKXfS9V4GB14N7MNgStM4ds7XXBR7tSPhfzobGCqC/Hfu1DuHGj/
qw0P4nC/4vIxHR1XP7FKnVWZXTzZ1PtujYimrzJ60Ta92hmOB00xyjhIgD+e4m7K
d3YE/PEPgQYzgvn/uzsspbRf1rNa3u4h+rMmkOVGqIef7dD7NyAQ4dW5uhRq5FLi
Dn7YuFMGr/AcAoCHmoVOQJXRS2yOHtfgExDgiIwOAK5MLWEUYvW1agMpe4EZlNbT
/637079gxr3Vq7WkXris84/SzxLxFzr0eTU1n3CSWEZpbBrKknGB8kOLCZrLKpqY
l0SAp7HW1YDMbs/acfElgr1IZBps86WJiAwTd3OLo3VahtHyN2Bq0v5B3h9ZtII/
8MwFLygurv3eRoUZTxng3GYPQH4HO9zFsfa7eN6wiyGi0hE0UuBYDrbxoG+uGh8v
H8+lFaoEYzsHuJ9j6H5e03H97CJj2t/bKU19xCOZLMd8Fti6H72bbKEnfJlnrWEU
HnPh+SEd1Kl1xdi/1LUrjamJswaHKr7AlpzVhEr6Uk/AEpj5EaQ+w7ZIhOdjvx/x
eHZqyA5EcMbBk+TIvF91nCDjmQXCQBq8WHzhkBJGFy0Ii965T5H1ZHEEVMQS7jDd
Ax19w83hqxxJEMfgRbJOoCaMSM5toeIRsgaSAaSPJr1OO9sOmEkXJqGDfBqXvFcs
+kMyBREgu4PJPsVECwO9mDRzYxWlZhMZbiNngHykAS67ETDCb9oTOyH/hZxW0USO
a15mVGKXEcp46k96lGsSmFkZzYsy1TJjjHrh2QPyL0VaLhhba6DQTJSmJNW2sRDy
bFmRBnIZXcubdZspW97rCasODBxyk9sPGDDjvKSjcizpjc7pmfhQgB4WXI1BMvZ4
1MOUPJPvEjszuVDbkznGP09Sacj3+8vXAEjbHaqvWNjDKVf9C443/8RtVTdApFqE
pb7t49UHePaHvIwvMp9eFD+J9XPIUNKQLS8pOvuXg1NhPq+4cVO5hrml3HhueVDP
s52vPb2XQP3vQFp07erCWNMd1/iffCJzHOMSlVqNhRqXcZbBPxlBhBhq6UTOADz0
AOD/c0Oh2KnBvH4HaXzf9blLIxij0JkylZOmXjDF5fH8PB8rDusdGfGmlfvTJD5Z
zud3ttJpw7djCZr4i0KaDThiVm9N8FepN1T6kxs+0z0qeouMuIUOSv8a6DUoToka
I9YsgbgWg3U7KP2Xf2oa6ki2tRtoZZfUfN8iPRiVeL9PZsIXix91X4KdY4mwGXGT
wi5nuScxVvXZlpqqzFQa0mvjwPbVkQZYrL/YI7Zw5CfuqnsAp5rVd+KS7DErGYtf
p/YR8vmNH6NuWJHeo0Tqa29ajWj5a0VGMhGK2ytzO0cgC88YGMV5bUW8SBQAfz35
VUIyfbRkrr5U7HlOTd9IBU6qO9WJ3Tq89pmpe4T80x6eeK44Vs+7RQ++V2Agrm+x
v0mQvjFH/VLydK8Zyrzx5M9zD2fu82ol7FxhtlOQhEsQbVGyDujAMhcmoTPDTspe
mV8mvjuHJob7mFuB4nirODeVhoz1axDRD0fe/eJi+zEJrp8qAPqRCQpGdDkMSkkI
w5ITm8BUbw+kO1J7niXqlF6FtDFnM/hU7xWwSDWAouB+RbdLAH8EL5pa/81DDoC/
0HD9gqWfhDE5clal0dF1Rs6gpvIAlwjTDENus7/dgbIBzwFNlnC5cziZJ0XvxXZN
h9EXXfdZF0sPuRcd98mDjJdTvCNNAeX2q4rq2HgFCr+fpvsbzB6twZidp0op12MJ
EfmZTPVT26IwKXt9YKiXgqF/NNkAMVpmmdtjcRTomhxAnmX+hUkXkqTQfRScvz6b
Z8ZAVECJKqGEc0hXwS3GO1wWLMKGcuvxpgWno2AZbUtHfqvjAO97ciwfJWU4QZCb
inGx0k0mQMQo5CPe6bpu+B4D3woMKb9Q9NZVC6f41ESqGKqB5DdtRxhT8FHwtY3u
QD1kQnMA1MpAXaSHoR4KrlTyBnIdJGya45leqW+UpXjUpF81YB1hMOiLN7T512Db
roPGJMgOuRKRqiv+21IAbPkzVa4Ve32+bo7mfxmb0lfnxwGC3LCYKOt7pCOhibiZ
ZQdlJlmzyeWlVSieyy9fWHdV483UcjH4Zdz+CzdPHZU/mF+E7yDFQPD52IMrlpzS
I19bItPDAIcKuAEziD82gUjFnpJcKChZd1rJR83Iy40Q3sRzR6cYdjrsdY2Ak9AL
6RJISWHWItg3yjDj5nOyxF5OGkrqYYw5OigFK0bNYrZe1o94xKytj2+OqBwYandE
1TEVe0VTmI/5n+zoE7+mjcS2K90pA+pS0BhTQ2YbmKWotgSGWhU68apuSHIggXZR
IjYBQGEp2TWdrskt3jyC6IuMJoDf3Z1+1uEQ3GBv05FhcGMa0QD2M/ouwrWfd3mM
uLzSgyQ1lLk0x/BtmzKtiRZAVauOwRcM1PVutp+ZVfjJMQq8OthsvsqWNOoKiiAa
eyDPqZkTJ0sVi4JhTuJCbvZ0ZjRQsayaI6GUpSIzWcwscS3OWxjdRfJWm2eCq466
lnt2JwVRg7wUm5Uxq/+7/mH1ZylDBx0s7cTtRO5wljmc0Z55UFDMwZZnf+23rdSs
Kj5MuCQaq2Tjj1Tk9F+9Iqy/0IkLD5W7lcZKdpPwdF9g5R4qji1KBOMQ5jMocjUs
PycSx7mYcdUw8BF1fYiPHayI2FvM/0Kvh2WHLdcAleNNcQ4ig/+dkBLAfZlGouvt
mF6+W1eVlElr5VbunHRzwbYhf5KcaP70ZF/35CYZCFPWDJsbRB9eRH5gDAMe2For
DBzZ1D0TTDkbgIljLjJC9wt43C7PeX2w0HDKqoabSh3T1yJ/vX4FjStJCIbbpnZ7
b9OZgr02JRtWNIKk135MIUOd4uHb8A85ZvLXA93FxShN2bx9LCpSrin6iroGqasL
5l6TA0aDw0FIasl5jF8Su6dAcRco/QjEV+BStYeKN+P0QYhjzidkh4RAlH20aNsi
EUh5ik2mf8o0hA2fy+uDPSC4DhCbgORYMgnw9xXeVVHFLKl53giE8fjnJ4yEauXd
YS66eEqmpwnTsGh9PxkdYT4ELsa1E0hnhV/zgRj84HLi/97W500AGkSEgc4CDEu8
O0dRG6lgQIUD2gmttpTL9p65hsUA6o7/mmyHNyeh+tBkUQBOtx/4obwyjDD2LABP
gzv5Klwac6idnW2x0vVRdyxzY5W/HaNNDz6zIO45i+q6YCmXA+vonoRKngve7WqE
NnqTq8zTiTbJj3p4ruDw1ikZX+ixeqGnes7XXBrtyaK7y1Jo5tzkouP2w/lSvsc6
aiNEBc1H38gTlbYRWwQifH7E85rvEFtZhayXwT4J8SMm9OEW7ZhjpXusFXaV7c8h
buHeoJ8chB/z3Lzm0LRxvotZOBUZ90f4ucOHUkmbYDzGqJjWmR1L6139bd8h/Cge
iRYZx6X8ZrgHNLnk8MR1hc9SQfm3m1zsbtkfcxW+mofBv5pbiH09m9qHXrlkPWU4
B7nth4s8Sv++UFpm69LznSV3kg7IGqv0YiSYsO4+EMiidztO/hKPEA+2EjkxY/rC
tn61ccGPo/B//cRcddPMU2F3BaNG+x0au7F6YYizVGIiGe7VASuafo2Wp4NQrJhT
xQcSTciIHc/PnYpogJ36lOcTdoXuOP4faQKkNzo4dA4gE4INdRZEUc8rqZiKrZ6A
McdGKERGq5363SLybY3z7aEu8FX0HXSediNfSLtkRa0YBq3ob8gPcKNH8ZjXM0+c
uqKFOgWQDLoZyBppUGDZ1uwnZa12urovVuwaklk51coxyAzc2msPuZNGP5XxkPaL
FajnxOxN4Eb1/rq653nAUHRNLlCX4DzkHLUNmSXM/aN8MU2QAz25Pa+sC1X+K3Um
V4ohpSibBPDNkFxiUqNPRf9XEwVcDHiT0cgrhtWARhG2w3X7yEkW6YcE/1jaEb/Y
6bVJDunsBykflqvq8tuW4yO3An4eaHS7DVP0YswpzpZoC9Embc6qlx0Vd3n3grck
DD75GVfiVBXq/BMxTuSvowC2ZsqbZDhxL7uYYkzMW0Ue2IMBC58zuuP/4lTCpduH
jbx/vabIrq4q6r4maUoypblwmOxo8Z1CV7c41SkgiYiQflKQhjzAYh9VnvNTb5nT
60nVnTEcBwpvAeAIjMipQ2x/pOy+Nf3/12PfZTN79OYhu2HB2j+7auoKpv4S7bFA
X6K+IZQ8zz0yldWAy/zhoE+WxVNhQ4WtzsNWrrgA3im8JFCXa7YaF3sqoHVBNOqf
+jraaEpGLqALgnh2egcbFb17ny75ZeX42jWGC/fxBri610g4RbZNE5Pa6mLGpHFR
eKUns61ymmwPGT/P6F2xGyNINdr9FrSVdpVMns5OvJxBZiiZAFAyaSdL9DsqwYqn
FSfznDw/pZdjztgNuTRemMuXF1eg9GINMaAq8BB4yOgA5FB6MO6eFIL7sPh1fQvZ
SdcnvqErpqbMilGFHfO8uJRYIGdfnLNrJOML4/NNaI1LZy/Lsrgg+5I35SXyfj8g
RU4ii6ZW6VICp+nrNLtZfD0nvof6iv3MQqfVgzsRwcPJEILX/A2UZarF32qOgD/s
1WJxdBFotp4d+STA3wsd47ywOV5COClhxXBQm3UeMrBOxxkWbG1MmC81pYFhIbhv
0We47m0WTfufn3HKvm6F3wNexmSgB2o4FEdTAFWEKqkuKis7B2N60HNg61tL2SvY
AnhZMIsiucuvr5ONOydfpayOcHglB/qgmNLw634HmObvhEuXtn75kuQWTFcpPDiE
NhqXFsh4Wacm0Sep36OXlbYfR5Ql/P8vw6yi/Q7FLl4ydn4ummn4VLyXZ6FTnjDf
A6SiwVWrKQfub5BfrCiOWbIoE76S4XpDZpoyI4cn99B08J4ECIf+Q/Og+dgnocMM
lvmI7wS4zVVqSFTd8xhZAOyudwrYJJzIS9phHo6PqDSLEyHs8JClcyFfG/oKjmjo
JoefD8ScSZUracBNytKbpkcwQkmYaNqT9V0Vp2Z/Q+b77Uk7xS7BIvwpUBBp6aiA
ef7ZP8G0W/S2jjJr++JWqzy8Wr6czdn/Gl04nuTaPnvSZq5Jc6YGeZcB5kb8fovL
Z9iF4QqOwHfIBiIp6+3Zm1BNJ2OAk9CmMAqbZWV5oqAGRyWNTOm8ySphMg2EEXLi
cvvJD9QLmD7CQPsRTsIf7DczXRHJFQ7bcoK/IpFQodglhXrABl+1BpCVE/mAjhwO
Xe3hWc7bi+yypypB8i2gpMrLn7EAX1hTsV5hOh8hwB1z6tPl4rXGRxEHGwUcJB6W
rJr81M+5X6Vk/TBREMGN2hNk1z6kpkccXthBXi5Ujego07QymO25WhrbhY8Qz3Kn
kLJh4f22tFvIWVbdnKQzCL67LQqDeNc+ZzMG/rEV8QkglYmTqkdo9OKJStCsTWoe
sKwMfe1iomBamXlT8f1hfAAy3r6pBy5nziCHXF5YeLuWEhNqm3fcZeyB3qDnVQWT
c8ZeLmq4DUtGIUodAMPIuh/Sbd0R+pClh7LJt9NEsrNiOUz/Hj/W/g6BihMNyBKz
3H23/4VL/DzNr24MKuYl0JR1Udl1eCvMFKaUCavk/5CG6r6v1heHwU4xkG2lHHel
EiA++bIbItb7wTLKWUDx8Uo5I5zj7FKB6rUM3gyy/R9KMMVPm2YfU22edoNAuv58
hE6Ob2SleoFzYgHy+vaOw9/SbXNbPCLC4rhKF61d/WbevAeRYfKNJyfR47SWq1/Q
QdZAK6yx4vpu7cyCql8tarvJvHqm8kTEx986w0m/TI6TTAllX02amTnDm8RgYUaz
DY68gJx0aBB1XbHm+fUQefiDxfH7GE+vOXqeC2v0h1PFvUOek2OmxoeCF4/k1x1L
0Hncy+Xvo4cEBcDvalRebR7G3EwIIZczOeoZENww4/uvPxg4hniPB4ras/v2s6B+
/Uf6y566pwRQVmexItSBz4APV9QWSPds5YcvKEFv+DyRA7gePWpC4MwzQZUnUXwj
fJaiZlKVb/ZFSmPR/JvcvbiEIdc1Pf3L9gxUyTee2cWXCfxVebSTEWiSnd8D8Ata
J/fhBRTqPuVAoHyKTHsu5980FJszShugkrA+obtviyxhDgKRPqC0AgY58dOupNpr
JgerXptRm5lRctxOjKmEVZe4Vnq0lC/zJYAXCVk5m/KGw82fSGt9kNsjV0frc7Ww
q9LvJCEZHbc/xmYx1AuMj7fCeNkEBTGAHD7ipnJd1oo52HJb22/TDklBmX8bAdPi
LHMVqyFFAjQTxmhgHvl8PovvdNSabfW95uaCIn7K7NX5KkSUfFpYDywPmSUeUtyo
dJSdodfRmm12fzp7lO4rhAnZU6n7UGwDKp7LRJO8XYygU8c8+2p2R6+RfVlSAt9/
iPYhi4hAcKBWzunLuzonyiozry88DwNXuCWwyBIV8ot9Jy5cFPGp+aAtxgusAmGn
Ck0zgG7DOhGlnFisWb/OVvwSMvtqga7v0Y4wz3zGE4cFUJpDCq3VIB+4mJev2tfK
eBOL+VMkTk6jnsnEmjbCHBVBqhWMCL0x8Tnqffzah8GO472tCNAfXoq9NM+yzGkR
zBRm2/HgiZ1sNaZPboSsmEBd9Gf/sKzcPqw72tdJodSmndQ8OXTCawyJ7X7BXUHy
tQR7DbDOQ9L6gR8lEot7z4ydrwrrDAjsvZM2e1ZaIsOB1rnLpmnhTaC6YEBr7jpM
ZZe1gLcwcQpnwwhoMkLxaJq+sVXxVnBUo7tgrkUYjrG3rPG8xhhQQnGU5AWucxYo
rOnNdlgVL2+7Q9+HF4lsg/267PfrKuv4A5dpCdBA5Flx7mywcXYJd7FjdevcTsWS
hPLOX7ga4eLAe39vsLt20cebTZdC62zm1QwC3bo1Os9BHHiyyLFMZdE9KMgfXq13
xYIzUhwWA5VbUSmmVEsPh9UDhz8mSCorFGf014j/h0yqmU/TsXjxtjfAjbOHvI6i
0a+TKXveZsMVKnccBlttW+9tRJ9JPsX2qyoxMYEibwSR4mL5EtVs44p70Sp2ksBa
uvNUGhnQ8qwCF0pSFVJh9OzLqmPQp1wKckBzvFkL8U74ow3dCNAaH12UADAPfKVy
Rb6FLja8lOWQGt9AGZv263IM7gDB8Dvvh9WJmlItxxWFbLv4sfpJQu13+KUf13SM
H0aEm1PGxV4qOoXFq1pqFv9/w8psVYMo6QJq2555bzjiyy/zYa/OF5s1Ca4/jRJZ
NYfGvgqG2reZL+Op4bTIAmKYvhr3ziKKFf6begPhD0vr7iN9MACQfNakpMDApZcT
DpmTAUijC3vQUMs2oxpPW4nE1vgAri/8eDlxT8eIcYK66n6TGnsqIsgIxN3YWUhi
q6zRi2MiOW0+DXRj1UsbYXK3dcYURsbGFt8RIFmxrvpmLiaJi7YHHTMSK0JJxyge
Ipxo5ti6XQ9cwL4+giX9S3bsHeqJwhQ0c8XKk5ujj5VTkZmsLNh6i/A8hh1tXW2j
k5BrjKXVx0EusddJ90Qy2nlUjtFNmnACHwUTx/yr0naVnQvJQzEREcBz9htlEJsQ
JRHgz1VymxwzPBh6tE5Bp0v+nw5jZaf75asqu09Jjd+L2McvXBxvSZEiFX4gstCs
1fo7FWTxCqrYWDDtKxAv4BpOrAoA8GuZA3O7KY5gLwiTZBVsAycZlBuDb1d6anej
qRv7HC6wNlP3oZ4Bp19sWY0JzDHxan6ghGnorqt8iXPBe6l8d3C2OLRJiuRgbPwD
5ZXSKYVsVXofj19XOXvDwU96SQo6coakEI6ERIkAIbyIC2k3AyqBwATOcwJUf+UB
zEqgiySj2W+lqQ7ODLMFItSfLdFo2KREIfR1iyD2YdXAFeV4dQnXviTNccOBJx6v
L2EGzs7s7nerwgbCljuDfwepPBZeKHRuthQWmKalMqFgQySmrP1NEBN57ICpRKgB
6t7VeB8XPKdPRHlkqyq5labfvoamfcBQQb1+Pd5PwntstCkR+FnV8dvi9V4EtbvA
NRTM4sgbqi4Yyrx/Cx1ZaIhoGOB6/RweScaPWrcNi8KHp2TmNQWV1eoiNXDlyGUt
6WpLEvKOMW+M79BeHOKj/dplriH3qk2dMBLKul4Oza4AgzKmDoQkRNyph9vQrnvp
bS8zpB0MrSNKOD/eCxrZTdiJ2E52nIkXysH3fnPWLR0HTj9SPhdyo/occBgZJzuD
mG0MoqFq0rpdVmRGcYkgsbFpRsRPamtWyK6D1EAp6+g6eZyGq+glkpQ3954I2e79
/qI/PBscoRoG9rJ+cyCtHeusTxWFCEtg2MNpqDFFFSnM/inUWsQiLCzI2hpF5fJi
bjxYu/YyRIPD0RI2bSMLJGyRAhdzptXhizVHImeLb6nsnQReAZJJU0EajhbSoJ+l
iojCqnG4BtMYZdPvQjpjtBBWO1X9wHZxLkHGMLwowM8QLFgo6Sd5rMpN/CzfFa6s
dvnojODmXMBH/30nDwYZ3hX4NBJYdZPari7H2TOkVu9zMI9FsY0YMg/eFrCNBf5h
EIzu/qGln0vZZc/L0czOwRlx0ksYQlPOQXIwWRkNEMTfp/JXjPvsMPyYPYY2/i26
+c5bapJmKSFn+XxiwTrd5koKLm/RXQu8HytWC9y5lVVBX9wlboGgRKI2j9swG0Vn
7heKwyJiFUVWh4cepS+Hq4iIA+iKq3LrHP5Fn9UaoL8sEB99j6S2tDiJ7TNSW/zM
9RQICSEsOEdBX78Gp4bfNXlSAvB8gmLARKSGB/9KWjMRvWNSd36fRImNg16VmjH2
0VXBKr9wGzf5iqe29GECIJMPY18cUJSi4KLzXNf6VCLheUw1dK7OtbSnPRqm3O3+
jRW2wO5ZgGWsoXaQI5tLNuINtujYLGMX+5NVYWa9u9LQHZCZwMP5dJlTrugLMXgJ
8/5W/P1zs1aKNxiUHXq3A1fHVmSEF+YCPWsY9a4M/KWcRLxwSty16IzcWP6aYGsK
Ipw+Nr43G77eC4wtqLUZWgbRUzp5GjI3tIZE8aFxplsSlGM5UnXeo4c/EyAg0WIo
UsRH1oVLgmv2nNwpdCfkfXSwXixc9KprLbV3/KpZTVw5TlavwDtQoC3K/nhjmgxu
PygBYQABIXZ92tWP+w2iK08/F4n9kSaK3PbX8UFCRYbkEDZrVuIBW4tpqDiY76KO
9nTGWQWZpuJCMft2WDyxjlO3+xJrSLF+ExlddBfv7PtEfL0OLIA50T0Ir9O9t9DH
cwZUB4KyRuLLoJAI9Rrjibmm7BOCRMjaAA6c9ihuOyWjgeabuzsB0cOCvoK6PWyb
rbIsP3bNSSqd81+jX3Le7w6iHkyw1J4HhywqQal0dwfZhUu1q9oZLqCJv9M3i/hr
XuCZzFd+pGiwCUYvi+xt6gtbMtR5VQIbOxtNXnV6jen6/qbailEgjtwWT7xHvuiW
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cWFyyZmF5qOu8y6G7qfgo42s7sZxFdX3dJ7CSbteuXPI5AWo9ixDBul3XLYYziYq
CwHHOPl5rnlG6kS5L0KTTOthyhcQZCiGLnHIvM4mDTKPa0SFQTc/795RryYGfpIf
c1Qr3yZu9bK4029l+xVM+CXQOeno8etl9HkMQZAdBC5PWfcdYmakni5OqL/ebWfh
/RVEdsv3fUEfs3cUL7DT4lQEG/FFvc0Ai35fpFLXvD3/l2cYa8oVUXH1LZwtANy6
LqFuUwjWhw14vPOvwmhSYtpg+fCMRsgXwp+N3wq1WxE4KBSChntW1xSGWjoSIL7t
/8fZ6ZqR7tQidWHILaFjwA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2544 )
`pragma protect data_block
Y5FUR78tdI5zYCUwoG8Kj8hwIryRhYluqGo5WXUV4d+MNXRypANCLB0vw59SetY2
5o9mSIEMoOiOO3upCl3AL1f9URUVJxeCjMM9mcNyNpoRMdIIAyJaZnlk3jDnFD7q
qAwQxQDTMosuzqD3xGJSnbGvliPo1S11lm3LJVlIVWa6Qd+GCE4GmDghm/sZK90Y
wxZlNhslZwkHd00Ho3o/CNvaq6b793SxVcS5TiHukqvhjiB7kRMnkJyfl41lOG86
vkjyHjjKOTQ+6UZddD2FqTOoE3F1QlTl0xlAgzTY7nI2Ym4HR5MkRPiqUwI5vBlJ
jjLZikTu97mr4/Cc77sAWiCjPd5RFl7rKT4W6KlXZGDXo0oReTt6K0ktTK02d7nB
9PawaI+1H/OVNTiVF7kIKMXpENFtm9dEB+NGfv1A2OlnSj13OCS5K+iVzpD/ge/S
fbGX2573uefY1B13dpR1izsjKVPjSyviRB1e0yh6pEkdpxwJpEj2d1SBGPGGp9Ib
1Mw2ROhsev0wvErgGEslg+6hUVBjDohok5QTd9Yin5fG/L6NsA6sNBbN0GePuEcS
9htESU60dlDwHy5KCccAA0MSsjb6NsACcXRPuwfuiou73NWkGQ3kyoADBk/cZVPJ
Wz2haEOefIq2zLknGLM+k+8uA6ErEEmtdxxfoUqazLc2p/s3PSz7tJpCRe5cQptG
x5sSBY1dwenaENkrfu2K5iGA4aEGP4BuceQ1aBWHwq430Hsh8dY1vWUVwgdXrMgV
jyxj5TJCnaDrT2o8LeNrWgT8+nUhQwZA+xntuwkLPSzpNkONEbfdjoYoMXK2yxlE
aEwXEe4xKDgesQ7zKwtRQlWf0Yk84Kyc7ZjDxr9QJ/eODPUEA9uN2G14grgVyafX
u/+fBFQW8Cf2hemZ0E9Jc0w//E/JYrUG7TtmPt89I4RaAZGy3DCKgOssytl+tJFy
Zx8XvzrJKYXheXzgseDjmHk7MN537oVaLk/Vsmu6yEVvb9fWRYhzvtGoR/1VnAW6
nsBdU3IL1S08Rhu4qkYikTgUkYHGgIwvHgSUrw4Yur96ewRMmPAGNJxC264QSpRG
r+yDUM4G8cx4tdDuBdlroVcSpm2PpqfCuZjHDTgwRaOUlhzvyxsftFdhPKZi0Xs6
O9u5EFVdNCq37tfqt9X374uELlrcXgckehUjfD0WwawkWWANj+inj9ho8g+fUD48
vi9D7Nl6eWqptESioHwoQ34JVqiimsia8JqcdfIyuIcpgryOiEPc2IiU4agajbcd
yitrrCzYKHIjavyfLsxf6eM3b/Q+Ug5SgIYD+XqDCK8V4N+uXc4mrK7EKnWKTJqA
GOkfPgc9cklTuKxsIniyFiwBGrRaXcq0mNxx2SYDsXMXWn1Pw3a7SXnTRZhlL7Xg
IrxmGQyF6MIpnroZF1w25PTibxzWzqthEchcY/h0p83OEvMaIlTvZ28qiAKx4l4O
kmFiZXXVOfTySrcTNNhpc6ovMvqIXiGtHWd+HsJZLmcnH0wQOQXofbYeX4T6Jxpy
p7boj9qpR0SLGZ/zEPFXGIWBUbJjZEiwR6FYWl08M3aKa3O15GNFnTOB7By2kxDq
Uy4GGkFMU1GtjZ1XODZ1xaVnOx+nngHjtqfZaZ2SmJf7aMen33ACbxYFJRoiEktj
FaRU2uL2HwJBqZt/kEnL9nJ5LVDhgkKWNEanSE8M6DZBPz0YsoHCdH+pNGvzJVnM
r95+JDQLQYOeH9T4POkJI0mSln/J0s06l/DFKOuE3kL+7Ixjl8Gli9Z1rtPftNcU
XmTKtfxr6U38KEIAmuPbZ7V4ihfgccZj9GKSB7yWQHYI5Ml08vJXqRQdz+tl2WTe
bwNadWEaOjCQA5Go2k56y7BziVntlGVzj6M4f9x7/foiGqZKQ8uJe7zN2yKLPs9C
W9yaPrXT2pSFALuERSkZViODk7jvMscrnah1BQKKEh/Rg0DeR4HfDKrybDC3AkiG
7G++50SKL73lbeC0aNi/LirqtbcDDpyLAeEZWKuljzaufwg/iw6aE7yu3YSa+RfJ
j2PjCkZtTF9IG9vBQLyjRsOhuXdjiuR6+SXMcsIoKj/ZbU9RuT1Wvr49L3ddwr+y
/iGgtu1z3fIpEeF8p4cfsOSbEj8CAdU6M15UEfWQtyR3tlxAA5hvU60upn2ePm0b
MGmkWdrYmCQAYLkLA5ruQmFD4UgGFSomX7upPhgBPT4buNnKiutE4KwhlTQ+6Tux
45gt9tSHaGa7cKU0OeTqnteJcsK192MElbSrgIK72CTk3OMGWtFCioVYfbCKeEA1
fcp6GyDGUt+dwgloUr4N20i4U6drNCCwqDDobsxkGktVuNDUGbjZB2wECXSbj1zz
QHL3kiJd3H5GMzBQ3eKF+iGdziMRCpSPKuL7ji14QOSX4ZedfcStdtTFGBis5iKF
V1mu+tfpQGEooYTA74k+o1H/WcKl9BAU1a5yKXkHn9TOd/GuUVwnmblAdy8k5fcE
63MpOfhaMmq6zV2pOqo2VkwiHQtz9XFRRNZXAFYhR4WCb91V/dcqJWWn1Pq2HXk8
9CeLFHDsSdAuYtovA9ZkBzG8uyPSgB4XEsq593qYQkpCLZYf5OhmvZsoCH7jKGta
OBR9J0pjh05QbBCGwJRDgFKrL5NwOzVcIXJr9uzlALvkDt9dS4vanuzvvnajCYVI
laobJwPEPtzqQs4+zulxUQjuBi8PteuSJzLbi7/I+i9RGZ2MDtLq4iVtcQw8p3Iv
fDolVKyHFMaJ4S725yNz0Q/9waUNH1nZkF0JW3qt2x6iLXULLNBmHeMNuB1sXRcn
MUZKzdbPVZ1UqG/HAwA1IyMkTRv2qlCSqfdGzzx9KarsCvQnpL1OZyT4nQbOpXIp
2fACMfifIXSK27zHok6cHDoHr5EESGMJ3cXPRHqWmCRUqcRUo+HJkhbgiYXPxxqD
S23Eq0sMNyudLADAEIlsX1kjR4V5mLgaxlmJhZQ7Deie+1M0/sR9/h0XCfTcgDph
BBOw8WVY/EcqkVddn5KQQAacuNwaOIpOHDv/JWN6OhBLgTRSI8YTt+Iw3qGcX2Xq
bj/SonOa0mcxnzSYPyZSRjeb07LhsXPnEeN/c+XwRmjGTukGlb7u9Thw59TloX3S
9hg4oKk00pOeLhrNJXMknOaebyjqxtt0AH28CTTqK6z7VTAJaMHw0YOgAxzd0PEp
knYmwRz+fCV87+c3gcYnW6iun5j4ZPixKPLZJgiaT9YMEhjcZPq1FvH7TQxV8KH+
3Y+EJfvGZm+/J3YgY454fPjYMVN2GMq/OQO3uleF9X7yAL4a75ytoWqoWEk0Qcfi
7C49p3F6vNoq00APKGt8Rgoz8jexhqwJHpsGCdyCru1NdB6aw4GRvXr9qefqtbQ7
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UNjeMtfNgkqeXI/CSmZBmsT8LSlVaOoBc2nwOXhfifjXa51tBXY69XHeT8cOVxMw
2MJ4HWrugtPi+sveHyOE/Pc7OdrNdolR/JFIDD8RZsF24v+ecsUlX4tzv2eq8DYw
jdUtw2wnr5WcGFxiK39GCeEqkTKSbRlYH0AIq+QvFjDjU9zh6OyrnaLeNd47WN/W
wQrgYZ1KG2PrFazBdr3JZgfAO7hX55fShHQ+//YXjnm0lssXNro8fGF/fYwB8cSv
QN1VbXD69g1/CfMWP2gmpYJOjwOmClOXr3h8dSF60UGRrlA7BtwVW80Dkz4hZUZQ
GztSA8gDCpSXc+rHZvxe8Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8432 )
`pragma protect data_block
oMuX05UW2fI7yOyoJ6gGrvostvQyZnZJOqjyx87GepAl/C9dLqihsgpaNLulSA5u
vN4qFpIjhWXN/NGvSCHnJMmOaXKCnYuArlD1cT8wIWIo8MPBDaFOGltWG4MeIU6Z
AzA1TXOTV5omEPLeA5MMDWwqaTP4VY/kvkYIRY75Ql+fa/rbZFIBkFvHRSFK7R11
POwxxZDRarQoxICKtMWBcgVYhcBJHcT17RrB0uNV+z2h1Zsc9XB6Y4gFF112DGsR
xONUI3/KOyOGdDdheHJLNi30NuiLg7+r8ITpAgNwME9w8ix+gpfgqT6EMscdpF7a
RPUVIteZrW7HzBrkyTVwcAwGaYLfphWIqpHT7uO6QgFk/QUrPdKicPrfzNB/NJA/
ecIDE+BOHI6qaqRGJ2TNdahupL+YQYZ7sHm26oD7c/KSY+CXhkATDm3nBNebliyR
klYKX7Y6TJGNqw4g9sizvENZN3QyCHC0oQWyR1WbXwJG4Bge5ldev2lIXZ9sPGJQ
BA+VAbQPTj+FZQAkMeaMv1KC66CSWDbBxvRqyXq3JvaFXxFN+oBiq5G+35UntiJQ
n8rFFzHx8Qgic+GHjNn9zb7O6h3IC0QKq87vdbdOjTBVJ001XyDF9RjddL/0zZ5g
bqWiN0yZ3FOxI6bqVINermteJ0tnhDxmjjBfzClt12B1Q4xh7zNvrAAft3CpklGz
TMFR1FhY/6YbvAV8VFG5+Gw8/fhyV/tOTCXJLv6X+5AVH8RO1jLP7DZVnHSyuakn
UnW2u4zWqm9oM9ueTaW8YkTVGa0GtmKlHOgGwDRGOA6qYtzs0P/KgTTRbtNeyy0u
LUteIAXtVe3CEtotUaC5wn+yx+4s13tYOr5o2fVejGtrcoBPZHTrfT4EF2rnD/3V
XTx6xW9C9CUY1hfmYrpBVAis5BP02JHZfHMDkmauax/nsoe/DqMuSRBuT4mpn2nE
lEsB2qCFiuD0NeUNIPaEzG1Xw9a2sTE+ke9AM/NvK5FeYDGhNBgQGFA2XRhys6w1
zANpOfQ3CLJ968z/TnVQaJfR1y7IGJFdij55J/miN2P4hORqmwuoSkTAtPg+ZT2N
5zcNw/pBiXrfGzoXCVkLTAEuMLr/jdQ4O5ljli2/zSu99YhkWOKYEZc8thpXgeEr
z6OmiVlRJTv9deqeSzemg3Mkjmt/yCHLFQvx91XIZ8ffaw9APUsJqhC6biThrqo3
mWAH1HPwKgd7Lrh6HTn/TaLxx95uYVwJiRZa2bW4uXbdhuLIstLy23uSb8CThXZb
7V2aOiEKY3RO+HYJ6iTRISASgZ/FYiJhjiXDrxrrS5F3njBlP/NLPhOUPQ6rT5TW
BuL16V/fK0UqK+E6UrTp07SlT52LVy04auF0pwvvRmBWG8j/dCyjJ6crnU17M1lJ
Wnnkx2R6hAgjtzRprw4SY4y982CjA5mW9VfqLDg0mXUG2vasDgEaMLT+n/r5Z39f
6Jccd1e/Uz+sKB4LIa/BQPFT4CDxFttJt1SOrfwKQ/pVc3GvQYle04HQWLmVfl9F
0jQhg3bznAVfl4L5rwLCQuOrk96BR7TNHhz0+GCU7NCTu/gFMi/4yVoDJf+DbIby
RizbLhkWDCgzalG7sq4X3vYxAof+95fUYiN6OzPJUw2X9OTBK9AZ7+BH9IR/LM3T
dd1xP+LTXd//1ZoMGbJ34IIoj1LfGrfTw+wBP0goLGc6LPTtBd8J8F8z9oU9X9eI
trwgON0HgyKxnsC9HLRJNXm4SAEXB14HZvCZ93W/XxHItx0y/IUrXOznxkjSRDvu
+DU6RJXC8Whb4nfGxpdYVlaPM9aOlb/E7OwlXdchw7S15e7C1AYVT1XOiEW5phcD
6/rT9j5b6kI2xUi3UoCFg87QnAnBNzfpiYSrm/91SeC695TsxqeeTR2F3Sgov/wp
QWf2/zLh/4oqbC2Lic+BrrlngHm86dkznCAozcVcJMOBNA5ClKTuBoy+c9DcO4X0
y5z0ueDs+lrKuVGYrTRbcQODuVmt09kFwEH58IFpgT8EaAA+ohzVZLPgOt9E3EoK
3Qdoad4SVhqW+OyLYLr58TlaXDFXS5oUYbsIEfUF9BYWSSjmWJb4+nMcEffj/gna
j1gZO/f/NNWSHRJO2Thj2klF9ovQxkTk1XOyjewHr8+A/oCxLfiXrPIHR6udpXiJ
uqOLqTTynJEyxSfXpytJJBHFlDDXYw2flDhJpnhGqJCO3bYaLt+lfxkVlt3fPNWM
xi2FvOtmp5pQZJQw32n5GievbtNJprOpe+i6oaM48WxeUGcBSvYs1rcduGqticzK
LtLb9+e14hVZXXfE4VYwdMB2ZlV+4hPfRNk30ZUOahQRizQT7R25jzPlvbO7p1QJ
JLOOnzOUZ5orU2n/m64zbuf84wjcv5F0VnrAzYCPEwwtH766AcKxx7lZ47N6cm3w
exI5LsEMJCUGM67JfBAuzFwcGqvLAaKtOwd4HAlRq5LAc+A6N/YBhic5SCqSFHmU
U9GYHwPilku/sbr+l9YeImNiI25Q2CpYgM95hl4KDK9wG+RuIvlKGWD9M8yDodSe
PB6KjT9OE0RZjvrGrmp1mu/G823VqsnWajg5c8kax3UvE8hTtVmhwmDJI6rkOndj
1irVONrsE9WJewjJGJX3Bzjdx3njWjUSakwIHWcF+ThEdU2CBA9/fvuKnEmJwpCg
iDY/2b7c2h5gY1g3XgfaMGWKnxE4PpJHL0a6zTf1yYnrDceTBC99rUOBci7PvPPW
XRKeocVuuSWzYwI/WGNy0DxoHCHMknNctj7/aRBtZ3uUkD3j0rYQTWT+LTseFcSn
hrWR402OeuH4bSxyc6+lvs8Go/fMiGDutiSWRr+XwLFhIZGTjoUZjaE/jCbfk2lF
TLVccKKEhbalINW2DeQeK6w00Wn7nrIpdc5a+ZqM32zA/YNoyxJ5hwFvhB6mF+o6
LHyvM/Kt6RYB4TNWlOqo0YvkC4DnZ4k3jybPR9CNZi7Zvs04AyaEW73sR2TD6l95
nH9QLQe75WY54KcoefdD6u8Pn8MpY8JH2EL2Fn9nASm03TVr9cJ4wHgRBVFA2U8b
c/G/VqNNGwlDG2F7bqiqD8gZAPiPB2hSNdfJuRiHQ9gOipQta5FtliQOqpWXP8di
RuA08YiGZ2cWI7a5JDhJcTQ4im+nfya8slg0e+FVS9uqJLrYlSTC6HxiidPQwb3T
Dq2nAS1a3iV3z36G1zjHDf5pD1ynV9LAAZ6o729cQ6jdZfcGNHIPkwyDFT6khliw
KUacb5IQ2nhjDo3Ht5GXJFdPgjgwurZgTociofdQYCeva3hlZ8Nup+nNwJQgzS7O
UdHj8tUSilTjy4HRhrB+iVIlOkxSljkykVteSCUPZQnmSuQG1UfbmJfq3wtEGvRT
9oYp5EGUKbQIUP3pZV4hm+MozR5Y/HS+R+YpMk0klWKyjkD0+4hnS6JALTXyHw2j
F0RFAktnLXuNG1z1CTHzaXSvXSclP1GVduXfLf1rjJIJoSRaf5mr60izcmDNjzyA
OOK4S5cn6wcEhIUQchH6rjMj3hp0lw2D6S9jP98yu2XsyyY6bO+TVT46eonkgx5B
XHmZDPxaMh2NCqkLIcTiWdT02i2TEFNpaWm+pCyoJe/bIoUpYq5ZxXt+c9yOm3Wk
I+SlJ8t1RohA6RpzOYU6WOL5+jKCPVqsp61ohInqSAn8AmLYpqEGksnyLFhesVN/
V678RLRSspKIgzjutUyMwDppeJnMovWRQ45fH8G0jPxFUIQzdKs+A6JFV+zMqKN1
aAZ88f8CmAkrzI+kZIW1hC4x2b/JhclCa6ttvNw+7OGhUve1W/N2GAarHatff9WO
kdiudbPfxr/ranWABYFCEwDNPF1aRgmttUxKobJ3s4QFn6CgokNbQ0CJCd1CZYuo
il41hI+5Pyyrn4wkAvINpThBG1y2Oc0FNUrMIOa6WRjA3+Snc/IXSHmYmWRoL7gL
55u3MwgykAg9DvqUELm2UIap3iIMWK141JN5nQFa19IlZrrdiJmSsUfza2vJNkOQ
bSBu2NG4HbsTnMr0j5MfHMADkEc6nQNdCVqek8P6v9kMseZj7CEbV8KFf8hFWgkF
ikr1n7PzrhOEsAmWJrX4Ia66/t8iuOxq1uiJVONBAtBznpQf0dAEstzaDLpe7mcc
RmKaKf4D70nXU0FccXU0t5CrnN56K9OustWKBdtPnXnLaday/JLAkXvHiK2JKD/9
rcuheRyd6m8fYCRo0wQNHgeTmNQvDjy1ALkiwXXTHJzrW1U88q09Wt38/PJ2wLnD
R64j6KZwQ/qRhmTh0QuxfTbHKa5Sob+cbil4eda2aey6ynPkAyD9znzmNUQ7yy9w
0nu+NhEKR/QgFv+YDSbAwQv4odt8MYMOm9l9/HnjlKvztMN+nZjqKks7p6q8qo9M
cngv+tx/Chu52eCEortNnSVdCEWROcBVlo6STrdtDbEmttu7Eim2XDt4Z+Wk7ZMX
gI2gCSBb+IsLFIK/Kmyx+nUU1SqfpJB/gai6SkGh5FWEnizhcIs/EM5h6VREbJOF
tYlOt9ZYj/czlTEs8avZYDOVrOSN+DpaxQJIAknsyp1aLbqMPryUYqPxDaa/1NNC
wKjLf+c+oD9aKKySTCkt55eRumzObvbj7I9R3T0LKBvTgZsjsiVDvnv7fp9hOBAd
RarSLE/+z70M5nnziHVvAW/iN7DaCgLyYN0MX/vZfdY4TckFW1+Q4j0k8j4n2jUV
62nkJBMCqg3WZ7mGBvQSfVqxorimr8FE0feJsDfgvWX8WqcLcmZUAEomzL4QqKzw
+s4lbozT609tCCPeHUbIdmNVbD6Rw1DbgDI4WtHV5s+eGbd4w/rXS5YEZancLWkc
IPBa36T6+CSqpT7r8SJ/qYDhLeMxIGCUCUach6s1SBGnYSoQnlPsRirbflMSjxE6
FPPJeCRulEGyqd41h03lpRDb60iEglMeRODEZ91wMB2KJM7AEUJ2SoLsLEwdLXl7
YIP5iSnFr9CkNa7kQV7lyTUloRSGS9rnOzNDvMfKGqjRXcJpThOWoa34+I0j7UjB
gfIcggV53R2sO9x+JQBLdo3UEipisDPdd3qHVQ1ItYCgo/E50G0j9fQ1mOgIS+Mh
dsZZZeUYQ7O6NoDiyHyFQMDEM8mKjVSCUZ50RhTJrtm1r24I9rq/fqziw5io1pM9
16/OVSFNEZldO5Enem+1uPENq3AIFwGczr0lQVVFF6IqUAq/fWOU6xUXtHPTf//1
yJvW2uCxlLXKj7wN/vszymT9rz1XQwoA9cX7EaCan4ynUWIHKWvquqUrrhcEnrV2
oM6wv7Vf9knlgjlKrF9ELGv6gaBssEW18EVHnLIEKBtbOcHQ94nDYK4OSj43OMzl
p8DEXb02bA1yrx3abIW/yYh10g4gPV63YztucvBhB42Eib0Tnq4WrdPrZf/TYT7z
Hho9lnxaRjKRuFa8NMvUytTcqi7XDhmaWCjBCchMYChrbzXchs0F71HlvqL7ocV6
TU7Tjel1KTy7wTIEa7SyUyODmf9Qf+sBW05+zYqABfxCt4vwxqbj2/GYH+M+J35T
emwjdgGvSSajNV/0yXnoqANXPB4P76R4XvRceDlcrh7uo/SicavB9PhMDwnCyC/z
M+/ljtAcmntA8aTULwgX0M7KY84Vg28s7dum/4cOzeMGdTeUgmgGwO4oJM9H5hfY
fv6Q6TnbivGfpF6cH8Apg8pJWxq1qMd3mlR3jNNT8/67ugGyEwVjg6shBMIYxTA8
QoY9EuYaQighifTBtWKxsGL3JH2VJaUyXrdpPpe1sOJrXS+m2iyDZ41JZgHTgz7H
ILr6KVIuxp1ZXw1USg+3lygISTeHCFw44FjGzSagyZcMl8M6XRtFq8dPXLOPHN4z
6PMP/J0tyFScx4+zzMleiS9bk6aGFizzDXkjXiRTt/ZEdS8pB42CzdZj1sm6QIwc
kGlMLPZFF/DO4K6siiHGPZojpi/wqyJ0qLkj2HS7HXYF3gt0AulnHYoFH+0a6ISD
sRcfvLsABJQ6UDdjj42aoWej+vAsKjvhPDo5lhAEI4p0ddapagIjsDEn/z7yF7pg
3y8F1mSn+ccLObbuG+vDlo6Tk5dUhBhvB+Rb74LcflzOA3lnjOMX3g5CZcbQ7SBV
G6WZRmLaHsgxD322R/X2rWMcettuaf3+jjhqB5n7v5kwuk9C2Ez0kEFT8N2NHj8+
+tgoqtm2Gfsk7TytAPHi+14xL72TH0OJvCCwIti09urNTMXbz+d0+AgVLVKP8zag
LjN7DCRD67M7B87g/P14t5zAcIwkqNratIPta45Y5r5SrAkKNMO0Yr56h9wiKBZb
cboGVdI2BuPLFxMr9daCFW6mD2croesFF0Rpp357cEZ1nFOXdFG5hRX1at8Bghb+
1ATBDwmQCiI777hD3oySrVBBVNrrMS4IAzsnY9rWTjqGy3ShCJXvtsu0F/Jlt/40
e61H46I9CVJ02fkPcVaPmhug23KADndClX5cGNVIVtMCBpCN1VclyWJ+BAg3xeZX
IOKqosjdB8Wq35CXn2INtntdF8twOSJ9SVoml6bObCRyoLrzWNaV2wCksm7nLmwr
NkftPOlcspi+pPISR7+Hrvu8BUoyfdRrDryxEoeBnmdVyvReEmZ218bQjcC8TV/X
XwmYEmWnaHAr+VEpFF/oNOwvQVcgGMBha6yvkU1L340lbVlXVtwwv4Oe4rpbUoam
6WY/SNCnHw5vlpX1u9oS68aI+5zDBHcOe0NRdh9koHfiA2/y6W3Q/yptfNcl1ZB2
HKQiVfxP89+KF+y06iPOekuHoi3+JdEh/Uo5U5b+UY7Tzt6LSlIhH9Sh0vfP+IoX
Pk2g2UMBhN/8w7t5fy8daC8oYqxy1h327yDxjF75WN0523vzLu43qfnW8SSCNK0D
n+Y8SYXWvPdJJP/xfOB1d5YXFeQ60OXUvY8D5WQ3gK0MIx/WyB0fP3nStVQt79Mq
W3BmoTT3nxnBbJ6P1wuSxcLwTfeZ9cSUpfMUW5p+lTMHPJWbSHeFwUDmYOl/hWmE
+BPkefEMSh/o8D1STI3w1MN4q9awJz/B6be3GnyXMdjcfZg7iWRLAhNAQ8Ga9L63
WJtNQNdPtWCnLOC6NZa+W82gJdRFoIekB/sZx+H2ZHRYlZWAnkxdJ4SYNQbJ8QDX
kQEuFIKS0eeeyccsJ2eoYR3mzrRuhbkIFjaRKEXzO5ZI0m7qXlRjSu3aaZjw52tT
KCPgP6jYOlg1WLqIyMKF+ZJJsVX7OOPbn8Ngyt6j79dy96lQEAhNrH1G67e9PWhF
+Rh82wnKNAurRHfNtpyUmvz07UOtAzp8BjukWOAUp9ksfZKSXDaMjOQQIWboS9EB
O0NgtN32fMHR6bwtU4uFEq87Bz68G7C0kQ5LlEUlNTfvv3JvwvPmfjZ8H/41XrSY
dTMIJF8ZygAAmoJCrVOrD+xV6Kk79HhdeQ9/hjXQFLMZQG7zdJ8P/Ixcx0yLAJKd
jywW6qxjCL4oEgSEgYPqTfw9aylO5PWSmDDwU6I1R2fP09ebciXp3q4Or+aE4ZK3
W/LkWqWmMOaFpgL5w0W8hVXJQZWdnXHPRGYlEPsyPMJZpcF8vjYmgPdCyWki/PAb
rB4khqhmczwKlc8L+I76+zWXOktbizn9hiwdG0DLafdSUVEV+sN7eIbV94j+AreK
/8vnoKyX//YoD7DlxwfRmPJsPrLyTIv7C9yAKS4B7vtRmwDHQS2cDNuZIyssBzoo
qww+wUAM+i6I8S0x/jkVhaokP7iFJ6rh+tLtSX5AMI8paGggqX8YRvdLvPAldKIN
Rkhjq0uD8sBbgy7RdmsuT4A4ehJU8EJSzlWyTmGqm9Wp6JMvCNGT56qKibNB8Ud1
zrg0U3g9YVGEpa9/KTLJH88QsxX7rRYOJ+HiXKoJdNPSM1wDTQBYYmCHvr0GA+O3
EGZzgrouUEkS0oapb9IhfAtfLdGOqj97njf0P3tjtpDaMlAE69OMErVl1RrqmnRr
zNGw2TXoL5BuBIDPj/I4udsd+uhXL0j7sA5gne0uk9whLWleWQvI0W0SrZUE/tBy
6ifF7V4aBRjForsJEoo0Tx+r8X+2rTTeOLVjHZlfoJ+AyZSA1aOmL1a58Ritbrtm
WzUtt6SZJZke3mr5T4a4VMPJZDSrwVr+b6RcSMEFGPdeCX7GjcO7nZAxpjAk4m1b
8ri+cfFddEVBwGzne6AgvdcotEthZfz1QipwUtOt9FfeqDT/2SXtjVIdJHjuYJTP
WX2bZbjakYVhmwVXJDeNtqdOsENylc4BqcCJPCAHyt2N1NJv1+4ja6jnuMcnvrRc
N5RIs8h4tTJwnKHl/LcSUh8pdhDvhqlVMgtP2/Kwzs4fzYu4LqGNWJSdJPe9bAbq
xTh9UbXlHdm+32xRX4yQ0kioh0i7oVnyzs+urbSy9Gh+sG9rzmzdPq0SHTcU4WJl
FEE9lGLVBGk0hiSuS31EQ3mZHK4riZOa99Q3rQf21qdKlzGJepVls4pdy2KBG8Y0
8M50BjCnPONsQxo0MIBldJFSx+GZIJB236gd8kBWIhZjW0+oWK8r573gCuzDzm5F
BafR8doAINpwo9Sj+QalhhId6u8VWYWqAR1KIEAYzxY2GTXnEUFzkZkftqF/b2zp
PiApA6Cj162VIR/sHib695pVXrw5Nm333XZ3Q4nigWoYEJ/VFdLXb+KetzfAGaBo
AF6/zzYmKnjRQFjnvR1bmGrb1pjeLtMD/IT5O4P20iTvGRCUdtjDvjYn2Jf39LU/
nd61R3MbCTCkOXUdeqeAXH6ehUnupvJLAuZr1iqa4Em3on3DuNNPwdw39hUuxmxR
LJspOErgxG1AhAh4uBFjdWM6hjr0BSF0GE0x/B7sxOElAM+zigs3OceBrwn6nlUN
nGfKwDb9vcT377z7ktNWuFQdlidju1EU2nv7ZUj5nxyVJfw3h8AI/P/E+2tvjPLQ
VU1yY1IZ40LEa64HYNu/2TRIEQjxLlAfZ3PC9PyAAJTn6CkVnnBHroJ72ZcHqAtl
78lqzuX9Iz7fRmKjdgrpUMyp1CF1cR3L4qUXRszML9jqfdfcuhYzNhl7QfO7QCtg
7qgccZXnxQxfC9ZTUdC0Xj0TFkmJEjFNYuf64M7M5BVqnBMDvxYFYJz1WoT51r1j
i/YEHRov+cR4Kq5xyt+f58P/In+pHCGGOHEt1IOZzEgZcxZGrsTtGKJ+dodIqZ+G
GWRFJMtMd5prw/kRPyKTeOC1rn2fKpOtciLoovbiaChCRE79tkn6j0a9788u/hUm
VlhnNwcnVICZaMMO7JJjsvw2RhQLzsroI6ibYwyFILLCR9OSMMUc1kUgF2gvjUs0
944fIlV/rl/XZtnSa9neudTB8CCKVhG4AP3BV5sxwh7C3Hqv2bx7CTDZt/1Xj8Nk
OBcJz25zU/hxwCx2hs+Jz/8D7w2oQ+T9junTm7NiHdRklZCg/GemfCrSqNhUB8YY
O+uqGpKKF/ZG+XmK2pljL2nE3EnRcQP8Dfzhl29tMnJLG/fgu0GyhNHiHgnhw8Z2
Uwnxp2LMOV+aCnHExWM077YGTLmcBPbJLoSpp1kIuD8GlP0ZKWTEEraVdHuLOgGj
JIZ0zD8A/VEQ2qiuFeNihylV2iY+A8cI05h0C7V6FiCKY0tGLJ5ulxAT+gIka5Sb
0h41G1W8JzpJGRqpMlwTbx4fR3KNeDitPqa7W18vT1mN4Z0CYys3g+FCW9fzZZ3h
vA4tXJEwFZW7uGSWBjkyEt8i5ZsCMk/1//CcGWJ4SmxYDE5ogi0Xk7NpnY6oPs21
ut6ZPx3NkNMJt0/vMLJRZLOYaevP/aPQYDOQHiBRlxNSZ0+D/CqYdsA/tSmuw80C
Q/DYTGleuf9Cfkby2WeGXxAikblLkjfjHoebaICpz/zfdyzZ81eXGRm3Zv5lPxur
5tWaxCEfI4zlzCfkz1RJlCInQr5EjW7okki6j1uRBNUvgnS8EcDOE2HdjxmJaKyR
HnCo7i/TveiRgJCH+E8A1+epKcynDdxLSJ6jg+ZxstzJ9NuGTyftOdnzv1LF8w1w
kUa9LTmgsAGtinqui4KY9gAmZ4klUGSLlt3DScWk9f26MRxiWZ/wvRrls2K7xPTH
Pp64ZSr78HVuUiVpfyx4SeTNexSMLxKci9XV2nNKW/r+ywQNBKQZICs66c4xus8X
hQC0XKE4Fme2cE7dSVGdSaoWU/TVpQVJaLCnrTKVH3gO/k7VLhWKBzK1nkx72zpS
/tax+lTEykCsOn0kU4H+W5yPh5pT28TJFziLHpNCa20VP9KBFtdWoS21Emi6SrXl
zFsJXPrWahha0/+LMvoNq1Rdw6Y/LNdSpKpn21MYN3taBj5QBY/nNx5YrAMq45Ar
Sososa3RGKTJ+E/zSBa1B7AuavpQ4uQmi9qu0180NhsuNnehWN3LM+TH6FTBy/Lv
H54tLiaKkKHrMUkuKAdXaqVY1+FfzEcT7xDqHwmPJUQ1VmPRtX2bB08kRBBhmgie
eyUsZg4ieoHzd8PyYteqXFw0WBGPtI72B8+5K4Jhdar2Gz8WFv5dSkdUlI9vH9a4
Lbh0zoyyv6pMk8Y0LFAOwHyn+MFeMjEfOYuK9p9EchdbOd+cYNpvjUWhC4bdkL/3
jFQ5ycYi4m0GRCVLehabqH+ICExekRLBdr1z0xS6V8wVIb5VbTjWGxqYl0ba8VKe
mm0HovCPwjRbxgdBs+mzVV3Au2re3F/E9DSz/0PRBVK6J36+4h7YGo5ENwsT2w0h
FXn1ZIVeTNEcE+8+5BJzyo9jtpJUUeVlNmuZoQm1eMTFK0c3ygQHRn8p1jybXQZe
LdFsKCGyO7I9PdcdDEIUqInLonMg2PMXtyyubCypl1+ZpS/dQCoN4vbngbqlWdcZ
77oOsPyCbHqD0+ZZgy29BLZBamlafAWtQDHs2nwSSa9hL6G9/OWGjd2gF5AmxF2r
YT/y7MsDyaq6uWqrxr18UdTyVfpzWttMlKlO6HLGf+7D5g7PHw8cmXITtdXU30UQ
LK3ULbpQedXJC+TUQobxmXj5yEPenGyEqEdEzxXAEha7KxsboDt9ALAWe6if86Zo
TzMM8NxP7oZ23dFYJx32s+l2P3m9Yugr3+eyS6Z9WLq98K8jE4oBK4KuZ265aGZF
/Hiucl0Ryb97pNrlXeOOS6XospeBxFxDeERdAclM/niRb88U9O7TAAVCXPRYMttC
cYzFLVN+wE5IrFzh1m06QR4pazMdd3JlPfUS5QWbQgk=
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EwtCDWXSU4t++fc8bxpeJ3+Se1xCvEnY5n3lQptp/rwc/sJ6rXf7S1KGHgsj1cgA
aTKkBMAJGbwXSobailnBewJHTavtBT46kixkhlQfrABGbOHAagWBA1adAhXPNUUJ
DGc4rsqQWkF3vcYBIzs4hLHr/qE7FshpsfGKqvQ8x927mM0BDdDuE6r88mqz7j30
BwiaVBGFA96GK6PiLXqG9StZukpaMH7RaEAxP/+o30cT5b2lLn2zoKvVViNqh/VD
TBcnJRv/i/+xjkUPIdm3KPJWWJjqqsWJ73K6Ec/MqmEqsIMFWjIb6CiAmxlF5yZs
ua20Z+DT2XiUW1vJyGLXsQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7216 )
`pragma protect data_block
7qyet8EhrJtjY6zg09Qdfii4UhowWAJ50ZDdKJyqvVh6JAYVZRgpUuYn7SybBBLM
kWAEqPkOCYf3zi+ZPmaFqU1crtVKxiEJGKDVK3XO5sTXmUMimU8P7GNUEv3j3md0
SG39jO3N4scm+AC3z4rxPjo6cVzTNXUqqGV8t4SiBtx/kZUgo7Bz3JxwFyZwpTmW
6JyGSLnC8PJqbWJI6cqvOKavx0Q8CBQ4YICbDvojlrxk1amo26cLFLPkGl31z4ao
G/fpcdTjKi3K4ly121/bOZSV3eIv7d3xgrH0nCeQcsfdrBqyL9HVPBUXSgqqFJGC
cpsvtnQiQGmbe8qyUQTL1F2rwb3csPhRfLOwO++cq1MjMzP8d94y0c6cQoywkETS
oF0WPKsfkU9ripb+uA4BHV5xxIBMOLhs5IREFWVb5fVj3+/lEXzA6/fum0+IIF1Y
bVGcrfqU04wni/BPqyDU4unxDUsOVlpdoZiSuxiQkhhLA0TzOiRdKFmqJCqxgo9J
4PlVUIOSA418JY9Ony8witUdvhV5/lkTT2n9Qj+T7Zi7qHvSk7FKRHJ88ESdJZSi
wmpwxD4rE8I6ZHrjLlWaPbEiiHVSOACMMrwkIub1MB/6JMCGqqqrGwBrvcO8br5j
pynePyAwmZx+NIBqX5czx1ub4MTXL7WIh57e4oEiJCzarm6fDJgZi/u8DF21JPr9
dw3+EDvuDHbonfDktlhjBsCk8iJ4Z7C2GWhGj4vKbTzbNXGfE6LYML+vgZzAbu9Y
iUkA75JLD7LnXzNDsy0onTR2ha51yQytnQWzbwviiDvj3GzW10JxOnBWU4Wbjfhc
SCr5ejDII65uBNHeyipJgIuHBviX991RCUygn/ipgPLr9HRZm8IHE7Ii6oAVHjEk
bdvz4cS/+mk14vCB5rJclPLnDrWiJXcNkN1ZiDQjAsjEG3noeq7b21JGoZo9w23P
Vi2WX88kQDzPEJTgWT3WVe9M/K/0NxCnYVoqKFsGzpSqewlCgdyAhAcsn0yyywbr
yIXky2lXXt4N5oVRAXeJpIE6qhY8eznh0XLncDzQz/Naob91s2WJTImYG7jYiMC8
M7QocuLYh7udHdZ3mGjABhslO63i3P0hZMB7GzVaCoS+Urktq4cAl2HXFGcsJlKG
Z07nPWK/Iaj+QgNhcQvKflrV95W7IDJ1r9DFfCqA+7PiDl5dIG5GZ7ED7omZ09fb
FZFRMvfvAJsrFldxz0a8zAD3SjirEMCyDyNn0b1FAiwahPf6loKItBDHA9d9KM66
WjAsEaAcheshmnyAbkjJjaiMn/YUsIKvFrloB5btr0e2oOw+3LGzlWSW1k5jsVpK
SJLSROv95ettLvALmdJAYo6nHVu3RWwPzE0kGE8M32oSiCT15O2m2s9cfBucO7am
SeHgeYI2wmUR7LO8yHzWziBUiOFURG1uchHqrnuZNfVIV5OIwOHtjfIOdXj8V3ng
r8FBcoyVJkg/kXmtoKjcs3GP50qT4X6SV0s5fkDsCEiDlGfXrNbxhFeFVNZQz5aw
gJtF440ALjG33mEN3w8dBUefPxqr5T9Qng7lUP7KNZQvmdvg0NDaRqyzKKetW8/q
x37JGBi72dNFJMnhS0NcUYBIrdWB/pLWiqQZfUZ1q5MgPf7lDH0NwdH+JOifunTL
eFVP4MKFIY6mVxcmOjVcjjNCOvTtA/pjaTW5fD2mB8DE8JKPEzAyMAPFq163Hybx
fBIN0zRKlCxBxSu4/tTfzEMjH1kJg3TPzvs+dhEc1hmnjzDQXe33lMJxlVFjbq+J
GUeQt3EOv5fYfrXJKVcLGLczDw3b2fes+6w92SqUJRfHez5T5mlZPAVt+ISj/LHF
WBen2RmRTdmPjmSkOH6MiWTG9QlA7IpnZwu2hcXmJd+GduWFHJt4MWgTDZM8+Tot
4MUoAwsd3V/fGsGajwEuQyn1O4eSDfGbIR/dqyheRIyww7e27ww5d1iIJOdmilma
pocMVQNgJd/Xp69epTSnLmqyZQAa6ZyZy5qngFRn15HMSc6fbN3v18IVUUeIa7sY
736PmRSPIPiP7g6UNJCBzkVPZu0tO4aNLCPp32jlfRykXZz2o6vB6GhpUDBWtWMQ
ph+9LlR1zq7JcKr0J29FtDt5E1ossq0SeBdge2rXId/7DRHI9JKEEqzRi41yv4lk
lws+cvfkuHwyPFVVb7b7Qou2De2ThB7Bbj5ca7HFoVyshKt9TtHcUOPGtjXbSMtq
pD9TN0f2p6So0x1rAWcEqG0njdGN9w2aM+SEQKE6Vd7PIsBTQerowUaLHi82uSaW
7m5l6UXCOLUK4eIf3vyN+SDn35Wx93tM/q9ypbgc5sVuzgJ6RmRdRNK7Kz5+l/Jr
nmjKzwI8aBp2hw6pbKFeJdcLP6GFzyVtCt4gCGdH51dWCz0yoODSJBO7DWxny7Zo
fNChvatbky/gthRgsT1fYMy43qdfeSuMP3FCsSK8+EGrtUrJwqFhPpOPoN8lmIYK
UujUh3wgNS3VsUspq5XqFHaQcPdGvbCQnP5Hed9FgiBJ8kFDw5Gl6bvCBho7kEXp
pgxG8fAOeJsTs6OGRip+R0+QznrJ/v44uxnN/G4Fh+BJxV2j6aiugQk2XjbDZxml
D+4YCvwfLndcTSXcwqR7s8fhP3luHy9C42s09rU4GE/aNRZyWzVJqC7qn7Ylm4+O
omMYjVZTx3xBnDLlODVjIeeFBOMASlsoF3KxMNi1fo+Q1VVjDPHQXi+e/5pmRkrW
fqMvmxmVJMGUruUeFrBBO3CtbbLVnZ3T2iJ8yduzsPmCIcSfkyIN8oSojbbxOCuM
Xh8C6LRlZvmkNcf6458jSPDaOLA4uW98Ve4ClkQyiZmVH6z2kwSvO8vlq+QdB8xU
NlrrwG0v0o7jqqnKZbNQlHpPt7L+yQrfUVHbIM727+5xrsk76Faw1fD/PU1rxeJU
UH2I5dXgc9BVeqAxzHCg83E6giWWgyX47caC3f+68pd3vEWMkQW+XqpXpvG2z6q+
fgup9ho35xll85qq6OMR//JhaFGR0Rb7z6R8/4dDTXbTzHgULIDJLHeWibQxzmm1
N016qvC8dPL+vBwzSOdUnA3QhL/oYgQEDeyhLqMabQ9EeHbiLUiW/UEBYO/vkkwr
FDr+MNJrnQFQIg+JLBr1HbxTuZDdLxOTrlbEkyjv+9spx+NRg7aoI8i4xOi9FeBt
2/NwGyeO+vkOETuqJEfeKGTPM9Qo3egykp+mSDPkQix67MKHwEGyaUDm/lAdfkTk
EV+ysgGqV1OFzc4/KKVBDaxYrMC8Z/4AX7D8XevYeAG3pxUvr/qyTivIsa8oM0UT
iRrZalr8ru3c3jt3XOJcwaJHH9SvuKPCR0M9/zqG5D1aSRx92s2i3mJ+6A03F+4F
9Sz42rb4KbzqNV60VtDtgtg/3bjF6twMa1fnSoZLmVfwfgn99N0iqv2zUPN4/JrK
fFBiTYrHZLuyK9w5mwlUhTSHsxUowCQ5v8q48hj0IX+dn/AoEi2TNbm+Zfx5mAGN
ojPHUxGMT05T00wZf+SPqke8xeiLcJvgjv3K0M5d0OWhYrV+AgpaKuqQerOv47LB
c4TLkL34zPNH58KxGb93yo0a5Q8nq7CPuxYIvvQ4/j0OM2f5eTid6f9bSui+SirZ
4bRyZv/jLAURftfGCuRkRIesKqkfl+1BOCqAJnN00s73rzMQ8dHJoM3uVHuY4eDt
imq+15EXR3F8nG3F2PjOvkhbhOxQCSF+fjVYJIhv2kgBAsMvlECnU1sl2FjeMsVh
uHF825Pz3vPtfIbR2SgZGxoBP271A5zyD8WX6w9Xm2b48KWEFYee2JU4xp8z6CX2
bVfXNbjC4U+jkstvbMCExs7fZqFYrEDa7ogt/VPjybr7c+yK6XbOtWcWk5psDO74
/eLjBlB5maxe7vhgFM0DyI3XU11uVkbN09xjcYJbHTZ3sWh1tgzbI4nu6Z5hlCuw
3Y72TxIhQWxmwPTHSa+8vfoDTm1Ktirkl2VKWA3p07xDVUPu9fgmVHYEvP4lEhMN
6LVWajC3MTn+yooD6cC0cjL2M01P+j1HJP3PcM8glj3xGkprTqXeRkrEHYGzKRMK
hVEq8tqabDKs2R5ToDLEHH+Kmy7sQiKFlmDJ2RBLHxPYsGQkEVxsUfmvw/vz+45D
8fna7hhGYsGLAbcOq3lyrY0JdBqPrCeMggd6QOlhL6hDWygSiYocUB/7YKgjQZ9Q
ooVDTXFpyuFUfExJl8kjkdNAve4Z4pDkr9tivWlRo41kJ+U2vsJ1CsmoezcozPnQ
bSao8mOPmaezpd45wxq+5nguu785fdyI+366NbQ12fQEsSghges4TUHTp5fg8ueM
ZKMZ6ahRMawYKmPLaLNe6Ez7jNx7guJOfehJtkFw2Rq2eyQRGi6RKb8CGQOe4OB/
vJD0RlAGzuN7x1QlutC+lTRaQV4NXDAcG9TVeHGarDKRk8cAvakqdGmGuXpXAUyh
/oQsixoJltwMUdQwgEIUlraxJYLsb5YsQu0F3vhNgVfNtvcCnS3nb/tpJJBDvz08
+2VYB393lXIJxbXyWC0hWva42evr+u3ur8L7BTzkuovRiTCdvHXajbIrYhYLUoee
69aoay94fBThbASaGd+GIgcS8aPCd3ApNFFmseg7mT+UCJvEJBcsGA67oFD+B52h
VB1Jg2YHGVy4PhxaYhF023ILCTpuPiqeOVE8tE5dP/vcQaRtW9nYipN40wsmdrUo
SPtlIhMfZRL/iKeS88xsQHIQueDJ41qWeYieELD3BAcK+zggTsVlR5tepgfygx8+
ubk76QGbP46haWCcm+0DMg6uOPfNEfri3Tu5iDe7MViY72cYwmgxloI/OFcu8MC+
vQ7f3GWSrgV49CxwP0ZzuLcLnDOovFeSiCHoMb0aomPo8EtOT+bEkujInE6T5Lwq
ktwz5QFWqAqzFK1f9eWjdLqC3jriLxaVnNJlSAxZTsj74eQQzvrQPd14v1x975Gd
o8rfbHOH5UK5YaL4ToSAE/h5DxWourNWpAtVUUaDznBmrwpLJnncPpSnLk4rhJ3Q
2VH1pF7Zg0lQRvhi+xeMstuPNP1Y8hpaKbFFjNAQkWSWuo2iDpAcxnbWYEacPsCR
A/spuz4x334E+gVhdweSy6BWRDb4cAGfS9OhzbvulNd+l/iyfpzXgSDsXIb944II
OE4bjy173aSRURCSMxaw5BBXRMaFjVyHPC/+H7F57qZO2k3zW1zNFCxD4QhBIoLW
rUgOdt9JWnS7YI7D8ZYDw1nEO5n+qmm3GQASwqqq+pEWZtkE7Q0GoadkkgyF23XH
B/mlui+Z3FtCreiJOJCO0lBuEl5z9IZsB9DVq0sBUtCA5G/yzsw9i8pR+Acah7vQ
y5kWzf1CcQaY3HbUZBf9noJ7AofZOPDRD2lxDm168MEBMXb/ajEv0UBu59I9wvgw
aRybHUboWWPdJnapOfugXMw8M/Vz4d2mACenDtEcM8TU2F4qlreCkem/qYPL8Pso
JtLmo9wXgXrDVG/WPSuQpLgh95U8AJf9sYrpgUj1r3FRi0n8yww0T3Ln4fcAczcS
Ml3odT7wlqgWFyBivsVqDKOURgCSHYhXjNWfOph2Tl4GVIj17FdcI9132C+cPnWQ
deMOAAn3WDO4h4PxQnvGNC1Nx5LxLS3J3XdbkKoqQ/DkA0lLuSs/O9sVkNJ+qoIF
21QlQv6USXaElYDanDO5fVCN2toUAx/G1S0uAK/DQsQKBd3IB4bUyQ0Qo0luFxb0
5x2eWNPHLKliHAbYFpo/9CVyuGFYQOa5Lxbg4QvM8X6oHwLGELulfjyWk4WDDrM8
UtmFs57Dk4zMl1kzpNZPOqrB/mWy/vlFbl1McsEUyiefDeEgVs2Ir/PEt+4nsy3v
nuc9QUGdSAo8s0qwdNv93WR1bsYAopAggFrG/qsRRp6WxFA4cYzh6Qim5/ArOMcI
zl038Z6glUfLX8Rl2kglxN6Pb67c2Kbk7dWqUD26NW63saxp1qSJ/9bMsv0W8t8H
JZWcvpxr4sCZ/N7Bf/ljN2yPWFHw1x9WzkdzA3haSZbNUn6x2FZxqYPfvBeAe4LE
Yp5RAjm0UY6w9EHGzR32vb7R8YCUvQEEbHqY3wKgJkwnxZ0EErxP9NNzNWZRNX5Z
qAJXKmLbK1wnLyooLrcjXeFvp5vpvncbx0MACqD9Sm/LRryy+WAd8lC5bIDnaby8
p9J8P/hIzmRXHz6qqr7V1sVfNRs8WSn8yWzhLuHUhL8rXC7BaokoYxVjrDBHBXfJ
6usA443eqynivij+M36a0rHX7DLI/l4LZKPwhwX7yqMNhGonXiuZR8ni3Cm5JZem
g2jBnNRpAVN+g46W2szgL4RbpPrEz3hIHLxh8wGgYjoFTjAJ/977Lg4u23LMUeHg
3qTPvHNREvjxE6ocBlIn1/8rBhVKur8BFn2lFptKdYp29PRpja12qhmgbTNPl7aA
mh4/iZnEAn1yaUaAtGtpotcTEAPMm4iLmQ2h/vU8iAK2S3Y8hBGawSd8CTNXxWT3
CHc5SmPARyFphgcujglrmngVcztOhYQ2BuuwLJUhz4QpdT5rakUPxdxtK+94vzpY
iWJP3RTElcZAQaPEWkrmwkYr/PnlgKQclIEmyDAQZi3GnM145BhyQ37g28p2Fm3h
vPi7yVs21XmPNwrbyysN5T8r/5mpBM8ob96WCGOZjMui/dh1zT5ORz/eTDLggdzz
38qt6PGrcrXsC1p+BTytmoLDJ2FwDdIEsT+ZhdJQBaK+KNgb6P8xq492J4Nh/tt1
O2BQydMdE4PsJsCVD0C+FiMBZXy4jL+28kgq2lTsXiTgu/CNVR9beugPgjuv0hsC
E+IBjXxhFSpaQGosMagX2px+43h35sspVL7xlF4xA/egdLosRHd7VZL79V6c1QNW
1gUuK6sqkpndNAsq2NM0fKNbqAo3ryHD1tXq2speDtvs+4TrqYLm4J/i+7FeJeH6
SB62odM/QN1yBref8Ci/Dl3FO4xcBgAcWHm/RZFj4yU81IJxo0bW0PcfjRRwfued
oazCZ84SW9kZ/xnlJuCYzFGI/t4HqK7ibWbuhMOn+NoCCLhRaEVoTpZT/l+IhBzQ
EvYG3BFk5E0V/2tbGVlc9Zui9A6W0xZngoBTuOIcSSJFKRaPNlV07GYa4pR6dpeo
FHRk5dHUefHqCnZHlKpzD6ZteI/nn6GrHnnUy9XyOCUOu3khMhZJzxby6b2ahxv7
CbdrV7kZ2DE74Dz74R99ZTZP1wh4JZXmRT61WNF3N0DI2hf2VhwPgDRf/XP1623I
8VVZ8stp9xXmILmhF+a4YuuKfgETAOyyAsHrQR3Ik+biTMTp8SowAkO6WUuXRNNw
S1wqweNuBmwcMP9pztUARR0F3s5IPrFtNCMosx/nPnI42hChRDCphUejOAOzAdX2
rMxxBbyaQKc93o+se5r4ZQ/OAV57UIdpVPC+LbAQa2xLnqMVBXrKBxIYuFrboeGX
sKjpfnS/kgkxuxKGeqIcZLuMappOIGzFfpgftioFtW7lgyELxrWNATKHSACKWtEn
y+geWQ93UmM2b3XSKrDI/ZuOb/bGWNZkRUTtg1X+2ILRK3OMZ1hnSol0WGUb82AT
uTjMG83+m2r47B1p+Yh1BbqeYsnwgPkJqI9loQAlYLxtBZ08C9Ij2tMG9dK5NHKz
GN0vQM/DKTnJxYVDOE7RcFEld/qBaxL4bEoc8F0g1499vLoshd2SLCVGBFY4+IHY
lQ/LpLe85yRigvQT4kA9QJxCroGgvWH+3o6yhG51HjlOQLaDd9hkeLFUoWKd7Jt/
E8Q7Y6c/flMXxXwuI5QKzNtic6evM+c3DyI3qHrbgZ87j/kIuLCIca/fmYd7vs9x
cPqqfjmCb8zrDmHuFooXsVRZoST4cCu2yJlkIOlIsybnnzjA7YoKr7mMdEZ3FPNe
nvYsfZSqNVSWilwzQBNg/tqeliIiEtrkxhfAfSV2fX+0c1dOAvb8Sh3rtosR0nuH
5qDttYrwTCgrUBxYhT9QLsqSC8A5d/tfJ9FgeqigkIOJdpzBZNOl47xmFrK2JaiZ
S6Q1zPxr9oIWk1nQzZIR/enB4eYWZS0sxRpGkogJcpD8UoCUYYu8I7813zwiJAW1
VitAcI9357tkQAik8OvrQV38XOeKFSzB1gj+BUKfUjEEsUr+SiVS4S1NROTuliQ9
bzl7pnN2Npvc6K63TfjUlawqCSsYSB3j4ZqfdhemHvZdt3qv2XJtsKXX4YmtP+hS
DJxMBHZORwc7nke7INPdPRpssG3h+nJIlqT1NjXZgJxhaZ5RP33eUHHwZqdYdOD0
orlPDzaLo3iX3ywAqmRYpNNXNO8Pviy2zPZaMOipelPS6IiuRyNw55jsOc4QsHYd
4o2XKAnOV20nf69j9z9i1QtUD5cCslEFEoByVE/TsF3H/rFQF7CzhBxMhnVzg+uK
glIGnBqRHmGY2r1rh3G8U7ufgcpRmZOndhOjMHnW+H8QUbhqpFJRLMpYUuQ9AQN5
s+rOGk3XT0ecIohB3HA9Bb4yoHvHwGUOYeNj37EMSlpiTgOlrgZhcJzr7ApglZvw
eXX2JN+4SepV5LEiw47o4B5YAk9SPRgb58TVpcFC409mPvhFzQa6osWzK/x2mDZ9
caoCNjuUUfBVDGk30+yxLG6+niVDLoKOE2gm51sit/iZCAQ1HdpbDheNSEaDFhse
8YHnx9HJbDL3895lstIa8dxT6XIyOofOwcxyaBfszOPTasCM6lkUhyJzpXk9O4sa
vswjOF0eastiyUWxRmuNrVLJkKnf3RwqhyMAoSMGv/N3WyC+im8UcWEvk461kiZU
Kpo6a9C+L8pAx8H+eC937+C/Obgl3/5IBJLWVN5PXniLfYTiyEqy4tM6Ng11Jzf8
xB9+MVa648jaqwcB2k8pzrmqzaA07fQffuDDJ+urkOOApvuaneTN5kLpM3DcYerj
/Z5XMs70omNastGJRvU4Zcym6rVCL7hHvtnb3fle0ggJdvc5gJoYEI/c4XE1gwuq
4mP7lFfi8QayNC6Qnd1W9Ed/qc4P1BE+CQ0QpeM+q1yiCqp4wB/g+C1TYydXKbIv
YtnlqLeZ8Nj0ZOMd7XXIF7KKXhf7StGUTmfyheY6UiHD6cVIpBzd2kgtlFQih182
5cpWBz71//OFv5YSRv+GGG6rdWa0UjFxhCXhHKJR/hjj5aHygnMdGP55VvSJahYu
s3K+dEzMmrqWqeHc7wJehLq/x7aJLmbRRERLuTJJHtAcNWMjW3IrRz265+g6Vt/1
FridGy2OC28ttluGhgpXW507zG7Nzp6Kl2QFs+Vtxj6aT39GKuxDfkKE7+uVe+Ls
PrpxVFtmXcHl5CEaDuxqNu1Xgu3Hj+Aqf0tUWDSt1GuB/CapaUWha8qErSs0PKWv
7JbVEq9bIFgI2PN/937sfs/kURMsH3j+T0u/jNChFE/jmugaEtF4NIgJZmhugiti
4VDBaDQLmnENAsMD6qy/KEW2ddJ9LXsKLZz6aOdqFRXnWEm3FjAnypFdv9SMYfsW
f+nDJJcdy71l6DlTom/8OtJbxgtPKw1NcM/4/jTqf2QPhRI8Od1jDNYqtHyQn6G4
LaDoNd1Q12JbynKrtYqx5w==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JSrfJLMzqDycbX+r1R4O+92eg386+sSf3c+r0AdM+uZvwV2yA/Sf2ADaAOVnQ3XA
nSmTquOX6hzMOSU4NvE94B2D0WTAD7cLecnntuP1QwRhyN8LnxerJ0WVzOhCxw7Y
ej02RZO6Z12SOQpnsXLG++/kX9RWSwlCoEqzwQ8jFiyiFE8mHscmgH1l07f3Ct4a
9BXly0P/4TrGF0Vz/s61a7TnJwWIwTnF/DvwyyQrD6r4G/0iEHcvyKE0Wd07cr6C
F9kAadcdKQ5KepHSNMeb+JVAbk2ArhmiXHm+LOin2E5Q3rltwSW+X6x9+gKCxSWk
ZxttLkHOIbzolssHW/eO+g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2016 )
`pragma protect data_block
LLXRqGrUuLQwaXca1fO/Rt7MUiMzlj5rVsdFbkaHcKuMP9Idz7HMNmriqvDuvVoQ
g+U+k0murjqUi9IIjEp6+qn91u5UsNV2MMCj5Pe8sKDnT3/4oTEtpG2MkgMk0Mor
k/Baj9BCLB7NCQBZ5nw6ju6+aCXqUiViOIW/pQ69ISdRojquGmzkTAEbN8UGx1c9
Oam+slS9IdYadlccvTz4peCvwrH28PAc7tU0tS59JQIBuTNhTX5qKiIS8MLgqHAg
cfv2FtrqQLA4BXeuHTXUD4IzXRSD+gNh6jtfkmAL/sUc1g7awxcJd5ZKSC6aH9DH
emEBKzlNlAMkJE4dfCrFupyJF6z1Sy18RLyKMwD6Z1wfii/fjD8x6aJrDu+lmo1N
pj5nMxNctx6miUuOjw5uOarTjekJmRS/5SfXUxj2g0Mcm+yVUBo4ewojjVXqsAqr
QTJr7w9kESmYHD89axIEiNR9Mptq3/9rY74viPjoouITESD9A9ly89uJRlvXpmpm
I3ythDwg/+7hrsWrvPVS7+OfuaXqWxI9hSF0FylqUfnGbJZRbnaNwtDFtiK5VBi1
PDg35quJKX7l5TU5m4gnfBPjG2Jksbv++tYCKACFjc54SLCsIhO0x8Dl/D4L9EgO
8jc++yGHjj0hW3vvY6wV+IVqWUrKur5Gj8kNO5Kj62h0hKoefNX1kZsC+brE22wX
tvf334mX7l2PnGYwi1kN1mP05/cM+A/ubT4RghzW3XH/Y00aECieH9IlV8/uUqdt
69OFF2Mtl/TXrCuKyjHBMhFitzdGYMzAtXF0t9KDQtXasFfCXp1oII1ikyHcZoY3
XBCeFNJBz2VLmU8AU1oqlNS1RCiIX/jWzbOenvMqxxY7KtpHdQ5ZEwYwweOUhbT5
uLD0KKB0WEjRCnig0Lh2wagU+/sNyK5yW9YV8Kxb+8xHaE4xrjV4Cr6xhBMCa+8j
W366XWZAoItgWw0TFJShYdpVRcu9gc+DxHWX+lEZ/AK5DVvwSgg5C2R3HwlAkBIG
gdLhfYvyELTc3zrrqp0jtBSmjE8vQLEsnvp8QsB8tDhBgrz8vRYg8X2HTNm/Zam0
Hh0bPxNm3ZjNyRpxjI1YrKEMeHZ8u5vLSbyrzTN7niv+RKncTdMRSlwT1izQPoG2
VNSa/5C6JSlv2nw9WWV4wJkO53MDcvxvgOM7dNFP4WYlBDtBFR8g8C0HQomDCOqP
fJwSvZjgpmu1y9N8cUAqldWmmiQHHE5ig0vzYUVEB7nA8aESkTi+PE8wAGFh9xW9
bkSeBfSJghWtWEMsTp+aSIUBF6d69KuH07PqddPMi6GR2oUCS2govfCSrU2Bfkbm
3ntuz+ijCvcVQVzRQMC8Xne6XuX5QfZ726LBK6rm3hafooUGNWvhAj2tZCTHmIym
0HLN33lv+OybLHIW9mhA8emKdvXrY3tdtBo2N5hTuYMiB+vOluXzb30x36s+O97J
97prHgJNNibBBXUvOULKYPwWVPbrFSXDN/DQkOTbtRVbqzaYsQvjJab0jYwACmhT
idf8RVOCXzaw+BDdDgAWRGQXpJPpLMQPixlakOdbv9tg8X6HtvWRYbvsCXS9K4rj
RMBfkuiTQPir7ZY/WSPiRQPBJIwVfAdjMCMzp2BmO2CKRUI48cRsFFNSi3FbxbSm
wGJRE96K2xQNCTVRdVtWjb6aqOz4OZDAkSFpMjipObTK5E6Z2IuCw6sJmt3jIK/R
4P6LFCoKjkeUYqe2cJf2dDn19nXfW0jYV0j7GzBB5gaYPanqP3dXJHl3lLMLTQoR
0dOsFcf+fK36ec0v2DjN7hOEAL+NACbzHJgFcT7lBzLndxAH3pldfE75wSfV6zoY
+7/UibXwORhHSucLI3GQVTV6MWr0RhvqczpH+E0pPaOLVP7QT4eUpXKgdjCOLFg2
nNrYh6LSdGbl79iZKPQeuprF7ybGqeu03e2aepZK69hck4U6cAtT0JNAIIKJDUhz
5XFDI57aFdbjxYytAdcJjwoDXhumR0Qpm+zGHUElRnCiIx3EcjTt1ke4JiiboBUH
1wBTL56RQcwWQgXWsyK2LREn0LkET6EAe9oA3wSm1lSstMn79GeHzTRD1O7jVBC7
G6Pd8nNom6JleD34n/Ck2NAVoHF4vGZgO1m2c+e6RtaQTDcpqkbCEA4rdhvNd3D/
LFsYOJMyZnLdQYz2e4aEfoz2AmJy3uAM2V0wxEmo0D3LUWCgIqRnZoXc7LwzTVsa
JzmfzZInH20WJcNnwb3JaWMVA6KgE9KXN48MMaHVg66qugAFJgLav3irWXuG6L8l
sQWNZDa+Ah2GK9VrEvMC26/ndIhvSZLUAgN9k3PqommI5W3OSBRDaGtxYrA10wf0
yO5M0ctVUZkr4U9xkzM9uLGbGCxZiH7DiY2v1jJkoCkgjhW1CEIIci6KPPbKWhO3
ogYwEMjZMMKGdpwZIHGNUi17kL0pZa7xuL7mZyuwJGQK7VYRIU5E/kQ1fQeWvMqJ
wJQc/NTLi+L8y7ZPV8b4YMQxyipbUXiL1RLn6oj4JpWPecJhfHmALA1EexKuxau+
N+ClqHtoZagBUKU6GMq3znYGkr2jzJTUqMQg5zcnr4B0JWro37oY9VYdV+Ss81a0
lVWPObXOa7NED6BfYQMn5RH2m4pvOVuS/cXrYbe7y473F+jJM5phhNKbO/Y4FVTU
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SSl/KX/uRh2RqKT6Ber3h0t5DKGYESWc9zR7x38Rr0Zx9NO+oJuKEnhhQ/EAfBtw
Cr+QPXHqXg62IwgiMEb6SP8ePGMfbv3+RDsiPpOxwqbfFwoVXqDht5fsQA/p3+C7
xPlMFS6KilBbg6gb/pDJL/xWN41O7FPfGMvKFL45JoqcXnFlbIUVbHitwIXptdNp
0rhEi8bte2fSL92fXEsm4/TH3S1+SzTGWsLIT6xXbpe4VKYvnStOA+mG/ZvLQFDx
QF2aglCMox1q2XKpDt+7114ZJ8asXhckRTqUU6hHZjZoefD30ke/vcnFY17mjAlP
dl+l5+WJpssp2fJClTPK2g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10976 )
`pragma protect data_block
B6RsuDHqMw3vndOdmKovJq0GMIDntvVJRdppQN1IBCFtyVD5pCVWdiQlgugUyjJO
D4XhwR7DI0XDwLqu0ZoJGMhC1+D+xNwBjjJNhWo6BpvwMJHL/4wZCWmB+LkJdvF5
ACgliDF+bm7T4GAWABUDr6UIYZETLF59cCtn9MnXSxmqbL4S/29yAdegPCvmxSG2
yMRjjSKlxA39CQpvM/bCcSxB4+BtpwA4tvh7sUyQV7tOvwelUvcFDGxe3kxnEP38
iLVnmT75Ex+fBbeKcLZTeqG3DVy1t0IatkEa4P7y/qydxA7rcReB+hzNP1grqwbn
ad8veAWAnf9PVi7PFhP8S4a4gdqmf3AUKHTBDe66zqp93ag/HhuGA1I59uyQwSjI
5mFSnjm/cYziE+Ev34w4lsseSPxwtpdp+eNBu1w3VAC4ppJHQfzib1hG1euSUicu
MjpT7pXoCBYK/gXM4VTGGaBf71+mEYx03V3+tFzP8EseNMJxP3NTYhidOOebL3BT
j4pXhZDJtcg6pjqQwgEcdX5j5ejQINV6Cbj03TDeTks89UjyuzdBqrH8AhR+WgkC
oCgds6Hi5t3bsxt7ogKNpq5ExnqUwNRdGfmcCU4gjLTSHkIokphIRnr8ObEk01pu
z40Dd23t5pTmu13cHq+gh6UVMfh1or49g4/8SKddhdAkavFOXojrAcetdpxdg4X0
YAsDG0G2ePBiwkLgrPEy6czmaqisdquNwrTfFfKtk3QejWocUBF6fEXXXMT6NXoy
NljWCapJtHK4iD3DjiKtmkbOKL/jxsdjS9K844h01kZ9rTPMNUG28bj/eYzS4LX5
OFH2b+uMXcKOJqVGpgzQfpDdEFgTxu5zB8+ZX/z7hQ/j19bgugRAlEoGNuzV2kCc
Z/cN2DQ8xF/sKmErWHYTj6zVKEqEDjTmVbuAlPrreMh+QqfKIkfd2zTtH7JsU5JM
MbdvfqURXBUZ1gwEjXY4zN8VLdt99zXZJuzMHaJnIzkW/l9srWY1/Wxq7gBb5Sjd
AIdaY+wNlefVpMbMqp44+Q4zoTUbQg9TsGQviEqlOD00RD0FhR2/8NHvWMOKn/oU
ASzM0gCLghTFG1ylqAH0koftF5oMRz4qJLLzb8hC1jXMPB/iXW+MGJPLzM1QmVUc
kgXYf7C9lJkVzA4xx7qSoeDnefN05qzRvRAPwEKtxIEwrhg9WYzbZQ8gzDC6tIKr
3HWwEOcr5zfhiRZleDjL5GB5nqGPgNfFqyQTv8L8rHtYICMn5H3qR84ApxZKKG+x
ny2rBXtl34CLhqS/Jfbz751vyjWVtx9rKbo/C6REXjc8w+odSYie9CnRMHP2E4bQ
3GDgXKF93ZDkZ3IL+n30bW/Y4oCFXmDmDvwOHjngmAFkxmlv8wAuiE4HUHOWJLU8
tC8/1AnR4/qLHjdv5OXnA5g2AVcsLuOrR5EmbWXeBAp7FMs86CwBLSarNYXbVvQ8
NzAhVt+UVSFiowenb7nHd10OGhEQn0HUV+ewte82d1z1GN2h7Yk7oLUeE/2mKBfO
la1Wu5C4FSGOPxeCf2RnWFkFBrQz+3JQHNH8DuTfDtE4BXdGkVfNMrkg+nHWlg/M
9zMOAC51ZfZmaXaAAr8WHW9Jfwi13AWYXZRw/fJfH3G4El02m6Sj5zQpL5UL7c6W
P9ZD3h7lAu6G+hGNp9MkO/LxY+ggSBOt+ioXoVYG9Wg/xUHQgLWVZOEZWVJ7RjTF
AX/afnDdJnzVVV27z2y1WEovNyaVburRc0kBF5XbU8Hz48jc+iZDYRyOKjq6mP4i
Fsjt2lW65KjSeG+XkssqNH8NTlwt0E6hwHQABKmuHCJsLR4laWyxOq+XrSfbJ31V
QbgEy8pMFr5+yqoiYAT6EtpPP7f9eWpmCfgGAm/9y5my+Za770KLaIJpG6EvqwCW
3QbfaNmAstqDCh+meTqzp2KlWN9WKHk37Dv3h/b36FM2KJaYetj3UIgIX0cXTwmi
ZKf7BqBDAa1mF5sYESj33gdrFJKa+gEIxIQ/amXUjNavtn1/Hub97uC22gpCgLv1
JxZ6hA6tq/t0S8eSrZqa0GpVvTEloA6MDRwu6aQI+7+cVLmEonSetYF4m+HnWVAZ
w7127tHoRgrWPBlK3AV4bydYbufvodG8ZbftTUCtciKi3RejizW0RGsKuaXqfLjT
LzZcDHYSoe1YFIuMQ7zqfsjTHHfN3Fax8wZ7UUKnUwFz1xK8v4b6K5h03EQX55wV
ITpitKkPJevqy4DGLdhulPtKC+XxNXdLGjsKXgKwiBuOhtJVMPjpBGqluVpfIbXZ
9GvCo3mYFK2cPYqrHSVESXtI7cp65HeA3BLQb8zcKd0xUCm0SJrQKruD68JcfbyK
XT5Qm3y8bRW+mAXcbBupQLUU8N18ZCtsE/iPfPMG9l3pjt1WYky7RCnSYMYKwU+a
kGrDDr8oM0m4b74zt2+bZ+fenY9mP6CWJQyA47Fv2M06dFmjkOmz/0FBaZEjLUWt
dciE9xUS6y7lnWNm7FunUB4xSut0S1M74bS8lmamk/Qla18BwDUt2hryxCf4oXqU
RLOk/x+rxYZ0LvqKqnUYWkFCiW8HoTe327U5yIA5p1pBraw8wWquAqlB1Qy4zy4T
sQEemLDY+wH/io6R9Sjdi1wBfby+xApAywWoLFrgk2mxrnb32m3RrQy+V+OSZh7Z
UqXgJeElSEJ99kPGD3E2y6XLS1XEGyz+JHQIQg1d9gKQcNPCClly7piEi5dw7Iht
01qlWznQBK0R8vhBj7N60JkEaRa0K8yASXu0t+D33zFFC174Quxi6EUo8PC8eUVB
FxmgOK7vpsWo2MHmKV15dzX6aVHkb7UR8QkNkwOd/Mn07mJhwsXEHNG+eAaBf6lc
iodq//6AJTKGZYvj7Xv9aJQW/nX5mIMIKt0QX1nsCyJjOxqmf6GHgczlaEd6XWnU
Fb3d5RBeRis0qjdC6DH1zCV6rXzujg/SHbQkzZxlb3nKq9XK25ubg37Gn4Kn8VnP
rSZvvge8zze3pLG5SxO0r4sy25svklpSl8o920XfrFi8Qu/ONsa0UoJXy5VwjluJ
izi6dwcEYs804/1LWFbeCsMF3fNENV9a8P/5H5vu7n92OYxqXvQrasAadQ01VuwG
0RyTUT+BiEW7OCDOjG68eiWrFAzRNIQlctz3Gz02dycLvE3uAvLqtkTAyzDqzokr
3jGjHEuB8xEKXRI8Pv8RRmOfHQayT/8yVq8eAoogQT/+zg8irWQtzmUgOnNA2/a8
WuZRu5C7zlJcaApRT4Rfr11anmQvrTbezYEonglwEAoGgRQx0qEscSWeexwhjrvr
udrBnFMtxDGuTMoNMqElZjGvoHBUGtup+YhlFWtbrmPlUxA/vN1G62pqyqQ6wRQt
IBfWTwTjweRjLdYYy8+xANEPFD2KAnCs3unQ4WiZHQI2TsLBTOC4y+gw9t2naCDm
UKehisd4r2osq1SiF7OxBh7HRXl70V/dzyrwDURfKzfDKkGnjqsT03WVgDHRAnpD
JNYbQ0WIWv4n215HANRk7lswe1sjwZBzDO1gGQJLnlJoTt0ptuYsFc8+SJNH+/Wg
11B6hsYQWN6Yv+uwhx2I3tGqmU/hQlROV84a2T91pM8/WQXEsQgBra+iuUGIv8Xb
mxvIvegJvoakaEcGIKq9uVJNJeMFJgvclIc14Zg0fNPNuNDZJM9oqiQfz8qiZkI8
/fJdMdwQp079lbJyB4g+SZQ55UQojmso//ymiCx0gHD1GODrbj5eRydrJMuZY3qu
hk0/DJW5PjLXXiJbLzflnCJStBmNJHOfg63ugSHBJOtpOyQJmFJvs1I/w2GjLsif
Pf8mUOIWrbgdbikPjZK09NYcoWoUtutwembz9y0qN/gSfri6afnFv6YOeUt1DY2V
bIC1rKGSbjo7aQsXcVUAEUkliPkIfdg2EL0Egb5ixDFom91VORMH8ufM8jY9QOKC
x+0lZGo2zsUkEr20TnOkO0+3i20uaqu7MlJhI6utOOdYN6mdn1qDErEH4QE/f6H9
GKn7lowaa1MfJsBWHciQrp5y1qXA3lKiY1rDuwdc6P8Ct8WMg4kx2p1C/gbpEVPz
tATRND5Unw4T7QTSp4zTiCdHqBkyC5WjL9acPVKaGmR/MHOTht6xvIxdxDtcbjUX
D6U5WzwMCI4U1SzCV041DKVIx9H/OId8iesM9JmTEsaDCqo3VWcE9eh548qnjX9Y
dDIhBrcqdPWAQwkVJWZioKUt9DE9IAUBv6zuYhHdxlp6kQY9HvUzDMvbZ/gF1n6w
N1+5mP3lkTT3xEBrqw7L6y5EE8YhHcXT3EwpUPBteOY+XyK+Pu1ts025Mfm+zBsp
I3IrA0uIaVHhVxEjt91piDf5vbdFN572iRsEYFF8U14Y3+2mi620mbhyc08lbMBJ
UpYfhvkXgOEMMG6Y+eGCXsMxbs7nlm46mZty0xVCBdANFJZB7v1WgIkg8k0GgzBh
oyfU/f+RazYwOb7/r0Bqv7ajquxQnEUI5oEtj3mRnThyzVJhvacUD/ifNVLalf2e
numOv1LnfUx8QxXAdnyBwNEZ67cmq6e4GK8eLmJFDuKAX/uzGQXIKQciItPvue3D
IHYKij3yBqj0gKlakJzCJgJd0E0NZXFbJrQ1Xn+g+BvoZ/1WR9wXhU9mjpDjYzhi
PGvYLCs337xHPtRfciNWBEOKQtveIrc5lXu8Q8EEcgLcYVhwmySpK02XIDwnVyhz
IlqNdO6+t9AwFOcW5wi5PPc+Ekl+dDFFKCHK3j78QfTwoMq0/FfzPhrRcjQmEuc9
owOLG46w8Hs6Dq6yAtTGwAkJnx3TFAuoBBSeq+Q+UWvOSzrmEOK3JU3tA0iOtWby
hVdYwvnhXWm9wSmYXA6HBIeK4iuddbzdMOVZpk/++fGq/On78mHdZnlTxcQ/U9/M
43FyL8s62zL18GzxT5yXXA9DfsxShzl6TWoO9D7sJugJFr+y1hVTYGhc+BP27I7O
g+zDOgB5b9M//FW3L94emt9ugelfqhJ4KHeBf/yndBpHm6+HHtanxILNUrq3Za9H
W9qEPbjes9n8pu0sXErqmEU+w3xUSEkE2b+w38WkE54OV98yY9idgAG6Iotcl62Q
aQVDuczFb+CV8tnnhOqFMrK2UN+fqgfom7bEYXsimXcWRSmCWoYPuvotRk5RRY/C
yttGpmNhaW+6hCqHJujCol4a+OdMztjCmDIvT3/pXfy2rOPJx9CzhHzx4TlNFenB
hSSzVN0DED95jGTmyy8H8JIDmqdvolqSczzlfGJ/ZAz8sMAYBC3DbN7Ju7ESL/Fj
7Wrzn/EE4yTHuBO+AVPJ1wy34HisHQecrgoDysi4jpstjJbHqKiA7Xlm1eM9PW6N
JCD5T/sgfnHovEPbgiCl2Uh2rYdIj9tE9SJ8crOadUQbtEKm7KfnNdoYDa6YhcK6
m4IiYUYiBhJG39xdCn/tWZga3Q4RQlbIaBwJvz/PL51CooWZoY/NFsFxPbJCukno
24ZA4IMCOQoWfz19iUO1omrL+D0SuyQPQlryovhZfXXi+W2FVN0M5KiRXAmbO3qJ
F8tJGq8K/zCVy3vdjbZAqk1TFd9qv7p3zb6eevHA8AnxYyOJrazs96X66v+yKQ8I
LSqmxWX0Mhh4yhjMW8lO5odXxg1HhePG4LBwnxhfwn60zA/N1rO/QUy5sma5NDY1
1UrUwT97ARyWsMrkU2I0WIH3s/k/DnltchFn6/+xc3De1CTfpKwhZ+ud9lhJf52h
rKDeBUsQcL/9bL07YPEfOLVPNay5Ma8mBwqMeY3mgXC3JWpPUZRm0vdZFRCmcD6A
c1++ahFsPx/jwX7RNqs6/tXoV4YSawc0DKTGvmkUlmTe4WQ7J0Kqhr6A0Vg6C39M
SeS3DQZ9nXKwm2M6fm/metR+MArPga4yddsV4ri5cjVtTaKoj4/Cp8KY7Un5pcop
SHNLQrHyW2Evw8K+dlftx8p1dm9ctCyrCR+SIbYcGYMsmvnTW6ctQ6KYO4yhd2xo
YBqnRjwzla73sQvmmQoRCUX854cDfily6uzZq3iqkQhXd8LZDhfRsxjSHOWi5Yuz
hAgQLW/E168P2eV8Sin2JS2YEZDZth81LNMAY3MLJpniv2M3tDLV2t8H0X1X84dS
LZEh/m2R2mlcZ5xtLz6eoW3ntjcTMp4EFqPfoPtVVd8MqexNMSbf9309sA6f1icC
soBMguG1NKECeOAi8PyYBUWLQut/L6OnlpIvfc498cfYM/egJ3ChVyimqBM5Z90l
iPA5M8YzBmeuA3zFRo+OuS1UbiMF/4PCseVTYJ9pGDs/T815G8KnkRKnkxrVanto
HziCNsXISLQTobbSAvZuMrqanozlFDdLbLxWzy6UWL+BCah4a3rgud10kOaASSjg
FVT3YTz87EBuJlx0gmlvaze/cCt53iHAeMVJVf4fAa3jaQ3QdZeQqw1I8tb/v5Of
rBjoUEV6bLQ7FzVd/mrGSMe/9HfiO3agC3BKkxtagiBnacIF6niBMRS3R89q1PF+
eEyTS0NBgDQnl843JSnyUGp83o4nC4XkOOOGk7JbJl4TeOF1bWnUNj3oVOyiLkgl
utUu0f4/IGqLixMx19wI4LsSBqhjGBC6HcLcwPpqJrsHieRjRJ+HWAidI8okD04O
V9RngBTP68GU3BUb82UsBG8+AxJznD7EsEJnZoJEeuMVDIvsSgiyF0rLYjkIRgkN
p7huQhDMHo9iQh0LjY/uydpt6Sa9NUYK+NzSBYGxhNSNNnCp7llFT8gP3V8EYAt/
BPeJUqCYHwxQJQOS5VOaneiNggH82ztlgRiekm3oJKA4LphR3vpeUqrABlLE3cDV
LO/VKMAY4y8lxWzAui5kDKIsPCDkFPSexZQ5Co1mMWtbruMu0ou92GHScx04SYQg
9b27craiTO2uPan+KyCrtr9ye1oj/v2npi/G0HS0tGPnzlUrqb3KOcRx7VEs7eZy
UKyFFPoYLshSf57qAd1oGX8v+A6qOlVMt9AyMu4tukSyvXTbZ+0sTDxNIBOwKDIr
sl5sJnFF8D6sfi8D0RVJQsWDT5x0VCFUMeEUeY8re8WNJCsd/Ev9HKKJuXJov7Jg
OTbKF5mkDKWxP8g/PcTrSqQABof4Hh+dL97g8sacyF5+6El4SWy17MBeOEKFDa1X
8XplXUEoloQC9bO0Z6bA6973uKmCl7m3uPC1WvWc7DgKZdo9I1wdLQcfR2Sq9UAa
E7Idis+RPsP7YOU2msl/e14stZAUbLJ9GOacRIonGN9UgcsLXtZ0a9Zvy+FjTvkO
zTpZq/Ux2iwORBLMY5N8Siq2PnMZ/28/JnRr7zcBQdt2ILFiJq2lWq8xhSS2isWp
srUA0OIvUgOXVbTjXH5tnsH9BrC/ecqG0Hd1IY/YRm8vZkt3+nNNTbMpaG1PDxQH
kxXFuR4+zljGwHOxb2aUZGFjNQVwoiMYFt08QHGvGRc+C6zLGKhQwjdJ7JFUTqHO
Y2NK4idgFKuGZCeMeELvcI/sPTsKzfOjyRmJi7zmyqemwXK2fO3ru1o4Fai41lh9
lDkczozPbgHAZ1P8UQkmaPS25VHuqQq9UHG/okeURXeuVccbNVIzFgVELL0D2h3b
jw05jLkKIHfU93JXle727OsgeAYzNYjARSo/96vWQhaA6tlllzaJ4NjQggSO/FlQ
zo/EczIXv9E7e2c/OuxEeTMhKWTnNCEsWVtyTIz4AJAO79W0dO5DyAl4hE397Fws
qzUvwe4Vn/S8lLOtknarcDHSw6LtT5ZDBLUG5qYTMNoTgRk4IFqAF4+fVaMiAST0
nv+3I45jBT4qyFGr0sAQE8vYRRBfEriQIRpn3FoVWqfDToPUhBFPfWqdhuHgU8O+
OO2/MmpxBySbEsZ+6eHibedCvzrhMmfj+B+msnbWfSLhl+MYIr5zyJz6tDP3cqTD
MSrAZuwTBjpWiI6al7Npzan8m9zxBf6AJVC584m/lyPD/qwLPOD7ydy53YhdcWRn
LW1FcXBMkExXKyXA7SOoEoNy+2rrTsDmIB9PaF9MxJR4UGhFYk5NQsWxIMoG5Z1T
6FR4YPdmcokvzeHpU3CQarDES0lZyBap0k2RFd9RwWLcIA4Vdc5ft3M2+/+hugTg
S9ZUnmgu1H/pZraoU2m5DF3BDI5wuu/Csqcr5uEq+HtIvw4w/8cZI8tCbmWjeCR8
eTD1NOOlISP4dExP7F6dSb9dv9r5TFOGqh2ji4Hh5GvAC3obzjrrw8sgHYxrbiYh
DwF65WdabiQjeXoZe2Bm78qnTLKTmF+BuMH/A3aYMGw8gDV9Hb6QNFavi6KqLjWI
US/JGHPbxtv7CfBqIg+PpX+ihPuORgaH41Gw5MWKKzwJm+CxhNVmliFvtT5noKh0
+T41Hd9h0gl6I4x8lb4GV0ZDhCO9w13V8FBni5HI+YBQnBDNPiJOu8kktnzFpG+d
5EWmyULym+oYg7tbKkYVmHhXDhJ37T11dh0nNmRE6Es8Y0d6hEuXVCPVtZJZdg5S
LrL9ZWOkBykS1eT5rj1oJHgFp3zFY1TO2PHCu4tbLkcCuq4I+NlVM5q4ida/JR6e
Lo7c2CwLjgKKfkefVUBd0jwhQId5M/gc2UaxNvipz6OusNX6WLv8QurLSGV41lQH
cyBn4AhycQbbas3AcFPm7gsYh2JSdgzoBYh0dvxPv8K1g34q8Oqk3v4guJh4YEh9
6c19sDVPmqVh5rU0X4SjW2Q94+0jsSPT1Ayc7xp5XWSFq95pSysg1yDzO6sZe1oj
a0WPkEG7IKOp8slLIe/XBWBjpfR+6knx1UfHHYEabvvk7+ttqFZpUX1m1KDKUFQG
bjGrGnuzofKcLQ2SjzwUNZgxx8DIK77YwEFQPpnrEAr5cUwV3Otnot1NMDCOOir/
xfOB9xMmebF0oxKL1eDZIRlwWcg0YZGCX4TeyO1GMFP/XOo3vF7fNjKT2b2mF03n
GxmHmizUqdTTBt3uqhmW3mZ2jUHZPsTB/kzAS35pZAHPltYRwPBqyNn97UAjl9m0
M3Omi08kKWFCktRt2FmJ2H9chNRDzA0WPHdPTFmFdxMsqfXUOk8Uqg35MynOkn+O
KRbyX2mindfEwcjfo4K7+SvLhfQ2d+ILGuFkV1szD2UzDkb83TbvJJ2C62Y6W1U7
wqC0ZNa/j74b8wPTBZ8BhlAKGiR9k549FDZgs31D2eoQZIr0RmPH4UzhE01+j1vy
yubEPOx+vrSxJeAC9K8eCMx96DbSZhPznEmT2YoGIKcDF5OsIgzrFlkOg+kwY5pE
CKsITWyllUHZiyRp/MBHV5rHgtdbEWUF9Xj0xuDxYxM/macvYUUmkMpC9fOSFOkX
DweOGxHyWqSCa6CW59VxdGPvrxUSN67+U1DjG046ntMP+VahmYVhTgJYli59kTCW
s0XzXPp2rmWoL6ZSd165lrFAwGAxpSTwpUdsbTtS9s8tRLzdcG57xLtKuGoeJbNR
t6p9usJOV2QYr5dyme9xtLSTu6eMJuP643l8cj4BXhVf58CPiR3ISIhhTDBN0g4G
clTB50hHsrD8/fZNibeMaRDr2nKtCHJ+6cjrELz/h+JBSHi0RdYEp/PJQIb8FxDf
vPoDRWWOz0GgeWFT877UIjPgI660R/EGta1bls4e0mj3KX3m2HWBhSibMyJuxVQj
M+/Z0Gd7sQ8b/jGq+e29oSz4iD55bTxiWjmdJOhBP30SRJv98dK+aTL/AF3Xam4h
Apit5/Hh0GwCv5fdjahNvlTekgOByyqM78PuDFHSFtrvm1JSzJ2NvkDveP492CJ0
6hWfUTDm/wQov1nQ9qd530hCqM9SwJt43O9DUeZSBmSEL8ROomUyjjIhzMhKJzkh
oofgWUn4SzXtWwU/ZNCTqgwn+EKHzZ1f3iFs2UE3QaQcyIICim6Us71f1y+22txP
uS/VcrjTPkNpFkAIGCpeqB5VsTaF81joPdhnNMninqrI4CngSxJYN6Ir6SGPsDY/
wHTjMyBew/HRVEafDml/Zg2JJ0Ry2LYIlRVoK3w4m2Glifim3G/5BVQTYz3mYxYR
wasLdtD0Pb1Ew4zFmuMlGPkEBYzru3YnDqsTgNJDA6pSTyeTNr3Zh90FAdWSIGFx
Thu3CA6J+nDMa+L9jgK7LFHcQnvz4RzCL4kST0WQa5fFksmW+Jo35+esgoK0u/cS
lholmaytl1aKsLrggKBkygxS9cO5ykse5a9JnLCufkEwlErPHP9Xgsm7Ym3g3/u3
eNZyAYW1RBqryEeXZZ+9bDltQAeR4Q5aUTIX7hU3RmCWcYByO/xgv6/+KbyKxJhU
TmsJypelp3sq1hQDKkw69l7iPztcaGEz+M25s3auHElWKJ30dBJ78zUUYbItzi5Y
UVW0ywhr7uaVrypL9fDPcyyy/G/4FYfj4r1u2VSAww1SEiFZDUbwAEqVq3mCpZXN
npjMbB0Ws/rDa+aPsiOZoU4ICROXxmsbUDqbo3aj8Sq/KZDvdTBXxTyqVjD1rS3W
WuMYtkipDGnAM8e1iZFDQITKaBHgZHtSUV1j0SJWpIwLkBX4Ensn7eylIgLjwy3H
VpnV2Y6baaorZg09eiwrWpwx4+rgW76ZioFo6zGEpQyWfJ9awGNduJbGqRphxuLf
L9Ji0Mekhil7rAwYbRPTTFcxMv7AmC0TRxRmGkQyXN/UVAduukYjGor/8NWkf5ED
CEbMF0kTGZXUqtjuvNqnQepBzp1yO0+OYhqpVB+DzVrBDbHbplYP97V8yY3N0oUa
IuEYMbhwKVyszXDj7+NUNCYHnwCcg2XBosK/687Jc5lOIjOWbkUWvubWo6NHP6i4
s8+6SD5mYTNsOyeZVySQBly74210KlZogWUDX7goRK9nkTGA7wxMaEdoRzuKlevL
NETXAvUTYguS8cEs8Cr5qcSHj7+Z7g+XEzF7Vl5IB/PwsFz9t4QuCArvJH4zi535
sYhEKBekGfbEuJ4sRjf9QYYvDHNhb1npk/pG2JI5vgjxaoG4K0e21nfJQQEf6wzi
IMU+03SJ5oJ+zYg/4Ch98MiJ5dI9fbEaq5fe48qr9q6BhVuNHK+UoPzFwoFoGFqx
mGPNG/Ez1bFlPmXtqTNVSHUSQ215vYj4wTPdfPCvCFtwqhq6IFCO/VcoxHzBQFJz
paNkqO2eZLZqIDJ/2wnClxAYi7xUcIMVl0M+jkyJvYTOOmFJjniITAxyhHBRy5pT
+x94RNsVppPV8uAqCWmxmSGuuNFnHU05N6L7A66gbWMafQFHrG2wYgvb8d7kdfXp
YtRtw9qusgKR+YfhgezWIcqhDh+0aTBgOgfzXJ5WFoXh/9Ahy/DRojFj8Z+NnfUY
KXbhrVZI4CPzyFOakGBok5KbYxlgDrTtNKUnxXPxr43u+4/KZjWov6d+Cd3div6U
xF41GmcoT45nUR8sEizgH4SilNShJPpZO3EHHt0DOCHwtslgtD7sASykOc820HlD
n8T63DuB863pqK5nRxdYS9c4W/88bUCAicxzVqPGSQZbgnxIvlWteoRGdBIb0ug9
+TSvGK/5Ny9ICpN+rxeLN9c04AiSD6U+v88AtYNXCoSVX6PwTIF/f4eLqd7y7vG+
DP3mcyC2oB99SlxnvsFMlvz3L8uZG1berR0mnJxitTJ8LPBJzeJur6HSj5xYFq2t
Zsr2PQbWWpzQ0oLjyVj7NJdPES/o3T5M6nFT0xV/7/3tV7QdYMjz8qoahjT9aub9
XAHQ1yhXlCAO/WS67w5LKlz2LSBnajCIRhgZntYzvvIeDeTD8YQrOzMdzKVhPW+G
Q13lipcbcmaKXqyPnWlDkjNe5s1VmbjMbg18AdBhlnNPN6xXWN8K5wtkUc20TS6u
1z5toi5tBOMQFRZWDiWSz6OeYO9zpTD5LBOUFxXccfi0I6MRIDD3xaRC++GGbSBx
bXo8t4azaw1LXszF5w83PnIae3aZmaYiPJxASCC1rY89rI/m5+6PnhVjOj+PyCG6
yaaTM8BX6UnrC2Vv3+obIyJWRlzlfuPsXLAhLIyb13Nk4GrGpzcROCvkp/m42v/5
EAhi1As3eKahOwV2r7EmsXe4EWzK6XZ9+eY8nlNctci54Y0XT33JNjnyOUktX7dh
NQQwhmN+v7N3Eqh6p8ht5Lc0G77TkJ/bGOkPN7zTf6UsvcMlxwRqY2dy4H8KjWTf
QiGaPDILDtbjc+MDzQ+KULvPINXeHzItP2AUxmL5SQSqscrzOpO14kxgZGAvfuE6
RXMruaHKsEmTPg+toN6fhZtcpIEE2ENUD6DAHb/1Q0BuA3MR+rrpKcdZRVnG4FPJ
Wh3AE1NifUntl2+w/8z8vkNiCZW91B/kySY8qba2DZmw2CT6k5e9ZgcYW6Soc67u
q45nUEYG3VcYSVSK6+QBIlOKQC+rsa4qTA8PE/RTD/cRng49xvreWFSjPxnd3Yyl
fjuIPzfpDaqw/VMQ+CPQ6dtcg11cU7YBwiiffbf40rlD0R9f1IfjSPdNj9sn7F8N
OqyZgzmpXwPBLDRqI5r4ir1r0c1v3mcAai638AM1c/j6LZhzeMn8av3GtFnSCBGc
OfLqSWpyXcXf/1ADUYtTFpT7RiWnhNb5/DvXp0geMPHA2NR3udRcbboWQfWl5Omo
yLe05hK8smfB2vKliQKqnOaNHDbmrVy2f7rU2KVG7YV07wFA2zCzvBb1JeCKfrQB
KGFwJ/Q71Y38HfbftrPMjdIFBJCvk30KWlaMbYPwN3rtw9qHK/1ShYyB51qACrh5
iENthcd5vPVDbEUSM/mqpCIG1gZnTUMIUeVVv6xDaeCy+LNonVSuCUpxKFU98faL
ZfksyUpU0vDvBEqjVUmEK9znVFw9orJJjJKDijmSA8oC+yDt8YnWpa22GJJFzN5f
0nwQHSMpawrnzJZw3Uf2incHPtqR8vfOf4s+Bxlyf0N1PmYoZRcMTZvcAp8HW+qj
PicSTw7VPElISR4f5P0WUgYdIPGasOURi/TVNdLZgB/gkb5qHe6Bko1fW4oZ9oHP
+0PaRlf7jM6KVq9m5hFBxws7qb+Gln8qZZ0YlZYhc8Q6tPLJ7ax4Mn65aVn9+O+q
9VqNikqt15N3dwElwrSTtKU+a7q6NFRRjaSU/Lu+PtGiy9yO2b0YvAIe2BSODDHP
TP5N07Z7/uUHAxuijiY90J2eEnhJ/4phNpiy6vg2MVb4Ily6fEc//lLIRC2GN5Q+
MH30MkKFUULdAzzELyCyyDl9rKJtUzdiQftRENljIwS6cJe+uJkiHnaE4pkvg84b
sHyOjpGkLpOIkBwp29j9oJHFQWE53vjsDnkvZaRMcVqJf3SIm/1dumTqycjbS8rn
uYeigMG8cHcq4bUDz+U0t3bM7BD0ERjHUzCUYXCtynmhcGnrX4bujtBBuPpz8C2x
lSXlUpNtIGBM9qgWI/C5SQvCjgikMePup6GqCT62CAHprkMl5ww50RLcqrVQbkLn
1VhBP5jLoONP9P/kiqtBXDTOTr0mQzPHWWs/Bn/iVIyc7H4nvnE/0yCj2YDNyN0f
5Juvc6Bf5ctKBSpFGWGJM4KcQ/fouZoWKTjSxrTIrrOwe68OmB40doobG9m2GFq6
LWQ6yungibYKL4+3+bad5B5B0ADEkKPOqrUc+6hQMRMcbtSF3AKG/KjBpJgKWAxp
VIw8HQrjHVAHUiRa81Kdu3Ugxfi/bdKU0mZM12wuL48EkfSHgb742JiSrno/IrIz
UU8Ya6JplEq1xJtnWBdxTTuX9P8NBqg7mCLWw3q7hd5HS+7zmaXwT3IYa/WbeJEf
LeRtlMlaRo8dR5FOHXqUZ7z17pu+DCXleQFuOSRdGXGXXMFkCw96tXU63XKZUmi8
JwOlJR3Xp7cNCOTxsl0ny1aePwGbOIa0jde74gIiPn2p+h3FeohDEi6tImzjAs1x
oTalzB6odjE4LFhSE9O9uWJep5yzOkAZZq9s1KcJM5hAurBSGL4aI1d21pWqOvJ6
pwxUjjPmAYe7B4OVleQLiiscwf9mu/NkCyWmW5/oJqLDbdBDqgb/Z9MspYRve9ls
lo4fZX0PNnKrK4JuY85Z+MAJ+WFWcggqCG7JexPw/fm4ki1gWYa6jRWe3wNRa9pn
Bg9hDTfrpF+NJAhzgDg4mMRobe6cW2gWGvu+y7MjYJEdvFJ3F9MphWsAonRlKLmQ
xNmc9mMpSkpYngMCKxhQ2A/gnHF8bcBKU+qxdNhboazx8Wv2+RGz4zWNxk2f/tAk
hg55VHo5yiQJ3vPu4piluJfHKoKA4YHTBFePbVigRjcid6PWSQgKppWmu426cuUy
JFhdGF4kcB0z7I2ZO5Mt1g9b1Em/4rQa5ri4W57SwYohwn6Zg0Czzs4+3GUKsFka
uTqWajFLqsfF91FCJZFHZh+iHN7Ct5TGw1w1a3BIzCWjwSD7FSlfgYYxwPs94W0u
KR+0+a/rRgHBtlf/CVgzRXwfvhJ4fy0MH9AJeyEWE8alfZgFZyu6jIE6a0IoeL8y
95zRQz1A2JmT1tTTVBboAnXYV2pNKsd74mxmdhZnPq9EVy5L3I21ryEmLmU4IbXH
jn1T3qg7UWzo/8AFWTtvQOYUki6OOuzC5obRWZEcMkLf21Yz58yNwlan+973gSRK
TC9WcNcnsVPua1FV2M0ZvT8/OjR2GsP5MTDwIFA3A90=
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bn1iOppJBLhtddAIYPvyaJagdfrOLe4k2gxH0h76fMs1xNFldh5hMK70lK0696Nk
/EszVOc1diUc0R3iOVTl89++FZz9E1mtzu+1j+ziey8riu8/vJFReyt5XcTlmXk6
5h9ZKV1qazOrkj94f2HvTeVMJWnV8Mcq0aNKDwQZnzh3eYihq20qKSHvljrWAJiD
fxOQDGmMl95YM3BQoJPNLS/CAW++xWyKeThG8yVl7HRkQavKYazf48HZnVL+Rig9
AOgRD4qNH8KraBRbgib9gNF7SghCmqzyvrU/JUkF6a/2NZh1AKqeZhwMt3E5IAG+
LP82fHu4FC1cVydnoq7WeA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5040 )
`pragma protect data_block
mUwBB1WDKvfKhrtLPT2LGn3LFG7wmazuP+zOEMJYeyY6pM98dkvqdl9jZ6/rFm1h
WM9sbhoY/k1KMMEz8BZPFkx17/B+hEQwkZYAl2SVqz31oa7PpU4VHJWNBOGz545M
R3suqdei+zuHMO8NhyLSaTvcPWLoDVf90ZC6Z6F8WCx2vhzmDmuzCRHQj3qFSVeu
65T5JBcJCxyNPnkQY75kL5WbT3QIcu87K1Yaz3+qaK0XuP3q6IeIyv7klBM8QXff
HBnJWnYJOm2MipuNR9mCu/twgQn5E8VdVAtMbqv8cvT8mT77EPA7cnYyeTE7tlsr
4UB4sWrsnZMhhtBCwxx22o31x1Q+vNELxifncKp2gPhQhjAj7lAeOdPoR/+T7swz
3r9YUuJEnRO7ANKPJ1Apfr9jd/QKCaPzm7A+C/B9WGofgb1O2kvKUB/1vs1MS7T+
/QKytn6WHV6pEMrJuWAL+g6tltcc8ZlWKOJl04Jxs2IdVk+4menXZPM1P8bGKlif
J+l/thZi1l3mprXyYLJCn2AzpZH/ni3FHm+3/tW7NQDXVpFAawygntjb3Ay16GEj
AO1PUKGUemTXmjrINfnhb9bjKK2cFnVCQTCWy5ONvskr3hYHRnw3tcRwy5nPlVhU
NM4bqf5BcZcFOUYZyj8ORVPorck53YCbzcO+Tp8QDaIbcyjfL75b64snDgTg0TIP
Nhxa+jTnYM4s1ukL/+JEATc4BxSU/tASI2gwvGBC9pepD9B52LlBMaW7IBO/s6Fe
fLKZBClwJ8qRyMj4uPFqwLKFMECYH/+N/QRM2CxmTwBb1zQaer5vkREmZ9GBevAu
3DdX0+r1LpZdxJjPDIT4rTveq9r+pABABHeiDutwAEakFE0ttHUyRLZyJ8tGD0zz
t3D+FUdyw4Ay3Nh022D8vzdIbCq/hMULrtv9eMrfJnPIOilUjE/rP6r/NoW0Hj5L
izTks316jF9fmFO+B8hniueXpWPC4Ctr9pSY36MMLIaFvalrotwUAaBSM2deBPJ1
sEEYs1AA3912VmeuycI7yiPcI9GcIxp3RKKWXkYLHJcdAgr9BSeJYJPRtqmwkxio
GF0rsYGyKw1nCSpx8igpHqQ7ydeUfliChZ4zlHUyb499b8P+JnFkmhTCsYru2qgx
nRJYaWotKl4/WKKyui5f8YPs0FeKEqZfDgBgi0to4Qx8gSorot3mSy74IOhUvCsc
cQz/u7z0jxF0uzZjdqaCRqy3kuEoY7GIHEfPSAqkPTly5JZyZRMLGEddgclEJ/YK
0vjfoaR7TaD5qmJdqSgCNZRdUQwxeIJjZkHPSqZsMVWa6EMydohnOeVMEp4685bO
iGC6G1Z0SN5GfecH5OjFBIO4nMqlSX8uyuZ3ppkVa2HAlwnjSc6UIEZIHMUfYUMG
y7Uhuv54+PfuUBfClMDI1z8H0GAqyGf74/MDOV3gkMboTIoZ+AVrEFlRNopO1iOm
H8rIDeL7XPKkzeyIXIdJdZi0jIxaKdxa8HC/etI7ZqHLcrfELs/eKyQfaaaSxbgV
Q++PdK9jvduEtNiARHiX30fmsUZTQ36JQVr7AWfa39gly+pLHOMq5s1EKthlB7vK
0IIdmAq7rkRMV6MwUhaaMWDca5I26hIKztJ2tq5YKifLgHgotUIAIbIVqgpzkZ08
INjt9iPglWDgy8fVS3E/sZCwbJWPrfUuJqIQvpiBgvkRUZ3mGMxRYEn9mlDso/AA
tQ1EiL/PWxVa/Rlf/U9e4prxZjeDzxGlK1VlFWEDLFSY7rKtM1yiGiKxO267cVpc
RXwXC3gjJlU/FFz6z9Klxlu2jmMhXXv+JEP8pzXpFzFypaOfh2raK3pHxPpo6J/A
Tzn0Ef8ouTUKm5UM5Kyh9nE5TaU43t5fjxDjZbYX2utCy1IbFetsAb9AnmfiQuTb
qiVzRFetk6AJKsbABZXx8N4kixrcGg2f3ZaaAxWMlTFezk8eGuF29tfL2eu6z4Qi
01QCn3tGJS28IF1WK2bcPHDYV8NLCj3zftKwJaHAwLr1DWY07RLU9BIYWzSS6hug
y46Qzlqwv6DI6ZWxJsZpZIYsVdo5pEWqJKYr9BRKwsW2b2ZtwzS/a07jufWk/cGJ
HOdByqQu+1F8WqwvEgh12bkxNJC9myzg07P6x78JGfrMSnRVp0JnmGYrpneS+Vlj
11/xQw6R45g5u4g/uQI8vOIQH8Q/Y0u5HgD47dXXoc91+jKllGSA7qBv4CAsCZhV
0NKP6u/Ls3hmUFdFOmZ/D7GAAvVjXSxo8CmXR9EoRtuF8e7iHLvP4FBkol5Jieim
blhHV2Cnv8fQAOcjIup4I8ETwBeVJOtXT+DZHmN+SFsAa1ZtuE9W6hyonibHxl/+
Jlqyta6fLIfIeveZQtJVuBjd7r1N4QAmq/CgvOAcIz3ASsmNPE5mFmsuOL0UyIlK
pzYrYFR8h373M+Jmj3jH5kRPgZPpnIdpKn40oooDaiG55NKRIWBrAhMLmrGEGcEz
SgzAVpU/Ua2bKYidzXglVwrXXureZl4jOAxLJ45S0lxEtkNfpgzG2YMcEozfV0C6
IHYMeOPYmV+Uoa2Wb5DiN4fF7zeqBfN9q6rdbsIvPpSR/1aPC/Th/0GtMq3tWJTv
lZyDX0JBCgIZPbK+VDmRCj2v0/kdEfeOB4jvYPtasEGRsPORJFy2fpOICtgMJjmV
LJ5giJzG+lZY5J+zjuqwKrm/q4BXdWydvk5yGzuTTrIJdOcFWJwPp8b0hp433MEl
CodmRn3tYwdsvJTM3ep1aUrH9stYDof6QJ61rfvHUhfj3gqUYxUYIiYuYFdk80Y5
kUGuntHev35MU174uOSl+snPmB1I+AOI+pKxrZ2FavBVSl4wzCZm/v7jUqqR2Dl7
Xz89IzHFNeeHsdgU4kVGuTsStfbBU6A+FPHhubwa9pOPuq49hx/vifue1VnKuiMJ
tXq5fb3gQ41DHwJPO4KN7owNpk3AlfCRfddIZ3I0VanmVTkRZh+SlJUEQMInM5Ir
f47m+vgeuKio07739prZKpQkMVnjiJGi4s8pFTTsx9bc1hsI+jSThnSoDV3MXfmY
aUJQFVo5BTyNS6ISuaaOHMVDp7YTQMxdGq8orTeSjNaNrRDo9QvDs+uXxnoV0d3H
wGEod176OurlkxurpdG9m/jZsggszRpGFzyYE7gr+tD5MVOwRoDqd1iRemRDI5LT
5qYQ6JZ1HMNsqwKyj4H/VOXK1DxfS2vpEh1iJ7dFqdLB/M/X5xXxdeFczKMAhb8A
AhaAhnk7BPaL5avbm0csGXRfEBm20zfRvQN8BqpzyQXiwaondRKu0C4v7qyemBDt
9CBBzqtkAEiPMV+26dtjBOCcdHgVwOwyex9lXe3wPkHSehf+lKO4nbNWWGhfo5t6
4JgByTQP2vJGm6bY+h3SW5kXBVtNuUMPWcV8bfwatpjfSWMjTkdzabWpBbSl0ETt
QuAr9HNQFS861X3NVLUDbyI4lUU0LDh6lFzMCZYVT+3eQn24Lu1Y3OSppO3W4630
e1+E89aQGuUqSnldGCdaG5GO/scWS9XmDrwbyKqLd0GCxP5TY9wh8KYuPP0lNicn
FVvtxLgPjkrROPgyupWNDc8lboc9MYTVJRyRgBQTYj+P0A2yseY93EqUh2L7bmk7
iCb8vkatL/5DILmtOcmWi+9HvRDJRWCKWHK0osVmaF3B8BjBSZ+hk4BF5trakRho
pGMS2rnH6fdfls7THCkyhhWDlBD1v7gU6/AoIjToHlBKUXf2kwSECoEk+jUFbM9w
GRgd8MYYW+SJXDLjLPU4qj4Qccpk37SaNWHzseMfYg7PLXIfDpWzJcvSGwiVRwNQ
DITHu2v94w5LCGlQRYrFJfuO9UibQXSBmJBiC+ms0kaHaXe+hz7tn4ZdTQOTPENL
dUoND9BA6UPfnGSimX+LRcI3e29077kXO4RL+7PpyAssYsVauLGrnBk+DELsqpdu
jpgXdTWBRGhu+i8R/6TZVHfEV27mFU9YlR6JuGzvysi8fX125AqoeKAQ6ERnDLNs
1NIMA3vugYnJNexZthWIq7BPWnk9cUyronnQ2RPWD5ZzBOap6Uy50cdeD8dC4FY4
97nJCd4OgwgtGAkgDoUB15AflsK3zK/UX23rRHeUtUS6CbTJR35aNprY5NK/MHrZ
MupIf0GrnLdxwE1GXwYnfKnbqWXa7i7vyOTMV+p2NGsY+smPmn4WZvOCtVUXPb49
J5RFEYe7Iy9oqZRCD/I9XwxRikto3ruZqIGwCXtL8epqoZzpMuXIfmo/HWeaMyAh
rKQgPshZLAUdKhCwNMgYWQhbNlWmjl6I4i06NoZfFyljxFsjhuFJQa9+MuQz9FB2
HKeU3SoAbU9tEZNN3n3xykT5dRfKLyF8o64NAc51r9++P5CW6Pb5JL2z6nUkuT+j
ib33Wf/Xxvu596Rg4lgebXlkg9hDhh8WlQ3NMwGkZrwNvuSKhZGzkMy9qpc5qqLN
7rZlj/eJHDIdeoIa4TCWDjWpnZg22tcTi3berdJ9Kgf9u7nAnt/32Z1kyHt7WUPR
NjIyqTQXSdDCmkKukFFMWi06F06vNY4iAhwGunBdmzmaSdwYNmO51QAYuI+i1JG/
Iapt86PiLrpHAnAGzYiwi2XA9IaCZdcCZpv9iBFJqtJNVkoB4ikZLHpjRlfYslLv
SHdr3gu61b9OTK1h6DgNhhVvihSPaCBzHiy81Y8/tPcWO/sS5ORNM12XT71/JnTz
wZoGHkzBgty137AorPK/U1C+reyzU71QRPQy96Zv7dCmrNZZoQ7rvqSkhycr/MTg
JO2NX+7FhjJqcdS9/vyl7Q28G2Ot2aTGaibmm1TMz+/7w3oKXOyAzuRJQitV9K9r
qExkNWpXVjsyKZvzGflpO7o4HhhhE9loawup4TgcbsxEj9YEgJ+CPhAjdCoQ9kFV
JI5VA7GiHY5cN/UFew3DxK921SWfVu3VW+Qur/KU8eBjSmaTzP7JCgMRCKTt90xA
+YjJJOzAjDGL0duC/903u2y5I+GDgmmlD4o6rDDt3fivp/Xiq3Yp+vKpkwfPxoqw
3CShMdEhHW0xosmBpblawKeyJLIOKqkSobH3v1frmSxSgUBuRYrzqlkdPxYJs4Ly
SqV25lnZMPDNRGIiAU1zaeLCoTT0PKXoykF9xc2xLnByMd+uEaGufwiRCMcB6n3A
ba2858025QWNnb96J0HW9KfNh3iIfeQb1L5hfJMsYifzxdrpamoiZtFmsi9GCp/a
EHE1O5zeBQQKDDEnnhS9Din9fIyIFTSOXh020anaGfHvfaJGFenLPdnZxHDKaRFn
D928COifl6daV7BzHp3PURa2nTongpNkURjxhr6VPRxnDJP9+aDvmxlie7b6Yaf4
xQpPpoit12xNpxbC4YLMX8Ud0E6SZpeHQSd/CQl5Sx4YxIGLWEuR5FJsoCqm3Qig
HcZqByjktrALRrHQSIkrkFIIUtuk4kUi+7AqQIjSE3GwFAQnz2jdRqj1tdzBXpBR
98vJW91YFQY1jr2yNMLsHqjqjVwn1O3wnDmlimq6+JVMbvG7xuE7QZ3F3hG/QNgo
c99yA780inQEisl2VYqgesVVT8bLpBza58CpL6LOxZzR1KbVUZrJNqMw8Y2F6EJ0
KS9StYf+oNOatU4NduYUBoBTflnSFM3j3+9vojL1tJtE3VZnM74+hd89OnoEvWtO
TNdC3Ka991hz2vrIwOaE3qkdZNRFIU3V86uaoX4DtZut0VrqfX49U0YncctRt8fH
ZwYG7ZOqJYWnsLqrVKL+jDkCeCzMh3vx4zjtymBru6im5jBNdMPydt7aN0GcLoZ+
GPe9RdPTjaaM7vyRQVk5Wnq+RFdUPcluEgkJ9fS61mBlEIsRjOuakRZa6CWF2WyF
SYdGM1fax0lHt5U2GnNVFg+9cYBbN721dOFe0VFU+nZxd643T+pQoWswmtcqwNQm
YiLUYnAqNeRZnMpEcqLdh5VTG+y5X9kvl8CdNaPVXtWfZqpzWBp2nIydvK539xPS
6IqgxaPa+o3i6M3/RYfQioruHiC9bDk3EJ49KPl5PuUTBQZ0FyMXJYxDzJMEGSsN
ZTTyqtLLGv+2d7Wqq2ueX9oJzBPCcr8kz3K/+vc3V6X7CZ8S+ljLXizRVOTDfExM
6ll0lD1d+eO3pjwepX0cnE3cRGueUa+TRCPKJGMBWHIWapSqzTsKKixVgC+AqnEI
x6CxyYbFx50ISea5iqfSfqHP+9N5JIKdg7wiGdBYjQwi7Iuy7u4tk/X8LUnr6fw3
ADgbaE8hxdokIzK7nvO1Fff4i3t2gGyF65T3PcMEEC1JytZquF2/jBYTjaMYgZrZ
wHT/q+OVOYASEkYUPbTlxsbt1/ORAFxeOTI4WLe3iNeNjbr8HabdrJ225YnxGpbD
V0865ClXL1+dPcjTYOUyv03Vg6Ipzq17TpMH4Qjk1673eakczQ+r4WJqn6qSQHtU
DvjyA5mfoYFuOqYHCJzr+AsFALx7WWIZbDNEmLjVhcSlmSQ2TBkpYmZUiUMzB0Bp
qApRA++fOeUd1JvkZk+06RW0/jOsg1evS4kmU7Qu6+gKsscYe/b9LWDnO4RFYGZW
2vQeCLjo0zBjl9slqTb/cJnDdcEuHC4LtK08ffDSewHwdvk7Y30xE/MyNUhkzRyO
TDs2Cc58zLhoP0l1VxnpSn3mzrvOnqBYtK46B+x10xWEKIdwvUm+rbej7KlzAIlV
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gmoAWkbAMQ3eD3WZx7er74gCB+T1ZKoP6W2fOzKGuKRTFHUS5C1j9MA90Guif4Gn
U+8tvYNB6C07aSrbhlGi/lXhT2yLES8vuNVE/q2RU3C8jnbXr6IjT1R/vdCK1v0x
bR7K+J1NXlQLCYLlZpAHXpNG+THTIoYlT+CqEQ/SsQtosLI9rEVZPe1YD3LJMdwU
AwJvBahNjEoXDZoo7pYvyEg/zVEGBttKvRSmo+59KkSaDBEOEgheuiteqLxDasE8
xAf2LQo2LYb/Lb/WO1e2EfS2reOsZhe+L+cKYMBCUQvozwQfv7+fdQPIHugMg9ag
vdhDjjfPfap6NUNTd0o93w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
b1uevqfZxGCOLbrm5yRRY5UZedppLS9Rh7EyqrmlUARmeUF4IqcP020aJZxoySeZ
VGrp1KutWedxSeHmh+V5Og+EnZs4gS/1BiWK/4J7DzaNDOrqzbjOny+2S8zgaJwz
0Wdz6xljHSVXC+k/fAWWM2uPZ0T4Mbp+glj5Zf/IgKiwOsYcnZAnxlnc9rKvL9bp
3kJnVIrDtj40tSb50AoHVmia2oiKuoQD3a2/i0Bn8vKs+1mO+ic0PdLiYWDtdd5i
2eQIbUf0fG2PTE5me8CXDE0rldWDeeEJYIzjtEK0MVQzOhjZ2uxoLWku7jdCRcsr
K58fC8ujcUaDM+OZtlREYMRss2bvoA49gh3z79c/haEKXlSO6y+TZ9fVMr5rgAGr
WG5JVJVRaH/eLiyEOnzR9dxv0agujCyZBAhPyAlmKGXXanZM9scMZozstmmmzR+1
cenCNbXqJhyo0UUauHxJZR1565HFY8L0UHn8ku3XHgyaPoaZhmeQWi5ay307bYqG
6gFutE/zAJvv8rW2/uF9ZVqtDgT69b7nBko9+xmTn3iPfUEksFt+y8sq8VuzFlNf
k2tG/vXrsB5HAZ5zB6if3DBYsGB/eJlLCC97lohcD+QePijM0XjrWSq3bggru1mJ
V1r5VWlWu+QeHJZCqOZBOTvJqO38vC/sveR1FOOO91riW/HMPMehIK1zZ9Wb+11O
Qatl2r1V0q9ZmZnmz/BF6TQW1qRT/0tuhm1Hb04pybsW+dYwa4TefWeuVnG278zZ
REdzRGfVEc7l9jK7GLLxo9IS/xxJ1uyeeq3WTA1Is0InXtgxvLAwC3lWExkGaikb
yiZ2Z4PSNCss/R+909ApT5eR/u5e5qgMU27GsJLhPL/Lc0K1uGhEo9yx/QLpt13v
Tw/tH1sHDCFcgEkAMrkLW98qaA9p2zhBw9ImdverFTk=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BaRhY/A55pkOPG7l111tbcAE3vCwesqpsDU0avRnQoRojvmEnl+7nrmY0Nr2K3no
8NpMgU5orzHQnavuyCjAotDx8iT8pgwmHGjVrEcPHjjC9J9tHHr9WQxXBlMco1G1
til0ldIfEKbPCU1GbLvu255vtJfshTaQwn5+ESC+RsBZsuSRix7V5bnfMDYSMvuF
1wMzQi8sBcvx96YKAk3kgGGsxFEH1b61RbM55BDoc2EkzzNAWRESSAUZRf1z2UVR
sLBhUao3EUUQIPZkNmNrd7PWa9I1zciUzFotiyZ8TC05v2jZXGXeLuaBfvizolia
rwkgCzaYIQC74nrVkzgVUQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1792 )
`pragma protect data_block
ONgE65j4AJe9laK78sNRkAbDNlLUnjiWiJwr3kw3Jvzlx0GGnDqP4LyvcUkB5Ulc
nhfPX2V41QDpe/nwn8S33Y6tagX5vMc196VRUi2Puue1edTIj6s71VFqCOoMILRF
flhFaFMn1JpBhSDWBsWrPRCt1anLlL1m6yVyVW7VEtOB8FIYuHHUbK5d+0Dh4HKf
b2SCbjw49K0G0NtJS5ehhP4xlXnsiKrzNzfCusob/AbZYkz6Fw1K+FenpVen/Czl
R9B2tRogZSrdpzsCuuTQ81EiZVfvklOJGBME0+q0DcdAmhnCf9Yi0l9NcuwmwsD1
lbjJW7l8waipnwdebjhJgUOTYesvfD4hqXQbhlx7rMwJdv2MlP9v56StFNN67DDs
jIFrWtIFuzKRRyiflEAoB31s59HmFupvrhEdbGcj79E8nyhf1slhxyGaLZGfuPUG
h4xFJnKf6Q10IK0XpBtoKJ8coRQG9Py6fGqV3Cwl0FFiggkuU2s5T1/kGqi8TmVP
+e6xQiPXKBp1IKHPoufiqUwgNBkYUkzoDZz39vOshKY+84oqNSdpLGlCzKIOcMmW
bkQGFDMhhScGM+y8Fa6lBPVPKORUp7JbeWnKnzALZrGzO/yH0DRlY/7T1xfDAqrc
/WojQSfVVn/1ZaYqFdyuorGEHNWTUa7gE+0M2YIxAHA//P1FL/eQ5AUbhLxV2zWR
/zczJyM0VTBBEQfTEURfmw8PYjX2PgFbsNjMEza8dr5+YT/MRgjFjGYm8BofuoSQ
ymTD0GS8NwdSwK2dpTTGBVCUSCtruiaQZtTXcEPKcZ8Gjg3exmgXvcyovs6dGS7G
0L0r4uMYEonjEVspAqePzKhYI2QvIHo9pB01qwuLuE2New0GXpe+9psR4VFp6MPZ
WvYPL2+CGdoNZKpOjimmAcIS/cpagpYuLcQybBsV/nyNHtTYSNO8v9p2auz8t5c2
qXCdLKu/8pT8dQI/PAutXjFCRq8W1cqXzoL3ty5AwzvPoZoWtQ+AMocETgIjk5KP
oEwWBAaB1MTuQhQn442V7BcD+gZoKx3oYzZlp5m3Q6nR43/Yt6OAQdcAkHwqpyrC
TIGHTExpuxy9OJLdl1bbhmUMDoMfVXSGhVr7uZme1ChDxVqAiwHG5N0EinjIHxXz
rRcpjeAqM60c5MnvzYBXTamJB9LsxQMi3m09yupyUQ5FxrrrFK9zGKY8ckb4g3rp
Vi0/ysg6pSZ1qzGRbyprL+5rs0e2t/M/FXg6Hlrk2f4TxvbZgyqYQOBNFImhGGn3
FyiO3WLNoJVW8REY02Knve6lYKin41CFSSK3ezw6I0q10V5UKRjvhW2PQC0dlEFP
+SYZe1AdQ97kHlBDuoexEsmQp6SOVU+d7HCjAM2yLNbedoviwY8Y3ZFpWf4q3wZ0
fJ3wXMoJRXhUVvwoIgxpZVENG4rMkAChgvrXd7M9GvgO/Nd24Ms5oEoken4cgupK
v173lAOQm/TKpk+MFqVCGV/hml4RGIrNnR0rSF+89oIRzVxlz8lfO/tAFmjuKumh
joyx+y3kf4hjhVwNMtoP2M0DbR9onQc/IAOhUo3dpsRTGsOe1qkNH93ElnOKY3oX
WN1lERmnVrtgtqZZ5PkTQyUQUpfsbvPbv9YiXYEUySgHMFnJIqWp6FLc3wUORtkd
hbBuJA14s/lJ8QsP+2Q1ohqUumBLzg5womX+BbsKXk32DQjhkIEGEzt7cpQLEsnO
lyj8BIMxu34z7LICt1N6jaXujYsFjZ0yEJPJ22h6vf22bjx8ZnznXamiv0i4M9q1
hd+pEuhCOhNapoxPmJsL+mfFa6wt6gLRu6NuCtFKPbMIAsrtbgOTe4nGoGO0kb3p
/v+9X3Ycyn2o5PemD/2EMD5fBBg6ik8o5UWugcXoNVCLLcyNXb702avLfaXmUBpf
KKnnpLvUfAJyj53k+0Ks0iRhgsIAH0OFK06+Lvbqldq1gVl/Elo536+tGJmukBt4
UJpS40TfSzB4hPqJo8N+OJF0D7CgMO+3zzi79zscn8uH426Q/PgDlgeBQTDmNhC8
t/rrk/Qad+2470o2B4RJXwOsf6Qx49q1bNdb2CA09UWDAwyU3qmRzNbRBASVmMrA
wZotJgASedTNOsORRq3WE24TKOqU34oYUuEt4Jb6SCFI08r/Sdi8IVWZ9iV41IQo
Cy/YDxiSXPNjbMaqsyrbpiI/Nq53x8jAw5I3I5KecAUwJe/TUhkdq9UoVwU+YMJq
o5AIUrKUIOvdvz35r5iekZ8oEcOWC5JiMd5XU6TW/rHgHhEjE4bXPEkM+J9ZqBjG
npXCYZO062YgNe60DgpfXt2Z2yEE9VfEPoLIi3qrv6AiGYr/rGiaKtgb97hG6lNS
w0/eavRMXIPAlt916ddvQA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SkhGQdbiBWB9cqYo6iuR1VqHOdWM/YLojFDMTln9Ir1zjerSQuJ0/QlZdFITT9mg
rWXVIjV4xl7PoeP5b9dT5YmRukGJWXPzHhyG7iBjNCsAew1kdMdvle4nMWJPU9wq
83EAQ5aP3CiiCzsFIgJ/XEFwYgHbQT4NdqX+BdrYRqkPxcIYMgNg5EDHA/3U21cW
ATYIzPbsloz9VlcTlada75qpuXY3YnYIT93V2l/mtg9od/fQ9I452BmB6qnbFMa5
RcXjY6FdH5nbyI2mvQbModTpnrvCLnHGJkelCkY7FCV4HZqv0eZtpnxCHKSDN7yl
fW60+yo6uCD/4f16XNBbqA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 30544 )
`pragma protect data_block
iarNUPnUR+lU0tEvWw9iZxidR46ZZMgMl78pZxtYqxOj2XecwoGI1L+2Xv8OpsYl
hAHEYm8SCPZtwNHsRJoIXbqLzqSPlufjvA92RHL5sXS2vX8/h82P1sph2ha1ZiMj
u7fn9T6k6yO8JVleSktYSWjqIS2z/KL3rQA7h/HI5EeSvlDAI2nV2kZhYjdVzSeu
qlO4KmDrZnBdt1ZLU6xptdTbcR5GCUacPQjINXpYMyHQDluBZ6MxIJrj5eWXQysG
blWwnfEti+bfli78O+rRBEXSZ9gifuCfxUdPnMlG2vcYi4b1XQi5S99NWU9tjgKK
d984w56Crh8fLRGCs/f8lEidXksGMxD0nfrqMc36efsqn5FIqb5nLdIXrHJ+MIeE
FfSuDT5WGHUZRKOiR1QVy/+bF/mm1YkLfMXUZy70ClUS1qdEugbfeAUWKLiS/M6x
N8SQRkmwiJXnvKq3txekEFwCdFebMkQqfQg7WxcqQt7v2VU30YdFb+auYYQomJR/
gXlv+IdPEsyDD9xoRbuVz+O2GJHacUbI69alPFEYeixmjWanufKGn/v0f6oIk8aX
1fmntCsMN7KTzwZeW7bbL2YPg1gpT5y4bFLvt+in58nglAbUls2MyowVf5trqgks
e/0usa8xkmMGOAF8yFMCR+N0VXlggEGhl6Qt8qpP1KDEk3qVJDWYAC76eckHjEfv
Qx2sbBM/nrSv6eEdGXMJw4hAzCkpZpsX4UjIZAdYHKL7HKntKNAJkt5u/QcUezv5
R1UoCVi5Pdfb271+wLc/GedmqbdoBVdh/dxAH63/fxZrRr17FI0G8dVsFvjVbdWa
3NvAbkkC6Nk4JPxgOIzuUDmG3fdTGJbAQ5A0f2uUdt9s6vAKG2rZANG/loBBX5WJ
GUIFUlv85zWNlT1gNbhGI6p9QR6xgdlXmJPqNOUQAmzvsfNg4salU/5oeVx5XLYx
73AVuDF//ZPTGvcV94zzdWb9VkXgkZ6DndNEzNjlBtMcW0rqiSTW6PxhuQpN4+W6
Re2RQYxptlCX0eHxOJFciHI+DAuoMDaa5WV+nwK3mZ7Boee6bFxgaLEtIkwUaIjT
g1JeOq/gejgmx0C2/Bwl0jB/Wy5nB72re2T2rMIxlXGfXaFvVWRfm0CT/xRXlkCb
I5gf/dWhZAqFKtsp1yUJK2i618CndBTjLtahPcKg+XzoyaPc3hO3du0PD6QpK9kx
XvuO81RhR/PHt59e3G8ga3MSdw5KE77e2cjAN+PvbUJ9hEgYaqnWk+hq0Gy2pYXL
FQriwZ3Ow0+7T6EKhNIlaHXp1eDlwl8jmHDZ98lyng/RQxJjSIWB7q0IdX/eEHre
qPj6zXIEym+WEtXWDlJMRwo/ovBLzETWoaECK/nViJdUgmbVSAs3IRlM0DbfZ+AG
C/WxY8Whtk1++cFm7Wfg9sgGChR6L+841LyYocQWZH63gHsXIaK7Qhka363OxNeQ
+bFcFt4otCreMQ0N2M4gkyWqNi+8nL3Ip/HuszbrQtuewYSMgQDdy7ZsUMfdW9Mt
qDJVS3jcMeveq4LVSWOHIetXe1IJbMhT3fFADdu1Hee8AO7Xcl2T5SAV9I06HrSQ
vRKdJQOu6+iO6ZGbB4HCB7mIAlCePXOuCdtrMqyRigUE+y/AhhQ6TLlOKh+h7b86
Fk8ZeIXFvpfo7muXjW+QOSH0++QNiCeiOXotMKygy/fndh0YDE/owddP+zvQ/aW6
pP+FmWJ3hmgMI1xcC+J1tjO7zffZOHKwtpC5nSvSN7blirivtps4nFm2BUK0z6II
56dYx+a1dsD2F6pNfR/AT/LaV6dq/TJ1sI6TlXyRpGIqCkwyhA6IpwWGgXgSYKLb
GpunkTUJX2kDUTgZmsbWxIYxf2hDHOopHQDY0AiAB2vxwgyb2VSGVVT8qifU0Na1
NUIFq5deFGcB2kMRhoyGs3ht07uYg1U4/AEcHca4IgtLg1oetE5OR6GaoPbowtHV
9MiEZu53JUCkhbhBj5MwlVcvUo2w6GMsVREA+3BBZXydclWtEDQKizZF+8oUYisJ
h2hBBgLx0g8wgOru0rUJ3sreAsEsIecCa8GIoRcLqum2RO5PDGOxYlJ6c1av2fM3
vjCiTaxUPmItcApfZIPbd5WjIwbU3HmgrsINOH4jCkR3lPBGbKdeTr9aXM2Ax/f9
HwPIE6jgfAEg6LoGSUlq23uZqgR/sLMc7L0A2TTTSGjLRUYob3xHnZS6BJhmAtGe
CpHOHCGs9uRxq0MK2VJgSYq9LeY9VtWqxH8+PpGPj+cBmx8Ldf4Gg2rBAUa+68gU
d8ZdF4zCOsFiLNG7LmCtGQafGeyXQBGc6sOzdp/R/iwbxN7m+bcGklaVI51rz8Ga
p4kIN51D+6kX6awz7OQvC41p09kTzjXOsMLJYOoJ/SI4E1Oeji8/s+eTYaIAw/3K
+V65WP51a8542X7ac3+FdF7nIYSORNlIiO9hBUZ2qID/qm+i0DYhLiw7yBtZNuPn
Uvq3s8xegKy2TIXcyD84qmBVbXKtxf18jir/chmOy4tkY/DDdeIMl0UbY1Bs6Rp9
pceIxHPFPk0jCFcVf+kjiYRuLb+solVla1CmkmGUVmMcLMwMGLxqlKk0cK7kV2cq
NlG738uNSpLHjTonI7EjQrrfkKG2gGDiwetJXgdA+HtlDgJVASORtSIbZJlAToxe
UzG99rUCXU0y4821VGs3gX09V9zgRNwccdYTrwfVBrcY1D73gLnn9kRJDt5DWZfk
8fU3RjWHkRNDtMX6F5DGFAi+fcsQtAkeAVquJeH3y/Aoq65MNwkNuMDiL5sbzCYU
zHHmvU/Qsdh7PN3XAp4eZaEN1giEdDxkS1B5wYAIvhDZDFl2sRPRF9zdTH009S1x
lt6yPxgt0U8uOh9CVBbialJsqdGbAmroeExB7FoVWtFacrOmgk9p9aKoPfya890z
4/fAOXK01ptvzIOl4cFUIjji8qbc8kkYaXM4XrhWpaIe1sGSkpfIUcyjV+vAes+M
1aBZhVPtt08UJM11h0sILu5tDvjggNqYY2pvEBcCXmiWmvPd6bkgN1Lc2/Pbc0os
kM157nGuFuyjXCFQaEbGYc8vbGjoasmuFE6nFxO86R13ibLeHR2Ldp22TG7vpKkl
ZdhmY38xndFB6FadtdaoUruKIk53PE1sCaHkFJ2bDic7MJ6rWIi8wNvakOoT+jTz
i5dmY8osMKRKbHg7XNZ0N7Mt59r4+qTTyWpqGY02GcbgUBJjE+VxjPwA9ijt8vjN
3rVwnfjK/JZSRA7iJROILzQrpIZ5quMiQeFO1M9FO06bt2QHBWBKkBOUPpdL9As8
2nnXiGBn2kQy8YEoqh27kRjTBON/Qr6UZkBhmJlU0tBXgBTaT6lp3gA7zFMUeCki
vEXidyTkn25FKsCfLAAW3jhy/4taoVrs+lGmtSGFrE0jgoyDQgPdgSUcpbWaKawB
LM0350nR+H0tFsx9G1EWvwvolc+z57TZne4BwQ98eadOz9exHZwaHy85Q9rblw7a
XL61pXZFc1e76KhdoO7c/hWpIwctUIR7AWryEl2lrWurh/I4jXXByapChY3L2viK
NToTknNdkY5Sa2Zdi3xYB8gJIsJqqmAfTyma/yMG7RP9mXCeFVjbesBDs378dRP9
kZTuAoqScBxYksnj6csA/i+5JRgvFXaXoW0EyIQBqTQTkC2TDiTHS80q0r2AGz33
o4YjhQI3/VWMp+OGc5/kXLAHikGtGDqiIiIU1BP9qh39CobEyWNCuFyGK4um2BuJ
ejBNcBp8i69Ui5V9ZTeyKFTXiJ798MyzRagKiQvJxsxsktMZLUEH0evAbBPuj/i5
nHfxolddGrioeke/f0CuO3LQ24I8Zhnt77VlPaSJYqgM3PLwgCG6ikMwSf2OR+bS
BBB3egxQ42BgjaMmN6vQKzcTnPbOwPu8iKboSzzfo5/KfdVt5ZHTvO8WRjbEetNe
bagC5f3LFamiyWC/xV6v52zL1dZNtK/BybRh86uLcINqd4creBUhaBk7mJX0ptHX
4vWkFxsnmQLbq26MyDIyRul+zYqQ7gM0LuKPyXNwhMGo4ky/mkGZT0xq8ilXf4sm
6luXsXjnGm7hbIDKdsLAFwunQ4H6AZFkdrHP+hykP2FRBAuE4WB/W16cjg1Kb/fy
sCFkjGAFWK214Q1FlUgeoL0CBVLj6aNWPachNUNIr0/Eb36NruBtcxZUPKfYPmwz
n4B88WWJ0LDtyXIAIvUxXJHeZlgvAa4IVoZ6Wc7ax6iSulNIeb39Y6IqRuDr5kCm
r2UejljSMI+0ynMya2CkgxDEySUoymfAYsSskoKr95s8OVEJPWK8HLh7g6a7Ql73
vAvrEOP3tb6HVznAQ6pmsU/x20v3dWshPSnQn0TS2lgnb4z0Q1ViVW4H/TsOCx37
9zvhhqaXk3RVSjrFddQTZV2aQZY2mcaWAmzu5epXyI2VkkOrrB+aW8R6DViegF+M
XZ+QFZ8lMt3o6olyDleVUA9/t5j57qJUXnS5f6fgmKkXifTJrQab4nmGJIcVqnkU
JPbu4eY/Y68i4k0938LX9LvJpu1KeTgoZ6TqC1a7gOCMIiPx33wl4BlsBObJ22xz
FEYKWVWEWC3mVLWRdR2hyvLoJZuWI7F8/BTX+8Fb0qXxGwxnW7SyNWj9u8IC2AyV
OYPg/VcBuxIasMWM2zBznafmS1yosfHloqHDkeG8mHWb+88ucsYH/gJ3U8bf4GbG
YEshoCJ3iwqoGj7pqtO1k2U5jiPisInA5MWuob4uGSK25OpE/B7IBWAx6JsJq1h2
K8+r2XwmnN9HOHk8nOM1KBiSYV+bSdjmRTIz41wxG2SxPqQKLPrcV6cFtyNtGKV7
eZwY6KVxodzPJnlQUjYmdhskZ7cgUtPMFw074R1xaliiXfKIXAqHVyw93Wwp6P0T
FlSzQtq/fJxvgs1b0MmMnOpBgRYYYo2sp6P5kVa3A8zmsK2QgrknHPdOy4YFgQrt
ZwEL2TaOF/ky0kKMrdUZB3ijaP9kYiiEnu4D1hcCNHZdBBVz0E5as+H3pXLAzkMK
K+/Y/eennc4/oBFjci2Bn3kSuUS7tCHYtUlP2wyO850VbAibjmuYlrjeM0dmrzcx
RVVJk/8pGssjvL9Rz0DU6gTyt9uXAYv0JxIlmT3JJoVzvFHOj9VwPi5FcQ1Xj32b
8Lm1C8iA7FDAIYoX/TwAXsXjVm1OuvQIqfyBMNegCyPvmCv3U8N8bBCvum9ONAts
bPspGifW/bIiBX/G5D4JUr//iGnCI1CaRApEDOme5vr31E9elqBoFyZaDtN09dP0
nrFw420VCqlte9JIFeKwC+/2nSWDoeHnp4xbTReAgY0qvSGnwcJB8zQE+Di04+lw
s6+ynSQb/2q9YXlvgLyvVxQ100yQ83ul4jr27V26pQfh7kZBtwkM2fbFecNgJrXy
ht7haq20uYax6iolEysv7ASu7HH+tDyVoCdhs3Q+IkcWZp5W2PjqDOMduADAPbbZ
ncFWamfM5cv++/hjwVfSe1fvknUKvERAsYdw0XJPsNB13KgR+Qqp8EPpmpSHdUmv
MEiqmCUEarkUKoMsjhcEQX4StBhMcbXibPvlk1i5YpVrTEApLKFgscn5XpB8Icef
W0U/U36qUwu6yFAfFykeP/Sk+xOpjbcBL5DL/zJIrQPEL8GE/dAtxetfff2mLtOe
qv9FmDZBnCoNz5w3dAk9/5Z3TcJbLU0ex5QyMAjsxN+a+f1mdNal9tIYf4thu1NT
n7rZ+jiacZbuTiv05mVqb7NrrHFjX0JvlL9wuin6k+qE0Z+SchVggRrn/Ioz+XIp
4nUZOvenBaMP7NfdDFo5RJ4iibrezfHNIF1G0h2BmNtKUUe59J7kpzxuBPKpupBy
4s491duY7LcY3as35yUzxqcsYmHTe4HKVjvoThJQQSkFwZSUs1MQSj61xB8dOeUw
6e4Gnq0uvW9FJ0pszPghT2e06jced2ssC4vjU45ECRqQPK+hTUdlGfliibUhNorx
AgHrQv+NY+IECwgTx+eNI+NarU4p6ygs7n3WSR9TCbvThuFubN7CcsLUgbHzZghw
mzBpyQ9BnpYJvVHP/FrjRbp4c9aUPZq/rCYuy+RmHNwPMkeugqA6VV4qL3DFZMb6
9Cuc0+zpo8cE0OIH+5gjE+IyMna5gCrXjRjBD1pfRzAxzKUK9t9EUte9dYlCQG73
OpwEKYrZ6inzLaqzTZR+/NlFJjAHbFAX2bZpB6fr8AdvhFa2ClY74c8AYoWOl1N+
85K2sp6QJnpKb2DVs1Hd8yGvPpDnsORtOTbs6rxkKSvHyu6xqjwySLnEoelIW4Lh
Kv5icPkGyN8Tm0W/UYNxu3Eo+66lyS+8eJs9znmggqjkQX1TMYzOd3imnUA8TI/d
/vA/NtB5bTsymvOtf4H9c4lNWZKP1ZZFDBTyoD7GpTnS/zyRdqy54H0rbo9PDQA9
sGPRkJ6HhDOuFF/cvNS3hEH+Q+TZlOqG9zYS5wpEc2r8/NUBECEsWgK/ApfBLtVB
+I0qdoXukrtLev1b5L2xw4ZM7Ep5GdITN2775GA7s31Xj/oSKmaNIehXiRNVRNSD
WpxkTB6DjJsNLJ1TgjcPxdjf5SIBS/2N3eqj5fK3MNQygc4FSJwnX7sQcUTjseCY
rTRIN6GgUbD4H3ubMcBv4NdusnhKCBHKrjUQjDU+ZCVxpZUcQU9vvdGif6qfgxK6
3XfgrIZSzQw9yi7zdYjy9Ay/ZMAuzdwAvptJSPpLOWAlfeXUyWDpgD1Bu6xPFdmG
h+FMbjWJZLQsro2s0QqptFNcup1oEe+ldNZ1tySZngev9zCDjLrXVSR+lZQse6Qm
IZYdSpnhNSbRxDZqzYq8s34c9ESF8pES7LOm0Awvm/NWPA2XJiUGElCL7CcOtj7b
dMW7cZr+Lna29NukNUDxCZ6SkzqyFh/WZi12RHmV8u23aRXB07gJUocLs/wNL2Ey
5rkWUPzg/F3UB73SyOm9jrIUVvPqHnqYk5DhWJljy+SO00z/l/JMQYaZF8MYFsVp
RSdtfbW8UeOdVhxngVbG0nwxw1IEnzOPtfuFh+JtT8ruX6j9qJ/dTxxPBMW3Q04g
A6a19NlVpezGprKqu2CdEJs8uuqtTY5SmXEZd9iSd2Uh/Oiqoqvn9UdfilHIb66j
vmNeCZNopvDoalIInvmc6OyMg+cbsyQsP/aTY4trmi1Q9rxPbrs/3qydJHublIRb
rSmTUg2cZ1WFonsqbREBosKKe7iNv+E+0ttfNDhmD7+Mp0ssvu0dQO5cAoq0Jr/r
Gpp9mYGGfdvkw4Np2J46moj5Zj3qnAE5w2i9zI7v06acGWxly5AU2a2nztRcK/os
VhXLEiRt9h9HlOPuUkWJeWHCW8obdHsX5xmBLnM7qgT/WuD865U2HrE7tieeqnHY
fZwHzdb20/AjJuqlMd1ExpH96PgKNxBu5tZ2p8zs+QmAVPx+OocNqcQWjBTevcQ7
KjvGQs9sBJXWTrKDhrIzDgcJJnD1/pub0nfHdyu6H3cwSjyXOmUJqzJUi4rTtbdY
L64WBrcXldj3ukdb1AMZnfekKXyRJG5Co50iAZPfuV7ctTVgv8qfWnqudZyu51Sp
njMpdwVU0P9eYqiHoCv9uwlNWGh0EA63R5BIMr7f0XQs8I9hoV2IPcWnCrS1VvcX
iZspIKgdlChRyT8nLG8M4alOlZ/pn7gD7mCdKhTZlMhdeh7MNr1IrGawwMJ1RM/4
XYqQk47xPzgtI+VbulWktfEOEPO+uGowUZEOESuDzbgPlGeoV7ZTXETIbs+AQ9we
rEJm/vS0rp9o7cbBHmS7o2V03ob8IyyQXSbjwXuy4XnXh56Q+R16q+mhV42rSEAX
yw6owkQstCpkEb9DYA9hOKg0ALEHdxFV5ic3ocYHr/NIfSYvM0u5HW2gt7+jKAH4
GHltIk8k/EUCYz5MchdYnB3MOBcQZVnC4Um+bUGaIEDN/JYWUL51wby7eFVM9E+6
kgpXoppVnv6S2eJwGOvaP7dY7wlQRJb68F6vfsfBuJakHTW3l0PDhl8P2K6Qf0X/
v1gEmn3KWwHNTtYo0+32W8Rr6Sf+MEcaYGh1CHz7scMprjQFCGGP9WYrehNaD08I
YRwI7DByudVwBVLPCWjqCTH5FLUyuqZAyAX/roc12QWzcSzERfCeITtiu+rg1Rxa
x191upvebLHCqY4yJsMeaCaPAUBm78z87JIz6mAjK+jGb67qvOaiLI3pDH9DR0BS
deLfn21Gi9I6VHvJ0snm9RVMF+/nHRjyHUZj+F0nIxe/bFnxyAauRV6bhFCR9cok
P+tUTvnngU70rCYjJHIAPcGGiLkINRKQkbx9Sp9ijSiA/jxxWvNYCrDvwY88SslV
MD0tDt9nX7a9kYVj+BjqFHS1lHzButbLWNpA3t0xJLsI07oqAhtrFLH22pxzqx9n
C+3JUwowQW+4Z1N9zHe7Y6A5U3r3aga0lSW8rRo51fWpvs0XNymPldILK4HkBQNC
DAa58N+ZuTPfgpgtdCzB9W/Fxmq53FmSH/Cu7OYshkhFPnlQ+fiVLJ4CNAiOZlwe
Lt45t6WWY/ftx+LgsBvWXwuT8Wxpx0VFBqfV9CcJZz0vBXmlWGac1Hz+doKZPEnk
KtqtdgX/ntKnbNw6ztiw2PGMA+t4YTssJlbfUsb9Mpyx1VsXSmwOyqTxfGrVEJmK
7iqZEpI/43HuanuM2pyWi2o3hoMZouqGtiyDtbXU884CcDUzOz+LihVQdj3pxkkB
XFzjMgHBw1qSfWGSi/DX9Mi0VdwFO1q7LpeW+OB8A0SaxIVdeuO4OwwM36IZVrgG
nJW9t3ut9CzVaQRdYQu6BiYQ4ZzVGYoUL8Z767hdrpsF3kWQGgu5bdInI0G2d1X/
3rA1pphGLl+pDyCxHNXb2yAGcaUrVBvNLwCCmwvBYv3uhOGnu6P7rG0zwo+r18sU
DtT/C4uRE8aSixHa1iQALBLJtwJ0gOmRdK1ru0J4wGcSOjk1nMzErVerhm6EbQVa
KLF1Qr7sWmNrNMphF83PLEzeSAE5orWag3eIi/FOSxT1N7/3AiNRt2ImLMYc1ngT
7Y/0Im+/tbOmWNj2+fFMBPNvhbcW87LFgeIzANTxpL/6p/gQXVi/CRNF72u7vKGO
G/J73OhuuVM1Hbfovd3dhbJ9ijCreBjh1TrtST/mcQLP4LH0PRTTpaNgOm1IxHiO
0z1gR62PFjyUpGcOIeZ1cTS+s0rcaEUlmNhnaMGb8vIAPXjAteri2eeIPAVuaXkI
oGEGzxw74RDOf2wAgMQPuY8DW6Ovn542YwOBw121QAfU9eaVFXAgUQThKgPEicln
tvneWXYdH40MOcgdoMaqmwROf9bF7z6vo2OtTxbiOO/7WRF8YxFt/oj8A9ES2v5j
LQr0Bg9aYBF/MKqKLkRYsSqv+RhGEXEc4zop2hgjTpCeLHxCof7Cp8hmI8uIcgb2
HB+kPXic8N8zmOo0dZNsmg1V3CV9B2SmCDTAregz1TT6nKMzOF3c5iOutcKAAfYg
yiI2S3LC7Cnpm7ZN1pvGy7mN7liz22BU1TBnsFYUD4dMcoseu+IYMYV3cJAEiV2L
14GNj8xReHbGHRBaREpY6/92gHXZN7r+Brl89blm9S1/emkJDlw4AGmYP7f8QL7b
mq8bJpCcVt9RSCSjgejIDvJxm697OQ1TweM1rRiUKSG5m1fTRi4I9a5zmGuVbhsP
bOGPDqYu9Ieuin4/xU0EXzpO/i9jY5NdoVpHhlBIBU8ElJGTAGZM2WhIlOEhQ6AX
FTbMb0WKddLTvg9dfcHgV8FUApNUhMEP/fftwFVnGivCKdDqa+/C3clzYxW2epfW
mHmjpzmj9J2mVpQVB6PhfclMHyqUE68LI3Hg1L8z4LkpLyZs8Bc2UrUkHPMDD+7i
XRLdSTeBW0gXIGeFiWX2C41FHfLC9jDg8AEmi0ugEcAX6Jk5OCQz94LJYM7eb3RY
FnfCaeUDOVNKJkJpBVTtI8uNCTr60O4yk6+ec0ziMnqGtgGTAULY7UlxB5uGNqOL
Xze0BJay92LdGKQjofzBIJ3XLEgn/DBqEHkdQy1jYkYyPip8C7Be6cxGY0L3Gymf
lAxfQLFzsMuuypHXhVjCw927TgO3ofcvD7hPl1bBvBBdm9BI3XOYfcvpuE/xCq8m
beYjmqVNOd4rRh11cGsjMEVzOX3PWebamFMVXLilJnLWBj3Ar1LRjiS8B6q7Ich6
arX3WTg3KMuGtU1pAZljrY6mumYGOQCtYIjXPcwRzZLRmFp5L1v6XKD0VjCz7wiX
BPaftKqeM3kmRNlU6xgpF8TkntryxKmAsULi4fnwpwEUUyBdxKYGP9nW+NOBiPBC
LwZp/IWFwFuEdsC0hQC4+VtXQldD5rYvL+SBxYTBZkxHMghR5QMuQVdOyodztZkZ
g28q90YWQSh1xzxusEaWQlCir30CWaoVz3eMSNKnxSzoVSkwK0tikw2s/u7AZshv
JItCo9s3syDEp6sVD2WgnNQaS6YWjtJp/uScO1BxwuwKhRpeeMkTFlHZFnkVlcvB
oGHGsGg+zOBtkMafgFksYVlqMqoxLpbF2zLyLEZ81UtNenTuLxhJ6BJxgHD1dzL2
Y0LIXfmtOO05cMl6vaGE83M89nQ99E4dD8KG6sCegZ1d0wq26oNH7BkoZ2IAzgR3
z9MyEIc6A9uoR1zMlC7+ELH912h4k3AjUmACSGJd+QrNqNes/K2vehmzzA0XBxXQ
a/xQ4V8j/vUKVAQg0mF7OGZTFzLdAV32os+BHGjfQ0vLpcEvQH0eL46GfeGYatzN
J+HdjgBm9QNEoNnNgyEkX4+NuIEdxD/Kb2UL4XiX0WsXd7AEb7VYlDDx4uIv/CpB
iz0+XNZw/oQrM6JmRoM5bJAtyRjKqGDZoSCMG+o2FVS/jyAOASK4LkhDjbRd+xcI
H0psNr1DsvKDpqeE4f33tI5iDy2KeoDb03t+GB5L/HwcpBmZy91//M53vl9WeteY
3VJElMqTkJSHqCLmlVfSoWOCvBRGHdLQBoVigpa6cQy8E26n8BJ4Xm0pg7ORbJp0
JkYM6Arp+TYR9wJAmLOBL9DqrC9xI9Dr57mwLy29pHq1YD6Anvk6/CkNWUyLJcdw
AdWCKmr/Q7MBm9Jfic8b3hwiWAbIDtXhrtb9a2Fl+dtphMT19I3PUG4ZWjRu1HZu
QGGdJh4piTvcxL6FKwZydIlPrEyWF7zMvSWjZTdt8r4OyIVdaDO4ppYQfF1mTZU9
0CGkyULAGZ1dwqZIdyFXrQ9Qunc1OSs9dC9GpqeRuWc9WudX+XhORZ4+kcYBm7il
JJZISsCux58cgsc1WGqm2GLkdOHfhZj7IODoHgVsPDQ2aZAAgmmXEudqbW/kh9VA
0xsZvB/U3k46x2yAS//cwcIcn9OooMPRxCAof/2GUyfuSKprZRSmo77IJKdVmBOy
hL7y/EuClolt7yRlGXsFrbjvTsBLWdxKYl/SXjod8FqFb1xpXCCiujT81/fmvz+W
nwjrgxfx2tK9El2n1Dw03x0XzlgrRpffbk3UDMaTqkoOnlSkQPS0LPyVntGaWOS8
OUfSf4FJ0kTk72tRbJaF3I0GptCy9ILhKlMpdCeGUb5w6Dhbp2NqKD9nxQP8OxQh
GekcQlHd2KUmcsgoJqWH4lIs1g/xs3F1lQXcSATThZFO7IvKVsmG8zBRJCWsSWi2
zhJsuhI4iM3GN/MZywfHJcAhXpMeQk1XjPGu8ejw27RadyydbmjMyFpPanuc0vFX
hr9LLMni49bbmR0EX2+c8viQd6AcyTCr0gvlG6gZNziSfqSSwqSJXUD34JlKGgWA
/pki6njQRowzWdZfvJpcDsToTDHVQiXwJXHFrNtvIGa2S0U3Ew75QPUTXdEwn4N7
/Z8qQlfpJcGIfC82zxZLJca0jyuh9+FuGDlJA8eHRbnPOwTsYmX1Y4jxacdCr/8O
+QAAQfhUc6my1YDaUjWbe5NnJ7IS74UWai7r5t/rHs63t7ENvCDwGlUw0CQGBDnS
puLJYxJz8w6jyPCnitma/zGW6vBtkO3NZGR/AgmuhFwI/TA9YRM3Aa51CE7X8alj
G6I+v1Xjsj4GMRHjLZzMM45+SeT1vH5xc3erlPybzDmIBXYRQIxNBGP2oPJaJOCy
4ZQq/0PWK4FWMKeg57nEJZTzE/NgAqSEh8Jgj93AWMbn8iFJaj/FGRkRQmgMbQyY
ElegVwQ1Ve0JNe08DHq/89dTbOlAZDTlPYO30+StRGjSZicbSGFeGUg5Tm/3CnFO
ULOrPPOY5Ikk7yR1HJbTtq1V1vqe5UrBpDjqprcYgmYGvMCwJZOI3Au0O6WIuEq1
nFHuwVUL+3wtu8YacRFWq3TgJ5o/AoDSBHU+Bv5lVQIN7I571Dx6nZsmsVnHn+j8
ZkPdq6rjMwSl+PeK4ejxzz4OigcXPaA2+EFiq90Yt3EsuDox6+YZUZNLZFmAOJOM
1uuVm8Gp5rMfSE0H2BM2CCM6PnNuJDRAapRNKaCz/CEMK1Y0IX4ryMZlIQv5aXFL
nU+pic180wbK3Z49MOrMPbShmPkHcUJVytH+3t5++FZIj/4zPdB1u7qHoEW9cGAy
d3UP2a2RkTp7PYgPItoQuUmhsorioMNrCg3kDGnSwVmiebJKEFLaLRkhKV8mvBGo
sy8YhWVXXa9B+y4EIILkx22/QG8W47vH1BODabVZ87whDLqliNRotQCDbj4+3c1I
KwXWGds13fi3eG9hRvhKUYpunlvnSoCZLfdJfABeL+HCPINK/Hy+CLW4fDu1y1U2
Dt4VGVIg0ijlrqppcTZaPinKT7rfx227m+82dDLeRX5LEpLgY2XVcmoHrmStacwE
Xnc67PA5OGiLGCBXkaVrLHp04lrpICQfR29nuqKvVoEpigUh4FMJokKZkC5Ae7Zp
b+lz1ccA17wwjHSNLbVu5hN4mVCCtf3WmQyVBtk2uRNJhfMnR56dn0sHGds6oKYI
/qscJKUbNdtJ15t3aB76HQOPB8oA4rfItdK5CuhIKBTGt1kQmgvP8n/WEMwtGLfW
PSOTYj3SttTL977kvUh9vIkHd2RN/ckJHLLt0rcx5hSzq4QhXy1A9D5/wG2LBHdo
humMTYQVDG3GKGg/Yx1kVRzM5m/nwuHxQuUT5N84IKHYbGlePsbrbExxvNIdrtqb
UbS7J7tWc6PEo5zCSHzRpC/DxkUTBNhj0Z2Qzem849gk+cCHRp+h7LaBzMZNsnUf
ZRjLxwM0FIaoK/M7rJmSM7EiiOy0ZfyjNOR/yVRrvCTSa7TcvUUnUTFvtBP62LJY
RyWy/ubU7oRxMHYoOkc0Zj3OiWLre9V+vVLuHyfSmj+S6+n97uBjNu+fY2zUZBgS
5Ci1uPzKlMolPUCPrwGGG3w+i++1Wss/kCzBtEhdR2zsUfGHlD8eT7xBcoB2cRaw
VB5hxcZDIFjI0tW6owpbeteIAjTHVRoYw1NSKB3NykKofGrDH900HrLljbXayKap
wq304qS8sVfFsqIOuoI3qnnPXrm1MREf9tvuDA5KfXXsuzuKvdW/yiU0KimD2FbP
Fl0PLPHd05+t3FCroCtSHQO5Hik3svgaY8u7tfRTADy1VgvXvGaHDz7dk94rO+wc
4CklrOy2EMEjFL5KgTKKgcLFcNS2Z57hGwFTQRMKSXcH/CpwE2pv+L/S607muIz3
dvPEU0IoG0dbVjPJcUnzY/0ygf/UDddd3f0kpA8muG02GJovgBY3Z0XWhN2qecGG
NjdRQu91teGRlRc+36TIt5WXmvd63uDxIC1iBWb0G3SVFWR7A6k4e6u+HLSpK0a1
gz1Qu5puvNJmI0XHRgGYOqaMRLehTHiLAKNlefJZ+LclTWFAMEEsDO7DFZHB1Ho5
6Jn31BwgpsLlg+Gzw+Gz3hoWHD829tS8OVLeuk+Ik9NxMdhpbZAP2IVSf22pqTUC
dCNjPg7taa4b4NECBjiPdjCOOucpLX/XJJngV4lKG5QvmWgIIs9LJXWant24RwFT
FgD7j7EtboEOAkcVbQFuUcii7Vce7geWHLOiUCG8I3feB/D2YpbN+v7P9Uf1aIzH
6n3qnAcnJuYYb6JwPAdQ/IaYxebt2TeEB79DoWdfqE23be+VgpZBXAFIlAHpLyJz
ZKKvISJPwATvRSp72TrQ2i3InwwZfTXvY+4RL6VxDzw5Rov3Zf8IFl3yAVUruUEp
MVC0KtHl8DrIpBtrkvHUgpQtdoFsQE+MKeXnbwo0JMt+kF9JPXCLl/faa4CofoBd
D0uvjPUKydTMpJQyPvhyZ70TdE7MWlAPoZWeXgYPVXR16hNTdgOAdgdkZEOOwwOd
zxfe22NbiMbDGM2Gv5WNA5O39D7O++CATrVLCZglfA+sjJ+ZF0SOu6OTg9o8qD9D
/nOrv8NKd3kqXd+FqayEPLOTwrtSCztISpI9mhZh35J90ZL3PS80ioTghwPbQpJz
hC7Ei9o5FMUt22PJXksnoh2qRX82hZBkRlPFyRKqUr+aEFrIy3M8IFM+jDM2jnRw
vJYeAFFleH2qVVjwn4VSsyBH/7vxjebcJ2sQidCabMx2HZua2Xi/t6SK7+HU7464
uGtLU8d6ylEVJKvpfL7BM9kJyz2Cu+nUOrbOQDYPceZP03oNJGyRajOY05uonuG6
gAatXsQm6z1M2hNH5L1SeMOdq1p7illzsKquXKhApC43z9+LADB5k4UoCjzxkt+6
CJPA5gTRRBE7ygCPf7JoNyrWQZNctpka4OFEa7DqtM6ue+crpKYvt4z7yloec1mq
lO1GRQtLvrpWt9KM45ca/bu9rlRi2N22AKgNvEq0/B6oyJKWNorP1wF5IMvraFq7
qjOiPu5+Ki5Iek6H6plMQ/Kr6lCfag2C47Ex2oF5HOlYTJtY6Cpp/kiyP5AurvMk
ad2RoLJuwOqfLdT1E3pdLaBy0sCEv4qYGML1UdlaGX6Dc/6u9u0cRraTH3H2l1IS
lGo1IqJO8ZIsHUGGU0WSi6Igu4b9z4qrPKVcx3Npg11uvbWtnF18UMz37/X5lAjX
sbrjvkIEACCGmHg6jrEwICPlASXapzX2DwwiUa49+kIkTxm/daD3o1YI8TPlmlqG
Vw9+gp1FkMZPv+lXK9Vmx2HNFezQed7W/aWyfkayivC6H+UTv67yXWiacZwzXtvs
+uJvkC5YoNSVG/r7PCO4lWDvx4N8BoadrUtjv2LYuUk8e4brOS2k7yHe0I9wuYGC
CpVgQdJLuDiOYep4NY7dZ5tPcgmuPkOgW+Y1SipasIIn6fGYdwHEi0PSrZ6jtCVg
PD+ML0aEKvvto9Ib7353ovGZoGpWpAc1xzv2o/g1fxeoludIvULCID09rZtxOaCr
lh3R3ILtnYwdYi3OIebJJdG4kWd/X5eLcI5Z9h2fZciaqtI07KXr42K392RGEjTz
fD0epT5T8vcwTH7t0Q+4vd3cxTVQS7wLX4Wq1vjrV0+/N5/g4DS77Y4jAm2DKJre
OqcJwSZl5AlrXbs+NgcHCI0M2d6FvCb8Xl/BDrbpuojLHyMCr5uQIEGJ1ShdwQKk
eJ3el9H/XyF1KiZYi8OMPcBVCS8qJm4ij/L/j62l7L9aQfDJjcUIfpQnVW0RgmD2
4WI7iZRaH2a0v9tBrvggEnwJaZ79BvcaVUr8JHY2KG+8nczAt73KygK6kQ8/tQmZ
jkVS+EjZ7eOaxmJNu/la5mAaQApdnjRhsmrpG+lqfdWnpcNYKbm6P4n1w/f6RY1B
Z6LrYZaSONiKG5nWjvJP58GVPkQ1XqS/x1Fvw5h1QmHZSeFz945xYU5hOCchyLxs
6IdlDxh+JRMgP+pUx0f7GBBmV6M4TQCCABlM4ZR8guP+trnZIFkJQnTmBnggSNuU
RXq4fUlRe0ufETer1xMzfjso3uyfbMhZBnMTmkofbOAEa4XuuYQwF3Cl49c0PPYG
3JJloYqCVt/bcKpJO8HC0EKEQNBHLxaTItxmkQTKskgAr49qp44PGExhRZO9XA77
2QH705TEXx3ROUU60RkY2FZHC63Ngqyy6YjPHhydskRWlac6JxyAPscTxmfBhHO2
AuiVqkQqSN0j1242lRHi4y7uhhP6ke3uinM4zBI22g0eHhYHj/ksy5JVkdg6eYyp
tgTNWrtZZsMRdsMIaS3rXmL8w4Wz2clqPcQDKrX2I2pbiZ618ygLs/OqO3kbfZHJ
HZ7+m4e0nST+Cju8HgE3p9SSCDf/Lyj9m4tEVRR2s+7JHW2HAYN4MrAbMOnC3993
3gYHDFy4oJAX3nGF88LvuNdl/wiP+4xEeAQ2WiTZ8JEe1yxTMxSNUHAaRklKTsWo
Ow7NTbQxiZwH1lI/YcCWDqyFcq786mBaXaiXUhMzqSIza5CNE8+doVyzbppaW84u
V/kZlEo8fVcwAQx7c8EVJsIiSFKHkDEfAQIkJR8Lo/9EyEzjmHLhV/OGQWOHiDji
ehmeDkdOWuq7gdjAJABdyYOLKWIVPr7SPJVplx81L9ar5nEBRmoG6qYEyLsgjLKn
1Qb/HMxLSNuLll/fzqZ1Z97ImntiA4oRgH8oCLydUM855iXhmPnKBRq7nOE8YXOV
Q+rC6hTUV4FhgLbVlfMGL5x533XLffh6CtOEVHpQPoLZ96omBbY0hXnvlmzIvcE9
0uUxklqH8WMxVgIExBwtgoG5XGsfiNO5DDDc/ZzkRBKITKuhAqwx+NTgkDqoJGg2
UzmHlzGMbdS1Ymjp8sRycke/0XMcLoC4XrxcvIIXK53s+/Bxgcn5hi0FGCyOAhSJ
lmQFFCWi4sG5EfD0qD0jnyTuOx6EWJr5Kzy36ad2IyTIPdxcQO+lRjX49S6HjrP0
PxIYu2bYP8WcfFj/5okRjq4R9cjBMh8zPst4ZMavKi0eCI05OimIRdmWfu25h4FW
Q96ttz2f2KL7g9fJz6wUXLb/PRSQTxMjwmY+dro6Vd+4CeYLPL/k8TwLWC+TqrtF
l5GGvNIppPzEQlL3eHNXJvCCfxLI9Dp5XHnhr51RR9/MNEdPIA1ynmOB4Hh/wwnw
isjmuwXwZDjwr7MmfWuV1YimAMWwYqDFMpZs6Nq/1IWdf2CGZ9ZfUZYeC7prViHU
nP9WWVm3qaKFNxsfuY5v7dBMQ9cHsPDgdvyWX+RXMX88SorA7XzMfCRETg5ykC3L
2obpZEBm1AqMsrAL99E59H2gmvcEgcuR3pBdE9krmcdX2GgdF2W52QHwt4GE5k4V
C7sXHxm0UfptfyiIooTOsDD2A9vEt1+wOtfSzv9M8dNgvKVxFv7voEW6J9LtSVXd
x2JMOZkaQQEd0CrkHsNfCzDZNEmOB1nZY5Fi9hXQAY4wS8S60FlqA/8VP49E1RV7
7iSv32MVu3Q0Uf+1rVSuWRQ5bZgxs1MtidCN7497yPhsgRz4r1VewdY/B+cmCdQF
L1RexLSsFt7K24QmDG7F977hXOvIsrc4Cjq2MzdbU41GPPJn2AIR6Xp+u5wM61vM
EVxWbOcmmJEdLOVzwQbE+ORiBBoBtCTLiiOkbEc9deicaX6JF0KfKn0HTtwwz2h5
BTD0nxGgGGlcW+jV5GbhU3zK6FKE/EJC/KrJKB5Pcv4rDCDlfzy+K688ePeMW2Ef
NQsiAFL7MsE7YQW/Fg4ZS1/sCDPlMhFyzoA8EXIjuYSkTPfLVP/oFHB8BVat4gXr
czQLnRviFrKVpWzToWyXckns3ii/L1iFrpadXuOXx2gq3/f6lsh7AnNtCt91+QaS
9HMlMPRfPcBm2lpCTzYlIe44GxUubX2jfCYQHqYFp/cT9Tra57/FW54E0DysIdiV
v48LZ9tevG76k1B43T38sULsEbY4UBkpwB0jHq0gIwbPZ9zWu68ELIC9GZAnbnLe
ewwC3JBvvM078GyJuRHbF9Kih83Cgdo5lMPrGhLQKrKkSKAALl/zDoz2OaJ4V3Im
7qIhrGnHdQ5G18KIIPH5Wvw09Nfoadvq82luZG0jh3qbMLH0hxc7OswOlHOAIYef
LYro6t9GobdfTnNQNwEyw35sLkRvD1uXMlkieGZ4co0sz0n42DdQRD0Zg14+UZlr
8ENhwnHWqzOWbn/GrHGG2T09oePPmtlG2QEnY12onC8OBKRThiQb3+zElTKqqfc0
MpFtkngRC55pWj/dQ6nRdnB2CCso3T0hf8jzBeIySCCbKCxXotKgF8Wa/zqJfNTg
Ol0cXjsKdDNG0PiKl3X2ba3RnJz904lVEMjcf3EunYGv4RXqX6RlAMzoJB4tbDRs
7Vgh+ijerqoBFYmHx8nJQBjnNsHHBFwwGxTeKvTbbalBq4qfimn3XbRvoRa++VtJ
uxANJAeFMzVj2RD/1lBm7N5HTX4zzrZdtEgU+2IZBNP6t8jqmYHFpjab5A0EJczp
nVvoO5GgGKKiRIMSIrEmKbWfJp8LBKVdvh905wcnyQX8SmexbeF8rTDfRYLkjsQX
lMVE6pgDGnqLCBpzHNzDdP2BNiHAIMzksX7Ff9zaorSr3F/EgDXU1Q53IJNJV/jV
D0neFtLGHL/odn63pck2PsBNwTu/53pJQ0wd/JBv4ljZKlnFA+7MvfXMbjKX0rGi
IGAsqoOcO1wUJ/nxDd+6Juhhy1MJQFPbTBRmOxkBHlSQHY0uBz/xmtNijZfyBtwc
qf5BELk1gVyKo0YQLwT1jyy+ui7WCysIxVbUUldTM8+9olkk05xBVrtPAP9asqR2
49W9DZniy3Rwogmr/MFnsewTfYJPVNxA+QRedJEhLolSqj7Rr7RGUhJxbpVriG9A
HnTOMgyivE4mH6ulrT4gIqcjUpNH3Ffdns1Bgr2ffWQCuyTMcO55e3sN/pFXImha
nFP7v3r/t/ix7ydO3vjHSMlDlXY2NrmmOpj8XNhtr7dl5dcU3NiVh/5beTXFRZaq
1VJ+qf73NlRo2DeY0600qn+UhsYo4OmJ6mdXcsrMO+mjAzLEEWCXaO94hwveUPq/
eK56RQntp1xinwDMUP6crVljddcj6FPCL4rtnn7L2Zhzc3kNs6eC77EV1173Zz8f
LfZMtZrB1s3X6nqCiAsKp+AQh+n5PT1no9JhUCIvdNi5JIVBgsH/ZBdVmTKdBkhQ
3+4mZ8IASQCiTZd1y8kbPoFX6I0DMaOoOCrgk/HWd+4/whwmNFyrT5MxOzrK6/u/
g/oGQddRWs1Xv7pniGdMkOW8yoQHa8q8RAP9DREzFJuZmcRKIxGiOIpWccKiyu2Q
rxuH08i/f8ZQ8gvranA6CQzvufZUoX/mPhvZUuVwN0Dkbe5vLiRc4Eqz0DjQxxLe
nFgoKtP50HVOMBDvJY5xwBHtsk9O2Xt5zKmZOI6WQ4DloHk9P+zQy/quXQwTJk0I
PyTemkR0b61p+C8Prrqj5umMz+2/3oAV2/kHiv+woyVVzXybejn5fiwZwla5kzuV
5lGFZjbPOpv3vp6VDJn6YOkU1gQHJjb2ahzqZ7sAkJcsAhg9o2M8klZjgJ8WuH/g
8WLGZfr9KLTiz8fS43LfW0O+2v2o3AMthIA7SaNtek0putGCZHO0FmgJ9pSEKV98
7vQXMlYPbSZbPxW7TdvIGEvLRNMYptjqUFzG4QVxGxiS9IB779n3qxr6mXSUHciz
G0HCdItb+WgDiPZdbd8r11wOT/KOwGzYp+Lgqz+1HQcc++n3nc7lOxQmRq0N8t/4
nJX8OBTpsmsqBWLokC8diX66aYhcBsyEkD3top1NCDrVF/R5iKoCfJVLs1vSNWbd
ZeQco7vWbyOvI2sVPTXEQs2VCzfURz36IUq6rNBQMqiZ/HtB/Le3uqqUiLKbfpGT
i23BYn0h6yezSuHkWDRe1PrToJlCr+qGwGjy+/BonjGXzBS9JK6PjHPS3tBo2+BN
MaYTiFObMsU16Um5UNwEsKqUc9/MCfMiJDO2P+JtJT84TbOtYJiG3nGMlTJd7pql
ohPu/+WptZ08lIOFOakwANOQtU3yjMEdX1Mx33l2BRkLAf5dnP/5F/+nMYv7xoLb
FLj/I94gH/uTsT9sVMrMzxoBwhp6cSs0WCSSA6W7ksQ/4wvfYEIHbTIWvWvWWR4z
9grRm22J2C0YRQMx4sPN163d3uQLU31hPS8poyVXTZPrDjug0W7IhkUcpM6Tmmgs
oo1izKViO/B3lzRoa5VTIJFR9xob8QdQN/N2CiCguCB0thAQNYPai5/Dp0NcDLUC
+25PJz+rHhC40ucvgYAG9+UsN3NGgcZ4/a5T1dStKCmuXRiTeZq3B2tEs3Ze7l0U
9LM2Koif5bg26KSdKPQALI3XAszYDtJ+tnwtQ54c+ACoC8czEq8msuO48eQVOMy1
w4Ad3KB2EP3A/KfYaNNAl3YmQtD3nNTaLqKKeDpU0wIv2zaoXzfiUS/sNCdn8MTo
FgnobNoLDBR8oxXVJqL+Mq70gTnaCLSkwiIyQjhzmZ0fWh7u9NFGUptK6sV5tL8g
sePS6i7jNiADRNLm/plscQ3aFge/HKfXZ0VraHZNW+r6uBUCNQM5jpeVG/1wAgh1
ZmiGGvKHB8w7Nv8/0BEeFvDBGyB/smo9uKqbIjqAmlakAo9EUNrViGb0OAB+ivR4
2H0zCkJwhtk/w0M80Jog5vGR84FHM/jRRo3k7IXVSY+zF0X9GWXTw4sXSwQdRUlh
Y9x/mLS8dHnELParcJcXTuh0rzZW2J2pYEqgj9UPC66MY1FcFn9+OXkk20aCbeVt
jLe2Nhg1zRwAP1nV/vwVbBtkr74gglW8smnCckuKREUbtHTQcbL8tM8YCk7AoxEs
E518G4LpfyhX6ndAIJUxAlrCbi1q7W56Ch1zvFWVb7nmrx1qQft0rk5DNEpOZdEZ
RUubYN/TXSUk91UVIp7lYUMJpwCQF7Cvsu6xKlC1LhrrNO6bckUVGnoA6fWbQMGW
fwD18s1dDeI8sfAXKOnYRpOy20oN57rABiMzIhHAr5Kw+mAx3FA6isJnjrzMVumn
o2WT/NDZ5oVYxxAGp/BotA3zvGUmGdMiMiouq8Xm75PYhbvVenv4F5bWjarn5+qg
Ag36Hm/KT/9F2cbRYHCffxdrvdc5f5EvaiLi/gtMAicNHM2qqrAVb0ml+2yRORzM
YILDTsk9BBa6w6RXnWS4hif85ObNgsCmkL7iwIO/UD1e02CWzbiUvyiF5Pzjo4YW
aX7zznDD+BH7CwXISVB1YJBkDsLMxMMk6a+alUagXNCU4ugXBY/M8fFvuOyGZHjs
97ryB1f5MzCkhJPTey3+OUXTbyedIPFWMH4zJFn14O/BM0Z1Ht6i1ONZnG5RYDsk
jwoU2N1cyaIyXRt9LaMohnJX6XpTTyStQAmR0RERkMZyy7Pxnv5ajyg8fTZIn1sl
Y3O4fFx+pEmwNC6/ey0bDyr+UPS/mfmyvuRdA11yFGzU77cb7LkyAn3mAA9bPelF
QWKjSwgWKpx9txrW85Ky1UEkN2H59UNzDRF31T/VEubuWCYNS/btEGPoSRQufHRq
tPnzj+Pl0A7nk0qscBCuHJyXNiiUoGnyR4xvWXAhxzWJHN7i2h3GvUHHs3FjZ+Is
llF1zyFn0yN856oq0hWSagLGxQmMEAsiNe5qMc5NwU17mEnwhjkvP5s3Wcow4Y7U
L++bgePJDsJ3YwS2HSqGqqvHyUdf57yGEpYlYDI/popRFPtLlyJaCO+gOW3vM/Gb
wARQH8GkCoXzRGxvrSp7+rizOoH0MKco6lpsv7dgVRIzrXkoEK8spQmhZ7OWzgW0
wm5IZZcpSXRw+yTQQMJD38kraA4fBDfP0+jhjQhvcLCaAFoUK8FZMETGF0zsGgr7
8H02eywLEnSdFGoxrCAP/hAcgPanhJYoJJKTcx1n8sbUv/2APZym1xTLZygwOX0O
kQrpg37YJDh7+2Lo2avwV81BcrTV90s5N1MubdFaozU6rsvnsTA+PYk4Z5p63CyA
BCzj0Y6OUljUJGuiQVFcIdXO3PcYidmpQ3fA7C5iREpLePHVe/nw8GBcAj7j05bq
ga7Al3toioClvCt0y0twYoKYUstye8MTqiOL31r2E27A14pK3+TIJkyLa0eBXeT2
z5wrkaMNnrCMGZ7ST+1jEyIjEv0g7vdJ4MCexf7gMm9EgKOcQATdkoqqLqyOJ8JH
n6WnknzKnPzGe8HyN1trj95h0ZvpdmjHonmFKKkjSUebUIb1Y4lSkemlgA0Lf0fD
Hd+2D7zcj61JuEsC5hdoaluOGD3Yog+WkYOnvodB9MRJ6D5VtZuqzaZj8naKRxs6
+ASssEpbozDQBVrTCzLmV82xIk2I6MO47vorueSLXaAWsHABKVyZ0Gt9ylcFVjja
qQgvUgo3xKQeDukg5fPrZnHW5kY3D+2nLikYIWtdFxdxrIDNSkXd9X57W2iNsYMI
+8JCl9woZZkX7H87wMh3bAboVSlBdZjpmgWSPwdcJ1yUQ4EIMc1rPmk15jMLLsi9
U9TUPpxwuvW1wk5e8vBbxlWOpR6ULdZI94dK+pptB+v0EajI71SeQFQyfW6Z3Q7s
99qtVSe4KLIIXK4z0a7PaFuPstoPX+XA+14BsEylUBP6h2ayprjGrviqTeeS5enW
z8i4aUXOFLZzUxTbGePWnC+hMG0Ak6EEmaayUctBUmRbkxpIixJSPO8GjgPqD0AY
MBenbB59Ax9irB8ttDx515bXjQ7UmC/Pv6B63hFwASdOVfRnIUe0M5D1FlfbBZ8A
acUeKkl7BcjVTLrKYouw6QyrzJnpfyYqzQlC/xQ3DP3AHi5cuJPeifTzQ0EeZLNV
eRYxot09D9OJ2QBkgsF6ECYUeca9CYX6K/kAhgwQVnegbs9E/ppczbbfM8whzohy
lLO7ybfbSrtvIo54jyS3mRwAyHyKU7rK8if+UPLH1K4M92qp6vZavIEhmIbhJBVC
wAgstWr1uHzU5nW83E565cE9iaQL+OkaTa5qcTwVkXlOEDwb5cgHv6swrTXaLCEh
dCIeSX18rLoQhk3E/2KMPjvOCzQoB9Au/cH74onjLRUzPlynhI8OCNgxz0U15CZ8
ZNwLkixwXQfMV8wKE6XFcQafFOnr6xjAgTn+HW7609fh0G97hFfXHB6FVEM1dzbC
yjYrAFqVLKRu0z2kcR/PV5Uz0Qphmc4DZjBHRBwOHTyhFNw+dOdh9z7THKUsCUAD
I6ghykcshN1LEzqk7tEBUsnTKFRW5tGqnUC/tovj3kwqqU/LehcZAMiVUwLD2NzC
pekm6QC18igSIC46uDeHQNpGcsaG4R/GMaub8FSvVBYZlqZIC7+nxlwvTPxsdk5G
dNSt3FRgRAzyhepPW3/d5UN2WXyHcSZ6BJxBtxoUhtSOI8D1kj68/hyzaBTuYTjq
Wr/kCPP8KIASZExfrW5eNJMIWWbcE0hJJWPhCtKaRtMCaGGAFRz5spb/DG9YUOp9
x8fw9RCxSNDv6+do2dE7sEJ8afbBhfYVkjxF1i4Mhwv/VYhO1KK2dl1tEfxnr8Ix
Dfad93J/TE8Q7JeYQJbv56rk1PSqduKgoxilQlQKQMHPioRrJkLdIeSlcnPAcnd5
fkYeqLmHAnt2VvqJfrM19AAfspG3W23QNp232euQiu9RmLqb7evhSQepbcaCE4wy
nFrJNKgaEDLaZISGSQhPFVA0G6FC0Kzu5SLEow7yoMJsX+O7NtZla8bN+i2jS3LD
jsMz2NQcuG6jSO6E/H/k+dYFEjmj1ddDMsN9aDd1gXDt80pKhupP10B2BWYGM3pd
qGu8Zee9xR5HLnsT9pwjkoB6PKr4EQRJ9US2RVMeJkrgVsa42aCQRJ5XBmOUC5DS
fcODqyZhSSvlab3lOOE7ko+CKiD8Bzn7JAESYhn+xjQ5Ayw4+Y9jsB39aupD4DQE
wZB5LtLWjteKMR66p9a7L8zsJkrWgcMPQC5ZZTMnAZ+Jk/5YQh8u1tt5CCs1pwbn
MCbRP/S1uwoNA+WJ1adUVYWUI+RnbCYtqiyidYSuCRhHfpLNU75xtWwg3ZaVrsGp
7VSQeYdPILdvEhdwvNZV/d8sQ6wcL5Gn+KrblyfPCERcEBQwFKXpPhvhue2AZM2o
Eh7MKupof3oD4wQ3o0PN2m+2wpBaJYZ+85waaleRBZ99cZ1hFpx6QkwryKbyCzen
6QPjVbLYrmKOC26oULKZDJomyUFHCQ8IpPgZwhRMgaZp3E6UuEINDfGqrIwTtWH3
JsRLL8hK8qHPXYoiRGtzcNr43xPOqEc5t82TtLYNbrmdAV5J2/KBy7/R9vfOrS5U
hpAN63+wKoBkR4NO/yC81HNLLG5mPVata2PyctfniyoBssCLso3kvdwRGxUM2N1G
xNSp+A/3LXQdC9uq4mJ/+EebxyeE9Dxc3+mlwbrW/lAgEzhb9U+ECfy2q7/M8xqc
BC8p7Q1hJSElJbrdXwL37EWTBhXkk1OKaEbMGPWCVKITmJucEySIwJpmwGbEipcv
MrRgPDEv1WUpOa7F02C3Z4NLE4dSF5KOTEVqlqz5gHLk9NQZegx6+QB6tLbdw0/J
9WwWANaqbD0BnMh1Fn5Ufh2x28Zl+c+bb7FXrYsqiaxLvUTimWjOW/8e49aJZR/n
2/eUdlTkU6i4r6QJFiaEOEj5wmlYwOhsu2eUg0l2LpTuNwlIsGmnGzTmXMeBVw8B
vSELe4e9G+YhXrqpkPjo1szc8rlEWBTKkK5e+i5u7zrv6+izje4XnjocMABgTwfe
tt3qfKLaAdabCAjTpjGkYl8a40NTm532bK5+BlP7WTcrdLQRay45EIZkYC7FLGbJ
Db+hpKIJOIcB8IsGsmfe/r3C8F5wIc7Nin6GFtKiYkiI2X4xEbL86YRlny04GfCx
knSIlIsOieWKV98oUCn4/6F2yxzrIIGY69V+4nmAe3jP+1TirvVFYQIYyJ5Ltm7s
fA4JodeoU5tWdFnm7S8lJ1oAHvjeEsV1ZM122DzLGi5RokCZBi8qZBmC3lD9MHbt
QJZrc2yXXdoJThZNNJORHqRUT1IqhNLkXtdZy8hoIxr696h3z+YQcTVq/OWSrHQ5
T4nglUuOFRh1QWw+Q08Xfn8nS1kKVE8IRSqc8vowuFTUIYR7C4/h7R4FIPlL19e4
sSrs33uIgyXZwCRN7kNWcjz7QRViZXSjGpNeeYNyFvxp1NIfWdlB4Pa29k8C75d+
wsfi6w5q/+msEw3pg82tapHihztaqJ49T9fubfIF8mkdUvnfQGYA+FuKfDd28DvM
gdLqRfXoYPkvj3/N7v504UuQOy5fgKXwzKRyehpC08wtW5j72VITekR5r+BEt47/
CKa4mshV67bQionkA8xH0HynVepdmWP1aPzHh5ZYH/D0zPBtU0dlU2nYYVWAXfRQ
+PNjRfnZPrNmSvrQKuOC5jzFfRGRTwiVPGW++yjr8bsMD+uWA3xA4wcoatKpH3mg
4a5e1UOdFOsuMTaeuf/jfMuecdSEIw8RudG+4lU3lgHD1sOr+7KjULzm+Sq1MDCN
HbBXcxb83Qm4coidnuFjYOvFBRchWY75joIsIYsv9es4IhsvOSY3+81OJbJeWYn4
ySuV/UyTg7V2Q2cB1kKx6GnzP76dUq/9+TF82pTfwZ//CySpWkHZNdKWNDaoA7sf
ReknUIoSIECZGQeoE2DXjQSliIqLBVQr1FTxpmxUVt7S6w30PCI0uFFoez7ikYcc
zmMeONRjeshFjJ2QTuSjV4pk7/rl7va9Kd1ubO5gpT3WbPObFP0vTfh0Ozf7TE7Y
ynxhELF7FR4CTHP386BF15MaUzd9/prP6BGBjqxoPvyAUBqTcS8Eu3jWPTZ4xqRD
95yoaHPZ885sAg/RTMFApEgC14BTmVPS+R7AdpTMbuSHITTshcM2hGXZwMwFY/fV
P2ScjE/v7h0FikiguWd9rygw9Y6usLuweKAitmvxONxggvNQs4pO1qiD8uWrDQZY
oPgT92vnt6PM04vVJgKlBy+YDVrvrRYWUFvcUdPDlUWS6k+9c8dOa800UGd6Y2Io
Aq/l5HdzMhirN7QxpbkIAIOiuAwPGVeg+BR1qkLyAcrWSnwGf8+gE82Ypa2uiNfv
ziotjgmhMOyqHdeBglAEdNWlb2KbKr5WJUIYgkdpaI/Ewwviw3Orzk94Z7h5vwA+
suVLG1Tg5R5RYvm0TTYOASdr/bZ6KpDVaZJk2KbPtLEGUzYFyvvtEo0NKMHkpMo7
lNHsQjYC6lKF1uc6EKQtZpB8nczM87lo1Kjrve0zukOIpZpOCUUloxOdhB85r3k/
D7o5kXmSkWf2HaG8V2thAowxPMwAfNKIca8zpdmaGgpl1L66c/po4B1jIKqJZtWN
ohYtDxeP5+1go3lSqiicfHrMKqFj/s6JpNs1cWjEKoKG4oqQB+TvuTGz9xkV95Dj
HuAZH7THF1z6giRvs98dx4Z4+3HvvYm6agTC1n10pd1m2Bsd1Pg0jrsDxMZyle8X
Y2TUszeAIuBxxbQb0IuEAQdgPswoIKWJH+YXhBVTe2TppxmsTGSdrHVq764uU4D/
RxT4Bv0ApbUq0vEPXNrseuZjkktIcXYVk1JZlj+yaPEERqZgLkBJxO4uBVexqCvm
kepyvhBD1mnWJwvJ5SH2ajb2WWlsRu6x8HpWglV7Llth+a7M5zgHm3rAZfC9IJo7
EdzcpzjrPNwRgOHXnsu8iCLj7y9krpvS9qmfnTp87Jm7TsAkhhZPulxQKsdq7Ngq
/IdeSoXSgdKNBIEaiz+iRvyUpN/z/+Ai+MlqMZRcVhKszCOEnfwnbkM+E79/f1F2
LgzT+5aBAaIwZocuGA1F9Uv6S3m3iHSnTsXiRip6EvBDAZ8OY/9RtQ1ge7QhVs/m
urwUg5/fR1n1VRP4EOVbuficsqwLv1zuae+CjGKiGAzr/nrphy7ew5vWzhrSc4xf
uE0V3KfuHQxCRRjRX8yUf8T1dsRi7ySTeKtqHlW+27euPaWBNhMFrRxf1XboSMIg
HLxJQspMxiMcbwhN1SqAXu1u5TAPZiAHM529hfBda6aJAbabI/0uuswKQhiMhRRZ
VauyNDCl0DuMOdiaSzo0/nbMMXWgNzbJAzCG7audY00vunjsk02xCcE6qnIvN/Uo
AQXucbipgrSBC7K4kT4Je8C/XYkgauFZBlxDjjKHj8ZqH1VKDtbaeU0YVxae2QRE
ZYjOQM9nP9a9CXObWfX8JDK/RbySfpFWAa60NjhEjIN47ht+D1meTU0oP1iQtQHj
UzFxS4Q5r2AEZq+mvjLvd4OkgqSGNllbwRLF+tydezwreS2CLQU+0cHD4Mxv2Ofe
rT0zZGGqnT3ET3ZlMWmdTI97gwae0lVR0JHrsMtYjtcSnwdbhg0fX5iVGVXtQGUy
kAtevVfI8u+cYme15uEO6+rO68v/wV9DTcjzJ1b0isJXp4qzwP0dbVn2R1JR4/9a
1mv+ICcTLlGJgpQHUC4JmfNP+aHTSE51/eW6D021gx0p8TwDL2Qj7gaF9j/r+O8p
ZgfEl5bHlbKIxdKPiaYM8slzOncgRQfdz3dn9ao0NPISt0uxJdlnSmnrWjQLrxQI
F2U9hIJXcAg4SXwlhY0faNtBmg6jKbgaftuzwgG7H9uCWbekbBeGnOzK2CQ4qjlE
g12+LogLocDUOfWYv0gkeasyFRC02j9ccxHTrEdhWgkVA7b6jaBePcFnn7LGKXaa
KRp6QoDEGgK44vbvYZdsrSApEDJTBWD68XKS51SIqboGjhuHt4NlxPsBRyfah3wI
CFqZft3foFR+03+jswPJPJfQyRErVgWjTGE7tGMoNY9HemxV5KiUPKBKq6uZrdox
WQTDpwP8yMGvB/cBRjaa775d58g5K1djNlW6MJbkAveFdu0rXXxHq6VrspnEtFoK
DVN+g4HnKw2nq3TWZFoKwgpn5rP32tNlPqqIqcxDvSRpsPuKUecJB5IwPBvnXUuZ
SpaJd5kCLW3Wdcrh/v18uLKcANRRj8qCUCTzXqoFJ5NWJbE33oySohnkw3MR8USZ
v3Be5FNZ9L3xJ7GrsClpsvgxvPZIJ35i2qOvzG1RGHXlMy+7mwFnRSbUnZLR2QUp
yFp0rukbsiLYiiR60igwk+4quqn43BThv/+uMqA16bpmzqXsixoyBmqKH2xybne1
YF+N0MIL3kBLbZ3BlALXRkkkdOo4fX4AdtWuiWdUhnlEdOFTi9FXLPssDpukv9Gm
oZQEZs8+37Nyz1rPxn9U9mo2AA3UWbSWdLClJBX+ThaqlCIVbMtZwxgoH5xO8Ek+
6J/xE8J9W3czuItWrshelkYp9B6TFviznELlgeE3rxAZbueKjJR/qSP+GTlvZa1p
nzGwMseqiewtdGF/i8P0aqWS7iqlUt0FOB5g4WbZZYRwPPXAdpmUuUw5PSauUgE6
+5rs/sndII4Xw+Zmfa0fQmff9Y+mbTgDBzQpo0brTdYyh4WlQ0Cu4RzGZFs8vGu9
nOWyvm/vTXOLsl4AqJ6nzu4+V3fBhsPSj+ROYL0kwls5cmzFV6XE1aU09xdQjDjp
QLsvzWXW+4zELwLPLweoptBCE13VgUrTWf1vUh5s/2R4MNXan1BQcL0ammckDkW2
03BNYF+oyI6gPo9dZGCeMgUqwCkiMJ+VtM2uEBrY9X9Cteb23tUi9R6QfEcHkXdk
IF0hm65kQK12PuZhPAHwZMq0hyipRGuddJEEq1tqBKloFreiGX/GjfPxRVJUckV+
N1whSccOvhZ8QMQlKqz6RqHwoRwVtLxHq5mNCJfq00IiQuk49TbA1uh+kc5qlvvt
NJhWdHaZJpolLDpIXNi2VdZMb5ug926zjHAN1Yw2BydX/jnHm50xTJ+/2iH7bcSR
M0uTeFFyuIvVTMl7YiR0z/NvD0W8Uc/gFRUCy/aqe8kmgAbHexUA+gy44IxlN1JZ
bCWXLWb89x3fOYRUi86qam1MB7aCwKq7sjsVtu3oxQalHd2qHukorRFDfJHRF84l
vqs/RPMY2jcBtaLMFZIYL5Ir9Hvk6IgzT0gwz2UehH7pB3C5kj7iCay1n9jpSGGR
1tsv19eBXYI3OdwmTFhcQNaPDXGHhcQeeqJO5o4spNZJroxqa7zI/Xo3eUSj8R5c
vKrTwm//0r0Tf2cGfpahzImYkyvsyHLp6XsGOlZxkBtwe8m2sbhPTYaa1XaGo87V
sZai73qlgERgm1vleIkl+HNkWgk4W59N6HpiGQpitxfeam+grkraY62J5+nBmV9e
rZe7yevYeVnTmXKFvuChcgT5OaO2WwWwtniXNpEhnX68RcCPPHp2ydBZ19V0I8V2
7zgKKmzPP2GP06DJbysX1cDuOg9isAB8Av1RJha0k3uZG4RqAq9QyxkWBFi/a9j9
8s9uW9bP27BMUfnuctJq0/NIga1W5L8WgxX/Dzj/IiOKMs4nhZfscoh/W1GeqxV1
UVjBsQ/eFBck3gHwFHTyPLWDLtS4WiD9iBjfiRTBz5qcqu/mwJSZOzCfBHeOI/Ur
wnBg0jKz3wCCGMaxqbYYDuVk8q4WY5MTFGsQRSd2w8QecwwCw5I+Dv1qx1oIWoGc
WWzlSzcbGOgnAHZ0kY7gz9EWHJejJ5DVIuuihPCTglEfTGYZq3Y7Ea7NltTg5hLV
Jvo0QAtHTbfc3kGXgtbivbgOmL5BmREHAPLNCp1P5bLomiRdxCectAwq6J+XXekX
QBDn3E7K4SL5X+YeAP7TnZRrBNLBGlvuEPugNRy+1Wrrm2BVFKMQBa0fnkb/XWA6
ZrDqA+OHi7St92YQAtILieTO9T2tX/cP25hFiAUEWfBnH7xejJkYZQuOP9/a5igB
mW5SIqJnC7l+CazaQWMlq5s8iAq2YAGqA5Yt5OpkET5n6iuKPTfuliDh1e7dTj8r
TRHzjSzz19rPeu4FlcI++Qm/flV3xtMxC8qQrMc1tMlhsU7vxD22rAZeY7cDW0LC
MHWkkb++J0A1voj/dAWM5ISnwNdKLckpdzeCaABdegj2WzXVprzfdy3DNIDSgD23
XW+0OZaFvn0ARtZ9kzxLjfMyVhksnBi691EJFHZOndFA1mYF0Ml6/kjIt4OeqCk1
BfhRbCMaln2x5Gd9nXxBehUh8+9t7jwnNYXSchtzBX5NrnmM8yENKcXGBLOWaag7
jKyVmk9TEVhw3PO4ZIHBtfo5BP5c0QbGufLXEPChlOk/+Kq1Gw4kf+h3OZPAHT5v
7lBkGcfAsBk5GiR+SYap2wJJOxgtdAbON6LJB0Pt1/EKuy2GuE6AjQDC+gAohhbe
wzglzxEyIrAQIKZ4p9BSM/+ddeyyOjeUFKe1qIEhgyrdmtTXtEQWQKCq3mKbdBWH
wh/Hei31PPB+NHKO0xdxjiXqIuBvoP1FrE0bK6HMKzsXnTGaq/BZyRYsl+Smch4m
sm8Umt92a45qdZYNhWIe6QvwcPBNQMQM+wWuitDfVF5JF2qxlOBQp/tL0e3xYehw
iIqzI7T0LP1kb9MOMYQdVpOvtxkVDipyhRqBl/xNAI3BEm/3xAhXbR0Xaqq66CHe
3vC+IFeF7KOPYQwAFNBjdHYw+Ib/owgRB4BJ1wD2Z/LBwjQindvkwYxGi2NCTTn6
nBWBujR3d30WXnGHaC06ix7np8C6FZ5X8SfEYIq1TnrNgLz7TdPP0BmIicbb1zhk
c4qdhwKr8FZgm6SAb8pAI3Zcej6trOsznEgY3Bt/4WqsqvkoR6M4SVYwMAntq5/H
Axx2bmbmfaFKUQYJkb5dYV/iJfcRFjCX49kQe9tNugh3HFU2hKtyx8M2BBXAbY1U
zuGMNhwtKTl4E1PbHF1dM15A8dEjIA6c+Iu+JAbltFSz2ht3wnXFYPixUuLhr5XP
RytJn1KzrW3tluI5DytojNWjO+LiS8gxAqs3Nv+Gimf/ZPm/DETabLKNNmJZw2zl
ud75cBTHdltaWG+Tiikr52Xh0jQi0cUuLXOiRRdIZ73Exoi4ExXEEnN5Omrldjnp
9/KLBbyade3o1USF5yVH2R07mb8/Kj2jIi40qqSf38OV0wfYaN4Qu/yZpBCWznZm
YdOqkEUZB+NZlwSN3bsVxGZLyRyQvi2pF9W/WrH4WbWDoihovOyjAMv8ZaZKs1Nw
NbMeul4l5PiyGhmt23DfC8G4erTkBAMGHruAcjohJTUzIax/Oc/i85Spjakqy7Sz
vg/44SnWzIuv+Liuye+Qtjnp2BtomGaQhinIqiIKfpBBZCIEW2GKeUP+ZL6/fmbe
yq0i0T4hN2ZWOSV78cdLfDMEChgTkzRTCHaWNHOJqnJRb5QU3ACH5sJdTkEv5ysv
6ItKijyGpRmn4ihz9h6IVzs41RuHojLyk6ZUerRqilBpLmaAxNjG9dwjUMRhxhhA
dUh+qSxnoBtEOVEt85zFF084G7a1P7cEyLIZ0yI0mRTwygWccc2XNArV1b/xdVUh
k29gBIHchKlwFt0P//cS+zvHBpKCAVGLEgRGIps2NLqIGlSo4RuekMCCRVu+VSp3
G5/zjSLhwTGZkGDLTxkrpn8axeisQtgpm4OuaTrxS2/Q3QAStMHMtBW5uPefhNh2
Xcrj4+tvHUe9ZWk7XtEyEF9MFwUa764EaECEGHaDCL0GuEfOZGGrG6aXJ41Xyx9C
Su6ZFGgmt+mqi3vYi9FgnmWSRDmMGGFme6venB3j00VaGckSNsjZy/ghjATxnLf2
QeLsLGmpK6jCI57r4ylMdOtgSVKhA5hwnjTETaMVrIYALG3YrqQnIrow5kTiPkM/
XbcqRvxfznhCTNl7Sjj9tcSbqkuGdl5hllxn8mCIAwsdzgmmxnCPkqkdphRJ46zT
UxbotQMCSNEjgx7+KGq0LsoAKdF7t5uJT4sMazXX3AWtXcIIP4JXsFWsvEqs2OVZ
ngJbRWrJhQbkOl/ONVWLtMX7zQmZKPM2lmJ7xS6U3w43kRhCSopCvt3DJf78IQyS
AOkJ5lnPSoxmR6ckX9dHzipIWacEWhSKwzGYjekS16pNAgMHx3xMNM7w4V382utY
E6mJyhWL/jf5AMN2h1l4BDtjnqoxMiox/sEGCRQplkZL0TQICn6qLvbHMTrzIzfl
LVZz0csfIBQxdwDye+klnJDE3e00a9Qn8PBnypk5D4MtDSZTg/wqazdSlNjzkFb5
VuCjmF/RDHXDIPgtuzKUG1tGb/oJC97WdyOwvnk2EAQ5JcioMHE5up0O7hM+5I6d
aPokVMRLXKNE5LsEuvUYjtmiDDOfXVQSfhWG/n1PiJ8aHWDO5j0XXMeKBjlqki2T
NF9VZ6alWBglnGpxgbdX6AHYYCcVYZlKRf3eRuG7ebLiFyTC/KqLvjDYonO1F2Q1
GZApXU/wzrf03CMGElP+Xrr0RCA5hClaGfWEVGWyoYb87Aj9K0B/b7cNpFieynLF
D9CJ/rx45cEsdp9UzCAFzNoRZDZaE460byWC8PELmiK53s81rJY9rckXnhqItClg
cIMduaUS1eO+bIu2bQ1IiKg3mIUx5zOkJgsocL53tD7Z1HubzQ1m/GGVc0VuSxap
Pm95vw19SmeRaV7GTGF0zWrdazzUgdlVyhr3ujMC6GbLFgaxy0fMKzpby35aOkJM
Q2SBVMaCC7XNm4ow+RnyZlnG0TIII8ZAgL8pgLZNHN5VGmjw6CeNNH8zkfHMGFKJ
WblfFqOh1fUPKo2v/n10VTGPdcyUzKNDplfUHoN8SvrU6IMZnVK9obgOOGvSjvTN
X8AlRJDy3uqtAmZCJOK1+b+HwhUIWabvxAJCnAD/RnEQiDhM5VFjkBik/dyjLUlH
C4diJH0k/w7kuSOFEOzDqppdKzJqyqfwqDDwWon3JBIaHLH/0iY+I/suYUNUDtFd
a7ATGOJni8V1QvQ5vc23b717SkJ+5huUjyWX7CZRtndksSuYc6Q8t2VYNftgMUMz
vagBYZDe/R7QcEfjL3ipAjDdMio49XAvYOsigd+Sl565LbO7iuOcvIkK1vIpwgb8
6rVstrumH53nXSQw3I5RzqyY9T4eERlP7i9lTsTEerXQnIu9BqMClFr5lfnV9ruw
IgbT5ZrgMFwlVpC8z95Fg5zqmzfaJJkrgGMrVLaT6p/g9XKK/7cN/EUlkDsIBAQk
Pl6olJkEFbkuh+s71aqvr/TJxbP1nEXcnh7pt+jpzcONElPKpCbYqZDMoJoC7Qui
0ir+te9RTzQRsDhBUYmIUyOvUesve1B1vauk/b8aoVR9bb+jpCEC7SbeggXkOaHz
C6JBr9pXgaZWLCU2EJAM2j8i6gmW4nDy7xrk10aAdzSCTxHEc7hhOv+U5vz0QX9B
FVkpKmUxb5tjio+IfxrA2olrSJF/SlzbEjPuzs/5oFsJVTSTFqNCKcNLjVfCG37B
idJWv5S+CtfLNkszcqUzTUSnL6iLqqAKmfANVjC8v0vkNDVlzovxchxOvO+mS02z
hfGryN52OvsEOG43ptd7hCyvj/0q158jKcEAtyW5jmkZhuOQcRQYqAH0ZycrTwG7
psCab9QIp0kzjzjWfiAQqgFD+oDQVr4iAFgnzYBz8PJ1GaoZbSHkIEOJe75h06Qt
T5ax12HZYB0O+K9NYm5YoyPimpTZ173B1oVM1O8H2QXs34rEwx6IjrfqGITbMr3U
pY5+UJdVIsaQoE92z5YkvacUyHWHX5yV9rHAYvfkrLfYTKJYsvvbq7UxvRulyIou
EkD+4Ew/kGF5ovngGnjcJRNfjCrsnoTifKw0FPVMLl0HgEAXOcIBpzR/awIKwkeT
rHOAWkmqDXp6hLQY5x0pxAOCp0Onl4eII55K9lJKICOzekAEg8Mb51Fj4Hi1W9aK
rSzu58QyyqkJZ8D5jL3Wz79+HQHo9J8O5NjReYm9Mv/SQ3eWUERFskey0WGNIQmI
z/Do8wkfRlJj3jwLtuRvcSRWl6+MIwxKfWcJBkgXBb0aRDBoAazRxrkStmhHAQCf
ccAyyijYVLex8wJYXFU+1lSknICCmIiK4BX2bmWtr7wW/8PS5p56eTS4DogIAjMi
uxv6DW2EdAlXdrrVFD2tquU9IGa58p+Rg3LREvsjHfcaT9bCxtrQYMDWdexTzjGn
uacy61LsKNT1XSio2Yq0s9+zomif+1pUchif2B0S6eFoOL0+hKILiZjS/p05W6mW
YAhAAOsYq4WoAysnhAUaWs0qFriqjt0rpMbx56GCS/84/+VX+bEJRTF5mY4baHqo
NAbIKk+SK10twKXwlanHHAsOVOHH9/Vh3LmXXQgUIIATT8DWYqwZKoc0fcJjAv41
WK3e8HqwGAC4XcAWf4VhT7rDjbIcjstFVrfrm+CHJ6NoNNmwoeqVdBn/hRbTZDIJ
aajadvx5ZBqu7SrDttfqQwo4degD714TxEZlcGOvX48HFvvkuqmVDWm3WYDcaouK
9h8xy6zr8bekMfToqCpSiQ+LZBA8A5ERriOlsfpQtjMbg3zxVsJo5TUOmfjSQzXc
RtLHHJoHZEFFLYMTWHt2VcR7vZaRIuHiBsf7Gqb+RagVHZB06odRKiuLlRsX+P0c
LTZP7riYPlWNSzsj559Rr/dbi+psIhVxEHBCcReGS8NTaxwwqC6JT20hygSkEWgs
N7xF3//opbKVKGBhfKRKqRM47MNJHCVstxhtYDCmW9G00VMoK67986tb+aVXUM1u
npVBNFZHaavuEE7xMht/ynA2WAtVyg7gCTPL6mCq1ffXI7C5OTxTP1C7VRP8D97O
TSYeM1p6vs1XSxIlKg0NGGcW+49t2QwgonF3/Sl3v1X2SltxMaVG20hNcYA/xxpY
KEs3fIkhxORXljV7h72DKNchgddpq2eYv14eEZBTLlxq9Fl9i2gB67/pK6FDZ+Ru
BJZbVh6GCAaIkCEThIONO6zYFRwxlIQN1lGk2/R347NEiiePC037uXClTts4bVQA
NDOE50s3Hv6RAk2R4nyO+D92o6UR7gr01tVhPljwIJ9jcVI+bM1JhTWXEYQPrhCe
4ZV68hLh3asnggy4UbiMfSsIqJpXc70SCxYBEtBNO/syM4new5A2uebDdRZBzsVB
KBiSThKjk/zoXPBK8tsHQmK67fET/I5oVAwdtFlJT0cxu7/4pCxqh0IJ3CNXfXLl
dh6PWM9W0slfSRciSx06L5Em7W/Ha5hYzBkBOapOm+J+s1SUwppavF7lJhYopU7i
A/gbOlD4y6RYqi4BCIrEFw6dlxWRQECxi99eccopfkh9o968NOSWWMim2CDIeFyk
ABLK6xsKSJAbwPlqCVRi/q0g9eBGK1Hz2bvaQJw3bk1eOXyyrv0CFIIGHJAtOnUK
W/8NKY+431ZtLFazrOeU3HK7JcCN2W/fejR4s4EKSaRomeyjTtG3A67PONPGPRp8
AbjPuHo+7ClulFReACGPwgCoyKI7MjGLhdTgbrHQoyk9QakR3pZSB/ssxz6wwEM8
S/Yv1UOlS2qgDxHZMilOi96zq4pJ32GEMgkRhw0lw9NU+PCChVRtUHA9DKvcwjR6
CkIwTAgkpBB5W0N85YUj31lHxl9/y2NCqO4AVQy4R6ijK0l38kEsQG1lfp6dRp9o
rC6cZWKI1p6b0VIDoVIHdcAkpGR5gtqqM66OAoze/kLNFFe5N/iL4nyUSJOmkJPN
0zeNf6NkGdkXxOZN25TGNuwTPZYRjPziDXnxldxbLGTsU74O1wFBAyRiS3JVYz+g
2GSA3ahxFOIckKd1ontm+RF9T70D/R4lMzQBEMKuD9D12ZjthN65ryRsjRZf5rsw
D71XAHAXhaevWv2ZVGHVDa76ikmyZ62iCTYSps/ockqlQ0rHJSbTUN1Kuo3/EIUy
GVm5Fs8ahieY00VVtey1IjxxpsyiKDOwBfOfPYnsPIgK0RVKFkqm50+AOfclusk3
doPZVZwkNYUQZ7B79UTEXbqpLKVjsthoeNg3T16xWmXx7RAugi4JYET2Dju1d/xO
OvEYuXewkmXzIHnxucyBa6HY8v3k5OIfLmamZ+sKsajX4bfxBUEcbqk5DugyZfUv
WZMZ2qLCWJ2IdZV9yuaCwSl33SytAifLMO5jsB0fWeJiSYCGT4X2tZ0wsiJkC5qS
645P/V5BTC36DHL3Y+HiXvxAL4ItmsQPeDJSTtXkivNvH96mtPpF5kbh2nF+fqGf
k3hFypyj21cX9g6Fup9a1ytt/NBnTnF3F8vPNxaKpbv+zkm1lfgVha/9BcQec5IJ
1tgJmQS4NZsV508Og7St/FcgQB/x5q433tl+iqXw3PG+c6/Kw0HaIyqWtOM4Kwd7
5FBw30VJNwNwt757xaQtr0qWlGpX+KxqTVOTYllB1vOhPJmPTofTX3bUeRDi4TIn
1JWGVkwqGmGYslnQwlALWUAyzfFTqI/22gbjAFURJLrEuvyYLDnG54HtJTUSMJRw
QldhQSH/PehZ7C6VzZTFTaKNGtTO4EiOFkPOBjIU1NRkO0Rc+5p6c/IZP+xjNywG
QPI1k+woxhyK5j4E9Zl8pRHDW/aoIthWSYpvda54bgZaljqOHeStw/I3hSsW7T91
aLTqDBn9ilrN3kzQMbfBxe0W++FMOonhbF8J04UTFjGquf2bfmZPqN0s3HJFrH32
ytcIpg2hZpG7O/AY+xy5jfDEtzmXH1OZ/YsId8v5pyXWW2TZUpRjYUCAr5iBKs+t
7yLdSjRSJCirWfrzf087BnxeG8VnrGIifbGeniFW1GFoGq7P8w5RjS4gCfo+r7Aj
fkhdFDkoInqWeG60QpuWb0v1K+Zqd0y43P3HpDRH3wS/MKTM4MJnBSIxcJc/u9WR
G/2vjE+K93fs1Hhhdbx4lFTkhuPQYtgfhHfes6QLrpCSZ1SxlKVQMr0Hq7VXrYAb
ygH9V/DJYy/AhsmwqcZlJ6jFpPsUPTvz19O/JD3hnfsBxQO8XGMuaJA6CyPqIcqe
Z4n4zdAf1T54RQaCx3XzwgQ8Ec7Ami9I97/97qvIhgOlMR/iOtzxbZsSYCHT1P9k
+F4zXYo3u7t+XXLBf0Sm6dzMDQrwXIGAPPCqWidgqSMLLK/wKExhQ6Lwetz48LpA
lfopFWIoj41tR1cNiMSVadMVK1fwvBJkgkMhLJ2X/PmyjNVVUMKA/wdIyeEpj1L+
JPGrKpOHDgWmvvtQUJsNIn0QF9xev8g64xvqJCUiSb80vivw0kEc3z4w9ybgUtGW
SSKpjg3uUbB+SzmhOCoXTvh4y/KQyKknWy2HZmi4AkmusCveg/B8rgyGny4afMDG
hnc5VWngSFGtXkeSz1SHofIEq3G2rU/CMFnHtTh7vGWaK1G/Mktkti1hj92Tbk1A
Y5z8qbzZvAmnTG8QolyEf8PKUBXbHDA//EHge50p86KvEalI8S6Z1iEpaPsRdjMc
/9KhA5IjCTMc0e1niB8fT6pej3Xne8z8+OwHqTuO0vTIN1ew77JNMe3fukJLwmu7
4NQGceuqXLhZw24tgC2J1rJcKDGseNxFvfMiqMzTmM7sEhtlRmVLQ5HTUuHs9TgX
6x6m2vDinfFdw8EYMOmd1F1Z5+krV0aBR2I+Tr1QqMRv0crvXHXdG61xOoVxFHul
ksLCJ7ZN1RwxT51j8xRY6YW9muqPQMUCCul3YA8iYTgz4VYHVwK1iqU0n2eSLavZ
vYzDf2CvZrEF4nZer+YHB3Ldg804PGhxPyWc65FA/xnsOg5FBZJk5+LDYDF6CuPY
QSA1G4DfoD44fsKaLgyHMGkN4ARy0uN24MiuNmugMKEnkeYouSDNHg4QAbEK3lNV
ART+SvgUVgxnJAhcAaxSiNjK3RvPARF+/aok4GrBKq/K61zPkyHchd2JFY4OJ1+r
VaBT6xbHDcfEataSBdEDPSTK1zplyL+EY1QqyLNa1h5uXFA9Ibe7Uw0jKDtxfTBX
aQI1g+WaoN+GC/ljwfb7/saCWJktfk2JEi4APp6RM4T/YJMO5Kp3whm0X0vbFXCa
ID8EIZHYichPNcYVsAMPxJPlGnBXrFNUayEnCcR74IkaRtS+UMqDd/4enAJRrXAZ
yp4hxHns6J1aNIwjhfhoSoMg3TP7TVWIbE+cmD5lE+v0yCLOmauYH/5co8qv3TpR
x77wBwIpe5cXQrYCGyuNG/O9a4LMP/r+RXY0RO6FO8CLeIl4fT76wl3U5uMWWkE5
TZY0rIRxYTgSgDqvBDmCpSUxHN2CftzOIk51ow49EhNW8zZzzUQ8WSwHFYTANi0y
iA/tj3kpPhGs6Qd4iPw7SZaYlQzVA2OlGNQdTE3EyDiJja50G4lP2v40AmWfGkau
4fCYlhgb2YRhJdoXKArw+0lTtodXn5HPC7s5J3V5Yju6+cKBKwwpfnExZBJDFdpV
7gqemYLwGXfIwI4TtajUXhljIRYZ8x3A+ctWo5akdR9cCocYkHQ8cz0+2kdziW5X
GcFofeKDKvYaRCUd2Jks9/k0sfI7Ru39ihpgiYRfbxZb9TMZ/AOKU6FNu8V3lWoD
2SIEU2UnVFJBNayKznDxZc9vTb/UvXHvK3S9z76YgGWi5Ma671MywX26iurvfrsf
Tuga2qrWJ+nbi9K7qnjBcio6QmZghvFViDjXlTACyYv8SsPWQrVpaNi1Yditur84
ahVf70aXT1e2tswscpQhg63Vl14/HMmYAP6OO7w2Jynid2tjI6ZaXdwbrT+7wAaV
zLrefjdNqvrSo1IG3k4pSz4Pe2haMqMp1ceP6+JV4NPt3MLZ2bcnqGy92d5mrLrS
U0HYMLyyJcpGnDUkxQMANoe5x/9ZpU4CW38Q0tIz4oU9dE/bN3sxdpHH1IjEerLc
m31Z7A70peySNwFfEU4Fb05b8Q5FIm8mh6YyMlflQhziS1pf0sRkZKlczciARMP5
ZwpwO2k5hg+WNhDYj0hHhPTNAVQyJ0eqimwPmqVvTpMGpxu7C+aQA5tfkXik2rxb
gyLmxPVj+mQlTe1pQz18kVzI5b2zl92U3ScL7cbxZKaSd0vroA0s5XMQ7bq183Si
BKihYf5MJqq2NNS1cosCN9uXc/FQf3Gfk4SzHTUX0a7toQMwu3HOuW+Ky4HdHRCO
X4d3eadUji1CHvyFBXzflSbx81NsXrfp+fAqlkI5BCWD6pma9YThxKYtKJB//QHb
LnfcqE/FvHoUFlqqJIPrmsZlv0ONormjG5xusC2c770S1yuEL4k8U2WLmTXbMksN
SNuGD7jAsBgDH4u09DWLEdjBq5HngJ3aSY6vQ5VZwh/cbM4e7+FZjsWtgWb6rY6q
vnjSAjdbtejcRQ3qCyDc7uau3xkB49lI6tdrLRDyYE7fgYRKPfilIEy6v+bcclW9
JB9Zhr/dOSB1CH0NFiLHwI9ZnPuhS5L8dGr+rfmwRlN2802Uj7grJam6jIR28jGs
vcT4YK853iySa/+QzvafUDKvLTXvacvnnN5vj3/TpO27ZfV/6tcKPsIE5/LtA0v1
coQqpQW7TlPZtPWsC3IvzLJc0NbnfqWdx+qOBn4vxqPc8/kwl0VtpmV5MnKo8DEm
4Ej4EIZVp92u6CfafQpGN8XBr8rZ5+1FPsoAyFzQ6wqzdGe87SdEDOehvpD/DmRC
n3qxL192/tyB0WUdYta4YoG3XCV2CESQasJaaWkcoratVDnbQixFLDb2VE5+gwOm
pRhh3K1O/HFu4BzS4KesY1wiuoaH08EzEpB5wc280x70Uxt3iW16NY5OS0Rdv4sK
iF49zcM75HeSo/NL2pLLE5+96+HqOMCAwC/ve6LLmO1kenM9V6deKLjDzb/CDLnA
exFV/56dcvjUyJ4aKmlOWM4Gj9IHgq3InSd7T6/deqUhMkTEjApxpbBZyfSCg7XE
YZPjZiAuk2xSBxhgsw9LZ8DPMNdTFnNtwkKrAMOjvroPdHqd9fExd02DcSGJDatr
aK7xU9c2vAKKIaHFSaxnG/2QC4zqClTyUWHmGbSwvui1AmqZtE/rFaXL+pr2k/Cy
oJ7oXyAUq+2qrL4XIJ1qQhynMF68OFYTayM73GQfMJ1rIPo2+jlajn3CMTmuOmwh
HG2yUAkvD1IE9G0BS6IGy71Yw/lEgNUeYIcPuza3WFlDdpnleqx4X77bEsnMG8FY
ILx6sqf/rtagfCEI4vVVKumdi57vi9QJ3h51tfHR7bFf8BDemeI0UgYtrvDAjTwi
yBqsUvUJJlc9HbuEaSR1SO4dDF3CrlX1BmH2J4kMshoASD3jN/9wgAtLQTUNdwUT
F8U6PbptgHSFAyuPZmqvN7kppwXMmaLkDRYjqkaByB4S5Ao61PUU2UZHCHOqIELz
JNOADjtim9pxENlF14rrCP7459HYJW3HDX/ymDcAEvcOe48mFLLJQDAavPtwhmTc
bqC7BZba+gX+S/Hunp1YIfcqG+4VNzzby3ztocPUIdIm3KfLrPmpQBvNaQr0HK42
ujjLdC33MnXuKbFVrEPaDl+cs/298JKpFXiPbROrgtVNtIqIu3O+wKeSdOZp69ys
3ZP47Imc0l5VOOwy8B/3SJ8unAMXw+vL/19V1lxrYH+RmqzzkXMw94MXOmd6vC4f
0Y2XJuukOO6Zu24+7im21Z+OIg0HppFHx870+a4IHPxv7Pf5GvoGPXts7CtkES3v
8Eh+IoBjTFJffqf123s4LitJ71MbG8xfpHnDZ2MauLGltGiodVgPKAZi94b20ePC
UHfvewww3nHcFesHn+7m4jZkxy2tQKXVmIEVh4F2Vxot17UsBlKYWXf6rDbRomr2
QpBRsDsy3euv+XblvZFCMvjXgIBJ0Qg9IPMr8FS3UJ0pMMrQK9SRPmvZkK6VZ0MH
7tR1Cdm1DuR4+WtBIJn8v2VCe5Jhp3XBImo15A2zSMTrmHbyBz/g2JuNULeHEHH+
V+sEV4HU/6qJkun7bzTOxsqHO4nV4Mq86++GvF9wJha+toK889YxbWdNt0oabQJK
edTlsewX6Yu4PDhCRlciGg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gc5qKg94wChLdHfwPOBLRmYyuB4c+gNWy52wIfMFIcFcL6nCKkvo0S569UD8HpPn
48urJGQM/Sga2G2wGMGDDW12/H1FavY+vCaLMZdOnmqev0OL6qDIx5UxHiJNiQwa
tJIULJbBhgEPmlMoQMzMK/mzqVywg4HawBpk9BdA50i3/FZ6X2MIQt4OD4inSfjO
FV8KZbORwHBjS/aAVvjigrzBTyn+CsmMJprvj5saBZ7wgK5l5K9oY4m3CI+jsB7g
qbhzBOR7vmpM3PG/iiKmViPauXCY8h6TvyeDnIKvmOPmNsopmnpc1LeNC82yxHus
XmlwF+yAcQ4HqJZ523/vjA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2864 )
`pragma protect data_block
BWPESvlsQtZ3NOs8amuQ+qQN5i8FGFQbUwcGQ/qYUcsGvKH+/jYwyZbhWbWpwKv6
2kUHbeolMbRecHOpM6fVuemplqCOJnRUWuXriYcdQarHfeQxO4pi9G9hyWSjlENR
HPlbu/VQteWmu7CoMGrAcBKsbJ/56Cv2IEwSk3mHkcjsx9jOlctAUJWt6MWb4BSt
6IIA0Dqe0pmr04fT4NSs+DOILqvAPrdAFKolaBGmz9HV/pPQHSLcdAs9waxr1KFL
F4qV387Y77d0veLOQxrVEzyTIUu/SRrP8YrOkYofZjJPdCIZW+L1Z6MwNdIBplUq
GFoxB6u/HFpPsZCPt4OIungwXcQYykfoifBQJxN6RMih0bEl0uvkZkUCOJU4sk5B
NEKPSgwzrX8c/JugWTaov1KqJG2AAWF8FRJzR48IeSQavkZRaXiUn39qrB0OD4Wv
Uqd7YAyBZRxodOGid2UKPDxE6sgiIegooIdVW1LZlYAwdKY/0RowviEC61Sby+xU
v2+D9s+T28K29K+Ifnp4obfgcgn32CC1qp9iub6idEHbmwB9ZMYD6djCbdxrfEym
RyJXJt9X/mnMqrLDcR2QOwqYEBNi2fgoawOCe/AYG0i1rJkYhJ43pu/tE5BuzL5B
YOKsVUGhjKB3JrQH/uXdRtTRYJAJr9etXPY/p2QtCyAD0JOh4QPAvVALpJmK6Zak
Rwz44skYRP2Xj8EpRFfKeXkTygCccMgtE5r6dpxKYwJ1NIUvPZD80oXfhBtGvf3I
nq1HlKfphZjLL8UPYljhLweBy5yStKFUx31d1D9ZULxZyTrlrE+4tvd/X4qup9E/
5Y9ozR0FTVbACmLPm3TuK2AHAK3lZfxMwJptTtPCV/8OALEP+gECIyKUJpob+Q8b
ktQX3EQEFD5X7/+gOLFvhocvPDFs3WCG3lbBJ1yrKwG0y2Tqxr+o6kNconipPpIu
JCuEW1369Tpa/LjPX3oRSlmmruacB+ViOKQ0OkBRdTrItSxT6cubEdEZ4d2pEoE7
qYwyx1P1Vu61/Mo0jaeuymZwcYBeIIE0MzWidXo4usXq05qcbcz0HefZNJCozO0G
gcZm+ZWRQwtz0vM5UNZhGpvG+uk/Tm40bz89w15QtX+jeuhQE2VOFfYFEiTVns+N
xn8RPpprf0sR2aEWM6AWGPddA5jk+ekWfzjw+2fWLfHls/Ww5WFdMru7f+s7mzTT
sNHqIHTMptFK6rkGvMpWpFs51d65pnZQgb5UeyB8Xp5+PpfrnXR4XXEBw9YUKNR7
UdLE0j6HfT6gSOdGABe/U0xY48oulLu6wPbRvQO6QizW6lTctdUuRypzyR9JdQtF
IYhjL+5Q5J1QPxRrOpGoDHaykCt+B1lJr/Z1VOKCcZSZTt2WTrIk4YcKCWMx8I5F
GrbLZrAt1dBhI+L66ePRwHxM6ZsON1E3/UGwUyTeI79rwRqBvG7n0PjDz5+KUVxe
pKmvx5IoxLJ+xMC55x32wTtrz+dP3VwueRt11TNwWtIBqM7RRV9n2H24tegx7MSO
mg8DrXF23nHIJvyEDthfCg7B24JutJhmgnD0EjDN1bzvWoWuBLbBiZHNzM+s+yDT
GN+7DM6fD4i6ArO4bLqYsEggPCsFqFLPjj4cFxTwKR+5Mdg3AF7ITCVDciESVN6H
geUw+B+EoLW0L8zLHpgKCEFuQMgRRGWIgXdRZ66ntFR7KFC0Iy0DyVon8mqlxe5F
fQoDCPEtwBgVjs07SxPjPVvY7Ok5lGoiRAb6My4itbUbjQXUs/MP9odgYGY2/T/P
+tcXB+4O9xi0q0qIsg8chIq06xSYWQImb2N+t8knH09bPK6ozGgZi1miQBURBefF
mZHiiwFjV1abGCDQyrmM1gobQgHGtWve+LYF1bVTmbaxRb39kiL9sb4PfLYKyt2S
Mw1EQ86reDrLMDrlwWQ5p01z+zTM6rOOknyp9+6/MxA6sCh9XqY0Uq6e7g9TjQy/
GL9Mq0HYfLetyDFH6pHFCrRvaaTai7Wlv5giv9yadYzowRTGQZRFfBLOCds1Zy3I
6BLS2o7tuNHBSxwqqQK4Y6EWwzvMq1o+RL8NhHt403SfeCErqv7MyGcF6bb523Y6
Yk1NuMHRbORt2/0Ex3zZnGDenqSrhRABaeZHgbjVMMFH8wzxs+WXGUVh96LfOk2j
6JduBh4m40t4gvRRemhJyvb95NQzTqb6+qC+fY6nLZUrv8uS6Tw0v5m9NMXD0E2T
0Al94gN7sHghcmX1udz41wCXkz6XbwxgmbyJGc160q17gkwoqt3pYb0TPdo2ngK7
Pu1evx7vBDZzglxkiu4L3fjInFpOM8vWfrL6RkLAR16tsUDU7wT92X3ORX/LYFPR
p6g2m/MeUkimDwNWMGXA7haMMNf9LPWzvwmCHI5uw2xg+c0gTWut2OxxQjNRhV+6
EqS15R2XwjwFogtKj2Gz2MfmcpB3t4R1cObl+piYFAhRzClfFrMQ8vFE+ajmS4Kg
nl4dI+sdpKTix9raGyRR9xLB+oGwZjL9fnVpz18frkRl4FCos6Khm8eZveDJao2w
kRQo5VSGfysi8slD/0+zuCxPUzk/dk0yVTY8exsruPKjUkf7aqlXzYwM3WXJ2crt
xOTccTszVRbLcrSeHmD/csSQGqk5MeBCvWwbVAvKm2VzxLk0RLI9SIEIB9iQfSYt
LHM3CSPzBVgyL7u1MEFk7s7aRGYpiPgPR7DCZM18PyyYomp0xBX2N3ocbrLqbURl
Wps88o3AlFPSCd+zRfD++Zsd3uTg4aymPDmE8NPkjCxgZK5yxFOAcbwtI47s+/9K
rvx/uDLAFrQQwD8cub02Aa6erpb4vz65ULDCjdrjAgC9EJvjfxJmgKflhpVO+oNR
3PkAEWtMepNb0aeoM0Jw9Uyz7CoFzub4ne33J0frHnEAVrYMKBXZAn8AWjMHzR//
vS0tmtEHR53gDUt37jfbK+aRqfhQSZvFnTBSEgG+kxLVdHfibQjs2wMjQcWNE5nF
6eiJ5adR59RNPEerZAehz3dBb3KboSeI2SQ5Hi7dVAyNXaG5NL0hZTiOR4SGrjxu
MXIOyZHmxkXyNnN/VwpGIA/kVQ1OPOpXGP4bK/G8LiE7jxVASczftEadBsG0vL79
hdfewHNzgkgt6ouMxaHCxhsSILw3iyooVtsF2thr3hHNXSjmTPJd8LF8qbdqhAr+
QcFw2gSSVxKjAffnYn0p7p9Vj8+sCz5r2PpcFnAQuhnny6YZXOmFQQX+rjtgaFcP
N6+u56V+fFXWcWXXXrmrk/wK9o7BelCv5b2ApKbkMyZDylNUML3eRq0Z/PSyBkZa
ZexeGlXj/OUxkcfiOqkNWl7pPgub4isk7VU4BGf6P6e3qwc/j15oFbJEvKFURQ2A
yOQ0TzCVWboOh3Mje7i8uGV88Hd3bqWtov/ErMsL+1AQrMYdnjEMMkSuNVshXz/p
LVRmeN2Id1rk/nIdYarr6OyW8f8fps4RtDx/QCkADCUVUFndTVj48OoKc7buFQs6
sEctJJkr+BofVToFCPmSESW6M9lJfmqdflOsk43qFaf25Bi3ReY7r91DEeDfE53v
yAMjHHsdrppU10N7lZ28CuAm40ZFBZTyGn1itx/rDKF+uznn9QZyLg9GQVFfO13C
HyqjXXMe9jwK1DGwWfVp/lOrupg034h6uFCT8rgACMmhl1wQkTwa3his6YY9Xt39
402un0XPzQFs9kNVOporX83oXn6qo3mHb+1gAC1FqXeBw3MF/atoL6qT1wIZv53S
sun0QpIaytiHNm5zKXQ6y0uQr+7Sww1IuuQ5HGhukCE=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JeeeCSX2kVSO4BzoquNOIwUXbksFcMUShf200+YTD2BUM7/7PGItnZagKA68LnTK
HWTqORthO5vseDjGyYRy5vA+unye+ofkN8EaYUgVKqEhtaU/uSZCtT68weH2A3vl
iPZDevI3p063mb/X8Ry8lvI03UVcUqSiZcOVCzlCYQzd7rucPj5w3Vh13ZH/aKGr
Pt7b5fTEIxdu4jfbisWg4bmJT1hHAcE/bjRSqyKLqH0biFw9TlvFvQ6kRZU2vYAf
7kqsPgxwasrTtvtqERgWt//LkYUqEXzrAxwEaWzjotUZ1to2kHz55duHpxxwU4SE
5wJG7LlD525HQ/+SLS8IHQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1296 )
`pragma protect data_block
L4ImQIwQWgEdWEpjV/XGs08ZbdeNV8PiqYJbtJoaV+8NrAnvroP5BRROFWb6Yxnt
nR3tpByTFqPJCQ5J0RLLu8mcxoHBMrAXAiJjlE0wTDD+Z+648VGqlaXzeMOW2yu1
V4w1L9tQfw4uIBSP9RGRVMdqd3groCs5/c7lBYVpMGI1/VNZ3jvG8QDTy2z6ffcG
suD7DBIIUzC3ru9fBUZjs5IAFXe35DxScQTOaRJ2nW8U9XNijZZoO9sFJwD2OUhP
QJispKq0ly8ZEpORthdgNCvfjfUHa1WCkzqRKQXF2sd5TMvGKQmXJMOWsTbZ29Ye
bcSDbpUuYSlOiCE2vZzK49Eye6mJRlZTNsrvAyIYChsAf+XfQWQs+7SzyVnozZv/
dduPhJ+4PvJ1zgdvvjNu5smsF8dI+tGbkbpXP17NBxVMOzuhhMwzhexLlONY2bjR
EA9F5gstuMPLGfbK/11MC9NrmA3fFXvBbjQR+4InnTkB2iym4EkpcZaDfDP6RkGQ
Go80+YV9bTkvb6m+xZWMJoMYG8p5Bqp42UkK2W7OUXcCrqOpK52YP/Nu4bUewnuc
yGs4B5V+TfYdJIF0/rmH+1bF4MC6KG3e/thJLaGs5mB2wikPPxzCIUOwWm8NSWVG
PjkO9xYwktp4pUEGZmY5FsfsD7YdPZkq0cXyq03+ubZgSeUit+6tMQxm0b6+aB7E
8YPmZGriPQB+ZlqJLLLqyXW9XfWupOPiZcDsjD3q99o98sbgqTcXxcVaO5HBn7Uy
uS9IOn6PR2vMb0X7BomKUEgiWro7x77P/w2sVCcz2Tx0WECGfOA/RoHn85JjdduX
WCfFmLq0cU9cK/zfwXhE+sxiDd4dJAlmviQcERA+qlVrvbdTaQU0Ia5uRck60fos
vq3NQlABh517R28ZbvzgvJemeoDSuP642KifgNjBJhfvI0XN26RNh3SOxI/xzaSW
qzR04DLh6/kp+W0Dukfl254mTLPzCBzcWHtDHeOij6pOj/x9e/J+sdT/IxbB9ri5
4gvPuq8kvJRRxK4q8zLoOL6RIlg4Zg1fZGaXOpd0yucEeuVpNM6GrxoZM5PiqoUz
6GlMRPzKH5xwHqX/84OzaeThftkGHeEDv7e85TnVoZPQub4t3EbAlplprx0igXfb
QF8mfK5MuHIGAbDQqnob7FYI3EHLjXJFh2cYVnjgZvKjUm7Z/B49CXjjCcp+g2YV
AHF92SAqCn4zASHYo9FMj2sqZRkqeW/AEQA/rXLmKUq5ACMlNsk08fgbArvj3jcL
u3BV5Lu9q7w5LJqEU3b5KlgkcWRUJfqidm37i/OjSogVHwRTMfloEzPYT3i0PINO
Y9rxUHi8iJkVxi9DczBlOXtkrxvB+dlQtkl8Tzx0hX/krtc1cxd27GbEg+ldbzYi
9dwJ9RK8aF2Mi0JdFezMKn/h2FvVPKfQO4n/5DpNd582M0lP9MBefThXRd0+WSUL
2ZCcl7kz90TJAVGJlXOnB6Atr+/LWnu1qwUT94XlkpfOvolQIaQCB2Haxh3RNyZZ
zuBhQxWaV0GHpO+FVGJhVZgj0GTshZ/BJdd3p95D78TjGLFsPeKUxLf+E+JG/szm
oUDwDHmKr4jINCb6PnGc8RXGWPH8goYQZTO581V1mN39q0C97hgPtaWj2oeegJYL
2wW71lclLKRaUhYZ5hlGiq8CnXL27BvxSPCd0WYA5u3ZlyfM3Zbn03V2q3xauVoP
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nUe28m7dmCPE8nMbGiZYNsgEs85MdHTKCrOrVKg8+NCzBiHuHfIATyvDnO7RxgbI
rP2bZ3zpBL4Afl1yGUoEUJzM5SfNUlKOM/U7vdmcNFkiklaKhN8GP0YmvXcSsQmg
OwJMVQr73nLFOlc9xov2tePdVnFqeKhJLPBxMT8QBB15Nsb2V7G2ayR9RyuZQg0C
czd3nkIaBiR5BDXoWWVj17om8d8ua9/n4hj662F52erIDWuZ+T4udOWJsDAiwkPu
fCiN4JQDmh6JUmHTtHFApWNneI5SwzhcTnshl1m1QpQnCce00B0+rNhmDvo7XPIU
A40wJIUagZVmHG/2W5PwaA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8720 )
`pragma protect data_block
Ceo+qjDoGq6/N3O+wVv3OubzBw3a94Eyp4AtQXURu6c4NuECqcxKPm+B4eHwoyIF
cKrPj5Zq107/3HU9xWIBx/ntKzNzShzJ+WLQOMyuezcJLriiYHmEovNf/o2hl+BU
yb4xQnOuRcR3VCRzJf+44ZsDXS870Dv4JcY1hj7M1+iQqgRkMmoftTEvXI+ma3s+
/rpOVfpZPJtsDB7KejqoRrjs7gIl28/voYmCja1RfCGzkidgesLeIQzlBGPuB+bI
eaNdaY1sEXcpaiKjogNaax3QJQ9XcIgzENBe4FpU+ARdlmjXcGQW61AUCVK36pGB
PAg6jFdQeSHdrqcMzwWtPsGtBzdxs+3Tb8QLm42YFYED51WSN9IKDoBOmVcc1MH1
Wwcwtz/mWgiOuwOLH/ylN/UPiqt6/Nm1UuuglApI+/IBcmXHgJLCwa6fCZYtSjlA
IC6al2ZKY/vkr/Wl5fZN6IBO62L3V6X/Q8FTdINyx2I3/J/+bm0EvoLBmP42gRZZ
EOPUhX8RdDGo36VHagVU2xp+oEmjDlwoo9s5JSWvbqnigmf4VdD9r9ptAK0RHxD3
X0hDzGiANAd1RKk2Ph41U7OxBUyi1qVv8r3yDmHfoKXPO2vb6gJ0szSvZDfVtecL
aTjUROdN3oN0Z/wH38r0HMRPa3MZY/wDpawBLx5pFPtdlHUTPaUNVmu329cR6FEC
QZvi7M4OsHk1VDv3/76os/7vDlwuuOaLWH/gdKdzIL1yWMPBlJ25Z2+BOGCdIJO1
gCGgkEX2csQu5MmkBu0U7XNK8RnNRTdvSfh2Aw7NbV2l4Uuzmx1x7CqxoN5VDg+L
GCUcAFLDBpGJLezqNuWIBrRUIhbdpTY6bbycK/KrFE8wYB6y8Kq2IidHcAjw4MEt
Nm7bjhnPlTSDQ7os2rPHEFUnpqCaa2TtecEzHhDNqKYMn9mq72d7TIzoHPPPbAYd
KpZ2LhGPyJTJfVqUsWqH34tSXNuC84m40dpnpUgRDSs0rxYIaARZIOotj4zlBkOS
DhXVxcpX6MAOLJnU3ypwZRd5ptlfv9mRzxKkzmCuM/mjr3zS3ACbUylfwlZF6RDl
/OivvvDlYpXVPXAmoFFALYt8/RtPX6Z3SUWhOKuJKXZ1SsQjNB0w+wAt2u7FIj89
PrQGh2pspi8fQTIEANJ0qXd3CtvoYoXza+BLDvCksqX2AnoM6OJxMlXj/ncTt+pL
hpyYGDYs6O0Fk5zWBOc+1gRyD3zkEb9pCbl8Lyl+xcov0fjUOkknNM/tbpK9OCTv
QET1CALg2i310Mo7nO/Gkhl2CkLEvtUWwCvjFQCVb9KwERsyuMOnz06LQm1nxjNG
52qoXo6XP9Zp9b/1fRg6DGQR9GZssDhCKLdVatepmDt9H3jL2jojAd7yXhkTQHPl
6xxnkdjzYP9Q5Af7/9b6MlAXRRQl6C+6OA0a7LVyTbg8qfnPBNkwAw/negYK2hVG
oJw3Jm9zsxxr26bx2vOJo68WxqH73epRo+b6VOix3E2J2a0F/hMrVwSI1mTne8wl
BiIf3GsTJnLoEFU7jqkmwp7ecKUXUnd6Wjyt5EmVTGd2MaqsQYT2oyUDVmiqW3v4
8yw+0l3Hi29RSj/7V4Dr8XbNoWLh62f78qPIF4dVnb8Upeeqd0nvXKp2J1I9VkvM
6yJeja28b4lxubuq3dNDCbAHP5wcyVfZ1Pj9NhPbNBxSFcyavVuKV06VHpY5i2tF
F6w8AnuVHDUfc/aK50MjqjBu6CdjU7/Wf0ySIPeBt+yKTVScJNj+zQOD2bUI8o8A
3meM5MIrQ8AT+OUGq3MA64uj2nsabRcGbsfbXlW3MYnOxsYl5kDogJzRoYgBRLXb
3537rU1TQRe/RC9LCq4+GhW45XS9U/4ylQSeK3TiL+dyQrZHi+F31PZJwBWlYYWD
rzX/EUWwO8oY0BZKh0C74ZxbMsEtEP0NUnphjxP0uIk3dhwqoAh5sFa4IJcf95YE
hU3GIXuc0W5qLdEDOzVNR2nxlCKbeKEsMKRRA0R91lXpIqdgtI7Ylcj6F2VAs2tj
sWZTc5Vj3LBQAg8p+6Mh0SoorgKcXxD5WIcIHWccQkdWEqWRaJ1AoAgoAhJVRPR/
0q1VWvW007XyCRyRfT6AtPcQoV0z8IlL/1YToQ2SAqEjTWqHo1KaZ9dM5luAADW8
TrcPWHVcxv+BQn7BkK0Be9FujIM+SjsM5IODNQcSqv/cqimHu9vAwcgRdUAREcTm
lGpVzSAT3EJysaq+XL+Ucr5Dg1rMGJRjT2s/J327nvgQQDYsJCMTfQidgnpb7ERM
CiEd1P3u5ANm+Bsa9PuZrO1bOyexozfhIXIT1g6C5nScTim4Imd74Pe+k4cxF3WM
x38HOPR/cq0jPXG8L00B3+vjFAgFyAcKfIAVnjCe4sjAYkiQjAEj71mrAvedrsC1
2C+Oj75EbRxhVbJi0exd7yehVPv+OzxT3OXc4VVK45zH7sSBn59WIuHS7MI462Rs
JjH3Jn+ouT7pFe45nTKfyGrjxMUS7+O6UdhZnUX9KGMjZ09QcJ9qAVrd8MlsMzWQ
M1i66KncGRwUrujASYWQvVMIxOuIYJNH0Ck4Uws+sulqzzzmM1m9YmFMWZpdLC5o
cJgwq1MOymOuZlzfjrSPAgDlAQb2aP0+fuQglE3cOB5+qHCJw54Pm1UBvbe8iuSm
pYYK057Anhf2z4C9I1kpAqWZaQ+qyqiVfDd6YFAAKWwX4cwXSQKDspGP31WGoxTb
zwrAR7KnwMI/J2Ox0zkbu7PhPKCSd4vszHUs2hQ/CkCVt3hZVgKifUqKBquqIwqt
Q3M9DHqqtdwsK5ZvswlYKBcYkJWZYY7QKqkvJeGnOwdyr3N96W3VxMRCiQ9Ljlvm
TQQVM2NtOJRI/9nQOAQZ6lLPTRWbC2c1kv/Pi/a7q3v9LaCpgnsH2spFBM3UnYoN
hdJm/cGGXq5JopJt7gvBs49m33sb2vlr8BC9uU6s0JBeJ+6RitycWYbhDCoeOOFA
24K66GHO82aKClZNQaMgME4ySMOdxoyW8gDOIOSFkCtMTPnZ7lSVhw05lWNN3cyN
mYnxQ/uZ8eg6vEjbREZfIqQWLaTXJ+GhVbUN1az9tOZ7wTaMZWH1khsdCd+dzlNi
0W+2GWJ/XkhKKRWFrz3azD6JIBi2L+FwMb/vxU3a3YwkuSU5xvHDBCjWjZf7Ip7M
ggz9mYjkL3WmCIFOrp91Bw3q11OcWfd/TPEKwTGXLuv4aUfkiZhcZw7XLeUEpDrl
QFv4zVJ0uEgJ4oYTVi8l9dSq67koV741h9IvthhfokWntO89vVgtzs6LwJujFSfw
ViZi71T+PefiLFC19oqrojagA3kz9uxpLxrcEynkcx+hdWPf1AUkqoEQ7Wlr7ksd
VQD6VaKw1BoQrGRDXO8S5ezAWQ26uroXD4VRhY6TB7cGocguXYLpt1m+OcQmDtsa
oq5YwJEMDf0qObuaazrc2nHqrqWF9Ti/ABPY5rTsnWx9BtT2PIhkF+v0L5GH6uca
4rXmGDOb1LffaxtGQf/mADB3TQkzzy/HW4hv/S+5fviy8orf5AE4FgI5Bqvfam+B
HpZ+6YSFZL3aWgyTs7hAbRVgBJerfD5ralUp4+IStqLxXs2wRX2airJM4Gki6euz
6O7ZFRH998toU+oI8jZUe9v5vNYPKx1QcNtxl016sk33drQLW0bQkDCDRHSUgvd4
BJvw9/BX++cvZoIhpGuei3hO9bugmroxFqUL9DQwEM4LzEwztrv47fR4bWPHACiR
ipn9lWssrLljuJRWiL8uub03/sg7XD4UjQDy1L9EbdMBOLyApaSazql7FNbuArQN
eRjCW4Mkh1SD4CiUY3k6rcUW5NNJXBP87uBxKIDWAWhNxf4tkTlo6Iw0KfvsWmiX
YwlwSFIprbT9csuujMCWR4/OusLKssSeJrK2nXnCQWkfqRcN2cRziderGf/MjXnK
MyKKUfACV8/AmHdv1gkHCwXbZEejIK0qeWoepSDXHWb6ZdOzRVk97v1SAckrLamE
SR9SySam0MJ+EaY/tIRa8xJt/KQQ2vHmnNQEJkV9xzpCYXxOHlhsYnGTzGo/4dYM
E4/zqAPKGafutAJk69LDO+jJ8EhflwBnMCJIPTFh/ixXUiLFETgTkxuvbEsZCmaz
5/ZVJG0P9mHNWvXZUmdcvTdvGwhxFNWq6h4lVN49i/9JpoXt6NFzZrp+u2SIAJuU
IycSqucSDSGc1+0OutmSYJ/T458YIeno1Y8gKwrT3efZEFBEHIcE8UMiRbcSgw+s
/3dDddzivccjfBQP1eR/cUHe6fgPD+Fxwr14nacettkedsjO/9+TIlw/yUqTHlmJ
nUx98U7ErnF4D/lv+OVpKyVAp0A++1bUkIcqvmI89Um+JWAg/1D/DaOBD+ujQPI1
cQzYs9dpuKXZdP9YyQNSyqn0NTuIySsr3POC9DkRZuj4MQnFkE+vhQm7xFvIvpLc
j2MqBSRBBfXVmhIu84FV2FyQ3MAWDyrfDbDM/rAh1FvlZ7yLpyEmJ6pFcsVz3Z1X
Urjn71GUvYNY3PK1XJGony48+d4MiPfjRWmmhTnJYMbrBOqzntNpB1XbzBvPYkDS
FaKldolbQRgR1FYtlxfxlZp4RIaGbbuJ6xyr503kBNalahu5je8aiYmBbdl4G3/W
9/fBGyaWjNZhsBHVwSkizKSM5o2nNLtwfz1uXSBC0MUyZngth04T8TcQG76F8oTf
wiFz9irZ0E8kX8wd+t/scMnr0nKPa2OCNwjayAXd5DPo0FTj97PLTNBdDTDvyevi
MR+QfxYWF16qYmVmYUVFQyFMi4/JCrzVAQkOD6XLfKr3bZqK66kWjySga+DT5ZcA
IWLcFBeJ45UtN/iJKa+4E+9PEd8PmYsBYWke1X/pPtqcG1x/wMk+NGOfUz8bsTtL
Id0hmtaheOgDuVXM8Hi5RukPKv86VXxKI/G1BwKL6p8tKyGvJHRsHfa3CL4CeDin
NvWDaiYAPjTquEQ04CAykJHMrJTn8/7c10qxiv/klxVYALtFdHHgzRqVFBf9caqF
HzzHjtafRbclBjH7oTpiJyPMIN5AbNLWGJ7bVTHOOGAW6ROsxXxdmBh7VsH6lhbP
X93m+pvp6jwg0iGcLbXFZ5c+1Xi1MrHpg3IsQXHBs7c3aQSmGWJatZ2eJd4t5deL
OW+zHTatWpdlbbhw0rb7Psb3qoYw/TjgVuzKDHEPIOZg5LQw4kPVUreA4zHUFTi1
czYhZfw+b+FK+l+9VigZwRBHHQ+dlRWjAXkUTZSu8tHgFRNM3hVpc5UiBhLYZdYD
BU0+fh8iyPTOzXOqK/D6D5u1TYuXkKuAqpT8Q1ug2JrfEnvf9vfftxurj1F5h7/O
5Bcsmt3Rny1H/Li728Z6SnU/hS+FRKHbRZ7/uhkBtZKFGJM+0ZgJGXsTwat0TRSI
7IP2410GR5PgzwNUhoG51ZX2ux6cpOnb92nv4aJIlFK6NMCr05jkpgZ0PocTMsCV
unZU2wjkwm7DrgzA8Ujn6LgHbbO5Z1Ex2kdrZZo7mHvLhHlt/hmS+BEdZLfhRKNE
3k+gdFuIe2mpHdtaCKooTkvMBrgEpmLx5Sg+E/Ddf48gEGN/Hjb30yMnVMrO1Qzj
tZwvAUQMdGy9a+MjCY5/iS0HcDUZZsh18eO57ugnhCtyDEzYI4Agi5+sf5tPBtpo
C9RorQXiUHnqA+YE8/KZJigLUlsV6EUhhI4Hpb0mDfZgGAsrAlo08dY4MVfdm2NN
DPSehJSejwQe4rIDWSjoigLm0cTWU2D7pSmGeh4CfQN+joo9cGO/KyefsW9y3Z4q
8SGV5pDFRctBd1SEw37EQM098pIdWEj5nvkc8dicAcLQ/55Vs782GE+njLP5f8Ni
zAChsulVR5qjzWzvGe3EOh4Qm01xAZ/S57t2m43uprDf9iv6F39Nl2A0k28q82vJ
0H4OXq3e/fkrVDnZbFQIdQMctF0VzzDwePYq73XTeAHNN7oGOiT3fJMt/c5Tr8+j
UscgKfXKtsrtDgf3RlWo9HNuXp48nP88pWqHyGt3tpF5IKeIznmGwebO32ZwtjB5
kkrCgDTQLevO9oAv3lAw2hPGjAKpKfhc2Zdh90VufudzvC1GMN4JGgraHh812yIs
zJzFNl+MoP6YkoUjAYqXttMmlqQmee4YhNj8DgsfOaGqjYpG1AIQksj2nPLkuNVe
JjLGJ374DKvawSMV24jTDujNkb0h7kDDM37KBB6GOzcDILo+FhnBCEDLjuPdLurC
oSvDYKONyCB/PRWcxei/NXOOMzNURnSEt0vNJ53HKOTH7Np2Iypg2zNLZlciNHco
C4PhWgB5aCKh7qX1eaKm244TTRF159W8EAjkN5HdaV+NErGJPtqfnTmcx2jQ2Gf4
WBy0W79PTNbUmDZoAuVYzjo28pHVG647O0sRIy3rukHqt7Oc0ixu0eomglf1ln9/
Wp5xiTHob2fKT5JUMqR7IkxPrk6TPDdbA9/GZ8/ejjX+WxB735K9mRx+Ndl1/+xC
AZs/15/aDD7i2uUWQ3MliXyXw+SD1C1DyriwdQaLOnWKPHtjLEUeQGhdppHUtz8h
bl5+muyzrl4likPTm7EOCERxBVG6rz0O0OJAdXt28cvwOCP6zR+gKiipkbO7AnCH
YqTf2nJTlggOkSshIOqzce5aQVSwWzweD4P7Cun+tDub52XGUHZzdl1XJ9FuB2yd
ovK5oCg/Sy2mblZ+HstnQVzb4Vr2OqsbsYMYpXyiZ2ARSc015IrKI+OCKWuBDRd6
MSRF2/4N61MMV4kPT3PXwQFjQXqsPqsI/RMulCqgtCE0ByKnhyMVMR6E4TYpIVKY
b5kOBANHa43lOEHXhJnp3KtCdFr4BFcM1IPVKypt+Z7mon2pkl5iO/gbk6NIRim4
U2FTPbMIlSkJQotO/6CFHX8IVxj3r9qKxVaoFlVajjiNROkcHCTUePd0JwUHNro/
uWVr64B5I1cCq6N72HHs6GaJWizAVIvZilqEmtT4chvW9qiiYi5wpSkb2fczqYZW
om7+pbZM65sH/eW/iIZixfkE89NUl8njfB6WkfNBUDVAIzIHINEUFfQvynAXA1O3
EwI3GK+ZSvJkj2cIxIEnIOr0sqRO+V69NAUqmo5kBupqxdpW5ZgGuQVbz8EisQuQ
YngIMd8K41TS0hk+uS7t1PWkOijdkMYRZndx7HVIemQv+L7k5SN4JNhs8D5NTemz
3w0xVmD15qw3AhtaTHEB0oMUNwQXGsfIzjI7nNbdSDij7LjsixU+1e+eF4MMxssY
MUxXvoJdE5V7dQMAwqrLyrzhHqe/sUsCjNIC0LRBZNDjs77NdR0c7xna3LgJukzi
igy5EADsd1eG54Rryekrze1hpHJi8EOO2+ltktZh0j0Gdp8TDq7DBVIW9pfqBl3s
s4JkkFhhyLeHumHLcn6dOgYINIOeNu4Zb6ZDMW6msydSL2l/4vQ4LlE+0q+Ws/DQ
NI0NMZ020WPv2x5L+gj8wbxiR6bCSVZHMjeiwH5x+IfeEuUrH/tB479mOTEFH9l9
JgZc5Mb16u3uTmVzkhS8rToXOXJwsXNuK8hRwiJXXZl97EvhqR/tTOBbZPtHh4hb
ZAVvLr0UZjfKh97yUX77qQqieavRRuyTDc9gj2ZcA54MQ07fAcuyloGdKtwblPMT
2iVp7yKsMGs8V3zeLgzxlxhMjCtnvvBci9GDRq7n+Yo5CI5dLTVwWMwnOwZ2Hyas
RRwiBqeM0bKsCUXRc+MuRUXadC06Rr5wJjk5/yeDRc0LIq5fjPiyIiGZ96wemamT
mhDUs9qL9DuMcp6hdS82yIjI71QLUyaZ6Slvct2U0edaS8ZreLvEzz1zsamd5S6l
L5cXgiK6ZY5pyeBnsDsMxRBN8XAiZ0f41zNGrUHOIUQ374xuNVB8itdawXp9iLnW
T8xfnqrf0FjoayrYnUrIePEKb4/aWz63xjHTjNURphGM8KocoGchLGNVABc2PBTe
t3lSB2mjm8SdmjclPaoD/syBOtSGeZk+jJnvvJhSxd7KJaxjHK3V2wVCWq8vZ0H9
pSFttRRmK9rtH6uyMv7GnLa7UN1ewfo26oXQSkkf407n2e+kX1VlGCRIDbJpLJ+P
pbbajUw8dtzRFmMU5Ehs/9EoWb1M4QJYaKzoYCqpFDKkiF/ie7MAXCWoFHQVznYH
vPWE0DdeegMH2UKtO4p8TP6suyGsaTZb73v5mZ5ithciUPsGiIdvGZVm6C2GU93u
/VGH0+YlCXBy2oITxo86DmuHp80ma4bNXA9QHsdlBqp4AJOK+QLxhgOH2H3QMDnB
mbgxIDwy0f8DDaf34VVGkO2G+H+3pf6qXIGtuiKyc6F5zOJGJXffbtAe4Z0A2wYG
hYvy/jyTFeysJBM+M2JXwCPfW9+Tsnw/1QRuBWJSbJUQG1hVvYVOsTU4kdyS4bu3
eXT82hMyaprNKUhnMyZtgEK1PaF8nYjCxhCW7CFc2IcdUpw1xLZM680iUcf6ZEKy
xR0U6ra5yN/ldYCp/kCtfM28jcguey9usUpuh4O7o2Lwaem8xjivXIfahieUHzKe
xVgkEwW81JZI+N7+z0b7dKpQ5GHjxuB1IZ8uTY3LABvpDnRR5sRkovuGC+OYBVPY
cUsicvLxktVSxLQGZ+pERFQlBkQYYpHX0Ii3s+H397EUtulGX26D44xXw+1/8OT+
t9ePvcwFqGMZZPE5RBM/vNfAqSbVLcyc9uVYrAj2kksu+pnil3WKdV8jRhVIU9q/
6w1OBHYL9812xW9j4GL2wD6Ay+BsMX/iXJ5g0umXdsCg375YYOOYLGXa0t3McVC4
GIOKSyoEm41YhCBm0Wh2zAcIe60Q1Y4ynZYJu/L3OlLo6hGRhXTcLCckyhfwBzwE
lwSv6JV2AA4zJjKJrJL6PV/BeRLedVyrh8vCpKuEvvw2EUV7Ucgiwt9KxLJwjYUq
Y5NcUOMxtpn2JUglUkPxI1Zgs3MULA/a4Xuldqr1anOkuxBpZxgLPuxF5IqTFTsK
wKAh11O+hggSqlYM8J/sloqi7Yq0lgFj10oVQZbyBJPPZtb4DtvE8XS9BSrZ84BH
4YbN4ZT4sP1p6Lc6zwG9vCLWjxi4LVdgcDeC8QKGt1YwBUZkCi5AvYRLBBbPhF4L
Wath4kfhSGMGOMSJ1zfHtSvCYG5wb/krzfmUGH9qPjohhHKepz1OZRC7YJ9RiEb2
ovP2221e7Jk7HXu42JfGSy5cZc9O2ZECgz15xOqb8H0CncX+Uf2OPERBLiKESqb/
0ceBLVu2OCCF/cMwls96hsFl1MnUStioNM6oaWkNAH1G3S43KAlBIQBRVnivHsYR
x1/UTwj8wz4CI8VOJK1vxLQ/1cIJYAxtXUA9zNMMDmgcFriupDOMUXvviHRK/wa9
cEBIdW4ylHH1b+7dPzygyaB9iTCHLuPGhHR75UBkqQksyLjkkMintOqVn5xIZVEA
Su8Me7b2Yot0gAyXGYXfP5UZtXeQXj2oBo0h1ZyjdPKH8nSSe6ibh6F9vGa25t6i
OPiNjzkp3x3tDr6+wo3IltEJlPIX2KoWIifj1R1hMzAz91fqDZtuok710mnXGzfK
ZYMG6mN625jMoAX0EsoKdGE8NDy90VsGEYEaIdevVAHqhtyLEqgr5BUiyh/FLPKF
m9rFMuqQDMhzC5OyrmXZkXpkNBF2U3fdrwp0XTiU9zp4PCHuWy/YTf/hrCqKym2Y
eXP91p+w2StvAFCQEmc7CwfMLQiOImjsZuDm1UjhBxhaRp6MB1ikOA27uH5oiqCw
ViYibVcWgzxK+zRN919s4TxN4tF+WRIz77i4IzB2fXNH3yJtg874mQzzafZ6a/TC
2s7cnXwT1wzZq8H6dxwGbhTd1//WgvJJjhm4qc0tsZfpwiJ0/15zStSG1kqrGr1o
mj0S9X/l/dNOIkfIRQELJHAUU3J3SAdqKkxS/uWUfka9zgESBRqEwWl9D+xj26nd
nr1Lm1D3922Igj6KSNjs5FA3NY9CAscYJnjPS2jFfHo0OxZGPwwTiR+ucfYWpBPP
W++hWdcXhjSxRgpnFtoqtiUUaUY6VvofT+605zbvUA9+vJVOaEuXGCe6BnuQJ13A
T6zPc9EmJSLASg0wZcm524u4IbQLalyD3dexJGcoJeI8INhMdGl5OgcEIb9pgx1t
dU1uXgA83u+GzlZ1VoA47lh1hiOs/1R0f08YGsNcqUG+tBwge1GKj+MXAyFwNK+y
LVAn9OxpFxe8yU7fTueC5E8Up7O9V0yW+4r4Qbuj6FKrfw4Sq30YUsaVNIvD+W6i
dRIPKEttwmCBoAMk3kuDMz4KaYDv90EVjdQp+TbXDsKrhmeRKpBjmngX56RpATcr
zy0sqzWwZwcuP3O0L6mI19cJE+oibSVVIN08hswElIt5OQ2+y49lSx/iO8QrduEY
HJZNz1WaqVnHimS1jDjG0YwbdDRl88ipNaJhQjPvmlJeiJX1+UlBJoTNlgtI1a7Q
CIm3JlV+NeK+M53aAbUZHjY5n2sN02mB0efI+EmOzQXz3EOhtwhBxKdPwwGdm2dT
ZxPVoYeYQg3ZLDruY399MBZvAC9nXLloMrud38yKoyi92RTuBULJUfDpKq2gloDR
M0pbq6DTmWj7eRHM/t1bgq6EjAyomENqyOsS/TXyf5gowlL5/yk4lDgWKehXizEm
4RHYQSEReW9gz2UvFtOxysuz2dhd/XAxG3A/XzYPnNpXC8OuI6kDbT/NRpLRcyum
/F09FdYDqarm7uTMJ0wSYxeyDZSOTVi+RI7/9Ma80O0itSS2uRSktCWIe4lV04Ic
gk0VecgaFmV0fASrUoGI6Kf5matd9kh6gOkRqWOBxWTwpepNNLISM6pkaGLS2GGN
D7lyNKeZyiZWu4eM38Q6dtpdxKFjdhhS/AZHXbL7SBSLTGspFhPW4SbJQa8j/Uvt
J+5gP8ZrSTMOSQJh6Hy6i1gFtO/x+dWzQWvYU2/Uj/Jf+F3N+CvUNRDdhnszM2Nb
HvAypun8QtHpFGSoaGP6W205YXR5A9FaeZ/q4HVI3eQwRWm6X8h7F9AWL1JOCoyw
dq65aT9VEgbS3kazc1Rv8Tk9WrE78iUPoe7NEsqUyVB+qjFFCYksWp3NjbHF41yS
Hgs3VjXOgBv7+q4InUffiEHsZeikoso4zlYocpqfgeHhP245tGPA+Fy1uU6x+8aJ
HlSG8pA8stDtgpFXPyxsDsihELly2AkpUvd2G6SVi5P9vOwYpuR1FoW2MqwtZtr6
pSOYsY5cntaXpHkGetOht8tIh6J+ADZh2kJQ1hjQ/dNT1DG+hBN/ivK7AgNJssF9
5kp9+ZMOmW08G3oIKX802RHzrAPJWpCly9hJcEwEjf2L7kLtcO036J0S/51whlux
TVYYExcl0qgmU4+zbaZpV9FOGCCJKnGZz/9X+eborL8DWgPkFOtAd5pQxM0RhtNt
SvjIaBxF6WBm/JV/rpZ7fZVmr90TKQMHrxSiIIhFWsgsCAq/6bAMI5+f0QB9if2B
0IVO8zCNE4C6n89a7w4OwYYzr6d5TVNiY2Ol3ABgGMZKKRyWPGu8dteWLE+aRz83
pGUD8sG3X1WZ2ArGEvFti4YYBl0xZVAGZPg4IRbS+cE=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RVKbmy9lQjwgNCo2qzZ7CeWwdKGgiPdu8DS0Xub7h9f9MEz7vfbCPwNqQxMpBLbw
Qgt75g5hdgR/Kx0jSQFuQtmwCbRXW1tKv1liX+X/m5wECNfEXEwC3rvb7VxzAToO
WKtZqhHB37/UqNRAMB7ZdXCj0jgKCXGse+apia7zk/lY7JNC3kr8E7ELgiDSFikz
qWpN5BNjdWRyv86ckKG7/Tq+HU9w/oGWouRwsT8RD3uNo09E2c0bvOvfuURRslBB
LZn34B/+iPGtEfPIW9Id5CJxpjHJX3K0Wb9ZTWqtm+rpV0ysjaoSTKC9i0Butb4I
GqxGq5j6BKAD67XlAUjFAQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8400 )
`pragma protect data_block
/0oL6AoS0sCHKqexxh5E7cNO3BGL3oE42de4XHBml3SC2ihXtlNOxsiqrz9NAMwj
zCHONehdaM1ZDW/U5YQE3UnZ/UmBoL6I5KLiHgSOJQN9qfMAgBr276wSYTaQ6ORW
fJydMm83FMoYtxr9IyAtKEEj9wyyJfpaHYkUsUEVVrFMbARkoFJmX8JvwFYuQxaU
q5F4fTERwMkPOdYwxQ72w9WFzZ8IhXAUUHEOtcWMuyZ0tGhKB17/NWaAP/aa4g/6
5KN3goHdB8HGF5Td7Wz9Asw5dOTAFbpE260wlh6TskD1V1Axevx7SteY34vhxbhq
9Q9N69a3dkt3aRg2xiR9icrcnNukdrExxPouwbiGsK5fS+crgQesgWJrWVoNwX+O
i3pcCgpkjGUVDNJmq/tU/uwRh0CK26605jvRAu+lUUGURIV/pQVUCGoGGugkplYg
hygZ71nq3NLL3S5CR51DCqhbkwQlMU2ncnrctdHx1xcZVMniJaaeKtLkGMXcle3V
qUXMpwy4CeulFY+UVrdlHxQxyLN7q69ViFUBqw+Pbbinp8MrVBlRk5GVUMeFwjhP
1w3tFYSAlkaZnGGmoXEyb7RTn0g+OYD6i9gTdxZAu2KIuwDW0bvdRSyyMVNJMIEQ
nHf5u9NFvODZXAfyMLCJvzAateRIj+Xcr/Q3b8922I4JttUPpl/tuBA2FsrREWOe
AO8eMjEQkWYotc3jRQX9CZlMJKLkv1WIOAI003hQCcfjOAQRU+ZkvU/KBpi1ZSKj
BV5FCteA6b6uj7RDnnlI6e+hfYzGg4Bv648UbHWUNzwaKWL8rbIBdhudvCpauyAY
2p3U0/WDWI+AHbN8ejrO0PdmHFicghMEJFzCCnmrdp8nFWW1qXucE3MZNpgnTr2s
hworeCspc3rgoMPlMMLMXxeq+m3dpu0t4+r2sHiGD5JeF8HULJ72XTENAeT8cf82
qH9peFbK7C5eMEktTE5RPu8tatNWGXEWu8phHWXUUyEwSAeOiB11vMgzgwWBON9S
jmk/XEM7DSRFID9zYboTdmVs06M87nH5SQ8FcmeyfvoFVraty7Htket9/aTK/j22
WeRrysBd8jp5is3T5CngtICc7X6QPM8JCD+POFEsBUwpGSOnQ4niK8tc5MBGT14w
RbBORs7Vm+8M9r57Vpnf1OFLDNjOtCv41S2gC798v7IZ6HQm4dFX5UkDlGFX78pH
oJoldT3G3JkWZ1IQHMhnSFX8fpZm5skCL76L1wL8nC81ZnLIa3Rl/m+7HO9w9Uo2
TGMf+LNSaiK3Kf1pNQ+p7WuRecJJ4RNvkfaZEo2JZ+AHljt/uB4x8ZonGSec08l0
zMwmdurAzyy1jqwvh76XVV/eR9OmjRApRS3Kz6ooouMV33ueXjIA9D30lDDfQS7X
X58mrzJgsrr3kyKjw3+vlPcQC2Sr5t2ldfFA/373uhEQmOHEnmeJ/vta7PUwYpCA
Q4CDLgkPzNS7vfr7NHz+GA2JMxDi57REybVLuo/5vyXnLMSSbjHaBAFgPYB+7oEh
xoxZ04bmqfzpaCf41qXmp4HfJKA+mvcVv3UGMLKGgmUoz/4Yd+l8HV52Ykepn5PO
2zBCndUTRpMic1P07ZTettnfBlFeCrug2yDycFvBWrPyDE+zRhAnV2iTdv2S//Jn
UC3bSjIWp0vtoTHLaxs2ZMh+4T934NEuMl4CNmdUPutPwhLvhawqjR2NEX9bJXWV
7pXZBJa/5MGMNHEMg2kUu1C/0wMMpR0c4CefOFEX3IMPVOHBs/396aQAiun/JhoL
Zoe00iWpubUuRcAg1grdvZKZnF+AkD2RfoPrgLWw0aYMrrteAWSCsQ9SSd6KPlVl
CuTRK/fNok2uP0lo+VSB3D3FSNvOl9w3rRMFg3EkpKuHj43V78CiWaPHZG97KDnZ
aUrQVzGVW5YoQyhqNt7eQoyKUWcKsmzzW6klcpHNBE4eUu6cscC1yzuXw3KDxR0F
z2sL3Mqr3vNwoK9rxoe0j+nlrxuvgRF8q2WMsbQs0Yj1bgQ9Gx4hKucVhOMU/G6g
6kDjmqk0Pk5EFUegm1AsWiJNSqhypXImcdIJAFoZB68dJL7uk1vQG9Wwg+qgqYbV
wpjU9OYV66N6NlC0QaOGb+VFrQFgdUw+v6WsTSIzhElyUJ+seoohxQ8fyAhYLyqq
hMkN9/Bw8qOwXZQT8PgHA6yhTId8DyV2TTQ5m/LSqcDxGy3DMCJlvNxu0tDgJdXd
MWaMqtCiFt5PdDLFkSWDBe9eTThqgyDxzvbJVdcCOcb6oBbKmkWxLoIqsHWrVziG
nCad6beVV+fXws8LdGNy3CnmXoWcRqfNRd/zd4gwfrlcdoXANC57q56WgEYIX13X
Tklszc6jvdmQ2HekaSB4cYmUP3fnISp/k0AHdmgT4GOhZMELb2IEqL8AMZuYqZXr
3M0NmLKix6q7j338+UOThz+6SIdWOebMLdUOgyR3jWXvWm9VghYzJyXu0CmdbjzA
bhNczeOTCvcORjlJkP3l2V3D5XKBjG0t+oZ4AljYDj9ZGi1aY3GrdaJZDfP2H3g8
mmbbAVcJqU3DQiDb6QfTs+PFMweAhJgLhv/pZ9GAEMSDT8AazfOHbowFrCVsPgjF
BeTd4MSLygHUM04zS0/t1gIShReAVlRuqmDyXh3KB9wbqtWLqj+BEjkBMqZvJGzz
ndy9xrCGaW9V526K0b7H6DrV+dNEWFcw3owz1cJDaYKRsXFYoSxZdfcj0RUZKcuI
sQQG5W7GOqfPN1d7W9WuZ3BF6xO7MiixJsaznn1cNyJw39+H4z+zf5KUfQBRIDli
oZKfCC6raj8TxsZpgn5q4GP5woYkWI4aPppPDfGItvBigUrhIfQe1LQWKDEw2GFf
zrukCTOqNGk2AgyGLGGpd9BiqpTIJHKrfT3gyxYOF8/sJ0/eIfvqyTpTMyAGDtss
jWPIe8CG8HvPO0TC8cRbQFzcP9E2/S2yHcAopLyzhu9IDRgaQCfqVMNl1/b8ZMOR
u8dORvGsl/deJml4U0mREqqxP3Mmz0EOgCWqhskhgyYF3gxgtF5m3GVNvYHpFYAo
yaTxt17df+0sq3WBcs6IHAcFJY1U9MUiETmM8IQrJYJ8SInzskmw/Wud7dI8H8td
rklsQDIhvNbF610TwWoxlFIc6iVWaOSFvCAi4F3B0tG73STQbRuOYOK8rqMczqST
A7DQg9DfXPommhkse0sdmzuZiMYtP7ldGKpOrpxQwt30kOEBe0jFM99cIDLHDAQa
/QO7mxrsDEXU57mZU5IeKei7lNwktUEKSnOxWlN5MiKip7tinF9BYUJ2r8YS9Lis
KXPEnF20XlsNtJEv0V7YmQLsTxjhlMt1hvzGa8TWcRSkWs0guDZTm1jNx3UW8oH9
tKxMyDfWdOi3G/FYjikTGiGJ/bIFrGunHrqnwu4GgVdjwXb5n86yaisVOZQW7rRL
OpN3mQR0kZj7+WdObxYCbMffWaJSFOUlgX4S5ZIKKrQC+KgMxx6p8g2j+iKPFSje
dLdJMmLhkThalsNhz3k+YET5SZCE70lQ/31m9TQoJuzLPqn1954Nvesyia9yRR4t
n6FMXY7jR8F04o3j7S2ybgo18zB3jdlpMcf+YYADw3z+yRw+Ih6k8ty6N4Y25aaY
/LCSaMemAOoKT5cQeYwM9j1Ab2i1paybtvLnOkxLSXck0bXLTwJ+9dAHdrCQLeCR
P2q8VxjwJU8CB/6FTxSQfb0SYSMnH/ujlegdDwksDJ7qSjv4vNIf4Jn+yMRTOQO3
sW9X7yym07yUfTqYUihJ7rsY5pDasYA5jY7Z4/rAEk50a4l/P1AICoHmrDna9guF
nGMW8U/q7tTnnlzeJka6KKS912L7vf/hU3MFFAjemcJO6etbQ3WmXiX599sFC9yK
hz5y5DIICDvl3uj1iLIKWHJ0n/JjD5AK+s9dKosGberRQJlBuKqwWDXMbxtWSMzR
BAXnDrkQJRBChBhUPDo/a0V6UJ9P14Rz4vn0e0i0U6OrFvGQahMx5yCY1TMv6+fu
CRkykfA6EKfBfNw92Rn+09i/RdrUUANDTsAQf7t8eRTsNwvAzWGjVfeuER+EHI2F
onGT6KE6QBFCbUNa5yePu3t1LFb4RVIxnT7rffNNRCd617NU/myXiVtgivDJVk4s
fRGgwWcND16ow/M/q2CLGS39wnDIHQnWRivcflkBreMPddMjzFyVP5W45KtyuP4R
OUV+Nod1EWgKG1TDOcdVoHt2184VoTZjsC3q/gldkpNMa4xxm+w3EEA8C9x4CrbO
zbfK5Ah2/B9W13zDh1deYEpg6WYDYNj0hqEUrmqcyTcBSH2sb1JMgAm2PcpR2IUh
L0RLONYYxaxx9qm3pEOXiJ0rUAR0YZN3H43ME+Z1e4/pRyoCuExiiPgbvCIWRGVB
ImO4FnihWfHIVPsd6IVREJjkwAuEdkCuqyJZwUVyPCefoUmnvQSXg9qrEaj0X2u/
xYUCZ7Jp64+c4hUHQfenHChvWOQr6Elqho290th3q/xxtXdiwPK/Fg7uoHJWs/79
pv6sSsP3D42Zz45xH7Aop59QmEEI6yJ9fbED7OWf+Z08An7KXcb3CEL3gz5klEgI
XfWNMEXT+2/zuyV0qeWDkJs6oh0pTXuKw1wPFFRM/KmXy3folycnEzMkCBrBOtRh
FwsyZa8M0u2RnWlqphhjJLPpdUhGCoZ3VYRriDR4YFG9Ai2DWeNINzn5Qm1d4XQe
13cqVaXoZB0+T3GzBAtlz9hg90pQE9zXqJk3EULaPq1kasRi8yBPvfCYeEImgn90
beMXeZ0iKVhc2wKNhSktqt9mMnjDzI8UobFfm701nWXQUY9ngpVv05iJP92+t5/+
FJUv+wr+H6YiGsooPuSF4xLfL11XVVdM6YtjOpYPwEUEv0qxoETzj9z7dcW6qQEu
eOMMVymoAy5pjXJyflrowN4rGsQerITjALSx08xYlj2YmOJQ4RE1KCnPtmDPbZBx
esh+lA9AxciZNxctR2NpR7nq0rh8DVhJiIguRH0DjjnOGZVP0q+6AelbNWHO2V2l
/yPhb7BNJ/YXX0Ni+Uzl9STLs86Qpuy52TRPH83rDseF8el/Ez1yjQ40Tesoma8k
TMJFZSyYHoBYtYM0g5RD8LvPRZRt+TCJ+4EZkbl2awypta2/Lfl92i+vJ7lcpSIO
GfqzzdGgkGg4uKzVkzoeXsfRdMSWKKXSMi8tbg7c4MKzYaeFzGqcPPYLAkMMA84R
5Q/+Cprcs2ivdsGuskkt7Por7fg8+VGQMu2MiLVVsrtcymPwvbAQWIMNA5aSrS5/
XaS1LsxOLySHHhNrZv9eY8+EJ+VipZgNuyywpL6uTtf27YbXmZnzXAGvYsgFohvI
84+9G1i/n8ZFhsl9LREVM4cCngBgHpOWc6D75lo7PmodZJnOQgmPqZQkhaVj+ivp
32Y1v5kHFAKu26SjBQhkPwzobsnvfPVpKCqEPnkYW3jUdHL5cGRl2zmCNCdRxsfw
4F6LRMM9baGN7l8hE8EmRSLNoY40SLeVSeQFqhA48YTUpr5b27fc8N37pTwK162O
WhQIWZfyOGqvfN0K80sjt3ZhFAo0SxhZObh1lEpql9gi9iatUo6z4aQ/nMNwRzoG
sGbvMWAfci2/GdPdzfUbwnJJ4J/sLdKYJTmXOO0lFvbMLXFquv5epAeDDdShKc+5
RerFoMh1RBM09nauoxc36R5iq1oRi+TXcZwbnaqMUuwLlNZcc2bsFnETnYuuJBU2
/CwvA5lmNlxrg+lcT8vf3agd/OrUtUz4STxSpwgNYpyqlCXuYRbmbVoX5epFILdU
kwovSyzpMilhFym3Mlj/1jxdaJG3M5VVIPiW6EHHIqGfIt+0VJYV/c5HMqGa2qul
bajttQh/pwYLgF+QKrof0S24IK4KvE6mIjnMAQxlXCY36bJBa893BPhwKBE7oNuQ
VBTlZGLhmkkh3xPlG+QRcO3/DiHjH9Ufq7MHJ4GVOLzwzaUKntcwsV+6WbC3W5wC
OWlPJ0KajzZolUGBKxvPhIenwidOarR4Vd9bdElISiUUUhuYu7FZYY1gvn4owFI8
MmW4thOiLea66EtvuRlDRKErU1tN/Iy7s/tu8yNCZZ8vURwdnUXthsgWp6bfE3bX
hZwQThHgNKdUy0AI6eYslKS9hiErldOJsbjp/T0VrA76DW7N5heEW3XV83NmgskX
Zk/c16R8Xx3jCjwllF6+LsgaeAqW30J1kt+oHG22+9K4yDdgnrix2rg3ABbWM8jY
hsT6ne4QfZ0/j0Ts06dIdWhUcKcVn5A2HI1dLXC4Olp+e5Y2THeXKmmyiXXyXDdO
oFdp0wuzITvHrxA6pNMizW8I5voviWWIiQ6J4/TeL1jtjMm0OEvm9w0PudFzGyC6
2Pc12Wvgs2Awoo/FSC1AKum7gSpPYtzYBWfO6Ui3s6SigOIYkaI8az8N0CB/53QI
1Iu/9zbR4eCeUJDiaEm9k1if9gECWRVrw+qHolQH5Mn7YM8H6aJuTtvOhiR1sXpz
xTq3O/DxwFLV8g4kItDAgyyoxPBp1/aIH5OVC8EfkoCL6KP9Vs1JItYcoS3G3U1d
l0B660XOmDt0nWEOI0SHr2O2wwi6lBNV7wgCrcVDY58YIgKLVn4U/8w4sJwFXlFU
KwaQ50WDsiLmeLco4Ouv2maHrM4wu7k5/FBvT7uxAu9j4PUaslw1pH20/4Xi36Mi
3jDew4z1T3WSTCHcfbvs/C55cSojioQSZaqu9jQTXk1TPC8RQ/CzCNgLmgoD3JGC
ojLP+qVujNSa0Z9I34jb+1kOhDClXjwp5vRJ5fKkRCuwzxs7Ie4vCe/89URBYH7C
QJX53udCYzUTPsB5oCZesoLgvQu30Rn0NB5Vm5NJwIMVCjqyTsYPpJBd7XBF96ur
qwVggK/4nNk83YREJ2PGh8x891cOrtZSxt2VuMYXrXELzP+QJZQ9XAzzN8O48Jhz
1q3zU1YgXPC+Z5SIh192UhtmbubzkPQB1pIAx91YXO5Qy3jFOcCY6E4NTAmtrZIj
hedRC5twfoSgI9jPdDcQZqYfb+K086dXgm4uczSs0qsRUtFmWdypYKeBJmIt1Ekz
EwgUrGyxDTUCtoCuTYHSZI0vw7L0iUDet7P5mbkWHV7azHOBz5JY4FGXccoHheK5
gC8M7DUn8tXzs0PX0M/6QpOMV9535TjasA1uNbU6+rDBcMj/VgFWrxC46EWWhvKJ
URWt1wFbkm0/WNXMDHa6u+s2f4Y3Vx9Jd0WFOcV2ZLhIV6RBGhdkTUv+sVfiD8bk
wjgL/uOHaH/S5DEq/u4f+n3uUVKWSLXUo+ao9UXsJjWOK78CKBSXcf0+tzIQSAal
YzeaYR4IXectUjf4vaUA2ETtW/DeZgge/y7+bd7Y1qD0hZ1JERE6NlH5NNoNTPyx
6J9/W8KWTNIE+V2ke2MZxe3smGbFLGEi9wCq4AhwYhzYZRdkKESPJuqxyTDdvsDr
+m51NfW2+DkeVCuGntxXTLJRBthCnVI/fH8+/IqVJi4Rq6LpLkWBThAcFyptC6iQ
0OEUEIjAkcDDhmRPQ10PJiGcakoAAi5G/dDXQRjfruRePUMdJ8fbGuw8rUNR1Fxh
2LslXFpuYa4It6+8kB1vTj231va6fwQnQbrdA7MHF2KyNcuN3nmIQo7NrChaqvsQ
rWM63tRF6eQWv5t7aNKfIKcVA3fb0nrNsWbaWLuw1UWQqE6SMijiWvcPP8/cPg+m
nkt71VozbLk9F8LUxEgpwrkhoDb6i4PymW7Acr1xYpoTPIqQo7xlJtdgw27VKJl0
j9wJmRmckyrm+fle4vy4bqfvoP3nu0r05cAvGbnR3B1VMy4ZOvGBgjXOAZdkAE7t
JpLghTGjG5dHGhEL8+17IC7vu1nEy3RsRFGB0tvS82e6suh3Ut8cjoIqrh2kGm1d
0mePHRHDVxRH74QQar79W5FjFhKotAk4qixomXsffTTntvUqQMsSh6cwcbtMw1zN
64IFG2VjdaYkHW6Sg8E+Du7WDfJWtQVa8wSEFO0roc9EFBITzMWi3cB5TtZYnZLg
9di9hGiFrJW1Al8/t28y/1LT6jqqpQmRUfFuN0y9uU5RGIAIXFn+QynIImLIzRCz
v+ATHFgqsxXKoiJuBrcF/J4SnEYFrmXF1mILJFJcBTr0LUMWpwEAx6zmkO1NYX7q
/HX9c26VbbJg5fDfwS5jlc1Q4o6M7kTnAdD1V5Gj1ZD1Fa/6Py85sHksCNEbo0Im
X/TH+17ysB1hiU6XJJvUCmkvLWuws7X4WeiFGkVIzRjE4x7lk44SwpP0zEV0E+aX
Ozz/nMbEk4RLwi+oiFMEZv2LBkJJLUaHULwAtZL/JJxkbs9XyFzSNdeUQsBu08tA
PSWEy5LqqGr3fzG7A9yOA+b0WbE1L7o2V6srdevFa0LOZLZkHDVlJ2qkSByDirCH
M2h7yuK9k/3wuhS9ooEewYmfteZUZaGYIzsUIrgfYX4aIdXuBYuX/SF0Qnjf7FEg
dILFza/CRrhe0sWTMD+CkPNdZRPKBAFhHG0QIUIVIPF3Ogs5xE+lYnG4y6xZEi/D
HRnUaA1ETj7BeDdPMYMHNtFBqqG8zhhysH7tY53brbpSs6UnD/9yYBwZFMXr9dMc
jw49nuei3+tb15leiVD5lm+VHD8hzytgv8XtYJcAb8bcdS6UzWEgnbre6bUxB+l/
Z2PmBRDcqbuSRyfFTZlprOp0vwINpbTUMhTqHotkXV1f57bmscgsjwZZs+YlIGMX
gwCXugnlXd8Jx6AWvX5L4k6YVx3Ue6ZRoMAa0gczmsq7artFcfPaiKFMqoTvPUop
s71GwDFQgQ3Fk9skKUHtSfdDWMCTOkxAw/+iApSquVtk5WefCZfTMPRvukB6ILHs
Q2qVIraF90UeWGxBTq7/qN/JAkWbN2HZE0/4fw1p/l4VHI29gDNamOdIwd20+P9G
Pe7I7Zx0gRd0ICds5LGt9q/YNbv3i6FoLCSiI8lQGI6BhZYDyS9T8Ow3T77e83rf
53kXpjdb1enfKjzX2yglVqTMMtjAwdshY4pEiBCeaVjowpw4lIOrT/iwsRISqTpj
wfRUpR1EbW98qAIF0rCM0vNLAiEeABVvvPTgzqLETXs8wSXwiz1LuwzxBLtFomPo
q0YkZmASO2Sq84avNwTZ9d6LMqXHZ3yBuQuaWGh2ZsezgIcs+BKcY5bdB+yZmL1q
9E6schDGU7yTqtvzFFyihLyu2dzVcEHzRGy8C3V6u4KpINuI6bP2Ixb3dDpAuYVa
Q50jI7HyDfTOs2Ent+ny4bcCFjcU3NMhwuB++N9ur7RzrYifPYcD2f83qthYaCaS
jd/nAtaUCKMfq5yedqdKHdkKRExkhCuNQkP6T8w4/vwNR1FwENuJDuJ+KuTg4fEg
2cquHoNoG+I46RGENSp2XJkrPikt0ysmcm06a9Sbo3lhsHhNwCbGDpK0KZqWNKU/
+mROzVRWtKj3C3yHQk+eItap5hZzeS4YaTI6CSAmDF5dQ+n/hxM7T7cozEhbrdGI
75Z+CpkYTQ0uxLZMMi0raghpkR4iCjQHPUUK9e8mWkTdRMU68133r4imbdyDhTJH
sE1uf5DswIUfkqqAW8TBSWpvAC7J5Ssq0tWNrHOlwtbGPP3UlZFinn3ECOQiC08U
rZO5f/pPSduuOi6ABHfMnbEUIf3UFbztdV8/7JAWWN4EzPDL0ZhGI8gFx41Adk3Q
lWyNkqlpUYjh/+btBN8c3+67cb3oMvZiQUV7y0KE4JY/9yty4Mftptjc1Na/YuwZ
9OiapRXKBWNVTxqdtBaZHCXjg0k9pSrnP4GlE2Z8CNElylDxj3BHacGxFQmzvMhH
OK7TmM5eztmT9jHO+kwr/MBz9BBIujIvOi03EtW7mc3m15BAX0Cy99Xns5l8u64r
RpoNcjHpvmvFdiNjRXqhWDsQUsFGmB1D5vac+Wrex6wK4EkHVZ0LMAouUXC3p6pQ
l7jm82Od7/j7FoMvpeoCDwn5v01T7EQe4nNAtfxyPbq6Ao4f0wJLlx8I/LmQg7n3
LskFRgK6gyyS19XCTJfBvvzljJWiT4jS4//GZyzc5me60bNaYxHgXX0Lg2VWa2Fy
dXhn+Ie7VbB4edqaUhQmI6uoX48HTbnyvk3tu1xCV00ZsGEIu8tC5515pEClEoew
Rv5pbnfYH7c4OiC8vw3OgD2aN3JjKL6iD2GMvxF/+Z9wOYfhASU8bVz88gzWGLzZ
7YdR2zJoWZBZL7vPfiLy075ZUBILf5C+/1nGhXdNcZ+XjFQZqWnhtJcYae/sOw3Z
k/AvEUBnnDyQs/xZM4GxQhSZKMn+FC8nC3KXjgiadwOJULPGBM25n+DZXk+AnGC/
q7NAqUJvAw+Vmqw7ofz1AQ/L+zUt1OaspnSHcxb6FNvka6hwasJEh0e7+QeTsQtM
0yzavEM1XagZpopaJNKT6yTHKb7P0StMTd3cgMKaK6c/ep1VXJ75cYGbcL+yyLQ3
OF44/gn4PPRYZ8rrDx6Azf1/ATHdemVqf8goyfi65llBqxrK8rVbisVupx4QTZzX
HCKqb61x+cgDjORqupWFzcjULwSLy8i6+2gIUMiIFEFYewwn7Z0VosqZfjrRPuob
CkHSTwcVlIVn+9ARg+WclEHni350RF5eG53AQ9osnlr+bRNi/mKxduE1+T/arZuG
ZTWaxuY0dmVP5F8gQX2kBOmnkttK9BIv2k0TAk+5pTP4wWNzGJlGGtp6F18bSick
MCpLpO50OQ9rwKu1eLnd/di87Frrl7IeODT6tD381Ggb6ijAk1kydOk8bTsE2aKP
Q6PN3HHqbU0V1gIaqCtZwDLjpsOMsOB3vWC/yta+u+TDgof6cxB6c5VGHJwiWbVl
qYpqT9kYUp8dLp1B+b0abqpjVjteQvOZQfAaym6o36JCKnoDnjH1mwv47EOPt8GN
c9++tgk42hSOSeckgxQ6KohQEDjEm3qQQM+mfSPMwDiJRi0sDUs0eJnS6UoqxDm0
TVcLBu4JZ6vWZj43gaTNaF1vVn4FpfR5e1lEBtAB0EY+RuESGGYEugHf3jgH2p7S
PSdrA4M0/TnZjHFadnkOCQxdhSuGP322H1Lv1XtgQopGNE1//xjM7wjyVac+wbGe
5PAk1t0uRFhnZQvA0w+IHpG7ztQduKoD/2UbHuy+4wQiThqOp0ihRXNzBMe0DCeE
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FFnBMG/jqDOPRcnGCu1Z8MYdf/sgJ8ccghZJpUmr2k7agxpwSgFyohuPpnSA0g33
hwWM/gLR3wHMOaFIl1z9YAwptFEPOTaP8OH4vNntxrL+FaAtyEtTAyZh5c3A2OaD
+yzf0p1CHw2s7IBANu1CBTv5GqnYPDLWQK7sUhX+ZNJvws9R685ZstuTQelck6D8
36m7Raqn5yDDWf1JsEN8Y8MBDiLNE6DK/g6F5FO9rX4tpbrJdCGJO5jKABABSPAg
qgOVRHMrU0klUHikbxMacLPALtFKw5T9oAiavhKwxyamrXbieofrZLuYsd/pZkgh
g4aFfBmSbllB48Kli8QnNw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9280 )
`pragma protect data_block
tV722P/yz2LrcPGlL4y1Z2d0h0nXD44Uo6WRNqLzhfF8MWay+6MSf/T0hRFV7Qyk
N3yWbgAFQSfB+DEtUCsm8dEGHnKL6Z8RqupFJlxW2cv7xy4DAq/NOHAEAEHIreA6
uUAVtS800uV5ja49r+Jqw7vaVMbCx2IBMTMVYQkpAi0haDf+2mNcAEeY/DW8wLpr
hJ5LijdanjN3+zU+X1IukjWXMDNMXHjJMYz4Hv60u3EVaol5mOsZRy/0H8PNgZx4
wkBpdJrfwcd+ftfaAIqNwjghX7TUkxV9KFd0mWiIvuaU/VfpM4WbmkCD0lXO/Yi6
MvVkXTA2d2fLxYaXC9ZFXUeKPJU7I3QL1j4pYwlsHb8ngYrtMRHYqVrHC20bb9PR
6KbDxGgKgXDXaWJGHDTvkb6rtDcjwVlNBPrDGNCTNS3mqzl0VQx8QfuXrSpVyOq9
WFganCxMCOInR0pJE6QX4zFohawd32zwlc8B7ASNWyev57v1/HQf5X94hDiNp2h9
746lVHand33mzUoOIFslCmH0ERD2/aGNE3E6uLMa4Om1qz1zsq+IYZUSDP3H1cUH
4+KROiME2U/9/l2TyTwePo6oVSPhPW0heKn342fttIKAgGtCFDX1Ic7CCKa4vI4x
XybjoBeJfnYA2DTz/8DYzI9mirXoNXoIv21G0f0cbpMY3Qk+FFi7U4sfw57NPHbX
b1CWuu6H3ZBRgGmX+9H5nDKoGCJRoFzqr7uX82xgj4gYeQFUx4fZ71eP2wuZDxap
yFFXPoYyNgwWFpNLAgXmsQmZsm0aR4or9QX62DE6qT7pws15MOdl+jSOqMoqCEFq
KlGWRqD1uL0rcaWiD4DwDc4ei9eX8dcQxoByyvQzwxpJ7M9pyB64qf4iECs03uP0
VGqA4KGbqoxmgYoWFzVN7kxz50ZFxV26BCIc5b0iyy5J/vN1ZmfQzkW4DWVFCGW1
8nRyM/ClVRVfTSXJaDOQctY+1tNwgLIT/2zs6Ymb20xF6nQddT2e4GQg9r35RJL4
Wo92xfqm+GvFpJsBV7YLU9fe48CSkqiPND2bUQPB68clAwu2bfZxfVNsXtu/IDvV
v4aVcEuZcEUucreXYsUMmWrXyikJuAn9piOPi4ZODQf9lz6tgeh4wvzHpMwC6qXt
ijgF/sJLQ9kWdnqnN/uhBO2HaJEjARXN570Bcd1ExK0huNvWS7I8kWeRRe/5KYlH
XJT8lqJbquFV6HiKtX769tyfZe8WmgHDxlIxIQuYxRJtNYUBM5Wf7nXbnMSTufwI
Er4d5INa+WyP9ADvoJvpaB1VpmMdhJnkn/eJIvojoaVDNMYMatdMsEI9F/C6oS4o
qqZTFbyitv0bL1Fu8VSVVdORaEUzS0LpvTQZLqb/DyvnaSIFMIM9u3BRTWHnxEym
A4iHHH/3kplRu6ggE20V+sPy0VkBMgac6Q0YM3hOJtWM6wyPoQ0+Mj6+MCIPV2Wj
61qdU6wbA5aKKVSJYMmIcLVO7IWzWMj1KBy8q5DBzBshyy3xu5Wr0wsJJ0cO96/e
jVHVHQY3rupSTnm1iHHy341fnZuNSoPpAQldGNGTpo/UB4jhtWQGPf3X9rVzoIVb
U+4SAeZCbTIDcjLAPeHzyUxZwFhRQKYzxpfLkP0Shwz41C0ICDNMjwbrBctvg0Sy
U0/2Hr5cIiHIrX6yd96eT5EVFSjiVZv7dsh4lA3A8C4LQxcisWgaTL6wCv7mD/GA
0wTapWwAV6BsJo0VlkSINNGRD0RthMDBKAJUYvyOtzkLOgVk+aFiZjR8j8H0Mw0X
j+ndm9eGB+6EkHwLDVBIF6WajTLDbsVpK1vdiiDF7/SBZvkkJUDrp2eRp0AhIn2B
A3DAdGZc3Qktrr4PgY1SkKS5ig7+Z8BJ1DyERVKcY99mY3Q0ISE22H4MRMUi64yW
YLzIoEB9T6WLIafEzXxCCm4XhkRy996ka5FJ0O1EyyWdn7cLqJsBQHPrlsyr7q+z
gnFRfX959B2909VcysgpuJpty9gq5RjeTZqn7S2xCd0vwMH/JKuY2el66Hz5f8wp
Js8YIx04xvavbVguDM1ykqce8dIHVLpkn0ovXgaHqmtf160J4LJX5/oWcaSG42WC
gdD5wNA1CL04ivrhMiB4irtoD254Vm5GHu0sgyI4uh+TX9Wh2UHxKCq6co62iWQn
r9j73SLemWaqgoleH+y6SZudq2t+IHylei3lB3IgichrjAC41AhnFsTK2ixpUb8L
Zd5PI6Wz6vheWvrFW+Iqu2mQ0duspg2nh4mym5RTylsmGj6PYu1KQHZVLOeW7KBQ
ZhIPesslGyGJp9Jdmvrj9ori3pgxPJpdl8DeA+RaA4CnQAgSIaJerpGKuDT9HOjX
QD1VMCT9ZR7vaFaJ7Beqhu0AqbiRmgNrlZjRxHuGh63eApBw5wpnE+QP9tMaFkT9
hFD3d/TAKhESxI4Ry59W/afwHUL9NtYUFnnyrcx168f50U4YEepOGPEW0sKRTAlK
E1fEk/c92rhJrk1926gkvc3KRl5wAiFTbK9QgvwW/nJM/NJ1LZeXKcOCxh1O4bhC
NR9pkj+Uj1B3Rx0mGewr9CPpkFHwsg2WXOCdlyfNfBPwuEFstVg8nsj6WrDUbmgw
0GU41QodYoW4ytkYxJ7z1JN6ZN20V63kVO7kMeBCHn3MASnrb9giaM0CXPlRzoFl
x1qxeNb4oAafpGunDrRLVHMv7CwPfRcFlxERwcKLfEyDvULVGR6GxLyMNojIvy1F
Uct3Iwz7SP9ZLYKeuW+8zOpUDVEZb6QjiVWbY2uwOCtPuJfxNRhcCCMkWM/EfaAh
q6we99EPq20jlYWwCMnWA4gJHS4PwEVtlF1mQXB6NYLJ4HAvCc+XX4O0RU/FvgUU
5j8oZwr5dmvkZMLcc1YPTOpLluDNpCFYvM9J/jt4ArWyT9EECZYhDQcp/e9U/T74
keSyqR3SLGAGCb3AWvqoz4vZMRcEqDQVJrrDELnmLGsNBEibHjI8EYLR2Iom+6K0
XxcoMIrYbkCwdZeJsxRSkRGN5j5WkZ8i+g2whJYWw4TUseuiGt01LUZjDiAhyoDU
JMJT2A6axipJLq2uRJRRTiFyFTPNMcTqDDLDEJblYWhep2E4tIxyAenpKlDE+9s0
+8ZRa4JO9AYqJctywRu093S+2wa72tzfabYMaWEckKDpdDVmjw4qUSpIIxcXz8df
7vcyxPHMbL8NZkV3FjqWdy/f7vxYjwp3XpeBWIG0OMzXCyoFAFee+tD98jXwo4uS
t90hIS+/B0Hs9ybc4kEPn/VKnw29oBXWARXB328zlgJGL98Ilh8dqtgJuY9DPlUw
uTNzY8kfHLBH1pkUrA5hxiWbLC23a/iHbvk8nwvu1eAX9498b4+lh29s697PyovP
w9OvLGruZ1p5eiPMUCNcVPyyeQ4jnameKMXA/EicLLimSoS146aijxNJ+7k7ouOl
bUamiEQArEJUhMd3XCY5q5vmoYTxImPv2fy0HgdD5R6Z+XN0zhdy+09F6X2FffzH
47NfZ2hj3FuzlIAS94BwNH/KQ07taiBxdJ6RpDpYF6PTJDdAgAGxZj8gWukMWPRn
x2mwNYW7ACHNANrQ6H+GejxLNDEZXHiN/CNjqk/ozM4rdOJAX6xMz0R5SJTdY+W5
uMdVKF4tC889PV407U7XZJ4c5+bIQbQGNa5IgUVhj12w9zkosdSvksiedIkfwYlH
krCTwWeHWCLqLBS5uG0BFXo/RMmwYr+bgBk903m/JVUsdEhhZVQYIpJVMNxp90OR
PiYF/KI15VA4LgIp4BmW8ZpX2OJXXF3EZSXbzhQAVXf1kpT+Xh3XxyiZdTpcaHOe
BRkYOghxs8gdViq6+Mop9dajw7QSVwpveCgQxqx4BajYmOcYBcB0nh7K4xyTvOB5
T3iMLi4UL+j6CRKT0XDRSYiwfkUrkC7eQMhvsbbeSFTUH689tm04Mkx391d4vxjj
3l/WwPxwMprVyueQ7xvJhU1JMhDj+5vc1aFKpcnoNssQbQYiFvQv8WqzVIBrwZiH
bJHviwJypqNsuhXtB1aqyCT/stZ5BMij1shKSsg31usThdjMsLXgR/0fguCnhCm3
jMuitopmShdq1yLYqufoJV8cSMCCS8dnFOslGXCcxYSW1BrzKVI0ai9VqciW505b
svf30WoKrvUe+sPFseYwUBguCS8zFBiKSon6SOjit4pCvnP/zxCgvRAt0wF7e/ZL
xAn7fnuIQMgAo0fUlEqa0f3o/zOfQ9bgQpTNoeG8AgC9QfR4SK0AevO6mL8ALlV2
jYUaELy2MTUtJhkR883NIr97a4uV+SUP8r9vxuueYBWALNBxdeBt4Zd5X7PDsEij
mhSrXdui93OQ9gvTd0h+WWzjhhFkE+S7Wy/h6euPYAMvxKo8eK7WswX1bZXkhVKV
UWSEmTDgbA5VDOE5vKNuuE0cN9NS7FiMdyZ2JPA4RWqLlzuBkvqexh9xWjGXez3u
4LpBW46gv9amwzPJqE8s+5UfURnMyWud80htzLs/28W7hRFCM1iqyLXOeXFalWs8
JZCftAPIeudptSEZiuN0+qH9L2khKOuEkkVUyKbquWYQgHmi+atKjnMKJJcYxECc
sJU3lmo9F5f3YabmRlNvZN4pgDLqOFQnhswvrckuoDgdnstZ8+38fFw3agAQgKUL
5d7ncOpeCZjs2Bq5lbucpRHS2k9OA10E0KaGAMDZ4bCY/ZfXK+QjkoDuotjU9Qh/
+UZYmawlYAvajxpuA75aUOm8Qea6PHkxR+ejuo7KI41VM4kdPkve9wdD7BqxLqsp
mKzADiBrQObyK6rxTehUL9MrNwlyamBpqVZ9DdU4xsvoCQOUp2eKyip2G/7mPGdF
XHOeIfpIAIv/xlVeQRSGKp8PrwF4iWbSP/uTbNrADIoNLhK+sM/IHIr7iJbupNrG
CXjcDr2U63EpwiiM7U2baPK/eH2e0Ej2P9tkQdAwSTSUoz5+oPoD2BS8ARfdYURH
+XvUm6HNYfQmKhoGzgqGaBzLz64BlsoNxon8oeEfUZhUZs7WOA8mbeXN6ykpiHUt
ttFXpaclygxZqmuFFGggbAzh8CITRUcdvGbzkFA5r99SCksLakSYq4Hu4GQrz3s9
JVJfO7i38XoTtIy5QzHhZkWCd9SqkCGZIu7zOtfqnNeVCIIXmM4Wzt7ZkWkSgI50
p+K9JUAlIr4c0FtyeJezE0do3zjs/8z+7NjIjcZ+0xaIVPKl6I5W+EWHeuXdFupi
k4uUsevkwdJGDih0cNGOdsp+1rpQ8nnli0ApA3tJIq3Lm+YryoSjrv2xfQNaH+b1
fzmGDlRi+ysOF+Usiidfq1ldHtr6jCtXCAEY227tBlSCKygEKp3XYJILQY2sljAc
W58mQ2SG2FbxbhOwxURFc6zBsICHjHnm2kSvSB8z1HDFIOLRZkJclnjv3zVyQe80
fCkZyrhP8m7WEzxrSTZRrWaYfgg4wgLBzF90ApT0inMOCLhKFYcqIYGsbx+EcUGQ
emcp6WYf81LOtcO3hsrcSbBQY+r19rPeK54Cq3/vwbcs+KVQT4a5DiLGKXLdpLPP
kYLt9wmrSsphFf2de+42RuwHT8IrQaa9Bpoidl0t9jVpGBeuyA+u+KV7qWK5fd5B
VJOBPKnAATIoyiws5/zV89s6lkrClivgNxesYHodlu0tmS705vllgOP0jXhAu4kg
0kXqfckNqwqFqH1KdfbJ1QEayZZY3GPxxeG7G7Wgl8DcUat/8fc8tKpieXntdPrV
otGssG4TGVUJWtrf7IQy46E0jVFPayPgPM7iOH+AZO/y4yI71dJYJHIiC9jnu2ux
TOXYN7iJCB0dcob82zn1QnAz2VR9DnKS6Rm+5rb6zAi8lwxi2dDqUWIghN6XmbAc
C5TLcVqJp3dlgtUCFWJnMjWTlrzrPkRXrlgrq6khXBvACPznmAqRNdxlv2ojpxMo
TYQll+hSLpAina12TVQBqZEtO5hNCoOlc+IuvzUWsn2xraLdfH7k14HBIF8+EutU
7MJYpd2RHFJZJHRiZwoCAZ7kKUmPgP7T31iHTqBe7F69Q9zbkxX4R1xMKjCT0Lpw
8EoNUAO3fMBgvhp+J4P6oPMiLRK8kTcodDFdOkmQXjdLYm73TALjBUDv6a/ugKs7
ybFjgOQKPzr3AaRAhq9MMf7Ma3x9k/rFohNVvL2OmdPxCrBxclZCRgR/1cYslV3v
0v0oZ+gYtXYoNxwl3twjiiHeuOMU9AbJw7f93FMH0CDQUkc9A3B0ifs52+Mmd0oB
Y+sbGu+cY1ijDqnIBYyv/O3TP1QMmNWv4S4C8pOyhuBDUNc/T8A5jC/AzpJc4b0n
t2/9s7xALUIY4uMJ/ssIZOuKhr5mzr59vpsB8Z1cuIPV2bVW33FkwUniUrEMOehw
lD7knBGFttolzmtp9rae+/pPEcCPQw9rty3A1o3Wo0MHUQwCUBxlcTXnJySl0VmU
jdP381JKNHtXdiax9umntCC2+J24MU2r0a7MpINOo4s5Mv48G7q9CsArF7RgjUvO
4MBr0QpMMlQNBx/JWTumJovXoUR8dMNzb7AIcGrBdMBMYqtUhabkEuvdKQ6xZhV4
4Mp31ttBJJqUyRfW4vayWyc7Yj5ziSpzFdnK5xJvveI/3LvNYERgBLKh/WweRFid
pxm+k9GNhx1UjPTcfRf7dFQFXL+mXWDBxa+i8MexM/ck/AwFo4RzbCIpRR0MmDE7
BXKauZS2cz6XmVj3vqsc3mqyEal+LO670an3MSW7oP1/cDmM66alLKRudS1HU8o+
n0eXrrVFxczDE95uHMnMYJhYFzrowiKSb0V0n89TgbJQUHBiVUaH61bGx+kaGXAI
lh/ESBx2CtAontucmj55YKLgXYdiWITfdNE9d/TSm9FeXoJclVQsn4yMrqdnmk+z
4Ua1JUU9/yNJxO52zdqETxqAi2Di1fZudU471X0v71i0oE0pI9t/vXt8YtSS1bpc
SwJFEx8qt0aKIhECUiytwXmbphlsI4bPTcfqyr2DuJGFBCrYlVp8KB5TSaa93BgC
tChxf0GmgvLwNrEN59DPivPD5CkyYn47bPKEbYkr7jjwdLIQAxKRLbSAb8qmh1oG
5ujRuX6Ma0hspBufG2BNMCXv9apM9EOZsd6AKrVl+8Gaq60nGWInSlAtfifBt+ex
0ViTf+TRKNZQxnLuZPxwpueumnByvuGn6miZTn/R7D1QfeMzk+u5PEvxSv2vUbzw
xoFlIlWmAxvEt/rS8A+FjWaXyWo3Eku01ywwB3skG6bJQb9l+aW+/duBRtdJrNJ+
lESbDcla5wFvGvWmmYdFIKZ3d/aGjeCTyNjNCzh5b+Vb5eRetIB2E7SXxYxYafoc
4vSZorqikBldPwo6B1ATr4dFo7GcpcAR2GopAnYA8yxR3ViTknaOWFkKF30Jo3M5
8xsm6K59vTOXAQ+hz6yzWWkeNtc0cqoZ/741j+bO7k2zYjwj6fOxgcnSQlaDGRyb
ULApttjM0Lvn8Z60CN3mSjTlzOij5i9fgIkdkEA4f8f9hoNrTre4YR/sUbf+gE5n
Kdg0EOfr3/zas0UvdbTzNbU8tqNX/CbQPoqHBIGHj2kjEZ9h/y5c6dlbXedtAt8z
rFgGqdC3ofEuG3O/m8tgOT2pvfbE3eIjaLgsdHbQCgIYOrBNd9htIQBVmDFzHrLr
9ng+rO1JwSdpuMVziPquAk2zQyFK+10JVSvgd3Uq/GOceLwlQ8HuwN+TB15lHWts
H1n/zZ+3oRzDgp6++F37oF692mzjKP5vSVliQDBa05KwJFK5CipG2R+NCzPgCE3m
q4e513r/ae0NjaLkrYuv9Al6BL/fKMjBPzHqd9qIgwk5WPb9Gn/bS/xYrKpLvsug
pB+y/nqSLKG+gduHLwUOq1FUG23JqCYpqxJUXjsHVZCi2Cp6mF0eOb+fUYTKvG7g
cUMIvJMuV156U686RpaxB/woeoDpngysuWPySzuX4gd+/LMIpb8PBA1e065eDluh
jLnQPFR+W6Qrc1Koz8CnDvP2nhxki48a5RjcDlyA587fY7v/pfdOExKekeVw2qT9
LJzlyNHdHtSQT79F4vFO+/QAZ041YQwHcni8Z7ohlhk3QBWb3bd61TNVGWw3i6Ym
eFYi6E+Svj4iM57ao1L899/EzJwrIFdN2py4A2Mw2raaH6j7i7EdtzWUEQHNVC7R
9yqFi3PeCWa2rTdlXA9Q+iQ9wMnmJ5SXDtr+7WPgNfYnKzGPmQgxPujUSDAVSzjP
W/9Xd0FTxj4AfAqALvga0HJ8udk0NrvpNk6zr7wRax9JJiO5C5olr9AVHm1yhAGL
DagkJBxkrw3YYohr2xxYIGSq7JrJVmpEuqtRaosiNVCa1OU+vrls0mLJofGlguys
SZjM9XEhNklcEPBeYmRQE4zm+E5UtPJNDIw1pPmnYqnRtSsePWIdpyeLuu5a/NWQ
0rSoJ2ZnmgTSCcPH2jiRFqLc9h+O4l3eOBWD76st72fKJ1c0cSk8TK4bTY+NlKwZ
nNMHihfWwD04Xl2rEiITBpO2kaGvp7M2nadIlvk6HwCc/MLF+2atr6x6TFyYEgNy
13noanRrZoOdSTaB5/tBsBRjN0dlSpO6N/qyg3Q1mPv6hVrFgmqr6Tw++KJKF4CS
pqmHjzFgairR9fmOOlzQKPDvL6LLaGIshah1Tl4HLGRPW32zxhhcQN763FEKchI1
dtRtgkEgj5QnSSSzbMZRxF6ZNLMMq1miG1kNELHmjPsC1HCyRLfFNoLO6IupYJyy
0B7SuVF+7wddb9m4FroeJdA0GddjeKKgitChI8RsrVfmlqUgO86/Z08c43dhlZnE
DTraYWoHrff0pMxOlRm/iydMHhXAdHN2rTNND7iS8iseHlHjbOO5S/9eQC3ATADW
m+eQaTo4thXZQxhPhgmgF877olbHKk1nWpgdlAcfhyytehNm/AX5Vdw+BWtqZo+j
NJu1Kc9l9JTgRICEPe5+ERraHF6aKNlP4mTGUaT1ND/hh9TDH+5DMI0Nn4FFr1xW
lTUVOiIPhYkelh9c4EbrmCpXy/+6VDdr3lj/Lu1EVxMqr1+o+xvR0JIMNyXceu1F
7fdxsfe7hguf8hXRZRFjX03t6YGqHMqb71lY1tAU9CrnTXemG1T/+p/zUp39A1Mc
HtVNdItEWCQB4zFvE+k77KlLIXQkLr52qAZaK1Oal7Aq9aFNenIDn9A9YdyGO839
DdiwkkUOXWcRjNyoLmrgjwiTGkUzznB0OrJnmEPmF1E6IYXEFW9LxXAIoKatcuir
oz64aILCWoklnGhZLjgCJrAdj2uC00lWPUZZ8Eocfif6nbllYFq1+Dv4bW772Lw/
fb3TAAGUK/f7U+J33NqoSPfbELek0+cAOzmSnAmH4y6/rlijF3f7Ee2AUPhgc9z6
GvBXBFwB03LktZDvZeSER7dxGBqjVtTVSbtgPeyyvojScpVCmDspJoiLGgwIm1Wh
456YLfMbGfyu2igvLkqPuL7hj31UEzzEgs6xRSMgiDaYd0P9ym/K56xwQBbNX42S
QvXvWxwq1JaA8+VTkzAsSsixr1pWfk2GGd153elq+8zYRUM+puISHWifwgNMyW5r
HOVOBsyPv71VlwgOYfye05QR4KQi0PsLsbh0dN55nW/bAAgABwrIFbRrtE5Jh8xr
V29t7aMZewkEF1tCcM4CeQ9FdzJaD99gRh1ZMvdzNyXw5jHRBwyUmYAvKGRjRiZS
gmTcahOnDfEU8kG8YcSteieszCa417xtZnJTeKbt1SBALZgbr4qVr2OYss86dgPg
VE/u6TG0zB8NSag2hw54FSJZNVKtZsqNynsmBL/nrwhk6MuFBJR+4WiMRWPxUC49
0PfgczwqaYG7weCeCXZ8AVsUePsqPrbHDujIoSMPV5NG6app7JvYC29IFlHvIWNX
wccX6xbmirDUfmky0SqKi+OgLmesI766rrphwI58Am65e66v38x1VCBGyhfapFBF
Td4z1WD4IZrGnJsKAdy0ad+GPKxjmh8APDqz753o34s0WMz+twcqx9tmBNWujjdg
uqls0Uc20Zja3O4av3XlkCc/wbL15l6WdlZ1iVMbgK/fJI80T/HI3+VHfMllt3bW
Yjy7o8C+PSJCcpw0DeW7TusXMkGBA8K/yupx72t/bfsqAXfV7WJmkIGWpRK/HdvT
OrLOULE/vlUspLIbR++J4gCJbTvmdSREKRZ5j69x2a34aHUvzosFtyd/XTmTbg/Y
dgaAtKIi0xlrui/OYG39e1fCHFyAP/QpdJz4u068HcgE5v42YMIkCLsONmGiZaod
ciKr+nyCCfEeunaVg5ypaHaJojA9VnOJYRtSn1fM18Agyd2824TN9F1ytaeLxdVL
FOzVOPrbI49v3fsnHO+6WXsBTxM/opqKvFTKnLWv31SmC84ifOzLmil78uEpJuSW
zzQttANsV/3xcTKo4e1YSCA/YPgusShWtAwbiBN2rLvsefCTvRI28KrIlpMsGxBf
4nLpVjU8b4WBanbcE1mN3w3S4lDJX+xTp3n1nhATjJgk69C5z2Xcpq7+6jWj/JE1
fK2XFd8SZ4iT1BLuw5d79C9jiqa/PvKKRjPcSfspr4T4D9eqiQPm3phohWC3b2R+
4c3F7LvDMoR3tDLrZV8rzVwj+6MzfOw3rp8a3BpBCalddfE9aaNdgfmY+y87NYOo
c1FGQLiprxZu0dnbFjUz+gUwG3DM3dSh4HQt9vJTGN31B5aMR7eVvtgWBWTZRhQM
EBpBevmBS/zeQfqrB43OlKWBusoqCNPZvHb6Ev6TUUZv//P7kuBWt9rQyteRnD50
LUTVA+IHmv85w0oCPnDXkFwm6sBs2lnDDtMSnaR/uLm921tcnTxWQzTEXXSkP/I7
0PQCmzM9JrGKU3FaYPjZW5jvexGtFLafTaXYdZjZaMOB4OHf138LO95sCkJcGWXJ
24OtTln9QZw2tnMQhhjKee63OlwP9FtCZBDSLU3Lb7bY6Q7rShklkIlJYiJEvvsq
ZYZx2bbdzR4nJ/Wu6fCCxkOLrKT9SX1MzpDrnc+Bq1Tcb4a9tJbpV5wBpUnVRptU
jh8vrDF3YMVWy0l2MjcGZVWXmdcmZqh0+abt97GFWdJCf6m0HDpAtqxBx7RO/LMu
TrblMj0fYyoKAmE/2PGByidky7Ho/S9oFqd05sIEksPyZ/FIK5hEtuLLT7Hz/VIp
pHhOAmQokq6oPvkTdWDmJqz8h7+RToOaDZVAoqLZeDTIrMxlLTV726YhfylAAHx6
imjOOpSZ7f1/p9B8vjVOH8Oic5sSNNGkv7LAO7m6y+GQhWQGWcx+ehLwh9hghZaQ
C0kYF13n0B1yoJsg+3kJEosVoEF97cLt/00H+o+GzsT17TOkMFMDFaLAZsHn2HlY
EhFciQXad88kfES1m/GGbrVWSDHUoRbd4smlplCgL0BxyWZ4AzxbClHfJZjpDjIl
odILE34svc1/W3O7VHfHUnDaCMCv5si3Ta+0qZJs1uK6xxC7HCuV3bJBFb4Cx18e
NScgHPdBijfGvYHrJK93Wkt4UPb+pUHXZsZIr0ka4uOrA7j6yQnkRMgDMREpLzL2
loBmo7ajwbYY1WZkuLAizx55Yn4UFuqtUOL7AuHzxQBvzSLeR3sQBTNi3tC/w2e1
XrRoKIHzOfmcAYRjX4LK3a+VXDq0gAoMwYfoeCFNmh16mGaGoI1MFrrQGPjuUov1
jZckuIHW7ptm1/1lIuUpeS6GW+egFEdjpdawopSkYPxg10f9G4qxBH/2LACwMrjx
j5mA4crJ8RyW0klgwitIRdobFZr4n8Fcdjc/Beg1pIL2sUlN4PAulEe/+ATrePb3
3U2fKc4LEMSznw/JOIRqoUNUS/GEjUKnMNk5oRfqeF9+mlCkNJwElu/m3gvGprsm
McL2g2xx1I5oSnL+rJ88TsAXsB4+u6DYVVq7AJl+yNchFw3T38niAQZoP3F7ltD2
GY8LSGup6+egoH1tmo0n+1wr16ZQTL4dL2eSjlFmmz+zwpAv5M/X20wIGXRmSp8n
82DIvi5YY2qTIp77ET+/qYI5DCCSAPNIxHo5XPWJtTHQIFXaE7Qg9LxGKwuWcE3j
TuwaZalBV7NWW7DolZar7I3/CZj0R2DfDVqwuBgy5y/pU6HTgLavHUYW+SyzZek+
dba/F/RdnCLlLVI+zDVBjjQrxr+cBLlxaPsPQpIKCwZtutIG0azxhhWXbWILVPOI
RY06i/2nWO2H/KJTWwQXMf6i/RuEH8MeM8ZP62ISvy1GlbArsh8ToHjwu7f1wdG8
idAGRNlKsNuOA4FzlIts+77U9+GTitrQet+eE+qpgQoJpbGYySchMiG+amKO66H2
gx4UUfbzbz1YLGolEJ6G5Q==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cV7hUmXJgpfflYASB5xJw32pIGq7kLbvUDEL0NJunlQAb1GYLoRGNJujfTh748Iw
DcNBVH3eKmUIqbPYNxi+ue6G7+1U5Sy2ks0Tg2MfQk7CG0pQShDAQerbMmd1yzF9
lKyajKudQpoidSEWgDJXdtt3yuSb3FeDd/edOWV7unBMDFFCHrretz2uKWg1iaHi
6IPr+C2kH3HQ5CGD/cMHOID27fjayiJwiTg4DSZtQTe+VXP2CauxVVDOOVOHOsbs
QnidDWeSb2OJfJLMJsfOuDXNUkzBHnDA3nl3PPqsblFbM0cf1eqZ042I9BzCNUej
6WWUvNOAgQmtDU9EMNLJdg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
VfTpskcli0NMsBHOsaUanCVpoLvil3BoMZ3EfebdzrvmfgvnZTzD+97Gkw7BnaW7
phQ0tr5GfRnj+MY1CUeN8CK/LI9weTIunyTvHvwYdR+hpWEuI9Cxke8bS+vbSd+E
/ksQ4pqR2xyvX20n/RCmr6JsRF2S1Vd9hGpzYSDke895PR2p7jdCjtK8a9eDwQjA
KLOKh2TLNqydupn9PJGwlIZ0RHvC4ZSgF0/beSraY1doMISUslAiMKmLw1TUHgN+
k8C3RluITZwEhgVoRvusf0dHqf0LKeSfliHwiC+6Ndj7BSuCRvAOkbYbeVXxhu76
72OhYRP8CAoZlAnnr5RyeHtyTKTgQoOPpHwcNqftfEIV+bJ4Yyh/9/r3F1KjGv96
iKPGBsWqRlTad5QKnbLYdCobSzMobTFOeRcvP9dfYFeitMSkvGH1QjN/6eh1Ashv
b+tJfE9EoU91ukfxXaxqyfQC+JB9Opd1koAHlkCZYylbqfYGuqATrr+QFQWc7eYQ
RODcDE8Ui2D7StHvSlhz8hZ8F1mXXg1+JvDRoh8lQrrVmj2Kv6L/mrjZskJQLkKi
N7m+ox4oJA1jxemc5mm6VFOKNUowlpRJ3H5/UnclHHVur0yFg/Zfw4bxcR8POL6l
ZZ4iTxkElTMK5F07XQXFmeYmXgTjL64qPC0qJ0LqEmdcCNJJ0oqwn4onpiKgp6Ds
GM9wyyy2bzOLlklRU4RYXwnBgsSH7bLwk1KQKHg3xJ6VXQ/aTvaCaMYtJyIJVIcd
6lvKSEJ1SR67U/WOdxUwyMTtzGl5PjlLYIs0UUrQvQxL83og0qqIeSfVFs5C7nsv
dBm5BHaUGxUu1oTZuRp3nuHkW1VyXDkjjQQjGUntJnOWjRRVwt7DIjZKRIPTAwtm
inWmp2e8tKecRQOfqp2SoB+52pCXdfyprROjHS8DG8+gKL81Mu/GJUXe1RlrOlIX
F3GCzQYYTaP7U7VrVVE2bTcsDe+Cv5pqQdor1lY9dMKdZpuXU4hsDbU7y3nBRk6k
m7LAjVjfwa37kp/nXprznz+2T5iKJhwe904axx4fTXVsj5BjkzYyrfjiPPXmJLPW
JlY00n065Ca1uklCgIGRm4nOs9u4f9Kz/BjI51vLbqqlmEipY9jX7o39VRxTG7HK
R2CFjCcz7A37lKjE0UIEI4lG0MwTzicT1xCN2j+kbZVubhuS60aL30P575qrmxK9
h9O+12WI7lKN/VNoz1dRBwPNBj2VuJXfh8svhUouuQCNUwhb+PAj0RoBwNkdnjto
htSxVaClw2IxMK2hVbhdXc1mzv2zoezwK6u2Y8Yq4gwpgchPJ7ydVZe8VjtFh3Rp
K/QrhZQDyYaqE/CJULGEujKpZKCevi4cn7961XKDD6aiWl8zgBbUz3z5GD9K3caT
uIZii86Kq7dqFpQ9k16jGrMHlfJTVvTbRZFQq0MxFOMwHzxSv9hrHmydPpU0xvIj
KxWOeBs7oMWNFjm9FzIupyn01mTvzd02STP6sqznxQihzgt9t0/TgBzaRwyZv3Nu
ncSHoWouFhaOluazI/ozgFY9UNVOOdJFIIxV/B3+JI5AZCUdOcKntpwvQqJVKxGb
f0CbKpPlU5ZGL45Q+DudcLR11f5qhh31SKrqrs4sSgplaTRjuDZDusdcX/TAws8P
iG6EY3il2DKhstBQKYRkav3R+rw39cLvuIN45bWmZK7h4v3gbIshQzCv8j0xiwKN
Y3VME89xkLIlfjiqGejd5wkD3ZOP3ne1/By383vhPks1JA4dvIbv8Tae+7vzmcuk
Q4+YmCDKkgV6JiCHf8tImTV+5GHuRQmhXW6FSIAj81L71MKRacBX5GJHezraqYLy
Z1D6UIg02AC3ZQG+DUBE/bETftwE8x7O8Aaf1Pts+sttcin0F1Gmcjey/xGKvwx2
fSjKR5Niod4PlIDUGZ/kOHsY/o5XeRqCxhYJpDP6AkbaGtxTqjy2eX+krpXyz2I6
mOgALj6DCwFl4G7N0VA3cN342Yci20qKi3S0Amb8u5j7zEIFb02oqcvscqrpPy0e
6ntglnZtvAJK3TUMDG8v2k63cHzyeOrhCPlCL3vivK6Cddio9IDPkIKo7B7YUoAt
JfsPbHJRtiqoTrkJYpHSoconHtgc1umpaYCvLAxmVsWIUQX0ZuCQtfXK35dT1FnP
QerIwsSAoKg5VDNG3fbyzOK8Y7kL0wucP9FOfi1gs2ciwa3AMvgXzbFNcwndOsv2
P1TdId8ut164v9yskoM6m8XbEIlwr86ki8nAWhd2XCdHh1BtDKcc8oJqPNjEN0mU
MCEH1sYA2AATYucYYJZ8TFm7Mnr/0Ynayoc0WtF8VZTRCPbCX0IeFWh7vnxuR7uE
GISLkhr2m5Rq7/97+EFEyySZMuK7qSpyXBX8EUq8yoZXitJC2nkjWRIbYnFAMvQv
tzZ204zNeDaxPmeLi6F9B3FTp8cU2sP6mvS4DVzo1+n1kifXRdXNzLKDSee0YQ9r
ijEevYQaMPBxPAZ5+H31wcQknvbkCJsp+NOz6VKS4UN73FWC4wPk6XI2Mz+r7fce
BcrAOnH/HvRFWWRcY8U/km8OM4Dt/g60qDrSwwKwn4KqP2FDsGYeZCPoppCDlUAh
i1g6yaeVWXDpbhOcloeZzOsB7c70jJVyo/w4TEdXleHQOczGXjvrUd0G8NVy12Xp
xg9Lakj9lcjL91jG8fO5+/He0ayOE0afnCm87hKYXyGY/NKw8vCwNfVx9xeC3/sM
LMkdjRTEpNBllhDz/OdHQrNakFCXDTlKJ2kxExQwNyQ+SBnDiTr5+26CfexQtdxn
E/uLr2s9fiBPlo4qnCvhvXs+qLQ+OAQkEftXobuWw8RqxnkDfjHjLOEBYmEqWA+Y
js80BmdatX8tpF7nmQkXpRzDUUPoVqpbxWbsX52BhxopR0ob+u+rLmDpZGQwCOSN
dV5MUmJ+kidnmE73gz0jBWTuMW9XdjoAz92K+YnCtm2uPJbkuEuNrpTbIVKIswBK
Luwpdaw6eMBWJC37H16M+J99+uj00EEOlLZABuHOPTRShtmTpAheWXzAeRMr52/N
hICaUbuWZWQYRP+1hd0BOpGEgGin1b38F6ZXZ0YeI7mZjn07ND8+Yzjqq2zTZ6Qc
ZZjyvwBs1zo5t3U7TFFQjuV+ovyevO0LhArdEsITl0mOdmRtNeC+6l09Ue2c2vS4
ebNPLDszB91Jn43iIRv0+5uv0MgonQdNEFTZ2Efv5DmlEB9gijabIfZdoS2fyjGy
C7KDSo9kErMzjiNbpkuAtMvFIl6GtrQAb+WxNdnS0mWptx/2JIfNwlH/ZgtoKOOb
Izgx9b5L+7lBs9vpotquMbFPLukHPJ7DbHaT7GNUTkD1zWFFb92e7XnLOdUA7hG2
+9IOYwg2mtVoufmgmatfo2FZf9uQDXuyssJa+b1CptVshp7XCfDUtPrKPen27plq
llEciyViwTl4asUMO/HmdeyiGwU3J7e9dGXsFFVi3Ke617SjgxpOdRGfpFWeqMcd
Laahyz2NNPI/iqnol4ty7FXkFy6m0jsVVwJ6a4k/GLIz40Vs8n1BUnu5zdEmCE06
luBUMJXvcXaHjodcQiGAuiDdSK6GYJdT3GHEP5CuAWR+GWnYLak+p3iZEnxgxQ8S
w0ryiT8+HmvLk+NpZSNhy1zcxbEkZKZI9baJXpgj1sfJBUgd7SP4+GSOpyGW6a+t
v+bocy4j64icUrcF43NYMKSTvzZUtGySOqtdp7MMVchxCfzwCz2Qm1bRDME2CfBO
/Un0XpHx3OIf7mKH+VVmYdHQcrPkLWAZTGc2boy6EJirlBirXrqmA54F7nAs/C4v
iJRrtV25ga1wx2vhPuJTYUlFiZqgFNadLF3fVbTdQGNO6eSbKcRi7qxFRNaRct+H
DDCIElJH7P3VZezTeLn+gHw/h1iOVfSbuL2255rGgNG6eLgT9XtSnRuaLMQRteoC
f649KFeBi4NqfUGuR+twey+yRSRhWcYsffIiVntYGcu8SsWKxP148ZrlfDlEb4YA
2b2lgDzHjbPMMENEhQTWUkwIeJmEMK22w1JoIjAqu9GPYZ5ATgIjF2yRUYyCnlzE
qr4Ee4f2UwaTR36p0aker9WbB7ebzG9y+fh4YawwmVfvSjwVOffoeMYu1tmHv6s8
/ivNfM1wEwajqXEd80xWuo0KBqGJYByf2nG7n/v9dwalk8HwKv15hll2JsOlmEXB
RIHM0WBhnLUVLLB87jTY0uI4dHxgO/nZOMXgwNgmnXsyWO/2Vlpc/QZdxCQjAJk4
YApcBnfpNI3cPFgTN+jsYRo0RONOZr+mGNowq0OGxmeBIJLLsuPQe0diEqmcP6VA
IxVyQhg5lWUOK2S4VzgvyxscdLOJQQRqPQ12cUwOIReDzETVqqAOt3EtEN0mLWtX
pkO80ZfYiAio6g5YHS3jz2Va+woXunPuWsFF2+dq4Yo2WrdTwxutyTdWW6X7ps4l
wW14Ci3pSPUZwiV6hOqg3TJ+4m2P7A63nABzuXoyxTu7f5G7K4hNNaliXsGyTdmq
wzf2izOm0IjOhxmqwk9yW8S2I1AwiyD2/OMg9wfWJ4j4snd19zAgURwnenjN89O3
y9CxEKxIQXxVR27geJB2sd/2ZMe+IWQMH3cs+JeetoVd/Rl5zItveEpGMy6zOgzZ
Z2vPjvkyF7U/HOnk2A5TejYMOl0L5TGBHAMdSLHfriu3fOq2nRNdf8LNAtta1wa3
M+0Ki8GneuWB84AGTsLFptYnq6XC+eWYVFOFdoZjKTMkDxr5ZFZ2aUWLbBDMBKTv
z2fxnm2WxXFw9UDRi9+4jilzGJ06LTSArs105x0n6p7BRCjfZFfzopkNkXApgvhN
4XRPMD6xMRQhlMBZHrj9YApvr3SyvNB/idy5eIkZxtI/la371246Tayz9WxCnsJi
2MPw+9ryOSgfkEWqPKxPUkn++4+6nOxXQ9Yz3cYwm94xzBJ65ECZydkqtjhr/w5R
F5Vzyz4j1UN0so2K8fZ2NATEc7AIkVRgjw4EyhnuQmRgPmSLi7cZ86PFvXKSk8ZT
qCAP+plxdBM8v/EaBeLuKvG3mFNkH0saFl3rLAngwLVWHJKBW3AYuattlz/elz97
OuBno4JEFo6yHzF5BJRqizAutt0zZJ0TL0r3LXAk+ERr+5vmXoCiyU2o7GvwKYpv
7jUHogbg4W9FGTXv9TBvDYHR33BmwkLJYWmQXo0xo+wDDAvmyyDPaIXu19USM31s
Ys+m2HWW2q+aUiIQ5WXvKIn//9ZI9ckvlqQstwcNaf57kmB6EQu3iKeB1F/7/SgA
W6u5m2uTFqyUTQbWMkCLKYp5HcdKaHsElxPPJNZVZ0/ktfIBLK71uOHT9WgvEa3q
JscUEG6st7kwyyGfK+4AhEb23KGTu5ObIjRpbQZKvXCxz+yOjxBv+l27bouFDZWQ
Yl91WcNIzikNAIarWNi+MnlQ6lMr8QsnmLpPCVZckpjrlC/HbWD9xpEtYHviMI/t
d7oA9K7JbTwRVHj23PRi8F1i6EJ2Jz9b5RATcWJow/vCAsGxG8ghEKXL4OhP3Y6g
lLPg+dfTEMlSnUlcazkc6uKDveCAX3D2o0e+pnt+ZiNvGon0Ls8fY9T8WzU5azWg
i9QJAey4ojvlteDskERjM3CSxIVntHq+9dlXA5++8CQznUKWiE4qybWCwnIErnIU
VqJfuE4OOLM0u2cJvdt2+s3ctOg61tITHky47kTpZZt8pZ8IYcdGyJTP+fmaps+Y
/3AbF0dgPaOnv9hxBey2zwrSA5R+LhJxn0RAtKX3uWNfyEupkvJMWpae3rJZzs56
2ov5s0nfdJC71G88U4lI5FvjZ50nR50FlishU1SU0Zgu3lgtcvFgoiatNMi2gyH5
I1yS35mEAewmTqWrCOYtHmSjim49yD18YDurU8RRmKwPDwireeew0Gy5c3yNjLQG
FfYkRrgkmTpWZz+wQbvQWzZUwa39a+jjnulER1E+omE/UgC6O7zZmnpIB8XnGbcg
yvJYrs9XsSkeuwBVM5Bp4ixAp8pg1vLI+JL7Xvz+yz5U68ZUdbXQPsXvyHEbOJmB
lx+tbiFJWQtFyEZSuUrzvyezqgr1haOfThUbaaE25GvgtH1jJhA2PhkGenP0DMF5
BJ6Qq7K1Gzt6OvpWNmuu9mKZ4hJVLSWVd9Eh7VYfkwXPaHm3InxSvH0YrvcNehnE
7pDfyB3qCN6I5tJitB7YQxbTC10nr8lg7IM/Owk8L0I3J+QJlj0U/MLF014O+WFi
3ASmNHc1HbnCDH1pYywincgFumOfTxvP97Aq4o4IRCf6jj93msS1MIuTPiKIdDd8
lA6ZeSKbrkyTQOqDw0m2Dadw2V1GwWbN+itwp2UQ6wlGu1Dgiot0S+7Jx5LuoHhs
ud2p98QDziLfTJ7OUeb9kBvH8t75v5NhWDKQcZKjKZznR6u9w7mdtsZ8kk2wtLZC
Ev5t7xG3uzuZYiiuVEubKazZPc7S6UN0bjO78l75PGgPXg9Z/SXLACbEseDBmsGJ
WpArpA9hUCAnRvDUPfuurvkB1GnTwmNXu6pvfRAoqIVMkj264SfNYorUMnGhEVTB
AurZz3kkSp8iSuPg+ll4brw9kuQ4BcjjWy9E6KhASnmNGRcdqDh+o2SwPYVFQ7AX
PFrNVA+7G9lt65bkZL6Ybfm9sUbCeRxNjzcP+BIbbENa4yH+P1VzuQkFhceHzH4S
WiDFnB/4QdrXo5XfzATOnNjJfxGdOBMfmxAzSyFc6G/RzLYboGBaNpPqS6JAg/jH
e65rz4RN1JmBgmUTGCE0cbtLeSHcgCkOwzBOVxoHvmkluIxN67CPNFpixKAauOW3
c5tAC/iSmlI9oQhbx470xdedfsPnGaje/uYcXAggtQr1NdIxY6Plqa93lYFt9zl9
1IsqVntT8HpOIyzL6H6i+pT5IZcLMBeEb0CyGosZSE60IU09jA5jgKJDML9oUEO9
bOjLuLrBo+Dz/5kRPqEh+QIUJjpS62M98tIH2xXVy9IaDSrnVZsCEEZcgMe0aTUt
8R+kXbInJyjyPUT76dMw2uJZokc8POs5BEVT5xp7K4trTUVPN7lBi7G4cn28kqnj
LBiGMOS3pwQZp05bl4D9enT5J03u1IjghmFLFIKEr/WNHyFYHNrppCO+ogVPlQP5
Op8ty4QWYQDA6+E3pLrINXsLq2BhlP3ZSVIeEElRhNkPQbrNp+P+LcVR2uaj/Cpu
9cHCuYmIAmai9dFCJ0QFEev5nDeyJG8nYNjEFkWZW0Yaqp2pLU28tJnYiPlfa3ku
Ve5/2oAXf/tBklutz+sFzUGZS5aih1ZdFs2H6Ird9hYrtP542RJ2ouminKyCqLNS
T6zV8ptOecYzDFqpar1XtH5gPc/0TSG76fq86heXqH43Lf2X11tzWUUsJV9s0jBe
tGCGTFRPzrpa/wN/u70plx1vejrBJmTay4M6V7Hw5SL4FEZtTNJAjInftFoJYcr9
//VJe5mGQ2nucANKs65qq5Ovg+UAh1H+gMqKkVPY5ozg4+IzHo4Djid3BZTzQxYU
15nhxCiGu11G9JAM3+XVvsSyQ4wSc8ICZyXXf4AEjpkmDc7v5znL9xV4JX/LRGAj
6LrL0ZGgGgF/bT6n52Td9OUqfXbMlBD3Jchp2SC0af0yRpkm9gEiyGwPix+1FHnA
6xrcjmi7b8idVdWlkL3egidWCoJx5HqVGikHbqI0X4DOBqQzuVignfw6GPdsAZCp
rmMrKDbxWi1NhnVWriCyDD8t1giYSfTJ1ePhyMqRmXpqtlpL4rmszUZsXj1MMj82
fG1lZBMZB3isPvPjA9fhzo3TVNkjKpVj4OesrhndXNsoRk/LgIdFt5jgr0GoaheT
b793Iutk4GHtaFzipkMZXCENlyiDLdZl/hgozB2GqrQrpzCt4hS2By7ubGMyFkwK
oCZ7y6akCstUrtK/j8haRWbRaAfNglDrcn2E/5YzufPVNII6QVEceBexcIhqZdNX
QEz18ASRDVPBjtRwylOGyKyqlOujURjEbCsEcph+EAE77R8bSmJ9OeH2ZvkYwo/F
53UVDEaX7uu4hzB6RKtYNrfvLY0e31niiTDppjYLlFc+WCBpBUYkywKbwOOdNh5r
DGwfGxGA5eiZro3FgsshaBvNVu+J2QPQ/y473bchmlqdhT24reVY9efH2SMZw6NE
2kbcaU6itj8kiHaMhNdpLTfx2KR/fGLJyM9r2Id3+A0BmkOE+99q8ZzlpvWFZBJm
CC5cKyXome2BF51OPyjrFO2KLeJzB1S239pDFdGMpbmFtNH/b15iOwDFG7NRtRZU
1pGWszIVJVXPcAzbovyryiwWg10PPDRDTreq79vTlcjUg4Xb25quOuqHEPwQBDaN
lNQgv7btUnfk3+BCmapWr/EootXMsVQf3PXA3k11xd7cuGmBGw2DYPm34ct0apYS
imOwp8dvkdb4r5oNNxJoDnlDCyXU4yA6rgef9SoHzdBQlPJFNaX/IS1a7UEWNKnF
jM8jSsEVTpmrIwcoq8TNxej0oqzGdDWTobCepR8K+xi3Qr+drC8efB8+CP6Jl2ON
PFjSiPsYDikcTMZO9YCbmH4yIOWBnX1gxH9M0ksNtTPnkdvXCg/4b6peVTjL2ta2
+qX2R1bDkyoaBtEPMru1N0dxqzwTi5JjeFY8FKTUbHQB1WeTsWwFZCWlRC8Vw36L
LdwSYnDtDv5pbc9mlZeaOvUtZqWaL0AJQiNAbCe2AK29LBltn4ZYGmdKFOcZ9GZ7
diWLA0z8FK2F6ncYGr/MEWVsDP0rV9tCsDPHtx3YHYXNRmY8ebrFo5juUaaG5qkb
Tk7VORQmBM+MoFYhNbEbiA67qNlZeh1OXkJFB/LwIs5R8lopE83cjCZLKG0F4UZn
t3X3mG1tzEniVQDIL+FgV5O/EdTs5sTqvmfie+tNeDCSMpRCDyMpiSCIPmZKajl3
xfxWz/ICciM2rzwWrweXCKsciTsr08Dr6SWZm6wvDKYTJO/5t5XZYh3U5P/MawJz
p2+Avt7EkbngFgwbeZNnMjPViYEMcejbLsJ5/crLchyI6Gb8jI9684R6zIv0piMb
6tUlsQUZ0udhruevtWjX3W6t+sweR8KTwASsC5MVdhJkpVzSGZQfU6MS5sDCgdYS
KjV3QdPc1wuAD2+Ae+LovxIeXcu6nd3VYlHGl3xHnqGRW7WNNZA+ISd1ks6ehhoj
ojGNyrxLYm/tlxaP7wVN1OlU83JZ22dfvztwrSPNr6bMwy8LkndzccLHAUJSxKtc
ZxQrwtUpIqwc2lhNlZ51uyDRA9HMMVk6fDxYTR/jB5UpWszbGdRhRuCEkiwJ0/GP
YablZlbVhCo8nfY4XhiiK3wxMoHSN2vyVg/E7W2ov6O/FgL6MCsEwQSQOWHDIggS
6CWrlCTnvTB2S0tSdFzXo1mUa+9Oh4tg0+B5rRxEVgYH0oRMAsVpMQMizUTkm6yi
oRha/ihWX1+DTmRfst6qJbnJN7M/g8bH+LwtwCbiNgkmjnRia9nFgEzuD9UIAfE3
9cp8OGNZ2QtdHJhu+TtPc0H0cyFJBFRFQJUn1zrsqP2kvaAPwHUHsYXuJO7TwgYK
zTAYNFPyWtm+BnK/QopDRUOQtSgVfv6j4t/x1r887gzPgDMMOluJNAlUkJ/SGr9n
oASv/B08Udr41XuO8R1lUY2h47HXuxHjG91OgRIZX6ziySFMdkW+Rir4LWxYkS8u
ttisvAEDWKKMxjWyJeaz9UiwEUr7H09ak4h/NIYORCVqqS0WvDrMjaRUAa2WTOtb
SgkUZKgSnMeMOW1tLk6JclUCb97FzJxeJ7jUvwga6TbR4wt+nJfrMgSJ/6giMaTR
S9R5t5tm7lt6AGme9CTFzNnZQS/e1tH/pBpwGudpDFNCa317TyBuYVF+Oz6KXnn7
f2a4Y0+42QNSQBuYNOkWRcutlGHBALhp6h0byAZuUoR+/l5vEtS6+zZKSaozJ2rk
ynd90odMFBxWxx5xswXrfzbrAJVlfriKIRFqZd4nE+zBJuXiwRqtdHReU1Dz5i+L
WYmvXtWCdOFvGi+xYDvhO+FC4HoKAQQrsmWW3u6KnkYUw5zQIQc46PMI2HBySvmg
J+FuFTBja/25tzhzH8+PmtaN2Gil6BZc3o34porx1s8CSuG4QYoR3Yfxv2Y98cqH
rJ5vEb6QOQj/3WPPyWPuuWGGmcEz68FqPqXWilkeOAPFKSocLugkYEpFke/u6PD9
X1Dae6Vqjy+IpaM6RKIjdKWqV4aP45k0HxMIy2T06Y4HtL5KbHgXON3J7zKS56Mx
oeekMcml0dm25Girgx9lfjttsKc9adIZE2gbBu0998j/GJPPoKUbN0TYNBiC7pGz
xNufE+dsL5mKfLMGUyIcHbNnINT5h7+Svr3D2gFFV6tJyp2fvblpjkT++MJMpL1S
mrfy92ZOvNnkpToXedj2fD34Sn9qd7HjExHqYG5bQRF6ggQzVG5KH2Zv+wkVD+b1
UWarJJR9Y7lg771SkLKd9nOl7byvWPvAOCd+WNWQISri/aDyBamAZnTHtIjsZ3sx
tVQ80AyCMI+RoxCWzxEH+munJNWL/NE5rdSJ9zYfSs0c2MOkTUNvx5jRHCpeIYEb
9SvcY+6uvQ9XXt+coRNmwz9GDmI7RDDoBuLIMkMG8TqhyaULy1af12HlGu74F9lp
1PEm4yIpZMJR/AZEsDNpOEM2rDF50PqpdvS3hUo36suu67K967UFNIj7p2FlKvuU
4fAX+jdRwEZ/dk/j7auPn9QOjEyuSA40wvq/7ZTUzbVm4apwxa+LFrpSpgyoOjGo
1zOV5pmVYUP0tsWvHxuNzV8oAOi/UQqE34VcNoPwo0akkHxhHuYkBkOxdrZYkSMj
HME0cmdUxCC5WyRjy0vJ3O69M/wToOz1Je5feb8ZEUOJi+eCk+7ElNFyu9a02x3n
fW9M8iIbAK8i/NP29ohoIUQysErSC483qhLeC4uw6rjNlyJUOvOOE2CDS0dLghFB
FGqGYyH8tVNFIfTxvqpNligNWB8JSliGGqMVAu04wIqJcVi1WZv/6DgW+mwQMmfQ
C6qvzyDSRxHFCiNfn5MPm9LBSc6UVhJqzrA7cWGUYP/Y+EM4SgwipANfgiLx51VD
/pkaPh0V6b8MJDQRXihSNN+CKSapgsFarzMR2FYmospKzqCs6Xumh15ROyP1Ih1X
DQIR0adN69c0Z81YQyq85g==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
PBhNBd2gr85ktAH5WR68s7Ne1uD6LzUGEAK9aWKEE38v5bLRY8kBeGgeKoCIlyEp
bgdZJOCL/3FcjSyWpjJfG8yMGwvUxyP4y8govlm8jlxtMdb1RGfX0LGxOA/Ir4sN
LeaGCtyij47Lg6M+e16h5cW7a6XKeItNCSZcODy/KS8o0R6vmGpEykAH6NICkaxM
i3I2xBDKZX+YO05wIDu/2rDiHuccWwWWPZkHc0xgRss+b84vi8D2Dup5t13shhS4
Bi9MK4X+kz0MLJUqB59Hn+mtkPbfvL+wCtiLLKFsPgXJetK7ii93q7bYTqTM0U9o
PiSdJ8z/jvCwb71otJDpZg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 27200 )
`pragma protect data_block
Hg6BJr2gxC2QAtejgQ/9034ZOR+GML0sbir7qW5hoGHk21cQmzMBao6H+mYkyM++
ndWnJfNZfk/+3LDwNi+3jwe5a2o1CuoL54A0pAWPu4bxEVCt24wUEHXRgKuWwkHw
xJsQDA+zVzh5ZAhtBfqfG288IXCrmL2QLGWeUTcuBXshO85/4nTX42hsiCh1WvZR
pV6ULAIrOV6r5qzVzz466XH0KiIlsf95IpObBdOBipzfObktyyamm4QNc8gEPSM7
1p0pLjVSWKh4wYbD7P9M+OpgkWPtUUdyxIqJTxx6KV3zLiNLQgg4OVv1yToBc2j2
R3e1y15gw/fAG4JdYtM4ghF6XNxiraRgIXKOiGlGTFVIuY8W3caai5DTz1xK97c5
oh7rQjIBneHmnBavptSRHwroE/bOuDkHy9Hzk/9cllsFiz+zkvT55xxtKbDfpg1Q
XO7FF1S8iLDL9qzC79sC9w+Os2T/Cbhf7SO6k4vdCyR1txEXJzoAW3gjvUkyko4r
LiRzwF+5B5KjNiEXJgrglprLQj52uVCBHo5mo3GUqXlnrYBg1+QHUHRfHLhnqKQy
3QcySj55aHf0zph7K6kOaAV1GSgQ9IFWfxIZnxR6tEgAxS3m541YmpMCJLveb4PY
3AQFhK5Ek2Lbgok32511IOlqVFciP7AeNtUS6KLIQVnn7p7sYjjfFuCklOIFUGKF
Cf3GzSQgMPVU7WdLJQt+3k9X8oXAl44rhwG1JCkk50NWfz+Mfd4svfOCo0IDcsVW
swFGWrQhlI6qeFD4KF14/ie2thr/qBNgDeO3AxkUMYS5ilI+SUzth2GIEsR6+ChB
mVg4aIHbcBoaqci9aWjtvp459dBDyKGsIlg755ei2ajjl9KVAyWpzhuLqrOHpUdm
lcKDX4upgGFKVfCEbo0xSse/KT393O9JCALLBtXwrIFUsgONXQRehY/DXT0xAUDB
nzvjb4AJbcgKBoJOS9AdYn4/yf2H2oGyoo04mBm55kb/5J9whBOOVfhPY9Pzqhyu
aCJEagpTWIbSZFty5MZ45E0+4O9A3ykerLwG4A59/dSmekR2BrYG/jEDntNPRDuo
5VvVRUIl8sNnaa3BevFUh77Rnw9ikmATWB6BhBlpV/pgwEGPASJNWro/el/CGBsO
vF0jE70KfawQCcxkeziViL992J6nNiNCIXpPg9M4gwUWtY0vJll0W4VtVVkCC9Iw
04F5E+1fcPcg1buiEd4g3pR2WOIsxsEASDPYIYA2XfsKrgHnTHS8K/eD0yJunGo8
p85XIb/DHjvR9eUznfu5ebdZp/+o0d07+GskZoc8AK7923JmZFIiFq5eE4KRKYli
05gXASYhIMcKNpmwTTGRY8wLKdHAnZ/+WF5EpboOLGu2XXGx002dqYKKpT/Kk5v6
/Ri94ZOkUvZHQyh/7dYMMYkHHQG3vC+q3+7wfQJ4S24jEmJsorW6fwvjWMLJBy4Q
Uwq5G0hWVd+FQOxDBjp2meVZqK0M1ZJPV2zAPFz6M+m6wyFyR8kwTCA+YjT8hnR6
B2AdlC+NokkWHlwuN97Vq4u5VMO8EuePUqumoyF6RQcdtReBPkdp1hqxU83C6yQY
lGJhgE78BK2A9eYNpaZH8XbGUzwcQin5bf3SBHZFprIUKA5OEt5N/3xPypu9jaoX
fgkO2tmVVEY3+sWH+jb/89ueMhY4cozu0U6Vc49G8ZVA1PEZe2ZunCetBqXlMR6z
qESvoWipF/GEc21HzM0ZUpv7l9nNe58meYEfATmNe6VZIogSGBFBcdlQT8Ocg+iQ
J4inssfOHghBNI1qxjZJ+e6g+/KPP5ozuvQwF1PvqxSVQ4IR0bRXgoAzqNnTjTMw
+hcZsobuXPcrNMUf6Ad+dfWlIp1JKbI5mj2YONT6+9MXaiev5zS1oztMsX6UsKpA
EctgEJ2BpTkOjd3ZQz5dNvv510fXRHWT4AIjXUWV+mhoVntSavCx7PspzNBUqZry
CacaKdkuSabEvAmnWOyKggJUPRFlY5irc93p9nX/bckO+HjTP37nTV4eWX+G1wHN
8Oy9+uQUjp4j6Ty1D4vW/RBbNKUfE8Ag5W4xnl1SWejHB7MR6jqlid52+OCLDbGh
BopkUGEZwZXhkT6R74ItUro4LqWpZgMfJqMHPjloU3o2i1Twn9zSOP5JyaP3Gkh7
pIA1OcBbLcEFR5+hoX720LQIDYKEhbCwRbv1FOFDOtXKCTwBXMkck6ilrvHkqQMW
c89Dcb/J4bumMQ3YiWmmTBeQNRoM/dyyNo2D8U/GvLbdYJKRpC1kdyygcJ+rOwuo
aoqVbTttp/T/JwvI1y3SwX33jDLAkrFhaS3X5luqo1v8ljwqdq//UQGo191GQAOz
HhjT2breGloYbg8zYkSHUB5gGLdWwzpbqUAI/rk45T9qZas+K4gvfzo4GBv4ZNMz
F20w44tAU/W+1y0Z43656+utWQyU5cikpaKrwCkYH6GQC1ol3Z211+69LiBsMGsE
Bxgplnrb25otZFda/0aKjeGgwKDPHRDrGq71EhrQp5sUGvK8rq+KQfZT1ZNgAb36
K2WLtiM7DjkBhXI0QAskEvV2W6X9P+KkD8ZF9Ef7UzAcAjKqx5ei1GgVfMoDqner
6Zs8/ZSAeeWTqe377do6LlVnGVonA4195mi5/ZZitoBwCSFZ0HW61Tm+tQmWDLAO
skvN27rbWtipzKgTbDNbx/EgXSxW816FGHgridNkosz6Mfu5685BztbNYKn/nKGw
QCAB2qQy/2AVBFMWJN+pRaEz6iXP1W8trlZGtfbaCakb7tOJIFN7p0axn5wOKuuv
/mvGt8gGP7ugx3m9V6xX61C3IOKcmcMpUTkCVs1KK6ejJia5luBbsPPt8TL9jeEU
8xsDOG8F/HRdxRpX3zdWUI8QoPbJ79fak9Tdwy7BzjhDZ+SjEtlhAa9aeCj54C6h
JxiImHtYFep6fHmafdjmm20VTe3o3Azgb28RzGHLEJXKIzthibXx5FyyaHNgK6YF
jQKuSWqlV/VBrOwp1HtDdAHzzjeIJ2fl6RvQ2Ya1n3OoPCYoH5z5iTan4c6ePHfI
pqG1Mgre5oWIBKT5MESsNm6IbQMPeyKpA1GKTj1rzrQoRL/GtDmbF+wO9lFKElfy
S+3WMNE6VjEDLB2yS3uG4/2bnPkOjRxCzM8Nr818/3w4r3//Aqfu0Wt45mhqiUSU
tMb48WxVWCBV2rkzxV00lPRVYwmNAxGxUGvz+gjTqjQoJzw8rPhLQkIJbXG7IthO
O4GJ8IKMKym+yPZs9gm7w7I6QifOIJN3euOLhj+vD/kvyRgpozpdBo7Vp+PQnBfy
80dPjF+akw89w1jggF05C6PskJywnenbVUSbOw+D7Oxg2ds+Vd83CDfZHfVc3vt1
8EkjcODRwjp2sRsdrHJ2inOmKU/pCUF3tLxDQm0olSu669dHfzU9P6zqcprbSl+m
/wFZGjCOPnjxRPU7Q7eg2gCBcwhJrQtYdJqEjm4SzqkXg4lmWabeV7I0RFoKGeli
eWAxyqmDtOvFnacGdCA2zV9IW9YJodrOJrSih6OQsCdwcxdbm+2uUFoyu4WY49iu
VOppegFqzbevTCpupu2fgVuauTM1FKf2y9mdu1i9nNoZAMk5XKwYCoAPdxaUCGq0
4PmBYVTxxacHNFqnBbyMZ8vu+fhkCsHUMNeFdDf0l5bnGVEb8je0ujVlxixk1kZk
Cg2lwoiOt5+LSLq4/UZ5YOFddYxWZYu4RVJC0Fr8RfN0cSJ+dNRR2juO8EJlvYnN
PklHKJhm/26SGR4DumNx5u56gIGD3SRchah7+sue6sODBL0jQO/hmYUyteSjNAaY
tfbYdlOukuxwU4fo9q39dNXrCgehcpXRAxdfkIrirP5GJj82ylBP1Z8MnbnCI8Ct
/X+bn3PD50hPc/1Lzy6v0WuxWFG7TuriDMDzIY/eqP94bVzy8mSfzc0HKeLMY/e3
fLIK8rAPiRaOyxL+7UwBZPpkU8XavCKehmKVjrd9ECUNNOGdbg/cessZ/BAOVnU4
NnjD4IrW+HGYQRUqxTVnXa87q4+lgqTMZfZO95iUzk9seuc8Vfv/tRs1DqSxe55x
+kkPXvEAYWBjVbh7PohSa/vRs7T7QahnRrmpBl0BoHoN17ZWM9BOanOwlfERLQ39
itz9lRJwbic0KGXcTOswgp+LnjsWR0j01lWbujyxb4lCBlARUvA6Xbn6k6htwrv2
IV+oiv5n8KId09dgGuLjNruQjbCuIY6wWAqtiy7Dpk1LVTXKNpsjlMw7Y27tY1xf
BFT4XWVhyEc3WGXpkZrnZTb3GkiZDKSyaIboTJIT3tJFLlXm+0KuI4boWdwmC4N0
639d/6dxzbp0mCWU/9oz9aUBlcVMBXAgq/w1X3V8eax8BKlkLqzd6kdOOjhglfvk
hfOkZZxJmVHjvHictAOrhP5ozVsxop9Y1NYD286Z20s+dtuO3nNr+syTV3jFjqat
E9SimXx0NZrOZoQKs9Murn+9XTBYuHICpU4Mdj8I1YTE5/R6lm4QpKoSIhO6SGiT
domZmK+CSYNFtUn/8HMj+64dBffxRVOS/Fsw5pEzF7C+v1xDvY11+FxAJ79abXej
tbO6ZvKEEdAagIc5MqwC3UOKJ4UkyRgk1MyP5u+iCKrHRXPvKwbzQQXC3acP2op3
jyX/88+AzSrZ7GUzRp8M4eHy9tpusetU7aisCxxxK6qufvs/cT0Q1lyrWbBIYjyE
GGY53Al8am14nz/yEQQuCezn6apLXGZrbqy4i6MsIrw8NAeREon5wh7m9PMKjPXv
bzMEcWtGA1l/iNdU9wWYQnHhB07woTs4+ZwcyxLe57dmdzjSDCjiRJmOBa9wm1Gc
f2+Sn/hP154aq/jHeo9Q4LFUjiBerU26zDAUgzZSsedvRybKytZqRiKiJ8wzbCzm
wkH59mljrOzjxmzzpwgeoZ8CFSL6UZ1YVZ+of5CNuSPEcBhywMEcISqmwNn8ltNv
qYucXVrd+/MwxaeYdu5K/6EtgGrM1HOVC3Zv3tjqjzL66XafgMaEUkJAFzkofiUS
uL/uZ07QGEcv7PZM7aoD/CL6x6VCeRzipdY8Q8MRSicSp/ZbGcW7BBY6FTpvKzOo
8fqoUO7wYgJcsb4DLGY7SHcsDX1tEFdQUc0TUpqOqFUNWxYtmxTEFI5EPVEv4Fn9
Cuu1q3jWETsWYsSse320VlWUuxKPWOcby9j5A3UYFRZbsPjlzMDUzjanEOWuTqTQ
ZZXeHEAFCrOwCW9GUBNg/xK5qjwR8I6imQTja4GguZZup6sLnZOrO+l3sS0klZ00
j6CIPr8tqT7h3crs17Z/eALJSIEvTO2k964rDl+hwbP1s2wYBDYw/31rA+sF371g
TtgM+qIDuKkkJ24GFgwUMfk8hc/Ehp5uxWXXtf21p/JlQKZq/63phsLvfDdZmz1X
0FxUbHSgfcIWP5VGxXyjG5JT8qbm5XZk2mm4DD6Sn7WBwjNCDh3MmFLMxWElsOwp
ykkC8etuiQ3XUi9bQsdMZ7oEsSuK5hTM6mevg0NBnMb5jJ2HJzAUeqVRu9EbW3eh
eTA986jPB2fa4VfpxTREeSKf1r752P4wGiVO+k4revtZ/3mNxWOS7NPmPOQWvm6r
LzYrH8FRToPydHIE78jEFo0hMDNdDGPnE56ZO2gRvFfaqmtVg+Eu9SM8UPAbn4YO
Z4WI5/HnwTnhx2W3rbRCRpir7wqTWxiEnM8+FG9GEtu42vr9V8Hhl86SzhK8Tfzu
kcbiTtjbaLkBgrOsveAFXluTgxthz3Efg0wVFGDjn3b+Y/0TVt6GIgi0wIJ3HAZe
+zvnGxO/8EcE7R1UnySQFXc7vPQoDgVwTSxCnPR7GBGCJyHWWWUlBpVVo20ohVs8
fLbzloc+Y7vcLd603xp9WQvQfvzWAMFw21OamNK0cx+xdPvJ2FpeNn7JqFhavWsS
7zH9NFJSXr6JDh2nzSo//iftLZ9a4Pz+Dz3Jxh+hiIrzRR8PZd2Inlc4JA7tznM6
JKLoLlk/sbcjY8znqO9wul6o6zu67sEAOH011Bg98C8tpR3+2xQFAYp987ncErFo
6GhjmAzfU6GBD11lWiaQqVxqX/13qffj+gOd44xweHSpatBCZzVqFNlxZLOl2odG
Gi7szRlkVxPNhCA72k/CUfvf9JMskN5RaP2Njvq+5u/MhCl/Sm0LB9O5pER27nx9
uwCygrZeWkXT1tpnLSkzZZBNnRdO10ictkZm2JSJK8vwel2etFcQcz+/1DglV3LK
URq3+Bv3Rmm63cyOCkSmaaiFSKDO6tGsllyaVbgT+HniVWHCl9BFc8bJoETjhEst
TTYuSP3DUaVrj6amVhekDYfw+9y8sOl7YSfv5BzSmr3LQHr++b8ZVc8XfeA1qlOD
b6Mi/yYoDn5JqMhbkLMIZRQbBUCVz14DnDfGN3ADwwqgzL25+ZZx5cVmpm0lZCqq
+Qgym0pqR12Hv5+7XbcLl6VOuPwwQI2RGaiTU41qstSrMJX4uZIH/053R1zrjvUr
2rsop+YGIpQ/QHC4eN18lnUHfERfZ4A/ZU0IhGiY2wiBf3tRrb60pLrdNS3ya7uj
gXsStzmRL3IcaF5q8QVCAUF5RcPKGPCy5TtxnYL34gE675HTZIIDvs5OfNO1Vi0p
Y/NnQP8t4i9/Ui2YwBKFHIQFeBkMasNL5P8LBOUrmXijpZqrpnfrrmXvyRbSCqWP
FwObtAOCglV/DFVtOCSlFEGBXG2o3mXEQUm6FI9qgQWEBBnJWe63PZCBB+oSi6rc
y39rEMO8VAJaM3I9YdGg/NUCdGf4Cvr5zbKyUW+p2rULcWrVmUyK1Y3SzaqRRwgd
rFBlCe7d8n806xq893rmLoTS7fVNE9a16JNgRv/KBbZLj3atkl5O4E8vrua+Tw77
eTFmC9AMWxaRmRbyJ1lxth4YdhGAnitTJZGPEJyqD/p8tb0hbOqENCTkTeDV8355
dIkVUKc3gQyX0Ha7lZSGElrVqZ/Bq0pWH9eHpRLqUlZua5Gdas9Eqp9OUY0SyrRT
N8joP+RInTH1SYg/QGOuW1+aAViOyLUg1rRLJw13WTP8Kl6eUNMFR9/DPU7S5dBh
IdX4w6A6QKjFZuxV7tsRRkERx21cMtwI9bPszGh9v7fzDsfcdheoviesakQOoeRl
Y4a85g00+dNIfqMO6U13YWfG4mhpKtwZfiGHzPoA5Wf4di1Fy92DIL42BkpbizEu
SEJaKhTWKo6rv0ATCCd3ZTGuoCaQK1RNkQghtHFZWAJUfovdXGtWnLwIsIJTFBNb
mLVUiMNkjVHK0/uNQ2jHzXLQ5YXh1XAgeMTHhNiPyKtGdC+497sHr62Jl2Y0iIqm
eu6FFkdpyvEXSrkeHOyrhUmdZ19Aj/+FfjTe8O5bk0De9Er75pjtZZAfixN1RfXH
pv9uLhXghEGpBwhBbPzsC9NBJFOHTRHZz3yyVofQVcbaagcUiC5l9QZTTl60Fo5x
0BnMmwwR+ZcDubAfygUYCVrlX3/uujyCNs3U2LhnTKf9O4/KMoJ3Ks8PyKiLNMfH
GakNHX+iRrBAsyzDa8DHBlXZ/JJhOwXCbOPcPn2ylDXjjDWFN3cK1RTSNDohl6NV
n7DGwi7uzi5s9oBN9U3/dUa1bDlcwjAnKofhKY9j22gJBzORxuecD4Xb85U2aOSo
S5t9cQKDMOQD5RekbohIARy/tbeW+O4Ee8hRQvSBeK+7eQwqSYXCymJbIRR6GY9o
DC/UJfTU0I2fou2k1yuILLtSNoLT3thsOVleXIPrc8plpY4g3KeSuz1xZfqJz2lb
GU9EAl2kjfyafp2akJ7rUDEcxQgRrNZP0/jBFux6xL15jvwz2UJNne+dJc6wBUX6
Pz6Ghp0pNOVq8nzt40vc0gNsWeLMUmFyFVXl8CcSlPHnT3S95tCwSDLri4XRGgoF
VVgd3ulNJoScJHMccmBxBEfymaKXL7brX8louMhSxTBURHwrJ29yBeal5pRqfl/C
+VCg9vWBUScD848ayjRGqts6RDzM+TYnnQ5U/98EQKfJ+Iucbtm0RNWTW3+LnB3R
Y/iYY2vwPfTdNG60CZM3KN5xYuVrIFQuwq2G/tTQWBZh/YsiTiEzxlMNSrITc5vz
/g4+AtgL7PwrfKwRw5fgyiLIw5qH+zvXyEJBuR9+dl9YShkM+L/Xkw+FMeY+9X+h
Y1L+AzfqdTdBTDPluRvDzF0vZe4iLBd0kUUHfzMQuyZTP4H+sarHlBB+QY1hmlmS
mm5R6TFX7M+0ojr7nvOykSQpLigGVlZ8h+TcghRs46kdxWZvd6dL7ThmTdJH1TgY
5JBB6IfppPcyCITDcL4Qx98XmaibDiirRRxkpl9hqSeX0zJg/Mrj5BWBFEwSiFGI
jaHaiLqDOXRUEQEYH277UM9mZZLgfCO2BSu/TYxi7jDNzFQq60eom01BRCgV2YgN
jvi06HIrbatAQbRPgiJZ50D/jqR8w/cd2GVfRbLTTbHtfMp9ma1+xp2EdGXFfoh2
Q3/wuAZkMkWA9nCebL+rs4TTxaLdYWIXABAT4seQTIs7xWY39LsgXQLSgkdun3ji
LWqbJgQ+5EnOFlQm6M7pQ98D+wkvZTh/WRktFV1ixtxT8cilTPvokv885wgkn8Ij
wvGyEdgbbYPSAHofKMus6hp1kGxc8jodgn6Jrhh1CiI8lY6BXvR69D/im4PvZm64
Ug4cdtRVROoBiUBUS8Ygqj8U3CHpgeCZD7UXMe38dtEZXLFO3cJLB4tUHw2/ngM+
nCPFbvagERc8uZE3PKTDMDu9UprFdsF8CYphXVlXDiw2VURWvusmfS/qwrhoUpBZ
dfDGXiy8GUEd/4tuMpE+Yz9tmbBN5A8mlrYaNp6uI5uJwc/w6JUyj3j/IlYGEj3X
GJmmqSnfH0qJ6qOH3lYkjCqJEhv/iJZdqXFQ0zTQANc9Fmk83dayuft2IsNIMYdq
xYjYb9jM6PX8ok2k12dQYQ6lK2U3LCzqXA+FugIw/FuETHqez+cQ6zks+OIdRbwi
cn8GAOP2mhcs93GG626/uT7/q8fmu65AKNoSLSpRMlV04yrpLKJNEW+sm2Ry8Gc+
AO12l5CbJBAd0tVx4TVEa7YKOzs1bc1EvnUZQCaMGJrXbimBe20sRSyqsaJ2dgIF
IuLKeY0u0QeagoDziaW4vCN4gB5OTsr1X5m/T+qjtmr/CT+IejsOIBJBiNzKr4Jz
2+LZ161C1b+GSsFf0XYPCB4MC0er8YbhaxVkZGH/VeVHuccL8qUIcjtruKHVnfzj
bpd61DuIhZ/tU9Ota+BwSHJB5LOUIDN4f5KUJHZiNGBytY04+2sOhH44Km3xPhs3
rYoaLz8qz2vsfqU+z5IYdYEZFSmceAdrJEweS+HJQyVZR7QfkNREkOwUZ1ci0o9n
ASEOkVurKyz5rYR+jrcbp18CI7vwIbM96aSRzeRH5WzI1TqStBhECzdityxwovX1
GS3grYKIjQpRfjIujG2gnQFCXtizTvcg2ddcRwWRczSjStpHlmEfIdUMG3Scfx2O
4dbSfMAHNhLpDskd0jJ6tWAy1gMgNs+H+584hPc76BCo7Ob9swKNjWeqtDJxbR3h
Yl0dyxoXJhH5Jj2m1eRTwLjbso5hQCCllcGybpifY/HdeHvaDBZSzxZu0kGa/buD
mpZ/hpAgYD+jZVAMOvuelChlIq9u6tGY+rwTTSnEQpNYrG2xesbZ6023lmeMbH3x
hP5vqjhqhRlSTtgmIivru2Gkgq0vVUmfUXK0WM++WeZaXRgCPajaJdy/ltPXQs/R
IdUoXQAFjgaSWzDAKr1Znm77e7wk2whLDnf4D9b5HZzo3M4fTUntNxiSfEyWIKYM
eYTzR2CXjGzrpZxYAfYeSfPc+yiIGRCVUVczY7FQkBA5n8ZqP9ydVasak69RUQQG
rJ96lGJA0XNzsx9ra9XQic8EE8L9YjRzqIYL/nu/AmfcA3nGNQ+zsE88eL8+XN8t
M2PY4zehiqJyQ2uTSxslsDofFCd0Ywr5lb0O7T8Js1OPlR31axriWrO8uhfCtYZD
eAbInGpgjc/6cUxLLv2WcrJAkE2nTsm1ve6prV4EPCx7Kbj5ZXln3gMSg2RylZma
zab4Hx4L7ue1rlNzr+vtvjB5QGNtoCF0nw7j+QIfDnVR6e0eNl1MBgbjq7mEvCa7
JSFsgKvn95tfHMnK8C3ULPFUogniTcjL+dBxAhw2p3mkX3vIV9DisP6rxuypEnDX
bV5T3JdAYCna3FqPYcvwzh0ss1EpO/R6pOgLZ0nyrg05CCzooAKUU18YorS6hG15
p9NG+oex3vcQUuSJuX2Wpv4kNIklPbpjFY57Nj6BZb7gtS1aBtKuYOnedClPDOAk
+lKTRUTn0PwMfd7+cGiejg87ZgzNLpX32DkiPWrLwFQJp5exEchhk33tjBtZEzah
Mtfnjdq8abRIzV+zEffjmwaoUcxY1dKUwPqvGiB/b+m8HYTStMXle7XCgRZGbmcm
zSuziwDX6G6WbfkysWG3sJ2r5mhOqNqzBV2s1KW3ggfM0Gvwv+1Gh0M0xVoMNdNu
3nvVJ0zfhmwiMFdw66VnTiJ+dnAOVFDFZuofTGTIoXjI3fNmaH4fTYpy/mv4Cd/U
SmpuImLRQNhWzkVmMiB1l3bLT6rkUYKlIyMYQy5xEIZsIPG2CMzAZHbpqBxdj+en
NXjmhVfAOmAtCPf5HJqD4PMuTgKt80M+S39z5UcjYY9JR0eysJ9Syxp1biplo/in
Itw+rrL9GhA02+PqyZGPbSHDlunpbPsyVB5bOqPP6CQMP36nU2aV4fsRUNDkSx3q
KXN9VlxBT4T+9IzZr3aPzl1HBqAeU3pfpHKF6Xl1MxHAAxPwemlVEXeeA9vqa5pk
SM3hjmcjVMGotEHvWM1vCQsA7iKKj7pEzHOH2CanAKiyoh16+mRq6PplRN5g1+hd
s3JPv5dT1428Qx81lefM4eP8cjcXsE+PpJZLR254+YF7qqqNJ/8F+syBaCzRUP08
3ZqZuJwsg0cVZxD7F2f5g6ygr/k5XpxzWGg1ROU/p8Kl8bJMx8stFockSrNh3M9k
UX+x9QYlFg5FlZTur8zbSC9h7SLoq/VnJzmg0fwkLB6P32vJsT3AvQxEw0nPdEGl
6h/ZprQZv0jZOCoj3dGcgUeeIqm1uM0gd5vsxCV86sWyGRolyOblKag9R+qgcEVJ
y5+7/JIP6PEG7yafOOfqDufTS7C9lsiuA1Ccanc7OoGWNsZgDOCKyu6vc5wO+H/O
vmSygyDbBT2QXlmk0xch2spvBNqjarD6Kjkdx9FhTNvxObjGqwosfAKVpKdIqhL5
/bWtZ5Rc4dg/0hOwQ7GOxq7j/Rn2v6C3T7WiLol3nuIfL6NjCcYYQDFMJJjVKYQQ
HxWniqGnNK87J3sU0wHHConCLNr6Ov+9ceFlVatI5jhKKIB/GZ3xK1W7wjC6Dmkd
oDQFLwE8MYHYAg8fFj3X5ftI+zDGVqDbm/0lrHIoy6FV+WCe3RwEluGzDjkjBoiN
uwPxbJjufa+QI818BZArYL+mdvJSzWtRbAnaAsCH7R30FGo0BbeUwbrqKzgZvcwX
HcLA1cunjNyXC6umujY1AL1d3l+lR6xVOJkF8VSktVuTPA6fm6pSccPAjyWsUjXe
6Ma3Ubk1FECnnj5mXTdZ1wGuWPtRfpqMmjwojc5cXIE6DeoAk/QBZNJBgwfcqAA0
XEdyegxgOV7H26YQr/rmJ5jdSGKKOmGg+kpm/aPCrLhW6wREgR5li/MsZv2I7w1A
+U1s8l++Dlu5vC+8vVIxc3SkFICab3mQMOfriK7YKfALZ6sQSjz2rlmEiwSpvp0l
8ZlAcbDpymFA+Nc3wpt9NxOVWDJeY/eNSjAHqYk7vPnJz+I7clAoNrXTb6hhVdzf
lar4wDP9urTC8cLqntfqmVuJAa5qoOaLshub+oD4CD4USI87ay21WlEv+DweUNmK
9X2BSmTOB4HkbqiFkZcz1DNwZwHGXj9n10a6aH8pyjfXKCMkKCaLmbjjdE7lf00C
SX7bSXMY03oe7zuC8/1mJbkpMtQo+/n7YcRrCH8maTexdpkPwS3E+7k9MaKPSw8R
kZaNDRqocWyKOyVRZP15AGrxd8ZuFUJYGZ07HLC6W2kXA0UKQBCTQ9uUGLY0fkGf
03frA87KIApyDwOcj1ZnK3wqaBIFB5VyA0YNMx/L4A74Gw8hezwURj+sR5Qr/a0V
Jy1HKbqrqv+4YY9FXcrb5sUOAcs1Oi8gGDsSTX+vEWfyLqJ5I21ohip3K0LXiQeA
/JNGrH9FDjiz+MKFI73kuw9O73Zcigm8crVopMe15rdCcrcAX9zyJEuHCfc3jBHV
518wm346tB0xE0Bq0ZzWSQF7oCctzMovTKP2QbXNeKB5QUWGhAHsdhxo5ypq0zqM
ajO/nOASOluBDQLpV2141dLn248+J5tLy/krRDrZoJkRdFrQES60tUt98yPjzmaf
8PSWC0vejKV2xBJf72gQH+YPblAIf4V6+rjAOWuZbFGsgEiLVPRKXRbgdIctp8jC
/2wJr7SeiNtN74sUAz31fp36I1eeI8ZhZKldkKsmC5oOn1VJxJ3bmTtY4svvHILo
2txDNnVzqVf4sjnz9zDAWo2z6SXmcXfWBgbrWYG6I5PpdOEclBvSH5+fgTOW4nGP
U+b/70MnJz9T1U5WZ+mphfYs2xSuYvFQWlQM7f0+7Y98grKHyccYb6htGq92TFWb
+vbgQWJDnNGZOoXdHtrmIJj7LreUzCbREjxnZSiG1Kk/o2rdjr4aRk3CPqvDSGeQ
J9w2EcePKfoil/7t9Es/JBeacc4GPucW+HaxqvCGHgYk4tuuuNbt7X2NeLE1Wtmu
cpMpgPpBmxW9UnVMz0m7fB+/951PDVhtxx2zinPwVKt4bl+2xOChIWUq/496gVQ1
5U5UkeK2m5lI9WB44K/FSxHivr0Zhl2ob2Gf7C0alB4w7OP4mZjswVFAAGqBGWuh
OpgoZ/b2FFqt0Uls+Be2jjU8gi2m1owDL5etGkK+RUuaxavZBhdKlVgkIJhY5vU/
6nfaEqJATNZ67qTc2l3ZKkAPIj8K5P5fw+o5Qn7J9YB01RYeW3vW5grisICocsFQ
TN+rsb2nYpDxomCKsct8CZEI7JGREiIGeI23hQWA4Lule8iuBLH7A0xu91WukDpd
nD/fDY7TCML7aQnwgk9/1SNd4gcGubtDTeKPjoRDNR/0X4YpUn5rX1sN/C1ONhTw
Hwpj7rDhCBwf6YDmEdDVZRC1Z4SZkYmG4bDFHZznLCe0v0vXmld9qE8Wu0jMe8SP
q7ehngoQnLNVq0LZ3I1L59LcV56jmb2LS8dyxxQ6mwpele4qWxvDjzLX9YMlFSmD
yud+JHypZT6aSjWPpG4XWVjU0NiGk6fscGBOIyhzdrss0OS0HYhdni53x0+QOIIH
xbjXgbzEXXHKMOjM+S6+v6kPq2ztrWuw0l2VpzqL2HaQ1bqLvjzh9eRtk1UUzjT8
EXU3kDu7TSMc+BHkG4DWKWl79Ki5PYMznPYOJNJ3UDVXdI6y17Qijd1XiA5Z5xkr
tpSoUo7lTLsrDbX0mUTPCdsfMhiWeazmPHSaSpK5t0M30ZkucGGAVY5Mfe8wKtlL
NhXO7oBj5hwzuoQqqJPxADxvBWJVOt0TJDGxjHWOnhNCPlXat1r6X0RR4BJlGQ4X
A9yVmF0sj9UGKhUS928HWI137ilNV5zpe2IMtGosK+6uMYOBKQBen4vhYmUwdLbC
3M7UN0EG16OciQOd5KZjHxzk7EgrFrZXNxCQNuTaG0h9fu8BGcH+u+0zWP+8mfbx
bMASBk/gBJ3CMhv3cMrXKczFIPgwamgQGyHO9U/CrDbCavui14Y8mjTUHvJUlMEN
PAGQ6tdjyX8cU1g2LP19BVjFrUU1pprSzJ0E4n3iAG0TiKATBjn4qnnroL+aZG/C
ICZ3ddqsX9o3/4c7TBciqNiUmsOSAYLJMnKoMHyCfjXRvwqXzeuFZ97zBWoI2fT8
Oge2CENMYrW6gTpqPQ8QOj+7xHL3AMq5eTsonE+K2n4YZ9Pu+xuPJx5hhJn4B/YR
H418MwUK3GWv0SHfJDUa/B39Ej/+1RpAg+pRTmx8Ln8q3qm5xmA9ElrGi9a/jTVv
fSVTeiipqowm5QnMywa2cKTQ/5gqpYscWvasT2HxZwDG/9DOxOc4EY73uSbOTxMh
GAt08KD8eEj5FktKDayVzoZDozA1fMAa2WlvV/BOmAx1ugGV54LNbscFzq5pPVym
v0JD9mzGkH+Qr66nD/U5shHsePwk9squteR+L3vcVwJKbHIVNlXHQIJjIltP/IaH
UT2fUVlhOH20t/AlcNEH3ZPoWbJt9iXbq6nrE8Ww+xaJzIZasjxRkUy5jD/IjTOY
jHjeicNtpQdMWUU0jI+VCW8EK6brmFyIwXEuo2kX+kohBqmzlL7RjW6fUqZLb0AE
EcUe/6maXBXh1D2Ab3mhQA4i/vyzN6+kPEpxgc3sRUI/s8jhRyIZowEc6hgzmVYW
TGJCr4H6V7p4MZhMmnC4jVWr8Ubx8Z4pPTZOKSdolA1x7JAss5TodP0+y33A5Ucc
DNVL1eb40OZZe+m8buXtKel10rgejSSJgDlU9Ocl7ocOxJ7qTeHg6mjp/qBQkJqc
LLWU4fhFMIuFhX6SDUZ9KHzG29y4x4gn6v9wjHTX9oJiIhi2/urAcgMBGKE2QWVh
wj3P7PJNR05lXJGXOlCM0tzX0D+CtGBwCvUXnBwOm9oIhx9ZRbeknu65KSkNP2Et
RqGUX1xSeF+4wEkh96j0QjLBgbGVsvoOlKWA9O5LDruABNHDFopAoL/3fQX5/Bhd
MBw5VZSrHabvbQ35GD+EfTXIe6o3w/K8dvKEnxk5aHmZsb2cVQTOZhgXYcMExz2r
0Gqwo2NrayZ6ivXSZU5tN94VQ9fxg5rVi63JxqeHuM/qQcer4M8EFHZ4De8SKS3z
bgxErjBT4HPLDzwurw6GhIZJ45DxDiMGbfXIcSXCodfCterIn+CYhvuMQYwut6H1
iLnmslFWuwNh3EFg/XsMytWGMojqU4fPdcKdhc/fjchQ/QCqY3JXwg0rKABCEcJA
/uyAZCOduIQVT0nCvjDtMoS+4EzNspCJzN5CDP5JMJQR3kFDNUFG4NTvvkF8jgyp
LWgE7VhHcChkZUaJIV6vi0VD0+/1K0aVKROKJXb/+sPBy3eT4M09UXHVarYOu38G
9BCPHJWsPcCBw4tkEGlHY6G9OnrdxWjGhVNyF/L1vsPBPFZ2+2ln/o3MRb8fkMxb
g4bRs3Ugf+BTALWAu/AJrXH+uRtaZuzVb31m0RpXxtxCvzOMb3ea1SR6A6BtqUWp
D4ypcCmIwv5K3YD7uNL4iQYTWYDtwKN46ADClfgdFO/pqWFDeNMpZnWgTxakhp4p
CmfhQKByoYeZ4SeYVaZOgqn7+z93T/MrXJzdoNj3WKEOxicEYTNz9yPRAtxYWYI7
3CcKO6zVcAEc7V+WgiN12sB4Q/+B3xydLe0RNf6i2XHv/KIsBW+Ke/i48a8lMNcy
N2l3X5vhE+VyJB5vdJaHIb0ug+Y7an3V6PZTahA1p9nS86SEazLRck4uYYcgfPid
udnyRh4FOukp7g8XMlEgCxEU2wSUljXzwdHBiX+ZbuGsL3cuiPHmzWpHwdeqwbZ9
lCmiIfxhhPgWo/UoVuyf5jeNxsebY05+68Yt5urzB6nDXNz1qlYBPRtfAf2amfKf
znfDvUP5jutTfgcN+aYa/E2V560rqlDi2q18L8t6uPfe06z4fYEjXOHjhP5cswKD
PBHe1iA//x7PPp1FMQQQSKF5UyTufWM1XbRtIUN/1D5lZTxxEbhxgFvk6H9rlwTS
OutvmpQIeBXGMz0Q3+lFCUiamBwfXnuSPAzSrPVpBOytSkBJy6MJ0r/jRDvsdNaH
gsWI9O/0uVMQqzoEwMWsskKjo3BQO5dt03taYQTEYqqKXAzp4dshkRKtwjAUoHG5
5p45XNi4Z2G21WL3m9bmGjSeA8YSG8jVZA302fJbyHIgJBhqqIg/TxgOfXgumFER
mutcZ8es2Xnq6sc9Rq7oKs4mFoUgVsSJThZZABIAm18vox1gwoMsyn2XM8kIaGyk
sqeSHkQVqH/2vYrSHK+Qd+goHDQdFaotOSlAGDWtOzjoI0pMSsm9ly4+HVfauRZX
SSjqL8GYroURIv/ec2puElrOcF33Kv6Evg6kDEYOS+LwRO/AJpmUW6oWvkzmO1bV
3hQ9XH0RahrAQSZmGTx5Je3HIJhaz6VGiMJfjH10CtZTVZ17NP+BkGug6FfqIda+
gjK20JT6dWzbRBQ3qbgSswyhjExvBSsj0AdsLYc8e3ise6SaEB2hkCBds1dbKlGa
WH3f12Cupzu2xJbt3G3MzPN5vPeAAw7BOslkk9wcjG4mEM4RHhbVeVEx+H6goNRh
aFUzYUsjnHh2DvPyn/4wqQhg2WWGBNyn3OLL/yfspS1NCjZnn73I05DdXgNMMj2W
JRkZTtronSrMuULLlZfIwmW1CCVuMiHk1KvE288YmGWiJZnxeGwYZpS/oB5jmxtf
p/JyMoYhQ4RgobUrY/8Sn+x/Or08PNLvKX7ulFaRpAa8EK45CpA4OcXXF2rTSNzS
YUuB93/xqXcBhSIpOGOMtyvVNClXQmGwwuStsOdX21y4jxVSIRKPFXT9lYQHpDDy
JPg802NYYOZyism2TUGQ3DXviEt9ksSvYt2+tpnSpGDRLXlvvu9bHky2HrxnU+uT
9mtJM6U3KEFYbv62lsffHUNpPLFFpB6jIbFZTgfxuUzrG9WxYHGCKKKIRiXV438L
EBDMm6AkryZrXcptr+QcZWo2OOJRgwUdp0b4yvogcRfvkjqRf98hvvvl/4GOLuti
YOT3zUAIcTNCJkK2IqrB8y/LsZcGOsy83hMEmMLlyFPNoIv6a+zuuo6LREXw6tBc
LeEiOyhoMBjhjTHjGtdJiE6rI+xRLKESO233A9rKBJJnwzjRF916YAUBSsHZS68+
xs266Pm0ZIWBPdYkrXQrIF+qXYXZsMHqoUXA2znZSi+kow4bZ7Wzkrp3+63Aqqwl
evDujtEL+aF5aN37hPDoSQVxWI+hdu6XNrGgMe0BImyVWvQbF66cAAskLTScDV0b
WqhajrQIIdeQ+2lXuZmtIB1TfUaOseMhMEIIzQgQD+OsP0rjJvUEpmbReyXnZhn0
RudmT/M9FoUWC4/2/MBzmfd8xHuBwHLyJQcgWLHTh09czlkPX/lepHbE/1piibfv
PO3qjZ3wwPoJ0rHHYNgnUfkz+XbrPovn3SOhGCQy7VOP4I6fU5zUrKmNHjWGdrCz
fuYR4Zn1QMoz8ofDe9fCXjU/Ll3NMhaWGcKEsRpPjlcf4lLP6pBs12apuHH2oTNY
/hP2li8L4z/+UGWDmvy2BoqHMDE2WJhq0yUrTEvvmH0kdcjqV/ciTAQqy9/IhGVs
HcIOgg+lQP5j+sKGVVc5y/FobAwDhlvHcrhq93BGZIgyxAo3h7RVXIm+aWD6d+Mp
a9xEXHFIecJh/q9jC1qaEVhejQylA9xh0JQkQk00Fcpotg1OyVZ9rHCTmt1zCazv
zSK+jP0YdLbaofNOZAPzgJzfX1OEvgalUmgxQ+qnIDPeH6QSlU8CCeCd8xd1oI2D
mIfJhZyAjkdpyPMzAwTbwiI94kC5DRAyMDhv4bjRmJVvtXchtbDBWmi/TupB1Wk1
jFF3pr3nLPLJWJNlJo9sAA/tI+VvaOqKgIFkqkMpZW1mCW53RnYCWDPOTnWE31+X
Ofjmkn8j33oIX1nHIuRYlItVGygvey5AXXvtTIe5qsOt+fb05DpspVLrxN95B7yP
Y80vobAMBVa0GSkiT9eP1Z3RrMKA+7HkmKGrXLVnVugJAkiK0eUV4UeTQtdTtV4M
YX2pL61bHXlTXnKJ7Pp1P8X7D5oLxrtKb5v84T273T7X7k5lCfhFIHel1h8eDShZ
Aj07opSIJEpt9uMHF+vovJIT2lqIYj4RRLRCo5dbjUrQxk9gewnVUp7uJ2wpvNPF
4ZA9RPQ16irYOltQlxbR9VKQF1tCoMKZp6zecH0T6jwpXOMQFIhQ1WQsFdgLZkOA
5PAK/UVTOlX9HIqXgZUQoO+9wZECbMY3RNbTa8en9Ay+yiZ9QrRmZHroZ3KGCbKH
0FvNqN95kyZkZRTwKIH8OmN4tQDSQDLfoZgDR/kS+9h2T404zr8xM7amQpPscV/F
NOXaKIMYfb8+HFwbrcWi/rasgyOEPZ/GFjRltTtlWFAXdsaoI4YKSoMWy+PUAxFo
DI9no7tDWF4JoRGrEUld9SASzh3kb+F8Qfu5rmPpNttW/IIZMOgGOa1oMpuhmpPH
2AMyIMmHrdunRJcsMmR4ijR0fk1obuRu1BWizU9xPrOQk69dxG8TpBO9QzENwpa+
J+tFMTLFBXcS6F/tbS9H9H3rqXijC0R+4QTfOJqjTdL3iKmb5cyv4kHN0r3P1g8A
sxL7Z8Ku+59wF8t++8OEsrLrttO6KMq0tnRzsh+xGdKmYfjoD4kb0jCBW5WP/6lj
ELPXAVY5IJhY8cK/Ttecqb5l63baEB0kBU5c8GbGFTIVYa/UcQLMYBcaJbHyAaZS
t9dXYNKvLOYWcvSaCejrULoktws9Bj99ks882M5r1hz0L6YW5oICcxjxS2qtZ5Bt
i0CXQVIia8LV+xYgz9mcViTackU/Si/jsUp3o4tXYoXjN96zlhBI8+tGQfncVKy6
oiiLHDY2+dbYlpUamfm1TIf/OAipFJYYsl1C5FJi1KFrVI0+PvLBC7BpYwPSEjBX
Q6UjgCsduDrXV+tk1j2ps7gDryGvmDrPkpEWcklheQIzHxe0ZpMO4d0SoC7NmguP
bQD2kNQTp4MNTArpraNhNYaG8w1NIm1B8RhT8Yy5iU+fiJtb9WLptzZ+g0BL+alx
+/Vr+7s1TWKXxrTjmr0MJV0U67RN7T7eofzKrbuQVG+C51JTj0jJAoNY9Sa8bcTY
jY5vSDkVJ3uDvFGH4cQfXo+5dHPjTvqjvOcnv23kLYFSEQ6HUpepnxL+3dqhgWnd
1cxplB2XMnSEP2TqEgQMC23nOIjz7lIB6M9A4HZaznenEDI5rAmzH7f+o8KfdBac
oDAkpiNYyQI9/F6MwtuwHpsAKtjij4mUdjFjACcpJOtAZGAP1wz8IOi1FO9tm0dn
FVTS3mHLI9Bz8Kd+2qmGo+B3Ttha1HQYjfQIIh8Vh6TASbtf9wNyCMF7tJ2trV1B
C48ISwnjKSc9K1HrxqhCqZNNasDx3S2UrAPQURIcRqspANgcN0JS2fsKU9EvLYEa
ualyxquuMFJIr+7iYgc1KcgW93NwlZ6SdnhUio1GQYtJrXOfo7TZnjFy5jnhQkTt
z+DG1vbpuRjZonnkLpJ4T4icA6DOnxRF3esSvcziP5LTN9Bo6+vpJ/pHqEG/3XsV
8SN1DsDPxmsQDyZGrf2e0tqDVmZOCZhp4rPQ6JNFp8oxhODJ7+V2MrV30to+d/ac
RzoK8oiy4rf45LhVYJ8wyT1Fu9rl/qdinLR5dfzpiOFR1ZOfJXRqdmAXL5bhvKU2
edeTy8hyeNFY9atTgLqfPcWf7IkQNuRG4dVyveG5jXXnMmOZA2CaI5ldeUqkXI53
OzP0OGCWJWDfEeWQmuX5A6YPBcXTH+kDUkPXinIO4BHBsZa6KzBGhYACery3d7fU
aCDN34nINszC1z0pcguGQE2xIXavlHtFfg6UWAF6MQirFjkddPdN5Jo8fnSQ3os6
rrUQsD5BwEco4WUH98PXM/3v0Ap5PRvR1LAL5xRqndd9n2lQFgCyUWvEiJLtNpXO
0j6wGLjxvFs/4xrfQEz0DJ7PG0j0YOTHUL1GTzACMcuXU/0k/T4iU1ZxQ08okMEO
fX7X+AWKjq/SfHNmv6Io0bBLUN7+OYTBfSLIWLQKxIVlxnst3CiH3e8yVJmfCShS
/b5iLSNfB62RrqDi53HyDsrwqzeVG7WHV9mZeLCWZD85HRz6BDR7SwjlBz5tZJoA
EWRJnLOSNW5jPka5nPXBGsN9I5//5rIFXZWmhxvXNhsGBuyfBqVztDrYdiwBbXx6
vNAQk99B5szvzJc2EinTGoHK9tJm3NAIfcS0LZgnxAqFtEfCuS0W3lc3RpOZbNty
LrR7Ivf8YqpK8iN8BKiMKKci8sz6TA5kRpUIfE/0uapIe5ytcSM7YKLbKzIRVXd4
aAfAWMuu968Qub1fx/22YCaxah8ntcUuFNRT3N7JRFMplJvhn2sbkQ0OTZ0PV/97
1M1n6bW2Ndx4VcZc2Wub6CCaxJgCjt6ejcV63eAjs8gyVPeQ3qIKXHNgVovGApJN
wNzxozXzDuivObucqhalzPuB38qRNdWoY4LeSCRNHH9csHxcH13WF6MD0NX49bq0
r/kDmSi5IDJGLiy91IxZ+tvLarydKSLAOZbhJsP+yEZfX3+9OhUP7I7v006AKvnG
htvZwzx18JaGWRmDCtHXyGFgER+yuPGYzVfedzQO85UDhHny+5auxJBzN+e1wOIv
KMpPCxEebEEGszHHcYvgM5vEny/AVe0K/qmRNrxeElfFbQWB3OQOZQcNj5LsuHLm
kFuL+YbqV0MrFGMZ6f96XwJRQag+wIdwRtnKKu1jSJPXy5lf4t5eJEDEf+7zd2JW
smoGz3g3im5afEJ+YxQjcl/SoC0JOx/tCxlpBc8k2rYxoG6TuPV9wdlVpkrGh8h3
Nt46E5PPiLashhxuYquT32vwhNnFdX1a+srlfj1EfnXeHM8hhR31bWiADr5Pmxmy
QfI1+eUIzsWF8MvsORY4gAQGxq4cIFe5F7+SxcioQmc6h3mSbdB8tr3fN3govyI7
xvqbh2vxYgMSjoS7Ay7V2eYwhMd7kbjtD9qg/Zva90GlLjynSj59vrJPKXIvOeQi
Xh1NdwQbOaBFZnacAzTZ4EfLcn1vrfdcYHe07Y+MczggP0tFQQCRztHzHswTc8Se
laRGSm8XdIew9OUyBf5uuswE0iS6WML3LfYTFRMWI/lJmrXCmS5jU6a+s/jtWB0O
LIeDq6LZAdllW8N1GL8P/OUCUbREG0fWdoduVsUKF9wq8mpGu8XdsKSaLeKDJr9S
2WNSs9lfjLrwcP15iNcq8ctouvGdIU6Vekdcr/JLWGo2GIAuE0H+Daa0bTiuDY4C
Hn6nuWgftw/5tKNWrkN1QbGndEQ0cA/ocoFrJE+hNFbiLz3S+xWRHFgamSARSLjs
ZAnfsFlD186o5BLfsmjSopsdvBJqjxgeHY4x0nF5KKRJy3MDeCfGnuPoMXjuTKsm
LnYLkku8CaUSjZUiD0xRaWEq1rOst/beVlOktsB23q3djECV2qoSyfRxb5T0ihIq
nxSk3BEQdfIi1z1x3QxF5H1Ej+5Xi9+La/sgLPHyR23hqQgkLoROM0/8DqUFD19e
dEfhT0JXyAw8QRRxK3fPqDISXs1zJ3+cUU23JaqQs74RcX2e5JnTvS1ZLU2NPNuX
C3/uMgGFyCINceo2WoVpgZuvjNGRn/4n5xodqkcoD286E4rJdlgexsc5yMAGI4tZ
6xKzfmjWmSQ3EmPjam3rdLoMWkiN0dSo7fQyMlpWoVTiVnXnl4afR6KFgue9dkKc
mzGnWpHRdU73w+qMkAPLNEi5UzBfjLvL/vVH5ae9tgX+8NP5J2XibgdcdRNxfcP/
wl4AKMya27CYommsCdyARaPXmGUF39b7bImjXVpn6kqeiRXirnHY3l+HuX0wog3R
yLZBNKxyh16Y70xDlg8+ueEfuqJiuY9ZsohHdLUYfbAppXRoZfMebfAkED3vXInv
vgq5kG33pWrPmx76QwN29JReTZKcSrdNkJoWZdMNkaDnAo8bX141dS/cJCNHTUAO
ud3+7lqr8WMs/xk+i3AD3V7jgZFTagm1srevKzocdcDICsVu2DFT2VqiFm+mVXIs
FbfF+a7OxufMR52Z8IyrDxhZaac/ZOUGbpda7hnBqejL5TGt05ncnAdHHXNMDX4S
AlZtTjxVjtttRO1u0MIMsb8NDyrKZSC9ahm2FPkW7sVywrOFju6goBh3jnUP0HwY
/m7YCSbCBsNZ0m/l3PEzJyqTrk5qLKmEePXVdGpWt17G4FWTUnNXbS3e+4gy6Geo
B2XF3LI/bKP38Rk3I6ftD/FSwZBeTjsLIJgzUQTm688lFknbHZ6iAiC7rYeudx70
vxmQ8ZW5rxXn1hCu0PSRsJWze5hghVQaR4XR0suycPp2uwcWrE7RgC2k9bMmMtqu
nIbq9rxJkjzqOAiDXwsY2Pk9pJXQEJB8SRYclVCXbHYUiN01Ul+imqUvEk+3VMKq
Oqfr4tgInx/I/WD2CJHdIUri/7UnJTyyCedcG5ifTvPC0Fm51p23tJ3cf7ZqXHzX
KYiZ7DvzdkAjaoxOorauPYVfzwIcBvOxPzkuMpXemb0ZfDzA3XW3sv+uhZdtnF4R
ki90PodlD24lSQ+CQPPqHF5rWUEg1qiYysf75gVNP0+bkxSWtifIbrtFWq7aAw3U
ZOkPMaEznbwM+LeP5lI8dCM96AaJ1qJZ1DePkEQjLkzwOcFx6pF7FcLW6lhVnfmn
QqBn/qYTbbdLCkNtUAxa6JoYd4Pm6SX5efnJPPiQV1RrAXSzL+IFNw5iSN1QaCvm
0Fxem0RspNBu6mHfAQO6jwA1T3ndGfTlYsWGvo51LXBF0JpaBL821QZJ7DbEDheZ
0kjD6tVCBJSe2bQ6QU4mQlgtQOHPxtEzhsJ3VYs8GPQu/nka5kqb1UZ1eB/blkGR
sXsoC7cpHPwB2MpuCee1CBZMCpBqKxmOoqMp9i/w5HcaiERaXWuHxPZr1ZAmVAT8
YW+4lMva5a00oCwqV0pIxJFPEwkx32I0FbtP/yeOMMWHFkEZy/LV3hhJSWPw3Hbt
B6a+EynH/LNLA+n9Vj2oLKHBjjv+KpwAWnuxLMHvAsQsB++cIqL0rshn+MTQdMUo
NWSXqBH0rcgarHqEeI8L5nAb8n8h6RVVuyuUaUfdzxjxaPNzTjHBm7XHCT+MGG8n
GZfjbiHPboofsTAtu29uBnEtCpW5Ku8LJ9UHK2IAQi3U5ZOLmeifPhslPD17sqav
bTX4WEQoUTPIzpa6zwsqKIUbCW+ZbJYj6fyCqEW1UFCrsJkdqVwO21X30am+gqa2
L51SlZ0ESA0NHi3YbLlwZe9hCZk/uz0BDALdsgQ4g23dpjb2AnZbtTIKv9Y8mcv5
b5YwPc9XtnAMOuqOn1UGqYlYqMkDIMHg8b+hP/RiW6rf24ORhoyws4I8//54UMiR
BQY92SEemZdU+/uCsyajIY0C4ICcMQPEU/jGHG4VLW0zn7Q4TSp5JN3YCf3SJJH2
I/pDA2zgJ6zt113YwDH9woJymCaUMRERbIzB/ariWJqdlK6SNxdsKCKhC9bKZzse
ASLGJubQfP4AfXODgc9c+lvblVPmWK63bCziuR+rXTDIwj9uLPmVGo1fCoRVpIVj
u/UCO8SoV3p2OjQuUz+a4E2ho8peit42yYGmamH6JpT8SqEM/o2XlwvuqgBkql3t
1n7xWpUeA2OY8/Y3jA//Y9jqxoX1FO3nEoNynCrrI5Awfqd21tt8bwQ35suY/Vcl
MNRUT8J0CZwyAce0AVBAWeCkgpQU2YFGJK09FX+Mmr90kAEoYTyhg0U4sy1pQikW
4BJsBvQm1SHyNtk3r6crewvU+nJQGA9KgjAlgoxzXSTkeTEVl/yXQDCjwbpfWeOb
AHaMf5jGQq+e1qM1FcIMPehQdZC5UGfR/idRLi3K32Mrto8JQ0i7jCOgymC7bVV0
Q0uj4VQ93qppYvvkMlLYMoNNJI9b1Gs++gH92hrjUeP5JDKZi+gg85sTOsXcqw8F
KAxkemt/9LJhdQ/oQkTqomUbU/PAeOObf2QaZmn5PGyW1/FEsRrYVKkL/q97AHTe
grzVOLHTfUH+UyP9qqo1LXMuhQow0wH+KaICTKBH21S/CUIa2yvA+G3/HSoNAFFn
9d2gpySjzDusijf85Qgey8a0NUIOVRKoNTriERw068svjdJOphBZsShh2o7ZqysH
W+Ps4Xvb40izmTWRy48mDvrb/48W2ys7600C/Blc/wSRebfu7UveqsLEyINfWo+I
WB3l1FCeGk9EfCX/qBHUkfMBZtL/wHGaZuEEczcor23FsoxEWjYy1bTFH+Q4WoZM
tqDg/cwYcp+HsrLUw04JhLBuLiQ3L2lCdy//Csgrg9yIJ1aF9HtsE3EBDZurWXtM
eat/G+4neFpHPPV6rlkj6HgmG30gQLkNCkJGPVHvk7sAyhYC0pbR9vACY+aHEeYe
leIUccU4p31LmLAQJx7D7bq/m/J9WIZwCXNvKxT5Eo8L8VoxfmL/UbSpO2FV4mtn
51srg/LxV6HaBZqldD/TwKWRI8/ZfrskK8q3IBp1uXuHsLNAaf0QG8iVB//EczlQ
SbnjVzLKSanCBBxf0Wxn4/dH7z5Jrc4VNCcVjWcCDCukW5D01RMGQzQPtbmdl4/3
2MBpcfi9+GY+eKTUgzhlHaQrFdtVFvNcb8DCCpIsLxGA4ZYgNg0B5ZQp3/kKIp9j
fC6ny8tfl2/ZfRMWFaz3HCKa6c8yQf9PUeoN6cJecu03mJOmjZ4erMdxxchkshmq
tn3l4brkoVI/7ysTvbnpLWIWQBm99+Aa5kFfaz4d+phsv8aYeGz3qimqBD1ij/ex
BBZKDuhQ6s5QiRtoz8AhMtFxTxuUEijyAsac6IA1ImPf4a9UWJLRG5Tuao3tC1pK
Oerxv1jsd8k7Seu1wjTjwnN22KomxSDj1y+jot9vNBR6aTyLd6J/wGZJvLA3JCAG
8AB/E/HYMuuYrFqOPD67bd+gsp/LE/UPjqk2WyfELA5c6XzW6mTWA0caJt+MF1fD
a+yE4MERh7QuBhHZ5aIxsysOzjoJug/5CdDWrk4d78skmqjcMeduW2xwMwm7E3vc
dBZpUAVAXBHRGBTkQWw6gOcdIOvwWNtfiH8LR78Me/dl2iotOqDwaeeO+VpsPAI+
g7oIVfhA8Jf5KCfVFcMIzK257bhP3UMBlMkkaz/3MzjgDI01MZWgepHngrlYsfEz
OWqxJcl3b85xEpj/5eqoEglic02XXWcOb7yWrkd6aIXbfalJwejftpuFvbRmDtdZ
dJmVJkOiQKLad66gVBajFCLFUUtXgtBHmHjAGI+XA8BjZpaxNiSvXI6a3pOgjZCG
V7nDhMTka1vli0+/u8PZseEtSugOs9S13aC5Fs09vZTcCOBtUqfv8G8a2EKkgfrN
VJgyTBuCNi3mWV2IiUR/XcafmNaq8hmXRS0S73cR1RvnBgoi9lK/R00ctO3mo7ZM
P230fbliNVMfpXKbTimFC5TsEUyYm1ITCSm1o6xOFxHbLpzjF7IAMPypPKC0xw3F
63LTU0OkiMTt15VcH1fJ2V/IpkGRhpPGmWsMXRuOvQaFg7sfPTGl4P1Wb5VDVQ4t
zQN1M8hvF24L7N7dSkD6nns+c6wIG80ZSEqkDLvn275W8c4ctssOToOTkRvPbApm
ew1L12SuMHydAozrEZXBx8bMo/q9zScWMZbPCXo5vw+BMFOu71zeoEYX04X2i+Oe
9wBzhfAipGTAZtntXglqwvLvRGQ9ZYxhMWXg2J8bp+5NDmXMENAsWY5gPpHJOVSK
Nd80sKM3ZTsqSezi8urzz9yPTuXtualpmnTp25Tydrj3t+M2K5eKHdScoIu6U+AF
PY0HbsrU6Okgdh3V+ZYB48RswXMzTGI3oz3QZ6hqkxw8UHN20rPek1ppU3y7XGyB
3X4hHtdDbQNGHS9VZN/jS6MljeG/+Bmv3VRPL6tcuw92ZS/vrOwimoSrPS7BrN/s
ROoTFAKcJkC0JeqmoTfuYVTaTfu+2R+1DbP9kT+76lt7JpIgf3FG/2UhKjqI2n/q
5klUOnMw5XbipXKVOEpBWQ+AaJKrpfdXnKV3UWarnmmKUkFWe/pAoWUYKM6Hp/hy
gyChtbMpNZUh9cfFzGj6pNFkbW6H7R73K74hT/6iVEpcIUqVCRqal2Pj2ofINS3Q
fZZC5kGNg0yZr/CluHfnAIntVa3ZelO4bwV6nLLhMvTIeMUk5jD1CVL7Xp2Kq8ll
LKQqS61qnwXc/0ApMv6o09Mh905+RbcrEd8W0LMNjZkLBMUMRpueC7pwPWxzdO8u
D9+xVYn96cb/o1pHIPVOXipNI/r+Lfv4w+PC05co4bvWbBCtw2idTiDlv+er+JWC
DIZ06zbdi9AYlyPr94ZPZyBIpUTlDJWN62un/wi+PIds/enMcxKavU6Cote+F4bf
yVLfweljh214T+r26fZ7xX2G1BYc33q+UCb5Br1pmRHPzBT2ars5BY0q6UtqrBMd
SszIS1AaWScMUJbjSjrP+Obup+Uf8rtiawCIACOxtjHseSloGYXJSLTZpev06gJM
rDHYaipVjKge4FRLjIOE3IZb3ZjY633dpyKQA5pAHsWgUbJGBD+4qlkxCXKy4BnK
zSLKnLXobcWwVp4Gk9bXwel+ODxr1lQR02B10KCp0SAO5MB9AxeysCykLYAMSW+N
jHnNa1q+VeyHM3EfUlRiiFE942Mj0aOgUCjXsmZqSLsSXqPo1FM6dKMWPjRav0jw
K771fDmL+WtFGtuZ/DTDMOJCdIHA/2VQEQ+Y8BFbdGfac7PUq+pLhsYN/nBD3baX
tObf+bKvM2nYgOhb9RezF82OVkjGhar50Yj5YuruzhWbCgz1mNCaqNpFgawW3hX8
rBUsNzXkXEBgAlWd6zvPnM3850FxBrcaaUUnPcfupEArPc6P+8Frx2JZASrX1Xp4
X1RKZYd1xkxxSPz2rEi5yP7j9My5aSS/PumA8aGi8OzeHJYEHTcgo4zXK9rBAWgT
Van1+Fgwpi0Jssh3Lbz5lynEfxMcXFC9/hvC15iTwwnJ7r9WVXfXJ1Vu2h17QgSf
jgCejcOSYDPWZ8i3QQcugtTukDMV+mp9e03iVdrh8X66jijKpEMCIyWfmzFrVbrZ
+8zyw9TLjzPBoOLAfiBuMaOG2GMoMTg0kjSyzZbmd6ZC39XcaPfHAUGE36yjbaFC
Rqlk/THiAc0WcS+uw+IUvVe4aHogh55slSv2oBIusNTy4nc3xvLTo+2cO8kMqSKm
duNP6I+gzezIuheB+l17/5otFSjYED+gocw5Jj0qKquau3WnpqEJuXiXngQiIl53
1kuNA4z1ONFfefrHy+ELrmH6suVXDAEYqTQOZZybJdbVqx5n7DRyl7XeDezgPy+A
O6Nvl5KQ02OInMSAd0cQ3yLoOYcXRV9OGMOKellpZwjBYNAVLPuwfheT3f3U/MRm
vpyFVoXqrdbufT0h08rqD1aojLBsjCORLIQuFWP3/KueX6PgcXEfUzccjutsKMTC
NKqNfMKEleBaX+c9+0nYH4NE3eyOjVsx7cInOqfa9HMma/tGMDW7tcnXVQNCyATm
JkKLcz/0yyaxeFmo5cltIpK0b5h8Aa8ks0LUPw3Vr7/0HAExoNdsXGUoR6aICIrH
bK3W9zirD5TqZG2aRA9WG0w2ULz32iaLzPZUgC4YfA48PNtSFNLXpKcsLdqSRBQz
1bApf+kIynKarF1jhsQlVPQaUfUILEwgh+RRWLaKw5SRSApvHGr7zTFIFpQXHKm5
DjuS94hSwFfQdNsOX4RGbrXs7T0Rp5M1KM9l2bvE6/sRa7yz1TToC+mDOXsVbvqj
aH6ZbuSZiHDKdmR56eAP3ZRVKRPsUPc4UtQtuHnGuPY6/OFqkk7hsEcCeDNlYmGY
BnWkXkhuujpahP2NuiVJ4leZFNYYtCdTWcsJn2lIeJC+x4mzM+TxlZlyrn3P1Jqh
kQv5YBY2lq9K4szbrjyU2V8zl5/knMHG1GYhauYZqQAel8J15Nu9Gl2Nrv3R6maL
B1U9WC/pEDLBjLYFrZx0im97V+2Op5bsYofkrjXco2sfiyrx/WMMfwTQjG2VsAF2
FJX+vhvUelO8o6p1YE7ze4L/CTCffBx7pRCf7jyE8IBVBh+gwU8lkhfWWZsFKq52
UGGNfecFuTrZLSIpb1V9FKHJQTHXybXJ18MkEa7iH6PivGpYX/uB9hxB9US6Sw75
erXlCS8fNmoOfgd2yvtF1wF/8sBR4ZOH71pDMq37Z9hbz182ltT0s6LK9cmVrDey
mjVLJB7bv6watUkSA23oV/3ksIN6n+3JCOpSDAfexXRUGRQ6reOHieQxchsVwMQI
gcOrKMTAP87c7TGMlTqz4e3fTuCMTENsia9fCxB68zES3hJlK/+ciwQ9Ci2EN1Zz
qJ3qLaBJ/hCHrYbnWpcI02WVT4zqc9pyjweaElcmMCGYEGmAxO4azacalC730eKw
CW8tuRIkuxpeoXTIGAEd5SnUUfw31V1ojjY9Fq2Yj0iEU1U0O9uihpWOVs7vAbje
WEieKua8cZvR4N2CFvbrmJlcf5JfIxAlLk+xVnbExpnI7bcawerfpU4eD+of4uAs
HacuNkrMIv5qeDVqHTqttw7gjt+o1iBe+V6Q/McYG7rXNl79IHdKj+cAGg+EZ4ku
LYdKsiuJPTihh+aaw4+r/t0j0+h2+FMMn/hIK/GMsePbPFig3yXgCwUUHiCOVivg
yCxhLyvg1v3VL4lbpHFMA9h8WJkVtixklOhp8sej5rl9Bjs1irn0OafB7JExOIkV
J4cpWrhcKb4HKXFonDPH4Wyal3ajrhituSUb8BRCGMKX4T2sUK/chUzYGiCY1mju
xSHbjyB/AqO7RF9u/Po438n0Vt75IuK2rr2wbYQE6DO/TE/pYOiASS1YvMO8tW4R
mvBs7UwAc8Mar8km9STX+q3nekLUiVW8VPnoZP2lwdI4qYbd5fIU2UiU/q6AixI5
2p9AFEQCnFIxaAKFhtSjzK+mzFiOv/+XWelhKQrc9PnJCzihrapZLeRrpI8OlclC
OemLYkKN3bOfCSYkVP4zhwvKaTOQqpLKT7mxw90nVk8ou/lwDM4d+5KIvaksaBsp
9YGe0uXUQx7B/5PgDokOCay58ibWmKggs8ejjss/If/NTtgM4RdSAFQXVpiZ2Rl3
eZTg/M0DBePbzc8j2c0CPXB4tIkM75dngzC07HD6i4OlhGciAY+KrIJaS2n1RxMN
b8zUCxhEjxzq9gyWHK/s9W55Qbir6PGmmoMqfPuL0iO6hAJuutRvQC2fKBNEYih0
cG7h/Ut+D6azPZpv5kI6nPjpD5eE6r9PKKO1CYHMCf3XR4TZFkDkHfy6DYI02Qmp
d0FgCK4OB0L1NQl23HYdnC96Of0GiiPG+dBR2t9Mn1Hx6NSXLuJib2Dem9uXCfhK
G4QBoz+xItDi7XFlz4Rp3euMxNa5xjGyYH9m13G3vuftMDukY8T2qKj2UI5gYvoT
E1fjYYVJpxzMDcGl8aTtgn4Xa8f2NGzRE9xAfg1yWvG02maREJqhbn16y0GID3hy
izXfG4zdTavS9G65yUOCBZs9kKrhBJcfYUXkfjaP1uSemgJo8RshENfDoPCBAgDL
T017yUrUYXUHsozO7pYwQFI+FXCGxzS/zJyeCVWPI6bB43HvPk+PS6MdrqrWhN4l
W+qt2J40EOlvIYwLDt40DOCVhxr+9UgGpSa/nLixl15uIk4nzfkLaytGOuXk6Ulz
iXOSKmRgtQrQmwpYTm0OqzniaQ/a25MLtRQ1XkoL7RePB70yinsX6v3UEjRp2FgD
vq1kHZGb+77N/gG2+tpAN7Cq1k158J7vI3q9N33+w/mQhU1Qj/dO8eUpXRyoTgOg
32yF3XiHOLFK6XjyehsYAGsZeW4BnkvDD56MERbW7sUIAlcMuspSYIhig7CplGpb
K+X5H9LyoT4PbpCLhVsE8HYOX+N7xLy3T0zsJtLV1zMOB4mXE6w272tep1UzStxl
eaOpw/nQIqW3YJELS6iAyRdklMPuD8vR3PhJBUJh02RvNeJCgEMgBX8taIXOXieh
jqyfKU9ggTl6S2wZtzDiuSsPMHcrV5aTVQ1ZLF27n3jBoHKCFRade7B48UcNQmgh
c9lEQ1msvrsrZVzAaBHQUNggBABCLv4YK5RAHZ2LJBRukRtPIgRGFRM+P1SEy5bq
8p6HQa2tKh2lhQenoYZIRjB0mvZWJSS2ImFDK8ecUdyy8FzLlus3i+pqi0qJ8mf4
4Xd3+c7gJYWBnnRCo8j4b1HDTGOllnrhCA5WPXNmBuR+cHYknDvEukDUq6xRimV6
dMz8nUNRh1mHV0Vp7P6vUGkyGlQZgzWRQbsYErAouYGtyp9BYdvonUivpkiZXDIm
Y3c4VhqeEzU7vxPU/+cyczxaWlanBrplOj8tG+w8NfZn/VwevVR2I94XyAFKwHY2
VbKlvWk3mMZPt8TouqoKeIT5An7sNWKgSSpcfWsCS0LM1lQfKkdxYd1IhxVtM+ID
hsBNwgB1GLi4jhkLeu144D/y+kMFymN0fW45pJWyJPq23auCvlGBYei/Igne2kal
YBcQpKEfiCMdYZ4pvLV2wePXDw0SLvn2BPTC9W51VljEuh2Q1NRut9O5uGOXx8w6
7ieiox/JH6Oyzgc1nGeVAmlCA+Q8VpWyqXXYihMAoOp82KeXiA4gdKsL7w11dXSk
YRwLuO2juGlmS58qi4KorEnOCtgQojUzUWn6GXg4YvxDydKlUQHvgpxa7KNQAjam
2nlsK2GjyW5lry85KnOJRtH1lRBzBbiLlx01plKVlPpQqU6CH81NJt1DU8HgYcil
6jdIv9ijPWvVQ1mp7DnC3uFdsp7Z5C0eiwkz9lTEUP+oT1PaeR1Rl1/zKrw2sBWw
Dl4DIeY3WG9Tu06J9hGP3mH1JwlNLYxSeK3O4Bu33CFO9WWjOf6R5Kud4H4ig3qg
SRVCVjoEYRYcHM+l3rn1yZiTuomaBjwWE+MQ37UikeMa9eSrKp1hdxyxJ9WaFeJ/
bDlb9Xa9FsRqG08kVetuz7VmsIZEDC0owyYqTZ9r1b6X0W80rYuExj4NS/0Vsspi
PMEzjgwfeGPqitEspzxFZrmmak36aX2fD7Dg50d5V0Z4VSzci0AEl0+m7JbB3Bqe
hGLl6d0Q5KVqSETyituSpgl70+5uTpR/ORCxLYNAsFDuf8sKfLYdmFaa7Db0iqVx
HnQUEJ5E9ENyrcUyXnvs2XSkSfnD2sxsFvY6rw9ZlaTQEtmr30xFDbwWwOrJB/Gw
dpZ67mVWVPQS5yKvvPovHxVSFxMTEogtplrkbImzq2rVyZXaVlxCdVIKavT171A7
0QzFVYvV5MlOkofzTDQL/SLjQ8nNdDTQvQr8T0EBv4FoJVzdKXA+46wFKoNkxnB4
mWfOVzEYbvtdRt5xEmiEz+DgcR+AzwCzJaYaXKetgyQnmh/9rGe7W7VmRY7OK5F4
fulsK5D1OpvxWZbN69qo4nBZiTZsR2a2VPbxXJrHWm+CAKZ4ffuk7lg2DA6fkyem
eZC7V3N1lkxrWXlWhbVUulmpK+X1RakCy6+0Hjhu5tWiLsbC0+HE0IxZpD/Flvgn
AHIBd+/+qI25J5xLQPOX3YmC4gNCL50S1WPM3YFOTJOwOmfcDtATGvPvEHzDCMBX
gFo4YKbKhMfK1DZOCy/pSkzTpMbD2a5RNVDJOeyOv3a5DysXYT+ojp2WWWqIoXLI
igaUk8TRK5FHXp70rOM9aG5mb6eY6DMQu1+vFy/wLXwnhjbXrO4FOYsSsqVeE70D
kHdVj1gDoTVXFBtDkRPiKERAmFeJpFKrpXWGorOFUnpc4GlC0BylDL2RIPM42U0L
BTRdy11UqRfYKVEuOYIrH5XofWkCaEmgvCXWJCb7npDeBWJ0YlEJxf2ESwspC667
BMtJADcamdskcy5s2snS3tOjcN8RaVnZoy7WDBoGAV7hjPANFUEUnVeqi8bFRt/4
rbEitwGos3UhODIoUyu1eQEApt8AKqPiyZG797MbY5Yj30R6fXt/c4+VzztGVypP
j2A+j6a16YwnUjBK4EGvRjNGUe69mRfkUFrL6YV99cwV05vzwnFMDBInjchQj024
dNomWKmXht/mPVYwXrEV0hzeiBaruZZtpTXyfI6vbazlz5fU+Vknhqt+UePiAisd
vuUoIuNvL7yM/T96chvjJdNeCPYBeQBLONn9VqLbC/14Z7yBXs82c+V0SHisMY0f
tagx6wVN7v5R3JBCNuXeOR2fA7oNQKwaOgsH6VjCpa2bIPWrBURl8fJcsDH6s76k
Qq5COGKy/y8c80o6hXWczim53dwkU7WJ/4U6dMLCpiyjCYh8j89JGl5Mn5SybW5y
z1m1UhgVc4mfu1dc7GsXT1U13fH/KfvdDHeyGfMAyrniKpnu7UQu3AZGg5G9fhKD
lhy2HHOmBulnONmEBECd40AsFlBYGOKH8oKJbb1L/ScU+0a5FhPeOvfauAGuzDry
lVF84nckEaxfiUf748P1JFBog/08tkeQfFutGIerwuVqGg9mYeqkLTBqzxurBsJ0
oh39qQ1XHEeNIpBycryRZZ3WqPIdCCFWJuXezIjkMrLIw7v/MdEYHfVofku9X6Wi
3DTXuXBSoWcwBMG8847ni7IKDGsCpchI6CKAkMSVc/Q73KidSHBahvPMmldL1+AN
N4ofT6ymmwxpnS6Xp+YIyvdpiftLxLvhtvnLjKj0I6SGHJe6ZTx84t5D/CLi6K9B
C3tPy6HWqiHbXsTBkn89NQCJQ11B7T6WSbwmdt7v/9xQFP/RiVI8z/Q6x97gBpMA
xk5eKcDibXZKraO/+8hRQUZM4QbHcvKytyH9sjcRqumaUTiSRqoa7bEPAF7cx5Xv
HbusqxLeWo+hqfuq95OqNNZknJUUK1CzTbkik5ijYpQWrqwQlH7BxoPwdyLXZrQY
uJqOrAcAu31NWfGEvSC8AKrP5PhJvnnxhADAIiTO0kTBCD/Fjix68+ZoRw2wcuNh
QNKTDu+mPuDr1TGMwEtg3ZjNXgWyxk0e7vAwQZ7rxG1ZiFQSbDWG+kEaSm8ZaE/y
jN4eYjUaHnUTdIp5qV93zx/zlDWU8h5sriacuqOsTfa3ikWi9W7tAD0QwE9eikkG
Ih/jjkGFUwm6wdf/Oz2SWvL5dp0rfzEaI4TrQYHKNF3M3gBJm8dd+V2XAs026HyD
SwZ1imSQbUoymEYs7YQjxI9UP4jsnI+NQw6tZn1rmEiWlnEXewR1ASeh+VCsuMlT
G0nNwCkn0WOa3BXcE8v2irupkBGcrlhgU5QSyFmNaywXa3BqgrRgNhN5rb1JNNqV
z8hezWB0FUgkgvURVqTvJ7hCCHuBgfZ5uA4K9QMxmIY2XZobka2xanjSOesIk0bF
xtSO2Q9KNz7P6ZuILJrmYVJlf63oOgUY/o9Fnzj/IudCPH0mvhoTehQ+BY2iYvu3
33Q5S117clDDF5HFDrNEN84HfW4USFhVdocl/TItnBk5IdXjCft5hvsjAoGoo3v4
Fdr2kwjPmp++tDD6aVnjlEGCBql7J+yqDFnbms/VeHqjr0dtfyrfSlJxyFfQ58kk
upeI7RTSQaSTeFxyXsEIBJ9T02NwRgCuIx7FUUqXUsLK9IQpABV95+gc/lIPNgEs
AZJrAXL06QoFwhCgCs0kf9TaO101e6eTOE8Ha5B85NZWAKTOUwgQO77oo4u71bXc
rB3zPeiw+PGGUPEWWc5LOJg44aLB0VbVqGcrFrNF0gHYhjAhDxZsac1DRyJRIuXT
fe4Pu56ofd1ECMYQpRqrvxfU8Sm/CxYPiQ972Yz81nk07KMcb1Cw6buutRgsqZ+B
W+YRbwk7zNCzzDSXWblJXdLHsFhCuNwKULGAIiLHvWPYDUwHTLpsLPn7aB9k7NwX
/FoVPxJCxQrh2FBpIrItTBReu7MyXVYhIc/wNLwexIkN1NYNL/6XoBdpl/doh4rn
kucsrl7jYPYe9tGAiw9BK7zHC0KpC3fWafUAEZvwpFeXjSNRtCdoyM6HXYNwOCn0
wRZ+949OIRa1iDqbS7OXZiQrIVMU/UMRAfV3/p/yVbAcalWKsidtcDHXINou7nCI
wF1cKZLxkpbqeOqTKkJZJdwBPafu+NoMV8qP7ZBRhMlITmoEmSm1qwdGp90dGIBN
vfZvzbYegVKEqAIKvPaFIxZvxS6uKSndsDiKgHRbU16lx+Cwdpd7KElAIKuzyZVZ
EyFGZ1NIsAkMhEXMqUJfXud3QGmt9BfBfWTj2np2Bp2/yHGPMG31+RaokbF+pZYo
VRJTDNYsfqxAzq02ugghJ5tcBijDQBCeL090N8xh8Llr/N9ceEYlcFnvqGCc6L2K
Gw+RM4kwMZcZaFBTjkZ4WZp82XFu6AaK9ovI0WFGIbhJ8U0HSG6zmHM1IDVqRdVK
Z+DIMKSIKCg04M2HzCPlwBdSPCJDI7FZQwn8qG5QIh7FqtpEQpXSnfRvnZWDAROu
1iaDnoZzyB7PLd2LKhqBt/0G3t0l13KkDvgd54jaIa5DtLCPWC0H/uKbbdxSZwS6
+hQabgaRSgK/4ds7brT4T1wCltVN5U66TEEWgxm2BpJxNRKDep/KyavlO7Mn64ps
L2RYUFHuEKIhstl4ifgLpq+131lMx2q7sBhoSgzbeMplc8EKPz9bpHDUh/VE9nhe
Di+ya0KmQWsmecViPTfTKZ8oAz6p7Gs5hAR5/sDxrXuOyqrM/URI+wh8RmyerkyK
AqydjFGExJrQuod0BWvPKLIZ3GE8UeQUQ/K/GvbSBoZ3e+ODAMeCNBxTn9IbZBQt
M+wujxsQQH+IdnBnDTBBQF+q5VXM3DMtLH8cgpCJyb88yvyUUBez9jArw2S44Deh
VXM1/V6IhrHutWpnpJta8iEV3wHXPVN0pHAlsPeYaEsWbZYS/6Qd2kqxqpjOYrlR
Ej/w4FKzpFf/Piy/CY8XxUkstGoHw2gwo72ImpWFQPzy5fFP8O6tir4ccUIoyT2s
AwtmcQHxxUqUgJumUMO8rVa4TSfmHsT22EYF4PtwGE4c5bs3J0wuGIYyfyPQwpvG
YGaTTl8tqRUknT/MQof2oHI3/BW/INY/EVPKXYXhUrNzSHpTWDoSsuNrCInA++9C
2BAuMyGBBHW4cb8h6UXgnd1ZZAW3RKQDy2neU9GbKEIYYnYwrNlJ9IQ0J9KH3wmk
ec8/GGsJWozKURMgNVREdEiWZ0JXLYjGpO9CEn/l8L7FcFw2DWR+Jktq26RA9mx7
HAaJBYnFbuAF4qbmnWqkO2iZY+rHSwlbJahDkjJ8CgiEU0WagNhAY7J7SBahQ7K2
H0Sz6atjSwWIWJ84tJo+JtmMLt8j9jC6C7POpcdq/aeO1RCDTsqB1tN5gU/Uzgt8
8ny5+FTrU4zSyHMBcL7xJggX1MC60vvmHV1OAapQFjAOpIRMyVPGHDZSvH5JphPq
1OlcDInlcFZg9zY32YJ6Ho1sX/3b1W+4SnPqNvgWCpq/weAFuwn/KEc+8BiUp9z0
IDdMh5N0ZXscNA7H4RdxuC9jsiUeQwPGQjquMdx6//57+0tW2eE9JZ1obefj361J
L/FkDdbArRL/aCk9wpwN6tJ+S1nncVkSqgER/peQSA13H4NfNByjwMoUGEdcaGJ7
OyfQ/a9CHIGen5cnRVgd0UvqjCK+fqTpF6NBJL71pW6xHiMQwro1+9wwRsE8PzO2
9DupKlq/5GvGDpIro3aDj/Sd6NoGb/yg9OMfK0sjHXZSWHX1KB5l4i0rqKnVdoI3
hwbDhVy8R2b8Ny6HTlbl2hKeF2S/WSwx/rqWL9sDrQ2hHXkDzMD8RUG+qaayCJsJ
6762ondb4eoYgf4eEA9DVZD6zOOkSw92E8u897utwbuerxZ6Z6qmSwBL2b86Y3m/
BwMzkHQ98k2hPN9Ham4WgnjVqiWYli2CZj+qSS/rfG6g1lacXanHJy652aDpuX3d
tjx5ShKKslZgwbDflHfLDylOhUdePFEWb7KIWnByva/F2w4SAdf1/nUM2cNTcbLh
TkcZ2Z517rTtc8jSNBe3JNVSyA+hUR/mLemV0f2DaoC95ePL84U91OpZBK/Vwlhj
pyZK6aunj6KlyYf/jQW1zo2IAPi9zo+TNzuJQ91UKL/TbEh4O5LBtSogouslwGfK
NiLeAbCXSJPDXtXWkHqeazQj4jIgbWBjy7ndjSlN0P1RmTlTCFLelioGQRQbMo6v
Zd5dXji8Lz4LEWhm0WmEJ1eTNILIwvXMldjocTTxcF3CzAfF2xuHsbTGw1Pim9aW
PUv8RRY1nKeuteadRFfi8JQsHHhQG1YlsYT3N9Lqp4PmEBactul9c1FQyHFFIAf9
pLCpi9XibYythvGWMp+Ycx7Duhe49zlLDQG1d/Ttj3g=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
KqSDpq6t8dH0Ol90QORVXsT6xVmMgZyHd3Aq/9AToCF92+AcAmmihEiMv1Uwj7+D
149W73X+V/8QbRZnQilTDOKbSHQhI0rpxhkJGL3SgP63RPNEpQHUBsNYCxoSkBo5
HlUylfsyTzwXkByKGn/Vt6CV6xpoK+3EmU8OVnGB5SuRC+qtN53d/EJ1gvAbNNJM
eJVB/6A6Fx1b4b+3JpYE3qOFz+gaVlxsWC5xGuw2uRsuGCUcIflnAAIO08xSBD/1
TDuE0vdT3Z4ciNb97C2UU5T+AfRXFTMISfxN5EdCPxDtwNyEoPzYbiEetZYLOU3p
6IhL6em8EbtS8++caQ5jOA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9232 )
`pragma protect data_block
1jY05u102hgW6bqGjkGU8RXNa2F/oIaWvK6y92dnGZOcrBy1vu97HCyrCxrA05qE
kQwhsGQJk6Bw3VweTQSNlqXaG3Dpj5xKETRA7DvjdSAg8MNqfDF4vqWq4xfiuQTu
TkF9Jr4wXTbIyvAGrAylEZwI/wuIvvv5K+JDE9Bps7CEeEiYfcaaKKlvebel1koP
0m80l8woLhWpfOewVKqoj68QiKAhy1QNF71kkOS6VYHdhHH/b888Ixp3IRnA+mWa
2JpONN4E9/nOpiK0gJe+3oXgCVvzK/jc4lgBHqp7RQZvbpHD/q2ot+b4Od+LEFTV
YnzBvetUUcunVauCczyMm/PlNO5Av/3Rz8cm/lL3ZB9ecSKe3XlIvPXXwK+fNNSS
XKavCsIN7u4ee5tCrbuMiz38B5jxZXRavtBNOnIwnbRyRgp/y3nVO5jOJ+gHTpqI
Olj/95oiHHOF9pVtDg3nD7V1fySAAYGeLi+cQXbgJ1TgfHxh6LrEwqkL2rrEXVOH
iE20ioKA/KH6CGSl4Z9jdX3H8u/8jJDoSAUYXs/5vPG0/FRzjobEYNxfRKh9Dy4C
eCk8yVfJNOpjVGnaMV0jKRf0x/61EAJDUgR4RLiZz3Yx+f6GI+wcNCvo/XJ0oKaV
7I1l4u8Hjs7hzv9IfFA1h1Zv8HYwGt3cN+0jwr7oIRtuhESO1y70RUKTDG2j+ek9
J19/ymNsxighQWeUyig5pSp+oD02Et9sLiiKQl/KhUeaeG1zndK6o9Lbc8F1mI2Q
ALokU1RYyBLlV0qD3A70zidfLFUQz4nkj0UwCoo6EpxNCAo2QAEuH+GF+AFiR5VI
RQs/pC5+I6v5xLwQLlfiEfUIt7iwL4ZghXnNC+k+s88JVPg4L23OmLS8K3dJufmM
acg/j+QzVcGbKctpSWIBk7b5/HqYBhmR8fgiRJyP9gJGw65sldDdFxp+YF+dkxN1
qlYxaGmwEn31i5mF4joJHrfmAtY7dOcZdM5xinPUDa7r+/whq9nPLL6Fpknmfdz7
EBNcM3BkebDOxuLCBTq66YLjVW7xdUCdaCbzJUmkBx9cJI+fZPP471QQOiYr1pf/
cpj4O5o+UQ0bWsWig2JoOSsUOck9oHqlW13IFpRbZjSEzzZQ1PPrpSG7jNjZ8102
dmTBeg7CbLayfAqX4aTeHh4u/n1BFaMiej4RV6XqQLNh+uJn/x/AjbdH/gv4RWxY
BlEg2S9o7N0wANB8Xy9XG16An7LU+lwxVSC319wBOLc+3/EHMlwHzIwGjDQOJUO/
tnMCaSg5tiuwhAnwf+5T3B3xyACUixpqw1fLpuNvZxvM6DYyFXr32UmYSfmN67C3
8T989jKY8InBoEMZnoXGri1jGpwSYnsoeTcjINnp0oQLigd02KqP1wkarpoNhTaR
Pjb2Srzuc0HY/9/PaLc3h/NUyb47QA66liW9PTUnrk1ABMSvFm9NvT2ta8surkc/
vQwaIH0wQ7/EL7udHA5k121dOICOf3J81PmH19Xfcz6M2Mg02CkDJTOfYooa5IHl
eJXpIKXJBBvS3DVYHO7oFOBBb03n4SIEmal4HczyST0YCyyvlt62I+Es1wVOi3mY
ul8zq67mfhdzwO0ktKjuBoIyQqkQIpiay0w2EyrbDpsO42AaVH34LNkgQ83Tpywm
rq7/CHRx4oc7aKx+RosFPfyPNq7NxC+vEftVHUSstIYlc+8BdiEw02q69+w0Zqah
onbxqOhjEW25Em2Xh7+rwYBsEYrtLfqqn5B0gMb6Ig2tb0GWJxSr2l46BwdS1HoI
8FQkzkLji1O+agqt7R7Q/3nbNpcAJfLpyUse5L5nv6x4FlAwqCXivRcV4IfUYNXA
viUCXWsKZfvfbIqLfHLeKr76gHnNJV9m7UZ3ZB9/NZ7puhXgyTu7u2TyUO+JwNSd
Ky+4duBN0lJSukFnSwJhbs4aPfcRMEtQmMtB/yhLu/1+AGIPBgagIr9BGRoVlNee
uF8X2NF7MIoKjhR1Tv4waMtBBohPLUv/iTpztp3tYeaFetAsay9zeEORVeNaTQ6k
Wsp8RYAvMUtvTYnUNLUOVL8QG0+j90dRUFc32FvpKj1kqUWdn34nlLJmaSXJrQeT
5lzEAyokpJzLP5+42L5RIsL0VnjokWnK67LTEiR9v8vdZeuB7/Uzjr0aYPYS3v1y
xXOGGMDJpYmZGxKDSgcg2WYYUueAZAjm1gS2Xsq46vmAxroDb51VKDCi0FNrqN0f
UhEvVJghV3rxkJQT8syaqdIYp6ZggZZ3D9yGJCXVpa4Ta4divZyfF1gCRezW6lp1
VCrhXXGgB5VUyZpLqT62OyOB9FIwBOTb//E+EWZbqieTWGz4KZ1hE1aLR8Mbo33T
M4NhyOO049G9fmqaarf3ZOnHt/wTIXsf6HUcfvNzrigX4373Rown/1nA354EQv5+
it3kvJg1xjdQn8cc/jYJDSu0mLQcVHHwz+JyofreTiJJuznT4+hdRdh0b1RG6Ah5
OBP2xPFHhNLd9asaXwvXAj9NTxpD1vEcoTaeKOkTnoomBtBhgYitGm+RoS5/Ws04
6Og3uqh8eNX6xY8XqvAypLfE0eeOznC1TTH6xwgcms+4farWX5WhtRs9ID9XYZHL
dfwI6TW5HBy3ct9Xz2nfOZez4r2+A1qz2+svXVkwA1zgky/G5F7GAVo1RNHQ3kuH
/T6m9vZMyS9qtlbpzGa7SbRRz4pfH/mA6Q59yPH3IjVZKblMKcOTgXFXbCc8+Sat
aBgr5LwbIVipDFgkpjNTd7qwMJKgnSPhEG+P9/dGHot+2H2mS4/4eQUnRZzhmbxX
y2tIKKanKkUyptW8xQhlvpSVlIo8ibIwwWhSGAoZhA2zAnrl+QVKMyOaNQYmeF92
cRnI9O9IiKqW8j+gjPurQX8tY8FEzuGx49g5yDvVp9NxxQg5qSGO31W3XhaQPRBI
YYYyVcumUiWDJuhBNhiH86D6beKLHYDOWbSixHvtJyNFTEO3bxzJERkS6QZBvsTp
J92tIvWusczPZpLlioliG6OsMadnI9iCfYSIA9/yvy9PZpHoIgic+zUe+pXF6Ss6
Auf3VKDoG2qmPxDZyvclV0LTHZsaDyVZGKNeCFqL03sjtNXl+t3Cd+ttfIZcnkvt
EaX90vo8DEuLxaNDQgiIgqinDSoOsyNWOkFYEXFvnvXKrpLLp9yX5xRYi2k23ZwG
PLBB4d4Dnza7odGj4VmD7aHSRRsmgV/5bdKVgM1aqKdMgxx6QMhGeR/6HHHXbW7a
WRugatTtMllMbYKczta2HfxvK7CJjqQPOy3DOuzd5U9YdajPTLFHYTtakElNXx6K
KzQHZdXpgMb3y+QyE8GY3sGI/QTyZ447F9a7r3Ri4Rs/IrJjmBD2zLz3/ldUaNWe
C/r5yOF0SkFRftivn42PbszFZzvMv8cdELMnFR5cc259r4xuKJhXW84v7HABuv4e
pSzKxHG2YUmE+hxWNAUEXA2hNeOUHAQWhFT4YQk7S6M6xNHoTXaDJGuuHBVpPGhB
l/pxdCVhf7qGJQF+H3f/mKR58RIZEKPVqqMcF/XwOmr5Bv+BC3+UEumSCg5zS7eo
xkmh+hugGpoWyRNr7F4K6hl6hrIneJ60FtnjxUyCtcCRdCMFmQdW2ir+CA75NEL5
XDdTM2ixXzteBtlK4Pp7mmrRs47HMFPJb9Kud4UCJkkP2War3Q2g5Kj5HHi8dCO+
bPrQoqEBBNeXnpfsNivJLGnNlPFd2ko+bYkS+D+3erFyxwggSzaB6KyZZ/UD6Pet
su9FASeh1Ol4HRpOvB+TgrGv/vYx9p3DxrhI/aCMWlUOHLT6SU7c/XEByd/qoKu/
k+CcxxyU+4P/cbMQ1Fgx8K9Vtjg1al6XLm1x0G+NitCVITHGy1Z4keuMURVoQVh4
go13IVbg3UciA2LRXwPOj6Czy2B3W5hDisBw61GnoM429GvAOXHgfQA6ZIABRSht
CNXZZzja5QEsZFL/xqhLJv3icBp1dGVOGBNtmcojzaNDKa8mR86tPo9ALugsZ/5q
A0yXJMcfNw4X7VouXbg5CdC529/fyU+CpGS2rD04+I1zgZD8zLiCtIMbGcEmHzER
8nnm5A9ZhixPu9SENVlD5NxbM0pdESOxpeYQU7+1JCbAC7TZQi2LNDN4aIaVQcpl
J3POzsNpIUMOF6uBKV/UMcXMtqOefws/r/PxhDA6x/Wx2w7qT4ok1JeDo4jwg7eK
2OILuH0Nk/2KnpZqmgTkbsjScqRXXWLlkaWEsje0sEnXHDf91D5MUTmzIBDA9l/N
sga89wLJ++QdBosPzuL44vd5iJr/8spk5FERlX3Xnyn0XIlZ6LsvllFg2F5bkA+c
eZHBNi0/6vzL5OptVI/qTRXt79TXDccndHEIBT7gjG5U41fGOUMqBfSU7Jj17O2O
NLpClddVMYhlX76UzLShe9WlHIsJSFprTJr6CU+YZ7ku/IWAE7WJAUvm6SL9BPml
WOWDPllq/CAyY83DaWr6lzZ4cpGnI/hv9/TsEiuxZ82FiquH99iCIlgxXX/WJwal
iaKX3NPQ9tCXjZL+U4kKENL/bFcdrtXuX4pZY9/8NqT5eeRccnibYeqW5eUK1lYB
tQZNle45qF2rKmCfOYYaIivJY2Ug/P1pocdFYf0HFePaDbYt1l08FV61odSWsM3K
1OjcNlMYyJ9z7A4qN30MxWVZmMAoEGEIRRuKk/uNcFowKYuEUzxpjjVEdmZ9P8Pd
4gcWrE6/U+KNw4gS4TDav9HcXyYVHLUEkXMN+JwDiuKodkIBvvFHf+7az+kw65St
u75KW3dAeNuh2v22j4Sxrf+tYoCe/svAidslcx1tA5GcrUkLJAtEAGNo71JFeLZT
4M+2f5COIF04d/VU8Qpjka/ySds9qY/MmXPYNIzU4vTt1XVKKXRwdObtbgwCyLXl
k8bXd6alnfxiIXOoIxGlTNUPm+8ieuJBKyw4Zq+L/E++4ojb0toI4YUl6CE99Lrj
3g5sfqk5CpCemlmdlVyF8zuQnuwiYxv57AQEbrMHDHUbG1TZLZ9bLFfgFQqf+949
tcdMQ4/ZFgySro/K2KqZ5PAlwObTNfK3DKwQWlo2mO1Wm6f5hxzdbykmIXzpjWcr
rXraPzLhNc8jy/L2BJkCufmCUQyzYEemX7oFggAGscZKzieS239FhMmAtr4CZePh
iUT5Au9Lk9RVc3QqJL6qWBNWL9szwR2P1qa5SqUQUA2KvW9jh9GTGFSCQ1myPziz
pECAexKx1uf2yH9t6QQCN4B5m4+wNnHjhgDRKAy3PYPv8JT4ErrBn8zOT/e4dhbc
PU/KRrQF48a1jS6gqgc8tL31UWX9kMD02tQ6mlJ2kKOe0Sbjaep9VHEZ0HdS+Zsl
6NJ543nR39nWHYg2nLnSRUQD4mrtJ0pcuQw/XcXKhkDp5gpF4C/WCbACq7vPeCkf
8DF11O+y1Of9i7ZIgMsARNwxik06V/t1qiV8YpDrpb3mBNkf/a4DqFrrRdN3lR2t
pdwd5JktwjNmRjjOb086Py7jBs1cgF+mVUvsMYhydIarknGrfVfMUkjDEkeQo1Bp
j20+rdDtTIx4yAR63aQdF4id282nD7THGRl8yyMVM3Lyg37baouODDwQlvnPU6wc
9sUZxJd1QRwyvD+t5e3DHQhPCVXysY9StqmTOkfRxeeZ23dMYoD+msZpz54Ex7XZ
7YI3wT2va9dbk3hjHu9zFhM7+B6ZO7rtXrBtvU2Rg/VI+KBbZsskSjnTcmM04HQJ
OqGFbd+kDeNEYIWqYIgBzk2DLiWwxf8AjzJqX0lx3V1Vg7RexcuN+J3aPvAaqmkC
7lkjz8oB9964sRZJO0RzIJyxRBzPYnNFpRpQINwm1fq4AACHtpv4bXlHE8PfdH4S
Njou34skR6KkdDOgX2njtg4Jt/hQCpr2vWfpjTRP515R/9ClFcn0jLlQNTTkF09m
saXAzasLsd4XNHSvQJ0IFAuwH2l+jNLPAt79XpC0sdCPkJaynfSTS4sAGZcxI9sm
bk71oNaOck2q8Gec/TmrNoW5KAFJdFneJZ5El18kLEY4FKflKMjeKSq+Al2F5d8S
NY6Uq0E5FatOMEiiwffWuia9onf5l7vtNziP79/Pw6ezEWkwbrzyXYF4j7TwgZaf
wSx5Dct68VPnvyWkwHe+OyJwDXEKyou+3Sa48wOPXJxdnWicaYf8aQYKEiiA2sh2
j6ly6I0P0+s31B/Yf9yu1yVozRniXrM5l0qrHihkiFv3ZCi+cSFgQ/lT5wF9ZbW8
7S8o554AclEQ1o54Fxu4hRW+VcRA3WP2zKWgdEB6k5/dIUCRQSbuG8w71CVyVTXL
c9mvP8JMhNM936e2BFWwOgH0V0gQaET9xKIaX73NFTZTlXHmVC9kWotImXGulsV8
w6EXJZZ19QWuHs+M72t0r/X2m29hbVSbXPiDXnD7AWecJVSY/SBw+WgLrrN19dKh
FgRS6SIyMqnrrtOVNEEwZ4YRb+0NLus49exsdalP03HAxwe/kAvRqDvRfUpkyflT
+0juCd59wZASnvPR8P/KiVX5lNfK3JqptA1ZaAgmnKFFAixWtk7Rt1xVx1DSORdD
t79zceFqzR/PhZ4Dvp01UjeTIYRDu7RhNU/psk88NkiFVXITmyyW3lZXT14nvH0c
aA7ET7SLtzKvY+2n/9W2RhKBei4umALW1bEbD54FjnnOfbEk4BP4ZtlUoX5tZHnT
VFDiPWIRb9U/vs8AVbydatHXvhIE0nlz+UNRbxaGkBW+i2egQWDLOcAlcgcwKxq8
lKGHPi/7cBrQdtP7/f6tKa4ObaJfWwG0TI8nW3oRi1Jk+ivSCC5XniSZxi+JnJ91
uZ3Px/0lEuDnvl8+h2F9uWDis4ryXgr25o8swUTvt6trXYTn5DxYMEkGZG39G1qK
r+aMUrgaS3nYznovDYZjVOjJAU+fcNxOPU9u90Ct5oc0dkMOVcZeGeS/AVp7/BI4
WSRkDRvHoozzOatc1QfX9T/pGI/T2Naj++dZlqKQwVvcHcrFNpNUSw0+pB1WSw2E
OGPgkKZpqtmpZtU6HZycfVNFIeKbNEJD7yXeE/aoFoGfd2cvx59dAohRVGKO7wCr
xf5tIxpKc7AOa1+6jKSkWpk8mJF4JXIS7mfesikJpLxBSIJ63Ye3tYZyn2BKm+pj
Hr/K9oAfNqmHiJiYj6PeuKzP1xfEjdMJcdJ9s2OBQs1ylJ7UMILyD940soGNjIdT
P45yWDOa6mVlodAsukWttcHPlzLo1nFj4FOKNWd3rUSBGJtZGIBztKbD3qWgkTGZ
BKXL7YZ2wf1gX7XBe+6nd8JGQbPdv5/Ck7esycCYVJ+JgGfI2/vei9Jd9Y9Bz87j
BfHuEQS21aowkikmsRILk0lqFOq8nmXw8OjhiHNOUs9zWEGJHIAWHBCzEf5o73hT
aHIsYl9pME5R9zMdyfNPDVviWhZiQPs4W5w7jFVkaZIIWhMGcCeL5qOCgPzzWw/U
Jyh8bTLdi3dFj7KHW9WJC8ZkTVTYOh+fvOlekAyqPPVrMPjbLEucZ9PKWf+uxRR2
7ZAQNNQUktI3tMsn7IRIIHiovwzjlUoMbG6Wo2fvxDpRDQxPyVOxfkKMBTFy3eF+
d49C8+Ve3ky40CGzvDJeX5F9MS/v5rZHrFz36fT3Xvozzlhsx7Zaoe7ZuT+/LajZ
Fa31uE5zbvw+DOO0B6w45FJqi0UDSABuWDUICbheD7zway825q78Q/iUPqcPXgal
3P6DRP05TxOXOYdF0lyUfjjepvHpZdatm3tdPQYago7WGbdT1OvntkqGSPGzLsTC
Y9BnoEKVG8mIGYw0HXINdMpzoYeETQJyoU/pwesRd6C+ckIF8SeLTKN+ozgNxxBc
wK5zucIwCr1ctjftM+HzNDL6XtV9RKuOzeYZpAVivcj/l74d37VacViEo06nEsz/
LFrlBPDxgqUL48MAOkD4q1qa3zXc8wWhKGS7U/qZammFyXoej2afecKGZLz/4JeC
kbuuwt822JvprSNHLnC5oXd+lk7XgmNscBMytemnrhmjSzXoLO00JNai8bVO4TET
Jorvf/hqQLHv70wm+uFJ50q8jCUbpks8gXW+Cs6jngbytPYrHBvCpet4Z7+Ti6Bh
dSwEyhl3ctMmFTQqz8JM2zh/nO0Ds+rS/JIIAxBKFhpaVvIqhH2TDYGUoXn4lBue
1SWEoKmSr1mQiVgn+Eb0lxHLNW5fJX0bm5PpUDRrhOx9a0E/iGcJz5KKaNAztbVo
W4ocYaIKhZ0qquhHnQmHxS6Eq109vxtzywRsF8zahUUsoM9ut/l2nHfL0Y1XBr7k
wcWQLgwpaNKpsc32Dsp7igJfU8XkVir3TsDt+1ze8qRTOjncP70DCEQ1zW7f772D
y3w9fH7xh1FBvMiDniM+PSSD5eoKVp2l4F1l3upLzhgYPwDtemwWHHA/mEnPsf4v
w57pgTlR63p8Z8Kddt6C5PC4nDYScv53BHujLM6wX5lfUgaSY/3oOfuyqaLjLMeb
UQEpn7pDIZP2Gd050lMe7S3n8nzQi+VpYhw0tiIuW1b+k/vOJt0mbSn6aiHhjg1a
f5en/Wu3YiuyTESV8bK2p1djSfXq6ADt1bTxccKRF5VWzujLZ8mOlO9AUh6U+iMQ
95cXRZD+qpEpDsb2a/DR2CUwxwy9dFyVE3cIj2xevzLYQ8EBB+DMKFKhLQ+Fi1ZK
Ziyit1NygaLdCl55Ornv2FFMsUU0qlqTgYPW50qMxw6VOQxikrh+WDfKPs5MrzfP
pZaExZsbDB22Pzw6N1SxZuxLgKBQLgLBYObm7NHA7OP7b0jko4xM01L8gKx/ECBq
Uqbz2TVdDSlh3ZrFeiy/9gtEq1DRckw1RRhfbasCj61z26O6EIoJAifJvKTNACuj
UmvdBHNcvw3LMh4pzIuVJ2DKsSIEAxTQm+ZF3kl7N2gLnKuCtPyd4RjyvioEe6G/
w2Day5/X0ABjIBJ/fww/EHKmm5hadtbURLfbwq6kMcRx7QuaYQlqiqmbKlimHU3O
uJKt9wA8CSvxUD8tb6CHxrbSr+v73skn7Q6E5z2oYYY49AAZ4AYtYkU8Gmbo4Zf5
a96P0LMySpJYvZcXO9YUPv/k2BZbbum8R04aOmyYbZZ20os5WZ3wMY9BwwYi2Sz2
Ts0T92pCGqnDqpZb2p9v3HsjZ39RVwBkuqZhrSwRenasEd38cUaRCjjB/9ldIm9P
Vbu452PyJaU/cv2Af+hJtfp416oWbys7T6Gv5CRJhXws4HxamcX1M5F+x6EM+JZ6
vVg0HpbOT+X7HwBHt4UUVFowovzfs2eZqvlRTm1/Um12zLYDhMtI8rxEzMnAYpIk
V0xsVi+k++j89G0pO/Ke9XzuOIKjFHGydMx1bLImxRE/+6nmiHuEm1rAsJStK40d
cmwGMerOdZP7ADVoGeWgGc6/0DijjIaGYMPAwoZT7U3ACfPCngutimUduzURsQct
4EnN6PxCq3fr1CAhSq5RK1347p554ySnku+/WwUKchDz4T3sBKQCPZGqW4WZcFh8
m7i3760lO8WuPYW/du7qS7xWFwWzxZV4AlzgzwYpj3+Iva6l74ATvyraUyFN01xK
dU+tJN1HOfDULrZ4O14JAVkz3TOkqahqPRGGXyjmQLkAgmUo/J86O0o5jg9XwD8j
S0Dq0TSIATWGoKFBg4/dZv/z9jek6wXJSy6LfqdkXILLf4rBQq09IUJs91WXFX2S
0nhou0u9FOF5AAQbrJ3ByaOpgYuqIJn2Xk/zbQriXtxbanyWz4yQEc2izx/Tughc
o7IVSTScWG0xRD4vgDZP9/9QL+2qBAkhjkDpjh8Se/+IIOOp5AKWJI6H7Q2Wek8R
uqTu39rD82I4Fe8eua555nTF9tgX6Ad966fJ0/EpYch+PmgI/LFTs4rVBxwjkvOp
JRrrLx1Bn41zDQkE2yFNen3gqbiRG/rWEf0Gba2R7v7OO5fKcK1KfRFnKsiyok4R
jT+Ny54gvadN2awfz+Y4ZEhhq4bjSsvrKxmMf+2WmHEEjxKYwanDFoqFiA2SDU0q
pYnL2h/8+bMcwXohz8zPtQC/9sdFLJkPueeo/+oP+Jf6ebO7VmCvrAq0KbFAVd8l
HUFQfEh4+jnhVWdIYQaJc8Ww7MmeDRP9CUaIjWRIw9SyZUDzf4ur6q1NzX9ZsKn0
DISD0bEnICxtK430Jdioak5GkzKIFdC/it62OEthnu+FwSMHWlzBehnq/xiksFxj
1tjLPC1+TofK4Ud8PyZIHyRFHbru63ccGsHnrh85nRVRz3ZHjTENCSzfGnUsRgON
RVVPU5J2lOm4fhv1IbhQJhE3JRs5HuoVENneiqkEvb7AmGxw9/NxUGzwGMOYVi4y
IT59Z7xjdYnO17awP1TWYArRcASb7iYbPMtLj+n1SJZtZ32xjzqongv9PrFA8+F+
PVFW89Bl3IyVFQVGrUBU0GSADUeoyfb7fHRaJanSD/P4+U+BEvwRNcG+3th6a6H4
5tyOylWVscFU1OEIpN5Av9jupXm3N+7q3luyvCbAEE/fe+mx1u61ArVst0mjXHs/
5Nfs84bxxAzJTAfQ3WVDf+lPBTrc49ZTT1RqdTLh7tkz/uuUvsNDimUMcGGbg4qk
0Hl8LsDEMHorFKYJxMkzw39lhhsDWkU5VWo4FCY17p2R4CIdBaKRm65L5fRVsGZp
UuoSidPjsimZ4cIi9wDuiwem2Qihw2UYsX3bde+ZR6Koj02MM8pRMzzSzAa904b1
4AxI9+VHZHgYBLH9/+1X3FOz+266uz7HMrX0JSkYPRf0uX4TmSBX4DQFuHE8CwWq
aw0KsV/mI46Axn+3NYIZzm0pW7QPIJr9MMJc6RonsM8VS0Ih+9+yNvOaja9D2xJZ
Sul9RMyqvnNHxz0MGs3fbl8WDTQJgaHAmPvUwIRhmdYTYR5lww9gNE+rgiESehva
Nx+nMKjhORFqcN7fM5Knz2h63EptqlCfZFJHzHbGU/pzrapGApSTV+ABONAvFvCU
zUA94VlnUEe8IfECAKC/ry+hSmu69UQ1Y/2nEEobrW+sCL1t2JTVWmSE6luWkMwP
n4ucryROo57pBIpiuzvVH2shEoP4NXwtVjhkaIPEKP35/oUxSY40eampWAElEADF
zRsTfQ0LaEG6EC3tfMoJJMAdAsH2pOtantM328t0+Ve6Q8EgtjwSnRmQfRhIiCvC
V0RPIAZOCZjldIyw5JkHL+yszM4x8kz2JOnVlTmDNtQAbmZ0j5jNO3Qei0p9k2ay
dd1G3vcTJThRY+I4OzWAq35m37fkr/sMUN9yRyKoJa2Xe1sNpoSQlxvI5M5rUnKe
DHs9NGEqDSZZ1VRzp2RZQg47kIOrr3F1QL64whZms0s8Eh1TkVducmHx8g/owY4t
/0q5g0gf8QLV20wEUMn97xOuk2ZFWxYdpNNtGph2POEh77JWXqVrIH1LRV7D1VUy
sZjayTn3dJcpM7BjcqHAhMduKhHyYbWxrq+YxeH3ySi1uBTzAED6GZHRmI1P9zRT
fJ9BdPG8AQNzq+IVzTD0DSWLXV2aq8D7w6yg4PQuGH4ngM4nh3sadPaNC40nCxEC
KJCMbSP1PQ5k4bVE8CdMlDZwPLAFRd3PqdBZ35YqKnwMjQ6d+SmhQylIVPMoxenz
LNjW6auOiO1eT1Xnlh+Z3TkRms4ZIKGpbQUdcU7ymmvSq/Vj4cZy08tMYlN397Wm
ME4xIzGXDga4OwGbvW8X+jd+exTsNA2cslY7UguNMcwlz/Ux2JSFGKzdh5Uu4ulL
OgIzFVma/FGkZMIfkuMwPujVmHsKHOaaMsexFb+5cLKANUQgpV/OlFD1FNwuPUQ4
wUWR7NOn2SBGsmhK8YSX8MzJgixUxcKsELdXYBw9Yq/NpfwEZEkLtCbEhrNoAfEN
qt3pfGjxyYcyleqeeDbNsjjmDRZgho/NaUWuYIIBhtG3J3MCvNxMm5n2ZpVnvLRU
KLeLXpUhIho4YFMKlmVDYt5l1PIsaGKHaKfkSzSpqfq6BrC79asLeLcRTZ84rulB
ZxXrSY8N9DxLT83n8yyPcG2/3+Jop6eaDy1E6TbkjD6nyTpj56PPuZHH61IvDut1
Wy630RJOKnruG9nRdZfirTs0hXR3OCIQSUfp1gEBwXI3D7nxmqAqMFfyCFEjv1I/
QaaJyqR0jrv8k1Yr2TNrnuF4s5xjMtrX91U2a6pWFgjV4aMeErTz/kzPn3STBCkj
MV2qMJezTYW+WGLpsRvPt4n5mJFj+Yz5AeHBO7MxV1MjxZ3N4Ydt6VaOPy0rVYP3
8u6qzJOVul9I9e18biBlOQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SGXEaJWRH3qzCpkwlrKK7RmPIccSp96VCiMSMsoH0tm2JtlC326XeVAa4AS2rZIN
I7sncOQyZ7z2cc3lpdvi1TJkfgwbJiq4rcUkFwDUhMEScKIn+76bYyxFSsmuhzXm
5YjucIpV3wJOQtW2t4K/ln+Mpa8n0QiJD59vVCWRs92iL2xmrW99PCK3hMKM9Ech
Yr9oZAgbAmZwdHwlUWCRy4HHea756mdWoxXZDXIP22zwTWh8xGfTrWpetdZTan+l
AugD7oKpGAEw9kN8iuNqcA83wvo99E09cXgkXk6HcoGWUlLuQfnQkFNWkbA3H2UW
Gq+srW1G6BqKDp7cGhkzkw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14640 )
`pragma protect data_block
a7E5aDENVnwpULUaiDnpROcgRL06+GwlFyT2eVVL/rXEo9iZOdRfmNW3WO9JPGHz
yTatdKXlmdi8n7bQ552c7dn5tw6TiFkovoNboKn2rG+uOJQT6KyXDOqF2+J94yZA
1hCcQl1QA9igEDGQttjGPLHs/Q2NjahBafzpdfnToy1jf3J3158PBO64mW2UEY1p
l+zi+431DOqgth6ie2pwOpg05+K8PKCilG4x+pa6oopNKwUNe97ktqvn2VInBGFq
cxsOJ7z5N2U7lmgt/8Uc0biKiBylq+fhXHywExeHIxPREhNMVv52Bte/GnGB8LGq
AtCwvwENrEpCfoRdCwy86f+mePZqydqq4NA/ZM4RggmDqXaKE/bxPBCcmEinoSgF
0t+X1GpaqQjR8B9iPHl5iHNXzA5TOmCtwF0OJFJrVPMiz5ph/JkjxKJz4PqB3rH6
0NC4nE1k2TLlB2wzdQrS/1no1jjrGzbxNL8EU3OPj9EqCNOcsESb68GzQ+nsVCoa
A/q+x986brJcq2AdD6S1rJlLOmG7OX2vAWtnLpXTey8b1/uFRtORjPZdXM4Jor40
nNeMJ8A4q5ZhkoAeVfAiO3pXk+TizYLNlrtpupCrBw8KYj5jXLPPZ1IXgCONnJOH
+/n9dclCuRVgULA65v248L93r5zW5l77nG6X8D9CiejtVxkVyrBMSZJ2GEStoyG3
fKcpOw0j8RThQFW81oyHIWUzsOsGkE4M6gUkUcu3r9rjv/SQUmagAoKGrTe4/uSr
C+g8ny2hL7kGqrOD+kgaaJsgFjIOmfLefPzW/QdjvEB5MtsQco/CXSHg2WVywANJ
E4qel+pGG8fdmktfvdj4vOBSCCRKeqFRYv6UotetlUiChIuI1Yx7Vho4/bZSsSNM
rwS3dAdZ7xY7I09pOXQeBI90ByYhjh3j1aYIko6hb1dVH98mLODupznNihvJ4EU5
dfrWb3PQOkkqX5PsFUZFKO52HL5y8hXclcg8lxkhCRoKUrN86fl9g2rx7hqwpTpN
fzW9jIrezSm2j6SpbyguPtqGmQ/WNgwyBMOlkCziynOt6EMQHMfP1M/N6CkSH16h
5GPc2w2NOkWGSB9izJI84iHMo5TSwMal50kZaknrV+qAwwqO1/ucxE+t/OlYmpLc
6JTlu9btBT6V4Z6PHbqqgtIqMHAzvqUB4zyTZB3TPofuIvqIAD7fLNCnbDY7pHrp
ck+v9d20Lukyzu77zSz7z61lBmlk+fkBghiA2hFg+ySqjGFIWOGc9g4xQFQu/Gor
ha8A60MOkZoaLWeUzE6N8XTQxAS0bDQAe0Nhta1fdnFbZY8XchtGWzvawbDbnPUc
XnxwuWKAggUQ77sClma9kdkfKcY6wCt6wlvocaUMSa9KLff96o6zCPlFazFCtcL/
3UmbdnlMrnG3iNi8yVPedTqHqHA/6SU5E8But8rv/XJsL9me7MDKL1dP2cPnKRQA
GwJLD7KKwUIfkzObA4gMqPF2GTuSSHcSp0QkRlW9z9J8G5q4enDHvMgEUgN3cKFS
KF/Y/LlyxJmxXsocqQ8z01qSmvClsu8bUco8jnvqjsIO3RtUQy/WGHe/JC3gDbWJ
ZzWLvy/Ix82ER7m6MOaclZa702u7QKejD0Klm/LFCI7fuNADZdatE4j+HEVt8X6h
mdFG+JoW/2reqQpqUdKPqAo6SwJmXtQ9y9eeaIx9wZ24QxnCI5NcEI8lypyvl9am
qWbK4RuOqEvP0MWwinuPGUrAj9f2/S/eV1lFOrnr+n/hk9R1C6T1TDqBh9StivSx
ecyhBKVvkja/3o8/IodvnEq9eC1LaIwVYIBO0wPWvomdAMcrs3jFu0ZFtiQCHLOW
tGXUXWADbLKg2DFhxQuN/c/IlnnDOtYEcw/F3EAdrLeqlgml1/Jkv6vPA5RoV9E/
ZxVjPqYOzlOagrtAUrIOMRt93Crs/Gca7Ybto18fMRg0E87T02ZQvFMac2ARYnAG
ZihG45yCnrYoy0apU0n5IrWS5FlvmY/Sq3Bu88esbGgUTyNv+tfFqm9MORx6nE0y
kqw/eJnb2ywpWAY6Vdz832KnhhWKkJ8ikUNlB5z+CNSplH8+Y8fN8XpYGFxDo9SP
QzsNqOelMXv4EUEY0Nzx2uJt66jiGEcSbhnHHcsaa6rq2asjfvfQi2AZmDYcX5/x
4ivyP85drIyCOiqA+CrFR9XIRrg2vZMPgDc8dt2eGzikRYiKJr1Uiz9P68tZgt0H
6RRg9O3HXl49ej6dgWtmIN+ixTX5VMkjlixoQIhREa+AyIXvbBeSRcf/S17ompp5
il1X0cgpJic30LIyQJu0oULQXLet7Z4+mV3ipEOr2Iuh1m8H9eOt+ZZpt4YYNNwW
dQqwPzhz4B5Nno04ZH994B2h8QGHrO+ypYmesUykSMK9HLY6f7/1HXzvr0omX8N7
qICaESlGmIDzD+A6cP2u6l65wbkHOExIix+PeiWQIf/pdBeOYRe6J+CmdtZf0rbX
OoEKPiLXHBXdpJG0MLnbq2LJ9Kb/f2VjjXhJz3OND3aX2IPIPrIXRubDKntu7env
fK+M99kUEkCo3kbCxBtML1Gt9p2JT+qfrR45CR6sym9O9Js6dc7zECYWFaHID2S1
PbG8dw/WjPIet2vBb/5FoppXKTm5b7FXnJsf9JPICrAz64dmIbpvBfwBI5U4hMoO
ofJOUQdhYjnjge/XUI+PweufaHezCrPtwIy45jqWyuI8TqcQZmk5Fz1SqyRjR0Oi
n4SucIbY3uUzgi9yjMRRQVOhAkdcqODwj1cdT9Mczw8opXdLHhjIGX/sFb5OS0tj
/Izo4BZRhB/QrlT7au946scYtrYI1UFbFpkbwDRDLgaMMBLA6gonDkyciCwzXSHa
1CNpbtl+IDNyF7bVhVc/sPNhRYobqaM3q90bzaVxYrGVeFvW17mud0Bm5289Rxkj
fbefeYD2+D8u5x5dD0gAnNAJNcgnIkEqr7Fx5i+BHluViIm0ImIrcMj1Z2d9h5Cq
eiMxVcOSvjzsF9BmFuwGUyDP2gXnPy55oufv/cFXBkSMVl3SgK8WW9FmNGNcq5fc
ZCi32FKLvw6fAIGFcYPaw8ahjMn+lw9pmz4fHMSOGXh5MBkqRU/WimB+83H369Xg
nUUf2eaaaaeImtCB+lpZiWgRHMGIBNdMYTKRhDJ8qI250DmRV2SK1ON8GqC7z3t5
4+fmntobkK86Q3TmEVJllI0f2Hh8+hQ3R0p1lpp83ozmrrFkdoaKLvXbJZPMtzx0
NG98zQTh8Uys5rn/SM/V1bS1ml/H5w2OciV+c674prCRyQE8j93eIWfDOg0rKZUG
AbtbRqKUzTfsLXrgnxbEhVlFIq0RgISdAG4Q00RB2ywDymnqsqPwJSz+6odEj/Za
B72PrmZw11VjSt4/ZVk5oZHnCubmAP9yu2J+N8+xVfapCufgwWRSzqVJ5i3eZ91y
OI9uxlc6oMkBqEALTm8ivSxqTtoo5XkWqCyQ2ENGGJdIvq7r1s3VqyuOuyocb7PW
1zAKaYmQS+yHCf9wYe8/26H1yKJpdxZP8iIisNJe7llnwBKks7fRvkrphg1Kpnvz
CjpV8KsIbI4hpacOD8s5AWUUSV2P8xU7mlWRb0OEtmS86vxv9Ln3CCn50nPGwbQH
inGxXCCZVMLCM98lC5oK8PRsqNryxVdCpxnVUXUfmvqSIshkY2p1I0+oFflzDG7E
+hOWhqfkCK5eCNHbD4ZFY0Yqn5THK+KbdrcaZXEmD/ySlSGD5ME/rjgOp/rTrSq6
M0gyCCGRHHE4Ap714cXORt3WArDu1jLghQv4Ks9575UxahQFiBOOrxdDZo2SsVXt
713FXy/Agfp7IkmAjwbE2dCixURmm+w29bkJYiMeUM2GGqTNT7lF3HX1sbFxzUPR
0YbRtXyu3JZOlsdqrAJwReXdf6B7no7OeCr+VRPODaqanf6OnK5vGkBEXYe4x3v3
PgcNumbMcaua1QpA/8QDlrzF+HCcZlUw+/SZBc6xnBGHxiBK0/oSCTvrpafDZxtc
/PdiCP8eVcfMT84XS5ygEm7+mEzrwCXG+D5f+4f4Ok8exjPYxPrNEtV20nGsZ0d3
vL0aLPKDabVd+4BkzkgFR24qD9KLQMBXfaV87Qzulcr0aEYMFlxm8/d4/X8CnNRJ
6ImQ91FTEP8l/XteP4yAvaQ/lGn8a2lkvsBUocxo1ZRncuwZ4Qoy1HTMgib4u86h
vPapaJqRCPa0kzRMh2GBXvmWNQoB/P//dQs0J/eLPGJ84Oy8VHY3FQZm7Dn/T9gf
Z079327r15xKHGMA2I1iq2Q/9Z6nYsMKXSYcN2ktt+Glb1PJX48Aqepn+/yM9u80
8YWBDmhghKOJze/OtfSNNPcMDoQfHMtfRiI5inm3BDKXMLEboNc7b9JdOaCb4u9i
v4vvo5z7EIxK6xkpcOJvMxWXx9fmYZWc2SbVxp6YqmGTSFAe4ZCHEHH/qV7c2Z3v
n4eb+JCz3mc8KC9DN4UAn8rb6Gtw6lNzCvKBknXbXucaopdMuCRD6rW5fgme6LUb
xlNaCswasHoeiRY3KKwuef7/0ZKaF9KcWlYeUSScLBwpwEPQ1N9Fgp4kafeKy+LR
VAdUWhosNV3NAuaZgHobCrMMPiHwNtTdz477HrOOqhzd5o2TKttzl1A86D7zm7Cd
z9o383mTlD/f8wQU0jg98QYxjipvAxCSRgw1NMK/TMPW75PCjccS081FqWLMxmDj
SbOSloro2UxG4XUO6QoUtVeJlXvF8ZaW8Rk7VbvPgWtK84KLE+NJs65aGr9MPebD
HY/wiUUr62UZGBWuL65SJfhlOrfA3zLODioiTA+Tt+yb29VcUV6OaeRC9ixc0a3P
wVlyO7J4X5bOslZ95ZZRlQV8HF6f8pQpVfySjbyMj5pjWXNA9IpxhzPfKpiMA6Y8
hqpgDbsVToEVexFNxahby+2VeRpx9ywNaxqptmcfsTCr3iers2sLTj3MbC7+jgjh
UtcPB2bsyrTQPlARv7mPPyfFnLjMCUqEOGI+VJRo0sEPyrnL/ZSxrBYY9lfYVASi
xMap8qYlPdFD8grVMB/2om8xzsvPcD7DMml35uPQbVXCXjHg6VH8CWJDB8gOm8xx
0NsoclufDmNtgtSPisVdivgcwKOkjmue86T1ZjoOR5tEw3lLb+eVTDGaKb6Y9stp
LndIh580+cJWZ+4zvDkMLTjousM1Us6KJ20+wz/GT2e2IZFzHuILHifnuXDOPFfM
C4lrNkzFl7tfpzwHfjiLRHnXv2LL+jFFyWQu3pstNlft/cBhfgWzSb00NYtjbFA3
udjVbmwZFqKQuojMH/MZXbZ6pN1fQLq9A3TX32XJ0Ob6xuzV8jPt41vJqIQl1tGl
XSFlOQwG1DDnuz8XLhFvYydH+fuYL9WRjPy0J2aHxqt3oJ16GVWCi/oVpr+yLXqa
Tti5AlLlPdXQV96ZvOzW0/eZWR6CBd5mxFc5s55QcqhDREf8iqbwFxsG/4Wp1snm
8igiNbXPa6FvRxd+4beHCNfth5zB4wxGe+1EaE82Gf6vQ9HOgU1R6QKEQaECs7h6
Ogr0khEpuOHBwASK5JAo57tTDOOw5xgAK/MwvpmMBfo6EXB0tq0BezIIJRdG/uqw
obHrHL+HksobmTAoWEI6o7rWtO1UZbU/jrLD3bxRBjvljzzqqs6UuJSuCkwigCWl
hlBXS+26cWL8dFsPFna1PHf0hgajq/LSZ5fv81VYYuMV5P8nwEGkQK3H2XF0PMUz
oh64tOEuj+xTvrGab37C8HxnbBNU+mzwwNZdtlJOUfQXxZA/6c0DOaSSWdw0NWyB
S/L4z6JinwCRVRaaAf5qJhbyEISVV5XB27d2QdzTQa7O8DzoOoWyFmPOKHG1v5TI
V1vZm5UdljyMTbZq1E0D5tCrfpGGpbQ+WAwMJEEqL+FdZPrYgzTjSfwfphsBiTGY
bezwy/cEhzYwiPtoTWaaxZf0Mk/xplKFaqgiNrc96MWjF9d5QkGVElw/WNU972c2
FRuHiLLdnS/BLGNHUQQM55G/9s5zg4C83u/8JddPN08YRgziL4laK0GOiJIWJ9gu
QNaKGkA/ZAT/WwofVnQr4fWQ7LgnmYEPyJ1jEAnpYVyDa2sVWAuOT82jASx5H/9Q
4aS4MFHNI9ZzEY38MnHYw5bOojW9xMVOXoWDl4CoPbgvHbi2vq7bp/WN0ukq0/tp
+wq7USyxRDh+26/W8ZoxyrVTPuyPd8S1Dl5wEo2g7yT6puAtKECLPRX0pq+t5fM3
A9jp6Cz67jCoZS0O2wFhvHBn10VfLQKLaTpYPCr3xXybBgMju3cNRkOhoKF98Swr
qOCrPDD8GwmXnlF7ioo8Ly/K7lEGagsRqVJ4x6TKEYhToTK4KHhSPdNU81gabVzX
CQ2Ibfr/LVG0+u+EAMOISfIwrBahWUlPd5hruMzyAAcpxeVtx3Ghn7+eG/rmvPQo
A0rfBim0WGCB6oDwC9m2u8qS7H0HqYrnwMyuqygsg9xljA9dYIfBkHIh08lS3Cd9
hf7C98nSor0Vzc0MYnlWmFCZln+30KjtqT7mnlRiIVUMd4M7UUCTIcBOt6QQOtLQ
k+orasViVlfWgT4E/wpOiALcfVnyP9He+3473hCVfi4HQ58J9E1ciUvnTiUILArQ
OLBz7pz7SFBMWLB/0wej7kYgUkfB23ec+Pp8PVVVXuW6nFiLu1tH5rYTi2IocDv9
FkMGmJnXE03LR8kR8YTGBBWehB6if6+rnXDMe+CIfAYvItVcl+9hync9QQWYVG1o
EL3sHSIr1YtSOcGFkhJDKNNN2FQtxi/P2BR6DmknH9S2JgUrlGoIs6MvMchFD8w0
l3Orj3guyUbcZKb00ediQT+Heuos7N8LJgUvWwxGKm9o7X5SfIgNHYVf4m+Iih9Z
+PcBHuVjiYCIJ484y86WR/QILFb+WAM2YU+sbn6RA0+k/Rh0hkzpvdkcfRDofy5M
qs7Y5kxHMSklGgcZ839oYcpQDDOP7e/bsymqpPyS8Y6694G0oM3VecQxX7D+sb+B
mKj6MMGTr/diHFb5JEcxlM1pCFEsuOUfQdnYxgPiiB3+ixqrjBEQcPN8jRDSOb1r
w3GSjrUx4yJkaI4YwsGj0cIXVTglYLE/YW9ro1moCOKOvVFGWzt17S2078OBD7Uy
0O626MHnBqfOpPt9XL1zU+tPHFb2UwSIe6EaLH35NYceTaCUvQFvORi0VtzMeR49
umriLsVHQIftIv3sY8nc02f2ZSr2atf/vST/PnkPKj6XTkQZM8cmdTMc7N4G0vwp
TIqnqvgfVICwECkmXanW6FMpzsoCWpKvzuXJcnCZfa/NChYjj2se5z10UVgLjyFN
E51JBzzEIBcfr3o9QWT0WkURK9yCv6ahnbDHG1SvfrYw/ebilFVz7hxlQ+ml3rJ7
X6YMJlVjwHrEzpuua0oEyU1BzGNgqUZKlwiythWnFmu6QnAkrtLKaa5Rxlcews6P
PyJIbXHRezyCCJp6147gK46CPq9eL2qkcssYuKsaJr1ijaSTgjxbKAIjuHV7Cy/e
mHWlTWCteXPYPdTBP0i1PyTXFpIcVbetijEUSm7zVYinEP/aEswytYhy9ldLJbnB
EpKHenb2pes72cUZg5U6/eW+5G/Ys90lTu0Vqky1lbFEOclz3lC9Nu8Qwn4CLnXK
1gBfKjvk3k2io2IMbkjkqPsfeuBN6AQFauxLEuJaxWpxHDBLixgrG/H35JbnIbFo
a8MIr6xJ342TrA3WB6+kUcYsHRCecINM3Dq6ZRpywzAqaQyWRZCJy0jpYYUDwCHO
yA7u85f5fN6bv6uNZ51SpPsqeJdXh8rbEORHTrbopXuQnKy+GCmQkKiJTR10ijUj
ZwfZpLORyOiiTjvQ1X5pxb2PwrOSOhI5MWsK7PEDUKBpI3v8rUChP9IxMMzbnx6k
si1WSHZMo1sChgfY/vqnjSUpUql87MNH1jCjJ9bZYm03SM+ZmQZlhfKz09q4Xhf5
uT30Cmo2wvnb6wYMQhi6MwxgdK13W5SIiResoPHj87ezpVaAZQJ4wE23U2tGHD0f
/kKQD6hJHDklEd57QiXmSbDSCXAPtP6c+xVMKBEJpUZMYq1oH8MkKPr5ZTSm4ga0
9pHn4T22bGA0/e44uoAH4szq/wXFmoTiagwKWpFqioWLioCBsp7KADlTq2Fk57AH
u3eAM0ewl1TD3qCDarLLrsHGON7wB8kFBNInXYYbmCQ0qfrU7n7fflCEaWIYqLFU
cgsIO9t6Zf4UfDnWyo6FZ56AWI02qiP8yeO3t7Qhcy4UdpDK5nS0FQdv9TuUzQ+k
vqSULUUN+xOG7xZIIe1QwgFaoryMinHQq7SjhrBGTLbV2XnEcHDYtJmwqqQ3Eg1d
4u3qqMu8O14PjG1l+ykpFmJnct+BBwDssVmDWbdZahCA1cw+oQ96cFjxG/bYFHU0
6iTntadIaKvjDKfvrf7ulXvqs5BSa41aGWzSNYUHT+LXPVeTnz0/mWuOmblsuLLM
9fzi+J2s+DULs1Pq/M82Yhls4YX3sfvydi16UFTRExDWAVzXiqtadP+nP5RA44e3
MFTqFwgEJKv/ukmaZoAkecUVmt8tU7WkwGQg9uyPouoIpEgeZMqjMA+YRpcE7y/J
1PioELqYNDbGjSqeP2sIHqsC/v6EuIdjPE54MW7v2mffmuTqAr1t9hlZE9oeQ1jQ
Qp8C94bGLStiA1Su8lbaiAAlqGyagYo+QH7lMQ4DC88qG8uMYyJx3TX/ZHbyPcjv
uqDRWbOrzHNOBnILds+ri3zWmtQIABxujCrvCAsynW6gkOJivF7adT+I8wQRmU7p
C8V59qMLnKCFMrrDqAMuo/nVMqMAIUBQSPTWpRs2tHcQ/6HypjdTR10hEDstDLbK
A2j4xcDQvKpY2v7GR1JoAXOmYL76usYUhiqaqS63A78A4mBJvm0xXmewppeYshFM
RwV3H8n8y8FzssXcNai3b1b2DPb8ZhqoFO9v1XW96RrBAQcvX58Ae4UX1rU8SxoC
xjSkx9hlQankvF6/VNBvv5SL65aQQ+dEfOdK7ffxzRhY/c30LxOCptODw3w9tzmQ
UoU1kFI1zi84a5fWhAtWcVnO9f5OIlTbOQJskcrdeQ9zbhN8AgURbyQl73QFl0MX
7eFWiprn+4a6sUpVtwk4Sb5V2xAMDHo8/5lbAm4fq5XBTTQlbDQsLzsEmi+3+eLl
O5GBd6yoInR7hUKfuvgDOxuebU0IknTZpD63GSgcmlaqVG49Ku3TTzH+bQWQQzfP
gb5ekXFrxGjlN3kkVQteQo9pnG9nicxlcJ1fIvWdrQxQ1WKOCdCPtnohs6DzkEEi
OLnYkccAUe5griuhoaM9KXvWBVOyfxfueTAZztVBkTebJC49KWpWH+hZmwdP1H5O
x4RssViU05xJlNN4hcT4ivp4mKBWpx9YMoLTpDFUYX2SAq0sDf1eC2KVEyKNY7fh
9JZlTuFIyVYMkpJhMvvPUZ6MHQqWZKjif9WowZqOTxcCrD7lo34geJPer7dfnPpn
wWAjsIln/5nojgk3yiVbl7/XppPXSxXUylbbxZzyVddjNaBUDB4nI+8LQ7OavpSj
RqTY5Jhi3RgHA8vjThWmr2VE/8hVUvyYZjlLoS+VVx9fj5T8p9ROR6j3ildAHkOR
ufq4CiF3+bSC5Kie1Gvld7pWSGipDoEO8OjQsT8M9u2jGyoym05ML4pgr7OVto0k
xPYLBO6W/LlohmmHXZYKy3xBcVDdfz6SsOZiNrcF1g3QNJFF1WYsLq6zR1HzNjYV
u5uYkjdRBX9SctIof5cbTVIsw/Ii1op0fAMnvyosgSwpaHM/5OXWoOlfwJKxOumw
HhQZZWpGbCla1aLefnXhK2rJ5/mNXEAozKypq0GZehQbhIaqYCAj2YHAij2w8/VN
3J1otC8yGrwSfbz8y6kYnl6jx8ovUinfC3WQLl1Zq3ZdK43W4O0Exd0HhZOVmyjK
SFC2yFRUUAHta0ovJohDHQwJ3fXPCNZ6wNPJwFdm1kyYtEaY4gxQUVn+0oPxZwS1
4PL1CUlKH7hhmwcIVnE13NYptgcV1AWto/fxosHfqpvuPC/bm3kCq7XN7l0HEYgF
4LZLAcmEUF0fNAfaI8MV7KsxsoRPxGtfEwq4vAnVy5/AFMQUoBjAT2JP6k/qb3e8
nYbCA9ZHrkRFSdUDuz5Bo7eDRxyKxiOlOzFOv5i4R8OqwqWaBzWZyYf8czJJltbG
lyRDdkJvtqWv7eCFnx+5uMkrsRFP6u7pQzaESuc6U1v4FM1SNiC7siuWM+lBZjMm
Ji0naoD/EfIzTemsbxYCh+arkvgqbbdhelX6Dpy+RNAp1dhHXV8SKuaTQTIw/pYL
SamE6BNymlDJAlCTWJ+UmNVTGVLAv+zBLAqQsrtEWgucl88vYJBN/ICbgGoSGnEe
L3Tfi7QwYZ+H8WeJDWi5nwx4csl93s+izm9cwKamlFAGXqAEOIxFF/Vts2uUpcNj
KVJxWSPeZMdlcGosohZCzyjKdu/Tw5BHx3J78f25c6IdmNcgRxdcKWqNI9Tt+U8x
/7sK8fCDYVVhvh4stDiJI6IHLz69KcrCel2JdmNV8U78TQxevuwREs8HE/Sd8brA
huW6R5BCwe1xoDZqWhPkmRcd1pokYtVeXciN2gW1ojId9ZJlGz+B/IRf+4ZGgiIy
IGFrLGgtAFa8asd8q1bzsAZivE94jQ9N3oUC4kt1E/HFtdgBcSq+rpsgiTwfQv5y
pC2IYWXDverLoldWotMUgqMoA90G1WK9pd4TfuejlyIESg0JqvTk9FhvPElHYkuo
U8662+71ZhAZuTwUiLteIn1rPhGlJ8aU5HJSWGZc4H9RcbhQWMW4Brx4xTB/q6ak
MHygx0Met/iYFPXFQ4BA8oZDql9hki5niStYID7e3v6P3405RlrYcbK/00AyOg7I
W6mC2imDpD7i57Unugv4xS8QH1kkzF5ld619s0rCw5r8YHvNh2fkGJgt2ToWdBJE
TC9z1GznqW5M54NoVbkGEF3dM/0q1NBuoAvC0Gk0ZatHhC83+fLJC2TuDC5QSnzT
SYlYJ4axXgvIb7Hk4g3/XBhrEsYBTENlC+CmsbNU1uVoe+SfyeVjaarUVgOH/kCr
XEg9CgBHHX2KCpAdTJwi6yUoOi1uHCtr9WQIheZ6Rjhek2oXCtJTN+56BnPyIJ12
jsb/L4VBEqxos+FzAEQ8vvUxiPd1Crt3WPvHnoUULlX+GKpamc3KqlZ+1SKR6kPD
x4OM6BKeYMsvp5PD5jfyNE2XKT+Ic4BHWK8haeQT+0jpVgdT2Qfynk4J1NloT72q
ncz3g96uPM+9LC7UiD5MbQa9AnjCpFQfe79Hbf6VgjJjMDvvbUio6lmLnJ4xFWR4
9BLTZ9RJRDSvXLLKJbBTS7M1kMhJkLlfpVGp10g1mbPkh5Js9Qguf9jFe3enw1Sq
a0FabE2WdrcqQGAu3T1zBRnBjnfox57c9iGSD64pFL7CAUhnYSxI0MZAQbLs0HB9
fLiz3jH0ZXqUf6rgyIchRzAVYq9pOsEAso2J615hSdFT1XBd22fBj2qOjTSmOTay
ZLE8So2Vs4SXNjfilKPtNWjezQrqaj0gP4aRm9JNnaPurT2xlDx1wGW+sYZgU3VL
ASaXvAV+0gL+OJbinQ8cJeg7PZMpT20zbCiUfnP0Cf1V4IGEEF3VEY4EpqzuktgM
8WtvOweRkg5nyOGbBBhXcwxPSlQiX/2mgZPqD3jQEYWDZqIU6++YPF+c4qEUAMHz
6UjXaP5OOhIpVB5I4Reg7tNuUGCR3ZNbTiBOAMgWUGFhf4FzRnnVZ9oq1m210JD1
tEE/O7ZiwD0b5oJjNgb+iyMQb1BDxDxvIZlxmpFeYt8ZD+o5oHyCt8Pr4wsGPUag
7ELoIbirBQ+0i7g2phv6dCwsbrRi0tivACoOvQH1jq9juF1nS0UPip5quefy7Yj+
4VgdiHgzoHWarfuusevC/IvbcgKfsn4VHoA/pdDEroroJCj8+w7hFoSvtuWUZ35M
0s+8djhLq0jPc8mnWvqEhMhlNf6ZgyBqEOKoamuVFqnlUA6JnxMJSNVfV06dQtuM
46HiUyIRpIxbxoRrt2YdaRSyqDJ7o/F77xgrl2of3rlha4mlz6zZzFCbB4S568ue
TM51iHfEAYlqflgVOLBH3ZU5FIHKrh7vq1PKgo0jWRiQ54VdfFnWJLT+Fa/Coi3V
oP3C55XJAedJtJhhcBPzd3OhvgutXAZrZc8NMXJw9ScyFsOLtTKDxwpVcZO37vmQ
cvX5F3QQqzJbY6s2BlvOMlKKk5e/KYZTj+TFarH0o8SgA9+LU04sw/ggdAMuyOOK
JjrZnuvcouw92/4GO0FScrJYiXJ7ll6YN5iHbtB/dXJ0XEBSnB0jv+q/8vwqWZZl
xlayqnqaj7/fQqpB1tWglRxuiKHJOgo34InzMTDaJdvwXKdFa2sDIp2+ga7otbjq
oCQcbqcAv73iwUZCInfnHpaPc7rc5TwoaK1X7V/DMXFXPPFQRR0FO+FThGugAXMN
b6qjL3cCANV2dFZr+VjnkeE81cnw+bgNwpMjBtqzEJ3sjBo6GdZKllgjBjzK+igr
G0H5z7WqYd5UcM1C2PQhzuvhc4KIqgR7As55z6DNvJCrOwUk+O5N4l1JDsm9J63c
vm+atD1O41FosHqgIzRkoNgqg46BKKWUbvivmAXDmBrs+sl90MiQTAzp1L+kw7xU
odharqJDrJiwoTr9mp3T4ON2ssf3UKlCmKOAcciKEBZVA24uCD27oShSH6m6NqIO
4NTkKfXfhuu69FAP+bOUWWMtDvuubl0Jg7PYt8gC43XKq66BB7cVxHaRD0DGE8px
Vyh416ti8jBpm0DPHxJ7BEFsCnzBZY/myEkhtb2OAJJwdVgjYC9IeIfCpO2ecI53
9b+Ku163T/PZjee0sHbCsCKrbePxYn0wXfohy15ghfgrOvQf4AFDnUkXTLjVAGed
VvhRTo0PysU3KuHAcBciP904SDWtMOV2UNNgbCH4x0NY4uKszeerGr0vqcej5Oy2
Zlsl6EB911FsBOE4cmTNpOk+MrUNNCk+PtI3dgxA6CeAGbihqzHdSHleLxrmoH0L
suVgaZTTLlYfj/rASfGNJ3HjauoLHklpI75O71ChthFYaIn4oJXKgDIarA1h02n9
JAIPJcBW8rTlj6l7YcB1rns7gsQ14FmHf3h1W2A5KbAtUZS0DBLsoWfxjOJx/aG7
8PvbLupY3C7o+l7r4OfyPyJaRAIqev7kqoLzOTO2AisDfvDWJUml5CoLUqEbVDe9
O4f7UJbGGF+2tvAn5X+j9zwneyBh2/Soj/IDBMPJrr81gn/E5zTeCTA5P7oq4gtW
8KpfEH7p8sDDx7drzuaBB7g69uQAOOh7bljchLzct9kuBW0IGu7UtHSAT7c0kltt
0oFEu//389QEER/RiYxDCYzoWkng45njqMIjX8q6J3maq8g58k/SAj3tQG06F6MP
B0eeX2Y2kj1pUpe4hLgXuZZZYPmjdQwk2ABtoRIE7ztRwxlD/qptaoQfh9WA+v/d
3PTRZrnjxprjAyS7EMriWVtHgu+83uvKMi/DUO3PQw0O9+zvt+0aPF9AdY9mx6mU
kKd70orRYX2L+CLvNZVEq9cKAW7ih4UDt6EOR+xOVngDvKXQ0cvcMywjNXS6H96r
lPo62xiw6HNzP/SIcnjA+hPBuJmAb4/iXnDoTpaR5pmMMyZE0PJmmilb2ENNXhMf
KxhFEWfSWfu/tCrF3ZABoqdvLHO6yPJyQFhHJ4TmQaMtPUJF4yqtYYwkL408yOIO
WnYiPqlAl4xmIeZBRgryhNerBKhu2CLpbqZHEL1tSI92Jv5A3Sg+769SDj3MAEu+
MlFR87JpVrpmZfOVasv1R8APJNwOAMYPXB6XbWGQlkdRdNXd7Lsc9UjDmKf37FX/
NKAvuMQe2oUsAlQckJRwHA8uiYxguxvCIY4aP/kd/YivcFFSe/O/vWlXYDh6fAve
TKjgV9bJUQv+SEZ/w5gUTgngwckwK6B3FWBp0jwitGMitnAEBrZWHJ+r3fn9yybM
YwE0kiurFMDN+9mPcP3IuhmzutuPQY11yn/M2fRQ2IkdbXykDVQQeONsvQhkwAN5
lUSOJqhMuy8ocf1//acEWWK/VvbBgSF37m+iHeP91Vl1TzSGZJzHd6M7ufgbaGOO
UAvtLJ0JCsPoJQMZziOoTLBsyC50VTVE1ye4H0Z1u33gnrTpUjg/8BvuzKAUecme
SLLfM0Pr6Q2J0uT/OIH8ung8iaVqggO3emJdWb3VRy0teGc0Z6+sfVRbSr0/1o1F
uXb4C8IQAAbrzr84PjWSCjc51mz2Wrii/wKru3T4Q/Tws4+pxVDlmP6pC6TlsRHy
5DCKKSXP98SLZs7O1rexAdOmlM0shnjnKPYEmFOG0c5VcMFt3q0WY0JX05Btl5Ju
LWdLu4eaNWATkdnR0dcV14gQP5SkU8WYHC4KytYSGi6IBfq+stHRzXjJRTFS4yMO
Sp8Ea8l8wjXSBci/XIzu3b5v2vkj2EuEHjL7dGMuAMxpA8Q+hE8uuFDBb3p1HJoL
DLFnrgwh9x9VcjqJP6ex3pVlglr49TpCW2kot74COHVAzyIeWMNY6lbtEFRax2bK
0SeIWlI0foy+0X4BWhrbSW/3Kbxc8aK4VzCar0mSHBEmg1zqDssRRxhN+qklcDzi
GLeyXLPgPdEH8NH2vHHvbKebShOWLXrZy2YMWF4CojQC5w8ZA+dKIl4mCEOQQYFe
JZr2yu8Tj4CJFTKSDTJMiuPHZV+Jy2ecQvGE8NOd2+CxdCGDLCYbZ7x3lDoFynWL
z3mM2DBnGbmYX3ByEfbz4Wzb4PlA2u0p3uwxCrZTWFX6AyTu6jcN1Ks37ZOpdSYe
B+/Lppu+FhLxcgDE41BKrEvvPB92AVt+Cyh9UjBQSoLE66OfTxmmVDoQFthyqj6b
p4pn+pZcoHbL7dnPLFcEAvf7XL+yWTrutZuXsi5Gsg7xAVFmF4amqSZ0V+DDuEAS
b0pMg9iT9DDUVjVbfgZQOa8JSqX4G9IUOWCC4EBdNyJmPoqelzUFnmSKtZe3Q4dh
3rV2HMHshby24QmZQlz/BCfDkALicF4yeEYdRdXLQZhur8TAeixNRvCxYnyXPt8O
L8FyCzoMV1e3CPbYulhAv1X2ZasWcREpBWFzNEAZET5RH/xj/G3D6Xuy1oGwQYdg
QTF9MiSE6sCDAaiY9q4ZpfGr65IThvRcUAfQI4a+PrPoEaCyFF6fZV2mZ46r8OX9
5xtlb3cteM680FRQ0plyRDdoaz8N2+YA5RVyYvQ0EB8wsuA2R9p7b8hya9TfNhvi
inIVLr/HH6MWA3WOrq5/Ci9AqL1fNW7vFS6UERZ8MXsvUdYH6MDO+FxwlPGS2bxE
NJcuv1t3De6Ml0ow0SIf39leZe/j3NiMJew4iNfiOA3IumCkBJu98kAwfjM/4oKH
pqiHvrCHzVcNwS2W4dqDHbunTg3ZAriXlA1fHmI6PCVl7SB09kLV0eDls+BO7ubt
Kk5Faivf5dZT+c7tLKo3dTxHk7HV9pzKQiq2TgM0E3UxgQzXLTcUo5Sdi6jBhjsi
kwP29ijii+zIGyhw5LmOKEICC47yGeCTkpXo/efb7cfPBpnm6I50M8nR5Vzb9MbB
I+dlyEbNBsyUnojrCcmkXnOCNk+YZjnqb/7Jy59sjQ3dfq9Bes6cz26iMJS1f+nm
qW/eChkI24Bzr8FWxFFGQ6vF1/E0i5HMr/rWhrkfXWmT4kaBij0Xp91YU7oODdtY
k/CKFX53s5IZ/Kt/nLtypWGoOUYNI0Yu0hyzrNWa0zoakP+ObP+csR49uCdFLqtW
CVOw9tTTe8aPXYIhj9hj0rTVBeyRQoONn2Dy9N5HwnOabcyxRwV6FAbG5dTBdUOr
rzB8B8hHwCluxPuOEWSprb/KWW2hBOU+Mw1CBq2DqWiOOGuzWkqMuHHNKsgYjyir
GqNF+DVW6gDd2NpkeNxuPZEPcvZSyOZllcRmoqoepEU+uEKGuicWivhYQA+fsLNa
JmGIGi8dqAXbwQtLMabaTzyA+Yp0AE/L4EZTP5tSxojJ+dapqxaWeNFjRi/Gbtpu
qJM9B4CnqlfQj0CQgip28q8bpqMCjAGwpjp+673X2BTuJUP+YQIuC+EMbppyi6tJ
8XY/wtSI58PqwOrKCEwTF0i/zcOeyMSGZQUIlX6e5r+ALkdnScLsUnXukJkrgNGH
ksKKis0Gxk49+OAoDXnkaXl8BDNlSIXvAXJTJOP0llAXPMxso0BX5N4HVHnbJT5K
b7+WxcxNSrJMjLwk8cuzalBPqZLwDULFg07yUWkERfLJCVMx3jfnCoDySRMkbvkA
/LBzoHTqrQPmUbGU5/LFDayUZ7N/9Vc+9h5ObrTILSiEpzNZ4FNHDJ/84gIGShAU
IJ6bLCwJsvK+rwkGO5jlHUJCsB+KwDKknxtGB82oot2/1hpPczspD5+wXs+XrnY4
drF+HuZp1dAFHCsYVhDqWtNZipcg9o/l+lSaF/FJHZ1f0QfWvgfcilplV2dhyt0G
NTkAj55rj9tigDjuTgGPdFDKX9YbyGnbZQOR5Hh/YpyoSRFznhPsN89hIsjvncy4
FuP9APlcqq40fekbZDeLcpO2lp1favldJ7Nd/LoQq0QsWjhicpsl3bOCyEDTaS8y
FFEKNAwUvAeqY9jtwXnY1/gyNCZtSabPtT5IxdZ6qGDYSyKZ+gwUItcGXymLFKSh
IUquKAn1Y1KsGrzpHF2Fy+ckZaE0V3yPXzrsTTvnOfMTmSZgCMjpPQKrc9AwqTMa
2X5XEcs38/F4WPwo0Pqc/YKDynrM+r0a+5DBhg5SeKcsUWk3XXdMBK9hyImu952L
rw8aeKLYpy0q6z2K+D4a0v4LaC0fZHBC9PktfdvxbTmj3pN5/Zq6iHFxTl7Ixp0K
kaOwAGaqboIxfgNXs0W7/slOmzwC9PU6nvO17TGYHWRwwi1vg/+iWsd7T/iM7PU1
gQ0eGwXF+k7L5q5FsLFbLJvL+CxqXe9S+tpwYOQM2VRvMt4aH+x91KuGeract5Q8
5Q9zN3i2ZhxezK3iOCGsV0Y//d0HOmpsAXVLPChVPZFF46x3pCKXTkFSn5BXh+Ib
B1r6Pu0+f19kJbPbOglFWniciMjVD3V2pRTNtFER3Z9Ah3vIR6lIDm7LogL0mOXc
wOONh28SV7ZIjFkxpJy7Txa20bYUWcul+wtf8Tm4gOQViMCBF0eqV0KoZSPNX5YU
fsUnMBqqryZxtWg3tZdFowXzQBMgoVvgDEpUrlKUMwnGv0txmUC1+n0qW71cSBtU
Tq3AioPzm+sNpyBjaQTUY49DmP00Wl/+coHViSNoRANCrlq7rQX2mjj2wBwboX6D
F3jpiKw4ePRnZQAW5vgBRK7UXIeI++sxKJn7UhSwlSscSyFJyZh/hkKv/KBgwhcG
6u1XZujTFvy2Ms2htXnGka0nTF+UCYGUMrVDT7I/BpXRNDYeKh4aC445SzxFFyo+
Ualraf37tEWGV1dxNs3aTbx/+vqT/nOh6TM0K8GAwqFQQo29zhytzZ4i7pKM82YX
UWNcWbmk1QLaDFyMOJjmolhYxCIAM9v8oDS1iPxHj8sa1cDyPrnqnrlCx2IumM49
zofRPSsVWaXtrUU8LDPORBJWIOXkoqoiq5cDBLmqHfcnoWOSorkxeI4YdBOIh6fq
v7yUWXjJwAiXQatKvBMA5y68zHC1oQoZdQU7xGDxHpo6Z1cdcaZoSspDtyI8uTNN
YAy0a0f4d91NDJrN1hOdzuw9i0wbIp+Jd/V+kF/hHXOe4W0B2L/G43iFRkIhrfCD
qddD6BxTAMzNVFfsCxRj/NqEMqxe73Iw1Hgec8sXNtlpEbCnX19Tm0JAm1AEkhsP
n/kJZLt/WILb93mltoWq1WYVt1B5GWk/jVn2BhwDyyUeI1br+bu1RvsdM0g0EISd
t/WN+Lh7ibfbw9KLiFE4R1K1rk43t1jAsqbI3uUMGsX+YPvyjxwJI10JNbrbST7B
l5fmZKrJB3lPRrIUrX7Wt+2ZlUYMvlLiCfMonnvMGx9JnM2OIWMtZsHGKGKYh2QN
2kerlKi6Jub4e5S4d8+ZGgNdaWrzIeVDrNhQ+iF35ITe2MV8rtcDn086pCG8JTeX
F+UaLE5lVT3ku/2wHJwn7PjH4Q4HAIvxmn/NkBEkaKHgMiRxaitekBGtsos8JeU2
Qk/09rKtD1Fj3g+Z17XVHaAlTlpN+wa4P0XdLi35BRTVjDaQez10QK0/WycPEaTm
BwQMSs50cVCOsBP2BWOn1vT3QXhIMRQ7AX7Sed3HE78x/4KYejXtR7EZS1UJFxbg
8bWeQLDABZmnK4FVGB/vhNYxUyihh9JcnC6wmWfU7pbFaXaGRmSGQwKF1Jmle1Db
oqqjZrVpt3Hde+95wEnbvnNzK0v30tl88QhJVqHDPP557tvChtsTxW/KC/jJveX9
RgqwYCxdeTvEohaB4XDIjtvhb+8mpSft0FL01IUY4OVwLEc1EqH0/v+pbUwSVzKL
ByCyh4j+1LBmhskx+lKFFmTCUNo10UbI59qGeHhuupxcUKBlga+TttpXHjiGgH/y
WRSrCSP+/6vXVowrk/sz4q7YvlebTKD7eusDnyvFoTDtqEwPHoCIoztnHUMlpXOC
sX9ndg0eW2s2MdYd+jiPY2suv4tLQsLd8VOWabFyjsrd8FZRIh5OVjSKj+VRzaBj
bjZSWBj7ROrjCgMfCK0Itzu2Rkhv+xhgs6XsjlkncmcS98IARa5uASt+owFRiALT
I/XAxS17QKlwx3aGY/lVuG0d+DSdFwEbg0qWK7AbtCpf9VUNtJCtefcxcwlQNXdJ
SbE+a4v6wWBPDhoCRwGENnmuQUBtlas7dCPJbfVRBHSvm3fwfKH/PALvdiYKFDYm
JP2mws5UduTzgsFVhxvKmWK85ec89kBwN9+BWgR5rPnYKEkRAQ7Ll4i3wVq0Otle
b0vCA0GHzfBmEh/wDhQn6BA8P/Yxo8zUkmQxmjLQug5sInOElxzzYRHHy+J2UFLA
IQe8c5nD76R4ur6YIcU4sUA20zNwz5Sw2BFIxjBFLjAUfrrLKpgeplBXQVSLSUQs
uD/wd/eDQVvmdJjUX1sIwBioaFXrcelXOzbPVoGym/PObXde/Nh4W2GJe8kJNw/q
mVpVaXM2NP/oSDhUHdovK+XuE7UYftvqVimoir2D+0M4OCJ6lPrlG8j/K4SzSSYs
U5w62HN4Ni4MPehcXDA4YePOlBttb7bTPSRWyUhMXtzzGFw9+32DikvK52Ic5wRy
kHTq9hwcUFVPlXn1ue3Ri9UVI0Bsx33sPkRiUHKT8lcoMPs96a7BMXeSf2f7S1F3
U4tMmaPkkrIGuAH+w329+LGGCyM7x1h3MO8fZb3Sy4u07Or+IqqiJeHKo5u07ubJ
JciNG/GxqfjsyMlxY4RCETWcar3O8/uqVBCQww9PVIAUJes1VubRYpzyxuRmHUW5
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
QhrZhL1bvXr4YLHG1qOJXjMeScvxkj+JdMkx3hB2ah8obm7S3g2KL4aXIf9+i+wB
aCRwHDOXX5+Ne0swvciHN/sL4oUx/nmKgOdGyp9P809eJ9tntYe16p9kqMD0xCbx
22OtEVtzGgYH4meT0z+MyoLF3ZB9MSNlYb7LQAZsDTSWy+xXFJNQvnWhaMKmWaJB
GjRhee5ceNFbPLKGQgbBlYU80RJnqnRggrCHTJjlL2mp7sSCteYg2EPJlwiUDba9
9z0kWZuLBcMfUzPM9bphGz6drMLPRuJ3y/THjSMX+sI1Ky0TXWLKJvECOfTQw/i3
AFB7/GgxEx92F8gHjOXmbw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 21648 )
`pragma protect data_block
1hK81iAuHPOaTwIkOeUO1R80CMLwe/R4X2WS5JhjghjO5MM/ZZaF4orUgK+bTDEr
cjb4e8L7JkTyydmNgize5uxWlvXZu0QapZcQeZIOz428q1JkZ62fE1v1lj6VxKMl
AeSu7xhp8wm16mGlBwp83fiITr+dtYwlwf+rkU4AGEAqvkW+OMEBgum94DQYAuxo
HAE34GL9dhkxPLfFf7uiHjYORWeTfa//9A41u9fnaxNYinnAnlWt1JAsft/v3Osr
QBCckZVd52M/HTg2yKwrmDiTD+3v/wglvYVc62Xu452hQsnEK3WNV1EitlD/a731
4rMQoe4Y5KlOsRzo9qIRyHGpR13VNyBl71P0/08g5cvWilyb1RAFLymGzXuGoy1m
77WLk4LKtPQZZ2gC/cfZQs49Cyi2doIefq89RtoOxS9Slnm1O+tMKrcWjPpVIqrV
4V5Jes3Qzumt6zdj8QD3WulgwLNM0d6mwAd0WX2emq6y1NpST+lCd+6YuLL4quF8
zBTww6Pf7zXe1dny5Dw9RRx+sU64k9Tv9ruEQOQthFwdpgumT9lg+pKoU46gslQX
eUD0Y8pU0tU0wBMEpwxkjOCCovmjOmzPBVLywdlPLbF0Mh6HFJXxrUvjCP28AIYd
rauiXOMN4Hj2/MIHrvLUOy0DSKleyem1dnd4baPTEciWDLMlKlXq2y7zeSDVH/aj
gFVgNc85XzJAoR3YWZWn/F0ROIzp1pxva32bAtPgOCBaOH91zQgpLhcBKPbQLos5
i7iqlgrmUaLV/+OnCz4jH1Iz0KW4TBgQ8HfGSzMyCoLMzTHLPjaG6okdkk/aVPu6
rHTGigBoLsmWz9T14ZVcTlyETdcgqDo3JgLVVRlzoiHyIt0T6rdxVd/AQlkH4k7V
aUn4ziaUXVGZyPmGdGWzUANrhoAot0tDnvOQk5dCp1JeoArlEjxz03t6Rd57qK/k
IIVKz4GNImzWj9bDTU0u2lhsRk50ZjO+ZBUGUoqDJGwRzDMrdqvwMck/OvBZ+AAN
zJJZF4QT/P7ABslw/A8Ta71wurNrGEhwHbBqW9w4VmvVAIn217hntVkdnAFCjfjW
mCxjT6ZZaidDyNYp3Q7x2MOhjhgCM+9JdwT5Km2CQZ2rsd20EoAojCi2m5VBCfQ2
YPJoJDW4p5Xbp9NvzCiEbkSMhOK70E914IEmXKpSr6DEy24RqIefNN20i0k0efE4
vZnMFOoee1cfjtTCpgBs1SOj30BF0GZ9kkSDLe67i74WWqhizJ7IZo0ymE6Nx1Cv
TlUJejeHl603gY6+tXl6+K/ZWCtx5MSpRXf5ww63sE27JqpAvK3Ud9wQf0hSws/u
8Qb3fHCFQfsPkF9B9Mz4MUexi8jG+oQk7IL6IkK01jES6delZARMH2M5MvDmY9zM
4TUsujLa3YIfFIv0v7IyL1awcsRJ6Ls0aVc6Re0qUuuiN/Yo7LtXSI2D7EBk5njv
E3ztpISMw4luQ4sdbxyIh0wA0x+7fvnfOWuAyJgApDJoJ5tGtZ8/25nWtaqRUDfj
Q7TYkBqrgfRqMfWvSJxLBUt4IaCtuNVcZ5Wrl+baeOWsPIttdKGg8LwLYph+WM63
TOWLWAYut7A9xIarjK/0XlMw4+CSkZrmxrATlpvAcPhRIEaa7QQfgyZo5tAxMlHP
PE9WM6uXDc+SEXSjB70ORhjP7HaI9BAnaDHmV/5MWBXvFKguEYW9AQ900W39MfwA
eY9cFQ6MTx0ieWzK2V0ckA/sWve6ZtUFrh0YxnLHGRDH0lLKbE7cJIFBMhXrX18B
SygPDT8VzRqm5WPtTD4qGd+hEUgwYYCwPy45bc7RqOjhR7a+IcZ74FBvSUdVpVwv
y08ItiVbVNWnbnlz7BbiTxJcts7TGc2ywjn76uEdP9kSMQVkdX07E4MyNh7fSYyU
Ar7eJTO61gWKmJdrI4LKWDhjVcnbDg188UfDsmzD8kOg95BOZuNYJ9ZaSWxJxFSw
rxx4FOBqVL3R0WJvhZ6Q4WboEUif4IS3KfzkEtZ/vqD2UsRwp9AS5yr2ChCh3klj
jJN3HHncTYMancpCI30meulkYYCnOlMx40AVy3tXYOQ+w1lyxK7TVCGt09KCumuj
JCv2BafdCs6MDWf6nEZF0W50euelrQrf4x1qc/paoEi+HRhVvysofzLBbtNR1EIf
cqVty+IFcdPGBV3N37Kj2J3wESvKxqwKTLw14P90kpGc4k9PZKPL1i8LonD9mjNt
KK0nYug9qgT2AlOVEpH6wHa99apRv84P6VvWPMaE5Td/cfU9LnoOAWwJxfCf5l93
aWxpKaJoFl1tlfnN0xR6rxLMmiJrn8FcdDR8d+aZOHBh0K89V/IMde+1+HOmrIjB
nZAy92hheWnMahkM0URHuoao2jSQPXst5aIiWDvIwSmCKoUU/So5tYX9l+3+CNPx
yUw9lnBs6mk/QY8Xz38dH4crgscPm2XlqkD4Ucf6hzUaFarnKBg2unNJLLyGo4xe
2LIWcz/DX+bhDvILoEpErg3BVjRiE5OEld74UOldEKh0wLnWiDDz/Cxn9ur0BjUM
FfjeUaXw73zwT9uBvmgcD6j0SX1Wb/BGeUHLCKsnEEDMEhpxOUU9A9PRiC5CFOmR
Nb7jcVeFVs1nFd13AiVm2THhSIvnLLi/ihv6O3kzL60beNmDE7UdV6UALGAE5grH
unsLrAkhCdC3WkyvfI8JGrbkYIMs27fxSyXBhsWYMUXH1bnj6ut9akXqqCmr/D8V
i0NzkdN/41nXHTVmQoUFMZ58822yKNyqSFFxT5qd78vJpjEcjLhLpQJPbIcmIPTO
Da0heiLjgn8ubyqFcr4G5ZFPxmJCC4CEdRXP14JQ6YovnjTveNx/wu2DFEhNUcZ7
0eqiBM7GYql0Jye7qmUjGOO3cshypbSVWIQlH9EKV1SgSoJVBm9Ih4b2p7caXPME
27t9SwPvxekcTdjmBmlo/7HuJASx/imTLywM6Gr03KC7EnxgWWwMLmGv1KwRMJaX
pdNAj+HuvyKErCIJh2Yu+Ok2BYeJVumApZDXASd9TzplvNA88pihAyCE9Hj2el0c
RW2Jd2WJTXoGT3YKt3n9SpCPAtWwxu2tgkePTrIODfFDt0dU4+JbRBbS9CSRWD7Q
WRNo/tMTGNyKPV+shGDWGoXvoi92PoiNEGvN0lmtudGJUByMpBVR6B04Y4CI/4Yn
cDPkDi81XWju37/ZCTuDz6a7ODsYiOwUP2smtxXRZzFw3RtytBOUJoC4TCHZ/jll
I4heKcdTHsV6svjnOKN7NkdHAwABwMj8foqYOwHRSRcMaqHcom7HjltsiGAuKfUN
pFuws3pkASSM+HypefbtdL8qKXwaB1bqc0xjLIJyDIfDq/FUgVMu3JiFYr60oFgf
64A/eUAM5vvzwKZrI7l3rvF7iZKTB3X9x/REPlgG4PjS5dknCPA7yEygOrL73be2
gRIMalVypQ+E9IlP5JXvOO3th9cibKwtve61AwTRMzA4us8t0AlM1nUtM6pYMpSp
5zVFKnGuMZlK2a/3tixo4leZujMP7HV/qzkPNfjVEuOsuix80OcjWgEODEtsZogT
q2iZBdn/rtMkS9G/bLHLlcRTP7QTTZEdLkMqXTDxgYcIor8VD1wqC2r/YufJ+j+b
YXscQ60InkS104VHVtusn7eBmIu5Aw4MKjcRiqWLR+n+P9OPEw97ZoHBAFzVgq5V
edWNbaZCFe8ONERNn5aF6fpxmcAsqDJWxt02t+M+AVJK9P9KFucylB6fD+CZiV2I
I/5tQWn++PAEneA+HCsh5KYY0OlHlVLrk4wvzYcJF8n4PlIenZu8wbFu/BInBifL
2VWgOzltIVLQj4xT5zSikYrjNCOikTcdia8+ri2prwRsy3Kc+WW/NSScDRDAX8Kj
bKTNjMxmXeuxBMX5zfK5f1+CPJet1Jh1drRZAb8XkD5NN6pt9V9MTus/Ca3vXgjs
qVw6iBHyIy0qeH24olsoHluAOMhaJc7KFeVRp4q8B58vvkjC0kicY7J9m9w11Yfa
aprX25RYMia4LNmjtBrYGRzm7eP3wtH688ajuRGbW/jQnqvA9QYhfIevAzIR5f1E
y6KGu46DL5uUxRPZsH/2Vai6xw+Bb7UF+BPzuDwmP1H5B4V32QAak+kd2L/MEeW7
mxcdr5JtBJY1AglLzeSw83AQxgPLkivsglgFDIUnXsVTb45Hzv2HRIJ1ePTlgMkU
AM/Jc47Pj2tSeSQEkaJIwfTuL4sWN8d6Isz9LgrRZRu7D1Xmoj/b5eRb80Oo2F3f
vTG+qAq413oBy++YA7l8s9EIUWHjte6NifZkEWnZ/R/eGuZH2DNLm78J9VUIGXf2
ZcDtBfoOX09fCg4GAwQdJAIQbrOQgtNTd0QLQbCJnZWxAVlXUBo0X844CHIihZ33
BD7Yh5Ig242/e0gt1tufxnRhbDtqTaeFGmTaN2Q2pd5KKNVpA7PX0doTeOICMfMq
ffgzpQ6txWPBkgPf2e/ti5EKcVUEd9twAG48NoRtPkFoj05ndsEgtruiyLRMhW64
lK+kEtFwdMCOlTIeHVTRJIcrzQulwKo34wK4QbXr+4AFBoO4ohhWbsDbrPFN2eX3
luDu1m0dpM5KjFiE0szzdJQFvysDVs9whcXw1todTWO4utD9YIYi6FwxRLj4EO+H
dZz8yvVVqvSMcmWiZn/EhFN9My64oSa/W4fGdW9sFbhg8q5i+cqmjkFyMyP9G0dI
4vC0b9fXNnrGKr2Inh8qC2IClKLQuiuGEqLHn9TldbPeXiRJgJd6fHtZFLDsN7VI
TeoaXXXv4lR6ljMHS0fbulWUj/PIHMfpZUysPxP/67YixESfISN0XcvRTDC/i4bG
kCAI3i3iErjgiSAZDx9AA3q9UqRvn0GxaysP0FEE8iJhwBmDWWxWz0ChCCkLLT5u
o4K3vUhKEH/+x3TcnZKRbhlorz7wIGkZ0TtRi8s10zf6zydfF4nHelOqEmECnxZB
45GhwVsPEn6MqOdlu4UDp2xWuWBt3h820TTGLKjojJNzE9aRA2h+JYsizx3Zwaay
ig4Zg/VViVAj6u8wJdKo2UlxHlsd3z0vfrYDsSFl7YQuM5zfPExnIlo8sL+gFGGr
Vpa8QiENmFsJtabNl2xnoE85k9lcXmtbbG8F7zqYvduXr+S1S+x8ZwupVP9Ey7+e
QHygJ3DxUr17ydWMCtlPRzYAeo1da96Wc9O7JrrqFQXVK8PGTJ21P28sbftzejgL
f003hPy5ygVO9ARt3rg94SST2aG0lggZvM4nbQuZR0c4uzKN8DV/FRvxzlDRx/+9
Ar8zir1/OotuB5wyQUsVxuNO2oKJPsUo3V6N6DO6/ePvw1MDO/NSrxL2Xs2EzOT3
zjMEkChy6MVLHPT1KiZocaUBa0vpzuuZeFoAbznWb/DkvF+ZQ626VkspaECC+yPh
WvKL/v39HgBBomjqjT96/K+k9AQmRJOL9yBzIQZ/HdJLA0j14Y6C8UDgUL7XBzt3
Jl/cOtbu1ZVIhjjrVgNeg94CZn+qN+1fPgC8vphSgTHZmmxBKOeOkO639Pc2Kyv9
1ZYa9Zi1k10wrd/X51iSMTatuDRORviCCO23blHPNRCRsv9Gsi9UTO4IF08OOhch
UavVg55y4Aj3xLMLl7hR8GxoI6/S6RQvlhTnNTYXxp4L8jC8g3LfO8Gdlf1+3Noo
hVm7MAQf69cBkxat1RmxusuDjtatE5Dr8Jy92+ITEuiW3B5ezr3j21oNmfucuSSc
4xxn8eceTyQkj8pLc9rQ1TedDnBKKnkZmjnR32eIIpRTUsCohatKPAPW1Hi/toAi
p8pdNSHa9jSwx5t4linbqD0YVo0m9C+gK3uQVeZgZEKO89ZY1eIcZEF1hd5x2Qxm
g6azcmGb4bnkkge0UMt6pyhG7WTbvTsh6ixWCXFWwPxAsjHy7UqUwmz0bgH9S2DL
H4WfIu/K3AaBCelsx6NuNdnbS2Zg6E16bPxR1jm4BLDcVlNGd/HM3C3cwZKubRv6
Q55xCIseW2AjySa6TU+1cogCSofoY2XooxTr2loESxSkBxTUCQ3eNZIxBcWgmaUt
68fFal5SligrDwkQxRZYSGvgz1fsGEtg+fKq+ZNQuiIM5zk+QPqUkOAVWpNStHNl
kOhX1OR26/1LUp1jgNlrWonmuAXdJoZRblr8qwvTlYS10Jr0HtJO0+V3crgw8sqw
0fBlkayEezpfzSRHGgRdRFqQLw//Q6JkU+8qk+XcyYaqJy4GYoFgb/gC0G2uKyt3
kuA50P02OHuSkMjnU1zPgffrGR4bdQjVkopgpFfd8YWl168XdegYQasKSqZ+Sksz
O4fHoisSpmVmkUPPyaY2DKfR441cVVZWAjntqh2EsVC4SWVaXHAGxj0Z5iRtz75D
bnI6v53VrFrEMZkKjcg/liKmoxwXQ1VyLWtkIVjdvyyJQ8z1qkRuz8GDM9r++pxU
geXrzY99ptWK8AhESxsSdUkYGS4eJ0wLs0/PQ9vI+xC1LRH8kn2w7Mu4PqyXkQCr
2R0l2l4B1gznFt1lSmWF/xeHI5u6Fg1lTblUaxAjch6rivrQV2ebolVPEzSNBSHX
ADngF2NUyxDxTW4EiOrtef7O45kIBVhFwyM11FXF2tPN59nPOpS6xIR8LvekzpdV
BO35Nz9zcAM1l3fjgdww8dy/Iz84MVDwefMMcMoZT7khuOxuEWixq+ewiaUo05dB
lbOG+DFYnTJ9p6DtMRJmLvYIabjwZbS7TlTb22L8znYWLIgAZ0ni7KIjxx6zxVKY
qg84CPnH0j2FugvgydOOL0GtQ/enRrACkTuhg4YEoqmBXwq5Aio3rf4xvqIsBqxg
YFIanZHxKLlHx9+mVRoozGKYOL4sZQNEH8ePuGheWk666bL65SCaik2SPAm/DFNg
DojwtONYq9V+S9UZCC3SBYMXrTPWqU+GSTcipY9+U5Ykbi1xWImnuKGmYIMpGQWZ
iB0tBLw5sq4EFPuVtEqJWo6DF1upTpV3z1tfAilhOK/6i/62amp2Qp7K9Z1bDz5I
VX+ctT2nEKQnCTHpVPLuiy+1MR+KRo5ZqOFdaSddeJfOzoanGbn5V/QGQevaiKAY
KuxpiDR/2pUq4CpezowVsMhC6A7sJm6GcwtoCydf8N0r/DdDR5H05qmGp67MmvSB
uWjnJ87V/8ulCPqHHdYF4cTwoNiitBjvpok35LuBQYeNAxeQfMjNaPGSfkZBV0ZC
ytFQIwj9RZiGrk9HZV/kxFSsLIafEn9m6LtP3ojbSuH52MqePqySt4xYcag2vOhp
MMb+gXbS6DGtsJQfoz65gsqyIPz0ujeIKe9pLbQ68+HvEoLLOFzPH/z/WlUlOZnd
0ptLAdORJVKdH8ipi8Wn2T/8jaWEYLC0M5pgKqp8R3URkwoBHsZcobnb/W/AMjSP
MgaVeKSnK9tPI+FyFWt4rlex579GtdmclGT2odlS/R8pmW93gkbqkKq/AIX70lLZ
68aoQHDW49r8n8VW8UbNo/Apd6cOxjYnQLIdXIL0qJd/czrq4ubbz/c3PW9VECG7
6Y/mFDItH1MpzL+2ZgEwcL87lsDzoPybWChH5tIGIbx2HXiD2jF7yeeJfZwIJy/X
G9GppxnNruipmU065RpFDZRpvcOfizGIVB4G6YjYLSGqpBThDExfd9eWyl+65WXr
3ScCN4cXBGjwbUJjWjyIx0BMuCLeaU60TMAhEdF+fGmSZHRW6hk2icPSqFQ+2bBR
6l7CeZw2MxjHIWMsuAtaXP9NxRU+a82se4l3XOuIIFpC+GHCstPar2fZe/UVO2xQ
0uNhWkHYjEBkfJLWcEnLchEcBttUSOUTa3eik2ELWepNuc5EG5fPO/zJibjxF0+x
tXhAq/H5rFx2IUtsCf5gyBiCuaGCRN/42fApwmWYdeBxq3AJnIiMDhjVzrkoJGaR
Ur5BaAwSE9fyPpwxsy5djn/znMGYCX+bTesc0M6+JnkCWuMMkv+Rv/aaq8FBXvN7
m8w9kdEDqqm2SHKXHoz0qGdJ2Oi43NR7Ddq9/ykkmW/X+ILI+UYdRDrZzwbXjksf
QBTmV/8Fk63L25EoXeL3WUXNE/5ngSH449Rb1VO+D3XZH31Jd0p21yu6cPmysyfY
E+jcFU6xaOZ64xXnzr3NCCm18ONY6R9FyLtdhSHmbUtTCIxvbYUsg/cTgQKyXeFj
o4lDVPMS//f8l7dLF8jxi81tU4pSERFv+hvXICk323v0Q/J/SrPjC39QuB+1Rh/S
scO7SDRZQk2OT+myRhAV54kGr9HU7/mQ+wFszREe7vZd9PshT9tTEW/hwgO0TpLB
wN/toW7zwafbIR9b0AAM2ZVrawrA+5LrDOPc9Zlv2Svz+YRUFBpSuy2bKa2MGN6o
tlcegGfuPlAyriklOFcGoqCenLt2mds7GPDTyz03KYVoqVIuv8X8cZbdKKiqPatx
PprxV/C/f28q54HOEKTiSWRvirnijLMv7pGdNTAArzEb5IrD7dvtyaURhf3cHtmL
Re/gnxRFOQwLcT1ic0xzJubgDHPZ4anxsivyun/OPBeRYBi7ABzUH5iVDhXc8W4p
Q7HPbaZwUMUq9kkHufCWUwN1SutdqpDUr+b6Te3YezFHMv4rpFo6sTViPViGk6f0
zIGZRCN/XYxlxWs06PwMQLlhYuNVOMKcpyXXd2PAA6XYDgxCxXwP9PTDNTd3XAhI
44EOlC4d6ub2HOftrn08v/1jBQAF5ldwyhq3j2h4TJ99ZiuMRrrIGJTo1P0pgsQk
5gWaNsC1uqsE/kBYm9Wk0TlmN7IOSeZZtsXtBToQMCPOaF5xI3OYfrCI2KrTxnMr
oxF3+Pwns5KXZExPogk0l1ZRhKVESr73CJ0RnB7tAVSBv1HrNWWh0Zi3YGrgCgiO
Kk4TpjNbtIJ/5kjxERlCUEJmzmCWttwOSK77OHXBjZ9kRcOwuC5KCyVol07Y4PT2
2SRkZNProGzh/+DEOsOdYgUS74vb/QiYFn2cqWDwKX+IspG2LID2ikg6n1nxaqOZ
t3P6Z/vZoD+WtnCHj+SnKdE2to0uMJxlYw99p69mJkqkW3+ARJINtVqvyNLXwVBm
Vw8FQ+qw4Twcpc1tFUxYAdbUawNcfRPGQBkLj7TuxlN/AFu6DL7TwA43ivrAwcWI
V7oLRDB7Oz4x/njQ1jiyangEZpfaq+ndYNIOlRrMz1EySHGZndlR0IlX02kjBO0e
vC5YZ92tj48l0qXx4Ogu/oXE+ypEs1f2CKkGkELLyNQ2eo7vb424D1mhHEb501l6
eOA9eUSHD5ByYF1n7f74m6PTqUnH/wBieLaVHu/iWwh3zhmgrpm/C8GGB6ghjlDA
fns8RhYkevcG1l1U2rxBsXqmQBipqexhxG3KJa7xmenCiClHJVc+bqfshYbk5jhv
T3YuQfGJPOcXBwuGlVylEHfpE7WKYiBK2G/obEEaeq+f5BLw/2uB7AkYKJNjFcEP
ccKhvFZ5q7ms5MloJTHLDn7tWHW4fQtFeuY1YSdtmYWyDJVdgU+LCKfK3LewAUmM
VsVSZauED2D5VacSTc2eJS8J64x5uGUlmPusqCtm/8da53DJRuNmKzPnOE1LjtVI
29hRRTpnaiOKCs7Swh0MMQaiaZ8uqipYO9mV0Wa8GYRt9dkQsV/PwGgHktPySuVU
SyfxdQ0Q+qWIiycMK7NtqjJ+iWPz1pMb9fjuHmbaN90VVuxnFl1l2xrMW1XbXs2R
I9arHP3U2AoGQSssVUEXutnoGEismmxnbhyKJDUcBoIqdQ0ExYvVL+F8/Qg2YPFR
kKt1RBesS8X0R33c+H8JbH8D0cHenfHq3fOMfP6WQ5OI3TQSRLjJ8+JiMwEsvstx
y6ALXlG3+KIXsX9XGmIqXTsslDL0Sy8rQQPr9pJa/QzWVSrV6T1q3FbDO1kQ24xc
vY4o3bD9+49b9dHQW9CpUNQrnUQqQuMh6Sn4gigls4keNMz7LiSulbBkVK/Sa1MS
fgburjROSc02U2UxK+fLGMkkKOttCT/TCwz/Xvspek6xt0SXlG16bnr8jTODoiL7
x/eEq8x9kMC36+CuDAwrtfFuitYk8kunY/ygaSgty1T90jySyjeHOERt6PYXT4Wh
24DOfxmnTMsBCgcV42CkcMZdqPOhJo/IAjuUoRHJHLIMS1Pz3sW6VBFQz3GL0oaW
y6mPhQ88CQJt1p6rITRzBE40/ejqpA/e4Q33FEnb1A8dAmWCA52VtdXJrANspNVG
5eZbU6kCtuhCbHXrjBsez4QCuWCclPCTnh/JswwqDE1H4UZAE4oBN8Oi/8hz0b8x
QRuqzc9t4MFwXJW0co0QlFaycxn57PNxRhjaDsRKqje8eBb/ocesAdXBZu2BpYic
4BlFgzgHd++iyIBgK1ep3efHKAqI6wV76Nu1FE+SBzxjG3ue8LcMxwpTihhe7rkD
ucDQDuA3DkaUduJfcO9julJ6nlDHIEVMZbrEy+GwymuAwywXxsCFfZ/S0im1vLfQ
vRrNtRx1GdO2SQ3355tYz9hLwVQsluFOJ8tNUZhG4vL+FrwGJ6giwLSHPLb8mYHA
JaSuHucKoE4Jm3DFIqUUv821VNCatVCq4lfmy7uumrRFoIzss/WZR//DAGR5DAf4
ygHiTdVQ8f+TUcV8xSqNnzrublsOZw13SKPZOlt4HrGCHZxfqHT7OfkZhcB+8Jfo
gxRQGp5hGhTD/HYMtkAVblL9vDgVb/wse/JUzKKPb9SD7AJt3bt5ZxBl+UxIWjtV
unDa4RbhAO9YlkOoJWmeilY8LZrM3eQuHEaux+064765JjJPDXUggK5NxGTIC2Hb
lpp4cxXGLoLCaKcOUiZa32Ef3cfbOOOInjGdljVNbvhP44w02CvYwg0D6h7SxZaD
Tn08qwJ5rCs0TL6p6aNzvJb2/aJpLabifFlZOhHUSIYu9OZOTjlyrQpq0zgOZz5r
dLIcJaWoQ8h89sqmAB8MwHimd6eVvhJtK9Eli4oAEK7OTr8oT+FBm7NA3sj5HVup
B1h/3It8igOSpxM58GDqhMg0nJn2t65HVhgR0qSOeZtBEmN67ghImIkH/UbIpJj1
FSaT/LYn28ECDOnPDRXQBzTSbiKbosztjP8QcRuJkGDllvh2me4VSqV9xDQtfK63
Uwl7jofI2iWNsZTpDa28PKprmlk9ydNk+adm1Edc6Gj3As88XWmX5Fqg1SPO9D3E
EurAYVcXh8as8Qe2LcJcCnYalk8oH78XFT179B/rhfE43iJAv7rgGjQzV/aBtoJJ
gDjqmz99r1YYPTsTI3xxLFbW0eNCGkfCSROsiMdm5RrK53rX9fKLsF/wSbrljRIv
Dm9uXrCJYeIRwje1y+pFI4VIUx54v9oyi8HkyNFix/1DYMU1VZDhqmBN5TRGjrpS
FEN+NBMJs/KKq7BTpuohPL0W7/IMVCWPfdVDYg+tMGsdCd3ZIu04OvLHWRXWmWKD
9gvS5mgUkuWMfVWk5JAd2MkyigbHemm0buwyvvXCHYvXkdQP7VUWZaBpiMqgP82A
xttdISn20aQZCBzA15gE52ugXx1UKEYdNy2VjgpTqbbmub4H/uWwh60UNreW164d
D/jD8GsXe8G9gqdF/yj45VxM4RF0MEErDdLWFjN6Phq4DiCDb6PYx9C+YhEvmhYM
8vgxRNEmysM2i0Q7FYxEFn8VW+tLFHKYnB9pX+tnsvqTOCoIIENswU1Gs3VXq6L8
lyp2NQvy72plYGrfG23fG1gSBkvMSSGJYverwYPVWNwOUa7gZ7csScuWUyVz0TU9
UZv1bJknbZGgCrbo55gcFHxrbknJakIzP1p5NXRB9KkkCmXxM15UDf88TSRaUYR5
g5m5pWd1PL6ETRMoBPQuCnaMbpTTOv32LEOx7XKgkuNwxFqawlyZVEN0ec7gaZZ5
drWQ+JDWxYTykU3/eLqi5KPI3b1IB9/4hgsOUDLNC7A4pdeU1cAEhPZYTeHZLF2P
0t7pHmyorRIGHlHhPh9awmBoZ7Q1z5jgun4ENhoccw4FUUQwuvV4+kzsSZ5YZ6QJ
ljcNX1LFhS0vmLYyCLN9qr9mbiDfOniJsIDA+G0hM3G5z5YnI7m4r5e3P5n6L5II
nhkYeI49YBCA5r/ut0nxpbIN4ESm9qxPEZ42fYHJ3fSrwngaFNOsmNfSsQrdthSO
Ip+wzBzKiv5c7PXXCQPptYibQXqFrkC5BVLvgYXFXsbqfd2qhVIOEpYryGDXy3a4
6T76D7kVUQgHM+W77GjFUwjL42RJhncRNyhxWVi26l6iGgXHvvblDMljGLU9zmky
DKzk1E70g0HTslCf8KQK3fvA77/94yuOvTTv+G4JaJsPFyhEFHuiH8roXYWyO7Tk
ioXI6hGMHF5qZUxqgzPwsQqEs5iqM59YwDS6vVZtfi0/2v/QYYbgzPhJJYD7pSzO
kazA9EClBMQVvdcXA90yJG0fRgmXv9BMdWBazmTAQxdJ03A5EuxJyU8uns0/Oisp
o23tbVcbbnOJRNR2kPo1dNAibgnyLokPSSQEBgmrfUTsVIMSuZDzJM5gr3NvvaUo
D7yJGmuC10cUMwT0BA6RMlbwXlOPnRng4PAu6bkHTSzO1/ASbq6WLAtUJroOlrgA
F02XLDFsKRjYT5EEoaq+HkpU3DpFeGKBnjoGIz47RwI+xnasKSkFn2B3jRicuRUP
E628WOfUyHcXwe6QbKA5NDEhxCaMfIAdp76o6gSdu30MFSBwMe/sDSvLMA1njllK
fR1oKnzZ/EQ9Xm/cWd/JWTA2+0RLgvfupcAhvj/HYdrwZ8cAXt9bZbAe7DO6vuD0
+kuWpZLlwTbVInMCtNv8dG5CQqMSpsUGtLj12tUkIY1CzmuzWDyg7jjyOa7E2tWc
w+b3qzdQmr50L8iJn+YsNJktgIWv0p93vZVow6Hvmvhw16AeaJ5lAMHM2jrMk2V6
Pu4Bz5EzVBNwyAwjpykxNwBT2aTXKudjIygwXEFwOLXaZtBjtrt+L9zDw1JJ3dyk
OHdQKZYmKzJUEz3Vl8tnk9VN7JbqXbZc+vyj9lyILhH0nweydDJ2b5lKMiNrt/ei
UVkyrv1iqDR3Z+98+mQ7PiwEGLzHJsbFZ24FREf7LJ2tqEFNH+F78pr25iKoquzi
RQVsAObKgT1Kzjf6P0A3xWCHSaBGFUXTnLKRdjtlj7VPlSpWTRTUsa+Zg6pWazZp
QnHhdskEIjvCIvFnmSFwJ7T4LjWpvmYyAs+FUaxR4n3cAAeikvuCf56qZ3tGlEYO
tKKfg16dGpcsyIIxhVSwWePvwgkBQ92b9jul0+Wbhkh9WKv5X7WjvSBMoV55psCA
ua32CP8nCDq5cu4Zlm7fNY691jpcUOBKnsUky5O1a/G8fiRzyobQR01g0M0aCHZh
Lt0sCsLZIdBMA7eHoBXghM3vu/5wkcskPGa9jyTFNcaEbdlbClPOv/ktqPmRYxRM
ZWUCSZ8uDtXt8GuWhQ2u3ex4euJmrZVHzZYSBQsyt97K3sp9T1cBjLVht/Uj80/v
XSTh14v3uj+Jkv4/Pn1AZYpVNV91WCGRVv+DiyQDJqjHafiY17wEaTo85dof18/S
89k1BWHRGAh3KxKq+obNBOyMvFAnpxkbWS8Mk0o0iJuA3bnwtbtXuGpr9d6YUwTf
87oAaWkbn7GJp0kjdXt4qU/pOoLl/8XD31lKNLWSWregH2U2geoKFwUArUSFsYRq
A2It2LMXY3SiSGOjjrM08jgreezBZRoG1AljeOPrBbk3UE3oWhvXdFKgP7ID/6DV
j6rh6AP5i8JEuPKajTLohEnmpIARVfbjF7IfzZceU0AzWp2dVlI/O4x2KHhA0DQK
XwvmpheX1b/P/Of1wy6LWqjss5ysu8U6wU3wARbpA7PenshKCPbnLnLCZtpZsLdk
tKhaPVI/neX98NNz0zrBA/K/n0jynnC19ZFRqSDb6bIgu0CfrVaipVGq5tm9rI5r
62pkXQ55WtfR2QR3U5k9V5lJKFsWTYdKJnSbzgISJRUd4TcKOuQFFVegeL1qRbEQ
kyU6Ep5nQ6SETCTcsD0dZKaLf6Fnajz5C/G+gDxNwZErJ7jsd6oveJMKb8YQ4EhZ
BEWSP1LIpTbRqq/NfNm19Z1uAHc88Urc5Z2eBeG9iPyO5NIruoXqBmIEZCERDUtK
JopvwpL/a0d0fCUqRFQFeLLiFxUh8IV05//rHb14Sz1PsP92hlSf8SNGnYpmQ8mq
SrHWeDRskGk18RfA7/6mRSFE8njKlEQi2ihtCj43ex8bS/VdOdViM/AJJnl55mRt
xAZiNnXi+7pvXrnEKmW05LtId8nY7rb3yUU9UKhFrVqC+X5efAjxYtn+cMt0AMel
4KgLpKKFjhqD/Xj3EQwEryDwMwbIvxnF1QXjxpbTujhaYHr3u7vHFwv5SABJugvg
y8gA6nTd6IJ0LehlxydJtBnc36mxam9k50wusP9Cb+OHEDx/zWocdsn6vtmFav40
e9gT6xGhusvc0uCO1BtmQjL+p2a0pL61/1Pws49HaWGz3/UgpEKowhG7TApP+uE9
zjrSQVV0mIkvmnWPe8b6fxTQdUUHYehjXnq5uMxEyIYNzmz9rxYa3l0UTTuT/tiF
F58FEH/DKeDcXfe0NYT4S8NpOzS/5UqVCjqsxBzP/xWhd/b6leXasoajPy67JJ1W
2aIhVJAh1lgQ4FsiCehmYfi3wA4jssKbcxnZSuI3DP7eZze/arJZKXxlR9CtqnJU
nqUdJjfmgYaHrYfJ7AzpLbgQA5H1msqQKojrAq8Qk8sV4su+GGbB7LTSTDnfShGN
Omu/sDAwDXUf4h+98V/3pddNhLbWN/OltOaLTQUGKLUGokvMFu3ZVElu4hupSUvt
kDs4P35gK/NKWbaP/j1R2UneAnn9tbMOPVCTPYvdGyIs3eanqG7ovQsGAKI2Cg1Y
nDE9fn7GpEp4Uk3sVLwFmwI2K7KgMJUw78hvnma1zgCd7bERG80gBspPljq4DVYM
q4DH/U9Sg0U5d8SetrFrZKhHeW608CsnVQKlICHkOsoVqx7BynfiaiKwBkwICluG
oPtJPy8FdSf4zSZGiqNGOSepANjSjUZC2Q+3HUApuBh+Ba8NoHCgeHethP/SvE/J
b1dduAZg8qvOWx36Pmcz4MrITXPJPq2i4T+9hlSwsKVOK7iouyjGiIuXxq1X5ZOi
3Iz1ZtooBNYtTcnfdH+ou6bmhnmApn6ZieWUFTV9O2tJnTVpu36IZQDV2lu9psqd
gFcCpeDoxcTVCVsHZD50fKipDg7hORQSvuCt9BhnlXa8cDafz27RlLOG3DO/h8+4
ES5lqJiOvnKlOPIdeppMhK59lfxMzqCnUtOW8RpJwl2IXVzTcftUP+M0Lu9FOuhI
sJ7EAnjToqlpWxDbJTIHczmdEXeNQmdzBBhIYiN/79772upQUoMmwYblOIVdzzCy
YWeRcAYSTF/JqOGZ+sEB/LUYxS6vc27vxAepSrHL1+rKl89ZSfismOIsZ4Lx4Pir
J9a0mrvCSYkrG6ObhgTEDCygDrkQRXLQ0QWlaoRR8OApy59QXCOePnbpfg11vLIP
kSpgNKSlEWy0t3a/FHQ5KE+Z78i7CpdmSNAOaaITCl13ljD7bZVuA203cgSSNGcV
NrvFzEKaV8Z8zMulDojc+5Cz5/L9pnG9gtjmUJKzcT0n6Ty6cbuXym1gIHrE7Ncp
D5txR+ZGGXj1Mv9C6USy2NPlg1JJ1xK0jzzTbmSh/2h/fxcnVDOuSEi4q03AP4DZ
ITS4ZlktuR8V1AJe6vKxm6WHKe1A00BlMJEXSiXkVaszCR/x4Jbz0e4j/AKdAhX+
jBH23bRYZxilUIu4DMxBb/nz0eHJeu9k+aPiWfa3yS1VtTKr0DrMC6rK5YLnc/2m
JzlbLl93ersOkJqLbCyNsxD3rbSGdhgpady3zPgYWCvklEW6mqKEyNKehKJbyugw
Np/x12HMTEh7uX9mvGR0Qqxov9arzOSdzRujQ8rnh6J8CoRbJRP0fTOluMZQWKtF
tDTy0vBk8EWeWIkMrS7uuFexZln3wle++mBDRGJ/qqoGuN1/ySbRsZiud8+mYrgc
leaNoDALTMVetnMVhbGoRzBZc5R7kzu21caGfXbyh97CVwQXkcOPUV6kWaAb8p8P
7wzKLzwO/rMKaSiP9AWl1a3ZZc+jPB8vUWtguzv+nXxuQJKKSg6/rGFQBLYB2T86
0MPeSLry5Q0Ek073OImWImvN99fWl5KOM6CbLhil2/Uj/uLs+BKbh5U12j+1ke1K
whBHCqJuOqFyVACkGiwmqVfvK5CBjVx69IMxblhrPcjrCNTvxUZasWj0Q996aid5
V4QnYpg9DtA9By5obJmHzo6eONyXhmHMgrHA7A7kn7Vb2Pgsjz+FI9pkVZ9m3qs3
YOATireb/GwV/ai+wP/KXPtB3gx5KpsB74m6yOdsIwa2Yh8h2iKZ9tOoXXh25M+P
wbO/TRE5Cyo4Ssfk2R+5odEEx3kP7U/9xwMSbZXx1s14pmiWXJl4QdnH5uNgjF7n
2nyX6hotMf7buQJsAS4LJzn6EPe6KAM7k3p8c6D6X7oV7QwUDoQrCWIpS3XgpFPv
XDVSzWDF1PTf3zG9vejSqhzmmSvYWJAtYHSOGMHYBfWqZAUmjpSVQGpiD6/lOwUv
5Rc5J6NpNkWfx3A1/EvYHbbaY82IFgbJmrKl9P6V93B2W1njSzhwU6J7Pu20V2/z
CJwIEcnH+86/ONrAFec413VkjK3EYWSVvrHC975MWkXc79z1OGyA49gtUOFZfVxC
CGnaeAzIGM0dfxc1UO2HiNFUwMIGfPTdteXEUqyRbkU+LwYrHXzfEUNX7H/Z4wR/
f7wxQ9tn/E1HSeeL6yUx/cGz+eeIgUT3N2kL1x7kdO/Mu5gYDYGFLOH4uzgVl7r2
cMFiy/4iOyCYeF8TOyTPGo45328i4UJ1PlA6A1ttLIgCGEQDbh4NJ8bgyWmtC+Xi
NL/SE5C1LGIz6epUqUd8AhqOqfmRfuMbno9duvaWu8adqKsd9xxxOqGgplqBp59O
k9ADT/q9fFi6DQ5OybwlkpWMp/hWQwwth6xfDaFlOdZo+oKY8Q0oDNS+tzYFZJOI
+vbR0ezmCg/i8WVKJarN0WUPqW2HraF8b2hweZTC/pZinjkUFAVPsxgrVpnT1RtZ
2SkVDANiPFkR7pQ22rNAtASw4yxoS85xs6n4v2iqqFVG/Z9HHNlLjsbL0/1J0m/G
OSTrtcQ5WLTjbgdEASGB0XJJ5rymDdVIseZe12NdPAq3sMvCVV/TfFrt/0VrtqMd
JNyyqv/91n+pm7Rv/3TmUToj9s0xz9K0CNOkRtnwVCBDbNRvb4VynGBcPid0tMf5
qpy0pn/AgIRYPMqhmarrz+hWmUrlaBKICSpLAPBGhWQEba7uS5Tj/v1WbGvIkY2K
Uc3RNPTj8v1dT3ukOOp1Yn7xcW4sRcZOiCNvWSvuWWn6XjiV5fAAgYK3lPwx6NEs
cNgwx3FTmvPwHJo37NccEcecrVOLMZ8xapmX5AeAEjQ7L1RS4eEHxt/E197GAb2B
pm8Hzh+dRTa2AN1/FAFvkCkmwulDPD7UmGICZMi7C8aIiQ5zEkpKUeLVRr4pKGCh
ti9SJjvc1dlvpbYlrLRPvjCjaGIXT6ZDNjyJsINMUDu+WvU13+oIcM40kRnJqMDE
BT0CiEQzo6JsJC6cSgRSZ/0twEOI5tj8JZoG5Vc9ch1LfQGJEB+4vDbi/feoJdUJ
VSKVRGNZGWgkBo6L9HhqKhZnOHH4qJS2XnemzoaixCeLOSQHOv3AGrf+40Efe+aN
1rvFUwNTB1JuNjn8rURowM7VttFUYXWPrSl5L5yG9vyCfow2rZvnl1bHJYimk6jE
u+Nx3i3mBrXK5SRKsu9UnEGpDPZUKAt6/xICIGUOAAXci7TSl88kH3UjWltv49Ah
DcNErDCzfrloDy1YSuKNnxMVpJ8RGR/6MTJ/BMqPeUt3X5cJfND76IoeJ6qgNqID
LV4fc6zVnAs8Xf/NONCKTSbvcCD6piMOHaFzGzr/0bhxZQBY0iAYRcErjiODlwW0
VYgaZMNMYX6fQH9/jfRDrn6YZJsPYub4Nqt5jR2C0pyAcdjNpwrtuijISnz9MB+C
bVRwmNyquktSoX7nJ42iKxgQauVsat0CVy0BEKO1S8yJMFAI6P++oe4k/h9ATqrT
foMMjtvxLSdHmC2qFr/NfaUiVw6DF3eDnB/QRn7hONequPoD1VEcFV/c1Gpr7NBD
tWy6yQMXmVjF8kFuL/xBM5UjOztTfXpC1HClvzPnV0rcAb500ulzbQYrBc6aJY1K
/R7Wf/5kaZ7VaIFCkxGTArshEtU5CC2WKFGmU29vC01DIgUWDXxkMTBcuQE3rBwH
0fpVaStTDj8T+R8ho6JaJzhb1uHlWSVz4Zp8D64D+xjtMYoV7iQF0S+WcDQxHLh6
WpoQIRWCwyFd9AeD37tTtiT+UHYeCiVAK4AU+kNVnoOfy3hVzazL3zX1ycCXNLeJ
58CImjmUHGxL7FIOtCq/5JBZX1uUs9MjB41nntpgYjLWFj66X6LOwtw7VIhT9GZe
Rcw9PlXM9N6A6UNGb5cycWTeT2jG/Wp//lYrvUSfMFIYH5p0f6BnG8n8+hvQpiLM
27sLQlap61G7e+69upiDOKv0VOpaqdHpF7JpgC9oS1yaJWeTuoIlzshFePjtkwo8
rv0h2UBL+m9HhBYwFWtFkUDAXPcBrixDdrlyyLWuTvrK8fG59kw9oQlLSSOjDZF6
7V5AdX4cq2brmjvYhITUA3Z6Eo1nSi64EPOcP8S/TSytZH/d0G9leWNRP6R90QMe
FhSvNu9vXrgVZS9uqKhr519ji+TIig4xb7KTzX5t6cgRBer6zISok3j/ef9y+4JB
oB2izKTZVBsRGcaQ2afoMvRH6A9DdYvqVbsLzJH9yJGEMOwEW1czM+Cu2/x/8GU7
t3ZdJmYP0CY7XNoWSCVMhVnJIz81Q5dyo/yV2bY6R5mqkQgFfdwz32+A8G20ctly
DiqiCGxCuKD767CmpWxWPmPHPlGd7rWd53dWsUluN6tIjlZyl7gaVKhgQkYHu1vR
OpnKlT/x60Qvvwd7EKqLhFhAXj+E5JfDT0fDD0RG+UXNZD5WbcOfLkIyCsplysDv
D5o8fOR9sWnWM0HZwnvpcqAZ2u4xZL1OpJ5stloi3dC/TPiB1cEktqHb6gyJXUYA
j7rQacGRqq2maSEflrB4F0QdtAqkxgQsTLT91rUaTtJHPuBKyj17xTLkj1GP3MSH
2Kec6VUkldyig2u8iL+DYjuZFDiYU039vJ7Ch5m9jDflZ2GKu5H7nQwPnqfgIICZ
5VP6bjuLSLzrSeYaJbN5rnsuBIMQXhc6kX1sAex/lFRD3yXbpDtK+5GEvJvqxzDe
0nCkRu30JN3yUfKFNngy6B9m6zpZ/10sCyQmtTcpAlpT0G6znKJOy3H1JiAvln13
KnKvJwgPv6vEYZlWpnXZS7xf+dx/a70Htf8adoYxD7fV5zRFk/+lBhitWpxAlcia
46P/1MR8YmrMme2VbVNir6T+6J00FrcPZVupMc34OGqqESplSFKcoYZgeLDKfapu
HEweoP3OjkLvkiQkcyJ+owXAU9NR9U2Dl5OvLcSbvAKTFzPkwHWe31OEvVs5bZZ7
7uogseijY3ukPWOm/XYJDolE4O0vHvotagSLee1jMO4bG2ij3pkyeOQLZtEHpL2a
+gwuESkMf4cS7OfPWmqMNPTRN/+23XmeJ113AvpCstNoCmF89oXQe3q8bznMjt5u
4JRSG3wXyPTHfcazqIvKGCgFfSZQ04wxsGr1gZTIrLR2uF5QrlpJH3IxQ427ReIl
I5x3uA8yTY1WORpV8cGRvLtPCf3cRzgkeyjbCCPadMQKBQOnWrNwrnS1l7NxjtLC
CzYvVWHb701cil/z9ElkrP0b5pAmbZw2nM06xAPJVoViHWji6PfZJszLyyYJLOPM
EQA2YOws49RVtT9sTQ9B2DxiPMlAPmGP0ttPR9HybK5bn37Cdgd55QCDgf1+3J3p
DGeVOHEukpUooIP1mHwVpmZtCCq+qEdIaxFuTAvyJKR7nLadeKTUafIZ+YzcfgMU
LiPwU2+05y+Vu/bS3XzgXKdXy1weWHp1kx9zwZf5t4h8cTFE+vW4X/enEAet/Fxg
jiFjrHMHM3V0l2wW1DHFHEykiydHr4ok9AFYBAl7jJH6YH38DyXUO7mwFPWOHgQ6
lnus677heAsbwNA62EvecOZiG6X8ceJ7/w8h7q1go8w30HE3FqrFiZCWxP1q0LqU
A+HX2dq/tBSmHOx+ISKt8qUQ1LEbQ582FVMzAdFmDpR4WKofWiQm9nimlOgosYSZ
FAPN259IL4gfSWAF/CfbU0Tw4nUkONxRLbAP2CmGSehruKcXnso6Ndb2fB62EyYY
K5RL0VPMNZnGQT1KZ55aAhs6nxgg/hU+wXkCDlfhYBEyTQFc27PxudVE1+uUv4KC
2FPZqoyR28V7mhJ/v4HrM2Ppq+e/M7WYAKLwzgjX6+YsL4Jtz9A3LwSSo6DOFmpQ
yxKGXK7FSsnd3KcOwqAw0qV5B0AAkP3oE9HjqOk+CBLkUHM1xJXR9WNTdic/fgPg
DQ56TLc9pIT7V167XOrC/ygwJMONljpxpWPCuSyjXFJWK0FNqMNzhbvwf4hlaNq6
5FFoazperHHMWG5XuOkEzdEGZ/a+sdG+U/4Niq9p5KaCoo6ck85GdBQ0KV1PmiOq
4XviuPejxyaBWvmkg0wZklH7Bw+5ctCe1vpTcetDmbXBQqn50FwDLD0jdYEUgkvC
9kXiAyhfaTj+4sfcCGXraVYJWUcJ+8V2KFxVqE+HoByL5onVlyEkdG034Rsnr3yf
I5kG0av6WhbuA7mBcv4Jqt7/djgwskqq/hgGLlwGHkEq4GQMl3v2m2NZqMqxE3gM
N+T9cQmaJJhMIq93I9BUlU+cKV65iOPkv9FhFUClSZJaDN4AI14m1f4w4ImZZYmt
oT3jcoEt0hNwLNUGnzjeqbwB1cBkfLFOEY9l9ap7mv7aibHjGBQzZX4HICNDv7LE
r+VexSWJObg/Ys2ILCnwxzc+d2mci9QLIVPyCbNdFlLdhbkdOXzMvVp7H9UwT2Hg
9A88iP12QkrPym2eJIt17vv/zYL/qg0XKVQa3zCWv+goXhxkIok5vzPBE+dTA7Pk
rrh9VhxlWnB8uWbYKFpXYN8/6gXhluB1tLAdeHYPc2rta6Gc3grP+3yRAV2iaUeM
tjufUKtZN3KL/ZS4v3BRTr/9bWQFdIlQLwTkZ51zA1MZOIOkKpZb+km3Y7vT6sow
lmObc0vdMDPq4WtbYbmqwTFtTFg6sai3Vfi26mf42Ko5IRx6P7oLqp/A4ecTREQS
3y/SVtlp9vQCicfEUJLBZzawB+zWMf/qucB/opEOXiMckZJRPz9XJjDpTGNnTIt7
V3Rr5b4TgUOtrJRakWpsGxtl3UMxjS0Us0+KDYe13P25eOU9bepR6eEkHdC9W+Sa
qDjstgYPLpjoAXd2au4Tzm4vCrDWAhVcdIB17QOq18AKRhRSWY6XOwTWO+Qxl2eh
YId473ZIrr31EFQ9aSlF223IsHC07qCVLPiQ1IyYahowJMOTbL3agvBr7PlohbRG
k5U9f1HgIC3AIBLF8HXs3f5MnikmnqtyDeABRMP4P405Ps5ayl08StjgGRdljCeN
ObElbFqAzTXwrg9B+pCCMJFhTH9JG/l2mk5085ZWge+ROI2B3XO13kaZ+uLn6SAO
lj+2JG41+MxDUaCn1oPGQIL5jk0hF4M1xztTMXlsxBIfEirX3TmrssX+QT+mcElT
BEgAnu3tVm8nXNta2m2e7qKMD7utvYe7+XHNlr8O5AYb+y2HAEtZNa63s+I6HHAf
CPLYRxevNH/OWgKxiTYJqvH3gQlPHZoo7n0SOuIEs09NZZTP2iQ7kWqcoAVT9ACJ
PNaIsEcnzuoNlODDDa//Ht1Pr/wa9LPATv+86ehHF69jwiKdSslaUR+ikJcK1Z8x
6C2jPfCXuOSCeYPd/654qvNSkGH5CZG7AMZrIsUAtE2sYl/ZNL/tjZa4kR/9cuBN
zHFwew5vHNnSg1V5Axy+MlRwmK4XvIjb8mT6I87XRTaucB88p9stbbnUvJ4DwmpX
MNE6+RKYBgtPs+lf+TNeY8QnoCPj3Gpop9AokH4Ya29H5kFYne8gg7kunrUDLmLH
bVQGnZ/a6Eg0Q5mgyH2rVRvrXdgaJlKKjPp+T1Z4SD8BoJPynKyFPdbzzgccTVGJ
gkITb9vO1LVvENizHnkb/pEcjnJ205TECmTX6nKGPcGPbcqUhBooYL337qGv2TqM
gwm4Abet61lLcw0G40ssGH1eLSspN+3zkUcN3BGgh1PNwPWkDgAxSvFgtTG4K9ag
2J0Kg+X0E906N/8tlw/lFXFxmjdOrHmR5i36GIDw5CrPuMgzhsUoKxeL7bvsuu2p
jnVSnrn+Pfpq7Fy6iTWoMeDhvymr3ocVJUNKnfO2utns3brBwbNUpcDAd3awJePc
1n51af6AYyoEYY1n8UTAyZfuS9HPcun0KmQ8d2Jrp5nxI4N8wwHApiV9BwyKUAGO
3GnOFaIJxopjakMKNQyx8AG9ocHfRC0DJIHAjG4WaUGh+WCZVR2U5zQmJrAQ38O1
473tsphGzCJ8QDB0uDzElyxyMsutLBsZL7JjBHuzaHGqKaY4qunLPQawHOiPXDup
AjnRh7Sibvx3Z8yxvTxfbtdosaA6fbS9h18xfEK8y21BuBUH6XdjVyp1Kyn+Wjkx
iCYkdymyl+oedAW3Q0jzZlZKJ6A99EK58b+kJxqkRAUb6rl9rg1IpZKueLqquMDL
D4yMvRBz9xjacADmySpe4wI5ke+uNsLY1q0Z5R/YIzS1M2kouxrxprjCS3kloAKY
764gP04jNRz12z3Jq2jMJ9BSgP6m7dE3/9sQsqKBIZF4BU3ifyB2Vup0gogmnv/Y
6Xr+Ta5+qpSIwCBpHARKm7rp9jEMPqbIZoTvgM4HmuSyt0iOZtXaE4rK0GidpH8W
XsfXlTnbmCwlfVXJivtkrUy3eQfCNlqfzv9hqtFiTii1a1P1z6OgB50etzRracU3
levzlKh70nkOdBBmas0QGJyrBWFln/QfgoYB8zfTSxHL8BW2Yx+I2ZzYVZtBcFyt
Wkd+13ijeUUwR/HgI6cs/HGO2bzpaJKJJzD5PYNfnwk/3WN5AdxttIk2DJszymg0
wGMLy2Wq8anskO4Un1LiUCIotMie5E2ncGsCJG34RtKDp+oHrcrQI5h39qUpeGvA
Aeba/4Eki2FsqDBhtAqUZcPgaE7RwA1Mc+OGwDsyuEDAWD/bpYe+oNAmUkYJZ6MM
Z2ezNixD1pKlnsnh4aSHRFJBYpighlrhWP6VEIHViSd1vIjsA50j271RZMoPsDRl
PJblIO0kxlkITzukz+QVoC/KWByay3kW73l9yiz/+lAhFKk4d0gBuTPVyEcekNPm
rXIiDx+UxdCzyI3JNXZmeqwPsq3IlzCADa3Q6PjrzaNV+Ux8EjY3SnbnEFfVeO2w
0pfIjPKnyvY0FKCtMayk3EvAyHVe78/FDSHLpQ0uOeLRZOJlB5n0KGoWTvAw/CoI
zPqLdOW6AkyRGaKjz7sXxuP5xSpAK6o5TnyAD95bgg/jMLxmDuXpL2NsFjdEWzXK
/sgw8VFhJ4QWrqXTkUxcnkAS5LiZiNMExpU8c1hrs90lm7B9OVRl5dl3/qYNNxrz
fr1y2m5kAkgSEX0gNdqI9Op9Ml4fdUbCxbisLcCbim+CGZmzMXYQSVfvyEdmkgq3
OQqR6om0hjhpG9Qwqp3DNjlYWAc+98nMQMURt0DeAmw8DhFBV43hCDEV1gLvlsvy
UV0VkiqaDSwshUksbG23UH8H3Xiys9I7LWh32B8nkf8WIi7p0b4jRT4uzN9ouom3
3f6Gyc0G2gnl/AE1MoRwm11FXUbO5o8rsMYvFooe3L+w1sy83Me0d6mXMmNa7j+c
cKBc+fqVo/Az6kO4RmE4bBa3wWts6xk10RsASIsKYwBUn2EVAHWpOVkWDQUy77nQ
4NlCHQeLVUuquXUwSpyuQ6RUQ3lO4QHFszlGGNjxMEuHCNpDBgIl0Ma2+w4Uc4V/
1UQl/K/IRDYNOFtnzSXoqhPbjU9a3PrFEewMK+fvrcHADUa6ox3ZfV101bKClngy
F/p0SDpcFbaNaEk5ndldZvc3/xwD0OlKFdmsmmpKdir/nZKMLBqMwsltyr9Ch09U
EMkV0B+YvoP5kXkk3n6rxUyQ+Yr+dO0BNxyb546P1Cg1ZzLOVtA17AM4F4HQpwOc
7nnwpiwnq8L2F0k4B1sAqp9Y95n6oeoWJHxet5qCjDCwf3kRH4j7XctlSPI35AD1
PpLl9LT0hx5bx+LCQP8qB5pIvIPG5FUXjwcCyFSQnYi4IxX4fX5S9OwXpElhbEIJ
gSZruoQL9efB3A3smIFCeA0noOoqceZUTNaOfnB3B8KyCE2jZoYwupV9NEzZfYMv
XOMFpFPLcXnXHJ3hVc2nE1RK4qMSDr1Jy4kok98WL6zRa3ZHr7pnfLKUWElq40vY
ETF2LF9U8KnrULBrdXzbT7GHYNWgCq0ELjVw+pELLan/Yf5K2w9zwmix/ek2/toI
d0eT8T35Xwo8UQpGVxGU8i0Z6BSE6STB5HTgNrcVIpqq4ftPjb7sM1pwVBSyeIcr
+htHFgjsW2r+4kfvooz9jdbQJoq7Bw/zyD3o3ixLL/4rJYfASYjbErdFndNgiNez
VOr2cFcVFHCx2IfpOkesuQWdCdrGUvqoouw/v3/D893rJZc3p9NY0haVzXbVVdTR
DsV7MCEpZszgGvlCMEoz5LEhxi5CUu89Red7mWiuW5EJAxCbGXZirYTaxEC8rGp+
QUGg7F7kQAemdzD6BSvhJwVvnPFSipzfv6yyPXMFgKv2++/d3Gru1ZDgZu9QobMS
S805hKm7UaB3E45YQ35JmG3nZ7gdXqIzVz6az7QQ+XdAowiMq1aek4WDWQW5+MmO
CluwPvM0IKSmDFoDljRh/1uQVnCgeuyZ2Uvy0ToWgcJ2VoSELm9TePQtFpFABi5r
gFCYoB9HP7gG6iKHbdghmyZIiNC47lqcv8s1kzoF0fpiBST+O+uahp6vjxO2tUHL
5ZVTuRs6ZqVW6wNx5K0LfnSil80DVl119U5VZLmUAylFReGuegFP85Wt/X4nNaY8
Bm6qCxauyLLSg1idAXG+LSvpleQFEJbMYb+Lj8oa8hwbNOowOxfpTdpLfbHPTrKX
sTd6SpidX7zQshw4fKvk2jBcLHJQGdhwEPiAed5spSWCn6pomYA3K9iv9ChOktgJ
6UPlVDTSZg/cjPiBB3FQe8cl+pVwYojYXVY3OZxVEG6CIG3QZkqT6a7hRIRH98FC
YO4PgStuXki/oUk91myXQ0lTnFdoDUkFBgLowSupDLdIB6dQTl35pEvaCQguiEmW
amoR+VOYhIk9pOtn0ne6/GSKToQUbO5dh3pJz6o3R2thw5F/nTadDvwi/4DoWTG9
53SfYkp+cnux0vCji1nTpMZ3Svb2MhokDoLdPuZbaH7eGe/krEXZO3iwAh6jp8z2
abdBpth7IcykX7xjeRS6EFHjhVf9zrqYDu2OZJ1gDoinrvdeJ/2D/jmqTx9maoQp
Y3ZvTwqTB73axTL2bv0i76kkRrJPXfqWz/rRjoDl5zYSNSjyAfgKBGGr9VFPeeHl
LEnX7vhfOYgFBgmzJZgHnlxphE8ASY+sOUktuOxqSeWECpOzxl6kZjprT2ZzOthB
6FMcrW7XFkKh0GQok6p7wyas+GuvRX0Al9l1hwcY/ThEzMWSa64hTMqvhUxo4J2A
0Kau/eQBNvBeGoUdjUARPSRF1OSoCFZPD4juYTGG114Ll4m9y8HFo8VviIJzf7Ca
AxM9I+Yy9LR/pct/UL1pY01NAUGyYtj8xPQ1AU6049KfGYprikElXv0kKmQ1SSYi
IfEyxdDFXSGjJjK4JyD/Keyfshti2H4+y7Hcpr0kg6h8ZLcjFrjfgZSYukH/QrUC
0J0ePzsjkphW/BA1DcIW1RfJJfQf3BO0lrYzq4rQ0NzY1myvKY2NP7HWOcltpXnF
MURSi6J/77o7iUwLoy+FK//nt5KAj2inMVSDjRDWbJalLZ9kPfjfE8fn07fKHx8z
RX/Bub17kRCMl0LgxZHup5sYSBL5OiiM8HRZi9VYxuhUAz2+srLvzgGKoFsx/da5
AhS7+cBCZmRAV3SoNjvQQMSSOvLFvZU/sN5WBTw17lSr0Q0+DSYqKKcz0X7wWmcH
e5DasBgx4+HMhNXrMKxZZADUMPvBLsf87boUPDqiAU3s7kU07JWy9A9xc5j3bMbM
ZgYfoiXf8PytyBi8GqHf+YTiXxQS4kx56MaYg98SwLEuJX+WHLhmKoJ8VBXCEtT2
4zo5KCNgJ2gC8R3Lma51aJLnffMld7esBr3Y8NFFDWeyev3vMl+y6TjCGMFIwT8m
VfELsRDyuQoX73RamWs7wSSm2rDN/7AnKzFyQIlMWw8fdG9fOuFN3nYrQStOjVgi
e0n66TfTNFI0bL1oRCexZVjJUP84Q8cJ7x6G5ef48xEV71I988JH5bzAUrm+vKEb
3NSKxliL3KgWc25NdZBBoZB5wUQA7jwVrYGKrz2GNxvFCOlSwkR6T9lCxS83Ovb0
r7Kme8T/eFaRaypUSbhNR99xlkVVGT8uUwIFy/5OAyauSCGrlYNy5s3YsobTPRf/
nqESDiJ4cO6bZCL4msr8UEyOyfwTWAhajjRJ9ouxDUw6GsUByOfRmnpZ3wKriWcG
SvF2AmHOB8BXRXnnObmVG1Fakkr1MaoloAllrhEUo/97GaAhW0HWurVlkWovkezg
JgpgQlc4NwssOU2Yp8yFCdthzQpJB78jiizQvGZw1HxJcqc1rX8sNgNV3Y+GuAS7
MdyJeEmhg+KMNy64GjmT3gF7CLLLJTyJ5Yr8fm6rtmZJMFdNACvd1fWntDHmL4Ph
y3P08qQXzFgKs++G5n/F5sN6DO5BQuch/d+CDGmQdv473a2E1q1O+7/mPZSXAHA/
Z0RHAZYxnSmQRi4GFZJohIK3HR8yfFqOROM1uqs3KIsUG0l0WXtG/ZFSe+8HXUjB
YLGbt2fRCSBK3smZ5kw9aJc1m54dTWCciCqJhNpEtkuwcbJppxqMlaAB4REKVH9F
znmSzcZ64XYstfTfFOKh8D165TNDaa9WjQgKU28QaQoIItzEFfY5cFpYI9WGpdjE
B0GWlIgisdTvHFRCXNif1D0g3aslLRS9ntQ/Mm6WWbap8wYhL7Ywgo9ArPMGnETF
b1gesV+6wJnEGC+Wg2EmDQIjb3nPpd8XIDK8owTZyP7yhmNz8AG9OGJEeU0jemWf
epnu7lWUwkt5WvZsJflPwf0gntUnyEBsQRqSoDGy26JeOqHzPCk5TasbUY11/GUO
fUq+/qyHC5thGBbA/ghbEIx34/1Zw27w9xqdaygH6TS+DSzOwL3Fq3efqDiiEEtL
dmkaghSKlWe30m74rNC3wZXEszqFtbOq9fbpI3P2YnOPrQIgML5IA78kdXed+GGf
Ao2nQg3bUq1inR2TOO3WMtZg/8fhfcVWw/L+qK/ke4PLb2SzpAMMtz7s5km4eRMc
8y9Q/bw2SVGWr8phP+uXN7NL1pQLlHEjMC2saGh0ksML0OB2c/OOHlLCM+9Ejcjf
Z4j4XWkOrzUydS0Z77Cs0KAo31ZvKYN8Ii0kgbvAU6djd6ocg6DsB6nqVKVwUwQ6
K59aJyFJdkQxddpyc8aVUOW7OO264dskcPXcGFxstAm5C2kp6mWkmMO32dB/C2Qf
FblABeXeIYPaxX6RhaaBl5qB+7rZzidW1V3d7BGmxV1348MO9akxfJY6JsX2FOzP
Kap1aWSyXp4QYtGD8uZL9EnYdkNs5cDDeyaeobbdYzgHH+AL9PJ/7vkHUK7sk/h0
nlXA+H0nSSlYiqPbPZ5a8IdCVm707V7vIbA1Xm8yA1LsIbEVXr913WNlbiSkM2Gz
wLTvBRHrSSfMsNMIxIdjN56AMTbYqPof4TWdXH6KIZQxrtPDORA9KJzW/tvWF4oH
nGufTNwtchHcK/3X1jQnyUZVT+WCKZ4F62qHpcUeIkwKSCe+cC4vqhudcxQdPTOy
ZxiOXQ54WJB/Qn6Myt0RE5sm1yzQkKC3w8dz8Nx9cgtTKOu4xXwuuRkEEEuDZZsp
tJhRFN+LkFCuRGswbScy9pYObHuiywmdAlbfO3ut8Jc015EIYwHEyAsFrOnNTtT4
S8CIHQ5jstU11TQDpRIybvL7lgypJ55v/dXSGZhr6+G9hVTUWbX4mVc5nmEM4E3R
0Awq3yO0Zgfl/sq9ay8aw5OYGLTIHTA6+fLc7PHpMOELu2XApQX1mb9rkeHETI4w
cyAKzc4RezdCt7el2ct4KBSZ6IbldCH8KRFqMwJwRbMsKBzpm31c/US5Nmn/zIP0
m1bm1I1fx+j1Gwm7YAy4kaxaKnCjtb/QZS1IMP4HG2YkAKBuLRarWv2zTV+/2tWV
ww6TnX3jBjHa+e7BgEnWvRWvL9BM7s0LYcymToUCklr0h/oPwTqAc5SzekCGtyKr
lZv8gd3LCpNMEiD+9mEiS8+RSHKEZHHwn9UEyhB9Sws0LgPimLttCcarnszjQ71W
zxhl3qXI68LxYEnxtvBtBcgNoK/KsJoi2y6vNDQoKwJgxDWvsEpV7BidMe3riDTN
NdAXJmYWBJ5dU/lOta06TwThuBzwvkoMs1PGqFgrRZQWU5R4CElIlrP4qhtYCqee
HR1fxZVrQhN+RNmK2JB/smNHNltBCOZmONtZcWQpNpaD6dmnP6/GxzCLlOoXpgtX
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
V2L11Gp74syGwY4AHs8dGkRH+MDYmNtTlwBeg9NFZ3OP+OATGT7o6lH+lapyJQi6
reCbALqENdTxGmXNfmLvWXqyl2op0trP7Vs1xPHHckL+6B/WPc5/3Th7Rkj5vmLx
Ig5f1sZF6ByNe0ZCFsQV9iKnM4Y4s6A/OV035FD7c4/SwOPDhQjWYDEd5GgIYP7p
eZnscMexVwwOIlvjFMoh+Ogg7YnivnBv6x4OVZnNqdVGKvmMKBy+mfHKpeYIpbfy
KgBBMX7l1D4T+fuxPNrtd82nNidGBlKuAwCnfaQaa70YmcKWmDfK8iN3SpKJAw04
j/ZdagQqZjcPmhURxfKiRQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6496 )
`pragma protect data_block
gMSes1UscqRKbWlL8sSpL7Vtcr2eOBxTk4iBBEQhE2X5u2yozsNL5TUdbYTi3P/p
HrtfXoo5gKELj7JWC2UmQ/+zHUe+dZxNnF3L38hssoyuR36xfKS8N1228om2YPXM
A8QNVUnQRC3vl7uAdjgwgOgjDzihYfRRH6K3fVq80k1msSaRES3qBt+peBuPOoyJ
vjIcwxThBzALKs/uumKr8vA8JMxj5e7WBRLgOf6Plf8mSoSD8yw1VjPcwlBwNOGO
hpujaT+36JiXiMJbMc02InY0xvLD/E7vfxb0RXMgWesE26JmYpv12op/C++U9ndF
jrpK2RV9Ky+vy/LAnYFkZuxeIJOEmv7SzmV4pE5zUCw3NDaqiFAF9QHb9ZLbULq/
H1/RcdHwv6kccXH0UHxFCTP9UMVLOz6mpMwPPLHwNkzsWt5jwsY7v72v6NfhkEWj
hlSpIdHGN0y0x3z5pVf2ZBLUg5gwKstErFF1VJDNHySWCnhQakX1X5MaFfufhrdo
VGhiffH4d+DGzxlbUJvvqWiJgmmb0clXA8LAyeqgvalOzFYu+XHGYIypBYv6eM5F
cl5bjl+yybgbB/+5xLNfTTKfmAOXcOyg7A1MzOCOStZRzwDt0SDzM6kh0f8nJ8T6
L6wSCTn6qLoZCgHXHYdHZISBiQIqrKzhW7LsMwriWjaQjIKC0bg5OzOszlF7/nOj
PRQqH3ri5BjdWh0Ldm6XyVNCQmzhMDq7gUPtC3hInrRneVFejc5km7TPvQfppO7/
dP4BI5Frkqn2y+xDQ0CogYHX4w/CLyRxMc2Bvhwgayy95lJrJiS4KcqlvxcWzQIN
/NnHsrlNwZ/6JcEtsU/h7jghRDwfA5RVwVskfbhFGGPB0YEDbt77EM7UpSvWdBkV
VRfVRMeWkAAn7X7KfKg1NLHtv8/q2F9AAb7FmMOk0PmD2W9ZE7Ma+yfsDrQu6SED
SiI3GL/J62Hr19l5oSRpiZhSTm1OupraZ2O7ixnTdovcLtoRP+DFOOZggCBGFMZh
mvlWABvOKGyH7GQWpmnZfMzYwGKpv6N/Cv3p4QOA/eupekra8AYaUJN4t+vcirA4
6B0VgDdwPU6QpFNYdEpFN8b7b4OdzYN0BBPDqgqZ7ldE74qVoUTrmqQZaBLw7no+
wO1RogVNtfIQmv5tA2ytRgFhxKnpeizml1g9pwkMqR7jAZnznvSK1CdpGhODZhx4
rnqQ6iL3apq3lrBbnSPemHb/LEoo3IcBIAmsW4zxYVT63WrDJrCUOfyKiJHBauAv
DAMCEDncJFAgMcE7ahOkmTVc4pXjjB6+XzcrgWlDxWTkznZ9DhARHGT5+GliHvGg
VRUUuvy9gq2xOLBiLu/6vaoA7RqK4bscnPge13eok+ja2mIeExgDKEHUWITPf6Va
Vea5eP1lqZzTpoXQHrSyVI/JeW94xMxwqTGdirMt7yjpYnlAmKhigR8Nohc7n5C0
o+OUiN6Xv35BqFPynVs6uAKh7z0TB2IG1gtysUqDcV6K61J4PnAskWqP35RZLGw6
DjT0xAf67V+lg/YXf59JvtA5VhILguXSPxgiiEl1W73VzxPBorAwo1MxsM6P9Q5z
zXhB07TwJu2dO6FQKIgVA1ej5Ki3u0A3My9VDGWl3Fu5jeeN1jFxeWIDexluOk6n
eLNfu4IvlsQFhG6P4prL5AfwtaBWoJpV5NyxhH4vqwfHPAS5d91JBknZfKuD7pLb
y86Ku6Dxp6OsoAHWOC5qSk9a8zgavvhJ95J7bI7ItGhgq20bxS1nh18AT4i83g9Q
0++e7512isgMP8FKq2qoT3ULId/jz7Yi195brnOrDb53PO61nROJ6ve1ZKhQyv6P
JfklttdhKRDIbZ8bVd9dNBFX2KrRQxzpJgNUjYFOS5aYcEh+QEKp9nf03+ehRNEw
feRY4z8xm9SSOTgUVR1d6CwrkHpxz1toc0Erb1YVIO2KmfOiIYlT+lZkBhXmghl7
jPzxaci5z2+Nei+rkCi+ZEvWNDpWA2W0LqE6vcXV7XY3aCgL6oKnPga2pLHFF9Dy
K4LNEJ3ptklzXTsla5CrzyAAEPFX5SHs9/5BdQG3ts8EPJXwtHi/yVb5M5bzHaje
1Au4alTz+Ee6jt66q1WiXzk2hkixjYRagIFzAZVOOnWmOUJ9i3RpPxmZjzjFmbNZ
tB5d4jfU/L+6091biX1dYqb/qTEh7L0IhTPQZLLwoIX/X8k7X55bWP/J8kEeJMvi
5tbSDzLYPcTHg/okbQRm6hEJXtLy03dDh3P4b3zYJ6iBKJz2kqnV0I++8yXmFL7H
zQ/FRs6Yxgq3R51TqTtlfPuxe7Ej8POIAtXvbEiYrDpC48cCWhq2g8a5iqo/xPYf
ieHI3lS/hgnE+3wPiHtEEbUDNxU0sZDXp7t4td8Q0G4VxXNwePWX11TmxcW30StI
o3ZFHugQ84DBmO4c/CixfXeCQzbyz6v4MyELFZyVLDSxJvV5fW1pqlpEJfRyGzoG
MAXKji9I5Nesixffq8xYuTDRTkEAaU/HY5T9wSfHxZj6ixb49XgWCp0hUAKbTN7p
9UUKkFinPmOgS7fHgFmuEWK+2eJtS/xDJfHp4ui40f+sCOJRShvcmyHVoPPpwvQo
mlZQuhd7J5pjvE45JI+Tn1Vk/CyKAOCHJUnuwAGJhpShmTsZz9g5VwT+0+b9veJ3
5WVb7tGenC9gTQqfOkirVvshsBX4F0pAZbsJb83G6A4b3pfOXqDeZ00fmbKIJPea
E/jCDeAL8gjCWjumcH0pnQGlQXeGnz/IZejw6ebioqRLgQiCvoqzzkdip7YnihP3
fHRwDRiwiSCIoA9TWfJVyQOjJtypiNPlnJ3eMdmbdFqJlo7DVd8qi3XUkBvZx/Tj
tX0NLkBPGv2cYXvUTgQ0jGfQl4rg76WBSf4DrFPeJaqLU4+OeVtsJlFvQkJO55eV
Kq8S4iAGBTOtWMio6jskOjS43T172ZVJbXRW2oGtcl3zIqRd/3p0tT61un5FcDn5
AEstqgFMpsSVtN4dv62aA9NERL72mtDnscg/HrzLHCgSM+hRC2xynsX1k683toFZ
+Hgz+R+CeLIlIVpg/VmqXoGnBtHROCZnmNgWGzKbVSYxKGcLR9BFzH3w96w/+SHY
J8Dl0ndKYEelOoAo2loJi1hdlGDQmcazNOcc72cO3hUd6JTMHSLbP1L4kCrBFq+m
McKe7seSLasl6VZ6nvV7Z57NFEik/KQ2SwH4csLlKb/eq+Uq+tu+JfmU8soSCki4
gowyAsiHLc9Dp82UVINqFBjxJI0fEuD2gcQ8ZkDucmXM8/NZ99YLrqUpk9+9xrrB
DqDU5x4I+u7192ut3qUwN3rSajz/XrxWq2Orw5/t13Fi7vLQLfSKPqXCpv6Kpmfc
F/hDF0toG9lAZgImsBv2y8ZSaieO89Fquj7Z7yu8+nJIWWthDouNjMWqlVMAdjYx
wNPxQ40S7WX3CjI4oHEOGVjusqgoUO/kMvDAipJLoYZzuVdlwidUj2aPQSBNceQI
gPBykCZqswGcvHxbNHNIkHh54PtD0VUiGuHxzVraR8AcsddLJEkKOHlbSvupr8zs
6iPjff+WkQ4abUklUWQc3/iT2GLDFfB8OvHcYwV2EA/VyK4Duzx0pJsMXx4qX6Pf
jo/QbPQP3UZhDBmw847a59LDtugcPWgRIUc5E2vi6Bp2/ZBOytrFe91gIw4AeOip
cGtCKaoOtWmLvPXQJhcu3cXKUq2cG81jmGYF57fFevG5gwajD8mUojnp9mHagWR/
4tWjopdBA8dkV4PONq/F/xx4K5hnNwg2zFT6ngSJiZkbLlGtTQkYxJULk/UnjKFz
cJPDGBfaQmVxYLtX5OZvKEWC7ZAjxK4MvjHv6XPXuGW6/GYTRt3gONJEvS2vEOzP
I47trBTTbG2/yWA1foUn1lGpsSiF2uCweuqXaEJ/vowUirCq2IurqPRLYVbL16TN
XJbb2+6jwZdlrIBgey+WlDYi4cWMECfmXjWu/+jI0hR8QlLLvUqM2nAahEcFdjo/
yPcTqlGQo5OoKxiwdiEcNFPhJXQ0fd9ypNVk0Icj58WwDYnPTwEEhj3ouQwVO3XZ
HgnLAohAnKokprMZEZU6EMMBNTy6Omu+u9yFMmC579qNMxSYE+HNYRAXBHl6s/w9
xkH2MSfF4xcuvUiXkeZDOWlBWqLuy6FNbHHausp/BgdFWnot3+BAJLiJNXMlxlh7
jwAFZjbV1zGfczqzOorgvI8xcb3uSj9gug6RKDLFpEQjKEz+bl27MQigpXpvWBpO
T4eXREnHeOCJQ0fIlgv5nRbnvOORd3kzj/OGdOhCoiIgwMbZhcRv6UAxMBYwgFIm
IJoY5ALVJQ5Jrrk80mFSXsrGuVoYPR/Zg1m+vvLQ/TL11LwXgMIyD0JK9A1C8hke
2tniJzMuEBm0YJudV8gI4hOPUJPQolw7ck0m5n3pYtOdY4OPjP7loLg6puY9m4Og
gqie1vNKHovwg2BOzIcyPtZu+DM+sstiZkjeAEMIhJBtFraBAr+Ley7EFU497iaY
GZw8KP24iZP/d6enyNFdAb7u3jpX8bbb/dQIB9gIhXehVezfJW8oKTxhzAxrTao/
yseRFmM712TZNi4c/tNO+6CxgEd1atvwZ95OFYnryG2A8Ps/MNTzdxNI3WzHwaCg
Kg7dWXIelf0PZq/UL2SmTaLFylmwA+AQL9upgaI+Zl1fvElBzzINcGJp9ipFaMhO
/3Utwi1UrXx2rvi45vBdi3jllfAZC2vsmF1WWJR0FGIHKMBcyIsjsMG156p2mlsl
7F5oAi8FFfQN9LrTHP0UQCma/X0/e4Hy7zcpvSJjDle9xHfjrslvfd+OXIvEj8Xb
hxj4osgExbK/9Tf5DKzy6mC8roeVw2TAalr7HQXt1HhjQdZvPwqw6XkB5YqbbMnZ
i0u3XfsEFs4dWZ09l7htW/DD684++0spQwpz3dGbJK5nI1unVQXEBreqkcIu06VM
8ry2XdGVVO9iiclI6rR5i6G6+o97EolZkvCJWVWxOyiO5xlvWm4xBttqK/LDKe9L
iUKujCyG95d9s6rLyqkFfdZ93B/8F/aac6IpEqJV50U4qJk/kiqouhfNezVfUh6T
ICMwg/K0ycFtR9KrSvFD0xZtUdjDhamQOLWVUx4JytOiyCa9WnLkQR6bf/De05Oi
O2MLQb6HbGTvdxgMiIqJLWHoP7/UgRRMiU4QQqwOYkEg87KSjNBp9jMSMMAnHerI
EMnxdcE8qWC9R2B4XTaIb7WL4of//vVFgVqlO70ZXhYArjiiW9mVAVHOyMat7xqJ
BbL+NUYbkVRNp2oiGv4An+F9r+B3689x6KhnMF35bw9JQNJOfXpFYjAzjMRZ2drm
Uv2E++n0CRGpktrJX9GkP2hesM6gPKfsabJcxmz2J2kaJvQ8GtHV+o3Ew6fwpRJR
t7s5t+w8LH2FXlKQVuGHn3skVfNAgpteeqxyl7BlmYK9xd9rJYHnho8nJ0glfLtO
mHk7M/sM8JeU2AifbnXIAddOx9apgminoFr+M8KQTz1kU/X23DA2IyNtQLpPt/Nq
nb4Hp/i9iB6cvzR5wMqHjEG8GFRIx6O1H5kZt56G5jNFbkHDBvZBnJQEK+XFyfTy
6YbvFYM78w9PSZF2KtGI5M5UgElWU2mLGsyoWeXZFxNgndSR3KNSLVtZS94Aedkv
646l8Ndkqt30Hb8j9Fa1ZUIknQQbhDHzX2I8K9/2ud1GLbNW1yraR8BUkzeNOl5n
7o6Xp+cAt9yhGbyTRhRohyNffq86CNByQ0yv3/enrf4x2pU+Xg+nAFozUaeVsONi
jKo+mHhXvz//cdCY9Q1+g9AYC+ZMfDtUxHhW4zD+beRVtpYQ/qJhFXuMYkEnU9LD
M220W16fNZJWVtYsL1fYfUR//hGZ1Glnsj+cQwH5fABiCjOrJR6pgj4dnSntRRT3
jMEbY2e+TwUAGo0kYKqyPHIDMdpH3W6avTq79VoZHinYkcDmgNqbgvfn5gFmK1TC
sS2uRlkRGcFaa5uBRuHopXd7wD3+9GhOQD3Q72kujZQT/kJFuN7ZUs+7yWDzeCJx
Hj4OHSUqwUGrxobOc2pT2FPlcb8DuF1gNubQOaQJiciehwzsm5mnsMdj2ldtyUBw
5LH06GZ3u70ySQtWFA1kZHDfy5fiNV7wo95EmICp2w4TQ2dLfXW5ZkbVVNTTPZod
tRTuLK712rYMSUjObSg+0TCeJh+qCp1zsABxL2rQV9zXPFuporDV4zn83M4R/NqL
8HJ2mWTelfLgBsp/Sqsc5BnOIO8rZ3vPrCmOiezKhTPaF1ejUZnhix0tiSH9DR8j
C8YYeuEhs0LiZb1N6DeMO/6cGnmtLwChhrGILA6P6AOzT6hr0eRsu5j8pTzMcELq
e6rhcYZlfsrQwb5lEpzTsBLDeyZATVxVxCCtJPxddpa3eVh/0w3s5HwmRhzqbO+r
dgrdyqnMMNlWy3e1WQxkO3bYIwLnCNJrkjAPREQMNt4Aokgcbf7jm7xxjICUorCV
SrVumQXQW8fRoquz6hjybKumzlQTRLCs+HUbDEkeUdVl1rWF+mI8LlnSklTnO8RA
F/PU6ZOcRg47xiYFwRPzyq2fHA0oeyaMIdQsER3Az04pCNV7Q8CbWRtBGA/Ym26c
Tupq/l5zPlmRbRqVpT3bZydD0wh1zmF8BWud5j3FpUfoUEBUcR0IjljpGBGxyeeZ
EnRH7YdqVOC0lCz8JfFLJ1O6rY3E7r/waWXuZsijVQinFzpVipdOSx+/XTqoqwfI
ltYA0zDJjFKXScyFi27dlKB5e1Ym6wII/mHIdCz7RoXPUePiBR4uJ/UzAXC1b/Wb
tVBfx6NxfMS5iD8lQQAnVgIf18G7KN4r3OkGnF71mtM4yottGY7dSjxYZge3ExDd
0NRQR6toe+69SKou3ju+1hYrkEsKxGVLjlCakaF50ze/p+stPf3It6+6eMEu5rMv
pz2tGuj/R51eg4hD72KRlBhoqT+MPxZCImNudDNRXxvjZ01EsW1vHoOZeRdcqOf0
hmkEk/uS5XmS30Jht5pxIbgePuL6eUSAavbgcZLWgRG6q25S8XjdfH2NT/neMNtw
kGmZHfmLeYHAdFvEB0LOnWffqjjXbgvpVHslRaiSYiTbNusQYD2uajGx3iIOFudF
eCjPddNSie17wMbDqXNvBI+0ZNvMZBamFnRMQ8I6mgnZchuf7E6x17FlFU74Mtph
3dz4Ix6rt1WQIE7IhdE1CaIypxi7lY1dmYPKD95buKpIjuvUhNXzAWUKiZhIDp1I
Z5NIewWGbmww0mv6dFjf+kogAK1PO2UePEg5vVhMM1nwHpeh+48JIWCIlptMeBJ7
t0+Cq7sSK4iKxi3hxOwQvU9TC1DamMoI8DrvZvMP7N4Fl/yQsWLlPTzu4bvC5EK6
8XgkCmyEpGAFLHyXXjyrZb9u3rKLbWn28Fc0q6nMhySA9t5Z7h9DevU8215Hegch
4MjlNFznRqE2M6//tDFD/Esy6iirtzPjyyEHOauZzrcGgvYLasJ3Mf6SSPpdoNkE
FKbDJEB3m7FY1Lip3+UIoiwLrllpeCRnAUIM7V1QDJWuQ0Wet3hFppUY5/OiwICu
4hzycSwjWUbFOWLi10g9pva56QiipITY4t2vUc/Btd23tyLnJv4i8bSiQK8lm8l7
MMYvJKIk0HXL6FgtpYXDplbegxWxJl5DmtJR4zJK3dMIIhjD327fbdZCNw76s0sT
xrEWYNTpBqxlrwPE7wEOEwTehLhyCtjx1myaW2giWBTEvfEiNJXgDDLDLFLqck2i
t6spMM+O8E9U/YTXZmsZ9eHBy5v94O5h5bg/eZRlx0PYclh6YzT7zCxsvSVKPNF3
D+EF+o8K6wR1CnqjIzcMjHeAXctJerlpI9U34j1VgPuaCZLhVSAwwzSPJQzOHcHX
ef899Vh3glOfO7I6qyWif7bQcxyQJ18tOsAk5tSGiHZv64z2ciEU2o9fADHgD59I
o+5ZABiJU+pbVFbS2v3zzM1JPveNfz4tAR1Z01ojgXl6wExVIAXFdgrhgOJe1lmX
puea1yHK1F1y1oc4STjRhPL1MH/rcbe5wJVgvwpYjJ/b1bv1eax74x1lobbojWJ1
e6BPVHguviuPuRBsNimIkxYiGFE2UIThVpkdY4lS/DFRohU2mm++9IKEinAzfOsS
8JkN6/Y4M64AJMRBHM0zbFW5DXJH+uFNtZ9lcTYjOSFreYgnJ36LhhHc2LWDBYMD
UQhTJToob/RHnmbbzy2MWM9faxCAd8Q7EV9Tz5iCKNZA+Ynhg7hUZPM/Z0evY7Q/
GKCdxMOrw4t1va57SZED0bB/Lxchzj0K8i9IsiiDBg6YjOnY8Nk3wW0IQimKtzGm
m7LaJ/yXiaj2/sc8MY3XCzpHcjhIx02JFUtalpYQ3csL3XAkylLye0YvgXhcG4Oi
PzvC48IdkODFXsAu45B1iTLKVekHQQ5jX/9ZSfRduxYkDVf6dDxClgP9vyZn+so4
FUVis8kZE4tg8I+G1mDoNimF5SRmMfiLhUIaYg/RYbi7I2S1aGPBb/S2T0eS4XPG
IIHuFpbQ84fa5h2Avfb26Rxx4u+sPxgKD1uz8g0W5FZ6cpY0oeex2xZbpadI/vYY
Sxm3hu15zDgpGC9D4Ki+dQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
QnhyBKJoe889wqM3BVC0sQfoyc7BjDCeu6/2GsuExLxBL1b3r4ovHxXgB+Tr3xTa
D8oKO2Stz+lWkv5PGkHXDMM3BDXggqd1eydG9+VXndFVHdB5SI8KABw+sqT0mJ5E
x0yA7qnHOPqFyfsnaE9RfzPdEnhPalfX4Q6E2vwai9BoDsQO/A2X4tuCV69vUwBr
v8jjjCKb6BuT74PzOUUT0gl9z1yc+RSacOoazD6RhDohGyPlKeIqjjujHvlinXHZ
0g2p44MOt/fy8LD+7kTvfcTZIdzvWZw2FzzHopOGi2DY1FDAzC5EjqvTjijkEvM9
1gedgGW0T3uUX1DSMeoR2A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 23840 )
`pragma protect data_block
TCUacorlLKhcRyJ/Nd+EC6DJFuBta8AZ9mRFoXSmwSO4BF/J7k2vZcfuYqgMrKah
iJHnDXXIrniI45azEkgaXZZr4O6g1PE+WuYmeKnWfDJBIF8zOsOYr5YoQ061EQo7
/kFvUc/pTA2U4oBOJkb/8SplbxFwaSd+rrT0mudzuMwqegT1DVUtvtMLHopWzRnJ
4Zgu5cHKKDn3rY1MnXb3Ea8fqIt/nnLUHem4dn94Q9fDWEEvwwaI9aJZlWgeWNYn
qsopfmwkQxu3kCn9tKJEK7Sy8I2HL0/njBwyt5cGA2WZOLa2d6TSGMV+Vr6IglMW
wWjygfCwOEvC4znxI26DBfh9M0i7Z7bn/mEKsN/4Cep79SvcSLDeD1vWVMYWx84t
zFG1hs8ZypfM43IrVPWmVGWQ20aIOyMB1pW9PFOyHVaM8EFFf0YQ7bPTMHNic2U6
XpQqig2uTZpDtZhem4XGPS9IWyJhSzigvSLPPGtxcJ3N0N9LfK56tH1g6a9oS5aq
ntT0McM3tVY40XkXKZgKs1WZnA28zJwejYAVES0Im/7uIjLtVqtbREq2UUrb21a7
QIjyKBlvQzu7if9btdSvG/BZjoqJwNCY/hrolTPBIeZO/9GexmHRm5rq+/SAtA8m
KxP5Rsxj7p4iWr3VeJdu0fwOfb5Vk7tzwYvomkdxYeHMA0882PkXj4FnjHzb++m+
DX47xb+9/b05tvVgejCs19sziX7xGN6Ekm/D8BUHM0o8QMBUIgUwHeAhYQ1LfQ1Y
uLUdBH4bbEwaptq2kP+oC7azK31aImWYLLcwxXuiB+QwCuZhp9hMYCgpGyIJoXA3
f22rpJtjRz3zQ84YC72FupZOEb9OYGqy9BxHSVkV9J40wHONKri7SZ4JI9T+uLd/
e9jTox23PgoEHHtPphGXakW9/wjxP2yE2F3QI4m+Tufc4Y5MAu76D0FtdeH8LAv6
uuNGioPLfBS5ViLGTMEfl6ULPg0QQvYO34PMfTwi0pG/dha0ui44y9S3hzW139Nv
tG+fvhM1e1iI1E+oYKbtqZTSOOQqb1L2paaDZZfWOoMBqdYcrvK3vRwcyvWc3nI4
Xibg1ojTfRtPcHhDyQLvRbNS4AQOAQrBFuXbyCvqh023dEsKMFRvLcGvEnpDuhoy
is/kzOoiaztBfkZDtlf2Ykrbo0I2I2zLIHzPdQEtwc6vrticymDMaiUeFS+MtExR
kAI0Zea0C3aHcynvX47SFV+IxW8EzIJ7WSLIdUN4W4Uzt5mHBh+nrmV7coGASGzX
uyqHmHWoZkU99XYY6hTQEQEBqXHu9a7OvHFJepZLB2yp/DTZY/iN79ZVSvy3Ak2P
kAZrl4sNfHyQIaZ7sjsZYu+3m3M4V9KHp+Ya2VzgYb4bnftXP3yuK85nLL+5nPuK
ee88Jrt/H2X+zP5ZlYHSZiV/MTborkOJ44aIxEfnFKYOb5FOc4ojVkN0oyyeF6Mr
dkyyv0c112htk6ODGBdBCmrU+zMFb5jhYTHXUhu5O+/zvgxjR8NJqx5dIUmQAF/V
ImOxLWBApmlbwza+QSbtQqvCuQgyZkB8Uvrxg9IKWAoY2Dpf6W5hseY5KUZV3Urg
Lr5Zc1Krm4SXoGQ0mqkj1tUED8N6lSGGAKKXYdujEQyKffwNp6UxabciX8hCXFQg
TL3QxLIGgR5Jsxy1YeeGhvXLh+jXf4BqQn3LvDjm7GrJgM2mKJmfrU3re0QcP5GS
clZ005g4mXWx9mQLfhgh3uGZmPUz6EgrcENV/HHrvXokRH8FQkT0vg4FQQ0tKyhu
BaTK36FJnDBRsilwDF1wfgnW4S6VMzZszFHX83+9sa1c7tnwWo/AO+WDReYXLpYd
sPxe1ghAydnOTEAfrQWaF11x3yZXYxPxd3USuPCtrdOZYj7o3Q6Xsx1G4hdAg/Be
Yh+RSTnfVT4eq8pA9dXVqhyCRvDeV0Cj4osY2U5QWAHqUqs/KjW+ZWLdtwJ6+2eT
fLi5whsDnbAC6+5H2KwiHvEnCjUfbxNHlRQ8QQIOeOnQU9S1nDJS8mJe24brEdAJ
pnQhvaU6esQV1lsqcQjRXLcR8b3gzzYBndBzXCVnE/OlziV8EB02y6MVs45nBrTM
yJqCqBAQ2BdTgp9BETtmye6dMWu1mxhYKqAf1pE0xiFT9saRufQrXthrUa44RMUM
lOYFWpMAY2eoCkH+i/oFmwSoyGlx25gWgdkXNu69RSW9D+TrLE0Ya9iPOehCZVlw
2wvSLtay+ZUHlWXGLYd7RNeacbRoTwPo3091S94G8HMph42g3Wedkd8Ijrmy7+1e
yYBG8T7ciwmwz0sKJKJ7hztaFMZrFi2TMBCuMr6R8GyfhSEB2a51VjxrdHcenZWA
cCZvWNvcAe+YBarowN+SFWpjIkxrl2DfgI/AddAKuy7Ctg5dwDoT9fvU3GquMh5M
iL/hRZCO/2OTrHP+eVX6nJ1RyJP117Zcwvtrf+BWuyjqYTMwZ0Gpsg5dUqYJZWPQ
SajpoZ5WoGaUeL1w6dUGhf8Z0zTsozM4L38wQo5j+8etefHK9sLFi5WR+dLZG7DW
o+4tF+Wkb6nH7dPPO/8ZnyH0o8M3WHi4WLFuha9T4cbUAWP/xxJEciSaMxDIeO8O
1lB4ZalIh7DMABCpnvmtTDtSlBF/5B7FSTuDdRY4rVx8ZTohOdrP4iSKMHMqXoia
HSH/bVgLf5p5zQlctYF6UlsCW/LDSMkn1esBNlKceaU9XlsK01YxaPyWGqnALEcS
B22yK5piQhhoSUW4cA5FjnYN93MA8+BUS+K1YiYHEs1mK60Y0euWd9vCPmsITkT1
2aRW2Qtn+JOfIIURvuAYoy7AzhxbuV8vUy9r3QXyuc5RHTuR9FUhZVrRdlxWZ2z7
tNGNv13/5LpZ2ckkM6d2/x9bcLE7SfUk+EvIEgvHKTb9wQ6YVUPFp7JYWxpkreid
u8R5pRmp/FfFXqZo2oLj39Dl5JEfE01u3WySAAlnF/mb5L/FnMxEzlb17ChgrKjv
SSm6+idO6gdnryd/ji5Tinlfp6ZHu0wd5Oq6JbVKuKYLFcQucZdtAt2Pdglrdmur
4DTwfQB92YKAIT8BYb3rOx555wriJTqDIu3ic1fFZkdwpjVWDa8clZ/YfQ86rzUV
EoTVCaS4fuNu6DeVUqFf+pzwYzuhSac/8p78YMIE40c+fQEu8rpRDeinWx8F41Od
XwobFmYvnsPnF2Kl4xbZjr5LCuJcgWLQtqytKyr6x4bvizrXyTI9AJ/0+zgIXFLh
vAgJL/4qoJRzqmYJWXwqMFccfNV0KKx9cmy7yP9Cwa7GMVP9dnJIJglMolpp9CDE
5Lp6wKwPcOOjVBu+wBoxq+VNzi/8gDuVHPXeIkLPZxdBregvukDbNzRM9a0AdEeY
cTgRE4G8D6HhFumxI/67CBHI+0awOUfjFi4CrXCQ+5QKl7YtAYoTC73sR0/IonXS
oZ9Lph8vC2FDQOqXdMYmu2WSepCTavkVhfICJxe39GjkVePJMciUibcY7dVno4A1
NRDsMnfAnY2hvATaOhYnO8g+iq+Cy0ocQ6pifX9YsZguSpORI0wJGVBztl9u+Ro4
vEotgAo58gOof5YEIY96DlFWItBaOFkMwEJNQAuZ4D62JKlIiLdgmlK19JltGVvI
RDP9eBjKCjSQ+Qe+82VTYbKCBIp/TJWt2Q67INZeFdYV2J8sxiPFQKaDsLF6kEgi
u1mT9e/E+YYyxmoDGrBSOwK+y19EkwlHqUvvtHPMahuu0wk8oLHPf7r7SdHmLJEq
FXd6jV0ROgrKFYAZa0WKtnwOZHYaHnGV+EP1acfAzUpTA6wCBkZvMybCPSgKX6Mr
zi2QeIHjXTDolkPf/FyzonO9Ls6DCNEhQRaCb/LkDjFqij3TqA+DJszMIwk20ZLV
Wsq3F8APISbzq7Qjb9DKTHslugtoKgBGFHpbfWK0d2m8bI+F/NxdZ9HhdSH13PWn
T+c9HsF1/nxtl0TX6Uvis+golL1dUBGACsXwINFfHzsCWbYB0QfB4SobXYsz5BTC
a4yJVjGSyxsJxUo9tHm/9oeNKwDdXHJixxWN3zZKDZ4un7a6SDpz9ZnYGj4++0fe
1j9m8VHcl5camOFdukshKoZhkEiUGeMIqBxL71zh0Bi27HDzsv5SJWEzpqLq85mM
3p677gbSkj+xRDnM5TV6u9GqH0G41rc1DQoKgfeG2r8K4TMkLFl6r9ZT2snlv2xm
6YvdxiqR/Ae2FpbkxEVgFTSNBSclDSr3Qw4mRtCCSsuMcuYPnVTX+iTb8DUiCyAv
PEvtPZLml4hSL4vz2cTwndspwTimnCgaDd0CaCSHmQP9atIqsueUITkRw13nHsJl
4sEzGqBmy5kMBqwEh2w9mG9SOl8cOikV3wsCY6ToElKK0ju/IMOYi8bhUb3P8+h0
n/3HLTOZsdLTSAu4PMg/VeCbygQUZBPZ5i7CfbwjppubUwnDDuwvrWSD+teR2lur
o2/4OQQ1bNf1jSVfSIObfEHCJsHTF3InvHsxK6FGQ2XHnkGLVtd7rIxXTPBCPxwf
Vy8dLoEIq/ay7UUr8GRywE0sWurpZ7k4wAe7Y35b1uXVzWkjSLegV5YPglO7CxWG
1MEVW9B0YLdUMzMRCvC2Za/m8aiUR/Zs0hG6XWw3jbpL3WcYbJuEzqurURbNJxFY
1OoPw/bziHYj8CKZZBaTeRCA8OvTazh4ZjVoQ59ANuQdulX6qqNO3FT+RRM8rCmF
aoHaZMgRq5o8MmuuYoE0djt2oFwuxqgiCvDbTt9DuUX1AW7f2NrEITB6QUNRygEB
lX3Rp7qAsWKiLXOMq/Je4ABK13uEcFPvBcrGQURCUwD8kA7vf4jsv2GzTdGrysYM
hNnRXsg3UZGQuRyk71qurgJ4nGZEL3rc6VTfKiSz4Lo19mVMRX//cZQAcBykITVX
+y/MfnOPMST4gqu6i56077ZWfga1VAyoQfYU7nxlzOr1I+eUJs8GCn8qRNJlz4di
3VYrv8bsYmggl+MNdDkrfPxAdez9sZUCYfRINmj4krETW6W0A7O1gBkMwBBRjyik
ynnSjKTGeBrKvfknJIVeYnM7IhQWAzIbD3UszZAw6ahBw3WmZVlQS8+LIPfXi+gq
yy/maKM7riZcRCFehzppxBPGaSMZKIO/Tw0Gv/3HQe1fhHWbVnXM6Pdl2VQaVl5o
/os9E0LaTcs4f4549We6e3PXOncYVn6fuxo+GUR6orkqb1Parl0E8OtXoxd7xXNz
99sVecmi4gwqVdVjm/+p6owxED29uNToyzSJh6Oq/02TLUPqJTm8zInqF3hrbOEN
mT6889QdnbWX/v0aDCMqKAHeCFDMPXSJX5B+rhNQF1WUcLDBH4LmAdB87FeBGiVW
e4l4JBHeySnd5qOQUMQl6+4YsA+aNqMA5SOpAh3ca126imwwamgmuDfoyqSX+Xi6
aGlA3EA9t/tEsT+ArNvRfrMgmz3HZul92ClBRowpwT+8C2xSicOJqXLiRmQ6VA1Z
0hTEWdrKwc9CI7iSx5kETDcnpcaWRfGEO7hxnHEevHvltz9FsnZghj+9nO30utA6
sunjW41uul8abH4O5An6Wq+xjXgL5BVEtyOXxC2womjcILASVasTudpWw6nxSvul
OQD6UtwYmgbNlt7SJzwzih8a3uzaipfUUdpnKI/b7QOTwLuJwgH/RsjDmo/CAHay
cuDqjkHJ6lYoFG+AMCIVqRgQWsoccS8GMGGmjgICmPUR7V7CZJLnwU5pTIZmJGkt
wgsl3QYnNZNrMC0MrFXkAlKeMFfHoRm8MiD8ckBbMbwiB8JT0fJqytpbbRPJt8Fx
OUg5awu3suqhGGmQYMbxYUBJXmLl+grRxH0lmjUmqelfBf0Sap4NerEKBHmLwYuX
/XUfCNrNtlykKRtfRpCZ2xT/FI7sYY2g+P+3voC6FPytwmf6Z4WJszlClIX48Qdb
VXd5MfXEOj+kEnuj8GZZPqyIVX0NIdoUc379JECdgVaMOHjiO6nca8a/qqrSJ/RF
pMQqjd3JLqDynKHbTVnS3iiZsXrBUPmotM7PabMCBv6yK4wlg34StwFS6dQFpLBQ
+CVM7MUZ3DPq2wNNUuQ8GEGN+b+SnS1TbF20s1X9p3uix/fKHwL2EJC5keCkKaFS
M6G0wbrpT6ARaanEIVkMewZVPRTELb98ivQ8KZ5pKKkWRMmQ0/LCmfCvLFD3jEUS
NqX+y+ZmOLBpZSWTo4ik9zJaWCFzwUP0Y92xLEqwiIyX6LmT4/nu8eQ34zghOvC8
/dBATUheHEUY/ePdU6QG1YggoVEl+cMH3EC96VE/G3jczjAdcX+iOPE1o5ovlpLl
mGlxXB4qtDJqza/2IcNGxZ9O5MJMhl+CrCXBtZK1y0zwe696z4KRA6GfTyV7XMXi
HZ5LLA1u69tdEH1U0HIDQKAVcnDo/uqQ2Zw2eH7iAqtv+CR1qncykoJorn9CFzHC
g49uwlNUFn/rZLZsdaOBBSJyyNQVrjghelvLUAbfN7X9VCpaEia3wzt64L6u2+rl
8wYa05FKT3C0CGHSY4G1qndKIF20qysbqaV9eDuWZAdvggOZYCvzgMADQYUpfagY
damXNzdLcSqe4uVGtth3aqiL1u4b/RkiFEinFdu/XS8vkIcOBgGoAYfBTYqi4IkI
qmtsPreVcbEmoCznrrFFHa6RMolBVo7DsZ9wog8vPOzJ/r4C6E8j/Si3K5RIiTW/
YHiW3w9jw44FgwHuDMi8Lok/950j05+pTeALjy7baOOtfRyjW5dHUo+AzUtEG7Vo
m+GiXRQ9fZRYrgY7O8bnGlo8S+l0tCEKQpXCgJVWj4EncTMu4ed3oT3vBbQyghb9
x9ErmuW/MU1gktHq54jqAoliNzCHTTnBcsIKBBVbKOGoi4RdDOWTtmPVYlZjs75z
Ki+uLuyzi57emMFyvTKafh5myyain+uiPq9CKBOiZgl+SAv/P1G0crJsdakphENJ
JXHTKP6j41DNIBwTcaP7gDalTsBh8Jlgw5TFvV532xea5wckAWZHiL4smjrJqMsc
kfMf/TCJoVPb4iRJ0annvaT6PLdQbhSo3xmFFWu9XmPhGV5qZbCXGhzu3h+OD4ug
sbAZPjfQyCX2eBL2CVoAJAI3YFq4uyNYrQIpL26FBD1w7F5UADDmotuIGU/7K1fD
5GZTLc9lro/aB08I4PRYZQzYdvepmMwsvEYAxVn1xMhVWyDcO7OMmDtLmN4cprHM
DjE3kaFCou5VMW+slADn6J+Ki7n3IRx2E+FtLMg8aWW1Xjf4j5lJJ+M5CkUquWdt
RG1B0W2setGposESo6cnWuglD99eFcc7Ar3hzWUB/zNXzg/WP68/fY5yOlVjAt1o
gCm5Kl3p/xgMvlOP0mSoMlhJOsEwFJh29JVPLWnacd/iMGvoUwvENEhUs+oUSq78
6XS2rnTjUDmCWrkIOm6/FePQttkQUEEBYcZYRX4aMwxYnxKWGmGELgNCFpfYBnI9
oEC6ZfLWRklFOBl39Y90Pu9slKo5e3jhvcsb5NAFYH4p5xzF2IIU4JIiJo1ewWw7
C/gy+FVWNdK8A5RrQ7TlIXvp9ahtqgcvxUJ5gUSx0+CYNTsZY8GRl+OwXXC8wHVu
1cp5A9a7ZXwVObI67VQ6xWuqVIwJU/ouOiwNvTvD9Gs7qim8HJaUJgM2H6JRTDD2
vPgyr9q6ZJcIlAX3SjN3dX2gd5LsQ5YA18gRd6ICz+TeE8YdPQSzXDEnTddV0Lyk
f9/9mfbw4pjaYSu4ij6bRzy36mBTFYurR9D0fYFNVjl7J24HFvas6LAmHGd1YuH1
dW9OLbluP1VbAMHdNQasMh1rFpgW4zEODPPnwxb0N7Ra7D9bTtH90U+D9NO8gYZ5
B57WOWyCAnY1irUGlYK6RVZFqyftkkSehxIIiBBeJZbiNytTIvd97KeDi37D9HPY
r/0xAlrszwSo65/DVc6bG2CLek2x5fqM+mClNliw8FyxgvFH+Zn5GEcZ5HHeMm/N
6rLevtqb09xZkbW8F1R2wGWy0hLC/2nl1utuODaT3Drfp7RJSmi3kvWZofG8WVeE
s7S8sxfch6j+jJ1Shw/HBlAZBQbXDgmbhSjChkAkrPd/aL0/WbchHymN2JAoHo07
fJ4TfdxWqIv9C8WlJTfy84DApgnLmgFbMOhgotHCBAFuhn4SQN6cgdFcBYCtaHGD
VVlX9lDx+gm46zypo8onEwDxhBfAKfm6dNRnCeAfbQQhg42vIyV++O5k6MHa3zd1
KY7T/dOnN61RViudy6xHML1KRMC4if20USwQFtN3huVMkyjaktRGP7wlxGhOmBoK
a3XNlQqHambhrnT49aS4+N1iC3FQxfgeOIoa9qx8IjwtRDCsAvAO8BKA88x5SG/j
Y2ldxGY4Txpa6hkMCERJw+1+FQjGCETBtEpNU4R+jT4X8w7X/SYIBWqYpdAQylzh
925yuo+G2yD8I3p7vhRpigKv8SCBp+tKB1L8QSs8ExtblIP2WlCwprkzekhVKycR
OuzmagPFZnGt9OxnSDHPn6Gy6YfF2TB0pW1Kn5+LLBxHAc26B6jQDLeR/edgDiXk
Yyqh2Y8m75hTJucxVj4orz0PMd7r2stZP/DPp7ksjYeryK2i89WyK4WxHqPHnOiP
tN8yOXZo+3XDVIrC0zHDRRskiC9t6Hr26nifB91AaqwGg+XoyX+mOIh9HPPMUHch
TibjbjIOUwV6bk+R6A7Pk6OVcUotHEoa1Nq6Zq1curjYVivJWQYXS9FhgKBUS3Cv
h2a/GUO3rDDQajWuNLb0f7LPAmrY/NclF/r1/woEkfmvuOTOk++fH+3K6iyG9HPm
RC9pq83Fccy5O33wcn5/1vHND0oUvCTGbZ1Q4rjDbPEGolqBoVjfcHH5dwCti8Ds
8wTgU3nUkw0jYAIJCQLydUaTMKMVmRl0mnTnyvdOIwD3kL6RnYfXTiBMQlcXNlVJ
GAfiiJQOMXF8kNpR6BMFIWL+Vr08ZhRIFlJyDUESC7z6+82TQXdaq+UI2c8e/zOu
jlN7dgjLgLoX6lGf8T8ID9p6F+nZB4g/CaDuTnvTVI7heMsuB9mXCpQjmlWx5/NR
ZClkT7tgbbPHlLriTF6suDDy4GDoDUqc7LX+GMePWNJXIZlT+2SKGF6PN3toqlIs
3Hd2JZoi29SfZ9EmCupGbI89GcnyGuWTHEMpU5QijaGv79gL8KkIZS9PvLKh2SMy
nlF+wL+kbD8hS+bH+YLTu0rIzh74ckhriw1QK/zI0YklpaS/b7lOSmLaHrIQoXlS
0QkBk0w4zuRJDUhvBUNBLLHnGcu2dSlJra3p77u4cuR/rsizX5auvpW5yZ3AKqA0
cwKw0rdt9ldcxcfD1uA/1zOr2FHdQkypqELsSDEcl19zmgvm8UlfQGr77B7308WT
PmqDYU3uqVRdy621PKUXsDxSB+gRy1w4tvSgfXHra0ejkN8OYOKFwR4XzIqYaSO1
x52mG13Jx80q0wQdcjWq9FCH51shQhcdEArvGZjv39SejUydVLUxZkAoU7v5QXih
cMVjAOKHCSJYFfCQmkurpuEH4Ta/rQcxL8UA6YQztc9+/KbDRVTzgYSnjNWijvUj
c4KRbAUm6zsWbw1QtonxOfGOy20ANZer4oQCTmaApZBuEYxt/GeY1tNLwwuoQqhR
bpggBlZ/tn53rLKH6TCqsoJxzd+Q8kUeWOYkPPtYTE38GLo0ciRMeZrATarXHXIZ
MaJfCM6uo4rX4P9p0LDIViTLqRtCzR89uLOY2+KfhgufXzOsIJFl1Oja4r06qS2g
INbA7j8GVyOlyeSmpY2ix49+DPg/Wp7Kome8eEstrGvJsabOmq5d6HE1KkfcfRhH
5xCrFc+CQYZssgdrMOFRJ3RYhGiZLuRmoQCbHEsXHjEToWBhV5MPKMDiDr7QnZAI
mJyfp8gPeGi9KOob8YE2rOtFQmMSRWqSi3r00pTkvcMw7nTY6b8/nn89e6ZRZkqL
PhVEtlQLM3v+Wa3fEt1WM7VYX0IzXinPA/S/UOp1ZIR3W9oGmvcArhm62SdSYCSk
XW9AAzqIMuYoj4MOp7d5LN37ASJ9Opc8B6HlWa7ofikhi12xE0RNyEUUxcViWYeg
Obie45GLP9bv3lUBHuAadmH9XEK3sdLD4LNqMf2quI5S/sv83AzXk9Iy6CV6z1ca
sGyy6c4d6NpLgxv2i0w4PVH2J8GRiEQQjozGOEVtZxYtNeHJdEldYycCy8nPucZq
GmrdQA2TiOMuStfdDsi195t/uJzTiNrE2H/+5m1XDVE7FtwIy19SYwMJLHCmy52R
SkVoAntfGk8jqM8MFSC3vm7hNS9xnUr6MuxHSIR9JgZgHCbqcArhNFNzxlb609mq
nNtDa19V1/nJJlBpeO2e6UuMTjSrvh4eXxYALadOX9WoeOkLkyw43p5iMQdb0aZ+
o2Vsc8+l9OQt68CQNFtQNHD7sq6aD7rJ8HcEVPBPa83b8BxW7TVk8I1CmxmDH3Hd
QY72x7bC1dGIb61EDrazuhL5NkGqX9rMu8MFi0fmq4tYWmPzGmE0Q2efOlaMLXy1
LzYd3v21vcYxqlsc/8dFTbgYQW5ljggQdIFo43zW89xxpB4whnLyFsb0cvB4+gHw
X4isOX98kHaqHCuvm4Gx0omA6quE4gMA5jRqQXgr4HLsApUjdTW4Y1wEDRCNzfDM
2LEzMBUvvKEKI7fgXX8oI5FQyrvabcbwxw+TTh/JZeEGQ20mu+C/GlUEUQ5qVbwc
8/fqSotiZZj7rMXY5vCIav/HSqXdVzrMtrp7fVjGVQGb/9burxpkiguto6dUSsUN
CC+TBJxfSm5HuaWD2Hf9/pHZYogGemhGz84wnZl3s9bEeS4d7ftJZY4BNrViVxJc
I/+uXiH1G6lqThNCW3+V5e72x7K1ww5oRhRIW+C+LS3pskAmt1zMRDq5FTSGC3bU
fJn/ZictB+4s6fkp+mdOsVzEwhSfYaUoD+ELyW7oB6OpXcMN98n55Tikvag6/vnm
S9qpDhTsh8y2zFGa/dZ7FI76PLdE3JckXlDRb/VWlQHT6worJ2xbnJjMnNzGItCl
yB4AAnW53uV5XnfCYrBi9wQjVJT21FjALZNnC9LWCA7vLWl3VLzMP4KAMnzGCCOT
t1jcKnf91svJ8D5/+2DD/q2GNf31UYTbS3dmtRAM42F1jNtu6D58x5Aw8P2BZv+n
OCeMRtiQB39VqRg5AmIp4Cs9KaK20u+8M9PTf0q9BURdgYykHRmMUYNgxFGv12Zs
zZIRENseVFFEMnuP46G8M73j4sSQmPgJ6qM82lqZMycVcX7+V75c9xoRMEpLQO9E
Us5oC+D1fM9SYlk2sgm5U9Srs+HiYsGJLZ/GqpRdSlTPJ3ia3cI/FLAXiXHS07EZ
tCFHjEgjXSYqocziCm+lKVJahma/1L7HtKmEZRl+0nZ99eAzqiJa23qC8qgH5urD
feHvP30yCeSKcZ9+2ww1NFCYR1jz34sLOb+Jut4beLQ4QY/kkxlqSbPkoMeCjiwO
295jDd/Qs7oBaOTCAphprQ9dahtjwX7L6HudXjdlUjjA2qhDXtnRbuup4Wsfpp2P
IgXnJ5VUed1aXm9ydtKB3NZbf2U22uz+t0CbgWcXPKHB3O9pFGXcsMOL0sd4J+4L
BSRxPXgepI48ov2pbMTv6Am/bYuFOtUU8eto7umNMxu0Tp4mtbi4ddRrxL6AahLu
j2dY5Ebna2UVyf3/iP7wXvGFSIdZs7YBO/Y3hOzYiVQmIK1BOx1im3Wy7TPrhwL3
7YK0o8ENAkGGCj+RJAsGgXtv1hVwfJN3TWs8KYGLySxroQYjudRFzRL8HQsydKpP
VC8AximvJqdjprkHTqwRGh8JHOHCuZCwHWn3mks7gCsxBn01/3feF40T2Ciy63qw
hc/u+Zrf7ZCXx/1giOn/MxUcV6yxpObenoYPAGycl8szEm4acolzyQJrpHjJxOfl
PKoT2QsclRgvTAbm3/ogq1n0oc6TJDySbaFm8EyrVQK6HvvbzOFZU6By3yGXzsFu
J9yN8l04gEHcHxmu01+RkUIgbLsgoE5DqOlrmJPV4snTWeWth4rK8mcygkWNxYPs
fD5wzMDlhLxaOBLNpI91troTo7Q5A/zWc/OGKoCeXI2vX5PE+Gw+bWQnzox5ZPku
9MJlQ1kvauuEaS3a8s4pHx33tQDOEgQRjoREnaE1e7qtRdQc6XV8R9YuRjyhuwJi
iro2Y6zZ7FjSFyv/BybxYKECRyCe5von9AEibPlsP/Lpz4Pl6t6UXckyZhwiIZFe
G9wIC14sXX04+JA06nvXJMX/sEaKfgHL+cCT+2Mo6cfgXdh73BbPdlvmnl2qAa+q
gp6lj+dI6EsRDfT18GANbJsKvGXHPBZ7rUFPIDjRdFL4Zc0RnDUGhvOdyIG8EutG
94OTa/7j6XfXrs5qcJcOxQTqv0o1abEKZ/mdEPu2+S6nmt4KMIfq3PQwQMOOekM0
mFSukpOfhFHFDPQzk6NyDjciRw/VfQwYqK2KrJVaNVVfs+HS25T7B56rRnbUgMiM
P4bF96a3tw++nkQULyCz5Ps7D3LB+USqjFNx8+eakT/H5PY3Oim9iPSdt6/5eoGh
p/WyiLttdWf2cFMN+mJLF6fD9/bRH1EexpSiMUXRtYGWNcuvhS+sqxaPUVd1H4c0
VLscx/P5LNCZWmYltWYnua7+4m/er6ufzt59efmHoiKDsYac1DHszbQ0eI7dp/R6
uXh2JDwK5hM+G3iQ5oCFLJc33NkiALvxWnaF4Yo3IG94KHfMpmSIzX5W9UjKZAut
vC9tz8zALpyCU88IgoIIx5RgC0wqg+BGUy7DpSeb2WzFgKkEztmuyHwCuityMZEQ
+yQsm+9tVgDj7dZWdA5VVrNi+EYkbUyJMUXmXXrbAx1qCeJVY/2Oa24hl2/MjMfV
Erorx1+Mhg+HEJoxcVrXlMcS3nfpEv/y/+orXxVPzNVcujRHCP2xNHrEuJsLF9/N
i295LHI0CcENZjdKzjtycSfbxRgXDQKcuNlIRHWNaLBH5PmSdHpVuMncHj5gtSp4
0X7+22Vs375emUI0zfBEtu7+IaYHhHAXNBdlCWRzgsSuJD9/LKKBL/XK5At1HPHf
xzYAmnIKZQO/BMU8aaIGyWqkOgrWXzl8/SE4ka0oH+1CW+bJmmRp4Gl+SIj5HQx6
DSlo5RJ+taLN1Oa2coyVOvBcF31D/BXk7hMKADDrwDvsDppF4Owh76A+FFguVrI0
d24CF47vkWKrE+vhQI0BWxR9Hx57naqEz07eJEIORkdRbqJfAaZnF55KMbBxqAHh
XftyOghyDCB1tLLs0gcZir9SdW+wbskXBXvQDXLwWOA8vHMqeX4BTXOyZCTXlJqf
MBMTryOFYRw8hsVTHjrCirtIfMj6lrwAVADpc8RaWyOQFi6D9ZhMbFW6v0hg6SXh
MTnCUY5Oy/cxHgUjQBO4d4lkJB7YKlAayHyNWyW+u4Kyppdr7JnUoq9/ubPrMuWB
WsakraEapLmn+zLBtdnKzpnNVN4+DHxLBQzvAQ7/t3DxT1BgZT8up5pl7HKub5vL
kE1zAefJmMijQFiZTVzlAvUIbSYJJNMzkHeyGbLendGi6m2D2G9G/hAYaY5kEHoV
jQ4gkqpMMIGSgZbLq3Wu45dnjys8cPwSGI96GeDiq5vxFLTJg6tT+9zPHgI9Xwqx
CONKVD9HhUmsr/w8jChAnlPuSvZ2cbft4UFm9V+bjl5UZvgyM9J43m0XgQ6Mut4R
kD3vNx3X2DxB8eHV5V55OWeb0Q2LrhSrcKUmYLiSPY9lJ3chMk/jI1EwYk6qPlMc
ZBVD11qCZsPGYSotD3oCvVZ8wWd0CVvaHc6X+TpbQcmvQxXopm+qx05NQejzVz4X
Etrt8xkZP5tvwZirfAQldg90ufiIoNTUdmW8deB7G2/MmKJk4JDq2F3Na0Oj/fZF
n6dhbD9ZoVDJ2UJznobqfPKGOAa6o2U3HMv+S35kcwRkKWpDTKI9kSsHrGdiN4j1
K7PDjmZlKNuomK44s6awbqE1XC9gaim2/l2Ui9AclNpNsOUDewUHNt330XQP2zM3
vOjAavSr/ihht3KaHspfqjIdzUC5G+LUeF4mePhF2nwIe+2DfFW59S0sYGzqg1FP
KVdcvgCkH1MuGRdSUaSPq8Tjoc2Qyb2CWzfimVGvnKLTNluLa8k3DbX+XumG8nrn
URXE8CSiMv8iuk4T+1dOZFeRsud79Kqtei0bIYJpOra+p8bb6wQHpyp2fQqE38u/
geIqTGqfDH5/fjZ7aqmH8XL/ecHSgxHU6zUnLz5tQp576Mg7cP8bZr3wtIDhdK+X
jPvTisHPuFXMoTz1Yf4ogBNzs+Swq+P1pZ+Ksw7VWOUtAnJY29PI0Ed2Tv4TgwWI
GrBxT1GqeImr8lARpntA8PlYLoWKkwuzsTn4zFfq5Mfoa2BlOri6ZNvWovXTa0kc
qLbdcA0p4+mQWaqm5ebPfvftn+QUyARhf9c0nRVnc/00PFzy11eJVoR5H+gspNYN
+faQiHzIGJLufljyx0RouV+Vp6A1dCq86lYNojKT1XXRETi54bhg4Il7SYxbno0a
LJQ35zwTkban+ShZAdxDZlq9UIUKkV7wSOiH+gbyydGwyICl6PY7+XJ5eHl27h6+
Xhdk2akxGM6kb+ZR91TNH3aG1EbBgamHm4sMELsCF63l+8ENCD233G7qTxTyTWHI
JENEchtjFcDCfFf6keov4Uejd2cNVHAsIhruW4r/TQmJa4Qz+di+wWrQMDXHGtC0
c8hKlEZIvQ3YFE6XnLOhl2ImbEXVdQPbiHy6Ipj9oN1vmAJNyQJh56/uxYuVGDO0
eKy+kE7jfgMoYjNWLa+c+CLhhI1gqi0zhuj9S42H+lz3V5NdYMzMXFc6xhyHQwvt
XzxIqtxj7pAbDpsNpFWyqIivGF+w98U0Gg5W5C5j9CCXEGQMIqKAZNwVOwUNAc8/
8ui3p1Vvzu2K5ELvcVljCodHU6aaXkH1YxakbNbUPKOFyYmA/5dmoZR//DjrUhhD
cbb7a5PTTVuuSViuCBUGo2TiIGO/YmPDlcDuvKHe2Kr9QstoIvVcp8M5kI7FhqWv
gH64jBd3HR715C/57IHryZB36pMeLmLekKsC1aUhVsHKbsyuU1I1KCmWf53012sW
J+TSazbakPXZJ2f6AJiSspMuHP+ccvbW1LQQat4SpnqbmiZUQLQbDvIMHj69RTMO
5zI2DfjUTpD/LaNxeUv/5sa1y3VdLy2dyEK1xT7YWZl9VviCUjSase4XjnzWWjGZ
w65KqW+uLe3+FadWSFHAwI3/x1mn2ppl9asHRdoYgpuVL1mAY278kuODFTLoFgp7
R/JyTkZZY3uXylvCaigvFls2LEs9qtuMj94eWYswY1MfBI1SwM87e7IM8SrykKBp
4/j2cO/TZF5og6504Lz+QZJoXTiGrQTk7hduE4HBZmRxm7TGN6nAR+n35HPH9veZ
PmjOBE8uXr/6WoPS2jZ1oV85Hw4+Bu1VT0Sb0FXQVI89QjyeWxST83X03YtO3+Ye
pDF3OzbV9E+oZdlx+kswT9t3fJCPybuBhp1Gc382sDGBLZDhMyFCkYDbZeYtohxk
TG/b24BGtzZMuYRf7hS2weu1dR6uKtaEg20QmAUfI3nz3oY8nS6+xCzooAkB7nLZ
oNTIQDmp7ihyUPsnxtHotQiNit+O+WmAkqX6PA5GnZiNwY04D3vS+IfZbg7PSZoB
UrPL0nBiD6a27+GddNsndmuwKQnFZxHT5qLgG10SlCdE4nT6HOGJvFzULGhlM+H1
9II+EqnBhUPVSRZzfBSBfezRWFx4VF56jrl6Ws3Kv6YKUnjexCYqqwM+rlWymTbt
YnOCIMON4vPMyaTF1JfftLdUpEAikAd64wjEXfBI+Wxn8ajvTuam8yTHXKPaNJg9
8J1uIOIhHw2GumM2DhwstvWMKr/9IWZo7lzTO7BYQB1kzT/HFHahApi7Xygq4qIg
vTGcyskNJj8/75ya0SLFSv+r+ykWsKpdLED+gnmfVpXsMJYbNs6rZgEWv3RP89eP
r1uc38j+Up0vR3uMlRoEt/QVQFYsWsTkmd9OT8pvCu2FANbFXdBtplcW5HrX+Y5a
5tLd4+rQw/ARceOm73ozeyC8vyz/eXJ+b8w7u6nJEEHRPHEc2ztBcG6hMBl2rSsn
NLUmQFNrdfLI58RWyERp28Q6mHs02O4OdiHdSPf6lE5Egid9eIb+/C9x18aNScOs
jQ2SY7szbEBlebHBoi6YnXgdB5HeY+2Z9bTi63QMJj+XZgDZUGIxVoXeWmTFS4dk
TuAjm/j+0zYsauyJCSs2YEhUzYTHvHmlS8J5VkcMBVXZ79vd5ay6OwQ1kuEV+EPU
JJZ54vrF3HXGibS5SOWY9mo0dRLhiIgV5HVtbU97KWj+OY9puJwivPZukq9/uLvB
qQaRYPZFr2MhiPMDVjLgCM9d6ibUiXLg6vsFM8T1ffOLooagEuvCEObK7pNZ0FaY
4ipU7jdSPc0tLtK5jURXVTsOeUilV77PGjoVcuEVv4wHp0HZlXMHcM/tdJfHs09I
uuYp/rS/ORWZ/oxaQ/p3xzx5yVhygZQ/lAtGgJwluMUQAf+z4bvhVZJyEbj3DP8i
+PkwE60FscvmDum/eSeOfpJ/Slu5MO5VxTjJe5+4lBhiz9bZZH9b1GoKOSGZSajk
0G9sK1VI67PuyJ6gnWS2oxTvXaPIsDX2AgsDN8w5h4goOy0HjEuuPqdIywFHxJB1
GlKqlMvvXcHiQNinbLhvXDB/V4Bkk5en445x/pIKXWlYcepX2YhlAL96bVTniDKx
M/fotW4pnje1gdW62z2N9SAGD4X+Rlxvtcn64QQH4enLbZ9EeBikkYJsGYkPtr1O
DLlhyVevYnRbU9Nuh6EVGFLgfugvNxMRxPxmNz8ik3K39xnoKzaH3YZcyGYCWgTW
fAYKgiKiH4yzqczl+8LKB7NZpa2MC1Sty4lMrWMaxfK8HJwU9HqQC9xnkKoczg6h
FX4Vrxf3SbTRolaZx06GaZoJjAc0lzdoFSxhKNYCqXKpig5/fBujtYh1U1UfdoJh
VMTxYSaEwED7YCMIx/xY9Wgq85MyatM3yn0EowYcBTJs+7N4n3Y5J/5djoegriIk
p2gdQc8doEM46ODclPmjjq5H6AZIQTekNjCJPc8FvniSSRqdD0t3t+7ImVkN5fD7
hpAkAXa44nbfeH9YgcyX4EbTLvzLqagsDwD1hqoWO2Vj6QIzWYg4watuvnB215ZC
ayesdA4ISE5g19WXVx2OF/Zb2C7OgDV3xlWtOFrG2Zk6bJsE47uPZ/4Gaa4eRd8v
+DbsIaUF496H1/CUGnnF0e++DLZ35KHEYk+aCgVzYUqERONBjwW41fRbc6iXi9ga
oJlaFsJz+zPDrA9bVpoWodQ6JflmtqCvLXmBR6I6iyyBytIwF90tZ5tIpJg06Jij
84GAcS1v8kd7uE39ieOYGs2UJUN9Jbu5rm6kaOhxq9LjKmQYt5cF0xnBWV3Zg3+x
0A5JFkm8mtD9joP6RNtlk5x+MXhcQZWHdSlKd7SqAhSKTScNdPkYdf2hMSbxM1Ht
g4kg38+8yxgHmcykqZnVar1buC+eK6gW0N1RvSuwwqJt/dH7u1shyBy3GyOR9OSj
Xdb3MIFhlnfXcoFHwRntmMKjX8z4NJ6ToJsUn2C8LNcYT5r/5aLtchPnaYE02t9h
KtTyAdXHbDRGRCK707xf07jUpt6CV6xzAPbnwQAo+wzBI+HzHQA1+K8nNljUz2wv
utEiu8tlEgc7HyrO8zBiL4gA6DzGCGC4K+TQH6I1Y/z2qw4X4K7NJVYncXtv74Q7
68gzRgQ9AqyHoJdVLQDd3l6050VAsIFdDHUnVusjFKri6W0EiI1UBuE4L3J9zDfB
84PD7+tERDSzSWLu0fNatqP5fD08mhTVKBYZea4/4SomvFSQ+ZK77YCGAOVOtjMa
z0t4896aYX8y2An7VWlB/nFlLc0gHfv7nv30yXFqqqSnEN+gUEkNrZSLXfHrSR6w
GTykEY42UMLKb4vDYD53l8YLRRE6zYK7NP6KrSyPOcBK4xlBFkQs7ElFrhw/n/Vz
DCb8bW16xuleVbmKKMk+/RZFEV4QY682fpq5w8uFGV/YmbJD5g/+3fad2ioVRjHg
7bJEF46yaVZ2TdtDHrlmJHGFLx/Npqtt1FCXDObTQnAC8vhWtog31U5a/i3TLCbf
x7+SrfCxHI/D6rlVkZ1dzy1xfaTkupZBrHuhfqzdtoF5NbnuGuOSC2NFbHszaMbf
G7FgGdp1SOqcijMqyJhTk3jqabsY3CANLRwhtgKN6wWSfkH1DsVtFPudiBMtFAbP
AHNyry9+Ah/Q6GdzPdO4+wCGSxkIWDEXTG6seSlhNHir1d6mG1+aQVUp8fyjSv8y
d+7CFshsBSWHDn9Znvxv3H+xQPKbz9LS+uzPzyu6pTRHj1YWcc9Jxu3szDZH+yfI
pMY1oQE1R7r4w/o7/cRRGHtapcRb8dyJSVrxUDiD4LvR61vZ6pM2NzHLFJbFyMTK
b5eCah//u0w3XKcAqZsOoTVNkowDviOtPvt1Lxtnyqvv285ufyxWfQbOA7SFnU6h
5mLzpH3ZU/pAycPO1b1HNO4JhWG56vm+4ZBo/QETN/ArbfTXt5rIFa22kLbQ8GtF
lzgoiZNiuCYfsr9JbPI+Mg7c+vK42xAFTj9vQFmOXJNP0xY6iOCrBEGhlIo8WxA1
FehEwnMo/aMr8fm0cYppRfWZNrbs5zvRoxMXkAwp1JhyWiPSV56DQzStjXItK9fZ
XgrrJTI10bT5cSQzlm8N8NxQiRrju84+NLAHacSG4w2FjykR80B+nb3+tjdtYO+c
vtO3qoWwRUvegzYhDthsVISSjp3O/vhR8iOE85GAH6c5OgaSoC2VJDQXuKYB0+Cw
taCikA+59iO9p12zah7yQ25DBmi+y1rV2aFoVDG+xkfOxBMePAeb2i70Qaxga2Af
JarAHEKek3ktwH0Bxg7QxjJnadKVEzts2GXzEilOCTRfwmfcw4bk2jzDG0sPi1sA
ij/+gfANg6g4J1zunrkpIIWpTpcECUF6crNi3gGmxA96w7ur+hTTNakVFZ2OL5uH
U9TwRVOuULYc4OEbnmEtEUj0edMe+tqkZOQZ43pI6HkLSaX2r5x2coeTHmdpSDA5
QH62dtQ0RRTRrItWMaLaSvbloB4ipMjTHg955mmhcy/hrQ5x6QWUuI0qE1MX0BDy
ZADFobmkEtv48fb+CGX3Gzvoys39TMhY8I7flNcSUiGGaChsCv1V4WNuyTIoPkJv
tHyj1OLtzQBTmQr2RYdYySRgY8Sjbmx4b+ZgfrG1/H/gbgqgBwCw2hgWwyaMn7OZ
UzHvIAF6bvcyM3WBYiaLQjxi7K7qz/s5F/XRVCI/P+ZRSYOVBHvS/P8mL+MASt3j
RCI6/LSMpEtLNWuDxaVPtv3YuES26X9fdaj9O8yqTGGAO1Q99+mfdS9PMX7EpDFM
qRhPTMKcZ6sFydOYzq6OIfbjUMO5N4p5nNlhIKB2TeU+LQq30vFCL3Ck96EO3jeH
kcRsholSX9eOJbRewdT4LvQXTw6Wzoo5eehY1L84IddPTuu8KHOwr4WS3jXpnyGf
mwr+9QOPZ/jPnr1IA6dMEgk1lZ/0mYAI9vly12vWBMvHFsmw8iOPcYKAoVIUVw2z
uFwmPLjn05+6Sshq+bXTqSaGjzJWK1UgMeeXO8QSJy4ipI/9LZuljBXM8ZgZpypF
WAduCJq9BN56xH0+3X5XiNeaJRr3oHP4R4gEjsu0KShauE/TvENYFWbDYP0Slbpz
rbVZF+mHqoSyOoSWqz1v0ptYVPCY1dcLL7VRoqgny1Alf+hW8Q7ALi+P3ECkSRpw
5iYEMdtaxQCtwlXSyqua/jtXuxr7xQPuxbumLJQzX1TLyfNQcGAyoxoKNkihSG9H
HrLye/+qYSvTZ7vFrjOCOfXqM9SWcOL7MfS4tvt66JkEeAdVhycpN3LptAgbHtsL
bbwMa8CBgDBW67lRCkY7cE28jxKKhHb002YZ3dm1ElpYCFA0TXHkHXNbIq0nn6ba
OBDAVoDpD2XU6I6SJ5r2OCxbb3z8i1Vi7KAqIYi5YZXZV5PVws/bMKXPaOBQPkIK
jWzFNM4VNUxJXZTQZRHZcRmUkceYfMBw6yyiLRbQC0Up/tbW8fmDJO7F9g9q1tmf
k61fvpRO4i5ehYT6Px5mcGvsRz0c2m0mSE9kjjVMGN4myUJxKpsTLfAka3Uhh4gz
tDl2mWLXhLfv2JKX/aF2zIsQCZOG7TlznAyIO0lNemd0CcQmB80T/fSOLjLJSjGW
NunnfXcVV5knzQcUrImENW2SejSRTZZI43M0hqYAPxAnAh7AC4056IyJ3nJmu6G8
gWKljoIFbLmz39Bf8tzAG86btnJ0LbFBQmkkszVbgHejB7WeLtTX8KQPgnnHwDvW
MFtqvc5GwRMMMvgLr6ggjATS7ESolGrkXQtmqEIwUpV8oy7JaM29O74TLYuMb9iR
vpI9mVWt64pUez4zTHE9Ams40r0Ph9lSrLxWvm1saWQzqn/RnA0a0y/JPwgs2po5
ZvfloueT4lSFoymZPEqhKXNIc5t9MHzyiiqNtpZKMppLBZYKCcDa008sZ75TFSit
q0glHacN0hodRkQJToctqhmrfKVd1869LC/pXL0CtC8biib2ksrF0yUnSgCQoFAY
/5IOPQ+kA9JpCLMJHyd7Y41792CRMrirzLJGboFO5U6xvy8ZtGbCGm78NC3LzvJa
zbHar5Eg4nnE6/81HndwTeNZdb4zgkuKgHwPDfr9lPfNUJRF+QPY6qPU84JDyxPv
Zya4fFB8crprUuCeWaiA5jg+JXWC/IL8RGf4WiC8UT4+UMh/TAx6pWGXVRvrQ6Jp
z/2omGQ4ySB+7q4mGTvdKpEKEiLl+MvulqC21I/dQBDqzlDgQEdALRT9MorvHele
OQYcSM5cMPpxjDuWGGV4s95AvD7K2S9rtaCyY4pDLNewrcD3CTEqbcF0WMBn65Z7
02kwZcrVUnGyKlqg/4CHO3lR2isyj9G0tR6Hch4Dp79qz8MTSnGBZIANEI83uLW/
NiwZnlP3PYhzhkNpXL5exqKI4gupKGYN7DYgjcjGR1xfbPHXVyHnswlMx55On64w
bLAR54fnVjq8OadJmnzL2nic1rO6Rw9q7l4W3DJeJIcoh8QgYsa7AVbqbovKkjcg
53MPzFLxwyLWpbWICyM6HfZ/scfwBoWoLu2TDUtuOyB3kYxAyQL837m13mwW8Jw0
ad2ITjfpjAAz34GWFBPPgbOsFewX5ZdJx3YoON/IDK55TDxO8jd1oDZakud1cEnL
bEyNpSWLSfLIkAc3vJj5km2+Q7Tv5qN5TzDLYakHEo4If9Ee7nySyGU75Nk/Qnp/
d0vjsGt7pU3cpKnxwJNcgWSfE+/SpsAl0Npw9OxEhf3WLwC45236waXpUaL8iKxp
/avppyM7Bb3MF9y37Mv06kVOHsC7wmlVyzQbqvQYFqSKxvfrnQZGSQoVFu7RYRcR
iX/CO5KX6KO9uUCEwwWlmbWzyPnknzk5EyqA1voPh14Bo9IOXJgEGD4fMI14bltI
LNncWMzityaRdLCLEL0u4HQjwqhQipPG9tYXXYHyI7n95r5a9HD8IfrWQ0eAyvZT
s5iwnJWDQk8081pzYQocsGdXNqB2xidvWDadlj8R3HelKlLB3JB1ynUs0DoacC2O
2wziO/auOxERrGmXoyNu/5lKuUjmMBdjYEYSfFhz9QYTLqqax6NZP+OiZEP0sVe5
9acLTKuHfL7pu5qZo8waBasEOqeGC0VZe+rl0IpyVG0qmrxSOxhjevW+e9SnbjkN
+J1W72brdYYSdq5IFOq6kfDY+obHLp8iTNnXzfBvVDnily/pUVvjW1rCInSdHIab
656MGnEw9iUqc76S8twGkKjtP2TFKi9+r44pU0WqPwE3Ju+RIAa8pyHwLB2KmIJ/
SbwdYFYaojfBwBUf2s+ynfH1AB4qS+eDhManYDPZ6YCPDrrS+Hu7V1NNtnWhCzQX
OdkaTByrDjh+A/mhh/Lb9bKkd3H9CAKtOSbZzC66dM4+f0glS92PXjpgbe4FB4BH
q+eJQz/+T2i1ltoitENGqjuSotlG/n7129CXbGNoNwW0WVYswuNKdvTut9iOwnEZ
0uudA8v9AY+gH1ioNBRF9g4KxixdRQlnuxp8BfCXIYrX2O9TYDdbFprfq/Z8o5Zl
8FG82CYwn2sUW/pysH8fGIWtlOERtjXCDTx+C43WAxgQwvZ0LHoRa0ZI/5c4HY+q
GJeGaOFz85Z1Mrlb7Xb/EST30Hlc0HwPoiL7K/EmFXbH3BfAl6y0w7mhM65FujFc
ZR/UTNUfEyXfD2u0vmF/xQ/RTF7KnJpy09J6qapbq2W6s3B718StcI3B++G7ZYyZ
Aek5zSk8manWyIJPi9RQ+RVVKaErKstaUekvbft6rCzTOTErYjHVaQFUt5v17cpn
L7iwYmuIZIUfBDo1JCnt9ZTfa0bx4W1pw6o21xyk6ZhIG52HEDu1ssreC2V/a3SI
BgFsEJ4SXpPWvFwYL/u7Aq4gf2yQqUT4tTRnW05kMMK7KPivup+dNKBxBMrI6AAu
k/uuMtPVnR2erNMoNs6YbQ6nkR0X4jVmNLerqve4QK6Gr2XOdxj3vpM9E59SkfHP
QAfT49h+lSt6/y/rtUMiPsHi6Dkr3soICD7D21lApQMYCXkuE8eX6qVJyW11+W77
gYMXmQGZ/PIvDuuADtN1QLKAGS+nah9KL0CTftEmNVPy2LQjCaFpm2brbtOkUjdc
DmevsTJ+Wl+r1+7+omBtMN1OqL1t+/qKiL1jc4Gp2hx9X4DbEfe84HV6qpGhR1cQ
GA1A5QaMxdCk/OJwpgEjNwKDxf300pccnLdmZ8+crt8bjywxjVarLXZahi5iuSrU
wrnGq3HNqOJs5VzzT133xe6kZd9IHZqpL49ILT3P49u0WpTGkFjCrlOVweh+ypPD
xgHlMnsUYEYJv8JyF0o7JA8bkzVign6wfzmSqCN1TkTHyrsZbzV2wJoK5chcErUC
wkoQQjHombxkRcfEIgc5y5/t1RkgqE+IdyStQjtUqGHIrjX1QlZ26qOUUFgq2Sql
vtxPpaowMpbBfi9T/8+rEvGNEBOAA+1I0z2qJmqUaytEXn2Zyp/HgJ7l0dBLeLUy
C2sBlJ10ouHU6XYKo3oump0t+2trO/Ncr+ajyvwO2590ywDhzY2ONozFJ7R2TLvj
ksLtVCh5iD6zCc+Rg9DwMmEI1D1Tyg/pUBOmyXX9dYgIyYBdpbnoxIS7HRHaLb8b
Rjw8lFT7VHnXfl2GwpBouLo1uSAhYxdCqnMurkywDot5ukCWzAW3W5biAEyxFOfN
gvhKt6kGxQVHRZU57f4xNYQxMj/8+oXsWybQaylWp21sf5XAveU1dGz1Ulq/kELG
8nVKuZzg/ah5K/EB68aJwFo4Nl9Jw3mu9jGfsB90DjRkR3R6EbLvpWj2Z3pmI9o/
PFeQhCFFjh6wkh3ODzIzz4LizpbG0A+ASTlHNdwXfg69eYD3eBARk9mgetg1qq15
NHQ7K1AB2yY2HP1B/eXTdWYhkmL9o2P3aHWYwRZG2Q+gEoYBlavRYd/hozyUd/3v
po51Y2X6qtSbKAG2/urVlAubjFtTqm0gDDmKTGGVVajoZPq00bkJoVfGYkWA6d56
0JHsML4p8iFslwGKtRkc3lU4SZhHm0hEWD+xokCoJbMoFEnIGeDet0+huqBYZ0hr
0R3sXN9C2ZO7EP/9aL3qqsCjEaqyGBc+uNm/Ijn2neMAmIC6NDgZA1D+mXsTpxef
2FAYEO9HKii0ugDnKTXGV7O4WYM65D661TNXa0uQmKKEv4EJFvyY0RtL9nBQ0had
yol0rdJYHWrtKArrm02d6hoHX36IQgOM4I9eCjCpTqjVt+ly3KrF5zjOWGZkztUT
o9pGvO27W9PcD2YxS5u3zW6LKMSAU2wrGgFzsG8VEcgeRpIvBLJTl1pDdpwL2/Cu
db6r5/acSGBLWkVl6+PbK0tJIg/HGKbYWevtGN3TaqD8sDvuMgOENq9qCcZKsHbZ
b3sqOYSMPhFYtBf1bbx0BC0OPP1xhFXw+mTmqGc4e5ZiUge014PkmfqpHFX/vYAx
WdhNKzVydYVaM3z9o0BU0b/vrh7vNJ+x64ZMOTmqTulANx7rAxCp/7+7NQ702ptU
ZQDePNaG17CxBfN4LBOQrNpENrcZIXQY9G+q+lRqZMeKLoRvDi+Xr6fvzcCJfJaj
tKsjcUDEv1VrnT40mpra+TSbBQ9BilZW2xE0N/oiD9+D41GSukLk38ouPFIPXNnK
Lqvp6JBQ94sJpe2oyVDq2eaX0DPizT/3xUU4lOHMhwbbUzLiI1SWFtylM4dO4Nt6
TTgCJOPutPvvbdVJHYVnbfwrmqnkuRzNhQy/ctLxdNn7oyjqDwfiEwyQDhqogkpc
dWqELbPnI7vqf3O0wwUiBUR10NhRSs8tn2Kd2tJ0rxs//Oswbm69rz1YfnVtKRCp
oyjEaKSglC22xvXFfwLi5paqTVe4l1XpM7EEE/xRCiBR4Xwx8rrAPcE4IHFGhf+6
iyMPXN860TCMrjueXXK7RbkYx3ge3T3ODatq7sVZCWUZR1g8FXvVRAJkZAMLOT4Z
+NBnwpE9/i35/AAE6paqt/Wkrc9tYSX/Q3f6FCbjjSKd5BnOsN2q/wsN9VcWHkgF
+i+x6gIsK44INpCwUO8oIREOsQLO7MygL5M7ZE48bvwhVA8EzVyh2LEg3QfE6pmE
3XqWBPHffpb3wztRRy2sLl8/pQy63IpZWI85W5xsdW/PBRzhY54oXv6xES7GyeqV
h433RJ6/irxSY+J+mzN8j650g72V6ocMhEaiYSQjQUBqzgDFYWyrQ7pQ95c5CuFp
tKpxOuko6PDdcXlmVqC6hpot0uUmlvKhpCa0wjFrhKCW1HL7roC7xqiFEgkZEUPJ
Bui4w0/COq+SUKsVLAfodHpx5nEjXmQ4T0urcFshoQ9mXv/9ZLtAcDDtnEl/WXfH
HmiAniqOdxejpDDd56MBiU90Ns/5LGWpRvzEyNYMY0A+JP7M7uRcwEMwBSxhWiXu
BvTdWbGdiyO1yW8PmC9xCGUDYO3rrO0hS9ewUBeU5Gyua2jyZ2RBpWfgSC8Y3VbF
vUSHr+Mg/3Fe8fO+jjnSeGt3XWUxbYjQ2Lk18N7A/wdo6/bmO73WpkmuV62UTD1E
IxUO0mWODKe6GWlZy0rQD4mEiU2Kq7GYECg1d6bS+8spUXFlcCyO/RECl0yr+NiC
1MOGfmQq9StvIwVRk2paQfjpYvo+gB2A66/DmyJbPuqIkRUJGms2/xp4LUR25OJV
teB93CfvqQDIkTkpnNqY4WF7XsCSnvZNheVCXrr6fDLMQGzyte4+aJW6rKzB8KML
VnI6Y7moQ2sSIn8LMXsiSKRws982FRywb2H60rnJP9jaAqx3RAwTZ4h3F25r8tCQ
5e+nBof63X8oHbfzX7l3vH/v9nUjiNRv6/ow5y+jozELV0rjFnr1uZnY/JjwPJ5S
RXueM+LHIQZpFw7ZbGJgZx8TmV0ksx0gi8dgOfNZ/tW9dVEemTvm4z5tosQbDZoQ
mINSkTkLPJVXSLrNyGKDxRDG/Qim7xrRw5IugxtZaDbKhR+C8/z+E48/BLQ4GlUM
Adfzg9qgKckM/aWPH1PqOWCffYzVfIy40MEqW9pQtMj1CrrtBpw/vwrMJpBKE5VK
/Jd1pkwi2bOYCS6hmyq/7YdpJKWM8ldfU1eQYG7UFyk4iMbUfzePDgCdRBFZwCDO
2lIU8YqsZeOygB5TKn8Y3XjRXjkSZwWL2w5gjckZfBkQD6bMVulwSwCj3FOtDcAK
yp71akIpH3zNPsQ0GeDpbK5ViInBaMRYiL4Ls6qLObwnHeJdRwqTqcWGGBPjBOyp
jDWUv1/w4dVQtVbb2+mXls/iFfO6F22Yy19Uj02tA9SAPNkeZTYd0kKWdhjpOAmW
Koz0EWi6yjCRir/vNqiEOP4W/vNFQnT/CiRh81GOlvNffDiQX+dh3UprhwAK9B+L
GzOKjH7ZSNnmPG+kemco+TuaQ0uuoXwGFAZz1HpC5vOyJAcaL5JQcloaBthGq6mD
7Hyh4iAZVaiR0LsJvG5Iyo6tcXSE5kCihET1fmCZS37OGrddQTOIloRR5NEgnOEB
7NEooiwxYNrj3ROKoTwFcVa+QRTNK3FbIBPmUGcJ0YZOf+ciF7K2U0xSJpJvzTce
WGQaI56saTUwH9dgwueR6kEWzWOB1+4Y8dy6HY1eJZ1O5jLgXHR2xMC871tmqQ49
2kpUhGiy3uJTW4E8a38/JPyCnCW6Wyq49lpkKyipec24AaRecPxO8yq9DmMTuyzS
H6+6Nq9pnyCxYgq+/TY2BZbzV+SWsJna0pI6rFn+z6QfuZzm9kE3mEo2B7agmJNf
HurkYcBTFfzS4hM2aTuYt7ijqptjxvGnM+KbDXrpDiM8hI3PfitXOhzBClef5jdm
oeTdUHP+jN5aeMvW59mmHqT7moUy6IkLNctxlBx4cvnc7ddOukn9DFGDYf5sFrbA
So9lOGbZ6Prw7BIZ2/RZDRvO6znXrmORc+pfm+a+oMkdLjV6WE9EiEf+BMJy9ofl
+RmNRcyB3vTW0C4I3eqgDVK2avqQQUxNKlmv5VUt/4qKg3FBTZMHspKrGi+jX5Ur
E5f1YwZ5Nr66FG6fxNc25LJ89I2R/wEATB5wErFcnuA2gcSvHLlyngdoukNgi+eD
gmXamCl3XWeotwq22IHFmN3NaJW5TCCVOsp/nT+b6ZeC2vQYijj1m9gYL/AZoHu0
YIq/ICPcXDbfZQ2MbAcgiJMqM7m2252yGJ0D3R9i2axnjqK5pRfGa7f8grQpB2hT
KbYuDxPesigkBmkHBrI5JyyvVlfABE2U5E+X77Q5f4cjemYs6rX8tTyX/x4SQxKM
Zf5t00+8h4j7nHb6dDjwEq+VY9T+RyuWOOQtcMIyoHa87mfwTdeSrnMBDUWRCPfS
sS7s/9Y0jaTB0IQL1MwirePfLLdkQAvSVcHuYISveyvAsgessYX5a0MMEie3j441
Sp6PKgylZrAZvD5HQ0Uj3HxkyAy5JaaOJlrqqlLuVEUEIeawao0gn2FEFmf7Qq7U
g2dKNVwUHGf/Gy27nl6O/5GpNzLfgHAe6Njdkqe323u2B5iPs/KjUVy2TwlD6axY
wyBH0iQAIdpDxJgDEWtQga4EnZWUkQzNYNVCEyulVtyZRf6nSdkhEz57hsWVqqoi
10CUpsjI0Fn2iJf8vcnJVk3Ed1Sq6YEEX3/il+1NZvHRNPw1IbZD1pTQuNyVXIPB
bVPgiiWCtRLCE585hj0Lr8RK3zI2N/3IO0VrnrHh/fYYY6XMsNcQZDPmjCGh9yKZ
U0aqwGdke+CFsKgvTCx3kIhpJEDh1QzjWYq9eT3YfuWyMjiofGmFjTLkIWwax56j
AcrOC4zwcdbqfojQN8axZ+7alm4M7dV62K0/T+bntARCh3hIqnk//pl/YrvqNry7
nE/YcNRBI1si4JDcDZxqg+eULAFvv/mpj58EIGaf9iUDQugO9rdwOrtBV3tpwiQX
WMOw1rb8ZLtpX6NTG5jsp7NnlDYZWTAeTKUDhdRgGDvJZ4xN33q2v4xBYBPNVarH
rIN+oWn4QfvRD7e16/eEgjWs9mmLPBP1OU9y+Mb19jgQEo81n3Ksuj0XPsVsIX/l
CuuJisQF56noV4Nn8/dEXUrmr75qk+cR1J8v1MbAmct/mDps3m8B72r0psOgHV9P
RK3P2jxH4EgzBS8i0wTDYRfeon3L6mxNfWxAokYVxETrVyNZ+9I41CgLLJWBmxUD
HZ7hyo1WMJveUmSkY0m3qRfAKVaSn1q9m9XWckOL+uFRLkN51/NzRBNM+f/N53A9
mB+RrYninaTY/afqvJP1fqzswoJP11bwRS+E3ty5BnC4dWmETQ0XiyEuTqGuTc2o
DWVexISnAD14D6z3LvQ7oQaJ2TstH46FPYmdbmsaTJ4u1HYPOpgUW+1L3I1AX3w5
c1kMwBh5+/UueNSk6gBUtxeoDDBLeCK5bXxDRQLDyhleUdGet5n6/tQ0HbEsneWi
N7gCgZCiA793l+HlIWeO8x2DXSGNy5m6aaAlHI6AqtYWuagmXJ34GswPnj+ol9Q2
ox0jZcFWHGX5SQ58GG0yI7amMwNJalKIcZUxOnsgSye5rlMEJ9Yk4K5h+VarUSRc
XjPFP+4MAHMexks6lXU4ICZ68JTxGW7HbTakhn607EDhthLHBMWUUY0LvygxGH/U
ZGZSy4sOEK/lYvDcn5arYKTqRfZhs5bZXpYneWUUq1UUD2OxKbGws4hrjj2ITots
Oop34BcvnWNZPa0Q3Ac2m9EoNNghqhaYIau63jxy6SHCqhnaa5zc/2Qq4S64Qiv1
ErPm3Lh4F6QhGRpo1WMZY68ySqcOQX1f66/VJO8JXLOQbCF3Lqqj7ARsTU9LLhzi
NdLJtgdnGU+FiiAusOG0b3VFibTFlOzv01IeyBpBMOn2Y4hfHmmWx6CwB+xzmJg5
5nAKhczBO0cW4IUdrId0+0S5aokjjpvzr0/jvLHCVftr61GWQn6+3mxKuz4gOMx8
34tIF4Pysn/CA16GH+XmDwqZGCPdBWTvThMNAXQfshBlLdy9uFmdmxiCTDDYTC22
GlEkboGBoGRNYKu/dVqBoMZ8gjosVZiVps1nPWDOb0Tnop/2hODyA3DHUOCQ+S3H
3gVjPl3ia19awaiimnTEto2RDLKIMDYptn/3UJ6UeBbxvjYbyQQT6vQ+HWLrsQdX
f1+NiRwWyfHp+R/CQHrR2fzsXJ5t4W6eLlcmy9QenyICxcyGOzqS+Umj4BzEDj7R
Zmd1uFSysBmRgmrYnS9ITBQVqBfvvMm77SAVB5AEOvFHDTP4ZeA06siv9u/EFBCL
WgDCrUZ8lDY/2x1cZwrot5xNqCsn9NJPbenH5X8vIzgesFIvOIXExmIeDn/gnFB5
XrZVobV4pEPW/I7P9aoyaPnYI3dR2uf892twOjIh8S1g/n7BgAUJx0lliGo9vzBs
3e4K0n9YyDvElF6auFl85JUVuLyBw5dbJbUl8NrZ5AD974MUTuC1GTX3yQWPZfWC
wl4a4z/q8WJI2bLt9ts9bLAkMQ+Z3E4OForSDyZJH8H3zMaYcG3KNqeh17+naWqO
ZuO3yXIzu4ZCVKrQntw+vnfvAc0X8CL8T9SciBnHX4AoZ7al3b0dfZNsoHvAHCWE
l719jnpis+TXhdissZ4QpwrLlWKwOOZeCkD2+BZCNxiGXSr6k15ocwSnNH8Dt7VW
iPdnWeeBuis8/J4n6/6VL3l1haqsk1NfvXzkecrQIE7UksYJSM0PY9nM/LlN8rYY
TSEqATk8QDr/HpEKX8m2AR+DfEMGYKqzJxZr1AIjQecFb5jCu0NfFn5+6CjZT2Gw
xe0OzdwJS/9ovm1hqAEWRSxXcb279tc5He8jtGiHngyWfRMN3j/mckOdNlzPXDjD
optlspOS2bhisCwcgx/3o8DX7+293blmoihHkUHtEzjhb5b/H3awevNDVz4wRyHd
J8/8LCRtaSQpMIgw07djiTnLg8ZA+GpRaxtsEZUEF8pC6F0BIosYWlggBupANmqV
HG2KS/WH7MSmtlhtDNJSAGH+dZ1N5F3k9F2/nlzvIczN2utMpAVo1zfnszzb7gn7
LBrXzHC25dkJZaw8m/mqxdyYaKCwZz45ObZBP0Tjj/urm7MYLm/DhOQE2JsVPAz0
BoLQAEi7gwdcpQE76I+pBm+g99ezpVWVenUBUfzI43PxpwpfnZxWxkN+1qTK8HSv
WXweXYeyqkGR7MEQD7oWM0tThI1OKVpFAo+H0PKeky3OZNx2R+fTxw9PcLSvL8jj
BhL11/av5vR2b7qaz4sXWrwbd2x9ATEebmCzyHF+vfvkN4lprT9cE4AoSOMXNS9S
yU2TFs0CgEb4iiWB8T2PvtMqLAr0FNibQsm48yttWjbFpRm4QpAv2teMCbHLGrgw
p71F8xq+wTxkay1kMHeWcXEY6Yrk6UMgZtdflq+3TVPTGhcWOI083eVsXA8gU/ne
aixck6DjIjGjHJNY74/7YtX0csCvYwIaK4oUFbjLcPSlPlN8SJyyby9gOFCS4QWX
UO1r4DcLdOWow9kvDLYlImRV4BH26t22SFXYeSNBh4BEWuO8DfDsXgAnisFKCf5+
QOAZRPsqzlW9Cu0P24Ah6gdZg/+cBCHb63ZaVcIhH2uPxI5dLtKUewyyYAoaNIZ8
8uNz27tJ0knGgVkGDX4GCQZWieUn6xWcKgJdFJGED0e4pNsMtq2uJ5VBYSXjoHjA
PuUKAbED7DTP9qglEYjBhuWnAMjOpXJFO7Hf1Ji2YvxhUgfdmqLUpBnYITJBsOmn
vX37ojL2LZ5N+ijRM3wRMvp32ukRWXZMU6jyvnwzIHCrBERG+uRT40DQsTcTE7aE
Pj/gKlKZUrwwWIQ9ufs0IMd9vyTutSmsNEhvPtYHzI+jlvCPKO/miuWZOLSZCS+j
atUafK60nfyDXwJ5W1qi5G44AUaYWFh4eh3cl0/idCkatWAMoAfCLbHZoa/jNGFw
R7guJ+YD+73GAXtaHZ+Aa2JCsC3uweabJlWBy9i2WVpeM5DwI590jgqOeBY/piEB
Y/3dsjbbybVkcy0zqGk5S3Ub5Jr5EztDSlrfi3Kg16z1nnf6l5eEBdllfmACqTQL
SILuxlMQ7bk7J+12t9xv3LctwGQbCEhYhmEV6E9R4HQ/jw1ZCrtrGZnSCkgytOE2
UbtLU9VUUH8UL2EisvPMdHiDgG4B5u9jGc/IoHril9AWHE2QSMT7Wju0iEsFXzpk
IR5mcRtQSBx+/xRhc8lW3hE17MysMOUOFix43z0JBUuL4Ir39C7hcO0U28xVYQF8
m11ccpwI0Je82eWe54Oao6kM2upHGST7YmBofg9tYv4fcS8w51pZIViw6vuVbzMk
4PQWgvJ5VYrF+DeYujFSxGw3OQ9Jv6JR5XvgQGm+cQO94pYvY2a5ejuCYC1YGHLx
oKxiytXn8wCFc8qYw4C9WRfmdrZwoPMuAast+es5YWndH9RHeolb7ukJRUansvxA
XBzzhyMNB5nGpiB5D0F50+BnDyu/nVrFkxL6IYueyLPwD1sLXMxs103u8uoa8Sez
0paM4ap6WeS3sWgL8buDCsnIhoHl5VRQZWvi+Hm1sOWVbQ47FWWsbkRvM1xppseU
trEZBEE64+GGIjh860+C3CZg53BzQoUgUo7lEqCVk/L2Mr+vGh4Bl4snZy7dM0ki
83NkvKKalAJ+K9C+hzDiGps4ICMhVzjlr1dZzPPqeR7mQVRkwIhS/pld+qlPd2Ic
VvwhcyKRDYlr78VhELdXrZtuSVxsSu0fQ/EwHltSlQa2s8CSQT+RBdMOeC44RAAJ
/cP40lybe6yiiLoxHjpkQ+G6uuGd7jnulxU7T/8QVtf/N1jb+v3ovIwtOz6kXblf
iThfuRBoHoz2ziJXB9vkdoqKJ+kV/8azvRQzV385Uep5fYrLi3lm9+PB7Xxx5ukK
ekNgmX+ncCI4ZlBxhREN29QRGt+KEf+txLY7ge8hEjTv6x8+xKKpQDhOQQYqOgmJ
9uGJyRBMjmi2+xkHlkHO/qumVT/oEksC8FwZ6Pffu4P3fP7P9xrudL3l+bbCnvAy
nYabMTB8kVTiJGpMFyBcpKKX6JQeRlZiHSWmUNJUe8Y=
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
moWCy2qxXw3msHbMBVz75W9x+c6NWo7x8yisoiEXweIiTv0UJTsPlsYoT6OZ4pq3
2rqN4evRw2nC1G2/YZ69fEYSIcIq9N4yNY+MtuNkeT2GrQ2i8JEmBubn5OHKGQ9c
3BaWfgCPpY0e96Wxtwi1IQxnOmZQc68TgE9JDEJ04OmWvgop/XsqKglYe/l46RHT
16YdCHE71S+mYamdL0gOXq6eJiEd0XI+kTFS+snEyhHNtrsJO52hVzJ8MfZQjBVO
n/vGu+FWCFfjDaxsOOVJB2NquSj90MvFGOcHT7yTa439YutSjBobMWfIKqAcFPEh
r4z/ThVs71WE1Myh/7fgaw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5104 )
`pragma protect data_block
MkPzwtSdGpU5RMsTyDb2En/AFMMp5VJeT7H5EMFodfbUEfH0q+AU9fdvXevNJHYn
u+kDq0eBEuJn26gpT0YTwmlu7nstjCn25PmAkilpymEr5FCYEu2izXwlgYhpdyKx
gZ66vmD24imMl3r9wNZmfz0pTMc2OjuwjpLpP6913/llVxDOBA8cJrKS2JhfVFCk
uhacEloiQiM7HKwxaFXsbIkn1OD/ryF6GND9qhCWyO4PKnlkbPbuFZ0W9Pu1AOrX
DwQSbBYZGCt177gyC1xdOf5WWvScyDBlIgZmebFTPXMv9sWKJTO60IBl5eT6wmaD
6SSvm/ajPIQySwmGcOrCHKxk4zfU42p0YfhEOPqy4Te5KoWDe7rtY1iV3h679UZi
TA/G60Aed9OG0ulIF85kDnwtcqw5gv8ZiKO9V0r4S6a5418FfD3hX5J4qPNXXUyy
CuQX1MpEKatxGbDgjcgX2lThABXtr20FrGenIC6QStNrk/xus+Xy7ecP3d9JgtF6
4ZS+6QQYN/USKP1y2feBqtxMdd/fIQcl4oNQ3cv3s4VIadukSFwZS4wL1YKOgwhE
uSxlowciNThYjqAmSa/aBqNR7OPzqve33aUElJVzOTiwJayBz/PsSW4lj5icYagf
mc4PRLacqbGRHvnllgYMahjamvJ6goGYQFVf7vqXT4Yp95uNwDJXu6w+SnxlgqLk
TRTMh1dnAAkzz6JTlS5cYVp6r/rVD5y8uCS8AKrdiItmoWSXL9J+5Rqaz2VOteTs
Wu6nBbSrO6Y9jD7cmGnYX0sYLf0Ca7aYAcasRurN3sM+y4qccPZglQeGqlc6vyrP
5/Afhzg3QJ0QichORv7JtL+ydNNmgY1uOppFRl5qXo+MEwOMIkrNlrXJkz+NxEfR
K3MdnF3cabEzeNsmExRx5Uhb4EtysmLmQ0Ha2q1Gq9Kt9b+lSmFVNUfUhbeap2AS
DjA+VdcWQG2LYfGVRGxNQW6W274yPgzVcIuSAJyJG1BRqxucoqbsk0prd0QpaYos
DQoExRGq7w0l7jVYGXrVVuaF5hz9TpYRgQ3yYpeea95IUk9tSVQX4fAu2Cec4eVu
T8F9hFPgrPHJsGUu3VSNy0Gds9kftafaYp0sDfPFNPOGYraZ18Xnnd41CA4QwgK7
h7lr1KI07Dt/W5L9d+Zm46Vujcujtm/XXiRc6xCCTj+7BS/cItj2cjsacOHa7LmL
72XKUXPS/r/ohlTgBbV9KH8dNHUOhLgKPw0hPV5OiTaNlazGL2zpba0yvdzwuD6N
U3mGXDyDXTrSkex3YD062fcFJTuavnx557ogCJbDjVdIqv27+vUAy0vNZAbsonmB
LkUDKvUiu4w25RZzN9B/mAI623jMYwOJv/at09wIB9WWRy+SEj6hKh9vMcYYu99q
FRqXnLZ0kwWxAJ+o+3KtxaochVP6i8X1W2KrrGTz6dfB34RUK4LZpFbolz+0TXDL
3JXoNVVTTqzD01EaYBgcp3T/w8qTBVGOiihzyleCFSASDMYWcTaUO8mlN42Q+VKK
3Ysp8zupt3ga6t7J3lT2zf8sqGc/gKCQ2xeEP6DfOG9GX7ban6OFWykBuTApwgT6
FU5FBwPQAAzCPnmgIwvHfH8XsT+Lhaq/9LCLLf86Runi3qvBNERRLjhkRR0aLiPq
vwiL0rNvtGim5s7c+/HHgRyYW/pQvC1FUNtjXJiiaNjIkFUJuVd0RXtZR2SCAt4v
/jW6cEKO3ikXbWUokY0BcmgU/njuEHx6z67vtlJbUfyqnWiepLzvao7P3gDErn41
Uh+ARsaXRTZZBq2ikFHcv/oAANVt3MUmJCNCytA8qfmY+lPeQGD1fxWsbodWeA6O
TIzmd51S90owvG9Z0sYPQLyJHfFf2dwU0pnm0HGHhX8He8HDSQ4T0TsQ3i+2p0am
fNYUQ1k1vbuc1KV+KeZT4uYz8MfJT11QPkmHIcfwyZnWF/UVUlKTfDPLqAhMjFIJ
ToC/M0i6cn8PORMZK+Fgx0hud15Cc+agu7FXeMO3RPA8TtIHNT5l/mVOVpJpiUkd
zQI8F3Rau/UkeFuZ+T8U40E293WatahWptQ5GUIjoAN/bGaNpyOM/nDrzbgx09pE
ZzMseyX765c/GrCwEsxTiOXfRZuq0VtTNL4u8YQVlkaQoV6r9VIsYkRw2U+j92pq
lJETPvvIrGUangS11QiUlxyUiqsqOXH6SE7LQVeU4zHni80a8W1bXdMic8triRBD
HGDSjjgQloEEgz4bUC/e0r1yA92cCKe9DFmtgL/dY/CR3GQx1Kgv0sXS33awG5gb
afi7NAlKV9ozk3ETAbzRWZyZy5ecU+O3GXSgYgwtCwgnS3fuIwjhw00I7BX0698L
YM9QX23ez6P6BdeX5uu+/tUtZaaKxq6ThqlZ6QKBP9WlI9c53dFCosOMyBjGXUWz
TU5Yo9hoXVwuJaZvaOnlYhP3cClQ3NOxdpwfkQhpNIdWis+ewpwQE6+3kObxKpcT
gkmR+iduvMGcgvKYuoFlKaiVS3gpmz7winuYjfDJ5eSHCs1UQtKS6GrkJ3vrDiCu
rBBjv/PHy56iEimzZUVXojsL6JvIBEPF0LsocCFoogyl0b8sCIoHpq/bzYZrNfTC
c5ep0Rr5ZIPEPrBn+Le236ZI8OvbflIES3MpvOTwsyobPmP5SdgOl2wULzZTSJeR
zPqdlMp57EiOI34lhregdJ6ILzkY5+x5OTq+tne6LsNE68JPgERrVN2INST2Zslc
0RzdNOI3501c6RvnKNVLSei1IXLJjmWtEmIo5DC+xvi4C1rSt5n0MgFv8xGkx2KY
4/s3ElhRaymIWV8R7kL1q24f64SSx54MJkH2ncFULU12cfnih2eSigB0vdMfooeq
9UUJGanvFzJWdIjlSuhXnjjG8oFECOIbglubfHVnuWh0qzAvmlHMHA/NclGDZHKI
R7ZfyqP71P1Y2d9i5WsQ7JyYMxzUU/HMlHZ/7AOJbsLByKYs+DjZbxE9qARWUNEl
7Y0X6IgDXVs6bRG+6tacjnEyzfbEHBBYG7mVF68B8lkcto+M/lxJRLNONac9YXH3
fJ57BNQVEjT02+Ejew/nxDzKFeVSzJTE2yRpZBkSzRMCXtYWXwC/FsD3GQ6y8Vfd
+eiMUwzUrO5qJ6ySxLwLrW74IfbJke9Mv3liCi5JbWyMjqKg1RaFkiczSDAWHobO
EGQb0rSr+w/wqWKZGPbB9QsJ1rDtXM3QcmEf/0LzWYJc6A3qbHOoxsfLJZIyYZ4j
1GY1toPjKKWeE8bZmtz93E6062AFd8MA8vcWWvoo/L04C3NXCXaUwv+sUXzJHBNg
v26q0BK4NptiWmxldYCYBtPqDzF0jdqZ1hFA/fxPikuYKjlQVFp2cCoJeBLSXYxE
fY2zRFBqJtAFohxDoTcjV7GDRhZ5/47Y+Pb3YSqqmNhSEqIGtZq4Zzx4bIgxGhf+
heN05l9+QDmgPsOoqRWsHqVVqk3r/4ShUxSPYD8zHrtVADJ9ydReLhycEbN/ML/a
Jc31HTYF1+o3QVuGgE/3ufC9mNxvnAT089SJu2a7cCMDDymr95aVxlX4bEJ8ZFsF
AqMlrV83Jx35xarKxnj191fcLiG52GC9wJi8E34ftGL5DbkYUVnYEEsiu0Ls6BAg
KFNZHoniEEZ+0E4PEWm5FCQW19bchlZjypdkbq8quCd82pNvLb6uL7oG/dUZ/Ea8
CYW9QFPA51Igu65fRsKjWZlu+zfLCkuAXUMObpxkMu02wW7bbxO0iC3lAPr3+ClT
LEf//BhpVSSHPSIA7CjHHyXSMkPL2OUoiNU2KCQs624lrJpTwgTNkilX6YX9Mdca
YDONpDygw/LF6MCKON66E8vkHw+QRJ/WERVpK0NM2UoNBXEsQyrgxYKs3Jp5W/s5
WN0+WH+AIpzNgfld17o1NKgMVG0ODvLGKAKx4mUk+pasvOzQTkz68oJv0IFNBXee
t8t7YLHeL1pbamM45OyD7q8VJfpx75CTiF99xV/euC+sKN34TNzWGxU+7dsoWvMC
JIpTMoTbSaA/f2QdIjgeglfzhx22e2I7UrCgFiIxhMv7F63McoJpgbigfy9a1xsn
sQxV0pxqJpcxjT1NIjqYb45bASJ1UMsmEYsCeEg2Dz/UNDI8V8PqA4ZV63YYVovE
QMCDwaWjz8Ls+GCctdP8iQ6dNjS6WuzQsqZdyUqo7VLlSSrcH3NkXgcrvn1hXEvG
XRrWBAcABV6xeydf1szhRewN6xJO4VZCxUuBXHf7tfqOAhw6TPQATjOQxIfHdnlh
lFQSJLlBC5upFUnAgEZfvneoRPazDxpOECLU7JMhiIhFoJJVQNjXAZTzC5l5xrtA
jrRU5XtRsruvfZAAmgNJctnNWKObcTtlXQKZI4tRMsgyUOEofeYm/NIgI6UJndgs
92yBiCC+c1ojANlq7drPL0Oh5q2/8e7VqRfJNLML8XzjhXZr/CVJXUqc8UzJlW7h
sDHbVjtEIW51ocPZp/Tct9Bq4T1IpvF5hl9hf3KM4xeiydzs8SkFf9UfXP52kQJx
ypCLTCksWh44McEaRwAWmvrulgOBCyciJ0rVep/eH0J/muk5WJwObkkIB4Zhu/au
I/2q+K93Qj/mIxDEXn8mpu6kBFU6/XwQDHCJf3LxqK53UNpgjvrliEUqSQ6oovPa
c2xKhD7MYnIIniwrtROppi55xR+BhbqZY+hdZpFrHak4PnGw8F5TOVzCQW4OH3JV
3TT5z4nKqbQKaOXkVOi+u9M/rjzUsseh22vVN6ydQ4na31eaHqnBwsE79qT39vZu
GLWUO1ASMXXH4VeuArJNeFQcVqCWbfNGQZrBdmleZmEOLVEnZ2heF+MpmOZB+iA3
7K6y/zWTzGmB6pxpC14ggP4gcVtp2zpyZBad3JDE3xM92YHmd4Tu4CWXk1dAEe3W
741VgkmsvyyKxFUsPp9lx6Xz1zu7aPKPPnNTRLTQh/mgeEFuvxQl2voWO8assnnM
4cvvOrUKKk9YzLtW4wj5Qb2HLb2czfGvdaFP2ZduvUR3JZukHbl4gE8blS9fbmau
2b1/PvQI07KQ0XeOy1tpx845vMkHMv0n7IBg+mm7VMOf4f9v2ZFmswy5vY6GZqpk
Gv1XUyIUyWLcaG8WfhL/bngNcp7eXKRyq5y42k5OwMXXkRWWRu3Frjr2ZT6QUugu
0EPFRqbzXTlx7+WJtIbsWIJSwgT97h1ioqSUnozWzoY/SZB4DkuZl9u/OY8nZN5t
WWZa0u2A5SHqHBlV0yPohmjvApd4LX6hBH1eQ0KjwfgBeZkma96tPQf98flysA5y
b2aREiO2TGdVTU23+LFmP2yig7vln5FSLfD/xSfliY+yfxhfgka8S53DSwjb0URS
MwnKpLWh3z4XhgYZyN8ZEuSVdYk9UDr/0ZvgaUrNA9Qm/bP+NJkXvfnAEzSzDVj3
26bDVY67OAsO2bn8s5sqeN8Cs6i/1mKUOzk8obdUh9hZgfVdmSbyoh1Lkf4c+ScA
75bYeylseu9TohMb4aGnGbSmjVAy9TL8zP+jIHeYM3S/pIBJoQND1ZQhnV3XsFKG
GtCTIL36C5ooXAgXLdaxf4TrArmBiV+rkUB3MrYFPhU2XWGCJlluGgEF2k7WvIky
szJxgzeqXj7E5Bsyfoi5Nvnt5JJnKFgYEgnuE+o/jznvrkECzsd9xGY+08OlDUpN
8lrV6aUN1yO3qaFs/EfmYpxDT+Z9menWTCrvF8DL0A97+MzSlUWyYXYeGb1sAN0A
BhLdjFiDscF9FzM/7scJu+i8vQi9wFIeAvXdt9FpdDsQqPSgq6bURI/qf9jy72JT
R77+boF1GBzUe2/oBue25SG3rgmWcmWwnIJ83V9XR33bsAx6LNgwlpyKjkr7gN5W
OcaR7bhf6JF7xtfN0fDn/xnOEtt/VmrUFMAJ+6b7nKdfZ5/kjOtnosrggkiLU4go
YNHk1P4XYX8QDxP9mF9vpUEjpYflXNkwuZnfAw4Npqnh10iIXOXMiIE9UeM0/qgt
tEySIer2vW8E+NCui5Lm87KND2gaf6agAyIG208V+sj3gl86AxtPFsovjtL41KFS
YKZZhpwxVnpYh1gMEh9DKfz9vGpfghDXRKBwmiogdOXFN2TXdqc+ADyBipYzvTrB
T92Jm2xtrtrM0zgkSJ/wJwmxbLRiwWeh23ut72ntKj4VzmODBrqOW6r6uYSL7KbH
xvyG13G3yrfLmygUf871+sK8sZiYlkUVYJQrue65Ji6ixHxk7dNmmJDu0EmVylqD
bfsX77MXZu5fRH15bgN103fcEcTUePMJBAaPWjAR6kIxGdvDKZgf/JE6pbzxJnkt
RB8LNQaCnbYPBmKL8HitipbM8VKn3oVrytucJMD1Ivp1GZjskCYfFyXU+UKRAE3O
XX7BVsH8WYt2ek+2jXjlRTerTt6aUYlSpIOL3dZE8MNyYbbxdc/WSWtU3HImJHmb
cMOfQ65YYyo3Wtte/gHYOK8ZnOYVE80NdgmCGHFh1Db/2yKkn4j1EoDCtMsoVDWu
RvbUIvBlf3egF2vQitA5BAgkIOqPb9YjUJWBjD6xpWdKDRgI5Vp+PYKRgqn75kiH
3fhzmF1BLn/ofkEl1KIfaPUIAxZDWhpf9ZuDvdF+1dKcF0onyEG7877rwCtITAKG
CGNLPc9pubwsjEPzG5co9TuzHetuTkQF30VgMRcnbT1bJgg2F8r1VRLL7R1ShfB7
52vo//18Yh1ipicsyICwLeYgreQg6FoIUcnyVavtOYc7TdYr6uCQln29Y+QPOWmm
iLA5xjsAhguXkWGalpL7PQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RlM5H3zA4i7y7BsmLxwa89zXsI+Aym19nRg+Cs+iLf2F2Y6Af2epJT6IkR2HhbbZ
Vr3pSkcg3BJVhHscjcMywOi5sGF487HeNGrBtMZF439BqgmmQQe0OQiE9/Mc+eiu
AT6JGkFjZKjd/t9ExPThU9lekWODLT6/sQUvuQpbjy4c+Ja5boBLNei+HRYhG3Wc
79DGwJyj7iHC/8uuu13HfSVKSxdy6VOs9V8OXkHu8RqieOx6vozSeiWHqQwrD+iH
LXaUuuiWQBh4+07zBF5wHaLa8jOk9MjZ3CEAiEqWaAn9Vk6rGk1I8ByzAxUvqBL1
jGE7v4HyNKNX686kZU3DWA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2624 )
`pragma protect data_block
lF8Fkq7GIYwJpLHrp4/u3Af/jHrCYJ6L78DyO2EvRc0Oqmmca+RRQ2V3yR0/EJ6S
aHmnPQA1AZ7Xf7Z68UWdg6CQdagzfeJKrWOvpapE3S6x9ANL4lRSmZM5nIUdoyBa
1di7BsXO4I1KLS0ly9mlhOyxRTUKbBmAacW6+uHyJFSBta+a2jcApRSE70SMy0F6
5vVM5xr25jchgjQxQhO4k8dv/CqgrwndeZWG0v5ol8uGg/JaC2BAEqLg6+zFIICr
1yFZHilk+sN4XIBwrbPKQsUmW68VQ/kMAztA/K/Ducxw0IkxFM8LenrgLc8qGMYe
+/W0VKbNwcjO9YJJB1BgYrXeh5bvV9HEOrq6PWo5xAcIaMsOQjGdfyuF1TLURjSp
VwKJTBUGTzQjTZkjhgZGybrZoAhN8i4ZW/jChuZTx/LhC32BaBidPMdlMa5b4qzt
oOsjx0IUxCDn2Tc9RFwkg+0bapjwzIDHud/9S3mVRLfmWuLm/LBCWu/Hm3NKjWWT
mGd4MstA00hyblSyiqE5VHdHRiRqynHiHWmdodvKXs/rLohLKBhjH/ebvwKcehbW
1oflvYfVLGQN/FnGvAndHU5tF72XzFa95m/4n0MhI5tz/9296S4GkuWf35k52Wxr
DkO+/zrcnWPMkMuSjxQeW1vv9IZghwT2+sj9vG4ou9wo49t0qHAwH7enPJyAKOZB
LQSxMRCh17Ak6z5dkdGxrtH23xMxVqXUEOsets8d7m92RWEBeXhXqr+RoKz6f64Y
zdHsTTc+FAuwseChBkDFYCEFZBfsLppTJ2roEm6YIWgn6vwi56q8jycQhxoEGXAM
ASouenUrcKkZ7TOevlsqlfxSe3qoPOOdTukCJ4s5sM2fjYMPUlCaPnjeX2zq9kmq
vWF/SggRECvOl2EAz8XC6sOg1TOaLFQ6iLGYlJMGFwpcljxJCpklyBtQq9ptQjFm
lZecKYhXNonrBmFLrTHdhh8n+T5IKObdhZufKHTEiC7UnNlt3P4eWhBGlyZGqbRG
jZDDT1fovWuv1/oOuJhUt2hrV6j0CkbYl/mVwvnWVgUHW9raJCSmbDaLpvS7kocd
SZNQRRSqPSVJtc3PgpnPP/A6HCY0Lx61/5D5GMe2FM3k6QCfwYJQcvl3/6blqezx
C11SiWOwVJY16QvismSxeyC76LM8rIXlyEXLlcXFvJIh6ZwULqjv6NXLG9LkQXhp
K/1UwHQWiZYbGx0YI31o14QCze2NFlJHkBTDMZuTvslE0BW5/uirrof2TpgCP06B
4KEgB9AWEW7ZNXGSSaRbimBLNp1gBwsaT1VHRXEQPamJgqcudrQYq+7VMFeFylhe
dPpE29dbq6syu+O2B8O0R1boEM2mz/+iniD/1KnP6jggO7V/i0lG+zzfvK1JUCXP
z319mt8rHOrSWASxw5HejOJCbarg9tihOWY+Wrm+u8vJwjhlfZj9TeGnZkmPXC/p
jWDgEj99WQ9b+/vp+Lmkj5E3+3ldrDT7Nn0A7kAy1RukYKJhilo+EPJmnTYrW069
LRdb8nEiJDDdaGiKQgNrMIABnHSvolhBY0JOpkTZztNg1IRdkinbh7eCh+Pqc6sa
oHA04OVXFnlprdydEE0mjWq9qLhScS3hkIj7OthhgLhepbnlWp/E2COctrBuYa9e
xI3MElycnMVNaNOP+mtRmVUuM6zpi4x1siWFvC8iLzNqXg+aeNQxQlt8q7E5wwus
OkoEg+FknSFIB0DChdKPeX/0oY3XFC3HbxJa5Pfv2fKGF6/vURfaItAsxPyAV9Kh
Heji44O/qstNg7SGJYggsXd9nq/c+/Q2X0s5F1kAr/74cHseoBAQYV27D8JkbX5C
cPz5OQ6iVFQMuHONYUfmPHeFspFUbzdD8S663Pdq3K3awolOT3ohYv1rBx5HI3/v
vVNXSbNtKCoDgWzL0dtfvLeTdNkWrlpzfBdpKcw6BfALH9ix/Rjmj95b5/OnVJiS
01gSwhszHo0pYpaEzhUV2hrVWRsA/pmBEMoAZBTzQ/SUVDmuIu9QzC1v7Tbr8Lyh
FBnYwLj3aYvuC57PwAKHnyk14y12xTWzRtbqQkMC/V8zJujgtMyynO65PWNafSsq
Nc1vTGCyq521Y/fX3tSi8SHQnjWmv7ShdxuJheXqb05rkv0uGakvs6w1MsjJnzeT
HyfieqNqVl6u1YKNd7+LW5RJ0phfQTAMl8FNGTXrucEzxjtQajHJDA1GesaeojD7
Kf8XKDR3LZdCHH/c5hAWvVgYD6SJhKHh4Cyu0omIUp+MyJcLDjVk+uBdvptpxXPP
4UjoQEkpk9LLSMRqOxhZomXlkrj+lP1msG0ZG1PqzxRBmkZACwGsh86ydS/e/4Lc
ehoSMLxbiDMQwfjfbfwCaQj+Mt23jF++2Qi9qmC1p6fX6cnGEKBodUimcOBa06rj
ALCyuibYqss2J5AgAcmcrmJ/wcIE637B9IcIVR/EfliXeHoaOQk5x0L7NkIttV7C
6KcxrS1euyNFxhbFoIgMezlNijS0mXlGsO/z0qOCaNj5fow+lRWJMmdVRBxPHa3l
jvUq7Gh2/OWn4QgYNrSEvhgDzsw18+HZbFE8TnQxvEMvbWq6Ca23l8RcbWbkP63+
neyKB98Douv9N+0BTAfPSBy90suQ6u83zWLRmpvXLM08osAuCH7gqKmMQBNXERjg
OXdaquEVxF6IVL5u/xsF4Lg0cQqoJTvuBF2ZkMw0ApmCKfAFGh0DkYoWJgGa8QEi
NhXrxVz/SjG4LuAd/1ya6rGeZrb/h4rQ49CNCu7zfutWQvsJV6YFIPh2zr8rosgD
fs1r39exbiFVoBBFtDUvPFbis7p//wAdreYs3EcxWtXW5+tqQ0yiaPWeDYfmUrCS
F4gQZFH3s8dSK253YFDRRuGABPI4zFPqR8MbF8sHTHwGxq4e6J38AUnlv0vlTUm4
Rlgj0WLRHZ66xBoNfz1LLns+ZGmTpti1cpooJ3ZaJKdqGJvhW7LScwG9MMIn1OUl
fNiQfRpZsanc1hr6qRMpPEEEmhueqeVhmxj+mLh67e7pUxUna4yQj97Bxr79ofvo
HeR50lopjqJ4wPx6TEZ00tVhFDjtTwjPSlfWGu5moPDgRT8qxAn75mR6zj2ZnB2x
MCaPrxrc63XrrE3S7Uv43pVwdti4MMtdiOkZlfcRoJ4NnnM+MPLelwSQFfCpexzM
gVZl2q2nb1Th0BTRrfVgMIeZa2SufcE41rJqLZ3RWwAyNqgSR5i78Bhs9+JsUTXO
UnCrmCnu+wgCIxB09wr1K5P1KJrKhwhiJbS/HPkuhj9veiG1b6WA9+IICudwFKau
Lr0+QuDgD7TYT3mWC9I22Sn8Y3XBHGrGaAOFsrsqeReOWnv4szpIdLzHlUaItyrW
8YWo2euxEs+bPqv37dexkVXxm/e2d935gPQ49rWd7PqXenJNEXpU3qQaXBLoE1lN
2adVNQaLZnXogzKT3mZxls89T/PX0BLIBqNUmN1Ty6g=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
m4HncsLmmGvzxd+Ugk0AnSaWwO1r0zxSJV93UyctNP/N/Zqww4a7nD7FebkJjRG1
sRQf3DFQ00ea4jd+fDMIllGh+0MFweWkbtGg8cKcCHxgxVD9HAtlBrsubeEwhGvU
q/y1KgsH1EX5X4H16AAyJdNQCHhHAsHmBVL97rzTniQnNlLJb59/KQm7NMD/NwaA
O/AUvKq8kkN5g+WTOJwGFbicBVcqGWxkxG6Hl3Ed4Z59UhFHknGhFTwa3Yp/vcTJ
J9TWt0Dor2FDbFdQYOgzjeaRlseQ15sKNixLLjoyjbJboLWpDjPQgPqAlDC1X2dG
jYZRuhYNjNcAV9uhzcXoBA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17824 )
`pragma protect data_block
uxjcFMcXyOBV3C3pDCjEOZCB18QkzX7QHxRYMMXXB3TbY9VV+Ovz5kdgkXah4uCi
H2CEBQuHUS58rDO5Ix5dzpB1tdCgpWQOU9W65hPdoZwAqoKsLH7JpCLz73xG+qIH
6rvvXVNU+BHltuqXNDaWCbGqufcld1JwaeKss1SndWxKlaQMCtdM5ZMtcIkgFB1h
yma364TmM37P3zWdDlnb1Cwb4LS9hEo2rmcfh5yuSYUvyHsbNEke0L1XbAIIsRpL
IMYZnlyXHTrlx8pwSiDMfjMuoiK0VDqw6b7MM9FZYviFecP3suN0ZvSz080xEZHb
qh1yXqY5pXFRCCflI82jg15TDWLTTL9RsjxLt0PT7PyPbtCeHGpyJluGsnw3NR5G
PTw4hEcEkKmE9aoBhRLZQCOuHaG4R+yHUcLDi0Gu1hJWKvKp0O57l2yyMAKvB7Hn
LcD5TCwMlydRSQHUSJCjl4Lie78M5LAPCjj8ueyDa0/U0X0amQff6f3nhFSofRyI
v1BZa7JyFbQcJcKdzD5fj9bTB61k5PvX2lp7w1ZrRuJxNODSfW4P2wU0ID1DxqGX
d8vh0PSYRfzqEWSGV0Be6cMn6TYi0g9Um2jAXRFy5/nqjI4D21ahxi1r1g8jM0Ut
mioaEwGfP+zYjkdufvx9kkAmlVdIxJ/G0l0MWG9fC87WJaSaqVJukGDbYWvzoXXD
JhpgaCa/C2NT9D/Fy96Yc2qIbEDBtEckWmMsDNyIHvYRZjPxGKFitch9m7YZmoUg
mOd6JGxG2Ou7zn6JWmfGp4rWix70fH3CredzcUoGG/KSqJkaans/W9LLQaPi+AHH
fnSLZVdg2P8HkhHOjmJIayqtPtn7PmzRPPfqwO/XbsW8C0YOH0pYbXqjbT+hAUeH
pp/+/pe+tuk5PswtR/SV/JVSBVytqnfYF/Ku/3MtG7KTk0wAFzIyIBJQSn7S95b5
qLS7/bIAL5Aoig2As5MP6sfATMB4vE7BzrcrgdMXgEkoyPOUVBtZukzVCUdvAxG3
1jqET05r8DJ3fjQSvknn137facTnyuCjAu2CMFIJvhc27Iy3xEnzl2DONMrvgyjV
BA5jQiKaTBS7VSmJiKb5mGlmbO+2rsDE2pc6zsmJBBnmUCmTs/mdMf7kOkLVB3O3
JtTE2qh1Y2EGYlnAqqv2deSiHpgNMHhqRh7tG1s1MsXs7dgcSnwayXCB/MynRYIh
rFjC0GD7pcgx1bsJevyLsTEAbeXfS1xKpBzoBP2ioqKr1Y7QZAjZEgyz8p+jWiY5
YLjZj0XlIQcxWnMjHxqsm+0QihkRcfkWfIlRnLoNJIvUIuPeC8jxjbawFJkIh5Bk
Vllde9E1lRgHgf+0KAcFrhnnm60uWj4Xdr5CW07pX3VIrAmdbhsk3sqez61Yubc8
AJA47flc3/mWUdALrxbaT+cWQdKms73I0GO24U0hV1By6A+J5jsps8oqy8FSZeAZ
26/R2wTPUxGqp2afKl3O6kfGG8hYWt8W6bxzrMWP4DPVewYdI/4QVQzQ1NpADyiZ
C9rhn5l7qQyntBNPAmTNkDDnLKDZI+M7vNsLuyygidRuBdWjb2Zsr6GGrvMdCBbE
XWtNUagsISqOO5PnkZy54j8EDlxpjlhBS8n53reWkmVr8JnkkartQ5eqVp6nMofT
oEloaDgM3Et0UvPEoied0Ix7E2iMk8KCWDHQdqxp/FUS3ctQo1mF97hLNp4OcrXs
eXp2aV5fUMp3WJUqT9Qrjwu0Ulm9r+QZUYX66uPRdQncInDbv7ulbJSE0Zc34vzu
GUH7odohe00kiycKiMDBPVqCa4GNq+pDQrBH4irLArIKzLb3jCJY9gTnUvWFbeS+
SodqwV6ozkpc+aEN9b/8kAKM4ywG5FHmiwYsU8ag/AW/slrL7cO148iyZKKxHX3X
nxJyHgmfjUUhs+PEDkE8M3KLuwmQNlOxs7vVCGiGp2gc/U4m+lBiGwuurD3AU4Na
fJmYnwPs8zM9E5kEcOqgjZNa+sWV43H5DuKOU+eUWGrs/sHbquvlqHGFxpinYnxT
a+9UMlyus0dQbSc3KZdq7HrWkrIfBdeI5DzuSqAyko7pDERwhLX9u4hnXzZO90md
qqlHrDrciPMqL0UTEs4EetdCAuI6sPzTjk5nYV8lz0eJKrG4A1c2gwrfyk76UNg4
F6llp1ry/GpR9Rvj3tOUgXABTKRcTQVVRGD6RibZs7ejv1g66n8LnR7+6VDDUza8
xOdNgNwqZfvGERfGAoXlCRhrkVKfLfofETc9ghokGLAe4IFrU7My1DgBVON2l7+f
xztTsk/ReJ8dVhVgh5ffs6x3Rip6urYAQ0zVXDL9A3URZAdN5mlC9xpZJV43pNhZ
v+pWebwRjG+ao6JunNz/1q2vel6jNkQMq2W9xZ/wmDPHYueTSdvHQ3e1AhzHMKIY
o5jnJY7YGHCeFPcV796acaHz0Ov6RV8VRPIQrdPx2BxpPRtpHxifQ5hKU6cb1CRm
slS9Gx4oeNVxmOMO2xffYCV2JFkx7rWKw40Y7KDu4DwN8TUGgpBptIHmji55HMkq
VrkQYU4eqTl7YNvvtKRa63Y9ThVubjFSk+h2gKr7AT6TwI/w4DL3UnqqU1GVgNUX
AuP+J6Ao6qcdoyPtUA7LD/WsVXWKu4gmACZ3DQa/2psOjQb5PpnPVwuVVbxwIpFa
2OE4bkLQYZ63dctT/Ln/tu0SvSuGFHm/E1ufMXo4PI9aMG32IWFXle1r5xYOhWhp
p/h1BYG0/gyUOQcas/6OkNhrw2TvDKsoUsNUM+Ltn7NiZa3gRf/V3X0DKDYdvQI1
CFUiOXNO0x/K/R962JisQYMBYlPQxburqey14t6/fv27jInODYmjNM7OYKdLYAoa
RHSJiw4rb+Iv5JbwvPyxpkf8FA5i9rJOlrZ64XQBKSh+SMXOf89q+6ZIN+EtHx/v
l/Shgjre9PZZ3RQLUIFOkmadGR3CM0hmTpW58wPiDhYYXUZ50WJxEXkMUktwAbaU
6Jfd5l1t+zUKVDMEAXYZftAbDnpxGgVryga0H00h8C9mYZYC0uAatmOLqWcpoetI
QaoBXbX61rJOlozbYZzkRIZrm3F3NJOQvYLPi/6W3/2PtPo/JgUx4vEtGBGx5KZJ
I44FXUR509FGOch2PCaYootFTdPnlMCm0uZ3HTwlogBvDV0QWpjetfeuI6o8bN4Q
w/tfxS8t4ngQeZ9fbsYcyFWpqykTUeABmwJZ2pLPNQZEm0cTGt85Z0zHB/h8aj/v
Emoljl5ZVHjba8i5zUqSakloAZHjVluKQEU5VEZIedYP19w3Gy1sTAJc1SM7iWmr
DHQazUu7qRYx69uEOpbUCEkYJXYK/xzspGFTyX37iyQznnm0ESxyjvRhhZicrajt
zNJEAXsIgrvzYHK+8BKPeZFk3H9uu0K8XcxoMhPCFxaQpLQQDt5ExeEfFrSO/MQZ
0CpnrYpUcrgZNujEvFcvtBI9KfTpyoUErrcZwbgXJUFomEkALQK6qp8dfp3oRNia
DVAPNsZfyQ6Xvfji3RRaW5bumda7Sv44wH2OxbFDflJKeC1LKKpUZpZ/IMqcJt/t
A64VDB1oZaEf1TrADFN11ukiE72vtsiWLWw94Azr9ceZ/n6rFFwagq6wpPdNZ+L8
uH67u3J9B0oBL/QLPCt6t79KTN6IRjqzwTDTK8GstEVq8SK1xTkMrI8qomgi0ZWy
I8xpYiidogFBEml3VsVmRtkJ9C29ak4uUzOR27+8lTBSsH9vqt5Yi3Lnz9/5Wnag
b7LmbQFinD3ChAB+Wp5RWnkPsrtuGv960+eechanI7rGlPgfcsiZzHTDoSGhF3gB
QNEW8gXecg2UT5Pcn5IOhhHOz+vEvEdQ/0KDzi63Ha9+POdbpBQwgi3UxJtXB5J0
eU57ycXagC8FU4YZIOyZrOtGHYIepy0hITxeJI4LXC+TJ0qJNKDi1DcYqUp3AUzq
zPu8GbQ5SHNGlBSt2W0GyHGFqI5Exdqgh9tXmu4zSavEOcSp0fUvDQZsTssWrjpz
jqIqLjMVxbM3RJq4itKUon3MGGa80MMHi9u7or1Znox2e/8w1oHDbv17WL9OABGM
kA8X8l8ZsDIePTSXuy5X7khXK8KUVaisW/Am2uZaah3wtqnEhXFFPlPjQmoAtx6a
yo+RqapNbhe41NcvSaecrDRcXmU8iVm4xnMdMzxQQrKUPoHEfZqNOIBI+tQNBrJO
j6qgR8rMkFZLJHcD7P5fAcx0ahG5pzngWtFhV514ittQ+s/TbU5Zbd0kw/dhdzsV
z6oaf37G3cnO9w+qa1TvrDfllCkNDK8zgve1QF8fi2bumpYXINnim0dDo02+GxLB
+oKSfxk9riHgvNUprjQs/BnJXrs+aJC7NADkvSVNm47unQ/rmV8fBNvSYrCrkDPU
+suexu0QNdJ0A7TwHHDCT31yZQ4FsLZIMOh+TaN8ZKoVfo0cosVI6a6px8dtoybj
zC6XBKrXhDglLCx8T+2SVj3L/aZYdce287Vxsc0rJLwgeIzlzv9XufmVxzkuX521
ZpqYJ8GhZtcKx4mOryf2pD77kewJ7ENUu5HOX/1xBtmMk0uzoNpeEZe+iLQT6uUM
qY0we9B+7+NMoViW2JjUNTSn8+VxWa2Aj6gRIP0tB9Z52RG6S9dkvjj6x9TurwCX
7BxgS3F6xCVVHugb2qalJsMXU/rLZbybfrvg2KAfPcQmQ25fp/OxWG/PQMcF0Jkd
xWD1EqH89ReTTYSGVF90I0iR53SyXcYtpOpB/VTWb0g6E/+Rw56RtoJnrYSPMDmO
wiN0sweGeISQZD52cI6Kd8qmaHC41Fh/Efg1wHJ2wlj7WOj9j4obN1iIfj9gZkqd
MPdBI8edgyXVPMWGJjAUYMix3yDwWZbjF59xULeG/6COFBvLpEpqJtLXuAkj6Pfl
W2VRcoGCBkEHHzQiBGxtQoGONAHpBp5Ya6R21Wsv+Ru0fQWRjH1Vug87lDn8x5Ug
LxE57dQdNWlub7P2atACKew8Ni4AI5cFT4zf5mMNp4OIDrgM+2oJDgRGDOVDC5Ez
1bQP0E/tN+lxZgU95w7DY96H0098NxIrYSjVqEVtbQSA/y5DFo0FI4m4UPRMPOFc
WYrPpvne5tqpJRTBf8NwbdoD79xek44zKBNIvc8dTgZSkb0bj6eWSQ9l5RybuINA
+ZYs4QYalLTUvMzA4WRi4tL4A9oXlNdWiICRHO/eAD/U11Wlldg6EinExq/N+RKq
GYNdRWutfD/TlGUtgXlt9HcAMd0CXXZBhU8jdwcZLlGQUhYS7AISVAU+aJLso1lc
53jEdtNXNgDC7c7fStaLIYxSJnUtU5dBRjjI7fZVO70w/Hdulm9LhqYEQNAovCxt
az7eLtmJG99X8qtqZjzIWEDZjMDA9VGn75yJ0Kqx5Zneov3CUjCPeS96vDNGgNDx
4ctSTOLtJ613wZJyO279jfIk8NNFV8o5S4vGAMusn5TClppbddPglj9Q0sjVDSEI
3r28DDQYhQyVklqLzncbMTWVF/QYy3odA7zhWA1S3VLBxKC3bWVsMJz7eWcwgM1G
ffaDJrf6Kw3UuSbAJD21et+XK47BOn0OvW0i0T9h8kVsLj0AalVW7bOwuY3fkIpH
Q6hhXd/EX4aNGKIoKnlLVpUTJvIWDSuxx+gJ1mM6NryhbCvAoQ4b75BdnXNCEFeX
OySWTHMMEBHMo081nK7xpTaXovm3rAC61Fxy7zCRK0LRPV56r7QnK17PtkBVILau
4CmGK0T8/YQRjEUkDyX4cFRArnuUS/CXUszAwqH9BRxzQ/9ftk2AC98xzmMXchIt
HkC1cutP6/cYd5r/jO5y5NwiM6jXHrbLpjNkFNau1kEMCipewpcBSC063/bUSgHI
Z5gjts1BUNEitwmX9mXmvgDL+Di9KgJqmTin5TS5Vb6odq5Ie47H7rh0bMPjEKNU
uPqlvQWw0q1IZnIT7Hwlis9VHO3+4URDnM/4LlvqlH3kjTVJgBM+VSfUhcCRk8lz
dRr4ANXZd2fupJsXlti0+vv0wXUouA84OAMBaU12q+7I6wPHuRAMRT9O0g5+IN5/
aDUusYRgUflX4HHzop7BS5SaDHLg5KdIYh9eA/FN1vMP5ECqLLWUiGwaWgFf3s/b
cb6Thz34LUfEJoB0nvbu61fbyVt3AU1C7ULyrjgRxInBeEgM/74Mbji8q5d4T/ec
f+FS/588vKCkMkJpMiMiR+wU7v/x2NC3HF47OijOtdxqn/3CqbjzGdCg5KuYGT2h
qYPt+I4xKUC27BEG79Rjhw8Y0ZetLrRenFX7M7Q/LxCfXeVixpIrpiVmtgOEsTvm
NZV548ghdUmozROmcwrGe3rnzauAqusMBsrA7zJJgRSCiv/9AP2R7wdClUasYaZ8
JOv2+/c2gRXSZvrBM/A+hct81O1Lzjoi06VAi4n9O+v9MMO5hEmHoDGB/TYLjuXE
/q3zocYEZudvNojR/39DSPvA/XhJEvv22dk2C1Rir1KS3CLRVVfUndU4XRRMFidb
vJy/3376it2MJ8ko1B2lhilyDcn8GP6GzDdZumtAVdHrTGW+SVfTLakH63YqjvtB
6rsvxaqTGPh1Uvgd4i049cnUJN+KoxTcEp2P31qMPZFenTp+QXgnIv8yhHEv0gTP
XB0RhnDstVcw3A/sZn31Pty0QWXy7J88fePdjL60nZ371iGEtUqggtblm01C94ly
IVkAwr0ebauCAmNAi8g29p3UTPqigJo+s13dBDt3u+7QWjySCTHoh6dhMR6TG1gq
BPEjv7mUmi9PTCxjPmxpAqWn2bfC1WVnBZKLjYbPriXYUROthC5v5yXbxR2Qd4cG
Vwvh26jY8PfIS1erjUiGkDaA8vgzn3aleEtUEO0XivyX09yHClZf/LYVHV5yvqo8
JjmN/G11H9LAEkc4kzsNiroAnBikZ4jAt9dCqeoIZbVbGpL/PNuAx59bFO7KilwA
o4DvgMbH0/rzmNakyZzzl9nFwfH1T+BFwG5oiFo/lVgMm+MZcd7kvLh6OsIDtOD1
MmZ8q1YA9FI+voAYGWhoC5eqv/ZFXsuCSHAPLxyptvGbaFWXBPiz+gQ7ZCBn5PkT
RJ866+v6i/BO6o8yYC9x28bFGoYFgrSCnuLjDGYrWjIuwF3BOhPDg5n85d9jorqr
NVX3EY0mt0iWKVnvf+N4P2bCvM7Q8Gy36MwJ7xH18aB/H52QLzN3SYACRZQs2OsK
hr0lMFidBgdxFpByO3F+cNv6eZnYk5VvN4+joeihkp2NDVvRedu7TXUh5WD6m8kr
PScDJjL6GwAxhexCy0BW2c+N2YgSO0nT2cidsPqednF5Fndfdg13O00D3MQYArBb
hP/mcGLHRohd2QSGc/HjDqF8HFyf3qH+venxNhpXqGEGKE/ESLMMBljGZcGUVOsB
/850jjUh9DR/6/v4XwJHE4bzFLCuf7OwP+YXADvpmMp7K9fQqSmT7/tgKXGEgQcJ
qEtn1KQUVtg4qBXj1/48djMlQFGRxEhQBo4WpZd2C3bZ1LTckj1rJyl42FVxQrMc
+tAkttpYLkWLQfMnetjx0y+/jWA40Tf5mymlYgRi4OM/Ibg44NaNc1+04p25bMl7
5wwLdFIgSH5Ai7xnUQHv+6bV1P9ZfS5wHHyIy8DAZS0iQaPy+L7I8H52WboaNwRF
jfoAxgr6fQhKk/R94fw/68gXXGFAAoU9W1vh/gULTx+UGllveouYE6djeG5uy46K
6k6SPYj+aVMa6RIIs8E9d3psASJUzxXlzsyGCH3ekUtpoLlLcI9o9LxwOnaQ9k6f
l6tZvhcFBGUJqzJnH6Af5UXcI+BTGd2Vmlb8rzWerDExdXstPd5x6H0/rAA5OvOR
G48dIudJkfX+VR5Uj6FMK6bIzjySt6srXm92ipC4wNUyDjB+X/H4bhA3OwNId1NS
hTFmfT2sLDN8TUwafo19Abz67rP99aIzqdnBncRBE2D1VPI5V4XSQZSx4+gXnAPP
AKT0520hF/XYKdKVt+cdxNfrYA5UGUUjd+IL6GG23jOxw1F0dZvz9xYTEtvxhT4S
DsjXVg54iS5TdPC5RYkGEqCI5l1y6h/tjhpHD8senh1cVoLy5l1Jb+vw9VoSxEp3
Ac8AED3FhOaUpZCEjmP7dikCnDY45lA/JsessUwxw8xp0oF97qxtaXYS+qHhvFYR
nmZdXzDbA7HU5r9mnfWBfnnWFhuTNDAxh+sg8l1/3qsZWLOFt251Dky70t58PJ27
1cpQ6JuJyFTWFE2WCNklWvZHuhcF9L0W0vLQp0s18F41HkC7xlu89fF/AJ/zMzw3
VcvBAmi9wdaTKLlQbrmWCnAlp/zck99fvxEOJs0DCbtKxqqlm4zJh9cI39dBCI8p
dtz3Jt61A2skI+nVe/fUUqnZ1/CGQty16D392YdYmS8fJGYVROFEswSnSn23EYDg
bSG74uz5xEjbSVza87dO+qQUsK55jGiEg6IiIi9yN7QPM0tHty8pZls+45/s1G1S
wDrqJW6fp5bS1Khd108+tVEt+6y/XgU6M0wC5ggs9qPXrYwzHvmFVdmr9TNzfWMA
mHq7V/O0LliZNieNiUBPzVpd5L0FrtvhsD2a6YTG021OP4srEDdXRpjcNcSM+zJ2
llyQUAawrEMnfFaRSialSX1uU+jO25fqEiuGKHr8qRrDJPfIlHV6+qylhoLpVS+2
N1WT73uy6KQZuaSS+crEkDJpLTg9W9siev2Hnv6d93hsvvvvAJ8oz6nIWZZ6YypA
UDu0KcPtjG7rylVNVNF9mEcp92mQ+B2bvIOI3g3uSffIFzPtQZaPMdwpKRvwptc2
/rKKLmeGoAjKle/95K8niIWp3RtzWW1O0WmGq5eBksvyjPJQdS1OJkiDDpXS3Oar
W/bFab2Y+CNpitqNChfwKhVEJyuqs4lcSCzMFxQoLXB0iFujqab8r/VuMwrSj3ip
b051r4yIOJjM3IQv5V/Co371sDp+mFwOZNoQ2dNIsz4ViadlQr2E7mYpo/lzNl/F
e8xMAC5rZsUsM9V7LOi8aFsTWNj/nKBdXtP4IIAI5UmftotiU976MwCa1k3VxmNr
ZBlV2GOwG9DcmJ2Xeg9nkv/8RmkAXiw0Hx0+Ns9GXTxgVNsPUp6K1IodtmKu60ca
tWCE0ID/o6/iDO+tsLb3v/0ImJK9FRQXZBJCt2QNzoG/tWUjqJ9WhzMNYPMIiRd7
t4zYovGng9uNSQ95fdyLIjgC3PeoD7AX7IzjSwyFdd4L2XX4ZTGemYXMNOKk99fT
BT8k5A9styv5QXKpSerb9CH9/+++gUVix/pTNvg7Xg/QpG2ncM1m1JfSJEsT0Tj/
yAd4+XjLPd87r7Lc7r8BkVIJ22vKLkLPvG6u3zEBDY4qQZLJfhiBV6mbxg1nyMKz
c1o8j6b747wTAVXy1RHI16/nxU2S4FG8WZqRnjcvhmEhpA5i6HkUJH+ytaYywtYg
nM+Kl+jlRUkoGnG6C6stl0+A59dS9WqJcKwny1Ss+xpZCwAXIE6bqPThOjG+KaYp
rJfBSVNVLWfsxAEWDZxAgKcI5udTh6QiOk5MFFRxtlcHGgLJTIi7nPw2owNraqw0
L/ssMv/nkskuOVkMlcA311HHn+tU6pwG5RswWp1TDltSNjjHn6EftCdARjBnBawb
EMQ5EzHtLbw4ktKbSnjAXCN2abJFifbw0Xw1TI0RD0HmZ3AvxIm/mj3iwFkrBM78
QoDIN5a/5NjCpJaNY6I8eWneJo9L9W4pXY0aGoSPe4f2UWV8KAbOXluXiaOz35sL
svSBKqNk3qiK1N+LRKwx3YOkFThL6Xx6b/QAWkNsUg8UZXj5xTCPK5dvC0wk7SxU
F7sU6QvAQTIsJFdIavFtH8QE8afqt3i00Kfi4RC8QaKA6IMmTtRWYe4QZKO1UoRY
Vl+pFZaZWQUJWEaSESjeYozWBYpO4qB7HG0haJe3vWwKbkwfA7qzGVdat5r2Jy/t
VE+H07wBEj/18qlp/41o/6mlmSOLbktiwvjHP9CsWQtcjgBDgVNIqUq+IO39jDl3
HZiJ7qV9TpAjjvUhaEh9RB+EDMwiaNYJqGDSgwn1rqYgcIIaMiFJx/ZTzPlrYjVj
6poNUSzTYNaKsbEpE0HgmDAiP0u+mQKjvvbH1gFBVC5AhOVWICdoyHKagliUa6+l
gVEjH89zHyhYhDx8gqGRWm4YQqVhEs6pkbe0cmyqdWCVe5pP54cZp+zFD4Yjb/t4
PskkjMwBc6PL/e5uSQcYWaWcsWaAKvySrgHCBOpGqICJIK0l9zGOaEL7TJyHKPsi
PV4FubYiDKYX0V2d/tfT4/rP2wlWIpEzTY8IYGXR16j56gWTs9p2Tk9qIlOrgFfr
PgELcenws2SCiFZXD+bKIw2QTu6Iy9Oawwi5vuuS+pd7ZRNgzoSHn9wQPfNTghmZ
Z6q9Y6PrmQG/iNq2tIw8i0snA9QqQVz7pTf3kXbbAtyMc2VZuwmWzc58QhnsGG69
Xu6yU/o2oAbAHcb1/q2mpcKuBPRdQ6xK6w5hGs7Qy6TIhW0STyBntgPg48Xve9qO
a25oW9fwwwJEnFKjiZuv6VzKJ4YXsOsCBOGnYqoy1BHW/m2JRbBk4623PJfvq0xS
ba5cWfXu9iEig7LVwA26ZUz5pSqI/wOb8w+SpAG+wLF4lIbJqDe0xEbs+PwaEOMD
Y3JfrI1U6+Iat5g4OEg9L5B8w2u51YkzuDP1A0BwXc5rzzNER9vjN2mRHZICobMx
L8AwzyI6MqXZPas2mC7qfYk0AHO1qoZzW9DQpoHJ3ij+kl2FT7j1PO02M7FAGFcB
+R+poBzGbdOt8j8eQN1U+hxPt5A3jDFcZShE1VCtM+8pwaB9S1cB1fZR+FDy52bl
KyNsTt9VE72wq7b6I3Au3fXVzOMF1qpR6Kg7ldf/K2A8C2KBiJnR8wDUUEhP4Fd3
hfyVmxFyyTqT8BV31K4vA78qBY4R/wvduA8+XS3IaEi6NcOvsD3R/kc+J4qKO2Yt
eanN93WYNh250EYQ1ptb47IeMlBnLWm/u/+++8bJhMv/5/7V/s4PC1XHCSqebEg9
kefXdNyyScPRtcv0obBUmXaTbHbGuIT9Vq3ugO2pQsdpSskkECwDf7BL2RY9t8as
CDXsQYG269gV4sylbz776xbQi5xnC+9b9tjPuA0N/oQWcHvolWNQ3w4G3cBFbk5p
yuR/P+elzLmqOmbS/j2xVk3on+yUcDy8VpZ+1LaTEvmoF/GzmnMiBo7W3zIuDw32
7gqY/cECBM0d2Vqkn098/WoTy7GCNCVgvOjWjSYfkphx8qnb9cW966hu3YpZQxYH
TKk6zofAsfnUbJFi5Cu/o3VjHm84zIl6jYJ9jNkIghbu+ng0TyZIU/k8v54XXGyd
BlMCuVCsCaw/PDbi5sfjoaIuKFVVXZ89Rd9awmksLhImRfOA9fQpSAqrLixIkzxv
P/ar43P9VT5iIbPrjMAdV6jDAfvTZ4GhaHzr+7HiKpZ9uAsdm+0/blEvcqDE5WZt
YXESj86K0na5sXkCylX3HYUAD0wJAP6kNRgRnn2Ddv6jb6Q5hqHz/4Zk/H+cbv/e
36Pod63re4Q0avfJDyGAfYBDfXTaVPqkMqOmFbwSykNWzVZqEOpC/6qzSrRUK6Xw
zB3+EO8fbgp1A62PSjxnwmSuKz0Apok6ebS34Mep9eaH52tkoYP1LrfeTSdxw74y
MVMIE4cVu3ut69tfMRYOPtC3vmf7B75dgFnobS3N8p2EQJbR1QI7lgyO2BbtsqOg
bSgNqmTF2LMgIugC4nW80FOjowZl8LtK7oYNVrXYr6VHWFTnI5zmXbGiUijnyJwe
PYhvfrchyfxKDEqmcLwIobanF3FCrpQ/vSUjjRSz9jWTFHhxHos3i/J07knCNBuc
5cPedNHCk1Wvna/r9oLZXxwjMrwMfbHKvaOB90HID7qQ4v0dOMJMZekMGKCfP0m/
YD0+0Gs/9Pk3l8k1ogpI5+9pwGdYyBb05A+njDWpTMxGcx7Y1eB0gYSiPWBUNVRe
tsJdCzRZ1wlOH4cYaXz5kBxVJhbOIeBhgJiaZ5zpr0LC5c2AkN77CSAjpBcyKDcQ
5eRwJBmBVIR5WSFPHjInhAQFTPxE35PrcYmWNbb+pWlEDyZTiQzvpcv+oOO5xwL7
JyezZnZCvwZot8gbgUlOqZ6P6dy8h2IV2wQShDCJubHK8MUKjLvOuCtBskPP+Vp1
dPtQD4qxxptBNR3qx06BNqV+5Yh4feLesCAmRzpLygkjMCTOQCG9DKdyy2JP7aY7
ecLLOuwEqaVNB6ZykStMXUQLt/L9crxPK8mkUyquQNKIV3d55iQl6XTrhNGg6AQj
+TUgsnPUnHsIO+VlL/P3gORL2oQWyDgStlGQ06rWMAhq6sgf/NHSVSBBO00lQg0i
1zyWn70+BoaxglTfiygqnBa8rCedWqncZhEDYchKUXY+jAudDAKrlBNIFv9oDixH
4x71cSj+4MG5Y1SuVVMrLPAqSlBtl/CfXArwdenX4bw+e/lEI4n7bx149tcUReaG
SMhvga8M+XOOYY5ISJnJBiqkftqFZo0TOzyodIC9R0fJfAmN7uWDYcFsLzkt/yMu
uoKnnf7nXmoGNY+ubzbX1nwfa997PofSwD8Wz+TAeWCZD8lmL7sqYvgRZDtiQuab
3ZjScx+MJEaAeX96V3/eWWRMt0LY4VMZvMg9LT9UTOQXz5rAG/6kC0SlDp2sRL5/
HoggDPYmpZXVnwLylxl9Ndm3JMBFXdAUJsjNvC7FMWP3ptGMrB7miZhFRo5tPlFJ
dzRSayEshEuS+1Tx8ERe/twZhI9ddMN/4jBw7g5LBqpVN3xhPYuI9qx72n11jhFb
ModNqKpSsCKNXsE9msFawrtmrxzezWwENWMEfz907yXvGJXSHA4kfBukiUARlnIv
bWgkL8T3J40WM0/sF7firBLJNJ50SAox1rrikOZEsXnevZ4VT/E3UKTq5rRIrQZa
k8FSRbhUn5vWZ6tKAvKg8V0OctNmeGfvpBqSXjohd/gNmz6kOxYZclJy9V3tqM/t
SsEhDf2BvzP0cODt5V4gVeel5R5+bl1/FuYLP2F/5yrSBzTK46kPJSaxQeEoTpzB
QmEv55NrUqL+mWgDMp8SWq9JMrqovgn2YPW2+4YfSMfWugRFbema/QDHC/PJgc7u
/5/dADnSliRINw67Ge9vFvlcAodt5GFhhJmGrb7ayiKZJH7k2S2QDwMRQ0jqU9GG
0cE2CPiE89kD2GuJhQxtdS3YUJjb0gRqb8y9PDH7mAacT7y5XdArHrfVYKmJYrwn
7wMh5P6ABahjTVShuG7ORc6Z9aZaMPK/6yqewIaRfhVXFYnjIAGRkjOep9tBQ2W7
EOoiRtS+T72r0ctfkAmlMtOXIt3L3H0OC4Tj+vtbSLNtwthQ0+Ts0hLwkcplIbxz
SGmc13wMqxKGwZ6N2O2F84fexye88jYfOSLvOt3cXAVERKakSgR0i5lUj5oO+q7N
O4uOQDU4+SEoSGb6UuO5nwezoZiSsj3siffftwf2UEyB0CiZj9844gWOtUTprTD9
C9dfG2SzmcuEi+7J0Rr5svNc68D7RZsYCnluGpbQd87icNjPHFhJZyNoG2nWiwWA
6dPC4QSNO/5nhYqyAFAqjCb+r+nmUEdVtGIaU1d7eOjAn5c3HAFJoJd4DSfDn3Dq
4rXbN40/Z7Y2Fo6pjv/HUCgxfWBhvwEk+N0lWYq6m/t8BTVGLcArTqUZg0DBD5nE
5Nm84u9vhqaTSBGq4gVc7990jdzZzN2Gj8YxA4jMOxjVbUXJRaD6FU41Wmd3VLI9
5RN4Oxt8Par8L3nggw9zAnhalp+AS/YNhcMYUczAnJI/TQsVeDOQtq/NQmmwfqny
eyipn/Jrxe4OLuTZsffvWKRNN99ETuJbZ7YYBzBrnmYq9FkVeOgeEyVfdmp0zpTH
AV2SPA/ZdyRlgXmSsXdeNZ/INtS9JwecsrFbQwcWlfG3toeUM4OgM530fnMTbtDS
l+8UmAO8z4oYsGG9l68jJDVMK8qBcWSYPcNF0wWbaS9Y1CTVPh/OSrcaeLKtcasW
mDG+2z2jqE5EiNHZ9Bgxl0j19EYDA/qBiM8g1oWa5b39KkuVw2ClEZf+Zn/bU74A
8ZYoOPDl4OoeA5ayG4nOFNufs2gUleXRH2+0COAYXcGf5Mv8iIpiVqlZIb2lhsG7
DDdTWju+XaHCDEmxxeUmZ2mbdMwYbrsD4om8ZOHRKHhK2dvBZL8EVWOD5Nxo/ZgZ
05qqjqcPycT9HfV+iE4O/rwMrTEHGIXphoyq1aNLQW0/pn9dahtB5nvmDP7uTGwH
s8kuxvctDoI88CpxbEiJ2rutmzJVOoT2ux458w5MW+ndvzo3sHz8ygtxcQ/0Omru
7JbYH8MpDBoEHPwTxWO6ZoU0U+mZ1AfbgDgErs/nZlKnzA5kB/UaL2W+0UYq910w
u4j8g/0R4MuUKplceGrtDRZ3Xun0tkFihKwTVT7MPuUAkokLTw+cfw2Veq90NYqz
Kd+1vSfazwPfrVp+vRzUMg1ow7c5QtKFpEiRjM4jXwwHcjiJGO0AtWhgNAuGztXB
st7osXOw+aGiFtAGDE7rAd6hzxAsKrC817QWucVVXkcJLPkCd7cJY0vAuJR51Shg
cDfk2NiP6xGplCJ7n2LGjM8cW7OhnfM/7SnpDZH2OyHVvsJA5lfOEUzT0+ZVzdgP
nT3dX9BOXZhZXbBAEpc1ZBomg8pE5VsGSXTHUPpT+hv7OKhAf6n9GlKi0QumIgup
xZtDcEcm5j61Mz5SoCBRaSVI9cM7VFXX7Y7mOMsBZ5a/onq5WZRJQoCqa3nqp0T3
vj35cU2l3Nk072gzftSVMefj8hWCtcujOFYpKQU4FX1O4ilBZKFmkxwdv0PItfib
vcH7rD+A7+LQzvI67oSX0Tzs6liMwBDkDUYj8Uy5JXDjEU/5bV82kIi3Fzs6d1xX
Xz344fT0kmf/E6SsA+mh3E7+f6RR0FlbQTaYjo3/yTGs4G+2ZmjhuZEubD7f6F17
DlMUXUpq9RoRpEWH2bbz32CFUl6krS9CLMGGhwe5N6WkFG0Nl3+i3HjZkwctLXa8
eyJxGl5xHGW0WGAqrIKZiM1pnHALmD2GxLTgp7XTdtNk70e/0I+T6BE/0T9z918V
XT/us0J7PQ3/bteQmCCRS4ECYQwUK+SFWTgZZgSAuDRBtuChtjNPgB1N6D1UqDfC
HkiL9xS5uj08KkpgBb8edY7fnH7j+4CXnjxSogIl/BCjqOl+lKSokhm3G4VRHkwg
jiskr5ulWNenkZJK1+9tGjxe9rERRceLak3EJm9gkh7Fdj58t6A6eKVmp8snUzk/
ql8Q5ckYKRkUE16KFq+RglgPqxMN1LsMSWK5Es7NffmhHQipg9g4CyksSMrbvzA0
BFLm2+4P+dltApt7QMKMsTpz6Q3oHbqDAgZPSEPxB1BTgQQwtM97GN/5c+Ee3CJd
PRJ7Y6Q2Mkglk41xO+Qqvb2XkeJJJR4yyPw59egGh5NUMXaEZjaRZGGxjikkhsMO
4WU8Avg3qqMUb9fPne43QQptk9bI5CsiTDprF0EUUnsAN7CcIvd///Melit0Y9i/
TjVq/NkY1zBTnVAzHvWSlQSk7JI/mzx6hdYQ6RwItnWohQRoAn+f72tASe6/DsYl
qYYPb5NFxdP5Oo+U5M9WDBR/mO49BxXEPlE+eop6JDDXk+d3f1+ofsEm2b6OvRIV
S5GaHnki1mJwjQyX2t8qofGz5R3E854r3IaK14UqyTao+FAKWkRvqHZGsmU6yDO/
NG07Gc31wCNwwf4knqJytePTn9LHsLBh+qFCfAI7zls4nYdEXNfXJe78I6I/6NSW
YJTkEE5Esv00d2Yzroi5oKjqFQz4Ace1dERkc6eij3QJGJUtNdjIpMd4PWm2HMTZ
LFEqGYKXNVvVeVtecIL4AquBwduepz4zFPINvDkMPs1nrz3IHcyhH7T0+0JHeFMy
dpb5ZL2OiGEj5xD//CN2K8wghiS5uK7UpYyYsEwfc4eR4esx6aLVZCge1E7OUdxm
4gm/F8v/R9jXkjJN0Jzn0hKRW9zTX1atxAJ9JUcVzBShxv7rUUYEWeG2YNrH7Io5
uS0BV62H5EK59wS1cB8F+6peTx970wR+qWDhut+k6Srar4zGKs1uyZcfFPfhNlUm
ruGo9l0hgjV9gffNrGAFSWuDbeQCq4hh3M0kb4BeYzVrg3xZQKCL/XC5JgXBS52P
smxvEiipQbxvVKQCn+aHz1hPImyxC8SvfRrOFCBIQT5XyZf/xuF9QVcOTWXp4LDc
evNRBJLAURFRlJ6DcsuJfWuxFIwgEBPtEUlJBKU0Tfx08QVhmllMn+9N8Eq/E+T0
ZoGd3kwQek9jTmKWqKPY1Cu76Na8My5Dhbk4TaLF5Yqid058U6I3TEua3h3XdR7X
xrG3p0cdArnG52rGRR/VL1rFeCvlqcBAY0A32xnfWC9CQ3cYOuTK7/mE0kiFTpKI
v2hyeY0c1JvNvSs1e2k5F38NOYHYL+gtOPg1lipRyeUDi64kw99rJpMRfuTUolDf
QumQ6vXLZeLArF4wP5FlsKpeF0nAy80s+IhVwUEkadzEYQbU80hXL5HKY/POyKsY
RjeKSIQ/fJkwZg3OeHAp1VIM8BtmsIhma1uIs8UOtG8T3pbDwcPNLcmWU/iRBhgQ
C3GLp4Tn/PggrcWyefyKwL8Bbom49vdlosoyK+OyosopyTeC0/TVRVw3BH1djkYM
IfwtxpWeuutXN9QggMuVBzUkF9i0vAQLNqx+LwmNb6gYuSfWIIx1/xA5Qbgmcjxv
p1g8Dn1gGKN4wMxnMLtWUXtDnSE+nOq98WOx8zc8BljNgbmGH/oXRRisTMnDLu74
NQmS4B9Bb87rV/PHbgPiM3XkFjoogemF6+V/H6nVCT8R072tFXN9cMy+juEKIJ6t
qUD8/Ehb6fCJLEBL4v14a6JL0b8OGGGjUiQHXmgs8M1hMuQ3YVG1xYHyjWAb4FsB
UY2Ifd4lMuTCfayIJtIJs0pD1E+G8HWEaVq2XPEb9SmuMoZW95LbFsw9lDizHNP3
OKx3+N/htjWlomeGxT74+k7TmNIyeFmJhIoXTN5eauY/cgclh50lfXz+5zzMeWFH
xreNBq7h3c5yXLR6PJF/KV61l5hfaxRI/d4MBPqnxfo1ibnKRepdgjyqUxcymnLm
+zxHo2Iib7yGMpVwzpOhbzwrI/1CSiz2ULxm3XckKMVcnJVEl4M6RKZLB3ySFq/a
chK/jty1JfM8LjQACxThrndVePNQsxLLW53DsPgJDRtiDoHxI6gMJDtZJN9zdhE3
862oQ97P8O7GQYPLwbJgP4cEdf2olxnKJ/yND67BjEvxi0/Fmo7XEZP7/rqxUJXz
KBcTU6FtUZl3kceUOPRBBFfmsjExJarI1KSYj7TewWF/GHsTEjRrjVamLUQHuRZ6
v1sc7q1+6zUjsF/L/9ar+xJ3eIYULjjgRC122S4qHebp87VObiBxzJMZpmk3eJk0
R8cR4+HTk8vA/jqyuCZl4lBYoDj0D+6nzDYwJZM4tk5jA4QWZkQopXZ5iQ757xGh
rHy727ghSRd8PPhhtfzNd1WA/M17xqqQ9QyuTOq1IfSu3IVaNNr3+kLsYc5CsPk6
oyc05WlBKzZ/1aNyG2DyiZB7nZkGoNz5Uapj6xqeeysvj6kh3Rmc68Yn57wa1V/b
/egL5t27b8sNcnalJVir32YXr2oXAUIVFlXVmLeqbETWrRc6bwO3ZVhRtP5tuA3L
ahMyDpYObyY46yb5Wo7UyPtX+s9y7C8WeQUISMZWZ7hOIVI9nfy1e6rnLlOt9y8w
rNFTznXXNQuCCwrW2WTcyAf+EOUydBbHbdR8OT6cdeuFhqHedI5pPhQnKZ9CX3U4
1P9wffTc6A9oKKb1IiAIO5WwL9ntBcJ/V8JfHcIu9FAiQde7edFyWadOaJjWVuhf
y2kmGAZZutvNO/yidExoByEc4hsy3AcDI45UHD9gpvqr9ye/6ToSJpTck+oqpm2O
4UfGaKqNnT6YA4O1twA4VgnP9Il9okUAItAMoYiWnmmY/GBjV6AtVaOXWKCDINoc
Nj+alO6j/Ndqt2BbhtSbtvlUZfAN63BZmsjukCscyXieDwIL0onaedWNW45f1Bqe
MfoevzbG+YAeFKGYBuYzHWBxHK/OJxG93sQnPltPdTcQ7CATfmC9se4qpdk1KYHx
PEn/kQ0M/gXTd2RIKTNj7WQUXYxd54riVIrGOWI4wVaA8wxzcfj54zIjUNU0ifdv
o3amcr+YwE9tPsDQz8TZhNcd5U3hVtGcorfbjpQZc+xC7jkb+bvhQAJvq9blUj0d
Ds5tdatvNdQO0IGoPANednv8230gtA9KPvmaHoec9RUQJkWCWE+hqsAzW0YXo/7a
uPGtXh+I5IAF/BywplinAXJhrdHl2l8uboVLBlnZPeb9/qjhPQg19NuH7y3ga4Gb
3CIUk3W0gUTKzFOHHR0Kuz95CWB29Ygg7W7qpEgP6pIPi/1EG0rJNLFrwH6AspwT
QOuBPvzR70nUupuBdMDtoki5+QuqvHFNXzjl4CIU2IZkgoehsyu/U+6fC5ctMRGM
FX4VII8IkRFn/E04C5laukSKcXt7QyTKQQEahDjyQlfWKE0fii8KbpS3z6OipAJk
UJLScbmDgR6cKsOX88J48tl34Pa4q2TyWZeIWeVMjG8vz85LhQKYG9f4FAnJfVkB
Q3br/31SusAzYj5jd7Wx44II2x78NOfrnjqua7DDp3qodMwgvtDPts2mcWnvkxo5
yXU32j9CFVlJFa8Qytu3VlIa8DgXy0HQ/caUN+T2PyV91Djx+KzD2b7eWe9yqTBB
EZZUykHIDcJ9wM4DsIVPAMk5rZMFkM2UJlAXNIzFUEbO3B627yFOZWjvH5+vSMJe
/Eb/egX0oXoWNvnrTQRp/G4U8K1vomTfdq3pc1KdW8LtDcNmb1s67XFzegLtQat7
gqZmIm/6gIG4VFYOaZzFdQUchPYuohuDQgAKSaS4Oko19AbP81OFfk2ppIKZWdmx
wOvbXsssXn8zQX8W/LHacz1Mmx6LfiaZ5ga6BydNLi9JA433KlUvIwhDOOXASrDe
nacJFmhQxJaxcUQTYTfbjoEPO+6rydzShfnhnVuDMN5vyeXe1q4INz0YfUeXueSx
3uW/FfQSDNqKwI51ZoCHsVUCTxlgzj9WV0Jk/ckWnYP50lz037GVYknycMUfIdLb
jv9Q/gu8ULSR6pLm5Sjrzfz5BlepJaxvV/Cd+Few185yqpPbx1kSjB+YXaCNZ0de
3yeQ06rpmxH0de0yAtrUQJ/N4SuyZh6xspS29cUDnhwEdVJrtMmh4ZBi+THNj10b
0DXPJjUELG8gzaYll9sKXDmKgsULDLAItdHVF2voSjZBv33D1LHCVR/65YqtFNOp
GTSSgWF1vIxqCv7ZK4bilnutBqftfP9A0s3DvNUFoQdwBLpOiId4S/6D4pEY1gHj
Q68wYPv76xNKtY+IHnnJ4CoBk/8Z0UtR/kFcuf10aEQwAKrRhAArRcZyCaZ80G2/
T1f4kG3rHUQ2d2K03IQVDaYtLMALnG63XCg1+8NqREiLNEjiUNsybzLeC8L1hXXB
Soo9vDx8inTO2WDg9gXEXWvgZ5wDu9zY7b4xIZQffMu0Qyajv0wtW1mA+8TII86r
9AwT3tjGBxdnRgAxf4ND/J9ta0+B9lhhfmfqX8adDoZnjkoeJqs6kWBozGRJBHeM
ByayYK96v8cQbC1gPwCkVt428CVTip6O5q54poxOPd2k2bytCeUcbJG4Dxihw8AP
JL+2F87mbHWEtfI646fJnzD+klmF59gkBNmTyhN9SVbSak52c1tUIxAv/oQwlAgn
ev0YpoFo0Mq3pAMgBZIGqFw+nFU2T7ADXtZRzdq2SSATHNzbptIBz6da0hq6no4J
vaHYMXoS7PWomOrwYYRBYLOqYYIX4mUiAK/HKDJUHqA5zaDAxjLnKdTXBLQXkY4P
Vhff3wFujil/s3J5V1Hd04KC1GuJf1LXR3uM/AXGGNv71GkbErggEF1vqbvfD7+v
D019Z8S/ucwLRouPrR78MLYAkisllbmy6QLqkhkrOffpwSrgSW5aQsSdSrSIoWvo
BS6FK3rS1jGt/s77WkQsI+68Pi2QN2yQuTVpCXvgCqxY4jUOpVlEq1KupQf42gAY
BzoWEXx0nXL/VQvh3qhXAqwpjgsDCxP4DuG+LHHrgnGx/uxwqcn+z3mWaTXxDqBu
eSH6yeMiC+RhJofebXPdkWLKkpEogOJ8/VuGjNDq/3zYT+/RW07CVofMlvJuBXar
Dh+gkniSdozGn3i14OAR0Zb19N0ibqMD3MnGIZCScHtPSXsm8lRTE42DoXPN4n/o
u8Fbj7U0JBXSzqAoHjTg62FE53FacQ4xnqeQ/gdhf/MwdW/+8BgCYQiVguOKNCSb
LVVERYZLuMqB5KIp0s2YRCvs6mCnrzB4cleICVRbNUPKl0HrXJiS0gw8alL/Jp4f
plt0lBp5xoNTwIMdVSNrlLAMFo9T5NIz5zoL/pKTBIzSoL3ECjX3BpY6TXup7Xvx
EMoZOUT6abqbx/M6aMfEGRC/vuoYsYt6Nm7cNjb/HU3dFgLqVdwQM4tvXG3rmVvA
SYr7B1CT3fbk0HK1EqOhArfevUfQI1es4+DOWIF+oSGpMB9HVKrGg64v0z3Efws0
ejcOS2y77AX+pWYZ0ZR0ZYRnSnvzRMeeOIdbPu2EQEbOsRfIgcF2uGA2TajP6Hcu
hbzWfp5AlUimTVvQgMgB5itrofRddke3ygPsMppg0aDieb2oeJ8xn5v5kCPpBDOB
yNolG2YphLGn/Ras5UGWUM8FX4x5rQCA6YqYc/i7LhVZrGqYB9im30zv6PpQcC43
DzLYWzYgkxQESDNZzUuGs18cVLANyqarEiaPaUMJL5ZyD3iWJTG/JVV8jY3G8ZIi
7mw+mesr8ggWFhspuY+NYfVyJ+YkHwSKNIwJ6EMY5BSHT0eb4aktj8g1IjRhmFVL
1Ot862XXOOOTOgOLwiHuPKlSlrSLtZjN5ek3i9HElnIwx7CCwFcuJSuNrlMp4Iy2
fDP00fi4JJEOHo8Wqu1jSm9Pognlxew8bgiSR98pMhX9ndRCm90HJhCKsnzyjLW5
fpGrDnYJdopibi5X8/+XqWaMRxBQxjcrhExKifz9bQ2aLPxJmqcBiySBCwfVe2LE
T6cBpXKg3hnB0wK9sSzPtud1xDSncl2iRJ/Xrb2++RUfs6WdZvY+ezoaaYdvM4Mg
RZGk+ttBior35/Ecd/t9EmdBsDNaBgAv6Ch5AlEU4lM1MrkQyRobScAkIv4SaWhB
muvy/FNucn2pOHHAis8vYfg64Mf3omCx4CW1cANeR8rWYPxgPJ253pRSBCK+FH4C
1yBpW5QNRBROkOG7hkm9cd+KpJrNKe4sduTE5nur/aoPhyY+Uo4IUDHxz3Hx5RNp
0H8ma07hxS+gJaGFJyFPGdEtLam/ug6MBZK5qliKISfujqWudnixQZZNhqs0EaQF
mGItDc44PwdTvbR82mgCLKYeF/yRvoEL6hriIzo7HGfJ42AahF71IH1n127FDN5x
7J0QlRvUTtHY5Afsev7XB7fTOugLSKQftL/pCZetrFvTxeOw+DW8/bPgNNQ8rUOM
0QSS6imUwe6APav4kAeeVumVb/RoULj/Zi+D5yZ2L3xQ7K77KDv89IQn7iBXysLH
I3MdC1lzt1sMS7kW9Frr8BnNyBLzkpRsg21/cikPxTDN0waCifgxvF4ljoJJFrUf
juPL8cyrbkUMvjmZNA6O8XVwNRuu+sEoIcBtbZMUv+GgVbmJBUNWk+/MTVbBRjHx
QwgJsWojjTzhISTqCMSsNJctZISYvOz8/aH+d6gC9DKlLKQfRpOBXCY9lfE/Vj+V
TLJa3RPGvK4xNLz+2u5aSuW0N57eWcn3zK3hjmLV3ociTKXsR44HctoqznsyL1gX
byg3sWnEv7xWx2HWZB4j4zDtt/frnKCtivK2+lTngbcyTxP4Xkj06jV3bGbCQXiT
vxWwNULmF00ZsvstNrIDXYwk9699FADbuqliPKFGNrFSwOYFal7+lGnw6bR9xfes
QNItzt5Q2hQwxbLcfaLj5bd0Fw+owRQh5a5d7B5lP+3Wysna8GGuzmxg8zNOBf7x
AdkuBMC+GDFPZIhDIJjnH9ymePAMLlrvZwBgHYRxlzFc359HrxMDfvMhvTfCYGLB
vv1qVjuEhvqqDMllY4iUnaSSwe8CuV08ojyP12UpMe7QmuISn2lnZL7Da6X6k4o5
0EtJOoJnHTn/TsDioOdRf6lHxL9p5/Ey2+B1Yzts15GYlQ8rxMzWSE6mXC97OJcS
Yx7apSIL+C7fGDY3YwIzZ9l51uqdaqnocK71opiyiQ0FxApHOCC8QAHAyCq0rb8Z
OKXhZ7F0wvyYIUM9NF7xKG2XImvGeNHh7dTW30p+6JiwspoTXYp/NZRFIAm4HLj1
+srxXimzTFCMUY8JczzukCqmIGwSzydrfZf+jXceP6bjfhlJq2DHqboO5hcFCNle
GxYGGvoXBMCz4DDAXNSmeiUYdPmbbIyXTENjZAWnJj1vz3SqaLKhm+FcKap1E15A
NWR14v5DzjIXaog2z0QoUSxuVUu1dcUgWw7qfgu0a4UI/+DpHiJCsrLGKevoXKSe
/MlT1kiMKtcISI5b2TLFolvtBZP9UeHiGVTbJDevNepoNHR5Mle1AVjsqpUv1Z28
YwgyE7C9+/V9z3x+JBXWWGpMkV69rl+tbc9+Ynde7JK9Qp7juZo0jKsOgZNu5W+d
fXL/4lMU7rd3/7yNlcUYcuaHLxpIWWH25mi8eOGujF2I9Hr1DNFmn7dhZ08Khs4w
ipLX6dwNDO8k7wJh2lScF5yLzJavR94QUzbGYnw7ele/mpzm8KpWoRgNRMtRcMb1
KOtd0MUwXYLLe1PhIAIOvB7/Jbtq7T2zARkgaUzCRkJdL++73dZMj7ZLIZngtAg2
2RNH8iFIjH6rt3R1p9c9elDuhw54Wf6Cq/EJrhRGTmrnngw1o9RgQ9uQQwjddbFE
dN66bcKachvRBTnrozUklD7bvn7yKzc8fZjx7sf5np3Z2nHc674DO57v1RUnTvIc
UMqW+8w9zLQ1Q293lxEyVofKtx+bM5ffQSgEaVKl8efTuFu0HMiuoNCvHcq9nkzx
XzxlK+aE8q32hOY7CHxM66S6i8Q0/v0ISOyKIPCXwtoTTxhf3oD3cpk3x9f6QzOd
QWadXag5tPzFadEeiYHWiaR1esev228KocozYsU9YKfNrG9HtgNec1PaJUZlZoqp
MXcQo4d17g6H+EEA80BbpP6Rma/Q+7tbaa2OL0HBPm1aCYNXMWbCTyhBjfZ6p6F2
hOSphMeGU0PQWhasj/iIHF6vMOHW5+HaEzd6V36pCIZJxZn0Ik4seiyHvm1Fj468
PRHeZm7N/JzW/aj5q370qyvbauJjbE4sOwQ7G+sUUxv+NZ0OkqHT6Vmli/M1nksN
dZT53G65rN49rxTRrp9OSHBWSL6yIGdecNAqadIlbg93KlWwEbyvHisw9F5brkaD
2I1Rf3/Gx26Cf3sngMi9dRz3Gt8xwXIIt7oyxa5ydaC5QZMW+LYghZRNXuSahBbC
jf3d2CeB8XvqXHOSSfnc/HIGKCQb89m6DcLTfvvnEgQbSffzaOEa5JvltTUptlIl
n6dzZDz85tDt5+kZbL9CDQ==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
d60KE5pbOyYTOjgTFudL1JDeR7i+8F0bH7qKYJZGHgfut8+ZW7+VATWf4VH7AZJz
FtqeEAIZZtnuCpEEb6oT///F8lFb3uYzb9XZ2cVtLKXEig5uCEfDUXid1/+dzaGC
7tymCj3jOsj9n67xOGBIfw94TJPcjcOPG6QNSfC0dJFRo3sYVG8EA/52tATaQr0v
X8G3WXvE+IhQNrC7vBHef+G3XRhAKKNjzliqpvLxaOk5Yg32lTMfYkfP+qrRT6hO
9r8Q2sgjjKSDdMgC/WKNwGia+PbmveD8KsEgJt54j3g/I6Ly2Dif15GgpqJOQEKc
EqB1Ydq7gNpPNrOdiLyRZw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
i3IcqQr99BtgAlo7hWnFz4y6T921EOvDwvgqkus5XK6t9wTvKT97BLOtZdn/y3B3
p4U1y3J8hBOQmBLimknhS0J2tVldN86WohChoz23nay0yhxopopKv44FxhZSttEl
pqYBd8TEIL2brH9d0QfRx4vocKVLODfNyngNOWXpe+2TkybWynteNWpT/YY5JTDb
rfhVTvlMaQ27B4ycocsUsQVBNMcXIU0g06qJ/gLKTtO4AiPux05Spvjf+6VpCbL/
oR4rptZg3gpq4Il7A+vliSG3daEIaHJ32TJh3pl9PunZL0xfhxjQpUo0346trS/K
HaK3GAS1lTMM/Ojp8qitFoOER/Dl0Ts4dkwaNGIKcXbJcoCJq2YI8dsHP6XfvIh4
JRTAZXK9ZUIIEf5PbvjyTNil89Sr5w+OrPN+P98DYsPs2ieSQrxmLX1fUnuAaPIW
5Zg+UwNGoCnpjhv/UaE1UoTawJUFEisQDARbCHGvLQk6+vCAApH6EEx9rWGqe4lT
j9p4cvwnyuh3K6F20H4y2izSEOraoOcS904kYb55q9HW9iQYqQEN8Oe99pMUO+nB
iL2VHijMws2g3gRU7g/FkAOig5ozLZlWM9mwzWsX2gfqSRMuBrdw1Dq+aA1DkhQI
xykv+43dEzuz5YNiHqYt9hKtd9GkRM3cMfp+uu6QIXPk2hSotAyuRiPVLl5U6MDJ
ITREn8INU0gKEXJ+WT46+psYDQg7hxV3hqX8Fil/LRJrrYBl6uXuryQJaydTC/DV
1ovySnbvKaEsKVyPZCkPSdfO9uvWsAI/Yl6NrbcnI6HJ3s02YFdmtLOOD3E80BB7
1faNN7yKhEs7cTgN4UO0RbhY7Aw8l20J0uoZksOUbO/kNCHfS7FPZLSXlnHLyMWG
Xx1Cndjek5VngS04d5xJctDJNKYe/3VpsrNi1WEI84ioXVvca6sgJCVS82m/iHPo
4Q/QcKf3Z6p2rw1zW2Tt57QtJPQxJqZD6JlGMcMMfAItU+i2vOeGMeNXA8v5H7Nr
0iZUFtw0W91nCwzIspug2ueIxm2FZcDYY3DLO0JTWYjc8kpc7/62FiNVtgyaCN8Z
pf0zh9+CNpp+LBNxwquh57g7MqhA8VUEPI9ryMzgRFgSRC+EuszJ4FaTbj0U8sbV
Ym/sAjbd+T7nZmqKoQsL2I8b44021VJnhw38yWGJA+6R3+E4jtxdGfsckT4hoLgP
HNp9lqUZ1EflIH+85xaJtSzghUxiaqbgvtLx2kxOTeqCJIvRYguqsZICbQnkDiEX
FGIUW4If7KFXfVLoAXBiSnkjqIZVeHg7dzmE21CZsAaqp/rdKOrbkY6qQ0xf1LV4
FB7EvtewHr9F8ZUxb9cUN1s52fpH2sAQZxJfD2DCkRxEmEEmidyKv9hhDxPIMECu
RC7oT+iKscha/p+FLw81unST2C6/ZavQtbc/0hJ0CRh6pmT+xwsX8gGfMeIq2bjW
2V3frinKV+KriIQy1GdpF/5Snkm+RHvWHpiLdFUYV6NZTJeLpkA+VbFZvlT7C0aE
qIb/eyWzi7J17JZMb1SR0FcAOChQgycyPE75NxdoDLfrf1qd31Mm7isvg4ORAC8c
DWPGY7TA0/2UhXRGnde4MziYLHUyIQY0s5G3UyFFKvO/sHz5cNcmPV/So/2vmjwj
iVocYKNgHYobISe5199aeeiZjywpFvOgIoKX81YEuqaRGqWJjNg08jeQVNwHA1v1
SJVGM/v+TIOFwtn0u2pXs7kCyz9CLLKbXO6YpPA+O0tCXu0o5qblPjlAtE5SxTOn
QKE3gTx3caSc9tVhhRgcuRQ4AzK5i0M4CTHGbUivrHr27S2AO+R10L8yvGEaPKSV
OhTfMcgIgE7coQBD34J1nkVqi4lhuBlpsPJlYewAuDqc9hovwy9HrmNlnZ6oUzXc
LteG9oCFW/hxiqTSug3orITnujP9lyWbqvFFJqg9Nx5PZK1x9KIv4ISNrCy8aqbX
gs4dZvvE3/MP0Q7BioSLe/WNG9kvu5YYohbk5B6s2iBGtpcYUb6jeNFj9e5rOXgZ
vDKcnUjXZw4Z/WSEwZ5SJJKqOn+xgFdFkcVBYto0IJk3OscBB2yJegPa1idVjhg0
3in8t71tjB6FZIcPTsb99XXk2kGUjCkAIh1m6ahB7p24JJVfbul8ufozYUCs4mjv
wQYnM1m7WpEvm5rxQfxekH6+rKOtGjo3yszjzIiCkh2F3xRZsoBDG4ADoX7wrKXh
McCz8rG9fyf+aaid/VWdry24HQVYuLTFgVs94Zi7vok1dMIM7oCHk6PitIsQYrMQ
HWRM8JbV8RKJxnCFkNdeJaD+QQmsUAibmvIrQzbb+PcI/mm6LMd4pqvoAXtrkZ+A
AFfD31CXK6PDuWCxwzfmYCwaOzsICbnvOOlaIym9INQmH/lEYxOx9cXQOwbLHE42
I0uUq7EjRXp6kj3qa7sKY5wKwDr8JjU59gLtiJIdV75redqNHEzI2ak/v60wVhVS
Sn4uT6HoA2C/eTJg/4ro0LVNVlZXiC37ePJ3XtmQgjqfKhJ/Q0bgUXXL99s8REVr
4GxdHuLGFOiLFAevqM1oWjWktDc+teLTkMagftdOl24IwFJ01+Bxh7soX/wEQgGh
jRv+e2+ApcPvnR3bQ7eGIdC26ysENgFKc7aPjavAoG0L9xtM7j24ojxIOQq2cFMx
z52SErutZfEOPCtouv+2jzRrcKXlb6WzYlb+fy+fYz3lUgGtDryweDgU2PV0ibKh
vR79NUbHpGh+l3EjNk2TnJXumLE3qJcC9BpquU6Iy99Ixhp6vnHCCfFtAKY8ROz4
WWbYBnr6HbB0dpVounqO0RQvpC5KZHaAoCn5ctn8ahmERIW+Uq6cMxC1zd8uexqt
N516b7SDdcz+R7t+BWrWWv5HgFh6cwLumGC4T26q4nUOK3/ciX+8AhhrP9zLnXsR
MgmQd6XWS82OhKjBVEXCXRxOWgDW005fq7IKsfGB/4tC4snJS65AfDenIOtaviXW
c5pVBQCEWsugn3T+R8QG+zUkTeA2loMREHIlCfpBx+c+yCPMQUd4wfvTvvSQOgfK
PsciwR/JS/zgtsu2DsUqdE6+6YUPnBVCeLHICJcebKQlNt11Su6pfI+xmTP8LpIW
u2LdVF59PBAzTcudbqZnU5jsWfT5P75aSh5QtWw5yDoyJ+4fNeIeg9s/XScFmCnp
bWX+0z9VlfqcwF0tLQ1oF5LDyFwA4nbbaz/DFozJzmIIAT6IyIPhmNV3Im4UL3GV
q8zwSrt29PN5NmtyZdm8C+bdzbEXjS+bvnKPUr0bywDhjotaAwPo6D0ts34tXI3r
ue89h9ZRDDe2JUtkWrFqCHIUNja02Poh5po18018wQMK0BKK/xe7uf3Bnku/842q
uCvqgRwcDcxB6caDpm0AxaAPmNzApX2OX7jrizzpp5lJmoCKxcfVhhVx7Mu3Nr5e
VDj+ISKYuieN74GYhMQnSpLT5zAe+G7gDbqPyCKBFXVf2zVOxU6VFSuPCdUbJqA2
J5n3nscBdnSZ2gE3CFfsEX6y0JC4bSEiFBHOJwhTVwzTluV29nTD4q7EX1+AL6jJ
PEtlltGvVx3ZoUjGCNenaQL2MS8OLh3A+crhoFYWXfgin/1geXc9YZGKAAYaQOiy
hIUXtPao+DStd+FycQZqxW82H+NYTUG/5qjVpo1ZWYwKhT8Zsj77M7/hLIbb//ZI
dFjqdghM4JZ+ls1ISQljYeFGdbnelJUcw/KRm8VyHe9kNYOhaSMAdZjSNGU+px67
npDlebOmuZywRHG9gsaiK39PpahWKt5Eaf6hUV6hc7ywNTsuiuTyvBrcWh0VnWFA
H5BzEehk+buNR8UzsDoRKmHQ/E/OxxXgET//k2RQrNkGxcraSpgzvexhky45EFfN
x5+AY6nrE16FnD3Go8Il5e/GcwEDpqRfoHkTElTjauR2SND/6UI1t2iu5nZsh7co
yqYizWqbph7TTHG0LkVtp+bxv00IzHI35Wci1Qg9SXK5wrITIxXDb4xIRGIhIQsK
l7P7fxxFaL+drqSPZJlulp8gWdpxTtNIcovlfP5j+9qiqwzCkLh26s/e+kZMYZLQ
nMKaDIxKd7Xf6TKSmM+zU3k77a/XeqENS5tCiojDkjISdzC9a4y05Ylf7JqnSi2B
anmjYGs4ZTN4xhIqTYbajX6NlItOvWtL9qM/g+agA+Hky+6iaYl0hwLcZSY7FSDH
M2gOQvq1gB6I5tusKQuEMbBfsO1MSa28FO0BZ7Vd/OovlNwF09KxAFnwKHfZFwWC
GJhd4nvMs9H1XEGVcFnNVRUXlVBNAw+FmeInWQ1fbbuAk6/pZ9eJ6vOHtEhyNrKu
YOOoQzC3WoJ9uEfd2NsgcO7DAj6D+L9TQYLHk3sZ28vEXUFu8W5FZL3cPv5l29x9
vej/uW8ljIpfLv/SLd1bBkdpoUPDSafTljGGRsLK9cAKB6nGPSMCsDSBj5qAWI4b
dAdE9xKhWT0eyacsOaDiX/c4gmDbcffDbBtmTA2YasR08Qf4plDyr6dcysF7beZx
9SUH5BTTsNKnFowjQ7g9XUYyYQcBkVPJ+LqCMqaQUalX2NoH7jc291Mhk28qTBSJ
5fg+5mJ5IkIdg7zSH2Z/Jz6XMPETwMTvAPsp08CJreKlQwomGpOMrrPEunSPxyCn
hX0LHUuB9jz1TGmbf20MYap0XZmwYTfjy4XwORXyFNQfQWIFxb2nH+CSeGJENPtc
R17ByFGA8/zLt7wH6cRjwzADlG8lQN9YpqO4+nqhmXQoCeF3AKpjyf7r30xas2ky
O6uBZ3IKQ1CM/EwLxf5NVRcE5w5ffERLyVcQI5xHdPB6foyMXuHJCFxQVqUEFW9p
e6YiwGpNl7lG73zgU8WEoXQ1nLcpS8UmabD/caPpXoMtFov1Bukwkqb0nY6jlnRu
Vj4F6cAZN1BTMHthjUwChey47bJZFOq4AG1DW8vNRoPsWJDcR5jOrnyHoQV6QeHT
TRcBuK+xWiQDPJicQwSu/geUHJuprJ9nZkiMJmaU3fcvaYQDfMlysyo9mx/HP4Vm
OMPB4OLa8axk4R3AfY80JEYuNWgiP6BsDKKZKM1h6ztS8F+WDwTUp2KIRU3wJIB4
TSIcAo00WY/+TXhk7Zb2YAQMNvKELOMSDkE+s1UNHMrkAabXIq5UxUAYPk55atWm
JVT59pe5a3IZKwUmKCaf6J9TWB4m9rxm0f2ERKU+bs/P8OnmRZTlAS55OTqt/3dB
xSlDSAUGHLTogNu0XpqOBryS9wYM5ptPwcz0JvzJnQqB3llYCXQJ1N1r7WGqTE6n
dC7HWKaenfJzfmiAkr4fXULM3yfHFVdmtzzMmswDkf66CoCw8oTXaPoqOIXIwUGT
fYTNWJ6Ve4w40Cqm7PGyy2eVWFYBdNjy/+mMeaNAB6DJkMzfkXFC8o7jxGAxe4NM
KggrNG9i9mk5BS6bWWnaLHYwU3F7i505rYF0ITkeG0qKEqBTc0HsiM9lRA0svheD
seZ/tjRbKqOSUTbi3yfOyspUwvms0RNOpFAnuCzvhzt4dGZC+Gnr7OvinQkhE5v1
gMsTd4FNzw8lOPRlFUJ4enbR01YmX3ITYKJtWsf6RGHkMpTdwd+W6xCcVNoSeiRJ
e00GUDUG0Sh8ffWjQBpSBNKIcYPGSRhgNJ5zZqzAi0A6W/ZapSEgmAHz6VrrImfR
M82+JvN+sAbyMBIdgfqH4Wc4539LUwQAhXaNG6Cq2vR2X8zjxvlNZCLZVSTmIv4n
mwcvCFNhz/sCEd/BulSD6jsFpAtU/S4ZdPN2jrWZFGz535ttuaWXYMgW+u21jBM9
iWaVV+G0lJIH9XuqUtTQ6uR8DCoGXRyK+JI1jRyyDOIwmjir2kGh5Vlex+BIr51I
HjcTn9ipu5anfUJ/gV/kypZQCDT4hcufGB5Y40nPpaKsDJ9gRgoanbggtPlDBZgj
UVvK5ZEu4p3ji5W2TxT+SjOmKHbqnPGz8n98q1L7JHcCd8gej/ciCwvApX+jWsBi
5X4psF1zM6Cgl/IhpGyRGIdiIH60aZEPd5ZgltM6WdhF03QXY18RNfLxanOIN6WD
xPvJDjMa2ojaR/Hpyzdf/H4cWPLANHJTnYLmYYC1Rx4eNGmzMmsosYikhFjmgQLG
OxbY5OvdcA3nxgpdNlA4c0oa+SFO1YW2NfY6bGlZZhfjSEZDHqc1ARujbcP+jjef
OaQ6aDIHQqMVp48kuPjDiAmEnZLPr+LciST0gi9b72P6ZogYFj0lVAZE/wfSCQTv
xYiB0XuBJ8wc0mEmviT2yDzxI3PqsFZxVwU/WVP5i/K0vW67rBDWWzSYxtE+Wgrm
uTjc0GWUskuW+rkXff0zl3GpO8GPzBkUviVKpkNNAU08NKbmzDLeVryOkjcsnKEh
qEOCGJqVKzG57OcekNqfE+/AXD94VJRBFvDYwRTBD7lnh6UgktW1I3YMUkZIkCNk
dXx9Umclf0OQ7g/FdiPCm0kDEgp17ZVlNaGGTa3o66JS7TrJn+J8/KgHeApWoxOp
m2NS1Ge66d14vpAW/OIny2pPUTV/yVfPVm+sh83CAJXwZOF1QTTTIrAKJmIg/TVk
iIiR75i4FtXULIA5+6TCgJQR5xkGnOgnFdm2iUJ93VIhgKibYtc8L3M8tSLfzxlf
3FBpG7cidmT1fSSfkxJ5lg3f0zzF0EyD8nyHwZ6mOF1FX22MKHxgiaoKp2UxErbT
wpwFlnIvY62+cQdLl9XnBubdnNLpAxBfiVDpDZfeBuxWt5kxXfjJC00sH8mhbs9X
yOyUw5nNS3QPmElhgZynLlEItjwWwEFQr1l/vIlNSEDAT5kqJnDLVca7VzVDRknE
ju7G9TkeHyGfULOIJcwNdlf+Aj+OYezCECou9QekOB0EBkaaLwJypJRC5qQ9SWaX
NRmcPywmv3brgOzelqhB3L6NGotOLJXACLnE/uzOycBOTVtYiYS4cs55p2qSNYBA
riitQDAkrD+GldQQtm3/gISeTTpxCEXH33+7YO5EcG1Oc9LYiqo+NO8iaMR76BQn
dCrF0G9cc6xmnx0LM0tcUInIlT9EnLPuqHFYRx4TvFR46Iv/ZAwR6+dlQrEPMNba
VyIM0ecUL9eBn5zE+kj0455hO4XMDHuLaUdPN5TbaCybjmEaWUoBtQ9tH+mbUXJb
jKwB+8bml43h+SjERkXJlHJXcKGw0ZeMhZbkKrUF7+37mXCtAgwEyvxDiYWdGHta
/B7VvdMsOZZLWN5WnCMM+KvRWJBPQQl41kRNykgUJDFe4P1B4hHTcI+K/frUHAxE
ud+bE3c/LWHblpVhL/H7SBDJO4KYg1vKGr89bEfai7bvYXDqvYC282aMqToY16DH
2Aj9OiU1Ja2dVsMxTFFUjcJ9lBGpw//EO5fBUsGXKHIrQNwSK96/Wju3aedwUf9Y
dq/NQThCrZzX3a9lvhtVc/dmkSGbaoHXi0FCaVWitOG7yL+RULE35h2VJN9Ivxxk
4bcJVtvEHBgZdaErUmx3lQQKjpcpG11iL+L4rAVFhBs9vAPWxwlXLm/zZRilYxRm
STmEQOqyhFGeXTS7TY4r1p66GFHiA6AS34KPFCsNLGB93aR8xNKECLAqytu/HPe0
lJmjmkY3KA3IXG1O2YLGsT6nAvJMWdtTm2k5HkWOf0aLt9R8i9dPngHluLZM46ov
hrSMsB4BZ64Y2ZVdI/OhJYULdsLy5inzm5rHq4p3YSVRY4rx7OMsNhC04LE/cr8z
qeLh4wG81/l4lCLDXXll6ABThlEcFQaUzZXFkVHGHMyRh2YsMnZZoeHpsjQ3konJ
uwbERD/esN3Q0snuMvbYJaaWntbKM2dn9M/E5c7wR/OJJWdE8sZ73q+OThwxI63S
x52qG9sM9qMaxcBxmRgJ3ZgrDufheXPxnKugNAp+qB0CPCpxRzltH2pv+10IX5sK
wyj5r3jGjn8Jwp76LP78Nj/w/062EuPaek/DoEJr8/w1S60LYbCdBkvDMNVqFani
UBLu2G4pKuE9ZW1u3D1OnA==
`pragma protect end_protected

//pragma protect end
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gKUD6r1TMZxFrHsfnsEk7xSx7hdJfDdWHNjpcdy3uecfluvDriJg8c/yF24k+Gg8
lzAP+hlh+Tgg9O6g61N4Ppz80obrs2IDDZo7YPX1qOqBtkC93U5vFobVQP4foFUu
t8EhepM9h9hFjqt67Jt7IfaeFDCqOVra9YneFpG3LnXr+xbEmCxeks4t7MinUABk
fLJuyzDlcqf1VW2wZz4l00uRjheNyzzDvjZut+69Q/YG/45KNptHlc43AIyBOLYf
0vC2xUHYVmLtBjPaV2u8xaPYQAqa5Xd63Ri8w4xcWI4EjeE3NtKF+fgfUKa522H7
2l+vKkw0mpAccttL7G1pqA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14512 )
`pragma protect data_block
lAWmfZ02dmcAsluw7grcz0Vy92/LwAqd/ySHcUUAhJZG2S0oJeNb7Z5k2115MSRL
/U31oxHJ7u404FJ4wVJoyyPSDOjckBtLkRS95vewVzBjjgawJeivVUIyL4TKqmOe
Ks1pTl8qmMcOPjQwLFPtfZjxQEZHPto1SkR/5ZbyYpVbK269uaEVOhPeuudCqf9j
mIJEkRgwXvJ+lgSse59Lr+n6BQDlqK0sOExWKxlxfJkSj6KJzUkFsa2Y6rS9AR5N
QfHIfWMgd8Gk+mLF6f4I3Xu2R7LWypXyyZwhJSO1ByctVgLstZiSOhzv+RgwxXSX
PDoUTwuNZr+3fg3RbCe1dyhn6QBJ8lLjs0dAA62pScNhcveqFhMnWaVq89ktfALG
g9utqSWU+4V4M4LdbnXk456WjKwjo1d0Oy61GOX6As1AkMTzVfFcfbh0wuq5x61Y
VJ1rPFaoeNBJebncKy25+v/A9OFFy9oQ1pg9WNnBajqf96dMtCiVGf1cqD28OcDX
7yayJmRaGbaiTzHBz6mby+9HLwfSN37JJ/CCJLvKQkF+Nr6iN2UNFuWPdCuyDd7A
XuX50ltycFyGoybU4z6Y8UnJLipWsysllNqUv3P1qnuBt+mma3f9A8GolAqDUIXX
TME4XX2uBO4ra78EfyVaO+U/rZ5+ovTj36qb1cuvjslnwCQ2EmfIz/czFVYWM8Ui
G4l8F1+2whY3QX/GnMGUtINhdMrVv7HUHLJFJckrdXsota6EqGS9ELrX4qv/dnIL
djoyO6ZWSLX+PTKG3SN7lWwDG5hKoJylm4b9ppGb6jD1QPtAoVu4nYha7FTnOUVW
zk42ixvci7kRQD2Ppp5u6z3YSAFtRwjg2ppKvqaJ/XsFx+MtA+rwe9qomoENZCnc
I4eQrkh5CqNLNp0poFy1stX8Om1/OhyTSofKUX8zxFMo9XipXOU69Px/VREHLpLe
ERHSlvvINYF4KYN6Y2vZPP5wm/C3/1TAMCbVXdLY9CwHuL39YcxnXnysXsE4GgeX
7ophqwhBbnTvUnPYOaqeJdYDbIbqv5DhrQ1iCaRVSeobiftayA9wb558cPxpcXVn
IM7/3Z4xk7fvR9gzE6+/6ZQJftAkVeRDqMFgeeAxggVtz4PkhvL1uN6U5qoELU2C
ZwUNm6Kx2oMvONYwO5nMDlYGzFON8mchIchWj+JnADzwUw5h2fLUi7gO5+AT71ZD
Z1AjLfOiJnliEbvZNe3xO8nt45vEa72UAmSZcL7tQTJQdH03r/BBn/UN7XVUnT1P
9PuHcPRLJqNRgzdSZLd8tBcmM1SH6tZ8KxheX/BVKWwmnsJfqD2ZaPy+awnC7w6f
S9bZoUdCehGMg3JPCyXr2wfr0LYrfMtlTrLWVDZ6/jT2x9WU4XFM/wJcLxnJtNOd
N8BUfp9RZXCL81+lMS5AxmUU18gm30bj2EzBPTeiYfD52GfQ5u/ECigpYSWIpOrm
QQKYigtkH9CKlKiWh9rjt227ODO/7RV6A5ERjF4whYtr4RqBQVmUAYIm8hVGYi8C
0oh1NE3DwKQIkt7HKongWDacCD6XYjcXgKZEzqI7L6qP5UJWCxYT12mNsFlRdjfj
ku37NsBN0wSsCcMJKvSA4ZI2eQVFEIz/sGisk2OD9ex/Vw1LGkI/5JF5enhSyXvm
iuLsAb2J9vymDFi28CdgL/hSGdFtJKdGWRUycHdtsxBuF4LRXUhrjAk27kbQ8vaN
dGhix+vpkO7H1UiUP1Y+nVDRLPPtIxA9DavxhV/+FIQ4EQZkd2M92qV6mNMrQeEQ
iIid0OJl6UrWNx4HoriqDoftmL0fwijx8kjy9E0mcJsKjXflfNinNxQLIDwng25T
5Ads5FCHVIboLDIkWm1IqeSO+mCg1qpSg0TrS1cgjzMUfznKGBk6VKXQAITAP46z
vtBaqCQdDiDqv3oYKhA+Aa5xNYQpJl1Fu/tQveZpqBXzz5hQyn0rB50HigQfXyiq
caKAwdjkc52kunYPIHpoeNmNRcpd/Nq+X0+0h/OhC1mBokxxWFbMCBGmXbLKAL40
SNq/lJ/d647GmjQNIYTrOUiX/uQvKg40ae6HP0KTQVu1WlDrLaiXY9LRlu76RqTo
XU72qIoMAXJOAKrRD8Vw+ihAvmeiu+QOyxL8LxJKbtB87nckPay5yV5o1pVYt+Gv
3q5sMUkloOEEqBEKv9ZgrD+X4m+LLpwzVb+/g/c0F+zFztq6MzEWGZG/+zMe3XQA
d3ITym4qxDPHIlT0CQQJxWQSevYdcSuYGhPwQJF6Ll8aqslDWTAnGxmtYxE+MORX
c3UYtMkgKrV3JQQzaWkl/rvlJPxdIS/KrruqwpZhejVPHBQVA48JC5rNNOjmSb2Z
Lz/gHEc7vwt5bkXu0Wzf6OCyQy5s88qW7IG4ELwsncx+ke+au4/cFp21LuSTW5ap
DC87Wo8TvmgomHCTo3hDA8Z7g2+G7ki9zcgKgSejdQznI6FLZoD8ARLinkWg1GJ2
97iyZjRjju8LlzVNs68oo8rdgu71fFfMtifM/oHyCEwe53wsQ3bi4B6LnSvVrC8S
+wAevgOUC2s4QSS916V6eSq0H9GX9HbncgXRDd3iZ3ZmnGaykYSqTGJjSeNW9GOV
sOzHxx9VbRglKwNipyDd8YE9mARNsdf2RmU5RDcUKZ3zbTZfJwcOMjWA+R2cltz7
ES9Kojjeg7ek3/msmiA/Sr18qB0xjRUwZxVSHRCXPklh8s4xgBnsOEdAVjkeLS8H
azA8ddWz7Qd6pV3aYG/+Ma2wt4GgsZ+Qm/20NIvoF4BKsrw97x/RUTmQH2SDixhg
9oNBKxpIbVR6zG2x78pYP4KBkADCc3FaHC3Npzg++n99RO9OLV6Zo0QzwLm7MPYx
ibUV5o1/4oWkWFIaXxp4vwunZiOkMVGkeNBhIF4QsILZ5+WP2rksWxrI755igRqM
fyy54L5lMgeclGOEcRtSELQKAl8ZiLBPLJVWbADX/z77Std+KuLBi4skRlxh+xlY
pBcaD7jBOfUsYKVJz0QVbGCAZDX39Zc8llF9CotrimTRRbpgJ8fLP5rb3ByR/aQa
ZO7dVucoLObvVpVxzht9aSYxru4rFZPXQ5zcOl1RlebQl7DP/Cqf/cM28l0bgraX
+hyhArn+yFMOqqwRUXY+uq4uh5FR25FF+DdQyzXWkFPlb6W5Kdbnf4GksuMuxv6l
/GotBhEqP50t5UnA7QycTOSVlh/Is09c1Ecr/EBGFHm/jDCeOGd28R3D3wUUZ6A6
iQEjhN3WidvBTwxeZaAyg2zXjx8/tyJwWBQYh3+CuFAE1oHjvCxFPnxaqE7JJghG
ZXmjaAK0P5LZnFT3dylVaF/yzoaWlm3+lyw2oqW9F2GnFydOG3wcASfJmSXclfDG
oyuzIy6Kzt3w/XdVDPO6+4iUDnPSEu1hnMTC3z/Gg70aMZ5d+vBKsL6qC//rsJso
54Pi+0OEszkVnXDExWtMECd24w5DaPk1vSU2BDkXSS1Sd/toFdBUGFB5esQMgfH0
IXeMa60GQtCf8/nr2JQl4samJZk44rmEWTJh6uw8PQoRU5XVDJr9pGahOuyrp65t
NOe27ORFMhh2Dzy2t/Fz//FwHxY5ti9p7S75o2f9QS118TeFHRS1jzTW6CdGABeA
wZ/JpVEjZGIreQFbCB+y+SovrPPxKp3+aOTtGsR3Bxm64Bo2NysbjSy/CeFavN9e
edc1bd33XvwYPvAAQPRpw7BUKxGjgu12cKtsIuV5rpJl9rh+jW6wnwH48ObD59XM
HjS49Lgxr3YgLp/yIMFd3opYYyyy6H9nAZcgvfHTBjxS0lano3I9Z2+rzOW5g4QH
CsrIHoT04sykfGudNtE0HsfeFKqZCI0hJEBmdiYhcfWUxLtY+0BCn0y5AVli4TAt
bVbyDwZslKx7JrxpwPwKkafQqhjA20A2xpoPFFny/LQcqZHjfskw++No/xxTp6+z
xRiApzBxIpXIm7zXXqfNvUzMmP5bk2cjNugBLQughSvIlZeLfSsdx83S7jUIyYxo
49cUXblC/nz7hfKLG+5LMNm+YI41XrI0M9N4NvYcwcQS9RvIa7jILf3dX4Lx+U+D
Bva8A5Eitov+68kUIvcIyue2OXzfUO4D4DvYybrDxDfIG495V8xJTuRfzu8sDU5k
LtIPh4fYkVC92fRyY8B086odkPvUDFYGnfmLVlsmv1hOilDFU+WfJzuaqF7XE+my
uWSC8VzXLwV0y6cFXo4FPhmFUvmqCJ3+mBTpfUO2nt6f8zlEY94iH4YiFfasgX+Y
mXwst2kytQjhPf2oH2Rw5g1B9jjU6a7y+2NCl8xuxc9oj9A12LTRbO5WW8bNQEKp
DjLyNZu21LwYPqhfuSt9mXjGVCv0yhJnA+gKRkDXQ3Q/Y8b8gK1uvIkGlzwwiimX
n0ND3EzQpQANjDsls0ukDk9/xbrffTfo1TgSISoZKNEoEuJl4nDQF4l/8rSC3579
Em4sdE2IQ9tjAlNQvggf0Ig48Um3BjEN10LPEi3IZkfR3EvktYKB9FI8yMfit1c3
vKDOyJDWU07/whZR0bMg126hgBoJJubwNlpcNzkubngWN7hebRxwjBHZzAAW59qO
nS9DWeTSc+roh5OyNewMcClkn9Xi2sc+JOLxXzC6qp+uPa246IWZTatpHB49DItx
tLgCZEe8ORyzBbXmW2NhN7ijA8cw1T5JTt9XxEBTDHUs/Sv0ykfXqrmZVF4b7+/e
IvOC8gZKeYjq6JElY+aPAD2F1ZRtiHCU8I7oBojMwJJRTie+AR8+OLrjom3dSCtV
B3TOGed7zeu8Am9JdeioYsJLz8KNfN6J7V4TxTSJ9dkdkheW51X5VuDaYtZ+6rYs
naG64WB5jpS5K3eudW7p6lh7m5LEmadEhsP/eb7W9hultanuAFqxPWa0W+PN/xJ+
zKGwvXnpW3p4HB6M/hain0fbsRsdD56S6jf3enVqZuBZnVW0K91QJs7zfP4bZdEK
G/iSaqV1+3XnW5okcb0B6/00+a+fLhm+QT8Z9oL41NGA3CfM121vj9+U/rrHYZP+
mEwLBJPmbLtBziB+3N7Z4Ezlzp918v6LsutkY/Z3QhsH5CYKz3sy6hus74x09EZ4
Jiq/AOcCJ8Bwkp4/njA5Ctlmr2gs0wCqEzIf2zzRZJl71jyq+3P4DNRGqno01hXz
5iFE8oTGZBvwJJeJ728eMxjBGWcXBj0cCBffAqfbwhxufaCA6XvM/ObWLN1l6HbA
/3vpvUwgDUrFqBQDSOP/SNZy+l0MgYmw4XgV1ITZs1gRLgRTy9TeWtYb1UTirN0n
cwmbdkweW/+sWHQCvqjrWGtyZXsXZyctcZHOAO7Y9WnYXxxD5Wvban3DRQoOq6XF
hH47sUzYyLK9pmGNiGOhWvh6FdVec7qNIdL+UrvnEo6jnr1+YrHfX8FrLRSOHa/6
q4rIMUOmYHjmmjZcBrVQrMPP9BH92hpHt4GFO2cH3Kyk7VMxXy1TMwq4wQsnFRRL
Fq9TppmKUNNyZ6xCjbxdWwAY3BOOUlBcJsUECpp5VGAp/anN8q6GM8t1nxrQqrHU
j9PGmNJaZbFhqEj2B/nyq8u2+f/AC8kiShKJp8up+9ckVZBuABDw/DZK4nm+ZrYP
tKpV6bWaTJwpDDJ00iiL9cRaNf8ujjc5Q+LrxPD9LlqJ3A4ROB5q6ZdzHhbsTvO6
LazQgBBPnSr/lws4v3O3mLy1DahHfD8WGbS037OzI8d9jl4HFWFoXzmhUV3NcVRG
mit2WF8s4o0nXw4MJnHr1VBjSmIXvc9x6R4Odg0n1SLYRjSz8nlsioP0FwzE1yW3
M9Ddj0/jJzqEYpbihUuC05jOM5x1eKb3BYXerA55EKCpPVBwGWMk1XigOTaKjH5h
q3e/8NLyMn4qlhSsOxPaEOJLGnXiDA/y+/+QtqGTE9p7UvUMa5PYPZH/LNucJw72
Chfvi74Tj2R3H7j6wYo2//SSH9f3L1/Lb/qUAuoFR4MDXn6RPUqgQb/Jork9vu/z
HTTnCWWLIu54XpUJkEDHYXHEJZYJ5W6ergqcmgC72XyGbCuIBktoS1xdL36wLqVS
wqqWI88sQSl30D27DYhuhGPx6gm6A8GbmkXkjcP6uYnFiPQNxPXo+6FdlJCjDYD3
H+uij2CRnUIAbN/1RykNYLEKcZaRQ9KhUfBNgfET3I7WvASLNaPMgibfsOM46V5G
jphu6W0jE50BHORl4PWG7KLWlHMDQY4uNJY9CoaENXn5TCAxtaRee7PYtmCThfJB
laGwOTiRbmdUWS+83kKO4iRKU7+unY3Yh+cmNCfN2oPXom8X1jS1EaCFE0wKaUHg
Mlbrp5vmbJOR+pdWTk4bUdK1VqEHWXfWOPLZMDi7++IR+7ChTBahGHvFVr0Sxi9U
jRHZspwftiYLiMu2WmnDcu43ZdKnPDmY0POTlf0SXwef3mql1AuxxotUwOenJAIo
YjgT1zIMGLcOTfbye3hiCQfNMBfp5bx8+vI3iQ56FV7IzIZe5blG3Wli6ZcMdhIX
98XJQRWoMM3F/Tsr+epo/ElbcfR/yg72qteVdNwfSinPOkexmF2TByyOkbDLYZPB
5nrcXILt6yn8d0TXi814415WHemYXLP+hPwODPxR5M1l3ACE3Vy6p+rAaCyQE5fF
Ez7YKzwjpHjWjfX4nkIIPPOBT1gw9CCAYEqRyRJvz53DC2SkaCPo/mEEgkEojIiN
o+ZNcO56rtbve7O7IJ6N+e5zuFaDmv9amvlEpMO1MietYqwBPvdlJgK7j76PgoY1
d59B8Dg3uRcmXmVE7It7LaEM16wV0YrxmGbQ6tcnTuyvdOeYhez9E08RoYb5MtB5
FAkh0jKBH4Nm7LkyVz15tDHtzCujV5FXkPxV2BZ4+qYSRwi2QEyBfR89uC+fheck
kFUMITSmll+nI25bAXk0OcIfINgOV0cSyfLCyb2KZf2mrvVFQQqwAvB76/TQuJph
ssE8x5sOO8EvNrpinhbvLl2bc0D5nvwgwfsk6nKdAYxq7++5vPUjTNC1DJXs7v1l
ivxcAYa+8S3vkkuP6cql0Ddi25RXcaeZ0rDvMCzL9lSLQ6CT2xMNiIgq5giO/IgA
a+AvvI6GWH7zCEGTMXd12+zozS7YN11bWHWkf91OL5aX9VvBKQGgovcmC7qEZvir
eFz081s+C0h0xa567/lGuyRzoOi9QZbZYOOw2+bv51t2Ea7zpHJdYliNMy5JH6f0
L/EhXjrQf0yT3OwnUwHvEzCtY5OSvlC+/ff0RZUeEmowBJPh52V/b2oTjECN2y6k
7RSCykm4euTMaHcjjuR+VkIvXOAs+mX72VCmsZ+TuxUrd8kRVVQYX3jjCV4sn47f
nC20Jr2qArhEI3JG5HtDtR6eXqJS2NJFIi6p1/PIRCzaQaKwCchVtvbEKsHDFc7w
264F3/gKko3YSgISYRRYE1sVeUbXCwgz4lFGpKNXHZM7sDBocOOXu2Xb8w30AmPM
/sF6Qf2lLDbV2f0h0ureHUaeCwuqbCS4KWthh5AEuD+xl/dn3k6B66KURX7eW3gH
GZwc+QAdrYe9vo304jbj8WmN7brbqS1bdoQrSOn6lK3XXg3q3e2jPG7dWNjBCaHB
MfdLr6iP79bFtwnhQESRhpGBW9wpP9RqnrPHZVH9qVieywUjprThakkhIseuQRvo
J660BYTdTGyL0Aaucsh1nWzeBwfMU9EAp1AwTnziaPhy8r1vf5OaTjbW6gooLMRk
ziojOWS8hFIx3mWC2kXkbq+YmSuw4r4Nu5csrM4ojHrBtIrnUbrnb3IKnJhNQacv
dnHMcvDe2jPNmcG7Y5RLAwVPtGsTAOLPXqipCr0lCnHAaBwjNm0fG/Z8dWJcumCK
MHpVtP19skU90+0E/tqwAKHSytcX6utkTlffirvJdXHztebt2ruUu/DjPq8HiX8q
bUL7XEwqETAyjmWIwMyzVqNCu5b0AFVqr3pYkVbjuQUUr9LcIi4KFREtzF1tulbe
1VlVTaFay5m9J3Ha4akTrmQ1PbhVZneRGmUFUz2XWs3w0qFmSI+rqR9x+aZhRlUy
kkDu2UVGi6s+upcpIQYc7/Fr67H1J3lRaCOZwZFDGtKKCPn/hINufvlSHEI+Cl0M
JUTvWltX79sBozWClj5F46lkGeczkDOx74Dsf90vmY1cnNSjNTubA4JX49oTw4CN
s5dRaKUVUWmRmSRpuhKjxsZL7azeXNUycMwdZGJS9rwflgM1Zxf4TlziiBheEXGX
Q7vy7tiT4gmN/nz46xI/sCCjQDDzDERtFlsUwD6toGX2Zh2GEtdZvRaMCFtm0k+3
ujluyc+k20VNLCgZPbWFJ0c33j2j01kQA7JF9+kUvZ/pJlQ4xOHNMsYSE/5ziPTW
NE6FD5SJBvQdwwFKmjhTOAs00RHOQaJGc0lBDf9aCPcXIYsea5urh9gcVtMUPwcp
6PUnPT+/N20W7SbX32f2C92QTvEsoufbxabsy1Ai+4vfbthLdr+dr1JwroPMt/Ek
cRngFbJTk/J6C+ABGhWqP/N1ha/BLNQTKSB6o1+NOhAv4tKceVMiMgUPljjDDO11
wtrfNedKFNKtq2MkQHaNKxnVP/6MswH5tOwy2e9eJFBD4UfPZ5pi5Ml0jDn8Gjkb
tw6p0xGWc3XdYqF2cr7j+YoBWvu+QLaWtTANXGQq57LgKxKR/xlbQNuPcPY9bptM
wf+65Shw6JWVYdeOYpx9vOIKybB509h/Eae2PnGTEcfz9deyy/XAsS0Vw2ICVKlx
VpjRY9i0x55zeTBaKZY1/rqB5AA+nHSWHPfNKa+tik3KwMXWxypOFQt5lsF8XcAb
ma/qQEMLjwt63jl9cszPex3SOFpwGO+iUxC886sHqpgjx1mpo3H/BBe3qXo4B2uW
ovlqaprXOBbImOvEhyCsevnhZj8P2W1Vuk+oTtVAcm5BszlT8RnrTImOIi/I3xoZ
sCe/R+cXBVkvOO0Hs4XavAJnK6yrvJICGEvs/eOG1m2f3IV0YeKz2nbtRB2Ho0nH
EudHzl+ivjQNKJAYWHpe0yNZ22BYNsiQEZGPUYrizQqtVHvXsuP8PbQyDb4qA3Hh
LxUQ/BHBaHISvAkLXoqvANnA4TNlgE5lvmuPie4PUSHoBPqyuRUB1HEECO5BDLw1
LBs4ckTvviiLXqFSCyxePsaXr6xAU3+mi1dEA3ZFjwPlG5aB/nnPVrtb0xYTeugy
djbVh+4mBN7FUccpqf+eprrH9QX26b2tFUYqy/Df0g1MabHj/empTPeWFcTa0ppo
NCZwo81NdfsaECufgJwcUxMQUwSUcg4Fn7yCCzxZxXRkW2Rbdmt9Za6O4UryQZjK
GBBIkf/bVk5wVQeIds0+ePQyfReQ4x/B3p4METMpDvFJakeKQeNFsv3h5ptcHUHD
KUQC+1DX/+l1aztTbqRZeTgYdTKqi3AYJfLQdSapsrlyD3Rji/FG7GD1Z6nF1x1i
P+p6fVcZclzg15x4tliQ4wMHOJ60iNWuEAviZKinKDOvhhlaY4wPzutp+yfo2E9N
Zwg3gBSUkNzX4MCQz5NzCJ7GpD9y7t+rcOc+1Ont96S5x7KdujXlEbgWBnHNPiPT
nDFepfoWM0oKOTuRliccK6RHO9Ts0RDcnDHFJe3TPGmwFk5iM4xviCDDVM8DRVsc
0DW1+uPi1VqBV1Z5tVnGfdSHdQ1EsFAwB+QrEP8wRs1PrGRQbYgwOpclMq3J2dUy
l0RgudyJOvza2gNriFlow4zSxQ+ZdXZCgfNLWK0v0ZbH/hvCHcZ54ZgLvdMf+5YJ
iFsj9E4+IXG61TKa75i5JxPqBNmbbRUa9dvSiMaG64tEk4OOTFuRWZE6wmuF4gFh
rRvGIMJ7ShQpBwzNIzsIpEWUxMTcsnVYGOnNH+t68XqhU+jX5cDlQfJ98qrBJjY5
BwfE8eqUX8wAiohRxqsKPdnNbJR5g+Fraz2Ba7sMe+1IHdlaaa3feaqkXHEt3hzz
C09x54PFbGG7aO6UQFjXpfybJwp8hGizbn+s7IJDWzPvH6Q8LO3Hr6x/6vis7jUp
yrffXqAf9Wn5m/OPTqNF28+ufbrwwnBxbK6+GoOXquVaHAzeI7DnQiZ/T+tMPNZy
hlWKhIvf/Sxwpdegq0SbHx+vzL5b0qXiWMqwvroV4fUFQ60i+NT4ONeAIgsLEodb
9stubbhRysAqD27oCzep3vl1zI13brvxXTlvBsm/1YmoWvkTpoH67Desh9J4NECZ
GO2qe5C9ltPvS4Z6grcdRDUmtQYwUInLbr/y2Mg/w1oYzxeJVlgRTozfwcLXhhIa
NU5tigRHxZdVa6ISabFul4LGeGGS4tCROdsyrWdSx3tA6vOKBYXUoJj8oHJIzX5v
bfFqTJJW0VQLJzXkjaUIBfTN15Pz8z1Q6RKffSAYTdv1sX0s5zVmkDvjQCUJVFVK
csoKFAOyYw46kvakfUu84AzozLbhnhQIzkZKfL/UAOVin3bWDea9CWMHQKg/K4gJ
fzbPFgQxfnHtwwJuFhPgbkSlr/4F/vYTw59yuJZzaWHvvnWqwcnsv6k+kks4gezP
DOeLZcfhvdpKD4W/Jo60lf31jOBwatOppn+ePKSEtIbJ6uj4WK3bzJo2wcPZ1cfQ
dk0V4+fccZZxWpzKGjrvwjGu81B98ciqYODnQpy+/vFDGBSyTtSVovYWBMQYst8d
+iLUrE7DB05IrKD3+FaE74PQE+G8SSYwtZBigr0eNZJnxyZ/XsEAIauh7wcgE6hK
Hj1MDRAmfVRVfNPb1iTt6eZWXN4Vp/sbmFVYOpWfRNIinGzhMAUKH2uk4fziIK1C
VxDm2VysGWFVV7xw5vZU41DU48DBp6+aKNIFRw84/4tfUnq+Sx6p0SysOaHXThJk
C5KdQ6Di8L8WuGaEXWowar59S5F3oe+2LANHP1DXQE6ifNTh1xu4sdB9WUZOWUrG
u3syY/mRjcd55SAdMpecON/c+RULQP/+n9NQtBjolTJwRLAqUiXftbXG7F6L68SP
q8EywmZy5iu0UAiBBBkacsUp6KrGBHBm0F2Cxtr4BbZTvxyz3su+rZWIRW+XtSA8
K5djhaX/vfeqLgNzZiZ5RUwidIvPhK6HvzhAv9ohroMCcutcoIz1sTYF08PR4EhJ
kh4gesPQm+hoDpsDFn2EDoW/cc8IsWONeN6TgGQPKKwwWnEeRdTdd+gAVY8K/iL3
VFEm7H03/HL61C8SQT+2lyIb6WhKocp1KVXeTmV4e81uukxFJ/slIbcBK9lJxfjI
fr5pcWZ7AP8rj9mPzmC9w7CxNCu2WKqh7IBHfK9CzPV5MB3OJV9Zi9GlXal6PmS6
K0Eb9PdN3mYp3tikGF5B3hQm9pAOzk6XQKLZPJg3thWTCzJ5YpVMqpj7SG8V+HD3
MElXdpbpvW8dNvZ1eznk//FfH/dC7qEbpZ5siU6T/jEdAAvfxZkfmYjc7IWElohH
ra+ohk/FcthrYiDyplXZimVNrLohGr69WC7o/v2Snd2ke9dR+U5ciGXFfTUVRq1L
K6bvmk/hpwa8dSSj8M7lAUy7cLxAC+fgyl6MbSMrihJvefUL0WMzGLYgmvhUY41G
Siqog4SfrVKQejFwaeyqWxd3S63ceHCzcFHYWfV5EDjUAQJC3ItniSVQNKceaCe8
ZgIPshSvBIelUfC391VhqH00q4bGI/bgXcd/nP9yoZtCB1mRnFhCYmkmN+FmGv4U
KYQN9fiiRdHpbwxTw+xlahPrxsEmEXkI5OyOXo8Brq1xRmR7BQBqRi2qSVr3vwqJ
hPjRUZ3QbEanHtUtJiBnGBmd1Tnml4+o7VZ4aTDUk0Rb48ppF9CAQpWvorIhXYEi
j9lov/OyrsrdGmzg8jEUZnWjlaM7ekxIWYUyfPCFUB60mPx3fOuoE6pw+tZ1lrE0
uiBl7ciafvxFGV2YDfB8JtXpKowps0DP8KEPKWlKyrUWBap2TjzP+xIoFitiZ9gx
HcdxMLyOop69OcALg3lIuyoDxd3mGGNkpRK/bJZFUQvNdjGPbDCtwEbB8Q4FN0F+
5q6KWeZSUBV5K8pxEAO2IAvLRV3hYf0VoK6sj+UgqrQxjDEA48JxPMN0XEtl6NSG
0vUb656EESuiLFKsHROzR96AzTN1VhncKzVkd6TJ4tOJ/K3SAyK1yLz79J9HV9Rx
7Cx+REKkkfClhgvaH19azT02FN9ni1P72ldxy2a92fM/m1vPVeApyKKjeWyAHwuE
yJ2u1CdTEmO1KuZfhQxQJn+XMLtWRWGU1fyLLjCabwx/ES9n0/Y6WR465BeWZ3z8
gfvA5804w+3ytCoNCYIj3ooTBqNe/BbcQVECQMuUoqXIKRnuQuF7OZhYSQHAyNGP
zIGp5kLBxrGYN1s0W8KFPYvZZeD1EXKoUCF7bPVb/KTOMk2+sXH5+fDSrmjXifc0
zadR2hJ9wl0TENSKVHpZWMEGW8boy0ssRGZZipJNvMTV8fIyO/0VaYjjFhHqOqSm
J0/pjfH7lMR2cb/jHCp4xU3b2d+vmKtM2tvbCTuqjifpTMDfPMPYMg8YagTSSiEG
VBaBAmh932g/W97fQfAMfKn950TXBa3XS91I2QaJ7GFvXK+WuBkuinBMRBB0v0+5
m0OIHcZB9cWmJ3AQ6rdRkzOjjSjuDEwyXxkV/hIggsm8hND7iO7rOIqeiYNxQt3m
8daFdrzRzCpEHiGwBOYmB2Mhhvn7I1zh5ZvkZGDcoNpGtJZ7VmVBLa3gBXd838L5
1PUN0prJXEH57pI/ZUMM8v0GSBI4zJBNCtzNSSWy2+kGpk2v6UapemfI/s+sPc+n
skxhNe32vTOnQATdUa3Pbs0vDIKoMZTfy4oBDujkc8gY5PSxYYVlCuc53rLJxIkp
h6ZV80jYDkxj5owlfhTMIGKLniRUaiUVg6FHHvP+heRHfzmuTZidJbcIjdskOLaU
Lzx/38waXn69Aj7hhu56v+e0KzHu6XDU7Z+MFN77VF2g/IDmCW93XQaisOVT8Xau
hgWoi1yktU8dOhgjZO+um0NQ5YG4avqEv3e6Tp6x0fAFaSfwPxELUHDFOa4bL0WI
a3fLrPTRfDNkXum9AJpEmMITriUXTQDAwk7CCiXy9jakPWLi1eFp1uaxqTgjGf+d
4nCdOrEkQa6OZ+t/bmhYODkRq3qVv6pAaH0Kl3wkSTJ/ZDlncV7cfrKVUckCd/E3
/ZOJVeyqxOqI3puPR5zfQeKwnxJFRblPKVqz7hhe1P3RVqILE6kpkZ1OzsVb33aO
pcPrngmdr6IXvJ/LChCsbr0apUMJ5sjMEwoe5aTAZymmii9W/UneQkQUF4wSerFQ
ykA4bLhuesfLcKhk0rvBfbYDwZIeKEaN2iFKzfJpP9jk9gDykqDn1mJDsZd03Y8V
tOWahC6cF+oFqP44yAvgJsKc4DaT5BGHbqd1gpSj8Yvwl3gng0DuBgiF9ghBD2iY
y3PIlgYn+GhxjgAccV7yKrHljL3bY2smWJywkHDDKa9PUj25YIDvsjxLmDy1EvnP
GnZUmpLcQTckoALfLTVOMTOhBMnN/8Vve6Soey1SphLysdQQ4da3At9wcR72jg26
h1agaqpH1ZtzLi+DDPcPJfPq9NtzMbX/hd5/mPP19e2Xjmp7NDxZ/i3mYjPjeuFS
lACfGb3PAT89wmn+Wbvt2zqc0gjmmj+JLrIE9DAvk0BHWX275lccXGPGzMNcHUPr
etkeZMmGN7fw2h/NeYon+sPESg6PPElOG/n4A4TFtyVIeyTfcoL7XZHZPs6cIyWr
ZwCu8jevvDEWzEjSIKPWX57F2u6Avbc/C1h49ewBVM9NUM1Bt6WW/cku0nWwQxwe
blI8s/BuBlxpVZjkqgEQvk3AeVyxz5CD/jHGmA5tuxiVOYoSYTilkLDb8xxnGJ3/
Sr6lMoPXWJV/RWdS9bbXWwJENWbT1GS3S2gWDue93Zmw38ssJ7BmXuAAtI+HdE+m
4s7s6Lfuown+6eXpbnhGMbW4wtCNPb0WLnKvQup060W7R5QqfD96ZEJhnZ1Rh/gn
V7XJZYfT4S6fngvw1r+6milKHynHkdzSd+x6nVtmk/AS0r7dlbYKei4NgNX7l1s7
RX/kFbF4Og8D7o+J8ZozwFAWqTWtMsoqp3aWKbbzxhKlmu5EyV9K83EBWQQeM8uW
EOHWgWSppPmrfTu1HF2MQRKmYLnbOHU0z8a//Nx4QYbZgm872blgodIV+FfMCeMr
zfjPk/4pk8OTJHs/8RYptT6pmVawrM79aIqPgykxokxykJyr2ZBK65QLXJig07SD
29Ur1sRm655T8cniDjfNyyw2do40TRWJc9HApqJp3uB2/433zM8nU/URR/qqpM8I
nfLNUijhSEqWdXJWiIpAY143l+2ol5AhGiECXphWzuKxtsTSz3BMmOkH6F3RRUPS
dIToJXh1rbb4WtOI9wrDhhTXkcFX+Hh4xydBWD10lJlV4vgKGan6FsM4cjTpIzJI
86C6ThzvZ0rLFCUVeYJKeosM39JNs0htHeTM0frG7Tjnvt619Z/SyBDPkhJVwAF5
ccvoI7EClGqlumaQa/wKrhKpTtlag7PruAYdcfZ4iomu/bZ70bru3bTjz+OLTObX
A1dbQZWisF0bo6JRCQK/GPS2WblB1/v15HC6pEETSDiJQMeZs0JRYuBLC+HF5kwE
yPVlYaadlHS51PJGRV87NnCHSCIZnVPR34jSHAQI01ci803geTVpCnVlsxqmBWqJ
zh71jYvJpm2Jn0JxAuEARSBzrkCIjthd5uZGYrdthHfo0L2qEbe/DTAgAKdDEWW+
hvQ82rakg9goMOFQPgy9Pk4VJLi+IsIbqi/X6rhfzghHUOJ0xECDJkL9MoebQsbU
y5le/FVykic1xCO8z09047MSLUsuT4TUvefkt43E5mmb7AI4kwuXezyC4H+2jPBo
DcgAPxsE988HcHYBRuhl+bTx4avMCMj7tyELxrPFVhYfOsfa9oSBxAhvs558U7+1
I/ll030s2BUkwIfe1CVv/3DQdUFEtQ8WqSNS2YdwdakTHsnAFQKaIHDWs/als8OB
jUuNJYXGuIahlxV/IPNEsYoq+vk2D2E1NfiCfmzoHDmJOmO4SB3U9GzEtNcTSWS/
kHXQLrQNHDAm1WrjPIqR8e27A3dFr/Gfz/2WqEauxpsqbgMSKm07+m+MgyzOOvtz
grq7w8t/Tsd54Sr1DiEM4iwSTzrwJ2GXf1rMVIFSk7Jx17ZolHwELNDn/SX+RwrB
obOJGJX1g386AVRXAo8HeHr99LIeIHJFz46II0gAMvImfb2MoZVhpKAwKgKjqMMZ
WOXhiJoBHo6lB7OFoUrdFniiEQ1k7gjeSK35087M9yjZDV0z6DjUSgRvpgOR9pei
gBc4LVcQorYQirNuczhZBCGWBVXx/jbOIz94/EZ4ky8sBPgqxKJsi/AHijhs562w
dyg/N6Xgd/kJyM7DzNxN539ANIuOFo3nGvOh3CzuaUOO+knOmAe7cyrmpCFTuIk9
2YROrvhwU4gihys4syFTILKO4fi5EW67yWogxxFPo7fFNjKCU31DCYCCK+S0Io5P
iD0xVuGcGzHhKAMpY9/+ty8oSvCtstvc+RVaA6ifvNPf30brznyHP0/5ZUd2/fnq
+Iv2MVbUJlTZro277yn/L0H9Ba9TlemCe2W4s7sUIfcSBXzlAqllHoU5TIBQScLW
k0R6tjkHfxA7vGuxBmGq1ErHufZ5YWKg+Ir3P6NMrsOApZwhXuinAjiUB62VzlOm
5TBqk8ihST+3tIi7srjechgU8i8PJtut1bDrhPhUQA8brLHMh5vVObPri176XEO/
DfzwOYeYjILgbsjZgKB1IZWE0pVUlsB5OHQQPkd2QiqGVG5FhnAuKpOMZeN4ngkp
oivO1xCsai4TWVKlcvdHaz+MzVaF0vOwrGzsSjANzRFtO7EoDNGv7WAmUIZ7R2Y9
RMU7xCSS41VEerZTm5GUnHFwLe15Rhu70vrofBC1MH2iuHTWHcmzdD5UQA/rxo23
9C9fxzDzl10yGXezCOuIllnQK2bXQqzJC8oShmyDbFJ+dx+KOGEpbKBHAPfHKYlv
tNal3LS6mpj9b1zfkMTMqRxr6gue4bxvtWRXeuYQwGsWqd89oac+oEvrPpMshBPz
FSvpky//l50gh2Th4eOOJ4bM3Mb0CxclYhg2uJuSlmuOf0sgunMN69XrqfdH8k9f
vv+5QCD0JaARIRLwO6QDjiZd5+6Dj7LKjT1CEPtCqlauyeydudmplziOD6jBVQGT
xeAmqAKPovrkwRNc4CP1sw+5j5GZbvRgXN7stBmjIzKxRq5VWi76ldKmm0y6Gbmn
TV6glqYeuclvMuff15XQ90bx0GH1s09pxPj/0t69B1Xc6RfVXK26p4NLy/RxnF5F
dukGEifxAuGVH2yl5Mev0sq3CXcFKCswIwxHrIolZtQf2s3VmvSbDifJmi8ASz/T
4KcCzoTzh07P5sd9n9WV4q4isDTl67HGzPslqHW0LRWjrdoSZ1lbcVcpRFFvg2bw
Y1MJCtUj+PJo4+fUoV26VbAlHqykZaFJnpBH9dgmPdlU0pIjgJck+tRt8N2mEghD
IeBTbSfWwy2B9/IzN82PofUPp+utNZmNbTLyeQaUuU45VRWs+TjdwqIeM3GE6Mqa
d832HCro00V/gfizwZpg+KB9kAK5k6Ga7sybrw2G1LmWIqSxlzVwXa47c/e32AuK
0o1z6+NfWuVJPsU0rrTtAcBW3TF/kLLQnxsQkqjztUgW3kcuv8Z1IgRVUlVclNIi
2MGI2FP1XEOEzWGYE5hgT0MjMcplYHEO+W/spje+8b/qofcwu0efWEf2+x4FH3N4
+CNQsGVkXvrtXexEH+ywEqmt6uPXMaQt7qAU3O26YfDx4jX4M1DgMJhhaixdNN0I
zGqHvDvEF1JJk6NYzQdYDjJ1nBX8TTXL9VImTfGELNJHBbuX4C3HwXS392K1dr/3
ikTTDIMpFoyyMxW7su1anY/0FsfFmScHupMOtOAjqcvlga5MteXcemhM5vw8e/k9
OMGWkl24WAHSxUMMWw+anyc5iUXYH4KdW9Zgl3E8Glt2UcO/yOKLRUewervzDQbW
f62hoFcaA3pIxMle77o6LWOV9Jky4humjRTjZjHuTSrXhY8Vmtnmm6rDkLUbrYXl
bwWE9gyGdXrWnjTMjt3gBPuBWB45v5D07QYEzx2vNAQd8xzSr82lZnyxKUSStyU+
Wo53/tFh2m0GMeHjIEOgamHrq8yl6vG2QYiH4nMH4NR9QeyTS3RBX8A2XXDSagrs
aLr/FdjzfIUCkdH5AWiCVnK1eToECmslbOeTS5u0WCtn3dKOp6ldtjekaHwvhcPH
+jH1GEdS9Ox387eZXCuj71zQA8mGbd4JMpSNaEpAEgCcuyrJtcN913Ul4pSAWGHP
hBx0Msg2305EDS7t5TeZbsbQmCj3pUhrsyf+VFJVNROBV0httrLoUOoG8UrCyg0A
iSyOKQC7B60WqER66ts43Z8zFX0AoYfaSQt4t7nYlgRzmiTHNe5pQWycZgNGpG8w
ZbGMM1gyZ2v8Hpu1AnH/sRAQA8io3ShDyAFPZY0ppjUkJjwe9KtNBG/GKJyOGjD7
cwrZm3zCQDz9OQdUatIbaQAbCm5hmnZ8tazbm/KKUQQf041xqZFEG8eNmVC1PRY8
vs9f0nrgadwuPZ1ZQWQjpKRLQ07Yg3y6OYdeqtHBFpC+Pxuw1kH9cSbDipyhh0oi
m0fR8dvRKoWUKd6o2l7nrSlTwuudLizv2X/0eZpBns/a/fFoWxCh+jZrGtp33Ud9
uHtugHtyf/lWdV3Gs+X3kJDblZMO7WHCuZX+BLhcH+ba7F+0Z6UrSZe8ykVZbSU5
kzZQYsbxgNtZ/12HiomW9qbB+cSMLncJW5if0nbsGDMxozw6BvDNiyN8EZCnrs4k
wWPrgQJEaJBFJRXWsns7iVbXfHt4KtxOD/zoOuvGRjT2DP6yr+IZzzhw52EQPvKW
DbvUVsJnOW9iieglL8IMoU6hh/6/1PHfjO/Nld0xkdSk8xl45ZtCTMSX789gOaFT
ZcrNJtl50jFRi7mm9+pUXyMYFLOieG/7d1+Y3sYStNBpOkg0zWi26r49eXzG2gs+
Tchelw1OJ5b6Je6eUyq6ippT0I+lQp5MxxmrW49NQz2hkEGegJKyczYq+b+HBqBL
rMm4yXN6P0f/8Q6U2PnpoiWI0Z5oROuJAG4gEn+OjYyYjrdpmg1VI+11TVf8eMV4
r4T6pVMeWnpmKT0mqUcuQGuvnq38dyA6aNU47XRrTrTXplEp9vO2ZVchCCh/Bj1W
GLsqEy36Hsel38B/+3gcU1BOVXap9KeYuGOsDxrykz/yyo/+9ZJBbvBdGiY78n0c
Z2q9SatR9FjuyCaXrO+d4hYHRrqVVcWYsMXaENSF4AAaM3pZjDIvmPRMLRcoB+F7
3v84fHazBgYB/IH94jol6+KJFh6TjKOJhbOy1XCWUa3y5Ku9I9FN3Kob+7B0hCGO
5qi8/8lOB7sAPffh5NwoddKtb91aU1qKvYICi9elzT4eERPQiFX8gARoOPA47aT0
7Y5GIVc31iz71392MDjEYCG1wOvuzIRAppDXsGxysSzmRkrmCOah2dZq2vMqprlP
ilQw06cJDXFBO8WC23egC59A0ubuf9eInai8IKJ3UHfPjBzue494/uT/Eh5Hlwm7
aypnaudbQah67ZH25+S6ABoYuT1ooFHOEtJhd2W+2nMWjWJg18PMZo1s1DvJ/a0D
6v3pz1yDuxto4bZ+xlxAD5Cqg8pIXp78x3YBxoskNEWHrtlS+uhOHIFpikdpNU5d
TfBVM0YcAZ0VdBNZ3rphk+CvC867qrJb2cNkeb22XusazhZlB+XSmxGUNlFUwbTD
9VdagCJlXc1PlunyjbGBjRv+0cqio0nFIAP42XmHQYFsX49/orOtZP9j2xQKu9qs
92oKD4vGG5TDvTgzeU/vgsf14hqImV6U9j4lFm3Z36HpKDlNpgesfjGqW5Q0JnvJ
FFxJtsFXNlyfXypzemQi8TwkfBUXNkkZ/AUFUiBi0RDW1ChozVOiSwvv/56o8DaI
DgE3x43TcMgkZ4imtagl7YuyKE4+lY7Ludr8OZqofmSlhHXT/2Gw3ICtJSSqRlzT
bLr+x5O0riiLJ7T1Pop/45+IzP/7j5xN/iKIBkmI98AQaF/ooVWxQD4d83WSd+ml
CNasNrQVagEg+D4B4SB+qfvyF0k3uXQdWe0lwNbkSSMbmvZJg3Hiv+EQ3WgyS4SL
t35JdFhe0H+PXXaBOvauwigWm3/7Zj/xT3PyDFL7M81qrwfmDqWbmSt1d9xXocRC
Cv3Q3FvWPcC0FeMovoGNcg==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RZWvMefnYvAtK4riu4PPYW73xUtMLUVBXXVbZlsdg5Op9rypeLR3AwXbkn9qjus4
dmQ7k49wYWaff6Iotnv56mbOSwqLGHcIGaXUN+t6ZQ1qKRD9zKuUpofwb/uRGplu
sfEFzvclsPsJgfCEXQBlZaWtqY+IoloVZhNsiSV1SW3Ajb1/5YRzTLqW0Q7wZ5Ak
6ZpmOMu68GE273/zYDf2k8D2yZY3e8wfdqIotqR4ANNR6OYV0gC1Pz3pY54FHlDj
am2kaXz5TIy6MTdw/gJXBiyQZFJqIlxmB35UkJcTq2II0E+zP3/TS+vV2JG7po2A
xiQgiTk5ZE51i4ydaezExw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8688 )
`pragma protect data_block
6KW2H+IdpFeX2gkVFJEE97Hi0R2jLkWIwiQM5BUQhXMLyRCL+9ub9bYzBuD1k29c
XYD2HcgTVgwtJMjRgxnJXqzrNhFGJD9VHWH8BiMef8wDSKpkeau4vZ48qOvgq7im
ZTn7fvt/beXmbx1SNnJ/W9u5Ftadb7SmS275X2d9CBTSPTzmaI47C0RfcGS713q9
FT/Uff1GeWCLz04UE1dQkWg+lfM+NXpnWZvIoCNWSQZ8GGfQP4RgRbEmtCf5w/9G
s0UjBjg5Iro4rwwd94G2LFpABZqDzjaiZ7Km7d0fFP714gE+4Wf0OZZCPLoKzVPp
nOqPyAIRKjV9mw1AWc28C4vEBD2QIkPJ69mcjMnCzVkUVOQcJJ7IdzsjiRkjrC9i
+uFraH5eMeuWFKbCAKJuCbCyctk38wbUiuWmXuJP0JJx+z6Gx31w7fqQYLGtxQ0r
TmN3W9sQmuwc1FMMUq5OqFKjH6L+9PMdD5S1Bl/lL/I9RBPCo3qHJglrebF6lNmX
G5u7CpZyGT3SQpQCgALkIyvxbNlkklL/sweISRvlTu5inXk65V3YKBJXEascuAKj
/1Ik9BSmutdYoZ7NRPaeWPInjyUJiZfqVxhQqgqtdKt63O982FQx++v6LsF6c5wp
kvOgUj3SRJ3pOohvs2ZbhGEXUKFxpDpmh0VvdOG+ZXoW81Ep6hlQ0G/RJKnkmyr2
mwaBW3xat9YZdYpkW8G0QhMzjlUqtsKlP4BrfhEx4jpunu92psbvE0LmRmU5gZog
Ou27S/w5MOwfq8LuLo85yGg3rwc2jHpOeiAkO61iEHvI2Uio3hbH4rbcUunZudii
Pv2HpbuxdM2A3tYoO6vu5dLj9hBkMoHpJ+WERX7aBRD5srtT9yKi21eN+dMD0clJ
wdlAyi0p4ojwhCmyukvzymj5To5OGdukNXmJVmbwWDtjpPa1BwKVJf9xePZt2uWx
XP4d/iQoORcXbKIWMH9m6/MItLEnLhIUD4moiJpDbOp/9pG5303jwo5x3bzrf8UM
0CM/635Ont0t0uwn/fAXG4+0E/xTMyvqgns7b+z5tt/RN4lLrpqyT6596KRJnql1
dXIamugKKlTJb5TR/Tm+JIdfkDAEHT7lM0s1uQUtEWDPElMvPcjDfBKyYbVGTpr4
04w6eWz4ySuWTsDL9v/aTr9R7kJDmsGrBjB8g0eXvHluljjbQkw2OZdPtwHgnAjf
bCk/I2txde7XxMSDErFW7i0/y93OnCFMeKHbTkCafn+d5g+TQpGXAmDQgZ6GM0NM
RGOFA5JilxO/vr9u4IgljI47Xbi51rJSEe0B48bqWmPs7s6g3Z8SauVH9+6/15aT
7cK1drTrlImlVuoGz6CjNJy+iiBR/cBNBQc08sSpCl/ztqavJIN+JFW29sYPla7o
UlMQwndCmXWqkjfUgmcMMW6FXrVj+PDMpPGVOfFGbBrAO9YW9GQLaT3d+ZzIMQ6q
ISbNkfZAXl+RhH9078yZJKgkULM+mxuk46W4CRKto10koioks6RjBmW15WixUbUa
3gmPcwJQ1WUDUAGcHJL1ws45c/5PwnsxWpO7C9LSvej7Ul1TxOILUJJZwwe5EZ6f
1oISllJs5kDuzYIIxSen6hOc8LnPEmOJKoa32g9gagI50yVGUKb4ik5JdoqUp+/7
M8Bju3AztDs+lXOhKBkFBjo9edzTwpzE3qKMVYKh6S3xqmLbezhqQMU7lnjnqeyo
MNu9EPueP+3/KpWHcexMjU1QzpzmidRcF2yh3xTpbRbCF19ItjYl49pEdXax+Tjo
QmSD5tWusxtpeiOdbRftdSSETfpVZNB437GK5YJIGX0ljGvShLvGlj40ROczBxSj
Dtk3aRWlYnfqfZhdd8ST5weFLDmvw1XJOaHwWPxYsCfrQjsgmOf7APyIYnYI/nu4
6IltonDq9tNa1gr3nidTCAjI3AS13eN1gDX8AZiZ6n8y2b2Ob1qGQnAUBLAYD8Yj
b2zkhX5f4inXiyejDljUTTdDG5Ma1o5L33UgJyUwwPkshomCpDqMNsQlDrOcfAHq
8czy490txZZpnS9KD3N654W+OtDkGayF4AlSy6eKGrZXDwWoqAAXnuZjJBuZM+R7
+zk4Ozv1jquCpMwvbWy3NZHnBBwmsb9Fg8qYxn2/vahctxS9Hrx2HF/dzjDlB291
87kcTejGZ79+g8wl4dXMMyK3/Hu1YhgAkXlBLVyzP6CuZ7jziVAPDvcRpgI+vvVQ
L+PTqKIkZ92IvCcG1jabyQVUWKWJ2M5h5bLO/AdmUvBURvGIPnebFxaamDeAb6Xw
7EOaV2Edpffzs3RjYGiakN6LBdIVwsWqSqgoKV9xGuF9cG5ooPjP+CY00xdRpyFo
toPsymJkvvJflyFlzmCsKd3DDi7GwC997uM6qzPqqNkRAnZgj6IFO+aMUc7a5Gyq
8m7+Xdus3sT+3qMz9HYEZnZdnSg0bayS5nsjZUtUbSqSnUTewESZAdGNw/BQHI17
dM4HnR5HmEBJXvMoSJRWU3hfdrpC1zFumJVPYEvftvAoWheDwedsuEocErMHWZHY
C3287dWocfJeSR6dOdHMtsqRLyDm8f433KN544gVfOGXwfsc/C2Txiq3Ef1Aud5t
JCdvSHFqgsyDQM5SKdnaWW/1YAcejdBruf3Occ9DKwac/cAyTgwjHeAMsbS4knzi
oABsMBX2kJq//Fdla2+lb/v8Jl4rFrelPvfKQoQPABQLLCFdcWKZG2iLXGN/qUHT
nw3pCPVblFfBZQ3adKLBncE/EBpH8fo6lsIbEv5TFBPGZxjb+7ATdkNcLwfN6sJT
IT1zYViashgnwpimOYhe46xIvEnmYmo9QDRq/40vOpy+I+Tgx4397/BwGMccbrj7
Jd8aJdDwBs/z57HzN1wigXp4owruBIibJ++KaWY3SDEsQDvAIZfTJVA4a4EWnoak
AnsLXd4m63oZ1kfdLEiJGnToljqJfs1Nc5EmTenBoOGymbCZpEMQAL7ZaCDSMgoS
kROY7NdB8RTrZ9utQZPZdwQ/8wSmJCJCYofsRStw1NFwh/9HPCd7Zotr7lazl/tz
9OIPsz6/4q/LRQz9p6o17yPobyOEVwFWRIEaj3K5yTHiRcIsfyOUyZ1JXGHg8Fb2
UX7v7Ydn61Urz8J3LqwRKlA/wIjaEHTF5DJt1pRxErNYX3LFCE2ll8sU/l5n+wBA
IponjLTwVCjQ+xe2oMBIJuRTMS4vHm4Hdycw7PrATMAOPzlkhLTmOrAhRioVEGaM
wAOWOdBwsE98zR+RYsKpauZcGVTDLqEygTyRk1UEWMuy1Jcw+wAu73H7M6f/AQk2
aHsasvCdnI4Fyvr+JWzk1MB+R6fsaWQ5bypnDWc5cJPdk9b9rje9HSFgUdtSocxA
HPh9HlF2KI/RBjMrKNqnZLAWi4YQcoOxuYzzx6k7SNi+UcjGM2jtXpBO9ysyh7aM
vFXtieSpW2HkQ3GhaMGikjL4dqyP5WojWCKFkckL0zWueaimIzSgDU5DRr8d8z0c
e8OnR14tDGzIRL5m2N9TlfiXxeYxEv6srtjYLFmC1RPs7ktm8pV+6kG4jFuqlU4G
RVPaK6IvV6MwHyoFKg8nSEVuAZi18hfs/2z41r3dXWajhPb2eIYB4mz5MZHyuC8n
FQZZtq+yNjBCY3G5T7Ya3xDuxXK6wPY1Qbe8y5ycHekRwxOf+aXiAJtVQPDOZS15
jheJ87WHbpDr+3fVdEhLSAGI8VeeYeoU7WZZkO8YcPJiOgYf1tk4sU7p8HQBiRFf
cy4DsZvSoj8vah+lUzISOvReWbbKvx/gDcSfonJjP6ztTPalqATbKbLhfsM3LUBq
sMrHr/H4o9qx37gObE7xgZyAAplRUa49cc2tyDrnfYZg37eicRPjND+RZXP2rpdb
zzlnunYjWJuFl3HLNxGsRIH4TR0XcajwgZhWxNCa1fenaM2xKTY2d0uPENaNkbp/
u835btKce5e4VQgdVkWUuFD4Mc3f2zAQ+eFsCpn3xPYG9245K3+73J2gvzRBh1bk
WnwAMTP9AsF7rl3CQfMgXvvPktuC8qJI5yVldYvyB7Qs1kwuYdSbXUVaL0l6memw
bBEmHGR0CowS7T1bvseog9x/xb52vHaudahOgeDdoyeFQCEGYLP1dcnp48wPgt7Z
LDKd3srSIA14PKwbDbKVJC16dv5EVT74cCbHnkqAtwa2jScTY7MeJc+Qx4sYwNn+
tglMMOFsu4WVDUph/mlDm6Ybsr8Kansb/mgjv6JNaw8RQmfLb3cLSfOil3c0B0lJ
Uh9EEOHYbxkZPFoatLFWckopUYEdZBbgkzr3si4PoJn5qY7Rkckze9cpHRsZW4mj
XlYKUHQBrybp5TgA1Ux/cT4D0m4ZuSWIX+ePCkHXl5uUjPU4NqxQJTZhztVExmrK
O3huBjYjL7uHbscNRDwa96tTry8P/EQ/avcozqTMtbColbxT4ALxXPFHVcEO72bx
Wm+jpdgSaN1ElSfmN/9J102w04FpptfI8Ty3kW1QJQX5k1XSkF4dtQsffQf4m7Mr
qN3RiwvHpzbVYRUPMfMPc8VD+HB933RV4Jdn1Ae0YiQplRcuNDdQHeh/GE6awOoO
FMSCOS/SVWuaTEYKTFETZeUQBIK8kpsBIxwfCQN9TfCm97HJdntw10EDV7fu3JeJ
ljSHGnxYsDATlRa5eQrLLr5Yw1jiN7sG7LG9VuwSAlEuyppiKj4iU5rMA1d4cnAA
y6T5eiCkd8duNr6DofTiMntYP2po0vdtpsGeP3cfVsgV1yW0sz2LDMm4dUCsm6Ny
udPE10vjpuzWjLKGM19dgjTglReD0qKXk29ijGWFaCHjtEv71ihHdj4+7wXsEyHM
Jv5ePVIAlOsL1k+uFxO3h3vAEVDK1iRZWPgwj2ZBuheZX8/M0/Et3FtL8yeEb/vB
QUWegLy4Pb512EQ9R4GXcJOUpw8KYO3eUB1kFshcYWaoPPER6R090A3/gLWB0PW3
O20spiJsFwuM7E1jwoo15L3wPFtHUroEcRNJJV71evWxEZcDeXQljMcr2To7j6YE
P4RRFfiCmwVTpaqE7+HsP71dO6qx6ViRFAY7YNscO6NV7z8BU5TohU9V0n+trDOB
KgHL/Gvxk90sz4bJkrr22w3GMAkWBrAif6ngJeNRNR70fI/GU7gzUVbbCqSRS9/6
jeRL3vU6ZgthQ2ZREJa6rs2eyYK19Ra+1686OJwOqCJdPo3gRTJ+6N3kMfV7FaZu
MiyddjOZp5EvOLuFZVvp80REp8fszIP3FOAWULSBI7KUojZK56nhvHD8YQgGLit/
zmMNCE4ujQ5QRGzr0bLRXehtwpQ5IInBJYDoGRVrYf+stUih14TPDu0yamqKlviE
LvGaE1GAqvRFSY3yjs+bvGNf+POqYODmCKTP6K2fkjeEHTOIfhA/PTgveXTuWZeD
qgayR7nkuJpePCdyeoq0jYlU2x+DG7WVZzL3z0KThIeOYA7f6+wsPUk5RF0QkHPg
U22tScCmev6qAAfftE8qhZxmj0KFQYH7XofKogEEeMZcuUxI5pxVSP60kfOByX4n
bsKQJuNChjcBk56bxwKP9WHYqeQM2i2F2E99+4MGAN4Y4WY73KLakT7tYadO4lhj
XLn9a6+wbRSYaMwN33PFWbTZ1YN/nYJcCVWfs70hEzkHwQOxSaiuqhAQpYdkf9DP
lV3Ye8CXz5Z1XAS2O9eKeD7/KeMdMtApiSA/1RYp6/FxiZ9xTOGZjLPP2cGrrUti
KY1QhNIjmqctemKheEt52iyguHf8kVpnpuQ5V+prr26nyAZO1ncaGLvqW6xWZu7x
S09Y2uYd00Oy4hC/fIyynZJg7kzJu6j6KeXT88ummN1fohkEMBJx0/KW/9AqJG2J
hE54AT7pN1dl7VUShW2XCJuGzkVS0EmIQZW+Y7etpJq688I9Wt1RknY2YGloGzVo
VGBS6vMdqOMJuYUShCAMDvo4fnnomROj3GkSuuMJemUQNPh/b61gOnplhDlJsGhV
L0c5iergG951K6UWRtXYjtxrjjRMpdNZRw9oJd4VHmiJ9ZLNKdZ3PX8Z0Qq2Ks+Y
aNmSzR7TtjtCc6tD9KY15MEOAX7avTtFLy3dpJ74Yrbzf+GyA0jLyKPe4nNKBnTx
fDv9g22hdqicKV/2Qs7t4X/iOK0oJYKDNJ9gamLUX3qLXBwti1ogj9OY7uQnDnn3
BfBlIezeFu+x005B4C5WrXy5fKUTbPHTRStPHhCR0Bpy7nj7wCeV/JLv4n7X8jYD
bZr+/nLCzq5SaikxBXEVKpkDB5YPI8d16QyDQxySy+Ib++WVTze5RM1kDkfNKEhH
rAUM2NRyq8x+L79sxysNiT4ngzRu6cZUXfZvsKcs+5UwQP1k3iuwP6DClERaolm4
2YMXhV6zd1KqNpjDzCoHLegEUC0HjaLBGIPg2BEhIO7dWk358qIwaHfXAYqyFwrR
cnc/7woiQL+8M9peyu8cIlh5zdpLg0PPwx8iU1I2/nhm8ArG5ctAqpG9H5wZlcap
OWWWcRLtQFStibaaxZNF49mYGsbNoa8o3eb75YAAa8FJzwKHaMN8P5ObrXOJ6XtA
XWqfeaWmgzPAMCU9TkDq88AVoqnAItmSBucXJjiOnr1rRQKcA3DkPorcE59oiaDn
rE90jSd55ZZQN/c2CfcX6PtxHIfiuhvxrpcBAH+nSiIA5G7bicEjSb6HQzbEe5NS
oYAyMD3GvNqZV/N8elbEEq5mwAnYfPeo8p1b7GMz0QMIGzQDcSM0y0+SNwhDM9C6
ff+tC79B7EOlme60+UCyJlx3c1k08iA+xQ4vrkZ9E1SVrw9ovT/XYgdwoHz9H4y6
0Bqq73vPRpKL1vTW7p6y+RwiEeKhCdDC334qyGqvjYBt5KcgZwPM0t1HYVdv2HBH
0G54Pdc/oJgGVj8qO9HzTl68xYmiigCahvvaazK9iuTWvcRDIne46uAgv0kUEq6q
U+3yrwgNHS5rcwcaQ5t4CtF9fI4Jhetge1T400RbOdqLm6pT+I9raijZ7XSIBDgB
684SxHuMdygqN7MWr2RxCXNbwO+uClZSXuojmJndGavrZB/47wJBxMOwrT3KRAN/
afB1tevzRo/UA+18BW2jfhCoZVLjnJ3op2mhTIxb9KNCjaSvhRLrV9OmO3accZuS
/J9mQcF9R24i23OWJVw2odTIpoKTWs7Ed7D8sWkrAXZQI0aXXTVz9hCifU0i00of
+uQz/V19RWVT3Qcay6x3612dY4Dz0FT+VQ3vD459jJTARLLp6urwi2mMEObJG1OA
rCPiQUtcrRMLUaGQgs4upRItxiIbbBYuNoslWDz5iVPohwBnXib4L6rsZwzb4aF/
rpizkIcr6ewZ11HPqOHmCS08wgDhMUoORxpMmi/40X1bM2oUat2znSj6ZNsxxldh
Xe3jcpPAd9LfiBVCOsEgbDKlMqd0yR0aasVAtne+n7m5gByXRr7ASclSAZQpIaMt
fSW9xdFmtYazOnB4P6IGYhUo/I7JTKcs5ahOwI/1N+jSj2XjSESaf7MCfuI0H7xV
VOtEjH1DciOfwzZAkEry38Di1p8vH5Oho9JYSF2nSHjH9p8DDg7HiInhT2s7fqpZ
cmnN9eb5IYf+U7xk2J00sPepUkNTxv5a5MvQhodgR6+LPJj+CFdYc8QFt7ncgyQ8
wInxrMmr+KbmmAxGoYNGumSUnUIdprpyiNeJ3182CjaJec3EDrxGDnabdneUgJQK
TyqHmWdcDQ22ILlGB/iR9Jvtab+4dsqpyKhwuGFSEjaYoq5ckiCgZ4ur0JnLgyWO
fnloF3PDFtcxAAJALOrEnbY1nMOiDLhyhX8ow+L7PzOHn+Uf8uX8I4UlrikmQ7o7
gzGXvagm4oV/PSQU6n0muUfe+L/XPcyV+B44BT/QY8k5QZcBBXxHXZUfZAmQUbkw
lkl/X6SMFDoy26lkeJ5QT/mlftG7TlkvHHPbxgwsODfhbj8swAaFeqaxEDTz25IJ
nOBsXWEJjbRQq+8iBBNaYfhgN/+rsR4DDw+Rp+fuixB0Djf0o3Wb93tEImAfKRTp
cobHIvCWGLvQ9AlZGiRIRrDVYYKomE+t4REpN8W2IXIX3m5U1Cq+n0QnCCmu9WOr
2iiwyR7gv0sU7GDjMKIiI4g4gXUdpFvLpfm/RlbY1Aas2UTQ38FHOtACoNwQvTKj
fCqHPkflqMWcw8SfUhrdo9ONE5jFOTEB7WkCatAg7XKPlBZLhVThdKgxEposRyYP
QfNgkvhkQfSyOVRzyMDIWG7ygQfFpj3M/GOOwfHg/IGMZaPNP74xpRvz9psSulej
IQyBwl1HYrD5qiqZkm4RUUu/eJGhi8tyqk4KTM9fl+4+CeLi7JyfPd6cQAD8an4B
ya3xVvzGXFanZlgtcD1MVK2022yfCeeI76HaiNDLhZZ7jlOE7BYN4tG+3XejQeNe
CAq3oxNp4cyGdyX0RES8TIvxiHEt4Od4uD5zNARl++cvUYRAsQB9dfn2f7MWvV+v
UBySBplmOeYSjG7sKefRKpRsL0XAG3oGyliBkV10mK30o0J4KqSmRaWgiUOp/mtY
KAkhA58gSeyQJJxvy3cRUHedw/L9dpDSXvrGP96JZzk7Idz+yU8HiiMwP4irCdxj
yhFQ6gGbrYC6B+qTlOM3gx4yxC7HC7NRl9mbCTpcyPfXTe+ZjahwcJQzJEX3wxRp
tCjSD1U5YjDj/NGxkSTS/DPM3uCO/NeuGA2quUcfKI7xXO14maUddzNKauFlSYDZ
Aib9mvra1hP6QCRlrzro+Wa6vrVwqgsVhlsWw4O1j2AkLFgp5i40I2AR2ysk+B6s
XHc42HFLWTE/x0zWMOvLLcKqhvGZynkZq4mfdXzQ4OXEhLhMnG0LmO0gZpDCwxKY
6EKd05gKr+hWoNEVT6KxoTa6GXyzmIB0zDEqW5LZGA6xm+tQLqnFzFD0xEEB9giL
hMsa8Z1bGnF6aj3UcmU0hyV/CmVD0zVqVIUUCRQmLq2JS8BNaZeA7Am0hASDEq9x
3dLVcnJS5BspNbYXJBUsKRABSMug6z8VzKXEa5IK8SjnpsOy4VOrr6WneIUQk3sZ
lgwkp5NutvoN8nJHhcyvINd44cfvSWzoDjULauiVRFIgeTZfBsZ2A1mQZsnlzvGC
dsLgK6URkW/s9CacgOAoI90sT+od1YKSjBezNogu+4UcqPdBOH7fldTAbdkIMCJt
pQv8b0wGeEohFAGSXByQW7tp7MLrDWLI2Xpl8mNikuMixChsxYpyt7uIfPDeDsXA
qyqc+vpjAXeOPVVpUMxTtFMuSEHdB7S8sxQtCrgHrwasGUMh1OibFQtEs1x83Dwg
/a78rxiL8WJwGeRXpyC2jfkG1KBw9Aiy3vzau6KVlGkAgcSYFPOvnX73Sx+N0RH0
g8NSyWNrjaneyg1Lx9Z+ZKKSmEs41g0E+h9twWWYYP/qOqag5kht+/7J4M3lDKTG
HibC3BL7LYKuEoksRIEl2idjO8c1hUoTEeFdqbe2sGWc4lLGZaXd8qBm8JHBuV0T
a44j2eOFVPb4k3oqNO6IImmHilLj1MpuBVS8oAikey7JIl2amdGnbyxjfpgOzL0X
x41oYXFRvyOM9yu9kc6Xrn3lXyqi2L+yLJPVtlCje/pMTzI5Y41AJXuRJ+eAjgd5
AezbI6yhDys460zFV8hZcB61khHZxm68e7+k0cr2SyZ/hlOZPLB6PoDZX4yKzwQj
wUTCQdlhimZ6XKUag/wO30XcPH/CtGAfT4sX9W2gTihWblC2tOnSyBpB8xfK1eqH
RhL9TAISZzfYFd3VG6thwgsyS6c9y5ttg6H2bpzUB3WBlQZ0RsrQ1WwitJKFCR2t
PreYSxv2anfJ7xs/JElA7gt/uxGb8lNZXv6x0XgFQmiDOCQMEveTlcTuFwBH1C6Z
ePn3hljDZdXvWxaXNxM1E5F0lcZaunWkWbolrqpYpkRNjO1giELbTYghVr3/+y28
ptQ8/n9BfJh+fleEiXlZbqPqjcdxqoxwUEcv26WZnWy6aQ81nz25S//DcP9TYAo8
I6zfkJpGFQGKevYT2b1n7g/HZZ5x9erhNb47VcylYEubVqY2K5H1R5WA7tfxn9IH
tUCJsfMHH7gaZexz6EPLtPDkFsWCJSKutcg34mpSt7VmcC9xOeeXPiIZ0YCkHWq9
D6wT18qQz4LYxQoX7rV05jD9bncSgBEghp+XCAJ76INGMj/Ifk1Q+90H/H3Sdn+C
aoNfnjl9yYv4s+tz9nPJAC+HNeUWx4w8p8Hf8okUst/2ugheWsHiS9iqVbDKlZlG
wKiiVNWv8nMQQ5lkMdo0ouEZfgEdw0Zes9/r6tvgvVGEVrlgZkhLMH2jIbWA8kRb
IQaGWk/+v0XMxMbrNUOVD8EkK1BiQ7Ky/rZoBgdQ10ia8xW7vfPfVzwB8fsUFuQ5
pZqLXYsjla/mHQgPOCX9+2VcnEJOhiUPcz6mZXrR2Pm6+MiSJSrRxdcOjle06wY8
X5k8oeoP4TT66oECAxul4u/mdKMi3Y3cvQK4lsIwLXjycROBrMPl7TAX93sIgGZP
fXBUlBHtGlBuHV9ngIeAPm/o8746G6OSGV7+lZLbfkKwuQV2ZKRwwa49xISGrQws
5usnSBe+GsluRdthua2gDdsODSunwsgQoboKaEuhRgWxVy31tfC/Af5slfCvB2nI
OJSr2AenKZ+kwe5Qs8H635Uzd2t7g/A58YDa0qhn5H++gpKewaBMoiEkE57jt0a0
2pHCIweqOfh63JUsoebrpbLe35WmdUSCxDj2sdfZz588fNoSeuMxZmqNDGhGblHI
gkbKtGJn9AGbghgBBje6/9BeHwl8GUICLDskkYCuSEuX0JjXWezX1MXgLvx5LqoZ
L1O1qW8tYwPTd4LCLw86O7nwy+Mw/Iq1HztyTssFHHUlOuRgzN6B77o9ERAf9LR3
CMZmryhM93OrA0j1LRrGQT18SwKW04VB2HA90ZkosqQDRLWO/+koyk1IW611PM7D
ZCgg8UEEy4Hq1g7fCR537jeCF0qBXHbi6DkMqBRfub8UYmcj/crlcaJcJLdeiCeD
upa7X22Q2rxoLVYBbANfHWLtvHe8F72a74cQUflHcuIZoBDic33fiu7ylkIb0qhP
Mubp2wTRJCp5Ybt9qnhhvYDeWWcTMqlfxzLKTZj31l7hI5h25x6Q7CqTcTlB22NX
HlhG8Z+w2IBtmm/MQkjS1JhjO9IuXacykUxGlDJXoUHgi2kWvIHiUjasQ57ALetB
K3IWcJJxnd5SgjPqdWOKZjLPNjKLjhqcOsEmNbaQF/0kFWIDkgkSRn6qGAKcibrZ
r+zPsmN1wg3vYgWq4M9RyvOCMYEBUgHyfA1OXMvFjyTIw18XKTgd+4FcJ4BehczG
XSOMKB1t92BgPKcE6+batAZYaYpeTPj9k7/jCsgjwdPobs4pC9eojny+goCZispV
L0tdV80zIZQpif6BjkHB+8hEDNyq6jSn+VGCEf9t3DbV1mzHEsSWcw6a8J9Bms7p
MPzaMjjC0W8hldDX6tYipE2pOMhfG3LQEjTVRMeFtvEPDx7bG+RHX2onJ5WJxSEC
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jWCM2MztuKsE+vdxRD8OP+7NfVpVFXUXCKOg8y54FX0qPjG6WNpyrsJNZsqePYDB
70NJ7i+6GDAIclgtire/UB6CUQNO0MLJ5SAO7GPGnIXptlBfRJ5iOjgF/kmP/F2W
crKc5n4+SuBEp9YJ2a19Wcxqnk4tWd5nRugStZGTBBGlIDUTkfNvHwEPA5sKhHzj
CFklJVveyK6V8ZqIhxEo/6UEIl0xWM8LQJ4WYGRUcVmSugmIr+sZPNLeQg6HGz1D
nqh/LuvhRbugMnjjdzjYnyWZLkBMGYK5yfYjaPNxDiBCz34xKSFYRIHG2kwTXT+b
N5JKLbdiV6bQWA8WtbDLgQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
ejhB/mruDe4jOybud+bD2c8JWNx5KOwkcEG33lQvFveAdouyAjTdrs27C3mf6iZM
+BCsB51Hb0hbseCKyeB5ZinfpSexVjAcwvgBYUemBjm7/Z4OSvmCH2ocGJ5T5q1/
m1UKfK+l9pqLL0Ak6qsCA2YTmUcRzciYO7purZduMsl9DkxvcV6cRdiVNsabaVvb
O9ogSzUn3J0YfjQdmasMnT3jtrsC3/a+y0rUzKQWPucU7hG+oqGYD0n8GZzwcq3h
M1krfg5ZSnrT+KMSDlJ33xnZYxhE+cClVScYEIZCaSKDw0JMVnDTIKaXQAJwiLbd
MDX1yPgLuEZ7CIb2uqJc2aKutkaCATBfy3/tznxoTRfmpCQvhzODVEcHjT9dpL0u
e6Qsb4R+xFnKtl4/YBSOFTkpkwEbi3C3gB1nZFTm/CtPy5wk+z9cBDY/QGPDeIs2
RW7/ILYnZnzJ23VEEzyQLX8B++u25Q4JRDodLdYJOhBYIhwYSmFAThBWswVXSq7z
wrNzzD8y/XVw9wulD2hee0oI5GgQ5HyJeFxQqWwQyTi5fxxfHnsgzt6h02kRzxmx
HEcHMAT9pE+MrlFs1/TBQkWbK+k+QABQ8mZQe3XRe4BUhDoyjUxoTBoN0ToLWo0a
xv0Qc6lhbtv4WDhCC3m2lq5H/ElFfG6AiCooIcyrVM4FrI0RCyAfyb7NgzyCioTa
dlwKJSFx0L3dnTk+il5NVf4KKrSgcRSamnzUWbhR/uoXLTPmwMw7Lip17ZcC+j+j
0bk2pKjM99e6V4btTi1OyXxv9fOGeSLJE3k6AjrTiYDQ/AzrO5IVU/IP/W7Bn8rm
nF4Aw067t0o+17sAeYUriHcXJsQVaXJJe9lrReZ1yjqXxhYoO49QuYWziLuLJlUj
9wSfQWFClyvy5akWERPGgNqcs1Wq15vEteZXpMi2EdpCywTVvbvGxYKcmW7xvsX2
Gz2JihzwESDy4AK4MoYeZM9WsYX6OD/YRJwvbckwdKz1p6gpZBy9kdn9le3PlidQ
vMhcRPA22CxzyUFW7exNvcTVAhsIKRp7WcmrjqVQOwxdFtcSv7ykkqlgjztgBw1x
Kb+b0bBRyKLb3Siv+8dHmVL6+2I2J66ZzZ2eBT9KkwUb7qhS8D+VALEce6nqBZlB
PhyGKC1p4QdrgGLef+GOnC3CfItGRrWsk55Fj0h7kRuubYFCoZ8KBTiARyoXjcjn
bj3CnNuJIsYbn0RAMKnxZyka62uoqWqcSRIGNrD5wCwxJrszvdVeQQ7GH+h3ZqiD
U1pHmdwHNInMSWSuvNY7Y/BKzZkktNmRT8/1rTcFOtstRR16cixmyfS3tnu74KqO
hdVBa0G2wH2w5xvMJ1wOmMLDGr9dkxdBdoohevpjLDZeA+TvZMO7Eqcm9gqndoaX
53l0NKZjwm3jUMtUYmiaRuR06yxvjeEpi0Z1GZV4pcucOM9SGhR+NcKi5J0iaPZ8
cklTYEZGZ/7R62FGjndoyJq220VRkTLfe2pJjj4Q427D2UrHjGXoSS1XniEMbBfF
ZuBdeLTt3EekhOh+4kXrIqRuPRCtJJh9akTwX6o8RqmGrN26jEyAVi/E4oZvy1si
sgP7teqlMXQnyWdku8J7NRdj70ugouFASxif5ekNJSQRbHpShDVUX3dJjHhHzkGR
Qz/b3JS9k49Tw6z6IhEdjgHW3mkngj+kf/4G5cDrABA2PFK6jrKsYfbmoLKSBiVl
PXtERmwqbJWtgLCs8towTlGammfu9kC599dOVh8cpzG3a87wqsCDX3Grrk+5vYXL
U/037kpJosIPcwBGtWHli9rSCoNcQDv9VrdxXvt5gWNqDGJNyxWPbprUljZT3J7U
YdcqqEQA61pkMza6Z+HozuT2FoL9pJ7CSPFPsMSrIFaN7rnyCsW7noWmUFvmapam
v4bHfi8BeHl5vPL36JCewZyocA08ANplHky8hw3n9uI9RN6IMxqzfXsU6azzjWcl
HAFzGzswJmxQ3rphIFMOXEP1VYz1W9yZMEmHHkDdqfPnhVZ0JSl7AS1VouKIXQXy
HXsemE9dthX3Qolp1T3f3lqp3RLy2E673PynYMFUsWTNE4mqLWZurTISPjA61QfR
BaG6BuyUGqZn6WTm21XRloCGcfjcZ7RTIcEKREbXMLhGVPgexAsslnUbh8TEgjMh
M5n0WnTY8Qg0yxqZM21YARM88lfLMa35oQDb7ZHw9ZKKSU55JERNLWDHnOjQymHE
mk8GicQccJMYk50/6HlptX4KYG48d5AAlleNd/38RQMwz+1zBCy6n8Kstlb4kw3T
93p/mDaZk/vWqI6aAWO/DHjWcm7L00ULzcyBqric+cNTDcv4L7gs6zr0TXZT1Umt
sEvZDFhlUCrPsTg2AjQZEszcsckBB1isxnlPb6VxdpHacdsiydx/HZ5kXwVEo4Rw
pbYjIJOIcg77rU8VEtL21/n504hpoMic//BrHLF8XvjdctuoB9JExnajjP9RvVB+
dIxbbTueKF5HiAnOaT1iBNq/va1uVnbZQowrYCzjl07eR3xO0wGRF3UJCj2FMR/0
nyBocrvR6553k8cdlp/7sCGzgN0wAezTXoZPZYrtUjHOhcty+/Il1e/NLJs4+jIw
DevSb9DYPtriJdYCgFQI7Ec2KrNYjKepNnbsNOaZGrHsHMdmuZICNpIVu2Ozs/x2
yY6pcNQrQGsJ7DeDbHTCN4vncGeTxGQmCM09IPRtfVnMUhZ+m8c7DUu8mrB+lm5Y
rALwhg92qjkBGl1M5RNWCb9au7QTnd2rYhynMfwWWTw7o050Rzz9SrOjsGkzlJ0N
KNDRtOMpnraQAPnYTzc2Z4Oe5my8BkE4FghJjZgvg/AkFUIzkDaoMliSGFHRXUYl
OxjOgTUiZowdsVWRqWdn8k8cBsO4VkycoEten3xnU4m81sxzYcPTM5pyUIdJDpgO
JJn9WRu5dRX44UQEB7eJNBnL0tJ+bvj7FCV0hApH0OxiM49NptPYW10rrrZ5v4ld
/8Kk0OHUk9pLYN2n8/5Zoxpc3DJCRNPBqOE7eD7NJpG1IrE3P/WYerNC+VlzYkKb
VaLaUu4mJJpYNREDE6QzNOOoSCiiva4eBssdomP2Lo8mzdYYImLAYqZFoKflVIvu
a0J9yBCYTvulypLqQPKaAHtMpBdYPHwO3LkhUgttPPFn3Cq8ULOR1riWK01ckmTX
JIB2GV8tp6QTR0nCdN3f6Xx3MCCtQBeuKvdLWYypHwwZ6gJ+cy4Ae9BsfT+hECch
3yv3WYMwDA/JZSuMFmN0QVoEjz6bySamufQvyJMx0ZSXePN/T7XMkn2hIaq0l20i
4zLVOEDr8DmXZUksIHsLN9UfB1n8rZgUN7712D+8Av29l+H4a18LgxHESOBup6Am
ihTNa03wvbkjrky5yw3VDvcIMyTVrbgShjWL89uy/ptgpB7mYtwd2NN7jdGMmSH7
9HaFJNksHWpPpu7lCyIo7V5lgUc1jpdc9zDYQCH6g3GoJXmxmppvEvMlUQ5mSbNg
4vHeudjLq/E0g9GDcwLjZKOYeDPF0UxfEQ26gosfks8zu+ZGWPNXjhA4d2p0tQMQ
LLIkHir7UO0B+Vy/TKjFTDDcQiJkIGDOljHqy8MBnf9holsE9MF444xXEHJU8r3l
ESMT9Zk6HChIwD/GnvswrsXcCabnCdWPT5Fb0pUDY7sKUXlcw4SEbPkAhAaeflmS
KXH3HIJFWtkBrdTN4W3I69Iyb8WY/tS8UE9ivjdddtI93w4z+IpNRmKen7Ef1pRW
YLhdM0CCMPR0fpmtTMiRvictPrxgd0F/cOgWP0liCdOnpkTjVHw4poMJGwPT0fBy
Ur22uDYMWpS2iNl+Th39JlqwFCJqi0SvSj4aVqxid5ZsMjcpgxaOQrn1yVhV6OAG
DVl/TrA3cSMDxlkAtmLdYyy2BWVTBWsd3YN8EH1208nNc4UXZ7Hf6w5z5elffovi
Lu5GToFTBmAku7EgOOWo5apdKUyGawzSaXyV677A5sY1TSMqf3a1WrKq76oXt0Sz
oq5ylV7C4C5d88o9Xm+JSTGVS2yFkjVkCJPR76mo2JjgeG+zEhxZfhwUUd/JWoJr
QtCDnElZQSg41u11kI6bTAq/sv7IbQWuuyLPrUQ/ZUvJ8hY6HwVhDRcdrUzfINER
Kg7P6dz2HKaXSFYGEH0Z5vIsWtUfDhTmxP/oWyajo/u8Y/VyayAbhixseOZWz628
VAPJI7GJlWLxDvK5OkfZgUUTahzQgH4uniGu6QmCFhyNr1civnD2V2upGatHs+g+
5ZN8DsiYPEi2rYileIS2EZjhgX0gCggQsNRy5OW7kpFRDmOcJEDzRxhcekbf1FE+
+eWNUt9OwuS0uR5AiGySIzP2h1l13aBuP0TOTWITCq7EXoOf+o1BzEm2revm3Cxr
a/qL+hdxi5gxLlEE16AuQ89h7OYquDXcMwRQkHKHf52FttDSh+ayx0fzj8kwoyi6
/wPHMyqBV7sRtap/lv5m2cZVvmvaCYt/J5GdmSYTP7pDIUgtI1PV3mN7Rw3Fj/SO
uR43K3FapZTKejYS/QRId00hbOrK638RM98hl5wYkVhLuZNfEKheKK+Vko+k9q0a
0hHCRsnW+F1/3uFT3138//cnlX8VF7aYYVty0oiczO6vDZYOk1+5WPlZvew/5yZU
tlhIfBzAl8eON67nIhnQa8/98K3HH5zhl3YXvb8ycBn2exLApTs8/6z4dsb9LslM
zyIM+EERiSd74K7mwdTpX3SRmwEFDye3IMutTNrdb8wPLo4KiINOmtBZe3Yigck4
nrAhBLqUMQqY09eI1hAT83tr2TXHdBDaK5/4pO0QmvSXDUbs0jrv2BKtDzp18SRq
5LS8IGFpUxhFj7Zl3iqgnW+gtReUxCPkztCUt4s/7O++7OuRuvOicXNOtR49uniC
wXao8P38hhwvZ5VnjczJjgNLYZ0pUJ+LG16wqNQfUKrnBHXqiGlaClB8Iar0j2ES
WdkDpoBVOXjM9u8hFR7KdjP0OCVT1QsTEttx7zqmnp89R9eX/MTBHpd7R5hnteos
9elXaHZTFUHTK/3PMtrFz71+f2nkI8ja79fclBG9QQY4KNW7yu4eCHmt0GiakrKL
r0K07CCQFZZRYXhJRkhMXhlgyLm32j3eeokLFiHV5oM=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
PCOPaNyxnoAkmxEb2hV9UN+I7KcUx7pnPi2RR16fRn16mMELjmRkKwo9YvryEopS
14pVM+lblCFhhdpa74OMa9HLrmJJThg+teyc1XWp2b8m8yfTFXrdHhr66hJ0Kzy2
shVajwOdTH/DHu/hCTFuiS+g/miCRX7gs0Cp4DclL3lwh64TpR2V/msxWcCuBLWP
oV3AkSE50yT2ZFQbnQyFF9evqS/WYf8fp2nQ4UwC/j1GQZoKsSRtrcz80xMfE5s7
1XFJZt9TLx+F7EVXa6Qu/RTkvOb+nu9uFzHNXu45sgbE6RfKKe00LENVblM+ZTJH
tFrCR9M6FfA3UNzSryZPRA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8288 )
`pragma protect data_block
+EV8797KnNhyUWW1yjX4hQZyLXOeCXmG1ADQstzqbQLwsyL77bK7VlTdYkCFbC7f
FUXAqO3RYuVFqbUkzu2uY9tSa1yagva603MQCVeAe2DOumQg45ZTmWUuReW+ipXL
t0vhcpra3Qq0GOpUwtGKHuMqTywmWCeRql2CnL6o32BmDwXrKUVTwbEPVph4VLjr
rGrER8YTqhoVaiYX2v+JlaTvc4clFi/G6G4TTHBeVmZEWb0lc3EWDjE6USacDRrs
mvWNHjjo8ToXs35PZ+n3Ythcff/tNMr1n33JQv/s9CS+Y824xTRbSoZRPUgPRwK+
QiioGBLZ3JoLXkrwHTWUMU4a0CN3ieLnuhVRYucap8y9t8jtpq9CM4f25xVC8Bng
5DaVZhjXgSkeUwUmW01EecRFDJ9xDb3gKwM9KQjAJLKnviFrKbregdCbUxOMuZq+
fYuz2Xws72LFUZWPx/VTKEhDfgkMvtYf0AZXpMMH4j1tZEDUOItLWNQvBdyKjbEj
nOnX+jQDuQYV+YyXe95W1VXzFwVouogD+F2DvMA+mZJ/3fb+UC58oK3bJOS/PqLM
HDTJ4ZHBea4W09K8ZknM72Pu7VRKWtwIBzLaaEytwYJ9WJKKP7xjkgqs6RGEQrxV
MjPCOaYGJ46YVNzu3ugWoOvchmgcH1MwagbjDD7PWeHNtUUfUyS/wZrxr6mz7axl
b1wVJRfJobbsdR2gO54/+vofIWIRFOc7PdxJK2P8Mbzzrz9KGC1He/o0aMfvhI0C
geyRFZKSJzbr5IJPsVoG/eSITWGlr5Un9f27SR67i9CtIds0He/PMNePAC0fhakS
8vVYVhOL85YgcfziwcSBZW3BHASZ3KeAv6wFF+fIMceXdgpXgn1FAnv8KODGp+Uh
AIj1dav2jR6+pbTHf0EFdy7843PG7qVu3lsjutc0DbukMQ/0dW6hpqnyeANkBZGk
mvND6HVYFi6REuX1bMWPsqxE5tbc0a+lkrC1+DWTsAhuBvlf7pziQ+4hAPTgHaGr
J1C71mp6EX+u4oddysTW7JC4d76WZ4NjWfYlvjVIELQS82mHzVvobvWNU+UebYWc
KM792wro9JNnHyHyezM11kayq5VtoBfAxr1yBvU51B6d5d9Z+W8hYtOs3j5VZG2J
f+YYHyROlvZ2cP4IWyEhkR5FexYtlk1MQ1+lkia+HSme8Hay8l+vK8mqNYkcnzun
bwejqOkF4M+1v/PpVEvtYWubi1Qk43WlLdr4iAwCOrq/+sg0rF2KHnuDahbAl70s
4C64ZXlw8kkuPk0GTYkC6tsmCvEbYGkimWKYwXJHlEYlYXdEKeVelGpgSsDIVdlA
AAKrR0sF46Kgtc5s6waKgF440zCg0OqRDJE/0bVNqkU1alpeyfxCCsQEQNf1vJrt
mx08xE5gKa6aZ1Q+uiKWxrOht+9qQfsp3KJj7GJb5jnEO2f8Hic3UI+p5mdR/XLF
T06ecVeAYyEzvvBN+Yrc7OSlqCx/ZENNcmJHCd9EC6N/f7PpSwMYfXnY6j8Oiaib
LtGcCaRfF8dC9yOHsnWMvuzaI59rzVIp0E8Zsg8XvdeO6cw1To2wzb+lW+wfYj/C
a59wZEbTQYs9l8UXE+dBb9fGc7tcfcIyiKyudVqaDa3zIMlvILT1I8FK4Ewi4bCI
dbeduiEaAYbOcRanFmUurr6C4AyglClm4gIfiDpWmCTYJkA4BaAATVEwM79YQijM
cc4qNdpG84Eg7bS+onjkk1sb0aytohtmm99Anyvn1S8pv1Iu6ef6blJjtIIgzUaj
yQeC3YSRlob+Si7xUUN3889Ff8ku9EoozB56mKDtIOZiIKRSDvyrHmMfgvHcpcXd
O7m/ykXXckYmDT19ChNz2CvahZOaPQTJtv3LerUAeSKWjZJx+N9crVboOEX3rXmG
DHY4N9dihrH9kF+fy0Xtw+baEBuLc7fsMKUmBf5YbNORZ+POcapCZrVf/j0oubr+
NZP/5ZK7n7CyY0YB6QvVnLtuOeMLpxg2npRk0iY2Z1ZGMlt7RnxJWL5DYjGJv8qn
cY20Y8gKE7gW9S0X2cjAFSN/enm3wIMVBQux+TcljZzAqegPd7kNuEhWgyKmeX0h
8EvkbwzVhu3KzbRsL330U3jyJKqnib773xH6WUkroBR/Lj54u29CT2WG6e2G36Lp
Q1AAtaQakASwZCXY215/3xTs9c3/BVXFOHHNiTyRDd2x2wEVUJym68qwUXU+1NKN
KeOe2znvCgylepcR6IXVOWQqoPZT4SOySd8Za2rmN5GRj3HJnDUmU4eaf//Xvy11
U9ZxTUouVyQ4rHYMw6Z2nAw/0MylyprfYZS2q2fm17O3TGx88piLnFX1fqvECA/d
8ErNM6i6aSgUky/21VfBtIk1kkazDCFGndsEuIFkBDp5zwkkxkCl3mkhKETUGzUN
nY6O46ae9Q6mjSdvjfzrRro3BA8vsfIGapEwI96R2iLfgdh66dHCte6SfGrhIcXz
51DFG9FRiVLY5ew2K6+zA2p/VB+obUpLd3xyCa+94fBW+vSaBr2ScQpJ/7k9x3z/
pTZpLErnq88KEUchm9oawJyUwWYws08SMY2mZ9U637SMw81iq4ucWsoEzaiHfDQZ
KQp8vWSC4XAocQ0x6GqG1OlltosVt71oBovYaxLfzCSKTCyNSKDpDUHMWkanGaKa
LT3LPVY81bvXdV9r96XDPZ06vX8zeV0JIzmaUFUTNB5CbZS1nEIkXylEIcihO02X
aDtfSmNJiw+j2pCVqajE/x6rk9HxxDV9807eauGtaWCHTK6SMQ7ClLzwPLq8Kchd
fx8X4MRYKW5fGd9lSBI6sTwnVgXTX4rHsEG509/hk/g1CzflisOlxabEoqcaKL8d
y/6kDzDqk3LcYiQ5qwnByE/wGSomnnMmEH0LBJD1zpTOu9Ay4G53IKMOuu2iRH8t
BP/TssiJyymQ+9nZfUcseOh5sJOzPJYM+rN67wSVDdQ7cNnLMrC6a7etJJIroffV
eZyt0XoxhfQ6VVhhEHVvE28qgq4Gq3LYrMapBEZnLyF2NE3NDQI/p6qEDu5y24z2
qiiUNN798jndgvPRaxi+1E3K1vL1ej7UuATCmGaWaxn5bOYk6jL+2FvZ/dA99PlR
SwQ5DLYJ231ar5h2rlN8XOe0Ojn/Kbphlf7VfJ17DKCHywZ9oHS5ea0//IylQBb/
dUmNMlUlej5znHUPT5xmGm7YoLLo1eoUnBTDOOhG39eWhJKYJKGLfrAqPRSvUDL2
Q/0gnCB+NBa6yUQXdRaqOYgnLpftvusGtKcihK6BTxoYQvLN3hTRvJOnmWbwgQqG
CVkrEpBJmUw79ZloM/gEcy9HjnE6rz5oYa/Tl7OkbHSISHQqIKf5mDDfOyCYrtUz
DD2jbj0rR7MySuzUjWXH2OWU42yd0mOe9GeDeK7CScGrbtfWxzkbwjhcMhd1OF4a
mL6VQjxrSzmjctyX8BM1HV4feI5QPM/I+Y1qO9jSz+0zICF+jwX08pdFC0px2zH0
g54LVw5NiyFcQuywwWDin3pENBIwg3lwWxmzGGyqEXzI0EeH2+oh+jJt7tU4ULwK
RgAfMer8ZPZVEygXIBc2wIgmHMULHXgPzq0OxngmB5Ya9NO7NjOFcIxQvAHFfnOb
7VEhAEXmuvldlN/HPE6k5/Np23gkaYm1bcBKcTHz+0EnJk+GRcQea1Y5uPpEiC2j
VUyaQoEIkJaEDi6xtsMzA63QEcmbdDG6x8QcQDM4ozo/XcOPwYnd7VCUKaHVGpUn
sc/PaRIh6O8032NHhGfNOV1KhG8ZRDQHA4WHjMxw/Ga+iGG4FKj7oIB9pOi0uzIy
8eaR0jGP+U8VcH1bjXHSMdXSmCuhYDRkwWbkOHZ7DPpT1s7STt5mc2V8ad0d+inX
3BZ0q6LeszOl9ko61uPGrWinWnbArVfKPBNP1tgOiSPBJ1bKK4w1pmjkSlMyFUyz
Npw9qaP0a1HdQvw+Gi7prmXz3KypM7SP2qLqalPrloFtTtndc6ljsf4mG+tglgLL
24Voa5W8qbrRJCRXAX2OJ7I8Ex1nn2FtT+qu1y3pi0AG+GUqeNxODZ89UmugjWO9
rRdSSkY5aAmCwPbVOE0s/6gNTKR8xJioN/jzzbwvU44KFTh6JFyAnBCn7/1h+buZ
E6zjleBhCjqibiV7rT0S7HYjDjJGekhnCj+rQ/PAFbChCZbHmFj9MeAboSDKQOrT
NGV7Nlhgzu1Pqx2zPHdxRPBA58nAt6l/XJzFbp70dyXYknE9aILRz+6KupkKTZPR
NI/lZeIlAwfph0lRZqJb27WppXIBrEz304Yq/eFoOJbM/bMcBRcIPvweJ3f88d2p
cC2S0exzUFXpzfABkAnBHHBeJTOPuMxZyXBO1vDJIGoejAAv+pZAnPvDHuGIaJtr
rbhkRwuRGyF68iC59/lrY/SWWJqj5etfE25HgciwfMHHB+fdqEKcZxJI+na+HRaI
huXTJfkP7kpxqzdR0cg4CDedn/JObDIHGb9Iz1I/Z3DUMEo5QAqBE+ombzB3Od0m
wTkTCyQZfu9vJWi12WgrOWy6cDG0otKm3FD6RZBpvzK+lfs5gWR2o7d+A9Ozd3do
kKsfKUHKk5m59DsUcyqn2oEKabZyaxM4RV8w0JCcYK2NrqlVINZwcrpi+/oUUkog
atJMZRYx1zunt8UJVWhh2KPYWibdcPUQq5+jJPySB6XM66droNpvktv0Nqz4hgKF
Cv0WhFszoZ2Mg6hgtywE6ufPbHfnUKAKNkqL6N+3p00iI4UL67vsgrgQ3IyYzSpz
gH3m/GOQ7F1ufzIf4fHcpB1QJqDAyCNo6qgqqk0upp1XqyKXUIZC6fWKkO2LcPdE
36seiVpZ0g/Z0S3Zayh25+SluknLk5ME9EPuHSqMD/oh0CZlVSfWXk7+hMg24yum
9RgkcnxysuFw2tjcKPskFK9oZXyUnRvvji9q3cywL8EYJCUObzvDzXJw7Lanv3bX
RiAYT8OL7DQ2EixXu7RIwE8VkuxgIwFhW36XbPreBU4LdvVBtzN0+NjWjwSSS7TX
aFlsD9zm5biCtzngVoWu3TOH36gpjCwmkxtQTGUs/1l0uiLNqnmj1N7E1yCzlCCV
f7KtbJiOelyGweBluEHdab4w/iQ1eZImnEKB2fbl2FhozuoiSYtifslyU4vVx6V2
y9c7mHFzC3+8CMmLUZf1nbUWZujCrnt0BbNnyA22TTulwJSAM6YH+WMmZUMEApfw
JiDkDiEhe1jUC33ZGK8IlpB0W830/beBgUxyT2uGLknSu3hvyF7f5jaH5UHm/mC2
5I4mHoHQ9KQPg2fpzgF1ByjjINoCeYSPt/TUfUccAfzCefQlvsZ7xLBK78ITCXOH
1sTdtMFc5a/lw3xhnBQrZ3rt38UAe7Cof0zN/RbdXW7PaoHRUsBKWHJ0iXBf/ncN
Ypfxv1enemtGjN9xylwoiIaU5QzXv/U3n3cWJChYSAoAbgsSKg7KYeoxFu+aATs4
VJcQQC6I+BWqThS8GzrCuGtuHQAEIdahSjdYWEXgsoKQCkpi1TmCL6XjDsUg4bNj
3Y/geJVaBSboDVMS7uJyONh+iupoB7aNvdSBBWllXeDWMN2+y7QhldfJ4xW5oXTt
dQX4Ww6xJSWDYRnTATzc3NwcmlEWDdKx/3jIo3qMP9yDJczOuP04Xu4W1hH+udak
DRz1KlWSi48UCR05Hq42tC1lZwr3AdkiDZ7gbTh5c61n3npNAl0re/GIeUxjTEq7
GNgy407L26rLfzfk45TSItLHVLYb6+eWYWJTUUN5IRkoF/CJR2AkeB/pT+4tNC3/
M4Fqt6aB79KaK/5Ya9RedDCvkE++e0eEaD0w6uT7n3+KhE5yvmEss16lM0IEMiIa
JIb8b/3d5jTpI/TQqAXICDBzEk/Q30FEMdA8EqnW+/FXUI6oMBCUIp7bgi+6h1KO
1TfttcJDzWMbDSppcAaByOtVJxKPS9TLIu5qLSjzB4rOQajyHltR7WBMofMI0hjn
5ldXGU3FD4SQ8h70oEgGpR7NaixXCUNFkOO14ulc99sZ1/kXAcv5y5mrQfMir/CC
D0Ji/Ab7g1vBtUtJn9s/Z55ZCWFxpyHcMQstaNRGCLDiCdFZmGOZmKjZag90cuoC
Fa+HqN8UGw5xKPqznjl7LGxcvx3ZmkVkHEc5v3qopns8SJpyafH0oxolb9L5JvvZ
mPbPf8YIhB3rPBVJJO7sJU//XOV6LVABSQcnEJYgqAkl2sI1cY5HmofWfvTytSBg
6jfxTH+DDQ1Xneq0Ao3oPp3/SMGyPiBZMXJd6o1+ZwIo1SfHCj4zEVd+NZpiAV5b
28D7rjBPLF4MRgiLH0p8+YqzJ+CY9bsrdqiukKbWb7BK6gF9j15em6FOouW1vAXD
9PO0Sq8YXkO/nnGPHh1Ol3LvENDhH5Gr5bkuAPRchUyMJiyeSMWv/xmMutzJdLmO
PG7PRfb9K7bVvbTehKtJdd4SxfHz4xAxPZyv3FbYP79we1gPmNrgotLocsIdDd9q
yNMKD2suDGO4CHYNm42OFPKP1gBa/zY62IDpGRkKhgJ+6trSIRdBk7SRtls8g6Cr
spN6IhV0Cn/58n/30NaFtFbx3FcaqJuB4HleOOT5OLVCLMv69Zp7YBpXaelbyYCG
rfAEr26huOeoFazg/g2JAtEd5J17MYCBM/HSPMXSIAXjxxhti6gYP4iyWxwFxZhw
cOEjbqHV+Jk/7i/9DcXRRV0aFevMoS+n18RJBnIKSCQYnwcrMfw4ox56XXcUyNir
2PitZGoh8027zWQWxrBqRv40LFS9dfl6yrflbM9kvDY1kpq5N534HB/jjY0zKCYl
yjIxR+x/9GrO7sj8BbTMLwVNJXRIVt3z0HNLA9fTsX51/YYEF9rvtM/u7PCtmyqn
kIbgbEYRTsMb0hf/kgk7j+om2MJq8/TZ3pjYahSatTZQpj4an6iRW4RoRwN3c9c+
nSh/YO0oX+vmsbEmWxKaHkZA0UUJHh1UxqtY6nK49gF+oURK6s2HapLJchc5CVQg
F7EClEJrZ/zkrEUyFl26pLsjnR/fhvDGWyfjS2DL5ywEc+TyCcXcMZeTMBRz7Lv/
Rs3DJAHOmHCvoPAVH9QLBgW/fRoJUeUcs3ncytq2nQrD2PD/Viug698XX4/wc9pG
Kj3SkhRx30lD4vYFpy0j+6EEgCuii5UQdz3He937bRzk9K7bJy6wXEwDsfkaBYWx
nB8U+nVIIT03Zz0UqY4h+ZBPIEOAqlGiG+oaYtAxoz3snuE4xnm+WBCOAO0Mr2bj
wqVuzX5LVK8vUIJjf09MAUDGEy7LSDKqP28aUcbtwj4Zt1WYONn3uYYYUsoHLDra
AzBUmFGXGCB+Ci70nDfWbWXtY1olGocTP7ZxhOwSZtOLO1fw6nBGbQpQVe8nlCHP
7azDGsI5APZgDBC+5VEPvJEUJrUbsPaqxQBRW10dqSYipn/K2hm745rAtUsTYuJx
N3ZP94ApOb2v9dxff4X/Rvp94qHoNBNOXkMfldpCTt6n+nU84NhGdGNdQxH8/yw6
rQj4ZCAt/aSKlrVY6/cn1SKzbRvAT8foSLbiWxkbpLurbYxPOhq4QEiTOP3ktry6
/8XYoKt0+uc03XtLEWHT55EbRbs7agY4DFf+WzeOqI8soUPTstAZqrBAGTjK2us1
MQuGVccMcq6yY2mus1C7oDHdOznn2cmO29dS4UMxMfZTTg7UnHw7a0H9byY4j4cx
ZWWP9bKs0ZJk7ec/qQN77beEAekipuJ3qRnSNhpsxQZkicpbQ9MTvErDMNdaP4NF
J1yC4DnrCeQBFcFDCbr/IkONz1HqCiicRVul31a7Ot+eBUpihziW9CjbSW0Ogw4a
RqIYWrARgfEuCl0VYLoOxTdHB2NnGijZOXSRkmoToiSZtsQs6e89VEcyirbZhj31
dmHcP1iK6DCe5cZsrXS3uofikk3tAPEpSqBEAN9fZes7+yFIWqWB1wM6XmNlKSeo
BLUUWyAtdHlJ/fklLybjA6hSlLJ6hWbPJazpTzXkhTd62hRYWM+V/9Y0ghv+MK2p
r7e+1ndKas6sB4m68poixiktrzeLyN88/c9u4nBdVppQNBchWSoFKqX7pvEtxwAd
wD5o9ND5/YpDGAEvvJVL6HYvccnJ7qL7AdLPtER774GuG9SPcZtxPJ5MKxEcryio
5ZemRjvkSRKV5Hmn8cDSXuli35F1l2ua3BsSWwH8t2D/0Cj4bcpAgZr6eawwhWAU
ZobUbXJMTUYfWlDSGfYEPvmaFojj5PzPbkfA91HA3ohvIotVyNCzfLP262vjzR0P
ExPcMo6bEbbcd2pepfJrO3axc2KORZa6ZgLCECTgZN+F1dd6grU672Ez4RMCnlqf
lHkUk31sJHBZ694dMjqNbEg+3P7IOjLdUejwS4MJFgqdqEkS39opYje4iwzARYMF
5MDLr7vNzMHUmMXoosGNwslvKYXbUzBLbI8dINLWW8MdBUvK1CLRDv20x/n2XUs1
eq2zbsnYITqdQwcyYEZXnuQ6iw9ZJuGiRnnR42kJThl/oVsVny8Nviju9k+2FHD4
7+tD7/sKaOpaT1Xihd8RtJpsECZiPCUfsGNW+4CPKw+5DGYP8IhuonBFvBr7k+xn
E2UZNM4WUeXeAATfZ9jVHsAH85pynsxuuLu/sWafHl4vQzo1R+bhqSWJzFS+rvYL
bgG4jSqxCXrn3aRqeAM+jm7BeYuEH1FIGx55X2AMFfSkHinkz9bX7Is0/CcC/1BI
12+GQPIzioQSCN1Ie3fEbWCwIA+rPzUd2Pn8hgzQcWbbs0qCh3NddJG5EMKdc26y
Dne9m6pQSkvRqfkLEGzT0Hm5Xk/C/noX5dfCOXlRL0RIvrIntj6y30vjQWNyHQir
Mcqt3WatCOHAjewlOTi7zboTB+cwtMPJHchd1v8K+mW6ReQTSJwSK8DhPmp4rfLl
jLH4QmHNa8DNJLWJ5rq4/8d74gcfVBmrJQepKGaambsAEcHbob0Cn7uvDwujaQul
U0pBDMIUm/hwqPImz9ytyZe2WDQyI31my/sJPAVt18im5aCzVIqoFmgdmGiL/MN+
z7WaTGmHUmpF5VM5Q4QDmm9Jl8GY0+2pyjJ+KaFhJkLgvjdpgY5yxNin2LmfNtgx
q+ZHFLpv2C5yKZela7xhdLfmlg/pnG1NtUEQlPP+5JFVqXBF8q8/fxZ+T38ubEYn
jptb1H0XRnnrKSiElKlM4FRxPjP14q5VD4Js/yHnK9qaYhgLw3cViQsv+2OUSQ1k
DfD+Hz142sBneXqIsv5NR1bdmwPdCZ90nWW6uVqc8a4DRiuxy2wBx6swlEneEppZ
RHd/IwLw3Rzev9lUO8HoyU3GMQM3NKId/k4wFEGbNlIkliBpbphSA4bUFxoxKfI9
DThRkf6lK5PhCU+ex/0iscz5GdZFXLouQ9xQb/WKiuUKZO4RX3kmXJEPtFFHSTI1
M5qpScB/8vA+JI5gv9CzH3duz4+ofpFh0D57a1xRic2+qMqfBY6DKiDWvRs5TEgE
PZ31hNFFQH4tDCeOUIoMw2nwZkOtgpmheDzIFuurrwijmidd6gqyWl6XIOKfokLJ
1fGYqj9IGvAo7OpwTyALkLv5PGz6NQjphL77h6oE4RVNg49e3AAhN3ZfXmTubftP
+Yy7q/NtHvo+YBPLJ1BOu61MunqhcH9B7BQBJiTAgW4Mzzyih+avgu6J2OlaJd7+
PHYmOYiVUMFtbqKJ1BsUwQ7an4DsMDzXjtJFkkTVitIYWB0EjhwP69ZNxiSF49uQ
wqRsLHaYV7izxFpMnUJ2xJEFmmizzC0YsGwxlx3DegA2YVlcukE1Hn5E3JLApxav
p9nHlocyaGNJaJmoqEYvNSddm/yQCtKIB15WkUvoppS2+Ek5qi/4TOeTizGMPcRs
sCAfSEb6k7nJgzQazPwBz4bbL/fmKtBnI6c8dprVCmuaQvFJWR/dWYutIv/sA7Qt
CkhltfTUYtFSgii2KfbF5R1uunslrjo30STkWUu7k+Py5aZ6/FljK5RUZHYFmXAW
JbGcxBTMfn5MEm3lMeOj3Sf1SY/W/anSgiKTeOrJ/1xbmtMbBlh055tiXY1jzy/R
AMXOCXo9r9uX7Ck3Ms7uBG1LM6Hek1nB+IbAs7trZ9fka5iyQy9xNKq5WjYlRhlS
TptVaAL3k4FYRPNfT5ZYkvCC3ustemiR2Mj7JTJDxglbRWSL/Xbh2WHsvDYyONVu
8FTVvpzhNeGg4PMYRRK7EbNOv7XoK7rhi1/oyHh44YiXJtUXscWy2HKQRZtYvsds
o6mcUurSns6ZBFTl3hCT2Gb1OiTPQfh/BT7bYtmo7NIg36rATX2MjUlr2oVgC1Ww
vvi9mMSrUgVvHo+yZKZo7mDqTzzJRl/Y0OrxubzTA1UdtowxN35YkITLqr9Zv4N4
gynA9GzPu6dfl9JarPuWJ9983ec1Y8uxEXw+u+NS8TZgfBmmh7UD3sKRIRID5Ozi
+H3C1z+08P40LMUkzyvErCdatHuSqmF5OZ0LGSEq4U+caRNXgJo0lgVnw4EyAw/2
04/Zwdil/AqGovtU3v82+YI/S81JQxn0ViT8u74ak3Nj5iwz0sTX+Uf+E1Xeagdk
FS4SGMjVXQMUuf71FKTYfGjGX9L5J6MK/s4Dsdi76LjDz25COuLhKbVy+84PJiLk
6WYygDAD+uPZA8/MMhLcekz83bNABejIh+83tAI8Vno5Cg0w5LWmh40cNsK/FWSi
JnZB9WIurLM54X1pVxs9Gulsti4lEHzchy2wCUEqETo5/lFPsatj8pgU5YM08uV8
aOfdRtLGYmBBrFSVr5rQVcn1tZUcG9t1t02DB98qgkgwcazlQJFHy09KYUgjJmE8
La1neQ3pp9F0ziUVjCuiX+1qc10yrZY3GXtU0mmdTLydA+UVXXCnVS6IUbiNiSQV
4cXQtbF7N2+r/wLzUKj62hp7e8VR279MaQ2gQ2gK2+2Lwk4JxxmFLPAnyzz2mt5z
hR2gKYkR47MbZPUHUmOVSEfsemurgWumLh8/LZiljhc=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ClxM3U3CvmhQt3GxoUtlwHxgEhj5rFCy+9H5lYyn+Sa2QuMA5PmomP0fAjHjnymm
+Oo9iqhw/+p4qJ7tUfmH351XSVkhG7DqZRUrdV8R4qFhdlm1FAGGPmYkzq2Usy44
zbUJAe4yPoEuAW9U9t0TDeEsQ1x8hShyF2ld9m5mgKfZpafpSk1u7YPCK/+nARwa
vqQklhkTct2tw4O9NwRcvDyURTGzojmfiFvtpvJ7cvbXdbm5Spip/I5NeAMrapOl
g3eIZBaYA+9RtNBvZg3oH/riAcVoTVd8PqyGobvk6+Dvlb9IY4OZSIO6h41JwILq
mB9XpgXcpsTnFOwltb71Wg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 12192 )
`pragma protect data_block
Ce72smD53WKtfmIlxhUBsinfnPwy3ehDiYXj3e8YgowkRXCw8QNz+35c0LXEtOyX
QqbM8f/2/SRZTFfg6hR06cYRsM+jvQPOnkVh0tGT3xOU2bI/OfrPHcsmm7xPUbmx
SfeMSgfkyW7qSd2wMPFUMAyR2YIkw4VghtinHIxsX5DKCYuPXE/vCJNReCyRqCOh
OMRyTxQ5h9qjsXiPjor+Asluv907cPq2+MeBmBO658qE9z8UeNB3NL+58kVtZlVi
Ry0Vt2sjUvZ3JXs7YGAuI+x2VhqES5/YfL6rxW1GDkP7Z1f1fgnd6PbqG/f6TmDz
AiK2fHX2GuDSQG9NIydvwRII9QynyNFdGcympcMfmvdDULfJ13VKxuLjw6jEguhj
YRbfI++DE2znfE6Sdsxj/5EIuEf0oHiBPY5l9ucN6f1cgJi0IrS1oaKaKyAK6drc
PTX7yPcn6qDMEW0P+TZzTIJ9fMVP6U4Q3wAW9xDmRu8x8F136ixsjX8sotlZ1AWK
JHPwger3F79GPlROtg71glZp7E+d61fhMnP9aetpVokzcLBbpTh5+K9pkRv2cL0p
j0UtXwfOXGzJBQjbDkE7Hqv3SGveLa2O7L0N1UiouZEWpkOGqmfxrJ1M7V3naYGi
GMv05z8i5bQpDtFgekaIjcnLnQw8DcmoDi6Mik1ySe2nm/Cy8ZyBL+zM87Odi1sF
xIi/GigNiLtnQDmafEORrIw22PJvaot3EAEb/VOtsuWOD5bGQHYMWOZzDhKWZZnB
kFRDR3Oz6Tl6U+ewon5LNyY7fpm4+uSS3V/ZN+h7gaejZ9OIQWhH8SSewBbYI4lz
NzMTK8gBqHKmDYzBf3EW8QZBpV4+GffM7YTQNrZg4n8vxhaO3phb34C4jjIpPLoy
UxHyq4UY8GUeSZKcrM3d83Y2wIMgCNCuxbU1G6zpluDCZh0F0FndNVVmWXm5tiGr
IhlLpkIcNGA87G0grcimiQUiz09mpebPGpNwT7lvaJgEe8IJ4BhQwW+2wTWFnvsx
s0sTxCm1i/7oeLxjKYDqLdNeVREzaslRmKrC/jNof1CYtrWGN3Cft6/HypvyBren
1s7K8PYca2JVnr+9/B7Wt8AlL4d/w+xMiV0TvukPRjE9rLNB3XGMK1XsjE2wvS77
i4ywk18lSG9G4w9YWqptRgWr984FEroUEZd39rMrzTYizgg+ALitEyQuMzrsYxYZ
UcM63CD880209N/94uE9e+U2Q6WJ3+P+j84itMhohB0kxdqoOFr0iQtwfpdG8PdW
6LyGoVjfBXZ1+YJcszyAw8pKiHEHODJalrPpe1Pc0ku7uugBO8J67y9xLxvokdeP
y3wltV/HUwqx+ihStYUo7wx5XKfi3495fk9m3V228OhNXWotcewN/82G9rr0Q0Uv
9EkajatfGI+MbUBhxbC49C9/hQdgFDOInxd/FQ3FKKhI8qGBA/ehMxotNistVsgj
On28VgUG2rJVoq6fOZ2yNzClK/xWmmSSPoXidP1IpWcCNBkgVFkSz4O9fzXOQjKc
hrkq1S/M+I63VlkMWgx6vSfXUGgl4zC1NqZLpMTLjZtRA5Bc9sSCALkDYlAgBlyC
0Annh3I9UsLVFJQIJ9zPOFIdPlPbNwbTHaE5eiNVE6I4a8nXcPpUmxpaKA6IcBzs
wfC1+J75NkMIwWvleBpTc1hS2ATC4KbNzi1f2d8Wq4spQVwS2/hEG3rKO97uA+mo
UfGKCUm73Bom+EdE0/nFvi+RWpoST1kGIMXDXkb65UrFac/Y5RF98N69cIziANTn
F4+ezSAKylL6OiMbaKoNTR3WiiRoepVxphLjc0WdcgsI9Sqo5nXe0ODpJ8Q4BgNi
fNloLuaRA1Efhnbfb2UE1zNle/HalZ0zAX5stC9afE+rz3YnXF1quZxO5kVW6gow
p3P7LSX6fp3iekYaWXEnOkhDaN+nbZgaj0ETISFHTSMBy6G/4hFbxGD2J3//haLW
50aHgbvMwNSfqyDYuIVH2Bec2LTRX5HKh1lrJ+bdKNlAx6/BwvW6dEUCF62iFpTz
tbr8MB8b63yasSMq8OaMVWkTuhibTXu7XL5Yo5AYROfB83xQt/GXRmHK9uJscuJp
5He25MxuBFVTk65/3EUmb9Glt3FgRPZQIG8kXslD81YufeRpNYTnDdDXP0xbrzpd
U/CwdzJXrWEaU3ryfzjugEl3aoLn6NlMWAhamjhI+mut0t8vz0IHXv6rtETkPXr1
4qMr+isDatpzugscCPESlkhfj2P/B0HDP4jXFhcl2y7nKCIiJFFNScf+diq8mP2U
HiRbf8TivQK74Cw9sqBqwEnRWOsoL8d/6nhapBdWWe0zTP6QAUyGlRd3jBeC7pA/
wq9S/0GnVDcmdtnNFer4dutL6pRBaSM0h/q5ckXGtJ1xkl7Y0rhRLXIJMgmXr+k5
FF+Fb5MziwuBr8r/+Sx5yeq45/cE0QFTbKWgf9HaQa4tuHR38IUxCSmA+4aQvZHE
pUslL2ATQq8mrqa0ywFcYrKc/d7qzcZApJJOwE4DZvFTRZgAPaldh3nbVd4uMZbp
XE2Ov7+btvUvAD8tqdOAiUnBTtTO7sAiGRHsoL4kMlAmhVk+qJpq5l9jfZYMpaQ7
tmY11h31e1onUOU26+mxAJq/I0BEv6v1PBKJ5OEZ8dmS5urlIw3vy3dfzki3OMYf
BLwlNDEPEgVS+VWjjPUIbo95li/A2BTp16gbK6jqgqQ86h4yG8Sy6zC5zWlAhaUs
Avvtzifno1MYNS6LSEk8Lk5MyNmMnJ0DVSsthqqNh9QO5YOd93VtxHPh235j9vEu
SO2x90u/kzluExXLJ5PSwpnQO4N1eMRJD7cws+TI6EyL8ZiCzqH2cKo5QtovTLT5
dVIg5zuHcF2oQXljnzoJp6kcvLK/ljviMMU9lRB75xnxkMERkeg/RlC5Ld8V8uMK
4exJ0dGGAjTqz6CMDbY9APxr37i1ZskIrUl8W8jUzXg8aHaLe0sQU6cC0Hmo/nWU
Egbs+xTj9m7yGkIQ+aMZfMA0Vi+tyHyXBNzCoPRubI9Xo2RS9ze06jgZCoGDgG0v
gf4iNZG+sRMvWMzth3yujQgOLcOUzJeb8g0wooCWLewXwaCzWb14xZitzM6l6V/J
2R7cF7KPk6U6R9iQnzlw00FXRF1G89cGxNrae9Ec55f0UeJqht0+FRvJp9K5ATMt
O2oqaBu0YXJghLJBsgqlACzZmptPZ+iSk4QIQJoS/UYD557FwSzsqwij7OTdjczD
HH+mAg2s3FnN0J8cPia9ZVvTWmW57v7UcO7p2A19g7LuuyeYDQJ4Ra+3vU+aB0fB
/HODRKTyFa2Oic2UMfjzmWwX7xUnhj2KoZNpzG567LY9D8pDU3xaW7/LaqOqXmaT
DmYHpspJYryoyljKVDeWOQ8R2AX+XWx63HuWcHvHksK9J+e9R1vzNTUttuWmQoep
4hnezb7VDnGxKd0CjiQN4EIDNp8ret5xqRpkCjGsxiG9GKbq/3nYjM5NOcp2oMXX
djB6HDeaCJEcUIrTq9PfNqSh04lNHveeKOU/FL65Fl8JeKIk7+iXA4heYFepCka7
/baSzfCYQEg20gr1L2OCFdATCdHYo3hzvZOF7+Ia3qBlrpY+KsXwRJp+PENFij6r
+O7pY4DNs6hbR9uW6Tl4EtUD+d+zZauMO9V1L8U/AXxZhVUo27LjzK79WqHKqqbo
0K/1yVRf9nGeqUl3VX+UAPRe58g6MYdGKj7BAAcdUN+DnoOgYyMf5RaynsWbar0v
4w9mM9tvs2Q8JrzxuiZSk0/0zbN4s7rGLsLxvg1Q+mnUi2LtMjxvUw2KZAXhKF6D
Ow5ftcgpyktQtE5oUtPsLCyMaxk+VmxmUOA4AwQTlSiksbUFt20m3KxMZZ4o7iD0
4QgB4P4084Qrts2PvSbNOrCNtBzuEMGMlM4atttFZfeIHU/sxpmrg002QZZct/ph
Lc+OPOKf5lCYF/4AHq8aDinJ1IYpLAnrR7ScZO0XEZmJihIyNAEQH+sldVReWjEP
yvfLrUSrRgE0IYuaTLuaqZJHdAvS0Ebwm4wEcG7yUJsbbGDkOuDdNB9A5TfbshqT
cy++fP8NeE32ZI793wUpD4kjBubFFOLmkFvpaW234UzYJ+DaR/Xl1XTtuzh/qc75
5vyf859TS6K77Gt801vxXuKcgdb6S+LZEK88BcuGiKgV/QU1kRrxf7zKiTekyL39
Vn0xesom+W25aJrM9KQ8uoBvccLwnefMzNHDCHar8frqHUdyAntxaEXeX9ZxoaiB
MAe5m8BK7XnKj9Qc7X9g86snw+AY4+63C5XRAhgPp2t5ZK+5ZMT6SNq15isZB5TF
KlJpCXjCxBIA07XYifDPGCwyhcWRAqaJS3Ln1l/EPfbJDGdErWOmoK0bAunVrge1
eofh2yfRkiqDolcy9xRJjNsAMoQtUoc8Izd0DRrzFNtZ+IxpNL8ZSMTcQBvO/uXe
O5mm67L8k0I2KNy7I64+q2St4v2TnOlM18UDE4uCTqIkT+qi3p2gcFAz83+7fvHe
hJCRKRDAA9t0A2V4MOH51WsMPyGyYPazC8PFycqI3qBxVJD7gbfAxydeKm1fh4Uh
BgZUXbUOC6ifGGU1VpOhMn4fKNX21pWy13DRE+SE7CiF3xZ6HDEQLXc+IyTrdv8r
lEKHNlVCRLRyAjMcqzAvRSbAIzN+4gTGUcDx3HcaVK+Rh2CIl7BwXAP3EfHfs7S6
WK0p7ZjByZdMtsCqyFCuLt55bAVm/GCPgubCIGyR9iaCixaG7mgM4XEWRPj0UO4E
qaLUEhXGBsRrVLkowHe7vyAnHx7vOwXC4nEZUFRAS4LsArV2HyZ2X2CK6hGAnK2Y
sZlNXj34zT1AeHklxrfxFZJWgvKYzEKkpvypIg7+zzcayhaMcLJlRWicUywYdbb8
AjVVAb+x7brjTHVHMmw5zlqtamLIBxl8/UYuY389lf90MtIelSmU6rxzNWZSS0B0
FYYcO47vQMlq012z9T6QClS+EAIsad/obsSZylI+YVvWm09puSPZawORjgp+5BbH
YyesjswnY1jmT58fLNZaKYZw4vB2RYmGU348vWnfuj4iBqJol6WZ2Q+SCGehF1Ze
UBeA0pCf0vf6chRqRJle7bIix9E3oQVdjKHCrjzkyw1y9ETgCHJ4eBvtJ5R1DxJa
+E2LorpDFbTMD0Ewm9sNgwWAOP8GnDSpva7wTtF1SHveiyBvzMtJjgBgDWwAWYNx
A2B5IS0Hz5HcOFZvgkkI9Np5pRLi9VJg/iX4WbN0BY+uDnr3llrdL5YdvmsqiRYo
5BEUJFVgEhzxmbkUBKIwEgqXKGj0RicyD1NusVK3nNQ/8B+aCkq8kdi3KpLK+JaL
5Tuc5p/39qxfA/9giDPLTAaK7DM7mIDokSA0r/uGEmKlzba1Nazg3v5m6EsTVR8c
rOIpIbkoFFjr73SKmE079v8kirW96pvu3IdP+A8tY6I3zQKwifIu4N2eHkf+6k8n
TqHeWZXjYbvYaDDsI6cglweXJUURj0dN0pAblyhbTeh79FwrTV8+KbgUGjW54VWL
zwuyrE8MvhrD1oxNJzJpVAijc5BFIoZ4+4utiiMwbGgf5l6O5XvRAzWmuHkA6HHu
HjurP+w8HqO3bYKT68Pv1svbBJ4X9mio3VXB3EtHuC0GRSUxHonM34xPixCa5X6B
QRofwOwWFWXq3eOFmvpD3NwS79jo1I6+0RGC0ekBHs3bKwTwQvQloO6NTjE5KZea
XU6DoaqIuedVVjUN2PsKYYZ1Scu1XwDDepmA4R7R38cvqqw1yMg6G1ekWvD8h6tc
obz9EgqDdL3ptCI3FhGzJ2L6uS2+iyuy5sOgl2CH3Grt21ajJLz5UEWbCMiVGv82
zzAx4qDwbdKHtR9v6t1VSyZmpzNrhjFm/G/DXBvZOMh9GyWFq97ThJz+cmSSkRLH
Abblxuz+O+K+AN9XyQIJ1nd6bd6TckrwfWyedX5XxGdR9ula6KHofQOxkfBbOOZJ
3KKFVYxPJPiiXwanUOjktmBwU+8b75cGzgs14/rXROVq1yLIv06Jep1NtxQecpXI
ND73e+bkZlAyObgfTSE9sXcKGaXdCW0fIfXHsuofhjlsrwv2HJIBDemrzqV+Ykql
vwullvmz24UjFllte691Tq8zazJUCjZoOEq7qtvfF0zOckf0csiZbsPVWPNZNwSe
LmsHHAKY/w88kB/sSIAQB8Y86Ng0Wq2GOFJrY8q0bki9k9YEFasMwsl8nkdlbyG5
1yPceYwnyQpVoHVPTFD7r6JfqvJ1hrKw8j6afoqWA9kNR5nrEqS6HZimhCYYPCa8
LahWnHJoUhAokkwiP3X6A2ezvQRjdtPhVE3XFb0iIbAhcjJK7Rv+C3b1u8Doye1N
7YHc0V5CFW2QjsRgMmn3JeYgA6wSLPig6iT2rHMsJBMhrI+rC+aNbkGHf335gUMA
Q+eGi3WAjb4hp+LZjkv0ra3ejqKu6CYubaqIl6W3iHaGwNeeFttTr8Fb0j+QGK0l
n2wVp8WWA1yxz2G8YPYRM3XmnwJ+OCOFWeP4+A7atDNaZZMUtIcNJ8aEwPNVS+E7
Gy2IHRM5HrlTVvmSbh5+6V16SfQFF/djO+QdL6CveNnfAxr+OpkbT+lpHk2QDatf
+JYyGCj1ifM7oRCWBKSGpRnz+ey8peyxlMMrQs9bd3JoJ8KSDHAwmRuxEEHwVogk
V7PtQnc6eOZP9fxst7bTJh8ELuIap+iRjkDayi6UK3nzK+rccmOGB22oaztWUR+0
EzDYMo83P7PQRVFc29daASrtBcxuIOa4w0a0zUDQSKM2ZFIQrDILSMqAA9nxrFrL
HF3PbGHfAx00y5GS28rzRq3AlNZfVZuZSaKZjfG5IE8NMj1/XUThqmzTQZC42/jY
e9mJKxvWSWrBxVKj/2oQL1VIK4UgHRFhgUquH1F2e5FknaccWyiRfsS0pLqOjLBl
N5/+SdoFSM92X73EmY2+w5wk81vVauwEwEcXogXlcnNEHQI+dbJGqbIvB89nn7YC
k1FMyfiAHIBnB6AtuAWeKDTnRhdyuR5RDgxzBxyGHKz3jkSGRhxOoo6wdzAcN5Mm
rCo1KoWRKXp+Y6zVC/9VLk8tRyfsGB+OTeRiPXyViaGtRDqx6cdm/zBlQL9/AtXB
P6C779LaRTdyoEATWgPcPUPYv78P7MwxHtMd8CrJUzEv8Pb9W1iCP2l8a09GDCkS
GRLIoXpX3KpEzGSjMfk0/KLe5sJEb2n030A58Yj+hanbjLLbtPNuLMz/IMeo1y71
u+gGMTNWJImr1mfUO+imzogscwh0jScfKhMPAkPkk0mqT89Rh1L0YAVbgRGpUxyG
fqp0eJCCA/g4+9AfN8Hig8JV9ynqgAoVxjUwPSeJJL9o38kkx3zRKv/BnDKkU8q8
H7eQhJqdPspIL6oX2vbX31OK8V5kwFzpurH1dUv8AnaD6lf71RR+Mb8QFs11zkCY
76N2YVEGstf2+44ZKRokjmvhJJb0ybBmKGdZjK+4RBW/bYncc0JyWyGld3TEA7XJ
upAOwLOMGR0cFE2/zYiau0GuaokniolfXjJxX4XctrK5O9E4QraJSDQLKba3DqGP
ThAmIXHGt+92N+rJmNBkQGl1xEA2Q0Vn8EISHQyDH8wpgFca49zG48pRnIe4OPV7
D24i1t5JJbvJiW9GkekCM+zHMrUvP2MG8A/Uj8vGh20wh7rHcSSi9cckk5qgpXpG
/Gn1kOjiKmTv4CSZHgS2BOjecPTjrH8MoI0t0BtadNNSfLV5rKW+K4ip1NnHii4l
2CXjuY85f4R2MJWc0iVTyLvyrrT0evSQp9YqHDTAJQWqg+uhpnkLFMlojU6KRZXw
/zDgu5Gt3/SjCu8HLB/x93psbCsb6sRHZKOHOKloFb7Nw12t41PRqOaYAgx2hK+e
bRjkwrkyWDFE6RD+HkZFkYTYgzCOQPrbkh4Opm46Slm0WV/H9SrzKv3RPvL3/HSO
iJ/a4lbI51I0/IhMCb+7psOq5anR1XPvHvVb7kpEWWLJb63eORXaFkrnYotpcfia
DK8c9lXpovFC/W3CGaWj3kdCsQwWpYARIcAX6F7uo8OVUDqbJJbnJl6C4GbyzNLx
SlYIeEqJd01w+TUefNhokOlucHX/rcbAAtiuw4oAB+myO/d+SkJK/93Z5AVw1ZG5
gZWD0p5gb3wQJP/lY1B5pr+RHiS9Lu+2XVO77ECS81vcSmnOzDEOb2RfYw1p70Se
Tk/lBYJLHJS5WjQ/3J3p+mAaH5+g8m8sG6dW/YUvX4LgmmaDrzvZNosrtIAZg6+Q
kuKEDSxcebcxlGDY04OOZTqSsGsMEAjFWDohLyoZCy5x9QOB+Wj6NEyTPZpv/ZW9
e5C8Va1paeX7dUBD6EdBMmGETU63skwRUuhj8U0xiuIFbfx5xpPeK3DrLp/fx7XR
gm2gJipB6tCM8aS9dilyQ5LhdC97x+QV8Vs8TNGbsn5qz435RuQ0AJbvTr2j+vQH
irWQwGlq6Sd//yOuOU5RaPd+JTFnGMvpsyG8NX9WyiBJ6nmlY+iD0ZFLCdCou3Lt
tHxHWOb3vXkz6JzYDS3EBwGpaL033IzL9kl8+e3wf2w977/Khp0J3BMrtw3CM6Gw
quwhpddAGLw8Ajj+91tDid2CFSoWtbuTeCdUmmWYireR3VDKRPqyVk7Hq6XlzP0j
IKFmb/pJuejlPhzO7H8n1+TrxAkQFEgGKDntX63TZsccTVcrx4xHCSXD+T5IpQGm
nH2+rfvl0AOYJoAsQzIkbdwsNa4PJ9SkQEevScIwWusn+rsreF5qfbn8olPLhj9+
yubQ1xf1eDgwIDbbWHK0HkmZ/qySMhsqmWR5t8EV88ItKVN8dZpKTb06upQPXpds
AnmP+EUcorM4wJLw6JzfWxCGZnvYdIxSfVQz1GHus5HEX2I2kD3jRiGVMpEJTfZq
w2EdpmqoAhm2txQvZ4JLiMfAebUwzLOtel98aiBu7otmJSe0kITyYRrDN3ts7G/J
tK4EpZb51rV8Nr5xjk70UFcs5G5FcGRVsQcKI9xtjbeED2WGUErIOAZhVcUQ9saB
41ULFQ4bIA6xdMz7DcHDSl/TgpAVFjrHWAo7wpgQcNTlTMrksL1zYqr2TUmtFeXQ
Yugjhrw6qjQ7Ira5IX928a9L6Zj0na/jR+GnG/WatqKbsuN+7g4wVwuuW3c08yJ9
V1YI+X/Sa7uQhPcZ/LV0Fi2E2SrXk8GWN+ZVJRLt/AGlE17dJfGW+uqkNyngs+x5
YZZ/kFlJuJKoxnj3XqUmlqr0Usv4spE9HSrSBU/lsioTtloHrHty8cDPte8NeQGo
20QH+F45AJft/Aff97hKx5GgL1md8IxfUEWk2zusbm6HjJgmMnUmjFt3FLkqzfMi
F551aDIpA9/FCf7gFTjS1eZ2PxVt0QmY1I22XovXSNDFD2E6EiTmu7ZwHendBzHB
e4PUXe71A32QS7Pbl3pKCvIq8X5C8ceZFM2zHnerogtAaCFvvrXJ6ZIw2E8BkXGT
RuK+7fgPt+4UbeyTPHsSwydFLJUGgqDvuew22x9dcGl6xHM3rMrNtalAWuAtjlry
cFpLshS49je4Wsw8/lg8bEIiAn9Pyz6cCQNMklgMSMnrgI21Ir0DQb3xqiPjHlXB
sgOIVpIKX09xZFX5fxdHicsaTQX7ne//sGx16tFApJOLelh6Jf+Yn2BGTH7Zi272
kvuU5a7rVryb2A/rO2W2fu35rOK0EhEc2kQ79ioxhq6YuwyYBFVs+/DIWwb5Tsv7
NYXabjroFLOiSoXSGkqwLVMLaSX0D7H7774CJpGhpaJsakOGOVVtce0zKsD5mjM8
KKtbpj0MjxU8fqp4qwMojfJP78+ugyg6avGZQiX4LSQUM9GUxf3oGftyhV6Oo2nS
Vu6Je9jfaYAAA3ipXw0YiwxXCleiMtwb9F6Re1PAq3jOoAzeli+oBbUeBXMqPeW3
Kkf3C4PwvgBUsdtdxOgK/QPVELEN40CIvGHjFDbe7h1oTXwIyo/f+pPxpj5m6NVK
AH9md4n59iS7yVz82K36SoXLcO3DRNlsBCCzcShAusFPUK8S7ViYVY2RrMqHXTFa
IX8O2zdFs8DqE7fyi3ENVLxHxwKsLcPZDvTKw+XtPbMNWoLJnxa/5fpt9QR+RIJ1
5vjUAiV/9ecTnucfUDzd3OHtz4+ljyuaFg4qzIVgNKobzS+gebHtHuXB84NxUbcf
J9yQmnrSqBgVd3G5vurWNnlowP/es2u+X8FyCjPcvCA/1vhoTjOTmfX4KZNQw5iJ
ArVk/joSU3urZzGQNcWIbQm7m7E4FVjllyu7XEM5F5QOM/Rm8z4aH/jnbYcYEAGq
itEHEJdBvi7QThBpRMceNEneQ16s6+mOW1rFpEm6RkyVb0dzojFip7SqDYziy2Gl
bCxt2WodL0o7mS2r4vf4Azpbv8FAAxJnXXMBqoQPFzEmcRV20DbeUM2QqY4oPNy8
h/grBsahQnrDZarpKreimoytYn447LpgOu9E0oy/2pKWg8AHZzytDC9Ye6uHGfdJ
WRH5TxgwlZVI/xQQK0nkPFbMRM9/u4Cbau9TPlTC/v0mYUhHeint+dZ7UTaGQMGN
5NPtLH8cRRrFIKYj7k12Bpefa0Dn83FJYiml1tf33hZUHEOBlSshEmFRU/KIOUTF
Pgn2HyipTSJ5+S+vv5hit4LfbD1gZH8aC0Yz9tA+OURgeF+DAk0ZqvBhysS/PwUT
FzSdCWB3jnIrqFv8ZXSoq5qwiGO+pqKrmP85mVTExfdztLEgzlgzxe3uCos9N35C
c5e3feMxcmK4eyZbkRtZz27Q6zL+nBNIQs/gi4QsxJyW8OBXw2Dt9o781ed2p2RM
4jcrbKakR+i3Zx0GITJUYnX91V7ahMKP9kDxOmAJGo3lJC7jNitwdaOJbL/KKwLR
etCx9q4ho+uFMxBzIkAHREg/goa0GLfJ6NBIAVFLWs/N8KduIMVG2X0atEEdPeOg
DAKphAKFHIy6Qq/H8Y/DnrS7SB8xVkG+2CvYwfcGCUmysZdZvodQnRywdxrYbnRe
HXQBKVu5rvrQ0171DyC0p47yALRTVgLaTS4IhKT+cGs67TD1BQnyEaM40GbwFmuq
eK4uh26CbKClE2vL/JKGXYI4G5+CpfkliXpiooOU9IjUJ1M51oIx/KfV8sCnjfLE
KUjsM/GosC+nxFooGzeMgFy7oobUQat/8hgP4b+gFssBJRGEZfqRTodR1vY1wRJC
LlS93Sh+SGKlEVx0Ya/ujwRZus4b2TEdV9GMF9NkYqsN0AiJSAk4zG3Vefx8kQF6
kwyw9YXx+lPCI4IJfEdlTh2VcwnJu9Z9G3FbLkp2WA2NnYLX+dVRH7bwBebSD4Xz
loVUfhdm8mr4Kb53LJs8O13t6HT0+k4o38KLiFjQwVenkeh9Qi8zRQOspERMsaZo
3aG/UoTNbwOJf0vlcIqDkvccndRZaDG1yewXQjpLki4NS3mx+XfUyYNtvo+OKdiz
hMQSTd6HBj5Ez0ZbT+g1D9BbfEjvMRy3S01KGwjnANToHPk9nsaNev//YikKHtWN
Avad1IQl5V47oLwjp5CJSEd3oPQAwHmYDZ8LYm2LvSvRQO6nLpzS4d+K19S/9RvL
OInVBavsXREbM6hrnOl+ibp/CfDGJXIRrK4vPRZyWNhRUz8W7jzSBoV60nTk4qO+
KLLvy0LoQg5OiXFPelpTd9LyZxVqH/W/AJeSaq5t3G7k2VGek2+QzvKsAp9McWzZ
7xia+nqjiEeCfJAkMpL3uDBYyK7nECFDKrGaG8r8cp5TzApHJy32SDIH/CVwu/2M
6jHMziPu79H5geJw8Q18vRKFUQcirtjmIWnmTZVPmswxFii1yzL2UKH+kw0AOFTl
BHFJWKnZbyBjr4+8/UaxlDV+OTgngbqXJg6cOOas10aPQ42MkL0j/BDrQXVqxlg7
Um24QJABsO+lBZfYsCzl5MvO+/9hGpA93fJNpaPsRweMDpTlsgChXF7yFb1lTZQS
t0wdgBBOMRuh337/ahO1Q1fQ+9HpxeSR+dhx+Rt/Gg0rEpqBfTyekNNAL8d5rFeA
OEUNDVhX7haXTq8Xe9G9dLhj16aGo79bMUPKta5apmFlDBzHJRPKNRh/IJcVxKZS
jIlweb1uB6o+zIsSH2P7+vSB0e+6uzk7ciNziEFEnOyoVrC6lInlsH97bKBG48bw
DVOo+ayiMpJDU3wzjE/O8fgSbWH+h5/owe9c1OXsXSghIM+iMmboAkFIXXFBM8DA
aLcXNa73iQDWGXRjHSozbuejYicUFLpv7mcIG0jkCowV15uvgJ/ZmbJHkbkV0Iok
mC6kQHCpfTySJETVH66IzSWXbhiXCyX+L7rFChTnK1Bc6qCKQ054jnudSh25ltGB
zyZqUuYh5zfMDPXOVlReEFYLAaZpsa2ZDS9zjF/OTaupP0NlX/OdyID2bsByOMvu
O3LpWcpVBwadPX1QdtN3KBEqCosF7o9uaaroQLOeWCrXSiP4eEnTobn07wlcvX40
ILEQeFEXvMMTY1/sjquygbHIePyLb/j8rwnG0n8p+uiJXJPoZ2vgWBoPbZWPwt05
e86r5DPkHWg4usoTzH3x3So6Du+l9eXADPdhJ5ks/2J7gVZmzjeoI8jxY5FFoawj
i6GsykNWymUYjQ0tfIKRbEVcwEt5+SmhlxlpXsuiuT+2aAXkON7HE5yaB/XfSJrO
82XKZ80kwIADA8v4gawIDNY/ZlkJnNDjjmjal3xNRGn4S+7dw16ebzsJFRYJIZm8
Nny8TrAHFheLdeiELbF0tXq2C7DgV6Lw6vTBr+zjxwmsEmgIeKy295ntdWe5a4VI
aXM0TVFS9lRfDGhy87/SAMe8mAi2Ti5UfI5thDrBhjltK7Kc7zNS5R4yYeEme5J1
ofDFa3K7ng+t5bBlygqD2ELKbgK+eMExFGL+SWYtzBlQNmgfFIfHMEhXQju7sm3b
64rZdHtwzU+H84NHiGkHBURPbC5SJJBzVaHY1q6zPqDghtxBnpfsemRSlcd5jTiG
160bOze9rTo2oJf2c7sFSoU0Zt3vRzTfaSZk5G1LGwAqypd4+8gFL1KLeLfOVJ7H
llIxXLJLCOcDyqhamjUHY00AOVCLNAp/YG8Mk09mKdL+TmvbpN/d8P8d5Hea4wak
5lszuhmOfJ5jdcXdU38oUp9WV9+HC0r0k0Izt5WmHuPCLlgJyB4FQchpfveewbD/
Tv5mP0NpzNoxPGknwdm4YJGcX6LhThViNPm5VoGn4eM0Rgxssg56byK0AoBmWZ+d
ZeJErX45q343T5rr0siByg2HrD9uwx7EIM1aIZCX92WXQwYYH3pq+U1ibse6glD4
E+WhTLGcBwhVLWD+IXX2DOW86HriVLrShokACwSk6HVz4ArGfGDI1ZIjT6wf3mDX
htIIJmjPj3fz6bIVLQeL4LvYsSrtJo0nY+ggmQoBjdybxYAH+XfdvtZ7w0XxIRwd
hfDA02Faw/+Bqw0hLTWRkCGhfEKBYih8q8aH1CyhpiJNY17E5PeULdTk0cgfaogq
K8qyVy1zyYkmVSC6MvkA5IowPH1CRgcdf+N1zoss4OrtUKy26Jkeo2d6sZtNb5B9
5ykPnj+EjLnwdJJnNcJXuj9WuBaru6BXjEILNr9ZNcBbYuZPCtDds8EAbvpJI8b8
CDv6SvLw4qc2WG8Nx6ZIlBaaB/T4t7GyOTrRG1vLgZ/knQP5n8ntZBDZeNpMexGp
EOLJkaqgDCrMKRtFJUIqWfRRTcnPK3oIcjhZ4otvR9BJXm0YMg0cY7sSi0sKJXB1
A8/LpxGsA5mrPK7hhOkqnBX8HQ+XKBzCIsQBERfSpyug+YfAUuNU4j+MmyCjBCd0
sKhWWM03B7sKb8CJwyu/3qiPEPn3Dhl2NPJYzXs01OIQFNuGIfx+5Iz1Nkxg0BdU
B7aeeRc3y0l7sWSePIYoc9BIE+ptWwvVpEe8jddhompHEAh+TVBs2m/fzN+GfWVL
m6Qn5G0WbrmPyHjfzF+WH1UDZSpFYmSYCFeTtbVgbBJgeiP/JTZxFML+zrHzYE99
fgtHUs5c9VF8gbgUSUJSktQ5oAoSk1xyG3102jCkvKCxGXBUQjCQRi+mPf+6nzfW
XZQ2syeFtQQR+HnG9/rWTSG6g+NFnLzLkfKJ0DrnHOr3Gs/qTcxIKnvzeIKriPq3
we7CpQcrJtAkRhQ3+jL8yTdo0QFfE4/f1kNWBvPRaI6ki1E1v5mHbcSgisMa4MwK
UH0fHBnjcDienpZph5GK8CCBDAryO+fC/lYifAELhqaC+/3nbLiEgucDRQLcfZRN
LAkCU4E2bEXDBJG9Jv+n0JcrTDZz5YtQtJEj+1LNHbEd2o9ea9gyDoDvaEFahe9D
5Ia6WPLbkC4TGZPPqJmdizhucch98BdJwQzvvgjoxyihl9xS6OiDtQNGbm56DmG3
nGyEw9FeuJ2DQCYNoUdfEqC1wr6NhpMnzlWONOZUISbtmm/EypFw7CXdwys7rJVw
HVa0BH191b5drSqbfWRssmE9/JZYKrUXfHLpBGHAGkmN9SY6P5V/7IV/KXq0UoN/
ORsiA/KaXlW5CmwimbYmFtSeEENOFs4tt3V54M9K+CvhMBI+iZsXYVozaiew41Eg
5CItif/TCchLkMiUleRF6ZV2/6wKU84iDYgVI7+8B31gNhYKpgOO66VoWmpLloTw
Uo4AoE0xl7Crglyj89oYca6xn/KyfYdY0N76tNhPP0SRR+Ts1ckUSekJhutMemUH
koflidTO8p76gzzGmIFe6ocqNw1vXYMGOGlldQmh0kQhzX3tlnneM+5rM+VIDOlc
IJTS8r85JYarDwC2izl5TldI/uyOxKzfqu4vYeXrsYnEOiaGnklvBvTHNkBUrM8z
ZUHrzmjOv7rxPgzCw1vgxGNPc9sdKZy4eT7uR1WBkFe1c83fDhwRChLOW9MV5e5E
9mhywCJ78I1lQHhmu82AlfooerI7+nUgr8NKiA5Y0rmJJ+ls5Iy+kmlYJkbH8XMF
2aDT1MDn+rZOf/6v3butnv9VvLGCeUQNE1oyEb5GTGgVdVA2lJKwteBItFIut/7D
96TUaCMhjyw83szAHPUPDvP/FGNy903yZM/RO4/gND1QBwC0/+Rhpi0GAxDBlZvb
OLseMgb4C4fM9gQSW7Xr1FnwxzmXPCWxkAM7Pbw0+bCHTCGAgqv4CrRR6i1jl+1V
JBfFWKLepRXMVtZBtVK3fxEwzxkwTSZySzX5vz6GWSEZMQUPYecBQV/GevITQZe7
kSkQjjz5tSnw1/Llu21jn3dgN57AzkU/fS6yfiavP5C+44NNBMLFd0PkAYaqsahy
pXTQT7paAGP9VrhWM22qC6cQqZmtAowiLtAjbzvu/irl+lz2e+74swNBeiOQTJlu
1y+LuCljOM3UyFLT5wByd77VlmwXolLyz5xl0+kwZlYwnWcwAGz3OEb5biujXEjF
zuu2i20I0Jhj2qKEJj9O4rav/obe3lwGV2Hzt8VVdms0ispG1aMN5cYvXJubURBW
N9T4Ip8+zrfvMFl9pJR+05nDXMQm5nc0YS5i2h67wS1KBOIYFhPSfSK14U8Uv5gI
/x4Htrw6leEpV1vZu0rdyQ5CGTOYr5O0XdBUrLxYCCcQ5QNfO49Qel1xuv5noK/i
NgcFv7aLIpMgrmVn2ll7rmN/CgJMdl5gycnCZQe1NBy+GnIELmUZQoV6MU057pz5
wj7QY2UqUeNENhrm4Vojz7WreMXDl7HENK9p5lyPuaA9hu5xS82qzaJb/ptRt/mR
YH/gCoApXxpsTd27TXXo1As1UaNhD+5VqGinZfQ7aeB9eo3RpHKni+sMyA5d8u7x
0eN+W+PIZ3oV4uX3e7cQmifffDiKXnxOW/3Luq+6ZN5siNE1pGz7KU32Iho2877N
QBeDjZBhcMDOfATq5ylYITi3LQFtU4AkiOiL76tolF2UgFHahFZWv+jOwR85sdw8
UMKvwUOtKN2vIjKN43fznFQ5cIaKJ++6y8OmW9IoIylLnkBwLXRgJqeHpa4qLT4T
Vs3HSXY/n/V/Kh4+ykn+s8LqahR5lPZ1OL5qXB7WUte2Yn/4hDnVnLv7fHKniggG
aUkxF4TJvEzckhvqS4G/GxwLfkK/6gCT1f89jULOwT85TJZ08KvfL8l6jVDo22Ee
YXzSfMX3aIR140lOQOIMHVVdvz2H1xFA5KJXjaYmtXkKhpuLfQ0RN1JDDGiW9zFT
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
axLrfFbKKfshbFa5EWQkhYHIIPYXAz59nmcrTwpud9irSXjAb28ST+NilztXaORd
toTNwPzuN+0YQM9D2CB6QpU1h07XOFrJfsprJ9M/yS1Hwg5Yi04/1mcZcVJl35yc
ZEe+YdJGMT6RB1ZhqTMP7YIOv4S9q+tiPMUXHJfVJzpd5HpMKTE8udC+Ps5eG108
MbhRuoBLdQ+30QESsG5LILqNfAi+RKu+nROFygw50ccD/ZcNtxcM1HrTeAPID1B+
O/udgpBRlVaXtJHe029mrHglWj9iOFNQOAmaA17FSQfYZYEOU0fT7tQvYlCjAAq4
h2Q1grPHkErAzel60kZO4g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2720 )
`pragma protect data_block
RuogQVnjbi2ka4Apt4TzxXgTU80Qf2sEbEFmYq5gvvL51umzy3nBsaPHpuKa6RsE
JocatatOSGFA6wiay/UpC/4/0fniV9cbETfQxT77k6A8eJOaOCFv6zDXdYdpG+0x
u322oct6zURWjN4LzWBTseg5IapZ36djOqm8c9OpSiSjkAfSIuDGZZ8uTSefebX1
f0mSLhhBg0nPQqTooO5aSW49a/0X+LUln04tzgDZZi6zRrfzUMa9SalZ7agDgYDk
eyJLMnYh8VFq5k0/COjiWgFgvBRgs4T68Ww79MWdTrjLT7Zb6GySFkAYUwTZFlQk
zmOHoOCwyG7WmiOnOKlnSXncB9zZwPw2ruc8tN1Q7kdSBU/EsUfKk2nSl6sMUB86
vfTXmMpZdsYAWenrf2paIvZ0GxwNDLowFuFyigY5+c1v06pblx+nVK7RPOiji0+W
juFNcfY48T7q4HuR5C4FGdt/DBIX3OYXDScIUnE99/ZTRxMP+L1UtsKbBkQOxdMq
krLf8pp7fFRkd2r5Gd8BgIjAvVH6PA7yPU6AXKsYEf+O5hgrT7qt4+mMz5y1LUiF
gjkEJ9fNbPuMLEvCHhRI5N4UcJsaTfDd8dFf0hr2rURnIoiKljDNpMEgpLxikLKq
V5KeA1UpeVontKE2JSVwA5HVoWYD/Br0oBbg3syePst9o6MKDt+aKCZBsYHAut9g
s7oxnY0Q2I2j4RS4K9ghH4++mwvirrgn+3IAkfbB4XBSygP6oieAMyEdAVPNVdLY
vKjcSpQ6jluopC79HLfHTMP3F3acQIvYz5p8KgpaauoefPT5/yNLayLWpug4E5u3
1FbraK8z2A44kT2SjnhWbzwONiMNG+5ZiPddgwXR4Cf1BWk7rZIt7uMCxJQc5OuA
5xCva7Ggao8JsKCTxnW2ErJkIjpuNNBeZ4/V8wVeY4e08f7R3VBJLQziIytr0srP
HkU0sjvC/pvU8/l1uLhcZBs7zu84mXdMErI5owTAoS0M7Bq53uCxPcbYnfif+p96
pJzfEOFzRcM8DrrAKN72/aAAm0WQhvvhnbTsdPOXf0vdKr6nITUG87pDx/HRrdbJ
hEA87APqypCgYQs/XPiAjwqX7png/jydEFp8RyDegSUG7/AlnhQJIwt+awYv8LB5
qTliHehoMbgQPcz3w5CoGX0PS5oXM6/s7XqAnwdpbWhBOckVd6TDOxZ+FxI+Jkyn
9VgDwGm57neBjIG0p+DuNHz2yoUxwJPmXtnLkwzLvPBbTTmdV3ftv8AlF1/Xuu9r
SxqJL66CWmyT9ofaF8gV45I2Y5CntRCUUgqczNEfC7j+odL3eudNL/AjSbO/0eiY
Ru8FRKJqjwAgC6c8PoVD14if8yWW9OXR2CbsKK9zmUa6+Kwrm+k8FW39vyT1DTl1
HQJsvEED0y4LAj+yhnMEp4BZjRAsvifKrvqNOT56BZHV9PAItxKMlOW/F6rjwKdu
nWeDm1MEdKIOzhu1CxbVwf2lTcoqKi8HS+YJbbt2ydMvdd/N06aUsQxrcF1+oTYV
oeDBSP7dE7bF1UEUofAGwdyiCT625DReUyi945yFJQOawHDjO9UzpimWfItnTEmh
nIFLnixSY2fXg5sWBayudGfYIapmfbstzCqkLkVFviGtPM707v7w9x62gXJYdXzv
s0HFAXsSyLd6pohyoCQrI7jIWfDo/fYhE77pkfdUW0Sgznr+ODPGSYDXc36sSdEH
GMTj7kK7cj0GKmkLoKfDnCvvjbIzg+07UI2h7DQEcgrLfl/jrm3y8yHK893jfg3v
+E3rH4HOzHVRVAzzaNhKMtoSE0gHwOfocXLGjOYWzNeEfXNtBRBBpc2oi5CVVb5g
4Cph7Nx9lOs6HDP9VhbtUxWU8IwbCMQdDIxvd/QkICtumQkA0e3eC6vxMnGOOnwi
3oQBJiXoYp0VmAOkRCXrpBDDUbIOmkZGjXlmLbopOOK+2G0dDT5EBmD4b7nNhpWR
Y3k51DUsQu+JVF92J1y/0OIbRGwkFHrdE+IjnYJT/E1N19cm6MAz3/JCL8sa6Kpq
U2l61mFGSC7cQB0ow5D4w05od1Hs1qs0mZv648z5AjxY3o7cTWwrLLZSaRFMyGPt
3Acd94PaR59zJuAG+Q1DiBgAWyULsxteFYBEu6h/EPfFS8KfOF03VgU9dtOl7S8Z
DRwfOdZMdeKE4ly/S8t0gcfjnZNxasXQ542oY9Fb8rFBwbiFcKBvFAUMLvy/RpSA
yMXI/e2ppWS6jU8Smve/b3+OUR+SdTLp90DEfH3CS82qY4wOS+4lWVqj3xUmegxs
ehX8ztYxaBGHBqKRzKDyJgoKOKLEWAdqhl2sXs4qBxEUEAtnov47lzyhENvskxik
auZKDdupY6U3wiRXMWo0I7gMKVg3MypCGSheRNIoIxAChQB5nnm9hlrZOxB9oNYI
rkjwdmGB7Ru/kYFEq50I6p72hDSbslMP1AOEAhll5lLpPJLShii9rhGkHO8ucJPq
DEp/J2FRvVcxphkG6bke9d3i/pCVgXy2b36C37LzfmXwP3QzbPTyOLP4qSQsSR8q
aEcCEu/Ow+ZVUy3k/VVyRhv023TlQ45MsTRCJ5IAM1Wo5Sq6L/8i02LvumZr0GVL
6g1oUmU4bCOmm1ca26A7xGKWD4arFGZRx60L0m+YGEYjH7SkolBgQFqGcSPpJ+n2
Ydc118j3dxRUDV/Fy7UtQj1XMGGU76Lf8d44fz60SFkGdKnaPDnpMM5p+CFeLaDg
l0kl2/maXYIPEBjr8Dnxjb4gQOU9Hf8zTVcgtSJgjQrEfoCB53oW8/Ptp4b7ht0T
aJHgSGGuyX/yWfSLThs6CNeM25fW0az7zFvlkCaikNXBNXDg9a3mc4w840XpXCwy
qQuGy19vrzfAWwQyMUWPhmAB8DRpznbzVKFQbwX/ybi8hBl1P7AHoc1v36rsHWRz
Miji0G0BWxrrb70dWNIIsBRcgFNc2nkBuBF8unsL2+b/uK7glIhxDlzkpQToT3FR
Qg1esAnhgq5vKLN3yTxPe7etFLiPXUZyRDu5c2Wko5OcEAjjvAPjyn69PT9YD6Ii
42LBq5yoyg20iC2zQGDA7PkFAJ4Ab2r32Q7oYPwiPJI7TVmwCkuOXIb+joolSIif
Z28tyHm5mdLhZjU8cQdVWzrvd3QMPGJXdUt06QtlTbVw/uvjTE/QFh0wTuS0qSak
kUABxe6q3mfrsXX4DNL9DJUpCXxdnWDKgYvI58SwpSWtTtAVTsMaJTW93v1+pZ/+
H97yQ3U5YW/jnapB6gO+6PZMbK2hoPL9EDVLkgOFYQjmaIL2i+WHTNFvh6AHJv3O
2WLWpHqX9X1pgeqKMCZIvfH3PJjvhTwe3zvrWQqvT3y5OMHQ56evQPVYnW3NAxzl
Bo1+P+FarthiFcBsO8tZOwCe/aPewWyOgWCjyfpUlXAVfUMhWfeX3gBLbjt6CYdH
ZHHaQhOG59s718ZlHmvFqVxl8hz1ny3ypEJmENbB3UlBnqlbJVtOiPsPwPTZLNOy
BgKaoGOv9tKUZ8FZtBuNpjEYzhE7NDXodSqMtd5tQBGA1ljuToVTIQkLFL7k8e0q
rQGiZmnUvqY0FPsCrXiRTdgr5q1rrr5l4e1daVdUe6s=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cM/V82nybE8c/fc6khVCkvUwEECgSXvhr4/RPwG1oR9u31FdHY+enMh1kmXKtvX0
bOWTV/lcGYf5jTK/HWCr1oxhBqHIHyix+zvgYnrNy/62KPsK7GsOjfs9pCOLgW4W
tdSvX3nKsK1b8VNiAMFf9Nav5Ac4Xy4c8QmQ+GnfzWJr5Zco++GFf7d7E5VZ3FXK
2eTSwmLthNNfaLN7y7+Wc6MOpoDt40xqrjr8IqhIH9UMD46VIXB+jZxlz5MkI9En
TTFbZWeQXs4hF4uDRdH0vM3klY+v0p2Efj0rRSFaRScPd9u8Z8xjeBli2pLaOnVM
XWLHHCXWpyqrOwDBcX0Piw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8256 )
`pragma protect data_block
KsJFjk4eWLPO7suryQhgEGRrFbGnIrKNagzGzwfYvZZDdsY3K+zqb3U1sOWozKmc
cCZKUbS3HuoFiK9Qa6RBoLDVWC956/TXIm5oQBy5wiOmmBHVNSTPqfyryEnytzTD
mJORFFygHcOB51njKsyRPrv9JJvnNI158Ov0OQj2APEeAwAAecBZizg9tGEH4waU
oOfv2ZdO1a8jITODvnakSZSThwpLPuimBCMHqCPbFuEScew+16ap6ljM0E9bapNw
OX7pyBZJCGwyaqqj5OfqAIRzQOMCCmCdCqcJKIURbcM4PTpCi3Kuo8FxfmAKxDO3
3jP7qza2ru1Rji+4q4zMySCe/PgfSukxmG1DE/gWd12zSYeiqaolBClc1V52DRhc
pZdSNBZV2DIUAHhq3tyGLvE/sdoWfRkA5pR4YzKiaBxyqDrcaEA1UiTLwQeOc7tn
tXoYIvhWbGx+e7mEiZDp5tRQmJ9bv0rxCpBBcLVz5jbbCdb/EVqBBAI/sCcwDsx4
AOhMMBa52KSGsk6nS4mSBV4UBsBNF3afcW+aIniIvEBFbODiDS8dgju+7duTC0Fa
pBf+6R35KwQEfbWcctVPx3OpQsgt3zmAuewg/4/OolQQzaZ8ANTDQ2ylCIE1rtuI
oHFRIswXaACRJijfUdqQWuPK3ZT0hDWZg60PL53XWSNb6DFMR6pwXU2LAXvTO1Wj
VnMGgM1LnA09MyzxBfNBMpGSownur1LrcHjdWj4snJBn8eogrwP1HuhEXDSWAvy2
NC/GFJ3mV3rEWES+WsY4f+vFt/CodaxmBi3rGPCJ0CcVi8SFBf+l6ajFriMrFLud
D3GVT5q16r0zZjCRG+mKyHipY2ZQIT9A2+i5YqgJYdQBZC7wK/rZ/MUduhn0OLE8
iDvYeWWbUbwf37iftGRsmKQNl2lioc9XSIsC7kItTpYfziLRkpCng0ZAj6n5Azjs
oKp1D3c5FhMpQyyRXcF3Y3q6xr5XiOO6DaCKwaU/PzZc29v45vXNxvaYnf56o2ya
Jks5Ak/cUthWRULoPLgkltko/7F3xhWlk0yLyIF1rSi8kmvz+nWTtVNv2K7YlkSE
3PbgAON4pJy7TqzHH1PAToqhdn4p1MbqnqLZVX34zWxwiZ/K5gFNrJFpynD8882U
vK/NccabHf5Z+VY9K+wz2Ab+weuXI/vs4lfNTmy96SDnCY4Q1hBGw1jamBy0Qdcz
hfhHge9svX3vpocGuvkE6qSCC8Z5ssvI0SDaJ1dHR3F1BRAvUkI/QRBVInyy24VU
bx/XsmaaKFV9fTMAU3KCkuT69TmOltMtoUnM130CNHRPaDRDWH5Y2/EmmPqgrUsC
pXdx5hBPJoERfp6Z5yPU3iucLmO1zY8IEDkpDdQpffW+VP8sqvx+f+5U8gHreeCm
OfaRZEyZeQ90S/coz9+cPEEVwuve/4T1pkRi1XJSBnDhsOmIwUnaM1baOILblwi4
rD0o12jl+Xg3IvIUxQblCAEWi58peOnZkBqzMuBhtVr5ee8wItmAtieoZOxy4icp
Xy42VVjZCpJSfavy56FFBMGxyjeYpSwVdYP6gOGU56JWssbaKLYbHv/xaLCQrYXD
drIUqFF+FuJsvPhSn7xE+hk3s8rHN23EVt4dOjPJ0Hk8GOEnZik7BFwOEXc8exh2
9oz/vf75o592odHTr2rsO3vnPUQOLBBPjjNsG2TnJmusg/Z+U1p4avbkBHfQDOou
X220c8NbUoVddkcayJvRBRc/JVb5hysPQaSDvNX7LmnvISb03DeXqN2TG4lzCd71
TUpbaIISQZJw+7ukc6kXvUOxR7nC4clbhdhl5M5k0dtTMrA6lLLfzd7+DQylm4fw
QMzLunR1THomz1hByRR13CwKxpdFx9VyLR7UCEjFPrL1xPEzHzAmDTNIWqXE9mfV
jRlKGTTf9aLGwCqzBgMjgKBQP2ySCr1OEqjAHziz140wDslOLEztDAAR1Y60XArU
d9dDPPnKEuEX16d83ZC/S9m8LHumacI03jrI191ovTGqDu1rwqrrUF/QCVwIpuH/
ivblm++c34GCCK95b9nxziaI5O9g90hv0NHtNR8gVTxQsmI7ljil01/l6/U8gFnL
RbIpvdN4RzYcu2usXMvv15FZ9YCmV/YC2QqzC86LZE1XNar+xl8ern0UV3GX157z
47t56MRS/Uibp3J4qR53FLnDrESOREAHnY1YpxqaqI758figI2UyiVyTMyjXOY//
b5uaxtilLNVBnt53pXgGtWHfChXWooQCrYmhFbDw8bE1Wq6DF1rfmfG22PTRxEyf
IzIpGpAWaxZpOMi3MbtLsn2zorspI5K3eGS2hCL/GSIDc+PU0hm6oSkn+yW+c2F3
Em3rn5iE+wRzvH3ZbSfgdmSkCpCrP0aya2IEE3fIThGZ5CJdqAb7mN7TfE+HObl4
+1CJsKl2Qrl2u0jyJYCYdUSqeZ4jPcLoLU7jd5yUiJ9cO34nW5D9q6HhZHUs2iRN
qtRUC/9bQ+T7D/qZTNs2y4lnfct+aaKGA7SPtQhRXnisGDXa4rSEvsM3h5G6JMLM
Si3SblIKRf4hwnomi/E27OGnblVaF3sIOhi6txKUtXKp4tSHBaY0amSYQX2Hx4Hk
7/p2+MKU84zr6cOoOXcCT1Qoirs5UUrbWOZMVmHf6mgX0cNW3SPgnSpZlaIj+Po/
zq1EDGC4T/kL+9F+2e/x6Eo8+VUmdY5UexUksHzY9DgJLMieGFOWvUpO0owa+WrW
w8OkEWX7DhLmVUMfxN/4Ak+DEG69yuNA/5v3odOTaCg1C7Td31FewIxKMKRgcQdN
vmCtn0eqoydKkoRU+OQv9dQrHFNx/9wk6xOTi8H6iDjntV1SwF39QPfKSu3ardIE
23Aj89gtELUoLmqFQqvfRrZVimo/d+/6w43Kuw2bDB2JLVw8W8EQt6lNe/gkW0Ox
WwG1J08x/bgAi57bc9QJTihAXEeANnWkskV91SIdWJsfRmeJHVBhmFqkjov5gHm3
2yTvijCxHR4LY6nLCu7IaZ1SqMC0mHY6i+MbASa60lvzVJNmX521vR5wqiUw5dvd
4TmbAVi/zCRh8w9Imaf2OgIB3P7y6dtvzU5/mgVSCMS7eWo09VeggywNYgfBNr0i
kjACpG3kDWGMsceXXK4DTAT9mwua2lcBh/z0qzP19BgBuyGqlzeQ7y9m8BbNRs/M
W3PWmrvs+Td7o0x67N9OqUtYaWvJnag4QiKJIOHT+13+mNifR7OZ7GwkqBKGlimb
8U9TiLxDPQPqKm3FoCEHexs/ELWRIKDp/09e7tt6Ndmdxpabyy+s8wAV+IlggYT9
ZD11PZDcp8g54O+nZo+kGn5MNhot0flu1NIKmyeqvYMZiXFqhVs5yXkXLdv6lIMs
f6AfMMZWDIxLATXbkd/SN59LqG3wMGBgvFAsy4gS+R9YTIBVfcXFkRCwh90PYs13
xtCkH6m3r87j8opbnlLot/5K/2v6pvgVvm2iKPfled+yeEpmNfowpIjigRdA57l7
evn4BD+hm+1AW2GT9RIaSqX72xP0R4bd3HUnN5dG/OCIBJWlc5x1bVnnU5tUPpxb
FMmrYEIYldmPO0DLpQxuOiAjBYtp5F7xRkNLHb3JuYG/5xj5wMPdel9DF8dgthTG
u3KYJvHWyIolbtToE05r6E/M9mbfinut9AJYPoR/lsu8ZG3pYMnw0FR1lLOvss4s
3G5Yb+zu69kWURbR1rEfMhlZJDs+X+i1/UEP/WfJI4Rq4CBt7hj+cwos5lKpqR1Z
moKRoapkgDYkkiITe/tH7zfxE7Pj6fWNmVwOXFXIeeKLJ5StGYMM8gefYW7ms2II
5Nuaxz162ooC8txiFMVRcwt6Kr9Z1kscNQa/BCS8pvqz7syBbfs4stxIYbpJ15hx
UcYnUL3rOn5yAUmh0bnAxHgzWfbxe/yJsbVZsNYYSZcC6OhbzNQ3kgNdUaf3ppug
nQuDK5Mdh8eYvx1Zt71oXFe1gJNlbYTNFUs/NTD092yi7QeKdFP5G39sv1vvw6U6
wwqw18AU3aRuPVZIKjDeXYEjHdr1RZSh/VRhm2KVXn5Ynvom5Lma7o4ViXk9Bd/n
PS+t12ZT16Urj8mZvLmMV+sO0OftNHIebShUvMJQKW4ruOSG6AlTBW7SQ5+EAYyn
ZUfCUzNZg9i8/OPv2BZKBqLAVy3MYJKMt2Jc2B39XyZwEYF2TQlVQr85htcVTOxV
G6YkPr3l+m/LorFOgaR3rtl+KCfp+c1+qEJ9eAOjSj/xd3XADfugxK5p/2r+mNSF
gbyAXbPnX8f8klMnM5rFp8M71e91vp9EsF0gRztyFv6hrbprppIuxjROjAbx1D0G
48j81Vg7yKySjsTxd5SqtZY1JS29Nv2Q4GJeMHK0RKsFvL4AXvyzaNbGYfc5EtTP
V38hym3/UfSZEWg603dOUXfJOjYNVGGJRluntAovQMpnvc0c0L0qk97DygIFD1An
xhVS5de4mee3NQxEc+Wz+lhP95AeciPDOFEqG87Xxd89qO2yi3NfvGly20S9jfEh
feZ4QJ9EtUlDDjV2bgvRV8spYPSy7msLnOi7D6ZpYtWnIXA26wXieZe/ftiABWyM
kYjFVpkXDISBW/DKCnWfJe7JyJtqf0VzpY2JRvWHG8Hze0dHKUZFsL6cHWPsOQZq
voc8SdJ3NG2qmklLeQCdKqo4TW9rjfaiSlM27YZQXxrEJhA9ZvgsBgzrs33G9dbD
EG8TEGnHRmDlY9scWJ8GFIoYJemkhslzMn6m4tkC/Be/jNJwo/8FpMnW0N5IRx/H
jz7Z23QA+qTzRsp1jJ+SShgajp++KxFOCg2ZdRCzSyKukD2H176+27Rq/SsXvqY8
cGStUhn1MKHUKDouNVz0uPLUB84r7syEJhE/GDCRXQvuqOtba8/znZ4iKdeSC6QX
VaheYfiN8Q8k45qtHO2oy4ZGJJeZHCNyVR6JbwIEEHMsQdwsADK6v+Xd9Si/1EqS
Sk0+p6Rm/AKy4yefOr1HrraUtUqBcn2StUzdWbp7lcKnZTwJaEx4qYNVWpfgtYVP
T5gVv/M9H8DYkdNjfJBeLAidOTiS8sxYy+yDUJKYI+TQaNU3c1uJFYeDHLRDzYtw
TpT1+UkKhgPS8hZceYXZueprm1AFbZV7vcwiPsJrtkCWm8rylzcUPmdsdc1KvzgT
J3OkNi4XuW76E89cbizTu6jfcuFTaDlasK4D0jKXl3wibOY3BYaNEYfcQ1lHJ0hq
rFgD20uRHRrPDVAUHkOwgN9xw+ed4W3wZRVNeTvvQa4rAAjpbAXvM1QyfvVkkTSl
4TKKdZd3n0Vy9UKfhANZni6ULsu/5+V+ubzdqn1Ui/RFJ9mOhyzyBYVq73cgRYZk
x1qiQJu89SQdb3pwDeGN9pfsmM5ER9lvkE7qiQDQ+9yVQcJP7dxBfSg0Ck2Tjaym
7NPjd3W7YLAi9KWFSS42KqiuWNUXb3+A0kGNg7NKLtBVy9zr7noILfLguF2jGoVd
2CdNHeBb8fFPwYG3HTNGIwSraf7cjuxXuY4Oc5zpiajR1dOBjTVca86+H6L/BIJs
wm6YsfXAT6pvqNWazobsfxP//Pm/n4/ghuTLH1CJB0oSL8oPTUVaiom1UiCPiE6X
pSs2jFEiXcu8S0Zey9aop+G0ikkcHwYRZxjX9XnHfDVvo2Q/BSYUSKUonOQVF58r
MaVaKPvirsvcfQQzuNITB92xOZkRgtEEHPPdOQCwrmgopwlN0VGQy0LCrncLFOYh
kYI/D+YwoOFGSbqIbcj4+eHPY9ztIDHj8EoQWvuP2z2fZZuO8+oi4mDpCazJTDqM
b7BaGQF5thy81RY9ygSWYN1RA3O1Z38SZ1Qj/WqwoFoNrloEJmnTKcTDQKJVtODX
43dBSWn/pOH8HpCSF2Ul6dpt49efoLbmIwO0zOJm0mnLL+pM6wFDVEm6+ALGJ5t3
9tMDDGnKZzCOWinOqD7+4pzWTQtKatRgem21noTyJRCl/EGAGtz1kM2dJUGp2aPb
3icVqh1sPzq/zhl0n7XirGJMs18O3bIWLdseOuVL5jGVciD1WDZUwt1DQmWPYkDf
x3ioHyrcwyEt9iJdHX62lJp0Nk6/wIql6FK7IQRUUFfb15ekmItshOe9FDAbyhog
P6r6a7sAO8gONp9n+OzMYs6tEyETMi9rUvwJwE2mEqvzqqQqhZlpFTVj4JjaY71G
+0jjj3mgHBW+xe+3S67sxreKtDGBdGxCXagzDcj7TRKyD7fRmguQvSyzmKZsBCzq
cQ92s1VHKsUkbz9PM14o9gozdLx3VKZ8/pTk2AtI9x31baXKFtj0diINzau2s4G1
AUzsip9Eq/HbH/sMw5mvWQeVr59CfAqlJV8eDMWg9Nju8doSq86+ZYG1NKzdy15x
Jyy+fr9nZgAg1xzpxazQz6YxJiChg57IMw+zxruOnGC+z27mnY2nec3JCDFng+hr
CaU2ReGbi8sE6K+oN4pOmWneRE+XXlrXfDBPaLh0TUd/hsTxH24oKE+1WecAFvwf
gwl+i0j7ovvhwTBzXPJhHj2+aY1VYtw/blF0ovQZRRPBNa9Ocmw8zfcqhyxlRH7j
E0MBmpJszy0tMuA6TOYpU06cnL22CwBX9n4yqW4+BgVDnVqwhl+1lvtEE28/pDq6
SefrBmc5jHrrGmbw2WZmnonHe65V6xZY84hx8c7QuBToH7/j8MpI30+nz5fg0gv5
OIg1uaecEwmQf0rOg7RNcffAiILKhXsuwZJTUCv574KrLOHcndCFbMYL67p4/r5l
d96Pi7j2Kz7cbHGzcc90Z84DlHYo16jJAYnwH7Ob+QTdhRbXmpnMDOKBZzQgv9oV
hS9HxaKfvge8Bf+eR8wdjw3kIkGpaFecIbbXP1ON7K9cpOOIQslF7mpNxb7O9QBS
vyRZuxEbXZYc3HBnamTqgv3MH+zVfo9olVgjQMtMTu/Ux72bFjULRqgbkhvoy0Vc
1hb9LT8Th16JITtUeqfItmKTk/f0qg+8NJUR9GUoGnecivDJqE5c9cdi8NIlvmxZ
inO1RIQknLLx6+qecNuY/U3ewH7YpqlG8Grl4kGe4fpjiu1z4bB7+28Bv5SisemO
ZnZEtP+lA+e+jtwM6jmbISEnVGBqWhs/LSL4UeysnTPg1ufD2W26rhXn8Qhk0nL8
v3wwcxn2jyP/de98IzBXve4SFJW4D0exrYnGATlOQbCsTPCp0TGYdznP1JtLSwMA
dElo5wa9fu5wJz6hE3qVk+I+UvU3ijfsFdak1lJf9e8r3fcdyTB8D3w4eqjEsPaO
539L5zwWsVqIzuCbOb72i7ei/O7PDYThUJ+dADGKFSULb/izUkm/G54tpOhRQHHZ
5gNE0FJiYwxlp5u0vaGrNci53nPOE46e1fNnhiGmFP+fFqtx2T3Th03oFsPqD4Ti
KnnAfFY4wg9v5mlEq+ZsIXrkhDTN0+KNUProF9acZmSp0gudI+k1jHQCj3NTlZHT
sydveTO1VFIFwg/HtJPfVFXNNReW0DdQAYuNazdXFKh9VZQsfN5ypOyEbF4ohEOR
ZQIo3x2f6JRhKd+zJGv5kNQwx4YMuUHkdRRuuplQAUweQ0bmoBAVR5BP69qU2hev
zNEFTAj+cLJuo/h433zzbu/BH0uaimjZqMPTIplCG0t6B2dGcb0Ash0AoO39YPkE
vVR4d/2T90nVz3zldDKpDChJ0t/ZjcZZLQ7jvsq5nXSxTjuw+otzrcIytXl7qxMv
tLNITPohe28lfFuzD83lGPkmKg1VywQlzEYwI/pAgEUUvhGSwKs4gEmGQ900FSGO
aV8TqfkPvC9t7HtZBmrSjVS6vFGK2sUadyvlBK14YPom74YSLoXCMDssKKUetXxJ
r0jiTpWVZsD3vAMPce9qoaRpFlnGlLyW5eO8TiCIDIjrmHJ4/Yw3YDssHtVyPec1
GuW33W+IvsbRkvvXX/0YpNDCHKZVE3bD1llpbeJlMOBfPOpLsIRje9dSz27I4Odr
rrL1XtwcFzTLO2bZF/ya5kvfNXuZ+G8/b7y7PXg8iKZf21D27KLQAzUoCIppQSHp
CbNSmwWuZrh1enavPIMOMW1iT1+RKps69YAXiBYBjHfoBNRXNb8pwPU+ULdGj1Zb
GQNFykRhF8CXMqbf52kofRGM9brLZNKhsCZ015rQSt1Bsi4+SRegRC3XPV+TRxbF
ULsP98l+4W+cLg5VhPzVtBUF6BTlzdC8VRGLnQiF5bVg/G3+hnm+ZS2WKEGEUsPI
18yDPES3pZufkSWov9KTtI1t/NFr40YriGsn7vEe0O46vxVHBINsr3V6Kf4YuKZi
MdGsA/5s2O7ZdGQ7IyAKcdrHPIkKXZTTIwQTzNscy1q8GRFrpQ7CpQcCKaT12jDO
694vHsbqlS2F2e/mc6Q8skUU6EwDubYCTM+XlAZL0owI1kq4XqlKB27rJogAxGjj
vKJyIjHLi16n49lkVSnfBbqNugSfHoWgDF1x2IKcSPUZsBb/ZqC2BdA5WU1nlz+h
RApgumREDoku90grt/YZZTeYLO2SXf/ZGVtXD8ClkzsG/+bLpDnFirgOxkVAeoXA
HICtzgUTN4N1gCMLzawrvakjrC9zziiOYScJ/ltlWvN906+KnW15vYV95kaIPt3l
Qc2sueii4zOKBZ2f64JMckPBxCsklfsrWGN0dYwTvtDUdEXrIMMFHFEilc0/tl6P
c5JPKBrXQvyZGDHZItyxxBC0GGMOMX4WSVaeuzfA2HxPvdVn7tadCX4KKhKliCLE
CBYLHTFheOL/A41E/aB1oLmUY5tymVonRiKFPc9ZyLGzmwn7+8hkJkPAHxogSTrI
WtOSXF7X6G8NjJUPwd2TJ/SGPa86D2EtgRwEf+BXgBwq+t2hlw8phIvM7gZha5ar
GmG0U20b+uuh54RTK16jZ7K3BQAaDyUZFn4QTPfV26TrKSApNZQkoCu76Z7el2WP
S26bjR2XXJlPFMo1d28O38GJPmkxMOfHrbyoqY03C6CcAuBR06joRY37IBpZcyrX
xZCh1wxd1y1rK6XYrnvPTbYzhg9I4rOXav/mvKI7pTVd8B/FQk3/Tby6BggsNHNQ
CblMobL+UiBEWYqVBf41Gg4LunRRTOmrYBxYmiwBn4vlwdtBCI8r/U/CMOh9sZuG
MJx70jK42afV/Dg3YbabBHaMZaWsM58n2TBE1KzMklC5gy8iFCyMnDdJtgK9vBN+
MXHEolzfS044dcr8xEKLk0L/KEl/47IDVwzGvAeqGoew2ozg53X3jiR6wvPMvBEl
s6eK4C5vK8PqxJfvqI28LIdyzav0p9X0XdvQir9HolOig6Vpl4IlM5+beFNwX7Pq
wI9HHgEh7QhhnMnw8wzL21gRlHu04bvVBmYqQs6pcp8MHi+mvCzCBmmLsVKDbGzg
ldV5mMdN5DFLHBKrjblZkpjAruLmFfQKMm0qlOmoAbc/aQaZOnCDS1ruAvwh785w
RylgVLeiSjNCSGsqkdSc/rnZQlJGPXfXUhwI0o6D4T+W08wDBJHPw9rF7CI3/Hpw
OkXb5jkhmRu9IEJDXYzEm0KdvtOY2nEpr516KK7fn3S94uj+/ZhwEE5F6vf+8HJB
paAwj6pWZOLg8sBkV3Tf9Y4Q9fvLGZIxUiALNTwA1ASlVIir/7SWwmppi++KOIZj
9MXd24moJfRpTCGYhXi0/rsHxCQ0+mhsfJpJAkkHcRxCWhN4jVTxoG6FWTHcawzM
YPMLOzgNL2pENaHjyMA9HG7kTtwj5A6ZIbYC6GXAJ108vimGVjSdEge4DYxJpW2+
rOq21z9xtaiqkE3CfSQleHZjOTqyF5nhC2oFkvkkxLAMemzH9OeG61UTqEy0vkld
KvrnFyWzmX5EnzFzG3hZwNfqPAr5SrI8PQbxSz34FgzLZTGyHZAO64hy0j4PLvUs
WHC3Bj592sMZWCBs1/YutmSSstBbmjV0z031CYy/2uvN3CloS87phhaDG+W9z0M4
AhvlNYG7TWd/3yIWrFTtFnRtoT0gTPIBsBlcaUhQWDqZ/dKyEfmHQELaApeD/NBj
+okRfkhAH6W0TBuK1ElDnY5H8m54kT8lHdNC5BGxKNoBgRDJPRi1XvMcFSaUpCwx
a3RO7z1ecQ61j0vslkfnrYmNSuJfXhraBmzqoTlnCKKSKufFpboxOayQXBLJK+C9
7DH33D1+ue0dWc1spKTAsUV8ObvQ8TQ01ottWSjgWeLgz+DPFK0lRfw29/aGvhAr
j/w8iQ+23xiCZxfKf4chSnaZg7Z5G2Nu5nqxRgIWh+gVBc3OFuKOkLAmBPrOB1e6
eMhoI4pcS4PaocSTjuLjJsGqYAS9dYJToZlNUW4W/pjPyfRk0ej9OnlTCW93oPSs
y5/Qb3iS92mWyiteIzROk/oNNUs0l54Iu4BJPi2eu76HX7H7l78315w5IYtrnVR+
007kfJ8igqoTATbFOAb+3rZPAGkljCZvMMbNOW3aqjmDTfwxgQaIKvfazUmET19C
eCdDLy6RkyVWG4ARDqNuWAt6sXW9rhXaDSD/PrGBHNN6gX67ZbYvKnwZoznoClWk
ykp0+0Kr8yBfrcYbqhBlmUJ1LbgZM7XdHvFSRbGdZKGV7kK5h1gJpp2C3Va8P+Iy
BeXePiTWRES78jRt5DOPdiqUKxNUlxGUj6JiahsS1oUlII/6LSycszl2M/0A6Vdn
Jz55iEmHF+jiecezcswY0oricfBDvhUbdP+SiRRomIZByeNkggrd9LhCsOsBPESl
KTo0lNqlPaGStWx05DmdKOYxs7gQNgWE07BzhhFKwCc2Ydgj/vqjAoCnrYIDJpBO
77NgMYZFjwhj7uXyEoA/DZtqvsM8quf3fpfdE2RHoubN/8jyHJxDxza8B6NGrU5A
BMe6EsXKa4YulBPVbTzK9L2X4CaSqF7liAojQ0Z5MBqJPNui6wSoFFQYnjBB567X
YFCFfs4sGKn1UWM1jtd6gDp/XPTbYnCiMRLiPh18WjUxgAiFAbaSeJHBVaEoP7K4
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WSMV58Nliihjh11Xi/oE+3EcLVmKYrAf2dgqt9fbaQGHF87QEj1+X4vPnqlIxQUk
qGsq6OXUxG8apO37vc0dhkB50eXikoainWDCkI1fKshyOVRpWPIp2Hmzztc3u7FS
E6YFEgxbCfuJ4i8naFZOiCjOLJDHekcYAZi4Kh8+lSubJLOkXfGI2llulOCjK8vA
iMgrRbEX4vF8czShQKOwMcvf0MT/SaHjUTXxhIUAcMF3SyAkoBtOjdh0ecpUtSE8
y2ccb9kstxcEfkoe6c6HIFzx5m4tgyugGeQFApMc4tN8M+PtKOH3FiNeCHofgoLs
f36mnV3cQT3O2Y4hKWcwDg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2672 )
`pragma protect data_block
eVe2XwWu4WMuFAoN/2xpnt8Ipox18qadoGqukzmvLAbzZF5XA8qzm+mn+Ssml1wk
a9lhhBSia/7p2VvCqPnsKJYydPbNxETFvGpDW52CNnoaICUuimCRCD8ebB67XM1F
ONCD43w3JsBbiA+P3P3Mu43rpf2z0R3d+ItxNCjGB7TUrF8eKEXQppbgEd1QDXyQ
Kv3x51LzEa5qhyUCdY/bL6LITk2MMaUsclzQdb8U6VJwkpYzbnI6HiVEmh7suvTV
s1UgPPNQ735DTkzyl+yPE40jv3N1g2+oVjc1t9fLpBKwtDADLE2HPmQ/Eux2/oPz
INPgdfL23xSixZRIHbWW3UtvOikynfIYXW9nyr+MQAi+Vb76NbtEAflNcoBNRFoI
IBxRn9bZmTBOhPym8RkI+ykAo35c+Pd5QqJ57jNb09ugYA0nM8I7L5QOuOLU2YcN
mIOZ7CgJQlNIeX59x8IjSf1BERYzXtkCqx4oRi9m6+d0Eukp+ixaB/U4cE915FWm
dm//u3YKB5ajMs2atR+pPlND2+VfrdjpG0bFAXFCEA4c20THW0I5jlGxca/pV1Hy
pgh8l+azFGZmH1bma5uozcbgP0EIpd7/fbFynbHJ9geANGqAO15TT8DKV6ndEF+H
KcocCpPXn2PdStmouNedInu2p3t7gDJNVJZKhGEtUYOA2KQNQwno6U3hqyC1iRnB
Ron6I9JJRYDoq4hJkdY4fTYEPCVLSroI66bT+wjfkkh+SgPMlN/8Pgrwl0Izwela
BO3C8GgrWFWOagrNCShq1qgTur0FG9mkkn1o4ZfCEw236dbly3PQyaTTbTO6kayD
dv6hgkiPZA3tTQ3pwByCESzGU9WJk9rhOe2R0z2h4AzzRBVBQyevpommjhcrxDzV
NDZ7mpK7DYE6f8svcmLslzHuvsKPPQ4TDGcQlgvdFjOJqUpfol6IFu+7muDolIon
zClO1HVLV2vMUQsSvRyXJZ+NUBagm/rG+Qzlu738B8lcERefUtH29DeLP17KwzcZ
VJ0BaTpbTdUk4SvhnLn51aLiAzuAkbK3Dt+jcaKYT+LaEtg/WMtvKP3sqDsp/Rd4
2KQY2fR478Uw6Iz0sLH1mwxO5aJPqn3wNnoQCjppw0C6naVQKZrIPUX+ia4YfV+o
UY8taZVZkjQAu55m31bzfqbYIR/mvvLcaatLHoEViP/eiTfUe+NpVEbn2YhlAEWS
5im1hfWYfK14CpnYt9rP21VNODyXDdi8Ic4DfkLk8tNr+QVbIf1gBA5FiMqj3Rmp
5/2VBNXPPBMooCKu5PTGrqxhTgKdt+lAHr9Bqqms/B+06Huhoo+FsP4BgbJvOZUX
7h/mURDsBCpJpU+PuDS1qpNMDafC9G6fRisP1hgNEjCVpi71zxMno0HOZcz9qSXK
QKHit9AdZEP0EIQzmc/WCI1q2YoNSfsnUqdx50mjimxL44CPu+UGuI8Z8BdN757z
SKWe43JNda/ucESAkRxrATuavyKifgEUOy4x6revve2qWoFLFUo5gUJY155Pr0CQ
BXF6Nx2v/YlwROgo56oo+1L7jzV5sAicIkEYqDIPACCjX6PJnoZU5rWv4XfeBtwr
KqvlaPZNiMzkawdDswD9PiOZrGB9hoL6+f+t6Ycg2FE5CIepoGnLw+WX+HzpuQPf
5IsgH0iWvLN0GfG2RndMYvPSQ3nGrlSQMpoL2Uc0FRlmh1KwgpRz/l9Ly82hmpDh
YzKo0ceUnGXRnlKsxZHGcomk6MGQZ3qTg2gUJI0h3P3HJT02e/qkuXGEvFRKjIXb
xrqVGTIsMTkOhzAPOyawdXGt5J/D6X26HcTs7riPictloNNTwoEJv5qjQTHg7L6n
pFdOr2vKHAxldrbBct4HexG/oA9e4l+U0Qy7VhK8eZ0ARS32k+UdFP3uomvTnPIS
9s9r/tMNG2XnVO6bPVWYRPZ4T98w73Zm1L28vfcxzNjUaycJeexfQeA43pyUWhBm
ecFX7MWFFfkiBAb31z/OYGwMpih7xEjz1acYsLW3Ay0A0EQ9fBPE0JpVz2v5DrQ7
7uaQlYBroSRPgRuAG9mt8m9hRBefQKQCBC+hYPM1ankMGfxiqvp6QrjVmfnlZR8E
ZO9z2BI7xd/QE88LKAOg0iWZjQWjIaC5bIaNsfovs7ajPqi6z3tZ8hXSEhhz2xMR
5GIUZgcTzwTubKmlQDMBWAXnFzJjX/pCy+gzPMZQ4925cU7BjzJsmTEzSHd1kE5Q
KAJK6nyPAIKwMucexT0Dv1DwONtwRKpdu5UVHvHdMtcraOmnlwydLDIXes1UOSaV
uJEwLGxBkPl3ttlVGM2jbIKvjAIrTSVuaECPfnxraJGHBtjq6goUgSgwaAZL338j
HQMcYi21Ks+UYeFgQkllilqxIKNjyCJiaYGcTbNsoTH3Le1CJGwYmopZcgTyad1b
bGu6gWjgfBws+DJQ9oR08bGDrC4NRQhmS94fCxBhL867RZj3bf8RXV5xhRyXHXCJ
jV6109EdsSo7jEEXE0BUjAnkLWoj3Wtwu33TQP6BgxMT2gGsKsq1JTXHQ64I0IJU
hqjsR96wCoUfnICl4o6EZxji5OSS3mO3wfAguod5EazVL0ryg9wbeXSmFcrtDqlB
t3WeARC3EjH0WOa+MsFNOMkixNCxcvelaIPcVQ1HJRtHhE2TwEpQWYW6o1CD8Ry+
AUkbRlEmXmU1nELeKW6E9MjV742ST7QMdDQZe17wZVEd/Tx5EWOVCi9i+mP+VvgO
8HGNQXuNO8NVr7ihA6YyMdOH1qiiXnte/wyec7AN86ecl7eAqf6C5dPHLdQfP48P
stgrk+8BVyiT3m2jgOv4lkAAoFY40Iwx2S/PDBJO/7eM+OIheiPgmMyDZQkkWcT4
Q8T0J94ZwqGiqvQ6xGbqiVXuIGtJAKGuQ2d0aGrkPDDyY0omMglxQO4yD5eenl6E
aNfNcnxi4/XlYDSToqFmNA4wWvQvUyXqPXxVIPzHDtHfXYC3Coy+oHbNmd0POHMW
uyBVnzFYs1GIWF/3NG9KG5W9w+0zXT/lALPTd0s7QQFVR2NsaUSiwM3NxqZ7ss5+
iLVfgXpB5AlpGwiiDMnQGW48nyInnLxDUFZ4ODcfww65bYl9McnIvbKgQFCwraV/
3OFwxWrEO7oqTlWOsvXEbCZUXDQREtO1u2TH1LD/baqdMW/uo/ImEO04bmr4CiGq
VSyetrJZPOlY0SDaaBdJPqbr7vHHBcz8+YMxnEd6YnpG6OSntXs5mQF+3NaBzVdt
+0+8AaDHTKabmZ7ob1aFNvwdlSmj4ikWLtblZ6kNUC3HFKaVdmDi8r2/AEjs/dup
++2vsMIViZAhHl3Cz6ZhUZzqWSUW7zdYwxjAUKk+0J77au5EbOfMbRtUTfiQSXfb
pcEkPmPIhvfHjFn3XMMnTg/xbcc3mb6fvdAH3bq0+fIbptPY0DNUgAumGckrVE3q
Vk0qiS40P/66TrW42V7Ggo3thSQHWvrCnj6tinxQKjJaXxBniMWW44lYDtSOAQQL
G/yk2YwyXK5djVxwKa7JRsb5nvXUHCeKvCNBqNG4jLw=
`pragma protect end_protected

//pragma protect end
