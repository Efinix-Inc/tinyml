//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2023 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = tinyml_accelerator
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Wed May 31 12:01:46 2023
// ***************************************************************************************

`define IP_UUID _990a5962222d08a75c39d9417cf39c577ba9ee26
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)

`include "defines.v"

module tinyml_accelerator #(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 5,
    parameter                       ADD_MODE                        = `ADD_MODE,          //Only supported "STANDARD" / "LITE".
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,      //Only supported "STANDARD" / "LITE".
    parameter                       MUL_MODE                        = `MUL_MODE,         //Only supported "STANDARD" / "LITE".
    parameter                       FC_MODE                         = `FC_MODE,           //Only supported "STANDARD" / "LITE".
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    //Convolution & Depthwise Convolution OP Parameter          
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,    //Only supported "STANDARD" / "LITE".    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,        
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,        
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,        
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    //FC OP Parameter         
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,  
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE      
)
(
//Globle Signals
input                           clk,
input                           rstn,
//Custom Instruction
//--Command Interface
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
//--Response Interface
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
//DMA Master AXI4 Bus Interface
input                           m_axi_clk,
input                           m_axi_rstn,
//DMA Master AXI4 Write Bus Interface
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
//DMA Master AXI4 Read Bus Interface
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);

`IP_MODULE_NAME(tinyml_accelerator_int) #(
    .AXI_DW                          (AXI_DW),
    .OP_CNT                          (OP_CNT),
    .ADD_MODE                        (ADD_MODE),
    .MIN_MAX_MODE                    (MIN_MAX_MODE),
    .MUL_MODE                        (MUL_MODE),
    .FC_MODE                         (FC_MODE),
    .TINYML_CACHE                    (TINYML_CACHE),
    .CACHE_DEPTH                     (CACHE_DEPTH),
    .CONV_DEPTHW_MODE                (CONV_DEPTHW_MODE),
    .CONV_DEPTHW_LITE_PARALLEL       (CONV_DEPTHW_LITE_PARALLEL),
    .CONV_DEPTHW_LITE_AW             (CONV_DEPTHW_LITE_AW),
    .CONV_DEPTHW_STD_IN_PARALLEL     (CONV_DEPTHW_STD_IN_PARALLEL),
    .CONV_DEPTHW_STD_OUT_PARALLEL    (CONV_DEPTHW_STD_OUT_PARALLEL),
    .CONV_DEPTHW_STD_OUT_CH_FIFO_A   (CONV_DEPTHW_STD_OUT_CH_FIFO_A),
    .CONV_DEPTHW_STD_FILTER_FIFO_A   (CONV_DEPTHW_STD_FILTER_FIFO_A),
    .CONV_DEPTHW_STD_CNT_DTH         (CONV_DEPTHW_STD_CNT_DTH),
    .FC_MAX_IN_NODE                  (FC_MAX_IN_NODE),
    .FC_MAX_OUT_NODE                 (FC_MAX_OUT_NODE)
) u_tinyml_accelerator_int (
    .clk(clk),
    .rstn(rstn),
    .cmd_valid(cmd_valid),
    .cmd_function_id(cmd_function_id),
    .cmd_inputs_0(cmd_inputs_0),
    .cmd_inputs_1(cmd_inputs_1),
    .cmd_ready(cmd_ready),
    .cmd_int(cmd_int),
    .rsp_valid(rsp_valid),
    .rsp_outputs_0(rsp_outputs_0),
    .rsp_ready(rsp_ready),
    .m_axi_clk(m_axi_clk),
    .m_axi_rstn(m_axi_rstn),
    .m_axi_awvalid(m_axi_awvalid),
    .m_axi_awaddr(m_axi_awaddr),
    .m_axi_awlen(m_axi_awlen),
    .m_axi_awsize(m_axi_awsize),
    .m_axi_awburst(m_axi_awburst),
    .m_axi_awprot(m_axi_awprot),
    .m_axi_awlock(m_axi_awlock),
    .m_axi_awcache(m_axi_awcache),
    .m_axi_awready(m_axi_awready),
    .m_axi_wdata(m_axi_wdata),
    .m_axi_wstrb(m_axi_wstrb),
    .m_axi_wlast(m_axi_wlast),
    .m_axi_wvalid(m_axi_wvalid),
    .m_axi_wready(m_axi_wready),
    .m_axi_bresp(m_axi_bresp),
    .m_axi_bvalid(m_axi_bvalid),
    .m_axi_bready(m_axi_bready),
    .m_axi_arvalid(m_axi_arvalid),
    .m_axi_araddr(m_axi_araddr),
    .m_axi_arlen(m_axi_arlen),
    .m_axi_arsize(m_axi_arsize),
    .m_axi_arburst(m_axi_arburst),
    .m_axi_arprot(m_axi_arprot),
    .m_axi_arlock(m_axi_arlock),
    .m_axi_arcache(m_axi_arcache),
    .m_axi_arready(m_axi_arready),
    .m_axi_rvalid(m_axi_rvalid),
    .m_axi_rdata(m_axi_rdata),
    .m_axi_rlast(m_axi_rlast),
    .m_axi_rresp(m_axi_rresp),
    .m_axi_rready(m_axi_rready)
);

endmodule

//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
G9sOjA4MnyQuuCyERrt+1jB+vHyHzG+Lesxl5qwlxAVUyP0fUZkioJOiGuDRPmns
bOeLuIePNA1f2v89vwmB4GG1kqMwQsgxjydPbMQ7+Q/LgNaP+eG5GB1rtHNloYQu
BGHBVMp+9WwQX7Etl4MoHGw/tW1ux0IwwLccRJemXPl3SGmGmth6yhynBvtZVGR+
+nmjjuxlxXOVaPkK9CrXt7zBWwy2wyRiW8Ji+S2QmSh8Tsro2jEgK+ykzVf/u86Q
Op1pMPencqw5PIlb9jBuI06r+/yilSHVwv2EZ98Kthkn6JyVbXf2gYuFLJY9SVWZ
vJjSvCuDMqqPcTU10nTGVw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1200 )
`pragma protect data_block
KGn7axyAB6hvV20gTI6cNA3FxSZD+fZ3f6ev//XBF8oS36Lird3K27eHV6gtjqH0
rn67PtnxA8N/ytZHHtU1OL4PFRYNE6Gc6XvKpp691OdZDzlGG8BzBe3mNuM2Mv7S
rEuOtVLsSztdx7Q27Lu7VMkl0FaSQq+PbwhVjk+eMkvBVXSFN3GXf3B64MyOp5hi
ecOf7zPiyE5xlgF6iJV1fDr75oCOYpPb2rExe1TcLRkFByYpBO3CAXFn597RovWG
G5KDZpq7fzthE5FRjIdwJqHKcbPW2aEHSNar6/ObihiDviihSlBcC+5JGDhz2e2G
vourREX5dnu0rzpWu2gW+TNyvw+mIWoc9R15PF1gMyPcr8IJ9FzDXwSw+/GkYlly
SZPraJvtRELyVFZcyfJWPoyoBzulCbvpj6pPdPl/0NW49sN8sk0nbuigQfV7Pwlh
FWV+EJ7kPMaMz+0XtdJ0gLTnhZh7YMN+dvfxgJZTXQMmTVW8L8F8gNLQj6/JMthR
2xFavnZEnXG47vMpKjoH77+ZI4rh8Dc+iJVt6EboamZXD9izU4hJ3AdWeQWDa3gH
l1NjvoGwzJp18b0d9aD32O/XqfhsXZsPjGEYqOqkfUrts1KeCDOCl7dJ5NGQIvBq
t/aZ6XhWwlGghx6A5fCbDn3kl+dALYrEK7WTmLLraJ+N/ajdRAiqgQbDChrLSq+v
oinJm7seN9fRQ6Ru5Y2Bpj8XV54qR8B3zhouknFi9vO6kw7pl6LLNBTeV5kstUrI
Yrfz4IAqSLeiHg7VKjcoLvFgrTH3vcTXqleRgprMKlCrABRdBzBqie9DRm5wLveg
XjVSAC5CgXjjO04QkEDyuq6r1Ti0xiUZEpU2w6j8hBOdgux3NZXtKVe3NVtDk6zd
DZ5JjsPwKDovEr0wSXo2iWf6hr9l7Rzc9yNDHlWlDN2cPhRQWIa3tcvTwO0cn0b+
JW4LVU5zDayyexTmj5lJq73lS51mN2VelnmkuttHH0ny5EHJqv/MQW806zcRotEk
vKgXEkgTRGZfvWn/kKmxRLkeiASYHth7d4SV0XVBtxwSnMQdGKRgyouwqH+4+ic/
AjqQtVAY68KdMnzEPCiGBrqJRzxa4vnKMaqvJXlujEDPT8ZzAfhR01z7t+jMMpGy
R4n/i79jQnIDjNS7f5hgSH5jA0o5cgGVG7nytLdXeXEqzoyDQv+05gxIMREzMZVr
cGPzSGnMYUPfioILKHI7M1eSvcP7c5JV9Rtl/xihx7+oOSEkS4NoN45RlF3swkyr
6CUqfmONJBcynROzpz9zdcGLYHmASc01cLJa6ENvjeh95ggJDEhS+vV2Ww8RTG9D
yS5apDgrWNw60ogjHNFHo4n40cTwiRpEy8RDq0aeDBCDDhaWpc67cOoc2dTKNmfY
M6kMPLPqzZgcImEaQkLYAZlQ3pAvxX73+nVO7uvuTsg52mngdEC2KbMc9de5xWCm
L5cMQSB2WhDuDL2b70drRtWvzt1JC52Ho2R+L1obIkgCiIaNxsN78KFq+Sn0K3sa
XDV83XvLMKhoqXuYhyO8TDm0hW5P3C9jo/Q3WxD3Xg3nD1CwSCst5dNSzad3Q88c
`pragma protect end_protected

//pragma protect end
`include "defines.v"
`timescale 1 ns / 1 ns
module `IP_MODULE_NAME(tinyml_accelerator_int) #(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 5,
    parameter                       ADD_MODE                        = `ADD_MODE,          
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,      
    parameter                       MUL_MODE                        = `MUL_MODE,         
    parameter                       FC_MODE                         = `FC_MODE,           
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE
)
(
input                           clk,
input                           rstn,
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
input                           m_axi_clk,
input                           m_axi_rstn,
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ib8TU1dcKTxVl+qRgTDISvBc3WuY6oe6kMviyQSRoREbkSFTdj/UI8e9csRzc3p8
vOzsB4BIoTESVXnbxCmVzesoGwICoN/6Kmd0hVdAMIk7Jwhm3Ab6mVkwA8c43+bu
j4hbXNQbBIPt00lXv705eAKQVey9wDc884imtRlBW9MP1yum17U/IgM/ewolwHo4
y5/z88iUyfJpJYacqmQP7GOuzqzg4zeVEhaM6jvpUL+6UoeDuGwRXTGHcqc4aBEr
6obrvIh7kI7B2l7huB/+ZI70Lu3vqXcl1XY9TyVok20rQSfc8+nCv3mWAhx/Vzaa
x5MA8GlvlNCxbJW9/7agcQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 51376 )
`pragma protect data_block
bGdR2HiAT8U8K1HuLpQ6La5XlXV3RIrP7GQdFEy0Fcbfov6rPVDLArY4N8WaOXrp
hertpDadddRExVa8e+PTj2Aa6xhpcgKDR9NtoghfytQoC7wtL6U/xeDbgyx9ZbWJ
xiCKz7LMwmCTPzA044yXRai+0Pho7ROKCf1CvToqez+13uvRaf3cQcYDIFI9F/pf
xcQqBNNqd0yOu/PJJodAL7CiCkhCLyeEiEN0aoQEQZb9nelc0HH44FqnfpHXf2m2
sngpyV8AUc5nq4qHlYHmNzMhBDn6OLZC1kXkq01Mu/E4tYTr/8hXZaCxZRtcYctU
I7ZrwVEZKwOFn1AEvwkKFCC0gguNDwdPOVMmZsoIFepiEKffe70vMNTsuxpHlJ30
Q25BxATajQamJTfB47oP44CGFEjc5aP6we5xLWWKynkqmelaCg5mjR7J27lqWfx0
Wch6k/a2N/BTnF2BKWiJi5/pvNnvHJobxKy0FspeEhQIQ3Uu+KZJJ85gqzdcd7zL
D1VqLotzHNwnaSWf7cSNmBO6ii0DEAm863J/fc/2QlT1LZqPUFUhv4et0EVivbqe
JddYj+DJFQEtLqOG8Rh83VI7C/JhkwWdvb+MwCLYHwgn6YxXttsF3ilyP/PU0X1P
US7yInJ2dTzxZTPZfRc8WB2dZ+67XSkjRJ4WwON/w+7A52k0dakf65mZnxgcmTpA
CU3A3D60tgVeAUmqIc4Ngzz5sSzMbTTB1+c2X32zLOAAi1+Eio9fwVUaxOQW4eD3
jhgWAI45jA9XDAs4UfZoyIzKIXy8v10uDnwavMzjAAWE9i5NVGUOPxuKe2O8OQKJ
1eI1lDI9/f57UwxaEunAMT2ojZwVykFiuK/Nn3kHJotkr/SoQBrK0tUWeMu4kc/o
+N47PkXBAJHSyb8WMS+OOXdiXrRNs8pFbCcJulI0ZvnR5sgbwb7emAhWnmx0qxhM
0DnyEWAUFpAkasnxK2758saCBei4m17Yxu4hq4ya1KqeevOna0FSXdrOJq35bKRQ
7Fu031CD+iLED89ghz1hAb94KElm4ZZ7H2/4B+/wRmHS0ApH3P5A8+53yNV8JY/G
GGQSs+DEy90C1x/U4dQwPHk1VL83TGYbJFGQs3WSHz7LKtL8JU2Fr2Biy6XAuME1
HF5EuSoEJQCRJUf0hP4Xwi6uek3n9HyYJZd3egPIJ3u5gwccXMHi+OXXb82C+2kS
r5ayxk4zvnHJuEyquGqOqnjyv5pEhl7dTBp0+HIidcYk3lSlMxbxtUdKYv3pwhSA
/enQAAuhH7BzEb7HP3YBhnnvPcqCBqrYFPcFpiQ4+Z2gbjdhqnONh919S3yoU0eC
npa6rgawm6XojKLfzlUBRwcW+2ZKP9XhsD3teDuX9k4wdWdc3XDFO5ZKmHm98BkS
JFl2hE0gs7AebnM+ximpSQRz1oh8aoTz5FCTgIhIA/DOc+JEEGrtVq++AobAbFZV
Tekq21TwYOoSw1/abue5WzdDRDK4lPuTkXiXPLF4BZmh0UPH+GfAzWbdWcFc1jSi
/g3/yFKzpi44sCg3ABwIv8YkLDoDSgyT1xDMoBgp+PYAC19wIUTV9TjNn+Pnqk0N
lt3ebqoRh3EtYQc6eoEMFo6qJe7Ov+oKIopKS9P7E+L8s9m58HAw3+BJc05s8nNR
bqSCYuIa9LEG982eoX8O/xkrVCFnPlJ4Q0v0qn167Yfxb5FWePtawdj/S4ZHAMCA
XLym8hPfSIXt7QPi7DttnFt6/lVyAz80bG1wBYT6k0SRX6oOAf54O7C+gN4imGzd
imaMhbKDgHeMlTWAuPz8O0bO3o0CqRMYhBJOUW6GSEwI55T17qZWc638/Z3Rs9MV
6WAiXxLKgqz8eePnzGAG0VM/LbR4hZMYhA025MqmaVW+VUXx9d+TtFsvBkTe9rx1
+96EwTv4DBq//30+DznsJ1OIGs7KtcQpDMRfrAhXmsH6ZY1BKI8JCvK+9Edyafsk
wqP4fB9DMEs8Hn73KaYWzAea8yJ+AVybsLraHQbqT4YPPIwQkJl6MhI9Z4tg1n3e
KSgdfmYq/YgEae8yMrpAuOhId3qBpKUf1XCpHIC9i2Oxgr6baT5b9PjH/9e++Y7Y
t+i468h7f5hXv+kuQgmq0tCU06mgNs/BuBIsXHIEIDYDI7cu68aiD3lAG6vNmFK8
Xm39de6RmwAlNDQBy3qD+/AFOR5fi4SN7cxzaWiZQL+jqQCL7VM7mw/Q5M0DcuD9
/Ie0DZbf0dUncnVcpgvfNIjpspKSk5kGIUKsekPZd5+FJq3XH9hirF7hzTWCQgXZ
iF/8tdNiMZODbrIEwvW1zIUeYRZrM0l5lmBi8mN2CwWFsvjTqMxgJHREmkoJtGAC
8gNjZ/pq82NHyaAcMybfMBOl/umI0sKRnkdpSqzVlNf22HIjXotJItze9x0VfZjO
bXRHlxYdRiy+uhzW2f3iI/HQHhyoQjDdW7NDnsbGnd65ulkKtg1Xg9shcfH4Exa1
eVfs7NvMR9QqqDb/D9nE0EtIRqpd4B3NzJVEHVpT87smiYDwz8EFhqQYhzDbVGWa
+XRPyKjLL6/NPJ/2oNwDf6L95cEVeRSv6xQRXgDTKjPOV0ol8DBEBnGcCZsvi05F
FyBMGjqVQVo+hD5aN5ap1nh16DqbylDBLhRB2leIsHKBzMAxvrgg5b6vlGhZF8tw
MbAWgtvibG5uFpNRBHhCLWK7ohYaUU74FV9/qnN7uETFwwjHGMdLLDdOAFxN8YDY
3xtP93er0ajyfyhyZ8J7fAk5ZmeP5YZSiBXFUmYPWKr+onufT98e6g5E6Eeg4dot
yP2WFb/HgIpDiKJCGEicYl9LnAjrvm+WIYwUOu7cSWg0cd3zxcHpUODUuw1J/WGu
2gPpBCuqC0Pj3vqofsj6yUn7p2/8NBCM5r5PauZF3cGBi8VIPDJ/+6MfVK4Td93s
3xGRxkwxL+bUT/C/ewaFTBBrFNGq2Oqp5jZ+023bqBOuaAkbA8aYqqOotT/43zEJ
MlFRYZMJJX9Wve57En8ctWBlE8EZ/LzUf0jtxYSDAfINCJfMIH6Fk2HhLTNDfPF+
muONCEsvCGVl7E9PwcfLT/00k/UgvHVPlSB4D30VjR0io0idJWluWXmK+1sMWDry
caLSXqQWjPrna7m6+OEgbdXhFSTujuDwEt63z3LSkgZM0JfQJC1+Ntg7N4GjLGJM
1nU3X2FFx4QOL53hqC0l5pyLSX1FfNmadRAIg30XTqLyrIR/Y3SXfLQ/zXz2ikkb
d1xAozqjXMxp1xaJHVFJHjzE7D+X5exQ5cpQlrCrRkqlYwMU692BH02BBSXVdc0f
bQRPufj4wdGCB8kmQ/szy/+HmFx41yE4IxgSOxnQy8ote+BK8aJ2LFE/ZHMOzAz/
9ZmHd/s6sjFMkOluS1t9eX/MjFmC63WNv+59gJOXReQ0zVGzRfxsG99M2Z8ywabv
GXfWImqtwhoNNXrnXIk6ItGwi3h5iKuIiYfGXWG6CkU2Sq4avTgCK9P4p5X5brza
ZbJrivPv7SuzDTRVEtBdeyN5AqhFwGOK59S1hjH48e8/6QZgUfndROsg1W7Pv+u3
EKP1OAkbxKB2XopSJ6pD5A1GLnuYxOb42Rsqe+u/vUp2F3f1pSN8i1gfgCumLrAQ
evPmBvqCLK26x9aijQ2V9cTn/g5Ai+NmduIWG+1dd++r0g5TuLoFLIZIeWVP2h5N
PFKZrCNGjcRVc4/EmLRDO8ZDsANGx8oIQcWWgzZ+EUBwkYTrUUwxpO4F3UuzdM+Z
aM5PhuElvWqo4++KX84zYrxTAhzKJXDv29Fn/aIfYZP8Ab2mrK43k3uLMC5hNQcP
m2DcRJi722UKLGNUpg7tlLp17vRnktd55ptNkiixSTl6O1EDuULtlEcpg1BZf4t4
gSFhKz+2apA/Y89apIrQUIgUdHZAFHaUvwer6XjpLh250Gkqy8byqHBrJPz+wt4Q
nxh3OwaRHkLIyrB3rovlwf9eVAv8GwK7t984x599FBNdSNypCtSrCmlI13VL5bso
Ovr+og7Q7NvdrxAQrx80bQExg+NRqFXZJK1f3PLek021k92d2Sh4cXas6c7WU5EB
cVKFWsE4WivqnzTf4uVOjZsWKCyexh8gidNx8HbPi/dQqeTf62/Aa66gK1mnB2Cv
Mov12L7AWGC67pQKnaTnTPRE4VtxLy4/5Wu7XZL7vXDlOVHTBG8ClYL49gnMiYq2
EqIZWSLultHpqc4/c1prloUzK/pjSeWawaFsUy4PXhmdyK9JO3YMb7I9tT7YOpYx
nAtZ0BVfCLMOK0tAwKr9yDT32WBdfZC19sDvaP2+GXkojr1xo5E8SH4kzWvBs0bY
ZQG7lWepF/ZBS8Ovsha7vIEQ5dRq73HId8dF4kgyhUTi6faTgWvbPWvqrBbUZKKn
FbnNoBORxSPhsT7KZsWQYdBh06uOJtcUtq4mcpvxBwUqGeE8P7gfv9ujyZwIQJlB
sfI4WzZZ+vZ/bjbdOcg2/KMVNYyYvrb5qSaPVRQ+QO2ATRq6hES6GMMY3g6U227r
A2BUjN24uC5DnaeE8Jsl1867ubpRz0wc293JHWAteV1hqnRt0xO8UclQiclLzwrz
BO9QdNiYwtU00WzuvzPsrYSrH4aFf7bP9V5BNTionI8eOaIHi1600ng7D6YBBR04
YoxxYVZXsJi7P+4nDq0X8gc+dyPX3btvtyx6am9fgaW8yoOd85PploIi3ZXY+U84
n1MCy4Y/4nZP5k2SoBFcVYJ+QQD7QRZCHZYBZ1prbTNxAOIuvk0faY9UDJvZylj3
8Vacc3B3hQv6ePGyxJFNVMFhZpNZClE2ChegcG6wBUMI+C30SXQTzi3MANPwb213
UQcRQ9S52qaNsr1dIO//YlwNlDFoeRpWGvbT0Ly+6MbHWoyPNJCf4KVB3m0lFUm6
gqT1dkNwQYTzMSLOSSH889nzSrGVxsDF2Necl52G3dSPh0qLI9zcjnkkQLPzY8xU
wveNY5hyLB3kVRxduDaHoTCSR43HFVQITgGqMRTfVcQyOSqV5EApX3NdCs2rnmZu
q7klDoCt8CysgtDQEdPs6hM2j543No0GfXbEHv66b3Y07MWpfs4VcOJymjUFxUYf
Kt1a7FhpPGh/xr8kseJYgA5JWuDddrVYXCR+FtMpB+stekqTBqF9orc3/NyA5y1z
/qBzHqGbXoqPrsuXlqYE9VYxLgu76RYf91EYrIxd5GeJcT4P6L2aHweQIdlg0UgC
+yXD60EFkbbSVCGPMftomXj4VZ6bvi+OAx4IO1ceK5hcWiF5IYtfzihAeFUVFYMY
n4EmoeWJvaHiaXdZyvW17Fwm+K3tm3ioCzAhDkrKSox9S0E0RaFFQ5/w8vM2NIkX
Wab6HePzop00WMh8tbCPcTulxvN1/qEDkFHLg+EiBWz4fS1gYjjPF+8XRBx/EPMR
pljTC6yEzo5eZB7TrAn4fsU9KM/3Bfmuoj52v0mBZzPumvqcZE9nly8qVtmvm2FP
5RpVBiBFqFjYHFAzIMCcuB8BVqX/KSxqKmInWAdhx43v8jr1jAagP5HeoYwH2L06
ap3pzvvdn/VvDe4bAc2cWlKBNRB+9gcjYdfp0hLtxcYe1IYa5rOb9muQiGnoMjcd
k8kZepRGe4oWMaMK2h8sRn8cu1MIUC3oIdXaiBzS5c3l60W0hoO+Avb0kHEWYFIs
ast4zeYlSl9diiNo9XmosFwHlAXM5eUYfnyP3JPYn/8WuP9brnSnDaBQspsgTKUJ
Nl00w1LNxIyPmiQMuJQmD2fyNxkDO1prT9AXpV5Xw41s61W1lBTDML76Lis+8LCR
ISqlfg806mhIDpSjhD0bOsl0XhpP1ARdHacQj0ctedXg4gHX67qFcPnOjD6Q/aMb
7W9VOXOQ3SJg75mB93yBylpRgnY9rOzKs8fV47c9X2tnjmIAcZWaFomDGrJU6aXu
rpRmvZdaL5S+eQBryhKIkK07nXyg/abNgwweY+mfKrFiwYRqzbTRo3ucG4aWfqam
snjf9YGbWD8jVeNP3Hhhs+Jr7y79VvvgnuOZqVdSEm75EXwysv5+5CyDncYKneuO
mJpK/a2N1EQw+Ng0l73zEK9DmCciWYkD0KBNzm4u3xc1oceyIQR/r7fX9DPXiySi
dadBnRi0M96w6sa7mjpVbSZ9QGzKFoeLZh/uXBGlTyz/7onKaRlAIDXz4JiooTuo
bfjFGzeRQ/hR7bPzIPVNdCh9wBUe1HeDo/lqH3JkfDn0TrabAogWofseHhkV1DFl
Tn9Z6Oqe7c7EPB4qJ1+x0ZXts05FtfoScABL22JuWq+5TXxaMAz90blYo1nD4Knk
jAABtirujBNo09Hdh4V6wStFbOrobfnDYU1Bdba83/oXR4ZDkb4YtgwCNUlTxxkh
/EyewYvxYFINuNlefidfZT0GN6vTy0Ue1Vyq6AW38H+z6kUrwgqv1Tr/6uLj/ZSF
D8OloffoYqgreyQVtO9dL+MShQCAWuy/qSTgEzDGHalZQKbD3+GVbQy7DAU0hx7d
pZVKz5LN2e4tdzHFjCbOq5mcfkm4FRLB8lRB6gmFo/w3NTRPSF+RsVChSUZzcJ0O
9aUoC5VxhtPhjbXJRZmeTZkzyrgrZcqOFaND+LBLST0Mt0sWfKM8DcZJeut0mIQ/
StNoxWapNjO8vRSmBsnaf17fmqZloqFSyP1EJjNBv9PzL1I37n97mEzsbDaFQRpH
TucCkiT/3eGHBe2V5eNTpV962+eGzEATtJM5alunQsXMymwvhwZgJ4sqHwS307Dc
K5pTa/a7Is4Rl8ujTATKI/3R14QqXEQpzFiPiftfhupSHsc+TBYnLIFmeXOAgYPn
Z2uAZh+6EQbbfyw7P8kbmv9Pvam6NUWmuCisRe/kdriAU7i3nPyg+kqTjHri9x3g
4ltnyxSUsZsRPY1vft/K0lu6y84CQDqj/URyUNux0d3xZlUO7rTdPeZ4AWr7Lj13
+uljF3vXbMP7vRNi++ZWkoi9qXiLf4NO4OwEtHPhBepK3qrBATc03ftsbgYw6ROJ
bmY+MnH3yZQaiEoTdXNKQlxau5TSnCehytFrPzVv+b0FWkaEQFd041wqtil1F9QX
enle5Ase4oiLlAiKYR+KE+Dj0auJgBWTKbImw+ZXgVq44spKuKQseUDaTSvQXblp
UqOEA07gPgV+CFlmEn+UegtWHaj3IgXMRVAVrnjr0JbDb5sz1+yah4ZAH1hSdIq4
jZTe5qgH3BMexrcMnhPY3O6sQqlCmfziRu5LlAcTvJmO3Itjts92+Fi9xh8wrNJ7
vPTFsEGL70dbuiwXQkdgiXsHCc/6CvPjP8KfDuUKZmPM2o/Oc14Aat2RbxwLG82f
ZIciLA0b+JTnuv7ZDUymtH222bYzT0+GkMlHTfM8EYsRGpf+6u1/4F57MK/rKlmo
pf5EGqjc5mmfTTAc01r4UYVJJCBeg5U7cOAopL5WvykM4iPT6dst2WYWM5pGAM/I
QejWB5NkLD7ViaXk60k12gCtmYt2SGDjay78oR3HyeGEf9xHrtlKEXUS4L+hsF82
2IWlKF4bwmam2hc9eCl0HGMTALHrLnAatahkH2hucHUPYy9P6QbjjCAqzI2OQw/b
P1pGQaMw7DeecGmDbV3WOA3TWhuZNpdmAqgiim4PaYObSx6s39N3HaUd5mWCJBsl
ZokEHwZq9z32uXfMGCihRNGJphv+n80qqyoeq5b59IfY+2kVxjjTXDbmQjPYL5Co
RmhZJmfQ69upugZ8EoUep2cOWDq/IBqkFE9HI5j/JzfRQi5zPd5Y3Oe2t5A8vYzU
3bS4n/lybUE+ag0OJPvR0HRG4Ozv2lrsCxz4AZTWVwb0fcV6i3Z1rfSMGCIQVAdr
ifQFfI18Xik/DSPLCYjvSDfwGkQ+t1Vk9/R21RABv3D8zah5A2Y5pPqbwUSpws4/
sLibJyKJGw0mXdPkxG3gHNX1+WYIkg2fb5N3crxAtYZoy7HWTTDJmjZA9qPTKy9N
4OVXggbsY83UWc5+UcD89CJvEM4+beaZWB+AkbFII+yvKyH01KeLcNmvEoOLBjbg
mjTb/ojnDuQmcMP38RqXZSbDPc7gPBnyFsdtahbgMo9hFzfyvG1/txZ87+pkUl/F
sKIfU/07ba2Vjh1InLhnvxYSQM9ir0kNXBXhJNd/3oTS5v8Hp8u5RgpxwLJ44ANB
WAYOs1bOXLDySSDdHKRFodOKtcvRPpptqWwxLjo+0jBI4pQ+0Ut6Ch952pA1Kjwf
Zbdnz+ieYxMLhO4KltSFDPRByYH/s4njY+6VzyDUswbVDm5N9bSOilcI0z67TSmj
zF/CdKs8x4cmxatghBhteGguKK5MR5IpyakLhE1fplpLBSxKKVNqECyCRPkkQjsb
CO2Bg2+PsOis2bflQANLi7w0nvGU5CZ+BRjD9tzyVzhwH7KvcicAHlgOr+U7pQLE
v9mApdxSML4emWKCb8n7zGOYHF5PSiukT+D4A9KSU+mvuOZD9a39VO0/1Zgajn5e
dALh03W+t1wRrj6DukCGdEtr1tIbqTXpmfWEsseYcBMNaldNid9jVhG9a9Ow1Myn
By52jUPZfxZs746VU6r3OCsBjFCkGzoFMQy+TZzGjfC3hd14JD+mKwF97sMQLIjv
KhuaQRQMIb4r3b6nS2AZrRwwraTcTCd5UJPx42TcDFqAOGpb9gqZH+2kdrqbIznJ
Tn+SCbP1daG5C//VReqhfuDIs8QM1tlqUkIQCRL/vnKw2G6g1EzSeCOSZT/EKPnY
rhQKuxrCiNfi6LNDmBZQKrnUSjZgg2UZZJ7tY3MQEow9OFdi0ennjknjTJK+tc74
o2qix1hJVDbzrmAE10KqDb6zRcW8AYrkihL0i6q5CSd9USGmCKTwx8Y6LB2aqYNR
FT44r4zKhq/0wLEJEHwfgLnPMKtapaU2B3/nxEfk8+rElTbaRdwHaqXsfl+pLLkj
VTPcZFah+6wAL0tJI04Cm9RxVwYPbxt7/S4Bcuvenf6GWMyr9wDJ+JHvWMCTFsqm
gXVaIp4+PGeMfH4aj7Li0/ZdL41At8hPzU/e6pDOK/U3iAChmI+Bz0CUrrFcjQAr
NdmkvIrZMpTCw6Oh9qv4VDjohpwCuHUPe6giBQ6tn8mMREdS03OfJ2Qo6onllUEd
jhS9DgPxYCZ3LYsz8CVXr7uNiA9Gjv20l23bCit/2xZAft+1FKodpr+qMEwFk7+B
nLwkN54AdTaEvPDIxf+Pwb3+AvTXo/IaXFjnJBfPw3+F3Te9I/tkEDw8gNBfB2c6
lnVSqgcrXGQVZ3V49K6gYzoTI6W9OdvpYbr1AiXBhJFIyFJX0yVJJG+2ALdx3YTJ
MGLTIr1SEujMbmJP9p7xoLcPaBoJevTmmzUenQUfzNlCqDkE59uceAo71is+Y8y4
v+jrRjlPJXidmtWby63GQEmrfkUSlif4MOb6NnyaYvQilWAQslf4NMN0mTiUHWBR
+iHaPDdMs4+TIwsXtvLYtsnUllEit7eWs8CNkdI52IU7Buka9+zdT6cQ9GlxN4uj
5u6UZh68gvWb2yaJ/oBkABiyhxZDdAyaGlqqReEq2zWJhFMkZoYVEG4PLAKM8qOe
Y5113t21j1NSSJ3Vzmunjcz4sWs6kPqS4YK08h5J5iHJMDxYIuoTqwRLJmG3U9Rb
yZQlExfEODBrUHBB8G3vxk0sSYkrC6fjsEc8sYEQaDXR86IQQuMqoMcL8SqjXwD7
/EITOFIVPQgPOvpLEEo7bVSm5rI9Dpyof73aou3pEmzvcv5Ehmkog/AQD6TRakHP
qDpHl05YQX37YDjZxBVqyFj7KPSTmXASei17XdLGrnr+3ei5M/dSQG1dxfPT1t+1
vm9iQ6fY3vZvCQWu5yHepRRe4qiL6xydPpIYZhyOv1GGrScctF/+TMmoUTDzV4OZ
3RdgbhLFWJR1S4iLB0xEX+XHxX/01rqiAC1tTd6rUieQZ91wd3Jn1QKkuJeRD6Zn
PuzridX3yv7hvGKSSbaSDK/6zXUxHF5f2ZOezie3YMHoMLams7wWYBwqaPhsxcYn
Wt48nElhKolyKdF369x7c16MwEmxU29/2T9adXlJ6sMNON7Ju2HJUuM6Ifn7Zrg2
Pn77z1icehA68fYnCmLLgY299XlDZbo7s+VWrHIshheM/9nZr8fvQ7aynHQoAByQ
GmQmb7nJDKe9qCUNOPNrZWgDK2DFJwV8fVTloBR0jgrt0myUmLCK8qb5JhSmJyTC
s9fQlBhdBW9ch+6mAEwnQbO0d6YZjowqffNquDhMDWXmhhZLUv6tP58HHcXhghwA
kyjQcMQ8EpURRNU+uD6JUxk9K5zljExhWX7Cx8iv+A9NC/3/WhzMgjAhASsDDQ0w
afhdmAsUD918ud9k/+px3KIIwCSnWGF4vo0oMLzf9tG9upPDHc+ZtFbX3En4zVi0
ALBzLxigztMEBTfEbbI6wfeiala0iUDfPj2qaQB053GAnCzSESkSGpykpTgmo40p
8i9sDzAkO2RcNHPIuUlvGp4yAkAdLXDQW46Rt1P/mTt9M/6BnMUyd1Kky7vpg5d8
5UIjRVjxO4lT2Ah3zuuJMpsTzq738qiF07DCKd3fF67MkxBellMId+2VHAKfIxVQ
upyoptw/DZur0VHQEXGjXKyAR94AGYwJ7PjPTqIo2pWEWEH0DsGZkc6JZ2LH2+ws
bD/U4z2+F0jV7WOra6kt70MZowWIOC94Mvf7PvB7ebmZSBWoyJ/K7LJdjfB8iFZ9
4jaakLG+VT+Px/LrcythU3WYuCBdAYQvESmm9qCDRIzIr/hUGfE1SRl9t/mBFNFi
i80UO4l98VYgQzFMBLUTNPw/Du7CX7R6XRb/pvaw2EzeUL1slB9FKCSh8TpxHGZi
ZBPuaIRtt+Tr5D8U0sG8eDqcKdt2k24LNB5PrpT0lej0jtTgbnto8cGBYgA0PkFN
2iQj1YFcQ+4cMSrw537WKRTvo2ADg53jBn7iHrH0RVK1Z06eCV/579mj7YSYPJ0S
gLCkWO0+VyI+orMcNYX5UsJaR+quaka6I6fKzOdVJAXZjEQypg1xA5hI3rBg1Jg1
HQEI8JfBsutT/7O3CQuU5a4iTYmX4XrbEjOTQ72BVQEZAelaQBspcJlDOS80jYjt
Msu+TzrWqT/lBDOt0ol+eQr5p6WO++JVODjzKREGOrB5JfJkGkOb/mt6ldnzEQVy
pIrkMKusLxonDJB2mGQ6gNt4u9CABnte/bg8rjAblnneIaIV0avDEoYBfIZ7b27a
bYZ+PQDAHMLWRsVAVfT3ymM0aFbGKqRrD8vANfc0zB0ryZYZTjNyAf8k7RoQT6H9
uZ1kl6AG3sYoAzP2iIsnZWKiLPKkRy/vOicAvnXke3qJTO2GPxLsgxgYhYR2oviB
Vmi6qMboVpShcdpUdXijKkmeLkrwUM6ZnhuCQ2YY1KOifbnfnhiWwj3qiXUEzJuz
pfTbf6RT3v5TN7i6sFTSEDxn7Xw82lO/ts/AkbjwM9MnuCl4Bz7YEqpISGvv8tqE
1z51u/BXsLsDyuC2MgvBwjBRfJ06yZFqb9cWfLUnPrUsr7wyA221pSyuBvdSqyXo
k0byRQRAAkMnaO8Ysx0SroKopTq2ncXrLDTZuzkre3fFuqaB/9jjk5p1jqphcoGW
gUQ8UNXfeWqsjV/shA8X2RPPW/pdgyfx90RE9p093SCnKYnYnnSt8Gynqr1l8KfI
PRCYDsD4XGOvVvK0XbHJypVB5nsBJ8JBPryXcYGZYvJerVE3WIhFXFzm9CNUir16
TxjmPR0100m6RvjxDyceO7LhbaF//SOZOmuyxxhamx2R0G7wlAGyabUTyGtLKtah
c0LyaJT7U5o5G8tqKOXhR54YcT3NEkk1G6ybWT+V9S4IEnE3GVfKZyONEEU7OLVP
sXEHrbokG6Hf3J+jqvrs0F8y9yzHsFZh3RwPQ0v84d/6N53L2g51DyutRNVyS9sl
PhL/V6Ka3XmpjF2KtupLNyZdNYjZd1DQUvLtYCK8c8mtUdb0ZhA/dnclODk91Vxl
g8dFP2erTY7gvCxorCk57IuDvJoz0PK/M+dHfqtX6AL2ggVmFEJZvRjL1JzLLEG/
36VasXIZoElxJtYemOz7QqMy6JuXFmmLOu8FCQKFR4so4Mf+IlFnb8JwMbz2RIO4
JjSGGG4cnMcBnBQRUHc/JsT4PH9RwVD+TD/IdEsZPrKTLhT4S3YpS1a3ryQTQWTq
sk0x9Yc0Wdrkgp0XcpO6RGM7opD56ypZrTXrzds0VRErYUtk2YxX2QQhV1SRfZfb
mvtvZB3xMGP++v6ld4TfsKyQv6/ert8yQzLeSMuoDUEAOyA/hnzYtM62n+3XlgIO
f1baVBAgsH6ClEQakl00/6q/zVFzeEjZcFzifyfFmG0STczWq0fejORajDoDIDfB
XJ/IKI3QQPUHzh8RNWqpdzH8qJm8t/T7UxhbQHP6XYdAp9tyBDHGuh0O63vu7pgO
pACwM/J+bRbOF6ccK7WBRmLG8rPfmeS0xAGD1yEFTSNKESx/TpjI7UpvWDBwVvsZ
7UeikSYhnkXn7j53qT43q/qSwaTOrDCDAXt4zBXev08S4haFXWE0KlZuNhQ2fo1j
v2dcHTlM+Da6Yt6RJclWC18XvX8Eott6XPJ4vXzttr/8ZUvf6eomaPkWZumhvfKx
WQuLcaj7zYGT97RHdjh0DWq8wqhzFil7hqDdlDgSePO0JeilsMVnZsTBzCI4mdgZ
gLdzxS+f2EZOJnCh9Cma1vggeDT3jYmLQwqbNspU/W2vzngosyYvilU4kFUYpT9S
XkdutOps5EZIhxGMYb/XB+ULduCvfJU65ILUF6VfATz7ZSpDJjU1EH2/lD1RVJ0C
VX2jiELByil2v3gdlY0HwaRviIC5NMLGejBdPYRt7wBRg9RUha+OU6MICwhuYNSK
e1OLDaWm56S0DiHUXvYjhGxFbJWj3IfARQwSPXrMwoT7PvtQlFS8BEN+piOdVC8J
Ba+td6b8GF/yQDpHvCHcO1F65Vb4sZdL35RM8VnRD4Kz3NpaWXH/UP0wnK8eFdIX
DnDT74u2OG22QsX7bnA1UJbXdZz1bCvvTSRFwoL5L2g3FqqAbg/wzv8EcW+Y5r1P
hdgx3+/u2GMCsiRBg1HtArcEFp+ujHL+ttPsebOpP58C+s+N2l+NPems+9e+DNDE
ljA/AU9MhIKkUB/GJ6z9wgs4APHlOoIciGPI6w+eNqoOLM8f8HLGqfjVq/C/QGcY
Udg2P5oPJ+QByGLxSdqphXOvHrrjt2GRjgbI+5Zf15G+W1sEZ5OBWtG/S6eDYN0D
if/6g54dSVuKtM/knncNpONm4YjkWxM4WCBqR0szzU0fhk3YyJYkGELB99QDAzT0
CFo9JUCtTGJj86+oCJr4v6QiQsMScJkvBUALZW6cPvxHVf1a8Mw+IUI6iv3N204n
g0GKuTrEZu17skYGX91CJ/adWUHF9vY7909kCh80gMBOHuBDEHobmgDaHulUc2ck
LhfzzY0a6D88B2Jk2siUg2kzPLnX65FV625u8PVmeGs1xH4r0xlm6xLyACjqrsy5
I53QZaJF6aKYbDrKlzxoy8z7pbcR0DXnGy45W0gZc7AaGBhAvxrR79yQXesLxOI1
dh0cB2q9K5Vyf5yw3yVO5L9jvjEO2NqThWFQM8dbyfSkHWoZZVHmLIgGVJkGHsID
21UPeG90PV/MxsDu1cNDInGlwLG7oRAH/4l76lDusgmU1O2NhWKf+/loewDteal/
3JRfO4uJlrQZ55k5AN98jy/xxwYf3PA6DpuRomdhE/UO7rxgYbSBLBqKWG3PYHFo
o8wsL1X7JVSYA/bojULdJJfsgQX/mLJG4wE4WT+eCf4Qw0oFEOUqyaiVDK+xijNu
+tzzcYwYFlqW27qBBSbRoEtoPBUFa4zEr+kxtOSRKkEuyR+Ici0DCrD7+Jy26hIZ
78Z8x6R/PCDcIA3CVef2mYRIAuSgiJmh7WxMIWCKJmLvwRVpvEG3DZsfoLnJsfIE
CQV/06WM30RogZlFhcRYXqfhoqaSepajAm3+Uz2vFJrYNFKZJ3fbDKUmrWkiWnIU
rko1bUs5vcP97fYyjgr4hcYDi5hzU1yBzSp8ua9dGSDUkHmZ1B7/2NPyEgZnLVCB
fVibRzNA9TY0MneuzHxdO/qvPXTxwabalKtP+a6/cG8dHe7whO3Scn6TU7C+wZZv
GVGSKM/MZcgKm0N+m5GRLme2FrqAD7QoTZ2iaAhE8poNDGgpM0R5CYxBPsyEH6Kh
aqWkkL3BjlLos0fn/ycOQghqM8xBQ80VwI0OAonlDzdDtp6X0fauauXLhuvfFuVX
acZz5PDtQtJdhHLIkLXcJoVqCP4xTgvKvHRcPCypoS2GdM6N2hkuRNGt94cZVD9a
zmMXVjGKXy9mXKLG0QuGc8W12wp5zQK82yfiLnO0sW2Eu7vZc57jFGE7uk4Wq0i5
WxytQRZnaKPCnb2CVpHkVdTe1aCLNt3jFhWZr4UJT8okQT7cBxT/VXDs6+7oe7dx
7Q4Zf4vDz1pIWsWyaNd7kspHsm00GVfc4YLTqHKaK5F+TclOKsE9ZRysThQxcnDp
m6VVo1YXL63LG983US/gya5zc5OZSVzgWvQGdxOw5DLRoI8D109/HP+moIVTZOiH
ro/VKZk0QmPEASFRb9/vYcVO3DraxcE9Yd9QBFNZhPtnvp/Ehpn/eiZRbOMl5VG+
t/O1Sr4HdPnziYmIegwFIJjMyLF1aRmXPyTsXcBQpHTZu8ZVFYKKfkvtrdlgCsOP
1AzLP4+MeZQsX0D6HNR8F6mw3iOTOL3MzMes0N3e2YzwP+kMhoCHv5o0t7ky4lO0
fMyPxzR7SR4WcdDCyM/sKcqiASG8YtT9GFqitihRJMBtblXJgr6wthdw4jfwPdnd
qBH2OhYdW9hJvJcOHkR896QASH+s1FvTvF3vuIsX92KxQZfuedoExy9UUhjwFGTg
IVZzqojHtljQfX5h3/AzxsuC6ZcJ1RJB6uoipydv9B7CbtDOHkFDEZv/NUDRVc52
cLfa3waFmVPTdBZQM3OSnrugrNaynSoE/qUvSyLb2mqHV6KwGNa1nG2zZG/xvC2H
qyUp7SUTbJ9AwUq/ZgQJMR3L/iaLUVi2Ep2RgjfPuJjiztGXrxNZZ3taHu9iRoFy
ky0XyCR0J6rs7emqvRKB7NHNvEhN5TQcLTHQqzregNz8tlDwlzDalG+fdCZeHF1V
h8vqXBRjn90nBtmdVuHoenVyk09jWf31YO7PJyNt1Dnf6PbhBaSkKLYGK/qni/U+
2/h8b/BmpIfB5z01NGxVHUU7ods0ygdxCMeRB/VLqgcbNCn0YTzlqN2FxRXdB5oi
VAs1VtsW/baldlO2sZiLc3hQPOIaF0JaQGmVcPxAVKh2HY/ohEIjPuuTeEKwuXTq
kVTc9TcNTl1cRh5V3ob3DC/p3QE+CNRBgk8+HmQl9HlU1DzxZDPh0EiFyOcbbAXz
dJMWLcx3tIVCRjzO2KnBWBeVfo7sAfH6ATp5pg6FAi0kK45pw/6n1OxdHLl+eoDN
IO5HKfv8ymkPRNrVz/w18nhFWQC1vTLUDLAUPsNpaYBiknzO1v48dl8/KujMKx+F
WJFqfP28QJ0NPX8bPiIrL3EEBtKbvmzprhGwiMiuE+YFqzHbKL0YAT76L4/7WY2v
TMxlhn0fKNUUxDkRaQxEXJLrlDiXeoamE6/yF0dxP3dAK51aU3B/hotaKawwaTNh
1QrEcpsEEzbUeqNQaI+Slfoz66BKaMkkO2r30PGI2alvNWcTxfrKGX9LFrbTNpOE
Q+dboBqKKNVSsOtLXhD9r4t4aPVWOkW2Zg+6XKt2RCSaCQj3TvZYa/EKXlLgQYQ9
t3MAFfxlxARKQVpCxdBDRchBGP9UrZMsCT2u0w1LzqW7wDv0yX92N7wgRtrVl881
H3xd0jTm2gWmBpRPhmcSAz2D+V57x5flA2FeyGAGpevd8N1fk28nRXkIvZjJI0HX
xHN+pi9LsV3lqPTY/RhFYacGMDSyZ4rNECkqWAnRIq2wDCfDeKKk+kwa960cfKcl
FN5KUp/PUCUBEaQnmS6wqVtnH4tF6uiHmAMKFj0eR1wjC4gMsQMHDGlkIrMjcohS
cIrxBGOxjNm62iJXF0dBgWQPyqa8f0K/HXJpNKjaZoWn1SNXsTdTGVwYMQBs23wm
pEO1yZ31mMhMNngHUnVmdl/JXla8sCI8ALmzkr6/CUB25sKC2IbApdPAtdErRucJ
BVRwIuIWoKS5Wo10rRjTxRXKsysJGV3gjdjy7+y/0x2pFYYSC2/kM93MfoYQF1Ud
ISSeETGWUUrofT/Cw0dhuDV5gY5KsMSdMda41Rl8aeUX8y9N8bGJqlKwaYjBJWZY
JYf2QTczF09/W2648x+QXn/kvJlaXHkUk2E2f2Z4vXc/z+oHRBpsuQzwWfGbxuhM
tfIPLkMnl4so6OhlCKGgImyTEdr9NfrjS45nUZQdvz9zOFDhG9NgtllbR4zGIjlU
qvg1oz1m2pHFr3aH+VoSzRI9yivDnt/SfygkT6CKKiMdrGeu3KNFBPmRFntTver1
ODnT/3oZst/4qrXFxuMcmFp5fk8asM9fcdHbR5KWp9VtYoBrlwVgEUBDyJAYCjB7
g5gZBIF+3m2VjjBsWEtF1dee5nEbLo9rEj/q+weRdRGw1avjz1EhzWkAVhZVCYR/
XaD/9CqkxDQID0NMhBerp+mRKfSuk8w7ZzIkSGZDpoURdvBcPF2uw7M87JhQzY1r
PIWzkjlnzUlSxnnx+JRCorQp+1rGHPzvJSmhfshw4AnDC/rtu9Sg6n+z+CFp62kJ
mAWcOCuwTMYSpswKMV3WUYz1vhCgLpM5IqYQ9VzVz6XmHyJ6qsd6yMy5ykGVizrR
U27cXG5EAAdTLO7c1Er3PuiXtpSHLY5rOtp5wOY3Mca63P2PDV3BLVUTvujANM3A
oTuJvFt/s+7UWBWRO2HBd3SV8T3yvjSYb0SkNmiLfkf1jz0Hx0sMy8bpsteNic5J
BxMEVsobdYwf3gAtcONkUD8FCNx0G6IRIcOyIhvVP9BizraduIlDOBlNnIlfj9AQ
GQDyh1qBfnQJgNsWj/ZUeYjwcPgg4IVxuA2MjkYgxjQgC9GvyagICFEDym194Kcq
WtG3GpwtR/iQVuprkL7ZmC0kGS0cYWEk/AKSQsLNouUAwoU0Pyv1vsnUeiX5rFkj
1OZeSuQ++hfU0i2BbSXbQ+Iw0xL9LeFBkij+YFGKuTRKsX6LXiZzz/JZxtOQ/eKZ
OoezL1S3UWgjolHXYEvhcTJIcorLSBzwUal8KrMFicXF1ecQR9JYtfaA0cd1ZRhv
ilT6YWHoJ3iCdsJjmQijTxou9Hao40vJHrtxGib/8HqPb3XWJmFAaKKQTskG5aAx
OdtgzD6zeLPXYlWRQbOCYa817BNXjSm2luzB8YGqejRVjWBsiWMC/GTUpB/soT5N
4pYDXPV2fKPlN/Te1gt7Fg+yIri2aO/bJ/p9Wwa3vDPQo1FGbo+oLaOlA0FjfqY5
kGH7G/mepk+yThG17zCfqu0sGWGP7exoP+7t8dUtiHFl9HSlwQ81OgiSQ+Xuw7QN
+CSQtJnKM13gyPXFoLbxiHxAIdgjV9emECnDF7rzWh5hEQzTFHLYchMGz8mlavjc
Di7HgTS6ZYDdCfBW49OAM5ebkF3Ec10Odf2L8sE0HDMxWYz+eCiA4zD/dNp9BGu5
GijhFJge4Xl8xteFrNF9bklWfO/91qxmNEM/KXyCmFfswFeZgnqc308L+lcLVRnt
heFHdtdwtBaeF8RaSYyjJcG84TDa+yjiKZwQiStBpkxzZqkW3ok3YLvUqDNAu8oR
I6Qe267nZP6iAvIcJRGuaEdGYorBtj+58O3sBu1SikYmlcch0iB5gZ341/96UVm9
t3dn9b/C1jmNDeGxT1v7KX2denQsiiUQkRuNze6wOIqcIKX+P4aJAgsIo8AGKrWt
CVDIYAxMCs8OEavlP4Mfu58iXvMkWthqrEocfqbuFiO5r/wmTY/ybw6tNKfBfob7
DFAgTt4ALX7FBDXCbtwLNgCTiwIrK8oWNVsenLLLn31ahSQ9Xz6iVutng/OPfUIV
d2aLn3psc7A0sg3g3ar0wGq9GmubBE+qKZx74dRZ7NsFvM+3N6Cu6Nf6uZMbxtDx
YAlPKqRpvm/t/my3n0nYg2mprIU6K20AkRR6jimhKXalgfQJCNJqHRN71SyEYtPy
2Mp2NKY7S3Zkaz38OqnzLaJ1k4mpr1ghTUV+fyu4vpMjZWDGTuOhUeatuf7nF83D
hiCW3caMfmLzLeiI+5vOpJN/86IvNjHVNsKAvyG+T06+mts52WFISPZ73CUDKKPH
8UYbxeROwiUnIGna5T4gr2ofjx5XRicwSyVfsXJBVbGBOSn8fe+lrgLZ/fDimEf7
OY9vi+kKonzACzHVq20y/I3U4iyRjb0Up3StfoLDMnyB4/hectFHVppH+4kmHB/i
QB/57DcdRDjF4g9kvqn186zJu7TslgfCr1Y0svF7ngfFa1N5CZLD9SQxLXY6Qccu
/RNpZ2aqD0tniV8G+o4FM+2IlVlDJdzOQ+Y9ijnSBabvpUym4RD/th3buoz6a6ok
dDrbCtxfON74eWOtdyq9gY+p6lfJWBo6wgONFP+NrTZ1MUddDlr8bWRsxZrVO5f4
0MwOO4VIHvwhcbYw9IMfmbbCo1md0N2PJDjdvFx3iAcBjd0aV2QyZXVxS3lN3Znb
k2GYW/p76B230jHGBI2lm9aV9aV+Yk37wA6eeemdYVdSk8atFv6QC2YhGHxdrDPU
EgZrBJ6VpV4nNmcotGe+4aQB/OD97FQDzyXGZ6+O7NBi+TwSMKamuoUoTk5PKqM5
Yz3Ek9ofCjzSWd1JeXjm90jFWM323/GjkbQMQt7gDxWAv+futRD4XCY4geLPqZCl
68UME6EuMH47H25GPZRD1onpD3usowybAvpasqLriWQyEe6PcreXtUqlqNiLtSeo
79LEKtAfDxAH73YZg4ayfXVpgi/yK0Qx7VgT8hGp65UUIrIR/hw0NByjedlWtH2y
HWWipAgYIsYN67uEMcj/mrUSpFu3cWNZm4fZleQ/aaTzMb0TSndZXoxxN0FGW8Sl
KqxavEa4ef1kLn0di6t4BFOox3Uq/xXxKznbj+fL/J799fpW7wdF9ZCocA/pzDQv
lA0dFjiFMNW3E8Cv3MlrASvI8I9kn/UNBmsbx4sEUAi/VIC3VKXNL8vftDKEUH79
vJXhpyH/aluu0Ceh7bESgESNbToLs7LzoIdlzUgzwat/OvtrXheXBqrKEc9Q+ntb
OWdPl/3YsHiVSbClSYDgP4/WLvi7iKr3zvqePW6I+KE4j5qYQfwCORYhGMk0+1hn
8jeDnS6esjFqppn/YWdSZcINxDA6Jjh/8StvMaRtTAtIhJ+UdtEyQQTS3lYO135i
NqQfXndJSskKxbQbOK+jInc4gyjW5vFx7XD3LWzQZUf5aznXbggEVZ7QzkwOkBcC
mK/QmMy1JnDyAQqugIIuyA+Mz03gZf4Ao5Okv6mu3VpH1rI0lAe0/9HrIJIS3Z2F
q/68pTmN8F//Z/nwzNzS7MLtj3MFgpV3jSWaPU1wyZ3q2ntjnhljD6Lqg0NtXMwP
Hg77v609qJyvSvkfko1i5aijOkkkTzcBxXrWfGxNmsATTxoEzFBcgAHLn66ismtB
Wqra397scBOctaAepFXOyGtexrepHJhGCGhOuphixZq3QUClrtfzK0oicllq70hb
/m0VA1T1YoykxxU9iOjTz8eH86igJdGP9atMlStgF2iFAMqcIkz5XGuDIEMjxgJZ
vq5viSDy7IaL4e0OC5oJZzFn+ou3W2tsBZdC9BH//if+JehZUY0iK2jYPWS7g+am
ngkA+dshOL3oxu+iEQh3pbPD3TBC2s7wvwtLsGL09V/42XNosHmWpJhdLrhDEDvn
FzmjhvovS+zGeKLwRPEgKocym0s+YsrK+41gKPSvg2Vny/FsTMAHrO8R8zVU5V6H
IWBUurLK1X2wKM1vHgV6d2IZFClcNbi+7QoYtJed2GZp6PK/enUNfq1S6val54kx
7fA5uiRR2j9z3LW1Hels3sTXBq7K8iF/9qCvY4vx+b44gHkwa9Ql4Xmd22RWymIq
FD+SKtH1SnT/6xT4IqOuPU2Wa9PtBgGayFBMxZ9VeueicvYWmyNFFODgffVC6g3A
iXXx2KkcjLAT4M+39OFvPWzUpDaUwLC1cMaR8UZqM1Cv1JAAMJkLmCXjUtF/FgrW
NO2nGr1ncR014S8OwYGGRZd+DPIq01hFcLj43MX/E7WJLbJt4SZRC5VU6tD3Zz/8
9wQAnkwHWoDsdX8nrEYF1F0v6qfBI+Yfmoo0VQhfVop0wltfZ5uFwdaS7ch7Op5D
qup5IKztio6xvcQRL+hqh4T0q6jE2D9NMob2VdExtN2AXJj7IlJVVlqV48KumvhF
XCyfRrIwnIPCmlpKApxQF4BsENlPf3pJD9NCnCCpwXyxgtU3+APktLOPU+Dn9FZ2
xaztEEWfsj/MJPS+0wLn5rWpjyF1iL+YvNdUEMDN2dhjMnxYZbP3QS1ZwnU2otdl
TsqAmfDnky3eCz1wBmxqMuVbSC00KRSM853C2UGBcoRXP8qsQ/3/xoNt+Ld0czGN
i3q6TXKqFQ5kNYKeyZCT6AOwk3Hd0nj/ymr18i7eXY5JMtfLKcZCfQiv36Ggnlns
WdjJNB0u9QgYJ8WsIWGup4cw07mu8f/MmECJxQAOuqRUdXWk8Uqpc00yiYJJMEi2
yNrskS+DM1xD317AA3MXiVq6atl1pjAw2ldJ1EiUpyPb6xETwJ0GS53eQ448tyXN
vMFwnKDDoMLhGlQf4mpcSj0qhY3lWF5+tRKFxbTXSnCTdNiiIVzk3BiPAQVJ0uSZ
uuzRupWzrjgY8GZ/l2xIwLc7uacWmJErtiIqkg8EysP7iHM5Qz8pT6z+BNYlQMtS
T0YGkpsPRV9sAhmxednkSDNVe/kR9OYQB3++9B235J9iT/ficguLUeUw0qlxgpMP
p7jLzpL0bjXenfmB1qA385Ws5VgYeb8d/8p1MqtSVc0+9JXdEdBZDvmh0+agxoyu
1KU5xR7lWm7pBprjRzcBa5GoZPU04ZcWMZqSd3mPJby9D09N0JyiH7R4uZ6rCU3s
nrAVstWtoSUaa3b9axT3NeykXx6z8EzPOxbrjbbNConMJXu1FR+NOlgFb8p2/Y70
7MaVjNsHLWscIDre8jcXdW99bie1Dz3YzEF+D2HbvTHWYd9ihLAiH7F6bZpznjWj
7xkwMAjZqx2z3mlMYNbbhtsQuGiHNDsNezYB8ppu2h3G0+02/FfJdLUpFkmp9DcF
BShUDfrF1JIGnG4DVRq89A9gdlkaBYhLKVvc0ikmtUdRmtWzFq5B3j/Gdoml3j3T
zeWvYaEc/lNP0gdpxlwteO6gdqChIAJ+2jyjeZKzDbbNMWK1s8bXFCb1WxHiLZfB
kQDTkLW4+NSZUvYj0YWZyQPhuxa6ckyphbXI5prgYcy3YpvptC5UeE6RRzpjL12J
fEb/F9mpbBUspWshgIsddErCMO5r9y5EMo43ILNfoQxbCoIG/rAPvE+cMLsvficz
RZ1KjMyj0JnL0vAz3Z36fA0b81AFBtg3BUMeIsCc3T8ehznsXLcB9QHwjQkkmPok
lcU9HTAooskhlyHpg04Ia8pksVsq8kjOZBWGAa0RTonIFREJfvUSFfvwkYQ1b1NH
GPw3Wie1iYs1wk1JTdyl/7QVtX4MKfCT+9Ur1rmN4KuSyqL9YNPxmYvNx5CaMisg
8wnlhYFHZFPgJWG3ahED3VQdwn1dsfN35Z+gy4rk7+uO3Jc9fE9cPHdSt0cnZxHl
DvutJZXTJj2jLQwlPafU13y4tkqWKrz2skNTTygexYdSR9h0ZR5YV9JMZ8vMNw5R
s77KfPBhIKsjR9rplSpoF06fbdtHzcTJgEH2Drh6oNMPDHS/USpYMOkdmUIbH49B
Z93WD/+f24SCBApLJgiIECOvyty1zEHjgtx54Fr0fE0FXIOHY1jzzwgbRF2is2S5
yvw8Hzgzl+66RIm3Nfi8CAmbGwXuIZRLFaSAZJDU+LGdw62PpBfJOm/JBSxcg+3M
3cY78juHpJK2wsuio+hkkM1baG/ypLCDwuDKW1dcpdV7CCBa41rns/U+K9IGYCX2
ei3j5oV0jVE/+TSPN3WTMA9Z1p0voJ2WnbwX437l+AGmVAYKKS8y82S0roP1EWKU
6dSvQ5Q9AXn94zNK7jMlocYDF9aNh40K+91+Cei6lO/bw1EjMWLGZuA1CUpPRdwv
/mfpvU7ekU3KXnDeOrKs/+n/rkrlKOMerQdjzoe2HUo5MY1Y465KEaHano1yfnnS
3u/nfFCPS/f7IqPv91re7OhCvezW5V7tL77KgdQg6XS/QPxeZ++K5kRng5VADxzv
nr1A17sPRKJB0RTJEGW3OZud5vfA1bdlRnR0qE0HQrPfzbeUhCfzjZdiD5ywjnFp
TRPMqrZPZ/JHZ2lKFcmIZBoPEfzyJhjNoQdP4hNm+Sb9x96s9ZplmfDAC0izMcEp
qFTJ8O1mYHTFuZGOovrDdj4cQ+MvGjcPCatWR8ZQmSUNPhDf4SBj7m+IeGHNdmD2
0LBOD7n53cLy0XVMBgNbR4qPBHWVYWp8TVPeqDPR2aQ+GW0TMqcx3PM1cOkwsX/n
skEq80tVlMtpnpVVbTSRPCtL2rdA0Atr8j8HvVrPZa8Vuj56QIJYysW+QlSgq111
YRy/6NAUPRC4VCgDPJFqNzEA9Yx4lPkAJIS/VvysISBr1i3V90pB0558m6bMtCy5
fC+5dow4l6k510K7ArHwC6jENvRtM1CsiADGoYix10/GPrT2ECRYTETrirKgDRZn
C72ZuzuIMmSTVOMCn/AshFrMmn6uG86gMDrl3t4GZbznuaFxLoAI8rGxqgqgR+un
s9gW3ZvQZdQ2QMtawIRQTpdUUNlvHBrfAD7HsfFlCBJrjzRmTPjDbt9LqZygyVjP
CIvV5Q386s3kobfcKiWVCJhPRibxK2lHfGii2Swxm7P6hDyorhrwZ5iaGXMO907U
yOoui/TEnufhVvDeyh8L7UZTIQ3pVyVLyhHE+VTCm7VhFImdmM3zBB7ezAeBajo6
LfIOch1yrhrhB4DNhlyQi9c02KF99hj5Kh86Df+vGywIYFC1w3airdQU5JpOksFT
WwcloFrQXyC9qWtSdPexyH590Tomqepvsgo0DhkpH4u4Mf0FFS+dK0LEihKBetOp
b7G/MmI77Uu8uq0q9ZppBo62T3ad9ZqR9Mshvf0i07m/awgDc0ef5u8clwawQTBB
CljufFU2QPUpy+6k9zU/Mrt9I+KQ+lKu9yL078T58KbvorXdk+2pSw5xvdGWeG33
KQIjXmryZCaHGozlTZmEsRGzriOWF3Hn2HcDs1gTAkLzzULQj5aD7WXnvIL4LAVA
lS9BLiDy4fWJ4NCQH1OjAtf5HYe6gL9v2AlWjFGurZ9al60e7h3UldAdFETO0hPV
9m/dI+CSPjYK4E09gYTlOhdmCHAvgu1S1cHyw2q5kl+VgXWD7DEalOlCOlLOnphs
KblQofBFTJFr98fAL5POEVKhNtXzMAX13NROFXKervU1hJ4VvpEJ67Jn1y2oZKNn
KHizFvl/iazYEAFZGytp7IbgyHA62e8EUuOdQw/9n4sq9+s9otmC0eMWM7eelpEA
tkdVo3C2B3jeiypI5Sd7O6+7zGjuhZBFe2rUdQ3ncHhfIDPYEHQFssEWNGfdAiup
ZwK3aXOhE66+gsG7RGiaNmtTADjni7xY4YeOPjDUt2WDgK8e1CWYKqWZKe0EbMLi
dfg9QS8IPnBp5VXYi5mx/5V8B0VIe7NIQzyNhncsP/5yUJ6woU24TIYa9T9u8nUF
yz2aTfrUbuuSPtHc5SqkSBgwU0Ch1+EZNcsbk7SXST3B96Csp3LRcx5+yZbzB9Xb
GFpagGtZgRHwE3IFczmQWqR1mJjJodv5tDJGVvEQ5BYPfE2AQ+K8EIOJYMQg45o6
7bTJiDp0JAbscyNUUZi4GsE49Yc6b5Rr+zhta1Qd+4OE/Hx7WSL2r2tygwISSJ7Q
WG0a7rwBfRXnLNhvNbKfZX/P5X/NXLKSVTqgbvL2TdOq/bT52nAfkn6Qn1Za4aLW
Wuc2IRszDkRrflXjCGfU7dX6h3GP8C8MA5BLDfMLPf11aolgD86SnR9yVZElNniV
8fd8ecTbO65frnIU/oBPC9hM3XjRabx/md7hBR9M+LoJPm7eHgAsL0deM/CB9pqG
Ss2W4uToYAqm2RDpu6h1sr+jaKJWYlibr0ahasO5W1oa2CgCPHsOA2Wx5cZer7N2
AS897HmqeGyjGk9JXPLJVhv/Cz2jJZSxGKWstLBUVIhw/prPQHCHx8YrC8914120
xv4vo0Gck7fMepbBHbtPeZ9ZphiFPJmldCSSdEiVSVDv2gxditCG7tSe35flFnnY
axght1vcE9QzqkNZFWCRFbaxtr4MlbHDkrI8doGcgJCHjoGEf+RTWoZgOR+YJrTc
zC5Wv7ePCsNT+HBkfIpAYTnwLZ10l5jEyJW/vtt8aihoYPeCFeeqkNELLAImUppc
NbGUjY2CoqUwPVRzQWdyDPq2KAtUhVo4mWAi3CFNx/jvm4Ks25ZAKb7SBwnLTbAH
XAMgfji8g+fmf/APMVJ7GKp+FM5IrZde9TWJ2hWMSWhdL5pR+vrJMcEKVhwth9Bd
dByJwKCTZd5ClRf8qq/3QPmHJ1B4ysq8KDaCNu+98W8rEkvehy1F7HZMjJCOs90n
i+3fkXTFfEFrKHzYH9yIRx3c+QU61r9Ev1/r1QBhzOvYc1MBvXev0RpwJi7swP6j
FF4rIdOZrlrXXO3PTA7uGCvnTL5ltLBLuWRjkjOOBEjBBHCVFrsG9tu0Y+n2h/E8
tcKHANOnV0gg39Vgfi0S2RoldiI5isHY4FUFSTRY8j46IyHzVhMgzUz4pBA5mUAA
NrKiQcFCUdqcyEzRR3u9W20xZs071dgj8ZCqsYLpG/YrKiUEsHdHnmyPJValq1oW
80k4frGRB6b2eTSi8IVdPic0DAhzqCGmfTmESrFM5fm6ThywzT1KUBPQ9sCGbsHD
wdLSIpUcTo0JrimWYXhLQg5uccghLJbZ1LCetC9XScr5+7k5z4gfC6wsCJrNaUoi
v/hNKTj9mHNTDF2GMQvT5rZR1BxHec/qB/vyLWxJqcICRzkjXY2c2UW55EONRe0W
1DSfn16ibvL2xdFm3pnd5ci3+NnjFf9BMvxuuV+bu3g2OaAyKP9jlq+J28HDYF+h
h/UxvIX3funMQTV5LwgvyoxtdubmdRsWdZvi2LwLn1tddZbZhrwYKO674cEf3Uj8
A60hpbmVKkYEy8XJ73MPb/6BHZnfxWRqqoYTP97559BJ11j5B60TwI9ZqC9Gzd6G
h8GAhlCRc0kHMmzHmDElO8G3snldXcLcNthUwjlx0xRYCqcEYszjdd31JNr42IyF
5p02dBs39bn0s3lQGW1p3KtU09HwwBiU5PC8/FHJTCKzrFpMA4AE/+uJo4VN6n9V
eYdPYiVUWa+HABFKnFIi5eZt7M3A7GRPNq4ZH1G8q+nMiWPjJz1mohG5CKG+R+rz
l7DBAGSu1trLWE44tXrWWnO5poSbq/D01WFvm+aDzXj/4hxYWlBYrUMRW0w/Tsd9
MijS7urevE9Y9SF5CEXe6oj7h20Zorf+WtrWGEXgOJ+vhVZJbai+w8cStGWyuaAh
KEwcqJOGznuNzm5KTmpx2nnS/3RFQWgYIndnD5w5OlChfh+tl08/tT4qLflynWAX
6mk2+vYTj8ZMIku4sAllGcyqaTvyb7oxGCv2ByekfJ/lVdVRGTp52c9uF2NsGLMF
eEXslO1yH6Gyo+Zlp5ypfXQepxW+r4Q5pEMK2FmQ/GAwycaaV84TiNc1zlyuD/ek
L0qLb9+b0DjwmhMQJ1qjLpCk2jb2y/9fMv6hiAR//75xVRDZyjYl+maEncnxXbzd
QIYgW+p+CdNjk8r/DesZ3icLgBbuqYzjSVJZbWhCwl04So2fIO1dAuXeXYYYVKsl
14MyLaXpYVo4lmlhVXqyyNDulwkzFGvgA26j2w3X6jcYEUcy/LDKLWHC5LjSid3C
+BMhgzcLUjTu4UgVB+Tgs/NjX1RAAKVtyJULHMw9v3fbrbv+lY/PS403FMsE+E8T
v1iQYGTKcbd1lkGlYPCYFFxDmkbkXfKYRoAozWtTEXktusgZUQNiTTET05L65avb
C+bPM1IBkoMcHclRuN4lqQpgaX9qLg6yCuFxjsuHyGlBS3fweTi9kccgV9HMDvEc
5U4ClOhZuprCAamRiQtzBs2EiNh1S9wnUAqGwe98sjW+5UI8bRDyP1+n+uesh0hj
84oKIyW8VbmIggJhDRRk/AN2TRRmkuc8OmK1E/nf/gXWMRl/6XhWdiJJ2mewhgbe
9ORrDJFi25FdXVSPy9/AJtyQ2lKaGbCSXtWlkzPrJTeP/fJGa+A4ccI/2ZrNTJJP
QY0eEdiouqm31MY8mIC81bvFsC5ndeJabx0DR6qt7L4jC2o4wPte+a+wvxPlVVFF
av7FarnJfPRYXPWKfz8R588xhxVbqlczfV4tGSBEbLcPLaxkxv3W6HwXTD1haAGN
1t/hOYJzsePk2c/Mb5zWBw3cqmE3OLfPEkovX0Nhp2yTgaunuH6hTnPNsFoMvVq2
r4djZfIZOwlVzlG92eKPXZ6/P88LXVpf17IGRDMnvSp1vYZpsJri83Y5lwh2czZT
CRaRWsMTDRX4fnGwOVsIQyBL/NhSkiBudNKH06Ei1HauOB4BdSUIUv6yNv1m3PSc
AqZ4lkpzV2xnOJJWnGlzvii8LbkJTIP28XXTE6d3BKvdwGpOc4Qv59Dt9Nv6BlyX
1LMRnO5QLQxyNreQrcGlpxXLBQHz6V54u/WYg/bYmPx1ykuEZwMSMtqqZJ8Peac5
WCsGZnzoZY64ZHGhorSB2nMXlNjZSCDUjyaJkkT43/Jcxy8NtRKAHXYgbQjk5Nk4
EfgbbOTOJMZRJAJNgHY/U/xvtfXkAWA+drzOXRrxXpdHmLUw43/NewxLpGrRwM8w
djXFQ0dV4z8nWqgIvO63efsOsMaaJbI0BRDoPuThUtZ3CjyXqT7HR+fg6eBQsiqQ
5OGIzD0LVGpZQpbaod288Cge9u0cIUceBIdCVJo7b/6qH+Xjo7pEt63ZWhgmF/2k
S53KERM6FSOVIlCNwCjJwX6xNh7Hs3tRGX+oBjgOXMHgz+WR0fPvQRiQl9ccVSwL
NE3HFOHNpDVJ2l2F7NhuvfDHdEZffxFJAE/JaQumllJnnn9m4MQ5jefpxJGIJRtM
LHNjAhHBuK/nOoByY0fBQT3gmv7JnZJ/QYsngAp1Ye72zSRLKs5jTyF9tLAylGdN
wSIEBgpndOJ/GbKgCcBy/6fPlJdICLjBzZVNcBBDolGDgcEx2d95AU0SPt4TAU7z
noNI7nTRV08Hy7Qa5EU2uA7IkotvkT+RP5//EgV8SPDzDnjVU85x2Ev6ckOLGLKf
8nnKCPKtD95bPl7K1lwazC6zDrHtdrnE63Ilu+wa6mXBr2GZdWZkog1UbPxVCyf5
R8lPOmMCS0v88ER4qzi/VLVoJhyYybahBCJaCtXpCwYxJRYEfV0zdwpWYXZXVN8S
xFXelDMwsAc5rSQaTYKTVjdkBsWeRXJ1+X/Z2nRqDtPI4oSm9haW+D53U+0rjoD6
Oau/ySBzONcDg+2rfZqM0Q9oYSZfB4NfKlkEczSgZxV5qXOA7zbZApOqAe6Eu9kY
96XWLdyJacVv0zi4WYAZAcRSxDckzoYO5JiE7JBYAtMr1YKv1q8+pstsPZ4sYqd0
dbLda3EHTvqHiX+oOtZSms+W+vQ9xUnyKbjD93IaGoToTj1u1QMqgmVWSckv5CzB
AeX+sy8rTDwugt8CO3pr8eFUtIti/CkBNMA6tAlIk4nud1PY9acuJ46R4BfCcOQw
rz+f8hyK5EW4i6elaAaKtSehQSaiCz2DEfi4sgKu2ZiJgX82V9KUJprGJEU3Hqi+
tETZf5+12534i7hBcNWbK5kqHDM8Mlbc36aFsr5suu3w8f+p+1AZ04QK954jIf96
m7E+UkU5+MyrUKX06YID+7xxcvpD+5tfp2+IBLXSJ72d8kaRrZXiOeZ2kQgl/2gb
BIOsYKop2OJPCUn0Xy68FDaAyy8P7lXseZDefrYQK57yM4fG+ih5nF4DpSVFBpmW
M1V5uhp+jEtPAHSAOBWc8Vf5WjvZP562N+j228WnQdkkkit8nQ3AETvukgSj5/2g
dD2j/F9s7AOjhucQFWBq7Z12/J6ue2yK4LNBH20veBAGxyV8FfJlyyfm/TlI6iCb
B06VwCcUb0Q47UpXjpNx4/Toa02tuZZBtOXzcgvyk7eX/6huGIRO5cFF6UMSgnvK
udUh0fsA8NcFERpk/WQp3VKPbtSVV517l4fEh+vnxu9iEA9j6bxnuzIxdF+u3IfN
4tJKXJ/qwuUn+nS0BfJROW65qvRiJcBJoXeTts3J+lQZjxc1S6wOhF642ecYLXcF
fERRNwZMl+6UqTUrzBmQhCNbJ15i+jDZQvA1Wqy4mGiCvyjrfM14lJ0YvOHsclNk
VBA3jNcHs2oLlUt+0x8s7BePVmO03to3iXjqCQ5NiP6v5VIOQ4/qweYlbhCMe6Ls
8eQuJVMaP/aUQmist8GlZTuyGkMZPqEYhxB2YVrKgYW5jQ3AT2f9XJKvrq0Bg3dX
DVQihsQAwu6e7N+HQn0wHFYT1MmUElh31tf8NJrmrpdG48n7W0cWhhjgmwaRXP93
G9aVBc+kqA6CJZCP3c7mfVa0pUfum7/4SfnJSFze3i3/XUb8hHtEVV0auBpo/Buu
iudo9NSdwAOeLZNp9kzfwGm+PaoZVrKpd2NuD0Q2Dl6vLWNIhekqoDRZHo18Jpml
F4HHSHL7OHinF5EJ562h1ATRK6DtgC87mRfvD1tJjYkw0CWKB4Uq3XCGbxCN65d5
NcLpeClnPgWwWn4mEOVq24ROtbw+s5USZpMSBO73zFbN0D4ulfE1b3LoJP18a4ht
eVDjAU4CN5XBO6+4jOhdk4S9LVwp9XgIRPpkNsLSKp61vpwcDtNhpkszHqpQ3uCn
aLspJM9sN0FrjtRoPymRcrOKPzjTrqMUgy2rjbhRKrAs7YyaMi61+UupMd6slCPu
HKDdWIE4M/a58UsYIuq9zPBMiNEqIZYJfjDHEMOx3q7c/QrSQojxtQvdXcmjP7XC
WR1o6ErXWrwTr6dpu47Q/yr2r0BTyOEbkLJl6kosVpgy3duYxs3GhYcKiIUu9pd1
LzDNNCIyHuE+QkIgCIG4Vax3Z34mc4/NtrEFfgNnn9yvclp/+CFtM9IfC0UELfE2
iBrvxVxnZBSwOgYyLjkaHYypBoI0Wn7SI4fEStYTEGw0FFkQUk4vYAYTFlMbVpiS
2DK+BfgBioolma+EiarwbzrlSGBgtOrv+Z8RRwB9IRz9esPi4+nkDMM18yESQd7o
yMaZHK9et0EOML5jv9CV4YAkps4tFiNtPVUMX9QI958By5BAgsmc7Zv2DWiaPUPO
5e+lZy81fep2ruDKHWiOAlEkv9KnaM6kRjm51tLCpfatonJl9eG1QAkYN+2OsQuE
5MmDvKSQZDVEMrHylYd7r/KVUNeMj2feLdbtnFep4SVQWn9UzEJB7vXTRtLMOhOF
mqkEahyGjdHYdaROqM36/2AqMGQYWvdWM2XXmAk+t/KB85XJLK1P4avu5DMPxE0P
7Dv3VXcBFip3hI31jyox6M1tdc5uf43U6BVaNvfiXL8fVaEW7FUa189fnZy7qNyZ
7PMsWZdnfDSqR/77iOKOrDMG0fIdJDpIrB4J4iUyNF673N3qBhsDnPeRzVpXgpSF
z/g0RTo5l23iaqQuWSnCu2x5Gxw9oJ9z/8dycERE6AHaYHig3fZb6uaoqR7S4Jo/
cSushab0MPslglMNv3KLFWw9NrRqbHJZoa7gFBx12qJvNQQ7OPXbTdOWFCQzi8ID
P7tMYch2u4yAWAEUblYxqlLqyAe3JBT3Wd7McIMOGlnbv71fHYhL45W/I8q7BjwX
ZeYZm2W1KEw3HumoDvJviU9i0xX7rEbmTWXPJdde7YldGZKqUfUplcEr4YLLbDUk
p1Qs69QG/xcalVJcfB3SNKQTTtMIQbU571kXRW0Lkl8qZSkL59v2ubwrdbSPc7Al
RdP+75vpf8NntRBwHavnZmzAqf7WMe8umBkDb+vh30KBi+H3bj31luKXmCc92c/b
24sbVQ28oSobXeu14w+aftXjQ91RWxmJMOR4QgBo6TaD1LaXGtfip0MfKTAnWasv
xOUgN1JQyPBMvtTh/i6sUYfUEyxKsxDOFyRLoEgB1PHxkOwfIVDJSevvjvV5Sr/B
655X7NILLTsp4KRRGAo3W4pFn8quq0maii1PEWGFZtQp1tCOvr5lF7tO7QuoItrX
O4KC8/+WkWbZw/vsmgXk8vLgUiwEDHbCf7Z5yEg7t7w6A+V49Y5tqSQrhgmSHfr7
ALdpM5Wr7JRA3rUS60mFUX+izIN1EkEcr0tFUVr5nXo48XKFGkT8yExkQj94Kqv0
14q5OGofF9C+MU4vvih/rE+URnn6Fc0gkplunJzOUoGUyFVOACMHh4qGvHHwaJEA
d/0knOlmYp9OyvFRVcngazwrJFE9hjWhZop7mGmj39v79zPfRWPncUodRHmtaF2F
Z8j6RY/EWd4xFwiPoq9SFs9/rPVv6CKuTlJSV5C9QOWtkCERk6PQuVCMZh+xo1jr
u2kot2agmFqTwoPZ7cbqNLhs6KwHDF1mU+0fYrkRNjLz6OV2xlZpSZRbKKuCjo3x
8LZi8Tpx54QtZIn7SkEJcv6qJuuw4Wok2fLJ07b8zCYoe3rWHe3CZuGq9NGXYgQh
SUqdal20XNbuqT01nhbPhOPiHG3lgeu/tyuJX83uhgLG9ZnWOgbNkXAozSqy4Cf1
9dEs6TnmmloMxqK0lYv+QTtoJX1MlR1fkbKeXZvnFoLhufRNz2ZPkg2gwSiCeGsZ
hjAscN52p2SNEdgAffabjDdzrt/+SIsCRZjEFY8L23vu/04/cdz2CZ58Pmla0GHM
TlgdUixV9WO3lCZ2WjVOuyWIdzzO613kFMZ8oPzwfFDr8LwRGOOGH9kvqmh+9eu4
eASfQxLm4FULdLkXwvMbhEBbvBvE166rW/UYPjRwepxz6NVxqRoAa7XEycxNUw7V
Z8tJUa4RNpwyyKRMcJcgDeDXzqy9XI4Fe2Kq0WiDecaVhpH1g0VKUTZjxIgtqwJ+
lLBCgcoyiL9jVpa4VU3m212JKmadbu3HMJjIG4rF+AcMQZo+ZvoPunJ81WdKbJxI
wLwn1WG5BOPzgu+96w30ZR3ITMRVUyshXtBVZj+X8aQQC6Z2NJhqbJwaAYsXEXkM
bx+9QebTfp1cm1u0XEFm6Yen6Y47uJjOaR8JWdwHi2bjW2wTdEZqlkWpcSfKR49A
Q9zeJkZgvMkZDQESsF3zsa2ArUUXFAMJGANiE+Qjbn5Ve8tDdkwVm0eV2YwpqRyJ
e9VdyHwy/Z8dYAoyT3n54lakLl9CGcwFMADPHM5N7or7otpNXnLuxDGxMZZHuOiV
YwczbyGEW1uYG4n2+n1/ap5YS2dQ8MzEbRppcrFu356J5sH7+JdF48NBOduWZAdM
jRZbSJIQLnrlYN++VU1twpXqG1BrLuvWXzft9d2XortDpTdiEMXyI0IHs1Gxo5mT
FoW/CAGSsSBMhSdMAYab7PH2J9wcTAc2JkrbOlDo32Q+SA4oa/Vu1xTN1u6XPkEw
53KoNZ6tcI9106XfXFyOlHMBxwqxr6ki3/PmZNWrG4Qwv9IHHarvKmuiHa5VRbb2
P8xLPjYJAgdHzMMLxWY2utgnAFl6ziW4HSWFoBTp4FaL4PetS171MqfM8QO6CKBW
iJ9V+6JTk3x1CxSfPV5RY8U0bkHEQp3xqtRtyf+3gCHAddXobPjPLMtGSwY1QLW0
qAFqkgoy4ACTTgZjLjAtVLxMvRo1UX1j9tm3KrGhoNy769jPNgQUx1S01UzeJL/D
lzljcmmr8X5rph5tNZSHNFCvUJ8QHWYaIweIkYS5ddEM9bjWHJ3xZ2Zivm8O04NQ
EH/j9EIkFM8C3bORyFyuSMDDhJ1D+8T6aNbcN2FE1NUyn7Bc3O9HOem1aQENBMsh
UHJuBPOOHBR5T5fW9TBxiJniQIIoG3cd8I9xOKbG7DPD0Z6gAt757N+wtzbNxvT9
4IN4GV8d3Lcb3unrH7mMnOqe8odod7RQOXyse7KNEddLFnbioMcTVe/vM/cTcH7u
hLOcdroe1/7TuKOiIEk7Yqrjz4iQRW5Rl7/GrbHPsp1UczA3pNOVOEq6HACzo05h
8bPK2728PQ1gujcniQf9BJKDduf5Rbr6/92I0ggFBvePMkUacwTbpCAcgkxz4CfL
vbU6xJMC6Y0DLMBPPtaQqpMbK5j9Bicq9HjXlBtdJzuVfeTxSBhWKdMo5I9j6Ro6
ey4zdilVYe/t+GUS+UsNjKZwMWeRU86W5rlLR6BmCfRfNZRfhQx/FL7sXzLAXHlN
prVm/s/fmDbWg/dCH0HchW2yXXRjO9ftWCJq1pSh73Xydo+R7luDHfdyMFx831r1
Qp90PbgH60ZIlg6HqiPCeONHHIz8cB0cQJH57Ocq0eTS9rVTnFOwD+yTIFVVsyWM
kXvL4S2YqxB/hj/aMm6LPHJk8GKXlhN8hnKKyG7CnIxtOCWvJPQOvwzetXi+BCOW
HyUYfewFVxnfull/J4mfoO7Q8zOrOlBWxixaHzSsAa4xzLGJWFYpytHEt5M1d28S
W8GiO6eQKTPjjg7EirXJZ/CbW4iws/PUWPEsZkLXQDH7Wvhf/VV/Z559q4jM+VBy
WjKqeScNY3upfKiio/uEo3FIo53HH6Gp+n2yYONRsxeeufOdNLT8mBawCqPmxTyL
zhOhMsaNiVRl/7H11zt31iJP5+uEwsq+TlBmFh26RiVFh/tGd8+Wq70cdETGc4k4
7C4fSm0EomwrwlNbCcr+P2Br9wec0bGBghn1m014Q+YcaWoNLVdxK/nRTf+arH2p
MQb6A3dwCIfa03NtN9oEmIhLblyO/xaQ6jPwE5BIL3X/a49kPohBi18W/DRNIav9
OJtFflenDRzzEgY/wmSsXDKQOiNL5vRSz1JRvtfTQyYhG9EJHZ9yXmNhEgVDokvq
UHMYnkHoPG7/4A+DXcqp/wgYtmlnlQRREEYM1gUqJhNfZvdfK1frYYHnjTe1BRii
IC7P3fhKIQcVklGewe7yS1YBgAmGfG057nDX2eeAOH5tJsb/FmUu5xtk/TqlXY/b
ooRVav9RxjF9SpJy2k6vkN/VvnDTNdk6tKf4NtnlXqZKpzaq0ae1wp865smMiMYJ
nUYGOR6GnjJILEDN8j343OgROn1aQP3WEqZPDCJsYkaDasg+SZNh8zopk7wjXiT6
eZJoVXGkKg9feATvNT+0LT+SO4ZDI4Z0vf8RUQuGTzt9LN7M53oputj7juj6PIRg
F9jBAcrS99QsK0zdGMWOPHgYj+1HNRBwIW2vNnGf16yUa6KLl+7w5Ie8DrYpNFZ9
r6tDueX6hJr0+8RdpDGRgpjDRmkfW9cbI9SMhmX7ivYmWbuDoQRQTAxLGlrkFDwh
uiD2JCKJFcTc95ntFYj+UxrPxNf0KMKNIITjbTWhoozOrgM3SRo9w8oyqRRKML6R
+97O13B9Vb1saY0TyzVwlGe4MHEzO87X5v7lj4oePH53KCIem3sgQQIuLvC7R08t
wPRaYBnvbY1LltmbFfuSeVYVcXhCp/piHFEpye0t6xH6sj2FKXIF3PjoaocVbJAT
ctcfzV9uunCQmobI5jsZ9lMDu8ZIxAwn/oth1LZYgAjBO6jry/sC6kfbQvB1V84Z
rr2P4Ojlb2iFCi7AlvjpkBrVwzq9WcnWUBdqT3OdSWlMwWNRpx6vY44jUW6NnmPU
pwp3BHz4aYUReTMjmfsGGlcZR+aMmjVBTjXv1ufi4xmDWNUKOSqJOPfm1Ti8RbxA
gAHB5NMcJcPxPBQAz/+jVqCLCnVN8VYUrG8k22Mcy9Ge6HP3xYx+ZSu48LUhiN5k
hf+s2KIPHcrH6wEuzwBREmgYDy84QcrSWhyflDbfP75o797fvq/GogX0sV+CRgi+
pQS3GTTx3SqC3RzDdLgIxSPOvaB/siuD1xjyUy0OM+NMoKUErhg5wztsLpzChjsE
ZnqDwj25HZ28p9AS5WtlFw+cXK8C2PLscWS9b17YhJSfu2l/tDCovJfxmNIBVUVC
V/IBUWQZzFu05yUvgCodKkotM/DVnFmpxwa1XzozowtRKF6e6wOIJWXyxugbWqXF
be8xgRzToqZAn2MG3vrg9Yx9VTYzoZ7PjF9wqu0J4o2ghlKSL3j6d7F3eCxoc52Z
bEd2EWha2+59EXzBLJTN0CtSp3m9z92efHMt8vg3oKpdScRBARDEWn2n86U+Yt4l
Mzi4Y9hd7Zjo9uesSJlgHezQIasfmwrvGqWaK0KQYCVBmg2t3V36qFpMiv/80b17
hcm5PsUtGTx5j8Ak9OQroQja+8YTD+SWXEnYLTVO0YJNSNTcSv2UiLHWvtH15vlH
TyezwMTtDLt9Bwk9VPFGcg8OSdap2aLEiVGKwPy/IjfUD/Fhe9eNdtqW8roTJTun
vihSmxfPL0Avjj4CRholRI9Fn5ld10Wx9OFwifvYJXiqZ0B1079+RRriOr3L1pqU
89t0Q1NT7pxFduPvoMFVE4q+E7xtx4b/v23Kh4IJBuh/9/LsnWDOzdBWLWf6xdQo
sywosv6QKl2tjlpM0Y8bpusWLl83tW52cngwNKWan2q0NIaDjc1L4G/11ujHyZSh
RDvwSvwwMmr8ljdhBen9AW5Tno+YiLoLfK1J5FeRMW0MP5yFR/xJDw4f6gu5QcP8
HOCl7UBHvJFzJwbuSysbY54EAvVq8ZVxhqs9etkZs8ptUVmrd1tMLsQimUSEuLC1
rn1Xh8jCbf2X9YJ+JnZ8OWEO2s4SzpKcqCsd9Cvi2MFTzv9XzXxmnyzBkKSNhPSx
gQd3odkWNJREGz0tgJXEDn2ewkUA02olerKZZ9xEL9uZEIKQiTwt38uC8auUeZFn
D/EfkT9V4FPis6FnssPYK7MH+f/oOWfdF+uZgeEQmb11x/U1gZKIYuiKY4Zoan7o
EppeduuJyY4h9a2hrVuX1wskfHZ3iesXMksld1kX5daIydf0OjqigMVPNl5RLVmH
BVhJ0Zerm2GE8pokAhtiWm0RSbLV67OcAcOAeZABehLDR+ejnBSaDEH3A8XXVWsT
J/gbVAC41BiXEh+ghyYlzuga89vAqgtvtw6dZJxv6hFSQ1YzOfamBR/+v+7Tf6VG
izBmatC4lYL7ZnpQwl4vX6fFLI5kA8j6aESxJB/AyZGx/7EK1B4FMXPpOnDlcidr
eCfeULTPekrIkK26qgtKgLURjpdJ0N/K5ix2TznU9Oxe8shXVEe8cTrgeTWsVvSg
XjlX5cPJbhCmyzkbmVKvjMmWVdrqahEp9PFgukao1q0ZfVw7FSUj1I8BhjMhxHVp
C0Gb2UTIwWdG2pWtC8bi05/xPVripHfQBxHx8okKf+OQWb7puPPo18aN1TtceRQ/
EFJBto6n2ky3Nk7kwWaQzt50vyLOMReyiH4Sx56xzBpVlldAvMImfEyz9H4zzX1z
I/roEmeBgHdLIYoEzYUxuvNjWSw00IbpVwfvZc6SDDvOj6E+5+opJJ3ExQ01JbkY
WiORL7Vwwc/o8auVibQrTwzaZzM7Wq0lYYzdDJVTXJGkkBF66ZascrHVzjL+gd8a
3m4i3/Md5D1GpQ43omsuIry/mGkCrsTh27ZBrWojzkZxzYcSNdSug+ixAIc65kEZ
trDF4a/92AdKGc4VsIvNIjd9ZdGgCqEwvSb1z5HsDxL9cED5x+tPTKWqbTrZd2c/
aAiSQ7ZxUmWR7UZYl9V8hwQcQQwggn4z+3DUdxQzMQpwXRs46yd1CsdRtp/guaSJ
DtxUJtM2XMNFGX1lC5Pwdnb+gaKmdVuNG9jDYSFesDNAYeKZ7FVTTLSg0wBZhBpJ
p31HOzcM+u2xrXaJTpaveyO13buZ+sELR0Du/VuXLZHYFT/VK175ThmwY+ooTMCH
6o2bS8XCiNa80GU8KvW8rQ3ncDyKF8U1ey7hk6D22xo9MSoGW9yd/xw5Kv3woOu7
xC4Y2qNpsdfHdH8zrVaYx/7Y3w0iHveBgHFReftaU4s205h/4UVjXy4nUBe6Ao/t
PSdObir2cERucYIztFnK5et62M0WyLNFVw9QLaLVvWLxAzjUD2Rh+XhN0jG2pt9K
D6OeQ1XYFqzCdN/qYH+Yu/QNt4vkzguJ7fBRhgdU4OZzqwlCCJCDt5f/c/S2w+2P
1HslF/GUGLRNsfJ43yDmEvAgsKndMuXTyCVhH6qvdYOZmTxU3LB42z0EQqk6j9/D
RTlncZJMD7lJOi2XrdMzVw2/RhVQm/71NU9wdlYZmJ7+ZvZJHv7Dy/xqCTnbEpGC
YQopHkdTz7GecJgv2Ucpc9jfYDMi2Q9EhH0CYV3PPf+Pw/zUitek3Z61SVvcF6Fc
6QNIDEbqjkIm8a5oru7VsI6jcTyvVUm88OqVfNOmHJFQx6E3QHlrlZYSMXjfDQfM
okxvBs11l3oRm8KBC224J15npxIp5ipOKQ8cHiQjrsMqnNj+dK3kUpiqB/TGxGP/
ZPpWOUG14khpKlcWTqOgy7CKZIYniIHtf6hevdb43vd+gjYKncO/BHpJHEytHGEQ
zt4nihC5RkaS+PTNpIIkXxBo9luiaMl3IHuXryyIICCQcS5/Jxa+u8vJjb1CF3wZ
T8kIoHRJ3WxzHZFRItbMm/nKw9EQ9ecOz4y0+DK2kT2Ni7sB24SG8lKUVFbXvpdL
sJn1T05nBsPjEU5CSr1v2h1E+MKhxZ0HqPA48YQrVq0f7KrhstJyj3zysr7Q8Gwg
TvyfLINezst20BUR11LQtsxSgzKZUwM3S9f459N7ztDUju+llKsWz1uCrR3sbtrj
TWOd0Qx473jbzTVHYNAyGDU6DfThw6tJFqfhUwDRhsNHC2qF+kx/fdYTxKGwqbzb
5n63SU2pOQ4kyZFtktndyLK0TlUXNrdaMv8tyTnLHk9iI5za+l0BWkGWxxTJylK9
xZaoX2p2wD9xYlsHfRJ5CnRbV2dHxhrswNW4qfyaYM2KHisEil4C1u6ZftEuTJjb
8E5IbDagbeEGH6XcQlTd0WMo8swoJYg8gSez0lufjvatlahrxtmjUIsBxw/goaG8
PIfOJToJXteK6Y0orOUuxvEAicxb9Y2bmWZevbuMdKyaRitIPZVpmKOMP/0HnGXZ
1JOKpMb0uBZ4Y9yRgZo9GscimamO19xmhtnc+dL71oGuaH8qO8kSs7NiiKPdcKBp
I23QcrGooIUdyH4+9PjUNOcjaUUZoHrh5KZTZ8MUQA99zClCQ8v8AgOj6G0O9Oi1
wQ63uIJ4A/b0U477shIMubkxg5yG7nsDc9OXL7xwSYZR2mKuVURk1XexcfKzE/7Y
LIbnMsSQchnm7IsIJfzWwGbEp3iYAmEsrGDLaGt3OsjbxqRPCzwOcv4OriPIRkNn
AnOl0iJyHAt/yBmAqO8I+bGEL8zffgPu3otG4Sw5TyCdXH5FtS3NeJnlgXU98q4T
OrC38ndzx248QszwQ4EK4JDokNfeImqg8vzrCUI/PmA/rzhAe04d+qiwLQg1jCOL
Or2YCGq5U7pIOcTGgKMUIUkRBFGmgLVnQEUS0qrqxxyZLQZRlkVWxFldDJb83hRV
fbswBgV0OXviUm0842lx0kqIozksSthj8vCS9xtB+Qkn/OhhyXdqHX8BlJLetoU6
py66E6BBxDKDC4bFFbJjjpqBQSfCCG/j82eJGdK+q3huXUU7ClOGoCRLmhPV62ZU
QZzLsYYZgiYNhGDvMi7+GGYnL3+XxOkQCKTtLgRaCEMaDjfxBNHwMNtV4zmQOpPs
R9d9fqzzzBJZ5Tx4Dt92evcpQT7hQNif4cmUE8GUsjfHLOfVBwKP6ZgKU4C7W307
nRxqhe6OumhxfEZuHXqa+aeduA2MsgLaNLsn/gUTohpsBYxlHFTonoNSkUKeqpK0
qaqnSeC17fg7JIxp9dB3g0/LRXO+457zcgcT2xH6djEW5ZFOHwbxVbGRgKMfWEFC
+cUD5Bo7gaYQuozA/Lnd9ba76g8SsBj2tLMty01c2GRmZEYVBVmplqrqlS4zyS5v
YzBXaoksvCJkLAAJxLsFQbykkYzBDBosJh3lkAa7bzDEHkXPacOop/jX2ICDeMEA
lUBMMTWlMwrrofexPpsBKQqAJhZoqjaP31jBFIHbsfo7i4+tE52So83MhTNCdtQB
WhrghK4v7dt3k7dkvMOW8KyjoedV5Qew9ssJdQ/FzrVtKiQNtv5+6Yw8EHGhHW2s
1kpYX9wWJpyMAI4X4VJWzTCRaYqUDfoe7lDx+If3dYW6eHGc6VTK2zIJ7itcVuVE
3gF0R39Sn7ZzXNjeWq96SOxOUYVtMdSxvkavEt0MwZ/eAOmiod8dH5l2PSMdAkAb
W7LWxcUC70S8UQjTyEZnrKX7PXmzFlC9I0mv1yTZsTXxBguIDcLWg6GJ/rPFdNyv
bs46sXj3JPWX7Tw4r0cXPhr83MMEWlwbBk8kCiLqxwaQ+43TYetoYI0juRG6w4sn
G2ZCEsEZReBJBTDHAwWXXdnyyIlkv8JtVZiifPRGvLG5Nic0IPPCbJOeFiRSSuvn
xiKNkQPmCeVdb4WjfKv7sxmFM2p4a1Sm5lDggb6NQCpdDTaMBrmRfztlJl1y5acC
UdE9hOqEX4w0V6NvNsY5xZGbphdREG2uSYxINQ3BCLk+PD+Qfi5HhkianNaNGCyc
KToMEXITggtuWcW5Dkn5UKQE7BR5u8VFfGk/3EK2SYrhuiSK/0uh36l9DKHXh+Jk
/2HOkdeWkddYWSkVIPNsplPqYnlWSqwZ10Qf+8aS3EzGMo8u1qSbcH4V+U9b1rri
2ax2TfdGC0SFtVZagpVZUXDM5kHWwg+g7I6Uym41KWCDBOxP2Aw6PIfU6Dg3xBZz
paiJbhxZNmfm7tI8O5ea5zTnO0HBYNzs3ncBtRKJLPueCgwu8XbLRDV6Kg8s5kJu
mjqSYCuScfVVaClWlb9dby6lyjjMBOT+nGZ/SJY+UgC9iAC9xOYNUbulLLMaykme
q/wyAa1OkzoKHla3SSuafE7n82i1ruxgL+j4hxQJOJFVrCeAPlIebmRevjWZtea/
tbK5abZvR2hWSQECTGbIN9tTPKKKzNbgNe8/e/TQSoynfen6qOHdBOUVVcZDuI/5
FOlH79STGwCYjhcquOV7km4L5JhOveEWDH2NVdhN4MlYkFUF3wPYPAjwcufKlhRc
Jy9LzsDD3FqcbTccptfHBPKu+CUcdAk+Yt/nHyRdVudTamFTw0jgXnPHaQoyTgh4
EdGSc20402vj2mnAtVImosFI9e/X+A805IX9+pDL73i21TqLHNxNpTPNuq+rRlao
rFz3+jEkSMZaGoCvBlC3l54AyXNzs97mo6wr26YLo3lR+RQaDvVVVFIOiZipM+HE
TrVr4YmxfBue92PT03GnPZdimvZ4RbEhbc/8KG81r9NedGW6aEPfaZ4Pnk9Etlpy
6Kq2I+EjeqfyNqOksva4Pv/zLjd6A455l6yrdlJnLWJ0MxNmpE99cb5ZaUg3Tz3E
dEC9QR1tJQfh53Jj8KiUV7YWBMTEmddH0O5uTkYcsBe6+GQBBQBMo+HpBR6EHsQp
lhdpcJ01IoEU6GSvoZ1RjYiwpktdCHPgd2iGSX5kYkWDBs8P/SWfzQ9xfGXd8z68
Q5/rj/pk0OFsyG49Uszff9rd29kxg7W/Xhws9enbXXC5U3Kdv6U9EH7+0dtxuKrK
CZ6gC+UnCabjS/yyuXhqKd5T1ZwXemfhknT9JdU1b+L3bAHZRH4xbpvf06iAhaHS
KrcL+SBHt5VazkU+72g8JH4eG6nmIatl7y8gfkMVuGB5mvoPSuUKcvDDiQYdbs9w
5+b6JkXAtR7OlpsBq+qp1moopbd8GQI6t0OtLJyBGTw/7SQuOEfv44yeFC6r30TU
26MVUOCeZOwO0u1xzd9OvqEO40dDMOA0MdZ3G41zd0sf1vjv51w+I9Mt36R7oZTM
3Kb6qwx9vGbosY3qwfClF2e2p/geM5MPJmbupqkq/yaVh0eUlMH2x+8Q3ox/VQq3
sx2F54nl5NuGMVXkCv9Xery/jgFw/WHf0vlVsufGZTrLCHrQVTqRzdVfkLoVvKfy
EPZVNL7XfGm+zsCrmHZggGTGuMEM5E1p3qtpAYu1DSh4wGJ3FtkDcmBKcXBAJbs2
FJAX/Ji62JYCpd/J6Iz8FzzK9w6O0bU1l2XCJDjzOTVq1BYrT7o3R9HqTArceQ9p
Bo82HiI7YRqfArlYNe1v+U1yJgszHWE3BDeiHbRQQsWeD2xXTC/wF6uqvGinwU8+
EKhGFDAlLumuzR8+XNO8NJzEakT+YhZ8TBEbA3NXZH3f4UbuTgeEHZI6z06T/8FU
n/kabp+82tNCSJIoOq/SH+B8mxN7g/00glU0ofv1dxC6lHvIilFZNCDc/gXMCmZV
JlcdcNFGqe+Yhb07ruMayr5MpscE+v4qfRToMzbnbQbzXePDMIGDTpiDpBFAUZBf
6mRRE+R4/cQHzHUDmHmcRtMYF8nqdV+AWWKq9EA4JWEX9GIMnNvJNzlM9YRSlMKS
+L25XG4gAy0abF4AwNl2erbuiFTTrdUOz7jHwGaOPxhSi4zQqw73LFFsih/d2qqo
WAlFykbcz7xx/Do/09q7mo1r/lLt51DZyz3kYU3gh7T6NuWPpOWujDKsCaeI7vwV
1yL8gRtPM7BDnTWBD85OaVKl531RYUWHbH/DWQnWBILQSfHAOVtsGnp09Jrll7IU
mB2bI8KoIAGccbEXSLdNL/6nC5KUsUCBKOTX9yJuVXcsILuVuW/NnENtv2USdMWX
JnzCa0hdVQBazFQ57Y13beQ/4O7JgCoBboXRTRGkap/KmFcT+e85N5cAxr1f8dWk
Wd9ZdJJ1SYOwihYARiDmWQP6dHcFaPyiSoVJwGAEZlA1qNn47sPHUWEHkdz2J2cq
aOMGRrsR44f1HaRnz+nVZflDLBvg+R5UzhNEXue6k8q/Qd1YgBBU6Z8J92iVFsmN
j377nb9LjYS67hgxw5XfQ0f8T/WzLv/+dS3ZM4hC8GmvJ0cKt+oP/zzOzAvfFmIp
JVcIQuFcgNNEBfS4KtdkHT4VUoVWkeq1KY9YYNGbYLyZLFF6apHaibfo8qWi4yae
Kn5zqdfnh3TMc4/vUzsjN4XCHwFlh80zDhJ3HJAdusTQqMZc7CGvdwcD+YlkByYn
h1aMp7b50OyU+0xggaNxYbgstMydxVz8gEOkFJt8jM3L5CROqjgXTWV8QSWh3ZsO
bB5lpfFtixvwor6CGgHCs0/fvRamfOe6WcXdBg8+Uq6q5D6C3lYjYQaqGyyvKnR0
9fpc8uU9cUqMe5/toAvwfra9sv4oA5s3VPG1p/mkB5GMpVvhfC7Z0DHHfrRYKWmb
y3AItvqoIwUJ6ec6vyurp9O42lT/WIuJkMi8FC+cUq2xuvCKc/+y437ybBDhpiZN
xh3t7uwFml7Zzq9tQDk5A5GdkgNajTE/jcvv/Nt389KqM1WMIMljRtQFRtO1bYCS
jQJUJIF0a3odN6Cw9lV1hSc1229A0psMgEhbgsaww/wqOWNGoCp4+ZRqrZ5Ds2f7
a8KpSg9Nv94kFFaLbSns+WhRDWtetsYfjefs2Stfo4h1dyqjuXEl5au9k+LjDQAv
jxoZaqT+4rrnmriLBskvgU5rndy27jZwQ6yUaYIXKJgTfPITgDsF1s5HY1X1R4G9
vP7fpmkqdgWk2pAQS+vr7DXMplRWyYUdhW6B04XBz05mZAqaBtsZBjlkZWoBOI6d
kBso7k5qy4+o0cTZq+vOlzbCcS1MLGWWxwplEziBArSgK+1Hw77UHETTei7v9G11
amuQfPkR9qZ+opUR+u9kHkX3FKAnSEJjEETkRSnqtD5ilpF6jFwF4f911TT/07+g
Vu8b8wvzEpgFyIpteTQTMzpvnyhslkHVIhJkODctc3gMsX/Nb4McGGMK/s9t0CCi
1rNg0jEALbtyBUcEWMkvnTUyBc5vxREEvOLtzhpdWkmadX7OgDLcTH/GhkwYH0ZP
c8Ge3+RvK5YIm8dlzomAca+6apM/GSfX75WwL2gwMyJaWHC85/JfbJHXBsFWzQd0
SVx2uPpwCjHY91US/2Qr5JRMMpGKI2BOps7fkMsdaoEJSUQNs2vTvqojGsDLV+Z1
IvYsZLLizqC8sHnlFJS24bDI3sbcZQKImlcN/oTuu5m77I4uzpvbVH2t9+a6Y/Dx
bG2nogNMfYauv+lhUqv/LUhH/ksKTtNXy5uqnRMV/8SnzxgzTmC+qvgDrDXzs/zg
311iCc0fmZX0aOass5vU09e6Jp/nsIlz1LwmlkGvp+oKedcF9hybXigkCYbu43uQ
8wM1TO34q3fV4/Ai3UZBFZb2ar9JzBobgeqzyaNKkZzAbKeMf5kjpa7A4AyUqUe4
wiNtUytav+IO+afo3XSFYNbKdmm135D2qTWvQI+mgIMI7HYtgGvMviMmnUnQm25V
LInUpfNPXBu584E4oUhJhF3ac7kyFRjwcINdtIjPIWPiXHzhsLKxMFNwXo2NEXfv
besEDyVC0NarCIk9ULi5bxN9MGfk9yTcmADXK92h1BJ7usvAGNH9cUREqWR5alKA
ZC8zoiQs8IaPdsZtj/QYTV8YspnuS4BVHIWBDWLY/lwm/4JFhkgs8aVC2HIba7Ug
m0E/WCmYhOWbMdAI4WFqwcwNFOnBrAzGB9wxkNCsV9mvzTJsLbvMsMQJIfyBKjJq
Cek1XjUkcj8zaJU64ANUz07fmiKEUTIcellME6HhM7qrVchbvSFv45epER3Y9rD6
XXfZknbGbpEbpteAGAyc7JSskMBGgxCTMqau3nkD4YAoLobjyUiEH9zQH9b2a2L+
Rks3RXMuykxKzpMNiJFT4wQBpikwjHIdrkvS7jIVDtK2i67eU5jScgU6CF94vkFo
AGWBL+VFr0SzdukiuX1gwuybGa+DY/W7I/YKZOn210sXS0OTII9DghqDqvRW5bBd
Zo2FBSg75R0nirHktI4gkWt/l4Sm2M4TrGd1XUWBSUo5yBULqhp8BBbxRzPcrqDe
TqS60l6AbYOiOIrRyoIpYltwMy5k36xoEwcfUJRyCLZWXVJ907YSTGtoLqPrpYBH
dacurfc+0jW0i1fpMqzHB8hIlbTAb9XvQJH53PkEtO+Mi6rK3z2bJ1QwFfTOUckZ
QDfGCzyLFvp8sN/uJDlfAlaGjb6PnTE8qdlGh6P96wOjuCIzsnZP+HfX/kDc+wyt
7SQU6k6s46g5NGNPvZeHGs8Wci8dFhzB2KkMxW5Zn2RNaCfGGG+ZAjl6/ePQLtAI
VLDJzC+WePv/3aY7/QTN5q5+/aLj86TN9pyJoRcMFYIEDTHFbF1UvrGdB1j6uYDx
v58+3ZnyxFIQHePipPqC8XqXWq9Jr6Mmra83YLwtact6i1W5VnUDHRK8RcFYxggT
waKiNu0T7TDA43qtJPBiYClCikzlY8upcE9fT2qb2L1moWAZwjK18el/Vx3iezAX
Snhl+1yQ5gMmKOB5LKhmRPPaYiIHgA3dawvnUvq0O7Tioj9eUTD8Rm0TMXhUsWGG
Kqr3z9sTZ9v6H6VpZYfwSDnRZ8rtjZrIVa3/rWhTGf/W3falVIOq9+N2CIJCHj3o
eJee15T4dPr4m3u/LFP//wYZ925dX5Yn2Kh5y00RGBCcvueA2Mpwb4thygjXr2rU
6iK0T5MdrskgGeV+Z8jKfEys7kRyqZG+UOuHgauTN4fJp3BWp+gjPmSd68g9MrOW
cQzbZDPCOP/XrVU7bPZOgHuIRBSXBFmQxXPvRe50Vah9VRPsISs1OFDvz3AB8QMW
PnzFNVjgxi+GBEd97VEV/id+GmGEFHPW8bu32+56BMRTCosHzb3DkHdviN7yUFmV
9D5191DgVDXIhVqrWgHk6jHjv6HgZ4BVpCQzM7a5IgcTk/hrPxMXxAbv/IWCGAzY
3Zr7WBQkdCzayuxmawpPpSpQHSmob10HxgPyiIJVLxuG6vleqh7VMJw41snU3ZWx
SjIg54+HWv3lAk1vswNjxatT0K3uOT4AxiZGXuJIdaAZX9IaOChUxTBrZ/7TSI1c
OOS47LQtSrk9/vlTTheWDC3L5IVoIsCDjB4GV1F4SyRDty77l0Hvl3UBKg+GwFKW
FmlK8ynBiGvthsTud912OxnDyUm1MYmTDy6osy4XB7WrQT0p3es29X8SBTCylGhp
QDJtCg6xtURnr5Nf8nOSUc61amzLGbZCnJRSlmgybwazQ+/TmA7k/0W8SJfZlCGa
YtEtIOnAwy/u5hKb+DCdUoFjR2cmNZanllVBQcPQBGMkSRZAKVG5SYPjCyMmYIJ5
NufXiNj/EnCBTxQH61ApQmFo9gLmE37Jv4wIap1Qe0P7vBXRY+iE5ffmyWFIRb/H
MSUoxrFp7lI+qwpdHFJ5by6No9TtuVB02iP1O1KA2RTWVd9Pu/zt5MRPc1XVrMsy
D+jNWAE6yb8m5ujPksECUPvMHN1WZdIXgR1rboRn6xvhcHQQTEREdEFolN9leVzr
vEOceUHFvde6Di5L2lOQx5S7k4mnC0Ykd50G0R02eeZ6WaoInxIg7U5eZ5/FH2M6
3BKzp515Vg6UXhSRIcZ+5cnytQWu8uzPM9SZz0QDr+cGoFhnNXqOlJjfXFW2EtNT
DIvfKI5l/PbiH96JvbokdoTxKcsEfp9nezjZ7O0za4zFlAocVRwFNhONLA8LoCVU
RpdWAU2vJZd8VabM5EFD8LKl11lj6yIszZSzCKyxnEqA49XVnHXfoxrEJMiiACl9
LjgAeWkgZsKKboxSjWXU01EnkDPnBUUpap1TdKQmneMts1pYJcfaec4vQ7oG3p10
SAbw5dj5oWzh3x3C1XZ9Ii7GglkU/GMutKJoa5Un2F40J2aktoQKQMJV33fe0bQh
EdXRsIqu2K7YXCAXzg2LyfzGss1dhK9CwJvldNxluWbsd+tTHC8iV8n78QCtqPDC
4fv6UVus8OhAow4UGkDSrp6lk7jy6UErmZ67USAuKqM9HybsLbA1c0tnpRALUZMs
1lNfLdontw1znFKePjm13rBSneCQdKABZD1inVkzjZXntAMhq9SsasRJf3MyEXmN
pxTWhj6DqWQ9tJ03ZZtMOPnVO90Yz4PB8eyUQr293ALvDFOojNTeTpkQ0i5RRpcY
4X3txVvRZzdcIXgGszZcBCUukyXNmHBwE1xSlr4yQOvz7Rn3lzJrhWb3BR/9Jc+I
Fpk8mjP1R8k+AptvRi85NkdPVH0NXWJZSy4Cc7GUsU31je4paOEsPv2pDOSHEcPL
1+up/Jlsl9m6cwWmnk0wjoFViqvrW5USXbTuIKUz1P6v9YwCSi2Lxb9KdvEeBPEB
KeBAAaZINhR/j5ZPEn/EeO+bk8rorZh8Kg6F9gX+Mgrn8wrAoDUfN8eO6+KI1vx1
FJX86kw5SYi0IPfm69RsC2/3LE1sqNbk1FTUA46ZX7APAZHc0dxFoROwsk5Qc71L
Scw7RAO1xwEhM8UEegUHZPn/GDX+ntXGFcrh+wqNSedKxL50bn7QJvuHtPz9YO3q
Y7+TDbIgYCLp61z5F5XcNPWv5vFRkQbbzCb0OXpx4b0/sF7+THTiQUEFtuCYV8Am
z1JHK7jm1+98EuUqHjP4Y3vfdsOlMXogsx+LMNn8XfwyCW360x9ewPl+cK6dYtcg
XXhg6TzdpW0hsHSI3LwOM16OoQoxn7O5ljhzlfIbgcPCUxEY30UsdINvTEEp1DoQ
iWV6aZ5Wl1WyfOGze0rLok7cE620Ft3XpU1MXH/OqqeqJ+shYhmlY4h7hmwey8bY
f+4rz9uaM7yk+3QTzTZN6q2oQlYO+ATWMTeeR/vF1tB+slo6C2O+OACEW0Wa6EkS
IkV3RvdJQVXv7ejnd0xB+3vxDi94U5IDASvX7nNa1s37KYCcC2PxjMDQZqer1z6q
lHegYuSy+7kuVOgFTFbteUOAKm1C7HD+fx1/KXTyv+REaPLwNkLkmh3xENFfGZ6/
IcqTF1ni7zP21q8CdeerDQVprWYYi65fGqGj7NzqN3AZGtVKmIJfcSEfKwLxr/0c
f142ScfxFBylnbBIxMAAFXZGnXm+I/pbsH2yXKhgSzdpPO5wk7qP9R/w9lXsyedZ
WdrIUvXZZFaE5oCgBbzd+fQxwAr4142YNaQ8nvWhjn+VhCgFDdS/LLPA/v8b0cMr
UbBmIH/zRSLn1gjaRiEFgUGoRGh4OS+ZjRsFRj31kh+9xVtoNyUJLcZEdNMYlSKQ
CDUcxgBzLVKrq9UE1FEI7r1FsedqBfqo37fJZY7cl7o/PsBxP0CXsfGodBGFGuII
vccny3dUQC/RrST36zfY6Bh5d1/K1ubV1eHQilzf4X3fWdgVL0EEIG8cdtGcqpzG
Ffp9QqInAxMp/HJjShYTYVYloqx7kh/zSejeAGgCfbgBU1RUXn8s/6oyq6gYNXfq
gJD+gSTl6Z/Q2aWoEtlIIFjutqF5/NOQqcjGD6T05yiTSAj4Z8cRQEBkh6TpqDW5
qBEGQluPDKDF5S1nm8UEbaB+8ty7lzIY23BMpFoPQZ8MOJXLEjw8PNfVG+JYvaD0
jOc/0O1BFeo+8ViQpPq9pGj/jQCaL17w3Nv/koBw9Isw28EEfjSfnNfx3DH4VwoD
xxkmFi6ekClrHUEr9WyFiE1Ir1HlyJopQtQ16TkOmfdkkRndmspa/Ai/OwCN9jK0
KpOnjy1XxeKWaCNptyf/JXFlYknDEnNgXqKHjBWqXttW6C6nd0LVmmsqs6WzLpPJ
hrTzb0lDUnV8GwbEN7sUS478Ty4G6UEgT2dEHQbaY8RmWjJICSQkieQrkWCQ7M5F
TGiNx2mQMLweJYd3q6LrfcNK3r96tL9p7jFVh1YHzKiik/qzHDUxOzG/JQ0R2J0+
GLLImULjIhi4CJxCHqgbFeCoMqv1YBCPsK79W3ZhhhdNyf7Rjrhs2fHBtBmbSuSS
5pULJu/43F4zE4ATJwZ1LxAmsRAYnh/iaWW+9WsqGGLrFauZoUNsmM3vIx8gkQ/A
Fh5/cUTSKi3150f34CaFqZaFVIeLxgHSUCl8Tu8JxTa9AS4tRIox0CKLrdyjVMHZ
egB+a0SR0ppBJkyd7I2JqofGFW65qyyPe43nzpnfkRSGjAJVvQu0gKDXdnIKXPUL
BcvDgDCtknpil1VGbmpJBo1QEgOGHG++rRzIoVZEY1erI4IQbYodj5fo5qKMXedL
Oe5U7M2lSm6oD0N0Rp3Ejua+oz/rAjIU3oXhfbFjIbViDJ9SpnGHymQqy06iB2hl
kgYqMNp8kcF1bQK0iKoStgqp8LHJLgMEEIpvZvy8vRgaeHOZGVLYYeBTTmkty7ib
omJvB/U0LfJAnc9+LPiHdGfg/HojC1wtGm3T+FvifuV9J+nTZKkBy8zU9+k8WELO
R8YGLc2DeCmVYLx57WpLWTsi5ZjdUm6R5paL4AvEUyOHos/5MFEbM5JWOwOCkfKV
eRDIXOTEewPSd7ZO1R311G3+7jvTBbfmISPEmEAKaK+0sITBZLkQRxk3OX0CwTyu
N5zKwmULRfnkxDWvrQXqm53KHYDtU5Z0FXFJ9WXeDil7R0kKNZCaznALZ113bJN8
G5DS19kwlccmBt2kWHpq9LfFslc7AYQN+9nMlS9ATyZ77ZnQTCxpLQxWSa2br78k
7WRqTbqi/0eFajY1duCbS6GCnFRMN6zrq8jNBS3hiN7OK5b6ZARrXqYqHFvo1Uch
NAJ2Dq0NBhYjfG4/3Ymv3VqClk4kT855KmIdEIoVh4GlYUN+0OequJzRkp6JoHKw
SjziS/R5xv/0LZuEG9l33OFRfxjq5G5seUA2uxkRWjc8xpMfUS0wEzIMPwurR3kd
sCO/Nl5Zh68J0k9gxNqPf73E+QqN7ZA3zP0I8+UX5fIE0l3cohLt187vTmY0HBoh
DO7FP3LxmC+gxfHgTSMJqVFcAPiITG5V+dwFV4lNf0yv5ydxJxNtOZLWHP+My1/t
ZZ5uUc0qE13fDmLnN8x2pf+CBYtD+oF8y5clsvLKtvyED0d/9Bo5kd4F0CMvmloY
RrAW9XeTKSYqtjLkCMYo+A1QWhMVahyh7BeOYy/DtO7cUo70s1WpgyRu5kHw+9cV
0GiIYHpjKZ6DoCvdyjSRdpSh6YxKQbizq2t8l3XpvijNhbCOxzdqzqGyno7WhzWc
lkXwZijXayOCRsZHDpdgzK8pZJo4NXX6G6fAjwQVS3sQTEtw43JJj6fooUBNN9rJ
RFZe1NoWIvjOxqAEJbk+ULqikF6QcWv3SkIV6Jy4UJGz3x3Cv+U48CijPf4bmf/c
m7JETGUOT4d2n2KZmHVeBojNNJF4y5TDbbN1SCeToUmrZcUSkBN8SiBBe7kjQjb6
3H5bI29Dpv/KRfYYauNFvTImVqUMub0aqjVXMUhCrF+adgzrxQcL4roZ1bV3rc9r
E1qnKMBnaxoiDIBEz/0Rix3XIx3niS4a8HWFGD7cRpgmlPNjKjW1J9IzIqna0jpU
8jBZXKAlYDq9ruiWeY6lTZVYB715Wdoa2TR2NwsIEznYyNUf1id/Fl3lChscvy9I
0y4yQ8UmJd0c5IIyQhKL0rSePX9WUJypcxXh3tBlTpPNPJvoY4vS7tHzIDnjXowR
IHe6VB0JV+kqi54xtozDTCg9CGFQ/I1DgVXGA+NO+9z7e2cM6JX/OCVYXRJEO9Vr
G9BlsYbd1D7maUy/73o4BT1Wpc22buimCUiBHXGAdE58ZU2cuuzIvuj4e9QEk0pK
derZ4e7zSf2hgIPOSydCIHSOhw+WOzeHF79QEq71oG5g+dXibMKXE/A2PCLEpGAT
UkS8bKuWrxSzF3EOhAId4RXFuJ9PBSxwGKdAo1aEmxM65mmFPNDcOVlVNMUkmrIQ
Sa81mPH/IFVFdZZc2Zwd5YOwpRbCVhZJvBkCXJntscCemYMa0bvsMRblwlMQzkXJ
SyA5cBQh66GzUbqIQJNX5V9apDJsdlMlJabtiR1wtB0nW/F5PclDGIEpLcfVTLA7
SoGmFhX+V5aUXErR2kYkUkSpi+L2dzZGv7GQNzmTQpL2imqzY+9mvE0WetpLIbg6
N0pZ2luy5N/0UmDPQI/0CV23jOckq8Y8Y8dF3FGz6TBLGEYp+Bzw19eF1QDoqROX
fY4zBR+pvaXH5fPkYJqARzRXUL13XpdEIV5ldvG9vl0tJmCOkqI/B/plKtZxbV5l
xvw/TR6kP0OLA7MJUtFlxuQBQUOJpBhs4mbNpKgiqEsknnfucB3xP6zxwq3/bGkR
9feq+Tb/+2FiwTBScdTrlfkXgAN6wKgLN1oOK8eJ0NYA7GuK0JCkvmMjChVcfUWn
/njxrgt2f0ueFTctWN+ZP+/1s4rWASNOj4yWNdtCfAxYPThtugmTuqVPyAl3F1Wh
jCiweDAqxnhQfvNwO51Zx+w60dO9FiGrEt/VLTQbaporM/vfHM59o3UDRXCYuBBA
+Me0IxakahijNqgluTt/W7PKTRNxwCM/ckjvFNRiOvzWBFRUXP46NpPEJi1dnNeY
YPwElsZoIORv3XKg7d2hZWaQspSyh7JMumbIt3Is9HPOydpV6V3LILcrQjV66bGR
eA4/khpKi4lqp2Z4dcsYGOW67ZbyUIxiWjhODnlxei31k8d3Gmji1ce0U67a2ETQ
m/flQucRZk9WUzQZy+j7SwV2NkioLEiAFwFq5cSvwWNeKVOJ3iJJhIl7m2s0pg/T
0SlKT0yFmUsGjVHKqRbu9/pjSpIDJrqVbCiWu6p/094GTe1a70Srpy34uY1vTvcr
7UraOENTn27VgFv0ZirtbefdteFAQPuhZdtQUtFHh/maK56CsafPIWTSje8DUnRB
q6x8LZd7JrGEjy7oQQ5KqDNJ9jLgBuHN5Ggv6stz8ykgwohGxtpgKKpn9NFCjxuU
OqAq7n+89JEGwGOWOeMjH2IYlz1UwHX9LVh9CvrnTYYZoioymcTe4dpcrSBa4YlA
MqdZuVFMhwlUGXb7P60FXSXHj8Pnmhl+es5yiRd2ZpClwtlWxOSqhI/B1zoqTacL
YaYKvg07jRshPpFon9jH1OMgPAr/S80q/mDYQrXa0L1D1pQ9DZQVJ86mwF6Oo6F+
2W47Lvh64LP/CqKwpKzPgJoUmKZVyvuSqMopQJqgjVT0Z66LgZhARPkqyAcuJUeW
gT+oA6E2pAcyo5wGhUbM/XBaOYcGp9iTBbrA2emZqyZpb6GfzX3ntkHotxW5Z36m
784oOhbUkPRi5WNFI41iX2vaB4MwXo9rSs0hgP45mW7jjR3iwoi/W+pAizbB0EPi
4PShxuYjIktErXhbZJ1gzHqmArUuK890DKaq7Itn5Wqa6J+2OIkcanUhhH7edxUN
0XbDX/PwIw4hf3pf/YANZJ7OgLMhUpIUsNifCnKCp9XGbDfa6sex4IQcVsG5xT7Z
J0l5486fSqX17rF+oqRh8wn1WhMcjZLdydGJ6t0zckH00EY6jcc89UdHK5U5fUBc
O61m7Zo9+8HEGF1lK+c5ASS4/dk/QxA+cUq+htFocKBXTeiD4IDmN0kXqAcFonNJ
AAb3Q+bN5VX5ZiUvuxudcUCL07x3SYzP4d7l9fIHfrb5bzwuCUt87QhZiXbqKSmr
+D7tBryFGk/15O29Mb4L2F1u+EyPs1WyRLNf3eR+SOTsz3jovsk9nNBadxulvKkI
DzI1asZsJ+EXvbcJIu1q3njyIpU62GX4LkrdbShnLbeUFBt9Vv2r/l7XuOd1Zdra
4tzEdguMAjqa5QpqqQtLWNyz4pI4bQjLp+jZTRyeOKyBTzw+YPT8swv1UOVOZ1g7
wXn/KiHfia66Kb0UCk1bYBdC0OxGuuM54bhy5nWmsdOfWPm0vHpuIhYYOU0AZQk3
tPdih8+qPZJbO4t365B4swKL/wqt7yvJVD09aHCWPeGiyrev8x/3aYmt7YXLR8yu
7Tqaq2AfAW72zrxzwJjF38jR957HtuUrk33oD41/ahtTMfZ1jINxq9G7Fs2xC8i3
/isrd7vi1/k99tpLS8tU6jgjV9VaTee76XkbfTpIY7pbL8oKyQ88ly1NOzJkDS7p
3kL7Wu0NC1zNkYgN7MwgDTH4yUOZHoOK7FsHi625wRRck1mZ27gxAEmWvHMW0N9M
DS0KURw4AhDluLluIFDU8ZP1nt9gxaOz7dVkrh6aNgCEGcZS6AzWJA2YtrL5Dq2z
xWXnbmCIoFGGQbN/yRXqRq+IdBaQHRDvuZxBW9j9LZqxdmDU2lSp2MdFoVfTVKe1
BTvGUKlqcTObHs7t25GPtymwqFWqudPYyw/Ly2p9KPJpLIxbnTe5VRSwLdF9AkMB
ug7UQHz1duYm5d1Shuo32YT4nyNUghvia7JCtSDljh45CWC0IofbBkwiOdiIXUcc
eXVy8o8PD7aOU3tAIzKMDXIXax+o4hz1t2szMYxD8V5Ve7ELEjo0QKjJxv2fOGaP
xEFhU+C9rcjJv2MJzvfZwl9ymsPq252WqcLTZdRQEj/IKnU8GE0Bxhxwh+yYED+y
zFJvmZHFF0ewDlf7+Og24mquA2AwMgt9VDe0f5nNj7uNQunmBeECX2nXRxcLKhls
XJaOIT8ayM8HgGRjEgB1D0O7qjG74uva/2YxAFd+NbueYg6HJ1aSM1awlyk2RdwG
k3XKs5YtCPgL/U9yQ4dQEcLyvPcFzW8Cxb7r7sPK5X4XeLzgxAQATYyXeA8ba+eo
CpB1Fk3mIZnbZkBpLlkfRTZ2x+uyMNm0RIxSG+Hwj7WewriWiymEJvMDAVisFJe2
3zpztqmJ0olQLFw4mt6zM9eBu7oJlrI5oLTPonwPhsccaVZnecJbjIT9PbJemID3
kYCIXLlOrmdKXW/fieyzGVjFGTnpYRJiye4R0kDRc8dP7TchcmTLOkZ1x8asCY5h
+vJx9TbDyIKoz9gZUo+8rcY8GhWalHFqmxsJx74hEn9yXGYGSucjojdohAlWG9aU
9sAPMbjqqD89JkvxyHT7UgbdB/dWTvEz/sLRqgTRO+khRK6NxBfmxXIDEbqSbRFP
BzlT2O8qvIO8/FBCYEldv8hg6ys9b/FOlhaA3/UQ2QOu66NgVajtblNKrknQmNQT
7BAam14PTQR2ahT+wE0KlijevpklFoAwFJ75Oeh3m++4eaupby2XjsJEz8jGyavg
UTxSuE/G9w8dyOS8C25Sw5hn0PjGacFzfIRJzECAelLL192JhIelhEEJWy2k1hf9
ucNhGLjT98RXb7jQJ/B837gZ1iIFK3zV38cC4I+r80tXVUVY1W84zhh+z2gzYh4c
PU25tG0U0Kipx85pql0Zfr3F5mdTOqFkYVrXudx/YkTn2SglDkqJHDh7RmvYSoLK
29+1Ic8N3E32srMgXFJQxxjjuHV02TL8bFgpokyjkLdsXzk9C9JRuV+nUquerBsi
xKJuqbljKqt9o5JQjhBuWLbEx5lpLlfFFfrsGTziOYuiX7oq+dq683sK9xmMIqP5
q3aVZ0t3YIBNj7hH5JCnSEpERt5BYsh+LqnrkUNYNEgxlHV84e9FkaFELRdwOxP6
J4hFXldeUKuNLm21yrzhT7JMW6di8v9F+Cllb07kC8DmUfoA0DKszTb9LSXrLDOT
Giq0bX9kBNm9QxT39r0PrXkVBsSKM7t6WlqNJe5zv4twwBqF/duu6ykRIRewqZmA
lSc7NOa6+0GK5FQHZI+42owx6gEYVF5L4oZ9yS7bDQEAl12A8YIoJQ9NKWk1Iqx3
/pS7G4Y68xfannbGlXjWtxPa0QxzPcCaCWUD/08ln4h1jxmRMR5TmPSb0gaJr8vz
CkYzPIh6RYE15Bwnsruv8KqddPQu+OMOGUNE1vra2opl+WxDViJ1xe7nXyCMPaez
BZCSFovP/JxVeG3lZQPwg5spyNpXtQZlw2H5svZleRM8B2NNBy0eI1yLk3d4P2Ga
pYU8DrA6AI65NGaOd4WnRHTOC4fcfy22j/82jHcc/CTt8KyFrqpTSNNKWZmtfwaZ
ziLWWnsU0w+YZfvXGoouVoeUCKTk9VqiT06uzKAKIVpdU79z9QOMzsfwZqlesOB+
07Nkrex7CQQv4s7pbi6nL0xfXOztzqBF9SRw/7MnSLdsTkPcR5ez5OCdU9rCiYJT
EgiBkKmyT1jXZCtMYThufFSVFrExfDl7JeoyEzJbB2bjEhYCEMWfLGNxOstnBFQN
LCVkMlzuYs/PN2ONAjkDOw+i8CKqwn338fB2Yl99XL5rwSPRJK1d69jvwSZVDyXY
OcHCrZQt9xbmj6BlnKSZ3UqnLYGOlkLym73rzXaGULtkvEjBwE/07ThKbjeM+FO+
F8pgYvYUpxt6SrCP6WZZJLep5xGdVGQa6XDpFEJC8WsoDGDcxDnjgLPgTYAMe8xD
dcje4pJ9JXUN6dPuaBgblGUaM8MmlBsEir4jfP6ppGorg/8pbxhnD4wl93LV1ldR
3vXPiIBtHEqGonxxVY73efN2ALhUQ2jWCbosTvDwc3MK4bBSfsiV7q/3ASafCsME
RaXwcgoaa4Tau6ZhZzz5nciWZarP3+VvRVtRcPjcm51qr6Gllov7UX8ELkQRh1Bi
qx4c7bXpinlXnA2tATd8yygGBio/Ojvddk0KZBObfIrB7jg4O899hssD8gl269d4
CL5goE7PUFv/w4pw55OO60fLSlS1s+03QEoKja4adNZFhqqH5oZAiq+JHK8whnAJ
dtFwpZdUYrlEjm9DpkULF/53GYyiQGC8y5aLZ3z2p18jAMz7xvS2PWPqdJEQljts
mxCGFI1CENQoUqgTttK60K2Jl2C3eKYt1+m4zSwliCnrisAztgy9PzPIFlHxdpWe
JtrvN2PRvy5C7cl0SQgO7sY8hwUIyoJwQODIsalvhqlD/jUsUSmepuC5b8N1r/Jw
YSmgS5A7wScYViyVGoYvBjC7D4ZKTgnedwC1K3ROK1Gg0znYdUytJjimaRdBwbHQ
DMq2M9mYAal2XjdoL7fwMRejM34mIDIKcvbJdnyIS02/BSZ/NW83IoX6qNVVhZ9K
3MANpXxPJPuZh76tf5B6IrTvLLjA4iUyKhNtjkqfVX229mRdnhTtDrrpHhvVWPu7
gFvVKUhzJeNrFpirZ5S8vKnPQ9+gJXEP0iK7ha9FHMeAz4Rkob0oAs/uW1gbhCWd
m6uBWulg/SNPQXPzW+ZwdMVe5LVJggodrPE52vJNvyjgqZFZJrIWN90O3Z1r6+Nr
pwYSZn7Z+bYA2rzlYa9Uo65EBV1Gr8TcJQa96/+uakf+YEScep5MFV4SmmvwkWUY
2IqDLbk/oyk1CkOu7sbh09jVpypH9XFrPqhA47ud1hrYQSsC0rfpshe0lGraX3X3
yRK1lQHFIHCiyPFpo5MsmQZ6QtvJvbel9ra42Ueqzvurdga9o4EHuRXzFtiyZ27J
XXNg3uecGE0qhQMwOS8LHr9QLYN+xW1mXEiA2X4S19s/fq1a6N1RorqocQOlKzNK
d5t4cCh/OltlH4HSOIGtzxM9sGhK2IzJcZyQWNqZu/u7EJ+f+Nj9W54Kg3AX+/gK
Tc+oaE3G7UKE3xxypmeXxDZXnuqvo5nQ/qrOXBX6JnSYGNoCXKHa2UB7FKFAlBpN
Gg7VnVBKTbtanvWg2BRUEZMLddU2pJGTEyEZ1O3C24wlQQLi0tlC7McoIFGJkx9W
5+Hrupa5/qr497wYz+f4G8t2ctOWDR5Y5hSNam7SHBetch5QeMeF9fOsWBJZZvz+
KXNBIrpM9FaFRZWZcVplX4CJqMNpnNZZ2if9IGpBQvtdZua4/SazqJhkQ8AZ3An4
Jo5T/2P/IcbU5B7JZ4Hfdz2dCa7s2Idn2pkRCeu7MgDhUba+s/VwlJq8UrxE40Sv
SUKAgGPuC5oE1rPEmGKgGRF/2eCOMN96CgthNuiGxZ3ilWc+mFOaFUTSIhxc/51p
6fJuFhanaDHCqNYphTPiijVaEX3sZwyAiwpGzkFZyZ/BUrNIQVdt4TvBpJu9DKdx
tdKq6amBzNBqJeE7ACDouv8qjSA2THjlNTioSycUFBYu/lKPAW343Ccy2qi4/oZy
M/qprIa9YSnbrbnnO7Rm9omLl2gPDrjKCtbWWrE3HWzXFgo8klsKXyN147aBVmaO
Lpe3c419zfzATjq3A3dgxf8HWLm4AGc1CKmLSWnnO27n/lCNS+/lz0C8HySDBv+o
39t0fCM6AMSaF9+jErjtOWu6tPCtjYYLoBr+a1EGZjv7z0gDnuiwJ7XvVJhZMbX+
rwb6YMDfjFCyN/2TmKRQAemgwU0EWvIREPoZXhVKzmeL3Ah/iePLz49ig2LN8CA9
dsTuHke/4aVpWG7X54lBmnZhEzt5heSMHr3I7Anwmg21xiQapplsUFgJXR1lwgXb
Q9We3QmwxlFpdiwZSEyos9UQU9w4RK91KzbM3jDTUHxHP1w33FLy9wiHIHF13r97
9vRXdAiX/8ALApBoNrBoSlhv6+NKgC3+lLBkgeZgdQ30D8HABJP47tYBwakXRXvF
n5qirh9BpFQD7/CYQo3ReRUagWEHcNY+QokZZps3Cidk2UlP8AvmW/ozMXSIsjjs
KJ4zrMSFp00zFfjP10Q/1XoY4Bic82I5n/yntaErM++NEFvj0CsKg89Qk2HeDFb3
p1rTi1lWNKjW41vagw0w85Lz/2O1qJPAItSgs5Axtdmj8DRWmQH7mOxku9oT8XTR
7EFktofX70wgiQvn1VndG6AsTG6qXMFYcON5jEOvRL+/K1ILeyReFjaXHBbuvdOx
vAnexvis1mcyOtMZAfaDJVAT8JmgvRt10co6WB2D3rjYWXvECS+Qt9izAxhFCAlh
3wYhJdSy3qCdpBvwjAWsIlxR5HMzyogGD6rqg3+lNTSmEXCjF/s5sMmbB38iNMda
ymki49EROK/bFVREscKfZwNNAqopx1i1kucReQwFkLW7eib1jLtkZs2yki8aHNsZ
nBlAVUYvwu9EZvHY5Pc8uLDBP1FAAHltRhbfb1JTituRYIfd3RFeqxN8+uOVMIr0
KmJfLOh12l7d7GPAPl92wPUyQcuompsjQxJ7Br4rFKc5kcenuDRoNqGxORKuLHPC
FRqBxauoO1tMfpWWcCAz7TJKpx/Nfieg8P0riASPR++ZVnhDAmtGIUpVX6XQl9t/
x5/npgn2QGbA2trcShn8UBEkrYnajdF4+cMT4ZbuTOzpzYSWz+drGrp4YdH54RtY
0fsEVZkHXIkDJXqwUiPHe+FAJQ6ReCdyzUSip8r0bJCagXHV0U/9gD1FjvEx+9y6
hqCtJ2HhnHCJTwkGnPCV3NSKQ+fOncaf7f7jgqp0ums0lhSRWZq6ybn0XmN7495P
0uU/FxA+Zg3kTl1ux4lyCRloaH4HPsWOmhTHiZ3iDfQTySwvex4XCO5O1ZYQX1vM
7vgXTEY48DG0SsPtWh1Xn/iSE3d+VvkncL19OqZQxiLIx5cFmtYqJpr52EBO/JNo
qDGxwIxI5dgJ/us6dc2BlkprLPLX+TlGqRfLkVDg3jBc9VPpqqDeCbRclb5IlVm9
Rlb8PdzodMWBosZyy4RyzQ28kYCJGDS61m9G8ytyobAOIAolPhEgDGlpciWj9GU+
KQH7eV5CDHMScPaUpUcZz48HU4JyUMRa/sNM0LPIG81tzaECI79W/vP1zfvNRLvD
gEJ/wKuCJib39OfzjefXcAC/Pyu1LmXbMx61T2Kzow991pb2MaJl6SHRZxMrFK1C
eCs1qA8IAO27ZrRu977a5NW0mrsrMHmTOWgp5KtiOkuKC2jOHOuBiSeJ0lSqMjlX
Z0+RrKVjP4F3ZyPjUQd+ho0l4+dt/r52ItUnT+NVr8YBcTwaUlYh20nVZ2T+D+AX
5AJ/qEl3RpSHqZnIpnubjyHwdpW7/1Q3s5wyLy707//w6xMCsFEKIIX9LJ76uWZI
Cr23YU3Ar4jB5FCN7XYLu5CkpjzDuLWvKtVR/Gsd6veqK642FrwnS7cdJAclhvTI
KIeMY6xqIK9JRkL4YVigZDDgeFUz+suGH4I/TNYZhcUN9DpfHIe/rFn+RlXvjGrg
Xq6t+Q7i/oUR8Xrhy7L53KafVzopYtTOyD7ZXhuhxQt/YVAgMIv9icj5a/34GQx7
24Eg+n0+S0FRV6Y62Qt6fqMFSpJ5Vz0yNnoKnX9xleXOdnENsBo4TmmexuFpKQeC
oJ0AxkR5bUJiczFsgR5AFkjJtlH52Bwdwwbg5DcenQavhMkSMcJFjp8IIMoCxmfQ
7vqH1ColTQiLVwU/USUVAbbqfJwzNPaTEAtw69tEP/6bvk90bUCuQMtwKhHTtaKE
cKVxnlby+bekCGRiVqDC0+9D+ZXG2jQRqmIcDTfAMijC0XGkhVxTkLRmUbY7ArwA
LntaqEa6+guKxKvL2qWOMrTBYSttMYWHaNB+jL+zmWbViklWObahm4rbrx89LCNT
KihIa+chJO33xcYvulM1cA4fAeMohaTUgHxdM2FJwOQcpUUC49gTcbYAlKK2sQf4
hkFNPlZj2IiCD8tC6d3Bok9+GFfJWeldcRC8x3J1HmvF8m6Y6RywJY1fSxnFgVwz
dQqpfGUiOFm0YfUizCyMurYo6rjiSGKD3kB5dmgp+vVavRysQK94BoS/uBLsuBSu
wCVtD3XJfaxpk9twYcORdzLB3jhI4EVnQ7pFmnO9eqyuLpEOMKQ/Xg9KcI5uoaxY
BODKPB7vsGumzbXBXte9PkOTRwliLol3Xv/n25h5NilXCBRO4hjT0fUNPyBYVFXl
uWzqjqWc5nRP0I1/solimBSNPUShEAJmY3pZcdHEKWJjXfMDPHJZitcHE84+oxE/
jjj5ALjKsJtEohR6M2F+ULSwCK/+9NgDDJo3JCm09DDBfP7i5Ypc0qjT6iwllnLt
7xMHbUg2nNpAvHX9hB/aVhsUqjLQfe5CToFs+JEtqCMGzeLbz9zKwnMnXGk3Mybh
k8CVoERNPY9K6tRYzQqJ1HJ9aSV0X9femKgILqY6YarJtPHZtJBxM8XVSqu3vYcp
yC7Bt/Wo96ONflijA9CW82H+1DGNdH2N6n+pvhcbk9KFzBd7fkD+bBBxrPtC71SN
JOqJw74v3/F3oDEdlH6k/6uHFU6l+UqUXfA8eQ1CFbXIcx1xIAWpWUJyD8kMbGmI
fKOrwmBxEgU4wlz1pj/jQJ7qREwE7VZyT6shoNGLsunCE9+GNj1NKlHYt4yqPlzV
JPLGnkEnjsYd7xA0QZnr3G4DFrKqNBoqbP8hDH83fNZXf1HNsEDHttGfETOIyoyZ
x8EylEHIV9Pa61PQ33INFOxVGrv8N1Q5niBKXChSYEW0ooUjY1bdyGM5iAyxj4sF
dEird362Amy5RGIMFpOQY/bWtHUifmWNRANDjlWj1oCWXWhNCtJER9CAjlp6bHvH
j7g6giAeSlmsAXNRZYRlrzeoInF8ByYUtS9Ffd3ur/gkePHBUpz6I5LXYXcgm4zh
bzlAYJoVfoubK4D3Ke1wf21+kI4WUl9A6dpZuYvzBcr/jPSt1SBen/NGkuJ8w4wR
wUl+es52DNW4OJ1MYuk2O1TClt11CINBAbdvvSqrbj80pq32p7eekX/7Rhr6kdpu
bXI2hV1n/vQ7zdzx8vCFsbG4rLHcg+mqBO2yF+PPEDG+7bH9YMUDqZoKwUGgC/e3
Ohc9OnQtkpOYWgjjDVUInMZ90rmPiv94mlDJol35fUNn5iGzc85qRNfgMlUtrXdK
+0V4k8lUVTYf91fFDeedpnUMz+4H9hmAEF7ZPSaBRHWeW7gxwuZ9B2ixP7fXfx0z
IbWGL5w7eEaK7R9v0W5Bzgc61O85ADv+YBgPVkJ5/O2f9tK8KyAQBR9Do5wBregH
rmRLesR4Vr6MSsy8jZGrVP/3b/BAMZI9vCGMhsmnm348pUkiuVN+4sm/6ZrtvrFe
iwNY5wJlWxTP1N048JshF+Fnv78oc4cp5lnU1bHQ1mRGjCeyrUn4Mapxwcb4LR8q
XwjMBgvsTtDKVM/QnvYNX4zhfOKEIzSGQ7/zqTGuy1SW8NStpOdRx1fAyhSL//aS
wTew/d2QbQYtJoao8j03DE0YcXSmnh+h3THOAmBagzZZIHpaWU+ZVZD7zvVOUisl
WHb6/SzRMBy3rQ2eflzooFjEt17/nPQmSdp+7zkeyiOSx8HIc1vmssDKyrEOPbU8
9G2xPQ0aILII6lOaYMCDGiyVCjCyq8J1VQsYxCpkauLlH5f8IsEZ8qaIXQnLBJSI
WvpC2an/GIQo5qVAoDDxLONxOXPSQkd5MNYBwWoMuUOD9fdm2XlmET0vvggBZvYU
IBvBhDFrk3oh2POL9x9EQC16bq9JVVbJzdUfSb+La1sZ5quHs0djjW692OuEtR2d
CiZNGp/+Q+iW8xueurgsZhQ9fV4WHrHE14ftf8f0Jdf7L1ToRpCenOBQUMgvdr+J
k7sasKBMoJ8EgVZRx8WRDlBHf/cGbhGelZzU66Wh+4tATIn8AYrrsu5NyScPfv6H
QNwk+jy/ZL2F1pilY+StMqO5yJhrpAjq0bc4fsCV7D2SQqm1zytrIJcRJAkkjgwO
wH3DR3TGDZnahPh6/JzvwKisjIJTfy+KvPA+WwwgKmU7azdYjIuQbtGBpzSfnMGM
EUKLL45DRFEtG23a4A+3gTjMI6Wkbg2JdZXYnYUPxbxuSSzl5vV5xmj38FLwxWC1
P4PwTcpvOmMPOGnFGA5DEjrorWMo17rKrZaIfgcPRrrOAacptrZvoEV7il0fDkIE
nxxC+xIRlbMphONsCQcVBKul/89fBSa1DhtS3Cx0l8q6lfewvLMPGHsdEyGWzQaT
n/hqVQZtSCkv3mE9ERwBRS0yYwJwWTPshuHPtqIeV7M6U8ufGb0eNJN4qS2i2VdJ
xaS+df/yX4JapWSTJJzmn4bu5IBdZdLGiU7qSVNw6POmpB1A+Q0l9LKSVxvgN7vO
iggSC9asUKXVzlXuCu+zrSkwDq+ZARs9rO3olEIlIYFVwDZolV+vbB+/jFEfC0De
EUIwBQmjAnksNhIua+Y4rleeSjDnY25Kk8w5LmaHV8x28/2va4BC3zBr5il1qWQy
LczmDUB3N9yj3Mbc40rKaOz+vAB7c/NaSJNes1nan5RYEcKLrZoLMXqLo7oYkou1
DgcjtLaoCTkfpCvvQJ11fCDK7zJixcqgzTTwn4+Foww061PWFEurZ/GLuJUZzr01
DGm32enr6s5Qm1y4I5ERgYotixz4YgldvGiZvbKdxuFXHxheYcJvSPcnvX/i0Jx0
saqL+bwGMZxbKi8M/CMJuRlPDcuxwNCU72SOO4pA4pZwbMjCY9PgBGSbp1FCLmou
fkglpGLGBeQPzcbmom8bdWpPVjbgQtY47miiKgn/4FrJ8cQ5uhqf08NRlKeXt356
lOo/5wkcTCmL63EFHoyMg4xp6hQinZwMCuWX77L4UGNYuBgM9jpfz9W8R8MeyUJQ
dgpa8XQhuEfzYTLnbnCIYRze1kLPhXj5v4JTUWb3AsT83Vv8IRuxYmii6ziqah4h
gHvKgfMr8DBTLuE5UyCLNtD0SjrkMDCIgeeiF+0Vkz4UlDGVq+4ycLIgid4+Xmem
jXCIxLx4fZ31IC11S5RpqXtr6+HZpJ0eSlIO+6r1D2IIa9CFvFes5S5dlDKTV+PN
+rElRLCfKlTWT6fj9ZvfZZ/DURgAHefv1R05IvTWzeXSdOE23933rLzmmA1nPhqP
tv1AtOQM/ipcVYafGF+4yx04QvASU/1KlbNOW2o6Lahl1zKx+a9i9JfaXkfI57Om
+uBxlMjDPoeQVPnuCOEUTKmbXNZYaUoLlXUOQufLtzHaDjQPxyNWsHiE+CfWFr68
wu7J7D3b/gpNVAH60KwtkXPSQej7ONiGn8r5Du0Ut34YgfJCnjKNMLSITZ6/UqWh
eWLDjV3+xUskI8v6pQfN/O42y5c82ZuMaM102V5LzqPzkey31aIStZocO/nVs18T
m6rOSn1JVtX9mVU0U92MPKQir2QhSYEHdRbXHABSvGaTvbuv0TX2EOxY7f1+hywd
9nPuXd4RS8sXBA0AaAKqxOcLuw6PcgGaQ+tJjhFyzogA+05qF/R/dYGp4zP62R82
nsKCgr9lGa+vwM3+/a8SdMimNllVk+XQTaEBYzb8d/0/p/ZsRCJu6eJhVSriQyf2
5ECQ9+bBdqjER6IqNbBTS78nloJytZ5YEnHpdKeQqip41Qviu2Ts9Pej2FOl+vjs
hz4KpVoCLJ89acFuS7PlgM+uEhgeYpMjGFFmxYYBCZP/mgXJff1hxEF8/ZDXsT2y
OSFzpJRpi/ukK8e6qe/Yg+YseG4xdI15dxyTNjoiicLITGHhuvZQ3fNEkKqhWcbI
v8mYmnLkteDJ4lAXQTLz9mNJYL72fZJrdqU3iezieYZn9kK0J9P5Qhewa1c7vDsh
x5NOrZRBPbu/hPT/RpuRgJMm/bh/oZqOUwW5G2rkJ57BARb7dN7m9OXI8pEFFYct
V8G8SbZSR2hCbvKkBJYkjwHZlu5w1dFmVCJbWIqioYj1r/LvWghiP9xvD6IgW2Yq
SJml9NRlvn4a7SEAXcA2NUzY6MVe6h3Hq5e3U3+HGXm0btR4Tq+m8SB/EPPA05CB
r5zZ488CKHlXmgNAe1SvSTGkDjkubCSu19vAckHMtp4v4rtBA2vhi/f6fxEpkHdW
2X7UuzOF3ZabEP+3XagEfuPoDn8XaRupRpKq5oErYCCLGO4KU67AMOxm9OPax2Mv
6vJy8FgJhUSxoHlF/C31QTYiW/Fs0yqnrW7HfepN2376ZfXnEVgWiWNEyS5/JO6L
xTFsKxwRAW9Br4ktGOXo1PwbdSBeXhqetPR6Kkmowy9M2jwmMwnl8pmcmoNn3kIY
MXb9sRkvHBhY1VfxEMy7Gky03EHLQI2Tt5ODvFY7DLqfaI0x9guvfYfkudZMEoSe
L3wgSV7g1QKS0nG/sTYbFvZnre1VxBrX00USL+Xz9q7ie5fBffcRCal2U2Aw229R
sY3RPSZUWd8rj+W/GUsVur3YS+amnziQRkUJ9Fo0Vqn63ojhitAHUHPw7tslPjAr
wPQKdZPoXb9sgnJBvqvnL3cnh03YDuTAYrlX7KDO/f822e63Iu1P4MckXSSCmw6H
t8PfM8eDOKvSvMf5u4ZyN/1VapgsIdaTEmgqw/36h3lUee0Vs0hav/U8RD0LGB//
ySC7FBddxBSwi36PTVHBfOQj4+WEhpXoUdfrEbd4Cgk0OfY7h2IWBqoHZ89NGCRH
ZN8XfjUM1PGSQ43SaVW29/WJaChlSe65ag3yyowD/0Ys87alLkQCw4NnRbqBhIHJ
3nM45UauXVYlt6o66HXPECMIVjSKM/m5Umaou/kWUYoq3YrPtD/aw5evU6nvIgFj
V5PcB4joQmSAt/StfF2k6x5LTX4nMjz7JDYT3/vqKOmAcY/qz87bIROU/5ZTGnGg
ipOm1xPTXDDpVpdQ0h750WzgL/ruXhn+DSSLtJ2Aewnf/MZsenyD0yEXWpLo9eR9
fiW9idqnnlZ6CPh+I5WrXGOfztJId/4oiioYssA/sudygOdXtjho1SWKXjw6ROr3
li1C9Zv6rwLoB/znhwo8cEaMkTa38a23rIVHpX+qRF9mwFpvxHPVLYMFqKjHjro/
YHFN8WwprBpSSl0Hov8xXUVmLvwd+F+Ntt/HrPKRgd2qIc4Mqu2gQkBNCOCdH9W2
CU3GBX7paQLkRBB3lTH1qAzRLYv+kYa5YVtQ5GyO1WUSPpuZITJtftKyRqYIDld8
6njCFEAao5mbU52PJClI5rzyLLuSrg+xrWLO0kfY5028/Oj7Lq7Oa927KDGrc6CK
XDDZ3RUT80twgnPQXyWa+NG1gPZmAFE4DYT/iEdTFwNCs8BkAtnHnMklNn1lPf0/
NOu8l/NoQhPp0L7GqX52LllPhhjkl/+FmZ5F/wDGA4wPKKP5vmwmllHm3Yn1Ooy9
DfS9LU0vsGA3l4GB3kL3Dg6qCf78NhfPDoWvq0M2XQxh8Zh47aYyuDwKx1PpA5id
0OrwKyjsvcOb4vGsfOeTHbe6Ft/ApMFgxLRQRhDUIOTgoMo9cSXXx8MXaJsRlMlp
z7JvYS46PZxvY//DRKeVmrBVAPUvxQLU60d0NS0aUyWLlsyBlIUlLY5VBnc8mTH5
bYzt6qs1nibzk3bQ4vUVCPxq+0DbRKo7Lh0cBdjDvLlsKDg2BzcGTjk/6KvjVOov
Zpm+uus0+a5B538+k9oCxApYAACI7cgNZKEu/t98BC8ux9+B3Rs6wpocfIty0HeK
7+87fD+ypD85ZV+LKYPYHJK/3SwsJeKEOQh0a9ScbHFFNfwhfOhzO7gDll1dZPm/
KbYykdbrpNXYQTat5WMp5HuVV8DeiNbKH4IAJgqNmMb/nFPdz9imyrDuNzhczDnK
UFTxrTIsXCLuIlDAiC1nBGS9GST2y5ohTLKYaq7OH4oP+OJtAfkexIyxoqaO4rHB
jqONArZCHYLKOepuEinriYwQywoNIyW7AG+ExygD1bxc/o0HngG4Aza/HK5d+mH7
v5fxzFRYFd++K/OTCnwXctucl1n7frBw+z/6RiNSP0ere7evNWX2y/5GDADJsnln
bagbXnqvteW1o/be0P56WriDIdkMc0aa9ujSPIyAYJhLSZGLi4xI2XRDeV+zRJ9T
lQF2YUKM8xpMIUwoL1DUM10G+Qw+iNqkTKPqYNzTjJLisDkjabFoh0gdBT4D1ME1
/zUP+t/QHZXQrBDoNYHt/IxhFvMjizqPyJqYpQm2QTrLgb6vYzRMsK3XMTbX/Pfx
kocovmzNgRUnSRsL0PI6lc0fzHl4sVgO7D+GAC31veHFp3Dhne6o+yAQqNrP19Ih
41S/hEAURACI6i9I6Y1NBAXf9K+apdiDHMdDhrhki+oh2j+MKuMEo0LpiLItRxXp
ogfUuxbiymGvS2YLhBjy7gGbTOICizvrqXk5lMYx+Kn3ZwS+JLd4/Jgj44iv8nYf
SURnKrHmrQk00NsjTHmGidYhlmXDjdlMGUNU92dswjyLBbkbchvS8BqPVWxd/aBm
ra2y0xEDMP5sjUfb4JZcdVGIPO6c7ZPWP7uGmxMaRRLoHzqiIWj+O3UQs7VjXb31
uJR2KgYYecEIUxXz8yVS2BN5sL3Jrm4jUr9O03rR2EZv161P+TsF7a4iOkxAc3XT
J/4lDoDiceKpT83eWhIaFZCcVQFUtbfEjfZzggKfS6AjZx7CJoNC9WgnAgEhnS9Q
J3AcOA71zh7q0+8hM605jBfYoVxxKOJOF0FO5TQP5HOPNzzzTxGxxj0y1AazrU0D
dmjCJruAi83RhV4/VXgAOY6JZ0EqeEMxKtwEfZ16KxyBohGfGESOxiEnWa7XEPaf
ns7rQDlGylG0pBvtL63qgdQTI3XKW2iejbaqoUr6rVNRFMQ0TNKrreEGhM7AvM6R
7YYYxC8B9Q9XB2mSOvaPOFL+SYthGb0CqkqebhHXjPlFrXpjTSjQmMb3cGFizfr5
4mR2w6Ft3skZXtjNpYHrd8YUebF0ZJfAoF+QIPucBSvZRQgfm/eQulrMsSmqhp3r
vatI+kKY3F9T7Iqfmc04jYkRzv1WSLXt7l2NSHi5Odb2gItJRBvFykXd+r/j+/hu
ezu83tKPqCwR+VN7iosnj2yD9V4DDb818uK8bct/e0/8XyPj/kPbG3J5Qlq1JeBz
C/WYIYqdQTqDlGE5bNyqUkB5RTuAIDW6DQ4eab3lnS76jig1kgKyO9NCIP/vgNgA
A00c1JX5jkTh5ya7yWTKC46jmp2C9szfGnDIHPWNN0b41orGtRQHBgg5YUCv7fdF
egw6iFFAwUBB0IQgOV1e/az0d9gTs3CGlWCCBrgCXAFMcI44tmhs32kNm5SJ9Vsh
+vQsFzIMSb4eDKWPHQWJnurgAJpuNUWOd/qS9hmFpBAZ27H6eBxdwVCJ5DNqp1Me
bDKoUwDv8n0ukmF7pbU1FCqOMgzU+Zxb7F4b7L4+3hYERuQcJKEag0jZvXBTfB31
8HAORKox3F+s4tsiEJSu9OoZCHFsirEWiKuJkkx4GPp+w6BB+Qj5XfwYazhVIhx9
99hcgp26NRpsn3uEDYgi0gA8NpARsuWXk8EwNViU+d2yRFCqguljNweGKIs6ga75
DLjLfE6B5azYs/UDIKFXc5WIomnXRK4hgV4CSyZzfUsp1qJTLq0D695R4ruUFnl6
yG4eML/xIAIIrB/P/Nd8ITG6c4HCuj3UOvMJkZ+BOIEAKYfMpxevSZeDx+XN5urm
e63fdgpdscfUoFmlIUBei6yrmpE7683REB6Cp+Ff+HuBzPMoqSHRaitaRxmEId1w
zrajsxmoP8HeRk9T2E2jshqaHXO6JEQQVLDGWWhj0s7rfgdGhw7834WmKN8Xg+kx
S3n7tjimlD8fCp8+KqRKlPZGj/+h5aPj6ZOr+JqL3nxQ/2bye/TxUcxLGdnpN0Zd
P4gWGTuFWEJuaoC5EamYS5k4hyujonQDhyOwE9RFwHbmZQiY1uE8D8qxIBHjy6f7
nNgE8iMPWv5bcHq9KTl6L/nT7OFp2u0PV315dDh8eiEgEbStBRYAryGPKuRooO4x
4USRGRCccSjDD0UU8CkBoUaqBtpYKo7jq347gcu6a0YVf/ZvEtp0dzdiWak6bBDg
JGfXcVsGMvmY1uMvQNBgUiobAeJ+gK28g9nGv4kpVEd1MjHO+qFmKzMxG3EADPtx
z6r++rQ9I9uB1fDnr2tzcI3KwUoy6a+ASZ09vR/hwAyWXXuP3arZY5rF75Suw/TP
08/O8owCH1q1mjanFnfnyUJS+SnRP/uUbv0ooDST65Ek7/OqrXpnkCu8HQAa26cT
wE1WMzcCJH9k59+4Hw5y+FCKAe6FoqFy38p73agP7h21YFncZdCYEvRTBjw+6suz
B84rYg/ImL/E9WaKqTvWJfG7daCELNM1k9ZcNZFufAaJWG79mWeds+eE6A3Zx9vr
6+iq1y4sFQCnsOUvMHJefvqDQLLwaE9UB2Rstx5j0sfzvwWlmfUhxpN3L/dvuC0/
ZDj6lF+OylA9Oovgfe2V3u6n8u2rDaGkr5WyzBeHpuPVKHUk2fDbpJWeru2aOJ1U
n/85oowR30tlfx8YtTpMQjiFFbJGjcZoFULxVPqGMGgiK+YKSoH0vQElwiRrJHrK
ODhxfVNqbZv+yiocv7mhqYSIMsc1JS0atJfvXVntgMfHdSwL522BeOVPUc7g341b
FnvTUSJd08G2BtkeyIS0BlP5saNtcnk3dIOieXCzMJXeZH/AJFlsx+pjJdsxoXzs
sSbep+Fkv/unZ2HCDHVJqLoQyZEQ6qRYrWUHj877tcrnhhFubbpEGe48sY4Rogs3
zJks0sGKBOfeavqHCNbFqKCVzMkHyEcEovaYUUzkwfGB+jdyWGxTJsFyfLEmIKF4
XNm54DdLgN/p1F5SlzTDDMbj00xb6eVJSbdJd7X51e63D9ADnPkzghN9RXYrd4d0
KbI0gWmBF5xMAvMn3p7xVtSRjvlrCqZCOPULQxK6TpLBdArkQtMau6ms/ezSzRdn
mwhUHODRGnY2TBsR4o54ZpzOBsIkPwgFztN6iTNN2q7NVKz3FRzEpQ40KH9pGvdb
ynuRjWZvT4b6kBQzszHb18tCuy8wrA2gQlv6Jvdh+dVcktiZ+xkw9GbPIifyU0PJ
jdxmKj8/pqyXVfHJBIwpiXzgmPYPIVfKnJLSAYq4zl2tXv56kAmCTXOWGOeTSbc2
GDVueQNztQQzvLwSFFl4P3P0M6xmqppvDD2lLZ8QDXV92osmrgPSlT18ICgpNHTZ
Yz/igMryRWCKJLIbIPYhjUNZfOwsGgwV+BAk7QRfCmMqDzubiA1VcRlcfSmvKpO/
20+hdqPUodcVS4dEuAYVHxoHDQML2p6XM9Usg0eATkmhZXQRTJc7zQDa5jAsaEXV
bWJNiwiaz8Ro/x9o8aV/IW8dWdEcQf7+YHAYcGKZETZZbwgGxe22oYaJaE3lmxp8
N5OXXBdns1+hWjJMNThUA+ujh6B5WXrXbV/ctD2sdJJgy8DI7o6QCVx9dCh6faGn
PFZR2xGpTThpt+o0cLVzSkH8tWRb0PXeEVlMhCfKsY+VW+PgP1g2JM6Kz5dDfSDh
a3RK9C3QARutkIYALZ7fRgwxEh3VEHgjbKI5B9W+iF/iUe2YbUTBWudBSsev+gGL
QNveKxiNgfq7PvoDN6rTC/jDkzZJJMyJWIzlODOctG8vevTdRCR3njIc+1Mb9s7c
FYrFEknht1jXIXuZ+tOMADDRlo4oDa8SCPOuNKxvlwQwJzqf7Ytp6XqTgcXdrvNX
/am5LtKQ7leeFXCTGRo2sh4RZgmRudEmDWzwt/2hhNMEpYpMO4ClKcgJvi5Tcv3V
ewxspUBqvZFB88B6cY5xyczYhwmQ6w6jLSQ5+UtXjsFwGUcPsEi9q0XwqUwLMz78
A5dboNontQK2ehoN06LI1C+Vx5wGdIib9va3fw/YJhNWRRr3mj/Bpu+s/CL4Fg5M
AmBmAwI2sSW3mN3dP+5xBcep2ca+uZ3EqXszklosyQ0zvm2ne6SBeZFm9NQtfabt
5J6ffIovSD6kTgSj6kDAsJcBdgFiyxAFVogPr7v04CfajC/0VdpnoBiHpYBJF+Du
sbMKeroWdK7JsZVS5T2n4J46iF4qjQFWM2m7OUIsqUDtGUDhkXAobuCgVapwz6DA
luMWcmp/pEq/gr9SNQNuFT6av9hcsC/8UJaWsp1LkO/68homWelrsw4ryGeuzIvH
GJ7FT6GoIU0ZSIYVez8l3wF+MKCwjRqN3CSqlaoKF7zFQRZUPAwwFAYCpctGnVXV
DM/kYWf7a0b2NMu6SzsxJJL/HCL7Aj4l8q55FMIifAUjZQhQlyUQWV/qE4cXJrJS
36KEsjbgm7Dgh96cyfM9oTRkQagfdeb9P5FrVAGMxQfdbP1wHppJ/NEMS/3Ql415
fPgI41tU9qKkUqlvPexAi6C4AtNw6YSwvnL+2AG1JyNS4AaDxv/ls6XBlDeM8T/v
gKEr0w2U1BvoYPZiytFwB05ZjhQ3Qv8wfbGg82QtciK2vsqESF11WKPja5iQHyOz
HZE8hUBPK0e01GSd2OcGM5P3mQbXpbXRY5BBVh1Vi9bo3Sh0E7TjFldVVP7Ojg2r
nBpuuQzxKM8viIbWEl6GiBlI098dfJXfMSMhuZroJmKjR0PqVlGTO1+3LM53kXHx
oHctkxJgiWfBy59GD13cyGeNhO1/8mjtG7xmZUJ9Rx+zunVrezuLphSt5UMBoAyO
35XjL8ixCuzubxR8bGkuiA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GDUve2rG72U1odYz2xdjKD/pMKLmwl5X6DM58bD4xXkGPdWMD0wAVZdrrQ4IOdJk
KpgAS69B1iUtw+eJLSrlg0X+1gEfLfA3DAgS8D45Kp4U1YJdGn1NVz8GZiiyQ1R9
tqSjEkYabRvsRgkiv6zhWCz20DKbTfE+Yn8zOxBdUojINy7FzJYwhhbO5UWvbyM1
OKdBwyrUYSXqwyhQQfu3yiFLQ2NtPqC3c2WWyUd0UB38IHb5Kd2jd2LtZzZZC2MH
vbJ8cmlNI+b30Ln4zvVj6+s2Gx2hmO11YD9YqpBwacPkoV01PUuI0fqJctFzgdXp
kzGwEHIYCBsA4WVtVXAMcw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4672 )
`pragma protect data_block
sJ8bIlyXSgdCLi+dmCiT+bKGG/87F/Npl6ygNhDWNGOwshNluObSlS4eesYF5j9F
Ble4slhW08nqoMJuuFAMuN2JAEpSygK+ix/2bK5/7VUf4qchzpyw13bwtFufEJOV
CpWq3/zeKztzVvICZzRIfryBaI86wYRUowMvzw30gJgr5nz1RB4QJMx7peB6g/bM
B3mOVcOqJPHW79eO24GjOwuxjzPP3wE6A/Y5p2itce9XTyYdz55GUKZO2/DfLNnw
1+YEHR2NtFw/DChsdD42Mt7XuDzhp8mTXDQNkePhY7SBKfjfdZeADK/iFa/JH7pW
LeZENhLboF5DfAC9BtpsEnwATalXmEKsQva5z3NW6je36VLRI7jGxkSpFuiWaQb4
X2yYb2xGVufJyZF2wRBsdjyzy8KpnkeLxOpaIr9NvjB59i47tntWYHNBOF3GGr7i
QCeq6DixWo+eLHNaJu6FMlJO8PHwuTwnbhb7TT/T3ipQ2YNQltoLocA3TzS6rAZo
nKxgTsaUvWfli2w1D6JaIgYuvnCBMHIst8UvyjbHqXgqOAl0wuX84xRpxIRXTIqW
YL7evvvVCMTwoiG3qgb7BkYFqeRhx5ZefowdqOeerG/ZfK4oyd3Vg1pwotgLkdkF
xlqKxXufIL+q1F9UjaJ2WhdZnHTb3Ks/NdPAxcrQy6OVy/z57LJ6WQKIDfOHoCkp
0idzZaBKsuh6J3afB9Mrw7+NCHs3coajmE1WorBx1RP/F8A7RtMS4ChwvaJH7N46
nSEBd061nOWVu121zPDOgWbs9PVmAZ4vR8Wn6w6w+j0K+p0620ISRXpMv9/QfhCx
hcJW7X5X7rP2PF+YtOhu00dQInrOdqIymZwQ0O48JZTp/SUAnELV4neB2tZ7cihM
e4+ki2ea2E5v/hXkmQXJZs7omHAMVMqX+klpjFAKR7iycKjqKThE5nt+8uvU983Z
iR4D5x07T0MDkuikqGglD3ztVmF5Q8TS7aQ1JesxbSzFyubWkksGjkFmXoshYkWO
8iO4HAxUfhIAWLqFLoOSl3f/kgoPLKe4Yf1zSf9liAk7+NO4fXOeniJttYDt1IHW
MTldgYNN/hEkdsaXiRg/B9Hoyn2hIXPl3Jd++HWfOmK8QU8IyIsr/Lib2hR6v26M
1wRC6Hu7qikLAlSc5SkX5VWISoIHw4iJn+AXaKpDfyn4HdyHawCj/FWlTkG4eRea
Wrdw9pZOqcUEsaOpRh+KOkhuEC4VTS9CGbU7k59/9B+ZM9JUSJPnKRHETSCmP0d2
F9I7GFbgKPimGmXUGGFOhAVtGBkyU1lSTGSP/JvMvFYqu7l+JjCfUwShaeEDnwCY
G5CJXX7R/CvS2gnrZZfoIDHhnqkmwLay+pQOgnecRJLOSaaCspAHo7wJbpkvMS6B
lkoJYbLSK2rVJek6rxglkvd6U6SLVYiJaVjYAruK1WApYwaz34FTaMfvDCwQ3EC9
Upp2d+Db8WG1lxFc51MXNRx+0zWwWOhDzb3EPeoOuxLN9nYOjLIpe4ZD/uNlfRH/
Ns8w5ab+5FIVxOMa7Ht7sPqXq9o7n3u8m9Rbp5QGf82/jjNp+sQYASm+RYsU44nG
3fgt5SljKBfgvF8q3DvD7vhR42Cp8L0OilEm8lyr2u11H02aty4cVSvjQ3dBWCAL
LWMKeHVFvjO85J2tVNTfo8gVZ8Zgs1Eb4lPnGc4ckvshQqdzx1E3f8nN9Ql+A/t9
iHy1khatJ7dNk+jKOS/E2bLovrNWuSjcpcJE6S2udiwRXi7eA8wHMTGpXL1qk71d
ocBdnwEMysu9q0Lb/1MCod5VWtkGEhN1gjt0RgjxURJ2ZJX0Y1eKS6j1ZYaxrG1I
lD26kc1l+0lP4snCPLnVTcRloFv2XShVCMX9d697hme9otEN6wpfZkFyMOfg9WDF
f6pzsGM/9SsV2+fNN3DUIF9rYYlf2vg2YvdeVA0G6lMdp/jlwsSzmvTDTXF+Z5a2
hl/JGG1ifRqqtKJw6z+aOygcr1NgqMtGjDpX1hu9AARS/zSSG2mWaBnuazHw9xEd
oVJ2UMxpL0Xfko1OkLQ0uiu5XRQdulKE5zQqGf029L0hg24cfYQIamEe/2X0nN0S
X9cDXmLkHyxKqZ8ZEBRb99XUKNK4F2UpRxY8QydZli+nGnZ5lZ6p+9/b0Gwub+yF
TsJP7WJ6u/REGMtTcZ+IgnVh0srlV7Jub4QkG61UIkA5tiQP5liPxZdZGHNfv5YY
KLPEY1wxrtI/WzQMz/dELGfiUHMmwkUYSSa7iZFxxDiOCtW/JYw+BORRCZosisPI
Ocx+k0y5WT5segzsHQIrtr6lwO2vTAIKhDKCAkG8Jo67f7Q1ipn1res2gZW8tm5e
7+ltpM72YSM69pXNd9jwZpxlVDLnGwUkQ5iS6SJSUdrm2BzyRECUhFaKlShg9W/8
xqRNJWhv2SU17z9CEBg7bdxly4/J8f/fqFnnsjzXsAJvO8p/Xrc0EVGa8StiVO9T
XgACajl7AcIvXjIQvaL3cUXc0P1r5t0HY2KN486QyOW0VtdTtPLsn4B/weWedKsz
8/ZJ/1pPFbyhPsYDkUQZAYq83c1ccLdRY37M1XhOt04QEboWbmuX5+nzWUMC1hq8
YizIaqWbDP1z38guXu6FDcymkLsSR2qdLHwL2Ru1RN5xXWzTU3Izlo/NYLhPGWY3
+R+lgMiU37tfObe+0bK8eaIVutsANp6L9iBGEsql8LZwVwuVFjnP7gMBFUvf5963
mVznMxMzYUfSbEG/1KLe+AR2PGVQfUQWhcmdcdcb44W36+e/0nBavSY/Kiax5bA/
+UV4GEqftXrJDDrhsuvEh7HYZ4ghg1Wy2xlzmVQNq8sRuaxVD7Zm/8QYKek9YuK4
5SLm69ly3qAQi71xqVO88XGquRcj3+rF9BJEa7Dt26Fxfge0mKe9N7A85IRgIWS2
+1fbXZLVc6DdyCODfOKnzquB5jaSkdeKbYJc7nSXeMwl5Nw2sZs2moainFd/8HLm
E9J6k+Ty669DR0RACJJua0sRzk36rW6T9jy4HPKl3wR1aOZe1YmcFskxMDn5iRk0
Uz0Xgv3xbVw1q1OagvzzNr5pqRiTD5MHTOChSg7RCSy943s27/9wEGNaYVUNRCeT
JX9WrECfOWN3F1JYexnPB3dYfgUwaF7/7NAWqT+ZAc7RwM055p4H1uoPhJ4wmf5F
+64Sxeb5TZr8eMLzbX5lfbi0m2moxlUd3snuAQrvas/xeAKe7WZ45tVN0GeuJTUK
DxZX5Q0VqGq3JN2jIgKM0W0yP4kY9o7wszo0Zwmx3qkaKiVpYo9HAO7aTYsppfmk
qyi3Nx6nWF9+Ct8Y/BVxS/wtKU8DdZpRENTreqNlJaByW1T0ebwWDBeB1fkw8koL
cn2SjUvWa/zMeH/dtu6rmrXsFKZ/5ostlaJjt73vw4HbOwgCeb6zEGrn4sYQ3zD2
2Q/Nn2xIat/r3eBbpyTUxKvgFn+/mG9a6WEjm/5Q8XcMoSFgi6n1P3bP6q9vkbvv
QSmVFkoFZrJLhTvThdQN2PzBHiM3XnccfriQ1jgVOjCr/+wiDkMKt+3Nf00iYDIo
reUyzUXOMaEshT5pTrv2mf+e4ncWmC+JjydxLjN0en0OOeGYiKjPq3S3aOUcLbsf
FAZdEP+HiGd1KTCl9q7W0iXsMQqIWtuoabvpAUYbvUgKVNgDcgAb6doAGLx1XKdJ
sGcB17SO4VDSKUXKSaTQtXi0QnVNROZBqZKQLFRq60sJSa9qIWRVr2/2SK3B7tv3
q2IPkY8VVCGNP8N9nwAlO9NvQluvUV/Vr1a4T6HGASFwalzL7m8X5OyqNbZHrorE
CAx4aVUSIF4BhB1ra45wXOTuUxUaWZVUAeEUWntYK6q/RB0cv6/0hl4zd0JJlmpm
xVRhXjfImlJAwlKhTqe6i8bQcOBSqGfRpM8pvBv3A1vXLAwoxp8hkGBLjbbgwEJL
o59zdFVGA3rGFqqGlT6zyfOQjVp7uO2PPZ8DY3yI6eSbQ6A/afZHwLyPwlBixs5h
NHe50+/DjJlyCqGZU9W1sE00nF5LnV+9T+yK5S6uv7eyjYCL4Lf4IxDibgYtTn2B
YNHkTlEtlkQiS5fFfMTFdlJm0/QfJMOD61dXn7Wc5VxqRHLs+QwZQ7r+p1nYys6r
U5Y4q2DC7zKPuYsUON9WPIpsAP8PSdpcBmqNJK1ejdXNuj8xdDri9mlK4MHsL9A7
k1KlQYYmJvYNOuv76xHBHNSANyY+tMQX8Z4di/Bl61lqfQA1juf11zgwK8Ado+uC
XxoQpdOILk0oJzbYiWJBlPmnT+tYiNZUkF2BdKNUnC5WR/1lvUYuZcrxDM+OjNpY
noFI9+GN3V25kPT9ylPhi6SEKlo44oIiofZUA4l1I/I8z45J6RoQNbp49dc0r32W
HRpUd7T8kbSHqrsXFqY/OA38quRw/TzyFgw5zHzxKAoA8/SVOBb0ksPr0BC7itys
j22TwX2M9z7PKCPj7XUO3+qGkNvm1LGSS18wYnuBWzw3YtQOXFVn8kCiZ/G1uLJJ
S4QaIjiRoiCE/jqA6LDEHDolNjsCrrF9KDBoaHcaMvxDA1RTeOT7ZLYYLU7B6IBK
y6Uzz61j/aQf6kAnYjGsXWqmQN+cvughgcnLg8gNDZlmF+rDFCDtN+L04Koa79LH
AOIv2tgCKzWy4k8D96N2i5MhZe4MYHes6KEZk2dwYPrwd+TME3QK+m45dPp1Nn2G
cAvXPBwl3lvGOQZDW2Rd9mJYx3ET7QAwqMqmxNtA7XBkQavIt1p+kbCzyaXc3vJo
TowFX8jFB/ivjZxfajI+My055O/aFPiP7PDeA8OZ6tY2e7VUoU9FATRSxd6UykYL
VEWBtsUoWuYpZpTX9bZNFApMUaWh75dDM+WdY22gciRQOiMtrrOQNXP6n8Ra5Hqm
0x4nyYX+b0aANASR3co09px0GJWZ7DAGqnAtQoS0yFfqJ1YyEhGwn6Mn/eEbRsha
ogAeQaJLHhs21u1opEgLuZkMtfq6SeiHpfqZf7H1uY2ZTvtJ+vEiqxG07BLsGbXw
Pq2/eJSaJ+fxiicEPJcPQIkag6SDiopY00IEE8rnFFZWJfa/EelpxGuCRVvZiXjL
GMk16BF9YsUSDxDJV2Pf1t4L/I2fG7RMGrkHRyPPyZEN1Wr1p8M3DC+ZZzwnKP4R
n+yMFwjhjQ5fNwtf7NhZ1DIDcAv2DwLtTyaX+9lv3KGVRPjOH0FJ2yZeQ3yWc/Go
2VyxBO0WB7rNyRpIHdOKkC8GpkNipAENVYPZrYcAsxUCkKMAdMfbK1iUjyaCPKqA
eENtjnF3dU2lUWdELna+NBoPBFcFcgBGwBKC4HUX+UFjtcf8Vm5niCFOZ6g63jod
MGwxQ1EFVTVV7vusuSg6bvZj05Z+yfhsyvCGa1QTMV05/bBu34kUXM+A56DaDLBI
VSRos+uNb9z5E+BdVIVRJO9LlR9Wx7rwmXyEZdXIZLUwf6lPp4y+J1n0Mt/4J5Ed
jrruxDWcaRBxNKsCQRlJ5An06T2abt64KXw//Whx161HstqEPFQa/TgHlZV+zihE
QpRIPG+0GcnANKDCFlLknTmrX5r/JZthM00jL/lYPhENZgs/K0XYPM/2a3gtDu/h
oVQY8b3huxG11arKceQdcsemx/9IbGfiEtpFsfRIP+OvwX0iO2Y38n/GqkrU1pae
E26P/6egl43fB24ITXpJhZavgkMR968IyspmdPkjMom54TE8dXHPOtxq8siewG2I
pmYCO1LzAHTcsrXLBqUEXrGCGTCRq8rIK1jvNRQrTod60ywKObN3mCMKigm+5Byf
6wG63VjrCcpKgh0D6wwLYNOOd7q1FXRMXIWBRo9ju2vJDCjM0E0OncDZmxn89Ouv
jsOk9UK4jSjYb3G+IOzidWdJtDDrLBTmcKHOQPwE2BlU/yyHvykt4IpQ4DOZNpo5
vYWoqSrHxZ0xZ+YxOhx0W09fb8KdUqxxLUGZpS8nBaHV000kGt1QyDZ3FoZn1+X1
4kLAYO7U4KtftEbB92Zbbfqg0cmJaO8zwnYCKhuROoS4YIx4T6mCXhVs/bqOj3ZZ
3GNzF91sM4vaGL+ncz4El6E1mOAPJwHaynET7CoW2UTyTt9/4eoU/+O7MzXGe9e9
xuKW0TqvWcZzJ1JDqV85CcuKdIv6UuDHLWYT6Nqs587f0UupE36WsFCu1E+MtKkt
wsJD+rVAYA78zZ33yIBYeA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
fZngVFobkxwW5NDGLQTXaqWKkzfNMNZiqP+na/VZuPdDg2eBEjJsoQaoGP/zcBOn
3lUcoK/Y3xLprftm4BvACLiGt5bUsi+UA2at1eYOPn+pp3RVR22UkkOy4VnBcLHC
PpKaxzhWRTDA2TSaS5M+FmwDqz6Xli6VZKCX3gjPO5qoVDLX3ATXG5cyXo4/t1/h
BuKUAubsIro8ZIH+u4T6gj0RmLfvAQnZvcZVDRIglSad/J4Yutl/o+Hy3XM34KWw
4XcRVKixMTgOAUizPmtActcKoTlaTnplQje7GHJfDBdJ1GjQ2xaKR6+B7BYYbCMn
M0MM4Gg4COrSmyKeorY05w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9344 )
`pragma protect data_block
yp6//xoJGnEwWN/OyC+vSV6JzIbrZK3B3KAcQTlna3XSNne3ubI+dx5E0nxe1eb6
MOdy6kZbT7r8cjX8S3Fo/aEQZpj8dQVMIrlF29hwSlnSXRiIX5EnI90a7015jO1r
fUvd362687aur4UbMbDTPArOFVg2Er0GoIYz8s1hzwpClDktFLVOfyExzMR2sjHO
GHeIW2daOeSZfm3YKrJZiUPf+ThdHaWlvgkV3pr7aJdeP+a4MSVaxptfGnGGjKI6
+a4yrIDMqL0qjq1o9buDliDkYFKMFf1udKW3LTW02PdiYeBhXqqkdYbjNGUIKes0
inqp0DhS73/+X0htyficJ1+qt79DxD4jM5nJ6/phjWE0D2wFENvAS5mjhjX3HnxP
j/jcCCoM2cyAAZrPMMCF1R+rxcyZ2ZlHSHvUt8mJMbXLyTwYk7vtYnsILlANkKMb
MUf2cJYisJY+V3aIlT5MJq9eOU+YzDl0DYEdOXMGADGeZeMCHhnsMkCMEsfd16KZ
dGxhw+13GIViofcI4u9Q2JDmZI6zrnAtHbpCFW5deYkbTJy+SM08rYqukQejWwr9
uKxBIK6a2JtWWBEEMntbayY2G5oEc4ws0FOJ9qo+mdsPjupBlRf879YLlWviVn7r
Vnd7rFYM9Fzc8e5xffdeYinIfLgoSNNJZTB2gr4DFb7mX0wMLwcRLUZ95KpBltmL
4YC9Y/tnerNib2wAxUv5LnCJrPPkEUBesrfPrUEV2WwEwaL9Xo0/KIfmKFKBKwMs
GIpnXYotjVLDEZaLI1faVhtTKrpyT72WwvFBK5srfuH78IBHODPJnyMe1/eLXr1N
znio5Ew+GXZ7mN/30Fp/ymGMx893YrATw1MP80P0JycyBPeIgcdpMbR9ohdGYrlp
hMjtpM7U/Xde48Uq7qSNwdG/ra1tb00IqgVYlhEoeq2vMTk0F5m8UAaZNYt+MMES
u1aTbO2NOOvzs/mow6yfYsMUtAcf/5JCBSJYlk0NeVqIHIOMjjzPpF4RrhLcN+iM
Mv48ocSeO1n+Uz9QcEMhJkUPPEmDg+4e+Knkl7T7Ukg/RdC6fQAYdEVmseYX2qXE
2A59u40terklwhTbpymHcBiwLV5ZY1LLvA3ApNVTs7RZoM67uQ2qxsOFc2adlO9k
w/LmgX2PWabFQbpi0zPoyLJQUX0wTgvXAvJ8/luWZPX1oAF+WC6+O8xqPJfylynK
SesJN3gX/tStK2jeNw2sAaNnjrhnRVjvfbbv3GlTROu324pVyST0BjSqWF28mqy6
uuEwiblxoBoy+uv4Mb8m8xSfvJ8kg0PoSmgjQl7GlZN0HAHkX0fWOd4RraFsc4kj
36n+laACNFhslKLiF0I4qfiVlne7fjC97kbe+qtqi6z/ZAC+TGrgTsVKuq3NQ8me
jCbA8J9QBsn6xvHbGiC3ApcrPMKfgfeiCy9J3lKH3R+H7Npw6cmI7SV/Yi08QbJM
kXlHTZcJ0yM1Hqmq3R2FniFDY5zYM1gWy2LLHGJOXCwb4mhlF+B3KknYbSaPw5GC
Yeacrrb3W5lomRwHvAn2tGpupr5ec3JcKu7AapmaVUZ2M3T1rYgnOJAeoT6Bh/vI
PercWayyzWPQo+KIGqxGN19hULjcy5Gvl4gYEmOrEkLNwtrjfKy7jmZO2nKH9nP5
Oc57tsBIGDSq/iSdVAQRuEQ9/3NwzPN/FdfMG5bXWDSabsvsInQKZFpnZCeeizdP
GRFf7NE9l1C0q+ly+CN0YSg6Gy2I9hygEtmxM2F9eUYJCWYt08yyM1t3OPQBK9Hv
b0GSoJHLiDSzPY4JZA79JYLeSLw8Re/1iHAh1ZHd/kEda9aT5k6HFwmU6tqcUHmn
3ZgQuIZgKgRNy8Ygik+8j7wCbGmx3RN9F4Sx8KKCJ1ffWxcS18bzo6uGN38aiSzz
3jZ2nmk5YlRHP84BaosYQvq+d/cOQ5f2U1dXxIlVqcj+fc/T1FYi6mTCUVLlp2wF
Bo1EYPv9RPsydID0uvvN0IagT+3QR2c4NfkQ+z43vAhKQSnHaUzDONMg2iiNtUqd
YfmmguoLmClSFD4rH6LIck4RUbJ2GSSv0ILh1dqEL5FJUWLRKT1ooytyJmTzPdmo
4cRKanJihoRWQ8Ml/V2MW0SemU2qpyxOEZS6aG6ca4kafcn0yaBNa9sDFoR0KrGy
w7uPrn2xmjkpZyPbnjXKmuF1mip0aK3P9SI6mSjDBjtsoQ6sdpIl26YHo3EcNQSS
vfnFi6xTBhFAT3AU0VCM7hrNSvqQs6rwq3prZ49dEdphbYrJ0Uzn8vZLhm/o/Wle
zq8hIbkXaoRBFmhLGzkuG16uQT6TCyhXVJFH7XTq/cyuGqYK1yb2g6hrOZYpqVqL
n8ttAXf/OMXRyF7cal+X+nUtIt1FaoMEaGWxr0RGoKSD2vcPGwp42+u9NSxrIP33
8Ttq3jgi+41pNTHTYh7k5ciVO11eMPsUlGgwS8nFDV29GAlIckpNBuPS4hBJ/cAl
JjP8W5n58gWC1T9atLKbfNWa5G4ZZAlLK7nH1Dlhrw8xQvtju3LBoMW5lBKEPqqs
uZlmEP8IOQqt4LddY2IHfEoaOasF2htfAH7qEq/0ZZ8+O2OdITSSw5+pYQBqTxzH
YfNYwsXgOzrdSS4618//DnGmPfb9hR15itO1ifd/kAemuX97oTcVhLmPVLNAsGL6
JrUNa9jCxRZ0toR8Wxizi+LjyAnYJttL/NkSu4lA/tK38QZnVs7lSPsXlcTjd2GI
15d3bKTj9KbESbYOZcO6dCX9sjcf2II9iMMEx7W1lvgH5ZgO7y9SrF0PbJxAyenp
kosskS3OrAIwvkB17pRkXCOMgENe9GcAnWrUCMfPAdO720i2p6+Yl2b+DHewWslw
IbESkojotwU0+izbHcAl16Tb5PxnoIdiPAHMO3HQh06zqPccUp2j14FXNcS3lZBa
CNG1Nkx87JIB9puKdJCv/qIxpbxI76PyWhzp9cSp31ocF+yhNtg43KFfNygU/XHU
QExQhSM1017fvEv9r+cYUtdIs8TaiCQjwFukKleuezocMMXqqHe0z4ACHJLs1NyY
WA8cbgg1V0yKQFlpGnIWV6ragGoqSiJ8H2vpDJwnH9FzmbOHmQqlbhMdkLfrnVBJ
S2IjRKaiEap2S2+7yE1yQmjBEPFqx4QP8vG4L3Fj341hswsjknlZCgDVecl8X5GU
R1WlYp31YdtZma6GKbv8yR3b3rbsQvlSTlj+6UGMDWvwvsyGAuEl+07BQMqxu8GG
UEojpVl8nhdg3vvj5ZV+KmQz3+IN0RC0oM7ktCcRz6DkPmHWGSlSVmfWWh8JB9eB
J3XvhbfuaS2wvdoHOptLkgqx66a7N3GemrqrtOEU0Y2WE7arBs6RaOWbyaBHdKrx
/k/yGLl83iOvt05lhG3T2FgETSTFwQWTuTIQplYCjyPSJuLNst1Gfw4V8/k6lDi+
zIUmy+sPZEcjnMhKQWlAQEil3pKb4LRJO2yFJPQzK0xn6K3I1/8dX+ixaYhQyhDT
F3rjdK5rlxnlgVstRnfEHB8VylMqsJsUo0rgamP2kgVxVJ3q6GM/XA0bpcl/9i9j
U+Ka5bb+S/CAgyQ8hPJH7/JYWr8rGOEoC9+AN7KS+IlpteQX5aW5ryK30opE+ivG
00g8e4wnejYSV3D+LJcNXqI8TVegh57g3263/5xRHQcLqX87GiZZ+MHyNeE1wDOd
50udU1PHsgFgpUuqw5MdLUHMxu6IjRn30WXMoEHrUXlKLJdKoxGO77pmkLGuMwAF
cUtvTID7gP/i/Q5VYFmb8csklkVYt2/fIIxYP1P8Wg82l6pGH5WFn/lsSpVkGvE5
zdShPIBnKdKzgakO4Mu7YqUnxTJr31MCIDy0t9UdOSVriOwWNUpHVEJI5/MdRtQA
r4L/qIz3rHZeHYqioolQsociO+s9U9chgG1Micc1pQJoKKpA3IzDQm0jNhCT9KID
+uji9gfUq7LtzbBCfYMPr2LFFiOKcGBXlw+sdeQpXtjkUfsHwqKjkcwtkQvVegxH
oQwbqEFT3XbHZxaOavhz7Y8tlrD72v9WWT5HVAmAVTGXJ59pHQ0srzOdB3Ao3dX6
MmGhrRd8uoJoweJf3TDIr8Bxcra7rN1r0Na0HJtRfF728DfBCP2Xd/nqcVeatnbh
ohNS6ra6V0kN30mIGtui5HnomKaEmCupWm2OdQVt/9ELHpQOSAU1oIFLOGvUBtPP
aKKSppSYO905LLreIlucZuRZF8f37sdN3kObKRf4+bho+tEygtixVTzrcWxjEPCz
RN+tnK0CCJzOqGXef6PU5kWOM89DP/V/pNp07QaQUJIqgkw4l/o+b3YGqfL0Vnnp
OvgemHyR6qDgkpL2K1qP02d1QGFtfih9lBuNLfEgBOma1R8V4PfPLLSxq1/3L4qM
XzKuwLRw9t/Q3S0GPZfxWBqcFxh8f1fM4xQKb6i0Tm6zccMo015hHi4x3NRDIgBp
ZTLdNCQ3/luUMx0qvOi4BHtfTHhRu8b02BM4JiqTqR/0FWYHH/KxNQKdeVHqMbA6
kYtbwcT6Ub/MZC/KDPCYmomVJwIIYwKvJPPGb15c+fcvEaQWagMDFcLkWpfRVZdP
OK1J0vgBQJoeGyAENtpXZlXAC4/upp3qfc5ZzDRlHORV7viFJvNIJEjW8bSbBEo9
lS3D3b2j5Ys1ZyJmtv2IRPXYQmGoP910yVxlmosp+ey0nkGk+uwrik+HsfKCbPtG
p1d9jcEPEY/FoxHxrYXP+DSeFc5sgd97zJHADVtWYraFMiKpphsi4RQ9h5D/HfBh
20olzrYdSplxRftZOmqzg70shjPkvNeLkF2gmk8J2yqvzPkvZTanESOW6vBh8chh
Ad8LX4vSvpp9lMssYbNdVBOqzBZe73rWNITYd39cM2xiXzmUH5qld3P9wzSqHJ9s
8zjpMTsRNA4XKLP2rrdv/Z9X9mIMeoMX9VKbAWHaPDCgNinoevZ8/0icyz3Y+TpD
wU0dbqAsKwtPAi4UJe2VCfYKTOPDxyiZL80nvrdwrnGINQc4daYRPoTLLODyM0GL
dNeK2fTRUiPBpDH2xJRAXroIccEMKEIO8SMRlGVoxEb8MZOhsgW2ueJ5OmXyEdBz
/fbRyuy4SeUBsnJX7fzLPgkXEhHI/R0LAO+/LiHcTCEFBvLDt6YTPbRjI9IcwKzv
QSxslhh7aFnYv0xs8zpM/FroO1oPXi8pgn0ajP8l69JLuDJtdsa0CyxQR93KzrUC
SR29V2cSoL77yVNjxZQ0Ey/jxTw6qnp5v/eqEtFR4RI4jS/QPed0h/DkV19Grxk9
6Wu7fCHNTc/GLe+e0GjxLSJvoyMfy1KTy05rGhpmYqXEkNK+sgXEJLI1aYNEtAX4
TWIjPy3K/SJ7t/+1MU5acpAEzMhKZ7QxdIYTI2ItDYLuARhNEq/s8fNT2GFQ6Iiu
s20XP4opcfnizRVJNADTZzt4zgYK4Wlmf59Dlhgz2s94l4juAw6n9QvQ8MTB6hs3
XiULH5bBsCr+Z8VIVAi/75qPmVPh+OLz0JA8kCS6keThXPAsBb9nnccn6ulJ/VP6
wSH4rVyFPyuEY6Jz2eXcNB3PH+nJESlkN2rH9tdnWZi3J7L8VEfOKsYdtlDEGUC5
jGTt8KPSv/ax/8ll1JynWcOo1gDhT+HEGxwMI1m020xgPe9ZosI0z8rY7/S4g1d6
9273WUnE8OA7dZwzqEIrUADMBC0vr/EyBZJMbVtxl9vk1Yl27KBTIWV3f6mPsdoS
ugZvELEw8k9GSDEv4oKMa4CJLyZFasFPtR//FZrU77O1aNpF2/9GUkdtVuCnNiKK
EwQWqmG6+EYWkFFtEK4jf6WKP7f1z/FfqHWlu6UDzq86vQPLuCLj4+pdy/N9SBpZ
rSVc2UBu1GR0/aSofUUGqeiQpitMJHM/NICa7pOvNx4EBRuhF+oYhCryUjZsjnrJ
98+hD29PbL58nGV8fovslzqm1TCRYHhPpXT1djY8yn1yBvsCtFMHx5zKfJmQkzhl
oIpcQyDvwWYYrhsNx3WyQKczJAuzS4+iFi9q7Agr2OYwUWqsHlm2j12Qem9yJA6I
NLAYF0SvkFXRDJ/eAw6dHNY3c89OMKnKCo1oXpexsNd5kRGFVATaIQRlq537n3JG
3mNNuft2A6nP967baAMaRtbjXJnvievA7cdZTPVYfcRN7Pjfcbx0bPHp1oCo1OXw
2NCYWk11/niAKdFrE0svHbqBulD+RiCLGKP0dDFaoA1J5XpVMnkHYxTiIXuDOXox
bb6k0WD1R4tYbnmZiIrJ9jvFnY1/Gwpftxqowk6HvLG4OMt0+4Nl9V4HvTxXVa1y
sEDpUf352lK2yz7J+bnYOZHnNtgwA4mcv7OFplBHOxjtbOeLIwIBRAqt6vqEatfm
weP/1pBN6WXDmfp2KtpLNgxiRXSfDK5HK6dXbNbDdvSd9cHqDbm7mLvRL19PL/+8
X1DlrS00F1bxS706IDsbOavqzY+cYuFF7epXvX2+nOqJKCmVmTewCZ29B8lMaOSG
TVXjo9jBpEfIDMfL/7T4FH2C9/LuRDXVBeB8b2NyBwy+PssnzF3a0bpGTNHRCtDk
NeBXmSi+pFcUBUmRbAqbBHFqSd9E6PT1biIQsQgEtRCwSqTLyLUahyVYBvbKmnAA
/BAWJuUPqg/XYKpgj9tfYcVhji50G+f4NcRal/c8nzrh3FktQFPdhOV2CmcGhyBv
eq1jZFJVt1BuLSNuD4wj9VO5ICceDR4LLCFZRcuGGzXUeYNxQPzDm8Um81Q85AkJ
irpUdb4hYseuJddkrEhodv8dvPBpBc73Cp1NNPzh1asytGOl6XLc7PJS/0FmThsX
CmSTPj5AOk837O4xgwPN+JJr6x3eHb60xWQ6M+NIAmB10JSA8d+kWmRBPckbvrqo
tbXg9i3Xj53y+rEFCcJv7NgiLxBSUxMCPvtQRxtgckWReMzglW2mjKVNlvDKDijz
21IINEQ9BrEekZjuG5mCoCXFB1JtWBGbLFVb7UKUlcbrO9/WNJ2W2yMR+TcnGdUc
fpjTD9A0Nh7S2fL8RmcQhZVZWaYRbX8H04pqQa9rnFq0agYtTsKi30BVEu7PW6oT
4LUEC2xbNR8c+NC0N3ALYAbeqiVKjcKcyC54Axne1gb3wXO4ThTF+j1koH0sduTZ
onsj1u1686qME5KY4SOF/hw+w81ffwjmX3V7UyD6a2OK2AvjoYZKwZVymohg7R+j
26fdHdx6uHcn29QBrEUXnIL0FszL0FMKcmcvWAscDRpQzbFQgBHNmhHKwLV+UCZp
GGkGYtV4OZaW2Y5QscWCKnYTXcBUrJFYm3npHK/6+piJkQfOW0u6Q4zD+uNaxkYN
JQJkalHN7RuTLRNyKjhcnu/LeEEWFzKV0i3m50ubEsa5cdk0wy1EqQKZWIm3FV4V
L/Phjr/45NiHGhnLROBR2JFMSiH/KNOewbyIet88wxOTKEiK+nvnxdPK5ozREkH9
Ev+wGsAhfIOJFd1y6XL9ynav42HP72I7WU7c/WEcYTjFKaEs7MFRs/qpvzQKzHfK
1otHWCvQGelXyTr15pLqelxZHpWSS5omN82p1hdEHDgKUMq9XOTMAgU3jvz0xRco
LMfa4A0TezOb/oU6r5Mrf/nxWddqjjqw7+pLO49zkB/NaLsq9x9fJmHFBGzkOrkG
y/8F/c3Dj+6GOtZOipLHjl77hDBrJ46EXA40uG64t0+HH82dJPGoz/zZRaldHl4N
Bhb+2vCrHk1sVKVugF1qISxDNOBkjEucu13IAAIYjboozZT/9/u9lI3ZT4481K+r
+RVKMyI6IPBkGGxOBh6Sj9JAzlK34VKz835yRRmeVpuZ2I6qS/ebdiCR185/P90+
e/wBnVci2Nny6LQqpmtA/Vit8IbAN4jYv7K7irvaCAtyfhuR+K04qBfwYVjJfVa3
UmgzP5BrXLQcrqv6111d8kS14OEhW/zbpEiidrVN7yJDHHIylpQ1ggVslB4coFVv
GmAgioTThJi9EBCr2+j+DT+jTn8dZZGRhirk/qyqoU1iKKIqOn+z5nYR8AKW7cCo
1nXC3vf7Ggul5rUDv49A9gcZe5d1/Ndf3RJc55gINFtYI8MRjT67ZSAfcdtMJX2b
Akp8MKfetz82OHsnKwc2bhTRoYJa+SXFCAdACPoINah/7K0WlbvQnypnBQZAfY2T
rUCWA/sH0lO6JL4an+5kLFL09mRopp8vKqGbgORJqlGo9i9GRJ7bJXWUKNvPhddT
HtVN1Se4X7INgY5P7P6A1b5TaU9H1lBU9r4fLXuSi3CGIihlfJe0XPKr/PucdSr5
IlbCSAuuxo/1QAFxsSAfuc+TZpH6eEBNiVxuN+3F6tDGXbiPQAHGA97ZDL635DNI
BjV7npBEGQrkqM8jBOc5ETk4Lg0TqpcwaYo70bPGzyVZ+ofSUs9+xpbuA+/zMTEx
gOmvqpdBmCNW8DugUkUlGySVXoAWC7SGDLWdA4qFNlpi+nV1oN1Kt5sL8RdOO7mM
nOFk1Jtbj+KYfsha3f56aqdtTJ05LI8MCN3ofSIUmQAwK1/CHhVmKbD0Ca5mlRal
rCinZmZC0Ji8vvLlDRq2ZZckypVgzJHuy7WLmRxkZtDzUt/92jGlqpV4XckumyGk
ns7MuwCdrqqOIYQiCTWUU9yY2cUdLexpjW0THGYuY7dAWYKe+LZH5rMByunHF6YZ
hgqe9qoQ6eSHDGt/HWBIIGI5uGeAyxXUh5vXf8EnHltMgaB1xmLYvVgg7Jf2GaiE
h5+2BcY/PDEOXKL1Xl7xIaJ97zLNl/Y3hLX+osxQ8dfRNeKmricwRq+mldtMH3Rg
LgwraQiXBWnryztWq8AxDB/3k7tjVvDDsmB/b0ipNoBnhG6bWN9ocaX0GYOtwVYD
+tUEwJg3KdSkYWGSTTI6U/9AbVmKdpJ1w8qZhQqt4HiPP1JWKWQgf4o5hGeO3s+d
KrEw1/a0pt/sdNp/kb9JUR+n4IiVMcUr2WyLoGEOIfk5Z0HxgcUF43FfA8URbZsa
LytopA/e8/KCRma1ZtHdXwb5ie4TR/PFvSX/aUF8KRy91QtkwJ09CZFnRbtAn34z
aBGexF8nTWpICclmYJl5EkdC1EVBcQAeCMaMY9ghxMY+xkexmFFzmcLAkfPIQa89
+gm6mGeCwWhUZtm8ENnim1hvnWxUEdxBg7P6IIZMtPlrk14a6cRawLgB20I/JOaD
i8R2TeGnWCpUESUn5D4ympXfYJ91ZfB9BT7DUYQ7JhwrInYGuVh9CemBLLOpgBTA
6eYMdJxnFzSvl3wKHqQtUWQraFH9jmoVmQlwvOk3kGS57SwND2MpJWPcQNbl9zvc
RgnEbZGXhOcdqPtzSxghZtMSinPkGqnFZZt9mh4KafE8OYJcA7lKOkTlpxel6PHc
7TicUdawFLk9nHDM0dJn41r0E2boZ3esbMf9QBh6Mku1jBbSxULRr2JuWVJRnnRs
/TYTIw7/MCR6ASksGHjBQ1XqnxsrYZF2yETyfM3D+fYe0qCtOxBPW7J7JksiZuH/
w6HaYtvnCOj468zv3wkbZ+hPQ9VNTmZIkQM/znAl087NwlD1P++7alZWbrLcPZnD
M8Si2C3wwAKz/rrTppFzgBZzm0ZTcsgrP85lp8n+pyb43Y2kgSANzwinNKdmi9NL
Fs51w5Dvvhg22CSOI52lXdJxlvyr2MI1z1nPMHn8S6phWHs+VU/fgT8utlCIVSbG
s6ASeTMxy4jcxosjqLQbC1zP59lW4DarTTsbuBJ2iN1KIvqSKZ+pDQxeUWktTum9
/18Zorhiy3fhY54suYE+fYD0k4079RVZ2QSZo6lAkjDBMG7FTtIct5t0ZKiTAYsv
OgZf3XeROhGlKenLqwYXxiwLfn1LwhTIIU34RNs/XZP4Nu1hN9Y7ZHmoRbgmVlkt
qrufGdFOqycAsFxmEqg7X4yb7ZhQ+kuMYu6Is3Jrr3hsfeYLt3IWrRjTgQB0Fazm
Mu8wu6rVptrHjFK9nzbQmnyVn5VV9LtnIhCEdQZQN46EqtvspDbXaeSIPHp1E6ta
SQCVH53PuOfyH7qLxXTqqt/fxZzji+nC77MQbEAU5LTBWJXJsiPayd0rJYpaToeA
hY5Mm05Yw8ir6vkvDkkC/2t7uQrVoMJJS2G1Bc6sArrIbTRi0U3ke8wwEC/GwuOi
ZkFo7Ry2i0MllVBKsY3Fiq7UBn3rho3zjBLH8oMAaR6nexitk7P//DGQlFM7JDjp
g1oLvsZLyEkzCnkN+Rpz5R6ukGoUIsSAmeG1RKjSchhkhdXx5pmgMdV2BvPB1uh1
2AFq9BldlkPhN+CE9aTRllS0PahueCSli+19afKE4iJK61agjOTMsAdbZd76j8Sz
USEN7xapOb6eW2ZcbFai7lKjnP4LBhzBsTqOiFiRC+GuLP+UwgNmY01/JGSuEn6t
bsYoGr1Yjru6apMLUvUmjz5SmG0EKvziUIAa/tS8qBAD1KtC0U7Vj5oWuJxy+qjW
CPJPZtxKqfh3ltgWZdcZh9lnR6yuwnn+JhmF4/xptMumUbcrYvIhslAe9czEeAUG
QHYMIOHzSttRaAwx+Uw7LzxSpDz8uyjjVhSVPMVJE5RM0lLOrS6/auP7OjBOlYc1
7VAJm9OJ2r3b9oNh5DeH9ZGE5qSo8T/bJCGnXp+uH2YetYijWQjImvnF9kO6NhgE
PNoe791WeQGSAsxbGhgfVRwWpnKnoHls8r2Z9q14z1oQ4Gfjk2UqWXz0CPTDpTOH
Vi5gahMdp/okaMjWDxC1Al72kkYb2Cfdf9u9Zu1O3mZ/i4aeQ7Cn6LCSeMocRIWq
35VP/Hk3Vp46vTzPuzPbVnUhH8+cgOtwozr+XYoseEw4PoX2+T9NzpGSthSgYGrs
H8z74elmAH5EX6vBNeZ8nrlqjCDsqZyomNX7xnD0a+4FCsm1xAcSQcT7xWI+6W7o
nVuXsdPbP6YJgMG/lTfCQ4yzx5kk9B14VJHts+6mNvzVogIEBC9UtstXu1o1Qbgv
jqpr8QXNJWNRPo+clPe8yq5Rm8ZXrhlAhO4hb74tqga/b0QC3UdZNXNnLQJgiJQu
sKln1RnL3a0mTdj3UL8Numij+91qwO3TLwvUWuhy82Tg6rbbkD/R89Zi6DLIU2mf
Sh/mWu/Xara/rBhCvp7+dnQyTi+BLIGomVgQ1eiikpBqjpNZpAk9OSmoD7p1/pw0
rJdkpsjZG9BG0/txUg9ax++EPqGRPfK3Ar5+Q+9OqXP0o5eGYlLr5o+JLarPSPtD
LNHkNbLW1+tFUxxjtOEZf9a2733axPSvkHsxbhBQ26fjwF9C6kGFVnpl7SO7U7LL
9zDn4lua0RLHHDn5TcSGbKZ/Z8vQMtJqLsXpQKaDipPsHg0OBCGbq7lbTpKTSpga
M+BtJ3oZHazzGUCoRpoZ6ZulqpGoJvvAt8dt2lH4Zn3YPiJJ87VUiTXVSc02kHp/
aatV6zpfgJ20F+6jNNqA1fZgrfjyGqVK66J6S62vwuvsfYrcewMP9plWB02+H96f
bqE6a8gxoRwPdpkICxIPzjL/MEut9Jdw1l8hHdQ4iKH2Ot9Vac7LEdyu/8I5MigX
t2IIaCMTTtkChKHWYt8xYFRXwQC3oPRh0jCXzDLK0/giQDhzbNCVdKUcNcfyoP4m
/Q7lZ5eSaCJmFYswz27Qf9Hm3Rgu6q2vZm/jUL1aayg5zjzjktJ8okWNTY4xbJ0a
MQcwhMjCEOEpzVxIBoRTVX0qWTBYaTLVc71Y6HRr7+gKT+CLCxf8A8RAEnejfOHs
KJ9P4jeCeEL7KyU5qgMFoWLcSSbu7axNXuhqEth9WE8xqFEiPU3NO0mal9t5r/Er
YuqxmYa59Vsm3c+FUGEbkkiGV4NiL41Lq138NDn0ePomzE6VyqIWstxd/+1Igdvt
hBeFZ/ps30MhOHBOIGkRe0HaKDp2Fc42pn8vRUoPp3++OZeOwmXTj0lkBHyg8D0n
X6a5hHPhYUtbzSTbfAt3m+uh0Y8Q9uPstdZb9tX5kCf3wnPKvwJxqbn6UWolJpGC
qE0slD1GQ1yPtm/bti6zuCSvnZ64r4dR4fAepysufnmSpeaYLcaeZQlq8szFUnkL
IvV/rVunygOVSCJbVkzJX7btFZl+eF7wNKacl8LBGWIex6JNZAPq9wB/JOA1x+p6
FiXxX8jBoJy47qJcQOJjMu6O3j9nFui8XKXB4QJaooiZtgi2C9y0fqWa9H8aiyBM
AQyPQVleM+4bAnLEnjMcDY/H4Y/WiP3kxu5lxouiMn8eMUv2XF9dzE6yeoLxPSE4
vpnJ1V+IBLiBQQmYrBuVEuQJUN0jgU7RffkTnPgn8X+ib+2Sqhxdt4KE15d3Znst
VBwU72Ca3WaXY+AJ+nmCJekyiuYa4/o5LWQLb4eqKMns5IXl3TuRfZvvqKsFXW9M
AKINrNGgkdwNy6+3+NnKD5/gli4Xe/EkYxxCd78Pi/Q=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UHSJBhF2ca3zecl7qwFnEF/HfDJxuYZAmAxh+XsLml0hjoApqtGM+7dCcW+v0nZw
vtIhUQ70AOAiSnV7F8CIIisbA/+VKGg8BZuvmXz4+0qfOla7U90kvciz9+XHGxkr
V+mQTxiy29gSE89TWvhFIe9kPFi/sUuQotGaVZJWgqJdgjeQxoEFDtgLWNp+gfMt
y+e9vS0DgajD6up7Vzn23whCys2Yl1F3KJRtt5bs8M4zea1f7/3fDWbjsG16gqDh
PRdZGXdKTuTeNt0mkD6HO4AdStVwuh10dCXl1HS0JTfzQ3q1KcU5kSsU3RKQxvgp
EEhmL3+38NSsfLk3kMg7sQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
olgf12Fm9QfMaBqCBRarrTHLWM1NfZbAzbsxyuaM4CYPY6dJXg75Dzh6eZ4FvFjd
Ewf8giZMTrD0I2JiXdw79+Q1Ek+Y8If5APESmAoy8ZBDmChPI7kFR5G9kll2+EIl
HDHie1ApI9/qakwNgKGLJPUq2kqh2r/FnMMSGoPkuRYJqgQIozYqZO0X0qTWCurr
EfkJOSq3KBX/N5R2EuzU2IU2wFey6jxnxPnvtHJFNyon0xjuhCAb1h8sDzYuiy/7
fnH2dZKyWIQYCqhBYQh9nOs8F7nEoTEINbVGaxQiK+/6LlMZK2VDLohopnxK6i+P
gEFeREBvN45jNnOSCG7BHJtgQS2eRpF0TtzE6Rc5Eyqq7C4Uq1epIVz0ACyVkKLE
t4N0nGDC8h7lNMlFbIeTqwpGooGOgJt684Q3JkzvgzDL2haEaDDuid39pcLV82tg
igG5mtClShlQ6odOrl2YrREWAj6rBBQlE7vSN1uHBIl+b9LQO8oRztNAHspYKg+/
BJQN53EK4rWcspc+e18r5AgeAnr94DNtrE8szgpWtZAI/8s0SlOsgOMGHIy1+rNY
REFeMSYTweNqDvYUbVLPXO0SSkH4zFw223H9N0EVJ7ixO4rKGXSnA0ixAdGWxmSB
EElwmhMZ17JkgAZffPN+DN9ZUelLGW23BwzsGZMuXYWLoxhdiplpBDp5YVpoHUW3
p1hHDCkO/mQRDwKoK987pyVy5jOlb1a9IURtKz07w/g3I0Y4GmmCVGVwPlFajKHB
Kh1UpRaekrqFtYHTa4Tsz4aRo5XfGC1hixokL9elSAKDmy6sPpCljyQtPFBUAh+r
GPz29/PRq1nepYD2NyrSdQJBsVXrAb7fRDUqLIiXY66mLc1jnsRaMYtuxRYa4C8M
SY3U0ZEPcas2NxI6wpYknXQhonngiUAzEZHTwmgiht9SokjDTjxLlBfrhCwtyfSn
hKxVyxGyCCC4GQRD1cuIU6wxIoOkhY0mr9UIvyCPL0BY0Oc7xUmcYy6iOd+3dUYM
J28U2XFfJ1X/7KjjDsWtcvrIi/XwituE+Ed+jGbNjZ6u2j+BmwykGvKFMvxE9oRW
a0r83ipHKQlXFznb+EDuJwbnWb0u6B0FzTfX6fexhpKQhu914p4npqfqQOwT9dpN
HxpTbbWRttJYbV5uHG1M710lyqapFuENDuIrpwZa9oTxKCZ55igkayrShmx+qs8p
ufqKzy4yKA7UwuWcLNn2H/YyAR8MDC1QRLIYWgToS7KFxOJk0l/HskSsW0C8dohn
3trp1ENaM1mavW+nVcUgHaRU+JsRt6XJx77kseX70sJ1Gkw7MU7+Yg6oHc/FKJWM
1vgZpFauvMjqoAz6zHZ/hl2OwCs47G6oTOY24/WDmO7hrqZIkRG8Du/G0JzVLLVH
Hbf2cw4dK8JER8Nfwax/0lHTh4Zecf9RKIgJVNs1q9JHC8IcMDNseipvBOmnIjpT
eIobvLxqP8w/xoxk5QHFhxZqRYSByevqpfyU/IrEAziuvqK3V/R6hPkge2pje5z7
k/HLskMOuWoDuuui2CRfyjjZ7RQX91fxsumpPjnuVFB6jGIWKwG9OQIcKpsz/8x6
fAtE+rzE0SwO2FuFn5mBzCKZkNTkMlswPtuTwoVJ8b4LqOeaRuTibCkbGt4g3KF8
9mnuzTlpzGzysReADxC8O9hhcx9vbrWHDtJRUkSdCzQ1MDPr6RiwWlChJyb+SVmG
n7VUThPKR3DzJ5cOPQ+X+TKbXT4zRmxq9PJLWq1CWfDEgD/sgV/5O4x6dpE2G398
txocAUTLcLmhgTN4MSh88GEQ1aRM9tch6weyjkLHxqyIXSrB6tql9omN4sqmrigk
6LOMPZgEQXRvWpY8zf/BFUVV1e+EDe9WlrzAvfd/arj/8PaAulqhgbs6+ZUIFYS0
9xSLD2JI6mxJmblHLR6mC78z7JboC2KHbkDvNBkTCR5vH1CicjZqFna+urQ5hA/6
4+stnoHltMLe0ivcRKtflNd3JafyDQPsR6HAUaDYJt9AKheIyPZSZdWQdVI/qDkK
B9h78+wxPC2FlTsplm1h4GZqirU9Lrb1qhoG8yBlzP5Hhozsj8eHUTywyyRuPPsX
5sgFQr0CAA1096X3JEqgddFyt5QwYahX1mSOqGDU27WasibN2l95n2f3mnp/N3Ow
7P07wCbVjN6L6RM8hsVwJsw2e/8mDFj+tz88IPNUf/EMCfbsXGgpmWrK1Gg8woCM
6xxgpcFc7YfLPtEc35LwkNnmvnQseL/Qoj5HuRVBUmxfRmifDChsZ6EKzHo8zMOI
4PqVu1v8LERbQs6tIoci8IdrOpzxtrDaHAXrF8y/NJxuBQ7DdxTBApGOpUXf5hKP
DRzXOR8jumQksA+Lq2rxrRQUsTvAWbx5DRmV5SnkGSZKXXHYT7u1lbLt6qjGd/Mr
IEBuAyO8IuPuZHJGv9GeVxNk5ayyP/lEadd8kBNZvY7U8Kt5BzO/uZQFWhHwaUXT
AKYZM+gr5QDjnAIe1C2Hf37TtE4jogNJGgMru0k0cs62J0SwhDlDltak5dQ5ylT1
rjbg0mxLTpXxwcYXOFu3iDzI27GjBmKLf6DKfIXF8f22n0C78u/E2zbEK7qf68/F
xNmR0yXZOxLSwnTliRQjxeLuXbG2iUIapoF6nop/nabdlQFxU+soeAeHpFrn0DXb
01kMT/LxrX0yqothwo7/0mG4EMQV6jKp9WOsKhUNAxRsbBsWDgHYldGQslrc3in/
6rHPEt1Errc/JrTG/Sw10eWYg35gXxgx7WVXBk+YYclJBp2bRqIFR5g3HiAg3NPh
fL8yTE7OIJ/MqoexqT1q6N1XrpLPnkWl7sXMYXuQyFCAwcRsgeyIfc5WSla3gsJ3
OnUOvuruKyqLkClf9O7RYtr6kCnxi3Vxpvu+9jUa50lYXyDukP8uJSSd4RLKayhv
NRIBZaoDHr7S/yuHddgBAd2AxDNtpJMEJi46hEkiwU2Dx48BgwFE5pxobBp47cGM
l+N9nhf3EKOoMYLCEs0/0l0BGSylOxRrajWRVvstJKqVITnHDHMHq0Qm3VaDXe79
FJupnf8KdCKs8LLFzZfkg18CgwZ0o/fRf2siKY//IMXcEhTSFdIbxJMbmV+J+h9l
E85KatRppvCBBTrwxWJ9fgmRRWF+DbXuBXitrpGXxrfhxib71cFBZ7p2bV65DsrH
ocIWWbw7ZvySzjZUjJZYuggVwr3VTIOgUNyeeS/yjzQ89DdlNzrJyAHLf6O79NLJ
nDYYz8ZaPgoAbDgZ3mZ/10UoZJ9zi89cUEGytKhkV+5s+xGujAVTRv/PsPl/3PDN
h7tBjnT3hLlWPLi+3M7h/UZL5/Q4l5KgGBBzpX8XbxXdpOxijq0RiTZzF/ut1N7a
q7Ojnv4k+WztKrpL1pq6BTswNRXH4cdvtHjx2FJ5JI8etnZ/Oi7AOILSpPgb7Sgh
rYSE7JlzLV8VMAuvESUgnkx2GlVfOWGjLR38RhU1RVGJHc0TzNyk9A3B9CL71ytL
EhYi/Dr4uPBT9Ju55iuUtU0ycX15SBF+di8duRnY//05ARTtjWxcxkSx8fVkzQez
JA758dntBeY+0fSF+BWPPPPJ3W1619O+KEcWswO/LHQThret0nG9qp5QpvrJW3EY
hNS/fUKSG+pMbwC+ysIQYryNDzTyY4eowbFDO83DGrQTsua9BSWeqCz03uclIj3O
IJPCW3/eZCE2A6e7VjTuk/m6Hcj1yv4UHSVbOQSwKAE291HpyW0wTHJwOz4mGtwi
+nvq4ZjU6hGo9daotLcLeqxUKrKWATQyasFhOPYVeazmz7cwsDkXKPjhcBeGHJMz
UYGnDTVqFA6NwzGqLMDyZrW06KtdAu2YRdGjoxnQu+bUJcVO+Qo799aCrB4hZS67
ZlxdAd0IA2b0Y127BQV/wJvr19WkYUOM8h2lAHeRBft1T9atm89KdwGlXslPYe30
SGoQD9qjbAmeO1rhca6WFmdinPlSrL0XAks/VDtJ8M0X8n9bsCfL/wvmv/Jriixh
01I8Yxeb/VK4hNHPUubtmNLikAWscepVdTn8v2HyTMD4EMohVf8eQSpZVi5tl+a0
2Cq7oBmc6MxCnDd4ARl/xdXueka5OAaU1HSIpzh+qolnz+j+2fOJgts4x0jp/DU8
NrFMi5lmmTQIePHHZqySZTO6gzSZ71oPpEFrkBhVNwrhLS51DZIzgeg0DHsWpnMu
529pF+UYgZ/82TL6AItn5ROQz1ljx96WnvHBttFLA4+9Ibb6bOOWy7Wc4kOWRMHR
XD5HeY6ugVRTyOAfsF845HhcJBOH2fsxwZVG2fPI+JX5e7n2+OE2jtE8tARlAUsQ
3c+cUsErbxmrr8nYpEVyYLYzyWgvGZbLCVloSeLAsBRNeyN6R7qnaY7yKLa1A96z
dyLu4Li3GYyaGLJ9udaHjk7caEi+VFYhfzzXgk4uBO0itnIjoyAWUjp4St2/Wbph
0PCDBbTDSsnx7ztxcWB46RlMhE1GWHtm0rS8reay7C1l/ooOfGUGxZ7yuZLWPeok
IUKoJiuNUoLnqXfZ0K19goQfzWZXTjirMfzg9ce2TnJestlD4kOKw2lQ0nXrEBe7
xMvlffPnrJnX9BaGE45FhBEX6g7g2MfFqBMG4iUAgtWAH+1qtYM1EzF3qdpY9k5Y
c5bUY81Qv+f48zGZ/MsWsy4TWM21698wnq7/IPpvmXdnn+9Dcq9oE3GE/6wuD3Si
CGK3umVfcxDbd7SjWujvH0ylp0zsbcTxvRN8433dwenTsFmKpBEac2JQwWMyFj5X
g5BDaCOS65qJZ8lybBPxjqYE/PwagLTrIcDD+H9My2HrnxUDEpKXt+Kp36twy/Rz
pwPIUoaoxuzgeMxg3303Et8/ZtoINfKJVVqe4YPQ+ok6xm5J9TBxnfrGG/g/MZJA
pVPvRyLSrikp7ZuVpPzu6sMjnqaFMvdpJ3/tQ+y49PotUZm/22qU4sPr7QyhGPnN
IKQvebXRPV3C7V5dEjgAKVq12eBNrfs1cgKTieX6TW71TvcTzq8tmZebPmeA0I0i
4bx03fFp9LpU0c4oEQdH6MiEZhMAWitmO++qlpecLMaJYyb5eYrXCgqi7wBsZyRM
s6a0q181kP/yRj6O0hb4tms1C8xrS9g/D+FaITAQjRQCHg7QEfhlVukdnbHUUQL6
TRDfIS+zJHsDTpqzM5lk2V5/kckI0IrAb8JGSQktcoGgZj+cOn1FTYXXkQF2pkvI
wa4cwl/KsMqjDzku4yrK4rpoLDnyKrV+83j0K5ZXvfzmCzO/w+Z0JJiY9tCrls2X
A7ecdwBRx9vILOGvGHdlE49z+RDUPd6tj3d0+HLNPKXy43CSLPPk+81qp9JWuP/u
64ZLdMkGQPcQUb6dxGeVa/wGR5thJkGlEmFVUkbK8BIKTwVkUWIcJsoZbYS8nA7r
SMtdJ15w5y0qPv0K+HmkCOYqJldvzwgwxFntM5CZ6ETnS3Yw+kepD0MlSlsTpIQD
Bi8R/uSgrayaWHN1xRFAZSA5OqJnTsfh448gjf80S8BzGBkrhqcuafshSGAZlvkz
abFtipkzsNZjNcQ594fKofa4txwSPZQ8wKNDfLYFOhANR7qMWi/bu8whoyNUO75c
mVnhVhqeZ61frCh76+ZFWS+r6PItBoTluhUkUJ6BCQVa5/JP4ZkbnyE+KY/vm4mh
ZxfHtUmkL7PI+vCNEqEbJQkPQLsSYMAZHbKJmklYF/euGYlKkQRFIrt/9/iQ438+
e5GpX1USvmmBk6gu8GCqTdWdqCIhAfz5VR3GHQdwmVSlGDYXAeyl7QPjGO8d2pcD
++VcbLrxkiv3ttEoo718ObxeyoELgqlJoiuyNhiWtAmsC96Fe06/bZdPDalWfN7y
Kr/cg06IpmO38yUDtMxkFEIKTj2ub3au4GIIIdUOewaYGVOCZiyKG8ENBQ2CacvI
MtTi2VfRsTyTa6sB0WMHrzM7xovF7RPkF1RoGaTJTfkVKLYhvY3v13GgJkBpoXcu
MdaUc8ysGg2J9qIJF+BDfNyo2Gb4HLzOkWdDziel/iN1jkXrvg/MDZJRQ0v8L33X
789jo5q0FF79heUVDDcFI8UK5R9mwaCyBkzPRYvEpCpMylknUzrqOmAqB+PviIG5
i+H12/mDE4DTN9/PZNfNdMyt3COA/amoJxXHmfeF68fNe+Ya0/SadbOrWQPRjC7M
4V5Zm3FdEnQ2ODlZsBt69J2lgw4dPNpaVaWyCzn/FYMefq0cyZ8KLtFlWxqMQkce
ZmQnmghnWVq3BkDdV5M5IKZ2eZzKsQU7kQrXJIpk2iYOh/d8SvC7G8mjcbW5lvSj
Zs0qg5A8rSb/E6/RZlMbHWiG9z8vixoRO2ByEA1jQbFNZFJAJgeAYYVECU3DSWiD
Lg7/B67/l0TOdwFWuHNY4N+xxG2/sKTfmFS1MfHjvfwQ44WwlsldHe2r/kSBmI5S
nNrnc07jBMQkidvYTVkpIn0rT5n0iOf9c/EaEATugpZ4IFWZUO37klHnsWgeAbV6
0j9kb+ScwjaNsZr5oh/q9GGX1JTBsMhrpARRUcBxre6lDoTVcMRJUda96h84pK1x
/zLhNpNz9dmm8P3COuGTEPn5aqPecLewE1B/ea1QmSSJvNlwvvxoyrHbRuFb0JBZ
wUx+vfo36GyJFMxIzMLeRzGjqAufacyH0AhCTkVfAuHfZt5pnCNAmVwNUWHu9Tiv
dwuMsOlzq4M4Rj6X7xe7oRMMDnmvqNZbDfQw2tlsvZBCskW/uNrc9D8i5Y+geB10
qm/V2Nyd6MmCxWDcg4oAGbiBK+Pf+DqULVOOw2lnxLyOg+NNsENNMv/YfztiYCh5
g//2cSxuniFKHPjfYKTalvJedMTHJ6h4GdrKk/udwLC291smC80AOQPfg2DCHdd6
Ymd9KdA2Ah54xJx+eRJsPWImu2cPR2u7fkpw6HVqkqRlVBtLyTjFP9QwbJNBUZy0
P6M2QkOEJR94yhgCFeOOzbqliVbUEME+zMPoIRZg0l2Q7MSKPd4PX3nyKjfw/sJk
m54PrwMvo5kOvgfon3NkX2nOD2lucojdqcGLtVuAufpZ5aVroShYGUL4xQPg301v
0YtrWJ/4PpFPUuRkVdt9AyC22Mu9EOIhHleTjPmX67gHuHfXdi1JDc4TJyxZXVig
MvxOWbFeEC5UXW7Y4Fml+dyjsXpxkGvEJRnDHQrXkPFvIeaZ59L4BXAi2MnOB7mB
tWi24S9g4HGNAJgSqF++BNocd8bvudPeInZmbJtIF7bi4YOtiPDCpzcK1oG5xxrP
znVjC9PhJ2qi6J8c3XAUMsC/GDkJEk5dpZzZLZyu+YFAM+8TI0l3dXYqJEjCoKwN
5yCzxC3hVU3mkcNJ6vK7G/x0KHBs7aCNgH+xRxYR0Q3HjHyXGZkbxwR+dRlAgjjk
zyGlbG8zPw3HeWOSTrfnCYLsFRmVjPoNufBNczgkZclRIGX2zWt0nE17H0HWHWtg
GiHOMDkr3hfCBbcZ7MjAukA/tmHECUJMc3wkdoG4FraO5M8zdFlp0p6FN7F9cL2t
sOKgd3lbwblJmUfl2IpHMHYAq5rnlOwbd+wVhcH2IfheH39+o4MHwW01hPjf785F
pElKB4dD7v9Xe5bUkbKoQ6I0acm4OiFj+OXa0W1W7AlBsZfMns4e6T4UuELlmGd4
HVjxh7x7VVBFkexPBJP+F2mGo/9FfTi7V1GIegRoSTMfTYtSR3I+ZO+8C8o9bCA5
KWN6BvbNw1+1bnR0IUYhFfZF3VuV70VL/oCQ2Qt2lHg95AbJ/zA1MzKuMhFS66ll
Jsu0Ax2xAjQbXcLGx6oVBBfqF6x5vy9As8LzeEbTsTUDLfJfe43k6ZzufgMKKL4N
nw62/Z1/k1af6pZswk/T8zxxHhCobHTyrJFA/72yjcf0G/9WFSV7gNLb5boVPz3l
dCIle64/4f9p/A48aUXHfUJuyvCKtlMEVpxoEPKkfiUQThgqRBv8QuBoC1zyUike
z+iSUCOr9+LgHyMZYOefGkkW7TS6SQSLFENpARrC7ymyT4y57wvbFrBNdE17GbhZ
GeNfK3BgyrwYQH9HMQ0pQg0VB2eT96ZPNWgplxWBB4+8vOR10eJ2Wmpu3cQXkHzo
JNlJq+TsD2nzHeO6XVhy5KrowgXXncQnFUKUn4lfAeZjvZ2xDEDc76pCMODYUOUa
uS1rqORcFvpvt/awUmB2P1Sy6zpuTx8dnY4/M5UDU7N2k5K5f1jpWy0c+jxVINmk
Sd6QQfa3jZD/5E4PdqD3xZsoYY2jbsShMAxnHLQ1Zz3lPafcJWI4hoBERptUsdhl
MNFwRWGCnCuziGN7TG/CvsRQBCSwMVYLrCyBTgkQLyb2uMN8rbPIKJUmVWrGEv1j
2dJDlb+eSj+0KLE7BvxggA6YRWUOL8YoPNTCMSr650txpAxakcUXDUcW2P76JjsX
lLrDKL1aBoNpKn0+FP2Q/9Bb6WgCtOimuQN9S6dzuuBA1q4BhIE4bW1lsjG4EqiV
XuxOBu8aAjKAUJxowZwQ6xizWg8Wb4OQfP4e5GxcNCoYnsmppzmvH3GjgS2Wd/ub
tUNeJ+yOLsNmpTMA7r3GqKPne1u2JNIvfDxvRrnx9lqDAkMuB+RItnddnyZDE02d
xpEzzzcxJIptKyx+9PQSfEcG86ak1+Z3mh6cV/Hly6xdFmVCr+KDXPhOrT8eOoNj
9HT16JId4l+QKNu9B7ziV8oKJECGRSI0/JeRmFZhYlz5UPgln7E1gwEzYS6BRZ/r
qvfVPLYQq/yCHQDbggLYDZ5cbMmsIS2y7NPtUGDmFzVcQGkoJ1ZXSShIJmEOag56
qB582gPmXUdOGnmsJY3Dl9D9sAdY5KEbyHs8mhEVwurtUJ7Xq8c9bnuIF3R94J7K
YHVlDQS1EPcCrVAeSudGr3PWAEZV2iR6S6Cqd8IKxwhgB1LavbGPnVMAF1OUmXo7
KOirxmcWMf09Hs4E1C7Mwyem97UUcw6Ta81VYWOmILEMFfJL0Vjp9uUWwUw2UXK4
c3ShwSpXLy32TL4js2i05Nn+0YV1+Z0bUYzGwaWHcEInzBFfefdb9tZMXvw40ofK
apEil+nOJyzAro+GZ/AbBWljAArnlyhtt0F6tBH5rgiOiC7MFvu5vfVz2UJaYwwm
wA8VoiqAqxBWy8+1fw+iPylmH0ZLv20WeeOXvQn/itiYWgFRuk27s6s822Y/RtWw
WU0kImk79SCQKY04FW6zooNKA51a5waTmbSe9Ar6yFluq5jBiTcKIds+G2i18WL5
lH0hAFMGKrfnY8eCltNXfW543QqkRv1BZ4/rNl/sY2WK5irwlfxbSOolPpI3OAK+
4h4gUdAuxolVymaoIBFjJicZc412HdS1cyarevBrWvky24PFPJqLAvgXpOYPIscJ
dRuoPh1m9uU5nkWzzDSvpZPubL4OyXQRR7FjfxmS3DPTgrPJaf57+SmXwMdt4AAN
RW2gHKqISIU6gDLjlOVpC//ovote2fdsbOqxBQCHLJLab/TbsMfUbUNWNhUa+te9
18ddofuwraOsnUbrR1vBHsj/lpXhIPRRkXNNfjp/dSDsHu3YIS0FYy6CvFC0dTiX
1zYmPMRzDFx4D/Cbdw4CkDqQ5fkgSrR7ZDAzUFQq0EFFEarc7FqoYQ9Hmv8wB4k1
yPA46cE5JJdfVGR5IPWmVlap4jeHQsegBiz12iKiXlrjl14EnfJ+yadCdF91xBjg
iQKzKThIFVyNq/gcrTMmFaIWrX/SF/TPAxKJ0PRqXr9uRyzRigPJmB32Spo43WAN
c+WmggLuvBvVyRYmt6K4uQ6h2mVuOJ5I9rY2+33fS0VKLmJMTpVN2z2nWLbanEns
oRHKy16pVwhcC0lvkCFdajt5q1so/sYehDCfiawkWBQKcRUsY1zuBtloKqLNZGiW
mML9AxyQts8ikUEunohgOM3bcbIPYffMVhTnXh5aP5RvX/F/n6iJq1vnNEg//FFz
49ZccPkgMzRs78VwKaP5ds4Xr1YjLuKHQlv/NIicOzoQ54vo2pWuOIi7Q5MrrvmN
2hcasVvkorDzwH3c6GsoaoQsNxpwjwPGxLSzbADjrICDkAZa1l+WiaAKI96ezrgF
RtiQSy78CbwrMtmD8gCS75RlmVZ9HL0hudmfNrlpinW4kpLlmwFAiePMABGosmlC
CVNXIsCmdkTOixWb6SAoziSDHRyHN1MondPaOe6Otqrsc3yYBw/lbOK2/i5ZSe3i
9D8ewhrB68Br/hECTDusx2geM6v7KzTd7t5qzUyZ36nj76P8Y26adgyOd8MkRSWX
/TbC79ZMxHGq8t2aU6MA4NQE1GkMpDWqZbptyonK4FRp/PXHw9q6583cWClW4V6V
bYEtVb2XKgX0hGGecKRHPmF7GVClD00vf3vqjBj8evjywhQIM0j7/TV3rpMOG2iy
3aB2oQvAwzYg+Q7/qukVuDrEib980eoK5+lmwWohatTDU8n30mwUBoajbdmFaF9B
xr1aq68haLza8eGghL9Fl6k8/rmhp13A5jpxwXrNRlevaQXzBFwi1o8dhktBhseA
ZFlf6b85bjD3mQ8vsx8kQoF7hnduwp/P0rSVHdrnj764thdHSD6IkHnTtIGz4D4Y
J91FCRnAuL2UGrJYDxhC5jDIjHAlX6d51T54kFadR7JRSCo07WMOFUieesjJ8kj2
V0/FJA1rwDDmx+t4Czbzd6IQJMbe6g55ILd2eI45nK+szyYjlkDgDQp/grsCAVR+
wKa6MJYsuw6SCcTroI50RaAlfurN6fRWXQ934SRGwXULQLV3qda0TPzJZwm6MPI5
d69h8nYTLI5RR/MrkivVwnF/LcjKBtIeaoO5ZEtPNcQN/rL+TljCnsezp6sB9Vqr
ej95lwNaRzm3xr19skYNj0Am0EF1JjbC3hmBncm9J6Sow/k2Rv1IHfkO5JTFQqm9
8LsCHNezHCUuoNTPAIboFfSPeiG+aJlA+G8mXQWgCP2VtdaJ3RMxDus80ELlnvJr
IEnNjWy2mVEIe8a327CmMmTBjO3KYDPLuyi+GeqeBuGzGPp3SMzvBidzhpc5xCMu
jRsC7Axrwj+fefoZFVkXNPNOvEcEXSHgyT3N4+zOTvMpvn3HnM7bi3nBr7EnS94A
7U8Su8v5ex83xUhPCjbbtA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WaQNC4huU9b23Y00bGsVFd0HVW5JIm/eFli21Rt4ar8VZ/SGd3VlOAXXgD8PtOlR
6qZ0YxdKwP1XtkVEeaC5lpVxrfbfX94Y7NFh82s8spNB+AJTPiafZ+3LGzOFDkxR
C73CYfyETohCJohToPm6jJhcdhYp3scDKgAFXq1ghQW5/0sUaz9y9oXc2XOtCPMM
qqEjqXojow6+TbjhCeXog3rykDw5+Lg0b23LfSnfto27G3Cm2mjJFZ7kF3WhE/cx
aOLIa5gaALrEg98FnWdPcQiMzuK/f3U15xdKMPQkSwKg32kaIWl9GpqXnAIMj2Rw
DorUNpHE5d69iae+yS3TjA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11952 )
`pragma protect data_block
G6E6G7eWg8ePBHdyxqJLShjOf6vbDlk4KP7CjkFmuUszzG/wlnpeGqYBEFKJRiPz
zb/KoMbBVJtUPGfB+xVx6mWsBM57mRFNDS7axGfUGyDJkV2bZnRgJD7Nuz1bKv45
e6PuX8Sr9m7enQWjMQXxfRMcjx/6TrZRMff4efzVy8iXbdX4b2ZxuOi/Sg7gXha4
ctVAvkrkVl+wA1Z2YtvCmzz/MbYhvOfmE9jPPn730yqyLOtt2T3ZGyllKaW2lMgX
V5h1FHqGzVla8fjPIiAM1l6tuiwTLjl4YkQGTjeOieCNSDmlRbYhrbAEPJndu1eU
YSmvkiNMML4+fVZ12qxyFTHbRTTwqK3my1ZowfWM1zSD3feWj477XhWQnAaW0kc1
/qrtWDXRjI5N3EzBL6zViw5C55HNfo9wVSfr0EWWHwqbWUfl66/UrDr2cBRGx93E
q/JbHd4Es3FMn7Uxe4b8ta7wrqxfytyeBKLdIrGjYzjYkchXf1unaLaqDS1Nierf
a0WbCZhnT0Nux9yZuYztIWOZ7ffzl14adeHcregDoe3j2Mr1RoDt+z+r6jyGnrtl
SBJuoC5S5w1cOqDA8iHSCsWPTrLG/JIA+70bruUcIDxK4ODurqc7Er8M0BqeoU2e
WBwnd0JdK7VU812Kcyj4BgcqVLu7lVtOz09P9i8AC/Jhj69uIJOys6fTz80lviMI
pIAXNWMC3eR11Knp8YM/g2OOmX43uYWVR9Z2Q5yhqIzGMAPvXCEIk0CYkUvTEjaJ
PmhnPNSHSXbTItyr8FvS8BIWYAf1XdG4erYMlbSu0G/pZ1nAOqecIV+C0hzsWVHp
EDS5VdV3AMGCdyYWm+oIcBsXh3x6rD9wS8M8HTxwxf/NkCGa6LGGun864ln6U8z/
foYeMW5Sej8ALmX9DRkMkOQHT2GCzOtDxS63MiVESa+h15peSPyMRDfGRPLrAGB3
rNNScHiclDxaF6YlO42o5hVMkQXBTWj2R0lb6LMhtq3+CtNTbhuuEVO7MNRa/lcB
5rGY/x6JFKG6SAbeopJrYURc8tn5wA1SJkl+fthB+vrJINNiBzWeKWvgOa8qwRcm
w2JbmxhQDEsJCzk/omp/6xRNOZegjilsFz4YpSatdTqgiNckFs1+DhSUjarciWfN
uW+TxpXAWwTRkS/tmbDJfiHguqA1TJEE0+19yIhdOGAmsFpmoYcEKVKHyvvbontM
dbOdh+MXsYDSCNTbYm1oLtLzrnysjr77ZOFkvIk9b3DZHtSgYayJdXfQ5Dpxasll
6OS15D4i7ZBKLTn3VMwtgEwfHtaI5vWBLpfrPQWAD4Yfu2qTtqF6JLjU2ytcytGL
7HLbOuD6ZT5m99hz1ZXCPkgfLeLKq9tNf4Lzykn3lnJfacU+ImSNbEFgZHes9Upd
PvCkr8LoB/q5JUWM7del/2fQZMFvtJRwU02TWO96nNKu+P00ZBpNSfl+PYp7dACy
i//++ZCEjU2LvgmIJdDwc7zTYq3XAIsDkF5IU2sQL95aRdvo/X+4EvlNNDSuelHf
Sv9D+sB4N9oDj393LQJc8LrAY/0Ve2WutZkcYmjgqE9yIsH1dY+XIL9eqF8BJGow
DdusOQYcwEKjODbB1gvLqq8S9giQHtLUui3tpWyo3IZJpdkGDddG/z6NFr1Uy/QG
lznOusobSeOI6T3e7eXhHv1pDCf2oGBBMH5XWcJfPY+VtAtluy6p0oe9OEh5oh8u
fdzhCyitRTwRCZmy8WHkk3RXHwxI7e0X1RnisxTS02xUu+D5PH8RlYlL7+foT9dR
P2+ZaVnkaZESMyzQQB+7J6+6YHYs8QB/6A6OFrQYCFRLHDXSAbYSETy8BAJ5mz5a
k+MvcPwSenuLEiy+p8S6T+myZP9ZiL+A7cYKnM3uxWQk2MMhiFXol7XAdmRsC9/+
gp27TOQ46t7JRP8ZbYqacPOvxpp5Q9JawfmE0WL5/UysIHeWw64TEkuS/AjOixIK
C8dQUUZ8NPUpWk0eUokHB2emPa760B88PR984whZiSAXZUki6Fagd6cTIt0TPAx1
dtDJh/aZ87F6XXmLADw+bznbjbPo29VeodQS7VW8XY4RuPLy3JJsLHW3V7x370Ro
QItWzEL30jtmcOVMsko1jTpzmAgDcAlcY5fTB7T7c1/7XBUfBN4qXNPt+96W3dyJ
DGTUVBwvlo4bRsKj9aiJXyeYzkaM6vgZ7XbICJ9Wg/nv6TE25HGHvyMxehWUJktd
A0W+FnQV6P+Cjlp+oKvnABWHCTqRn8aQ8Bi5VkKYECqvfvySBc0bZfSA5weYK+dl
F/l22sR0bdSJRj8IHnHQvZikyMtEHBRckIYzdUdDx58T1j5zn6sWTIKZQhb3xVbH
p+hNypTw/CTYFPRrhfruA3WzOg+RpaK4rkOZFK0jGuxXvd8s0g/v/+sUjq6FklTv
Vqm3Ao//xtCYGCGV2NLn6Nnj/QEciGAr4LuxHC21WvAkVkmENasQSngolayh/nj+
j0GaZ10qq/9AFuatbyJ607ZX9wihsU4DBqs9DkMZEKtCsF7wd33yd8xKPAiGQ3Eo
vhgvnSaqYFhwknKAdMy/AEMCcoJkK3YVjU5Nk/UnzYmx4o2i3YEHDhk1XBSLnIEk
P67bqVL7Q+aO6MHmeFoX2JPuazuxG19U0d2at5790Cn5ZgLeW6zrN0LN3BOVLfiX
VZaifxeM2R8OxUVCfQfdjPIiXlPo0AmGUw7s3jtSlPvPlXYOrBCIFtBHUkUxj6Et
L4J4/8lgKKtrraARJi0i1py5aKi8KkU2jx55n41tpFJZ/Nel4COtfdqPfEmHsGzr
4qbXpEkQ7hz2rDjhkIT7G/MEmEddMuMGO/md+xvjumV0SsiEHpytGiW1/66fXjS7
YlKHk+0A2qiu5SldoHBQtELx/9T5U9aCT3B1z+ToRxNPlCVm/F71zr9fAtRuZqNu
9wl92P8BSIBykraHJ2tcTO+KfQpeSwhCiiuf2gngoJh5WFNv1hIZVJ5fHaew24Zh
E1x8uiu7iiYLSqlUzxfLxSwuprUjnBWXkcn2dvEIniG6m43JGUO7gzO+ed4F7SrO
DiiodfJ7psrohT7MGhIMRDPQzq/ZXC5bnroiRQeuLbtNLeJ3ZBgv0MmuN1DDC+wq
1alShhUMP3DIRBIQQAKLrrru+Y3qICvn0ZwKztNxBxcpIJxtTyMfxrKCuTb29hLg
eZiOqTWOz/Oj6e8Lrvqw58iP56tv9te9icKN1iHHTXri9CfJwROWJC7RpKPZ5/X9
ygY88vet1JzBQscaRN2/gCDZvS911JAAKmTYQk+RGWuhatO589IJkusMIxDHNTwj
PcmcTXyaUWVsTr2m/BalsWiFw5O4qpyxhOT4budY//Ky52yuFlgOw5obrDsM2B6q
V1Mta1BmFEhtYIAKDq2o90iZOpnopnFyHh5mWstumuk7AJ3z9OyLBFMKRXEpj5ho
9HRaOGlgo5EE/YDkOvL3fye4+W4IOnMQR9HhnAF5FY/NMvN7/nnYA9AaUXGs71px
/pVBkeUZY6LSBZEzbx1rTNV/aqxtEyGL25iJXaJ34PxscxIW2szSt8oj7toesVpJ
TJ/duEWoDhgtUY2kQUX2eq5MU0kHJescikV9W4FG/vFwDRNaIuL39GLwBeDiLwD+
xlW5WDCp/1fM+Ra8dVx4fC6OEuQ0MUdQJyNaTA9IuD/i4n2fIP7MTXFFPZVh/wah
Yg7sioYUj8gS6cZzxnONOJqRHb0klqsT9uBqNP/mXWGLkbZR+tmfqqJksYnqZjTv
z1ugYso+0xK3xqr3fpEC4jHBxrHZTHfin/rKNBgcMUHK4BbRO7vnbGxpS+iPW84M
q+9LGXhBWNB3DVo7ZKBnbmPhi7lCBfkjkpp9UFnUdO9g7KpvPHnokUrGij302TZ0
gjJKuuhwPCplEGp0+3DbTb7kQyHAg3aXsnW48AaBF7k2oaeWG/DqWrsejCKHwzIc
dP/gkF5oZpoorElFmF73NmiTzomL6i0+qgED9aUyUv0GMw3EBOyvJgqH9HXImuaM
wS/y5NtmgpZ42ND389OupP7AyKQhL5OM8txBbS67sMzSG1KrvnxRIEeDSokIDwSo
DDn5BjwYLu6//h0YbxYm8Ez9RQRUPXUqpmN5zrE4eChMqzjexuxRmUBNx4B5DRGi
Hgvp2dstc/ktgUAUL5fhA13/sS2hQKAPTh5HnFf1snoqyv+SkTWm2WfHaoqA2272
n9BTBQwjFQv0Tuz2LTFgKAk1Es2kiBlZBA57XnQbuIvh4AD0E/dbRShXpN5zqmtI
q35/DdDJ3M3roOlHlFV4wN0M7zUtQPZLYY++fJjoNhBXb12hKOR4psxYaqF00ZOW
LMZbQ+Z/0K7N73EIbsvx9z8oqqb1x75LyGM244oRc+9dznsd4pUSuOw/Nt0DWpQ/
IahQg8MOcX/8gqAf3ADgPF5oR2vhvVBGGngpYYiVohx8CeeZrR6kSDL0NboF2itV
bHH9nrMWmGvFhP/8q4I3X3a7t7YGibBCwztH3Sgbxc31D2nFX3iG4K6BbS5CE7en
vn6ikJyfox24B+Jctwcz8X5tqNMb01gcFsRoOqHqvYYACCSnT+mcXZXSd1ZAZ2Gg
TlSDfmrBsM7DsUKk16uqb+tfohjCebFKhlHXb7YXK9rCJkBxWKD7uXATk3C9ARG6
JEZ+zHARxpt8zYrKoGjmKt7A+y2c08HA0IkGHBVsiz2AfvaGf8upX2KExjTn1Q3K
HPsybzwqiczwHMOFZEDDHGBQlW8WLbiAkGZgeUJSbl7phCRy1CAoNxqfK21bEmOg
LOZrNrckBGB8jOBcVAODUK00wxDDnVqB2+ANQPifeVQ6MFo6WpAGYWnmhgHP2UhV
STfGweLbn1PZeIUMLBaKCiFOTBAsU4l2bST3toRGfsPEUC7dB2CiO4qE7+hes7+8
ffSjdSacFbMwl3tNDX61+2mfGez+vRsC20Hp96QnlbzD3TfabCowCaxGwNVAc8cO
N3ToVJNXp0zzQ4dMhXuQdrllniFFY/0yLwas4bl4eznYr9M4eCptqDl6zr+KjSON
6tPzaUX0Jp/11mnijwCgmgZafYz+IX5oF71Gt7a5gu6E3rJBeLGA/tSEarWXl8Wj
3JG4CNqtvAIIM6BY94Mhs0sE/o58KMdvwqvi3OnbZfXhDaVzyRZiDnWJvIgWDWMD
MHSlfszrYSHJIogOtWsJG/g8mF9Uj48IfbBmi/nvZOdrQMXsQxSmNXGVEuXucZdX
NkepYF0ADtxOkYYP4kSGIEwBU10rr57wHbEpcDx4DeQ/PY3xOqPrBEs86PBbgRid
iSvllFVxZBpGELWpNWQzeyBYrTBAIdcZNHtwXAwTx4SL++T1l2KR6fLtHMnBTyjC
p9iJgnb+mAEarPBd1ukA282gTXa7VDfDbmSZj54yVKnZ86vIiPTWqVBFMx6nIpQm
Mb/nL0pEUUe+IbfFXamagkzlsiOdqIjlI2q8GLe/0kkCPT60zEp/p8JK7l0AUtCN
npKBUdF4QWg/nbO6hQz64svRQ9+bUaMWy13Se7A8pkDJ93O+nWR4+TOOnXoq6nP3
D0+yrlU1a83/d9DgYEJctdSWAcQDFxvigMooeeDCSa345hTu/X5fCdIdaBi35vyf
gEN5fQZKeFtvbXFOZck7P0NHVXbJRRVz+BategLqaRcYbgZfNvFdNdxLntQ023qY
ETKQAARtg4tIM5L2KIdCsGL0T08G7q9//OkJ9N2kwOPXUM0ZyGx0YLaGVK4ThHno
TY6ROq+RpfTrIVQQ1B7Tyeq0CG7MERoVwN5/+cIuAEuYSWIVMNgzdaCwI+P0mOMX
B2FG9PVbkF8QI2pWG8RwzGmANVX6X8qLcslNGzZVl4ppIBnnRumkx2H16kUR5Mci
Th8RohR0jvvCnBtEkGHaAd3DE7lbr3NKnle+4FQZyVIwR+DH5r2H5MQad+A4WnHM
mjDMcgJF4U75YYgb5X+YCRmYYXOhZM+wt8BOjV/iNGV6u4csaX1Ac0X4EhNiACzg
GNcit0VnmYk1S3po3b8Fuakv/PL7DxQPCAPazsD/k8yZcbz2R+cY8oaTtLSLvaMK
WuRvESme1FdCUQ9sLXmXwrlsawyMgR9J7LBhy87BbUSfbUw7csw97PDI0daeCCyL
32fW1Di8BKv6gdZF8cQ4DO7xgH3C0c9LYGfRIUAb5X/gNAYXxIxxgYcK0qviBerO
L2RlGd3cfp892tOkEoMHUQOUrjMWWX5TRkpqP1da/To4k/nCSR84q861TkiTENg3
61NiPkHx819oNO748xWacs5QRmvmPFI0RsOqA462eowmWFya1UIo4vjx5ewRYirH
cgdMdekIZEbki+pnrrlNPpl2BJqOShLZjMV+grNSuOJkIOKCuu6yXVHSWZcL8/Xq
peu7Y9i2tRpf1nhpQtUlU1yInWKs6aRCoT3bSnNgdp2anyhx3F5Co46nTX6yC/6T
ymZCRfTTL+Cu3b4azbLpq5uJc+7nJTTzRj8PYJgLiyoO8bjiKFw1w8fkAdW4eas0
r8pjlQvL39uqrB4rTLEip8NLpbTd5pIzp0gJMYtZzzDtcd4ehaXa/O1Pkb1Ghrtu
LkTwz0V2RGVfVvA7/THw49QcMuBK9eun5m0aViUWkbha6plj+Lui9QkOoz2JH4Y6
j+MmqerPDVmX8EsYe727FuwgL1535VanPLuctca9y8UMRNI0kAA3NsoMNOKwQ5hn
PsTA49YzybbbECe5ii2Piaq6dskK4cdxUxpUFSHq25OYYgJcy3Dv+63/c3vF1JEh
ugMtFl8R5TSvTAP2cVOl+HjAxeLH5UDMucftCZl9xmjZu/TnkmBR7ROJP/JE1Ps7
rJw2ej+3E7iTyXxMGYemF22grOZLeN8obROl5l9U4w+mtQp+Mw3ERJb2JcGQNXbE
JhtG0So3fJ6Ji9nFLD2yQckJH35ehl2hDaPIpdHWmjucuqG+8EgCUfBGCCKocspr
XBXfhYYo2KDbDyBy8WapbB3wFUFMRhmtBDcLyphUeO3Mk+0vmh7kgVYarZl9VRCo
Zoad5QfJHTixxKRcw0kfw0YMekPczC9euI6Te40NUXcOEyXEVBLhWrL2gHbxjSh7
P/TGm9OpuCFMfPia+Uog+506FviKBnKxpLTB+yw9MZ2+C4PnypUoogJ5/pBvu9zl
ryp5jkvJhoUqDsXwzQnZbLkA1csxUyLyhV9Idf+EJS8mKbATdJleFRzgHp3xGtz6
c1RsbkSmjDJ7EgCXe3uD3PavleA5OH3pB8+ECMUIi5wQBakN/UtR9N0pc2siiACj
5m8Z7h+Q9xYh9wn73M8ln9kJMCFbU1GqoQwdfcGL1KB5A/Gh3R/QGyQpYDHRX2OX
0fLEvhj71fDVhJTOw5Eh1ia8gxFxWSnbfyXTGzyqGlvk+gZFRSVSRlTMk1Pr0ojK
bAki/bu1p0w/9Rkhgpbk6/+/fz3tVYUtFN/pHEbdNNJP4UqetTAXlGCm/E1w2sR3
PFu6w1TkpaEkxMlc1A8v/lkyOb4kVEcjaP/2rpVmDwio8ueykq1w5VUQY4NuGzYu
6ido/QoycoO9kEHczZS4LijcA1ns2ndfzo3n0GsHgGWOgjmcnzAB4dqg1KVSAv1+
BmMCzB0MC/3R9AFQjGNdkpymEXg4bvUkbEHXQdQ0/pOOkpCsZLaJO5an974iFMpJ
+vC0lbi+ykCobpGR8wPYMIM7EBAqre/u1CZEH83Y3y9LdK9YR2v3oypYhmIhFyYz
CG6/0IglKeKs9DpmM0HN3QYgnKoXa6t8BLZibYKCniqsDxXGGkDLQg9CVwE02npx
bMtgOefmpoiIOfSzXo3+oL0dsplUws/qz2gLXQy3dfPMBtAYTcC72cEPdGtGOGCd
UH+kio5Q+KBXMjiyZp02auuCzz/0lBMRrWAGfyU6e47n53SEcbRaRAFzgkDT1gkr
A1M8BfQbk3pItn3R4MjdfHTlOcdHvki2lJZdDE6vFfrSw7vm1RflB4YdTyueLTLf
LZ5g9Gx3Hw7rI5CzYYGq1XLk9IQGBUu5DaHiEi6zlimXHFp7aOGhM9CijoqlQL3J
h9nCcHjdrhklfFXGqpb2y6UNHS+Uib4UZ+Oy4fKvj76CSvwSdo6iPyM4g1eyE9jv
xZkfR1jw2tWPrBXrk9QzoCbQqfF1Rx3IWtVsAE2SkVelWgH1z2Dno2nMZS323UPx
6ofD8i8uZgn/ye9crO4CGScTW3qOuF9f6hHpdtKtw+TxlRZmfbmfIS4VhcIMUcSz
3awi7gxutouKd6MwGYdaQGvKDxhLbmkjWtbAe/4CNn2o+Z3kA2mm8Hury9mczBTG
d7zg1FGGC8LiwypGW6jv3ZkoC/aN98idlocEHoGVtsc7tWMbxKrpTnFdlPYXzUDt
9TL/l9QsvWAc4Xo2oJKol1ZYUMHQl6nOwzH74bx9uehhFMEgRZxAm6IlBhCbyh7X
DsA4P80o0rEHr/SFCPQYSzqNhzCRSG3O7Hv4RSrCGg8I+oBACioYj2ffXxRkTg5v
0cQaEw96jil20baWsvKfd/oUZ7yDXdWRejPC/0EsJRHOGji/N8EfcYP7AYkElS88
VJ1Oa+ND9kL6kUHaqLTHAkDGbdNqdiKRutHhn5j11Pro4JGSAq2d70PSaix3oWIC
rWWNgFvII6Ju11xy96RbW5Dn6d0kE8Gt7MHbLzDf0b7aH/GEoyzQoFZZ+vB2McQb
2JaKRhGsLdbi2X5eCyAmLG5ZAhnQgaK/cXvDHjLm7auacNof+4uflpJGdki7/zLv
ZwwJSBwCVzDHOQ32H4IHrE+3DJ2a5P5nye6wMHqTXxNi90iQMRKRte0U/DIrR+d1
sL1rjQe1eCG1BazPw3btfaspyrj3nENHd2hSH41jJYQpZkNQjUiuMyUyJc8Fw8ph
gXGzAOih5nvTOfwhVMSnrTrMxYgz4Wbno8AVFW/mNjX1j1Onv31L2axjayLMkXgV
RtwtlW8qFflLxgE9Nf0QBf35i2PP1PqXtoVw0TVjf2kis/xTmJUJ27YlTaew2Jcw
Y0srpZPX1CMq23wOapjcA/WXvz/cWzV6+G82KP11VPjz+y4OJJTNdOO7Joe8lXEw
T9zA1ZP1ZdOlH0LGJ71LfV4cQjbi4oiq2ecRHz5F4Pvf5YnSTAyvetoZajMVPt6v
9NB9Ivawg/iYc2N+1bfYJCy59X1dv9nYbM3kyfy7SyOLRGFs4JAza7w1OkjN+lhw
gpXteHWpZ/hIpTdQlEfP+Rsa6VU6V6tCvefpUWFQshbpvADHopo2inwSdjEQAfHB
/VhWQ2X4Sxb2+l062Jn6hwlakAFli85pO3Z4jXC7A430MFMpc9KpdYjIN9EGq6sL
oK3b/2pPTsCvZ8KHpFqDvxRdfE04ana54+c3R4i8DYREn9FKICS36Tc2lA670ofv
js4prBkn5m8U/IBeToHPcIXnWK5EAWovGGQAZteHoSh/1QtlQ75xGyTjZaWanArD
sTJ0xdVONguD1XQ0wqdhGJup3b29ftoXuQLokeWgmRHGFbPKJ7rE3AY5XnOJDJjn
Zhc6ySV9ehKbMeTQw0gmDgLpddQxNswLiB19fjIdDN/ljVuVlyDw1Wl9wJt27TVO
g0wUFQ2e76fYBh2CtJvkAP7AVZyMkpOOIQSJrRUf2ChnXyS4PMEDTwqkYErsVzPI
50gkWwaALMXufWguafrDkaqgw1dQH6wwXt3aw6SEF61hUNiC/lw0/ErWZ9hsX2ki
KUSQXtyoSiGswnf/c16fZxFex4iiQWEBbsGiJy5cZeEkWJK+941zQiAsM95f5eWV
+IqJzc0wBUJfp/+b0egrZwlx5WYvmPJlelOrsldiwBHrt/fQ4Vi81LzWCkUDmjhq
uiHA0Lt34+v6EjrdKj83MrIdtl3VOoO6w4j3rYXfbUi4kASmOR+TOyFTR8K6erT7
ft/7elzvRbWlMqkGim4WCZEN1SVQiLxGZIimho5K1+djz/N4LELuGG+7xsBMDBsW
7aJGk+bfvN4qpGUc+HSlNEkrfQ3g+2VnaFVXHkgtErq29klW2+8MSfNLwnxcIHQ8
BM+m0vFqIRK19LLp8I3Wxj4H01QkMpcGsp6ajFLb1+Jp6lZhcVb0n6/izC0EoWfr
0l74sUdI4MCjaJNtCxe73hCSlXbilIVQIExiJXCRC8H0eMebg/DxVmPQkTDZZ45U
naTfmmQOnc/xJrgPd6hl1C1eMZ0GW/CWa8V9/8YNAu7r8IUPpg6OSGyxkylBBIz7
Z8f6Y+TdEwY0WWCdNgANcx8gbqFT3O5Cwio3J371RtF6uZUHDFB84Q2uinsjH7Xy
1/TYim3OV7QKTENdGe5eKC1wXK5HDird7eH+NVefPorSenKWa3F294LjAp5Z5vaJ
8UC5rt16PT9dcMAbMiZLZPtkBjrD7Xm+mUnYMjMeVkpkE+szRfPrHJCmTUdjepab
6AtO9ek/luP2xkQbHQhXAxDy1iEB2YLGPdr+jG8+lYgMH+IdFs+1fpsaBNRYkA9I
UKQ7EKNwKHXNPbpXnT6EjHeXcF3+puA1M1qjxDg28OqSlC3wUjN6Kl10GDseBpBv
f6n03sf3llorV3UOv14eYx/OQtL7dDGs9HUmWaH8pNMwuXRpv4YTxIPDz06Ocbyk
DZaSU27M6bGu3C57T3cwyeejQooZZP10GtgXSHAEy4T+l3+KYY83ga9VOdCrDmny
UMVcqdsp0CHLirLkTr2jRfKtiDwPGXJ8IUAUDgvpfFosDLh4mIRQSNFxvtOEQ4iJ
nnaLPdH9Rd7HP0ojZLVAM3wHaY9i/1xtiHWSzZj6AdyDJnxvGKUuyzW9oDNPT04J
TLwA6b2cnNrnYWtrPVH5Px5cfSAGYXvXthAgvM/KA3T0hPpzoDxXmv07FeoDhQFm
5PftyvOFen2UZJzad/7annmvv91HkcE6YeA8WkqByw9a3wp9kQswYVou9jEKqO2N
ChQG62+XC0btWa5kBzXB2B6vd9c0BjSKJJ2CpTPvfdUfzpumtTc3V633K1a5RYWM
yPJ3RfDymVph0nrbhF9HU9xpRE9JVAxZR3wizuA2HJJzfiJLWCMVXVXVHWY2Q/96
xrII3SmYnD/jVWjMjTJsZE+qubTAk0UBZiKj42YE3QbaZ7aari46+iMePht/uJbK
LwtPOsj5EvD7RyiYzaZ6aK8XUFEfmwvgsVTsVWs42lLm5NCUH6X4KKLlQhsc9Pse
7l1zSxqnCiEzTJIhn92B3Dm/R9K7qYrcVJpoyTuvUzJGGDybrdsz1wHB4xlqEd3I
dykMepNcuMviF/MGkA8yQfGCQsGC0VknKfuO65NPl+NJomnCMlFYHv4knTl1aSjC
gm5mcc2ap3GDf7hsSIa88WdrraieZjBSInVTSWJwkP+fYfWFkEN/EF+6mpMVJyqG
lngdiUpCeAFHdF4m8QdzYtS3RuM8sdFZJk3jeSkXbyaJlg9Im/pMa/5PRLAhB6G3
eg8e+Hc+UYaUpe1Z9rP4yJd1QgSUWFSUKu62LDpjmHp5qUWpUoU38OoW0PQgSy2J
yG6f2f1+a9A6I16x8vJNDpBrRooouYVHCZzZe8p9FuC0mV8501Om0TE5fRcelF3X
RHozOX6Ifpm68scKl8fEZDYH/K34L5yYvg6E9go8vFXNc3cf1XaX28lwQYLac0mw
Eel9LEXCONviSO8M398QfcexhzHOgtlddIkWuLzYDwQckXT7G8ePsOHeOWMn6GbD
hMP8CyCpMQvZ4YuDYDC3q3ItMFHN3R8pM+2cjh/H+u6MBcW1tmhDSMWHyp9YB+ha
f51rBomngq2Rml068yrdZtQ35f3TLYKqo+sfo+TZcRb/2Cba8YDjxzNWXM5ekFo/
dwW/g6+WIc8BFqXp6paTbEW/nz9BYnN4+St0UqHcDywN5SnX83nBPl7rCqDRP4c4
4lOsoUm3mD2WgcBRB0yxOlVW5anlUF+ttffYZbqFzDWgs8vH/vRMVsjuBJl9VVfp
RKDKqIH114+Y5riPAucYex/RBIigl4u6nnjJv6kKv/HuH3d/w+SCuPQe3plwpdKm
p/hJwLvwrdhiD/KOaCfG3pfMron/cFk1aXIYDoVYxTozPooSsGFhX8iHxL7MajU/
JikmeH1ad8uBoi5xBtwxMsk1cWAW/893sNPAzNXJVr+har3n+G6liFYV71Scauhr
1XRGq1WcQ2PyldDN+NbCCEEPKyvUbsCvotC1eL0K5CWshg2HapxB3bq3mmkDhrr9
wadeYOsoCEEj5K3wZ0QloZuUHYnnLFej6eDqD9TiTqiN141cqVaMIdM/4vYA0CFT
jZmammpd1xmMxkgc/RvqurFo20IU91dUnI4FozOLRdkFxrofJKOGuIXgawePJdia
Qkapx8iOpS7jjfzjNPN2dfJ6rLTMxjdL/y08sHFIWLG7cxptoKPaOIajn8nTN/gE
dGazcYMOZb7y5FS2vMQoaT/K8y//m0Y7uSosVvhQvl8iIcRg1ITUZKVfH1WNsorb
w3DODNO27KLaZcC17UICamhraIIqe4Er/Uge6ciQRKPKpT3xX8LNQVwjKwhcOmDL
+QV+Yh4uyGaErIzjkAG+JreH1YfobzY5YQduEY6Wap+ZA5QlX6+TGTdMlG2iUFbj
rBw3pcNhsaIpuiX9jxN/SikrPgvfwBnoo8Ly4T+SQB4CQ5tmnWm5+7VMZgDovGM+
PmRM/MztJz80VadF6kelkZORaDTTdF0pqLamCw6PP5DfOpgEUkrIln5kxNfoUcQi
bExiUjZfZXTFs1WnYI+V5yoJwrbMwHmdpWSdOQPxjcGGdqg+eZIMUUSrnRy1tGid
gDGgzheFviBwlh8kRjrlvWWDDVRj7XCKkSuc47PMJon4e+kCJSg1FSe278clYEke
edZX+3qjWrSfiJMm50Sh+jbxNwVic5tUMDs9dcCSo7AElDz2ipa4YG8ow/tbh7fU
/wUTeBwXxoKh/ibYEC1hT61/m0R0jTWLwq3qXpWMPtR4+qLsDCLT+6vcc9E1yHTL
yCaB8sha5q7DRc1P3loxcKdUZ4QCzYmmzxGoq34CH2K1A9HKETxkKGXLByVVob1S
k3rIg9/Kjjj5F5op1trPPW+Jm6GdxaymH3p0ZEw/+baB31IU89Xx0LorvRoKJ2Cg
DaemAWRHKTIKiGP8275kOAfxuMzpwumK5StmfMkVxPt6Tbl04wtRE63L7ZJ8V2XC
jyIKhIQKsNwQ4+h5OEtQz00btNzCtbMf6fKO54bGtlbDR+mN2DGj23Kwr1ibZF5q
esMwhWKJ/KEysaW02/CIrqKPVbiV1MzhE7QKFWVC9RZpMdloyVYit3pW9YlkOkZm
WjuYMAED+Vtot0hDZ5bwMpedSu6gyuyD+tyAABT8EK85DxYCEgY8VTa7+WwPab79
I+NYAHLJyYtiwvCIPiwr7S8/xu19KZ4ouLgAWMqmVNYpchZ4oa0T0U+dsWw/ANT7
YMcmZmBradKvKLuYigztNZRRSBhrtp+eiVU+62YNEBqIZjybkaEQpjyxpF5pvXZm
hlNaYt47zquUHlwF+p0TpHvAwRe+G27dPVpgL9aqv6q85H5G/eCdU4QLahoIBZTy
LwYfKc1pev+fvPBA5oRjhc5hzpJ7JON5nJv7qSmyyPMPsLSSqq/NqMgjhRwSa8p9
V8eHITxOxHpQQpktz7DzPKYRrnZ+ND0doaXwW0HRY1W/0MPeJIZb6sxyBTJqJaBw
vByMp7ToMf3N+KK2AkEifq0TKSovv+46qMx9zFU7Z1vT0pIedgJ4HiygEa9O5dy7
qJY3umN+luR0Wy1ESB4YwYGhYrIMgZMT4VrcF7YBBewp9jQ1W1ngBDmR17CSRYyd
ynT0rEnHtnRv55vHvPkEgSYHv3uSUmluu8T5eccsfn2IdS9mTXsYlu2mwE3cZZnq
tgZZWQNawsnjXdCBw0XLCaOazPN5bQaiCOLNNI4o+XPzc/xta0bPAnEUwT3JWgks
DTF+xDZ/vTNXDm8lTDKKzXzDbBQchBL7wWlFrKOTTWX4VWaQ7KYbTHAIzQZtvfrK
aSUR0CdyaFqGRUnnAn+D2YsuR/3BRNjLSNcoNcWZtDwemDYhPq3xCou8ZwP83BkT
9EZ83F/pZoWPXTPIjP27OiMS4oLiTI837IoT1tVwKluUTcxnWWVP2w96J7RM3ZBs
WlsWcM87dH/xIaegfb1Up/RorNETYxjGq5MwqlFd8oJZy5zYfuYEt2gGUU/8UQ7D
+7n8MtCEHex+2BfZG+6p8QjaxQs4vwLP9CdYmCy8ZvmfnXxllAKUi9UrlVMyx6y9
kQq0IvvaVtQKj8WUXYVAUVtPa617qpK8iQf0vign0LLnFnfqGbZ01ONEdU86SwZL
rpPYkFT9v+xwiJ6pUMp39RckPWiFhqVMZrl+OzvjTx5YdAyJWK1Yn7nooYjy2wZs
XOdZ8wBIFljbAaImbKrgpN9m2t2SE8ewBAAg+So7ioLAruOk573I7RFo7nw2D8zR
FgMSP6mYeTWKu1hTwt6HFclljUqWnl7JP8GjZ+lkYWXtp2r8SaaLNxc3715rm4YK
Gcf8ionplXDAeynPnEbYHzBuJkni4BKWhOE9RjFgOGrYfyad0d9wGVKdXQjZoiGn
d6mLCDMdGIicbr96ly5qfKdn+9B/mbeV5tUb4Uomjw/paOxpkcTyaP4J4bytTdzs
9jqedn+bqGVs+t4YWWSW0HDd7Jz5Q5ndNfcOsz5jcDvvhqC+bZjYzM36ioc7A06F
4pQ4gPAFb7rio9HdTfXhZ0xsnaRxp/g9FOOnnynCq5fq3i8tUriwtZLxPLo4mJFn
x3eyHlVO7Lw/4tP2zKOYs1VL6K3WHvPLAcdyIkA1tKYpKG2NoHhySCtCRisAezS1
I5gOTXouYziJzCtKhC1E/nSXY2eWYuzNPT1GNztURWY3e7L2SAwCO5cX+/qxC1se
0dj1CLbjDH1OSAdSwU1nJjIRDPWJUZ7N65FHCnB3IHSJcqevmi72qcSWWvMc2Q+5
QSTPFF733P/ROC/1ORnCAbhYQfK+vJwqv8tRsExrL3X9ZFW/wCrRwwDrQ6DEONsn
F+z9cBy0+syYYC/Kw+8wjExxjlD9bYbMj13GCdgLfS0HfKFBZmdhZZF7OEAz77W3
ISmB7ogTou6ilPP4W8EUqoEiME8x+ekDAtft5nkSwDtIjLuzW7nTamXD+m/UVag7
t1HqhatpKkBcjcwl41zJnQ0FUZow1HKFrwlQxfRZ4ju1O0sJdmEUVC2Jcl5fg78U
gwoJ9fVpeMTBOHLjWnXDkfQ/RU0kWZDqrxwEBG/R75jGISZD0qF7SxdbO5jF3Nmw
b5Ru5axBAhthA1Q62ndSGr90bG7srtAPXr9Mt4B9ceGvZOELUqFJVu3eQlXuPfhA
+6lnVknYYz9Go8o9lL0sEAcHVa9Mg4tD1Oh/BYYVi/IILCUsZRbX2+amwAhGifBO
wllqvDzdqbGsMIvtQNCDJUILNC118ZlbwUOYy8+BCrRlEoq5oh8sdGRNSrjSXilg
jVgLdszdp4+39hGbFytY8PSwxiSyaBg6WS3cvNy6T9sBHJQ32rlXYNSOnNKuymsA
W3z/ERHv2TD53A+sF2hJBuXP1LM0lyTbNmsKSupcetHUOSefWSVQhCEIcUdYsyBw
OqMp9B8nNjvB9Jwn9i6205q8SsvWryBf7uPmx7fb9HBHtNtFNzppmQIGAtwlNFEb
O9zBpAAn9ZxfUXuwygyHNLcgdTmEAsKxo/XcVmQ2CaT4bBJCUDmIuOhVf3i3zB46
rOU4K4BCsOavuuTyOlGW6Wx+qItuI1n4d7wbJ7O1sD7lOEgfJhILKybgAB4LJStG
2u0psLOGj3k6zqXnWvEHqDVM2OyniODajcjZa/qisXYwDuiwvvbhiefu60BiYyBT
4378LrQxZuXDEJVeG82CvuG1FOfHZwFpNqRk5BRx1ewFE0/sDOywtH5yTLx0I/6S
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EDFrhRKTet3Yqq1CzUMf6OIlmEid46CWy3Q9vkdf6QgujXnBCvckxfhmawcJtRiU
ULemsuZVatiADOhJqiuugd3tO6/geALw2QljkQiaD+OJlPbMl+z6K76OtExrtVuT
lFtBVb7iX8uzvDGimo3x4JrmWB51YREmf1qru1SnmQ8VgnlBj0svwlrbNtGlXDdb
rk+GAKGiKI+9zkmhbE9ytxhATj1VyajgWBgDGtRRGXBmWcPeulN/lns5SvIp5med
ZR70QhNNb6NTmhwPo+bbFEiq+FiRWFWh4P95ocxySE8w/vr0pinO0j78jsNg8SEk
SalwObLKaXfemGrRxpEt9w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17376 )
`pragma protect data_block
7YBf2ju4jSfFsHqT+M7N952L4qgQ5jZOhYjgjCtctDTfVAeO8EeNKQxIkowpOHIb
ujNKYYoTqjaDDlThkYp91C6U99HW32JT5pomsrR/UVOJ4Az36Wfiwg4/2LOx8fz0
BU2OgD3vd3jYl+YdLHL7HgyoVCxmqvdj32i+0tSXB5PHavU6lbv/FdyzZkcGYLOC
zPnHHwf7nbCBEhJWTqNY2+pzykZjkZxMeIynS/ZKpTZjvvYHb+mc6X39v/icVI0E
hsNyWzMwL6SgD1T7iMzS8oM09TkXtq8lrKceDJ6BwH/w3T4yiNwLKdDXwGMpuHSF
+7+/3YiAWUxCsuBBU9indGJTXG/OdN+xlxf/+gVXyf5JBHOK6Ds7BqQ9iJvqc8ii
b3nqEnPEK4fasIyhNKz8tr+kw07XqcmGcWzw0aNiJyKtVy2Nf/uCDpL8HqFx8O/C
S1Dz+3T1GlEzcQmy7S8Btg8ZzVo7guD/x6BEm4U9n+JbjL1zU3KnjBL4hksJ+71X
Y9hVBpSfJN+lMWLbBCW5yWEfueZx5f4DNiRHYPQQ8iNonPAXKgU3UAkfzeketsuP
IVNt6HqMZPn3nS4ORd3d0Zeh27PBeM3MTu76IOWmuVlqGixvh5Q5I8KpZHkgRcTC
saxweXxTkwd7oI+zGBscBTSWe2TS3gt2u+nxfYMNxBvYSrWfFFGK81HfGFWKPeDy
juwJ32+5pq1vp+t1AmiZGVZ53815lxW8YxkewDkimu8LQ1WA64uRazoZmJMzfS13
nAqeFr+sEkaU6GfFAKqQV1lsopCfU8T9zk77bGLBS/ukiDOZK7Ede7frEbAh1kXt
GtaJ1x00WbLXZZzkCIz3KiZfG7HAParU+SVP3Q9XYO+vNOFYXKoaUfYRz2fVaT6w
qj6Nnqbu3FEIp5y5lOqXnSBTLE8aMgiWq8WRSNJjVyho9Pr32fIDl4SxXyQdgzva
PwhrWGBpb7va6azJiQNWAk/SKEBFzXXrZLJBlGEywkn4wcUh02TaAn35V/OYLy1q
xiLcA4Db/JtxevnC81GhsiKGcaautGYx+EkxtnR7O4S6+gIbm6lZRMQhLLhmLJyT
3aJ1eZnCJepINqx3reHEKVsGVlvqGkRFiZhkFoP0TqPE3tpaOTbmFOwdpitxsCNU
GmArnCd4H30QOBhE/PIwVSuzI+vZYyXXam7xVB1lmjRhcCVgzBP/VNcvnm6FLh8R
i+anmGBZmlrJJ4yYtopMmc8hYSeg1IweM2lKYu4vWbVI7RSGTaxGpafZcHQmKX+9
Q/9Js6jMWT9O0D65XB2McB8Xixb99cxU/nEZC8LI0j6DB4LdvJ/XvnzkcCtnXSMZ
+gnY+Zw7BUkJhlinsJ9EFjGnjNVtlvBQ7IpTkVuOHFjXhUSsqnBEfbud4UEVNvBK
KesxOYU7GjM+ddmDbN6dxGRFRsBMzOEJ5fhYvnX2dO0Xpals3tuiJspkachEDk5i
yYlTqNWaP7ONRKLyn3QzgzfJW2HZF4onBDqeJCghAZ2leDpsZAATXateH3OzIJ5Q
MVtgFDNeDwwwJLQtHcFPAahkFO5H4NE5mB+CJO6kZLPzMOWq3AG0Kew2S+aQYWd6
hDlcG4Ex1XlaH1X/WS1Y+1qjHUHchDF3p+3U3Arh1FABamW2wfs+BTXWjLausOmc
ZeQYy2g2nPALAndB2yMoCMX2Qy4GmH57Sh4yqoo4Z72dmUbeUUZf2fHr9MwclPmb
eHSdaCjN2RcIrlpBUd6o9zksFf1bx3IvTM9eQ7mT66DKKhPII6dFUhhlF0eH2bnB
i/J5EWy3tI01Sn/pRJSouY9dhDklZnwZNOrQ+8svv8xSrSv/fWMzU3eOiyq23Q0t
AC+WWVlgT6qgjrnx7FHG1qShaZHramvM5OYiR3YExeVBWqCoPE5EmHejmZmzuF7l
DiKR6U67XqkDPr+JUgm8Q1ZzhkHo5qoXuL0IMDEkg/VqAWWNygATOr/rMJyFJCoJ
cpbTbkpHf9hukaa1NC2BpqHmOl3YTKXEOC946LjBpNDd3OzWr7WcZJIq63eHUGNS
acBPTYMCFWk/DwGGjgSy/X94Zaiwfq9nPirPIH0ry06WEgnj9vjS9fnjfIz0ivhL
5QhWQ/S9aR8+epDexrePZQItKa/8hmZ79Im2AGyoKRjqCeh8h9yipnoIgnpb+A3b
VYIeBHwnVlhoPrv4szxJUJCkCNJ3ShpTcNo050IijBl3OKP4ysANavkXX9c9ibKt
d3pcqdROpN/uZfy281HhPbGvJIkXkkFECiGkjCOazzOathS6YIcHY5C5VyAb2tVl
BnVJX4EWRQuAcZkTv/I784CIZQpVdTee9ULfRU2/HWt/1KmmglXBqCWKXeVoigtT
OaBVj92CTKWH66oW41VweXriK+9dXj8hOyDoR3EHzqm/AFDh379D9KWSoNNIqKvN
KrstIdHj2E9TPYMeIPVHNt4va38tXdW47SpAhAmaDj9s+cq4YsRoj5x70KtDTJWd
r21SK5QiO4Yrba83/jLHvGlQ1eeh43BQtsVWeDDdhW2Wld5tYE2dNw2SXMpO8ojf
W/0WM1DimuFwjSRlTnXVjdznMvLNLg7v2ns8pORNVW9C88y3+gUiA4lIOc3t9mRa
9P6PsZoL6XT7305VYG+C+HXtXR5l14ZimM9+v8QwPjCAx01/mcs674zTeccKds3B
+jPgUSEwz0kR/F+DfHFkgFNdlImY6m4IuxG5gYfrYClyg6nGqicmd6qfDM8ZRa0C
KDMrat50F23240Bo4NfjUFoimnr1sjbGiNOYpJu72/3eozroS9HhPqttD3pPnoY/
91lhcXSMCtM8g9z5yTLy/jmnIED6E9Ow7cRe5/gpk5Wm5IieS1pViXC77nC970EZ
I/SGT/CI71Lp7JFA5XqrmMWSf2OJOFcxuyxaGFdNYAPoQTEBqWYL5+nRVYr9Vq8V
wV2L97BqoeqRWsUsiOO5vQGT7e3MLzfwYWlfgZlMQRsH+xMNzmPeXOAPSQG2fNwm
+GzMTSILePA4OjkUSjZTolLMb5WXDTWYvzWo/igvJPPESUgYra0WvTLxq68PT8b0
rW4yerMgwi+KGvGUd/LNzd0xCEkmjOt0Lbxelnuusy1F14ldNOB33MI/0eYQA6nn
y0q0Qen2PNuEOyGXbjQIjVad0t0KculpjCoLtWnkxHKWmmkEpCd+rZhMBavYm/hu
cSKlJkhIKeKiYheNc9s8L6Lvl69IuMscCiy2ZHnMF5T2PoyNJQiBMl5ul+hcaogf
zf5UvinBV+lrmlN/sgMe7pi9L/ajRgfFQNNKbXEps/Drl6528VrlpdrNte74FOOn
ioBnmyu6KeO1mjevnXlEWPMR7iO66C2aOYJEwS3hic7Urf+G6faw86V4cdYuiUsU
B8387bo8GVtkl5/5CBZDkSBSQH7QKOZaiEnORx8AQUKDPWUyMtVjodzjgKIAkCnx
FBPyahtiBiPqEa6iFkzRPyG1/ipVe7/Q21HXau80LzZcBrWvGQmnFxxekuGq4O8n
mFEFayqbLnCqxP1dL9GKXDWvrPVeHJ5pXC8izYYPnSPTv632mKbzKCGdnof+iyfg
1MhTwf/6yLTNNE+jg9BYOeLXZFnuY0jw2I90h7W5eNKVpx5q8GCMetoXJrgpOg0R
l8YVv7P/IOT5iEsEZmXhlI7tu61V2igrq6ijgGQaR37yjYwRC2ytTA6Kgx5bL7nY
WjNFBIeDFvXME1XWH1M1RH2bHRnSD1i0d8yKUhSMrumxwBwskPsnovNI+kcBLmFS
1FxDevAvXoOXlqQ7n9jFdVGUBSzCFDsEWaxXOFFSOc7zT16Zko2PbMcNXiOIfsNu
0jOuj9eS932ZnupgbNqym71WCNHA9garVR7frCbAXkZeavYp4MyMQu/po1j/vnwu
vh3zySY9GBYTtQhCl5BovuCXM1sD/ctIwhhAnuqqKtcVcbQfFkNz6S+WDlQw7VSX
EWHe4Py8Mm1lwhBpcUBz5yWIRhO50zgSQMYCpP9XlJ5Ud1/wZIWWse44rj4BcmHo
g1M7cOl8t/Q+P8yeWq5Sm9VLx/YH6de2REkBOf7dSlkICHTFiKq65YQgPeVIicds
S+YaQ7RxXc3AOAPCmYP5IT3D9ZzK2FBeloNDRCbVVfLLd88TtFka41+hkDRXmrs5
VZofKJyGVG75CbumCRIckoTO90U0KmSTrZuuT40cPeAGpYnuTiDYR2GXKtYJrO49
d1q+iTKa7+PAqZ6cR+nNZ/Z8sxJQ+O/CLvPlcLjNIWQEOzn6CR9mpuq84StGtr5a
DUDMvIYyR+NEwIFGdkZgeboe3D4hMm/5sxyFr1Hj09/QVJn353skAhFj8F+PXtYZ
4MFKQY5ViTjXxHc9Fxo51sNE/9dFybikQEPWnuVJctpu7To1NGBxG54PGNvSg0Gd
9DniSmASgDEkmtl2dTmDw5eUPr2YHdIcAWsMzfkV/c7aHiV49EIa/rkVxZEdgV5Y
MekmcNo4plGP+A761mqYDBt4yR0nnJKlWxYfLiEH1Vj2eAAl5OLpPyFhnxG+2DC8
OyDgRT2C0bRZ2HRj+bVt3FG2Lgo5wyKcRf8uGrT61O7Fo6LWEALT3DAV0YrE3lcn
Sf2gkaFqOWZern/tSFnofvpXMI57kjQ8nu+r7Bh141ZONJqy8/6h9UTI6jFzGxm5
7bGuf8kO9BMUINa2sa/RexZkw33ivvPSXJX+3Ak5kMgn9ggJr/d6GERYDfeZxbjQ
o6tvtVB0AS4y8L8ZGYHRh0umOue7uHwm0eri9B2SKai/d9KtKtUTq9xwLysz2v9B
U/MqJwFuUb8AlEEf8+aMYXz7cnSwBMyJQL9ASvcDcL5JObSxQaeH+ZE5+1NJH/4b
mzvD5v/8+q9x/WfGTcKxot8CKrM6r5BKUVRmgKgAJHWvWb7ruexNKZh6cpPa80fL
j4E+KLqpPGZ8DMvlDBxqK/V5wSNXQB9zwMo3J9d/AFe+PzdHwBAjv9L8UkW5aH8r
/P5VnUeXf/PTecQSTa+elXEhlSuWO0dnXo5oFppWuQ1F5TDBaI6oj9Rn8lS9GplI
5+uCgyglbJA1x5rftM8OFryy0yxEukS/PHdROhHV1EDNLr/byvSqnEVhRM8zpbyp
82Mkz3rM7HKToOBYvVESsrlSWsovk3xSLm+6JjEmj8NhDw53ylZkyOLQ5P3EGhdI
od7xGcfOIa712SX/l7/HhW8zRDb1s4H5QP1pjo9oWy8xmiBi9VHX/5XnKUBw40nH
vTHKMrEd4LJH3bYsZ4J8KeoGNxzisXRWMh1C8QgVQ2iT85wnHjttT1yknWIYyoz5
2Qg/ssHc6Ie2gF+0EuLzI4yzP9NAnDYEWNTDP7ya708Czs2ee626YAnqhJ+L2tfQ
Eph9Kjgz/q54DhSJMoz352Lw/NUG5tiOYVfHGopqEprKenUk6AGrmTiKckg9S/g/
8tveOdbWDErw5BxZaqJLaVVAPXgnudQcAyaJCG+c1zPPttF2exY9BsFakqE8POuH
KEQ7B5zlAzeSypwd2vu3YYBAvaYLGQCDs2p+zpBjTaOUkX43oF0ayNvkYCvbHCRV
8kve8eTk/7ili1S20S6yj01aX72xvqbLbAcLNpBG35/+AUz62HrdFlf1GQvNTmUs
J9XCvkOXjM7ZJjeqMI0qkw9FBttz0tSAmZFwh/X/vZnZUoCjGKA4TkzlL5Ww8uKy
VsOj1qhG5+Nk8uLXL/voU/wM1vtzvtQ30J7Z7dg/cskIUNtxgAwJDEY6PG1BzB9b
lEYfRu/e4y42GvxAN8hq3vzwJBuHN0cndjH+qRIef6+rHCxWVa0YuMIWvRnMHJIg
1h83vWl/SpTRDnovOR0suh/JPfTbdLQwQ9cRdHZULIUMeB3EVvnWCGSaII99v0KF
MKR/9gyQaggzNPZYRKw+TOB0hbSYS4XNcwTPot8hAiIW3RIAso3qPWVTMIB/Dwbv
S6HCCIYWODotSh0CRwcfYocM5qY+7U+vNulg9x1u6vfmocxR0BSDSaCo3pKzXIzJ
KLWcuRetT0qR81tBWkUfcTzMRD3NMJMjT39HP0STYA++ulVhnXIW3zNiK2dAzDMr
wq9FVjnGbJuiblcMqC7KE2VZzbpWxVVH4SURqrGYbnRdZx5M7O9rxAP5scKQmUEP
9OJfwtj3L2QoP5GgK1qo1GKUzH5wD+REPEI6EuZXqtCmB4EoUfWMp8uJQFv63fWk
tfCKPtrqyMjGWhSZBeNE3Py77uEQ5/RYtyBW8lMBbChKRhGjrf7T33BRRj5Kv20F
tARWFPPofC8VLJAb9vFdiUK+OCugiszXrbLlegmSrfisfZZObda6lxsgiXnZ1Hsy
8oPbEErXIUFS5F1bMapKzoGNn32cZIIyqU6BUPN9Zd56HTWNleecgj4dOrcSglVu
Nd1YJs4YJmgHmVxCcsahoqB7AbCLrE34eFbWRCEjnUqWgcF1dT34hPPgI0SkvMyW
bGr3dcJcfx4e+EC7ZQm0jAmOqgrkIzDvfjUotfpON0YBl8CYs72AgoCtE+d8iNqk
SfcmRfLA4+7tNVmUC99/ONKlZVoEPWBx0qHPxgeI4UyEgu78Vauoo7U/Z7HPyvwS
XvYHcF82X3qMnbsw6gMOTksp2mC4dvxxPLSD9Yo3G9RKiZUdJUATnDkt/ScDVUUH
RMXwr6XhhoQpJhPOgtHFEtM/wtw6GnOTrqzhe+m6p4jUGs1CswDOUe+WKIJorWMb
2MfWrqRn0/sOXqHe1B/sBMqyXNTT54a/+ORbYOx7veJEuE1osyD/gFWOQKdplhX5
IxsyS7YdxAZlZq7cDYCHWblkYoidKYLK3TKAPtf0AxmqqvYh0JgQnEP+wMISeuA1
/sm/CVD4knvWOTSpMmeVpx46ec/kg6VbsiGJVf8M/2r6FO7mQrMMPz3u1OQ9JUOj
HPcZ2QOoMb3V+QO1BCWFGOZGPc6zVUOrDXJLY2iif4AMmyePWGEu/SwPMe304NbF
S4R5Cn+f1JfxPDSXQrj45/PxrlPU6oKRmTVur5hZA2QiJcvkrBFzf0YpjZsyR9u4
S6tXNBy+Zv8bosUFwcjZ3UzKkHQyAk0/LrWuuOgO50tuDp0pPHa5UgpBhRlZrm7+
igxzbpdD2PhtzIJhywhSwE1Prn6mHZWPiHzM5KzVA4y9Lp98rXYw0lLpY0pNHVBz
9mVWBO2s0RobykMqzPImZGwIebTa8MOpBBfgrz5FFBSqc2IkCW0oSTM0VIC3/Lpk
iXUJxkrNUDUtbqajONZc2fSP9eNqyGmmtS4/iwr+0hmeect7I4dm2zrTtHiwwaRj
9LsP38Gh+i8/X3oUafh2Kuag2XKkdqCVPPlINobYZaIPGx9BHOY4TvDbGSBVzF8A
J5sCh+gMRJnBhrqmEQJzXn03PJtHJb29pkQB194+74NU9/ZsfnNB1Hmvflhl6Gv0
VaZFnkKYCCOEgOUCLCNu//YIH0Mz+dhcle6AZRscG6KAAIhcqyBgjJriZNjUVYiI
QBFg9Ye8fZxmtiKlGm7sf5rHYFs2g7l/U8hM+DqH5QLNO1aC3pwLxHV4txNV/gtm
KEKDAiLZ0wLxwBX/tQYK1NhCv+O9Oty408Gd78+LFjW3EUUlPKLhhqjhAlGz9cPk
0NucsWL9SBb3qhpSKxMAFGW2N7MTCwAt0Fkp4GE9INFLq3otwAGh0Vu95CR0wZ+M
fY7+Pnp/BaGPwWCSEnOcK9ObIVyWpzbtVckmQDHCNdsqa9XqWVcdr8oJP0E5tkmT
HzW5gg4jVKF9BXJc6uJtWVOc+KEyE70RlHBPF/sqnNjogeSbDI86E2ML6sBVywiW
Ltf42iUpHJa5FSrmerflAiG9/fF9RpZdaK4noPAcrAgSYV10LkAqnjrexD/rOSs7
YCKrzrpHHnO05IEFpnCusxkhtbKssmUI25Foi/VrqFqvu7EQWhG7uLwj8eoDwgfX
dtov5QRkyVkrhxISKiAjPdDaV07OS+zISOfkJi6mKxec2ITO8Qa/ziUY99k2WIpG
fbqqR/gMvMtWpz0FK/qR27OLYbZWP2b+a0oOzwkYiTDo8nUqinJ9j6mjLeKXdwXe
qXI2Ik+p8r6J1T+E3SfMihCC2t+BZi7RzAORfFV0FI9q7vzEJbdUk6mb1uNreAjY
xfsO2ZtaxBxMzgOAQnl9r+FL0Q0u8BH0ebQsskPkbLLqMIbR2My3MaCiWjTBw3Bf
CGakVXSKc5l1MQ1ViWOPOOPMZrntAkCdM5qPYkw1lUKTuQW9cTJcDzGV+pu4MJOl
nXi8b5uc14x+OQpb+9MCEw477ueGFrSjI8Q7mn82LGi3zgGYgy3JxgTIaIHw3aRK
RnqHeixOkSLAjoI9SgRjbdrWUwiQ4qLgJ7ChVCWCXeWyXoex162Qu8vlTf9mfPnN
MLGtkP47E/wsbFLmD9KZX7PPEh2PerduEqQtwQO4Z6s1ezwlrVp6iG9WoicLvzzJ
goD9YX6vEFxSWR6e7trY8jA2d3gtwR1kDN2M91myGjKr37fcIdJIDZ4ilgxIvXdY
BbzLqbgkt1RDG2x3vCQZTfWK+I53nY3cIW5guZP8DFEg6xBwzGz7cE6pwbEAefYe
jsICnBfHbx984sBnuXGiLpcIuFx+7wjFeh56Q/Ry6oMzF6tuOm3f6BjtqZ2uP9tQ
fSc3ouo36s3qi2QBXKUv8xHO3Gycoyx8/Ly3QvsAgQPUBqKEjUENGt+g7u6gk6BD
yCTh8mnw6Pw9bEpA+aKK4Q9RGtpV6pZfAjSPUsSrdaIdbirkhZBK2hOX74IsfW24
cfYKrpdlvYVSU0rFmd/K80a6pVqo6vjpiBt4QjUhj5UHHvRNe+2sK9HSzeAlUIw9
FcfDr3QWPO3ExjIAfJox4SerT0UFzv+oeCnCYhi3aQyXl//+eNBUBuryPX32ki6R
8z/LiFfMM7+7fBq+9XbM+GG73CNfLu9cRhbum8A2k4CMYWBzZQ2n0z4lGnamCZ4t
mcDEBkbivq5P0t2eG5O4P4yIx6lIYLh/npI9NkJwN2CeOIAitheur4th0+AZcEaa
GD1B5RH1/JyXr+YsmAUDptI2g2OyV8Bny8KAwTrmjy4ilx5oxsiwAJGTUxWhiHyH
plOC8U7I/mAT2tY0qsAF7R3cRzBk9bUzIiCyzz0k7dZ3Sy1Xt2ydOnpAcflsmAhW
6OLW2SQAmSIQf1f/2qTdsr4ZQKjHoJihGa2+GYoW8VVZvnOZEIT5qGcnwm9Eh8+O
p2l6IAHL2YuECP4IYDcncDdDXt426q7YDhq1YDncg+m+WTjBn0B6G9wNPczPdWo/
sh3rsZoD3O+gs2CoweMvMGQomt902HBwMNQjPiGF8xtfk7k2J3BYV5rbMnPJqk/L
WqiiTMUZ7w0+bkIVc9Ky0nJ/VsP9i2xRSo4a3bIutN0s+kjQ0BXliv2KhENFOC3R
amJB/gmHs94dSYlntTuuV7IwGkWghdoq3Id3wUVoAx+YCzu/wk6ox05bi8ciHAO8
K/Hug7Jgz+yOotcO6mrr9ugO7dgZbWXZxNbvICEB82R6oRBIMrkBqhJU9Tql03mm
h05SVlKDyIdbzCILKoib2p0lsSTlb+smmhotaXzMree/q8ZPtzcUo7GCN3DA8/Cz
OpI5I7xyAgZhaq6/YiEvcmL3Cxi0F1gi337qaQrmOcRun/P/RFpmDDswelx3Uo1j
osIgfbX+4hIpNAooG4l8Ur/UxsSSrR3xX2n7O9Xamq0HAlORAzwuDNPkq3VXXNGT
lDx1TLmfB50znIv+UdT4s7Ipa7/Aa+MhofOCSGgh0459ZQ5Z9t0EgvXyJ6OPqgQc
0u6qXyXDcTNXDXYqy5q0JB/a/CF3KsGKXCiYs5yg650dVj3ziDDGyQlEEbjbiihw
Ldbl0rfwVVKEDs/D+j10Wi303WWJFAtoqnkJlj73235S1CCVmo06sJ16PC40PtLQ
J83mVEdfpLTaDTCD0EMYfUXMJ4YM3MZVpg9iFEEPQKsHlNp/oOJjuaZ7A01HS1q2
1xnTvwvZm6Pv2L7R8CnTWfw0xlG1S3uzN9NiAeJSHQ/lDrOF0ax0ueHQktuwfTdS
mS4kXhOlZKMuJEadoQe+sJT4dEZVGi8kbzUTJUpUmEkZSrVQjJiTM/1iRL9ZQuDw
f/ZwxypnR4UFgFJOYigQF1M+TbCGLwNREkqeV3A0AV8zJ4kGA9lowsQp0mbRm0jj
dloWGrqffSw8jT1pwI0RlbQ+caSUvPzi5688dTX8Q2UAeywKNJl9CU5/aeVxEfRV
JHoKHEsMT9ZHur4ouwyoYebbSMWAEaVaBHBVKSnVAgDKNg4C5u9wPdmofaU5ssMF
8CTtPxyHTfY7p3OrSfUAIvlH6nu9EalU5T1y4nFbX+gi/c55pRVID/3a80GK4hON
MzKaBtfTDOVPLTDX4YuNPSZXK8gEk9c53Fmpol6Bw/prYZpkOD/l9mb4KM2J9ql/
EFLCndi0nhQhc/202259/bCgNF+umygoVLV/E8uGXaIwS0GWNJXd3Wc5EtUGfH5H
BH7ZLxwdISly1bEG/RBCoFCAS3+RU/Rywc5R7hPVi7gUm77gi9EWOdYVEszp44qs
j6faxjZsvTEnxD0OX6Q3IusGA3IlaFwRnfyODYeC1u7JNa/MIFV6PIj3sieQXHGQ
tG5l5Ja+Ebo+HyCzBdvIU/NL2Vw9h8MSbjRkk74E4aI3Ow+TjaKPmkgycGepd//r
nMPrW25zCRnKTCfSZUUIIwOgbTmMjEHvsQFg+eM8djT5truETvzmV1AAap6e6Vng
vol48jWD542sE6AXKUvq1j/ffBjb3q9xx2QiTF/Bx5WAOYhCNvQJ92bBsiAQ79Va
G9iBDb1LfoDJ1ZWF7d99UGLVHsRfmLpfClMljuT8imxxGfyw3QZzQgxiX5xWmLNc
aVYzbwh1PQ/7oE37ShU/m1nD785FDoM4UQJNlq7GvuxWKxHnOdHrJDUVbnaKTtlR
KEWmfe7PT6vVuTtvrkrFMEaSwryuwpvB2r09U7AixIVTZA1OeDeHK5jU07vHL9N8
9ZmR/jnscJCY7ihdIYPeFg1Uv+LDc4FWCMDx1MXnpIGtQTssjsDsvd716lP9CJOK
XXO/BQ3jRj7fhE5axGnpyf8TcZXfdo3PbG2jZ5mPWV9+4ixqKq614JdPiXEkjeKY
GdoHCVlvSbuKeh7431Gfzk4ziex/0b1Jp52aaFeSAcQlX95kPBbrIhTpmW7I1KPG
ObjE8Axt05zkHzR5qKEHa/p6VBK/vApOkEUxb+ERk9pOutR0LUtb9h0e50hQdFUu
uSjQHM1psSo4We81UBsz89Gl0jSYf4e0Td9IwNE5rO1EY63kK67eifyA6pRdh9Oa
zuv3Jw4Zz0z+mBSP+wYShK9tiyPV+aZqhvc3REy8MmZg3NwXQepVQRqmRcIL+MzG
GtrDyFlHN+oS84XcHovYFPYIES66zq103SFUga+6ZBzCq0a3KAL4gdKRTuVcPwuJ
rlJONCdoozxv0n6jHWv4PGc7ZvN2YO/kUIL+HL1/XD11yDvUsjCGlKeZ/as1ACmq
J38Od8T0q/hSCU4Kh8T7R3/X5nk+UvWLJFm54vODDNDIbMzQBOZ7Qd59YEikhnfT
ni39x692g+r8atVtFrZfhs6Pg5qolffoG9hvFkddoV/U33lPaAWibfRSCxfWfidJ
Qx5BV/Z+D+BkrNb3TJZRfLoAMwlXZFiOf8ESybBd8uIrpZ5/51akQSq98qaE6Gtt
bvf/axXWFhpTs6DUr1g+FTzPwRhrsAo2mIoqUmuQiA1soaievrfQvwcuDfogCIko
8OHm/HyAlqRkcNSAYrX5hswQncCLgep+PNfuHVvuY0q6ORKy9GWtcSOzM8apLieR
GbJV2Xoo9EYe+tWeHhtk5jZcAbSJrlw2H9D8khYMmh3AwgFCuuF51fePNTcEcsmY
XGLL5OBTbWZGDNx9XdOEqSmmQ32b/fMFtvImaIgrtoYCSFOUT9AiIZog1P+WgYVb
CGPzAburmyQpNP7kfyd3QPhmaEkJLZXupBojm9tds5FdqZ679Z4f2VuTRHbGegJK
T5sZnTb3mmczOhtJ6uACjyu4qhYbhJThSwhHWhOvRWRubn4fpZ9L3CCmhUjtWmxL
2ylr5SuSn2kogkQzeiZXXdb7bCnSN7Tk8aajtMl5EqmZzJcohET3py0ancZwY3BW
WTCFRejQneGGtxsak4ba7JdO+tZGY1eHDLsrJJz7YUqa0KKO/aR/8T51s/jaN7wb
fjA/6+IKCljoHgxyphB8P0ayBgqE4QL+AK7DHZYzvnu11jag/ctRx34KJ50IiEr5
q2LfPTcbIQOxGITT5rjgtqUHU5JUyaT8tTMd4U9D5bH8poskoF3ueh3qUV6CayEV
NJJzJuvzB/VjAPZwXaR8MJmRJ9jw7uiwyIHqqCLzXwPj6HHNewYldltC+ba/TEil
feYg88TYpd0puGCe/QrzWQN+czVpLPuj4M8gXzfYzTC8GYHudqQS25i2kytxuFkI
bG6oxED099On1pMLR51Ze3JAaAvym8QWT67HY8cb3S45eBGUScoY8eopVTArsYue
spCkqXSsnVXv0TCE9qCTEAKz8ALsZN0kQ/HvBheIck3V3RZUK1CVvkhHPmStbvzH
bc4xaiXE37z4tf45jbxNknrGU+m4zsU+SGnQ7FBM98MVzQR+voa12v0p1lEGmjQ7
f/gjNH980nsWmy/cJb6m2ewDpTaLm3V/tE8A1J6A9OBuUtCpeu2N23EUP3fs++Ev
FmURDAEVbbmHXhdJA/mHSMkmD1AJfWXWXpD61peuxayk9uIxODdOot4H25hf4JB5
qwsF1c/k9X46wgB4c+Z4cxYGnM5kHXMIxOn4rxnkdSmI9grndIcZNRCyOFzxW2ya
cTEWui+yWIXoVpXIb/RDUavGO2hnrc0yX7UIcEzEBV2IGr3M8NRdOt5SJ8sCCJli
bxqI51aqif4rphdysjhXu5momyz94qCA5GC/Bgg3I658y1aoGnPmGIdJDiNSho6S
Ii4s3O9xhekyYly5BXIgqIfGmWX5+sVkpgOuSKRGLnsm3+8nytqROMHn58Ec3rcg
eBIZTpy2j0Tk0rEXngB1/DfKNjimUrur337vcPequqIGQ1b6CjQnUHDUZq2pryll
7zteEQkhDWvcWN/2zENi8gQqszY0IZFq9xuDfPc8G/qrWLE1/8CwITdcjLO27rMi
eHMr/DvdfHrcE3ljQprzLjXu6g7LPMTpQhG4GKV+9KQ81A7tNIOjk5TD46nMCPoE
XsEmFauRBRKyeZSZbnEVQhaRnhMZDtb6K37oooIdlgTENgI0xsKZtcoKjEHHlwdO
WfMogfWIYuLuGETdyhfoAx/MPZA3Hx24wUyAdL2Zj7h/Z7kwYKtdZxwQIFzYnWC1
gwGv24VdelRtRZSHHDQwRdW46FDgqbLgwICHnBYen717NqRMRCr4mj9PzL4D60sZ
yWIl/F7W46sNgOdPr+Y2ItwP1AGPums4FY56RISqTCA2sRP1A0jMnEWo2A+NRV64
dn+rfUpJ9zJGGd8zviUBkkHl33k6VIKjXRrkarau3YHlEbeVhdlV7uA9t5BjOx2s
sEGNqD0fLDl7pt6Hqj006XX8q2O9KSieZ+7Bv/I5pleRQaoUeJrp8yUFIsyRQ0MU
cdlyQHPH8kpobGlXvQvmHDCuGww2SFno6RPPtynVJEA/uHxXUdLIeve916LpCg/v
4q9ZJ0u54/o0juV3mLh3n5YhIYRnIWzuXg2pwHyttiTrw6TLt8b0T05rTvtp+gPZ
isi3CAf52P51Menfwu8+1kl3t2SEdcpM1wZqVczacbgyECz4w1zHAsH4X45tAZSx
2k6wB1MzlUm8bRCtQR21bJDmxNaKpAqR20H3r5vnbjxaP2GewKvY0uYk3Ry+DlzY
A3Y6Rki2RObaw+lg/OJEaavsMxZzUkCdUxY61iMu8apKIKfH23P5I0Tddjc8DqT8
56F3YFev/BRsEvUc+/GZ3Oy4YFPVuDC3/InJkqssALATU445Z7EZzkwrgQPV5KU2
VnJqt+Si6KW+fvnXJ3fZJ/zwk1/RLX9524s8MvTfdcQytcvq9JRelhbcIgGMpqWv
u3YHQk6r4CuwzkRAfZr8o9ib64oDC82bOsBfTDlm7jEFu0wr5Gl+XttMpV2wzzaA
Mt76jAk0L6rVEOmEEFV8QJ9u3iLOZ9N4+DGCAFLLLfvmVwY6baOIjgffskS39pBr
LXAD6ptqlud19NorHpeja1SR/dUt0/aSel+GEmQ+eAaV25lEeIyj14PEnc5o/jgy
wCC3267VpcIIAzUXOn6/Mh0lsx31ePJNfGqgJz7r2cEFYUm8J9q3j5ocJ/tKpJVN
HbrpDTJGQCRLNogCmTU+8aKDIDbZd3ksfUm5IHGrnLZ6XJYwQ85Y6eKZQ83kIZAC
//wFgyw+dAY02FR31ePBOjdBJCXTX4w3GiRmqZKp6UKubsvH+IB2jsJvUMYSpXci
4fngKXMl0eOpmsRZBSXID8RtLa3NWzi0Ox8i7o9iky4OYs3i6fiFPt9eaTocbeGu
1lm8P/qtvOn79MnyL4tkFPWirRgeg7F/ay3jyDiW60OiC1lm3P0pbdxVfZ+3QqZc
BTwDRYY0/0T/7VsWzWRmpSc/4KDZ9G93Vtxj9CPQm6ATJByTDFU4nx5j3CoR58Kc
TS6JMxEiyG1bnur2GJAG+k2Q3U0eZ2o1PzCc5m22Dv2o0eQvr0qtG/4PO4m7VgIW
tkwmOnwPxQCqFkRwQ776XZaGxMTkFvg8JXpev2uRL2eM+amkq7eM18AavAHl8QUY
KS1So5+vDMTTDcg0DN2OdbxY5EMTAnbJZw1q+6U/ayg3R6bc//IXJ+Z6izOqibNi
kkLmC8AFW3I06tpIZG9WhfcfTvIPSOuksl3STkhbxtdqHgOanWE3naTHywsoynk4
vBIp7bDu8SzzqUQfyrbUpZSN/PKJKi7jzCcwH8EQdVb57Uz83q/eGtmfPiu40d2B
2cfB1LwJjvD0v2QaNT9xykFEZYdsoIyw5NEJobZvN/ywekx3IdRr3sHA0wVnoZeM
IPP64o/G4H+KmAc6jy8PMpbF69lpVR110Uf0SXvHuIED9INqrNibEYQa4fmEs31o
7KEO9E9ciaHInNdagcFNQrnwAE8tp/V4e/9EXg3zodWqXnTPJuxLG+/Xrh3VbRE0
nLC5fPCJyHiZyfkB0QJ5adCDWnzVQ8ttK5p66WZ+MZ9KmpEXBU1o82mJQui45NCH
gxzc0ClKUHaq1Hnr4RWZpK1kDFOsUWc5BKqPHTZVH6JYXNi6qq3FKeHu/uIoz3QS
heilN1XHB+fYnzKGrXLsIJ5bj0X3jIAzvhllSXnOoZAYjYjWqWQDWgs1G+xWqCrV
zEU2hdl6r4a7e5Abw8vYZTn75xHqtY82JVc/Q6KF9kA+dHAdwas1+HFEdIR2zDNG
MQ7wmrzeqoZIgHWFRU+4cAdsH0AMSzyFJyNw6XFbtHxbPbkAcROp2EsP7TMfJMmg
8YXdo24nAJAjWuLaZHZDSsB2XZxO8hmDYLcD8PH0GofYpIXF57pBDFZEsuUxS/Ze
C4/2RK5+1n+X2oVdNrKBtLxkHyzgCtwgaaiO/D/NJRCU2GvRU6Y/nL8njIWa3bY1
dOlryrXnmesxNfzYqkJCqnjrBFyIlMMBEyieP536lm85WZfyM7IJ+ijTGbrK3Rse
AfB4HaDOf1XDzdQlSFf4mQphSb/7YgVj7YHvuWi8+UjRBRDHPmJ20lBjcmaVYb37
a5sHKU6/YQeOCnxfp9zFt8pWZVwxTiMv88vZIr91FO0B0/ZFdAmMiQlwhTqVgWny
3JUCwqznmtU8QaHqdBPwV9WVfiFXvK0zTO+36QnAbFtnSv/WUN/4JgBgdBp1Tna3
hWn53uRgiQ40NOfWNgoazdyzLkFcAEfUmytlxW+gAzMCqnYTDNU9UNYAGvh0qnZV
tvBRAxG8VbVcJnl+2SnVkRLTq25DazA2HOuShOl0634n9izcjb5iRgxH3JT/mJj7
ebDLGcRII/Sq1ZAwJFGfv/6Hd5b0Sm6uT5D4Ps/MSD/6z1GhcXSP21NncwxuVoEZ
HzEJfVG3IIEwpmhGexs2+Z1kCgApP5dxAtwTm62W5k4xznKP6mV0uEjC7abvAGBA
8kci4MtqPhGcxRJ9ggmornfy1XGwf78EyQB8jka8kkyKUXL2s8erMZf6RP58PZUA
3JRgaGwF1LwGcVfMQ9/46EQIrE6GrwBzrGtB7mNkotYiOxjQyCeIRNV6M+2WhXKB
i+fyZ0koiRA5kUfsFQAW1njzyTqcNRmiW85Vcg0NQ9Jjef8HmVfNWbkFvFsr4oht
Yn/X9a3wqgBV7Dz9nTskFS0ASsn+eB6CDQJQzn3L7kp7bZYuKwbJV2OT//C4bemw
yEvDUoSsSmvUZw+Wv98T3zyCa0qkuPX5uSCOqETP5RrP45GVf4S9V6JdRXm37PmJ
ajIyFmLCQB8qa9s9seCogVNs5eULdmkkVYN2UuMRxcqkNd69iJ8Mhs4N9TQKPkvS
KP+JrBdzGSnwVbkvF3buT7FzgQpHW/rplkY8ZRUSIFoIecljvPbf9EVBt41CSyAm
qiMG19OO6un4viZGDt281njmbLnPlaFpFXz1VHaUU3Uwzgi5gjcHezVf0reqK/bY
Ddi5kIrfRKSaXUPhMQzJWclwEfhjewO/W0CRzRFoZEo5znhiCCiXxubzCC4O/2pd
zAQCpnp6m3SWIJphI5AQ/avrLP31xH2GJ/bSna8LmQd71cxbgJBDbv84XsrnRcaO
PNeqepi6qyXjbYv7uf2n3kzQNXp63NZ07Sq9MdNjeWL4/eLO0yMLcfDkiL6M7/iQ
hVbKm0G7VnC/E++Dg1fHGsqXYdA/UGPpvsiyYDSdDhHScdPxiHnenVNSYFLe4GYu
UNGWbz5AWAOJBPU70qTWn+Howuw659gtivsqeUrQRrhAEyMNqE19mvomc9PJIu8I
rQA2agFDiEVD7oK00blVb6eviDI8t6oOJf6m8wl/8xwbcmBspbCMXn1+TCn8IihX
PAiUDWzPIbdsJp5EGr5tt6FLBuQn+ZEXteptLpuB5o+TIL11Mansi8FzEUNFlkq7
7pf3tTD2+2tEHmnB0JahCiv0vnEaP8zq2WD+pWcYXD3pQPWAEvQDVLUKdk9m43w7
uHLm/R9iRyQoIH9DxtFdkXQrGNJE6b28t8PRo1Gg0YmzLJ10c/tWmnEDoYjmVWgK
5KJVaxDDoS+n/PmKhWX25JpUAGjwL1YXnCbCPqdKOg5zQxWQ+aWI+pMx2SRmyR1Q
BTJUMWr3YwxCsRJqic4Ar/J4/5Hv3NnKqsz8nXozNDpBeUYQAVbwVlDkYf6paYF8
OGh06fYXLcp9XpUdabWv6yD5WNU3DTapg9pFmAUJJaEUB6MskyZDm1brPXXop7Kh
6qRkPTZ3rLd5/cMah0jPQpv8iR+f8jWsk9hXMsKy1gIopaxegcEHHszPnprZGNlK
Kv7MdzOP0UWXgy3Kn/+HjH+G8VGYycAX5A6U6ScaqfOnvHcMaTl3pBInQ+HNmT+O
QMKx0AImYlTlMXTFCbDE5jeetEcU46cetcIbldWsAqCq+ben1l/yQTgs9ubQvObr
Te9+e9cg7VyotLQwrV3YiZowCbpsF8GH9t0TlEq+zZ8rWzzC8QAk4OZIjwbUPtfW
g7P09nRqdJ44HCtqheil9Mqwtwj3PXqqb/0UMa6nCo3CTAODxI1WnCCKDhDLQF7R
AqACIx9GeKPpNQThqPgPQGer0c3+ib1UZzY26RlXiPCRgamH9u5YZplrrVXWLrNW
8aimwMkjk+HcKKYPj2Eex5C7yo/fTcqcIFsLH/bk2cYjNjfvNwY0+3e+PkGXEolM
TZuYG7yvFBHjY2Ko4MmDQexJ4LKQ73XhnYo2Kzje4JC0mX9DEaq0jyQpZseVs3pk
ilFapF7FagdzHpwOY79DufdPiGAoQItIZs35cBuHaxjPy31ADIaQ9YVKvnX4/OS3
/FEhxW7CuU7TUqhDs7tNzJuCpC6kX0CoDGzFYIqGC21UM47Fd/JkzmZ2zQiASyZx
hjO6oxsugVbJ2CnmirJwkhX4HWt65Ac8OdPZD+deOIGQWD30zRBhI6C7LxK6e0D+
8Vm0/BcAmNcxx7tsmUh6ZY7HoobxNd8UlstM75eBiCrDP8ruQMynyU0+svcqqDGw
hUAiZLQlQbsJFA0FeP4yLYSQAb4Q9MTLcClPzuPTjxWjNNZIr6f6AyFWTqIWmUHz
CJpVP2fTXPjBtBxwyGdhq+nABDm1iiE3jtCKO0x9SRA8KS0VVENCsguWQn4fpHtv
k45fIq9mXfB+ZCmz6snzX1lZVIBssfHf6y3PQp3UM6Q3rCWiWSXJNVNxKvqQ1nmG
L14Ksd8TQva2IvvLz2294MsVmPd2LIPMaH3y1EdDAbZj3j8pxHqKXJTj312+xPFM
zL2JEGwLh3ynXp/jinr9de4aBTE1YpMZ9RZ4VF/SWHcR1oVRggjoNmFyDDJk3opk
l3957a66RD/RuYhskEbcr3FVSVPMNQM706uJ/wLXkhuD+E6gtWggeQgte/x+S7GQ
Ys9iMuliX1Yq48oyssu1P44cuALl5d0BxJ5hGXKoWXp8iBR2COUwNRjFchRDpTTP
xQyYIa2RmYs4Q37YT6hnJbSe48AvqJjZm2zy8NPkZ8X8W9K/P/8HmIAiNLsMM3P+
DSFgmXEJ8k9VKCp+o4jjBkft39XEx9Qz+pZJ7ajjlt8VMOtL+KjqzAux+xSG298n
e0kWTFyYoHAhr70O1i4oXzs2YYp588Xj6uU+OZCEJow4SsrRj4FihjXuO8MpC5CU
Pd4xm8nWSZKzVHFd+CCWP/CbW4OVKajwM/FrDtMTyB6RHwtybirfVdRCFdkLfJU7
F6yzoZduRzzzDj5vcozBUP3F275L/I0hQNOR4zyzhAtqsQqM+w4/CcyiYZCbYQGR
kkh+1knlLZFN2KOGvWGmVQx01I/Er+PXzJShBkgCfJXNrCniGgqemmogTT9LHw8w
/zrPBw//0drQ/6XxBUyJjSkWmiQu+QScLxV1gl3YQCa/ps1fnlv1WGW0JA1Ljed/
w51q6+LtjMrssnZu7rY31n76TbUVzHO1wXqxyvpdapVMHYRjAhn5zjqL/Ckw6Lkf
aqg9jgtUAKp4Ss/GardsF1/OMVqkTOnkgDLCwg60uN9R6izFQ2tU7yn9COUJN2gk
9u3CLfcMcqbmsMDen3p4w82wlu8QEQymSK0YeQAbrJw2uWhMFNvHDopUE63oqfVO
F8C8QJtRVT+15rywVNoR8c9Z3oxLMeC5HD/Tj5G2H7V+ESOJWVa6SuSAQTVrC7nY
gk0yNhov+VKEwOiQ8i6llrcvJsIrNAxwwFq3WqlFn0PeR5Q59HXhP5/y6t2ZvyLY
zUoRLChvDvIuCiUHZSL56QORGMjYYsM37T2p26H15dJOiNZKd4YoqzPHXAxSwG87
kAeW1Ld2AmX7QNTdKRmpgfsuyd9gESKKV/X+jSoXSIO1JJA1BxW0t2kp4YIWnzwh
TRRtxZQseSi4HIMhG9OAKFvEUzG8ZumO663ZE1IsGPmWyaXXnXll+b6dGaD9MQfD
AILd2cJJflCiUAG6pp3sDJzliiZ1N8+STrnhF9ouGzyabmj+7QV0NRCbjwAviSOL
aTYym8NpO2Pu00+te1b5II8abXiy4SjSE9klG3evvRPZEbK7jHksAzyeyBBvpH5l
4pDZTL7IFiyyumCu+enhiLEso5Sk+jTN9EdvabtvbB+EInZgWLg0t8PKd4er6Asf
7X0h3ImpeBROVCwpPJy1lMZBRbo/1UEz6z8X06ElkMcOJhSuRr8rWG6SEwFjHhNl
FT2MFLMEP9cP4wpzpVynRcv9qeEafxOTZq1w/aMRu0vc0lGoqWAZwN02oyF6TEak
m7PQHPu7fwC9nYkGct8MFcyukeQnfJNdUZSItqVP33YL3E2GP6tnNyL/7T53FuuQ
kI1PwM/j93UH/3lEPCC1jFQIXcvJKQiYk2ipOGqYRWofaY7JNUzenRu2fj3Pwmy2
3kk3XRS4ztBVSnRPaqVofTL8jPgEe+SHlJPtlf83Pv04MgW1pc+KqCb81xW57vNy
9KXf5/qq0dl/HauGul2jnkPpp0Ue2TLQcKaPnjIu0v5FLk3JOyCGkP+8wU9btiHa
f1peVOoAOWnp4j3Anl9uqwyUK/3yXib8BpKsMyRe9tJENzIqnZ7Yk2n721hAPg2F
e4N4ntNPIAOk43r2vuxVZ6UXfIaLyFJ2zqtczcjo/WeSZ51Fi1sHcWMh/SxwMPFn
I9J46bIaIj2F4yrD4Eq7cHv5QfLb221ikzog9AGYdv394z/QV+YrD5z9wxRAzbzJ
Ma3x9Fi6b/Usfb9ZQjTwLevb6obuxwqbiWG8EPTC0DP1sojtoh9BEwvX/XdHVPCq
Ye5p2DTzMnMNlkqfxpWZNtf8YWDEDWKoLX9TIsATmyqNFDuulMF7l2cI+ek2lIHN
DS3UAkFqiTKAfXlHL7bq3cYCiDOgSV5gJFGskHoXRQK2yZAuYdrpQ26dqXpwjQx4
cACFsMpnYDaz59tDHPpXRaftWr1h1zSU0jyjVmUEesqyfOWrc9ICtQz7kzqweoXp
cUmlcwZq1TMJplScVf9ShlfpytS99IjqxvpBvyK/x1c3XUhw4FzbEahEeDSZJxOc
jrFvgXOhK8LYRn/UGlmxXzxb7P4ubCeCtA4zx0py066DMX/SKut9bFFagUSRIbIb
WggoQJJ+LnfPfE6/HXgyvG8yHwR6xJRD46dCrNUtNxwqGoXCEuJEbkHfffYOcBSE
W9RVakGd7nFUJL8KYBV5EDliLOKUBU+wJ0GPF1cRZI+pLsbtTLYFnxOGeoyf4pgz
oT1JdP+APr6xAtal8xebnkGBQTbLZ15QXe79Ak4UNKdLQRsMXI1rOsxKHK0+yjXS
NRZRUJVajmlKNJs7xil7C0MoVevAHgn2y7Xqszy/2AKVChU3oqp2t6h4FmGILBGx
4jqxcbI+nycjSyhimuG/zxpH3RPB+8OZo+OzE11VS85tXdBC0pOzL9bRrysrSuzG
TAx3kZABx/3tvHkReq+2B52BgjBPfURhBaP8UQeTipX2Y2vQo3zlWTQE1MK4KTaJ
olz9ZnOflZk+1I2Ls31grjQaKQUFHSDvHJeicosnDUO+Uj/MiEnznJ7foKOzJipL
6TeIkeOwGQ7U3Xod8JkqWuoKhxIS+8Ktb3zJ9ZbA05O4Y93AiyJw2UaJyvVWWGHK
Zhk4A9BwsEC/jPl5Zc33F2xZstRUTGLMXENZ/AJOFa+8AaAL+Oj5sg+E9G5CBKnu
SM1VmLPefHTA9Wdp7mkReFQxF1MtXp6acqH6Y237zatlUpo77RMZi2tAU4J+dj+z
+eu8UVCyOwbaMdpuFMQxF8pWwKFfp3G5QMoNwP24CCYsMcKznaF1MDCCG83i9Srr
rsZcfZvTt3tqtl5vs2QBF4+q3BY6VW1BKystGA3bgoRL3IeHnCPRyPi2Hgu6K/3f
ZUhLm1Uo1wABsdl5HM9nXLnMPRqXIwcqjfzQRrM/6DwXl7YyZItzlk3wwtS4wBEj
gRqFgeCb5LD2CEGSNL7k0fJHKXmc7mVvqsi2ZZKMbyU+FqZaB9Pidqtw9DdXjs5K
LAt42Ws8OZgzPGCmxxx8o4Aa3P5uUmoAVyKXVlLSTDVF1MuwONKbaJCih+9OkOOO
4/TJ2hNO9q7+8q9wPYpdNGIDE1fHjePoqNhk4VSQkT02Pi0oH5SRvcllEbA59vm1
MoytB+FZLKzvNGozE+8GEyPtBt651gNZ57pVI5AnqOYR2KSCZ/kTFaHciRBMbtWA
Zm/zgtlB2FgEEzwuHk00QCetMMX8gk6BlvTDTeB2XZOORR0vT19eZc8JQhUhVLGY
vk7KZ2+2I3iKSOg2VEolFJU9sv3gFTW6IJCZEjYgMd6ixJVeke1IQnA0hWnBCQtf
okNXHtQh1HTdwqX+djwSCKJrE5RZ7R833LGHZ+2k8GB/t4gFaB1uM/Fiw+pVHLei
BIo4vZ8JQztyozyNPhC9AMqNu7QSrc4xxnKVfNbCxJ5hLKFalp/8UI1hwtDMz2mK
GpXEkMas4PUD9weg25h7fwSnBfa3m/sJsq41DJ0ioAZrwTxqGrYTAiu0vk0gJMSw
AEP91BTYe2iZj6ljjT/ZPFeTO8WAh3luhFkkG1Sna62QQK8Q8XQJa2yfEFPnirJ2
wldKHEVOi+28LuXaOnZ09by0GGDre1kJXrZqYiOhLvPMz4PmH7cwRgzQV23fptPb
Q7Dh7DyLB56+sDIXJyG4X1GGMFTvwMsE1GiyEXtI3iF67MoOTi3iEebckEWvJXXh
99ghvpV7ali+ePj8t3UB5xO1ETcgfk7blF0Ee5xi3ZJNUtuC/7WLNNI+aF8iXeAG
9md4RVq+VJXCjKLUUlFJEnTr3R+IEuo3zv7z6XdXwHQTv6Sg7TX9IzoCRwpF4Gh3
BHpVcsHdAKdpJJMM7hQRWvYz/jlWaC4vQ1HYlvcf2/7ohOjb1rv3fYXTwRxtAjIR
+EnKB1IM8scq+csOl6FCXTCSyzqgjYhGL0fuJPENABbTUBo+0ZwzHvmU0a3Ft7B/
2HwXhIROdxlllivrLVze6iPJ/aD8pFdUNE4DouVwuptAMIAPBqJOPNaWiPL3INgw
DEdU5ZII7Dgn9DMYqsLpuNCVlsqh5IOkbzZW0GalqS2/XNSqNh7ih8joTt9gvQV3
B1+JC3KeEpF0XonvotPIWPAKKjJobuN572D0ze79Itu7p+C7aCCgTcfzwwIwb35D
BVqys7rmAv5doluO9QeQRKOpgduGWDfsfitsMtQ8vQxLaDe0W3eJJagercNdilaD
1bNyBbCPSQpmkPtFczxk3bx85/JiHXuBkzzHJFFuuPdzK/cfq+2UkbZwo5os/eiB
IvQRPlcN5xLTJuiqAlK3IiwluFM6/Xa04uBNUN/f3eYRpm5zfZ9ceoBZbpV3HFhq
nztMeAuAr8C0ErcVop9rIY5IXwA+KIv8s3MXjv1/dDO1W5ZAnYfoxB9Q7nd/EB8m
Vu/qafZohN8TBjpJl2qhHTSNWK5fUMO3/JBUOv1KLRPg7JXzxROeGLmHzBKMXXIj
i1YJ5kwn3Xb6pz81w+qOTaunKZezN3houbY1LT3JhirqATiVzO8lfoyZhN315iTN
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BGu1whyEkbiQhF4L9jfJGc1+4URXNE8Xe1y45fUhC0uy/mohQn0QUywMBd2lecAh
uuenNx5c5qlP4eUkN6aAhXyIIxo2Etrcx1A533ETmauMT0xhVcRcvRrFplHx//GR
vNnK55DldjzMFKuuRX3NUojk+YVxqLC00y61CwzGnTplXf2BgmfCu+uRGEVc8ngN
C/rYrZsPfR70DK0NXBFLRAIXXhTbVUkqo2WOsZA+jXs6wcth88fc10Q6aygHp2gi
5p4BTXAjGJZh9Oh2pV+ku5hDND505hw6X7UljyinmMg5mi7x3L9Xok6k33uJcn61
XuQdFv20zBxrbotkChaCOA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1232 )
`pragma protect data_block
Hyx2koIJvL0TG2FTsiH3MIHK/ZBfM11vAhaOPVm5Vk7pDL+N9ofoitRKChY+WAmg
UipPpsDfWkSlpXrksAyN7QdKnHOVvX296BYmVLBoJdsyttttOmh2j59AR0GDLo9g
dqewxDz+1TzHsC+C0B4r6/0BipGewGlrJ3Pg0h+VB4/s9khSOTvgcxG7XuCHVE0G
Dc3qIVSwgIEXaXCmgpmaADD8vcdz67vult52UktrWZH/vFY9rT8D0jpbdV3W9c07
qwVqlQJJjNNYubJbIrkOyJY1R7wkgMo/ullZsuNglXBFOipgjIKy40KGLbzgyAzx
AyudJvSOxpKFiDnOshMI0fSWMcuS7UlaWB/sUOzf+xoKWobfR9GkAcrUBLbOKPPl
myVau9rXi5J4WrhRQu1bBqOeir9XXC2hVgCviomOXXjT0h4vKWs8/cOMvHUKSgmr
NCruzNJOGF7+3t3jLmhsYGyrR687dBBvptKX7HTkwaLwjtlRuDsKLNfwsOCTabM1
TziziD6IQWYo2Pof6u/9tpuqvRr1ZGmMbcZQ5mhQdssGB5aPtUT/a7lZNlbEda5P
LjbQ0zwwUn4QVfJMBAsw3je4A1w01c2uwijKGHgQ80q/eYIGJm4YV2iRkcuJ0bU/
56hH0aw1sVFHAoZxXVCZLeE3USf1Xc/Ixe3kbEppWc5UHR60jhmx4JzUDDlo03rF
S4A1CvqSzHS5DRwq7cEGd4K8uNwhjRHA6IL3Ozbd0jsg2KCEqK+dDwRWzhV3zUrK
ph/8HRbTyEr6cq9QluKjjphHjxIuLWPLtmnZrO4VhqrO/NpAxTuGuXAgmZwoSyrE
mRFYDMcECHgGNA03zvrHGLWwjdLjnlOVFAKIzc9ApzUn9ZhrqusL9qF0sdMGRPxr
A45XWbeHypJh6c056C+gHD0wZOFpBt0lMPlQ1WN/fvsEsycOf30RR4wc6o2qSXi4
P6Q2EC1LFxJUFsmwSS/guyGIHnAUWzPu1aucg3u0yuFR9xmVwRx+HnhihhfI8GMS
u48VS8Xb3LQK8srKKnf2+UnyH3GFrTlvVOaC1qrVyKm83QR1bZ0gAwH10TSwMfR2
KH7gHEuyDeU7YR5/Y13UC3A0ejSmQtWXhBU2bQXdxnUzFXj+eVhx7aAyoQ5YV8zg
S7G6267J0jTLGkfFRfVX/Xc3/RjYI6IEpGHdFrEwbDxLzka3LDFpN5X3LgLxEl/R
gtY2NSnFxlfHDqwGrhwr+DvlXYD+jBVNJw/rjmhqZ1hsviKf7HlqUjPW5B+dUAtL
zCDwRYLOVNjl7uX8Tis7cAlR0iORh56vIrT930fYx698UHkGgWuoGMnrJcNFgcuK
RIW7+iV6q/DFfw8QOmxqF7N5hVy+M8O142qsbFhTO7ozh1elPGGH2rasaq4gmX5M
0zUnccrytd7nr+HUjfICTvzrG8wDmsb/TjgfSqHSxg490Z0yse7sAivkjq57hsJY
clJgRNBh1Etv3ME0+lD3jqMS3eopVKEGp9/V+6P7gq1YS5tP/Zf9p8BMRrz+lvVr
j3nK0/Zxz7Z0IRKgHQqJV8elahjizuMsaiO+wJygFN8iL1JBKbPGIlJKEC7r2czk
53uxLImEWR3LTtoEuWWhkxTmwdX8Gh5JpLnPk9FcCxY=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
P0+ExW9d5VTaNPppflKf91GATgRWE3aHWp1QP2SyybT2BkHBtAcDG/qSsbonywws
w53R3ywIyqWyfzGPHB1OIiEpG8TEEaeLEf/R5/W+c6YyEagbJ1cciYTOP0cdRvxh
0qh68Urh+eyqB9m5nJtV8EkjfUvw8fdMFVSFnAf3epUjncUa/CpUtv5j9Qctu1Vx
0soboZGw5LpcdQM78hCYbIFxjj48gxGNn35oFysK5XjleNYmPScNFX1AOLM5AEEP
EUSFH7Ggfn23ZdESjIpKxnwnVItZe5s91Tw/mJ6vK49+g3s3sCBZKcD45tRID2Fz
OvQCMcLaJEeNkSYu8kL1JQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 12144 )
`pragma protect data_block
b73GgxyCzD7pg6aPusXRHpV1AFrNadbxXaCUwxlYjl1dy5dhQHPe0NRhHzyVL4pa
DD1DtFUPsLjoxOxaXhDkuAyjQDPHz4b/lnXAz6EuXygdcn7RPl9KKFyoO6okb+r0
5L1tCE0+i5lBx2HiVrd/3UArFei19M4liqnysEwVf9csK30AX1yPF6CxvxHU2LjY
3HjepDotVR4Njh0wZlcIDBYuw8i5nVWwJFywejEW0+4ZkIOvRnR0UHP9eCghfQi9
VnYMA0/6OyB+y1QTDCV3e5wOFHWOcq8TwAw9+qAUE1GQszd1uTBJ5UjJ3FHkv+Kx
+35xyX+biCMIeZsJm3bgbRjJ7TkrV5BqU0EU8fmpFW2Wx27comQW97DKiO4xnlMx
gSd+ZpsJBS5gMSAxxY8Dug6ThhTwYbcXcF1GYm/BKrQhkSUtT0VdtokD9OqxHfu9
6tpDRR8JJ/e4GpgVtQ//Z6ziQddEtoRdvu404bCQxlOaBJ+CVsQ6tT92ikeuZ5gZ
rkbt6cg5qFoJKEHg7hioKzm2VUQWzh6wYWA6vzQ0NcOl3O5RFaFcxguoQBj2+MFY
5lWrecc46BJ6NitM1EEcDIbC116biQMzZgFf29wX8iTmMONVZuU71dXkmO9aWSIj
1ipcMC1NXgwxF6mCVZG9PJ7nBL7PEn8lCNrNVDAan5aunfzSilP4Lb3zjc01e29f
urAAnmeo8urXj9L+isTmvGucwomV0jzkmQOCmNvvE+vNuKnuhZ3mdUH0A2sqyD/H
tsPWckYXrId53PBJ8zUAkgjHBEqBTYugmjDtADJ9QcRGFr4GgAYOw9WfiysjQOK3
puuT+oHdhbg/OdIw9xbqOmH1r9zyw+5Yk7gpxlBA9/R8/nXlzHrvwbBRfqEtjvgC
RkSOZVu0WmlJMbeTVTouvr4shgSz7m9Gok+zPOB1X93IaEEGjOZsJHynN4zx/yUq
3qzGwq9e7u/BN2lMBuw2wCEIqpqTKNigvxKjXTHvJW6Ud342mh8AifRzgFl3qXSP
oNErZxt6U0+MTPSPxsX44cR8Ig38iB9Xdwiml4df2RyGzFsyZiSTt23ShpkhAAfM
f+XLcogq6AqPjbFXmEGZoYwnNaVs7qcoFNZBM9a7j1VzrKwyXCX28uieWkuJZbe/
+sO2h2wQv4sPnRjw8nqTna7H6Qkhb52aX+Q+UfjNQyMpTIq3Z65eZ0thQfO9n7m4
60Hmli40tuSnA2ihSWfzW5ZrEwelEmM8EYJeukJGZuikZmY1JKrk/yNbcOVggN2Y
NJ24tcYKUSljWVb+qVgc5TgDbjENeBT1cxTxcTVZGiPOV/deSqam5AbnWQlGSn5m
RUpcbhLusUcCo7BsacaMcYuDBosdUSfAyjCjoDVOGGVsn9CEy6RHEVvDTPpGYuGT
u4HjKDFMBAsPSC/pbWi4v44wAP9i8NNGyF26FitNr8WhJsKkfiheCrSKNjM++NPl
gh8vzEqmkPUoM0swwX4oc61Ac11BlmNbu5uGYoHli4ZJOcu908pGsgtfYm0x42qI
dKHFZz2LWiogIH++b2VI5GZV2EG5MC+m06/z9f/NoMsU543yCCfbSkUfo9QddtAQ
WI+hueh0+L2Miii5JAHMGErvn2Wakm/59kr9uGx/SsYuWNA0SDUoQwEs7t6Enuf+
w7zsZxNUj/gmLQ8bguPrAgpJD1eswLo0vBlKC34X/YrruFxqWqwhrd85JusZskey
tVPuNyGx55m3kZ4V8IJ7gTSrjGAilYiG03EO9mhfG/BUbZc4QQDB1TqU9HdJVik5
qnXVOgaejfQLb5V7XBx40KOSPEMPLs+n7Kz4Pq7d7yM4tOMKUl6NTqFUgmIm5NER
/Q334/8dV7MlBgX2srbmxn0MrXckZMkDdIg1yHfgBzJ+H8iQYKhIbZUF/1lwWbCl
RaUny9Fgxw8KqT982KLU3Gklp9+3HCuJOitl5SUTF6C13VFFcTmF6jFd56djLrJh
dqT/47c9zLkCW974FQNFurz9phPDWVnOcCv1W7t/w6tRge2pI7gBH78o8zX0E/wF
nAp6UxR1clUmZAwtyUPNiFx92wiLv36OWKiQZ5jKUQAwdmNidbwRbAFKbVKbXtC9
ic1zmD5TtVgBm4BAMK9pU+SEKeI/3MEx405HnoeX53woPYMEWougAooqhUXAH+Q3
DB3Kz68sJiFWZq6L3orNC51t8MfGJV/UOCTSr5Jxi19EDcSeHzmqDbSNh0twDDML
cwc1qxzG/h/S3W/z0C/8JVJKFZ954ZrkFEUke3LDfIqam4qhBXtgjh78fWoal1No
EnVIs/jpL2fcuRwHvj6BTimSV+Y6xu7C7/wGz0FaVzB3ruCaWs7U9QXquE30j4us
0Nngw1vKluhK71txZOWBmcbzLGqyWe1Q00tmeyw2YbO0FkeygMXD4XX8lv/Vgcwv
27PJxsSpI1Ebe/UUgPZHX4/sI6ljsu5WFLKgqCbLkENEW2efr942oArSMTk6iA/F
n13Ncgua90Gp6WNhdgUjbZAdF2X9FILMY0wYE6J7U8FpE5uCpgdO+XaRHv4rb5b/
i4SKnQfWOhzX5fgziq5/EK6WU3Ep94yHCoDRxe0MXS3WozVVBFmiWHjmqDn3D8Fl
4fQ+pR6TDyhNYCrCoNjvD8QvmvmyQRBv/vnCJmVsCB1mtQLbXk0nrwzZYqtSVgGc
cnF0vgWDDbZJAuAOisfReMq1pnEoCJC4VvFQP5VRjfbl3o6R9kULkUWdHbQbSBcu
4+pDKh4+PoNEMdUww5rYtfA92qMQMELU6fb3Syme2y4M9pkPl3xsfSf1YAFiLWTX
ahehxzOrR1d/eiJv8+4LJRxEzH3HCNRUd9F0+pbT66TbXLOLYUQVysQb03UfchId
cghBJtoFDJog+AFQMlC+JiTVEJchQdRg3FSfMVEhELKru/KAKHK2AjY9iIe5X8gI
4CXxUIQP1jUcVq58h1FoVLQYeFYnBBB43thdZYaFjhN/jXeQYi3lLwn3mqvj5Acg
UQVU+kXtgkIoa99ezT2Vvf2M2isAXIoS9HDly3QGyRjF0El37z0iRvkZi6tXB9hw
yOqhvch2WtTUr2nXhTxjXKNOUuCOlf8X1VrfHjwYaYZWvhXqoqhx3sYACGBfUT3F
wCHi09iMZWb8PmnbfaRisR4eubmKS6yKg81ZY7zL54yc7Wfv6xncyvBJBRjbCfma
aHO0Qyh7ph+EHHLVo3ET50FZwmjVWWA2Y1nU2QWcYP0TdkXLInymOEI2pELp9egz
FwmyqrbB74tdFbMqCesbTf+aN0Qf+p1sADD5JZVeVGvIFcCIm5QhnfKx6J3yOxXW
Czrd/7l4sOPrPOEpUSkYuiTCo3u0MT8+WYxXe8M3r0vIXclzI9K7Cd64ifB/TIIw
BSYoW/rZ5vJXchWwv1eh6TK8G45U3aFJ2U+Du8MtXWjK3rMnzZ70j8+aOUNiWi2o
RDJ8tI3XgOPm7a3RnXow83R4CE2C9S++Omf35aFW3D41hKQhpk71jbcEceOCJSWp
fl5/uMyDbAOfiJEOTjQB7QD8rMeZ8u2Ex/dnhiYX8X5GlJKi9fETJsgopkjCeUfs
4KHmIcaowO+BvBwWjux/jD2IeHx1pKAQT39GqmdctT4i8whToWdAU3c7WTLud7Tr
qvNh++Zhliq3Ki9S9g8uOutLSi/quLv16nsJvgR5lDa7cDUHYFbHzVNWNM3QYkpj
848O48uP8lYx+VBqkWFfXtX4BWhuN8SGuvoenbeZ+KprxeyAoyPr9PzaSNRItavr
kmVgbG3PdeKkV27HEeilgBu+/Btz6WSBj1ifUr2XUzB/QyNwFOlf6899KcfE7eBm
gt5hTObFiyNEWRx6bDKPIfe99EyNBJQYT3Yy0dl80Vmcuk27ibQSHI42vSDemCqh
mnuQUyqxzDV5sgVZPDfxbg3PgvDJ+fWcCHdDeVYn+oqOaWtlTQzzkqvJ3rVajk6J
N3i4e7uKzf9TffryL9bvESdSikaHuG4Lw3rkMXe6xTQ1ATSy9bt/LRnFKCqKhuWV
iTDgCfpa56YOn8Wce5qOdmQIqB9n1A1l5MYY4aAkkm3WvTa7aFS8+6ow92OGWCw6
AnKisDoR9PPPEHv1odye8WHQkrdbTun4xXlWLBqgZfBL0BFaB1jGERxicAizN5P6
3v6VNQClOeNtKqY19nRSci3z+r9ui5Wr9+zCsgvgqlWmPKhIMOVyiLGr5wK5aJLb
tz22QibgMqzcC7doy9kEHVWHFjjIqiMeG35qftO6dOW06CnVtOFhEZI7A/K1HFZk
dvl6cxynMuFCjbZJOHJkU4ubAyaPaNehQBXH+JEKwKjlnAMUJxu/VhSDZrrzin87
TcX+eO/db28s4craNVGNdiS7SLEOF3/uQv239jedkHv6K4E7OgWDZh00+qPUoWSv
xAIBShdlSTAooNvUWpxEzn/Gxmq7pe6SEZe66tPs4lA6ExSOGgpqffDm+6WJTVYt
3oMVySPBfiVRMNu5BrkxQHfhJlODnXZpMuvT39QCdlqAMC/FPmEl69Xk6rxlwQ6O
9ZP1I5rudFOWTTpVx0/4lhVUVH85ie0Bfy963F3eRlTVGlrUHDPJadCmF5FXXQLR
EJf/psvml4AtKfy05IYQtGmr/JFRijDziWZY3bnSL5xBibB2A5wwG+LEo18iN+xc
UPTFlA1nvaKUmdo557HYmW6Tudx79fXvJhFDk46Qpq970c8YnLF3OZGTxc8yoUeP
6hDB7+n81LSOlx2nYNzedEwe8mSvV1PzDqkr/9ByR3JIAuSPMbTegwgoPjVmwUmc
cPrQ92FoG4sa+vqj6AOnlGy6Iwd8fVhbGK7Nyh7K3CBT0Ruawm14ryt154ji1pkX
ZyvFGxeEKvEIaQhCyU52Z6rhmVSWndsyh1dLS+U8lOrvp4XiOEkgzKP2M31vSTtH
bNYbvV6ZLObXQYNSrUD8GSH1ftFvvpkBMs9Eodd9iUkEMdFSLCRCYYRQZ33eMCZc
Ila9VJrKxkHhIna6OoksC7BkU1pAzL87Vi24ZG1gCQvfh0nsccPqEYK1UX6imyzZ
yuDL9WOjX1wQKNvSgntfZdApej79sFIYv7Ae2oqwMeceMvJSSFn6ZWlHMuMhaM7G
Yg+ls8/j/905MCpBMchzLDjctQ+YoJwl5WpoB8wc7asP2IParS96Swd4TJ0MgDU4
6RZXuBvwVHZFBh1S4JZsEmQlk2Wh0hZbq77/CnWjUEVQlIW7c+mnk2fnf626Fwpp
yCECI4naHUrElbSPrI4YvPNwme8gk8PTfXAikqAq2aAKDnA8Yx5yGyk+a2wb29ec
94glOn+SXERYhlvfTfdmDp6ybVYQD76Z+FOWvffqJssETVfy4Q9Z2bNXf4UeC8fy
ASZRbIchlvRU/gW72+gZESR3g/G79vQwT4CsVpnSIgYAJX2D+GV2MEsrF7RI40LG
fAMbKN2SVu8tP5PUCDNyQaqGVTdNQhdH0p/OPWdoOvrej6lqY25ifUTM6iOWFdMp
VK0KN+jzQm7G30I2kvGAGiGtA42ABqtHUvQ8Kfb6Q4NPX7Iyghsn5SDmjXUNJJZ6
nH9jbro4bPtCicli21u0M7tb1URP4pysD7gyxm5ZNYXVUj8KQZz5Vs6mJNfxGyWF
9Q2eQcmYkigSeTqQVrF5G05NpBQCckFvIapHMyk1XcNrJBYUWUsNTxhdieLgcRiG
Yxsn43J+K10tiDhHVwryR3ozhLKNymfTbKVidP5LSQcEvzMfbOYECfVGI5XuHeGC
1eZZTBNPJT7bNExsaJ5tJx8SAokbqJoKp9bzAV2CTD3Jt3tkbtFdy0hSxuc4JE+x
T9ov8rKuxkklh10WpNJAT2PeSWQpNi7ypFpi/08DiOgYaumOMuuTaTI52o82x+lO
/33igoxPAFaeGVD4PuaGztC28PRHenIESmAnzzqXWta7bbjMTym+pmh2d6+/ggUi
WthAkcpacwr/5CwO8TQykf73UR4bfb4G2X2iTpWVexc/XIZKkPEESKQXV2j4ETKD
i6ZTL5Z5ZgrhLbR6s7XWZmVlCBVh4knbmy8Xz2m5EwF/rPjeWPr4x5fnY1W53Ckk
tBTbaKtq1R+Bclxqy0VuVnpvtSquOp8KgDSU1YdoXH4VYhu2j30LWMi7KnmXUCMH
JPmyTSG00qChhTENG0eWXI2lgL315LpMrUui4VowM4b6UskLm8YG9hpB0i1MWQKz
ysVbsff8+0lp4aRkwuo1xi3on8nF19mDoh+TBTT3EuvJVjVrmRi8vxQ5VNl4LTs8
uBQH81v4kp0pCFm+XUIWH73XaSZeWYXzKZmXb053AMLFCff5mk6MSjG+jOpFfAvN
gMI6NGWFGAMCQRodt18mEkdXyjF6bv53YCwqJAI78DrJMrvK37ArR7DAj6XVwrmq
RY9i4gtDR+FUHEXeJm0YthEMP4Rkfdd59H+xzmuDOwFbR6rbRYUHpu+PWMBaaOZ+
Bi5Wey1RFJtGc2vOC2WoMCqZKxyVQ1n8aQUMnGVJ0iaWja5FaIRXVrRzZDVnFhDj
ALmZhHQmvleglvutI5sdkL4Q7A0H4iuKnxXlW7HYdGk5J2HpMw4ia76UXi0LsGzt
exgeqHFM/FvVp7JhMGnXUfkxMSksPpYvVEhBnmgj6q3lBTcw/HLoSma4WDDHHlae
94Ke2ZHY7VIYE2qVmdOeFNhr/Av94963zqXxH8leW4OhS7FPUtFIeYLmfh/TZ0AV
tarI/QaanCXX/B0CGTkTTF3n+nD92HgWtFJd6w8KwaWVy4pyynkxY6PreqxBpxah
xvm5tP5qfPtEYfs/lbfV0Ppg/liHJKNQvFVzvV8t8jVl9qbKBzJI7OieKjMDNkCV
4E2g8N4+9+BtWp4nH/d+Kkyw9FphLTXKJcawjkzRBeF3UtPRsR1iyuTqAl3Ar/og
xasv6NzKLTZ7t79zmHO9JyA0oTtSDTEPwm96WiW/HKYcgJSlLitmGYaHbzckCk6t
oSZzaoBcSV0NxlL+Ob0whwwvjIc6lIm6iaGFfpdsAjGyb4UcdQftgYrK3+cjoqb6
I25ihATv1qBTjw+w2xSAnvylDusXLL9jKLFK0xSNWCd3Dokw2rqUXvCa+hYmbLeF
8ENJcQvitAtZ8IeYmEBtTGNyaK7983YRoc+P52hgpP7tZYNGRVfx43aAbpa71a3I
QZr07VkqCDfe2NMEd56jXHSo6DIJcxvv5g8515Vcnjr/Dcx6ohmuSzbj7QOtwr7h
uX/lfp2mC1KKJAS3U6HAMA2ANu4u74fapqpAUppp7RwQx071LiQB0HxhjHv4SMh/
rzueawEOJ/P6Vb+1ZIA194w4strSJKQqww1Is9W9L0jokKgZHbGXtWLI2G5Mm2XD
OHSHT9WeFMWKFgwcFwmV+Uywx9TzdEGGAu4CeRPmxMVHewSIcvuwc/E4XS7UTGwv
WXXQNA1Mo0bZOlMvmcsg3hZFVy0IxLJZf9xn7fle5raYOM+Pgq1v843xuyS/mf0n
xihlKuGRJkaJvG1MQc0Qx8XE7zne34Uq6cZWkfwt5jDrVxFAOEfZ9a4EP8k5Ps0B
jK5MsPEQfRzZ6K6pSvz2vauBJ6uuZkwjZrPL/qCkXP13bGndf435oDRjaUpRYsUL
P2r6kAgSqMasutdREEpIvZklp2dpbzr6wRyM63BJCyNQNQF7j8ILqEm37JKk3JEj
ZUl3PKRuhDaHKEpNdtz/GRVjr4A0wMr97pW5fZN/zjE8z/PAxSJp+IbeF3lx58/Z
YM53RtYlEoG/naRC1S2H+G53s5F3Khyh8DpQODVhspWLP6IRCuAWVMeHbHTjozQh
ocUO6ZL9PfCwK6TqZanBA1R+UoqZkAekEo3i75Chxy/yAdUA+9G3woyEO5tsgCTo
Qhz5lkWAmkNCKAdwtgYqYcso9K38r/9TDwHVO5UpHctFcL/+RUguA65PuTAtQVHF
Rsxd7CxB0C0ZaXa08bWImv9yXZjkIAIyCADEkAFFFPpGOLsBAzSBYkesDOWjlmsp
YZXB+Eq3K4b6NOKJrLe9z6wnZ6HxvSSmOXYjN5yZxeNSQtvuiRB1XnoDHFZ/Sf9k
8D3zCy9x6NYfzhJhFbaTr8Q+ghyPeV3uiPMDgiraRG/hnCRF7pwXxqPK+qInqTMY
cyAf0qPPFNXPjiyBbDoFGZnQp3ngY+JBdq7EyilXldATxkoQdd+ko1RdPwTlnlHP
Y+88xQXSlxKDrxVN9QZMNjcquGf8b6Z9aZDUfWNUKuE/DU+skNzjyDipibQLDfJe
Zj0ONcC84NcuzaoMKwbem7ZM9RVB6NvigRfnfx/x1h2EfjR23bT3mM2NRFd3Eidd
Od+OmSnUdmKEjzMvsK7kSzMTn1f496svxCsxOoNuCuCqVeh3H7Of4O0wIdtzR4Mu
0PJ7KsjNEDlNt6/+e6sBSNVyzGxE3S5eiAqHJ0XI1Y+O8iPffZkQBVRDE2sjuBUD
ZxSpFWCW8xiz02kUtSNK/Fzx7onr6wRZe110mCFry8XNOQhTVOtycUDWBrt/cz9R
Il1IB/vMwIpsUShDgfxXAKwrh6t1QauHZRWM5/cs1oCZ81bCEs8Z+w2oMxjUmZ1m
NUu9CSJr7eqrmmbgHKI+bBCrDaZVKr60usb3WP/OsxRHovrS6ak4J1A4Mib7Anz4
4Xl03A4XUNZucdFong9fi9PgJVMwKPkp+KmHoXVMFD63Tnheu0nx/DSSUuGzX1vR
5mWjz1e6ELZEVqt6PwoKTwfPke4QNj3Ev3jzAa+6kLkl64w0niz4TeFApVoTVWZS
NNUnjpDibH+G6muvBSf0HiZZhIRbtIz38d+3ngMzLFZdFnHFzl2AYMwHSP4u+INm
R9enwnRw8bFzSnvadeQz6qXJdwW87EIKMOqGco5u63Gxb8qNShBUaduGNMTlAAo1
FxN37uFX5S9jg6YvS0/7xNBLem2ZWab7Z4h6n5sQZbK4N7KEDiZuGtGpJe3pGzod
DepzZQL7jon+gat2ggX8KMR09wP/WlF8GVl5/JcmPpE+25PySpZX0yTQOOjIT9vM
lxE0IvTYFzLPBxsncCQf4nKO8lAcfLczxsSVW/FuZFqIhPxnUScOC1Su8WDSgbK/
NmsELY3l9YBRFZewWNdGaPLTHg2I0I0zpt+kNX9FT5c0kzRcaHa8wbra+iNRlHhw
rtRxoZbwKTEQiCbdMH54ylSPm7Oo/UkszcYclD0A2NPmFsCjEwHlXzsSYB/VXxsp
hi5V3VAam3DgVn1BaHHpmwLHJ6SNixq/wBb/RRnUOW3Uh+S8a5ovoNv4irDrY9gR
3Fw1qyHkPet4oy6hbuHX1vGQAf+XUdEQEALOA/yGamtuuuM+IS8AvtFr/Dvb6OHB
rJhyQMOlDZaf3yh7PXIO8z86xPFW7I5mx2BxsEhuuXPzuKVJAGXZIp7+lf8ox19g
uc7FebD8Sk5zbf5rOrMT/I1mBRazRtXKlC3iAqTJeCTIqcrH8+QedALK7igI1kyk
Azim4dWBtVayMY7NqzEG339yMkxT0OpTXO4PVi70Z5Z+hfpefZaDJ9EuLLgfHHiv
2tLJ9YAF1wIBj9x/xeZkr9TksRtUMqSDO6zAIblbs7FMdd9mugxj14W36TZcXIQQ
bGw6P6059OPq/B0MZfac6ahJD/W/Kg+Zv8sM7pnQvAxHiKSfuwOMktB4Zdd7noQd
wNZukkLcoMKBT3fH6CbAcuLk8mROIn0ZNX9OdFE0BKekxd7Fd/xoAzi+L2yNRQdb
Nlnhb5JelMriFgAoydvGyqgcfpKphny4W08WMNb9t4/JfVu4FSR7uAlVAt7AH4Zl
je1GrrrTgeJBAu84BZ9GicxeuOMUotDAFUdlUJsXkyJE7l02tm1XefS6bZVzNadU
ZoET4Ez9DflxqGl3u3M0z7BeFoUh66HtYbYxnSkzH0RhLX3LcH8lLsGR3GXmWoJE
6e7BfVEmkHDvrPwLN+4zH++xGGpOvH+cDzMtHxZQrS/xDNqSZZey1Nc9qLDLcYne
qClacPqHgnCuACNcW4zgjPwSqzZ0CX9fwBkD1s1l7XXS2mXPck1T+lxB0SV3nH3r
m5a/jSINeMbZ2fQuAuWzTH85gWfkahuYaruzb10PSjxRbg7m9BG6DK+nJamKvxFh
A+dId0VUjJLRqRqE0dVzP1zRS8lJ6FxEbJabqVKiMoimrQ7DtyAXinH/9uT3ZyvP
qBh+h+hnatxKoO6QPAsb1gEWAL6tgncOCntNnQSy8kLYSqQRph2gzEOLzoZJNGsY
6MwZhwS7TJitqfic+upeHuAj/aNt9iUA5mN2zR8XeShhpTjbWYeZqSVoxM28ab5o
dbATose/b2mFb+suFNp+WcZkgaAPhDJpPRCKDu+9CdXEbpvY/CWx4D4DilcZMo5G
p0berYvWiUHQbPnJ2cpGBIhSieRPiiR023GdkvsNQahOh5Eob+BBDgio4WYCitog
d0wXjU4Wn1PnKAo3OBfziD7PMUv1eFtg1H/efb1wLLf2aVeomTZCLXdNyr23zZc/
TVNEuI37zV8yUkd+CnC1QB0oaxtZKfU37wl4ZQi/RrfahwucSKjxL/4l74r2RJAg
dtaITkcmBKO/O+kcG+cLdJR49YiI3sVcpO/XtkZ0F5evtavuPuTa8Bpy46xe1Sdi
f1ndyBlsbNa6t+x+UvrP1MFwvU/CMMYxgTBV3EHYCMSwjEecxemW651/Ypii97OM
o52q84ukZMjf68e38Bv9uvuFqT9jAruHzn1a3hO0zq4f2cPAb7eTIuIEvPJDsvQd
1p5lPGIBVhqnr6BY9lg3tJqD7c8PkVCPNTByL/IWPiCcvwP8SzRYwcWm4eZ6JVrO
gF4ss+K3XqifmGlgjEDlaj4HQcfC1ddWc0bmk6TX7B0b8rhYWjT4Fqru83NNuZXK
HSP2PPKHFV05habJkZUzlaDlGeanb/DmeLhnkmAWhndICPlZ6dSlso7GGN/5HKgK
STI/J8aN0e5PwkyMB1dHYd8PT4dEfT3KNDAnq6SACgR5dydGi8rtihmEo3HTKxEJ
BjnfZEzRfUQE4yrAY1+rqrdU6rd+2RbR2V6SiPe1mw+XGr0ihJ2xYVhFuWK6QMaY
KXSutP9wsHOhIHK3QFDdk9qwWzxNVE80VlZ04SoeOZgJhADKelwLoXcih8FKFCYn
n2OrxOKkwaaWUQh5c/yV2Ss7LmGaCdN8LNyNQJ7Abbmo2yW7yeg3pGRhLwr8lBIA
BscCB7oL0rmffgZp6VkSkuX70yVZiGmwbFZvAOZvhmYZiDquAYJt5ogfruIxDFIm
nh/cXBhY+K9TNClbc7elvtHbk6tFe2fpXs6dyjqVl1rhnVp9Uczd1vj623AffwRp
cZY00kRKEhuz4SY4TQeTcmkAtlXpoO18/HPiP9rhk86CefO3EOUd+kk5uvWYGqgq
NvK+n2IaqCGQxX+pDpQGgggXN4Y+OW3MUM7yXZZ7JMSBanIxqFo4hN8U/hN52e32
pM1pSFbxIFBPxnfL2u0qqDndGKBUILWE7tttNNE7or9ubJOdo9l86A06ldKyYszA
xLz1weTwSr16SLJ7lh8PnnQ1tzH3uIo1Y6/lC3sLCX+pcKhziDcNTONEEzLi64rB
rtkYYoVz68F4YGLokDYK3Qi3Yb1yRzEaoxbiGo6OfG6g66/2xl/KduRjS9CJiAGS
CHD8CbFgdP6bVRmkdkKLjSGXplwuHG6IMRhJDpRvj3xMKeCNuZtCWS5hg2gINFfS
rLApoIJjMJBNjJ3xnxyYHSNWUcquK18JDAOvvh5OAs0DAt44ZQiA3wV9V1UfWbl0
U5Uagg6nZ5nVSy8DxNXEKALm6Ss0dxeqkYewBiv+jWZHxEHRE8YnwFNW0KzoITkC
GwSlpAI9d+7BYlMC2aJwcbmKA9lDzQFcVE04Vp8GqOec/REH1O+mdnPmba8UilVO
do51BLWDgM5cTHqGqMDsCVcTLoznyhRMBk1Wvc9flzq49W2cNrACad11I2jZsyR1
Fn1nZAMxZAyyax5+E9Bw/5ayulrfBVwUwfvy+HTcgY+SSE75dAzctG48hDUgsYWj
g5bdn7R34K8oU1/7f9rFFRqCNq8XM6w3nf9cJGM1+45/vKU8U1bDKARdduCT7cFT
Xs5jlUskR83KbH6sy/uEHVMCDnt+OecJUZnoTxFtLr7VE/i4NECA6/u3f1jjrA57
sRzfJXdYvUTrz6cSVKdDJBHAeD0TbyUXPiYESb4TloBVrHB+PV442A7HJV/nZi4z
CVSgk2NBF15FIEvVZNArpQD6CGQiJ1wYxVXNayv5j92RwgFTvpPi6XBdZNtYMVbD
y3aE4axthP/Z9BebfnCrtHKOiyuegTBNQZA/e7Wc9Zi0rtqcthDvdvAIMcOGAiqF
bPCP1qXEYGLs04DC7sB4i3I90UxGADn3fuBRiTu0rFZnA9HvJFk0H9c5Mve50c0o
IN6eulDCR9JJU4JRCER8dJii3keT9iviP5vml7ytWsExzs1Nz4h+AuxbkHrWU/4/
xED8DAT6wfTth1XNiOlrMYbBfhSi9euQGFrviiFzK/Sszl3xx2ASJdze4Gci87td
xMM1PeC2TkJlHbqjkwSgYA29ISRmIkqEUN5zxr6DH/DiZIkv28oEklSfJCZ//sHX
hNTT9LmiPrNW7fInuvvOqBYOykn3ihV6xad1yuaKcUx9ug3NkV3kKrSgivmdE/qf
Py7mEi5NHt4bwLQ1CvcBtHkrWPhuaKHDq++Q9zc7GPa3+1neQX3sX3bwR79gMLFf
1Vwd2ZFzkLoFIrqBdYciYOdz+ZdG0MXd6h3nznFs1gU0JCclWNPf5nb0Dg6v9Pxq
x0wOCwMAgxfenPdGB/6Qj8QEN2LBF8HjxIxLr7jxva0o+Z1DRNH9miC0Ij+b6dgZ
qDP+O6+75WiU6Phdks5v5y1xtxDhewJ2+FVKzAZC46h2dGhgNedRloPoaPEnTWox
R+PzILRQkNO2x2PvhOW6o25xuLG7wknc2rMOI3awibVNQ2ZoU8nZJPSjDTlYWUh2
W+pPnwPs6zPP0uMF0vf7rL4bM2zPljlRpx2CDwFiLDN065JqsbkzbSpvBNEsiUq2
3A5T47jf2MHt89AdNNZwRcb6Erot+wbM8ZiK/7MC3XkJacz9p12g1JMsxnTheqB6
OS06CZV4hZWt6PID6meWalSV2Vn0pGI4i2RvNuay/8V908eScNWFreBzUiSMDbjp
uppe90Q2Vup/sR0iG52efxpOtWQaE3NSUDRvSt2ogxsI+KH+S8mb2ctsjOSi9k+X
y3/c9FCBN/EtXfvj2/vJiiFpyy/11RH/7FdhWv/v8AmNJf1BF7ZhOjNWBoVw4SkO
vum2rGSpM4Tq63RAYrLEdJZBHedpgcjBUPrxNK8lmgeGX/BokCISgJpkUBocnSHv
bRGxzjf6eSAiD9gHddxa1aDP7RMdJ2lHLJc+uoOKyJCId+LSru7o4tNHAKStmpHx
4n5sn1Foz4WSfkJZQNbKZ5yv6mlaE6EWMcYzU6iAkxesV9SwkSwHsYSL2A5PjTL8
sI0a+wzLgT4qqJTdjmh7u0fEeWIzvodXafCZrqmfkP+qIJa78xv4jhZFoTVcWSRZ
Gv5c8L5y1IinEhsqi3oNEp8cxN6yRFJmWF+G6c1rRoWlw8b61+95dhfxM5/sBZr4
9poYj5+sPP36tgtYayoQ8Hz2OCeUJSBnqBXtPfYJb3myRaq+7TSpUOAJljgESouL
PohdhkRD4Q3WW2Rxq+g/UxN702dVbBcE4RkI31nsIdhM9QGBc/cop5LLd9OSq2Xg
Y9IbQQ2f+prbR/ua/SDa4w6XycJ37RTgJZ4/+X4hEX44RWSXaLPYd59KkyRkIb2b
APunbJQooIYa3macbx5K8gm4rkCoLyYKnyNdDulT2AYxHJDzImykU9mfecH9dCVZ
IM4hR+v5YXqic5WY2nFe1LeGf1ZOIZ50fAwehSAneOYoKsMDAyirzBVEN1F3FAJ+
8EM5Y4/Y0tqtNCByNV2emkTgVr/sQd+n2ohOovRyGREhiUW1PDVPRVs9mPKKtfea
cLh73bUkLbOpek7qKaIOm3GsLhSNFXBmLXhERogcUKMOtjjO04LLPHY+zgeV6ycc
gMKnZ8Mo0q0hhnDAdBWzaUcVVKEgjlyeIHJwJ/dcfjQeqjOFgUqn71VU+P+EXXO+
ZEZaFK/Cl6jZHa9IrssS0nSBe1BWisZZUFyBKGFuYJ28m/iJuhtSwyYUomneQ2kX
AZi2I4HxfEarCiLAZUsZMPWewlTc3u2Brlt9tLJ/iKSkK4gslFnONpc/OL6BRyHK
0QiA1BSciLAr9TApOO4hlGHzcTtFhivvfEfi1PSnF7LOx3lwrtRTLX25nvVHX71w
3iXGXPvzTz7Z5JvXWONGAPag59hyOn4mv7/6lHq2XUKBH5d4Gdh8Z8vur6mHppdg
fzh9B33m+fUyPjk9SdihV5pPwlWzdHEOwjdNfWmai25k4tn6/5woA31A8zFDscGs
aOI1fO0IDaHLUKZORayZXSKrayyYPwhOfC00hRb/SFkRJ951UXjGaq0fZDm8vmW2
XQehk+ANsorrSazSy22Ys1Cup4Wbyt5VQ32Qu511F718nWNxUFKzMssURWjZDJsb
sI6d4Ac9d7315rCi72J8rbSestpsrY9I0Ovu5fvrhfdx8uVJ/l1XToa8OGokVfKq
y3UFN2jv3AC/LmDKcnkeboIJXcDL8TpaHbhN2vWAy8rwXluQ9m0ndqxuj/5FwfY9
hiQjCHguOUPahwssoEv4i7P4UcekSSZAjueMHnHUw27PgfJcNX9DAFns5Pg2h1gH
haONKR/wMnG+k0UzHWtWlLgX7TLBgjQUv2xSPfgneGSNuWLjfgRgggzue6CQtP7y
ni+Gxvr7UcDkMxp+vCzhV0gRmK14+Ufp7RuWTHVCZymvXpN40QD//uC1GJpnYIHb
80SMAFHRg7gWTeJpgdWRd4DKez8jPbsYvsKLvE0IVKIw/POJUREZkBKc7k26yUjQ
k/cUe6Tj5u7Io32SHRlvOT72MZUXiYJlXuqIntffc0LQ2jX9gqFVyC+sGh5Hku8b
lzelWxpZnYkX+8NRl/x91F5ldt2jLDOXZ6rBAQlyxPq0LOccoGcxs3h9jzytMgJB
ZoIzP2YDFDU+QywtADHnQzc+RAHAWqrQ0e9dMQh/W84t7vDPL4+3JcgyWH4x2HOs
7qur/m0BdcfcgvMuux45iibZwrxiNDJb3jj2V3qENgE/ZHBYQEvVqwCvdO37jCtR
wIQHxQiteVU4F1bmbNi0e5yMgaorWtsWkNFRncb9gMM/GhATWhNt2o72eBmtamnK
3yae1LwTxsrUWaT9w/2cn0lUUTyfKCazWHE8mnyEw/pWfuZEtnxrJsfqdeTF1RwW
apMlL8A6z3k3yazZ2vqlBYOmEBtfnhRCBbSXRQHD2Y+LeRDXob2h1D7KS1YHvHQV
EYkcQdAIqug/9fvMpjZ4XN9cFYFIw1MUy0Rs1I4613UZ7JoRNN+8IaUdtXrulSxo
Ea5Ul3iFiWFzjRTrLHlDHLwp9D5gvTPFmU8BKvPVs+ZU4yq9dvid+uvJbZ1ZvaRx
yzf8DJbMttWjk+12rK5RZuZkIz3wNlOmpjd1Lco2obYWbOUrTumqJzgpI36McnX4
6V4dYMuaCP5AMXP9HCbkuqsHY1BMs5qfyewglsPBs5uYBUpI0tpZGzv3/kKNSf1u
foHBQMlAH8a4DzUebZr5BUkzVGoWgbA9Gq2wyKQSN2taNFVXFb2pOzw0jPgGwENT
jg/ML61gqHZnK3IDTI2TUYEF6qxNSA0ZuhsUbK5kSG0l+f1vmpRqcLI7mEGmJHYS
s0mRezIpQbERCcrIwXyB6ZMlXIc4eEaYz1zgOTAAsbODYJZ6BBfVNnabz9ocVga8
0xEAYbonPHMJelnasioBwzR+HqKwYweT34F14vxYHIu7Y2dvyZ+RRFRYSU/1GpYW
AbZa4CYeQpNnQ1X70Ddx0f4u9Ad66Tn8Y41/LbjPcartDJ2K8gWssfgoi5P1rj7H
cBILM19yJvs5zMUFomUrmScTJXC0lajeokpvXN6vzNm6ZXcjG5R+kHv+TPJMiSlK
ndFzPV51fs0LfsQGvmKyw7Q4rxdlAN96z/t5JVaRNlDyCN7NUtNo7nYFu8gdpIjj
ffQBAaL2Xv16YjNce033jfKFAT87vBFgjGCqT7pX5LBl3uSReOs3WPEqHzFSddmA
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HtI5vefd2YmzwvVAKxkYieak0AGeSg9nB/3vbBwxwsYBiRdSeKjdJCAlseXJ3Na5
wrfOe5TrrtkLc6S7N5fqClTye4MNoeC7mKcvvxr+3/1NTLYQAwLwVm8Rl3hYEl51
BcP9gE2IqiNWO4sV+jYreAmIlRRf8sggfi7Gn8r8CpAVTpGLG+0KVEX28rb4CbjF
OtHJavw+TLs4gIB6noz+teAGK9i9HO2ZKq5p3UxuqBcb0mhc99ERavWgQiJzJO5o
DSzQi+fuCgj0GjVnucYq9oE2xoLTCBFDy4gvoBRbL3EEokS2UDJjWCQorjGmhKFL
ckBBzW8AMrmOaV7vPw8CHQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4528 )
`pragma protect data_block
jbNb20z4dMft5NCV2fPngTN13pEB35SOi2nbS3tGHDwvn+233fbCwtXtF7q7zep6
DeotGdPz5ICoilIkobd2pX1eujmVkdOaAQwJ+aBZ0FeHn8BGciOqH+Oqct7UGzyE
SUYDzRzAFaO41yJCibl4YQOj9Hw0FhKW3rTy/7rmkPQSGeGW9buILhNLKdEW2Z9J
AGShuxNlP1rvT+sJhXxMckb8Pc8fyZNu/gfbQ9ze3w6uJUInzuVAFFSvz2wkNpXa
SPLOyaQuECQ7RF1Pyn/n5eL/kVVkP5JhfXlkcb50j7mtxRUrQgdZEBl+alQWund6
sEb6A8pXUV9aqT1QnUJdMXYEbwpe3M7TArDDbFjH0uX7Mmgnv8Ou++UdbapOioYs
zvaHpz3rBh8+Z2jB0Q0TU+pOBtu/33u8pe+vl4uj/SAHm34SiwdPu3M8w1LFDqYk
OOFKDdbpD2IMzGIRYcHV7nch0xKWQwBjmHbdo1yqzOxqpl6z4nl/3KdFg9bdOlAd
g539hNWFLNUciw3NauisuWh5Q68FtuN4UIDdsX/6oWQJgraaJYXQsfRDnMM7yytT
7gZucTlCU9KcDAT9O+W9ATTyPtLuXdiwIz2Z3yMhOGpDUbQANgcjKiTXQTlgIY+k
/Je694aVF9zF9prj/wx5DmIBvalEF3UUEkivnt/ffdXECqTDpal6y26u4MwN+g8u
d12KXsilJRoEgI1sNWqNJyl5R0xQgEUJy7B8qoS4F1e2Z4BUHBf7ofbr/9fYIKjq
AtZQh1W6E0zAHdISV7P8xxYAtqZ60orHLMxZMow1boWmSiy7IZwvuVrCopL8+mBm
mGEQYaZBXjikSFgLh7XSivd+dS9i8HSdtK0bCgwOLgT8SC/xbvQBO68zUfwruevz
Eq9KXuVHxbNwlQR5mGjpMxQUlUdT6g/FqhEGTy5drNeY7q8bREht86Yt4rJ7V/UH
Fleezv3cXz29mPAnbbNi4JWIFTmUlwbLjrVCkq+EMdjNTQM4IbYZ+DbzCRN6zyok
QJ4ofxo3g4x9rmVMupTxO6Wzq0S2pKNC/y46PxKzfWPTWGbvPXlQT5dbPDMxxuay
J8DEEAQODZJRTPC3A3D9MVZY0R+mpK97np1K0DakdUDQW/cSgtDl+Yz93DA581Es
wq2JVZ3gVFeLlFLK8mZ+Ps+46kiaFEUgVvJfpp1cYiMts9OQddM1ZoxxXQCPZ+SM
ehfE0lNXKL2u7pjwPb9g6szZRkMqkXQ8qEZK8MGAyN5arDGJGSVCOrB9BZc3eIZz
UYL+NCLvuz0QT8sd0KCDIa2jLhZAKRsX4KeJ9XXgmG8RRR/g7yYflL9NrvQSVzT6
WOY7Wtp97fHtiAJDR5hNYAfW0+eSLKWb1UlMKkf1TIIdcqJsvLgRWjiIKv3+MfLY
uSdxk1d8lZNwu+zu9/qoOXBhAs+uqHc+2fTYxHmZsmYcNuveJeYd6dKYBghrm6mS
dPTYaJ7LCPLtUgWVUKDnMvQYkz1YdYknDWaSpwdpbmhZ/8eDsFN2SlcD8LntWLuZ
+T8ZHrWPhBhl1nA68zs7pQtUR3RUwq5By90sANAsQUJn6ClR7vr5jFk7eumvBPRo
EAwk5t3iMCjnQYK1ts2HdVDyVwWkQT73L0Q2CJPOouOx7n6CdEuIP49tkDTO/o6C
iYg+PgLbL/xjCtiB+oKtAbMRewZik2hCbqeoYkzczPHx+Q9PmgY8snmNRj8OL7On
r48ZBo4gKJbvOyI44Cvnd/su8odWZTbjJkcvNG9CkWedCHcOqMVxP2jKp8Xp83f8
/QmRgEVOr789kxV56TRdd/1rd0xBxUE0gaR82i/78IcizVzF04FZhx9ZBDCcxEiL
orBKWAfOrSADOwNJdOEiQ0rIhnHhlPxkhuSPqZmfhFrIxWugwStnNjPyJqVPzE+g
9sy4lu7xoKm8n6M9jtskzOrxu40Wdet9IqQgIhLqAqwIVwkJjbSvY62UgCZPUB59
NYEwNPtyM1SiTrhrSG1O22hMfEPIORMii598ymuN8H6cYt+rSMsaG+wygU6ET4BV
aBV3K2Mf0xereNaXCYz5fz1q7++7NeYtYaVHw4Wt+lii3J8N2UYsqGAVvxlgUHXP
QN8a2T8wwrjWqYR2czNV3YifCn8qFNgrKvIzmvwKTvPsTDIvricGGgFReokumg6V
+f0jXyW0e1Qnafho1xBRLpqZVzR7Qz5O8aRegy4m2+sE7kIhpsV310060AMRMdIk
rr8HiI+l2niODmhhS9rW7GsvxQxOZPqLecP7YCCTHVmq4BHTVUFX+G3m4EKjjXo0
jRgiFvmQDpbYPkAJUYwdRr4tRVz2+PXzM9QvWdkMzPn5f5QbYocUNqsTgEFTnBx+
rQ3W/baFDHMze+PX/OsKpATrmMNWbjVvedmNOw+gJ8y5WHQYtKzu78mWjXV4P/jh
xL6KNHZfk77HJDvl2vJebdMUuOJWchL8f5Db02qEB9DjQoYld2T5qYZutRSbkaVl
QCUu2vWj9xCAOvatKJS8nFtpQC61LwY/AGigGVbNotya6woxviNFT8VQ4e7KNXEC
JtmMlYzwidoatAe6cRm6iOCPnx1O7N5zJzvAnbuHGwgAzw/9/8v291YN1Brzqej4
cqcOoiy6nwlyA+tabr9PX8gjf1NERI8c0rq4t3Z8JbJTQ2bw83Y7qy711Fppg6Sc
TZbJsPleFkw0uqsq8Du56agsWtNR2t95Bi4FRm3rNL7sEeBZbpRfUTbSiVXHWuPj
SraqPXvyE1FgcTyDgmGaQNcNtEUXYhGMCSaPHn6BjpKLHV9SP8/wy/HGuKoygFsi
B6AshMercv7k3h8cbu9AD++iQ4UOP63Pqf9hvI2/t7BgW1KIjr4CNiF0ENEwZn2N
pNs54rTLulpeqF6TDFJPWsrJZYfYTz4qQKRW45Sa1iwtnIDQHMvpuKr8O9tEe66M
zdPQYtJqJqv+IYDhnTn/IO585rX9GRsLL203PJKS5oCCK20jyuYMuRZTroB8zt5q
vannQlB9e4acc0LO2KUE7t9g6jCrJuMs2Rl5/0UMOpDFsWEZ+DUvql/v5M9A7Xmc
iNyejmDXMyYR83ZA+GninMQajsF/lpd/GMh2Jmg999H2dikqq4zwP+sLCuD/1tDB
5TIL/kH8CStRXxOO9yprxKBiRv/lqeJX7ofmtyGuWkClNy4MnSDnKVgg8t9/3gvT
NQaLz5Kz9AqKYRftVyVJPL1RWLVJcQeCXm3iUBmo3q25p8ZaU51yE5R4eteAjdK1
c570pMtDZyHa6PQt0rG2tGy98fI83I9p+qzrk7lm/tm93ZhAJ7Pl+KqrXiXhT6zU
6mfOXsKPrSY1c9o90gtn7+BYvKgZxNN5o0x7itHsd71gwVIrHlLNpeJwkIAzXVMC
3H3P/RpioigZgiT19ROZKEY8RJhs2TSfi7O1HHWAB/P8lVvkwt1KGLzDAA5fkg03
zEXa//IQ82s4cv2OoUIWS2mRw+wArAK9/4EvbgvhGaqFwRtwr4C5EhYxmuFytgjD
ueGhJThbTij5lySpR9gjXbhsY9m7PktFgpGuDjZ1hpcqMBB8pUwXQf6vhHA7cizj
hy2LOuvrslCEW0eSsAQ3tS8Y9bQyZKAJk1689saAFZ/5W71fLjMR5VF+iobG02El
AD//MXo4GRKhlx/6gyMuy98PtnhQDCWhxj8G5edRyyPf8fzgDApUN0ANlW8SgaW6
d6UJGxcRT7tvBfGv0l/MC47PjfOwyX+nJpz2GuuF+K+fwaYwg+6FdT/hZApoxFHd
ymfaV/7sNUQI6t52WyuoqJYeTn39pdBR7nGEJEVXMhIVC4mBu5/k5yvzFiU3eLky
6ATxn5gt5hqXA0UxDZ0c/moKlfAxkis4cc1/gA9G660+E81006HUtp3oipa6LEfm
ifq0bi7ZwWXhq5qEWKHlSxEc5JPeXvME/kp05Zh2+dfs2KacmecHP9aKgogV0NcJ
QLdYYeQAs5PfE1LYWxPGSVdmHsiP4zxeUjuF5IRc1vmfhHrXveug/OZwM6hoiYBn
bTaChZ7NtcEnz65t+OYNMlP/fgUQiziqnqwpLIjApMnFKBrhriqv/4VWFmVghJHM
5sapLJlGxrbJQmqCXZJ6fMjdV3GH7+QoyE41sLqmrxuNiOJ/Bmf+BUAEAdQiv9SL
8rKUESQdjJ2hJFyJAqIP7AalGcU1IUMv1ZMyRRTqAKBBkN0dpIaevsEShuVb+pZS
bPo0QUU31USeIYaqWIAA2aAANAO90O0yOLoxZmOICKrznKs+aqeAPC1W/46uvaUO
hoVsvQWEHNcIoZQYS9ZzxicijX8GpOFHCVnDIoZJFdfR3wa9QeF2XRug50uP+yOP
+sTzQuq4OR9CqSsrhC+nyr/ev66XJCZdiwUBfIPjuwk0M6Kfu6QB/dbco0pKKjJw
1HJRYrUnNBoy/G95IneyqL8U8coaiWq6o76V5ED1ImE8g2jPIFDNSsO6ocRbSEPP
BNEC3Y8ePpmecpf9XXq1SV/wvfkmpXODJf0Sxred2n207AKjy35hkuyMXOTY73qV
ta/H+9sOHIcid9xEJ46Ik8V0QWDKAxGS2MGpXZNAwjY+5aXGtVTT9hv8AR/FDTHB
q8GHo4MSjwHSnlnWLbxFI9dotDuU27o1/SkqmD88/Z8DA1PCr0YcFgWhzJ696Qcc
rpQE23rLcOlXKwyQaX7cQr2dh3aNCuveXv7CxNn6GOOXOijG6z06nY/yaDp0jwzB
bVAin4L7nAIXJLkFOHwoeNRGbt6esTtzehD+iy+Cwf1bZeJ98IaV0IkiT0mJbt3R
ulI+DofgyVwGXL4WUW/gaVn0wem2uS85SqDSutK4T8rl5YBcIkoUAPA5AWUM/Yh3
HJ/znAVi4zUwJnyq1qATuULJiEvStGreHPWXHp/2ie7QnIIAjo7xEa/zqtHOWnHb
uo5wHJGAX1ybSGBXNvQc4awwlyNRcga2jVClcUDsNz4dEorg0xMZ/BFzTO0n22b3
L0sTXgtlJmtqULptHNrZLd4PyghoGtYmJMSO0Z3jtycMM+PpylpAK/fhnKOwfs25
28QL0/P8W9c3/UZebNmk4uwQJFxouYICk18Ks2PkMVA3pdHHyc4ThYadVpXItUd6
dKsKNHBdBFQPEABjJ7mT5xc5D5sADrmZu3b2gXHWDrXNsu5g6KebtcFzXm5hMBip
CNEahqumSXGjHrPqnu4L3FoWdJlPLD3xw6xyhSASURMpO6xOi0cXOvmX2tUk2RDv
6EbWqPNiz0asZ+WWWcuwOGL4REUvHdVDi6vE4ArWWiHI94CHb9q1wsHChuWYjd4U
pDq36VmNjd9UkyUj1KBrMpGmR4omckPHTYTmUuDSFrgT2wPob6XnAMhNBSlEFP3r
BSzi2nawLycPa0DwO65sugM71OamAW7Q6PRaYdITrzHjMZUOdizrPfDy8eXp9HRn
++bro6hqlLMm1lyEkUV34/J3Peazb4XzoFWl2VqSq0Q9mRKMPQSSZZ/z9IPFPemz
crPq6ySyGasnpnJdAAmZ0nx6KSrNGk9X2yqzOi9+DGQHrqbjiMalDbj1CSPleO1f
1K2WmgOGf7mkreVf4AhLec2SGY2q4zw4MywiSS45t/9WKapoQWETSqtz34JQC6x/
gV2Vhsa0pFUANbJNxLvl3fy0nMSSDg2+jt3dCxtgLcoQ1tzdof+DbyGGxX3oZfJK
tEPWKcDdNVN1cOIRQZeWFoNfcF2wKus3vTfL6rwK1P7tNVm7W8T7oBKPXw5XUtnC
ajlPYZ8q+aUWXFkti8LanlTCxvepBhYMGSM4zU77lvYMnC9s6SSjKCeNXpH6HRZ5
c/TeSG8WmMIF73srcUgZPlrDmx8aVY2Y3VkVN/liDyHp+VV/CNeLHh7DFoxstRsk
HZ388n5O5f+XdmL9n/M4HLNeNV8FPZFChC9dmh31CzaF8qBTuyPMdZWq4rrcSinG
XMQzIyxqb4BtUvRikRJ/gBQeneqN1pUz4jnj28kda85k8EkDoJZoxhvBtTd/GVbD
1IZtwiDg74Q+Sddd3ZVHZQ==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
n4X7MjCoEBEJq3Mgyr+JUMQAilHXtqdKo0u7lMU4vIDPrsJrPI4rE4MyD/BdvVgl
OCtP8FYf1SYX3M92/CmmDWqKnbFo4RNQHD9uH2j3CqcBgrjpSjuA+ivID6nF2ReH
X2sV7xZOxHusK2+OlTTsRyWKfGTUHeK/TFWJONojQRN4IYpWcq7ULfuySCFkb/BX
77S051nRvQ3d8KbKwllZKLz8ODq0P4UuTxC3DMGCY8tkl6YEPdXrf8nhOb6AZM4G
edxwcBSgN8kHWPSu4T4ijTsu+CZkpM8OsfbdMm6nUlga8rqXSCsdLDzpiK3nNBKJ
J8fHIUcrH8ELVwGxXWTivQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9584 )
`pragma protect data_block
HyhCt4MdEJe002K0Sj2RHWGlaPV6JLI90in8Kp7Wl6tALIDHsN3Ln4oQ8dZqIOYT
gJ9dRhkHUA7APEtfyX/t0ZaRZ6zbTTcAVW3wGZURT2tA7uPWIpsONz7RVqF5tkMo
JHrANBOsquaZKLJqjX5jlLm/IiDbOYB/ksmLuQnmGZruaBCdgJDVoPuFe3Ytc20i
8Dn/PwYByxC0SFnTWiADpyEPFds6amhtHkH33f8sxtkDThC17oL/EBX98Y6jxzDK
qxWWHxAlU+Lo6zIHQ66tVCLZjeKiyzZwZQ0FbnwNNg2rTPmiIyUF19z0dVh5yDwq
Tp5PX4LeMpy5jw87PW3ep6AiuRETdyZgkQr+vZ/cXe7GjjQfEyCvObrWoGPyUY7/
Dg5iMcMiqpA6+rvBbBsE5LJgJ8cAjffAqlzZ/UcgQk2lWFJGme7Q0ZvDyaYWgUrv
7MSgHDbJxeoLrdlKuVM1N7YAcah0H4PkI4eCfgNMgVfHmnLvH1bgHkUzX/h82cTs
6lGnnOQRndJozd9UZ9E/A4FYmObaheheGapWl30d2myj0ckSC1aQRnQN1b+p4YLG
tNWUSEKSxsr7yJ6YXGO7+N6Ot4KdEhciweYM80P+ePMVhQrL6QOYNMrWSuat8Rv8
o/YEhbqIAG/mKB8CGqmgQcjXFSa6KWbe/4j1h5ygxHiBCVMWAO9vPnbp5u25PpN2
Wqq8AFvSOONBJxrIuVeOVfPI3qelmds8GVXTw5WmyZjZN+FIiCK1N9kVfr5D/BxW
PqyVFJuAqKgv9sHbInsHA6pWY5uUbB48IcnHNePse3nS3DFBMpPjxq1me2oS0I+C
SCOFf5w2jbmMbPjm+f3bAPpZJsUliZVUdWZJPBcG5AoVL8R4sw1QLm51MTQb/Iuf
eAZeitGymHJQSxfjXiXrQ3/onyM3RFQihZfqxvoa2YU4l2Sc4L/9sizDNCm7Gj+9
OE9xu8/1mj+NBP74s4vAkAdzILjebzB1zIVOq+Ua8/W7A0xea23tCvIowXaG9WGM
pMd28TOSA5ty1g2D3dK3tbHNokuAxa73d/r5ZGLn8aGGFfCBp3cdAQFhXJ6RaEme
4++z81ZYJIqIVZl3VM57D/rS7b7xiWjY332jGNs+syqy0Jgmw2wOtdgtWDNjVbrl
SOWpLSnhaElYzzPPwbkJ54l/h1RWJzyJRGRSUmNVAF2cOD4/29xR/j0SovLQkzSr
2Za8lVPGsBCl6Qob81KcbJSoJjUPErzyRFhDP7UhllNfjoVq5sksmdC0ccGAjB9h
XsvibRX0H0UuZ+0eXKYwbm/CaCEHm1EgF5Po2KkR8e7DMn+TP1R1jDuBRsJTv+1X
0cUN0b5dHq9+QZj3DLZoh2AZWx5uNIJSCCFE/hJf1bCQdT58H922gteP79KiYiER
qV9a39VXCpAW0gFYCUhmhd9XO79jY8M2h44omSKURSMTxUljCVXYnaYZl4bIdmZ1
2fLXiUgHBp5NKtpubbSqJkyptl4cyPJ8vQnnxndg2Awvp+w3/10uQOLlT1jHM/zu
iGOwXwYOVhNHB/dni+QseXZWAlPEEaeZO71LBMj2E+aM9M8qQw3+n6RmbeNHwrFO
NN9mO5WyoqbAyJEA2ThD8RCdBWqgU3RZr/gq/u7XgEEA7dB9LBXOuF8/v+l8qNQ6
gl1FFF4liOSJuJyytMoQo2DxqLMYp/488o6nsX15CW04IlDbeMsQKxeqbXJjDa6v
tcIzC5Ipyd71gWZ4X/zHTnRcUzG2yxlKsBPZm9Bja3EXdj6AmDLzqnwhUSPEJkTb
q2PpOtHxIhr4vy++igsUJ425aQmSMXxWQ55F4EGTY2pR4dd4p5ZHVT8XiFcgu9DS
ZQxnKJiFJzXt6Qq2aCIpCr4zZWhxHM95v+K2mumxINZssXSOlEY+V3akh8LA4/yh
auscc5O7jnZpuuwOKNS5wCLeU/72fFChIWFrmDZ1QIllNeuCu9Z6wJTd8GAdStUQ
GtJFxD+VQZ5vlUTjurV0Y2uwMKdm4mThqRexSOo7Lmeep/0TEdyP9evIMCv9FWn0
ovKTOjimkBg4pZlZg1zMNLjqIYvqCKKoem+357B/7qpC+qS9NsjvU3BCEbWANpmY
YRFJpuMbiRYYhJGtk2nZVLA/3GztYDmkUSCstpL9G8ReCXMN3iFbSe4yI8l+rpl9
FCAHYvh3pJHfSRwCwn5IerqGIgPjPg4o0rnb57w2a4NKelojxPwyBjL+MwJhFcR+
KlcRdiC2ayyl3ElWOOrTm6XQUSnUr9fxTlEWj/NzDjFL5F1jC95Ox8HLdmq7HaRf
ltPEwii5CY0Np0JkMMujOS993GE9bVQMvUTjrHqz+X4XV3uacfeItGLFZD5oDpio
vntG+JjCnCXfpzWu2sJGXxr5EwQYRPFUeUv8mRf5uke6d1ROZ5gFcNVwWX4ihNOT
JyymZ26/jjbHSA8x0oawRyODjtnaLyU2meueUgCHN42RyqJhMwMNzpvWUp9Ith5R
sjPheSkFDpwBMX8qm/0Eelf8Dyh8BxlMelw8bDXL7NzzZJIA4INiI77Owpb73UZ8
2YgITCGTlMQQBMfJkZyFcWCwIYDM1vbCbMRUpIPaeJagw4QfdH8KCQYqD6YATxea
LJOXe3ds1L79vL6nF6lm13w1vOacFBAkWQlyZgQ4Nt5d75Ta8xurvHaVQktgmQCy
S/L3UvyiDToWsMXzEcVNK17XsdcEJggnDEbuYJ5xB6kYjXsgVDJRMIMh8iqu5+eV
AQ33Bnh6xbBdKri73mYuTasuZUw7shBeVLQ0lCapgZ4FFDVTrpstkEvAuPsPaMK4
Rbw8BuE1lGN+QW1EMkPEdyJaXmSND0Fyea5uQHz06KmjqSTFBzZzzLPEmaiw5QrC
0qWOtuXsU6Pmy407acXJpmIrDVuZjTsROsjwcItt02qnmX78iSRzMg3G2R333Bo6
upcwIQftrXafb3n84MtPR+kiGLjDQc4zgWmT1b/DjfLnPYA9hKoHxYB9FVmzQDmg
2XoYar5u9GIbIqAzmPAT9x0ynBsb3wY0osQf6a0EkRD3x5Zu/fn09AE6L/jfcprB
skTgOhwtEoXWTw2j92gqqA4Jb0w6stwKWKNqRHdI/SZ3fvzFa7yvepuOHAAbcFYj
FqttOYfjG7cWmRKRezXYVT9XqSsM+SgOPBl6Y9Po//TfDhbBKqDOzH0thg3V5ouq
w2DFt7oOU4iUJ5kXIx0itOIBfzO0Zz9v9h5G1/sUCHvWmwev3t693nESECvbCTOh
avjNgUDPQMXeVSlCtl+SvovCQUKy6vvG4C+gEwaBpWuJqq9gT9ACWRW3kZ4C1qkW
+zUDIJqVFayQcc7spO2cnAoQFyin1wCoKmFgotqGkiDGrMZsIKXdbOSn8KrTJhGs
8Bl+yJp6yRnX2jTeQ+HTVxhQUBkgLX87waXy/XIBLOqnqAtQKoaj6fI5Kkknm+O2
YNd1BdirtrvArq6BYG0t6dvwxhlO85oiIqVSt5rgdRieB37zUD6DQGzck2YwiksN
Ig8DjidAMqMxRDKniExzUfVTr3nE70qOfgDHRTY9TxXG8lJ3bTl//6ugPa5MEwgZ
PCvbKkQJdQRKRX7Vx/bozEQmZGzS3X+cL3xLJZ3UrnulHzdS22EQx6Fm8jCOZpb5
NPXXeXjOSM3NYUUHSkZMJg9NzdD4hJTGiWmWa5hawa4iRBAeg3LiMo23/11XXCq3
8mrEIzwC0rqTFHiL3Ka7LpsNjiAquU2yj3t6cYlLJXSb9X0x+2vmt90LMA0p9Wvl
o98toWgBS6HVvclYlX/Hv/BKTvKbvvrgUs8NNDp4yQYGWZROdtW4r2KbWaQio6Qx
o1Wz8a+Fcnr7/hfoPBZCa8stQmVXvWFOK14VVHJQAkU7QOz6T2VUM6lpDD61YnWo
u5N8lclYSGQoy9vmIBEHeugnhHUeyxblxBXOyjSbro7q4iQQVQ6d6nFoBpgvxjbG
8iMcAXrpPpTAbYDE8ckvwFJAjCgF0lhK7Gky0+l72ZEqxKp5b6G/2Pc72v0j0AYw
JgiPhkIcJJ+XJboPCL8WhWucVq7y8VKCXFrRZm19hAnwPGY+HaC69xEkrR1yxfeV
hFTjebDllXRyhU3vvZEIj5r+bk+eByJvrdWtiRRXaVCHY658P/COCuZU/KxshIHg
Okm/AuTjk891G+upr/S/IOxGXLxgGAVAil9B+v0aZdSSE7GaO/xxSjRRMzukw9dJ
/rcpeY7ZlOuYksn5zYp9283GUTgizxWxl2EsDWcC/uSh1BtK/dyJKUg7WD5ocI8d
cx3ozPVEJ4HGXXMKiGJy2FSkBeBtyTYmfmZ7mdp9jJBY1DWukL4RrOGCT0ydY4mn
qsRSVGsq2DAkNjamHQBXvaQsBxqfXVFR+/bKgkwdofGhaxRrxidf2G/wj86ODChg
pa4QI8IM5ny/GdsghfB5jB+R8RDFcDE3MVrP6BHNOb2i1CE6Rw1hd8AdmXjtjl/T
PBYndFKN8V3Ejmx/mzH1LEhNHonpmC2yOhwy3xipdUeBcGilQOAiGJIWQ21ylEKL
yQOYG61g2pmHLBFVp59FOlbn3ewdjBQMoWNX0ZyXHdGDVua3/IP8zm78Is31PbYu
Zlh1mVgj4rcjvEX2/PLam601LDt2gXbOC1iSCrSfb1M7iS3RnsRy9aMFrQ8tZFtP
Cu7XnZeX6lhL3EI5xF6yIZUXx0LcwBcD5wbh7sjJhNZBQ0ar+kjgteyr8HxI0kg7
sRQ2JbpBcfLaCXc5hJArXT+FmJr/xuShstx/n0mA70Yn4MX3aBzmit4uzXBuU9Gl
IEAoeRlkpYE7WUDDp6DeeMQYPVMYIOlVfHSpiTZYQ4iqqEQeuTWjZ3rPWkWqrA2F
VH6hteDFDBfRaG0cuQFwxXrrmwHPssy/5/blSiYrwNQBoZmEKpCjZNMejkEhyVDR
LDkWWFDBzGabN1g+b7si9JJ7SNJhkWstUo+W3htScRFU8BXidv5Zp3e9l/zB0QEk
WKdGr7BjTQe8TmjuT6xG2t2Wd/wQ0QqoXWtya5zu0WCrWJh30MOrDslshr8a75fk
+LL/Rf8TWbtI6B0mCUez2OE0Chq4iF7gi6vBgcROjtCGztKBwp8r6R4VxK/iKZkh
F3mHRJ/i1T7sg3+rgAyxJcemtvd10Yd4lwmFUo1cQCmIR6MKGAtwQHlFq94wBXYx
Xm6vsw/2MhU5TRRETM1cBGnHm/xIiaBKjEL0yu3hO8OSa4jBx9LEOJ1vOaeOiXl4
62QVgEjPkEhEKRDE6ft6IgM5Tx2uDFLFBMTaokvj6Lv2KcN5mSzrn0YpcVM5crhd
U0mM0wfl04egIRKzFOELa3sI4s/wL4t+qf4YMHqnFhLRHyT4mizWRna4IaCCZ0zI
roK64G7+A3S+NDVncbTMfzF5uGpJbs8KI/oqGMVo1ZhOhNzl7PYG2jgMuAXrP0KS
LDgAH95JfbLV67PgojWFNtGLue6H9x1yvLSoBOyw/Oame2mWysDFohfxasYAbdBr
9xWSHQBT1BYJAvU7O9ghTB4yXm5AeZAN/mpBfzTJW64eoZfvokjLLY0M8ZyzPNUj
Ep4Razc4WZzRoS1pcFosKIPMNhz5QWy73v8VoLYPKvV7PW1mNC12eUnaDLqcjsSF
v2j6y04gdfaUl2s+W8ry75loW9SGRnDMaprk/8CPVLIKwFDmSi5VZZpH3DSCIsVo
dQZm936WrwSX89fbZikzLytEtBo/KBpAaLRctPD53Zq+QWWQVA8esjkhm1tTo3mi
DT+e4Xb7sGYy39KS3Mo6NIDC5Yz/Kb7VsxRAtQNQz1w1By65iwlfM6blLfrqeZg1
Zk7gfBXJE+Do2CCHdVQy67w4kAXmb7I9DvwpVflLGIUUFCJ8nRNkJBJrPg9cVz9U
6+Dszido62v84hPni01V7SMx1GKRyz2yJWGgMR/v0Y1gJxCFQWNANezgDxoa+yOt
oWTc40JdK13Nf4Q9s7ekXSLMDUREwFzuttKfPQQOBIgyLOkKoWCXCKbDXeculL35
EHl415plWUVkJUA7QWgVluvpl68GKGh3rdNOlv3/Qx5jfFP6LAKnOHQG2vPf1ivT
WdZoE6dSVshGzxP1wsSkeXNRDm5CzWMY42Sfd1FAiVjYMc84SfFdZr3Hxst4EhLT
7jpSJLxPHI4iA5GwuAT/VencenzoX1kZD4k4fVA7oQjfwV/0Ye8y6L9xUc2n5HDW
9Td9V4cHCXOTBdK/H8Z+rprQUnDhenSVvALllG9MdexYRTFfBeDxD400u+cgMI8c
cbSB5BZq8V6WoqB/Ke5pX0EIxhXAYPl4qmKUT/Um1ZzzM6yMCdvF7AVkgLBofRcG
p67/h0Vm1h28tkAgWjGqnS0T1oy/fg354VtofUHWB30SFK9mlYkSyCOP4y6+847K
5jXSM+AAcnSD6yaQemuti3r6esPLg42jEHQo1K1YFmRly0jEncXWeQFTeHbDp8S9
Vbkl08sLxMbVjYpDhcQQyVyvvPTC8e4QyLDbMUWCCf7aj26Ix4Pta/Ksp/+mZ8nI
F36joCp118I/VfQIY3e7bKoJiDEch98a+Qk/Y5iA6P8fi6sdBRdFNNGqoF04+xP3
m3xBdPQYW0b3ZPmrG8dPe6gINbZO3StVsr0Nr5fE1gszBwpCtxAR25TVbFXIXYuO
qSdWQj2gYdOElfO+Dccbgxm7oXvm2UfM/frD8SXU/EPw9pADToBMGvRKGDI3QG+A
TWO4bE2uRxg+5lBmovlm2WnK+bnaGusEjxfr1fnG0XZWXEJ8eZ3zf22vZIt+S42a
bM6SxFY4Af4doRbHH7Wzq/BrUaS/L8ax/V4TAMxZ3w/NpsB2ftpbe/fOha2ZecGi
9Y1lY9lybCRjrkqCjqxoemumUEw9LwIrf09lJywi2/FoiQLSarNSjK96BePJHcnR
sHPBczT0Mpdxs/yxm0Q2KhWk3phs/+c53P/+Yzz7TlGfrmln2jOLN+uovUNgEtug
RUk/cEpVaaIkHsRCeAn6s2BtOiM/GvAgXDwYUmcK7WMZDD+pCvDxkSZCwoCLaWtd
cVzp8QIKUT6gBNExyVmPgZOlxe8OgCowxuE3Sp+oHw3B3g9QneVCdPZxlZXGs2Jb
hq+mEVogqCp1beA5bdUmE++7OT+0FM3WlNAsTSSPPjEhDaxIfZZjQlnhu7KTXVLM
odmyG9kdHWloHI2rv4rQAfVv2ZbozJWLLQ7vcj8eL4CsbohPsb6hFzujPHmTpoR0
9toA3o7gn31IPXq/y8af7Pe9VVHwa3ct0MHp20WXqo6SIzenNEURcnQrqOc92WbW
KyO8AH39WpmQBHu/Qex7vZcF7Ip7rbj5oN3dN6JnL2sivnQgHF6qpWiU4AO/dNIB
AKBC5LKdo5adBRL2BCD9HZr6+tm6stecbrHwYohtDqt7R3ovPUkQtGL1juytxjRO
ZNQxc4CysKFE4PNJuL7D3jIiNASBNLz8h5K5M7i4w1Vuoaw33dHpOQm8iaeWFMtH
d+BMLPQ86DjCg9P9Wwo6vXCDTL/WYovPNGLH9iQvHrbbUb0u7c5CgeMNX+8S0Xht
+vTBXI3skZlB+CSFp8evPSiX21gtkKIIrOci4oXxnTshjsFDI7GxsQ7ryyA569Ly
2lQzmZl9g492JL/COfTx4tqwbWLE3gHjVdDYDUMj1OBSnINEGgNlb8C1C3WbtyyQ
vadUCKNUm2C4r0Y1a8r5XtcTHajESWwT1vQqR6LmhPD/9pE4lQrCYGhZjyQnklzn
XP3ebYlq+KSl1Hq7tExvL3ThGm26mf/5WXxbNylBWwsZdy0lyPIQtDyiBlHf0NIe
uys41SSYFEge+hwfpxaDTO6ZSyLG7YBT0LZlF831j2xoxmj62yI02zaMe9S8bDmK
WJmErzy5DyL6DjWLKQNoCtR6WDEM1O7Johj9enNbrTtWBjCIg4W93FN6Y4zKLxP/
ZHQSyFUx38aeQ5N/s343J5GFDgLlQnlIGqJ9gcaEDEU4ZpSL0Bre3jv9nCEogDFY
EMwZqmON86VaUKGDHdLmiMsorE0BCvH/IZPadyjOIq1TgbTCeIgER5MsDXAJ2VYk
13y/FV2Yw/NgkXNCRDGeGjMcHEi2JeoncSrIe9CGfic5p8XRgqa4hNFeKqp4oeZY
JfN33qBjTpldj/myeJkF4tlipvjkGrm19OgTT/EkySlcA23qRNdiXMPb7nt8Xc7+
0p5Diiw8klbWv/7jrAfetb3L5/p79hSFiuwsAmOv2O+ukYN0YpipyJnQ4VO3v9/Q
HXlo/D+XyRKdy+SKS3pONkBWQ4Bdc9JF8GO4FNB3qowKvSjLr4OZIk05TQD+V0/L
B6jlBda9IMyY3pPZXpJQh+VOxpXD9ZxMZHZreV0niVyql7odrSvXCmWpa2kKCT/O
FFdv7PhIuB3EeFZmpkSosVQebpX2XLugNbSS5tAv3rptqz/xCZ0HOcknQ15c2eIP
IVun6u5WaeIZ+xl460jE4HGxvG+GV9Ik/grPse0xmA6LBsuQJ0m+fRvAigKwUfU0
mB61QNblyYHb5ULBjY5kFgxBhs7yp7cSXfWyONmF4HKd/j848DyEbkcLpd5MBRTw
Xsa4xhXoXq35C9PV8+JE57BSSfPyoqjGn789W7t2rk/Yvh1I1qve+LN7OMv5krkC
2pFYmgCjdK+8shan2bc6lzNUrs4FtWHOAWpoGtK7/CKQcVJgGRBmqB1FD7eMqOP5
4RIq8ZLuI4YmlXxrrRGUi6DO8yvETa9NFXCFa1GEo8wwjesoCoNai9nM+3U8F78R
NRUT+x5gmkO8h++w+qxNj5iTEnaVth2xP2mVeIKZ2YN6dw8VuWh5OBBEfLLCnhSa
Ng+iryfclEb93W3/ipgWAArR9B3bcyMcy+/Zd1xnEaljuf6iJny624SH0uIRRY7N
W/fSX1i3laLEJ5gf6mNlp5Usp/2n8j3LZopER4fxIqIUsokS5ywBrXyX9u7J+9EP
jRv3C0NbcH5XncCxNFZeOIhqspEb3xzFuwXucgqM3eyzmkYXgbjMbA2BrpHaq3MP
w1GPByX3hUpdynfucWYGu4A6XowtUNhID2sLy2VXQmFlCGJaRpH57oMWi2AaN4hm
83SI8FwZQrSZpUZQmcZoyi3E5DrEazPNFYODdRPkz4eFWigP/Ntad4i9C6IBPhUd
mNr3JV5YNHO61BNm+J6WGG2rxbZ6SdZ5x8AZwGYsUhIUkLMIJBq04ToPY/BSZr5Q
ITl6DcZT4rEAWaYfjb3YPm0sORRyCAYXs5OJsChZ0Lctt11FmRwZ/tmTulAHJOjI
kqPsfCBCVxGzAVnisoqySY9jhugjFIxTHRku+AO+SUtZHiCUVh6cOCPiBH9Ov0Sn
l+PlXEvAYxC8yBCuYzqlMQW8ojHM+2oscKNOk0s1vJPuQq4rZEjjnIqzW+o5FNPq
NUEwUOflaPPTAdeJ1JOJ11XiG9cSx+jODQiNQH6gp+lLzTnuF/kLB3oAU6TQ9cUl
vJg7U+TSmiBsL9I8U5UQMwCPV5Qumtu97YX0SC1RhmoLTUUaQXmGmwwCHcKw/gNu
tgL1U9Drj0UXUN9GHQ/9hXWn9rEv3sDqAetsyWAu9bbht9iE+PdV7LayJhbdW4eq
41cLugfNNyt4pZkNRKeyCIDFewvocc57b0QOIp+O9aIoK0jHxNrmVra8gdCHU7mk
ap1LRMaUbOjDPuh2RM8dxUj1b4zPfzqQx5YOP4iqiV/N3ekonJ4T9xwiq5jzXaI2
GJLOawCmDPeW17jLQglHz1KGqfkR7rCjnS44xi5ijaebMGNRFnSry7iCMMbEtH52
mG6/zwBJoVxkolyNcPWENi0ilkdfurJDPvSVBUmEtALhPYtrcBRVXnmEQt52KfLK
xfw5am+OZewdZ7K1CecbvtqMMNZC9bPAzxSrinzB2hyfoEP3c+Yw9l7fsC9tHvtB
ESjYoks2+IEcN8UhXnBppaSYfjc7/u1M0e29k6Ro9MfQnx/olX1c/YWdXvHahl6x
L4NHwL2NI9sVetQFBoGzJNT3vAPSXSPa1eISYv7xjpiI1swe97II76bpZCIi/q8U
Dfiz6lSKtp0ttZKEbfAJYcN1IQlH0yeCZNdcwkVAMk3+sNZxbADSbF1D07QzIQpg
SfftS3MgNpUZs1FLwON3nBGfuf6FtYYeVHF5matK91IyXkDSwO5Ekbq5XTYW6pC8
C236cvqaLlZnlVE0VtfrMfWeibNwbzYWCCkWhfBwkP05G1ssndoCsccIR0+s4rto
KwTDTyBvZSU7NYi8j0j6/JEQliIEAJYxuWXi373ZvzJigiKl7cP+zhq4AdneL7dj
g46zHTLHjdMNTX8lMNY1IYjPrX6r+1Zb2rHDQEGGufXSPm0m/8kTJ2qXV4w4K+eZ
/tDdJZ0edpk6Qglq7NllfZDNgQTsvFjTLzGrmV2WZR+LsBMaggAszP7yjbZnedzl
BbeuLK882qZ3ZIl/u+Fqh1IS1Jyv0nNP7AX5yazS0dP1IsXEYEH12WDZNkQA4mOn
gkzajE1ohz+l3/zha2cUO0kWPkrMzA8citjWyw6LOcRNNeTkKV/30ff0XzQfgawr
Q/Sa57cRkpzQ3hIQlj5BZBZH3fCICrxJUwu9rcJ61ii0Lw4idTIXgocgARo4nUQV
7u2Jt+GMR4j4sQmDxrI4ypuBF3p66EqFeBsNo38CykNi2fBUjWN4+Ze3ACO0UTD9
H0puJQgX4pQSpNWl/s7aDmh2GyuChuYWpWyHDBWY0XMzvjC3agKAtclS5kEcMO3p
a9nA42DHnzMHbWMUG3cRu2T37CxCyjRR9Fo4yyfQQPpG++m8SCnvXqCEDyBJNcpP
j/8SMDS/krwfSiHQ36hFloeAGDE339ZuoStS/CLDWBnYaLeTVZ69VG5HRSnDdCRC
1J86N8UJNExIM9R+CYZenO3kgVxZ6/ZHLfUrvgeavVZLryQnD/GgqfcB+nGrNbg+
GLwa6UMSc81Hfz/SRECqOVRp7rTQct+LOSW4mHMpJcGPiYdFQ0OSCtCkuHpeKotp
5oYJVXK49Leq1pO2tQ4FyLw9kqOiQxKnLAIZk1QbiMMkr5G7qVJE2aKTzH4+Gy+Z
XKT2RPxkrdOwxJPG6rZj4ycf4upYxW8FuF87C/v0ieYRUat4GES5JnUiTJu+n0nA
Wi5M73jdrLwvz+fEWg9SEJXRi1uuFLELwrOy0st45/6c2aXqb8wdj1/Ofc37359t
3REfa2DNGqBpYa9DheI+I40uIY6v/Wbqvni4M3OEC4JvXvpugYE7LGW+Btuch7E8
ef/3NmZMtTyMJB+YgQsvX9c76SrZOA0C4TKIVfuuivE4w+PWYJh2TrATmOP04DZW
0dSHSZDHSsXfL/U23D1EiuGfBtWrY22aEIqqvOSnHITYTtWOiD+kQCsGu2LY5YQ1
hG+7VvdQRLMnmh5UqCDxXfq81COcBnKWQoMkVbZ+9lm506m/7GEuwBOPPJwNwG/G
78b4ghUTtEozV7RzQ3PnWVA7IXlZZ+lUoKfvVv+TjSCNr/zRzX+Y7fMoPaXppId8
IdbgxdmOtQToeUsU40fm13Wjc5cgWq0j/kuSCVArsq97ipNIzVE6aCEm35kS1OPG
6t51r5BETJxXmkDMCqJHfeJKoS16idkBrPqwxuUEz+61c2igsEpqGAiN7gkC8sAx
mKkXV6QlR8Uvrp5cCg0mEed3+ampsPXcRxk8aRkyjgxjjr0inK+dXtuC9ToiFTWk
zboQRDwyXyU+z1jy9PfxmG01geVVRcWz3n7kvm4P8gIU2E3yAegrzJDMh4F+hM7g
Vc1NODhqLYV/cyfzaEyuCP8xBdqtypOo18lunb+2Qxc2/jd5zcJfCxAX0z1kzN+w
J/x5DHVqr2ngPxd/6xcMyeNX90PZYWAF+T6ApCDYZNSm8SHS/mi9nkDb3av+IOeP
270VqVI2I6mgfU8CnWI5PufIlKzLTOIGAdJEyrnPrX2B9dn3vZPbKgrdwKuOMT33
1CGK5TCpJZWnd03NBHor0RGl3qaOZPWxyMwj3y8CD6To/HuNRq0hG98eHirlPmwF
lKff0NlWOdW7LT2mp6Yp/11+/f2aGvtoLBNrJ/cN+ecg54baMUp3vOnymzP6WAai
icHiUz0ov9FLFlhsSCs4kBPe3py98AmqebhBuUkesH6wZc7Rjz7mbqFhE3tZf5tC
M/Gjld5C1dJXxc7RBDYY+c+EN1EBrc/2PnJ+bqktSOHCZgBXyLnibJxPtJBJFUxu
u7b94m7wN3TJt46k1rMu1PIyr1uyFNBfdxXdXlUFWr7RnWo0a+7bWJb7JmwG2pIs
t72oAWAbN0T9pfE+UTXt9vwrOVBZGJP2JsuCZSFOSOx5+xe3hGj1482fOimWrKh5
t+7MLegvjXZ6SZ70z+iLFwRe/NXU0kyYdDl2gZXPxrpkr5QkrZmZni4mSpo+eljW
rnjt61GO7TQpos6ByqAsBMia7b63btLJiNbk+30En4je9aEdBOShCtO+gTgQ3wG0
zGKzlg4OWjIM3ZKTML7YIJlrBxa5oZMyX+yaJGfRQYe8qhqroxG6IiDSNAqivkQi
ipweRu1RsJ/4VQTKXbeEV6GiCOSX1UVNOocluWU/9SaS9vo4GhpNmPG2RcUV3dlV
sAocOlGBbquqMARch4BzosTOJnJXyR24c/PEC0Tp1Y6jrIkNmEqrRjAXTdS/LtsQ
VxLpdxbsigFR/GJ/Ol2Ve9Q08X1MhDFUwnE+q3OUUDDPSiYnaptpApj9wBzpSEd1
ypaahbGe0ALZMsvvWz5xTaLEjA0FOLi6ouR7fL9deXc=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ejlVU9cr67DuJ9kqPabnC5ORCaEX+P10tkih9FzBW8b8IUnDc94ELb/M3mOEXASG
Qe87iO2NKVig34rU8uaSUGx7ZO3MbQsnvlj1eiw44NLXCwts9e7XV8JN6e7qarSZ
HjT/5k9BJCf4K2P5xoJfUdWTR3jtpmTtaX35daOK1zZ7qCgXi8BusKesh2bEXp/A
g/SQnN9xl+O7Am4cBqP0TM3FLCvLMh8nStFByPMV6wwOsqdeTsNaoP2nRcbGee2w
x30O9Ksu+Bl4FcCKahGn2AUEwZ+JiCUScW87UVLBgEbcq9qSWG6TR5OTbDxiRsBW
G9k6Qfj68HKX/vaFoNiF1Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8096 )
`pragma protect data_block
z1bqHXKsBvJtyioHyr7oDwkSQnOQ5zMCddTWSxwIuYKkMWV8GcIg2HaZtWMGBZ/p
0qxKq6UUI0P6uj5dHl21SKmhgQbGFTwQ7+Uor/15Rx4AOmfC14GkJP2d44f67DVE
KbA7YPpB5/iXTh2aG+5s8PSMQGl+CeIf2F9FfLc8TEDMNyHgrbBdgfvgoLZiKJw1
uL7sO1o9/OD5ZLtcd+CBOhn1v51y67M84ul84Wr7T80kVXUTwhyEJ1Vr1tXtjwrk
SuFotcjALDup3QjC500P9jXokJhefIjR/ZpmhDTTT7qgqCwsF+EFPvkkl3W9L/Sd
msAB2ZUKFV67019PrZk4NeYt0kNIaTBPBf66ZjVEGdeV+O+xgSoSUFJGE363Vb0q
TFaB29DZsgcBqfY+1RaUi+LsJbEGmP+OKLkwbevGH1fjrwHaYdYPg7MW3uV3gVwW
vpmtr61xGQ706RflaWCCpSbj6e4EGuIwwQtIcu5UUn57sEcq0fvj3EZsrMmDxUqe
IUi0m3kzF0Znli5PVGPCzsdcXgF7lcQ0XItOs5lF/hOuHHTJ+U2lvjpVwxmYRAW0
VPLg590wzRumVAIe8/SqXU3EoGf+ADWnQxTt5ELBCwBMXEJVpAHWgApaq7StqVju
L3iKOR7tiojiFtMSOWYekK1Kxv82vjVNWWvEseXmTPPvoUdMbLWbSJIgQ4jGgHR2
5NTWXuRqX/IykQTzHdFOgO1tY+uUV5th0R9w4nqNncKb8PoMa/7DcYtsNG3xAgSH
ty/7jq/Dmn6hXsOQuTkFjZ1QqHDQFuOm1SJg4BjwJn2XOUSmPrbC4jjfi4tAVQVW
YC7JF2ZjReVMOh1tixEKygtv34/gRd4DQVoLJHg2G5Bg3bbotAa3Vg6adEPK5+PH
JhukaqlRzw44+EUnhqobS/vIzgLMYutSHdqRMwFXluCY/XfogfpG8ldgFJTfO44j
NXrAvg3A2rQ0mi1+AXuB7cRN3CrAyCmyOpAvJvSoFNj4M0/SfAOHQ+jYJ1ikEcAi
h177O9+V1xBOaZyt+GhmggFpZAMAElz3Wzo1rVtQJVjrgA6vZ8tnhKFji3lmaxBr
mPkCdHQaa+iiLdFh85kA+MBAUQ9TGTA8/643kO5qCXWcwTAUmJTXatDEpm7mfbH/
5UviNhbqbRT0knwCA1CQDMoshXhy5Yr5IToKwiGHvBaBcoosRpGigPeUhVN7jtxU
ETl9X1mTuLRrK2p+9SDniqapXD7NKgwWT9o0GjqmlXrhsu8w7W6aezOSWwG6z/+b
Gihn37XS4xqqgkFOYox9yXUGDmMOBDj7G1JAb1zKjeZcf9kdUsjBO+E6Wk5iWInL
mow+HiYGaSAAy3MUrEtGSxrcUHsY2fJ6rVDQ/ES7x4g9OwVOWyjvlQ0IPmOn5861
5QKwpZ/vpF0XXSZueJVQCN4hnOcCRFrjRV17tsqAtJjL/CXIt8GEcoI1Q8Sf/rIw
E5XlNJmC/a+cjVlqUWBrQnwwYF8zk1HxXl1OgbVJ9JPSz8ZgY4VFxamHwHKm57j3
Ky0+CfLLlC7YpdPOHx700PX7nNnapFCfTGBHO1yWs4EsC4tAUv6U5pd9thOqIwcM
DwkOSmmPmZgphWSnL+QO69SIAe22y5sJn5o+QLEpMPgc+xx6G27lYOFo314MhgPA
aGZbVnkGW06xpjDf0MNKbrfua2DkArh155ozZzN5kPVtLeQ0UBggqVEnYT9OS5YV
Zx49dwGFZqdpQFWq7+hGjkTYcAjTiDm5Egi46iQ9sFGctqBqSK3SY7pudVOpx5vc
ghWKPxLwc9FT/yCGsgW2+HMGtvbyyvxfAPfeIOj36k58/P9FiGPOVcOI1LtdmlHK
damIO9qPs4fJoXdl4V8vhsF5dpFVsgO8N3rHsYHU1EWye1eSU+j25WacqOBcElxy
G5SxLwJPzgi3wGH1qO5L7YJr5bAUrHjAhisL2YIUd6Vn6219SB+lAB5AD4Z+Eln2
JQKgCaks3soel1cZhvk7RZ1io4WsD54IGZYfRZ0PDp6eguZAfaA8C8EHDLmMJA+4
0QAXXDdLFZXSOYtsbUNefeDfgKx8qAj/UKbBFZLam5wCo1RSDU2UiXag/xoL83W/
fZMVn86Fn2O3nfQBMfE8/FRy5TgQklLlG1GMVn/5o1QN6t25fjGoZO/a4cGeEYEA
2tmjTBVYPj2hJQmNwwXFImkFkBLLmmJVgzp/6wfUdUO07yTYRyDvtbgXAqq2Vw0m
Ivl/7k4KoybBKfY3GYQerVMsaEOa0xDi6CyEMlfVQwRLUn9VRgZxskTJ6jOc+Yxz
m5zsAIRspRwXtp2egsyA++plvO1DFnkNJpU67piQ1TdJc20PYEeQveQVaJqZlBNG
oar8rMZpejo89Z45/2AdNwRFr8OY8FGnUgZi38yw5loV/ippPE0beNttT0EKXhKg
g9LYPX8a6gLxnfS4FgDLW9G7dnH+IQCTRWcwXnfTvy3Dd17DhvWlLUdxIWpK1zUJ
2tTiVISsUDD7VlKq2IdBwVDNCVU1Bt/3DwlDOmwbEB1XPVWTDpFB9mEPkRecrLHt
Bwl/rhqvrAY+/oWEYpD6scnYNj26MdxngaKYCh4sl41R4UbRv0CibnqiDkFrQBru
juny8uIMJ1c/773sV43/lV4nJxS7M/3wWjNxSXtrHnIo7eb9NdwMDKL41mUKmZLU
G8VHmopPYSD2gVsranDn4ve4UHIsZjrsRY2ruS3AyzpiRvt0cJsrJGDRqZiF2fDH
FR/JboW4t5GVifycYvxjib1XH7nLn9S1ENMZbpzOSU8uvIviBzAV6LG2loswbmCi
fs2w8UlQMqSC2BAwpfujcyzN6rSUFpsXwpClfnvk/rB2pEbcrGbfhO9bpkIVZ2rC
QPGGu5AZ9duOtkZBIfbispuO4VjkCW82FPRJQ/0sh0ktt/VXunBfzFJhRIOOfeCf
2KY3xNVncCMO8OJ9c0907bfuPpF4A5O29WX7dz33Y//MXna00noWd5j4Efjb5QR/
kFDVxxOBTL00ajGI1eUl6aRL5WgD1XVB8fcNLNz72mGgdYU3sfTIYtJOdXJ4wRIC
8S58skca9yrP/VBMSX///ALPOKic5Wce5AYGCZO5c8Kk/wZoa+EgyJPHjHodKbmO
wj+yk7gSUSKlSbrWBNljuhxybi25RuWwTOPHdC7hKfr2pMtzaOwVpdZ1pfWELxBx
78Yoi16bQu5jOD8aOjFU/nO8GkJUZvEFawaMeBtUVVVKYccb7MQXqgXQzXU7zBRR
V0s2vEI0bLQ7mimhYBmC1qr1VwaMqKZV79JXGQ5xhpOPWyZZy6dk2ZqIrvt9iDY4
R3UdF9g/a65rOEFa/M0PeVTKXY/a17bzR9g9O3zGs9O/u2HRijkE+hy9mkrG2/AV
YggarpR9r6iw85nOV0sRRUiqwA/O3p2SI8XDMBd+THTvXtLdQdGA98SDTpwJZA6t
uLOJR0fcTscDx0UMUoJlig2Mb6PVhR7N6LrJuPg5WRBDemVEq6DY+HKGAXHXepCt
IaKAQPjkKYItSMmXZ4HCtuiL8KdeSpqU2Opq2DHLY4DMEfy7U40uVSG8e9IdD9/J
1Vxx8KbdBsyVj6cWnBbkxrBWMtDrR9S8/iTFXmnOzuVGPEKdpJq2BZElhnC9Ay9k
w+BlqFyIxorAUHUtjKqcItDjUWmjP1Ll/1tf5V6STW261dxtcJywRtDbmsDOtngc
3GHtNMwvtQP5Sf+EqkftXj+6Jtdv5jbGc1HqgTOQyLCDD70PlGbDqWU5n8uZXmdz
ESXQKpX6huwNjEjdP2OInRYSXSRZAB7J2kIfZLfddBx0rwtgabAs6urV7hVrcviL
Q+FWQWlSXkvwOYKATJkFu7NtKKjdPHN2jDSEYI1/zccZdc45WXaLUqFObyZTgC9+
SNSZ6knlgmRi9hVAi1hU/8RyheqZ+ZdE2a9J74QBzt9EbNzRx/WU5H3ilYYMlTxF
+qfuEiuW6uQy1a8GW9vU/Dm0Ts+8cRnK3x6Ysxvg4hK7T6uisya/h5xNfSj75hMM
WkGEc1Yvu9yr+BX7d8fq5jrrb9sG7Hp+HF6CS+7Kt9EJVDYQHurhKhYEyTeJpmlZ
uZsI4hTccMYR4Ba0H+tW9Rfe1DT52jlBTCiL8B53f1+ZPoDP+337Up5VlO7/RcTM
KKrQ+LW4y2NqM5Z+OS70rAuZWl/e3ZPNuwIzlwFrOOkCqjR++kxqn/bob2w2PcNW
frE+oU2Oi1g75r2Jh9ZaIMtnU2fzCFhZjkC2Z/g3yYLmLaknQPvZlR+k+Mzb5LVS
2Me5lL9HGKAEXLQe0KbTdsQA0enNQu+ihQEMths6IpTypCbzfWl/M08NUvxOT+4q
QzqH9aoBZBuSX/aCoV/icfczn1p80n/+aSsrgFrCU5JdL897agDgFtB58bf/Vh1u
OpvI2WBxvVZ29iMNmNa6mmBRn3ig6BLcXMBVsKwTJRbvZ8Vg4FmeUVjRTXPxIjOh
GvqTeGsYnx5gPxzL0k5yy94btddOQvSd0yo+vcPYVaifqkGPjOTKlESjJUxRoG8y
Ra9C7CAYV95j/g1gGyMAGEytU28hL60kPsG3ZkYCoOMEqCKsmu08zZXiuMJYuPh4
jWlfuEyOq/lV4ZHIMIb8Z5iC6wybSdpLgrwA1PORCgIMJcXO5D5zMZK6Q8xAqEA6
WTxgihJMZ/dxMAg9Qw59Tv6AznmNtZWLz42OILJTVwiehKe0LjruzILNWp/0P6qi
kwvU+GqVmBaXIh9f8H0nBbOvUgpMwRpQo4VlbXFcP8m3kki2rAcaCyyk+jgMUrEQ
pW9pRf8VIg1mTAWXUTh+sFN7L4DfQWYUgaNujG527GVSvXdZARocLekpCFzcGcrb
38bW//p5xmRTCGPcNdhtM4QLVF31u0A+rOmFkqXn69MHw0AkEEJb3Xc6hgCUVIwM
AdARAoU7aORg+XrWwJ+zi+qv12J3Tt2DBPXswKiNhZO3TE84GsfGArUBTrpu0sN+
sJmIkBAPId8anSpKxUpr9R7EqUNfkqeYFWqkDDRitjUwjW1arPM8UUgo7xv64fYc
2/RcrvA/Nsnt7XN6eZ5jT458gKsx3LgZqQZj3gsC+Dz8XXw2qOvO35aMbsYe8L5f
NEYp2ffEoqvoFoJMiQ/YmUjmBzO33C3aPqt2NN7xbGQD8stkFYl7YpG1P4PVuyp5
sD2pSz1doWVnvnu8IrCjcZpQmADqMOYOA0UtsGIwBjT1AP0euPNA/85MTEfjuMG7
G7Py/j9cc0pUqBOwIqjX+DPPwM+Xur8Q+4L0wPk1iUagynwKZ2GuV7xkDAV5/klN
rrJi46nXiCMYUHRZ/ykIUksX0C3pGBAy7RnVt4vQPDuEYeH3ktcQ4eSvxa8JSycb
HxdPPo4jt0u22DEZOVF7f7lzo+q9yyhMtCQNhiZ4qE36IUbrAPN+8uf8fbvbvvFG
X0GYyfVETu3ML3KTvDmkqGGR9ao/azBhmoc3AkuNNPzCXSi2pEEslCv55qmBBDyS
bNa4VDRbMsv4bDFkpiJRb1eY/rEA96nK1QnBraqUHRdaJ9ShE76K8Py5yYjFyaR/
lsx1phpO560ffIx4Je5bLyDxpr3GGRE0gxN5s2CBuFofQWbdA8dpp5lc/cBxPX2G
A6Txis2HkhSo7/7aWi1yrSBdVlrqXdSIQjLlvss9DPSZIJa+u2NyDMY8veM/EohD
0eJYHNokXuVZeMdtssOoF6QqOSpllaqDfOzEQ5q/h4RfCreY5laRuaoyurQNPP8K
VR5MgzU2MtzGoq6iil1Jy1fr1MJWTYU3/3lH03jkawJmXkm1a7KK6zuGziTgTIC7
4paSfifX4ZqIuyZLNWvrpioikfZu24UXfefwaKqD6R8+JuWlnm0ef8hbbcC1tHse
kRrmORjTvUT6XBe1MWZ6lmZddqGby7KzvO9xw3hHcq1plWE4zencu8D4O/6K8KFa
Sep3DGUXSD6zEvNSbHGhZeOajwS1B8ofCvVVDLQbfjdv7B4KyQrg/69Wym+Tmttj
slAKNbDunE9yCsi+BtgDHqReV45ZWOQXr7uaoBfn7EFWWo+vr+PEblLptEXkW3qh
LfTydpkogvz3BykzZMYayeeeljHccu3NT1uYIR+GT7DHZrQFot+hLngVRxA7PlC1
yBeBZ6ZKjj2b8lnzwSMdGFz9blQ9/KjjYiqE9l++KE0Wldp0WBNE3vMEWjAJJTri
y8RWTv4QbKCY50ZrJqJU6GHiZHBbQrQXugSFXMStOBZ9YoU/8Ek9STIw3EdUE/BT
gQIcEKDOHj5YZTUDfiAPZNpygpfIkRpmykMXrEAY8G1L8j/AASZ7J1xoOKcVTdOq
3hFP5ESDqTIqk5ga+7exV3ANLL0tbKGtOPzYJKB3AWFZOucnvpQ2g8qfglPicOUC
ejwJQk3T0oTmCnvKsk2xOi8cCZEId23g3sNrtH/qpZFnG/M8U8UC/ISic3P/UnVU
FZp99uI2/kwugXSXX19g8Aj3mlFpDxPmjpu4cz8PK5tZozGknf29SxW1RJQAyK40
CTxZP6QblkkeotJyNExJgpybgwmycwl76fRatzscZpgbad5SdCXJZsgu0FgsuxmR
xvXQ9GoRSmH6nRYF+SLFLf5bkzDjOylIy6ULFqA+ryWOT6rCRRHXcURgqwjPsXzy
/4XDaTzLrFulzXWM08hRus30jQDvq/kxlWI2aRRe2XKzhWujmr///idMVbFIHHME
ow05Slnz4oC/S73d06t5V67U3AwbTBzJ+mYv2xmtZ8noxbe02NHkUJ3HPufKU7Q4
ppVqv4X6AtYfGiJuacFBpWD8eDg8vBW3Lk+WnKrVw2iDDkiGmLLk4065Zyqyy7+G
20f3tEYuxkJzhl+8W3F4hPKHTeXKcgYup+1IuVt2XrLi5Jvo79g+OV1MHrvE9NDy
Y5Z4IPCVYcWvVhT2dCkdF195G70hlR00zNVhwH5OH3tZrz8MRtfqskUerN+UTkud
55xmRHJSgW7f/0hXViKokDjUBQtxOkvltsaMp7cqJ3r+4D0sJJy3q1ktZoXaPD6Q
A2owfXZvOLeAsR3bB9jCAY/K5RtZpvjickWQvZF6tqMZGobNZ/U7zkmPBplRTKcs
mM1YBcNXXGMnxIC+yGBIgc+8uC6NSDPAyh7pmRes9rl+bI3aRzMGJEbu7/4Nt2UX
1xAnvnBeI7+NCkzwjy/oIWK93aeZGTquVdQZCMi/Z1NFh0B9/lkZPfE4tYMqxXSw
ItTB12pWL0NyAQiLeoLsFRLvoQyhHnMnx0jY4Rviq5cIln9RaP5Xl4CWHlH6jYio
PZPX4d0XWxlaMmB6AaaXzYifowgoiBh41naWL/mRjo1kO2w+CparMAftzx2dhNh0
mfa4GoR4AtiuJugBso/GC2QHYIegx0KeTRB89w122YDvjUmeUeMLs2RqZKExvaq8
FRg/3cGA0TGyuc9TcPKT7XHzYXytlk2AOdyDkVYrg+sTLZX6QIGcH5hVWG3oRgsy
rHRcqx2474JPFXDg9TUA2lHl+DRPxuBBLyWRZGgWrZ5r2cX1yo6iDiWFFaf76OFP
KtvgyXMQe0ouXc92gl0T/2hpGL6chQyHc7ehtRgzhsoQRD9F3JZBykYKL+wxd8Fw
dcCufjrT+Pdwj6LG07q5i2vLrSm3qoNO6y3NVq3w5Z01Ak+os4ycd90UzOrwDwKG
oCrv1/gOIQVDxVrvWn3+qTUEbdI+jA06ka1bSyqmWrelzF2aHXneoFiG4P089iFl
wKREJBeWDVQcFaRxGjq8w2p+nhgTk5MKWXfhO6Tdaq+51i9WwKR15kYjvCo1bNlS
arlYovLlNXThZyoaa3Kz4LYQi0ejzFEYY6k0R5PPyyRou3WFATe9BQm892f3kxNQ
aL0AZZzaTKwFzqDwf9gyNMHL8wxSpkAqF9uXHZaYwtSW6xyz4rh/frhGsRbMiB4X
/y0kApr7WHWT8WnVp1W3NPYq9Szli2p9naF34e/tQqDVciLCVGRGXOfpp6RAxqn+
V0aIu5rRlG/iuKywvV6npMQWk+YHH8BKLyoQr8ijKZJycukFhflSlfU3THGFlnUf
Lyd388GDNp2uwGCO1HJrFQwsM6WOYFQefBcfqhX8S1i2AiNTbHvV4iegWmaRFxRI
qj6Q1e9JlGkyfTuuL/CThFak8uqeOG2jFqi75a/cBeAaIsk+C9dRIJy50C8c0PQ6
3WWVZYP+daG1vytylFxR02LF7urXacc51clXuiiRdUjY4kdopHeF2XJhER6bklxc
30XCs3phsxNWNcWdQcIC60pdvYH3iQ4mMb4q//m9l7h7LN7af4cLICAuvJo2UqDX
aXeagagWYh/c3k8uNDxr7GG3zWa33GeZk6i+znV8yiR+Qdkn1cF0FDIO52MDLmsx
HU722iS6bAFYaD6eunftHRH74w+XY+R8i22fjKvUcWSoxuoOtrnjEMJ3PQOMPRBG
HRszsFBgLkSemRqI7mcFJn/ahwTVM3AeOdD4SG40mHWL+lATUecOsvzWYrXGNfFM
o2zi3lES2i3h7Oend136cFgV3jrTSzp5r13qBgsRLkpl1Fyx370Kl9NJFA+I2Qgu
SE82Kz3piVzRkzyzzVkTA9ZoPyBqGKBHRHXxk1MBppHDlVK3Wr4X8t0kaDNQY9/K
PQ3Vx8+Y9rYZG/MOASmqnZpLzqQcF8mdIVKsty7twUL9UkNkf1mhOfcn92EF5XRG
b2p8S90CTLBw3MyY7IYIaekAMVXeHxCI5uSEWylo0iZxBfIcIj4BdOMdrQJny0dq
vnkPfzHdJxrUXkVZM3KrCNfR72pym9fV5cltl/Uepx0KRG+siohBi2gtRbN0Dv/O
GQQSmJ4lc27Mam3E1SNVfesgAvaZFzlUKtlaqDvx2bspEzGIE6rkrWDfbOFUUBS+
HrW/4ThWTfWq8Yv1fXyRAMsaAkp9gq24/rvjC6wABolvEycsFpo13SgdVTdIxq29
qXfXTpw7AZlgDV1kyJEn/boCviWZVKbOR6iZNmvb8vpfNH302bMit2NHFp13dJ8h
SB7fs5ywipdfqTKhg9204RShxfMeB50Qlb3fBekJTBE8iddXFZggu78iEHyk8YQp
1ol/o3voFfQWS2INje4sevC/C6PvRHS8J1ZbP5eStNlVWmDZd3E500qlGJ/knb+O
sxLd0GMQELvf13CL6ENqR1Do5mLLOo5o0Mq3sY/qhP+BkdXqVGyMkCgyCGObgLd7
aT4Cfx4rKV+p2r9ncYxsJwmtSeahpNYwgdmTE8GphFOf0ij2CVB5uPWYp0LlJ8FR
WA/YsQYSat9dN9qF/lUbq9E/mxCX+rVE0wYFl2NW6nshwyS9EeDLuzoMAFdIPSPL
M79xeJ1uUigYjrDsIerWvIeKkiYHcICJjrb6Qbe/TuRO6p4GaEsL09WDOCgYGtw0
acTUKTqQ5rQ5zDHFi4VvHO9ckgF3Ui3gs0jcZYwxtkLKfX1UBNbS4PbSECT/9h4A
tfNzMEzYBwRSS0WuPuZ7E0RMOXcj2pU5wO5gEwD2RrIXr1GNtLoGl8tm9NW7gCx8
4XhCDdeLfKGsOTIubGjNeFAwa6gXCo5exGwerx9dFzclNZCdKABnKX2gvbhAmofm
/PHqRa3PdSgnBP2Ue8Xim21Is7frvFOOPff47TF6j96ogf1Ndnl8a/Zy2gg+5od9
2RPFa/zkuzvGk9cJNcxOlPIQqak+q4PO1nQZGT44QzzVR9MIyuMAsh5OaI3sifxK
Cx3cTLxJiokBIAkb+IRF/9d86SFIYfbyssWmY7Vg2Ry+QL2VmZy/zMTqzE9mPtv4
6rgoyNAYdjll4aDDZOaenuyv/LAoimteQYXW440gYXTkwcpv7hAikutE6ENvqr2h
4FH6QhWvglYBFvmGSruATIYHkMXBxeaA1HWNejL0HoySq8icdeqjonMPxOOtWrFx
RVFvpM6N8GbqJQx4RQyomWGuFvkHMt7QywoCVHmYtOi3hxkzO6MIrtytI5C/cE11
Bz9BZjFeacfgmcbOiZgFott9kZujBOppWFZ75GFpbJvhRecX2c+K/1iHjgntFm/h
hBBF/SZfQE/mtlrukmnvPsy7RI8+lH/2e1y2Wb86ZV0Gms4+zYoL938iGryip4RN
m5FHac8rLTQR7+DIrinQCb2CNxteQ1jdfcnyPHS4eXo5E8o0NRaXS1eoX2+obubl
VTYld6eMwgLeG68zSp1VK+5KBr/BKDRoh38IFGJ2uztBsds+mCPExRB0WUICDw73
SIo/MfKX5GCwfFRZAjzerK/qO2JluTJZ8rFFPwdc6cybZ1fdTvrOh3+z9/KXteSM
cMG11ENda36mEo12SmMr3crhEy36xUBwMhrc/pFrnAALvuUWu2uw1pfS53NTYAX9
UcDVX4KkD/QcYAW+bk4/97uNIx07IFFsuv0kvNUmJz9Pgs5Mz00JWCPFfvLBdKqs
r451K6Vm90Pmfdgz4QGK55yPtLrk6IDaOqL7SBOTXmtTigTEHGGkjCGIz26CRTnK
FA8IlhH2KUokS5bfU7uy7LBekaWlxGfybSsRog20Wq8tYIEmJ1fowcv6BhiS8ga8
1eEEqUeXAHFTnQ0ptM4oOuHwIug05yRZUePqFuE0YwHw7TueZz5Y1YPDEbuMXB+z
4NcIn79GNhPLDKIz0UvgKbBuvJMQEKAK6NNgzgal8doZ9xaZE1TbE2BNJgziaRNj
UznFxTvHmevBYi2CdY8P/9LV79iLJzK7zAGHIgLIJ9iX8y3Tp3jZb/xd7PBqohCG
3fWLdcxLlMZiCrWMMGCXXkGLfHPrCZWdg8LgnwYfM1g=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EzfG33BnvjlJt6treW6IBIEBc3nVBNgIbxzund3cl9dtSmRRoibP0nVsKPfUhXPV
j2TakqaBt9KOospcqQXmYssnBO9W99irdT1IyGbhAQv3atTfFVWPL9iZG8g/vkQm
VSAd72cVMLmzmUJyBqQTxoUlOZoKhZNJR6hz8pGkDJ8ibWANpjPU08M69hjK4sWs
aEA/RSAWZRyjDNruH2BCt9EPLjN8nAgVn7mcrqVZi6m3QWwCsBV0UjuaIWjNhd+Z
VJ9r34iaoAz4AM9ZXpPUeLcr+mFPYGmL4aV1QYkm2Zcd6Rvk12anC4mDeK6SebZ6
kVyQjSkRzgT7bgtBsSR4CA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 20288 )
`pragma protect data_block
OocqmmQW7LRuT2sJ/zSySdDYbY1UeiH3+6QvqAe4JJ83IIhnROPO/aupzZCqoUWd
3kkjN90/kXkstfARg0cL3MbQic33s0y95yyoRmbhhwyYqgmPq0+3p+6zkBLhOIWD
pThRA6yroqt+YBz45sG43L9Gt0K8O3On+MpiKkExL+543QX0NEXtUcCl30ckcO2U
56JVO0K3I1gUjUZilxTlRUn1GMlscTumn4kMsOGLHfU/Jsj6xQj1VM40atZj9TtZ
ueHmQMgiyUohg6U7gd+sP7oxzCgxXdDbCP//wipykauFiZWXR+BIAZtqEjTLXcoZ
iTZeTa5eSuLU5nRW6Kv2Ekx2j4PU1RjsJV+GRZbrccygmxYRnrPEfkya6M5r7Vdg
iXttpQJZ19+/6wDIvAQvTtJiyNaKRbc+618NlJVbjffUTXumdeNX0rNWnPVYqEke
Nsk0w1V1xWPLMO39e5hULH9j6kglbz0CZw/5rCJ9GahVjBXzzGDuOEc9dHkqBhU4
9VzS7cYCsaCidA96V0mky+Luezsn4jKckh85DPh2dnV/3vatV+Ek0bJvkuQH+4An
qL2vGWF/lsmOSzM7/FrJhsTS9f3GnuUIAzYzc0xvN6qYfnsCSc+ucWpb+W8CD+2y
BUTVUybNKfASS6oiBn2xUzc9M6qxSPtuv24/gEj7Gtzzt3Ocgh7vfK9lLYD3+drP
5tYfkrqv+pgXbHlfZzITuDsLWqJYOp2jqNePdnuQwDo6BqLXrRCgdPSPr1Q4Ai1x
QUd+qPstqOfOJ/1O2z4S+7zgs2vYaloz6S+iOhpEcmxsH7wZwtcDMpqHDflOC4oC
k+/dB7kMgXPRhxnETApl78RhzRlSPhUmI9z10hmwPUc+rN23JwDpK5xEm5gz5pAc
xhMCWiZNjoLrfHk1vApjBerw6l8K3xKGnEBcn/L5JlGH2ClvIb7XRQq+ZxjXLWLi
pzmt01YVA74PRZUM6E5khK8My5KmlujGqw5RNuyskx5LXzsmoTkx9GOKRIg3Zz50
IirrIRslP9HZgQtx05NNorpLeEoBQ8cqw+Besj/ux3x6Nkb6wCxot71X3ltsg94l
tCGM6YcxtILBkmQ9WnazBbbcKRPXxUg/+wBxPK+fAcBZ2ZwB36eJsMCotSPQSUb0
b0ZZrh+FR2W5ZtpIKCXRIzGgaFmthciVZHSkMYYeSPROKLUi1762s3/po2WuPsOU
gPGHGk/RpPxRuB0JQCqI8N+PnqZEN4twgNr6VaUn2w3zDe+78BJZB/gBSD4OCRir
1boxbqEySe72VYMTfBhDDinoU/O+iqERLrW4r1ca1sP1fU18EzHDWMFYWdrpV8Jm
sdsNZrzXKWuM5C0YjhyiuzzHEzeVpdjZBPaFvHCKAJt1fgZAOgyEVrmeNkoHn2d/
SQE1AOPfQ4PDbvYP+UJLDwFhD3RCQtcW/SQxj2VJ9JPdiHkycQGH8bgG9wxkgO6w
Au5J2BcgDxE0GasQHOMmrqoBb8/X/j/VbX1ypFiTpaRNev34YwuKMfee31odGx6p
vJU5fZqOzHDdJoXywmD0k6Zaj3foSlZJ2YTW/UbQj2C2KhPNBg/AgktIKTB3Hcz2
SHT6ma3cItr2I0FYTSJOEixzeV0UbBmYVeSJhXVujLVsoErh3JbwE8/JzMKwaZex
Z0DJP0DXqgQLHRHKeQ+7mSJ3D1B1RL2RoBKnWsVcmkb+QxpLrC0STX8Wem0qLvIu
t4YomijAZbSYP+RuoMNVrWBs86fg9l9/r4B6ql57R1GyOwcK3SV1amJGZWTDjeTS
2sKTlexmrGATg8lEnrRMQWh4cDGuTP00x/9G2cPlaKRKJbfIEPMSOpBzHV2pMxyF
9jvNVsB5A7F8Ot6ytlyOU5vmBdlknKFSmEyOnvW3IbgQc20trlQmkoz0fiCrQE39
jHmh+LnWF8ZmD5Zlwz/oSYtAQsVPlGWijnNNaHgnPcFpMcT2l0HF1I1cgnnvcJrH
xKpSSzGbc2JMU6fQGFduKzBP3FyBWY9rzGs94WkVA0m9QmMEL0kEb801JKGxo+9a
BlMZsRCaTva/c/lqos7dhmeVzdyemhX/Pe8uNGULWwCoXIZREr5LfzaW6yFspCl6
PDuRS3h0T0Hw1DtB2zginOCSBQ9WwBz8mGYYqu2ybf9Vq+gjsgWiMwHtU0qJG5FM
SqSYSetVJFQKk8pdbcj7bplcHExbrfumtLiONUKItb/Z2gWOPfIybqS045RNZ5xS
ZDmPFzYFlItF2iFp3qMFHaLi30cgnlEbs/l4lQ8X6ZoaDYSJgGUPv2hbIktsoxnb
1koRd+qaTbHC/gftj5AJ8XX4lHxksJ483yU91JHmy+AMl/gGl1BvMJkklaiulvS8
tyctGmzOnakoq9eap6l7Zj51L8qR54OYz2tiISnbUCjG5F6kiLSKMPkXxrLlW7u4
7UY9sRekyo877O3XDxj38OjssgEJ04bKQnK6BEUAbP2yflAP0qKm4VpNcyBaqR/a
Bx0DFsqlm2sg/HnSeP+jc+O3n9KgIcPUyXWg8+hGFDrh/4E+9XonbDXoKhY2CKNg
r+VlCdkvavjGaL2OW0txbHpAT2I+CUWFXmM26FpC6tZobxUxkngR1jZ8D6gJQC+L
lFpKPuVSEWP9ruBU8kRyLuYGtI9cJmjlWHuGebCzKy6iyW+Kp0+ZFD184FVhQ5Bn
WF2Tb5JJRXeSNCEXshRSmaJZ2QZc19XYrisLIP4mxFVNSNiaYiM8rlPEvGD2Krvp
BGmnbaur3zsKqMVQ/j3HzojsspJWj9N5Aqx0g54KfYnDjQfm8LtF0uUUiLsVZF+X
SPGA+GWthPjCe72xwEl3VVL/Ch6aoimamhh7pwthR9ND3XA7wVjkaF1SByoYkCik
DSZR61Rma4GY+IFZMj7VQFPhy8aSWammowp8FReUaZD4c3C59w7/piEzl9W9uCjr
VxFfKHep3i0OWvbPBuPDDr6l0zb8WsOgiNn4bjbSn9aG2gEDQxXNfeuGgIPlIQ6Y
yiqVqLc5IV4eXfJckVdWHRyJKuL7W1uwRpZHQRk3xqVzNkyFzGo6rjzhfgibXHwI
jQ/PMpBNnj8MGenBTfylJwNnX0Mmz1LfT3BqzUhVO0a0ZN2dVXsuRCq2lkaqJoo/
fhmyVSF+n0WtMO1Fy8jpP4TOtiyIobGzpw/jhsyyMzoeGyzEJRAi4qydFzpspLyv
RjxOHz9om2FRqxkbFTsu6jvAjfJFOH/cAMPYdTLbZZMQPhnsRI9XkuWc3KIfZZQ1
dnU+d4KxzPK21FfU3TVFqtpqJS9JJK2iHhYFCd/IKQX6qABPJF033qTKzpu6rCJP
hgywHLzfyi+vWxF1ruiYFoEnCdl29HU5r6D8NhHpf3cHb8AzX75zmXR8nwm8dr9h
0NXsw85H/R2R9162YbT5SiSRBkSY9DNfd2QTo4MN3VvTFACgcpWhw78Z09Ot+/us
LQETFIEi1x4XB1V6WIpdz/3qprcx/ky1OITUwsUOrwNx8dUbn8s5hjvnHNcluSDp
5KwTvk6vRVaS9EyqT7W+wdMML8Fz1Y/Cau82HOXh6jBpFMub3YDaGxxBsiysOUcy
r4HflTobIuuOii1gaJt09gWFfW2QfXJSJLcUHvVahbdzZoFOO/7UhzBFsh6kTvGx
NBLGOJtKmx80L94i/J/RX0qHbIJHSj7/Yzr380jqC7pqNRjMpWNhgZr10WXFPZWx
xnVzwrLnA5tCcAWdeWTDU7pMVzU9S7K8qoyFgS/TPcC7h70xtxtSFE8tSVm7YTle
F7UsTFWSr8hH46pQ6eQpxIvOstKbVnlcquxIBqZCXWG/y3VKP8kqOM0N1iqvlG08
5q8Hlsy+F3nIguBGB2NhdiiGsVdTSb7BYogQuR4WMaFArK9j9EPnAH8jFv6gV0Og
U/aFpLE/WzTI32iKGBqfX9ghBlieuwUnHar1ePHnJ/SZbtjE+3FS9uN9kNuR6OHq
s+6ghTD4fOWNq9OKRHV4bM+sShZQfUTdVl3vdio0n/ArIMZ7F2pVU69FC7G6Sy1p
tFPSQKOZ5ZhMQUmNmm4xUG7CaFgxM01/OfQkeyuohoWhHelDNcf+cBVYJKoOA+Ad
QHEq5G8E2jL3BKPNzNTJN/fTcxf7JQlxpSbUliQcjuIxZwd5FUKnR0P6wYSQt/my
MLUZF9id1YhGzvx26Aqnx7OyzEHd3ZwIGAFXPwNF+eRtMdWCFS4jfsj48T9LBq+q
gNNjlSIMgxcJ1CXkRZidBXOrPmEtXJDXch3Hpt6NzJqitidah0Ty7ILeUhlvVCIj
PkZsC7PIpISz2kJCXQYUdRxHRaNSwyszXm7K5cCYShzaUP/Xpe/ChWlAhUlblBEM
4cHYiBp/3yQPyery4lUX869AuiGfBkCyD2Q3ZTpOUBZ3AfxV/0sawwPMkR8h0FmK
0ORso32L6BqCzOa83E+gyQUoH1TblaCMTWnzHkOMEtkpYvECYqTEeYKwSquePHbU
xsVuNPlBtZ9LEOFa6hsOfTaz+QoF9EeXEsI10JsrvWrNEmZydh/z4vg8qtxeE1zx
P4230zFsRBRSHwL3oewIuMTLJIyNKiFttZoonY6BbZ0DRMM7oQSLXzDYXS69vPUM
aylSKjsHsvQyPHNMJAiOgQ975gKGeBwWs1xL3i6TZHkAqnpx6ZpkmTdzbOaTjMGW
+V36xpxXklv6iI26QJvlEwgWdyvfdMxeM+wAUKgu8EKQ0yBSg153JaR4E21YbAND
Sp+g5sRB3ZGdp00qti8zTfkOIQFQSanjQB4vmi/be3u5on++VM6scODqTWrgLOrG
5gky+0H3/o2Lf10KjmUp811KzbMm3arQdMzjqenODbY176NkVvvik4/m8GNe5j20
Ljd7cY6JXnm2vXTGXhM399CgkJ3bfCmrM/yQzLNCaqodzh8q/9cDJV40S5DK5s9N
lxgMPyosPw45kWnsQhwVWuf8iSBOXQWGOnEMD7jCytiUxmX9FRZNkMQuHhCp8UQH
pd6M4BEwpTkWCCox37gfPvPbzEg7ckINcv4OsuPAab/GnzNcQ1kTqmHXm26jSSmS
GjcLTbXZdh0nsdskLB+NEaxz78KIaxGHXwtCQW1z6zC3WBzjVS8e5OgmyeClwUif
H5A+vLXqK8f2AyTM2VvWOOKXB4PZAI5x9dv4oTqGHJfERp7HXqwntZR7EBUEk/kH
N9GNK/UPgwvjgMoUWOTQVB+CcEbWkHUPtbus/Ydidxt9MBbQPJfZgzoWfrt6lOms
94gB3C8hof/lYzE9kJ+aa2nIAeubEfTmklaiZOtOGi319K9fptJgh9proxhTNqBF
aN+XuZQzOFhekU3G2ZJSy4QPhwTAOTx9VaUAe6FvWQp8NfjYYDRxJNDZDZaKnBY4
6s/jVQ2nac8VjFZHeRQlpFFKOPI1MgaQyf/HL9YoefAXK+spyE45NpRRUAgu+9/g
LXz0s/FE0VgMm0wZCPREYqpWt8Z+jTe6KrLtds4wWCwhtbC1jK63YMopv4KxcAQH
xQwKYLQWBm+ETP+U7+g4YXK0mUnJCyfF+KoWc9yxih40i+FWw+55hrkC77C80WBw
/DTtXW/vi4c3LciG1afEgRVI8qtxK7yQEpqRr71u7fpjJH2ccdY4JB93CWwyDuVD
2j7edhiwzZXvKkPpasR3YK/tNGIyd+rio2mKDquRrBA4oDnRIQR0du/EUAUgRjef
U0q6Uz9tTZQsaQ6m/4OnwTZigfAPQXSChjVdJ39JS4dRjbf6ORmadZg2IgRzao6k
LuyoEeDx81icLnN5PfIwh/BRxYrZk2/FwalrHhG3Oh8zqFd1wx/HmyqzxGW1SdWn
RapnRKkxycFsasfCNozGn5zfBIUntwbMUp1TBZ2E5qyQ3f4VL59Skc4SW8k5Ugi1
V+65qnZv0MHnGnISifUV2Suh21vAOkaMdlwQJheJ7p60z6YNAGRSDtZCaI1/y60P
uqsjHsQ4NPPfF9PLwji4BMKFnGxTiul4vg1fpYZDU6VaOyaf+96HzbyMvUYskcpl
h+4//dCpYGrP6P6nchSidhzXZhKfJ5vsH2vCsPjRvzztQj6VOFnpq/BBWaaVpBL7
jsk2vIGqkdIwnfmc35L9zkIKK9dGjrIkqFyVr2qB5Rzkj77QioetoperprfxA95D
BGl2Vm1j68kAt3ccaINAYb+B8JUtfmN5PfSVc4qC53y1UlsfkHmH+mSfsszwV3kV
ILy5CcWyB2uPLk7LfIA+03mhW/tVAL8H6TCK88APLMti7O1vKLlHXrw15qeFLmLg
1fJYkiQupb1BureRxXzvhCIbXMxy8XzP69xst/JjaIbpVz8uk57g1oU+/NwZd0Rm
WqadfiJrpAZogQm7vjN1z2z7qYuIDyzOG5UIKZOYfyUHSwhAN5N/rr/2E2s8pLPt
BSosBJlr3utEM1DwWerU3kMSZPl+EI0hqKjB3Sgw8tGv9Ih/Q8y9GkbV1BoIxD1I
r2wmdfINTJZSWDq9SHVm7Xnd7UvPuN2XPQewTNNKUZG1VI0z4MWeDjX2TSllc18h
l3ByG9lAYqrGukjZiygGb1GbqVEM4utpRMeDfs83M8rSUWYFmAVXDvYzR0ZvsEqB
DaaSrZv9DEB8iCzLPIy8jqjW73pfAU3NSzqLwVgiIAExqW4kTDoEg3XRLZGrKY4r
gskkcU8HujqQm4dxFLx8AEqQ0IZ77qZQeOMoYPuwnGgwbFcr6yHKRzCE1v1upklZ
XosI4hXzV9vCUmFsecSQlTQ3z3Si3aKjaoAFCBGK52MhxtcBPndEQdRwXSKVlpjI
QUVxnZojW0zLWEZQ/6ZgzwQlC1V9hQAn78YFRc7pVHSC/Hg99tO9MOFxwlytfJ5N
Ae6MseJy8rVm7qdoDoG8Uuw+KT4t1qoC17M9xzWCZT8u2KsHN4c3/bNH5wEjUZ1E
7u3GraOGNWD9M8Pv/UWz5BsxBBKF6jE6bOQtG4lOYXMxPwOMVakKXmFOnskBDolx
hkKxj7fQfZaZ4oZlNB/CdWy430DpCsgeiVZVkQ1wbgd6hXSz9gXjhsuCXkskPZXl
RVqMkb/5u5IxeW47hJZVBuonK9oOVWHl1dFYDwkJ5xpU4wZu10dUEzDwQnfmjGoo
cxLsicryViHLJgJ47ThktlK7qFkPGEimSxOWqJ1xDkA9QA8pNfPbm28PAkTLcQ6K
qNZjg4Rto4LNxmxPrF2/6tC7wuqdPWB+657wKmmwD9d3qmRuHbW3jsX0P2uwLpxy
u0KctLBtiLJCuiHLnCSh9d76yENrMVaH1/0kAX8RQDBfKeRMLlvQuzC5KsMXr4wd
pcRvc0kMaTC+1R6id9FkzigeGuwfczkiwBw9TSQ1J0xflVvwPjuAOhYTDjvFaiie
i/CEva8FE980QighQqR1afl/7doXMizsDN8ATuX/Xo/qnZ5SqLAf7jICz7P0b5O9
OyDZOQUyqMCzdIAWjPqqAfILzkjtDFnz28KrsAFD1eLN6nxXUKCLzktjbvsgBRrq
HbVdeL93QSveBdmOYRAjT1IHE2lEHPKMnBGoz+o0Fzr3tvCCECkFZu0gchmBtn1i
uGn46uDQPp1TeEComtX8DH+hRaWwadKabcmZhDJFuzf/OB5vfYd47iiKd6Aemvkg
8F7V40egH6Kig7S4HIwjLNgJdk3+SKXNDgF0ojNUzq7oAdwRDLBtN8wxv19O0ZUG
iDMXSP5fB0VlIEePEh6xe5+RrQxMPabXqPhGJ7SDg6eP0fm91eleUfej+ohRyqro
Q84cjokRxMXB1FpknicuxlvPWCkgcSHiAAwF2m6dOONfK01BkTJ2JR8VkfUky64k
ur0CoRNlawD+O+k6OymowOiNON4KPh0CxPM4touJyjlb4rDo4kxB/FbjlpJHgy+u
5O/o3tM2DYW3NRP4W+7uZvXEZu75wdfJ8GtRdsvy4Zu9JC92s2bmLl+GbyG2yR7g
vCaX2LEZ5ps5wLZGk0pzqv6HO43ddCuI4ofgGwBy0FXLSfqnNn9ICB7lDYb1qRZC
Dlgquo5csbOeAqoCshnCQyLDxPra9BtNXEcP9m0+yx8mC0KljuHbviAIPAqv3+O3
QKo9gmv/bCmPWX1IpyMQKCVPuPh6P4ikYNsCyl0sfmBrbV87R1aVOS0xcEomoJ5A
Ayg/DA80H2JQGC9yT11YLO9hXJ4ELPSVgnP/U8ZvO6NzqwBcM8CCU76/EnLMP7fi
j72atDZDacLlte4oZAhPaI15EDL5TeqzpoP+04oalRedg8YKQUuz/oqqZYcO/o2L
UMlHeQhsqPEF0KbONRDOK79/hifaYeqqwzKHGYjzih0tXpkeJOwOVATJPiFQUZZJ
D2+WbMeT+3xKFksT/dz97fq910OqubIXtxse5CNg/gWglekcpkK8jXxMEwY/IMc8
Pit2sPHzYuc04bIbMap/2Agx5dsOX6QU0Yx9muZx6A4Xp465jcF5UkwfdYgbZskd
4dHM7+oBxzAMsmgaKbbpwcfg4vfQ+bs/rd1x1WOj687dfeTNwWUWqnAIpoJgJnL+
tBEaxaHyGO4o4fY9gDCv0/ZlFc3Dddzhdk8Zt4utAFzq7PCzNI3bV5RW3//No7M/
cPMpKpwo3tI3ttjwaRFlwaBaO4heZCsG3yQRjXBQjNd6tfDt3b4CNhcEeWDr42ks
4x5+8DCb/FNlCpxntp5aqSgaodJH0pI0rgZoQKBCcp12rH4KJpfpYkATN6eAvC+e
kWYQXoEeyPvwE+QLGVNlR80e1GzyR5aS1vXYe02bOyQdiCHAALcfhCqZCWT8nMZF
KkOV8TVAajLMWGPrLTlD+YgIHbVrCv4QNyXWxWzDhGHwcHZEWQ6dWDpibritp11N
k01p0343uAnNZFCodF6wyvJ500esCWi0D1xs9QDP4CLnL7YFSOM4gmB66M4BzBgF
clW7Rp9sFO9BtjSQOPJ9RPSHclYdZ1U0/koBlW/Z5VIqTCNLkZPyN0939W+Uw8pt
MnW0CXGHEVpo0AAw7kn4cT+By8uFfEXLTOG6x5h0m5F1N9Z7TIjq3+j3uJ0O2kEO
14VT5RdsNhxilb+QYJk6cDmSugzONWI03r60XiAKFyWmgUBX6Y82WqSF/XVvxIBy
YyoW4Pt70jo5RltrgYNdXxI6Uk9Fqxe/we/Vg9ISKiY38EKnyNQBuGDb6tA21nyY
xMcIei9pGzHby6iyU6zrSS33oKU3HR8IiJBVY906cubF3DvZfxQ2CVF2TK6yuoPm
D+1MgQNgF2vKJ5Hut7NgbPwtflQMp64/pkIenwt2UYy4Yppuyk3B4fEkr4cIfz4F
HtQimAvuDKxE/fuZ63iYcWGXA/EkKsTEO34AihyQV7TgJgD1TxlvEG24Ujk7c7pR
FohhJ+ZGwb01WZQfWWTBoAW/LrAbqtpJ24x5K/UIWBCZZ1slU9gXaqgpmXCOO87A
54QfaFiC06sdZUHA6rphDGXaDHau3oYewoOK5iSLOSRGXuVCSg23dKgyyOiy6vds
xQ7yYWTX7e8ZYNYISkzH6AzLV34JLB92VBlzGDk3MRnXavzBWALbAtzPqZnN0Kv6
Tk8gV/0CmmBPoayL+lIy0Tz5dGttwyZ3ER4wZ2nMWZjJT3QH2HgIauh4bJpPmwxu
3jtBScbDq5yTV1tT7Jgec9f9Emml0ojpAT1su5DcrVNlp6B2ASz3qtyJXPZw/Vdx
2BBdu2G72gpiGtbNu6cx1IXwemxvSkrRq6MBFcSxIP722lI9mGEMW00Sn8hUp4Tf
SGkfRF1pAVUZLFDmjEeC2pnq4fdXuIQhAFz6lBHXqeNqemZK7a6fJbSeQFJfg6v8
TueuJECaNgev4cMMs6wIA+AdCxml2iTPyV/T8rgP3ks0Ko5GRR+GTPLepGuUQPjU
SymB8HSA1pjRkpcC7FzCZghVxS+2GhHjfAgleQof01bEzcj7ylUd7OW+mTxh4no3
YTQgW86CDvgA0NbsD7dnGwFrBCa9UFkgO9FdK8UbA5Rc0Zj5rzmucWh0maOdrTyw
ex4wLBgKrPBzHrgcrT0hlgwciKkx6Rb1SUFyHwf0nygZ3KZyRP9igQ41NzJ4eAfp
+tX2/9T7Ycn2esEfdB6ag/wkgynZnDR5drVThXJgGTxbvY5l41Hxz2WCOMNgzLIj
7SZWT4CSreQQWRt4gH96S7lM9kGJOmXy37ZR+rjX99W3hBfFlKXx9ON75ZSQKEPX
KwYX7HkUNRxGmM5cdWOjPo1UkXS+9C+ZfynkC4w5fIXvlz2/bulltQzsERuM2tbt
qzsc3yBn0b+5hnXxslpUVr0qWitcxeur582sBtm3iBtuX6WaRKu8Fm4/9zbyGOTw
dfalCAV+VjvdK2qVQ8j9IYRaPJHC6zt6m49eqdw/t3qn1mqeKWSoTbTVtyjaOHbG
yIcn99QAFoN14OzBVq8n2Om8Yle1br6I+8SklZ4ZboNsrbbw81BQ6pDm9N8g8pUk
TvPzob9iz/uggabNzX11qOSneGcbEWAtVMhJS+e2HMxSnoUlqHlCGlMQ8/Yu5E6l
lfOkr92eMkX+tz5Hn0CzBI6Hnlj2MuHqofve6Te9hjaWkdonv5bT5ekgL0YGmKaY
cuGfSp0aS/G/qfqG+L5xwgr8Czn2id8n1pUzulfOZvScKT/uLBOCVzhShzLJjGzT
W1+XZHL0jrHrRyWeLChI33jf/1qcw9+G+5VJHPW5QadPCS4W3kEP2Oz41YAifTqk
8apzNIE3erSWYt2lOAkA3M7k180AhOa9ZJGwCDzV0EtWCktBtsGVuKLPKu4BFm+A
0SlGgmOa8JUJUc3yC23RexP+2LE+SYsGXJNKShrgPVu2XT/CKWwUxanCoLOfO6Y9
SUnUUkyTE9K6R9oKIDOs4NMwSn8MO77N4sZ9VniBDxb+/y+3TuRl1VEdv0anUUsQ
VQ0vnnbaBozDefSBwXLUralmqwzJuzaBtjJKJMzSYvtjQXxhINhZTSaOmJEaNnch
pdF+Wmtlu4D3Igy/ZgEeaSIK5dj5pDRheWJlTXP3qV2lT32o7WgxDBXF369hHccg
wPmA8IKuvlTY5jDLCfKUrQ6I6F5uSIktbZYd3NHjS8hZ4CZDr8KNoLD0mlQkyc3U
/YHSGIL8g7rVR9dBrZ2U6sAbYGLnnP3/fcC7IJcqGsjNfP5rzgGfQWAZLOe1d56S
mf0Aj5QCgzKkfAcme1Edvj2XtKVhAVi8nFE/CL69KIJyOqhRV+I42baxQ/Rw9MOU
H14k7Q52M2mofO2T0+BJq8U/eUnTvHo8JsgrIHgQ1xecu0D0+z2Uol8nFvCrvmhl
0svmS5O2pv0nAvL+/0gMgHHlWrrEkUat2KUQOCFYRb08ork3Y0CZ9xsRZyfM8VXU
BbKkKqhpm2P1SAYEFlVetkZ8gE7stqf8Ud7rMq8Ntqz8V+XbqjcXATiWC0TBLnhd
mPVAuuarMaXnKqyERR+Wjw/MfoAoT97K4xLmHGSAXziAClQmOGuU2Kue2QSOhaj+
cyBkPtCrHwhRDyabX9CGD8hJaVQkzD3yRQd/ULCZUZwWOOsb9MOB5w6elZ2a+9w9
wp1wyek/yRoYQ59bMmkhEE7LqxSiARWIawggelB4Jn7apkSxpvBg+4wQzoHpxAFW
KAHVO2aTaXL4uM+AnCuGCgT4xbwO3rbSiaLsdzKoXIeNdZIY5hBNWpko+XVOllpH
6Ghyo1qcA7HJmJrUQ5O7HhZ4j2EJaP9l8NZ46PizzNtWStsZ3MQk9fTN5BGwMulK
X8qX+TiOrgNI9oK2CY7YvHVoXjfeae5j+fNpaHkpW7llSaBllR7UpJwtTpr//Rdf
4ktuZzIjH0eXQVO1Dpl06dNjW847TbZ08T0JwBJHfx+aXu7rSzQiO9oBlc/rKHgY
v/SnUh4PcKg4Y17qfRS0pha+Lu8Mzh73jsou0th38iyJVm+W342y7/pzx99Z4B6g
vLvOMSUWhEtQzAvJ7chctDusnXqjJYBIW2CICHWyBi49HRvIopRlFiWS4jTLV1Fu
W4OnK8rhdfB2IMxSEbc3AYSarvjDp/C+csT2Z3CJYCvgruHqxJqD64wBUMaQNiYf
NWD0R38ZURmnThm+ORFFSsbBtWyhyqalGAjXGjtFDFeosjt3PcBch8NmbcjxnNj5
FKuk8uhlj/TbTz2dGa80dwVbLLrg+EYxvM7mujnJQ9qpiWXNPjE3WorFO5dbS/DL
pmStVZouA+1WP9z+hFABhBqj6Mzf9TQ0tCVwBnV/9qSCNOo2FkqSF8bVflCLA0XX
27EDLqm3OOZeM3GInFWPuy9son4ZBpKMjXRs+IgEiuZ6LOfqleOGpzLuwVyat03X
LODDVxJikPI8bVBR4Ku241ah/DutVTkHQUwBhpriHQmwa9a6khtbUXSVC5uDyGpg
AhDv2Yt/090tNmvESys6zpUEL3qNPDlNH+trHdfd5pw4DuMKN6/c7DQe/ej7TQSw
qRx+Bg+/mU68SSBl/9FPYhDNTyQmr5aEJYSsWZToPJA+WrmGu/+DqsHlFps0pxpo
fLtjjyjwjsm8ub0GwgdLAco3qq+a0c8+zLeDQz8aFEKAJrVaV9xEWI6Fag3omtbk
kq5sYRWcc3RMFHSA8HJMqup1gSOkBgWsmuksFIYd+h/QpfCqwKbgunEDnz5a3l6e
9hfPMUEuD9UGStf+Hizby6Y3h3TVGp5uWBlAwPLUj60il76QTxXDHw2X4DebIhNB
Xzr0KJV2xnfbDGG+kw0UrUJhj0tDpVnuOiIKfYTxcFHDOMPHfXP6F/u8zjspsjqr
MawA5QAB2zhUv9tzUWIEz3O669fgVmWt7dHu3auZMyjVtkwQUFWfHaAbxCU7E3j5
M9sS39iEr2uSOq26y0Ntxv/fg+IYjHWRP2hepwV+XB37XL4Q/EaMecV5D9mSpZKT
Y9yrHyjleZ8azXxoYOB6O0KzGGhoTm3vhQADBapEvAiof+cno+TuyjOtRrsbV31P
puLpn6vtLAA9LgG8lj9D14WISyxSrdKzCKRc5a6r1gE0Fv9xyiWaakbEYq6FD38x
J8NRA4BJtHtnJy1J9bV37zWtUDx+C2ZQ7Xin1G6puMYiySxeYxgXevfWut2TjIZK
MHTezee6YWxCm5Uj7Ef9tYtENiNRJ/9b17B+E7EjVQSq4Ml6rk0CqI9VI6JB1Wrt
d2IIKa7WSDvhCzhUUmC5AZ/4aceaOmNITN2lXHLzfY5nhXanIRqfaQkv6sGI2/OM
44c6PgJARwqi0vevtWgKF5mkRcf4Og+GwRe3o7kfIdsm9wPdvoJ646c4AcNsHd7p
ka5G4Vvs2JiMupjsynVYlL1u8K4iOTESbLnSk2t3chaw1//Ezfg3QU/HzZfdBgXS
K23Tqm9OfVcPX9h0XqEsJ8kT7IN5vKd7EBA+Qhg4jIbELt4YoOUlENKsML/yXh9q
bfqQSfVl308R9w72xm5V4w2aHN5R8JhvhyDTYc465yDArFrlRqj2xc0AU8M7RA11
FK4FwEDyk+Opuv+K7Os0GTE6IF5IhhHhtZuO70CoDH9g/qDLe7eQaNfB0MVXFxtK
p8QeCpq3QNQ3jf4Vrhw3yMCtuOqn2j/LLH0DmhG7tdd4X2f9BJ3BdG5OEcOYGHlD
aXWsYXInT+qPi3hc0zsThr4OWy98XGB0yBd2yIuQ64KGVkvcihywABfhyaeYuTok
1SBOdc/HNCTCzB+w3O8fVZcP91cjAQDzu62LjRapTLjOE4/kl1AB1gXkMYp4C0rd
pbFarllpthm7KV5vi5ofKeGy/kmu79MjED3i+WriO/TyxZLZAR82L2qrcG3ebRK0
BmGa3mL97+NRDtP3ZcjCKvVJBu5gbi3B08iet7HVVKKaja6IxMaoVXrpbZcMVbTI
U31YiTDdqLLBRUfHnJZFJMdBfh869W4wGNtCC1uPXGEHpjR6VY+CWvF5aDj/w/9N
DbNXkIwwLaHvhp+iYC+eAPtuKYPimhyzniuVIabkiJy3HzRe+w4abOMQWXLS/6+y
WBxjKAnZxBfpEALJQUomsecISbusSujIV2CvtDryJImH810uZtvwXid2ZODHXCYo
ZM0jpHHmvwpUVJI5if4MY8jHY2W9QMgcU4wqrXlpQOIZGzpm9+2KuHf7H1z6wRP/
U+ip5kzAywnO8mhCSM8LWvEQhYBV8Ny9/ZuDBF2UNHkW9LLO2SB1/x1rx1SNfYtI
8eZf4j/7QVipI1toivCXdL9BSXintbe+BIuPFwY5vOeILxpChBkAZsHYLS8/Ugky
OeXUavII70bnPVpI0qFXsTOUdueHv+rtyoVDsjmkYGPghNIlwWZoPk6ro6Oil8cr
mKcGhlLAORsiDAS0r+GFtK+T7JFXsReGs5ZjzW5oe9qaCzpvnXxoIMVjOsQi1SLA
itVLHZvSuVrvxdjdwu1FH+KTZzE+x/iS4RNM2MffVvdgw+ZOQ17R7mAQ1s3Qz1U/
1Ix2g5aTBGJnt1t6WsljDtqZINb6RqUBco0HjyW8w1zWO72JSZxeob9xOI7sVD+o
m2iMl9hLr/NjC7p6TkaNKESQUTeDFrB/wCd2XmEhQ+N+oSepTL8r1f/TolKso+vs
ZK6Ffec5Je4mdMVTgKgTuoAgkWNrQo7FRvmvz6ww5UwWhRY//SpUpkSbJo0bpKGL
TUl2hpxoMsdoRL4RCn0+x3koeFr5bVUr2Mo1PtTum+mWV0uUWcRuzy8Wke1DYHzf
KIS2G+VTzuen59OTM03dkV2WQ51JjtwYRHDk+bshnJocFUbdGN+bIT39peCkU9Fc
u7+XTXF22lRdWD+he3m4uDtv4dK7XV/pobW163Pjxi6GJPkMTZHNXeUV9lPCj+Fl
XcgHH34RoxfDdSUEL0nRo+cEJrchfdQNrQy2JYCX9+31i34/iKcT96c3xYk4UfWa
p1IxtDIrmodI8AHauKcrNxQEmIZgr+xpBnAeV4vshsq/L2P2Td8etfwgf5oGzuZa
c6s5kEi3HnKd4W/fqGWE4oIVpl4b4oAh9R2aUWaLMHKJt+uBfjTw3q+/k0jbwJHE
Rpy/rm40QmF7QTZvVXrMcG/BtaJSDbzMr+ma3iePknm6lW2I8Z+z6WwkU6FKm3PI
8yn+o0+odQ2Qn9iybIgtHna0ZI6BE6tPgLSbNTpOcDv5M12K4gl0KklDrJDfMsNV
bLnTgHXMneiR49QaXvHWJxV9CqGe/GVTUslXj5ckGMfxhEJLmCV5KrrcZ1SSl2P1
Lghei+MJ0VHnTG9wgFUsPi3xIoUXkEOCoNmreDpsjP9RLPiiChbmIa5Wf+aWb3+c
wvhk2S6po/ySquLj888YMGdUmDSGd0HglWsGIG00n7C/Rb+gxC2mhW98RSyePCNv
3/3qspKwwekCb3ILaxYPU7ubQhdGB8jrNJerSY9pl+nj5EAjMHndwTPi01nVLmvy
GAT5OQtDhG1h7CcbAwE43WdHvuuzxBE8hSSq1hx61xngVBeSg8EWI/n9GRRNMjgU
PAPhZfzJ/NYgQlvAQjFEwJKMsOb9ssapCYsiEYYAPZE8D3jA96P6m1xgTNizVo0w
GA8L401LNexkJ0F0Es52A2BqRBMa7W8M0sy0JkmEsq1+NUBcVfGNtw9eT6FBysKx
Jp7rdN7ELoNV3ASBvq3KHebkgcn6WCZ4gpydoNt83m+4Qck3xUoyWSIQ8dXO6wUv
SM1LELzB7/hQxgkS5ILKdmFJmrCbJC/38ckvF8YaeytEZ79OaZJ8xqAf4zc7SnWZ
iaa+QvJkikuUxFOMsMnGyHOUElp1vejKPhFXLfJVwqs7KRPO1a5l97Ur2Fkp3Li1
rLi5hLPIVLZCSQOihgTZipKYr5XS9JPD+otmvU2g8Snfafei5xOzcT19WLdFF4PO
bVWVXaZFIPbhleDljRBOThR4pyesIqbGwGhoI9dlfQWV0GPkw8rLJ2ucRA2OaosQ
W/vHMWW7dLNuBCA36RAUIl9saXu+BGrVBdU8+IyrHTiPKdwIrddLKDOE4kuGGO3z
UBTSt5C7yGQNIh0I3y4geWTnoJpIq+kBDbqn+ohl9t2GtAIkKyWdry431GfWM6MM
D/POEr64ztNCofWEVogOhIZyvJrXgOwYDRmdZsvrIEKxy+P/+Ws78ykqOvecO4kz
6GNDjKvbVYu9/bT7JdxThlNCzZtpFwdpl+0rn1DL+UOx7EEOGlhvPclvvZ2bJFqy
rHLo8SmBL/rltLBIj/a1/PzJkY7JBPUXpiv7sXaiwkKTPF04gcJPDYNhUF7c49rm
Q0MCHvrQzGhzo0nWBHqvE0GejniAhyFmhaPXy+YiHkEbQbasDQBaioCiuZrRsXdg
/mIPx4cxwKs7vEjAk/WCqbbTnXiFJw/C8NJmtPh/6Y7GzY54RPvlp/xnB9bQInu6
B6mj4cQ52WTWw2auuunw90XfjPlTDuKGifRlM287TVem4/mXMQnwNv9R2DSnJORD
6jFhPlKpRpDA9NwpVHDrJH1yah8O2eBgs0Igw4sqREq8zWb2BI6L8fh5nA16KLpk
9aoWqzQq9SAcQdHE+QWjp6j7EBeFT3q2TYswUA5M651958XpMD7nwlCj6Toafz1e
K5mWENuVfDRZKzYUYv8N2aRlgs6WfdDgfii17YfXxHfqD6Yy1JWO44e/QfvEqPEJ
q/7+MAIDb+pWbZJGpr9nwZGw5e4vIDwa75VVliNCP8YFZAsvMANRR2ihUJPkBdaM
zi72lEST8Q8S4HwZOnkVRW1re260ZeDmt3OeuFmz9YQU2ND12D05LVNYudru+7Y2
r3rHnNw3s2OGATRdx5kqrwQ5rAOjOLLAJHPEHJu+GAZ7NEIkjnr1HJ4FPefbFCn8
do1ddd2BstLHBCAYyQSAv2jN7/+Q/D9ARswTsQSV/LYa4cFdMJp0w/VKN67oHJyL
KpDU1XZ/TTAuIBROb1vzfVxuzNaVfLkfIsJ2v8l0AeBrCn2E4dEL16lvxs6f4B2n
mNWZhdcYbieqUTxSsCrnP4AEf7zr4bBsLn9rFmxNdYDohhz6WKYDcD+4m+ySCqI3
R/xiOaef80nSUWi/8xtuPr33/arubcbA1FgQD7GRpxCDh+Hq/aCAQtHAay5uZpAp
YGBBhuXNX2yy7ppDDzctSFGJ/T2HhYiWKG3LCF1CENU6LnZZRUuk5LZLaUtWc8ae
0h9xZl4uVRKr7fbST0ee+ssTmPEe0dHZ9XkG7Kajxi3QzSc8Xifyu3dBd3lXci09
Fny1F0bupRYqTeU90hW7la4ophk/9tgXuQAy769SEuUV1HHZwL7TcnIcS3qBf30B
JgCXejanYM6TtenfzmKTiaMIjQdR3dIEZvp6B9PlFdohds0xKiBGwXp1Ymq9aPPp
WT1eD0G7wyvPySxJDWaqW34mq7PE95qj5geRKJhnvuTFS76i2fGYaR3MbSYhpXPN
Ht0d6+ho3mHdYKdepUHEFHbsceDwykunu3OpJskwxWqHphX45O5ApDqjHSHQPxu4
8pCFPEGZOnJTHifI6PWVO1vu+411Ol5l5YzC4NMqampvcGmNgmdI8hrL8h6SktGB
rE0adBDgQInvIk0Uj1x9LXIJUqwQLPWE1JaS8Y889sPRT1bF+Lk9mDCHMcSHdRsz
EdvVI9RPPvje/S/bxx/wkxFzbTcd9ISqEqvTItEV1TIjZldSugWW0ChJvy9GT/Fu
TCwHzeSqCrRKVWgDp/GYLHseXpwrWWcI9orisU4k169IkJliVmR2d36M6IDbhapn
Jl+VMN1sfWeKkrN9yLz7TyueH9PRHEx+sD5wPS1g45wnFehRoj/XDn0meEBjO4aC
MjYH4iY+39Sh553t/ckTkiC1fLIDji7qX64ISxOXIigRJV/9R4wb09a0Rb5o7Xv9
NIYDEFstFTCi+pGyNv+ava+e6Tz/Y5SVfwfsXjik8tMOElFu0q7YW8768/CMIUb0
cyjOkvdB95JDrVdVEeXwLyWuJ/qbJHYZ6gGyzoE9YrMWhB3+xeaY7kdjRyfFxP/S
lPHaYzGqEZseZYxeEyKyJkE65IK/vy6xTE9nqz/Ha7py+Jj6nCKo665u7c+af/UN
daQG7X/HU0DbRbGmH3k7YD/uuF+eGqOXncgQXJ0j3VciURAvvFpOucjXB8ZZ1jkU
TVGj0W12ebPpFD30cpXAw+R3DNsAIC3r0O0pSa4To2s7pzPZJ6bTkbp2/8sV0mEJ
5cOAQUNDwwGsJHlxyjr3cUTNGdRAQFFw08+mEb7JkZQSKLSz/WrjQBZWoocT1vrZ
Ls9prhIXAVNoVRagN3UPcNN6TaUvae+JsEcqtsUpZRTVu3ZJN6nPGXacFgNr1Y5G
kRnqk0D4L2vOZmhfy2n47P4ftaT6qAFonFUXQ5c0c5ooeD6NOvfzHGoZmqBZs7zH
cPbmiqh3XIb53oPN5xEAx4lSGvItW+3kG2mgSq3qrzmvBFFbCRnF+zQQZiYm+luS
0Nz7QTunAsYgxOGZiB5K7TedIMUvJSldhn//c9B9T5pzhZj9cLxFar3hxoQe/FLK
qpsBEV8F7KJBEWrLVGA2IY4vVgGe0TZE0RevYE8fV3yuIJZAovcm96ZfWwDKAl7F
bOmQLpx0eX6gKvmjacdO+y1t6QOLhB5ibhHxkKplB/r4AUnAlFcZc+Vud7cffVMa
LcP7lQ+/LXwhJz7MzIgjBg71ZW4tRhk9FZYhuZVvIAm+fP+SPlIG+aZ6txSQcOlv
FKgUUclEy/gD1Kc8bc96oZJm0gbMeSfWRUp1m3gTlnQTHTj1dbOB4kZZY2TO0RVi
71pSEaNgqH/VqQ5ksgmH27DIY9HYnnNHzSfwsy7dw8UER7+0BoURdeoL9NU6Ipew
2+uyk32wI1mmX1SilwM/ovV18b63WQCaxUgNLkN6v+DY/2m6x7HliYbQ820LRDDK
PBb+2IEuM5UhEOZAoFP0EdOJY7kbXjH5kAHl9NkLJOcRzm2N26vhnOtHLRCNnfs+
93uQeeTwN9yO83gbpvL9gear6Em2wiHe1AGhmpo4fojk24l3Y1LCk1rhjUUlRD9/
00pW+0dEZsgjg5o3DjfLPRgDBMQVCtx14n869d/NbwqboXuI+/RLgAPmKZEtr8Ue
rx2w+O3FTvN8RLx2cRzLQX93CRAbObCevpJurF6ASmpd6lD6MWyyop6dMzg22Tio
FJT5C5Mx2AbY7YCEO7SkDhmRKWHDHEJKVmLfCs7gfYnjPEtn3v9CStxCGk6BY85D
DFa9Qqz+iWlxoTZxJVw0vl9rQASb7YVlOzToU3uKNmyUvfngonZ7BlRphFoXMiwh
EcrrWdytolQU7OKS3h5yfyqwpK66xB/6EGpWKqegFJp61p6DPKntgXOL74viZBcw
QNfruY4liCwijSawmPQ8y0uTj8H1Jlq8Jxr4JIEvAu1hYPaQNC3u2WoBH3ketu7Y
yOtAmUVL7TfKSJc4UlHaBYmS0qe24URPECdvMKw9X23dfw8/hBhLy+vE5vgFwGrW
cjrRde/vVwYVtEq/MaNT4NHv1GPLIGDGFmauq6yOddV1ZejgwNj707GFLyW/RY5A
LGo7abo7+Rw0Rbpms2WWogeqfH2rS6Z6rM5I7ON3+VlL3/Cy8lbHNoUumq6Cdc+y
jP4+wEQqoOhg+JQOm65acXBPjyvQewNTfK5bLtxytBNFbeartwLSs88CgLUOfUMw
b2yWMWcl36tHgSepmJPuZ+sXxpftMkQBHCBFx5t5rQaEjyH89i3L9+HugI13VeVw
yqKIR4AyqBqFNbQ8iODSrZe8xFkN+3vKtrKGPrcXbyDYIy4TGLheu/Ied6vHtj1D
sgFqVTeNYKP7CVP087gGLny1yhvviCSX5hnApRdmhKid6R7iwBLCJcZx687JmChI
yZGAqwN0oxlvb8Q5QDBjtM8C2t7fgZ32rHTYHz59UQ3GWLJXa2sBltc2Q+xaoqHn
xWBid1G93petfRvAluCRsfz9G2pxUjr5WGU4TNanj+X/AdKMsHdd+xmr84ag9eQ1
E/ml49hRGCBrt4zF4lGyA3TvKKBIOcLLX+034PbeGTke82+vkt9cAopoamuLgbT3
E5FlplnZiM2sSo7qgAxm0AQZnu/8MJQ2hgO1BLfMo3BHPfKZRrsrPNPq60qy6Us3
GbKVjm/vq4jtcVtqDDAYoDJEi1fMH71gqSMiXepXFOpfQpO18wavYaYxRdb8KVb5
+VmBeufqAxTRe6rLUXiZj/INuzO1dUGPLhmQk8NsZDqo9Q6pT/N4V6dDdd7oebEY
Hcr7mJllckUKtGfiHPeZqPH/tCfpZlvKs0sHxCwkrtE5g/zIicXxHgARR/ZJk8Ey
XsjHt2mOz+r7K/epnn6B5wpeZtfzSmVIf5sscXmYZzhBO0hdjrupvEs/c369QJLn
ch1gzwb7jV0q1XFQ/fpX4IHPNETk59lXCtd1vnyqXswf3Afps5+kc3LnmH/8ArJN
fS7+gFJH2KZpy9mTHbpG1jP/Py5s1y1VQ/dbIGCihR4cxLwE2DqhEZaH0kH9oIqc
XegtGELyNu7EDu9yF4KVXtx3mUL+sHIJ/NK5tTQMF+lKTADMwyDZzdUV6RetPcLO
UbCa3lkFVBvLrkXdBFoFMWDWb/EeLOmvGGBm7nKqQZ5Cu8BbO4RcOVLkNz4AisXO
fWlaSfuYhNOUAtc8Cxq8hr4tJQqgIiS03jIzIoHb0VwpVrlG4soMz+novvqYEs9G
VHlAe2YLJ+dnOkjFYiqQXx93viTliDYdEtNYkcZ7m8dtrB7FJsM/rI+FElD2DbQ4
EKH2fZ168lirto5Rz9mKbVb7I+ye78Aot6qctqchThbdCwVLunfV3geWMJSxGHUZ
aI3avqNfledwMxCWbsGtXj3Pod4f2U0v/IHBRtBJvRMGPYA6/cWs/EOXIlqScOf4
ryn4MNhsvy1HVs2Ccq/UV/Emgr9fsxPZUW5bHO3/+M8nwCPLR/crigM8U+58wP1g
ohOtaVFOqOvcMeWf/aXhde4OhCA1HMT5gkMpR0T1aQmVvtODZKGYtU4uAAdJG7Pn
OMHhMUxpMfzy28UjiJSCJzfYJin25Yk5O+ASw0JUSvIzqZbNsYXXCtptOmzeAw2d
1WX1wrBanLC4TXil3YkyOMAa7gHl5H8ZS4g+3ThhNieswVbM8I0gOoXYPAUH/7qH
1hwYeWwOXxpUOWF35SrRqly9MjrYNzzsWgwAmphXMFQh9109e9Ifv1NSMq2m1JZp
9BIOPpEjbIbQpxA96TlbV6dgc5B/Qnbzf5FDxALy/DmRe4M4P4WWr9rNyMBWyu+k
flMUP2UGBZ69aGf96ZiuEuUSNiP2IQGAA9bHL5rHhHLFMlHI6f8GHnGZEHHVSk0W
l9bnVHJrT2R0cD+0+tMY1rud385L79WaPkrBADNctt1vztZxvyGMe2Zli6ndtn/C
EzM7848astC4uTNtLIyc3dj299xHIMh5ytwhm2OPwIRoup5JcrUx3k1FP2A/ufJa
YDuonedwProvS7DI8OPIVsq3vw/AYW3NJOvPR7eHAkV7Zu3lY58WONzbr64wrWUs
lQxoUYjcK26/NuDIlNSfrkg/Lfg+8AEd/5HNcm3ELU7CZE4/BhhZmnDlECRkNSyt
sICwWglyHXpa7OuN9nLRz1ZJSs9wH5ZO3uKoHEM66GaTKhRnuKVYKDVjfubiCG8S
zGUhjLtUDCG/gWDkfbR0eOIjc4qgp1yttx9bGtW7ZMyISVNH1IQ+FGt93COosLP+
j3tpkoPFtU3ddJu4TqNBNVQlU4W3upik6Crt6y0MhLlfVs867snunbmBCDq5vuQV
NPW8ibvEXvqd/BrmBW9QjzKMcLGy2k4mvBsiL0IjnHjh+zALeYg+2wd5L0w2h/BU
E8lu3X5OBbdwsigRqmgII0dzYl9i/dO8gU/7hp6A0lh6o4U2UR55XGF9qQXB5lrS
kpjwfYfrS+5FSyKPFbqKZXE8Ryltn9FJr634rXdzYgISB96HzIYViBz5ZvMr23Ci
UQXa810EL4WefvYTW40QkMaCbMx8fynmfp1cL6+xSaA5KT2H5fZxmLeUL748qfXI
fsIp3rk34ELI7WJXKBAdKn9KatYjAG74oyGKFDHrQUuZAHJIgTWR/fM3U1W6K4cQ
HES7Zj3sdv1BxKtzY31SJM53awKQ9uwkXxtDsYLaCIWqDpezV/2N+MKMbPJe/Gq3
8OzkfLxHNuNZII/zSy2Zh+QqyBLLEDPjjGh1blqOyobaeY+LcDMPVkVhtnuKtiDQ
iUGAYCskKI9DFAaMbIEsU18iKV6dWIBUI8fi/lKk++XCq9N8gLFiTljUKmXEw8Du
6UgucLvexDIFAg3hGfT0jBCL+xUowl6ONi9k/33JnryxA9ZyJ3ZGCTiZdSlobQjj
5GPNEVcM0a2ud80J0RRC8eqBHjmOsx8sRriL7wJ3MHsVUj9KPRVIIGqODPu/LB54
6HC/oqCR8XY6J9MN7svqU7aM+LS43QZNBcrhTqUPDye+0OcCwV1TE6L8U1j4cJWX
VjU6D9IyrH0CW8v1uupD1lhr+RzEkcOlwJjivSiOzc92FVwLcPN+/BD+08rJg+7e
IHqHw36to5rBxwzV0PWk9y+5aRzVFAQQS4I+vXU7pKeh7gflwl6Zz1HYGnWiKSoG
YcEaB5poi1Hps44EO8+z9e3fU5BHoMhplr0w4k9y63W1jTlnilXW4/l8eP/tZv1Q
P6dPtfWS7YeSaejByq5J7ImMr6/NXWXWKp8QJSEa//XNyqEGqbfKuSGzb5947jeX
udl497wh8Ar9sbYqXWwbNeqgyx/va32nav2k0Ec8V2fYsEXI0emv4EH4TdYmnLZC
vNZQxo+94DOH4eJ7qRveMb1mhaUc+K0f90tTZzCpE69xnrJJ7h9fupi3cYADvAwR
jCPPtgD+hUvdk0NMxzi/BAvSh+IDm24j3tEvUqReaUMNC7u6L4OBAKgTrYVJa528
Z3PyIrXsdgyu3MNsge9raoDcGC7dbI8MXyYzePghgU3fNPW+bCy4tUO97Ii95Sic
fdz6npzveEs1TqzlKZSHpnh/WBEV275RPVyYy8rx+N5AhoZzgKAa+hzn5fJ1TBdT
bVNhji89r6taH0+H2GuSmZ0KNE+693XuaJvctM4lAbmSJgu6Z3Gr7CWxkQFZoCsO
qnWgngNygGtCnpc8qWu3Oe6XuRlzK3oE7UaUm8pFm87nZggLYWJfuDevmKSdPFq7
U+E1r8sQgGXpqxfcCf+RwLGmYa+GWlwfG+LxQWe1NiO441xIjyk/wbf0DafxndDh
MJiu0WOnyIhWwpkXraULVEPoUzUf1zLM5u+upgOyT/xM5+RMD7CpLkn0Sn+t1o/S
RwQ012ojAPwH1Fdp652HsTfuUDtQX9zXQOVsaXcfsO1FsX2iVjkfpyeAm5dAJ8aV
44y1qNy1FY+2tiCrjLQ0g3d+zor+QSN2m7CxZSgT9n2jgt+p8vkCM7y1YNwPXcig
Jt+u87++JOf8Gi1L0cg0WVW0FuJ+hPVUMSg3Z/LRNIevpQhTyDZ6CvBDw7LbZTTE
olFkwCoOpyWdesaPE6xqhQqMKXUZfluFYsh2HRI2abGgw8soCigXwGmTbnj0yXeI
haqIuH0yNO8gQ/ytUVhKeLQCzjiU9qVlMWPSyWivY4zgMlvhJ83hdEPprOv6eqeS
CJQUepaAZoyirllGENejxSwue23eDkM3NEVKrGVLgAVtVGZxEF4J+dp1tHpZumNT
Vpg+cwt0a3XifRyEfYjTGvCruekT6ZEsuBny2Rd0qJpHWBmbfBckFOQF7969k/Cy
NuZIvruB3l3L62RjuX+2AhJsuCUYcP3LYfvXnI5L+qlcKPEZSv86uH97DNMO450e
nsTPE5XT69ZxY/TK3Sf02GcspqZdsqGSfYX4fhrH3GTk46rKJDPZjIV44/hbudH8
XMOqoQbS50he0Jd9qlJ6C4PYIuDWD7vf/djc8E5z/Y6lkjmoaMd72m1szlmc9kDc
m4JO8Mzw/KfeWh2KEsOsm34pS/L9tCtXVBiCkeFr/qcS6U+cGYQ1XMNJ9GtJJGxm
dLxqf+unT8xGjEIyAVZfTWEjKpmwwVTbdia8gtGAjYNdPVUzIgMJWRfZLSUZMFTT
j7NEx7ji35zWjOrJzGwGXYC2hrlTP03Nanfc4kZmkWHZi9IeHiu/CghFmiBsr9Od
GQO44394xiylAIFGh5tQc3jnuIyWW3k8BlxfaMKaU7QhPVr4q2ugDxwsY7OJMJZl
fdUVghXuzDrrcBkoy+i4T3Ro54Hp97yyNdyA5YubcrrpON2ZV7UXdmJSLT3FNPq6
SAlodVxCTFhqyq66kc2clBOzvcqPPiDUVTVXDEWivh4R3gsnqHORwVuOqsVp1qUH
UCLVewvpoh5XJGqi8/8CZw5ubF3LPbS8JdTn+NL7nwGJ30R0/2pcc4GtY8XEKacI
N+nOpMKxxHfm+NwKKR/Z5YwGVwfBFBsMiRxukGYej7hqU6tB170HE/5fpYW66IXd
TjsVdz3mk0SUK4rtA5Ysjs/zUhuqUfJmcxPZnPmaR9fkulOJd3jikPlTsGb8BA5n
n2nOmVxPzimxwhZjV2ZMrDJQVSc3n4ThGYdqex3npwD4aK8FaSBIP2p1164BG/Wx
/XXIuMMB7t3SXi/oQQexh7pUriArFMT8KRP/JKiQ+67QaZBUyke57o3buOfkxrcQ
Ps//Nfb9U60ryqXbwUEYWs2K3mnXZhOtxyO9thMm+tFyK+bFj8K3cInrihQIEuYX
gKJHdrzxcrV7GgbllC2xXIONxN174nmHRhtcJEAQe9mEP6yU4df9kBvLlAwhhQ2o
/w8bN6db4A+bICWpKxMVrEm/rtWXRDYDwXUpZCEz9LfPY0rPi1pA1gyQsFpVwexl
oYfPlkHbPKls8rDqCVRzYQvLVbUV81u641r1lO0vFMwgEVTUT8O/uUIjdbJ+QmAJ
mzP38Aq3XF4aN3zl+pCKan8cgXaSdBrZUjiYvu7TX8PZ1VAfPe/NN31WN3iAg75o
x2HI+sIsmMutmR6aR+nfG4u8qpKy64WyIRJPHpzf8s8x0qi7g0kfS0iWaVQwaNhy
7zd0oV4s5ryXT7qh9xhIwi4Bm24Xln1yzMFv0QRDQEHb4TiIuNLJi+9aVjR2OM5z
ZkdBESHixwLdCYqdAdoC+dGwXGOiWO+kx0Syom0qwiQBCMJgD0wwBs71ngyzQrrk
UoTlghBLYkeZ46SZz80/TC+NFziOFMzmrvB48kIU1mXabyS9bQpLNuZQlijI0N2F
NZwCEqeBtgQxxTtyqdtk1+Qrmt7FZ589++egg8ydR6swJBG8W4h2PSiTftsCrepT
hgutqWtXIZKAIVH8b/1f9bCd15+6fLgvCrGSpDCz074iTI21ObiI4A1H0VcLBv+5
hVfRLbpLywFEdxtVydNO7vuJBQIDOPQqWejiys6W+mCtuZ8I1tuSxfOacL9CG8HL
KyyzOYPjmokcAclwAllwAV4GvtnN4puw/OKaiDC/ZnP46/RC3YB9Qo8cVa/dcrSm
7ZTE6YROBabJ+iuhr1lQ7LAEOChtkA2C6P4lrpLmP1Hm5vpeOy10xgW0z4eEZb2h
BuOxreA1US0fzG9uOUQkfascJlY34Fa4xg2jXeEUBf3dqcRzhYQGCgKohqkF8Ivf
Vm7jdU9VzDyswDTOk6zr6q2+b4pBuSvNtZPo0xMChHxpIzx3lFZXQeSYarAvne/2
t8dDuyoFl70qD+yu0qgf+ai+HnVKyxTcMObBZwLjyk/aewPRezKdQhIca7NchdN4
LqmQS/EQYH5x7KcX+57EjHf9MrZlvHNxOAqbP+XoJeJIKYb9nWLrnHcw7nGqDC1H
F7a1rCDrhD50fS/KLuw4RwobMW1QQS8dfhyP9HjJFv5/PbejxCRO2g1Ga194KeXK
tD5PVf3RvIQUww45uy8tAHdqEp1vt9I4wMRayznSQUknfQIWOnSNrH83jLFjtXJ5
HnqKMGdJsJToZrb5KiXLvKeqcEkucGTlH0SQUJdMalqBcViGeP+kmEtvc/VnMIjG
IoVPWESxpmYG7rhM6noDGC0LEhgFhkPiF/q4aiTGVoY7lWJR8KqXqDiaPtqCskEY
00tA34dMCdwc/wnu267VpfHmAxHoQAoIqv2rSICmO92bTvu05JazuIEbPEVtdeuQ
jhxs82VwDvRE9u666n8hURmNnIpUtsWGTP2yDGFP76diSKHCZaf9iqarVoLTVnBT
/sGNSBdL7tjOa/ZDoYxnVoE4fa+krlU9esOrJWHm2JE9H6OGftTbSCUGiFjt5cj5
f6hVnIokOMRUfsMY8zfhQpyvY2iXbDyXJn1Z2nGkEH7HGWwH8VU3DSU8UQcE2mZJ
KsK54eVEE8rBpu90aJo4cQya3NxNGuR7VHL+d832Xqo3dx+SN2vnpyfJRq7PkSpQ
8CioXdxTLh+CSfc6alcGcruQi07nQYbPvREeaxujCRAclPTHa/FfYZNdsG1layIL
HvK3FjprJRut3aSTFOxAR1UMqT2cxQPCDQH7sogTguYnHLjQwvncVWmn1JO1t7xo
z+7L6AmbJnqAluItiGvwj+fb1IsEMoJZixZ/plEqgp46WlQ4sVADW5x82I700KJK
Sfz0bdfNma0U+tPgrxS4wn0RkzDuuOccX+iiZBA0EdHinCXMZs1RyxVdD7uAjhbT
Hps4F5NXFcfdrmtYK4OQsCYyVY9AnxcO7q7lWffHLHKch0erRkSYKRZfmMi/xcAa
1MEDArCIZjhlGFVqZH8Ebv6og8X1kub9Uh4sSJLdXVhzSPcRZkOsyjPVzLpDUyLf
KClP8yxuIvKm7IIrNhs/dRPsvGqKzVPDn5P/VdXNxfU7cUaqvXkm2Il6anAx1wwq
XAfXOl39Dr6jBHRMI52a0sfOMKIkW4IP4Wbz5c4bfIj5OjLGONp1AJz+NyB8awSP
OEw77PtISKzM2/92aTgSboP1lUaGRKHWHqgVqPDWtrdKIF4GhxzocV9WIST4+zIP
PsA6E3n/wjSW2BYUjtR9y/JKaSzcs6TdJ7RqFBHEfEoyNd9EQYO+UvrEAuwHqU+T
nxOOyQQSykJLV3lnmSjhqcujflIrwwPziCVoYri2wk61AYR44XXU2wJ6nPlzTOnY
xC0neF04lb8RxT1UbEDvLHtdBe6cU+R/H8utD4iwe9g=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nKEw7SdKA4lO0QLekPNL3ew15dz6arPWHelecy6ZIwh/kA589L6Lq20lssA2LKoI
5ioxh8Bz7AjIBfnfJj0xGQ7WL7ZM8xy8TCVvDux/fYdZO5S50gj/GxYS65S3964W
YB6zgWgNUhQjcrflI1hinyakU240mjPd1vVXvdezNWBFFlsjLLwVtRKueQMZVpce
UOjCS5/J7JCN9WOi6czPNjCWu3Mp//bvMGYrjSJOLSXT8JHgEusc1ZJdx7RMAarh
s7HQl1sCZEkt/mTlDtEI89olHZsusaKlK8iMGN4ygB1Z8uNVzRXzGDzGWb+7kue7
strQYaYb18tG662atRoO6Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 20368 )
`pragma protect data_block
4szEHw5sd4z/nsOs07eTzYHNDrSmGinvK11FrUkv4tqmDC3CEFSoNvq2L3AokFj3
RKB+o25t2Iq/VwytPDsWVL4Qj7nMJgL5K29reSBup1V0HqwuYi8ZOJ6tyZ4E2cuz
dJWdpeIPyF3WRcDScEaNQcchID6vZ+M+LimbyedFsPR5uyDXzDHhZQdnzpUrxLmx
uUqLqEBImLpw5mQfEcFZxHLgwv2VS/yujGX+9RYqLiD+ygvTJu3DmRB72kr3D0m2
cbbpOc7XIQL/4cS0YW/6WVOX+mIUXvF0GT9UZuubUGcMmn2oJYYfvSGoNudpDVub
EUIdRIVBFymCvNJL0JMD7dvutBCEu7V+pszIpiLddFSFOT9+6qZv4WbGtqomUK9L
tt5tyY0srrZmCIbx5zSW7ldPzLJzYEAwfxF0XI+j/rEXeMwZIWknlF5ExsTX5lId
e0gEF8DZtP34kjxa3FAQ3rasPak/W0Lj0ObUfhWOQOExoRMYUAHkt3tXLo+a4Bs8
LfGPgGukhXtYE2gd6XgQudzoDqqXggW+GdwjTdkz9Uvnq7z17yuN4wHzZCRQmkII
qo4mvIvhwHIv5uX6+VCqDw6vIKg7iyxLzOfDte7nSjEHnpsHFxQUfq6g6vFi+v4w
9HgIRnuozjzu29SKJTUhHesWnA4/7fbyB/9BHuWtrS3ecrzcWRqK23xSyiDYPIPe
l8RH3vnTqtmulLxr3BJmuG7DxjA+PZOT8GfF4srNP2WNsbkELdY8fbjYOmonp1Tx
EOzUzolEY3thtDV6LE02jdKPGWe1OnjXHuzLrnsJdfCTt68twalKs+o+w3eImZaQ
v5cM5DubpI96AzWsgQZ1KyYJ5PaRLTb93oItbirMRS68eieaBcTmCjECR22SiL39
ps18QQV3KtJtUbCYtUHAdTNEAxIGBggxnvleIq29L6po5csm0YestaNnjD/k55NO
xzRns/jp2tExNzaSsSF5ZIdGWStu6O97u+GvNAAtlInhShWXV3VOKG2vPftJR40P
mrCd4ui9L8+gwRftLpFjUXWBqxY/4FUOXfHo3ww0Eq5Meu0418BLFETwR+PLJzuV
D/x054UCiX33uUznW1OooieglmWbdhD85fQ/lfQ2Bj+au6BvxFGbIa6L1uavgFt4
67AfnkSRPlt6VPqSEq5hwXM5gifWaufY1NnPxKzJKnktZr/f+MZHIwStnkNqUbCc
DZ12q4h0yjC8RO9nymBygxg/X+u0yaKJ2u3qxojCh3t1Nu7PHo4rWEZQ/Ku6TgLC
XaeePTYC5kiaapB4WTW6bLn1s3p+NoREpE5MEgSpD4xKl5fB7BKpdil71dhYF5Wx
XNG1Rhs/JuN2wJW3IpVKLyg4jkgvGZiUghhiBPO3xXxcexR4qPbvnfWDe3xwIrRp
NV1vu67AG79RYu3IyYGQ1XQrxa1bn2z4luM8UOOVKLhzLOrWo5fLOpOZb+ziFplY
uTouiJVNk5j+Mo0y6YjJJ5OFM48AoWWgocHYQ+nLYl6pVxbDJjFEMxg97pGgXDNJ
1hqBxFq+vUVew+r9h6pCLPCHk8kWbRr5GZCKEioiPw9XfDc6YGhiWvjiZrISj3/e
Rlt/vQSJVanB7nW9IIbsV5L0uGv35p+kPnW7MNdALR/+GOYhxNuoRYL1Dot1Ox4N
hLYj6+wUBHb6luRvKAKuLTB0RGTsrLvEJ8fVIzpPNf0rhhTumpbFQ+dWUrZ9Fnw9
QHkhud1+iwG9qiIi9rNe7fLkkcC1y2kfm/YrxJgTOFIkz84QOk9wsXmYzk0GCUWX
WNKah0oZNiWCmr/DuIeClLQT+GqK+KvR4PIrCzPU1YqFOs2GfZtSkTRcTP3Aqorv
nHjBMUuoew6znbayd5sUtmPQBoRotGoQhee14T177OI0C7xcrualHnkqaKt6Kpi7
pTGaxmmP9XBtdvHMzsT1wCjEqISDEjFSaRrXV1Y5eaEplA6K6Ij1+VVoxAGdzG+Q
XhKIctXPVrE4Eel86YaYcb5DTV4MJi9L1aonJXbSLdqp/I0QaATwjdpDoc1tzia3
tnl+VdVCEMq+gmRP3RGjjgmlwzHVZ8+sMhvPTAFtXiQwtQ2neLdzDAFvYJEri/mK
EIYcedm1sYGVW4H5l/X0aWLF8fe1ti6cEjQBaFJYMCGmQ2XiY83S69+Umfy+SpYr
3+1VeMSfF8zE26X1v+n0q7Uj4aplxmtph3SWwv2j4GKiYeUmX9DNnd5Qvd/Mxr4J
Z0tZfWpSfZS/ERE/G7RXJKmVT5q9ZVUmMnW43b/4yZwkxvlDvGy2gq6cikzk5B/b
9CH6/dbWmztVQVWOUhkBN+k95pTmqyvzo+i9h7p6bM/x0Xj6wRd/aD8XcMFQatzL
LFUD/rMU95BQwaX7WogucHeJsIr3Y014oKxi5ZnX+TJ4l0LbwLxuRGBO44etpec4
jlS7S2r26hx9D266qbluDJLna8ipcOgbuUFrl/RfQFPpoK55t99rvmdAVJn9Ue+Y
Z/2/0IvOSi4a6pZRMy7ygYpp6G6FPmdy1D81oBZqKlH04bW5cAZYkhznehZHWh8W
FRhHBf7bJRIHCHOJeZdALH+gx50fathCzvHldTNh69lDNaP+qKt0+uBlbBJ2JZbd
j9PpHAEWQ/f3U7FQnMT+kju0nE79w2gY1ndtt84VFz2KLj4nRQi2435TI16bGLu8
rnS6scsAqig+I2A+nd3jdtZMGtzmCBFxQuYWdkvpVnT+Xt1GqM3AnBBB+FFJ4ZLu
z/GWP4BCLv0KxBK9Ho/F1Jlt2pmNaRZNq4UE9dPVVM//e8Jdq10I3Mt9fo84e8A1
ZaTBFicR0INDldY3dGqPS6F4ctCQPACQd7LnZM/jbD75IWsBjhikWhTusi6A9BuZ
dVxWIPHKWOhoF2m+ZVlIEv1Nm+ZATV92ZP9HwECiosRFVyZcw5xYSfhI0PUg3XiA
vNSK/zhyFSYGdv9iHYrPofli/SaAPJHGJ7go1oA+M30pelDwGNo4pTWa4amGaStM
nJ567a1CDq9hGl7LSZSGUojwhJqT3i4ETfKhETE4IYcKOmtuGzothCVJcDBTAAI9
oHfDOeNfqmZ4Ql814P0IyXmYGouruCoV6gHjJ991w9mjGmPP3Y8TQdK5oN6qfHC8
39uOM5Hw4CdorKTBxNMduRMJym4KXgPuF6xtwXWAgSQuEX/hdJtFGT5mldT49HZS
t4X2pAY0gTxKNy6iILwXIoKx4FhRXZJBT5J+IQlRVWx2QmUXdoXhzMctY2KVhPMx
nLwAkLaSjoes8ZdpJ8kqgvX3JnfI/7hr8WlErKZMKOND3gdRgXvbqYZpq/dARYg6
dO7KD0RClaLzWrJo4VzVbncTIxQXfordDGgjmDsYzlaM5tiMGCwcmUmJd8pacshD
vD5TCQdS7GDVnE9/ZlTWNMmp5hKeC2VoHaWwU2vtl8W5yKbSMxXSazesLFviv/Y4
DavsHSaNAGrutV/uk1SNpR6Vg0p6sDcXGA8gGbekVLgsZz8mkisE8iRFKzV4O/Jw
GLSmHLiCuONGp/YDdAP+vq6Ssdzu5VxbGxvhNlLvRQJUJZBIhBHyfYLixZ681HBv
kBKKmwk1U4HGWeYDmeE0ik6l2cP71GO55CmzHd4lU/VDCVSySM34GDSs+EtzFOww
8PZ7sPzenXXigb9rK6nBxUiqFrn2ypOvCHuNGqIYlY5VWPxLglPbljAoOLo+TKUJ
2ULSUiAOovs0a16eiaM4Nz22tzGiCli3hErxkv8Q+fILVWD9C62rvATChwCrTosv
VVluH1NEXM41t7PqMUoZck1nas/9cNAagjLEx8QaJauyGXETmYwiEi4QQlDGLeF6
ax35f8YHsjItOQaYMaqqv+Hf/1+LLrZ1OHOy25VF7+jvwWpvh6nWQXT+EuRSv88D
uQtpUeZZqEffua+Fmk0C9d30N9UktDRECgz3MnmSjNJfEq5s8KhvWyYLON5zfzKw
wMnfRmvtAbJQTrQSI9vAYJd7XZcAgYxen6xVZMqGt4bc1XVLM4+bTvvEylH2IjKA
lxTgK+qTjGGlyIajytKg+Ir7Y3QNbZs3k3FRHYVHAaIlNp7ugwVOOcHUx+MlIjTb
d3QzKwdXx1n0AODixflUlXK30Swwx7Wdt+NpL+gkkCbdISXmZxyWdE+MD0Js3sWl
wUdu4kIsF47s8p1ndCZqqnZX+XQwVwrEdDzAL2Z0nOi5FwLIC8dHVR1P1TWN0k0r
uENJSVsOS5OiXyxCzWgZpbHeh8pBpHxIZ7rPA0f7sEbS5kwGyhb/hXtL6cJvU9Tn
+8YOiHybWyUOK+6OLThrmAxGtvalk9voumNnkI/9SzxRzBM/a+xKe74fufY/QcL/
RzgHZmeRuTFwvToa7RrQVnkyzQJo+lEQbUdgTvRi06mndhuoRdFbFPpDq0vO/i7P
PyA5TveEyvL/woNlqL80nd9Bn2sgqm4HjF71SRfRnVK8lCNlHnlBJwaQnuGJe6uk
yTpldPCRFw8T+B/Hje6VvJHsjjUT6xsdynT6TgJ83u+wvlDbp/d0vaMeEqDffCsr
OSM7QFZ4hgGv3GhgC5qHGPESxx94laW17uyic0tAoej35+6VXBX889J/E6mkm2i0
zYrFyxBZptcROwdLEE2tGRG4oHMAz/WwQgQzw7NEyyTR0EZP0vop+R8WAcCpG26N
a/xJ4HnDuk3gZgv5ZslwfdICJCiD+hufDg4gbT5dly4WZsYKIBEllQkyplUtA16X
pejTkk530NOZJjEHzzdMrc2do0gheR1jcG/gB55MK8eapGlLjJE86ig5Tk4bu7Ea
ACaYQKsn0fxu8B5nJWY/ajhRdDI5++C7kycCRYf49fLchZNj3qyZtkHeR7Sikzgz
7PYt5XozI54sN22If9RGVTK26CF8YfwJ98IZuro3JivjUVkQSxV0I6ucQqNTU+BN
+f65zA2gwFsbBw7fhA6lezOtzTDv8jmGrjMY1mqzJVby1jSTKwxLRkbo9Y08VkfB
NXtD91xSlUovYD504B6E2EKF/AydvHFWhTIO0wTFixercf+yjz2Zbi1RTm2k5s5u
raUkrnh5hl7bbqExK+HCDYLZ+U/HX7uRHg/j+hXPKIlQ6CCwAjFWAt9g/MYZcwtM
Ij8JRoudcFnudZc+zl5aFJfBKBu0fNhmDortWFLtfKxs7/1y+p3Ax/E022KDGBmc
w7mCq1cedkubO4+dRxFABnYg9SFJVXB/ElvnNLSsGs6/3VGTlQVhpj4u60cbi5bd
/I004W2MOu7zx5jqaHQyPZSXAFmIMhN8uppqStuTebCM+uZyiWGgHDzpWZLNvQXY
kgw6pKxzVj6RQCkcOzw6E3Zg5XzUuDZPo+E06N1vmLxGf2hCt3fzHyUbRhGItLYt
yd8db+571kA0ZAqsz9mtayFycxIBSAMkAjGakZHHyaZlqjX5HbJ2lVGDjcPXumim
purGhp/tJtIdZI7GHg8FAPmMGrItr8qaaJd11MThzHHGwZ23N392YV6EsMpVBTb/
LVLX0paGa473wBJMqkGfg26Vtg2m6ExsRTepz/J4IUxv7oodDtVJUjdbPDYwx9m9
r7Dhu6hpjHl3TonGhHwskb6KufUuTtiCLFWZrQ5IgUfRbW9l59M9B21AFzYTbDie
ScJW8OSeD0j1hO7oJd2ibBYsc1tH2DNy8FB0fkR10AwhoRd/wNYx//Pe9nU9Brb3
kW/q4q0rIfxb27onvfXC5ei26eRcNOHLX2sO4u3eqwkO/mxPYgR4fOX2Z06hu79h
GD4RW9tfzUtIElhCApDriuhDBWZMcf7/st0bevwlmQUIQ/q2RYvwuL2dsmPI+Jcz
eFh/FlTr7CKykX6QAo9SSkJMLwPw6yTc5++Sw03AfS1RqE8XMujYFRxpdLj+yJJq
YR7GvHo3PGJn/9PDrQL0QEC1Gbx7plEomTzz2pKPX7aUl7k9xviC3b4NzohqWCx5
pNb5nyWOulRZKYrYkdW+RhYnjNc+jhwml2dMFFFDeDITDIQujaJjwnPWg9ls/MTg
tlfAeW2dx98mKithjTyfe0fiNSZVpcHT0cT1eelYJnVJUJYR+5nuiSVVzbGX1IGK
+Lcn/8WJNIhDWmaZNjQrpMhF6A13s/j5ICvdgAWdO2o9EdNOsqGMEhsbkJyvKIdO
odkOXD5fbkzCuFN/f6h6Rqx6uaH2wNPOXGjZy0JZCAyUFLNuudc5euwsw19hh8Em
6pGZSY5BMFcGYiwUuhj8R7lz4HSQq3bArnZMz/w51icGzxKaOZtmqNlM3nJg0lkt
qO50Vv1F3un8JiZeXHBB4p3VRqNyXbIPzxYjNaLnURo2m6nYTdyXAP25nheA4F6R
GOXc5vvju5bWAvJ2sw6Mcs+YK/X0+Arc/zJlW/Wcqf5bHzOYFkktrvloVeZ+k085
AHwvEpsKRxFoihDhbirMSJwAYJBvA/d2BoS1Q3snfeQnKAbNM03xZa7H9lOzo5Ij
GSAkXoEKIePjMb81Uib4QxMAxLM2VoZba67QmFV3QHNHSP0/9Bp7w3XuYUjrefkr
e6qyxJyA02DmKYSr0tG8cwCHCH4+OPUhgUh5X6uZ967ZGN5b0D+fvkjgy59r9dJP
fO2RyPEmr1K9+xBK0sg/pZYN3nNU6TaeRh25T08aY2aydBa9svfi+b0TbudEZerC
KsjDmjILduX2KaT0Whd+fqi0V7ERTDC+r+9TZ4p7RDBOoNxyYFYfgZIlstXCIKOe
U0IyHlEYdSoHU0Rl2ISKHiryZ+En2i7lm9WR34uUjecX1j8rdg31wBJxbrCsOlVV
lxZx2jgWVfs107PkoP5fXTNPSC74YpG+qdPIMgm4eseBf667sOKDmghcVQWqzWRj
vM/bc3viNj1f1uVPXnFdNBMLFSyUuGW0slszh4r6GRkugdkELerWiqeqCosEgSO2
McttZV3PQQlyIbTZkH1Z040A6E8U3sUh3YlUZO15whADNri76XlhnCn2QN/9b5hL
I7pSij/yAG+SkSlG9OAPUeIhQ4A+ViLlFjZbhFC4HY1OpB6X/c3z6EgDNPorYKIF
cqE7JEwf5mjjXNSPlIjiToW1cKLXNYZx/d28khzNpraPWLy+Fqb31wGuVaUcP421
T20yp72ex/pRXS84WbIAvHaLw+DmWPNhOyfaJJi5SwGIbhyGTVaU1teP0FEyF9X4
6Pi7dybAIOeepVJyamSkSNESlCQkIF5CA9cTCmEBqW3q8xj/iR+63kjR5mGyf28m
X1p4yaIz8IoGT69x6c0fuKuFAr+uL5Iot3T9AFSgLyKsB2MAM7z70HNXoZS5Pp32
+kB+BFAKZW5BNth/uO2FwYoJyq5UGFSgeoyLhksMTR3NK2JRynGLOfhRV3kEec/r
jVvEPzvnliJkwos/ZqLyQqkXEa+WekilwzMM+MCbS6nJD7lfSjS4vb5Z6WimljmR
MZ8ezRhw2yGsR0m1MB0c2VHTOiPn4krBC94QunaoDdHOTz4LlL55YvX7M3c/b+4b
T4/HGEoBffsdlowIK2uHXNeiKefXtH5epxDAUXcZY/iN/NK4+7NYB3TPk4+7QRQI
w/MaM6MnEW0lhIHJKseFUASraYU8eD703TmCw8RWGaiANGM+lCDN7ewvv0fQjcZ5
ub1uPXYqB4hJmLN/dq/KmqQTe+v6SHIGmRcxOZD59ASLqEnKMGOzLfBfr0L7xZA7
n6SSzvO87E8GjqyOsOcW8EPfRZaudBnv2uZRXkwsp/X99wU6zg/BaMBsCJktdbVf
nN16fZqgzzPEHyG5ugVjp9yXHqUD+QyNqlG/bU/DTXrFhwjSJf0jmoa5sZWpVHd8
QJodrcJZxpR0N3YQFdgZffZiwcM5BmhRoTzX1a/ZXt2/PpJxoxOyH8hXM/JeGX59
tYGNZ9isrdHFTxDnxJcB7Qu/d1aFxbDUo4NFI9HFzoCQ2G9XnFfgmUfS1O5uWvbF
AKwJUnFGwiFMbsKrMDw+Ub6O3twl/gaULkbbmnq7guXu7tBQMPK6LxjNxektPdK4
y3sMynOigpDbNLNmSjQMctdnax34GBr6S9hjLsFEmUl9CLi7LW+1CtSO2HQjpI1Q
l3/SzUrjYldXp0jodlDPtxbfyyP1qvFbvqYum0jbayA9OT0NoKcRpPT4oIYGSTxS
92VMmFdPERfq2Bypy96k93QmUWJby1H49d+okkZk3wi78trmbmld3IgBUw3fZH+3
3mhEUpb+DucuH6pC4kImE9V/cQHTWpR0CeZPdai1pbiR7wYi58u4HKrxu0Jr+T/S
4zjOkRq/svWUyg4pToHBmAV07c33Pkekk5bhdd9L4ti9tEgnD+W1wld/Gu/E+sFA
jU7IgIPDNmdSTjxcxnnd+SbicwlZ2Fx24/l2B8iwRSWsSVp2um+g89vktjTXmsr3
shVN4x9a+ov7g7PykrrIlYNB9Ufq+QNVDUl3/nyANIzsIP5FAk3lGqgNgvW8zhPJ
WzK4sGbH1J5PM/jkT1zeCr6oqEUXwf8gD7gCSnPhDj6mHXOtlVDz9IgMytMBIgrv
JG6tyPhmzoI8JCgofRcou1dZG55DmZsegOdDZtfmOd+oXBXbgr+A4Gr3LbfCPX9h
fuZYGTvfFRBaGDM9MtEZRSV7DbHVBjXn+Dq70EtP/7CQPigmYGKpNWv40GXAEr3x
a03FTK2LEX124/xd4mRt5lXdwGBLU5CgOph9eF7BTvXvJBDKZMn3VOJfCNFSuGlc
pTI01boRVJ4xeuB3qEhG29vzTp/SVCZPGpp+zbXZP2bSzOhKHf1lGD8Uos+t2K3e
9Sml7G8hhFAWWCWTsHSqHPbIvp9cXyT0QytnujECzICG+yu3acNczgsBGJoOFjk0
X9pTg8hk629FkRhfNG3UPmBGM/CGg99VfvCgJpM+aX0G595I0xavdsHPQs5245iF
3sPQl/T9wxZ79JymmNLjXLi8dBRgEemqg8SnQC68jPQ9rrXYU+dgLK+AzrkO9IHi
qwe0Zrt/zhXuyu3PolAYa1+5iJMW0oChrNoSDV3Kd+V5fQBYFiQ1XQhQ1eHBGryp
i4qKE2kNjv3MkKgibAoYrIGano7EFDlHNJDKZoCG2ew/luvHpaK5P6uv8aqwAn5w
ICqC1fIgwcJYh70M61kRymarytwhNTFpLgEX1zNGHJcAtAagENQP4QOf0SAHhjGi
WgsMCYpOZxK2ZpEXypy4LyMsGa5Cz/1HXGkzPLdtLyO3RRfRNRzFiLNi919kCyeJ
wVGB/GHEb7kFupCyLYc4NrO9QcrdBf5uk2+EFal23D4I5Pk2YbOGU3uicsTILij2
alnNpQknjUrzCyKObxFtUfLZTErFh/MYW8szGRynrJqIjnJSsTlG6vY7Yo5zExsj
dVEk/D2+5c0XFgPQCKs6cVUlIr4hOfx3EhBlU3buorlrsLuqeW991yhEAlU2Oryv
F9X+jCFURI+OUFcWdG6vWgfG6dVIto1u+US0HOBt7XYjjndEdkiw43/j0nk1LDeN
nyAei9xnETJCJ64lJfpxzMgfJMXUmpHkUdXT7FWqyW2flnGKZykb7cYeb2zfGiiX
1CGTYkKGIBaybUAFxTz43WRnQo6xqhYP8ACrJIcyGvWOUSP4p1GjFp2VXJV9mo4u
htodfsutHb0zzBM1OeNOpSkGq12qrGgpO4m0PW2iXirCkfJiCey1f6ds/9V6n78f
SXSZxaX8wtkPQK1duf9+3/3ESo6/H9bf0LYgCt0VLiVP2npRBCX/OK6k+b7JCVEg
01kXH4GJhBWJqGX6mUx0+C+xGx/Pm0SRDY+pM0wWn+Q+YYvuOga6i60jFjQzgCQr
ByaQ/vQ16euTw/JAjTsSUhi71V7AAPmNk9ySoxrexULzPwJBOEMVUpsk7xaQOjIG
7+SVPCIB4GRr7S7wBdwLWKsYrajwfE4s8cdmjUReLkRtBBflshwFdiQrCA8QQr4s
/AxXJ7m4ZUL7pYOGALxhNSGCt2YHQZ4B1tVTp20wh5jxhTGWHuI0XxxhB7EcLBAT
9tNP7vEMy/o1sJ283MvfJxh+nZ9apaA2A5qd28REH3ONp91th2eCJxErIK14esFB
Td0C5WqHeflu9e9Iojk0fLmAh8iNWN/zYW1frx65PnQGu5A+HEH8XxMXMFGpHKAc
8cl01qvgxzCuIcrPXFyVNRqsd1DHtcYQI03VrMqarHCHYSWqr2WO2cF+Jy4F4fLB
YEPn/3RM9K4hqtGqMGUydIK0ZcRypTEZ9hCG+9fVgrBT96Mc9G3Hi5Bl6Nqos88w
pL3kRSCAAJI/S5DQ8Ul/5q12i6JkoOOlM798CAUoQAiSZBUCrVZb0NfxLKO6lgLC
xacPZR4SCHzOj/VzqqqfHe/Xl0vfeLk1mArbxmzR0tlRjEwTbcGoOavBcCIUmSsF
wjWvPGb0PtG0CQLYhcED7KMmLIAFcePhifAvFL8k6MEW46zM279vA6TgLX6P2A+b
orXJxes4zrZVU6i5YelLKESMjD/ocgqFEQ5eEQrnjCJVOSE7JRFKKUJf6xBwMMWF
C4kB05EYm2+wNsoHUzOoyVQeorazjjsjSKYJKIBE33ymW3Hk1Vx2bvnbLOmSk7ni
KcByvmuY92yvJ3Le0wZEvVed9sx+JhbEou60dUikYz29JPI5wCXJJpIduK4SQ/kV
rZZjQYDIzEuzpzh3sOoacPb4/IaVa26Afro/7uQtbKrEJJKFpqMVAXaK5OCJ06wz
G5l0et27dz/SDTmK+i+SxjJtqrlHXJyikKfMYpzeqCTk1S0tWJBOIkruOJEqdx2h
VRa2FAGTBzwz6IT+FeHHD0Q4WzlNbSbvgGfB+Fw0z+oAh1kLAp0mQTMhmp2bZHF0
T11IVhY1FeIhNWOq3fyBxSNJs2gxn13wVbP7xhkeiJjb4LbxEdSz+4GYIvs5KsPo
aQ3emcuGPyyfBkNrJWAlXS8EEakFGIpSXp1ul0f0K8ImVNfEhRqw+N0n4TWEy2mm
Zte7XlBXHUg/NrGFssMhCZgUVi78a7qf41cxORM2momWRWpmgicXuMM/u/VloNkz
2Fcv8qSqg0oL/+VyFQgrJTGMqfQ1OZWIpw0urqPYjdgS/Ly+dVSYhyKihRPlYdF3
i1ZOJaGgfjxYI/23Yo/x0X/+uJXtERp8y6ttYwDvhI6JOQBl+050u9rCUR/hBOZO
dB00RrvrvhK4Oe02+NOOBqCYlkxmaB4YdnbjaBf/1ZRq/IUL3eB3pG06fupD8Vn3
0FZBcflhLviSIvQ1wMy/Dmwi3icJApMhnn2T0E8q/yqQMdBvtHuAFOmMWFN/xyG7
WrLMpdkIdbGNersJLuDJhg9z1uDgs9hTbZWl6c23akPtS8RgUOFMOBKGNyBb9Z2q
V3bpPdlBME7FBhVKA7qs1FhO0Gqvc5Fa2AlQMCG32DWRm4Skb7wssdTI4GZpSxKw
Ba5jmHw1Psrmm7WS/WJ64iQFJ5izKg+G3qbHMu1TUT4EKF20ibu+Wn3O5MmHE1Mm
WGhA2SNCeidDQnycFhRq9oJZgVAoynmsqDWjvw65de0uyhmz2B9rYgt88kG6h0VF
hgiRKpDpAvSzDT0t73wp5ELImNPNimqLjKgyL/PN+zO0armoHbqXlOaC4IuaGlqN
RZ62L2vgLmfSSEXJv62JntJle58lnmBMJckoUfd44DSo31vD6CS4nPjZdl0tjsX4
z3fGp+0YQBnr5uQBNEgIv+XS2WC4jui8KyaZycopy/H0L6m7ktg2LzVgNt1Bf9kq
DiSVU0/PWwugsbxon8zjf4JUkIoZVixd5LUevC/+fZwUQgufF8BekimxlK7aqg+n
sxpYiB65TOkWSobYiC41+/+3Uiaj0HDS39LlACNXheNJ1H7yfd+FwUWB46jxsIaN
Kugmpd6laQaH60U2zPycaspOfA/4LNt7Z/06h9G5yPzG7E4nMc97pDbwjk/jeRDK
G1IhjUFX1dm0IjRhVyCd2Dx5s9Q/mMYsJIBT5pfdmvFtzGJxFyNM+5mffxooMTIs
x6mT0NFfajX6m3uy2R4L4G11iDjmYvOy8dyoqUYBwqs4QEw0KNJVuo/Nar27c0AW
s8k9CjaubYLSWMPcOFN8Kyy7d47JcXFR/NI8mkoqEJ0Pb6PN0c5p/KMDTz9AHzAo
vE9+DnoFTBrQdVrxmCh+r/wf0zllReFK6P1TEnp4BpZqpjnVJ37uHIALG4NfYxl8
w6IWuiJGkdEDAm9TfBISRcd5azWNaeoTiU6fLX9r9f04FZJqsBNMOrOWybaekhNN
PG9euWZmzy3bOEtH1qYbVvl+Mv30u8whT1IYsKww6E8Mn5x4ekjYvsV+KUc9B621
0658EDmJxVXVKjci3oT8qAwUlfRPLmV0aBx1J5lPEu8jdcmkMBiekzbC0RXWMZoG
NZaGFY5QaoxCszRPNo0CxzTgBLc6FPbyESlJDLkmj4yWyoTNcm7ixZGHkdpsf0D+
YX/POTNVqe8sKRQVnYpljb/rvO1GMh3oDkZg/sEo7BrcM+R9Hsff5aa3Xj6ysjYM
A5i+AwMyOOJsXrchA1r3kzGMtrIOhPj0ADfPbSCiFoidy41ByHkZsR+1jAwnqNpv
tGsuPKqPAXh4omSF1tS5OrylplC6e3Tpvhc3VR1y5cypyEByr8zt9j2Bb9PZiOZ4
BXPdN9H1WJPGfR/FmcZ6+XNJEsrhbORaiGsqWe2j5NBvzNyD+3r6fysaAkii1Wan
uu32JkpN2nnG7EoUaRoMFuWBpFwlILCIyecj51uV8FkkDQHBYfdok9JRIbSmdu0E
pUdcLDAamNwWbl7Sf2xkzqJj1snJX09LQh++aW1hUKU7IqDaiU7nLDzUPRiw2PHy
dkxgVWMstQyNX8F+Z9rLGc5MmNm3hNsTUGUxRxI+WxFWuvd7/wi8JVkXcpSR2eJ9
fdIeLXH2nzuiV0tecTV65il1hK9k3VQya9E2+DUpllGco8rMEOPoquXbJx9vxoIi
3I236tOQTNbFMgcBvXe0ZJwb9s6elFeVEtgiwQwVTueiMipvYGAq2JTwEU8l5gtt
49Q4V9zC96cBVfIH+jWFStUY4onnt30lY8Wdv2+b9WaJYV1ycCNH+7FL2s1tiCll
9PO850e5Fab69CayKvzTWAfZt+dpPycopyozJMguAX2XFL2w1RiAmJkJgdHdMWSg
U1pCGubJQu4XWdfzY83qdfU6U5hDwoYwzXAfDj7I4Nski7cQN68omWZmRZAFyVpX
BwiJiVOdg7ol8+gIoL+gtJW2zWZr775opsjN+AYZ84KWYvHVlOS/mwctghn45bGl
If4fA4kduf2OqLEYyxIToNhaeqJEbQXWQzbgYFuIyxWNQyDWmsV88FI3cFiYXSMA
SRuV9HgjlkDTgY7LnCzVNxur9efxXQFzVSrDUaJIm2RoUBoFDLzyF2x6mn8dru6L
Cc6+apd8+kq179Vi3fbNHN0d2kYDEQgQiJYakuPujOVMXwUEXDr8A+QNp83JNYcX
4xtD3KwDYqUYwz172RtC6ZrI8lqqo2NSve8mNFMZ28RsZ0LbR8eF6fHEU0t6hrZM
otiTEcJXZP3pmipzbzkspwsuMOgmbL9ZfQLIhpATFJuP2FhlKjxK53LtSwpcs21P
jWOqU9Jeoks1z5aXoc4broMcpEE6fJoBdPItmkDgB2yoRocgYmi35FH4dxO1f6c3
r0ah2rkphBVB+zFRru2AF26OiIANvquvFIcB7L0ClFzj1V66r/0CskabzdcmrYgs
6JhD5aIKx6r8OUHc0IgsZPJkitRn8HL/kg/a4mAUZo/OBVfmlkDXNDQLcuvmUieU
ykr7esSLIJ/x1LNa1xmUiWB1BcYYmddYUb93uKuNlbtikgviagym4XXrLfmFGW9e
46SYOls12Cmn2XeV6R2IIdgoWg4j8cho9fbQGTG1vnE6VxJLCpTm7rApXmITb9xR
jiI5zYpyALUFl/WPDCFFl7RA23/4Oamkr13WSebJ/vOkFldcLH+wC705wH7eFYFn
b0vWGu6XfUKwlNZditcLau5untdjcxF/dBQ9v3pRXpo1A7YDamyTeeta+KDU2V86
AS83MOSEvnrdqmMw3mieQ4MXG59St7kHYQzukI8/NiGbEZEN9iNDEB+ba+bFr2mh
5OXfNykF9sg+SmGhUlSqLkUuSHJkLQnosVVh4C8XpDpJ5qLnufmrz93bik0gFWuq
BQkBgy4wSpKGIEHzv2NkxvxpTlpvzSU1RsevRJvc/0XQZ2sZqCL+CQ0Uc+Fy9yZ3
sZFFK7vcgRPt9KvblVW5MIiDZpwpuf4yTNMeWzfRD5Jp37FTW+VfBs/KiVEkB+5H
U5VTbsWSRGHehZY2jDZRTPhOiPYNWHRSkJ78KXBsoGht6tUpvVSw+kHAqXUHOEyO
kgC354LIKQ3WlnKD18aOXHgZviNsq3uKE9rKoou/Ry0RGQR2Tbz9yEfqVH4ej9lb
eWqU2QvlZl2DtkWFzuVe8/G5pRXb10tze5exynOzR8tekKutpdHXrdgyyRCtw2ST
lLsnVy/Fj02tjDpHh4j8AGxXSMzgIunpoPtTy2acBbV6bXR7xyRluRQFrks09lrB
Tzb4NbELGFTr8fPnyRMHGTwBnbRC1ts6sKrmKAE2vbgO2cBai+uCDBUNHZIlg7XG
HRK2JyX6QdAlD1UaP5eYFk0FRFksygNTsN4YZTYxaHwO4WIJ1FAegKQoqvpYDlL8
Kml1r6PJcMEltFPhVmcKFH1op8KK+99LckE75VSWTvmAvSZF6HnYyaWsiC61zRYs
f1KTnAns1gdAT8ihczvMh6mroFeF2RpPHJJB5VLEAuHinYEXnGlJO1u3/5ySt/+4
CiAUid0BpHV7SjiURPi8zhXP4CBFGhHRaRj1DHJvGN0V1rkR3b8ubxLknLEPzdow
zfz5JQ3heLuHub1MahyMt1THsDUorYYXubKqEbYxtsq0uV+KWVKXyoSQWNCgQuCR
27PRewbTgFScn+sCeA3wJp/Jjeh9gnvA6S2rPe6HCAVjgSHBkZD7G/2Fon9gca9p
E5zC+b0VeqeigYBt3IZWHWO9Fii4LFPv/B0JMIqZ6SLC/Y9lMSnPuMy+FiwVrn49
MpTCPLtFaReAVLkNPidvdwknZEPaA31uMSxNs6PVhm9Xw+zpIlvDt/M/iDx0xYo6
9w5izIaV2CkYxgVK/zwDH6EOIiyVD4Wvs2JEk5MXljvMsxsGXpGqHWlDsbRQReX0
pb9fwIeo+7bwjoMOMhZUEadtRD8p0jegUu17vIM9uYyFuV7CsXBKvFVbU8LPtWmI
2VxOheODY8L+4Fa09qRoBT0l2xFomiej63Y1FTYsZukyZz2VmTnwz4Fy3TVzOAvL
X81+bLMTIPpuBl9bh4C4nuTf7orHx5CFCEwy9X8Hg7v8/0L2FIIx9hEZUqdhVEVJ
T3iFcZU7P6ECyUkd5MuC4WjxBki0ZWJw83AcK3b7TzCZmwQlATJtABWXiuh0knfY
Jr50F/dTBThZbRi5ewSZ4Ss9FuoNA/dwCwbIEPHmloFe+t5EEWi6BbMDC1osnRAv
8z7ugEEVKrX71XUrMeokYSpdIZB8m41P/f8JXpa1mOkvvaDiucp3Sa71CMeru/Gr
ZXuPsCadU0xcBtpWFfT/ZFXRcJg9X4isl6QY92VCneN0MPNL6DApfuDomzhGHUtz
IyImZXHYlpY4sAcw0iXd2rPNLINGDTF50fI/3ItvEJo17/IL3pN3BeZGsMtGZAET
GPGhmMSfFFKJNEJ6OLSzapmIlJLe3DuFKeqy6zOC9hWTGxTQQtF0clGNYxF+xeiG
c29r2jaimJ6/g8mTIaoOStiRWZqMh2SJ6WPQeVNxTtHks6ffUKqkQ5Uf79Plzl+a
V0DEGzTb7NyAx1ipeiCHia+GNMZZssORtbXyQIjiTqBt8YgAORkxp7AYbhMuAmZZ
WNPjgrJTfCXCNytLOlDjgBK5udUUr0GSgZ9NylHuN+utjpuD1VQy/WomIMFYORIB
Bbg0yWkAik4qCcp95MT0UbptawhG5fasKRaHbhPeLyQZOkOpuaS8vERZLebVwrjH
pvnFwyXCQuPoRO+c2q2ENky566GolBZ7Q+Bq5yyHjaEQPySABrr1PBfw/dVpbhhW
LxBI6cLkFgR/DJKisvhTkTKBkMb+IZs8SyiAnnwSR8jw84zpGzYnbak29Yf2DgNv
uDQBp5I5elGmxhC+uS5832rGPL/eBczl8mL+I3EFI7y4r8U/Trab/Jat2OMtci0B
QQX2MKaW5rVy4hwmo5SM4I3OSOmI6CXjeDN0M6sKI0tTDUcOJICho5uekbiD/YBz
HqKyLIWnpmCjDNuzAYdA5W7aVkIdYMCcVUQoyzLpLaeVxWqmUQQOcgy3SjkagtS5
gqleQsYe6JGYgHScacNbq72D+nimNmK3iwz+VOvo5aXXdVpmu4J8UDh1ZmLW6QsU
X5cF+QWYnAHHMUZnHWWGBXmsenGkbCB8v/bE53fYuhYq/H5V8+JxxVZ3Rjf0++X5
IOwTJqxbqRGUuty2rFoUJrWH5b+3HV/WFrvWTEGKSD3mOmfgAOclgqtER+QGoXQd
TkEyGqbrZthdMiPJJb4J14JLJE2zzVaXRKTYu3zLZ57DRliGAf8ROG2U8zx/O4ds
FwIO+CCP9u1KDjZHyGtn2vc+OgZ/LiZhPt4G5wRH4ctyn/0GwyOHpZNQl7+EIoWh
XbLUk9/Il2OUAdsaJblR2nVRcUXpfMlLfbhsgynHfOGu74SZBR0Y7/fRkZCagUCb
q2CnI9Kh9u6Ctux62nbqJsHR08KIApvjYlKxo556KQD2tUY/N6nyLjA5Xdpti+95
VcBK/CzKTxxYyp3pVVNDA0BT/1R5/Qm6hzBXmrjU3ytZxWFDbJAvMZeVrGOS3Ai5
hVtTv2I17fOGnIBKSUIf54FuqiM0n+lv9GXMyuVBBXi0miseyEmeL1mZ6bni7y5I
/LNZ69nFNdjJLGW+CVOkc8g6ffccpwzGMHM8E140YQ/Z5CCi/jixrHSE3SkHzPLL
lE9SZyPiY8GUm3CIO9PnMhfqJAoxTXNS1HrCVaolxeGA5akeCYng3P+nZODEsGFX
WHEFC+j8P0odTRF6MwP3SCcn+o6955snP6ESGCPhkNM1MpKN3t0BM+tXUAw0UvIW
TL1YTjR2bshrDrWiBuWoOuAQ8vY4GzhtorbY213ocgax1lYIRRGyaYGikDljc8G3
IINIrvbTmRG16gDj/hz8em2y+Sl0NJ6sDKs1LS89eOY7EtDek6FpPvbpKnnGigwb
6dIX052P5huD+TmxyITduuS2e5CVKsIpCmetrziZLLrG9emqH+xGcxMQtPsQEoVD
5JwzHjTpi7i6asfqJMWXrUOfzMnzkdXthLr/w4+d5DEDVHKqWKgrSgVsj3+3aiMj
uzY2IJtaBPrd2Lnpz3elsZM/jK0Ime9bmbML47jj1bL724g0yd5oupOAyy0oVtwo
0oHnjrBBxNTlcIiRcqKwtY5rBpVSDU6WbA2PvM1epcMAvbub4haLtPW9TwDuAq8p
h3foQwGj0+7kRZmQ6YFlGF9gVajW0P4oqAiG2PTJ805tIfMrFNcIMIJTJaJTtJz8
PeHHlJF0fiR3ovPNRaRSGGWdvNJ3UbMN6jF7Pd1j1UiE/KED1KVTSQ6dS2Ox3F6T
DI5Ty/y2jvKvik8jFDqHBNvzgXsO/KOQjWx9L6oC8rQl0TcwWGm1Sm66wSMEN5zi
ANf244X510TBE8m445AlISDbvCoNTq09/LOPFdKC1qKmb3W54xzEeGlEiMYj4uMF
OE/8qRm01KguynF/1UOBgBDBR7G2EkgZyuLdA9eBkoFtD0AlxGpeYAGNzaowWqbz
4A79CahMvcyQLPrN4UGDDMqJYh1NIXYYb5c3SEh8xvCGVnaodXsVEYdYyBFKZChp
ak/aq3F72zvzzpt1+h5ccF7Qmpkdot/MPtCkJvEA9wTykXkC1MT7ck8rcTGctGTi
pL1UCpARUp8E3T9i7+DWOb4S7UDD0siy3oposQPu0wdrlOj9Ynd2b1Izh8DOiY03
nAFYI/h8TiL9ScLp4Rb6onYsBlkudpkEsQM5BhqrJVo6UpiqxcQrIRiMzy0efNNn
hCQnXZbPmJViYCAt1lK3vfIRh+qmBaCreFlihUeWgTu3HkudaLwHh3aaxqw8YbiO
vsLWeSUXV3YW5j+ZNHAHDarVL/hxzDADrkfff8WHSB9fPyx9n29gRx7ig4lLaGAP
Ev+anx2A2SGVsXCXfmXLzqYJ2F0BvlygwDgxCNOBeCKbmn4/JW+7+6h9NaucGvHV
nTIq3U2V3hlFgE3DagDv6/XH/2HN81eYxrgwqZ9PEWTMK0nbcK5gDzM2VRiwSRNQ
ww3vvBoN3Vwo6p6gOQeFAd5eR+bBctIQn5XaocuguXLnUcO5D+utFGAeEe2+ZM87
wLeDIGGh5dBliBkzVs5ovVnf45YyOl3QJk7J2w6BzrlzqGfxt9klnQ44yZK6ZAiM
u0ELpA8NGMZYnZXrnJMseFOs5lmLDh3ZQnJlklBDSz0BdS23KOwdGjmfJowZ8h5e
KXuLWWSCpudiwegk1SJUk72vwLWuZmoY2pKZnuv537q6bPzYJBJ0sl8n52Ma/EZM
Fddxg5Zf9oyMwaW8hYXPSqhc0WnZBgVRiexwGr6Uxb2Rh2XZzHnEeL9tAfEW8Cua
qGPP81uT8FagQzzahTUXLXa6DrLVcuinJrbC7Lv0mlZ7rPPByWOZQefEAGWwOJoF
wLIFSGbMB/UmLdaAVwYouVE4lnylUzB/otmKJ+QfQoiAOCJ86YvOg5LvrPVQpxLC
9s/y9i86nfn54neYIhcF+Omz+SYdeIjR5Rwx/0sYTlmYY4iFOdx5ollm+oKKDxPR
B6nKrLptNbJsEB+BpMOCYZJwMQRGYXHHT8X111dkhAUFbqDkWVlll7aZqqi0EMNy
Zu8vXN5OQ7fdSlMECLF6k8UGHt/lTYScHeVFwZW/9o6Em4UT3K70LWVpctn14and
h+vkXqVR5ICRKoykTxIXc63ENS0jKkNBh6e3a1R0hTs4qBRgKlLHQ7VAxRjz959j
T9AgGvCx/5ZEvleTOgwtj9lYOp5aGtxF+5Q7KKtt9SOuMJsujpvVf4yFbsE9qau/
Be9u2DT+xyhnBNQ0HBIQTC95I17wHdEeivhC4qdc3iwQMR1iIM5HIXEw0JgA6io0
2K7mcHOPdfMUqFNGQcji9KywxdPqeXGqdQ1AUVr7KkPwmt6kDLrZLymOllCxyGtQ
Nxh+o+mmhaVRnZUmbsw/yp4fig/lTI/H7YjRQvcHxG/TOUiRyqt/9g5IzDDr7X2W
GsbGg+fII7lZkmePt07eXalevhgWIuLGw9yqn8JANyIYY+suI/5QJGvf8ume31S4
+47fluPgYTy+yaZ0/FgSdlrMUbvd+lBbhfVV3PPIgO6iE8Pv3B6wMxWUs6L3fjVl
DMzS+jT1NiZL2DiWR2wtHWNV0a9VFee7220QI721sATtqwWx9nROfSKyAR/CSgLx
+ivEP2Z83zd36lCr3KhaigEdm1Y3CFH0UE71irAQalqPxVE/or49Puj7cccLQqin
8Lf3Ya4or9dEMr9iJIRbW4LiaOkSfjNLnZ/3RAur3x/ZWIJZ/FP314fOW8/zWNW7
8lx5uZBSuK579fRnV4LzLH2DMS4PpdVDn08ZGSWgw6YvKUIB7ewFko3MQVp0Z4+G
WBBzMDlq8JrSXNHZkPlIeqRWQ0j8kLoJe6VXrd5v0+INpjtBQ9TXf+Nw3TNe1AhP
uCMuobVMBpg1JHfdWLT+cEvvIyhfQNSUXucbhn6Q1oOQLtipk7BXfsP3btO1s7qH
HqfV0IlBzst2P5udRGpuVPpOJTNL/Y+VAjCybJRt/LGl3SW1U9ARUoAKICNpbVxy
6rV9J0wKIh+QnwlEcyKAz8nrj1unNmcpdChgCidLF7Uw/YDn5NnPD7wG2ZjJL5Qu
vF3KKHVHQCBGNcatNRdY31OOT3j8ubMjr61knZODcWaV/fFF0yG2e+ZdLtu6nYe4
oWjPq0vEO2eZYI0+4SlSFh4MVFoqAUCSWm5gfdsWXYeEhQlWPoT821ipjZ7qJz4B
HOY9hqZvy8zd571B+SxZbqm9puMLs/+BmLlhmA3hWdEJEo0qmSimXpIjiZKGi6yH
tR2aSFMFPa0P2ZPEcv32+V1qhDV2Jn08cgXMaEJmCGrV8ma+78/lRTOt05rPY4gc
lXGKfJ+C2IWKT6i9HXU/FH2Bg714FTAT4Ch5N3oKpG6V14awtAX6ZZ82mYCfViEQ
pTIkXCVfNtXuZ6rAXCShuS+uocum8xtCDQrzCaUudwYYFclmj/qJRUkVn0RHBN7n
lBlp8WUYs7vVc9CdTWy6/KpkocTe9ZCvm3+IugjvrMlsVMH+eQkeqUXXFMnAq1Jk
mR/+aWj5xysftashH48oR1RvFCJiLLl3e1FJhnF7nFofU1rQJDmYSMv3xLZaxDmz
jnEM2G4DcwyGp46fpUQ/QBodMp0+d8aySIKyzv095Oxmc3fjMqdEmAYR069oucBk
Iz/e5UC53PD9wN2xrQKUy2s3+mDJB2WRGCuNWcrf2WTY+/h/BOHOjkO630o684/h
FL9CbGx4UyH6YNei8do3BAS6XDZg9ZMMxlOKrOelSUvTsT4xKO7Dcy3hgL/4xc3C
BPpjVdIaviiJTYKjo0ju6qdbsd74WJ3O05XM7ND5fcRszp49+drTX7h29UbFZrAy
MxD+A6xqHEVkaFQLSKN4X2OqamhK3BWlkQ7R1AHH+0giyzS7aRWKMRrlp+uwQv1S
qzUXRo4JVH+aA7RzG+yTx9vt7mScBfnZztmblaOywAb5CXO8lCxPbXh39WqNB6xI
sOag7NI+1NJvuXncmz2wYU+mAzE8f7xR2ESovbQS2CyDlddCB1RpyybhrkC1ikN5
1LFNf+HsqTJVILqN9seHkkdli5lPQ6tNxf7J+rdrdXT2ZpLVTHDgcjHZU7j1wagj
yeRI0k4p35DPQQ7gD1d84k0PfAo7vftRFHPwK82Bbd5ytliRj7fFE6ORef7/lPsJ
x9odwvIfdODG2ib47+mfL1kKHbxO679JWumGHy5CNw8Qog1L/Gmrj6WXpWk26Qza
0M0TvbwSHqoqJP/1yOi9t5ZtyshjwE6ohJF5HovX1K68K/PheuHxPIk+F02lTfa1
mYSltKNUAZ54u/aSsy+dbpfwFrl6Ofo6e7WpUuSTcjwNi3EAvCzUebD4YxXhEYHp
OPkyOj8amSrAhP1OS9ImE4JRxy/Xsp7Juq7tKjEoUmRhicFzvuyFqfMZ65kc3Cnb
LpY8bkP/I4zyZxX4N78aaK8BS2BPycbkGUt0JWe/gSV2dmWtYJYSOb1z5sbLk6l/
W868xU21X0SDrcxIn889UJWjCQXkqP6wVON4W7WzWBydKvAfs+tg80Gk1HVUU2Cn
pX6VDob1lN4Kf/djTOV5nCdckgFPHLV+c6FuULm0Jkqhkj2N3sbW9BAz/t3iHKvz
lQbEKxac/oFp7xoT0sikJM8FlvkZvR9DyAPNG5FAZ1r4mz9sgRG2IMFIn/RC506z
l1pDyCcMTeJdPR0r9UDSww4tAusPoSYJKYnu8Vko5XVoJwGN9htJEXS2qtP9staw
CxAP1d+vKsiEXF2gtAy6H1iWnlCQm8BQuwnG6MJo0XaOjhBaC2+HCMPpyXlwwvzG
gsdJE+PkgENXgXt+DcxvtJQ/m+hHNZzyfuqFhWCvoVMK5lbtBgTUqjJH182TSwNl
97rI4EhovCnXLZslVMoonCd7CyWVgWIY4cbvR/hDQnriwuM+g9LZHi17pPUCfMV+
ORR+6rEvfvjC9EZmu1+ar/aYN9P5mM5o8dsJBSENckI2kp15vC9h98qyk6IGSt+2
qEp5yHoCwzEsfhv2Ykstx6JGGCUC9qeRYgR06AtuBdjXfQ3RKZiffNsqDNcOg+UL
84KH4fjH9jlUVkOsdxGT/sw80aUS6J3WdMnpbJIW5xtuFLuROtmIaoulUpbyj7Oc
haPQtDGXsZK874XFr/N5+badCRX1MZDrvZTvr+fCeesB3BGPIyoyHc8+Ua2LAclJ
2MDyxMXmf6kfDC0M2fz0SC113nIRTE1tWTDTIdD12eBt3KmmbJFMNln4RM4N0X88
NZeM5cqoiMdWYLkZM2iK5dZrRZ6vCT8B1FJa5pe8CMNj1OUh6pZQ/BBrSDoYJdHM
szm/rK6uvWO1OCEHlccnr5FyymdMPOqjkVAvGBab5PWNtPaYD/BEY0qsrhbzjAm9
+1dVl5pw2yQKAkwXi08MCisxXTS1qGNWn+0A3gqkXyUuWKxvByH044VbzaHElQ0Y
pLIklQWzp/rRd8nojWwBRsMjR9uPx7ao1P4Hh5JDr+wehB34b0Jiz051/+z/d7hN
ItCd1GiThl3ppz8i+c+iIvHxwVK+WFBkb3m4VMrfrLAWIiRYNj6k53Nz2qInj7bQ
Sk+VkbJPGmsTrJGV+tXbRdm7JItTO3WqXErsvbvjNbTFiR7/JCLkqye6TaowgTMo
9mcTVs9xdm2isKz4eZUIj3gpqLspYOolZcR+mqkVkbpS6xiWd34oA3kV0GGah7sw
qblWnOQsJZsp1VAdjJp9cqulKLR6CTgLqPVgupgy5ASPFayry7cJA1/wvEeMUuan
PW4+y9urXgv6EcOyV4kFL1VFC/g7DdElxLk9S/Y+YIKjBWYf3y0yuDq8dM70xnMz
8fVAQouL61slg6I+Jy+foIZV0y9znl12UAin8xhZv4HXvmt9UliVajnQBP3fh7mm
t/75p8v5lafxCF+xwddVhQafGwmLxLZCI0zgodQmKCrTUEt1vZ7jV13b+sf4+T52
u78N+j6fTAFbCfE2aaFPtrPIPg8oJ8axmlk5WUu8amYdHKhpi6M4sJsKSzgz965/
ntfkiWPjhHCX9+M5SQEgyBa+ppjsZ7v85GFaSpHKCFtIowGXJ1WwHnt6fZ/6RaKl
w52n/IEqotzpAgrid5iAE5ZX+slVd2244kUexByupX5wBLU9l6gg08MPEQOOc3ox
yKXPHUkzJk9cCzereD8Dvm1wCdV+CzyN7e9mntUQxCJZzNGTJtSgLwqRsErHgEWI
NKi/QBbrVuLY36Y0LO/Jr5NunNoJTuUEyPgaZf2lqH/LXkn/INiNd7+lC5NVJgVw
6xpUI89c7yR3l+pCQc0uhZZ6DLJ4sew4WA4p0c3I/iRKvuUIMHXVlWu3mgTx/bOH
WvGt9EIDjFshqtdmPDXEQD68F3PIW4LEQQNmTTt9aLFSJ7sCpdy2IlKmTkkTcsLR
T9dRny7JO2TjTxvmU1NYkPeKTuymvxcZdsex1GMAcFSwQw3aJu5/JgwaqzYwQpDT
wwVo/OCy5W2FucWOm8r4VqKxulWxRx0d/FsOD4MN6FB65JzD6vEgwrEIOXPmoOA4
NXA7iXBz8XvQPzhv3I1JDJyh4k1HwsGDjPAU7NUwAjkSNshf8xZC/q7NJzyiI3EV
u34mGVRU5oFGI4WHh4JxNGK+tEXYNGxJI1x9XnbUmYK8N4prTL6c/JiSI3b8YZuu
jpOt18aIPbdVs/qv1irMcHGFE3GbvKdji7NDZqm+paN/2mcZ2Cc5b9I0uko7yX3j
D1YJxMHfYSbW4lCBJ090YgIaQQ+wwcyvDXoz66aZRPow+F3ngm2JmCLxO/G/2g/z
FBZ4/JiwgS60sxWDX6fzNN7Vkcp2fLxYXZBzJDKj+MvV60rHTgIMCSiuviaz6CGX
15pQ9YCEXaZ1SaZLWkStux5MA/PoysP5/L9kM6+P3rUtnQp8Wogv4WZfgH6I62+X
W/GepWHNn82jjQJBtAX/8sMXYIOdsrTAl0wMfl1jBnUcV+13LwE29vD7n6jNW7gK
aq8M33K2oxWf2PQIF7nizbH8bPcAk2KNllMRB6eHrgEvNG6t7kCyW6GMEVeCST66
71IGSGEMoDJUKYyESX7ayDZkglBw6JG9iha8pqbHtEziWv8gyKX93zsREvzWaBG+
JMMWUUqbiupYXaLKFVQCadVTwyhssLnCguuhGIih0J10DzW+Uy0zdu//7s2lDkHN
OSU6iYTkQrdrIxKpD/V193OBeTrO6Ms3HT6Xn/UGuFMlQWAT+spsTTj12u1uMRX2
lLaoHh8/Korx8HwHNJkLS7gbWZvv5KUjVJ85d63gRdTQZHr0Lpm9EfKSbFawsEtN
PtOWM++TA7vNqo1d45gjZ37m/njz8chApUsc5xf+0n8/oB//eHJ8oLH9kT8vLozZ
h12xs3NNLMBITJGLlB4flZNzF3TWxiIFUhB7XtCXTemgb52/9rSdDCOpOufgOEuw
7ydIJidBZ7eE25ERVlA6ialB4L/84HrZihv0v/4iPaWpIU25gIctp+Cmmtfh0c+X
PQdqx5i5ouMSLjd+0fY56jqLMU0FVmlZidPiYfeWGx4HNLwxm/KPPwwGcfQxb4As
4AjQKVTgLB95TXnxLwBMd9/gzuKvx5EI+RADBR1nKaxg4dR1VwxRDDMxGDzP8qR/
siWO2YoAN91oNojdHcwte6pUDWseb4rPmizwptXVLjbSRtRov5nr7wh9XQchGDMY
MVz3yNAQ98zvkVQKKbyhiBvmvy4AW0WzeIGw+r2ZndJHnSsYZ+KpxkM2kWUWwJbi
nojoQVGMbAVg4mMHx0Q8ipoZpTCfuwoRJtdhC8E0gyHfWgp46meQiTqtL2/UDCjF
vsTkARaSu9r4SlQ9IqDb4J1abUO3aOcvlEizak62vjsAAMA0U96LEK64fR8ux6ah
T32L+7kWCLkmNAgm7omU9VlmaVx0jJGsxAf7BOUWm3bwmm6XQu8S8GuiOQR3tOo/
Wo3T4pbD5GlmUaCT55Wj2UGBDDMl1ywQL+qWtHWgR0sr2FCTBDxc0Fc6P27Cj3gb
0bDoBIqrOdxB1hBM6TQKQyfPqPmiwOSJxklc2RA/uZ5rJdPwPQ4jyPjcqGDE8vbC
ChQGgGIS1IpNBOKtVA3yb2AR9W33BgzsR6PLEL147hBZIvT4yhBN6vWIv+pa/HST
l8rqEjATfLPlHwbOUFZfeHMR7kc8WwUbrUMVlk0/THzwJiXIlPGsrYAWFLU9z0bo
rqlpvnCCCvbPddE9qPH7OmzZR31d68jAnX9tYwBv73yMMHyX9P9xDpxQfDvDylQ5
EK4n9WyD4jldE7L0xTdEl66V8ykCQquXl0F1FsoXo7kGxMW/WHEaVxq+y0uiAbz/
lFwcE59EgVwicSUwTHhKwbTUo3iM8C67pTEUTzE6X9pJyqGhKkrb+HAC3aBtZfkV
rHZQco9xlmIbRwPwWnZTY08wXSTETFRZn9WxMucIdnJt5eguHvRV0Ksf4/htV8Oa
YSBQlfY0PvMW9UA2fBLclWCNslf0+PFp+Cg2RUAtD+HQV6nGOmpWhBmpb9zYi6Dz
EHzrQGUl43CIxvyAP6I8+ahqHTKPp28eEbew0LmJ6ii9dzshtloAGtU7HCnvZEFl
pXNXysxNvEnfLjxGTEmtbFVcqWKz68+aQORazZE8h1HU4kRsR8n+F+ezcS/ZorNE
ai76sTXU+tvBX6fkRUXOfk41aJE3ag4Ufb/346fuk1pBBHmhnIn3279ofBVeQqgA
aTbr1ItOh1Wy5iCP4iZt+DBQHWji1qvb4iySFpOUify8n174IsPwOHoA/AgbXlvU
i9/Uk2oVU4nmtlFBM3gi0nwQC42/nMkfwrDfLk5xkdPgnHSRlsFK8IHLd/8kbsxU
5RzvGCwNMblAR0lbig0HgE0fRLEz/gXw4wtH/kNiot2jyavdbkVO3lvQMz9H0V73
2p5z46Q3tClj12XXS6/XCvvjbD65hKSNPDMdoFuDo2Ev6E4Fdu9+pDy20W6tJAjY
yFZri3XvGpDdX9HNhGQ7kt/57NOS1fRtIxjHy02TUrSV8R5bY//3FItG9R3sIRn/
PWt9lrkelgeGwU7Qzu7BUT4xG3ipLzOemtmc5sy3sYHlLVwKk4j1tpmD8o/70XcK
1xgtzkpC2KUNxq6yA1x4/dmu8dQwxr6wPqAeGJmKocqVhiHgiurMH5ZWjLofphML
1qx5DSFcbYuN8gD7cp25Q710rr8RB+vi/pKFvXIf8NFTTzpXVKHdNGg3gwRirPLZ
tD1pQBs0HsKNhD5eTcNDg30z47Xy1X1XAt77a8RP1El1u2w+vNaaffSrm8kdwSzn
Yav09wAZP1Uh8vR9rZXjPZKIzOkRg/p/7M7bqxnLsVoI4CWdL98ohoshuVOrhUM4
qZwRm/C5hAcov8bRAAUklYVPwCENGIJWyQA7g/ul/OnDBtq6WzNqO2r68fpmFDRD
WhSSRRtuFRlFt6JHp7nl9ysk92h+Xe4UXcOqVedsV1OjdFvvZU/gstTf/jxgPk+9
3WSrEQE667BEUeEHD/+wLfA7ThOrSK6lPvdzlEVCJ7NOgh3KDXbyuaPGw8/7WEJM
AQ12lzZxL2nQjSwgLjPm5ZNjCy4GMCTdBerAIRpg4QmhoURXzuB4OQMi3T37jL0z
xWu03NtbChnbEgj4A1pay7c91M9SzeAgDR4vchbxV6b7U6vlLDT+OCPulQXavN92
42DMvbRVkGfUREp8PcDYI9Tdsu3HJs2KgEQvPc+DbRg3DYUrIwEXoEsTVSHfV939
x3+PylHGIPJbbz97B7WRCDkuzYvMcamD4k8+ET/H7OX2b2xXPHcJb9FBOeUwJ8qB
DxvXHJOvd8iJ3bivDeOrEj/YKCNVj4yEHnmI7fn0Pf8hqe4xoZTqDr6ILGMZw/0a
dM2DHdwzkQZvL296R4/ZYw7x6bDP012GOY+BI1zsNQor4lgVzRLNypi8otD1KZAd
NVO1zTT1kQnhtzlSlYbUKkO4EmmsKxk4wAfvMvolhyCMMT8d38jcnhySWWAIXt1j
I6NspcXrulQYxQ0CQz6pChynqRwgCta8vKepRFDMWCo+yVlm4hqXTWpJMR2QXy4w
oRw6FhYMyL2BNYP1Fk2I3uD8tscBjuOfoMrXEqNHEmTqRebLbwc4Ofzuv2F4O8Jy
bZOPBsaMJwl9Ale6pEFhTN5cSP/MdUyWgJmEe3eViqEWjf0wODhGDhvxELUeeAfc
c9OTlgNHp3xo/xEn9QitaFf7q7n17hw8slYq778zqi8m6qgKLVUx8soxM5iHz1wE
ZphtpOOHZfChwDM6DkDwTfEufBxN7u7Ut5SJsXPfutIgyc2pN78dKMY5h5O13qK5
6mCrbiGVPlkZ6YSfLLTiZQ==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
I04IvgHMJ/hrYLsqnpxwnaTWBRWi0z2Xadwa5Cj4ldas9oMUS5Y+NtT9zuGZ6lcf
fPAEsRMAM/dPPgVgyGUz/YSzI+GNQhkOAhRuWfaMvqpUSvRKfnpmXeUvUKB+yocY
XCjVJ95DEnUKPGGqlBZK4aEQVBGyoIUxBMWpumJRClTfTW6Tw1gI9i726hSJ54Ss
eF9urgyoddsv/FT6K4RSt69McIEuRfmxcWbq78an3zpKK3CBb33MtNc5H+PIIJ8j
RZZdmQVfnLa4X5SNIIAPrjrxZFTmEMHIHBLEtqj2aQAhOHNV/75+FZz0Jn6voOWQ
g4MhDlz21wspSoAOkpNnNw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2016 )
`pragma protect data_block
Xn90bldnwumU7DD4///VqyKhTS/cjqg9cPxWaJZygIgrlar09w6tr0UmTu0OLTXu
lQUokGVQ3qU3XLiidPv1rQmmhWN9Or68Lbk1gl+iL1B46WA7WIcqkqXWN5hJa8Wi
qPPf4s40ASNFfdVxVKSP51iMGYSszN+Jc6bgZTESKCj0aDfjF9MID/odUWjKcxoK
ywqk6iZtaLVQSLRNqFK5T3J0EbHfjSrTYla8YKxhxZepVj1xH+k2ACiR8A1lYz6J
vdIIh1el0F++L657NDIjA1EksU5CGWJU6s6tjNCiX8+rdD8Ek+sya+Bc34ti0eEG
1VoY0tWfAkeW73O2lM1S9b21l2danPACXl2gPTTWd2SKzQHr1sglJbe6L0tCwkPP
HrBElaIQ4sQyTY+MWDd7jlkbbuXlJu47Q7/hHzlqVtH9HYcf99pfagoEL5br7R3q
qqKDaI6S+KVLXakMaHdVHspmHvlPP7BdKIkIljwgD3546Z6S9M9peznFqbiyGrYa
LUYfXuPJYeebYuOmftltp+D46YhVK8EvMFHzrp3smm9G5RBQZ7wBOofsheOl+EvX
6wG914JpkFH0yBQEzNWm6hUj3JYfbuvgno9B4+bHX+2PduJSDPkNjO8WSBPlpGxZ
ooh1rnkhc8j3cOVmYYzewfzV0hOSNWm+YzD94g5auCo8ULSjYSYznL0iFNlZmxkn
wS3o1slS1v63UOs5qWwCNzbDOcaTFTuKfV1iUGgydNd0luaMobX7QeCD/0G5TroR
IL8t8Zsnaa4I2jXCGQs2o6tre/1I1yq/eJ+B3huc7Xn1/PDSJMsPhZLW1lZUuUAk
wAfUIDAGDrGRGRPUaKLqFGH+KL+Ck/3Td3mXp53HguGFoY+NXi7ncgz0l4i6/aMn
GLnCBix59XA4PlEntYC1Ma7+1H1BoyNqpj46KlXv/lgEVev0agFEIv1tX9Q4HDt6
XFS46fbgdCZo3w8KgvD0Lxj6Oas48CMgVXOqJf5J6miwMYBfmDrp8QCcT1BQIxx6
oByF2xGPx3kl2Yx6EEWF4PjGG/R4Wp/H5e+5W2ecPrKNcXcrMXsP5q9fQ1WnEbRk
RhbnBryREGHlcct13LEDpPwKhTl3a8zp5Gzx9zOuzzc1xEl4LMNdjh/Sb70BLKTk
2W3IsA76flIvieOez1nZGtl8opodiqMSv0If0w2puC81+J5UnQxkX8bg7FSjwTo+
GyJO8Opc5J6EyL6NbG9CMrkd0R09Fh3VZde6YHfdJ+mMgvdSvxbSbNxAeZslJ2kL
w0gKN0jKo1wOZIx9qkf18Ry6SewRc+X0HU3fyU9otEGhIDkAX/YKwdUDey4imfy6
XHeeQQcjQPIq6ms/uljDg2x1B4YJzdf5mE8Q3z4YrP1jch/nWkmexR6XStHH6SCb
HHBcbwN81gL51a3+q5ihgoCeEVVQOlGeG3uDZwm9+jzDcU9vVfyfh1DRXqV5tPLZ
2QkOjzv9qAKlv82Md+lsADyTIfHBynMSU2B6XFxu33rwd+gItP101O7hlZpRBXk5
PSNqn9zZX7V/8nIM1ixMn5CPql536+kqDIiMWizEGBMZEGjNWwUuSH8Y9q7gvha0
unnxoxtxYYydQnrPdAkPwdolJZEMaW1k3gHLTF/hWhRsVxKbbk2/0JUprSqHV6z+
o0AkWpCeFEt0E42UslY4dQa5nAhJG2tZ/Hbz+KLTgrKOE/heCkLLNZAqqpPARL9b
eFtZCDh6aAbvFBvrHX2fivqC2WJL+82mE/bxmTvRbEtje2jFsM1NkPWRqCDCWNgs
znetHAN0IhWPgHzOTcp1LsIvgHNrf3Or1WCCLMwVidV1C/pQTfM4pYwL35gVwErn
8r/9GMp9KkS2SLVD4+bEF8bnCJpVPp+TK04vLG3+Kw8H/dz85DgzILLVbJGsoxWT
QKPiyK/F2KlFgLeCrBWlShuQsFN4SC5daPucm5ozFDrsy7FZmAdYel34c+fkBYzz
eD3ANWn7jrp+9E+IsuJrtmYwobZuoPnjvZyEr6BXhigu/uGPpoBu6wlf8YJeaiHz
2j87Qc0vA7E1LwNHq3sfE9iA6VvoBQIa46p7IhvgC37d1XP9R5jCPp72nDSB7gPW
WzxbzrufvhG0iFKjq61b+P3jbj/jfMfFGYWGiPj5faN5CUWmDT6hPQkxEwS2HZoN
LaIdD4I1AZH/YPUAfLCt7AXTsuH/t87+UJOfBXF7OERTO5qFRRi/ZugQy5GiIuhZ
CLGjRLUDCESQYqzhRI/8bvScpznj4ngfVrRnOQrYzEoNhKKpiCgchlHaBiwUzgzr
9VzC0WXburNhpWMpyoKM1cL/n+LRFvgW5t5xoiRPcUdKm4jx+5qqLeFTQ/GT9Wkg
S6JGCV8Mw71P8+9CNx2Vi3BQ5bOT0/xU9tbcxzaCgMlqCGJXZvSE0h8Xe2rB2lzX
rsYivFb0NKSmp9LkMOC3yrbV+h+r1I0VNiz7wGVz1gE7RcEKxBEPv9Mdq24FJ7yg
Xp4vqteuoWQYZGVM2x2ytDcFEX5Ju0qNpz3xUC+ab4gP3nkWwC3aBU067pWcEU2X
vu8hPrAf1EeZ+0PHEl6DcSkPFuj83WrmMto/vAK+hsOfGyWzSeIIpIIQlG3DPwj1
4xkzImbbDP82aH3ctOHFKVAbXzZjeNbKgsk6gUMjs2sy+ats6+YpB9wQVB66/K4/
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NRgdNGog/ecEnCXuChhR/HqWHjTn4GwWr8i1MEIx34mhTKofdvEauppIa2Dv2qpR
2E1OdCLsJTkOUMEIfDuPjXz57VniyXiKPnLnGXAJOARSkVIp2q7ekN/PQOubGl9z
AzluE79CcrPlvV0RazCAJxdQ/f0HnhDqRQxWwBn6RMJSerHN54DuKqOJLOLYx/Os
O1q81swFK5m+xsdbh9ACBrAS6/K0zLbtAbqlu2DMDLqp2WnyCx1J/PatvCe7tsoY
BQa3Ahyn4nWmihISV31A/s2zaznHwfanLuF3ITqKO9nsWtg4uAq+i3kXKvE9rUFY
Pxf4HulZU61ZID0XutyZ5g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10976 )
`pragma protect data_block
zFwd5QikOmAU5tfPd410gw2Isc9FG2vd4SDOIPK1vWfY2TURObHCgAMD2Kt23Ra/
u3qjp8b4vbVb4S0TARqah6trqWeS9jR/nCYK/Wlavhu6r4BunPVsJddk7LCl203y
hlQJzK8X+ksuvO9+Pm6gq+2djox4PDs75zN6rC6K0gxSscFgQvR8nEpJrhWynL2B
dkgzJgoGAE/upgiCYurrLsV9GmDTIuu8j8nCRUNsueXZzOFKFxPriGdGvCuFGUKs
HnGEFUdvyo3I9IlvzrDd2MiW4RK0oAqAYqMyA2CRkGlVC6PdzKhyf5cz6i4DqpKH
y57iJEgnwQnZ9B5SrqvIMzmUWffQ0t6U8Fq1OYAGDu1Yz54Ne+FpM37QSDcMl4m8
t4CEN61SDP2kIByHGQ9BYSAU2C4MJv5lf34I92JNOVxERbUqPvm/oLD4+roxo6eQ
t8aAKSH+Vxd4ATJY/o90p6ILO/CiEdTN1vqlbBN2G4uq13Q17oSdXABzC5CEL+I+
lUNSDodRyqwtPGNPQi2Fe5vVdHC66OdUo2AHf/0BNVY4rE9qAlrSbRNz4+/Z7vYG
gwcgncAVMfDSyqWFpQImt56VNBYg854obnZ/7o8FRh3R/pmEzLEJN+CBzvO7Qn7I
WZ6Df9ZFlZhtdj5jhS+qoMki0pE7YK96X/89xiou6zqX2BXenUIewv+QWYFzGB4A
Ws3K5v3e0ikfw42rUw1VR4lgoUW0h/jDlABfbbCKfhUN2Z46cgY2HIAF0xUtr1up
rZ/zbLzav0pVfj2YjVPUZYM3+1JNk5TZcVNAyRZfb/9hoNeOMlg02orSiW9G9jMp
JDxqF0opX6mr25EFUJftwjJTIZDWDCCjN87KzaeQ9/QqLWGyJJCOgzyuw3h7k/x4
AnDcLXP9cjEaFyYRb4Ym1iwhugy/mVy3rnt7BzITE0cdkRhAPJP0tB2GhwDyjlel
b9IF2GKu44UBBfooyh/8OCpNdhzQzlk8ReeUaCVQ99+OT1gBs21lQ4+Fv6fQhl/2
+BFK2UMdMZ//vn2lLsvrBQlyCoIYCEPK3Ub9wyT94CJnxNQD4HSIRxCuLMK3llb4
i+GJAiagTdvNdQgD+wYONoAJnm0ajSPPTLr/SzEBQz0+OTt0WqGuIBtMy69QaE8C
x1u5oDXPXAYEQhjn5ekPDoQKrTdiHWeLO80sKEhAOIS5NWKXUlpi9uMXDxejOz9M
o9A+tmQawLk+Ait+iEvq5+jDI7OmNlKtpJjGfO0ddB8eJDq+SdcknF14lWQ9YzfF
lwJLwA8q4+W7GaYWCCYFRsVgokRe7TpxMLqRNiW200awoVDNWwxPJ3Tei6Pc+4z/
cT8ArSEVRm53GnDcyHhNEElNxHV2R7TFi5MMbZd40TdVUQCCeX8N4iAdOJv1IRHS
9DZHEOoT3tYgAToCw50MeOOnH12/J4w7XN4FjmbioicsxJQewZb4l7A0wo+fQb4L
5jIWYyBPrx3uh/N5yaTm2aVuvAchRNx5uSGF5+0/DhUGdVXGpQRGyTXef3U0rbJa
3teRSZh2QzuIf6QmlxuCZfhqxkxdlkRdRuB8NgsF2EqijTVGYrGGQZeH3rmKLU6e
Nt/TH59Jn4+YZVuYN0aAEkEOPOtIVgSvrgy/cfwKVj0LqDLix6FuvmY42f22yf+r
Y1DaEIGstQTaFqOgSL2sFVTkplzUebj772innA5I8OJatz/uWXlmq0KEBAKbGFf9
h7RVybUXLttpIPq9lL6Uyhy7vu52vTrKvtCyxekMKY+cBluFu3L7SZ7OwyV2HHDI
2SBxa+b59gBl/kVUOa00+5QYxOGAbvkOOlIHPNuKTRIajlVsb6dCBGKGNiUmXQOQ
BZFlOQD5PXafYgadcJyE3YDE7tQNtBh9KkKtM+l7bdjyGPd99tZg+x80AcxOkzKp
tSgMFE/VGAH9F9Vbd0UPFYEotAHjgROlzfUoLsFv3Z8+M9tz3Tlq3QwRhMf/mcU9
Ap77wKHsvYQWvHhjtgrMdWSBXNKi8bYhVfuyHCHZeWsm/SspS7ChM2I0efdG9hpN
dZwXoyg2RDCrZXc0+80sPL4t1HnyQgvwvsfOx7+nsxsnLFB79sTzLbQO5xRBKTx6
12KiEnqvDTUiuhKdn9TkvRAi53zX0VO8D1I2pdIWlHtyeW5Z6rDM+QjXF3XtjxHh
8kl4QdzKJVFCJIK4fftq8PJSnEekn7+oCXdQY71OlJr8Hg1pqbxaudLe/qJK3XmS
vzEWty0RIdfF2NPetvMoYZYBTw2WSeFW0RqymY9FKsL53S9DbIgQ9F2+C6v6hJ7o
fPGwMIvstri0Qv5wQJfQNIg5DwmT5gs5Vw+uCPrjH+xNVh2pnt7HXbCHdMjcsEHL
N50txFaGeuMVMGMm+vA2rUq3CtDSkxBDJZhZXCo+pzNZkqJPFOWERoGlwb0GW1Sb
Rk/ghzfhj/0BNcrDhBswgpaR3F8dN2a395uS1w2x2tCiA+ss70Be/hSiru0W8iH6
jLrbpsY+YGJ4zSOC7kXqhlcuLr2IzhhlnIKbMvIIPjShrmfiMaU1Tjpj1zGbOfMs
8ktwwwlM2TlZSWRGcJNZdUb6Od+ALH3YUSDV4PbsM6DnM+Aoz7JSARKro+jXeYwH
UpBY90cP4v3V7xdQOXdtvj6ipci+S7xCqxlvtWVUjk6O22gJlKlm/Vfu7FJzLxGG
dbSjSI2WMj3C+FDhtBhgybuy8f54REUVzRatbgxU29f3TVWwSQHHkgYgq95uVflf
Z2ScwfTub3CFJB5fekSxjpQvULMfy383ljs80ERQOwVFOCn5O6g3DgLhccARUD2t
5lyLtdLZMR5ZJrbXmxtossLg4Iz+bA0kuiM4/IJWB0OQRAMSr+UCBcY9dvCcIU5q
BQ8BTf287oQyK2P6Sh0Kwl1Lrs/ja3JcgN32b4wFnPjMLMAFZDEwq0rZwKz0UIxw
mqQ6pfZxtK9FErGuYIGbU/8/cm1nog92QCrF/FjGsPpw7yVjXBpiadMZzU1e4T0x
rQ6nhMpAB5jr8X1QfjJH062cWt2czRGDKKqYXWg2oSvirnzPAjDb18d4K7NkXhWC
xcZqGh00/YBqQxQt0VqPIzGUBz34y4FjJUmDCmHDcR/ZEG7rORP2a0ieFDEa5+Eh
ybbXl4j2Qw9UNKX5NJtwiZcCSr73xbmOOIjZOVDIbaZVuJenPPciYiIX3ycy9fKZ
wkdw6bqa8PrzlkBNAVBMqsXrNchmogkr2kfyH6/zshnty6z1DP3HsvyEgkyDNszt
b1wBs9TxhUj47TyIb9aKu6nQrsddG/Ot2bogkD0VuhaSlZFLIdfDWSSJasfmcW9k
I55/D7PpiTAVj+WDqeNzNswRcyiSFoFPk6x5a85ABN3U+4fM6kw4QoY23MPpKidz
oBl0Vb5YGWhX12vX1AyjNicz7MJIu5sF1Xf9guVbskLQH21k56WYxK6AA333cMPc
lmaZd0zcS91d3o2lGIhG0tx9A5kRmWUIcgmML4mNYojy4oOi/2sA6Px60O3UfPcf
Og6JHwvvoHpCGtZjIvfLVDqfAnFhO6CejS33WikAJq7Dd+OnSPTV79gMsU7sSzn1
hGK1r6gtoVcj2j7Z5yjHGBGLySUs4hLdm1PMVUVL03aENQZTwK0fEJhxGxq7Lm1o
vkTKjaK2fFmdVpTOXsjZFyhWpqit+Q51owo2xl0HDgVG1fjAURT73DdznYRMz7zs
u05DakBXK7VnHAgIF+SEt4dNzBtg6xHFck2LTpk4p1TPy78pDBe9cPAFTrN2rfiL
PRH2U/mTbeijcmtgoHGo6rBhXJLry9Az3r4Qu4LIVStNZnxN/kXLd6iggMyanxWI
0FtrSNkOiXhXDdwVJJQmM5Mv6PfNwuLnFqZL+/BkoMNfAe4/l3CAECBbi6wj3rJr
RAr3dv/K1XeA/JcLPg/0ECAJTDVjFtBa/2HNjCbr+i1CBTsQR4SoWqTTY9kFo1CF
8m0t7MIUSyKhkyzdqNjptDzCr3Ees/r1n0Ug5M9710Pf0AlDsuHkdCpVrX7UnZzb
K22yGYn9HCE3oIuAAQbbq4PHI0clS8VxsaZ3nZOnzfKNj7Jo3wl6HZZCdMMhmvEP
ZNYANKvVNWFSp6DPXM5e06Zf7O+P0Lkqj2x/9S1KIMoUfhihPZWVAvjowiD/dkAN
4SyPv7Gcg3H8KXeksiC1HEamP+T9sm8voTS/zF14HEClf+QfSajqCTuadZylqRL8
XygURNi4Mwx1rzWVWRqEyu7Sr38H78qlTmjhxjj2A3lzqqs7SLlZCcqZ6NS4FclB
NnYw2v4Ho5D1K82JVig+n8sVNoLdo5k+gJJdDif2fFoRXr6uknL9bbUic9k+X0iE
xRFGyzq5PuTmyNE+IY94hL9OlqY9dCXcfm4fEvK2qJos8kJ8PhwyCaD7ZpMvXhai
e4xEtoc3L4uhHFsqtYWQE1XFOOq8u7v38p1D7S9c/Gdnx6cSdJe7A38E05RKR/QX
YmyWocEVwdQAW84/F8sKvY8n1QHVq+/8jThGaB6t5mu2ryoTnyINqBzhR9ADhjkE
qLuxkUqAI8HBJYGh2ER+jsskvqcf4h6h9znnoZEg+RwvYlT8UkGCe57ig7M/dJ2P
AK9vowUK/ceejC11qUkQVGMrEt2BpsJD5xqmmjG1v8k/m1RIvAUcev+LlrXTCWEc
G1UGv4rFjYrs6IG9GzYKrzX4SQWRrO7/MszpJlXBGc0Usaa3Ap9DRxXM1YfGim9t
Gy7vCQQ63I1EtEvvdbbkiHaMS0YtJiRbBBLoGMbYGegKz2zcLAlWvqxcsM/9Uu5k
hmdTmUTZ5ob0gk9yvaF7sgqaITBk2unuPy/sm4THWeaLQMJRAgH2ZScNaRdZ/ao2
41grIiLdpuWeESZDJ+EGShjm18CpNOVtNow9FQ7TQVKJZNHkG2eTRXOEm3Ygd7sK
L8xIpx5E8cnSxz5GOXTViV1qJcOzcPUhZ4+G/xLSYepK1OZJoYJJ6oAZnakzP6Gs
2ws7gxNQzIb7KM7f4t1zo17jIf8byjQmj0G8JNh7uzk8zg1MzkLEqwg2QOuEbbq5
tbz8fjFdFka/zOcXRLqhkgiQJcMeidkqUQCuhOFoXNvNHqyfMZufR1j+UAf4rKNm
1VKYklBOryEZM1RO+Nw64SiUOyPAJM7aJn0UcplLIA8MVsjEaLe1uUKn0YXjf5Vu
o80UmIripJui5WHNK8eoUx5HwnycIYd7jjaA+8o4o4UdCD6A2ncjt0ANQaRTIUEC
9NEKgpGWf6Ig+dlXukQOgyucI35FnmxjqitdM/8Wu+D0laBlag1129y4GCPnzh2i
SOl7zuuKny7UCMOzRyZPAN8veK9jKP5M7ind/PEFelbiysw35aWe0H3tVThlseqX
kQ+my1tEsYRclKoGvdEQrUJFcs20jdHhyDv7xtzUI4NPImwD6xHV4t8YrlnPRuyp
wh77h4CNjfKzXCz/v+BdZWuZ3q7dgteMds6fRJLH9EfoNl9fYD1uR0OVu7QV0CRj
Yz3IxunPAprqUFa/1SVIaCXWePY7JKwPZPfjJWa2dz/P9u2LBYq0Z85g+iqfx/Ek
+JZt2B5tgS2EAZXMToU0zZfmVk8D5P8I62J4EDFn8K3r6S4GAuKi0U9ZhFkssBoV
ddmYFVpVyT7VF/V17Xc55eCUfSYEGcswMEuM761mSHI14LPlThBDOhJdn9nShoSq
hpvMPGe3bS8VVK1eXjZdFkZN6P9rPLQsfpfEjm+Lq3ZZ+k2f2sCVQ1DWcuZ56OhN
bH01ohm7D0emCeLaODDTeDaS5So+zInM9peaBTwz4GQh0jAALg6TyO0gCNB6MdEF
RgQOt+RpfpRKaAhsX/+al4RrtPlofgjkVvO7ye3pmp/m86TuNkztzb5o5OqfoTij
CZiqGbdZMNhagP2KnZNBRDI/RtC2m0JYBvekDWoWthep3cooQfV4IkFzFdCmb2ne
AOgkGU1zd+CC6dNRkxtuIYp3J+5zG88sSRADjLY/8HsrIB5bBClgDQqDGG1UaOYk
qBkzCOFAuDC2B1zH2SbrINml6K8Ih3RcEk1vS/Qmp5tBZKGZqtIIn9ZjPyFPQ81v
6P8HQK1+5wKQ8lJ5mhsEl0m2QkitMd++mV0xASZzTWrGSUfVxoKdP0byfigyMgP+
A5t3gd8aClGS5v2dnngCxLrOUYorhmAVHGJcpwisCXaowO9xG876QqbVrRhg5jJS
s2uCLfVmcCki76x3V422AIgQkm79JpP8335msk4j9+v4lpqCrPVkshK5IWmlVNcD
rdnk8wDWr2dOt4+nyMnqpAAdDeOwm8zzOrWyCPOMv39+P+ZXqsmDKi61EaF9HVEi
MOpzur7Bgmqx0b5V2yfDkPudFvBy0D8awPcXXfgRCAoIsbacn90pMEFyOGQs8W3r
wInTLtb2nrvktr3rJ5VkGaf+217Zlt54mnwGENQ9EobUmqBvTEnReGM7cJdEh1cE
toftW3P+0u0LL1c5DaFjuBw3dRp7dLqUafYd1T7oE5+ZCZjb806SYnp1eSlkV7CW
uXBEt85zW9ZDFuejU47qXjw5SeTxv3/vSNl28cAVlTwNdN6CGPJFCOTsyn1l0MDX
YDtTrtHvuzWjjWs0cLLuDGa2aphM8oPvE6xvkYeShouYyEkTb155/4vnFJfZf5hS
EQuI+kxdJd+ednrug/prqTa0g01szNMFwl6Bm+XbeB1M6TvQXlsrkGW4qwjYkh+g
326vjSY03GUsbQFUraRfxx4IcIJcfyO/rfP8S3TaZoBar3IdtomgTHT/BIcYl1YR
D+SjndgL2HzbhEZO+K2YkPYD1Vnzx5HQbXsiNQnh8tqW2dWwgkcbLe14Bm5ZkJMU
i3L/SYaPd+uqDhc/32oNIAAnrntpvBbsN8aGF2l+sYogzJw42bmY8cC3iGNYSmPu
l/kZnIykGf7+2/LqtyRiMyYbV/AF/zxi3g8JdAPIDsEnymX5t0zdgMmSwjXHw1g3
BVf+JkRMMDz6KpPikpaGxi0021N47hM+dyA27x/ZoJr1pybeaS5NWCa3XGRsoCy/
HoGok9vtF3pIQ+oQXMVXRyjO0iY6PhQLM+oSpSYjAi5PPI8ycocNO3JNLn32wH2O
jWGsIEqUcmYV8TnJkvd+FA2FKXLOMs6ig43WYCwmjZ3+5IEGanOulAEZmL2jqo8a
72uaerwq26itQ9ZHY33pPnG3eeYs7AZowFBB1z5ZDvHpU19BstrbeTt/edXX0sFA
l25m1RqHdNYR4N4IV05Oro2BCzncws3TQ637+qziZm99OD+K4cR4chvkvN70aHpf
Pz2YYanYWZxJtRIskeuZNwRNXXxskd4/dEVBU1vAresAB/fToC9sMSIrlhwkiJct
W/PTT6h0F9CNv9g1jYLunkEeeylgVsu/fvuxVP9jOEVPAF4oP67zzh1eW3mQTJ33
3xrIv6Ls77C7fJNnCWtwU86jE+hxScEddK2Mwjriz1ZdaFKsQ3u3pNRfE73Ktqrc
Zxu1TJQt2V16mcTCWbO65S4AQbqQzsylhUVD3LvJ6ofB6OxBQO/OSDTZC0FO7z4n
p3W3e4a5eph9Qx9kc44sK5sWQsaKG3WNs2ZpEpkuH1Mco1esM032Z34QAPz7Va3b
zAVXqLIUsCj0j8dtdFtvtQCKQbrUm+p2QQHxoGb5KqB1sq6UVQRd4HjeggJyFe19
XPdeMzuECVLQNjX04d0fgjvz0Y1Wy59zeNVYbhm5vLCleRMGjI+s3KLBQUGum3sV
FanU3ZCRVy3b1pkIdbb30FsER7EV4ME/1WAIeSz1T8jSKc7/jep2jocJXFRpev1a
AYJuW22NT8uXNYzmocz2e+6kxT7AKbbQfGtAG8fo30jHCj42xpbJQzvXZFkVgfAR
62goZy94j80NaDgw8/Pd/AZn/J30UtRj+2u9np8oPcGkMKBIaQqsCgb+Q64iwnjz
9uJehG3VqpgmqFEo79enU3Im6CnVPWPuC388GXZ5cvo4G8MQXNP1D55RMYW2Lp2p
Ca1cACfs30CkzAiYKiHZdIuOIyFFu39twYphVorrtpA2Q695oDXXlLFOEdpaelOc
8YAb6ie2mDBCKOYEtm/AFn8xkKzrkFM6LOT/fsw0wg1MOhhYgAiEPQpP/txEdmew
AqLOzsYQr5F60hq0C20eOrKlid99n6P0Dq7LiBAsXb1JorunCi9nX4o4AqtMlFCW
Yy02UAJJh0PiiX8fl/Ev4bhLxSq6ZpRMwJxSViphuANtAXjuAz90UF7wS+kmHaaZ
mAVmK32+vuz0sCrGrzXoQuErXHEOat6OV1yyRtr/VTlHYxVwaHrqvDH4TV4lDoJo
PnVZsHIA6W803Zk3AzdkLW//0euCO4VaDpQCX9HR/VoH/wF3+yjbANZTYd7SPmV8
HDwEJcDZvliRYf82Lj5gI9gevaVqwVDZhvtMSeOMQWBQuApSQ/5GJsyXGV2zQr8J
oBD4Wxsku0Y5st8r9azDbjpADVr5mFmnmrsYc/+ORUMMJ/FLYGSeJAImTwd+nLtd
k58JXYoJRrYrsS8oXTJcgRYsJnOBpCcJskHNcmFd9rCEl6BKY/26Euw/YM5CK2lQ
I3f7mdvbOI7G8h3kj+w2aoqaFxCpuRqDJoJ7ItazP8cgV/prMxETK5mwQpVhbhSM
3RMB6ViWbEprXItScqxlfd0gJxCnfuquooHUkAPOXkDphoAAzQcMGOiW794q2REl
AjT2ct7DGBJRiLojHlPYA35HMhQ3gFu5XwVMvVlHq42Zvk24ope3ZE4y8eXQKxao
FsTpVWqVpGRIiYTudJctXT21FE/YxDAhuEojsOmOr50ktq1uelkQaMT6h/FYR8Ja
97oaAQn5eePci+S4f0616S5KH9RP0mm5vMtTdHmQVwfIIB/1H6VXp6v2589pug7n
1+bydhID35hjpuqYqBGsJA0SxhAmGhVMkBptMUgSMqgM4BfLt7+gKS8xMm+5wTJj
fKmwAnwaWLvVtY9NFuioJ5rHpVIwAfZW5+bJ4irD+DhVBVGXxhrQnSkrChu9lxpv
Xsc1kE07MjKZTyA76GtSROOgn8pnmokgnIPm+I30N/Yjot0KC0Gcc+TIG2d/o20g
pEsNsnW61fX6U3skGsfqVm7WS6G0TldaCi9xfQIGGXRYCZ5eahFZdc/BJMZRLWqm
BZy5ooDKcGp0SeMeRLNuOdV0roBwIgA+y1tTLg6WFD0O+4d/DfLs04F2KY6DdYBX
epF7MOrRAIeCxzghH7+ALY6t66N92NO3LDaGptzGorLFnqWmj/sTqBUn9gwH8nn7
KvLumgErzJRWuRLneBpZx1TfRajX3TWj5VBs62j7xN+UDxsGTKDR0Yyr8bQZ7DMG
fLSyc3tRbIpj5N2GqLa1xMVr1dciZe1Ls5CP6c73Vah3SObFuvPet0QxcxHJsGMj
4nR7Gw6EfF0uPxUwlDT86ZZdlDaKgvdjHwUHwXjkbS1TaPBeaAllFxGHT1SNavgf
TjIA68jnx92BGiSEQwfCyM3oUJJC1+UiYIqMojtXFeoBL4TRKHb3DJem7W8yDghm
7S0PC4vi20Turs0Xhg/zz8Syb9SRODFEoRBSLOE9VfUXbUhvSHQ4p+yF2ERTIJys
W/99rV/+l06TZCxK+6K5CmdRJoewmjfxazeUYUoInf2Ze60c/0dq6ieau1UQxcMI
XGTFPL5L0wzyOwlojg0gqbmlm7SHLEyrGdnZ4B+sGdbxfotKVWvRbEHa955NMiLI
y0+BnlVUNcjeSmBeIVzv9ka6wEcsUCNEsdIVqXUyCbBBnXghaWhKfAiLCYGp7ya1
DmCi7GJItBWHhNaPT8LIH8KjaYpFh8pPkvSWkkOtx4XGx8oQZfwueBU31kFflbBK
tk4FS6bxUkut4K5hSuDNp5rTwRcmdtmgc12+W5QPcqIpnZZ4eITJsRh8uRhqyY4j
/DU3d9dvkfMKBtYRCtjVRk5FUtYaibD6WJkH8yKtOHq9CvXhKyehpspBlr6O2n+q
7Y53L7UAmPidQVk+cdICHRCy5ARAWmftPXTkqGBbj9de73CokjHUITW4e5FVmVEm
tGH7sz7kBiN2R/iC/o75I8GSaI8qdH6/irkUjcw4xwaSMclYULSwxplj7tUKNNnn
CUTyvL+R6s4AiLzK5ephEJRhAZF3dDszsbVdDN4ZDo1XNnmyubXhrXIy/q36zYQ+
vukq24AMzM9u1UBFrjaYaQzzBc3cRjDU/72+2aVMtU18kIpuReeFfqYZ5tRgFgzz
p/+4HC3D+7W1RBPxNS+jna+CRtMdy//ITvB9WT1ze1JS5W9K2+1y1uZAyQhx6RGd
vmr2af5NLq/ZaczbwWZlmHESkaxO+DCMw1rWfzjbNERGFCCn92oCPp8nPrhA+0Aa
CE3vobilvX2/wLNLRJcUopWeCEqpwLrLyQGZly0csUIwftnn3MgTD3Gw3GRI1NzP
NzkBCPjDeGfC4ZFR7+jk3XednVR8dHDX4LHiPFfEkWDngeFf8G/MqbmoVKqKOIrZ
AYbLiHjS30fwHxcWwiZWL78JiIWJPosQpDOIq65gr+F5zGhFf45XrpyOTy1c5vBd
gi8YBb5NKZNSXv3O53E2cJt2khXvkEvmQ8t6hz9gSNbrUWC4cliCxe15rdOip1Qf
wNGuHSmHN0M9uPeujhzsinDMuBMibwzIUKHq8rFWlzWlZrul+02ZRJJ+04/3jdzQ
mSUz0+C2ZzbGvwm2bl2UGchDQPYtLjLjABaoM/FSpwoUlv58R53pUYSfNLewTsMr
I9Cq7H9RHwTqIMGejQhoRDPPCfHAQeFOnq311AJ+jR8xks+vgkyyBYnqjjnsL8vo
3xFFtMOpR1uG8M8hkGzq+J5ImAE9k8a4buOuQrcRp4NqrtFwLdsKrn9RktHWatls
k0zHIHeeg6khLRr8WV8OVbmDirANC8oHHXrkDzw8okp+BdAkoz6ijJardvxx2A3a
sHRC+lHxZgi3wGcdzyG7nKiA+KU2b+Oy4FHwf/fA+G4ZcRDav8wEIsBpdd+awZho
79xD5qHXpOufeubgGGWcOOTpDYU1E+Wn5B1FBi3HieFpLoex3F7I9dhhuIl/NRJ0
YXM9uvyr1KBpIsFFK+x2CnWbbrUfCCXKZfWQYYK847VDkO77b9TtPyopzXRLTMae
lyMckJiQVfYLcqGsEoG4dIxszbN+XS8AQzxkhxNMcOgirsllr0zrDlmNEtbBpUZL
b2mQhIaMOHTzbVVhZ5ArPhPSDHNNxNC+a9sGpN2f/ibz8E3cfD/+VOOxj5nyuqTE
J/KLBU148jr+BNcXZOL4v4p1I/2YYkVmrwynWnp/ft3Cvs/fGDpMULoryjGNJb8X
RgHxm5rV9csE5UAaDeK1S2c7HkDRyZRubFg67rVYpt1uzdOouETdPkLipGH6N+tl
yJQn2vh8ncXBbE3CO9HBwCrsHPiNvzkyQaguh3p+Kk3jyy1hD4VRQtHcgCFyu2HK
nFXBne4JQjc+c54qW0NHlptaFHO6V8GPNGGVZQT0NMvUyvX5DEgjWq/YkGOg4rho
51BfVk/j0foZFkYL5NofzjvfadQZIVTbcqw96FhC8FdGrgr9Nbu7xehexl72Liwc
cz8OWlPPOCLl1nAadwElfCr0a5m7/9vRyLCeLmuT5uXs8MIX+4seeCh8Z0PobP/T
z5tjqZG6IyOS9JDneMvp6CoF7+61xzkopHyN9p65sj+Sp0P3EiAtyoDSJx5L8dR+
h++bFcKXW2VMtBr3B6+IWLk0104o+vlXNFANlt2RlUpZpFwFyI85EZ8T+O46GZaT
psX5SWQ5Jr3+aKiYuTfeAaXHzS0P7JW86lQ0KGfLVhoObRpY5CyKlLJpbfYFVQQW
CRPQCMvuIZr6bJhfxNl6YmB1dSoua5q3lULW9UxJl/p+rEL2W8PeU6EMrtz9j8Lc
rUQazHVyGrPodWPJ/fd8MViq89E01kxDgBnXvRP7DTrXU8/VPH+8SJjYDfpwPKLG
TC4Xm5Pc/zDX53zgUXo4yOH/93z3EhDkI0XQFi+xtw/ojfiQqwfWoYLxBH0w0EgC
O6eC6MW2edf3FYJ3rHl9bF5+H3r6WVw0qR5SAaNKqI9TQXQaqDuwveD/7TOUQ3Bu
Yh4bph0iY+vEaVoAXnQ81EuMWy5+za32fwbNsBG4Ztr6YMXLYDiSca3fMqc30MVj
ZcFDdlB82encc8FlkXeTALtRBeXhwy7oQWlDnqqfka52wdis3K+s3LXSb9rQ2stw
YEkeBvI2nuj9vt77irlsI61uaAZZT395esoOsAmKnM7cqw5WV6EBBCmHcS4O9eov
V5e6ygy0EDlyQE8rNZ4aT0Dto/Lfzi/tZo1Kdn9MFef2nFoV3n5Xvv2sDh5labzq
AsCBwQ7k0J1oEzjCxLS33PO8pw9NRu4ysqCthJ3IX7Rcf05KVzVXHx4ZhQE6sd1A
M0oWJDqTRHuckV7EqD5nUYP2JRTrEFqRHTyyCxG+3+W2Ach3yjiwWKJYZUp0qgVM
jkeA20Td/219OigW2a2fXHUtwomRZmlczV/BzD+zByy2p0PQHkDdZs6PKbmJSipS
qnzZnLqUtNNxAU4ni716Ep9rCfrL8g/1r+HTSnQj2IOmvRuSSNYPj3XNKsgBIQm+
aXHo7byCLXmSyKLztK48+xZ3cc7ENcx7wJysyWvA2+7OFgxptFOtC9U5SmFmfnvF
LtUdJoLx5lScUipfVUCo0ly95dmfFEMAz18PpHvCM+Xt6+UP1Vcaj4M7jhuijoQx
gFsdDSd16Zw6J1e4zP6QOiBsK+GJI9SV/LAHfcvhP3U9p6uJl8oPBkpXWo6mmIF+
maEf+clk7KznEcNhh4tAlh71/jSMo9P1U1l9cVqL4+a9JjTPkcDMicz444DYnayj
an1Uqg0OWvuxrjpjVONy3KLwnOd0Ch1E2cgZCW3wZZqm0gU/BxYYO9HazNBbKqC6
LgBb2uTrDrUKC0/BYDheGUDjqLdwBc9EFMYUTpwhy3uPmidmXDTmXUI3GYENiROV
jjZHJINevjtXtKuA9F2e936MllqKNzU7/Rks6Q1P2A9MKVEpREItGAa3Tcf+yH3+
SltdHSX/6Z1zTfJFQt6CNQP/IcEjHG7TbBu6+JBtf75VdLqzgdoS2h1FeKDObrbm
8CRNw8y7JoeyCxGtFm8b5HABBKQC1VvsQ/KfbtH7Xe/H9GP18Z+UmuchdsS9k4EN
DHsVbg0vCvxebX87Cnwl9XPtj9D3NUpLU0+Tfi0BNMiF6dGIcaGKn09x95DSZp/L
0soyexOJ5JtDwquTs4VHvYHZ6uybROhFZ/HRHeP9eM8sZNWHCQWxqGQjpIWTozlq
dlrPOsKiHOACcVyh+KH3A9RVriiMwf3hZrlFuDY24M1HNBZcAhENw+HnbB/VE/w+
3xXTAz+evg90RJlpqp3pQH9r+Ut65tdybk/XqBPVMq/RCoJJZkBmEW1Ca59YYnqC
LzvqdsLzOvE2tkqQto1b8OhUHEXb7ZVjtgF1gY/jfL8zd+RRivrqS9rv1AloKiTb
YcJt79nAAwqdyKLi9oL68xGpUeceS2mv4MxcvF30OS75hatBI8MjyMgv/Ka6m7cQ
2RnQFGrNqXWM2taHA4lOtdzOLXiLJJMco8AfVUBx3Bk+4qukTCxrxbcTJBFzt7JK
Lb+f6+VgacbcFRQQv2O6b1fGKldzMBuDC/bmtQDSrJmDyZI7kx/Rlltfbrk8CBgc
kL+5Orf7St7tBIDE0gRZEmH3YwomfzjzbJm+w/yf9HhPled3ul6QQlLGoFSZ7Npw
6JDv10VBpeca62esSw53W+Xro6U/5iQ5SQhCoiAzGUCOOuizV660Is66DM3qfnlw
D7TzxWsm0G9JeUrd8EPn63s83MA0H5jCUyty0zHYlBdJruvstjw+ME/9yNXU+3K0
EDwM1eb1juA0H+QGxXWABK1l+QfLgSHXwAO1lJrQUljVPCVGntAOvlkzTN37NLM+
CeY1jt7e3HUlDRnoq3ffNwDeVZh7dsJa+2uX7tHsZbtpZ/4XyZBtk8dsAzxnL+jI
nKHF/KZPCbhNbRUBVCWyYt6Kwg2/QjrlKWAc4HZmktXrj64SsWkw9I4S67T6z7J4
tXKu8pWkjmiH05rdy986cELyIjNWBXzjRmT+ESxAFeyNpSxb0/wHkG1tl495dk9q
SlNsTAj3rhTyxU9dmY5ms2/q8rFVD/4utFgd5FfD1Yi2t3bZYEyB2rlOtEzvxovG
P9BJfm3RYYGAgzUOU/yIalxRyReh8OZ9QJF6QoNccUAFutydEtQv8OXYuZGdenGG
SpgEVd9oJ+dptk6cSUL3VO4AWSlYgWCjHbByCJw8iGrfKrFmfnvjL9+/kmRUwFRD
ChUAMyOo6r1ve/3fK5huCLSjVVT8pbMfrZ9gpVdZ9YtxgDdYSDjkOINYQp+qx8sp
nZm6AVLpYq1Oo2pKyM+uWuBbRpX3D1MpYfXoAJTlNiUj3DBygNZZpYjczxDz6w1C
s1cRlAv5MV98RFZT4F6xpkg7kgw4j50j5LS50ps5Vz/Xao6/rOl6YGsS8Y/YoAIl
ZPH8MzL9/bvyPpukjiI46p5qOlulr2d34cgJA4HtvzKseSF/PP+mqXW5li/4QxME
Hq6JY7LHdrpQu1C2OWQ5A5ZBXBuMx5EYfdjkR3anra0=
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
c7NcA2oudpvRixQdRfhsFuY88HMENmfIie08+o9o6ugIqLDdPIiAsiA9lVUuiorD
K1ZC6N2f2Vm9bGHNtNL6Mqf2Q7rI2QiKbpaqECigrEQpjXPmk6yu9sJdIdnMVEFf
4f2JRNpQgBX/Is4cZJDwOLyJdK0Haw8wTPXNr8a5qu71uA5GUJJiApFehQ+ze/J5
58znY9Y1nHgqSGFzliHvZxeLy3zpIIhbkQJNyNjmTikj56BXvfTOQ9pJMT3HaZoT
jPD7unEs9daPyu9aGT2+hgdhR0QbDYKx73ytFHmKQytn/5wSHKQxktoENv7gDsur
0aDr97RkDJx7fIw+4L7dDw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5040 )
`pragma protect data_block
LoFYYBKyNabkyR7jaKJqmY5RsuOwqOxPhu8Q27USJmOqE6PKNfjpowZwC5Z4Ft7J
sIKYzOrv3s3AFRdkVkn3D0TnCwI449Y3EWXvz8HDLvE2iKKR0QE8rofVrR5sg4g+
ACoQWL4dOGqxp5Oyg/Ac2j7J53Ar/1KScRiiB3zFhVjzJZHRHFZBw63ysYfadpNo
YGAhnYM766tX0QtmY13Xa6mTDS+aaaza7fZgtsP9KBuoYKSmAY22+1aEbaihZzoR
pz099fIXQGgNOmnsnSBK2bSEyqMdsRa3Dxh5em5usoApGwCFrP1jk/QCoTc9/JXP
O/5Br+lbGE7M/2Ad4i9+JdhHWbHFkxx+nxZTA70dcL8zcpV6K3iFJrn3zzdnP0p9
DUbsPG+0sdrNdlBec+Y5xbzRSa+9ok3aIaj753GNtb48GGsN+Za7Dx63xRU+lXiv
ZmJRAfQEoE+joV770/tP5odglVsJnBrbe6L5L88v2tujmIAgniSqww31SHoYDkJG
WobVcaShW23p6vEuzu7ia000b0WTNAiGOwzHiXGmuLHEsBMa19ZGtwR/p9v7FMwK
taxHEvXr7ASGBzhZjmJeXavIjzHRRAVrOodl+lPrZX7THbr9X42pcO5frYZcTpXy
F8Bh/9DSvheozjsZcy6pFx+jNx/Lv/TBSxyTO3V9+d2V8IgD0OBYLPnN4WeTv+CL
EfA3KQE0m8x9G10/xd7s3h6dneFNoq798MMmeBi+ofckhiNkXG3TJUqAsuUTgNHL
nIbpy/y5tsDGQyp6OBcpHn1VqE+pMU2uqW35rvC0vc3XHzhseljlp9LxIRPFneaB
dXFV6oOnIN4OZFSUCsrfP5UGIBu490lsi+Kz9CfcxxJshAoMSCtE/Wo32XNlehRO
L/0epPecBZUc0+JjAT1TbBBCCT2vSwRJsUVbWc7ajOYpg0SUyQMyTvcj2rvlOeTD
hHd43ZcamcEUivnbC32MsLX4LY8ytohZG+h7Q3emxuZpuAZpvOWNnrdGO+Dbw6Oe
wL45hPc+vZyCznAZPrBZur13g0atjhRAG6ees4l2+2bg0Gh7BVqthS3HbVYAHjEw
ZUHPmecz8esJwhVcBMXCnh98dKUWqMyh7rbNrOK0DR16c/n0RXHRVJxbzL26wTjt
PafRcGdfiSZnMxhnqxqdj6nVpZTQui87nYdOAFBwQqIpvH9EqFx2AJFl3gtUgTdL
d+J87yQ3Fwo2329wOnsvHTAII7U7jDqpQrgyDVRA6TcdUtDcmmJCEtE0jd3UcuZt
LiyFD2HQBA6sREgi7vPUrGvJ8ZiMZfdkA7LC6Md5I4F79uv3VYJSMZ+C5zkg7lcZ
vPcm271bFhFWONi+iZ0dkDnGgvBJIuNP9O7iCYBPiYHguvC0X+2WTRO9eZSepQCw
UeTDx3CXPFJXAWLi/f6KzmiKILN6wArjrCCRgE7xan2xMePvQAdl2G+jgiH8LE+j
cWHd7j4UPbn+IyI/4AL12mxKqECyyCd3zgC/Va33bAaGRWmOwh/2pf6T/m428B40
2oftB1BQrsJCK6+IeumgEOESYfcXTP9dbuFv0R+tJFFtxAlkG9x62sbOklRtu0Bw
g6Dff2f6tsjZYmE/PO55QlbqI9TrKLGDa7Yx+9jlYvtl82Y10oV5jWXyVgYwEmxl
UEUbqHU2VeKbmRKU1avWsD5mmsbNOVScQaDTr3RjaPxSu/pxZFZeYD6ZtDZDgHHF
WzcZ4PG6iBLRCmyQj0w+ztUH97b9Zq+5q9KAcbEbRt90asZNiYhmOs0Qp1/UF12B
LTUzgkMNh3TMHU1uT4f4qBkODW0cY2CQ9ZZgFw0TvbuN19ASd0EdE2Q03tIAd0QL
JryxWcvg2lwJpvzf5CzwJIJ+WX4x6flPqenjvMc9uG5Nav3YnM/Y5Tm/4/qTAxlB
B9R6LRpD2tsN01dyjWerE4ryUYvvvfT3m7nWIOiNQm5H+N9LpTMEibWSp8qX5lqz
+r3gAXu26smtGT57BaPZg5gIyg+tgw9R0wOd6JcaOpaESY4GOJWtAe86EZywTKZp
n0VxKq2iiTId6QvsPH7lBx20uLssqP/4a+LVd6fXQ04JY6SoapB+IUKkmUoGG2uC
SOIZe3RvJq4GRKckEzr1dIZ1g14p0m58yrjMaKp9dBLkioaF4ZKClzO7l24uhomF
2kZHss3e7/ZYZjosLd1SQceJ+7xhlSJcxU5fP/VbBKMddhJw9MMEOSPZJQRHBoP1
/eZ8WH2GeAONEBDeUEjEk3lJd8qGllMSdUVx2jrxv7PFwvAcoed+RNlT/FssjQJO
93okLWbM4qhz6C6lq3SxHQG1pT7gJoNststF1Wiy4nTGsZ7o9oypn4jKGecu7CD3
lvtUlI1sFKTpXX25OYVAGRw2Vi/JjGuYVDoKXyOK71xDW/gHSZgKGW+oMmHB2cSx
lVl1COJ831540zUbJNto+GiL8HB70W0yO5VSQ1fRZO7FiKI2O/NW8Iz+Eznbk/Jo
r8ikXbla3iMqHrkKb3haBLMoigbLWAwVzo+6fvDi0a8Wlo8vonBDqHDiJ+CHRKFg
ovvxOgLxmnvnDnKM+pyn4f+wnCHICRIiWw8wN6tTMn0+aXi1zUWpon8xDbZNJvj2
4naEamnX8cJr8Ls/F+rr0kgw8nmMxKA2q8i9ubEcrPE5igfWdC2SCxx4jhPV5Waz
A1l5/ceNGVIIEy156NagoX2mVXiHYeNkCAWPMz3T4UAr7p4PCviI0L2KQV8Lzuda
kolD7deFKcc2RulckihrAPHbRkOPaBcOwE7Lfjo72+UZ3JO6S8M7UJ2cDQF4M8H/
KZ+VN2eE0KJzZ7KyTRTCvg+qrUI41S6ONF61hKru3giS+znngzkOi2tnCnchiW7D
z1bY1VbRHA5E2DXlhrUDEJR0D0jNx762i4UEjp5ib4luTaKoXzfry8e0/7H4pG6P
HioBuLe9LCqwsz3+hTazAb1+/Rg1DBzagctjTJuVUVvDhySPSs+ryURjKk+eK2uz
PUBPxJ4o+8GY/wqeXjUbzgFcpFzWwJ3Zbvz732OQ9+T0x52V0xFdiip5RT0oOZQl
PTg6/RCrsjtHz9MZmLDcYeeo9NbV13uxZ3D/b2Qc9pw8zyWkQjgVcc13G6v4zx5D
iYiqzoAUHKpECupZ/B7+9wyZvjeFEucXAZ05bGCyIm6aNusCWB5xa4/a8ORzOkc2
0ozaAbGqkUyPrTMlsQ0PpP4W1H9EtyaPGlRaL1wUE9Eh4v9C5WoLqNWNiapu1CHp
WOrByB68cKc8UBRltDhwClm3dxITH4pluFVRG1H7UBH/jb0LvdCLhj///APOXSEH
NVCUizp7sZPy2MrU/DxmiZXGyYRmmFQ+zwVBsh4R8uXpcNhwTXMfOZ/9LLmDhCUB
jyt2BLG+pSKKnRqhbZyVcgUpReRxtD2aD9VEc3CWANLe9Mj905VNVGnRc0t+PxLJ
4CHbLvHs5MlvgEG310mrxLfXIDngStS420B10nnJbQhZJ26ln+TnRNPJVFabB2VG
N0s0xvqzT1nd2jaVDKWb8ZCH+/dhrNbfDx//KlRV/u5fovXuw+0sfIfZIyUfiWxy
DwwuG5Zp1ahvJm3MbqjpivsXeb5Nzis03tSzIeBTbpe8ywelZI5ruLsJ778aosG0
DPnyDSFtru9sOu7s7vqUglXyM0iospl2D7k8IvTag5ruVHdULaVsR6ag2gi5qLck
6rfL8vhQ6YV93jLx+0Xle+AOSQhGPGtYQ5oZkWRJ+4ZQa6by7VzbYsHFYAGOdkxE
hDjM9QbE+qZzb5KOgcKEi++RIC9vJCn6Lw/YYFxSZZL0LSyAId1yF2D9UToE/2gc
hvZyJRvW56jvV8FQLo76Bubqv0LJg51NT9aEi0iWtFwPkv/vE/PfpV1GQJOxNTxy
t7PEtbdiITpnrYIpRzRWaSTHGsSjqw//dFCm8I91YoQwVDy4wV1UnDlLFx1gCA9k
5hoGhkjFnyT/ZTqci1qazOYOgW1BvA2HY374CJPbdl+BguF8ras2j/8sN03uoMVa
5EUHqj8Mm3VOXhIIDhCm6tP11ebnUvu5T6fs4yDCAvhWalpblxp7rxCcVuad6+e3
3M+BU1qgHEoGzN0TTuM8rWHvDz5s9R8g/5aTgJT71VfwmtLxYpPDM4cCUPwtNY/0
epeuqBSJ/ZGf8tBAkco3svLLL9gppIwc3A4pXeY9ZknN9d2Cglw1pKkpFFw3lyab
ZZZf7E1caG2GAWL0Y0tBUTmurQz5sHry2a11olhJ4leAnf6pK7oiweTwjNmEgqQO
dwWDd1qmSe1OLVR2yQLRh/rwWXz1b+dUhhaHcUHUqnIC4XVAh0qKXl57YjkFvPT1
vh5ktxbLrN0xkfv3lynZFO4kpo+mnnWhTarGpu6YFV4kVQ44HYDKo/vVQ4RgS7TA
L5xCuNZlqQ9Jm2H+LQKa1U3H9LfyxsALZM1xEPPBXfvJKoZI59E2oLIpUswXSgT3
D1DNoRLziHxXL9Pp9C/U0mn0DQIQH5R7TZLk5ZBhjuGkZlzf1Vz+wdvpZeWPgDiv
D+V4CSPDUSe5+jL9DXWk7UEfOc/JhWMurk97MCSEFbhWQDzFuwodqY+JAQN7Jyny
9WKqvXVcKBLFr2naxu0IHykfwFMI1nJk8O33LpyEn00qGAUKh38vnvMg3bsOcxUA
ACRhWf653k8q+yLXwutJJHWxvtqvI39AnPfS+R3wDhSBjxUPwfb0gTf4ErD68OuL
7kRerGGyNucolVXYsqUbU31uEIgXXTVX5oVfusJrHQaMwz2323SixWKo27N+2SLr
QvbAYaUd7hCPxpE4NhUDJdEcIVUhPU2L+fvhoGbGhpXHlJZPPHBFXxRg0wt3oVyV
QgzSEBCWoT7aZtx6JgJlgGX3evLENzmQA73HZKqKj9LO8eS6QMablPY1TEID6ENq
1f9MnCPb64I7wclMjb26+m+nSlnHTzq6D2MayXtjptUJjvcfzNSNJ3RWtVuD+rWw
LIkIBj49xqTK8GrMDkxry8NVVEB2WH1SW1ircsmSXzoSsI7a29EbXWpSe4ggEmge
IGI4ew7OBzvCsD+KAHAj5+afHmgJMWpgVZnat4CEeNrpoGrq8X2CazqTnMyCccQT
p7EpWC7Bif7JziiwJT9V7BwuUDLPUF79s1prns7PSV0junujFtGjHuYEwrzRZN6m
ISvVMG9GQ9ZykoqVnrbJu6SXCbrkAovSc7hyF8nXi0/H7tIphzFcSYcF7soHfqAt
II3XlBeI2OhVH+omwQCCSlU6/odsPXjxeY44xgASWSR3yjYc86LPCcYaKp8jRO1Z
XSSMi1HJ+vFA4kGxp4IjqyVd6b1RIZw8FKZpkEHWEbT3UNGGT/i3UyL9vcYRACRo
x/uxU0EBUIlHNQFN2cK0hpIwxth75+cz2z+Ev1AVQNGHpZG5/XMeNvtrolpbWhCE
tjOZ7Wl9fgMtx1zKSUSIW6CPXG4lo/zqNf+K0n+ANp1722SMj1FzyyoN7YWIduy+
hgcL+o6tY4MPSmTl335bGa63DJl0ZakLXRlouW2IMwFpR4gLvPVmAqi6neOWogSX
cenEZqi7O54f6hMe/Qb/jD47+3pULBhP4a/ALIThDHgeqv/SRczrQ51oW0VXt/XG
XGNhwBc6aWkSVU8KI1Wfxsk4vmPNfC/E9qjG/ZpSZy9vA8PCCD6msQpzYzunf73/
LuIzYneBcZ+2s+eOWIAgzU2SmOWou4Szg9GWsg6SSBB7dq9KIv+Rfp9VhoCI+k1w
0zQp0J5vR3GklNqgE5oMF6VI4Sl92ADyjeHF4Iv/MhWrZNYWgFdRq/4VSkz1zV21
rNQkY+8xClIuU37Skwh3b2QG9hbPbDFV6FbKkN/GeiCVl4GoEbVoCMc6rFvVA+IS
DcgTL7vPufSzQeVrFkkqmrlWcP1RvSc7E5xS+TTJAWgV4piSxxUMPXWhkHJWtMSN
0LSPa7qP44W/3k+D7Uq02bT7Wd964tppODRvFYCTPbP40AR1BLUG0bOMhbEJWrPq
a61thblG/nIRlKd/CpcigbCWXutM79+dXZpv3Cm7dxJiJ2+UXrhbNwgNSpR24kxj
P63F9jCpWkxQ9P4NSoBUCfjh4tgB+juLXledW27ZfrF8KbQAoGgweVGJqNOA//C6
U9IW0Ehl+6G92Tdi1WowsGTcfuzv4kJ+lEwQfCxeWMpeyH6OVLG0SmZgrv+fa09j
da9Df5VNrZUNDbeLYzEeBX3vWwQbqnBhT0lP+0uw+YpMDBXBleS3GHIUMvdT4NsI
j4Q35Ra7I/64ZPwuaukgV4ZNJDP9HmYUmWT12t/zzX0ZPAkikd+bklntGHce5dFK
1249Zq7NL2fxEsfyFF5lCxOjqA/RvI/bcWdIuKMD9635UI0AmEChzB47MO6Zwi7h
zAGXNOcZnO1bhpqS8nW0hIHT3vcXC0+E8x12WXu1eclNcFxxIGfwu7eBG0WlaRjC
1bgVCzlc9KDoCl9WkUMrxTn9PhD0tpRZJF/MYuAMB4RmlKgkCnGfvWYXMMIqVX4C
mviT/obglZa5QNp+e1eXaNQO7O3OP7tPMty+R30jJjAIsY7ulkG3TQibYPd9DGyZ
N0zg1Mb8NoXLMUhXa8hOpglHburBUHWVaYgwCobIXN4QulefFVldL4YQSqrx5rb7
uLu9h7bWBtf3bm74RXjHH0mzrzW7Ef0x6qsxESx5r+v4I2b4bQY2JIhTjmwNTQz6
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
kxNntTDgZeLtuzwrQMAqJbj+Pl+45t+dDyfumgIctwoAxa1KhJPROOfqB4gyuuyo
lOyuaDOLwfUnv9gda9Adit7xTcXdPJz+HGnzptTmc8hf8KpNucHpuui0aszdV0sj
bBLJj+Wp1r8XdLLS47Fu/VMT7RTdN8SlpcBP75ghYSifh6tXmjjAh1D1OHVkpyMV
G/hzT4n7ORCvbO9+VMyYZWqRdgMApiBmv3plqKnlnSfvtMkhMkRzwlzpMLi32mkX
m3/CADwr2Ur7LGf+/Q5LmLdZq3+oZrpdyvc/6vNZo5U8ZBE2KSp9QMK6aoEcdeXs
3xkP95Tshoj8fBnnHlz0Sg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
jva446sVBXkMe7jfczPSmYWeOJ3gGF1Qz2mJI5F/FCG9zPnGq8kXb1J5D2z74ib8
8ZKa6pmGQ0Zxey8ohDGUgtXpriaSIRmwmltXyN6WMplG8IDnxoTW8DrcO+/lYTjn
JypYyHtO2AkOBVZ5lkwq3QvYKM49eX3xpXMpc1/fEfZxjl46nI7xX0abU1gJPqaF
2zrour5+S8jmjVfEJa73guQikUHwnfZcBexNeJpEFXt/26MQHWeSm+8/vx3bZNzY
9cT8LjagEtXXmBrONX6rgzJGiebxL2U2EcyZzyNZH6TMAss0S9sjDeJTepN9el1v
JcLuy6JyBdEGhhMPWf+qc4SDtdmmKnUjuFLsRTBL4ifZb/kjcVJZbMg79yhIFn/k
qxycPBun4U47TI+9LbA/kL+GiDZRdRpU31Yow+mRjV3iZT1fpPOfrmznsvZ9+sL9
sLOkaDQqTOrhJCO67zmt2j8pFaSANxvOjFIZTGtnXDle7TzNLc1c+UmPz5ikioAM
cOCWwLK9nFlkuNhq0dk/HeyhJWN+KbhZ3JyzCbAJlquYl2QeSxusLRLy23AgK6jn
Hq3G3xkuGw1guo2jTzqGOtISKi4oUM5hamKdnmMKl0Q10PIO/NCow4O1+OqKv0BM
0+6gW+WRmyTWunO7edGFGGTUR/CBYKb+CuovTXs+8L39XO5UdxVZXwLL6S8YcBLH
sR7QBHIHdJZvQ3EfMSlgFm2aJ+/MmyWyZTt9hXYobYC38xRYsmDpSOAp8vmtgbwe
PYbgaZzdTijBkgWukg1PUCR7/NpmpKAmQ86x5PtzJaux2SrsaeZ13kQ6/nFxxHRI
6Ran1YVAzQYoeqoUPPW8UoUJda5FOSsnYEy/YqaTwkqNQVmBQxw6iNOGyhTeiki4
D9ujLUrYNRu3+Z24uws0tbbyuf6sthWK8koKdYPGN18=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HC/FMhrHkf9iKglP7GJSqh7Dh8orBUhsQ0qSKcYIG6E0qvUt+JCrbJFFfgkTJI+x
tCBaM1lMfUqsBvjfcgMmoOuM/8akSPVSHRFxuP+CNnvueZvUnW5IURgX7klIX5/V
z/MrL19zpjKzwJBRlMzNRntyXia2YspFiVmS+1lwQ5Qobxn/XvOxsQwwJw+ccrYQ
7SyuFUpVxfWX2FXvf6N6ZxRFyJhNmikSEYg+UoXq868bG/PrRwq1G3PKZER2O9P3
U31bDYtHeLIQl6Vv2UNt6BT4G7ZVULtm20g610LvjxSGlUEPgkdLBTwvaUuzLfM4
aAlb7JTWpDYnn/KqCKbVug==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1792 )
`pragma protect data_block
fUKGPT6XI5kX1RnLybVN626IhGcxoktylFfnGmQWfmXS2V5vF747dMvj5hb13EyG
ImYizZBuMk3frXJ7GjJnaWl6pdmM99x3V0BYsGKur1PPGYvvI7ncNYn+VM5A9jQh
GndUfFCxNsO4FTk0pl7/wYuHn8P4GecY0JrYcO9OzMaNsTwgVjFqgnxYScgo6VFG
1ILNZqeMq/2j2hE6Gn3lm35qTSTFRpVTufV0GUGkmPu1JoQaEv4i4qY7B/K6KZTd
hOvag/FhiF3GDaKBlmATW+gMNKQe5YMBrx6E/B59YdsES7ZzYLAJpk0Lhm1KPnag
mBBMu7EwRiGia2ZDvMC+V69ym/jt+HeMzTS7GaOkghaLWzO+qXfKn3GiIhBRMr9M
GK1yIMkyiZbKM3lpQ8llJZ0Xc4iHoHEJyjWMwFPumMfCtwkpLXR8BtC1KSQQL4vu
EigOqOFsaurLCP5Bh/RGjte/rSXswHTf8mhBYB3D/a8w6o7m6QRITYbzJ9F+VmSe
di8I1ARDCv7YdDr9eyqH7DD3bduKPlIJdhc9frIXBsnhIEhhvX5MHLQhbRI4qsjQ
ZT4YISd4/YofqetPbsiPeRl4xFkZEsuuTqt38NlT1f4wrhVuWL6qNSfXT+9q9O/p
LMa4G4RMxOKNA3/6/qcR2/+Lc984xa39ZbHTE5iw9mv7Io1MCSIQx4lLwSc6N6Aw
u9+G1oJy+a6Gbbxt7I88mLtjhWb5HNGc4m5AcK0G1bfMbloq1QXnVK26UwDAErZJ
X96vboqaBQqw5aUxAse1cG2xCq0iMF9PkPZERkKP38nTuiCLF+vRjR+0pPaCs5ot
mIhlsvEBu/5wsf0qZDnYtYVty5rnMNly/QaHCsNlbrPE1cpoXJyjs1NItHtUVmof
eWL5tMmTdmCNVoXBONnvJBKvKMvO5M6Sdb6TKvhXSkkDYpbKFE0vHzl0mPRHW5g3
a0Z+H/IrmtG9NYWN3rmDaNBmnd3USDTV87PjbKMZI2RNPcWa/Fva31yoz1Xf9Svq
+a2pS7MbkhUzT+eUB4GhKS7yoAkIB/7S9fWXCilJ9JOmU37iu1hlRls83ef8AQRf
Tx4NckxiA3RsbnGph2Ekinsy9ZY4vtC+HQGs7kn9w5JULWhjX0vrqtTdXEFX89Sd
f9xY4j1vBti35PLqNv9xARp7Iof73bC5tHgf6JsSQVMPMuqXNVyQRDGzqWFFcxxx
N6005fgIVUDUYwJwbxwxvdcCcdnpP7HilDgcSH8h3eI/g6kc/P/4plp5FtR2KEfu
1bJvg+Fuqmtpxm9zT0AK2pS1iMmWSEOam/4WYmBjHvhTGyk1epSQw30yAXQsiuqV
Z0lVzlZB67xeltahTzws0VGVU0GTDa5Uh4qoaMPA4Yq1FfIFs5FWGyD5/HX+Sgie
pMlfFCcX5DcxIcQY4CcEjzNBIuIImEE6h6P1gT/O0dEqvjOyymq2al78Kp3cALEt
Ks12c9Ku+GdkaHfZMnmCp6/izqRldI7Iv6WMHpH3+w8CLSBb9hYVlBqxqXdiT++Y
BgwNMtrvImb4sC99aq6BRKz/TNNjvzllLR1EtcxHNtomidSRAAxeRq/+lHuE3qHT
rV+3t53E1zlPvkcAu1M8Wkgdwe0n6D+RIOQZciYHdBUcv2GBjhhe4p43cfQcPYja
qyaScf4WOtfGup1LvDquYJimWIf4fctsNuGYXdXG7QwqYIJfUBiTuShVwRjVkUFc
EUaPmEeHVtUVNs9Nw1ZeuGKD3en9ySUSGSp24q6VJF0o3pG+8jYjEcF9ohOKKaE6
kF88L2UVzQ2caJnmU7VBm4zmkAzWZ82G0a6WI9F+o2neWmyzaDnS3Vk2a+jQ23hx
wvq51ZlLYZNrZoE6FDTbF7X8FDJRv5m98bBA8JpPo+we8nnF6ZDRM8eQYWbF/UV/
xunqfYJornRci1Vsqai6treqgybYuxHi8BEda66fu2cHzOzq7j3x8ogJYSEbtMHs
mPodHcKoDZcWYLV5Esd2o/1bqp623S1tFRnaOYqHh+N0IIFzxdEjJ/dg0/F+Cgbr
4kc3+XsqYhcFpOUcSWSQ8j4gD+Gqjt7aW8ojoGVpB/tC/e4urlQeW1NS9yOzQADX
9EKoTJbe6EflqV1aQ3LtZsUG7Ejzvrl5B7WAgVkTA8XJgDJhFAbzFDMmZjIuDyXf
6b5M5ARydDGmIwTWQ+bvNIbmFiqryQit6BzaILMOLZKkZSbw1xB2cLDE2izwxo/d
DVuox7wAsFGnFTOUiGF5wz0Gec6448rK9VqNZQFiJbD1BscAlycRgMf4K+S1UgDb
XDg6PPfXlfqXh51hGElE5KXmqKLpJ+6r9EgZk7+tXt78VgkmLHUvUDjxBqbKY3WL
J1QPBrhpDoojBBYBQ4vmSg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GFPbhCXT6nCzrdkBPMQdGlRD2e7IcW3/i1chDT9KiZPqDJen8jMKsSKEZ6RGU/fW
7e1ghEmiz5O3A60AxqGUbIens6F6SWPOg0JC7JSPpww7eiIGNmr5Wlx36HHfbTM7
Le0RJ6pcY4R60aqsiWG2TQEnD6AvGgX7YUOskx3sVwpwDm6bMjo20+misTcc9eLv
L5gfaj/OYBSPz8NDLpy8WhMAoGEOtuTgzyr5Vf84op5bl40EpER88Mkhpo5qDNrP
spLMXHwNjfIFh85BY99RYe+yy4tjD3peq9oUdO8TNxv/+KFn4Ca0yqBIXHLplGBW
L4A9HgTIY/M4ybwUacgymQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 30960 )
`pragma protect data_block
g1pd5dWdBxgyjxzWvZW+0unsVflPGvlhTtL/aYKbmjCYGnrda6lgtgJ4rmbXbmgo
04QhzdwCAVQtFaE6Xn9V/ZyB9Lc7sSFFFuWlTLhvVCC1/4hnQTnrrVQMsc/VKkCD
4JHmlZS4+tP7x1dVoBqDt2wuutbGCl7tIKz33sqfYDsJXeDYGh9d0t1dZKV/qK4y
XwN6PXRrjlnCDm6TIpv8msGBEX0H8fUK1ylkLhdz4SlbcFKT0tLup6TaLqDVHOmI
0AvdBAegPVAQc+Ym41zdkn7/RUXSW8Jv6BLMH6eBCVxIWgHUoMHUDl3oCqU7grzW
49YZOO7m4J3Dsbfi9GVSmk6L1VdcIcKqGy1FhMJ9BaWV4PYJ6zBXyIflTStMWcn8
32w00qtBa3ylbK7HcgENFB+M2eTuI1NTszzrd/AmmCvoR7F/DwtRl2hARLHznQx5
bglhHGCsZFirO9ARpb7E1j/2Yj9JfYEVST7AFYBkAj4Yut9p58oFd2ibjn/mPG/9
2E5andNf+5z2bvgMEw3eCIyz21Qa3Zr1QXjgV7pewaU2dUO2PrL7QZVG4FldYMwm
t3uAPMyCAITJIKtcIwIGN6wcFkGHyioNTDil/WeyAp7yQ3yb/hvFZeVTMv6N+DP9
ep8y7QdBwVI6/lvtCUMgCExFw3W5ZH7woVDxt+sLYBaxJ9p+1co6s3cHpt+oxdDH
t82hbmeJur4X0iqKxhwG5gV1LmuqPnzEA1RaWazwhBWTBs7kJxOxtsM/bmavWn9z
YYT87SPZYeAmOUtZbVjdrpb5W5ntP1LXkjphkIR5hu/LiZhBTdKUq3Dnnqt+s7KZ
ownhFsQef8MFCpA5CXFYXF+e1Kdr2Um4jYbaOjCnvM7UGRfiLXGF0N1lH5DCDVCm
pLonbnUrGOkAD1jVhzOBLTOWGFGTjKfZUdzJZ3HzgrB0p6xmmFO4LLkazh51snQ0
2I6PM/elIXWliJpOoDdNUsIJM7x3LeMlr7Ql5L8TfsDFmejkS3BJCQWZQshmmiMr
/15oehmaKmAWBKs1K1WQ5sS8+xRtd8mVvOLYHE2rDWdBT6EJOJLHFji5GyHamQNx
YMXaxEvajnZJ4wIM1FTgLP8X9R8TUeoCcjb229MZdrcA3PcKAUu9vA6nSU0eLTva
91qtjcKxWAQ7AgmPtCWAHMVVEQcFQ4NR9QaKNrtbdz3qTVIUjloDJjvaweHzdzCx
OBzBV+MhYrwQe2TjClcR2ZzUx7oZyNVqIqyfF6lMdbEDxzF0igyKNsuSxyD7O946
tu75P6xXkYRH/FUwj33lovDqhvKnmzqLsphsH+GVjo1ouaylzPW0cHG/LYPr3dI9
2qE8H5v0QeqXXyTGnCd1fNdNr7HhjFBXarnkDQWFtP5qAkMsEb941NqeeX8cwVrc
THoSk8caE4wxqIpfTniu+paee78kEPvNSDR9bJUYoC3vhmP2larrwtwIWlZuoL7i
loxOSpHcEwoFHRvqqIg5v2oYhBLw53v0vg/9eGrpSW1op17245Af56yy/84bn0YS
WR18kcmAsFShzz6KRvUvIZ2MbCbsY2EuWbIAIhtNdPUnJx1EEENInsHS3vTfQWcH
SOoWQ5tbu0YpaQ8193IyDhvNBCi7UMk7lblM2mcRf6cNxjaM2jK26m7ztLSOcoJL
OyU+ozkkQXEYooUf4ptHZSnOJ5habJqSNpa7oKuzjVIx3kgkL5uJYbGu1ybGeckw
V5Ad08JYYW42Pz1RDn3j3ggz/E2NBYHQWhjEHK5EiTBHjfKJpZ8jub18viS6UYNB
qxQoxqqX93TALGY9v/P+a+OsEEuvEDWTlLUe3/s3jvWIBQI3EKzYkw99OkgsAdHR
1BMq2AeIafLP+xXpVJTspkuFcDTQcumatnizGbiprc61xRs7UlfFwlAHZz7PzP+P
kb1I3a2QqOtSvkQzLweiw/WWIFUxg2WxTXt0Jb/1AV6btEB4hAguXJtGXcY86MB4
I4jbeNvM5kPj4n6xIalGg1wdPDU7SEdWHf78nSvLVYSHnTev17OGOU+ENq53jVFe
hiiT1TL4QKZHR7FvZ4d9CbPPE7qSyIq8qV9VBVrZxgbNTC1g68ePKAUDqWqnlEAT
oUQEnQpEcRdehd1gTqk1f5vm6rweVOk2W4AywLWYIcYU7dcTCzF1yaFX1JL+9gcr
fBfLgy/j8TFWQbCbpcKnnPfTzl1aZWAr/QqFNgB2a/rNo1LzRA3mBDvl08wfUl/X
zYlgNYDdqZsYEcdNSdr8uAffh99Gz/7CxkzJMN4WuR3l6Fkz8sgBLS7dxcOp2qe5
1x5taqe5QzIPKE3sIUizmoxQ4IR4E0XAfY+hQbajOVNqxPaeyZFvKlRjUyMcdydf
3BhMvpwU/suDM/lgNypVLAZrosYYSX8zc2hS06Q83DD8P0hbhfSyT0t74implAqn
fxVatvd7nDeg6hCnm5POslQ3husyZnV6BlEpLCMV/VvUTcaXR+HaWmKQj2ODaxMY
xaIk+6pug95KvEEUIZ7jz9jzwl350njdXN3BJDK1ylYlGw9w7OPvLDJ0wHPZ3j58
A+uy+6uuDEcbLQty8Y087/ahn/mxEeB7hC1Xf0opmI1dNN4tvhne51RkXnLQcp7c
lxcC0BY4TqwPqdnTuJyrnUYXfquq1QrFLdAKOwGIUyegApU3qNvqHa2i8BjZQMmz
ZXBT/nIlTv3c3BiLmkeRRT54eoAkc8204PXgSpdl3iinuzHy0zlhRgGOs4fiYoUz
1y7dirFCFoHhn5bYck/EcWOMDYwVKVVrtqB0sYW6L0GC8hIXoHqzh1KZvFW56NAg
YfFFOes2cpo2AB+2EHdojpBvVL/MO88LU+wy+58Axz88fbY9lX+k080lZuX2x+Wy
SauvCHxuGmGZMUjQno+lItRh4ZtRo0tXGHB2EQU4ADOT3AZKJviZKBYRihCTJC/a
vgVrv1U1h+ggisYl8/9+0U3hr1eZ1Z8HlUUKSpeyz+pSZSE1z73hG98sr2WFxZL1
axpt7v/qctjyCFh5Ho+LDnOyESAbR48kFju2xr4NYzSFissuh0BfIaXRDLPQdCeS
MYlb7QUvt8f/2716jRZJUn8LfEnOhaKuSup4tICmwoKOzm1g9NGdurplH3b7C2Vg
fUeumdesnnudiobc4cEn3gFWA6mtpyuACceHjLnwTJj7JnPrX9MD8hAu0Pwh8dud
3U8KSWDG/gAq8hDgpcJUojUuOQMhUto8VbQ2LrrwAYSWZtDe8hfQRjml3wES3MIP
42eaAvI6wuLOyEUlcN8IY4e+EIxuyra/+Mvm+WDWElIYOivv+p54Q0wmps9w2j2K
U3fsEAO91bBhX3v6ugosI5CGEHAHDJ733gmu4qBzbPllTGN/IoaqhsRDRI14wgyS
QUbq+LECTzO7vIl/gMAe5tLaoHKQzkcArF5Zt3n1XOkr0v+rSeFnjLsaYwQCxhjT
AzvI0QjkC2OxDNRJegNv5pkz4hfhlgIuyv6W+WBraZ+M1ZID7pfog7lIXs7P47dn
XP/XkaX/2TOe9T6JDffzOsj7PQT9wKcN901HbC+UMVnJtVUmwP39JB2cYYF/ewml
B9e2QcL6aC35B0VDQjrt3AItCZWixgqpRRInjLFAj2VnRK5uErfXxVZbXb8ycqlP
nDotk/VGEXjfyqVX0KS55swhvhUKXlqlO+7CzUcK88Jf0YKhVOg+xTlfVzQTJWNn
9gNSH7cexkFC4WO912r/6JrfyRNbmItGyVjakQ8x529yVEsF5v+VzQhv8hgTtyAA
HWYQDIqsGWo1c2A5a4WZrmAd7j1hglds/1Fip+0X9ERV1RjYJhaL4m8vHHc90B9k
I3Ic/B4/Qzx49OA02w83MmubQ0mHHwtOYZk1COnWpCQzhFA3QKIiGrWYy+pPnPZY
voS7biMY4g8UHbjsZp4GgRirdA3YsIA1SsjcpZfEmO6hyJxnSehq8Wxq4WXmAKNp
4n8d4ERN0zQk0HjImvpvTsvHh6kxDkmRuS7kB48/kG0QVO0mQuGMVG9hhlhKwR16
s85E+Zv66JHpGYG+EYdKl1oo7PGxzjwml8lOuUc1pn38uZwOc7JnjDisWspquyMh
jhhBRlXbD1ye4Dt05DcBuajb+05RiQsGwiD5IyQyKcCb+a3UEmKmdHo9ZHhcfee7
CX+EwnropwI5O8JMk6ds+7DqUubemtV0FYmDXkzcV/Zon+NYPYuXXTFIjXlvMTMQ
7sjZ3qd0ZRFwUHeqiMFzThNJnB1wkubQoYv38/5TdVy0Ux1cfQX0hj3rhc4uwIQE
sycZl+GQMObKsufEQW9jJWhIcy9UqHeMsK/UQlmpaOFyu7DQv8Qx+dpme4BeIG6X
W/wKscstI2YkNxyLotE9c8QxjEPlSE+r8OAhdE97xI9JciOLo5q/qZXXrcZNYV3j
LSGwYXsrFkVb7pGRkjEBxcijlsS25wbjS4CJlQ1JJx3EHAe+PElCtBzfau+4ndob
ycNsOVinQjS1y4r0D44WKrk6Y4mkOQNQD4O+8Hfb+I3fQjZtbpFx314rAM9tGV6J
DKrJAxkPlgH8i4MKyYGNVpCWG3yrqIUGgfBmu6D3EOuOCJrIDLMKpAKenXFbBuwM
BYdIVr4pgR2h3mMrYNMhp/sEu1vnH9DSGLRCO6eoZpM3RvxT98VnlKyfYWpBjWSs
REbeMJsAdHfHte/r+LNz5sZKUwAcaeplSMtvhkeIhGfPCSUjGdAbIU5XowHwiUZD
o4g4Vvh8MmKyaE5luaRIbDAQUxYntq9RnsBb6ioBdZTrrAz9wH4RClSR9VgVDxff
iaDsVprvOq11IQfaHx3chz776Cz7GEKhlA6bj7jk1ZCqhYDG6K2Kz//QsBLw7fGO
qxQh/V+yZi4GBdRNhqzzdkVo+0OCOwxvvxvscZPI7P6eQC/hJTDyAStfz82c3At3
3h/zPpVO3yroJ7GKLqB+C+YAIUnhMmcJpiHTrn+Ri0IFRbhE/5Uth2mQBeq41E6j
+Ecfi7Gj1bOheXn04tGIYIFcFkyMvYL1Fs4dyhPIoql/MUISrOZTNtMykvl7JDsr
Y66Dif+J755E+GIrQB9LDOjqMs7GbNdUPitXiQjY8zE9qAi5cs/kogZ02LlUh0KG
TruuP4ynb+bUrCcofZ+vPHdLlTtItnJYITfAkG5vOzh0jhga5TIQyvSQ+vnk2vcJ
YXZj0xCBO+8pglFM0FEGY3aOnkaLWprYBirnUV4yTCM3Hh/eWRgAx0gi1ugM7R4k
vQxw+4d/juaVnvnEoIKZk344slRErfd+AiEyfSU/+MBe5YEhQpZjYKMEg26J78Wm
k0ms8IG9GUhCtfWyUIObM+4UMHu5w332YB+8lJjTyEsm4y3klntZDrdNro1hqRLs
jen/8RH+k12hRuOZf3PIMgn8OhJP21Fk5OvQXYV1qG/hGiPzDlHt2JGCTkYv/YrM
E6Yrkvk4sZZJI/tL5kpPA0AEJN+WEHJwuFPl7wa5tmBtMm/qCMjSvYYw9tk9wmMk
dHwFoQvpXk1Mf91mvoGhjn4JW2QUsf8uF6sqZhopRUNZPzUgRiVDPjpWnPtgwcFi
lN02/mckAdbGoIVOxlfmUddKGJIcE+TA/9/U46yV1xvm6Sdd267Szw3XfS6In8yX
AEJlqQSqFl2Jg8TESbiek/oAhpOcU5xh3q6MJIXjMrStJTUBAKuIBiHvutHRRoeP
+PZUiT5pMnYMJLNQp1SbFVyOKQ37yh3DNT+NXCI/wamum+DFMgVV8ON6GZsk8EDD
zyGwYVwxGAGGIxIhX4un0jQLypVuMacCSqJo8KSmFwkaWUsZZVPZNVMfrMqoReW+
7TJ1puPgAwyOWbzblanzNj5Rj4dbt5EWVtbyGX6R+OnZe2a8fQg88k5HzM+XgQlP
FHXLpi6CepZJdxCMwRLu0DEymqKeiZGuEG8OC6DjiJ4/UVTfuUV8/lZBZsVdKpMS
bvirFac90woZsjWGXOrFybCm+Z9H7lXxwMKKPQ+/Yscpp3y5qHt/GMWCKI7ZxuHu
PN7zydOnVceXZ/0i4WAJqWoac08xGWNII9c1lZJ+1wDx72CPd6ZE5E7aVPm/tgLh
9u3CZWF5H8lIp79R2eWuWN256cmee7bh4YvKS6VfG+W9neDX6ctyaancOGAqK8nS
Uc9VApAdjPgZ/Zn6M5YEQS/wcQ/rL7tikK11GiLNQED2ahz8n62JemHMG6f1TN3D
KrbkS7austnya1sg8oZSPyU3m/BlUCI+ffYQPXPlO3M63WyqtvdAOMITg4tnaHIo
Q+y+D49dSESwYxV37TZ+fQWqSDGuMlyy3s4fXxg6P6nSuneaQ82hBbF+5B8XQN25
7OG5wK60KtYzpycs7gSgnNpkHheTEkqa/GnxHoAmlcrJoSgUfdv2ynfg0i3VOAhr
0cCgpAIMnpcIHavxQ+ZghyBckg89nllPcWpTnliq3qwL/1cgEcBZ1nZ/qWbEMRWy
GqJg2GQ2fGMKlal93RA5oS+PLi/vLh1WF+nWRNQk0jWKqHaiJWOyWB4ssx2Pd7gX
YT2ya+NNTv3jLYG8fEUf6EjnuCu6qZOjW8IraVVUiktYWhlI64fqDPHCtMFEPYl9
un95nzjrsMtan+GkgJgGpCSDrsq5hr2iMrB+7raSauEQow1CubES4fBBhtzTdDvf
R1Xnj6GbdtNVviG72XBIxCnEDFE9e+ADtLVGkbpqnNCYX+YamgzMQjoINTeEAqF4
iXAGbo7rZBSdmYuBh5VsejCv5dkjIKfADBM1N+7HEZ7h3G8S+oTUZHci3E6DBaEb
xUWyNJrRcl6vyR9V4dzKG8JlHCUYvhbPrNt1JDRWob9+tx8zAUqfeoMzpHBRFVxt
/ibpYkRthntZ4o71gAH7Ayi2IGvxKP+IGQkapbApAuOckNTrhlt7VQ06ZRuhS/NF
3PY0Dt37g+1tkSLDCAbR5xhc1dvF5h0pjqcVcWVoS36BtT+0ILERlsVHb6rYjPsV
7GjpY60mX2pByrdSxfDsIKQiVMKt12FqZ+tzHxV4hBdV3w054QsAgqlajPxPKT2/
fEY6AY4aP4rTxopHFk8j9uzWTopxA02x/0mIZdRSGIgwe0iUqrRcK03C5k7UrD5m
bEBGtO9m6mxpGTDbr+1UMJhcQLkATDHM5rjeM5l9M4nIFNrsmxD1nY5BObPrSwll
lsSb1nhPQ3vhaiEYDLrdxPUJTCZQcHdolL580DYxDHW6IsSIxrgjMxk6ROlYKGKP
gdkDOSRH4q3VXIPH+H5mkf26yUAKmWvCnhDYmzh2Xd0SKSPf38+oavkhf8nELevv
dj9FbcpttEUTfak29ME/7YUTym2P6GXpJdrlr8KjCU52qsuS02tweKe9jcrnarji
gGX4oCdZJUiOfCL+c2o0rrNmm8OlbHO6skW4rAsWlk9NGRMkqvBuVb0jrDK2/BV1
xRMrdNG/ZIO1/9XhVULLjxoEUT4q2AJbqZjASxED52RnzTHtAqlrTE19jSYaO6fP
VKk0aH4WomoH0UpGd1FF+qsP1f2X5XBB82ltdg0dekXh7tzI3fNkkT2ZykID8L2U
eOFYoiFg2N5j5785nFHsvixXMI+W19MaL4LeG7yuhhTBjDsa7xn4XXBEGzMqMsXz
J3NdZKtgOfpZXE6YcA1j4OqC/xHI1s5IruYtWrfr5miRfEJSzUXJoFM2gk+Yg5+Q
2DRA5BDfy+zvG4CAfvQcd498OgHczx0t/RZH2DOpQFVhIKtIrQuOGNFXVuBkh7pv
pqTSbttUV8J8oNnwC6U+RfvKyd66iFKE2v8V0uVmlOQxNTr5fYF4JLYpzO8I++X0
3Fz1/h4Bb+wCilqpHTMpmCHU4m6M0YHXKf3BkLp02fCewKiHWNFGpmbRLh/D0X3X
RyFHQt0mODqe2M8UBEsItTmHvPobX9N/hK+kDL5iskC/AxoCGmZfh9+AhXZtiiPS
cQ/rye1EwhStZbaGyZQYxvcCqOAapiSBMAHDI5cMIQpBtmuCD/zZZdD/gyANmDgB
2ftsJTMKOMIgeimY8zDJ79l0Fiv6PcTaoZFSuoetL7rrM5o4yZ8bwTCvgZJlBH13
PSflTu9JbQXnBeSZXYQFO59dvgcnbnDWHsKEhSar+mm4av5M5qjKnFsTqzcDy+mn
8o+/kBwb3iizX6eh2AEv1jKhzg12yvWp93VBEX+wHGpjcn6ShkHCFmPsK9+fOvfw
09RMkSRBvFB5MZPKGs8xMbUhJK72CrdLTkSmHe5369ehQuwRU+f8BEkOiaUXY5jH
02EXJXfwlhubZr6ExT4h88ehzj49PPwC37Xr2eFYlucsDsal7wG5xyoOaH/xUEWt
sQ24/EoUIMWr7P8dmOlknD3vaEff83SqA4WZ0qjw7PCBjt+LXMwmqVkRSEiptYR4
CKU4KjEs9IH+QTAPg1PCu9H6dwH5WM31pia6mFcOZ5cDxY4A9bo+fSgpvknUyCoa
aUwmOJDuGLiWGeLGxvuCab+vCq5GqWUIfa3Gzom2IrGLhmFvFsk6OK9YMgeex7/V
gnjJVnm5l2TemSm3qHXtFzY1AuUTspDE81PVofJ4mUjFdcwQxrVUhf8ttRu8MRjz
Koeys59vy0/e0hM+xi5tXT5ZNz/e6p3BFFbOWv3vlFdZbeF1c0WBCMSlbsXjIR5m
cgp1jDhv6V0cROd4npEQuIaCins1OvRbAAtRaLI1slsQXfMF8Z4K+S355dpQ2c9H
7DqGkt1bnPa2kSOZ7CMDUSLtwC4313UuMNQyic17tsyeMPrDjZvFh+Ah5PTVWRkE
BsRiMznAocXVF0aQwix0/3959xJB1z4P5Gp7FMY/Bd6sKlQV0f/Cfx67qxR9mstM
z32QbDIi3UqISgG1Aglrc2HFGJYOXAlwl3IEVzyIyXz/7N2ujO71JVjzWBTsQ2aA
IuC3oHy4lLXcgdQBoWfXq/H2zkYjAOxc8KhHU5qgGBbwqksogihHhAleCaLBQwkB
w0vYDp6XhqFjpWh2t8Pn7VJLPeLu8gExB9NF0eUF9DRDi7QvXedYgtmmyuvk/bf0
yxPvIfpYL7UWILgmOKzHgr42yj0032qWox5zL+Yp7lmLAzHWYuVZDvnpd5lcCmWB
tqmBOj2GCRmX+MxBNcjT0+s7XRzvTKtMELIV2adrWHP3DGJ0dSUrqTijOPA021FR
fP5iU+kI6qIl83PlYZQtqLaBTbWPAUBiODqzy87832lmQ0lrzehx1ChsKJSOS3Ow
BxDVaW6KvaUSDHOG01iXh0cIls/xplE46mGt6DQBkWiD1JESWRnSmwcncpjHi6cE
a6I2Muf33ZBJPLQD+BrX5EcDvRio9s5yQ8YPUd0b9Q4r1doB6JIQwLX9ohwEAZ4Y
TiVCvMIzu5DXnhQkuYw/0VM3Y0eobcKn+Z1CaBmmI9gW38myG7cnQX/tMHTM1wav
SPg3n56Puyvz6EagIcySZi0UEIQUFGt17VqrNuLBedFNToVwDwROOwUtGPh3Q/Ef
n1O8KjFb5DMFbi599zRGflAkcBGoB8ZWQi2SYZOQXcJovyxPMWa9HFBgokpN1UjB
iM3qDV0dJytqhoAk5lZB6MShZBpO7DzX30o/PD/+lUb0pzsOscAx/CePPBKyw1yL
GMdZG9lVLJ9H9BF+9AoJ4HPLP80M0CVnk2DNu0kvj6DTFbJWMjvg5afl3S8Qbf7Y
RgWZeN4ZwJwNvvJAwvF3VoX5Y2LgE5vqkK2EHxAe+GoTXozNh1kY/Oi8WiH2SphK
Qv0JlcsialoW9D+JriLyGpiHwuEK+psIdSNU/HxxY4MRuU9jvBog8jGSbWtT+l0c
KRfEwuzsgUHU/L92+zSr+HGygDwefOuVNYGncbmRlvUOSvjZk3msC5GLuxsysHB2
LfjGwuIrqm+T4sTIT/iGHyjKaHom8z/D5Qt9Ak6Jx5XBxNseFlNmdBrbmqF8irtn
K6fwzwGzxLtEpolUeoLOd9tUV5n+McjBjCongSd89kqiVLTGL8OvTBAE2vSa7lBe
CoYGkMBc2khVq3vVaWlCULN/OTPuyTOsDap9IiJYHXFnPLOAgAQ5Ik5rbGtEiY5Q
0GNlU2SSVP4JRkU3tQhCcVXRoqsFjxUdnf2uAvUNuOn7rXXLozEN0zBYKk9XrfBN
1oW80xR6JZpWP3C7m3r1yxGar/z1jzPvSo6DjgRLQH8/n42slL4vh02FRdbXBLzS
L3s2ew9BFcaPsKpdmOmmxoTnYNht99TmHVlpndTw4ElEVffKcvywA5Tc4l37tZ3K
hpu1JZUQ/EnCk8GJHTIvs5zKPph6KTf54KAQ2jXrf2figdV+JVAOV6PIFcIdPpT0
ffutuXbTB6nsdf8OmskeTuYdoREewVR4spZLz1H04lqxRkPsGB670AeQ77TsuWrw
vAhYIjEd/oUjF3KOpvo6v8R9FcX5BeEo/7bxgXX3WPOKnUZ670SBKUpFc/Q1jhhV
/G+RMKHaT3/2h2TazB7hLmP6ZFfiwuSfrXtF2pQSGv0jNYlvrCB8vmB0WIfwRh3d
XjWcvIY2BOgZzrZycFH+yDr9Mvs2hnCXX9KF+6ESZCvrxYYICq/YJyoI/xbYzwmo
cW72oa9wAIZWphqGE0XP0cVU8xVjgBpXCt7T+3GaERZnPR7x6zIxMaGD8RZANve3
3C6mXob//zUjk4SjYZm5h9VEgE0L3caG5UHsBXVW9CN2J7pydo9oTR3Ef0ssV3EV
GG5BgEQfHlAweS8+4DKQQJ6AIq9DNO4TJ5o/QdkinTNXvLE252E+Yci8kBKEkqwo
+ToZMe5dE1Zk7iYW/29mnOvbBJQVOCMOAn9HILZvTB00KRXxBT17deb1CdOro/eJ
AFcq6mCUY/0EqttlcCjgeE49ttdWBRXgZ59+IWlFGUL73h0gIvphJe9gH/RwuT8a
kBl7Plv0FsEnMmqvW9Fa3m3Y7aQVXBuC3hKjQCoYgfPHTmYdl38wqrpgYAv3vlig
d0apMsUGGvrVAqBP8XZcFcpzqLfesPnUUZeao15qxSuAXHDAAXf+OtfxyB7mUJyh
+WOOQ/Z9r8ZrHGaeLzy7ITQhO7KRzgfKD6yBwyUqk+duUm+7UY/MeS+84KXId1hR
UVs5nqandxFCbWIBihMeqXKKwz45qYvKVMQzA6w6ITHGiD3lyQDZKNafEDzmXctP
4T7vCiUSMrSFZQs3k8Y04hfS7dho5Y83ElXQ2J3L0BovfMaVBK/xkzZmFBGJ+Rqa
wJQ50+sRzBEtj9axVftk2KzmROOhyPwr13lobHsE/nMOSYlCrE3ya3VzeAIvjESq
os+IyzKlUH68Wsf8D3nEurOyno15JJw8IjWu2SdDUr7nR0O1MNXAM8iayt4K0/vp
JF9ZMCrj65vQVej/uZCBMcqazj++mn33TaLAHSYu46LVh9+DWmchbmPPCdbTmgHH
yWQMM/UO2oP4Mzbt4a6iW0fWGC7GUMhFO0zJ2Ep7JpuGKe4hiCtmDvZshpV7f67Y
fVYIp5zLFtjDinysrORaOi7L8WLdsY2vf0MrtPiBx5s1Szd0FgwcWAtFwf2DgXTJ
Eex18qwSRV/SUbzuv7VAwfw34wQG13dYLgtTpGVp/yXYTkKOWY+PWidSmGjBCHVd
Sy7O1k7YX+wkEZAazMCkVCWYwLayMwXhJpf9Hx9DELyF8LdXCKptdoV1iYRTZqtr
IkzAHaqkXfW8zC0JeOe3yCwVc68XLjH93BDwZSRSjEBwMGLhtuCE/B//GYaYrBO7
++s5f1oUH/N3dOSj8RUHXMImmmss8Q6+v4SmJcdayUDhH6uFu8hYUN+iYVXcz0P3
nMKnpehPkNmjWpR+Ibhsqd6mEegohBAvzeTQl3XyJrukZQQsMnh7KV9Omk1pR9FA
y0PAJ+xMG9idxtyoI5M0PMoxAlAc7d0+F8KRI36kjyxcrOe1A1r7znWoy3Yr/F2f
wLDtXmwKK4n6NGzZbRK3U+wEHLjMMfbnN/QHtuw+B5TJ33ZICEa1RmnOBmSdoY5w
LxHaeul9yUwbg0FfPwOzgrwNkxRW4An5qsb9wT6FuD6i2D1OCR6LY/aBsXtky0ci
CrjchDZWm0DjhnYSl8dns8odTbImS4K3ArvjtDj74asQCY8QN+zwnA6CcKvzNtDW
qeP+g/SFGxwdEmKuiDwmYL0Ahxucss/2DFq7jESYR1pKiqWVVXso7wqi/LRAoY2y
YTrQeb6umfUv/xbhUVjiOuhwpB8kJgwOgAj6ceYmOp3Tjz3q1RQjgfYisdt4ZTom
AOatcSFhwIOLB0XLpobFd05n/xzKSuu0vko/45a7sR7uATJGUBswD6hZmEYJfz6q
9b7F/lEBzpDJTJvG2aN2gZxs9U7DS0ooI7DV7NtF5ARp2+nTwAPyKg5BGKTwaLtk
1eUeh/+ab8FHxdmOW89T9vbpGQB9d1YLp/2rhW/lbowV1zKKP0H0uMQZRLIMCyNX
hNpv5zSyVxkMFIjmgQWsNqy0EELFqunD8gk/c/QjYntEeKS18KyJo59/Bu/hMBg/
9rLModaPmNZBEk75wsBwwByeGxxnjNYVYyc42t6h1cAtiEfbda+kA1o/gYrnJdZJ
MouLETHdYXFEGOJF5DwCsn5ui/EKdiE7Of16sl9jJkMm2cE5DgjZSvY4H/RET/+J
lkfTYs+dhGwf6IRKTjWLgeq0PUB0WNOo7hOcCXJqTrzNjXeXYr/CvKcmBHPlXay2
bCwgiOPZ8fdbNROL6vd7VlzJ1Hnvp+XDvScvxUwJrFy6VyYOKv9aAxEtw853qowK
MJ6e31GRr+H5GtWbHcddcPkuLglUQjO+v7MXSLz0TW2y3xW7yoeYEKlO3SFRJbOV
sOqftC0SjYJQlIQvv+pB3XssSDgzcV6kt/EXL3nziNS02A084t0jZIGaq1iL/42U
ABaJ1s1EdXqVCm7RE8AYyRhsl5UivUDdbd9ZAey5nS2XTug6e8s7k7oHDrf08CEx
68HGabpb/AqXgnLZsMf8UJa8/N4T4SZqtu6350KlsSj7gvW+/FqaohP4qmIbbn0g
uE4VnJDXj3N3W5OKjkZ4lckmGPU2FJHlcs8FKbNFlWwnXh8tjoUoFxn9U4dYTjhb
xFyRpHYS3Bm5i9XaAs6swYL6fJM71HC9JvCKsTGO3N5z/LbHpvn0hLI3NDxLS9eR
FKNxeSnW0RsR9meEgovLOlRqGai8bU0qak5l+zLmwYDLEZ8O/g3onq14XP8Bz+DP
Mr0T2YnhP2T7AzNJbb2DeTIqnThDJt6/7Bu5oWbKf3CY/3qJUr/hDQl8BlbTq3//
p01/Bnb0OB+lpYkiSnoDfCgJT2vi9zp/ynS/4zjo3C1C4DOdzG3SYZRmUjPWyZKd
d+uQB5bWA+uPWo4h7zPHUgNPfoLyB/pmQz9QvijJvN9Q3j7jk04y7PoOIHrLHMLK
AlEQgnzkLk7qLq/F/W0KF+4EkcOI5qni72/vKprSMTjcPSS4vdCoCwZZHEFScUWK
8rqc7l4z37GrGLftPDh0FhszzAoBD5rm+lzAuyCLg2Xi8dDcVqYYg5mbGp3VJ9Uu
AOKNDj01adZkvN4z+rF4Uan/aNdUFZ1nE70H6C9fEi9uXpaA6NtR1j5JbM1cr7Sf
EQzMbpf4MR5Ym+O9MdyOpvoTb034QTvcCVbZsCVizr0nmB+QCPf051ftGAUCYIjb
sZwT5kH2ipftV6GShC7Nd0aECe/J6h9c8dYG5R5NC7qqHvqbQPhOBHUOtKBF1KdE
fk/z+9ykFSgzbeQdAWKpEzJkLbwLhZdyMTHp0ZnGb9vMf2RttwWffRw+m+Fpg1zF
YITTnamuJC6GlxZ2YiK85pH+3Mz5TRJ0WD7COawlRwoi6s7pdhbA2Wq6Vm8vCKdR
0TBiBzVmdid6N+5tm3MhhIFH6R3gYv7fJi8yinVtDOF/z+yf1cZKT8tOpF1TJObr
ZAHWyeOYln0f+2mHbxllIdoKJVfQVjJRNBn38jU+Y7lmtPYnlRmLfFnH0AOrj5Wx
HDf7JxvloEDkUPmqoYxhlJ1oCGjLpuWkZcmeSrwLOScTEPd8E6i9jeYnEdB+x9er
Dj2JmcOi54QXqyAjgx6wUf9hJyWVSdXD95kDtXvPGpPm1cavqZJ9vJ1QOPPRgFs5
GgZYQsWpnyJNGBcMTMv41+pMSG8KA8x+d2DJMkUXSXfkmmWK+nCf9P/m507JU374
MYTRfNNgO43gKd3epRSDZfjX7risOSckgRewgR5EEfxRp6J/+367qf8XvZ5hSoTu
F3Sf6IrW7LUaYz+VS8kiWvyi6K4dC1byYTSSkQAdYmOb/X2pgYWl1pa+eD3K69Qh
WraiwktsR1rgux7bBvRSwAt5RCTRQ0MMn7+YyLp8gdWbQWOJWxKLJbzwitJuBSV/
41Lrmh/qxXtQ9Mrl8PYMT4vM6SuGwIBrpMsTeVraPGJ8xX+ZbtvJa6ZQTdwYSVwT
jNlSnsdrxWYVVFy0jy5GzHnqqZAdKDZpkhBPcov7Mwqq5coRM0eOMZxdaxSSophj
pIba5ASiHmfCqV0EVPazb5c0Aw8Lb8RqIYLmA/KHfZFPXjdmgmHNmSirZNMCI611
0sUhQDC1GvN+1T6ibKfi0JNnZ0ECpIMevACjpDnO9v/kfB4eX+n9HYlVTKl+nYR7
/a8+uS5meE4JDY2EVr7f+VE3Ht4yzw2V7fzXwsMQYTJ7O28A00T5DR9HFYGa6aAM
q3a/Y2MbeK53Mww5cXLPc5hj/ZHDYZ0m+oty1LTJcs/UPKM014uF3mzgt9gJHTbx
i4/zhrbawgV6eFW4XjNutjUQbDZf/Df78W1fiC0iPR08Erg4VLQic750zPGvr+3G
vNEe784ORltLW2iTn5ULx8JgvbX0OGthpfRef7HlSCCc1GadES3OdWYa/wv1LUQH
kejuetWhU1ITmK8BXVHijYEHrEwyiOe6M07uiB3E4ba3DVehs8g+gTE2ktMfK65/
sZurG7B/xLyZ9/mjXO+FuwIc8b6E+SNfTf0Qo6Lx1awaXjDUm5gZNmtc7kekTGvp
H/86uwPKgphxjSu9znY14u9Lw/J79IczvzhL26nPeLJTxuR7b1ccmkHyvJesfHf0
LNYwBNS4FAiKrS4p+aTgJyKQpdqPWRjcqK2Tijf3EDoaIs/9K62hoU66qTefphBH
TNW8uW8ceBzetyT7jBBlLUMwFUQb6JXC6FgziQhmoyYkm9uFF4cnqwp6OCEtoTcn
Sig5GgqEhKcgwipHTm2tUcu7ZiwV0XpBJr/4tMn7BZUAdwUpgkeMYT+NKEeHs4ca
fPW7dAKRg4NPzpY3RHkG1yIf0SZjEkxTUYh8IUfvPI/EJLMdM1xWYnKO0bxXfciO
+L3jOMmjkql/bFpa3hpd0uhXQzwTY1GlHZuNhlciwcMB8TVz8vPYhcZq1f5fRwKJ
8ZY8n2JOgC/ScrRPZxFyfoXwUrXpKV0eNerDbfd7gdJALlGgWYnhVa9K8Cd2K2YY
sx7SVS4Iq5cfzWwNMilvAW5pSwOpoLaZ9WBXhlYgoI8cCIFL6ZUBLHe3WLPLVUD0
Gvvsnqoym51i/jforb7KRKdi7yNPD9L8c6EcobOu6lyCUMJVp2ZiMpdspdYUEEtN
bmnZ5aooBa+i8TzPw8GAAaOW9KRsHWSRNdGbvkewRHjlharLCZ2P1Dr6oQd1N+5C
k1fTRk8C+2wmwq5yxi6nPc4AvP+Uc7wX1z0xrWOYCpez4TDWhMofYtiOiZjnc0bP
SDQod3EodUfZNsUZ3cZcQ85G9NeHQcqTE/ix1okt+U9im0gndWWsNAeKlBPLh7hD
QvfOmTw7x3H0f063VDjPamIHzZvPyhbFWyG/Kz5yRe8CH6IFN0ftgvP3sGFEz3BV
A8R9UjqaJZg/WRgwMDwHdcj7Yym3YQHA4w8wIY5H0Y0bh4uQr5rHwAdy6QWCOB5H
+SFal9IrG4Hbrm12JA3JCfQ/3w0SeDvmyjcVsuCdO8KLMZSltXC580fXTf5K7Pqm
2IHnq1tIIkJ+zKFrPLko7+4sQlFkUrRTOcPK/j2DCyT1L5swjzAFC2csD5bifFU8
inkst09h7/C4VAYmpynAUq+u1xl1LWwGxu5JNXwMde3iZqpKGsNQVE8bamqFLM55
VEJDAs3CIEB0GrdrxFrvwSSi7I1StdsiAVsglJycTkqQ1tnZYaSOCmo09DgCJPbD
2zsRP6ym19F5TIbkRyNFusauG0XpT4zkMHUvoOtPFrwHqBbaHS91z3C+YhOO+EPZ
CMPhbwA3d0dyTY5ZYkqkMc/E2908tF9Xz1AqKBKswqyw5jJJSZvdUdo/yAy7pJDC
Eq6IMRG8cP/YB5DV/MuaQLF7spVbaaINy0ypADbAI8OMQ0/603ABDEVsXIALzhej
D0zxsDnsuX8ZPEZWgV9PEsJ3iIppC4DYcTKEY7uhw3gKyTvCXPwPj9/AJErVBvNq
m0J5L+yJ9l7eljvXBtpGwJwhZDGxFeJPbCZ91TvIZ3rpz/yRwK1dZumv9mUG15fn
sOPycTY3kjhVpDhz5QoyzY61/HfgCnvukopU2GZimrWAZk+CbYBYGa/9ryBhtmzl
zkqVERibONcLs8tiszEEKL/zbTmhPORO+m3XBGUCb2rvMUg6x/5JMXq6cyh6+0Jc
qT9sIJJENMIYg2wfl1CT3VsJ1SJgtTabG1SuSONKb8HU8EvwgGozeNvhQ41Yc49s
IrLUIPLg0xEF3UHwgvvLhnQIi6EzZgBEKH+ejUGPpMxpwLBmjf6p4qKIwRTMuSAb
EiTm83WpXf1TYs3VrK3JZh7zALohYEyxKmTUsDLaN3mqFr/hP2dBGeFWw+nxq58q
FNjZf5RBihaHmpWCctrgU5BM6gptbKPjZVt/CB/TqO8nZ59mNpkEjeQvDEokIAHt
dlTyFtgK74FUfr6RY+659CNPEJ0F5UzeG6MMmm+p6cQDfOwnWdhQMn8ercDJDK/o
ILDx0xvkVW9IafJ+DJMBp9jM7tVjVKVnyMmfqssDV7hq+JSOYOG+Vlsw3f0mOLyG
C20oWlR1YvSpIPytWBDI8HWMxBfB3/sk9oMHoKwLg46Qk7ZrHSZuPTVgcs5E57jL
QCIBI+nmEbn5g1KQUZCe31Rcu9UVjF1v3kJHQJCkedlo81w3gVtQcPeFIJsjZgfk
cM1BAXy3Ki3PeC3Ok7GLWjmhiDkVfll7CmrgMJadpNdrhSbAUzv/05zH17hudgTV
ucLyGMQha3XCejBwpF+LH0W18zg8CB6PwZWwWMj65MCw2C81WcatwQ0gvyvpwgdb
iI11hJ/TGSE1N38nMHMdwwM/CZeGCtNTgueScZcDB0mM8SgstOkUJ24z2ulisALR
WqyFV7AxG9FDsnB0OLKhiNiSsB7XaFw6IXdud2H3w/zTZx1uhyaZuoLHTRZuYPm0
w3GcRlMpfEcb1ogjeyAGHxVEJZszjUkUgssufyi0Swb9dK+mJrkW+Km3MTKREBce
hzS8loFarUnwrpr9yLIruRcId1DxcVKhfUeDDGbC1L+ta09DRIw5KrhHw5vDHlxH
OIERJ1tSegRsWL3R6pYJNlf/i3sxIBRtiutCChEdKgWFRl3pFyE78yr3E9E/Qxtr
nXbvumTzRdG8/Lh6CEwlmGpCgAjSFt2mp0n1KoXFnxeGDpAhb37CDZiSbeAVJQsS
gi6PdmweQK1THIenoTtChK+gX61o0ZJuKoku2N7Plf2mJHEkRNrqVACktDyXnyFv
H7qJSsD9KgCUKZ3JGQkXrPgtyZ+e7pXTDlWnM+MrBUM5ieXQqMXMrRVd9RoDYH6Y
cTYJURQAfpEPUeAdN+iT3ZK+vvEjGkoNYj8P7dIPXXXZSzQep83I3KV0Il08zQwD
Tl2ljKVJTOaWEJBPSutvCY7roHkRzv0WSHb1hfE0+GmWA17uUcgi+G/PffJCl35v
GDupUXMp1LUjUuXL6WEymSb9cU/HwYBxIwKooDf1I/3ezlSm5+DqZJcuQeYYbuwN
XCuItpKpx2bjWHHLT60qF3grUuuDi7kIQ9APyv+jPUjA9wexyTwqanRD4xsjlwed
2Iu9PQF+DL8Au4+T3VqpXS6fK+0sQkxmiRDZYZIwfehgBq23krTfk+Wnh6ahmzY5
H8jm/tAYf+WU5ez5n5azUwVz3HZa9AAs0FHgRwE4Hcffz3T+cdHmFMF6vQBAD/Nm
c2rH7U6GUri6cEej6RQh7usu7rwjH7KdAv3oq7p1FkyBMNr8xk9TwH1QhiEvJf+G
UdmnMh6je9i58fSU9dTe1DNBg3gxynncTiIWETzWxgUG3B6w1vphpd3b8d4HvmRZ
GHusnPlrtNy+A4xFoQO0yM9qKf9WlS8dPRaI5a+uzV7FDKZQ5Ek99oeFIInA6vtK
REjxxWISLxzaG41SGojlEZYNNtDulNSThs7DHzvyTRFPwF2yqBjvSXQYIn0MKIWW
1jVcGcNO5i+hH/ch75fuiX+LWyftJYijnkXr8FODlb2FUgec3Aphlz46VW+XqDw+
1teCX6kXKx0Q+dRLeRMMNRsRfruhALUKq3k9Q/IHotazqoJdzvhes3e1fec5sTan
/4lS1QAc5vbcjhHYFaBcxz9VNu5qwDTVwTUyq8zJ1b+1fYnpKDnmOPU0/zIVg5ts
3bQt+pGJe+mQgMhtJwHQMoYwqjo8hXqqQgdsi/cQ/f/p1jGaT/jfP/9Q6akcZ62q
uneHvmQGDYFVBL5luzA1Ma6VxNQPknl3t73E4rwFTuBkgsiAS0zji6SACdDPlff8
WkQSKiVGLussMbUAPwLryh/SaXVvjyUufLdd1RCfPFL+Xy0s59EvxfcslNU8vHWC
2K15EeD23Aj8LAXkG1EcBDdXkrFOLe3zkSzQYfWZFa3EKiFz4EA+coFqNdWpO3Qw
DBe4oh49hudHj7ON1dSIQVApzo9mJe4r0BmAShhr2I0dizs5LffbEeHDbxFKN28x
uY/NpKJFJTybnMiP35HBoBB96Bmd340ztN9YAwY86mnhs7XNB5u2oxxNDShu8j63
2h5YcQa8g9aAJkYIhbwtENr65n7dRdcLWYIw8sva1xtr/AKOuV+n18LnAQnq17ux
t6Un5go77s4u68TRQrGlS81k5AJTsQsPorVm5jFC2WhLUijVkuVYeg2NuHCjIdu+
u5I7NQ4OwBEyUa28HIvqqGmmGP6tpg7TC1ywlu4rGnxWKcuL3hCVt8Qpl/RBs9FZ
dv5/iUiwhdhPfXD3/H4yhO+6Ftr6nzrgqm2Y2Zskvzpu7qqtcSpeYSkXyjJjQaGR
FozC3wVKub1PWkkUkUPODMNHM5oxxtCcRmAuplgyevcU/+L1/UStEirDtayY2ibo
nmyH+fmOH8gg5Ib8bAVeJsMM9BvyxIfeYr9uyGFdOrEBTy/JujaO+swiKbtAoGU/
1v9R+/+KWBkAidrH6C8k4sECs/2J5kKKh/mcp5HhrIyQzRR2jBWFBUa/enTFxvkY
4wSz/ChQTfRqe/bk83jNGYl4nlwgSOlQOxFbgj0JT7/pktF442ZPvotwi7cD1KSg
Rr45i6sRyj7XsoZXi1hrEgBrABJA/5IktRb7ZfkrA9pM0RSrGUolqYAY4ZXKMzvp
6div6QdlSutIjDGkAKZuuiQZTQbElBlpETbdieCU5blDSRbfwNpPCfjKd0HDb/Hj
xOMeRW40zOzq44Qb80IFDy2DCV4HuFL0wvGUMkEGL2kwdRAwRYqgApEjKis3oGH1
LHOSZ95e8jVBjY2cpRSczF+IH0mT1+RegTUbA3rG7PkTDLCLEkU1RFqVp+9lqdD1
vDNR2Z5Yq8omu2pbb6Xvky1KxT8thxgMn1e/wI53EbbAIFv9ebnIdcpdi1+LNiIh
8dNs4qeOh7wHpvFoBZeS12OEkLOG0mq558nKI/DvakdD09kZw1ZQRFn6eAbushwN
0sBF4wpu/XV/nn0XiAQip7FQ8e2w8dYH9Fm9l8HCH/cfAxoJuAFE71o1TzBgZ8/6
KBquTBnl0JnqX6MgHK/sxxadwpRIKcYvTaCtKU6cQ34An1dtBKfqy4w5jDox0ZgO
R6Y5lPG9xcyRny17O7K21RPZ1hqcasonXgw3EWmae5Yb0Cw/EwYCF1E9ITOEee0M
jtPPGT7/SKxMmUIpABxClKO8gHsEgYsC94HnM7bhjuIP+KWwYFkScZ34/8oAO9Vq
cppMjc7h+SRzIfZ91kAecrx6DkNpbY79PBvsAJHE+fVl+9dC4AJq7m3ECA1MNJ1Z
xFSTSgKRdqZGUHLvi2LckDO6O+oxrROJ1qnU55keTwOOk8xwWPSEXLu9dQqKwwpv
TTXNotl0x9ifjttNgY0/NA8uLHD+6Yz4diwi1ADu40Z4V9gvqTLY4ucgkVYj2PfB
FEQzSB2wzpUZSn9yOhQ4u3Es2mqgr5b2HZAbKgi6fMLbNkWYEiF9pzXmWJGiskVn
QlKNQCiDjGQBZ7ZumTLTJ1hnraOrmLwS47v2eTOyzhqhGszdTFTfgCElk5MEXVlX
JXGvGViNYlVG5R+xGWbmIQFfwvvaAXhOS6pQedB7EQQ3zvQWkk/gk2rnEEU2czS3
DzL7TRUjHHGF8NYR/U6DzWlIQEXzySkYaNwhcYl0BUOXY7dSgwGlmA6rQJyPrpYm
2uBjxLCyluhJY66oTo5zX3nra2UB+relmVVYD8Px9COBa18mTGBNhVwqDb9EZZEn
1BDGlDBcY7ycnMB//h/++khDgmIt6PLmJLYjd3qGL4FYCnny/T0GK7dJeyUMYxRV
1kBQswuqCBNiPWUjCJRYM0Gw2Xz4fTQfTff6HphvgeKt9hwAdYlnLe6y2pDLlvSx
UYyVf/gAsBRZiTwVpq05k/bZJVSPcmM9cA8J304N8A0DZrOwRqdzUG1El1JUzIyY
HDF/bpT9AxVzIQ1ouL7+v2xUykfBnkVGY0hbHcaFdAdofQTCt2H7qaPhQOf+3All
T+/zOIw6baXJMwUC1Zw0DDVDcxHa3YRyLOL5oiT/L/8KGN69XnB0Vi59sVmPueJP
mVHh0bnkloiKDqdDe/8BxOfPR5+b5fCwnb+4KXlPW4u+KhWVu73KjDzbS2Yb3wM5
G2MQpKj1WWKicNzFJbhfCnNqRHNmpFwpfqrIJyJX0EyBssAyIKIjUUEr3AA8ApZI
CLhMpxZdQrxk11s8pek6Lc52XexAw/y2Avca7kyQSRRc0fPiLiPQIZwPLgKZtTj9
rpXwW7z7apb+BDvfGFI5Ns2CAzvFZRbuYkxD8K/NToQ2L2FI1SFdZZvvkuvXrlua
lUs3iQbwITpAL6jdtPpjrmqo6M4OC7hLxQHVT6kB7jI0qWGNMOKSI+JlKUAw7ES/
+QzuNC1nDBAuK4t/gpxQRZTmzeEfgZ7wMdfaXqJi2Q+FgN0Ga4+KmpTcfQTyHpg1
rSRlZ8U4Dbld67TJjuyqGtHSpxoood4OKmqgcQkylEHzPgf/H2PdiCT665560c5b
hKXR4gxMYFgZXbDAUO06lddp2K2Km9ZkxGvPBWEMlyblPTH5RDRcm4Szlf/V+zD7
AHW7H4JIHWD5clxONfyjXT2qsb8ajEvA3Hho8/HY9NIRD9BEJNw2rzGeGcDX8l01
H1uP4zKeV2x9yqeXW+lr44lX0UcrRZuQTE8t6Xxlhz7+g3EDzm4pcrtrWoqdWu9r
nntDDlO+nWIBQ3SGokIN//CVOorDD5bJR3eZvyeyCZ/KgHQvSULfEIeFudIqycDj
EJAODuTv8OJO4Z2SuXx4ZiXVfMO8lPp/KQUayTS5TfvMqJqXxzAX6+UoFMZ+aLr4
zm4PMX47PypC8BTX2y0TSucgqhzahj7axRdTNzr8oQUn4HW8HKRoCZhlvEKKgn2R
mI9VHBpcH8EIbFHU9WFzfOZumtp4MVS2S46iogwxqSCgq8aft5Djfhl1leZLyP/v
k20/qgV1XMHCg/pa13DK3FLY95M3kSLVw7QOUb5V07dRdjZpS77euO2FLH8JuSLx
L04BaqYBbZBS+L8lzPcwQ9CbUgEccyenIEW2RpFS58L9XzpSzg3wPy/1cXMpxIBX
7+KBkJthZbevhh4sQkMjSBfG0OGMjBhYZ/fqV6y+71f4qBcmX3pVHjvuZI5j9LID
AVNLs4ZSf7u9chBtHnALcfuYZiVT52Z9PCZlIubOzm0blV/9QWzys843VG0zyujY
GQB5pEb+fxD5MdHVo/X1/w8lyEu2pV6R25omw6uU23EBBUf+2Y3mWeyf2OEhcz23
rHrG8yv/mjU0hRpw8iC4/ZAw4IhZpsntgHfyjceIvjBaZOAcxA591kRMamTC8S6J
E15FVYP8HIsJ6D8ga1qqUM+qlf+xXaziK5M/i5i9dOxdNLYgpN3VnThvgXVBUmZ5
Qi8bzHoVjVV1y5QS32LznB2g4oTjjwxTlkXpTbmJmIetSwrRg86yLddrlmiyba90
U2Kvid0jcdov6Z8Rv2bDCMoG2Ck9kBqdSCQJBuu/yBVjqXyGGnPp59JhyFVmiYkB
Hc2lve2ETIyjbBXFQqJ945PgLidRkjnnCnsIY50/aSxTcPaHfhtpOGntqd3WwaYb
kMxlC73dnpKBaJ+oYrkJ4zLaga7nD5d0SoShnoEE1dpOu9eRSeC0O+d8tS1UPhRx
xFIgz/77XP3r4M+A4pgdnygCRXEe8Dkx/h5ughhW3GWmC+PmLpeGzN0bZnn9Rpxu
i+YJqc4Ior0IKVCHQtfRVAn+fRuZDBB+IfGJYtPQiwgm0mH50E2ctDaBt//3uD1Z
PvgXPgz1SLgk+4Yocw36AiHbJtZOPfIW3fYj51Gv9NMaj/XZLT8xPf4gF+UnQlQJ
Xt38cN0BJOign3ysWX1QqBsGsqim0q58Xa+a5wemIIgeEzRYm6IANHMBSMhirM9C
fPP/EGgz9Nx/rgj3VUpJJrZIt3HAcka6fkmUrGt/+aqfygkhFVqm8RMiOpyBMOtW
+YwsIjVa8VnjLA2oA2r8R/opRNxHpNkfPqaWHx3P9698k//9IQa+IKb+/rVQ2QmO
XwniatHVWxczlYQQlQ99etT8TgLw7y6fKrCqmq2fP1TMbHRblzEzSHil+mdvYl9s
lW2xGYwblSxwMjwqo30HIcK6NZnEYuqjBHzdqP56+QoSj4sTsUGn6UDIX3hb6rJ6
v+H8TWKxrvlPeUts4liBaxnngpqkoqEWHa5oyrP11+Zy6/8GMZnIp/oNVTU0CTWi
ZXIMCVl32qgzUYiWIz2jwMsEYFj2BmAzRCIeBj6bkuaimpEIY5u23IpAOx9ChYYO
aI6UE3tbAM59WoQqgbAndLWiDKzdqWKbuF9+CWuabMrKgkOEVbp8W07hNWD8FwdT
GHVP1tmkMG2tiSFziJvCEVn7zVZmMnJlLgfNbQcUucvyLVdxEyfKMFAxuTRzlShq
Qy8LPjH++uVAbGF+GS9nZcH7fm3ScmrVQncmiJYPkF+ROejaEsy3yrLbXfnWLq03
d+qvHSQ9OpoDn4+q19y4rfJ6B38fAFHQJofiHYQsb9Zhc8ukvmMsd92M/Z58glkv
RuTaVnOj0MWZoteJYP/IqupEQWPcskKWO3uKhNrPBS2uqk/jk+9D0BL7xGx5zX0W
X7jtVy7pYnJ/mGZT4ylp1MORNT3dRDigObQKBVBoQdk1Oj2LU7JX/W3XOIC4yA/1
6GCrwv05notLiLMoaLHH+QCjRSZKGEvDq8jSMvDeMfDVbsGHPuUocqP+YQZKnKx7
ZoJ6pTD4U+vTXa/vbhFEgS4/c12dwoJgzudSCREth09IZc+rbLj9a/8UJsBPwKbB
MXCaOpuRn3l4Ggx1BAuXA5pf3zF9GZjOIqluowzAAfLjCEM48afPOurkElg7PVUq
1BheY6W7MnIvBNbUDcIUfRE5a5aGClbAD9FHVTryPsm6RbE/060QKcPAT2jGCQQB
SCdGBWmSoN5SfSvVJAfWlZcV3LfHRwM2OAM3ZaKHN2dM7HZjKsje/VdShoJX0AYy
nQuvbJfIqfY9tO+CY62DJxtQNl3dp2OXPmOGOxsRMZg3CJHbK4OoL828+JBeBus+
4Da1P6HnKWB/Yyxm9RIjbk3PI5jyNAICPL9tGoBNwkqlRE1cGMGlFwYDQaSk7XPX
pTQlSP890TO73BTTC2Lq7FrDGDcmw9lewy/8zEDe3bcdx+8MkIrhU/2rxaUh1XvV
PbixLsrRUF7m9yrDnBkc5gW32UBWK9PUIuX7sT2DT9XWAX2/EMnXQOP6KcLNcTuZ
jDQPTCts+A9YRFW2M4fYIFSPNZYPDto9Om1JrUSWBpmgsvETzEJUQ3mrnz5VSGaG
HMQlTyCcvu8epweCuaPWCWO0tc5mDlQskwDJ26OcgkcSVmnWc4Ebhuo+pd0561mb
mY3wmxHK2mnvdwkGUd3oBPMQruT2NabZuBiwFF1LhZiORnqEHdbKNxaOVvkcdg+4
LiL408V+AfNFIQG5xykOhDI1me0FIckQf9SFi7G57Nzkt+t2wHn97vOwJrQ2eW55
zBFCrioPDH6kCKX8JWUEQd/xYHb0wEzRH0u/6XKGobdGGAGeH21QeqJWnWXky4zf
v6i/h20VtLLwsPKgFKoiFCt7slxpPzIel/Kn8p5088UjPJ8mXtQlH5EknjlOd/TN
CW7L2rrLFmSi8U7woDdkNM7nKS+sjOX9J+qhwGUHjqF8IkDqttl+vMlFdusRNFqI
2/Afut0+yryn4kib8nGmy6u3tZN2jAmgZoEegfjPUajnfJUgkY0Jl7ZqwYJ0mivC
rcNVuWxhaxviXKM17JrdLcktVQvVlAmwfLqsTFbfQTl8qomeMdEIG6rBQhOgjJXJ
6scNEqwdasJEzQCsv4j8QCvYtxp0ih+t1Z2YfCLyBCjd70dW7UcH2hUe8DqLQ65X
tM8jPJjj7waEUcrXBzoyXD8MQALqf+UlbR7SIrSpvHoDcX8Oc4WsP+4uUAYcsSZH
WLNL+TKElkFPkJ54qjRyAqJN5pL4pVv6cQbDYv6mDICUHfVIlVuoX2EWnf+ZLrSC
5NtHCbnPS36Q/3xGTP98MEWLo7b1f0hhgyJaH6JKy2fuvzVbjwnfVBOCWySRf40i
jYWoN+BVTan+05Sm1hSfAaLGnKkljQ9TmUVUMd6qH/Hb1p7hvdMnLugrg4TxvpZU
Do9qXyr/gDC9/Y4A9MwTbeUduc0+3wjuimm16FWy8LAendPtnkAG6VTx6EyYxspn
AlZc/vjhmTkd01E4qL/omfyEy31hQ8pw3gE7MA+7uaHEPkuvwu8IPuGju2CSw+/S
Ih8SwcHN0t+9d2Amp8ntPpTXZlXffznvWZM56LpIB+PITqeqXkHbJrvDj2495ntP
Bm3jNphrcwujeIARHjMbAnFiZG/aq1pvb5aTW2T3jja0wNbhVOvWNIjPpmecLPae
+lVfWNKef8epfzQwD1fGAB/FMdFWNsMpXNhkFlv8wMGhLDG4qivKdkEZOM3KvyKp
HT7f4m8rQPmdsT3cJAe6MaPDLWcmQI0vvpNty1bc8NGMPT9OiwfwrGf1G2fHgI+f
nP6lrstLQQsnEUIjm2OFL15Wy3TjQh3Ktn/cahN2BOc+3Z+KK8Jkb/aw46j6VCVA
RhfqvC5Ol8DF+vDKsrJP8a9Z0WuNYrWLzMxdtO0wOCLqb5qwaaq69fLtQb/yGAR3
sNY2HG/+Tw2w4ka9aSRX/fkWgx9zXlpvBeHXZpZ48z1AXlFjSS/b559iY3k94LAc
zQsg85TzFqDNgXLYkz4rrXLTLHjczmfQ/G1NbhTVW4Qc4IDjc+IcWyruG0fStZLR
8tPmq63OVe6o5q0gMbFLNLSQl7o8v8stEJLH9t6uUNYvr4s7YFtI3+EKK1lHboBE
fkyjSJ7jXH9z0bGzvi090DR5HffBZty7OiocnxJPyjGzp0vXRZuT1YFUCJMRUB5n
f6WTknOxDJ/pdby5a4T+XXm8bzHySGQgSfMp5STX8+PmQBse0TYtsipnW/RaQ7T/
u7XXLkYJgVvKBiKIV3pGposoccQ4QLkC4OFiWHxOXxmuisGr5Gi4AsyybWXMcOg0
MJP3TX6b1kpCBHypG5DiXy5Ls9xrCZljL5FaKPzK+/UsxMSSK+fyu+EddOxxT4gH
lt2lPyuIa+b4QDsLlv+Qe4jmaDj/eMp/+4L+EhFezhd/tIg5MD+pEnbTV+e4mSeG
RNFmksj7tb6KDm642m218nweMGiNFTcHqR99oQtVQwHZxnerVrK33e9TZqKTBVbN
nv730qFabxA2y9rcAXMzQlzo2LiBeAJJRIao6mGwakKLErnBQjpmJxW5pTPuh7Ir
M5YUSIHCjBnrYqxJOQB6DZ4kAb+dCCvy5UJqNgkgcvo067pwEk4QETtoombggzp6
NdB+NDfz5Qyc8EhnPvS/O9dPdNXAIMvTC/wF4v+T3H8dm9HDWolx/quE5FTuFPaf
Qa3NLTtr12eLa15GLCqmN/U4236S0jb4nePFQq0j/0blMbBuPZR9H0ZZ5uQwSNEi
/vMsp/Xh7RW4tH+50XqX4LLqpjy1gMhZWvin0iv3zrxkId6U37gYZ+s+TIuEvjeg
Lr/Kmt9yJyTqh2FmYWg7D6VL4eQgJQ3fWzi/xv2V77C27ImQ3xq8ds9Noh94zncH
lO0ojL6RJkMUmgy52Wss6cRrwn4Mmea/fowVfxUq69C29cZoTdx12eDslKXITBK/
F8FN91rcER3h6W2ly4u5w3o4IuGNyyEYeRLEQvyary42M6brNGoZdBsgNLBN5xip
R6xckM6C06GdRbMn5GcNnEVVM4EsZmlfC9jMUf/otu4AxNUKg/xdV35zotvzBXUE
uT/9j2x6RbxbuE6BwPQZ1I2WJ9M06Yn2DK+mYSU+TeDVGVcORH6VSTWOnS/BDsb4
y9LWBSWooLETIKMq+Z5p7qMFk8Y/h9X52vcCVgRycqLH1xvet69xfgAmx8yORB6e
zjK9zbtD+SNCgIDRfZmVywqH8xPsG3YkE5GLKoNpemtL39EYn68xozsCUwzN5ls2
05sO8ls7J5sh9rdDxx7NZnmxJbb/tUHGUuSW9tvyVRtNBEOazW/MIZMLiac1avyN
dGfgg9KGNsmM7W+yLTkzyl2yzl7aWZy38JJ0/RYP0hJ0iPb+y9uEiFtMeD3Z05zq
xinzNDjke2eA8pDAmPH379Jf7YjGsOvmjHcd9VoYMQ8NY8UHVO26fbkjFObNMIrm
youDRwx1vIGwfHhdtDfLEcAo2X37Wn6kQIji/1gtNOBlQyZgZY7bVgBdxmJlaeyS
9AK5+0sdqsJ3BUUvm+fFIGxZDQbdTn/ipgaHjtaqhlN7KwBa207BuQQLSegy/AfB
0UNlhPwkz8RXC/zNDRH9lFax2pPInYzUpEYgOUwwoG6lEOy1KRKUvdrJ/RvYlY11
jxi1OmuL1bMxMpXIdA+yucjQXSxBovToC9fwvwrEA7B0KatuzF7GWC60epm8enUr
woDPrDdwQzkhMOOY+I5bwK1y8S+LVO6HAYEBfC0vNcu5Nmvadqtc7if2hvhvuzs7
9j+wtVRdRl239ZIaIArwyKwim06h7ZkuGGmKYEBq85wPT+YDWdU4+0R0KCCfcDmK
8Rx6lxUmjIyJDsK020hhyhSfPrcTdMqWoMuFDhSNxuv8q0nt6NZ4U9jVV2QYaock
LAlGHD+e5pMX+r2sXfB/9qh6wbaT5DEVfBxURTaikVSQJ1XXDbvR5p9JKh2fH4K8
pw/n9PTvTOoa5Tzs5fUZIMYrqCWB/IzXarxjpQXNJUSyJG0hLJ3/bbE/pye95Ypc
GX93CXVG8l4oYR7q4YnlPcaKx/YZfqOasRQGsp4Uz99KoX7iyXpnIdNPeEdrAJSG
0qJ5ZUP0ETkOR+n4OTAe60cie0K+iS83hTFX4uqvBh4rgCfKb6wVX1ZXxR0AcIB9
pBLv1SX3fR24Hyzvh++mbC59EnEGtwzwntyRq/hn4pm8pkKOTR3Q1YrZ42JuZ9+P
s4FTWZF3tOdNVk9CNybS3rEsPfvpHVwCl9pqQZzlps7T3aH7+DdItDw+gBcomreS
TsRo7WZhwrG9I2WsAALYZTP+z6GtGXR4Psa3FqEIGk4kdLRSXrbBKMoT3RxacWHE
Dy/fMZS5QgFeGvCUD28dxUjnHuECksh3+ZMEqiwDtFs/zObd0iJpbsFKOGM1Vivt
78qnqUQp1PyBfteCM8/TzLK1nJoK1ONIZpI73lcc+TEIRdb8QCF40cxgeta1Djgr
BCDjf/EztfJjljadnD7iXbMMwV+vugtckYBBfXcXEAhKd7sb9GMFsmUTreA/vIDF
c5qavAbVJN2/EhNm+xlXazZG8Xj3+n3+k3j35sw9e16nhAbE4ble6OtBPA3w3TL1
aCFuH4oKLyzgDhbRHM8k0VU9mzAexYcaWp0D4PBXYmN5oqUHT8jWMGNKjg0wo/S2
Ktgoz5ZY1HRdQ2e7iQIaM+zFE7mP+lq291BbSH9ohMQ9F/fJL5u2zdshsTwsvWkN
D+rvpnNJUpSazXE+g9hccsCMiwxPOko9gDd1DBBZLJeZTcW0HhvDi5dEJ7e29UgK
0m8iN0SMzMasuOYvbEh8U+pmef5gZj6vV3MIsymYMh/GO60jC+BL6i8m8nIJJYBW
lS+zRM6VhYwa/pZnMuoLkvD1YZRIczqn3iH/RjZEQ0iKOgMwUbMX2OMKSswG2qvx
x3vrVuLkbRQPyfzJbRovpAiv6IFmrG+1YYbf07k6sVKMN42imdmp54WVOC14xsvH
wdj2LTjlPPrEDJSX+4bjgBJmzLjP+TcWfiGknwP1FNUARBFzXg0C2WbZX77fVS7X
N9pN8I0hDWm30+NGdd3BauOfjezSqnaAU5vXOXI5gH0Pt3NmmhlTc1+VuBBqO+KK
G0T0GOOg52ynWm6SCz7fGZCW4+pAdQMJ+RwQ2A4nqeawHmAoL1P7Eod/KEWhqFkv
QjrM8Qw45EDwBtdBJixZCa6+aG9pnHnEmQ33e8HfGrREo8Avu9nflpy4ZecZH3ic
wqVY2zNlNInbSuKi/ZW16MsewvIfWvsia7o0DGmr+013SMZ4RB4cKrhqxOGvdN54
/F+VsCZRIwTOQ9WGRIGeMAoG62Pn3WKJxaAFfvoNvhZi3Kc/6g3rT1PxKpjK7Dj3
OPST8S8Tz0IjAG6A4yE1PrOT4t5stRi5VpX2uOCWDLnsWVmz13uclnEcwh3d3QIH
9l+KgRrfXp43fXobFp0l3kPD6+Th/Dp3yy8azgJaKoll+ElxAemwkYtAEPGqXsNT
OEpIdfPKQY6k84+kSQauxlnALiXeGqiNnwSY0ulCEfhq4YkJZMdMJGxrREVq9Krf
ed42cNWhR6OQh8rv2IxZRTRnZJ7kWr6X7d02eRuKLjAHbBtyqwo+uFitHdeCHz15
xxm51B3lz2HSUdTTmaBZfCcNQqrdvLyO4ty1P8E/o46f7towHRHpUziRY6o9tV6j
c2X5N3e1wUhHzjYNAzvak2RziWJsQdCG2qzQxGzpvD8fqpvx+6D1vPM0cP9W70D9
lq+oQxuEplDokWxaBvG5KqMdoNfAJSB6jBefhbmAkyCVruOUdcxKdXvitCyqV7fR
TMC1YWiW4lxGYu3gJXmOHHUgJbRM3EaR4lTEbcTFIPVwSgQN8Zwncg5xHoXvdjNV
9V7J705UvXJ7KNLeT8XfDxkKjmq3Bp216uvHAEKz9E6HlIzjQHmkicF8DS6PdMVx
qUB3eC++ww2rNdbSux2gNk5fjJ31I8CIhGDb7ahGgv9w0i1PkO6Om6d0tM2WoJ0a
Y+Gau5Qzr1cGxG6kd04lTQclobLHZu8SoN2tJOpZNe0jxcqUmCd64dqjXlX7ypEC
Ll1VSBb6PQR3yVM2A8A7tmCWDgxPvoQ5O3pEmT0hHAfLVlbdqIDcNf9lE12eKO/4
Kbqk1RcN/cDYXksKlB9J99Mj8j1J1dcnEkw08czIkucUxRhmyhlBff3rZWtGyFPg
Wd55ep918IfFiKF1qX1K/1FYpKALD4a2inK+GOEF69M3rBMIILQN78krzRFWe8vl
kBKCuYMgiNRWHXcZJSdL6CAE537W80nwjWYLp38VMFAS2Gwh46sORQ39PpX4597N
kJNbM57MEYweOGotP99PV9i5lIaIsXYnG1wNW8CNcGH3ijlWfW1GcomVU2uA3SV6
aITicGKCfmT1LNV0D3ANpGeAcP8yb+RJBye7w7b/sOcp75CtIKdUN+YXArT5dKrq
oioamI/v955ziUJA4L7CfbJp5LWVgQIJ4zykba75DvtYIdqiku/Wap9GDC4mRHJg
OQ22HoJUlBTv1yKdV+vXISc972BvoajUVXsRdLnSVrwW/olAt9nkAQKDq20E+kYU
39oBITpNkLp9Qrrp9laPo13+2NT6Btuh1C1WBHKZ7m3kQUEsnczQboXUUtjoHGzo
TV0K2IC2H/unvEfeOH36Qa0rm/3o+QnQDVpxBMwFeoc2j6XgSV0nfS4fSo+T67tI
sGd3xshwXmkbSZJwJi8b/QKWnaWPXv7Lsgc8shQuEmS2AdYURUqtWihe9zfaRHwA
g0sjRkJpAUV+V/B6culs9bl66KJd4DUgY0CtZxw4C25xCt6rPcNsKicvdS4UlS14
MwiVQdtoTr2Byp6PG+iIluwNN1K6Tn2fdGEmeJtnPLcKhgj4ehrNiV6W1xktN+fP
kR9Su0OffWCsRs05Q6zJSsMTA3LC/ceMit1XJ401MtbzAfHe7a9OJJ0UBto+XTO2
OUwV4BLJk9M9smTXY/d7LWLbWUmb71rfMvYf4Ws3Xl1Ipz7c14EauBeBF+NfxORC
1mKixwGb/oBdqQbf0qADRPS+MzOxkZszke5d7l4iIHdATzNGP5B1xLfTVgMyhLME
Do4EOkgLYwfB45FFH8Aqr5Cd8caEmZvBuBsNkjTr1pvCp6JiCudE5kmM6803cj0O
npfd1vLdNXIRWzUmA3+rnxv1NcASUHl47Nzb9PxlTYTqnJTQLzk5poYZQ4Oynq0c
m97pbrmog9Caz0GWClR1PFgaCJbK8FKLJqEryQw+30CnqDhcf83ZjkTHIC5bFNlg
xJNEiRbiN9zpNrtZ4mc2wDVDC0GstRyFR24WyG4rP/oy/1RePoJeDSTNw9772NGp
kYil4eZAuUYItytPw2/VSAMn6hoyoBrmXjpDiHNG27v4GgsjQG+VLtxh3sJQzqOy
gYehy2y50KThHoL188b4VXqpMSN7RB0afEok19BeVoBJ9/AmZHq57FSikiApMNSQ
REqgdPl0ESDAcA11FIE36lOQC6sdGBKTg3GmViiiSS+snL1BsKnuQITA9aV3HMez
eNWT/PZ4lw2AJNmZA+XcrjjCuRwAh5UMksgZRN6kGJ4tzd5/Py5V1KRK+1zKfvvt
BGxPMVGmzrxsTeuj0H1PfulB4NyZvp0yc3dWp4nHzYEPsCr5i3qcN+5au2ZtB5Tm
/Qmj30jEu5MxphZW54geHIEzJO14lJmslCXvfLGTUp0243WmOl8vtbYPylLLa50J
z5QL5zXzeTn6u6ZSio+T8BQMBlEpKdUAsVKryzCLmDsCaYHUD3iOiz1/OL1MJHs4
3lHjV7pEpNHKBSxcJO4/GLJO4wWDuDEDDiPiyDWlHzADqISwof1GgChP+7XwdO29
Dl+4wPARXpd4U7yVIwayHwgRh+iggoVzFtFCGb4oY2Dmn8hVUDjN8Gjvx65tpvI8
O9nGZodelFtNUi889r8TdX4bqF0jPz/HEBJDo8QyvFRGBKefMI8J8nvYMPKwUXTz
VagXmKed8jQZEOnWsvcCN44DW/UIzWzPqFmGtM6xOUXu6PBPa4qjHKhApJTJ1iaE
blN3K3e0H8i6ebTprB/a/gJfW0faeicoGX4Qgeti+BSBhPveYNPlT7AGkDMgveEg
3tDUeK2+z2a8Y4G5EGNpWChTtJcJDIo6I0Q1CkpNbOoO5c3NAM61RT2C3S7eJGyA
+80jjgpwbSjJvYi0Z0CQ11lUwj9gO46NMEll6Z/wNwVlUZ/ycbDyGNL3/6oCYnV8
7TIn2bX1isI8mV//45zCYvcIZubdnJOexhE/gYS50ZVWjtXLXRiis34Mg034DF1o
mFPEcROgz3TFoLwZ9UCgTkKGeIEWLIAtNhoq5Ix84dzsgR1yCCqs1Z80do0jivHL
cVbwFybhX9xdVrbkd/re6TiN1CkG3HkQyc8ieqT3HMlh7sx71TCVx9BSowp32ssT
i9OQIU53EVPk8o6dpibysyVJr8VfHiQMND9GHIHzPBDLEX+Lh6xhPDZY3lunQN3t
XtH2coixwLuexEdj6kD3MOV3LCV0f5Dj09U3E+PSsOrG7B97SxeFUg1XD4Q7ldy/
g2IiakxHvebQvIVqXx+RZZo6d47S5r1suKaJ+uMorSoktdvFW+natUirP9k53kMS
79+oGgYSKUiSNTLP8+pxslubBwDJ4y9ySPwdUeeLX6XqYF6ZL5Wn+23UPs+ktKgy
EfkRoTy8RApoc7CvKdOJwjAErL2AFRccY5PLMKRv8NEfwKQ6Z+5JmxSBP14M1SPv
8mSH+5Y8C87i9j3l/VBFHcmVksmOitXCkQRNY8OTfrNaydQcHSnrifINTR6aj8rJ
W3gFnFe9xvb3IWSIcslX6VstGkePh0UQSP6BWvkBU90Gfb4i4Ijoj8w+RGA8jXF2
bOrtFDRGrfkHYkHuTI1cmgSz1y+RmPJlfC0xfXb1HFhczUlNv/+JX7c8JvcwsQtA
n7hPPHkNmtYciI2Dt3MuC5vgC9zqmtZofJHHmAR4b4OjULicymAznGI8tCZ0eBrV
5JrVOYsIgr4KJYWjeZf3tA5wG7f+3joofjPqz1g2cLOdt3BC1C4mHPxVZbG/G57Q
kGpglIU6EaWzwiXyXFasCFu7NNvEsHQoSyFdjAaYbGROExsiY56HJeTWFgZO3e/6
25eagTb9+Pr8BkPZUvT4ATJT1RiVdRpI+mf2htDg5cd5+IdDMvpu2wDYAseYxFyK
hr8Ly13gk8COouJgQF1c6Tlqqni1SFy0PPCRXo3owOiJIWqjgWiR4EJT7k3g13Sh
9iZPkm8izrY+CV9BN5YVAl79yMoT/A5810EcYQGwWZs2I6ajIOReY0kcEAmhHjmC
6iz6O2BNHEWNB7Ygq5FGj1JI1IgLpFjXLDr+vJo7AbgIBtcc46uWmNug4oT6aaW+
bbgk2N5Ql9k7Zbf26Q6RBL1IEQ9TjzaA466DC5ZpJ8xQIRggOMMrCFKItEucngRD
qNvTnibc7Prlk96inGGjFdv+wkG0LxsKuRPyH8fDDj5gDfeNWCxQIBq2jlHYZ+7Z
yt+mmAYSUG846qdwBARDok42Tk/twhVzT2eGirPzo7/X5dCe/TLrqZSeR/wiJuxY
TP1Zdq092CPAHO02dzWfugSYeEYEz1fEZzPSRB2dPed2MD8MSUOwixhYAUW1tg89
9gOAZ4LY/sKzD9qdHh6vv8z05PSvMNxSKJsROo1X/QBC/w6SsBM8WHkd31Q0o9Sl
KoHSlS+aCBL8Ejwrf+W9Od7AcXWcYvh/b8lmxyAhLZOkh4oZR8aClmpZqmQLA8bB
jsNmiK6XRzwDvEv9I1dQyCKvvXHLRI8LGczCEv9V6VEWm7JoY+rzr6SF9F47GIWl
ng1RWxFwJyxVEArQrsV4+QaVm2O14SujqvKqJjYajg2aGTcZh/+xZ+JOcUtQEmF0
c+oeMTBZc23yOzWgIpHFEN8A1mitUhL0a6T3YMC7oYNAe8LMYUsDrD0iIoU5BFiX
WnINTMThP+jzjSTPtEpfgrGIubLC15jn4fOqbipbmlTkcTPQuKjg91olO51pjvkh
1tCoA1BcLxzGRkPzud5B+sAwMILZW5I6cgv5x0FcBapBAFluVo5pk/mlojy2TDXk
LnnjLZH6pp75tkGZti3qp2TrJWpEnk1k8QZ05XS+fhGr6jUrBoN/yUMHif7Bwuw6
ELTPR7raDXSMOzPw4coQLD8XCegAZi1DFotfdu3zR5y+aW9InYD4pjkkiCCdKsVc
MC5HrqGPFZ7bRpMfB/cUStDUaWy2oYe4cO1x1AzIzNpymvwNav5gsCWqNVS/uxL4
OKHgulQIIa37htmEm737PC3t3duN30gSk0XSIa3cL9fAR3Jg45IreSXs9MjBByXa
FnnZ0isJkK2hegHGPhRO7VshlAT5UKITolQBWnSiW+6zuWb/eYBuXYbNmMk0CHP9
KEdTpb455YCi9GwPQV5ejAwRm51uvcrEwlze+yOY1o+up0PB32K4W8+2OzW+9PGn
MYs20j7uueWidIDg0wZAdhNhIp87IJCkeVX3+r6lAcOteuYxAcHS38bLTC0uImIW
HKIukhnqP3yFr3Ds5sO9XUvTjcd+7AORkVers67OnLwDgw6SBeBqlKtyBAubYBOj
wYOg142OPbJiUt/uhZUqAAaUJlu2IelgvSFoCxVuiH6ZBTW/CvODNQQgbgkgIKCJ
c++9ZQO2nezs2vKJFeCoW8h5urCZYDxoDh/AQhZIYdelex0L9kDapc4nBmw5yYLn
kffRYZ2qvNR1K9Nv7Utb1jIxXDdWVqq59/vsX9tjULa/cPzwY/pJk/FF7WOE59vA
ZqSfGqCc8PPVL25Ie9ShbpUt7XQQI3X3gRlwIkGbf5pJS7F0mQRmaK6qYqSGHFZo
8639u9sS3O6vqgNhl78GiJYPfSZA8YTELWMfBHLQTntW2Jrpfvl1HgynjyiThYNs
l1gu1Bps7SrlNGFoER+X4kclP2/GfV+pF+YwrxMzExa1a2cKndsLL338miLv1PL2
kt6r7IrrQY+sqRub4S0BhwiM4UxtWGPPA0AzZFzhSIHLl3D1O6/hYuB9UMlYm6KZ
u5JxiY5Mi14ACU/RolXQ1gCO8N/SGoIRQdWBiu/uZdCZrPwclUaBfWbD6JLGCbFP
NhKW427vTq+CnLJVX8o3GtFQp8Z4Fr3RkqK4f49r19kh8e7xVGrW1jmLhFIBYQQo
eeUz8O95zDJKsgrUbp3FlAq6SFAN+Tq2w+i4G7boMM9HBekCXmbrveyeYQggvw6A
kaD+yDfED8pdWkexDW7+sSILMwXbFaKJ2kHaTdO7gk4Y8cWvWh0xcOD3ed3CwTHr
VarP75x1tA9Y7eSHJoskGIWkOResKketF8KY11u979RwpxCxGCkc+T7xNBDVx3Un
ogynIY0viAPuPCZeQijf7LaAKo4ywLXs+JLXEPvHNkoiNJwIKU34DSCPekCWL2wm
a5ibKVEHBH6bznmGTmbo/m27sIX7MrgyHLMo4N1r4VjZChoaJn5RSTG6qwQet8rl
PiytR16MxlTwPl/HhRzUQSq1ZhXaaXuuXBt/OcD9QOkKeV127eeKnnuGHARoS1Gd
FK9fOHQXbKRVql4uygOZL0ik8TmRdO9P4IXnI+J5ViJaIUJuQbS2Pz6E9pqPlUgL
R4lUJRljdXPF5xsrk7kTzZoTomU7bBq5WUKC3yV/hBzrkhepVCv14P+m7brNDLRP
ABgmiAIOANf7hL63UMWhDxAnJ7uXs9Ym8yLAb62/C0ZCNnBVF22zi/EQsGk/8hZY
f5pNRVi6bxIwWoj0CSZxlfUvuCuPuQK4DBDVjbuKg4P0qHpEPkGrVB8GeDsva3BQ
prV5dWVUelg6vINry7tlYGyo/1n5bLB2lepilpKWMM6Va5MzoBwibbK0dACid/9N
31q4tv5kJK+P5sXnUAXB8n06dfqCUQlJrQES/ILvltWaUZT4/KL06XT37hnh23wz
+arDiQ76U6cJoIlx9wz9c8PZo5i25XyhETtTsJ6rM3QjsTDjNa7gjGCQvbrFKaVK
No988nZJfNtTiD/mb/Erq5Kn2RIq9IhcyKS3hUB4cVAe9e0JqunK3QgdTWG86HTg
P7KQKRMLvdNKBah/9oXwFi1E0cf9c/649WEiKORtTH+qrdCcIk4r0pxFbZeBUBqp
r8B+PgcE+f5DfGE0Mfz9wAHl0kT8tST5k+o1e4jnhV2nUhLdUw5iYOHiZju6zXow
6A1HPhlN/W3fO+XwMVtfSUSoWVu8zPWK/TMK+vS96K+eOxinRmdb/R1Q2mMDr+X1
B0Us5osfmyB/UU4VsPgWwCCe/0zOrK2kFWVF9o+Ja958t2lfs5OBC+SMzlm9pQem
zkn4wBwuN9o+a3vkSYR1XGqNUr0vdn01tyoraVTEsfg0jBeWgUx5pNbfhU9ls13v
U0yL/qaNygyvM/YT+FWJUaaDFKx5zpKzmQ7m772D0tF/9H/a/t7B+kMO1U9TRlVZ
7leT6vtbMFrmFVnEuteT7Um/9o5CgmULWDYDEBnPdzrtgvieiwL+tiwnHtwnCOsC
eX4y5HmK0IgculYwoN38ZWCyhDi64/MPZYd8TVrCJzaZifZ4LtbySEO8Ku0WW7be
+b2wjDvjPu4fuDXnPob+9U2nK51Rf6d3nm0yPZGeGu1l8H8BSql7h4AyQOMUpUiP
JLHIqZz4nj4uQyvcPbAw/Nq2piXnmoUehKz5UVOJ1qGZUaSeIho0J94XE1Kd7ItN
ArWoz/a67ww+3CF0sLKwCn4NBDdNgNBiqY04FJfS1SZQ4lGTvnsdYUr1yeT8uyNR
aIdKUz8Qq3iz4hart0RvQNI11ALZ6luQFlOGszP1NvI3GXY5aaN/GGFtV1STRlOV
AFiufxMeAEJ03S2VdrCLV6mXVL+rbdeGWthtmaTOw/NQpjkV709nVaXBT+9uBfZ2
QRJMsDdJAQrbIZDV/WcC66yNri1N0dcsz7Aw+c4fHjBrorLZ3oOgHRq+KkSwAyIP
Gxe5gVwp67Mh6cBCAs9E5fP/QK4fIqkXzpcwBq3FGoIzArnjhOXw9/IJydzMEljo
9L+O0+C44vJJoCDh80z0x+wIfRksLACwOgB4EYcGR0EvjI5KSK0iyIuN5HLLMM61
3Wwi84+6qQDPkg9hp13UF9REyjsJX94LDVlibh9iXKxddh6d0+TNdwotd9rgK4E1
U3YXD8CYfSKSh7X/9feskojNO94JJgHlhFsXsWBIsV2oGUVa/QMQX7+RAHqHMZAc
UH6KnqsJkCjzYOBVUTLXGpKsmkUyXIe3bOLQJcFnhdtCk3YfKjYsLI6opRQXodPr
UYo7WbA5WUviQkmnzl0m+uu2+B9Ia53kUkk+GeWxFPlBOCUjI1Hj2kqDIckvJ+9I
2VoXuZrvcfHZYJduPTIYUff6ijNfkX3lBUBbSbs8FDfUew9AIr4O5VROOct3aK5D
B8DEoeJsrPEfo2GaPJIkUL3uDz5NrrnjN+cMf03Uz0ivmmF2yR3d6OfIT7r7iNbY
nRdX8/mNElKM9LoJXjSqAiVbfQoxew/kqUlajmPglWSOLsEGGLm8qCR3+ej9fJ8X
matCcs3DotM4XOkhrGUuBhMtQqVN/lNUEGLF3GelCbClWRRryhqSeSMpXH/zJBmv
KKsaimmDzrwB4ar2eyuJz8/pQXUsagXDIAP4VwzjF/C6iuEOMYN1qqkU0fFUIT/5
mDEn6AcPfM/1ObqsLiLu2aTFa2Ax7MWBTkeGH7aFWaLDPr3FaICziC/A1jpSVdGX
KO4ObL3OakcmEW7operv6k63JFywTwsQ772yUcIp4iOu/xg1LZZYkUqTF8ZhyLd7
bA/JhOATFg67hG42u4zpoL9c2QbbbV6ZDXbhsP/45zRTvAIR9TsLtJCfuQv6Yees
TUqEJ97/BLZVwNRdLamv7STnhxIHGHeWku/ACe6j/kV04BME3FScJCSNXGb8dOV3
Sugfh9HxOH0mWwZRPoeWZDtnOMnfIilWIpihpjl0G1c9OP6rP5a6qQIPOiel9nDt
JgdnGGxJr/ZXrPGuJL/rJcQLWluy7CnWg1Sdvg0HjkkAQN3VHABbSfk/UWdG9GF/
VXm7Mt5FrnYluRUt70bILCdx8cmcB1XmORySM8y18hOwldYkiCeeQGZZmNeC6FZk
JNoKxf+R6EAWYl744rCCZxIaP/+ivDsBd+jyttOlyKvUMmAycCZBsh0THomhkfYf
ONv07ZdSqwQX69QPqpaTz9TFNdwLa+JW+TAOmVJcyWaUV5zQFHK71VKNyc81AXDv
eLhFA5nLopD9lM8Z5UFIFLN3rLXpxoSCoaTKMFM7SU4i2QixMtO9pe9vuQvDQUX+
QzPFUvfCMu8XEpXiItEYL29fhr1UgkKD8kiPqXiV0+mct/9G6c4ylZ8yAebJaHog
xX0LbuM1Eliwfl3fXYEdHGc8pMFFymscbtKddeUy8wTVMzSnf8ZIW774IqP+mOuk
y4Pdo3y9oZMClFS19Yq5BUeY16WMD7csC3WTEm63v+K2zI6LkJQOQM0y3ocrhXzk
hKRA7YRYYBMwEFbLTAxsed86fxJUwifc2OakoONkJD+wqzzOjb0gTYj2cyRbF7bs
2cac2/iplh9tP3Tn7pvVGP3FugektfKQx6b/uBDP+0W/YILEShjbQpUPVnC0ZM27
VZFrcjYz7yVW5tAhKONlI3RJDAomxos+l1cpmQexy7Ssr/dczLe/ZfcL2+YMyRfU
FZByuvEdvEpMHaTnj5U3sgUjBMx65uWebUQYxqA8xJU+5o0kAKdqFxK7xLO3yVRo
K0tp5OhR7uy+8L81Xzrxa4GR9C6cYaHVc33t8qQR8TBaZ/cgE3kv0IDdfEYjjCun
uZ3qB1JGuF4QiRkxbXvSSeuuUEjE9mH5j82A44As9vme+etmqex1QBCDqBzptgu8
PvhvvqcKu6tuaXv3yOLoNpSGujRr0zuqUrVmZbGZ9rN9+03NIkI1sfGhxGTxC1E6
vRkb5Iir5zztvM3NA4GjQwEs7tWfsBIpyWf/UqzPhfomkjreoGMT4CRZNeTQ/4Jw
jPUhmOb/wEeXVvI86sUXp3RtXBwBUDsmbZX0sJQDrOFD8SWNH9+cOZ2juEQUARJV
sHDFvmsNOP6YVdb1JiKAo/b+qcbvG8Sw3fwWW8m+rPfyhUPSugxUy1H14gDkXOLH
vsMwm4KcmyQAAAFiu1OBOJ1xRXlBYaahFS7EVLCX1nsMRwCm1hwhDxTi0rx8SzU4
iWpYxcog4XrOWSemS2H9+icEBOYRlHwxunW8ftpuRqKf67GWPuyMiZE4Rskh2cTL
spQj4Ssb99KMCIQ2YMN0NzlQGqdOmU5x4+szPlHiE9ae6Mw+0kC/bD9rTxf5Rrje
VwacEWtT/g3ekRvT2h9iPp/CkDu5Fxfx/+hD5DMkEFWtwO26asDupsBwo2GtG1aE
eiwGHK1WwWU823bTlY2OlQCVVN8lV0zJTv06tCq1Am2iQt8iTwR+7buYwbjqlxGL
ld8EpE7CdyOA9lsH8F+hL8UkmzIIORK4H4znPQTFdhxcB9kF4ofyjVj36ZVay5Of
WrlaLROacVLu+laisdRCpd6YaGLDfijRQ+oS1QaCaTt13Okiz2Rc3uAnae16TDcG
NGEAipRvpAmv8F/9yOdiGO5RrjBcWj0/x06ZKBuLaXdaDB+8cdZCWQNTIgn13/9M
nUF+WwljkOqTt6EJvYgFKDKANS3FwtQJRtsHVxvn3NE46fIe1h5x0B+jHTbOBfUl
LpSg5QyJ/EGut+B9huNbQD1cLMBJNRcFUZZINOW4Q5QIWCBVt6xm2Et1hu4v5Leu
0vkC6aczEiNfehLeU2N3MtOj5Zprd4gQ9laKOMAFgBWkhVZDrvN1iZzwSNk3eT2J
0jbnoeqfJOucAGfo3c3v9nHQJIYisxU9wjFCKOmoWY92MTYO4jvtLWKJ0RBfRIPJ
faiHENeAPOh8abGWo2/1KJ6mKWhE4ZjqwKRWpFa7+UcVeoaQHJQbQLGO2SSIsD9V
RMFngVqYdQom6swPwxVDjzKfVZvy7Pcc5dey2IZJvrBL46esQ0ieet+3VXX+4xO4
O4iXusWU/DTpLIIueihwdcyBykcavPiep/ly9YgjSa6qrKRtR+crYHii2xVBTi0e
FqgAqio+UFMOqP3hnc1VtjU47iVtfZDTWKrJADv39++rD4CMzoB28jMytF+J1GfO
U2CsVsFxj7fKmFjSMqwynObzdOec/erp1pLK9XZ7Vfttc2LeCnM0X3xoyjN5esgL
DidczFnKd8LuqxlpR58OLkbwRnpgh0WE7OBwHFvfhCzgz7LXlW2/1Y3kTSgAtuCF
aEAlSsaej9Fw7nbMAAhlFll+/3XZiB5aGhIgFnTD8cYTNJRpO6J0Y0/em8e42u/+
OqOP1XBThlwqUQ/0NQzNWUeapVrr90ZNr2Noz1lmGm64Wzphkvq1dXa5aFnRNUAV
Aw+rbD9mqxEZhACfIwCfUuhHMgtti/+yM4I6JsUp250R2fNpf5OJyQwKc3HwEDCj
3SFMsZTDCxv2u3IIkXAGv0fbruVuyDoEnjaVXA4EsRj4pAXKRpUBMFa+p7znzWYX
lRVr6Pzh+6Ju87fYxpzVgqU+caAsdk/G8kX7VoVkR6sGiapcnwHOfE6M0yxTarFh
7RSF6rMLqY9xIzy3CsAaG3QvsnWkwmIL6sa5hsu03oizAeQgOZwtyQlSeJG4WGZq
3V10DQtHACiqeVGrXm7w9Vj0z2uwIo5+Xg5RaCb0cDpQxl199TlGGXyY797x/R5e
Y4phoFmlPNLDn5+QwcCRhxaTauBJZ6ZnYIEQzE0TYBURJxm61A8p7yFQFoPO77vw
rxbDSgqEDP/LHVOugJlHW/Uuav1pmFN11iSTw3gnY825uMJzZJPrBzIYMSH48kxp
9Sino0FUCTdxB0Dp4lwL0K0XP/dW7NrW00ZOkyMlfSFNNNL1888cEO4HiqiZGS/L
UMS11WU7qrZ8TO/+LaWYEdQU3QBl2j163dmno6hBt2ekPVUkDxSeSUERh4x+PqCT
Cth1CLeV7JgfhpU6K49wa78F+dK6y8n5TNLrQVJ70mIUsUFT5b/vWh3KRUaiF1FQ
SAu1L6xNGL6vOx8ujsV6Eu7bKkXdE/WNyoFZiEPtaEyHG/Td2JTwIy9HbGfDZ3p3
EcCR21Qi0OAjPUhBifqSFGuh9uybnl0bN5VVTncwqiLRbZgRBCX1s+HDlba8X7Up
0n8OxcssdAgmJuupg4VqTWpb/HF+AUyJxVyJ/iQ+eKVSjzwpAgyc2kvcMFEJRkx3
2KI6Pnctj/HeJmqqCTTEgw755Be1ZtWky32DMbbKKDA3U4btfowHbtkoLipps+29
MyBQOC+q5dUfZZkrCyI3WC+eyGmdAf1BT5muDVDKNOQXFNIBLnrVAFdSU8aCfkxN
Qf2AzUwvOfqF/MaL84i4HNoPz5Cr/xrusKtcXnlU9NYEpo2erMXkn1zja4Gqg9Ap
PlexVCokVBTf0Jyd0f7sJZ6al4YPCnHVR8SBE0QAnL3LO4TpdEa1KVGbBluLCdtV
G//Ng3bhMImaBFkLtjqiCrOy9N1JLhuvtiAs8HHpT+iAI8lHsosziZpY8tobfXys
iewsK7kGuTX7bTZK9mhpo0neBYH6mORIz+UzcgjHteUgvcNsI9AGjqEMCqM/gzhc
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Kl/bL7PR/QC3UPvheB0AShtzcR8E/KCx5qCGbcZobAEk5/rDirQjkR5+LsBJhm6L
XzwBHNg55p2cBt5xoGHxwqZ8GOWZ9YLgFcyBR7DXYIJv1sG29D6b5ZS8UcWA4l6S
gvkurCPtZrXwF1Mpqba9gyltZwVwDJo8smaTN+lGoQ6gdafTYTI5vdwoZke+UBfc
6KGZtI/RkoClTiMx4Xq+t1JY0Z3FaT21H4fVafMN1OUAGqgPb0kls9hyDCB8t5JO
RStvdMJu2041hjgQX+YdsjknlNtkqWSmJWnav4642lx08dAbzaxnRGwEKV2NuqBj
O7zByU3olz2ymj7vZ0fC9Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2864 )
`pragma protect data_block
BVuNTcs3K/QoeirH0MIlUWYsuugiVsIPYuKQorEF4oqJjt3D0mNvTk/hHqUD45bV
gKBps+BPvnnOQAsYv6YVk6XdFJJZpCD3EImfxljolPejrmxTt5lZMoRVUfAFsINu
BeU56gRobgcv3Er9yVK3RUIKLkdFuVYbOBaW3ZKyKfM8xnxmBzo1gCiteGuN63V4
3BUqTUsw3JkpL0ZDhlh2JhyptXP3jXcn4+cEavCheX77uUFK52PBkM0pDoAfq/4D
5Jq0rFnDSd+bnyaHBJ8cJ6rFrAWiDlKcYZKHWq5lGg/xxVxFPpAjPnOxNIRNDz0r
n0/MjHlqaXFbX8UoHWG2jeAL66YylMJBiVapZt0Wz3bo4L9R6DLrY7qrXlPj0tZ4
Q2BG66D4uE9ywN142/+4Xk+BN955CWaJqGuqePXv/rs090ctX6+j+KqG4YskNZ4a
dC500Sjg3ovVwdkWK+oDEVVf2SEPqYNJSgvyvgSt+HWfTFRE79xgmE2Dts3E2DGu
KQvDRIsZ2Q0SdD8v53qE6Eb28XwbJY+ec0TI9dSjfp8jyEcfPGLbaw5sQTcBXkwO
0iXstA8nAuNXRthetmwS0VMs17BiwvTV4FMnWIlUOSWclYqddPTazXtOI2BdWw4Y
EyGzDKk6KciK/wK+r2SuSFt3eEtJDkRAbAlUseg6wFaK/xGOs4aesBp3bDGM8sQp
Ppvu4AqFRS8BbuM3sJwQqNInEl3xp3oyEAODVlbTkKP4tUftCAPdFhsdY/2mrqCw
o9mATyCWjp5cz5A9ZOV9faeKJixrAnKmnUWgHS+AX/3G/qgKN/MKmUXg6PJWpi5f
VWCygArJgrjuPHZckl59uQZMDhVkZQ+fLsZqClxi+HG8hgmhOZnnlL35fCZuyRpB
eUQnDtq0twQj3T2Koq2G/I0bSeARY4kU+llRlsudER5sdboqA8CcDprIhpoKkVd+
ef6Vu5d3HKdWvQM7/kEcOt61M3M1zcElvIrcw4yU5LnoOwEYWHjBNpj3kXRRAthH
ZC/jbcA/2xIDswPooWgwUimoy3yjBantJ8RIbqBTNkno0r3iR6Xxp4Bwx9ecHqLK
qtH7sVAPbvirTwHk+hmUDK6Vp7mvFBbpftzDlfWS9gmpvuFooFDYI+NIHyse35M2
6zpHweoiIcjn11i2q2toZbXR3ZqbpftA6q/ubYnuSrI5DBoXX1JaLSGJiIudfwfk
fAi2Gkv3wnyNqRCWYxm1qr3MIu+GPvZzaPv2v1gxjkM0xlZryhBDupopcXczulzg
H0zjLS4NLigqKj6iblYbbXXEWz+AsTivxbnJlY7bttH39DW0499yvQkqV5Q21Df3
uZQ7t0PtRcoJTXVzmmHQmQjVVN8SPl9e+bccfKwbOboAFdarrPs9hWX1KW9J6Y5p
w3PmW6JgMsn9jDFPHCl4tBs/1Qf/rhQc1QKOhXRn2Dw3Im+u51d8/r0jRfY1QgQj
xpDJca79SBvVCnQ++Ms4cLUeJaEvBP3ZpSrVJAeC/+xzczXsHRUHR/vLMeCJYNqF
6LXjXti0z6xsA6RZj7rzLGVTxuLMJGycuBGY74cyiG+tpiaiXNMD5aKekDPll8F2
BWoLAuGlFgIo0FBa8tCtxLsrR24baH5dUUiGfpYNwq9q14vq+szghTvdTWe774gK
Ev87Civ2Gk+aLpBzeL1uoOdme4Wv7rfjBIKjm+bxclRiPA/ny3hisFlsFvAbd8OX
no4h+dZg7ilAfp55l1pNTwFt76Q3ZjWsIQZ63l/NQO8yPTT2NDrZlGu+ngCQp1ka
W96s3LAsuLRmFJhP6tZlzGgDFAHXKcHhWaW5ccLMqjLvkDQIjaRJ+ZOflLDkFXlO
XpKLD+49ltAG10WJTWcH+app8dYIaeTQWefz3T126on6ahf2pEEjVynl2uAUuLSM
SY6h5iw0PS84rHgY+mJKRKRxo05ralor0cKCtYMvYTh3RpcqogDq4TTfF4mR2rXf
jUEEs4oPCc8LL7FSVKcDD6ckc1LZY38S9Uetuu8LKLho5Llhyu4ga7V7gi3yMzmj
DRzVosVjMgz7fJOgN5HI/tDZeL0pPYiCzom2OkzodsqgxMVpO1L/KZzx28qepjYy
IyaCv5OLCEzrYmiLDvgel7nGRhoqQ9pxezh15Wj/jPi6IVxpWFjtTHemCzSbI3eG
qG/1YWFVh++lfKuH2xJb4TrrVqoPdS2WuHZaNk4SJ2UIH5aImDAbD0+vGTtP1TpJ
TsxarWXhNflEu1RgeKESO1yOqf360tWdV/921WgeFt0jzwrfu5CPZeYU9cPO4hln
wuVHcqXcKHsAiz9d5gGgZMhSPW3kSwqQeECmOQpyYVCgXbqD509KhkxwzEEl7/yL
vnScitVPMAb2zOJllHcxbOJQdQc2OF7K8PjIZYUvowTYCZ9qkr7ZqnFB2V3j7NZo
cDZ+NkKCVy/YBQbDhxleiUntiiaAaY61mdXyQ0Voc9X86J4RsqHptSymXWPfkIAO
XO8r4B2D8XBz7S0QDZN/y3RwuGffXnnl8TsG7Bc4Tta22xsGLcHnAa94r8Kpwslw
HWuJa24BtCPUub8Xib30koBbDDI4f22ZF9Nn6DXXVK0wYvfr2f0Ks42FjD7JGd4a
3j0D7QfytdEfMYabSWSnbxworsR2aT0jINn71aAltaIoUWHqsNF+9qLn8ygnPc0l
jM7gUGoKXldT9SgKtdkKc6R4VJSps2h+2nMU+SMjuGcNfDWFDts8omoBBJF/nud+
ffODiYIrYKBVQeSHHLQiVjlTv2LeIYDUMMwrUFjXpfGFJystrPsb02KOe+aC8Esd
bW6DQNY/fe56oqZquBt6WL1nLA0GDUlO7EpXI41tT1gEYbeZNXo9yVyZJJ7ifzdX
ELBcEwT06a2ACrlG0zgkmcRyTsf42aDrQ2EXalAzymUEPDDwxOoCgRZhzb8uGklf
o3WhZRaA78NShnUggStouq6MdaFVMLCrFd1026edcZFmg1THpkZhOztYacFEP9Gt
7927NGtmTnqwUE/TltNApNLYuHE5ZhIiNHxYBDvZUahRcclXrVGpDJeeaIyxplUU
oX12JhedB57W8SqzNts92z5lBeXdU5WvabEjVEO1r8P5Em2vlvPyuxgTuOyo3Yqj
Iry4pUcmUC6Ham+ZSoKpXQZytAiN38DDA08umos5a0LUyxYQbfNUHPcTCsXzyWvE
x0gD2/UHChE4lFY9ltAoD5kpusrLgQXw2cYDo9pV0HJAtyOI9Y5NBg4xohBvpqxF
DjPcfkXP7jNvecPjAm8wGsjhTLIQjJMQidUEKPKcRN0Yaym0enTSbXN9urxuBSSa
V6VoXrd87AMSlS0RgR9lH/fG8G/k3q5P8YXMop4vwWm2Ubub/lxDux4FRPE0QwrI
rXyRDUVrDYLE3owFcxb9d4hLgmSCogJ78Ix9+RNH2HdkbpJUMxEF8uIup65awz2W
vStMYytdZbf25uStiMQKVABKTJlShCDQxsTYM00NU64sUMm6+i5+B05Dr+vbWRuh
iqigp7RN2crdQQT5F+SpdqH5IKc0VkkGmUEm1UlzDH7m1eOoxTEOGEF58+bJgGQ/
oKg895Eqp3UBb+Z7Iq9bPkC7oE5Y6I/A0dfCQ5opzpO+HwMZ2JbDujzJcvZFY8h+
GTh8GgmMp/6CS2Nn7Jg50PzEA0zVPEbZ8SMThkJu6v3dD9Ot5TCCmPO2lznqUN3t
oYLFpK/dwU9pFgb0iIWeMOoYycdsuHpSNtKB75Ynwa8patHnaDWQzxndc+DEG915
Coo6tuWhn1o5rG9nepJQaED2Ioy9An3E1/eSCCKgCsU=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jHOQXdeY17FeI/98w+KVSc3mmwQC4+4/jYjOx9VI3s0Ex/tmdx5oJOGsYxIYBv1k
U6YbFvjV6pRpdfXuEmumc9eGZ42FhZzAVwbgwlfOmGeoqNcElak5l2aojPfYfIJr
RcqG2NEJeJITEk4gpYYN/nfZPVQxj66Xoy8darxBWysdrZCuJBa4STy/NxvX6UXR
hfmHi0h1MFlJO2FW3hdAP6BjH9qQNLGgK80A7xWW6Dr+HlTdFaWYaAJ4ZY4kEKaj
X1O4XkvUUmQnQH+/4cC5dGqqfH+6eF32Gxt3Z1f3ZFOZU2clQ5r1jnXcTmG7dE7c
Q8q/w1TjrB574qSA8I7Rpw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8704 )
`pragma protect data_block
ZZQYAuc3LSJ62j/y23Lir8y+Pjcud1Ie84XZYyxHSl6pZbIX5FDRm7xcj9OSXg9Q
WBiiZbLldHZnFVM/X1iggnxjUQQYYYR44c9yqSfjRAZkMfTiNjhTsVYgKpfNk1bT
tX2RF+Vb1/chIVpN8oURaKF1wLNtFVgeVKaIAPhfuqOHb+lzvsHoJ5oGPvQbPtzt
Rmoa1Y7h2e3WqiVinXWEtq5EFziE2gNC7kPrXDCq4DkdCvc/h/bG6T+6joSzVpAb
WN8iHStIREOfotd2u3WT5ry8lUdfbmedPAT5Ig4Jx9+5iD9zg9+tRCSpbZ34GS+o
35NJQ9mTWVSybhUOSnn0inXBpYFS+79ynuLAdyh8FcP5n59Q+SSOmbJJQCh3TMRf
lDCSqPakoLVlBwFlw99m34IlLGqbJ+aHvqDA/vGBkYwmPUFzfLXTqeFyvQHos1SW
v3f+SExJCoDcbgCXOLiKhoPNNm3n8sJYxwvJIP5DrgZAqUh4ghyojomcrYGCAi0c
9Z88f3HZvLRKSIv0R2ZzXraknIdUQS8KIYzvO3htlE4VUblQD+ACJyGKUS6QLUf2
giBh3BqDubV8kXeY3DJgziAl8BLV+N9zn/7BFum0r7BxxQX50FBuyGIMUT+qyYq1
xz4lUWnjSFPKjjXKuRlahYri0im8vd+NXGakc97OQk41v3qvZr+9t58H9IFX5fwx
rLBa16JdmahgkUb8rpX5+OppSRChdRMlOryEtEhd+91VkZlGW0mrYhncwa6BKpVM
TaR3euBs0GzXaAk7zlWPfN4AtVuxhUsk2o0AN24Ia8VD7ulvy4jVU/QOwDCQmrAi
WSUV2kcT/gIpl1gLlKNk5jdYtfA6dFr2sqUcj7X4BGI4OT6ZmkITfySg6EYctuGN
kr5L13Z8v81PvzoGeK6k2XTmRukdKOlJAxIMMxS6+zKS97JxdI5fKs7onOx2Jjf3
GZmG/UvME3m8ooDTccya3kLtkRfeQ3PaUshvLr9RPQULyKeA5EFrRKD3ogVUA+O9
0EubTcaruN+AzHVAdjZGiZChGiVWaGOIEVXZ/RrmS3PO0MtrFM1LKtkyqIVF7uu3
Ug1MJx6HIIlFwIrtBcjAF8ly5RkhAXpWDfgJkZBQ9z3ddu3Fu1ak4vL7emdi+XJu
8ob0/yuRILrC+5wOErqzdsnCF7H63nZyFtA+XqZOUo4jvyA5RUyNEdZ9R7vnrYDj
RXSAo3ZpyvOkpD7V3Ydv3J41VicGNySTaVzVm2v8x9Jd545YyPULwrb1OROAyUGr
lo0Cf2kTTcAkrVvbxpnRJ85wZdOCBppbyA2pHOIynVqCHA4YHhs4IDmzeX/AQ4TO
Uoam6a2oXyG+qWK+o/0DjV2oq+EpU4Lsu4pe1FBdJSOt2qcVyPzL9spyFe31eI/L
XDz9967yi+gAvWkVSse/4Nb/X1grHgwZl/3tyggtpyraoJ2/BuebLfpH54Z19xeb
VldhEfeCI/D3LLBVJ/2fmzjHly8WF8mwMef6PL0lgtFAntFJcBycrXshaySTNciO
cOi59gnW4dX8siuHFuEt3dFlttpHnhfzlsWvcez7qPKGyH19LPx6EtDybPDInYsy
7jY0BjA0rnu2yAmFEWbJGv0dFlb9Ul4y8GtUGwjak7sjnLB0KX9HkisLn0Utv+AO
QYhS/1FZSv9bV/c5r5pVgOn9DpCjPDk+gbjqCANff7Ot57XeDLJrZXDdhKgWf0yf
Bdi+JnNoydscysvTAZ7sNgWCrAI/PfYMvXiBWvRY6pUexG1cEXXuNmkwYq/iCNR5
B3jVwu9WhenzPnoAdYDyQ7pNPTEqNm6LRtb910DK1MuR4spKKPypFnkIpjn3U+DE
S2L4chwrprCstpwK/Iwzn2jS9Va42TUm1V/Qm9n7uFMDcaIFgpmZoikWPCdRNMkE
e4jkDimBjMoHo10mm4iCR0vQkYBk6+jDd8PprX4V3VG6nahNEO1y10NE7ANHwhsX
f+LvAx19xbkkeVk/iM4iB/5BMkR7enrC2IHagmYmXQR4gaqEqmBYoHV2gERgcjzP
vQWa9DBkkAm5y2oFIDl3OqALL+CvMRMfkUz6S8Ikz8I+NOxzQiS0semgvgL4ETo3
J+yEaHdXZ8yVKAUv9kUR+VaXawt3ywc4CSrmRUAaruX4Z4O2J2xEk9VrnN70pcuc
usc1k41K7oZTc6J8ORYpcESrEcXLcrxhLKYjXM+DwT25eLQYCrM6rwoa/BOdQUP4
si9g1Htr4aPn4geJmiWYwWAUdTHzT5I8FC4uHxyKCX9y77+zSM5IyIQrp4lvRsH/
3LXv807lsk6zvjsbNrlodop75JtaXanJP1pO6ClZ2ci7eaRTp5E7chKkQybvBMyj
8EDywULCBp9qp8SEjP+HRTKQWeIwvsBSzMul9gqLSQpac6F6ySjRrG07zmK7Wp3n
1caTdNUtfQjOsrRWMyPkIzWTz0NVnfDK9RKUb7KHUKzmNXGxm9ntK/j2p2d3Bbwv
aqtJXAXB/w/z9jJ5SWZ5ImDBJqdy0XK+pW0GYrn4qq4LU/1ou9inIp3otRhsYcIL
jOvo3EoJAo4oKt9GWhSgIepvIMijD/jMa2jl1kNW0O/8dDNVnqOgO05s5HSDSbiI
Bd98xd7Tg0s3SObSLCcyJv9VoIlKTzpFBKJAjC9otvejOJZcdEZcEOjvT8olf/SI
wXA3KHMn+UNPZQS9Lti3dR3v/AUfiwKtyDowFyxgv/RaUbaovvI+HtXiFPyHrtcH
LK76llb6AL7HtFdtB+hno/ZX673I0mdnmnuZwQlm9YyGQp0hRtqa2r1WW89SQhU8
8y0FAB4hy+B/X3ZOHhSIc2Qbx4IErlyd1RKF+TvKtBpqgEbjmZgedDs9d0/bmQdh
6XzVJWzWsbAlq7YAAEE1W0nSZpMxNg7pUYc8SM4V1aWBvEgMdZVf+JmopF0aYuN9
Qd3kT0rJRCNSjVL9E0Fe0+ttOoxlO9OXCUGyKkXR1wZUNr7HVEh26e/qY93ZEGqp
Ie89IAfQN6mXJ4WbeaVC7jGhWNt73zxENg81G+0zEEFZmayjf+heX/bGyn/PFogS
+xZHE6udSODL+onhNrLO4xWbrZFO3ifRGLCE7tLN7Uq91xHdDT65DbOwe2w2E7Tu
Vcli2T4ThCvAguzDsShrA6yh3hC8+GHKaufsc+IHnI1Fizak1wEl1bT2JcrBxdhI
YcYakqyCXv3y2LMsTzONRcLitdKjBS6bRXGFJTAHL+d6UnowhczAvPIEbrGyEuV9
sLlxRyMl5JRDu4ZS101ifHFcdpFgnut0+jHNA30Fv7v9HqWQMbZiWOrTtk6MiY2S
IffumPx6jy3DK45zABC1Q1vvYIcVu7KSFyZilRnH1IxzhWIl/4wRwSSxaiD15PfF
DBFCUwzMSLLfh53JsBMPkhGzzjmBQ9jrIMxMuJBQ8fiX6RiG1067AEJKuwLdWR3f
jYurRd0YDe85XfJ8w9JC641csbCvPk58SMHyyfklbB0jfEW7w8N1HQElqEfG3i6w
UVhxQIza8Fag/txdrfJYLvMdBCjUTHaUrtQlHeAmniQJbtngX3tO49efPuK+7IDl
iPcPYVe1pjtwXyav+lC1YwRtoE5oKOrzhd9b/UIBmMJkbBqkPwAlJbnv4yYFz07M
qn+UGMWR9h6LWi/L5hKp7acGCtOp+1m6QqXGgbsPkHR+dED9LfoKdcJoVSkK09gg
ZvoyjOVzpxBafXHL/VcNTD0HpAyMVzLjn3wwBO/QTdlUy5yrB8mK/84xHS1uvNzr
eNb5FSddROj3PWKmM6zcpJuKsC1kinH339HpwlOgl9lkWwtZ4Qyo5wVvcEMEZXxH
AfaCW5AJl7JGq9ISZ9C86R+kK7ePfZnQNyhDuSP8IqzaaiO4yDlQ24XLtHqroAzF
3NIg6qqh0pOgbq5FJLo2bBpYni4trGo2VsOySBtbAb/lJtOmkICPOjKHdNJW7TMZ
2hZb3JbUnCYQfOJINNhm7jOUHUKp2ncVP09SgEzMyfynWLB6t6TpCpCaOlGuWknD
RXwqAyKgU/WhXihMpP99P44DsRxdhwTddz+COO28To0LxhlqzEQ6S75oD+BiV3Y5
6mysx8QBuMoentQuPjZ5iZGct7R/2wgjs7gb0FUjhDAby7bgBgM+mXZVjmaHBqvS
8fDVRF25Mo7eMVHXtcm0jzU2JdB+ciKGkWJD0fQdedga4mmBQVRsndr3ZavSnCcn
eYOlkYzvMeuthKRKQXG2x6bSsbP6aGZgvjfvPLCFVd/TqQgU9tX3a9XaWaVsqbz/
tzMKy5tyoRpJuIKD4/XgOfMl2VNu4y6Si3dF/7cW724XSs5fjFXW1qVH3AIGYHt/
nJzrR84tUDr2M7PVSojxdJeul1R/Ejl29no7RWbIln84BE7TPnt8ggfug3ZnqYQC
QeuFfc462Q87sLJO6eJXGLRj8wyMZxUDkC0kOmvWRHFViGL7pzsYOYNbuqUS4EiC
0ehNT0zIEdrsAouKM6Z2aBVJBsuykssatu4YrRiZe2/u3YOhkXcjMp8gZ5cXkepb
USyNKa7NU86XtsX+ZA9nxBER/XoXm5LwK67zcD74ixbK0L+jO0nZVK7vYrFLdLhS
Rq0VI9OTChAH5B5f8AQZoqjMkyj81yQtbm0VotxawySGn6NEQtFLIrPdwfL8eIll
0Ac7bP2NKtY53kqnmGq1HLx5JhhkHuQYSfQAHdYa9U4+suEAg/Udwb7/Ra0q5fX4
OLpF2MULAct8NkSvVxXfftMMT7Hu8CDfBBSdznYvHuZMl+UAogKrx/K9PipYTDzG
T+Q7VzO0sFq141iY8+VXWJ1kA03kJn/tR/AYtwvKJXtfcYxw0HY4UTl6cqgrv3mv
DFbDJptd/HIJtAnIvZ0C7FpEpfuh66f43/ug8BcdO27p4uHKMAip2OH9ywfqk1Me
BFVvYsrWgWBc3f7mLRiVNaJfPTQK1JlhvuA4AB0q7hus1Hp6mjb/IwsGIeA7Sa4H
j8kNyRME3XJn7ntP02toL9TQRR+D6WlUW0RoaqN1uNScD76hJtQJwRE7+TkmJZNI
FZhERLwRHWBZBlt03+41LGjWcbOdyvwIv2zx7ua3/2FbMyjunzaeubPLRaSrAsz8
pF+zJcdg0aWl4U0BEiM/JzGlMnqVDajRvJaYaUSbcfIQiIcCkkxkl+3AkwqLb7nU
Z6c1b0o2S2DMo5ZH17w3ft6BEucivmXqX4g8lODIYSZP0HHe2mnP3jxg7AiSLwFk
sUoZmTEivifJP/KjAFJDNdcV3QZkRFebthN6Aj7pbOWq1s09w0ZQTTO+ypCA7whj
h2cqxATkeAT5QJwwJUhy7fxUygnaYpOyajitJg+HiBcdZEljOrdMm+G1Xfs1XUhd
Ncu3/2E+yUQ+PgGgikXW0vHugazC6Yyo4lYuJmeMYFfdPeLxAFJA/TzgESoKeJhH
0Ff2Cy5NV0xdp7upx+E8ZGqji8qKw9D0uH9gRj73CyVXhBbl6vINCWNut2K9ipRH
rTrFeSecqC6/Baz+5AXVLFyEy/nmBDEoArFEJYHuvp15nhmjssQW91BH6iQfiHum
4lrKZ7miIOcPf3dQ+ckQMs6FvZgbwSFoS7wtG9GmMb2v4Wq/UfypLfP9UIPS5Bh3
mhoXjC8mGV9H7hsZgkm6qItDH9ZpOfu/IKXeaNygYd8U1SQ9hQ6Wos39J9ai8hNd
d+Z42xKqzySw3b7blVdxuoNZJolzYXPMKwutLn9yFvg2n/lqhFw/QdMaIS5MKNcA
IbWlfAPpPr+IFxqfZN+mq1GLKm7EBWQWfu+g66ZRB2MRlUqcVVBynynYg/aQDlfB
khze7bjDcwyORmNJOBE4b1Z6Jkd75lnNFVJAKj2FNoe7rHv5xQX7JKVBnHyaNlMx
vbztnb6nKHcbI2m4zH3AbZRkKdbS5XpbuuY/8LtFMwbtwv6idUwym/bnPK7C69i0
yUhj4A84TKVSPltxVWXpS+AlZDKrdHI1VBaO/GAKCnh6a+UX//4vfShrBXGM9arm
sFp8lQAvSa8lNbgDtvHWL8WQccGgT+/iFE7x7lOu8QegruOgPmR3PLA13Azz9U0J
Y+KkzsZMaCtIG+ByVbY/AJ/SL3RTw6KWlkVR6MoWDyn4GwOvT1c9rGxKguBwBxrd
VV+l0Vck5BwKUyRkDTICkX8rla47NYfAhiZ1Rl6BItavQ6iY7INtw5dKHb/CKBuq
GQoxvd3EpUjKb5M1gVv8EjDwnaa+M1nIa/i4quzEZNpQrP8VpjA81kDDR6CuO7iK
mMdhmeJetDZNWf69+RFc2O3CI+GvLEexLhfLb5kAZ1FjzimtcNtwHHneM2sOBtRS
2FnR2rcuC6arG/TH6wHuR0B/syzseYqhBQSYkVBUITeLlYTUxPw+WcsICfb0hfDL
D8zXqEckbMqDygPLMitxVxH0j2csZz0+fongVEi4KPDgfWCgS1GEQ7v7wce848Z/
tlP+cQUu2jVQnf7LfewmciTUvldLJLcj7fVryn5yjMLMwiu6sA/RATbo/5P3lscU
tji5Anlu1zdC9kP5nA/AyGOf2j0s/tTsa2rhhHOV+R0Rxg3mR5D4nvdggM58XyFn
QlpHcja1D9+jVLCAPT0FidZlDrTH3RwdnUHA6su3+T8cnO/wt9Jlg8bJ0dfo/cqL
74WeB2KCTA6k3euK7MSpHf6Iqu4mCIzk9WmozBsznSQpyFgmJQObPMVW4xhI5Ggu
gF37S+tNhMe8NTPr1ybh/Mb3/gHyp9LCTCoF3tK2SrjdiBSVp4U1fyFhM9jh+VfD
GQ5tNUAGRIY6zlxlR4gfJlQc0jgIhfrIPeqBa+eBHJbU+Uh5xY3io0eydBOpma93
ZA3kJVvsqAGY4hrJWJRZMYfROCqkv53DqoqMSt9R6jxfkq41I56oMRmSj4TisK58
zsj0DZnK5BM6VwqkmFTtbqUGjGc9b69TSb9ssylH3I2wrwcZ/vx9YK03SI5B5LxK
+MNhiCa3p/wwGMAs9PvxyzWKmCryom/YpX2dQrdsZh6EV6EuvCDP5lSn04X6Q4Rf
xgdh4wkur1VoJil8Hnp9xaGdLgZCMkDiJ6zsgYH+7OqwbC2a4WuoaAVjxd7SMJG1
vqXJQnXlnz3FZ7w/Jls6vMV00/1tm8grnDqlo7Md5L2yLh8H3N0CubnltpkRF2k9
YHa75dyaZQsH/Ki4EbXU8n2by7Lfz9bCMo64bia2CB6vR+l2qA/M5JJPd9nD9Gu2
KFQ0sZ6CWSaplZdpQoyPoWo5Hw2j6n1g9TjYIyiuTJkQopLspWHHD0KHUyykjASq
LwQI+sYrjT5aUcAyZNx6HpjmN2s5LiWtrjDDLdWywKyxEu1GADCU8HIOU8FFeFiE
4TgYGYuRpksw3nGlc/SO0MfcC2Ga5z5/5R3lYrfiwyNM/udc27GDn7BmHD6N/Rgs
65qwZNeOwgLojOj4cDhredu8RnPLWMttLIU1jXuTNTl5+uBQr8ZG4373T+UfFmyk
qzhjSYmQbrnKajy3R4wSx6ZgW008pi9zTusvQtTJGNnQWJGEWEezLwjT+hd7XL9K
wQdBoXpn0xr/O61FgKC9QlHBgLGo4jU/MU7mbstTvc77kEqby3cidL4KqaT7UuPi
QR2AXsU9NQiI2+8uakTruLbjg3bCFRQhsCTawsz7jTdkL13Se/NRjU6W6yQYXTMK
IAEgXTdXJk0v6/ngQ07J81FZrbyb6defqHDAtBU5C8L6Y7C5seAb/dKod+Xoprt6
jXB3QBCRtftIBA0nvLMH8dqFQwXyFWH2VMVUvIl46++914WGZLuw8PeWolstqMFc
00o/mblr7elRw8ghUFeiBFaIazj/cqqQ3Dz4kn09yaRtI9VNncrYwfM4NAOzbzuU
+/HGVxugZ/QDkByLXf6F1z2w4Bs/JT2HmwP9h0BbEbtBrBcJb5106jLmXhRQVMzG
iEBUrmumyrQ6lE8QIpzaA8maF+KLM/F1C4W7sJrzoAHU8apt1ZHzkLI3zqjiQ5l/
gZQJ2mIVfPw9SpUXdcmYbHtGZ1X4Cxi18fDrR1kJFGtXuuOfRabCvEBAuk5QZ9Pw
GjL7jwsO+IjkuEoYxiQmpO28OdY41lyGj5qx9Mr22fOa3bzSyWwmNH+FA8abPwNX
P0y5Tjz7JyWhPHrvEHOiG7OGwvjmR2/oBJAyV7es3TP/22V1SJCO4HB5uiDgnvfh
dQS2v4K5jEDm3gmUnciaOnzA5Ct3b5nLnGjurbH8zE14HGIp1s8cHOH4vZNqxKgo
YU8vfBGH4SvhZBx4byWVT1fBVBVI21k4xx5CEDn7/v7Z2N3KsTbHm0mVF4Ua9jGL
YMxVyLSxmzNlW+JnTI6jQ5olA0B64nAjA3txuIBxAITsENRBoDWW2N1ZmGe8WAsY
OL4NSpJ81zTyqaU3/nH7KtYYc+pZIx5UW4BR6X7vad7Sm8oZSQX4FI8pTqoVXiTq
rrc4ksf+GTOWZ1UKKXH2jGt0uUn/+p2PtR+aAsHUx5mwQ6swtdxWFrDvuOMqLa0g
0PVS+VENehnGB3dNdTME5Ag+zn1+AgNlnxE5YuZveDNkrFdZbsRErESgS/wYjOVD
qj1m3UQsXGgyqH0TzwY31TStkiikELGT6DPc86ea5HNyJunwrspFenGAtfJ1xEyb
G965LWUlJixrx99+sxxIETCFK2LW8TSzP7cwrcPE65MAQIugGKVFyTwgzVybKOhv
lxMQNz0NwSb9uHIyGKGNOy8VeImwwIc1quRsn6BPX14nLqnlcatNMRsKkKvAnnNS
wFwi1YiO3UPD3pntt5m6D4PZ7aDv0zRM+0Q8G55hIDjQTo6T5JRdMHYJrkoFjq2p
2o7kGc3fTX5Xj0tjDHN8lnvGL6pJCQy+5IQ/Yny4CF2xCjuvVlx4Dm3AP7i4hEQN
k4fr4HeI5ulBfqWqzmrTkT2bGpne01olUnuZoqdCwlQUqqYl1M3RFXBIH0Grps2b
9BICTAIjAtEBxIZlcZolsrng4rcF8GFZcQQMCGw4RzCGy/hZNH9EFZtqSROQkieR
SjsR3dQSf2AoHNo591Hcvp64TuirIehMP6aDW1rpSpRPAcZyyhFKJkGMV7ahPPJ7
PppkHqbViW0sg23N8RSgSXiVd9czqND6+n5B5RMkYzNHpWPfON3QjJzt+7xtF6E2
TfexiZnU/OdZWU5jP0DQhlp6d/4ld8DVpXqabKxU7puBHac6I3ZFPAyl4lID9JXW
Vk2E8LCwUUMgIfdK1zzvtslmwhhxmURjZoXkLChT+H+pnozrfsE9WyqSWRCf1DuX
S7QvbuO7mgLmkvMFdtLC2cDsdYnb+Tdjhku/Few4/K5K/dqqkRCdcC5d2ik8ZZ/O
i225zjxGtLJt678NMBD51HMl/uX4KvpNFOb2zrVb72PRkA5LwVWaKlo8fwczMbUN
ENo0upOJJ4ExUyInHPJnVOov3gxN4kIXVBjgWgHmShCSfwLVejxFYp6WskqCZFv7
MFxkLPlbpSc3rpieBVLbLKX46zWoCNKmVzEr5JWDps1hn1piFl9456iFlLms12gS
NobzFLELaow50Xj3XuA63VkKkVJsnYNUEcYXA4JC2Di6+HzeBSNd6hF4n4TU1EoB
SmImy9YD5c2L2YeBSBzJ8JhslwPtxdwJV0H/7jvem6ibW3/7EzH4HIGh++KVZbGY
GsxSV9+bxRa0vqxqt7Z6LTrHGIBOPtHDc7lzV/uG+5ys8fjCwt/8QXOksJI5BKOD
gSWE2LGBCsO1XkhxN+zrL2lBSFlHA/uHNOokLDdVmqmclSs6fgZ7ZN2V6JCpB7Cg
FZYUihc1pg89ZwhqGWcqiIrHx3IctSwwI3O8H5oFYszu4vFxVtli9NuC4pvx1W2K
pMNf6sjt0aAlLqikXF9UTP91piGMRNWBTUkuiHu9DY3Mkp9IFkd7rSrrU9T7W4FA
0o/0eFLr4Caf76y6SEnu06pWkHVeXKYxEOoc7J4KRrxqWa3oZGdLryNoNxjxoHy+
r/gPoLCIn16c6LeVybnhkFg9Kk6MifINgmaK79+KYlgomJSUaAQeIXHD8xSJMs8i
VDzoPwM3L+tJ34yK+ja3jsmyB31QCoJnjdBZ51PJ8fVoCAmAGDfAcTAqn8dyt48s
OkLQkDGG7+2WP8B0vm54u+O+lS9FaSTAguJ30ALoDFJ+EzZ9mPrAhq1Ch4ALXR7S
xajvjp8+RYz+nPn2RDOi5z/EYO4YykLMLHnghNhIjSopLYtDG03iAHm68LetE4rN
4vqXDzB0DTKV64qze9a7v/RwxHu9BUW0Q6xBn99X1xSvoKduWnhvNqvL5hZQWdYY
o9BPc4zj0q+gZNpUROoHw5awfIgxQq9Ec41pI0XIDHfK3o2yB7I8hjsgucctkXUv
2UfpXyG4wl89A7baDU+/DocuVyy2ghCfzz2YPfxCRBJGJu4qPjH8pAW63nXdkIdq
1rcKgRisU9qPrLIdrEFklwHHZd5crOAJiquPggesFBmwFfK2s3ICVG65s+XbQk1J
wlAq4LjE7G0lGntZcOLrKcyhHkBMn1lr2o5NObdbwjO8R5pzs3mM3w10bS/htWzv
+u4Q+zrgaVsOesFJG/uDWz7idZ3fmbKlK9KA8wFO++K114qP7QZcbUvEveWOnI1X
VvtGlfMhlJzAlzMNCptgquWN21wDZ8mNe3IJAt2aKSFlUqSjAkBpPr56+YGjRiPh
O2tylPdslJH0LX5lpNdemyvkp25D8OIBZeYi9ljyMQaP4dvib/uKsRuUAt/VBMzY
A43n42sT+YXods9RQinSvd8jXMcvsbHFjJPIDHvn2/2MWMvEznFX7U0pyCrU8mov
7owxByDsVus8elvePkRRA8P2rD/+AHnOoRDvewX+btPpbZtOud3gn29j0TUlpOju
FtubOvBjdr1yRnT8GJy+SGIupqWFjE6DJr0GzUTrVSJimYBEYjr74lnrPbiICCpG
/o+MKOq4SDkNVb6yK5vqmQYBXIplX0hj3YvmmI9iMKB46QWPexF6wAHDTcIJGqt5
IyYeWdiKWtP7s0JmWJhb10/TyXc1qs2z9b9X87ZlutkvXbKhb2wWYNEomDxDmD9V
SCgiQioQnURqF6QZ9Dsnpc2vLB1SPzuJiGwO6IptJty1r7zCeYuAGt7bxmlaOHKY
hnL4evQbf4S9/VvoeIVyqmG5ULhdiQXePZneweLEPq3UEfykqFq/f2quKAv/Yj9X
hn1APnx3XTLm1TIqac9HkBXGN7y7oP0bMZpy2OpckB4ak/NGEDhaAwOyeKX283W/
uIEkXAQtJqIi4IFAH1WQHjq7PTy0eAz6YwRvRWDLd4FsRtGzq4jnhGPqFQa26Kwv
aFRPtTbD2vgo69QTs90v8gBwTF+SxR6GbKCzAEuKggtFi3bZOIivzV+tVgEYU8XV
CK8faEcZkwd5ipJlN8uZ6ETr63gsXB6vIcEggbgVgSSOPAANXZNy3Gk7HtVt9jbO
gtoW+FdT+bQG5hotLCdmteoxCxFHSpUs1Z+qJzs3zrerNhZbnOXM32KNreeR3rFu
tjFf4OrwK1W4Bmwz059wvErxQ0T49xlbx9/K67SHvC72Z4iXEDDBgxjLOqf9AAXW
eH9Z7lu01lJXsnG+qlb4bg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FO/kRFpxx27ELS9s9kWJRhBaLZ26G9FaJpu4MbeDBny9mJtozG85wEx6XQUM3Rs7
rtEoD/nv6/6MhMmCOIVwrYiW7dMcTQqlrlFx7Pzh2qK3TVV9JPIz/eFSHnh6MCWl
Ifc51gmqwXesnwClgbCG6RF64/hJisLq211wpI+N/Hj+Jjx1opBRGvPfgAbfwoLf
QfFGmvqnrsbyD6iheQTSe+hnFCZKv2oJxRHeNPnj9O3tca70nQRsckejuBUw+ejO
V+TRfZGRTEJdFWOXmQi25HL/aOh79JbLKgE9ScSiCASSDoHqwaXPx62tbyqxvkR2
rdQ32cf63/8mkQP0F/UA6w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8400 )
`pragma protect data_block
+HMIf7RoBmudLkux7Yr2sFu07ZjB3cubqjTrtbkBqQPllNMkZQWaDrzCb94kufMG
ti6C7U4j9KjFLXUevn6GnD5QPd3Jv7K4icYz9aG2ppHB9PgxZa+VPdE22VobrDiB
RNOC8HnUOTl/uTTR/WHaG0p0n96tze7RnrodaEIS7PuuvwPZ4qcgSgSzahkvcteD
AMU8H2AOFJ6bF3+2v6T4r/mvcWAHMJeKanQwD0mA3MIKRJCIrZfnq7Yk3ig+Vl+l
L7oyqobeHyne+8Ah1QYgOw1Olx0jvgikXwvKOA+hAXcUxKyDvcM+uL1KjuPu3SDB
yWEaS5EbmD0tEwuYDVEycaIgbFsF3UGHeeZii39jUUT+zeCA+DJYC+OrxC+6vojI
gD6GXSn5goRAhKNgu5h/G8XAhBrgd2YMEFX+hrzl0tPe8cvG40vkgmvQ0L/i0TmA
VRVoP0/F0GMk9rljTH+wBdlO+lV7/Jmk76IZdt72E2RUl9z2K9V9frkb74I2OP/b
isq7CpcV+4DYJaamDeBkC3M1xCYhu/pqV+SG6R+iuX8uiFXrv/chxJ/WcS8LPyDa
xslWwMpWTmmSxskxuhuF8r7Ok09XBJkaqd5CvgD915EXmSmoMMTfpGpbK8javYOM
pY3vz9wKG07bhNjWZgRknFRji+g7mt0Jo/eIFG4eFOOzkOsDRavTvNwPV8kRs3Z5
DLR3urlq15EqR6Cves6xhDNHxkyEIjCahUErwtqYgrzQ1l/SiNhwCByvdU8Bf+XV
wmznPkAOPlIDNatiUMvvPelDU35xlSnR/YqJajhlK2gF/yhf+ugwOUjdl0Fxo2uN
ky7JQQAfeU6zcc4wu2Xa5gkOWqBbIS04TEsb2qTDtGEXTQINd/UWiv5/4AIMcGz5
FAzvX2SGhQYuP8W3xDWsSXcfASJsDxKHeYyJmReW9IAGjvaSspOh9WByj23ZwOvE
hksmW3O4WDIxUllfqeDJnJezdqnxfC5Bay4DUcWb7UMqtHxO9fz9d5/A02yiR+iQ
K60U3P35vqizyImSqGNs3oxwxFjCU1zNjim0BEKaxNKAYGMlQXas3E2XrUTYEPzY
jQi70uJadu4WwBVrZC0dE5QCeBB9PbOBhR5RGi7Lc2XCF63bCIzO8h0PBK9aamU6
z4tVpBBz5BfZjrqaz09vCx9Rx9BLB601JBk0STwET4hCd8hIZPHDb1yCGd1hE51K
FhcRU6FhQRku1ZkChICP5UgMf8rLF4nueo2LjCb656ok3pUqATMLjSXhM/aY5qW4
9WphZ4h3cowhSHr6NEfLLDIqcWByHfkN3YtePb0p0OvtL96L1cEZMUVirt+FWflE
OeWjQfIrUzsGt/iQTEMkt/1ugmZF58A8eDgkOsmWj4LMTCN1b3b9itITcssyDl9m
fzcHwjM7NrwPXTY6e+XBl8jEeAQCIGAe0/8mXgy2BH6CxkS59sS1D1A+o5mYFweL
5IBWBOWe6JYTTS+lyw/5e1vzCHkhcfvZusXv1WyNE4Vzt4eWgulJmnebMHDIXohV
xlGXUM9iMOeNM+8WZG9tSz1RFW9msDXtlrSGIPNq7YGHxTG/b/2AOt1dEnayq0k/
RWfmT7/2Ea0MKgjk1+Tc/rO+UbwN28E1IsINGC8Cnzgea/sEHMiPm3c5OUPPNvmY
/G7i5kJF3S1spTPQ92JZ7cHiDdBE5gSNZsPuem+MNbNNSmkXQHNxnWhYkUulsa0W
W5SBTptaKTSy8/MYVgMehZOxubNQZEMBR3EY9d7SpfMlKY5/D756oOxVI7dgGhAC
LYmWzHimfvFwqVXlJp4nlwLDruxsZqnhlV+TzNRvB60VZWAoKXJe1ZLuRNeb6A4Z
/nqW7ueWsELU32B+zMrCz1indBCablNRXMANUBrK1vgZ8vtSH3WwXn/p8/aWUKUH
f+pHheAAIIZUKwPeBBTLJEst1B8fNprgKF3/ThrnaCWbm9WvSviwmLucGADG875D
01RsBnvg9ZdGZA48FDMYshO0KhlTNK6/l7CY4OqGRUnbeOt8g5C7aRFOHdLt7xFA
HrfQXF7kifXldH7vnbPyoO6w9qIun0Q7TsU7PfZGigcYRFIhQUCs4Njn2cjO/s3O
RnJpE4uWv5ZJdissyx+sqFcJRNLiRxrUmvqkzEkX4ximwFENUTHZiYuedmkLX+h/
Poj7xZOxRTeiwzQAjPXY1Bkdhlhn3G6m/ap9QajWrdH+PbLAvKk9PIk5LCEc2u+P
cFdUfVc/1XTTwDVOz9h+jTBhUNS5+KNGpl5lmki0lBfXqJvxzfP4tIAl1Y2O9I/b
2pAmthB1m9MtN2db6IlugunhLvGZ8wYUJJ3XGPrG4vtV4AB3U1lb6sVAQSBuxScR
6qd3Y5gKd6rBAEHIiGdesr3u7XVGuTStZtfzFZLJJZ6UUVxTbDDqLCHKQsEMKABr
JJZRNXoKxZvNwNRwq2D33poohJ6ZeN7hcjuFk7MsmK8fQZwcI7YRNWiWamZVz3pq
04S71rFOy2gYOlWqls7ot1+dv3MfyabVF3EsAeWM4JMvzF5ria9gLlCrh6vOcEVA
mzUKV9HXkPsh9+xbqqUxdN/E0JPMZmP5/Dn+9vX2RP2nM3qNVZ/6f2ZLmzHNATWm
YHSFZQEcCnXJm1yfqGInjaXdOv/aQE/r6ak6lseh2/pgwD54psdVTapsfiD4i8iG
9PGs+RHZE48kSvrPQwDXtFXzTDLygYEwLoNs41DKBN7qIvW6D3+1Sl+naCrpPX8x
pfbscKRPl3fswr56hDkv4eTDj4FRtAnbB5sUyCxMIqCQf77jqRBY2G3nttBEOs5m
HGgqluaS20HFoTdFPv5I6y9BWGP5ugLjg4ALtluOdhvGSoWlD/tUjuIkcI2koGlB
zHyACHY1ElUV/fwZuJB3iSQChdoUFg8SvrTLwRtDfmwiyW+WAkrYl2ps0pto1nmx
CMhJzOMhzoOZaWwi/+O8KIpAseoPECPw+ABBzjyGxB7KK5o9K77updJpPAiEAKKG
LI/t1IjciYLHFTIdturywjFatqi5lTS0r4WJ1EDUzR1uteOF7ksQC8Ky/jKOtLyJ
Qow6Was/gULuaE1HFVL9AULn1W2Bow/aZoIosziEqkQbU/NC8tWBXSIMEnui+MaC
HY2mrU+BWyFGcYIwgdHhlHoV2YR5e4UEonw9r61W7NUPQJfPB95U33sWG6tdJ6yw
esJlfYR7FbqqOskh915kU5bb/4+EHhvvrnFH1OwNHGEIRVxD7Do14ZjU/PvXzcWM
J73Il+JrAqmzHjCKhaOw8c1im4Ou7fSQasyIXljy/yVhRCldhZcAnR5NMJqzynOe
fC9dKbReYdD9CaNQAvM+zqEzm6im82pOk17hIc2rMioQJ2Z0NFCGoHZVW9kfnuU3
hbL0jCecjlS0/Acl4sCU1LM+PwpFx6U5wbtNa+P+Ku+IIqbtvHMoXoUJ1h/2+UN/
P97wUUuphrWW+mCb9wbb0thspd2q7se1dHpi9rjcBGBCzK6KWXfg9UzH5OIqPTBO
bYkWXCZAJS21s4X4xSurmd/VFWsS2orokN1PcMbOvbfXnqQzUKpt5bNqTHOsXewu
nM1311Jv/dUi3uAvCRcKf/qjCHqN8NP61CEEzj0ZL/dlsdY1wLt8ao8sBALdd0Eg
lvF82+FH8M9R53L27hYrE06+XgInQNhv/ky7PNeYRy1w4RcJPPU3zSBptFO9egid
DIMWwqxtzhpscP8ac21TZGEKRk3/47Cs+fVP4kKdiRJJpWrHJ67jO7yAde+R63JU
rFpeQTkAyktS9AOeK/uXty3zQbOto0PiML02Q6wU8xuri1OJK1SaREyocCtsuMPb
ngOhe0EqYcK7uAlRVj+3c6HHOAyCRlqH5JgqJh3WuXmtrFyOOh+7Ff6pb8DTZjey
rcf3Uo4cPbmLSblPD4yLOKQTdd84OhpBT7iXJwWYNs7GX54ajtNPKc8aGgAuteOv
ISaEFFMZff2vWQFyuWyjdJKRxSa0A1729JRTYNQac++o9Fxnb7S2y8KJXli0S+IA
vXmO+YxoaQkeodRsb3LL6901bHcIYqMhMhtHtE/1Kki54lmRusPD51Jf/oa+utdB
R9uOiGf8ysyflov1Iq1NrP2ymV422EGzIsQu3omCq2Fk0WrbgiPFdhS3OaGzpCcM
uLHczdS/W4AfkORiqtbOm9Rx0ws8VuCMMc1mmMiYw7RzxpabHOVpqCbZtTETH2xs
4unjuIX6xUJ/ANAL4fbwue0SwS7sRewXb3RgPqwvhiN6fghc1+Sw/z1bV4nHCE70
LrZniccGB2ze5Uc1AH/0jQiq/PPOgE5XeoLUQuwqN/+NJdJtmQizCvokQIWa7G8A
bJJ4paN1D7iMK4IwJV3CvEhi2W5rElgcJoSC1tjCDSnnTSZ6pOWE8lqL4j3Lk/fC
UPCy7bu3vmZD9Lq0lY+rd2DdLZErbczrxUWY8DD8GNL7jTQo7bMAmlsuB7ojYPrw
wmpHwZWKSPeOC1xBZNuzpOuw4MApYvyh0ZvJECRGqXEU/Wj+NsVokgL8CTfVZnlQ
Dx5jburCD6hxobOrm5x+21j50x5wD2fAnTZA37Fm9DAS1MezEXL2I4xveMzvf9TU
2UJKxSOthqWhH8VkdeXbfP3S6RpRJRh+xI6mJE9ZjqVN7A/Sm+JYLwQEiiY+gN37
eY1foB8Ca0rBcY5G5odQAlQm09t68dqMQpoeuNSBX/uv04NjUkZG23n21wRHb3Yw
2s7xzIt1nyqqBgICMXEP03UOL6Bj8/WextIRPaWcE6Gx1XAB7lHpu48qimrvnQjb
ro9urShh5BNjUCf7jbCqygb64wITO6TCu+/XpUIHPtP72embuipPK5BRhnAXvKSM
6osLo8a95cqs9ue9AM5NOZvrhlOCWlWIuAWLKQzjCkkwkX5Avt9IlJ9QzWRgamEk
Y02wbqr2hRTbvqrvoILsWXtNCSCeThDdHYLhBZB/ZfGp4C5UQXrAhB6BxMRXnq1R
lgC7OpqdL8J5hIJx5E8sCatSM9dS2OOI+g99pApf6Yj6iAApt2aqy99OGNo4b6tD
ZxcaPto0jM5vguE0ZZgB85HKXurYhiQS8F6Ya2HrIUSnEj8MX5aniCHe5S9m9FiN
eBQ/pydzAvrRcz3x2I0bUX3qvQaJ6CjyiQay0bXyfAFzwUrHKXGVBc3aKoW1PTaG
n0t9nO6O505iYnWUhm1ToOI+KkDIo2LvFhKxKEb5KWQ7/E0jG407TaNsy3HeDoS1
7wxvPZylRD/AHBIFA2xHpyFGcx50ImpQAeqjY1DtY6NlwBeCldRdRsRG2cnxikqq
EBKsOemEvHHltwABWYP6Q6HaC5UpRR71OPjqfexrAtAaDRDqQAXPmiaBsFSj+pl5
+7FMJvyHccJeGKvRHPzRL4TySPxnHAYCeHTQqNLID3G9dkuQbUgZLJNU/ylTBxpo
//QBwBGvIW5ww+Y5oUwMKIEJ26hZO9swFAHUslJBSllGHugJsrNYvquZL81MTjGX
JHfgwWBakmhAOMYc2b+xazgt3vablf7Ix9ZE46/ZG8WRgMVvCutOw+kFD/sru1Ya
98UltDFlbQjk0wIxMEjWtkToiJ1E1iIHalPwuHy5nyhBwGgpfiPckyKdqPgGTgxC
2LU9N1nWddJVQEMXvH8c3W3pplmPZQzGrnKVoaUdw8kXMffS4Gn/4y45jemhTljP
kuTIo9t/j7qfC8xeGaJ4o61Q7XLsZ9VG+PyqSChm8Pe4m6CcP732Nt98vDXaHPAG
vK6EGqvfnbhzS+u6MjSUXepaTab9My3Z29nc3KLwddX18975jrKpXFmsaHB0blOK
EGXj+ZNDK23QaIOfS6z1rIJt3aV1P59aR3fTGqnJKOpLGpStRksXaVn9HthwsCrB
NjvoqiqWlIVGlwWu3mj6vNq9+ZD5fR7ne+iaO88d0GbY94AMPofparSdnfmtj8T2
89PkiFBs+sb1jZwHzGxjbiCEwzENJhcMcNLzpZLJhDw1nxxj43t7hjQ+VCU6TS8O
AXOR5liWTUTErvG0/FRaHnIQBfuDZfUz+MK7gDGPOfqgycByGhVVacs8NBfW8j0l
H1rc2ge43Kg0zM4Uf9O3pLXipx6ZBfAjyc4J69te92BTash1iPE8IvkmKphO1LBe
Qt3NTXygWRrwwCM4eWDP9GFnBrYhuPiF9rIth3a2qpkBjzST++4/00b+m0XcBXUB
zUxios9DzmOHORsvKJqejyoTslBNTkx5x31WjqXl+BhrKiaHO2jotKsX42RCuWHv
TaJNceKKlpFXpeCYUBTg1c82r65aMHVSNuI7VAoah4OJf9N7JAbFsuEGw/AA0IbS
GckFrPezDDkSTOEiUg/HJcAKnFFK6Mu4Z/VpUnMFYqw9iaHhpyTzuvfFrFp+Tdv2
hvN1alDurTOlPiPtOBtDkSgArRAvdCiapia+Ol1GbXcSXcBhA2mhpPRY6WhgKfPi
nvw1cL9jRYr38HtczkM2Q4qJ2thTrielFGmbuSCDCUW1sHR+vi/F7qf+zCaXpyiN
PTPsIIVnbslLUYwHBih8Tl3w3SjJtiaukYgeORWcx310062aY9zf8R9CXID5GLia
98U4PsKG0pVp5jY18qGvEgOBoEgpmUi1/PV5TjVbtd6j5gja1vFqSRwGLrjltEG6
neniNY09e/Al+7HUv/u7x5LgRhK2i4rPrflCOC6iryfcTHB7YXU8ys/tCrkeJtfC
GelPVNVzH2d4D5Z2vo87IKybmoyfZhvuiRk1b1VK9+M9INHTHZUe/RxKvggfmlq5
sKJg9IYp4ArDn9DOZvTjqR7j6qip8xepQljTOA2Gq6D3Avw8EoASt10Zdx2a1O1b
ltOXCOoE/O7RZhOBdfWG/PXDiJ2NGOjG9pyN/KbJJu4i+0DXIyC2Qe943V7gXTlA
qlXmi7bmOUqMrkpFEw5ouwvnyScx8XWya7VdAWL7HbdIsalyhQYY6Ter//eyazGQ
vkIOd0iXl3+G5bzD1D+kJZgSOnRyu6tr7h4mMywhOEWf6uhAXuj4FAtNZWSPgsJE
r6dLUrHNMmsKtFnC9SVza1nYeJPLgqLvuhy/PcizPGf2Y+VTdoUUNa401vn9DQJV
gAyQR15cNv2zmKSJTfF9/6QXMGN0Dnq1bO/eLrIkd0vLJfL8/+Xu9mDh8DdIvjPK
KlblXd+WX+GBR3OUoe/KO9xnQBdYbKHypFP360Mx3RvnTnCENtxLLX6TUwMmfr2D
FMV+6iCeTmSiRDTyMrhGAJz7+5tpppoJiY1I0Xa+zVt1oEqqPfnt9UfHEKurdr5h
wisMRa4gyTOME3qfcsydqegy0gA8OrSaV8RzD9sfrYOlfhOTBnl2tJHZ3af7Khby
KNgOjcVp/AngyVK/pbTDASwnQTf/tNlWM5rBTyUlAWvs15mpTEzO6Fq2KOaoUw6o
E356jpZzoB6zbqHhbLdWjuGEDSfcxrsM7V6L+MVwHOLeCiLOvh2H7VWEti2dByy2
8Zat+iQ3T45vzUckRTVRfoVpQZIE0JWzQhDGrnLjT/pdVMnCjC0VVoNJTiu025S5
UyL+YGsFEjrQ8PfpAGibHKhYWgg2J2BT6JeYdGLhZrlskUn9vv/0SttX0BszLW1x
ENVVb6EeHFQHsHZ89xpvHDd0vOMdUX8Gdn+FnxwIVMHUWJjor8227HuPb9WQ/a5u
9oAjUk3SEvMvEHxt7gg1FuvxGapLtPtHGMXsFr1OhFgFjRzWUw5NV+5LcmUSGO5S
xM74UE2gyAGiJPYJyq5yG9VFZdgA7qzbUbzNoy9fc8o1BqgtVSQTSYvfzlYldCZs
EqF8BsK7xDaftCWnTKu8KUbSrkWGWjdm/Liq2SgeB/3/KRDpjRBj+nWhauJQjZSF
pNwaxQzKN8vlNKV5qw0SUWNGN0aGODRWOzAnkfkhJpSQEx4ZlXBlVY57MUKrCFe3
tBzKactFXRNwAYl4aJLgGbR+sM10bz9JVhE4ktPeBIGbAJtypRjhVM/FEZTOx1Ed
lXOB+dvwsBl1y+LELh32Qe+DDXKLfGwf4c8EJEMQ5YX8uL18dJv/9NXqg80vvYEy
uAEv0urEEd6jL867qboAHRCxujlH70POY2PsaDb5DgcEQLPatMP2OQ+i2yH6cTv7
HppVN9/ilW3+6jFZvEg1jo3q9wig/Qou7s/wfXCV7a6t5KxI+k5936NSXXYz2lNT
rukC1kAT2HPaYxknmzDLTWhrqqsprENdq5tuMVh+xeI6K9W0XSOghQacqXIPjQ3W
bVd+vDlIr4hRCTLJybgAttEs8dDU4d09meqflxDrPP3tIKMzZ8YR1wZaKeNEkslJ
QnI0npOFzYa3aVS9iVtOn8LpovwFV/2uON02wYxlpPE2CtjIRzJz7B1w37Aiervu
RI09u94FJj7DXOJyQmG1sJEfPvGpV0K1b7zNQKfOf5IKLfYMjj91hHQwP3sBblNd
T9M91vInD6FUaQxkjoc7hFfDH4+KEpXFCvFiIXhmOa/w2t5pQ0KyytPGKYHHkdX1
R4a6HTOE5T8IZW2KaCxEHoLrYYPdhQBIafAGnjPn/CujiE+szi1njEEhtACqmzgy
2zRftunx2zs1COh1Sj1D9ti9It3R/+nl0CqPQRT/yztcutbVovKpI45lriJLM4sh
LOKYMHr0d0zDQYRUsaQyTRKigpdve0xRJgDd6tdXW/4Ikx4L4sISNW1P9U0KhGB2
pKzYp/MFnZAiMyj5aBNxESc9zd/ozx3zyj0/FSjjltpj3Os183a4CiX8/TGoJ+QF
hKjMxZx0M3ju3Gg8V4z6/dCZeVo4q5UB9m5VTiHQ/S6A205I60ZupDXiWMZ/Sr5D
ppKTeZxbG0vWFJkowbKNUghDupabN32kbDB7q0b8/Hjztm0Mw+0YnwydIKY0nRSX
tzUzUPISwO25nnoYrWAtGqolqBOPFjQZlN0+ZsNlN4x8SQ//0VwheWyDajDexYSG
u9XuY991Dy2i3buCZifL/HdwHn+OT2jRrXI+531qZBB4kZZ3i9Y3Mdc1foCEcQMB
RqYFmXK6tGhYtEMnnqZ0CdUuSxaGACAEBh5TIdYpNjPDnnEuy9TnyQrbr7Oi+Sei
EzBSWZS6IcLvb742IpTroYvG1hwNvV+mHAqlo1vlH45fZpzWcM1E197H0VOhr56r
cQF7vCAtVmRNXm1HyR51V5Wcs7V3r21j0SgQIVKmYQNXv1u7oEluGMAOXhyQRIJi
2SV3H1GCXQHVCPiJGwUfFoyulQHfXqbYFsKizL2KxeRZBPzsDabRsIUaQ73cJ4tQ
cnVf3jzGLtKEcNPTz7JMEcye5HQ+wcS9UvsuitTSxc2j+0m5t8j9KM3uqKVp0vdX
zmzyn2ZaYgrP/lBtUPdcsTDJnMBZ13ylslz/pP+fIQ9y0BDiNZvCWGpZ1Bwr9pwY
3vmm1bkVDECjiOH0RHX+04qBaHRRA3/cvRRDZnc+xWD0zq75dpiunC4clPGvVce0
2m6J7Vr/dFQSZJ1s5yrrfO6gSUqHVyeZ2W7fuoLhxe5TAneJgy4k8UHufT+85yn0
vY9UdpMRkndy0QclITqN+UbZ1yXA0cPrNHzZOG/uoi8byMRqmbUY5ABqn/x1Py35
56cs5d248DlM+7+9FsMiebG24J/jUurPQFTKH67fkg2Lg+Ze/9cIoPO2ZjeGQMjY
Ro8ICQJVvO/JWQtPy3eotjwcU+kiYTEBwQl/W36XpP1HXhrR5ySoB0VIrYEPYFlC
N5xiebLcwZNyWfxEdxkk1d5H1rsdS/jGNMXmEq8y58qWCz71fjwxv2ayPvqQQteU
4Q00Mfj5fHhcvDMNX1zJr2Q9rltjLWGTtVgxSwxlSLi+bVT6hH5hSIPQQbE7q8p8
AYVTHgEQ3tKlT4N7loSoQmRVSSeurM/BqxrIzvgwGgDmT46kHsEujhaIFg0zd64U
P22BLZnKOu64iZObmkX2dUpSWtSrhrL9fJQwCWzl1XKNVdPWMwsdPtxsWGGQi9Ql
2/MJNh8jrpZt+VxFA1jIj3kYrDVTLsdXduISSRUZ8B6CDgvR9fBIxc+jOOTTxNjP
dqa4KjeoRuMaLZq/jwiHqnm2HygWebK2P0Sod6qtv7K/TDs4rpCHFyr6m/w5GqY5
RQ8C6tSghUDD0NurOc2tWulfs7+Hg0QC0zYv1cBxeujopSYQskXsmuzRY6sRoWVo
4vqaco9zRlFsaZutpToSLV/6t21mJPGyl7QYT8TEaA48eRzHAffMlMsw62zkUHyE
ExaItqgV2F6gLx+Fy1phMMQuiMG17HW2BER76yCW1posVYuZA78HL2L6tRFwEmZH
Hkc2ktCKuga9Iilusmk9/Ynsgxlka8vZ0NQw5NtJUNH6XY8wl4f6r/3i+OXQmeSQ
Gr6g7OeeFgFL9iptpCPAagUhsMS21yzSF5TYHpPb8zBUn8Fm8NgGOuTx/lqdvMCS
QG/wOKezDzACVkMBpHbj6jF0rVdmrD89wHtG5buXUCAOlPrZYDr5LNI9AvdTPmyv
W3BwaKE87wFh8N9vI8Pl/OdEOiCgFM5OlcSNeYJuVdrCYhc/a8QXNaOjMerFkJDR
c7SDWjQP5hB0cQJLHAwEKhDKSxE1NPxPhx+eVHjE2M1RAkbtJG1GOm42XQTjI4c3
5ep1rbAuMOIPaSma18mju8nFsCDNVmxLwf9TdnDpr07Z2o06E3aHAJInU7ctIMZ+
d5hfoT01gaPQHgk3eLQdm4T7ZX+06CNxXXV5xmqYU+PbntfzwkVHM9v4DDwCxaeJ
NR4/Ysu+Cfzz4RUKwdi6v2x4XwQOQtEMtElOrkRgDWjrfrZiLIGhpqeGPrfwHbpT
VE4FiFcUAsDau8c3eweosQ3MIWGRfdpqZwlOeGH0ZXTIQKgB4f7jK33ACqR1UXDq
MZsGvjP+609BiixMyUA4/8rVkw0+i+aE9yk0XkbeWpCW+PxudHtyM8O4NASwaVyH
GGryS7rIBbR8c5oB9sVZgkPWW53cGu/RZREW+o1H8kwe9N71FupijRWJES7SVPBX
3MLfe7Z4uYd5UiB1YL0ucgX8M4s0CWkBn9HgBm9F8EIPZNXHra4IBPP/jIqBi3Fj
ChbxYYcUGhrnRnMcJHTffnTi6EebW5/tEv+umrR35kbe2QXETlYCU4iXJn4CihwG
3ddYFz12DtmjysoNJ9YtD4AlJCVRpfICkVLagCAm2XwTDsBpHX9Lgd+6IaEEoHQC
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nhtydikaxM2AbzQHG1GdssA+HF4SWjTO1Fk6vRumlAtaphvZzm5ZonxmKmWNtFBY
6FDjn3kfLM5is0g8+42mOSJGQ8Uwp8iwkFXF2Hf7tbXHOm1dtZZ4ta6TsMIGKjpF
oa7BDw9lvlfo/b6Za5DtvzRp/GraUJv+DYs8DZnD+te02R55OJ2eJksiex7AkKBg
q5eWSKBmcAFYEmeTcjC7CgQUCrN/izTrW02srQoQGndG8/TUuO1LQximwpXffgxz
roIcEu6BcBIu/0SNVMn5TwYqf9TZQf+pvWZQirMolRtJ2MZpERGb2gO/nxa6Epa6
QRZ3GoMAB0N0vOb0cCVSCA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9280 )
`pragma protect data_block
lRvTwA6llRWzVmox9KtUApGcsxBmU+S+Rnb+SsLQvWWRlc/OQtGuAjyJMNZu4kS2
qg2whhgg7Oo9CDmVEu/rCTdjgN4Bg642dT5aKgeyGkGI5uZHz676H/0B8n+dp+yB
WNzoF2O4HBwpCQoc/f3qKvm2PQSzU3+frzmf3C8pV954Qz/2lqbNefKEx6vkGBc3
VTqsMm8wlF/YdNWIedmfAgGIFMj40gMDxJiLmg+uOwThWxNcuQZ48WmGmgcEJTa2
So114BC+yYjXJCPQ0ixK7STT7/KEov6voS8Sou7e0V+x1aLFDA80v4xOWm/Ysfva
BPNNVSAVT/uoCVxTWSnrUmZ/Oevb8w6l2sHB/nkHA1t2nw26K64JaUD2OCsz5Qsl
5xr2bpaPcXmsM7gOM4c1Ut2vjQnIBNJky05BIRUC/+BD9rYVsA9owYV7CTbXcIgQ
qqHv2SshmSW0IO3QGXhOBC3IRiKqZwamyUM5m97Ct560HIhxc+Sx5fPZkndWBowD
Spiyr4LdMA7e/XnE4pLQLlPgXbeDb1Z15lPAS+T59AOFvLM6eRUc6h+cH9UCPuvx
PQIwDSaaXrn3v+dyzSxy/L12+IIveJ9P0JmKQ1GgeC3GxbfRdt794EXMRdw2jO9q
108S4xUMjb3q6kjPDXiTJ1rfQ0MURAcSGoP9Q7utz4jThzxxjZnZo7HK85UJOeyv
oyWujDIJgvjL/Wl91CNbASCCf3mvlfkb5gSHBYajjcEN75YM0qR9zy0BOf51RJtI
4Obi98Ln9A1E78eVXMIVvMGT0JGSbVmigXmXrG8o323J16anx3t3x2uXHMX6u/lo
niS0vQCJAjGUTlFvU+bGjeEF6UBw6lHjO54grlOk+XBALu3OPBWGMF76S0bC9DUW
ZJA7i6oqfL41EFky/eGNHe8OYcPFcbdH/aSWeOToXReM3kqjdp5njGdIOoA1CjhO
ytXqQeDskxSmxvV0iNGITz76u7wNwrKFVSyBqQsC8Qg4tpcBKtkWu8rW+mGLApW+
QS0aVFVygq/8k3TPQxZ+mHSkD0eC1Pl7w4HK+s7RE5IfI505eXddRVavYj9AK5YL
GrW/U0zFYMeRD/GFCSUdbwyodFLNmYd5hRD8Upr1dhuD+OvcfFiyfWDPgwf6eW1a
o12mF9DC2tIrpNKXntgZKnrs5Blmhf1HNUEFmLYyC2+0ZC0VctWh52VF4huhIbjf
dMHK+1+giiELl3kT/+2A6wuNCdMPc93fy80mruVESdMJqlI4rGIYdwbJe/c73bv8
8lVhyRJJopi+ajkhicrMxtb2X902TF4M69vjaiAygLf1U5IJ2BJpA9nMpORI0xQo
BRXKa6SzEYiFC/OW4yITChulvaU8MWXwgaql7T3t8zdI1SkFy/tIqwurJHjpx6U7
BjqzWHp9nPRwg6QMV8dHFMWscX4pJQNMXzua/9hDvFJ1VUHzUW97q+Dwf/pe6CpS
vNsTJlq7qBemjUcJdRknD1KcogVDmxxsQUARuPrxipJP55sJJzVEl5S6J11s0CUI
UA5eU/Q60PKUWA5ZYWpP72Sf0vV5oobzIVby1yi5zL5uptSPIWoKWbzYLzTmjMac
A3oKXyBZUKb3MH0TF9NZC+l2gQ+tgxDsZbzmZL/yQUdxw9YUs7jZzyABe4GZIYDC
YtYlDGeTGWB4nvHdF+iF5lz67TpslqejigDNXDF4gWb62Pvi1Bveo81gcSgJDg3s
UT9vU4ZrGh0rMltvfDM9SRzDXzCNR/Sjzf5oDq6XfuG9N3p9Pp5dZWl9w8vBH0Dy
oL9d/hc6SmJlbGoeOqrMmOjsRruRJimgK7Bm17rgiy2K5frtDSBwhR6/njcO1wKV
KA0QF8GkRTINYH6jQWqduZlEbzO5ZKAsjYirh6J5yi8VODkG6zskwaz/OQm3nyP5
2L1/Lsg8/JYj7rC35uUqGGx2XhSSJ7IQ/o1KJ1oL41pg5kzkuQzW/80iPpU2661C
fhTOeZQgZQYpClvspRfHuahEzhW5GtSOchbdPDNOYnHb5bUo3dLFGG604JaMvuIY
zkLu63uiHX+xMBkwFCoQsGMEWAfGgWSvBCymZs/ih2Bz9EZtzpSOlcbD4ljT455O
8sCuAqmuFvIjFQApYOD+hIg5+gMFDiTt6eNERx7AXV/Gi9UFo9O5+iA0gXvfY74C
osU2jqQeOzszQTeIIAs3E70KIwpWdEx2WHP5tfs6cfw2uaabls5gVpCML6WL/a3A
7rHAy8/ezEuhXB286rWe9O1HgdBHLlue8wNAegTFuAXI4gKOI9MyVzs31wH/1/CF
w7ItVIg7FA7DH9RHOFA5jBMHdl5PVrQaj50/EICQqVprf7iEXZwYX0zdQZqB9Zkj
XJok8otQG+Gh8OaNvQKRWkFeaJSOjbdt0M9FgbvMAuWtOU47jiW09HXi52QHNa0D
wzUxTmJqbw81thKGMBXazl2n2EvJFuWNhOhyL6D6go2My4YqgugwS6gtDOqo2rx+
rOtTJw+WKDMHgpajTR1YSlkP2eb2ocXQzs9wt3aC3lBGFHubVh+8vABNjuar/Drk
+vP4imeEQckHHo8lAKi/N0jXgosABTrMF/9vVPu2hj/NdyjoHCJJG2vTYwt2S/gw
lL9tP1bNwa3uTnhuD2jT0AXXKXpp6HwHM0AUMVdmqjZGNPQjjdY0rDxjuD74P4Ij
6RGqLi/nG3APWYUisVp2N0RNulMPOUoGLw1Hqrg1KFU3E0PYnE5+ajKGP+7zFkE7
QNx9Fcc7bo6p82RplEYc4gesw8mJCtJjnouHXbYFo1O0WtHbNgjHCFYK3uQT+YdV
KVQ/3z71i6yBfII+qB8uTS5gicyVhMkczTOdGmt4zsNg33+Y0lObq8hXdm1lAnnI
FB1hwBb1lOLOA5XO70rot4L5sqJONZ3o+t+TNqhk2/NuNcy7Cplw9ZmIObGNTpYU
gJ58UQy0kcuf59rsHbcep38qKYyghlTYYjay+Dbj69l71KZFe/e8sAFjygY2fjLD
o4APEShCh4PvJ9RCYt57s1iA7zY/KWxIG3RDDJ57TfG8Me1SJXdwrLLb0mbdmZ7w
1jgjm246LPHUoHgqpfyxr4mjt55n7thGBgAVzx8rXNRSNtjIagVxT0ZA+P61jTP0
q6V45HXnfe0sQYiGcxw7Mv0LrvamppRQEZarTb+E/WjLDTxEO0RLnWOqeQZnFtIm
Ikh4uUelPj0qC2zE+JuTqH/zqenu6hV0PmoG4EgAOpA8Livx2Jde+dqPCK5HTbbk
+09eaHvSQRayhu+u5tVqx1KjLZQ0ICWW6eieRLDWhsfEAVGOKk/geWBfsJHeU8//
a8vwrBxcJmBb97cMp2QdJREoNyvctU5aqAC13NvcK6Bnvn9fdRQzd8tNewMb2IE5
xc3al+qDaM7FQmcDCev73c2x5KCwMacExiTLwto0bl7IMFPGGTY7LrURA5H7JyAG
uBgNCzmTGUW1Q3dU99zByzEDzsIHo+1KjljCxDOOCX4+JKQb/zSGexg9JdNGSs7r
ud6OYwx6G3y+2PvQCvqYqYgYLU3mWHvmk4BodITzemIHaYQPg2b3quhjTnLBpX+V
CaB9AKgRz31yKDp+sdtNQkh9pvPQNwGL+/Pj4z2aRSa4vPCJW4rpMeFMn6khihB8
ruRsPV8r1dpmiWXFaM0mgawm/xI0Ir8EIJXS2G8It8NwUVaNApe9ftiM4ht4fx/E
BMPc4fZcO+SuMXhbpOavBux1aJta1yquyKrIOTQGNVFTkciKMrMSs2GFP2+LxRal
T/mtz+ZzwteEWUbdgynmK1djxePdbtE9sqIZ+IMOjQ5kSCIJlafbGZ9ssk1BWQy9
Hs1UZsDj6K3FZghzmZxd5KTpj6jpRuQAvF0a9gXBa5YRG8HlxNY8XcRK4rDzgaaM
s5vPd6ZNe7KSKYpQsE902yqpfFwBfHGVuLCP16Usl4cG9lhbxYKz+eNTeYVAcj58
uTWrQQAH3SwQc63P9bfHuDL0Yc0C6GMMQf2LXQcGBjh2F+FYpgMHKQtxNqPBNKFH
F0u4EjeSBmkVSHwqv918CJinp5SgVtRE/uEglbIETe/N2jKuRqYbLv7cJejTP9t6
O8KYdx2J3DZbLuZfgmohYRyrw0bIDF1bSfCEPDyQwSfzhBIVkRdkXQHyQaXqfBqe
FeY1EJr1wTsrdMacGYdJCJ6OtJVYPUB1JTS5Zz/5o1zBCTwgffRIfjZ8uM+aUTdZ
3xmYpfBT1gh60V/UzKxYDeDNsE4PlVjiMRSVf3dX9vfvQHRM+CXr0HGJqMy2uXA8
EfW4IZHR6O64M5d6/RyuOOowBWwQFNmq4y0oHTGSQ/+zK3aW4EXK5ykbgGwj5VPr
KMzHtoZqB952tvB/VNpgN6O+yce7ix89ZcH00N3/yPWDQhciZDhq6OSQto4iXahm
7EmMk5DZMkrGeE3XX9X/RyQu9DovVe321mQHlJD0GStwLvJW04p4a2LfNJ8sndtS
92CJUbjQYipppWXulX31amHCVilaXS6TlOz8GZwxJCgiKUUofYaJxAVh3wSOYhmF
tajhZOJAg5On8PBTT/hjHStMh3ZldRasLiWncb/c2MFnxOvYIzQiP4SFKVJtPBH/
UUUqYhwNgqZp1HTiVvy0Rjct5rzgljswqrDW/Gt18xA05JgLXrFqLYncQxABqjCp
osc+b/WfoYD5tLvEdOHXDOnrwKvcTgPlGK+mIhCD5Ev4OQkbSq5+GuxSNEQEDBoi
dz8A086RQUPT4ZsL55LuUuOBEYv0i6sOvWGO20+55yZXBOxhgW7DDufMj9Nn7CnC
sSm8HPQI11RWfMN+N4qo+PNzuKOaapGMnaYvq0guICUft6+5pSg5prCr4Lc7f8q7
jIaGHkk98OuogOltBJwgP5O7xE/OPmXON1XTXJ51hsPtrwr4tWY73ZbcV5BxXdNT
km1YBOEPDVAgqqSX64LKLnehz7oa/O2+/2I7RGF0fM6HKQXcI5kdqceaQOUhjiaM
P+d1/H8jBOp/oE3fd/IgxeBlbDgCrcMrclOanODVSlwYvr86mHTVgJjCvPrZ8vsB
mAOvI0obGY27dxzgOMDwiUvIdjrGnvSooMiZ0OvJCF25c9Yrt7MX6qq3K6rTtcnN
GTH7LmiVILfbuxYsC4jusWqOuQvsvMeMXsYYBxf1v+goPvjz/06gO5FlDAxtX4XZ
9G6UckFpaCl8YoAu8ud+Q2NrquoHZ0hlS0ynA2pL3RQLkPsQkgPL5uo3s/9QVtFY
4mQ+kwE82VMhD+8nN5JjHgqOLoqSqi85u1rL2xyqzihYwudoSayTF9xd1pjeTi9B
/o0rTUjdJ+dB93Y7WjfdsH3JhTPUubTtIQpxKsad8RgiUr4W6CEsAEQkHrjszv/F
UvJAepf/TGgUKo1inisyW8Nc4m9cy8wjrJL1d8BeaQfi5hd8Q+TXD8d9ZDr+9Dww
Zri9c8li2LPbssmqKeNFTWVwdLGGhB8Hg6V2cA4fD5tV3BX0/vh8ycnPrNd1K0de
4u2N5+NKKMcbDvsYsIRr4F61YDwTBwssRybuLKesUxNJ3IP+o+gIjAXrRwrpVnw6
WO2RNdbLc3pn/V/7o+WrosflRCFqLjaTmqTceRWdv4b920Ysdtbory4zieEySgsn
QfywNVIuvmYkBg5F51cswnbcw5R/YLn79NoqeTWVcTjtnjzGKWxD6sadF6UN8wFa
J2eaAbb+WQxNYXemXQtHtYHRSJC/755cH19nXXveyth0ZNUDG+RgQ8jZd81UFEvJ
4okm1HfdU+Be1VCwKhoh5b2EYQZ+FamKp80OfqcDUHiz5FKdZETS0Gsybucw9Lve
1Xfw0QV6WmB01t7V9oT9qqkBNBlfGwIhKnbwQzxcOXhymVsSDGp8ELDTB/IXB1EN
6V2//oDYQUcRyNujajbXNbggobGqABRNjNkg+V/fvqzbbkjNy3orQCtySRRvfsIe
kYFBcW375qRxJ6AC/3ro/4pMkT02zp5PQdXPkxdNEUG8o2Sz2afkNHeAdJmQyZPT
VaCvU5clMJoWXDCBBEjLrJaEGSpqB4Fddp0LwLlUsvkpsGfP3To1XLuBjdh5d/Dx
/rNA5fT/c6sw3V5S2Rfy/jIZaycHC6K+kN9aEU2eNzTBaM1Nd+LaAXmiLCrll2sp
TxobMFZ5L24B/Nkp1gLMFlmjsupBCaBfy+Em+W52cOVOmxmeE73T7GBTvcVkIpDQ
7bjFcxb7Q24nyU2UmxnSQUIoFtWS/3POiS9pdJyzo7LzbiPvSiTMCtqUGGTY6inv
ED7XBSKGKQldNQtpjBUemrI/MPsPJCCD1H+0fNnpzn8x3prZ3saoHzXVh5nXeL9c
+5ziC8reiMVggi4HdJCRzLoWbBjaGmFizbO163X+LtMEjXXKBd7AgfD3b1SV73Po
jv/eeSRvDy0+7GhIJ/DnQpwf5BWzzSEgCpuRGYO8Ax+6JZxEApIToDJ2eEamQpTG
TAojqpH4QV+sFKChdta+0Ndg8onC+fMRVHTjo1DgutuFs2h+4gIiVgOBWbt2Y9wd
3qj7zfLcj6QDpufuy/ziXHtvqwUeXlDQpqqMsDuwGFET4+rTnHnMTV6a/u51qejR
L/QhWxEBbImi1iRJ0OtdAEhkUGfaCcaFukwOX1Npzs1V2AW1VHkJ+4kKFYPvPNxU
Z2V1WhKfoc6lv+pUzSpHiqZlWPDaN3xSAcrZX0oW2GqTQQzfCopqPdbM4+3D+wBj
JDsm/f7uwBYj0Xcd1plZnd8xPZIRAUhdEgH4WT5wjIcTCfSrT20Ex9Ih38z3r+nf
P1EqLTp50NRsFCJPg5dZzPEBK4ZZUf9QEv3LA33uylRC8rgAL7MbjdJEi+Un84k1
dbGQQ3Q36L8KuaO1JH8a32Jby5JVUV9SuLiDZKSTk9JP6T1eyfglOX5AjKNQ/0n1
W/wdxEOnRoqkohXjKgPZv5G1ADaRpXOJsAGH+Sjbg1dWG7sNH4MvB6GwXqFP5who
oX2Ci5cR3TTcxzbwt/102NkcVP1w2glBmSnWseImfSrR0bXtxhLq+VVyc7PUsyGR
s1C6fYfv69Oti1PzwiuELOzf7cBDOWzVVIQGT+l7jDuRmuyqnL0N2PeSGs5xuMKJ
2v4xqyQBAMUKb+B2b90DaxCu/uaqGd/JgASXMuCmM7jmsUDy/hmrG52rynb+6qeA
vsaMIX25jMgmPRJnbZE++ApHhjBvI/y8tFr5HdYso+Ub9+byU9KbbOqMka7EfQX2
dpnRdgJT9R+mjVrHf2fVQTG5t2dbavk8ukGDXMHAlbm8NyTzMluL8JbekftvVwAe
nq/3y7QqbCCnawKDvzuzpo9y33Gm8A1UzEMHTxB+zjJ6/CigGya6T/twIJk8wHYg
ycGkroxSwvHuuBz/B1fTLw2ZiPtsr7ZZ7GeVW1hjvOvnm/6tWmKmwO8xAROzY0cX
gePX/B2hEW4Gkr9jrW2ywh6jZL2uX7jMAmXeS9mRvZ4BFcNm/znxDhF+D9zHrXbm
PIk9wVHerFirdJ1zAwjPIOaVjwQR5qxHsG/YWzRecCwKJcWvbsYXWuQfBKC6blRL
9i2sGqmEeI2I2IRtVxR8d3+MwhEWAIdfZERr4IofOSd8ABg3zD7yWe0et7PP283t
SNY/3+R38OBJjRbddfyqDX7kf/mufxlme0fU4l99uo37is/Dea0T8InqFrH+Oxd8
hPBsoUbqRb10bJSbEulJ7dy8kUikIj1diP2xQLSj8e4SA7lunr1vMhrIOo809YG3
yukz6wNkNhfaEYNW6lGLbl9A6OBCtyjQQXOM+RgmRFo0JQGsUCvMiH7p5h0zUg4P
9dVppUArJlf0Iz1M3YBAvbDu91y/jur11wWidVzisiFIaLmLQbWRShgX5/KRjw/u
LQHWubVcgtJg1pKtXSwQtB03iamqRf5i7vWMOzrHhIoZhZ2AiuueO71AeUPxErvn
Wi3fDDCgQC9Kl5NTVuwrsn1bVN/x4+soOOlnvuS2Q8uettVaQqTpSk1Z09QgKl4b
wFjZsVYebJXNxp7n7BkNqY3Dh1QViZr7nEwP34SB4evA+hwIjhwQT+0t4C5DpgQ1
DacbS7LZquw4/Gs18d4pyEMbh872ibWIM4QYjIhIz8FSfiEevs3MpISxMjZolOJy
zNVKr+ZtyPHbj3MHRZSj4PGwgXfLxSvM1sDcpvjOv9w3d4itp+zjIEt7TlYv14Gq
4l6/kySd/WVYeWcBPMEC1W5xJauHT3E7h614NZ4EjaWPX5WG/DQeLvgc7yxueTW9
wsgRMxAFMKh4TdMmDPXRRG8W1VoIeKU7WSpd3FJGCQyRYYUeHTZhjVVztz41aCXp
8wnuujpzhxVfNT/MJPkbcR9RL/IpXmByTaCjXMyElo9/95ImRR5NTMUiyRJBObRK
hSH2RVUWKzB+Z7XMBgifMIv3sEMNuXw7oHEN0DSdlY5y+kIWG3Zk++Hn++B+2hfa
+IhuDe+aaeD3G9xJ+TzctguhwOWHV15/UKdJWBhd3IL7LPJlTpS0YZlyy49KtB0R
B86zrMl4HBzmU1fRLcnxUsWd8uRrdS9J4iA1onaPuU5DG73VGSJnWpN/89eMgsIM
YVHA3JDcGtesWjD3R8/ElRIf+TOU54cRKr/evHlrkhNSjP94Lve/uX76OZtLfRGw
bLi+VhK7oZlB2v+0o2mYMscpOobvebyAM0+I0g6ZUM00muDqmRWkoeyCZM2+3ctB
mlui00mJFjw59xlEiFAAEwGSmqm/d+W0Z2Eyfe7Rakx+PqIvWL0urlP7jfC5gp9V
FZUTePKoNfkcJBrMcn1Pg5TfPRg9YzV+YPbnFScpN3VMIfQfyVS58vAwfWTL5cL6
5J20OQVLpeS62mpZ9tLbK+++Mh6FZkfo+re8dqq7n+YgeXWEby4y6b5Mv48BLlEC
xDvB5EU8vT3hbvloNJTV8vYccWjdfj44P8hqckndaWWiHlGa2qvnE5p6zDixAnko
cxKG/aF/4hk66WlLjqXARiKc6iLulw0Dq2ipnzPoIrL0JyPjQo4k3k+QpltUmB6T
QQxFReEygKQsdQykLG/ERDTXI+qmFLgli2h3SUXaOH+BMjjgbt45tiH9mifiT+hb
uYuGCSzIFJ9xNRVv+Dam1NTn3aCrrJAoQogi+gsA+3lwjIhDPSwgThLp2GGgtMsf
PWGkZbUOE1zTswpdLDUvj6mUqhDvu2WXi+PstYeQukYa0sNNt9jdourNF64JFijd
zFYBfq+6w2lySB+xilZJjGqBUPOGdAXS3BDfz5Siawz8kr7+y7+SFJmYOplsbAG8
ycblCMnGvJPCDS6h10V4kb8Cq7h+O05VyODOm4WLa1xeg2vP7jVrSvtKozOqpITw
4MQNFQsEK/BiSbQY5nPY5DeIWWM5BZDrikgusiYVYM3IbGOWYbUx28gjIvNG9RJr
gxsyW5jomSbZoBuU8Ho6SNRDvAmg3TFbq93ZEbV7AuUsvI/gV5De/TZU6FUVA09D
WbyI2R+OBKYF5y6HhEeGY3/VytdGAzIvZWslaNDp76EjElUSzik+h7EJ43IJr5rE
iqx18X726+Q/YfT9HyadgrI7GadSBLrGj2C7JFkc4ubFylaP5q77TQpqSlo97Oiq
mAmsJSyBsq5FoURP1+qfiK2m2D0rsmjGSvE1u3YH0Ftca770ZOydczMl1jNOXCSj
2/lzpXX5IkZwZrBKYABaKnXjQMuV3PFB2BBdmluIQlMQEQytYUxWfoEdoAcxYH9V
LnCQLl7x+ZbbDB4+mpTmjENmNm6hfxXSOw2aok3rLkBvnrOg3/px4+Eyzf94x6ch
pS769GK+RQ+pgpw7iF6EbK5X4Y2irCnVvGOv89MGT1dqORYfmkFbiDWGOELoUXAi
zSERGx1QoOGi2bacd/W8/0yE5/gL+h7P9og5AZQWHQHqwvoZ7RaNgU85zrOcUZ+b
D/uyEDN3z2hATMn2YZLusXcPsnlA+ubZ9vodV2dsRjkMukWbf61HDrA9F/RfIp0G
nmdCcs+BS+4hMYMukVchqlp/TveLSlVwzIF5p7kkCSswxV26Ph1lrCvmbnBMZsVh
NldDYrwRLUpz1SUDxja8fjwfsi0CsQ9d1YV6lcZrZfK0tg8C1ICku+3qr7TEnKXF
f+evnx/s0XX266j5lciclt7hdqOKzUPFTvhKXgNEHXUt621NkmTeGhnmJLrTkiXn
1y7f0zpLve5iO0kH17vBX3g74rXlC9OyY5H3gKr4gFpM3AGMOe0JKLPFHusa6BWD
961W+QAZMGaYcf9BBTTOqiImTw1J+XHhbnm5BSP/lXMn4DV2PUfypoPMkTbcwbPi
LJB6NYgDCdviSFy9PlJn7RCWOAG3FCMIG6Wn4dQk9XIXnHccg68XJGc3dj/tegmE
AGxrvRWATH6lCYKh+bCD12VUm/i2wzxOT2X7kS5gfssX1vjzRQ/O/G5KpCtTYJ9W
rzyLoVcmOwhb1fUcOqGVrhQU9eQucL5Y2qJCkJMVviGita+Orz2LTvPS/SB6yLkJ
YslFMPNqLCaXbvPcRcJQXkaA2u+Sa25RxcIEnFMZIbsZODC2SNDt+tu3Y0qjD85R
Ij3YFBCqJD/ERVaeS+yJoK+4eLmnnWLtNzUeV3xy5/K7HqnlpXADHHkj2oR0sLnP
Pi8mcVPDf1J3dX29o9KOqR5iUhafoPuziSi4aSgH0PYi/R1itCcE35WKrsKFegse
UeHpow7jnxF65Zzpz3PPydQysHqNJaiKukMUENZv1R2oKnAAO7ljIkZfQ+hjEjjS
9pqOCT45VVNERyDAU1jUUZVM3t0d4jZapW9ze76Z4AX9iPzh6ULWxRjHPC49MZaD
v9eWa+tfd2SQ+u61PqV18PsHBK9MZ/tFSwGzzoXm+V7EPQNwxw+AJ/uZHOmi5q9W
eTKZV7v/IiO7HYozwI1FKHXXYJRsPYOPz2zqUEXfz6QohC3FPj4HibInoaQPGZTu
E/f4wrr/Gx5OL7fARs6QxfnZETlMUx96Ky80JqU0DyQCnRR4bZ6AGM1lwOT89jts
JSoKmGN996pE0v6igu+xUwe7oGrwds3wxknoxm9MZDTBHuCL+CWHmOmDlFliOZbx
JL7Lgutd69AZGeUli0PgCdxOSuCcVWiAn8783gsDTHMWiBHOsGwvcDvcLc+YKPOv
USUgdMqueYEsgiowOIXxccUTkJpv1jtZLuaLy1drUswe9NfVhotaEOHDOHn995BI
rOTiOpE+A7MBt7EZ9EORFEUafRd97UGNaI3YIDvcWzmEVdc1tjCjL0/Tl1mxNXiy
3HnZr6gDKMGrGXLcb2/X+59OotNCbQGKWmKSoBLTGfsHYvuc9lcpZuVOPTF/q8MC
Z+ha59TH/+9eXU8hIEHXIqT4dXvf4dvwlD2tDMWJDlltfhMkXKgo2ehK+ddk4vVQ
5Ql/kIYA8RDrPI6sKkCe0PdFZfWvfkaVvZ8sHiWBVqynnp1l180GJ6pmZ01BL/Wa
jGQDrxReZXEuCi6i7ROI9FVNQw2/6iAzGqaUU5VFqn2fM/gYnSxE0Q7y+g0B58eT
gQ8whYc+cxFrlD9O1ym3azDGmn/Cpqu5AAccXM0D49QLPaX3kelbwsyjwX3vj9q0
DScUzBo7kBR4cYp0IJRPnIiw6ZQdFZedPLfMqt9ZOBm9TyHGaj5YliPxhvNk3Pzz
dzpktudlKHgMkq0WeOkkvTzlDYSd3pL/Kfh/CeHyt8GgNtsZLgYJAC4RD7wxjHc7
u1tGPU5DTv4OwBF3U80rwl3OZPgmTJcr82Bqly3s/I+b/6ixBlMTpI04q7MsJK98
lSRF93bBrOBsVOALz73hnF1P2oZfoJ10c6ojFGNCewT+wEI2BVCZfA++i1AzZacY
eVAqYFrnZX84Zjm9haNSlZ3gSWqtcbCox1j1rWTVRXxorn1TPTEk/6FElMjqvHBM
i4pxaJE1D+zB0Nj4hcGHp/bXhcvrrZcuFHyPD3RW5avc2y7r6w5AFf10yBoR1+Pa
Lv90QuYOq2anGhtV9qlpVTk2iKiQK700g+0Sdpt+/BiGnozm5A04Cq+9iIem+5+2
MSd7haMOb8vi/WHhGWTKc6KUtMs6VJJ3/vxsKgiMLqEuh7GqNwp1YOX9OpJ2DHIC
f3Od/y1TLNIbRqW1h5WeTeob5HraUZ4xelsCiZh8i3X/o7UIwXbHiE8vZCUv9NDF
T6RwVbsAvS2izC7VPRRlETjZJDNwN2doKXsDF30+fYtfP+A/a/1uwRDlEjDX2dUl
8kpSpjLUcnAnOnhiv41OvbfNFiIdR4w8DptEAWvFBGu6Z24EQQg8eflYixDegV3e
B4vse5Uu9/RYMvsqExwu3lZGhqIR9uo5dXaWysFeF+RvGN55r68Bor4+ia9/CO+G
6JleDeC/dbfNbpqJtp0+lg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ZGSzISojspNjyvu90QrjT0UIQDcZhzcxaYXM22odoCaqQcAl4USBM73rdqI0US8c
mYjBhhRJi/L9c5tF1GKyxXsOwpNu4m7nT2CQAHn22z01gqvo0jH9vMPUwEfQR5ZR
K5fBSq6fykyJE5lHQgLJnQ/+jYCP78+TO6AALpUrMMLQ535M+TNaSfmuQEl/wly8
6GysnB3X/cexf7xC/onWNhJGJsaa9BpFiIouh0NfVhHuszqnVHsHVjzYtbf/lvvG
nKxeJOL30H98Yia3OU0/GvNtjX+IGJCp9dPCCEliCLjPWUccfdgdQq5n1SEg7pmV
rS1L9G530/IcArCypx4cdg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
w0ZR4ZghBxgBRroyeB4Paej9kTplf1WMCVOjSs1gmm1M5wAfPOFHIpT5J/gCZ+SY
sZR31gk/ASNDRsuKaeIZ7sQ6LU4Oq9hWH0rGMAyDWyJivUsUcFro4z5jtAqHkp/y
dFk36kK4p6AElEEqV7wuDm1C14sFgM0CRRgOehYcZqslAGwCjnnE3BRJu5UlE02v
C3jPhiZKXt3/m57Ggl9u2yVrGc5eYQE+mHXZnOoHZzwWEskAtYn5H6AVmTMIzHNQ
JkN1kxcNJQq2I32q8LjV1tYUbf0hxWFcUsr05P5b/VDiDIQlJWZCqxgdmWaXPQLg
HliYIvtsjCf/CZt8sabTvoZPxq6Ex7YQDQFJ41M7APKMhx0RHzW18eRkyJ3uc7/S
u/XTgbJlvIJHyQn0TY65X7op5WSyO2bjgD8wbFxd8mk7SsXErH3LwAplcSLz8YZ/
U0Z9nzRLsZy248YseMHaitgj7JGl4Unl1fgZ1ik2Xr2Xn1Fl00jggFpb2jBev3Z3
g48LpjhPWGOr+qtPSHxtowikaYhR6vXV0sGCN6V7iNfsWq15wNqkFbHVs2m4Jr3R
AMyKv2g7Wa/7EKlghItnFmFZl/RH2/9iWARidsdYwXl52Y8VyChlEDnQTVZ4ZGU1
gKNS2RvnA/PXYb9LAwkvJbEGPT7vo6erb9nuflYhUcAQHk+gKMUnbEhqY/UcF8gm
TnIChYLSnLLKgMSgNVkaVKp2XEvbM4+el6v9dtHasi4sG2zRpXi9aZHutNEAtu+y
07msz9ibpwlDlrFOAAXyCXBBFturo8JhmveijmlflVxYvDNwyBwEDT2z8nDEG2v2
6zWYtAK9ipZhT8cGxjTq9ySN2mmkAXHD3yEIkc8Ab0KKIT5O+sPZq9SZqUTu61KZ
Zt69MKSZeZQhdzImklhrhwMhyqBZT2WrFYqbYEmuG1m1S94NMwXpBMiGFjBU8pby
nnDTbzdP1zoEhHIzjmk88QTZQLVPW6LdpODtiyhZFMDQu4rfgzt8WL2JqLJ46WKZ
JAuTH5+Ea2ri4k7YaM5snDgZUjBL8weWxh3rWqk3/FTlGkILkHQhWKSIesFBn8xf
NnIJzvqPq8pXMtI7BJk6awtEIGFyc0xeJjBe6WzbA73zBysNeI4PSAaANgLone5v
XV+uWDYf/++s9tUvK1Hz1BCurbj9ZdQbDNBWBTAO88JqVbvuvh5fS9r8PuU2eLCb
JuoFbt3smqCZCYkApgzGorEnKxSNNiblTv60waL/TsSEGodObucB3P4jTH7KOozE
/7dsubOpuZ/7hBUuuEBArW6kPW/N+rW9lkqCZfhhSoawE4KfJXYc4Dxb3QtiJwx+
ILzvrWyOpT+jPhI5Vn6N6e18hMS0PC0Kdelhn0MUUiH05uBIyzYDtwjuYpbJ8wXm
FqPpPGIS+RMt5PLyWfQklAZzwtaj+vMgmRqjOIIH8GZ7EAqfbijhB/UlVnl9htaK
PYTuvpJEuGHJLLrTtm0UP4Yc7c9LmOBDwlvCJhoNIZIpl5L1sgrDJqSz05GJbMa9
4tj0pGgog4anaPVhF7cySz2OA21PswUMxlqjXGBNCjvqyBWMGr9UrGdeD+KwC2zp
gJhEyHPIp4bMtfAO9KltLuIaHLtw8J1OoXNYJLL5OwlY4O9j8pxapgyIX0L5Hv21
QrqUyvc515S6yLSQm0CPtN7Hu3nM5NKuzZN7HdGB6UAQKusg5bB5VsEvc0QyMKWg
Fh0fGatyhG9/uhv/OJa3hcVr16VwUvTpAPWoZvbt8fRj1WiqYiw7aLk9a8ioLDW4
wFvDI2+XdaV3DtYRk8qbtvGjxGHiY2UBjlNlziRh82aHaDXPd5l1PEcOjzIcePA7
Z65lHK3/TXowI4eqpGBB+/lAKL/VaeYT9pc2/8KcPMLukjThkQwQ3gbl2b8ZTnro
7sPpodjJmSMasCA+jmiMQL8MIW/PsPg40v2+zvypUEDkSdb87fA3YttfpNTCpjzd
fAVU+ow5wR/YVZLP6Xk9DkdbUtNqG3s5/5eiCluz/fTLl3OmuXTxkuEwuv2nIn5c
wxw/0aHMUZ7lQtl8IWrYXkQqCFXafTyJS4yKRNQqinnx5h9Hqo2b4lBvJekWVnLl
Ag7bjJ9oF23EKfjGbJXWiXHteWxQGQA+yHWINq/IwLDlSJAvFyQJRLi5jh2eoFhl
3GfwA7o5McxMJXgiSlfucWLc4TrCvYarYnq0ZLHt+gBNyqlL91SVV60l0QexzpEq
kZtOnGSqgHiyWBAAqKiI+72aZLQUVioKOxAo5hCXSWi1kyRJrIPedtAhOfi+ugPU
1eIFb3tD19KWOiz8y1/nxw6VacMlmEO3nMbHI19O6hwWBDu1pcvrClw1qqyawuuO
oqIpSe+n2U7qjFNF68vFJjWjltiqwT53EgbYwHlMh2fUotE78h64eiaCtBbFdAp0
h1yTnJ0c6jAiXHecvzZhFxxBu1ydkzEt6cSen/2icPJPs83IKENnyDKSFfPLG4GC
ocxAUxkUl7lRisCwmnB9eTepeiWVGIBM3NFtyjvJL9uQSUur6GqKppafiB+pkEW5
dnYHfLCzA5HEa6CAcN+UdJFGJd+2aZ17dUpGLubzCIyQ7t8ZvIIfr/TXtt9ErKJJ
JzcBwHzxDT82nydErXAz5s11WYB/nOiGKA/MxSIBB+HNE6JyWWV/8EUZVZPjDhgQ
hhRUPpP2wh5O5IMjz4dnCbcJAdIV7Qsxq4AazTUQeACyEWOA2Cl/Wil1Qp9hg/Vd
t91PiGEFg/BpJ6rrPHngeEIMtSPCInmRpUypxHPnx4p+ykfLpKRy8Am24uMYt3/V
UP9HhqGO3UMRk1lyFw4uS/sVzS3O/gfIzuXJ+60/WDuJwox3LCK5+v4PMiYpqEup
c3U6zY5NXX4pO1eS6wL2nJwyThhg3rKzSKOyKEQ+OzOqJn2SoYuUcPqst9+Uc4dF
AXwIqktSVSecC0keCxwvxcI+EXKe4hxfFIQXapZg2WRYVoc7Tp8cT5XfN6jpKlsE
ML+rTqY0IQPAzVBCYKDvw2JonWMeQulzMct/BRuo1nDn7AM0qB3n0z1VD5VtYie5
vexU/yuooj+NQUOeIHDZOyh1eVG1JB7BpzjkvHCkQ+z7yK90mqHFU6WxojDLxh4R
Jroip/JrEtDF/BXFByG2UNNywyTlR9bInYUs75n4Ef4Ok412norD8+rB/PbtRIx7
gNYrtKjRzifEnVH0c+VenNnbdum8qG3grocLOZ3s4p6Hr8FxGgqYNTAEImwa+zMD
DY/o0J1Ez/pwrWhT+Cm57tyyhYoFNvs6IikOTE6P2ulIQqS4zl4L3XH99z4qKOoJ
MPABzeMtq84k74Qmg+iP5mdrxtWUNFloWCXZ9cqrY/HJbctxz0kyc40fNLMjcXjU
OSFSHpM59PydkNYowx+Y8M5obFNAjcGfpUd4rCRN3vu/98ebYl9YGxRJjk3R7Ok0
aIOO/7fcJQRiyqli1Ez0+yZGR7FpShEAJNFxIVmyLwJ1MOooSs8riaWAE84rXYkb
27AoI2s8frpVdQHr5Qsl0clY4/mdiSpOT14KDTjH80aTE5WQOtusrTwnq4c8pfqZ
PJqWSy9YgabAadyUjDasNvDV5o79j8oqr8DT5jelfAqgOqXwjh+idHrKtwp+oL2D
pDDH+2/Wsk/cdMmySE1aBA06B2Q9Vou/13Gzg6pLj9JL+I3AfZV1KN9krPX3inIA
CZ/+B/B+lpuPeB/3LBbxek7TjgErnA268HYCNJMrAYjXOd2f2J1NZtmljn1W6GHK
fzWk+FP9gAMH41taq4T1ppsKvWniCIXzueX8BWiPulirioOlbsGXZTbjUe0YykRZ
RQ/MDZizrMTfhWTgrn9LPu/3afPPcX/vnI6wjG6baeCYENTODeiBm1v1L8Q18HD+
WWcQ0tbtjRcI/7/Fll47w2BbFTsEz1dLC4kI0H7sXvwaa1oSoIVX2nRAhGxbWbiu
q3obdYkAVYyCmuzY4N3R4aoh9FQNtX2nc9rSqdjnHeklNcmEoQiy6FteFy2agsjG
ZYCtUvhi0xJXZIeBKnRSs/ofX6YxRxookp+cpnbtCo6QD86rwDV2/ymeDfKu3Ssp
nX7Ke18w+cvOGLp7xJcnnKlebxUJ+hDl3N13xx/Gxk9x0UaUDn3iN0Sha+PuGGdg
FyCXLvizTpKRqk4dSVKPJ0ieyOMv7jCvqg770AYTdKkE6KJ8noKI2Z40ndO9gLUo
qbI7gYBDnNJf0FCk0FD8eI/OK9mn7ySM3xQEjktnEX+4KZC7SCNGK0SSUsnaLmNj
EbT2QvN6mmdv7iWXpWOd7wCXvwUO4yMs6DqhXdwx1gIMVfeG22gpZ+bXlZhN5GAn
RMjTdBgNVCEQ9aG4LeELNFb0kftUVMKpQqvpLkzzzBYtZAztb/LQfr7AAKelTgV1
pNLu9/Or1aAVOLha+VXaFh1kklzt7U4/m9VQxkM/cYZOqvDrDbTdv7bsGx60u1ai
T1z+T5g58IdTvFEJv/s9MpvdbL6SlE9a4yWXro3mKmvv+pSGFOre/Ok02lMMSML5
yHDvpefBovdidEXkvAOI7lF49//hoyJrGeqUwOWOo/yPTLy1YxhFEP67bad0hffc
2NmAA1+sAYRLlMDdl7zOXMrQKCZ/JJgUn+QKIcU/LIcMxHQC0ENGXeu+uM6O4gL2
iVjvieEJwxpB+DYd1oG2Pl47d+1PqDR1P6mcIo26q0UXNU9NJdfZux7Y6mK9tsJN
XfkqvTd2ILdgV9nxRSBNBSpihJC7Gpg5a6VfM0FM/BY5ABExysiS3pfDMMJI5IYx
egVotDINyjaym1olvqdUAK5Kh6mWi4fSskO5k8Lu1kehN663BM8fwzztYW+2zwUn
yEpHhAt1DuvyFJczdlik5UZh5Su43fl3DeURJ3Uznd2CKQAgouVlau2ypgi87cPI
wdJGvJzy9UFuhDwZhg4kz0Q7wpGJ/E6OBX1MGJCM5ZsZ+Ipnk2eGzLkIrPquKzSY
HP9xbD9IFjySAAmIROTFUw+/voOgWAsopywhdWfM3t4aWYbOtHR1DApkk76j3YiH
XpHatUj9/Xy5uLLQYx872ftL1wQgL+E/sOsohDjP89tYX78H48M/gsLHTxX+Itkf
vWhR+NjR4SJ9b5GS0Dv2adr7DS59tp9ibRAUgnOoIydkt0HQkMhl4PAV3JToOy47
03C86D6AX9ZyKDYyBOzckooY3X8HY5DO87TT6BCtC2Kl7Ql7tD3DgOj9/OAZep53
13HiRHUoU5h3OVEahwBQpRP/rqSRKgD+oo7HSwJ7diw+Q9T5dHBRTBlnNuDeGINu
/+Cjr9xjto+ojnM7NeS1jC07VIZkJf7fOLVvWuOU4WesN9yqYEmS+nhar4eAc3W9
BcgbnlVfkEZ1/mGfSG4jharx5bLEhll3JHQ3dtfbGlGJXl6WjSPiANppTGaK14qX
CRXtba7XaL9DE9gNhihnNz1q/hnpuSSxca6RuasZmrKjwc5EiXKe3fd6CPFvbLCY
oiIAGiT3V/Zo6yONCnV5l3s0Zlq45FNNf7qhGx+ere4Nd83c0vF02cYgrqZ1NTup
CJY1UImaeGk/Uc2/kfgHFDA+PB4BTpLjEwIEUW7NAbA4Hme7d2KqmltG9DU3TeNx
GibpiajY9E7sZlMHKRXQ9yoCho39sfxnSvw66xtsWHDzbPKAUTu146lT0GakgR+Q
Z6pM3e0ZeWju2X9+Xo4cDzfNfndiDRgYjLlb8rARiso3lLt4yg8ovXghnkiXQM25
57qunBabJO+ykojnLWAQLLdIHm/onIDrXK1oxTDDbv+oxKY+tXAktvZ8pssfwoLW
NcewrlPC7gfn9MAlMZyC8e1oAQhpwBbH1lyf9YtFBOB/Tk+iCkz660uyM4ADgMfq
Df5rB6iVYlw2nJ4atwtjk0zpstmhQ6UxTxNdSizd9I3d7yLfauarWYAH1IgO2Iiv
N79Fn6M529qIre8xNpAbFkc9UsPBDqRCCcjSGq/QXhtBKohDAWE96DVYtxRHi8c0
Eu7oHATHhP2y96kmdZ59eJ0T1diJEW0GtQT+Ew06A+979Y5q2a2hQS27kTUtrHgg
4LoA8AXsyl31ra2rFJzqeMc3vy+mIWP3yTy0z8ktITfKU1BhIGTjnFkI/kY55yMV
uQt2nbYkMuEEUk4hFyO/4cT/oyaljOe5mOHiGRtnF6Eyb5eb7NAkTEaM1UzrmUZ5
uI6gK7rluv8NzDppB5VloVMbtDv4e+YgY11Oq47Ua4/P5EM2d4kUDUt8UCBqWCzT
OB+0DGN6cuz2HoqnfixATLRm2wOxbM+5HOfVnUCSaldBFfnAfdLlvt5/MtJr/ecN
JsnagCzhyWpGfYt59012l3xFWiscp9l2TXfT8QwxnNyiWLc+5p1BTPQu4AEqd0VL
oF6wX3br17c4/R1IKpvEqINAEHP/V4BFOAgrcHjR0Od6KiDZBUgy69XjEYppgXVH
E0cvZjezN4Ky0FyiIek22OOy6fnA7Zs0RifTH/f1vCLIRsK7h4MoJGi2JzWV7raj
9lZepd2k0ADicv/oI1YQ4hUDw4FeNa4okWfm9gsycV0EERZ9YrK7wTZIn4Z/m7VZ
oRpkWOyYNYUaKR5+eoFgMoRdyyT2h+xrTqXiEtZ+FThV4mG0Gr0uhnAy3r4OxnC3
6m8uZBGHUTOcTvnKsh7pp1IycH1pUKv/WTb37s0Sm0wBCPAG1Wle9feOcUknTA8N
fM2thRM6iOuVIOiSCXPS7DUP8G9Vs2+b36rX3rjHTHyIccGpNJ/zwNQJzfiTBM/n
jxoSwhGSsc2+q52oITb6v4rfRhjoqMiGEb7NNLoWoV/TeYcyuQwvPle5KAO6iWr8
RPvZLCT4kSXty+UNI9KDFhzaJVSa9lBWxt0vwzW1KamtoapXUrSDAc8U3YmByCvu
fnDi/Xg9jOYsfgSgqNwVfoJ2FEyhbeBS5z4Rgd6s/LXJyRhJOLCfQM+FB8GZXtFZ
oyjF3Pb/xlwQp20I53Qiph7ZYyymFMtqLqSgoE9kNn04dip+II5BZZ7lB5PbKYJv
PH6c0p+aU3dptgtka2jlGAzsfYVLtJz2UOebch1/dV+lCVpMEzVIqSo+sKCXzWiS
Bt49IuGE19Ygo1lEvrEWmekvjYsXovKDrMkbpc4dk7yitrrGXZ5w1lUnxUsOnS7Y
IFPyFeFRPWGxIcy9STmNk+BYIdPeDKFAaBWzApAI4u+vhaL29/QNIrs3ptY2mYch
LwUnnGhXgvVeXN3hoLH851+ksmGpP4fNn/ppDLy8Y6g2QfsGdH1MrUZVz3otJDsJ
MEXDg2loi4XiVx06QbZSlhxrW85lVkTBhbIb4eP9AmTTJJ7RZAV62rw1vQ6lE79x
hkvsZ1EkmjD4AsAzRsJGQUtXEhjhuQsrXSOFBU6yV18wwhWVvGLP4LGl/sTeofWZ
eXtHTvsL0S87yN2wZtx8ph5/YxqGYpfZIn5eq0ThdrqVBfspzbVDZNOj0vj0AbsN
kw7sk/R9kmH4xjFp5JDkZT2e7QwnMthDJPbbuseE0ZCxIoTUiqFQkrPuth3kmfij
xbyRaH0IjiYQ7HXhYxEn3N2F8Qp1Q99Q2IfGjpyjweLZ9xFn4lojaiydybsaPKmI
kXI/8P0GMA4bajWIUqlcVkiqbIGrQ0FBmtZsyAisW7GDWMd1MctA7QmO0xYCL+LC
cbF/Dk6JdCPShGOfvyww2Ae3RbLQ9cCDIM0O+hubHiekwO6RSoC3+iVNnXDZMPV5
BaKkq2KOAvcxxHzVUA+9Sf5KPaS4ZSOl48XYdaYi4mOW6h4Leiq2TNH2OYUUAiE8
Mv01lx0Bor7QoBaXkE4LiTDwHYeHLF1SOLf1qXpUwrS6egX80nC+fb2DMNyjr6BK
oDbaSThxoMRqgipexkkbR/q/8i+LOfvqXcS1/CE5e6VeCynfO9fPBJuanhH5VM+J
v2KO/2dyKrEXuNZVew7Pq5+EILDtqJOukoSDI94262Bx1zCxqV5VO0S9zIholH9s
gUrZftoAb3VCg+uMBjrEumm19IM+AThoKor560ydGfYB9xxwzGxiColihZfqHz8m
0N5V2t1ihplwUHnPhGHImKssKToUrmkKvqeyFsMeesGhtpomrf2E0xjlT6zJtRvg
D8Tzrl79FEbh9mBxhIx3hufXVQgC6yEKW2DSd5RHbm5dKvEBTGpYTxYQJ3J90/xd
iKq2JVV//+vo09xQegIcEASl/xTinteS4c0a523IYXQvnVgKsdQ6b2vHZ8DLw4/V
luEs+xOAfF+Fs4BZ3LjraLP/f3miypWVeAIRW8uoV2nlozoe4qqUAKBG6XiWH8ra
x8KMN2btikcaR1p1Kr+gL/txq3t4QzmQI8sXq16fbliuE6A00qPv+tFXxNdzl/wi
lxi1al1VJkhgatHEG/p9q9hrUNpKVIIL4oyIz5qBIYjeRni+6B2sPS+gNccNH5E6
u7RWYZyZM7LOPMVEFJEdjf6LbLyMKRkrz3Ov9qNqs4b+aR+cfXt6rbQOy9WxetkW
DanjXy3SWjN40ti0KFYHX3mpwOSMccOkaCD8UwcAfqNim7pNoLm7GX2l67lFLJA7
BtCeP+6F1wVv1UCbGglKLmiuRtHWMZ5ZQvU3s0OjuUso640a6x/+l90K0ikF2kIc
txLrXHQpeDaruoUnNWyn8O5Jcclv6zw51oXw1CLXXhrwvrXswNIf8NrWHErM0D8b
fDP4rF698NxoWbv7Re+2J4ZuQKpGkobu1IQYQ37OF2AhkxPm1sJrh3MOV92TDDjm
tUuGx+Kmz5LGFqkY9jWr0Q5sWH4mjzNzpMN/vQLwjs3DHEixQg1pY/kio8L2Kvsg
XqqpAMph8lKHGUw1qf9ZI5tF8nmy0TKL6Q5YRTqEc+oD5dDktRFSMokxAUv/Tu9a
An8/WuVT20QlAqKRXngxuA921yU55aufhfSQAa2PQI2HoPxELJlXLhcakQD49v8Y
p3IqUjbL7ufoVYUT2DOJb5lZOrS1bgcpUXYUXUgXLjZt+uEfptPwmrpa1ztabPeS
JXDh4DsHAa/L47T9Zh0ECF/ggE4hXB6agyqxup2g0ppRfDzabn0wFRbYxUoAYDiL
FfDOkg+7/N/vHYxGokLiNZL3I7gS5ZdtyRb3sLWha+KBEuKh8qDW4/57hLHZq4OR
Zupq7h+nlM2/vveZ6bsowBLesHY4XCru8ItD/7XhjXtsYWjEWc1NGiI9+FsSk0hr
6MH/Wr+1HpHOStdAKFjMBqQ6qTxm6Y8c20lxH/OTMePvYiCbdEaXiHKRWQUx35Qe
SxREyI+v3CCZCZgwq5i1+DAqJYQ6QfmfwrXZVhw11Xnu5FWD8w85sIowwtx5DKc9
1lJQaPnFTWctDMstItLq6LFsTXsOw4GW5FGy1L6E8y3qT2uMAkL/vODrvchtJk2S
3VD72YgRX/GdH8l4evmDY+R1r47rA4v02Wdf34fkYeJnD1Maab+h+Gg86ZQAV9X7
vaYHBjGTsCLHuvimPpTYMmLYsyQ+1r/+9UF6hnOZA8eWlPGSKZSs2f9NYL2hIVVj
fYVqKUt2W1sgWo5VERtY4PCxg0Jp9YelH1m9rRurzbkbtcEqc9GPPyObokf/p12p
DdJFB2DzhLuUuzabTPPq/umNJ3EnCotDPIianPFOJgA9IteUKYbsJTc4WG76dacv
o7ti5iZv/FCDPr4RTSeqLsbu8KVip7BnGXvrkvzE/cTdAbZUTMo0k3DlPCe+mOyz
dZbu0mUbVuWl4HL2FGR2wJusRZP2A0h7zuF1VTC2kcEWHiHcK5sm4iG6Z58pqJMA
v3SXt9OGUK/UEV/Pdxk/wtoMO2ew2ef+GGtoKzFwIP+78sX3tEmjM2iqIF+QmVPV
gBnw9I2FcjBoQ9OFu5UDO/uIbYJkNezeJNQg40oZRyAC86jdsZn9jkRT2iHcAcKH
gvY89W60w3oW9UI4RMkEKnXI2qZf79Kz4Tz6T6upMqYllWZfVI4x3NPU89kPVbqg
7nzusK/7YFFsRGmmd0PI+zixh5R6SxfPL7EH43nYuvUg8SasmBuIb0Zso813iUwA
/Ek/pq4Sa9Be556/h5/4MAVGpvJg63kzI7hktONYjFInieEMPn7xC/nE9G/0jrmb
s8vDMQil1cuJlyF1qXelC3o92LfYMkB8hFwbTdzzNPH7/pEImm/PbIgjqCpz0fpp
ZAuB1hMqPjVoDUGWQ3CkztOoAOQ96AEhXa5PYiOIeqGoMafoVyt8x/r2GlQ5y/3S
2O575M7unHrzuDsYqS+pDIuenLlz1ioO4hfS9T4qpydoNLAdfKDDW2uTPwD16Wq5
67zhGIJ6hpyPWW9R9Ao046ov89m16EIlQ0DAYnRZMlUqdCMp7JJELDwW458lbbNx
rucgxaOXj6Y54ANowkzGwnamp98DGwqNPSavCGah1Duxb9tKZW4o6sS4U2xfP7kp
784I9E+FekV/lrFG4EGObNtaLeF2gMMZyliUS9m2Nhvchuwxl21rLXOP4fG72r7F
JGI1WVAySV6ZzkECzu8Qxpq7wQ4xN2ljwUK7owRH5ac7PELkk+vxNU/dj8YAeWPT
zt6s6ZFK6nbSOws+0Sy2i/S/qAAPJqaOv/KEp39pKKSbdgOzFFEyEHaojvt3wVFi
CmFZhw6IcR9UJnnKZJtwki5+PGJWkkWQrhjVGxbZcV9i2eLBLqSGmd6GEJBEc1np
Ec+6JPC9ltwIPnLvKHpuUsy6H+7uKzsD/BqvO9shkvKTS3RSW3Y0bptJnIojnSub
q4Dxc/tr2grOkoMwALsQN2ZAjXlNMesUAah4OVm2gd6rpFuBPw4E8i0domiqc14h
NH4CUxP5LoKrnpm5HpYTry3hW5E+odijlyqzF+MIX6rHqE2RHBLTj+YsCvbtgkpm
X6fFy4huehDuTPhbXnecTdcrGqfCRgZRxYTJ304Kwg4KmR8Srec5E78t8f+wAzw/
yPJ7QvQO4g+G8F2jeLKqthiKWxpm63sIGr2239JrYfveiQE2nxipnsczHHmL2dsM
vrcoj6VahxCiqQfed81sibFSAiSAXjnIN7fT14hSGqJEFv/hquzEMJQY2ULV0PN9
7GiMzjHUUsge8W5b9FOckID0FL42UoMTwfwifVEZuAKQOm37hR1Viik6gxO1SqPV
mvooTPEBDhprerMdiThOWAxKOs9KZ9iWaJyhfqYXOB70LqFSQI3Kt+rKn4pJZMWN
lIHZ0k8UP4+5ulAET9Nhsg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
m9tRUpdj6YQ4tVP2+1dyJpUd251cgLZakqYERgmso1GWKBBo8AO1hJtVi0uU84oo
wj2hvB1z6wMiC7pDSCmN2X/fkPq/yab2kwBz/TUl2ZVgulHqvs6Q4tEeddMsPWbU
4oyhjFJYl+j+Qfnt5mo+Gqrz1hrTXWBpV8u1Nz5uBP0JzIirebhyzxawC172/rd2
fEyaIry+qZYYNEZbV/6bHDATaJi9Nl7/ZkLltI5IB0Tmap/rTu3deG2Bwycl/bDj
xVPcdZ39Pa6y6pDlEvXC/2uP3OEv16V/2tTjr8F+9sazx4aQ0KzSt7oR/yI3HreE
a7aPCobSJd922Sjq6b70vQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 27200 )
`pragma protect data_block
pq+T4ju6vwavEJ1Yw2aNknUgDXch6nB4P6cI5wBYOXRufvHHP3LCPKcsmadJ/aOM
apFksZpBKyZs7TFXGV+tQMbUyJqETZPy+R599HFoFsPG+UsrFaK+sdQoxO2/+7cr
kL5ydTvzE6Y/2iDFUvhIffIDbIfM0mXA5gzISvfcH77ZAOzCPRZk6GCjsTE/onOH
d3DnwRGa6iBvxu1ZnAjTjsREy5CLquli5UEjPWCGO5Ea0jOCHQG09wblxyirJxtF
W6SPM1YLUHV5sjYL5YibF/oaCMjdRIkutHF1g7UDl3RCrbAQRHxzPlwwbbSpKLZ0
PWH2I3b5Gu7/F6Gv5pMn+Y9seJY7j74AdCmu190B6q+IFW8X2/vBK4MDGU8Cwcc7
qeprmF3EcMkYxM+KiI7ZURshKN3H90QtdwbcPYQ8ajnG9VDP6nrtXoyADakKBuMM
3dQiPHqUXhu5XBkDT9T7KKVTNXdXKeaP5j+1mqCOYe3pIgkUmiYNFAqJSl91pGda
lBWKBUDLg1Q/zT9iUq4oqm6QoG6/C9mtYl7Pz6zR4NX2m/STgoQ0pxnFbjWhT3Ps
xO0Y0JvdrGRKyE/zP0p3EgsVotu/92/aStyLGb8REkIesxRXy+z/+tpt38qru/Ah
24Ucvms1W1QX6RZm2YSAGIjzKN6ICveoDdA+mrRY5QMTY6yycDoRwCGhHBVxzpLp
6NgpmMJK7Jz+cIIMgZ9gA1k9rprg2uXxZbOzKQ92+obndBu9Z0Wio1Wjyy9VtlNo
Z5xIySn/NCjQnOopufyULQJVvhw6jj++M09ez5Rm7AzWjXUhcQxzBKtZWhZ9a31K
s67Znt1VyfDF68gZn6h0Oy8OWAW+4Vm2gN12ozEZ1UaWBCqv7I55lsMeFEzhqUHm
wuTR+PfjgFMdzZEhxCVg1N74h2fVbl5yRS3WkO3St5H+aEeONaLLE3qd8DOVFuJ3
4QKkJEqlpjT58MmAPxidanjMuKFZWm7Rwa7EmemWGPvd38lqvRIptnQDl3/wQg9w
A7q2D1M6svzBfR0R9tq88IWpIeEBtShFBMKtZZ+tzvlHPQsiafkSlEVbB4J02Fb3
r7boNwW/TE2K9NoJ9ML3+Bnl88XrA1nfj+hLUiKvOtclFWs31zPVLXmEy+AN7xHo
qsuBw688xxa6/MC6vICv9+yw3zUXL8wZrTqdIvvfZlPSCooFvD0ZgOW7qlOK/UJj
okg8XoxqIqLQ0kr+F0Ea4vY1NvEBDP7LxI1XG/ZrJ5pa6WyrTrqXmrvo5arlsZ9n
/JgvP949GIL6dcGZBNQR2WuAeQIwwu4tlbbmc4OYFLvVhKSazEQ+3q7/VaW1cEX8
VrH1UU5b5KGQr9GAIRAt2lJ5kPbcs44fUjwQLGqwDpn8CszRnK43mMgmLhZ/oWN0
nt8XC7lkiH+JAPOuqViJQeLSgMVvjEPVaD7v0y352WY83BMBCzYn3CQOvkNzDjHn
dG2CEbY5tvzpX1ZX9adOo4uc1CSmpaXr5fy3zOSVFGt5hmlc+g8Ytp6Cpu8aJ34G
dtgqwpWCg4MORSxWXBeRmwqJdFDci+mo85Cajc9HT7gJuO0RVQH9X3LMQS90W9h2
fVKvGfuuAARfLkS0DV7Leobtj3H/4SQ8a6BQs4LaYC19RTkv1xxUQm2RyQC/T445
l3nUmuetlaZt3nt2tZPu1NzkwCFjTssYauGVFK6X4xZPSutcXd6y1CzjVIDL36k/
mnHRWla2ZsKUc13Mw4u9Bp8MY9qLi+SyK4r3eG6RI7PcCFebFiOPm7SI8HHkxMIk
tmTOzOGQ6k+7WRMkR8iVl5BrC1Rn8AH2DaG13mExattOPR2Z52C1ojOpK1TK/Z+T
ECEZjd8/PodZ/fbrRLxnLhDdf/Dz0rgtXxWR81v61X2z066iRe93DalYR6vtEhkZ
8hHw76X8vAmwOWmLTyZSMpUWFryFkCsnYJbNhb6YiTav3W+uWkMwe0p09VnyP5K6
WnJepSpvBL/Qh+UEr4+7GEkDolG3dxGUTAKBLyR+pL5uiQZ/zfJESnFZGsGD5S+l
RjEVMUm+DzFUJ+2dIahAVUd7ToUqlsqyfmETnhZs9FsTusqDeJfDcpQ4XBCEUXR4
JoBXsdNgoUI0vyJC+8+AbidHwS6Vu9WWXwQzWbe9Ly+Ww2t/yG82XHxubSUKFrqw
HTwV65m1vr8hwEjntF//Lf+lDZtFk55IJkcWYC+WuCWGHTV347cEUfDvK+SDIxXR
SLd0OT8FSfT3BWk0+yzh8LKmg6WuW0ni8dqwj2bN49w8KAHpPxdx93maTnlSVbH8
W/OT22+eWeb4n12UZ3BJvsy+mzqo98MsFsZwIilQDr9B9labCcgOG8SQgCFooATy
ZBR17xJiCjFp6tsJCpNs52jptPGSqV93EBBbmsp+89F8lJdlSuT3RhVUbGZchpRG
MR8DL6icJsdcZWdDb6jlfKtIRL/l1os8YKqi3u/1qeqUd0XJGBVXkaDLdccaE+U6
TKmU7Qb2DhhBNRfZ/N52OnZoQnGTux8Nlw+AqtmBqGs7c8TJ5cqZWf6lDjxqhs6v
jfUtBJyPgrNRlQcAO0V3W8ZAzDOHe0F9YmaNVrKhAh205W17lHoDWAdB2hpvatqJ
Zfpv30ePKz4DczDh2zM4mYv5mFDC4GJ3aYTOLpSPZvaXh2g6cf2KgMC6ZZIdBW6u
9W9MdtA+2cPa1s+1Hid7YGDhnYImAEqLj8yyIgq3cJzgxGIz7+Snpqv+81SeDXsM
6Al5PEB3TULuZFTUDlewiATiMarG4ttLYVOUWSRV/3bnmYpV2W0b81CSTFP6pe7p
tpWIOJfmmgoQKfjJjdpqeIADG1heGkAbwf3+HDWl4piNXA0k5g5PDDWQd4HIxAfW
dRV0pYHpEyhxiCzBXJjGnJFmcaFN1SPdW9tUQT6s42mpsnd2v3EL4mua23JTGDKs
fB8+IAKqSgf+XSmrdbv2FXKiq/9Log94H0nETWVWUEgnvuXcoVizrnMoq26/LC5g
svpq4omxf3Fl77MLddqGBv4Isw5q23aaZmjk4I7vfoUx/jV+eEBgcsGLIQ/4X51j
Klyfqll8Low9RXYPwFYSlUcpYwE4smPDnP1Pnhe0MfW83LKBX5Lpt/9yMvtuSi+A
vL9wEUqwLcCvwU1nK0zNQmY7R5UdBvZW4MWgBZucZ+6HClu91EaCkwJYxzi2xLu4
8nrxr7vuP5vBOG5BSV1op04WPYzUol1AuziPHIhwbMKOLK/Sxzn1nkuYLs7+Ke3S
NH2XkrbYSxREqaT+uFH0oqkpfr5ijM1SxVDP62e7G+HW3c/mwTeu912Aw4wQL5nu
ROWun9j4woM5cCoTTYv7R66CjOUPg//26Vf785NyMQLrFwK7AN4sGphxveE5IIWE
DZ+b73EbdtqjmEgF1B5JJS/BAL2+LEV9SDgV9FfW5BXNCC7i/NDN3ITJaJg/dubr
mUcLP6tALfGZ8CCvEExX04FkahzpZj4CihYi3qmaM5bGMMbD393ATXjGBapbOHZn
8ux1g1pw7o9PLEpypU9EcALl0ja/+qK0kaf/t0oo98sKWwdMPrt+2g97XO6m41t1
8aBHRUBMOgleEvbGENyfXXsb1yLpP0lAK9YJ2/dJFzn7UvjSGi4G7NNAScV2JH+v
Gsq8y5skkjxVLqeq3M6s/M0EI24brHRnxVcGC02dRQ3SJ0vsjomvEzB5V0uezyiQ
DtIIqaapx9sYBUJKhZn020VpvL/wF75BtKP1tGs/rtqcjft4K98hGEjlaZiOdCmd
Y+aOLna4TUsuWOGHw8y04TtFI0iA1l7zJfQi2fNoKCjawLP7/zjzqK8DAQB2Hqyy
EcBgGCSBgxbnvWLV6/X2CdIbjZE7aW5MkBtMoV6NfhngtXKJUHoQyMV71pp/9f/h
NW91+NNQUpCDZyybux0CxsC323hM+6laf4efWiThi5mcnHDaN7PvpRPARbwU4JW7
LLCqjEHU5tvTqLlP4LQAXsklPorgPjfz8NmVBc9qtnvw6eM1B5uLpz/rhuXJq1iK
59JywUivodks2OARYme7rjPWgh8Vczx3/E2JJJXdZqUBzjwP8E2fDiO7J4NyCP7y
6V07837ur24t/PAqWOkU5K3yUiJi/WRUwVADtzPKOI2YmfQEwduLK/hSq/ix1Kln
Vg/WzvjRNvm/W1yzxvgfbYVrF7qIwWdbIgUvM8tR2BuvllCXi0HInGws8i+48qxg
VvYUReWWjAScdEISExKiXhhVbk6q+yVrKigC4/YD+oLENEFZQJ/oahMs4gLD4Fil
0kwR6iR7ORTugyrGhjOG+pIta/BA+nQMB0z7KqJ2IEA64txik/lA94GlFsXVa+US
tiX7G446UPD00SNdh30cGalfnxc+qQ2D5yp17tjMRHfNwT7Dnpme+0tBDotTyiOl
g0Nfq1/gp74y/3iTVNfzMs0chWG9f2NP+182FtX5hO+qxWSygD9pSLcrCeRqzoCR
B9M5o/vtLUyxDtv2wSLRydZfmTSPKHcBo5dwvQ6JNBUeexItDTQK68DplZD7yaKR
Bdx2TVzVYn8rKSxoT0sQ8zQpwIKr7YJZk0KaKfuwO81Ye8Kpwy/JGrSmjSpyhhgL
v8CgZYIrB9NvA6zGsIFl/WE5M/f0meEdbFuiUj0FgrgcLcLGw0NoGqNXdwkIPJOE
G4vUjoERT2wqnIeAf0uNWYyMvXTWyIno6JLtHJ9vm2IoVta+JFohPibVDB/h64/m
zSpCTyPH2jc8ExvMp0mqOJ+ROYvqEaciaK6sLSePowz8U1KuDKX2LhBZATUM0GEg
Aud8xPYA72vedWrgRRO0pEIBDe5lmfCvo2iPE8kb9np6+1Y47mTSD1+5HAmVY3Jx
iCWXIVkKS31dQ+Cq9NUqMTf2WkJAgMzJYrQ//pSvMTLd0+/ZiXUlPCePgKjQhV9S
/pY1fdmWhXDceQEN/zCn7gZMmMtgmE8oVLJQJjiaM0qcQXRGF6vU+49FjdIM6Ovp
7Bv8RkNF8uIFPIhG/q5Smu8jvjm6HwkeYVH4XmjZB9HxPq634Da63KkUYTwcL3dg
keWpUKgrLBwGfBlCF+Tf5FuxkWQFrEmGZij+YLIfmJVBH3/GJ/XEx4/w2eTMA7IJ
UhL6er3r3GTsmS9PB+B/8PXvsuxiqM6j6kF3rjLMtBXhRViEq3b4fRydxhnNT6Tp
S6jRB80LQEw8mMkkn7X919PhRiqaCt/IwuB/rTaRa21dQDFpHkaBKG/fKPbIOkSA
LQ5+iXnl7yohXRIHByhno5krXiV2Un6w1qKcvTl3BD5Kz3CJhLiyjiTeexb8s3EZ
aczdax8P7WsZ09ClGrFkDgocK0uE2OdcCYVc6CWJ7AYowoskGqbWYaILWjWQgqVP
pzQREalIkah9geSITcT9V5vQHlvt3wGJy4z5moyoQpAvPVVievTP7b/2W8jhmz+c
HsVJGXbXqhmJh2JRRocqsOAOnTdd11z3WJZDItpAbQeIt+ITqjXR9ccxVPsQcxrt
CjqfSH3FbSxYbuXc2EbEpQkRygZiBji5DCSaV7elp03eX8E6B+YbfzqKyjnGf4Ua
DOOnxw0YRqvfCtSHalvYMiAt7DMSBnJsELyFVrnu7BsXDKkLr7h3hn4jPTzjJJr6
2NAkeUYmmnr1S64dPYjLP5nAg1lLBnBR0Cnl+rVXLZ6RiETm9PNh8BhLypv5Mn9s
2gmVOphmsbJrX/e+kGD9yaKKefSfAC6AEtRbAhSvZcJeypFhQTzsb/jEPyrWktXz
mHqJjSd+1q9E457gR7DSrKzD/D9CS/vBVJ/dKyaaLeTgYk2dHjuYT4JWmRTxfQ9N
IEORvTvVmeYdIilVZiiEJcCWxTCruozGPgr2uymic6f8tr60Q6dBEOrR26itJzXs
rgnilc0zhGTpJ+cFwcl2sBfrgdv48zrbT7B7s3jm6yCxJAlHhEwx76OHzdprvh8b
Oo8U5m4c2f2KLOWVOaiQXyynZkaG2hLE3HZHmMe+gNzrfqigjqautnguhImY713z
2CfJ/EqVXP/ZSeEHX3wtfVwLCzXM4htOC45SRXrP0oGlKcpoF8WnTVdLUAdLjKxh
W7FQcUFDoUz7mKcXMPX6vR+oEJiyvglTukBzulwTXQaLCO3J/6Y4K9U9JPEEyhXb
hTXPW00837knaSx/DZu5A9DWPLeWlWOxVUojQJ+hS2ZU6KFy3GXMk8Ekqfht7Xz9
EohXFvr6KAH6qTHk+4PTZNx/hCsjcvg3jANgRQvXpmTdV7p68AhGhm+WHaizJk/7
XVgoHLdsY7pC1mZINOdYbFkGgLh95ZeaUbgO6Tv+7CWD0BxkUm6LL07BrbVxYOrG
r9RZIsP+6yuatD2WDPObFoNbLmiQsqKdXAW1Ks5AkQRL5U7miAwGjQJc1YwGuJX/
1D01oMORmhVGFp6Zi7b/D/SKVmgLH1MdASAqaHxpZ3x34ePqCeRCwvLvjlczca7W
/KpafTtZ0vFMjoJVFXfeyVIUhRNYZojfiWxV6wJ924NkUt+R47DtsSmYWXcITNCV
jHTsu7VTm+i4KWMG///kt0dsqCkXG8P9KODVEjNmpbpUw6H1hnnJaJoKrUR1fET6
9G7zj54kHdw8twr/m+1NWN6/jRaV/vt6pn101pCG5kmE3rYc41wVfEOmA8DZYraE
pcZZDhNNQMzlBBDq6HG3cdPocBomU+9sU28lU59OJBcHFFC4jP11Uuc74Iwi2HkP
/iYiK8anqow03OfW4n91nAeECnnTwBJXlf8Vi0QRE1wS7RdoXqiLybcxzDVOmnY4
qPi9jGdBtQAJf841np6Btj2s5KOzBl6XaWz554F2dNwNzFhUUdnubGxCrwO8+ou0
xw99XXEutlIaE4sulunJsc7vQ903PuO12PEy+80gzW99vy00qrk+bijxbAgNtizU
NyGZ5aZnOvUlx49m7QGSi9BlcwaYm5FHqvr9munX+nr9evi8g+Q1kJ5fjUNv7iIy
VEQxr3Gn5sLX65NrxIc1oZIlikVYv/jNaMTGj3XK1x7qkEHMnpndyQupNo1S93Sa
V6uSjILni33Cwx3H+wXp7QEvMS8XWxv0OKscQDkNkKTgeiULbsajcSjhQwm84xLz
JtZANd/GF59vNquM7gWsIG46pfoVmlj/4c5TAi9YpdfS5it5lD5Ya1uZi6ifabk1
kaY0aNuNw2jvFMJvW02Q2gdnEPGn1YuLybGiSkxH9bqEThtYE2HXU3mjMQECrBe2
RMUVnJ6mqmbokpca5tBBgw6WqdGB2NMbBejkRERQ6caKoBDNh60sjlzTNS9YZABd
wrxIlSFTHE0iT6KGiPH2nIQDMiVAOVPiiXDFnGyTnwaXR63j+vOZlKlrNf4NldkB
3pF5HLbC/OGVC8qAjW44N/X27tuCpIlTj7iDsUZG8MF0L5XcfApL8Q6skqemSUDo
jKwNuMsIu1B2afO/GpNYrNDZV8uRgKSRbDJ38PfMrJHoV7OL2Vrp+FkdXkvlO2sn
ajPQ736cgA8lVTzIbY5r414BcOXxBTQrr2a/6FY25tUhzhEAidvJv44Jtl15SIyn
/KcMNYBXyKs+7D4LPtwAHCsHeFAIvl60YkjPkbu/k19DfbDom+0uojbZnVLhpms/
HlbGTiTxHT4rKdzMdeWhsXCRbs9Or289Lae4fyCOQsLRZh/rUWcG+B8taKq3Sw0a
bv5VNoLzV1aht+Rs76MBEK4jROpJLtbrx+ZMX3xZ/8ZhRiLPi1Vu6ksl5B8mqd/B
ARJj2mIFc6SBqHJCyJVMKOHHfPJZHtSOR+H/k9EVmFZGU/0ooj9Zbg9M0Cosn03G
PGhiUbWuPJd8etvMbD1/9P1jfRLgimT7wn18HpyOGSUfAb0K1tEQEASnAdfn81q1
xO74nN+GemHHI28h4pBhZdV8QGCsYDggHctEJRkB9NK85/tYwivWOnrEAAYjfFzp
3e/fV2EccmnAtajoThALOyRvRVOAgUSFZfrau4aAp670+kDLdIdiKFTNntiENDyL
2S0mTyYcdd8yy/nPgwHcY9zAz3K2qPy0dKdVb+hddFV6c9wBcz7ymcqQJIRru/ya
4T7tLaACmpX/IFbckC7XtmYmG4JfhwZEWDU3rQoz6hqmDoq+k28zfKD8/LUHPbVl
r0G8YdRh+rzbegV4G6gtI8wQNLv6ON0hlcjb6ZWF73aIXywrxn0C1AUNwQI8jIL5
b6gRDUknNxDVc2IYFqNzz0d+rWsTwJdsxTDizOiLbb24ayMr57VXGt+yDJwaD/SM
omOjwzmZs73co7RLhOexqaihKJQccAo1sHYFzpJ2Bnx1NzDw4KwOAVRIhMxAElNy
qTro2ZLKbzHOOGHxYUYxQS31aowHhySK2iHqa7wsK2Za9Clk7MUCl9GkN7QgMzrz
jFKY6AN/u9/FwKFXzzG4M1ol6N/Cz8indXwPsKV4TcLQxzn6Spd+rZO2V2xxrZCv
/0N2ZJSnKttat8eY042SIn+g47u19LpVOD9gfswuyV6KQYphlagLv4z03g3aSrne
P3evz/YwJM+4r117LpHgyp1l9D1kAGljuRlSN1Ty18qhSALIHAC9DDFoDslZ6HYz
EfQGWQoACSq/01kU0VsxWdRhJVd/Im1iSBD7Ax2ppYEnN6ODlPWTdzkVhqXs1sHU
v2wI11ffbpMlhRSNq61Luu4B+CHxVZwgFz3hlgSCzFoxjPRXouhjUjsWzgWuKy5n
eNR/QP+uKI5ie9ASDI4IB8Ss8bOaZL60/7oSXOM//q0IZC/XK1RRxoN59DaKbWMJ
PDbstyglwvuCNDmgsOB4BlyugRX3tD2fzCEfLbTPf4RTfehe+2QWgXW8Rp8gquiv
+Lderch9XXGWFt7j6MhASkHCTnt0WIU5GY48Iq6mKERIAJZEaRdm4byENpXi8SXP
6QT3BHoq9m94P7TRdzc+w4SD421Sspg1A8MThXshon2Z92lqeHmiYCu6do5JR7e4
HUADjD/syiYVC05H45/RRrdVzAKPGk30Qy9/QIGSSACMfXk5lygqnantFi/5reVW
Lr8tAidVw+Lj/eauUbsKPSU1GfjHrXK0GeBalSFPcLCQNxl+SWw6Lgu4aXfN+moi
v4QdlD3UcEFbJu7UyCd//0AfiSVe5n2DQLRgGwAL0dDscRxGM6IMLfbLG4E3sK9+
m5OrYue1OigBWd+QN2m1FnkkDf3sA9XulNC1OA880N9XzWR9PdpZtWby4SiR0TUE
H9P4x/dnwdiPwK7hy1hxZ9K/XuptQlNBWsDeCbdX3B5cekOcdoGNTHconEFEcEu/
UQBklv5hIaEKkFhhaVjBoZopiBpJgea7IT1F97UBUkVXy9rSUS8UOzQ2xKjUI/yT
OcA7PzR8Zdg2OUajNhMFSICcwIvLfqY1SOSME81QjxynmPilkBiP73on0MEo3tdX
pFfXRTo82fYVmxu2cBZFC84qNiwUc+zYkYPzbGc+74vsHaE9/HANzneIK8Bk8y1+
aWppkrjEqrLojgu60duNyRYPrD5cHiiWhchg2+bAwRF9pBSMofIAXHTB3stx2/zV
cPtE5zHFOhvInMc0kSZLgZxKwCYge7v/JlOBC4b/v9hht0JRUCtq5fVrmZLRavP5
8ooPTjSBvnHOnqkYacODNVWyLPCqtvZjKAZxI57diBVb58BeKn5+ozX/UukroHTj
G9uAKyqAyGxbElzuiCftoTcf0SeVjZ7DsfFhRMnMl5VT4G0DgUM7dlJtNZf8KUAd
wsExH5oWL6xPo01p29ca9X4WB9TU936lJDwWZR2//ZDDwM+6DerzlrQoS4In07oQ
GH9NFdgpncSKXfpnLPsexW5kJZBoL4KZs9aGOOpEG7bSyDvPFSLsYjrLFosdaOJL
kgSREiXfHRUhLsx/wzVU2Yq/Gp0nSRbfH4s48tvK0mpfF9LR1sbyJ309DocW6xgy
MHE8rHmPAX8iYEQ5i6YP41GX1x43aoywYmZBL3d6gm+c6M3bv+Ii4KwUWDwwSHp0
oovzhf5wqAGRQAatBea1RW8W3Kz8tKOULDRiUxh8IQ0sQXnYvSrYLU08XD7eWR8s
93iITZjRefaxzB9sdVFqg85FWlVnwifHBo22A0JPu5gPdOk8Zv/zPloaaq1rp5st
vQmTXH1v1V8uYuEVV4HpxFSF9t57/CHe1xJaxkwQ3TC//a3VIwG0Bx8tTzQKy42J
YD7P0B+pSL4vFII8fCQ3cNx9Hex830KYr+wp5obL+wOTrvdsAziZq/xWhumCtzBC
d91BsQr3ftlIFPvThkNJn0OcG3CZyLSwB7FvdIIaFHhn/7EdA++TIpik7V/MvkVD
py4TaX+pItd1vWC53nOgKP9O0B5IVQYQyQvTIv7qXerOAnhiheTN/G5uoom2FECk
df99tzpFh/5oi+2uNKpVpfC7DmBbnwuz0FTh6EviFk6sW0KHb1FPCfkAH1ZTpRYj
P0FhoawMZeL2Rf5njA/LGKsrKuu1svBitBa+ml///BSSOj1UbZpUONXTRUijmgCY
7k8YUQrmdJBxRKI6iFBfL/TvrvqedJvhSYh/BmJobUe5qRlFW/R4GMZMHmrD6xJB
qR3ijukUxxm88EcsC/ziQ23ChhfFnleBfkt136GYZr5zi6pCmL9UB9KJmzuPYYl4
0kjD7fob4yJHnsOkvVThxQKH6im0uV9bCjmB++xyLAm6Hc0gp63CL1A/M0QOCvup
3jbDYIwThcWZ7Dsm0V4vVgnlh6jdbJF4p/ZmaGtxvW+dUt9TDsoXHF9s4pG74p/s
ItdeP/U86p++y86Oj72zOpELSQt8CRLlbhvL+wNuZfnhnKrgCRxlpFqbjuVtDaS4
y+o6/6InV2jWHLknhgyZY4fewnoWpFFn/DilltGz2gSJ0UN9RXWbP1HY11pybqtm
RFG9NIyXbTYkcMMow34L20cvgfo3lQXocaOa7Ob8L52y39mNSYiemihzSzXAoOCZ
VuUtXmNNIiCYsUKh45Oi8mtDliQH2Qs/1unZ0FBCZmYuNY+s6TyXoiyXWXO+8nFb
GE47it7f++66zZ+M8E6kjNE2sULbhqMntIl05yOArOUQ4FZb5m/l5qvZhovfhSOu
jrwLPkronLruWY0AYK6m/T97Vm/2IagfIOQsJ8Fpjb3683Q7rU4Zq0OK/117rLUT
t8KF7VoZkqHJzfE3bIk6q2qWoLIc9VN1EABTOX36b9mVgAcQsu1aHeQusvz6VYAB
WrvISFG4GU4x8QtS+ZBFoDo/xOniGEF8Lp0LQ3gZoYoSly7hKb09Spq+Xgtlz8iZ
KZHRWv3vyF3vZl7ke4/a4SZmrDkaI41na6szVl8ePsE7NSQ0au5nbLtg4BE4GIyO
Nqs4W8Q8dOwj0Z0SxucFPGrEi7u1asUfETX4FLCtYEvkM2hTeJdzvQm8A4sAVP/6
MH8tlH2tFqX9MFfcoQ3RWaAF/IdR697UWZoF3dz/OImXYRxELTMtTYeOoeNno9XZ
1FkNgWLGbuHG6vI75B0WsEyAmhwAJ+aivrTrD5uort7XhqUo1gwU3f5R58iNv/3q
qfAzYWimnzKj2VY3UaM/dzJF9AK/72Bxl0fw/tpVmr9e/qLns1C2FpAJVnP5pHIG
hGf3p/baqJ9DlTI5aaRbQwxX70fQkpYZqkDHNrD8tnuk/oXcHth/B7N2EhQGEQ4B
Ub7PhTRJKSYYEyy1de9rP0YaCQ1q9l4+5g7v402VD6rsYcmlxS2cizYfHUy0dksD
Z2VUUXGT9X4590ROCYioCw2t8ILu0cRs2FUcxZ7sPHph3L437poVYY1yoCY/FWB4
MRw/edXdf8Ickqk18pMZBS2zHps3hOjjGx6CcO53KgnO/RCdCHMPbwC2A2g+xsZH
ne6gOpBlmtHSg4WXvk4LbAjQGeMkO05IDqpNvMKvdIRnV5z7oPabE30SfM/i91p1
hfiTVisbbirosEVTTNaUJRWbJkF3GLH8rh5O0QACy6E4aFMcuMKi1QiABWUvHpLr
0yn+m7Uu6i1Wx++t0S5cKhHTFM48TFljQ6HxscqWiyVvzQ43TwOK9RNtwDYBjlD2
IwHKeDKqZpW+T8QNa6g+Jh2KxasB/ntkOWJFgwh7jw1Ez1+yGZt6ez7J1DSSaBy8
GERzggsYUugy513EgHP4S2Wxz5ozWyH5MrI4TFUN+/XPKOdcqyz/XsuAFfK0ib9b
Vfea9xb4Ct7W6oxjGt+MF1Bac+ayl3m7ip49Jykjx8ubfEoqsw7IdVE0KBjwd237
TXH8/I2aqZ9nYFO2OeQ4OYFEVGoqZ2TiWdXn0mfKmdIXNUVRyWmvm4XBIzVZLyMs
ych+FrWKdsWFPCYS2I42J/HGyaJlr/oRCFfL7icdm22iw4k+k1b0Tlrcmi8oJf6U
R8J6ES0l/q3Ro2Wa76EJGDl69moh69iOV6LMpcqJyGM/p9v8PhqcnUgkO8K5YlTR
Ekp683jQ1b4Woqm1AaTvTjNZbQXcGm2ywBX6BA5ySJUPeCE3LwuDfRvk/ZYkMU90
wr/N6J+dt3qz1ACifrPkxPVNspvgAW/Kb+Dp5KTuH853G0Jy5l0NqUPa4tpBN14M
S9NWyvhXXQ9V3xSSC+7zXeie8r/sm7tzE78DqsmLeMUi8i1RWj9154gamoP5+kac
1KyIETsNvv/ku1UFm1n91hdynseO3qmuI8SCKz3WVukfjDP7nebUvUBiC4RSrLUN
O6SaBe0CytG708CsvF9MN+tKHGDKFquTjsRil0T/unmrKcm8sprPa8QRc+RvbDPz
opAvIpD/Rh3/FJu0A0vGlwe+kqG88RjEf9kDB7vlE4B6MXS0HgfEm/EACdK00dkw
C2ZdvVCw64TbVwxcPzSBZnoQhsELk5ZF72ZDx+/i6FS76/JRY9xWnKHNTOjqIpRf
JK0hRNdOIAL92qBVlqe54/k/0dnh+S5vcnGy1oClNPNw2f3f06cj8GzciioAJQbL
rMBicDMn9BMu28FrDuT+fAsKeT/CUJK0VSB5WDiBfZOwz6axLojgD0MjJJSaM1Wa
FvaKYDXJ6qrIwbb91VKBDVC6NHzNL9FXcmQp3BdelFz4VFsVqtu90iIp/E3xvpcQ
Hy4xgiY4OZa6S6hPz615y62Y40UvOWuKSKLH0SfIn1ZRyP9LVwi4J7kEDEuPK8dJ
eJL5RaxzOqPrCxg/XuXvJ4AxMp7IxgEMy0JKHHYHfDIrUTVw09/noitFkQj6zaMl
XwkCNk7emG9bf8C7vjy9a1Y0VvyYsToeIPHJgIyYOO4OrL7qXRDzI3IBtIKdAYj1
tvAftDgNddrSo75eea9zXfsgK3Qf7+0pMUTpk8ZDcu3zIz1cEFIpfP+Q7/fdAgSc
HRjD9KsIgTC/B43m9VjWbicvEyUQ11Za6Wokrr0kz7yUhxmaXWmPIav2jaL4w8iA
mli/YYps8TtXOHtWCMrDqpcBCD8PxYU3DQjUhPn6CJsCRfsKzF7jdEZkMNQN5qB9
XInvildJ2r3a9/kQhLJGiOSa76xVWbIbyd/YsjQJxTeDLZ3xOYbS3Bkf0/iDR+5k
miOISiifa8861GHGznMKgo28BfkWYtMX/YCbc4SwNESbGWS/XODbIOQJmV9V7s50
LqzoSf9qVrZYCDz3neb8jqdB+O/o7L66uSp/eqcolz4VsuAn56npP6cjEaqi5Tar
RHsci8SZ9quoPToc9ZFEde1U5GpyvnkEmab8NwM9OoZkWquV7jIEdKlWAhqUewkk
ALL2oHQeXpYQRZlb6TBEB8uWe4vpzjP5L6oRabWSkFsFPG7tYCWo8SiqCi/aQHlC
4inO4beMuUMpNqQQoEYAJBHhoU9xfIG6oS3KeFm2mhD6GFsTOwmsW/b1uFAfWje4
bnqUWGaJ/7dWJSYlp1F98/a9Cr/6vDMemCBh+MuW5b3ul6pZsFrQDbo4rdexUQzQ
beJi+f3l6DD6LvE22S4iGE7voocqnlciYtfVYCcwpBag2hyxZdciffAc8PzRHDUb
mVzFg0tHVhuBG2EC6VlGu6aYse+xP8Sc09i2A0Yac6UF+yoOnfshs5YnceFxP4HX
kFSJBpFRKEOXoXRg8o6/66RSumAKq8goMQNiAAGGtgpoloJ08pVEyYOrV/gVh5j7
5fdE4lmMsRz/IG6rJ0stsEjT2dG6OKuKuvlkEMKgMvuYq2xmF7sjW11SEABO5ey/
xo3iKrBYEs8TyHsWwlADidK6y+g7vHgTExJzQtkfwG5tFjX3UMKyJqNP8lgQlixh
ilAd/7fEP5HWMigaM9rC2/rgv6yMB8h9Zoq7wWJ/QqIAZCxZNZpMq8pLkr96QbdQ
Al+evJyvy8aHXUe84JpaQeyNKG5PKSDzgsYTL3TwKBFQXZrrY6edWu9JaDWJxnSJ
9hQOR3pmCO8iGNDwnR3PcQc5bhk1PK+cyQujjk8NTBUWoPCF5YKGauSXohWIlncO
IigfvA8amYRR7Zh8JvGhJQOirktOmtqQxDuy9V8FKywkHxTvKaXtrepsUmiVFNMz
HnSu+2eghFEprL6YhMQZnHagvtBnd0fKsegvmLj0MqZg4/PWX268SsNB0HfA0jgf
M2uax+JR5s9Fh3Kr+eYBdbHP/yKSicKMHxT9ALF439MluNeOUyytdqNejH4FPRyl
EykWP3rJ8dTNdZxwGS2hKFVVSu/CbtmLXmDAbc1fw/+sXnj/WLsPHE3wjDN6FWRl
M1kDo1gJNhen7LZU+sa0jZ+GtUHm9KsUit0LTWA+jUUHAr636L7h77a4lQyE72sf
gmWk48AIvcR+JeklyZJm5hlX/KXWUH9oW6rEOk9u0Qe28VkxLTuvO572S2DIJZ7s
4xqVEeduCR5boSmcFldpz5ZoyzwBRUOgr8LaFjQBxo0KVpasS4XGDDApGAOxz+gd
V7wXKGCxuguNsuNmv3t5BvWHNLJvEdd90dNJ+37sxGfOaIyArSiUK1z0X2VBLUeK
dN8BD70wc2vhZtOTiBHgDqZAKiGgNPbPVL/P6FmbjQKphYIKid16ReBjrl2T+0Ql
f+HuknT/6pls/cGobWCmd+gVyVgOb7QiFyI1lpZsK9j26M34f3yc74VmCNOD7Sq7
AgGymfz/MS/8ob1LweJHk34GXVGqBYkKFtEj6H2xhUEtQKQJaTrMuWlBa1jJ5pKQ
oHvr6l+PIr1XN7cOAk5SPYC/NN5lcsBI4Qg117UzxBrY73FMaoXaKNmi3PlNieTl
HhCpidn9wEChKIbQ6AZfAp6x6U92zYgEpcJazFO3vEk7svHhL9n4YB2L8Ef8eSMw
2EMSCV61f1ZfMJgett0FYWtPmgIKQ/NHvJE9qlb9uYe8bldNXG603hAIAGASUib1
HwD+VCV3QrVKtF0z4o4BLZvklx1hUtExrOgBE1tt86wTrzUMYauJZRbIKlAHgEBU
aTcKn4o7XBeRT8t0/XmQu3WxSlcAF4TjeJCieBvsh9abELzPJl+mFNF0dFOF9Muz
mHnTjeY1g0zhaaVdYpYVjR4BeWe+E6/3vcWePuCI0esmeLvPsW5yuKLcBogvCnps
blPuP6bP05otyAwISlkPoTtajaUl7tEagkvDAJoxdkJfTKTRB04Y+UDUg0J9CJKl
SshJVTL6dGd0smn+iy13+k/Rwc3pBEzVO0gYVbbOm5smlk7E3J2xunRbWD9r4gdj
kyNLvdvC2QZ7Scnf/kVuaqusw2Y4S4l+dDCoqqvjpMBkfDx7z+xrwEXLUUbZY66q
G72fH9jBwxJpgstyC/zfjgYTovJCB7tE5l44mLVadAOdo+ULwv5GYuwKBbhhfG+x
1xaQ70jY3z3LQiu5EO8M8U4d+ib7HhW+Q6JUDDA7aPG2dh6OQgc4V/kREtndgMM7
UCbthjJhfbcVaojSyb7LNCsDA7LhguSada8SJ5bKf+mk5MtUESl2IEzApEmQY2Z7
KlsrqfAPgfkfds/YXrH84Tl+pSCkPg5df1pwT7sBfv7NV5g+ZH3F3XderUcfuZ1a
ClPAyCNjA4mD9mPuLfgRRYJ/ZeeoItKR0rQbiYsamqsIHXmmNIs93ZC4xBQc7tgb
NpGu3+fJQ8hIGE73lumd0ZUqXuvHb78JX9aFMxxQbhIXaK5IfFo1MUkR+1azSbiR
kAG2hR75niM0gOT1v6F5GXUVr3aPk8KDVBqXdhgq8myEglKxdmOrD4xd8TZ6eOuO
rbx/nonNhJ3bJ3vdKNNTdhV6HKbT67c/cs2FdmjEiItnrMgKKEizOfXlkAgRZtOz
Mwdwlx9dYiFth94r/vCOo9C33D6g0Tvw2Torfya+jfMW8B2FNalW/pnJzzHqjxGR
I2oLeS/m8nriYqY1tNfwrO//z+1AzeH0nG8TVuoBVWuY8THgMVxEn35zKEQuxMXa
6GaUiZp3Z1qpnO9/po2fr4LN4PV96rwDk0fwgSkA0fuahNWPQuxIxG7FNmLxy4Eu
AXVbVQOLEzjBUWcvDL6JUXHmUFc7MUBPp1mooaJNUGtRvoTTiEH+WHNv6SM1mKC6
4HcvX+zwfjMvb+np8NjbuwygGZXuOprufSQAbsgmcP7MSZH9C0ZI57lI7B4qCykI
SCaNK03ag8Fxf7DgybC1zF4wjfFzdDr316qw4Qdi4wocWpPe6ji56gGXT79KWZVz
PvdG3WU/RZJOMn3SgnADTNgPijXOC2Sg4z2EDvY29PVuly/N+s21q62dUfO2ZhT+
L4CDFEmYeIR91XCl1CuAU7XuGvuKKrqYZ2SgpfufnKhjF/OBkRJ8THklV1s29NDq
zBfqHGHl2iAfb3WSICHkkNCVFxaqB1WwtjIJ2+FZR7lFQENP+dwGM3kOiddXrLis
5E8B/wIp8kA8XBwHbQoYHIapo5GWI8X0mVbo6N5XCuDE6fFLqBFzLqT+LidMiB0y
P+DBZXDRt4FNeF4VS1xCfBW/SkVE2N6gJEXYWo+r0i/Ga4WGOgWV+qA6BqUeCn6L
YS02S8PvIyLl7LfKuIjs/PQ+6tqYqUKnHMbmZTJtuCQA2M4PxKSkrQiHB4vrobia
KXEPmgymsgNWYLhAUn99PED732msI245bL2T4cGtgd40cUYAHOp5UUQDArZGpeCd
2/DU1QkZeBTvt4f+9wWiiX2XPJOTdiJgu46qR8dS2Id1xo+JcasyXWRHhfVzhHUl
gWSzUYAoiMWN1lkZXfLCC676cjTiCVbugZJIzAwZYarbEImuCLUAP1hVLOFuObEZ
CVS7oe9aPMF+VrNIRW9nr2NMqYS4TXKtbgV1088qdPL/HEN7laiGGrc18F69acC7
pNAPd8d11Una0wa/uQZORFfaDYoNXULbleDwQQaGrWtP172OP35e9EaQuLx6PrD4
xWuvfKfhaolrr/VRsQH0RE1+OJBmq1xL+0ADm2lNc+O9byciRTQ9HllEcjIg49Sf
ULY5l+1ofim7N3JWdfzWqXf2uZoMD79j+1OO/gU/y7eddhDCUdZZaF25z8JFiZT1
qNiWITBQ/wfDew5KC9BM5QMqqXfAE2DUNTig6CRR1qk4NLez6fcGiukWZOFmf22I
gQOT4TLC6JTgBc1CJ1hog+B5qgXm+WeyQI8+ta9PJxbysSC0he0+tbFZtC2wPSxI
w1YJbf9masNdz4cFafhz58Kba8bJ7MLip2pQkLW22LbvMl3pXc9Kdckun4LDv4La
wr9Xs0T+TO2KvvhJN7WOR7XwhRtfw/jR4r9GFTeg4PQQPXspGyeLqRrpyCDFA53K
kWDsTkGI/5kecsAG1DSmwGT4EQMTii0C7n1tAxojsUoqm8isWV/L6DjGjQ05geoc
BlYWgwIPj2LBL1Vu3bb1SNgwAKSiQZPpYB1iVMQ6Hm2HurZcwaRcUKteJrOJhZGE
k8MofFbdXhD4JsxqIx7yEoalWPipoVDicnkU0ehHe302zKD2AsQTQvGdbW1XxNrv
7YW9v+7dKwEdt4sMSWaWurPjZHD4VTlYmoeFp/YBBYXgiS2RJNOEfjT856lr7YNY
V9y7mbglvFMZwY+Et6rG4cIjTrX98RJkK1lEqqqzVRs7BDa7XcVlsCn0AqPDmpcR
p5nTYxm4dVTZtbWmzc15GhmWaqW8sZ6OyzbHQfVrt18zhP15aQ2UgNLITlWpxJaB
PgPjQw7tHSGEaz+R5hP5F+cCsolR0yfovYyXOWLsGVnMmRvofWGgC6r5maWbv1ig
B5qLtHGtXpcXQEQmYHl7yryGiIsJ+9Miv2JGDodvuyBT59H2EzOZ7nvnFCCti005
zGnyu2Nm3jYzTS2AbOceiQsa43b85NYwjquBlqGfvCWfdigNPREKvmWmIFD9mVrt
okEAFZt1nOxpaNV6jgccGpDlaZaoAjKM3RZxYPFLLp6JSboixpGw+87FkenARcv6
XJWMs7rr0O2a/vKGlnUX9NBZ5wfjdDDl7QnUKFRCld9UHiQ3oTHwRsZTU5MdEv9/
b/6jav3RRHwap7kqP5QGWLXNVtnahwyTuGiI9vdUaCtRg9jGGrs9yZWCMl6pAOBd
GrbyPH0qL7TGdfr9MiwF+Fzc4eTYT0lUxTRRmQPZxnf1ItfSIdADZvN5JRHzP+qF
dmE/FfjiKC7W+ddzMQAgH3tmDrT6a044+JP6SpidwOK6yir7H51XOumvj2NtWIay
LIIMYvPhyyGujkZ5ktURQoF48pRabNwapv67NVpPnRuP37ui2ToMYl6X5ucj9Ck0
4825QRQPk8OgAle007jCcGuyYAsXdUEh3LhRLJg6MzummwmE5VA66m+83oRPX9Dp
GTbf/92yvivwjwYkLy5qmbwkANxX175rLX6k4BHhyhdVIjFjGchlzdsg0S2FBdif
Kl11iq2555nY09v0Ej5PfS72TtvGbvWkxe1x00VBCe6dc8zh1AXoKhFYRUFqJOge
VSe8QRyjtl55fYw3rMd5RpJ292ekL2987n2PYHGdZvywZhvdkUksxowQYJOsAlDZ
J5r36xyOWxQJt8X1PE4T11DZMxl50xXT4RqWOt1A7jbNuJE/VwUNI05fsgS/RQr7
3m5UmGOw/GvrPwFnBiU6MfcpYeAqfMMyEPa9F6fkKyuRQ7KmyDwRfq6pMwRPdPMF
45N23tOUMt3GLY+cpCsUtYEwQBcMZctzyztyNR1DpAA98bjwXzdxj3hjymJYX/57
evHAJdQ2lwlr8XoNsRXDAEfK+Q5I9+EukeFryZXPBZwK5WUhKk1WK/PfHpj8ZPfl
b9vVoLYrWpXnK0YTg9MtaCsuuf2NBFxnGIVeu76tfdj3L5SlGoxbyo9iwWdZTGrn
s/K3PlRhoyz/QRODzH807ngxz9c1+FT+2WvnTWbvjWSzQE5gzSBc8N1n8Pn41GEL
bbV5/paEjqMbxv/yhZ3zZlXIfvltD9kVmiBazNFMhWQLjtASllwJ/I8IuxRSwkur
gWcCHRWZhvNOFYvX1pJ661ABenUdLAP7wjlToLn4PXi4B/rUI3E+qOaCzbUkPmb9
YCZmOSlNkQqJphHVWVIXc6we06NpjzCnZZWXTnzB3UkuA2P8y5lLqajByELW2I+p
uYFesvWmZO5hFkVhQxFX24sttaTRCnYuJMi6L+S4A7R+qbnNcb6C3UQhQACSgRwO
uGKLyd4VpdT485tTjicOh14j3wA9yiIXRNFyOea3YUY1BfrLRtfa/vdOQFHGhjxy
22RwIy4/trHynyrEgN7lKGh0Y9ZtSWcndwTsIwRJsPYj9wvGdlwkAb9tQi6u79F6
UVMGdSB/1teECBDviTuOEJ2mihFcv5geExwRVwiuA4o2CSFYjjxbPkl5tFIk2+qm
o9jLm25L9evgx42Ef61T3yLo6G7qS7Lj93aUcDZVNGrIEyu4uYBGBOt65FJfdK+x
2b800/VkUIQVR1ROM/cU0giE3ECjBBgIMlWlqWbFws6TdvNVpiFS9Pd2uo3kR9sB
FM+XHOkt0M9t+Nrwl1UwHkMkDNlpGdOXIn2J6Peu0v4yD5/sMfggK8u5fRzSRbWK
vLUeYRKa5FQySedokmJ9M8gKi2ksrkVua42ArJ0WYL2ueATUth8jR73GczamUIjS
xKzKg/SpCx3rgZ+13Y5aLLVbiOZgAoEcg7+E8NFSyqNMaF06zerjF/6aBvtNRAPS
m7G/AB6H1qMOGKN9pY7vJMlV/S7wphDFtjHzB0VV9ETuGPxt/zIq1wXX8XDr0NqV
xprXoRO9craXQpswSHyWKerf5BTCfqWjyjn3gzKRAPI03XpZ0lZMLjUpt2TmgWwo
lL6+NbiEOhTkrOjdqvL1fSt7J+bwO7inDgjwgHIzfvXzSbVBE28DLfOcfqS3ieYs
I8OI8ayiZnj9p4hvh08mEL5l7Zwu8OZ30Xvi/LjPkK5fIaT+a29EA3+imXv7QdAz
YvQsdtWw9box5OiicdLEucZWt8oUK+uUhpMt/6VaYduBedtwCkv+3MjP2QXfKXrI
L8dOhSat/qzru6sFiuTH5NfV5QxHWCVjpfRDKqtvXpckdZ7mENre+8AWAA/kYheX
WwN5Sq6ykx6GirRECqo7VfDgx1CHlKpwvZTza/45mwYenhaA50J34i9jCMci+KoX
T4PutCJ/JiSrhZjiVul/sdkqQwdMITbKtt8A2ED3dOjCaHP5/B1Mj1gLZWRgjdrN
7oyU0zJaft8y0XW7sbDCNp8nru4bNN9mpOMcCAmluwKA1nDXn+jw74winqPmXq0O
Qe1YdowfgEZCZgaZ0gOX9kj6IMm1o0wBSWwz8ehm9Y4gXUYLLRGnFDF1CsRdj+dS
wXvNiDXjuU7eeYUAW5ErGV9HRsMFi2T5sExJga2s6kLriU22g3drJqe52uDgyrMO
DGqi0LEbXx5HXudXpS1iDrBTojxjSnSXHgC4B+Eu84T2QfBafR8Is9I23dlw3A1g
kJDNlLuDsYuTf1ViDxi2tPTnno3HXqMdjQGZ5pF0VZsNyEys0JUEWYJiTDyf+Y6H
28CWo6v5hefaSUnCmzfdBntgwTf2RkgsD6CStERlHXaG93CJrDid5c5dlg+z+g3V
X2ad8L/MiLT5O6rQGNJ6x7oWONTJj2J3VFgaSyccq0SPYHSwjucNXfZygxVW4zvs
dkTtlhg/FVtu2BBe5pwv0/d37BTCDz6EFGGRvRdb1TeKpxR6egVc+HDFNiGO5xB+
rbazAeFr7TAh9FDg5FKL1dbm5N46y5l4Evaytk8aTuFXvYh8oguShYY1mGSXanea
pM8YExzcq5RjWvkYSl/B/eF6naupisEWLbpI9rswz1bitkTZphEnQiewaY1kY/uH
obVNZPCg+4/fw6dLMX5k3IwWoOVPGSIGAMQ1ajJAFGoUgqPzZL7KYvG0M18hFWEt
RLLxmv+LxSZvUWKIWiACE1N1K+v5w7Jkg1OdWX04nrVpkjsY0niGoVzixNbogtDs
raCvinJiEYHoHvg71pFNgyZ3BKC7K94pauTGLNR7yrP6ZPH5J/43dKkR1krDwcV8
oyGI1P1ZjRl5fxJWh0YJwj174MOUQyG1TMfixF7WjCZQvgn8uR1U0ugH0CNqoqDM
Nk9HOWNODOLREh3J0+/92E+E8Dv/9AejWmE2zM+g0ORXu0u6qnNIfk1mdILA5BSt
9gz+eQOC82B/sRP/NSzv7BHs6F1Wfeu6KhCIwPAZ2LC0FZop7TEFSTZKOlg4rYCR
OlmNdAGlE9n4jEAUvkGZxbGclyy7nhzoWZ6GeRqdBnEPrMT+eyNQplVvlruNXMc0
NnZh7r98Pt4sdciKB1FMQeNrW/u4gQT05TqefEhPWH6Xjlb72LPKwpGBgiPBXb8B
2WKWY/ahsXbh4V30ToGfIWhCFmMUBOkEgZOPQT942/znl9YgVWMYc4iOq0jPuENu
dHr33V/p5NzStNEZyVP8Z5eIqbmaMnxZSXhxxGMqdnH+WOHopjtEoPUMm+yBj+9o
IpPdJP/xX+8Z+eSEK4rebzBRdRlySEz1CK0WS3nxuMee6X4mSjmHZXibWx2V+quG
Ie0GDFCYlogOBYhlkYDlvpAmOaejeAUMV/swRrW5V86mfdaBduNzD3YSQM6emQmI
bkZR49NeVBuAnITX7ZCtFIE3zLgVszUCYlA0JhZBgJGabIdH1kRxQK5I0/eMyJoM
M1eetgzylK+/MGfOyzfCzf5QKwXwAN7NZ7MZI9VDYivTVkYho0Z45NqqW1n9BhSI
NArkAM6G6LSFiajLIpAWWxAxizZ21nGOJAm+GEuGU7JWT8fB6WIa6vYtLMrT/UaT
kBAS4gihnaO3/ST6wXiCAavQBhKNqyxujzyvarf/guR2n6KCloy/dif/RBqcd6KV
2rAHu5Rrj39s9w3tYQ3AqMZ6rt03omQuR6luxlXnPGx2IlXtmQ0U+2LVYz9TCN2M
UvdASreS1hVehIuOA+vdhum9Q6CezgeHaRR4vWUrmjVNFjacFDTrYfWtIxdbE1hO
XZIulSVMu4+kaXB/ogua3TZgkAPiwA2y1LGi74zgD2V/r9sfyF5MlKFTwjcz6HI6
gkxrJxnAzDZHHP+qOlW839VzTiCgTrVtwc8yx47RtjeGdTe7yGgKevyXCFBcHC+Y
OhjNkSY5IKBVnSPFbcIhbx7KJFtYOz/h3FJ7PbRzG7Obxlv6RacElEd/8ktjY5h+
6bHE5H3AGqpa/sQJSUi3iivdFU4HZbm9iBQ+wFuA+DwEs0dHoulBNoVVKnb5ZFU/
7bcM0mB+Y/OZVcGoHfam+P7xZD1OdZeYkzTdhci/m4W2Ebc5c/zjajW9EOevPu0O
3+2gCxzhumHwxLBPT2JsdQAGSGQPxSfjDhVPyl/eXIMDYTJbcjKoTKOaKKjZgFet
JXauGOke4wX5vQ43Ri5zS4rFM4vm1RS0KDBPUC585hD7pRK3Clpdg2xYYptgzWDV
Kt7WjzTvA0jTbEhDFfSezqWcW+CthQpZhosqIRX7/WY7MFgQufWYpc9c5FR0Xwsv
Tgax0gGxTM8FB5kBg10M1I2iyY6hKAl/xkRwWwXKXGkgXKEAKtK/obITfv81U6+5
EKhW6Iomm8ZHwft39kmqe7qwLJAKvDf1ZhIyc5Nul5nQ/k+XNM1AuqLjLfShNU5t
7BoBLOMq5jcvx+rZs6FeGX8hQpu70IyoFAUmGrg0myAebBAsiTdbZnL+cmcgylFP
/izeEiFivxBGOdEbTsQOA29c8ukhjcU7VIXT6qbgffXzYajc+q+6ihNpn2aXBWb9
UoFPut/x6lDiSqMY0gaVKaJWT7ns+GVAx0T+jmJwaWoqR3jkwo02jZ9ojAl0jCl/
UUhh4RTGDFr+Dv/uoOyFH/iIdYMzqgD6XqCry85gzfx638NyCNgvgTEIJq9v2cTB
TDmMA3lMlcXfRkr7o9RLEddv2d75K5rRovqT6Fmy98hO6MKr7KgCnKTvxohspRme
/uxS4BOKHz6rlVggWkIto68e5E5A8+jNSY8e5qBf0qrtEy1Ilj5QXSkzlAMZZaMR
TQ7pNB3mPBLEbe5fYjwHYkNoS64b8Hcar/cw2eSp8x+5MtDnuDX8See7PEPGs0gN
+A8WytyAhU7rUmerQfT+ezjEP76B5MIW06FUHUT6GP8E0hjZd2a007qrsbdH62PM
o7mmGTCKVMMtvbiri/4BqoDMdFWbITh0ByydPslOjYWELvfMVAdkVkdD4Ci+eQ13
/67jIdPkLsbH5kDyE9jZB+al2IxzIhkLa2Ju2d5DZVllEF7an9pa1if4rwmvGyud
E/73pRORJoA2Q1I3doHywGvPuY3g+4Npo8SbfKLWb/3OVHdaqx0PO+ezlYKc1oFt
NvE3OFcSLSU/Qr8gWDBaqX9Mkqokk7DU1n9CCuy9EOAF6PBeClvfxHGjZ1QE/B/P
DsmN4Px+h4f3fECAiNcBM19h2VxnKQoBI29YDis1gQRrT57pAbRAwXHQmaQpHzR8
Gmpw1qBOtzbBVoV0dpK9WoVUj1PjKiVx7PVjvHVEtsL1NO38uPgSiNA4lNu7DOCY
jjI+SV3fBZOi0G8F9ZeyiggzMY3FJjj4Y+5/mJ3djHP0AZvr1HWDT3fPpHua5HoE
kva9sBUa70dishagBXq/iMZoWAyWYmYUIwgP1ZAuHAWLjdB8MunbMxsGvEbqJ4Em
QK9RiTD/QqZ1mWvdEUzhjHkYMiPJPm1dgGV9rLdSyd8f5mbpPmSkzaE1Ody3zjW4
PkJ5c5XFfxhlWzhFrgQjz+2whihqpBpSCARzhlgI9twBSnadADUfpV+dA31Encma
jf8jrVQNshOseqllQx6IOPgze8d2T+HM7GqQUDkPCY+nhTP+QEkzU4S37h2VCGF7
+KPiRIcCTz2BFpho0gioA5N7SH5r9OIKameUW6hKw20klP8O1jWJixUPdAPc9qAY
f81zxabWKFyPCz0FvSqh/T2djn5MoY7ZQi6p3pxl4xfkItvYuSlQzy9v00icN6r+
l+lTdFdTd4OxCSgL0axvnRIDQnT8wml9cTd090rnoaqLM3hP/8WEJTb67m/IsuMV
I/qcCrGFORjNQzsPBxw0GISsVEM54zXaMUHHeKgL3BVuK3+utgLOnYsv0+gfWajY
g+wwX0s3x+ESieZmHe4V0dKII8zLavbF5g71uVmuMIy8ODXw9XoVRwCpF8SbJfGY
wJAecOUoL56wiNG+JeerfYj9QVswGCRiRHBh4cc60H9UDPEAf/63lVuOiAOLIIwS
YUYv3A22u4OAZPM7zm0UH0yVLWE3AdLZGOINNRfmqOr1URQ2DVpmCejtNNm3NRln
dJy5xlxCvNCZ5xR4fRiI5jltUzZJmVwMCK2mbeiVk9sHZQSyJbu8lvnBY247QWvv
ubwlpi3bV7664gvhw6UO8hNDGM2/RgpSd7BHi+MoX2T029LC0us4pMEhHC7ycEbD
aL4P/+YnWac3CCit4GKoYemccb9zRp8sgg2joJq5CubppStJBt3RTnvEO7lWXTMN
u4CkiGCFC74vtdqr+e7K67AkXSSWZOh/2jnsI9YoP6MsuGOiMyoTF7P001QGE6yK
9Pwq2QI4LzhV7oIm9bsuhnY9E5Vst+NaXXcP9MWLl8g2DWGOB5TOWWvxIxE+U2+T
BsfhHx1rLy/GFhEUnZ5eMTNR9g0mRtXtrcSyn/UlFUP38HPK5jU/E5fa6HpvAVO8
4XogHck87C64kK7bA9c+2Y+vhnKaCrGPLlWV5AkjV1MRicBjXWMxkfedhMjfnH+r
AQa9B/FVwM1ZMHA24NM+7v8j4KfEfwLdH7j3/hUUjvNy86AM5r4kYdWaoBBD7DkI
4qOJyIo758TGd9g0qxo2U6HhZRaMPibXILMIRsKQt2R42gM5w1/Mdd7iEgz60lSb
58GzwNsA7E37V77WFFE8LFNh85WwY+bHqMybJeAVlwfRcA3p+KTGzaDQyZErWBqZ
+uRwBh/DFiHXhLTbaNFPmV+ehe7yJaHKj79CRsX5c81CIjWNj4j3q9/lYhBirbOD
SPT+iWvEsp5XfGcTR1XS4QzIjkVBZ5V+90JoN9AwPQdVNHbSUCcY+aykTI5/WIJD
Rc+lTgQLCazogrMJEQZeTbx0Ql2nO61NegtsJodDWOU4kTCZSjckUEfy+BFTwq9n
zvP/dUkIemnR+UgGvBSBDRJyQxvsCS56O4xH9U5TYWxikO1Aj1ir3N2XjkosqjGn
TsXDZhEnAYBI9cdX+R84+nJ+Q1gwrFnh5sRp3k1cg9f7FXqbUhVZ20oHqcvQWRU+
uBnMQIXVVi09vCph6uzlYvbrrwyRhkE5Jf0Dp8HdeZuzzD7vt34YWvYKHoIZvicl
QjZTucGLVXLo+eP8EIy0BWXKyiZY4R4rT8Tm/JWVGu7Vf4t30wHqHCsaLHxLtHn1
+WxkD0tjXz4mewNoL6v6MvEXBX93VI2SD8rAU7t2sj9gSYC4h/iDh+wE+4ZLmTKo
dj7I1z148b3vCq3gK0O2gIy1eXV3AkgERHJ4Xc5IbSCQGGLslw2WqqVFyRXYCTK+
AkASeaxtfZQGNwCLZ2N7atoPfZkDcCSlA/KsnjyF26x9g6bPNC/x66WZWNV4NJ4o
6+E7GJ7mioVBM2UHlneaHYlyGjclLWebmo1aFSGdLHrjLk9J6ICe4C/6sFNaKTgR
/sguxhtYt9+vWpaAqvGK0b9X82/1GkWOg3SUhpmzEBt/6fYMbhkJ/B1BBkx7er5u
FbcTBiRXT9G6QZ6cvUHVrVR3IT9gadRNbemxbTM6/z9GjmVoRTGvmwdSb3loXzmc
mEpy30VapoAN8ZRAxTuU0FjINcQ+z51lXbjyssugW0fYVJEsaxsZEfyG/b1h9/qo
HxB/dNv9exlVFvCS7igH5C3JuYh/vhY3QrrOJ4YXQt2sZdh+w4s1srnNIgcOL9E9
aS6gzxmdi4AURNd9xYawxilKzOLhLWKfKVOcKAzVKP/wCFoVWJTIvn7AhiP+zv7L
oexsUPeEf2q6kNZH1NJvmv7wJdXHcOt/pyY8jbMT9hiv1VEN7ndeaL7XSWmJnec9
LV6NeALkRJs6qeMIFpbc7SfyMOrR6cILtwfTeulNpMFaBpeCz/Xj3zn0GFEZJT8g
2wLuNqr7oplRpkpWG56OUXTfAV+rV63spSJDAnmz6LpPZ2qMKNC6XLJNAQAu1u+4
FwIgwqkmA6RWudTnHtbhvQn0WOK+vOELSp/UbZxpLBZb+NzlbHeN9o2z5GNR55ji
e7rAh0lj/iMMDCFYas+M6r+0mhnmD6c5ZQ0rbEcU+YvS3YfCbt4BeaazpI2YMkr+
6gJO91xfDlziFEkdNpV6mPKT4X+7MIX7FK57AJVphIVOKOj8YLGfppnsHCxPkdLM
KSsBKyE0UpPDBlaK4LjNNt5dB+K9U9yrgjnvH/Qh0mNjGmh+sKih3imzK4UIqCMs
JcclxeSC7ruMuPexBPb8JonziWG0+Pd4Gu17fk52rGpLfs0JTvF5Oo25AhYZQFDJ
6/jHjtncigv4AGyENDEVmceokEhWS6XcUBT45ugWT2UqDLB8kh6kJHU+6oY+fxZi
Rx6RZqm6KMDzxIkr3bXXP57yeqNIeV33l1EtDFh1kD7MrnU5rcr8tmgKbKWciM4L
pKqebmRsiBqHUmgIkD3u4oVEJ14ASKcNwhm7U8c+heOLUnwR600eSwnsXyKJ4hdJ
K5ZAagh1GAGpzwEjW3kcN5YyZZ1DofLOU3Z+RxVO3x4ILeguCBYDzUt1LwxIgcLl
E0ezfisduNG+fMKbcfrOLbmK0e9ZO5ycFCVNU4Azmjv5ZIiOA5afGjBFE3EXzEFj
5lEcdReFltBldn9n4PahegmMBICCwdODaZqvcE07LVbdBCduSX0327U7xRHXyzPA
lDmSWs9On8dgbaggmDX3lXDm/RlZ4v1FbvGZ/xNmz7YWTba876obsipfHb9MqrCc
vKliro+n1RMIGTGLaBNGz59uYsIKoACdTqWR8mJ5IezOoiEWFKoZF22+2hbCW+EU
HHEEJXfBjOQ7YUZH5BYsXP3+EAZ6BZhB8yM6AunNo15yROeKFJh9Zju4XZBb3MI3
LOg+DgynevMdqZQ+qZxkTLC+lHUybtbXutSSBr2vXG4hKs5a1I3PLaWOt3AyBJt2
v5pzs018IracSnoPyMINWFVOlbupcKZWxZrBoRiQ0ak2ZnpBKalE6KrJaq1YX3nb
6Mh+b8i3ArB/RejWNMBIcjcUkd3qzB72f/GNAJIO4j6a6kpPCLAZhEjXBfnpV+XB
Yp+jSS+t9O2mykdiqWHoxCdcEKwjSy2HKS4PHchBrMuc+v9ihtM5RTtW2E2sfJ9F
ipnYY7l8U3Sofd56fipZPsZmFfdWiMy8/aslK8FdA6N036Pfem9aPUIas4t+Pofc
zNysaxzwlFyJx3a+UvJdDLg+5z7d+DclTuPr8J5arpeMPWGywHTrjPGktjyPaM4h
mDiDN8lwdfGdCFJ12rjfvnkHxe4wn20iKbuGaJylu8a4VSll44vHKMkVeqtak4YU
mvs2sjNMN/5iKUrWcb4c5WLKXmUeY4zbbQaho972jL+JgUL+dQKwtnOQ00/omrab
jU+8ITYnclIm7qkW8OhTW1t3Q3Wo/zNBKsCinSn4+3ZriLpOl1QiPyvTAR1t2HGG
Yi5qoP9UzXlfSzhc1OwzsjaVGXOh6+ocHSA61WszOt9CjHiMjQy/OP1fA6NJB67+
T0PfzOxjq5z+RXXhI5X3THb9HDCUI7XWDWvit0ytnSRrjC8Tkz6BN2hddkKpfvdD
i5FUpJVIsYFl9IRDqKyqMTR009+noxEAJqaqOqgst/OzvuGIH9i8tMcuAni9sIeZ
CNE4Scb9ViKc1Rfpwb+s6sJ56cM78e2S0wczK8SeaGnN1eh2phgfPzbIbCsnMHMY
otqvn2Eil/s5STMW49sA2dr0hckMB65vblF5BhJg0g1HuN1V7Hhsb7SbY46menw3
BnASgL1WnicVUquWxJGc0tEvCzOaW2RAbSO3Fv6vNZoMCZAhsUms0mdGMgatF4Vs
olv4if9W1/GRe67Gws/Bgs5DguNUEXrBbNspytbr4jdlsS3hiM5uRzs7m9hxG/Ub
qObuPQYdOeilqFUa/uDFQZkrtBmtWCbfuMZPXWTzwhK507cjbCiH8wD3tGV2qOTQ
lnnDNS1EAWE3vI12FDUmmnglxeV1me7oaeGih6gTzwlvBSKHRIuW9+QjbeGQlQ12
Rx75vubDpVXFSwmKdk3vNG4PZi01N8qOGR3EIWw/wjEth3z7jOExg1M5InsPON8f
5X2WUo+ZzyN0nwGA+FTiUXkd2B3DSn+B0K6w2kNFaY9iS3B0qu7YqlxS2aqdq5d5
FUz4Ly2Ts3oxWPaArEIQJJoc2epy/CFvHvupQoKwbh6+G6GzNwhDaqMFI+6ZpDDl
mUqf451P/XLbWS22WSZQYHHTQ3Aeno1+cGeMpRtgHh88PUO1ycW7KwJEnGXlrCkW
r+uPlx1mLZBrGTvE7kRnhX6WRJEuiB+Kn3ZPSVBkwFxd/TFQiAArY8vqEEJjl3s8
i76VfTwLa2IvnaiBT+L3IDLk2kSVXsUDbklYx413pwlDKroMvNYl1erXqPuCgQyg
XmgXS1M5gAdmBF8PXvEyQdlr0K0uraDl8ad+fgCdroz/nryqRjm9fTHeivOihdaf
+lLxW48CqWZHyI1wn410GhJejE9ihWwjVtvSS+xouY+h8Igd0btwQBkqJJR2fl2V
beJ2ecy5JNo8+oFM6vao8ITVrzqfuhstOvCQ9Fk9CSj/QA7jL/sYjjSA1dqLIvqk
5m4Nexq9FI1uLN6bZbEF75K+EDi39Rmw5zHN2VFf7Dtg+wDEfgao2nEV/QhFjPUD
DtG9vti6p05zyX3XJWEzEG60WeR5u9L+OAEHUUvBD/o5xeT9MSwhaYUalsa6/lpD
yFd0/St8Mm6Hyf1wJ2aZ/K9BNFs/Vnnif08mlQG8ecRJKooC4Fj45IZfhINHS3Ys
o8DP+9kGO3KoNsAbfHiYu29RWFgScUcr8+UnZ3qjf7itBun/tmYKGJKtthFWkQnT
Tahrs7UubIeqkf/bjZeMOo8tdu+52gcHRSJbGDcEt8LeEDbP4KXO+PMQ8M2FqgBj
ZfyLSzbvX0gbJ0tUOI1AB6QLYHFzW+mp7euTtibOU+2DS4AgYkFH3Fdjb4qwmvQC
X1Z/uvPLQS1HD9SRm5o9H3547WSOKdHhiThuedXTA0POMJ6UIb3ScdXSOItLhWSe
5YWTSmKazG1DNIWpiZnJyfeN/4Y3PedReh4aIMmJIb23HodlR11uwxxcbBqdnMe2
pU/o2QDnqybQXiWHHBeF/lwJLqJn2mJle1F2Qp94So7+So4SCX4VgaasAKYp2vJr
V+z630BH4LRqAPXFgrAHEMtBN1ByRkHYHEaeIf80QpVft+tDQY8eITiuvSSeF6jg
2cp1FVzYHVL2PBBUPsWIWw5WFmPQSxPgZhEpimb63GtgB0jjK8tXuKkaVX+zsN1h
q/A0PprTcNXO+Q5c3O/xyZ8UyN7CcqtPQxzW1Q61ySmVbSknJdJyxenFczDYqr1x
NtKFy+wrXHxzS3JKfFUFP5m1X7fTPfW/fki2RpnNJBh9zXWD+BDgADkLQFKuBVsN
5/jOYugi0/y+rjCgumzII4/JGadpnGAoOFamF3d9u3nrEdDNFU38QxK38eQuw7dy
xDWuLHaN0pri5UfnWCYRlL40r74+vdUmqg5QCBuFefroACIk8bf9hepYzsPTxpKb
WabKKX4MmH7vWbUd3XGFxPPAywi5Uj7OhQKXH/W4ekT6L0pAfTAJiIvLWKB9SefR
mVJwJR2sbHryv0+PLLsC7PgBtxnSCvlikSPK7nP1wDnNQF7+agPdPTGmsKoQIh4m
xIl/wy6mfPXA5tjyvoHYe9aPJdO7P7UCOqV84DUcAkcmDo6MjFjqnBQ8R76YBoZ1
/rYbhX2t4pLgnV5wf2kb6EKmr9Ig9xBV7vQEgnyJE7ZzIEBokiHPyUK7HkjeTA+3
Mb7rYcIg2ClGVkajJfTZKjSc/1ScJ6YqJvtpVYw6uUhb9QI20Ruqmfzk52JO3k+h
mVj5LfdtwJe/LCwMJM/uvOGf9i09nMqmEMWdJHKPt07VPO5+hUDeF5bIG0Lscby2
hxOw955/tCOxUR1OmHrHvg9Ju5Y95XiTY8TNRghOxNP3BWZO1oJtq0DLTcm3Yk71
IVJF5KU9URsHcrE65fxAxOD9E/mrWQTzQCY+y1a4JmsPhbR5grNcvo5p+qnqEHN3
zmkAE2+TOkUP9B2sCu4sC0ZxTSqvkB0x/FrpMBOk4Zk6FQFYBvCVuIRP7JtmD7rH
7wFlQ80354iiTMBWFFEzZOwwUkbniTCl51BiNzTf2WJovv5J9kYy+LoBr5Qak4Nr
Sv4T89Teo3EPTV3dNHpGcm6z9SW2OkYP3OxApqtJlt1E6vApgMj/S3LBWDJ3jbEd
J4lD+fLPPcSw9JBvpBNzZzITRNog4MlgvwNKu4WN2eJkV5TtPDQD6Q3tKash1Zns
7205+Q8f1GByPl6iFkuD70+PTmrHx4v0ep1/BGZ+piYBbzEYnNBC54Ew28HILmE3
Vh2dP5iUqwTZZp4eqY7TJ9ucseeAzKRjXVaAc5JkbvLlGI+CVtJuRu7SJK9W1hqp
sxSTVfUxlf+2ZyVp1hmXg/nencbrPJmuy9QS7Y98OIO5/cNb2Yv7IL2WwbNhHt9I
1iYrbu0isPkUcZEWoYBfJkCN4W4xoh0y68gCAQSXCXx1vVXxqwpZNnSXEG8T7Upi
5qV+c2IF2kY5LZX/qSj5Jdz1AEj6duI7gPOhnl+37lTBAuMFsgWK8DnqzPw2HGoo
i952NVRvR541CdjAszvAA+WGy2dcZRUSZe/AiX7Ocp8mjUK9p46ym4mXIuIuRU0k
7k/ZFI8JlOkrTff9NThOnA1H14QFSKXhsGA68l2LCERjDKzfH6HMmN2WF4DlSvRV
R6+savQ1lJi/OuCavCH/Q2C5nGgV++LXXTvh8nIdTuipo9ToAswqSnOlvqqZNeUM
zCi7YVwXQ+G0GDLI9Gx1R1qSsv6z+n6bXNSemxfShC49mNp014IXlUrP40RsakMk
vZsUaqi+GA2y5Y3rn+aiFVB0edpvQDTS+93dS4KFlhKYZVM9OGhOrGh7W0AiiEaX
o40oXFTBX1NWf/vtATy5qi5WMa+2RyKuX9EDRfduZscI3ivZop5vNraBV2vPxVDf
m5FZ/x35hhiyrCZqRuTIw8eJ2thTj837NnRidlKrAdcIBaxwFXu8omoCMU1hmb7h
pd+AKTCLtEw7PPQLbwY5aG3c9ZtYC2eJR9I1Vvk8NuvBAqWnldp8RZNIFaUvinXl
TXJiCcWjHi2a8nvDuMrqCNJTajIjmF8N6O7U7YYoIXHFspV5Rf91a14yvBqG5hp4
4CybJucOVTwuFFIdpkom6LO8iThXOxahzZZJ1tJ6fF4pQ3m8afOGK25MdQp16nOW
MmzRFXl3ff+r/LA0StzmwJQdDzzvFLg8wO6Qv1/JXufDVBnmpeUhbZR0Oa8YaU81
25AGf9kyCEsyvuOJo//6AbOwAFO2OQ/kVyUWI5Ra/VKL+5szXG3n42hgjlbIuBS4
8AWtwf8N4FGeADe0VU+4BaOC8yI1oT154v1VHt5ANWdi2WtgvXrI0aNKgC7JIwbr
lz7Jubq+Slsr4OY9MObrv/UGb/wHWsah3t7wJmuBEFcqy72BIW2Vijzqg5+wMafP
kmTEZjPgDSAeIVaQBvy88yVNQle5gWhx7hRCLzHL9CXdKZPIFye81hvoaULKZIqA
MvKZoTCrQ2Rx8Com9ztg7XIqIyl4DS8TJ9rel2Wb2O+Iufg0djGAvq79QtK4orQa
ZS6MVCHCyC9t9MwdXKPqsAv91tp/aN2P6ZgeH4V8XkufVbwKNIqzdvR1OFBmRwO9
Iyt54nxjiErYcXthp9ItQ78XKVEu0yDgMCaVGi0GugBQYil1MTdW0anG8ZTwAodO
q7DtU/TEoNQM0aV+HCipf62ouKuDiCX4R0n8xuhfrmCrgGN2163mn1APBu5ho2Lg
glxU/0VoM0ZWcrXTg3XWLndcxLpkitYCyOjSLvcCnVsQN1tyo5pc3TUeFdmwqjOy
H/EvCiVbYFRhj4L9lw6A98OUwK2m4aCEiA4IMMGXn0pe2NF+x5VYgRFhBqf5txku
Z5IqfEqnFZj2HpJgR04p8bGwOC4/c0S4pKarUV/X4o/OCHe8MgH/fdXfbUjxosTl
CPKYf2n+cQWZo30FPwdaHgM45w8OYXI3/rVYPWSM4/ZbOGpPcPp2sSLcBoqIfk1v
hhc7WBqCZyO4tgFzNERsVmxSuhdyJakhfZMqmj8sQzSqR2rIhmuGKbmdf8yAnSkh
xK0/ihil5HGbBFPbHFF9XEqLYw9ITE6D8gAKDX1Hj+Hoa/kjryhIX7mNvEGCcuUL
LNMbgw5pzGvAsqU6p0Kr6u9KwUlHN3niD7CGCDFZKWGnROnL50s5GO5C5ZcxCuum
TU4dyZOB8Ukne0gHM12PT/sEuSDK9YtQX0YhvTqfTanaZ355hW8Xg4F5T/UgEn9a
xP/yWxXGQJjhdXYZOXvTaja7TJf2AFIoxsDJCU0KfR21Q0iKv3FuRgkZChmvpf1g
ITI29xLTznzklx6OifnmsBSozF7kepX9cW7XA7XIffeqiRnTB47ha/m11WiQpGZ6
c8/7NHen/du8avQfKu7YFzWMMLRGYzG3uwuTvtK4Z6khp7mGz26laUCldqVrdZd7
0a8jUwT4TQL080FpItpp3FDBObMLZ34VT1rfulnihDnaFNf49nQYa3yGukfO70Zn
OAWwRk+2jcXAwJgpLBvUldVX2HLcUwojWFjuOqlmsfQHW+jl04siBbfnsErsNdcE
06HD3nudJQm9lAuXWIPs6VKOsiwh0XTT4K1AlXt7tco+UMaXKP7NfxYxjB82wmp9
LcnjhEvw4of3gkiEIpm1MyuDCyyFtDBHfFGXjum1P1ykYqQe342ms3SYhqyt+qml
Vku+hzMYzul6XsFDyXRzt0kqWJyIAwwVFxoccdYRSl+7/p0raNJDWtIM1q63qh3G
LPqiCS/9saqr3U/+1eKOMd11FjZ4RQKHlNFmXvetiX4R6qgADyFSWCRNnxW7MPN6
9IlPF3lxh8SQfKaSVDdt4qJd7kfDVRlfDGSK5gI8KtrqyBMas7jabvfH+qySBBLF
bB8uyVoeBxaiWuueJX/R2+uH3Rw2i09sTvDuggWX3in0DF89YHCsRF6ZPKCpDsmt
juFmKjYNk+vtLexq7sIHpjL2uMhVDX+/SSfa8sNJT/xqT4ORJ6L27/w5k3q0SDij
ISXWWQO2eh8k633WL+YIkQu/Ubo/7dv5JPdi7qNel67AiQnHWeEwXKKeY49urrnz
mN9XKc3isFJgPk3cgGRaNDGbJchWDBxwIT3lswWE1ZrJ92seZJNNWukZgmVt7jn0
nrOFqN4gw/TUMYyNrUmvsSUmfhFoBJwlB1hF4YNsDa5FfLbYboCVlj8p+9/M6ofW
FvuztLucQAul1YPzmdnyzBjw2D9mZwV4ThqWsxEeZWsP23Ajmze3wapLw3WlDRwU
QSGoWEW63fn51myp7j4tutJ/2H+AHHeA9B+3mwuSvl0RcZm8DQ9sAcaxunrQEtDy
X6d5i7NM3kNvpb+MN2ULEXt6GbowM9ESFKuIon1UFikIfo8V3FIWHuL8GTicd5yl
IJr2N8MtFProUNo0oZuYNeSgiULigifN1wnLa6AFpHj6h9rHZkFnri9+dBGEp8Qv
nMesJxwttfSGmZWUiUfAngbvKOPLcqnLWAQf6jjlScOzKbF9cRBxWETxIRj6tjwT
UXDSQ6tu+Yv3yEOJY55i6NHaZEtQFdkZupmfjx4RxKQ5mom1Gouk7wIqlkfoIWVA
O5OlFkvISxUwiympexUPfSRpYecCWgL5+XX+NmFUdNGQVGpAh8aBhH0i5ITDMy5r
q7jP4du0nXgGG1vfBfbu8sBhqSVMkpI7pReJ3oDOZ88/2x2586QYI3ixY0tQ/dlR
P29A9vZS68G/hjYfud7URj0NhT887IeATWhavoxbTItdG6KC4daa3p1vRHfKp7GL
XZYF1MkPB3I32J8EQmytyk4+Qxbir9OoaDjGKWfSyRU53hoiv3tJsXgOOC52wi09
33HQ9qd0SJBmkNINIBr5QAE01WXz3Omzl6IzXoLUZRwobURoPLWcafBM0pbX6Yww
R7xjDUGQQEqWKKIPtoAIjibKWcOxW9b5B2YwcNphL1iqnUrVCPxAY4+p2kKGhrBP
5KyCPS5ApV6m8ZPi5HKnPeWiBHtJ1v0qvg1f9r4IRXOCEzFrGzC9AykRZ0RUJC7b
+/vOoR9ExsNLdtDbQhlFKEIv7+HVizk4VgwwLNaXesr29qEMID2OV/NhoiLH8yf3
SxFv4sbkdzIk0XbcQIWJzRrCQOhTVJDolIgUBD3yFbzuBBGlvvwF+FYzM80oZ6XP
1aX6mMVBznTyz0EX8fyWSts0sBT4foZgqK4mj8KjkJ4I3RXkFqoA8n9bxiy0J1il
vgCgZHrFnlRFkM8lOCETrCfbfrC86V+Y7JMbJK2HTG9rsXgtDarC9zxeVIVBycoa
xZP5WNYkIrDlzmIR8aDZsK2CZrqiB+mxg/N15FJwBKxkv+nAGup/355hhP8rQmH3
yH4IqxY9yJOfvMsGSLbCg3TmthWB0bqI4PGqARxeRQ1qmBb6oUr+u00U2sG/zeT7
NzqYa2u7XoOrCJEYjujhXOrMy7uf3ecnaXKF75LVcAXs1TNOOlj13HYpUIhTI5SZ
zcfN5wyGWdW4lNaZ1JIGdrEfywUAgAUQbOyQU14ornETOnasatD0fcIRZF2jmROM
C2d4Ar6FlL97OvIgR2hAWVytDBBAgDUxjkl+YO+vY8GHyAWoIXunuUUIO2NMf1BV
MMlGDnc4DPI4SAaCfDJigkC5dwT50VfH0UuAvuBEJ3V+yNkRmnPVCTvo7SRQ+nSz
61JGBPQsKR693PXU6UVjKqBfKQIixQz6OA5XFRBH/chATj3m62iLfDt15Kommmcj
PO/wY3ax/5cLgb0bSQw2vdGTInUNqLHordNLqZzchOJ2A675qq7fKvHsX71c8flA
8JJolVULFs0hN58JhIeeT1yTuNurEnOR89FgOJJgj9RA9iT15QLCUOU9eWbYWQl2
Pf/brOEbxH02LJrjEDoziBFofi3nwr/fHgSvAyOSoCJeNSMb2mjLIU/3yASP1vkY
DmT4v7qrMUIy4xCeLxc7Zw/2SgkHWfkhxzBxLw61R3rsFvYn5u1o3neuELGF6zWM
R4CzgHXgwcFO9OkY3FIjTWFjNTWb/+J0lsG0pEGuH9IiNigGtFC2mbv7qBesdlqL
es1pWloMU4vIu3j6vf10h6jEb8uzJA9xCq87l6MdtfZq+WSP2zSrbQHJb/4qQOYJ
6VObLcJUBKAtL+MQ3xds/Rlmxli3arUk4G0CeesjnYXZmYjnaQCNxknumnuB1jiT
Pn/F/sDM2EXJObWlQtz7pnBk6uixMzzMLf5jHHjaFTSygjYhE0PRuVVWcw6tw40W
owUREUxhT+wLvIeEjnvJKrZC+6ojz72xDhlg/JmpCZqEfh5QBKt7ogF87HB+FtBu
SdP3dLB6NueXFmCYPjuV/SmqgTt0LTOIyA2FgcZNOTrLbA+tOTWIOLTXf4C+DDEP
QJ4lr4yt1seGs1YnxkTquKzv0LFCYbKVHBxUgxxj/oX3uJFaZwM12HGdz34/xKlN
1kjlK5QUKKhM8nxn5SkGTawDUz9Z7Yi8hwm+HMr+h2aDWbj5I3Vkoqu8quOEH28+
ugauuub7z0ojxdPuOexaIqOVkQcbgrm+Spq8DpG+u124iyxJ2ckz1hzUuKhplcyu
HrhGMIAQ/jK5GNZb2+PJN0Fj4XvCi10s49EKKUEYGgo=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dVO3SJESvOvVwrhd2p32U0iZ6nL6uhEidxCveA7naffMbXZS1l8W2gmDnUKMxQXC
+zUlnt2o4tdVC7JrE3sCBDfmRlvi+lxoo2pf3RX9pKUgIcjHSkVKgI6/u9ie0veo
Fs25z6fNu9Gy27Jqo2I2L4G6X0eTeqY4/GdjEgFP9BN5pN0SHUGYfmfRVFRp+ABT
0o1fqQh9CgwyUnKdj35G9wXvR+Na38MKI6J6gtWIbs1iJ7OmrlBz1l7moUxTTeoh
jsLY+j4onthluPc72lYI3IlRAbB8m83CgZsOtnIZpMoRe33fCf9Hj8y+UY+jGxso
Wu3BB/qQpJLDwBc/vprm+g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9232 )
`pragma protect data_block
3q88htcuYJYA+3w9pAqjJYLPgEsAPXUGNkG4ogN9G9McV4VK3PyYnS8rYdDfedl4
u1TWVisGPX6tYTgQm9t6cxg2n3+9/IImVa/7OGzq7CYtGjRXgoCMTBY7Ej35rFsQ
dkTzSG10QfCyV00rsCCmtlWv4LkXK/GdL5c5NnaTaW4jBimnZ/KGhYNYLPemebz5
0fJnkIUxURovaX0L67bxnNoGk5MclunGVySo17pjUJvthjQ6aedWt8OQ9yIIka7Q
juexqV4kpAlGM+VJ13m+PgJqoEx+3YLg7aBYuOJWJWNXe8jsfPuzfvJFU8wJFlZc
U3GgWcYHAnaTWlAn3xAlE3LqoLYpho9heIDHXC5VR6g1Uhsp7P1SSRAdaLYj5YiZ
LF8IOY96Q+ghUD4qJd+ufW7bWAMI6a2NmcFr2twnZLWMFOMdtI9yU/heB8z9TnR4
PJv5r9TUrJOvwqkuwytPgO2xnVvQ6GKz/NpYIz8YAi0bcB1G1ILrfk0VO9T0SoEH
F5NsoguY6vtjcJV1qD/alvENzg+iC2I8eaA3JbPxyYnubZj3Q9Wp9vEA3gIooz5J
7RjiE9EzhxcCShxxj9pPt/pKamYvPtK6GDck1PFLNw/mFOthpUbJbzgtnRzh/CXE
GVIEX3KD0g9Z2R0i8Z9pGX/WO55E4CJ0Z4haMb2SLLr9LKT8Jl8t6SpXKfgiymoN
mhwx+aN26jVaVpivpstv8m/mZqGfuXW4oid+OpquVNfhWtKd4fJMibCzJRLX23Lk
uEig7HWH4ywHzwOGmSTHwGHcqZNjbVeQXPh+OcWtQT5ZSbCJE2XrSx3eXvQOBSbI
ehmPEFzKQs0p6ijpYkJfvxWu8PxLJT1xYFx/fVPfsmtLgH2d7Wi+QnxQQmBkmG9C
/TpmT/XgTQyqpivZcSYA/CVsQguAvooKit13BDmKz3xonxLFUm2lTkuYeqOgi0Bm
I++gBqHFlwXNQFDxfzY1ps2hspVjWHbx6bwTupggloBFQpiF3WaRqydHpaxoYFzN
t6WtuPwrggmP71CFww3AIU4AYwByfa3Lm64MQ3/6On8WNML/Z0lbn3JQnjgvVKA4
iUIP0HOvJ28R5GR4M8UVU7PMjNZ7zY+4uZu3sD1W4Esuo+EIRGIQ8gaZUWPKKIRq
Z0MMTkE8Y8DeatZT05iGBW5pi6o9IgOsMj1OWTxa9M68SM6isvH6xA34lijvkZsc
Tz6gNTXC2Op2xBemiA4QWzu+GEbvRLl1pUoG6X1udiMX7oxkVpI2A14uKT7jFOgD
uymrdNx5G2kOwymo3whRDkkobH1dEpeMlWhb0MtexGPEridP60ggij3+21DTW1s4
3zj7ggj6OvvlJuSG0ZSAi9x3XToAEUsOpL6z8skrlVswsJeR/Q2O/alA8FF+XMxJ
ezz7356Q413nc9a0YwZJLKCB/Fui6POUkzTyF3bryoPg6DGw7JaHtqMR2sAFm6YW
LD1LwJnuVB6ZtZgEs7W46PmwlQ1VHJdipXdJf7aIpSqlOWlQIlXOz5HFH6COYO5C
tcCmt3NY1poFdVPqnbd/XEJ2tShkvCNS77dYlxDoAm6O5tOiyeznZpQ90ZgcJBWN
6u7gT+hfHtxN8GYMrBV/lMnaaL8nAgs8AwD77ubTHYp0QVGq1M8suHMjkYxEEtjs
s5n2jMr3vtEm6elVQj26CAtvqQhB4HagkPnHd/uIvuhDZl59c3IEd87YmGMufIbc
KTmh1G8EJd6DZWFRrgTh3riTJ63X7Yfb/AQne68cU+CP23zPZOk4Fh98I0zWgqPM
sfxQVAUFfv/Xzj+Y+58/L2NEU6MG/SRp+SDiW2FijhzSMW0C3+7XHBxKuoMYtZyI
V65hKvRNDgl+1Uqfp01r1p0LKsDBM+krWlK1f6n5ox0mgeNelNgHc4vYs799g9WP
dZyjr2bY6L3blEq0Bw/QUrYC2pty7smWNt9u6tuRJDIbcXJO+lzU68m6I3+ue87B
9SFOFNf9aoiWOOj3b6VPjjA9iOrf+MNup1jHCerC1bwiG2lUigDgqmkfH32T0uH7
3HTsANXuA+83wBoxMO2+ZLonXl0PMPyLM+LF4ZvE8eyHKeNn/btFC8aBs2LdSgyy
sMMw3z3tFma/lHnmC2oyzDl8qY23X28KDX+4pX27glZ6NlWJA4ZPBmQr9lkAybVI
bm05um5decIVHND7dGylTK2YPhNBnCdrcyc+XvBilNmFff0PXys+nZnAd765AHcF
zFuSFbjvjd3Xbd2cnKl4pUS4DHRKmDkNGR0zgdLcb3adgfZa4Mujt9A6BJB2QMS0
wrJp5NjonsRR+F8sgsBz2vRnNnLzx8iXmViDFOCMP6QI6bbNXLhITqg+ItcWb7MI
FTvlWyCsnlK5w/q9MkOHZJo2NRh76Tpwpl4HJpn1iT5850k/vGEJUNpuo48oAmu+
NIfL7yPpuNhBT9BPoeZp560tF33AWz5zjng246PwsoMVKO+etn01rwmZ1TC96/oc
zoALH8h9FJiWDwafLAqvsQM+c/Pq44q9rqBo1bCrm83bNAWAeZUJ1OIkPlzOPa6P
JQxVZxSlP88GvAwuiBQWj3+vwX9u6Iwn7EuDyadzWEplze8PrWfp6pkkmSKMrb+Y
j/CjY7lsJshxEvVKoEY19+C0W1ls6WvF/PHwU93m4qjtlhwovXjxjt3Kk4zuWvJL
ahDkzas6+5tna0fSeQ1HsVXG/wqxBTwmy7AvNfwa2+rmOcys3NdHo84RLhxbMBBB
dYRdk71jickchn790gAsYq47KFjE4Rbo/K4jFyVzg1IJPSex+0ibHPCUUMKAWZjb
FouMVTNJDiVOazlifAc4dpYYAhyV4DaFnVSPVtRqpxvdFEaQKgvVctAbHehzmTen
RleY5VX8ZtJWlHWK5knEAgV5XC6HkIlLBu3qWQ1ZzOJJ8R4pqYQ77qsk2uMMKlwd
UjzQc4sWvoO8D6teixpQ8lnvuNf1N2yUhTP5pd4UmPW55iKY5tXLfmZRfVSj0uzN
7d4jzjGjZI7llbWjh8s1Ec69sm6s2s4K9K3O4U7X6IRASo3po+E05d0eCctRqadH
Kj4Hwxd33l/B1ny4Zl2FqmodAEjzspWJCFIL3zOhWTbXr5PpFu8/QL3/JgBnQVyy
mz1AYI/X8z5J3xAl5lZFwdcZfZGNrli3zj4vo7FtrcX/31c/Vz2xRvtlg6pHWUUe
Laanbx+qlOuDC3/feKw6Ej/lJssdx65CNwqQLWsgYiA81Xh/9I/nNbvlGMgQM4Sg
h2uYfo6gk+PDFXSuqceYWijNQ9jwowTMOfz5CF55pzqgQu13xTH1LvOpARspiSsg
uqHM7eeysiOpNwG1kD87X6yuledWlllj0P4w47KVDIGo6St8MBCFvSn8UzwQsEWq
5x84jAHhF1K+thU2yCjXp2kUo2XpDaZFNJ+M6Yccs57b11kizPjYR/C4Fdh3WQfh
r8KZBGSEGBbqjU8L2fwhmuY/A8bqOUoitzbVsUrk/4Gg6Sz39ui1oHMMlWqHhFUB
HN+ar/B8MA0rpgu3OsejmDBhR1vdp05feEBTe2N7I7VPLlfGUmK59v+n3g5+XYT5
STNIFODA4e1FMZxguwi8AYrJrTD3tVKsF9yJBk+cAHqZXEPEU0Obk88wG8ffAXWk
HJ1XkM5/rbJTsfGgZypmGevrr83gDwYYA6igAJAZhi1bBK7WPN3EX5Ijb7klJlcw
3n9p80kx/MC72sM+m4c4GZs/HHTARZBoPvaRSshme3RAe2x3RIxLMqi4PioaWYT+
FNfx0DUJag3Na0P2OYAvC9I9wWylxK2J/jOvrry7FXMEd0N+tgw89Ua1VXOgA9ks
fquLm8l8NV2fAsPByxZL6uea+BG25Zb9XSldN54dHUKjZyt5hn9AKHW6oRC8+iis
y8T9NZSgAeeKh5oUNdFEm7HTeh9sta1UsyH0TWkXRNkPltOpca0ducu/jysh+NIy
tlfd6SaTPhl+GSFpjXsucbnmLnSuFklQSjEDHwmnE7damMRNfJkjqdKArDwTKX6x
smjR08JrmhXDnJjpUJsIMmBKtcy6jIHwfSMTuiKMTXyGzYnrscmQy6gSB+Ljm7N1
hCYvTTH4B9qHLWKuzkuh7ri0b1VUgmmSsbQXfM+af4kucsuAfqmIl6xprR0S14Q9
pzJvr3wqVFwa5rSeYzpWjJ2+b2k/P9j9Z67r53jy4zcf1ZGHXdQXITZ2zxalwJvh
Ne/Z1uKoAIzSnN00l58qBYHHkRnJ9o77HCMsPh4xkezJOAvr41PB9S7axY727BeL
3fuic3g0nrzBqwaZhYpizJGQ0pkCTl8WFJKzrxXFkpI1oWZzuiT82NhN+KgJV9lj
IEV+EJ10zbr0Vcz5NxgUtR61Rj0slx6Pgk+AEgX+9pRmBsfVYuiA0sa4WvrGbP/C
RvbK2ms/5dSzvsma3cMZVMOkhKsVe9u7D0xNxmjUNCWfd5974uqUnCFBCbn3RZTp
iskVSKZf9LomSWFiSJS9oAfT7iQO/qe+398bXGN3LVvt/r3tlbbD2c9Ut8gh3I5O
0K8Ki4baTam1em42UeyS8EO/R1F9fk1GPUK1Yx10IT4k74smdVnc5b25mvZlyDe2
EzReWLmVxoUtq/cS3maMKNO37xpsO0gf+8DLUXxYdPrOMX254++Pdz/+MPIObdRv
JSISCNDqdkvrudaCNNzVrB0wqdBD72GgjTyb/TA7XqHWWZvc/BlBwGrLNS+LogNK
KbKJbVvwN1m76dpCwL9kX3UdM9P0mW2LhEnA5C5fd+uB9rBY2lgHe9bm6D7MYeiX
01NLNSvj2PgdcAUWt0F91BJV8SOVIeGdzFv63ncUlneN1zmuAgGs9zfgcU+HL9ag
OxDb2Njz+PZHS8pUUKX03zitLs7cxm5ZFy2zvWlH+ps1MRYb6CynRq+GcY57Z2mo
laE8s8FlDs545HQn3yicnReBR30nwtfs1Ydi+4kpT3cT1pbqqpatfFULiZGNuxnC
9xcKgaJ1xH9Itg10qWrBkBBzgAjR85GmMPmeoaa3yhDZE0nLXVl7nG+ezYG1gIOj
Elbg+i14kqsae3cnhSP47eDZDBFjC9TX8295OO1a1jxg92yJ4bYHE/Pqyzfg8K8f
C1XXSXInmlieXAlMVXB+laDQGld0XLLAp0bwVDpxDsLfMQC5RscC03gYyBb4HZ6z
Nf1Okb/QSv3GOBxizsP7UTkeWo2axmweVNzAbR7yNhEr1xwwr1ZxpjM3QB2efHQl
/EuEt5JRK5KljygYZYa6J+JRQGvDl4wW+1gFnuZWRE/X7lKnU5ekBzrqsUoWBd3X
iJZCv0NCwRx4rYQXNzzQbZ07HLlajwtOiOKimRx/OUnQGt+Fms7LIYcWMj0M2tT+
oDfSnwbKi4NW4VJP4iIAveGxoOs07cO9I/S3Bw4tdYYu7xywtHQT87GuSGlLm2wV
p5eMzUgyXSn1tRabKGRLRZTQ2Eh98uEB996ZACjRy1JJRd4dpFHq0XSovXZ9gidO
59UEdLxeiBZr6ac00bDu/RzW5o9SBkd2/LnkwjyGBay1+bZvtdA4dlBNQY/33qlw
PkrVKScQIxjbfIzoIHmUq2uWfecNILeHRp9tbHuiAeKlllyXV8cfoMOCQ9UgZXCw
4pPbNYSxR9vk84k4eI/smNFPuktEN45xiFzXCL1heln5St1FZnrL8cqEoa8S0jAl
7AcScVdljBXAqEcWfTN3NBLfxlj4ZP9+6VnUvvpoU2nIUXheWnyBL3DJ1E72cHhT
8JA9GxNJti2ipZKTV/QRkqq2YW1VKyGlpkq+8i0x8ozn1y4ELMyLyS57yrONDTbo
vxjkHPPrxsRwRbuqZx8G1h5LofI4nA57sZvX56eDUdlqsBgjR0Yh63Er3t9+Q8yI
ehO7dbGKQOKP0P1ugkXZEz0WRnOmmEL9ZFjEc85oHB13f/ls/atwPWjmCFmiuWRk
j9xQ4v4nyQ0DNRvh7t0xEm1CPNwbAEfdfGRso4w5dEdzTcJcgOy4XSSHN106NFAO
glIpgXEvYXuT9+iXmbiLd0gdfDm92eHtDXz6nn47z2rytX7VQAxeqzw31puC9TgT
KYLSighuQJxMpM2xzto+42KAbKYGBWIXBf4IBy5QIADLWsceYS0hJefcbxJG4Vw0
yv9thJ6bYzgulAlk0glbIy+DpL/3sBWGOZomDKm+edS4IQB0TMUscaCRqVSL8VIH
PUT3eHLSVgahh72LuRF3PwA9Wzx49l9gz3pQL6ElmugYnUPyw6yuRiWPBV5cwics
oIcuMqqSeEEVoTpVAJiHbyetz0C9Fd3ghVLZpbJ227ng9dPPLAL0DJaYLHl6GGF4
o3mzWo+F9LnL5iTOKSNfU3jXexOfzEGQISbJKcf+CV9x6IkTxfCxIqclWckH3Ghj
ZQVQ4p43H8+aoHcCybG/o9U8J+iRor+KB6mPvcObIymFkmyggLXQIoArW4jlFuFx
GzXTzzxcFCwWjRR8mtVHUVdnagnBSCGlrMFQmV8zyH+tIYvqQUEamSD5EGKnoamV
ZA6Ov8Crxvan6g/2rSOib1AXhsiQ3lPciq5ArYbGlTE0+YkG5eA80vd1WjrCul5f
zD9RZYOZ1dOmBR2IiqC+MfN1bVZ05ywaR4x3W7ccE2djvAnl9grGZjG3r989hsNT
0U45joDzuzTU3LMNyJY+1bAikZbF88m8KRvFGEx5oIQUe8gcHUaEnMCHvk4dLUdr
9wcYRkE3MZXLpz+bHm3iYCY0kKYPG2Pp3BNXO/fws6P1UTpgf4BxJ6+vJY6UAE9y
7kC2jHgknANRrHUB0tvxxrggUDbj04K6aBmgk6suk7JxNNwP/+yiyis/dItVVk1a
pbvtkfQXon4Mv0U57zKx8OOLoYlZ3/oktkgYmRN8IvcrTXtMLKCY5mZ7v5axoIaP
a6dWRlwkCDE0cvTNXQbTN43monwI2kVNfGX8yCcAFSa80Ap9k0y/OAyKYroa2j4i
ofu6B/go2MjG5B+mDFiVhbl9yLcP3i72LUd+GIS6RqgbKk/WBqZNJupNQRobs+Di
tJ7XSbddtTNivl8PDsMzVZJE+WOOT4NIMlZdBXAwFlWaof+rLLHyMyP0s83GP9Xe
5T3MBBpOhYcPCLChyXFgg6RVX12d9N8gC438uFwlu/PsCiLCjAdfCPGOPvAFnrsc
rIPV5y5ySG1201nKEX30mlvpLRZhqaX93u91t9KLU5DuXBaAAdQazEiAoAkwFkDs
437tX2V1lYOPnTyWcj2RS8QjyLlNeIJy64GbeANOxidD9FUpHpl5EL5y6PR8oDem
vPEcwWbcG2/E9jht7xeQxqkJPbIxqQKPAj7mCycOBEZRLL36yntBStEoilVTvzfX
m9uZAyAZTa866kU36qi8Eb32Ynb+504sTfUvMJF2JQ6juC4IjxLfWNzh2LHtRZ6/
yuRcLCkS/tTqzQ71mxp2hx8Y/TZ+t/FxnPp+8qLcH29mIa+mg71xeehWhJFQXFl7
POnduoZW9vbZRue2b+Y4IueMTmQf1hzwrzW0++NNCFRbzKvNWoB8M6Hl84lQyqFG
kxwrltVGAKCcJfQ/9TDGWWRHlmwkNzSX2l2EIGQJfrIcf+uZj/IqltBPXMgOTulK
tE/YscIzw2XuPKqP+nnKZFTTlx2QgeBHjVY3aqnzhaBC4RubCJBZf6rl8lo1SSF5
A3nBXidt28fnZhdd6/m7G95RpQ2Ly1aQffdSUi2aqH/8RARCuXHY0tgMT7nTNGS9
Ei0GL1gIIOqsKS0dLuA3ZzKuoA+FKPIcsj2/n1lQ2nRa1UTFdrP08cJ/tsCqnuHb
gfjUAx6+Kn86Fed98icpI/rNkHGYuKvMcHPL6OtiCv84r7m6dtI+S1x3rHHyoz2q
QRsc+opEPc/Nq55nfR6Fu/NAQ3ptirGF7Utomz3/5DbyZ/yWUXiLCiXLSTiwMSRd
Gyfiul+SMTBMes3I+lREW8Xcuu86nWOzJUq8gxWaopRJwimuiIWLM/cWSyr/r2T9
6RDtgTPFxRHVGMhPwrB/8YHVOgZdmWTQ6c/wYh3tJesUHoLxu0MAz7MOEb97k7pj
Kege9br9WZR5PVGY7TQXCWsEBiifac7GY5h16SYg8qU/RRrh19+bYfXrHqSyAVqC
NuZv7JG98ErvCXRDuzM9oa1bvugTLTf4q0rxzwCrABEDI8QjX1coUtry38a2j3OC
hCeag/3NVtt0AikzS69flQ+1NOLwQoumQt1dgTwHHfbiONJ2BTz/+g+Pk3g4GseO
sOoW9qkwca54daAQVpiRfYjZa8tqKBoPcKBO8L4xf6Ow7mP3miONfbGMCzyeuGiZ
btdeD4zHQOD2Ke1mTlZdI67XU0n6gssyFqKxXyIjXkKBgUXOq5QtjpfXKfrVUpuc
FbPsUIOBlVOAsC/s3aHZXyI1Lwlth3LL53SRI067ICa7RygtfuKwGdXVeZL6zWl6
VJ1nevJ7bR6VuR1c4sNcCP7cvutBBHpsd4fQ+ATGt5NBwBn26i0R6QqLVba8kDPu
sSWTz4PVayEKZR8+7pPHX1iddw4YdiapM67k5RhsBwy7EnteYtx1SDoxtxpTsRT2
Hj6on+Vv8hR1MOWpnJahjCWPdYnAzehsEWlaxE1JoWMD5isusEenEGUC5oHtiKRO
zhvyuzGsbNFZr1E1bNSFZGO9tvKBBIIrxVLKhE1TosxOtcDAzcefXmuDpXOTG5Jm
lFVkaWqyVR7lzP9lxctfVjJgChnFjoA3a4Hj1EJe8ndzYAOUnrtjrz1/03BTGl63
HvhVLS7fWTyY1jIGLhqcRFc2AmCAllTLtMNiu7mOYdKTXpLAJCMVup/aG3F/NKXo
ocJJWp5ShhBJtnDvhOnujIrUNkbbuXD1NwH8JGvy0KgWnJ94eYG6d1uCd4O1YTos
WRL1xetJ0n2DaJ4ILW605rOS0Pta202FqzyEbuNlvA1odL0jIn1cxognoyHbLExH
WXrBbqjZeuFrj31JiH0EURD+sJX6fpIpEtbf+O2HXeiFItDBumDBX9j3iz1jQEa9
SrGiUUfN078cR6+QJdbBs+d7wCJQ6yS654QOmoFFi9Te9XAE5RfsvNwPC57I2dq6
BWtv+JUs2FXJbbHgcD/rvmm5ceVuujOla8vlkmQD2u2XCzMqlwl5dgkTM9taIlvV
su4epPKhOHu4DxxZAlr3Foda/DLwShBCn8wdIGRLG1R8I97LLgRFb++nqU2l1g6Q
0ZyrhLkhEG6Ki2Neg/XUnd3MwOdUAuQQazIMPazPnFlY4TNBvrgq8AlhpE9mb3gw
DmHCsbKLftu/e9yEyW+OpKz6AIGuzWM47FjxqtEsNFGEvAT/kLvKm3TLZZwyPRBs
/IbzEqlSup51k0m6qeP6HEy62cROFLDIBcBefwnuSgXY4hpVYJxsd21X4F96iFht
95nMqfY8bf4gKkif6nqDrX/tJKS9LzXHY0KXMasm5QiMovVujH2Y4A9rXIME3odp
wpMevOow9yO6ra79fTR0ccD7huKd/aM61pitiq+VR7mXMoY53zmGyhBVvwGWyfbM
aDh3iG4IiqAFryIuI8oAbHKc0mVtwedPMeuINaFa7yPIqmhcSHjyv/5AdX+MrWel
07Y3TC3buIvr6HZz1Nh5PNbczvZVlLPrx2519r0720Am0x1ZSQ8yO+7yMAqUocf0
SvGBUkFFMb6GF0HNljbuBZvkSsGOFOmrstZXzaomhLPqy6mAAJs6SiEkthkYushI
EihT0lC5TVxpjFJdTAAbWsH/zpfDgLQ11qVwh3id649nnyKhbpE+qTkfG8rAt30G
4HjpebZYZvyt9wEQpGsFezAFuJVV6ZMWmXQIheSdiW3Y9hh1C7HaATBycVzl4s3v
2GS12RHA+6Mx3Qp/PETGFtJaO9v+BVE4JY95jpOA/wxa6OtbQ8Xtiry1rOfG+04y
l5L2olrCRS8keu1dkLOYdz+ekydxsQff7W1dBc//urYYR5X+K7Yw9+KCesc6qTBU
DBT33E/OLp8AbSwEwCL2i2rJD+CjeRH8egyRIf80BbH6SJJ7ofxonSipn18qmOuk
Dj0pcggm66NIzSJfZUCxqsEfHJFtf7d/vDDgXhJOlN5jPQpnpo0CT6zdylP/I5QR
8Ko8PxvnexUsHu6twTLvrRHY9mSUIiaj5YwzTINq3KTNKa2Xvxw+61kU+1qjflgh
bNS/qBoxdIp2ABQZkvlVLVtVb6OWkDZOrZlz1ysETHIlvaDmJbSqdfGNCc+dmXYq
Dm2GHUWf1+qA/QxBLBzi85/V8zwEkw8322nNIE6Xt/+rQdhv/km+037C+7Ri5Oww
dWuczsI6QVeNPwpRtE0+n5lT4lijziev4jX7R0x7Zz/a52LDnWsMQ5tAkkxgsbry
pDewWEg1y55IiMU+Wj8E4+tP7LehvoHLtq3fHoA4Dlie+By2kWDj3OnmxmZmCH0T
oydMi+aIccdselCF0AihA1N5ZrrcKnIzQCO4GnyaALZKiONo/SUDbPViF7nI9Omg
Z1Jz7w7uYq/dL/lfP5Qw9GbIpPDY5My1eg3c9/eH6aqRMkHAP5/BWe/pWdnd8XRw
SyUMBWm0O96xiBuB8P+Q1mVyAas1N/uHiUnU33MNt4gAAPn2uBriCiHEU2xrM60L
zUo1Sl7hp4kk4NoXQsRc3Zn6fpY5TNclXBvKzqMOzSgA1Pq+T9CjvvhVeLblb+nG
WgFzpaQF7KD01A6R12w/sRtRP3vXy1kbxgQ1dVIFKC9SgTV3UXgh28cZWk60K0AS
VJWM8GHpGB6AR220SiE4V2DobCJWBruz9isCbmA1SmSvdCVI3Me0k9en1/p63bkU
1GK004Ai4/EwUe325mpHvSmw6tOsJ6DdRvZTB9Lzgm5Ki9fTP7s+GzJIxcr0syZ4
TblUKxg6xH9lKAUKDKtQkhzhpDiFgi6G38rtbwn0nj6raachMEZhw+KwJnQTaJIF
QMekn2rAdU48zvAZ1Dme/EO1KWIkQg1ohhfz+RBbtKeNM1IzeS4p367GUtSKQf2P
gFbkOwSdML7TBEL2mRJ/SQXOtSSb5rM2dn+ASHZYj/atg9suYDzGf8IrZRaqry9Z
iMLfQWsgUZQhrQNPWAcSs4E8VJJLncY3S8nYf2d3t+jGEZ+TN8Qw7syNZVUEJ8jm
eDlYsMqkpQK1bf28hcjdTJhNlUW7VxjUJhu5sdJHhTyG4RVtBliPqqHGM2z2mVQQ
wYQVWsiXLIeEgUR7jk9g6PZxOBkniWxJPiFmQKOnM1KqlUvBWAtJVMarQuFNguVy
VGCC34rqaZRgVJ71EBbJtjp3AZqIZgFyifBv2qOJcHJXkG4jpvQEFP2c8v5uH/Qo
PPTMOF8lLmMc/D2/BT0XxnlCP4M//acKLClqCYkGGni0Gg31PMueOQLTcZSnos7+
Cd7YanWxsE3G2q/mj3RoBI60D6l6tgIhqDWPaXdedfRnKXEZUbMIG6V0UH8M3gUC
ADfxAWDr/59P7VX1AKsEPHx/k7UUQMfFLf/MxHvB4ju39ZuyX28+BDvGAIMkSKhG
nWL/xSCCbKOKpafhxB4XCOyiEC1FSBX0oT5qRyIUv8xI6tt9EHqzTbgc9hd6+HRm
a7PNomy6YgK2W8nzuyshMljiWceWkdwihQDLCzg34jgLBx4+q0oLOJ/8ecKWVnoN
vyPbD2SYu1asS60oKcM+w9Jcpstv7nOLQtCXcgty/f2ZBHICJQ4p5HEh0oJuYlVG
mDCuOVTllBPz73nXYQad6Z60XYOxOg8zVvTbh6ZGol3auede/ApP5F4JJZ5lFbYQ
A5NwVg/4nziLnKqazUjoAXhjdkjzGX7WJNSvijEjVYEAtD3nz5ngNEM9DF84aKie
v6mvEAaCM19dAmqWB1V4TgQo8GVcdQtjDA4Hb4joF5T00wYo5IGAPwEykwwHcbEA
9BHM97XvWM4/y6nFgV2hELG/HiHDQJgKqnkecAx/BYgh6qz1pghBvSmtyWyNK+0c
/J4ZBa+m2SuTqGF2mNNd830hBysaOzXtOfqrxIP9OYvGl7ND0rAIGWmMNVOcRYEF
89JW0qw73SAxcTkuatx1Vvd89Kn4y1kcGkjWJebvokQhW0qyOf6hhZgtkYJwqUCR
nq1XR1ZmBXddJhSPdj0AVherVA3XtDglxe6bky0Ngi9b1mNKH5KkjvlIqb7m5UvS
9ztyj/Oyevcib8qn17Kb30yXUJSsmlxVwPh8T7EKAJuhlpX19MQ9X937KbmuCT5l
TB7HY8UQyQp+8q1qo3lefLpnozI2jU/+K/mYmgghSR5gJdNVDqhz4/sAz3/wBMeK
e8RoSxYPPLnA4mDJ9T0IoQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
PQr88FmgrIc2dn0/GR/hWao0EjDxPcZ/mg0ntOJX9bDSNnyiwS4jEB5Nh4hMAdl0
luAsx3XdMGoRZVyMMWZKKOEWObL5XjZL1ktljUY641/4MqEu/gUNFMUFcmZWds9z
DaU19artx37DfctXvlclwPy/sB0z7/XmxGav6WuarpB8e0NwzKsVuoXef2p4ZC7E
EyeQ8kjDCIOo96Ql6euo2EhgL62MenL5Cq0jb8Dyiui4aBZ0lr35YGbFXl2mtIcc
KCQWwOtXqL7x6sB3Zqw5yB5T2SrenYP5Dz23njugll9XfieN/tQb8TXmTM3Rg0ma
0VpL5cmAJLv/+ln3AkLyEw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14640 )
`pragma protect data_block
UezcVUvUFHtTACu7keKUOJoBbA53pLVI4z+uO/1clNhLwlsuV3Xb0LC3o2edXUG+
kuaOzVyz+IBgXJuId1L7xTuJ006H+xddX0xWXRte+NVZYm24qUiA/YEs95D/Kz0l
fVsGfR41EY/0oGxVDNgZiST4GrfJk/R5Gz2Fh4XnItJPXlX61PsgiXvFURH3Xax9
Unub76OsWinBCsoN9YX4Ls8nVp8JOOxLACSEdyPGrKG073t96XEgkeYo+gAfm8q8
ULJrU47X+athlPTzWjbyQE2KMEIOWlZPg8XpywHdOSrseEQbw8wt4HgIJXVBbkT0
B9dz4JpQW42XfGnzVNZti/uVN8nvHQWNRpLZSDZsGtUoAr6TtIDRc2Ab92rxC1zo
C+GVI8P/AgJRG65lHk7WjvwFzHBShF3YPqhTRagRMK9Fh53RtRCrm9+LHXThywk4
P9BXGauEVZ41JXptkY/EV0VLLg/rlGHVq3B74AvPg59qashDXDxbIp7ZaRK5+0ZN
MS2L8UyZz8TBbU56b02g4ymJjUEinaquTzriCmeg5lwgy4f8dnGS2JkjJCLF5TXJ
+OnhO/tn2kE7YuKfI2yS/OSkkvfXQrCDRD6JNQtH5x0crB6cgVVhHbPUjzYavc/z
qUPylVGRRAMzbTe8inIo3tunYJnOj40vdsR+WPu7h1u5UHZX22qvW3wgOtzF9Qak
q/h9fAfZMWk6Zd2hjaTH6c43QnULp59OsVzsXhJIKtOew9lLOccgeqZ03F+Ap8Vq
DaVUmV2htTMJ/dphEThX+wm5Nq0FpsFFlwUQ5UyWLldBuTMW8WMRBw5U+fUQmNMv
Tm2IZw7sS/kpB1BaafMqJ9vERexzhzVsTW6rBSNToBuIKtOqPiNel9dLPYveIVkP
BEtRXcXrufsTjbc05eiH2FfReQPZf2GokS4iNyxhuqdH3VH5LFm0JC8Hk4kGWwHe
WLMq2vdbLukKJu9RIt/bKZSfFawPTVQ843HCjSKKHdjhwoyiYHGqOIR3nM71R0AU
dPxOZInnemTTMKERWfNCe5njc6uex/V3OH+r10rkdhc68XDZHQ7XjB1EOEEORCad
5l68kjeLMo8DqHjbtJP4wS9R/8yWlxz3fD3TBsmHkoYPx2Rexheu4TaOB1rv3Rt4
4dlAvQbxSBzc0t4XGmQzvSs1U5JEGtFB08wJmV/JY2sT+vMUnPfsLTLx/z1pgRqd
RPcBMnv/UEHNFuLfGI3lzvmnqA4CsdnqAvw1NCaXWE/w4aXvbx+WR9ZO8bmtk4So
t9GF290w4sUDjeCChmNpB/ia2pWTW96kGrl5qLygiHV8mVt6mExVhmT/D+lU+0KM
N62mj//b/Y4uWjt3lBhniORWrtWW3mAFCBO3Q0NyFhiNDhBfakf5xkpBTi1zxfqr
E3RwvCbq45Jlty8oWTcfQ5lUwdXvtkOP5w3ScQbXwDowxmzfPwcGG0CdN317sZUS
p+SktockkKsAHHQQvXZwKTihZsJLNbdQ1sBZEF01mFUpIij1sBOh4hwxqwy5mlPv
YHuMzcKMPtg3xJvVgKwdRU6ddIbzd0tw0ve0Z4njGcbm+iCmA7L1MOm+P1ZWoAcc
a0I9NoI2taXx257l6i3GfeuJ4wBpokPmSLMc3oDxZ+lW1lF/WfoiYX7NJaVWUfBx
7r6+AvvJ0AcjEBoczdroW7WdG8df8f2O+YVWiTosiTAF+XovzHhTqfX1efidlKMj
6cDMTm26jlwpAfFrAzAjFfKqB5NdJp9UP0ur8JtSUBTKWOrOch+Wnh+7iqknik/i
dzvI3/6SEAMiGcU/7IlzYIbWIWgE00NZ7RZcC+x1l/sm7XgPS7mu7vZsH3lvP1+I
yOBmBv6/54htGLi406Wf5+zqsv/CQ4k0Qntp9WCmyITZ8vXx5dba6pAUdwxgxxt3
YeqIDgeBrkr/Lvy+0YCyvlwfn+XTXx/vVaYSHd9dq+HeG1oS0Nj2KF42VkLmHoQm
JKsh7q34Lu81uojBDnlrvTQPJ2TIwqwDWEjqpJWY71vbRyME9tQkKzFHp9Q5E4IE
vXztLEl4qIcynXor26VEQORRvjVMosmS0rYe8CHh0kRbSTrpkeIhb4lKVdKUW3Rq
0JfsyA40E2xhkETlKZyCcVgF/kJWLDORKaqGMMIG5EACRg2sxxRnJePVUUNWZS6x
cgUo60Dzvd7gXSHEm+HiKpfCntHVaVWzFu1VwExblzfEIBsNbF9VxIr0Nd1Khqgl
eyEhO2a2rAcA941EZlbypuT6UEYfZMRo3o07VL2QaZj4P5B7R6yj8T4G2/K1LXq1
fu+jIZU9Xs2Sg1SZP9ifpHfn6nkL/BHu5/aRw+Fwtp2qxyFfK/+zowuPrzJaNeMU
4/we6ijPO8FcT8LydRsmoTkedJQvU5tdLQBYnuRWrslvUKzGwP6kjb00oz0KkI2D
/WuB03rmcv/Zbpqc+CaWWygUWPSgwbZfIfBKZZAZ9DbM+YhTzCgpcNEjozl7Rnlm
wOVsgyRonoEasQsjHIxDUFFesFju/m9JPyFiWdNCNiZ0mXxJeQKEA0+IAlV05Zm1
xqD0C9pNuY72gfuWiAuES2rcxr9Y44O9d2pwTUcsyiPswCYVdq5hLBPAO/Utoinf
3czT/5kEPqecUjvaH+paDgYHbKs6kfWZ/kVguPB4WvU2OJgPFOn6/e25VZxAZ9lh
sOW5+MO19wR5cxXOqltQBIjpT+zB5GK9dH4K85vHg97ZqUzlgFM0TN6ndWK4q9v/
Gywd6/GOQfz4WRCuzaEvYThlxNnpo5Ifyo6yLOFUo+VxnXs3EHjggxGrY9ln3267
PS/crs33SASRQAB/KCVLflJCV2BTi0UnXkkjnWP/ukuUJeHbQo8Txmxh6tTVTw0g
5/3gWHZwPZyxVMHCWKH9ZeI06Md5Ad6hAUHjITUYMiBanfsCRweAPo2p0IDMhpvJ
BxTNH++f7O5Kqwnd41AuKqhIz7EgZQfrHJw98kjYhD4w3FKMGtMtSiomLXW3HcX6
pUuoihNxBWf0/k8qO7mOtXw8T2a8bHQPVXljWUnHsmBqc/2qi3//skDMc6jkBuJw
IXTWwWslaBZb7yYcPwEjYn+EdWRz8Qe3xafz09BFENKBaE9aH+xKbO4Tf4Sjqmx9
VuuqtYgTvNlfHdqVWV+EXqqStlcQvBwAalYbwf2Wa+SG65D4RLgXX5L3U797tXpA
+u02CRdV1A//wxhhw9Y1MyR7haPP7ajhJ/VhNhOant6GK9wnqvL2lNO9qgzOgrDy
5h9KoGY+KVbW2fWtUTGv8I/gb+d6p6K7zxoaisVSJOUuBb9p7RtugKaLkDvORUse
qH/SH+vJkqrlv3ai9IFZ00dhzurknzurYn1Kp9WFMM8lvQo/oFEzwgOnajtIgd+C
vtniwbDM6hrPNEDbFIl3NyY+juHuS3iJvF3Eif+pFXEMF1iuQcib2Hj1SoYkEZze
tk8z8+q4HEanIMwKGKf8ail01k6MONTaLu5ijaXW3kwVakatC25mYbdLRzEnpCbQ
rdzPlvnT6X28XKhMdu7fUv6VUgNCQNuY8SzaqNHZL8P5hcaOBhrFV62V0T74rdGT
cEXjtRevIWi/GSQKJc62OlipxGMsuZIClzGFQokagyKPI8JKeuAzFqrb6RKzjgNs
mbn+YP0tY+k/oBPHJw61x+e4hGNuKKBq2lLp9vY7IuqYtIqtZX+am7DEZJD1YYzo
8LVpod3egkGs4WxkbE70kHQr43o7k6SD9Zv+UPMhtB/0kZ9+pvRYU/vrhjhU7ske
yxDvrvPi2v1m9CGaogSFq2Hio8TMBANbNHRsX2U1ZTbN1GQYTfKjV7NGsRMA27/5
0gqD818Yig2z02MHJbqV1fujsdxrCiffI+r4qTGvwpTCDizNqWKUYSqXuEM0JE1f
dOApT6VqRTVC30nJBa5JeZzokYqFXDU/3VlO9mhc7nO22L4OiwBjD6QgbRtP8uXV
JMkDvSFd/ZcGQUfmYr/XmyvzqHXbNL/z6RQcu2WcZlRdatmX6vgSstrQbreg5EcC
XXXtStpUUnH/s5QkW90XS/ezdDnE5QD/ueLbTs+SFayaqdj6hR6xD9qtDztBceLU
GqCbvKk26qJGDKddz8tI4VMVoL6H82S7nKbqbTud7OSCZ+mKxWhpl/QW2djbmKbS
j7yAGiaJoO2ClPfF4YNxvitiP27XOMiGFNa3+qJob3r+qzGvVu2zW7wwQHA/mOKy
AHT0oluMf4u71LpCetXywFZTMqS/ojRNWOUnENsFvqQ912r7MgGCgi5lYP4RhSEr
yB+Lz1lNmL3toADVStWsPC7IZZfh9cX6qAtnWqce1/cGb5WkPMVfLeIoQxMHTdnb
ZXCP8DxFEG3rLlIQgKmYGdIPdHBtEIluy0RfIjNa2BI8bJbDFxCmpIZCLRSfNhnh
Z0f2FoLQsdzSJcU+OCbNHIMGwXGym15v2MYBASwei5htdv7GSyhBGhRogT97+CEB
nkMC4ki0/ZFxV+nIgaQko8Ip7bVJkjszbQb4tyr9c0QNbi4837Az66rZTx2yvMF+
/ID1SHOqQpCyZP9SqIjz8mk4vizxLbHccf+FvY2DKGZ8ary6ivZWSsJzOKnO9N7B
ORZJ2jDYYbz3Wgm3v4tFpPAT0l1u1epR1xCmsWv8yYqKga315jM21Ouo6czbKglZ
8SWDC9nl+lqDc2i+jTG5FpG0+clxsVc63hzPgNy8lGpjLRLevs7xkyraIlfjVoKN
w/rJRHYBRjgX+WlO2uK37fRONZw6987LVdb4PP59S9lWi60oV2C+/KSQK0bqLhLD
Z0t7xgY0M5I2HLrcTABeJdNFpYjPx0jCLrH1e/ExlkK4ubVzL/39Tx0+BqVWf3jp
onTZox2Z5diSUMzIdwuV9jHdj6mxJ0s6SQi4uYF/bu/AABC47WCH+OxIDHigsh3W
jcugxXKh8zGSIU2aBfCcOgs3pmL/9b8CKFGkohc7CA50lKTHfYaso2gPBuOqqt2+
CDI8et9kQZkQcPsto+nJrACu1DROFGTU7sw3e/scwgPTpgoRLKF5BYND+G40LM4M
cRPrC3PAKBL9ACoSOOkVuULXf3KZFu53nurHHWunSYAysriP9k1jCe/FpT41paTf
pTncQNI7MvKBMaKfndAg8bqbsvq2eB1sXGtIjrX10NXomOhx/cbkuICWyXPIDBqB
tm+UO0ntHOs6JSJoLgKG6DCESd4pjeY5tewqQYcCH/5qnvAXHNa4r4fvpHCJlDPE
MvQ4zqLoAs2H6kTt8YmVwdCjRYjZS41uol+EzAlYHW46V1Xlp0ZcFi70mscnyaZK
t5/Gy9LQ5ZF1d3zHBTr3rbuJQkYKp48pboHEUGW+Tmb+hJCpqmBZHQW3u3VSnDMW
zPC1kYIemvCwKqxY2haWV1ispbrcMSDhlcXsqhSpsy8CYBUOX3tdP4bRlR1ULI+o
vcwJSwC7c+R4ahInysaDZgFXGVZsCPsi0oWcGm4s/ZOheSPwfi88QcdzP1oGf61J
jLt2/t1HVoa0vr1r1Afos6mbotal6gao5mUrFEjuUmMYbPaUVBmn3DIaOSDBl4ZG
yj2UGzRWe5IgYcPtuRlRwKeVSGsff14jshHsUcgxmj5jLV9ny29cZ1qbK1ebxhaR
b/Un0xa6wutFkgvTOn42pwAyIGcAj/vwj4FJhwzqUF6OSHR1rVyTxSKgvXPS8mkk
Wzd6rt9TALQ+EbDMyk9z7q6H8/sMmv7i70p7urFnqcy8h7upxrtt2KEz8yIp0CUK
YhQJG0OHHuV4MC0qHiraiO6UYZmJ0poYa4D61QujjcUbgVtLMs3xi4GYRn+S3kaI
CQQPUd6bg4z8vZGljsHaSki+O6okoc/2bSH3RYtD0VWweCnKJMNXKpU3WxmYLe+v
BvBbeCbjFo5uYA785qXcPQqDu4ARsize5MJqdmyKBtO6QAAKQMub2zVIwGOJY1Cj
KF1+3nkpyHQk1mZEa+0VfCmF6WfqrwBHHz4GMJst6JKIEzMk39zETRdXBT2kSbnC
sx0V7nxClFRv5ZMlyvzXRkuVak6cP4MXM3qEt6t2lX0hs9AUsrQUiCQvIwrgke43
k1MaXFGSPZD1zAb4vHvZKLGfxoYEfhsYkbTXBJpf0t9BWraqo/vJGEZpMllIATuN
6bU+bNYbfzrsHHLNMGh8RzaoxWyDidxRl0CgG0zManYJqfrIf2DjU6Za/91OISPP
Ne5B6lpeciAMXxcSrT/ASmKhSSeTTMWmdfmEQ6lwDZ1bEeJR1XTonVkD35j0tKSQ
oBc8j93BvamgTx2eB0Kk/OpH8WTsc5ZYY2wm3jTwSIdmJ9eOdSHRgj/gSDSmRWXy
8j2rQ2Igc2m3Oz5uZZyuCWKKn8nmXWVbQZOmpju2eC6WJPVdJ0WJKYzmcxTys1GW
B5y6Q1e+7wJRDgu1xtYv+Qt3TG2qAmJhlho91GsPY04Ci6eSfgfxP9RlVgmPyhan
fFroLMRaSd6nw4PsWdYM7j07E+XOTbHu7HDjeRIx0qq3FIIFcL9QLl+GrLlzxGR+
KnbpnwfeFqrak5VBkSWOG1tLseQ/qfbEKNu27A1fYvVicNLdY93xuRKFtP1s/nPE
Nyh8g2wCMtDzY2GmmyZbMBvKBgm24iwHKqFecPEa7ZKOUN4uRBntXbH9mKv7bUhS
Hb2mHvzpv1gpITpC2p37YNDoOmsiABTgXBOjTSbEXDe+E/M0LiDRc3uhkllMmXsw
qAztzG9qfthUDZKv60g36MTMuFD1rkc4A20vZktUJzqNuO5S282QAhURVy5c3Cay
DtxhQOUiBMrlRigLgWhaaQgSzEdHUCb0arZ1nbfv4VVRd/z+1NvQHCoBeC+atTBc
Lz9VfM8k5JRSXJa1GWY3HUdZrxZbbX9Q8nGn6NdvxPNKEmEl8KNH0+VHzFaSU1WQ
M95pzPLCUwzhkvKSD87zcGiAYMVnphJh7uMRw1WHVnUJmn1+b4j3fhXTxtNGxMSQ
8JWN1Srdvc2olHCFQD/EG4ONw9yuofFgrISmeGLyhXPO//HA6EkUwq85OHzLAOZH
xNVVGiVzEljTHOJT2m1z4x2XfXk+y5Tvy1OUPU3MyIx354V+Qk7y1KT4ya8oWcnJ
Tn6itGH4QyMVCrW5aXrDm6VwFHu9UkdKHjwsicIRiBhVNT0ktfMvtfIWD73jBFVK
MHBdKkvMtDEjlGFvJNo1MH+D/5XIiKxLqXaalHHvsI5m6UfdqEecFU380UX+lt9I
nuPbDNbzW9j1m+0Q14NkGPtBEOX+3tdfx0UAgn09ECDjr7//I9IbRlmECZ7QKsbo
FBDj09ovG1iJrl4flhj+c/nhB/AfCRUhGWLGTtHs/p7N2Fqpyg6diH5W2mG//Vwl
sc5IOgN7xBpyHRY4TWyupvfNlrDV/A/03XOk3sZ2+PkkpXbNMGo8NheImtFqZqow
d5s1tobjUG5njz/pAuhAEkFgKwtXOfntVQ7m4VWabH5FDZ65cpVzTI6n3N806FNC
7tcGmP+pyeJc6SWTWZZeJjUWl/T9gZ8jCyLb9vqPretZFGOauCxlOCIgJkqgrMAe
428oSsA/Y5f9Uoo2Yl+qIz4UC9U56bZYuKnv2K3+U0wmrafpmRHoYvjJ/z8YOKil
YReqCItxemW5LPWipzPcOacNwKqYg4BhFngxXxnPc0KMjNLENlnwAw6kZpWEIAwj
Oip1DQIg80gta94m3/XdLr3NzmVieo6GNyuMCuzLNilwkp/o82mxVq9c/DwSL4xV
HQWQ2/2jJgSIl4NQgeWtW/lAubnazql5/COYWHdS4ZqBYZCrF4jvAEhREc5ykord
h1jX4tCVmXztigjaeditUGYbLYoX4jU+ilN8bwp9Hm36UliHRTp0tblk6ekDCdZm
yWcejLE1HJAb4Tv1EXykRwSZzwgthf5jdiYE4aYs6Xct6TRC1XhgIFPn+y7/x76s
WbSiTo9/8QcSJNuuLLI2ohMfb3T7lZQL+tZGwZ571NUFgLss4WZaly9lQGQ+yVy2
ukh5qbAxXlxX3X6Q6pjBsml+FRhq5a+YC9PyBViM8tZFvHUx4NX+YjvyHPYNYdSu
Heg9PdRcFHz7qHmMXFdmdKENSFd2UQI9zBkrVzr3VO5RyOSeVci8Yn5Vw2R0aL5S
gpq193xM/Wy2Tjlrtcch9fBPuCR+FvpTN6JGltkuaEBVoDSL+wf6hN3c2QNcirwU
A07r14Zhl4KiXej7fqfO9IcGOHhkBTIYgyMiW0L0sHHe/bI0Qep8CjFbbT7voAPu
lrRidPb5KXivf4jhrRz4fTm7cwSkLjiyQhxuQRp6S20rq2A+83ksE+oZ8pjqcHvP
BiVJO/nrXbhuS2w9lj92rB2wyGY1hw0bbdt7qcDhA2TCy7h1r1wMbW4Tl1JMJX9T
3heNmaD6nZWRqkjZ6xdV/Yi64E1E7QpELYPb+5tTFJpuG52wZrAjIn49C7cjbLAK
kDiDxV3l3EOSy72B5YopvbMTxZo0hvNeWjU3fPew3kd9hn0czlB+fPIrklpH58QQ
wMEYFfMVwYummhFHEv2GZNCngv9AV+StoXoWiFOamIC/Bqa/TN2tZfN55U0AdNQj
N031twixPx4bMv3WxK2/xm2nzn1EYr3bUh9KMiUps2/S0cnYFW2u+UdI6jKUDviA
/sodxc2menm9rvy5A9tkEbU83gJmDlEEqFbZAMkgjZ2vLRruoWL8jGTW6LjbQ7qW
EI3NpNT4KUrO9o6+ldkIu7ERqVdPKlgh8PNEYpL18p4xBREbSZzhGAFlpnDWu6D8
5PgSw4gC1FlGl3jroEfKPhvgsT/ew5upLiAeHr11wTZ2at52OYaqA+5WihHLz7j8
TjAqJSixqebwLVAr36EHIoENFxl+xT9yADlGVEKtfqLUbUb1PfmLmUkvxgL9IO8S
ct5LXoBeR3kHezRdpPrK/ahTWdvjfGZG0DOk8oQGzj3aQXta8sjU6AcSNn0NCLt8
Whgupce2AjxUc76Tg4g+GzbS14vxnNCDh63rU7b4t+oNDlFf8F5xZJvr2E3YJYn2
Fh+XyqfSM2AdbALqDm/bsJ51BYsUXI40UBAKRuGH0SaiutlaTepMSYyNe81bj6AU
txRxemXZBH6CqkHafuB6QR3g3r18/EwPRTiHFP9H4+pqBYMf6HOfujDELIbZoiGp
O+Eu8wK1rlyIBrkuGC9d0bXJdW+vQq4QCvgCcKeBxDlqDS4DZhNZaIORNW9eWrGF
1oAjcZy3cW5OowRp0y4CWgjxkp39lhpxUZicUmRDMqgDhHPm6pit/pQtXdZJMXYL
t1m8deWc/J3u0/yR6VqZ7ci6CnutaDV/74txqy0HWsrXNsahrptpJKeofLLrrFbr
tCGS08pDRNnhclxaauYTTGWlWrfZFaWNJ3fnqU2lzeLDChSvXGUbbbkvbd4+iFXB
X2tMPMeJYbrrkQNNZm5umSPAh4spZYoGaSHzL1Xtwvz/U9pKoE0QgBcGpLYIZrHt
l6qD/5t715DzjX1hCkjec2cfiaermPRBs04T+wsH7JVdexcwpb2UqDvW/jFc3Hy+
Y2HzvHmpD1KiuUWHUWuRReVETJTFmOpIQmKFFcZ2GeD6TgjRurGlDToTcbU+0Hne
MqpzmKLFzN5rnHleaSuuURhymXAMkh/Bun5BvaBI1hQvu3v8EmWGpd3+aKv3cjqc
v71iLIXLsRwOF3sc10hv1qhOLWKMffhwWOSJ9L9JEggkXKABu3L1tlDnyWeAiBX0
xxodAYpRyJSDTW2QRxq8qX5gxVX2MboubxJNF1d7QnW78v08ZXLmBVH5IS0faTtv
dAm2AsGqoVMoBOH3aeZKonZG8FclgcQTr4i7F9Yql+NfEUIS/1Yj7nPPAGxoaaBY
PJ6n6CKD+c1KCZprQM1UmHwguaTrqn6squ3bRuFx+abN9LRk/JCJm2+y8vwEh6cs
q2kv3jm2phwXWc4tI9tkeIAnQTTex4lhIIG8LbmhXuaSoDd2/ZDVTC2Zouw+P+4d
A/XadtfN3BoUHw9ASm8NjZ5iX9Ql5HGGBQPAtlSf7cr0I7gQvpC63LCKWzT3mJkb
Nw2BVQdIMFxn17bVpYxRgzqY8s6N73tr1CfCptidqNIi0atmpSSlP9ZkUdJUCwbJ
YMMm3jsYI34IKTdBcneYlofS6bCew5BKGY6wJRFeFCYTgP4YUxUtORmR/qnbXUml
zbpwlVixAwKIFewjw5+NsDDmC5BW0IBVhCNIt8GfHE6fcSf8zCgmBadqb6UGWFzq
WFMBrViVQJXjttg2qqsOEWk1A15XHum8uOBCwLvSO+1T0YC5CwqS36vJoOB5Sgjj
CTR2MTZN7tOL0pbbLGsGByEZnA87kYqRkMZJHW60H6omW8KAOtRlR6pjVI1lhwb3
NrGtADWcbbwDLzGaxp3fQN3sjwlCEBQ9jn+d+zh9gjatR31IvAfj/b//RRzWEvNV
jKY3hjQAkE7r5Oajiu4VOsL7hOLq7V3MPuIjn0E+EafRWeHM8Q9GuWZW1GE2boSM
9uFLWS106ighy+8wJcQ5s802UcDWZ0XHVcMo/D169+LHvCNoe2T/EXiwXrvNT7PT
lQdB38CN9dxPFCDaWQ0J65OohdB8vp8GpdN/u2Mq5yrET3PQ7BtAsmdWoQeH2eQB
Uat+xJVBgmpnWEg4wm15128kJXUKkC++tCpH636R93Dqv+zPJ36ZbA/IOcE7W1kD
U/bOSRZodgoeRaREf0wmT9BXr4U8A7FaKop3ptofnX6ruQjTRi17wFNsJV0ZL4e6
94EfsCdq3rq5SnOtFq6DFPVrEhCLpGwwye/CgXPL/Aq3mhMZr/wZbKAXfefkZDLo
X/g56rVVtbhTA4wKE3GpqLhxjCnIz0R4VjgXu5wHWZLmpWpAavmpYezuvxcRhQ8l
Vnc2Y8RzD0ZAHWWMVti2kZdnLxNgZIqN19XXe+QLNM7ZSDICMTG/MslYt0NezA1l
3ZRP3vxLYOSZdoCC2eUmfUrba++c7I3fR4/zeH3TfUjSe9rRZ1EyGY4JWsCjO13T
twq8qc9fdq4j7hS8z/LUKjO+lQGa78WUr6z+m6V/VG/tbkpaols1LC8BO3SWIv6B
+p3ABZGNRXwUjKdQIF+yY9adrWPgpFbKaRowDwpyerQcOfUJJ+ZTohnS15sTLRfZ
Oftup4pNgend0jhJE1J/DbrAymwB1DzYeUoxjQoCHy5DH2ZiVWxM9M8BlS8xbfsl
xBji/silxiaZA0tU5zrPoy4sA5MAvD04F126rzF3y8NhxbMP6Zt72etIL1sEouLR
g5RUIeJ92B28GyUL1rdmFG/Bxbl318QLyJ7YWH4dOQzNqBgP6aqDZxP1nZv1GWJ7
E0iKKsDiv0cwq1Z53fGLXo6Xg1rphAcMHqiRKv5Hvmd8MjXqCVAzVLnfu8PxUc13
Eys+ZxMbJUi7XmeTDw9oJW88BtfkgClvEBnlbNSc5tJEmDgWt69IKtKSn7zmNRNA
Yr0+JRbj//DSSyVFFuWo2FivwhPXzv8MYPgi320TSjmgf2Yv0zTalcPiwaGD3iAu
2QNecCePgHziec+Cxbc0fHd3VU2vYhTZtXxqbeNLDZ5sdvWm1kIwpZaqRnUxtnY0
498Oi++ijta7I64zslBlrAAEDCdJNcVqIXSm5LtaVzvY5IQZZXnyPEogMBfm2zFc
W9Jz2Sn0RPp3TTygeHXq4Pmis0g6AwBZ5U6QeMPWlnLF3J6enEzm4Q2plm0oc++2
74OFt5ZKCIwgrbuAG7cuIyFJ38JYVoz/GqUHFGnDD8Skz2q4r+xdMxlkefal4/Pd
2cthrAIxkA1QOABeUycLULzCbvYZhADPcNaepAN0Cp1fsgcTTYE4AzibWa9LNyV4
R/YUst1dFS16W7tGCoAVqJf0AXyuFuMaE4VOxq/xq9Ap9dihn9Jz3cRuej5WMfhJ
oZancpxB7Cx9NNpS4qd2q+3/fLEmQfS7v0coR6e+bXj/FovY22ES5+UfrcQ5Zavr
K44AePwGCL8L8JL5ZvDnTJXbK+HY6QegiRnPDvN6wx1NiO0Z18WT6Qyp50RPxddh
+3YgYtILC2Z28IwCgyEX/sTwGeLZN9+f2Ps1V5i/JdAe48McJJu57Re9vfe9OZcr
kxhlkh8jcAUxTy7wbsTasdlMXmBV/3A4jlt22Mwm/yIV5TwQAMdNXEx3ldKKv8fx
gsxzLTAOzjNjjaPY3toC9HMF/MN2MUgeniZcDv1liIXhAFuj5rloHMKSfw2JUG+G
IjlgYVgP+FiA9zlJ8D2I9BFOwciYcNr1osN3ms2fEhOMTjJITTQVSbe8MMApNxVc
yZTW7jcLso0g3CXiimU/UyG81v/p7CG1Kuq+9bNsle2/YPS9PoZiDzFUBc1/qgtO
89Fg9Xd2BARlfEegIwJRpRHn4GgSlVBSxjYm94FVQGnsGEnfC9Q+VnwisQQaHwGP
HY6p91gSQUfePkyAXCZvNf9MGC9mPYNTfrflKncgcC+G4bdnwsThoIfABMzQrD4g
ljPb6jZIYYkaRLEk8GVgF1v7xAdFAgPYZAJF4+D6DBI0Qjc5mcKSZNO4KISeG3aM
RasdrQY11M5xGd50pS5qILxWbLI/YTUEUi8m7MDAb/qyevfW6ABK+6ZPN2lwbQva
eBE8m2LVTqc38Os9FmDcU2w4yMsq9Is+NknmYtUhtzYG/buZgrpic+t7jzS3ml7F
xQsIaM4Pt/TE/fcLxuF6keDAujNip+aplXqH/hDCIjW2d6fMo7mFUODJHGSOJjIV
k3d1lFdHWeDE30xlOH5jHGRlfIpdqENDUEc/mX9ODRC0MGb/xTiWyBDChz+/bSEP
SsERg6OtLMLeqB6HPXmVrmOGHHkUIj1PvoiPGRNkbzh6qitTOBP1xuyGkS6+fySx
P78iKUF0COv16HcN3GrilNiBMS7adbEUbyMZKSuVrZ76nYLLP0UcHslkA+xm3scL
FQfLOSDj925UsAvulTTEnbJsiBzmUnNbqWJ5L4JBKgjNF6SXj85WhD0E5NvVpx+4
UsxJPucVftq9nzrOx+T4XBeTHqRJ1ejSmbviIW8wa/bnP80ALyojqoEp41K8NpG6
LW4+I5KPKIsZrg0zApmoaXZrrGs7Oh8qkBsO8IvnfI8jLImCGikvykMHu3BmJnh8
UdlPICbCx3+9gdwKGsGqQPp1fTO4wA2Ea4ensRaqFMJZXL/y4a09GFSeqGuMWSCm
SY1MsKmbwcOa6RDk6TOLq4cBwKCqDtV+taYT2/xCO+hTF4LQXApKFWVnJnCESDks
JEtPUcuABfRUwbQbo5YWBTnTEAql5Jkds0ELprZzBs6+5olqsUApqqm1q6kQ6Tw0
97xPw2OsWeOhzcTASRf7nT+u7mqtZxJh5uSC/fj2hLyFvV4Udiu/U7+FXss2jUn5
Lb9IZ51rLVtf2dmwTmeb1fHjLHIDzHaEm7EaMazZ5IClaiceOlQ3py2wBhJdJYtw
jnC6EmyKIsDU4q9u1bS93+XYl7TOn/+7uYGKmNa3k6D5mKiFplD9nrErjZHmcsF9
DzWaixjkiY/Hk561U9pxvA58ASFIYew/KD/0Yyq+r3pj2ilRXmbmbxKEx0K8BoLR
7TgTIuzMm4FGpS3lFO8fQE7ezcNI06+TfZ8BSiARpYE3/+DLrI5BVocRQ33ebitl
wm8JD3Z9PlL2nyJ1TFD6E9MxgphUYJlA++2KF3hJWs3ieMzbNG6VbLCzIkuRYMoY
tVz2HJiGQ6JCy7dCmYhYCaV/i3sumTBn/Ja4vi87B6bBM5bmoefwt92kvTBh5KNi
+8iAAPDw3i+awTch9ES5ZtxPVy+Ym3XbSqxSjf9MJ0lkfSjNVND4hs35g/6HZtG4
J4SowT/zX9WoubY4BKGSUdzt6e4B0l98aTgA/8VEEiId95AoIEuWV9u3e0LbIPT2
nzSIq/nZJaNPNhowIKL7MW2q1DJSutOYfgr1o3JsSikjHPuhwdWnjm57hMJZR45h
lZegzRSnxnwkZGG7KmfSyjWCLQiXF+BXAihTYEn0pi24bQBAZkr4tw3vS1fDYFPq
b48nnz1L3ELG8nfJCEprWR7VD98Y4XhEkGNwYNdbNkwMEAA7wvQf/d6siiBE5K2L
5Ky9FaMXQr/V6QAmHyGGXLXCtVEDYYVmiq/NgM9rSO0Rr+7FAD5PV2bPCNOBJ8cW
7AurZqZDoUfqZ6LWUtZTHzHDEGB/ACpwlaaF8q5GdsYpaHycNtmPAhhNf+84ma5m
uXjy2Hu8mBAUcrv1l/6ewaOtGmU7KoPw+U7OfvJcCLGvdX5GJZd7djOnz8UHy50i
55ZqgMsFqStVCcpu6hsGahpqbnKBx8S5dhMu1xyUqy9/IGFaNzIXRzfsH0NXsf1T
U5YRaBhrC57lLRxHx8mlaN6wVdazgFo8bIOoLQk0acTheR0DrMsQHMrBbaPrKlzj
0npH61//nuHKyKFeP3xM4KKfYr0kCCpSlo/PKvzm51AiW/7usTr92X9d7KD37UGW
g8j7HvV+mrR9ivBTVsR34hioQQvofFWQ7eVhViHDghoymtvJaDIV8Yrjo80jrDzw
ad2lD7gPWGrHr8rUF8nirY/40VsFmMx8/kCwoqnKhD4OKtfUJYw1YDzRXEAJbdrK
Fwx8opJZY1Ss+PnQMnU8VPlZPPauWJ1odn9XbuLBbO91YgBu8XJnfeeo//9FwkZh
RITr9jsMyDOiERo8jg5r/vDQCvc+1a+DYVL6hEm/IdGFZG3tPvhuwBGB9ANPR2BD
ca49CKd+JLcp40+0zuKkQoZQJOoSzN5gYxz2FA9eMvmeezrzFkBr9xkROW/yHK1X
0h1+Zxwytq+5z4/5s/TbEIR2SnVQfJLd3Z7iB8Izy40Oi4R4X5rNyNV0mXFaCOVP
CZL5Xlio47K4GXTWRAtvlYSOA4OjZQZ8E86JGczem213Wqzt+SKwNlLYUjb1T6DT
07CLA8NPSzIrgQbAU51sZJ0JnR6tGlKE49FaFJwyCYiIXKo4tNVJAmJ+5az6N5ar
ZpQA04fO8oByPweIDf2vZkNC/V8qRylR9yuWv2Kchv4GusrflKwYgVsWdBSYVfAt
rZOYH0r0t75ulXsi6ms1ewfWI0G4QE1wcW2oECb6kEQ2ZHMkB+stDkjARvWc906s
w+IJhF9kJmnMxW3d7jOaKS9czHw2o4Y1MjBmLyzTNTL6wOmfvptMBg/Xr6au42t8
+jGPeqyugnDb1OpJYFg8dm6Jt0TGlFyWzXNS4gcgvZ6Hr/IX0oya5OaStO8Eb+ql
BpVQrtsTk0iVNJQ3irUezWOgfLvzAaacJzC1ldDox4hD7oamNQrA3JrqT+dHfLwA
0IxIve3v8SMMqD6r7/9jEdrB2pC4mGLQtRHdWbmX0QONP5Kp4zGamFaiFiB/u3tp
iB1LMC+Dl/zezm6Baq0mvMv/SEoS4cCZCdfGpzDN8lEbk6Z/GgPtnUofjUmaEt4e
enPxyDVhrb+Qo0oTgfgv19nBf5k01hRH2GDQd8sbHANV8Mxc8NzApix3SJkllZbq
cU33YNBtViIb0julU1LwMUvFVjuBGw7ZbdAY6SCmII1o2F7uMJ4jztRGIZcPJYnA
iH0uN5m01bcgvQmg6A+k4O/NeGoIhT5c+nuSwyigyhe9FE5eQ6imoRhehHE1TWz2
TBNB5nYcYT45wfjbPX15QANyoC1Reciv3xVwXbWCxqA76pbXMa7xVC/Gfhdn60V+
qHazxWZ4ZLGlWT+AYoCpbRIrPbGpTH+P4yIcwLFZcTWPpyxDvttEYyCkmUDWWGyM
NpWpfac9G5Eoiecf37hwSEnpSCuovtmA9d7EdQ3hjg/RJCWh0+7gDfIbSScX+GIC
whKapuSGIYc77bkFMOpGNF64jxwy8h9zYLMgJ+uawJYLg4GORY26hW3q7zo+525m
IGb1Zz7oxTDmp8hP4xeBps1r2Tj/Ig8KlQBydsvOebGiGFvtCs551gvG9SzqmmxA
MuY+qGa3t6LD/Rn5H5mb9fMVDJlWz5oAH8z6rNcY18M2b6gseWDRVGIGlXGDc4PJ
p3/IAZ9E4tevA6KlQBu7l5ocy/tfKMmgKxgHSiFISJP7RZEXIj70CTKjoWrtMbWd
5JhUAELLBQtAzNKiRUUPNpZvWpORSRLxfEcvtikkAjyyeVK48lbZZlhkcsxwt5V8
uYPwoprV6DK1L5MQaUZOfQRHgzVeAY9VPKx5QWu7Hjula0NG0qN62TaSZ9edc6BV
eWi0E69fwFqKzlUfDDM6khWxMUXmTYrTUm2mKLWayiU1ZfiPXvl8lDjdt/0zy75o
CtMC46QCEmdzT+zNZ0JUb52Rfb4sg/78X0Aw+3o8Ttw3zfUTLHI8omzFF18ysqx9
Q8w83MTq/63HGG0XWZD8CBVkWm3Rz+jkWRsWX/zmTCzZGDEXoXMCqirICzNQMrzf
8V7w6V4/7S4mAlMTI0mZr0yZiIOl3qiCtm7eeklicPKPTeEobHE/QGUIGkTrpq6u
CC54uEceLPyHBfxWwV4TU6DcG2AIn4L9PZj5w8ATYk0emOwbf22vqCYowoeGqdau
mtkw8Zv7eaSYc8tnGo2xFgf94mY8fiI/+vrnZmPY+MkXJmt4cJTJowXlpIN29eEz
WYVd5Kt8gSiDV4g2MrAXzpBnKrTJI4W2UGGx5tyDgoItu7j1prVlWiSIieZpoac1
g/CopNnBd69CgTBYhlVBQCdimW3pqn2i969WK0xZPFcX2PVu7zz3mvshJWVKUt+w
BmHtIVfL6gZmKr+D3FXKpq+yCqf9EVam7uLHiraKcv4JO97y40xAl65Vq50ApTtH
0+339Y+rBTe9NH1o1tAdDqk5Z/qMcCCoTdr9K5Iyofd11ns7B1rkE+O/VRuY2fa4
6VlY0w1R4sepSS0zcx8eqBBp8X85NDgwNQGatDaCj1Mkx4mFit7kI4JMD+Ahe86+
8Va/TWIkr5+QV0PL7fx3GsB9097BgJQ+KS/uMYRJOPVJPyOJxPT5/2KGB+rzEf2c
Wxt0pJ1i/HB5IpYGp11l12f3nD4t7dS8GahlRDeb3xuS6E/mWNt0xfAJJf5ylpJR
KcglAXmaNNNzYektPRIFiMsC7KalpZgBop6mO6wm4ncWmjKjFwiiniw7PITkt4/d
qyyWVlYFaWkDiyAzNMBP+KdnLhOeqSqUHtGRnEoTv/mKpD8dEJ6yTByRFZoUKmTy
xqUGRrxhvdkHsNsHD7GgGrwQ0sxlO7tuHowCbQL/cY8JsokfvjNLqLEztCkV5VX3
BmNpybzoiE6k+Esk/vGMhDsCcrG1forFwD2gv9mKd94DdWTdqaRl3TAsapfhMHga
0dbs1zlNnkCtREYl8EcF8d7NMnhVwIvoqZBsb9Z/52JzIq3n39hBRg4xD4iex7jq
ILbO4h8sieh5jc7hv8DAnZLL8xdcwiF7q9YE/alBiMI20cFDm9XYla4BB5rp9ah0
qp3ylcO4hGvWSLjH76Y1SQlju4UGEasOSJniCdKWA70GGL+mJ2rsjcMA4WaNOQK2
eOLzRehfgdHWMr/0JIuzbsI78y70EZvXamcDJWKusX7gvi5zAE+PrmLlPVBWC2Uf
3bHi/JlNDu0xvyIC13qQPg+jeZrqb2MoLoKk+WFHdvu+IPNLh9hRzYSBBjQ5hgY1
cOpXzKRqb6iCFm17f6MNFdsVUX7BklcDZeC69bOELtXf1ZzmQu9g1+iiQxYLMbnj
UzoL61J6eWBAyNeuzYCvGabuHDqwsCF9vJqG2q4nM6tf/amoKJJ70/+PCUlh12R2
0KgXSoLuMGOiSYKKi3OyjDEi59ERm3ffmYgM3BuWwGhAOigP2xoefdc2sbfq5lwX
PemfMW7VP22QNPidJN428tO2ntP9JvKkirbe8vu3ZkoO26FTkYhopa3gxeAasPUS
2yqwcm8DDaYNMNKFMZi9Nb+Jb/+tRVZ42YqT3apIZiBAG8oCwiI5rBryHpU3GGto
EFynbHYb5VcQYHzO/0MBMJHFHtUVgpCa9IMA9p9UACUj6SaeYunB+jpuS/cHrcCa
3ZErnEsFKawc8uSDJYqAvvL128aeXAV8wuSkIISrIXwvDrp9+reN7y+KFB2VgKOo
H9A6wO+T9t9c5NFEK7LkA15xagTMCNVPRG5vjOmRDkO50Y9ZWpDOK292zLviyD85
u0xKMn1HCn6qhOTuRiKajTkQEyJXxI6Oc8rmwC5ZCBucjNLKSgo3wLsEpsM0rVvS
SfgGblNhUr2ETOEx60JfG1V68aySpJl2VVBpIsuAvIpW3xaN4ZIBbBGfodx/JGmi
iKLJ5VwLgbYiMdQLwizYPKYcAKuoDbQbuxY+Rb+93T0RSByZbtReZLhh0dCx8Gpa
eU5jBBiCAFALfHDJBVk9gt77ZC36QTVXRKtCfoQuoz2bUrxMcPftMpZLmUeW730q
zSLkS+fcxNcB6IXncjg8eVPfoP01OomVPw6WNXI+huqX297MogG9/SQrJoY4idfM
O+9M7aBpm4iNZnu8fqA/ZbfvwpS9HMsGTlIRUk6j1Hrox3QyQYDUSCkCic9s5UYm
3uT5iaGYJr7/j9S6prHoEPaMwgnwXxf3GccuI0ZDkt/KE09ZxtGygjqT2tYcipPA
XzWVQGO56lrQexMCo1GRO3lBvaVrB4SBYwxCHJDrvnGR6LmWIyUDhEAmmUoj+EtK
mBZSdc3TDqCGHThW+lagZciDN+eif6HRnhlqd59HhdbNKsckTk0tu0q1boP/AmoF
wFc3DS5IthFz0zu2Lb5e1A9nqCjyT0fyBHfmL5LzdLMSExi0Vq6mL3Aet44DBBW9
z0Us2rYw3Aw8LT5A40qJ1WjUODsiijZx3Io295xH1HzJjr5ItPTsaIUGQQzFCkf8
OVfafQ2ffGuik4QrJOQVZ9YQK9fxqNlK05li06sUFa7vN7srRytR2LKGeRRixrd6
kUVJEw/PQxH5u67iZI1HppDrpn9Rqn59HvXu+3UZGGNuHxFzUfEypB8lx7yl4trI
xt5Mhi6sGcqHkFvInOUEw8uJSo8fX4+t9Q55sxTj+wfpMJNbPzWTvstHwD6PzZqR
yesjGarH1WJDbkg1OswU7ymz3LBkrxvXN13QnA/tgCFCAi6HzuMe9TEIpcb2OvyN
7jbVOJw3ZRU8TrZQ3jO1ye274wFkcdl1Z+ckBDaPzXyrDI2od7UPf/bdCBLHHwOg
c0H0qbK8E3sviMBmL7+iwoEL4HS755rsP1O2/nxHMIMvPtz/rzA3ieZdCOSso9BO
zBI2ju5rCPwFydLQlrbAzdthtt5SG2InwEPULBbREjcphrZ/GsApjMPB6FdRKUPI
fycyPt5gccuf2NGCpDOg8TeJEi+Y46xtd1Nc5Ts2CEVONFgWmYy4cy8mxljtmhzL
cpQwpLnVWud8SgMIdXycb1MHKK6VZE/hGGmABxdKQfDlKuWmV8Tj4mM0FtJL3i4V
Tpu2Qmg3FvOHVLs4R/JCZzhF+B5AuTjXzWnuHJq3GnbubJJZJVrsCpT5rVnrQjNp
Ip/ul9uE3cLqI5V5ej9yTqgFljHOBiAetgNEoAUb9xIwF+soZ1IoqgOqOy54TwNF
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
f90GsNR5mPHQoHNT55khyEt0NiyRFiRRMlrc8aywK334ChWhGf/93anDnUH2dyWr
nUKSPzp/i7AwarfUIIRGlS5Nt2JjDb++ktMXTrYKg0bxexHaokS/GuQynM58eXc0
Tqmz1gBkDIGIZGamWLd05g0UsWHsXU4AGa7TSYguApHWmm+8zC4/SMP3ixV79oW3
r4eMZrmrqJ2GrebDWYNqZQ24FpvC+20y0w625RKSrbgJjgagv34cNJv7DPiDV7wN
uLZHE6u7RHEUdaTnth0VRy7pxsg0BKGGoducGu6eENhWvlD4CeWa517lUUTYjpA8
iJXkP9/1JOHyAbIBenlZJA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 21648 )
`pragma protect data_block
lDeVruBaPUgBU0I5XUAboPGFkuXZAPhKQWlGu+cuNRbql8rJnlxR5o/HMMOwuQ/K
LMUAUg40PSI+rviEj36NFrOVwJ0IZ4HMvsJKkL5hdEzONaiJWPRxYrQIClmawljk
uuQHq52A4L03sAIuc6PhBG7KFdYYTpHWWMB3Gij+6PFcXsBfuBYsJtQ1GHetQH5U
EYlNyV+NQ6K5+Zhpwo269jr/wShk9dKjbz2hu4pj1QrFziXqkWquKmcljPJo9g8C
kcX4Ga8VhWyapY4KWcnDxtFuZKrfBeh4B+0s/b+2yQVnZyb4SymqukK7kd8SoWSU
RFsVRxKfGaR2fXJGOsZR4C4hp1F4imSDrb4dVprknogwRP3JX4zMMwUfIBP3ebou
aV2XLr4b11OHcRNFiYWlzeZtaG7cahRA+u3kMooepSxB2T0Nsq3gXnkoTNXLjSWU
X12eoh6ovaoavoGyBh1j7JMxhSMjboiAMpUiC1us3UnBcGxXn8ZppFAma2nayGZQ
36PIwv0g7fEyStqNkuT2XNSi5mTwrUVvjU+nKIZtCRW65F2O8T88zWDiYqSya8Le
WkRTzHi3cD61qOZXIwQ90khEs6xeyS4K9Zt65jhmjW+SVAM/+gHoXT3VN9c1Iy7e
22RVxRcncdScnje53szkL0NZX+SIDxMkCnPfkGbEsDR1oIzGAAijQjOcS4Cdrzxv
aJ+4P4uiWl/SUuibkXYXqf+eSamkkhl3nOCCFDDaEOW4LglB9IEOnkK7OGHglILD
pU3XM9jRAAbKxmlsVjPQcxcigWgIgb49fr82VSVjZ1fudABzN7ejTgD/BRp//3dM
4b2nuYsUxa8ohNq2mNmXDAnAhyH4Jd62N9cU6G2KXGScVehaDyLDZRtsVWyqsAxq
O5RdazT6/FzerPLV7PIabxYCP0MYwwTPrxbFOJ3Ohe+f0pY2cewpIC2soPHPOhsp
e7AECmkI2enxxlEm96znMR8+Sgyh3RgMFkTuiqaphz6xUlUrursoNLzEILosTnVG
zbH2ev4OEoHw2TV43CXa27hvBnEahVv6cRV8zN/WJUaEErzeU77ch/1r+//dkR2E
YA5l4uB3Shmz12w4HsAAwdMAIkzpmdP42Ad5+lAd3fLjTF1gy20woNCD+SLZkwsk
hRGPeFYB4jNQud481TbhHXL4jLmz6NQiedk8h2fBrvoxhuzuxJpGel7QZMZpvQUr
9ua55eP1fpyjA7e1q/1NTNOUSC5kgSzCGPXs0UFGyk40MKp2g+ryGqPqUflccE2/
MVIh6gJ+UnqlgQXEDx6+4xxF9ob5OPe6AJxarPfyhvCejfErlVsnPffyu9mPWok9
RBmutKgznK7QkuAvl9agIPS7GZuV1IqlhiqPKD4ekcCOA0jiteP5TVBP2TePx49I
Hnok4xpclIDPHiViN1rWtn+VZZQHU4IPMtT/fcXnjBH8eh6EuFsCe3ypEwCp2d3g
OvXslM45KsVlgm/M6xbZNJMYJLTShpVSiVzxzWhv/qB2AuRiya33jkI1HaeLE10z
HLhZfNbzItKy43qQxLml/E6iCJvPtywZ0Yhz+EZQlHz923+488KhBDMviR0vGwOo
5NVp3NY1/eCH3TSEvRI9SJn0TpO6bZPWw/3OgDDU1IATF0wi7nRy333//88wlcp4
6ybaomhYyVLUtA9XS97BbTkii5OaasYtM+k3P38tKSIt1QlmIkznNKwXIWOdar2F
gvwRuEfd0ZtNHzbKXUSBwaKqv6RlUaESGmKaKDFkq3h5eMb0wl5zOtM8xqyCFIZs
tnVwtwkWY5h8Biz3fU9esWngbR8/klaQY71osKF5F4OSydEu6/j8KwYJdcbO+3f5
hrypZXVOQ0b+Q7avXrqeB1UzmmI0YmhbZBDXy25nzOQSOsvcqj38UuBna1vOGP39
ifa5iXC4cKDH7RodHb/HIXQkd51zN9ewuw5eVOgpl2yxeCvzo5g2EFwbn2qss/F8
yZwHzXsL/+ExdfBkXRYhk5xppegM9EslzKrXAfKpctZu/IkXDmPOPycrxl22VAp/
+8F2FpK93xBskavsJpK5FHOwj9mZ+c5Zf0eOS/q4DAe4GY+fD1Eb8nQe1XHSiUjU
nRE+lgKYBnCPcNAXfq+aEhZ0H8iOrOtBiaROCsQn5AlRPMel79nBLdhYRSm/ev4X
L+nylK1JlLFU6ADyKRr2J6wz3D8htY6VJGNihLz5SrQlofK3bbY0LvnUVXd9LMuO
hXV3IOQUxVGpVVXkYX1mTpfl7ROxVSHeVFcX9Kvks+VggJ/eb896AOla5AuGHII1
u03uBDfTzQQVNdf53WZ6kqbH6kiSe9sLLEHUkWAJe6hIFkVrBAPK101QwhV2ltYx
ewUSHIDgI2vCF1W+Axs2KhVrDxwnQkkLIt4+7K/ldo6KwgDQlNUSVIyY7sTMa/p+
SzEkLQp5/BRcwjBRotTwt99p+GWSnXiXzDWtfx4oJC8rdqRhaYYY8o2ug/1r7gmE
En07V7mtZgQvLw9Z003H6hybSIEwe+X0Yb/X+utuOK0YITrV4X1NKQBWUs4OhkUe
irvKSwEJu/25U40Qt42mjUZBU7fHnImdcCscT7bfj5avs0iO5zVd1EuqXJSwX5yh
tmP0+xLsWTe4LtGgnx3PusOWE/s4NGMLG1QTc0nyxvKRPlHd94iKz9fCG0/VEXS6
M/u0pW3vvf9bXvNJJ0NnaX6c7VtCvEoVke+KlPsakQaGeu6ce94q1N0VKkUKMDKv
VqyY/TdJrZ+h1u0WSVGT5/wWKnwJHRNXdqt47+4w9TmUao7k5O6UHvwV1VPw1QsO
MpeSuvE83HXd5+3e5qZaEJWgNCJTA584ZFsBxDl4KfLaG7nO9rZBAtB8u/5RBu98
WU+HxbxCBXzvPsTqdMt22eguprGgU4adFTGwDqCY9cvVAyoM30A1rMTJhUJBO5cT
QtDh/5YXtsN6pgd3/h1zie7kCB7iXlrwLYkue32xFAtTy+/ByNnsq1P3NtiAdMb8
8tlcdrFYgZ+sRienwwbYS9Qv15UiUUU3qCIOrs8VrqDxAW7/783bk8LNNa6V9s9i
I4bZO+V+0m7ehcZJ9ov3DOo1sICgEg/AE6zVwDtzEOrBjP5Jvr6sdyxaMx0Gg5rr
DmMTtGOkQLgf6Eti5GrCVOfLiITDIY8SPSs749rNTt5dbZh8rcIcrf+7fSWGzYUV
KAojD1gpGQycIrKMr6BodrdzkPsI6F0pnQUS4KwdLcTV99bnE7EvoDQNaiQGUqfq
W/qmL8N0kSd5/BlUQ+tfw92rLEE5diUuHCugLJkvS1b0PjRhaB1nBVT2Fudnw0Jr
Ip14u3reY039nW95BvCwctQ97oZ1t/aI60leGaqqT2Oi87D/V9j0RdZhnWs+S3a8
cADq5Ezktz10SldUtpk1K/iTc419lBWtWC6kTxEJMXszlfvSXMj0+XD8BO0FtwvK
2zudr5Y40630zhl8gMnJAgWibc+qLdFC4RiOycJr2p4/nhla+2tb/UsRsIhWb89B
hFmYypIew7U3/4H5CIuIid/RlaUme7hYHAWUATNIuf6yxA09hUllHYFddLb6JhYU
eChpw4CZjFMKuK4aprYz9Ne7sFMVIvOk+qwCwyoo3lqzoxGcVlvhgeRRLZ7X/YvG
+qYJtBCrewVFEiWGh4OyPr0W0gos3j3OacYr1W2SEs5n7etGszEi3VwVzTil7zSh
rcUaLTNQWo6EQjUis8ToJwNZ1eGjauVOF2ZR+j64yq3V3kZbmyU28LMX94lcuett
BvcWUJEVqcpb3aNPtsS9v/Y2r4PwlvRmuZf1A/j1F9qLvExjEDNkBZb/Hgjk72nl
bun5MBk2bKHFjDMY9TCIwGZE/Q9zKA6IAOxnpOCzwkQR7LAJBeo+K7RyVPVRRGOh
b6l3YGke+T0Y0RtUV5brRFLUbdYVS+S5K4A5XXw0zlxmoFchp6ff/5SoIbtzQVaG
owrsmMc9NLTh4MLsB3L+zmz8636aHZuhZSQGDT5eNjc2xjhEZchEesTtZ6D9r5fV
t1CXaM5yIHI7J5TB/9xADyZXGwENZm8+y6MLnrgZ60QQ/oYROXn3gZPoehNJOll5
5qB4zhvzoIgFgye4O/NUwQ8bCtextanrTGRUj/e+3Dnnnl4EC9TZmMlftmroseZ3
25Heafgjq92Qdft6R1p+tveaYS0t1shPVrGY0btYPWro4uHuiOBe7Fh9Ryi9MQ6y
zF7R/cZxsqSsigcPYEyxFkNNLJPw77wX/xPL6LvPNxuC5pmPGPSgBtyBLn83n5s/
nGqgmsWNBnt6aGzyGW9FZcCYMI5ixagnIw7b8X1HbO1kA8Ooj1zSNhkTAX9zfXEe
kR6dO1ZFeWZCpuZEz6fpxKzJ6qKFrPYo4w1Q/c8aVoAklbBjcMxULnpkAmBbrl6o
EKFqSqJ4O+W/5bfTswySiCZdx34w5XCvRMsurJZpELc+mWTVundW4thoN8/GtSwk
JqOGmK6xEeDiLuomFzsNz5/jXJVXISPF0a6JVs/eTsicOKZO4btyHctREdv7Wf1C
eV40h0NoqkOAY5gIaHW2i4VulvgI3mwjHp4SK07GSv/isYPR6VQ50RnV2/4tPcgG
njg5+FsNcSeJcDlIYVfs/AO+3KWav8HQjjAHGmHF6yjzGQFjXyk02EG8tWePEn0V
Cr4VM3DNC009F2gmErzNwB3qtCmUBySzejHQnjhugpoWb6a7mVv7grS8gACRnknf
xTynGUM36Pm1kRQaDTYl20vER/yPZA04b6bKpxV2Tt8yXDMmDV4Av564Y7pIKPg1
q/9nvqTZjkgDdddFzuk0KgFkP+ZQ1iGY8wkhXGm/v9egjCIAQIp4rEt3gX76kN2q
wXD/0wyIQoAObO7WILqVwQSPUS0tVfbzQk8Ek7mp/hOMONihaG3KC4tDKdd0Ryt+
5E7QS6cqVBHrnSUubYS8TMf99dpiCKcvnGUYMqG9yHjBg7PT89bst21zqE0MTYDR
HeuN53dfGvbcTwrykxeYMJAn+wjPYvFAUI4cQ6MQhA8MWO2lSGMydyp+uW/BcAoG
PnQCie7DRngzYjULQNcPpKF/2kyyeoqdsWbXOhSMOwZWJFehOrj0sC1m/Odnbgdb
RAxDW9cFoncZRla9/+vBKYwXk2wWanSjflWYpMIzpFLvIPqVHhEeCtgjmCMoR3Is
B6HRvawF1QlBi/oYNTHOtmXvp1nXBErG3YKLCqB4TsbYyBNGqwver7dEU2cA6Kfv
tDYYsjMJECgEA8K2n4ZPioYYcZ3cPMMM8GHwR7aRHHOG4gX+ML8BFDKjkclUbq2v
tjIfXa5dgsWgEYSSIfR7bxlIG2EogbdRtHgJKj2zQ5A6ABrxEwJG9bpbskswJynM
v0/bmvVj+IrFpg4McUUjrrcI3zO5V6nXwLDb+ckwoCKEP2zkF0oWLI2XHbhGUu6g
rAEIl5WCc4EQ0UWezfBJvJZkaHFvAjLA2rPCF1cKhLnEWRftXaesK4HwDWzlCD6G
f5aGapeg4Bm6ZXIw/ChfzBp3OigFOOivvdUZVyeSBd2UZrzAcBy9TQc70N49Za+b
8Zi6ssp2mk13I2b+navB8drlTsnSZiQ1zz6q/FjsturC07fMR4k8UfEaTz8rOa2x
B+xGKn+85GzIeBhUSn/2WzQimw/g5TK3erbmkfMWIIYA84kfNWhNB6WQq8Iu8oYw
A1zBZIalCUYLAYpRvcam6/G6EpkoR4P3TKUzJ2OjtZX2EagSPIKnKjIUzDlyrKxQ
ZhCuqRHUMfH5SfKPvhBROjNCdf8WyUFjrchC8boOb8Xdw7AmvM6oyN4+ZTJDXQ/W
9ogoUM4GJ+9A+Z1qF+hk9pMkg9mj80aayZndlW/o3hS+yjjPFPkN/PBcKmpn7Q2m
EZjMJz1hlujqHIwBiPOZbbzDwsbQW96znoh4ARB9KTGDgTIUflcyOOOjDbGyV1cF
XNxFyLCQS1Nx+NnUR/QATpHep/AKHebccmtvPwF8Hjlcgx3hr0iFfRKU5b9NA9E2
9K5Tbr72IlwZGEPQf1LO2T568mDiIt/VtsdcdwJJC3DnOH1B4fpU0qDBACanPBBe
BILqtu6DbWWj4tn3DeFBx2kDqlVGPNwTngRNazFMQ177RsR8hbs22vCBRCWfhc2v
fgLdiPyScTgA9KhByULfS7uKk1dS4EJNELZSkpp2S52+pnClbvAolwG5ehCcb9VR
bloRtuia/pcwfg78DWoVhZrnwrLMsQrGSufXAiv5KtIEqD/U425BFRod+OV9fjE7
hACa4btcXG3Y/q2ySd+3w1Cci49R3zc0+ZcRVzNdOrnp7gBdAiksPElKSBS8fqSb
5Nyp9iTtraN7M0O6nGn68R458odZZ/tyotftgS3gfCflZKYcKCTkrtzMMOWwvx+a
AhOqcaIkcyLsVBh/s3pzLVTpmO//fULimYs5nIkUfKN/TlS/VN2nDKkvrv2LX0LG
su9z4SSlJe9j3D7ISAc12rNOnG60gAzsmb7CWF4ha6/V4s3dq2F9F/vpcUtxKAPX
GQWX241/hCQhbKZDEw1y3fGhJeYaS7I+flyooey2XFAF0FMFT+7oKUzSklNdjHcb
mgnyl3jlUSQqNISe5DOuXzbLCqfxVuffnpPr+qVFRWsPhBGW/zjJuK5giZgO2yuh
DMGI5F3EiJWwaWA/8SvEwzBK679Q9uX8jFCD871I1rhg7oiBDzvvRj3ndWUMZ2Hc
5BZhv02Wb66yMoPwisuvGdsMZxkzcgGApa9azpBdFXgiLS8Su/+gnk7aPlsmYeJc
hv+RNZFP4oJO/XoFVdhA4O66EX0RAmZkHyvKrgx9bgZpTjVxljwDf5PClDqmJEnQ
Yb0Hl1xzTTi2xHblcBeSpNSBplKLwAySRqtSlHOY7GWn628t/7ydhdmV9n/MYIVv
+XHx1w1dLNwKih/BM3HEKwH44ZYNUAuypZtcV9b48sDS4Jqt+RrDsJIK/4TSMDaH
nI54gp9LD2/5Tt3cwgQrhxGPylPY2S3pp/lVmA8wHjQBxpbTsUo/Q3pwf7xz2zW4
aQj7PAXaMGO/Dk35ELWykSP9gfe5mZMa/tzYp+HoxTXuujQm66lgZEk3VZGObrm6
EZVDwhoUgbVrTVpuh4Vf5AzoE35RWrAnjYfFnyffukaV11xVsx5iEBB2ayNzhzfp
YqTIRdu/hQnvf3jtzd7ZMQfsXneQHXIOp11R/S0FBJItn1Q6uanITeZkDm8Mg+M0
Mj9ecy3B6BriuBtbBeo37Y2kM3f8ofg//FZX0/1bUmCYubPoWPybEuIdBRdkDbOP
i5TnUOB8ypeFe6ggBUfRWaSCubQtkRZbAVpKsA9XH+PIJ67mtRU11A1otVNs9ue2
tkqCdoLrqy25xhk/bVtmXQrbWCTbbXLTesgrM3SyukPxGIQ6vR/St8w0buXtSvE2
PKZVKy2MQgr41fKoJya7e9LOX0//CdDvsytkaHVED1bTaCm19vsDJZM7MrO9i24Z
d0Z9ErwKd4/kMk+NyFG4GsMoYDGtZPSCz6HSauI6GlOOd7IxzZMCcN0I1dL8Tq+a
FEGsyHR5gNNfThKyKoKHTu9m5PxJM3iL9DSQCoyqHZFl2irDh69g0H43dLyGGj7e
xlTPg9HM6McT/NcRHbIIP2usGwFr3cMRvNjT70MPT3JUXsxN2YX0/bkGYv7e90uw
onOWmNHLbVxzFz6yFsMM9KJav9oavEJaLNlo+1wxW9kz3lxXSQb5zY1Xj4BZdauT
fUvswaevbXY/GDcOOGp6xQ8MStk+hqI6E8wThyyRLsX0tIGRRHX/EdVznxnChG5Q
sFG6jcSeda6+VV1QIHzaNaL+G5nENQSNJkuno4IUudx7vygBOidmXD8fZaMdW6dY
KgXs9DQn0fhCYqLfL9asde5WKm7RGTbQZ1pJyGkyUORzWVLqvYVZ+eohFS9uY164
II8p9gfHU5p/fxefSnhvIuSyLb3oqBKGvjzgwuD1Y77v2DkncCJg3Rt984MmoEuT
UZCuMrohuU7u55S5dzX17KNgVhZi9y0/IYEba6A8ljnPN1h1N0UP8b9dm4W/1wTP
LFQfv+GJJlgAE3ZT/t1A/QyjQdl9lejFzXn7EQFA1XVJxh1GF70KssBx/7lVRobI
JqT7iNNBHfS/S7sAN6RlPwp3hgPdemx8lDMsn7EXTDoC7hta4nbszEX3SBtvBZ5p
9WZCoXuVaBeT2Uox0ClI4ZfzaUVd80yZDFPEIa55sDtFBTbRzLXE9M+WhsfpmL67
c4b/SGzmo3cp0tMc4HN4tj0Q3gCxhi5mvRMLVFBL9hwlsCly0h/itv4sKAR5VDUN
plYKJHfYim+Ao2eLavaYjdZ7O/0PVZq/WZs6hpwn2FPrjfb2gvSMwwf68dqeU++/
E4QrHjgJSWuvx6iNgQrZpSvbomHjyzHSs2AKTclQwut7nm8eji9madK1kzY7Rmhg
dfz6upX51gjZchMfTgSAZqTBLX/CMWQug4g+c1BsysZqnqBJdTGX4zVibHvEYM4t
sqTdwqHpKAcs7FDkUjvO6P0E2dRD3Cvy9A3Oedh/jwfPLuWlk1GSU7l7uwcb5KKY
1B/mE0/WBYTK9TdWXcYmQdnoDF6Pjw6PbakmvNY86mG7lHGtm7h3SeAIPcyzR/+/
orGT1JOVjyQibHA8p2UBc4v+T/C62kYJXnJnNJW9UGaUqSSq2rPhB9V2tUaG0Gug
pGIY0innK4EtsqPLJoiRQDVX+v4qK2kN9U07VWKg7IiwPo0beAvcalkzXnFHCEZg
AiZeaxcMsonbaUYVuU4oZEeXXE3rb3iSeQhaoJ7pCRfgu1NXwNaRHnuGn6Cyn/6l
6kxQRUmlK7SaMNk9DXU1tJ8slkbMjme7EFIJzb1hkg6mHBKX4d/ob5hNfCpnpfLu
DBDXWZ+XTCPcyFMQkAMqA2UHJRq5RnCR5D3BdyVOXngGY+2PteDqsaa6luT2LBfq
2+qxJArnpSXJwstDLjQCWBoISTIKCwWhRpwa6hKJUStE8XTDIEEq/ajVEkPxcufl
PpGUU+tmkqQU1HxBodR1V4Esc130v0AvEZsNHHaN8gzKnVQGxN0xn0BmVhEfVat2
STOZnJ5mwktxVdj9eSM1yXNGI9tCu+RaEGUBAgl3XGFx2nzK3Hrqq1M/a60I0fzv
ZNroDJ16XvkMM+i3eaJeFfYtbwFzfL1KAgaZ/97UQu/e6GustnU0Vkg3Xx0Am9oW
zcbVtvTcFeV3xSNi5q3vP/kLfzM+HpObLg1uQ8vBk+rhqVyVPwyYKFMra06Gny2N
Ly3xR6ctllJmWJv6aWZbx7RLJ2Hz5alHW4BQrAwSV+kUXTr9XLVKo8F/d0/C1rjO
NdYs8FO+K0sysdfgkU3mwuWUemP8Ltte9g/KkuYJ9K1OURe2TCKWDlUkFouSBAMo
CI029FibcME3R2QmHCHyLnT0VN/MhgR63cTAlJC8VPbYa8KsgOrUZXm3w5+gkyge
tdYRp+hp4UnzZpmSGYpk5K2HE7mAhKrU7xCRbsSyQ6x2kT55v7RIFXDOBoa53lQs
ryZp1mtyJObNyVfzIM9em8BUpkfLHWMwlFnSj8PUg4l1WN/Sdq1kykwjkTBrpIgi
Gsm0B/86DqvzXwBldbX53+NJoxaC2ASSSfn3C/FW0xCDBDkfOCOLzXiJhIbBg1xg
Uj89BByvL4+x/8SGitlnN7ufxjqL+wEopF6HQzRfnIF+bsjg5AzGvVdUfeTsxrMg
oTBXSeYoRf9vPGFs8ZtdEmPI8P+MQxohWlrIlUBK3XuTaREFlow7kqyt14p5Sp3o
gKLxOHOjw63T1TfAiSDvnU/i1VP3BdmWhBa5jKRQohoMDVwdHRBNyQLN7GV3A37q
dFRe3GoHM/28rMdEmA+5SRtx1CKo6sQpeO2QlUpC0ggLcBuDat9+uuTXiZ8WpDf4
WQ51isb4OCHy6Wd39mu3s5Z9R9mqYUUwis13nVSHienslCGaYB/PAGOWcBNMiYx+
l8oyXR/gCWZ3y/tGl08HUuYBieGCywcyg2bV9njAlSauXtY0luJUt2gtdJW32S/J
06EFe70OF5U0lRC1zuuWbV5K6kALfjtcmHn9hUYWFAEnzV6/Y5oEO2wGVgrEDLyi
gXPhqMzCMZ9jIheTZEqkyjXw4YZEMlP35zqt1aQ5VklCI+c8mhPAoCJzDVhfF3OS
bGLLYR0wVTBxHLZUcY0mRSsy4ouxQ7kevCz/192vBwljGaAySsQTr4392imPN+NS
JSzEqtT0ZDzJo29F37iIHeO9zJgMKQLqyFGOIy3B2U/1/MS++4Ma8H2CUiWX7JRT
4USrk6i6Fl2HY2Yk8K8Ikj2J1bCbqmzrAGEZSJnVfi59DhpQNOgRVqCvSJh1iY2V
lfPWRwO4SK88kaHLsBSq/bauLsLi50VfPu0HFmrNRm9kpAcFyvU3tdBk7ufzab/h
1pqzbNLEMiziSWl9e+EupT0e7iXEoY3EbjuG1FHEJJQV5+TGDf6CjqYI4BvyNwUT
cHr9rfU9US+jFC+u3mYdKUtpcQdbB4ga5m/bSXs73BpRFl1lXshsXhp9djXbItsD
Igmrja7eM5g1WXHtE8xm4SJfY7sCNE1D7lXesjaYss9NzhyavScOBcRLKOUdQr0O
S0SxZ5912Zs+HfvNTotl99TeNCoDDz+Czzd7v6rOE9wyvbw5fFWmNHHkHA916o3Q
D/g+btsS4gMtNyDq9XIzBdKBwqbcvgleFDDdnRzhxSpQunR7ekiC/rcy5RRPR4+j
4LfLwD3GfIijlBd++EhJ9T2voO130ZPK6owydYwSzlG2/w3c46T1KLNzg8gWxxE9
HIf6AIHBnr/NpXnkS1rA2ZsvMRhOGDStn7OL4Y4g8zh4NfnHl0qstxWoT/AeCeZF
Rv/dH2BkDUoOZ0ItMy27oWSXgOXRc14zEvNRIb6DC2rUBWdsjqeP/Rm33CiKrbDm
GvRWwRjQbMmxnWs6dmVlqmS4JKTTEaBjVAMJTlKLgv966OYp+ABcpxbr7AideQSl
9LdN3FH8CCVzXiYoWJYs1mWPBFU99VKqT12ts3gatKS9hskK9NUva7Z6DxXkNLQg
fEyEuyh+2vqZhQnLMV8BG0+qEnjkdRhsz5TtlVX5TZnlyV5W5CZksjhAOxC86/8p
80Ou5My4CZlV7S7F2u3A8YurtOV7UvDQuJ6/3DQvdFZ2gJxtV0EGHdJLRLturGY3
4/1SGueRUzbHgHhVOUKqGm0Gn13whEY8suRV7q1mjBrh1ibGujF/2gUoIMny9gW7
i6iMcRcBZYzVy6uhKHOGqICFfZjUIv4bHvQapNKQQkgeljhs/trOZd53xg3NpDge
ABmkhgdiaJIa9h/gLQCcAfaz/+p4s0PSoQL6ACWx3fdKcyAF3+DanqIw8JXI9CJx
ZkrQY9oD7fblUkBO5YtP3STRlfZ2KXSPVSmAjjnzdcGbOZlQJCN26t5m2InXDzrK
hyNonVSgwUXhEYxhoPaKzEyf+ThlX9Z/pqjInwtBHzcCIfoO4aBA+6AT12mwVKcY
nxYV0JbBUW8mUntnqtXvQQSBKSrDtq/qYRop6WselMbVAbcppuJcB3YzLWiztI1C
950DwEYFdVeMhNR0eX3M5dgyz4DrUtO70RLQhdKVa5nvnNtaHrqRZceh4lvwfu0d
GhmlQPwGHl8J3GO9pnPOTKES2DGtWGqq6P3XMwJtTf8NKtXPouT7hh9tqlBiZTST
2xtwpWexLkVQcddb790/HT0XK1QHzoE4OJ5maMKszrvDXaIRhidDYjeWwM4CquB/
/9B92fnosbaTAtYglmjirR21eLCJjv4sMhiMxFitjuCDl3oEWSXstqq2tA9aOv5F
XWzgDXAebxsT7pltMXfro/FpptPdfUlXuqagHB7Da7sStPph8Bdopqpx1cuCc8mi
4JRsfsARdRQ7yptv1C8/K2JHUDqGrA/Q3yt9Ptd4wYY3ij8g9oXgT5FFTQpjbtYe
zAS8DyEnfrpeiS/BF3gIEgQ+3BSwkAoO6nBSpH5FLYt0ZqPo8EG35Lf3klTIyzgI
T+ZadXpHmqKYpi83ixdio8RLC/MDeBzQnb1hE4WbrtJAIyWZK9uV7Bx5rKk8m+Za
9Hx5bkQCdGa2pXR4UX/m4UDDzXluVHzJXwrDZWg4iuiUKDoFz82znVkBh4t1XkNk
eMVhQlNRR1hUqFMe+Gqag1BdPGwlaniZ049PFRseRITPF23uPSQ4D8dwJfsVUDG8
PeXiZaZd9O3VmBduzMlgbC9mWsUaZ5Vyvlth4H9BunIz5+93aaKSeepXQBwzs5QS
eEuvSkygiz/NEwuXFWycVd2Huej4K3w5XHXFdHPsx8YNv4+2rUVd9u0UUn/yB4nk
erLTR5qj92HwRAMGPO2pvua2vOClotlkN7a7DvmDQvscjN2IKAm4jCmOY4WFplRp
zmMpmKfmxSftRKSINwpFmWBE/EQCtOqX9OL8A7ghq7vfJaScGtwWRFMv7kAnqrQP
IHnHUsB4t1Nq+zbZuV1ijeksRtMEXRGynY2DynqKUbBrgKRFsuvbEnjt5ZkSiYee
65ksfk2Rp/zTBiAthwYGY6moc/aHRIp7WDXjEW3TtXrMuL1QCgAMSbLLXuWtr3YJ
FPC6KGGXEQHcymz3vPDnV2nKQK9NTdoI7HgbtPKGddPxl2iJX1hBxsv6HaTANUFL
f9FAsa3V3B7zxF308BJI1wjCNN+pxjDuLjQLzLB3z2zOo8UKVmIvpcbhRRRkV7MI
UBTJy0FX6LG0jEar59hOlN8cSJ9hfqQODYcQIGMw8NcdqlzYQtfXvClUPlIR8c0v
v3aeOGJeaPz11X2Uiq+Or7HjExudcm79xlaplUBWHsVsLd27mQqN87Iy25vlmZn+
g7NHmttkZLxtZ9Bnk7hELZKz4MW5FBiFXcP3s//UBzAeSNO0gHVoZ4h0HYmeY6BX
XGrNSKZdV99he+8tJ0RctrfIGhso1ctriIxCxdGUL7xIpUYU/MDnP5h4isRGGvqk
924WZo6oFf/LDPf0ZoD1zDemQqwm1tNkYHDuNO9LtxPf6UlQD4dFLBY4xpXkV0Th
PVAAxy94g7iTA3WxQc1G9lTJSAtHoXxIW0za+Wr2XxVKrwc18WYyRy7YjIL+zsVr
pOzjYcTb6wI/Emxgbhhq58JuBWYAPaL/vADItxqETOhlO7JWqC8j54haEpvL6LIu
gMKf5NauUzLtxdcWGKHvOdOh8KLI/SgM7fFL62a9sJLnYLhHVIZ0q/y/jukD7ArU
Qzov2befdnyd7nhFc3bUI700c802LLX5UEqmGu8ix2Ij4Z5x8YhMvpFiEEUnRmJX
5SDewmD5l5WR3auVKp5q39eyLNMOJu6lPPy7skAqgIM9JWvmtiWTrG0oALDSXG0b
//H6rxXOB629p7o9fNb5yXTbv1Tjs9wUbX9JWTms3cEjv2qX/Pq+w5ohmaFlOhKT
nnOub92dCnKUeA+rjjIPrcsG53jLTi3K/tiuXSZ1B64KMDhSXnVCdnnO5kuSTlwk
jixI2cJ7yfgHoT7M+VqU2umJENYNMWxhOvhHj2FTT8cHlsXtHtBK4LEr71iOhVcL
o0CQ5JLd0eWJoRPDumkwNkb6fZUslA5w7ybUcxvHrVsKCUKrTnt/GxmAr7oY0L24
y6u9NBapvukjSmga3G7Nse0NXxpV05JdcXdUYr/AFscfmXQVbsZOdz5kxjN3xG+e
FAT9ADCSArSVS5tIjRxPX/E+NgsSIRdKuIOycX8sQMbeu+5Yot1bP+4/CZEVIMau
jiXTZSLedb2H2qBKHs9IyNWwUX+/2hqqoieBj+gC5DDS3ZKN2buIMp+2PPPNgCz9
df5ijTrg/UqiTaCuBtcjcPsRL7D56EdAeeo5/7eKzJHpQQclOsSRRlnQDTbmGXWz
Pdljgel9WELh4KAbQlZYreoiKOGdoiR+LcqZPKml5OdZwCA+KSmyHUtDq5Dn0d1r
sVH8el4QcnfRNybCaqWL6Vv5ViwWsaSdW5N5FBi50xJvY+JZ7LjvKvY170/qjBou
WIvWkQKuLaY4hkEP4ikYoMTPNUayVMKTt1WMSxwTfi1UHS2zln8MWnlkH954Toeq
uMtK70o6LLlHNfixrnyDtsK7NKCxlChzErfYH4IJv1/6fDgdHKof2ro1JLvnuUw7
EYUAcIi39w5BwgU2tD3BLjQQ38JF785JyepO83zBHNlLSHSiRf6s0fLB91iiX88S
4+1WpzmEbBCHV9qRvAQloFDH81wdIXxYBBJ8jv2vepH7rhyhQqq+HRC6oIptYE6O
XlU37QF1JqDLvxI/2IpvichaP1HyXwKI77GPg43hZwM23DrKuOMPcxevgnpLzmK2
IWaQ8+v0ZwbYrLbygwtEY9+9NG/+//Ps5i4BvAQo6OQos7BEux4zZEJaTpaXDHKg
G33SKaY+dqa6HtD912isHDql+vKASB+FeImLS7/QMuxDQKeXVQLjbVrObZOlB5aA
CFgyzc7L85rYqilV8DkgxUm01NHhgldyI4GLX9QvlP9QVlSJtCND6OODiPfKQI+u
Ekw+jiaTshTO6BiVf56EQUzDvS+BUCXSmSBlU/Eo6Yx+lwAnh58/JL1DV89ewEHf
/EW0JAAIGcccUZtqay+E5+kf6fJB19MZcgWAIXmPiV+hJcVe8D9Yf10PzhcM4srG
7cbc+Qa9TXTcuGdyexS//VHI8D3Ez3AJU47wWwd8pZtHAv+dpCbefVYQogEV3Udz
q+Q0nTRsnq5Vye5cLIRWkUaUuGwQAOJpE+JZ1qiCJnrQdYnRtYPYpEfIGCbrEPLu
tv0Ce9fWRy9/Rn6EICmbun7nrwa8BszBSTR29l9rkiTcNSIpLptHHZyySfqvFZvw
RSqsIyiwhsakyRh7in1bUpEtjVMKvBhUfM/jKejqkr+ecdlRePSZsUm3XvnUQNsm
MzaiWheVKOIkrlTlx6lSWY3QIj1gtGtXbhFbHfaHg/ysnyLFTTALLx0AKT8vGC0u
1qdbSowd+sSC/flhLy4cWvRujEsGjiZuHVD63Rx0W6ouBYBOT0NHmCluFzZY1SvU
VcZUdMDB2X9tM7EOwKLBVtI4ItPn8u2/VQnnvbdf/lDw0bpvxwAbOgJoSppmwL8O
yLpleH++7Ti1xfQkrOiHEomUgCB8RpdWAJyfU1SuAoJZZhPjHpntYdDkPfOGf1Xh
DsFarNgt+2/S/b5X/wKxfu1VMbEPvjVjrWUnMbIgQqPZqi4nusao+LbufvA5dyRt
8bRpy2nPv6yORxSI6F8jkCn8LBguO3D3+/SLHej/KWyRLeBFTV5waRHViAL0WwSx
y8wA2OFnNFALP3rU/6tMRXV0aBOY6CUscRnSeiW3w4fL2ObzUt5ZHhYAfShHWfPL
VoNl1zJJyTMs4QT78ZBtcNNkQ+aMr96t1Ms3cZRCLqVOE7rczhI9zoYbeAqpAuKC
hANwKhv3hzzus9MymZei9a1WKBIWGhvq5fyWCNOQpxpWgGhm0piRC9agzirzWpvX
3KcXDVnYICEcpsgb+5az40GGTi5VR9qDOns6oktAiemTd4w5bY7BFAD32ghWO/7i
J8TMbKChTGqFy4qOrtl/NiBqROwqErBtwdUFKThmOXcLKMwycRk7k5EFsk7NgHEd
ZskWOo2CDWBvXGX2z/I4tlc0GIhJNPJ4ss5bXTWSSj7ItGkbEdAiOX4OAY+EDyMv
nl3VthOKWURKQ58P5PpNM86tMPi8P4aKcc+rFnO+FJsKUlqb4RtQW2FwaTreD7wG
bmnjv1aCyGOtysNyg4E1VkwaJy+xRDKC/vMSjffPF5eFK2Tcc2KmAmFuv4MnPaIC
8BikgWExzpNWUhR+oFjxFy76vXkOZu9EoFsE4qOQlZwQBbwdQvSxIzmiGErx8eX7
9KK1TcNcxJUlk/BRvheCrzvLd3TdclGpo+I3ywqvMbo3XV8QnzfCHSErmZlRYq5j
0AEvO45AJFmTI9iEjqge+qNmN8Hhc1ikEr183vnskN4krAkMo7krK0sevCh0r5pP
9dVKTsYtO5xqMxNEkDI60z3YqUTOjAHxp3L+DoyLVVz7yWBVKm2ZyTpYpxTYvVhH
PjEpHzu1Ojd+NM97uQ596FjhRgwf0i4X+bEwxKXwz81pEb0a5DAT5SnPDBVX33pV
lw03WmoQmKD47j4GFhkTvvjzptJTIf5etmlNdVig6dhpdQm+fxHDmFaQyO8UFMDz
HGa98rozxajyrCro1Qwly93jUNlcVUMAActB5jDU7tq6HYZ/eS1yJ2Lyh7TaXwQ+
U+cHerb4XuzKDhAOlgeDBsaG7Rb6uyPBAnL0wMPQXNr6NZc4vPSV+g7B+LQRTYSK
2Y6XuBHZ9Lr0gfkfGgvb95Es8lz/xnKHdJmbs3tsfl9Iv48/ZrXjT0GvMd26skOB
PZggCGMHi2rftaPXvowv7OxBkarOKU9c7i63NPbaT3LIdwruRUC08LxoeZVT9ZPE
+GQpb66DLtz9TkROe7ycLUDDbrq9LIdDvNOmVdEjro3NIKeF6ReEmVRADFXgT7ps
pSkxbTBRCcCKAY1+szsSsec0Bb3IpE3V7rqWWDAnsMe0V7OSee4UnBrQD+iPTRMd
FhXAZ9OLNTG1lnO6LCiPgsfmDG9yPEZ8Ta/qtLj82rTEMuHGuRi87MAfBL0zYIwy
ZnDWVO5PaOC6mUz+T8gupdlH426Sv85I2CXVpXdJzBHtaVNhT/zXi/xT5Wk4BnYQ
uXA/7suJLymbgxbYtHQBO31fxti2bB4oElmXqaVK/1MmuBRZEcImQ5Q+gLMeT9GW
wxpdD988ye39jq6GXq6OteEJ1PjG5RJySCpUtfhwPHeO8rzqoI0mVyvvV7KSj8bV
b8+tQVvQtWTOSiCb1TCOMnOZBB90GnnvEyOxyboAYvsQX9GJKzG7+UuNcuZ0UNBe
5aTXc1+ZOl2yTgeaLr6jbuFsVdujGS+FvTUu1ZPn/hBACQIwnIBg4+kmA7+bNr3U
nAGSZoxzoniOiPZdSDDI0k3xii49i6gU6LLDnu27kH2rjpE1eKQPj7NJmd9v+pHT
PNUOs12QM0GPFTesSKKbBdncGo40iXzWRWAlOqKKhFRd2uyTGGI3j+5xu3hALDtl
i21tj1iH+2hL6pTdPY34NLoWDfV5e34h9fekVxj8fk7AXzm2b/I4hRfGfkP1ZWi5
d2xczGq6UdtUTPfU9H7wWuqa7ZgSJHnQ0Bjw6QD0GmJfGM0/g1LH5LuVHY1pmqZs
xTbA9G8xNT66DkN1TDEjTDhh4sd4R/Rrhidwmw5/cs8St3W6XnhALNlReSBvYWdE
8svvRvHRd/+BNGMmpnoam8bD+QufLhaV0mFQ2Mwxj49QNSvzFCDZma3ieYq0d9YJ
hB1l5fVf1QYXCS+bx53dNYtvKcSo0lVqIZJXe41CAlK+RyKxNU6/Q6/JdKiZkei3
3i6R22CaT7RTT+JK3t3oKarG+cLU9uQGax9aMscQiAziPkvsdQds65Ll3k5UYauH
e6/fHIKvyHhoziATbF4SCP1t7TICTXxA5G7TgTQW2gu5LapQ23BJ/D0cN4FFGnXK
EQ8NZEEeMI2chFcod1Yyxx2KR8D9Nnu/xpOd7ZFxldOIRuD54pd5HxlWBsnEeJ3q
N6XoHupUKu3h+xuuuKSEFgei5lcmvIgAuNE7wwuVSvo6v2bJBG3J5SiQnhtFgwia
KP1didVfoLRRX32WqzWCCqjlphX/B+t2sv1lXLTcNhUfefZie0O06QLreMaelzFP
jfcSefjPpfkpdrx8iqSJdsddi9VdawWZgijMsHJawmVlAoYal/jaGhAr3MRaunFO
f7irX+M06SGoVwxzSS24zjQQVWEcIBtmWamn99uIvYPmW2CKL9Pg8Pk4Xu3771Lv
xKhnB55DzHYQ7TwSXGRAHhYRcUO660JexPh5Aa2rYPWBhUMM78v5WjsNlx6WJ03s
BBDOjB6I00FcHsQnzi2QGJLI9aMjk04qA0qw/Aix774o0CFlgNhBrLDplAeQEMp9
6LaI31euHz5GcCN5b+xF/1ud1J1oO3gO6WhEwHms6uqEJuhSE/LX4NTTQhPMTlL8
6cmViC1z0vPP2xdWuHqgee7v9J2r8CAC05pp4W9AB6J6ZeQqPpRqWBor6ya8y8g6
tlKiX09OKptUB2Amaab0EZE01qjqqB8ujlCZcSwFqNUyHdEIlRE/pFFgnZHeEhpM
xWSk2V0APF2u1FThdelKjk3UkGJoVydAZRNm+tIDEWprpcPHxkvREjybYA5n+4kO
6gCk8/cXFNXX7b9jJPC6lMVFnRsTxCaNOX4p6COG/2W17rj5ovVK13/F3DL0vl7Q
mvta9cq6tSp8YSV1yaWy2tFRhooYxRct+exa1JQLYQK/NQmZ6nWj70/PJ6TXHNWt
xhW17S9D5Mto9SK3ftFw/LBvFODZx8klTKbga2/mpI1Z0xdm3yEvtK09fLZDoSqN
x6vPh0zjWBN+h2Di7Eebuy944IcCAEx26uwnCU4VQd7KyCZxgsYrDChXjUcQicmi
j4fKsfQuoncw6QYokjtQ/fizLoTj3KGqorvpGe5IKXWPbQHUs3MeU5nC0sLg1zwR
Y50+DH5ccyQoLOC9AagbgnhRuRe/TiQYIGerKrfDYpMHn64hMOxleUddFNSeUHOX
i+/ofJgTH3N+xUdZ7GP7wQNfeMoFy8gSiNm6lRNnu8iGxdrPHAISqPfhpi29pP7F
RhQ6qqPy2IFCQXq4kYbYbBjBRCOTOCQxDSKa0Z5tQ8TfHiXVjDXNOegJc1wiTRuX
HkXogrVct0enmDUIpip5Z1yVLbK1m3y4Y61d7MWazjk3XBCkI9Hwsz2erEZ/0Rb+
kbh2jymdWuqLFYf6qyhMQcNweZVfhGl3bRnndNSdSIb5dawTjYm8xAo/mqnDUYAR
TCIv+QA3U+x5CviTMIS6mioSipukgiR6oBMF7sqpobmwTo/DOKTvUrdadV2yyp4e
LHKh74gEh5JkX6NZNsmatGRaAyzBRp7rx/CTUAgifCSfYF9SDwuywWzqocG3iTLt
NcUoLyYfEsbc3iDtPDL5JR3F6bFfRPbA6/n14+ltLPtR+Y9ZH2g6vq5yjFwf9DOO
Zn6Nsxcjt89zgDyROI1o6Vot4Jdrh6/a64/njKzIJEsOxtbRKJC1z57+0QdiNG9S
VcDgEYZhESquuvNPd0gaG3nBkprBLaedSqV9yvkp+rc0DhOE+7VM3yMGMnAUWjlo
8DaB05iZfO6qjlP7kuC7sxR4bcQxNKgjiH5sC2mWGAALes9cXXAHhRjjtZL+pjAy
NV/fvmsi3HOIrnWjLYHCrJilL5weqNa7fuVFgnCVMIFi77Yo7MWvwZheNKZbXDwf
TFakrZNLVj/EJ00hS+nmUdMqECdEtX3q6FE5l3VfhiixGE5FD2SIllXKaRswWAJx
N5IPeOr5vl6KZ+X2zTJ48wLjzi9M5UOqGjyjYpqUXNPaEspVfItCJVmZfXtT4izm
jE7dqFE9REQbHj4+PTUcBg+4UpFTo9VRroaOBkRk7P1efcL155OTxNb1WUhcQUq6
qAKDan/o08S3FF7SfKvTWvck/HzKpfH4HFyp8fbE2wgGZMlIIucw8qlZSkW8S/Tn
Rqmby3chrz2ULZ9pdWp34iJUDd1YD2reD5o7KhUcZL7g4+PSrQYyy7fdet1Or53t
vgaD5vvMfynQ+jrjV7dDKL/wwcQzCY+1GKy84kj8Teki3FDM6cTglzy26rmMlLQ2
XAEpDUBvRLgaw4HAylV4ztf3VHsJg0z9PPzrK9v2KEp+trG6mIB939NLli27137S
4OruUeKYL0Ca8WHyXOqvKU6pK/G/3W5TMzuBjDvrJkBlQO4E4wmcUfdvR3GpPOV0
RI6vV+8haXd43NfBboEKXpdsc4gMj7pJzX+p7vAFM1hTgAbBaoGnA7as9oK169Za
Vslg6YNqcB+ykSxRtpIqWlLrsIeYTLnLXIdupFUH0Z8dZYjR5L9XqhKX473zxdHY
Jq3mNXmpffFl3f/MCXQEUprRz/Zv9IEcl8QQ0o9dE417njZ1oNs+3bS5q5CSG+Fk
eVmDhCHj+pL9OafWiTlcg+IKruF3ZWko6vxhoXRl2Pdbaxb89QwHMJNBvnRmpn3C
mmKAyGJqKrhl+PEWqeO/fh2pmZeH+qlhhhLgzQsNL4NV/o1skidr2RMK9jLxeeew
EdPFwxkHXYAjf7++FPjEQ9LSNFKrVmTU3iqSGMs2EYknOiHIFg9vb9aUb20Hb7HJ
q0CzsdwaCo59H8TMqnF1cgLfaG7fJPiTbWn6Y19OXX/WZ+s0Q/FpNQ6b2EsHfzep
28U21Uyk/OxDPJcPIwd9c79W15gkNpMdHkWqtC40RI3M+E2mNnkLnnu74v5/cRc+
aEbgVlr8CfiOAKbkTrRJ1dPjTvgwHPzkGpzuswD/495Oj8lmSAVkd7Ul2Ypq75Z/
xkFN9lWLJjASapA3QOjHsuquqbvRuNiK9mtKtfL4FUmQ5tjYBNyKB6poicEMcasn
wSjrcgIZtjh+uqzfeqbAnVFAJQKofISb/IK7QgCLVOcxe3QBrHLO1s9NWvI5eRJr
Br0ZFdmB/jWmbfhMr3/SLYBCwT+ZbPJLJ65SyrLvxLYy7+N1ihNJzdLsvoRYbPTi
udSsG8smi19ST3A1s30OhEJentIUPSl+2hYZlLNXPf8BUEV9+HI/XQVlK0+OV2EQ
D2yUHrbtn87QWXeVUDrUhmJ+POZDsDUYP9g16E4MnFgxUVNg+dn3G4z5gZkmk1Dw
LxMtAIoeEWSTwgJtuzHTXOM7whLZcFoOMWEyxm5mlKzTspUUAPKeHD0FF/Z7qPhZ
ET9jK58iGs8aOr60WiPqC1oWYv4SwKxlneVrSQMAxQYaL1v+29eXPI0MXg4ID872
ryRLbU70BDAyZvfVwiJ+DqMGY+giOgkXmtDlJTUpng+71yZrrk++gCTeWcRsyc6f
9XhJc141wYTCOQ76HT5MbBOjOVcZH11BgfpuOxvMcSFjQyBOYJ3fRuw1K9DWHAgS
tMMeuZzGKpGN8eCNZzdoLFTwow5ypOVuWNRsOYo3RXxhZLxi8pfaSPY+wz845Sk8
8u3C9uUs9vaIVehPEP2wjM4AzmpEMS0ekOqivOl5E1wFfrkkpcD7zc9kh5IRyW4q
Xp5V+3w5+9vLGhcOrHo+4T45ODemViOgRKAMn0JAdiU4Z/amx14euTvMf3GYb53h
xM7wozXcgmR56H/xwafe3RTTdAtg8sX7KmTC7NbwXyfAYQsFHQ6GZupk8T5X/OUR
/OmZQ4a3qvL2o4TkJ8mYRf7vNZnXnrUCBhgWB8/R4l7gvmc+bcynlSTlkffBRD0K
ZyBvspVL3xzuTz/y8GSu+CD8HL+R3Q7tnrpFtT19h1ZRp9wgNe9qYH9yn2CAWvfU
8Wey/BKxm8xGlcoCCeuxyYYsl4BvlXk0fRPFuI4aPkF63ntbXyTpSWPTan4ofHhF
BIFa7OLsueGB+Y9Pl3s2oLB+HB4Tdg/j11LNDUZYWC1vpkMjwuvEWr5MCQWHSWM4
ERxouwXUZS0t4gelBm2tsNUo3ZH4FnFvCA059yNUvrGc4OTiTMn+KdzhT/VED53e
FsRBZHGzDZ68aHK91FdpqN80nyuA1zdgZ8g9auI5tH9bzl3tilm4y38JIktWhoDo
DvSZ7aYH/laEWKQZYmZlpVPQ5K32O/bE1cTpQRlzGLyH3zBJjl8JwfCfBl7CW7OK
omIOjNgwlTHhGEzKVb0+oYTCOvPQqqGt3bPaRPnI7ZO915S3AvC1FBv/CJ2p3loC
MLZvUS4ocik2iqEkr8K4sbzc+I+OIa3TpRHc8PUuMBUXiUCHw/ImmA3MxxVKquX6
G4W2jf99PFf9hzx4WtKyZg0Xj0inrYfM3dSj7p352G3U/Feb8yunKbLZxsRlQ2iG
92oI563K+J+snMhrTgRo9Qctk2CsZ+YXMdHr9Jqhs8cXqqIlUHnrld20YDBm21Lf
tvDyT2TdfcGkYdI8+ok3w30cQU9+yJUsVXkY77WKRd601t3R1fJKWucOFhsjnNOI
RsQJv/tOTps0yQtgxhOxhf9O7C5wLqG5QnAndO3tZ/MC7JNURNreLrrJ31iDtm1R
LYxMW74tSjfAheid8yPOqyzBvxqPC+0z9D2W6sWKCta/A/It+BX7RphP+QppSK8o
glFYzoKxbRtd0BXzQ4CfU6z7uKb41Z+M6wmwlODVrAopcBPcTMOBUH70waDjGgwZ
24O0RX9AdICMatEnfJCrKBzw8q3LZfGA0CO88bRJpD75+IZYr5iQSucWEPhI3GGu
lO+lSufvu+2kY6LJ+nS+2CucAFpn8L6sZOSQTzH+KICNn1s9Luce06flPK2jzjkm
yW94kHgZ+AQ1XivUJX3jyQb9AsWsXRyYvBOPsM1c64WAm7v6UH6mi5eOz+ZZjH2m
DL/LcZysaFEzQWKzWiqNBJcIKnqZncBqxcc0QkM863xo80zhb7H3pH6cO7gJxjfM
+o4x+B4b9gUj3O4VsKj4ITNwmuSgK0ySX3UQSo0BfYHdoq//HyniOAiriRWjC4Sw
hF3YfWFZ+NHeClO/qSlcTO+uNSVes3ezFGqwCk34fBeBicxttCvT+8HfNZVNCrAh
iCNHJB+gRIlV+H8r/V8b7RyX82GypiJp61fMRjpX7hNnTQtl13qRZtKQdFzZ9+y+
5TrTIW1oLPEi4Bn9Zy7ea/OPLSWFjSik/Mfq1hB/E57Ur7fbWbHzp8GngOrB4GN4
FZywfUxdTB2kzFjJ7y6SpOHK3Dj0NMhzeDDCnrlICtfFqJfXhil4D3qmdKHpIuxw
iXbcj8yJ6WJRqNbnjSuE6YslaIA/+p+YlFOEjFc25dmPVEYsRFdAnxypO44Y9Qii
7bb4IiJhTt+/F+rE/Odu6htdKFzain0fks8h+L/1/Y5uzXQNQbF6lOgq5Z7nw3HJ
lX7rz2I+fvHILlBLb9bFsfSg/Autpp6vHD5pXdE1iw+wNREqyuZuobiaoTKTXyFc
W20ddc1WgMPaX2Ye4jb9exJ+P29KOc1klwIZQeoMCYy5gbV6pGPqZUQ+j8leq2YY
hNg6zrWBLl1mikHbPW2FMy0lTSfPSHGwS4pRgcWm0scNh9Zat/gMcFyxYZWMGxq8
rNmUBQ7yqnbKOA+kt1ilqGuwOjO2rW/nNEJ+ZOAFxS04KdwlinjyzScM0NSnXHPr
o7eOVmhJNe07Eiy+5f5yARqsxBlR3H7C/zeCbu2IpCV8v4y7HRBGQ/E1JYEFWdE0
MpTXL5P4mL5aqhBHPFTvCowJv10ltCpYeazrHt+Ir3bVzyzlUaKu4cfiywvvOZb0
70ppZkmdeuoJ555Ub8RK3IXuLEqftKkrEqP/tnHtdvE5W/GprUDGOxufC/4z7w92
YmjVqz1GWQJ+WuKnlky4E9+g4rmkyvElUPNeLqaYxb2VY+inn32o+yBz5ZncJAOC
o8/tfmpR9bakkzbHacz9i9JAG+76vdQ0840fSqI75zqforUrQTV7zVlVu9ID9uaM
vjgYi5s4cxqw0VKQaNZdEM0tP8FjNHbg7jftjlBkyqXmR6oQoooEQEhhZhXbY+0F
+vG1V3ibl/X16jla7DdvY+X/tMOdEoICzbj1b+xmpnFFvzY/Nb4dzWNnl22RncCS
cZ7Gg0cTv6ZE45+FtJx2NS+w+IBbdvLFCpi384cjlzB3rIlOTlOZpFMnKSL1ucQO
0jZwR5VXTfZlGMHYM7CoDBj+gNvepWO0RhADUXraZ3HDhLjQB5YAo3NFcItSZdMB
JYKdAD+P5I5J9flxI7jEM3L/0nsqqtH+JFzUwq7fjLv/wV1jqz9DfJjnGMTvJotc
QQRtmSuI4rV287CeiPp4lzmaWPEMWiiYBiZDapGjDTYu1XUHTBzuehp5G1eSNG+r
Lt1az86JBXQk6wDhMJEmJgh7thdq2MlP8QWxy9oAZYxEaGw5Cr2P4SORmonlKRQm
MGwpKeXH+o44OVKeuJGEKFKCszj592rI49Ynbcvm6v5IUfCS9K7/4rwLI3z+RUn2
rAXqwGVSVoQDg1aSX90e2n9JCfGadzaYQ9tBZwOTdPtzk3xP49Z+ksOxulVFBThb
WAMSM+bSlcz/jz7HscmFaZYGDfZn8+yzIhdiAwPF+R6AxxKMwtiR+jrP8edhuEH1
TwVPsnCE1fIQohs6BhVW2dNgg9JcWzumzij5un+ubfPpwRRzinvI3w9LILImuWZv
MbN7cAUYbR7FdH3JaSOPTHJNRijj5ehrJfYUs5pSNdAfFb7E2HWxNReyUVr37QTK
TuJNs1gxp+JNQiyccR6Rloba0sVYjWJKsVpzr31hdBSiY92Z6BoZaaVnWCBCZNdD
1llcSnfsM2TZUnXYHt57kb9RkR9dWNbEKW+NUfTrxhdONhimT3jw2C7+02tNS+VH
GlcOnd/iUt8uGZ4gWzOcGn9mygYCJOgSpoEpF5Zv/8nSvOQuFTSVoEeGd2P4MbyE
iikh1buC56cc8nY+rQlt4e0fj8Kaj3sAvAJqcBwdgJpLyXAjiSAVeQuox9zWa64f
GuiaOYXLcbxXPbf+p3j72eOInsDOMcrZfZthLXl3ceYalRjrPJ8zXe4lvX5qeiS9
+R4PBSskbNLTU33QHMqJqyVenzxxTsZcGcncO9674STNkE9qDS0wdqI0WtXEkUoE
Ai15n99PAIi0rVwY6cEo+dWQly3MfkDY17ki7itxHBTvlDsE35Plf1Lgtg//KrQs
bD0zguPMDn4nbegp0iMr8pq5G5xcsjscNmDWm6o19PeAMI2Yk1KKXuofpyEdKCpA
4JdBenpZznObFL7vPJmFfHZgYX5nbSz00HTlvHZoX2n5Hgd8o8qWjhd7p268vror
qFv33UktjqKY0T5nSddMj/7PPa0pzBYAidyg67lx+aZQRM8PxFgXqhd9umDuXNIi
7myBTzNEX34I4fesofvFFS9cbzhT42Fpdc1+roIP4//wPHDDY6uVfjOTm2oK2OA8
AyLdR/kmddXwrBMfAiVnPQRGrToYAlbRvgVTCdAcNrHYM9U2Y5ixQsFRa98JrA4u
Af/jRjmkDFgMX9LWJE2B28PD85z3oMpo2ValkMqx+a7XW2xjY/HwDyO21wlNlrOZ
aZxe3+8+QWc8m1qink7NexweXFosyfEs3HQAz0iuCKfOzab9cwpY8NWNDMg9V5Lh
n5/YvJdIDrHcrYbSJBJNKLPiCTTHJv/WdKKgXxXgZhTWISbBmM5ZSLGVDsYYbf6l
xYNHgk6EmgfSFEtpEpjH6Eqjg+ttsVj+XVMw5wHRiKvgfzkvkHA9/36wRcm5VNbe
RRTtLRJcy1Ic8OsEXYYcQuKpcZiUbIY/yxWRA7wCRpRl107rj2NhO5xbfhNbMies
BB8H3gVGoNi+wL1B2uTypp2CUeHj7beQbpoozaqixT9PYRBS2LbM17FLw8lrFGGo
M7nZrXk0Z5Jlki91MQ6laZhaI4WOdjB9EkGH0H/llayzrv8ESFaXNv95I5BA6qgC
3BbiJH9/wU0rzFZbAYwsDI/3MTDnU/LegZWf4jJ0/7b5h2o7t36WCivlilHNcKUm
7Mg7qOokT2fCLCi/MEaJo29uFwb1xW8YTNSJZsuqWxy/oxYoNkIPGBuqDJkCFeXu
iV5IVQ38qWyw9KSnfEdIYfMSCWF7C7cMlIX/SdI8+VSZk6Lizdn9z6zZlpzUr9t9
iTUgujam+zE/6OcJ0VxQ140ziuWAhwj5YFJzotSjbYa8bo7/uKfkcpceI7yF9GwX
IB6qGI+4OLUhOehf9zZwRZyQDXw7mrKA4rbLrCa5eG9cGNImlFqRoiHt8mXbY59m
c3RQYP09BKws/F97SwbLB7sG4e0+hDhB/Qmxe8jI6180VltmjScwF5bNjh7BC4El
P6h6JH8ZkrkFsu8Vkwe4IrO4gNyr4mguX1ZIkQ3WY6V0DnT3Ua+/CXjyTfwOtspc
hQzCWDTW29GeWqeGtuKaHMVMpWqwID6Sx/rzqUMbtNnhsLaGNqAnidhmfDVk+Ovp
KKttf7m/+b7SSg4QttqfhMJnaE+7md8+yMF2Sn61GOiSN1c98T3eti3HqJswehz+
dSzu749UzcmPTZUyXjY11j5DuOxvkBfhfZew21k1GFZeexsgG+tJAeNyCJUIx/C3
Zy/yHsDx1PO1IBTLlihOVbb7jhKIEG5S38EOP4bZj3NTCRo7V0iqQf3MB4E47/sp
muXM7uI36dwCqlcmAdICQps3ppscRHRzrTAAPcnKqgZd3qWOEcKHBhEwVL89lNo/
zARc8qdzBxBYyYWBRZdVqeCBARIVRSFiuXo138LXQqJ07KW/4HFZGyjK09XOE0SA
bFbykD4FgnaxPis5kqDdAmf8em5DTrq6IhqTNNnbhvNj/Qe5t5RwOPTf4CTNbz13
U0AISGQl8a7eXzLRB0alIsJ4hPW8xcHe40/MtSQFDNkM+0rLg2jUJ8kiXW5xaj0i
ja1FenZVFkR5u0++knKUd81B4Kv5ynls+eh6bsyaf1eYDL+6GAt1m7nAmWN2/d7K
X70SJDE1op/9h/rsUpc3snnIjBgoxd8Sk/42nwYfOCk9P+JTM5jJSL/t150ZtsRW
LzuAGvCdBpd5Pzbwie85tUkV/+BQUlGmD3iSfQYYuFDEHEst/xcWnsNtURkbi7Ju
Aolc8biEds+Yxb3toB9WNWI/5sxRXMax4UihtSaRl34dlDHB3UHnDDoavfRZm53b
BCOkrSI7vLZiWMpm75y/okZGd/9+Km5s5jmN1wwC+8TykMWPI+C+Abk/Ty9Pc9Dk
5GW7CS1wpYX6TFVvKjVcOMcMyp5Bi+Cx6Y8VBYr1kleZ08a8EC20RCf49zdB+CtA
dgMLvsB2fCwNVWSovyM/kj8RBFDDG3HFWwFBMF/S69DKVPfQpJEZABKf5g2Ui0kQ
pIzvcM9oUsB89Rlw/gDYwpoPU5BDBwhYZcopqT9qA7jeV0udrc20SumRo5imRji3
SAzj8exnO//VeQMSKmqfUqHA4PvJu9NPb0jY5W+ZfxTvtu0DCDXoJAAEKQYfrTrp
eaYehuwyBrHTVqnMZ8sRIBVJPK2X/cFepX+CnK0qcgJFA6bwPK/d2SpjdWXJzuWj
t0l8WIfQ/yhFibF0LLKV9ve8NVO/a3p32wG2bWuAHqvNi7NXCxeBvVmkXM1CWzVP
Yr1RTqciMpHZcbUJ/8mGePrnPP/j94wMQiM3exufLNzhlu6V1PxBjQlAFBIHDcrg
DA50v+wtR7KCjroU8+RRlrT/fq95ncH4jfDP+plkkROdCmCWHDyPl1TNuIz1uMVD
aio2fLuzEfBGPgqVB1qD6sxBjH8nJvz5INypXrpiLTQtMIs3UpaxEpw/7xKqC7wE
XX1+nFbK90xzyBZGtWLTuOerSZjUfsImrvo1CBXJ9C9bApPh4kceoAsJAg9mT7Qi
zqqma8YhofFoF/KKZK6lfOP8vH2ihSD94SSlUYWEqBCMduTO5R6kv5MoHcjNYzs8
Y5B3+9uxNDIjl7dDT2KjNqYUceM9c4ubW9gRyEy3Ova2EoG9V4cZcKos8FqN+2Ca
JJZWrYB81NQKYtO69BgyMiYypgRFJksZOvZ896XR/XmdJvJ8GuqiclAS51xmkqIB
a5IprQeFwDJNu+p0SyfkzUCG4+yKDHBKchf3fb/M6AwIkik5uO/ktO5T+6v7tzBf
XUmjMvHLQdIHkoby0SuKHflX8ptK0F9it24sRRf84Ym8xLe4e2chG1Kgj0K0KFFy
p0sYEehY3uuezb8LPofT8+4kNkO61u49ITbcsOqenG1ox1FmrcP7XknG2nq2tPj4
725k3vPvrwQGvt4dtK0s8j2xa1wBxG2u9VLm/as0IqYiier8WjOKyHzBEQhbiH3B
+bDhkdnJJXhZFNRBBGi7Uh+H+ztNyAbD1TAF43PTizrhrDZAaDefB/dYFRp+zAkz
1KoNq2362QQvOI1NApnHJM8OxQNLcZpYI9AU/zplWQRo26IS/eDOp4CzkmMgSsIe
yJU6J8mqCwGKJvU1/IjLX3rZL6Fe0UOTGL9cqDYp1nQm/Tuwr0iMYN5ZDNIXO3Zt
UWmG0NFxvOSrYcq4/n3uYgxmRmPqBe4pQpwZPr2IWFrD9dkvjWaRU6ZjcqSWKUMn
cb1M39XErKUw51K79EFvy3fRc4Azf8JHZMMilMVP29tHiFbRVE68Tj6LZBp1EI7U
TTkdlwAz8ns2YuvfEu8Cj038O6ZKpl948wbgORQ3AQW63YTD6RVkbSDi1ZGtYo4l
tcXLAKxB0GqKnNGTUiz8XbINlN/kH6Dgl1h25wPMOoytbxBt0UCGRu1mj/oD2272
j1Nr9fzrnghLVAETPMiqTkkC7lMCresQYShHEvhHH/fXxhkmUogDC4T0bAXPDQSY
p7gS+lsaruNa6QIFD0u5JF8J36xeiawL906cLT95BPaClPwPwAeG10RkN3nYJaT4
DcAJ/iboPU/pd5GvHV/npgNsuLeG1T3UpdkgQinSvJhomay5zj+WlWF68nlxOTNx
s4MOia+c2GAD0wJh8OtyJtGovIocaYrTvOHm9T92kaqmbBeiySr2ZlGDEo3XFK20
Odc3duUG89r5TWUWyuZaukKhfFsWip2MH4nQUAESTIdY0OobanBHlz25jVv4PjX7
uo9pfz9R7SCV6J+rsqNxqi9erW5VtnHaTtSaQrD9zsT7bW3QhylfmmIlUDz6actm
QFEIg9UmJMSlqb2pp4LH2V7Xs4OKWYofK4AX/sPAPbY/APRGVbnKJjo674mgSSP4
kn/nj0aRvcCFR/HWOynwwR+qQ4NcFOhLYsuLdsCvw0gPVOnhYCPGRx7p4sYOLHn9
+uJufGxqnd2hZnC4z4GE+kshR12aoK5zcRsGAeR+68g8pN/7AcvSnMs09j8OM6N/
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
W9FVp5u2+IeyNKdi+pVombmngC4ZoKpw6613wLwlh7N9XFEjS0Nj7zR1YgfoZXuC
FqqwQ1luPos077vtfkGABW3TwwiL1/uKEr8tCMKUYIlix6YkgKuyW7EkHEwjqlLY
yI9p7h0BwORAXt36SO9UgJM82B+USPEVLPg3lz3315LtfruX/u96L6Uv0+OyRzp3
JtxIlJXPgUwRJXmuWcNc/L+EK3hIb4NLjbT2X0sIi6ed1UQyh7MKs3GLUyr+Q4df
3AB1DfVBJhLjuSf2qvhN8Af67FKb7DdR4VohLr65PkVzw5rWQ9TpZ3WvFtCpYLPf
/zFoq+ZBWsr/KEjl9T6RIA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6496 )
`pragma protect data_block
q0YCLUFFRP/IzVJymskyJ85UK1XxEi/3rMAofYdWst71wIvLc/EUtRC+8R2Kxtj5
ipXc86NCETWqOPpFki2RkJjn1w4bem3AqiMjcSLfUDdC9LbPMkjYrO6bz9MyHU+Q
YMj+LuMh7nAAFGX9xVfeHehr00NXv7iq6RszBK6W3s7jOL2TsZf1eP3VTpYsTCFR
t/WDc48gJT8YXjrEdpz/RVqmwTOHRT17brs2EHFh+sxXz0ATA5zrQh+2OapcuvXb
rW2NUQ4bn1nq/rUSykHc3gL7XXzHkaU716wr9XZxM1phU4UMQjifi74ii5c3qn4k
RWh5oG9KnMiPemv4IuTuaBagT7wQJA9YPImpTrQOxRjsUYUaUe4Ps1NeLrE/kVRe
EAZieHIbwxeXhA/tj6FsjRfKo8JNm3IEoXST8EYuANg6C4gTz92c8kX7kkPTVITY
/AvZuKCWiukpBbgci+l8PyBEQW7mnII7/v9/6KMGlRm24TQAFhtIbEWWrdr96pTL
UnUnrJ8H87kqkznfKrF0MpqEEgISl2rHG2XXryTYnrIC9fCL7jFhTY8+27f69dXp
bSPXSHHCEK9WgU5f0dQJWx/Vgq4rpC8fq1a3um9oZsufYWtF02xVJFInTg7TdMtj
DGWQFYHuDS53vAfZDnY4DYOsCmWOP2S8dB94puDhOzZ7VtZOdg+AOLXESN/kJWmw
y8xOTCHj0eCmKErRaLAfSxsUD4tA4Fu1FX5vT3uwq3vtkpmmmB7C1WuypioQvuCo
dMFZpNdwra3i0XL31A9hu4++YhxPeYWrtRMeqGDBhCebqvfhR7HSoK2h+YCyE6Xg
B4ufV05uDKQZsWI4wfC25FIUNR/l0npVhA+ACcTvZgaxLfao4vuLLuGLQFuVklC6
pp38VhU1WWjuOvPHt6QhIJOiMabr9korD3S3kNxP93++gFHVfGy5Wmu1zy1TlL5I
lNPKhV6QvLH8zxCrYUUQNfsKi/jGQXYgEn53ADWEndsKuHPPHpuiH2Zc3j0yGA/K
G2drDvbM4+C21wM3oampft0X5Nm9bkhR/derhRH63REAziinFTzyDqEQneSZL9Rw
1tLqB9V5vfTqvpDgwGdI2kdhoOBC6iv6z7KNY0OB1Rfq6IWukRaBcfbXLsWswUJj
qG3hveaqPERYX7EV6yMIjNjZy9b+N2fn7uaO4HmRc+uW0PfPEBW4yfXwYDZQ2sOR
Tse1b1ZgBKBf1khWlDXTBl6219ChudCWrx4dgGN15WVPWzFtEW8nj1LtvsJiSF0G
tr8UYqiWLBVyxkYKbxIdu7uIOErvScGkl2MrD1OcayeBcLOM93nbVglv7k9wVeGs
TaxNN1G3PVv1yVRRAv3Fl6o/qITkgopxrsL7BHR/lAv0ODQamjlm5yP70Wu5t5E4
volKf7hM5zkIL+QJvAxbntla1MjEE9l1giKQAUeMAhLC7t9BGOttv7pTEFLqAPgQ
gFNHfshLW4qXMtIPGKd8z0iS1T/tfc334mmbg0hNep37nXLQ0EvbTkQGvo0f52Wm
N6jsq3L5qw30pMvMgaOv92JHymR/rYAv4MZkrdBAK0Yr+sS9VUnAtvtblE7nuddI
nlp3mgM6X14Q2chs8/mXXZwiXjNZV0IQjTRVOqBZWms7gBQ7MP1S7Dkjs97EcHow
HFj4wfKqzm+rOpyCIb1GdYkv0LCKTo262RFaXCiUSRhPiMMGpqkYS+GFLIyFkC01
TniZHO0O9VkTh15hVPRCgMlJF2zYRmVnEfXyV06W8a1o9+xGuqVqmTUgu9pTKeFp
d+dqnd1y5y1Jkk9FxhW7tt4D03He79QbvIFd0lH6h5D+/aMX0ioR16A/l7BMFx1G
M3owzgM+3yswOVTshk2zi4jrbrEQa7ujfMFWm010AFIOCyhqgTaM8JwXLJGkcw0h
rf9l2qwFEO6cWf/Z8lFOxztPEiqBIyPZ0mwdICdNImd+VIDQEJfhyUR/v1tqJHRH
EtmW4k7DfFsdgNBLcOzDE2A7VZbRzkjwVGaQGqs8D8nkkjaGWpQOFp5XTigFGVE9
X4cyHK6pllyK2Mrzq9XMhPo/2+jSWtB6YgNOzUIaVUfL8E4WUOHDRzBfubw2Hlkt
8A1hwfIMHLkzXnYEXl+qaJz6jAcZl5CpJE5aJ5lkxOG8z00rB0sxWveskYd8KEYd
kcZrTlDGiMRyY0p3Hlf7MaJdlG3J3GoWSHBWDW3old4+BPuiZWMCb7YJxu6NhDvi
3BE21HDWC2JqXQqZJL41Rr8vmWBDl6CHH1eR+RH+fJou9iLXyihYMA4BghvHHgsC
jTSc0IrBJ6iYc77wh2qejhqOrDipkUUT/FRcf9AgmUyEub73rieX3twSv761Fynp
2atveoLdZUBSR5wEPPueG8qG0ZVAnG0zwCbIfh5kQdYrw+TwiJXPDLS1lkT7YnVH
Az9xBJg2Ud/TXkNIBPJDE2cySwOXqMrGM2daST8TCkl25p608GwQUzm0AVI9923B
p5LbVYPkNnrsPim2F+B4u2eNXKUfp8tsRFY+kytLcGf9xs1m/2ooO//qBu1DPLdm
LH4ziXWOAEaFCcgUKxT4cqUEMODyE2QJvDZmD7mCctUpBO0unKAF3SHDDSekAmjK
iWRzYAYbiAoD+684XEF2BOI24Y9dRwziV58jWUeptRdt69grS7a59VpVVvZ9vquH
vCJf9PB+4Lov93dmrARIqCQhhd84xGUQmVwPxL7dZkz0buL+icRTB9Un+JAIkD/p
YfjC7GuqeLidx2eZRpSgunibva1kBADYQ7axDx/y6Lm7Big+l3XR3jiJyog0rUPy
KTG38W6/P5ZMpvswexWKiN7QFKuWIBkF6Dv6M8DbSGtHa40V0soE3zhHhkERlUTk
PYe1dPLEGr39OY9ahfq/fJqJc7erB8FFXm7ar8meVO5RvJ9CDI7pB0yw5/yMEuzk
uVrtM+DhD8p2Ajc86ZCQCJyZV17sVSfv4CYC1ReB9LfmR5ilPZ/OAI/kqq7sI5Xg
q0v5LXZkryrb9E+oeyABKvg3EiNzJXjJoSYX89l17hXq6XYrM6BXYFs2dNxbic9p
KiUWGXVTzeItvYBX9QxWbsIc7k+fj6bUO1ibo9cRsRmLT/0+dD71jmsxn0wJACo7
JW8y0eKeJS74DF7fCmGfje+d4mjUVuLrc3zKnprSyFQ2hcF0sQvvh/DTwi7+eNws
7VRskUE30zWGBWwLsvRqSbJxXuglzkIspw4h9Re+npfhWLlStq9fvLxb7w8uWo/F
+QCMjSCEBBKM2KthcfIxPVIpWENnGSmvtvzWm9PaKPRaU25kLbO5MQzQeMHjWzRh
ydQTvCuUOVyZoktqkqPmYwKHc4kbSEGG+oujhcC1hVY8qSOzJy60hoG919AvWJ+r
Xoyg5tX5TSD7FExHf4cp+UBw2kq/FRoyjAmoqNmDzSaelfcOIE9LNEm8Ah+m2Qg2
mMxup2bIWn6sK5YlppmG7J3Y1dO06t9PL/no0tC6eT/oD4m2Um/C7lVPR/iDdbFX
O0UyJry6cMrVwG3TN/HJbKWniCckak+pdxX3b5Oalgau1c7U0RUn/5immh+QG3Qh
ALBmQjAuw6sZiXlh2vkuGrq6UFSLweSee0gwtbRFh964g497uFKgzNugNWI9luZO
jGAfJYG6P5S5lrXKb8fBS4wwFrfLbdTIZqRTS9rKIat1MYX+c8wP/qQngk+6LQVY
ll1AkLf6YnrPt2S5OLYWYpuG1ARGya4N4pW5XpuvABOAg/0OHcoh70zDSPHer0uS
g7dhKj0c3S6JOQv/jWJeQwTv43YJG60WiP8Z5UP8/AaDb7AjMK9AZ/n5FNuI+QG3
YYwDIVeghjuVKJVF3/A6EST4U9GTLfOptGBGyVJ5GJJLApBEjXeXOOse6yCmo1M2
bYmg/ckCM+YvelMksgIJntc0vdANPsbxFx/jFGV7BfkNNr8olml75OTgusgAGeDl
5FAYDix7aksibxy1wR3WbisEZwyx5UZf7Dg9AAVFBYqfGVLEJRCVcnnIfX4WAI7e
Vb0KylllTWSA3aJD9msAUWgQPwMvd8unZGqPSCSm0wrN4XaRSyv+ckjabUMLJnVb
t0vNuQMY3RPkWhyIN//dwp5s0DSvXP1OzXcqqjEls6v6VLSoJIZXsWo2uKu3lJKQ
ax0t24T4q7CHJKuzkHIEL8UTeF3QuCfX7uXs9++48IdHpqBWqzPexFk96pu6bgYs
qIj5MLcRiDGYgBTLS4zLZonMLRdpS41cB1G8OgciY5RwhyuP0OgTi2NYx1opBJ76
CFoBcuj2YmnbcSAuX+e7IKZ6X84OcU49zJCxnQWNwDwYS3g2dttorE1OO4ibCmjb
+q8jEuathPw/WcglB++GXM9lON+uzYmENQGT8flNmizJ7450xlM5WEEX4TLsw0lu
xTw5x0lWiZb5hRopghdX/KnlqrfLVNneIOAWrnkA//lFj3GUcXtJotJUiBfMqUdg
C90en/mQeoxtYTuYlRO40RkcbcqCmf43oTXV1aAxthCqadKsigrcF2oJgGFj9ydt
aEf9xwfUEUo64TY/bR9PSuB1Ucy53h5eiC+7GHPj9LdvSe9m7Kdeh3+Os3veGHRr
P8Inx0+XAyVb6TWvTV3XAoXc2drwTJRvq+ZY2iVhBJndBqt0s2oeLwAqtLCBdKWd
FnXpY2vJNPoZLVF2GJsQZGkUJqj/3O3RIEOhSk9maWnu2ikNP7oCqnPW5tzzsIff
h9W9+D8Xa9oeaYilmZ+u98IdXAeGs6L8CHFpNIzNVsn6VIaGKb+e3KJopWeSa1Zj
27PHpKKNB5GBE9EJcl7WzPKPNq5Tf8e3+jiNQdTjP/2cUJ38Eo/H0gkgwqGNfSbT
W1hSonqPEPr523jPLxSdnAazW+qPgblTiuWmKNwZj4C1kRKSLToc2F35Cevlu5G7
5ykOEMA7taxoiNIiIyDob9m85ZO/j/z4oPkIjHxU5Wi7aYey4bENzv5+muuuFsrY
72jy6AtkrvT4BGTIbgSxXcajnUZeVohmyRxlZ+DIbTQ2WXQDa9yMvI4kbIMqZ93b
cVW8cLR7OQnLeru2O3CQZ1vyw5llJ8AVt+qknPRibOX5hZYBRZnNSBv7R/z7xXt0
bQi8UyO31BuobAMPREENuaumoCKQhFHRP+/uy3idBEUoKHAmjrv0XI8MrfuqBdku
qdDDA0+zQbGm1YQ07wv2lrmALe0AUrlalUfSeCl9Vis84cK20LYB75b9aX6/8xt0
5DKbwL1JuHkw/0nD8oGWGMyOhl51k3ULjEhoIcvsTiDsNB4/ldfCmhap/BQqZLkw
81ZyxnLNqiAfr99yy640qTlbIbKRV3wNyyn5wAfQrdq826oHfH7YSEnaivlkIeDa
O8Ck57phmiwY1gsR8YO6qEoy5FG32af91fqUNUpm5R4OSj1G9pFkb1oYcne3T/YX
9ZjFwzw8gY4o7p9vCDJhSz0LmkpSEm+oRBaZ7kw3Kscb2/OQGjokz+rczk6ojMvQ
CfjbKKI034KMLFhZN20fHQfDbfczi+5rSPdQE/h+0Sxzhy1wD+AbqOpOt8mimbMn
qiCc4ghfnBeJLU8IHYaW3l2X3K0mYXKr5k4degJNkzZny/8/QhmubdfrQaZ5Q8IV
cI9gcsy7jvfMropGoJREHzfHTyVHk+0CWnAJmHLYyF6BS6A4vQ2c0MEOJngMjju/
9BpBCIQgJUXgng+vu8+ni4I2q8vbaZNAxBaYs2wTvMl6HLp3r2cOk2k91xKJqm6I
KjraxtplKYj/4HqZaK9q5u6lsYlTMNoaOvY2kQ3a1o6EunyURGOHwh42aDAvVucw
shAvE/n8wa9zr/iw/mnPRMwhCd4txuYxNU+O9Z5plIOdkOwNJ1H5vey3k9mje8z/
C5Ef6oZHaSfM3gdgqKe7Ikr+WFmDFj2YKD17gkqzqddPyDJCsJadeDSda+FMyum8
PMPLvKeBIBQeBNxnGNu/h+Bu8sBAMkbUuYWg8ugm5F1vTadipIE/aiaW0nQ/J4zU
m35ZAhuGKS6UPm7UZbL1mSF38MuzX6tE548arJlujzgRz6uYLxOJCb77O7bZl5/x
du2xIPXzHrEyH7JwnVU8YuTDnmfcF5wv3YpaeCAC4/Z/E9XWJQuKmCnGbprWLyAJ
7p7KGNAGiL7OFYw9MtdQupWtFiIUDi+cOQ/WCIJdY9+06JqHhZiYnhyEtPzMK9jk
SQ47hiv0AgFia4M+RAJQA9qCS2ep/uA0YmPIbd3FHXZZbIphG3z+6MIAnyV1Kgbw
TNL/CPNcRxzKTURIRCIixwi3rMp4kcBTtjJgP1YP1Ztkjf+TM0/6qg5KT41VrVeJ
dzCCItYcAl33k1Tc3Tzy0l2IGH5Jic8B96II6YBMJ8A+2IbInuvWMFtamkS1aDQJ
2WOHbA7WVe1qAOrbJ7dbkhi/zdFbDnz6GcAaDf3PvyT/EIdEhEVrGC7rNFOcfAsH
tTHPRDOfgKnhznf5LUPfTWIeeoS5x1WZdNdH2A/48TfCunK2qrIS/kF8VbULCuKa
VQKjbE8pm9sHAVfDbqqydKtXFZW932U/mKl9Ye+MaVLzs5orQOAOwKY1w9B9gvWj
q60lmSpupoaLBP9B7jffkG42uZL7UaUDSLCPf4205GN6MyMDyuND0uKEiyf4SKip
MtLBQCH/muB/Fg8z7knXZXMFk7vRQAA2+z9tCsAPYRFNrcLXXwHM7a3wZI9qHPh/
18B4FcaCQ2JSAWNsdbtPlnb+JN+4DvF3YzlczmiwWnBbSd8fO9JvSgbaM+uIa7s3
rXhN5zZ7PMWnTwaJph/+UUQJVH0VzV4MfK1Z05dI+TqCej050xPPdAiPMkcwufaq
hda4n7y0SCIk8qazJJ3UMy4nhWpeC7Be43ui8IKu33RVAcSrJK9BuwZWYh4pPtHa
zAcJJNpoR3cVeHYbowFF4zokSun3hqcSvuzaUGA+ngzJVFqcrCrZFoSY+z0+a6pX
ZoWluAI+w1HYaOFkUTvPN92CEyRy1Uc1+nQS0z9X7V5RjEhYze23HfHBhIUaZNMZ
BnIWBUX5WIsaDb3I33Q1Ikdbsx9GZf6Wg2K3Y1gfALaJHNiDIK0179Ta/YTXvqS8
1zCBOOi09ZCJkqNrytKQJV1zLBWtdA9Z+1fuNYN1pF5dTNrAleg1vrT4w84a6roy
EKi1fQ25mrQwcFCbWk4OeS2j5+at0yqHd+0SzGBumJkSSWYfuFA6ShT943ptuNpo
ePB/Lm9PPEQDJHlgtfRldXAoYm51o9mf8peyewot8Vk03FbDJoCsFPXkk1dBC8h3
fTnJjKZLhxOlewMRiaW8x+kskL6/s2K2OKkyVn2Ajy3+GR7mdGjbHEjEl/nf8XR4
L01d45+CrV6h63FOaVSbH/SyxWBWiGiJUF96i+eMFgYv8WPN3exe7fiZEZQyPn0L
Wye0zTA75v9i8tENBPMzgd15qeWlhSNvyYaBdBGhwwAsgkCyI7K/c6IyqdUBjlYa
55PLP/7E3zxGktzVxs6QgNgCyXB88zaXzJ8Pad+/iNXMFYv3ymswMUqEYthtCKf7
K0aaUFmS1/jmBafZr/iQI7O7b0KYABocw6uwkKKCsUEEFHdwtQ0V6CDgPMDUKvZQ
NbIwO3OdqZIzooi9FDSjQvJQ6bEw46rwwYJSnJ8CB8hOXX/u5Vwt4weJmJh9y3Fj
IIalijm+PncsIQKZcDa37y31WcRYZcZbEWMYlC76Mvn1n7qUzcbF0x7Sy+dB6iqw
cH4ZohEQPFSpPMhWbVzWKEH/cFQxgEcgjgXJCZ58Sx7nXR6sKV5SuyAhKs3QEKbm
al2NPcaalU5QgvaE6hYI+y65D57TDSq1CDZsYfm7SPuL/u0/Krk0zQfLn4bbNvyi
/uoqSmHweZpARrVy9IxjbsC6QFpVBjRj7KhpEM3YZruzwmudC5Vmvqr82tjK2972
gf2AtjZ2x4onahjAlf1AsBAyc76wmcXbXmKuoNn5NoqXWnh6CVz2mMeEGSdB6GhR
zpBDOmkI87zCZu2n5yiJkYoTbc+Qj2rK1yNs6kbTG7K4L3RuBz/lbvQfcFcwVqvR
BC9UWvL8D2o/4VHty6P3CjP3hw8tHgFOVDLzkblWHUAb2wwYYkyk5Ky1zgxNAIPu
JdyIgcR56ZpWezZc4rCseZKWXRFtpQWcwkBRla716C62cP04FH6AQkg7Yt3dk14l
9vh8NZezz3KjAzh33spjPfquBKw2a3u2sYk0bpGbdM9UvcnX9+kYTS1orZnZ1z0X
mdGGRcSUTRoTE2U3YlZChxgBVfq3rtjHIxzhCAHKXSWTb6UmVbyhWtiHh3S4mz8o
F+nApPdt6A3rfkk6rUEFdH8kmrDBjI5Mm3w15SN5l6jB6W1T7EKBXvZqC7tQA45h
On2WA1AVVUZN+CdDcXJe9N//mze7Qn7FXl8fFgqcnqorghQTGqSCglAboeZbYXwf
SmJvyyvlvYAujtSap2t07ylUwzokq5F8HtJkwHn7/1Ko896aLW33H//W4IGfJ07H
8V69ZTmF+8DawcPCrpiOrSEnZcFTjUCnEu1qL58L0LQnJSQBcU0Lh7ufR7F19+/j
dzF2xZlBvRPQEIgzaUSrhEHB4O/MinEVigAWk09B0vy8XQnG/1mF4JYOPKf7sZko
XsH0mTar+qbBa+m+Rtj87Q==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
kfjERdY7SSJfUdzRP5FP2lRfWFInse8WH1Cf+31PBF8HGD+92AMsI8/TwTQuXcK9
iuezSR7GbrjIbNr3QTk43WJXRFOac1JNdzo5QzZLSL+qXA3htvYVff1czQ0iT64g
iaa57eAXE3veABlKcNOruZEuwQq3iIWM3gTjLjG3PgbXX0YjL1DGBIXWzDKXCrOU
+2GrOij4H99XyAoQM1anUW/xz08PvmAQv5D6ntf3r/87eycdWOc5K0+hGz6YkS/k
gbWL69eCimUsGGEi8nFg4mrE0FNA14EhFLSs5b4SZg9R5ShMfGJ35OaNw3RSl1a0
vNVuFibud/Cv77LK6e3PCA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 23728 )
`pragma protect data_block
xYwARSt03x1OCsBBm/Tjr4Zqe1Y6n3EEghREmKdjG4//bKdaNxl7nfU/HnhXLhXA
u+BalDT4IflQfcfU0pfvZGvhrGMAjcVZVj+OBa0a4gMW6VBT/PZoG39YDNwAyNYE
FdVyc7P3FqaqeCX0CMceP/i/H1dPpkTjkLA6QF1vCwZitZdMrlRUsWrFGtbyDLZt
0HGdjaeN6r2t04DDuajp0vTc6i7ElvtCNmpzxTNMXsz7OvZAXBRd8WZN4LqPre1f
BrpRLOrGHaabqtaFP1YGrLNYnQTdh79S0HvkupvgHEQHkFLvTuQKFfIB9tt4WzeK
2Wcne6pu4S4Raxl9OFja2KvXIvARA/pYuzYW5WGMO+e3njVtF6zPXblS4X/oBgzp
/PTO7MN0N/bb+hb20lISBIdDx8y4JttAp6ggcA+ZtXj1MKMcx7u4ymAC3SIDP6GD
WRqH7G53fytQM7LbSBhT/Gk3yDBAhKN9bED2YhuYpIKcQ7y6sf75rM4tJrONgnmj
jjACNt3cgwF2Zm6M0RTqV4uv4IwtsjlaNxPsiNpH0HOT42IyCXfufjG6yb0O/Qkm
ngK3/gaVwA6QdFEdsBaulbMw2r0ODIerdVifoQssU11i4idlHnL6qeb6tUReK7r1
EiJvL0g9bEcRwSRAFl2exgD6X3Qqo0dBsW+0zaxbnLUz7D6IUDdOI0qwpHLLJgJ9
uw6c1ZbeiFKjszmr/OVyRUCp2gELugHDDrQkkJ035WjClh9pUH6Es1Q6vDio+9x3
4LWWKjKtbOhsg5B4VVlgeWz93/VE4/IfHatjeHtHYdKqyl8TzqG/tGahXWfrEdWq
tLS2IJx4dZdbVfSUve0T2u5s/qsZViGi1erk5OtBF0trxGbrYEtNhXuyCo4YHraV
ZHdcdw483SZvgLfO5G27QrovndGSjV6XgMYLRU7r2+1r74xjnkUTKp3s4YEJ7qiH
nTfRPXCz8rON3bqbAFOlSDlFtt7r2+tTbkAABnNt0AaVHS8c/6U6jDNvFZz+nOcP
xRK3TSh21QzgK1V5xc6PAVZe/LceOHO1cwwZdig7hN0QQPE6DKisLVSXnUfL6d2A
eOFPFlB7cZ1wR/baTpSy7dxojeBXaETObNFOkxmiP/C2s2OGG5MQfpSRwp+jpF8l
uwXZ/Eb0oQIPf2PNBsN8hYWBXdmX0g2GSWZdyXJRRSTwP4UHUDoEl9ahZSv3fz33
OqZWvXW4j9kEJHjISLk5K+ivaeGbF7xy3HZlG4gKA7M3C99dKweJITq9MJaQcGkl
bm1CjJWEo9rwRbixmXJBJCgynj9X+BGORydW+XsO7ObgIM7veDgYljir2gfzFLvr
dPhQdz0C2+l0BtPxZ71wOyxH7iHUjLJQjilLXtb76+U/zaxAaRp0Q3YqOQhT09Sp
JstPmw0gza1gDHWRdc72d+2cHS8Wa3zAyI0sl6vVmkVWvYXE5uQJuBEaIw4Nu7Dt
y2c+Hil2p0OlGUlEDnY04DOqJfQHIr2xdau91XJpxzPbxAaOagdFGfhR5ywnn7sG
BH6Ja0dR05nOSkVrzS/G7cEg8vr35y20ZuBx4S0mXlXdC3wluCZ0y4kGOo3ArETY
+b1biwOOgLlBU7miqUHXjT5Rx4QbSNDV8fJMcQb8JMlgda2VCs9r/BAW3reJ49ch
9K1UitOPZfxFX4HscPH0gsk1bXDion8WXF5wcRyORZAJIgA7TokGYqL/mpS+pNob
sT2iStvTVPCquGOdYj5DshTM219d8b73g2FbZZmVdtjosPKSjCCG57j2CJsPY8Gb
TrEHJ9goaKaLoP0NWqFHmNnXkju/SBzJN/qeAs97p3lkYyrmtGro+V4AsQs9mU0b
T0ACJ4Q3c6iJvtIYTOS8SrlYmlkdNVLYH1l0veZQeSvFuDwf+euRLlYBy7FcLQSM
uOgGQf8XldaAfIdb5Bmqr7U5ezd9gO9M0FqUWWrKuxfgPSIgLcxLuuS3XUVuJhLb
FkNnR1Ksm3iN+bfhaVAQlo6vQJA8I0XqdAutESxdg8bOPtXii0RJvxx98xEuwsgi
H2jNxiPcTKyW9p9Ds2zZrwofksrEJXr6AwGl46yUJ/iKMMS1eNM1wOWt3cH+v3yW
IjMenPLxZxXiYMnfd/RHp7g+XBtQCxgYyY9PY2tla0Niffgm5snSlQznIIkeM+f3
1/PldiZZ73/FI5cCB4gnMx2/3lvv5AorI/yvBF0GHr2qWxb9vOE+CFpz3YBTUCxc
QN31VTuFAkHoy7FwgdiIZX4lr8SW+oOuxguwVsH0APmgojFTDJ5BUGbxpxYDIXX3
r8j3jMtv+7eNONaYGDC3X7R6QUQcQOXnJLUUoc15CHoq+y99QGBERfA4/L5+V+vR
ACdk0atezG2Yy6IWesQH1dfGa61M5hpZQC4ekaTpvJt8xk2QPzMxF/ncNCtp0E7r
JLR0ifnKxfr3gSzY+TjK7UgASsSvL+khc3htFGxA4aAhdcgjN/rb7eo5YGRZDenO
vD9o7433fCmmepL2LHEYJvVDftDOt7qmQWpfj7X1XInW5O6b1IEy6zAPvPm254vm
Qya+NgpClv/r6H4NnceLVBv0lpdJKlXRU53eZ903b/xSct/K16POsrffoZpBIhlq
iGLHa8JHvuaOlaHcBphLGv8zY9B6fzkKoZf76XARhjw3DKAz684h7Sl3z2PDw178
ypPtMO6viFUsY49Wi6MMWwDIrGzeQccqwRacXmpT8OXkWJLmw4AHgFZjOGHER702
7pHH99h8FOMxNw4YQmPgRHkG5XT718oBLxO2ik3Qcout6KfRLa7cq5eObnmnHhaf
zLiBY73pd8rJZoiETNfujBjOzkFLNBRkZ5LTJvtgyMDekoHxkzfRX9Yx0KyFDy3f
EtuhdZaNqlnIvQnMbme7LRPQOUJZcTv6CrxLUMf+GYYbMa4+jSSgncm+CafdaRSh
oSVicS3kmIFYgdJbt5ccQOK8crOTUAumMTNRxhJQnpiNyMtKeYLUPkaHda5Q+Uax
TW4v2shopwYKxNDCn/4sk8O6CgQ+x1GQae1fGtnGjrw1cu/dqMMEnP0H+oeYc2qs
qtzRDY0hbZXjEhBxi6isn5+yWcpBqw/EyCkaKO1SnDAwbbFxQm4vnNbW5PIvlg9s
evQDHxy91eXGYByYlN0yzAWxnhU3zU5U65NfHu4L+Zk4eqad5+JshNFg66S4Fdk3
+E1LbuMZpmkYWaAUBMls1vEUTqjPr7Y3TPskwTkVSoXvJKX7vxsQhfw3SqWTGPh5
ZKSogGLP1hHPSqmBiW14mFMIdzy9Ss80f7Z6fIRvr871wB0lWHUbDqwUTOk97jdd
xBZCUoEz3KbY1n7sAIo9bXWObfUPFU/+KKhk1B9D8xS7nrTnLzQ24PFHCz1Vmxwu
BvF73IPGYflTMUS4AZxSkMutppUD/04ddg9Og/EXjez3e44HqlOCJYxXlM5vafpX
yJukdW3MnYilF+xg/bPucPMXj+9ed0JzYpnQGiEczehgzgn9DUwSN0lQgd4WwR33
fYdLQtryq+O2vAKuVxMFF8GbCh5vRBBo7qD+lmRASHpiaTnbQP+Wl+HIVjJ4nMD2
HiHvszfqHhS867Vzb8MU372uc8XmiHsAzjfjhmiUamB8dwRJ73nf7MA0UVJFVk1H
uiFRhvnrlWvx72fSPqf76hDPygPyMyH0Miyu99OvwicOmWnZ4kRIIn1HpxoIuPXr
wlVabr46xtW8rjkdtzLNngKz1XSEMGbbl01LWxqeTN3BEhQ5QxwGoxBLrlxLQ8rq
cNSomOX24vCjf2Efe0qQglUGfgn4reQHKEGqk/y9C6jT+zc6yPKl39kQKIFHklz5
cIIJ8dJQVC6buAl1S6Vxtxn0rfQcWoU4J/iKRGVef/tPgIZdXsxDJabiDlOYFLpu
chSqZO3XlNYgk8IpUR1tLvhv6FJrk/ks5VZnJAEIYMIF/p+tTaHUi9CwTnNozEtn
ZmScMi2cHt7iKi3akM/YszFrG7/xYvlJId1N2W3rGcbz0uhxALghGCGQLwZtLQ3y
T5J49cULXZBDwtc5ipqfmxUkpxdzJXhnpjmrjz87MrPtuJZ0JOeypTackg7BcTv8
rBIhZAstP3hOfeg7FyOpUT/j3OVvR2jiKfjASu5SyYhD61sGb48NBNjv72vzeX6j
wAV+EqivXiV9oYDwxCERsHTs6oJ5j1B5ep/tmz3wKIDs1WnKE/UTtfDQB3Utyjv8
iK1u2P50B4KzN9Nic+xJEJxEx5uVz1rXKH/Mvvj2l8tyLEGIqZoFWDLNkIRC7zPf
RVAH74OLZZoaD5LswCRsS0r2iLwr0vYYngeN3JtAQ40TL/ulwBEKRzDtWpBjth18
EndgHMq9PPNx/HdWDystOobCvXDDkVrlgpD4ZKrtbtY8l4GIYDQlw9r7blyxpXrr
TTlC+BJheivA3aoVwLF814KphZqfMyV2JBvvqSmtnIeEOQ2WEHfZKZ2BZ7ISzjKP
QkYTY/ZSkmUkxRxpxl6ptbJIEdCyFP29/q+dOwymwrXyXLNrMuKEnhXhBnarLBC1
LvEsJ5SQ+tlurRY5rCpd5D0a7VabJW85wWKo42pwkLOc2Rg0NFDKUP1pNL0FGwyo
8N3AWzuW3eRHJnR8rzxaQbkkMW61ZBycOOE6+7+KIO/TqMejEQdIRJ1zUuY+y4+l
I9L+3QMWpVkuAgs85CNiUTxFeUuoCVt57zOe/Lf4YE7dMMuncqrYOgZ5Yxk8Lf+c
AytBfkDpOO9lLnfE4DDf/DFC55d/t1Ptcw5I3ClmgpmCyV3heMk9sqq1BcOYpspN
J9ztHJw7wLD10ntsFusfxjoXkdrFZ/4T2a/TDPxWJjonSJubBls72S7/fC5H4XHj
8wbDvSH03VV9Zdwh4EYdjbLX7g8pYryDil5PW4z6zKltREDQlIzMLIpwLrpUZQ7Z
81FCX5tUUQ0p3Xp8Nm2vpY3SWt/4F7O1A2TvAo77wsqYlf9c5kx2weJRqhCHCifF
5dxl+jEzuUPX3uOMGFCNup9U2ZLjkkF/B7kN5hR6Ye0GfGAxsTqJzKGNls29LTQw
B8+cTzJsyjzOdV56h4ckHHWalgco36VZAX6FxM/r9Yozz1CdAXjlBKcCKAG1nuqO
4rh5Pwsuz8ClRsvO3eaLMPqtXIJDE7bxJ9b7qDkVuHXrI3SoTjuqCZa8R01CfLKW
nJ46TFaFyPo+kcneC1aQuoGibMS47MyjFmXMDt3V5XiD4RQYBmGoPCVA8HTavRKt
O4/q++LcV+NPsVLItXWhzZQNRgZ4OqhIsFdSEkhat35/fcSTImAgY5pdQSWzmBsW
JGuXylbyPWfgfvKAEPNvFNMAwMgCI5GooozkDBMHDbut1tJvoFdU+K1ymfBw9jae
oB4gGf13QJ4H2AvYjxtsF06BmATr3yx3xPN8LhbMhOFQjHfA8ksM6GjIA8eFIwf0
vUWafW3DqrYt9mH5+dmblw2Zuvj2Vi9KYp35vuu3mkl4ldZGvzIIdQRKsWOdgUDz
lJLYwfCTRpg2dz98frbQtYtL3zOq94LDJ5AB+SKk5NBz4X+4euGp+Tm1l38wyxCn
WkllMwO3UUlO1+KIvXrVUqu/Z7tcKi6Ib+96jBm9f73jCu4BUBXDLWBVsxB62gW4
5T+TQobQFM7I6Bs2FKdjH/L9tRSyqYwp/IriJVgHkf266kVCoTAKKgun+MkWQbP0
VSDrplbyJ0heW65KNHVIs4DWVeW9st8tXitwm9QmH7AUk9k1RX9ooMSiSkKBV1jR
ppNDW9jPejv7iFiqUB1Pcz5AWbi+YRVKe5VO19ufgVq+f2qYEYvGTLzlfqDffHo5
Lr8U/2EaxjZosBooq49XlaSlT1C+MScSuv5Z2clgn23rxyYEwJBlUzVYyyHsstJA
mUCt1xeoR15Rehl0rIYYNOWXwD1hNxFn/EnvzNAWcYRZ+03H6flhok4siDEmyfkK
QVM1O8FVXuf2gcPN1cy+glMGf4qa7zFje9Pi/sSvwX/Ep+/7gFiacZb02GrvVKp1
LKiyoLsMo4ot8vRNkLZSpfCPOEhkxPgQ3nrijWloZjCTbo97yvS4Z6mq3p1945fP
kiMrgmGN8NyG+1OKUvN06NNbWGPnr6Cf8WT0k7BmxabPIrfo/2Bz4BXW+N4rSMzX
di63B8HtqCCZC4Osp2LRbWoRnZlsym5OvddfxJ60pOYBY2jecsUoLdOMgGbkFSHf
VN6a6ffqVrm8Iz6tZs/yobS1Q9MhLVoXqjVKuH1TH9PAQiRzH6wOiJ5Hc3VTUosE
R5aZBe3P/HIdALPJitL5mSGlIE3PYeiVbE63N/M1wBa/4dnS9AvgC+W8/JhP1mTE
KeqMl+qWtXduiT93le0d7Tyaio9WPKneKX0dZRwqIcZfpqaZA71aUDCkWWj544MR
GVvrkiKvthpr11DANY/VUklmHm2s//QwNf8d4xlZesNBF63hapZ73vOg0NEE5hew
xHuiIGs3xu/QY98CGs91kngfFerBBul7aQiQo7pGkXtth51gsVaiYKTUmWRekF3m
z9kcSueLbp0225FZfIUr9sntcxU+n9fzwwhoxhZovnigmhDehITfL+mUDO+uBtHu
QLCZ/mLU9O17tC+11A0PTKFygA6o/Q1P7eOljvEWrKkabXdq3FnMXmoN03WzwR3R
9Y5DlUdj9eX5YXGRpN3rvU6H2N4BF5HHzh7FzdokF86zNYhaYy4ptr2pOReNVifL
op7mT8rL9StvcMOinMaJkV7sJIgDz+1ryOYNEJMQGJic8XsbW+t5F0e+OxOnp13V
UC3a3XC559P4tWIJ7MC1K0s8h9LHiX3Hlne10IAyQHBIKVn8fotBKm01ZGmQ8yIR
pe0o8brS//HTI3JPuudSr/wYKIF6XhUuLZE9eBmaaa+Lj90rQLAbdwcO/lUnUc25
YicPRDsa12ZlABAWYIAh2z5W4CCdHyJgCNtpA1kPFVXggDxOdgm4T+b9IJpTN1mA
Jr+44cIMeZiY6clZzB3KjVywwNbhqppe9EEB3Opj5BEIaEADM2pUKGM4CWoamD+p
qvSYeAfBplmY5fmouc2lX64FIWIP61L3mM88pCmI8RPNpTwe0LNjPogPkRv1saF8
5RxNaZm6y06rUASvMZYDcnX1JhkxtGXyL8xNTGFywfal7Q1a/JNYbU1ezt4nw4eX
O6N8jVsmnUYWr0pujujSZIFtIfjRPzkLrNkQ6W/gsZL8sDGVGFIo28fG/Btbu6vx
yliK0YoxolTmBMGu+jcQQHZSeaVhEHlBN3KnTdJzZF6McoGzuaUuueJKvKKPqTsQ
CF4WaawwGA/cYkQ+G2dsZ5i22YO3vVkniSmNIsspfJSgTL3qQtGIPMRcJhuABNyJ
YEhx6P5zA35kXy65prAW8rqk5NWZnaNzkn88a9NL9PCSJF2GUv8POfc+jl0vcVpY
pgWm3HhVR1dwRq8BACtmpPAvLcNlUZ1a3snjWUyHzndRPS0Uaj9DMrHXHqKI9mhq
eYoN9+QKhMEfcvP89WUEd5ghjI1o33e2iVxZnLZt+0pM+kiUB7QTqu+tOlKeubjp
4gvrKvZHHVjfu93qI+TOJbZcwGXtaYhYmRfLMV+4zRb6nGz78mYmZWdjYqsABzX7
znHjBGA+fw2qfKfIHi9WAJtVLQ8Q+W7PRnkXRDBUso4uPj+yu3wxpshgL3WT0PwM
m9M3BzjrQclvhCwsjqWbK5XSmKxGrqFGwG3aOEihs3g7rFq6UtiyneNmbNbHzyss
Qz5lzHr5+6CrC9xqcO0NMSi8lqu9D5+LTxokkTQhDofqDCyqA6FYQiggFaG3JhAF
7UaLStFaboc1rJxQCoipajwJJsWwZmd7SJKp7SN9sC1kfPTJtC0ePI5nSCg4Lkyc
MUq49c0dVg6jxtR58YPsriTiJkZ/QkL7E2+t20cZBqf2P0HdzH5aINroydsvQlVC
08Dg8R/ySx/SyBzqNxDSXw9sV143zxcvq1GfngkXC3HW9IFyifXHEUj+Rfz0h5WU
5TdAyOfg2NQU4UTXIlzv3KgnTn4ywVE8uXzmPzsvHqQvhbpjws62B/QX1e8Ze8Pg
rpTh5A2tGj2MdeuPgnqAzvjVlz5XXJ86eznqm6q+LERf7JOO/BrP8ezdYUgaJF87
aJTh+BW1M4ZV7RPifj9AM7RKQOuw+KcKOQtgspZqH6ZQb8aAnNDBB2W1DVew4l3W
rJTA25AzUNHnziTEm3f/iZ2UKZe6X5pb0Yf8OIqjqoiu2eo4aKDoPodD92sGHYfr
SzUbxEu1lC9mNNy7KPMnenVCAT5avt2RwHAIRbYDX5NzpylZAOl1fTsalO72A+4l
hmBfX8CqxQPF7QpQ+cGwDDB5G+s194/7oepH3HPFM6u5rd2QGkl3nAXKKkvFCy11
CUWWvao5OuR5UHGKZtGDCxQyzczSNGwQKjUpQvDDCykbcRSIzQkz0/gov4pZr1K2
bpZtFwCZx4xVRLqEc0UzqL4JflYIWS/ndso3e3bYIEavwSJUchaL2QWYZTBPWWTn
Y7JuNFRFwgTUlnk6H3ueKPY5WBtKlJ2TslsMmb2iT2TY5hG3Mgh4B6ULKsGr3Qs5
yZna/SfwwTrDb3eP99IPC1Q+4d6qo+9+7/nyfL4BKMR70rSAo8s/YSVRmfqj9X0+
PnS47pjRTMFmPLP6VCn8pReZaJSo/2c9h3i53ma7dU4zAUVJWSd3TAcpHaDRusof
2CT+b4PX1saSjPBcmX3+FYWScYOW+IwzYkZkKIRtMHzyM62ftf5U48kKlaMCkS+y
4Ik2SrOJ4+MfWF09ICl07zNMNHfT+lAPzAmfipPx5BwIz32E3yH2+Ll0NP5zW9TM
o+QCMKjscNN2/aFuLnny9PT59y4P6w+TSWU58y5s8rpY16SSAVcoIJmiEkZAEQDl
GxbAPYjf6BccBnDYyv/jyrHGh4hbs5rTo/wts5Dwr8FjtCZtB947iD01pxSWfSPh
zSTeZXama89k+vQ7f79iNAhDlzRpDkj7TJZvDSmIwzQPHk5oPNUKf71mDvqN4AQ/
pIBkZXAqy3DsWzX87ygYgqa4KZtOpbYL5dy4nOOI8oUKqIX26tuflfxxlv9862az
4fHh6I4TLxazZAvMn2S0TW7AiZgogVqZnIMjbEDarzvtNq9nWlJ1Cpg686NSZcFx
aMCHxxcglpJ4ZMj9Gdm5ZEzd1fCk5IIOi4lShKLtUKwdIO/RIpTHaK5lFPoIBhSb
io5ay1iMXNudP1Hm9+qMBKwbonDXDenNC67Bp0ZtXImNlJ3UXeZs+i/227CJcqz7
RPNXeIF6TeYYho1uwg1I7By+1CFWTKdYye8vqK9AfAAmJa1srn8XyYnYCbMJeMDj
leJi8XBwVqHZQQOi/3IcwMYlpVIuz8bM4pwDrbbHCKrm5A6I4j1aFwTaySsmN8WZ
4aFoJPFik8CpqtHhj1Qnv67BkY2yiatEazd0/ThWfWyOF35CebJ2pFS0zdmjUw1H
aHxzOeUeOPvdz9ntvKq+kh/Rxl4ZXGTQ4RZVN7qAswMxkIX32DamSKit7cOChboE
s5ePS4ozsAFepiguQeC/+yrs50X/xvuaSsj4WDQ786dR3fbfeChXscAo6ruJcJPH
9JrTdwohDWet1nSdk1i4EraKn3OY7u/xZKhsluVpBuqvjayRkYysYOoMK2TyNrEZ
wREgyJ1fgwsjz4ekZ9u9p/4Tu54qTebg5UaxDrMR6fr3WXMsH3qF7AMdBaYYB9fR
bhIZjmy9Tn833jJrUzdAqLBPSLKW76FQhF3RmS9IHhedlcIOwQsusp/4fIjFXkGT
ZFZ79Rlgmz/qP48XEEjjkobT5P2vzniSJFD0ljzW0/yrTdZKti8+T4dGbqC/mxvZ
w37Ak39KxVSIg313J+qyR5n3r97abbhYQtEtZLeJqmrX+dyH1k5+/rPJh2QsoZ5c
3r4aJV0pRKDv8ZOumBabNYK5kyDNyj1JVg7iiIhq6u0h/o1QiH5w3tCBs5TJDYyC
Os8/pufH+p1YvI7psIDc5Ir2bjY6BsFiviexUNwzvg3bG+SSgmv45zjuLSYFafDQ
diw27khWLIIgIyYuBqxhRIVeN+7ybtgU4rqnSWd6AgzjHJEeLmAGnsV/80s9/mhQ
sQHrrAGgs9I3GEs0omOfpQNGlZSU6HX0IkXUVUq8A4RWaaiJvTDRBmOFEFW8yKUw
tion8llsnRoi8yjyi+OOPOdzq7uo7s1b9ag9P6KsPEm+fYBj/r+oUQjiuFCAiCSG
mh5M1fPMGUd9QyTTbspnDRLzidgigyIwlHN0itJuczgcskTFhU7ar8hTu2foOt8P
vwRhGlW3pLreQ9zqStJ0fgM95bXij6o8mUo/m7BlZLvntHGKJiV1g4Dgq3fe+KRh
RiHsAuci0GdNXoByebeGMxEpeGXOYHh78xxNMWMewDMNeNaidP2Pmlk8IaiQjF4L
dV4QupO6yskkoZWC+HX68KATs+fLOlUdkuMLnZzZ9kVn7Vn3G5eD2PrxpqF5x5aI
Ge8eigXn89Q5NK92dUCenFE0k2VMfh8LWW53HSe6x4GEKfxYkdYa1ADEb704oJit
g6CmVULIEFkUz4oRSW0LstLw/5nenMlv/EIu/8qCbhx+I+Y143T6p55S1ynz3EE/
9+DtOKi8Ykqioxf8f8u47DvO859NTPh2A8iR29wdmkpxmUFwM00o/uakaQKFoo02
oOpP0LRURCbl+1Husl59edTHHm/0ap8d5Gcr5PlrynZPB1thkxChunkViagDWW4u
eh3Ad9fK6JmrMTRr9MdPyUUgs2m4YB6YBWFUnLYksNb7TmV6UqorUMpdx5otwEF8
XogLHIX0UYYoh047f1WTGmCKo/71guWWdHcVhROsju9vZIxrLfC+5Vy2DI00jdv3
wfjzrXoFCjZGSNVlmJs5MRbv+zraKV2+m7HsodkugRSDuwTZ7P6VQvWJKxdt0a51
j/L3/86eA0a8299lNH7TAk3Qlr7OJ+yzYVrjFFaZXBvJcRgKBUUrUa0zSig/y/1L
tISHjfkl7B0lW8sShJYljOJ+XMRCjcbFIinP4lvO206eRQsOFHKkduDBO06jt2PY
wvMn3x6cx/Vuz/OH17MMFy0N+ij0zylhMxr2VVJu3vIIeyeNwCtXZegp/XLm5ZfG
cUUiMRGM23wCqRHlO4PhFTRXKod+Urv5Z/aWXKa4OyGNML8yQwe4C66EBi1wB2Ws
AULuyzkyu1pDJSCMYTfyhs6lT0EujPVFfesvAIhYBsm+uCuJa/RBgZYSMh1Lbb69
dr3A5+U6gz33QUQ7Vap5xKK6Fztw1883Pp9cf7+c4XiSCCBfHGz9KmS8U3g2xi3G
hJ94yywLzyinVK+7JjhlnjZ7xJATiOxx8nz8F11R4qOQu1kRJlDlTxElwvKmJEOi
j4h9Ns5zMniz09e0gC3OgnxVaZWhmilUb4rjxKPhCG6VKI4PUPwbbhUJmj/S6adG
ePCSI44c2vB2Sm9Uco8PJC8KG2fvWIlnHjrJFgrb+xETxtrFSyr8C6RDJCGOHP+3
60K8DPIODMmM+z9WRmZAUlEwj4r5BhBK32UiTMQedDdRmr154rJ2J2xfby6ya9Ga
6Zy1puG/lJGYFBuWMhyGNmsNXlzBvKG/qrSjaxcKmm9e6FYWyj5LPw27VwRHh3SS
ZXiGQdeJmWWLRKITUoNi+R0cT4zUZoFGkJH5RvipID8FPr5v61jUo7oVpnrL+Nb4
NyTTFvy8Oh01Z8rGBcPoN98bqWpGnSf9V0m5B3DBKhb5ggyf3sUC4NjvoY46w/NU
C2Zqz4JqmKV6+y6Eg9rcwFBqQH/UJ5ciTd246RMdPMrg0fTwRNaBRlYZuv64TJFg
H954DlcJDjIOaV7qhASQ+JCC8iGpHBOF5DGYTUTyVT/A+nVewwiMfRIwojSP57Ob
4k09rEcqwBu9CFf/NQmxl/XzaKrQr6/YkJyZqb6bhphhY40tSjqG8fokshHNUtOR
ZQtzXCDmFNlWiJOc9vohLtg115WE9KkR/Xx+fJkc9ybSZRQ7Fn2z2EGueqzqTpIy
vsifG9hUBwh3uHql1rUSi3UkkbNmYq+AWiYRJ6lfW5M3S/mV1zY3/1cMzL+Eaqej
Ek53WDPGI7UiZff6hxjoTD/MTLi7Xu6FFDqCxGHEyGKHhG/OLi7YpNP1HvN630R9
po7X8H/pnCV/R+kF7qNDsu9AbxQD2bT9RvfI2DoihAED0Lc4LyWuXl7jq1e9NWRP
nPxfpaDYVGZlN/jQ5XCzaxpa6hMGSiUY5BhZSX/mCzSTS5+7W6jhmR5wM2OwQJ+/
og9QP+mvgcy3o7B5BhIL9SpnRbi7IirR/wJeVGSR3WeadmFpqOz/zHTx286Pzbc4
6Nrv28pDwI5/xvb6bykGUHzCKN11wHYhq2C093+Spm7wViSXpU7zBgzwR0TZDDZG
leJqd22zUl+DobBHKbU0GY5E6WQ2A2xNWQwMqdR1nG1440l4wMOWcQvnnjCGRvsc
B0Z7xR/5RpjH7t3OqEt5Nx7yQqxZLhPi0eOxA+mfIhFQDHOORhTnWLi3KzGNWxq9
a+09ebx1QTa4AUxHasQoXUG+RodxWjIhIpr2duA8kwElNh5rL8J0xNmAxH7Rs0nW
8x5rXyZtOJEMe9jcOUSvY7Fq4/1m7PQljPnVNbYElW5AWFrY6HKRyxg3CHtGVOFF
fwqKmoZjq16Cmw0TPydzcMnOhPXOKNwFBxwpxbUvsqWFmC3m8yl8Fg8cQEPy6CZm
B7n5TILd44K1bauduSV7Q/3Q3wmBvGFd+dqwyOUmHPZUoZ3Z6T3N+HObMc0Uq0UA
t7ti4AZMZvtyHeei34fxMcd0vlr/v9TXvL4LaCHINRUZnrve413/48Tu3CxSucVS
0AF66KX99QwPdaXbp6HuVDFdFPxjEo7+dh1089GLncAjD0A0e50pd5h0/J/HGY/K
BQioOGmd183vJu5DFTXf1YTW3PTVu7HkBqi1Oi+V7HGdH8UbhV4yc3Qtgs86P2RV
IdSm/+OkREKbGM1xtJNzrqUgVokTSl/g9A23j1h3tB5dfggPlEJFfCIHpJhSMbVD
HUWggW6vp8t5fUstjvVKLC717pgkw/9w3ElBlELOnf44xrNeMcUWqqFWOKg5l/ah
aRFBN2mwYVC7vXrWCZnabwVDW/F9/xetlKWXUvDyUycApKIa0f8YfkoiZtHzlwNF
5xEz6m2dbyyaq/WLB9uW0m1+4u5LIJZ8nwubsQ+bZ2HeXY2rA8xChWdlXn2k14FG
tI0cQ3nQrQ7r4FwEbvLhV8juLYGuu8dS3UssBvWfdb0ei1v1ItVdzw7+cRPTWeEp
h7414CBTwM9Msd1Bqueu7lLxsQurzPTAUUHU8I3K378+U2eHdiCinzi7AhgHi6i6
r/l0sEFNTBFd3zmIcLdQkv520qjkGkciRrPu0es2d6s4mnG89Dd0OP47G2sr0jbS
uYRmEIWLl3T3z1Zm14rkLMC9sw2JRVaC6JkqedTOQ6tUxpNc5pngS0KGAK94rJKJ
Mhek4d5su/iGBY5HA+6PAFzI9bZXazgtm/9AnUUCOQ5HaUCf0G5KV9tSIm0iGINv
v0msdd11wpkXqEwRREh6ALmEep0GkBLKcrk2WAw1PCmi/mItoIYD6AnVbFZ9n8gK
HBQNBYZ2+lszAZMKQHmbrE2JGbXZBKXGD+6njFohMgamiTeK3sWY6XE+y9V36MZA
LNvgTc2TV11LhNVREcuV5hnT8S579OLevb3sx6pXxbet8ufbb83PqIertY/ewa7q
Gb6MXtKGuChuPr8jFh3C+b8t+zlhKZbML1Jbt3ZyrKKtca9Zbsz6iqIMXxW392je
BbnOrpi0VEkAtxlIZoSHPSJ29Fiv7ysYYA/6nWTIgipiCVzDCbZULvcuKlCkx9GG
eZ2Sj8twDnbi9/TWQVdlGB+4/DbcpvWBeh+WVzELn/UnQ2Co8mKPP4yvZXC2OLZu
ZGhIPOqcnLcl5ZK4GX5ijdfUd1fiddH7rADE/FRMJB30mhY/ZWKevTGAaxNki1th
FZOT391iz4EKDVBCVBmRYS9kjEBm9M/p496goVqkYYDheLl/K0ip6x2Yc0Ch7P4Q
kyKO4FxRzb2/xG13Emwg1PLYA2WvLUqhga5E5C0qcjH6Ihxra/Xzko5wNhUETgva
fNEFXKA+jBVaWRjqyCN2xByKqBFp9cWdXhI+YLX0uyjuxuFQV4QrFzqzis5r3FaF
0SBeq8bk8PZwNLfMp4GQ0MNVJJjsAtEjYd5/FmYAdUktojvn2BFKtLz0Bg1pLkyb
uFHrxzu39qlEkZQGk+7VtTBH4p+ojj7haxGqa0DJZQ76fHqUcjQNAcfB3BHxMXpB
xk3A2n4yPH79Tt0rhrKsQikoCFP8u8TSgJAss3wN7A/38jfwb40ozvx1KgRMOzo6
TTxbbdhrE6+9/hEzk/0Z0FfPASjiAT7nhd52oLNdRYgDMf0edeC8o3NouIG2EOYP
p4vKLhNNhX4fL20yL6FSAbQO0oqm/ibM08CggdXIEJxPEHNSRuTnTRUg2kutRWoh
zhtbrgL5C9bWGXetwMbLnXHltIKdf0I6RVI0D95QpdiUuXlwj5iKxHeh0H5cBGfO
sYa6Nt4d4GAVpH5aO3yL9OEOFpF09HrWmdJ/w7YAXwjS2zua1kN8L7iP6J4riOcK
Zt++vH0Spk7bQofU4ZV8lCMCvLq88trsAvWtqIMd9hHolH6vQ7CSIxTXPv6UooC4
eL668/4bLw9A82IY5rFKdGPkBZc4faLvth0GxKcpwD6ZCK3xaPQrMVJo7PWH/4FX
CBUmneHjAYIg6u/S3e6JC+385Ccm/Xm3vxh1zZT29WIK9KTroV0+z6oiQczXDGfn
6e6gshl5Ry0WcV4qt6kbeS3PFxxfCUUIY1pZC8MG9RqzwZCZ4ODa4iMStBrAGvuA
0cMc15ttUvN3KZZZUiY+ljvfobIxcWP8pYjIbw/8oix3Ck+2ovDWH4N0OYB+DwfA
i7XrJQ3oGLsW0XfYOHEHgG99w5XrvVEdQpmKR7IX8RYqHe08rrzYk2UEWYeXPYSe
dZLalJu29Vg+6FfwMbiCfU/tDzbqVr0U1hxuSBaCP3kzYIffKO/pwZ34OqT+5KA3
4dE/xcQxZqLn8N+akdw+X5ulUW0TZ5Scp25rqu0OmmBcWKmuNG7G1R69JfaeP2x2
ah0BkJcvjzce6OgdGUZaM9+mO7nm76tJtgQRxWCseTSffFH+t9Qc1de/oGN/vrYM
WCVvWqPkHLX+5kTxmnH/9Mw/hZV5A55xsYPX08SUtc68v4br15gldT4bNDSQW9V8
m5ZzWGKqR34Ir4VsvVxwtVJr0Egc+K5hnZP2FL4TI9uXzGsF63FiDO5NFzJ4mqrS
o8gUjGqIS/VjRvLXs+gInRMyMy4jdh9xSTSH+19a4krpmErh+masNveJ7SpccefS
X8Th85qdenSSTIvDOdUul4cMZQmhl4VKvj8qz/SZ4YZLRoslIcpYBMJs150AqvJg
lOgRLnAzfCSgj/gFwaAU68Clki8V1KwEBaMNMb652uUWoJaZOKIO6p3N5dugHylE
4HScxWrNJdNE9BQBKtDqr/Oke76RbmS4yShdQM6g1tOm6LsNovNqehL9NtrKGox/
4Ll5XFoRCOm/upt9KPaPy9GX4DWg0fiusp2Sde63vd10eUeGQD9vXUvwn2NZ04yA
E03/Y/72JJAp+ufFQlQCeaVv7mMGZQMicLCtDIck4yG43zg62dXo+C8TEMwOrIOe
kVsx89IiNhGECQpymGfc8dn3n+i8jECtxg9XBjm9mhRUZrSvtuk3I1bMAFesxmnc
ZRSRoh4iNxe4IW+ijLqKfWr1MQN9tW10l6yBXcKOI/2IZhUEcQZww5o0Eon7ueyA
1SdIjyVksQn8CEJK1cQgV6QPUzwi94ljd4VdFv+hU/FAoVxH2VF5101xYrwxE7uj
i59l+DARh5a9VX5NRVMtbELpF0x4uzvb6aig7lp4k1FZnbwzkg8POAQrtJCWTxBH
iolvFDX5WtRhHEr2JpFhXvUQ00rn6kNOUWRkMc3LqHraq963KjsUEquizSbI6dRw
08foLysrxuoG7zAW814DdJ6eSVrut3h24uJCbFOM1S+o/1iEXANoSTMqbATdRCp6
Mhpc1TzD5AKkCCj1/oHt1XKY8/h9BPuwTFRksqs5ebZCOK5bPJ9yR5vrUMEfZPWb
2k3RMEEKmwOOSgIOgkmNF8YxEQSMe0SqBP+iQgyp9a9/lHoIHk4jxGFMIYeQSBRN
m0hgtenXp9LC73bkzQGs5M/XX3iEiQqqJh8tlCMNdWbeW8r4OkXX/FLOOhJs7phO
NZBgjUfjXt/grVvU0p2Jh7+qlVHEc8J1A4d3CVR/WQQrKF3jh2Jzl6bYooiyLiiA
j4YZ7NWyMWCcdVtim6AQb9Hg+jdvJc/INb6xR2vce+AbZNs2mLsFzpCPA/EHcv49
A5fFG/NkGJ8jxcKQqjUr0NfjogHt4RVZUUflJLgtH2VhPlbvV1FUxlGOgJwsZnI8
qdGMesbWY1swdcZRoUyDV2EKEakinmaGN14obJRkcUF30Oj5e2w6WmVmeEtse4W/
Eh8+XwS+p1sOWzPI7aE8TtfuJguerq0kLyWZfdAN7mGTzBJJSK86sr2gbKw4s5K4
EXSmiMGBz2efZbAl2YJ3xNYj8tsBuiDYvEtUW2YUkm9YJc1OD8LUVuyURt63tuXE
SfyqyPmG4We+ZUMCXfYX+2rTkLMOW7LhmvZLVRSXtd3ILoz+B5i9dcGuNDRNZCFT
n5B9w/Y3mN0AzIUpu4Qc19JjuNbls3XQoP2efLgiGXq3NZlPjtJ7CRy6aTM7Tms0
e6V74a1MqiVEmWxk2dbZE5q9lLXqDhOYZeWtoaO36IPe57d4+QHo1CtW5yk4ocs/
TzMU39qxVvedgrrcRQWXExno7cVcMn0sL9p1YrUdWx06w0ZcLl6g1AmpL2Cy9vyh
WsU8Lqs8AlaXABcRPFgSoWjmovo7BVIlhEkv5o8neADwmlAcNsbdXWmn90DHA/jq
g2xzk6o4CtKTaJrbUP32Mx09fpuWZZFQhzjyq+jRnWz+8YwHYEb33Nc7k6pTKf55
RElsrs+BMz4YTKneB67imW33NNBMya0+NUn13npZahI3P7L6Y+yTdekHTR1jvVux
ajtAQrGpRm1KG7c4fmb74sTtx+IFDDBMtz/F5IH7ZgFboZJPS8SkpRjVb6x6yO9U
8FyCVwtIaoWvJ5THf5JLXwjDKoCSucnCv5+QCnJ9MwhFXqCj4ojQWt7HTPQLzgQH
EEEjQSl0VRvkYCbGd7UK92o7wl6+yZLulDKwCR0Pv1h0TqY4kI4sY1Yt1pJ0FBOv
RZPc54G98S4ur2zA7p2Efg9IeVA7jUvjRINQ4HeKgNJPJRoBlMNMFfHXR2j+CNr9
zpVQT6MKAHk0p+hXjANlBSDxfH0ZnFEw/z0IsyljiDOmWbfN3meuMXSHjDhC60Kn
BXUBZyMxC2HQl/iY/spuI1KgyBYQ7QCKXO1WX2/TFjSHEIEMC11WNYUfyV0fpeuJ
3B1SFUN0o+NaL5w2b0Xw4Z4CFFN6hkaiq49i4JYJBmBbhLzkrUbnGtkDzsUoufeA
7uWR6bFGVnqsiGzKRZPlYBULNnwMpr9CxHq8pxLIXhQfYQIXgR9qLDLmsxioEUSG
z9ef+faGzZyJCOtZkOqZPR1aeMnVWZhTK3K9YPYXrnFcOGfVaRnTH0Bz/CEk4SWF
zqXdnumNsrfeLOJyoPsbFIChjvdzLAdlqzV27902laQ2uv3RVDPDenUM/2/mOeSL
n3cccmKwnThlpJIOcYTBeRknQnl7Ww32zt58cTW+fOgNoi4JYmtQyptYvBFOFnl9
p9iVhUD28jUf0n/wgfhdP+s+ImWAni8ezk1kiw/tdEcdDk0qNCGrZ2kUGr7y8zQL
yl3Lex6G2qwipdL0Gbpq/Gffs8OW7LNyay+JYGhk0lUki46rRw56xv93FFR3iSRe
735fNN2aIdi+ixXWhH1LtOIfQbx/0xM4Cxk1Wzeacsw1iOdKvLY8h7CMyknOokMV
UCqso5XnsBnt0CRkhLy2WCep/7JkDrxMqBpa5lp4DaXfkfPo/VbUVmyAGJa0sbfu
vlgKwma8sRBYxkjuHFUgi4ObpUZI+ifADdcM4B/29zzjcW65x/OCONu3oZH5bEF0
TPVc9PDCgPERtDwSwwU2CXdDYJPRLwFVRxesazKBu2vzyEsRr1gXOO7PaDf7T0At
mwYisRjr58aAxfkb1dojA/MiSU9LkVXuG4c5dUiQsLmlCM3TEoBrbQI+lZuzkFxu
dzcDoQeEb9SAOwLj6Os+RyAWr3uCA7tUlG1Vqtmxl2px3am3FlJA71cWqaMymz/d
8rHpee3wp4PafE0T4HtKtRPBG3G9hCp9J0EvFc/F5ie3JXG9qSDTN8Zr6S7yu7c2
nUS7qLhrqc+3WV5pyHHfTyOm87c/bGlT8kNIMMcnpelQOKkb/VBzxIWQvt+VmVFs
1nhNwPkJn06mTO0LdfVYm3b3yrTPqsv3U+EJ0eiEGF88Q+fKBKikWBaJSfNS6Kp1
ejxL5yRrQGnxnanIpgfIWqIwsJIOalQZH3Ruhs4na7JtzcHPi8jlZEexgkr1wSpX
XIzIbs2yUkAH+OPn1gxTixg8zyjTbSnfDN6WalyQpw3ki2IccmE15L0pjjPhg80b
hUouYGLuC0g97dB539lsNt6hcpfcI/vEc4f88atlFCTuH6rS33w4ogOAaOh4W3qy
k3Qhj+Bo1GGfwM738owi316wXlYosfMcSOaYgCa0IEt61VipbYy8sPYiBrpNdR+U
tDjujrp5HjJgcuKeQ/bywfwXw7xRJG8Tb6x4EPe9GNWR2Kc/VOqsGhnXYXUBfezO
FFiYBS0UTME+cxri3M2WBxL504jbg/nUdvLCvzcvirPx3Z0GAZbysbFHBJc1I+oi
JsK5XeJKiJz9JJkFqVgoy03UUArZgFZiBEuKC5qsFeYwvGt8I3BYQfp5lJJB9VCm
N4w/7xCZz8yjx1jF0yS+wdZHFt/yPZjTM6DQ16P2WjCe/8HbpJlowr1l2GLR0dZD
M4H42LAId7d8GKgy1DyUKar0BB7mclx9q6XkIKlmJ+9Mx4/bwwhlZLSzcDHCWKiC
a9kke3vlaizWbc5Ny6hg0JffFNHItub5C/VKlLQ1s80q0tppEst+f2bcHJ82geAU
u4uimD/tzBu8lisLQwpeusRRm8nbJP1SevijbAXhZp2nBv719pk/YUUM1dJQpS+U
IfjV8U2x/zLTBcKgTw3it9AM9axMO3tcUlOp7F7jEqqNiThf4ZCXWGt5kGSivO62
el/HC01ITBJL6ln8S56LIodkxEtkNB89fF/RqcxC365Z6kmwmHVLan1aNQgCZw56
M+00+ZW9PjPOfeMyNasG08tJ0duSDZx7+eQuVat78BcWo0wWUSH3ZE4lRuUhkeTZ
MCqOqoruHnsN1piMmSzQ/+jzd4KU8IirgtgSOCKEFTQe4ctclLAaFIkN8ZQ2YZmW
HvTN8ef5Q7HwHDrqaYAQM6oK0fHKxIDLbwZoO0+D7uBDn1L6wSSN7wyWKDjyUhOo
OSb8rAC2EiXqTuGogJlgEpe8cypupfyQ0sHwSNAKSUzfUlGv0dDx+O8N+PBAD2+d
fysRFZivyKUPUfhU8nRvcigjROQj423DOlZiNV0eFEYxKZf4s/Ovu7bCF6SbyDfJ
19s6PZArMhHdqoteAkH24coRKG+qFnC5nI3oyqBmH4l38zB72zaI88DC6qlmhHgM
YEINpxrUMgIch2npf5LaOjcsKst7mtrzxsKniFLnfzYUDo35f/5JynrOhLDQZPjd
ORnDF5m/U12PzQOMA28xJWvITFUJZfyWokX1N1NtNQjAuYWFqLWP/bJUhN9L3sRQ
0C6346S3cbnZteh4UPuJFrKSQbQqpJj8iEp1iPWQevnFlFlmoFakJrTg5MNEjiKK
dbBOw+ZvEF8w6X0BggLaBw9U3LX0uAxjraSH2owbXOUNGTkNqsBfkUfSCG3Dw6Cj
T0i07R8xd1iM5AYhKOjWLyVmu8jIF1urwhHuJvTBJ4c8SS8b9cm/RaYP9ECkV+Ow
PK6ZQaZS3uQdQIjzAeydlontB/v9PSPYdmKdeKr8XkkKKgIIGdJZOiDlmkVGrr1I
Hj9zDVC83cFxj9N7y1p3613PBGclWRd7DfM8eRoAN5/HIFicYC/BS2i88Swed9Ld
uo3k3lrp2Cm68TvN6/lIlNkUXM7Xev/TF8IJ/Wq2hRxRW9ZhxWUZU7IizMR4GAwn
GCGKva27LOzAOfKFvpFSCiPMGbzCV3jbRMfo+mA1i971BKgCQUKEi5AcJKH3VSsi
8tA1TOQ2lhiZhgZjR2062Phyni7M5Ga40BKL+G+0GRnCPmSoW5v3iwt48UXWJN0Y
3xJL6fhk9nzIfUV9lqtFDVttrRFMo0KSVWf9wYqTrldTPmRcs0kPdifj0lZ05ibL
pm571S9bSkw0kGMb61/0ZmcClMbvfcFEkmTYAXBn08Pv14IMjXqXLZ9a32N22hyd
RdqixE9AO0m0y3LMsX+QJPR5ZtPtKKB0T6RBYMN3xAo8SeoXFlp1I5CXZEuVjHaf
a7hVyfXyvh6NyGM3uvlKUDHxR3V18tOX6VobBhI7bncOSrqZDFN+iEOOndqNNvfe
enKNt+hmHhotERbBkbbqisGtKjp/808FdJNPHwG1TbE08/GCkmHmNC/MH2YaUVym
sfHLH2+nuW9oBFFA/qPouCrgViBwsy1d+olgichBSplZwnPuwEwJJmdsGYoWCkem
1NtLAz5IsOKiNIa2GH4gH2BC6uiM0RjJ5w89BgoY+jait0Vvax2Z9HzrucoqHs7s
IoS22WrWkZgU6p8/iCRuIXqwTtRfKmSnBWk7uRLgY0Tr5qb5po98nGV+LlNiCkD3
Nhe9xqee55pF2jKbfU9hdZeMS9KQrWUDXLRIP+XXLgG0oqE6XHxRAo8HTMhey2U8
yBYLnlfZzjIApp5znf0mpYhGcTvGb/eIFS/d8WDex5dMknF6zinw1t1Wa6ZjSlcc
xwS9EJzOzZEGEMzqWm3eoGlCVrDshqFGkmaDdxAN1iggrdCxqX4wjAvjcOAedSBH
sqOtShr/XLVfXB++cK1hdGmo0Vo9FL+wGyu9jaWnSOSXGHoGkml5CXkyF6z0deVv
hnmZZ0JNXkeOBsaq2ZBKVsKjG2hzViu6FuuxPzZjl+07NKJBvVmwBymPdvuIhmui
jcHdohhaTgPS7gZdBf/s6a07PKWXmhlxzhiOu6raqLmLSVQQTrHc+pMwK9jNM6mT
XfRZn82Kyf268ERlVutqMUSLaWHWUOs1FvLB7rkZCWny/7b1tyXrJZ1XPOCi13yp
EJE2XMsf3L3axm0AWtQrBzuRb6DeQaJ72qauKcsFd8cy9LrslCfjaexCdtf5E2QO
HVfE3RnsH6sMU8uEDoYyv6QddQHk1H+uVqw7CmO/JfWMuKVj8JiJQWZX470GLaRI
OERAwE68OwV+b/HK35SSG23ifsyHNoAoquWLHjgYKYbONmIm+W5oH6MxbMOprFHF
5yemiT48ku3J1NFn3Om91aM/nonG4ht3/DmJgJRe9BxLUUR6BntAYOCwhD7pS6ba
8OeqZDgmGRixGjt4ahM7hLpmgsiK0rlM92Dx+asrJeagjCZZ8+FW7Pq9oZYdrY5m
Dg4qX8/371XHKRvX9oAOgXWMzeagBakvcodT1R9phZt63E1SbUzs4spKq1Pc5ao2
dWzVQT5i/R9gcRBd3RSw3TvQjLop3f3Ghg4J7/fKMsD5JeX7RITEZD4FxmFq37mb
10mAwOtv6NtVhy1jMKPufnVisk+bmHO1Oqsbc5MbTwh5A2gze6zWSTOWRih8wo/u
qNxvbdcAI6ut2pIjsd4wmYJnFlQlYe5YAs34dd79AFNutl1TvjLS6yi4TE9slSYk
Lkolztj0TCK2gv3fP7eNaGvWr/Kc7Ur2rGSTLjgCgXtG0wS3ItsRy1ddu5T9g+WJ
PZpjQweS2HAPkyfJ/89Hd/65GtghcsuCILNCU8RTjFyY3S1WO8gTco3Jq7urpEgn
hhUL9LDdo9/gQWnmaPKEM8EyIh3Z6O9Gz2V2OynAh/P3zY1b5SpzxBbU7TF+whUi
d5aVf9V80RITqrHqtCr3TmWgYtt7APQMqmjpb9UEJY6iYROScEhK5ePNom01lH7e
P6+lwnZ6nL1sl8zODhYmOGpMYrs698Z5LyOS9DiYFIC7/CHQChWadPJr6QiEl+gF
VzWSMN4bQKjfY+50ZS56EIR5FM6B1VgbiNptVMAcnoHMVUmTF/RdfLROEybh3XbG
5mC9P2L6sry4bSA6FcNbJgYMqiBwL0hgWtm2yqTghzcG4FBZZpBtKEEL5T7MoK4S
yDzAWGODCaUjQMstghPa3O7bNUJ4Ut7+8xzJ6STi8vrIBFSCWp/+1jpOL4+hH/NU
PRmrM2Onjp8axyCa+6IWBuOP8h4xQ+RmLyWlU4rWPvy7FvAA3GHmEunlyUaz9Kbi
7zsjM16GiBJfgaASj23KQP8zxP0KWdYsyd+UA8hhflWL7t4JwbTNJG9ZjNs9Oaof
5+3e+MeYNsJU+Zo7kmObNk283nb8z8Gh45F0Te6VNeUY0nSr2h9F+m2njq31dAEv
LLYyDyz5C5NeGb2dJCK8uXo4kmOW4QZLD3tn2dOabyhSUCU+H2qMFIS9GAZwVxzs
Xpz/jVJlF6lrrNxfkFb9zKG3VPOeah5g+3N+VtAe+E1GG6+N4sMlR7PXtNZF4QJL
Jbj5kBPQ6Kmr/wrVCy8ajglYwmSFq/qJGZqCdmRIoKh0SQSZEFylmlfGu7In7iyy
EE5uABWK2TlScIvw3ASVqk+9DYLHc5FDEYk+dlh63NNqwb2Us+xpQNkN++IpzIGM
Vpau6WaljiSv1S9m98u98Ow5xRAvz0QsM1Kcfas5zx1PSHV3vDiuhebVRKu0LRvX
B7fbkZvyb/2pP/kugnJPgAIQ46TEk59xNfC/hVUqpMmy+5O/fhQAId4XUmmJrQzV
61GpASogIknllQpTQZ7LSl5Uv8/zHBPCrjkZH4I4FX6xAULfRcxClxyTDHs6F5WF
Qft/mFlHO72pK6dGCKmaxFzbQ7gIC7b7ALNU5WYoeAdi3t7iOsrOvTo+/b1Ml5cj
mtNASGrPSoXIuxn6o9PlEwYBTbEe/SMwDE/hOr691LkqOT4r4+BwfeXsNzGQhaJ+
M+e2EuDEo8nYJAZAFZvib5v/d0qwknlOk2Nj9//XbDirCpsj0jynshFNW4svaXc2
N4RORRvOqhsEWZ52YpSLFs2ULO+hwzz0lnYLDfQUeKhcwH09ZR/FyZnriP25jPzl
LZcKqVKwTjl0nniP7GAg2Z4CBUPGiXmY6ZdvYcS+OsEPU9YnEvBrZwdpEj8wk5C6
y8nISW7YJDv0lgBnkL8pmI5SHuoSSPa7FiwREhLtpMybHI1TQZ2dEmCH2qDrmT8w
57Xfbb7xRuV5pG4iWkyB4WA0s4LcVV9l0RHiAqdgmebTqzVzTjxiHxiSCUudVZEs
tOiuVIZsOCHxRpzvW3zomGIEeAio/S4UyG7aRbYDC/5EgQYKHGTr+drN3Dlrq9By
QFquVqq3KGQf07CgSIBX07nqoLBpdafjI0ZAfl5Iw26l2URVYkfyksgDWjByQson
eQeRu4Y6/4use7fiQ/mA9r1qKV4ExC2X5pNPqkUsQyNXxr6ZiCSDsGmUN694b4bJ
M7qj34h1BW6phx+czF37UElsGwTDqx6JZI53iM/xlFhMZurQb9R/slgOlHN1I17+
sSbG8y1Zr15FJ/9HrYbDt9plSNX7wH27VwielISw53jWrrRmMcTl3JYLhBD7eMs+
LG+UVAQNmBJow1kKltijZNhl7sxNpQHFixDuTNdKVSUyiwjMq18hv9S8L0SV34Xt
uGEeEw57p+OzSiCmrNXYozLj5wus2HumSRIaYpYHV8x4MlSenRvVQdw7wDzec0Lu
w7uactKLwo1gFrSOWPWwPdYciyWkceEGT7yDEhNySBUdfGwQLFhtkvN47Ya1SEun
BHDS+i7wk5j+qNwjt46fWCXSQj/VlT8dxEI0S4YmdpfSfn4evHnQtAiMSMDsO+Z3
0OpuZOeaKvoMrPOJ0GvPdLT29BU46oAH5S5WUuZCa/LBkdttdjyTOOTigZTYvgqq
uTZKSQ2kF26PELrRHPXi9kxs85yrork5A8MN3DarK7Ocpe/zxhZS/hC/OkFPr86D
Sa0QExG6JnlVRkaStXL3BO6XQnj7cqVTS67ol5F7x3nVtScJpGqjw1IJ5inL6txJ
0h+5VIfIItJoIRbirB/g9wpo3yzANjHSR2X1vaL/dP3Oe6wDdpOqK4ME69HOfNXo
CRfVwsIAsMXjyAlvTEF/nhpA0uQOr8jO24vBQtSlzm/6noZyeRaEVjJe2iG7MdfG
obQqTObIDc+iMrtctIch11B0gdfmkax/Le1VXM2L/GjJbVBCQin4ukpg+b5qhoo4
s37uM2u6H3AdnGnFFF1F/cn3j9ZENR+FA9ELtRLr+AWt1v1f8kT1FPB8ZLZ0QjKJ
Ynk9hVwCjM3yP4sLJ6D2cD73w6HBjtqm6x9CM+pHWke1ybtgep1aytWCkCLfTnBW
z6E38AK5JkQi7KooX9WdribSpkKiIrD0qXvG3Z5eliDAg83gZZezb1IUterc6iIv
+WDdW8Gv/Pq/R9vyfW5xUSyN3ffh0g6wmY5KCwIX7oJEWtDl9x3xzPpaizP1/eNW
gKKZoQwOTLxHb+TCqC5FuepSEMOflqDQP3zYIxUnsnz08y+ImQ5JIvtYqK1kBrZE
YX4wqMCKWTUZw3fjHKa9PSdxP8yt6Z8uYF9fRzNIRqIpqzB9+6W7iexykSzr2zrI
ANEilAmsariYhJyqNgl4TbUulllxbbnbaAaknG1EsZtRYqZh6TwWIWxZCpJuSMfG
lTnvQwes0KoCAqjp8d/9zlrH3wNY06BTAKrKZ+qpdLNAOQC215ZjARxVGs6O7fAD
kWOLGKAZF+zfce4WZtOTGIsYTolgeriHBPOEW/Yj+THEa9XmWa10oanmkkvyIjng
I2ijMmg8utsWlsRjkPGZ5rK9csf3q6J7aFXVRQi8Xja3ZaCIdmMfow427sAmTmQR
wquR0dm88aXcKXnvR3PJDY2cV9Et2a/uuskxrhPqeLq2sfrr5rjZBNsZ5Z9jzqY0
fu/u302R4DhnI7CAulfCxjIJvOjIQ7yk4/rP1FS7ZkwB1LKjIfh1tFUjRNkhjRC2
Q+eGkouo5+BZJeid4gSiRQXX7BljOAhqSeuTZILnQ1UQsHyb6nTDNBxqpUFzWR3A
TMVJlMKeNWk3n0eKNRUyIOmD+0EQHAjpShQKoJvgSRiiPzv+JG7heWRW/FNrh3mX
7xbAMhjiCDe22sEVTqL8+nVo78M5817ybbfR5LR8MSslX4NPPgIucpMsOILEFcbE
dUltVY24VcZ73NmnqMW8t3QZxe9TrYfsDKksWSsRc8fKElDUO8ALo29JZVSabGSw
tejED7pSKFLINPuVz7pl1AbER5SB2LWl+TCPHlDtnHYLCw+kPp0wka3X/37Sv+Tg
TEdAVuSwFUcee3OuSVRLTn7o53N5xkLOqsqZMI23dEznvx/oaMevDrtilrXWasGZ
O5kbLv9HTKnVCDI9T+n6gcLK/71rQivKsSBPUdCimMwMeeiY9lEP8kyosLvy0ETN
67bzvxam80G2+RH4ywnbMnF953CxGfwIvGAJUkSimj4V2Tfyqw8XC2tQECH7I4/u
M7vztY2vWfEm4/Ll53dUup7RrHKCsRdpe4828/AZsMBldp1RGXBsGE7/F34mHDKG
MwAawoQhsZYTdl5N7F4EojpbvCLwWRPTTN20DPYLjVCE+UmgCxeNwv+MJ6Md9tyP
63+8GGzrK9dHZL7H9ZxlMDcFTUnSsCwznAnDXYyWZJu2eZv4BVoY8GIOpDAVSLJG
vL17dEj7s0FZLho8nv29tJIa0zj/gFHnpgB+6YZD6ElgKwVYd6X9ZL3hAh3Fh7Ox
zCn1zDAc5g2XNzCwqZqlrtNiX54K7sSo21W7Cd4oQEiAC99xHvikd+h0Ett/+DBR
Uw3fiRdfRzdlYha6Qqli+8pX5LQn9VR0GpS5cLTyweyhBX/CYvip4wHoDc5esnk/
oXkW1xrGZdQHA3t+pc9CLQipvJrT+FJ+Sz8A4J0tSYy8eRX+eacvtkRARfTJSF+W
EOIJVWCE9qLaMkAZRU6K/4oM9fYL/1pVaIViOyz5vzMgLriD8hCKa8AhI2PZhlhQ
pOmv0dYmbNC1WnPNp3tgD28aRwAsNP/b5lf2NdrpEgzdYYmEPI98XLI7G9L5ADFa
K7VH5xRWm2X0UJdehYT8ANpr+23QP5UrvqjZN/1iel0NAtOWfa85oWjx5y0Xlpj4
Rp/z2FDhOJzTcqjnTcOFhz5qqJrRwZsNTyKUuxG4ZgMTW+Pzc+yBlslVd2A4S3Nk
iYs5Pq8dRV6ziTMK3LskfIajOSvg7pljnEk2iLKRQp8brwHPFWoQiSvpEPhOFMBT
yHWpSh6KFVRvFyw6DDfwh+NLlYSKcSLdjAQ0Bj2tun2egfuLIxDxJo38yXoL7X9N
sLqX9LS0ZUJo2lTRaH1/LsYIql1E6tZFVd0Ox4UPicXtKMW4ZZrBHe3PfOWT6HeZ
j5iDIuOkE06PWcZUsfAoJOxe1YEHOXC6a7Pxyolls8YS/vAL5s6HQqEciR5YfKl6
0XNy9gMLivnTV3zhLsjLQf/EDDSat5aJZJu+b23c/Hy+4jPYn6XjfFf10VfVTDPn
8JMVfRMwWGxSEkm7WpxoE9KpMymfXnecQfzzfCc/solsn455O3wICgkqdP/Taiij
IC0HgsjE/u16WQMs77frWyyFyScJAmXElMb9oDd/Ng2NAdsDR2AWhVuokMxDj/Qq
vivWNNgxOJULsCTdCUsagA29Korw2iZ4vnPlrH3FfvMPXxIIt2871JpsuoLShc/k
9jWQym74wRkcaoqyLeiqCBFZKQD83qvIkm3cNEsKejQ83rhmutO+JLefkLWubrj0
Gol/7dwjigJbG0RuYVtbrrYkazOCwhN1CrWzFZiwymjLSviQ2K18aRil/3tilxGW
5hKYClyj5OvmJL6Gll6J5DdM1kmrcZMCS1nxzXXKEdXKzjRlr5qQavcBwvMNSSJ3
Agt/rfgKyoHDKuvxuqRL8+C5Hp5eWjtWR5JjGflUxzZyKs6GjRsFpogP0Zp2GOL9
hF3ZHt2z2Fm83LAgKEGlgw+e2BIPafBhZ5kq3d8vaCYPX3DxJjUvK5lGsycDcegK
P+MJYlbfwgla4+ZtqQtwoS7P4vV72TAc3/qafMsVUktYFmp83IzkNQM3f7BeplUN
vf/dffLPahiMhxQSKbPHp8mLdYaA5n/Dmd0UKWo9oMMV0JdTCxSVefQK80Kck+Z1
CXr5Z+TzCbHv4o6rZRqYj2btamg+Ousmp88JVq0TNmDiUVDh10c3TTt4W3IbGdbz
3WKeQtKb/V5vlPdECrwYxoNklRPIGXtkvnzpMiYRj76itvvOOo7QoxkrCcd260pR
YfFpu6ObqN6HpO6qq+Rod/M6NTSpG1jPmaxwmlnYNZzOoCTM45iw78OUzUtOCxSf
cLDaiEwK/pvxP4DE7IDAovKKtpxWQ25T2nCkN3+02iJ3apGIFWBpF+63TNHM1nyR
7ibDf7lEFg8YhnUBlwNavCk2nmcKvgE4TwXemJ18cHIBsrkSp5dB1qYrSLlByp7d
n9sGj/feNgGEAh/CUEMd2pEq8a6YEWb0DSbDPiRN5T1rZvDt6K5On7mZuJzN/cJK
y7xjvNEv5AM5IMpxGlxcWGeyH+ay2Xxs7zuFtPguMqKRsBlBu1DuXqWiLPNkBqM1
CltGJU8JR2GMtfjjjaDkMtn+dkiHKL4ukRvFfBYziedF5t1zRCsvgG8qhwXNOYeH
OwMKXTFHHQm+B5R7TH+jPqYd6lEHJPXQNV+PFqtEeEaXElJuOFWSO0SYseBtB8eZ
iHfO2ZHtH4C+qmUfv2d6a6jsEix638FYHcOuFxBQB9pjkj9rWYiCP8679Few05AK
aP7jrESbylHHoyOWW9ioKavVvZSOTgYEehBHOXE6MWJObTuY+DeO1UMlx1M05Sxy
kOjm3hHMQcR6nWa6SqhaveVMnyGlAIH5v4mq5kyo86SnpXBclrXJqXHPcCS4tUCP
j3600ZIVGPTrB8pkySfidaWeudHgC/0ggXmv/j7gR0+vqADGuF4MT5RhK5soypTb
SdkV9cBS7qHlENgwB719muBZNyQRf+FLeEbxadX1VSeDO7GPKNDrd5Ueqco6GFAc
75fnsRXstR2oBGQF8b0NycuRmwlM3PJC1RQ9uXx3BfXxVYQlPZBprE2uV8Wei93i
/NpWq0OKYZqef4oma9cogmEWAGnBpD3/RPHNYgk3yxzAxcWwHmLYgQV8AMgBfaVE
FP3iCO7u8p4FvaDYvr/l0IykmSj02gUxoAs3NNPoHBS3ZA6jGpCs6swzyK1CaT9Z
mpeV4KSJnSy78z13voyYB523BZjYlE0Vcz+5UsZjiZQ7t+VPUKHobv1AtnKPyn0o
keVpV1LkwBO0E+drC6M2zPLynKQ87WssS9fPa/aQnW5/TCoFoCZkXBRc36sKhj5P
J5o8NBWzT2Qo01EkpC3DvVRr8eEJg9f/Conizu7NDfd7rqfaalHFUc1kyG/coVCO
tvZWNf7+LimVW0hB/mZ4csb1OeyjrMF+kMZSfLayyfY+eEdITMv3InBJkG6gP+ZW
pfZSYedvJLSQyBhbjo7RCEbDj/BYx2xKaW20GJ21e2TpZEHRALDIMIaduzG+DLWq
eT25mW82/vLOD5gC7J3CHx0U9t/lVIAxB8eGO0/FXYO7ZY9GGw701iogT21W6hVy
QbBqjCmtyOJ66TzlcQbQPl8v7+PXYpXlcSSPZPm7OQlj4KuK9Fc1SXNIxe8bk+Yp
+NNvKSFXH29bs4joNFAZmax7BzKE5qnw78tT9Ndmx8wjvhHU8xF1HjhG8nLbgdj5
7JHhkwvYL13LFRUGIaCO3HVRMXzZ0YfLFURWPauJ+aVMQVGrGZgJrGVd8X1zJENA
QsZHLdc44V9PhMTgIJDguXi93bri6LvV3lpI5CZNKglQ8jPZLFTZwy3QXYd65aZ7
0b0ZdCEaoPtDLwiSxIJuK2Eucasuh/fhWG5sGVyB06Xp255GBm11rM/IBg6PRzxF
6Oe1fQ3EFlMFz83cQZQikzuCUHaXh/Ej0u28YRDZmOC1gr2ptAgVCB43DoQfr9yK
jGWh1VvaQT1v+elnmsCCMsgF6wSThK9fkpcJgC9AaS1FoLWkjfxZ+XimaZ8oQ45i
c3IzwdSoTbK6CfD5OlAwbmphIhS/2uMeJ6Wi9uleXHfW7fZ5poPxv9rvkie1evPo
i5qSgZ1iGs/ADTUaUyy3UP2mJ6l01gGTRK21Z5C2NNARe3qvUm+4C7gmMyacwZ41
ESG0/HVNJ/0qGEow6hV5RQ9fn1Oe0wU6tVW5F/DJF1yToR80JYH6iOpetQbIYvD7
9h/chnxt9GBk9jftIOSaR+pzCEQutDLfV7KBW3N85ftVVaJhX7kQvsY7nNtMyC2y
YWoDtbqTYIMQ++L0Ca6Z698yEXDQj2cpQTwRJz8W5pJyWPygUrZvk+cfHlEqXQp2
8mnxRLG7KbESTdgbZAwA+KIGVQ3ySBALsDfKHDNEVNBeYHL8CneSDz+U4kmSEM4k
jP10FYH2JbrbAOZsBjyVcSyUyZ5Mm/0p9kM7f8hthEquWE6o428gb2DtLQCSs6wr
prvSCtIIlK/7P3VhSWOgo/sIMELU2IpP5VjwflLIpEFWccW8gpNIhtBR2cVg6YyU
QFM3OK/deDyLz1J582WXpd+Qpd7ytkXENUwmPGOCJPgoyiQQynMF3T3P+jP8l77B
kEBFoTe4dVdcoblT5ymcM20pcQU4XUKTdGRWQX7nNOqsJnsV/iPEM7nefakUijMU
tEEuMkTmmbvwXjAgE6/MeS2QxSfwYkQ3CjbC0+lc4NCbt6GenCEM5UDtABZNavn9
IumoiXpxKd3LSS6cxKQ3QeCOXn1p6IT0lqrhATtsWGCo14vT5fPiEYmjeOhYdtVK
eGfD/OD/Bb71yN2C4W/PAH+q2kLFssfGgu0AkVq/vyf7FnZTQg498ewzHE1HhInx
fb1Vf/rx3FKyGjnLWsCPhqllDEn0mWii1C+xVQb+KB2PbFgk6+0TjiWo8+/aNNNS
dY5X/TgEynil0UlYp4oYeFHcx+6nb/zcjZ/9l/2OQ4Aon9fLjK8b/YmBK7CpiEnh
xIuzCOwgvKubYee02pywnDneSRTD1uYZe3heJiYFXtAmQFNzCLWi+ww2en9+Ik9K
aZwQlLFHsK/cyCwqPjINxzeWHLRar8VRZSrgE+zkkAzCHQZkqgSidccqInpDh8ny
KciMJef7RMGjD3/PtMOkeDrKZRQQ/n6V9MM42qic8ecIHTgEKu0JkZ5ry/6xRDjW
r67FafVDr2zDKf082KpVkVKln34EkT0F1mCNFx/45dKpURwfUffjlQU1smES5gEG
yJx128AKcIUMSSenjHwhoE65W65IVT28qUXxCDw1MDb8tAivd1OQhJBGEXMerXjJ
n9MvB23B4xfMOdKYm/CdLfek+Ulxa79twS/G4jNzqrygQh+nmF+9Pgxq+FA6HcHV
efovNlwTqkCtko2C4/HCkIOkBziVhTXJQTGSo7xM4s2SnXp4jD7Op1vtQ6tLg61/
lQN3Z+k/60YzDNytT5eP+3KtA4Q12W+crAp8tDFcoJ606foHfXyr6+X79F9volU7
qoFfuCNi6eyehTzn00I3Dtp+pbFOEzoc8WajUOp46u7AMWWqJsPZSk66rTNgBCaU
EegfaheRZu/9Q506Qd8Y7zvwo1gt2dCvtIn8venQjrsfLNT89SrDe/nf4Nuk0Usk
lPliVQ6QYHv37UFbfU9xwLQCxTAjoyhzJCwLkNFiZX1ugGhDeqce6r4wi6iWdSFF
7Oe70WcwQZoFBMsj2ytvDEFJFFrQK8Jcf54fAZ+aTnNbwuI9Y1FGNTaOdCj3AXwQ
YXgFuLThkjV+Tm//fRmn8YkaTuDE5mZBye1LgkYy47zPNNjzTaODLAKnw84g3ARO
P4q90XumpLTAYZSlfWicYx61EESqgHtBSocq3x2YCWVYanwX0cpZJpXbGjX6Pajy
DukDQtkl1OcOvyB/z+wZvf6Mo/hZIXXq+7+wG1INwolwSQaMoBT0HiSz7lGLNF+l
rNdnEoUsHLlktxy9QFoGokJi6UEv7HUgmChKQLdX0uDIaCNI3LmX552nEJLSFK5T
20MMf37IFR7h7WxrA6/saDLKx40+odSDWScQ/26Xj5tFWrcpMXy2xFK78U0+v4Yx
ouMW6TWw0yJ1Bf7MTBMNZ9Y31LgWCXu1xWYig52MwKlvk/biy3l/AlSCd+Ae3b6r
SoXO4MLPxYIvjNebv/NPKN6ul1CahElLJ+yeaWAepuKKToHbgyrchD7Q4X8VBkXN
qN6+wqWbfD5/enbdnuFLu0dfn0n0iU8CuTjvLG7hb2YhJu/C6AyNSJW/l1e68q/a
HODd0lPbB9QDb5Is+I6e7w==
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SCESLccbGyh9GpZ/X4g3AIEBXQWQnH7JTvwyy6USXxRYg/wz5wfPZFD6a1QZZ5cj
EuLxp3LA7VVSZd3ztzVpLUIc2OyKb6x9JgnvPT7jA67H9O2w8M+f41peDXKz36kr
4GHWUBf1lkBQfdDpgJxboXaJsDrcgjdo+AvY+PTqSGU2AgMWpvI6Ni/ZRYq0CxrN
WDUSALnmnWB38qWmxwWYOpXjOTxyoJqmRUiPoWtwyrDfGzOxHJnxyUbLRLTllCcN
Q4hBGg+hS9PWnBPvMpwQSWmEwHHhWPPoKTSfrTreAO9vgCjtmf0j/TTeERQLbWr0
6PbHymlNeZNKgIzgtWonZA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5104 )
`pragma protect data_block
evnpuLgAjBleejzLpifZwq3/JUKxSZlzR4RMyN9uE6uNGMFgo301bimDEH3FOiOx
yIaL52t5JHZVcVu2SxqTPCDxeddRYCzh4UwnFVRdLW1ky4TFXrmmlF1wWCOf2n8h
xn3jjM0xbGbvQoZ8FyHPhdkAummKYSBgHRJP+OrMFF/1FTGnkNC+j72vbg6YXKGI
nRhj+RLAmtg+arSnpmFBPehkQLbvqpk5vK0n7dlozN0fk1dZcG9O13faux4DPYF/
5zt0qtnL6AJMiLHe9Qe8gU0SJ6NojB+La7dt0vS9KK8cPvBLKZBQFZYY6HK0apxD
ba9lpH2ZDiSIO+QHWWpKjrho9+g+iDGW2nlAx770hPAQ//cd4tOuIT3NoGy9sk8K
Ch0xWzHL+jiDpxiOcCd35WiGiMrjYTGdL/qqsnxR87QdzLgoXasd1m1W52m6Insm
FyoDG4lKHnDju1EDlAuPApVjw4DmzaicNj8EhH1TCAVZdXYECxS7NGqFP7jPbSzY
95GlTaqnW6HmaUsyDo5OBRFK5SkL15kh2icojodz0CVfo/EDUy7JZZ4iSfOqfsBv
DCpP0817JVpgEfRtVN+iaZFDjdJyy2EwtsTOZ/HkQ1HP/mjkZwrwz4OYwnyh7CeA
QcOfxs2mNDs+bon1jS1w7v9CJD4eAK/++Z21oU8VrFrxYiPE/bkJQiQLV0aXxV0Q
zpRxhN644jEh7SBfz1auy+vU9NHzXhM73pbGUmDHltakAqJA9PtmylXF4i/HiHZ4
2AHUagRzwyXO22y7OCc5qW+Nd6fGE9vopgTeVMNLVhJl86M5bVqB+JwprpaEt2ot
q52R0JxVBPyuaqCwotmNRKFA4ZUxRc2MPgIC+g8Tnas+CXnA5mC+LGwyFxw4n8/f
ojcJO4ACln+aZah3izFUp9CMQg6bYYYrUoaVcrz9e9cujOOQIKWilwccPdpEWKzZ
zk/eeMVxkiFgWMM9jBuW41KCNIcv2CBaYtMcgAYsfG7craioBDePSIRUffW+rZDW
OZlUD1oFlV+gqoFM6f22RmXddzS3Jto8P25IlP1D0NZkBOMyqyEv8KGP45zKChls
6JjrmVLXjKTfG/GdTvd75bvlgmmIr520DtYWJtnH42Yh7WTiwGecI+JRHjwi7HkQ
F6wzWm3S6AJ9pFueiB71yJyBf7Gb3HWbH7uu1P+C2/gvucnWveYINsCWFNFBdg8M
akt+oIb7ItKTktcHHrYowiKx6KffAGK1ttOkmC8uJRo1OuyHVVJbt0I/ZobVC5MZ
GVkehKj6nflJ3EuJF78lydRwlZIJwi+m/AkFP/QI/Zt+UPsQLFNbscNzYKlsUsrb
5SxjMU+ms/NAO6UvNheNE25QtBt6VYxyUzhAJSO6KfBoFGlNl1z8sHGNDxZXzSHc
EM49nLalQRBpOVVmfmA4H9C92Dy8Cxfy8+xn9/oQZBk/TIAA1M2bX4oxWK2CEXnT
gCgpXzODWi2NXqtP/PGu7chmGOP5Nk9mX40r7h2S165wwY+jocOxXpauToGn0cKV
XBMvHqCqLF8PDOwPjkRpc02Pzsi/pzyJkYdfCTqYs2maYjiYeGC50SrgJDne5uhj
E0sDzu4ODnR9dJMiiOdMS8utah5nMO99AUW6w/aEO5BlPqkCPe0Gcx0Wynhiv6eR
8P93eMK+aHZ0H+FAqQZ1xKjnTPdzuRj8GqF1UnC6eO93NIPPLz/vrnr4N3si1Vm+
sKl072L9vgYRoKay2CqRCQd8B92X7Lm/k31HAuTv7dWpFZZJ81cZ3vmVB7hXGB8k
UG0hwcds8mw/B5xTg0MsqrC6jyZ5ikS6PepgsoBWX0N9KLXQV3CcF5qZVUh6A5xe
mC4o/r4d5TGNG9HMNFOB58oMVxZAyVchLEaKWvcFP1dITHlbQx9uUiCNN8dqq6Q+
gX+WTcVcUB4haI3e4voooR5y9nm5Wg/96FcSuZBoMWrWDrHth9dc8TWGH/OuNm2v
hPSh+o5lxJTcmmcsDIapw8n+OFKLE/9XcIkAkr7WUUqB4sHNBceXAK6D5Y4Kg1vQ
KPQV7AXL44Odfif2COeSjelE4AXGsWXleUU34H6jzc82zAoZ8q7SNG0iA/2GYF2F
rQbqUGHugYmyLfUQdY7UGjZeJL7cTWRpD11sQyeQqhOu1eqmuh5qyLA7IpNlQYWf
YvM8KoiLShKXCo1jL//c6AA2y2EbCLqb+aZ7sDq6zj3Qz4H2R4pS6091kslMxEBm
0lvsc6oZawGLKwJOSlDLl3R3bX4sXqbbN/j6dpQsVV/tCl4l7uWuqBETF/6PfkEa
dO0v5dQ8PBm3bp1GrJgoxB2M2SxjLHT6wXbPXxrNgOhW7kc8Koj+dli8I23XWP8d
PdovSpIBwC8olFiWwGfyELCVt0fLyAJpF4d+mmibm5vyFBUfKqn9R3g0/89D37uH
0tMacA4H9QS4IG8iD1frg+W2OFXkyKm6Wl7sGIZwkt9hh57uG9p7RWlOxedjlENM
CY7Maj0N3TUnO4/4cDwIMilZYeWn40ZYA4IZzqNcxJux5JHaNl05xfdn1lR4IFX5
JwygNXOPcbwVze2m9VHX1y6crDZFdu00WTRLJs9Aiwbp5T3pkaw7garUSfxDOS8/
qqBMpDw8p4mkSnyAZhpVVWgq0Cj7ZQfexspmjnKH3reFgTOkHr+e12OTBJytWlPe
gm70stliyD8SpD0d18PCZJBK4d0w+oIY9DZ3U30ee7828y/eJ+6eO2//+h9/eqel
BepO4rPWRvcsvcSexh5dpfSlcWJfHN2DwxjuApI2fotw0Uaa48s3557USJUQucd8
lN7grfGU0S0CUEs8miJ95uMOWH55guA+Gt+1cKkftk22Oi3WM4eNMylNek7LrzV5
0/gBEhNDRvZxBQv7H73RqW4F95ioFldivgE8VhyJDkXRkgl7Kr8X5gz3cXlc2Q69
vrbk5OePvvYGtmfiHVcbXMKTuxpyn0UhWN7IBSskVFmFPu6mtcobKcHWR/4JI6ZS
htVIJU8J+8DuPY/NtlD2kMxz7ijjS9sXKYdK+dTAtEmK/ZEn5XShMj01xZdmGQ+m
qlzbHMH0X4mbiP7nYzlyqTX9f+6dYjU2XhUYBxxyHThWPbAuls+36rbsD9YIIVGq
TRUE6FDI67nexcSP8lg500d+BoAhBq5uuU1QIJo0RixrvcyFzykYYOdxMfxIhO2O
kVxI9Kn8PFO5Afn0VMbxxthBoTP7C3mjGRWs5Wl1C6K57bEfyc5QEFs6usnOoyUz
xH55qdoXls79pTcetoDduA+0mwoDKxGNWYbGKVcNQNEQy4Cri1r0uAMMuJMcVbk/
gZPeHs3kG4e5PI8toRxocOcp1I4SOApiRbHw9ol3A6RVv8yoYQv/dCGxoYNXi9rR
AKta9wtKXMrnEAxk8gsiB79RmajAwHVH77KTlWl+imQGlF7SbkN9DU+82Hbg/DrW
y7Pb+kiunoxCdRejs9TwTmXyXfag9xt9glJl1oMKS+Wbzc4+OA9bzWGWY9quyGUF
YMcPt5sa7E1HuftakocinWCaVeAdmJEcflllScXT2ZHJbpQa+Q3edrTGRHIVwrFw
odecIhhj/ON9wUVrp/IXQV7QZvIOfYAdQMCJhGulGc74xn8pVzBPg0va2AM4HQES
coH38hnKzKaZZAhrqSuM5ZP/LycA6ACVkyWRjFuMosk9pMuapPyX912YSKj0PKze
sNePTw2xNXUwb7Ulf6DiAvkNgDbRHXO/i/5/UGvmQtEFrraNVlCJj5NPptA3eBNy
XLVGxxhUEjj06KRD9n9R3CCnE7vBSCAegeCTphW9++uuO5ufsB0J6sP/GyCxP9eh
lTjhFwEjNe1cLesOGiyHo/gUqsZ++XQIurTue8qCqbpUyHwcNcxGf/zIJctWUu/i
U5XKc/GbGLYQy7G8WazO4tjPxn60RN/svYaFvB7gkWmD8Tfl4JpMNtKXWcZj1KjD
Nl79dMEZWm1Kc/5BshpR+YsfSwTscuuaSUlOKCXUN0vxOuaU1acbRJujIiIJq0gE
im1rHG2BGY/B/VWYUt0OGZL7bJyX5FewFj8toLZ7GyGeKa5XFIvEyquiGmUFFkka
dPM8t0d5b2ugTt2jZO/m7IkeCUD4eQ/EILZXA8yNYog/8VxReJ/tJNd1njkH8GBc
G1kavTlnF+AhfZ4POSYFzyU65d3Dl6YhKciDsR/PAjaCFKz3FO8AiqUdRx1YKdx0
2Yj5wKXHJrdqCGSU+8o4OkpxFvdtQO+nJ1JSSASrZIcauNvutTg036u4RP8iodfj
Fh53yEqvlhJQ0AEEkdG+Tkk8bBG6W86Jtw6szeuSy2iyF42CG+UivtL4lV438YAb
lxvfpc9z0sn0AqwWcoi8QpYyKcViLaDzzINcLxkz9StUR5eEjGvygvsqAmoqSXwG
XKk3QwlAHNbhuIjR7c6FHjxJ/2o9bxvg11VieN2acsPxBBeiHgA5fmywervVrnI+
kmvABtVKPQ9f3LL+UDQ/XEuqRcrHxjsdGFnVS8pjCn3ZqzzTqXa+rYJQ6ScAV7UN
iHEDOKCYQCNPLzFVPBDbI2aEl9pHY2zoZqSd5ssl6/8C7NfAygyITrubQdABxieW
MozPlQqoP8SgTIGgLFVGWnkFgd+8CulFKq3WFZxoN1Fpkzuuzby+BpTF6Fnhtt4e
XaiNetLElThdL7mgHuFkTNWmoYB1w0hE2mnadWX1wxCP4z5V/s+mGFYMHTDCXcVH
jbV7DJXFYxS3vUxSc6i44Vz42WFkPmjeQNhwziJBB816eMYz+qM1qbD6LeIeKIoN
NSE0ACAaEvElFUtpNXsz19+a4uPwec6v7y/O49b1p+hm94dJ13r4gEAm5zx6Puz3
ZxvV3rPJSRaxaHrfgakkAnmfAxj5Nc2kDT+WdGRbANRd/QqoGGpBYr4t9HjQgMbO
L2oOzyayIzsG+GthnuN0xMx7XdkkLQH0snbIHDyugq0+RHp/B6dNcIftbfYcTqGg
9v1ue5K5UFjjZEUFmrKA+xcRf/Vgmvz+cT9BgyEwkIiwMg4d53j2CNv4KgtjhRkR
GYUO9vG6hJM9wlvLgZEsuJIJ42rhrPm9ZUT/rEJbYvOvVNELlqKsuiGjUEK07RCY
GUaeeu1Y3D8pb15Yx3RK45Aos9MgSRy7kexARv/H2wnhA0r8hmn7nf+hWOu6hkMn
Hga5LirE9ygEwFePZTe9uyUCVAK87XJxgFCFfC0t21gF3L4ALGDbTdV3d3bBXwtf
wPnCbSJufrCAs+3WpL5K/AZt26DwotTA3VlQjtUNutENYJaZzl3WVEhuE65pVhsA
5V7oShMihbT96lQPT/ytMzKHFeiKfEfuLlLkFT1rzXUbn9FFGE1FzeX28zEJL1rl
+hzIjVzcsbIqqWEiwwFU7zfXhIz3LjHHiu787EOXPE5z18883CduLEZdTRBN1Euw
2DqE1lEz8l1XYJazX54y1xwSccsRiVAjxKDGyvWy3Jm2PTMdeac6ziFXA4YWHuq+
jUv7EnVP+VCksbiz1iCA50eFTKi+8eI2aCTeguzsJprPdw7kfctYIa8uc2L1RafC
9g1Qjw/1CA3f02OWK/wW2xbpV0qzMTEPyU7Y98KJjaJCvSdAJ3TSkBtbDna/y/aN
LxvB9peAAiDWDqnEfG8dWaK+P75uoklwOOtuHcxJyV4vXfamM9AP8j/QmJtsJ31+
hJElWmQf1vdJBPuw02/HOxJnJZRDXWJPzCZQuNJZ0n4yilbfgiMuhYzMPdO8kICQ
6yjrZJiQoQLCrvw8PnDE7nQ6TL/8DU/RVVYIitI7gKi9KiFaUMvBPXn9xMgjNa/A
ELj14xZh+2pBfI8dodEFJkQvuVnIz+ds9igjL7etrRfNV1poeMjI11Zwo6SKK2Pl
BLwK0GffgQRwP09aYvPQiTJAYr2t47OkeYiKk3lh6ja6DuKjCzdQUBML4Q4OrQOx
TbXnC5HbylpJyRwaTchSU0geUa4J0Q0Qqt/q7miJKn7Pc/SWt6JQYr7nJHjWLPLM
+hmzkqnK+dMFYdyDEV3VuITIldkBDW2J9LR8mcrmnvZIANiIZQDmw7Rnl1bcaiyW
ITo96AcjTV8fOFKsfWKTRGVBjqR/kKaFwNCXDA30WxYQpB9Scjy4z7uGHwHLyskQ
+XnyKsj59ZXNw3soRa2YM5XgrYFHOt175m1LDDWoT5MEkn22v8xwgABvOkf7WihI
X2HnCIRyXKbYK+Qtn4N1Q8EH6knBF8eZ4zE/k9Jl9CQOOy41P8cLpKOXxUGOgHEI
LF/mCLs8I86qfPfktS+8pADcKvwKnGm40sFubfq4Kn8aalSxNsqc1zOh2rE4mMo4
IR+m4GZ4ZmZevXW+HA7XgslplbolOraIZ47GLbl65TVb7uP3FLtJszZI7QXISnMa
3uu8D17hZ4d0QT08oyPinUy6r9pKm7HuSTt/e99/BcxvT1mueTAi8CX4xUaJAVKj
9956awCCCaahNHF4GHJEe6P2CcK2H1jneEZ4cM1znASji8tv6CGUNl5OYimcK3D/
FH3w/YlX/64m9j5i8KweogGrGamQESri8L8gPMH0ZXXiDbFd0+EegR4dYiwcuG3I
+YY4xcU2kFsWCNiModUqhdR9ZZ07OTcWbX1t1xWoM7ss0bgGPmDccN20bxiXHxJg
/oy1pQ6eJPPKUyr+4NFQ9mn6qi/U4zwXCgmdnoqnS5cGMxDatxJrwubxEyYm/aon
9YDl32AVYopb8Xda5+28c0Np6f9QGQzvoUhhjYvtF6i908LcXvWXi9nWU9qDeZUZ
k92jkUAJ93MDNghXEN/liA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ikLcZitpxDt1VrkiLFksuhb+oOKQ2AVeNwF/ZBA1vTles7fYGXvsRy/c9nB3oPcX
KG3bGqtdn6UtC7ANafolAqjP+w5TexIL6ql4qK9p8bhRcMH/AVzanTd0QirLZtFv
9s5vNyZrR8shGtmtSYQICodlZ/jd7KP4ZFsO21GdnEhP8gHF0Um6DJyONP7AWYHs
+cPQA+SHtt22vGw6npU18V4YoDw8AVRROnVEJkPLFCGSbhXSsqsFGuMVJHKxbjZL
ILOpEOGlSXFomkkwnZxtqcqDDRcekfHF725OGZzk2OhMbhHZ2fT0eY0dceXM7H2R
GPc/cRDwOn0lAF6/25mpIA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2624 )
`pragma protect data_block
9aoezluQbZPJJ0dM/sWIqg/aI6wl2F65FS0RiCBSV0i7HTGlbN/roxPFXvFfd9CZ
vkWzXbf6LCEPgVXzADOsC7HCDqqTN5xS5iMZ7nK2xxOoKalsqBji9kTqVu/70KV0
ZPj/rCyaR9zBJmZecyMAkhtqCvYNheSlQ+8MzEkJuEQIF/pZvny43fH2LGDxu0mT
2+19iJLuXioHuGsYYog4XGABAHVXcOZqCTDsgY7t11HZC19oiMiqYM5Oh5Nt8+rH
s6w0WSFO2YAt8lCClizBxBB42WU8QXmQORyUbh/kfOs7K7fGjr22SHnAdkyJ8tXa
Sp4wNpYo3bK6GWuqqiIDb4jdK5e+FryDEyUpaTqNVHiKn8qAsbSlGRuN2XfvFjyr
t78CzLDdUSNEox2PBhyc4Fl7Z9Yll2zq9a1IdUSA+w5B1DR5MK4i6CBfFUCX5UKQ
dUCqoV+/F6QyLIXkTZyxpI6XhhSvTpGNQ2+32/Q1mtuBRoReWdgKqD2NwWelo78F
n6QmqZIiQSec40E0FYQbdxN2lItAjkPkYby8u/dPv7X+8TQa9wq/hge84rmjz0un
B9AVtSzPZ85e85hNeUeA2jFtn54T/ML2ZIKWmr494l2830jBmHn224ojNWXuwrJg
qZ9i3ztLHagriyL7SbI/gah8EOb9GQjYyTQP4Y88liJEJ9ddP5X4jUHMxuDm/D6I
4cvf9G2AYWR5NhEKb2+Pfff2hbQKG0lDK1dgYUfzO41+wxi8z9M6NbZwdcN7Nm8r
tiAUxDbzt4n4y9HiQQSeWmOip6i8B0xsX8AVA7x04+wdNYNSVHurFTq5TkZvnB1S
OoC57Tv7m8yOya5uxptQuIVYK3mZtrg1ZbFViiSddZZCnwcX5Gv0LKekiKg1FmSO
fHvlMzHUc19Ba8VsFPrNaICPLO8HIEcVpEM9Pqwcxvag3iy/A2nUkJhDft6tySgb
0kXcDE/Iecyk+i97izkVDqZWLE0qc++cTaG8WccFdMMDsALF0QdGqpgMd1Bg2VWS
vSdBYEhHBOVujDTk8rTGtoRpwUrf9YSdZR+exHVn2b0M7+AqPNVVy2WoZz0RPvKY
UNX+AnF1Bv2olawTA7aJo9GyjZanumThePnqBVY1q47h/NemNCa/D5D0bVV1eLju
OkUU+oXGZpZoycXwXVpuQPYnMnO5ZnQ90wkiiqI5nd+53pz220J6If1f/j2MsKJl
RC/XvXtpLEqT3F+YKUyIX+uNXhjliBLmSRaqs2HxkmSuRzfzVu5bjT1Pj+XROn6m
bHuTwFAXYKnvZa10LjZ1q5+sq2UIlpbgR7yj/yRs4airPYmiHv0p3KweArL1fAPI
1iTwkA0b+4ArevttUatt/OgVHqsSPQwwbs1R3UObbUQZnV7djR8hcWS7xIEW3+I+
Klvsvlj1QAitF/eNk/sngahLFH4iyekcZcxhvq8KA73NeKDiLG0U05SKZ/L074Os
XI9JCUOqmccW0+U0ixvGjmKuDfs8bJQ8eHotOreHCtPVXhtoBEsqgCIlFijeLV44
Pf1EhbD51Dm3nTQYJIJOBpC2moxbna2d0l0U4HWy2TvL5y27f5ToRch19amjdEmC
PdZ4ga+HT9VZe2oMVHyOv7i5aUm7sPq98QW7cSYVWkp+ip8j1w9jvkdydshhN17G
XmY1+xvD85Rma7uLJryc4xfVoaeCzVQ0V71WhVWlSuRbC9ESY09BdJFJDfTsDzHx
SuzS86YcL9Tq2BstztcW/6qA1v1YLo3DoueJo6S7hPDspNRZqFPIKNwdBcupGKLo
GdzyFun9JNiVTjfduIQSvxc9EmW7YB/YS64kIz0I2XrGVpG7TWz8hqBpMSZWCfRv
Lvu+N+Gi35QK48kr3enToDQuRDGQz8Nv8eNCeQMwPbdzZq3+3I5JPDsLPDotQU0V
dfGyZXHU1PY6TZnrHpm3lRWRYrKAvNJ332kYCXtE9yeoj1ylRR6kCnSobbLZCou/
otKFiUD/S5xRrcROD9eljyGaKRdPg0rH9zpiwajCcBvODs9GSOS+KsgTt80emuOZ
ReLZ1pIzUxbya8xSe7sMy4IR5yXZfO6WUtv7EpNoND97EF1XUs+sBGcwF490yPGe
O+DPC06WziEwQ2yVa5k6d2PWOHvFmAmNTb1uUeQ4XBKo1gCj3GqXRdqYSawlq2ox
Kt6DyVJgSStoY22nJrVhytLJg4/l2MTdPKm+lEmg7PT+z70TUJP7Dqw49bAdH/z3
Nlbw80A6N9m6ZhS5OrPmLqsJmgUpmIrE/Zt8sLt9u/4Tsb+5M4xodX+tBH7uU7Yh
GvMIHmqksEu+dAOAmfbBJHE1c8BaBta0vU2saegURFLlaoKuteaDbNwxjAdLJ39R
pdRn4bibZNokfSOCYLpO+6QSMhXPWJwSpZC2PnaOErQ9NenmIwuLKgDYqAJwns+N
Y7SXG/ecO0HeGyvqlgOnqukSTnGf1mjWd8BfDp1rFqWTZqmuBcCWk+n9hR/eFwm6
3821wheRA6Y/FQAZIVJvDYn/HkbmU2y3pN1wCNJNr8QttrkcGkdr1tDJioif5YG3
BGwbSbpNS4njJww/oI0KvPBlolCrNM7jrbS7AaNgAAhKFjTjjYbut7jYl0gpNM6L
C8MrpJAQvJfdWTQlagxBN05cdc3hHilxsQEVWMLpF/4U05y7ERa/SF44tIMPLt19
vmxb++swR7z3UXAFdPtlHs8TssCHllcwuITHZIt5CGD73qYV+/JvIe6EcS+uIWE5
wGBBIlGLpyTrNhUe5VUnJdUu74D5N4zpIYCAhdo5gsa+ugaakU0mzge6gE6M89y3
5eUgy8vkC0Z4sr7cygzsoHXV7KAfdPHKplS1UtAIc/wpF7Q3EWhIlZ8HahMw3yTb
1g2YS3+mpJ0jPCbrC4lMyIJh9iqDqL0lNL/VoYOdc4Jvn1VSYTJwATMmd6XN2g4q
ddpXIThQV3rDht3uQDTJiZ12+xOZRB9cQRlsy24USj6w8+GpKr1v78RZFR6rE/ch
qj6XWjjnoXCwzutvAivm2nUZDkfKpRX8YKdCxKhS8HQfqpo4TXkRdQ0ONLCGZTkZ
q883+2NRubJPgE1AGF/1P7m0RSuLJcVD6vgz75kS9mIPzOVrUHWoQW2AgRbc6tNQ
lbdY5p0eXn6SKOBHQ3s1/2c8VSd0jejac4Z2YCRButAYJOTZE8li/cmNgBE0FbiN
7aM0/f3xvM5Vae+sajinoSvdd7HxxgVDuti8HvkvrkzRZ7DLfph24nq21qeBC+rW
eGKxwNWYXCc65A+eLUjsOUKsxie/fkOQLK9z2/FdbV558EFevB3okTz2gSKzGpfA
dG/BBXA+UJRsq16JU0VRKtoGU3/65H639mxojIX3EPvNmBK5wR1Ltxb2tLwniD6Y
ZtwaowvNXyjg6kw/ilHTbot4MJ05EnvWdsaFavla/XAcV7/sbIEGp0vU7Jmf4Wrx
AkmgPfODkhvebmfDyEoh2xkbT0Sz5gw5D0IDZUR3TJI=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
iOCGh9qPi3WTUB26ZEbsOyBEsr8sD+bdPyYukU0Px4RtFdN/O8zX/HLYec2q/zP7
xWST+4+7WZ3YnkS9vnKWuQAUKMA1UPzOfouJNVlpF2v3JrlNMPfbevcBCur8M6fL
5pHW7+c0zSkvVcO9s++HBhX8t9S/VK7joqY09+ejulXnYLkOYsDdficoGW9jDaP4
ZJDPyAeD9OD1E/aU58FusnjLkI8PTl8CCFjlQiL3eTD7olZOqG7h6PGGuNgFwItr
RSwxJIq6XhtiNSe1r9AVqa/mob1mF8++tHWK9N/x77xVzoAs2m+Czr+6iZm33f8V
jb5Osg3vipY9C2kYx62cBA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17824 )
`pragma protect data_block
B7G4Js5rUBuvDSBCHnWz9zXmIblRcfPltRm7dpARQ3lLD3SzPtTpzsM/EclZm7Lc
aeUFYozUsupJaoXO7nykCARWz43+Y4oOr50u1fYfonRTEMPm7VEnGILCzpMJ1Awu
5vmJ7HqrqYvSEAqTNZNMcZw65szXV+a3N8kS+8ILAsjkOLEP3s2Ldp4RK+/rOOjf
9FUywAlulh/99yRWIJ4F1xZEm6acaiPbLkiEfPuRB70OWIIrF4QurdAVC/BXmtTo
3+CeVQG0ks7cAOX7Rcgohf5iDKP/3ECXQPWRAboXtHooBQ95E/55X+5zXm18fqCs
xVZaKf2oY2KrFDcsjkGCf3Vd32fWbvyGKJQnxs1fY2115DJLz8BDjmhFBNAF39LY
fcTLNmwMrCDVMcGEcOBZStT5+6Fmfq53U8GkNzYwX+RJfXTqv1xIl1dZ9iJqgKfN
39t+dvmq4MKr+IjPNxcAkM5ts9UdZQt+o84jTedL4DyzyrzN0KZ88ejrG0tpOLOw
btnUHlAtnvQBBq7Yxe112HrwfLdBxaXae1DA3uxDYRDW7x4kynM69LFnHMcU3xFo
Ub1JxJ/89HdT7E4HmbdfapQblmJ9NVzoRx/JxxDnazX3wo0qdchNSa2Mlhuqfd/A
qE5DbUG5p8kdIr6tzoTeIJiR2F6uxYC2Pff1fsQxP9wx0pNFMYKLL7IB9P1Y+HgZ
9VdWedzrIO1F8oJHaHEiIpwgUbSURXDkYFajqJTFncJfYYoYfbNAO8UgTAGBnHNe
UXgZmRr5huPcK+6X7OsqbRmnyjiP50UrkaXnu7v5atkOoGCOCwYNzCahFnmzkJq5
sEgZn9pNGiVd1aGG3uK30T6vbum/ItUMkoo99Bb9FlQWpzkN4biU6rde/vw6BhA/
w3ucMhlyYPDMpH4IWIl9etjpKPz1IjGX1O6l0UwitLLSxNBp2VDOORHbLVOIPLrt
+Ir3gXWmR2r1yLzDnCidgo+3A75TErG7bZvbLBmKi1SycqIZkDEX1sLdRSBESgpg
YQtYH3u3HY0z2qHL3rIppmYJUCq5i/0T0ueP/lp+EBAMo9HAkw/m46AP192uBBhN
ngTAn40104ZVDuYLriZaRKVbJ0byj8KL0v2wmRIpnP7JkbpD4C0DuZDWB8DwXsmA
VEKFH9sgErROQgwh3w444B0D2Oasb6m2S8bBz3Gsf2+XHCMCykzzXOlLLuYSjhkr
w1lZusqCNWkAOChQFe2WC3lx/qQaHBGcTYMffO/sLaJH7HyUkR7fupTv0DL0uKcR
xfJjPsZZCae/kLGB0/RXAfqFWI16emMCsm8+mc6sEVBAGh3WDLfmjcKWLSx+8sd+
oj42nUtSZKddj++nj0BaUT02ur1hKXWOfWAL0zR5KSBQ/qFEMjP6L4UWMmjnCyNb
/JgaRyDhI9FZncN5RQ65YB3uxWFMk230hK0PAmJiFgUziVjTti9ZcqmN/Vy4Btgx
V60AuH5qEKkcHcKk3hpH2XWT7pbDISdrdRiS4f3+8odTM9PhfRdP4YALznvA5gX9
H4odlWG97auTOTto35zNwwiL8kAngbILbgElo2kh6vSM6uzJPaCTRX3Oo8NNGh5S
mjl02XpCC+qYIcaLsQgHGiDRdo9XbDMGT4Bbe6KUQ8fi5N295GyDpFSYDF1T3dxU
tZfye1BmMuaW8kXgE2xwWCr5AF1NySpRqqUY/LvUOBaVzFslL79nOow1ypXrUai9
9Xt64haK1tZsKaHJoWnxOERhQad40SdwWPgPt/+53SqY6gRqTlqs4nfLdSsOPQ9S
p5XPYlsO3hC6OY7VTnX/PkYs5jbFcfvBdeZqsCfTx0AU+1Rk8i9jZZTiC9PA4y82
kRikVcuLBHLiHMvV/Rf/G2CzmknaF60wyKlt7+JWOJDDsxBuDilaMKGF233HI8/d
oW/pvJ8s1PsadhW62iz0bJv3d6orA7aCQc0jXhWn463rseo98gyRQumUvK4xWPlB
4tAoFYAitym7ngtj3VGljRQgejzzsQ6soQIor6bf1EzQ/8ifyJVUIYevYh40kw1x
ak1dG06nh4yuEuiSa7mub8FD88PtnXEBgrqDSP1P/GlBd8eFs852mzkQyKtbUnVF
3E09cTvmeyCShiXYTXGIgxopHWgXL9aodgBjD4lv2EgPcw+uGbe3twgkBH3VocDq
NdQ+pAhFMQKQK2WsuPxfdtXE3sAe8UZ8m4oH3wRvmXEIegd0WT2QYB1hoOI1Qd7M
oBrDWjCis1FVibdQ7dD5YlfqZNyvacG1CqbUKZrLmV7jk+8tIQPOrHnNPKrltpe5
ZD5ltZfHF/ILctDA+M5z5Uhe6kRhM4EIuiMf79v2ERKJXt8LxCp5Iplz7dM7SAaR
zwgXUkYJIP6SJ+Hov5hVGdtnmr6BCqDIL4Sb7dgkyMSxISr14Q2JuvS5VLcJmfMP
rK2GS/HmEnZKnJtooqor9HcHkF7u904eM9nj2BAQdWuD3z5taoBuSbsXX5EagBRc
guM0YquEADPWP005QP5v8m1rBjhFY5W7offpNFaCM37oDxAxIkI5QoOLOgN8RUd1
shGhm5ctsEErV0+uYLhEh2lu/DfcQbzmGcl5MSzRSLzHPwDxI/n/+NCPLpcBb+nV
MaUy2Oe9Cg3oeqbA3Gpzx+9FbVEksVT8U6GoUXV7Zf2HrQN0+sy2ZEcWYQFqh+mt
t61Zwt2y5V6d8jrJ1DHdoCgKKAbQuFQSmumhGzJfPVeUewAgiaSWeIguxOSHqeY4
EkbPSauo2MT0ytre0dv+1dpyrp2IOUdzpn33w5MiD5jO1Ef9l/E82b/nry2sdRQm
NjiaK4le2cfYh8omGsg7T4ffrvPy47VyuvTL/M4d7vI+NjGvRF0xYlhOCcyUcA4x
w4OEiU+EUUIXJO56zRtP/o/oh5fQz9JwtdbrSbHVGBwvWJOPUIEa+QaFYybMLxmw
2HYfkbB5LrXs8QX+EQ6csSGTs5xpU1Nwo6ksBXbUjy/C+XQmLq562xyklAfung/v
K8diqVRnGAyW2xkHgy4lfIa2pNKNHdmDE88GZP7573sspOBC9m6w2g19Ugk/ljli
ZEY9eVI0C50LaUS2Of7TYQnhzzpJ1/ngB/BzdWgfp96cyDfDIAB/zW1rBUaRvYxI
PVQlnOm/AC4qSxZ4uLgWOBUZMtIULWvLdcRPq5H677vAscRX4gjt9At8TAoTBNKG
EUPUdE+ImHzMKnWzMJ8ja96nXoGbCHGMsoITT06mucba0nrPrcZZbggnE8VKj9Ve
ybtpNd1KHhtzWX8bprfgS+Qt2iTXxoHH9sLuRp8xZC4xcSkIobSd34XZmDyIzeBj
A9w8I4qnKVudhsUm4s6mCZdF+MiAbfZl1SoImY6UjsXqG8xjQ6e0KM4RWj3Lf6zH
BWzrDAcyiUgOuXLLzW4zp3ZsRsnk6OaSEKpx3Qw/NqAfpDHNMwJcyydZhYEhJRgp
9LkjD36hh2Dka/5XBdrBMdVXg4/P5N18zJ8XBtRx4kHpUs7XGW2RJCnw2VFUor7G
QpYvenO1YhHaAzn9wjl3ErMO4IlOIBX7ukH2G1CoPX3HMRetovdBjXGrV9z0cbEP
IccBte/QbpSFaCAr+3Z62eCaE66TRaBYLvIOjq91nHOrnSr/FhDkmyDcWHUNcTb7
bs4ePxtzy/NTUmW0tnMIIbeTfSN8uERX4cMr6/4Mgwp5bAGrwPuU+BnYRYu27nJP
8pDctt6ioUBBaWt3zfMXi3tfLwzKzNxF2pDu+j8a7NT7J42U6tyewsdTnToayMYG
dam+nuIU+q5w/p/AVhkMpql4jJGEybxRDGo/aT9bdzBZahdqFelWJjDfCgkKaQ2C
+83qQk3de1DgK8a4osttIWlvLFl1SepUlv4GZC6sX1RQ5m2RTReEiSi7YWxmS1RI
x52E2o7yzVqCX+isHl0rUU5mOi+gvVFnmN2V3JxWNRX1iXKiA1QAbue5xltp7rqn
9n9/KjRZ39Iq5YN8OH8fcPl6HAf1hp0HTy2QN1axO/lEjgCefGUbrSrlBwMjqixb
RPpNqCjgEdXrmWr54FsmRfK7J5y9/UnBxMcTlTDiXYY1xfbH4gogRVhBDZai02Qq
TFFECtIaupc2bR/tSCpF3cUpYniPZFeaIP6u+DFMqLquzCmuuD2ZDE5dvHxHq0o2
sog5fMr9P4qoWbcDo1JDyPSU62JV6ia3bXIiaesCEreShs63aha9P6yFQTFP+o+f
yWMh9/YM6Y95YaXC/NQOqcCkSugLTI7TpsgdeqIhOsQCpERJW73MTmk2Gpi15HeO
HWkvO+4QBVzhqtkKG5Xw22GpPfJY0t3K1onbjdE2bjq+mK6pVz6TPaMzcGpvzILG
+FMFFjSfgyXkDUOEPc5Q4FSTQ7hVpJuIFDq5Rc6jcQ77sFosnv2m3ZxJMvwgpn63
6lqw7aKpOanUkU48LyxAnan78UPTU+8FuwmBm1dE99IQcdOBGf0/GzgW0GgnA0M0
5QzzX2swVJaJS7WICJlisVqb9qg6XFlXEGa2xccZzEUlF9py24vK27oE1sQvLFkd
IIdNaEmWWsCYVxTKoJXgxPYPtIAj+LV4KpwomyZ+9HC9cnMivtdo+LoxOpN3bIjW
Rx48PxUO+iA5/4IyiEBVOzaG3h/D7OnHEA+vmfkqewRE0Q/2LSSg+ya8Y2m6rWDL
lXTQRcUlgcLfQjhcyN4RxuCPwklfe32AmTz3COxST6HaSFbQt+6NxeSVn+nuLDy+
gzLNxUwLeUZe3djIN868UffQMNHdaWTDixLnn7h7QvhlCWaFLzt6AC7ncjCfIWua
Mi/E6a4Eh0crrBvhZLyio9UGJ1RqPBtHtzavyM2N3qDWAk5qExhTfMbVwqmUSH/O
KJz2aqRqeesT0yBsQ2Iwagw1HxILFS9u8PB3A2j6PocOXmS7LbQICA3C+Rc4tAq7
zQMK4P9X6o4kcLLKvMEA5QbKubYXGKVFbNNhyrrDKkK/+1+s3hH+BFtHZMXAzobt
U3GxFfeAoQWAYedDoRc/ndvtnypopU2uXO5Z4Ts0fr4w+mhqV0UcQ99hLY2UxoY0
cLi4YhGursoBub+B7Efghp+QSOZ+UHx7fLcMGTh6bsTJLGFj7mBSWgzvByW/V8Bs
5nT2qsBoL638jKU5m9GKpCrTeb5glR2krPB+mUOJxFwDP11GN0wwdQuKua5IIOoz
sYBQBD+ra3VrlDRZqDIFnXuUsuO7fCQgjkbBV8xexW4QIIS5lG21Jykl+DZK0hIs
oqLKIvklqZO87be3pMaEEQyg24rzq1c7Il5yRenUWFVziSsZvSpNoDjhlAiPKmE7
cdpiWtEfbaYYuHibGbSIa+5QOfI9a6UWZ9KM4kAO2QhV0yBJirXikfy4/jmLEsdW
L1wobogtT4FYdjOaZdChfkwHu5VUrTaH2sek4CuH7kb9EtSSAF0XuIj4YDvDAfoN
+d3q+SwNnknoy5iNS4NLZ+Fy6A+59mu/wd0WddC2FvVuMluCXCyLclGRuYR/kXzG
uo6M5nCiwyuJTBYtqKeMz63IBp7tv2s2/tOfwxaWP24W5/IW9vggjk2NW1IpoODW
tTyh0D3jdY2GjP6wlgc/1fq3+BqlljaRKGLJNG0hF5factirilaOEIbltEO1WKe5
+VUGqmZlOMiKX3GkZRgtYL3CV7EIVcJQi33W7f5x4GHa5DJ3ZQcHsavvjbaPQde8
B5Ihyy9JDU79AETSEwk34Z5edbiNKGPTnj4LFuz+f0JMg0LI0REMC7Hf9HZ5bgEB
lzEsbMzfAjM+Z/21qUexmFZi5s2dL/ltM6BkmKi+btklp0AgozKXxPyBCMLQdEP3
9AGB2892n1B6y4z8lZhUuxZJbR+1vrjcBgOAjkAlqkGe5svqT4q8FspVb44c6Qa2
A5UkdUcJtb/vN7ZdxfvS/fai0+IsBVH/IxX6zxpIJwBK2g08blEeHbxjwY3HhNXJ
yMVWK0TL02MTOW3i1lnQX3zh3MxJGQ+FHMzF0veWNzWrV0IVKPfhIdIa9q7eOcVZ
Ux2Vj9ulBre8nCEfD7LoeD5lHKWJMBGC2VR2f5Sj1jB2U6awFvsuq+fc649SygsX
y5U9nKYO2fn62lPKo6NENFcmBhfTeGle6V5cpJQ2iZLRwd373TwjH+MQgffZm5kx
w5IO8fadckoja44oXgpMcZiuqbDSPgeGiR2nCH/axV41RhibmFHtLA2JpD4S2Ion
EoqtdGyGcWJg7zNMpQp8XDbha1pANGwAEcfS6YUfDLqw862bxWLBKzuxjkZmoyj/
2NLTzpIMuqljZl1oJWVYhOWvCrlQ6S90k8cweulvELkHxRAMrDpNoLO7fhe/28cE
civYVKbGq67RCvlnNH76MmRsJyEMwIdpVKkq9bSZ3Skbs6tFJH2q4ymDiVZEKf6K
DVNnLV+Spa8fdcZUk9hT/sCr0O17qIUsi+MQ3FeiNGQkDKdtDtUP4/Fwz6q2O7AV
BFlmMyfzr0gu7xamtqGZHkTIY6EK1fL86qVkJdjA2z9gzM74c/bbtG9zICAXGSVd
L7BuQjGoxxUOxjacUb0PIexX/zxEXXcOthc2hd1jqBH8tIEX/dApb408CVflZ1Sg
GdD05WQzRd8TTVj5nsxiQ2zwj2TJU5wonQ8ibUmFgOKb71njVIW+pvbTQHX8/jW2
RJuIVB78PUqgjbkjjTXjMEcVcNfNq8TgdE2NJu1a7anZ4oW9odWVkPjW6dCB7FmY
A/8XPaVjk5Wm2odecBrcUThFnFQNI/D4FoVG1X+VjZ8iJLKQugacZbvZJgnHbwwb
9RxVa/d+rtM6tCjfEl2gKf83CTVLn++3yDsGdv8Bq9cxPlIvRXjttYgVbk4KBVhB
8QoXtn8YaOMfbpH+MX8Eo4MtbgdbSvd0AignW5nKkHoKTyNbLOChj602xB+CQu/a
V26bNEE3MOJpkxyuOBjUnLh0ACsW9WSxAWDImiKVhP7FgAgVppgCzxDmUkxT+NNM
kA7gJdFOwwvG4NEwl7uak5wud2P165Z44LZeZ6mtJTR2RHE/L9M7Mpx4G1yhW5Rt
mRHOma+HUm4QizuMvESo74hqKmCrY79EbzB4H3NbR18x1S9EpNwSD0TAYVE7wnKd
QyD42laQtmc9qfqCkpQa6iFvRMEk9zGFh6PBZYipiYdAtnURLGTgXq9yI6MxGewe
r14/Xr9Sm+XJyhgJ9wzMXTztsMM4L4b2G1IMJm7ZIKcDKLf+j27tQ93VDjVlv98u
L5dp12Ry2VNkRSgsn1h+FsiTnFuK/yZr6ndB09/NLW7yJ4+Tfpl3h5pH01M9aRhm
bdEpZ8uYu7EWOIPTwTR7iTYPv1XTaxhececfTAqobHkZFjMD3FFVo359D2EaGFWs
iTo0hotu8pUH98an8bTog21mdEa+Jd0m3qb5C5qaMEACWDPdIhSeJfTLAmR2z+R4
evsfssClOWFjolFay3xTuZMRkJYvV7lETuBLVRAKaJx1IYAFQdo6WaxI4M9yp2wU
UQgielp0QXBLsX2IrJWWuOSP1JJ8r3FMAeMh4iKeYOZBZnbX9CQXJhOJtbh4dJwc
Vcf53YReZXkX5rE8o8klLESpp1eEye7QM8OMzYV/NN3qzYUNRdOaydfYkBg0QWxQ
19jhAqcgKmYSvQyr+MtcLdiYHLCaEOsceV7ozq75ur9GbkXH0c/CfCwFsg111zdq
IsTga05o8Nrd7NZLH3AyU8e81Z0HHHH8Gn1mXwoOKSapO3RkBMD2cL3S30NCM5Ye
JvwHtilX9zjLPeE7/C4af7O45Hqt7sw5xe8znIjBy+WkE9fZJq7sTcI2yllCEhR4
Fns8NlWF1mzzOn19g67cOCDCdJBhBFUOd6LC1dM1HizAljCv94WLfLKecHgnHBxR
R3ISVeadv+XCVv1CAGE0bmM6AFplb1DXWBO0Bt1+drVgs9tam4Ir67SOwWQzF6mD
x8xxCeQpe1F0GHJLT1C3dtAalGkG6flIc9Nd6Ra7LzMFoeFRmBEXWv/Eg7R1TS3g
N4cbWaK0p0Bi3v61B3YFcmETi3jBq++dhD1P01jap2tGdCPvb65ad05aaJVn0oss
JTrczltD4zpenFUwjT90g+gkQNjBesN9j2LpAf067VAH74DJFlsH0vfLCPK54Vfh
/Rt8Is5k2iw8WOLOUS+rDng4iHJz6LLfcdQOLJfnDiAhA+Ukmpg3WCxNdveGqe/W
NIhmLNelm4VDvJUPBgyHvOF8IJl0rafpdi+F/AJH9l5FLpQpz/xfMCi/O8T2Elr+
GL6WpwXzN3/KHgGCE6XeSF87GkFK3EstSCl+AahGUW4ZfT/F+EWfS+PVg8LQmyhG
Pov3jytbtZFnwlpvKHBm/gRWh35xXbEdALWx75LKoO6szE0B2gPuUK0ty7u2GjMj
1dn2jWZBiVdl16h5a3nGSRapwfGlAB2sDxDIpEfjlBdoFtB0LSddh5a+9ivw82MP
2y0P30u5caW8jIMRg6kKurp6ps3oEFxwKQKSzWqGG/DVnWXdBP0Jgj/1YvrMZTVm
d/Sky/pxGtNWb45bHQKBLGdWbwcYYGJ246KxFCpsr9puDWzDuG8ThVPZ8s4m+OpN
6FbuRmVoXyZUeLsKJfPSkqlOHj7WxPLxc+hifVi8lL42wNiq5JnzE4gU+M5qw9fD
mjFtRJl2wqMu+OFvPvEwanOVRjBLYiy/B0v9P6i5Z6N7F8vo2/e94FhgIpPXMq+F
BBQWHn8li+J75KKl9nTX8V892pRWArTakW55939jByYc/WE+dRHa5ZLeI/qdTMMe
QC5S7cfQaOAX9LLJDFUJ91TLG9BQnQcSiOZ0BWq1xq9IhDdOjfd7nkPvWMQtcfdC
3NcwMNkW7UA4Slojym7jbETNOZP6QuViC0GVFYG47uTyfmoqMrhJfLZmfImBq+z3
IY1uDjyV2QHVfSHz0jG/wktS2JAL6wnrcW/QIEuOH7ZvioWXVUYODUey3dkYv9V/
LPtenJ1MelAVNUBef8C7jKw8uJpsoam7Ybq8BM8O54X6z2SMitFj7Bj7+qBOQqe7
G67O6ptriahg8FR+nCmrgPFYBjtxdPgtWXemq04mYrgkG0aVPpeSxZA8vb51c9sT
Ot4CB3B5yrUL7mCYHiwx8R+4hkbJ33ItrWI8kJAv4TPjpAS6SVuXUKWt8FNec0li
G5j1xGwkLKrc+oqn1GmjohCmE5cYrnJK6usZlpwSgfE1GFMC+mng81qlZ3kXk1c1
Lu1bjhs3mOlocMcuvWJhSgqjN29mMDFUqt2ss5eUB9vvLEYq707NMX9c6IwxTEv+
gl83TFnb/9Yw16BkKupZ4lid8Qq7koFI7y0ZDUvfkwdVBUx5yBHT2RstbygT2upw
tHrjdeS5FxuzLFqihb3oySXUH20oyXNBsqGSdJICc8Rlw4SSfsnIhMZq2Ndkbl6s
Gn9UuUsAjajjmaCbfe+ltCZaEk73Dgbj7wnyoD+lRRGyWL0mLSdtYnVx9Jg6uj+r
ecknO9/Z9IQpkdR5OEa6b5yf786+rVHo03xrb7xd7rnoyrv5BUreNtR601XfmOm0
VsFhSdz5fZhUVxVD0ukPG8m7Qu/j9c08nJTCizlde9QS4bubXeJiIf0SsuuTtvjh
5UICt1KfJjuSJCqLQRrWkjkUx9SkX5Z/G6m4JARi4Zyr/gQAzwV5XT4Cia5mG0lQ
ReP9cYX5uppAgyMftGk6YLUaeplI92i94+YB33we+8gIbx5hTkP6wNxcPSzswuC0
gl9165Ck3pbunEwlIpWFP2r0qfVuRb3XNzgUga1D8vxACNiGVNhxuy6Q3GgjJzAD
mGNA+Se4bmkqypp01FhHCm0uduhke9fR/njtJUHh4I5tBjDc32XBX9sJBgqKTyyF
1g9SRXDCSW61+JKAzCpGsC9hE4wTVb6F1IO4ozWm7HTRUxU3umhr1M2LwWQyFHAj
8t2ZKDJ8Yjt/xuWpWRs85UXTlstutHmb/LXI+/ytighLvvOuxjXS+aPX6wqqdF3c
eJlIyeHuh3TgRu3FRu9HHts2yBfXQ1VZ1oNdC61FZkpOOHnhMygNwhO0aMFZK8VY
PPEPROIhUw/Elc1DYQR4lR451Fx8U8zPnyZQq67wXDqI2p/B6FZ9YH0//W1jPxUF
uL5FZALa38SgV0Ds8fy48ycaGuGM4B4gBgc5z6QvEmvbnQXM7FHDR8iQ71Pehiqk
HbMA4qTGEhjFBRmiFQPH4TD7DsCVpqbvpQkqVbXJUJ8xHR9SmwN7oOj86IUTueXM
YsMu5QhrN01Ska7v1KuDiQNdrs/r8kyX6/LcB8M+8dyqTQlZOTYwnWXDWktgtPHt
pRUJuuRQUbryj320FlbsCHNdqnZlsUBQOhPhXbA1ysghsMsbA2Ei9x8Pkd4nA6r0
5h8/dgFz0qD8xQw/ezbx2LYSw2489rkPygzdi/2u5dXUvM0gfe3wcwRppp66q585
kToOvK6QLSsSpzBCW3lbBQUny65OAlynUOGk0T21/FaNn4LLXF8frAQvjOekUVOW
bDEZb5Kl4a8AELPlzi+bLEkxozWpHiBnvw7h1YhfFQZpJe9yomPwLQwcNl4Y4kUZ
CDOcsfTTujWfpNefwP0ryZiRUOlViYd/OeyFT4yV4m7QD6kXcdzMj5bsBqGnbiya
JFtOCz9NOlj8HMDosXjZFx1hnnGJKZ5Eah5WY+27P0zW+vr8ltE88Et0MfCQdKSZ
P8qorDkM0Gnd+wGyYqOfC3CMsCnuDNZcbzKHkNQzAysdn2H52gbXMI9F0BJaohzZ
xHvvEnl7yxGV7FwWUvpVmn0ck+3orfKasF8n4jDCxfEWnnbaSOESDlZmCL5OVrfK
EKVS+uQ9LmBoXfpVkH4RTLMFlDzotQj1+Ajd+fk9LGjKjNWWVqcD35xuE7x3BlS3
eFcoEXWaQn0F+ox/PTMfmV8UxyqiQadENWVqePqKz2n4k5Sp69NWwWKVu/U9mMxk
CX135jYXhhAU92rEfic+uG6ufSoPZfRGehFDpwbkIDudnEQUgjxzIiRngwf+NprL
zcxGJT9xt/Idf5taZ2b+rsLFgrNF60wxtDCjncwYLkKFEJe1+Q+5YPIXiybavLy5
yax4ELCM/6zTJNmlyMoFRpZc0AL6RI0XpQMD8bgBnAhl1P0lJufhMy2IuM8J0+U9
V/sqKZA1uDRw7XZqkOVVOnBtlrvV5EVjFaIZrfwLlr8xo3sN3OMoB/OlS+mau71P
MIrQHLHgfJenXmrILKfFdnZRnZH2Odtrm5M8FYDdvCGF/agvEBi04MQ8nlID15W2
Ug9U1PoITwc5ql39VTHimiS77HM+fXBequGVJeMzlGKOyN52B9jQ7p4ht5f0s8bs
QOCDROo26Z8CzMNUJAhTqJqRlyyGbX+r152hy1dGrBN+8JC3TD5+JJZ2a96WeRWe
ohsIamVfoHkPM2aAvj141I97hMaqYqIZJg/g7tofELm4KoceJl9ZVu2Wc3vtS15e
MsxIewq/S+TqphU0+ECtgRwywYO00vCf23S21pIDsIIDlqoViCi87IVDamZl6JHr
QOcdo9i3enZgp+PnaaJUOF/lK4qcOSosbsrZ+NlMGtj0VBFP6umve//7zgX+3jSN
86FDaqLHjuJLuE7x97NCj+r57ObrwaMSJ3J6xmyRZEJ0Kmn50E9PDzPQ5Kig7AWI
trTRukO0X5UAf1X0yBejv2gGuit+5+Yt998Y3GwCtBjPNPx2lgm5gV+sEyc2IldA
ks/bSb3ep9IDNviqGku/77CK4TcmMtTYIe4lo1hxu2meIW2kkMA5ZxBMQc6KLAS1
H1oODLTomoFW5mZ0HV3UY6DAEWaWTMg1TnZXI934tva/WkVpyKbocGClNgCwAhJk
SejPdtpH9xOTM1dMnV0hvgAniGIeFhrGmVTxZzO+nue1d5IQbEhEpjUIAXx7c6h1
riMP5BZ9ACh6oeogJQ3wQ4rYda/T5wf4VEiNfKrpBFJKM4UIpbud1CxK9hyj1q3L
oan77oaQU9gtuBFWwfrsI9gaKHRH4nMagnQf+1nX3kOqqlgzf/F0Eafsx0L4zGLu
TzwNVsw+BiM2Kp3vsCtD6gOgvv6yUJleP3arsdg0NCYjvEO4MV2X3BZfQVUUsRTR
9wthZl0fJDTO/0GnlrX/BIpDfu6OKSL3SeUpeo2BEDwFanpiNo7bpXT4doCpqe1X
E5+liFiSr52zCLPt/e3uExvBBfWMCO5UwPN+Pz4nmmkq1NYJIKnyrtErKtg/depe
aa9aC6Oa1CbYAYDAlifsNVw3/85Kh+0bSJb+dsfdET8V1P6xO41JtLFLcaYlw2Ws
4DBtkwHoLvrhSwALmi+9UBOjIz8RR2yWeMrMIMQUfWzZy1WYMZFfFDf2pfZC8Y10
auxX4tLWG6S4mGJgBNyqf4jGh57uyaZlMVh3+8RylcNWfUVug9q7RwD7YCaV3dNo
1cL6DvkcT+hPgod35cxvaxG/EZZy/7rXJ6cKCCotk7M9N74tAZBNc/S2fk1SLu4u
tDZBAJY1p0nRRr5nkqK7DgofX5lKZvbq1E7QV+I+VLB4cW99tKxEmwQQBxcSv0jF
QETGIBuInInXzILeK/rJidBlaxZPLfysLlgWcCHbKU1aEvj9T0gWhm+0YIBAxGTb
uRQJfqIlNYGOvTeFQw/+XlGTEWQAi1DrPKGZrNL2x/ngAA6wTaHTP+nfEcUGJqUW
SSkbGTLnvDSh3XKmkXEnvoNSa3xlu/z5do+28y60K7PDnRi1j4MzRiWMfCpXmN1N
BY41PzkOjihylxt+1rkYzh/pNPNIlD1NPnNXHAgLsW56bZmLR0bJhsfJ6X2xMYlb
MQNUaKvoiGsT916UNasNLiue5NIAR5oGN5gbXlBR9t8tj58CXOiDQEymhOtznvrR
gO0Qr9eXSRqhKM/F4Iyiuc0zxs9YKUwQn/u66rd9bnjne8RC0TR5TEHopb2viZzF
stlBKk10Jnpf0B1g6Tm3+dvd2+RGFwPJBX0UOeJTbOKnts/KI8zj67cRTwScBZhP
Oc+8WYu1bX6+je2G9ULconH4YkwrBw6bVzbBNzNPeHKjbWEMguzr1DN3xvSIf5Ok
OYR4ROMp8/ajt+GBibdxuDMOy1oYsSud1TQ6BJKb4XjxbL7Hij9Wbsymdl64iXPJ
Qglh7mhd+k6sjcppMsuh5qlznA6v7YAi1DAWtiK7TAUYADisedlpGcktMSSC0vMN
mt/tNgTrnlbI4RIBb2ddl7ONwXDc9EBjjEWsvfd02Xfst9kqAR2UT7aKyExjSLCs
PE6aN8TA+6g0s64CWPmVTwp3cBjx6DHA8FiAdb84kJZJKzWc1/wP2B3jaNwZzlvE
/5REZRaSeQ4J7F2+Ot4BWVEb6qw8OOqF6w/cDSqpZRdkfsMJbcf/zZWJjKQ3tj+T
PtQdd3GIfNxqZu4X94ZOGoA1Q7Ev3bHQOExHhrVXPE5MD8O/FI4wDEjUGRCj8jLp
Z9FKoWzraoloRhSx9C/X+rSAjELJkdI0Iqr2X7sEgPmgDcV2xfEuNiTigZjmaPBe
7RcS+jYQxUzxX8szK9B/5NuEvHI1zf/lxIbPWmpth/UnbDFgH7auv9yG0B54Paw9
Yjv276QjL5Hh5rFKNLMFh+kpuMIFdEbtLrq/id7F6nG5L/yj6Dzw4LxUVet74aZT
2gCi9lHuqVotcaH6wH9jmYbKGUdju9JvRpqIkH5DlTvs2+G5V3i8POSmWKkFz3aq
+xiSqZ6OstzyHFTjrHL80/j3Mxqkp9+JxYTCnBZLlKYmV/yNqZCWapgE063jy3tB
zxOEkAgO6sO2LdPNLjMnC/h1j9B13iOjQDJYErKdcFiWGwcjE9vu/RgZXbU0opwp
zWbo05hb4WHg/0XinbFSUXgZm4tva8Oobh7L4Fn0Ct53gEq9G06UNd9FMZzTJqnR
/xj9YL5JjPCDkg+l+FPOIW+4RvH+7PkRKANXXDjM5gflww6NaxmPplSKHEZlNVJP
8BM1jKgI2fB4iUpLJIkML21bsvQRPjEugVrftSyapA9h5AmyVNwZlk/g/NsIuIYr
OjFTMsGYD2cn3PN9uLYMlhEHDUNhjkjs5SGgV4MPhB1zlUEPgWwiVk4tKxaKP4bt
0Xa5U8ul6itkwbFZjpUk9oTHfuBCv3Pm6RdLPES/2ySOdP1kkU6wy+JElC+nUOxC
CaAQ5l4bpPI/yToXMDpIEAdTcQao4Yc5EX3LFxyHmQ2pMmQE28SW5xu13euF2S55
UdZS8Yqk2tPtEi7+taAu4cj6H+juF/tjbFxUEd2BZLw5vFFPbcWobAoiRmwM8UL0
rAx2GDTRtaAyWmiY2xzt1kOuCRMw4l5mWfe7Q2A+cvK6hXB7C8Nae1763bCQDTJM
wVl8Dqc5hhEp0t8YH6G3xFwmNzPUHvFtpDTniiFQipeRpXfCkjqljUEYsvnuOt98
CdiK6mlJVDO2UwSmrFS/qs+mAsEMLVbeeyw8w27cQxgDwx9+NmoNNFwq4/q5Wn4i
AuvukigyHPYtSQd0Bgk6yQa9CaQKTlCUVbH1FeBDCb83P1gZ97w/nJv5RPjGcGk2
3yYBerqAJPyqtlmea552KwftXPnO7TKyqfMu8IT10L0ewsZV9OAggBu5244xJzMz
uqyCGJ+8aoCDgPFy35jVkyxXg2e2ZXqT/oWzs6Fy+7dQx66A1tB1nm1TnT4ZEs3Y
57+PcAH3O5kvNNq2NGR9PAbzHN346TLryAuo7vqevQvyj1aHTEE4Y/7vmA+DLauj
EmNPfb9J1Cc3+rFsiAjvqn6Y2NoJ2/EpSubC3Abyu2+PrMlVf1ZGkw31citYF3LS
/+pFQ48FDZQxiqDogPDJgo/uc8a8w8xgkDAdSZx9j+R1fuHsPdOgpJ6M9cSPZvOP
BHtbYEeiJVkTDoK2Z8hsZJAYOkQKJuyGGaH/v0IUUKeGJJGGNoz610KceSYofikv
4U5jgPVeVFvacNAcis9l/BQbGMP7ayLfV+bY4CQ0mENu0MGgvgQMsD6PWStMuv2V
VoDQBJd7ApbIUXRtU2EKVM2bGW/mc8OFj7Y/LCuOtYaTJl1jNsNJbx24m5bjee4n
Ey8RvU+9uNpYheNGxcqfGBp0DAv15pVlT1526sDZKTyVaUR3J6pcd5ml7LryWTCF
JxCLe/vlTeJFnoSBhdYuuY2U1R3iNklBxoh8IJkVsB+M1dMfjEJUdRDCp+BjIaSs
712f+/6ygXHjfecrsfr1S/vo1yKsStH5/dJot7x8u5foM5JSHDNeSO14jQzKLOf+
Id/UJVKkYRfbnzopTLIaE6+5FJxrmNlaoNMtVmvXUULcg2sLBhR6MoXBSajIjNUh
kOm4T6fGz8fkXtc2mRsJ9fIkSJjyV3coOIr6t5fw2iKE2PbfQ90vrRUjmVd1YgdH
jbfNpT9pxV6wm7dbB6yaNW4ydFQHychTUqQ7tWiQDhsBr5vImj3qQZPCfh2/Y1ad
4yT06q2TN66r0ObNwQCoJgTTLuj8qP/+hVC2JKE/hNRioDlJZMaP5SAHSUZrQUJ8
Zo1gbKYQbAJxhOa8cDf31khng9OdXwPQdPBG2jeAt/LYxMKfaaFJ2FGkzYQy8sCT
H3r5uwVGkODCtm0A9X46zNhl0mzwNc+YBkyBnR4DidbGqWxQvvXaRUzqoLdfmaOF
Rkyv6gXQ8T57nQ/kSu/s45oQ1r3uvZjImyWywr1GsKZ7i98PEJX4DywJAmtSGiax
BgdEwxEygD06c6xAZu2p75RTBwYupxgZEBkn4RK3lmjBNJjV1lXWYb7o1KhjxmPB
GRvGaLVusmEQFnSO8f6wQVVLCPkmaL4AH8SjBcMILxYgBX8F4UkQ3cIkdoPXX2Q8
Yaj0fPLG+CYjLRWQjsSuoU+E8Aufx86gCDl+LeivYf/OscwBPFRZUoW98ukHI6R2
Ho7P0ytyE/CHdSw2BdctLdDWKrC8kJSeqbDKtYcZSvcqRRJAjzP8Y/Kvs4sulgZj
0NeJo1Zp4Uyxb+Tcf1Rjq6xXlTgVicfg1sMxGfnbewbqq+fA3HDegNwheiKFNyGd
IPKd7uWcZJ8hGGLVZW50IKKvBkpFSkm1NNKufpVwaTsbgqBdYWznNLevlIwO3H1X
ZiZY6OaTN+tZ+SkD6YINioqShP2wUerIaJ3fLcNhSk7igEQhhJyaXToe+G8OKHR+
nYokplTxahUiJ+bDqn8J3p/XXFQrEse5k+Ddp0Qc/0pLL3RcLOgacq9lD9Cp3Q+0
uqWToeYAnGdU70k3sAtcwuHnXPEpRCBL4nhBJ49nk9k/HRbhvtzIEcGIEyC8EQuZ
SjrKXud3b35nwFg8/8infZVRn2W6/MFq0wkQA1nIZknGOvjSxCU4fZGSXDRy8nQc
bXK2tYYwh8DPKDl2ZOjfO3+hbWYKaW8SE06lHUhALv6ZlJJV9x2/xApPYPWAdZa9
v82k3WMciyzCQuAaixL71Nrnebpb3XwL5Gq+SLDoEJIs4iibw5kElPB33gpb1bUX
m+rOO9MvXzYSNZZfTQ++hHHVHF57HHYkvp/NPSGlEM8fFe9ipdNoQES+IX/FDLLI
sfGaaOYGyJT84qZPlmMUUSCB7ECF98VKkUvxAvQHmGF42ZM7z5Igz9Vb70WrHEO9
wFodeuSsBSvxShio0E2QtKDaIy0ulq86GbnSWwBbeTj7vIYH0pWQMWtsionq7BXY
OYGpA5isAQPUMW/WpEdgUrDUWk3coJ3n7R27xU0zfaSids64zL8rVpC4fknxdjut
FLfQP0wlZ9067GoIIxplKgPiTKsrXKN6q9w94nrgegXpgh/Tyu4OY+CyRfp2waG9
epPhJN+2U/C6w7bdESj1h9C4fUNLC14adq0mSDAbtyQFMKJisROdpzi58+z/tUMC
0rlUr5pbMLdlPTQXC8zEe73hU59Tal0oh68izdokFS0HBFZTudtZbhsdz8Lzl6Ac
5Ra/TTWTxuazKDcbBqN9qCv/6em6zDosyF17p3X1iFpY0+jrd5HIjrhplUvPLdkw
rEKJCBsZSuEuGLbjy5vYRvUatYXS7+TKCzOVBbZDMOdr6vm/Hk7pC5IEmG2JICn0
lrDHl3OrhOYJX+WKzyskxB1ijDco4+BrLwhtBORdORSL2Sjp6EZkJL9+/ylmomYE
JdCENjpcUDfnuxvkL0zEROWvmI/JAmLjS3puj+Zzb/R/HeXYOs/mZ1AI3A1FnuOb
xwaloQz6aixq/gP43Lepo5SiMYHKHOP0W42GF/F+T/iz1NNkh7ilpjy5gk+nfP1+
EbnUivuBtxClH+YEs+wZYNT99vAsnPsE9g47Ws+lxuD4hK6KFp9LzOLHevbVkOnc
DWoZepVMSIrqgfOUPBjpLQyU+6Gi/5gW8R7pqL+ia1zFcLXApnp6+1cRi9dgEkJr
hT6rusAQGWvfUgfq+HsBp8+gmOyFojJgkKZiHqukgWYk62aq1E2zz3p/UUBcvwie
LdVx8x/6vrx6hEpa+K6NRANNDwxJ9Qudyd6daCTC3upn8pJRkj5k3iS+HZEC3CpA
YtrKkra44iUucS/6w5OVPY+kyvRWVEnP2Kq+kIDAS8I38y7agDhvXaD/v3+9Soxw
5gOoAXQNAH7IJ4pLjy06yx2PQaDaeAksUzUN3M6IwwLr3zoYEV6kCUYt1xc5a0sa
i7W6l5yad1bLK8vm0+hzIn9kqa2H8UB4bH95cTwklycUrEphBRmvSKgsj8eJ00LI
Uhb+hJryQafNuSJcVoaHOaojl6Rt1olpgJOP1/bWItKVfxI/W+jlLUPqr0OD/sX/
Pr86PV5p2ZrZ+sUxMJ3g+qTX9EDh2YrPtqdYlnwqAWE3qdbdq7fm14tgZLPS09XH
jDIKVv0zwre3PYfqcVd59KHBHG0eVte7DAdCA5z4UcaVJmChfhYISIYDw2JKpjly
6sTZDMQEAJpmow8uH42oSeA7/TK6EiL8gOQPwxV2E1etKVP11HW0aoQXGx6XPvrR
6c1oAH4wkwdflMQLvliLzjmetZhRl+0m/zJV+560sn19M2ZyBSIa+ItNT4thd5B3
b4y0/t0zbEzuxtWLp9SOHw9iMs3KfBxY2wmDkfhCAUgLjQj4VUa4ujd3yH8hk/Q8
mIAgnoXI0d2pXPmpO9hLfPJWe5SYCLuuP+6wP8B/7QYjiQPhHHbL1tGEWvmScgMS
OgilHJotys2JHYlW+1iQwlFE289vQGYKg3a6mPSeivz9mOt5GzG8Jxj8A+SXdm4j
swT1c7uHlwxiEdISmzTK5GAFJ/LyNUYj9xP1CRnYzEJp+T90Ani5ZHMQrvE88Mtj
ivfbjwThoMCRfFOVzhgozq0ISRki1vCsLc+V+mviDuWrIfSFm5uLmH6lf+5ZmxXU
u4loS3EznoAyfWpMmwbqClBYBFmSJWpQZ3pC9zGn0tHqzFCpCEXfV+BwFeF0/iNb
72WxvUMeOpuZSr0df5ODqMMm3QCDf+zXN+YZ+19DChsEBGhfHToyX1LQtHWaIlRX
a7F2NPZtxo3MJAWF5OcWp7VA3Pob8a9gD+4PmJtX5GmcKJ1KtN32B4aMiDe/mxVA
+NHzLj++s4rMUYNT4koGMFW6276IS+7YvVgoEjQ7QfTgAs9qMEltOb3G/nLRNKpk
NjZdeWYUS+RbkrKT5OS3MQFX4OQxlVaCCBnlXdwXhn3I952x+iJD01aVl5otF7/B
CiT0kQAqgYiJaNfTh6XTWAxexijJNCNXc47QT2o0tyZfeafz3lH2CbFSMp4i4Uhf
+o2ci7atuM0/YGXTliJ/49SRmBGxkvJO3xxGcYwY4zuveH4gxjmMjnD0m35ryTa2
T2Q8NMQ+W/UsW2CxPbBdxeXHBKIvwNu+eVcfswcTingOwlZZMxUnBncuXAFQvd0o
wPnZ6VVqiECoQRWmayhy0kIWz0ZjePu63OTUj/wbPntR1Rjq5/u1xl0QiRuc7+Wx
sDxYzYwpFjMCGEKfa1R9bdQsNyjkeiNWXr/iJAtI4HG7ZRH8vAwtCMjZUgMhNJuy
8dbJbU4uNRuaCkgfO2ueccB70uuDpsAwUBu5LWR6GnX7NzNwkkbBbPMyZNFftLQA
dhFN+5d4KOQ7GPKEXkhcSpKaHA8GPRSN81xzsmBAnkgz+nZrb8NbbNjBxnJPYBoW
XxuU6ZFto0Q/AGak9HPoSgpG/on4NL1Y4Wkp5Tyz/gbwV/kUYH71Rc0DKBLrEQvd
LYK7rq1EzYtT7aaYVJjs6JmBQtm6kurix56gBjfc11an4DiX4brNmamYE9JERN21
4zGuL/+1RSrbzkgxxLbzACAWG1GKU11V5hV95hOSmTHdCsYkiFV09D/N+RM6u6Yd
EOpE2WQ8v8kMttBZifaG4ZDGsqy5IofYXeFtp6i3XusHlQq+rzkG+Eh8xYnp549B
baMQMhfh3zyP8G/50TToaqnVod5Dq8GSK1xTusVAHpsw1V3pX1udtw2tx6SQGPZ4
uSxDluijQqiPZM4gyhKQZ4pKMNTptKMzvY/zfPJDlMSZ1a9fhR1cqmSSthCZD9Oz
e2RrYny412ggX9c4thdRtlbCopeJRuVHsZegnMqsKPBBSjleL7gd+1JtcuMeFthU
uI7hPQtEV0+HHvFS1GieJevPJnU9sr8H6du07hagmKy8VKmk9bv2vpTOzw5g7+np
y85So4sXK7nUTIU1nG5pI5ZQrN1GW+yy7mUmD8EhQ7ekYmVfEJqifZSk6T7sM0K6
ejh1q3B04NEqf55VrtnFDS4LF/xZwseOU5hBg17XR4PQ/op1cdd78FUNb7DfrWBy
zxOURZ9N9Ym3dy4gtGw7/7GW8aUU2CTwh5Y66hcWHl7uQsQcOW8JdhRUae2Fymi5
8Dx9mtlGH/hRUG4A40cRFWH0YaxoWuOBm4CpaEK39AN7bdvEZwBzUi+Mz+Fv0Gh8
MIn/blek8B90uC1HsRWibs8/oxI1yEBUtg3/93uZdB0WpupeRz21gGx0ajNdTrCx
HYffDkjKajmJOsvyyo8Y44cxeXSnAIhweb956NEMA2BlDY0hvC43FOZyD2dZtohM
iAy7iMrSMSi26SKzxf8QVltfG7a4LjrFSW2HNA+edOM2jCP10uJtcnSHlpojd0ED
ZheqvWdY7ciehFIT37rZwT7cpmADCTL4JL0tlTOYtMgNeV5sMzklfPtcxYJOc0Cy
0D+lOSlv15BUq8NCbe0+iXUnoYD0EhYWe8cbreuPVXPP/Q2AsPbd3qxurhABPxJA
mInZuH2Nz3W19V6Kg6tJfiYWbAHudpgSp41nrD4zuArDmsuo1SBbQ02IrmqiKiiP
/1ZMPRspHI4jih1i+SCVwT+ryBNzl/C5ymtMT2pHaBGHvdaP35rhEbRshssKuprI
O+u8WS7Jvb/lNPLR2n40HHxGbv5NYsbdvXdaoLILZJTT2VRsSNh6w4j4JyKEEtTX
1WWyDkyi7jmBizzAIUF8jlwKr0qUfcZMmcTMzCBb5L/24Bs23bQy8xDU9WMFZiAA
UoSsyqU6BL0pMSQ5Fe/BwSU9+LV8ypHmBYN0ybfkSDNBf8m180fy/QuJJwCwVgPS
9lpEmqWI3RiyZqJJTOCfT33+4MzHGNhXDAu0Pum2jrzDIYCa+AVQfBegzhZZ1/NI
62oh3SxpLo0oYheSUe66OyrBPkV66DtOIn0yQ+5GeShK1CESgh5LE/334pEgllUi
drIeQ310Xpmo3eYaCtM+/zbtHAgCST9co8q8884h8LCcoebWw6LHeu/ASSDnk0DQ
1bRQ16oLslcMnE/MV50yXWOXAxldGU0/lZ58jsVfB2craa9q/XtOJ6KkHaL6/S2q
JHeWc0YOhxrG/LZ4ouc5eBeDUedQ8Z/emIL0g6/1eBNFfGzvXOb3WpbhwLJo1kk5
mVKLGenKnk/R9Vf8VT20CqMLSj/rB5dXMj996RR+B4To+up+VIYHHbtRM8//HpgJ
au0dK+Iw6riMp3CoME942yzfqYZTD5XiGeveNtytniOM0QZn68GW4EWvFZgpC1ED
hSt3/JiFGoeFyXi6SSxqutxQlBDpdY3F/lvfxmTk0UygyXnhrwNFdLSzg0rqZfzK
3mD44d7xLd6bOjX2E1JzXAMUqHqYqk3/5QXDyk5UgroGhKwLLLtp77Pe1XDfownh
RURoUPTuRlfdZpY2/CM+ae8Eh505QD3+afEhEooTwppVC73MZ9zrPi7sPF5xeaoA
SAuJC3G4RNE44GLAjGK1ssVNCOiy8HAOf6aJBdQPdPGcFueXQSV95yeDI+pXJhX1
T7wbsyZsGzxfPmbwksp3BTVunpw4ElMIZQWPy1y6DWMZJSuouarovEhHZ1MdQ0ct
uMc1wfavjju1qRWJqLj2g17ZF4fiRAPgC3jZmv9L+6/TqRxefFRq0r7VliSIjy5+
QsQGK8QWoz3X6jUQz5UrwSlVZjdGf1F20bU3zP8qUn9COikNwiscQeKlg+yeBlCi
jW3j3EF1Z68rI7Jc80NzIasezVrstcZF/UsEidnUMtxT9/+As2Y8UGv5zykwjszo
vv7cn2V5p39tFFnCfb099JFDmDqnu/6JRHuPJn3E00Rh7uwzhH2ol0n1CciNsQRH
U501BzKxjGLHk6aZ8Lb3Rknd6nWMtjUT50ZAzfqbAJ87ns6ibzD23BPu4Cy76pkP
t8avjqkbkLq3iBewSJh+hxJkMDPEs6ytPlNZPgowzQ4LxBz3zNB3tGIiaWUdfSjg
OpZP3PvzAjANDiLgv0sD6Os1kOeje8u0aLB9YwW0eH/+3ow3kdQ1RiowvlPrAQSW
yEASER0F6cAhDJzlswrlVBFmlNki4dtAl5egll4vMhpNmxjyvTQlU3vccoyVLWtU
5tQlRhXkonBo7GuJrYH5xLv/g/VD1x87GqcWu5YsvCJLg4oTQH4CzhSp6h11TAEK
zhly4bQNZguv0Xrv8l4WfsZJN/hpFJ4vK0DHVaseyKvjSCibOm3EcO/vlXTPRyjK
iXPKqAFjErttaAAqiMnENvw4yBrJazLwhKMCZZCniEOf/mt5YqmP55RrCBmLuDPP
mUtiAD40lfKiNRz8npGDX39qVTsERUIDhrMz5j+xiFmwEHz8Uz67delQAvKFoUnr
lbOP57QMAE3pBOId8LHb51tO8W6b7uUPuQPlUjcVvbR5AqeUcDHVSu4fHtv19tzQ
8jq/bP96DpPSzBhDcf6aUJ5BzuKFP1j2kmDSx4E892ZDT9ueae1C98ythTFGbhXS
6czVxnIQCw+gVHFaBAloTOV6cpQIdSmW4ddAgX89RlfZd5XuiQAaZPAbswk2k0VB
ruEB5edf7R/9JXNXpkzGkit6JdgjKLbu+/2j5N72fh+kj0CUs+gs0RYcoOAf0une
mLVnysICcPliBWdeF0tG8S1Sv7e22eFhipdJYdexI41Wtj6elVSBEnWmkfWHVHt1
JiNS0izA9wrd1bi91kh2DeBtAKjdgDcZkroRRjmMRx0uND+VMWGYeI7onyyYXWim
dnEEtjoUcqnaJJTBJ8Rmv13b0zy3Mv8PXQqTo2gWxtDIXKhghwr01jttY5V10zQG
mEWiS/hSdaCzylvV/nTKpnUZ3CE7ZahWo159k2mWZaIPJM1ECroo2fEYPYUd6ASI
pD1Ra+y/W7TC4lrslFOvnqAwAEUzIgU36XWAPdZwXlbTUvN+MnLUMk1FcTaV2v2q
9pFq1X5KedT2XNXL/RRfCLpaiHxIcWdI3XmpRmBKgOIQ9+OkJl2w53DI/gsF5oed
lVskcXt9tZ9cNtRUc/Q4NbgZbMYL2wKZWXwD2vQhe/wt/g9HgTt4+v8IZOqzPROw
327yimf1ViG3sJH3X9kff1WyOkdYB+Us48MCY+fTmjsRDQQyJ9gBWkfc7nbgiUi0
RFGA25ZI6v1sqccLec3am6adL9SvmF+kamkvk2kGKgPIX7x4WoehteaOnUNTxPg0
RCiVPVwxfn6ljtETH5wJurSj2lWexGlJmB+o0Q8LFdqjdtBZtRycBfiA+2gkniFU
3R993Y2uO6hSQ72QUwN5HfNYRcJ3+d0EBmrrRc0uIyO5DFwVeo0v9eR/AMJunnpS
Fmt3XHpWIeTqUaiff2Kp1JFO0eYdN8E/ju035ZZA+Qnx2TdEqes8zmH5WFO2KDPd
IG5JRUO7gE+wfZVfW+jXE2P1ZVcFE0BDK7XBau6iMF/6Q/86Odem0zWet5HquUEh
9cngGuXpssTctcqT1knCFP1JeaPNkYOg7VBRIu3R7/nsIwPPmIbIKWAF25R6dYW/
UB4NvRw7fyw7r57vpPgpIPSSE2B7Zg37I1CCvpyrI3hgnNiUSryzQje+KhKU24GG
+KRRGDpYGPfm6vMAVElhMBkb2NSWeA7+Wk4EWcuGiw5fdyzznkJooarBuU9LPCWd
9/5ucsPAGW6Q2Oeg0ZYexOoLfq2CgRm+PBdkvDqyifZbICLkc1uBYbpqooKAWq3j
65FrjO+5f3GlTEiO5T/S0aepxB4WfMu7RK8lMS2aOblvf75Sf7wHX3MfZrDN/c0C
vJRWKy0CBj1GXGOHNEUIkKX4gxjvmk24zJSqUFibP8NjQQBHBcF6CWk+o2Q9D9D2
gvF5SM893vbzOixIm8zJMojjBdXfyBRXBBkTpU6TI+BiW2zSlTTAw2Gm1KUTgCXf
loEuMdiqy9NgXQQEgiNkyCdJLTXbbH1MZeFQ3kX7/abJJh3L3TFUTLK+mgF3b8OS
qjDtHBvlvpanf5A6HYOLgMF2+yEDQpWAHHS4QJvynJbSa/BgVuxdybkyLM0Xg8es
Gw8N0t7zHI006CoGpnLs1qnaDSwjBCI+rRc6TknqiDD9XyTy5NyR1Bk72dJWNrCA
eqzsp9AeYwiH0m/dIXReEg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cDLkA+axxSt4s14KEA3wYgw4F6cTEAL1YfUlWGNbRnH0fRE3O8f0mMMuZ64h22h2
zxJcxm5zV9ltTbodjnGFXXTPxbHE2R78/gF7UPW1cSXO551XYSOEGrRtQmvNOUOk
ENLpneK+lTFbMfjaWq8IlCwbRUNdrTPkTV6MRBCMPwt1n4MHeWaIjz2W130zEfOQ
0OANXlwvz646MHdjVlqWhAojXMEr8vtQpcUzaXIrIE1mpIklKa1+COunL3l6q6Yc
QDWAMgBV7h5QJaHiTL10EeJKpdjIdVTTris33wdGzRIpwi0VaZD5Z+IuY+Ekyg2s
njmeoIN5rBHoRd5caCuPtg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10416 )
`pragma protect data_block
sogY41UwAxM8wWM71KPYgdGGmBsRrjHAoU/rnhCWJo3bxuuC4rf521xwelmodpMs
YMzZnbixHcuyjpvDm1DEYNSPJ/JoNTXf7HxvX/k5hkPQJIiJWy3KTwrMRe9Zf5ZE
bjEZZVEIC46MAJ2JkZa40KlE1jQDLWnCCk0+bAify5NQubaUlBuOPdjKdkMOcgWk
iHTWcxi4NDlH1UhgGzAYv7W0uuC5DrXusGRk3LqdNGyxnSNU5KBtm8bXXavT/sCm
Okx/8Y8OHF20cWeOXdAVEPlkdZEYv/+hEc8Z83p8D/0eM/W/346P5HS5o+X3aY97
Menn8Xc9xVjNjWrdfZ5C3WVuQqPkcDaeLdDARS5JcaZCINjftPYQljNWA7HqwHlj
l1giuDlqKHCj+lcV2bchBRyOFXvlsaIRJVv0dpzyI6c4xiDK8X1ArK2T0LrAl8JP
5yLHIa6oGrcnL2lwaKRfVkYVf5WdArhOtCgoF4eoOT21e/gXvFrlciF57Yy+JTrg
XWKyxs6DWasD4usX2Vn4kaVCaQN98QDUV95zPfn/BN0nzgcynLzHTCil9F5lEnGP
OZNICE3CHrHbKac0WNooMHfkLPsHwyHGzf1kEa7NxBiOjCocPf+725BR7WgUSfLj
jLGnJ9yErXSoL6Lea1RiSBFYNWtQSRoE3K9Xm1Ls+gT+Vxbz/H+ENxyV4acWVLgl
kQ6aJXVzMZvKDGdpArhXJlTy47yNcEeMiTrpUlomH/rlVkSpv+3/oHpP8DdyVDL1
FaIJERoErglFvOH75th4ULD0nUc+Dh76Kyldzdp0NXvhzqmATYqqlM7EfM99joHl
dx0MoX7eGemomLcF/BDyXwRqH/RG3+zT2uMN2pg/bMGJL50wXL+PdpRa9oUadx55
0IvTJKo4c+JvTxqS4Mxgi5WzbLi6ZP9Rkl8RkNUa2AKtSDs0ztQZrGgBffTQkLRD
AOBFO3ZulwgnldKlyWd1dST7+L+l5W0t8TPaC+vr9SYRSfaZ4oAzLBawHzO0B+Yw
GlAip4cR6lTRsD877XYP+MsrBc4nQhaJrNzP1tzhcPkYk8+QFGDMRqFgnmWNOeUm
69WJMITi9IxA3mJ6YLwqCl9gzfTs3+WRzYl0USqVcxoHZ4lNrXxO0prT4+EEvhR6
DY5hKYfyf/W7Hrz9R9mdBTx4yjlNPEoxvh5KhAgwx3g7SS7NINa9NRd2V1m/gIdc
MfzVH+AYBvw9GoZhLUG36hY6GdtJG1dTtF+575GHIC3HXTzyub5OfTK34N25BQCI
1x0dF0EAT+/dZjN3O0Abfzj1CKNh0qSvCy+hEboNn6lnEek7YriaqKoRKcExdqnQ
Mhg4ZYcROYgnMuW+tQuiVUx7Cue7dBAW2FCFes/Ob3tV4xaYXAYw15qGzkmZ2rGP
gPq17PyZ3MCfpU012VerD1L/ZSKwTaHpQ5KOtYZOW/9eM9PyZBIukfO33vCJpHYG
m6WUabah9tX3K9p08mSHkQW1OVufKQtwJVR+XMQRgcmT/lHlLNGEZogwqZ3hfNGS
UwXtoLnFZ4hVzDOEYz5UAf0s4liajKk58m/sodPXT04SSaOVIh9YKOm6vZZgPbWE
f546J3w6xc9whTmylYWhaiyBkyUdfanfdQBMuSYyC2yCpOZ1NLoAT4/IicGhZgGg
1rBfz/7Fmrtkr7YVc2q8tjAIx7uCecZ6e01VRq37WFb1XxZ9cguTP13IU+7oO/XU
BkWff1y2DExHWk0yMeoVx8INsACflPIRggEpGHdmiCwPNN0U+azw50ntx8rXDm1O
6of8Se49rpO8nes9EFVyr7tdBFi0Dmv/xAtzOXBhZJfQbBKPRgOosSlV67ziEIbO
pvJ5d6dgn+qHxsuFkSGvSvpN/Ek/tul34bvxPeq0+gVoY7avyAovkAANih3WHW0K
YUCPhVm7GHBqWIdI1eod7+CBLXoYnHUOLg5el/yX3q4mvx8IeUr9Sw5xNXOeSg18
G0ZlUuzUGLiQznX+JUHu85DiepgU1X2lOR2Ckvp7mDI1ZjiFuLMrZgAAcnkKrTdP
TrPb85Su/9rvgmSixInbjz/rtJISqj/cocNAT887szbaC3xWtqzS6ssn+QBLvM9w
3iF9ggJQmrnfgk8CeHZUlNRHY5c9OnULwtxxeMY3aq6UvgEdAHYOJ095GTfyLCUc
N2Ll9t2C+OuHnHDuZ4ngeWHAqWpUBhqOHt4Pg0vvSyIssjQQjktPeAVE32gvl8jl
8j8IcXqrsfc7VHAT6CLjkpWgsUWRoieGpeE/oJd4V2zZCyDLIJJf73HsfNSb8mN+
ZuettfuT/fhqUZlJdesuL3i2gEWcb2MUkNIOS7uCRhdxJ8iUPo3MVKDiImxd9nzh
8myk0wXarwP6hZbYbb1grPu3n2FpAU/IJN9cS6rVGfhkZ9LI2ZKAlz8w3PUeBdR+
W8fxGXAIk8YkJGpCM7ogQ00eYC+g/ya3RFcqA8hD3nfrcOyWasbqjFIJBSL7roav
mPCFLRwuEJ8iNjDKGgRqsXSC94Cl7gAk6lF6vFXF+UAK9cWhWw5jKbVYTY9TRzge
lPxpa2IB8AAcCxP1gPOo1WSh0E3QSW6ETYC6J7R0dI6Hl97i4x4r5DjqZurt39xv
54J5DFpy1Q1jumXpTIWtZxsKUN+SI6uspC3MhSpW+P40zpjh4324AIyL2TO6lYMt
TmjrXU0BgMoeSy+d5MLalxeVWQDU2lvsnt1EcDsMKLiRO04hKv5DnDRxndyqtrW6
8A5tlzAQwPApvtpapWAy7205vn8S/Xi5PN9TMPrzHfnvmkuhEioi7QM61sRSb/Kf
DoHzNTtS1Q9tNOBDN0O7QpWV0xgV86FMsdja/0pCmZHOeKeJqpk/+5AR9XGcth1T
qCRs6IRij4UOG0fZvqHfKdGyvHsrd5gn5+ObVDqMbspN/vN/FuWasa/VkYyOA2xT
9pqQoqSv/Y0iK5CnBis+iZJKDseiNvT7eX2WoT4xHLwg+DMs4BZICxcTKQMPmBCr
/Wiv/BlHpcoxOd2UU2hJiPwKQP8Hr3EuvecG+poMpesUnhI2BtewfYc/KhOgzrg9
9XeM6r4BDIbLjTxX5S8b/E5M16RxV02O3jOKuv3SGc8AyrCVPaN6K4r9/or16h+q
7z38WgcKi4b4ID1EMjUHGFABjGNceJmYX+gWvornGKiQ+qIt3wTuftE04gBOAQCv
SW8yBWyF9deztVAlUH81Cv/5L/lb8nv1V4USkOPdSRUj3H8hGhrDySXMPvPEY1tE
mAtiMmQfeaVIb7IUhH+MYR/8dvF3sCf03FTxmlEDSxxW2s0YFwXvUtvBu6SxVKIT
M69gyZg96HeqmqcDMlx9KcqDz2S9aeGi7aF+XIQAoqageqA3IxbD6BdLk9umClGp
shJOxjpBuGDleo9G6eX2RBY0z5lB8L+0AaUwu6mFE7X46eQTmPtvV7T40+IYRivv
1Z2xKiz0O1Rrfi7zF/mjULiulJ7vPEVLRHRzMe4UEn6nTvTWq0budoAFx1K9riAy
5n57NUtOgdfwSQ+dAbrDiYsnsLCcrzcA8suRkw2SMEsD5j0Ws6t2yv2xX28rhjC+
PSBiqPsU6X89mwbeqI4iRnMFDw3s5pbxLp53OZsrWRs6JnKLC0c8VvO8mTxtWPAn
zZPmQRsiI02e2geR75NEfZFU+nfWbUD1Sk3GtFLl3pbDKrGOVXtT7i/PoPTgoBa6
g/3uT4/BRyyIiKHdOhDHb0b6TvD6kvDspHXRSrbumHUxBtM7rjjTrspviAmzPrR9
KOcTp1WXgLmiRY9p8GbSHC+2cyMZRCD9Sd06Fv4TSQMbG0lBTjpMfeSqPXcRKTi9
BEKphGsKIFBk0UlEV8icUCktCl4OSu/rlhuw7wiuOwclKnHJ50Qy7q1ZgPo1/c22
PZK0Z4QOSDbni3h/7ly21XfE4969d9KNYX+ZpfjaxQdV6jBoSD8qd7ImX8RdBKPS
U0UiLP6Wg75py0eOC2a+N20ZwjU6mvGlNGVKGR6NPYbYvo64ETtiu3+qvP9ViOoj
0fFvF8ydoH615GZSAmblhzEcbd0IBYpZGqdBTDYTVlkdjkXLdBMid4OyovEbfv5R
6hFLyAbpee8Xd59VBx7OxDx5aDiPY9YbJreD2vH4pcPLzZi+X19uGPtwOEZ7OewU
sSvu3o9HZj5k6wrbPrgzaRmWrnbSKiwx8ZGmB8oiuNhL0OtlkPlFBxCNiyUrlwpr
tsESF8l0I5T+mkH63aMyw4sOqF4oMivzRnUkzdBlPI1v6DQrUK9KpZI3F4NpGPD9
9DtJ5sGP09IwCjq+47sesHQ1JqAWN8UpBtDraeBxIFy34D70wY/bBR/Z+vFnF0hY
mjksZzapC5lOXmaJ3O3Aeb4AZFZwKdSdMi1z2W87Be3Br4uYmJ7eA/8k5byuJumi
3I/Yj4FWu0b/51qqrjIskWAaA7OYrtt3Y9aKxdjVgBbxEg/lLcW0NhSETlGRuFR9
60CCVI/bVWon8Vo+AW80Vh/QiPOZReJ1Dd/R7tFKoUuJdiPmhhZl+IC7nSQgHyfw
hcSbrStUuZ1INmh4Es6/9xEeHvpV/ebfiOYX+sTFPaESKXe5nBnkr2QdqfM12OVv
gYwjwDScROv/8oXbCQI9dmTdXjcxkt3hAE/4gHhsKEuh6tTXB0WTyJzKbPRKFoww
nrLtg9wN/S37INmUvBDL99t7xIhW7tw4hUWU2MP4uBTmd2csAiHx82P+THIB9jnh
nzI8M0NGkoqw9Igu2Tl2g7Ll307gUcccOynXCHd5BraXBWKxoS2nlzfoOja8OmP4
VjGy21ilrvOtCRWQVOpWsVkAqiLoqR51UOwjdl8Navk8PyJqI8xflBOl2iPaVFBh
4bCx6Xmact7S4g4fM9ngBVAxgjV2ktD9QoTL7zUJjM7CUzzNj+LZtgIE2A/os1F7
Z+Ct74lhOLhZifJHYs8/unO+QatxqA26RELvVTR9cV45TyGrO44I02K2yN87MLrD
1OwpN9iswDQICYplpTtNI3IoRUH+iNZMrNd7wyN9YPEBwdU5timNvHcB48h9KQt1
g6qz+0bnh2LJn9PUskHuZhDH90wzaKHPYoYp3qiZ6lAg14rnRpbvvYU/Iq+JeUlG
TVosBi/IT1nJw33Oe6gXXfmg1TQV9EBCZgnlQ+1BQvL/Qy9D1Tw+dkYkOkJUGW3T
tI2F53GpwI8vkDzjAJzbyChZQj+yJmZ2uYfxjTeGivb//NziRMngZzRM+WSnN0xE
saHSia8Jz2nvJiSdxlL+SxgNo1vkKiWI4vEAR3G18tVM6v4LA+dyx0KJZ6NtPZ4a
m1gTOvFESpX0lVzwfnW8OjT9x3gVLaZlj4mxLZvCtWekVHz406F95XMTdsRT74W2
ZpYF2K4rhifKwh4voO4ujUs5SsLC513+++kKMQLrMWOhy9AFdS05Isa0Okjg2rRF
rav8o0U/3n0aDTpx9h2X65cqmenATeiqc1JUlgI3gSvnSxiaMCvVoiyfILaXVa5f
4e2RGjZK449um00zYnrQbfxMD2Gp5S0yX8Y1v7AgAnTz+09oC1SCOc7WPkml2GSc
/M1ufP0CWuwWqDcLHwwdSm/KDarrPQ4oVbpGLiHqN6z66wcGOXzMsFLqjOkAH/y9
UINvQ/b+XCalBfx5uOqO/IjJBRo5X65Ph+hlABumxR7yFW5kNRprYVzMq1xJHRT2
H39EvVbiBrnQhYDbGFVcyVAhcA/5FRaK3RRO3VR0VH+a3szlQTX/+tgT/RoBfG1D
F/sHnJwnhDfk2K+WYFhRZjotT6/2MkJtzPcPCIDAf8misV7LJevuiuOUhaYPPnyl
b+uYUAhYRMSHGHjp8rbzzBJZ1ASor7cxY/OlP/1t/4gQBUDpSBEsjidMT+Pb/D9y
99DuwtvSaFuqD1hcIpUkINfIITT0V8Xc/+srYCQ8TbfFFWHgjkYkkWXUF98PuJd4
QqwUxL8VeVgT10J0baajF8EiO5QweOt/ft3tjF/1XL5T3ahLs//bqzqh0VjCbgQ4
2yIUJZtlky3ZerRZI2mGQq9dODATJrntShWMHYbPCwJ7zonKdtzvhVABqFIZGnYj
0IKLzGFwxPiZOgu9RxvMJC75nB0f4yk5dl324vdrBTn/DuI8tIVNb8aGryWyPRah
wJ9Q1km+HCUPc0H1pAiRd309AadADuLilYLtrpgVxxssh1dmn7BblEFVz1y7t2LC
vh88OXSANJzMefY8TSWI6/6jMla/Q/5VqyyEC9dxt22kacsivNpfN5Z0E03XDqFu
ItVGGBOaUTFx4TtVKBRCb5o2atQWtw72pGcyUI6+OKV+m+ebgXSyLIa+fn4fXs7t
Q+dmXzsdQN0B7lrcee07qqWe4R3Olf5EMqR52A1HDkRk//z/d5LN6qDaA3dkee4D
eoZ4Uc0FEhY8opH46nLr3EwG5oLC4BSgpn/R4i5y9fkWfjH9yJ/Ae3FTVqyGcjlM
ZsbVXLEwwmmKCNArn1eTWlpZZsY67IhIrTnVXe/Ks/OzSrX3WhEBwvjfVImEMGvY
3bE4EbF0Tq47rQNUv8gWkb7bEnlOLslMQzuVOhDRLktDk5hRS2MU4OaPi4TQYXfz
90hKXLbuoZLfTscIlEl+f05TNOVxTas15bVJqJLp5dpC6YeLrFfA4m29jM27WSRo
VWRQ7FxWa83piDxkKUagwZHNiKMEUYdPIC5O/D+hph52bXY65rUAGS6yLUXnzInP
eTssGttKGmdajsUUfsyO1fct90NHvCgq5WEowShOK07/MUZfSyVpro4itISu+rgD
4UVgnN3gsdf/17ApP05Pd7lPlF2XeNi2NMPfLNbEjNv+m/xERF0Zw0LP3y/nd1Ty
w9I0THfxh+HT5hNn9+qyxxJ1+1Gb2EmIZimuroczSAmkhRGxIFgay2wjVDAHUXEJ
CJhOJc5ZE19J1X5eu1nmba/z8OuOUWDMLvnIkv0wqQZrDTplD9PLcOMo8H6uE+E8
dWr4shVRLkJVnfUwHIWw38kdaEwOC2Raq3PjgNcQJ/Mox2u0vbryUEyWclCKROv5
VqjdJYfUGrlhCpNeUF3soH4wGrk122gTsPvRbnY+oL77E33xh6RtndhPRVLB8Apr
UNvwdFQFQwADuj/+u1ff1XiINrCW48WkGHy2N5kAGf5S3200uPvXVdnHst5Rb7W7
Aj9B+kXONJPL7OBsaGOcy19cEoCu5D0gtte5knJYgdgz3hQYsRmTQ5rETKfKRQbw
JhW8Jhvy2aHFFKF+1HNnkyVbE2t4Sbmhxh90smBzpP3fuO3UOg8w4GoR2QZElLl/
f1EUHbUu2pcSPNzu3KTsUfw9X2xx39kvz+a72Hcg8UGcVRPttQWcvjH1AU6ZkoXh
3LYOg5webGRWvCpS+tOvGdN1zQ33obNKeYiuEl2Uf41yyhyJHh4uCrZAUUZdkVxi
NbAbpUsHFxcRixuhUzDv9lv8PAOUytM9mHYFfp5JuvHUasR7o4LGz8cIXTvyjbzu
UZlpy5cO9qnzjaAeo9p5gqyablSnvMDQLiei6upcoDfdwVQ9FdpKmt85M6afSm5Y
491yt/hX/I4zy7rOI13oFcJA/+LIQQDDR58bMD1pgkJeA/Uzjz2YUhNG4RfuFxH3
xb3q2L4zeeAXUUMV885gBz+syqSMzqEkSnfvNlDcmNRkKS9BxRZoXl+UuBidNQlu
d4j4Vi6pkcA1mSVIIe1GUPjW0TNX1ZsyvDvKsXebnOjAPPjL3gg01Y2ECOz+MLUb
fpH7s6zhiNb1N7s9VtP1LBPWkG/W5NcR/RCwcA3o7Ca55m4APB8R8DsjaYOFK5qO
K0c6k8XSVAc9NTLcIj7nvu3Ja3F9rjFwoWOai8LOA1bQKySUWm3foDmXCQsXBk3L
L5R15nux6R69tg6FC/joh+0QYAFdW5AHrOM9EaFSSt0CAYmJJR9X5jwZs4IcDEBu
anYK9zntKoU8dw/4y9I3GDAS0UR4aoGZ1VLB2oF2rXq+LqV/Flq10qqp5K/Z2TkJ
D58a6ru+Ty5QBmBZo6C2cvmh1FzHaCnZOV1uSBFXZW1QCODB+uVHc8g4J2GS7xtf
oNMPxuj0bsBEeiajORpCEFkd6yOdQ3lpccjh78MWsS+voN76C472TOaQvVWtDbr1
e1l2RJEjc8Ebsl/4OA3o3TIAyUdCN+GjXb6cUKIHVtdXHVTqOK7DBR1sxQRTVeaG
W+2ZdYymCVkKFNP7cWOalTIwNJtvI3yCuwTjbJFbKKnfl1i3o7TpfgTsmiTrwfDQ
QQNke+sZ6sA6pwLHzzd42hLgYrl21OjlVSHigFIOMZ95bb2V6/dgONap+NyFsEcv
EoeynubX8YziDBZ0T9+9kT8Ny/8tUvx3415K+lULNgBkitzvd29wfGI1TxD49LxF
kgvtmHhlsptZ/KhIg8uSZptcwoymGdjz3U4mj7mlihomB3wFw7QtsA6Vr2Ld4Ige
uwuMb/j/Z8WspiAQ9h9D3Vuff8e9cr5FM1DrTFuVkjzZupqdGug9gYkBBCLf/f+v
jroWPa98XXX28leEr2AjEVd+Dhk5TijDF1V69vMFDsg5hwZHSxg1RQGS0UzWCh43
IBSnEBv0b8j2HeUU7AvJb19dTo9Y7hPRDRwRgoo4NOHphDwhnIQk9ABDuRih7+Yu
5M0qu//ZbcVdbtQDsreSas0bXRuYGCUe+CMQw+AhRMZQkaV2IK7zpp4arCZaGBs4
no/HC/4y6/XYipvSxp10oW7Q+FlM+UYpORL5sbfWhe917tZ1COzmo/MnKMokYWLd
lU9M4MEduqQYgZnZI6ogXirfD0NFAUu45reZhbqCNhIk8UwUmg7ZXzW1j3Oxta2G
Ub+voysm3L84faBq5zoKLzmwCKvC/0vcMf5rQ1pMfz11Eym60nEdc9EawxBi3nVP
bNvftvFvcBj/u4kK9PZUqzhcE0EaTKLabJkL4jkaJei+1RHFcOJMe09BQmoBs+ly
B+BDWpR6vJegWYtLicgjQ64cj0C2M8RGaN1kTd735g85OS9k7vpJBg8Glg30GM5z
rFMIWF8tfHGf5mKt/Szufn8Q52nQmhlds4LkDrg4XwHgeIckfwb9JGzVIlQ63YUE
zZghe2sRPbm4Y7mNgS/ST0FRjKL0KNRLrbwu4DbDXAa4akowzcEJVyvPJiSsnjQP
Pnt5qvRsj8NIiI++a5C/XA3RMwYkeV1iE3duZ2RLPSg4o2d4KY3C5IgsQOVL3xe8
h+PDBu1BdIWbnCHCKD6gKH7zs2VDcXcVuPuItq7xmY1NLbLlysYDr/44GxD2yWyt
iZu5mQBVIyx8B9HALWvQf8ZTGCZa16GOeseAk20MTh7ctjKRqCYRdXlXXaOebZtN
81J+YwcrNw6hwzV6o89cocNrSDiQLGCDmlEXAA1TMYuMMy/zaUpaTKdc0OhAg+0t
srN8BZUV+sdukyIZZQq6z4WGUqwXxBAHEGGi4/E67IYd2yBiO2AUXPCH/+jXEPAD
AX/WGksNhzZoDd1n6drgayQvjhgbhWg43SPmcsZSmvo67rU3nL7058oNWcaMhBMK
wgpM505+2m42L8wewyeAXbXSfWdPTJx1sxWIeUAd2N/8caMY6omBNMk8hZ5V07yw
cN9Yvv67mSFTdyrkKmp3ekexxXbmLO9wiJ/P/lb7q/Bihzp6+zVMzDfUHq+Qq6P6
DIMUYlhQyM5PigDkiMbqjM41enbPhYU2leqGg8XPahF9YC460eCoGRuACkmlQcMf
57rYmJ4Ey/h+4RXWjolIb7ueqfn4V1Sdt8aCQpmhEAfCRSWYa4OpX1qnNzD1PkPI
CsJBKoqpQInoP3MkJZT1ubRRipoYB3BirqqUi+ILJnLhV4EH9EWrPRgmOQaP4lM1
QIZe2z7yH3BXavL2g6xWTb42o8KMeffyVdiUbUOnIvmSTGAecrlERiNVGTJ1yWlC
ONMs18MstZdrYmZQOKeVmIJMEhb/tcuJ4lGkUYFMNFByqbWxIq2n+H1oimiFCNev
wRQMv761OxwP90dCuuzG+gaKwzZyD1wUQjkTVvrnjJzf6xQOpkPvUSWVmdG2EJnf
HVoVpDObNkQN2QH/I+wApZH7LFIllUu4+/cbT4u9t8Ye2V059szTKPVfwoHXdriV
BPZDmng3mP9jTJU10hKxTlBvhdp+KeyB0MpQZpLmyGeb5LHKpWOzeRt4Qthjk//7
KMQrPKGioCTqtzFADF7qWEsyi3hbS2GBmHTnTtODh3Upv1oCagSdvXRqwfjHgLP4
kKZxH8NmGhUJJlcH+Zu+etIy6sBr7uKH9NxM1Tpo+13ZZyhh1hUv133O02DDCd7n
DAzpGEYKPduUReMXfdgZUv2OofQYGYSQ7cTFbangBLrN9FniYKkLGNOQmGIQQ4bD
O7WA41W43ZgtNkS1C0WhM9ROHJzmSgmWY38EHuoO4VFt1fQK9knYsqJkPpoNhrD4
+9vyxXfqI6QgB5KLPGcVUnTLHxgw+BAsq0pdUcpxtryUxrszTlTGRWA4dQyXqj+M
hF9Cz56wG4trpSF1Hc4nThcl8rSHvfb2GCSrTf6U/JEqZi2xbRYGug5YXbE4rXiO
XE0cyh7QXLF3sBnbj1j5wnxFxMn303LEfXHLnk2pMmNo7arGhBNh8j9beTT/oGaU
Ccv5DfDmNFG46CTT8eC4MkcJv5sLvQy5LRRkmEA0fBkbh/CZKaVIQZV0E/3pc1DI
s0w1uwSP9GxnbzPW4oj0afNxuxljY5OO7uqADm6qkHnAM5EJHjhpcgt/i/8X60Ch
PRXO+YKxACP8Qfcig0gxyXl3AOF6zfjFC4s43uWO21gzhOg1HO2Zolj1IJrGIfix
hmfUnkcRA1XkHbnX67Oe+/7aoSzThxq97DVeU+XQFDn4mmsaiQt1uWIOzS0gkzCd
hcFpLXgZSAnPBWmkkycs0Xxr7Q4pZvw7U2d55AjUin9BdNWPf3T9WkC19x9bCPrj
bnLGcW6Vhiq6xccTfm5DN+vCIlVEJXeMSUEvUuHnns1JjSc26eUKIBw79MVjm5oW
ETHHm9ScdpkuUhOJqJo2znQpRa/qXyH0R9EpQhNokmTVwVo6dZQwiJGDlZ3jC5hG
JKs6E1waAXIlbawAQZiu9UPaf8jQrMbwj6br999GdF1FzgWP9QNs5y9UcR+8Ghqf
whWa4PemkNkUYaWbH2TsXAB2Qg4Wmp3Idi1fb/Tt0kewpyBTjl/bqt2iap5A8q9N
Kq4n0zVtaf6lUyTAYuTP+hyQ/xpwSHsLWeA4AqfLXq1UkTgQpyv7356v81a0QMtm
cjcMuN2cQt+8sqxDT7vKiPK+ulc2Db84YIA5uTPJqzZ+8/D0/7VMmM+hXqXcUg5h
b9yBYu8oGRXROn4o+PbPyzN6jNM+4q0RKEJ/X44rBeFNydccH84gdtqSLzUYmoVi
2Y6OaqNUgDwx9CJAyyfYLA0FkimHTI4n+xUFxLGdP2SsDWmzdYWT1Sw68E2Ewu/Z
n4o3oPy/6b9pium05uo3SVhEcCMu6x9/CUFBw5+VqUdPC+H19lSt2sU5FB8876P5
EnBf6TTbSGhMMoK92pl5Al1EMT42jrJ88XXg8SE/tnyF8V4ChXXWh7n20j89Y2AI
bJaV8NZlCzAYBp8MhmJAEtl32MowSgtrmsoJ3NyvUEE7h/yvlATJPUYq7oGSdTSa
YdGww9GHn+WPLJU+2gv4COMX9DHrrZeP5M9ZyMUV9NrYNTxp8a55F+4z3fbcetqy
1m6xT0bDGHHzjpyRzv1VZxA6Szgu5P4oyqGINbz4INdN+AVzS+LrYu2I0b4xESS8
KVD+z4YEu/yAmX5p7/ZJ3/YFu1Tk62hg+rZIllP8K7FmtoHB8UnDs0q73axbnOSN
U+hH1ctRIv2lZd5ZHqawElVkyrK13G4qk75scpa1TsNuCUqBwndEpJ2dLEkx6no0
Xbu31ayL6XLM8zTN96RY7HmE6cM7XTnrubgb2/jNnA35gZJ4Y0Si5Hl1edDi4M+T
ef4JHjxu2AJDHcIlh4x+yftL3ebKBZttI4VXIOzqeEkGd5VdoNMwiN0ZcrIhsEXn
mqgz5LEUWWvj1i4/VdzeJHo76ovaKoM1RAHg7U34gcjeWsDRynIwz0kdmkUw9+53
GZjcpPTvFkFJP/ZmFcL8GQaaowPI/xSKXsCx+fSm1ECPeGvuEZ3v/Cd0Kl/k9AYy
HXPYOyNqKe8qRg5WNksWUaCSnVRkQp0PQISeRQAWadrzZi3WfV3ysLBRCfF2GIZ6
rOYShaXC5+lKBIWYOXaETulO7zYOTCbTGCsaO2gyfUhKDPmul39I6jOlLL8QjK6U
vvPYyCRGAcAxGtdcSM6Olhl5I+pajpOVKFfazXYsc0gf7xHnoyy29YVE/74XvHNq
7p3Prt5q6jmBDt6YKcquscfcME4SjAV1Z0gYCJ8dv8UqYpboVaALB+EZOaYqVxAs
04hg4hk1zy5hiE2atdu71wvuaYARRfxt+bVO2w8yV24Dwuzo4hODmAZZ9fr3amri
3GvOrHnHgWvNf654SZ2LZ7gIy2pvd8KhWEfaWTDMGjh0/UgmrlVW5ArNVBC0YuJd
utHIRNBWoblHcS9bvEZxwuFXOxIh6cFteugelTMbIxkmO5Q8x6DzWynSIRLKE0Ch
X3JwOCV+YAPzNYgWgTVXO8RBRQ/Lmjl9UamNC704x4eU+QjnOuJMl1ZTeHY0Uv1q
kxJP9xVqBwQ35xNgzV2GoNYe/TiTzZvc8pVjXoUIoFDep4FIzo/oFKvhyHJOKXGX
Zk2fTyOI26rZnTKeUJUPP+jiZN3S6+x5imrpNwPvnf0XDbB7TJcb7pC6xMJJHhIZ
Flo9v/txpe/+Jt26n3c0uAyZIFvNEjgalnNtfGXjAgEJAyk0txJ2odNtOu5IcjMD
Bqm0lFh44y33m+Lvmn0zxvoX7ZZBcXPp4FFTgba/6XZ/WUEm7H/CUHLkXADvRdiP
qDY9AqGbMIDDCre1RBbyO+LQ0kkJPZhg2EkpNwsd0jWT3qHchz6Ye3X66mkYzmjS
TxWbRycIkYdLx7OP0+SVUaRpC0gKg62vOJ6KylUtfcOskMvFi+GIbVygCCznxg8S
H4LZNRArYvLW3/C0NUaVxSze03sR2LseFBriYYrL7fSNAlhaez+ZdTpE7W1k13Hn
s4DF9DiRaKpr/bzbLsOMKegLRGXgwxVQrp3CXWlwmUvHNjAq6hIr526OvpPSYPCV
XYEkaiSgq63Lzk0PIeFpCTRP3rIK6uivGAMSnFsZAAWnV9wkgj1eegiIRrvrp8qZ
xpDcL03zleBrC3k6qPNLR/8YqclpnZkPCTif/5mv6/Rwyv2z8tNkqcP8oh2dE6j/
+02MNcNT/j5IkVe9kXni5p+BZty2W3Q/cvfskotoSWDaCAtMa1zsSxM5J1y6bW0o
pgrQV0oQx7w1DAzAyipzOdK0Ye9zDCCvMBwrfhYjtV3lWKlpZlwtTHoz26XfuFFb
NfWn8YEg1GGXkZfFexxs5xCFXHwJc7LCXwuGkUaNqzpELv+Fdvjzxjdjdlq9mPrx
eeOD8FzN+3b254SYgz6KNjTJXsgsfcquf9qlCbZmJfx2C05KzT/k8QSb/1r6JC0B
MHtBiVhw9QsISZ0CKOxGuzt9O8gZioOBoDwX6H+8J4KqSlfsRtxdOYHW5DThz3pP
dMnPXQSx0ITKT6RG/WWZ8QvV4bxr/jzU2ormAfP6LnjhCUqoaaX5jL/Mg7s+56I4
A0Q1IBiIJTNUq1DBK2uNjrgkwmHyCnirh9N4p0RfXMESMMA5oPpFoOGhUq5XTDg1
a6IO6S2ngvuil/XRVSCUP9Gt5R/zlkGWXI/MFSIm8lav59DpME1jyZ1gRG1qpaKw
Qwa8r6EhtW4MtgXPW5G/BtirqZXLNJxuCbRTzrSEtlXr9iCuovvdWkte4+boAFhA
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WwG7aCNNRhDMNx/vtRrLg+ZfyNXn5sHChDgb5a5ES+ZvhUPFlhTbKikw8omloTbx
TS6fJ6Ddea898rHxJODsbB+OrAp3EhdYsohtCd32RX62Czfo6/zKfSTlyOcOd5bh
BiynFyarG5C4iyiqSUcn9YudGnXn/ZNEkZVGgG86/TGyQ+BavAeXq1cyJ5AjiSUx
VlSk7nnlgutEwYMc188ELNyJMOkZa8m5KOqVfubEuiKIrgz6SI9zVqJae7u9oKCh
v427VeVOCcmQwiPoPTcc4+AipRccxvhEG8ZHfGCEfx+TRYXOvZnAMDvtZUwFD6wO
OzZTHbCAB08VrZKZPP0Grw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
sEXkcj8SDRzHKqyHhjPdCnJeS0s4myC21E4n71IVSBddYtmyT+RIFf3sWWcyEwdW
tPJNu93/8KmReB4LXwzdyoHCGVFig/N0CA4lAelw49v31n1QIpMk61zc8L8O5B7B
rXfJ7xZNIZZtsvBTFGMed62moy2jq2oIopoMNSfaoMDs0tnNRfnvWUKo3oFQIfqZ
nxaI84WSMUuHk/ibt8Vedzmscj7tALbAEBgoB6vm8PIF6YLZSLC2nvVNs8bKcbdq
Z+RDc9w8gHnVV/Rg8oI3skxSC9/0Nm0lsqu15ohGJQ9L2rNuml8aNyPeJK33YrdU
O9BwfidTylxohMUhjBgF2l4IEuTXLMf/SHxh4xHNlDA2XW3Cekv7VdMoF8z/hnWl
s6aQ+Q6ZmmSk23yKMXInYhrSPYyparhDWDImO/WCuZOavd3iEgL9pOWPs+8GwDNd
HtokQMO/8/DFm85YMdqgisRYGUcSYy5Nxj5E3Z47HGxPefT24z2uoOTjS5vFz05x
TDYw6dADiWsXrVCepCer7sKYddkSzGxbQQ0STENqCldgNSWYXYd+X+e4lgMiMqF8
i86fLU8SmgNaVph2sQrWRetVh5bInB0GVJvBGhrl9jAoV1sy03G6XWf/UHGrE7JH
7vnPkaF3sNHkymMAwqnHhmhPnJfp1pGtU5tECfPuRIa1/t7P/ygVigaIYhRciip+
gnaiPafIz47qJzj1luHMCCOkZa4zsr2xlCwHheOkpUUFHEaZaJmRwIK5r2UbpSfd
iHeevG99txf7Jkaw8GZ7JJiso+5qd3HibINZASKAc9LTXIOk3qKuvMCetPnvCSJQ
xXjgt2YK/FAvnbHHOhdSblSAvXoi4bhfkQtOoD8I/Vzv11p/6Jy02Oim/RBm/uDm
bRJMqU2u6lgHI8hpufXnFElo34ktdFzUAYnruuA0OGSGEQNnh+9ZIiO4h9fby4XH
nKjLjJF9/77AJddHWG1sh584QEBZ9IU2uHzjis6vCvcQ/p3k9p7oosuUgAF12aWl
kyfJ9m/UqRfHMosA2lugetDhyhUYxi1Jd/ZompgXkSl7U6hoZqb6qxMzxeiK+gSK
JtWn/TuNEDFTlrAnkxsk2+TsgO5as8AGqQgDrQnzrOGs8CjxBprWwZRC8OBnYvj9
1rPvfxjEghBZFnfXePNfkDuoW/4bfBCyiimWbSCHPDToDGExewT2wNOUTZQ6/sqN
sRmMJ//vQ3mtKS6EKh73wL7k+osB55HJndLYGU6iyRyf9/nut+7Q88+9Wlezr0NW
qgWfM7+TmOymARhUahKiIeecwFbu5pLiuBE4IPWSr0gxOeUsXEm5UcBCtwmpbC8J
3LzmX5cjv2nPizi+AcDB0nBYaCLuoMnvVZpr06A8ohY7YR2KoxxRC8wkHfDQ1qXU
7Le56bgXsPQ0tkMSw2ignROfnrONraUdwXznGrxL9NXpNqtxogOBM6oJ11voQFgs
gJHI9dP7ZUEVbBZcO5LmsrHl37TRJQ/BqEuTNwI1O/yvOK1am/pg9NfKDz2UIs+u
5dypA6KRr4pE+KWW2nzLvlPp5YpS7LSBx1VVeqQ9NyBH81qvZn9o0bED4qzKMCu9
L3NCn6NXsXcIeEawtcMOS4828xFWZNgBS1ACELWlDHrTJvm/qc7g2HoTjtiJzLHv
U0+PQfyZLElrVBrkaqIp3ulZxIBHaDnRFD4Gd2CTKQ0WoDaAenimTCyTYPFh7h37
RX3tnrxPliZAVo+HAhB6tHCdLuP5DyqjRgjVUiauAslIZmsuc5DBy9mPB9bbW1sE
k81WjOKInxmy5RzT96LBtmg1gP1fpxBFaC859Thf+M5JW8SVOtCM3vlm3uN0bT19
HEZnDKzkIAOSCWSOl17DgmnllTdoLLqpBu/6z89DczO8BPbA58M+sw3mqqhnMVQj
Zc6Qa6yoe68JapR1J0mXtlwExrLmbdeG2NONZrKhkYkyn9nQxieW5oGhbBEphC8Z
SWmfBc+qI+DmxU4y1+8H4kNb237OGpID1IHQRVOoVFfI57+fmFCcnIkl2tMx2KBy
QmGh0nqBj9D57cbZ3ayfbWbQI5Mc+So0qG/QaCeXkxgjGXBerfVPihNQ30Nk5t1N
11BfvYgqD18dOlL9ecksTSH5nWNEm9PfLWoWe2z9OULsLqFrbIuU3ne64MEIbdbf
VpizAc/LR4E8MUP1P/fOa4X1DZmVfj1dFgdO8eYBW87H20EA9893p/+sAqd/0qKZ
mwpBD1UmxLaD9VRB/hl7tcWOArwb43VUp57YxGOaLzgBd8upFYcuZy/twj7mSuWQ
+uV1otONp2LwLoI5FQWYzqom/YmYveFHJF9wB66D4tUMKB6Ps3Ds806YPNbidrHf
AyyuMZqovLH3ArvmBO85VgzEYntS6IMWhU750Zn/nHULqjjAu0/ZpIPHrRlMJjdI
sWtq+kQiPPZRobmpMWfb7pnkFHtLyMVhI4N1PoTmnOzRvOoqK3qh6CbScNqodDI2
Tf1lG/kKfFrp4JvB2wElmAk/TM9uHsBqTGV2BSuOYvPmFmc1hlE4vIhT7vy8oLRo
455npBFo3qjHb0bJmbYKYAyj1bM98E5tV4G7du3e38Bz1ZlXvlfTZFBKY+unp7ww
SAeuDc0fCYxw/kfRfmjnoig2Yb8u4zyrEqiWycI9l2vbyxPFCqYJi701LyJ82HxQ
rW4qruLWf91bvnJWiYGSQLd4Q53G2I/WTsWATJqPkM+vEPb8CWo9AVN1lrQRGyqh
Z2M/9MvhF8iiOPnAOH6UlZnmNIhQJKIVroB8k14jh0sEmZ8mQCOgDOsPO4j+pwbh
Df2umb8gyxqccFAF80hu3//jU3R6jWSSa08TxvTafot6nW27Lg06Rd5ORCNqbo2H
TSDYCW81CTJRMap1/gETPHgWMR+xt+olNFR4TKh+Wgl4dl50joLWlAUqz+nnPm2b
KvmzbUQ0lczuOwYCXmwXcBuBqeraOsy82G3eMqo1iEHzb5eEp4PZq4BMLivQ02XW
xDWDZgQGKDdrGHVvkP8i3xIwHctBY3ZueVO0IuL7eLkqNepTqVSsQyV7NivDiJFQ
lMiI69cR3hluzviqly9EUT7RS5PgHuCxEMx+cCC1Si8Vrk7DWKo2ZxOYml0521su
1bmLeFS+g/alLcUW8yJPHEf0BzK/YgJ784Zobp3KVl8yR0j1fzH0ivXnLOozL48T
uaNFrpGfGTZLNhkV/kM41Bdh0lm2oMUnFE99pTNq916WWOWFtGV4iivB9v31sAwm
66C8XO5a/ocdKi7KJc2k5T8+iA83q4lJ2qa7S+UUh9J0AeLB92FQVShwEr7wW8kT
nI6eIuRJ5fk6VRiCvkK63JwRREI4BX9fcD8W9ctxkQBLbnJs44t/d1mMxt4CkCwH
PVWtHprJPwBf/V+itBD1igqqSuvIqiQ4dk9xe/zEnJ/8D0B6k3A7gJf+549RZUN1
ih167Lhfou3hNNTqoGay49U1o40jU86iysgQCex1HfxLjVGO97KcDpPDa8gM/d7N
rBJdcc+PLUmZpBcGoQMx/GQ+GuYcJZngaqt+ad6/S7Hubj/6xzSRft7pgwhy1/GR
lRbN/n3X0poicFwheUJUolxxi6p30Qp+kieweBrnswqV17o68ywUijRFQPByFDoS
BA4M5jNn7nWqkR0CuZk8jvouaGXggV6NeQtoZdMqoFsLQy5YTtn/gND5AGnjBV8U
3ovD+ljYb1Nb7tro28idGKCWhAN77G0ka/IyCFVOU00Ao6lmo/zgp7VOJ/xA2urM
5XQYX172ldpxxuuXneoLzEOK8fgC2NzbbY6hUCid+3eK1fR1bXoI6EAJDsxbOH1f
05w7SJhOPRIGwLSeWqMH8fbUw9KjCt5imA5/7RN1JBp3KLRCk0CoiHlgyvx2Zr5x
7CkggO1Kz1Eu8oPAjgPy98ugmlJV/Tq7+FLdk6TWAmsbdIsqq10j2sTwysrjSM5e
OnzniUTL/07RcOHzXxIIr7H71YdrBmqU8yDKqfN/ooRFB6nX0KIFz4s1x4IwtVEE
/8JGOo//0jgXphyusQ5ChesoSUN2jcXDiiGwvjJJTwB4JzyLHbjxZgcgSa/9L3L/
+ED3cScG1GqsZAb967ip7y4qzJpqUfTgrIxvol0VJNYj+NGJBZZv7ySkWMHQ8ZN3
rzvOWCRIJog0PBoFyhLKMZiJuB9y45IosF57Lxei9liWy9/rmZkt1iirv2gMNmIk
dywVzL08Go9+bzIkHadvu/bpaI/EVOIXHGjwyFefp0cNkaip66HUJTePfaOc5rW6
RPVjkATj4ycOi+KCwCydyT5iYU2UKJVOEwxEx6h3ZGkog3h3yi3pHdg65S2TRWIs
WYkyCSEEAMoCLvWcHSRbl3uFNJjG87GBpP8bldhZaeO57nc0JlgPwSo0AJHX2t3w
nM2Wh9RDWd6MQd4UhiUnb4vIkoS6KTeqvWWCMWiiiK5m3g1KGVBIU0cs6QEfTNVA
rN8CRz+wvUVCQDqQaKunbxOB7mCJAbQnVvTP+QdhnecVzK/s6cHynckWwXCkyHHm
bT8ZE+OWqbknmpuR4Ix/rw2iSqMlDmnoFTGv3Zd7BlGGe6R92oAbrH0rS/TU1d0N
gXF0Fy3LtkB81KwpMWgCVRCkxJhSAuYUx674cSdGkm8EiSoUxMavBSfFFxVIvXtX
WrLFb+ixxENlyQFoL8lzB3hN3uaeUc2PCYLmArjSt2gZtC06lLBUN/wVy4Wg5dB5
uoHySCKxIj/dgyeqVOaS1JzImjIRcWLRRz1qbZUGz7qfKOArVoco6YnGZG52W6WE
Havr0fc2BQbLwgzFwcKGQz1BgeQkmGtSQEjAZjAW6HSV7hVHvQ3FKpeD77tqyG/g
zEXYO9c8vLMc+pKVMNkA8knw48Sft7BMothYZziOKQhGj9Q+gp+rjUdpl5ezpCDw
M6HbfWgLESNqoJelRZBo+fOY9OZXjgk+4I4MDL522kOg7RHTEHE8g3b3nJUmiP+n
ci4BkSFYYgl1fMSPNBQxa3axAyFdls8xNt0wS07Gtk1B3h7BeOkPoLmvDg2NeEtM
2f4CY7PVSlkits0wQ8Q1wej9T2/Fve4tB3jFWmq6eJONxI4zGTyUSJXnVgk08QGd
mRm3IQu/tGgsiGA9K3FsKgTCfotpWx+tESZOgpKeJ4GJkKojX95tGXprcHDkBsXX
I+3EVldWNcS3ffl8RgP5Smza8LVlJYJsiEuzo2+JEnV4QATwdfTudTock0vpSNdc
MVbcYtT2MYW1CHAZZBrGxK/ahGHI8IzUoCUIzDpPPZ4qWEWu7A9n1taEWfUz2Y2n
NvL3saF4Mlj8WkTpr4GTjecp5daCuenQDRDp/diG8iOqtMOYfNcY3vo5/NAfS/pJ
l9XwZhcSozxs1dQlVlS1koRM169YPzU76r9NcE4lzrTEN51MC44880Fepdr53qVt
C6r18W4zvMyjbEgi6Ix3rkpbA4fAYNsYZaqfnqsQSNtbcc857ITehuJrFhJO7Lz/
n9IrgHCM9qJDVTz+lFILnX2tTkat6MVX711NxxTojz0FAB12QMq8DO1lriV7SBgQ
7iZGuYWxS6bDNu9rNmhVUG/ZNr3e6bO0QAlZ9qfzpKfezLW8z+CiWT88UrwpACt/
xNzx2l3gaFPojEWP5AOy3xMn/ZK73h4hsbskQZ04fNNAIPGXMaVYomyTsWp3mzGb
HTr+y73XbwuI5oGzAxRqrYwMkNmG0c4su/ujkg/37/vaidwMo1rOz3EpCYnefd4B
BWvjfukFvatt+QXbd4boisDnwll0ppiv4D+4Ayw/XBzI/yBI6o6cAclzGcvgswkk
CDN1HhDtioDxrSRsAjmF8j/6Z81CAAjhpw1MfWscnB53Xy/1fY3HI7LjXU7pVpBg
JoNhDySCw8E8PfPvTj8U7SKoW+WdYrhSYeIs/oeGpvWsqfTBztNly3U8Izwl5uhr
M2Qwp63QLmJTQj1oBPyjArcLwGSCO356dCxJ6NatKSXF759uyEG1UOTn81M2WjLQ
ithaUx6n/T5DTFhbYDw5zo6+v8q/a8MFGydcBjzO6PDhanVJNLDWe7oAXat3ALOy
d9NepgLhSyjdfdR37pu29QP4v0wD16k9CPKGUiJ35R0/EtrbdR4Ft2qRVSzxDge1
C4gKPb120wJiX6OXdTHNdAe0Z0DVkP+roOzCByyfSsmMSJRVtfaSPQA/ogdzpogg
zb2rCiJybNTdun4CGTx/Uuy0E/LGtFjrszjFicmxTWbpeYYDho22CoQJjJV3KsHB
TYJqwmcPvrfTX4woQV+0BgVA6SW911kGvAMyczsyE5VvmfGq3Q0FR7UvO+MivwXu
YFPBMkfEhZKqitC8HmEWz5S8tl90Zf+E1nkw2lrY74PicW2G1ef22zbYWU5EqIoG
BcCS44Og33Bl3zBgFilOkmVIegamlaY4q8VicPUlcuLWjxEKi8e0qg5FqKUK8peW
XGgqRDXZWwsiYGajp1n50JFnoKwwSt6+6vqvJwyYBV8ZNIsYC+6LAd4exznraWC6
JYd7A/qbxrvakLyI1ukaM0N+ckc6SKbbJOPkAe0Q2CY38EWyCw4Jyv2oASkFK5RN
GIm3Kg4vXzgCaWE6//ntAMsAcq+znr71T+v2PJ6JlQP/QVGFWpAIN7Q9uLMBigNN
v41wthhLMTOMfj087yJA4qhcH7va07/De2ZbaycUNTF+jUa+t/T4RTpCXljEz3ld
cl+gV6AiWuR/uB494ftO0aQcw8kAPiD7lSTOlEQ3K/jcDo34RGUASygnn13CMury
DQqxkuHK6/OPNGOePzk3q1Xp4hAmPaD6Pd/k3Fuv+V5sA0xLbTGw1gsfojKJIsWy
OMpfk09FzNqnp4y0wMUVkPQw+87UfW2x0AjtmuYWt1k+ENKX4x2CzIvRsEM1P7od
apj7BtAeSmGJMEkWOsaVbflcdyhcsGJd1fwEsr29/snnTztukwssrrLYM2seCDG+
vr3V3Lvi0DMoS0ycYeldG/rd6xv+gjAJgAhGHxSuaNQ8OpA2tOJZa6QnzxTIFRL+
XHu9lxJ5z7xCt73Iqgzcw2Kvv7E/6FMRlZ/UE/6JbeolRfAmN8iq8CrkpFoTANPj
OXjwNTmKa8YMMl2hm0/Jj0F6Ho8uNpvLf1Q04rzAiYv+hTF6slZleGxV8tHEXFDb
wqvdC5s+szgjlop3rjwaRJzoUAp3EUSigKgncDYQPtTRau29jvPKvk+0XU+rxmep
0GVsCy2IyXHbLGSK8Sr67ujQ28ai0736BrRcaFFIg8qdzEn9NL3LHDN418TyUiqM
iE7PLtTUrpSJ08jAXIRq5pTcbznijmEk9FGc95pC3AYV3FRfG54zD2Izlibn6SQJ
o5JA/G1VWvzt+9F4Vt34LwsrBbqBEUfFHaCPe9/aAjm6epTlmH2LDkuqcuqpf0KT
1OAU/krP6hfnm5wCnLkU61y9Oph5VPcG+LP9kGLz/9EmYrIGUSDT59fE/WFbHYVv
nlqqUuZXkN4AWgT1rrOejOc+75zCmNSGZ10+FM4K+zLVarb44n3jU4f/PdsLtWLO
CA7WdeDHpNhjJdecRCM2Q3LCPyEAEn5Q6088YgmxTaYrmrCw+qewR2Vd8zYWvdk6
XTH+jEje/3Tub+ODlLe+hboIFvuhoy4urcUVcaUxCg/gBYFh3eHWeiWctJLIkyrC
hXcvFAfeIcx3C+hSB/S4IQVpUm4PDP9qD1tqUwRgnxFPtc6Owc228PYYnNNSnP+c
XZxSGuQeO6jWlLE5DSzp47Y42fUAP8Kq+rn0829dbovN2U70v+qdjfA/VZsdX9KT
c4TU1zwt33c6lE2bd5GfnkyJviF27RdGGZyc/AQ6bUgeBG9Mi+hB0jotzt9vHzzo
Ol90ikb3dOb5PbL+DHurtBHhBADK/tUY/wQk8I6A47/R/26g/gcP8CG76ezETq7Y
twyyf3+UCoMTJlH4lk1pRB3v2un6QbpFO0rIDo8Bx5z4799+Nss2ho/PfeAEfjyX
N0GxSyRAIea5KQ8Fx98eYw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
D/h4doCkPxX+DDuiBMLeZN0p53bEECVcUQgTnjB0ttlhvpWJdrge7f0gdexTHp1x
SD75ojXUIjJoOQ8pfsYf1qZMS97dWi7GlYxc9TXvZoVMLLhPc6kq2IzWK3+6RtKR
kM+Mbmftui4lPYlopSMKeW068iWqqPA7Cgo3jYbvgg5VY6SR5GeCiD6+QryJQ6T/
2dViPnFK3KppY/ohGieJcPX/8WHG5xpp3xi/++qbUJyDy0tvtkA9NM8itn5r7X6A
0oaeXHK/VwEyBNbTujfNycw8KO9rKAzpSgvx9XkWjx4PrEOPdvNJGsTMhkpy8hNY
Z0TJbhrr4Wk0rXVUjLgEZA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14480 )
`pragma protect data_block
zNmQLqs4nxEaVibc/YK82XxgqdSDl7tpsjP3I4W7fVCmju3PThkCIrf9kwWJqkX+
dcrfmiHBFw4xnNBhuW+5/6ouD+qkcBZAj5H5RJxR3DNCxMa7/V6vQtKJL4LULZrU
s/+JszgGMAOiSaZDEgC7etb98AZiEFYfSvZbUM5iuksIoAYI1BzU60lBmX3Ju9Nr
zP4kZXb1PQagIoiOW8LZN2Rl87vMTDXsMzPLBWJnhs9ikaAd+0pbQaz2yXvKwTLd
+iJTLtG9PZMrog79ppzyXzDSRk4uTCmOanQIwtgHZJuEF1s7pIlqLXtjfjDiuMHn
YNNjnSUvQIrdfpDZqvDHEVl93MUWer233alQEhA8X+aDUTTHk1a2YzpMwzkiyzgV
0pzAfQshdm3xKIBIkkVEv9+gRVKwPF2FMg91Tbgdik6iZ2wkYvzuYMgDmOZdDDYo
mr6C3R8nvm+5mWt/JDrIULik+0wX6+0xstRA1N1iTZvqxfa4guMx4Av1aP2HmjDv
R3EWjHnxZ3U4EFfLA+TvZbAWLzsbB7H+vJQBNP0DpgDk2d6VztQLT/Lr+QsovuZZ
B/PaG+lUkFuZNg2YG3naAu5qOCsN8YF1XqCZShP21SEUwK5Z6QomCF8skhKHNHCb
8uz0p2/OY28q1PRqe6+v5h8x2LpPV8YLZKlVUJYjZnAn2WDDePuJZm9XkRaPA0WU
9dWSvZ6l/Cpmiob26hKG54iRfh+qHUWL29h3AG5Qj1+HuJECMHr2a/k/7SRNZD9w
cFkuX1mEIeIYptSx7TFigEyyXJ+l8MFocHJrvd6EAHCN1dNbe5v104iyqKkQ1UnU
D7U9knwuqZHi1cHfeXMt3Jw1pYbvmIQZ1PdCtMm5tQocD5QFRk+0jo1bTOTQnFr0
3mXVe7YG0eulXshYffSTzGKYqOo0kCU5wxV1gfhN1rwl/ca7AuznHQQPzmhSSNbX
Jvh3A0pnc3GNmypmxw4oTKlIK4UEm9kD9renldNHApIdKO6NAciiTILPr0zsHBs5
hXnCi6jKctYwa4SsBDO39495sGTVsxciZBl0x0w+SAXLAud8+2XESTGHBfPkBnJE
+KBShwp37+qI/NBsuY5i14PlTcKqVpXusIRHsF+71XRzbx0aOBIMKHhl09/WWidw
iupph2134ZYoWusbB+N4BUb3Tvy7pYFr0G9Wfknr1xl/GodYS6SEDc7QTETd7rSz
r2wLFe4eyHar218MLZNaifZZFatkTR2Xp7KXPuqspjSX2+OpVdmfK1ctjBWxyHbZ
AEqbH81KEa0fMXO4fP8quRq2F68BOeCuHwt/g1sDRDbuDuHtOKTvAFZWMxlu617s
r+r0De6iO9irwr5zdRtrNKMjuQqIOoSiekBig4vRvyxtX9SnuSe+/gq8sl2wn7jH
wJa3yITUZcRcC5slPFd7/haOr+AqPv1tD8Fq5lRXBzUjXfVWAvoGRcnrZMhzJ1iT
v2TfaUrAhn0tAfrJmBzjvHiylihS/2W7nPfScjEX1B00U3xdEdE+A9MUVDB64MJQ
2CgkihVlVYSeGnGLFIko22vqN9l4EYHByCoT1ZQQBIh+bWwAv1ewvJpRgJYS1yqh
7sMyi16knmSrS5RZ7x3+Vw4ktoRibB4rG4lYW/lsGA5wh+jmNDpjhjL/IpDrai4J
M7WqVMr7yRNDjujmG32NfOCD/c6rWZOvYVuMAW/lufnOYRph97gUwMCvmQwadWEM
KpTalF39TAkPrInc7rmuMud6EHU0wLfAUlbhD48n0iu7H6mQRK3UdofXtL9QwvZO
oTiLmY5KD3581C/STVGzJNvSRfKgt8Z8xHB8zzokn6WvnyQNYk6MllLuLQy25wvS
k8HrpThjDmKYIJ+Tp7syabTI/2BzmuFXf2AyBQxoR8ZH2zMiorS93FbWoCWGZP9k
XipFXyBt9P2qXzrDhKROsdzpPPWui4n32/kKGusJYQoYNl1GrTgsaPB0RvHtCGiv
wB1z12r2StQa3TB/Vr5T2h5popMl8GRl6XTfKsqpoi8+or8whfGd/H9tDtc8JNhL
XbIjS30MQ8BNhQSDycD4No47PZbAx+XTyHqvcvJfv6uITyR4BhK51kYV1tPiMGwQ
J5OJR+UlrV5CuwlNsH1jq9mIYvlKxGjrOY9I04USmtFHW/Lqz1oTfDxlPiFnx4MZ
Uxjrexs2/tp60M5jp9oeD1JN53oLFgvjtGysUJqY1GWxdWLjTFWpWOIAXhwnl/4s
2UKWPjo8WOFvYvEn2FJEl59tKKnHy1AbutAKRNQjuraj5OOGHs4OBcvtAi/nfMAO
B+yhr5duxkQj/WWN8nKGioHVQ9+cViDdMRZUsNMyACJrRFLksi+c6gNE8q7L5+zI
u9deUwGm3SeEBjwcVFJdZ/yXZO0oA97vq5Kot1P4AqrWSRrfZ9WpxQvzn7iG3RYR
+rkw2Krk7Z0Wdd6tdwPciV+zv4853llGzrhEdLoX6jPesyaD3om+o30FeU8R8Zmr
hafR0tJYsUnrA9iLr+NDPnfvwcX0/K1nIweHsJWhrurPMS6SrzGaxh+VeJQihX9v
vesDwGn+Id0u3fnDtyQbPyMEM1uHQBzNu64ls2nhBWSE9h+Xz4nu5OJUibJe7g3G
7i4ZhrBRd6f9uwSzDt6Rg7PuAew02C9bkN5rDTjZeg+fOAb3yUdbZCKWGhgXjkFa
aeQRRR+UcmnwmCbNBItsj4sHDAjRIQC73t7oimMDR7Z21Rl3abCLO34Geor1QbwL
SRTy/9t5sQJPHkRQERH4t3DtJHLCJ5MIk7ongsnhLCStr9Dxq/gXBGBA2Ln2vBPy
aDQJIcPe1yiJBbPJBhgbUX8zqcbV94JDP1SjPjTx6LErxXoWftryRuAkUVPqDPQx
4UFjX/9hvajsvl3hb2eZGp5Rb9E0wWUUcuOJjDHVvGaKjYIqkl0TCMzxFBT/FmY1
pknIw9jk2wEFzYEZ8Q4alyZfLLkEa6Pf8ztCrfJ8CU3UgoMdfrCIQLtlfkr6X9M8
Aoe3op8OpIlCLjIZqJvwEitKej67IpiuKjLvqq2ycK6OBtvP1ab7kKPelnNA7pxI
M+12OiRvtKf9jSFutBSCEyTEdyqU2jlS0R4dR+HJrbI6g7DglfEAY1CDQPnR0G4g
HG8mjJreIV9/PXGACMp948onmuTO3+vwcsbp+/xR90/fc7oW9EWv8p5qWxYnK72Q
eKPuC52/ybdxUXkkvqEvi6NPqzOtL8FTWweJ8Bl9L8VrDaUFPSYMauBs4m1rQiSC
rsbW5zGgo50ah0xAQE0LW1cOdQjafjSEs5BKZTUEyYRxvGlYOazcC3jaHjLan9Uq
mByflmulyAwbubuhQdQvfwE1lPnQd61oYW51BLxT0fEWSkxdOM5m39khHI18YZv7
wZ11DkOUSCNiWu3vECkP2He4noFRIHLXIr+sz9DcmLYGv6irszS3vxTH3g01A4gC
SN1BvxO1eptIjA1jF+ZrzDzz5s4M7FFMvdePae+13qsJ55wqr2bJaPC3U24Tt5LP
u1yghreU/OBKDNDiybfHBFaRRAGm49veeUr0B/g0SJIrs8hyJ5NmAYIIWfxWktGU
gHu5fL2be2WHThiJ6tUO/j7SI4SFa8BVEvy7VCYOxE0IblXJl8btQBlRkhUW37ZC
c+2TLiWmDF4HQeQmtYfOFNBjmyegAmtPGfJu82vraQDmJqhPk3fsEjxdvXouVJaz
2qDBHK62EK4Pt9uuFhRKNXj43JextYo5dIKPCAFo5Cvq6TiY6z8lX7pPC7BqIn4s
hz4bj0f18HFDcN8kPzr10rjmqB7G7kqMTCzCdqmeSkpLg2BZNfe2zQabuLN6RtaZ
05O5cuOFlTp4KhjTYn6iajLXk/eUvdAbbbYNMphS41Bc+QRCzxrxQUvseuhkcdEe
O4qY0zSPWUpp/ua70UCi7UwTkhnUXe6Ab5tTMLZfIADoAHEiN+Q/rQ7Z8WZas945
ZeqoJz02EaBxOEOr+QpSPHgDemR22hMViNCXeXELVCmLslntgvxmK6cPpSfEZ/S7
J+Yqm1EZ2hQ5iT6fdOX+0SjO1a6m6rLBKY23N+KUmukHd1J1AWFLK/BTRfpmp6f/
aA4OqWou1c2ZamxMeJl8sfVySnZHIiH+c7BhMqLhBp54kSPMGJHVO3IqPbMD1TyM
x4mh0FhC5FFGUVxAUTCB6OwpmV3kgtgX11At3dJrS5AzJVUCjNeAgpocvcTFnI5H
A06CFIE5xx+gMqQiul5+N6ShbDFqywImImi+1Kzt6mxdBNGzJxZEs2+SIl7zBZoo
d9h8RAb0nQiHbShYnDC0Urb5Mk8O9BOJ0/sjO6LjhFhoxyRZaJ7NBXGGcs5DVJoX
oGmeCO60WdiOm8yyMjLe10k/+g5ITAZIcVmFNkdVpfZpMmxtew/Sm4qjd8ExkeuC
fzc6pP2Dk8OdKZszdG8e1noyaQd7r29mktP0DrYPm5Zp99rJjo0nIazS2onOg7YV
ggpNQk1G3HFdy22vJfnpAjjq4Rr69GYIkfU+HMkq+S7RjuL5FeplzsRO8m0QOmro
8Z7szQbnQK1BC/CmzschclS3GAq/rF+yoCiHNYgKwIIDfxCUEl+VxVmBlLrDPVT8
TMVJwah2g7ZttT5wokQYt0E5IHENIYqrhkdVWJV73tZljnfylkEDOqS/s4MFpxja
v5IwWzCEvzPbDzxhViYXicmKYXzFXi3a1zu4rKSusZnA2XLFo30coVt5ZHTK58tL
Q62MACBP/zU98M8KOSlWI+s34F1ok5Gcw5uC8fj6/9WdGPLzh42Vtx6gJ5MPM+oc
1Vf/z1AnsfPUNezO4OY0+be6AiuIbV+I3rB53gOoT5BqaTe4qlmza3CFQUcali1S
LA0S1TZdAS9LIzlfboDnXkIXiDbTyWv2/j+reG2PZq0iNoVQ2fzdZUq1rSuiRv8j
bpoR/BjBvmyehw/RNmZF9fUhgTwQx83SwPTKc22bzvJ8dZOREU2CPOSter5a2jui
/gQjZrYwPIiF50lg5rxkU9+52TB7g5J3r/9R+6k6CBZ8WvNlMFkI8aciTfKaGjWf
FGVXAHEymAqiKv947O/muk1jnnCFG+n6cVeO3xHMPel4u4ng3MkY5yC0btmfgWcs
f28VFmbji0xlvTtaYj3pOb4c1N6ycWjZ713L8XKD9zQ/srUIm2+RLBsrsHYoh7fu
u7J+X1U1W+f/bsj0mpCMbzJlO+whxWj/eIOSSJ7aOlLeUQpywPxk8k2HmPbAWFxF
lvj00u3ouVgCFEDtMk34/YmO14s2E4XbaRlPIfp5k7IcvZ1eZ5VUy126XzhK9uIC
P3t/SJ3Z25iWc4eVU0m1CqVrj+TwDvhC0dYniHREzHlGcshY2VporncPw6DNS1Wv
20758N4pUYYekVnnwDv8/iOO3kaOKkrbA5Zdhtpp/dyOicR8lSrSPW9Xl+J4EoEK
cvAjSqZDM4sn3/dyDAn20TWAAtIQ5srf9RB9KRcRjWht391YMtdlhm8xDumn6XBV
zjCEtMHmAg2hF+0i2uH/jWyCtM8l9klafDrXHdNl/hqLTskYGA4F8yQ5+B99OvCA
Wlf5URSn+kWaIrupKtoor2IBCRrnjjYA8dDkqqlJdL3E/wVpxehzuOZpL2mvnt/M
ZULE7m2G/mKCYCsusktH/RIgP/DPZHdSar6az2g+eALw8BmwHR0FVzjX+vESFQ2s
1n+zGvWSktdO0+j8MGdc+Rwn0i5u8DRoFbxfe+jwOiDPm+LOsATAvAafXmY2VORm
d5PP6g5Fcjv+nihUaKOHbu0K+hiOGyXunnuXVr2wtKTwKxo4fg39eWImw25wR/zH
JYEfXwWwmyK23rJnTYV9IzIaLmAw40MaLTJyvXTgwV8i4tV7/wPAq7N4cwVoem9x
g2pNDGESRjjYUivJx3YKg6pt4x9x+96738c5cQ1S843h7Yrhw5kf2cMRpmcZyvJT
BqIGBbckJfwBT2met1rEg4JHPOxZFrSPboLkJLSU6ok8geu2plgzdGg+V8CgSr77
bZyRm2fE2YtyBd+ahNKlj4xEtvaFE5kfC0Y5Eon4BAcSxtjSpZv+8o1OUj2ctPjr
K1rBPi8BpO1O+KkEWSkSIDYo2+XNF13yOKR/LlXgrhegDKva1afGJhHRGU7P7/Tb
0fU6EYw4TtccQ7/VGwicOtRoceEq2LydnL7BrOt4UQW11T71jblLpu+n3a5E7X4I
zgvQAbfxI9B1gZywnNzSzeDtWWW8fKLpqtKPoyIQc/N5lVYJz67RLlNmFkjxRaOf
o2Y6WCRm1SJp+RO4/OQjgcpc2vFt91L3vnC6xYKzKEOls1DojUjzDcd9gINbwH+H
5d7KjGvTzraCzGbr5WLPQensa2QYIiaOaNRKw9IZXcflkqJkPQXRAA3V6aZYrCYv
yobOvHSbVsH8zxtJE64z3qLLSfvTWG8mszb0/l8E6QsENCc4pOyVRKyeGCC/WU1y
WeqTUlkwvlw3WdUbt2+91XUb4jAo+aqbfzK6N6eHzQweJg9j9Pu+ZHHkgMXcBpgm
XbR0Ffm7KOHjGEa2EiDOI9KXU41JF+fdNabaUXlZEiTfSMcMNy88BOtw7jTVeLLj
6gpptgPaGrhEw1nvQijZ5SDNDE7rCd7fIS6BGrDmQI4gs7Zu8NBy6DpWdte/Q2J9
bxCmdLmg3sXyC8hfixGRmuOFTQpLW8YH/8xCs/qMBW+s3FLMkA8q4Q9hTztGh1hg
kHJYu0aDvuDxXDYWUIYfgvi1+gNZvlp0CK5gsxIKu6/zo9O1elngCQrZy/84B3wZ
5oHZNOpp19NF/EoNAkA5vGUnL7iF6vw6gAJVC7kXDvX81hgBDI+LlEEQ4UoO6wCw
Tklbsx7HZoiYzwBsl05h/8SsI91I2kao1fVNCJwfxr01n5ocdakWGkjSPsaMQcus
x8Fl2wu3x8IjkmSoLI6n5/ImTxPNSxhDpVX6+kGXqtz+3pdEHqq3xlDcuD1CpfwH
SU0bGgnF89CPgqiKJyTEVQjA9wD4C2EjWZZ5DE3TRLpEW7XYMh8NleOQ36v9ZpIK
epjcHDAEVztCdAIS8Te11KxRggOHjcrmQSTNsx/CZ6Q/mSOcpklN6z5i13n8gSuU
hqarUZco8QPl4sLWN4+fM2Ot/ElsrfJeiczUfIfWQoXCqhbzzv2NweqxO5xG/dhO
VpHP3WRnchEHEQIGcYV/SR/z1X2b90F+Cytv4WHctfKssls518b74ziYseNAiT7d
Ff0k/KgOvkwaxuwdRmJEGna+P7mGUqwdWUbCbm/xSj+88O0hde7IcWR46sCwxaIV
cpQ2IbeOSmUh3ADwsMnDHFrGfBlzqX7gjQmWz4j3cMqYj/dBg+YUf1X9GS63DWbp
DkVrTDSAV6KexCYaUxv4znXdwnWd7QEAmlf4rkOW/L5J/AXSsBg4E/72p9n+QhJ7
dH5FIiISlQMWg7N7okrL+NP8dqbrLxcLM2JkVQ5iF/vpHzbmKdYLT4j4ioCtdmFa
gOW6o1dphBVOkcmOFEY/uV5GB67SBPY+OU6VDOLq+qdFETluL0i6DhuMLCNPO/aL
FIa4xOdyC3L/uFewoidRzys3sQYMcHrvnMHMs8UYEHWpGsFFv5uRxIFdRvoIgVoW
3N8w3T9WuVWI5OqH4+gWDxkyyUq/kesLdj+rwqBrkT+MpK8xqUK3tYgqYF+6zeq3
OavOh+eITZsSxEobypkL1+tAFuVSSKcnnLJ2JBhFoKsTzrHIzeRGRRQjPnAoVUF1
PuDY5jr/6ZftfIyHAxwmZ708B8Vv95egfq030gkjiVcVa67o5aQdEstxcJV0O9dq
hcDaxTFkLiiRBAtb355CCV0kPHCRtQDnxhQOCLo8codqcQDDAbc8xFa7HpRhaMTm
/EWsatNZjt9haw1o3peq7/6zIODPvG8LcHuLrL5aI7qbK/lfhlhRsJjpjcqbX3GH
iJ/X9nC0hqGddkRL71epR36BWASgO0KTozv5Fjls9SlJthIkOoEWoahnKjmrMJne
+qiwna4sXEJ3b/jRYqBsK0eNvUonEr/OtR61AvTlnpmVTgW56jBr/KSp0mMQhCJk
VUEwxWbQwUeDIzOToOaqVN0YIVOEEuSL1gihAZtehsOaai54kmmDbcYedbCQUJBO
jqPLXxVDSRWc+uh5/X378KpfmaPQAD94ABwFLRc959qIBaPkdSpz4aRhq4bikBYW
Dhc5X8lce3SZmtk3edUQH7sOsqyBzNLSowIWHT2+XfcCYmFjTu+IsCwPw0tVfTQp
tNd8EE8ZgBuFd3kiDUutXpaRHHBAOUSBj36P3d3Erz7RDBDgdKFphpYDdsfMtXMt
WAAH+9hovnPzruwKLyvMdy54sgZlwuF+3AH8hm+SLqF/zSoNvJtkv1oQZMeAm670
7pbmzeLXypd5MWVYDYYdAENVsJRI5LWtasVXLW0D7NA6OktxuCy5McFAFXvXCFk8
4IdEtx+z4GhyJNNgP8pbvhnb9k3oMwT3Jyo7Sgk5x5guT8hAz/4yoABbp9XLks2t
5iYBhTR9FAhEj9tqnFY+v248p9rQzSLW8RBV9zIgVJ/hVJRYg+vHC32/FCoJHCve
i5bH33m9MspLt9bgdAkpwNwLRWj2UDVGEbwr1QB58X2WO/S7UGb8aUk2XlysDLJV
6nhesMjO2IOmwgZnVbdJCI8JWlH894UHRzot28UVXs1qHOYqC3FTkzorSxS0d0bD
PgxU/jZW+/TXJth5/crRo/3A3NVHDvzHscok7Qm2xVQKGOTn12ukGiHgY+p2VNMt
TjdTh3B5Mb6KtzeZr2mHicns4wW9cwYotL1Zwrs3Wwssd79DrJFUISpA6mkCdMhG
KVv+DH3V5bFVUU2qsVIslPXQBlPwwFIk2fDSF8xqewQkYBs9nb0XG8e6cBaNi+VQ
Ma6S4CTF9erxSrO2OeQ2Q+I3ijAESiLWOie/Nx/QlxJlJIxNpApco0dJtWDtSkUJ
swIkGrectDJIHa21jGOxdaaYa3b7yYOcjhua76HT7YJzwu3KxUJc97rYSx0qmh7T
tLgnzs+3UVjUsJ7C6j79CIRVvgGro4+awQ/qiMQ+Vcz+3KfvTct2P0/WljuwpooJ
n6Z++b5u5tIw5SYH3cjfe561vfGSiBugkMphKXVn1HYgYrTm2fuLo7qLcWX8nESn
4DptFXFvW2CPDzL5512puXBRFujnEmZhDJmUdcADsWWealJ77Di3iJ9GUwXYAoZG
VpR8+0+WYHBRKA4TtJaYYPj0ubaATW/FIU11kfFlcqCNhcm63xV10PWFa+Z6METp
s4/VZbKrikTcNHGGXI955Sljea8/cBvkRN2vMjqW5hbhv67BS/OFSwls+X87eGjn
yAQZdf8+srvMCwYlXi4ziP6qLCBLNTnm9ajweL8JBHq16yiYpLFLc4yVJNW0gsWP
2Hwg1F9tTL5Hg4QaiF1a4GHCgjDFHn1C+YejbA4BEfo6zVj4rJn44uRxVKud+GWX
WPSQ908DmjuPvBp+p6FJ8fFkPWnuKNKggj9kHXpAXnoFjUeA+5Sp9R0y5b2/Jw5L
9zr6mTX53Yrn2JgYiEGFeAo97jecCWBsLP+acVGNMBR+JwlNhnMTQ+wFu8bJ+G03
LB9dK8Qdc1KHaSosQGG9Zf8XLdQbEKMxztS5im9pd/ln1U2ODuuoGGrNNz/8ndMi
fAfmMnhOreNWHyD2JN/tc3COH04VKkdCuVfg42B3RkZfOo1jfGq/DdzfU1mZCrcV
f/W9OhHVkFQUo1tTcKjXU8V4ZmEh5doXhabAQmtCVqFcWNbbP1fCPqxbqmgoNx9/
c5W/xlmaU6yMgn1UzDzIoNmxwYstRfZbNLm9bHuk6wiwByIrtOrkRzSNURVWC3pg
sIILejjklU+vhyWKsdtuu0YQGN7u/kUYj1agVTUHs0Dfwj56hEMtTdpcqLKvnB/x
uCkEPXP9Ayd4YwDVs4bfDiYN08zbtZgiKQ7TEPbOeGSkpKgl6FxUofByuc3GFO4T
iqQWsZMbylFQ5rTOA+ioI6+ir/PJTPSYPb8YD+ES0NxQWj4z4wjVBZNP3WsRIpI2
cXKyvLM71BIbU1W8WEoNNcEXN+ufsCh5lUqYHbPlqCxm7X4y4nHfRaRVtl1YQdT+
E7zwzXkEKoiO6jHVQ/fLw2hxLUEtXdU44FwhxhRDuL53wc2hRG+y8TS8HtrljbcW
3x1OFqi/eG+BRAvEJPIJKVY3vm2oHJTr0pTPchaoy4EWf9prY+UQEcvnlrUX3Fru
DTfL+0hYeIt2Z7nxu2LKVnWrA6TH6YH+Lf/o1UCqNhXjUj4mwS8kb7Z3qy19ALsC
coFL6eK2NEE87aCQf0aLa2IByDSiQ3ke2exsx4SATZ43uZw5pogkjmSDWmxmlC2m
YMWB0FfmmSEh1A5QoC0iITEM19vUUvEJEQ+HNgN5J7nqXBL+qp48cImo3+Ybehtw
ejGPw0qvsGC7PtUvODVCwA39jOz48qpb7ccyHfciDsjA4VxYoCP/GaIadbodvbcb
sVgx0ZNE9dGI2rm3xBo+kRyaFZzHDBhWLO6frQFg/xChDv8/iwg5CcHxAagHC9Zf
iVbKKX+o9jJ/GFGCFeP86GQeTDEBxBr8+H2DxlwA3U4J3QmHG3TLS9U7r0tn0CzV
6ZiYBjzoN+2EJYtuwAvakN7Pf+1HWWPGHRoeKDxm6LWitv0+Y6fr8axPpb6bzVKg
1D2eIht12B1891xLlcUfLsdBBRXJD9tCX+mDcWe0JqBsCizInn3w5RW+OOPrWrxb
81orKHH2OpgGmjA8cFcaqDBnr0oyPcdRGnMHgQYeFXrQO4k05J8PpAXljnIf9ivH
GFO34nff6YvUpeVrPatEK3X8MOhc6DElTfa7ZPpFPFYCNKVxbYilI/uUE7u/kqAM
iC2yBqGSvoLIrqm4/z8Fqd/h0fDGO/dnw4ozcclvFkG7x60wiV+8bJe7/xHW7zwp
jXn6fe6Lkmf2lCpZWp1hSl3199bC4jg4DwE/ZcBc4DxikFp0KhJO4751cUSj+md/
fUk0Eozxx4LogWVnBFOQQnb0G5PC40jz7w9PHIkCOcbMQwJm+DL5r5FM9EIWdW11
ch9pq4+C0C9qaQ7FF6VvrsYZh+JJyu5k8WaoXrqDi9K2zA52xyTj07o9IcoTBeFn
vyC20PzXf+bhBC+kkcgnpHYBvRgWCPi7hjq+jBU+UoGsKxs9Tto5F+0OpxVh7/1b
lUGA0OcSAcJhGRXOYnXUB+c7IfvZshvUulo4kiQg58CqYPE60re23UX39nKDaT5V
9Xa/n5iFNdTb5uV45XYJfjc3evyR31f6ibvJI9VSUcHqWLfElz43HsFB7GWWFvIO
3Eu6LPpddGxKRgSyqFYe7x6VkVgWFf922+UlbnDPdK8B33plIwCY8DBv3D2Ihtes
/F7C0EYNAO90aS3xEd4Qabg/FqpppUjfnck4t5yyuF/4MaDQfUTLED+EuFqsyHKm
B2lcdcujV3CsQF8yF/kNlAXYJ0kJvm4xq9MlYsnWfko7G4m74lIAizcOFy3IymqN
1vlGZj/4MikigjnW5Fx5ntUs10yD0rVZy+72Dkcx7UPSiQa1oxIf35/02FOHqXs0
G9R5fkcqIWO3tj8LbqCpQjr1XOJFd1br8jPIDe+T3V49z0LYzRLe5YbOj2Spft4A
GQnQwz0ewnZV3mI/uTiPpp/xjSlc0Mh5c8zI0nd2Aw8bvxRvhMr4YWZR9sNkHz+Y
Ug31eD1vphsFQ4FIDtYTblYOJXRE4J4gzQxuiT6U8SsO/3suKnNBYjE6nDuDucvw
KB16D/YsIO669BVE50QTo9rRKaW+F3mUBJpMI8q21QtGO8nhnms2TbC3IB9ScR/e
lhvg6bP3X34meK8sDikba2H5t5Kaoz4vnLF100GoI6X3KLKKdMuVe6LjVSM3NrZw
er6+QMKoHUcKnSAlInx84xLmkWLChyx3IJOn5KbLjAoxaYix945RU5exlcjxAtfv
uoA0oY5nvVXngrK/aoUyct+v57Aszb/K/rRoaeCFFJfealEASoOnhYz2dicNhFtW
MOOJt5WM1U6oRo9XPlUHnbXgouwwTMDxZTFIHtLEQ5cpIQ05cNT0qVMVy0YTeVPp
mDcPCNUCxwrhQCSKEu3V6fCqjKzOHy+ooR4OIY8DVTTGF+RzKiglVRHNljcLsR4n
TBA5RFeCwWDhQrEShp6GEzDVX+CfGuhzBka4BMev+LID3UCGHV1ZVWirx2e5FXYm
PsSu8G1E2K8poiYtZht3ZrtxGwPzrHXUcuPQtN7Z2nCkYWkBjioGsKUrSfg2lH5u
E5v/R506qw2Fnw/HWFmw8k4zlkj9uQfLqMP8UUCipyBIQjyr+FxaPtYXJcx/x7rC
W6ZEi/z9/sPIAQiDumxcf6//25AcbOn2VJm+D/dy9R3uUbc3SwclI8UNuY5SohUr
Q/t/c6hD7S8p3tMjEVke+sKY6SzLDep0JXCdz0j6yoEQ0HdqpcJSxPWHsrEDqhPZ
76bP0LAbuMaYIDvOg0FDuQoNcYnHAK7GYwadIAwqzCx0UmxjvffnAwxXnnshh1ur
Xock7OIz/A/bfYXejdZPKNbUfRXNgaz8hlOuy2QvdcoMokxsaVbr1Nz+4j1JLU/9
ABa6sWrgsYPirgmzX/5ABhcbDVRWimbhRDsjmpWY4HSTjnTulT+k1+glhnHxF+Pn
GzAcE/0oAKVkhZOaGfyLoYFzL/7zZ17tsEgGkpS6qNSVYMxrTg9L2SbFUWQ6ap64
i2hMvbwDZgHDHE+Duk5gSVXYTsDf35IRFfUMkngggHmBsX4cnLp9zDDNkwAbBnNU
R9zvpT+CIZLxRYUvLLoiw1qeK8QVfpVPelmpnyB8y+D6WaJGP1L9+baYYuWPuhxu
YeuSHsOgJuBq2pSejR5uequQTL4VL2FTmZ7DGzIOpo34oH1wnj8pTT2a9AmUfUj2
z4HquyPo2RCZbf42Qgc/jWPIiX6QHkIPVo2m52GPeNSWrAD+dtN4PNJhGh/r5EEU
2uFsVey72pCnj8re08wTXsLzm84TDEVunLxgpXnjRtXxYQ44FBUV8HgqqmoNAkEi
5aBZg4eRiirbTJWbYjCQhH4lK1/ucnvsS/IByv9yAYQfP6DDHbuaJqiylRvAsCq9
ivfbVzVYPtZae2cTxONnawGtyUXhAx3nlGntbsvRgOjMFuDfR4aoasYplA7wuoa6
5/Q05+fKBKSqZtlwjF/B/nmNympOJ7EBe55/IlCLi4IuQicjgxhjVANmeJB+rywG
VDAt6GlwoMFvOwJhu4m/MtA2gW9EPGqKZJoiFRAVQrWc54G+xjpHhV9QjYLFlKTl
d6u8VMo9ytNnvpBxwNLywWE16jk41iChHgLqIJ4nK+HK6rzO2UtgFq7nYRRL1nb+
5QjT+KY/WVdRXyoGwJv49yC5bU77Iqkz/CCy84qLi7XjI4jHixUGsd8yzkV6duOY
EDPAAvnrHqt6yiSvD9MK7AUeRAvX6MVyJOl4mFkYFW3vCNn5HvxwKQaTrehHvDGS
P6170kF78n0J74Yf/qUXDO8wralEQiHCCNmSgIKMSYf+xHAN28nLQBtrDIzaHcG8
qj7mrDs8wIbcbOEPn/YG1KNQBkalhgZ9Pu+26jtTIHnmHLmZrQGmt6T3Ufg5A2wU
iFSxs7kqBIElmUBxfnHdv/EykZRQpLDkFQ0GmjQiZ2Bp9Edde2UkO27JERaoK0/I
Tvw55/4rurPO4GvJtxim45HIeHLn4b1oRu0bCsKIhnIu7+zCnNDqDnboGI3I84Bm
33Slu9AiGhIpbhO06fnfw89KnCsk0BCn7W5At9I7sJN9nYHAno0gZgsPyqq3xNgO
14Ez1pylsMpK/hauhV/F1tLWn9LjL6JmioJPDsoZLealLrqW2/JqaDnWsJySFV/a
/+mCVA+xf75GYnSKfnae3XOc/RvDLQHp6wV0izCe7kZ6UfQJhkzsqqKh1DWpjpGN
VQniYT3ZTvyM0zOCSgxfpkckUPlE+0r+fxw9ae4o9mOkasQCNfQtPK8PfWSfckKp
flEfye/Zh1Mf2lz+6c4UjKokDkuvhZq6eRaWVFI/GhXOhKdk6PzhMqqrPgbEXBni
cD4WXzdABNL5kfnFiLd5oemrTmqd5K7s/CGfRDlMReHua69U7s0182BiVXCj81SH
RUfowDzK5K5ebai7UMZkylw4c1PW8Zv+6XiWI2FPWUS7ynjDW3OvouYRIcZ0ySbt
G0Jpr9G0IAB3kviwFQVR8vPHCVPcLSwDwXHsFvz4CjXAdfBboetq8XpF8fbwCqmY
ynchLIP/jP5cQ6vs9WoLXGqC7Kh0LxQ0HPVG8wiVFcIT3Z1kv/g72NAstKJp1B7f
9uilVV5wPhfLkrljhOsdGqc+V2Tu2AtH7SwBVu7N0/XHrK5VvW7RkbfKpUL4aRhM
cnluRYbZpwT8BBcOTOZkhAa2FrqRs64ErCRPPNsndlTlyFwFMepEy3C7ninNsHRe
uqsd0ty4rbUx2DLJA4YYopKvOs6SLJ+RhisKQWfUb1/KgEtxHM+4YLEdjdLNHK3V
DpgbsimwgqfqJaRHIn5s60pfngVERJ49Ozxfwgad82vOGbuyMtJwK0mjMZc1r2Mv
lfSYcYHstizRDkS7+VzwwaD9m5xojt2AUFvMntfhqRpfX7Vr9XOjm6huIaNBdpa9
qw4x3S5zHpIlXXHQfpRtwQA44ikKs7zthO2gnO1WZgVfqVHDQuQ8qvdWiWB1ZCt2
mb39tqrDjORxOBhI4+8mtJ4eVx/cspQWQht9vTpIY3UM36zQkYAXL6wIkD+TDGl0
DrnltT27sALtvwiY9d9FW1ibh5ftf6m4sf6zbDHyB+4KZfZqft353Zr98Rwy++Ov
L9Sfppf5BkI291pTTx1oIS5uW/h+saIZanTAc2LInaKnCi2EWn2G2sX9QBe3td0X
XqvkFEtQVvO4qhW4up0wSv3aIYGLMDWqsK0HMFaCz4/hTVrMcjzKP7isd2cwU46V
x2gwueTFqxujRqCySSFE5rQhgcE/HbAuibu+j5EmFZQrwpvs5B2ZJZi7XmsbR0fK
bLGQjfzSKM09ibkqRyK8Vbi06mc2S2tOhLJ1SA07PBoFOKes/LgbdBP6FjWHlwjk
o+eWWicxbPWId1rX1UK6mbhn1sIxMRRwq7zXnRS72sfQbFojOWT2UOfuat5HIhRF
p2jgDzoJXOv6P2ZmjXmB0XIZ7biV5SoSNL2PFV/TisJYdIuC/MVLAOEvrRSIakUi
syLp4nihzm1BnMcaOmObuoV/C4WLu53ZM2Qo9lG2dKqJvRs1tvtM6FyuoJVQDLOw
ft6UOH+AMExuxFsrk5dZ5hIJCcFeK+iMUcRuEd6KwZBwhmSMv4YnkKmAhPThfXHD
jUgqKAwj6pmOrbFamxd79bR3wry/GTo4HSkKi9X3CzC0kbc9zOTW/dmTmwos+BoT
9HqKIHozoYehLbsYBRHEGOwsQHGsWAqw5DXEalV+OuLIMRPYrvMdqnpPDnoL9021
Kk4IKUT8QyDfO3IvZukn9QyuCW/M5eWDWhKl/CNqq+g6JtZ/FsS1oi9Uyu/00bCZ
1X7wt7RA5N+i+YIFUrrftz5Xe6a+cO7/50IF5atIvmXfIX7QBNPQFeDipqvb5yvh
njZz1GQOHNS+w+MN9cqh73cWu67gNY5b1qCCl8OsIvbfW+MguyyiUx2XKVfWus3m
BkA8hpfkM+3xHSUMdmXqqFwm+vbfWK549EpF07nzXVkpecfj1iLLWT6f/kfoVDsG
5Omxx21/v/d4Yw90P+M/1hrrkUcHGqJOvNOmRMhCVYdy6B+82vyrmD46nJU1p5/d
/YFk+EsVtgj6IdyX5/J/94OSin3ZhBdsV8zlBoDGg8/PtGmxPmnCXSwU1vrYIqeK
7Pg2L1yitZhZZcj2glQwq+fSOA462c9/daHpRI87jgoB2zLclM+sYcy32gB7MRCX
Lhn58ruGsC6eQziNtSGck+/EhmBVllhS+HQckG/LieGEdOcPN2jLzSAkFO5ahnWP
CKEJRAG+0HjB5GgLjQGVm24pp8sPXB5my8W3V9AOdDlYAdAqpRNmzqM56d2vXXcg
0a7iA1EXrVJBuO5TFgwFqHZ3eQIBVxZ5es8wB6NcCYPKOTzMfBhQtoHtzY/qhamt
DGzEVT9TEm1JBEiA/qAi4kKk5dHH5rbZFoqU65FfSBygmvUBj2dEOF63xDDyV7nB
R+9PHqLfONTeruAnZtlO673I4iivVsseHuPWftqL3QpQvy3Rsp2us0YMIshwToAO
WessirJ78se+fQlnXjqDUmeBU8gaVZ13qX/WLxv2eyR+0QBn7efSLqCrEbQle+fM
Cb62sK2e85urX77+BEigA5RuOw/kyJttFlEXyRLPIWME7hlYjVyE4VsK13waoka6
MloJU9Kt1zDE4c9zUdDFF8mucUZ5Le0byWnZMB+Nxa6J0fG9MC91wri/8A61COHy
IjI4VTLxJ8CK2OujF6AjOoGvsokn57mnMvsoQfQCSFCRYtflbohCIj85Vt4s1GSw
Dcd1JGc77IjZphVE0A4eLlupUgqNvCKiZUn3rY5Jd5G+G3nq3rrluDcBj3/Z07bS
PhfRZFQr7eo+rU0xHTRXd/t+Voye/UJTxXozll9lwJ23vpnFpBpfmiPYpkmar9sH
IBlQgygSifmkMjQKxODnEKMxOQytw6cbuu5fpKITdjo92aew1TlkXt7dN+oPmfkj
FpcsjerIf9XP9o4d/B8GyNsMosQ4jwKIoVSqRSS+dMJ99dO91hdZJpUVpl6DpRys
XY0KTlYu5HHHtlinEmk2B8eAZt+/FbQKHz6BesF4gJvGDyqEkA0v9hlDMqIbHDuN
gFULk70HEwf/PA/lMXWxj8gkHb4rfky28BzotmNX8pG/QVMWGxhChNiGEFFC11O5
VRvgeu22xOXFMMGomyij0cJzSklg/kUZCk31pv60k5eCL1PHSgmve6mHOIQZCrB2
9TttaqnHNZt4XGNuEd0nmT3OuWvV2V5Fmglr2YeFquBYhmEchAyAs7wGSAlE4Voh
gCW74bXNjNn1UG+6HectOo88MYHc8Qf0On7XMWqt4aft90sJapTrfo7u0e5baA1Y
BbNW+3MgtDcPDhmZ4at3dAXywM2C6p08DLX9ATmjJaydtvfXbTIATr8ltuCh+hC/
y5f6lr5PAmGvImmbCyHvJmovOo0H3UlJFImHYsCIs0a0LfDvNATmdlLaA6NKtgLV
depKjMveu2e0vdIGp65067Vg2vip7AKQ1aVqzKdIxZ3acabC7CJ89oQjilKokD/I
dYSGC+s1kBeb0dl4KWMziOImWbix39TJHv83wA+i/248kFDyxTZkKE46QedigXcv
bFN+yzGKh+RfHE/eOH3YunCJGTrD5c88fxT1x70MI1IdVJM2neYS3VyvUiAAmTob
1imyV7QocyTF4IqEba0V2ru5Q2OJKm8tsKH3n10WGR7k/Bx7QFgMLSQLq+gHvQR1
CyYsZKAsgpFWNARuFbdojq5e5n+388QJ3rHPUled6YHR9xI1iTcutP9f9x3JyVaP
hBjYXduwAG8O+ps/7CvvWsKedDl9UkQlryQEOedcth0MJc5MQ4CtQe7CRl+Zg+Zs
FB9TZtu1mzj3HJ4xLtZshuSHiYppeOLKv1Kc6EunuS9JFsNZBPJ7r0FlTmmXs7Ba
zYFmo+rH1HRmoY6wSQdYZvsGusSH/b4Z1uwlT/dPrOgwExRVNIcunJ+fyqnKs2Et
8jRKtz57ct6Ll5bIGHqKvjVjYH7vPCPt1YiVJBf1rN6x9gFmNKkxgM19+7evr6wx
Pz86OiQFFMxNdN3HQjZAvtmHBOViddOBf6IhYirT1fAzhdaT9Vsoz3OFGNlmfKtO
6YnQ6RbF45AlYoxjIyBIUWWSvJfZM6mJPOQxfRlVOTDCWyQzdYqHiSx2zZqTRzTF
Q7ujgIDwycyPmWTv6kVj0ypkA2LrrEuMNMnNqjt/8OFOzebTtxpmxjjSclB+gT8o
OB+VBnEWps/GLWosV2NtK6sLCry5Wr7f6Et8zbYO+Gp5ppf8SWUjnRDlt3cqGfVV
v6NBjANGU9UWa6IlZLlr8NOm5o46IQ4ksr0tTvM619b7nrVNLJVPhNnrrf2qVXpn
F67WU6R//0aPh/MccQPqt3KN50klemzzAXaVBXTpE6lHW+Q3+3SMcSOQygjk9Vqx
PtWQEQildOpdY0uiDn+rNiV5Zdw0jZLTJhZGSi1w6DX8/zQThDe2WE7+N4lDIvYT
edO0GldJp/Knxn1MqTLy9uzcrKdVQbKwestApI8084osrT4Pd9cnDdbOTiugnOFG
j78RsjV5SORNdZ1sKMh37Mfns6wf34Hd9XZYGt8mW/Z3RbUZvDwdC0kjMXVixjnz
L53pWW4YmWIC3rAInnM3Y19D7Kb8mtNl+wl84CLe5M+LKbxPEVDF0nnjg/pOWjoL
86CWuj8tS2wl7Nfk+tQPGTqATJKGh8u6VQ5kO//L/iVzrXd/iUrEEDzyIuer0iwb
uZs6WR67G/1i4kCZFNeE1w+4agcGjGJuLDPMRiSloaSpNLPkfUSCSo1aLPGmruhi
2AJzMnGcCZ+g8YsZU6tw8VaJ1Cs+JJZI/xzksicXN0dPrDmwUgxPwJgj5d0EFr8v
o+25vyDuamhp4+4h0NXhwumGsNjkfrTY10W1jQqNP3Y5qO9OzmFGWLJGQd/xNgqf
FwUYl0LPvdnaPeQiuFZgxRvWdbBu+3cC7guL99YPTlKaKJHt90HI7YpisShhWFEZ
HYJDjtvCjCN3G91A1zx667IuJAqZu8zZrdXY7eh966H/HKNgraAfqqPvtGVT/ZOV
bCYTOc9S2fzUNhF/XsZUISoS3yC9Jl8ukFDrFsieEi1vedueojjKlQ+zz00GHqTW
wUHD0TPHhUy5Hjw+Y9miKrNBm4GecKRIZPrd6YsxxetKH77DsPL+sx9psLGke/lG
Zoh/yiJCtYp3W4qgxmVio2tqjSmLEZwrFuNWXYeN8BsW0LIkC1g7v3kEC1aS/Y7K
/Oruhouyz1EdDFvUbaJBpONSjlsQYm7HBOi61ZhdQ00nt18oDD9Htdh9J9PCzcnF
Xp0RMt6WH9vXdZN0Yhxt+Ms3bbZR0TZ6GIdW4X+Py5BlDdBYa0+wm3zxfyNa1PjJ
b5t3pU55EMdOWL2yOJOSaCk8n8JMLsmNDmnk40N9sVMMdSQTc/5ZuRYp8nVgwGY8
Am+x1SepVha++VqXDhHv7sYwnfQkXnBlH1DyNIC/Y7CS6eMmPap1wYQ2z4IqwQ55
Ji9LH64Tz8oFMB2h8Z50bXgfx5JpqFYLtnPmg00Ptls=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
KiHkvGjmUkKMLhxI2QYJD/m9VTGLAzyhwDxsuFvJags0zpmH3/hKg08dY76tJ3Re
eEoyE+Mw42IkrKaMoFW2V6RQFjFTKW5QTreZBY6pqiCBE1si1btkjhVonD90X0F1
BVsesWwaOWMXC3XyvCp4oY2Pw8Hgyl/79knJXs8+g4yOQKCgMC+YOOZJOQ0sWQ9O
Lwbk2G6gmymCjx/dtxtOKmVbzT4HK0+Im+MlOwFV6wEelhT86srGhw05mWFCrZXw
YT2c6S2tQRLpWmAZgrHUV7aYE2ewhlJApNvmX9mPiy2jOte6k4Rb2N3vavDKvyXT
hO+cJ5/hATGKvoRVyMjXlg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7632 )
`pragma protect data_block
o633S6+MPDmPxlW6NvlNonUi0Pq8Gz5JqLWOBPUZn5bGyUPI3IUMMNpm+gkv5kYr
OEL8QCNQxeqx8VGAH7k5B5mYT2yBIptEfdfIUMbAGRyGqWya/h+Xxx2jXZ3Rz92h
X+oaIFmR7ELTk3f4794FxIsQugRvNPQmM//kuYEcnkVF0zizg7FDMu0DZ27ca8kZ
ZDlRoB7xNB2IFpf+hwQY99BXf8Umv/VCh/ndkuKgjSGMYwHc/5zuZ4AQMxfHYYpd
Z2brIn9J0kGs5lmG3YTfazDuaGmlDCZNOVyfCBI4t7s0ts+KGihN1tlc7CmchkvH
aLZbEfLzn+pKzbvmwMtG7e03yo1ucCHbHVWXTGeWUywbrUa4q35TmvQ0M9Dyo3ms
xHMWjQvKb79GhJB4OE+rlYHTWYXLCI3yzc3jRSjQZvYuqnwXa7B90wFXjIr6opaD
gfVvKmbvW5RfnW/kwirIwJ4f1eTrLijYaQW2L1LiqP3qZgJjLz7P4AlnyPYVizro
xxmZPsJBLuXpY+zIbS+4PTtnVPHbeZqfl2ZcaQv00yz7U5WZ5Oolu80Bl23HXUxm
IWXBkyL+YNhl/bVYNsXY4XjCKHGeognMmz4HphbULY6PkmuJXQrIk/J0bOrZaJJN
lz5mYxnv5Ai/Uf8Y/xFJfU53umo+alEDbZkcJwymN+mE88YFbPT9do/anv8xNepu
3pxdZROcVd1mNpwW0xdFVT1k9Avzzsk0KWqpiZwYr/IO9UMRygeEkFLB0T74SjmR
IyqDLRXcJmP65kAUuSRt2ir6GoIkOPiCNTcp8MLdY3LGKicy5m+pHVOvwXywGmsQ
a3x+M0S0GEfIv8P4x0HtFd13almNsBg4xSncShHh1m37b3QRFDTMnZZD7pKm/+PA
Dlp1Gn5JBfUevYhI+dIt0DwN+Fs6HKUUbg3FyjyQIHPAODCTpPdunzq3eoy7x9aU
IVm5ortOFWxepQjuzIgH1e0nxNGPjl2wwOeVGokNk2Xgdd5N5TGVscslYVrBWtEJ
2cqW905QJ2/h+XILOkx7ZqXkBPsYXHQz0+6JWxexMiXLLaF7UABJ6Q+KSBrRPvRM
EzEfgR6YTWREny98UoJEmik28ZLxpoqs7hb/aS2QfZlDLWF4tiyJN+YfAAVjxL+f
L7oR5AsxTW//OBeuOnOb3JXUIPrviLFMfEi0hIKSKM6SJumIf2TBYx6qjhjLy+PG
ONsXlO5qAOVvtdPm2d5cpbww6BNGuH0aN2xxl9sCq6NjowBbAw0aXjZbhn6rwEFy
K4RM1GCwhWdosixz9LH+QHc70w5tFquPYFqd3vrf/S5BPFUBsbiZBZwd1Il5DbK2
89rKiKem2STg7XopflkZ5brHMMrkJC82wFkkp5Njwu+jm5H0jAHUIUAhEld3lqbM
JgFQJDJ5l1okZBltm+K7P/o1NMKwx5t9qXlSTPusecPCXlMcQP4tq1TqyGZSCk3H
aWGaCGfDt3CTGor+2pKpFg60UB8MO7+r75aSSNYV6qL67Zg0W8irvSGtDELl4E4H
HUXoLjW0SUM7CQRI9uzGUxQxm4UeclE9Ua2+wOVqB5jF0/FBa1YJDnEYTGtO2Mdi
p6zR6QT4kDkBJoL4G30XjnP4QR5IO4NxAYG4rkecBSb+Vf+0lDekmnzmI2SfGoAS
KyXnGyZml3eJ5yldYDGlxgWc1XKDmkjk8lfCnxjSpUKsKLtw2gdUR/IuoEfAd9pK
LFZy3aXJpWzy/1cAO6INDovMhYMSrPycDcWR8XFkhRoG8cOhmby2v8imkT1fYg2Y
GLbfaxsQz69TPTsULpMWKWvz5j39ksV/4DJlFKgk2BHPTWH2iEVP1NDbvB6khtkm
L0XCS+X360WjyKQhmRAQ3NIZ8DTsrd3yqIrua/XaGvw+TsCCK33BLxYQHMMIFLgY
5cs4stuaaHVWA1NJaPnxsTUwLDxJdGk488x+PHSBL6BnMytNo04NKcJehstb+IdW
y2oX5rr5ARTWcsqX/zPMqvU0FfYz/eAWpFtpRMxapwOILiwnBtYw30lr2ksncM0U
1Hx17riQI9yOdaLfErMh3pWIzoZScJnuXUnsWXFE06B7+09WnCO4slHS8RmLHBbv
sgDz14Se72zwaFH0nRqmx527pi0UekeVkGZjd2tuTNQae6FL95lY2Fi0wi5eKw81
MEYgNiH178h6nWB/l1bzAR5jnDAQpevGLDOzTZ1twxA9iL5xguXMWWekrhdo9htR
roDYQE8FY9vFDIR9Czf50odMnqinO+yLtZszfvZTDr27KvIc+UeAmwUKiEhCMGI2
sFcU3TTjr0BOAQyT7GeIDnlubblinU9otCpYghLjbOILN2jtdCxXwjg5MOtoSXxS
uBvxUlV8MYwE3RaOnx602Y2JP5Zd826ORXgzGwUzl9YguOOUNsASbW59vBAghp0l
QP0rwRzprf3KzmYFTqIqedJXtKbWfK9ptwgVfeRFzAueX3r5r3pbo0topDTSuvWa
FY1nVPjGrQRgK75hO4ITfVqDipBXUh4E8jOTIkdX5MRUGa+b7Gze39dwsGnu8Yj/
l5dHRiUZ6xNQj0Ia0q2B8YCK275xum/aTz1/o3St7+i3PcnIFO04wYLmP13LaRGu
1w+AU/IAVjc8DydyQ726FI1PUYlLQaq/h4bLHxiykIYUyZRnt7aG7pt7IjXKDQbI
G4RkEPPFfiVhStshOW9hgmKizsyYxXV9TLLYHNk1v9+trr/hG1rV9CZ+lylA+FY8
Goai0CISrIGcr9hx4jZjBbzZEDSZZ+c0opaVWm7w0b7IRQcHBmyWyo8tI+7zW5lJ
7X59K9SV2lDaljfVUVa+Sk+c/aEVMiMQ27eSXodSGxtoGWW7ml4mA2x6S9qynELj
OqMLPDdcSqVPiYqoNRZzndkOZKGhP93RlCtD/dsrbjzmEV2qudFQeVNLEsi1u68E
BRVpHvQkksdefRGZ8sDHMeWaBzi95VpmAcYgfB6H7wB0Chr8kwbOabmjoLR4IM19
alLm+mtr0iMfT+i7BQfd7KJgDSsEbU5JOUwTr28u72ccvqroJP9DNffeTW4cG00m
cWcDrTXCTq1XXhz6raf6PbNKczJptH5jjmFnmzl6ryj5Y9nxp+IyP+uK4Cmah8i3
3V0e7TOifjSm5Ag+PqI3TUWsDpeVzTWfT6+87kDz51HCgE44xY60EQZervARoknb
rXu2d4qvvNqFFtuu3b3nENYoTii2DE4eKg31v1DdnKYQWriXSq2AUvoBeZ5RBlwK
ZG9CawessYJHezQFCjRCgeIYTRZf5nWuAoJlqsiEoSGEYXSI9ANAsMv6u5+d1rGp
zjsw8gINPsUp3gTTku70FsjUiwg4GEnEy05c6g37EDCV5E/VT57b6byk08ruWfAa
hAy+Ot8MH4KuaVDbCBiJhOxnmiItX1GkdBpvHQ5srAO/sF9Ekz7HuPYUiis5JfuZ
D5wxf1gIuOe9x9AvLDQ2nqGvqo/YrjN7PbMsIJqlVRa25W+b0/u1KJgGWrlpYfeL
RUtuYC11hLCxsGseQ5ZM1j7DPtjh+qOiF8+cVTIRLW6SJNxQv5yaHQaU/Lk9GVJe
wHNikoVMuIHsXqDUf/xjiGGTL+FDB+kZea+nPCSl+s7hGZS491LNJo3ZOwEBcyaS
DgQkTiW6ObFtJzZbd3wRhfEtJWsbHKYJ8Dys41SPw4Q/lSkq38fNufJjV3gkk2zX
LJvEK40O9WD/mzwSUXA9wcOfOAF0/dH1cZhRGRSOCtvCLhtma/nAc3Hm4rHFp8Ng
m3WoLzMuHY1zvmZXUO/w2a6yqqx8U/pt5Pxomi+3fN+RqxzDaBbAWjeFjDYT5BoK
qUFbG2FbB2vlNTbLEsXhjptzOu0cN2YOoZkRstgp4DEgn04Vv7xqSKy19uf1Fs9w
/dBTa/owawNTrVjtb/1AaHny/A7FQ8MNpWV+bGDNBPKfzWtfgJsvDraxnZ2gG1Bs
QGZuxy7SMj2G/cEVUoTRHzeok3uclzKdnMlcb+sz+c9tWxInoos7HaSMwb9e9tCY
SkcajNcg4C+NJiztjLNl/x6Weud2zquwgN7Wi6xiWf7D8lXygNtCQw9kJX3H8obd
U511fn9TIgfWp1z8gpeMgvxp7lPYFjspfglfVIH34JE7PSrpEBYfhQC7EZhgOzCG
zDOjRLU3KEGd9piUkjfk9Yygwvotf21c9LKDwDSPMRKc0lf8EogR+jjGlLHjWSWL
Qb3YHocDukzPRuDY93wMAKkmiNEpAHTfVcb6uH2ddwaorF0THw+x+PZ6laiWJ/jB
oF1/0wLFoqE7L+Hs2F2iRp7KBwQyW8j97scnqIM6E/DcS0/XX/mheSIR/utXfiRi
/sxgQA60iKSvfWb9dEI2TcEyoy5SKNjllVXjyrYDPkJN8lz4ixU1In7E8QM4AFlP
WK3rW7KWBa7VahjJyD9tyxdILQlZEj3K6z+qSweeRd9xqy+qYeW+OGQkqWXxa2p5
+3USF4CNiOp58w7qQHdVRLVuh9ndjh02EFgZHor7rjqnU/ZP1YeQTr27M8ubxhn+
OPsAVdk1sBgulNzTBMG5jg/4eXaf7Ws8T4AckLCx7lipGd8Gckf9ptVApWa4YEKW
0vDCn+IECZ4rRc/IWfA/TOXcKRa9N9S4cKJU88HTa5lgvGgpwYCmr7hQZw6M9Al5
vTNyC3zNl9w27gUXRkHwc6zCka9hzRfHJWv+U+TQGJd1fHrXaRS7ZzLIl7mn7dOW
vUOWIDSJHuSC3Exm5/etB4d2+DfT2uNGzm219Tgj/y4GasuYAltTS4SdJg3vGwB4
6LCIwHSjX115sw92VWREVoNWd4VI5AeKVB2f3rxidfIdSRnPAlFYO90Z1gCkVlbG
rQyt2Z4oBL+RNDIMBM9mwjTgl8GhQ9RWs2nDQ6s3cS6J5UOsFqICCH67weOmt43j
kFC8KKtA3ugS1kH3kDoupZeHBF6FXAC/NWGwKBFprri45WAJ2tTahNYot4O9xe74
aNQKQUBpFGQsjVujzLDQtgd8LpHmsB/m4EvTqKuqBoem2sKBgCJxfq82UBUiLxXT
09mCnzF+CZNYKohSKhfke1T6uhGQxovN+KrTq4JcCqZVZ4oV0B7s83RGe6ANAx5K
BhfE4eewIQQWBBlFQm7WL6nRysdpgUx+5jvz/mqyZLfBjDB5bwk5/X9ea5S8q3hV
Pd8LfvldcE7boIIVFlqeiyrt1+BKyHlpV9iuRllAqw/nUm5rOUR7RcuXw3qndBQu
MfEFlrz/HMIm7MQBnGpa1tkegCU18mpUpyJO5yPqWUVqS0MJZpnn917cdXZN/Vb8
bk0ddwraomp99nuEVOcaRNTAd1aGQE1Vu3vAlArI2QXXm6ghr4xBlQAf5Vs4s74l
0XpGtOZ71r1jNRYp0unm9tTd6knkjzFr47mVL0ATTm7X0mxUaSSbHRerLO4XXBgO
TIJfg05fjwIFx2EqRmgDeyQFfs47CajhrTIQtJ6eBUpLRWSqV4rcQae6KECmj8na
E8GH/LwcQ78/i/qVOUdxRztgm0ACucTZ1LfnWaRUeijIupS+m7yWkmE1N9j1lLPb
K1ops/Fi0cboct2AB6sdgCkpxGRqvdrnHahx7Q/2rcgskr4aghO1fDexVC45B6L8
TZkh2LuATg66R80EhdywudDvGIBpj4gecc562+NQ07mqJ06MsOXreU8eCm9VCjSf
kHaqduhMfLvzeIfxq1wKoDDjntIyYbseMdPL4SZZq+rieljysZX++FLIk18QBg4H
wIONdnf5OfpHpegNqfZj+Y8JKnlAYkNJoMY+ghydDXHF6i7sUemwU/iAVsVueADg
vdhAfQMHbjfgM+Gcgyo3IbpmXg29iZojUtad6L46Z7Yk/+ZcPuEkwoE3bB3q92UX
zojgfkLrAI4J5MA6cYbRAjFTblVjbkGPZxnCgTU2jBKj//Vd6wCx2Ikg7WLTZTQL
8zqIOqpXCj8JMY7u/WI0aPsJfXbhQ1sAy2bVlYNYPdkKM7lXqxMv+hMr/TJ1z9ZA
6p6ZPbRE8ATffmrKwI7xCyx45LV6xK2TH288ibLxRPkOKL7xXu6sSSFOPT5FaztY
CoQspeJ6qpjAxOZAxAZ2Nv4478jy0eeL6aJwhHPVv3OuVUGbqI4i1L8Dpg89UXZa
9QDcE6PXX4cSDrrzMJ1tSvp0ErGlQ3m8snA34Xceawl6Y2pmBgr0GmksMHMGQ5p7
pQjACMc9ifVfJ8/yNZBGsZT5apGVmRRfY3t8F4Cwq6372yBBClxCoh2YZ5SMIy24
5PKB7P90oTuXiN6K1ncXfl622uBApIzS45k8oSJ7GadGt1OuOQ6uvyS6v8KGicda
llKwIS4IGIh+3RfGpDyPyI+6lVeUUH01AL9Jq5GO2n1lWXFLBExxlbJDICYxmC+U
MYc7k9TJkb4IdvPUUnEodIAFYEajOcnc0oYs6Sr1UmKf5EoEA07yYlvCd9MrezGJ
mlsIYOYUrAzio/ZCRTaCzy16bBri0FY/HQHxfdTcEHgpS0jHXAWjhkwJP72oPw9e
SI6T5/FTqSccaRDo8O7O6WOXoA6RasMPi5CsJMJzhNQXlK7V8NSli2RV0v8k9s21
aGEcRZZo3BlvRN4UvmlUtVmwbSaAEUHSlD0LGNL5e/u1vlvXwNNeWUk5Fiv7VVk7
nFOKjZbuuBQtO0R96Ffuk9xcfDqX9QN27NxjYE0w1K8MdQMGNwQkOoeAh8aPqdHT
XmnencaDQ0qEcngpupmR10rPDpsXh0EboRnxLy9FnC/1qwVavCjdcs3BykS68KaV
JoDNZoEmUvn91k06Kog1lX4raRWdJ9KGOjOo9aZWcEnbe42ViCkZmn5HHIT47f7P
hb2sudd1Ec4I9p8ebjDNkZdw3Rd45dg/99XFZ+FVQAiQb+qDN8GkPReM2178ADjf
OFgyRwFBqjAL+f+5EnnRK0zLDerwQ8ZWgJyzYsq9lcSj2EJ2CkSuNuy+GIR4cYtu
OKzHWF3g/tFwfFg3VAPMVn4kOkme5EBsrlRggfa0+dDMCx2FfNiyN7GkgF+/u3Ns
IklojLWGlufOVe35jcF0C+OMRwuOgiIciEO2msuGabzCt8cVDoQnehngoay2pjoC
OZFP2PdjWWNW4ONvLWjMQwNtCcvSP3+kVbYLlSfuTbD1+iqe1e4hxK6YSwyYL4ve
Rw4JMr3SgADwHXs3yAi0BRsXdeZeyLTE4/jw5XOWVkuCJX5fj5kNKZZBb6Y0C7gr
ZATuxqNQG9wFE2jBblsZ0P6UBCWwfwBFTKjM2J3x81k5HbZdvQwVvuwXvGJOu4EG
9G8XMyLlXBGNO7myH+Y1SGKCsJ4zy2jtu+V27Vt95AwWwPVfYsVRGnP8mWshY2ow
CIo1XIZeEzwcfzhn4XLHkodr0KhoT4FuyTrmAjy6c2o88qmYxsK6yBeekyqYAXLh
469XtjmgjKD10NwNjmlDeOtjE1fHgDkOOBp+hKt9amcZzmjDnich5dKly27h0RzY
DCyVmoj/nze4Dbu2gDtLxmLMged1Yc2OW1nCCGjfDJePpcA532zK7TPtD5JweRT7
QLSp74B/fyHFXKAcL/B1beh70ZlXbSq8kqbbpxWl+4WKF+h0jBMhdLZX6FcuMdy+
nzhhguxhz7QEoPsdnpy3VQesk+3+cHN7mZjCcqbtV+oSWSx3/zfm/ye1xdIwIuOZ
gm6Q+GA8rPWvBxRrC119fXF98rCLyMd86OWcoSkpLEiF7Y9zMXtdN9Q7wsHFFeQy
YHSD/i1FzRkobVqYJr08GipHWx5ePLl7ANvbKv+iOcAFH7v6nDupbEsbvLB6k1t4
+XLC8GGOmN1oG1/sVIGBJ3xc/p/A3mkUKEygUfbZYMZnIQirn5WXMz3XfR9l4hQa
Vro6vdw3wIvuPzIiOc4NFrz0Pr+/Ie9QDWcx+dVCMEY4saXZAcW8jRpHQDeYWDJn
GI5R5zHIxUbauWUI/xDnJz0FXy02fPQQ4n0uhIbDPLg/w8c19N013KTOIhXRUO7T
HQaYkPNk+eM1pVFk3/vF7CL+Tm2TtoiMg+1SL5vm3dDA6R3cUeatrlWeMHYUnjNI
TW8ViOFbwt29Non58HpThIuP8VyUPojNuaZdYypYaA/yTavPYHclGY2/kWLGHy78
qFWHkRdXVho1fYjwihjEDy9BLf8B2o5rN8f8rgbcZ40EBHSM+HZm4NKl66Y9vmKU
2vl4OEyZjBqSB7pUI5qXgVuBShpPIa+fDK4/V+RMnrEbpm8Jo67s0RKYiXmZvonh
2G/apanQM8IY4o9S4dcK+HNg8TN0pBUJxiJBzT+xNACKv8mFvQLVanuaVB0xgZ9c
S70mlgptuICFvHZ3Tja3Mgi3k7/B7QWa0CNNPymnwFfaFG5RjA9EZKn8Xa6uB00Z
u5IKuBloheCy+A55T8BNTvmy6BOexRdleI2hYWHM1BpeWdbnzv5w47tWK/C0gyVt
cJiw+yFciF1AQgnmm9uOT4ls/SEMhPiF8SVPWiv59UWEF+bxXcdOhhn0LCSBdUS3
3Cxw7FipboWBqyO2sPbQhWzHK3MVOO2VpKBsFPtEeccobDPy34zgarhuiAhRlFwE
BXHHmObyk/leFSb0QenfPznx2hecd/xtJmCAzanZ2UbFw0d8qa3AyybRjjFseGDV
WXbW/5hoVrElPqTcfnwvVIDiy0AH8WZaoAjTJHYbhzFkUw1qH8zxGU6tFO+b8oqN
F+g8nznyYtT9ArrrY+GQrt8uHtqIqciwTF5TkS34e1f4QU9ysoTwonypcnIbfedM
uue+hGFuEQ+VZtEJQwi/MJPJHWmt+V391MFUzPaWdy8ytDqWl28S/uM8gF9WXwie
dt8Cv5fzgb79H6bz2YeL+I0Xn/6WH3sOdhuAtWMmN9tV1Hrkuc6Y59GFH0vTApXM
viE6uHvGT22PSfOffie8AcN/FkMlBrQyk2b3yx3AR0kSTYRpk/EgZX4prMr1EDFl
KxYOdujWoOFxBhmex8nQbxgSOYPQCu+dveSDMRfRBa22Oclc712dPQsMmq//635f
MzqUMCxa5p2PJpwrqT/SBvoM2OrHQ7WO5veIiMPPp9jjb3v80nKyzxFgR2LSaBq0
N5X7p0iZWEMufGrUfucWfbJ5iI/a0mVQs274KZ0HBbMmqlBgWQO91jzlamAYATQp
QNxUqcoa0xqhH1XD57ssZ7Y27bonmkZwMXh8RbzI7BvXXffgmfDAeEw1WZLJdq4D
C8XyHGyTKlh74IYl6ssHCMDmMqCMTiRjF9Ama0I3aJ3qePbW8lS6OJUJXQWfEFkT
kXddG82TW3uUjdKl6r4c8eSfngn+caLg4/cGzMfEtII9QIIhCBfToL66r/CQnIhV
pSz5P64jICoQ0TwzFPzbThJeSyE5tFqTUMAjHQqKyel1zHDzuctTbRPUhCYZQIj9
F4ZQtaPub3HwW/3DzbyT5diDvx3qJVjck53au+I4ICgSwcQaLC1lMBdSE/vkI4j5
ZzFRhURzEkC869SoyNLVRHAhiWMUPzasgF8MKAHAYHuvRI9vUWu9OPfnEWE6Heoa
424X4J+H54kCPJwSLWMKM8BPYxzWQ7mlEVMPqwSZQ0m+pxU0Ek/7thSGtSp8SNFe
lPRwuz8Kg+idqLYaQYL0C61kRX4jJ3OItF3x24q5ARDgm2YEsMnXGnNxOPcPYzMk
aVLH2VGA0wF9ikN03g2MsDD/VmSUIVB9ttmGK0dUojZtwrZZ8JNgNkuI/v3B4n+I
hhW0Z6cI2lfOFowK2aS3GcTMcGt4gMOWR8I2iXzF2Ld0w3Rf4gBFkwrFYzgUpPQN
ovpS8euz+qikgOgTBY5iMrzRxvx4e0qgUcqKl6tABXikRkz610X7m2jD5MrW6NcS
zSH59m5x5V8rP+ZI13g7/ha/i26b0kux/qIRKFwgob9cO60kTyNXzp+MaRjFVXop
+Gvk96nYREDGWui5en2dXF7VsaJ4/Q/QEkyRei+OovdLnUOZQRyi6kUWfaVjEky0
JJyO2VLSYGG8uY6YvQTZJ+CRerzDPT5m1XaeC1rfdRUWnrQ8ZeXrcLBjQXN4RAZB
MD39N3/wXySLbXnqWAlY7NImNJaAHuu8W14YB1jf8QwWS/f+1es0E7G1Q14v/WG+
O5BzdGv0+SaiLg1wILffWFDVOHZnFrCp/IZUGtL8iAEYvWQesYMJ/rrdOOIFINYE
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hc4DjAj0I/vt6yFZl5gkRA9At6CRsco1fIZoCVNBEuRfucSmABgZkVU+ch8y8N8l
ioDoFDExlwIVtqt02xkSGWE3mjX+9Etd8Rc0dLRmFxQE8CiaAsaZk/arzSipWUZI
MIglK693lAXGRXcixbmMB3pOLZ0oeQaJD3svH2hugOf4mzpckzEHT3mM6sag8QoW
aBdV+UeRvViLnJ/jkFTr+j3A4bUG39DWaAKd9aFiVJfdPXJzh6qeRwF7s8SGKhtx
ku5/9BApWqe2Gbk3E2t+Y3nt68pAXnTncTyDsdHkwFeF/EVCgbnH8wAljAbOp2tC
43qLavljRIaQlBFR4NPfmw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4768 )
`pragma protect data_block
SGCwHNRs9gYpcKz+vrwgEGGrVdBnpffOEZOeTrH6yiyz86IDukV942Zlk9hoe59x
n9dc6zYAFa4It+JR6SyyYSEBSlcNGWW+CF6ogWWjn6pP3uMsNFmODXtZ1bHbhjjp
iogZTGxItRID8jKoOqwz0Dq6wSH3kTpbujQt/W/q0U28mTCLuLSpWXVXvNzt1VXH
Z22HHKsrQdxpLnCj5Yz1N4gCsf0xWRsEWxFGodyhHXt0vLbarYTeIAz50yp1j5Zh
tkDcAQDC2T+fVlRcL1tQPsFXWlA//guetwweL01AoXjYlvHJPSKgHT3eVYWR0Zvz
XIlrdLD/rTXarnaT5E16aEF1I9SEttwyEqR0wvjKMkEOMIb38PxHUvWt5zhdcItQ
+1n7Zc0bZc4a1mMzj/TN1glg/yiYQOpVHKbJ9WGsHdAWvtXSkVRe9gQ5i6qgbqjT
UymZol3qvixS6OG6owCAjUZEOywbjHSpKCGmqdqJTyIfSvFKZfRkNnI6W2+RB3Ky
xXBRIVXx/SF00Li9JDAMKJHOS1jACztnbJaxrIAtUKk4gecGrwfxlf3s+IJrGJ2P
9DrGuWOIRMaxmKm/wppZhE/EV/TQjzKpyGktMxXFMVjXgq9lGGHY/0+3EQ0xdWjD
vrZ0igFYA5/6qTURJ9vk49d+VphAfQ1cBlEtYhVmPFLpDnePRGpse3UJESci8oNs
Yy4TOYXGw5MN/4D5FcQWYFdSOarlkrZlkcdaNnawr6ON2rksyHX+tqMYqDm6f52m
vg/iq9KZlB7lckgN0QcRLPUxYQO6PyJFC3vMo9n62XZd4pYCiJ1rg754Z0jGCIPh
VI/iJ/gaBh99ioqhCgprZpW1NGqpPxiIOBcCzeW/c/VtIT66S4ql34x5lA8f1AzE
zM5Gvdf1DjhgMzHj6+IghQRogNFaxp3y/1gFVphhMRek4WAIW5ahaLBbXHMzqZOR
WKDzRuNwMEd6PHNjQcfXRRmFhlSOGsRWmkiG4WGY6pHtLhbo1jsAxBRev0xV0qTy
2EnDBFmai4GZpjNrzBQnk6sWIm0XPUyElEAdxhWUzKgcDWllN5w7a6vi7rbRq96E
Ptl7WHwhgjPog4PDojWCC8OoTZji5Xobzzp7tF7QGLExomhoRMc4Q1iswVDJ7ivE
JCxxDmRkK5Ce8HFSaqTgceW7oOaQCGf0TptwI2mH4glJzJNLy2OIXK6Gn0HE30WP
hPR+BSpln34N5aUvLq2H8Bz5qm3RHMNwd4S5TxIqfVkGGflYxS8JLT/5oTbmY1D5
YAb+0T8tNPRccvEf6ncjUxqF45akU7t9/ksjbuh4F27Dt9I3WVIqpYxemlx0k32Z
TaVz6OMSmyH0UUeIG+YM7a3k+3lmkg0bqp8X193gUXKPUprssIrhFeJsLWJ1X2Zn
nZ+7rZhq/Zz1Eal2RVN9E3DZT1MV3MYzT32im6k716SDqFOmnnwr4W88cOUNonK8
74ICM/PmL9ky1r49iAdGAd6/hFDHeXPpE2TQ/+b6HVEamKHWZwV5wo8O8zgigMPV
yLg/YSGLiy/Zyx7vdgTDbZLKXk9XwRLyMPHwc9Zk1pWMlTva+c7d6WakYUcfoN9N
TYFIYjwntU8ZXg2dxh5X4XqxQ92r+D2Zz4+N7Mu4Ir6gCxGB+aP560JcHx/+P1ld
nPCpMhnSaDY64nCNYj2WVIA4th2Tc/VxpPqH1RN41BOl5nztcbFojUU7UAqe49eK
fgwkU0BTYcj3NDE0WZAgiVUM4338RDntZYugwj7iZ4AzJPM0ThbGnjZzBeqkYSrt
T1FLVttGcaSHxCgAbDOcjetDt9UHwWNzcZ9bAiCdkF1GllkukahCE2+1yIxJlEaE
D6IGz2aQc/JPVMo6z22gL8lMcinjUWiNcfAmtJUySeoI6524Yh7H/6ar9mgjBBAk
54IO/+u+ESnQEQraMUtgLg0Wkxvsh+IuPK1GTXXLamG0GKbkJbtGPvkyrdfu7Tgk
Oh/1N1n5G86QIrZGj9cItUoni7uyfm6T1TxmHJcc6ZPgxtSL8IqLk639nAUWcF0K
+QxYgSg/mF8aeK65kk2ac5W28qthgHLiahVa7NuD6X85pBn+PoINdFJgGOkIZBGl
QbQ3Wx97olKbh3a/sCiIjudZFYtMHmd9bcF1KSN5IJ0/AihOLgWat5qVNPeLIk9P
Q8xzIb8CdeHpEqO0yrC2A5OU/S6awg2+8G4p+rBWmGgyr10yZMt6y0hn3j4OFn67
M0nE8ZSCWMcuruTpf92EsXXjfhDOIoAr5z+E7Q7EcOA5mRZ8Gd5blS6QJoZvY5dr
WdcETFlOYOcrtW6VgPrbsdaNxk3mwoEv0APxeekwpiNIvPeKbWZXEosd+dW+dQq8
zbvtuuGEKTpUxmEIhD/Utw4u/SyYbrdGI9lWx+ne8RL2BsEjYX9rXYsfz3RkMV2c
EmNmTObquwt3vkJbAyRoHX4S+gfruHAh347BYt4HQsozeKYk4203wHU1bujalUzG
1ORlrtGDeHR7Eh1+E10ax+anxlwVPX3VarP61xl96wzKtbfM+azO3BQR+AAb1/VN
fKmf4lQ37wvTqBRIkM3TExqa7r2UmzJOxUXWTEer95OAU0DMJKZjrj/lZ6gWXIjK
Kp4OqcS74BTmK6oBC0H02aT0rQKDv6D9J/MmNlfyHI9iM+pCN2PLL6t4T8Jr7yw4
W/rAnq4hjuMe5zmFc550dUjy5IvFlZlcZLP+tbEaE0UhHP2nC1CdCaM9OMFnvZ9G
t3dpI8dtgGTsWRhYuJSx7PKQEUoBXXSgdJNLOyDvMERvuY3VbPJYscaHn8t9GMM1
fbLvJP/hqtNj0m7cVmWK6E8nRvI+cQ0PjNtrhMjwQI3TH1sKSEqmm8WYhjDhcPk3
nuLs9Jqz78gHo/hb/QByokCps+JO/CRU1GKXATmxGorHeLSOvGukoREjoCqTM0kG
C9AYE8sCI+lnzrjV01K+m+sGHAQ8talmcPe4uh0M2vfQbLERJWmYTAURmZvms43p
4LBgCylxrw7/Nvojh1aFHJCsSLhDWRwlNPrN74nzI/JN9QaojceWM1FLj+oGUVL8
f4RVyKJ0IJWs/JHqlW4lHvFJRQjlaXI1Qet891VIyHinD2ON3bT5eR4IUPs5uMOh
swOZvDmdHUic0aDZyHHAE9Mj9bGK2UeED04XMgRMy5WTtOvtWjYvySNt/2qsy4LG
NGLmAuSHtkeJz5aFXlRG2/V2X7wq6RYusWpMERS6I0zblMV5nVPsxydEDoDTQCPo
Fk9kcC0t1s/MIUUhok5C7IDLCV2A3p6taS36184UU53nIEvBaozUaqxpGr+6mEhx
19knQmT+EOcBnf+6kyftzIayMIjdnoiomMi7qNbz+FSHScNEwLCw58ZkhTw6fXjr
JeVu/OdeEW1lO1FakqvbSMJZzhA2QcPi5TItRJ+E3QfCGycRbHcQATMvM3AXQpe1
MiFslhE0twHjXC52Upx3DoZbu6u3NgvB4uuThDYWkR7vtYpe8ta2eg/2F+b5GwTa
kgVZLAyYgs4D1yiyhUI7iFHf/TZrloNvDqh6ZgKe/k1mkdVXxut3Ef4J0n28tA3Y
4oPiHAADM9KIQGeFMUsdr+T//5lLiaQHLmFCVcCeHDAUd2QwYZd3/rES2WxDgRkA
zZUmce3lMzUSpiAoktJAmXiNX42v1jKJcqHK5gflIDl7oFcKKsh6Sa+/RhxAChdR
/2CaqNK4xPZBooLF9alroca3LYPUeTBXo/fJn2yDg7AFt273uF7r7rbcPbQGlNuQ
EP73tbP0SFuxBUKpL38LCHtl2s0M6hOpF7Vf6/MNKTlA5spfXjZ2TgHzjGZ4rvgC
F7e42nJSyDwB+Z9Zfc+amme04Hft6PZK/v2L8BVubjyV+7SA7mxUAPBRooQQEnym
irjew+9Lxlix2jnDdbnS8esdDZjJ/F46n4VDiMHDo4Z6UKQwfA0bW0b6cf1lz30q
rAl7u9pLP5GOpb/hLYW6SjmcYiFHxc8wLEtLwdrI1MBOimP6gCKaV/noK3k+XwlP
FZgGLrq+aelijs9KpxkhyZr1UXdTVi4UvLnQ62VAhti87P1VNM5YURHzGpBmgLJV
iPPtXiwmMFlg3GbGu1ISsS9+PqecdEE81DXajH8YOlGRcgV2iK3r5WywLtUqGuMs
JvE7cK80u+TOlWZw61/3TI7H/RxCICyu1mwuFv2PQ5zAr0aOJ6PzaTMyxYP0U8Fz
RyEw4h6UN8XWtNG+/hnPIkJGlEuMuCzd9temsQFfiNeVer3dAYbvSE93SGL3wq9i
Od2cqG/JG/mJnhJzP+xVAxO/lxMLKUcQnnK3Q63ksG/6bZLvDqPlW8Pj7HLp2r/I
le69y7TZ/TgCCXm5p2eS3+ErNKnEZvHOy5k3aTo4x/sf8dJHEEGluQVe8H6fvnNI
dcOZCtSjPF7342pkF/g70lLP8Z74rLyfD8ZsUyn6Dfqle1mZ43Y+1+mpCm5SaT8O
iPrvmTgD/JsNbKb+Se2ihIs23t1N16EL6XwDOLz8DSkxl0hOhbvXoAMHysfEi2te
WGJqoUqg4RUBVyiY7Sp0ZwEnZwSaCNW1FF0kTCV2oPxE5gC9p99WQgwtZ3pR7R7F
MlTm9cJEeCrAEWDEI3jGYdjh6NetFB3+DXHY0N9caQrQWQw07m82lXh3mpld4rDZ
ZqCe4Tt85n9RRJ50NDBJ0gDcTIv1SMAQvzpbtVKQhZWiXrbgA6P09rfQgir+GNI/
byHzA+Qn121VEpKl1z8CFa83fQYvqGkYLGvUlts2g01VT1WBr5EwbgVCsbHQARpp
Ma9ZbJeSx7PyU8gGJoYh7sfk88AHr2zraHATdsA625Y82DowzJ2rvxVQw5wGzQCZ
/1Qu8nQPi/kCiTS9PVXr1eB9uEenCtJWz9GXZQnGLsXN4pjfEdZXCYLTYQ/gGFxt
SQD56kNqt+9XUqC4HE4M3MOLp9hCPvq92jqwy8jEaFEswoJ+INqd/j0tBjiF8o8w
URCxG6Q8M74ERk0xXKz55qt0nniJv2/A+4AqyOAzt5+9Zlk7pqu1TEfoVUkR2DhQ
4vDPWCPGae5G+kV3h8+yFKZ5vAFfUY1R35/S6nGwLzApmXnVNF3Zr6s07TfAOoMT
DGRxcmAqD3ZPQZxvek42aSXfv2OQmZ2gkofLh7pF5FGk1/c74MWODv/uJFBBRp+z
AxZP/xAebmZcxNzVZUi5xbbMS3C3wKApbDlasapTrx2dNhDs07xfYXNIyW531qI9
UjJWZqF3x3paRDdniDIL/gVzusfL9Eci2GlZla1f0uifsLKRk32B3LuFdVwF5wmU
3Ba9grAsQ5c6egyRYmqCVBnS20tqqf4jVISIVPSMu/6cXv/oo0/D7//I1fikvgH1
rm1pYR+xtu7HVs+tGPVpxeLnXcGKoS+ameGz7tO5LTKyDp9osol9Q1TruuK3Kbm1
20qfbCIv3w1ZFBgRvngK1o/unF6N2wWEYN6ck4eHtX0Iq1YWPa2EXSwrqanG14pV
U/SyVem70QR+Bdo5IuCrcd0sIh009na+A556NHa/mJ8hTY+Qz9Lo4eU6O5dNgyMi
pB0peLtXQonS0/vHbFB0WIAXcyKnnibHyFJ+W1KKBe+PwP4iBZc/wsVmty/kxKXL
nj2o3E7xcv0rsqXCWDf+gKve6AH4xywx9/cJYiVoVCZAM7vu/pOfYCHUxVdhPiEA
qm+hUxVnj4Cq0xFFIUCV88Wkr3JACekz7jAndt/6OgQ/GxUKEDGQaHx3ym0HsbpR
yUmS21sii5hNUw68phkCXb2C6Kle/OupbR5btjpnInv81qGJLQUksf1Qw1FXzleS
A/eqwh4O6ZOp0kqM2GTl186ZDKKu4SAj8/8mGEyKIv1bxZg6o40DAqSgFfhCXTLB
7vSlJJDSLKJzQ00DOGMcOlX5agwCaptKW4Oeqwcxsj1cMKKU5HNA2DjX5/ml3ou3
P8UicQlc8+a15s4HBRDx+dRiCCcjhNLyrTfwtSMHS6fx2lVQZI4/cfSewV53m9vv
UiFOrswm8VlpfySvVe9lvR6Y80Go6GzTGcGQYotPHKosNRIxFr9P1HfaZaLmZF28
2sjBzUJDffgpRqF+YK56qcwLlQFaLlIIDCrk2xt07a8joL+aHYCahFOvoGIuQREa
L9pXuD41yotO+iJs34weZeXCL7Y+mKbDfZ7JiEkfS4MN/iq4WDTk/4U0J37SehIH
oeJur2YH+KCYmWiR2EwL3FK8jYusuG41J2jGx3sFSY3gEXcGimqmH22PO6qBqQPA
qBVc2Xikh8zvQ57x0Zq8/qLlGl7wM0MhdzDwDdQ7F1PjCgAwfWJP4eb5lBGAHb1T
Yw4VLFbpyW/yEPxEO/gf7w==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Km8lMmifqUXQHNXYmOG0f/4acEdKt/1Ine53133HyLgZC4LmCLBRF5K7BgIeqy9Y
yR1iRxrkfj0nqzV/5w0gIPuh7ulu3ljG+q4ZnPnBkdlru+biXKV8RGE7tzmaN+lo
Yv04XliE1uj741E8l6lPRHpzC622PdZg9j3+ImuZdtCfiAkrk1rUTZHattlpfW2e
N5Egj1z5ab5rtWcOq1VKkxfYXmDIDFoKn5LZAd7GGcoosVBWzvDvCzHHqoa22tb5
nuGBrSqzD8LB+jfe8g7Sb+vwF6UjO0Tk2xNlL+3w97hK00BbUyBOOa3yOy9N8iMg
Gsz9IXfftpuTtZKe6h3lug==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8720 )
`pragma protect data_block
cigdn/S407CGw2rK53aVCH2wCn54WJ2RpNN6mY4kmiuWRcios/Sq4w3fcgNa4Dzj
3HB37S5f6n7xrxB5Opgaj+6x4tbp90b0VqcwzONVth4gXY0OPzZJrR3SSlpDcSCy
SCZq/MHDsz+p0fPuWcsDHKT77wbDykjLzSH4NJW52zcmKdtJ1sqG1NOY3QOGflFz
x2TKTH4k0vawDmk4zRdBzszwzrmPm2PyPVSnYom0WTSg3TJGj0Aw5EhaZ6+fnRUg
X53OTmoGWdE3oiqFM0iiZmTpFeVNLKUfM5iY1hyOpPxV6NQ6pc+H6ur82g2eZlfe
DwTDNsUNdCVidWLpMJ54x0UXU7RFkcqQf7IUTLCKx4gwlvhJputDIdTmReNQU7u9
r2f2jOWzM/lg8xu1F0Grt9Ho3VCj62aFkkn7er1jo1NrlK1pitFKS7TOd3NUVdnp
xaZ66RZKlOnm56qMHllhwaAGRjbC2nOfzVEyZI9c2K0RHIEb1ulZ/s+dhReE7MBr
yY07wcqDTAWPdw4+Qgxv0HLcrCihtmyll6sVzeWDyqlfOMw39IAXPbkND3KvPRCv
lp0SAYFzla0CMo+98gDBR3Ha0j5EqN7IgbosoLLDlpd17jAkLI/BUA2ie2i8ZU/a
+7uuoKifZW70Do20FmUSs8uSWucU/VS/isHjVqS7N6tMIeRFUweWq1MdPL2uWyFG
+YCMjXuokxQYJXy3MO+RxT1KnZwG5vmavF9nA4BsD8blJgAIhTciIdmC2VrZp+85
+aJKpEN61XseWce+hnT4Zp5h31U+ra3JvM7AeQD/qSDeIFkxAY4Hj4MdFih4yFAV
ssob3VIs5RHGSmdlR1gDIz9/q7oa6hU8gos0Fjtva5ErcnfdkCK8+Bx1PiZHY1Kr
kTHHnEdv7H9KwxXOb/lY/08+ieukQvbYlrcOjw5NGgJ1dNKixJqf5HBQZwlmtj6Z
fq8iVlvUifbg3XsXrZvyybvH2uwyya1JWYbsrBuySNVf9Z00cTLf59TPv9EsuouW
c79aF3kykPSkMyFm46Kk28N3nsHVnoN8VJag6E4nlBZtIHDydaSeC7Qiq96PurpE
h3klI3/87XE+F8UTQt37QcI+aLSUGOjZmoALef+5Tj8ZpktzgDlyzxMSe2gPYTda
/voLDH1Kq1Hzh9bFBOvIgQ2EpIWC7BMdgRoRau6jCp7MGgRc1++LqX3nRBM8x5jn
7esNdLW9+NJa62EYenxd/k52sgmS15hstx1IWOJ7gvpo8rFDq0aLOW/8DMc431hj
ivuk9+MZOhd+sW9K2kvSkd8clG4wAU7WBbyjtbSlutZiPHvgVVhEpZr1l2EE55k7
/plIqGmFXI+5N+WxQWB4F694RXTRL81r55JK7/NzD6xPgsscnWHapa25IwfhbWc7
l5k6OJRVg0cnUou3LfCeNa9mZqY5Y6Rvg7YUCl5T9LIO1Y/O1P4sCqnGizdKp7Rw
24k55TZtlcC8SwvXm/ZNcs2XyiwXJUGleMw6aj/fDwmvgfIscJJk3gwEgF/P/+zs
m0qLvR/DH1jyxvF7xZH9VHnVkHSvdyUAIM7btPrKwDuGyQFZfiuZxOjMJJoMFLwH
k0SwQ+rznCOPFWMJwx3Ysq+ZBYH6gFblq/bRlbH4pq3GATg60fPi5U5mtCBdM1yR
dF5ki0PF4WcJiq+0SRojHypRKG9VyPmE1Y1nN431hurftZF3Zc5gPkPhMu7WQm9p
yN4d7MRjBDl0bMFnwSOZS2wefYZ2aqFsqrtT/ujUOj6WMMYbweAjY/LPTzc6ftEp
llyxML1zjujwSEASDn7RQTWvpmQ34Jv3KsXSxyU0bPmy/LmZJyM4MUPUGeninmjU
M4k8htTNX+VLm0B85U9lDNIH09yNgt/0ykbL3tA8z4x7WUK/Rj92E2krhVNAUey4
lxgNG41cNiFUggfw0vmog/Sub+n5G6gqpCTpySgdCJ3chavkYL/zX7qyoVLwsx1z
Tdg1TIp3sB2UpXaxrg/VGRmkBubZw/v+joQ9IeY7uYY9vOt6anZVuPGKlfp7AYER
tvJMZwoLbmzj5p6l989bX8H1OJJEtDqmDRBAWXI6NH3EOFYlEouB5GOrh45MeH9L
KkAR3oWp+qufLNGYud12DESnUBCmSXPCzhYkxA7dnux1SLZDSCnGiRjCzV80NkkT
uEtp2f7pEoGoLB/gCa356Gh2Ih3qZofAkSmpSb7NQyB1V40+7dyqvXNBKSDpR9Jc
7BEDXka9s+yoOkz840YiaCpOIJ5RdY8UPpS7Xje3C3Melsktz+CaWBN1x/8P5mME
goWJ/5Kx7iEkcxSHdbFoHzYfNYnE+W33O5jo4sEYF1Ap9vTgugDErm68Af42I33C
iv8bFFK5qKmgBPrLWM1d6xvkHs+fvq6ErFMiOG5Fgp9hhgYHdV7gAnfxsUJz02cF
95be1DhSGUY8PcXmio2WM3ltp8A2XKFAMqNtNsnvmETLAipgmngQmPu3zPBZlGIa
/qPW/BT9CjWpzRqzamQQTgzBkA4bbH+OsYC69VHQECy0yUq2MWqN1SD2nYOEECw+
PiDD2tT0sv4me0l0JaemcL9vPeF9xU2dZSeMvXgyoQtfAxoTq5lzcTuP606cFFir
felNgiHfffBsSX/H4jNASuBoI/p7iD/WfJf/fiMLShXWinsL+kmXS1MyePSCeq0r
xDSoWFT65mCo+sAqUYVtMe2ifm8BcHFO6rPure4WmlZmV4I6qxaPmVJE2g/izLKw
0HgTAVdWFVb5PcKSsbn9Yj2+mAXdKh6mgb8iayFbAE+5yaGuW1QQm9lt56ORcGH+
5sQJ41RecZJg9X5ntvD+DGjyIhRfiPDcdGyn+B5JRRD0duKntWFe2RtCz7qC5TnV
cnTCHRwXMstwAsB+7Yw9Fa6qCdxC32whz9B6ORy1y5tmnPSsoWwCWZGAl3NmoJHN
FV4YlHPy2oZV8WZIgovXEp4sxqXjdekC3sLGvcrvDGQbYI6xqQAprWqJo2pQBcHj
knN5D8NfWt4bdaEDmNmlC53o2MGKBsD5/hP6rEYYQGRwasq/05XNDxjDbiAYg5bi
4stSRgHM8sFFa0WjxzFousT06PAaYX4MZyvqLQM/CddI+gLOhzxMVrAUNZhxlcqb
bZs4jfb/Xzx3svVR0mJRtxfEeLAEE5/qzA0vEKlAwxk1TlT5FCpYXx7OfH4MhXEt
EB1lYzQjT69unnPrUjdZLgSAM+yqQ6Y7pkw6vzjK/d2v+8j4XBNJSG6g9jYghRF4
Vt+gZYTtz+1G/WJrpLc/ksqObet42VStNkr8x4mgwBCRqXuvuPC+Lk0NZSXON+7z
fQdoub6LdIG6dIgDYdA3RDmlWllFfjAqwFYLjxyq/dAHBeAljusUdeXAOwc1hg/V
fuqPllsiJB//rCiDtWLjuBpi/noyl9atD92UUt30M8bwNqe9aZNRjphF5Y+ueW2V
WKOIGqBadp6WL7P9GqKK1mXJC7KJbA3dkb2ZCfLFt4hqkNyuApbxZciz9Thn3VOI
8wXjMy+9pxzd1WMztrSFX2I7rab98jA5JQSk42MhYUkCtvDHpAVCSrDULAP9oGcl
kxw7kZ6GRBZcFkq8FUPU6XeriBnVMDI1emy0Lufcwdc36t13cJunEDWnxnNjJXsA
7I86f1a2/cOjwx393ORsHvkcgVUurdFjcCP73ED4nA6o2ycRRUzh0NK3Rfw0F8NA
QoOEvEQB7NcccE/r4KqjhGFw0Tb/OWiLUGQn3CRidq/pIzLPR8OZRWH6hDC6EgpT
TN+hVK6Y/VU1cUfWoG5VsHGWr0jUxaHIpZqOBtZKDEqs5rernvbwz5My3nitTdIx
dytiJ4ksKoVpRcccjCoc8tEiQdI32rEv2xrkQnD7m+t6cK16eLTpVSvsX12RmO1X
FYUAdZbCBcTnQe7KGuBj2f8SdeZ0fdR0xEuDydvyg6jaTAPwksAzaWPsyIXmR1Cd
74nUvSgDj35WLzj53TOlpErSJ6mhZPYFK1RKKmIu5CH2e0MxaMBzibKLaXf91ItJ
uAuBT9GFe/XYEnUBOAjLg7cXdyoIUqUy/aXIhqC55j0v2iQdEyGZljiDjL4qsGgz
HEu4ysczGKzvYooY2Udnsm1Y9hWoSWfe2mQc0X9FQ8LVvqvRnZ2EiLHKDnEKYH97
nDaq3obtOXPFNiBkca9yyX5FSvGSwOTC0hPihWaX2Qf77S11BT0lipswuXa5V0SG
UR94ABrQXe9K595zPjM5QicwlzUPUFDxqCrYb6GSApzdsXPrY6rkcOVk0JJwpAUk
4MxwQokNxtTt2+nuASjW55c/YFyC1sTQ0H8Ib6n05CXiEiGOfpBGbplknbY5zwr9
1nfT/PXeDWaF9vqFoJqKVnfBGB1phRW/x7uxIF/aLp+QtYYBDOHkEyqnifbUER2v
Y+ha6AmxleuNs4XcBWHUpPJWI8cR7jCVrmAKsI4WPZuM8X9KImq0gEb0Ma9s0+ia
mzSm0QslGX5FTM5yu26yiHE9ubPWKfUnOzYALgbpJ2gMwPPYDQeghCMJC9oyQpMI
l5w7cvTkEQ/Xm6rmckJvMhaA0IgTtLkB75YmQbDSZ0J0Kn398rsCEriOq4MqJuXC
6T49jirqWdAjAm0HVe7B5WzzflpZavcQvCznrYSGJh7bkcFYOI6F5X9nyJ/B3hlk
MRETgIZWhTgcYhYJtaA1iwEdBIPERYnsqju0bI5W3tzYMZLYwMIztigmwYtQ2TQu
u/I3LYz+6Scw7lXg5XamqCNUIqVjyZQPfiNy7AGtrcGHzfrPQ/Fl6hI04e5T4d6x
MIXP1ddS9hLK3TDm7TWSW+fUkolSX9WLRIaOKSEFErTkMTX38RMupvBmnUCYtqtp
rX71TpJF7Eng1HB7bS7Truv43XBGbsYUKDE7TL3VV/QeHdeVEIG/JtNPMI364Wyw
cd4ySxvmkvgm/hMcTUjAolMxp9hCMHRBd2zBd5tmOTLUc4wn//FdR2TFo2Ta+gXx
H3oEI7jC/2QO6XKJLziVncRcHqkSaXjIu7DXt9LNTOJ5eJE/XFazwIAVNs6O274R
H8zihu7roENmctdlTmLJ3w1TfoWXXeIcwxl9uQfIgLMOmLLflC/PsBj58ZuJOB+T
HiXxoLzD3MBlReWpxBhVXJQ2NNX1Q7h9kl2YuVqKRZXhrb0U6IOXsJpaGL92ESdg
JcRduikwpHMbxtjmwq/Fsa6nsGUjcazdUmG5Dv8ENyhA3JMge9Poayewa5BXOAJN
1+1vcWMeHSvdM68YJ/PioNr0aSbGBDtOyyrzJxlOx2g95uZTTSv4z+z+jdWwFP0R
dHIp8d3tnin5SNsrZBmAODdDUFsZAYYML63/1k6lh/xtI97Vg/2jV1yQ05Sn6dN8
H8naG6jroiaK4tG6IfczHrKrptDjq89C858j4DJz+ER1sF0hzFZo3uQQRRRMaWK2
WOoEdnl1Rq2pFoxUf/16CWMfmi1livd+JZc7te2/LaEVdAxy0fVdyWWr97ocb6Bz
QfuW6q/YtdACgshYrut6VbNf9oeyrtjVcFWLncOuAcsv/Sh9wC3vKN6hFFETxtmL
OxaFKME9OgWbSEJehP5qdI8v/LHxv0FDNXhkSIHgbWbXbyJ9BO3sRNrkecGB/LlE
OOu/MIMXV1Vav/0v0egggPQsZJrDy9SOtWZUd0/R77X++uyRXK6ej9b/lW3eVO65
MUqdboqEfCvdPWH3Fp2gik8he977EsXuqyMtAA/3ctLEGfJSmiEIeF8r45FYY3nE
M0rw+zdbfO8V9TKMVg6JXptB2NLztexrNi+WCj1cgu3aKTq8k0g982HnK5WgzssX
JeQmuuKQW2Gy/nqoRLElNjJNE02eDPgZo9QZPFTeb0xjR1/mVjcSDdzb4c21gH2G
iHvaYtAX0FxpI27V/edSc9oPMMVuRWJQlDnjBzure0Qkr1KPjj9bqsLwpXIV46by
8Zf5tljpbGzJB2JkiOVLKnaW+vS1J3UAJdx1sXNqB7YB7CdrFvLSZmdszQLJTTuM
RxYhzbnMQ95dligXBV72aflwlv4QrIMExaGW2KvRpFBEYCIR35p5Ii3l8ZBhKV1e
rlHE8q7MR6Ra49YWAm4YgQvv7iuexkkyXgWc0zZ3ccGh0Y2Ud9BZ4mB10SfUc6H7
2qUZpQkNR8OJmAa2TA8UecaN7RAFVipjwl2zx9ymem0savGwB7GUnJQ5BtgOLBWE
eiPvs6JwuhUA0qjubKTjCEvc7Ra/tC1+Vk/eWb5xFLje4JgkUJ19SLK5XgPooKJF
5MvA1ufBxEnI9xb9/Ffu90z6qWK7PG9dzFle826tT24fT8x4pxVaaX1B54Ucv8sd
TxiOmX51EptTKl0Lm7hVvZhmDi2Yip66uUuFwo8LR+/3L6Sa1ByPtmvnZ/bJ3Vu2
Jk4qj25tzktrKFGP89G8vy2EQvuzgw8WdnTZYKuwMo82lT05K3xIWrRZB8HkHpLn
mv5+6LrchAaESd0oZTjUme4P2uGonbGvpYhfqOEkEtW5Cm9SigVtgCczjqIO6H/F
25JVUYyaJ67gPSRn0IrDUDnuGvbpwNjfQWcKeBFZkhVkPcsyUOjg2guxNdKl6Ip1
b8bscmzFU6jwynlIU/L7vL+ho6unNS7w8F1C1ewRnGZpyi4GnsS/kppQ25UkumV6
fz5iNPVGz1lYGfGhPlKKNJBw2v53ulA11DIqkynR/2rVThlng7lUCsTIjY+/Ml+/
TUSncW5W3vlhPkE+9Gc73awSsCwsSBsBeZlVLNBbfQ1zazAoXMgm7mniBHTBb9th
DdwPKJllXZBRPa57cB8tFtd/BsmOrIiEjIQnTBV7fFso/YzY+T0Rzs/5m6ObVoqO
a3t6fXBeUL7nbyIvnICakKsLPTZVyslEO/LhaUmDfuGQfxHojXdGZKxhYzt1zGFY
4wI+9U6rKRCUCZSE4wThUycEiYWpku5w9QHiQKwo3yBCBXBy5VaqKRQisJv7odFa
vf7rFNn+vvuRKMbxdddBqTjfw+zBR2JxblJ16D0w+gyk7DhZy7NCqT5Tu5gzBJHx
FSI1JBcRMz89mGF1IGT6j6eLSlqe2IjUqTrt7Oov5PXDZz32VKgFCS9pPXOyzB38
Fy5OurXWkCA96tVuZ8SbfUuy8o0goV6cAU3UWAxfQDnmDHEjhRfsGMKylAmE3f23
c0iT4477SNMhaOHeMSkFmuUDbFwYh1GdT0wwlaYt9Y7eiD7STwMGGEWRNBbEiOYG
SnqFBncv0mg8hzgf+6g8CiGxIeU/ROBTh1/AGVP8O+mh9Uve2T+VGd0NJbLT+ZeT
Htnj5f5jeJylJk7QjYDan8k6CAOF5xkRyQa2fbuzpg2H8DcbRSW6kqBpnB4pdkqh
JUbdc1VzWOvz5yW8ADunqz+upVT0/8vOWKL85hxG7QhkNYPGjz8ngehxWyefOttV
XbHANNA412sRBzbEa0WDZq8vOjT9R6/U+16RQghU9VJoB/Qq4KWGg7r6KD3r42fR
pHgPmNTn6lq2MNRr9qxD8CcG7gNPSaLRhzJAwSvPszJUzkh1Y0ke5Cxymluym+Xx
HDwyyLiZm5jP7sjiE/8BEQiRsDpTo+qeqw/GdityJ96tgcDd7cNvCMcs4FyDZiIB
7YDYVPmk+8KJ/NbxaZ8dHMUQwyA6aqT5Q9xzQ/zrX6l8XtC52do9ScegRDA1K1Ei
W74AUsb0QB8vNnvu9bgypgrqqvns3fZSTCVDcoOCHys4tuaQlyqu2RLWmprMwuPK
68+h88uuowUz72AseH56dCxNpfM+2lj2z2EgcKtdmB6/DxvVai40GnM4zkKrybTm
GQdh9SiWlowm3DM1zUnMQqWXJQ6AqLsbCeaouJyS+7zuvgP4I0iKcJleQcVJZXQZ
q/esFWJrsmsovKXEGSZusqy1F7k3Hu8DOO2SRSfptUOnjnkYBpwAZFr94x4w7DMf
iI8yFdDXjCEn1mn4Am2t6DecL86BbRHtHlC2K+xzTJLWdnXpOu1dPCALlX/z2tAE
U5GTCRkvJQTGcqXt1W9yU82iIhqX/nlhW88hsuw35B8nQY0IbVaOxFw/2bO/PwQz
0XtBnNbRBN9UcPX2f9iYLe3i4NBgn+vA7f8dGJTwBItb+pfbeE74puYIKTgP30s8
ikxiGLn9Q6iXemEklYnTWZfajRc4rxx8KOu8XO3h7JD7YsVMwRdU+AHttSIPSfZQ
CGxtoHDWyn89Dy0FLS3dSaPgtdmAA94Q4bSqFXF+vrBuVOCc/fLTr49F2INBUqeF
ohBWlgX7I0vN5Zn1Z/uXp3F95FllTpGLV2Re8UvKmKVKjvJ1UTBX+6NUfTh6d2os
2nDXK/V6yZjnLb7TTvw4oFI3kTufRjfHn32P5AS9sT+vGD+qpmfTv5vwnk6Y6eMK
Zpq+iOVw05IAlS2f4OQHYg1SUVjTwIpubbjWIjUu9VlwibzKjbWT0S4igOeh3XSf
zEMO60gJesvSQZS8CdJ0xOWHgxiGVnBRaBBSWWZL+MUkVeSVN2/g8oLerWe2zSWr
jV79KP0PbaUOEgrWXlN4ldtaVoyTZm6HMUWOy1oODiewO5I3DeP+61L2MZQ5Vmqk
X8cb7U60vFUoY6Exoqs3jLuuTMjdKQVfVzBiTqE1ECgKCdGaqNdIvRaCLxj+g0h9
4d6Zc1GDIW+mUkByafN+w17UGJd8m69FTEFaG5vhMHe/6RCQyziiHstdd4xWFPvP
jAHY4kiCrOC4h4B0jioRLvGLk3xTcfbWgARshhwDqaohr2hU0hb4Mvjv1EBaHf0w
/w3StU83xLHwem43HNWdVo6GQEDXY2ytsHElpE/t11TMprlWRosN2+g/eXEtacTj
DvAugsgftzLIwj486qgurfUJtXTgrz7r4cNiT6KiEltf2C1mnZP7O1JIuwmGke24
s4nnrGJt89/zWvKJ5rPcqaaBSGUejR/pmEzWjSRjPu2oI/CHBeiWJ6TVzJuoDt9w
GRNOvmPTaGRrHvVvN59G8RF1RmiQo1isssh0BHVpfdSGFMQbKeI5RnsHmbl+H8BJ
vwlfYlalw70w//cn8FwxRSBvoFdg35BUbigCs04abiLATX+6miAgvT3Uu+/I54N8
s/HV5o3EE46EQ7hzaNR2utttlE5BWq0KM3DG1kFk3XGgbIwcY0stHmsJKLQ32zyq
WLPlrzDAgpunSaCTDRES6V76Um4JtqBmSooqCdQ3Gm6cMRPjDFPI6N+WpDXHc4J6
5xle5zSyXnIUU42dfyohRpU77GeaK5LYWtd0ZzREuKYTBH/gbYK7HIRRzLO8vNQ6
JqXowQ1NiWoqbw3+lMmJsqt8DRrJ0x86gdZvgUtprtoiTviCq41huXa+pdc/qLL+
yazKMqQ1+Ga8bRBOzlo9c+tZobNmKzg1Jn34jCdL3vMEuiabGt20hPf7v2LxqXME
3YN3HqG5UjjWGxSGav0nJ13UvpK9vqDM/eozz3rDsmXJbjKhndoa9oOIc8m76j+K
yJHib10pS8a+XLbpXwePNA9077iSMuGzNwQ2wh10UridvPmQtG0SfBuc+uZ+F+4w
SsbnlcDs/YW7blIGikVGlXZgUvePPbFIjQrixNUCWOYtpC6MNnDvYmM320N861Kr
jVpNPJeF8xdADAkMRYy8SPBWwP8EXxehr9aiZV2cFd0OQYCKmIStf5JaGFRmbcQi
iTgOZwLFINB8aitFP8R6vbmJV/wwhnl4dqvsihZtdV0zDLyR3nDj1yRsW7zTIYHE
Z5xja0CHLu4cjkSeLtN+/RxCE/aFaKQF7XgDaD7QtMJKpo8qQ813h41kTF5ow0df
ZOfcBWnP2vJfh1HwaUCW+xYuvsn0BtbIe3grSsJID5QfCneEqAT1USGnbteZ2MVx
GRjF7ENV0S+uiZhJcsZWftbKbi2sF9liUUZKZbzzi2Zsc49FK20pfnXhVbAYMTWz
JOL2irxUCFJmsGhtpOz/yQzrTbo3PlO7da17yM3Io2kEq8hDPdSiVujX8+VbHNPo
qhZeYz7557+uW2eoEpt0Zu+N1p2FF8PKjXE9tQ9iXOIfQiRPreTFO3UoXJKsFa+g
rfvPJQFLPVfjN0Mw4SvoWtf1GoLy88wp50q9lQY/Jcu9PrYFIxemrPCUxyNq14rH
Xlo1aY+X0whUvfm8VePL1ex2RI89iKFhbtaOWE+mci0Ti/bl5fk9bdamvT7YXQcc
BU7PhnQVdQvw1khEvmQkR3wSbw2IPyjJl7CN1I9O+/tf55ZM6TecBU0aBsTpxQ7O
COCqwkqlm+GeEfvkDVZUdiWoKGbZv8Nt8+vYI3+FFpfPcxOBw5jGK/VMracjS2em
0wozVRWr3Jeb0Op3h7/baNuIR8WoHCgDd8pGf+W0+yqvWdI7yFWvauiUVlJUO+/0
slVeZsBj93SvUaFXdhEESey/3kaZZ906Lr7gN9PIB6BmRmOVgnep/8RwsS8zlpaM
OGDeKMiMm/4krKRWBfZj0dzCpwbgVtLBGX+CzABAcjtEC1TUgK4dfPx/TR+GX6s9
gTT9JGsW2njYxUITASKjR1EwOjfqZMcVEh6rQEDdgbkLwkIEDxDtl3OrtEVRuvku
DZBXpHePR3Rbmcq7PCkENACk82ag+9ySFU2X31hJepDWozZzA3a0RlZgZUnelVhZ
hruJwBM148rtptUT5CKgSi6SCD/odQAodpx6/E2qJc5fKx1UjAGRpiPU1G1KAykN
9iNUWHl0C0gw+zeZMbDHiP11HjRBMED9jTIIyTTEL/50ocZyY9ik0OQox5huGBNG
4U2JrV4XRT4w66CCUvi/eB8vwI2k2EJ7seAc4Cjl6UuwRwS5BS2tbA0kWc8yHplY
0TfDYo5WK+r7Ysii8v5Op/A3GgnYnb3Z0CXEfygAoFmnR6U55Z+RuRQr8SK0u2jQ
fLVzxWflh3Vp8xPadFxE+bHf8rn7RnYz90r6Om/5DYC4a62uNI1YBpJ+KnRQIPTS
YjM7rpm/4VtZBnBTPK+HMo7YDeMdCpW//LV8eOG/yu/JgbYuCUFVx+7ILGGrpyna
W/GwCDEPTej+oPK4M1pIq4AjKq3FLXQ1ynYGrBFdrunGxAq+nDAvRejSmN6ykmm4
fBNACoCSk3QChFq2Wb/XQluxP3vk12uDs5GWf0WCbyyvF5bf8I1MWD3mOhM9HoHa
XM7/OfMp9X0Mh/b7x1dV+xjOFCDBWj6YU8SVpMJxNwJGhFqE8zbwMpDOPR5ClErS
2+De7JMBhLpRQe251bY9xuMQkads7Akjk3pAn7RhJmbhmATKeik5LovH7Po0kpSu
RSjCTgXi177eord3T2EXLhWX9T7+DKzxXIQiEFv8KP5MG6SSwwM1REjxdTiQdA5M
YwA8fL1Uh8hyqHSIOSJEaI383cy5WILcCMMgXl5JioxX3mnwRRpg0auktx/qdkEh
E8dv2jV/prNdgXq3m/28YJ6CCQaGWqi4BcTcPrGuPMfKyKu3ZBm5VqVRYMUyPj3Y
jFTooi5jSeg0mP5gDN0IDMgchi2lxUotyjIbqBS88Lvn2eZ+c53RMimLr3IY2TGg
DkJUnlVW3Z2eYLF3RzgCgI3uSV9kb+jlFzXhsKe0DgBXy/ZQrJ4i6cPkDYLCzgPE
2+DDC62JcOvMqs69KVkZDNQLZ4AR0xdqgxjnJOyaliY=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ASkcQ4kTAWVBL4ynYf5ZMU2oHG7ZM3MmsrCJnVqnS3FnNd4ynSgNQMwrXhvPTBGl
AJZnkZy00OMjpF68VoHMb1bN2kpbgOIoC/SXgd8VoZCSzSHCn/eIIejwkbdrBMyG
Am+xB/ZwrA+PnV82R8PrxFWXTsBmkCxclSaAfsafW8RZSjBtbQk12BgZebJJ6OpK
9afZQ+1c0mXGsNsNrcJaPiYP5CWjVhpf3hz+A+jCrzXEEx4HtCRlCybwgQvwgpIa
kwcEjWRh5YiOLqd8jXpP6PpeE7O+51h2gwM+6R3Tu8epPhFxc7y93rR6XxOfweoC
G84YjHVSMtSoI1fzKhBsCg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4336 )
`pragma protect data_block
0GHLPLl24iMTpCe4gSt6tamsy5KeBj0QJ4WsNCJKlzDHmgSNq1t5z2zeOc4F19ib
d/OaM0mYlzeU4KvOmxG15tRSYZKlCexwgeU0cJqesn8Msv311l2HaN2yMVJoLEvy
kKFka0ljWRUOLijTBdPj2hIw3toPWVMF2NW4OHI68dKzDUtm0UzWLHDsmaiwVatN
lEd5L3E2pE9sw0T2AGwcwe0q3vzYhjTWoIhVAC9JpbkrdhvceHwnK0fgOazrvaS8
Z9WBQ91KvKyZNfgSNM++mM7PhZ6128ExWjHTE0zelDLGyIgjbSI/xzC5eKfi0Fct
EO1NZbEPj/o09feWP0yZ/RxPSRhjyAJk32oBK+9F4kqn+Ld9xS7t0HIskK6FQYir
BMzQFB2fcT7978iaHtDjir3Hy4CBy+S3jQNLWEdFY31GGAf2MiCXPk3FmB6U1deD
Xr2j1EYm03kKvtb87BSw4WPF2s9DGdN/EGZiqDvu1aXkfiWJw4Pkk8wcrNGWWEC2
PHzFNWZ+AiqAximVE80YYh3okEUZvkCRjecTtPCMgee0cceNn2D2XR4GsR2ruCC9
OiSGHtDHenGZgdE55eaTxw78+ov+G7jXCMc5kX/jGbaZ7+IRaDoOUacT317LUqQG
IYG+AWqvPPoMEJr4crY7iOLdYBRJv6uo3I6Usa9fm7e7YtWbmGcZ95BdtsRFIiEF
27AStepTJYXtAJ6YNeCF5rxjJEf+CLjN/tYyyQrkFbk/XWs64sB6J3DrDsSpL4ra
MKZ2iqcyL6oyyxerr+EFNIHSc6Ef0DFVk/HKdQHDvK4xj2PMkZtYdR0u3VDz6nfH
Uy75rzK5e7XFOnmgC9zjVPLILWWt17BU4sVCRWkWgLePA/nlyhKibbUHOwotgcOH
Zx2gyJhc0Di8KGPn/SdT/JRMIx0iw/rYr8p5NM8GrT9XyvJ7lhGVyVinYwJhKa6i
rHWLB4mTkJYKav71xg6f8uZqcUG/1XBtkh0/3iJ6Kp4bLQkJ83UHdl7OpmXbufcA
1gvJg39l5mtea4w8lGg+GM6vHYv6hT5BcCSnrM5HV0PX1li9ojUa1KlJSyQU3AsQ
1aknx0eJJ8lJUF6PnbnaTAcCl4XBpC6s18G+FWsdSrvhSOpHzNp0I3M9cpURQtN6
6UyMCfWdnem/u0WjDdjyL3XvmC07b4PQeoX5uoYQQyeh8sdy2U990kY7jAHEle49
oCOWQ4sDtffvqv1TKRAkDLxNqwEQl4d5n931Iu0KxsN/gOD8YR/uR01Da45eeAQ8
bwQ18gg21QMIGsJpBJg0ibmJhgc/bjZcbKbZTmW/+orNUp/Ml7GdbSWKCn8x49J/
Nfr85Py3ueWCB0y7JNFkYgM38qc3c/N1SE5kLn/6MKI581RNZ3j7Y6ENL/hPE2/c
M6BW42JjWbWO7N0f8DB02z4W8Y2l/aRYjewx0XvCMe2MM3F7K2sr+UF3yJoe+bC3
XajJFodHqkF9u58YJ8V7LrUYNWtntC0hVVxawbVEEcZmxM27EC1Oqjb6BVmT2+Oa
Q1Dj/uoGObCAVva8rhWuZQu9A3zfApdiRpcso114NAh+YqGL/GO6S++Sn6TeUowR
d3oGMOJhY/PfD/Ez1i1EpBthB84r3Iv55ZZkIdeovY10YthYqD0Ol0k1K1DHzJv6
eZsm4Zf0YQfubz0fC5VZDwzCVjP3DpKiL/Fogc2hqHTwKIcMDsRW4ockJaWKRm6m
S1qko5UWJEOqrd61pAJuWfI5TSafzQLpJcbVnF7yx1SVX+pgPR2aOv2GgP9lZrcq
pdB6OSfkbT6oM1qH4ha8DD73NYaZKJywsiPxEinMwe2aekvpcKCtSqkF9jpIPpQc
CAx7Y7+HMuNmo73kQokVG6jvv+gac+ZVzLYfGvsQaywyKzZ1dxIEkVhW7KEnuYo6
VW8qRjkKzbNZYMRuWji5n2Kl7EapxMfVs8Sjg382FWJyv++jCO0Yi6WrzrYH3Sfd
ip3BvriJtvnuHgBbQ1BGpozQmaAZ+LfBHv88TJ7kSR1liRHKITLmyUvyGDayxs9N
VIz3cTeDgZEnKck9JuQiP+AdZdJVcRyvNf9ZgaVWPGx7raqen5Z1kE3dwRFi07Ow
Hq5UaFZjXWEgJcR+GXs3K0Xb5tirQDAPIWmAA7aVQNqJCNYCtObGZU2wNNmv0hF2
x+/JlnaxJCyqXmYxpALlKOIEwIVEGIdfKl15/lyyOv09ebxLmjYoS6Cg2d88voxX
H0YrhKbAPsAVRNVXH6qPPfPcGkBISjd1YzWj3fmPsULxjO/ipl4quIgHuvJVTZZT
hFYh/MqqT7kwBvkUeflAbclRP2KJQHwZnFafyf49HMvHS/86bhhynJuAEQjU293n
nfTCHneiZ0XKszyNn/icMFDb5cH7N3ZfIEnG28Dgemqf5zPcAuB4mawnXO58beu/
gPfhAdmQX9oJZS7hMPXxZpEI9qTvF8+rEY9lMP4xaMJNfSn18yNwucL+CHfQ5JxN
yS2NdpA3QlSpl81VP4MyYDRm4vw0PkfD1LIZc64J5sLyreU/lfdDQIYQRer+XgJ7
z1SB8n4QqYzqrqamFwrX3ammeKX789bh8V7KRYJJJ6I9lZMcdbMQ42rccYS6mUzZ
nEsaRyDoyavWa9QqSYEC1gQeE2KWaFnvrWiTcHOqySK4mPFSyb6CwM3tNlYv3Y14
7V1s08f7/Cl2/g3bZZwCLjMi9RnFcI7plJXI/le4/ozkhoLjGG0NZEScU40Z5SwY
ShGTLcnKuhc46H2r3q0ybFjByKDZx9c964WMOtk61hcVl0lrSk/LarR3lX1Xo/xD
X0VQ+HJ4ABMeXTB1wFvEHfMal2/XhmIKYrEgkA6CgQblubBQAEPyqo3tZSGJ9ouc
T59eR61wZtQ/6C220Ici6avB/QEy/ckEXrCi0bgxV6eU92JSHnkfyIzUpN6cBU6p
U0k3pj1RqFDKEKbDb3Df3DVtdPN9cM/8y2yrMCcSF9ZCboiK2EijT2JroQyznWOg
Vezmhp9SMlx4nJ4FCEdFnANgVRGYcVCTK49DPgKJguu2tO8IgQDgDr5KdRi/CKT8
xV14/+ruG17e+sumSKN+06dINdLRC9mT3iPukTas4lCQKasEvBSFL1fSI44oFvbN
Ue1ZhHVRgz9RQUsQPEqeEsI3+600OGEo/p1eGHQEI/AQ0SLeC4VXL9DKPM3ZRO6Y
5TdiVhiN6qmVRH5iq0MstUHzaFqFBIArUXdqhG2vS/Dv5xL+sZYxLAeO7oSR/Iqf
XNeTw2E0znWRhjTuA21UvrKeuU/nklIX5b2ArpRV0vd45QL09+T4GH2kt0RoMxcB
JqH3BKmhAD28c9Re6WKrcd9Xa29cg/rxlpQ57+1elCuKy0XYz/BWywIzu02YVFbo
bo92KXnv6iKwoQLJNDxGm5tF/QIu/v41SqoVEeljMasKGVOKmCgFFF0jeVQkiPwh
0eswKvaUr99A7qAnPl1AYqLf+Yr9maKILiA0HJudQVlzyJW+JHAQ8e/RvHzzVpLA
4hy4mBo/95s5whnJ24iU2++xBYjKjtS0r8Ka5TtMyVl+GMyWZIRDsIszHI5Dd1NH
KPVEn793l9LaFRZOgJz6EvZS7cGuaioS9vrG9UjEvlYb/FOn4XfQy+7EAx3VdNkV
0ObUajilVdC/L5hQEPpYF7qQMws/Xs/64OYpVdhyFzIDxHO7tK08fROZn7C8E4ZT
56TMZP9JRPBVv732x4zFejTK+lp7gLu3vWAk0zGRFb79slJEpHaG/B0glxAzsVVr
5NdOh4uSPM6ZsYWjZyz5hGI+QXTeeHVPeU+9x06MwAqP2LUNyA4MpczzKWKaHmto
0JTyw4dU9a8r/2KsVqIwWjpUnzCz6MyfdawDVyuz705Cr9tHGIi1/0BQsOh2B4cO
lffzKPA2qrITxYEa8spurqzYArrL8HtysKvCsk9tSbRaFDzT2kbXEOBQo8IopwfT
89U/gUtaDSM5C3/+cMTJLVBVh3PSHLEftbeq6hHf2+17cMz37CYD60c1AgLUpxeZ
3+LbJMTAb8BA96i7Sj8sxZ9k/ZAO/1sC+Vbn8ZUtIcAlV1cV6UvdQW9xs3/jqorw
APznAQcmZCyV3+SdH5ogSd6vrs8FOr45w13XEfoUaB1g68hNFAqpMF/AzyQ2pXGt
iyIPYME773db9W5h2YrUPgXtwBYzULkqsqAzsWb6M/2xUXC93HxYkM8fNLE3DNfj
kKXmuQ6Dd8bTxYn5DsINTGd5Rqlo9XpN7U3Xl2HrcuxfIgaMF0X8pA/Fe60mIN3H
HsWlmQMSJXrC9Nhqc8hPKGFq7Rig0VaqesxdCEx/0nrbVopNHsKbeAT7p1dEejv1
GiGAm/C0obES5pp0qStSFwPF29Nqir414rTC7u7cImeNTLQleXchmI8kjRaOPyag
JD6r21Cl1Osy+PyNHxGLF4Zzfyy9aYIaGQpGQ4GeV9q9CqxHcgYbqfLLeqJDCpJE
wDRxW8B9O7hCihQJ3tkXqZvJ5ZHDH8LmBfxtgZBLey2WxEZmN1DfRG3LoUERVFfk
CBayLg3dYEoqO5D87w/1aJME7haPsqXXKoPKcK2U/lC9lYhCjC2CsajkYrDBEwPI
RpSB3VEQal0NXieKnSf2dsskl+Fj3WgTyF9SQWzte9WvGK7dxsOp9HLvodaKPhFO
5JFPTCp8kjTSyfGE+XXPQt7Ue7xCvpZF8E+Mydkcj3n8iUtAfdu653T+B8V76uX6
hb/8hEWw3afVv6I4xpXiHxD5gp8a463lQWjW4myntnRWQjDi6aWYNCiPvpQ9vG5x
dUEpsBzLN68BNfqPQrEszbI54CGVXwO+NCArQ6++vY/Ls8A0AzksA3fzUsupYGa+
+/wVwpDEebg4IptkVnvCJpNCRV+qMcdViTiyRhZN7nZO7qvgnJjfwus0J4BosOQK
EJWGfLkkfuegppUW5QQih5UW68mcYwW1kkodY/NNdzLkKmHmLTUrR5HccAc3hc2N
2co0VUItyPrr9Kh8EcO/vrLkO84Qv409LSR7LOAjMR9bZRrXccjB1WmtMl2offs1
OxWQArsYd90HQBXWE5sg8M3vhJY+LnuRI+IWB3qvIAALJrscn7dr16iP7CZIbud7
FchlEP+ShObrh6TxtA5deo1t9N+F9o6HMqWMC1s3XbdRDBmfAZUk7DOjo9HwM1W6
GhajU9zqITQzYOhJ4WC6oFLSnJAZ9bLDuqWVelAwsmYyKR0G5CP46S6rrajoyXTF
aIuLipzHK4OvR0BSwX41wLIkNF72hhCLUSjVrsEwg2dAatqIXPerDn2n+ugu1hEC
OppH1IVwgrlosNwOsGCkCh7T+6+36MYUn796d1v3xViE5/vDuNNX1dCavTq/r/04
WoFdE+/46wH4PfM3pdrox+gP1SAhF/525UAcfUC+ZHJNpLtXZylrFhwXLVSCsSuE
FXjxtxX1LgvsM9JlqtGACn6gYnNU7TkD1ylvjjpyWWi1hFlOgCfetwAJbWOm+uFE
1Ogi20rKzywxTCvgdeQ8wPIx6n9qQIjLkn0CTHbBUOHjZM1wJlYcLUlGPx7MEi/h
QmXLL9/rNIyu8iG8jUGoY18cUVyOFb0oYTpvub79n/nwS90lcChl9KYCdxEeHO9h
reF4aoVXb36wKID5wgwWGif9ULGg0OaRkHs3GdT6WMhd8Ip/CyA0aV7PcOdYq/LV
iMX4eX0YZaevwmpkaay/R20voSdRtBcvQaOTX4zCgapmW5EY+S3eTLNRwvaekuLw
cfn2QJx5oe/p6mVwZIV9NQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Jt6TT6R6Y4sf5AfLAsiXm/RgyEv1p2QjtT5Kj24dLaqY90Flab/zzO6qLSQl0+L+
nF8396+94xyOdd9kk5cLKsgQvdP+pAATkKydTfkaDcp1IzXg5rlhuRX1xqQgM0xp
Oo//7kzgr2835L0dVFrxHvVk60tYZKnjKsiBVDDP39dDZZZUABBGqhaYXMiedSNU
icL+j+KdXsEr9rg9LFtaUjt5espjtbXA8qC7XRgU8lEH3Gc3x1KpwKNDL0VW/7V8
EXwxP5Ux71WjspN1zhhmOdOkYhYgPSAXJkJ6xV1pnO5IjLsHp4/+qVtUU9VmLOAm
wdZPJlxnu/Rhf+yfQHA2lQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6560 )
`pragma protect data_block
82YE6u4idb7tlBL/YiYnt2rxo95ErSvtMEf9XWED0ZDW6v+L3b3C9zHo6H0fx/uO
5tkNE5w9TsRX9H2I+S/HZJTQ+ARhqPIFdbmENdHw22gKbDavkm6Mrq0GjxCXzSHX
tNpaM8SLM1YOSJTz6nQnJqPuf7kL9PPQ8FFO3jWn13kJD4rdAJwN3Gf3k6yCGVLx
I+8Rqe4pALj9GhKbP8TiVTuDidbMxoyhY9+fXR0yeViHb1kuIGccJuyPys18CECX
xatMAXTROJrDzZHFDwUi+iD4WlYUS5ZZo+Zkvf1qN5ut8dBy+wXvIeyHzXsz2uJU
+f2teOMu7k9v0TSkyJLiIUAasNasUk5k0doci6aeZZSOoPbgYcs6MM7B3+4C8Bs0
espvreQQgsSKn++17yaQYDLgfY089FAC6q+ajB18/PZRLCvGH6wNtvpaV6jN3mu5
URFdxCwzNV2NilxvguOMR/qtbAbteWJi3N6JaDpztD0Y8LFsW5qv5Qon0fKbxWnx
kr/YPGefP9dgcO28wGY/djhfxKW65c64uWJZIJGv/dvFgdk9JUkzzJhJEbkHrLmJ
m/InT4/LscP/wPlrO8FnjBRQs6smcEAAT/dWC7mbwueQ5AZ2bcdLECn3ENU057ja
/UfaowsMrnij7pcgmnwKTzK3q3yXWxlaRDZe+axz3RafAUKuaMIMRvZFI1nY4D9+
p+FUJSNXU+veI/DylNhVQmljjbEKXNPoOrcI43958+TCBzOdgsGp/VTtLeM0z9n1
sIhnyAzHwJTGq2UqIH3n+VB2rQhTATmGxyUXnPr6FwLzGlW05kfYlNPXAz1hqwoY
quETEfUYFFF16oBidYKbWOlXbe4GESbjaZTtRoHeG45o2ZBCF15r7pzVukNPp9Wf
SI8Dm8W9qBi05KJgs/DmolNJZSLdK2ifW3I0ApB62zmbDW6BRbOPHIv+DzhRxi+W
taWTnzSAdDf/74SJ/tngLZu0ATaFUMHc02Eazm7BtupfZSQ7rYe7ha11dAO0C0jw
sV1I9PYH1BpzZ2N+WPV8JLwAWYhZdDVjjtJvDVNzEeMJMshbRcKOakPzXmJCkrGY
bagAlcr0iN8dsfe4uhUzka6Puo1grqJJy36fXS1VFWq+VACmS0JMTUp3J7jj/37U
eKxG4mYqVM5sAi/G2iT7u8tdAwgfaK/3OiWF/DPJgixnUePIi8DJVWErS0Kuq8UO
eqiOagq4Mc0ODB0pjYD3pB6q7XOjlVVEacY+j3usyTF7ZnRCpU8EMeIoGElp9ybN
YCxeAico3MjruB6/Fb/ga4cK7aLRhpeYz6zUlT4qWNcPrUy5DUnsJ+hkMmvurVZ8
7+GS7Yq8N4MdUarS1UiCJZfqUQTKZ/Eqgg1bPOOUWwlhRbfYOBe2o/LvHyCCcz/j
9D9sIAwqslYOPSx8fcQEP6Vhe+Q6FQ3Ghdlt0Gie9+rDCp6XjtC0v/jdItycZCEr
43SrLxrl1qdtjdgm8gbwnT3vmEnIpUxOK9k6bJKrk+EfMk3Xdpf2ZV5KEP9D4DD+
4Ulgq6CTUyqaqQ7MW7TiF8H53N81mDEz3jci2KBrpov4jGFquxIxQw4TDERxLaa0
0U6uYoVa+5qzff5P1+SZ0XGm3jMCiSEZfSvttC0WPNqFH2zVZWc8UnAHdDjKwzdF
VSO1ExomYfc2qR/Ky/IxOfs3Ec/aMkw7HHAh6mjOAaNYOJ9tQ0kjxpi1kvSYo5Rt
gnaacU0qLrnKxW3uxB5KiXOPJ4HlYHYICSO4t/r82N3VMNababQlYFY99ONE/cQ2
UzkVusKD0ImDTD/hmpX2wJWxpOCVqwGrEzLTE+eJTNQRVksPfmrf/72EnFdVaF54
YGiTZsJ1wb174Ez+saobEh3wnCYVK6dhbyBsunuSyzRv2zclWpD6aAIVg9K4DQ+6
B+843rcZwuZOuRyHSGBUcZsN0jzCZM5Fe//WW5p8bX9DeRoLSPX4xRxtxIfnAKNm
cFKGDz5u2XqvsOi9FGNA4R32RCr0dxVJswD0def7R1OxRZnWGYHQD7yV3QhJpG4B
XtEDF9oHE88Ob4jnvt3B00f3pVNtzwmI4SKBy3VIj4fgqEM1jK0pbs0vhAkESrmW
wagTV1l2RpX72o+zSjNqd82gVx55+LvGgkZMmOpFxefVWKOJyT2hQsnd3I7ty6h/
mHeWCU3pm9TdkfHgO1C+7sH9DJyFP64LkZuWSUeX/cokNvJQ2qqkaz7AOu2G8YLc
3VHBtHw9QNNl0ypZE5H2eGKcO6eI9d57IfhSm2x5SG28bRr92nooVD48yIQOa8Zg
Acy9HTNp1PdwzMoQhZJKjfRXYqn9bUiUjxIR20eJfQrqtebMCpS3MQEhntFtbk00
4Tzwf18DG+Ss75VC/2x+D0L5NdzcbokyYTM1SzKvR5hzC2ci67loHGXzX6jqcEDM
1zsjlzGgPa7GLduarEDZG7RndPjNu6RJbNX9UW7dxMHYhUGtJB1FTBH09EBUZIWc
vG+0/g/1A6Vb1Xg/70VdvKNpYgTmfLjZwjK+uDcL+xw3n2zb8D22gNiIUnrv3U2i
JXb/y4d31ZSBw1klaOQUlGbCF8DOnnwQz+kD+OUhR7ywJTH7KPBkIdQ3eq51XPR0
pun2XfJKhPQgi4IIWYwAyfGFxBOr7j6T/QR0BheHVuR6BE6NOzSfxrf1PKNGp4Ax
Ul+kuvRek/B6pwJMtfjy4YnFtLwGOtScxhQ3J8GHgyYOr3pZuii0ex7GYpnEcb2V
qJPk3e60p0dJccS5D5uG5IcC2iIypaVDfBRTCTwEYMSVrcwnhS3bVWC/7mLywEf1
h/Y/Ku+K1TsUx3J4vmU13C0ib7LuiGZJZd5eQym2JKn/E9OYSpOlUPY8PXAKXCZY
lUZu0/ZvxVGFVtukmq+3BZ6fpUkFsqfanr3o8S395s5anCgOSiV83SGqH+DwLska
yPKLiAsU7UyA2Pz+1M5brWXMj0Hilq35BT9USASAdPl/af6G6zbzFSUw7iWFWLHy
y5dbmpblzSUWk1UMu//xdqwSs5/YWDg6Q7rARgCMfWS2Bfsu0DmRMXftQGQFn7il
L70ViT4gzBQIvfsYT/XF4VSOPLcQgfPvqQGt2BYJ1hvoFnhg/4qWjjc5C+92hM6c
i/CvoI0SEQQoDwFCbzG/IoRIlCRGjU152p/ajMz0wijFFyUZywuB3FN9tduOMVqU
ysIioRx8dLIg3/X7BabhU+FWMjD0x2JnCpxUAbQMkugLpl5h0q3SULHEgXLMyo6O
YO7P23aP8NZvTQLTHABp9gXy2nsWzAdh7/k64jZOjMO5WIBa9DbsbKrHLRSQlnlI
5yLnSN0uk8hmv0pv8di9JhaUskBgl8MOx8a8KeqHwkzHRQkuC2eK/njvxgs/xu09
WSAWu10MpARBIXhaPKq5vFb2DPQc7l7weaRYhQVGIp9Bu2hHkDuHxnc8f+zhG55q
Fw15aDHQeptHSOc8WfJN2MFa1cO2ndL6DE26XNLowVtnooBlwSPIEDIhD10phlnn
injoPwXCerFsKgZWX0g1mqBbZoDCTgCqb02PUjxg61evu37HTLOTYvm9pc6VvVdi
TPv4ioYrAuJ8YKUZ14o10MIWGxmi+b9SsPmKMdBikxdP5O1KX5r7sxDxdLKDlskS
U6Ooex8q9RNHX4dVjRgHmhmlgIPBs6EqjTu0hcDb2FAMHSt0l+VfEBS9Qj7mMi1t
YLKlnfl6Go9XCfQRh04gX45LwKBO/b2RLg6AKfHnYijbcIznyTz7/0ngJOlieF7C
dniW0YBaHihSNuR7YZ1XUrzP1bdKS1a6booiY8+7c9eAHenSkDhMYZh84MImqxco
sfolnMhDOmxuBlkvJlJUcY3ApdYwHZi+4+nekGqmbhwdVGdXlidKTYNNbfAGfsOF
Gmn5I2abtjdwNzLhjSpzRF9vOkzLtT1pgWzaVAQYkot7n5ht/AS2BGyEzm8JP74c
xCeOmq5wTugjUOyxqouAk24sYrzN31Zt7OFBfl/q3eIXqWri7Jk3D8CGSdA3Jh9C
S975NALCI5k2ZBnEj0CY5UZSqupcpXvVV5FwxB27DbYZ1yMi2NlijRFwQLTb6bwD
LCaMaePb+vmGsXEL0sOb+12Gva5wEz1zuk5QW7t4r3YTJo72EwIeSmr389gfNgHi
z22JT5ns0djo0bdoEJMkO0SFwmjl1dJrJhvidzziRroFI5mbN9JYLrAnKmU5zu9Y
m1bWwL0dCwqyOQKTqLNNonzcLhGHDC+Qp/iLezEhGgfB1DXtiXfLnaDN5PQZ9OK6
fP3kGIEATGhWTJD9PGhORy4QcIg0fRNh+3kHQX20zmokfxPaquFi9Q5NJUFrsaI1
T5VTcW1EaUFMC/1pp+HXFPwB5WuZadTcsf7JrNBwkqn+k7PMKmPzKPtO8TB2/R5E
1gxDDrZHrbEHo9FnqGD+sXMT6S78wLHtfnUjnfrvPEGLKlwcQpDPNyBrVJjSArAH
2e0qXEJbLjysydGq4Lso8UjR0m6ntF6EQeagtQA88IDG779oRHLR1XicG7FcK1Qd
/CgGql5zPnti73b5cKqBPn2IZM4LNl/Yi7cn6w6/jZWRAHAHZnwIZDMhwE9n0otI
nbn/YU4A2RP7bUdG6NWERRYhKVpLQpkFHr36qKy9K4rWdk77g+b/SfZP3BmJTUCb
b+AMK9mPp705JlR9VQpqIxy4MG73kqTFVM7+Fw+SLRH8YPd9PbmJW3MobTsAU7/a
/+nnpIw4Tc4XYxryFVTqB4O4F/ZdnMQL36nOzrCtFsv6x+veo3qdso2s0HCOP1kw
uGkNAbYzjYxBE8KuyxO/sFINVemIn4jaK9GP2pyNjTMS5vR83bhIgleu7gL7KJIY
QaXJ9AGd+OG39J7X5y9BLRnhS3yduZEqCh6VSi/GVBimUb12VE9zlbNDtpLfGh4a
w9OlBqPpEWiKTguCHBTeB7FxWInMS/3G8C3EB6rz5tV2wydXMozbWW6MGs2E1c4b
hJmB4XZXPeUCBL2ZSjSx2E8Gx/fMPoxJ546yGVrHFZLtnZri4gkyaKG9MeAn08mz
0FPvOBQz8ZTyghxN7ClDZAMgBL+wnDCFhy55tcX09Ir82BO6ZvKz1N+gLylTRQ0o
hBo65F5IJdwVq39Npa5Z90ykx2SVrQEdx3CDUvTdwuM72/hvQO4T/trmKX09dHyW
ouJhMloV1m+37Gg9rSbwI5vLBGlqK9bbn5XhcdORqttG9TYEzXiWxZwyLZ9JaGKC
9VXt2pS+YJfGKH7cGv4+WrToAYHOWyb5sUnFNugnQDrVJx1outWQcmD3p5YJN/ee
pyFEhx0YT2E2hTbUSMWw4DVqC6cSQLRw0+59KxTu4DBQQO5YACPH1F9vRnET8vjY
s4rFWipcLlSVWVXzBV5z9hd2onLGsMOzgr+zuf1bGqBiGJBiBEuVxmPqhhurUhKI
0T4DWipH/zocY9yrfile0fsVCDQW0jxmTJhFsU+4pHSoNEGrATtX22RQDv6rX3JM
X9wuL9M4gOLl6E3bd2+pOa3VUf7zzdBqkJP1voIAS+BhIxd2xtmDdPKr1Yr+ynFI
6iIF0YcYT1fzQ4pzOvMKuPVYc4Zh8UDHj1OkzD8BG7806HSJ8G2hiZJKmH2MASMB
vmGk8vz0kqsqX5aZmt1vIURzVyXKpnUpyCZGCOxr2aGWX97lG3nXXvoA0Gr4HU9E
mybYXpnoV8eyh5857Sd+X6lqOdj2axYiC+t7werRWv+6IzCh4BpF16iC+fuMpXL8
Dxa9vdA646jyuiZGXhpja8pY2ad2wXkeGE7EflP2sMlpwA1/ZCmCOl7U+mpi3qsA
wKx8bOM9ZFY9qXBZkR3lfvMSaghoUwMgZC2KlN7MKH/iVVTnW1pMwzUsGotjEW17
O5KLCgHNKkqGDEWhnCpjdQrd0E9HY0mf6fxB2tY6x7qhesLKX6YBiXsRZoizEb8b
rhTHpoBN3fnaUb7PVLoQhfMnybZFUzxIUIAGl3iwNndwGVaVy1mcu6g8jsaXfH9V
ACi6pI9Qi38TCsQFNGZfDMsB7/wEsp39JxAcXOXV6v77zP7gAmMYqHdB/deGu/0B
XIJ2J9tHsog0y+uYjAtl1kB8DmtIMfy+8MppsjZlo/jh81SFfawaSvvgzuFXPD8b
MTWy26qMWTgIjGflMu7eeR2kt1UPgJqxz3xMKX2YjVZo1plLNsljELU/6FF6TtQK
q0ECke3W9fVtPV/hjVXmZf5ma9FnrRy7GkBco/ugBMJrfjuiw6TnMecM9iAOv9Tw
5dqGliIh+HMY5johKWa2wDDXQDATHfG7fdHqoYctl7LGTpJQ4+Se8KMz0bwxDJff
hURF5xqIT0Rmm89qUiclXMv+yA+gF7p5LndOe978XziTGxTj9+CD3ww9hc+wZ9ZQ
TeXdresCf3xG/EnjyBDYRnz4SsGbkHfqzb05G2FFARReL9nPw0XBh7NAIpjdqhqB
9QYqWniqz7Bdyoq5QT0qOY5LtNb8UqllafFFJDb1Y3/heIsilbYKPv545TeJkOvX
tZJxlvt3FGKsGKxLOiGCXMA5lGJhCZc/d97dCNu9RkER+fFAvRQPg2NbDFtBOMeP
NQdD5xPrpI2XJ/u0KqBTfzEtiYcmh0DuJJsDFTEJa8f6O7cRfycZDBmwsS5NeAue
d4b0lwcNE4AV8RRjBx9AQRUNu0OxGkzqgB8Z/Otufo4bL1E7YRPCpe1lX3S0va4t
1Jh3U/wb4aSCSWblaZc/RuyJIgMOFeUMejhI1TcGtQdHLSMAR0Bab7teAwSQ57bM
8Bc0QuyUA9edJ+sdecw2tyibbdSrW3Ipn6lSvXPUHH8eRYZTvi9nzZ1icsWO63Eg
XbV2cWsE/RFcBrkHy6RNd298X5/7Io5KkBYhKg9RdQj5wxPiBLX9a2+qEFxjCFlk
AznC6PUrLh7icL35YdSwbpMiuOUO7ZEIWHS8sRUNYY5Wj9VvemRGnZUSHLzOKZI7
onwT+jYZMRnEerQwdX7LPbINP7PHvgu131LJ3BqtMYqG65Ix6I7Mp6l3uRXSdOqZ
EwcXfy56cDj5Dev9xONTej1YdQCFRPlBYTD8KDfqGM8VozpEFm7mkPWKTHDaGG4F
p1MLkfjIWQMFZj1mSwzwjY358xb00+OXHyxK3uuZhaFnWvwuwVxwuANAxA2HZnLp
kbq33LeHDAPl3pRQEWFji2kOtvpPA6jUkVNMP8GFRkg3D8nBJi5OTBigecWQMlyz
x6GCvkP3xmuumdsTGMgbzl5vy5UCqHNabmIORHbwgVDi2snRK2foIa7+xlpEQadL
c6LIQ80Z2vQJvDVGFWquNSWMuR7B0BEUTTH5yopRxjEm3fvYimMegTI1yY3Swjid
/lzdOGj1DCHOg/ganiPisP6ojeYwmW2GF8vauYBmpfDmi/V/1ihmwQ4MD/qef/75
PAh57BKzz3exBYlsz9AKpG/30erKDFR1lvto11J4hRrkKWrrbL39WtOiVRA2VvdT
d25EK8IiIzj1BNdUg0cckELM/il5FRaKyicT13vzcTmYglyh1AYvusfpr8j5w+Sf
CLMK632FozJs8ar+ApxqjWVl8nU7lwgMJ3UXitML2USYKGBTSKMGnUHd/N5LNTYr
d4Kr0UfebnNlqEW8WzWY27uvrEZxt7gvf0mXL2FfMfigWsktTRkZFD/7kXJMG+iD
r54bJmmnMq+nInUBkdKREvW2VLTHotpxhX+fYU8SxVX3lxfqeVyuyXFSJgQLq1LP
c5n4hxc17XkIRQ7GR3evQUgG4TmdCrRccZQvTeVAx/SIwOjhm4X9vN/Uoh+AfHYF
ocwBidC8fTjCiivBPknsCbV4IXJc4iMWQ6px+EJMLNgJd6ki9oS/r+4Ih9fygF2T
8c2xyzm+oeSC1MIAs9mi+MHQFoCHSITrEnUa5TSPmmvGX6vAQrApbecTAhpeP8Hq
+g839VLnuCh/f0R0BbbMpYXO8PqYNayoXuStsGR7X0INtSYtsGnqQ1gmGPMZELIn
D2G+AI6I8tJe6yXKmx+BJ55iD0MaDkR8vQPVoZ4h3gwef5ZatAj/vHaHNbODjkcJ
yRa5BEz+fNilNlvx7Kdms1UV5NPsnSHkcI2tyeftxvpgLsgV9V3sZJbn31CM1+BK
hC00y1kH1eLmoAREChn5yO84SyBrL6t6v3EBQZgKgaRRnRPaonOU9jtqfOyhu3vX
3T7mMwbKe0k8feXJSarcSZ83Oh7SgaFgGzbTtg0Q85hYjz7Y7ElmbNVrbtybYpGH
pJlSAed6qM6FvvnQz/FEfjkqn6XOzC7+NegEvDds4FAOSsov5AQuabdikrBRsfay
Fc1PGPqVGz3y+NlHKtBCnLDOKi+jGAfDctA6wYyukqEtKkTtfA/0FonAHaoKP9oU
n4b0KdYWI7P58qXBh8TJiNGbuQQBZffetl7lAok8JkjSNloft7yW3ZnCWtaVCnUb
orMNPAIzz6GLh/2i89L4MA4SoB2QenYUtq6ArB6pY/M/sIg8OOXkXmF8jwcsXROi
9M8JOGqTBH4pY+ltOkCEWeONYPVMgK+8IjQmo0CgQPCL7a26lzycb22LxeQhZhXo
WZrOsv6hXwS152yXc3VPVrJ65EZ5kE8OtOIOaxfEKMtrhrdpOkpJatzZJsmgPvAU
MHvzBPGokRPLOh1YshyEFPA8aZspy7UH+yTr0aZkhOtZEq6IvlMSPt5DEZwwxB4f
JU121KImpF0b+GJlbkgorckZaO502jyNGFunNaf0BvQ=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
YkWZey2frCOWm5CGb5KbImN89mp1Xu7tNGNkCXPq9XiGwFGpA/CCvz58cxs1ZDZ5
7JEwn1oMhOAD7l8C6ZECkGhjVU347Q8j6mRtVu6XIItRyEGtW5RWDPbqW6uPrV65
wZG0Tm0QX/C2/zUT3XkwGkHk+pbD3WlrFdfm6hmTWg2/aSJ+T8WPCpvok6BBKC4V
YKgCAwXC2Ou06qkL6wrXLFbHlRVQmzUMS5N/BuM1icmWeg/b3sHOunxxdeH1nTnP
r27NvzEF7+kfToh1nfJEBxg1Jh83t7MIQlxdQqDb9iw2FPjQeKluPNxB37xj8eXH
TLx4neNOKXgiK/36Lwfe7A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8928 )
`pragma protect data_block
rm9Rne9olKEPmERjbq3mFjt0vF3IH2pYgYMyry8EbiJZ9ZDX2Ad+wfgh5bNaaEBm
QiPeIe+YFfh5PTHsFkqpegWhJ2CljII3dIzHuCuuknr8PC2O8btfeFRbt5hBKOxe
FId/aptTrK1pU9G5klAnpdYWVwiAzMYlomhgFjgNJWt5jq7Qx6BbpafGKYUMj2mQ
JkTArtybwtSZdAPWmYJha+xwAzEiuNdUuzC27TQ/Bz/DwQX1WvqIQbmbm7FPiuIT
BfdwZ/DlNSNjukg2aZ6BIBwo6k7ySbhLVbLptkf8ZOBzp9sx/jYIhdlxGgosAAQ4
LirX4SXcfCaN9ulTrWgiX7/UQ4EDLMMQyaBOB4j9n5IXYXoa6HiBlAS1uP87fqxK
+zJPipEIvLJPHNQV0STkF775WOUiL0Wi7DF4U2SR7ywpLgLZYsL2FtsHE85RXClo
y+OU1R/+ve8Bb2Jf3E4EECucJ8iiju6kjgrHZ/JLjYoJmdLYBCcdRQEgYAE/FVsh
D/bXf9oKDrPsdCtvqmdQry9wvWTh6E0p9544aJo7ZPAblWOITw8vTUuoxGiexEuX
E+YHSQRdX3QQeminPkyCEKYQUQgRLHWRYOzlPj9C9Gr+tRJpX/uVdUXy6Gw/zO4s
0diQOs/d1pX9/V4Sl9ohFGWypyoCK4yJY+G0buxxPurm4++84B+Wyu14K9+7mbMx
heraRbLAPz7ovohQdHkTJ9QkVa3Z8ObymxlJaEfCL4my83wSdEEiFgEmgooLWhx4
3i/sLAMXILXIww2iekSsEfnpRzvUnh5MF3dKvzKTXOGQlkHAFjkLcE27Ol0YIgHa
feVv65Hf1BydTkA1LCYKuiHiJqSpOBFFaGnj/CXLQZeK+XQu77y5zseEqW10kM1W
hHc1QXFTUFG3OBj0oTXwZXngkiNbC1jZmSTplgi1q+oR/AHas+mP+YiMyPCDNUFM
YbcW3FDM7cV8uT6PVmtQUiXn1gb7opqNcsE3Lo3Byhc9vXlcLBZWznAIZJOKknWJ
KPmj7y0XlVbkW/WeaK522MEmtfjGFa/MEA7gkQHfmDJcnkjAH2m0iCT4tiwK8Jap
hGtGJBsyNJ+k4YlQ212uGYv4zjT7GUO1BXoDBqTYrfYSM3OPOnOosH7FdnEZqrdl
OJuuxhQUDq1SXqj5gDD+A4R4AzlJ03swvMegzA5IH8f323p01hIgHzkr2q9XWAT+
kwe7dSSv8vVgXtMi6BIgaMpi0K06hE31nl4aeGYCfhxsCdlLh6Ud6cAdPGUE1I/K
OHJBwPwvGrv/sy8OxWx8GTGztQ2pI2Se3q5oYX9gyY4k8tOuthq/okZMbLiUkSN9
oPh1gQzEkjOwa4a68I1/AySdSi31+tDF3V++B1qWGNO7EcR2jKgC2iJMaXtzp+Pe
3UgBD9v6b2/00gHFYPPEyYTrb/izqyx44m0haprdS/xvblYehXnMNyq+cVy+Odld
249R8QdGYobZ7fOWXDfnSu+2/5iq5WgAsVjf+dIUQ5Orhp85bSt15/sa6fenK6rK
cy/wVOCVoYqk/Nfk86OtD2e/odBmZ3JCka0IXdRYHJ9j4KUy4KU/95Mycw7N/2cF
7fhhbiaI9V0YmdUEwxCVJYd6a5oe68SA+GQaBGk3kVRjCQMdbrUgk+Vi9rEyfUxF
flJYQFpv0oRgIF6erk27SpV7U1dStmFn5DTyiEbGyUOS2f+UiH/Xj9YyyTGJDJwl
P4vdtGi6KTpw/Va1eGEO3GxaX0Mo6rEvKoQnj4+Kcsbi8mDUMHezBWB6B8MYjQSn
zbanJrd+FnBYSDfzF2bLa7xqbvGL4ZujO3AeLEbGvcggH+P2G+AvAkq2hf+rw1eQ
rl4NDXVNqUK1psJ4cvGWIHEFZ6i4TiTb9MrplACI4xE7M94iyNylh1KcMYXmFKaa
PGH9z+XSz48LColztJcpmAMWPT0MOO61r7H228SQlah9CUUXDNlB318LaeEwB0jZ
pJrjyhygwWa/iKT58jONclmWUnh/aJ+H4RaWPJfus6AJxdcg4LE3CPR6jBUcAXc+
Jqa24cwhTD0dBCzHK90RSs2RriD3dkDf0L3qrm4502wvjI6TOqzc2bC448BDF93d
2jW2R3ePGqZr+WOYHaDcBQ/G0yDhnhAaZDqVIfKUV1+cdY6sfqxbqmo+yiNRVeDf
L83sskSLFF91Sm2FCpPtvaVBdMNxmtNr/4hsKHov0+I1jeqOZSPZKCZLXop/AWD0
nqTeYBWlIAGFbYzkjnFQA1n3LPbO55PSBYyUVer+rt4BNTygaZufNTICyCScuIbx
5jL8nU/0oQuY6lB8cb1spwLCCuU0Yq5ZkFveUQkG2bvuVl/aOVFTiN2I2SprT8i1
HmvUwgXmprkvkQ+hOsnMHqiPWD3XOKRnRbxrKQgTr8reMCVMIQNkmbSqE37b9xrN
piWJGjuIZ55riH0oWyNc2ngl6GNKRG9Z+NI6vhWPAB33C4ZseVpfTqC7ct6HIR3e
8efB4HsB8V02d0tGSVx40uUa6Aj3Wk2+WfUEJzLsEZE73QJxlcygiZX2tTEhNuGl
5laV1C6/IKZY+cHkJB1GA2MU9BzBrpRlQfmQ9RE9Oo1qmHVgk5k984luuPe/YGSs
tuJsvDG2G8M4Ewuo3Zli8VW/Bxi7yfAojAMuYqFu4SzC+xW3HeDaz2JGZDALgeca
eKiImdvpaSlDDqrd9Ylm6Nno1vpAn8I2usf057JVHFg/to+bSo/VfWpbYyjlHsVI
qLxUEwZbty+Bc97joschrTLA6IVpy9fozYAuy4ypCjxBGWGZS/YwcJ/9V4fjriiu
4BviZkM76tItW1ykOCLnXkPk+2dONEXAqkNT9RDMiv2DcsH6SK3SA0puZQFKV5/3
Gxe6ELle+1QFGoYIPyFi2ttIeu/Rk0UibdTIrI6aa49NYEMLe+F7PbEXyEcanTtK
Ld7/fu+d3DeRNz3tkYEqeMMkGVNWY0WqbpB3eEwkwpiLurwMPiZNA3VWpZi/FhIV
p1PrUv483q7EpwUe4H0gwIkHKHkRHggTfrY4M+p04MMEA+/bNvSd8yLjN3yqGP3r
mWfQoiJ3AIUN82aFDSdBv8nfm7Xzk4d/g2sPJ9v4pPjcrAZnwq2nYtkJnwHCDXOi
nczwemt73OIw0SwLLkL1pgYc8nRST1Dt4JLDu5iw+Z31SPH/47GrTAxHnU7uB4ZG
bKkpYgWcMMOK6Tvifz8Y/WMpyraCMlivrw0swbxPfQm0NYttgmgEhpN4ZiQU7o0c
Hax+vU83i6FxknvkcJ7B5zEqNZBn24Mc8Z5vtrq4if5jnQ3TNzwdzTypypOsBCV0
l4+ztbUw5OKuTZFuB1gtG1upKLUE7Evh0mNWqpwTr01CHTNPEy0aRSmQDs+HM7zK
zkYmK2KXMBLKXI+gVWVVm7nkqGX6ACLBDHxBzDbfYdzktJk0xMy3ejpfEikFhKCx
JISj9KRb6iuv9KV1HXC3VRYMiRthl4kIhWdJLkUAecWoQfUAKh4xsJkFbviSmEY/
AkEggiVG/wT5UZb3GF/gO5+0OVJibCT26ggVzJ2NndgYw7O0r2Gno4REVdQe+3aw
OZKGt/geGELveRFsDw9zvXZcFNPSkTwLg3Yaafv2fu3p3q/eHd61fv2HgaBWedl4
uzff/YaW1zO8PcL7WcGd3tVTuhXhmh+8tipoBQOj9OQK0azZjysYznvxfDvyNXUp
zWfS4JVaLvcyuCer9L6y5xXOYtNDl4t9rSDJVnZpkt99fIM7Tm6Nr1FlN3RzpQoG
bXHCRsJ1AjA00mpFAl0XcbORKsQAPmOMJpLTAmoCVDewakPTkOdYmL3WAFVByCnA
oMdPYRQXgslAeIOIhPwUViMz0tZnGGZqAGSVXvwq0JxYnZmsV8cH3HMSogAeIm7m
MUT7WnNPR99wsK2wgWHOTusLv4TTu43ISRuV7VhNccZCy6LzRSyQ7ZtBaqzkwpub
JACibDjx7z7stESbqhg3rSnuG/YacAuBx4wTno0F51KbhMV2tP4ts8VKDbQ2j2vX
l3dnmgPBh//yuXkKyEHEcWrdHQT48dQcZwqZK33rrBYwypbn5xYEHPcjE2ovESyc
tPCBtdUAW0YySBXYveyZmKmj2BfaIGUPuQCrc84QYmiy1Hy+NwUF05SCf7aBjzs2
LWQtSO0xto5m/pv5H0H6vn1HXM4BWaCNIuAHFmILLTTDs07VQj3JK0cB3//r5rLX
in3TgHsSEex82oTqXbgd04dd17Wob71oTZ6wl1tYB5j06h1H0OIhr1nTMIH9VToi
oUBOMSIPT4GAuICoiIf8+Lnt3tB7SrdA8opBwfMCKKpF764Ki/xAN2NWmGQGflz1
JJ4zju0IRJcGR23xqAtL7lPKZ1+jVFCTv1eRU+3cXnOVg56gueeliGMZGnDO6Rl5
6E73iSmH9l18PPq3hmHpYSSJRiHmNBvEg+TNFkoov1tVWog0dID0b0G4p46YrZbK
lMR0RT8uhskv+S0nekq9ZkIKd90uzJvTwYNIbyvezy2LVtiyPtyrZU/LzDapLdRV
j3WEV+ac7BPOb11wNk3F82sasuZslrcQ8fAVBc+wUiSUT/mKtKlqoboxynrAGn/D
emw6ytTvDpN62xOOWC08C+My2PvcTkBQuy5Q9BiONLL8EKl24fl6+0wVC1t2WL/O
hnuhdTOvzM2Xl1nTm/PIsMtKYjTHg7k63+eBXlT7TUjtwue19aNrLSwtqH2RukfQ
18rPSMbTyg09osC5odroz1oAM9NKvAKLyFkAObEw7xZNdyqEXTlOmRhvgYX4QL3v
usjr6epV5DtlxhfVsscfJyxO8rmHreQW4QMSH+UR7b458habvw2qMLUpJo7lpXXB
PajzefueUlFhfS2mOz7JPr/LsG6ForOrh56ZYI5tpS+ieFWrbziBJliAkxV4u6cY
PQwSVRL/kQjUjECIOBwKwNYXIRjVPj2Fh7F/5WToEhKJ4xlTTzq8N27HV8uwyEVg
UZEKnZYRVD3qh49/zWuExLbnLqhXmAAPoLniryxpkXpJ6JWCxXx/zCmMljdEeD8A
wJwM6nRcwKncb339K2wxSB7Bi2YdJXPNWiDAPTpuzJpemiydPX04jLm0qr3Dw5zM
2E8zX86rRueEztvl2KQXJGtj+XwFM7cZ24rurncikqMhf3MFBbMqRgRauHiB4NEF
atAK12AR7UMTgHwTqorLrfvZIICuUDV5sRWH8mOEKk4fZgh9Tdrrg/UYemzTOVcs
J9V6wBqT7U0GK9FNhdvYziaOw5v77ZTZcbiWwPF6viouSv0rHMpJn5FSAftUtB2M
MLMWduH63FDzr4fFgtgKfzQIuIeoGMnXXv/LYlQhvkbEZFYv94LCigxK4fvLs/FK
ugMOYBBJeeEh4UigHqvFdlAElMOAVA0EBGEPyaFu1fOaPZCvt0/lRDeGSoiJVSEG
vUImbLV/qWUzVcDfI2MwUjzB4yNQoFRJazz6MN/FFVeYOperB/1NWCRLwB8eX81w
L+NZpHwpMrvlSiG8QNQXOLqCpWJihIdGoWqChqkY5tn2pbpuI61ZG0Ln7Y+XilT7
P/438QxJeXW/ngMisYkqoWx5TSxHHmoSv4RBckdzk1TfvlepYEIed1rNvm0+BWD+
u2wBe5vlL+M4Fv6P+XKTt5pJJ2Qn0CFP8QcGUAW9wN45UevUaMnVPFlWK+aqj8QW
yDTalqZic+y47BXvgmteVrZGjXoYiJbpB1rW1trbRWwQCQimNHy2RvV68Ve83DQE
qHDGpDmj6ohu2pJOJMuc9Wbu0FZHJt2nkmT9HxoN3+96bcnyQLAaGvTrLjGOkjG4
6t8ZOvej2nhywOzFvLYzqO5clXE1feR9WUX8pEhEt+y9i9XFasPH3zekBjtze5cX
8nDpNfavF9QzPLsC04tzIjph2mlC7Tp4UwyytsQHJbg0K3dkSNsBWhJqkNJ9HIDb
p4gdeQv48XdArhDki5SNFCdwOuA74xx+kP2I/tl69O7kYc9IL9UHoPwSg/TA0WPs
pbraknd3lJ2LhbDmWtF/pH2Lt95Es6WeNy7YUai8MfcNue/7OUpmlEOOXtJlBgJJ
k1k51uDCtgyNDTp8rnjn3ZJx7HH+WPVR1YfHYqPo2D5S0Y6HYypdJzFsniR3NpEd
n+9xlIywVOFE8zxICkWx0AqUsr+XyLvbVpo3WSiZgsHBwO+jK3VV+aRNylwBIiaN
9p9U5iv4yrAQgSGaZVaZFMdoS+EgSDP3D8MRyM7gNpVIC9Nqx9gBBCDEzxuuvfef
XpUuNvJwallTqmd43GMnWG71ZUeHkPrkRVzikIZjRNsujUr0opSuCk51WVvp79pf
/uChssC5cMEqWoHYgE5k2wlPEept/fNlz1C4ZGnuCU1P/AJlfInRMcrneNA3av00
IkbEH1X3QW+4+xs4nm8wPC+Sydv5erf/l7Z64dyWSso7LCnB1mGtYg+NxrxE07we
YfvN7ElasjsUmdG0FlkSSltIPUk1kUmfkqOMHgI8R8/lwGLMoizqryMx5QQacU1T
eNiWw+WkxUWlqrvXSl6NL472UCFFdf1ZBzWe+4eFcYU1V3n8TFuOuRCUC2vfqw1y
GZMiu+yvVqMJdS8m4dcYlySu8ILu6PUM2AuYTbl2du/Z7lqVh26FwwzBpogJ8k8Z
FYLaByJFVtR5wWLj2EbKnHatOn1N0S3YzK1x7Wdx5i98PjQU6aZ2qW9mSXtHu6vm
b/qfQMXnQVRZpTsWNsEFKDKbJcIF+W/pytwysRwsyTPa1F7YYmObyVzzqYwk5uoS
GQOOXEFG2FW6rkp5lTRy0w06hLJNYnDOA4Qnomuc3eSI5RZP1U1L2BgjZ7uVIX/3
itM0h30xiabhPu3MQXwDm9qPbykej5MMTL1rPaAuXL+YWsD3o0n753Bl2xhWyNA9
Xb+qeb3SR0WPAV3HLVvjpGWVpl0vaQiv0tsKk8sj5ycHCjIprr4mpvcnxnVS40AO
F6taCrejBlqXV+evhxa1PuWKSwSW71DwIShYa2r9kcbDaeg0pX/nQ86Vno2HgkRG
+pZ8otPyxM6dAbHKs6/QW+vpXMI/EHwEciiwuzOb7KdfOCMeLCumPPNf6bJRSPop
WNSFZi3AiiFO1wPivURVl6hRzu59K/n2J9RZFHM56XuI7t1KAWTnQGpfhZVOC/mf
V4R+76VQd5SL9CPlefcuNGdKJ66ffw+xES6u9feB6+otOmYcMK8dHgE/rU/hBkX/
05zUwB73CyDhfm360eI8WivroqzKJBEctB2sLUZ9SY85nf3acfyQUc6iqxdGWVdi
oYUGIMVDwt4Sq+0QMNSMemKnUZEL7JjF2qibqaV4vPqLE/Xg2d7HcA0+MUI17DCB
/9venu5HYqA9lKDLVduhDgv2rWfQ+ELRk6dJlk7n4tLi72k+ZCT/OlUFpDq7WzNZ
I+EWLFYca37v+Or3c9iX1A48jEk7QDpyHB3V7XhcZ5068HG265i7wAr27rumFNa2
T+cb9lIjGQwuHocn5rTnTp33iqLGsGvU4hJjVInHM7p04xiIVHC58EzrVXE+E/0u
a3kvEshc2p/Fd2Gqx9tmX9aoNOrlDHJgrlUV+l/PZeIkRjkdZbXxIm0iZA1L9SIS
2rsGauM8wsOi0+XiF7fILrHqUs1tyRZZGKj0YtPY+KeqvlFJs8348+Z9z0W+bVph
N6R1WXLNVr4nIpVVzdMz/IMjUZRQYoHiEGEc5Px0dCPCRnjstC8CHvesMEpjf0Ty
B4vbshrYOBssW5gvWg+Yy0sQiUfrV+cOCpuYCxCugiKrQJqk3+LL4pnreNb3i1VO
UCZ6QN+1tC0b9/5QPWc8HDiZn0ABEDBLSPVvIrPuWBTETF+bEj5nF/jU7zH7Dbhx
+Cl4/MUu3Bq+8vqJ+Mpr+qHfyu+qpOnucZQmksRKvnrmb6ScYwVcbo9bUrE+Y56B
NWsktHsIk0bPfa6ZadiDT/yAakeXEq3mj2mcHdx0HLNHFAkrWIZXwAMmISXqzKM0
jp6LB+iGE0I2I+QvRiPaxTU+6MmoCvG638MvVEZjTzWkueFtT5kejBaE2XxggBnk
OrX4uQMJHHnhpdW7YuVRsIZC4Nm7uiAUHyIereF61immuzRZ2ect0SjuUQJq3FhZ
Hq9pOLDuDjudqUo8yDclzDDOFLrei2NhupWN+URgge+zWnYfQlRnIjhAJ1+HXpHu
K2P/ZbHv1TvVtpIsjd6DCalS9YUfSA80XYq1liTIBT/JQlcERPX39h57nfJDqe4a
5vyipn+Lu57VyNgjhzBPhWY1mXqm9XtWJiKEeQ6oTidvigl60J1t67dFsfgHhI+c
2Hxj1PpCUQEMTBMoS76zsuMC9P9Ri7lT53oFHSNqetBe9zA1sjUu+SLUL28i8xbs
QY43fitPtZAttK3dFJTZqfjxlphY9cR4VkWXQUTFEO1cqwJsLSCuedLOmNzP1B6z
IKCEs7irQYsTiPsaOoyNMyge/LtBq0D6POj4bneRvr6zoepvDqgRBAGytub0KUyz
yYkq3WPaj28DnZhT0+IpsxtiCZcpUFg8PIVq/q2C98KRjWKAWFnRkeZefRJxU6iu
99bHQT/9RkLpjTAiVoj06gMSxzB26E3RfiF/uvgfDtGxMgJe7f+kkRpTT1CailBi
Nsj5F/MDFCZxY6pNoHBhi+qy42pu2IaawO3UtNujtiJK9xm9b7b18UAU2/wDfT0B
Lwv4jRByKE9KHjV5YCnTPBreLqdW6aa9D1HFSWdGES0jJx/mJvtUlEDzrqzPfdTl
8eraxyE6J1oLi/IoeQ3cMiGWhe+BddKKyhk2NF82KvX+6cLpbIh8rmBsveAMlg8Y
Tm8NvqqWjHFl43UcbXrhMVZs+LoCJrUQIoTaNh4PuqsTXZBqrqUyceMPEOLhnXrF
H79rpD3DqSQpXE+7DPP1qL2nBYcsYjTwawbgIymP6G1YsMxWXPZbeEiISLQzPxK2
X8KSkdwVyIK++lryd5T9Sg9MxO6+ZUZn5R1epERJ4NwOzI3J4VMhzjZxGB2SgOI2
iayBA7CG/250IdaW3lUriLYfOkhRcG+WFqqT5TVly6MBp90vfzIdC0rsED0JVfI+
q6IkQxtl8IW8htnRoYEHa1Gpo3ZOv9h9BCViyoOpQtv2EX0b/erAlFXOkY6GfhBQ
9+msKFjXZ2EnN0n2P8QgzBPXYi/b/FHNWWchs6Ov5R1jSuqLrXlzBQ/cf97oELkQ
3sGpkx3k835O8EuSXdFJzW3kjMzqYr0lPPCua6+JYUrneNDSmTi0qC4X7ra0z6/C
T+qxthLY8F9+cxp6LroH/8WknYgc7q4VP4K92CJzr2oFRoKv20R/AgJpvdZTyZOS
l9fa54/nvaXvjMnbaoI6ZtQVQXoFwYlrc2bJw4oaO5k3Iu9xy69QlU67x/cACMCa
NrmPSLYZ8xlWREBEdhHoFCEPXsBkY/w0nVTHnsyG1NHnBdt4qNGWzTP0haLw5sG3
3qed6kjDIdLQbxV5cEAx8oMuWhoNKivi/S2aMatBlww2Z0Mu3jxzHwde9N6vJsRG
j0FosKxc5K+vAU+R/nlbW1ewLogt4v929QhscGeeL0YocCl1ds5yKa1jd7XU/MHg
VzHFWKuPZIybW13mvPi7UQGDO9Qsn/5adQWcoxHysur+Nxn3VEZO6FjTfML5q7Fn
nf0J4SKYOHEcezRTiXMNWt1PcO1FACBZpZf61eNECPDJtQPXn7UHn8ilQHq8yhja
H4PqBBSLK86KQlDl50cbjUoqm+KhYepvRwgoI0rrkSR3AMQW2QUeGcZTjc6HyGOL
J5aDONLNOQbExthCPGAhWcUwNUGc+q2d2DI+xGbg60qZS7i6//6guB9WElZHS70Q
kjYH+SiiScUTlklHn/C7rixHh7HPRKrKQWq84YxD7EIOMWKQRyI9ugc6Gr928INa
buZH5t5lDiQ9pSTMZAxzBzpcv2s0f8gBMe5X31NGyF5urELsLpOzNxcRlugKZyvd
a7erLmHuSZWWRL5I3S//BHlJLpjzPLtHnKwiz0kSB/LBoL8976ZK/7HFUEgUGbdO
iuVGZzoo6GQZ0d0dfkhK6hKj9FAyVD1eJoP7IrHQDPWq/XPSKGr2XOiXrJ4STZYf
YMdyPsB0/2poNyPAI8Xqj8lnYJCLhFjiIJ3Xf9f0oyxmUcMoqNNUwBYsrmGN+Pbc
aQd4eCZcZGiMW0/eWveTW7wJuzMugACqJpm3CyRPW8pe6CRbrDXDz9uOJfbyJmU9
yuAkbBk+nOtDEmSiwwTFQNirZOIAYea4v7snxHB/eCc7eUyGMqh54oV4ER8wf+ru
ENMw41QMA8/qH0yY0Za57q1eAZbVWYoJ3c3LQl87Oid2OzLxdtUfz6SVfSbKiESS
nL8QloackKNAPfZZIqM7k0t8/YvNNjAwPGOqxXZlA6K+JyhXt7sXAO+0Y6fAYRX6
yEX9R9Q+qiKrjzXzkElwYmwLMPVDEOJ888CRaEuNxPUPex9fVCn8blCKpe26ZmOQ
xxxqLH+JSJmXwl1evSEYZvpBrcZGnOyt0PJRRdvICy1rCUrGR61JnZulWZbTYyhU
dz9QXsJpP7N0IKpL8TP+RZAnvNiZyxBFkFEB7hyFQK4bh94f0vX5A5MtFwPbBXtj
lLFLlwdg37db4RB2k/fcGBhESnM88P1bZQaUshaumRaZyc+C+Z+9ARUsFHu0f7Sq
ktu3+046Zfu9ZulBslux9JZL73OtuNq/M2EKMbP1TjUSTALs5zi9PMNsbmXqWtj3
2jpMl3J3W9J8uXsArSNSa4uo4KmyxhUGK34aT4o19Xac6G3lzvhY8JAuYLqwnesc
txPw6jcHm608GpM140NZSHiwSCssP2BDN/ONsVBYGhHlfvxMcyqLWlE/Ix0rZ57I
Oj5YFo18U8DAwCyBRDgkXXVuqFgWMgliiPuil0AZl1iFIweXBQyRj09T3CvuhWXi
eoc2O2UxrZ1JjSRZMebauMqP2PM+CJuRi7XpuV2N3lXvE/2xveOoonKoP5Tp1Jsq
Pzy3Kr/Gzh4pvAwSMbnEifT3nPJYMFsmORRhb02TkrgwhYs1NcTvlnAKzXrZrWBk
7V7oHuZESWCtDEegVBAIUlilMLVscyOqNcPhbykiM10C+R3m7WJjHV7SMO1ulSqx
g0K81rwzUyRHcQm5E0x+eg6aJRmMdZX/3/dkoRXonbRmSKsDWa/8oWlKsYNuyi/n
z3F/BWL2BKdGC38OLv9hjHgI+2vD2HPUcrtU5YNADEH2zd9ghVqafR4fnr8jNY8t
qymlgAOoDJ1YVSwxPvFrURL8iLAcAuq3+wIrDc2zZq3gIr1mxvi9Vvu/+i9Tj/1L
H+/VY0Zzob6SpGoUKDFFgXvNGX/m7VfHpXENcsTUBktZvp0//ot8Ynlpy8ELu+Wj
gUecw1zhFooYDJn2UWvgXotFkbNiQLQljoP9CsS3F2jVrNCA7K/ZW9fNqegBR1Q/
HoM2R4/+NWGEz+9802svC3j+dYwyKCYbVkri7p2ZwiaQw2iGPmaf7nHS6rQnRnRT
yI4LFKXkAsVgNuDerTJyqG2UpTDovbgz1ubymvEL/k+n+vkPVJ3SPgO20cQMBeie
MfQov4D9DHfj1fjf4MFQsNoQaaUfALGQWc42jdNhWe+9C2D5Y7FyeepeeZW5deqy
6OLwqkAfRxaqc0VbVcHZwdHdVy/03jvS+cPVyvnzw3rBy4SU2KGkl8QolC07bOGI
yodSOnEV+jwpph396iZPldJY9Bsy8ovQByF40Tqb+ust5i3G1Svxg1onHj0LJVEJ
UMnbly7FvFVu+3wZy+/PRAuB3N5jiqkW9fMpoSnJODsxUaKnhihVXcIpHAyvzZAW
b9TL1dB37K16bZpZ6TqXU30zepLvEl6u6yvdQPYn0el3yPuyw+sWxTUnv6xjrq5h
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SOyjLihHpKE01z1/P3mqPnBgyoQflWqKPVj/2NbWQQvStmMw/nZXzPGuUf04kcef
F7O7FHV/+ohU0YRP2QA20qHuKXrRsKwAEqCh0OKxx/G8iFXTL72Ok2ESxpiYLfO6
rekK1hWKY0vszms2O2oGbW0OK9lC5iy3CkocBoFPbFsR9eZ68QNYvAHFP5fNI7iW
1G2L7TIapU+W7eX58Z22BrkaRmjGdDwqXqz+Gjg2A4FIy8LxcAiAzSm5Rw6SGdvC
NORZR7C7KawEwYoEeDyHMTEiJeVh3Znw4U1i9hxYi5gXmip2eYw0lBckUvZinXO7
nW/N0yJ+U9xs0MBfwzIuVA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2912 )
`pragma protect data_block
TW4OdrilzdjASJ8svMM8T0HhGkmGlRNilLRN9l5kF1H/irEPWDm5TNOLggM6nH9o
zR8gtrbkMgrlmRRfjvQMypG0Se632+lidK33ZlMrzfikHDooFZ1jP7xymjQYHRnz
DBzi1eC5tspe3aLZuDbgo8m9rcDBVSc6hRloc0Em2FY6S/vxTDZfP90XmPKmJ9kr
nh4PYg8n1DT1VdttK4aq9u1MxxuLMMOChaqQVnXrTbPE+9kOUV6mCKnfsvhugXWN
aEadfW4wsZDMHeW1PI0gxk6FTpENLckK1dmE6M4vhb3Lkstm/RdCUSze5pZKw5qK
9bFIwHFhwF6NVgm/24EKKK3VvV+5qFui/k7ODk6AgobejodNYk0ItV981zjB6E/J
rLExzc4CDW8K5rLJ35+tbkw1f4pwxvUDtho+YMtOkQM0kvMrxZd83GEnf74L/6YI
dmHhLDB1O2r6Vl2wp4coJg6R/MmXPtwG6scA4Tej3970QVsBZOgKZQndekI43eng
2y9Sd2PstBlKgR9VeEeaEkl2E2CC89AXDeqvXn6xFqIUP9Ddgc51jw4tF74c7Zc9
Gf7YOURg/wcLSzk3zZLFK5X5o/pzGNw8R7IYfpZUVHrTtKS/qo34guy6J9h5z0aG
AxsqbY0ue82m+qFy83Yu5xqN3A44bLPAEdb113n8Zxc3b9sWIBSLy13H1v1xFkR4
mmMeTzNQWPpqq8qRM+Z5HPh1qxPu1SQzSdvOWL77aS2MtbjGiU+HSmHeuSpgYTcU
0Aib+Klv6iR11ZbF7sy5hjlWjhd/njbYC0TKBet+VCZv1SuiYe8z2ujnU6Q9+Zmh
Hu/N6nOf2HBhhDKzFld5pbyl+DyIj5956BxB2aBOSBSeIE+ItwZZbVc6Rd+JS9ct
x9mDH6YcmJ6NpeCvqdMc7JPiNrcpfojwZHiqytQ908J70r58znR5znT7wpcj/vwZ
SzBWr56d+5KmkEZBKemwBJcMy33Tnj6TQ2vUL1NqapXQHZaOfNkz0+UqxUU2lzEM
f/lSf6/hoQ4kGX0Iv90iFdR0Tf64/M7pJ1FRBb64ItJKuDdDKPCbFASP2YAQ7hlV
/TuojV+oPXPK9XqW6yIOAbLApp7BLtwP5rtrODxTyGKredHpmPlJysCNqbVvMDAn
PVYLuevCvRXsFTYXLoZk11yj2kIxws24Hiib3zmutVLDqUtLxZmAoRybdiaJzX4O
rwGh0w2CR1r73tG5wwwzIWmD+cQDmFFKZZ48XumgDilaPL0T5h/U7xN0az+wyZPS
a3rGypCVzLAYJs9zB000IYuAFP6Livz0or3zczxfRTIvrzNYZw1J6z4LCZ4vV16P
/U0fivWvo1PgN4/Su5mLck9gVYjfSaMKnnf2ZrlJYbeNg7q+uW/B4z2aTvfIFDQT
zh+ECcLsbxV9O7G7hX3oU4eFvtGVEyRa7/gzNo9yLiYjOQ8iRy6mpKMF+Qv1DXQq
hh5/2E6hJ86IplyoQjj3+fhkCoK3jysG01ARAFjtgQBUUUoqR1OgSBfLMzKZ/rU6
YIKofcJ0sFmTjc0YhKjqpK/Ln5j/oXdqv9+oTH+X65VnZlDeUCi53f5ZCPGu8Aha
UcPUZJMifu0zQQ4lNhmR0bbHK/xhxGRqEea4/CLRBc2LtdlmXGyLxwOny2j0djEf
ZLMX+uAe0GBclA1uSoyqC85heI+II7xQW/Pbg+G8vj4AMeXHU5AjrdDK3DE9UhTq
APg0+sM9F5AywE52SDqc5Du4hwhgmxr0yPFCk0iApC+vqCmOZ2M5dAKfsdc83Kh6
23wUIW9mX+EfsiWTvXB3fF/7Nl+gBMZffT1ej0XilRRjK+aovIHv0ATtIgKGQ/fW
jl5+B3XvcKqBJTy+CYYapcBeyjXg+alszxRc5o/QhVraNg36pvaybM4eB0l1To4S
ep1MaoMvo9rh6L6H2DqwTQMClBF2xE+h1sp5ad5zBWf/9wPt0wFUdnFE2rK1GpSQ
Dp899X/4ShtRHEWMXSZpZ1amx9TPthdlXzPZo7X1XRFVtHqsSj9Gh0iCGaAYDt2+
tmGotFsUR+3jzdSlpEbTV5CeVJ6XdAKgCkWDOtHtRfKX+EC1aJQrYwRejyVVFBb+
u2mfx4YxGgBECH55ngzFzFQLZjtKRddAVWcbcST8A0Vp67Dd7PqHiyGD2/6V7Qql
34pJ9V8r23JgSU130XabmkRWsevnHo+Q8Io2R9R9vEiL6hZFufBW7f9voF+XmwAv
a9DBOrboZeMmkvGOveAW9J+LN1YiPFGVGMpzN4eZ88pUKN0vadXVIgbTWVWBtr+Z
4KefZXCUHAWYZ+0BrHRxMqyYNgt0frJDZY79RefrI14og1G6mW/YlACS4x2rZTeW
j+FZSngswOgkn9j0arq+VLe2gaZC90I5USOlJjVZ/e8VbPR0oX/ibzCgCzcQZVcu
7rSlTsfwKQeCInk2G9i/iYUUBNeBwbWnp5JljBVKn61SWibARhTXLQVzxMQ8kZiW
1ZI57mKGe722rbMCDpNWuAehWiFWlANW1iLNIF6Txz0Grn6CiWJljk8m4vJzatUM
EXvDjrsEu9myRydDQn55Rr0jp5GZReRsfzj0qGiyyaInjSNFEc4BorOE0AhBap6L
b6I2IYpksSt1PtSmY/jHsChkpG4xslsEalfrI4Tf/Xaa4PHCuWTfaeddWg2qG+FE
fWOjAhsd+hK187tZvSXDYgilaM0azao4WH6ZT/fWDwtC6KHBSvDJntGrhrq0UFw5
fhNJfKB0F79aIqenfBqN1AtyCuedMptt6GSDnJ+ERalrTcqYphsb2FW09As03R6R
k0XbKCRz98h6uLULrloRHNs/bh2/upT8sK+txpJ/LdwUOnWLVQbs/Fko5wTLnskk
doIDv3mtPUpA3rOpyrFisBozfNHeJ+eHntZr/YPnJbldkjuHRA/ssS8KlaA7w0Gg
AXFX2+/LzJWo9x04G9MIcCv657OqzGxqcZ0izI4caJr/Afcvn0SzaHOabI3MeEIo
1XUN+CDCTkTCcXUEn/jUs7FVwxMafL+ptaWE43re/gP0u3Or+dk9RkbIwQdKiyt3
mgWy4PuEddWIJ9f0uON8L2rGn3MAPO8nCVUBgzU7Al//43y7GQO+zqhLO0XbLE27
lMRhIwsoAZKFXDh1rsBexJKj+z+7rKsOpSS7Je6CcynJ6ZRCT5hh0ehpaxV1oVGi
PtRJcZm4aHwSSgQhrzNRJMqdHaIEvI0TKzxc57bUOUb0IlUwt6fgoD1YAb6i9Mff
Bt+8LsAAjRZSTAmudtVTFKAAPIsvdhe4ANOxNAtU5Lhsm6j1xSl4v8VVV5M77N0K
QjZQ108uoE+yAR/ztGbeQtQbKpTBr78OdfT3bkLykzzihJQyvMj+FKX3WiO3Zama
K5F9P6EpTHZQ4Ga521UWP2eYfYBDJ/U8Jr4flbYi2Oy2pMiBXNcJ496XFkabzz2j
X7s3O+k6I+vAT6TFceV6UNu/787Ec6HK9co03Hf4DZNCV9gBeyW2lw8SD9BLYWOG
d5RYPa/o7stNGfc9fMeKs7MGKAOPMumj4H5AMZvNc56CNYbm6yzxs8KfVpvrD2jr
9T5fQTVY/0+fTGA+asyBt8le0ObZwjviN7Nvu1iPb3SGmIQ8eBsm2Ud5LTibu88o
/DdAAZb9JC9UuhmTZnRCxxbcouPNbWKIckePUFEaA3a9T5UxLy2/zC7XTqTVY17s
7E7hVUMz7KFglCzi0zT8I+0HDYn2YYQlZGD4ByFOad2hsXb5B+rT/xt7fvTirMrj
MuuNbZ30rV4nuh2tQug0iXZcAdUWR4uWUdPtjYqhpNyyZOIB1lIuVGFhMbxhsS9Z
sweHFstoGdBcuM5XwNPLYItRy3EByfy7bGDscQc8xxA=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TEQGz1eM+X4CcogfGv3Hss4ZBSY3NUgYQfQgCe+iCZy/GVROIq1lwQF3XV/pf8eT
9+nz8JUdIVhSftGZswfcFyBHqWaWaOQ/xUTdg9isfjsnrJO252cX6c49YTza8Caj
uPl8d1OjqmSSl8dXApF35CcAM29EtLCTjeop+/+BqHf2ZmmsomPI3oqkHf0Dz62T
pqOCOHkgkXISvlCathKiWAGMikAvIA2hTRWcyFMhqPtY7bnoJtKZ4i6V79YoicK+
fSdm7IJ98yw5qeOM8i3Q+R1UsaPbTDb4ml+pzfbs8PPwGvK4cjEGvwrfGHxH7uxi
IDekXh+196wbfaUpNmgACQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8016 )
`pragma protect data_block
blddUqNze2VWte1i/l7wn6ASJQGVrMWN6PzEZeI5/UVsfgVFZJus7erzisrfLVtQ
3zApvSmfUyAnItASRk6bh6S+vt9ezOUrbkG0k6kMLsI3fvUEe4PiiWpRm0eb2d7s
Vh0/osF55hZddkajQzV+667yaplWrLhVRjBVCR2Lwt1mRv29dIMfxMpU0J4iN7kr
4hDN0xICkV0HuYKOQsDDYqpd7AgR3bB2uQVHfRPRKl+wD7FqFj4Zik8M2TbKn3br
GOFmW0oOxOhK147jrEPhve3nn1S/ZGY8KhCfOSF0ofr5T9wURYN5SwELJGpEaBJb
fNV7xIPdDx89Ybkpn/BQ71Gk0yKPaSqZ9vpXsbnb2FdLubXR11IvawFi4GzYF4Ab
yZH54BLramBaDHsCDrfW5k0zqmGXV13kJlaZqGVI0Xb8ZDxMk54gOjKRsdWM9yr5
WmSmJUKX9SNWtjnCMFbYD6iDooVVEaHHPwrIXAmKbAin2m0MZixkgNtx7i3VvygA
cV2gFKh7Wxi+BySsaiUzwhL+YB2O4xw3yfJs68HzEgO8pSR/H/b84P4KSEPuU2r2
sAMMYknRmchDAO/m+QPtQYoFPGp1TZe3lxrRrz4UbAeQkcNvWAr0XWfHuL5nqV1b
wRXhNyomEKPuFpywoq0ezHmdwtFEYfpwlNpPlEdyWwctkagGWn9wbCaS8vRunQHR
VWhQnYhJX5J4zER/XPvj9vZGZRfEr/QHizyQMw2aotEkdFuI/fCipTKVpZrw/KeY
fxAB2DHa/BhbS5ECLDy7g1bxtmwktwV8pcD2eYVzi8ZdFaeJ8LYqrtA2FTuzCbNw
PIFYegtHV38XTUMwL4ZdauORv+RnZYwV27o02QNqGiKO61ifaZT3mLcpBZFE+2kh
UJR3uRML/OfjsbHR0WXXzIfQEqZG/GcT2AolluaaZmlwxeXYxMkAnzarRNBTUHi8
X/klZ0mCgfEFir5lcHbIOfrs6OOgH9K5nDFhVjrq8+CiUXMHCXNncExVgt/aAoww
+UmDnon0UNQuGOc2izs+ON9y1M9+ZLZg/V8DHTqv/hwCFzOajtWyqcLL+a2HOBFU
WIkz7/ahhPuXFGJlyJ1edXzExuj1N5YCvtVC/42Ow6RM+sdL/2nzSzoq7xs0daXg
0v56eCma0obZCJiTzCdrMK3emJLzZjzA0FN1B9O0JhgVRFnLVVo+bwIXCDKnrhfG
Ivt/3LNR6f3pTh9+BhPAdXMk556J7jW4kMruOJHrHfjVFCiOmAvOmgVOLfUxFO1Z
rqXRbb52QvPDbrM4GdEnvAP16iHEszXhDBK+oQeez1tyPOjtAaEFP7ZOid8pquYu
2VTVvnMdMu3UnTdyyS1IHN8q0B5HDEkfguaErMR7vtOrg1gMYff9CFN3lQ67/HJP
GfMjEn2zlnVii+D0UHy6pMWMhVDNsi7a7QBrXZ3z4M6ShhtCFNs9AAiXsiGQPENy
pgiM65GLW9T/YSVP3vWFQ+DZz7Mej8cOGXtfq658Zz505zNrn3xH9aGHtP9Wxz0D
AmULgYezkKzh5aQRhBZCxtpFNBCLk8bl+XXufi7W7U/MJKB1ogFi/6I0Ox0FLfJu
vyDuXetTqtvgrx+6QjMQ7LkbI4cGWC+Hwr9Jo4fbbjYq5n9AvBnCXbnYbZbQhM2z
oqD407wXDXdEiZyyUMiO0I8ASj3xz3n15rwULguXwvjjsp+rxPTAdEQRthXmk91S
td+tM7DZMHUtb3F3nNQ4oQlYuM/1ney23oMBybYdXb3X1iTRhFBanCOitcNLpSgV
MkFw+LOk1y0NMAYByKG/06+1Y9A903hk9+uYlkm0mFq+6x5eUpPMi4xxNxHHNBL4
ECax11cyEbSuQep8RUl51ainnUfFgeGj9QwyXg66L7EvqLhnpzA+YhehucviRD7D
42DgwESFPywrVbVIF/ysqUtvV3ZPtY2n6TCmdjhovqF5f3Op1AH2+ub0uKzoIKMo
eYltaA4Z3xz+f5ixL4xAXr+Eim/ZhNOo2oH8pFagwnOkoajZKu3/5xN/ym7ihLg9
dSan0qFUmvq30tByzhP5r4tFprS8zqmoyJ/ywup7kKBuL2/Wa5G2gE8lQ7ShL3ri
LQdCI/xZJD3BZkEKVnEI8mf5JgpEK1g7JbzPFQdqhSVDtc40ZeulHNB/YeGVFPLx
qNj1FmbGAWxROdYj/6x4+Py6mHo1OreV0w9zMpkmDCLgqLLvdj/+FESGmD0wUu+p
rxC7gIsHTmZF+NX3hEVjg6lQj9yb3RVLezoUzrnDMXvUEjkDfr7/X7ZcugdnMeBi
jiRP1LmRwEkM5jQtl9FWlA37AS/nxtmfqkGV88AoPPtBOwjV9rihov4y7LTA3vHG
igEW0Q+XyWou3/vJMWLb8Pu7rC8EwIL7sM0B6GVpNER+NtV/kgTf+8Wd/k1DJ6pW
etAyxjTiLatl2lH2nqwJx+YxOUPDguuvru8z+YKdH7qmnTESn5X3PdKajqcGR08s
+2tHQvvxiRkyjlZDZiD4ZZ23KEJHFWn1j8XiCk9R14UjZijC6sxkHqM1b80IXVQ6
cUbbAuJ+n8Rc4qrgHWNSfOFgfRgCiDjwPOVUlM/074+PEQppvkIwLsmqt51tY7v5
y6RJUcnEKNb2WpqYypxHoVaNcV1+yVUQvR4sX3eoCQG3UsTqJ/mzPHRRRtUrp8oW
SBCh2Xco1uqBQdSHCA4Jj7JoiHCFRsOh4xs8GXO7aVj+UgYnbhuT0fXYXhJGAYX6
L38eip0O2J8qYdyc2IX/vftf8WlGP1kflXmBnxgadX+qRkZAHk2aTTC9k/+6XPGg
Mz8ubq6QeBkc65f2kVLhPMb3dwVOLpq/5CmTYwn3+r1Q6LAcLDIipgBvgIxiqqnq
Tq0SUsTtYRV3K4Q0TBCZEKVJxZsEez+/30o2sUuPIhjUHZl0ZnjxFRX/SaxOrrQJ
GKNke8t05bljEvT7EyrlnRTPs91ZY9Jq7N/9JzMKjVOFviv8SQDxW7u2xCXZG7DR
8a1zGPWv+xpERQsz0noVFSkOUm+gaULRaZUy7u6+m11nB3yT0ZOTtK1W4mNGwaL8
bxKf/sx2hyN+QC+tWpDepWQnG29+RdU0LAsyYbc0GRbcZs43+5JPSRU319Uuty/N
8ZeWYI4v5HETWEoXwekaek4FwQoZUOeynW8sb/bS8NiWDSidvm1GQizJcIrhARNu
bW/mmc9ZzI4ZDkBc49Brjnf+UP77MPWdBRztoBdwQiKI9y7dDo61vxCHZu45BGci
GsxEIJcMF7GU9AqZKjvqV413hAGUeJTKGRBr4aJsjT0sHVgnrpfYFKB05kyT4/LV
n3NuHt+KNx1OQL6tVM4XbNslqkz69e4yl8mqOyuUtT2nEy0Rk/xWbSCgafJLE0pv
/o56vZE7AJAplMtFxdMqU+Ay8bVZivgsXYlqD4KDxi7+5rZVIkF+eLCCBGSAhpe7
a9WqxkP26DREqJpdCibLVErJ9sTjWD1RgEhhCE134QKVMsCqiat2AbCUMlpuTCJ6
CCSEDmhZInKusWO3dtHwtV4MDRTCtD3dawe44+fdbdJc+Jit+rOCxJs1Nbcf/mDY
4tmMMl6LdOZDFM6M//50OVVVSX+EkehMILK0agrD1sSy7aHy+NVDnXr3Fhp5fe7t
MXUNZMstCIkaKSPbtqp1innT9fzfeKSNR3ZoLdL6plUL5wP95xdI+wffpl5+dKkU
hPny5Ky1zeXMh5KX7wFSdEC9BctTvMaoVnd0pqfj4HdrOOalFDOfbSUaNIs9Kqkd
HZ73qen6T8TtzA61CqT6e2AgiRVrg5g7MeaAL/LvbqkyA2H9geKsSu8DgzhLP9sq
PVwgU1pPtu3csD+siSv6gbSR/NZ72jYaCallTV+gUUMhRMBgu6zqeWREhvVo90st
eu+4++K5VjgmMP4UqQP/qeerDBcpE3Wjxf+C1q1/eOlgj4MeZ55SpEaNSxdXHB7X
GWd77Vyz1Ae9LIE11z1yxIhZaPp7QXXk7iOxSkL/Sz7w58BtlgdjKXJCGYju/e7v
hFk0lTanO3iJE42c0qEHkMuQyq1rSLb5iO941ZQnbmgA87fK6guXdCSaUKlY6kDb
fZpDhU+r+7smOxSHNG8vUNaJf0F6Sw/G5mkWYom85Awni2h5QSig10xEzqjuLaXc
sw57wx5F5K+GEW9yjyJegUv9XdRoMEsg6ozG3GxrEoajyuLvqsx82zt3i8SMBfb4
O7psl9PDA7P84+TqALqi7inWDPkAQb6lMTKs8GKfU822qi7Mnf0zCxKFa4rglPCl
0az+cyxLnEbCEtcV567oynwhLsaVC1S9xQUtH059tr6IlViDFDqfeevfbw7U4BrJ
sV7VyWxdmAUSkyfRTnJfaj7yzLMjLHJRxOj8WAso2o9XxzJkCnkyJs+H6FsBWWUg
o2RUdc8PVKuFt1o1jXaPHwcQeAT/tIFgjqqcpmE2Hr45b9XIANtHBWGoopH2Nuf+
UVloemBT1vtCKeB8VCp8+Q1lOcTqnlx6S0e6Qzs/Vdv4LVf5DEBXf6DQiaXAR5e9
gHKCf1kiJGzcgUAtv5dlgIsbPxKKv5VYLrDM2VwoUxYwVezjEmVmy+AMw5wEySoi
7uZ/sZ2uTpJfbO9mSD1zennKifnSvDEKwwNPzlKO873Onb5AAsbncuCBVt6bzp+B
TKBi+jqZFsB3QMRav2dNMhdg+3M7p26B/MaQLp/xD5zwbyuWQLeMzdjR3jQd9Zuf
26i8zM3VPjrPrdpyIf4AaqgWUG3NHpm7fIcyf+r+whonkmg2djCXdJz3JyLVIQZu
wWCWq93CIh3+JQu6XUQAbliLPR/grPOqyPX9UiFUsbStcX3mj1LFwcAQN9dofQTz
k0238g7Bi8giYRYLtxIEtRzRBL42CnoQSYFDIWkddhmXdQh04UJhessGxcT3kBdO
qqF6Y6so1EpECC3pDoVDCPXlDkXJ7lMHMr2qu1B4JdZUqaA4otStV/frFaymYaoy
oHM5ScYdXMv2K8SIyV4iV+pOiK4dfvXrChFSbImJJzktwxiXXT1ERiTrn+WlSg9S
aFjmPyAdMbpntVMBzjBTRSsD0wLXCDKCBjL/PS8U/qAliLwA1ToI9s2wGgFguHR8
/j6O2X1XeOOOXRoxYQ3Yr5qxHXs1RyWZutbDKCPOXfy5PKFA/CYItrImD23lVINc
qWg/5SrttcLCAYEE0WMhRtYzGcPDa+M9jfVc4lq0D8JrV446G3h5Nbg1H5k3C0AB
r/AogYVpOQ3ZxhMi4bWLmBkUXh6qbx8XfQr1xZq0+7FRTLaoRxYwBG5znUf83G0t
wfsLvAMo16PkcaqVefC8g/gM3OX3Fyvu3ycjsrWRmf+HgQSXhkLgJf6ireaBXu0S
tLhsf3v+J1DyJk2kqoMtYFX3F5GtFiHQDFJOS4UvhOqaLlmdmFKLodSKdzKhbCyf
D+hbPPEyuebS5aBpPSLynv/BTAzORK4oE6wY0CEEJmGf19QZe8QcQCtYWjQLZgYB
CiaEPUexvHDv+JpegX2iSVsIsFTQkVNyJSe+Fqh/5xCfbe8c0f0mPxC1YneJyHha
E2CFSvteD1ggUKF4PcACivMLKAmdRcU8A37iSK1bMX4/JqQ/vVbT166rtnVGoHMU
C70NUMSfLHDSEpJ+AFiAULI6Y6rUA6DrYqPLxdZYVcP9LRsg8PpfcSm60kCd0p3l
aEa6oYbZwCircfhoOOwRdo3I2inXlIrdMGGbnYvOyfmzn5a4XiADzF6nIyCeGT7O
sNhXfWQhClkp9mL7QVy0RjOuPDJr3CMMZ41ViK4zM6HqUsqGhpyGIwzm1ztrpVxn
Nj8tOoBix08xWBbDVVAdlMwdFJe41X16BmUO2Giv3Owkexn1pydjglPopICPZ+QS
TAQfEeQF+8rtdENb8tezRcXiBEpCDxIg/xcvSkDjedN4iybtLgwt8EzjSQ66HP16
2GmiZfi+jWxMbIfP0n5mhvh1gYW4qNk7paXo1ea4pBijzN+wrZBL7Y5QUKyXEDer
7hH4d5sIA9BKoOL4v+BHrXTaeLdNfoe7FL6zyvIUusCKkCpUQVRxrAJuXb0Am8cz
rtKuVARlLOO85e+3l+eyHdQM6ge8ygTrt1zA7x1Lk/sBQlmWrXjCggn6aESNq973
rBVBOXPERKofyGBZHWcDklYYp8gKTYsLPs/4Ub6hFHlwgRsIP0QAItcqvY0lWrqT
TAIG+x7vG9G5oshUpIC1brRVwotRZq/Sa1DyTIMXJiJ8aWYvQZWgMLgUeeMUxP20
B7gxXAEgs82I4ohbM0/OlI8c43bed466Vpv/LM04Ry8aTpYE21lqNi/rlseUw13/
dY0/fRz/n3cmhVdA26bBTch3wo/916gc9On+nXfelynPUe05ZHWvQzrUsqhlhRxE
l3pQjflMeHe+MQ1lowTZdVOm+jcBGigrqo3z9eVFFl9SA+pgMxYCTNgmrW9xNXBc
NwuJmHDFBRfy+eiek+kQ8BHNAXqQcD89+ctIQ2/T4LwV6/Hw4spzxaNym0Z9w505
9hAuwxzOd1hrq3WADyw+NLH81OjS6fkDahUuJVEDZFAFXELwsgv6R/uK4DlntG9K
bMASQ+SS+UMGUPiSCwiTocg0fVHn8wL9vHiYvUki3O8REqI17UJ3yXAdXsPny5xW
aPK2rDjbLOZt19VVOk7xTb3mK7Yl3jZRfV/V4bgyBUWEPPySUdkXAnMJZeAcJsiM
zTxtz5mUPxirXU5o7FKJyGTT6pJiKYsORmIdoy9ZdlIPdz2Zo/MxjzPZvTxN473m
cP6aAYBMoU4W32E6RQi88qTyrntJiz9qBasaGMbodi5LVTMkYzeTchC+4wJImUaG
a+/JKGvb8UIns2px3EZU7rnPA9VNInfOAXgBOV2Btmr+9znGu+PyBD1RuCh45dDf
BCbpllg5CAiD5VLiBVL5tSOvcaficurmNACEd7vhD5jrjwqtjeFBlSkBqgms0wJu
4akhnnnitYT4UKYmr6rOITBg2Ru6N7GBWk1Zfc3Eopnc8JQkH2abmMz78Uj+B4iT
a9OdvyhEGSoKd3Nb3fjmuZVlrTe8BQ9KvCcrC5oU5M3ZF4UwLEOXB1b8JJC2WIP7
ezo7qgKgpDqxfYUsCXIhdi8Qn5msACwRUdcQmwNjwGanK7Z5FvHfyfNsJUWub//q
QeOiFSRUM5BmlzWT9nH8nvgOJvAAvdMQwYkZwv960cueoQgWcjOoNSusXmKFIvdj
QrDFY4hnjjVO2nSmm8ZI2KofG6u6Vo8KTMrqtKc9BeWpu5dbJvRI0Bmust3pzSwE
vcHaEYjxFeajI36CAorUxS0zFPxrbZmW4HhVURAiIVvHdxm4pc36Dkv37114K6lt
ez06vaV3XHCHU86fBuS6HZ237vel2sXMOkeJ2HDgwX2G+Z8svO+I7ryJfAbrHBXG
XkPh6rC12cKbK7LE1zW2oIXqMmPXl/J0/cd3fXj6MZu5HO+7qJ769+7pTbWc52kp
g0i9RfOafb0MPBLsWxxIzdhKBbNhhO3GPxKUhwhvboYJcK4Prm+pkfR9eujVVaAG
fpdyKc5hl+mTf/j0686mChv1hwHn/GWSDU5l3kq13Og5+7FXUjwojaSLUao+ZiZW
AsydPleNF3Y7+n/pvBsAZEGgUlg5pnt+Z6ZP7W7C02AVzTqhQxypHzWtvkvLRV6D
Q74yuxzMSgszDky0SgFrGPilybkD80ayGOesh98ZgvLZjYFYzkwfld1YknACV/VR
fc/u2D7NGZ01MwwXNdv0ZTJmvkRmS0K65e+WcyITK2l9MkKy7b+H6Si4wXaD0iZM
pqP5S2ppHVIO3ZaEai0lMOKC/5E2PIxB0XdhaPjAv5pjqHv+WBrIMv2qneN5RGYH
sBrb2fHgnMm0JB8/V+LTnBodbHh5u0r9+Y9hrFUe4+flpnhK51gibjy4nnrdAHyT
mPFYUX0kEYvD6YVimcDFtKOyBaGvvurOjsCFOP9GzpBM/73rlV+quXinvrLf3JmO
rBnlaFsRSiIqPMUhcf9PQWMdIQWzTqqXGn8TQ+kQDFtrsW0xSlZQD7pbmaExV8IY
nqWEISkrdx8TnQNIDkCi4jHwkKi2+35IJCnDdk3Ptbc9LIA/wpKLr0E9uPxECNUz
/abLma30oMs+3fKyk1pXgs+ZKjU8EkTC81cFbnbSslva3W+l6fMXXibVmWtNqTqu
wvQ35QuAuJkLHSPhsdP+roS25Ir3zX3GEhByVFjNMTweIntic9+Q2gqjANJAFWzF
ClaefUdY6H8+3mqfx2UHXo5m7lc57fO/6R56d48/Z5/SdPeKkW3EJ7eY+bERf+YX
Ar2n9D3PhVlI5Zkmrni6njzRR/5UE911WrZTF3Na4G0Jj6TwA+yPeDKoL8xK9OWk
UvYmx7uHcu1MPwT0CPQf9osFBWw9xNZOPiwRJyr/pMdIugaGBB2nlyMcj/eKAvwr
0gZfG34cSUNlThy9MfP9Vq9lzyafMjz2ICb0epO8pbuA1HDG313nnXYyQwDLpxD8
pwhTzZT636X/uPJouRBt5DGhe8FLvaLnTjBZ/caBqGvIfx794+hjZ5AUIatNA4XU
2se3j33PIm29Q8GvhR6NOtthEus3aHve1LtCcz8SiSB35Q49CD7g8lVBnGtv/wCl
4zhEHILWeFhjPhS/qoCKz5lQhh8v/Y0qiVwYg3g/I4HSy7nhuD8MjNho2nR2EKIG
QWHcux+7/GrCKwBdfG5WrARfhEWm3Df425MGtk+X32zHCHjAsYenzFjrWkn0+PKQ
Mousl6BMYIXToUn2mpm/5QiACKO7k+kB+bkT2wR9rihuZRNj/q1eIzaQRH1Dp1b2
CY17JMK9wT/mbw1RLfzf3GUVBlG3LF4gD4qBDaY3pG5mRBkRZ4FJnwbG1EyfCzj2
Ik8zE0x4V2ILdzPTqDz7RmuI3mqy0Y9ffMvQ0HS/lmP6FH5bUp1f7SBBcOcsNGW9
iltG2ZpYW6R+frZvOHT90KozXh93jb3rg+ksYICKTtFG7D063BXF7Nhp5bnxfw9A
koqh6JXYLyh19cRDqqn+xZzSIobMTymVuE67E277XckLKobFzlDfvvY7k2S9hozv
ZYS9XG1hmRgDIJySyvPhSwfWw93G2PDRHxok27eVFfE0GCn49dHYykfITMAzeIvz
W8RJfWJvc8XCYXe3MtOlI1Zz9QvXdpwUiNdJtv1xh2Cd38+ZIWe2VhNvAoOYZQKP
tZdcWJjNAC+2/Z1aYLACZTh5OfYh/3mbyolEPxkFV/LUbSHyNxcT847poLgaon5F
hs7mvrZd58sHLRt+vPKnTtuOV44yfE1a9khIZcA3KqCE+/vfSHY7IzmpkiswkW8E
tr3BGUJZb24dz20NshOD9z+yXjLmy9ph/o4eUYSw7qQxPSBvWK5g9jkFa3lGKQNs
84C7Ob/DbYh37rcFHKUQrp9R6uPo26hOAHsD7yv8/2kdzCUh8eg5QfVvuTj3x9o4
/uK7jJBAJc373ujjtzsMkyQwsEbNAYDYBw1lr7S+bPm+W1cCkd2mXAzGVRhH6bf+
UVw6EnX0ZJGrj1Cfh61NUrP/ZkLzd9UW6aWcDwRqDGok1939OXZnuDVY9WSAEMCN
imvz2k10KUMX4maXt5VneUkRkrCFIsuOA/eaMxDvQ0Q0lpcqFOfu5Q/0vmKS7V1m
bT5Ln9VrjfyKRXRbB7AwcvQeEGZXsEPvyN1L2RizLfANbLyPfkRlrOAw57XOCW6V
avboadEOmoWsn0Cx8/CZE+Ckyw40Zrvxd7Dn0muD/T6V/1u8TIrsbx5Qb3jUNNCy
euegZGAstKghQyp/uVnXSqcwkPaoElwkEX/hERIa2qmDDoC4PiaY8fQdlVogT122
cToLbHfR8PNXURfiMhabpfc6bFU8hIgKz66Leq38dUglBmGrootbKjM6oS6iRlU7
KZAa2vD/+6KASOLyeMiulrNoLXPBbWBaoKP67t6MOM9mzl75wIxiiI2vBasgd7wj
ON8gkjSJNVEsNJNh67E+wEQirDRia8JwTy8YWYXCA2c+OrCjeMW51KxvA0ffT5v/
HcOyp/tSKD+2J2LPVwUjr+mu4TRPyyzCMl+lA0pXQ6MPFSHePfzCTHH5wDb+WbOm
7NJwTpKbIj5q+kUl0/zvMfswbKDDRhYBW1YuOnZ8d0b2akohkx0lpqIpgILwCo59
KG1XE/qt+qtUKK9AX1HV9Pnb1wDQhVfLihC0Mac/ZJ9nfGUWl+jp/JWXGAwCl0TR
yVikkyp9UfF0UfrUj9JgvlizV63fZdpu/D9RzKxSAMV/GpaKdyZEKitZQKkhC6RD
ZNaQTQ1hgGWsGf75H1EUdHcQa5bnKQmPKnd0F9D4xuTuimYqDo8aI7xBzd9JV6vW
mrQN5qxfibl8SCs1QG4pSPg+HXyeuI832inBmgfZ8m5AYPqDGMgb9weaWMUTswLf
z13do8Gl7FHTH1cyeeeWQbGKJEvoBbg8HUHpTzMiic2JkrqDi6zp4FPzzAAlqhZm
9WQdMlfquQvBFnSZSbkt/lelgeYCJ69ues0TRvBpS8/cp/MDELbDSOYUaDi6nFqv
SgrBkykl96fM/fih9qtEng3Pyz5MZUNkgDUBwesN/JhzEJzx+V1iVqvkYT9fG8MQ
0JcTtceU0hPh0PCqbqAcyhLPXNbSaAgREEtUl1aCEAoXuIyppI+K0onN1YGJ752y
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Q/06ewqHsY8w51Ydoc0UOE/9CrAoiakm7nKKdCotw1UturNdzsbFDfj7YXKRHF7V
jahn2O6WM6JQFj+V9mmAZo3D7gxXDEF0PrOA0pybMT5zA8pCnBi/VrOmKOD00xC6
euHdgUVtCGjoJkZWtPHLb+RXY13wVjqTRc1/P46qjNnA7lfmQsP5eDwA30JNBwFU
J0D4zUrInMP5nBzA0xeY/ZQrZPkZYiMr/LUVmq8FjPD3Vw0NW+oMmpfiD1rtI5Ds
CWe+hdvqUWg9cpz8khSpCJ2/xmDTgd0ZyOLJ2m0GX2biCRz9FqWeKVxOuAdknC1r
WnL+3H38nAMY5smn35xgRQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5392 )
`pragma protect data_block
mMBckLbdStpeZt1eISj304+OQ2/eMXu2uq/uUujNgMgay/HHuKIeMxfFZj81HwIX
qZpp28zjLJU2lZPYuQJyoXMcBsvvidda3PjYRArBZwGqJn/4AbIIA/qwq2tWr6mx
6AvJ4Ip+zuvymy7y/5mHniODlsVWtCVhHHnarzuSI7XMw4Vy241AOLoPCjFf2e80
0ewbCjW+NDVuw47lETPsok+ecvOXTxVBd+dfsX/3nhKzLrVj8EzhllImHWG6DSFP
vZln2yLfFDvnNZDwJv4HDJAb7DlG8K8Hyv9S9QMsvWckP3gjqEpnSjs7R//wWM3C
jYkql72Y+ve/LlODUPTkGk3QloqMu2wLCPiJcu19dhoM0AICt3uOt2e8+AAWoKdy
+7X71+UV2ERX9BQoIWLB/fZ6TKzxX5jTDvsO2EB44FOnF7Gb8wjR/ee9faMqfX0c
iYcmvqBVumtGB6/Mzc6/7uv7t40RqNWtIZYT3bVnXmKpjRR+1kTZgLHXk9LmsXSD
XWNLq9G5R2Obzj3MZW91nXxW0nKGYTbKukLXIQXgneGmGDcpGMSIY/DnSag0ROMI
OD+u5YpKqx2XvdvfKBKO3wBJXrQeD1qvIPGe14ssm1YejKLuFjgVew8YdwB/PrUj
9umVT4sX1f4RbA40rNoopqN39PVJuqJcKmFQlgMnxcsDS8HGLIaFx2n3wtd9h5eU
IIJT1yDnf5ZDlxUis168dR1jxoRqi9jZ1zJaDry6ziTtYE1aSbP8Wh2jSUvT2ZPO
OSanAthx8fvqMhhs0nI2qyGNJ3IXdROS656DiKRy470CegULkMMvPkJ2ERx3D4wj
xvgvtazB/QIcoV0bXk3/OAu9jBzgv26XW+iTaQZD0TXQp+cLAyFIJp04iUmsXTLc
PHUk2UBWTEhGCsN+TQ1BSFeOUzwHWVA/Lrph+enTMBYiPVk+Vl+9iNZF79foEiWM
uLYLj02GprLC4bVnsc1CwYLQzY3urVNah0D2Ryuj3Gp4AY6sr/mMcvAGsiISqDSf
Z6oBZC8Tdagjk+lZBcEYfgMM4ktCsIH6+iFoB209gZdDkve45fV9V6A99DnZUIbq
cx0oOwjiEJMsLeU1KXbnL/wmM729z7wUlEZtHJSDhYsgrw0b8uIAeclBMoaYByEp
FVj3HW8Cxgen0FfmXjZqmoM4eWfEe5wMsA3cB+05QiPBQSXN22Xka0TGVn2h4f3i
IE4KqE7MT462CUmnYpFSryasfewUHC5k1gs7GZmxJ/ISFSE+2SLMkrz5DH727/T/
lJnGe5p70gVDcazLK6o77GnF29JIMdzGEe+mN8PyfyTdtn/8eOj5d3AxFcjc7aCm
XTCd4vohqHQ+rQrkFpjEG+GN75b1CplQ67IRGuI7Ck+9i018+/Ic5xC5lV9EWsjZ
oX9p7WJCdeAjXaflpKYyY+dbFdvjZ+ME6SN9rXpGYf7m4qUmmYP/7NX/UPV56sJ+
J9Qq5KW1cjiWNLIuF/a9qcM/KhG3kRcSmTTmTWqe9Y/mUKHdrEC9P140f9qQfv0w
M6ShkfEyqJ808p3wHFMjdkpDuaRjl0IeWS/f+zvIlF5SvZYICRxO2h2kyJhQF2wt
JMV7vYrVowm0YVSHfoN2/VZtW/61KB3pERYUkxieWj3DNe9Kw0io+lmubIbZ5jri
VhG4xzRxV65ShFKcPmcVZIjALMZGgxFORxKsNNr0qbl+qWsVsgT0FKrZ1FL0zVZx
2NEymHMaFNd1lLFYKeYVdZs9j0aAGDWCJqVoYpePT9gjMhy3Wvd1UIeOjCGvpvs5
+zGgcMt2tUI0iD/lhJQhhCzn22oosm81PQ4bEaCPninTetiXJUrcr2/QtSqYgDwl
nJ4D3K/lCdUnfyPKcEkkvqq6TZCUzv0gNu1h8zDyn3groPtZmxoMU1Q2i2jueewY
KIvfJtsl6fpZFJFh0ezhofEu4QFP9A/ZTeIz9fILOKvVpkulX2kGwNxYq3KF1g3A
YH9qO3h8G2G+w3LcBxYgty3rQaALBeS4OvqQsi17wl13y08e+oQuz/CKJGYzDrRe
oytFQ4qqt4g+abVIEPocLh+KxaHRgRXfWP5KQN7yDK/+8YS4Q3RRNWBIYsLOsv+n
VLdaFDi8lOS0P/JA/1jNyxvKY3ZvHqMWQjyiW+XoQ+25yV2Q63txDcz7fXpAd5f4
VF1w0bGaqh0YB3wzM6mEAeKFQQkhHIctsARx4hNw7KjylttRpOvzmIsfw3v+OFGM
f+Q6CLY744AbRH0LQh3NwKBx1LdN+sJVt+Z6yiEDWGcJdriLfJZY7WtsapgjL+ro
ss60pvRmGHfBkWo5EHyg7ubnum1boVfB59sA8nbEOMWzYX81VUbXuEyAFRHpPkFK
0qICLr4+tFCT2be5D/CeSnOk4nt4Aswa1XPl7u8OlLdCXssJZVL0YX7cJXJyMv9U
LcQu5Y4CKpI6SMFYILlPVN6+nvNdBqupiplLe2TKVU34Y8lQQ55vf7TSnVxF8aCq
klR40HbNImYIUiWZ8mLllw4wfqsGtT+sgHCOrfCGzbC1NkAG2n6lmO3npjNPDwW4
ocbAB70Uc3ZCIVxykaZA1j2PwCKlx/kfZC51VqpEweRIELiZChavcRzIcQEfrUNP
jv/kjSCKdRXhgeK0fjSI4d5Y8XbGek5238K1WpTD6393Tf0BmX/o9n5Gb5kZgrlF
0IOr93Nii5i13yhPQlFq6toHAK3+Yv84KSRXe3ILpxWLFIf5S+DERCoL7C3e5UQ5
k7TnJLmmEqlMSGh+U/CvLqI6JbWgVNZtwwGlTGd30dm4YO3xLh9/Ei09+4daz4PG
x+ZiXtKa+U2GiItiZ7ErMjLvVXSUmqh9PL3ITQbmLmdrQLsFJozN5SA87FMt/BHC
UdC++vcJKdMYxy/YsSw2wTgfqIbZKgHsyDjhHKVXQEu3TY1wSxasCvBdPRigvX55
Tlxty+NCeNpNkyLKI0ilBQULYmEhirMnEEg6J/95BomhN0OS28xognZwATQfHarr
bVJwaw9lKJ1y+Rv+oRHdLZqFDppRF/7cEHv7DIpULEdltcffkSmP34nCSIc8uoq+
iVvxMyLKyu4pyYvZHvZavDTuIZpb3JSxjIMJr7b1zwRzGkPVJcBweH6OqehYVwwJ
TVGPHZcqohKnb4TubMCLLSc4C8Luy8rGrQcypvp4DV9Dk59m2NSFdWQUpWHXTFdZ
F6u77VVfUbENI1rAl36MCUsVzP9EFShGFhRRmvb+Ooh3enG/YcyuZo2VgpgyRA7U
LhRdGCQCXOmpbcm6dLh5EfGTqKywRxoWMDUTrva9+nc1ZrT01r8c9VMOy+THFolo
+9hjOUbMCaWVeYG142jTwoSqzZdKQp4uNb3qIF0B+iiv5C37rCshvLPhDjkfSfnG
RGAihjGtP+X+eBYxI8MVTAcCgDnEDeQFvZNbYrJFMpMHih8ImC/PKBw6wBe+XvLg
sRXsYFZmqNORDCgjad0hT2fZ+7EiMnd5W92ewT0OsKCtJIHVoE7fWvSHipAGJspG
xT2UaJO6zSjfyzFT2g418kaANwvHd8Y66bPJQNyKtHKzj/55/cqa5Y7MEtOscWZK
QG7oZFcReF/B8n9cf+KvCoug+/fc96WN4O+gzOyGXaB395uxoKYyyqlV5lsReRPa
TGqHjTRY6tRb8DIxTTf3pC6P7wQLGuDH8crL2YwTdvEklQJtJAosWbU+d4yJ7N4e
zJ1H3EZB4JMa7p3WDXc0kwz5ZZHSHhCKNcptGnn1z4BILUMJHguNiSAdEJdNSCMR
D6uECxHy3oPXx6VeoQJgNe1e0A5ICen0RnOG/sgVd+dc7qPcqbJCkbGgY6OTu7uP
AT18jlYrXHqzthdjYG29w4gtkB/wTnKl98SFBRiL+GVvfyoF2IN3GZDNponzX+wD
OnvKjxGII97vqfPqJ8Hj1MBXUO4UJAWyzda65MrIBAm7fjDMAWSPZs3fEcn+r978
WgEZQHwZTIy8cm2rGJv7VvoJKyngmf0CUlVNPknCKrpn2JCav5bYXRHsxTMBZmjV
poGRVkeWbm7QlXlJMYcHnlDQ4GaRZHDpyRlocwQE02OB2SQxagrfRMAtqhGcrIyl
kKfRlnK9rbTk1WKlEPThtKAjFdZnmJ3yNQFT6z66Osc8uC9YFdTemnT08RCGE1vg
xepYkwlsZ2DT8rFufXfYvqsOeWlIpIiRX9ZAqxeF7A1chTzvlesaTi/+yUwgXssm
hl3dd+XMhJwk2Py9lE24EfDLMihyt3wu7AUb6PeQN14YHCUG8lpwxpdlo9G6xYpn
QkXLH8WwMjAr2p5G9Ip0UlGJKFBKe4kLygMMBWB+jKZWSVE+ZRMutcx16fvuUQqv
Xp+BzY+09UnqlBWoJ7dTJdo7nrmvD7IGVNh1az4z5HW1iafnQZkXppnDES5NWyyK
diS2KyLNAwJzyLXE1HpsANPRKbLXtCKG8i9vQe4LYZAdXV1Ihf62sM3Z4/UKtCe8
UAIZ5p18y2vl0Lnp5AR9SUGS66oHD26R8HiD2FIhtb4+y5ktZhscB16USXGLFNfL
BKH2It75AP0GDkE1y41RrElG1AaXpJPX0owyKB3pdm7ooC6US970IfeN8DwnbdKS
BlVuf0FLMX9RERK20lceLyENZuO3BW/AHR4zSZcaIJWCO7TijvWFuHkoW+HSr89C
0aal8QKbvH4Xgw/kl26VPCjphQ5MeR5eIJFbb+h2uVl9ifKaJHhHa3bUFRKjxtxs
ebS8sUCLMUAUmEbL75ecc6qFEOD228KnVNOhfnEyQ3IAmSJTBttFmtKBEqt4oL5E
JsKNdlc45MwFdFOEZOXxMpFIAtwXIopfSFdqT5ek1QHqgazMD29gYBIgY1KJqNGe
V/mXLSKqCOLXPn5hs/gqYcG7cTnAhNcvuVjDyyMS2PJg3qfktiOO94hmtYSznjhL
NKTclzmoPUFRtxtPa432FPDrpsmDfDL4DVXOxMCV4C41hQ5Q8g/mp7RmglpcALF4
Ug3hRNQudBleA9He7wQknd96WfhEDd1W+sGuT3pbCs9Na+CHJQUZ1zdPUFx2iRjS
famsPGgj61GeE4S9yvnCUPK2oK9boqncA18bqGwu9OxHPZ9DEaHqkgEb698Ikk3i
ZHbPZtdXkXmfhUNGjpjEEXOhGuM9SrBEuA5yEVUi52KkdESGHUJ0wADn8aHJSVB7
LFDqu9gny2sK0vHPxyEOjZXZzYrQxKy4tY75WcCCSK6zk5IMupSp+brLXvXcxbU/
nizCq8o7ioxaU6R3PNHk/BOB2prT7q5R09vZvb9t/azDB7U7dqxtww+71e5LoAFn
ILSZE1NW18GEbAw3WzdoqQo/JSV8M7QXIROAqOp/JyhmRRThgkP7jTEgEXo4Uf6K
cXE6hNW+aXX6VFfEciP+DXW/9AuBU9+uOXgfQvhJDQZ3utEtTGoINkd+q4y0bl+m
vM+gXabdSW617N06RSXsF7ddmaP8/NpXeAYrKyZavcaZ8tgFLH7eNYmYNV14GSum
1BwFW6G5Io3S1pR6yQOtXU52RaeXGrLzQwIpSiC4W2RLzbyTT4Eb9QpxFSlGSXX6
vW2L5vH1XX54sPnQgXjlmAAQXS73q5Eo7hBx/yBhXWa/MFSt+gfZi/wOux+2XUNp
RZIH9YIItq1+oNPMGSdh4juSprQRDwRaAB8EFkmdsvK4rMrI29tVzdpkXFV3qMOm
hbHp7K+PCRXsLM3kq3WFTywm/1pZrxcWT3f2D/59n14JGmbQQGFxmulGdP0bTz+8
VXmks2usNkDX1mQdY+g1HtRLWiYoiscd1aIk7SMiVN9wNWPqDyxvzA5/ED1d56UU
Iqd8xTHbFgnwB0x/tHfMDVc1LlfIhNOKsldkyOsZIjLhzMgi0n4IpeiTU6eF7GlK
yQhhu+kDkdmSQ0l6sVe+7Sb3TtW1vDbS6F2wDOK0CFAFM4cjLhGT5KsMZeaRhK7E
6H93MwsQVCUexc1MrlYrSakiS8IgaNQ7ujxt5ubs7mqAv0Ox50hjpYvdOTQ6CwLb
Vmx+RjS6ytYTCip25w7sMIVOz2FD67XMO1NDt1KDYINBOQMiE568Oc1R8rbhow24
7dlo9TssfnJBdgv/P+TEQnJdMs/QulzOjoPtx3OvkTTm502LKNXhXdkcWRPfFlFt
pUT0PWbRgtxavjV0cTwE1wRm4RVT616t3bLj4e3D7qXJXPcGUCmojxWcbrki5vC7
/2CHQbykfA6MTaTjM2SSTZCpS6C10FpZgLLAQkfvNjiZRWObW4BPL/QNhn9yrl8j
t5R094LSlo8gIdr6EJrW+dWkFg7dESqsU8GVGUp7j0YBuoqga3GUpMdr/btW4A9+
oRTM6UMgD9zBsmbd7dj1TUP1X9FDlRJ+U7k2vTkjA54qDTW8AxVZKmqHciB7ab8a
lv6xbS1UgJKgSiaKlEbCdCvD1T8L7PC9gdt5rQR7zlHKrGbyS+fLDdU2o9PXAcQz
CZKoV2Kx3GGlpbNTI6BNXj+NMtxr6E14xpE1kwcVx8DHZt5yLl5eXogtLNMfkJzn
cq6gi8nY7+3n2FD2C7tNr+L00AHE4peH6H8Ktl7cM1Dr6Ga2O7R2upla1PIZ7fw9
Sn2UWRmqjrN/SY8OqsDlMa17GpfDtYBBrvUc5LIr/q6/TmIr+JOkWy1OvKkPcHB5
1shHEUH09plHmk8LWzc8sHPBAKrhdq8kV9GUBMNDQsTTz6v3NufXn8KV+HM1vXOZ
+WWqhHC0LTGfveJ4lshYwzTRQDfBF3W78T6P/bZTyt7RQIrAmup3b9kNg7XrgGEc
E7uBBRkE3j9w98slOESypLm1Qn8tIdyLF6Li/zhq7qwckkNaj3jqJdzrQEvxpoez
2t86CKnqguEnS1kgCri/MqASuUPdgOr4sKquAW8Vbe2sZa5xwocyCK+WDVfUVl68
dpJMY3iJAPTS74gk7L6981C8dYwN0tuT0Vb12OvKo46EoT42Gp4+RqMzo/btsEVd
H1j3QpdcESKvljpGcKDFXRNiKnTIu204Mk71TcAAnGwN2OCtiUTmpUz4Te1zusbM
q4Fcot6lDHOFgCy6T0D3HhLoD+28ZzJ/Iu0jh3PC3LTkRtHMCWpNtjI32zn4c18R
AST0GESwasM6aDygVK5TrHSL0BMQeOZnMEt/zqdh5yB5j6d7gHt+l/+7zdR3i/IF
b9r/HbwJRMq/zf6ykbp+Uw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
iFn407QTQuq31SFE0xrqd57U5rzCsjFz7cVpUmYXOkPZKVgYCIggAsxdbNhDKGGV
AVMQ+dUzkQL4TYAIZnUH68IaS0a/6l+T2EFLxsYWizNlGE+KKDNYjJDae2BmhvzV
54O50a8BHMVFOB+EHpsOxks1I9IDAW1dj1XOg4R47yqRjuUjlFcMuHdaIoC4V7MU
azXzR13DhKmhCp37wciEqdmEBVysdgqON24W0hmDcHVG2/e0eix4khrOXyb4TX2z
c/awtO9NqIhc6viQzlqVsgGaVPRZKvpaluwAH+lQZ88alCKdCiHHXiZuLGgzxsBX
03+KpHdtdfpVr8RG18ZoiA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8864 )
`pragma protect data_block
ylvDyBdt57dw4Tf5gnXCnMnSDS2lWDxVJdgNXBuSgIdifqgEpmCUxnlXvbfVyehM
S3oofA/r+dAbJRlSCSsq6EBvTssDIZfkr5x1Fjh6ZcexnEb+Kfo8omuI7hMUr4Yf
p2CH6/vPqyIS9IlnWCvl5o2UMqvQ9FSjoBbNAasbn5JHj3xrptrsJByHQVYU9YlT
0as/GEhsYL8C08mMPlVaJ4UvBqK9Zk2FvEqn8cccrTvhWdK4huvA5wF+7YMx5VNA
Hpd72Iu1lAQdtCNP1f+AMBl4Xq+3Qfrn0pPZZl43YAc1vPP0ZFOQDZV1HpiOM9YV
paaHngUjV7w2BiiiU4eFcPBGZoj38JZhNBHaxd9n4vjSTiBNSZx2Cn/hsnvlr6gs
MqhRfiyDVxIA99jqDK4+b2DbSaPzuIyJUMvNT/CicN23bT3rgJWbOShBbX2bL4KX
lesqelMCyuelFIIkohe5MOM5fk1jh3gQP2JwTmaYPlmrcp9cv12E8LSDsMpGzxeO
7i2XERtr1s9IgZch5ApwXIFkOecsrT8oFRZog/uyFjj0l1vq2pstET+AaXkQBwHb
IXAwdLr2QEkaGOW6xeEWG566q6eoQq1Av6AeY6VctuAl+ZuXOrQaqUfI0glRLBoz
gZ/3JTr0Zuk7LJWFDlxVI7ClnknBxfqfSbjSm54RG076aAyr778H6g8zTFokmxF5
m//zogrA2c4Po3euSXNXBC7ty5fd/fMAteVrf8dTfiVIoipObFIHSMU2ubzxT2Il
xBYfy9Ry/zaP36cTzcmyGX40WDxlfp9RWki4VkvErpaanv4TNr+X/6BoVGrrx+Jt
qpG6r5IDYqfZ7qfOJCq1IH7FfR1dE4aLAi1fOL9l2IDqkuB5s5IHUtqIFAERJpAf
piaDxD14emq/yHtyttOly8G1bjk4kX/7pDaDOrJ/VPjwTsC153Ea8VKpdnYKVscE
T/r3/cGMA9ahBgVYR00gb/FXU79kMsgU/e7oL/thKlpQ78qKL8CJsZfu4Wu/t6P0
OdhAhOmnoKrz1xyC/4HXW+kzj+2A6VYJk0l4Nv9h3NL8xoHtypR51bwLZ8OmTZwi
+yxURnLc5A62kwx4XA6K5IYlb7LmotMQ6ADKJEdWXosgienvjwdRjGsAue56FtGV
/rssaZlaKRSCxWlW776uR2Nzyh2ljN1TGmIiAr5/GEnshhIW4EbEobGRW3ilSIL9
21uKa6idM+Lyp1AaKTdcidfHokTfULMOJSXRTIj+DO0L/zRQsdmCLJCOuPdjACj9
eizntZbD3zjm7aMKs2f25rXD7ltftrSfe6UKbsevVUCZyt7FD7POYTWoc2YQ8WlN
R3l3b2+HIA4y8OKH6p0VWR496JfgHtCslgBsXo6NHtkqrhSfe3LCdbUs9lYSLxmD
BbHiN0GiukkDkLgG4rkH6kQTnmzLhY117bSU/GL0dIa+RjHXw0mMOujrw/tDwiV8
4heYz4GbMhZZ0ryLJbXs3xOGOSKlDG8rBZgWBnvfz85WfYmyitrIGSBroCPemm6p
qCn0s/iclOH0hPrB64BI0yHKgvXAABhW5n8wzJknAecbzwu7ueZBHJCgTo0SHxJd
+THirRW/gjGQlZJTMYTo5jk2iqQklWpVrJW9kIJPEuZ5u1ZSQzBz7jWuR4nvF21x
M0ubd1DlGP1dpuD1vOYSqGUZY1iNvuzKrb+JO+E5Y+24XtmTEd3sF9quhUYgq/Rw
RrU48dSwx68oY8Xsur5Y0b4vh3XbUWQZo5o8bq6WJtGfbsKY61NUa2ufySo32tSg
z1I33Rh9bZBbEo7XdDi1y/RVoc9fZBUCMtY4VNlo9l4xC76dwbLbLIA8WKLZY3pu
/4IIA52+TL91AZYFqrJ2NWdDi5DpEXrUatA8BLBiKozSfZveAaHsaRu6B44ewwuP
GZN33dciJPkEaoEx37F/7vJTOd3D7qiPMMizMrJjJRb9FP5g7wDN8kdryFaAiWBB
nlLxeMqlr/L+u+FGHfraW7rwnb9M6Oqunr/8mgjHHn+KXwosCQsAEAmUq1FkDQZe
qiQ/n7kFYbC/UeSjreTosZubL6I8bHCehN1EJOEpwilkjEfgm/uVHKKdFD0fov6F
g2vbmPMlyElQzqUUUIBRV264Oz8NvHcXLoueW5M6N+j93ygjOu6NvE6C39itdkef
xCblYpa3zH1hutuYKYf0XYwZTVLSsJko+Mkf5WoCl+fnBJmna13tON9qaofSPf0U
X4pLi2sDdr5r7E4avGUbg2/nietDYs0imZ7qjeBj9lfMfWPqsirW+4HdgLVyKfvh
LLftdnR3llLgxI9xJA7/DUXwQV6GC8AmYQM7S7Ntt0PrUknYHviWgTtA6GP6BOpe
aurKmhI9MZUvjkDQpNE1slsNUfz2jXIUsXBt3uW9U+of96HO4PMsJV7QSNRZXFaL
zUEUddTTEKvY9p+sm37RJm5qIooeBfhZ2XcvGp49s75M22dUXSfcvqsVKNnKyhe+
qbQtDZVkerk10IWDgBsFx/UMw5bqsgeV3w1FwEnZmpocnO1U3IwE1WVeZ8OiDY+M
mD0d2R1EArpUXs/7OIyXKtnVLiDENY97y0lVtzvh5dpl79q16liQUQVEHvzuPBO4
O/XGoxHkZ+IlFkUX0oMO6SnkaahGxmXi5aZuRD7SRWwtLEfkztbYoRSRxEAtzPHn
EEqJAv4MshSN4YCOT/VdvKxU+X86cj54VhU2kq0hQr0xwTd7Jj0NKfB2SvA0tbmP
TSBM/R82Y4SfR4snsI5xMBqlm50lqwbXy5+3xJt8Qvpb0KvmUnk94x3jAasafvz1
7LMuOFqocL1G17OtBHmfvfCy7/XT+FZfwkHRsKiFNA2qgSesaL+SulXcL3+/abVj
cbR8q7xMYh9LekJG6TMNVIp9LivCHLijfZWNEVBrisCFTR6GZt8QzuRmSFJeWW2h
0UaSlCRgumroXtv/Z5KpqjYWGWAEHLcWbS9FhJE2ctjOGdG8N1qQApKR0d5zSkcv
JQSXY+j2o6ZK9elzuf3qD7lVFaEAfs+emaoXZ8KCLOpBwBeZhFn1yUodtq7Zm4Z3
fD9dNgSnLCkGeZBwHKTB9YyTX3m/ojWyqwJIeYre4wRzDMXjWbOhcAAXjjuY6d+D
fu5t1X0W/msl94CftKuCmn8omVK2Y0fc518NTGjzaiMxjCfSLkdxvMj68f0KYZG8
mxESykU5/yfsRceGc0rkjH4aoBJP1s4WMTVdVAXRWga6KYkOzhskzluOK6008BHU
qFuadyRKRNYp+CFIRa3q7/ylzTAsj6pTLZMByOrpjBdCCFS7AQUxuzGD8ZYcr/jF
ZSkjwiakomiol59ZesyZNsopgPQXrUPnenTnCwDv1OFaU2uh1PqXc689m4uv9YxL
RCaA2bNXCrzH9AMlxNs62ctO3BM4xCWwXov8rjB1h9wvT/KIn03o+RFveiNbHsDo
aOqaWXq0GvJiBbyEm9q2OwPQkGq+xxK8i0Zj1ZnCb63KQ6C9Q72nW/gp2U+9aQ6J
8kETY5oYHOr+ykcPq/HfRcOVm6Z84dgmW+hLG7KS8CJzWu+o1AgNbgrmwEXdX7+s
tHnqXCrOe0KoZ2ouJWJXVIpaOSdkMlSfvwbmNt1HO9xRsAUoYqmWm6c4RrGt3HP+
yhlH7qyBxu9rGIxozGgKmG5RmzxVpfCU9a9A9Ig7iQtmZB9DAf0oN+v20kraqAkU
XcGlVETxbr7brbaE1PfUprTLWmbuqTqnQ4cmdt/TC/UiNtyvRMNIwJoTMwKtMwKo
c6SqqehmQcP+Y5P+VZbvFCJuHxoojwU9i99FZTFUxSIu7S9Qi59XQ6H/24W2Q4kB
rCbs3xf8OELmwx9OdNj5mMgVYtKlJBK9rrSMGu1fql2he2UgDnLdcfrAatiQ/GRr
FgLkATEiXjRmU4cEefBZzyJswS2SFAMfVlcU2ojQrhQ1iOE1k2F1Pbngmg4CCjyq
0sTsAB0KNI6leBK3qgkhAwTRaIL6hyS7DTTjDDCreiI7ZQHoY37bWdHd0rpX/7Al
uSw6jzIwDlt1yYMfK6EGEamjIhnDbazH9n/zV+nKrlBSJSoRm4v49VFpgNP+Tx7e
RRESqFnUTR0xXzFzlblcJ9AnCk7QDlDMEyjwFCnxShwHcJrXX921KMlyP65ifjda
0JRBX/zPmgFZh/SI9JCoyplB0uSm+MKlsuXSQuH0eEqs5qaVh+z450K7CjEaJrgL
sSUqxnI2SIWDxkr42xA+z1uPrT1pYaHhgh99gIGtswfhYk17IxmBviZ5TJSoOcFi
fjsFChosHbxSCkTm1bA2R2HwNdJ1GaTT3LGhpi+D9yDCUrmVADUvkwc6NfVK2YNZ
fzqYWirG8oj8+KCWKFmwJHMtIFXVYICUxEaLBzW8jqhlX1+h0uw4eb5jKO+PZ1Sj
ZuxIs5B1P/nAaTOLrLqWE8Kv8PCItKkfKXjvkzaPwT8a+o/Es1uAWaawvNZIX6IO
U4xEMFwrTpgc5lcIySJqiCsRLlSctLT7+xOJlO/Y/Se1sgxhkWPzmDU2ojfl1/b9
L2D8DHFidiLV3CIcM/v9xuPlV4MNTnvlZK7+TlGwV1mGGEAQkP9VVrT80gv8hnAc
Q5GBS/RzPKzLoNLbR2trey15Ek5NwawjzO7a6oINzbjGDc7lXQSGowPRzBSpqoBC
88GYhUniiXpay3rMkoj/MrFrq5zGXj0LRJUTZznd6OHEy+ZG4C0PNXNqPQqZuWFz
mvuy5s6WVC5DVmZIwQozUoHR/yEXTftg4p8EaqouXywB5frgbv/tslALPE9vVEdk
3bL3FyLcU63IPeQIb8L25LKzlhB1SjL/O+YIU10u25/FP9v4E19QdYopAcM7rqYv
zxS42S255oV/v5dCFeaIw8mtYOWD861vipOrU7BXeHuAaBWluzxCJvARkiuan3S3
wg55udbDiMXhKWEp2ZF8U4jzK2xR5iVSK/eEoObn223ayvnUHZUTDlXvvBm+WeXm
LQrkRRfpTJO3C8zUBqVgNgn72Yd18V/h79roRAHhm6oWNXH6F1K/vXn5NWYW3YYa
zzzGoyK5SJrq1KxVK0LQqZAnAV5olQFAkmzartsIdY1k9i0sGzYejEb1Es3ws8x6
FIU1Dd7DgynPaNvDy0etzknP9xwnspVhGh5duTYymInODglZzMHXkwa9G9ZBomIX
nft9zxa1UTMJL9BAu/jb9uUUTHBMHS4NvEyTkpjf9+yl6OuaExF6FVx/D8+whOFo
mMO+eo+rGk7AMEJj7WzLmn0e4SXtpTHDkvg2MuFQPnvI5Yo87V8BKz3ihT1723/s
dYFYIIk8+HmIX43+O/qUU6BvmfKiXb7Z5juiW2nzEuHpuyc8gh/hHGuM2D0c1yf6
BuIk5bXR1t3IQn19boUNBZ7/NTQCcdQzLIJzdZhfQbDnrJLzTg2JUe9Ok07x6vwH
4cgS/8VNF/hMJl6DkrhEFTjcbkFQ6jec54Pn9qoVc3NFf+IKqAFc3BIejCbzXMTC
Qa2YeBcO7DvdiTIU4DpTFyVC2A3ySUJfCiDHBR7Biv+YpXu06HR7s/EAy+biIq0w
EtTGvSWtJpaoujwQ4zUfkM53tmB1Z2S4g3YZaHpYi6VZUS5jYPoPK7qj4IaEXyG5
qkVfnVBzZyuGbryxurIX9Cepx6uyt5qeTSqnwEl+QY1p1fGEXpvTfNRmnhBktf8w
OnJNV1xMBRYLeKKYt02X3cl+e4adW9bQxokHpMhDVq4J4hW+oJkYbSBgKdhDkSUA
PEZBzrmzUtKwl0UzeIOWHpEWP7gMV1sGoPr0bJOGnZrEPI/5BiCQX6i7NpdTi52R
b0JnrxkRE6H2v0AhrLoVr6C2oQCBcjxOrMI593wIxIT5TUmqQMUmOxzZqn/Lzswk
7qtTsITWxvTJuQ3V6AARGZ46QDQZk0kA85l2+PT5LnLXi6AGfnJWjDEtAi1mHTme
od3hlaDEgGDp4harj4okvw6GisLHCWr1Z88eeujzNp6d+LYZbzYZxxYjVP5PPFN+
7pErQU7b/KsF8s5MDE73BJq926q1MfTfmtrTGFKrNlJOvCAvINBtH7i4cuWM9dF/
qI2fVGO4n/kIRueLm5j8aKNShbzFcFL8/UL1pZi9/tmuO+H9rCgLy1EQHkK0FWTG
H7b/dR+QgwA0DqJUam8eWRUTJlK+kSN0fpVI1Nj3ZjesqU6HN0NiWefHsH+ZD5q9
p6v0m3jVTOu+IbMS37NpTLBUa2TOWHHPoCtdAhKokziGYkIV2YV4MSdnJAVibqeh
GoeZfW/DMEDu0kp4Tg0ICKqGgpdrr1SW8vjkVB63k3DfiL7RocE1EkmWzOxUvVDi
jB50W2P8kVL9OWCAv5BoKakHTn1LaHQLrypZzWIgEs9cZtImGBcQYktX5TeLVWmf
zJvPBQ4XMio8WoOcgb/MeO4sLRiSEFNCNCC2YKAbpMJrwvVKNO3qZiBXiFryB/+6
EC27NwKEpzFs/asxDBqPhjyGBdhnlSuXLzKlvXBjYtvZdOHbWRrlF31SGgbpvtup
8+BtDqidWNd36KrImNp/RMeBXAgBVXfa5HxCqvcf80YbRyaOGPbAJWe+rEGmzyPb
mqFbXEkvqU21p17nKqVoeXex56FD1HjXx4oXoRc1E9k5ZhibskJWNM1uttt7Fi9k
b4Y1zdTUtwg/jX0UNJ0KiOmanpJcu204elbh4BQ3rlRGoZ4wMemqAjWN9TOM7O1V
GP7G/qM7lKX8VMw9sr493uWWiRJMP+dwTCezzmxKhIbf59Hh2/IRyZmwYnEN5L/k
Fe1kuWFZVTl8THUWt2vt8slgwecnsnqRy81bGODGluzxRVrLyWvUIfuaGJ8QQBCc
AhG9Ua7tPLpd4ngAl6nMHiTxwsjqTahs0Q/wzO31XUqU4y6KGIk6+f9PW09n7W+q
ON52nwtsoLzmriNdDmSX+lVfWyeCeXk/pjpAKWGVHxVmMGXe3MEKOkWw2Wn39cyV
jM+WLZhy20htqY3e/+NBE0DsbExg3RZ3+td+0VId9S7jLMyduN1TTobEwWCPNCvw
c2F/cVleqDqcALnQfL8KFvh+1vMXz8O/k+ZoW1S4afk2LQkKqMdDHbA0a1Nt8vvc
azy+HVqxCnGUxmMLaFIflEkd1dIYKGAAfADnq+hwbOMVGbALGDuAyQZBqV1YCVUs
Ya5pd2H1yW/jdx+Q+tR0QqNr5/VqQS/s2I+8WCbFLgNPmn4bFxeTrq5MH0op/8hG
bHPXWUdmKZqp/Ag4PTVIhRohfkz68k6vGp7LursT9vCVpJrQqjWkGSoBZgCiJSDT
RnXnZwKiXal1ELohaqQz19xbFoKuftwOS34l4L9d1d1AwI3kwNMlLXwX1FXAUYfX
D2zQMRTO0EsTnkbfKM0EDmce9xuGB4hSFgIFEhwp+1S+3uXWGZz4NDuiBO7JlgiS
hXA3dLLlEks8mZeHq3nGDgUGMiRW4hND/Yy6poUXpzu7v3ekb6aLn61aaxb4USQ4
tIqsuubQdFnPZ3mXoDqiUb3tyDBQpu03qP+RFHsH7H0NbC49vhvc5dKoenIh4jyB
VpmO4Q0VGxWcYWrjJNnZWc9QEMLjk+Q8jEgZYkhI5OgIpCJfGSbgWHkxF3h4YO/g
ATQUAbl8LykvXCDuI4zTE+oPL5q3doX3cQ7kT/DTAwwWUECDQNcBSmlxZFF4JzC3
zEHGYCyeD3j5L7qDUZg7drFLVHf60ONi35LMruVx3qDoRGXdHydLYDC7+XlazFl9
RHaIHTGQK16179ctnLJmXYV7cHPZ36Au4CEVdctMB4GbQnTIUU9h+WK5rMRwGTAb
JORRIa5kQNjyVcrqukTwm6Ot509zXA3kP4QZbX4eQDs3E5d1rfloXCgqeLD+M9mn
06WVYjBaaDT+303kcvz8JAAUjwhhkwwbKLQ/AGBAOuVt7kmHhJ9qCfN4nShvQ8Uu
rMbWoq0gQufAoETITv8Yg0Nz/OO/i5DfQNnVs/1GvzwdKmuAswzaAbxJDjF9lQRq
5LogbQa+wqAuyU6YaaxNO3yOopOxpBcJo4S38Tjy854bUA4MrVSMtTM42jKqJAyn
KlZbwcgW/nN1KcSIOvXr0faR5OCyIM0mgG8LSr6i1RcX88ZuYqJx6aqI4yJDlVtc
pa9wRhewZ/SXpkNcse4QKfvHhj+694mmMLsNlzfebF9D91HyHhkZFEHbdaQcycQd
KxITdwmA9Q8CbfTwJOSxy9s7ifFNKIA/c3EV0OdTn5ZqWqifWI64g8IFsjube/RD
CdsLIvsaAgU9rncxawr1dAdgcihP8N3KTGMUdJCvR9wWFEF7nGhwUES0N0wt9/K+
cPfSO9q383U82Imvd4JGYE63JsDwVCKVhWABKIwmXsGXgc1+H2okwAmRsfkjnPEr
PFlR95N68RrOCIdcQp8irWLw+aH9909Xbm+7VG7r/ST0/rwho1xDwbJpl8FkhCnd
gX3FvSbClU18Q+Lkn+YHn3JWhAQ4RAQWXtMyyjwMMe3iO4npNirlTk7FRpg+1SX2
ZfSA5/JbAwNPhUb+wQbkPNX+YjlbNmCD83VF4rTZpAVBf2XYEdkr76qOYJV3AaDW
iyre78RGOAJSJil6d0TS42x+4iKtR+LsY2VnYBQyzZg2vi2/0DijJiVVGxifqfXx
LJgWwRa86PNggS6LoexrBjWzVaPsCoMZk5BYOh1TwnR/bd1tNMR+mPslFWeaL7nM
GLsYU3qpEGacqcNrxS9MS0XcAZT5x8mgQpwJqO+OYSAnPCbrJIV57JNIq08By/Zw
bMOnhEnZSct1cEvStJ6UxCJLeCRglCS98/99nbOYVdHaF4iImz8m5JULKe0LRIVt
bO5T5cvXHsGH30vPhvCbxG1rrDT7vMWKl88HBSIgJHSGWvMBMml073hlr6eB4qgU
bFEshFx/1TVVYWA9q3sh+V0GODlMnClqrSBZn81biwvTcxIX6V9Gi7r9RvsxsZ2O
ezAt9DK6LzC/TPkuQ+yCpq41oI1jwkZxnpXkNAaYq1UfDfFqNa3brynm1gWiR7+f
G87eTLPVGGwYJMbz00k2t5wUgYLtlYMkPU/7usCGwlM59jonGnE3uQx5Aal1fWDg
JaiFi+lSZtorlEykoqURZnmXsN5SiEGMPWgO5JKeB3kUZW6DQqux2+O3D0fjQP+b
DdC4obO6nvTGuyoaXbvvBBYFklPouXR0ocDt+WPu4qtF+zVOVyUV8dSjpuNSfZ2W
h69LYIj0LHw+dOsoLDi+oc3UyY7wSbt82IW/jLC6TyPvFu9EQn5aRomLgFj7oOHW
h4xBk9bovHRLqWbv/z13pr1T7yzWnuJCZISBd6QleCDRe4ZrJVQV/RxGhwt2zMey
sFDUn39X95mU+A5ZrMED1v213LR4oz89tSKu92O+kTVP+mlqCufFrpxu2qSgMXVB
2CTjMAQcqJzjq2KSoJ638PnsXMdWWWYzI6noKk1sCrQJqmL10EFBYZV0JTrS/g9D
5Pia3LoCuBrLAHkZZdOiIFQ0IJDNb1BKtPploZgu/6T/RFBc3o4kJwbUPn+TwZ5j
+6yNx6Q0Aqr3pKKQpgAscmyA0FaZPjPmMgMsOp2QhySLvWP2r9QpsijGxixUq1Ms
uyu64yMujmSSBwNrE4nNkRki3N6CZbUK5rIYB3xzEEyElF0oO7ffJ7mgNHDsDK4F
mbyWtDpZofXd9efd+vcQc1xIghDop/fRJAj2YFx6paqJrUoRFA2e75TjMvziBSgv
TiJBLRFAgcZbtfSGdA/MTCpjt+YqZQum+vlt0tRxmw3rCantqPfiCl4GBDaBmH2B
kkf4e++dS//boZF16I1e1oac+xDJtOBxb2iTrPt3pv/L3J0iamBnE5AElDQpL6ui
TjQuvIqsFbeuOBAnxNHO68fMRTX89SSPfjUhZ5ZpA0xtNqn7db0UaYC46fqYKZbB
KOhSZrgBosA8bi52dLAW0fScdCMZoc//YohOwd5560jZIvP2sWOy5KO5Sgh8st5V
UPCaaMhyan3U925RtKF5YGGqgukN2DF4Hp5ZDbhD3fEsHLPJ+VgBUFicD5sFupSi
qSxIoeiEbdDwc068Wx8AxIG81+HimgoRL0+ODxg3s6wS8cPd54wYsoI7sHDKr8RI
ofuEnIz/q3T+Oz7ygVL7QANWj6GgGrAh4rDmAfpgc3v6h9P/AQRITQ9psds6+YE+
kjG3AcYqt0pbfnKSqf5/fpDCxAq7OIRwOlnQ1X2UcCF1KBPo3H/N8fOvPBTqr3UD
CLO/CH+OQt3Zkhys3b1qRLNWklBrykLPhV4z0KYKVr2XkAHniDLgJgOMxCLO446F
X3jcVPrznvRkvULiTGPvWShNR4pjsdzwVOyxkJ0CRrbKFmtUWAKpg7SRXmoAb7Md
XmZzkgO2cqddT0AA6jM/piwkU1/GMtolTNcfhkk6svDSHVt3qEn7D+tH9Ztohu0Q
WKBS8RpBZo/nKr7XGScRVd3fgg/7+jMoHHEcBavZK6ZXzIaPkhhARGHx3XXTSg21
EN5Tv/rXsGWO2qxDk9EWJkdLh4OuX9GcTILoRv5JFdix80WTnqRAl7s+eL2RuOsX
AnskaCsUAleoKO+LXfE2Es+crVQITK1oL9D5dKCgZTHPcQUBRwZTnCM4rbHm+7TM
uY1pMCJRumpwqVSiDaDBwHd7ff0MbnoJ1dVcXV20MUuFWUbMTZfEaAg4CMCkFDrx
O26V6UVqopiD4h8Q1N97TAcn9hao/vNQ+3Ei4AUcDajtCSHcsCuNbBaeuEdWoNjO
PMHqpslzL8r36IuDSB6XrWQTeDuTsuln7Xp/eO5xF7JvLA33Tt2uHLRCIMJgbszh
Cpjrt8Pzq0JZnNh+jgIGIfZMGCfxP3hbgjtYnxLYb0Woa7po03Xgw7aSW6G6eQEa
aUZX/8dNE0piBg94hN+4lT5ixP2iFSmLyrkrHp4GquqOfcn/d2ohTDQVzwIlxf4R
FmRVIeqiZ9T05kEBFUY9YjhYteOEp5xAG40uaB6xwKTL8mCWWrQ2S2YFWbAqSxwE
Llv2sN8B5rmjipQI7atJoO68zvFual1kHh0yilPjAXasL79fqTdWEJk+mbSypK7W
npygKhX6H5xv+faE3M23G8B/25X5FR60Md5hkJSInu4MQTxDSeC0M++ZmRalpxUA
+qyYeIczhcwKzGH3MEMdXxetUGPlJFxdwynYr/GYijNzLev0dv6CyxYlvV1OUx+q
oXnJE63u6NqITwZqHJqVuRX+ISwJ8+gbEPDmaUaz4bU6BYj81Clbz4zy0gWdAnO9
wNSHC3SbioMpESuSpT0mjmnMFGUhyXPLlB/UMGwWK/e7nSaDFTKQQM9mD3gH06wW
vxOP28UD3EuH+P2eF5ZE4ENW1MFnsJViYUAOF9iopJWNPFGf0MPSkddgXe+XKFCN
gzupddmDqXca4q3VfbSfE/GFHLxMSMSe6PE8ASXINzLgnr9mCyBEXeE9UZVF92Gz
TuRS4nJx/iIgWPMQ9o++QuT+TGbKyQYiZvLsljZxEeosPoTMtPKFkYMLOCvIT+Ha
U5kyAtexHwh16goBBhFFzHpTarx5sdYenVdfukQsnUW413jDKtTtHq7sG8hK7Hvg
+i2RwPwlCye1eEjfJHN228fPmjzPZXmc9ZFjylbH0T1+XVjy8I6LMXWL4k7ZJ8Yp
6LvZNIsPE/s7yLSPtk3JfmXMlnvYDF8IRyipLpmn4qHn8z8qioDrLpIzO12azXeE
YWz5QYOcSXhQlr9s/d3pF+dTISqE6/VFgITGhwjdkCa8ALcPFQYR/ZwHVbjahinL
Xypqt6LrpnGZR8Inyjd1R3le2rMPtb00bEfHIzqni3U=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
B5n/0CroiCpcBeA9Ox4b3oX2kAhUCl4BEb9LYttrY/eUoAPlCiwqNizRFPIdoZm1
hUGZ1p2pwyGDDsgqBuhQVB03Qri81vSNDJms1m+3ZAgJhz3n45lnyB+vUT+ecLFQ
Lbmw3sfVnCbyIVlaAglSq++66vl0yTdMyPNYjb5HT6dtIadSkIsCXtrfmPFh4ipm
JzlRQf2OEDWP+ibAKgx6MLKIqlr3GmnYm5ZDTIss6/1GSHkBYoMkeFYHIE/ar+sq
/GoDe7otrf6WNJihVvP8pFqF4g/0AhpC2ivmL6vgVUB0mGbiutYtzAUN+9JlasBx
aDfybUcHz09kkxfPRJ9QMQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
Qz43hwq4qeXaBfAhIZ0Dw5IL4hWcv6q0mdJKIQ9bqdQBZ+shthkdk90vIX4I+vwS
p1louSTa5Bi4BQKEdNtYPDLnIXT5X1LyEHXuZyRLIpAf+djpL/3Kvzs61XwRfZHe
wVVHNZaWWvcCDzVJEQp7Av2ofebBdzPBdLiXjMc8ifUoruynir621Z4jFlOTOVOz
PeRsFXV+rnADE+VJG27uSgt6yu8xIjBtWKK7WglE08v8g6wXtyy7+7Cvw/1WjmRR
lkY4DWZ6u/LglLchxFC4GDlPDq1FfVga/geHiRXaLQ1ZesvVq1r0adwLo9sqZe2Y
/vMT7RnW+9vJnSET1cqV4Yux88ckO5bGKffcz8rgLd52J8ZvY5NWwa+TuoaTwvqb
7LaFFZDWQRexhywB3d0UNAC/JQOhyG+Qp++TuNCAG+9SjCEXk00Ojc68LADBg+OI
8/A8gqdvq8t9EaXkyNCtnT92OO+MBl94/ItHB/ZIy25zteh2AWMHaEWS20kMjKNr
9E2RAA6QEYjIwiFezw6UQgQ8cfSDFay05u34H5cJJXfsjtGI6e35nd9Dt5lpxKdX
/7FYt5WstAxMMioZcOYOpp0PwzBmDTG77uqYidgLOEvePMZumOrb3y4Q/f1KfrJR
feV2AwgjdtGQsN4X3RR57Mo48I53UgO4Y8hp8ZGSLamrZKWdHNIjg1dsa4odVqpe
MrqIgq6YZnmz39il2wITKZAPinbtlPj83xZH3d8cq7uTYysoAaBKXbJLv/teB+WY
89RH/Xj7avfGwHRZskmUrNVcuhtsDxJB+2Jm7Ct9Q4+iy/soUeu8nUjd1OXN3hYM
LI/OJTTUFBbb1nlJmCXPAhPnN0fJfrfRzjGuqzcN29w/wdahnVd8I3/7NXVXz1yq
rL5SiYT4EbH76jDf7plHqrhBasww1j6yJAzXKsKldDzswmQaTFSnT0RciwsURcHd
VDcjSORKtxGM2x9sUD2KDA+kJQy9m8AiMp21JE53bM/qUm95qNudfLs84UNDB+Nq
0ddXf8S9rHfsCVs6lqB9SiXZULIUb+fDnfkgRv7oZkyO/aMZQq43r7PIqcB2Dqji
ecHvn1YpgWx1tdtKGUmv5e688urBb7mQy8uq50txNFHzkjVoIlUGeMlyJQU6frW+
8b3xR3cRZwzAKBolBMgI5545jb0oidhHDDhdBR8m59vsXAlUfT9BQo6LLBxjrKRZ
K8O5RcUrBSRbb808p74FAj9AIyE7eOZlbhHOLEc34FeFtYDuPsaX8l571qG+hFpP
byjSZVDII/TeTnTlFcbyw1n2s0pwt3iGVo4yIy8OctaxRkLvZRiXFhvVHWYDojPR
RZ0dgKdW25gXofsEX7FvRveQH0bvn7hYCZNfBCRYhFtAJoLQv21yabmIQPxUsFIU
4QwTtQ83vGMcRjjftp2gWNeH0x7EqWeH0cGlBWjrV59cwlYQ3a8EDPGEGCZAEPw+
IKpwuwwZiwHKG3QX9pRKfrRyXKR+grfD8/PREpu/SuViCcy4W8O+OnTmgN4R/5Nu
b4tJdn5RDDpYRd9y2jg5maoxxSTSx4EAk7mqUpIiaTqtoaNzL6jhMoL/7SJ4vL5G
lp1bpIKL8y5JsefLleIB8+/66esebbeZ8HhttDeNnLbJxdofeWjSPqxwfU2t8yea
oZabHFbMZZJvOx6Z9R5gVNxnhmMBdWzyy6MW5GMFUzDQFQZDGSkLyR8W5uKIuNuL
urY/yNVHpoqCYXQw/dT2LUO3BfkZPPQIHMQLZYGplLjlkt/cXmlxKZv7eLducAD/
gpemgVSKCGSij+TMCiGXZ7DJg2dejUo8euI5F1aSrTjFR19Yi6WoSSyx4cZz9bq1
vW0rvA0hr1dH1O2I4w/rOlT554tMBubFz9LUz1cLjqAEe+9KIajtdTPgTyQAsC0W
Y9QQhBOYn7NkMaXqeUpJMn4FrScDP/r2zGRZY/7wzcllaW9fqODwlDoT60QeB1i3
xrW0kw4B28k2S8FBRsbrnr0dmUQerfreD9JaN3GNw7z6Gbt6ET9GnsLSRTU5fsge
n17DYAhXKkMrDADgJ+rvdHnA8GJBlgzDviXOEYwJJDgoJ8GJagimeJDs6M9NS0Dj
cLz6NId5rd+iwvd56F6vfCK7y6edlmk6p6FhspgchTz3Q0bLaAQGyTC4lObZvPYa
KhOKMzAOQ8kZJVsCTNejsHpnVh5gWeRr8BbKHQk8m3guolDBUJqz06X1iBxx+ka/
ii4pPJ6I9n+NBuzw0mJzsAbBVQYJDs487/9izKX31HDC+Xnew5bQsITBqCBdSZub
898di6LotQYJHSYmnhSv56wVZBWyi5KnpkyAzwAkvAzFI9H4csZk8Tntu3ItfynX
FGjvrBCGebQhIRyaAjYPgunBzyb6hDTkLdUNDSHS3/fajlHKdGu/Ioms4LbWKvGj
Aw5GgKg3brYkJOqcP73ObmWrxQV3Y843ceG4Ct04bVjRcoGcdouOoW16Gqr5z3Yd
GNQPiRYKcLvLqf8Bc+OmbwWrLoHfKGn/hqknirvC6HhPn+avGP/JYnkWom/CnFBB
R8lc5CE/q/nxTz0yp1YAdwNpaRiqoLpUMBgCscczbVwBMWdqYPXeQDwFUqJrdpN6
z5YIsWvcytcsXEbOtJ75QFEl4i3P+GddbFBGy0Gg6KllmRTa23dFvYf2bLsqKdpr
b4UcDfXzAbDWXiyCPtSHXe011fusYFEGU2/BInEPBBZb5TWQJbtwHYKbIh+OpNBV
mAX50lAV851CJ6BoNmkKozho5fex/bFtt7KtZXyvz54AUr8q0cOpM5MDlRjy+mhh
P6M/PFGnmD5Zb6/s9VZZCn64al1oE8BiFElOkQ8AOn7OlKrtytAp3ZKK3aNrmQwe
udv+X4DsDZyuZ/km41nyRPzhLthSggO8yopbVHhTVRdEUIy/dbQSn2/D5Mk509Z0
xzDo0s+IUgGIrRIuRu3aSqDDG72cNC79aY1kPsF2rigOBRJr1wpLQXdSlifoFm1V
Y5klrjgtdzj4Xi8HsBv23y6whdRKXQcqfgCQkNj5n1SpBiMf1BaW32i4Tj58LxA+
iuaxIt8KKQhH/ICHtxSgfjI1VuFPVR1ERKSzl7GZVG6ceeQJxrUuoW0Ykb00knZJ
YcoNni9/v8l1dWtiuTWFT+w7QL53QHOxsMwL74b56cxqImQ0/vCE31+5DmrfEfTg
vemOXd/XXCDvfSG9JWIOWfFX4EbrEtkoZrz1+meGQ2hgZDy7ymB6ez43fBw3TblW
3NRKWGt1U1UNNuaKK1h2YSH5HC91cuiyekgJ3dki6BhraHP4gNEqteACbQKZk6rw
dJciiOnoIpoIefczFSNUQKitfx7GoS+T+XNbI6d8INWavN/HXnnuOk2QDMG7Plty
cSAt+u1+rLTy9vstqzx8XrrP1O/IAS7cXQyE/uzXYg67SnD1WdI6HfGxjDG8nBA/
goq2Icjetp5YblAIXfUDPxay6nYnPd6b8K4O6n48hb6MWAwZCbeLfOD4rFkRrKzA
FYiv2UQpHq8qij3+FkzIAqihPcmYnYQlQY2eVWnZLLDV6fr2gqdMo0hwOLH/wKJp
tAwAb36cXbMIjpZvYuZcRywFKwg2j5tb35LlbOaUQVVcEt9//PCDdE5oa1n0NVog
0zbjSeRoTILZ1yKzFu6RGBJlQgVdJ2jbu6gkINOpGKjz0TxCpm+EvVjedJNREIz0
/k7SdopM8PJbdi5dpNIXRvHZphd9yyUqequOI0uxcbINiNlNi4eOwKHcS6Y93LFc
LiLP/RzRa2sOqd5PuOZeqMFouthNagSoCgx/Sm0HoGiGQs2C87hD72QUSFhNjAcE
gOlEzhTGiAJ9LksihPeLypittHgWLNKnaKmU5D5Xd2EXwSRiVnz+fAtElvTYTIPb
gFBZl2YYv3sag2SkyZeCCH9V14xDcvKShp5K1hDyyXS2wg4Xqwstz8Ixubs7cjR7
eUZpl3rwKFewAEIvXGZJBr3hV/7CFdbOyl89TriMw3EsEvPA6FTFE9SE/CsUsqXj
IHoe6wTD2fdhwMvEnh3GU1yf/v9v2KbXnYtPIu+H357UBEe8MrdvDRPxzGP7u/Yx
wrbsTzRdj4YZpxoc/QJPOu04sRuVa1SVZMm9Yj9Ns6792eA3iiyGnIh1yOiICDMT
05nvFUYkK307Jp17ZySsJ4nqJ2zOoWdY+RvFlkZxPvvSi0HWd0yrAePanKXNOb9I
gfJNp0cIOvQxvZa5kgWlLdsFG9WdenqFuiFhiV5GBMbXBdv9b3e3t0W8ylcCYNB2
dfJcKpI5/k7McL6LvxB9zq5M/Net12DQFyNOcPWytkpA1Akv5ij1YtJa0vqTsT2P
dW6lt2eiMh8w0tkrBY1r6twdu5XOxFgLWjdf6J9yuNGvFxwsxn0SGoSLwhUfWLeE
BRkPQm0SXkD07UznmQBkJ3f1k4BCQywbNPe4p8Ys3mVxhE0Vo0ZygreLL5XsNPdN
OQQ+9Cz4jAhXsLRux+b9B7/OX+g17db6lIUMWX79425SMI154rg8ghdGdZEPfw8S
9p3CcYYMoDBJTk7qlZRNMgiKrgc+l9UfucxHVXu0AaS9h/vujmN9BabU+99PEtEK
QnEgRb2vpfiqlYtf4PbGEsvE4SzHigMXBLubfAJZJChOWYI7z7CYIi8QiUAUI0Z5
GfjrtQwJ0vx6weDZrceG4O3Z6eKoVX8YDxXWpr2Eyc9SnIWn0N68MbgS2gYdhRz5
W2u9g2FtMNbLh9vqU+qT0LMUx1+B+obw/Tsmdh08/o5l98d4XGYu3EfbrHckxRHf
sc7TZqJpXv6obuALCpWq7Az1GSWjxByvNGmEOKqLcM+wZyVIEZF02BBj/OJRaqRb
VCDALwReiw568g8VHswGyJkW5lKpbGKY2wu1ZYaSKHaaO6cPtkp3MNq003JV+AHb
ibVM0iZsJEZx7qcdKpe/l+utIsVZmQiPaiPC2xAgw69Ed9xnK0pcbd/wHh3Cu2Uj
lXhsqxKaZXtPf6/6v+BkTH5FhTdNwW4Jq1KtO/XGMV/DM1luDv6o7WunjaV+k9Vm
jwE9reSSY6s4O+AnDzqUoHEE7lD3BhTnUh9wEYDNwqqqFUUAAZ5vkRb3eVagHDyh
3xu9P31M0AI9IoKNUKf7t8/v7DdQQf1BCYyp/vmH+lo=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ebxc8pw+mMrmMNhdBF+iadBIKJe8aL837jJxi2vm3nBy2ONRKUo55nMDtjYeG747
uzyJvW0RsM486Lzl2sF1cbnzSnI+fu83PEkE7vE6l7swBb7hSp/XTU7Rm2mtNuXG
JraY+fUqZbaVt/G1HuUa+0OVl53JXpZtKVxoL42gOI20Q8kkY1rtLyEM3dPYLFPO
yE8APyZisaYk0eW0GoXD5pPwrLZlfSPUQe/KogZzF2mcfE8Zr0gNkVt8YyetJrXS
roSTPHb6qMLKxsLNPHKNZefHAZTaFbqHF/pm/5pRDFscRfz5V2gf2s2F78i6Zfix
0PTEfB1PZrcsr6vMIKp6MQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
71hh599liXYULCyPeaLKd2ZImhHnKD5ewnP/TCVG6c5T0QdXhXIIvFD1vYq7PkGw
qt7BeIfRpQpDYmCBG0XW2bxvTzYSdGA5kkIBtLWw1ghs5JTggsTQvKdoF14NP63e
pminp8cNWFqgfcrDtgbDo9H4eDDt4JNvavAHF/fEMprrGbFUXv7OOFmH3zxvpQJn
R2NhQ13RqKEz/ROpUpW1JvUZYrUYoZxKI78IYHLItFjRQFVNFfFpXEBApcgvLyoj
GNdcAmJcVA8CFpGArtRTZ0cawrFbzNAxzltWaia/PhALF0jzvkgawNNgQ08Hbxzw
yINqkWoPtjjrkEmrTjlSdPLJmGod1XQs0fVslXFg7Jmsf3DCOk/NX8n70hbEwkHd
oSYrP/oNnrqa60ShaNT9Ggs2x/C+WEh9sD3ZBY2YKMa2xQKcxPpzFlP0DQWNZK3X
dyuBA8ooJBL87bBrPO67AeN1bqYZ+k3emSRmDeRrEoawhPb8ygTQ6nSpWEMLm1M3
GDPnmheIwoLdh1w0x8hqXELDyoUnqfPBoGSmmKqEDPwFkT90ZPVAZI+bj+2h6hql
DhOaf6hMVGABo1nt+eydSsh6mkkEJkVp9EIYyvjvATLd//5p7AW80OqS3IqEaUFe
6xIBMNy4u4eGZj4vxdy/1VQOlSapXisveFVr/oAYRx4VKaB5oOF7q5iylCnGRQ3A
PoktyjXC4R8oMZxXlskZXIdvs8umi6OlA4IYKyQmap/m/lx+UlYzNgkH0da0tAL4
3RRLDaf4frjvJpoNcjvMmnbOejImc+2meHqiuHY+VZ+yerwW2oZm8Y5Lx88LnSiK
F0FK+JT4sRmgJs0oI+7AFyxJwoPzI8f4xoulub7k01y/6bsFF4OXPGVP+FWE9uHS
8PksOYksoEoK6dqrRySNV1SHjYSYHjcsae/h+yAONTjvt3c0sTIrfn0jvEd6uDbh
iXsNOE19TPEF09qyqCG0w4D+vcpr2XxcpxmY1eJbxOseUnbjljRziE97TPRvnKXE
+ZW2uhT2YPrXF56xes1mWLwu3DX8vrtXsylWsH5sh0FeQK1E8+MAb9v31NWqi48i
VaZihWl5IlPs/Jfi+073Jd8XOoR/451waUQOom6BI5rQ5pgWVMcnhfhoZAYLcmGl
xKRgbGAU7Q7lGToIXkJXYVGb3QkGJnxhddcb+MCCLDscM/T1dE7EKMYNLRf8qDs1
c28rJhCVbIm1OHuiYFkDTHri9P8F//mNerHJ+Bent40eZb/2qAyUWb2HA/PtcF+v
zoyrJO+25ExphvJgA2vfClsVimzawpeHfviv3lC+7AxxmyJ/t0AWF6UncxblhAPd
3b6N6ddNzasxizdkFUJxNUZ0ojwUJAXgXO6H/sRoeX4QB7CnHs/EhQ741i9+w5K+
6mIzOjfbpe1OuQ1V3GzrKS3ntuMW6y4GAorhP3lf7q/aPwq91DCdLPiekNNsX2ou
WVCeo0+znLjpp9m+6+89ULAwTN6bhgl6XS6Ab26nrTLhT7EICchowVkHgb4rMA8I
V2vwHtPYZWyeZKjM4B2XheVmBKh8oQdEcY3uE4ogEPZBLBYvR00A0jVXnN/oZ7kU
mBDCXvx/y8lrIoV9dlPo4RXRpfX/UAKM10IoNQasvRp7/YqZPPo9IHco/TfhpusE
vunUgNa6JyWjK93cUzHssijLQVm13zrXZZJ2i5UAVvlyMenCGF7aj97/3q7Xluag
Tm2+L6xwiNthI5bpb9mpgp4WGPZo27jSbisk5VeBdc3EwNyljU462odE1VKabjqK
cZGrl3RpceBuwi8AqSmtZq/MHfgKsjyIgOrXOn7PjAj6GXhydd5HVZxhiYZbZNUG
eiwzl/FhxJoPEE1xJHjXcyR6NocB8Oi9crsjCOUHdb7fluPGDs78uWe7Tnhzmf2a
dbutVQH1R6+h1F/UMVPzOBY8cT3p70uvDwgEqhon9fTfWbxFIAULNDUYHGPk+T0I
lHoLz5LU4B8ytC+X9Wdjvn8jFd2uAdZikTmoGF9E/Gbb8OjJXJrRA0bwfMQbW9fi
sNv77A6PTKYF35+l2SlXXl1mySq1XQioKpSL/z7mm/a7UelwOwWFd+QjppCAsyfi
KhkZ0M+IUg88SXkeJr2I20crH5YwpPJUPO6L4Pfhib2IDRK2yR3xxxXQJyic6B0w
UVhA43uf7d27PkMOOv557/Svrw4ctwpgCf0gX6tV9xum/VkMpKVPUxDDn2xnzFO0
u4Oei7M3HhrTMYZz6MFN3HyqikDhBP7qj8cRBlpld+WUg0TOlW6ij8sUF0p0lArc
hvKDKxCftvY+xsUmNLCKd83KC+HdI5RLaCjASfVLhztpnGw8mnyLz6LzsJi0k+UW
O1Zird6AlEg4aRz3IFnTR/EQGpoU+xJLj5lyOYdekQ9rIggTBJhNPnE+ji5yKKPZ
RB4C/qzzK3GwRULRr7XVjnJjjqGpk2Fw5NIwVpg+nvYa+j4iivbG64YlRi5bLxO/
NF5jdoEaIhud8wtXgOh7tXq4badv4wS9FAX+Z+c63+MIX3/uI3e/ZAfUCtkjNmOc
WRn5ihfiwfsEN7M3aMwhvgnc0PQRH+TOY8wbDduB2B6KskwL7k6owhnFlT77YTiM
218o5+rzBr2Z/d5/RtHCbbwmo8HbFHWE4nsBuaBTrCDU2CFXtOYDSWiQYH6P50lJ
RDPJyenu4hHjPxGoeEVYBwycyVQj8qQZ77gSWfhlwbFkwpCMxjx0ixXXaUG/qF8Z
QzP9CpJ0K1Y4G335sYoDiG3Xo1BRGU6TysNnIArrxGXcXjpRJ6p/nNTA65pd3zG/
dbJqCiszUDnzft/bzMB7/Gi2JOlNEVCEm/phfz6jKM2tkucaQgEoS46Q2k4SfpIA
luAl5gYGSZ/TVmpkm/ZvJUlsMlFSGV5GhPOq3fTVizB2zC3f9yMhDS2Gokf2cmZc
J+XeT6Lu/0x8h6MZeaMRM0JveG6eksIf9OvKarJ+XLpuBPKHYw2K7WmicOKyhVGY
SnRagArqGZjkj26TtI9CJDqCUzR9n4z4HpRN9+WzvjTKkBc+OvWEbPavQwppVbKR
phSN/c19VXDQMX8CUz8+8yVAXbfYj6xqI5RKO6oM0TWSVlCet/NRGCTu3GXNeAyy
PnE5/w9FduqmOUUt1zbE2kTPmPU6qpkcDvx7uzfrMScqBdLYl+ThVWEuX/Z1lWnY
PeDXDmY55ZYuwjbpIpM+ru4SepJisrcIflCS+wWpxIgT2Us4L8c7ztULMeKhQtFi
z/vxa3OGFmREGBBoQLRKmA/zr1bGzflDC73uXaF9cY4iPTa0juqQr0PAk1SlVGIM
SfhOg2v02wqyuVNjUEcOvc7Gw4uSBzNsF4WMElHcoKFO1dqNlGONbD44MTnKq0Ay
wUy49GI0wbjPDsEJX4Vy1RuJS3StMsClRtopEyFaGDSZGMAZzDJKACvpFsp8NnNK
zVmrmIqGeZ2axEW7aTDWXqPeQvT8L/aBgWuywaA7nqLSYzll9TPajrzmRpIdArOv
RvdTbwQSNDgPwFkYxtFYeuGLcUENyo5P8wJLjgmSdr3RedmLBJ8i/pn8BJzqywfJ
ddtuXMhtWQsH2RjchwSAWA3umse7herNzgzUFBWi9vnouVF/41KSltThax/U2/Sy
fMJG17QfXqnyxCEc9VPiPakF2zS7WsGiyF/MVqOBlX8AlS6nswq9OMZocphoJBz4
ZHP2GrdMtqtxddpSX7L8+fMfe/Ek7HaiAx2m+WcHr9vKlnPrzau/oAWeAJDZ+prJ
w8p0cB9m4aG1wg6XwZyQcZyqn4AIk1oQ61dNOFDY1orlb6eGE2FbfLO3Kfxs3sZG
gCFNp2BMpMHID8/c+DepOAVUWU3sV0E9Wfr3VKCBxK5QroOO18pXL9Jy04CMejv6
bsJDHT9N+W/yaBmarxD4mDByTsnLO8WlZ4bT7dzJjAothHRzPZFw9QW5X4YmedNs
YH3Ej/IxxxFTkWRMZ3hbdlCO6ysHMdan0FbtP0nHo2qjmjznLSv292As6upxMIBD
G9UBdFDeQlzWjQ91UKVUNJUCwjWyX5k+qjqScVw/oVvu2LS16I6GvrYz/LHOMFzG
G1ZoJvAfQDWpaG5CjVyTkBKU4MDi/UcPQNrIhQjdHvdokm6dX1fg0cXEVgSljNMj
IZJK9Dod2FRTbp9pGAPEH7oJgPRGLBzRKkr8XW0ec2kiKcW4Q95QiHOz9OOpYpTb
NO6EDhPlVOuQ/qmokxxr4sAEokTAu67rXP/+J8aPmhzSKj8poEG9cFnS6CyWoTg7
YVbcUYF/EdMIRBpMwHENb417HOXPqVvs/RjgVoX2dnq4f8Cd6MWOg/FKwLuwTOg1
Z6fdMZcz8oTdtB9wPtV9LnoXSaTOEldjm6GK/k1tAIbxeMUnJM/1ypvmKR6a4TMx
AgNjVgxUVRi+PiELT+qcq4Qe9d6vk/mCCxPXlKhHuum92lciSeBVGIbWd9IanyND
rsDh3BumxRu2iB+7sIblpZfFYpsFG19R+r5Gw8Zvb1Bd7W56DaefHiL4xhmBaAt4
C4LchPyssnAiB3MvPnFwJPN8ccuHuOPHJ8btxAPPnLWG3Lrn01c7y9iPjvuYh9+e
t8SFtuBkRCZV5C2450nLOPYjKX3mOtrCgLuaiScLKS+VYCL2tIgl23Epk/Dr+k9o
Nfm9/DfF7r6etwi1xyAUdKtd9aAV4/MKXXJiwhj/fyq/6PO/49xRHOZlWiPrqnGC
MeZmUY6Swvmnc0MqiwC+2Or17d8e2FGUmt+YjtyQaEarGcEmHzztfJoJMuBSnBNR
J21EyPY7kKGy4wVWeHTA++xVyQiDZP7fqe1YrD/72PkHCo+NIKICbvvjIgV3Ku3R
FxVKisNmF2UCJsSybGwrzumkI4tbxV8lU5RRUfqaFvwFmoBfCMJoLI7953eSNaIJ
qrgpQlhUlQuh4i1LqEd3O/t0c11kiFy7fV7IrfOn878zYmHx6wVs9Tf3fYw014lb
ya3yohAXlZJ+njNwdP3yypoFXhhm/2TNhrbW5SRoOQ7/5VPkTuC/l7/GfztaJApP
7A34/89wRP2H4gAiF23SxXa5dJAbYXe6a2YhxrOqqfoE2h0dCmeZQ1WqKNiy5h+T
v9NDnVIx3njtDY3skC5tpTwxwCkvHfAI4sz7nkyjhssFvPDQEtkoWhiyjqVUotvk
GJNke/08at+3Idl/iGJeJo7XX2aFAXm1rw7uVHJns6V54FNiaCVAnqImrk5MQwlh
I6PhODXapPNDCdrInx/7Y1oTCLOA0HkVr4cUS8RAfo2sihk6uUTxpl+SoHV9h/GV
dgqLis77ibq3uai2s72BUd4RWNqYrO0hZlaQ7az1w8uGEHAHWc5xCyJPBCjzUDwd
DdeFsgQWsxPemDYKbYrQmYug7dR5YrOF4laTWEouAcLNVOK6uFO1buSnSvL4A14u
mrndYQyiwF8CFAMCB5IDc+KHLwBFLRlRfPqQz1o2aB6bKArWX6TCAoKFtwhRE5WF
LHBSAZctwRj/0/EmRyhXXizoRXkbjDJ5O9O8Kzca+bLx8mOQOpMMHNqa3K3/mty1
tW1bAfkmy6euSVX8ijQLJBthUSoc5gP/4PeX2rWjQNlft6U522VLM0X5tV9xs7VY
Etl5wfkAN638fb13gNZLSSJYNaGGf0H4d+a+glOkYC0yvSs7GKBVtv2aEaCkQ0s3
Eyo+qAiW84elSqWv9bKLNfAqGxmBsblzJcpc1+2YPVoyHznNg+0JO0ZTULQ7+3/w
6/7U6yqw3xyCetXTy3mBcvRdzaD971hTfcBt7pBTxXfpOFwPz20Cq56U0GJ/0kC5
H3oqvfCHVgzlUGszKd6LzWKgXLza5HQFBuBo9OHz4WIYyiZyK0iTmfmuVauk+HqQ
CuLuZmdn/i+z7eur2/r5AtsC9hB7jqbJOxXXfegx97pKJ4D3nSzRRxRPBDBkGsqL
yXUTqBm1sJn79PpmnxJWsx1R7AywxkevHNZ77RLDCZNEgAjdp3WgWRZVsYCxq3vn
9fAGoHuGxZ7xQS/O/YvdBfA6l0+jdlwQ25NmrVL37GORKqX+4Erk5qAOdcYymIMI
eFPt1fT6Pe7Jsp2cyOU1aNF6avILw4HaPO5uQmz3oyJgjtNQ78NsX4cfOSS4w8mX
7rhsl1519tgXRiQ2h4ZC2vdqgtWu1WYegUIwFZx3NaNREsrH4HcaoTvbRSueQRtz
orFAPjYcbR48/+abUmzE0t+HPHSYWVibOyGbBrfLgV45uFawZ3se+2wxtNouJjFC
mhxXF3pCDnmXdd9F4gyObqiAlVp4Gir8F/YZ9BjubaMmWvmolAKQScrcfrowAk56
hOmnszJyo5T7WnIOqJmNp0mIqHi6JS2R8lCfq63CmypCOpYEPt58J2gDdwENNFzm
Od0E+OtofgjaWJmdIwBJuEWpX9cqmrS/qbJ7luOlTGbEriAsjnYpP5IUn0E+VVyu
edR6jNvUjqa8Vpy14C5lrJ5D4TQ3u16nrLB+4QbN2Elsl2GdBIRsQZhCEVTKTLyW
rOMcywBiG8Zh4jKoWFWaVfbUL86Gy1cEgs9yMOMkkQo7O2TbUht6PNEZ8uRFdGIF
aLq4zu/uRZqzDDqRvgWTWVCeJoOUlQJyoHjlERJTA2VdfTCS8dEYE+Pdtu19Y1HW
llwTLhdezxEvuoCvBQmYYZKV/v0bLwq6XXp5TXtbkaZSkDfkx24wlyrLGDp923MO
cRwKvYfck4soRCnA8ndqjcZpZ7vNoV3mEOmJ67DnJxZh4SkLCVni6b02fmyGTo9R
CZgDJc88LhwqZLrwVmk9urpHaOVZ5yeyiVMOTKuz/PbpzIwJstCUYovLvro5fLrC
SaE2Ta+xohl6Q3Ri/DpxPEVGpG1cO4YpVkmSCaouhO7OrBVEaEHerJtK3/TwSSrH
5xRc5wyvrKaCIjipOQDqwbaU/ibS55YCKnJuE9SGLqfhvzrjdjVcmEDfUpEZ9CO9
VGesJXquWMf2OZ5qGhYUL2PBIqVMtauePCz4spoty1e6S/Ky2bdLme9H8lxV7mft
ms/QCqrQGG54ODuPgThj6PZVsG0j2sMhSr8EOoET4SH/2PUyefAI8S0AsALt9woC
B0Pce/cG3P0Dmf0oxS4/FnfAGfSLfOLxNTVjNrng3La6jVFCtuGzQtx9Y2SlQuQC
FFMMjmyrAU73OgaW8CNrhg2b09P5jGMDSh0EkiG58RD1kfIsEb2VCtXWvyRojXMm
qtuIGwPic4YP+yTnD0B12/VeHIrjcLlC/rcQGV4o/IIggbYJPfL3zc4asFjxeHhx
q5zujKZ/RbVihF7Bu/DmbJmWLoq2Lsw2DZJaCJjwX3XoAtEwNU95fmL1p+2JJ0xs
q53bMBYLYmr54lWdJjjkBpVoLWJbCe4mcwDK2tunVVBMutokzw+lMjS1RTZ4Hcp5
1bxI5ioR3uKS4tMm+n1prRZwmh4ioUMY9JoLxfJxALD9RZ8iezEUClp1FvICT8DB
j+xGu7Sm+dFrxITF9/t7gTykktd1TGbCF+Bru2wEM7YPZhX3j+eWNhy/FhrjevMA
85kIAnq3cQFyNAlEzfDtYtRVnFIBtEl4aiQEaFZkwPqSXyrx8X0zpRJVU3E4+dCk
QqfEzTtA2jdfckbASRmvzxqcWDNqYFOim5x9zeuuRVzWqYFFHn45vn7Zi5Ugw/6m
KmOl6x9XsohDhbYVNNLwhO5mlwbjDgOzq/btDHYUzKIuB0KwNcOdMteFb3zW+I7/
9t3Whp3QuZ1Loo2UORtN6HQ4JwBZOWF2fNptWSsutkctURuSF4AxbMNL/98Xk5of
vZZQkiwcVe4qrNyXvx3pAEv32kRxRBlVanR40X8POrBn6s5By5gQ4XuZa7dyNhWZ
vYaiEuF8eqWr6gTTiS2PclPC3PKjmNX2akycdx5+6/7Be3dcVZ4UDSppjwUfZxY0
lb0vVQQkNM4czVsNsATR7+EFl0vsIUHa+OBiU2VVYxbUL8MkjR46XpUXbxdbIHSW
1lYq8/hsex8jCY6PCQGjGTleb3+fz9rhhnlP+odVdA2dN1EvhBJbzlGXw4DKvbzg
gYbqAANSglaAeD6DdqX3FprBQApiwZ0N5CmNj83M6clUH/JbmA+6AlLnH3ohzH+I
dcOdZkVOtKiKR4Df4HdvQz+N754wMI3zM8Qfiq+ROuIdUgsaD1J/2pFm0K+Zbz5A
7EqMG+9r8l0htbvoLPDf7rjy4NqLt+i200l0aWkGtye4du68ztmViqevNU9OJsiS
LeRYRPdz3kj/gwX1RinoXxc5a+A4hmsBTDlWMXMUANfrCbnyULDIX1kKlwvNochJ
E5cXB9SigMG0+b/UtaxjyKr7ieNx1Frw5VrY5CKBDihrfWW/EiUH/UyinCVsBwdB
4leOHfUqxxmLs7AtfCABR/3IXzcHOJRawcOC/cGc7ErC3MK7pCQJluiEHasU8Tu4
nm3oc71xG3NkrZxAkQSrpJ7wUftwxEjfvdRcbcKYEmuNotO4Y7hToPRsrzHr9qCg
PLaWU4jlnY/N/EkZcWUwjg16rlH0Hg0+bTB8og32KcQaZqbbKEmAtctiOq6NoERS
jph4U6FevXcDz89+KlGaBqrI1qGBIRrLAX2MBVxn1zm7UD16HsdNvzhEfaVuxzuu
Dm0wiWJ2H5+y/pu+vwCNNoGanrm/AVlg1jvZCT/+IaVcJCFBKH5NtvwuUylOz+tu
Q3ymqMAXZulah8EOpMw733zIueH4Pi9nnMktpytPZMbVdmXZRfPAlh/VpFSi8s0U
blVG7TbZWDsgr4pEKiLDlbGn35TzboWQpvxveu305LavzbjR3fpfSI7WdZQzvY3r
M2RM3qfqC1QDcyQrwa3hZgy+0/P9GKKU/4/hcGxBR1G+atSgPlBbVMlKrB46UNlQ
VDns4mNWSX0BlMo4XR2DcW8kBncQhDJaHT5dMza6mLgwj94c9x3RcksRwWGYZIzK
AaGEvNh/0BA6KXQ9tFmW54FUQVFwaixmkMQmKguVe8Tw0ZBNg3/HOe+rL013t328
x2uCvoeryoveH+R3PdXFc6qyjsjrg1NpCybEAeBN+u2uqfyzhphCKOOPJaAq/OQM
ZoOAJTMdAmtMiLNhTvp2H7PL0k4BjyeJySm1IGQnnC65aSUubnxKfpog7DgyEbbV
SqEwKsyG5s5vKlnIUCJFjosFnRHPzzRzB1c2A3XXJmczw0afXV4DLBE5CxHoILQl
R1Q6sGBvwzYtmvnUnaFVSitRONJwdlD4woepi5yXZQ1Rg226cUJy2MNfoMBZbxZr
ce8XI4wauH0Wjg972n9Nqq3MW+aNSnQWFFwpCDF5RmptpcrpqvRthjbDeprHle68
LMCeUrwRhyn+23+RQKxxKnAqnKWBahKfDlbQwTI76jxEdNXS8fuNe59TA7b+1kgh
eBKCyxot8tSRRP4RHeg0AB8L+2RX5/rhu4W3+ITiWBZo4yNHBQRl1fDt/q4WYCmd
UBhosYUlaM7ua3kdYdq7uT7sLN6yRZg5jJ6Qv5zbSjZ9T9aJqUhwz6rlP8B+BSuC
vMpxeGbXAGTuDP7UEZ+YoncWNtxlJ3H6PxMXB63Ugt+UdzkMc3pOKAMqAFfschb4
M4Rgvdr8BPVovHfIHnjdoNlhRoO1J62b6MKxqN5lebQSQdrcq+IVjIhYymWF/fix
XwLDgY7gWku9Z0apE/eut5DgZssIlg7aIQoGuqmWXupTQLm0KAnoumYGQuNdKaFS
IbjcS7m1xTrgV49/aVGQ3FOFCMcVC3pQrtj8R15sZmGFUVJf8/EJEg/hBQwtM532
6LrOwFeN+ZIGEIZdqsmvVpE6iv8AaVX70eL7pRLVCyKmrKnuVTHi1r/k+4LXeMUF
mP88v285hdgcVJboocHja14xMrbWSM0UpsN1zLQU9Ct18qV7yZ3I7gZErsEaNocQ
SIgMgd/6TFS7rbse2rwCku41EBLo9uxHN5HCs0SbRTrcURJHs4BNgTOBehinQ0tp
fYkHII1PfX4cqSXpQRSOSnQAYdYzF8TIlctYhoARxa8ULyc2OZgf7BqrrRFW823J
V9ShbP32GcRA8d4EFoIJXp/QP8uGkQhIL6jWox6eyNecJ7GX38jNY9qw4pqw4+eN
AUfwvDBXykmbHlnI2trzmemNjYrNemfZSYEoqntZGtQRtvFYGtObVo1GvMzWthG/
ydgZNiq+/bPGutAIFY6F/LGoEaRv1eLUT9z62VcL8QRrgg8+x8PHAsaCdsPxFebC
Og/L8VHvTAfLWuTwe3/SJ0wdrqmz8A4lAGitv9PfVfLuILpeZJARaXq56JwGts+2
8yeHYrPcKOQXi+VG0VUt5Qy5/zAgbrkDk+59l0NsmWfusbCT5B4zwwCmCzcxPQeh
MIiHsTIL2vSbuDa2yWmpdqpn5p8E5MmTDfLS1YyZXOIxMszbr8mmR76XnaEokUVG
iGLAu1MJdMR2TkXvigoyS8fPapI+aimsMJr/EN4T3Hk1Y2tO6fzQdqqqJ7JXPJEQ
hKp0DGFeK2avB789cSxmdbhIHJvddSr0R93vkoEGmGhHgkIzYQ+I5/c3e5ixA/k4
gm/DiuOT+HRgWJRHADg06IYaYFsA3LpdRm/XwXP/ghrnq5/MEbDrmso2++kmtkXM
BTp2mh4L4OITyNRhZg9k9rAEVbQyLxUtWJW607c8MIApK/MzEN9Fay917yjCETeZ
PhwyUL2s6ehgeHcEaQ61vXN+ZoptwTAqpKbS12owEAJaTqJxXDnfVimmgqhmYVV0
3oZ69D3XFfVlfWAMqL4zstWTBQICgySyxGYsxogsLjYIkb1RgYkD4ODSioYpcg+O
ATU9JIth1iZ2ufChn3lQXhY3sO806OJWCaK9pzFybM93IOJm4/rnXOJlS3jDGUxr
jVXQxdHXY5P4eeEUYfKufCb5jPEjd0mz5iygYDjeiLuwX3AENUW2aZzMbXS06VQp
q6jIpqr7NerqkRyS8RluiIwIpuh+sZRGItrqNqR1oJY/DEy51Jf6LxDNW+jDQ4+D
yVJ6DifQ0Y8W07ulV2GpjQFJ8gk9Z/xbFsBdOunm105cGNxQpKmnEzecZSsDr9xV
ct1YAFJq73rbPywoIbbx/IRJJsWL/lr3yS5yHQ8ytBXdsgHBcvyYRvAt7IT46y6U
zLnUqHocLjA+bm/1znW4PQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
br+llBlV+3AOMZmuS4EMLFwbgh004x4lLj1DRSJ916IRWLXQdP0dtCzT3l592MBE
xv4HzJ049ZsbIDjWe/0HLJCkhMnGeCooKsXa/7LLKukGk4T64BSb9Wsd/M3A0D/G
bL/Zq/ji0jfeBllqciev1muv+5LlaHVdkFIc/5xNTYJl8Nh4ypQXPpUw2pYtrMI2
7VzOGTukI6Itf0ICwgSddqd2ALn5iNPbLkMOWw/nSf1pM7+qOrDWIefUKpBqQiuX
DQVkgkbu0+S7/oOIIpmuHVpJs+Qdu0YdzLLME6iZUqPesucJO3vQqFpQMg549DUM
VIHJyoVwc8H+wJY/0vEbfA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10640 )
`pragma protect data_block
l24EELemxCO18p2WF8Y3dQ6RA204sU3H/tJTR0IanMWtKYB1RzCoWMTipK0ctqVs
lcZv0/ElYv1PP5Tsx9AlqKAffkEHD1C8rtgADR1S1q3fjxaOoUuT1tWSBJVRZYNU
tUP/PKDlil8WxMnQHqOd12eMECpot2A2eMNGWcY3Q5cYKI19rVuciyGDI9okhm1Y
j2sgXyvCf3VDCCWupH4EbANOsCG/UsOvSXpDGgYrs60oOcnB62+3sSz8QOuukwfg
Jzj0BaVA+zliumRwdulqVsBH1Ah2/KCXZSA6mn2IwphPBaGPsqdCvGzdip//xGgx
SYnWg/5Yo3gWUmvAuHck3foHxQ/71tKGrtQH4QJxGwSSTBXNajavYhpQTIctR0t9
9g9xokLHkUUYkFqoatzutL9DYaqJj55N1UvygEeLEYHYtD38kdUSJ3TbrhLt1X3d
SHY8nk/uehV8LHyJkJcLDNaBfb4zA9wFcc/oqjym0a2ZVInVcqP20qArnPjtK4ct
hDl/OkxFT8TiL2mZNl7rRfdzwz+zUTaQHliy8+th9OfsfQPx5xd5tdJMoLCiKqWq
pGNTcnjHfFmE32n0OUO3YY3PmWXjYYH/AM0H6lp7aqPaCXK4GVfpf/rPv+zTZMvl
3W8Yt8IGYFa7SWck9ucZKY0I0YE5noDHF+WoMWSd/vwQ9jHiVQUf8h8dPyNYnula
nDhN36MdC/1tiFLFUxHdEy4ZSz1xkSyBO72+mgshgE32OxyZC/GYKU6mNWegIsVz
RbzQkv4iSJ3DKxwjw5reFPkuKCL5jq4xM5P7UWBJH+jieCcE5NjRcVwFnIS20MXS
L/hbXUerf7AtFjLbuZu236YN9HhI/XiWDgXbsxHH2OXaGzJRht1qIzLL7AfHIvaB
OSc/1TyUyKZH/9QL0iWeW0p0v5/SrfF5Kq2QNkHAqL6HqQC60SpmhCbbBuRKOZ3F
dTiPp67TNF//PeGi/vGWs/ZPc1p/ompsACD91P0SQ+llVCMyUB3lkJnZRO+mfzGs
3OC4ebYfuPHi45KdVUb9+Yp1cFKw86MFdjJvl9uOB6oF7aY0NXpOc/Hnf779sDbm
JzpVOZZn4Z5vhpUXCNhdxRxz7aG8i3vnm9FlhhNhs0qygKnrHRBUzYfDFYWxoA5j
dQaebtQEivA/yhrh1k4O+nhkSRh0pdJbo/3DgGFmgHsXMGomlh37FtC6roYpGPXS
WnhNapElFpi+wd2Z6IRDNK6At3KTX51Aa9Hm0O3cZbShXGzy5Czv8cQC/mi5Jsgt
kkGvQ8xJtNrPTAOsVtGazxMpJ0oC4gu4kSx4jDAXN6ndWwTigEvLhHoiov08AnYo
pDa+gBkWI/ZrFVu25mdV7I0BlWW5FcAguiFIlpaehlKrhJmn5IxVg5k0ZbPprVJL
3XV8gWrIIu0Maa8D5r0wLxnHyGrplO0S0eeY1cr66U3NgzjM/iCA+krZdfdJgI0S
1GCdfRX3apmD9quteS61+1qUZHUpDxfM2XN1fTZI5mK3VQPNHBtncG+cClHjx/t2
wL9y12fbcq2Voq8AD2kAtozWBoAzDewQhEec+9nQFUqKOnpLDVFZDgprPwGWRTzd
9UggQgKRbSivv7favBy/3x3cKbuK+DtQhTPwLOsLE1CxoMyng54fX+VKSodBEafn
mGBBaREYncG5Nrlgkw7Rw+l63KuicV7RRabm/e2rhJ0ETh2jNuKi7e2G2O1/DH0A
2nTx25ii4NNW1lok20HeH4twu8I4sN4KplEBEEDp4kWf4gnRc2J19ihEtkwiWDeu
u8gigdUMVTVRfjXWzoiLL7LmQEcxASv54nOWZKYV+t/KKzrJhUVQ86UycH3pjC2K
ZBfd6tQfJT0OHaKoJCPsiX5Q9kLut1LE5p0+ocXeclV7KXgkBJtOei8OxvdskJRK
32FJ5qZ/VuHpy05AJL/QWZAxzCKFShaJgrHJ43ekypMWNRiAYi7H1ByVDL74vQjR
xXsrL47+sunuJPNR+RuYwEHlrH8oq3Y1poyNvF62+ZYkzGz8PciUpysE3tfrcVL5
OxiV+9qaMViu2ZzAfOz7J9kw8hn8mzzsBkuOVvVG0S1Y4K5YI1jUelNKFJjgxEPT
Xnm+TbsEc1Yu3VB6As62yOyWw+bslJZWTTOBxmMMM6JvAjJD5jZxQRjna3benMq1
LtGyf5NSl706ud+2Yp56utV9OIdx4HopMVqtOM/OR4bVSCOiUiaKohdLlp5sbAxM
7/b3T4r+LYJ9ExDwHm0pomiypnoXd/utqQvwsQRIUVkMOZ9YXpCSB3w69teHJVxN
ybGlTEavdg2ghZgdBfDNkypQiHtlsI+JXz8onSEJDCB6bRdtIQE0qO4Ip8BA7AFy
XxT1wMqvdkrdIlqyf+xkrdfsjsEthzOP4Fv4HS4mXIyNpyKe6GD0hSK2Xsd9ZHjd
GA4vBztC/X8Hlq1wCUg0t6bytOX1YJDCATaLARtSgZ0AZ0An3CEkUu562lLx+nqW
ZC2iHTC9nJVQXqC6m7VHpilZH5oeeL0GdllNAnMEvkA9mheEWHQnFdag5Cn5sXuj
Ho+6cACdXqGTHOUHYHWckpKzQKnaoN2LAX3Vizp0c7/zendax3D5fPdx3HFMWzOc
24tDlXsAFdjwJSjfkkPyH16m1cOY5yOhVSsCathBDvM3vkr5lzRXIQ9HR7SjF6Wo
eQAErOeM8G3AyHaQAc5pKIC/duwXleB2XPgbUlEsUj/+1+1oB04QvmIoV5ivFyB7
aVCm3oQGFDlkh45V7i//m/07SMRaWcHU5FrmF8qPLgteKdBASzXbPbgzB0DK3Vpg
OVK4bqoac4+aD2+1KvnICU5LSfrwTGnkgr+EyDCpHuVbMPM2LNAhG/MsY8K0JI/+
0uzpV8YXc268kqwtlmYZ2qIEilpsoZp5MD930u+7F85kJR7RkeRU7mjhB5YKHcav
ftc7o67KM/k5eyoBP0Cka8oWROlJIbmMpIuuzRJ2OzsRGe42cF7sVCHZzzgHnpgf
sQJMwO/cyWHnmfFGqUGfTcBsQUG6/PYT0iH2re4DYQ+r8Swpkt3M3CPfbOu4Eich
9wIdNfZ9yHIOvCbF7XUTc/+eI9feqey01vPN0tS8dBuV2JViximUz3p7QKqEFXOq
J3SL7s+0k2KSj7sDx6/cD49K8ypcu/S1ooFgQLUhmwufgDyAZBqWcKyd7CK6eHVr
I3xlSSveVX4pHOw5WOxGnX5Qi4Skiq/yXVLR+vLYmDZzaAEz4b7y23nXfL2XFk3P
1mCYRIcPJ1uds+xp/bdZRW4pvWZvQUuhqq8yDCxlV9DY2548FZNsUZ9rixqZ3LQq
OMndrXukeoVRk0lKMzkHMTyK7PquVMc6kudVSHahAnPCtx5nrr7NG3Y/1gLm3mFN
3J2u1nBmYuyGwCTUpPNZtiZwFEE0tyDo+SqfhtBBcUNvXJ5by19U5t4RriJgCEzM
Odbz5EW0Wr93+zf7aJL9XJ9ejgVuYwpVtaJoR+Mp9+EsPe+mR/Ipw+UIq+GqFIQ3
jk9eXwtblo/O1EUhbNV2MOt12RMy/Qq0eZjG2lcu8KPF8ZGvmrR3eCCt0xHD/XEp
sEK8Wfk7xmdWpq2tHWmL1jtHlk4JVkqGuP2p8g2YF91HnFskK8nF38K/5SnqqTrp
PR768XqZE/YJirXWa9DAvBF1ezRrUt5uibwU6CtYBEovJiYQqBi1jLEnGNjUbSix
WOFHoKOal9u2YHt4lGLvOYIpoDa4Dhk2Cpb9yr2zsvXJ2yU2BextZtlwti+ka47c
sdqBcDV7edvVAwXFBZul0PYRoKb2s0yfsixCjR8CISYxkN0qQz3vtzJKg8n2Svzc
vAY08BsppWBxR5kgLBXvkONYguubJPjx2OLAZQv3b7b+7d9O016th3mIPOKw4IFK
jxiYJ7suSQtVom/x7jOrlYVQmlhVWINRMU0HW4QAwKXpDaVkWma/wFAMpEiagNYt
FrsGHmNqaccpe8eJ85sk97/qfhjUr0kvesPW+4JbvS/OHLAfplhJlz4qW6inz7ix
lt4r8imA7pJzCJiX8rgQyDZnEI2fr24aMW26Vm8gtPu99pGfTA0nBpu/lH8G8T3j
A33vxF7WRaSYK/CLLgvUuziWPLalvm1dCfbmzi3aqfEE6hk04j/bz2DmmbpXajbd
o+asDm6QoAwxXIn/8Ofpzzhq8ecL5GwvLAwdWuQJqQA61tEqiF92mbE9cSYJtye0
WXKU5byCX3MbqRye/pmWJeOc5+tmwCHhyNfBv40oY+9EuQmd5qPfnwrMVPyihx3o
5zAjbANLRtp2Xu9PMYl2Cmkcfz6lzVf0BN589V9+rytk5Xn2uPb9A89SJRRwJM1+
jx+6gTIhFNw1RPhzgPS51SFeJFMtS2k+RT9q9UDqq6tZZa6op7lpHdIa+wFPPuFU
aC1nd9rorkrQtiJTDlBMQOX0F7eURRfOmeG1/P1NieJdw8ooHjB/k+Wj3weuUn+I
3GgCGeNWc3PHnUgrvq5+VQ9/xHODpb5Nwt4N3PvcPcZM6DBvu6v6aynbfZ1AbPsF
brT/l1jzbt3aL6fS10+amWI6I7ghrIIi0bleBtRaH1G77vraZwmPqPsq520vnbWi
H1mWc6U3Mxc4MWd9HaWaxWA2esVn0hevO+o8R7VKp9xuG5f8Pjs4OeYNzKQhXvsh
i4IOWxV3Zal8Ao2b3ZHaEzpuqC/b+Wj8KAlSOhprVeKX5ZewE8PKvD1Unjnh70SE
KlzzPp+ZmxFHzCgA/clOeVyQK0fA+lb9KghDwzYebUOWLcNpoqJBoAhBNPnNHe8Z
HRsMNKNijJdbpw21TjwzqE2bzDvecOhPofaFADZ8qV8TZyWkWzmo6ebTUEkK/QYS
DXG48mTjVBOPWemRh+q812I35YM17cTIS2cqS04K7rudNLgcugM2pqqdYM7RlBXR
6R+v6RPbrVttVHqjFbQw4CAoM7/RNodfbX/dpIom0AvtLA+u/0o38U2s0/hm/pe8
nTA2lEmdfurHDOCzNYbgTJ1zQtNYbnmYyG8pe6+rbtiy/INeuGZr2ZbYf1tXjT8l
4Jxq+9RMwVPJG42WbNjNtwFQ2Nvq5m+I6gC7kVHK6t3lqdePJLnD1C4N49voKDuL
42mQN6KO8dr9iVWOsYnc9Qc2HrVAOEQ3sgtbwTTflRamHyQHpvfokaW4Ji4BEhpE
duc4HfXhHrkntWUf3wPmLbXCOg8B3LOvSvRQQP9/sQiBAjbt2Z8fUOlXnIfYMMYm
kjObn4OzHIh41/YMek2wYvce5/M5yxgaom+Nb0L4nrEgpSTvpcfzuPNP1zC6etJR
qsN4Puh3TUurZir+NdbkTGAWh2PO+JNA30ysBKrVKC+b5npwbaXURAydqmKBkDSB
4cr+L8y9+FphfuAmMTK+QFkNHgbOkQnyZNwzNsgKSv0Dxiq+dwF6/w9ciQrRfHkm
VKPFDH2kbhHWLK9V+AR1Zr02mXMjEVQKi9+DYrtKSJrbnfY3dUh7ykL341Eut7JS
fpfW2sZQkQkXMAIw2Uuza+++w2D+hFwb0Z+d/3i11LmdLI5+N1mj4pr+je8wSeto
2eTrJ2af8Zj40Grds2Thx7oVdU9cWsSdHYa4+yTBxEcskKB+8HS0+VaoVSY//x1C
wPPrXWLE4IO8TVm/WeHp1wNrtT9KvuVmdq/khOgs9UBOm0J5bDv3P5vVOzZ8+/0v
VPOzGgAjifXTqo6o1xuIGSllNDp7IEvi8xJNUs9nmI0/HmaSYMpsvsnOkAVG5DZj
8xvJlr2l9+cq6/owuklridsiHikwRbDCW6mMsZFC7SmezN1Ti5jh6GX4APXjOfBh
CuPuzT1J+BZUsi6k0JCjT7BcOvIHU4i1WVE3QsoCHGPN5f77HxVD7ZIy4yqIfM81
8n6qb4NmsS2Shv6DyB0tIwNWF5/kCrfsmutMreOeng5ad3xGV1TCNC7CREyQpCvt
w01sxD3EyMvztKYH58NfX+kNO/a+AHDedowok4glgq5gu51k/+HQG14M8fck7AVo
J3bheoZwVTAeomxpne8vKZB85iDNw7si+Jk88K4mU50j5A9wMVGOu788zuA8o436
LWKqGfro8lquNXeNC8RK3ogEOnWnTwv7LQEP86tPZ6+zwAm1SEViP0qHZk+Qk4ZP
DlmoEF+PoX1bqkb4hEcQk12ioUaHdvnkevpgq30HCzBB41g8QCb0ztc2NrhPoRLp
DqjB4GLVqW4I28jfBAJIvbgDWmwQ1Nai+eeslayJQuOyyicWYex41QOk1KBeaMU6
kHX+HOx3PlWmOlxkcksSuiBgwGdMw2CJ0xz49/J7bHZt8cQU/ZY+vA2AwHQQbJkk
a32kjT9ejisjMB2hESHxmlOoH8yYluzx8ZiQwauZiu9k6NdfmWHyk6xxHsc/SI/z
KjvfSxgbYA1kagZewVNeZv/jxsuHf0ovLnR5IKK0E2llnHuGJK9qmO80DGtndLmM
oAFy3XT8D2Fx/b/tfR0AKwCaSGa85jfDffHxwmXNMBTItFzsTb4QoZliDOoDc2xi
ccF1mp4ekSKlDhNCdhZttLBe5458ALtHHOPpGWyhkFhgFyKK0vE6R7VBwsjQSiOi
g38hXqUNoUCn15dCIGvV5l5FlMfAP3csEEgRkndFTxATsYAPdHwegbFXyajxs3uZ
UATeX5+sQiYOet+GkLRQ4DJrxHWE3ejr7MdY8C5vJNeUALEl6Mo8Ngr7X5UJpcSs
fIpYUzBlt8oxHiHBs4ZKT7j7orqC/LbwYhslv6VznWF6bDz8A/uXqi+AnkpfeI7f
VaySsd3qpmb6x1cSU72FU3gPiD7pGNJ9b32R7G6X0GpCpPx9WgMYSLa2ZxpuRvhg
00h20ZqjI/P1CtSNt/UeeRoNGX9aFQdDY4dJtBzF2iPREZL+y+UVEVxSExIdJOXC
eX/4O3mvnCGDZ5s0C47ZclMCnjet6xx02Pj+YpW1UdotnsFYv+qLt2/0b99OFH9q
hRXbdTGwrgjnUJK1/hOUCrkHR7AfY1SMllgc6Hvd2Dg+++ilIYQfd91Rpw4LSmzF
db2dWdSZk+u218W/xi8IdCU4gGo1+Tj1kJku/v290zngEr83hvXtq1vlHH52TzdY
rUuBkSU+Z4ZOYc2IGy/8mIVSBbLgdlkSktRBUpe4zGPqQ7x6FfosMc5DzCs+b4c2
jiDfJUTfI2gS4Y5OsmTKa4nnUPh6itxFdNupaTJZd6D8XiNcov4/MdwodqbQAk92
EAkxvSDKoWe8pgVFf5elhhWku8xGwPju2DgT2LYqmA1lwe+WpEH6qS75oD0yipCn
8gajI8abSg2rKhivcPtB/JquuFi33HRxa1xqqza47YiQxLZ8xhDQLyoV30RMc2ZP
IjZhwg3xqTxc7/CMoQRhfc3JgCdSzwD4r8fKVjel54S08XgYwzEaGl2cPfWgtQHl
nIHe4a/FVLjL8uj8VP8jDNpUlo74rdOLJQ8yCrLsSzLLUZ0PRRYmY/ej0L+p3cik
PboivqvdcsCRlAFWOGVBHqoNYSoxkciQV6jnlc3DYRMJfLrCz/Q7VgBzYAfDuQhK
f9dAdPGO4bVsGJ1j82UAHv715v4KUYReXVc0tnkBpL2ZHL3S8sQ7tEuEwpS5rdSF
h55fExu44yAUSNgcIykOU6dJK+IfX4ovJPl7BtoZPxHg0FtVOWDFns01gX9MKK0U
00Bco9URv36BrHJZSEqw3Bu97f50Cq97UAUVnb/GZ70hfRCBMPBK+yNm42jC2/Eh
vxKEIyJAH5m0oHbFKkNa6OfihTySVRaWc1OY4K9q9cM4l1PpDFfQra2C2PKyOMwd
pT3pvvTHtFNHQ2LZEpL9mIBhHx+eWFXsQk4Kh55YgD2/PQQb1y37uS19DkM3LKrs
1s1fnHOetowoE1Ci/Z0tTycNkV3SaZvXcU7Qzxp+x0ZfVe84h2IoMOWGu64cDLDn
Ccr7Zm/IVcrEt+iAGmFnC7xvFVvk4Kj7B1YBiStphPo9WEC3OacQAVbHnwM3NHBC
YJyIJ06IroGdJQk1GxddlxjCPLqvaUkrJu649MRtiN1Cj5TF8NytA0vas8Gga1b+
PwDwJ3NMTsMTtdanUQ+EBQs05KWED2MxP5t+3cJeBIf/N0c4Rn/fZkKTdgsVwgQN
q5DgXBzow+lDBvcpDprZfiRDg1QQGlECdDX1DPTb5yickrDaQtkpvVCzxuxvXka3
iCprnyo9nRBE2D+1bCanxKrOeAf72CknVNJdQ0xmgJUWiUNxMTImDm9YZzFy8efT
SP93PJMpDRKnztY7ByzCnd1zUIMSq4nYDTipppdVb+oS6kiWXvDlPjLOr3yjLSZI
XrX3Reswsp3LtBu0gApNZo8yg/l+EHhiVdZm41iHjpdD5SzTkTvvrTLKXZa6G1bs
ig24d8KzXDHo/PYruJdIAqmZ0lvf2bQ00uv7s9kTLbCBKXrIRgPEbgSoWbOXLOUk
PpNFTn8CLHFMCpQmWmvb0BmFjK871Me747B9QDk2vkGn11bY9Go/+hr374sZkN+S
/I9Zuy/gccIJOzZST6bkZcvyg3hZ8skDwGBze9Gr1LiNZxhoBtfV9/wJvRfE+DgT
G9bJahtTvUfYgwCAN51D9dKBZ+IhEVtjGdeyN/zkjCE6jNXyJzI6O2WFtoWLVwY7
2H9rWdjKHoTgst2glts32keqigUmgOFQx46hsh6yILOkQAO9QTe+6twy84/Uqz5l
5n4j405k7kmuFNob4rESvUMMYgIZkzwVtHJrB4BMdiBawuymj8wCAZ2b05deLcE7
DJTt2sIfQkqswQPzKqzODDzi3gKhA+n7GblCJA1i8wOWsBABqGX5fTl2gNrK+FXO
m5KEDiulXn2zCbRb0V1nnsX5gJQwhWUOy9F9GfVh51x4Uy0WBUh/fU/ryithGLk8
wv/KhjbvGp0O55tAjbSACEFS9WK2sYIfbWruSSCA6WSgenaJWzxg9e0MBK+EWvOG
6bNkRHyTj44yUipt7edt6rJ5eVCEilm2bh9nk04R1Es4Fm0lG5A4wRbJm6J3ZfID
3YbxTF/JVScMM1HUBCgdIgKsDqCW6y+NTB1946XXxEb/hD64rj+stG8MD9ugWsv6
wtTlBZusJ1449QBlZ0DtwPNIbjujHSSh/jzoIeptjTWQg4RAynNtHhlcziQWURsc
BAonQcK/GsMBavpq8P3IF8XPyiqHTIRBxAUUfETmzsY1gFzlSI4jqQiczxSRr0A1
+Tjnu/c1oa5DNVaeQZYgacApY+Y6ZoXl2J1Ah0Zaw9PnMDR9VurFE3lBUYeY2tzw
Ab1k/6llZpTenzJ3z7xwJAsBdhCV2GC3bxvh65I+FVqjsaWM/Q1W2p1mH4hj9+st
y5SlaW7mia9g92yr+BhsBEFpTqkbpB9E+crSDQV00n/o/gybsN3g1+9gbB7VycRs
PR6Q5lkk7ODWXWehKHO8DFTx8Txsk1EmvO5GudFOMCDmZClyV1esF8yppLl9Q4VV
VNff9zJhdvqAZaJoD6V+T5iqyR4sN2zOkZhaLzgHdeOKWIhHi5zAMmQ23RM5pR++
Vx3GUWyforTODVkwtONpy9riNoyW74xOhEQ5g5H4/SYk/QI8NEhLOLeqn0C7mo4m
OXpJjpzphr9Y+A01DJH0eK6jtQRzWB6vWN2/Ee2G34duq8F3nbrx0z6hyJFIpU+Z
Va1ZTjxlZq82IuBJesStrwmGjCoVy8Zlo+3WpaYkPTztZlHRdAfLD4Gig5fqZY26
QEvXkHQ59zypTik6ulNS6TmwdjFR9f1MVC5US7O/o/25mD4jcjo2mOhMYr6qxwl7
rMMBqNd1+Hn72dJ77TSNGifH88is9ytObq3o81WyVBKlsPM+xZ9uuTPtuzqHCYh6
NQn0ConmzwN1XF6jJbi/Yw4ut3WkrEy5NslsfAiZmGU7b0UPNJlksjbWEWaxeoXr
zAR1Gvg/es203anvp2SqwSOQuEEdzV8UEX7vYN30OCYCdWMQFnZhqk5LJKoQUoEP
mkizKWRmJojB1U/PNC+tT/zvatcowKk74dwYpvG8fdKzCjidbiNVlkhIxkGCxsLN
SkKKHGGThAd6c0DEuBWR0Y7fSShW2Ch/8KmJFTPmWhkOQn5W1soID26tjkqPFHw6
V7jFYyd4JpnJpFoAllgWW7coSrqRIMO0SZErx0Pyr7c5B9lK+Nq1xsY0QUMT7hZi
u3Tdk7i8HZmZLaOC8XA0GOXeFi4FK1UoO0bJQlqik4SFuunKSkgFC1PW/3Jcg7Xt
VKTxLP8N4UMHCEwNRbtQH8RkYZ4I0/hx2Jz7+f69wUDhXuaDvp9GziRUKJkaNESD
EMgXBwTYbRGGmHrGGIVjLWY60Qf8seeByqBnEPx5/M1i3h6VEF3HtCsZX3Tl0913
FJeavHRdmRSumqc6ECyaInDfJDT66sru4z6qnYdII69yTwaiadoPTnKx6p6S5xSP
0Qc25L1eGzx6c2s0PJKt1PWYRu9/fDulvnQltIIfdCvlzzTs+pWtB5xUaDhNX0nJ
TVVaZGIzm4Ezg3PYoOA4O6GmXOj4RjMu8twL3N4Xa7fzwvqKbSL13y1fg50mJBmQ
Rr48BezF7pHXbkH2QGhu7EKnRoVoWV6M5X674zxMfANWNPx/7sSSqvwgd/dxNLDc
OS7YRDn1c2cnmAVN/vyK1WwWBO+PE36k0+JM5sEhGIdlTbrmNul0yFQ7hXP81UlR
g3OLem2sbt3GSN9PkSGB/TCCA7CR7yBZ1fRreebPwsrkWPhGDdP9LgxVL/sU/xwp
xyKhSMoYP5e3VJaUVe3lYZnX1HmICLlC+TQjsukgi+c4233JZvqhKwCb42GBofcT
zgZc9xdCKjc6V+7qkQd0Y8yKhaLh+rlE6tLcTYjbwYo4QptLN0ygJlCm7Tgh7NhP
YKwbA9DzfAcf+FxGd/1x02ydCjm7SBeIeLU43AfRZ9Fe/XbnvCqRn2e5PgzUyeBp
QRzlWeh7+dk4FR2RgbdlVxJmworRQFQCpDlZzubFpW7i0dsKAHAtspMvSCszopfQ
qBBkLHLROw5vGIv4cy+jFKvJfOxywpNkZ1P4vESRXuAFNGfT7Lb5E9a5RPTQSdcG
JwEexmpkIhsI32R2osWX8wauAlU21ACnOvxXpfYJvL4/UkLyCGJ1WcsJAMJEY5u3
Bidw7TyDXrFxg1n+AuOLEmBoA6uG/KFTnjJRP2txs4kHC9Epy+kxWGSOCOzJbv/l
eQuIX3oYTR6DMMuoKR/yVsNMLw6fxerTQWEOL2B+5FCPw6vxIOi/n24od1MHiCVM
eDRTOuWYkG73YGv1sW9d3WlZ8eK42FrJmzsCNyvhJL0RkujG3aMld5/kpinMRLWc
fyBW/sWUQPulA2uTMwJIQzACr82SJ3Tv1fNOhiUC5QopEvT7l34M/Zst2uSxVwEt
yl8u3MI+o4rar9jCvVR5kPE2T1Uzy6xfB+wDIE3dTL2rvNCZtt+nnHyA6xiJYzkI
mvBcgwaFWqhl9Hmq2ziNwqMbNUWZTK6dsFHvigdq0ngbum7tyf0g2icuTQCiaeaC
18SpKHc8FzINTMRV8JWyXAZQj8vfj+ExMik09rwIjrBXhKcvkPckOwBwi6xZ1KM8
gB5DXBVrDdK/j1ENsi4RJlgR39Xs5uZRGWrM1ukPr2iAiPKRB0lox/rzzXteWxSc
hGtvaSuUvEHwE2ImK6F8dvBfkLaNRd3+ft8USL9e+sfAqeKYhTOKLx6NuyanL2mB
Na2ypbfNauZkjsL/rFiOZ3ifYJO+oGWOQ9gPW5TCnFUCb8wVDbnecdG8NjSiKder
31tyo3JSGw8T7Vd2vPIUezqNVDaaSr0yl3/nd0Ga1TXsUq04b7VTEVtdDNy2Q7hM
iGgdU9KyMMDuUBkXTjJcMMilsLbULQp78vMP584miOsZlIIbeGlyE5CFoe9reWfi
6VV49iH5nv6f3Vx9YAViSkrHIc9+Jc9WqYCqKQDhVfcVDDwv2ND5THlkIxQHvdfv
A/D+zH2Ld29/hFPUpFCKJ13CUnipklek2nh/bzg/AxcUZXxmLQng5ONVFTOYAcvJ
P73A0If7oTjXotSLcMzBLqHh0NtE7yJAgFoF/CsRD8iQo1W4YxIg1MoUy7a2KBlf
PkgKkhDVqTbrHdAX6U2VOG4JhMYMAfQtA3YoG8enTz6JxdaJjET4VlbZT76mt9GW
7dVkZ2XJRrHkQmStZdfSeXrPHbBzOKF78AenuIyxBLNIOAIK8b9/HMbnLmv0KKPG
OwQbXb9l6KVzcKDrz+7NweYsj/Bc4MiMwV+PK5WGjHxdDSAdmdDkMV48m56ZpZzZ
7/SuyRN6twWPTyW0tzWXAW1W43tjsYuM3Ti8PamvrjDpOHi6D+zRVCiCa4zh3U+2
pFXSdoS8fBRI4ZuwNrS6/r2BvQ8zmQeIFC+s+Yus06dEXwTeYij7fIXOHFVnRATQ
obYvWs9fspVVnSqnlk4eIiIcLkE8tyMeh0TkGbQwx1KeOuzh+MrCF6DIEMKqAKaE
HTJq8t9GrzA0lTcmclXbCk+33UnWxkKIVnmS2LM/A5WJ4xgOFz2iy3yObOGSoDCH
YiZWzv3m9LFWaAcbohfW8lcStOU2sOsrZi+TkwAb57BZNIW1CyyOcc8S+RVH1z84
GfOqdiRe6Y6C7W9+zhZGce6ciRJHJIwlJ02Z3GV3qWpsOc5/6636pkrW4EaJm+yj
1+rNHcncUvVPwDKJh6GairkrZHuKWBNlEtR1VNpXyRgIPT1LVTk66lBtANdHVhoP
28I83HZ5CpdOxO/6eMcfhJ05g7x8a1E5XZIddlvjssSHCPrwF+6V7FA0O134MJq/
KBOih2gTxkXl1GoOayy9C6F2sEdUtw8RlCIj+vJ5g4Hw/ck0zgckeRMp7x0E6u1b
CzzKvt1awRNsNHoiXQJ6khW6en5WUk/OtpKHRzFV0uyZTuSHn0h5gKuEQEPOEj2k
dEXkpyWpkrwWyVHSy8JayK7X99EGMYUIw0pTBnfO7GXLKUvTOYU5neKlnlyqcumw
S3bM9UnNokXOdtgvFEypo7Uw7tMOhETqv/Q3W4eJiXA8KN9TA9mbcXFovpP9mdad
KOZoV0QM+jXTW27EtArelf5NLrIG0cvaOb20QPBY0U5Ise6+9Mk9WQWUAm7ABBdn
9lsXxOv+PVLTowHJ6hXjhYbH3+huq5YtNYi4wxxSI0q59WoFh1dHxzbJZy0p/7rE
zxQ8kDRCA051KLSPrVW2nILeWDHZaS7o8ERgA9TdPHgKqESAUG/saiHyfQknWmvm
+JU19a2JY64h8/R6HpPX/xvmUq4gS7Om5aEW0di35fN3Dw4Sy+VvqrRETt2LdwZd
yvvBbwvJtnnuncMIaj7hdzASJ0yYA9URK0JfRp4z1fzmTVSG4jzoqBz5ExCjL3iM
8BzK4R5+BjfyYa8WxMtRrar11keOkzUgk8BtUUNNI0noPYWMRTliid1XJytiTxyc
zVV5QwNQVlNeRcqIK4Rb+ltHOqXTyleQfdnd+3KMBkiY9oM/EE9mM86oFS7Trant
4eqoCk//UBWs1Dp6e0d2Z+SpAZ8KXPLZYw/8sdpmIS8q2nLyJ3c8+LP4itch3Lt1
CKxgLtxegQq/8sD0vxTioHlB/7KV1G2qub8n+2b/EF8qUstgFPLzvPHpHbZ3f7kA
MDNStl3dUs52VfdNbrRgMwhuMLnVZwK9RZ3GeyqNtxgrdMvr6o8JXHkPFnHFUckt
S0Xfv1FWfnu7kvqO9DGv6Pt3yyIRsiBLlRJJ6VhJIUSMVwCZ1a0WwP6XYafu5oXi
f8+oVjAFdjMD85tprm64f6eLp+vUFZ/J2MAOFB46/ZLY6Nb1u3HfOJq4MnZZlMMk
/vq4Q4uusvv+GgTA+bKJgXLko8WmOTpFGgdDfHr6pYeT/N/ZQpj8oIIBUfWbSr1f
NLvAK44HCNCgaBdVL04Bx7OZlE/XKSAvNgWr0Frh6zqBtpkNdjTko15BQ3kq5DPD
OK2oobwgEPM+mFdoeuAISvtYLSdK6uwZko4JqLA6O+jvcRKFjR2S5pbjt6ELCKOf
zwPAx+cPmOvQMI63n2YCQut/r95z/NXO0yAxXdoPFJf00y7Bg7wAK00BdrntB+tL
iqCtdgAORewj9tE8xxO2ms/nNBw1y3VIJeMu+k/CL/KD/FWje9C4BahECaksJ/Zk
y6rdHkg5wh3h0fjby2HzdiORmVFiAaZNOnSoB1Y8X/Y=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jhZ4hxnJbTfaHhhIBapu0y9WZ9K5PMiJ2EVOoiSnOgpEB5EbSATRXx2gymSUjG3j
h/74Ms6Q4/1oGqqy2Uuuxqj8OGqs8AaFzZgDnzg9ARydBCv2o60i/jpZe78voZhI
eUm4cSAzWUL7DRuyFsWkYAMYEy6EyFGjSBsbcUyS5RyRnGhBeqmkn9zEIFio41YE
ui/XD4Z0jXDQhfhOnQ6vhOVXol2kfxEbT68+y0sRnuQeB7gXe4MLPjckpGxqje0o
pHxqNd/RSBbwptjWsesoCq9DK/1NNRBF/pwhGZJe9uz0fVSOG/2ciGeezI/YIf0b
tWqq/mnCZ+WqJhOjs5kqow==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2704 )
`pragma protect data_block
8li3eFe5sXU5Yc1yriFwDL4YOno6hy0iv1TEPh/URS09m+QF0+oDa3jVzKcg5fei
HgXySjT1+sOtLnVlcTPF+pFbhUaZxaj+4voZqmyPdJIEN+tGpRyHXwfkVlWb9ABM
lFi26Lgmm/Vqkk9Kdo2wIUTV2CnytCeZNjx8exTb6h+2qLw6wcBLE3inr1v2ijq/
rT5jISTWwG0y+wRHpExdAQjM+jSm7CryXdwS/AlC2F1EOvI0JpUmqdPmqul6bBg+
G+b6sJGfGny6f/r94iZc5dQpktzVQiPhsx49TqADekWyhs/B7JMqgfwkQmy5/Qaj
JO0s7LeBqHHsqc0R0GgZW/0UqDKBbUb3CFTyQ91Uh9KyVl+tIiiPXN4a0B6C4nFO
b5GwFovATVwEc9q/FB+/b9G5YYcqoi1ZqZR6C0rE3YP3NuTcGFLXRWtC87oCHcpC
/iNpsCCBU0jlaKdb47OYN/6rKM6yTirF3/QK6g8YtUtVI+idmsJvUsq9DWtWYx3e
wMAYA31mdKrfIGeb0hukrj7+x8mb5O9bhmSFRB5kLAdQd1dZnGOw/5jQeEb8no1P
nBoYCDWpXQkQLs41Q6sxscsiAHbMZN8RUG7aFIcrlPKIVi4O4K5EHS2sN7Y0460P
EYk95pkNfGwc0BFoI+fpzaZAPxGzImuHrkdnqKsqeEVnj2/2TtTmG9CEARYsw5Xn
N9spih8Hp0LWdyH0vzo3uZk4gL28UEdzZvcUrLE/Jd/NCitMSSkRCTcyghjz2ho2
3yh/MmL6rDURNLsE0YC17FWW7BGvWH9qwak0EI2Nn66Q8gkoUW98oCx67rHKRPs6
6vFrmCyRwoTYpycIUfp1pb4js0k0X3ULeNGOIgBujqefSJ8/cXnMAP2++xHLLl8n
Y8Ykd/rCQVaDL3hiWXmrNzRy/UuOH+th7EmYgUCGuhcj2z6K0aN2gL2Vois1r6U2
17xKgQ14K7lioIPyXEv3ADTOyxw1yM08wCBUWPtT9gPywQ4zbp/63USwELKATExt
VxlDvaDQn1wT6k5wk3ZLa+pjQpBxEkESWGAXVN2+yPN3KrQLeiAW9J1vS0R9ve9M
Jjm+UwksP/NDLw0dGy8aTewkgIBNegthmthM3Mu8HikkUCoo4ODa+M70+GDcndtU
QSMvaj/sCw6/+YXYtAOJj5LQftZmT8B+SzWpaLw5Uqd99GGR2moCWxOoM5pxpsCS
tMYfbFPbR+Id8AsT9AvSFfuMrzqzrqUE05ptq1seKaIO57u2h/vxgOUVPGb53Llh
EQvSr3JF25fUupvIC5evfICRO2rBgGkpoeyQI3J03wCFHsFIOl0vv5OhxQVVAQHY
/D6xwz4LAqoc0AGEqtjhfzbKo2vnElLc0VFVmFhyxYv9ohotDRzy5htC6iz8KqQV
2U/A/eVAFXDaVvl/BicbbFY6pB8zvPN+lEQTY3iRyRqSuDtsfCg0gc3kE6wk4BGM
QwOHC6eMrGU2QX8QYrckowfHwtie4TVU/7N0cn7X6/l9k0PhpiJogFANzBafC3R4
3B+5Ma6uP3xKdxi0d3YCvQKli+KvbCzlN8zYjVFH6DKBMH65/UV3xpmdLXcLgL8m
nmqiih7NRQ/TfKT/0KqJOvI3fFofAzsrbbOcButwutCx+JjUfUx+sFRkS4oTHo5q
Ow6qxX38dlkGIo8+/ToIF5yjKNbDatD8oj0Lp53M2sJucwWS+NfntOdUt14GbP49
slpkIJDBnXmNCaOzwhiqX6L+QYwx/VuKpQ/wYsG5w3P7BTh9eo+7Z5Tq7p2vFqis
vYydlpdKS/ZIheYAhUwMT43RKEt5cxGGy7FD2sFE7O0MBtrA9HK+ch7zTQ3kzcpO
5XqgT0FcaRmFEGWXpmQjB3Osyp/a1yGKsQkndI8susKC5FMemRV+bg0Fop1ZLqnh
1Fmd2BPIdYoqYYFFizsw+lY7hnuKlTjVZK0VA/9R0uuDeK5X1XebW2mlSI0B5sN0
VyozS1tOGJpV7U/lWie+uK5i3APy0Z6K0uyHD3ODWoH6Jmc7OkxnZq3DAML+HVgJ
YKdvO+C+seu/2MH5wvhaKB2vGmKVJwiBKMr2ZZkr5qsacyU23Y7yoYiRnfWcYlsi
K2X0jdgk5iYy3Rhky8rYScBmbBWqh/eDZ/X26OJzyKq1J4bG3qgnxnZZxRY42qln
o+A5HGsF3cY9Ps9Z5el6tNQEk48nJTCEHnx7tinF1UqXYuCYNVR02MlDbtuM3N/H
yXhW7tIQxNxPIoCasTvRkPmiZ1ba3m0F9PehIGrFKFUdP4eGpHS6K2KwF20QNqA1
miC4fJvM175ynIj0SxyL5E6OePaApzbuXm/x3hlj5biVe4y4ZwXQCEmaAHuy+ZSM
nbyh0QhC/Ig/w18pW08V0t6wk5+5rcGN2M1C4D750uZs4Uv/yYE1qveH5Z2pWOCf
8jl0176YqicjwW3Smt2bcC3kkxNaxFis1rQwOENiPIJD1B2R5D4NGdESHAK7RMK+
dahIub7qm9TKI6nkIz+ZR0HRqLICNKxWvA7Nlxg5rRdkKmbX8LnQCG2IwPFl9/x6
+kyG/IhwI/t7or1dVXT0mpdRtx7In/YlHJPT5dc6Q1zkAi0KuNn/vJXGM8f4gzNu
TzJoWzCFtXzHfGi3sCwgfRLMKOJ7fwSlfbekauYC9siOsjXPgcqhAUk/TS19pIOp
QcD0iQ6oGzjcgvescgXZM472lJYJgyFJ2HA8WRdGVKjPkgUl6P6uqkjhKWeQz2TF
JMbYCUsjcOsUtYkBTCZOmGXPjNiMRsNm5N1QX597KzJ1VNS3jYVni1YWfF8NbeWl
NovEAAmB5pon/6lZbjbXTxE+BinOSuIqYB7I8ze0UnGbnt97sDbjLYS+WmuD5q6x
LwKgYrxjwh3MxAg2ZAACHnSO8XfblgWB8TkxJKTQXcyAofyubFUo7U97APln6gBo
H08KRANvKeBs7m2pWIEPC/MUgRvu/i+Q5rpSuGaYtrMEZZO5SWiPFt8GwKEiH0V0
QE296gnrJs82PKfNEGIwGwQclKNHRO6Sv1o2Oe5fXmN/fnzSwf7AlLX5e6fdVXxt
kQmGGDB5uj/cG3tsJjgZYo/3SujbSYurslZ2KvPxjUFu4ZgezIdKDjrvHuoAvxym
x2Xh4nQOW+FwIew4twhL1mwqO6fTIYMlcUQqGqjX7z/sOld+t+VbQXH6t21/1xod
m8IcTF+5v+F+wzLcfzoRsG0rgKh2X1LKLEL1vPl6c01Oh19ehtTPccPNiPbOXOiL
GJH1SN0dupkjdZeRpP9yVCE9ETC6wlVBcAU0vyN4WDAwD+S142XNrKwnbE3k4LqD
gmGeK/8O0J6wcGipKg2zO+rZC2SY2Kq8WCdCRuaY7wdlpnN4PxLo9FT95xyXG5V3
hUeZQ3UBY49hxCfZjbwXaZxEeHDrE8LEO6vItGamfaWNGmOqIwk27kxSPKxHSaUB
QYdeDUn+KdvrEdA8OIJDeTPKY7jYWkI+ZCbnvBw/db5XJiXrFPx7sekX5Yu9+2fI
7AHS4Gam2uVvOOcZbWo938Z2mW9HOuCtjhKbjmUxmPvgFetx8AtwLaKi3AobksoA
nm0/+wHnLkmqJbptqdhC0A==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Zaq161sF9X7kxNLJO3Umjcw/rItuYG2qbNRM1j/QW7u2ht9gXUAspAEdGDQvJ7W/
EfNJaZJE411wQafdeETf+aLVNjMxXr7WouO+MKLph02Q3l/O5uc22cjPTmCIy2bh
ClE9x2NkWY/YgCQGyae+CwU177A8nr2cSvFkycQfgdx4cvsRDOl3JbamerQtNevL
e4FzftD5pDMlII5u6ZKvqwhaxVmABuctGwOBBdjXjs0jOkNfPKNufT/fClrm/fI+
IrFOjZTF9QmNwWqAnkyJlPVK8ti+8UTPMxZc7VK40JvMGN4S/gwo4v8vhG6ojP+X
McThVC1a4TZ+ZX8hJggghA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8048 )
`pragma protect data_block
/eZ+1BGrYp2jZPYl7I77T07PmmZKmVqEQKnMyV8NGyNer6x2XqToG+NOjy05ZAYZ
/lhrWFLHXpGaKXGJIz7nz6kCB9APjhlXR31tPDBqnr2T9zkNhGT9Zsl1JpuU5z9r
80qAfWjIpuzMQyqIt0nZIkNq2QaAebqI0DpPOYuTii7tGOUrlQdaNCfFidysx9KV
nUJP36bL77QIQKmkDs9pFj5MCaQ8k/NnG60wWVyliGBm20ZACQj7+F1vVXS8ntvd
qLuS3oC/ofJvbWB4aLNl7hF2iOCzcDu6TvVGBgC6ROTtYh732DUKw8+rO/uHQBXD
NUzMlem0CT7U5HQUiOoT3800g7zvixNn687HPpCLNOKALb0KnuSc07ElcKuMZaVe
nXre0cHXBPSk6mnj+POqcz2Ve7vzILc3hfxr0XpEShVbyHu2E4yE3c3yxXI8HCzA
ZqJVh0f09rKlcX4wuq3d1epDRyWZ0HyktiUACsvfoNZlZ5/htZRlivV0Zr48WiAf
AQLzeXpbNfYxiqVBQWVNTt5NjbRddQU4Jt9y1+Xd9G0SVczWMGTKcVg4NFOX1ldj
RumN9PlAI0y/SWz4HmRBpF9vf7oB1gYgN4WwlM0tQPsexdn+J97twelC13qyPEjN
hmta8hV+wXJps0lwBL3sDgYqCvWblD1Zhoizvii3GKVJZeSj//g6lBm00Q9WgIe8
zmAGN/L98NLmWpBwj390Jvt5k1AngJDe5ZoUVsekPUeX/iPNdLZZxgub8tb1gXz3
VAbI2b0w2J4MLTShZ1AslRIJuThZwTBOCnnTUu6GtSx4eYvrDRHYbUsws0hmyYvG
5iqO/aUhS2ccLR2BbWnxwgvjgjVYUZKNePu77WOPYA4MtBvqbgSC3Ur74nzHoR+h
iHHfXmsRt7dSCOquC9nsZUbldU83SnSfANm0QWDDAopdb0bAvEcbcpnbg81myRra
XEiOPO8zAeJeFpZHVqHHrxzE/M2ADWpONdWGdBO6Q9q1tktwedq1cNbuFFYaIdcp
66JpFQbBCrt29bW4UaJQL1AANtiYE5/89NcTaJZ/LskBlJEYoCYVaGA3BOtAVzrS
SRy51oCoGyIwbGhJsg/893qlPdbKsXL7u4xADPX1SP2+foQoTcZGfwWhU9valsum
aAhRUVShrG7zwAye3yddivyWEOumztqp/9eRUIRuWiSd9Oa4ALyg6EmwwU08CGQO
0RDJlNQAuFKgEKeRAFGxRZpHpqqAVV1pXs/0W/LZiyvqZvsBv2Ll0u7LdQ8w4P2v
iwcLq/bR1uA7xF9oCSpmls/pYkridHGWMHznxXGz6CebdreQWayHtrkNOPPaR7or
Re37HoiZ1jTzPjJ4s766Min0ol7f0XN57MxTgCuax2+IcE9iWO1+N8T4WagisXae
86xaLVvD3o/HHFgYVQHAUP/kRT3Qoag6pffrWwvxWothLJEE7+eKu8R8/aI65OcQ
w2t/ZqfXGYKhHyMbKZMLwoRXim1gsp/LT0D+b0WkSqS028QdSoW07KT0htjVdt7y
uOImHq+st6ZwlVQtHMG9UIHSrKjVcXhmgHpUGpND1jO9zQ8EaLXYzF0n/xrgFCz3
OD73vy15vPp8WB8HIf2CYLJ9hbexDAMqGIapd9nITukDxWHtMKBSPUAhK/etnAlx
uTHiBsAQWXYUz/glShoO271mdMupwUqtboBagxOLHbh3G6EFrFKT78G4y5BahNiW
eYCmyFFnszlSfkuunhLIJzYxOpRj85cvg6fu/j06e7o+0cD1Sa6TM38SCoL65YG2
QZW+amTjYv9PwzPW+cw4vI3k42QOQtRMnpQs+k9wTMWPkvLdXg4MDRTvBz+v+3h7
OcpLW6kvSmpAujEI7iD/c20/5ubwaK3nFux3HjP9+PijwtHyXnnYOqgRi6BpKCFe
yfn0jvY5Mg5oVg5L30z9wGWcokkApLQspP1RQRKAVG72GeiivEZfPWvtXZoHl0mB
OtnU9XSXuYJx+rrD0sNdRGkenOmrozqdlGLUF1VKKVK8b6IA1v4p4QYAkhob/eXR
3VFPae/ZKSELX+PwbOOlhC8hriCsP1c1Kll+SXdLFG18dey+JK1seH/BBnNhOA3u
mWdoeqIEtSwoVR0HPG3gguxBSMObIOst2QR3eedkhgH6e9FfRpjB7cjPa4Rq6HFg
i0aALXVQrgzOd/R4Ta8EC8Y/ZtTHYnZHflVYTx2p2MP3FYe0B87PY4K5wdiT3KyM
LJ2yGENKhmuG4R6gImS/BA0DZFy2XV9S71lRK5aS9Ag4MBeNOJqgCMLuLXARMAqn
BWJcLQgkxUqPe3gfzDI5seSWJB0xkn8Ux01uFE+o9ZI0IBAb6T3WjMwZhXvocM0f
hts+aNBjybQc1edROzMlyFc584RRemIcxmw8/73uIWb43mTjxRWPaDLKKVk+kDWa
uWf3+mwT00CrGQOHetbt3VoHhYXATyA+HpgPlbrIz453pWhyUV+uFenkrkytRi4o
/8em31MXEtDAf2WVN0RduVOLlQACUys/BOZyg92I+yy/xVpMHzSq+RVeviCUuSPn
nVaKO5zHDXGJGr5wcZLhcsRCiVBYgO9pzZPiR1NLEuZNktqS/Bg1P9ROarSNXBZE
KzXOAakZypDg9yJ1+PY29xfQqYFs0RGIWmcbFqODWgEhww/U3S4dgri/a0FoKNI4
RAo6kL3fk1Wn6JPZ6bu8J+u2nmkasyCYtzvxim5AcIO/ACtAMCklPFH/zESYegob
Nq2EPeISyVL3nDf3jnstSLC2Jytf5mCp3lwBkrNkcsPrx76XyTZc418nWoImV59S
jwKMUWTc/dYSPtHgyqm7jK24RNaO5Sf3XtOr/JI1i20zylEdOJeNCtR7veOCEocH
rRomXmFLozac/8/peuHncuzztukOaiaOFG71E4Z2nsp7R4dCCV1zWkO7Tnh0vVeW
wENQLPUNNY0R1N2UwL92rZknNyE4UVRatz/4lSmZYqfVsTWGRAdXNXTpfjHvXjyE
SWOcdscs16+j2RQUCPPi3bwOa2mjb+4gezIldmpnRv/FdyidRVvu37wCzeX266yE
5JAJXt+DCDC0Rmxlm4/ZBx4p0w9Y03dAZ+ipMLm43ho9aQGCIHGy4trmqkRtjTvG
QZZ066rugqvKeiPoS5ThZatEhZya2pPAMuRnMaRHY4aGzGuhGFg3tkeLnTu2AOoz
2V/aYbxrhuZdqOrDNruPY+3fcMZRUKx/e5A+WtV38tdPJBGWU4kwcCyzCoUwMhz/
USJuoVrKBOL7UQm2CkBVFzbw8OuM3dU0YKnPcMg5PgKzIcmdbmMn0B6EFXjicjhn
MjqYi2OeTawLNuqHAF9zSEDTxblG89OXV8NlCdRK+BWJ2RU5AyvUIzH0T06rklvz
OjIJPqM22L5M62LXamEykAuAkOFBpawH5lG/GSrU+tSxaG4/wyh2IijOkzKWfwG9
lXyCnbMjoIPB2gl8G0diaWCj2X1q6c1CKz4ZTTGrcU6Wl0nUSQFcrtzTaH2GDI8X
UYoUYNMPXDy8IAe7iSaqtdlg5Y/16lsEGLfgVUJYiY/S68W5nMwnWKnCqbiUb6fN
xnsOSno6HvpPMpfdrgEgJaL1CmOIsG2VIvKfSj6mBJe7UblijtB6ip3Z6+cSMI+N
QbRKyqzC6E8kW667udIhNJ61EPw+rq5EJYAfYB179m0udv7BFKpnAj8XoRu3qkew
0p/sxITpzFFEicb8Jq9wwDRIyuVXoUlDJlQ+D++rOV7k7Ja5R87Fx2iwz0CjTR2n
GdpBeYYHqDHvhicmCFS0gQmNK9tQePP5Oie4f5TqiLa4i/n5vAA45yK1r+pbaRIg
jVap+2MhT4YDS4pvFU6Khx7xDrd/wEGeUm1ShvApIIpSvPOYKFWKwLCStJXmQWcK
v6vAgWm51oFIKLt0rM014fFwHLJZR8pFyusgdJmlvr03DaMafapCW7hqmaZrjUEV
JrorIHecoX5roPhroBAfI+ZwT2OombRAuxavrTpaYmsN0HStTpjhjhj/JZlIm8KC
KIPxnbQ8ADuv82M41DyCsIq4urfWVgCH5BMuFrs1BOuHEpjr/1ZVpveaGG8c5afz
2LjPHUev3xbY3LTR8i9SiuyZIl5iiW+1AOSRFowmQvkGyj8zbywlc0ZYaE+U+sJd
AHCwTVeOdw8zqKftWabIAPCfLZRIxESHvVdl3ZGKh3BRAwl2dAux1oeUi8j3ASCh
n4LvwUOS3Jcqg0z+dICxqVdZ8wDFyBKAMRUPpIZQUjJ7djMjtRDbKph9xpA+2A9G
axlD8ZELOHrFT1i2pO9oLN7UxhCV9lMpGrSRCh5+tej89rEHVWfJ+PuIUSv1UasK
kC149vFDT6rQca9OJOofvjeoJNmLsoR/Knf4dLSeDLl7ISdP18CItna77kwmcUxQ
rFBfiU9wXBe/s382UgiT3TvHqkVfti9lz16cN2FhE004NfVmvXHw5LGLo42rIPZb
QSTw84dQluxdBhYOL2vrhol2rPmjdE6eFaqvVvBATyZzbHQ9GC2sAtPihuVN6tOk
g81S5+tGfAR7o7rck/Ae+M7YMC9A3dLeF3CDwGokh7x0flnSER1RrDddAjIOaCnC
70K2RUOGQzDQ6Fwp9e1bZ5Ayn4ywomVBdYSC6UjdSArBryD6TfCeh0JVS5meHhNo
ntXaTK++uw+u6qzj62CTH1vbX04Ks+AC3Wp/sAgxAq1U0550EMKV+KPlaTry+7Vf
q+y2ZxsZZJ7qH9qZSHoEIS4BKgANZuzQ3+pB4mFRds+Ng1fgEG8imHyljPuOZO0E
BrADdnKETuii49Rs1bCacRyJL+sVdXygLU4/zcxWZR0KzPcIrIf6EMB433NFvPE5
tBw3WFNcejdPkDEDvdwJzuTcrX8IT3B5YjlqnJoKXcZz3TfeueOQkq3gXnMMMtz9
jZ9aXVpdYHW4JtVTDkSEtX5hHc7XMC/WDnDyVh/Kf2XqHsq80d2NKFTJZVetFKyB
ArgwkpbmC9Hs1X2lCn3yrXvLt3yxTZsb79vxTuKlOv/VQxVLxuI32nm9+VeIFcsm
7TLlscvAM6Y9MH0n+p8OC50tjJNXfRSg2bXDC64wTevP2ZDf2hYi5iDVFRPUugsP
gCRhflFFlcf7kThoVO1EG+o4C3jLRIM3T2oMjWyi4X6FjiAR265vhv4gJJZh118u
7hSBhKlf1obZOzPSO1Ol340uvwudujuXZHHEw7unEerryueU0hAPqQN+BckI5oaR
8DQz3D18jXZkquRtN6NC9kpcUBaVpKiNKJihZSWrTQPz0JiDPTBQ/HRqK6nUZ8nB
f6HkAZLvQY2flY93CQwIu97zjT71S83V9kf0iwYv9WP6NhWANtwPOfvfLgtlt8pU
p6B5/K9l+xRYVyiX8pNuhZ/1qcEqP8nnpgpEKQxWlbrdsv6Z+4j9XlQYo9ORcOho
NTxBdz1xMyqpQLkug0C/nV06tomV+RcyGeu+H4o5SIBs2sjspr352ZqZGWXUL+Zv
77yfOohwTawZv6ZDMLz8LEr62Pj1RuUkx335pMrq5v1emfAM7Rzo/jG2tVRez+Xk
+SVkj60TxFGV7yXnTo1IXvCWaSiTnCD8W7JD7USbzxFzkqTKNap5KRSPn+xyQR8D
9imY5UWLI/1D2Z7ZwS+s4iO+0QFyowdabuk9dFXdaUVbuvysS0fvO5F9NbMVY17s
ra+A8SiXDlcm41L9AcPXr/u8P/QHDTxeus7O0+N2f8Yp5uua0MN7pOjydT/eRk1U
1IV7chdjRiGIyL4TcndPjJCbmdW4AXeJhcAKJ85wzUpn2eJQB5leRjSBzZooYMVl
gkY0AAC3j0SZIM+DkjtNf/6Qa0ULsEYz/PMXSdRPX/TbCrkQNMk9pH4MZ5O3S9jp
RnlYATqHNOWwqI9yaCA28EL/qfx1bM634AgCYdzSIGn83WuJUJPXXWxX5ghekBE3
i7IdpTPTp+kCP6a5fCy4o6imDgAGTS2T5kRSL7i0oTTyrlY2YyQ+zWAnURGIAHn3
NMNyKesSO8NPPqDpqE2q2JJVyA5123mE77z2cIy8THhIaJY/aC0I7YKF453rPDX2
xzSiK/IqUf3u2IwIBYYy+kUPVhMMBacIWBVZNb4GzK2uy3VBXWu9qJ+S4oL6Xq7s
uauOBkQ55V44OgA2NcD/Ui65pcR7Rf2h7pSG+IAo3KLTh3mc9b2x7gqWWojXZDZe
lr7U/H+nRtPJ+0k4+ZCHvhv2QOhppvksJSjGeN7O+LsfU9TcqBjHyA/M0NzPbfCh
AEYeK4xjY78s35D0ypJYmUZtW3Z9EHGmLlWUB612X3J887UXJaqn+YdDs25yYqED
/xJp/EhbsufHVUNRvK7fTtbW0drgfp/y0Wa9gfJeLGONHLiFvzOBwGZoNF3HjYRH
jndBsq6lWyRtHambI/bQFg7zf1TduZv7vMEqBcl4FNl0dqOyPyc/pJ8U7ZG5zGJN
uUqpok3QaDGynjtTp9lYDsfPZeyvcrMIf06rd0oStqH73gbHlghfNFs19TLX2H0q
X1ux8uhgpDVYyJhLJ3vE8bhlbVl23KEGV+1Er6svo+lOICrGuEmlSVNelXHH87Zj
bKuRcxxgXWIoVL5xR+8w+qXAArVOCvueKcj2eLnHaDuABXitqiohvJO5Na8E5TrE
gLwbforUgwt3WgX65y3bT5vPKxUYRgM4jacJbuyGTuBFt/L6DOZa5IB1Ae3BynDL
Uwl+3u61j3WMMCxQDYIMb9u3tfZQbKDJW/4ColzgkTHYB9zqrcCyzpgHYb0CbwsY
8RGMssSFffKQ+mSePfxyN+mxALgvt0U7m0k1PZWefg8GMCEoaxqy6VHQ2VkfB07u
HrOLn2RgJZW92zCUxX0EkiG9XgWDo9Ed5XsLWPLOL0Vqtuhja6eQcTeIyvlmviMP
3uiFMqgJF/dQubiZJWgKidkzeyjnsDD3KJDJxg7Uqy07X4NY0XdBcIGUY6TDyAEi
AdAXuQnZPdxPkcNGMEEMFe/QBPVpzkXgvOrxoZiXFDNGUb3a/37GYfWcSs6XHVK8
MaUbaOvlQ+w7ZbtWKg5gJcAbTwQO3T+UKIlGkc3J0AA/qEBqIB4zz19Qv8qe8/CI
XcAWL95c/P6+9VhbGuUDLTIgQvgos5OLj/RqLZqiBTOOqwvbs9FP/NFN7Xfc3bna
xa9TFFW7cF5vPXimJ8sM9RKcquWYLApsnHMaCGst3B58L+nSif0/Jp3y5MyRCkV0
nPfjccikswyyVFVObMma0UYfhSz5Ui8oWElcvbgXJXWp7o6lSgi5mei2X3DaAHvN
dSB/jmdlbQG7xpdwNXC5biCYo5Akx94R51MwkgY/coOnIibeHzvCQNsC6KTq1QIo
mjxB/Wqb0kbkPpQ6UMjAkr1S/R6Z9sFYhiyqXnRiHpx4E5nYc/4rTZUy8nc5Y8Kh
2pLC9e0awOAq1rlYo3gKjCq0xdTF/IpqPvPJjw6H+DBYhbsdrIp7rDRm+gGvsEJZ
/AV8/ZuC6+QK0xfkrTyrsrfZU4BlAT7c6RUBP8eWgHHV+rQyPLlTksNom2MMYH6z
XlvvUzdX3HzWsGutpPNjfYqIDv0MQqvL03Vdz7pcuKfiwz0qQs8gSsvCdpafdJZC
zr4FiqmQgB8MzHQU/N2rEhJ84Us4d+ebY9ozJqFCyCCkvGne9U5VYMPM9Cxsak0B
LeUNJ9yRBOMyi7v2UcSwTn3uY02GwLr3Ujel1UycMqYLF8pSoo4wuiUD86k0jb/K
/akyiA/H3EVTvvSBMEco18qOLd7ZQ3YO6lw/b5wGRD93bryfPzzqZj2BFAese4YT
iMk7qXy1AfhRb0ot4uJtg41syJNNsoAZ4JlHaonVJCtz7M/1Dgl+oWz9TeT05hkH
1SDsktsPzsZmingoiwYxdUCqp5wELGxVumQfNjT3Ih9Isoi2kd5V1FwVve5dN51u
lLnkm0Mkj8LD5ku2RwdjGZdOQI18Pcs6mdl3KrnpXvSDnfP4vX+ukXlsQ0diKbwh
5E3ixkAVKKB566YFHOVTLOthyoHkJAxjnz/cN6d86jI1aD4hQNPjVtWMofFN0pX4
dow9BWFRfuIsXMQbk3Y+qsqadudZk9yLnqwbg4MTkdmzEUnBPA9t2n/7nxF086zZ
SaZFWEQHy3eoJgWwKwCSlwN0vGF7hdYfZH1oojE04nLlgIrmJZ5WndIZbPizeq1G
My3owzEFxtkcq3MUfcIHiER9yDpZhQZ3GokKp7kHpNFBXR8Oo9FkLotbquTWJUNn
XGaAXQhZRBk/gm0fxw9xuSk3/+BJsOMfa2gJlF5SAaLIC9Hk01Pxk8Bb9aw49ipS
c9DwgC4+j8NQqnBVNizF/Gj4GLbXE6cSXBlUcN0kb5AlCrQcLfFXp49QLeFvn3bf
n5BnutZkmZyeXuBCr6FAUSdSiiV3el8+/vLTvF2rIuWDL4dkdzFGvRhljyknRumw
xG3DHOYdrVMztvWX8+Pk//onjQPidCi661lX2gaDQlKCHLznAIVlMRF5+jYJ9akz
5+FbDcdaxihQQAlDrywrbs9E+dJVI+SrtCC8LUtTtchilxRu1ojSEIJe2zi2kMw0
8IuhK2cVnHY/+WCRNTkL/ZLL1yGLrichwW7QWyl0FbzjLpmCGyo2WLUWkBjqZazn
wQ5dXHd2CCG0VkP0aZOSpCRQ5q2c99C4rP9z6FPNeKQwBPReaPy3Tmt+YmHBZXQZ
+5gyxqkiBvjL7eozjji/qlwdeLVejYdrIiDIq02lDb44FN4KvXm/1intcsUo2juz
y7swYsrk/UkfLM8vyvkT1grMAAkroFdRuEDQqvflcQ1/rSNNVgJSuwmQS9RYv+Qs
MQXMu2pNblRhZy9TwGVPOlSrHsj8AtHH7N9e8gTcB3XyoF0L9YPTLuO+RLw2INYR
mA0sBFNsrBzqCLlAsem5+KDepBk9Go99R9lZi8ndT3DCQYvg0EnpVVrsgPw01Ar2
5UbWkQHl8ITPBK0xaaNBX2j3+VpZ9ed+EvwfBzwiCm3VeL+U4b+pJKo1SZI8+zGF
3Gvtuf55fWhscWu7Lv22Hik7Er5qJiJaVdyTbiibZiZOxDffeQxKzY3OESSU16yR
3sHfTpVJr9xf7htWE/fa7AYuImMb8x0ueK+fU0iiWM/Zso/nc21hJjSmg8u5Jil6
EFnBuEttFAc+mr/eo6abQMu6iUafHtSRnb0ZcRWjt23/ghjkaFXArb4brXCRWxnF
ZiPCQ/qJxwjo8EreMs/cvEvH5F/KjZKsNdzqIFrdL2zmkrVMZJ26GZvPecaXCBeD
DaSUvy2uWskHhHu3Mzy1Ey6CA+cDcobM8pUJkS24hsKJKJa2JKqpRjVwrKKlZZ7a
4RGdMyUKGLAvq/sncJn5XsAGLGEyZegqKye4P8ZVpr6Y9OQFfZSR3nm7B/zqQQDJ
IGFt2Z1qibAzsk1y5Q64N4APgHCxZ+2sis84LGffbgA/BnLD53DzY31gp3WVFU2O
Abepl2yM3sDlg+L4BDWsM23GOH7pjp3uyp98jH/XHKUKuN1h4bZodlZPp9awfhKm
LZlCZugI24Yi8gAAfmTaoyP1TLd+49+hYlaKTw93fsnZ6RHLJnuLDcIdqJTwpuhc
U1BMyD2ayYH8uMZojctdTGACVPkNsxLCBKMSSXeLBZ8aXDOQviIkso+s/4wTTK1x
apoW9cMovOkSnvHCvAORK5HQbcZ+9YwwuQw4u1IbTxlWJXj+Odo3q6hv0hnV6WrN
zM0+qCZoS0AB3TM8tpPICzxplf9Ltdtrg72BiFOgNgnAQZzqZOWefISRsCwdUSBv
ir8o89k0ve9iT6SgQTTiZYf4jIiEt/jn8MN/9YBI9scW7a8jnKloDQpVyI+hUhRe
+AL9FCdHhkOUsPAE//HTK23pjgB5sB/stOlOV+Aaw5eY0d+PTJU8vG4vf7vYXV7Q
ShZrwysVIzye4JmEMBTS+YIOCQYVeXhYKQBbbKE2vHbQFgiULH2L5ZdKbeER1Z1D
huTPjS0RNUrX3hRgted8ZmfsLhPA4JFAZHlBtWlEmizsYw7WO/Nk14nOfP6eoNSN
R5dTMVvDZ8oVtmeccgh6a788/TM+zm1qE7aVTFYd18XlhbNDLv8wubUgNvT+z5rN
umiFc0wTNcxU939H+hlkiVnoi9qsK4PIDz0TeAQy7RO01+72J63fpe6qx/Uqv9hL
sfB+M2HlP7Ob6EJC/A4D/PYmhOsD7TIm7s9b3DpVYuO6mMrwsGlyc3gjnte3NL2j
sUhTKdm4Pgi6qYlNE72HshjHJA8inP2VFmRvvq0/I+eAvPuOGmr0T6GxaTK6pZbK
u0KzshzdAqz6JVz9jccjs0JoTwrTy5+/PdhonzgYsbVkVKhYG/ArzJrGY4nqbqy9
jUfctBgYIQz2RtRmvsuwIcSBetYqzdmUNETRsnxUZND7Rq+NCB/P7tkHwjUDs5+5
QpeX8EpLxQgBImDvQC7YHFNUJQiaBhzjwL522EHcYi+wWMR2LeXWP7QIrYZG+FEg
jFx2bQgBDKInLoatSlv29IwpveEiSWdxsRNaqbIWOjDG7s9K5/r7wR5ybe0CGw+F
yaSN9zanvDZWcBFwFWppdT2TMHiPQ4IoWrvpvifKZvGQe4+ELMaBFEGeH22hKuNu
T59DrT4lFMNlEtgdLm8VZD+/lUbZ2iG5G1en7CWg9+YJVhi3D9TDdzFup077SmD+
Qi04qOKBnA0bOaiZGWLHn/Z2+odCx3p/KhgTdFNTzZ0=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jryF8nVTBW1JmowivDktSsFt/d/YaY8M0izN2QtUAmGVGufwlPfWcFuHjg4V5IPZ
pmV6TFFVwO4rNCpgb++r8limNBhtkkcmLXnYwQn29tPM+uuHc6a563uqcfIMmqal
04SiwgzJtasuGRk4qPDtd4eb8qr1zM6IXG+viTuyddef9xf7K+w8jhJ73pLxBTs+
7vQXNsjaLDUTC8ZsJy8ILdiwl9mMrKBTNzk1QbChbBBwLis1xfuYJimP5OQDLiag
SZqo3eVDatpzXTqMkXpU3lrJ8804Rw0+fYWJEzA/E3mGMGI//0B87nbeQ1cDvY0l
7WdatW90oZiysembmJ5cHg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5360 )
`pragma protect data_block
SiML+DSDiu1FSGRrbPhCBlXb1MluWs6F+RzjM3l2CTTIGBPt/WYxY7CcQBoro30E
5sXkuVhAhP/MWjPM20fcPC89pTV844M85uznaURjzTDAUswmztNSOt5B9nJhKq8Q
vn2X5lbhpiIy6myzUId32vOoM+URBqucfFJEWdkkUgvL9aXEt6/nnxIthhwSnnDc
btJkZcvAJweD3QIMB3EkbzQWaiow51dPGmr1rdvfb4io9+E921nQnPd0wo2W0mZz
3Wd/6CsGbl9zS1Witq5yvbG09aVlXTb5iGJ3jYasquxyIKP8Ex+fS35yfv7b8FkQ
xR2hKwuLsD7d/urxTdJjMi8e06Hi2rUNAX0Ym/4zwizJnvmmonMC0XfHO78HX9FN
z8jXLde22I9Isq5AoDX2F/Zc6eOT6/CdWKPgBOfITGBsJRtl6MBRlgv3NPtmZ2Tf
q3pjjM7QI5HOob9uOnT5hdJUvwCOqcvwYiila2m4wo8KPiIZ1YD6OAYATvD7RfYe
ZtudxfqOWmqO0obEK5FpOl4AT/gif13lrRQug7uKuSVb85GBACPmIEtJKewNUNyN
gJJhmrcWuXfc2T8XKgs/FWBxw48kgHpf/XEAXSBIJKyA86Rj9Qcf5qvJQtwOJ5IG
HeoyYXmAZCROMDhW6DCqWPLFDgJVLiDYpoRdwZJYS3MYeZYlCxOEAj8b7rHWhZZN
1OfnsNuWGFAnj2qxcPBFxWsUvAvnIAJcNebjWogyPRVgmbUyCO2YFpJZyciqgT2H
RaPwbuRPslMqRik/xjYmaPl4TvBDbnKLGtCs7gwF8kGDF8d1w8XVPyKDmXohdupZ
tA5GXUU8Ta1Xrt+8G8hg+Xgav5hVbFRERLoe5MVz6ha0Z1t+uujsqyYE0hMWeiFg
Eg5xtf6hbmLbJ6A4/uay5iTwEbaikv5E+94To5NMRHrY+7A46EX0nkh2bkgDKMC9
C6+hHhmmGlmJ/rXLqUqWWm6HicJq2Gej79VHrmTQE4gIdg3/v/dHHQdzsENI0+15
sr8CsjApDvgvGQMG59WE6XwwvW4GcB3PKDpIq6cBCEgbM28e6PgZ3EOCv8YSUJGV
pOtRtAysUYckEvXJrfamuHw+VNMIiMLIRr/cjJgttL/CmgD52h5o8HwH56PEQPsA
L/Jmv0jvHWGQkR1n61kXx4OS3E65RZvVgj6e0s9WmuuZPJaY/kg8NZtYSDDCp1OH
uOxTnIZdebGVi7Y4Zy3sIxRNSCyquTGMpH9oesGv9VU7VYUtBsSAEMrHv3zHXqdr
jZMbRaEMRspmmY79LWDzCltfSf13ihXxh7Dc9fZghs5x4uH27sxva7tQh2AFAPdd
vutxmWS/qrn+rEhhaosyPzCh6Pey733BzEvk4a3B6RVKkfvXDSrstvIxScWGS9Zu
HS/T+F7MZ9k9JwNjpou9YtPs5hb2m4tQMe/xoRupmM/q9o5h7caWLj5xWY3ruR35
WkIFlpNqaPZ16brvoMleUqvGcmWZNFlYSl/1fedJQvz5YLH2XThf8+fbRKjCtAdm
m7ydtsouHPvFfEBk9svmCXpu1VSdbYSUAPwWxsjxzjs1TgPUP1xxDdHPXz5dOWjq
iijTbc7Dxsw7UNWW+EYGvnkkzwK9KU8OGhqZRnbaDwR5jS+IrIjguBuPqWs6fx0N
1ij4y0z1pDTM4tGa6RTvmuannMwns5VG2VVlPzAs2blgp6JtTl63w17NQB5/j+Iu
IhHIuiKm7LWU7RAdnGiLoYaq8rv/ZT37PIlqmokLpzLnye/BYbITHYOuEyiJHmPm
IP7ZgtAb/Lytu5W7Tp9e2biCuMo45NIvtQPOy7ea0e5u6ZcIYoydhT1OHDUjvc6g
aYkzMBd5VmTUZXE6l80SrR4QYXD4VeSCbQarJ4VTv0hO+s+u4DYDDmD5EW9dDpzI
koeq4EeTv636k2i/RkNsrYvdEh7bseW9qakZvWu2YvL7GATC4burghe2xdv8QITH
MlTTHN7vKDsg64C7iTB+jn+olaxWZQp8ZDR6wiNi2+vFhTMEKL34pZPnWZhw6crX
Cgr5ei7m12VKNt38M4nXL5CxSS/QxqM0kb8eHO/kejfdRXvCB5P0UQVXUvXXuTbw
9eOA2p4ieDTn7RoBQWlcjQ3z/TT308Ae0IMVoPFMwlVe80ZONGufsl94tbeyiza0
NGgPGuPC6bkosGEIXVC47HJFe2cSIajSgdoExYvNViLC9Twr1T/K2JWlzgT0YtsL
00aja7wQvstE2kDefAv4VRLA3hpPi0KKzd005mJ4AB/1//PcKC0YeVXSIsJpoxjl
5LwOnsu1vsHLrIa0Osea9XlrihVkKamYeAfMCIWaFWgosjMy4drrQr5C7F1o+U4J
V3Gf8DPThMsLABGCqXCyIqKucP4RavSZesjWMyHdxT+gOus6Pv6B8xQLrcPMKhX/
hd0MVxUJ85ep36cYCTMQS/eVDK0QmK4N8D5fzKwYKZfPYAWD4zODfZnNVuLqOXA0
aKYod0amYxDrxZNLCGe2EocIYN7PXnuMqyovqpBB7vHIkXA+N54qjykGZvqAwUIO
nJ8lJA6bcI/HyqLWSXgAnluHQc5S4pZBSv4wZfzeyW8S3XF9/GFQhlnC+nN83Rk6
USbi6N0G6ElM3tU8TctqvOv59iFEVp+rDmSIjhx+PuhKBEJAypfl6MFJx/XlsKVq
Nq+E5iceuiF3p/Bb09bY425dbrv/NXfuJTRs/JnL6AHsx2/eIt6dqlorBTG42C1z
k98exzvsmdE7zLcfTdjekU0+aUPBdCbeng/gwLjQdzt9MTB3BoR48Kax8yrn/CHx
49J9m9qd2Z8WXT5JgYsT7hzRyaDcp333XAlauZ1nOc/RVczioiEQuuZvx46n6cnQ
KURySSsJxajPmByfs4wxhkElLKpU7w7tA0eBmadFSiE4Mhr4k8x2NQT4pkk/aJ/A
eP+vkgA8w8Y+9AVsApu7Xxkw/BRVxc7ZO/wJJqIgatzLu5KBOYuI0s49BDcdXdDB
T+GV5ckjd+TVxCNNDdQoe/SY3nGk5sUMAhck47IOnSi6Vg5cCPKBMdw9WV/Pfz4L
XoBGKQ+L+WfJ3chFEMjWbI3m0Vj2q5iu9AjLS0BQCAPpCis76GN+mEaJ8yn+XG8M
bGJ3aMPCo+oKX16DGbkAGPSTc4I/7rcA5wTWhgTz42V06bEupD2FpiFZ1yXNMJdM
8Mg1a07BYdsjKQpfbnZRrT1S/+qDS8Oy5X3xauH2BuNEGPeFT5PM4jIHA1aY3CSi
aj7jgc37mMlNHimvQm9R9PrNIKBsvEJ5KHUkse6I0Sqk8bySwr3aZR6LIc0ZpXjD
451gYF3S74eeagoV6N3pddwL/k84g1OpgUr2kpLiV6IHCUg4eRH1917XifT7j0rA
ziKyTBcJgEoVNfHtoQucGXgii37AYOaYn8n9dXsTGY+/Yy91PYcp4NGTXsG42qU+
oiM1mNDrSjIG1eywPVQkbTGycUBwFzzIaBL9m1fTfS6ezhJZ4cqKtOKe9mJwxIFo
SDI2GjfXT9TqFUZxs9p+QbGA5nk5KW1b+pYn5x25wJDVXZEQGI5toBWBAiA/9sdC
VY5UfMttX/sphiDJr64kQ3UdxgUut9rdhPfiJpHB7kYLosnkDuSL0VSjQzGEKLFV
550UUNita2kd2zWanekCfFyfO3Ks+gIt1YSXwzIwJh//jgY9k5fbqlHxDX53kRPt
rnRgQRiqd4a+aJPDl/mzxOMtTdyy8wI42+XZLOJSQyquBE3WyaejvBfpfJUMaHg7
OD4Ah+FOREX6yWH5Ena3KtiqM2UPWhARBIW829ktkqTikX8nVAk9RZpxAXUMNGxb
JMQStW55EYpHRlH3AUU1SrcS+QgtTC1xJVfgD1+uZo7hXw2hwwjbEMmVM0wQe0tW
u9N+iQUyXgo29/nBigBzhAkPzW63GZarQyPCFt5mI6BCR3OAVFMdf+2wJZverCwT
bpw9h8sBEYo6Bys2sKd5b+dFNJBZ4rKDkg20T7sjBdak3HnidVerlph9RmVAXOik
esFXkQXKvUY6NG58fpn4gJWX0jpNr6TjC0lJClNg8pHC/xBvDlGoeg00bZ4AT3dl
M22B9abTdn5h6eGe0mOKQUtX7N5bp2k/ZIZO12vdksSdhycxjtlnjwVpv1RVeN4u
pEGtE8iJfQ+AWhKNJDyZRwASxgM9U8xi/Eh3MuU9qJdxNPhsb5dkHe5I9f2upkRV
vqJWL7flapEkoLLi12K66uLnPi+irgBL6DqjY1JA/WGaMPoexBPOqya/6pcEd/8U
/TfpBV2+TKJE3CoSAZcfHJJhtlI2gELtxN236N3Up6gzSk9pwrSQr4isT7SUvfPq
FdBWBURgfn4q5TaBfe6kPro5f/LcnI71JfLRy8abZwIeN/eOKtKxHa/srl5fqbpK
PtKfk6X0SJrPH8AjQFpwWOcrPXfLYXbrMfVA6sfJFiET7ZY5C2NjOv4XBUeBSPu+
0GeltU9WYuTCuNSFd3qk/+GaWHTOpvfcjFGhWIGA6UZLy+Xb+SqTpdYCOPJIPwyf
vfJOBdpZheMymqcEtrh1Jac4VAzEyytDiy2opCXMnNmh/fPgZPVfS4t2T5BlomHV
7Dd/vHKFQ+ZSqHfZKjBrygmJeT6gy+nHt5yroADblioLSnDKPYz2NOjdw5psa2E+
/sIdlbOfvvOYHNAStMDRQ38IRaDk2OagOoQTf0lLGBg0vjdc8rOelrwfxBUPMFZd
gno1bW7Ff7fsuafcaTVtrEEYem3DzBDrREkqk/pOrraer4bO4hEf2q/0WBShMrED
9WMN4KGIB4u1EzHJPJyrjUr++4OhtcehfVs/K1sREQtg8OqH/sRTE3KWO/fWjiNN
8myF+lnFXMnyVMUu3L81JpHEHlG+Jysq4mlOB2Zii9mwRzt4xPz4mFrN99F9oQJa
yRA2Rl2EuFCN2/VUtgz0b/aeY/7z389Hi9YYFsuHQf6UZpG+GHz6jGSp7K4YY/wP
AjHo4WfTsJWthDIq7bzbiloH5/50OZGwLhYBWYyWGYeQsDEtc1MmohO2Kjxopuwv
z19atAs8SyudfrtS2yRi1ECb+S23SIdIeapuEr6WrT4HXLPS66cpR/y/9580A6NC
LpkswtSKGqaZQG9ox5QAqSyUv7A1O5EeHfxvkFA+ExDduW+c6hcSvWEC8F+bapi5
+icfmixx21/PxZuffndKyQ68zZZKApEphG9vKmMWCRXfLXgnbmjDa6MXioct37dh
9f6bnwS8CexJtf9jdtag2xK1uwLS+qtDeEndQ7x0pHEJLFplcTOpf2UszNUfreQn
8qOrVRxMCce9BXbxhNdcDdMQQkBy8I0Dk4rJIAH9zbw4Y7ozJEydXoTcToELHm00
c1jAJyv8/lrl598ezQ6NHywFOSh2peJNkZHkGmzlagotU1zBpIReK9BVoLOE21MS
5XRypU3X1owena4ohSnshLMDUzpwGymWW6Z54MtEk8PlWLhTlWVaQSTKrHLTeBmG
Z/rdqeGpxiz3vNVSEXRC/1oyDMO+GG/zcQkR7i/KyTFvKNgHMJjwbKjivC+TA6Tn
Jl8du18+AX74XrfMX5qERYYfyGjModGHZnKjQ0BY4JVhtoGgQlg4+kRGO0blV6K+
foS2gkc2Amew8/0ShhoTikVhNw7xBioJAIf3qudV/nZW1NTu7zzEEvdyyauTVzit
gG/yMaiymdjYfBX4i0Scz0QlQOIoB5tF8ARvabtDO7+4Y2TEvB27GfVaNLqocm/M
GjdXd7hMySTLLQMg/WgahfUvi6rpg+81lOMc/NygkvBJ3slHPvk5zNTjyRHFw/so
eWY5D7zjsGSnPAxRimTmB6Vw2cfwg79GYA5aIm3AQWiUI2F3JMUTA+2eDsd090mj
7ZBDM5oKMMGYsfDJHPnyozY2W78BDliLV+MKcsbVqx1DReTI+hsHREruxQA3+ErG
jNMGOGu4g7ev0A7fO/gH/tmQFp9qnFJAS9cWZyDKogd5gQbjjSo9TdkadFnuiMaX
WsLwp/9GDqxnDgpzRD/cS/HJI9IQUHB11VB+v/6iWmaMjHVJs93C90oDMI8DGRv1
lqLPva1ey/Unr3Ijx+Te9rwF74MZqCCNPRYxNojKRHrnuiFJmsq9Jzv4HcdvYWkj
tyuqi74eRuvUx4DDtmMg1EaZpmKkWY2Gm6Ey7Lqby1j3ZQ4hXNjgejBeY4fYIpCP
z2xYsQ4dyXOEDxxVCHALO7BJ9XYQwZ2a5pWi3L+h0c4LAfAnQvzXh9Klv1mHwERm
HHXTMmdJzwNbEX5iWuZqCjlNS4k6VbWDJOHr+Rd85u0GPNKwxIZExaXQqYDm4qg+
gq0JJU6/P3d/7JxX3UdH/DcSnanDagYuphwlQMV71ME6FsjAl4h/1vINDTTv+ARS
IxKIcNnWk/bU584ApOEka7yhKnm9kW0WCCdydijJ7AXyyNHuzFUUzwPRqacapa8J
Ch9cYhoCyAOZ8snfjH4//Dy4iZ/sOssQD4x88I0uYABoQ1nwD8RStolqAWFET47s
9sq7b3KlBmXySYxrbJ5jjn8oMGFvc9JPrr/78KNTcrk41hbkFDWtZEgHmiatvm0Y
0wlIO12N0JNoWCkiRzZ9lL9gLlC3R86IiTpE7O6JYY3SqKaphO+DWioRDIBpQvuj
mBMQKMmNwYhcCVRzMUGl5EYkeGq4aJZSTq5pdO9A5e+OgvovsaU3nklD36nDCBl/
PvBqx8YMczvIHbK761B1vUdgiZ51nlzmTORvS/dBsnTFmFyH5GJqJOB+szNbyVpe
S4k2cX2ZJrdkyUEx3E55j074cYw23KYHCoyTXYl+sopdRDjGTIkBEne1D1Kki8Fl
uJ+hgr9y7JnMPBPoOKpmh99hL45yuM3+wNrkkDyB9IxKctSNhkj6ulaYIkX639Wd
OuMiAZjlSl6aNGMF46LeMX98p1XhhxBKmfLLphyF2NVQPcNwYXGoGC/+tbxkQ7KJ
SN5nuJhfTQeNIhRmbaI1uLV8LIZ600NXBx/DBCZ/3KHBhIGVkV2qU2crO7/vAivB
ULnPEbBKHnSZBBdkNyVRzlXdPb2aFem1wg3FS9/Tx422Yvr3y9GPYbv96oxPHtd8
1rJsj/pnYgSuwnHXh/JUTSAUTFQzkeXLde1KxH0IJBM=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
D2GMqiIxM2vKpKOZWzwj7n4yoqLnllPJUQr2tHI8GW7yQFZ0KTHZwLBc8fol0F2x
M367pIalGpPLRRMF1J4zwzqnmnR5xEoO6WMZcygYOQzG9jSrqCa2UYdlWXnvbxa2
nZaahx3WYttZLUK31x4pGpseR7JcUDk3KvB2HBIuOrC9ZV2GmRri9sc4oYyzEIKS
rSH4Dc92bbZVp4IGyX7lsIHpiXrvcJwtnbgCObHF1xF532IlGsHPaij4OziZ7ibq
KOIrOKxspNnwKVU1L+SiwCfRwk+nnVp45OWJTKzx6HkY0X24glnpfRge74lfVnyL
B1sfJhtYc3I0PngMqDELAg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5904 )
`pragma protect data_block
9TlQpUzvKb0eTULObk3wgT4WJwCqhTSHkNVbicmYnyxLtYxHDDO5LiSNie0q7UuM
T1d6v5VUQUN++ioK4tPaUyfuDj8C58QL+WkpSe+MfxquRdMhTqn8Yc5VdYh34dX2
nOycaaKOojwXQ9OEihN93z6uf0Bfq7564yhAv+pHtIlHw9y1oZ4klmN5yneqQrrZ
nCnp1VhYMCKCjDaE8m31nRIZbkCFe7JbSKgYLSzP1JepZEQzbUlKrmU5QYGC7lix
DjyD09Qd6GYmBtfrocRG9YE0VU6a7FsrqhxuA2W+ht7Joctwqrtq+1wPcMHhPN3U
5CbXcfG8W0Jner5JkPaE7QhsyLI1n63Tsuv+p1X4AeIK+zlJF16M5i9dLTqCNMBb
1vSXQ3+NwQIhA6qvO584sCPSwh6RdU8XFopGW+fadxVMB7eSGH8+wC50to06xbGo
KvnxDdjlKzSIcJ+pXKNDZOyscBQQunyzOA5S2JhHp+DYXjTQeY6ZCPFKrpwjUlMN
QTlz6/TUlcLtks8kzddLGGCMo0m9dmRj3pHf/faicux6fAIjYsfkGrr3Oq2KvRis
kwXVYNPPcCvgnB9CM0xb2JFt8ejFjKhp2PMHWFAYAVSE6ZvDHiNmsHNXsix2NWID
jSMXPItEuf2MWTobk8RrFWsVwxdFoRcwyVgidJFrbKa3dI1QD3M0MLukuY5mXjmB
zNM63Pzn0NPinWou3j2f5Q35+ctxgnmjM3DBcR0Pux0bfbZRBqQF71JhbUdQMdxP
SFpke6qMA9UdK0ByN0wHrxWjd/jcZ/FOIMsiHol3G7llSvDm049zc30mW39QK3uC
1p1xNGjQ+/mRDeWhH9disCYGxzo0uZkyrJbC6TodG5XkzanBwp1E6UPu8SxOsRum
1XLEkxWd/HtKpUVQLOEdDNnHLcCTP1lsdkrSrwlbJaa8f447z3WJtM1XfNSnDEV7
hNjWbDU4o8Lai/zbbrxXXoWty/RhRy0aoU4pfx/DXEE7BzNWi1fggP7hKccxRayj
nUMaKyPxZdN94kgrmbtCfyKY7LTWJIOUrFY3UpAOlIPQxiWhM/72K4IRxqJM2H5+
/5mvZHTjdlqYu+cFiw5gECLR9O5+ZU8U7m7aY7+uZKMzTMykl8Fsfgtivh9dVu8S
Vh/0oWSlUvUlOK4Q+rOSDPul9fyEbVmy7Wijj3w4jIQCO5d7opKuRlJ4jZ8xzWpZ
v/LwJvTqY+4FmqNvVtrp9zsvyNXeu7LN6sOJiNrbh6vaSCPioPTGT9OuswNb0iEt
NHOrqSFcVOV0fd3qJ/opF+I8i8ABaZEOvIA2YlzfzS5XOJfF9SrW7NfdS7gd0bvz
U6AOI+guMCIsuYS2RHXOtmEVSVIp/2hy4+7kh6yQr5aJ76mhHODQ3d/QgMtwfl27
3RCRzVJBh3CM3oazeiEyH4vKiXXiO+346SZGJachbAY997B2GCH1Xoto94cRPNrr
OaxuXTjm9L8dl1phKBIb9rWvFMgFi7mjoxUsctZIPBdFi+s9ynYj//BMEQHzchBY
brxx2rueb9wSECjYLh9A6gvtXYFxqbtpOpGZASDYUJf+l2/AAbecv3hGOHpj8vvR
fOTKXzQcGEmIusIhzqXo9aRdQSVMUpXZxPTSalofgSeMDH4pBu8NEXUocdueBObL
NELF5jnKDjWgUzszVbwgmLr/5AIDRICdhtJgF50jDo0aMxC5Av6jtINseEtyG1uL
AMn8yv9fk7FrG8mhDh16/X2McFhecadgV84yzubdKRkKILjLJG3KoD8WvowTEk9w
P/3yHHxpJC+/EzPTGYBbaGw00NX4yjl8Nx624AVOv95Gv/2JdtSnzYeTMwtOXr4t
kseCHqnABb/Wp58wniwZ4fv5mPYRoXy4igLLbVxigv/ao6Ud/dS6feqKFVaA0Ua7
lFPAFrjDVPEuX+WRXs6W/kAkB/eU3GfDAVvprfTVeWSktuxaQiES8d97iV47csf8
kPRhHLXUHa0UqklPVqdfTK+Hc6vA9657g1TwRImj2a8jhCXPcejcykIL0e9tB5yU
1/Xl0cgYtWjCN3SiFPLd5daX2Node13A+6VpdHhI5H3Qm2avpF1YbntYAWM/UAUl
hmlt8DUKs1LkLLalT1ilcCdxMzFL6p+jWkF1OJceFvoGOM2FenG3OFKYi3EZfSb/
2rZUfopxs68jQhcdZwxrDa5uJ2gunjgYpuIRkQ8iq4Auyw8iyz1OU0C0llPHkyD/
MaHc8s8XAtPlJ+MWD8GdsQex186L2wq2Lfr+0hIMtrvU7qbjcGRzk1MWezVp8M0J
NF/mFCDT39i1Wz9ZpRLXyrdXIg0joVwD5HWhADlk4mh4U8GngG11SJG6AaA4cVjo
Lf6uCPjPpcN0vS1ev5KwsHLy0mpT8rKiTFjfxiDXQTPxc7yjBA5HBewy3Y9ZvHVx
y9LqSUgWK7yyv2MMQqpD8mo/k1eU1HdxZP5T7ZpylvH+f1kmcEljfArOUP7ciFcq
8Q37HMiN74i81OmnD7aWhIEjCrMtEihR8UgNsoGyLTgtbSDBnbIj/5hoc6K/Dgpw
k6V8U4DpvoJEaRKAWaI7pB6+eXxVnuOYU/jwMPmZi2GnFtW4piEw7Aws/lTjbyPB
HE9CuEvqVFACXF6/U5bwY3IWKj4IAm53OfEYp3zP8yoypRkB8RHmQPr+i3IioE3g
1K5dcd9/fUMEFXYazzhK8fQrxrGV84/rxQpGB4e6ENBJYuIidXLFs5eEq5fJmrte
jnooUHXIPGfonFXkJQ5FwYdlMnOk0ZBMrrNTFapLGcHuETdBLCIwOxoGByz65/on
Qy72FXd5gOXdrFnKsttEbg2bdBHG9OiG8qWeFcNw2/dmH0UmGxgcCNi1mXRYrFqn
20PYzHcw9xxOUmmPPW2dvbg1t7ZsLvZ874bvBa/0jkbOi19K6+ha87+0otB1KXB+
zvCFKsYQF6ZgyyfP/T9h/wHg1ccwo7fcSVSlU56U/Gj0vFSP2AtD/bBG92SymQB2
oJobXbJVw2+PIRkOFRlQiF/11EnMjhAu84gp0JIyuxNDK+L4Ee+YgnX2p81+8Ssa
p+omzhCka1ZKDP96mPvax76xufVsLME6908UgSDzhPLXTxDFof4t/YeuOMO4qA41
4M3AHmOB6ZBOVb9YGijrkp5jgYdyD/+D9bFglDhosQDvRi39cVFFcaenABFy5em+
4nlVlPR39qVmHinli/1Ye7rVi+j1R1Dg/G77jmR7jNthPnzCB9RKn4IeX3jhKWAB
+IW3Z71iIjkpl2+dOSQ6DpCw8et7gCRwnMuO5ATTpfpjEizwQ1XivPT2awG2GKLC
38JM8GlwvB7c52lo/hfxRUG5taRgSjuFezHOcE+97y7c51m/D6QQ9upwsjRd1pAi
ipXvJhpcCG9kGkBzZEpB2yAvSYAzNDQcDXKKLUeUFRzIRG0rymD18MW3gV7rxZ9x
/0KxIi++BLeEa3cdXNp1b6R6sauTQYaS4QY0lFRKiMHoRHYxWppAnn84LMiJ+Qit
hvVvtaXKbcgn9JBooWskV3bM5ceJEJ2wLOZB+gpksr1R+Ftix6n0nnvlLuoB70h0
ZfgMhcjAvMI+o/KFFey7DzcReOq7UMSPc0K/ELmMC0P8ONPT40WRIFrB3yTWrHAx
rFEtpLR4i+xGZk5IzM8pkspoxW+ZF/+6K8m2FD8CymVcU05HaY0/ccS7pcYPO3VQ
f8f2THS+exFKmv4iLSWAqy51jLMDUYirquEydR6CF9bPHtZB0nsnI9YMJAQHzynw
+oQ/vA5N97LM648LsW572lMWuCC9N2tRXLCMFDaQ54VqoJvG0R0pzfUBIH2y7sbH
FCSLg1+WDUnH3lBGg10vTK0K2G4mdL6mduHqBze3iPARWfKhvG+ym3RqhVI27KN2
aqbX1ESadoUstpuIonD9u19+yhirRs9Xcql7z2sPbf5qjzjeEP0rGu6rqnx0CdLI
4FdJ9xazxS/zHurCSP2yUotrZjxBQ/bLpz3vSVaaLoVWrjtX+/HpIB3TQ9rUAJql
f6kpTThoQSKjk8/CL6b8iWz2/bN5xx6R+LeA86MqGS51b9JyYGrpcoVcw5Vq9LqY
VmWhOyBctDu2veuX2HRrQVX5ZZ845y9PjdPtMTP3kDpk45PkaFwT6AcTGMHH9ijO
uDoqMcEjMaSllRp7EiXDbno0fDF3ai3uVjO4eaWIQZ/J9lbvz+WO9OOzKA6NxYe+
BkoRnYPnwOho2T9sMh5eDPCEJ3ykxmtvPbzyIFQznR+SAlZGCb8IuvAiesJtd+NG
Ub0S+w0dGJ1SQb8dDw9F4x6VotuWDi2H64qXUyHHZbBEuv/WLnVEDcmAyqRIEjsT
x+zzT3CJIbZpvinUlIe+MSgoO0GyxcOhrgpjdESt9xe2ifL3KWjOfOiwX81nypkh
TyGpdQbC6dj4jvk/kTdVXuJT0XXE6kyEyvrJ8ABz4FKv7yac0hMTqTUKZ4HN2CCy
U8l1LmcpcHQGKNcZTLdHutyJJyuxdwZcEYn0vvmgQMzr4DkHLA7p2iy4ImNvvp8v
C5zNzoNj0ewiUM0lBPEdh+tb7rRRiOgKSzhisRbbz3zGiP5c0iUkRwEvwD0uZIxE
hfuMHaAuIxLBfxy4/li/ijdvtS73+5aGDG8nWP8nqJbQkW55XvMvU9iOHpdkeI3m
ujp8pyF/EOB3z0ajXB+fKoqZoCN7x+RBotMdlc25QuxK1nye36RDzy8ntCqCI/Bq
YIwRjNdJUn7mUFNtmxzcCc3TAZ0yBHsCQ4+tKGbfOXoZjCpMM0OfdNHywgKQ51zA
9tKiL2zuiRNJEKhH6+JBr093lhUPfAjwFhIBZZUNie4pkPXrbOvBfGvzbItHkZHD
wS0UZg15Ymt6+W0YGtjrrtkHUmAm71zW52Eu4loPl5rLsfJTPj06dcHi2AwWxvYJ
WVQOdcG2kC/giXf5uf/a5MhkAV/C7W51w7driQScMZQmmi4Bnrq9GZ0dTejgdMTi
jv2jutrMp0eksQMH4riMjLOw+Ki7ZuWcU+Y/YCADeWyGH+praU6IrJrMKDAHVV/K
gNQ7Ce+PpSdVbK7tPDmMsRcNt5E/EyNTK4ipD9QmUZ/rHFTt/Zax0hYy7KREvFhW
XSdkLLsU4rQiGNCcxzrUaKMFfxhbK8/vPZ2yCJII95dVwyDQ8ujvmCflAid1UAQQ
eEOz2I7DOm0naYS2i/Cz9iptHfX0PcLek5mJ920cyS72CARWOvwc8GPdrq7MGQp0
n34nnhNZ01z6k0bTLV61qJg8pUnxA4NK7EFGgLX3cemoN1u9nhkHltXKNGdXdVG8
PoUKeIUth3rYW0EbWtwNuRe6qEtoRkzjGupq/QDJOMGRz1P4RF7QMstFy4Ql0fwM
UDXjEv1004XcE4TkW/kpPODEihcReYrJaNOuE9LCSb1/So8NnzzTboxY3YMImGwW
rYcFTu6Y8H5/BrrE6pDPQCBBqVhlWo0TM/x066Z6ft21tW1WVEn0jIS11YJ/OqD5
+vqaha95rcikvkfWF6WuY5bV4WnQlVEiXo8m0hSlUYP9EPxhS0IHWV7Jnp5fdL5q
wM5rFc9QguEg4jtQ2qZX+5NoUVVBm0W+A025AlfD956mkyU6gUaoVlOnPxR5HlzF
2r7ugPA29cpD+JeKU3XGy+KX4NoTCRX9M+oEZR8w0m/TFdwZpMRDbim0/Ukhpm8C
u1bsPg9DT23wtq85n+wxqPnhjvsNaI6IaBtpJkOD3osxn90suNGi9qZr2USTeewP
LcIzxUBx78bpmFlesHG6Bq5jnnxXNqc16Px2UMR45YA3wVbZ3IHAqrN8yUqPZ+4Q
oWBpZ88IUJonMqi/ogPJ6CG7AzWy5F2ZyRPx32Lj8uYJQ/CktnHGY4imm69QzKOt
jMHtJSutR1kOCAOp8lu4K/ufQUcOfLWvL4gcPSTm1dlSRlULi2FgVU6Vqk4FRlwB
SzYrvyXYZJOYyvsD+emAdc1Wq2kgitnXnquzDKhpQutYkARCioHpcaxdope7VsHU
nyaZ4PfkFvYkDkcwooo7CG+LRrU7WKS65vpgWicV99WynxSPAvD6pvrN9VLmsmTM
fEqdSpikQ0oXPxEI/kFZPKELKCxQKMXAUSpWbAOxtBY9Wqc2Bqc3OEpM6dow8A2f
WY/YE+ys47cZxyu8t8zaCYbSX//nfBCVLZ70J7pudVGQXLw3KFzaLHbREHta9Y9q
jvvqMHXpBb2PS+AmvFyo160RfAP8pV9kkjIa1/b1Eb4O+D5GXVJvBaQbVRVbCB/l
gkqDyHFv9Y/J/5LW4Bl9G2E8/jhVjGvlL5VVF8A/XqjmNlVhTTDu/mnx07AifUcv
3kGccNRemQN7rKbE5vk+UvsmHGOzMGTGJlTyQzWEGCCUveFCJAdxHuOerai7e5W+
FMy1OynMGW9a4w3BeIMBVV9tCb71sk40BftwRJPRuh27VhIpguH9IGze/4f0SoI8
qxNE+5jyuTm6gHP23bx3+AR/vuyITfEksI/j7DtSMOjb1srtwm4uQV4HcV9rGV93
CoahAIFAM6R10hMcJMHZWvma1km/DRvd3n7gWZzgqZyiKPpgLmMpaJvGy39azeG8
Jgo6ORmsi3r/kV5NaNLy+h/SaMwzLB8Xlnm9lBkJAg4p4RTXt3IdtB3rH6J6i1dF
z2yf7RJMpD+mLmvq5W9HZJex37r2YTVMaHBFL8mR226uCKqKFzDYYDiI2pxtQFgN
npxGeXdPxQ/MYcdyNqI49q5Yyy758tkSJlODTBr9YD+SKkWRpitTIo6Cq2jmnGme
+Fz+SsIf0g2eMj9zJeRFnMVt9+VIijpCyJLwC6z6dqxGfEPPrNesjc0EwfnAoJSY
4zh993JtY8tmyZPDIeGElufmv0cq/yLTihXPLPoqSX9pQBgi+1fpoXy+F5WR+mQH
2M69TU6RwjA+hyF93gUPQGmBKWzI48BAqQcgHZBYhShAEeeWuKQhFsAjih+uVjoD
Q20pHnixpMR0QwAG1bpxYDmxMOIUgxDXxZLeaIL7CJq47D2w5B/Uz0iIfChyniU7
BwhsQgWM9jMW3g/pTmX0Us16yKHNsc9TWN+bF+xMc+PeVwlz9g6vVxB5TraYmxEm
V5FmfCq5Cn27d1FtvX+Xz2Cvip88bbc/1sGk4YlihfD3b2/QpK1oHBeAfxYXnGd0
fwKnlx+0xE421R9DKZmc2NI//EUkx2bhGT2kBXH9s0r07oaHmxqzQvv7rdyKEbca
pVn9C/FDp/ye8RE8PlDQ3IH3ElP0FBgJ82pBpcXxLR/i+oJaTLbahd4yOgPY/U/C
ujYIj6JpPeahM6TXsZIxf4BRSKPLSXWZVsml6JX74bBJ3xFllIOuYX5wW4C7HM62
XWSts64RtEfcjzxUgCQz7DaGPJhK6M1MJjJ9OfX8szYF0tuV1Xz+/1k4Ns/+mi9Q
je8u2boiBCEKjS2CXNP9hD4fxabWWFmP0RooRg/7amSnpkt+5n3Vn7s5YnoSpgkW
Z8UGuLmfaPBQCrvTdAZ7HBIFHI8UM9pjx38PrP9kRCdIwp8E9r2DNFVl/1SViUG3
JrukE8GdJY74pnecpIiWUqIKK81xOdgHbUI37vwT/VUF+4y94qcWnqzlxo8Vz4Zf
IlypMFopduvwKuH385gvoviPg7XhLQKqJWuMCZrsmLMVMkOMR/xktGck80oJ/xSs
AVDtKimbFiuqKnVuew8yfaLjXF5stfTBnmbuNFlyTNDm7LO/oAOvpnYPxyGl4BtO
SbdMAfhjQug5Nxc6+vanhF5QPhxsjNQYiy/jYCBJ3BgZqk0ve+TZBLAm8xg+U72f
ogc+u7MBGBQrnald71gy5EMmAqVCMPfMTuZ3+QvXxBmzBdY3hs7wFeA7dpBIArlZ
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dUqpES5eJX7Ky4dH2o5mjn8yCqWPNODo8YXi2XmJ9cn3mq/RwVSMHM889Te841Mf
+C9PFVq7UFeeGrEJQuMDrSGH193vdDlBmooOV+82UFBiztncm+OAGa6VkvPl+edW
1sUnzQg1GLXTt98+MUjHy14GwI7mYLn13dgxCR/iKeSVfwRIuqqAuI29bdOAVGSA
goKIgcBqrPJ4dLYjKryXZawity9VnRhHQkvIkb/xU3dIsqZ54lWlL43V9FCodtAI
OhmZ8FWFfszeomnCOpv4Vt4Xs/6yZ36tvlV7hmjCbhqb7x7XYucVV22Y+P3CDBvD
9xIANHc9xilBuk9mmXOpfA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7936 )
`pragma protect data_block
/b3E2eZtMjC50/koj4nsu0cGGqKjMAVS/H5AsLFjD5lFn7bSj1gBK5COzTuwgik8
CwRVK0kZSSfcxcjzfk4igi818OwskAPXvzJT0FX/spQ12MqpI7BQMjYCXPsCFl2X
8Gum7hZbJPrqoh0TY9SRyjrZ7rxXpMwP++kvL/BGA85p7FmVCUuMbv0Z6ncoFb6T
76F6MX+3Xd2y8MXabmyOgaUYrqZSaU9XnXa9n9xv7f4dU6oqFbjhBZ2zpGKNDJYz
148Ml+xbipmTtyMtCL9VgEXy8U74LhkQ4wxCx3oaK3lc0XGWQDecN1ASk0Fp1eKV
3XuhOP8lTUzJxsvMl72EHLT6S1xR2wRZPmOq/MYqVvd61sO00GN9alLO335uaR1l
17nMwsGjQJ/HRObZ3Ye4uUYFcPWL9RJ14eypeNC6vCJt1ZRP9aWXugEcSGQkGjFl
Ixt5OXmgj6HHilSL4Uopt2u00Kk8VsS6e77hEluIgLQKojP/oDAxo3489vxReFEg
IZgh2q/soH8twOk/Ia6eCzM3Z2M9nR/Rbmfmxp1APLSg6pnNnHekOa3IPZPBDVWv
YanRGkgG+GndhbdwKr4UB/TTbVgFxI1GxMjW99BfysgRwlzUkGqkTMhwf0tGW3xS
on6oviPnb0FpqmDcIUtDKFIWFvs3/BzHiQDKFJoAIn+YAeg/1zNQRVZwTyStm06Q
SobuxVtmEdHWcuHvBRUFsJzA15gPApCd8AlSss67AMDMZunzB8LwscyKoTsO5yw6
J0ldPLbuhfGt+Juqh77EBzf56BH+W9+xwPZnCtvPJRAKGSwUU2YTN4BRyRrAJmvy
zlF3bBtUN2cqq53FBsnQjZOnFoTFTEQ1ZK64lI8z8vzs/3FgP7aPzUmjfp7mTEcJ
T3JudUmPbc1r2JIdZM8TxHuw3rhGbHccNeUIu8gZQktOvQAGMiQ8b5ZJ5WqGqH0r
G5jHFLRbReb+WLvm+TUyC1oaeYO3VqVykHDk/oD1ryyXIhjFjqOsbPwJASZ6MYOg
vFi0jvDT8mR3itdUugLvu7DL3VpdDq5TniRzkX2jnZacb6dT28RxpZmIVuoGM5Ur
YM18qqxDjbBw0yIWpnUJy5UuNaqHQNJod3nqbYm0k3w1Bwkyr+uKvRSehBnh+BlL
ZIWCZE2ThjezX/XuqmfHBeRTTClJ43bcze/id3jZ2rFnpoac7r/ozyG6ebzKIO2+
danhikaUxw3zi9NbkioXU7GxsNU+taKll5LwmCMvvPNPa8A4ktBNC6GJ8l2pZZA6
y4IcaO7rMJ3EeRlixu9qjX2iAY5M9xWHl6rX6mmKkhJjj4b/QCqYftLg3gtVwMrF
5b5Jth+HtOt4RBKyepEsh0d4PUDWk1dN/Oc71YeaqYkJBiSFSr7N2gWmKEoRQhu3
5yfXlD9WGkBXnIbG9aREEfUdBNCGRF35qFexVDIPLszlvq/qBIU8wTBDirL2FIN2
QJuioFMSgLK4eP8/52e4VwDKKNIKLInOjKPlxWwfeC5Hsa/BVN1tf3IB6I752oqF
bML4HFlg6vcpAY1SwL9JqXBE3FWAjSHDBmjF0bgH8M+W63+JDoXQjYvyDsxA7QUi
wVVtBA/56e18j1kgo0qQuaNiK+P9x3xWTZ88n56EhRNqvkGzJzMvvvq9NtwXo8/w
6nwICckykI4wYHQZqjRs5HmJOZ01lOkzyxOqXXZ28gzzC+gEnZab609eMUb6w3N7
DnVM/+2fAtKjhLeOWtXIh1lnPevbVPi77FJvVgDiqNnGeobvvwT+La/BpQ0tSRgK
VXFctDsx1UTbGrgTnrn/vtzBC/uQW4kWUxU2jtM7rBd/470wJXZh/S0q11A5oZe+
q78xvjanWCySRaFLNM4/34sYH+dJ5IQUWQSdlYBybUQB35tyvl43nTKdDfPvLPR0
7uGvJltVHaUPe29qxUZcJZFbW8JInv+wSy0D7qdajOcCemA22CjffAczj7IdOnVK
3tJYKPCatvU3IoFVyBKZ2yy6sD43z0gCXZyEMjnmFRl0qvfj0U5xsLwkBGobGSJc
BI5lkjT4km3z6Qgqyhh/JsXcbcNhp16dG3mFc18oISNsj54VNJ/J9w3WDMQifXap
1SWE6aA4M2h6kixo+tBnbNA2N5TWKhz5psMKmT0xZHqH1a90A6WaLtwFGIRfHEYR
ueJSwJ3MjkuvVzO9PuuzmPDNNatY1Rlv3ni2HMEriCWrH4Sf1sYeWhtwkrDuCoPa
NuaMf8qlo8apVY6nVcFAlxdlBD4C10g5RECMhB9gmY9GlIHnjBKgkh/bQ3tbWAtM
ruPoe/KfW911Yfd6hxQZ1dBJBXGV4EY8B/zXAkaDTeM1fkULVZXWdKbzbGfyi4b+
KcewIPBQ66qx3/nKrvdROXCVwTE8f/hPb8N2PxS1zvCHe6AYdPagMtWpHh9ET25O
q/vCu3aJ4+7KYWRNKgBiPgaO74CYc53ZQTdz7xYjFPBTTSPREwBjqjhy+MY2g7xT
4T0fJFeSh87JbSVgtNFjdC/LKYyUTQGFJzyHhIj/qbKytz03pJCzyKneNL2zLxnD
7pwqXDlRHfNfgsd43+hD6kHIjjP9KaqiF8y+LSAJYurX6kcMITn6zTnpb+npR4+d
/F4M8lgP33jr1ZOFs4qnEZsnbxjfSYe5W4Lfgu5o6tyyVuVBpbTQ4gBhy0AwgfEs
+ds95JMA4KnhSm2YIilbc2SvuMe2hs0FfsNwl8WhrzhHpQ3EDpVFVQQKW3H5aT9c
7xFdhhzJvVngCXOZQNvBEIQtbEclOFFqklC88TdifSvX1yIEXMy0Za2D28epejXU
0uoJUcB1HpC27N97r/ydAEIW5wnQ3yHzQi18Eq3W3wnBjyx+1jnyHxHE5JQIJj6+
brrv80Nz1shnhj4P6m+409cQiOJpQX8vF5T/IhmcQ8dAusAjkukt6BnnuElrsOMf
rAGmcELuXlmSOSamialBidHQyrImVa5F5cj1o87svKK9bQpoZvOQMD45m/O7b38o
xTGfkeLHniEyyE3Zc+35HwNeuy4sLxtyEysXIs+6ZZ7bPtgsLY+p+S7jR2fsRfFW
7u+bV3fkk86r0S9bbyh+kGIU+P7pQDkCeE5/54yk17JrRDk6g3Ytc8JAmAkx7s7R
dTm0A00yFKck8byeS5Ngm4Y11xpHn6fePVvib6uWKhZo6SkQeBcZPXHqg+0RMJT7
+lnZOpECagSsjx2hCG7WxGhvkWWDVSf5RBf0Hmw0mDrXai0p6PdIbac96nYgVNnh
KRGp/ZCykx810KxMu4un0Q/7Xcbpl5ue1aF0SYibJuaefaOWsYK6Rb979MfZJqZ8
s6ts4jNoOTyhlh9KHPEK97bBzaPhsySW9PFYmt1dutR4kMq0BMGPn+EKnDonlj8v
7het6Ti8dwjiVU2K7Q0F1o9TDhGzpc0+7RkCWYKO8xrfSZ4H6ol/S5A0yW6Uuu46
/LqNn+WfYadgc3oFOy01Hy+ddPkSbDAZgLOWGSL5GzSwx9X+BIOa8kC9kSo5frjt
w2MP6ZV8pj5dLb10Nyr+cP1teRACLDXQGYRb7NJWznTdv2ybQD1/TlRqY9plpRJ5
s21kpWKGuaE5lMsBqYknVl1efQ8CPxKcvK0FeUV1ety2qpXc5J89a/zolecZxlNi
F2uBg715raoEllDLyE9SB9jDEcoFwC05NqvarwfAzBT4LcBCgN2ndRpMfLP3fRQd
jngphp7LMaCKy9cpEH5w2yi0uU6CxPluFsGNXEkSLcEVWhNjn9PSkk7WNC7RJNQC
UlnQ7VpdBtFGCdU33ljk40DbU07cIauvPVNvcnDApHNhn539YtQspVoBZjOzU2j8
b04dXR5Fk9K9KRKXVIGT+t79BHEPCCGmev+ffc4tPOvFehvMRey6r4DpwB+nQrGj
/+5mbMLzAj/4Lu0QLXOPGGag9PgGq1ROVLt7dPXp2ghIabSAwpXtOieSJVDxrP8v
Xna0eVwM98VP3nickYA21sBbe8bzAQ5rHPPanYvZGrt2BMnmajDloAfvZM9sWkDP
fyTpMM2eF9Pl8EzItRb6sS3A9WwXLRmoGBB2K4ggwMBFFm7RlNCvrdcCsgHtbyJl
SIXpw84aENJw33f+fyyGz4wGdCgmNJfss2Txa4Xwj68A9DpDFhCW9yTVVq1nKybx
66TTE7W8badaEhfOkpGU+L65ubxiUYV0ZZ9p8k9RKdpc3dn4M/uba6/sPM2ndmf7
YV2Tairl/q8PJROIbgurW6JxemBuDHaVLv3+8ipIhT63ikyOv9+fWBE1aB4k71ja
qNqYNGM8k8OjIMcUiChghj2kCa+iX/Doeh20wIU4ziL5MAF3jIkLAHFwAn7RS5yY
dNg+lNDPw23fuziD6pWusxJ2aWxIaJu2MPHgkbnLoBRuw7BzTOWTtMtwnjvoFXkW
969bkNCclpfxpX/POZGN/x0QlW3r3Xflj0X2C7KLptq6ajs/3u+ZKGbykcNjVdNN
hAFeAT3qtPo9qoX4AP/db6C+4rVFRsD0ZWUu5h1VkKLdjfqimxkNjKf/JIf9ReOu
mTIBmDcaN1BSQffaTa6zyu94WvDUrZGPunwzP/1CIYz+i1SdCFrnJ1IpuTOYheiy
WanKttQuB5cwqWtU5qKzRcZaj6IDTsr5+OePaUP0tF+F764B7FAKyFlj9NdtSmi4
nuZER1OamgPhKBwxbhyN2biipU+5kkwLC0skIXGKigadwZJBrCfqK6lVcarxx1Qz
vFFf72N/0TDYgNR28MXIW1pDubPXLIuL9SXd0LXuvJZEpBOZeJyH/fQGtMB+Ejo3
j74ZLC2xqzPASCW20ZQLrWcbR/Fsg43oPvOveKcxdfl6j4dNIkc0muVN1pzrBysL
N+nqcso3NHRKll3XM8LSki/jIBHYndFeGXkebeYQKiuB//XAIbdwXbMHM7EDWYoF
60FlpPLUlnRBeq82ZhPmFj0YzMnU2jurVEzY/nLR/gCllZ/VaE4PypyaO/LRcbsy
DHvfZDsiNCdoosXZtXVnZ5hpgDHxMz2TD0DRPBdJwp8SBpAkpVTEjYtJq5zbC0vL
feYTdXyXGkPuotolvRglD3pqGaP/8ybxiuY82qORNYByqo41lBBhcSRI+NYrtqIk
2obu5WyKLnUYkBVMEXQUpKafM+ehV1PBgDSr2P+xSp7s87y4h2M/q6ab+m+XVSQh
HWrr5yuxg6wcJBSEQhohGZcf7rLe3kLUZhlpk9FSJ+AZY16Gufx4Zm82dyBvg2bJ
egxxE0aNtE5Z7WXggwZKhLglHHOyuuSyfg+KrnOjVLbjvBr6u4R140XJhC41STNp
n0YoSBw5YergdVaokyr/v1GyYJsgK/k1+LBtkNnkRjG6ngIpkWOozPiNXYQTzXV5
d/ZzzIa/y2BGLAhQk/UbmHO+FHk0ABpXLkj/fAp2EBOtpES4joBQUvAYzZnAkzHW
EoJJqXkxFRea2osEU+7XLcaB791FWsZdoIl58yyJ3HMMY76Z+XChsy5Tw1QqN/3p
Mba9O3xvawRL7Yx8H8B2Ay+Rq49aL5vY5xaVoz0omRYpQsTRHT9LRqdoX9LZEfye
Kw7i+h0t3mXo214sazWmDvtjsG9YNqvsgfqog413Tm5c03jWOD5KJwNVVif9tqR3
P/7WizIkIhefzYRLu9ONpy8zQWt5OEbXaxOUtaoMSqjx+11GMzRpLS6zgcLH7SMC
vNQCZmJrc7pV5UU8LI10dyDfaCZtYFs8b/lacqQJA4VXZxGvh7hDrIGq+q5cnnTH
PUgsemUm4xFlyt7SVY+gbDyL5pSmhQpXDUZRXGZA5ZHoGaP+hg5aoLFiccu5yR3h
jsmdkmOaw0pCQahEtkTtZ77QWr94g3M+O4/tlfiUdl1sXtrb0EmhNaEHMkU4ZsmW
PSTkJ5nr+l0MmzFeiY1wrZbUG+fZLZFf7CP+NaEqGOSJQe1zK0CDiDonnJ0QTkLC
Tnw/IKKOq09VCtaflZ8kLI+MBp99EO/ahmVomdTvtPcJGIoEMpTIZYsdsoyWrZi8
xozkd2A5ISTG+KVH000tBEMTXc1eoeu0R4lxdwm73Q+0QRVblqsnAmDEMvcxV7sp
5PMBZCrN2eNy5WqRJaj5fQ8VP7egWL0w0S1IibYKVdHarwgcLc8HCUVVR1WlZAR0
iW/7qrNgOsCf0VhD38A0w+A/GAubATw3PG2boE8CCdTe4eu0AvgqtLYulr+R4PJ8
xvBvkhliWdc4x95bQPJqxd+cTKTBlDG+e3VPNxkPeYNVEzjrkraC/8W3V39o+JVJ
1stNPJnXmbL1jwtJIxIiTKCozODvGb1r/Fv5Tw1bi0tVcZcFCdxzFQUatu8WpcxQ
8NRYOt4O5SpCFNL765du89gYWjb9v2MELty+leITP/M1p4hrOWVa8oGAYpUbxXSb
7sXWsP8at1j7gXsm706HIw/45P4gvVzUX3m1DiYAANxV7UD6UoexXS3AkDlHm0v8
yMChA6jW+nrVPrHQlmEqQ0f+A8Fzudvihf32hvTapPdIQ8jZ/KFWUUYKZaXImJ+E
46MkVYCUKq/nkTs6QmgABoZ7DFvDL7hKdNbHBpMSVIfgp55Jh/hY2ez6kJUxD+Hs
b0bvXYhjCbRp8y4ct5DnZO+uVjIvjSM3s72dsuALcC0QIt4VVyg3vIBn9GgR5ulJ
wxX6yhPFEtTsC76cB1fLnWc/WxNqDk+CAcHSqlWysmaRK8oRHf4p6NWbob7wK9O2
tVIX++VDopRJQ/NeZ4ZSCKlVcKG+5Z6KoyEXwkMsnLEjSioHsFMhn6eYqcVIwrgR
FwcgzT58Ff0eqxfX8wNiUUoBVSH1OYXsnHjeZR+s1hd84tPkLPWO8c4+7rvMw8uZ
do83D2ytidawYd9aLPYBoxkBL5rj4u4T7/MrWTqrSUHXptD10uxR9JglemPfGvAI
18IJdx4y1w1JBT8rnFoW1kd9A18bevk0UH6tSyPwwwPgkGTwQY18Qhby+K2wY9Nq
IsTob6eCUClhieszZcT4/tQ9qoE4TxJ3ES0mCXTmOAFGjmFbg45GLBglAEkIrYrd
p7x4PSg467TDtZNs2p7HgJW3O5j41D1tHwTzIMHWdR6cyH7yF8bww8dmeaSHyQ/p
4Mlw9nj0fqwG6+XMONt4cRXpMgpmhSGBJ9HUtredUgttxGWCb4kARUv/BPck6nS+
AiJK1GI9bTA2pnWENhP4z3DhLh8//d0Ac6pxqetPY9Km1i+NfRht35OkAX3Q9/g2
CuPxWKdOSGlS/IXz/y/N1U1t2cxUnds/M6a9Ip7BBENze+L3LGctXfsFoEuF0Z5k
5kM5izuZZjfWtZxXEkHI1SSSPmFH/ZHnZYhZC81PoYc05cLNbvj/1bqoxuSz+Kg9
iEwrot8SIUjU3cNR1zLFP2625AmInezu276muCuTWGsMuf/if0lNBP67KT2dNxTt
0YgwkX2wlBBvHQdtgsQy5uqqP/YR3TOQqlRZQHnymDD7sKQY5M3w8xfhz4Cg//ck
aIUecn2frg7s1OzrJFPwBPUyS6VNAZp2wX0ojG0fsJ6tJyGiNj9ASZSQraqd4OUe
Hlprlx7lRKC40v198ZMlDzNUKIF7zVPlaJ7k2CtHBOMn9c9nhgzQsRFVwAKqjcbt
3F40YhmznrCJkqjTN6HE+WaumVWnq/mJfReOAvkyRplLOnWgtu8wUF2MVQlrGHx2
vSa/iheZkrrKL7U6JtNG4lmUrQJHxrQiC1CXg/JjQBOTGxEJYCtWdIq9lccm2Tx/
b0dtTbkQpApEqvxlU9FMKBGsWOl7htMxVs88M0EcDh8WvYY2uvVR3XyGMCHrbjOA
ft1O1fXhxlIQLpjfkunHbhGGkzBiL2WYo5GBXqaL0MJY75yMi2LBypvQkVhI7GWo
xeSuIygbpxkOZDeWnbhXuheeP9+ypVeZ9+W9mJXZ6KaE2zJa4ZGGpuilXx8IJgTb
b40NMibWDdIV4BX7e9bd69RsuKrOSfjwRbQzsI052WZiexwZMRkCvpBTB2H5jkT6
jIArZlOtOzeAPBDofhGJiecrv98odHyEMj8ejiRh9qL1nbCyn+fCvM6NcADOj407
dWPcdqNXMIPAopqc1tUhiBnvfPPCINTiLvyif2BZpXClpvLN8RIqGI41sebsTuaX
gbLBYPz/mlO4/VE741hcOByJCH6IN6H6sNx6URGJddYLusK3DDRdmFKG9QUmnu8A
3LhUV4dyPweE3eil1YR5uSkNv0Jf/9WLvjyxjNJi4jFZSioHkc9yMKezAG82G5cC
DI9b3AIRGcPoFyxW0SDfoYBfV1YV4e4hdQsnAHuIISdaBxiXRjsjfkURclx4snQr
hOyHgvoztP17p+wOkj/Vdyk34I9z9X6oPxH/Fq+2UWdLyD6REu8qDTWZrQppKu3w
Fr2GnNDuDiBZRa6zf5l52IUit3mzT9qUCB0oOTyrtDy7/mIQoauWcWINIDg4oLVJ
dh2O5dopopAPsT3ERj8Howgk6WaXIMNYO7fizdC4+JIwi0wbyPnqjGSZOQc4nsF/
6wGdtayCdmrvP1aR4pa6NqyBHlxE1aU2rUza/QyivbcTBiPxGbhXxcH+aqLczQsI
GL5vr3kyIT6xv1P+bSe9ZR1KpjaH3YWV0BZm/0yucsxH6lsEqlObQsVw2bm7v22v
NJ1eQc1s/KPcX9wCiR8Pp08CZA5z4t8zvERW2rcYJfyCuzpVKpRGrJrvIgfIBFmG
Kar/0cdHJ9Q4uG1eWQX/6IQGtd+JyhkHS5fbqa+63PQAIh8gYz48ySbLcTgajzgO
pL3pE3omhgvFvZLdqaE8YcJnSRoVfR/U1qXxHjiAhzoLi8E4cx9oEXt4dSMLsEfZ
B+ZniSV0MdJbOvl/B5fjpk6HxH8pF/j4/7L10NjuR56vK9sZZ+1c823iiftjxQax
h9D7BXc1t2IvmI8B2tJ7PIRJs0cH4KdHUb6+peT0KjSxMl6NolTqbVSOZTwwTv9A
ILiV/3E/dmTpz2xHHNk6o1lj/Mtq+pwG+pVck/ye2UcLWrHkyVBEriGR+PA4y8GV
Ayy/jluH/NJ7CCpZrrqbTlYfCmJgyoP3oAON3zOlR4TqXIlQD+7Uu/5rAIYSOAIe
M4OOWiHUbHeoYXRQBNzGyaUILGqD4L+ntoWbMLexT0Nx7mRayYBhX2fbGGDSXcwQ
Hc+QOLtFAERdqgZgE8WUUvis2LfAz+36nL5KiyJWxkQukJMlc49W8rBP7Izoq2Tv
3suTRPThxEoNJQ5naNG+BTN3qUhv98BHhs9+cPavuvLmZZAtq2bxAa01meozjHq+
w4KkMxp5H6+l+tOGbfGt1FP1DCg4Te+dLX0Dh73kH4KkV4w/6kch6Rn8KxVip8TN
MK++qI2j/qM29gQQqsHqWVcAvYH9ZMBeRbl3I285WjFaUQLh7tRnTHiOLNz5eFlF
75aqy6fLUGEFQ3cprYAfnkObUD5E7jchrXLECVj7b0RmQO/qzGr8YgIVyaDHNZhW
9JpWVlFio9hoF+ZqAnAfGIWF5Oei2bHLSekF3Pe+1ItU3V0ILp/tKDqn1w1HGL9J
xW6LtDPem8Go4A40yYFBkVIG4YM8jisZjmK8Osa5BHg8rytrLI2eqoPdxZzjosmF
mNdvehNO3MHYrXdX7MWRxWwfcdrR8vtgsxnukYmI9s3OQIcvm2ZpPXt6v/XeL2vM
K5g0bD7FwI3cDSgf5HWl4+eb1Wx2rSr0/0UDiooSGs7QTzSQxWqKunwEURQqVA4z
j8sur/UT8wVnC0jX7awxNltSyOROvJX8M+LVbyJsVmeK405TFbRHCTgPjXbq4u7Q
8dtMHYSc4HJR/wqyhJC4W1njYfC8HHkicWtGpZAzYXYTIQkG4y7sjleotI2ppvbE
HonafDVomcWrmXWNs2xWi8p2HCDs8zunqp6Oqjch5HATYhFMqHfA+vZq1NdVnJqf
qdWpjHtm9NxRJGjj/uUVwzvPv/nekjdxO1PKGGcCC58hvFChEoklC3z8SbdnwYWs
binAgBrGBpRnu01tZqPzq2WPOm1KIe9/JGeE7GEhn63R5jAh91z6lVHIgpMqCkPw
T+SoJSqu7Fs4KV7boFJCR/MbxtFOaw09uRBYduaR16QffwfHSfRY60oXjUZyLkJQ
GaEKJQMBM4XZTE1z+pD/TQz5oz1WZeyIte7iI5UPs8JU2O9CTRkJXPlTqoFdeiTi
haMqwqHZ+J610ep6P1h1XuIkuPXE5dQB1I8j26g/B+x1n6AjkrHTe1UZ78bsQt3D
CgcnqDNitU6Ry26f9MVj2q6uHBKdu2M1QRQ6uEroT3axU/dri7ePMMp8bK4S8SCI
Kox7gyDDWOrdJc/9dzSVQ+8Rd8XTlzcIeUbZ4Xabv0kRc7MGIhf+swSPnJrZwxT/
Xy8uW7eYR5Nzm/PwCLBHhiFICKyEn5hTNos38I7HBu3QUhuWjOBQqz455YTvbFtr
TaDInXdp1PlHjX6dd6t1MhY5mrufKQx62f+8nMPOOZ2bvtY2ixJABQ1K6t7bV1iU
OV1Tokn7Ou64YXcaD7+tyk9Gd3XknR8RxXeKSaZ8/RtIBl4iqaC9cGevok74keNz
AI+F0nUcn/2XeXzO0rKEJw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ZxwPv7V3lVxHh6MP0ObwZbHMSsCalOfR628oSOuwOOpXNuXD6QY3xjlaO74zntJ4
ls8lVFUKvpmpEwvCqqU7PtpguxYJUV4aht4Oas4u2Po8iRgeZz/NIA1NzTYZmWyz
X+n4gxmE5Ri3qMzwbk/ipFwLobHJXgBxjXnsv89yIDRea80xArG3ADdHTyxOKipV
neEAkSl2OWtBrFHZgQJp4VE6x5CGHZmC5m8kvFOHusaGGJgSetBpLfl2eb2SQr6Q
M59a7xktAwHFZG9ggZ8d0/eA/mLanNppzwZUAzCTn9MwJ2V7ZtStdUVii/ViLH8e
jh15S0bGuDtSkxGz5Z56fQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5632 )
`pragma protect data_block
qVtfGWmXs8WWPLJdjtbUWe57GT3fV8JIAX/1xhfktr5/ZfpMZ+2WSOZ6HcLPKUQ+
sxSZQUIqwX1eNaxaRMYl41OTrg4AU/mM/PYL+S6P+Z+h4bQIRBGi+hf2Kt0/zAi1
NKcnSH9wwHIFh4kiGTLHlE2v5ZEvZMJ8qZ2z+bj/71Ov2+D1nsSd0gJ/NpavTWca
jRXO7lWy4WXHrqdIvnFYGBrfeWdPPVDUtriywN23D6ewfRS2hOcWWspNC0jiUKdb
Eobwz4vYOA4iyawenGJOqLk9rwreL+Gv+xag/npYNeqc8ltUKEA7l2aqdAz76iN6
bVyiCr+YAjlUJ6YvrkGpKYV9c7AEp5eYIyA+fm7nqoWyLHlEOBwwkby26mZ5Vmhb
vkF9FDBOfFmwRPv7TSGsaR1IPWIfG7+YjXWWMTiYA7dpv8MdTj4y/V0PFvdoHLe5
wW8KFAvO+0w4Bw0SONcI4ce9UacZcP8bpKsd03EPwPguOnQ9CK4b5xGjHiM7dXqN
7umNSCDK3Zbks3QmT3YulRJlCWQEwy0hgKK2KFxKVD0kmhN13ZgGJhA2sne+2la9
CtjpbMnTyM58+wdFpYufQxan67xyoHZsbbI8KyPjC0Hs6/ad8Y2uMO8B4FDzg3bP
88R+JswJpKWfIwbDdIXrZsxoSfeJ82UVH4qZG5lv5ZW3x95cMCG9+dmKSebs81Qy
p+gf+RrWw7o3lj5GUKdskaVSxrUib90MJNX9pUHLlH0mkW9sJO4CObhPYNlo0d7E
N3zNJeqI0bFrosCpNDGYJX/+DolJ7YmnJ5MElqIJ16TyVvoMcz8EqaptEfKa6ylt
0U+YfFVuzJx0VEaX7j8YQozgkwK9523wq8EK5iRf2yq9EDzBpMl+p6M8NaNGalNJ
4ra0yIjFvQm6KaVc7Lnq449pb9bI7fRWBt/0Migug8URmdktOZZ1Q2ZBA8OBnqzV
+iOJtHG1mWfvlavcHM68pR7+3pGRL8fKnK7knio5CyQerJyoEr7L6Q2U6lBH6TG2
dhgTLoWwg2er0/lAK1HIgcS+QCyllfX10ZJNAR0WOP1UX6Q36oaeFE/iGBtdCayQ
G1D5koPjrpUhcPV6m8iS8CuffBqCICsKdJbSHJEKt0jbIWmQPqsrZFoLztawfchJ
qCuYaqV4F85IW3HOkYyWEk38HdJ284Mur6bXmChklv/Z8K68kdld7dXBN5IsDcmp
9HuaidvMjh69VJGC2DLDUYbuz4dj+bKurSGOQoAIfXiJEGdrKahRI3l2h/Loz4kO
gF66yOMjUxSxlh2LnSx1o0Gjltv4eyar56tDsdcBxM2P0EmoQ0nL+pjW06QuLLMX
MOWkguzjsQg3G3PFk0Hbjyj6IO660EhqEA645s6uvUeE1JeP6iH/mKI64p5uQ2Op
cyus7fZfIgHILQ2sVB64ISccn0yJOtBlY2cxKZXN8Q5TanSHrMpGtt2YgCql8lke
5y7TnG3NHppxTXJvr1v10UMzMH5xCcsxWoU9+566o98uiNaSXHPIFKfcDFtIxF4W
2dgwoDAHVthiOOKi3EddPLjPh7aSrfMTR8mJqkIXWR67WK6bn+gsbO0xCPgy/S81
v80ly/G0ucr+mFKq8/qeB0HdlMhbaX8+lpxVFME28YftkPO/IRJ+D9310YAJUeUn
P74a6drUDGP0nfJGkBe3XNi0gzKoYSl4FgMz7XkGlJZznvj+hmZvRZ55fRqnZOH0
HLqegDJI7qCNVkzqu+FVGzg/TkenIXF8yxNeo8d9UKbhD7kDWBZl69Oalneg5Nut
qztfAmtQLVWa03uVzGaBjFSfbV+ld9cVF7ZDa7LsgNTye3jR5K1ZxPTO19I3m42O
4IcsTmXVXbBpAYKzEIFusSzgTXjUQF+tpL/ssaRjtCFF6bVaPO0r0CNnDocvCT4I
WnVvb+DL2QKQ9d3Hddd68Lp1noQloDgZ03Nm/kwBuXotnqTECQBHxz3jXUlTmeSe
NzDd2gICwcOM+WbhD34xiz49JbpC8obAeKIIDf/1nR1p63C4Hacab3rzCUJuK3WV
4s4OBbqCq8SGk11lRYesDOcAzF2vA7cfzqUEZHu8f89KxKvyU7yoWy09vTOp5N+h
q//aTJz34F/p9KTfnlBhDlguGqOaT9natH7tP/37LQ5Y6J+0I5df+lJOPAo4GmrM
msXfB/YQMPh0dmjCtA4us3gZtPE5356LQojrdI4oUmPH6xJoMyttTIBhK8DioXU8
3i9RUqXDd7znNeXa8KOTIqEVSTY6lTD/9X4ufgicBbf3N20Z4swfEE1VCKEK/Abn
dImgQhtbKx40jLfSUXKUNEGw9pWk/VO5QpwxAnyhtrjrd4IUYrOqnq5vuYgKNqBf
I5kDrKtieQwsjYOmK+0TyFMQjIhA2n1hWlp8ZRDZzMGJN8wJit06TsVc+LyglD7+
0YTaGVwMgL3ogPMg2B7duMg9trnXVbHZtvLEtWeC5SNt77+3jhgnUd80tseN3S/y
WpAAfZxSaM2HthGIEKimnpt4RXcCADnSqDrmCN62JRerTpve8hdKOyjJGwMEhQZy
VgmxKi9TcKRtb+uHgHjv+F6COCHuVInBBIORbT7vuQwoY40aUmVQfBczolXi2Hc1
pQWCG8x6qDSpllAeDZyUx/FVVP2LSULG8YzwWI7DX9qirXzCjrzCdsgGfYzm0xEo
OyENcPZjVNSQGOlvZY25RV+blPS4AInj+fZjYP/ZEg6hLhb7iPnoqJQbXAf5XDhq
re8Z6KGLLhsXsYzuX9DvCGYvR0D6HoJig1FSjsDp8J6PG3dYPpR9OWpou/CpPLc+
H5oOphSX5jrVYxXXjhFwv9h5Q+bKahw5pEp2AMBfwkW7eZQi03lPputEsOuNn4Y0
h+WIHjPy/2CdiLg075wsFcfKa3pKYi1r3KlkRTwc2lXLe/SArSPi7oSm6ZIvmXGh
nnw1RKqvQ2uJtpNExV2d/53fSgWUPuEC22qL2IkFq4x/HvuiTRT6VF9/btQDA0Wg
7rGRMJbfyOsTvO3RXe4mTUJg3zPKbG+qIWBXMrd+tJ9s7kRb1x8DpRtd4LSgM40L
06B+kuSr6UYdL1ctkFi0dNcr4ZbCCmXbjH4dzYXSO7TGKo54d1Pi9yDd905h+941
9A6q+VUng4RWpyNYfpLJBJuKCvxBsyVA/NYVxNsdJ2x38TPdBnbj1X1OvMS8eUrS
TvWOfwwjRlWPgh1Vl9g7L+raG9kh4ImhRxmSHUpC60EqFOuFjyo8fQ0z8lEAfIay
M5vZQD00L6Pcajx+FQQzhSdlolkQHaijZPLmkOwAg9Af9KBiIQgBZ/0QMmSieLvZ
3b9/cOFtjMkcd6v0oJ3wENpbY+ypgOJSDOING5DOzKcfJCcHyw6FBDwD2e+9P5qS
CwAebZx23qX4w1PxSBLFR9SqvAfFg0xyCUxoiD09F/vphs53qW2/NtfDJm9KM53X
uTcGyboC5fuEh7TJiIjylMY0goDItIjdFn4hwoEIdZL7fe6dFhxadzBeI7h1P6Lf
LrAS79/nHwO45ZZak+9rqXcTOntpjEHloY4dcvssWMrRUvd5Xw3weOfao0UanFN/
9+JMvO/tp0fm7uzyUa8KCHenUGmPEiVDnPgw5/ECiwYxpmXrpE2fv3dpPrhIvB94
ef9hHYVCLQd3mJXhRjpTmk6uyrXeCUn+a6oUGdjwu9i/cX486QShWeZ+sWqk1OrW
5EynEQNPHFQJ3zolwjSseLFP6IQtCL0HuY/d0pAU7lw9BNK7SQJycQYMGOrFPB1t
2QvPIM7NI9I2KBjwYrAvIciTLq/rF35Ieq4SEbfhDj8O1V0EQDbx4ChjfU3EKoGN
gJaDdBt8ldU4O4kw4BNMDl2sDKtpIxGdKc/Zyf1qNhh96jFbPFgKwsBKjmlz19x5
nhhIvAfY4VQbogEJG9EGwzlkrJGfe1BcoKGVIl/L6OV2DNkfMMtG4CyVAUNdeNhE
gKiy+sYm49pdFeYCONFUlqrnarWszAPUWOhmSphW0zIGPv39oEQDqKVdOA2SQHDX
OKxGXfqrwyZVZAlQZ/+ZVpguswHFPVO/paVbDcImjmU/+S3bAhsi0zON0Ou9kJoS
wvjLZCeiysLQK4hBQmYk4kSAG2PscVOB9robBWK88QCriTaI5gC95/AnDljKipBT
DFJzDmeXO9D4SLNwxf2lBMXOinWw/uZmPlxMeOGjMEOolP7QmvEtzR1gBOS/KVEO
TDMOmDD+Um/BRgnQP8pmtl6qn51ZXTuwpAkJ02T02mjskpNlPcmfk4LXnx9S4zTy
7e6mD4lD7kBoYFCSCgzHB360jou3uJ+d8NfzmltjQVyBpVe1gbQZ1M9SoCPIc+no
kGhUL1sKUbDIYAqq3Rt0YQPQOEk9rhBcklPQBnPKoBkMy9hN6ZWdW+G4TRmhCTgc
VOrt4VH0YYoNjx5hwQFv1m9HsSvsHoEDrrhDNvtvlVAnbF9EZjIqmdL6EdtOQpD2
qsLbJL4GqE7bQQyMjl/pVaCT3v9KB/q1/PvWghyEiCYxhLcTH+Raj/jDeQ8VF0M4
KoPry1GWowEVSXHvkUn+I17s85JRcnvnSIpy+Wyb+nvGQvbGJWuHOEOU1B851FFj
RuhkUZBtkp1STfdozOKjCwU8f8/VwyzuZehkX1gY5I95MGg75xpYEzPR70x+/ZWQ
eGWLV0h8Mne7jgPJXM4keTxf+mSGB99rMk6B3fVlT7Qtg2zz/TLNvszCZsvtBNcw
5ocgX9QxzPWl622/tR1/rIRFv+0isUh9jxw3qsrazL3VYRWyPPGsLRIPSlFrc+Nc
8zB/1xUbv+HVWp+tdo9VxWJIJ5BMQNxqsjOT1mOYET21GvD+0UeVusWQd+WgatK/
OzJ//TYbE5G4X0fPWmhIWKXQ/nuf1Ts53qHqf1u+DyhhbwPD2aC/yLzqd3qpxfGp
tyGFWH8W7g+VMSw8GSlDjg6+KPO/EkGZIgDhFHABK7b0m+gBjib3/mJm4pvhe8dT
xQDBCSFPY4IGbOlkKH2JdRTlhVvrN7Sd1dJAqtquuL+T66jq5RZgyW0BveUdVCF6
KqGc3P69vqKo1lzzLrgxLSb9PYfxe8m277LytpZxLzWoM1xjP5Sm/DX1GaVq8OgN
kcOnuM3L6O8MwsgNv680Rs7CQHb83zDwS9mcdnEqyoYIpzVmLV5dIY8cdIkTUixb
MaYgvpJ1PIcUTymOSTaNTjBYWgOwJ6OG70mhJIxQMiIVel5JBZqJVe6JxoOBeCYG
vGUOGeweMNjQ9GO8PQuUuJn5mYgvRHLFSSqNqeggq09pp98SzlIa2RZ7dBlCU9hL
vuIH1dkamU4iFCVRIoQiCpUDMflLmeyNvQuaJ7esxktBMnBfWmKF7FFRg4s8CySD
FSSYl/ydaKzYdTAleJzfZs2gQg/coIvwyaRzRPYk05+r38MOcGYQNEHoXbTtv81Q
6AOqDcWIiuL5UkZIpAfuan/ysSOF47h6YICFHpL3dhNQn7Q9yEuITn3uwsYuMqOF
h+11joqWAfIW04JmmrPjucgZzKxpPruD+ixcowlB7v24a0zEMqgbwqQRZBlM4/2M
8l/PdcO77wmuhUpTnQrGlhpVY2lSjFQlkN8r0Vk+tQaCptFH/JiEfCYEeM7IsAjn
ljCRAOFXe5UoraDtTFRcqxqe+Ag51ReH7WW8XCSnbkm7j44/TlwJgYKTcujpEoIb
vfA54K6wOTyRMwdHrCjtz1C8J1X500Q3HPLosWLVJMlLsHQc1Cd1hnKG1QQCxs2W
uolw1SKGVBlSd8BXz1b6KbwZYBTyxnxXuxW+oN1jweB7qssJdTx2+8b5jLSxIZ6y
6TkdA8vUwDimB8c+rDW1QqITXeWUI8aLN5GV1WxiU3y6970p59ZJYXnxfiTaKpgo
tdEN4CUx964yZk8OeVbZCq5U/RzoZQ2pMiCTp/yUuR+Hi6HBf6c8gX0RoBHLh0A1
YKBnJp2g4F+ffF7RJd3d9tVCXPkliVwdZ0eFWbK+NSeJMudMhMBjphmXZsNU28B1
vxEwDClAzdUqmWHoCTwsSZ1IE6GgGlZLucU0OuPcOO1kgTcrq+Hx+tUmRnpRPEhi
v/fGmmJAiJVyvICaEFYP9aJuXhowq4I+JDC+Uw2tXSBDbmlsPra5dJe9R6+5B/ta
RuEj/zilJ/0pNl/Ly/wmVGq1b9gu52oTdtA01X+D3cc9M495poUzB0j4NBx4zbYn
izy2aLr+OqdSYYmLIDQSKnyIxPX/f2wfvX4buOPmC5EpIHibziMBxoUX1Uhiq3v8
k2tUbjU4ctqt+H5USU6+3sPtBn/tgAjV5+dSdMWQWiL/LjKruNrBKJSYV+Vsil8i
ZSoAStR0ccLq9UoJyZgonJAZ6sHR4JiVZbZpwWe34FmPWGxj2aIFeaYDimEepDb3
LaArQzJdECR8wLwMnR6QIhj+7HvrWkPOKW4BUEfmekan5/RQMGkEdJHECSxhozk8
mE27zI3ODFd45HtvIHKE7eeXYbiXzZ0nf+5z8kFe5Umq9dcprgJ17LZkOtXVslqg
+qbeiiMY+P5LpTCudxgnV62/xt9On/UOSDbGYXSP/0oXkrd8dyTiXPUa54di/mIQ
a5jo5SmijRkRuwLwNb4u0qzHI3ToD4n2tZC4vO8WNOLY6xXX0HIYjlTob7eL9lEQ
aR3lNqE4mlGAJU9AjzlIqckQWCpX4R/oJxBfUmCSfAaMl5bTCugG2k8DB3W6sDG4
ozcAadCCvmr/OINUZx/h1walVORqptizrZUIJ6AYl2C0BfJh7I2ROTGSxHpFg/lY
wnDEHMTUnv2SeGi6aqryFxFxZut/yJ5zBhvsxPnzQ7Yxy5kO4E2Y97BC/ODYcf6r
loVQcvnz0cHaGJrFo+c6ap4qHXQ24YkppSyMTVY4ZzYONHvXSRt5K7xttVOHkc5R
YD+lvFz0RFf9+myLmEm8PECu/k9ONTixeOKO7gxwPexbjTwZF5bSM/TBj2CNZA0Y
szL+4CJcAcxiX2CLl6fXhrSWVIc8g0TX+obBFd1XyGOAZ00rTYAV29d5UVUGmIIX
BbuicIwlnR0Y+jOhrFQWBRfj/vurmh5OyYDQlf76DxTBOZ4a9w1ZOMwJLzD2slmn
fILzz8qfijjMCmd8CRhJU/VsfK5g5VsG7r4Hkdk2QcLMlEhT80P76orQVAN4zR/3
bSS/2akEf0Dt8fzkTg1wH6n/K1dwhC9VgwMguxAY6+nE4tqNbeD6Fymdu7XPVxNX
q0q97/GT+A0AxBfHEFFRfHYTgDlutVc5KAp8DmSatroipyEQ8W+VIBIMw5/JoRkh
e9XDLxQiZ6x4g77iG+4DdEFBVRYeZ7z7sKTij0GqOjaXvejeGu+SGrTVi5BZOSoy
FvvIRDdcSm7BQKWdMen9NrK3E8UPXUlxdsiz1tfTfMCAYQE0t2OrbFPK2svA4Vof
YfPQu7THufLdgUUETvi4QVkh5wgbmv6FDZvvcsENuzZ/1w1TD4wsWCdfW6c3MFlH
M44bb41CVD1z/iiL3NCt4A==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
I43O5yDkIcGdN531Y+BymihBHqK89Df+UnVI6vgTdFo3sBag5UhePCkVQoTuruTa
BnypuROw7/aFg6Yuidnf59/AUdP9YeaLjy2aWtlHNzOUaQQbxix0SGtFehJ/vUV8
bh7Z//wpNzdSn/Ft/F2zEmHjKa7TlM1kGuaDONOaKMkgflZs5leKUeTnfEDF8bQ4
4fuj4VSnMDn1witRebt4t6BJYf3GGvqAw4xZ1KSmLEWFvIbhsuT2HbFLre32ZByu
bOoCX7aq8b86zFMCOq0mA6ZkSPOMI0KHBHjwkfbQ5O8I2tJOwjKpq8gTxZuDQubu
Cr2hcYnh44oVghWHJ/pNQw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4928 )
`pragma protect data_block
ViF1dqPd3VOv+AghQzk2nAcKieWAKkLud+omFgwT35rnt3io1uCBUGkoid7HFSX8
tPv8Sfpn22yxv2bhusOHMS8zl2ZMc4KNgr4Rs2ThJpMiUL0lk1SSewclsg962jFc
eXqpFYszq6GxE3Uu/tVmQWn7MkohTJurWhek1gFKyf7pebKfThGIGlmV7JQ5Amqo
PmSb2TAO5YMNk5o26udyj/ro04jgvAlbuVfV1XWoqzNpgzuOpqC8K7efubqqkREQ
LKDfQi00G0rZ261tN9kBC3OY6xpRi8upearsthJmy+vUyZ0JiafFyuuodETxObqq
jvsbKw753F/kPg0HEg/BtkEOhaCH5fEhaylQczULRYw6RLm989artLBX55GoBsjw
vlG8vCojfY2TU9dGdBp0Nn71GK9B7tePpeoCyjZmcJUpALKvYJbp8wfzn4XMi77j
3RayvXWvtvYdcWYNwSgyDJak2CtPhwf1lH+FPOydpAnDZGjP6wRO3v1TuwzTJ3uR
l1uFl3NQLU6tH8dfXdlviUJgWUijbePqSHxYvQMoBYQBXjfvDyxdyIucNWUg5Liv
DZCKuXsRVIgdeNMvYzWVW/25OMJ9y7Q6CZGRZWSCjg/17c3EUFXCXziqWj6U7VQ5
Ql7BY06QykKwYkx8ibO4dM3+vkqd3y40XIHMgLb82LDTbDfoIEhuGt25O5qU1vad
2qIJ7OLXwZZ26Cz3hQbc2COxdYRiwX8rFGcMReukjWaQsvI3rvKvtw102L6DGRZc
6A8TRULzOkGvxQOLgnDaOahTztk2lqlVDdsiuz7E+WTDZFoWEKeo16X8Scv7/Y19
JMiz0spg6U7rMlRB+R0cTwM79kIt6StiyKlcGwrqDGik/q19qzBLd5q0xduDEQIf
JlZxjNnLu3jI+QX7xN6v8HO7RFMaUHH7Tkehdnju/U6+z7zgpN6s92zJMyxlXRN7
/ugGJaHN/CMa8p24gHeayrWCWTa0byTiUW+aQk0qHTO+RP35sGGifpps7tasUyNz
9V338xX4u06yofewZh0dstdbhhJh4EH1wa0L/VW93lLJu+ycx9CeXlsoIi0Y8kEP
SaZeXpnybg+KLs2wvbOzjMVPDju3SYducuDe6WMANUFQtpNnq4NhVVJiKxjYvYXI
rx6z6GkGMlRnpk7SIOUYWt+BMHUXm0Ri2Onpi48S/CBr4FvTt5U2t2p35WpJWBoI
Cn682l04JY0xWRpJ5NtAwaTwEfJB+meSaRQwXFdpjGzKWlw/Tj1zorRKxQ/0pS/f
5mQbcKUkSLZ4WJOqvVKzQnSXzYEuf+Mq7ady6ZYDwqt6LNxh6ObfdPUIenHz70aG
+hbysZIgLw/I4Jap+lfzRsZaIfOwZ5Of2aGbocFGmY0gZ68faB3Rh7AcqZJmyQ3v
YwVPUD0cnq0m+ynvHS91noghQWHcRMk8iuDPBXf1N5Swp1ZmEUlK/JZ9Gt2ogR6T
nMslbso+7N0eQImLRhopjMXzHW0oI7J+zwqS7g0rf6qkOchD0S1p7QOpmwhllkVE
JaALADcb3L/fmLnq0UPe23gOxUk5QZjx+5xUN5nFHudxH59Tl7jvW7c/X4kCzqJL
eh5S/+upfNx7JCA03s+Y1zLIUHVHqCzr/H/6KJqZPUiBsbsgMFcW9E0ims8oQw1Q
CoJUKGK0noie00Yt+E//6SicVSE09XWqG9ywlWqZhFTRchK2ZaKjoN7ky6R/e1m0
MqrujWcBt+ecWDwuh+WBp8G/1oky7Gzf2TiJZ8t2DCfSLyV+MMPGPNN5D26yQxE7
G6nOOz/LaPgnG0ulB9NDOSF3hs1mTR7MojvSnWFiRRl1d92o+evYzp7Hxp0HiEUp
irxVxBNDf/SQTcKPHbJhb1k4PXzYCC5IkM5XDac7JvGWOqJ7kepngboZTTfs9w9G
STwLmraSAnLKeG06ZiRnYTs+tCKC0pYhyJ4ma7OuWwjGMoDw+bs7s1Yk2mxCzxKd
zjjRGNCB1Kib/kfUYPILNiMOM7KToLNgOw3M2FiRqCx1gWiT90uV6IQMPht1Gs5k
GuUGiw+xvCbY6ZE3JXkEARfs6Dp7Bd1vBhQfCf2KBIKb0WJnnq+b248pIUCKyHvE
H5UT8tZ7/uVhWBsVyauEygcFFBSb8c8Xmm9wcDZN/zqWSRJ/JwLYYmH3PAioNnbs
qYMk/X4lAYx0YvKAGobcnNeKgiotVBjrPP2TTtjMM9xcYqkXSBJWFh47kpi2IH4b
5rBa1TLCJaGeBhFQpmhHNAJ66m3ql07hHSblgaX2dc6uDappmuc1p3m2OUb4PdMN
y7cJ9nwV/S58zvPRLShx4n8dOpbw4fEAMJoKDFBxaSkqzej5ILKmgMI7A83lACKu
VSU6CRkzAoriNhCsM875XMA/H0FjYPjsGOcMfH+UgGTlV3NqFMX5vOnp3FqV6vbM
3BWLDqjZE82ypdXiJMCPCYMnClRQEkgk+JQYFSSZZV6cHmdZ3TXE4S2ST+ijNsBX
MKoHC5DZKKvQIDUhmewb8Yr9BRe5D71RBbzlWBLMUW/Y9MgV6bI0y5KHCFGHXYTU
oRhyAzfIb5QT+wliArjmp/zzPOkkUWyGZYRVz1cdjr6xPhg/ao72WPDqKgP8z0hN
UjN5wETDu5zdVv2qYHaEBCLDtMmLU9HJtHheQFVhW6P+deh/Ss8tCFzpnlZDRbOu
JC96iDtXXMJdNWbpQGz/qBm3A4/kOBvzOeCk7GXdEHBPkzrLe1WBF9iYX1iM13td
aCL7kwutXR/pTvU9fGqlrj/f6Rv60eHtAWlb4BEEpsIBlwDL2WERUvVhR+rN00VX
W+TTTpgBW9k7Gb9FcQPG9ZjyIQFdRWxg8t1Mx8yCyFc1EAV6XebAj4O5/ttdIQVh
XkUvhQD5vSOSaPxVes6GJdD/s70U4feOz5kabTSXu/v7IS9oV8VCFbVkjpK3rOqG
vH0+rQoiGbw45nVZ9g9bRbDP0nj7ZQXMp2rHqB+lFKWF4+CmJZGxl64+Jsy5Gkqo
tY0epSPzmycBatpVklCSx1uUu4raEKVwXzL8WJMBcmoy90zZp15JhW0oPyv0Ejyx
YP5CI5NGiO36hNRwjLMaPeLVAX5UnX0axmgn8Wv/bdqEBjIDZXbnKraipLCIaDg/
0CpHMM1DaC7fahcm9ZgHTqQaLma3QB0u5Z10yCfg6y6VIlwoxtCfDVoJrOgAynkB
5uJWb0uGl9SqiOUqdbFhDF5ROnh4PJXTJEffRgecuQJbJhxrTT380VcxBYgjxzXt
0fGNM+7w+bm22s5Puf4UA4pHQZEadVYHo9Z3iSdJ88cWjTVlXIkcJAmQ2nakN3Xo
JpLyaqwxltFnmLP46LmR+NSZblX6u98XVM5HJY0OzMWCypoU41zszgKWai3aeemn
fbEtJU9P3TAyiw53qqJG7j0wvuNNRYsQbd4P8aIeHrb0PWiDm4iAzkrb95BGPSUD
AUwKUNr/mBWwf4xKvGESCrDXOl+aFc0qtU/dF5Yi1A2NUUEo304x8fdP8tZxwALc
HMMHA0/iXlYnFKWZCaJyLoFZB/S67a7owNLaemtT5YIvePWYM48+ZJO2xN95MCib
buh8VuW1uh4McPBszDmoOCSFr7h4jUFUWE7EDhyWdM163IM32aO4VFPRFeIuqN0y
9O1E/XKnt4yaHBnxmGPUHXei6/Fc/JDOZLr9P2ZIszGKiFG0ZMgUSi6b8PyGAn1h
QEKAmvCpykFGnfnIE9tVNff43pcP6N3vLjlGmvdlFASkL4DbD9vKcyQgPUPCA6D3
nPoQWtsw9KGw6kiGrurO2BSmJLy1kREwlUDpxBFN91N1gggjBXtzIywYXr0n2M0A
wNl57ykwNrQi1I7Tcm3QoJ/n6/TsXAmYjIg/wrS2fI3XUnW8wpwnrHOGJ0mCG9Mc
zREap3sznp+wPLGfro8zwpCQJxkNg+BdBcJxPrLt1K06gU503g23axi9aPobB8GY
cmECV27Ndm4vf8vcDzZ+RKy2TJeccI4hMnFuF41rV1B4uODF1AQIk4oC5DTt73vG
T5Vlr/yKnE/o9ZOzlyBPLygmXD/Rx1nGFxuX8N6vU5Ougn+Hfl6UnOiwsukOSD02
lKGByYQ6M0cqiuW1/7wM6kNZkcZUScwrx4BMiR98m//ZSUMPwW+clgHX11bRLRKX
+g5nSfbMLgt3AvVDVISd10DOofUo3IGsVKDr0VEzLUBCDBzR0W7DL/JyxI+TPG9a
05CHMY4fRgXRmbmsg8IofX50truCgUTN2/kWVsivAo0eZ96A+v1K7JAi5itMDToZ
uAqzezQRuwjTvlFrVRnBeEZaLegW2GTbh9Gs5BV8Dif/gd7qtq+zaYenyr26ThSS
f/QuuZDyi8jgmOUlbiANRwYA11VUeqP6BM/vMsfZhS900wPmu1/xXb0lQ+qwg9U0
uIRaGbp0ahk9VjFQ5aLuSaUGcqLlJur/GsYPTZknHWWNfyzbWLeelo6URTTwUB+S
jVatKOjYf/+3jCjwqep/Zt9IdrHwpIlWf1cWNCJcVYJN0gcdXmP4VyHFJqSJWa/r
VgTsBNYFTrBb0TAPSD8/V/mswip30ez2W3J14+nJ5sxDfaxOkBSdG+6M3WDhpLko
K8VjdFyfSO/++e8HZ56MBGeshPXTVV50nxWEaUkV3lFnNoVbEj0ePVNxjUCJY5S0
BEkztPlK7/dA/e5T1nMXOL+8APR3Kh95+UaHhcDyjikx/fossAyi28tFNm7y61zs
ilndO8GC4hRo17ahsdJ6v0MszJgEdLzQZO2+qrapzNa+cmEDQB1/DsduAl6HKBhP
HUE7nymEDFceBCZTRdw8z1t54bBLtsSMnICNyOmjqwtfGlEjpv0vz6ycbcwKEtmK
QuMggT07sckpsrRwF51j8IeKHKqktNl+KMpzyUf0ulukSFe0R/HGdF+oQRHVaPwQ
evCSSDRrcDgMcArXmRgy8ax1+yBeNHy1ORcQGVf0Y0d2d/O3YCufMLZfeZh43ELr
GafKJp/38+hjDGwaReW+AiWRrWjJVBeUi+lVL30LJtzSyAyuOIrt/pcvHRbxXJ/W
aTp6DnasRR+qBc69AW8SslHauZu15Qg4rC/Kkf24sU4BPH9VnoIwDGCXviVtKQKR
Elb9I+yLqYQ/8orN+IhCqjRkkk8mkFCCyP1R1tAO3mMoeBQzQWvP2WZxdKrbLDhn
IETNG67AgMy3r92jQtZ/gTu/7lwXkxob6sNb2V6ujYpR1akI4aP2G0MD7Elr/OIy
a1Z+JhbDhYESgo6W/px8WY0D8lMzeACTPon+VCqHOjgZIRXeZE4AERBO2C6Odtfu
PHGwiucq7OvvFqLYpXXCv4PavEFayTOCPUXqwDhoqyG1L80veqho77AKH1au+JJd
vYE2inrzB8kwMUVYTF9NaM1I+UF1ABOvwi1FYfRzIzKDSkGMqn+gNHI2Oiie0vJs
Wlqt0OmH6u3ThJKa0UEGB9TNAiFkSRDkVH1gfcIh1lS7OpbUqnS5d4WNMV/26J9g
E7Em8wuMnVpYCslRYGytaXDjZ0lMVxPc1Ho2MXdABs3HuLyFbIoC9IdimeeRhD11
pI5kdDL6QUcCSTScCE2a0uxznmiojjO7gurJBgCfJdXShUmTS03VUxI4X6Kd1n9F
3qxbAPwGLxHhXJn7W3+qeiUDzLbWEi/O9iJZ2ZOvJxfltC2AR7iXlV+OMDLUV2W3
DNQcWGkBm/D7AYSYW7D287mLq0CDYlYYQr3wZpOik40rO43D3eR8gQK0OJ4y0lMf
fjxsPNLhHHsYVE0yIcf/qkUiSKNIJtPpu2z9WD/+syj7h4nXRfasajCrZDoztwTO
pn8KIcCf7WtokCyheHE+5lXaPvy6Ak0UPhg4lTftRl6T3Lc3tKkWoDUfIQHPAzhk
0ND18oMqyT7TLvYhtmvADbwJzz/UZhqO9suCG3Qss+1a+jmeIkMcjfR1aULzt68g
sTnuHFt684aD1IPRq+ecg5n90XNT6bKrPaIm9K+BQyMPeQyxIRw87RKBpa6kddWK
/7FNGtjKSIWYoS82wreqFwZDNWXLYvAko/CaNjuJ2egAIp4gg3H86Q68yeooOjxt
xc8jkwgQ1CnfkgYFfm5xZ0DvNuWQ16UErwGhfDaCKftsiAGR3xSUN17azd8zP1XI
yN+trX4T31mtP4Xzey+ZoGgoZVhCmVNFRUCtGWE4e7Xk/WRQmgml3IpAiRAyXM8c
4wevtluVQ+UCGE9AOFIlv4zhHJzbpQWQGBF4+uW5JsrReZgQ7cycDOSpUzZ4FE6I
wVqkilpsc8Q6arejd5kdv4cTwxfBJFsVIW+SdV6OV6OVtEZjBRcXEiBAeFOSwGBu
yUyApeW6Heqj2+x8HMsaREXzHx55yBe8W5FZm5/USN5n4VMSN+6MpnDitkiQRX0r
GBuuWRmkR62SVtNgGu0p8vsmrQyT5qWZbFP/1Azb0FdDwRUt7AoUXWBvUOUznXzb
KlOF8Vpjfm60S3DgUYgBi4ERfNTeqpuUh1bR3vaHsvJvxorX7GG2fz5pxarWVI/o
AYq0yVABzuwTqIJGVKZQJvznn1eYIRL1Nvw4/XNAh1Y=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JCLxyvEKH7IFze8DRJ6YowMw18CZt4Gn6sM7Xi0xA+8jXkVRQkMEJHfd5H4v+3LF
F4qHlWhxUUyXu6iSyQb6TmD3aOiokCPSnblM5D+mBEBddgXMGezS0584QombVggT
rVbxsokD1K6Z5nZej7UgfcgWfW074OX9fvtY97c4iRJMXKwdZgIwPUHLSqxAALYE
lFYVhheCTDqQtZDbO2VQSVuxKifMkQyePjg32wYargig/IJLgNuHEmvdEbXQMVt8
GxF/+p2vqOTZACz9pTnmCn9171CALvV2iiBKZIVXp+OG4c0cKV4KuCIMNAXDvB9r
ZOLUXP8BD5ZVZVI+3iOibA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9792 )
`pragma protect data_block
hGWhC07M4rBVc0yHogD7vNnMC8gE2fWmxiwI4tswTe/xnK7qK/qQ11991S29IYbf
KDXEEWg//w/DoOdSZ98/NsgZsSnjfSSa3J9V2EA+O5Q89yOa8qhIfCpELUI7saxn
91iCnc/cQdeOA6Ea4MKdIj1zHAY5WyHhaKam8mM6TF+88AMNbjLBF2xTM3R6jP4Q
gmHCwdrzEccGUZF1926TuiTdNvgrmgLcbXOn7AVTsEwxcn2VUnvvT2oXv710GDUK
jDg4UrtTcqOKZaPE8FkcbVsYDxks8Y/1MHn/FyrnxRI20jlfsZHAqWCehleMBmth
+hiQxKFBdmN9Q/QSdlNlASYixZbfpkW2IBaI9k+tlvs37S9FglIB34rPPx8CSQdw
7Rg8cU1wAnacQOlqde+81iIx+K+33erc81jRX4ntqtduLy2td2t0wEnW6tfG6UwM
z7qkIBs/auNU9d2/7t6PcMk42DOF0ff7dPnZnHL9F+RCIHF3TmpDhAcT006OG/oP
XkNWYP90xXEnY2MfAFVM86PCQ3gPNKOFErnfPY94kcKRM0SF4zzXTcuhFXUkS1Sc
a2cgkuhFSzADRaAMn56fJZQUPub590EHj33a5j+QyYpznVlisYJs51JMB0POTlpD
Fj+asPmuGkDJmEMEWY5uH/1QiTs9YofcyBBnj1Aze32xKQAnkoJ1uHo5h2AieZ71
Bv9EUtYqjtSXm6iab8QonWrCfCrNNXJcYTGn3L7+miGAS30D/k+4xVmpswJgoxUA
WmxS2+YnxMS2l1cGj5QQ/crN40WbqUBmjUUtlaUuqG+GGWjUNLmFkLAqUW0L/LuB
8Eqq4kUpifP9Yt1JMsxasp5GGeVByrTSvtYX/Lh8813M5n+43OQMNABcTSOPylgB
gYc1qJeZxwuZEFbncr66dFZxkWmlQbq3MBFxELa74XCgewNquWnoi9q/LQbxs3pa
jqWXp3jwlcGMwc9w5DV8NsGP4DlW3FUn2Rahm6taQlWAN+IFJYA/+eus0GmXolBS
HY9tbfFe6RVHBr40FPwjoDYCHoX5NQWAzhQ3brfSnAJotNuESeQNKM11753ARyqW
3qtJEYt6JIW0CWJ7tF85unYYWR/TsO5AhP8r5RlNAhe6LKY291nwmLzcmYNbDpQL
cQ+KTodVMzQbhltuJV4e/RBXFl7oweTG5q9ANFERrBQZXGmog+3ScFB3xD3nIQtO
ozcc2RvH2RJomF4rV5iE7dKhII5I73oeX1ai/4chNONpMU9RbuVfyHPKQGzeM6E5
odJCYcj4gZCSlq1ubZJxx4a7FjvadE3MQ7CFWEk9zb5SzFvWzUZ3WlzmqxrNyBLH
XYzuqOZe4FZ3s5+177EMUGzqAbi5o8bTsXuwAhRP9FSDxT6/FdQRa4XYJ2j1GwJ4
1lg4ZUv0Sgdo3aVAYbV/DLt+N3kdLHUVLH+VbM3hXNibeO2xnH+bUGcM4Oy8ixSF
eQt1cMW5rBq4HunctReo7nI2qheVCqC3n9XE4BHFh9S/be3OWZ1o/eJUu1dT8663
MXhWGHqMUbXmK2C9p1tGwAF8CxiMbzMGx50yKtYtGYTO/FMoYmL9AxfEGvdzI/cb
aHIquALhZtGkvGW11ag6Hto0rSPL95bMHa4WHExxXtsDTM5JmNWJ5C9U4pe1YZ6Z
5oJnlnKj6FNu5vpgT5Uhr8U1LowkWd7FunsP/socHDvATuZHGaZ0Qr3MDGB/kj4T
AOl70FY2+PYgA3ruKme+Rt+YmUcV1uimlb+1jtobDitGLoaVvXXWxroo4f40N2PR
/r0AUvrv1oWwofrKtBxgUSVLIcNEVaghJH/7mCMT7Sgo060olo5eUvUh/Rwl485C
3SjsraS4yhgUTA158YLmNgNJVLX5a6uSyW13osHqlRNIBTNuE8mcld20Eemt0eiG
1k7gVFCKuxStoT5rPFMtHcPAdPt6U87qQpNhPXUg7c3XI6kIYk1+hAU1pAdXXicV
1fPZExMG93B3cbld6jh+T559fj1nYgdtY1jm90MVpuKeKikUgf2etLHAMakuBUXg
rVMwzx5I/1zL/9O4gFFploZr6iuGe7TJF0CDRimv3d6ED29f4a22GBqo4ESbZPKe
6qAiLYogQ7zF78VnZCPDcbSe7m9BaoMnytApVRy6qK2MW/Rk+UgeavrNGkxq3zBA
d8oGHwM3D5+UT5M+csMCe3/vBHcP/9CmLxVZze74V92G6tMA5E8ConaDIvzVjwVW
f+w65JrL/sMLksAnP3WMjIj/mvqCNBzjlb79SWtBhTxmsgZ+CgYxFOIXXzyTi3nN
wxkxFl2y6Bx9o4btO/e+NTuGy+qqlosswyrO1eji/zvZr7+4NJzDSxCFxu8g8E9Z
bElfMShd9ajREKfSo1zkSEWL9w+LbQaje5qu8dS5BNyGtKS5cWP6dfK1VlxhFIws
TaCNVrPvFqnpKaq0ew9aZvSd0gXhyB6xnTdd3Fl3ht9RdFVIb8yoLCXdcCcImRpr
DhQf+eOKxZh0RskCWXBkojfOBsKEALCMV7V/8x5gvUDIuxaBZEsx7SNWQ2wdx/58
oqLXiVo4eZrgr/QZPm3V7mZSKFfV8FAJetFKFGbijJSLIpoZMGcCD7953P6cLfLU
SiVizGEnNG33yB18fhBlQ1waPqZV1W1veMiR8CnPuJKBs05v7/sFUhhfCJAWTmZX
IVHSc0aXV8crT8NOYqkHTXY/bd5RcP+qqyRmNnn+SI6QBRiSwJ5qaATSySlN/pOg
P5T+DUSrFP2sYkfrN/mmv0x2xNxWPv35NoYZAHxbUDmKimhPGyu3JjNQG3t+fU3+
osaBKOGSqCuZrh1z27S1vqvAWa5fW4pFGWpcjK7d+ucfoYX0kMyO0bzHfKgOaSlc
BpYdVlutWPZ33BtMmcyoT+m0V3RZYOjLHbd8LciyEVt3B7XvPeOXrxWR1f3TeFTP
cwBhLOcuNG5u1udhzHgPU1HypPhR8xv1Xery2HLFTEdhFvSEB7yCxbH2K0pdUNjk
lNUI/l0NugXJV+KLP6hZpkjJJd/Jb8B7Y4M1GCNNzJ6vLWHqhFWN7XFimqztS2QG
V0bJARZFVnCF8gx4tDUQHGgYWJgsVrkQXSbqrBx0TJ5Ccuvd0YwZ75O7FrQ7ZRQT
k8keJrU6VCkCQi+UagIP74G8RDXt9Rd5/7wzMqnArExjozcLhGz9J2FRFv/WGA3L
VXRZIAFEKXHU0QQHZvWbAVjHTV9QD/2U8prM2P3XIF1UyFuYHYBZ9AXOB1kMty/s
SFfidj3WrPtmn6C4zFctSJNtcEll2Ew1Gax1NuWa1EDjgRd/ScKG9EzYRUZgPvq4
E6V8uxbDleVL/iVdIgUYsP2SqV8qgSGE+XfS6lMXTqkvqa/C5gQxwPTQTC3njCsO
SNoPfl8Wo+jTKzoSYLr9j21XEYEg1Hekr9G8dibFPEBnmKMI51+HNXdoSp6MZWwm
sadSYk/GtC8kHvKqn7xdtSo+xa8vmQgUZghsDxX2s1iX5JuLTD6kj1Jbv8v3eFkD
rQejEm5CegdcfQjuQS3+N8GM3uuz/B8sbM9Fp+iqViYkiu42g9bhsPkdkkgB/uc9
X8LmXgjknt6Ld6pv1Zuiv03+jzBx8gKme+vb3pNZWFWsXTGxF/rJCP59zVmLlWBt
h/lLAxQa4AHxWhMm+2RDsN1tawtlLrRADgBxMqmPSJJyYE7DDqs0Rg9HINPQ8R7H
M1lmz3jf2a8BW2Dy107092h5xnHq24wcY8fZhrWcGB89K3u75ftn9gqXbWfhlfCI
ymr07uXxTCuWh+Ecfi/6MbnhIWoUA0aButZgg/Y7ZESAADya89nbn1EVF2MYmVnK
BxZFuXEPvVpA1H4cdum0BNzHqlpv5qA1iapK/gFqDUESOpT9lNqOHJqTwYQZ480C
MtMMHDZvBU/XD/KnUjwwdjoZq9Ob+Lja3V8aYRrK0dpnQ2ogD5ChgNQfY/8jLm4T
RAFI3HqQBcb819ihN4viZAnBMoYZRECr7nZ+U4c/4PyXC5j71CBa+l41qPLBmN9q
b950kctFqYZXm8WYBHYN2sA5lxaYKSRLrYqJeTnv7kplSKEv+ZT/G48LmKmVlqU3
xfHFom8sEFSUW0Hq6nNWMJ4wDT8Bkm7OlBcCNjldpkjRE2ZwwmT3m/fX0t5ApJKT
gGuc1RTiOY7xva0A4Dwt00/wjqrEC916cJhHXztAyVYK8tyWS1omHl9zsi4kOOKK
j6lNiX0ofpdlg9R8i+U09X3LuIJFM8qyBEjYi/yVaoJWqhtx8KmZRKvYi7g0dg1w
sZKpAvCYqjMO8wFZdQn5EZlaOciy2rIWNJNGpFejNfikvZBX+eLUOYYsFU5PnN6O
c+XYU5syKwUEs37Gi2PEiCAFexp1IZb2BCX9E1KFtZ4QSa90htw8VLDNYU/8+M1x
ll+PjnFHmIk/2MZmvzIXi5+9IeJiWftEUhvXIkc60lCKMdLCNkJajvK3WdknyKma
5rANkOYzDJhGtxxizgcQxB10/B8xdP06cHQ6Q/7s7idnR59W37zWZaPxH/8ndN18
pCiUrYpdN4s8GkYRHNZhEHiAL4KojkbCLzAwx0OHeTBXgzco0wgN3qUfJh6BmcdI
BPahN+xC6ER5x2G27rpip2TEsNyFUcKjK6lUGS88yieRcBWwfqhjyoOBaZlc/7Nm
ZTRF9W5v3+LF79qzCnKfvRFsMWlqtmjk+ayAphZUjUe9wVQoiWyqDIr2NNGESvwk
6dHP67bzRRS9mNgbjn22VVIBkiF+92Qv0J1yvwYQpfNsl9Lbbg0o6IIS583dQI73
yhrIi62A/7Fc2IvW9GBZcXsytbOlJHN0I3WYuKIbzlSsnB7WUj9AwYd0PlLL3goW
2jll8scGbpOTAyvNI8IFagVy4yIsF2xqK8890kUyAIpTPAyLlKiUAU4otirv4sIR
fQQ34sogSigtSD/V8J6ql6P6m/xBuiYAnqIr7TnePu+tN0AknmB2WVBzqW+DE3jA
tRGSUkFTa9mZg2RvXWkBrM0sK25Dz9u+ochitHQ2oYWKIQPQHwsm8x2RH3o5NyHu
iwY/l3XeI6UBlMSw80ETCebPwT8otQ9BEndM/IT+Zq2anknFmxqWG6qEY/2m8sxT
AA47beIsVbhKZBcO2JstSksxD3YiWbxlg/KjwJSLE32LqH39pRBBKMqJ88NRcIdZ
5dMy3F8XTtv4JZHUUMuB31m7ayBncifUVJK89R5J3GoFiiSZk/KLihIbHeqvxN+e
lfCI6HNABv0myPxBZv1iccMNQ8wwnRKl/DTKWobNJnrHmujjRIYVZ45SycND7kS9
NBPAds6XHZOTe+glASi4uy90PDrax2J7xfU7dZP6nej0Njm6H1/BSpJfhmparKnt
lf/Pw8oSuLkc7xANqMSe/8Rg9WeHHKJx4XTHs2Tnw1LfTqKV3fC1FNwO3RFSIV8Q
4hcky6i2mJ6ySr1ziIZzbysbAwwtTyo3E6+JbvEjzZfRbSX98zXqzOtewDCcz6Wb
8LAfZJd7DbdRncIv6+jBdT6iYDiGf76Xwa4dAXf/OmpOiTMQPxSNDCIyV1ev/2gS
GOgKihJtLpkpKla9qTxNK7Jj+V5YmjkTKTu0K1VwacNkxzhORZhzjXkNoge+Pi9g
3EiGvYop/MZJ6wYlYiWiS4fbR4WUJRR6r54H9dt59dJICigLTbrb+mW+qVy/fogZ
f06pnWfxmB1uXU59AGkVJFh9bmXvHjMft6xKed3JVGjaldCGxa3f5RgIIlEDOpC9
QKeQiSlhxoFgsr/atddsoDKId+u+jMc7cQCEsNxDeIQpBEtPfXvspR4cMg8QblHZ
3B0c/4CMsfS39oMOZ/+wNX7FZ7HszwDwIRoHe6Wca8JA56pd8vySmg+xC+7lS4Kj
G2fDMB4bJOz5Ztr03UF4mrSwbOD8up/flrNDXc1qUiHQwllk3BzwlZCKVmrBvl+/
ya+C3Adm6tVNF9L4hiHjEmDeh6LMynnmp3eeZ6SnWN+3OHShm//rjsU50lBqHVh4
tOsDVcLGhaTbdtfODt5U1EJ1J7OFqhWjsWzBo8/EBLaCYyV/hM1bqU+qZhLk0GBY
68gOZ2NbRZP9lFX1iQHqDuNsRajBLZlWsx1rxzj81TuLveuLVEhRrmsNgeI98VP6
RUiyAJAJ8aD5JucwkJ/SqikJ4/xCq9gLLpYYRIZ0zg/spqS36Botn9fWloafyLzO
KazND+07fADODN8SgRy/zN+91wXVSvl85n21wLDked8w+474xMd5XDWK647NkYa7
VYZz+t+itOFUBQXuD5qTXYSfVoYenmrydsWBr5UJBSK0fYxuy2TFSzPYjgIOYxCP
/W51ZQCFrgyvU22G4S8lwpC3wMLReZCnZHzqX09mEbJ97smUHE3TB/YZKYyC+33T
03PxeaBzJH9Q1Zl6oXXKy6GQQbbYHMsc0t74Kp4T1v+mQMf1U1Bn0qizslu1KLQ9
IE6GlPIsKp1mR8ZmQ5IrOaLzg7lzBh5Dw/UolwXK9KfjYzDxvkMT8nOR0Ka3ZEi+
bFdr4ta8gc5oI8ZhObjGzIPRJITFvdaE0Kqxgn8wHDuhCtjTLhhi+zUl+C0EGvYg
4oU8be7rpmSJIpWgOCelEvMfSa28A3V9yP7Uw/tLInienSNnemzBMY2szD9FvDTS
UtbXfVEnK2v/Hkj50J88l3v6dnbMa+gbWpbtmAzfqDpBXdigzHa8yOMF/NfxgElq
DUTzOn9RCBrvaMkeNomFV4dx4TLiVyKOnS6SWGv3oZo7tr/SDMTcagVR9+WCCbsI
iDamkIyWurJCA38EW58zBVV4RaI/6L7BUiOkl2FA+a23RFNld1MrYhhSp1uHnvS3
mzWbEPI3xFEg/YFPw3BGHmT+SpFDnm/eYfcypX8RplEHsl0empPTA4pg7TtLCgCw
AVSuZdqc8xurGvJHl5e7AyHyPI0utha7W97hLcYNcXIRrhoBwI8mYJzFu8U+l0HC
hLN6Tqpqm1B1o2qGZCro8uj+zPdAMMJ6TFqVZDu2iXEhIsO7hjsaYKBhCBmzG35I
RJ3jpDjynApFUggR2gKQIZl0a2pj3+m3uk2wM90aVa3TDdRX6ebxDakb0R/U6MH5
4L0dOr9GjIYx0YMLt/lR6sUNrRSa6NUYghWi8kZqWTqT1zNxpT2DSluz9A5q00h9
DJp0ZUcWcnGfNw1YJA44E2lqL9S2fNQSTTehYC4RmUR3pUzw3tfXjdUOriPZ663Z
xlCtLLX7zXESQRNaO+wiGoyJ6NxBy6jGIFfYKdqqcvdxMoEw+NrZfaAmMvUkwjnN
tlHPuYwAyxNVVbjqQt8ugw/RL1ruQZvKCV9/Ox6KGqx8gwjHxkuJbKCyfhT2ojsP
XnkMjy74JPe3EcTTVWGxY0GHadvNoa2Hui+a8JhNFoD6l+zqKej4jfDTyzlBCM1T
3ZRCti4epNG90uYvlmRr6UTW2c5AFUMVl9SgUfETxR9/RhMaym7AZSj4lZwZZSZb
W4F+Mdjg1b327vgzsHLA2yQK2zpChUcd6yOBzbbccTvsozG2Ju44lGdLloK7I1Dg
G8keoygtzyPvIov9nM+0Do0jyaOOcV1UmhWzxPGK+ibTqYW86bw/yPx7ldtRZ4H6
XD003/fqQ3SxGxLxE9C5y9uE/rQU5F4nbYYCI8oeRovAD90o0000TyZw5/doL9mR
zWdV2KDCdwFcVrwMls/P6roV9QWtoolBlPl2mPR6MpI2eeYc4+YjV1QaODwhjN2o
hwzOknsxOnqoshD68BVysy+FORs4RZTGrSd74gD8N8RCMeuC8UsqrDOw0Dye+9s/
soxt+Jo/TgjZvpiPpezFTfExZf+/n2nLCptMlB8pRkPgr9BsB+K8d7dWjaS3JOS4
W0xj5Qv01K+3P1Sg0TRKgmNh/UBLSzLNYZeB8DeHySPAmXPHmtYcLjXA2rMWy7Aw
/1VRvBFYxSPEXbq0EcWkfEjTrR3KwRRDrmVmQfzNANtrhNS+qkYTkisv7a1+g94M
46tkptXuou+UvHjzZBjmfCWJBTLOBMDZa6AQpXvUzSZ86LVA5+ixNDI6TOceZtQ3
c7eJegfNuZgr7+N2Jg6oMQsUcK86PMqEZlnxe5Pv70plrF9yTUBFBC930RkD82rP
RuFO7QLXvZUo9v2/u40bL1Aisz7YMjZ8yYXt1uBvHFv5LWoqsfGEPtWuu6+es9Hl
f/n7U/65Nk5YFXIDvTGqJSASxV8BmRci40bNaw8eeOn9Yb8UU7m0tm/FYMb6rxEe
A8kNk3+IULhJTFiIprsjaHYPH6zaLNZLFiT3ZrPE6mgF5W2t9g0+VBdNidB5x+dK
kPn78mVhGTwq2IYN6tZ85Lz+428CanVSqUnfo0u9qVEmOmNSUFDj2bYvIvgDC1X7
3Y85GCidgH+05T967zGuZtLylhOhH0AqpgFudJeUAr6L8m+Dq+JGqy4pPOWoHj8T
4JoXimekaljEMD6mQjWhfF9gTlM1HSkIMX57jNzRwLm+097F8cn1shnBSsew/m0c
qn+1/BUJOSD0l+f+FdSHQmMsXHvEOJbvjKrR2ecK6F9ceuHkSyKcmsf1mrXkEAlQ
iu68KNnl33NLoFCEdrB/wvZ06N0M4Jy86Qc7DsSCctVpYncYLC1IQqlNTabx8Uu4
WNpkpd9X2BQN+k2oTEjZlSCviXw9uQ7UOhby16Oy6gYaTVlkfNInQGdu4E0VYvK0
dxmpEek1oNJ09ZofQCf9Lv0isWp3Kmm+ywNr6ZUxfVVBnrKrsgFKvMtk/ju9xJi4
7ZYxbBTsrhXDQIvU867A6aRguWWQozojv4xyJlhGaz54DaH/vUFvNwugH/Y3Zglp
u4xdSGyu04ePltMaRTtS9T8nS3eXwINocGdlS8eKow/byPstCvJptVf/QeMd1t4R
gY2N+daGYa3UIh0z+j5A+MNwkITn5HNMQBrK5WrztDAxrgstqbbYlZfKqWUFDGYh
r1Dd0Ex4RBg0+JRiaF/bCwyIlzyPvZ6xth41d2IDpFBNS0V+SVWnFWaDl6t/U79h
an49AtHCziQEFX8O7zs1jg4P8KY/H+lY4jZ7e1QFB1V5tsgEXGffaQhL4Dda0w6p
4+YxTraOIJVKSorabN+pMdvkJaokbmX+SZpLPoXnYF65jmtg2k8ZqZo/LivutTwZ
6Zeve5sRHT3OvAWL/yqUtzg0/bLCMKfTU0OPpiB3OYIcIpVixsmPRTdyjyJCyXfy
YqzdL9q6epbBbyKwXfdGBF9RxYQJtjngNnZgiunZj86YNGeQLJdd6FdM8lBDJLnJ
Zj+ZqPmZD68Snem9Q9pOvx+O8cXq92sFLq0NH/FUIc2OZippRan0NZRaGPlnDR3E
9UWzjFJn5OfzCJq1I6HKYJgtqGennIVxUNOu9D70qfkG+3F8EvCp9GaC03JSPqbb
J2w46G1w54RpvPoRBN/HhfagoDr6EufqDqE7hx+VGH9+76bVEJQAZQQ8A8b6r5uK
8rpZrZL6eh36HVb2fzJ/MqO5m1+e/w7s3jE4MjCS32Nux4lSOWcA+wCGopPF/45r
nWyNK4HtMzOfGCSqoeP6/j96ibl8oLzAUzo4X/6w1lS905LYFciH0Z7c0OqB/NSR
fMZ3/g5E6Dyn5+7EnPZdin/4XQ2roH9EXm31WQRVsflrUEvdRHrC6lCcBZcpUWxl
5M/lxfXZTOh1+WSyH4vg9QkDqiURGLL3wkqEd3V0Xw4WzMkxArjk7BLe9rG7Xm3U
h9qAuFRUXqN0IBsoGU9cYkAosPhxSwBziWwaRu8ltpC8UJPb0HiMHm4F7sholwgH
fxS6BjigliJNxwopFtOFLFzPhNmx0T43DbsnE8/058MMDLYKAOcuyUXGGPbXDmO1
9lV/4GLfbh1ZzSNW/G78Z+cC8sGnxKFOJwMXBcR8V/o8ZY1AIFJiLVl3mdTYjEQB
WZ+vpiXCa3OEurWiCGlQLdNupYHOAHasGXNw5wcShHqFsFjFEcJrwIauRT98y8jX
zs4BsUKaVVfYid0EOtVdIy1Eroq49RbVFkcG+S4w16v2BCYKBWqgXN+QyfnLTFyE
a9KVijFkKrQsRoE0AxIhDcgoOwSY5GLyJVSNloGU00mYh+knKyXedvWMBsCVAv4x
2PoGA51+Se0xfWegM7ctk5VlNQjfz38LgbQqAeroUBBdrLAvgAR6HD+hwfBdAorY
2IJ9C5kEkX7gJK5KaTiaY+J5ijZ9t4kx3BQM5f6Mc8gKxtJGbslPPlWvv1hK/BX3
5dsPVkCv41w3/ZQ8G7bU1GhPZnF/90QEk5Ci14bTc4l1B0+3GvQt3y3sN3Ic3zJw
7JYpj848MkaiWMiyL3ces1ozVfHnDKBxY5wZLdQTrBMW9EkdlRXUZ3emayWWnO3v
PS/a0Nn8pi5scT4Ykm3lBWWVOxiAZYFHLX+zVcGgkPHBeRHdDnVjAh/kcWquLmHK
LlHIlkIYvweiA+2wnsaGrTzdhUJi03Ep229QZu6NOeJ80PQT9H13ZspwUJOAcu3W
XXhpqcBS/ceaWeBj3X0gPo25578gP2O4DCn7DPO0494Ds1aTxuujrhmneOuBwEPJ
KteOkiDfuHxyZR+/mVOlLXn4DxroRQRpUxihSgsLJi9IQHJ6lon+j59QQ9Cv6jbz
skjIBdzVOIWo3t6GDj2XydqqO/9HCaE9Zn/+604iviPH8B2OU2NEX8UV/cFzBG5s
ATf1LQJgClspisz6Ku7S55S4Z6+Ki6XgfLZaqIp9yjE+2O4/lyCxlKQ9a9zPSYbP
4xGNxTdlsPlqGDFHqB35LeUEFlCEs3pfKcU//UPkqgJn4gtFJNdKzrNpOb7+vr23
vHcFgm4i+IDMPjVj5CPZ9xv207Mucmf3cwdF/cYt+RxurUSXs1FKA3zfFYfqY4tc
/mTsdOBsqPkng4Pr3co2BiY85UTxu4/8m1CdquCnBghl+STrpSqsRF7cnrJpys2l
/xChcZ63EfjKPHTmXWv+UG1kBpi+ngnITewLOCbuLvfeeBFAOabZR4BC8Ua8XABd
qjdzF2BY6oa//xXYRMyu/NxX+o7GBQLm+ePsg5p5pkMPHoper07ZC5+ay3o7dUIx
TZAw5nVTM/jDn7COYrizFGyCCii+lG43KDoefazw/6qiZDGwSqu2i5wkzbe4j3N7
QYiP1rUZCMDlSdkKoWHkeDjNa5ZmMn8ngg/pGo6z4eNdsipbufNceLmVK02Xwmvb
8w83yvHlUme+//AOTwg5tgYwMJz7Xi67D1C+XSanVnrP7EA1vX92wt093Jv+NHmC
7LzrBsnC0UV6hLSuRCzWHAS/hzigY1pHim8cnwifLGKhwo2n87RLvHR4B9lXhP9D
Fd/+kZ9ufQz6BkGaMzdORq5zLVokxm9sMdh1UW/an9hmJaGdm5K5ljweydmesgIj
FTJR61w3VLgEvoWQcC/a9lLwm7SrqR2Nmw2Gab3DpQkCS7FPpsykkxUxlmjm7Rth
vYOc1mZ39+1tKVN7oj9XrByXt7OyZvSRI2euTQwn/zIi/kq2kZgVW5c5bsQncOcy
8CJVc3Jj8VGUPb1VtSx829L0w5cPk4ArYN6USHcP8oCBOaxL78CACFnAbDGlZzEE
OlNFhgI6yOOCkP48ictlQwVYSuZ9ALKEUEjWd7HEdIpRVq8oSLm3WF12EVZw6I12
pzHGHZwDZHjZS8En3guwBesPbf9C4uiYoO4jYwSj//IMc/FHPLqWSDlgknt6Y7II
S71w3kM4S1N9S9COZplkDZueFYkgwcSW1uI5OF4urLAV3M4AOcN7H4shPMuRsSlL
NB/kUlswW2HBivp1zGobApXdNP22jGZrZfVmCg/0S7JFonAKjwCAK9ck2S+xZhPe
U8jvajzsJWc8HdlZ7PFoll+Q0u3/m2eJn2h9bUc3lMsDBNDTTbUqBVoDFvswIrDU
NHa5zKvPKunZJY8OBUC1+dPcU1EdN3Jyrtu5J0Sqr+zEnp7R0wP4QF3GBdySlnz1
a2AW/j0Ol9v6UM8Bvx3sroAVSzFofT5thWYouWGrrw11IcujCk8KRwAJLDikecKo
jZtBTZNXmDSK5lpq/7zNCHK8gtC6ws7hEolyniTC9Ve+5wZl6BwPo5V3NDyzTWgt
Gl2dU3M//LWPi421tyF8QTpYsvdg3JaSzw7vBm8nfEhCbiaHAKfXBrPYFrg/hCEy
McXBXdevEjilLdODYh4IK1SPd9nhj5qDM2mZmwg3eVbhQF3Z0d7rvW3qIakeeHzE
VSofZpV8YFnUeATJnI3Se+tedx0I1qyGhZSDmUSKwBK2Czz+TvWmPzvZfXL+3tBk
gTZSkeJcmZ3mdxIO5ma/bIZfVLAfQKGyirtyN2xlXLQ0eYhsOnWXyLUWYZdzyM/8
pulqcejf3o86fn76cHXsdC7cvRlMCEp0KlHIbECjbbKnxgQR68WLM93DfzEZNKQs
vNJpT2kSTx8wnI0BO4JM+V9eykrLrb5bPUL51dnQAQkcA5wyqauCSz2dXVJui3la
Vpc0a/WdIm6PF56QDmsWSQQ9jhYAhc691f3HJB9+e5OdtJc6GmwqDNkzNviI5tUA
kCSMkLWW/RTIYLVcu/OHvRI/7g11k8Ft+RZech3Usi8Kd5DMtq2Wlpip5mYH3z3L
Z0UePFkYnw6SPlRpquTo/gpGPSo9p+5w0OAdbRht+DAzs688fX0r9XpmnIrX3WqU
tS5CMqgy7ZZFnCuF8QhpXlrTO3VbGc47LwoBrIYoCJqKT32WQEFbchmrhHIt5Qwt
MsJeHXjV5oMwdY0bu5+Y1QBcGjhLvcFOQYJElWkUs4j3zZHt8FY14yKciOq9vL6M
RecmiL5E8KbflgALJ6m/+rYTDLaS/e5cPUUK+j9leuyu6WwZZ34A1tqNKe92vTAq
mVH2PHuOZHGWZzw9DwFJTvC53dv25nNn4utXuFiyDHQq7ud8UH/j9cZ0/tUbI4Vl
oAp7ZPIv1hx4//p8nvI3a6b53WgN4FOc7VabN6OHD/YO9dTzzvRaJ+hDN77JHO+f
IKq2IuiBdf//0k2uqbFkcsRaN70A9PRot2GK63wDMJfzJaeqUZvNGZw2KhXkFpM5
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jNd9v7FRv0es73xJ6oYzFEw1WFwhNBYgLfY/BokqeuZt7pQxrGPu02e63fSW/wM6
jaYyqsL4ujPySM/Pre9QpTe+AbCHDI4HIlgARzLw+UKFLfYpr6ViVP3HAsPpbmee
sTDt5EYRUnFWeUasfphS1t6r3JhpXaX9Eqz2NcXTuJezqlzwtFTt2DKC9oZWpV/K
H/8HoqwrOyoRda2d3idSJjXGpAed943n5XYh7X5cm0NejtD5yYE8RXm/Vyey9qFk
mEMGrwmwwL5sWM8ke8+5snMbTtg6pbYo8XibcpNzuC1Y8sSUyT/ZNgV74c9z5Fuv
UYM3bIgFb5CdXOEZ+l3ohg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6240 )
`pragma protect data_block
AvUBzuCL9fLUivz0BZmjeoXPmwFiaXfjHAhVDu3i7yGLJBNjOJC6VqQPV1X5HxGO
VtLA7b/Jd9Ht2nt+yyBN5JnWxrDApJNupQT0i0tcIpQ4SLEVLpT5ji3ZOBSHz9sL
iZWnIch4OuoJgjL446YxigucgmqsYdeFP2ym41CvK0r/DUDW36oEly+ryCHrCohB
PvyOZ2qpidHRQcnRZ6lVvmSRKNU65gjAAw5XVh/90XPx/pTAVHVSFeOMT/8Uk8ow
40/JRT7eFWeg1WnrI2Q6gdeMVmcKGRFfV2MNcyV9IwVQAtzK7Nx8AyoZh6rYPc5J
ayG5EJtQor7+YexpRxdkPgYL3PeB3ms8Eivhyv6h9dxP0BwSUgyWGb3NjBEGzLVQ
Dn/S/bGtNbiHGzS//u03ysJGX87pOMzKPF/lQIqcvXQY9dBzspDhqRyjWW6QLs+1
uyTKNX63BjJ71pn/q1Otk6y/fAvMyY3PLg9S71D6QssZg6GyEnJ7O/4+QWQXnVB2
WlANi7U0NmxD0o5+Ngj7IuxYtb223JaawDfwrV5Ml/fMs/fS9WBZn8rO0rZtWjny
E6nERUc2CaERFWQmVL8/V0osLc9IKuknLweRceZHj5bkmSLcBiOD4jILaipiCWBJ
rt/S35LgS8CcgOV90s3fOjCGAzaezK5HAb4c8Vo0BSThXZ4CO1d+tXo9IeDiHDwh
x914Www0D6uJwnkNAOZX+6kAr3trlxz4dm9oZf9U9LRq6B6Sg+S4x5TENQ6Wlsfi
Dzw3QUVCkCQpdMEsgqAGO3kvdRs6y/wUbEX0exoPyOFeagKLn7Y+3OGPJnSzuDK/
/RTQjCwfypFGQv3w9YaTew7PTIBIq9izxFcx7+6LAN30g6MyjX+8GTfgw+2CPorq
qLdEwO8sVSwHYyoSXd/HZDJivQs/XWRBQf4GdzS1Oss2WpUy0nqBPptPC7p1MB+6
RzPS1bJpk7pzQO9a+cR+fiVkBiXBkAgpItaEsqBwFQrdJy3hEAXzAbCEhP3O4eLw
kawkg01YgrVakhwHFWqgj0J9IGxHEBgVTW1HplXohVQbqMnfeMTry9CWOw5duO1s
nVHZKxGmylA0uohI7R1PbeSOWGC2iZl4MGoXOJj6ZDWFO524vK37/CQt2LD+svMs
B3OEAxTcnb0KuMEj/DFoWAx5vQAW2/dUZRij1qWGBcYVisnV+xY+F1g4IMYi0+d5
6D6SQulu4QbBVKMDJ5qpXyNn/iQYtjecHArpQ2+fKkdsRwLCAD3zaGinBwgISGCn
GKl5Zc+nhHxYviX4E+xEdwlUDI2fYLhwSf/QYny/eHWquXCvMrFp+TZGln/4rqw/
Or2BofUVu7ZPZ6gJ/qIrIo0ZP+7vMk4ozwzWrjrmdd1nlDmA2J6v16XFWUVfjq9u
1UvOuuyqbklQP0DP4CvyAFh5CxBZcQugPJ+ywbbSl7ONDRmhX7Nq1mwIoFstpspW
PQBDOWznaKj5qJvLZH3NPoIc811js1O3e0ecJ6rO/5Lc9CYbnwLjNITJ6wjWkzC6
R5jdcH4Qr1o6oX4WukUgaESpS8GNpgRmGX2eBZqtCOHGzXtkF7cBed0q5/cT/20G
qpYp6n3LruvNMwzc3mP2oVdjhvGQDLOq0bz02psgPUiu0wI2TG4krSFDQUHcDnwm
egaFeroy88IKvzDo6fmIjp8qCmfUjikLJ58E0rU7Xb9M1ZRXVAnQI7wP1rv0iKO8
m95f3w6q7Ty9zY2CaHfngCGWnmbXNVs6lJlNnVSu0kh6bBP1IkHIqdEJMQZNqIi8
WEIshrqDa4MRBr8IZDqZBU7Cy5l+KZ5vRupZifQxMoog4EXCB9AQ7Qk84VNBB1ic
LOeX/kCUVDDFgyUTl1vjom8VwYVbWeozC6psPANDdkoUCvV4ZTyQGstTb8k/quer
GlMv36xF/vq5TpghX+M7l0uv9UrMAMcvSGy86/huJ840pFoqA7m3O8ZjpB1EqhGO
8jf5eodL6JwbZnnD1yxzkU61b3CbHZyyyqkgV6jH2RrQLsB7T9CHtPzU4SllwpSc
eEfFGkGMWfPRslfzEgi8riGkNRR5eAnh+fEsrDJk3Onk++qc3gLrsQ7dhws8MzzC
6bQGPXc5F11xeSf1bskHjrkB7jVBwkggz1ESAf2Axbb6EQ2ZsaSsCjnH8ilXC/5u
Jd0AUUdyP2b34qHmYLs+qeaxQGatb6czK3N03oC/zcGqkhLrvbQ639bFfz5XRNGX
VjbJGovzoD+w0+GeRk0S23LExN1LrcSTZpcAPN3j4F6mBhcN1b6SX7SzUts6oo/l
rGMlrbWvupXZ1ZcuPGgx7iSvtEfZesa/xUvBZrw6fB25pqdG/LxpCAX8pwH89TYL
/rJfnAtKKVMV9RnZDe/U0fP5swmyYjmGaACQx3shlKlXYWLHz42Xp9KNWT4BCbiT
c7OFkKXkFHG8o1uT6kGBMejpyWLIYiSFI96SX7unPwnnIIjyuZfU0PGGQya9pfxg
z3rX+63m99FddLd15zbgadspmOKwGwnH9QCBKALD8Bigmgip35ELGpNLc3zZLUZe
XS72qeZgI2KajcJdlsqxG1IxCJ0ymC1dJtsnUo4kLuby4DERjthZjn/Pcx2dlhcq
cTzV3lZw/KaEAKSQKWneWlrZzTIl9ENDiNqylI9cZEIm8OCezfyT9poyyMsto+e0
QsZ24S9Q4dHVAtrgwfHEQuvnNq7SjEYgT8I4CL9hIgyUWKEJgHvbLYoVoE3u/Zod
WlWHhq6Gyk1Bsrl5uME0dPYuWBUcrBXfPt+YVPothsLPDSYNPtpwC0um4bclaFaE
iauOiOPkD+3mmuqS0xJ4x8CuVidmvhciPZkEZYCSJYsUk6Rggf4715S+zc1mLsSl
h6bOtr2V3EphqjQvXkZx8zySp1+8MahcsoO4rLEyk/TPf+Wpbp6Ohe/vA0d0SBrw
yOs6rfVD39kndgIRHjfGWmVLUbxzLwa1O22RgDyvG1qcmfMhleFUhsaU6h0mG8Pn
LY2YTRslaFjejGtEP9F6ZzuHmx2tbWts6sME2LA+Wv8vOaaQXab61oKSiBp4vmxm
UC2Tke7u1OZeXwyTmWhaUSHPlnLYmdYrAjHgDDLZ6TdV5b9mijbghARrMbxZua4C
Ae95BE4s9rKnnmwYcaymqfGr1wBhxM3mTcQPsxqf9K7/JcCiv10MYAEqQH4veUe2
bb7XeMQy4XdechAYzrPbee+KfuWioqcCX6H8LzOf8RrmJxwnjfoRAIFL2ygqU/1A
X39w8Jw0gyDViABUEVxk54sAfEChkxuWQpICn9tV3NxHb7bvaDNCJa1FLSrY2o42
rBAgxULgibI5hMljC66O3a4kfviHbgC+prJ2n8L7/dMka3UhPF927STiyUmlnHzl
oSIFegsbn3U/Cp8Athd9I6L9nwnTGtCQsznZdEgIsxJSXKYXaRrJQ9JpVk3lmY4Y
6IBtghwNjACbRayIBW+8wFks9UnhdgKU9vM/vKn3MeCee6wQDL2o0VWk+aRENxF/
FXSTKDRzyOm/6QpvdlbF/tjE/MhFyrk3V45CKYwb+Zzt7h2YGEAZXCUEGh8pOqsX
h6xtMawSnA6eFQO7as6e+Mc1FVTQaqPE/lyRYoZLGS1UDG2vYXEWmfZKJZ8yICT9
FeHz0CAI8tYdbzelBZsMDIcH0FQLCl8sR0RdyHC3syoaAt80MEIOWS+eswthyVcN
R7Y6o+a8v8HtSfGIqXfKNDJdqs9rckfntjJy99A2zbnjsMYyo7ZKxj6dzgrpkCDD
lFY5tz99IC5FX9064EzMLR8gPMoontLhg/PPa7E9JOOw2YMxFo3qkh4dYo27JJrC
8itErJSFi8LEjJN4agpVrDyeldVSZLKo9GXXUr/205UL2IYDw832CKcE9EkUvp/g
+SWTs/yk+REUQPbTBOEtwsVQCQNNUXhVn8yzRZhZXWp0I2+WBYG0hLUAxbqe6rnE
GVLOTIqPXFK9dJB6YlY81x662CYc2sbntmlw+7l6YAyZAQXoGjCpLJD+ykWHT6KS
b9BeTNjTo1ZMILBHrAGe6rcm1cRHtyoOpwkLxFP0humF0R/h96pYpQu8MbCnI66Q
9XkpqsGodGbUVzHqWCBMwDvwzKnuowqzRRC761rbo7dhbyBmtAA+mIIv6C2C4VXn
XllfV1hKeRda2xi1+KaRQi+zxLSueVX6fdz1p/Kfr839IMiMU8QP+zKL5H02wSkM
tN6x5A2FKFTe/RXlSrfanA8HIetebJkinhXYNXWo0BUTvX2MZD6jh62ssW+Zjx8g
eYV6YxikVOu8QuWGiudRhlXmPjZmT06gCiHz1O3VSw9K0oat3t/TQ9uaSaZh5Kc/
grChrV3Lq9S/+XEZJaAnlPsMTYXv6dJZ5krHrfPWh3mS0r3q3lZdmOIjO4/WRGas
Yhq2LsLz5EVeAr/e4OvZrJrrfOEc1QKy4M/OU4x4RpmGURab0nrSbF7IWsjrP0OB
picShuhZ+do2ILjsbTOFsOLtbfGzomqalIgR08+8usm4pyCROENGBYWwiN/Fdzur
7swInpNqnyDS4ElgACGTj0KTSFiBWRNhRqVnGm+bcN78kRMvVp57OjIZcWPIaJiT
p66mE578iS7cZ0+nAcs9WzBHABS6G9PNm0Ry6D70/1w44yyZctHu3oGejNzy+8gY
g6FAyh/qdS8U2ENCe6nDFISVqIF0v91vBcE/8CWP88sopI+KWAiK6AyAuM1PdoqV
dHlMsrVIoLiH4tBKSv452oFscGPCO3KWA+e1pDq4L7A4dxm7SyuYEkzcfl4Mev30
/qenCXBWMLmrX48Va0bHNlLYYw6yiF+O0nnVUj+ihQfKQsEjOPJuYQmbmSyWDzBU
GlHG+sfWWtPmN9QBnH6vG3fWbLFprLt4zwtDVqbsVPsSViKfdZdyhA7hrIukmr0I
0sZgbF9F3LMPTJqBHAD1/en0oT6A0OQWFLiH46YTttZ2HmKnjJji9kTL6jgNBV/X
C4asSEXNlcq6EuNCyj85rBOcH6Fwp1CJJEOk1J7eeKEwiry+DynyLACS5gmNC365
ETOaNL8uWiqUUC83y7Wz0+yVy1TyJhzeCyRzspOFHGQCXWFoeHllvEhFa/JNIn+C
b9cHEIv9j3VnUey2KIT4DANgZOeJnwD44qQ2cSyy5wuMde8IJeJhDbZrdYgm3pPe
pHqv6A9nIlHGtB7fZaCd3uBVLfs3z12UL1C4NT2GVW4zDl+RejZSsa2U45yaHYnM
A8hYeR53FpS+3S3+v9tLOuy2yRpnXbb/2/sH/Onlr14UPHEVmqiHf8MPRIdhQdU2
NyuwTJ9Dv5ukWYLjXLKzo0idLTRVmsiHt5/iUvsMAojpCymXnnuE39xVKWx0rs9r
N3MfNfwM3ej5VRJ6zK/11Nj9J9xal6YBwo5DGnImRh92X7ibvNutTgsycpxuxI9m
NvcwSGOg+0bdaqhNLczXMP6lR1WBkkSFeSnpxyF8r7xYpDp9ANfnbLFNK55uUDo+
Vh/4B1AOq9AWpCcOcSYgIGZ8WPpinkpOvyQ4WDvdY5x4Vk5seqbcat3Zj+SktWN6
Wwz9kyZnAcYkIKTw3IzM0AhEqriuNe5hfiAY3AKbGkpCpQc1qMzVLiQUj0LRSdrm
Rm0zEpJheYoOUBegno9fwTWQygGu4QJ8MOJi7E1Own5zXVGb7dA5EAa8tzQ/DEWA
TVgRH9kz+Fw0PCdZa/6/z6b+JOjRid6BUxCuEA5Q0SaV7ZbnzNGx0r/4hncUAXUq
qNTgPhFLu5mNCSEFTtkgVofN0EYs9xj4bQOOeFwhbiR4qun8aulCi5MO/oc49+Xw
HFs9hnqhxNOXkobF2h+/K7sKL4U5tN/fxfc7nb06cYCeJDHudkoI9edf46s1lE+x
qZnws6FI1LDX6iR9LpOm3973sNNgM5CTDdfrxXTdEcXCZLNseaf7WCHQGGcgMH6k
Ei+kHSruI160n+LRAqaeg1K3DT51fSZsNEGZVkiXJZFV93FjZKJJI35tIule5XiA
NWECXIrQA9Nol0NPLtrLx/Ujig7+MkVYxjZ+rKv+FYM65XEyiHpZZqPLVSDOvmOW
SXLx07XfXlyeFRxAGmOjmawSX7eN9SeagM41Rmw315KBoT2oOQLs+YXeWi3ykioy
AA4K0cOywkWcJ/wHcA9Vgp0t7DJhpkopwoOd03QlZNaPrH+w8Rxt1ynAZeKu8rnU
cZlTtKJrhef6IwJqPL17AjBbXFlEOftBqPIyAA4SF/aJ4GtejoCg3e9YpLE8WJhW
JnBIf6fqm6lqfFIfqeolwBdMLYwxQDz7XCeSLXAVpyI5ItjAxDrpwfBQ6djSVXuA
5fxkaM9dE3wTYWLcr73UsbvhUqCPseZEndyI2SEXhSLpBaUu2UMsI50txfXAilNe
y0b9wM+th83GHll3hWAQPBmf4/AIMmcBMT58VEyyPBXLiEk9PfYt5w25hxZjY5ld
Pw/Q/h69NkmBic3xFgBLOBGEDwfASWpY6dMY0jdrnDqb/PBCESMFBqiTYUHeNSht
v2jHRVHOUy5C6MkJSfvi/qJos7yFcr/rgu83G93RFwZm5/1nfZ79jG0jwFUQR34A
ce7vn01LWC7m8GjKdBjQYvxvR7OsnZn2SUe5iFF01i4aeYOSwHTSCN0BhROzoct3
ST4cSttQOFZIqL3GAGRIcvOYIB5zCrBPQMJNAoClPtlxet43rUNi3cFqtM2zk0eE
5x4H9w3+1f4egIvbv2Vkw7+RufSvpgqXH9Kohqoq075JRSAiUxou3WpMyJArnVCk
pQqyPWWsSNkLrNkuI6amvn27a1l+DmxK3zWh3W4+udB5eL34XLk60h8VrwmsIzHQ
v+KCmUIL28xMdShLpJ/A9xcdjD3+4lDvO/UBa/Xp9q2f8K1+xQn7BqwYiYj0pw7r
eyR473IgmOBa3cjOXXUPIF4lR/O13hT/A6ddknp4Q9mWLxzdFuP/4m5PDk/yNH7h
xcC73Or6+iyfNQEmZ8HRX3X+fUTXzSJt0JQQLoaswEHDPCllZqJIufXJ/nZo+uAv
Re1kQXjKCyc+LZBnM7FvNs3/n6gtMADdk5doq15JAkOq/PpTiXeCI/D4I9PTnNNq
SSpBYj6Nvjd0FVyKYnaNFDRMnxSJx2Ft+1Q4khC4CpOa2jKO7FqQRYndMhrED+UW
4M8aJEa2El+U6+G3iPJYh3zD7C11LJiKls0WkqGcRzZSNx06QQjdipLNGsgH108A
BwIRuJG9x54DcCerRziRQ7/QLzH/VSnxunJWsBTvVu/cYTDMyQZ0CyiDt1+SozpN
QzK5QGDEFvOI+kAOU/scNsCx5z8F9ZUD9AhgDI/vDeErK5wQ+CmLtV6lWrqY3OLh
HZrKtFPNs7df5r90VPHRHPoTpRUQB31MM8ZWm97fkV0bYuIhLbsULEbdX9ZkS0OE
gB8fp7UXn67hRuNafc6CqnnWowNAbd4VvBocn4chRRZj5Wt9w5OZR7TelEDtfL4R
R0jZDMfnVLAi2b1k1FDpWwhHqHDZ5UcPEzPfn/Wsbgqhkwp/J0f8c8aUFkkOnXuW
sLuSX3VZF9KzCcGjY6YYQj1cFw0YrvN6HYWRRAO9HJIXfV2OmVwkLh0cMEu6Y5Tj
uZXuOOvKW25I/DmueKKiexpjzATK5EggQGOdiA2Ebt7Zy9rajEmJVu7cxWKcqtWf
EFCpbgQKWsD1JiJGCF+/EFNBG+evfU8e/NelLE9oOgOK215t5zTEgDnMBfHt6ULE
n4gdxDKaZunorSOdRVyOtNsBJyTALu5sIjhsGhhC7+sYT2bUCRKUg+ZPLED3GR2o
H096gpy+CZJv/Il0Zei5j4aNzpR5IykJsWnxalkwf129pDtP2zgAEdxNUw7rM5b+
Rnmpy5h/8uDd6Lw7S11q6a1ttCmyJcM34fv3Rj4MjEa8OpGU8SfDabR54/MyeZjC
qd38yV11MBUTDprw2MoUKWtK3AZEQvByUnIGJ5+9iiKHfVUYf4trmEzVhbLZu25Z
b1DQnDBEcbr4HlxYJDwW5AN4QB4LBKNOMjJsS9EIRHIQ8YEX5sWse2QSfdN+NREk
q1jBPRCwIKeB74D/hSl2H1LbtY+SaqM5OUmjg4t89fb6wSPksEgEaBtJd8GiwRKp
n/ZU4f6+81bsc1+PMqkLd+CTrK+jUuZQETXF3A/lQYl6YOPSt+ulW//J3gxQbVND
9MaoB2wItWtqC5PcEGd2xohMGP2j9vzTo9pZewf2jYS2NKLB8bp6jbLBUQvzxlJw
gDI2fZBuvcgoPpDzUv+h1CmBcp09gm4BLO8INcBI/C9fVzS9uAj75ZJyt4uHstof
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
meHp8gpNNCpouo9uvt4xyuOSn6Ng/v5ux3aoEVHgGgaCRsahFuhx9/Jz/qxXUzZv
pP+VyHtCUQzHufEMmNM57JHjz5ZIp3N1ZzZ7K60RTrYEvUiNluzQQef1MFHCzn2F
YUlb0x8NdQsdvRGxq5Pi87gk8SARVxlZFRGv+0Nwf4kOO03pMJveE1Yh5Myubzyi
/3B5257fyW07ttp+s1G+50xFBREiDlzwi0Z+zNyFt7knD+s6me90zzi1+OsiRVtr
A2Ebf52avQ7p1bWo/lHScszbvXsLeoWPExQgeRuiewtCrE4ph1GkqEtkF1MfvOMq
gQjC8BXT5m82Ed2FGh4I7A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9456 )
`pragma protect data_block
Epx3YUfIiG4yPuy44p5qhF5EkKBHoD1F9IHH813Q0Wd+toGXq+siWAxN5WuERrqW
ybgn7j9Qk8o81fraIRq247B8nuTAs2KknWdrd7ZbAd4mq29ACMr6FErr0rh8cFGe
r/uef7YAc3PK1VfyitNqU3prOo5RJTeiU0ITc2vmeo9J3YVLKBoMix7c/Oe1JpO6
KntsyKs+CyvnLqDIwfRMdGTu9JuOR5KsYX4VQut0apyMHlBD7IoX6lQUX2A3YWOp
U/jqHCUUEPRTz9hYVoFOi2MGveyhJFANLyg9qgDWdaU5HnyK6MM+pIhFiYs2NPQL
DPo9QAujcHLgJpQVkRvyZlK2mbwMGdhvnQdAbepJkX2syLEigm385hoFH6zxnxl/
Zz6alijVtVbNliWP0ZUc+HqvS+ekY5t7i/kbf7tDC3yO65rtTCH/Efcgvodd/AN9
2okFSLyBKTeF9WnJA4q2wfOWmi9fyQyBK1F1ct6VNAps5GCp8W1e89S84M4j5bHw
9/Ckrrw+C0J0h5ON3CYtNDJHw67MjfgI3ubEkW3mUSCdUPyBjcCpM3isqVdcFxhb
l9Enbo3kVThJlJ1yvI3uJ3TzsCglXfxDqXcMCueJut3NNeRWc9pXyC2wS/+jiDLg
ZFsNndCg0JS0pAEASaUgcgoCWyJF6CrFfwnbkHB0w7KfsqvYOq8RdHrcVuuNZpXg
shy0FhVmAzOxoPtqf51ocrN30QYqAjg8Sahou0jhn2vzqvkcnm/Fdd95FPToNVvU
R+rjXUeqCXwIA8h+TUHIHvHdSWDPX8tZU6kDxk890qI7dOsL0qH25whByBDELFwL
flLIMBPhGgjDZyY3upGmQRbRmvibsq+PyQouA7yQix6dNK3Fl1DWJoKGzGJaAr1z
0MubjgyevWkpgiTpse2kwu3vusWFa1mHaFPvFmEO/6oS92dDweJ0wATEaqVBuDhJ
AuFTT05mqdUhM2beJzhLU6aWgzXiCwJEGdF+f3RoWmWSnCN3dOX02tlFliIMQKm5
nvyL9epRJW/+dNamAxPRDZeTj8JNSVCLByC9++Sr+pxjjHOslkCC8TqklG1m1UgB
Mz12aGJlhWsixkxcKA5gdGOBdbXFLm5/p2CXcS/VPCaFvMDPL6KXueMCyxJb7NqU
q6hDae/zCHZryftp9lYtWYb72Wa+JnAayHgrdVHTYPBACjxbbiyPvE4BPBNbKT8J
xez6TsxcOSUvm7C5QbXNc+4x2Y6DvI7fM9UNIzJqpL50pXn0cL9hMJlhof9gABi9
6vir5AGq5gD3v0AZqehJXrTonhbEvpRbONm7D3gyTdxYpiNzGvZAjuIabDC3uWpZ
6svLbkW0mJ7Z2UvsXZTILmn19LtXjfJOH8nBM4aGjTMKrS4ghGN0rjQrwmcZvFKT
Pt57mygqUa+Us0Dm0TM9O+ajHI3jubfGE2GMc9exWPeE30KdACIabi+mVWswOIJN
bLQgZD5y+Nem4SJ0YlwF5SM5+r+CSFNf7VjAm4o5yjAj9VoV/JlPdXZ7S2+ImvSg
wJ1TsVWLym+wAdrEdJxnM+brUS8vPKzgD2fij+YaID6v3YmNhukEBwxsxevqqe/L
XVp+ywy69e5goknUVkNFa9YxWQz4eXpJQ4uUtr6gSYyqn2G9bWYFA/KuQC2le2iV
kDVK+kpX+HH8IShJruS80tV1VJqGZrlOyfVnFjiKhDx+99jQEmsek4hhjE4+w953
PoNdwN/+sm+bs4gHRJWh9fRr4UZ83xpaiVrgvWOskMKdy1QR87QHHwaN1lXEjEEK
LSA+gJtsDB9C58+/8P8Yaa2BPzYsOkCuyATdvM1yC7NVcwWFvPnaVip65QYaoiS/
pZCNcyDdBodTDqWYMc/RP6ywoRnIRe5S+i58Gw2a2UUfuxVMUYVpo+38/EhWWBvB
kastNUXjybTkTWvmMY489hjUV2U4Mio2iTvCb5hBDRX8MKdkVa5uExmwj5xirui1
glzx737ucQS6gKCB5IRuns5NAxqRhSnhpVsopu3YzXjEW8yoQp4mdGw7tcQLyuG/
2nLOYDMTzXGobWBcQ6awVGSegxyzVunrc8yDFenEjDyQG36u/lbLukEkvFqlhPyf
hQfCqWoGIiIhTnCCM8igPBTaAL6oDtC9fzRP9AnV7yFAVrDLEZgVKBqL0zH2e0HT
Mx9qDx89mwrII22DnTqvQgB6xxBJzCWhwtrM3opsUTNPIw0DS9r0YKoeTF3qCvCV
npvhkoB10W5J9+DVFzOcj8+zpdgbbeZdWwyU1vgDyxIx+DVA70cBwdrphZUz22VD
bDzeUzh83eQzpdZtvWmleHsIkglbuo32xct6Emh3PzwmTcQTW+Vy4YhhLCbvBNxY
xCWXu8G3QaIwbzRFL+4Xbsg7ytOhmx6lpn27UDNvAJK9ZZmE3HjmL/NFwR6Z0A+s
uRbPUaj6LIjJAXDQp1O8Jjy5Z5fncWhmSICmeJyWlld8Mxq7lpAJcHH4KqTqvT8r
GbDF3liMDOfdgrAaTVjLLDO1Xq7Y8oEPVRLyP7BnIijAMKTk3CrBw22Iii5Jx8BH
VtSFlNveThVIv0hb1SbyoxYh/BZKau3jDXz4/i4PzIXU3hEmWEM2ovXjMsC4PUhH
dhEGLIZl6G9MsDIcVagHnoHZk4y2rrDCmvtR3L4l1rvKBt8X/rZTYRHlaSByDF7I
VbW5c8RS+IOlBZqJSBEuTOgbkHwTsLfxyT2GuVABw+zndCFsNAEX17l7cOr2JVum
92hHAjadRzPV9DV8I62dYDZt7d7uqo5f1hdRY43UwKDYKrJA72JYDR0GoFPn7OOQ
24Bec8YTVPWC4Tz526z6JZ3YWHkn0box3fZVFblCEHaMjTMdgiHEHgk+JIcz04GK
Y/VQrI5OZSjm6aHsG4Mp6N5gP8e6J/HbKyyNDqy0apdbs9n9i8t2GznddBipQ+ft
K9dvRYGwCxRs1LVooaRtexmzadKT4itwaawZAQ2T5t8lrAzBNi+GDCfMews75Dmy
rUm5TttJlrdPfG1zhS6WZFSMjW2d/ihFWPETbE0UIUm3SpvC+/2BezVN0af/WDT0
gpkLmJCRZS3wdjUc5Sb0e3vdyebY6uuUOAcjALQSlFI1UA+QbNWOFT3gOfWHtXo4
JFg9gNN+v2G+6GdJFretHJQM8XK2DifpScY9m/8o/0iis6LpPQWc3yAaSCYN+BEf
eLenle7z8tyFCdYIBDlgI3anerOQEKJxG0zcJKQzEZuAhVDnt9QnMbbVrBOSe1tt
9jrq/2vFyPFJ7mbMfAltymAX1IOlvqWwa9j9jpFvB+DxJPs3JL21Fm/zcWpPMu4+
HdDJnwNvFyBKy6aIax++d2t5/BEywV6QFQEuwIeNIxTnLBcInG5NFXz5KO9j1ao2
BZnYzKsoH6eeIkQRJC2ezcN/kBxw4ryqocKSpcYbFxY5TB+iwmGMsGEvbeMLBPFl
vQx5G9Xru6YIQMgWM7QyVFGOHUBdgSwc1GQ9IZaQUaEscL8VobGee1gTj+ahCDwW
0+db5ny6BQ2TOYiZxa+xjOhwfn+wWNNchQti1XxxOC6FL470GMoqmlP694kgTF3J
sHDMB+B+sEziWe2FwzNq2Ki1f2F0v7QT01VleXTfYV16m1spU4V09OhqDQjYmnIw
bS2K5l9WDCMC92EV+7ZiM0QLs44Ohxzhfi+L6PgMujYkxseYSLVvu2ix6UTTzwq8
oRxH2TD19yEaftWjWiY4g4+AOg34ftjIIGeE6M1lfvwaP0rmQvzZx8wph/TAjPkr
RI2ED/izyEI0j7DOKkGadX50jZ41nvr9ouOhGSuPcMeY9LRs0qMkUCYpqN8EHdso
VV6bYYT9TRBWLYb7R8cqa9dY4YxgNnOznvKbvCM5jE3URZiV3SuS5SwUWBysZNv3
EgtVA3BR9egop+7JWs3tAw7FlhYf7hpf4q/unlsli0abmu3JqhHyq8UjrnzDd0XQ
KABIT3L+V1td1Y/EeiUHzyCqbDZgVUyB7PNgkOaCGQt2fWa/0IeB31XvBzbWTQxO
NCPGMOzn4PswH1SqC2PP3gv1v49s2TUyM5D6qS8Ld4dxHNw/tKIbX0nzv+1Wz5vO
kijussvUqtRiReCVZxDYqfPFyD2FzHXms5E0oFOCiSuWAlMbIrJUbMxKG8H5a4RR
mjzeoArkgKsT77o3gNmJm0khSnE1yA3KvTybHVcoek6r231/6tjzNnr+PC1MoEWs
OcEN6uMxQFdSwcn/TWwmLcv9WHHa5dAbQPnHsMCv4ANLYDM/cHJcBOY6sOtdg11q
0mpOdCZMyPL4GsL/IaK6GtL9VCkS8KjhXlUYmqx6S3hAiMXY7N3e+WIuP3HlYZBd
++9SdWLf1F8rvtzVAOqGZnGnC7KxL5mPaXqG3scY+smsyjkVlWcGyiPyouuQU1xj
PAI4tfxD1Z3aJroP02537dMlgf+GxMtd/DGNGGA9fDDB7KTtvd/gNGtyNyIEufri
ED+8w2s7zEY6Qj0LBMjE2u7P66roe/HF+Upzg+6sdFbybun3VXnCzRGSO+EwtFK3
9ptlmWDCWBQecyJmmADNGiFFPCnFo0Ju9jaAl+mIJmJ79CV0IozlrJpD92v+kgUZ
cgj/YI6d2nGf2YhrbxV9/L4F5a/2hunXO2sdNA6FfNDdbO656drI4DyPcKGxq8Gw
VhRrmyOBULm1eIOsdGsI4XYCsNtKsFD+VRI4xmFoF27VSvKb2D/6MVvuh7b/M7OK
Nkc1aec4OokpYBgJUqMqOT7KC4zCA3qWLrsBow7eQYXhplGoUhbu28nmvSxxqWxD
DAT0WMdawerxxrPQTCLWh4NKpVZQTGZke01ahCF2e5CFWJDreY51fB6ppUnHBEzS
byLccLM4H+qw3QheVhlDWHJLwCeiA9jVltswcrdh6eDbvLH03hbmZmMaNBl0ZEWz
oByIcAxZ44agWbVgXlW67xVEWE5cflJPKsQ+Hbcq9Ems4Gy5gQZ+s0zEEo4kr08M
c72ce0QG3s+CH5LLspPUm8N7CgIvej+GN8qozlv4eftbudSfN1Wc5VuOlOGXGQfR
PPKfL/3qjIkinKtysiCQikZYE07hcFJ1fm8z4P0mkgF17rpHQ6wbmYJGCO+L3eAT
nSaj8xAEl78QnRJGMZOBZ+AvhmnhQNsDd83pLiPJUDABxnh27bQd+e4n1ndpQ/WX
MOAQcc5TIFPS7b+Xt6fhJcfUPETPuQPk8YaPyfGFR/G6lZDWgNSgiHU/0KioktMy
JZj/V9bVpQtOriY/QCE2lFyZhzifSrWKJNhyhAXmB1YHCJmLrCzpMBYWZYh3iyvU
cvHpjG2yk13B7sQd9xPtcmSceHS8hA300CaMlLLW4kLSXxfsiJOE0DHoJ4kl1nvx
UtFgreruAxKOdyKYAbgiXLR56gcX2jWlY1ZtmS4Vw6XisaUDGsc+Y3Pa8QHhy2TO
xj6KJQGcbzjWe4pkNDOJUuqGjFfCaXa8G4bSNw873vWUptqpTWKD/ibHDohCWVhB
xqyXbBqmx7PEsxgNIXXNK54BW6FOcsM44q02GeBwQfFqbDnm/0N7wEJW61Yizh5c
6w4QyyQsmVBXKx3ePUcvHATXDCLtf+oGn1YKM4fGbmBp5rKEj2MeX0/HZ21ErwBy
zargybjlRVSRoqZJPoBmlpZcfWP8kR/cfp8y8+yGlXReTksYewA82xPVKj3T3wC1
M8cLMbxDPidzFhWKKOaPAQtdTbjeqcBUs0u+HB5RcRkiJVRScolk4QkFnE+bpt5g
Y4jRckUk+axs7OFgZ7N1dNZlAJPviTBC0tut5MxNVqKuvvVbPXNNCIH5n44Q4U0P
FwDdMItTfW4pBQMvSx/NQOE/HSXiiaEjqZhoBKzNJ4VTu8/lLiNiwiGLbIlH2i6A
icgQWm5TKvefFUxgRkY2HfyB8+45AQjv62sgTRI6mG5t1AlNjlwlg45VIKyrTW6q
3/wCm6a/Jqghpjw8W0RhF4QaxJJ+zB1DGDToellNBPApGworqJrQ2IwE5UUoqjQf
vGIwf9SMvIYU3ZK3Llqj+IxhxeReILAMnycZJhoMxIcKgXj5pEXuZ8IWnyKjXjLm
A48AlpO8H5BYy9Mw3sKWi4xyfpWiavvY97O4o1ldTTuaMKS9Lsynj6KKhQt9dip6
LvAlpMR2UCQMFYRDWCQ2LQUfS8NEx9aBaO6egdCf6i0v59EZqWr30Dl/GJ3hD7sb
7U1lGnv1H6aP/N5DJ3k7CeZloKE06VBEbb/1JG+ikPHJcMJkUPLw2SthuCzRAGGh
6yX5Aiu+AOcYe9vxWGQyreS4x2IoDulqqxe6HUJFmOaHWz+0IBXKZ9nkLLl9FLjt
e0Ju8AOGNLx7vH2AskLRE2ZrJKumqwHROgbzFjIDpX6N6MGCO0rYzjtYnyPEPZnv
PZzwR/9JY9cv+xhUgjzjCaFOxZVxXnWPS7akP3AaFQVBUdFxBxA8LyJ1XCOM19iK
0J+oeyLXref/rn1VkjKZBZC1nHFW1sD/XFVES9GQXf2bL3Hpo7iYekVJ7ixYNUtQ
6RK3FXW7nGF6S/NYZaR3Eqvf5nMWL54RtTai8QHnUy1w23rlAqx7a/a8mJO5lwpI
d9yE3tLnK5Y9236fFntap6S4lKfUaLzjaZLKp6C1MCZIrlfragSEO5rpo0cp+gjc
KTRZXGTHmcHYDNTzdVgfF56epZ57rcOW4bUuPnCT/lZ669ltNuQuBUlOR2vKIu3x
gbV4wvAN+oeeq88bgdH++mRyrttsKqenVp+8+KZXp0x5tHFkQl70xbysjZEtMu1N
6JIwXXcVs7qfN15HukYlnjCJwZVBCj4ovMfnEaSrBVszVcWdopUtLXCTbmwtMtlB
+FkYzRaQzRRSWrXkyAzypVmHXlxElBUpEb9GEwapJj8HZkKkd5mZnDZv6ipr+Bou
E43+hAWgXlA+Vh1C+G56H7hOhR+jrJFYfJBzXgJhu2YzZsYajWsJJWcZT1tQidjH
KpCLTWNh66DOEqGas8kJNZ2YZHcMu72qweBTFbs/11j6nYKvRPvQikvgTSRAk4E4
o5/6hepGQqVHnhO2h/qGo8XYVEzjIr6/Wr0NAuas8gJamesNeSJcbIcu/0/fE+v2
E0lTRusL1L/fPsTSV+lxNviTAum+V8eYXg1g2McQK5GWJpyuj9dLlMeYc2/81poS
xdTZWbmsNV9YOoi5A5gbqpC7EC4BQFPYY59O1o7sS4dnedO1ENTrlt2EuB1OS5Dm
Xe9f6lCVhu3ZCZVtw/pMQ6gQyqPlbOdfU9FVxuzF7DN8FZCKLEC26U7y810M8RJC
yFszOBjpxCf9fQxu6xrmsCYrYkLtCIsm2Vw7EWTXBaYiQiJkz168vHUSTObTqTot
rTFIgIHphdioqNPAjvAZJYM4I+YQ19bfwfa7tBRiPPV6Yd9E6IQrsLzWR9Z25XFj
w1GOgxLvBjN6NeCFNC6g2E7p8jM0SpOonqUjVlV01Z+48RmrPRIVQK/ZvqrTPpr7
WPYNZ++HzUDla7e3Mht5jo82byc8WGQmnYH83qY6VGp//ExtCYTnoI6T4KMrdzpj
nRSxxH5eaQCdWbnUSwwxkEGflrv+732CgfuJSLgYnhb5FOWO7aguhzpuq/Y11hrd
OLkcEK/ux7PGQkYtUpikQq9FRlwhXwpj7fzgBv8YgkIGa076HmLJbokHrRMMN5ZJ
P1vafb/5uYxxWo7ccV2OTQkSZUGKVyDSQRDYzwYKi7zBZd+zMqDva/CnLJ1Q7YvU
nZdY3t0bRu+h6RGytt0Ox+6MKWt3JDUkRsqE4krDM48WV5uHRWkVs3OxFoQdmQU2
yRkrlWlA5/gEcrFNFE8HOlVOkMLZp0BJGC7XHQVlWqSU6ZtS+vMtXFi/rL3o3Vmx
BBf11gszyLC5aTiC4lw9yYsp8bx1LQKDN+L+yAxhqcGHoduZHx6Ql0V0YcS+7r5Y
QJQ9MeJIg6ytzXZEzQ1SZcWKg35/26Qc7V5vUvP/FJCu6p0oB5BT8OEApcyyP9O6
NcDWTr9kOVxkE9QQBnde8gP6Ccp+EdYYuY0krtUbe08f2Fh/2315iGT2WN+cc9MV
PA8vZ7+A74PrD9Tx/ZU4iRf/yak6c5jpCfVpRl6K9CJKNnXKwAzZVUNzT1vl+iP6
v7Yp0Ka2NeDf5H/rUW4qziRjMVBZMnb3KX43bZfpD96IpdISGt3C68SNSY7lm43J
PFP5wK5TcG5d8vpZ9LcZKS+GPAiww6aPHZnhZzLgzAbaNdhQBk6doQwtDR3LagUk
KjBIwoPkD4crq8LqTd26XuUgqHYExarfmnlKp0lCNK7CoJTZK3WT1NWJ7m4HAvCD
YmcrRNkAM4ZzUGAIYU5IxxUQ3ajfrOYcVex9US47AWn8MD5rEpy9QKCinh/Jjpkv
3CmPIb2uqH+6BpFcxBjiMNsLRazhj0cmVL7n0WZc0A5BqOSpyF4aUDoilW5zOgOO
sVgiI9cWDhONAKnIVMjHWpT85UY0CFtRvSh3R6qFC+qeidVSsNXjPKoVLURyFDcU
ppI0mC3pqmDxNY8Z4Q8ZdmmJhI8VhfjYqSa8y1jabIfTIGIuZJZ7aMmw8Sp1jGIJ
w0QU5cVpz6zcO9sqpzIU5YFMc+H7GBHNm+IgiF8KvOOsNM+ZNCD7VvPcfms2tgbd
Ak7QCYRrgmtw8UkryaH+GLdErCB3F+GrA3zVBe5uoSZkJttOdPRvpzWa7sFIl/xz
QGre8Q6c/qepJwnh/dE1yZOzUBtEK+4bc2/VorabwBlRi/xHySe5nL+KlnGFVIXB
wrBe3fpKYrpOJ5caOh1m++8cp8xy9D80uQDgGs/4NsrJX+gh5QEKOWpABrYMQUMC
xzPq/PqYetX34WSdbNeG+r0RlPzCcUKu43XBm5z21vz1IlsFJjq52QJskAGcUDBr
iYQgisys012pGLV7up94/BsG0YZs733KlE5Nwsqa/wOoy9s/AzzxOwnT4t+A45QY
hwXYI/wRRfJ/OISu713kwJ6dp1t8VaShFCBpKqzluVX1/eLU23bQ6ur7J983Oug5
DYH11qzSqPlKigF0iCraIL2aaBYeviaVrawCNBuciCCOaH4RRgk3pwYDQUDBkida
sP9EV6QwaJrcYu1PQnYiKt1mk0iYgwfCB8Egp/Lrc/zvkyAS7+jFRNMBlw3DgDaw
GvO3T1OHRfQi+CsA8c+RKwp86Fwp33Yo3r3fWHlbhVyvdQ8+DmDvKI3LlXO67D1h
0FXvRIQiWREr7laq4u2pIbyftAlSoLgh0xQlNlmUd/1mgTIL+0pF8Zfe6EqykBGa
/zTEGYkrFsryI7uFdV2eV67o9hc8Iupm966Ru+F40iogrCxH8oi+5GqNnYOqPLY+
MabxuShw3M+u0QKcZcAYpDvGJfsc/Y2rkXwR66rMIgSuNBy2ofLCUQ8mTmCUGiLR
0r0bQ1MgLbI9OGd2siinchPlXN33XaJqS0R6KCd4W7sXTzKvh0XZ5I0pZRiPjuIx
S6m4j91Vxbc57JG81KQSOGdLMGFJ6v1Y8sF/EF/FNj/i07S4SWPgXS1TRPT3dedj
E1VRMAf2XzdIPwqph+bDmIlqjSBNjVK/FmM/TRYX4rWjWI3WaQqV1+oajSHQzAuW
2YmBqVECXTm2ck+IfUO57kxhJ+uLSJ8qWpG4s5gkjoHa1aJReJaMF8npuOa4xNpp
RImfp6qcENRJwVdl6gTmSNZWR2hbBBTF2GWAHWX4bWpZ0Pl7Z07cBDLg9w3xF+A0
VYqFSSV9VJvBPntFtTBCgLMPgJip2UtcVpBmnlnjSZz+rxHek6X9CzEGu43CBPfd
X5MZAo01OV0VYZOc3GVyPoFr7d7K08MA7hWqtgG1TvnXvyn7WSR8SY+fVxcM2AzF
Z7EL86NOwpD8bwnvF/bl8iUV13CnIjRq75gB0PyQu17CQQctqdMOK8EL1N23JI/J
jCP3Gucf0Pyx82M6vnJhQATpJ4cuHVWsDxinZuIWtKDLIJ/AMdRcCfXGelAS8w+6
3+N4jLHRtjeX61X+3V4NSy5Pt/jTmR+9wvbVdAJEIjdxsDYr5ISuAfdQPHeJgaPj
j8BkOydVtrwHJKEH//D3iOIaVDGO+7ZcUHvYBgn8Wfzn066M/dN766/kvbZcx9ne
RVKxTDrQb8LBgr3ErtmBI0RP8ArbiLOnywSVTI+wEFYvD/y2QuFBSuGHNKvyQEgu
7w4alk1ValtAgfMah6P5PfzAxyousMUARJHXys5QSa97PRDO7fi1mkeZ63z2C1RS
zkaSayyBm9wSChi2SM1VnS5G+7KecxMKytc+C8RAtnQEiDY7Op3WEjLyI6tHE8QS
9PpYje6G3SUBlbEmsPsRqqeWjAUomLQAsYqDFAUtC1jIzfIhn2ojrGYa0qkNuXO6
S1cVENfEqpyIAnNn39xmhJ5eK0exJJWkHTDi/kW0Ak0piyy8PU4/ZCD00FPdB6Fe
usmu+a18g5u17HnG8TnBVKqjPeGoX8VNwje5tNSxs0YaakgYtJmrqvnEUL0IlGTZ
c5RvF2LYEv7FpoBf0XddYQowB5A7Y1Kz/37JypIqNNBjdp0kEy97Ib+D1t8RYpSZ
PBGuissCg8oLT67QpQMaajAkV3nHlG+Yzo8hSysrLQrS0VHVLMYIB19UCXoOqCVK
U4XxsKUUhLVNUo+xoCFsT7OmoqCSI1gl3FnbfoCaICe41emIRGVcgqMCBKnU/D8+
qSMdigCPNVlkcn9K+ghYQm6RYezV7K/F+seyNWBNMqd10XOmviVAnM4vx5b76kff
uWvpFFQ21k/9LI4yQ4ULXT3J7bJZrIDNcCXC2IH4d/f9AczUssZ6e1ZfDESicVhN
+TAhfjO1TvP/G2caev1fQFpjJatp3ipARn4RD7mrto8h5nAWZGbbh9MQ985gYxhQ
dTsekjddJBZq0lMFI1Hg2LHmsvd/ZDb1HYs4bg8izW5CtMSE+nT/3TDrWIH/I5eU
S7eriztcwymoYjEwdYrUcTzkUeN/W1c0PoqiNYWjYqGUTm6wleKgdHZ5Afs2qDVi
ju/gq+PaeHkbgBpAWegOwL/N45cMKk+Vk2RiD/01s1tk8Jbbe5RoOx+cjPBcx1F4
BmwT4d22rDZb+SDQPZtu1dykyKCEUtkothjN4wnYuLSv2PSvvc8XJdx2BOonLe9/
D9Kf2ZRo5sBPVBuPp2F8FPLiVOzXjfrpXfOpe5yA7iHNgTL9sfvGrB/x+utPrAjQ
mUzC0Hm+t0g+6KfklNa/PYdGX1iljEGryWuao31GF94GoAODldIt52hQTKAY6XuT
sVzrjNspHE7Y2MPiP1wF1qQlbpyS3WhxRySH7ENqv1TyUB+RpthrebRlOyirZKXp
TYbIq66/mFfOUc2FsUObTlq+ypg2kryIIF4Ibsg1qs5+siY6RZ8jYNZYy5JHePHC
ULIiTJPKFGkUqM7gaiKX/ALqmhMZt8NUH4jW4U0OOVL2rU/lzFhFiwxjDBVFuMXX
vitVsPszrABCz0xRO11uVR14/8UZ49m2hRJPCvecC5vlK530PWehHsKIDHPWtZRJ
qrrPnEsuBKwFzQlqCWxrjuZgwjvr1ciqE+onr4s9BdJpQCSBSQpUdtXxJo6uYGri
cJvbC+kDpHK0B6Nob96cjfA5ReUTnbyhW/X7Ip2iaiMG/DZb35x3cdC6++BA7dbZ
2REylBU1rEWN6xW12PW8piUuk3xTYne+sNlFSSU3x179o8PwWbCAMvVBxc/wwAz2
BAyCax+O9GsPVEc/jt/JlHdn295afliC8/nQKfzZ/K6dzdgbw2td9pD6Isdcn/nf
uiRmeXqQEKoGiOmZzmlM7p75I5+lH4K3BIeryFfS4T4iLjt40wjN59T3kfU/nBUL
ycXFh4Cf2i2YqONOAcHjkBTvkkZbJwESgCybm9OlhLfU2Z/Cwq/h3l7VxLlrnO7D
EwMbDRkMdkTjRf5qDfr3LjVpWMhfh5zCBeCdXGgHSVveK7jwck6W/4e9AYbFud+l
bEzv8/iSrSA2diXz2ulM4BdekD1x5MQ/ojkAyF9q12ZmQ1efkKFc8iMhY1Fo9kn3
iAPYfbSo2wLt7F4ampcVhzBOPftRt6arZKZu2Al59QG2X8ZSiM1Gse/H8qpBXBaa
9CiM1Qw+s70FPJvZSQo4n0+u1cGKRHQJZDjx50sFzAIejy6MKZ63ftB7Jwhw+V33
1EywN//VR9zzRuiFjM0Ok0stfCkkWUsAhIg6xqshLk6P8XDueOcxF4rH5jgQBx80
dHzTi1jdLwXP2nDNZjhRgstEW3rbYamJYiiJ5ciig/2jbAtv2kyb5fZFHngKpRV6
EYtwziH10rnPVptb7jU2VNcSRlHxkpw897law6nS+bIsNpVNlyQFX+l684B3g2Hq
UaIerRtyExbWR81+xdak4Zh2Ih+KjG2N/hdifFW4gbkU3kCKWnaASDGrkIIjMwhI
ItLQyPouKJyPJUUTEuT2XUEmM61X1wEA6DrQmCeXL2yhhptOx22mKJj37zZo9ZjF
wY2DTVGWANeZNKHqPg3TUURx91nozsqIIJt78DDm6/9EIy8W0eBLWmvu4hlvIgz1
ruO1g1I/xnIFSPuywajXeg8mOnNJziGisKomEgpdKkLYbe1WW+W5dt0M9jh2B3Yd
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VfNZrnqXvndUJljhvlZw3bFX12eOdEI+JzFROjYbStADOkKM7Ex8onbllP1Ozgm/
+FokPLQJgQdoXG/wVsNBUjuQi4wqUn3Qhv6w6O+6WgRH1Uz5giOVU+EWPGElu8tv
oICtDNhXHtJCVytt3CVhPZw9YFvf5A05Dg7HlUx+P4TwOS95wOvoncCjCUJfP9RG
NyH0MBkA66XCpAy55GpOM4EFvuSgIhFOVdNSzLNohw1Ugc6GDf3FxJX2ZymQHiA2
ylA9EYYf6yk7jgSZdOxz0JZM1IYQv7dV9AQsMlqokPoCRVZv84/9V6hG4UUXJIIc
XijDkzgZLcDiN99pkYgR3A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2672 )
`pragma protect data_block
YroV+MO6cIIy5njZS2T8zctWBTUWPY6/JFwsnKwGDLJ6bb5PHhlSucQWZNDFkDa5
L1So3smniA7ALoXiHKYceiauaFnlJhNS7PrM7uousjAEoATqHFW2DqHjvSDQoAe/
YMxh3Dk8r7MxRMr/5hCSBN1hRD8X2zGTqVzTdbEkBY8K8lSeO7yHci69IphpIlEd
M3It+S0IUdBcMG+KQNzVrxix0vf0V+GkFu0FoNf+hL9M92siHiUg8eyE9qd+OdXc
3mW/an7431QP1LG6jumNjXGtz0jYmUurw4gnVIoJy95VJYK2vSmsiS7LuGq35Vus
kobBLcmrGy2EHnZbAfHfglw1kwfxUlzHWvER8LFi9oBKaMPJEvQIBIOPlO5BwjrS
da0ngJh7eR4tHlJ2A5dKz/uWt543riHfV/SCEFeV0p3Yt4dd/T35pNPFbWbf344k
f/Lt8f0PNyDPtSy8ZuxLQOYBKEZic7gny5VtenEKGTZItNJF1DTL8LryOdORqyU6
ICAO/vHoGMX8Ts3QLh6UatQgooKv7zO0U11fJuQ57bGF9pE3Kg9D61YiJQrlW9BH
pxliGbjh6h40ZNFYsPtKOtKIH0OXwFOAqb0FGInTnxkO/PfbxBSTxyWfEJOvSi8L
sNIin+5Fnm9nqBdwPy4ve22bxOI55v4eWdiG05ou4rQ+6XRTMrkSVGTXIMvhoJ6j
Co4MNp9uXZujEj7L/aYiBn0VMRD0CwKW9vLRsbyBp+B35pERXeGnuCwHzOIKpuoJ
zgCOeDFQnJwCtFyd11o9GCfshjKyCywm/mK5aIGt4sQTFZ8nTBWmifjfDvPKRswl
fZnuhK+wHDu/F8NdfE7fL9LYVjPX9tGsmNS4L/W4/ZAf+YiW+RgkodlQsgZCjyc3
Cyo0VkaqXlNVTmaiO83DGQfMwE9gXQaBQlYl4IwztoCuJ+s7TctSgju7hv/2BjBf
XldaXzi1bHilSqeXwirifuUvWcqJO/NiuHcTjUAnmQImtrYPJeZ9XzbYidUYX4qL
bxj/NAtFeKNBb9aYrH2tRV2bGmYTheNMW53E2GdZ+UdKG7Vd4vdn/Nvzdtar7K5R
1QpxiKxqBRmP0NAdqfL97AkNWzmnSUrCr3UoKQnc1p6/Ja6AdSmerbLafGTyuTiW
5ja7EnCKwciaKlaFwjfY4Hpi10Mno050hlJnxetyE180JNy4qrcfYXo29iKknopI
DCDpwOiDyNyahqMe6wUmSX6mnSAZy3DtAX5bAtAv6eMYEhIY6n6SrvxCs38UnHrl
L7e4ruEJoPFuNvYc1ECE7zjWz+wmI5aZmidieOcGikYb5xwk1aNrdhcHu2bJxDSh
MKJ2HpFeenrbaGoagscSwyt6TfAR5XfoEsUo/2Hgh3b0917cgu1tLFCujWDRdNdu
DraftSnehFooPEBOdPo5pcYGD5L7WaDIoPqiZ/WLeAPNF4UqZtUDilkehyMH7W0O
+G2Nb9Ng0vwD5X49wFq6R8lgxsOTAkNso6W+GWEZHAy2F6e0BVvP1L/8rx7YrIxl
/nD44ZoHCBurVxYnikQSdPkrfVIjlLFgb/DlrJ3WFauZ2zFFKhmHCzFCKeJKAsjN
gy5BT10HrZ5fL8Q7diZ35eq1ufZfBq3tfUffXXH/+XD/j/Sxvx2srH3FV18HSxSU
Rny5KDNk6/v/C/fLEXCOOl7cuwqgqxsJRBRDGBOc+5Ygt2rlf8YID0YM8XzlfQnP
z9iR/tsCRwujRDuoexC7bDdpt3TPtM+uYBVrmAMenzPgAASQ7obKTSFnfRbl/xZs
fcgne3NKeaNhOEdkIiv2udhGUHzEN38rs1uLQ6fqcH+/HivCRRzh0NLZdd2PbtLp
cwHd5rtKsFdUyjv+PPUlg7YvPJ0G+aWJcqUMFNYWCcmrWhk98z1Hm0tsFkAwQFl4
pjfu0sgGu5HkTHmEAowOx75Bn8uilxDuHmFMxzwcMn7uWbUtiPyLETLtOCJCQh1v
P/XmUQLCoswiYofrdoWwM+QNMMFg8f5uBic1XyR5zWSaHygF+Bqj2Nkt1BzaFcK2
EeaKm2Jc9vQMWX522p/+4s5VZz/uRpnK+PSUWnw6NXQ0q3zaYuOtqAgwfJ66wkCZ
/cLOzaF63lhdJaDmpzZYV9dRBzMJwfuLNdZGHibvsvsMJSZphrAZAwLYVyAdtjsB
lGVStN0Ys4ucQ4g+/TteyeoYBowzK3YRj5xdMfMlma35EHUK/D8pvB4esY2kk/Pt
Ku/DTZoKUUu27q026Wfau3Hp6qxggGZuHSIGlZB98rmi6zO72M0bhAdHpbQWYOx3
dkAihZnVFLRBfA8X98QQgb/9F5wzpT9xhaUrZMc/5EDswLa2VY52fTtFGG+Wzn0Q
oCSp6Ms+eLzkhqDsbiyTsWNMYavEz3Nf7B9HV3SGk9Z7YCVnqXo0nmbL4zvtE4PF
H4R1tR+ZmMGkVzV4uuASqBNEgFDQGRvkY+80nT967RTO+OmOcwgicFEYYkC2NUwT
m41QxkCErXNEAMhNPGL9fK6oxR+MAwhhN5ekKL0ZflgKiRnJRxSNWBfmpeTNX3+E
3nY/o0B7GXsIxxerXc/Tax2izcFonoQWJvp+E/9qAU8NDiaxlO/xi0ZHIqer13K6
RpZFlrF90A3ythaKvIoH+eg6FECnxvEsf7RHrCPdV9KNjKc9eNQEKLpl96TtZoBb
jvCGEZ8Qmqc9BBM9yv4/I7+x6xoivesQsPNwnbOBtk7lHCgHLItCeamDhs1a0EDA
LFGt6KCZqzhaypF4osFtPIExQplLXxJJJFUAHE0c5jtXxGPdM9mZJB2H1amG1fnT
XIYdQzioB6DPTRnY2LgrRbhTsrlVNyrQnU752KaScXdhNxtHFrcf9ZvsDvip8llF
ucY04ntT7OAhOrenNTfTOkSmqAfMUpTak7U83F0NnePMXfqZbB5u3DwQxveGr6r3
GrDK4RX6te2E+0ZnPZxTXnHWc/yXHwGfNEfnjI4a7PpbwJ+OqStHmUCkPraQ+XyU
4mFCKN3n/xr2iGHlnZU3qlAFtwyX+f6v8EiODP/wlvmbmvXy2pqtUv9EqbzTNh0R
q4WgUo+talkXsfzUXYniSjGez4pwNGFxr57UWAAEuRiHEZoyavd1Xu8hFjxcVZ09
XHBG17ucl4t9awlReVqGC2BtIKOM3tIIaPW3ng8PoGwyYEXPMnp2GU8apGiYb5Rj
uRk8kpiQhqYNnCWs9jcHAGNY+Km4vvPKXcZB6Xadr2m7gdCKTEG6V2Xa1Us4+1oU
JzoBJdx4JVA73/vhFYNOXUyXYN4sLGxbOoKeAtTZbj5m5ZMOA0J/zgUk4VlWYDod
6OazTP9VFSn1uIhWbDpBtR29OWLr54wZW+ALKWpuiUqdvCJRPiiSqf1KHWULMKY6
j1NuuIjvp5eyTmDvPYAOiC3rSx0f6K0logaPVS8p1RZemPAFR1OoJ3pqyP9Y1VhD
IWs6c1b8KVk0KmbipxPO168D3l0RAQejxmaGasooXMpR/p2ZSoXXVsFvkdRtT01O
QWtMSI1PBKo8RkC4YVuO4A+zp+Y7sOBztKX9PyAaIOg=
`pragma protect end_protected

//pragma protect end
