//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2025 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = tinyml_accelerator
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Thu Apr  3 12:54:15 2025
// ***************************************************************************************

`timescale 1 ns / 1 ns
`define TINYML_UUID 160'h73c81d25824e2a411de1366acd73e551dfbe85f3
`define IP_UUID _73c81d25824e2a411de1366acd73e551dfbe85f3
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)

`include "tinyml_core0_define.v"

module tinyml_accelerator #(
    parameter                       AXI_DW                          = `TML_C0_AXI_DW,
    parameter                       OP_CNT                          = 6,
    parameter                       ADD_MODE                        = `TML_C0_ADD_MODE,          
    parameter                       MIN_MAX_MODE                    = `TML_C0_MIN_MAX_MODE,      
    parameter                       MUL_MODE                        = `TML_C0_MUL_MODE,         
    parameter                       FC_MODE                         = `TML_C0_FC_MODE,           
    parameter                       LR_MODE                         = `TML_C0_LR_MODE,           
    parameter                       TINYML_CACHE                    = `TML_C0_TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `TML_C0_CACHE_DEPTH,
    parameter                       CONV_DEPTHW_MODE                = `TML_C0_CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `TML_C0_CONV_DEPTHW_LITE_PARALLEL,
    parameter                       CONV_DEPTHW_LITE_AW             = `TML_C0_CONV_DEPTHW_LITE_AW,
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `TML_C0_CONV_DEPTHW_STD_IN_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `TML_C0_CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `TML_C0_CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `TML_C0_CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `TML_C0_CONV_DEPTHW_STD_CNT_DTH,
    parameter                       FC_MAX_IN_NODE                  = `TML_C0_FC_MAX_IN_NODE,
    parameter                       FC_MAX_OUT_NODE                 = `TML_C0_FC_MAX_OUT_NODE,
    parameter                       ENABLED_ACCELERATOR_CHANNEL     = 4'b0001 
)
(
//Global Signals
input                           clk,
input                           rstn,
//Custom Instruction
//--Command Interface
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
//--Response Interface
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
//DMA Master AXI4 Bus Interface
input                           m_axi_clk,
input                           m_axi_rstn,
//DMA Master AXI4 Write Bus Interface
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
//DMA Master AXI4 Read Bus Interface
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);

`IP_MODULE_NAME(tinyml_accelerator_int) #(
    .AXI_DW                          (AXI_DW),
    .OP_CNT                          (OP_CNT),
    .ADD_MODE                        (ADD_MODE),
    .MIN_MAX_MODE                    (MIN_MAX_MODE),
    .MUL_MODE                        (MUL_MODE),
    .FC_MODE                         (FC_MODE),
    .LR_MODE                         (LR_MODE),
    .TINYML_CACHE                    (TINYML_CACHE),
    .CACHE_DEPTH                     (CACHE_DEPTH),
    .CONV_DEPTHW_MODE                (CONV_DEPTHW_MODE),
    .CONV_DEPTHW_LITE_PARALLEL       (CONV_DEPTHW_LITE_PARALLEL),
    .CONV_DEPTHW_LITE_AW             (CONV_DEPTHW_LITE_AW),
    .CONV_DEPTHW_STD_IN_PARALLEL     (CONV_DEPTHW_STD_IN_PARALLEL),
    .CONV_DEPTHW_STD_OUT_PARALLEL    (CONV_DEPTHW_STD_OUT_PARALLEL),
    .CONV_DEPTHW_STD_OUT_CH_FIFO_A   (CONV_DEPTHW_STD_OUT_CH_FIFO_A),
    .CONV_DEPTHW_STD_FILTER_FIFO_A   (CONV_DEPTHW_STD_FILTER_FIFO_A),
    .CONV_DEPTHW_STD_CNT_DTH         (CONV_DEPTHW_STD_CNT_DTH),
    .FC_MAX_IN_NODE                  (FC_MAX_IN_NODE),
    .FC_MAX_OUT_NODE                 (FC_MAX_OUT_NODE),
    .ENABLED_ACCELERATOR_CHANNEL     (ENABLED_ACCELERATOR_CHANNEL)
) u_tinyml_accelerator_int (
    .clk(clk),
    .rstn(rstn),
    .cmd_valid(cmd_valid),
    .cmd_function_id(cmd_function_id),
    .cmd_inputs_0(cmd_inputs_0),
    .cmd_inputs_1(cmd_inputs_1),
    .cmd_ready(cmd_ready),
    .cmd_int(cmd_int),
    .rsp_valid(rsp_valid),
    .rsp_outputs_0(rsp_outputs_0),
    .rsp_ready(rsp_ready),
    .m_axi_clk(m_axi_clk),
    .m_axi_rstn(m_axi_rstn),
    .m_axi_awvalid(m_axi_awvalid),
    .m_axi_awaddr(m_axi_awaddr),
    .m_axi_awlen(m_axi_awlen),
    .m_axi_awsize(m_axi_awsize),
    .m_axi_awburst(m_axi_awburst),
    .m_axi_awprot(m_axi_awprot),
    .m_axi_awlock(m_axi_awlock),
    .m_axi_awcache(m_axi_awcache),
    .m_axi_awready(m_axi_awready),
    .m_axi_wdata(m_axi_wdata),
    .m_axi_wstrb(m_axi_wstrb),
    .m_axi_wlast(m_axi_wlast),
    .m_axi_wvalid(m_axi_wvalid),
    .m_axi_wready(m_axi_wready),
    .m_axi_bresp(m_axi_bresp),
    .m_axi_bvalid(m_axi_bvalid),
    .m_axi_bready(m_axi_bready),
    .m_axi_arvalid(m_axi_arvalid),
    .m_axi_araddr(m_axi_araddr),
    .m_axi_arlen(m_axi_arlen),
    .m_axi_arsize(m_axi_arsize),
    .m_axi_arburst(m_axi_arburst),
    .m_axi_arprot(m_axi_arprot),
    .m_axi_arlock(m_axi_arlock),
    .m_axi_arcache(m_axi_arcache),
    .m_axi_arready(m_axi_arready),
    .m_axi_rvalid(m_axi_rvalid),
    .m_axi_rdata(m_axi_rdata),
    .m_axi_rlast(m_axi_rlast),
    .m_axi_rresp(m_axi_rresp),
    .m_axi_rready(m_axi_rready)
);

endmodule


`include "tinyml_core0_define.v"
`timescale 1 ns / 1 ns
module `IP_MODULE_NAME(tinyml_accelerator_int)#(
    parameter                       AXI_DW                          = `TML_C0_AXI_DW,
    parameter                       OP_CNT                          = 6,
    parameter                       ADD_MODE                        = `TML_C0_ADD_MODE,          
    parameter                       MIN_MAX_MODE                    = `TML_C0_MIN_MAX_MODE,      
    parameter                       MUL_MODE                        = `TML_C0_MUL_MODE,         
    parameter                       FC_MODE                         = `TML_C0_FC_MODE,           
    parameter                       LR_MODE                         = `TML_C0_LR_MODE,           
    parameter                       TINYML_CACHE                    = `TML_C0_TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `TML_C0_CACHE_DEPTH,
    parameter                       CONV_DEPTHW_MODE                = `TML_C0_CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `TML_C0_CONV_DEPTHW_LITE_PARALLEL,
    parameter                       CONV_DEPTHW_LITE_AW             = `TML_C0_CONV_DEPTHW_LITE_AW,
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `TML_C0_CONV_DEPTHW_STD_IN_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `TML_C0_CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `TML_C0_CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `TML_C0_CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `TML_C0_CONV_DEPTHW_STD_CNT_DTH,
    parameter                       FC_MAX_IN_NODE                  = `TML_C0_FC_MAX_IN_NODE,
    parameter                       FC_MAX_OUT_NODE                 = `TML_C0_FC_MAX_OUT_NODE,
    parameter                       ENABLED_ACCELERATOR_CHANNEL     = 4'b0001
)
(
input                           clk,
input                           rstn,
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
input                           m_axi_clk,
input                           m_axi_rstn,
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
g4/q8kVSkvJFPnMyLNYzdJ1Ra1kTUNRLGs2VwwOqpKSH28/KCjNfel8sWP/Hi6zF
fyGtm6U4qDEz8Ob2zRQ5wnVAdyjSIfFnTa/N8tU/ndFTu++IG5wf+jxkxNP6ttOO
N6zqHNnNj+NVRGbm/FQtj7ejrVq32JB9rWXuwtqMkoFK2GdA0vigWyvYv9tAiYcn
6tNcup9xit8Og2mIoICmJ7VbNOoVDI6F++riMrkqBT7jQ8T40gpwV5poR4Z2YZHS
mu7VJo6wYvGDWIp07Ca9hDyDqE4tt4Sal5iFGJWNPS7wqjyC/vG8Ckp+YKOC8QhQ
OGN1RbhPfnGTyzpaWnckXg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 61232 )
`pragma protect data_block
F+UjVXH52tnJ4HZnfZ26/BiLOk8NwG5GH/pwmTcAVNHPXBPpX8pSsCk11qGY9Gl9
lCIa9sCOOAH64IZfLYSy87fIOtdZHi6p0el9MGbIF2o3kdY9TVkgeDZHivul9fu2
TyAWhqswwcWT0lkXHPb6g/fAhbZe+tnK9/yHoWXpmCp8+yu59KURn/YjUAmDi65N
fgKYRNNBLXwaemhdxhuqI6tsm6V24Cq/1kXm1HCQ6Q0RFFJOV5svDJrMsU934UZK
4NwbU897qYS3+dc1C+tLgvU64MOZP5PKA3DJ2k7JgdJm9cd7xtsQsnwC/oyFajSG
/D4BoA8P+0ye1zsGXSG8um1RHaUD173td4+p5++XxHb8xPaVLPXNtZ3SsTTaGnfa
QjO+9ih0Hb4znbwaDskwxJYEwyqLdb5oN5O0dU0ffErHgYQ7QRBaQHUMC7/FTeVp
bYmmklz/HX8q89hnwNC1JJMHb5fgAEjvOwdppTHNU/i5aehvCct8WNGYUs/BIHSx
YbDDmsECCgrJGqwW86NGfrvUvzsRPzDq+AVQBg1QPidamtQsKBSCVtq56kWIhTuI
u0Eumrbbn3ml9RQUT3NMtovyJvwcaPEyTl4dQe5Hc/1MVn2MAdcp3Hn2OIZhLXzk
y2fyv8ESnXSCd4U++kjHlKJYukv0iv3VubZrdr3k5xjd5Mw5EGTZeQDnaQTsxSXT
3ph+tqRJ/WTBWpySi67KsUYfgGn3ngPWAqPJ9tEZSYbea6/TI70+xOePTxMYM/WJ
rxHp3dZQycSUEX7IwFQDCOxURfXAuhy9+bZJ9HVaX/zI20pHz73g/7H8qHcWlWId
JDoM9DUjBTI4UgRX6Gmb/Y4wwZZYwmQcX/9tHyG2E7EzjKkmgfs4Y4Ul7HidKP2H
XaA1D4Anmy0rwm0Y2dxsXzm3+yDubv2QzUvMpqoVywCqBRsJNsnSWqeJJ8wr+EYX
4QszGCVFL9sIdOn/6vkqOzNYMlMGU8xQTx6pEtz7yIFhg4r68XRaLOP9wn8IKR1m
PoRARKzPIyrWbOmL5nNbqHW8GvZC0DQnfK3gk8p2NvnfG6o8oxBWzbybcDD8yKVt
i9b5S84Ds6S5mXP1ZS0YNx185li0d4F5mc3oZ7FY7usE6fOyw7d6RNLnW9dx37xo
1FW7yQujDDDhcXzuK7rd7PVXFmysuMCAgDnrKjN231Xi2NERVnASTkhXeSG+S+yr
YGpR5emw+fkiJ8YypPktPY1fhUvpPWJhYa//+ANqLphoGL26Kc3ZayNtN94emVJe
60GpuNFlF3jEgqG7QX69+IiIVona1l8Cz6r1FLdLDoYS7Zx2WPmYIPaROE6qejsU
4vB0Xmv7k9+UpJ12Y5JtFlKpXrzVPWV/bgUuio/hBtvDWQjAU/qgSNBhzZNc9znU
ujNITT+rfKJZfch0+gFneUsLeYo02TRzOriEbP7uMLEapRAyBiFrOK6nbtpDzYBt
ZTFm8cfZDW469gPzYVFw3Lq8H9bFiThssEhN6w8vRciTvHNHHZTjlCWHSnTIp0Ao
tnYp8QG4Mx+x0UD4ooSExEnSA20fHbmV7NbPbEL3mHWkn4VABjRchMUQArdOzOJB
cOt3ycAHrOqWoOBGATRYV0s9GoN5JtZRAa9OKxBnXBVX/HHrqh/Cv08iSSQJRGAv
FbSJ4ipnsEHc3XJwPbEH0MkBa3WmAjqZ6kb/OcpRinPgMsmcHc/owSkc8Ptti+Ix
W+XSz5NPJ1AiH5qIyFeagjejrBfbj4fhEwpmXzBHRaELCNHgRzwbRNw9IGDfWIUs
LONA2/XnDa2cPWmTbSV9ExTDaloVaaMAxH8rsl7SMTpejQTAa6Pv0WGGAdly3n0C
oNesXNPQtXywA5GTOs8XhWMZMO7Bacni7bX6zRHH9RXnvJC7lNa2p8kahY1WpG1Q
5e0PXy0aSun64kLJUoU3QLdapcNG8kVDR0KoZX5KJl8uqj8JHUQzbfoQiuU00/fm
x1J87kopvxY0q4w8fs5IgdBvfxOxQYsFvYeA2gkHx2cVAcw1Qz0b0Ha+6xrNZzEr
TOGsW+b8WPYQ7ZM3a6lmSpRz2y6ppyBg9mnm+yGBrVrqvuRjfYmh1Y/8o/Gtdi+p
sBsu9E59dlv/BP73vuOhcKkL4vqAXPiOHb21DFIMAtH2ZNMycgf6lPjSGXudSxDQ
V/FvrIb7q1x7/LD9HVxzqdOXV2kVbkhBUNcH+lr1EVx4l1Qtx5w+ZCshOIktjmbR
Sf8CAdBJqvFckrDZdESrN2TLqiFCPmTmWCR0MTORHC8I47sRJLNR+NICLJmwPw7Y
7p1M8J9EQJgUak5bohVPjSw6oENvypx7Oz0LO+x7y/hCyBqlCacE4EDIq1GBfn6E
+BuKD/IIm5jTDsRi6KlsqVvMi6y9K1r5l/vTWd1PU5VAJzhAcckIJaYQ9ESBWxFJ
AxnbTFZ70NYjfBRUocQBpIxJPNqQmHGdCPCfVqSlQPXCZVlLRWShmmUqmRXuJRVA
XKvjbfvqL/3PwKe0S3A5xnfbxMUEdxwmPwxAbwjrC5QUwL2uUz7hPgYKSbE31DlC
KdW4tEcbfbCo3O7r9aGftzFbZdxiLNQidMUM856WrTEG+gfxcHkCSwq5Q0HiMjNg
XZsHW2saa2GRR6xLoxgpf/70YKNwdkM2fLx3t7LFbCLDim21O5RH+f/FgxqAY7L0
g1QU1uQhB5D1PNa0GCrjra5fDi4F6xmLQxEdoHFUNZsjdNZL4lvcl7BAqXa0e1eL
VIYH9wRHphyuA1t/DXXgxGYq6tS8rEgDphfbNKezcrQpcg+vZUhNAsRyTznLneVP
r5pvZHzveXPEzcGHVK/asJsk5Ne4CmiIyBHWWKQZtjWT+rQwMAbxua+fA6EHDIL6
E+fk9UowZhuGOS8F72V4xvojL3mlfkSdJN002rjFqQhfftswA5TZtGAMdr3Md0ei
TQ5nmEn3bZ+U+rQhP8FbFTklB+gQafkxs8ND56/kCi1CVkxOdTPiU22/Lo6ICf1d
2ZM+X0OT0hjdtZ3mW54PJvXT+XRnmogMoDi6Aj0ac3SVS2/ZNZ5jljVse0sWlQMP
OrDdRbKxuXfVbApbsgfc9G6MrP3ISkMGFtWJr3bcs3l4Fl7XFsdUu1uV7FqIoYtw
QTvSX6iH0CTq8AAZ6WKgUobAcWq8zacqfvHBFFMzDlhVIh52T494+P0kge+VFrbq
jgZPvjVvPZ23Lae338wHkmDZ4iQdSZFW/M92gPKP37NqAeeFAjma4BnZ7xg+4v7x
s1lrNakfsyztSK+NKs95pIO7umFicSqUxpNjeO8Uvh6N9HKuSDNUKsK4VCf6ltZr
zJQpOoxX+xoty1XBxxeQ4L/1lLA8d4MbahzCLzuKOKZ/Beb8LyS+xPi2mO8qEQzr
XPaKEirCI+bbnu2kallCM+b/qMvhYrXhV1YWoaxnDJzoJbGL17ZfByaS5k4N0tEr
PzmtIdfbI3/5xgBlfo/E+wOTzyBFRkeNL7lLVMlRmmgqlFHrKxdcDXhAjw9aRdBC
N9KPZw6UFhKmuVwvy9dF5BTidFbK9rv4eXHekBQSkJ9C+UoxuRC2Y+B5Dm9PKwB5
7QPc0xtO9VUSK8EgFOnoStN7Kjle38XyRSjNcq8Xip03bV+jl1yY//er4zmrWC9B
cZFOTRzjnwquVB2SAjJ1Q2leALiedbbHCkrArQbVom+cvn7KatQY0ZXtTa4oxaN7
8ptAZAJXzAlxrA5tN5M/j346/DJRI2DDXRfvfxSIP1qP2H9AQBlYKAQtTVHdXLak
RP1XnukbUech/IDT/ULcOMG422EtU6XH5kzx+GDCqaiF2xwavWF5ftHHS1YEcO4x
E+d21jHig1JafMqSHHUkgsHV4xYhuvIEpK9velPbp7odDZrf6BwaQJvNSp8vkSBz
FagmZMTAEhXbZdYc5wGwGYzaoH6op4wKFoWpSnANKISoQBnlsj//mgdAIp9YOTH3
MEmiWP8TgZI/ACR3OJBqQEoWLVFzbXUNgtXAMu2NW1n7BSiLJb80US/7B/O/1z2V
RbqGCmzvoKeGV1eSdl9WaxyWg+guwv7Q1YQq6t2W8r0pIg81PTABsN4xTOTKNsSU
5secdkRql3HIhMLs3/Hi/2jyOtI4bxbvaNaZXSAgtH16Xvvxy3Dq/CGv+vIAQ/9F
dKLBFZjrBBT7KmofETFMdB+4fqc8D5a6PcVaxLa2mr5s5rZOKELUb6AWfmR2Oc44
Z9IEn92nq1hZmDKGAbecmh1QJjnOdnWM9nfJqGN8vPaYulnvzOlCiSS072hVEvAf
Oo1vyF3fzT3+Y93FTUcUHR84DcmfrFGUNx+blX2JIZGjEmyBSRRDOXsu9fEsdVd1
2IIudTRPODWIw2m/uiNXdxbfLVXNJnRYt1poEXPD67ROwlumSwgmeC1peEe/46Ts
Ib+whKvTEiSZNwOPt/AE6PruEai0GMWIxUt3uRBAsvJCCtyGaXWLDYrdGRVhSQQz
u3JporkDU8QejKCkIaFSNgOCRBkRhWUukb/KTu2VQgx0OxwEEiUqiltjTu+I4DDA
JK0K1bA2jX1lWEvqavg/uVZOSc4Q5Es4oBqwGwv0p3U5JD0JfQvxbN6Udcx7+IjM
UKQ3m2joHg+Nx0siTHvRjrQ/4g4HScaxqkZ2XTQOds9b7lm+8uIkVsOlCMnocOZe
BWDvvqCzASULkxtNSyG2e109f/0HdVy3GGOUgQDCq/y8NZ5j+KxxnTKxIdPKW/Pa
pxLPNoRNdEpM6urN1cTDwgFafUIC8mJlrP33jtuaLUNXN2y2fTcU6oAwpni3H/ii
5zABW2/H/M9MPfLya9oBpEcQVDje6WnwUMsPf5/YoTHTXyF07o10I4a3/qAyylkC
mNakygihmVym9SP3nNHtXUjGqGnd+0ntlWlMlPQYaFZDtphtBMWwVSUJX2qOwcYV
V7gchzDp7olrybBYbDqy0mso+OK9dOo6fikCbMh5RpCO/lQRioQ8JVYTlaF3bj3H
/CbaeECXAJWQ3trV1WB/7d7BFS0iCAopMwSuuVZiHIiJ4OrICUbYuYdlYaLFEqBy
zfa6A9MlCs/8uJEsTdlRw5YBmZEkiIqqKRfiiXbevcM1Cfyy9NVHQuVsFZhCMXkH
q/soK0Imosc8Al0dgCTMgDBMV+SnkuKebRRmwxu0FqBNkJiEuLbOFCXty1furNYA
pZC0NRfwrSSmyY3K8MXx/qTsgL0Y7Lvk0eQd6mwGEa57BM2YmBupQPUdMTTFTDpe
fYt26DMQlhTA4V5Ann/WWdXVJq1cws2D0i9kq7dGvROSvNFrX+jsicya2vX9JrKw
Ap4fyRwRJgcFkSf+a1bgXhBNl5MXR+paX0RFPt5QuetF1i5kmAtbv/aFRB+n/JMl
OFQveF23N1atssyCNn5oPcojRODEhw9cLq9oHaWSw5obY4RdIIGgzMQdfRcXoeZb
8B1ahUNDDyte2S1jHka0gWqs//0MQJyMOPRGZnOhDznA06tkY+jhyTgoPeqiivP1
PvuzyhJN6LyT20zDpVHQY/KdW9dtbh5AzvVWEGm0EG/i1LY8PZzkK3VmK9VJJbGz
+MgTtyA/1xeBrc314cDMVJkUsavaAwzOdbiq003KfuqgF9hQTAAC30rDvLpwWTXN
CQytJmxtmm4Cn+XBAZRQwCsgSirZRraS5ck+6Fr2if2x66kSGDemnAvRa8Qse/ly
NK7bYDxcU7B4X/EMdtyN7Nc/06brdrIMPSkOmCLvtWJAAjsFr3zjvXBASnqRFqXR
HVm+dQT4bZa9cIABOf8YyJOUhABc9m3Fte5Mu/5Gd4sG/KkGbp9+6CuQl0GM4/it
hQfv2ya9i2exJRWKNrYQLaNvU4Du9YsayalcOiPTDrxsE/j2PNWWDQGaQOS+ikxY
paFLfmFo+vChNKDduqTZgXOQJKSDUM5SRQIvU3lVzEdBf/7n8cQ30sqi3P9LzsOE
4NZVa5pKlnwGZMR56N4bWEu58yJarHK79uZGSWShaCA1Oi+U4Edob6zPmaepZN+n
iwmN1zP9Ye/UHsi1kYnVkSwb+DAiJgKdWu9YojKUkrFDEh13oy4dxXou2rSj5j7T
im0Z+WskMNkiZF6s79q6GsJhromEFGjLxFPg1lbxfxbGNvP5FebVRC5grllCMVOq
oIwmkkFuoOmXf4dctBf1iOYo/e89indDpTConXPtDgIv4GUp6q9zzQwl+lpOmRhB
V55o1uRPz3cNpF/2/McrtylwnDr1AuYAVbg8gRaHhpSynd6AxgmtYPO8xNo2/8uD
3shtZ6H+CGUh3MU7ywKVhEq6lwJJ/RmGtkubcR5zCDzyKBuhzQnBDevD9scZB1u9
9gtn0+jpoc2zfEU3NgnbrVTC+nYqhEx1VPYWNnqi+EP2BEGAeFKfkutHHR65ZPey
6ihDJBJAR5wm1QXpFCAE5VTVHDJCN+sPcwSj1gpWCvzMJHPNzlpAY/IkT0tnQfIL
JeYuyyV+id8E2o4AS/6gIbn5JiuqiCcJD/JiALDJATABzOjdPVWEpISmWKwRqGcw
Ekc/qM/pCx7EMsCAA6afh+Gl23Ga4YTYbgMLN87wIweyiy1PsKa/gOArtUAf0grM
TsmYWTG5IRmZtSX8q0MxZ6GoN3x0OdIcRjb0MEeLIj82wfgN6jJKuWV8QeCyg5rG
5vjJdJlU6UBg5iUZBMnRIftaUIK1TjzqFkmLE1isYNqvaKIyVrlWNxsl9gYkDv3X
bbI7LIzA7UAo+0uauwK5MSjifbj839ZqBbsxBgpKlSTw7EVuW7YMQ5eLhnRRTE4l
kZshyIlxey/ygZeoLVg3eZjqa33pRONb//nRlpsNgtwvJ2UMCeyjD2L3GOi4ur6N
5SFgFXk93HJTvxkD2rJGBGUNyjS0bYWjop1WdANZ0KllNZjbR/xokAFcs41RYOwB
SlI3odi4ALdR+DeIMiVj1i2GSODFymxrXW/L09pgM7ql281N1mocMEsun1/2pnNP
5MeDExD0WOL5jplZb0Cv7LWPa+PppHodtfAZMXHD2xTFmB88sMhcSrRaxTP9dWrg
3G1lMbfaZSDoB1fg0wQ2U2P1J3TkvlsSDhFR1M8Pn3TKsNa6wKUWg9sU378cdAaS
URsbrWJrMANfqfZMB1WPb9eAd9BB0NLbE5r6V2RNm/+048iwJC2iV1h7lF2gl3EQ
+OQOYWr+uGRhTC7D72eU796zKrAT3dOrdVm4LfbK5JOL/p3DeXtF4/yl9dZs9KDY
bpfRX0O8Po6uxl7PrmpsngZ8OUVHrVJKd/ew3ZTdEEakKFJrYqD9ock+QqQPOI0C
7pn+8OvW2UKPlq3mZYPt+G9g+eKS7xiAXCTdFKi1IoqB9qzKT+s87PhZE5sIRs77
kC6NJ96D3xWjIpQbNcJtrJtjIVYdyppye5ZDsITYFSUIzMFegPHEoMqn3fwXTzHY
TsRTXyh8G51MBGMNaBJxMQjIRJvcVXhki/N5PdxOGJ2Yj03vE+IA3LFsiOpEa0Jw
OPIgoXJyFdeMiKB0nSpNVH4sfV9aw7SP7R/9A3iBVSWy6AEAHa8jzaybvbTNOXbk
w7PV3tmLqYIxU2YfMwuX4mNe5h9+2gZMGo6UtPEXkRN4JN0VyOT1DzHpBVVnv8Cn
SwtZRtK9Iv1eHYKjf5vJIwf8/HH6eF9zzoYrOHxb+yTlPakj7PubekInWlNvg9sC
xO1KRUzbmrR84RlnToEOufE9wRIM5JvKRR1V/jZ55zSEPpsvMh/onBFoutrnEW/f
7gSP/OJKSWaDsUMtohitQ4gJ4tdBsVMSdbP27Srx1t589AKdYZgmxBYVHCQvVZZv
B5jnQO8pYcb+JR9MIXSFLfjDIa/y557vHH8gO1770h8WJNSS7vrZTqiVXcaxegg7
ZpIXVjiNWJPkUM6odRGyfeElR5TUfwWLJvAY5m63fcuKr1PRfIZqWlyFXQR0mDXK
dvvPpkKszO05r/3eASIwVgEtwV6TaMrrH6ziqvTGZHgUEzHU0F8V1pMfIz+vXick
Hl5fKZqwZQtOqJm/rQfZvYEQZa55N6OhHL5YrTEyO9OqpQQ4m9u0VMz3jK0OFgKf
0/T+9Mk8L7Hvh9FYT07lrWfwWpeGP2aFNuy83YnpSxEtiQIk1MfVXuleZtMk3fDA
MI6VJWDekh/UJcrQxG6aKWPgxGrwpTHbYDoBkPoi4/ZV6sh2Zf/JMcLPZZV2k3wT
yX06hpJZ0mFZNi59ZuSvxJmhP7Qp/EBzjxBCwQ1CLHJN1m5BCs5y24Zeb5/MlZAn
1VGp572k08ur5JeT3JLAYFvgyhM0UEQebw2oJVT4R9Oc3NFaZtc/dl8h+gebiZzb
y2Mzcpv7Qqy6IpfqeYq/mBvpbd36dO/gGhSYnUg0iKjhpbdSk6CUsWdd2xrwospq
JOB7e8il2NN4cb2+Dp5E6ThSjogGhxkAlWkroJZxgYHYUtW29f9VwIjLKBrsYN4t
Kb6fFdo5+hcTSlYzEVy0Naotci3xanIQ2hJyuEZn1UIgnRtFrKYW723AmOc4ZFgU
7bZJkZM4xJAdIBOWyTZS/3GeoUOPPLskCc7Fj6+Rj8xSKexXbocGmdFYvMDJUPOl
X3w748F0aC7K2k3Ofxwel/cPE5VBAhikZlWquXm09dEihYAJb2KnIO7MDBCT7Q79
ADdD64hw5WRyzTDRIqQyEfoKjoMmWT9fIUFr1LsMkhmTSk8IBMcJoKct9miY3qXk
nZWp4u8qnnMlcyh72rIT6TQ7X3cpBz59PA5ZGBN1V04dO4bRhTN24jKbRoYG+v/s
NkHTY+DvxK6ZfzTrQBrc2/DVBE7MvJgE6JB26zP/Z80/XEEDtFzwnbziQGGaK04W
bilWziZNN0ljML04nM1R9XJyoxWbfVR1TwT6R7KKKZJWaX/fWx8WK8L5vNpwerMA
d+BhPvL+lB5m8Z1zLuUcAXLzZyIERyUdvMkfEOE19NkmPbukITYYrOU/LbGr+S7C
hiQh2En42p52OczCDuUf5r0Yz46uDJ43mXE5M08CPgBYB5RDMbXc91o8yciv86hY
jQdhKF0w/qi3gcXsC8FinUbukQjcr9r3n9d/5npT6VM8EuvT0IODyTJGIKwMQUjD
yDwTzrU17QuOES7oh9KoRdOjCRNE8uYSsatwtzWe32l5EsxkxB3/MhwoS9vPf8HB
cUWsCUhXDLSJKkKL67l4CdAz+HumnJ1/pUcgMqiF3FHblIG61uV8prH64QjYC/R4
tHCAYUaris//xnFSyfc+UnRNXt9anV91R1k/dS3O+MbptyQB4xTimmEcJLu79VDf
5lAtSsFwJ9XRmzIU8A+oTF9MRHHMf/r+OolWZNyCSihXtJN45WCnd80LH+AmUV9F
rGcuff79ZESHnC/ft+OQXWSJEzm75VnBAdWPujUjSSGGq3vKbihKeNOjzz02y61F
nu0d6ktcEZoB8iKJSMU1KvKWfg5lg1vuSfGwwY5SAmLUaGo2tGsetBT8A6Oop70x
2PynEnk6qtTIhXIcZJiszWZbsY2QzqvF1y+JoMts22+yRFC9vFxDeUwKvkbki23p
L3+E7wAdyQnNW+0SCW3/4tpfrTq+CyilHBIy7f3U+k4R4zycSiyUu51IabbIuxkJ
9ieEbE3jJB3tmhG1VxbJp89vrKEU+TypoEJqF4Ki1/igRXVMzDKhX0VV8VZAyPzf
eAKeOXqg2DMRZWamRvAU9rki9QZlUXoYZFgfHunYQtfGZ3gccXDUbrsYNDPn14/0
rX64u9khh7SrutGxwZxXjkgGwsdwpqxOVMb7I4y76gUeuHHr5xQm+fwFdtPbm1br
icF4Lc2QcPIfzybpJBQMwSMCRbKBjuqkox23X93FkHAAnr1nOU3g+hm+VBlngeqT
zLBtLXufBmdFdR6xuITTs6EKAmipPb7qgR5aa/ZcC2PMJ3cmXzS03qWkmRQGX9hM
W9Dj+7AYP+iPlDIvaomdn4DQWLxcBffsU+gwBN6hJYYlPfxfZTRAFNpLXlwZqpTq
VDO0MYMec+T8nwJCnWXx9DXrRGEhGUTGig909cjK6gHr1BWaejp/mcjw96MZ/5+T
deR2zc+RwOH5/q6LrTQK781lO+eBBIUHPzp+v7/9MP/Kx98VNb+PJNfcPrG6vpLg
HFJuwbOs3TzyAaJapLEd13FTjQYhJZFiHb68sKRS+m8Sn+9Xsd7kgFJaJx9kdxQC
jGGUoPwES2/osyBQExpieXYe+xQxgICTVoQlTfzUkyc7G2TYA5jnAwTL0w3mjkTU
IH14h3SURfdmYFemZqXzv4gyU24u8+cktckb8FcvNnBRscSJTmAO6R8qPWGR7lB6
LGSIxMNNuDLYaO8cDwBfwh9PBiBVVMjnRqYQ7xk8tQjTRk3OEpPStSo4XTaqnWok
U7GzcacYy2fUrY++s+88HxR6dawGJSgkSUjQtQg5hDyLUKBme0yCIZWTUvOZaqPN
ohJwIxXiHuZjvx9x0gxvbkzFyN1H4CoJmR4x0DSGk1MkyT46KVP0+VHMInzuPgCv
oF9qMVAoGt8JaOGahxZh0bHc+NCc7RotJfBBfCkCtpmYaYRaUg4lWOkMyeb8237o
i3rW2aTLARcdy51ZjASsJpaxjhtqm+RUHgHHAMgWnugqNSowQFMU6NVCDPZvhDp/
/70cnUTBzw8JJ9AIWGN/o01OImrI9oVjw8OGXEBFZJ08qlTZQJlL9hIqDe3HHj/V
kwHwNgpumRtBpAcOUjsm54CTn9aJ1HAz19AvYkhUgB11aF0oHHS7ZYUXgnhyyrd0
n/WoO+Og0ZEkm0/T1qvPfZkQ4zAT+dvLhBVvkPcJIKT7GQG17WqDtv6cF2k0KG8v
WtzssiNsOxmkpw6TqGfUp9oeSO7cWxGGgGngi/AwKKZnuo5pQ7bUh7kYqPJapjN9
qfN+a7GvEnw6RPO8dJDpOzr/ixVnN4imrXPVnTLmQsZLtC8B+Gz9uf/ir5k3gC7p
pvGgjTBhER/I5QF0g3tjw8D1p9VmEgxgxMFArFRDIdN3CD1C+guJGaCkzpA8X5IU
irtbipko3eQWoEuuxCfZlpsmDxfyV+UronqGLX0BUley7RIoTCoB6aDJbMBGSpOw
8ZQ1dcYestQr7GsRIT9bC00sX/Tyj+RhGMIGvX+z1rqoZRPPFxSz0qxEYncrdfUq
D6KwjNJCIsiUeryj7dSul5h2qK/zDXiKInI+f2KYHPlL3AM5LlCNLeDHc4uGa6Yy
VlTc2OIsF7xDDx1IQyWOvihSrPxJc3EPodpVK7c8LO27AkxGOOYRDN9KcFF4Dyuz
O2z9O1L9++YODXPYjGIjCRnJBLgLrDHr8r5Anl1Ja2yKNzDO9UPawmIEEnMXwF3+
jrx+SPxiiIKfINwmTDtwxpjZCYtfSCDTrmlb7paCUvSFYX2X83/5lc2dXPJ9lTsz
TzsLpAZ3oOkxX7UcZTtVA/z4jMs4Z1r/IE4kBdSnM//dfIdr/79VH8XcifvEKGsG
an5nmiwDXta3anUZZyU9TWntlcoyd7U98y1AwRHIODC43RPwmTm5IBqccvz82CJD
CWakhRXMShcvU1smMufrJEF9Ow10f6clw9RqbWn5otH9zJOYxemAEUrNxQ2mPJzd
zSkzLgJdIeYMzklYZbXZ2hxldd7jBHBAltf8WcH50Iob/5T8GAPWqg2PHfKIWvej
qFImT0EKKcjbdJuYn78u9l2MgpoANDeHbhPjoQQhO3w1+tODwveKxC50U55k+e9x
LM3E0TslddDumIVqxW+Lhk9Kj5qQ64EEDis2O9mq9vTFL3qjPsfwj52gbruowQYx
JxmCfNIIzUmdiXpRxUGvKK2O1/Xd0UYQvh9HmoFMIx54Tp1iQblewtQz6ORcbO5a
4Z7EY7bJn9do3SU8VjnADjuL/53UVP+OfFbdlfa0AUhw6x2vNcy2K1BTdJL49OfZ
tBI60h053zAZd74k+0iXslHlptJKCRsx1hRYIrcmM+yB2nm8rkopJaSxDhAuEcWq
kL07+3VZOBz68455Zux/R8jL+Q4w4ebR2hD32CuoGyt1SWHgyvTWAB8h1Brk3d4K
hSYUVC2KOaX89XYcrBt0OkKAuJ9kkiJcAKJZ3i1EfjwonpktMjV1D2I6KYvU6ME8
I1ngtc6kEb75uQUFd2kT00+mohwcTTI21KQVQz264c1Yl9wAfOVrGPExxAes/AqO
fRwmiPCW9Uo/TkJdZ6PhA8aXfsk2J2YiJmiVYXqqv1/tVgmritOKD4mdVkMI4pig
iryK+kpDRaztjMJopcWMDNqjPKcj0PdEe2ebBuscZEMMwW63zE8iEhmB24t59jkl
81LTvxTF2P97hblrZtlWJIlKU9KDaMZ7wqv9oQhFOYQNArcDzj5gGjha7KG5el9g
RAEBW/3s0VrubX5IRVn0WvZljZTVwCkiH/4LQvbdbLD65FslKPpNtbZ8tFj3Htjn
2ztUWG5NGGQRYBktQm+DbLVHBbUtZy4/ppFbeqGr2JIzEEGmTIc9btsrmaTsB0x3
Q+YU+5WAsDXc77jjaCJe7TGBGxz0kX4tuSaukpfoVU1RCa5GfuyMZuDEg1kaacHk
xy1JYwMxb/LaxzblE0dEXlyWD8So1bqNaeLorcwShbH0eYZBbiscvggCQ6GVoZTM
2uoz3WvGiBzwWDDx7WVApFYnBp6+7MMd0Qm0Qo8hN4Q4xy/Qui1IhQ0uZeFIU5EA
nHutHAEcjgNGzxurxHnTuxQ+PZ73qct2XHFqKGKbvd8P2BfmCARyFDR2MZQ9s3pc
wPiAr+km64SNLud7ariPQL799TDYPMTqwP6CghrZHLfeh0bjrVZVJ79GGxxjuqHs
nowCrvOlNmIjxVXeVv0wJadT8vsgPnjXga1ssfB8NoQfeNC53fs6dmFa8lK3AFQl
QiuqPPFbyGs3/Fgw1dXYKDIBMQUMyLi6OX2NQy95LVbLuW9JM5uY8pUtYbvdbLCF
vRcTHwF0azP9a35q/LtWNjr0Jqri/EXx0L0N/Mg6cqqkDdNUztPYV4wZC7Ykv/uV
nO/Jc0g43XA6uRU3fyM3R9VCg4SVYBq+54huudTlhPz1+vhrMBLNie5C1vM6d9XA
n9gAsd1wENtw+9AIf15QSnUrYih4C8uA4gaVyudxOUL8iLmBevauZ/pVKCh9B+6J
UxNrfyFGRDuhQiFufS0IgekVxFuihcc+aLmUKKu1BeoWfD2yxDD+JptBvQkTIBBj
x/wS9UHTGxR/kxqlj18Pxo3fz2CSur/I33iZx1mFORiRvLSX4ZjQa1h27s+gI1On
RihM2tjnx9tzBgom7CZXsGapG+2JDK/cgm1+W69y5Z/CS3Sna2r0qG6cU9JXrpng
5eF2c+IsZ2zJHptaHJOl79Wbyk4gjlzJofasRxwbOyJmDRdoNHyZTdCPTGOEFyGe
8goFdWV4TQtGf21krjCb2Jx+kGHbF4d5yRbf/+N6GHim1VFPqwMe2Knq+KYK8TpF
ZJqIap51uY3FdKDdmr2GzZPLwY4cuQl4Fqw5ok/XSLeUeS1PPp6ZTCely1ZxKCUO
UDaPh6Dhxlri7RmsdkOqfNKA787zBx/upOolsW/VWRHZljH/I2Wg5yXpFCFRQGJG
StNqrXjTqgjpGPhXKz81NUtIeiguMoY9Av7tMz4lAcZRWPsUzOKux9+3RU6H7Z9Z
mHSSyp0vJ4AlMlistNEfejDZvvkSjWdjXMe2bNlptXk22VXgt52myIPOEJsjVNhO
sbuDqG5E4+Kg7mV4O3ZjJqE5Gr/ycwV8xvpE5vC5wJTkn7bJeqYTQKVuoLzywl+H
8QHDnzHBeE1ygFEj/jkS95+mVQFP0rN0NddhDKUEVSF3NnCYTzAKOWicBd61RUkx
DVsJgDRkTrS7/KD0/ahvpa+pJpXTbYiNu1yyX4q9BtbmOrNdjxpl5kkYUGNomjnq
MLq18DsuZRtdgqg132zp7Y1Vpv1/6tN5gjlY4vGjrwp0KFNN+5NABfbIsoN0DCsn
8znwlFi812+T6YpqToLIDCHYElPX/RVn+1mysXcl95Pi3ZfPzp/6A3yke+ke9qhZ
8qyqC5lUG8uR9Bt4MBI0tA0uA5vJDYYxp0HrScXrsOXO2GKCDZB/4K1EQItemER5
11xp1qEB0IV4ne2nJ6eaET1SF1Fgc9+SAe6l20pJBr6xDFsOCfxXIiRXFtyUoZNg
5as8fUKfKad8161JgSqHNR4gUu0g9OTKVxLQt8/UA9tT0P1w80JbzIFhuCyZsvl5
DZGvXKn5BHOCYYct7ljKuLRYY5PPBZHCZZ4T4UD8ELPZjQxy6sf5yslgHnqB3kNI
ZIdo9mZfHBV4rpD3JpkaCt3wP7yLGhzNJXoSxwyb5ZqkRfJ3ShH2m04+F3qPSZtt
zzcu5w3kHo2v2TOAmmX9DuVggQWwopf/YlnKIxzhvKRFtuZC49DbZmysWdzzDjLR
F94Z6nG2A2nG98D+1b4HBiK8N3Hq2z12FDkaWICA8i58j0aqRBRbXrlccrH/2EMN
2qBbPHmimlG0jPiVA31IbBf+IaOEfEmaH6E0Ztbre4SmmhtH8dV0zk+seyzeA99a
Ug9mGuw8k0/HPPxAwSAyQzGXF/Pur8hZLoSY5HBVi2qZUpCiKg8PeZoydGZAxw7O
MD4/cShCy8qBn1dDJdifKUNEsCO+BU0/DsgNV+gHr8wIlem35r2+idsTxUjeWkip
VCJ5yUnVuN07z3VHBy3b469Cy+upQImqzvqucZgqIrrKu+yu+FRUZIcUtN6+d58s
pqW5wTBT5m5T0zgwZ/O2RuqVaSFPvxGmY+L3ChMY+Xm06Hy7w/zseIHy4Dnlysnk
fig1l2NrWDlioUENVtPzi9pJvuG/2QX55X8RIdN1qwmjzDm6iiBxJEANwjb/fLXz
Acfq9VraKFAzHY024DFj8IURa8DbWvLHqozGnRthBAIC353FBHyxQ3GU7YFmHKGr
uBEBHFZdgksksifvXuEgJu5OztiA9crBNaU2pNcvxEpcNStZGpl+Fvt7+XwzkQtl
JiRx5sQm2sQJebcmMV9DKgfdIM0+dZPwT40X+L3WViKMsknIUUkowmgG2Vpl0Vfr
iOTPoZ81yYiMtfmM7iKQ5EBAUHRicy0DCbScBEHuU10Bp00ZvhqPKi4XKoWMUuOp
EVWNE1f1dsZMwh3Xhy9uh9CXL+kf+dAOVHWexaNxOJdKwJMgTd8qnTYM0z1HjunJ
DsFIMAXRXH9vzwH/IqCeEbVN+UWhHA4up3kEXsIoxETjSLgXlToP4Z90m6S8auIF
X7QG2xU9fK+f63h5Et1G8k2Gh4qHd/oDUgYF3VWx5dRi7keadKzFSTkipD3nurNs
DsUFlsbnWrt+GPF5djXOrL7mL7ePlquakrEP0nJDVLM5W+Ox24w0ymvaetPut4mF
7WhUvVhMN2R0RY3KOERJdXi2XRXT2AUcnEh44WggOyeePe2yRj+uGUqm23XD5+zK
ALwUnavTtse7biOPmG4rXlpFjVTy9mbtOn/UQVnEz/smhyk8Gw7QhxWrsw08GnBp
6EX+40wE2weaRjwPPIZ5VF5Q3o+d3CUloIf99thqvYZzG3CJ3/IxoQQOGiUM1vLe
155Jmb2H91dKFxOBSw5Wa/dVcrjVDl09xYWM+11ptZkITZstSs09QQRoK6qn2Tw+
1xg7smgsS111HOzwWM+n7u+qKcxoZW9iacJwPHoBkpTQBt5GAEG0TQUY1HdDPiwJ
t2urkl50fw4Mi5MOnXs1O9+OJvBQ0E94AZ+PwFNC7XVr6Q8HQspTUNNe/cVAi9Pm
/JYVivnxNV12zRcok/I2A3GVKpfoEHHaQ3Oum926qKxTsZ1gj+fzFYLJY8FvAK7K
geED73kboj8NmSsxrCAsqmBUCqE9XIUW1zRihfM8MNhtkw0+UIGb+H97+gssVGgD
vwr1OeQ33BFk+MCLB87dY+OdQzwGmtqZDw++2WeIYXLlhXaooqkppX13XC+pv2FU
4cXuTlO2Z+EpR80mIYxPmsAEI7O1DcpWU3LWc4OSImTXxHXt6CK78+5qTmkmPWeA
8eTfcSOLvbmOj3BDvUEHcr6thx80O3Iv4bsW2ya5QBTA6Iee2PekVoHjPF6e4VBu
bHNzVWZHnh6L20JtYPpKg5l0ewpoWrFnd1OARPxKXd0kfLM3f48F8vYK+DqVj/jq
jk1iTI0U9TnaTPmJmx8kJouIzbt/M0Df+WPpcT5603/j3ce90V9tPd792fW5G69u
EA2nhGm+RLIL1khODJUzabA4lcbLBHWhp0mQH52mHluEfevXIF971NylLF1CxlyT
nrGWfUbWt7g2aN+vm1+zayFQmf0suBkokmZ26K/MJ0pNL+B17EuaK4lbjD3Ec7x2
7A/xWawIoGH0k6fsNMGLHrEXqIgYaC9WQy470Ih91vm5VmPO3pL6YFIlquU9dcW6
6Rz57Y5vXBLykhlg3zkoizhVpHyJL2YkMigTlYrRPujqOwk1K68Ms0AlyXopWfea
X1Xphs8dsSHjzV3YcUwDj3w+c+5+8CeM2SrnUfTJScCm3IBSZYvkM/jbp4eLLfPn
zkBSXlPs6Z62dmcBFc5oexpw9dRVrLGfU74KEvnzn+Lhi211v6a0RCqUhyrDLSQW
e7lNGOeoFUiST6m4/X5hv/64v+lKQ5K5pmhUdzg5QVbUfLpKzcLUdUhGZwLqJyax
CC6FiFGzIAc1xssz9aJZy/LUJwqMMzoOvs8K/83ZtLTMgwYmLhytVMYmKASbz6Gs
Q0Z8Ap0l/+RbZOj/WZOLsRN3w9R9rr6+M6R0yZkIoE1BByDhO3EHaqlkDYH7kZR1
Kp01uugJbkSf77r+JkkL1l5GuWS27J9SGABnJejitGqUkQMcTyG8f8QHGPm1XLRp
hIHnqwGhzPNx+iLeZf1VRC1Ar/1fR3yi44X/n645g4f/JffCxskV2vdGAXTISlFX
I+sa1Nk7vGLlr1A9i8qzD2RmpqPwG5AGfDasLHbq1WEnnsdHiS0rFeRrUs+zggl+
vUhNUT/h2IjYCsK7h/nMm31X6jslz4Qsz1irlutwHu/FFSJbYm30c4c++AkAhV9x
9a27Lq+HE4v7dOrfz71uChD1Bn7Lf222ICumZczkS6vLVBjgmlFQAa27dOafb0Uk
HiyrJrXfeY0D19pA5a7PMKt8FwbIhxdtIh7WYDpKR8+AN3dHYm1kqTymQ7JEUtbb
wXwLrqYjpICzzsRFoyUNdugRm7pVP4XY4QRgOEAH9z6h1wZkLFzVpy7FlyLsZm+G
0RQVtuNSy5dbXG0TF3Uf6DV86uxjwvgmkmZDtrkclRQqoqpXrrWCiP26Mc/6XX0V
F1B/q215vgITpMJT/DI8NnYK20dZmXzlbnVgZceIYVY+WdG75Nqh9Dn18UZwg1D5
QQHy6xMDtzaOqELj/wyQosLTkf4m0I7PovTxMjVJLk5YSwY5nZLcTxcgBhJwCwd6
6pJAWdTE6i87GBj5C3tMVIB1GLrkPfiZIhRNezpub6cXLKefzjvfoUkCTh9kogiC
6V9iwqU/VmcQCQgROSk9vbE5xf1jmXJs/9UwXp7qQ0DyeuW3wVZJJ09fmtemZk3j
P3tiwjg4LNuhBZt/F6TdH3GUguToTKcPGVWqQ+pMPxpvBH218w6JaHXtrHgRXiUM
3YijbR8qssM7TXoNc5eUG/a0dmxtq4oBPGx5RKgbyfM2Qm4z24qQTAS9/qGgfV7y
/cD+nMHoLJkC7GsXLizeN2uvc5zF3DHB2S4mkwaEGhOK0ko1QM7Z60gYprKfIgDh
DXycg0fG60c/bkQGdE8f9ZCCXBueQPAZnzO/XXue2CwrikGIOIY8/CBQqu8GK07x
VQEP48s6c/jQaQjPIxEtjvrmAwY4uUc0Bp/EcTfGvgD83opPAtzP4o5GQUapR8aq
LXVE25C9pe54s1oLr+24keCeYUjgFy+9mrCR3hhcQpxEu6ycUmnMUtMqSYDGN3v9
thIFNJa39AKPEwG25ZzGvotR7qjId50xi2z3ue+6PiaIonoCJ+IVy1leNTra+ilh
p90XD3MAujkXwjhg9UQQI8+3z6o87mkTktU5fM5UjDOFQYxUlYuiyutta669ocLe
F6nAHA8rtNypfzKm5WX9GaMjiGUAJz7PwDyfbsFaSPZPsF8SDxc0KNAu72D8r+kd
84rZL74odMmIjqOoujwr3v7EHGiX7WqjzeWewp01rnNCX0hKT0motYEwETsxqiY4
EKGponvEBoZv8YTvdz2Yj7nMir5bcbTlA+yhhBanXxDw9T9z7syZRTeE73mdDC5X
0GL3M5mwZ5gi7PSU6FbqRBbHwKf0xpFCiCPJS3Z6cvlUyygE6KUgQrT69V2MT2jB
s24sqNuKj7KUVjmq34GGC3011R1grVqUYfdPkPGBubt3od64Yz5idPM9FQaXtghZ
lwMacEFbmF28s764g4rr6RqMbJayN/AUMXe/V3NGRaEDgbL1AqcKLNuMvtnatV3w
WwjelrKOuH4dcvDmYBLdvAgdxHCHaCPNj6fZebc901ivgtG807o3egX+SHrp9+9q
TNrXEm5PtwS4QXR73Yq3+XjlfLLrhvEGkQ5ZmJmU23ZZBfUA3bA920FLequJJBta
7Wdg6YDHhsOV5ez4t57DxpK1598ipfubPxBMLuJYsbthFxcobkK1jgdCVhlxLV4z
JJR0H9W5f8tea0qrcniLBskUHt3neixBZkGv1yzXDyMQqxrdhjYjsm1D2g44eZmM
XNXMKA7h9UxBbv/PB8ABBR+gTCkUAEAtCG5c872BhSClOYrV/dgxpTYxUe/0lM2X
VYxXxE8q0ekb6vOSsNIksFMJUhfkfyNU/0mgGPJpOg5L+7OGpJt+fAMHuhV+dEHl
KRBIeMnNARk6zK9JN7oFekhL19Ycctc0ZkfIByqKauY4vxZrmdqkSoqsYywjEfqb
WO8MN7agK0UXfBnA/nfxwxxPjelL8pN4lFqrsHF8w5A+w+L9cvKgsFQkj7q4QCFS
10tx0UqOKNcS/68CeTeq2Kt1YF/8UMl238uhRhqmR0bg2XvyAIga3/6LJ3rEYlWm
tT/NHM4r6OqQ8+uQdvPEkicu5F9RRyHIa6IkaTYB3aLaNtBTaKDJFEhwuAnJwXDs
FULsFUaJinNjywKPlx4hb3w1P30U3ZdvwUyFsobGc4c0/H5aM8g6yCAMxPdNGVh9
XD2a+V4MU/5VkjiunGT0UZAC9TC9TyyylvMmzUZKeFV6U6b4iohHcAu145gGDdB0
HG65qLZPZjNQEJ9u6flsNT2BUI+5QMHfDn10kphCsOvPY0oAtm2p07OgkCrVTKvv
yDVTlgU91HbeUy4l1KzdozqYcE4aE030YUo4Slanl82NRTCj2YRKy57/bC4yHRYS
xq1Vmv+GgyiOKhF/CyrFFfixtghp0ljiFiG+DKRRkgov7mvrNjJ7zOIXZyYqVtxj
XGdD0O4b3SF7uG/ReAKP65N3Y7mmbpU1onyuFHSiyny3N2O2MdXLL4rR9OMqfHSs
4nB5fqB+tYE0l+H9DZnLgutfXFvzSTbl/RGccpOeXiZ9g6AU+al8V6V4IA7FzH+P
P4Q/ew+HHUI1/cM3yuNFuA79Fc2kj4cKRHQOLLXopAMeTRGytd9JWcczEDa4xrXf
i++1mr/UhRc2xT4n1uTLRBipGCVHmQ806jYZXUWMqB3WotX+QqXIo1PuzUfWOFuy
rhDsI2KPYfGhQZkFUTDz+7g6K1hPmvmWnvRhlSFz7zElclEtMfOiDIwr0VGi27iz
AEI8Fgny8mekYePrdUstu5IfeE7SkjY1Jhd3arOYVojSkDFjYRwr3pgyIpf2QpJC
99OVFsTx+ccEGItKk2C3zURAE4FiVs8XaoZCX3K70P1epUUlpLQdty/pUtCNl+t6
4ZeMfOnEjwa3ACo5OyC0Ra2y53kBex3piRnj93NGwnZF4ts30tuyasv/p8sbf81s
NkPw5sJapDtscF4W7Rn1AN0FI0IAjXY4ooddiewHuIpm2wWnLxa42tE9y6hLUXJw
WhFofKQ1CKc0B8j0wF7aNFAmFsCL9t9iX0cYqLQvh2wSXtLf6oMNs44iarVYL/Vh
XUQ1prMVEJa+Ee8tDtoSj4hmqthW7FpRWdis36DByrz1SWt8AxheQCuA9CQlrbzT
IsPHRHVJe3RSUgD9PeyZG+3UB3BynGZ5r1rlq5UDFMd6SnDb/SUVq00hmzqZPwub
ck16XUkheF5FT3z6IYgxJFj+O6MX3itkT7I2E1Zz6syx8xrQ0UKYEAyYMdxjklmO
oLGFhFuue5sUDEPiWwF25hJiO/UldY06Tp3zsjJeHjSHiLnZ8BLVwsEpX4euDbLJ
KP5E13Sylqo+eBEE1kDrQjeBYjoInHk/PuLISb3FraNk6z34vHBqQKT+7yvpU6YJ
puEmGFZqO0OjZIlEn9auAk0aReKdYF6+qh1v8eHFbATDe3D3qfJfip1vtfBnTbY+
W+Wd8jBiVyw9HKXTyAqI8JMZjmhk4Cz0Qph5sRjEA6Alwf/x1VCr59+m7NKgGJMT
VmXsBD+ljlSFEN0r/U9Ovt+Y20DDDAJsd0xdUw+nJ5sFPDP05QOpO7XsjQDhcgpE
HxgZJO5ZcYzfnHFcqfTdDhG1nILm8Qxbxu87d3y2pu4PX8wSQk9JmNqyXJbKPX5H
WFVugSBPE2lw+pRHQaul/P2H5cjRTkzi/KoVXFCvq6yaSeJpBFq0ATojksuOuNr3
QZ1jSBAntIMh+YC98MZAgdjMM8aBu+M8xQV5caDmIIAtB62RoDFotJSDx5lL/MwX
cVnMdpdGJ/Qde5Q2lMTbtz11cEgjpq64aucTYOdEj+21d44ADMlNuoxyB/NZxSHE
eHrVs5fhdvAlNSg5spOYsUoowSymmI8YHtqT9kaB2bSEGAXgqjNmYBW+SqsvSnjb
ClKTD0st3m9ZJ1sQ3pJvwWoxaVbuyxdFF3Z2lrwQLLShZ4LgqGzhUno4sd5/NQi+
SjIya7+8TOCktYIyWqfV/0A6nex+BtPEt7dLFOursNrJErbw0kGttfzwTrDEQoyD
LkHCcqlld+++jCvPZB6dZj6LyiFgxMMpir/gfaGQLbY8KfYlLi+4jYiGm910lVKi
Qg7FAtfDdEdaNv4J71l8FUjbJVRjzwf7V+J7EtPxTro4NMTPHRiXA8O9LlUoOp/w
G0cLnWJHF1T9MPoL7wq7ckWXF3rIp8cZxptmASMsQu9da+U6i8iqNmvXSnLoal64
WpUxYkFGb7GuRfuw7QFEOEYTmDVV2i8yI8U7B9bvo/k63SAl4V8Vd/lvNr7Ajfw1
52Mv7y7mn/6IG4mDfl0+uES1XcjJDDYiCxYaQA7unSOKNrqvvJvr0GYp91u9ULcW
y3Ps0KO/LiK8buzR5+q3CbHOIOf8PpU2ihdryQctyq0DsS5FVNylU2VVzdiAMI4X
jtsRyNyNGdikSrNRV8c8gXO7jM3VqnPSZXj7QieeT0vhofgBfUff+pxlEjkcB76d
MVtML+19FN76E2sQdYZ/RiDO4H5GP+h7gD6FpnHAIQRn0XJS/k/P/OHu0qVE5DHM
DQv9QTHJ6kljYIZo+zUbEM5zP/VjRKRq/UMpN7wAqWxS5sshD7kcoyjlPS4gkutE
jjK9yAaiCMrB2tjNaJdch+1cdTz/I0jRrnSRbCX+0VG6+GeDB9I9Q7TIWYpusSP5
o+wAek4RSVm5FaYvLVRRXSLRCbH/DqN/4NpsdK4P+aXYG1pulfpCOHI7+GgHDPwW
5P5Aoze/wu6xtwAgcv2zcAeeZ1IxvITkFDmsageUWTyXa7uKG97bet2HgMMKFNTB
6on0jiSi39HMINFskJ+OutP5ciYYlPrqulI028n4GAk+YiV8fOUDfWIXzSbY8e1S
EcfJGePgdGz4WdQzpU9Z5iFUCT2FleftfhH6WNlS3tO97oofWLP4XpEXtg8i2HH6
0j/QyF5jzVCgeFBDcduR3C4G6jyQBWKRhD4X6AgoBGBJyRJK/Mi2ABvoHQG9Xs9v
Fu6a1Aq3fD74ZwVrJoLOf/HNI/+ASmeKssiNbyXDj/ywr+sGRBWODCuYdsqv3xcJ
UPSscTiDvQH7NR+GqrtIBgcwub6R7ORvga2J7YQ/+zDUAcAjVtpIW97x1vwnDMbu
fCpN6QYt4ZAH9UgjDGGw6Q+n5KM0CJd4yBqUHYQGQRRKn4IIANGI9d/y2xfQaIBK
Evj2hitwCD7CTeiWYTkHH4C20+I7h9Qjhle2FOWDzKDtBU9Vc5e9nVfwK62g9KHq
IKTeY7lxph2gAR8tdD4u8lm0+3zkgbm5iGkrmG2e7bZ+xwo53TTUH14LHKw2NXnX
JOUtknvdW5FnPo/Hs/5EAkRQOpqGekysaNXZXJw1lOG7iytlQAnVKW+SCaYniGru
EevGrq4KGn676nxi8f4eRrVxD0Qnp43zJbEPoiEzjgaizjLQY9jWXsIm7zVlpjsb
2w+jhuye9rufd+/4FqRmAgdKxCEnDdbPxbkFLzBd0RsZfBVUQ+nttXH6aBYnaaHX
BzecE/8r2WQaWf+Fw6ZJv7ilF2/lCRK5gG5tdgOF3rOM9gNcu0IMrxcqb4ponUvo
rpDIRyExqlD1J1z4KJepnkXvheiiAyxLR8+3uHUihPy1MJBYxrf+wU6tXMpAwfa4
XrrR9aupRTP5e8cwSjAsOYzogb8oALo2Gqz+fux4Lw1yJkHXXVZfgQY8HdxgvBDD
SVzAEl6Zks8AYa2gaEi87P5ldZml1OhlJpXr/as3s7cX3J/sZrQGTG3yJ5i3cs/c
JGatpU+BPLwSZ9SyVap0TFRAi5w/nJGmWR0mkjUJyXEuHH0IA+Bi6QmxAK0OGPxJ
MlgqSiiygHujytrgGwuwitno5H2q/EeUMlNPgB50vsvCbBEXY5xBGM8l687CECvg
ZggmaSLSXpWYtQy5OcloRHYXDTbVK1+W3BT5rT0c6p2UTFkuoD9HOjyJz8QB8RQj
FWTFXYLkbZvhHYG/nyHX6bsgvQH7NwcMhZiGa0J90J7qkfbMgjWiA63jqjpKnvK/
SkazGd359jO2N/Me1nYDOiWTtV2qNO+R57sSGJIW8kfyPA+hQgHpAai0WzbCialR
Mc6Ats+CWbeexKwyueT6SPZpqDpJMExzbW46eL5tOeIjGQJTRFmScOnDLKG8tE1i
I1PkOFG/QuiXNyGY2a1lzeDxWCzilhz0AKrSHWThi82x2trMFRC3YB6Kpm4lmr60
F3DvuJehAUDeISSEh7A2zZHci7LD9DLzV4fvHn93c+ygZuRYIc1Ws2JNG2mZs+4+
UD7I7d2pUor2bi48PoumXgdO4e6xRie9B1zGuaWn0NbR+VfP5htGpEhyyNAgwAOe
oAZYvfJeblTy4LUJah5oH4LKmhrRFZ2K6lVEgrPxmapMdU+3gbBg21hP3B9CRIaR
xxbrJPQH583SjZI5yem/dMCbuLNBSGSTHbeb/0YLxFfffOUq5Wpkjj0sC5oiR0L8
T0Fm28e6+eAPxWeo8PvfuFFXVbDKKo30A9DNk4syOpbCNCcKNXJdCswoJlVE+XZr
Ag1GnXIUs4tLMciFOq7S+DMpJYQTNAI2PhpovlORAcJvXWdQV7jPLkaU1a9ayvaW
Zm1hdxvuPw7u5Z4fQKaTuRXlyaUN9P9D2bQTci1sYVH7EkiR8kp5VI80vqGSGBLO
vAY1H8byhJBjeh1Rkpom8hQkGCW0CBDnLnJtpisqb59LkaPBmbXaXgJllrDjRkDG
bi5mJ8EGiTTYKN2HJ6MpUMyy25h6ooSsmsCz8fgXPjMCgEfCC8LPNZLq86SSe5Uz
k5UXxDBiLu/l0Y8uFzPtdw7GMAx/dxvXfrokvTgWfjCZXutIAXwWApdgNGXWh3mX
rQdlRcEmvRVHNaCw+t0Q8S5wzJl2IcahwbhxnuuYAvQOYzqzxn6tjIvNACO3wQ0C
t7bXYCiauPXZD5qGT8k/BYK5IVJ1AAx6ORoFjuyvTRxrKVgb1vVNqm2F3olNYpat
k4YGmj7o4VI+EG6rPyFQJWUrQYT1HxlUk0CdBq1n92MMFzAL+Nom75/UPPSbW7Pj
VCXLgDHSNSD86u5QaCLHeXf90Zlf6Brrk4i8HUn7zH85zqYf3YJXVlbEuBUDrv3C
rEysOfGvYJRyHrlWC7AcA+JNDZwC9JciYF4mQywoy7u0tEHjGGXoSuWuB56DHqtW
Mo/1XpsEc+dpk8pj99CsHVMJ9P04533I+WaoHcQ4d/mjx6xb3rwMhngy4mJSyDwi
qrmtVlhkInjPKrpjV8xx1F//UEH2aXoE9ST6LWroG8QX4OML8x61UP4r/5sGvYdC
AcgvcJhBms37hw8CH1rlxEirFdgi50h97uJhVI5BgrvBzqWfU8FCtOOzewBHzxgU
lb4DwS5OWxog5B9gKKT1aQLrwpxGzuKcuBXpRwe+iE+w7tQ5SlcBuFgFzML0EZNs
6CqpZsLhCkarUqMUtDLyvm3o6TqTzfOiYdZo8gicavYgfx5h625ypHJIKy9uk1tu
8D5Xi2dFv64WDiotT0+EGXryE08lmGIx14RlejZjxz69vCr89RbI9oBCgLnNW+Ae
ptqiUN/bsz+zIb+6r9pV7KmnJwTdoMuKKkVhJps34nlsX/mMC779uS7dNGGOpT2p
dju4Aktlg6RMgwLOPxYi1cGVpz7YiYV0tQh1+cnEXcjUtiyxPVtDVXrVqwSoELFf
XdbxcB0RRtVNQaoMYkEU0chB//7d3anpR8fxOFFhrVt1SeNJe+XTvqF6tSuSvRCo
/pqDJDyB/69f8RK9Kwy6ooXDUOZBF9hBsrx7BFCy3ABXzbICSgRvTnyKpPjHORzg
IT670RN6hwRPSydZtsuGpRIkTtyUMSo+1IhTUdu81SuFlJWjg/XX6J+VXl/xXmR+
gTjtEtA8yE4UiuPEa+GTo0OrNswi8NIIOFWowxc/BIZ/qIN7psW9YWoc3mcwWdlb
ERber7OotqnrW0gWyWGZsqnKN2bVhaD1ne0dFc22qpPRCRirXt0DuQNR9GO7/KBI
PzGwCr6Z9+R3ljKZdQl4eKiQ02Rszft+K8at/mY63piV62rko+ugs+CHK/m+oAUQ
2K7dnMYuHuDVvrvCiA3i2xjalsPsH8qvE3pTWfVoi6Z/uy/X5BFswOIx0gtENi6G
XmUoT7biUhHdh2jX/SZM6Y9PY6NzYHUAsWlm5H9TM4N1uQnw39DoNqfaqoCqr5tN
qOpVjGj81XdGFwJU5siAem/m8F3Cy6+jPgqOBK3fV8Ww8wPhrnsoywO+BtLWEQ9/
99m/B122U7jQLuLdMFasI4FrIvWo6EmopZ8F0udzh/9PhmzqSDoG3bDoVyBGVuWS
NMGwW2bduq94pUiRtl2CcEJ/IoeoooqlW90IkeaB1A28KJIR000htZWbWT8zjlKy
n2iCMMGGvll6zjVHTwYSH7MDJAhTjpXwePdxAcJGvy7yHTDdfHUzYuCOkWrl4ChN
X2/3MOKMzHAybX66lcmxqOvVYf3vc7AxihddFVGXOwIEXt6MrJm79NTSES/U/i1T
QRWijf8Lj8lXlisjAOwDjBPzkVHuwg50gH7qGZ+BzmXDHRgLE7c/W0RnqdZxVelT
p56b8qyPnwQQbTpirYFYNKyV+KWg613zqLouAvGMMQNoMy9/GbTHzz4HfND8AqOT
KGesVLpznt4MjWNZcu2i/j+17NQuM4Yze9JLMAlhLCZSRyZi3T/+OUf5m+eakckz
V7z7zgxadKTPbXLUDkoZrlSGVKKynMtG0+uXWNIFjhtR44TF/fbE+M/eIu2TD9Iv
IzSrkwOuahN1vgbnTRtUgP2ScRavXUCEBwYj8U8TbdKETEnAPCHDLh8/mD07fGcD
V1hVoV0uhWeX4CvbiKCozXpKNcQfeJtz10pvE7j+t6bSF+jIQx3ByKvGLtk2FCMB
Hnd7qPiC2+WSZnJPp9pf8CIU38+thWg2O9UCrNVWl9gLI18cdlUOLv60mQng1fZV
EjS7rXv0NRvpcyyAFUpVyKtiswqMLBaT2rzsTx66ddmp8v89p+oYFy0GgwpK3cRW
UhDSoCU3IuD+Sqim4uS/R1PuT3zKC11nrapLZ6xTavENs7mGFX8dQ9dRslA9QA5X
XgOfeImdrD+Am624K5Sv9gUO6qVBlnT/XsGc+iRXhbGwmvbK5cjKRQUJ+o0CkFw3
lNlf67sA+0k9XrhZs6uKd6SxAR1FWJx1zDvyak3wXy1PxIoKTk6l//aDFMRuuZze
KB+Qr1o/sk0GZ31p9Za/eIj+FoHGi0NRWJJYTEF0V8XMCdl5idSi8coYYNZ8ELdj
cCABPxzBCZT4wPKiFscoaNFz9nDTRU5lu9Bfj4fgNLIoP5YmtwEiamuabO6OfYzN
tozgqom7xyZM6FTfMb4APCXvuWyP+7KCBnK3VY6YqWoC5Zf2vTogzLvRgj5Bbn0s
q1oEsFMshP/neNktLUbbiHcIe+IZd60xYk+5DvBM07vlyc5Va6oUkCYMS1pfjSDr
/Hv3+ASEbw2VnM+1RFOxKLxUXzW8abRJOE+XLkTKoEqSNJ9rfwfCuOQncmH0xlZm
njVDjid/ckRu8CMt/65F8GSAo1CKZqfIKKBc0VHNEX+YI0o8ZuyWB/OCKJl34oqE
gYZLdsHpdIDIDa0QH2z3pXrxyb1pi1FKS0WsmulbB2fOH5Ke340o2ZagcYo36DU3
YwI04SWhlzXr9GUzqpQzoPHI+2SAE2iBNZc/7LEP+frPHwdK0SA5QWhi0sD6BxBk
d8R8pMAzoSbmmf/NSFE0EbtQdVOVp2DQLLVvh2CixIfeFYvhOEKOZKSG9I1V9jhL
i5G5CGNwa0Cbp5HNsS2h0ZrhXyDaPAvzlfJwWJ64VgF0SErrOVXZrxH5PZwJV9GZ
zfBT9mHQ3FZ+cHOCbJ+pNl/hlxPZlWCem1WN6acV+sJT3UhUPCnqDZXR94P7gWfV
9h+z3rBqaALUHtFM2WbWh6aiiRh8UJXvmnqZ8/508bnZs0alN2NDH/m/uDG0w+Lw
yUHIC+7zI/mw2xOsI9Jer/Kv4cD+9wxbz7IP3jkbGawMKgFDDYf8GvsXWiqqvyQC
mdpJP9koRYSpufzoOk1gLdDbr8IQnJrx+tQlr3nv0yKWPEeBLBK0dP8GUyvAp7YS
mt52Mgvs9XPMlmbVBtFpSrDv7vqINV6BAxLbv2nx++ayIBi7aZQTN4w6bvpVK/1w
bw1V/+4Fuqkzrcz99XX1jQZ4EW3ToyxQq7JzKRzKAiDmJ8lZlxStl4XNbDcH9zu6
WoJFRpSa6Nem21dM4FH0gARaVVB8sbRMeU0+SOfSOGDomjH5hpzOeGq/4f2UH7IE
PcHwBALbLOhAg4Aj0jmq3Wj9AwGG6Mzl+54PmaKEE9hVOE/dqf8Egpt/vPdKbY7/
0FjPIqxM89g2Rx9SmH73Ev18xQ5xrI9kKIzaeQQsKoRj3dgZyyOdMAoDIuQ2z/xf
XefhxvwXyPS/2Jc/VuTvphKxcU9q6r9tEHH5lcgXK/w/8NHYvH3/KCMFMIR04tfs
nqZ9IvJVi82eBxP6lReetW/995ghQaGfkR+2vk0pdjPc/gLuOjOWqF1f/sCZdwX1
bLQISDJobB/RsSVF/FxUeBJsE7D/7fsVtPikkVlmKyeA3dUV5csak7Mi+UfAS8QT
mB+6slk7vGfb2hr9dacsZEUFB9DcZPaS9pjB/scL7hRgNTvgMY/FvMvB0Ht+GlaE
1tTd15SCkSc4xjtE/9qejbhk5EuHuM4Wjnwqwzw/pYRoSjVb40e+wMqtPLfV+Vtl
RTl91GRby7FeBmaMYCMZQWtfVw6Ms8QYUCysDgAsoi5SvOta+hsQ5AA7AOngtRIq
iW6D/7Jm7fQTbUQQIICnXYjc2juL7ID2KQaQeYQvCjn5662NAYZMHHBrza24BKvl
VEsXkcWCp8IZR9TUMZ71ZGH9beNDGvvvSUV9YRLGAk+llVT5LMD4wtAZNSWHCM/6
Gt3fMBJUs8c5qaLq2kBYPHBH13rA9Oh6by40uJnweIgg7LBCUt5eSv/YzOz371oE
CxCYrwEhDCyJCLdz28AQ1aYrAMkRRFeY0R08hX2R39u8OV9x4El3xPJ/EMCfyG/X
1l/WKEBeypqYqdyu5paM4ZF16H4yOMcm8kp26YxUMqHyZ0ncnF5Z6PV6VrkfECrq
hnMCo0gseJPfT6OdSLVnjNh2Kpm2C1zKd0ozzMihx9K8F/UXMlJdwDxCBvTg3aia
ZhkUaDg2XVQAbn/COt7OYgQPJ1dNKudXwTQ1QwL6UdAG4Vqzlua6uJoqxHyQ2PyV
icJ0PhL+1gx4+vlFPSVxHPXEXZR3MUEnOqGW4EjJDapjmJQ/sD05j+E7of6VM9Of
ZI7RPU100q0jM3ZSN4gurCtRaKKDr10D/et1HHc1ZpeSTdH+opML//DNatQTUgF9
hpiMMt7T/UTRCjFCBmdgLQD+l/YiCmgmULqpDF/adtRvVgFsynCeaMixmBPDrfno
5sVgVFlML4dNbfXwUAbZG3hndRz1BN+FMqsEHu5ojGkUA/tpugHfnc3Btqo0RVSm
9vhVH+q51vis5lImg1c7ISObzJytBPZNvgmKAm3pu6nFqGORWegjhdeUhnKtzAhj
rgCpx8nSFP7LYxdf4sGqmh4hDVgINpgXmQe+oxHc9N5t/PfqJZVT+eYDj92Nuigj
PUvZwoXabpU8VkCNULoce5MAufS3nIAAg91aWFWVoqZHaTb3pEyYEOgdMZk8WycW
O5jDJRTrcNmkpRouUWcPymIHd0eMCjF21TVz7McgapH4gBETT8ers2z1n+9g522F
idCSXbz8vm1zDTk0epDM7cNcIYaCOzQtx73/AWmTGgUDDBVtD8wBSuW+BaDSR/jX
EPUzpUKFHRywR8HsWagoLKFJWcioK8ravwFk4LCEJNPOml28BljLS3wWLfrny8ud
1hs5jZpKloUyxp2FJEIRDRq9c511pMe39MQE6JSArMT4hTe7Dr0Lwa7JbNC0IiH9
KVfWvDnpVA4iKVKF8ytE8U1CvkoQh+CXqyjFZ44F/cld+PUcN+xDDHjfIIbklpgx
EUfBrtnUtQ4Y68P0U81hI1kACyOR7h5lZNnHoUkg5csP6c8cimAnspaBGgbJAs27
8sYEkiRfwBEbAfnelyYdKW0g5BZxt7tIsVsolzGhFXvRwF+rQX6T0gKRvxsUPN9x
G7v4uMFy+g9z3vTJEbkkcXqEHxMFgNentnehoodRodG+sxirOPtTP4aUaCSovzWw
JQe/yBHErAdKaC1fbtktgbVh4JAZsAhZZrQ2/P2UKTEleke6PzvZL/uU8nHlycIP
UeNl+LzGpDp2mzxhh8DiLN2UrR2SxccHr1qo4hNFDTGyv9OGHGLCyUSO7mvjD+Tb
S0bcfJttyEooB/TjTl1geDSip8e2nZDEpJmrEHgjhCCR2OGYr0OsCF76AU6lyNgz
setC+eZ+yr1cWRWjYQp+Z8eIVrpo7tqXMuOMbS7fvIhmMPzXrzMci+CGj2xrYLwT
YDB6JRypMhoysoUZF2Im9bZ3A7VhN+wTFM7YdEiobXnYW/k8gttwfHN9DGVWPZIa
5BagoWXgm93H8Hw3/gacbZUcIYSFw/lLBR0MtbtfkhibChNjwge8A8BbpGp/Ld/H
HDbRhsEMNYFC+Ihabb42T4ieHtvQocu3/XnAOgw3PiJdVZhJjFl1nKjEM9g2GAkB
ijBmd4VM9YxAu73JVlc2zbgFFQiPB9M4OA1rUTCJBRZ8A6/TI7U/5oKm3ZRWAYBB
N1S5GasDapiA+Dm9vQghgmFkX4vl0TmXCq7P1L/LACJutKFcsuxuW6yUoX+7ctIc
PuwDufGafZPeev3Rkcez4Je8wzuPiXJlYXVPghxKT8YYUDhpIwqDP1CXgJw+9zdj
3zxEv6vFtbCiU5F//sQmMp18as50YnnR7PukKk+6EZIdeqK328XtCC8B6qnYPQn2
x3WJzJbprMEmspw9/vnZjGhmXFrUTxz+uIXTCNJc0Z1S9FbN7E5+h1fZyUypjZyj
uLaeErHJ74qqnhRHW89HCzJmHS09oSnAuGcSSNf4Qs5eDtQBKA6rSlMB+gUswJJi
7WPHO9j6xfYw+sEAefod9FDzwTuqXGOj7+ACNuHha9m1V5hoRfZpmWigidlaKyLU
NjpPXczFkKOC3v5YZJDBlIQLEIha5XH8DDqYzhUsyRmVTodaGhDSnAxCbRcd1nYZ
nVzFjJ/KourTsTxxx7XXCN8Cu0RvDRSS17WAlaiZ+qAYHGI6U3soNtlShL4/QaKv
1bEyViWWo4fLFAV5UorP3hoNuTiP8A7jJHSbfMjJXgVTucP2Z5na9EOOMHLy71Q/
NXEP9/REZojXtq+dZhC8+ZrQrfgGsNrgl04D8T6lH7raXVIugVZYi4xK+uO/SlIJ
x9KEX+n4Uf7wLqYT0wMgISoPJTcv6zqC5h1uR/OgvHD1OJrvtimqrJMHBdfRCqZZ
dYJhFVfqVdPC/6H3tqXkwfXZHr54WNkOJ9bGh0V1/kY6dh9UxBbfMQk8BxY2CYjX
0YzhwDyoKazs7RbMKbWsCvXoy+ZaeBWJvfw3LCJ3j7B0m7/4sxQBxmzNEN6KNMPN
zWPDrWExJUKJUtm2K/DPUbmZFPX7wzcdU2Nx019HGO3sy/V0j+cMTxRyQGZvLrZZ
L7xXgZLucgNNJGocdxzwmuJFa5WPjaJ23G/96/MzVjEaAeH5fa9vpNjwRlDHgfR6
8Driqr9J7vZ+8xzbyLTDoKPm3yhaFVyEvQSOUVMf18j74kX0pTD/B0JVE0Onjjqm
7ydSHbp9VnwKBEvB6N5UCilBcjSQJcfsRUxOfOtbieAzGFUGj4Hnf+2z3CokPn1Y
nfQgJrPopXyujW9pGJlmOAt6rRGIRiEsyE/Mx/WzYNnmgxaF6xCiGPJOrG9LkhFn
lbu/FmHgHSV+0CAxXmS5s88QVoiTtRqA3WOWbVEh/xcmr3QXsGkGmguLmu4Y3S3a
eXYSTxTdg7WH9M36c4qF4KJkAP8p1nbKhc6+XyhEmjkDIR6+e051tZGOthp7Husk
jZByypjUEFnmImF5hjKNLObQaoOYtntVYHRXcKZUqXy+mZXT2FIVg7sM4WNySv6I
FXXPYUuXkvI4vuaneqFfi53D3spN7+yTJAAJNWYtfP/uc4gZquizrwUQEP5a457K
G2cRbQdPgBsUuRqx1uzq4HWQD3kdcit6tNiK/AWKWO8g8XjN/QNA+xbZmLG0dbuB
Jmct5bQWwIYZP+cmbqWXuMeoeSwmLqpOtlV9YltSte2Wdn4yBsi5DOx8owFJLYw+
sApPCEdoWzfGUqTiZ/XYCxZFj+vYhR9A/HpXitBRhUpsEv2haA7zKI5B6wQ1VMDT
roKvzZKiAPQ48PIA2KgASe8oTZ+id+qh+TIyr/fIbcDkmLsWZeL8KEURMv/dci6c
T/wiB95y9+p/GETCr+Q4hWBF7J1foTN5fgqrE4kH9RXR4nkFYVCP72JBZq93i4Up
7Ekv7CNm0y5AvF/GnuYHlyKoI9Tp6XlitQs9EnTDsEiS0UWxJN3SpXlKJmPVj5UL
JGjU5JmNqal+oSHH7jVLTF3idAaD/kdT1SrY1VnfRWS0/cfCSCkmLyDarmkOlcuW
MtrB9rxlbTnZxhpFM98EwnE84lDMSLEqYB6nBSgHLI3Mt4LE1H1UmpHJQNClmauM
d15iwHGsk0em5a5Dwmaz9Npd3udNwvC6HKL8dG+XILOLDrcrzh9lSiTpF6WaQvNd
//FCjScbSat49YJXUu8FlSDvGTxCApfvyL2PoCoHhZ3Dg6VEdVjXSkiLXCVuOi+S
CTk3rjN8teKGtfA/tsB74HNSPnz5feK4YtLegwFhRKhKIS+jYk9AmVthWdy7xIRM
aqyqzZEpDUiUplqhevTGN8U6cTn3ihKTTChIZNW6JzqxCKVyb/kt/MVb7QvvaBoJ
qM2RjKYzecft/wLMQUIjGY8SsJw62I+bollpFWfIeCFIjfRcKPW4LwImYMklNJpG
ID4jEnte1QyKFrlJ6H/M0llh1dfbHVA3oFC29XKs2UESwAE8FGHgV8iVG9+ic6mB
LCZk6FfJ4xaPug00oSvTultq947Kl1MRGdzn91ffB3mxg+110WSJt8Q14GzWFZ7I
E/LU4l/ZcMTA2aR+49uwNZcLYm5C99oGOYtqZw4POkZAaUrqDBtJ/lRZfA/DIEwC
ZxAz03fW8D/wY9SJpCkEL49r812p3sPF/pZqt6Hy8UGhJ2/N8VhX7B59eqRCxpk6
CGzilHLS0+3S8A8fNvXCmYFg+na809wwvlxaY3CLaLjbUvWtVD4b+MwWTx1FjWkM
qaW291n1CNyz15dv995xiOQwhAccqnfOhisV7yuINAjWkcbQceQZ9c+c5zg8sW2R
aJnip9lkeWxV2wPoZb5IrIkpu+0YBeepnj9DFgq0Z70snI/7lt4yT57kmuHsuR+K
AduKP4lrwuWH4ems2Qr4yKNrpBqCwrOh8rSudNiNi21OvGRHtGDLXO6P8mgO1PiC
kTWh/d9acx4qv8E6eYbpz79/4zyIivfngRy5+6/KJ6hXt1I/0BYB/6jZVkCSVTcd
NU+TKw6SZ4u9x5E9Zm7d7huCWPmwJgngBhdOE/Fzl+UgoihnzuPD9tpkE+hXnIQ6
/pP1aFNgsD052xiN+oQlkD28X55DkqqJtX6+fUnrE9yWXqAKNgikCik5nSFx1xy5
Hm6DX49sPDIO1gtPCd4S+mLw4K453ftffNnLHJNZfYu/NX7trd0yGtaILCZFZqQV
dWJj5NRVLjX/nl1pAXiuvj2sWX/jYdBPc+fBRyrbS+W5BwaKAU21sqi0kSXDM8Ui
aXe6o1JdXmgSp6eaoBreUmFWn7uKXKHNNnwEP/pXQ9ImM5tzbgwvB/fcYDDC0XYV
6FZXpScI9CGVhnfIhMCGx/gyFFv3E/jVj5H+h4w5j4Zbzwj4q2Q9jFzaWGGAEIFH
51lcA30FKf/QUsMwPJB7tRaX5ZpseGtU0Q3AGy2Lokx6gtQP+EpzCO9ovsQwGvNQ
FU15VGZ2PN7SSRj3At+m/TQo6QZAm1+96kHYAgzyP0h4M90KqGgbk55dmbk/xTVG
jm986op65zKZQLYebGa0A64CrWOYVrEn0QRNSh67EaelEN9RztGdhXyOsxs4S8zG
9yNY/N0i2yTIi6a0MaWO2vJ8gAqWNsPLQipdZoPjdGvZoM1jvRAW5E7ICSo6aAuF
3NLlBGezHRpXeLJ0nss3yeufBoz5Aujxt0X/2ghR6OI+4DXEaEkFYSKJgdrQSPCT
vINpKY886LO/RyLD0y75FXdL1GXat1jI5Q/V0DVIKiv5wUwIPw5yVoWEp/Xi+d2v
ryZ/QU8Z/sHgSNn3xKrr0ub7+yeFNIINK8+Pe0Zij8x+9w2bGcGDn+8VIA/QhaBB
3iNfJUpRxzueptXyUJ5WASc3HLdLoUMrYAa2wLPn1PNSxs2ugXBYjLt4J/0euzFj
TpKgQl/fBsvZmTrNxGZbkqqbcam5RjXSA0HYMz4CNM6QlpGv0hLN8ZH4W3Ysge0i
dRT76llPKaeJfT1UvJF3j8QNO9RifZ+gt0aoLc6gOBILXVCouz/9w+NMyqKk7qAp
MWVy2Cbb3JFxmjd48T4yaRAhCbkvdIXgJtHW2zvULmZWMiRn1cG+sNOjg0bSD6gM
Ke2jt0QfGnjAcuux2fRuBXKfjQBOtsA0hrQAZEyGgRh5EmR0z+7qs7cYb/eQ8XdV
Ci7vjvjXnzuB0QJcAYcl9YSjBPKg72aHcuLiPg5t2ulZ7LuJpg4rwH4H/YlsZVhq
v9NzlTll+fRwk5vZY68ORVrZ3sEoEKpwzV9XhGMy3PjHza3qnYWk52qUBEPREWUd
TUQj3sNGp30ecHt0pZydUUUMNH/0USVzUKT7/zL0099bi0pI4H2EYsqHC/qZVFen
5IiE34JfhIIVUFwUcj507p/eNv3aNOlAV+Co/VsAERWTdABC3/BlbC+BctNSP0/V
hNkQUaAv2gAKGtrwDlwqimhy3LzZAfcZstBrPPNIq2im1bTK+OpUhJBGyDcNT1nG
jM5q2xvqchixhTZenTqcWB3ldcoTiFCx/BeRouWPELWgkzUfQntG6llWSNFAepFN
7BQYxq00jXqdH1hxngMeqqTo8DKjTvYkAIib1Wrl5gvA5tvb8kafeGtKuwLn9y6T
JKs4VF7pknpCHISj3RDwdeQe5Bc4vmtrFuBPRNPcM1oQ4VHDVEC+ohf9RtjYdqez
DkH7JQ44uZyLApemdXXl5OqSRhoRI01dTRwbBJf+eJeXENV8J9Rk2sGiLt0S0tf/
+uxyMotRXKLojtDHUMPgcqAl4Apid6kEeeyV5cgfcIyfGInD8uuZKZG1tIWKa96d
LJ+SomNLF1Ovz/jBBRtGhTsIQb+P7mIx32DhL4a4kz/XKADUPvHEkPEwm2fE0QHz
nnvU8O3XzOUEcVglpWs9d7f3a6shzQgWZwXKKVOlXdW2TKCnvCEoeHISJNTj6HDP
X37onVynIPfSX0WlU3Js5/icrTB8Ka9yypUHh8yZnwFaKNAKCEAKPaJ73XayvsaR
XrYmFVMg6URi4NPzUU2IUYqBdCwx43c4sMO2B+VG7wW/SlngDwkt9rgLRn1VctfH
GgrsGu/WG/z2oJFK7SYOzBODVrBOr1yzOgGqmCXj0fvqbsAO5rrDCWu5koCdUYSc
rRjyNmBr9uSYv4U49Ddsh6Ma2UNOj+AFw6DgYSDNoBworOKhUH3L2Z1Csuc8nipX
Nm0EZpZE9n9Z/Z6LB/IOLZuBZTFlLfM41jPGNhKrvaeqkR8lXsP8rRTQ60nUpSuF
Sn9gh1XHTOvOf3IU+XgmeiJH2K0VWcgRyyW7TYbfYV9zDi2nQST4z1yAeKq2PW9E
qGMb+I3ChuD77lVEtBbgHNynNO+I55j86WYsW1JVDFHw8laPREyHzVs6p6bZDBgF
EFA6+2gVxMGbTIqIT0bXKvASsg3FcElzJXfZj2kCCKfk7dvWYgD0g0D7nvAmYVxv
LnN7Lw4Xjs981hoQVr+fmUXYJQH/cPd+7iNr6OjF3iKXmJummTMJUElbshqFXTW+
qkmZP6YGcx7vEFEE8HyR3dFzfTGHuEheUDNg9nhkck1OHGbHTXtmlhuR3V4bj6mw
lgjr517QTpRCfo28zRTT266qWjug9wqKbByNMKWz9B/lpnUHwEGOr7J+Kdu8zl1r
JbGcZlHFyriwfSmN405dDb+hZuvGIoFzAX0v8E/3MUm+Po6NUSVxTsIg3jmsnvvb
QbcyNRDP7boH7gVtY9jRCh2hPTqmQOEMEjec0xzzaKofhyg9UlfzCrYtmI8RXvs5
IOcLwyDQx3FV6nJva+2lSqFY25bZolf0KhMXFSMHRD2RIY/pa+p5vdVA8PCao7s7
JoIerYzX/E8FrOmxOYZPA7dac9qAjnYF9uKyehzgSsxk6kDN8S6pDDrPeWYS3903
QjQsSTrdWlNrMHEzoNFzHvEiyj6QZ1JPT8UunvhwB9NuORAClPwT9UcbI7pheKj5
3z8Nx9G6L2v1KArTaNqOVv/xpNU+p7/WmIEMYe21nb9s0aIZwHdDg7496Yh8HLmf
RRGl3qaLY4DcM/wnxK0hnaK14M1iGk4/wxb42dV09kYvgdQNWdV/EbyjQMHYcwSH
5DWwE0Dt4n78ZA1pV38gnSFw1IfWGAnR03QCYt5j/FO3SnkhE4vbE/JFsBgRmZis
lA2ay8Y4EhfUmHb5DJaRFzECboe5QGCyyIJ0pK4qsG6rPbGefVDoX3+aoAt/20M/
q91E5umGNy+qvKtEQahbLHqjvA0pDDpop+iehHovZR7tV1ksIThAJDy0rMlvsIBO
XMTyCi2wh++3gUa6b/JNlwd83dGx8RfeW3Sy10lmQVlFpx54ZPrkPuxg4fW0E31y
H8fhQUqqjG85lUctaUtdRxGxxqGxVRC+yrzqNx9e1aPvUrTB88OWh6r6tQ9VYkPn
NMh8JqqjAK4RPn+6IPTdlvrtvsiDFAeDLImHxUZ12J00Jqye+Nq//vgSQBtEUHZm
HpNZ+xw0P2O60Ofkrzh2J/YY++gH39aT8BacoNoJWLlr+je5rsoH/vSVbcL2uGKb
DxL3uZKZIkRtARKiDfBF/NFfyIMGDnxy3/uvd1ETOYOBHulMIc9WWQBCWb3EysBx
bcsy/U7qA1P+gOStfEiEgqLQYzh0EJT7rPSC6j8qCsIEy5DyMlGOeuUT64nMZda8
05Z39jVwRqxoyd0QCshQYdklkhqUtdkfIDOWHw+JCE6DLLsl9tpY5sCH2k7byOH2
YjpiYTQpk2V9JhNR041Vt5I0e/MBVWw4INdJMs/WvV7wqx83SnwIok2NiVXRS/hZ
K27NkmawgcsdhIxd9ghWI5pWvYpGXeNot4IBJxI93uUQWCdmhhE2C2CLuaXdeG8O
oko7vGjuNciMkqObQcBpid/NeACp0/oGaotdjyob/uaZYL1WCAetwyxk1XVqYQ3E
1g3Yaxtb/7OuBRsQoMpvfYy/svFeZ031WynpcqyYZj/XhaxORdyLWDz620F83ZpA
EYyEoYtzYD/Mc7PuJtBGzwXvbQK+MOM4Yi59fXF6KHek529xDrikwCwNsCksTGIC
bAMbpXwL6AcJyrMLjh4Cw+j7hS+5bH2ts8kvoYvsF5z35wGH9XcumniuoZv85Ofu
+NgOUoERfqnRyWzo98d8GNcUDHqkghNIM+jKMVzp+VUzqgtwaolOBH0iC9SDFGVq
v0sPYh+40BL5bDxrbH8Xm/0/EoJNWdj9l6lvLltUr6Vh6oDTCNPDotNp36nVBzO7
v1pml6hqeEXj0YBZ5W5oK8Gp1doEA3DXPp/q/MlDWnIGOI8/CWI555BKYnsuJ/Dr
NEQ2nMHLiYP1OKQa79GpFsXzLGH7aQXvjI846E2MgzNk1OhBPP0aB1SJ0yJe9Vgb
NeRxx/a6NUqaXLtg90dqCfQcwC/YDp0iKv+CUB8CbpEclBUjW7fs0te5Y1qmCxGS
18R2dl79ZBTJAtLlUFKLZNxCMPy4PguIAkYhygyHqC5wEAdqYzkmtF+hWT9DyN55
O1/pcO/mIk2oozRYZ5NX8v0xgIyX3nyHUYPClO8LP+JyYV88KBnExNbJUlta4093
f8C+Fjbd2WCfzZ8JUDt0pqqW4DMBiqcws4mhD71GWvU2i+tCvhTxS5+Jed22Q5YK
Jw82w7R255NYZ3VRGtvRRhmSG3qm/iPwd2YUzfCLM2AxvuAtHziseGviX9/yns0r
RWom5IG9UyqbwSfQTM8ZMovKqYmxRJBbL+yt50WEy+NjbMORsI0tkUGdlFt307xE
MkXKIxdohd9LImzP6o2s7jmdNYvBupR/xROSJvjdZDuHdtxyNv3PGn++BAzv/+qu
7GpUw7uWj5Z2/F2RBknZxSQqiVWWtx9qwXPqHsfWeo6pkFUaxRJa9jnSTReSug/j
nefSt//MIIVTHh5JDsrUQ4ehxtSiarHRKdTeUouMUK0I9+0gZVB2XA/KbHJcg9F3
nfDpxzcOqMkhrg09mygLWXuY0nGgD5+mSxzmYMvZiZqIke4900DD05bIcMJKFIVY
XrLL0E2V5HZE2UaVHEcm3wP3PHhxy7lA0z5zV0Gt25dmLx8dVqvBtpHgH/o5FU+x
LD3N9xO979+u9onIFw4fEenoG8Q8BlWSGDfajXDqaI3A7uRGnzCNkS7J6CBwdohx
tymvw8lO97lLKpzp3IbyILSKOJmVgQ5GLQACSHx3DtmlP8ZeMPzgPkLAeZT3fDkm
4ljk32X9SrXbrkdxBpgMUOgjBaHljzabocYeamcJHzwU4xZgpxwBX60GP/7U/nJ6
EGevImsGrWoX2N1xCr6ohQ/5UZTlMwABPfpVDnjZ9td1PPXQZT+dG+yDQyz/4V8o
JcAVzD7kkvmAzvbTXkHhi04/Ja9y4coO9eqh/f1TErwraxv1Ci1TzLu9ln4sVdG7
o8LcoCNB6EDMogDR0YbYVm+yZ7mtOcLsdnLLgC/qJdBdxKtnT9p1Jz5SHdWMchbN
YXiXsKyRjvoJStgfuZcVhJXH+LC6WCsokZInP0G39K0kF5tT0l1dbTT7ReTNSD2J
9qby4lgBlpR18w6nswtYvDawENtLDlZuODUealsEdYxbptsK74b3GMolw8QUm9fS
qt4Qk0AgR7Zyis+I/Ddnk/X+kPjBDwDYEkY0KlRYkaxc22AFC/MvujoEnn/RPCw3
cPCajl+1xbnTVm+SBrHpIepf5+qHsDKCIP+CKLNWGcvteO6DJg/EHviF4ycFyIK9
djebaYY3ii6K4KDKpFHTQptrQduBgIeNunoWELlp6OS3EUZSP6E3tTttN9Hce4ko
aGJ+zFB24Qa2apXto/l7hfrgm2UIHB4t34iWssoWVn0M8xIlDU7NANgUS7eIwyo6
sic4JaQILO/0w2Ufljumg/2mCYUT6Ve3m1XVBvDQxNkZyOGCm8EE1aMbMc1bX6pL
GnAtTZSeuIgoq4SBdMQ+Xc6Cc+SlS+ttHg6R+DD6/3Iq9rsM3byfNAQcXHXPvWuW
ux4nCW18YUGZMh4DV0qt94yt43qG7Fav82zAlAXGaDpTw2VQPhVpmQwKRfyTIM5I
7bxf3O6w5Qc9DPXxAQMHHWxp/IXEnzqys7nsvCgRi8byM2ikau1dGPSVw64rm4in
g32yrdH2u+7/Gzn6kxU39LK8qe8Wry6Pxzp5V24iy+pR3bruVY5be+wPq3Q1lTqw
QCd6gdMWn5tqHMqQls9giiNEmJkrf+kLzLbVCDJfnANtA6g3LPz06MMtFGvLGnwM
V492xlQw4wM1GMqiq5RwgHCBuH24zKr41mHQLsGFIG0eG0YUp7zBOpyKlpyXbrgO
4nsXvyuc8T4DtEPk/QAw0PqDotDxiUEmcfwjCBivH9qdoMRt+ve/CfJU5PR2TrgG
y11d8+CSVICQknDCCpj7ww+V+NkUa/NubGXDm3cp1KWfYZE6U/iAHrN1T2f6zvCe
HiUn5CK6uL9M/iudfpgzGxyD+N8x679ryF1z9dEULybca3vwhg7TXitVzwT8jEO+
9KVbLuC8qS83EnZKSZvQ9JVZYm1HwIl2+yDzbSDw1Ys3iy4qupv/mDaqWqdHrV10
oewh6zIAlFEIudf5pO0WD9j4RcE54IgFVT8L9DMDD7erT0Yp0y0h61iK0j+7osTn
3Exqny9Fy86EK0O+w7q7Ch6d+d9jv3siCQFlrK4k7Onpa+DgxPyUo9vs0Y35N8ZL
VW6gCETLLYV93ElSy/5EqCCrRZtQISiqTvomgF90K0AKiZyatcOQznwwzVT3bdVe
djVXc3Z1xa5WnLm68dSe0Dd7nO5Rfkf1t0EK4LfjYbW+jBrfA9mIUvGJ/xJvOXlF
jS2cnbQedR86ZjNtcRYLllS8OUooRLpKrRmLNUX95n1bNXVYq7+9ZTYFQ2Q1sN7Q
oEc0T+ej2XhWP3OcY7GMh0B3iRsyNVjT9BNSJrW5NQZSZFuvFOy4YJJFvWmVKAVI
CDaIwrpBpkkRphoqV3l7SGykvumHhC4QD1LZ6b6OsQvy0DEKnO9fuRh6X5AONnRv
LdjCKwoWMGK2ptJ5U1gTuksYdbFUj232lTURwV1Laxiw7kdIBMTrJoJvpiisVADx
rS+OMmrPsv1MVFMOFMsOKtzCuM0FeEhZFBicpLXjr5tJeLEss/uvLCq0VYONiPRZ
76uykr6cW68bHYUuHwVlIV4P6jey+giITeH2zoFT1ckyjOqzE25l88Z9iCeK0VOd
QGX9BPA7nILrz3k5HAizQd7RFCH+IvzxHqXXW0I+oOtZq92oNM1Rl30R+Z9cZMha
QX5vV1I3Ie7j0yD3OUSHYPS9ZoQjBi3WD4eIVN3eXMfDVFdbklcI3uHtaXY3OU70
2/TOOS1E/YIWWMaBiV0U2DQmA86+h2t6wSCERZDBeIpVy32whnQhscEY/kf3JIY0
nvirBqBZiNL88q1vSVhlWTPnDyQc7bQadg5q6DrMgqGGnitOZf/0AxkvBe4hJYTc
Ix4IGf7qdyVBRs/65spIvZVPEqmNwQXp8/RpDCUJ+bx0dbUiSq5bRSZq6M5f0299
li/jg4Ku/dxC2yv4bUC3v/pEREFRLVuX5tqxvQ6p1uEdb/QP+V/npG0RzOnaGrjN
wJuNmGDu8mJZG2+97xaDg7PK11GseeJ25l+c+zz3Zc2x2R7X/k6vniFX2s4e9a7b
Y+kBcpNiswVBwiX1Ckw4r/xWxTCvUf+6im2tydWMbxNn2UUC2kl8JJbUWiIhf47+
c60uXEaufhtUvksqanGZnVBehx8Vzy6rPpRHLlM5FDYJO3boLAwiYPqXzM3mVus+
cjYj4Bc+wvWa/nfeDFaGbklN9WTV02Ow6HMA4VzV8X6mikgXpNuJpyoNNsI8kR3J
6EJ5iGP4X+OF0wQEj9fzC9p5W3hDLV6pC2Uc151lasuUgEnjJi3FVJsJbxMLqgFJ
YVw9dgObpp/xD6vGjb8uQQRKATybgmUiuUd/uTa3Mm7M5JB6404k7CbnJwV+ximQ
xB/DouPigmoqr6IaiY3JLfDG8DWQzs+xlt8sJfgPRvZ14TjeqKRPUraLuAwkEqih
+i5EUrpLrGsv9ElvvGgT88dw+27T5O4EjKsXRJXaY1y7ii6O/QbxJRCQ+afby718
xzxDBRuBHXQxcr5atE4Yi0yDZCmNUI1DZuMccdX3xQS15aKwmb1QlZNjme0ecr+f
KdqsTPso18HHDGuLcGq8FUTAPsmW5GCsE+D83M5vF3hFJ2HxkR0CmwBavqPnTYRX
44WE4tsaJNEUZ2vu9PnOAaUDvj5r+/l0bROkzIIW9JjmpLC36i2Bjg60SSHcvNFk
LktrZ+rJyKTTDhbvWBZbJF/8hSQygl6NUSJ6sKjzdWQGX+4BTLvzc5WwPMi4Iq/a
7s0u+FjAjqbhG/0dCfPWmwHq10cV+jg82kp7ge2+Eh72WeisgO3B84tNPtsywc7n
aMDcuZCYUD9fHUmMu/X457vydP8K6amHSxAiji/GszPHm7aPiapY72XIvv9A6Djm
dVEx6RM1KHTb2WlajLXKfv3EZBzVf1s4j7KPGmhXC/tXehHn2N5zBwhrvTT1nrsX
a87U+lX4NM2+qjtA1ziUvFNkGTe/0L1rp11MFxBb6fYVRbr9ft8yvZCCvM96R8vZ
Dt6bt/UswOdBh3BhJr8ky95cwraz5AAEvsOrjiqQsc0kMON0DbFspglhs7rQpyhf
63PNW605tdDr8RamQW18Oujc6vFyPSfaMlohx/yQ+vAdm0in5zG5OU6nalj29GQX
Jn6tGa66Erw1swsaNVobG7RfeRuNCU4xK1xHguNAvQhSWct1qX2Bs9ntNouhXtxv
Bei7VJtDkz1dXjM/GkZ8GTZ7dT5ENAGk3MXHaGtGaGRQE2c9VCRlY6cih1yT4FiU
70YvW+vbAOcyPdLWX0qqrcU3Zcj9fHsDn8U4owJHUN7AaWC+T1VsU0wDmhhFFlma
Ft8yULfkbG6h6yFLZZvk3RoN95GZ9tP/QYHhfErGZXj6AFuW4e4Y/1eZWH0QMExs
zUJ9bkBOKSvQ20sFfC/03u8qUp412OTFuiYSKCjRytoBASx4qk5oRHhVeqq25c+U
Wmfa4K4yqcDy1PiCDU0//mg6a8FmVB/vLw6hmQ0X9OzZ2PImR8th4JGXxtmxapKm
E7NnTpkLQZiA34ZyKkxRbaXLzr6yvpxpAF0ZstGKSnAdrBs2aIvUoe2qCU+JI5eZ
KIiFoikXyDNwz7Kjl63Aa2XMVKKun1y87I6BMniHjZpkb549y/L/N2Ft3bAcNOYt
9IPWXrosuT/f/eSg3ZSTAVT+51+PehX1V1PXtXIMH9ylWuDnDJerrYKs8XKlUFxr
ZvYczj6Ndw1d7eTkX2C7SGLqBZZVAKLRvNiaxSPh1IxIVEspdguDPbP6MLGdBeFu
D8F38UX8JinZvKkRS2Btg4ea9sTfTK0raJn0VunApsV/0SUiPvnMdOSC1/XjvHom
OHppXCQ+wpmp8kRzfoE+VhB7xzQ0PrMchdTcXKwJko3DQXQafRo48BJKHIZ42HTz
usG79yAfrZN7j55yB4xXdNlkeWagNWrFFetloGNrjt9twtBMBl4pNM5Pt0PTO3zS
0SXo5eDsWt5TU/QgArt45j+bzL/sC8qTZPYUg6uATUhT1AbxMG3CQPmrahVKpvbe
3U1pq7Yr7OUDCjzaz8bamP0pP2JXnPbRULEj09nVL6X1TsGxmx2uy1Osb7ToYIpI
bk2RO2NUi2eOK0gQmL2EL4JRIMgGAShALhxQdPH38mpmnyGqqFtkWJVZgVh2TqmZ
8ictwLUhBSULw1/pYtPJaWtGN2O+wWZwYmPHDK5D8sZfPDRJvikqy+nfRvcw+sP5
wDV8joDlfshjuPAN87lUhoqwTSbtSEurh2DWl06GnF8vScQ+RCW08w12YAIa9EyH
Mnp2R/RlHeu2lsrYDQjZ+3pcJncg34jHePus+ADENoBG7YX2VGmqREZC6gDXHCMY
i9QM40Rd0ktcfp6HIBZDcDBLr1GFQgZRGUhUK+zzz9tAiTdEF28ltD77LjKvbhfd
biLCGUUFbORy4jgfkBU3a2bOozMTwms7jngHPmBacjlahYEvkiVKA39CWtxGosqW
5Op6Wzlsxh5OtXw0P/7pejFLWvhk84BDR/xM5hychMCGkXTswOZlGpTz2q6bXKyA
gEfeQ8I7ghH+DxVhKERZ8LGCMI+x1BqLduiaoQM9to/xKvkrohV7jZ7IOVElEVTx
n+TA1bUR/WBmVZgGpjki1crjsSZo3S5iDHZWyRVLbAhLaXtU+idnydknJ4+jJ+yk
HXzrPQBG6a9PYOeqzQylSNqC4y/djVCPhwqfNd5HNiVuzmlPS2pFJzAZGMshiDQY
3B4EmhjO8gbPUlJjNDjv3e988OIZ7dZSjuQLQbpBIJTZqtXyts9Xqxk59AbVr9YC
AhZ8uV0dQ9kGMjSWeU8FniiJ3kH814MkdsgmvUKWn57vyqNne23vaR0X1mF87xpD
6tMglp9QEQ6sVvxqb64kKK6DBkHQOR/xa2US1mbELJSvV3dD4KNurY+bPIztoUwH
Bd393Eea7bGwT3JsUSTbPqzYoo2rjv1y2ito2bBi68Vxo46nBiAyQiY1LY62aPlT
1qU/AEvdI/RUh4OTULVFhr1H3KD7EXWGW+TvZX7oNj0szJVIORH66rbSzJ40Xy9P
ML9PkHjFbw3NB6iVJ3wuSSUrhnxoRZxW579E0SQZhRwSGMYSATZweWAYgUcALRZS
BlUBN0OmkC5CiRVXChp7BKspdnI+SQLnSu3AxTHR5/rIpYlNMeX8OH1dXVmKeQ+q
jQJ+SM+b2H9LYEKkntRTu6oXMZ+2GTITW5ar9hqwRRfW9vuonLT/25UgG+BbJLC2
XCECviUbtuKQ4VOG3obOah5Hc2X/bvryHJn29EDxuFbm1nxy2oA6PiUu/Sbe9V6r
lXcDHyumFDR/X4XpPNdF5iNKzyo2mJ05yS/lMEDgbR9U7vOsumLAbw33pytbK3g5
7vxlGZ82F2ZZI3UU4F5XVpghQ2ynKGpiNlaDtUiwbEyLAgaT4sUUsjIYoUHzWEyu
P2ORqxi75Gl6OCPsqDwGkdsd1JZtGkvUtGP8efH5mkN2UxKnPAzem+8ACdJpz0cB
dRsDRAeSZ7usWaSvOjv5g6R6eHlU57/NDSJ7P2qdnJUS8R8rxV+cN1k4t5MlVRdk
8Jd64y4Tlhbc3IKAwxfljH4fcSfTAdXQEUQYEXv9gcA5soIYBD1e9H/sriuco+O7
kSNOorkt9QdLuRNN8gC2PhWhtVIDWF8rLTyOH1YPfc6NrHHniFlWWk+GroawKLNf
0DAE5NRPD6WLbBYBiCMgKezZ7z6ZE/0T4kcAI6AFBIFQap5ddgNfFKAX40idX3uB
O6Xqmo1FFbham5HLDYTkn1Jmw7UItHWMJmTt8DWwDTVdmul2IeCC1uHuFGjvrqFG
y2Z5wV4tEvVul87vmOGatvHZeZI1McDYHiqeJ8DOrupEXFB5Tc+bSTz0eCYAYDu5
JO/+tpBzYdBWHzyQBBdWasoMlxV2NBoK5Szd6hKk/1HyKz26U7yU45wI9Au6Uq5X
02k92jtZolqT7obm5xo5B1yx6ryjw4pqD00dD5kEYCEH+PVQIxmRfibq2HpyTFX/
tFv/cTpPmkYB9IPwpBTlN9Ok0pVdVrvyzFbeAe0gXpLoRPIQPEAISIlHVKqAV+UL
oOtIkntHKAyLJLH03aPuEH/GF7KgAFWN2QhtQOOeoDC9w+tznkatdUTqrUmlD/LB
UegsODemgoXwQN90j/FJJ/BmOyE7RQ3eiVjNa5WpYgs1XZ5pWpHa0mpH1/jzG2jh
J3A38On6zfQo1d/gkQoy4f4eL2i2qQzQNXLTB+pvSikuUqsHZ12LTVC0TYIAyCoH
vG5Ym2Z4vMMWZSRVM2hMtBYZ+LPDUUmg3RpebUc7RvxOQrZzg72YtEuDzPbSx4+3
QtsRQ+j67+xLT8V/gsJ7TvOZcdY3f18HATsd9JaZJJ3uxvcV0bd98NcBNMlkt01D
oAyscYRlcGNdpHvbfR0IM8hFgGotsRtBUXTRUztMqAD3Hhw82mJ6AvcI+YlHzKNq
xRHoLPxij4mqXX2qev3WV2IYYlmXant1v0s3MqtjZ4Ui4mWXutVvhwfYazdJJXdV
tHvXvtF+GjztimuGuO7ueCc0rXle+CyqS3ngOA9MTEkg5lh9dF+KfhMYmj/6pd4u
jq7oBfTx+Qm5rDMqKf3v5qs2iL4HDuVQUPgZw3mg7yzsaJ+1RjlV1FQFkeFA9xDP
sM/+O5Mlf9cvi4QkZALOTXApKIuv0ncGVGzuN8J/Fudp/qaW9bSq+SzHhDkwvV/M
nCt07sBi/VcaR8A1peIvK/cceSQjmWNB5ZY4pNkuqmQKc8vrlfGJw02leoZJafB8
jRkCwn53+ykI0IWLGA6vcK2lNFBYQKdMucI//CH8k/t/MO1JjjXwmC/bjVdpCLE5
LUuZgP9kPwNXaDfAjwn0aPdLl1WPLQL0oGySffEo+vA/3uoHtgqSblxhsfMZ3o95
9eZoJDKUAuuh2nP84EUXUoEbx2D3O0Fh0qBKwN0CXr5vKCn/lHSwfHWT9bt+RT8e
DwaNYKxWx2c83KM4Dj/I3bEYyxZO5YwZkLCqKhX2PRsmbURaw4GV2cQjyrv3Nfpy
8tU5OrO3zXg0txsN5Y+f8kgzxmvi1QtI3HehQ7rqfzJzvfXW46Zvn4zjZp4zz4Pf
2MIf7/my8z9p9s4TCUGmqQ1ckxrCOq02+DqzjqSPK3/ice3XfQkFSjkmQTOxZuRN
PaUch5OUwaOyBRiePXkBEyRTqn2BkhkWDOlL29sVHtT54DJuGTNFFGuVf7Ds6l7m
m/0zSjX8fA8+liwt/SCzGQV5ZBjR+B96xs382bvxE4JvLCYh4B1lGBl5moToaizf
LpbxOtgBlPaGzwmh5d91WDyRvzl9w6s2gKAcEJGXXw8bWR8m+y7TcL7VM45LQUc7
HKdrpNQJOeZsk806rtVQNH3Ltzs0iQLtjsYKMW1Axx2Shlw0LOhaLjkLM3ngR2pN
+pOz6/8SXXL+3sARTPwiTAgUUVy4O4yCgzOtP8Z8SSmFOWqiebnMI64Q+Yf96ecw
xKCDMyLlZ6KH0VNAH1pLTpckOopfjGJDEun8qgLHikUTO1lgFJRbE3hiLmE6AqzM
/QJPoeRB1H+sjhLbTb0O/gntL+fq5so28arYDcaDD7ZzBl6iRI5SdkcRgKcgHjv7
g1nQqCQmaekt+0/LZmBhSRs6rtf3brevHvjCaxUgUSIh1wndKIBzYz7GkvQ4rYDr
iOX6G/WdaBCdIuxmx6DuSdDC69sZ9N1zDw1sSGp605nNXqpOCl3XVw3OIghPDocT
2pTfMgKZ/PADEfEhP1dDFukGWAjccMUp4MVjI8erreqygzgP2Y+vGOsHBvluvIoD
wV27pw6lcm7JHaL3Hx9GcxHXEyVX48W42J4OOlBCiwZZ9SjVx1OKJ+0zFYB4hzfz
DRBTatHfOK61XvEIjZ67OgCnR3cP95b48UrIg+nmasF8ZbJ3fpeMgh8rk2aedP/y
RdGQfQPNP/2N/HgSTy/avpACVG+9e/7CTpihv25XtYUHduYb0Y6Qlvk0kCUsksmk
wiR1G1Cvg4Ev+bBvRVYbLAsCgMhxB8lPIAD6RUjufqI+PpHAs8+VBx72YPMR0UYq
e+tnra5788MwDV9kiKccjGdLSAgxvsNbiNdloOqrhS3JMikCZTqUBXeaaLQFuREi
KJmN94Nj/Ssn0J4qYAAXWknHFLE26GqlvGaNFAjSm8aOCRaNBEpTTk8tPg7aP9p9
raCXwDb75qtC/FPF3jN7sr1r0LAdRlywnKNSqUt8f1b6ju76mh4k6PB8XfMa0TX5
8OboRHYE0iZFT9o/PUFM8vyokZERmnD3WfBGLb652OzdBp8P5VlmrDD3/bMdkxfg
Lkdos2zUUmsefy2gcSpJErz85Xqkmu/2qweouqyeWdoYiQvIaLsVmZv5XJR5gGuT
HaO45dBZBGqOemme+pC5hM+syrjevMLr96TTqOmLwABwx/DEoHOaGAMVsrXEu8+j
ViiJKulWn70rP03xtUikQArxC3sxKuMacbFeRrTyB6XlvqML2oAM3vE5Mo0QPf7U
3/yaYJL1Sw7AkGB6/9GRnWbkxfJzxIk/N3YGeEYQfR13kjb4Hb1mpgnT2+G/J3DW
nwL5MCVcpJze4UkurZC0Jt6vfCsoBH5oN2NZKZiYos+BUBmp4P+nY7QPmM9R4NWs
KZQGIjI/Meq51H4jvEQkwW6Pl+wQ2u9c1xkE1RQESlmUXBrcdbFy/dCYb7EettYR
4KZNtPGDqFiDalTR2PZQXhtt2eSWqz9qZIk70kJZIV1JHpXTAaZYBSdR7Zzporvj
6z9HmBvvLJ86yNsFA2RtShZ2And6dyYYpN2GL0yuFlmUYkhgy6n88VUkkU2yoNkL
iBQtcj6V7StME95mS7RprVUuzDNittwK1QgoILzuh0u3ZWqqgsWapD/pzIjkFOYx
spzVp2USq69lJZO4FLEiS7GNGsJn7DNKpC+mBflgdHXd3ZV4z2VSlvjOijD4Og6Q
iBWFcrrnyv5c8ZSZvrTlQJdinb86wabIqQH+n8fPVRsCSY1tWgg4eGyHX6iNt+/D
Zq8H8ro3uhGWtZklTH3x/sswSYFZqvBDdm16//7zKrhWoU6t8SNUbm1d9Z0aR2lp
dta2y6J609S5ewEAI5MqhWknx6BLLmjrMxKOI2VaLwtq3guRv1R6wgHkSCTXKOeQ
i1E+JhEyvspiDLOmuRKws8MYZaYf4SDmYqHAaisZ1x1qM2T837K3hia1bQdMdFPT
9SXlOQEhUFgiTs2pwakatXb267XZNtfOqVg1IfOljLlS4fuLx67t7PZ9w+KZSnX4
ndVfNhIcq3Tdk/UbEzdSCglKpruk7z4mtWomnQfMuTQXfjg2LzEjoNrSXFemZP2U
rxNMbEWaCIaE99iCqRFcEVKxjv2RdgCU+RS5TnxuTM/SSKg9NZhWBJ7wJbxYZdUX
Fu2AYZSX1L6gY02oz7JMfyqAz5ZIRGYS06H8r2wXLegPpB2Me72L8I0mNJSKXavN
2NQUEv+j+RsokEkL+JQJ1Pqh3CS5vfgcPBNyr/jc6TbYP/zVEYe4fSuRwPAA6MIn
sTyWw7WK6WmS6GVdtdhaN6hTLzyhlpii2PhPEGkivbkE7hI1N2a0Hy+tyefq7ybH
D5JeJbFQBselTNLeTc6R5C1sEg4YrrL7jBS9PC2nItvfG0/akZJrcCuXwGD+NyEI
nfGAGhJ00K5b47YkSB5uZxKWV+oJA5eqDNgagw8G3U6H6HkTrnA8yxxvwun1E8Zo
jhMwiGCiPq3zFoE5ThlSjCwsGVsYxz7RbBLlYArr5MM4wQVECxOaDgzD1IskglJz
U9Je7R2gfFYwFshubFZclmdIcAx4zFdXfuG8UWDLjTeRuyCdHdWcxFEWgQEXf3RM
dcHW3iZcWL1h0C7XZurGoYuC28X4RhwMkInGFrYTLlig9n3ryqI59f6IGHad2GUc
Kg0+GHFLHMG+j414r4IrQShQa9v6+zaoj7TVtsmKuzcTnoggJBh0jY3+5yGquR6G
NGOn+MXvZJd2W4+O+4qFVBRBpC7yeSgd97JUkTUijyhqHGduCdnfmOosaHaJEtyL
bdGXn020h25RIyJzEmD60uq1yKDxXDyxiV/fgL38TyOFs9Wq77wPa0rDeJ/q7zf6
ItwT8f3AyjR8vfwSzOEuB62SEdNC/M8Udz6XH0nouBZxc+km81KGhDYkn0WCkm+q
FGZkix5CoHilnjv/plihUPKV7R6MEyklhz+Yzf2glmDF59BId+k6PlluDbUUHyFF
WeLPD2nnPRo61iIuMfcaK2RW8PZU7a2aruenmX55BIn9+lbBpIqqeuX3L+H/7CUm
x9dzn408PS+jU/zl2qLtOgbKbozbUA0oUaEMQgSSvLXJk4HKpf/KKtl9gE+BEkJn
2+AQ3y8voi9NIdBBMTL4lPDItV+rYMgJC/nNw8bFhl4RhiLchv2VDh1jISFjiGyE
uil7x5DhDnqitPgTCRO893lDnhiVaTjRO1lKRi1BsDjQ4gNwuy31762QTmqa4rIh
Riwjs/drGfVjZKkXMNzmznYzRGzDuU87bpmEcebI8e1EB5VP3aY6btc2vXt72tTN
TAhj7A3BrEHC+IN0L+btMshAIOu7pS68UYvD6iYBm9/W/N23W9SxMotR0A4VbUTY
GWIT4WmhcVrO+NbUq7q49U7JcP803020mt7Z6nysbpTpZPzghEcWrcX0qTPOfThY
ENev3Z90C8KoO1rKQO9adzM8Z8V6jlUZltHI9EPk7y83u3LwyYrn/M431NjuRyuP
lqNCVHAkp0NaQ3zJ2KU6hZ/iLUxT6PaCDC73PQMTPi71pB+28uxl8TMw/DaLVTsX
wGYZkvI6Krt/O2Uym7FOKdrNC9IuJo/CdmipwbgWx1m7zbbDB0Txh5b/V9W1vohx
49BqFV+Ka6IRIxGAtQ7h1zO5IhDa3A9L99K5h8I/eLgh73sgKBxdYBck2CNkMXxy
KV4Qqtn8cltw+85RItHgdCGrJgxWQU5qYhW22Fz3HB2nDxHN9xG4wMTwzhCK6c6j
uEANb4SElGdcD/Hwny6lCGmQbra3RQbCOr/iJAfovN4eqKfw6POwx+Dw/TAPZpQs
HA6hMhfTP/k/7dFVumzfXXuyFFQUudsu6JfXzYbtN3EPdE3X25TOK1Ms2NjTBLp3
0spsbJ7pdHaPlyZ6ktFN6sU089dqO6UzKI/sVmryUS3PX+z1ca71feIVezC0LkFD
qmqECd1K1STKNBDfLCIeCIHVAoJNlEGyrH0tsAdWDBq4t41BiX4us7Giqg0dG9oe
4ke5wwoO7Q9NzICt+Q0ZEe5IYghBIGt022FLX+aSbgcJu41dlmOfzvPfQXxIpWQc
TT1wFIaZG+tRI+jM8b7R5ihScxM0jn6hR6BB+3/lSIVIm5CQKLB/wrTS/7YGkea6
+IU98q6WZMQMBgmFbFkcQBFLRL+XimRpaNHGNjkJSTKDHLdp2O9BdnWcVqZawKOI
ZrxNZg54qtHvzl4XiB98H1IP8DrMKV0RY06nIgFv8XnsvBN/USlXVw7ivqzoLpsb
fn+w+lU3ZXdr4sX/9wlSrX5kamhwS6fIem/goP9Afs9tNQ3e3QjvT69OkwVfeuPD
WhqjV9j+Rt7++w8HtOS/WBEJFrPQPGZIEap9fd2F3zN+EpiCvdVdlvh2t94B3ZKy
mT5kY6sPW4vZ6e0k7nIR83lIVsRwmAojwaAJG5rqvhpGumL4iCbdVmmJZ1ygsr+d
O5eg20Mck9T09xRP7UZtjL1keKEXS2ryZyVtx0zUuTSxPH/3DKFvGj5/zjv+3sVU
XgWvXDsz5erX5MmHqk7r7JMIAGmEqzQMbMck7kxmdALfoZKauSh/9PTFN8jWKmyy
udemgu1M2DvtlDiBghV0IvdXA787wgkAttcbsYu3WcE1TMxOTZmCmhutiGq8IXEX
9Lmjr5eFcUD8eQ3CiQ9tAeYLQCKbkoH8+5G1pa2HpCdig7fBopqgjD/T/PPVB5u1
QFo41CFDpaLkK1vtKfnaSEy/a/X8zmyBek8kCqL6eR3ETUGKMKFlgbvabeZpBphy
Y86meGJIriTsLBEmjbKw4lY0L4Gde4oT0oNf7m3TsMai94BA5dX8kNoQHIYMaVAr
NVwySVaiO7EGCI3NsdaPaeZoSE6PbLxAM5t215syZpjrZ8cSIG/dQy7ZivhDAwtd
kIjFfhClsgetKiTb8VetG5zGIccIycu2VtQK7PEupj779FxTAJF19yjJJmGvETL+
R61f5vyscb41fMI96ksG80Dh/LdWsyDIZ8LY4KS/Y2d9EqPGGBUk3fBmIrAut2Ss
KCBVltqMXI9S0N4BCH0ivZEMxwELRbikJmPPTIiPsg5m4OJabc3OjEDjh6BntbTx
aCR9Fe4O0jw6Sn6pQml8rpKCF9QuxFx1gh6S1o5a4nHCuH+FWu4VC3RT6ECVlhHZ
q6WhORh0HyOEdaXLlYWtQXr1iGmvmcHU5U9C3AcFJ+4iEOXIy1fVobVEqCx0Qcbo
1dZnxY0OPAkqz9MLgnJyNboxGIZfNJ//lVCNvvFtdKiN8aYFAoetXeS+350g1ZG1
/rI0QBSg05Iv/gWTC+9X3cZWvEHXlMvGuwbFr5Xty4gUU7nflzzoOwnZ/B5G9nq5
hXlqZv24CEeLBqR+8qyRlvXVd3stlKMCD/1e1X5r7OCFisNv6wBrdkuAX9N4fIyR
jwvimt5dbkYrmskh+y6+4fv5wmAt9xfwytRZvuXhdhCQfFuAbCTemW2xTZa4rdom
0seUHOztO/OGZOZ81OMNBEx+1o68t58hnIhe/Ut8f1LYvUPJioPdHsyQh6rtn7ib
2qja5BlitFzJETpKsFFNfunf9kWSrcZl3mgq6Gpo1E8tpz4V6myPHdrI/o9LkxcV
XyHOsXOd6eeWoZFkjw3/Z9dCZreUccAVHM/bDgJIX7xzQllEhn9J7SkHQBWd3nJF
zL39fnFVF0gJ1zeOEME8u0pp4h0CTkJ3p1sjkIxrvsuxkV5j7Ui9qmztd5pCGavv
mYPTFH82koViIisaJoPo2RKw3UFIIgM0XRU8+OUMddxglt+b+BzvqYNxxjFxcU2c
jRs0HrzeuqBR/THAdqB9PhBfe6AM5dUZWf3myWIwTBT/SrTabBs1sdrfzq7ko1gC
3QrVZwGQQUo/9lheVa+9cIwQmA4jMhv6CP4uUfh3zKSeHoaFRbqf1o3DAnHL40dF
8ca4Ug01kDl+o+NE2QR+JCcVtYwRZNqFbVrdVTbtHxJRtyVBdhWhrqE56JED0A+Q
7rc+h/Qkh0ubirpAXi4+IE4mRgI6U2F751+X7kaFDMpIwV+uFbyVwfbSsr76/SEk
oEypW01YiJxZhlj7E+uUAipQfnOHA3MXjw5dJt88ySEzgcQJxePOxWvzCmfLGQbD
B2oFvtuotL4gMLcNVZr2ypjRTBLLPrU9kojewR7ptKFrqKEzgLYZS/Xw4xO/NWn0
NIVKYWg0DXpGjSv/wpsRU1/fsmnPvu/VShoJp6/QMag3eYn3k9oCEJdKIoTMAQDY
zERpXyATtbRJQdAjhsNAsGR5OGUPB+beelcXUPfofC4TaNfLowFrO1Twhirvu8y+
tm+/VnFoYdFugmmX42ujCz04GbJngg6j9IjaQcT9xERNA/HDUWBTj84fu2KYCeDd
5Vwf5fVLz8xqayfJlhN6Pd7eyASg28J541or6ReXq+Xurdvcedxq+a5MHtKIwa1l
awMa8WzCaP2cxDQizNOpWdiliwg7K/b0hnwQDYYw/GUttZIaz6L3k1GsBtWiPhNh
WI1Xdcvq7k6JzxF5s8UgxpgU1zYM4Mf7OS2Hy2dxugwsL/jL/waBJ+oohKK1Zf2k
6O1bFq+l7KB7XpcC+IkpndUWDFAjSe1XlLbqz378LBuLo2NsvrOSZ27ytKnbQQWJ
qFekvKm2fxNtssW2ikopowoap9ayGLCg+Jh0GMkKrVkgGdGyEGQ8I00U2rO3U9Qf
2ra4ShuRSjChx3+XbSv/8osv2Nb7mFvbwhr5cJ4L6hHE8zvfV1L1AgCr7yCofyGs
K88SR+fftq0hr4xVtVixKzaB+WYnLsTNfF5zCpn6cYbwTb6Uza8i7BrAS6Cd+4gr
9l32kS9rb9WsJ2orqAJ0+yicywpZtCe7m76cDTDKSkPfwMLVNUgyL/jDYVrXfKpK
2EieX6WgAtgDhquYoTjdcy06pyPNOxwCV46s0J7k6OhnFXdQ33Yz9FxPWSc9hhYn
vYcuxq82bO9lalidYJKk6uFuf/accEF3694jaxBUgBU3EbcQXzCqyccwGnucYCR1
9riuc9r83/hy6HRRE8n0Sxd09AOGtvSyz+tXYXNypYoeEbhpjzT5f3PZJRb/3mg5
rWcC5bhMZvGE+JuPcCX5WTlikMY+TsPFsHzfpUx9XwkMkHfTCOfe0GxVAFnllFFS
BtCeiPWDiNawxs5KypxDnGOG20hcWTM34w+EUrym1clEb3XicjOc6n3e8jt/PBPd
RSXAc4BdHq54jbb5oxFEGt2BYMuYImnF2ZFOp4jIr/fQi4xe2huNQuyanikUauuE
ZU3kz32Xn/t3ivYy/dY+RpI+1fcY9X/eYfxh2ySxpyNExeXIuGQi8R+BVS21+ufa
Lq3OWNdD6WUCUyD69M3Yuos3OBgu/81G6E2g2RsrDS5WGT5sIu680VyY/eSeGR+4
OPNvkn95l02rVMmxOzNovfKFo14g5KeJGGeP5cGr7+JPQ2JbcyXNt9RjbsC5630G
7MjftaSNysvOl/L9AUkJNyN3Tyqduk/bYG49IFbW3cwa1UHSlBpLSF15Ye7XlEc+
yuiqriurXy2XzzVVcKJIXUfTnwsC1IU9Q0pxAr8VOgmcZaFsw3V+FO+E/uw30Bss
2K9i9SaqF2XyFoiEURvgYvpNtwTTy48DtdVZI6XyjwotOcD1cYgN7+WmlwKpc7/z
4boQ/B2c4PW1HoLDOECvO1lns/B1PMPfFWebVUnlsOS+5LSP9FUc1veA8LTg316s
xUb9JZx1ZTvj4buRswEumTjhAS0pD2/jXpEF5fnOZd3CXdHegk+OSIzZeMsCMO12
fj4Dw2putRpIISxWtjPGviPK8hP+UkOpJT34iRRpczFSuep9wTzeWCs4pkGi74Tu
/cg4dAFOgPqnHqlvjDxYTUFs34oVH2pFiQJa1CKEmDw77BkR6RgCwF9BdC/pYvIu
jlObjLfkYklZ3NeuGsBvapps8dB1rcoDlnlntGIFdjMyzXSTqNOfVKqQShU2U8hn
uNjEF5PAGQUPIxlntiiSeJ+TRyJYlIizID+fhjpPEi0MSJpWGGB0qBLVCM6b9lc2
jQFnhtPaYmEoGVRIHaY0HzKy57BjQLSF7xHVYW/ar04GyzarHvUYTZnIFIODGAZu
8Ig/U30vYR6BDFKWBBKAkobNVTB+eh4z+FLHElwkAJrVIUdmlyZ0XOLaplHIuUpz
3vgCG0DSqY/EnUkj1qLC8LZo1gGBiIygTEMev5lvpcT31qzdwEwkoaXSFrm4cewD
5K96WI0d8BVIjotp3zKShcMMIl8s2deF5q1Tkv+wohLKU+1ZxKQQ+vZrKBxFdZTf
kD1vydE2vqG4Dfyg70xuOY7qc0/wiSxveRqPP6m7HWED8GUkvr82PE+lMeM+ViiK
8UcDwRiiFNMXPBfCwTm/xXUbysznhGBZzzI8MSKvIkVskvj4RzRopsbyk+XLrWLS
Y+ChfaGi6qLiAvT8R1QRXPLJ+coNZ5fXcJr0ABfokCndMMck04yNFw58bzqZEwjv
myhOvKqJo3IhMkHlLUmj1p6L5zF2Z1Y8dluXmPHmmgnUp0+cmOs09Q/u24nsPzKx
ZSvqwT0luAcgjmexE2MxYlANRj7e6mq1zND6aejceI1HWiw2FWaEBD2ms8o5ToYq
nlKqO9HzwaPPFJH9LrLSE07wXOjh1UpNBOTZ/ch1F/UGbtFfodQeMHk4mGLEW512
E6RJpXu1FSOIELCs5H8XBpNDuK+3e3oknpu3voZZryf2R8y8ijfXQ5CjuC3n0AB2
uz08t/+jjvVlFnkJ9381+gvM7Ik0bUt6bGqHwtOilOI6AcnTMNf+5kYieKzdUpti
fg267ZaHeyO1QgWtiPH43iqQ2ORxaM2q0nkwQ69DKHC4paoaZqsHXe1r+Uw8QYLS
VNvMzk5pJVhPCkgMGtgH9EejayzbNtOBzsKt011P5w20yMNaiiIUt68DJsXSB68Y
Fv938qs4TDkzBsNOHq1FokUmfDaGsLBGLF3mF6OsRWB8C5AboLCLfnjkw7wljsai
G1tZm/Cb+5VzZOzDngH5ClNIBLk0a4iyJXga1NYD+/4vc4Tq+MOyNmWilE7MTxGq
7KGJWBMQ3992ABc2Fjs7osSWtChd+MNlTk9OG6JLNkjvo0mCFUJCXF7l6b6EB47m
vTtxHzI44rlZ02Vbr+5+Ddm7NVFdUPX/Il7ao1+SE8qMBwbH4Ol8uwAnpyp5kfg/
XltT3w4OM72ZX1fWCT+ujswBll3UP3TpLg4Kcj919TNPED3ICUgxw8GxBezg8rvb
VoovoGOSsRLTEJJU38811QIprzV68Hi4gP2aoRWG613DMfMwBUe7welzPOcpHMOs
/3JRM3q15AFEpcf16p1W583i4FfGSezITCHVC4GgC6xaFzYKCWUnFDR71vggHOXh
bY5XqXSlh0gCP+dEelerjZJTeH7l+upfFM6xwn3DxiQdySmevCi6MFJ+MI7rzOk3
uzgS3dF4tpH7qJnixS/50Q26sYE8hl3I/FFC1JQW46OLu7GRPLC7b26cqNPSrORg
7t6BICilvzlJ7ak/uraFGXs+RJ/psFtSscQyKi3oSXkfhZgb1jXV17gX0eN48Uup
Rf8wnGtQhvNpgWwYKaJusSc2w3spK2iUBvTlcYkv0tUntV+95vCftFk8C8zi6a5t
2Nv4hYXHdxpT67SuqjLJIH1WTJn/Iil3wuzROVPA47dFpwftYii07M3S9i5VHgRj
YJNJM5J50ihZdZAIe041EnIVmov1VDSxUTtzr5jxpVo7WFj2yLT8SBXeDLoQWZCZ
Omppa24JRaUo3eAVwMM/x1BQmXGV8JR9dM8TNRj0i5nBqIbun+9qMT3VPLLoLq0G
qAujnZwZnhfQt+qL23L1VypsoRwsQZ2zigt5MWcs7CMTc5lO1FcQCoTcYp0wFmQt
Q24c/Ktlg9wYbXEJxlOhWndATTVboLeIgE5hmxA983Fg39Q6IMwjTqZ2qHKeBDn+
YeUJISWZg41PpRuNGFm2EyOilbY11bJ961xvWixqCU6+M9+RByL+Ay+mCYTw10cn
IlORZ6z/Ww6wsiHTmjugeDEyh8vzlSp2CHvK/00a7zJH1/y8FzTD/jazF7JHAq+F
8L0DLv6tPRaFs+1KK+59GDtVCHQ5OGIsdADP+dbo0xP5T3QjZoUlUicaQW9kIXl7
o63Gkx5pKZCvZiIjSWADoftWqB+bZzL9LV0Kvm/LnaDWtUEx/86Ta5i5USgJt+D3
zOZd7Upjp7AKxJOhOYPWaPWGXbz9l7C/iZC3oDSX3uc4Squor9g17yilJOP31WwA
yOEBp0edaeHsP3JXa/BorTEUr/Q0HDpB00XY5jphtn8POHOI+CiSKcprfXX/KKjE
V5McYWh+EoBc/MevIrZZKYa/PP8WyD83D7YNa2YRuVv1OyArD3fjAD6PPrTyvc7X
78Rj5O2Bx+HORxPuI8JHK2ek7VCktn8WCEKiK1iQatBxuk51F+3dCbNhLP5/5vf0
R5EGfiRXiS4VAPgDtTG7vn1OUvaMI0bVrZcjr7QCy0+KRj+QbSIB1AEX8Lcq7Xx0
XUdtjS9al4T8W+dcpPWrgsnpZx6tUK89qUVReG0Troq+HUKVDZ6NToRvUKK/G2C5
YmZGL0DyBQWeBP8nRzbNPffk4+rHcfeyn4eU8PsmdHEWIWGwHxdGFSCcFyvQGgb3
dh92XplIsXeNLbnXvy2ZT+eiknWUz9/LoYTsSyCz05WVnHcMsv9QZMQ6G2Y7QTiq
l0cqirLgcjt/FDo7/mUdZrXHzAq/lXS3p8Stb+xCJHI1qt+n28us3zGMyxEPVa2h
7NLDO+SQaouEuWhrvq4zD8cthQDFiTO8VsWbPDWBEMDdpu19QbWqXn8NecNL/DgS
aMs6Mg7aRiQIlPozjrLDitwulOfOS5kt10sYE6QQWCBCwbYIIYSY4Aj3mFpa6vbu
/3GOzA/HrErYh42EMVqXEUx458tL3tlVjkem25w2C5bOgYfrHt8OIpj+GbwjBJR+
OwmKS1Lj+zW6+4vCVbLcWa1mKWxgZdnjFq+vzSaY4iENrHieqvB6jYIseMmO2Fmo
nmClC9X15AwTtgkCJ/Mv5nuTBfdpWHYyZeuS2Irb9Sk7rfrCS77WDhcCv6oJg6R3
r62taI7yt86RVCQvt/BsYkwCRX6oUdbv0JkE8ECXb/5bFwGThhsqQoBHiSFI17AL
PgmPdRxjj2vVD00AY0PKLpyYfnq4Hm11ZxLAeVQfjcrBFOVXiySZGXI68/YuL2k8
/S4lql5Evq74RPJvHq07mYoyrMVQskRuOpw2nRFU/9js8sY0rwYcOVBsPhUnrosX
L+GLnrIjae2NOB8skdrlJ5PILbZEjZKRxZ8zmGhAOW6um0pxkYfrEn/VWVGeg/01
SwsjNwKQ7D+IL0OkafTL9vIP7INlwR2XjwyfVX14imjLuHG911u9S7yElwEx0u6v
C1i4/hqCb0iN5BzjafNABTHoNpYqPxLmrHMzrgBJS5cfD8ax+40sadg/FKVN7b74
jSnFjsxaR9MBzarnR1mNoYfNEK00o5NTTAH9Zt2fUI2QgaDEsCN8u1WtgIxMn71o
FjlMw9LJ158McBdQ9VZqCtv+7Pi+Li2u8J9jx8h2LaW8B1ggXgToL6sd/JzDSG96
OhE8dgyducm4BJrhsAS8UAUMZ5W/V3yLSEVY11T75xjTKxPbr/J0eb23Amu5WErc
cLh5erjHFv5hj0OyHhBWUglksuUWyr9/TOYbzfySrx0ADCkoYnhAD0UTDSdFRqHu
r4FgEChZbDPYmZFnHljnlQJWZyUF04t95AMf8GWh3fMrA21q1ytUY1rLg70Im5aU
+KgnpJ8KGQZDJf0qj9nRmED13QpHnfmLJ1lJC6QrOSYNwAI7ZX82BOS/VqREnlKT
JMGQ/cbQAB52oHqdC0ZT3UbmJ73Jzxot+gT8z+hf51FYtGbyXco2LfyXUXlQazxP
3GEFxtbkdKlNCQjoWAUOAoIq2s/CEKdwayRDL9w+q1JGMakS9B9kdn/4CK1qSNRx
Z/OS88CtH9i5kVmViD2RdvKWEkVm4Po1o/zDPb/GpUqiJkhC6Bcy5rZYpjXfHTcB
R+yNCa0X9+AGxTKJMdDz+nIUCLjsTaEl1dRX/X1XMTzPD4cvrrPQgb6/w/4o1G8w
5LEn7JAVo41uUI5CchynDa58IzqP04vT3XCxJB9YM2HooCjkP6YGRbfAC/DH/zwZ
jSZiMqKrfLA93S7P1RuRWhlH2/BWjLUbRjks4pYRDcjb6DliJlKS3H5283Uya3Wc
7PE9P6EO0W8Y4pEb/fJhkss3nWaRo7ZAQMbaVhYULnkDlMkEpGWnEbJ3vsEQTRmF
Qw/77sgTn9o0vVjA/jw2eC3AKOsG3kNc1qE+FJfxcVybV1/k1o3PiedY0Mn5IA0r
rTqX/iIv/n3N8GbAAT+5zWlDyHy4wULikG73e8VfigEXknlRzT1zXrhGl1nInZZ7
HIUjAD/YY6q4W0vqrw0cbhcFxmbVhuxZBUqq7LMDNjfsUWu0wOBvYpjTdkKCQkxk
bvGJZIkjVQqXzch3MHFdatFO8YK3F8GKr1ZomWVaR6qLsx8CTU3QvdBa7hgfkviT
UmuxpzwW/fTShykh3Varkce+MqZ2j2uHShl51DHUHmoBLykf0ECeBgUQSHN+w+mL
vkDGHvDiH+/DPQhahb5H9iLtKfJHgguuBRvSL/sNW1bqY+BWgN+tWflYe0jHsHcc
yspegI9gxUWvsWS+8TfZVj9vOluqJr67XRJ60Pq/DAadvpD1VOtopEXt0IYit8Rv
Bz/zoLLc8fRev91WHXEqnFvO/7XMEbuJkC31VnbAAkFe1OB+cixzJmmaM0b+aNYP
O/4erftMMQJF+bbhSctUixrvHPVQ4/jN4yK2iEmTWKMRgzNbZsMbTG2av/ubVel5
kwtXyRzcgfX4wCnnw9RLPihhXdlRea7/WuzXUcrGXEbGT/VDQsL2BU8K4ol58wKf
FfbUOHtXHCxCnAgU6a4NW+9cMLEgFrlW//jMjlMNSwHN7+r+hU/XfHJqTUzV9L+0
6AXN4l6IPabiNaW2/90GtniQKQ6bZgFT6QKenhjowHQEe1In/dJWOVKbu/k3v77H
2gI+m/iZ0fX06ORh8f/Fodo0JqZiDBu17d0LI6LpTJuQbZpDHilhJ6adnILqdrf6
8rSU1xCjDvMJL26aLle5PYkaVEXMT8sAq4EAsbmAfh9wD6BKbRRn8Wy/GI7QIBDF
1haFcm7I5I+/hTRjyqfnyn3842tsnz1LEVnorTTUS4IcXXebv0ifDiik8mhDuO3k
2gJC/zuzbkYDOElyLSfi0hbV/9PtpRmDaVehh53PMvA4SV+NtETDTZjqpTYH93yt
HpXGGPEHJhpYIOPxqYRyKWSFQvfn2RUicC446o4U2OFV45877qWBWDqo0g2iGvcM
pTnw7j+34udmeLorBMK2e4dR0OsPdiZDGzjPj4uE07aL14Bibvl3MjcQEBo7ocKb
I/hEjH3CQsz5Ygk4xfxPzC2Pp3TUroEIQ/dyJ/uqIXIkhil7ofPvDK8TcPSIuRpK
P3aRZm9oWILklFF9JoA6sABPWnlJOvW+vGbtS0IO5yZyHv6huOR2mO6JPDOoQ5uT
ooeJjZaMjjxHrMK5LwpstatXkfRiChNWGGAk8Fx3nTJDIXmGe6vTkBEHKZOXYZXZ
COM4g+miDkQ73YfE35VdemX2FsciQqViGI7K5vKS9EY2bjxCFaVaw2mjFMFLGMG0
+M6VJXcOQulP5ZsJJSe2n9HDUHj5V/LUqpjhGnJ+AJTtxuA9LqJmnv1ErttwTLLc
/8bjXDB2WolpQE5UUwR+9s1psKmhfu3d84EC/2zHv5ryEtjvsJZw7q5we/ywrjif
yMdhdlnfKaZCqgqFnQ5m8AAo2GTWfGFkuXEDbN5eth/iSONmTZNXl34wkRs0M61C
YudClXvC1qqV2wvO4oO6Ew7tN88/g/AcqE29UXJGepEmdUvFcbs80sjMs47q4OWF
GZpRo3PM6kQlJSNV42vrBnKwTwqFGa6y3c5b2hQWaEYdIaR0daxEEN50hB5b3NNy
TeozfubFsG4KPCc6kAL/Az/OGrqvoMpZmn0ygCwx0gul34JHgm/C2prshlFmCp/N
kkVNBonMzAFBgjGHFoDcvFlWDYNt73WfypyiWtO+J5YtK1YPxq56GzZWcDPDyjaW
hCBEzho0QLYCXPR9ri7AvcnnIcF6kgXNS/JLFwuz0MwzPJjUV2b0lul0UQMrg5AI
F4lejU1iuKHhPclgxsLZeII/wLWbhvkjy6R/4DoXYrlB6m12Q7YSHGsu9UhDQygm
5x84umpXJfitkeCmuT2xUEkbPeTMbEqN/rkXDm62JP5Taz4fzyHUaMv/mFNBIUHK
2m6XZZu0YRyHuRL68u4auGrEhDKXbaUl5GhTsH8nlEw7nXeF6M001vEAm2yzMoxR
F2UFxB3BJj3s0ijRdKAIPaXmYGvlzFBR/qQ7+rPv7UToZtWn3EpSeJWDKL3X+4Ef
0/cS9Xtt2Y3f1Z4gNeRG4wW7Q2hJ+CVxUrafx1QFGPpLlrsiqhXOcKk5qlYr+5Ad
ZlXE4Lz9a7/0PVD7HtCD4sR/gXzylASWs7rqW+HoPb2oZvgzPAa0ktXBYLH9SneG
GMFXOs7qgZ6VI2RMU/rjH19wI0KIQxW4uHAwDMPj8FCdc9OzlDzWqANdvb3ipGMl
n/R4ZnnuUVYlhoA2HvgQl1ZstXtz2BAfKnpIXcYJuPdfKW8kE2Oq14XE9Qo/Nwmo
HfYk0md7LKJ0ixZSFGF6i+pi5H/4S4+JTtYEjvE31soKZm/JpBld4oH4aD+CLWAV
M+4FONJB2yN0qsbzRKoWSZs25BPXQr7/rsuRiL9ohvEbnVf824YU4BiVShDq9vVS
r3h/P/YQ1m8TQT31WhkvlvWPJAXg+2zzPVgLuAw4+VJ908QJiLjAayqmWPEYhELS
PZ6MDzSt/d2fTv9EGD7Vfes9mA8z2Mz5/Au/AVUCNhJCuxY58kH9e4XH7jX2sJPt
evyih2+U/UPLaBkSCZ9HT5m3N7DsSjGG/5i3wuxLOK3gGj1VLuYcYu5vxtqJl5WM
KHGWBsY82KB/K1CgM1b/bakFHJzBWfoMTIuN29SlWYPK7H8HUmiEbxhgrCl9DfX2
r3pUdqTpi/HXjYaRYfF1zpnfmGE4zDjs1rMFMbSCGqUYBVFV7uDVd7VOqhlJUT0I
l6S9Tk1cn18pUJdQDSZgTosx0ERQvnoCjCiqU8Z9ySz7ihJhP6dm6aH1cEZtLTei
p3bsdReW087QlnHDPN8W2iwgAXV0uFMBrP9qI0oeReghE1ID7wbZDIhjPkmJmTSY
uJVb9aAigGuF5z48AiulHjoPWCsgqziOl8T4iHD2AP/sZS9z+rjZdQGyi0CqR4kl
UQqA9sfOCzW3yN2jU3DpGWql+db8OerX+1pZCo4I7EUG4sFsgrRdP5Bmvl5Cd2Kr
l+gQc1xYQpJWuaS5SvogfG2aZuk7enzhRTaoVOR921SfhknTP6LIT79KmNTEfz0Z
MCnCbGSkmsX6Fm8I3J/ZrT3YI4fPUdtw6FY/7wjoKSHRBasZOxHRJEET3I47Yap1
G2iqy0wBr/aiE4cyE4PuRzmM2tR0zzHCujrsQEhY8ElD+uQXOiMCdSxmQusOwGJ9
du0bvvqAvMIlEUDBF8P+iitBud0GgZs0jCLNgixmj+qcWLjrOaQMMqoLsXkPmTmA
npXgOHG6wBJKRWhwaTEOok2LIAT+A+Q7C0Yx/RTofaEwjUrpXDqHyQ1ZPU6koANZ
X+o1hJNdMECOXunirbSYTosgEH4hnGINM+ElhJs4maZbV8m1A8hVaMu0oL0L5cY/
G5xnAPg8FvpxY4bYVAp90/SeGfVCwrx+lRtzEWtcCO/eEgtBeZRsN/OVqShL0yYZ
hNMU6eFmZRnsfgER/mT4WJmSDi7FvNupR03JikrMRdNseOMZmhV9LUsBODj3YmZg
UQ5VUqgDXFlMVpks3po9U4QkcNK2q+1OZS5mhqDhRxKrsrrxJuOVYsS7zBOw1oHF
y0l2ZNQXBq2D9UVbMB2zCAQQxklacJZjXt+iTfbPYp2e0xlxLy2r1s6JsjVSPlH/
yTD+3QqLe6kjGk8KkgQieB/YPDCuIPEOQGT7JrvO+/ygwMO1sFsFogr705K8qoLf
LfPvn9PdCBagtYYNuI+7RrMi4/SDVeBH7Wxj65aYYIzOZi7n68x9rH8QjZHDY3jr
jpaUQfR3Dvnt7RHl6wlIRPU4e0rNM/y/Y5OMqlXdQRGVh7z90sHV3EB4vw53VVsO
AvM3twrppR9srCxuZce8hS4OYMIuw2YsKphzoOpLuNr6+0ddpltg0eCuPEmaeO8W
aw1f+lM+tuPL8JBCRpACR8jQRcVqulb40OukgYhDxx0CLDrUrrjraGpetCyjQm+O
t9mBxG3/PPAXbqY+GC81SlZVNgpD4TLWhZxAdgKhQ3LDjN0NEka8TNnG15E0lPp4
Zu37MHm/9/CAxyoy//OcuV/FflaqwX7AE9Slgqyv3GOGNba+lTIkTFrAUI2nkQLc
HZPInA8n+m8AilGdTxKRfUFKw4JhxRRLuXLv9wr+jRYWCqOGVP6PgfGbS7+M4w+C
O9wuXwXrpH9qREC0qFi/cuynYrKeoagsjtw/wMb4vKtgO+Ql/rAD7HMBtYDlKtoo
UgqvKif0IhnKplF2kL51aDs9OO6yGE3CdIRz6LgEy4+8voTbNntYSiz7285NYvN8
PT/sTDObb8JwZzST7gjhuTiM54iprdH0BieK+gNbDXnTuGmIZd59RshlDZaSVUVJ
S4o2+ECOh9nVyxEYuMD+Gku7FPdjKVSyIG1do+CxMSFCEoRsyzzcFLgYy8lovsS+
8cawFs0HF9XHK/1BM2HxO2VYs4oUPZI3+i9Bmdhk0d93BGOXH/yKg/eJTkK1sdF8
R2eM0mLhb5i6JlAfkFUM4OOtr3q4/bm2FJmCb1ysu8LcqZkrWqmbAwVnvAkXIbPe
QL1byEdyNPWXRi7MxKTZ+UGifdXpnwBh7vBztGVvBqb4NYKQi1NFojKhVtqQ+9P/
6yLzoDZRVila8XhfSZDbKOGkSP27Q+13jzTSK6+oqDv/ojdwJPUw0xb44V90EUwl
3taS0MvJhgZDaINd1FwPv3VQenz8/QdvZfjfqMmBdTb3Tl5/OHSipmEmMZOUj7To
DTg8jv3aXEPYdLBj2qLjUrV+68UAhk63siqap7m2KVew56wJhPGp+uxqOs2wbtXB
BPUGFN1RWsPNvuYckq8vMDPYa31BOWTRMRUpzcMR255v4766g16gvFVMCRfW+CBx
gwdI2v/gcEbWRZWYcHDkIGCEytHthYnnPLo2VbvDJYincIUEz4FCUatbSFnaJg3C
Bz/kQhNyGXDnhSA7eJiUDxlLKF0kn8MAPdWqSuzP31u5NXrVnWAZPAf7/oZkuBNY
MySm7ntavIz0r5qoVFGucc+QDZUhec5eHORm7yFAT9gVokqWjvKWYuvOC6Rb6ns3
rxvlQdRnEpptTxQ6q8JPKFN+rTz+pUc1XISpR+Uvdi4mYUAzk9gzyNMoImULb98X
EAZfOG91eFF7Mfj+YWkmr57VeSGLLc6r6i3XccuBQLk8E7K/OGdq66RcbmUV+3gc
GWXI1GmG7RciT8QgwkkUrv7jJHk+wOZJUSQZnVS78KEm/yNEqCxCPkWxZ54cIySR
OwpJA3APLZdEs3P+LBYf+mH9AJeTp1xElEsyivZw5sl58bnI9kkgFlUnh1UI5tG2
p/sAQCkCgD1bTxRZnuKEOJsVeb07LCXy2AIAH2p9i7Rhi8Ao+SAZizYWT9RWgTPM
d8SMKRJmPKftCl+w+gPS4+/GSAhApm9oA9Kzmi2f7e0H1pq9r8XegjrSP3G8BuJW
6TwVs9aiMpWlUXZ32/nT/uDKODfh7Wn0fGyERdNUlEto/dfiGeWqT4zgFlK+VvBs
m8wMkznWmLSXWdkzZHApyx2xLXzi9ntFFmMv+F6pfLzVRdLvdCtH2LF1JqtmduvE
QYNGkkCG1S8jxMKAZOGTDn8Yg7UExDtzIsFeli/KjFvbqA4UaAw5zZXUAtfsY2sp
L/y/ZzAJlVc4Iae+kZ+dFwPHwMwrBZbr0cP0EV/CpCorQsS4m7oPY43QbGszsH43
UkuFwA0aR0AbFu8Sw1TdFuiCTuRSKqy6qmmojuC/JwKQaWGKdZBGuv3Q918HLZeh
/haJcJZ7VwmYMvMz8PK/TiAjUlQ85EVU0oXUqOKtm0IPfa82N3prwMrq34EO9Oxh
JGgwr9fdo7bzStzGiSpdvFBT4sKRR1FC7BAQMFJmV15Dp/72wwXDqCDH8K7Zr3+K
9C3j0/zfYU9NVx33oyj4xK8MKAc4qtU9sIcJRbfAwhVzxkSIy9Ulc55cCEQiE7wq
tpHtOOwsSCwoXkLHkQ6xiStgSI2wwN+xXYJQ8Mde5l6tHZNpCF2unU7hVtcT1qEM
fVsFUQYcl19lQLzNUUcWcBFZmO2G0s8el06hpdMg6vqUnYEGMVdBHDToazMSiqrW
ckAoWPU7wDvrHweN0We0TTwkR+C3BOWWo9X9z27Iz1gYbal75KpQruVvUVRaFXbA
7nFMsrTRtibi3bNdNxQ6E821ANdOhsIfA9oCshZrE/Ovb75y1dxYX1JE8n1H0Lut
b/UmqB9JBq3ZUA59xfv1I+YsmFnvWst99seTtfdQGhx1qjhgOId9Xa6TIt9Gt7wl
O1DD1QyNXxaRS72WoIkqunb4UnZHCU8u3fmLuI8cxbVha1QrpHcg2pCocroMmlud
q+uHmotSGnOAjjDGwSPOvnQqVTZQVR0QtdGqLLkvIOuf9VNHHVQljxCRxlMg6AxB
IPljwOHnwv4RsYz3bXDBHIzmNkQGtnVyZ2/CQozPG++BhWxWhBTkC63HdT5wkBWJ
TqF3dWAJCzjixdShnmgr17Xk06tNv/rzJaIYa3FMXAr2iezfORHAllySYP2z+Rb8
rAXWWgQ81L0ZXTj6CDs4R24xAZfuaEnHB+pg5DG70yJrW1bULu9DiMYa8/TBcjIn
4DLC9/5k/pYvsgVYqyettBT26N35y5d9r3y4SYjTz89VdTx4rCcXXTWKsAcAopch
+G3Qkw9rupI5tl3gGvQo+vNX/QXauBV06YruvsQROgqCf+UAS8TJ8RZ+ClPE6lnk
Kqe8TlLx6nE8AhA9YO88NwUEPNRfJxPsa+QengMEMJKX9dUszFiQLOCYlmvYQ/89
h+k8oDDr1mDD2Iak2ciJQc7lbcfcgHF7F1+JPsPLRMc3CgqDNyo+upGjAzpUzlAu
UKNbDjPOh23IPRUjRtw98XWZYbOLeb7Y1JhTlQR37eeNcxeIabxQjGC3c1WE6YcF
s6OxPPIltqO64K7c9XLPZVgeWwbrTEoO9Tk3CsqZ282N1PqA4U27aDJGgVLJd74z
jjwLfbMEIlGB5qNemD+twnKqYHm5aXNMCCKFbkBp1Axn48eEg+cyj3QMeyvIQWtS
pMP6G/cctlG7uxP2AqjMMHdNzGRmy0vP3PRENCzxsnvscVukTbj9xvMTknuzYnHx
iJGaU+m88kqRSa1YYfBpToOia+woLn/m8MJz8PF/PtECO+Wg0yho1cWjjd4rsyOT
s8MFdU8kPin5M19sWS0ocMDcyS3+oTrQOc6fIS4J9mBybGHT3MlAbyoldLvpSRIu
khyXknX7QlVGSxXV7l5dbq6o4SKROC67ULcucR7kL/j2IDLmZn/zUXpcySqbnSxd
/unP0LY26iywJpPpYAPscPlxFoxO85H++DsGQmnDynORqFDKYi5OPRzjQC2Feci9
U70cub63HRCgluylJTJF9iGZy/EQ6Jvb9EhcxKj7rSs6fqv0byAIhs/4DbQcT7AE
RIIZZz0ZYjizleWiaJuVmMtXKFO+3bdfohsnHI0LM6onjMvcuZzM3ImTyJuC1yWB
u+nbayzXwryAq7Ffg7Vk0n3nAowiogb7aHmGF8JDAXneisrhlNhylY4CIpgZ0Sje
qg8WXv4jQK3cDV1yIBiP/jFEgAJ8jA9gmKtNVmN2IcfZ43EoFD/KwVnVq3T5fVGc
CsT6zyV3HgZuNlsqmnwaumGUPDnp8j+Y6wD+tadXmuDhy9wkxm2HEyp04qMlytkc
qOe8wvue3tDEoobFZcknEbDcZSmAWZAESqzjdMCmwDSCvp1YrtXP0pN0Yb0wKsbi
ND6vCn3M5mEqe7cvFuSpMFAOoLVD5+hUbijYDIQiRaNlLsOA8a68uMSvHxf+gDup
1U2g2oZGIktIUiYAeBQwOSCiM9/GZbwts9M4XF9utqZm0c/J/Fs044pan3nR/w98
7CId+6CNvMF7R4pqOv+1V7wzMzDAYObgjLrgoTUhG+vi+x2TTHJtS2X5tU88QDhm
bMqlB2bE7Wai9QUiPCWEr+K/J55LXkiFwDvimcs9RotR+Al1dU3mo2b2m4jZuh40
k06K6nAK5MUoS/YIkHr+Y/y/5PDWb04VM3dbAU1Z5k3ykwEY9tlgWxR+iDjjOG06
iq21WF6S0bmStT3OP4WFwl/MhFWyiFyiZpJBQN3qpVd2bBKGm2g551esEbhjZFCC
nD4ggcsTGmfYGMrhIpIaePZePNY9oiPf892r+DoQNASZxKa9KtjDvrT6sMGwC2pe
gS+BQLZDeZZiuopneQW9QnZhF7bzjufJQ/pt9rb9rOWOjTT1ZS/XBsZGbjddHRb3
MQJ/62Xe796/mxjKXpJ9K9CyyXlOsv9YeKIQjAD/mlv8drvu8f9opZEZ/XBdCFzB
UVhQH/Wc56uY/rES2H9SJGiCyLM7J0aUD6XOs1/BGIWG/kjvVA2k6l7G5XIL4Qnn
y1M0huMjEw2FsNHxNT3D0x/9dH/NF+COMxy1aL/tqyWceNDQINEudxpqd2/Vlo8b
I1Pduv4332gH8w4NVtIE3IreEOgByTw/5jiUFyqef0wTdrhVw9uNewlpgtqHzXAY
ShLg6LFwAavEG2IHrTme+P/ROitnzSCQYB+6kjQolSmR5pRwJ5dqCidEuew4th51
Tl2GIWDNhtWN6pFhvReF384JoOje0l6PZp9ZVjPf4edfgXfWDWOf8KlV/b1qeOBy
QuRC01sz1XadbxWaUqf65QKVYGZ9cGLgt2gYYDDfqM3BPHRT053JSOMrOqNRtDkp
xeBvfX/hcDvOa2N6+2H10X4Jcd2y8Yo7DyJP+621V7RcbAzWQuWW5MfyjrTYukkB
SkffTJ/Zux9DpYtH6JQGduLWDcMPjv4A1IsFhuaKsokUtJGYbJr5dgyZHFKLbTga
0Ulz3dhlEp1sKS1XakeNb+1WxVJguhBwgEBRJwNC/Hnxez87Bhqz/Gv7+CqD+1AG
q/q89XYw6EEqs2W+dneJqGfVb601QOfV1k5gCyNO1qYml/t0+VRyMJkL3K5rG+ac
afYCKOZPQJba1ERFGRbVEl180fFR9YG27RILn5tzPN7rvwg+SF4FYUz4lS/B17jg
4KpQGkwb7s3YF+6i483ddQOVO+goTKnnptydEAqQm/wYg0/exIwnb0zE6FeUOPsz
eBHjQrD4TV+GVG8VTOFi+ADopSWErFQdxGa8+AWcXWcnf6kOJBmD/42TEHCClcqQ
/4Lr1evqf+xycd52gJQ3GXMD4nmj9X8ZUVZqoTtbiYGa7B18gUINeB6BJOBepIdW
jRgeuut4QmTo8ByegHp0pf6UyU3QpFe/+G9pc3edmNa5X23m1/AG7uWVYPPWkfV9
7fkR/bpWdXV4MlvwmcVI442MSo0xYjm0fCvV4HjFQNBxC2qz79+RBbNm4fRuymTp
vARjhQZFSFHYubzCCkaOMxmu3r/V8s6U0pooaAiF5RigATktEYmIwwZNxMIRS9rq
zS57OI2CNplpo8ztzEyqKqhP6iHixyZ+eNTw41BuWmjcS1GX3aJFIczgGXkR7W5g
LuTruolkoOyFg5YJQ8roL0AM3CzHMFKGTgU8gdBX+eW9oCVpAxGtMexWOc4/EkHD
hDu0lGoQX3nV7kwrDThCTPa8FpKVkxrzZMvgFYSh3Ht6NzNI65lMueIeQoqZZvgb
aXZPTID1EYaSBdb6SjDwbPVG/b7lzmQUdPH6YA9gQ1chZSYiMxy9mv46M43Nk1h7
um5c80Unr1Yf39F7Ca+LND2fxqScJFkTOCUuyrGofjaMV0bkjx5k24hbliwojDk6
fP9MO1sjr0KSz8XH1PCqgHapOQO3EXkJcX7DcEb8Kc5GSc2geheQdgUG56i/WJVi
i5qkebrYFcbynBSRaHl4CgkEaSc0uU18U3VMCklC6tqKVK0tgvluG+RVFQ9XHthb
SaOAr/3hD9BNJ99egv0ri7wiGr67f/CjEMUzLeG32LkWVs7ikKjmUDyUfzt03fcF
GcFJdKln5Fk+UrEBB98MHgKDhd2wa59VrHkR4L7Nx4/YcvAXXlX7dXzPzoxvFoE1
Uw3TfdxH86Qwa4ll0fhum7i287NS421EZMD5LFOVBkTrrlCUMuuRoIS3lGpnBEnM
uFvyb04SeNFN87qp7EevBBh3nR+6I//JlUXzhUcHXwzH7MhaixYZx2+j/lLiaU8I
l2hVIHuLidFsxFp3IcA6UaueX66/t+vrp20H8SeqMQ2c/6rom5wY98zGXl8++i/e
5x5fstZImUaJzLCyk4v8ea600d/JHQOlTZbq7I2+036RjsUzccUUUGMTjpIlAUmC
dBmmqDKXawyHCXA0BvNCZMgiQn0ECFR03Skir28emqvCWL5q+TKB+N0vG11tTab7
KLgj/4tG3QGghqP1OjultJr/vT8vfHN6TJqMG3BNXcHrrsYBwoqz3ykacvcVtI6o
xwL3vVH1Gt0J30mEjWDG7HqJHOmCBGCtGjaQZlaqRp7G8LvPtwl5CuGdaoYg53/C
gmpnDq5UARLlS0d6a4eeu65td9KmKtJoJQHRzfROeeIHQAzQEILkWly/JASWxO4+
3SXiMBgxA88BKMxMS/XVFxw/1/oVbGro3gSgK2md3Kn6p5agrn0o70KpJNhBRR3p
vzEClK6ess4upyVMJtRRtZoCBugejNY2/JP07ALK0MLbl8fIRmI/AL/AQnUHxd10
y6XOu8IgJaC5lehEiQiXGmpoYio6SMMGj1Gs0vG2HJvLLdhkjXq2DGGJZhnpO9Km
Pd2jNy+/6PGhCtSq6FvmSnwsrv2smOpOmSig1coMFS6ychnqgX++ARv3EuZrsbIh
83R7RbUxWJ100sbAlAhYTKdStQQrPfD8hNQiQKhycbWlTObCgYOfGWFDUMNnHn+f
0elqmvuzJDZ1idOoA8mGHBRCHLs3Xft8442d9zOXJig0NbbF0fEw85ypF86XD6SW
mYJmUmEQcrP/nPG22Ze+AptQ9dYK+hVueZqaU2Kk/0s/xVbcnnZ3BesmahL+38aK
w9/Qhppn7tdqcdZLROocTKkwyYjqJnJK+N9K7RRxS35bq4Y79oIbxJhmZdHT7uyI
cS3NPilDGZueUsO3H7r2HuVsEMr9I5YhwnyraWKMfYhdy3I7MwfAPBU57hpqakhf
KEGXg4MA3Hd53iC8tOJgY0oM8/HZDrrbsnYfPC4z7Y43fI48RfLfJNOV6WUvEEVK
di7Up08VovS2j0izadZeVy3/C+9KYbt/qUaabNohZCSmASgYzQVLDK+wHb38zC7K
/PaR5JR4IeaX5BSFU+QETGT17g8teb144yAdxMGtltCmeL5OLZwz0V0+ONTE5hPK
4kdG/N4QIUVNXL179SGZkTqOXcEXgNCKkNXTxXHi2OdmptfW8KcJ0deXPKd3LVVn
a3d7bh7WzpVcoSOCTdI2FD8aThVqXxgDeqTBOOgbwzwwoUV5IMK8U8MRfQb1GAK0
IriECt9Mij0fQfXhm3tmRgjdPZKsJIMAQb9+2YYh56dMOVYm+LYSJueRBsZ+g2QS
CMm8ilP5koHxADmMNh8Xjkbb2ZKZ0r13vNFeS3N9TKwW5Tyqz7b0ihVZkHKUIQS3
6jf3ESrOWukqJvvUbfFWZmaBlPv/t8BxbI8hjq0X9gCc007CEtPb7JWJfjqCXCYm
of39rTSslvwMg8FIrEAnF01/ZQOkJupTkrEsMJuuz8jKdUf8yP+E+le5D2Pflipy
UW3QYUDYzbWQiLuzJ0AfdxD6tBXIMZPrdUFciFOo5++uoOvXfimMwvIo1f1MTyj6
dK6nGu8xcuSsqS6aJDNhzGflOKPa9ieiKId/cKDJPmahNLp1uCoN1j4JqCTyqxmo
o7ep2tHEO2pZRYFLgEmt4jl84vi6VcvYP1X/WLRTojHZmxAHdx43qKvdCge/TBuU
2wbIwldNJok3rFVaq6AiO1NAKZU0Y/TUfRM7Do0cAjO/CnfgyKLyGoxAnc6Lo11r
EuA4ZdM5NmC7cLxV2fbZwVkFEiX6OWD1EGH4PLEWQe15SkPDiAf9+PIR82VaGheb
/1OwnYnpf6MdhDsfDVW42Pe4iPIsFFc0O0KVxPhHSBW5Ts9Sv3dQMTKF+nV4PMPO
yw3ImFtoaf5s6FOC9c8n/G52grjQmMGNFNyufEm/XarVMSfzQ070r1WHfk6detZs
jCSRR/+6f9V9EkKuHHrxYc7CkbOO/2mTO1GETTj5K8ezRlwcBQwUdE9OY4YAV7xc
16PbMlxKnR0p2wR0yzUdhaN8rJpK4LeaVIihsccaM9JEE6b5XsPbdjYYyJFHL0ZB
Dyw9eEMTvO7ifVsfbz3zRGaoi9JtNc+vaHTYK8DZeQvLH6Op9TL/1ZG4eBA6AV1B
zxb76Pjj6nx4wtgO6H6q6QJaxng3MC5OhxVf8wOkYkn94OdrPsTT9DY33Gd4Fglj
mLvKIpTG9/MOYVrdeO+Ls/LtbwHftIauSK86X+a/j/cTNqNc/E7eunXw4l/5yHUY
yjX40Ch5O7YSIJIshi9DpW6csYF8ONDX/V2pj4htQ/v8XfmgvOWraIHdMC23Y4Y0
vslXbfqa3ue6ciu1mRLP9XlI7ByNg3vL9xT0ClyKwbfhtDWQb0NBKcAWo8vPUtS/
69pWuMS2ggto6Y1Jgqfd+mllqiT5ufvzLX3hjTSCppxm9HqImr5WlHR57nS1aCOV
O9M8dk0OzaX7dlo34KCWnjr/Ni39dodTafgGlC0hKR+oW/aK2Qhje0hHT/l8Ayhc
+ic9aDZeouQQRePTs9vZ5adItQMBGtrnxt/6SiXU43iQSsskeg0Zx0OwpMM+eHJJ
lLBdiAZSW99gvb46yRNGFL+1WT3YcrMzPqrewI/Ndssn5jQPhjy89sa9ztyMfn5Q
QKrBOhpkQMdWRZNhQ1/xrDgnMu1bcOqRbTsbAYDRDcxarl99iqK+kDUQqD+dur2Z
UCOjb5wNHRhby304BoIgrwlaQUWf3ddbnWwEuHMhfgL2uLNUIsgfOY1aJHwr0yMp
M67vr6G75ludJ0ipr2Y+8YEkugva2D/udRMwdWEy7vGQPqEf0uVJLtEZNnxBlQDU
/Ot9pZMhiB9U3n15NoyibcpHeSWUnU/hEZtCIlGwVO2A5mHO0/qJSqZOQ9Md6/bp
9RgDvDj9eSpWOhk6sjjkMEOAypYJeghh+83eXjDT+AtrRik1hD+fA3iMovIpQvTg
MDdB6nkMot1icS9Yd9Z31ZdWcT0s6OnToYOaxCvljoKBZc7iXq6R8XfQn0T+okGc
ytCLzbbyY9EVKVdxAY42ZtFhlsaU691RrHAeiAySFSUbukQZTWWL4CPIT1SZonNF
eKie8sGm3XtkFDFPAp3Uq/jgSAQvnQ0hMHipv5WrBRXHCJFNdbCmMxJL9CkQgR2c
XtRZ4jY0Jdd3+sXgaxbbxtT5sW7Mmn2BXc4Pyma6Ebg9YonyUrAfkkM9ol5+YjWp
s+4RrIBCUeIB1dnSCliLUsRXb1A0uAj62sMh4tJejrqoB3JRdfW+lcaC58Wdyj3/
y4ocS1IWTV9/aQGzU5anMHxqQXaR6K3Td+80rMoMztmzmyFNKl8MsqoBtigkCe1E
oVR0SEeyJ3Bg532KqTwp+SobKbkno1NwT8nttiMngBfP4aC+hhR4tiF5QR09rU0/
AktM5+E9k2guRfTyyGCnetkflnttMJUHexMbHjS4nKm4er5em4vkBlI+mPuLHcfA
+sNqF7WkFWZPyIltkDhqa7o6gfYuVZxIzEM32PyJJvVdtm+sdv9ARSvNTQ9mnU7B
6dK0bR5qxyc3gp1SL4CrmCrUTshB8MK1RsEmUaf5ftE+0eZLf+2Q28xFSB7RYmVz
UhRnjXUhGmF53wgeCwgGG+2gt8TukIroPQhBEv/61ZvkAcS7mtH7r6XejGX+aV1v
7WKkYwoV67giCbyJJaNbareOHu0hYcMC5M1kec34UaHPLqu02IMLHRU48clKepjy
auyzHeZzaZuD5FZUuW56/Ct1gSiZTj4sACuLEQ7jKnFubALstvKWb7g+I9V0ly/I
/pySKwLl+9xRHIHe25IIyKSu3QzadGtEIt/c3aedc8OFevg+KiS3S4vs9I6M55OX
kTbvGVN375YY3TXD3Q4k1HSJowFXRuG5nMF9xTF/C3clkQ/iPMIDyfmE/6nZ7k6Y
8/MF6DI2qA7gQWk9vNDxsdCfxPOfNvq1Zp3TQmfDLaQ8nXWEHeZI4GwmT0o1uler
+lro1Dj6Tf/UWhCPxXi0kVIGQ98dUOlwV46VQu4ZZxpBa2gEN1cXBJ2lj7yHVOrT
RKVLT8WZLx3jPd2i49rRlxvyg80KxbJhKuhzMRF/vXsBywLAcioNXBdyEOI6WYaM
4a1bfsAed0/BA54bj1wAeLeISsqyTXpmPvzwA/AMWcG0Yy91R9xuTEmzDwU1eDbg
nOpdQpRrxyqjZVkg9a6Qas6Vf1HSw79M6NlJ+Q9drpqkFAEz6uYWUPMoEy9crVYN
V+xFheuOIH3XfP2VLrqNzKew5a0o1XfOHuTOinWGxsHvUwWK7/pWW9cIdo8cu2z2
LL9LIGHauWbPzzJqJTZbCwvK3cn0PyG1Tq4s36WCByK9WP8MfGkdSD5THBJG89sR
R1/OR9mqbQjxpLNiZwjfwwVxCbPbJszv7ok3mFUtXwmuibk9P4J4GmyPq6Nso7wL
z8eHzL+ts9KGXgowHOI6F2zO5g64nCwoanHZGPueoz+7/Aa+OkM9dyzk4G9MPejQ
ZNmXL2ei0lIQr7y9Vkj6m1udzJEWeXD/F41bpDq+JX9vEu7lSLYCQIQo6iYyvoox
pOIBheXklsWyOuit8LToVHm7glUb4/wXtpDF5LwwMO7AjyVaT+G72y6Zxe9NuCoH
QOglOu7n658WUHjuST7ygo9XDS3XTPRlh39EV/ipueNyyZqowCPzfWeeb+VkNSj2
XnVPDw6t3msUVLCyMN7c2uaFyF8UBb+VMlKlAEKvfDd0pvJKHDWnbhV8jFPPDUH3
wjnlHZHGVk5UDs3/ml7D/XZgynq5aGd9EQJzEWE65CB1DfsfvpXTw4FLJlC36pRu
LLIv+4GEkWku2RS1TY6j6yVkLJWi1KS0Akhyb1XzANqCoaV1FLBNuVXuXJTr70TU
mMJ86eO0Pshfuz1oi3Gdqp3y4O5XEWKcaB65U1oVkXFfFmejifJpQU5f/Ek9Sf2U
q/T1UHBei6aeauBE8j+hnM62vFMOtWDWSZ2eTnN3hzQVp5QWOFmEkzs0zMgSKrIu
JSx2wRXuZpk8cEhQ+TIAGje0cLGLCWPiIBkUMfNX6DfXj3CJwaPBq5Uy/WtV02TT
HDy4GMFyLXAJcuVnRe6yYKp2qWNWCsOY1IuyKRXdctk8zkIeVv/dV4KZLkEMs8kV
PP27mZgtAIZrvAwvRiFm2e5PwjOq48NAs94numpLsvqbCfOtEU0Z/T+G8I1FwNiS
plzEW1608u8/OkCrFCYZIakurEymnlGhY+job/mxeksQMRM5nZDZZBblBU63rLZv
TNr4lVU6lY+5mBir22QTal5coLi5HI8pCSHezclCx6FCbiC8/3l4yeMxODq9584u
uBpzvz7xeMdIWIsPrABHGX7akn185XQm7DxArGpI6olBV337BAxypvgUIeJSFMqH
KBsdPtxUIFfC7KmyEDA8R95a7E5zSHmsWsicDvhPf+kA0SVICcD5LRt8NGnYzfAX
GKEsPZUyoROLVgMLII7ZH41Kdh60oCTdzJcvER2lcOk3ZOx1QLbEklklVgsxLqLM
cqk+JcPTGGvUDc6om4Ul0LGJT47ouGz+tquqtZIql0V7l+b5A8DWV/icsONXoAFD
XEfnz0m1hdH4iRzbQSdhGNYz3LJounIkwzhcmnmnTB1P6bS6R9xEUxv4rGcBlce1
D5EUVZIC38+UxJzVAsBp/SFZKMUuHmxyBe/v/hH8WezZ2jTK9DgtL9UI1dy/4TMK
DC2Vcx3xFr6UaPsCbWzh1Oi4euIahJ3cYuxnzb4AM/hZahCsEPm8xcVYnIZN+y3W
BYj2PpUAMN8JHn4yaIWOlQ7BISnGtEqU2qF5293o0W96VpdmgWk18/Kjq4C89iLS
JHZkn3m2xEWO/HAkzi3nUa7hrX3U/yVpJfFMcwjxOrNocFr1j1xoQwl/viLv+jIu
797fH5nyMnbe4UYZkgKaDbcljmEjGda54vQeJUia4PrGOuwhOk0Kl+aJlIwl0oKw
PyzAa8ZHfL8GcPbpQMPl7ttTNdnI17PC24FJK4XE4wjzTz4cDV1AqcroGX6dnwUQ
xWpIod6v4Qy3SKD1Xc/9CLKltUYlmf70qWSb0NRGmvt+7mqpmLcjs4jfmWPon7n/
r+OarPeZgJTG0GMSn6UwR23FVSwAZtEqNWTEplma0tF5lwR8euBZdj32wlr0Gd3F
YgtA8z7V12OVeGIpCiyWb4dltJzJnJEFZxFWIpJYgb7VycDWTh+qo//KW+acxwx9
9xz8mTRHq+HLyQ/Ym1hPwSlBd08Z+YZxVawPu3pvUtp4PhK6oEi424pKhzJVsdMe
a8aL6veiXwmOY9oS51+qQslDSyerWNltV6K9iDq8CKlq3iDgSguJszbPzRueJY77
Kubqvi8z4ZRm7iqjOuF2PM/yp0N1JW0qLixHxIUQ6ncd9PjPTRpkTWwWALal8LBj
DTEoU44JDpfdpxVdNfQE5BGjy8GyB0OpjnOr972FThyt1trZNYDIZNDAZ9+62+j4
b+Pu5WpWKHPLQuczutdTGSHR9duP5RDVt7JTEtiL14C/9v3vaaQ+FGueIsVJiRcM
wIY+fcZfsGy1U/SOfA81KMXcOEmZuW3Yho1Io9MobhROHskxNXJhcGdE0Vif5Miz
62mEpHPEfu3yLQh/V3sihSUKcwilzN5j67IT+Q14msr7KMYKXVbOGTbiovRkb6Hd
p29jJPtS4m+f+Na0PCqNywxDDXDL9osBDTY+JTzGe5mODYZ5mSNV17MWO2r+v4PM
TP+VqSrlAcSt/+6CTS8zBRAAggjtuKt744AO/MiP1suREFDSHcWIl+MVjk7V26Qp
SJf4fRCBiuYHHymSsqScEMXH7iVQE65T9R4i8AY+N92JXJ5jf4uHmEUBmlRU3/xn
fwkkCsFRFgG5K8OdlX4i+BDnxkSNY3bnJq0kuoySKHCATOVE6W2zbQbrwX0JYF58
HJlO6+donCFRUV5RAyoSZ+bkBDcmtmbHRj1Yy1rbkqLOa6IuUxB4WHnaRiOdZtJE
cJZ+femJaJagudfS+v8UqQWZuc8fTIDyVHs/pPLSoE59mCxSIaL5KGGDwrm4MuxK
WdFKmWKEOKCg7lsOgvq3WY+9UQaivyVp40095Kf4unjyP73Ax2U/fSZYD6jHNeil
Pa/0l4bKPyoUkrK9Nd7XKTVoPH1PAPnwY8Iy9zmQSmbeTTvU8WOZMRlAfebZt8TI
0TuKGBLhUfMyiRiHsMRxDqcO85pYKocozmKSLecr5hir9OcEA3+icigyS2HJjf4B
YF33AoY0RinzvCiGYRhd3z88qXn2zNC384CftW9ZyFiMwjmf5l+xA9ofRQ2iIc8d
bTica+/O1/xFGYMzfjFWEVbOWFNxzwxsgRra1K0gzgKalEyb1p5wPYgzX+9qz46y
xxUzjDJm8RshFZixhK1mtEEXIQaBi38V22smcd3kQU6tyXIYPjXx48dqb5SgYFsw
Rku+n7Ow1nIAb0FmbDk4uNFUhvAmj0qdxTfnBcZHwXhwaxOq6PDe7JQMKXHNz3xQ
PyqIl2K6jQJwyBA2d0jDEqK8H2ZiyLure8fS69eD0fTXriNp2c9drEOxh08YRDdu
/AOF4xWQ12R7G9LBZg4VAbU88WP1PD181d4reyKRhPSMUZJbrRFHID6TyHJYdW4h
tXqXrqPAOfuuBBJmP5fL3Qmt2/0wrG+Shoi5DEcPMMr4lPzwzP02rX3tUFS32VfV
tFe3IrXuEbatHT5590n+1b0JJuDemJQcZTicCDhMBqsdZEVMxngkBjGKH5rwDH1Q
mVdUvj9og6QQXZOCUmPWnCm9f5McOAxNRahBFrqxl+zMdQsv6QOmb9lsrJGCnGp/
FOZm49wwVuyG0Ep4/yfxgFNl+WrpuZ4xs3vPmwV/zIzTwvZY7ogsi3nIdHiTPVoh
ZCl8QT+bikoMof9OjM8NWqk8WVbRBSgGLO3Ince7ZcEva3liaH9zyYUNIz5sDLrR
Fj3bNiJK5gbkBDNw56IJTMV6PLM3KLGq27NIyRqlhU+BRAdvecToy9KkPt7Hz5E2
3bYox/tj7wyEpWymkCatWt3RZHQL5ee8/mB+2Nu14CTesV6zXT6+az7GzLSr6CJG
Y11e7AyYw0MPfvv2qT1WypZ31C4OrBf8fAx8ndxQNuOqcnGPbWZsRMe4uG8hcGZy
A7804nEpVWOQpTEIIyvYp1DDBcI2+jB3SI5VnlT4ZBcvUUHhDiCf0ebBbQuX0+t0
w5kLE5z07SlldISGPHhMMj441aFTzRRRBFZ8lq2laMaMgwfGEuYqdef/RUeBBve2
K2FyUzDFHj6qhMzi9XmRMgC0heR9mzpN7Mappd7X/4jc0vdr3I1GkeVD4Koi6PFs
gTRiYE/jdkTKslthjIKq6qJRD7kDpoMQEnY2BhNlXm7EbNItqTQ6nz7rfIDh/ckE
DtqN0GfFVzUYSzklnHLQnIdc+FOZNVhBr9MQLvtZKHIoNjcDXFm/F5pzRDLohKBf
HPz/YuCklLoE9MdC/C8Tmw9Kv71Sz5Lg8mXuOZQw3gvlZzxvJOvXxkfoi7ZO6BYa
QZvo/dVXRhO/rKdrQjqimZxXxsDKb0hhtzcbK+UIo/3EY48/UAYQ2IHARXW7dRm9
qroXus95EsPHvBF4JjZaKC6Xlq8pC2yTEvZzyU+nYbxPaGNZO59E2arAM2mJ4ENU
u5dAuxwHm39GE4At5H9Pn+WnR77DIARiujLmD59L4W1HWdeVGeFmlPlqGrVCup04
XLRoNT2lLePKBKFPRVpWli6+ac7Vx8BjqRdxgYIFLW5JNHhzaW2jE5WovLwN3v7u
ygu72iM0ldpLTR2/5w/frmigsk4PJQo3gaKQoFGwVHGSoLf9fga86PKqdGwJyfEp
AiOs8rRMIWGY9zkQFdMlq9QFHvFtRNwJWF5+bAKiKoDYolciiwa778MMe+p4A1PV
IWwwNE1EidJs+IlHcoRs8xIz8F6/tIj782+5OWPIMbTWybs6/ZhXRnAjkh+BJLql
0deehJh8kXs+gMK25wP0KaVxBhcWR9fYUDTEPWwg2nyeLa+XyP5sfoaK3XMlpgqW
gZDWT7PBc93kNV2bpLVfIl2M3JpC87sX2e6jpd7SOtGayB0u7Ehh4FKO40JO56+w
hF423J+2i6FaCCOZ9c4Si5tTe7hW5wTaPAaFEYkSqihRh6nxbKbud2hwKG8HMj2W
0SkYIYoP2HzVkVErxqxqrpprnhUxA04Ul24kq8EZ2di5JDbPPnC/EFj0ORUzO/k6
ObVO19Z3NiYT3owLhDoZFBmlVb780yvHAFxay7zyGJnrmMjFe35PrarneLBQ3jBz
ZGDsOiKmUfRTXZbcFOZzcfrZs6WzuU2SA0ksqYr+/Oyc5ry7va6+iLTKM8RoJBRi
zAbWFp1g0KAUFnT1ffuvT8C8FQIGGgvXWSBsWtALpb9OeWHCp/i7m2LUlubrIcQK
ag902qXB2t21YhGrIjQ69RWErvUnOIlauBoAc3zoThhSUrbJD61V3YNchil6S6XC
G7MozhShsLEV/lGlVtCw4nX1aeHdKjIuXn3Kvn/y0IdFxu85z/wSM0URvRtPDg4c
3NHWgsX4r7Lr51owTqro/YkFQ5Wxv9ua/t354zJfkREpl8Jxf/3trKg4Nz6mq78z
Lz6+JTkca2mnp1rt0zxaR1JcR2eeWTFykOGpuiKR+E104ZgAAh3XMGnZ0QNrw6ol
imZJsgNqALSy+tBleU5BTEzTWOCXQziLb0DIkytHFdfwaR1Ovv5dKQxlOWMG/pJF
KZN4qR9gEAA45o+qDpxRjhbuMsFIw6yACIzlDUPS9XvM0mmdXzTXhYHRznz4jWxD
bQDdaL1j2E7EXG6DROZFYkO3S2P66S657V0IDVYj6a7GqsuSfHOsCDIWLPyldNBQ
nbwS/ZLTr2Vmj4DXWHQBxkGBjbUSV+vGbkzEhMSfDsMEDq7IP+pmZ4N1+JlKevf2
H9cG9DJxZUztaRP3Lxt7ROn+2QZWc9LtiOcrEAxtZXdYfuDHUPWmW9jbJY3CQb+s
2akVJ2z2XFsV3eC8j36+4UBrUV+k5iyj3R3g9wTND/2BIRLMYiQQ0YEFMbKc6bVQ
fCw+KW5lfH+SeB9WW3E3wZPqN8oPTa+UmkO7FXwd9kB3epRwdNlJaChZJA3u5wxR
MvXn0VUAbEp0O6uCEXl1ti51funt1NQTXCmLVyRMtO0GsqElFiNah+tCtsJDRbOv
xoXDp44NIquyAIe96BOBpgpuOLiHkf54vZMRpveP7tODlLQfswV9QVBE+u+C6wge
Bu3wzQRsY1AFsTHfh2IpS7HY6vAdvL+lhgzDo5NNe9Z5UU5/DT0CbTEmDmsXVhmY
JvUhMT45OtRm2AMS1THPseXLlxGt2jSrNg+q440nUeUiO6XetzqVqH7WHndw80n8
iUOB5aJVC2XYybLWkW05jfrTwcPkGbmGFeNpoT/VDuZ3hOVN2yl0g8f9YSohPDhI
nVO8uEVOb/4HiSmL80NEnFfcenY9CIcN95pQqCdzhYPVV+SKRFuH+HP8UMGthd7h
twMFaTMDR6Rjs/DzskCW+LiVBKrLcM+WO9xOGujfORLrtzzJ34CUewWuvZmmdHRv
tLri4qsAxMiQi1+zWxW63/RfWpnyUTdTvLWPPbj8QLyf39AhDh0gSic5HgFXfSOy
c3jSeoYmHMjksfThFUg9sJHVB/rocOytjHWu0Jm4mS48LiGVpN6c2q16jLtYMRmZ
ENVa48KDinzlWPeC888i7ZYv+unCr9wyC8KBxIvBi++up5JD1Ag4iPMKnwKYWQgF
HDV2TEdpJj7t68C2tDWO3DABcAkrCeO3SGMHgKD7TAi5H/m0EKWWwOUC/C1Hngog
xj5oBDz7RkaAwdbrsIWiCbesfwaq8PMu03KG02TB85eMnf1i+SAwJJcLytubh5mt
BJKkTUXcg+R4UkYMbk+djJpTtT2XCAbM5tSYfllVncw0Rcfjr36GitiZBouo5pUn
YVkocOOe8y20EPKOVwGSNaHAKHqh+lDSCRNPyvb0IlVqiJjvFyF3EychMzsXE/2B
K1Ow9C5yZ8o3W8ZF1wZVULkNDqmJQ4Xsz4G/ic7FOsU5R/qX8XJoXy9Ucyyu4XWR
FaJHfIR98HCh0eYcKDezHCZuKlBIeJNjL7opT2s9ygVS6cdeIas4WGyZOW6eEN/X
3W8XYEDbzzY1STrSjID3Sxi4/q3FMBSLTW2t0nUDm63ZoYgNbG7v2U4jepgo5SVw
4BIu7nnwC+rUsG1FtGDcbL4U4xGjpBJmyFGZ3Vwkaeo/oKYgM1syQwrBPc/o5OXy
jsyL+BEdNz847c/J4f6Zrz14fPyZzs4VQrCUsPk1FBP23WLzvvH8eEjDIwH1rRqk
9OKH8sfDEkar8o5Bw6F3zhydQSKItjOXf3iFt24Vx5PFVx1WIjvvLYlr+UoEfPZA
nw+g/Pv4sd0QgBAJwKVW14JFh+iXG8wLzYzzWPVRd/ve2A5qL+JE6D9boY2a3rxM
5EEtjxMz+etmnV1iHYTnPsfQx4uRTjJTkBzBVe0Hps+z8cdf/BXyLrjccM6kOwW6
du39tfSXXnMBec7VdSEHUgsuCCyf6BnQtVUc2q6zz0c25Go1zV19HZmpxj0rsu7Y
0Z4cB8c4EVOIJU4MN9AFPtrvnmC2bUb99a8Fm7kGeOhWOaJOkohSn+Tqx/qWH71V
7g75ox4fKTaijaupEISOg1OhqJSvnOC1TB9+q1zMlcooyuaH4nOz9zKvV5y4rjrB
eRI7ir4KUP2WRH0BRVn+LYXc+t5QTMZOTyWO5wmVt1Lw+vEPT9RF5pwo1VubbxNf
GwASGYQfk71FQBIddg4JPgX6SZYSqHqVtRddeChFh3WPUNhVxpUfNZ5bunNd4gAQ
rSwADmXLpR6Nkz+gh7Y3hxgQ9XGosUcRl2w2P4iLYIYM9oJl9pXkc0cXgf6DVonI
t600pO1sX9WhlsuizollzJ/Yt5/Vr0FBuEnrehWgJUN9L/FIn+TW7EMRR9kkfgnI
Ap+TrpfIskS+lGYC8vlT/AfPvqwWlgU3b+BpsZI5J33GZd3G6YMsaYy+GZjpg/HI
EO4JwRbi4LERxdmS5tNPYkjYEq1BLoVsc5jVSkUsWVUzJdMYaAkbN3QHIX/Kzk5Y
IPRsQoh8eTKpV4VkE7nxrrZAduLDG5fPWhLDdtn3WTXUjii5U8ZthQyLmz3PRRL0
Yp4q8Q43tiWQUyqQGzvGZkIRog5NFd8Ay3ZEPPT2HnS9qv8LZWWGgUrL1P42lk0k
smc0V1r78sVFF49TqunxKH/3e5Fek1jwiSpDMt+ftxXztJTyBEbh6Zev+XkwSjDP
K0dgVEOPDc+tD6IIUgkh4scKzVG2RdPaH87vUDkWcs4m+UhjoDr0K4asTS6KYgSk
Eh1ydcbNc+OB4jNDWUhRBU8OPPPdc40uccCc7gGANZqkxD+lbCzhHWZ5gDvyezXt
s6+tCLc4EYkPQriCyEwAwunJ+RGnQerl1rukF/v6xB1tarPwc4hdd/frZScXdPxw
fWsRXVWS9L8Y0arp8JT+HC4FP5F5U0VJxKQ+6O02tEa4lf1Fl2yu2ewy7jl9h99d
vp2PJJweDTOwxGY5hyiJPG3pg82wybFQzqym+qFis/PLOzwo3xn8TQo745yZFHsf
OWD7iXfxq2/rOotQCcOT9/pZ3HH31bmsoWoJQJnwEryAiPkbthY6/TcHZbj2tbBB
OT+cB/aSf2QXeJT6cMbhzKeEE0lEQHqdCKzG+7KRidE8HnjSq5HPMlI5uaDRRRpB
Vh7+IIAMj49nQYSMIt5fyNW530b1LmdOmuw8Z4b9fj2wEMe/qN4+83XUP6F8XH0p
QVznNAkck95raTfCaL2iCI5lwk01r5W8bMf3y8t/3fgJtnpm/slCxZkhI54wcRwo
d+eEcfdpXlV/iD4WrYDd/HBWZ0vlsEq1ydXli5D92au61wsgVHMe3ccKkK9piuL1
QmlnAqWkLaHPXxJd3QZNR2KiRszwDxND6wiAFZumtHVFePBY6qfmeJQtPKEnNLIL
HtrNTjsBYr1fR9owlxzAKsN7V2O7jEAOTXQEMKv9MkWUsiCBQqmlTmKMbJd4eYWD
k0wzfHUPo3jhkR4JiNgc0P9zUEQ8XCwzQP8DkyV7f4WCFvJm9Xi27ANxuBRjgtY8
JzNJsP9zqcnbAINlWEbgkxWXQsSVHIC7u0qL4R7E9GtcZNglvGggnpLs8S4xM25G
xKffJw1NTq5fcZgVCc6RddfaFk9IXLRVtPxTAIyOOhn3gsH0dSsOitptxIKQUMT0
NtMuR8eYz00eDGK5VZgoFgnagv//stlYTi1vuvYPcbF68LY1EA+nNRrKKw13Q3yl
pZfuvVMQ+D4bZ4n4aRnvOusSMxhWM6nQXsDLg756fTMrGPuzGautuc7lqPMxC+dJ
Cxqemes8qMbm733kSvWJMel97FvXdeDguxOuWua5mdq6vy488VmGFrDhHmKGWkpT
dgUxxiwBQ/ltvR7jnxr6L8tHAxsJA66F1NuV7hiNJJdy04DKmpzle6jRVu7a4SR4
7buiMw9brGVNBfZw9ZoUcVNFHKL0qeN0/FIaCmAEITgg0Tpf8BOxxzWhMChgeo6t
YDjV/ag1aRXpsWR+GXgRg9Zqijd2G8x/QSb/Ed8hVn1ytFnM6OH4yE4Y20mUcL5n
RyzbU0CrkKjxjClNhttmZHPNFCaHembj+OLeCmO1VBQ=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
CN5IwqG4Xoi1Rbixf4LDrf06F30Vl9rX/iZ91PzvEYYEyYcr6PcGJ85CJ/erwQgD
hVlWXfMSGTeEBAZXDUfrw5h+go7DKgww3NxXe0Ch+nSPXhv0vQHh2Npxl9n37v56
pR6lYmvAIchnZN7+xDkQm68d2UMnW9jPRsCFm4XiDTyq9bM9/+bYOfie5Ug7oCyB
+gp56o9mPe1mIHsCEUvdYGEg4t2G/9gQ3nNmH694mH/AQH+NW+hfOnSqK3JGoZsY
ysKjNDhWqB1tJpPftfl3bbO37GKhUL0mHaGJgMyZp+WaZ9v5fDMRpgj3oV/OYQI6
6jDmVnEKrU2mEuBys2iSKA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1200 )
`pragma protect data_block
4dvFzG3Vh+D5UhCyboJMjOrs4H5KSSYcFXrfnLt4wirTcThjwdgkET9YL/YXiCzZ
Nok/RuAvugmHaOC/7dPKUWwkMjU7oMt7e1+BUb5/vvwvXol1rtc70J3PAs23Iy4u
Mkh1LZA0SEQTsh6Hx8ecHf3t1YfjSbmHSxugfMB2aZz7782QmdCzl/AnNLRvxXK/
QrfzWkeepneocRpGMkrDqbQTxX06FxTEIOhQblY+xZHOOkJEdwXaz3+sZROq5cnG
8NG7qREY817bCtlBpJHhR8kedpBVDcGq5+HhI/wcF47gmRwO1xSNKwF1w4AzCO/r
uGeY9dvE/1SGWI7MuJzoPYtI6oEfUDA7+Tn7yqiJ0O6Tv7t6AA/PZsEGWChEOm1W
PVfR/2pXgDT+Jqiq51d9eiOynCLhhqGAh8yVG9zC500DDgqWuB23zU2INHacdzTE
msUprY4l0V1MGGYUrM83JN5MM8IPVt3J7wp/KiroT+JSR22b0fLRXfr7uJ96znaN
4YpyQA5JhfmwL3JUlQMmYgjhOaBHN0Oh+9YBZwIdehmSXFZDOqOlNMHE+5xK1QXF
bQnT+1WHPTjMctkeqPa1u7YzPPdAua7ia1LVrzdXr7mXrMBKtZGLI1YfXIpVQFXo
9VDGdgcuieJhFdyYRwTPXEkoBf+Y9AvGVN6R1w+XUNUshmzN/geQw3Q+hiVf1hMP
Uh+bMJxctUiNhzj/7O/H/jZZuIxLjwWPEY+K8Pt+UMMpEWNv0JEs9wG3enIpn+Tt
LpaKoDY/sj/yvZ87VkkLYTJPuf879xfBU4i8TkXGSdabsSNB8esvbQe1Rb2pJ3NY
/4h0P57ojBbXYpReCOjFnqzRl+KVgAo/l3rSSW6dH9jncVWPv3ng6kyLvkkmxjRA
u+PtQh+gM7mO0VrSvzQdKXJ3CSBkBWt2sCiS6ZmKJNmLDbzuWi/jHbD0LmjTnW6e
O2q3CbfWv96kzqq6GeRicwGCSKvY3FXv45fwdNf//OlnlbtSmt4CbjucCg2vanEW
MD0mWK3eKS5prYQ/YmRsseWgKeiA7y0VnbuShcoVV6pxc2Xl3z6/DeZmvb+1aEaT
vkI2teIh/CQKDS3SVn5j6kHIB4Sw8DVJEpCjMBnMi9EoY9GLfg3jWu2uEU7qMujk
GTtsajMwNVO02hefuYJXuvN7709S2GdBwKTf4NKCF4Y8Xv3WnHV4xg/whx7MT2fR
S3LGmG2zDNhoQ1CXyj4KE0oo9PD58LPs9Xsau53D4WQmy36K/rzTTd6JmGNqvG0n
ehnvK/biZjHTUfwexMc6EvRYglvyH1ZBgql6RHuW9NZ+HhVt1kBQbU5zBERY3xAs
1T7BZUhx6uiIDMRyPB4XXr/zcrr3gbEhSIeEhLKnE6K0TFc5OxsBRLCaFlWUYurx
BZAB8tKPj3bGN82IDvOwjWhNsv2nbFp+QLpeuDwPtncEOX3IgLruGhG0l8CaXb0l
d0oNR4G/49nrn64EayK1MfY8Dijwy2cj5yqLKRzdaa20LlU62S5hicOSAMY+AGCH
gpZbNzc/fEGEyC5lw643C/LyeBgtwEEwZfuQEwxams2XccU8VZo3NsqMg/79fxSz
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Q40ZzNqA/ExjBeCV0BJd+PKEJ+nsE1YvZzq+TxYRaLsSaWwEc1OVs3y3BOf7EQ7p
vKmptuQuXsEvO3X2HmzY3bSi637tUe+C+RPDIeIkStlIfMhbrmRTe2DECBd2e1w7
xB20AnvDMeU2n5RHmcAzm9P+HuuwVukTLOcGBTgwNOb+NDIiKhZgvZsIEdF509o9
jGGyPpIxhMfdtm2q+s67e4sZgMwHqgaYpX1pWp70L9KXwzgCw2U0e4dLyR1peH5M
wUQpOs13tUwbiQ0eVwx0MZ4w8KnHkVt8u2BLW+ofz5iuQwAuWlu4HZ5o+Z5Tn+eo
01BSsMaz/IayU761PK7B3w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4672 )
`pragma protect data_block
20R1q7ToBiVHQTlMi8JMcB4EYY2kpaCAVRVyd+NYsC0Rq/Ms0qvEwnY6IKatexr/
5q21OpBtPmHZPo3dGEbs8LoYjf1/7OTlDWd9pFyWwhkT1uydM0ZuUT/m+DOSRR+B
wmXz6phMyEAWoaT6MbuwxC+rYAyqHCDcCUl02POpywLl7vCl3ZsKSlahpy8tePvs
Ld97RN+uRIxHjJwjGWyRE4BFNNwM6XxC3aNN7XqmRVv0rtuB7gJPNDiJfePsjFnP
+C7k7Mxgq0kxUcH7oImv4NM5Csu7BUCgdMdqpgRAPR1HeemED/P6TkxYagAbxkw/
tN3bh/gl65Q0LT0OtyhUJIwN2RDrfp7fFu6HcOCAU/cJvIvuUpjX2kjtUJYlHdUk
HB9AwwoonRycN/qJRopvqCJZDZi+VCZQ8TIAhCeJY2V/4kbpDwB0vBWi2OsOpw4n
hIIUudrfZHtIRgJ5BzoBhlmsvRA1UaxlvLVHCVU3ytuCLs8AnVZt4Rm8wMTTBNmM
ZO10lZ6fYDlJW5KwicLuAzfuhHXovIAWAQ3qlbPd3sDksy5JYEai5MhkujxWx0+Q
TqzQLbsMdxpksjsYbZ6QAH3pN0VGTw+lWcFxswLflB11dxMKtjhiSaW7vMw8BSof
3nbYh++Ki1wNdDFkfcO1qpIvQDqxDCuCMKGucD2S4pdhwY0X6NFnJnrroBuRfnfi
30x/x6SVmW1Ln1gcIh6xpN6feGChSNfszgr2yFTs5NHBcXkUrubZZfnDbQNCkMLY
bsw0rP9T1y0wJXBTVnJjiZuh6To4aZTxCJhms3IAd+rvkZCj5ncKsEGHJVDvyV9d
jSj3TUorn+9U2hokWa1XRr9l9QrqSFWaHMeSp2vzkCrz9PP4G2lKCqpiNXU0u6zx
H0q3XpF0n0D9HhCXvLoUv2InbtU4y7QONHACQebyd3Kov2DBpUVO2/Pr7kgmUQ67
NpQIb7Y4kt0bCPA4efpljCcSS0FblpNo031d4HCtK5Llk/EbbuL0N0OU6V6lG68C
NvTi45r87O/I3DO+ZFbP2Vc+FfTdUgO+00ngJPow1EmcS3leItbUO7kmG+6CuKcg
G8BEXQwSZHMGQ+f3DpltgYGfpkajeHXbG6H57Rf60a5cZr6vM5PFAhWlWtOgRqdG
Eq5dTISaAXoIkiv96+0nQCye/lvWTUkCup2nn9KXG9z58DPkPUx6CvwWroEV81Mp
pcvbQQhmup+C8SepMrrH+oLEJZlWFDCqBcl1E2xcDosZa7DZeOfkzdYPS8egUXTm
ZutxiRvsXti6rvRUdQdgfJTmYYWdHbtDtole4kS9doLZShM4JbIMnMWTpqDAuNW7
ABPmP4XDVPXFXS9BoSn6A7yRiEuK5TDa6Q7b4Jms9w3UgG544gAbo/F5zsZBlN4D
Ikm+6PNyUwOnRAOiQdPP8ZgavoMGKxXma+Jh6NeuGmvQ8mXQOuhlRTSVv/NROfcL
6jN3/mW1ZmDXIOJK5p6GdtTwE/uPRvEZh3Qg0SHxCXAY5uiW9c8kxvRze6SNF/nC
MtSxMR3gtMY0TO9y9AI/x5FSztfCcbHVb9Ct987BZgnqmud1sh5WH2bOhLQlw9IM
orNdfTL6xPvFPCQzU6z8tDyrsHSvobGdUtPdsAXXxiRos1+xDVcGuxXY0Sjt5MvB
k+3YauB5h8C5cJXa86P5NgWMeCn6gOZuntD2FWx87M31AUAIOopADQZMCUzoWreN
vZ671jdNv4a3tDrPc7aMsCsJ0fVwjw4TwowjNIK2tgpLmTKpto5zP6lB5IXEOTRQ
WoGaQ8eaGdUL4NGXogBvNAr4tWHsjsp8qbbWOEGJ2ASn36kAykzPbKD3U1zOBIBy
miqJW8dtoAm2OfnDyMcD80rVHNTko6aDTcTgunf6dQP7gJuHq61t2LkAkKWosM4H
honUQRWAG1ME5mrzJUjm9DUwzkcATiceBldKwhkHOXps72WksJ8h7sUK6Mv7rYd0
Mj4pDJlq0OOGPqvDgJIZe1EsECoEs21n4WzPj6AY70bp/XgaQ6Sl7k3W6CStO0sW
XBR18pH0QTR9htxmG0VYjRvObBNnFjrwQa5X5xzgSs8aAAF1/widbjsDILZJ0JHk
dtUjAh5R6ut+CuNQlNzZz2U9JBQrSbAmL4Nh28MfMC0xB/6i0uj9vEwVBLXU/lV7
cShT+/FGx727dqYQj/2VacYZ0GEE+RWNK39HnXMus8N4gIGdL4VI+ApWBF12jkhe
ZVSQLyQOEb6v9IXdv6TRIArXz4maHEVuTm144afXaR5ufXzgO74YThoZmAGD/wsw
8/QTq/DHejBadC/d/Q/O1ffQUgg4QmcpOAYeeed/f5n9yEQZxBgTgWFNcVVAWI9t
mO2piickdwi3J65k8II8P4AdCPxKuutKsH0iS512Q1XgSwnkBwCIo+oAqmAXdOLn
lgA1ejc+Y/LYnrHXhW7+VsqiyuUEnii7p4zFFqvqlQKfq/sZUetXVadcCgvEfe1M
ru/SVnnm0rgglAj12ZEBQS3XGfgrDNtOZuF2B2h+E7ccOP5xwv2exfMQss3E+Y4s
Ldi6Q/ShJmcaTGMR9UElg290dmTw7AD64m2q0qyUXsE8EbQxSRugfZyVA4ptoUmu
+1mL15Y0zDLuBOEaO9CGMyA+27PgGkYuJi5+8A/QcpGvEB2GhUMbqxOYtdu077AD
ywa6LW22PPimiZFRozM/ZIHpxcVgr5JsVFsmxjHLr+oD113KtyRrpo7EJ9hnX6NP
cOkC0wFOUy6Oh9Yx43tuQpZ+8jRGRK5kMMXpxrqzeEpW/jQTB2ypeZMoWnnVxJ9i
8bQNM6CogQbE/zRTnWFAHDUr1kRDvQnIeq3+9NvPswulG+O4XLG+nW6lqLB06l2p
MqvJv1HGWZcup35J9Ay3lZOMVSZvKRPNPhMUDf7b5LO1sdTQedfsekATqn180ADV
HI4suiRVpdmw4pXpVBpajtbHQ7E6pj0fAjFiY+saBmuLV0g7nyQXGWJYXoP064Pm
iyxIvSzCE50D6mud1/z0vfIgL23Xu7PF4hTjYO2A8dNDDeVk+e/yKo3mTwIVVO7J
TTN9MgS3M6upRjvHoQkbujAuN8KFJ00weKHx9/ew/aEBhXL/6oEQDgH32JAfQORw
osZEdYLrYtWyeS5YtVpZh322QDw7pyLQeAhe66V8S7GKkEA34IUlNe0mRyJ/ixvm
mwZJcI5v7C3uuEtt52YRKGDkt8YZJ63YeFmmBeh7zAuhMRBCGFG4t59Pw4+rIPmq
8pQIrIVzUxtE4J3BEumadjw68jE8xR7Yifwr+OXh2obkbFw4nud757gwKhqHF6L0
Ddlw/BulHLY4xnA8bYS2FOZ+yCTgQwlnzkk9rZ78fe4LJPENk3AbrEp48o95mVh3
p5CH4N42AjgaCbTrl+qmLDDse+YgZRkqYnN/p30WpQyIkC66Hf/0nYObdivtPTyV
3bvNCUTmF3wYaBkbinZlk9C9QW4B1VH6meR7N0CtbUoVqb790eiI6bV7idJIGmH0
rKwzJVfV3GcI+eec/rmy3/Zu0Ga+ZQd7y5JIPyhUSwM3INGN3w4GypDVMUcpYq/K
Nnq/sgF0WaECE9ol6vS8fuPU1g5Ylop3RN9otj5IYOPdEFKs7ErKO2EEb57cB+/S
thRn25/D9jJ++2ffQg3W4j3Ps7sdWC5rPFu9EWDfwRA0XVTvExL2m03SBEO66cfV
DKMFO19KfNp9xn1xsYcaB1qIiN7lmkZT9PhQHVHiQ5kLtjNfdBXYHfLRXa1HWlkc
6qUryeTHp6G05c/HMgFvXob2dKT9y9HdKsuG25B4j3ZTQNv22DA5Xi991gmb9KXF
tcM+6+xUghe/YAOO592DQO7Ccekb1kLAWAMyWT9HSWlC6Qc3bcVFPR181QiOziPQ
ev0sRLB5OYBXspr6LcNORyWn3DnHfwOGLviruVwu4WF1hREeZYb/87p2Xtca1n2W
vushwCxWyV/tePOo7Ka6E0K9s5UnI//t4lT4WYbAJSm0DYqV8X0XfF3XxqCwX9Wo
43l+hfNJ1RBmYUy5UN9b6Wm5lpHiKTkLGnsqXWYnXY6+YZcVY/AyKhaE79ZB7F/L
PnINtR+jjnE/QK0XRxk1692Oe2v6KJBMy6lm8S+5aeO7roq10vDlSWknopv/Wtrz
R4r97r0PplvBQFhR83frZyT4G/16L/Gn+pXmP6VJIChXQXPwm3B/hmQvscSvGs5i
QGwskEuuE2atYzuY03vZckj5vCTf98ObyM5qccDFARCbCMtHtdrk+6rNrgfTY97e
mD2EQHzqrOSvM+fWeX1lS9lLH5d3L59VJQ4swcyN9zsoVKVt9TMHOxVk0rWwyd6v
Gk9kT9ecBvEFhdA4AnxBa3QxKsqBo2VZ5BMxxqYomZfPTxYbMZWVNLE7UDcL1/tD
6FO3nic6Wgx33r0yf1CRfBP1z0TgS8Yq2S3SJelomZJJamaiQ8HeCE9SiLRHZ3Aa
Aq5aC2u+qZSmKlekoVU4b3TFIcj4PJT975QkoL6TtXzzEkGxTfFz4bzz6qxfb3KI
5KhL36pGJCMuHS3jtDXRu6ZX3/x5/xyP/rIsqYKO9xOdmWMN1T3WcG/4rYgwTLO4
Be/n4UMWJlyrY06qfbwLonlRkfmytMujFdQ6iN9jCANTfnJB0UXeMIkD+B9bXKcS
0AlED08UANzAZ1zXEnB081jfuQ2pbiT1F4OXJkP0e8zRb+BXOO2optYzmyQoHoQH
zrOzHhDlJ0yn59EBGud7aH1FVgEo1StKlTFqKliMXmsGqwp7i6mBLbZ9gkWk5FM2
rF0VKky8LixcKSOuAPiM+T31ow9ncHW4I48MSf49cobIiZVNRcPkJqprzXR7ivBu
mGGE3H6JdGLHUCYi9IM3k/DOKMLRRE9uBNIu4pSYb+yNTIF4UyBYeAys/GWrfobF
mx5URuLdTjpFY5+FB9LuJoR5a6eZk4QFsoZVqfM9OQe6SzRZ//fJz+f4hixthlTj
9LRixEiZXsgQ5AqJrV90Po9uw5YvTUSaYbNqriyXvUocNZeyZgVscsLHz7rWeEaP
KXc1QmrUbAbbN0oyGBObQ4ekddpLiTwxpPKtnYLy7EFg+8jUUKVKjdCy/0pnp9zC
ZLlhPdgCnH/MOTOk3pEWVOtNMFL8C6qzCfG4cC8TaFwGssMp0NDakjLva5u5qYMp
Lr99alRtxs5M/7jZfDLB4FN3XIAa1SzgKktAWp174d6MnVAcZqEw4YAfx+5TIuZP
wf6O8yXuq7+R6OEw4+ocUVJFD9TFXmq7jvhSxbCEkqVzRz+ErR4D7aEnaHX05QX2
P4IzwDtnGNFE8NNmqZNqIZrAmxbZt+aFNNHYuveTz48UJuq3w+kwSN9UPhvkpgHN
NXxWgpKe/4hll/cKWxaMzdA0NCtpHUBUUpP+1mZvWX5AcYeeHL6fszPdugCcWNq8
cUHR6eRubtXL/BAgs3jC2AV6IRkCCnsnTm66rcWxUZ1dn7igjS0Of9jIL5C1WLYS
GzhelkBNanrj0MhVvxWC+GVEMYe0K8uoOFZipxqcT7fbnLdMI6O0LnISDyuRUl9h
CGeNm7ATAfovtMj5/GSFovC2J1rhdNN84fATL/zmmUbvO14D/Vyo5vWOEDoAg0i1
8OVmTZTls0LEhAUxmu+9NlCi2kFqZtCkknWVjzqBBdu39IrVZMCEdEg8m7B6IsMy
V14z6q3jWOu5fT+vAdaKItacdq8CIoyQIzhO4TirEPWmCR+o4WOd16UCX9C2rg8z
5SfY9EwYFEKfkRpHyCW1v5D4SjSprzh3SCSTkWOwe9kJ+eTcPdeBW28eS0w9D4wx
LUv2jqWHBL9ar4o+45L7Q1+upOlP2pTEnSAwnXoDwccIV98Co661W8PE6X9s8/pP
CYdbJRQdVtG2upKfQann1Ga1y86h9+66aTgh8+zd16n7o7WVZgHUiuH1DE4X4GAM
McSG5Rmd3x5eQS+tGim60p7jbaWWREuuSCx2EoJl3ULNIaiEZwelcWswyzMbn3iN
baSjkHXg85m/EAXdOOBIlis0XXo2Xqzf8WmVj8CsiHn83HWpYrwu+2ESVek7QhdV
JiKHwIqNQSFVj/bHK9+KpXXQnSmiouazzplDB+DyMpnUZ8WyX0DdR7cUryNLBbKH
AazuplQ8ncfCvW/1KFCSnTW8ANmdCIOZ4gLbg2be7FktlANqpacb4LbSf6ko6BSd
bW1iwhcnPxmNV6XE+ow8Pg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RStP1X7Gr0gQaoI9HhGak/+WMPnrwav8MYGP5i+NVoucjBoB+jO8x1jTn9PtvG00
rdbBD78WuamPWL5X8ebYoyqEHFoynxTfH6we1scQC4vyzvn1hIVtBcJX2+0GK+rX
KF9gMFTgzGn56p4uZeWAcepXxsDHxFzR706LwJqTv5vft/0+mQLiJHxzwG9uocSk
QzBqWiMCKbrXC3YdVhPW/JkNOnMnLifE5Ekzocq1olhiNkDdKapOfLqxZBSyp93D
b0I39vNKUQ2DeXNvxlT2HBVTQ3QZirkxMCyP6RreVIVsagqIf0UGS4McDzNyD/bV
OZik3v+ZPJ/J4ZOwgnCSAw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9344 )
`pragma protect data_block
ruEsdQ+bySuF0gCascVuEiNLnx5+GVORXPsmK7HIfseTX97KbutrjDbDhg8zHF+G
SqNwuG/JfaBSH0snu/lDoNLbUEIUp4SuO0TL+QSpC+i6MBD+V08dRarq03whgfSH
VOes57vnbrzRQPKCHL6FjuwcGKbFsKFZ9jDCS7l0B2qC95j6/VoZgQLrRbvn8Hn6
sPc6LwKl/HbXJYwA9qKf94DxLxfag6iWsizqEg49ZvGn7hp4+kUMiJbhleLiIRio
o42q3YFaeWF9y0TSDCNum/2l3fOCQqEUi9QZBM0MmPnH4w7rnG2bk7T6Vj5FmBRA
D+tAcKoDBFL1hajMeO4fkfmp4lWMNoJAdcgraVsdadYT5N5NxjnhFtZhg2Yn3mgi
SQCYfLJfZUZjho/LhDrSZ6XefJzqOEGSS8HV0wYvImCPQ5u8ZeRrfUq1J7zR7Cmw
ADyhpKANKKJO9/QGUHjjH7X5eR1j9JqGu9PqJCqYfpujcp0Iud4wDxeLf5ElGmcs
mUC1BE4ELb9LvHfRMrpnTVrvT7IVJcxRJeie/GPElwTccZfs6vGVn6GaMrLM06sO
wp39ITYsQAJOdAwFcc1T+196EqNDRuWPkt6beWt5OJhm/VbthnKVKzg+8zj02jIJ
AT0AmoWPvO4xDsUrpGXOrKgOEv+ly8iuWypmSR+Rjc+HXc4EdJNTF4NPEFkrkKQU
p0i4FYchtpBJVDINz3i/YheipVwjzHCrpWLw8+ErSf0lsIseEb1SdSqiq2ChtJ/j
MvUdmKRpG7BOFlEBOioMlgATvWyOx5KEXUf3eMLX3WlpPZF04FbxR05JvX/H21/M
yXmqlrEtSUY63C5GKpeFyXteIb1slv4K1yNoUy8791IvT0u5XdC7IbcOozjUtrZL
MRHAYf9ifA8KsQtslxyskBt4cg4HpsHOTWytrI3ZV0R3sv4B4z9xjrFor3vuiW1p
ipycLO+3TvO944Qm9m5dd+OyS6s+Th718B/lgP9CQqJfjYd7FIPIea6hejYUXVRz
UnMMVOEvC2GKVIhsi15nMw9f9zExVJcxZGscizWOIS6CcMlH5miubeccj+C6wyjZ
QduwgxKLRofWH1+LS3G8Xn1hnGW5EHpQtLdXweh7Pv7K6sJ9V9oA4cVAwbafChrO
T8Qop0G71J5Y1pElF5p4rHfY59+eK1CHC6HdtxTFNxVV0anG/y7etZKhr7i6ZBj9
mNkemhU5UejO5kKC90gzR0Npf6YJGVzdsSjRPRG+CX+bSTa4rZKxgnevp7c+6fjm
x0PYDFJEd2SvNFfGcJe2gXp3RGI1N1RuPPbTgnUx1otBfidEMXM9Q+T1oR/jbajG
8uoK2sCbJPucMhBybG6ddmqeb80LeejKw7ad9HtNSVDW+6U8gbk+G8jlzdXVLFuX
hSRShZR5faykFd/4qqxYS8kx4jNEH1ItGfOIR1vbxnB3Mqmv6LgacRgGy8oSv5cx
Nc2TOxxPjJ1YD8qRVo+uGxlISP1Hn7IwTfiB+nVKrjyjOT9rupvGZSenIM+T8vek
1AWPx+QYJtVOfV8LdVuprrRo0vyoIMqsbJlravHuXDDaLY5hJqdHDLmYZpGLzTXG
eFRYcMXO1Q0wdfL6TLPS7McHenS1vms4lAeVZ6iAHAtVaaYnAh16/ynBiqxWagmd
2CIUzxkRIdW4BH0hzkzFy/JaX91MM/FCIzJMBng9kS/hgNjzhfeHPF+WL9pJc1ef
XASXhhc3sMP3g+aikJ97eYvwX/k/LpUV4yPgT656uo2Adcuv2dLYu0Dl66G+FZnl
yKe46e11GvfSUdmZHqdLYu9QoXqIO9gNumXdG4GufOon0Qs1f8xViaDpKhVOVZXg
edIiEgYAkXDpa4whOHNHt1dpz+YgOLqZXbUDdHbkXQ7Nb1c4qDiIWp0J4oZ+lbBE
qIB9W40IHKf4gb4AaZO9GB8e2gNfc1YoWKgeooPI6vF938XKHoTh3oPH4uAwdpFT
falJQEUF/x2QoAVBrx0/Om1CARpKpl/X2NKzmvEMqRhJilUOo8flagAu3nYd7ILL
BdgMBNzsBejgbmGTmFJFRLnJttxaecBIkLwnE0g4OJ3xzTNlgCL3KMyWv2R9H+MT
KXDVfnGbQfPrDFtoXb0gAj230WjQqJLj5ed2waj2qX9aIt8YjXB2J2MxL53UaP/b
Tf65OmOaCkX27MlljA/60tCy6dB2qgot+kNrCXt2tqDsRio4ZfWeWxmup4HZnVJG
sb6bcgt5Z9/3wAP/nbBEoXC5y1i6zJmp1KKahXCNKLSVHAhgCQESVdVNFYaWBWZK
NCVOQiQa9vEoIEwhfMBKKyZHDl/MRO3fK1hlyaBgNannzEH43A9vDfHsTO8x5Mnq
xUT46z4RDwVNoXwjVPhBg+TQrFxogFHM/kqWVtcp8g+Oz6BOGvNbE11fXzT53nF8
xnwabs7llil+SWy4vyIWN/19T9laj44cDDf5e6WpFMnYkZ+ew4dAsKLPVuwCbicG
jfBc90zRfzCOpDusnMeodD3c9GXd0ALS4xRc0SEA3vpYwBCbJHpLF7sfASsS8NQT
MC1gcrG1U5qOkvuUcTXjXHKiEthv8CqlUShj1hMxj3oCx+4kSbWldR7CG2y8Ac8A
f3GxTSPYyGG54q5Ldh8GlUqpX/HjbmoKYuoICcgcuRkqgHCBdADiTloq1kFZ8dEw
CbLRbV10K/yudlV4XEyn1KQLSh2hPd0274bcwWb6q4iEmOZxJKoIS82Z8fRXUeWq
zgnGA4pq1Ujs2GA7dQWCJ8aSCbu5VHnDPRmAAPgi9uxHTDdyFHUK7eHwkmTuYaYS
DL7PgGOguPH7iCriXjDHtgwt2BFP26Tc6dtzfMn2YPjmPndBfQTU65aO4ZIePrlg
bQDSaagyebLiywotzl0OA4wSGj3Z7Lv+vF1izi0ztKipmmNC59VbQutSFYOwQR2Z
hg5lqt0aQsBEoxuarScPOdWXyDZX6bSLXLnTgdTblQXLJdjw88Fc/KheelGdYXfm
4pGT2aD582c8qtpaO+ymqQurmxMd2VEcjbz86JPchZ3KsdtgMdg8JPMEkdE6cxD4
m1p7l3xxK4J4VGWb43JMngqxv7S9Eo5zOIBED9vviWNS2kxKN1RaZeONaQTAfcS1
wYODbjcBORdUFWQD1CW0tRMRX7hy2LbyzKlSe/LUSX5wmEALLLsVyQ+4XIrR85ew
/CD4Pn4m4oKhBTgIaCUqlLzJHitlu4Rih3ghdmUPu1XVbwjiVcAeKxlf5YYc2nk1
YLfdj1ygkFLmR+OyAN0/Z2y/ZgPUeLgK9KazWK+bVmAT7iRo+zdhDxKFAU0QBJT3
Q1O09SYXWN5UqnzqhuOOEb95ja/zVSzvfbipSoyXc/ZZW6Lsd/CEYZReLgLlBZPJ
PwC6TI3QYVv6WTHWWS3Jx4mPhZlEMpPD/CjnuZ2MuTkHf9IFmCxKNTkhdgyq/ygZ
HC3LvafbpXgQCgQmZOFGSNyb8yfrlxXDC53bMgZx7vOGB8X2ScKEG66HFVGZcGCy
nwOgTTGgtZmk7TU1BJA3tG0qon/x2WbgaBywC8//jv3pfJcY24k9qRlSLFhLfPoL
2g8qbWHhG6oJkVS50+S+aFofjte3BHYTaBwCai4xb3pjT9uTfeBELdy18EZto39w
Va2x+7eG+zrQqs9SfqHVsfQycN4sufJgmQnbs4wkCKJ8iQWp68vZ+ojScxYQs7xb
oNofVk6oE/di2SfP/vlbf7ynoJTahkgOCP0kxweG8khpxjxDxK+DLk18jRAtSjii
RipDjkh4FT/H+HnuwaQh6ShvZhPrYIu5MXd2l6oyyjNMbWjRWMPQ3PppGRDAemXt
7Hu0oMywknF78ApLno+imRjwajjAFyn4ERFLTAE1CUw5G0uDpDB5pQWOr6sHyeL0
fLDaSQKUqiwHd05jDnn3Rj53wxOFBHl3rCWe0ev4OU6FiL7S7XsbgJnvucIkwdup
HOssiZKuTKki2hQOol0eI1xlUQPYRbEqhTOpL+4nifUJ21fzC1q9qiiwqREy2Fhg
Juoe4WLlByQf/cY44erkFfB1uVYqtLrcVAuu1ET+uQZ0s28Rbx9jiD5o8nXs8EDY
20jck5wke+5zb/h+FCaIgOLGv01gC9ItYQ7EgiORvYfP4MvcaVzJscjTQpQnHPkR
+E22u1Er+ElOv5t6k34IRujKVVwxr9bZF1IVAVXjLNrsNC8Y/JyB9AJ1St2N0PZo
YVAlZGCG+BZexSIqBsZ3OhK9QEn2+dcP69Jn6azofrsL+eoNQkXxZk6nE9zxSeen
UgIAO5tjDLxuSyomhZSLBKU0l/da4T0dpj1HYCEDrWId8tQ6uaADcaUODvWj1EnC
XS4YXzN3FuWSrScjgJoMYCfxDETL6cqrsuHabGSPWN4vu+VWknjl9YDF/jJMPjVj
/2Oy9xRu2PMt9lm1+6XIuauYHqZdqZ5cOidhzgGrvhYBjxohZQg+UNqAbjxNuDUV
RYhtEY9i8FKV2XtpdvEjZUYfvLDpCSLdK7bonloe26jvXcARCKt9ZFpeLxM/wArm
44SJ9Zkz1EZauIVPtlAbt56SVbon1PsEc5V9D1xPMum1YbbR/bSNLqjSqghnwSzI
fdqN3RTwvJ74t2WuUGMNZ/hoFCkoLZBd/kyQIYIxNi6bfMKFff9Lb1cYbSywfHsT
vrmH4eG0GL8grWx/bpFpmP8m2gI5P2+N9ydgGQbw6g+tmUtmOo111M52wocBNGqG
LLIt3+BXksX/JyCYvEUWIVaR8syQ4gejQyYpcRQdJJBc0YKMtpGNi7u4jLUxQJkp
GXj7LvFkysqOtYUtbhehyN0BliLLbTVPMNzHmOoKkB2q+k3mm0SSCrxLV+2G6eWa
t8/yQ+d7JKE/6pNJvJ+35FOUv5Uc5NS7ORSFACUf4DBtpsN7XLEKsPGSnK0SgIZ1
ewCFk8RTLFxgSLuwC2RSq5WauaMXSNwCkygl8HMaTCtr8JtCP90BvKpmWrR2k04f
H6DmDuOjkW2FGivrcMIf8nHxRXEiOacovcLFAzkGcfhKPprEYqCCtjHYqgU08bZT
u5XpqU//CkfmI3Yf6S3mm97QFjTZjHNfzafPJiKRKSypdsfsGMpvVMX8iQ9s+jeY
BXoCgQ7ZF/R/vkk29+mJOdwI3xf7rU/CSa4bVUbvAb4tiwBobRxCiHpxt8ooSUM5
eXC7vKAlhzRcrxjvWKkwylji//EGuY2vvxlWGjWC1+iNKxlMykBLd1ZqNWkdzu5+
yPXNnKjpJX9mqS4M+WikbUfbU/4OMdAwkyJG9ISCKKKCpjIyJ268JIR+M+wL+svi
WWoNF4pycGdyHWk9xdyiaatwTj7x85UD2LblMtRYWFgt6Xnce0uudJOlcjtyzxls
e6++mHcIPlWODzm2BfkWcxRa+hx9XEkQcvx4elgl4O3Yde9ziSi6v8WniD5NTmS7
CN8FKQJY5LkqaxFTUumnCe6wE5uFolTD4xc9UZBnAiOkcyD290Gb7p3qoDM+bR/y
GCzs/5A28yOHltD+4QJCCXMl+USDMOMN9IT4gB0aoi4rLAZfNoSJMqLHLOkR7md7
cNCcYj/l63Q8P3p6GbEpugUmbhlFIW1LKETtX3beyAUCvKv0OuLXtyRmTxQCenhJ
NxomTa5Lp9FHVtD2vHf58AgwkufTZb9OzOjBtennjFkQel6oQ/ma4AoxckgFEs7X
SQYOWrq3JzjSqBUcaFuTURxnmLpd32gwu2teuP3rzNwwc4J3gRzu8aq9gs/IjexK
wG4cJy4kLzdZKaeyxbZJxcn8J1UwAxpdnX5/jW+BzM61BSueyDMkmfAg9M0eCPdT
wOgBboB1qPGtQa+MYU76kOckv+ivw5NcbMFwTC0oup10l8goKjpsi4bApEpuqbU+
OcqhTGUiEupjLbyqkP3jJkNdh9jUkL1TbcHufIEkBNc//AbrJv4gq0Pl1XoSvHRe
6+OCxsHajfueJ10hqWIgaVRRzN2UeOAOUsYX1TCqZQ7x815vcIu1D6mrRUuDt+bO
Iu5oaR391oWkyRzdVXCM5ZLJEDwQy746G0mr5OqLI7DIf8yuevGKNE52BtBIJfOi
dqZoEWayu/LSplNxk1WVPlOtRIpONAowWGxhQA16NPHYy2yS7FyEyLFL69AzDKz3
dRgHYB1ZKp9rNWznNau8rdl51/HQlKs5+2e9Z/UMqCjctg+o6r5Pfweb8xiG2aeJ
UU7r2QsSv9uLiZGwH5Df35R6rdJ2QPU7GrOT5fq0iamm9wpjeIpATs9Ba3ibeWGc
9ZKyPdEiSEpYtzD8/x71RwgdZUecPc5dJlIWGW+EZX6rxVTovdSguakWFNiQRdZ5
s3GJ2rVW08Yeft/A+Ne/B6C1O0C3nupMqH1JmrgTgVGqwemhyBnmEI56iuCfygIH
G+2kG1vpHjoOQSGjsX7zRlAQpK/++drYvnLh4I6ARnYtaaFG8/yZIWFStfR/sohw
zwefZxj3HodCshyxjJSBHQZrenBY0Y7D6p7DzFtkvaGJiYPjhYY+3kyZWDwxVsoF
/mwljlY6R+cN6Wr2fiMc3hPpKPXvFbr5K+6U4wKHO4oay9Fdt6DFHLeQ79m/9FAT
r5FTLKelN57Hs8j7g++A+Dah3Nfv9NT6oOXm+hhtdhzF4brBvSvM4oy1ZcIm1pYw
cuWFRH+MderLQQcbvzRmKAo8aEYJRPEIvB1X/O195m9GWcsqH+FFgLfjnRsteezi
h+j0dWWRLk9gU8s4opWXiaLnZFX/OVwmQNYuXn5x/GIc8iVvyqo0wxG9EeN8oCKI
G59rTCNjk5YG00VKBrzdydc0ndkh3ZuVFdEMcd0eKUWLfUSryQAHDH84OwS1dWYP
bsCzQqcYN6RtZKG3r500rz/u+/QW14FuJORGuGpkCXo/GtWt8nOokA5fEfvVlvKx
lOw3BnUPOTmhh/d0+ucmqG5PPZRHMAqSEe0Mdd7gpH7Ul8CLuk+LepSUJlNZdCm8
9LbpaOqJ1rVdlvgu1D1hYJ9u7eye7DU506qRsAJ0v8id3+SiGTjtKpnkm7CwDEIG
5uet0z4kG9zYm/61EQfd2vrSODVNLNu3IDGhoFLtZ7+vq6qCXbfsTVMsZs0R2fxe
5B0O6ICe5Ecm82t+GFLg6f6mqiwWpxiRDgiChc8ojgsEz/I4ISLmZJMd1yJrPakC
OdIQ3WjipWfmJfPh01/mSmDMsnIgZ7kKm2WoK2wJ3/qyyR1Z2XGRaD7eSwwFB3yC
T+47U8m4V2F5376Breavcf+ql020Ik3G5r4URElcGL3aCcUjWL9AtcJwynWDHdz4
Axi+ULCDWR4AZt/IQmV+ekJBx25eKdMFrrqvQwHheOhz1aRyyzSc3kr65+1spl17
mH3Yrw2607XitL515XjbLK/UjeOXdT+ZKXYt6jBSYKgnYKlZ4XDzO8RySOLeeKmu
eR3nEOUC+QQHUsI0xmgatWEQc0qRqhHN+kDchJV4bxC9FeYEBeIL1lWwnnh1uGl4
vO/oVnowTTG5j2e9SjBOtXEiD0EuwY2G6LJhyQMg5aAaH8GLZDlhl5fOiRH+VEiX
SCmgZjaVfCtnTtSjDLRmzlmvyFXMIjGXFxhj3J7a6jVKxYH5IxeCIdKQMvI4tBUM
Xz3IoEDRbKiHCx6Fzlld/qre4iW4q0gKLCLgbuoGDjS/kDsxSHZlYAbstclSj9U+
+FkJKg9rf3VeGqRPhFCiPvn5Ev2scukEIHmu5ZA6pTVbkQbF8NiAmygKAbmOVwMk
JLeD2Z3Yb6sfRCkasnRh6KFHVvcZ49dOy+P66J8BKn7EhFPIx3+oovWLdCLNqSeB
PIQnJBQFiGD4efmcwm35i9B42LCgFEVcqNk4C+6P55p1KUyLJMaBKge9Tke9VGYK
ffLPtfPHfwrhdgR52VirlEhbhBBc8nNdJssTB8hXZXDqn5C6lGECYZRbCrPHgz7B
B14zn/MevFM27e26CddzF9WnLJrdvJg1NMEOf3Mt7lB3DqQ8rS5xYFt8fobjokY7
sYLpz4L0NLX6ovTa/Rcw4gak6k25F7l7ukaEDHHEQdsMYbaYxQ9a2QOczVfrbJrd
CnbxyiNz69LHsQ51aaZhd1wFXNRAINew0zRfeYfVQA4KeOdwiLs9dntzsnn9JG6o
WWjXZcHUSEF8YUlEH6DD7FyR1SOgoSVB0XSHBVtpBWfchZUVGdj/PkSMxpw811qX
naL8qLKv/Gj8+IKlSDqTEtkoy1DA/2a5EOAlRNRg/iVmuHB59NgKkDeneQyZ6DXk
39LwDrKgJ+B58jm6MXDYXk2vcC//kS0E4DttFbqmL43Mw0jDKX9s6OZb3XdcR1ZH
MFm1m/0nzcvjYBMhkElSNb2VNJJH1HwAe2nxYQ0dwCMGo+jzJLknu5ETxu9hbHHb
dQGZoxW3fBiRzHqeU1U6bQKOBoYD++5fpBp3veYvYITR/rHXVKfbP+vX7ohenTrG
TXRGnWVUS+W/HtxkkTZP/cU0P8HKM5UY7IpsRdCBQnt3laQQrP9jZ4aPj2kyPcDg
yl9hNybVpiQLqSnyFRwnRjmJGVdtuHiLw+zkciuEQbr7YiUdBmkYiTdULSf69WHG
hh0uEm2LZgp2qzf7WOEvjrX38uXMzyxtRGfJqz0i1RXJWiqNAHCNFCanC682j9Me
tvURvmpelKgkRNNMpcrtC4EbodMdvisrG68BgumWOYfMDZ9wNOhBnfpL2DGD78E3
3XlfbM1HqUzCKEo15gzfYm1Hj94yg2VEBV+UFjPfCb4j1LlPYSRJ6fS5HhLJc+4I
QIELzbDGL/ofr59UUAW0mqL3V8vEedBcqlyAx2KWJqMj6vcbAUf4Z4SZYzZetLeb
FIgg9HZrninXKKR+XqfbS8pWUuRjLQlC1uf/i16jIMRBEU+UMksxNToxJInuueNU
tOo425PXLERbnNFL8LXqpWeasfXb9Nd3uix9QDsG+6/xA0sliAm9kWbfGk8NogtQ
Mcoo0WfqOegJPiFIxLa+0lUwizjz9IhDVJ/e5ojWS1AmQqwq9/OZ6DK08lZHNog2
jjkxM6DroVktq7Q1PfsIz6A2RHXV1E056MWwMLAeQhGpw6CWSnmcJxW8+GX+41Hc
v8GBqm7/Gcy1k+hVJYSo0O8c1yUq0OeJeKnMyLLWUd25L/L1AXkcTj2CSc+Te5Hh
9BGtE+4pTsJ1VWZiYqF0LnBxf1NSLLl3a75Q7pHXwDhI09CqRSC4UqaxLpXR9SVc
Zv7ATD/rGCbo848UovGxjwmMdcO68kmE+7FmdU+CujRDi2m/5oLVOUW98SBcf6EG
SI/YrDzHfGB8n3kGHs4Rwk62Ntwsh8B9YmheNCHdd5le18VWMTYT+oPK58WcKvsY
rfjj4fysByz5QSmgmF/5HxPIU30ckoeLwhLYhFcx07jdGTHn8rAkcl/8PLztndse
wC/qxQdsZbSYu89mb6JicdYMB8+F4CFw5LqwZbZe5/pEjbQC9RidjfQ5Ie0IhhZA
RDSckNcOvEuLIlF4LvSLGTJboC/bCzmUG9UT83B/WlYEGTYN2Zuh92oohG18QmwK
mf+h/QvIi5hGcJLbNoqU/VCg9nEpV5I/jhXxrtUt0CbRJM6XRRR/qj7cvA2djt7n
noK4dA1mmLMtTnNz0i8Xw68Crwny93Mnsf207UzT8SKGMY51na31DEQYzKy1UysS
mAlLDlKKyuKRjIBCNTFC3GHRqjm+muxKcSNunkSR+mp2NZ7CQr3EX5BoGfjGzcMi
vIFtHq2K78eZN2G9sQhHCTg3wFRCWRFe1jR2Seh6+yZR3JrMc6jLK1E+5yN4TDbg
5XElpERlLQSc72GF7v5+btzK/7sLGF/fqYU24eAh+5SpQoNcGYYSvX6WAiNbLf/5
dOK1A2UuF+VlsMSrNR7Az84LNWl6VqLeU6RF7OQuJFwnZMH9N/FidSx4ccpkQshu
rKKENeKhDG7YWEKeJ3yCBrnDeJYccx7iNBim10GZYxfY4SSIfe7Gkq9wvf2Nuz7B
QoMYTKvHgdFctt8Orgbgsaivby30GIc5utPeHwIYhfC3RuC17p3U4+LFfoaU7Q1U
e3UX9gO9sRkYufn3MtNiMgQjI/G3EumAoaNWtgbR1dOkCoIL+j9H7NMJO1pgRjP7
N6DjWzsjSzthoESzXq0jH1mgl27EeHuEa5W5Unf3hEEzOjaYNTCrjG90o5LEgWr3
LPUKwoeq74j2PUlSTSgP46wfWcCBvmU8VPtYXg8NK/HfmECMvy1J6p3tFm4bwesp
iORYlO2B078qZ1+dpe6ovDMFQbZ8sCRWe0wyhpnabAqqB+PKCBdGTHh/VFVOrtKA
uOMe9ripYNmKYRAAzC0CwrbmzHY3hCXKMrYm4QMTPJ81caXok1xzv2nGKNbrF7DK
uRwMD8K9xxbFbEvOl/t5NF+IryZxuVulh5XR0LHeE4uEZn9Bbr48V+DTYWU5hg1n
tu2gnf2hLYXr4uvwugzOys+tdkg7YbgXuEISR/wpZuUt8DSe7dz5AbvboGQ+v0ce
17UzCeLQoA8GsNcDPMqnPqU46Jm2XVxts2LYM7COjWEnH2Vw7lYqJHrbwDj2uw6S
EkVCl2kiv0Uxvk9YuARn0AbwCsL7z0b2UXXe78FNzR6R7xfCpDl6DbGBYHq8CqvY
FDKff6EHtsfJDM6u1g/zPC1D37UNad0qoS5A/DGToo8S2dmoH+Z+wL7oiHQjEwLn
UNdn//X/iWjLDOwg66yJAx3/aO+x2tetg3GFT9m4Hg5qJsigbzHJo9CX9/muASDR
vaHh/DQ3rgBb8djgpjgMTUQHvJndqq7IXpI2Eb8JvKgPZBunGTpsrzpPR+Tc1ux2
w/lRw5nNemagnxw6rVEJSGK4BV4v9KwQrEOugokMP17vf+aBBBrCoQtpSjguru+c
WmLsVtFJAsb6YjKLUng2EA7yK7hpt5aQ/fYf6KMOmz0T7p4Wg7Ca3nyRrh4PaqBR
50yAGC2nEedFTETTnZa4iN5pS01UeolhiscPCa/4dMNeLo39BYQiGK8tD5bEVPWB
Qs0ajVqwBzwmvXzMfOnj9Io61c5gCmhxkP8CHhZfQ4mLsj/2AhRotkqTXEdIq2t2
9NGNDw9BG6ibXq0u5ckeG82ChTf/i5X8cUWL4Tlacl5lbD7QwgP7ZAYODsm+DPIM
yAT38ktj+0CyjuZ4lMpLdAE0MQjjjbpJcXUAJhQgeNwvl4acxuv/d1pAknS6Ax7z
EEfvRuj8eAWTiVsdyV0CUpLNowp+pBKRdJ+8Mhfxqq8Bwk7sijtfAAyo7aRKhJmi
KtK2fpGbCC5KMiO1J0yM0vbdj9B2ErvLybmC7ZLiexuGPgdIQRj2SA7pDnH4ZR45
iOBFHwA6uaIJjIZmPWSfoqGcmEBhJCX0U+1MbhthHwaoFPibNVW8T/2zeEBYx+DA
Q4GHcBp2UgHQf8svDn8KIlJrIQCftn397el6Yb6Zos4WCJWjM201k22o2vAlDk1Q
Tg4Ywv6pBduwqp1J1U6CLBW7gPZGjsPbskAjquLpwi142YR1XBzbUmTGx3t+P1aL
cSlkMBVZav3Kt5gzDcDjtPd96TQLBrGWZFYt2RZV1JxmS7FancmHsWVeIZTMqYMx
RQ7uhfZ+o1WCpxTsjd1HOU/36atyfRdLZMyHd44MMyIj7dn7CnWKyYfEWS+PQbCO
JXgDqb7WGSQ/JCj8D9ZgfyNTkRlbUSOYyxdXrwxHH/QVoY5Za6+nHk4ZbyqU/8/g
E+LidJjegRcXdjoHNX97dbv3K9a1wf0cF8bOF0cRf/6UIVG1yLTEz1Jy6s52EsuH
7opMyD9OQjM0x3iXcmyTzibA95Qk5+ODsFcRyzZFVesXHCOhon5aJTR6meq5uj4W
umpkdprUVE+Qdxhu2ZMXppDv16X6RAoP/RNd4GKjrvqAT0lU6wKW3KqPTHlVvolf
QEhxYQ5iHoCX2JZIfD7W/WigNOeMW3xiA9Te+AhNcUD6+hAcvknqqCZ+6lboz2N/
V1EhnIuRCGozaE2SkRNPNUkA8s7R7XrD4tT8O3XhVzdPqyaEV0DNmdIZzc/CX472
PxJAI2Zh0lFbhcgwEm5iCr9Fu9rycVtbdPLLAazPtupxNdkoqNz7hD+OfSxcA42S
wZxX2zJgqhNB8aPnUGanY4ama7Ih4rpcnU1ja5S3nSejBzqpX2QrH1NCFWvFGedh
dvRhoUOJDvvLrpoHN293ZhLY5yaOlSBfHYAd3nM0RRvqp2xbFUhLi1pfjxmQKMcS
eFzFkY684/agTnq/P1CWBRtCKcbWaEA+E8cA9z2ZhuJsfGW0DyKPrBQ1cW+gKqIR
vAlUH7ZhVNFuVHh21HMQQcrVAhjpEAHXLU/uT4zT/2+bmUtaLOFo81HRm39qKpeG
kGZEv1D6UCvl6pV/zmgZlvnmJ+fMrLlo6SDy9PE4uv3lZE/wA4GQgqdo4EU4fi5N
VSF4yvutO9NMHPS1I9JTjF7bRNXHyHLUVg7/1QszugM=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ceUNNWMJKFZ/jat+jc9ya6o9UcFPi1vkosl1hHof5/dUNHHMOFSQYGxzXB/otHvV
zym+bFvUR41WgT0jv4LeDn5i5A9u+RqDWiqZMyP01e+k1lKdsqd1j0kAjzq/DaDi
Hpv2okriHw3NIktZlFULKD2tcXMN7Qv4fBroz4kPUf2BDBKwDZ+MAYRu2VJj9U2l
7Y5J1SIniPAAmAwCROR0MAZInycevHVSGkAwCpbNgoVPOyL/np92VjXi1WgZrL4+
RnpnkwokYGsyJUWBFwtkZdtLzjD8PjAM5N3WdyBjHkcMRxsXpK4i3AM99usTfVcA
6MtgX/q1rHpZZ5aWvH2taQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10304 )
`pragma protect data_block
9z6Sss1DSvX0K+A94RfpTg7L/69lXHLmoo3zOBQ26VxaDJozAqvQSGWXhje7GmUF
WlIrEh6Y618oHftsDJFbfWfH/Xmu4s8/us1bIfGTB8OVUr7xprsprCvp96nhZqPw
PfeaPLyFZXcJNtLtwYuEd07wGeDjyuyDaJAsYpEMetIrPWyX3PV06NjIM/1cQq9v
7w70BAeB4QugZU4fESgSjWso9/L09CEwRPPWbrt5ckThzox3QXy/Chk6nSUdXoux
n7DZcjjslWIucIlxtkc7a9OkXH4txQWtPQ+Q3CMQ0wkZx0IAS7/9niRHUksvIL0P
y8VchwvQkMc8ypnAwEnrWhAu0L/3+DxU6XaxYI3uaFNxLhl+46h8pf+QhIaeJLqV
s5Qrwu/Ox47ygpoBaspqkvbJJQJj/61QEw2IZ7ISV2C8vzthlawJpRE8l5118zIG
La17Y0WefxE6R4KmoM2S2OKuKCvpFV6DI4ur2gk/bfjjDQWSjhwTr37lI+V8dh4X
3whpTr74HlkbN1WgR4H2tYx11FbKF1NmnKsUZ1+ZbX6/qtFPOZ3rn5G1mrD5PqS0
Fv2bWQrZCvcCx/yXRxKJY7VzVpzhnpuElws1yCm/JUlqX7rx1j2H4qGsMkUJvd5j
kasYDnc4JLYbaKegNeZ58XVkyY9+MGbb71ZE3Rl6Cnx2BdOTYxRLN9n75f8B5yE8
8iM4almdYKn4V0PIse3yfPhSLy2ULxoK9IoT7itgv7n+XQfcJseyrOm9n4OBAKKe
fiHgetZWc8Od18Ey0/XpvQfdBDNtLjJAS3Zw3bjkAaCnXyYcresH4GY9BryAgYex
HkcejFr3W8LfwW/54KnQRBZ3rHQ6XxQ7xpkoREmOMeUwmXxgzjFWEbV2oqyH6vAr
xo1tNNS+81j02/v+TeHrDwRfrz3+D+qbAzhk+H/HlcV/g6I4ze+Qfisq1E54EOKK
Uyj74UDOKiIosHHxMhPRkwZzDLRYkJ3EP0KNJxhjQe8RbP8agX5CMNi44BjbbDPP
jwNRq6Nmc05/SNKAxaWTimCAy+Z7xbbNGWY/uowGw1PnQPYfc1+8RHQWf9/xYzB3
BhvsMLhn2IcFTOp9E8tjEd+hjYnPljhmkUZ1wWq7YLYgtv6+bw0bkBphh4ykVuNo
un4FEKk3azOij6FfcFodP34BFdhI+kYntKMmZDTD8Y3f3s3rlGj+qg00G05B7+Sg
YyVtvTl7gHO3c7uWTrUke1LX3P/wU6yI/NjzLhlVry0CiomJj4L6xUuFtbnKoPeK
TNgT7Ug6m0VpMKsBc6t1tXQ+sTWW/iZxZZKxbX/LaNhaZ2RW9VSYvEcEWwLFpkj+
z0aEmr1Wsrjg6xjxAIC8aCEBkBCWueRtUT+hAyg8QSxG7PX9TAo2K+wO13S+JbJp
wmX5/8WQPilU6zJI/pIrvFMVTeCjy4totYCp7DjMXCuM1ChVlFyF1cToC02BxPqd
5YXBO0AWyqZX5sSlxXY4zkIxtiNXnLOHI+FW18lOcu2uwNkIrRcupu2142++mdsm
mzb5NI5w0AY9m7JDKwvYD+nnd0fXvZtkZyYvVAc3WQeipirrMfkqNOoJKb5sy/We
tG6BjkFmt/NHGTtxmwTySaKiBCas5IXWbREfSqIymx5encHTwrokxu1SA+e5pCEK
brUrYxZ9WnYpEbdMuhjh60fxHnGlO5aFj4XbfpNTul1yrOHxmLFsXlKwNxx8fzwZ
PZ3v1yi5b6j98Pip9BU0NtnjRIte4jR1ILvUk83Bqw5JDiostyqE6d46abODUmbC
v8itX/+agTyXXFEy9j8KPua6J9QAk6ccHe80nomgacgdrUn86wuwadH9EEFjC0xG
7p7YQmSQWCDOTM1jRi1344cxgJrEyO8xsy6KhXRa/IVmVqtF0jCVJhFahdGvp+/Y
ZKYCqI/jrz/4HmlQqVLfBviIIYaOitQ0Mp+aJQNxPffXjI/VK4lyPK+zVboaQAms
q4GTwDcbthZ9kyhjpk9Mk7+7+3EVP8g57DZv5onbLIsYHfjYVMvslD7L9XWrIoOy
/CAnoMKPC/wPoTgyD9hcTtlKudmdk3IO1Rc0FRs9KysOPFDXzd5cmz7AZOq8kHqS
Q8/izdzzRGBrQBk7TdkvVk1njd80rg/2ia8hgtRjoAwXRPuykTvUxVxds6rramVX
htfVb2hx0f0ypj313McYZtfKL+vEEyXt+uZ+dm3zdj1MeGIH8N0/TTuGiU3ZvOrM
hvDOCtOaAovJq4kBjoQrA/rCNOSFA3frczvjqmilLTxGBk5SbL5T7D4KWOPe45eC
jJ6DztTMdqNnL2A4zLoj2gcBTJscAc0PsTVRS5bLE3Vhe8xjt/MawlkTDZBXhJnf
fJVykYD1dx7RbgqYsdbI2dxAq1NJM1erGc91+mAl6NCr0j4F/H5HbT2aX5dVsBxl
dmd+vUd9p4y4eRmqYsdRA9NiLsDB0NVacVHkHYSXTQxQSjbEDABP8tpiII0yRwhw
tVReKSQBoADSHqNXtcPIpMvVd46WKFGL/xmuZGbWbnO9veKex5sntNHSHgsJpSh9
qn8riDsEZpQfwp1yT9aGN5CRYiaeac/cy9is3nFtAc8dbJ2FMnRam3hhJIZ94nqh
y8Nb1/SJQZxKPYjpid7TsHJnfyMJYqsrT1LrTltlD/LWHlLzRmBHZHgArT7/QWGs
1BmdWjk8BjwyHXGkdKTW4ecZDSkaVNfpmIvjcyta4EmCpdYhKj5aIXOjtcA0D+gx
T0FlzzN5JpEY2KgGKTC0eeSvUtg0P7e39KHMPX4EFVJaPTkgPzDFKyV3EV6XR6vb
lyhhryvKU8Zn2cWKZP1JS7KQgF6pi8ou8fQ5GCehNTtgJVTElUdMhJNjKMPS5YHu
RDR218niUkjemHdsHNz4LH3S9CD1dKIIkfDDYBLDeVxscU+LO/3lFEvqEkIhQ5jJ
SMiR063esHThhtfJpMqoDR1d2UCmr1scu6PQd5H16TpHnJePogi4e1BZbau0SCkp
AirFEBzCqS2sESgtzHdR6spX4LuZtMKRRvrTf5oUezOij5CbNgjJZoexBF8TNy0b
EgbLuumaW/NIJpP07S/5nH5oHflQ43cy8dirf5N8WaIFZ1RaHs0LEAoJQa0CY8o+
TaPTCBBX32tjRutEGjLI/E5TjZ88jdjPQTn7KnaYc+DtoeCF1LrodZ+kggpc28h1
rAY3EQ8fY/xy6Rt+Ju0WL7kkij8P0Ao7G3dMEFmt7jnt19GZaFTOQ5v1QpbzrIkv
h4i0W20BpgKMMBDrc5MPlVvSMXunJoTOlcdr3DIZdQueOOAEqfzSy2UYOmiu5qb7
pSI9aWu3xCWxVdCb7u8kY65Oa7CcTSd+PtVns9+QomuDDYXTMSkIMbaY9W1c+s9j
WOF85Sl/SwB+loWR5xYQebJ86SEnCIpAx1celHWZICYYb+qpv65HLwrkZZQl5bfO
HLPVN2H2+Awcsh3OOZZSS5ZrUiJBxB/0W/+a3kUvT0VIByxz/e6BOy76ox1gSK6Z
op9bcGYPdIor+pU3o18SdIUGBQEqrF+OT0BoSg0Gz4zHw4OrnbkTWE7YXZZ2DKWY
o4PI4NrG6UW/h20mJR3bQc+IIeZg+iLLTjwjSQInwIie8Vf5mwFDYWWr1s4qa0QS
zPh60cnYTivJTdsfzrd9qz8ZLa7RniS1uwOMgKeGmdEo1EDAFsRTau0i60ComVLd
CFssav09w2o+UP8/Uzu/nQI+oHhz+uHJyJKQP6aBFtMsiWS4bySAKdOBd8MD+FAK
PcqdaO27WW6BKtp/EgyKyb52yrK7//VndDglYlf0BUg2lr6MNIQZV0JNOXJT7SRn
cdCH/6CIvOSzQ/t5A39yczZcf8/awpOlht+CHeNCBlTT0EHNocQt/XACSuTFawlt
RIf8yazB5jGxQpZkedH3lImXzKOh0YIDx8SZD4o6cXKcQvbXD6OvRlA4rdj4gMy4
M8Z/yrKrE/GNeH8clFMg0uae16Nrbt67lymSqP8pbgYvJ+1tS5notskr0bw3a0+7
LexxdElUh+WBy+8cJpdXVGjXXNABhuML7WlAvbudTYQlroC3uU8sF0+snf5t85mH
ARyjF8VEFHrmcaDX1Vk3nRawLPBmeCoN/7KDHNtWKMJMgq4XFKLuv7DGBuTKYrX3
1ehlM2pRglf3U+ihYcqeeoCCWb5BQ0wjqOxYKbflIp/ndtHQ72vYAnv9kJFd9X5V
tt+qIGhtDX0SMWRZCz1HrldhAbDKYyUC9EW403ZxI/yBWXehIZQfceRMfsCBinF4
exVxvX9rFYYf/3alXJA+akIs/7j1mhiD7YTWXL7ceA36I3QABiW3analY0KBSAeS
9Y96eukJ/wE1Cxv7G18xaLXj0ZipFGBwq7ck1VR59Eg3zfNNa/82NZ8SEkP4bKCU
AIAF2xovPCAPmk9vHrBclAZMHv3+XIlbVmrIUh0+kAXUyyD5Vks4PhK/IlIFjATv
lPsiBgvRzT7yECjEhS5ZpuTKJRG7UxX7yGUXwGHGLlqBQcPpd/+rbje1R0PhY9I2
LLBuCjg6awx6rHeeVaVB9dWMhpY81IBgRLbMt3hMODN/0B7U+h8CUxOguYhrn5n5
EwL4U30Al8RjwBz7PjffB4yanGEFEMi9IPimh+5qNIfUUwAIeNkuchfEc9ldKyiS
+j89+s2zzIj87oCrDNgwV6CnrnumHFC9+Hiqd2v9CqqZdgRitRJmlz2PIoK+iChk
aFQRAjxjXSlw5FziB27w8fAyjTN1RRRMAali4x+eKfwEgYnakHoiQRtrHF1tw/Vp
yOMZhmm+k+ur78g/eJ+KRcEfnMifBpl03sSEvsaNAGDIibELeIz6NqWYolZrmZnB
i5aDVUT1qg+P6k82oRJumKGn+BkuJAoMyB2OKNZUSiBFtNxzPp9S6HcAKsc1GCoq
7rQMGOjLS+LCVcnIdhYOG40t10unKtZh1N8Awm3AxFz7o00/oVBC2/KmqpppDsbJ
P+kW9larx65dsoGlv5l2rWcUfdoOb7G1jo1f9p5XnQyZFb0ETDAgQZrQoOkLBoiJ
Bp9nlpKo9HcPwRncD8i4ITYLMIfdvFnpYZ589feQrh2enqKC53/XrE/jdHTZnh2n
pF4oZyxiWnkvxi0eGxckJrR/cyaomgToRTB9oO61EuzeZ3mioKeIgEhrf9ekREf2
xhUqT07dfKlgjZ1Zz6W1+87gEEbZh6q6TJyG8g71iQmUyDptDsiO17L03P1o0lep
emNTFESn0JbdHug8hexOGri6MZURwmSAQNPzZ86mfRrPH9ws1Es/agnLrCf01cIa
RoL1sX8SdFpEyrLnDg6/xDiA5hdCCjtvpZOVicqXHD6gp4q7lE6zS7uJoVpmoeDx
VMMDEMKTtBthoo1/DbLwP8e14g1wVcd702JTiHYSmzrkpZH7amKfZGD/jRdGXkPT
ts+IbgxCiPau+J3OUwWENFtbOe6xSOgOOrnpYYhZLlCwbJaVWmpCFaReeK4pB9cS
C/ja0cDR0SPSb1Zr+eZQxnDHEi5HorBMmkAPBf+BuXOzBPHK/bD2P55AxG1Du1N2
6iZYWBWLnMvaotGFjdnZi7BAsf0NpiS/u6gy9lvu43/E4uS7ruYZuPCXHmda9jqt
S1qXrLgEHzvBaxiODT5pIQRir52Z2+K/y4uCR4nmY4WGbGRn1ofVQGu9CTYzE395
fMS5QygEUzTUXByOvuZlcZv3yR8eMdWRsPPlagFYT9JLv7E60hkkf+tantsT9F2N
1sKpz9r9qbbAXChz9kF88l1Gi1G9k2CdatX/g2NIbU0aRnjVn/rjXozl4U0mg30O
DnOkePFKqid7WqJlKFb8xdxbQWwD8v+rLN0oHu8nZWmKf3EzWLu8B1DcbROfkp1h
kTcXgb9NGctDWLM/HaBQpIMmQkCORKKzcacV6lxP53JNZwyUJJ9hcsP82eXxJM0O
OIRm5VBuIJ0LZSiBlulcwpcyM5rY1Ea5OrOZOownzoiZbOe0Q5w7NzjGRvLxE77m
dAfnoqnpXlNtoWfvIacJwfeEZ7sZO/ZySELA/OtEvdq3OOx0WiVPoJ6eeAVepe2g
XiN2Prpz/JLl+bc/FiYPOOd0Ofs3bdbLt/+uPAJxA0ONL31bgs0Iq48kTE+tPCdF
0TilDjfGNlv1n9xMnzsvHFCghj96nnYbk57zzKR5HKszWYkKl3g6kynL6CEgc04l
mg53IZCbwIq/hgfaFumVyHlwDoFEgyeXGq1II5uYo/YeWP5VMAOQyMZKXb0qUfcJ
F/Ayp8NUYyk6c4x/KF8Hn5G5S3L3C7dFpYt5PA4dr6FYJ9RxAErwMPbUm7sOcbpS
lWlgGKrr2m0oz8VbuPtBQcLQhCF5ZeWLvZCAt5rfgSAgHoF1g2kW3mL3z7mzwbur
Hf5onFhLsQ6LXBXeBtu3TTdIBchtt9B7LXgJ+AIOyzmRno6ceXYUKDIlYkkzZCro
K9mvYokHw226Xms6oT82uv0jRa0RiGIKiOsPE3iJjRAtVP015IHrzPEGHUN8nbJQ
QxaI6kzfcaH+RGKHSwyNZfNIEN4gpqlVa7lL1wJxxho32ZHRVKPymQBjXr0LNYhW
RwokXxnZbZfQ8PEPTwnom6+LlFRA554uKwAjfJ0iX/4fVxaGosjzDReFjkMe7dCA
GLeTtXUWg9Pa4ZMsxeq99hNJeHKZm0cYUMVZjEWG8o35uOyi9YmmQd5E3qTXD+2C
UspgVJTbmAZ9iWHsfpuPSlv17pvjJhu4a7Z6m5q7bG0Lf5H4Teq8TTahk8R7HVQ1
Nrl0SJz8L3ZQVNzcB2SszAX2JyT9LcDkDO1m92s/m/lOOcAtrghaNy0YWHkRTVxv
3y3amj3BitIlJt9MwJtzvitbwRV3I4Bgn7+B0TkkP+bYhbwRYj2iev3e68hsGUCo
w8M1v+fvDc+wCRe4BFTq1UitV5LoCsMIrl4Wnl2+vx8XBHAjQJ+4/7m/UTv+JK6+
NvD5yu/Mj115ifedouT5PXKggih+ffqp4ONCA+GjSDccMllR5t3gmXEawxifSd53
DHgV7YjPUOBkBj8psjuQ1/QdznDSxw2DLpsfo954zGO1uMQLTGWtX8sQmkE2v4dP
wtFOv4HAZmYpmPK9KGxeXPiPsyafAmW96K6JMbq7qq3UQLloWUbLz8TIspVuKstb
BydemIURialgsOs19hkfv5EguIBnJOINPOGam/b0c2GwyOCw12Onsx/LLyU52str
SVbIfJuxKkisrp01EEeON++XEd51vm1KYBn8nUCrDHwFhU+7P6fV9sR2iAeXNw/j
LIUU0fqFEH+JfepTFluLjMPbNYee4JqmKLlGeVw41QPIR+AZ6APnzCY5QlJksPGN
zfyPoUGA6DV1EW+o3uCE2WVJINqwaRQDnnHme0qmhnV56nHv0OQG9y0RtNxll/y6
eJiqgJA71g7odAUuHDd4XLZsUJXFyhQSRVGsMbRmG4IS3WA7jWxNDcoSnAlrk6G0
n+Kuch2u83tir/ihFYdaX2WNcBrZf0TBOUXc2rttk4NoyBJtx8dP7YPiaG6BMKg9
NIoDnHXZsiF1HZf92Zt3j0DiflEj0vBEXl1UJX+uPROGHZo1vVlhoTJkd5mowlYA
pFnKVv1muN66lo71F6Yc2I++/QQVhSjilTTqRB63dTCG1b+5z3xfUgEsJxENogws
PfpVHE8D+fDU0yTXgq9h2iRMIxBigoKLyD/tPK5Bnocjrt9dfgyVCkR/X+ZqFL9f
XvCBZub6FBYn/FoQ4ZRgNQ9O3jTHVMTmHMTa4yuinYR9aXbUgxycJhlncgMpSJOx
1WwQoYcKJZdJVd4oEJFWR9ick+xbuDy8DhnudHiol79WnFW4XhMCWviN+rxzxTHu
peyO7PPy1vw6d5jTHtUQbH1mjG6n5GtBxK+MHw4L/Ma480kaihaCwmArXEbiVjem
RlMVlGPGPHdDIoWwqIYZVZ0B+hJ3n4G44XlKD5F+J3FYEANr7vVNJBSOmnkbdGBW
uv8TNnMqYZkNsRYWXgNvpOjSzSd50SeVVHLB0fT3cG23dY42s6THW+NUnRcdpSmq
k3IqHj4SSbjeAkbxEhTdF0/HFO+FNpX1PIAr3VMTZYQMWKthVbyL+z8Jt0Fy+zEX
a0k7cLo+NB8zYJHhs8RIJgIvqk87Xuhpu5UyjZ3yJeghgwcHg4dC25YbK6F6mx3d
9wT8PL2PqpGBc83xOFV8uVMGpuHuR8EQvjK1R/MZlNRviwXHSjzibW7AVkQDiD/U
eRPj0OYEw1DfYMl1R3Z0/EBrFj2Nmii1WCIZZThrDPsusqZ4II1Y3YdkWrkkgxHB
HUBmf44UOBy5kMAwyQ+0kpfy+mk3XF9SoYZ6n83M+9yKyaUBW6z2mI+nOEBq+STs
GQdoSRqti1Hlb/XLSfedpGYeSS+kCiyRk6VkRx2fVAUfIL3xzw5dNU56q2DsXWEg
iXnpd8c7LV2kMiryuhU1DN7vrPbVYXt87fDphvGF/8g3+uD8ZLqHP7wt/uK0Rp4r
TUUURuDy9cMYOf5TZGBNz5jKx8F4cC4RUSYI1jIdDR63sZBh/oMcH7mclMkNPOsn
h4iuzA93GWslGU6MwMG/yEhHCpQcsgqCkBXfSvCFUpJ/PlKXiyxriVeyyUgOV5Bh
+Kv71o3KEvNpBHgx1YX+JNbLwKRNmd3Py90snF7li0vV3GXvmm7dzfQJdWtgIoCA
/569ljkpYhBKyxdFAryDfzHlX2wX4e+2cttL8eJ+R9GSisqO3gu6FdhOvsPC6Jex
2810XqzN5xAp6xtiKIKV6k8n212vFgKI+/G7ifZUx338N8nNsI3Y1gNF44fdXGT2
LV+XCTpDeX04iUBc01LEBg/+fOZWWrmpQVT/ofzf0cROzYxKA+caM9KJZyPnxNDS
/3/qIcbJS6rg+/7XoEGA1ISA74TRBqgrnMkCJcpgxKjc7QVyuZUOXnglB6EnAFUX
TxD6ZrryIzFDgLMHHn8XO/0Mf5n333jdscz05EnG9hkY1XJyZgJ1uMurE58ZTM2L
mqILDWorTD7U2bsVjEO0PDTKxcGFrNtK0kA6p0cAA9SgacSfmDmvFzpNJJ4u1K9L
S3O8o2qzS08rBgpPvRpDoXpm08SEkTBsTx7cjXtF1mg33wwCHJDfPuo9Dm1TfLYM
DuIRvhMzVsLxsw3qnX18PN/367+1oRVibPnuiUOdm6lm7IJWgb26dAj16QPyOilc
EJ2pulvqVq880tYn5sd2TnrSzFBXGdmywV0iGOwldDVgf1fVpYPC7L6UyvWT7rGm
4bN8QnhSo/F9Nk2eUTRm1IfDuPuIuwkuVrqWc23QeTRSEo+naEBLWmRWvYt9KXaJ
iXcITslQcXQy2JXGk0kwbQ3ay1MJ8FZXVKPKoOfB0627rifT/o1BQiIbSmabBTHi
Ng2K9GtEj/lBq2S75TPnSAldZn08kyePabx+0r3SNFmm783QOkei6meydGT1nTbw
LWJKbEgSNu5dsy3lKQiW+No35msr8FQ++c+2zNALK4rSvCBnLJIBONVWnD0vQ6xt
O1+h5tq9qnygNM3kVufnLm7AkxagiF4x9NCJmHYRkQ9nIpNcm61dQU/h3SIRmgIP
qTt5HktAX96XiKiEbnLH6R5OMBEpA7VHtKBJ+f+Uci5w36qftsGAtH4IDZFqQVRx
pFNN3uVkjPXMDMs7EX4barE0jCbCa5xui2H4Un/rorqDNNWNrA38CG2rjWge24h8
4L405IuUTodO8ckMCzIl6crxsiTN5UIWAbqYtG6vQAmsdb1xGYlWm6QR4ynApLc/
mE+O6oVWQhU9FX0+y3x21VuQTR2t3+zDUM0JaeodP+EZ6NeDTyPkYyKo+eImWzMz
rhrFwBPcbd2Rh51NOqaS6z3gWjiFk7Et+mR/sFkzfAoecXuoHIY9V+fWsfnqMAU4
TMbO1LuYy81rS/i+cVGd7FblzuH9AHwuWIH8o+tbvk4MqexLetZ4JXz45ybFcCbC
JY9liH2k43QEimWo5JSjlfK6NQrzE3Eovw86vxrYnXiDx52uNWUa3yRXuQ+Bg9LD
UkewRu8F1MebAsljadB57ZYEIEP8rotWhWt22GzS5YvJEyHtJGu4vb2H6nklfbTM
LIwoFDvUuZebiesEhC9gB/pLe9a4OnqCDYr6yUb7J1gnBodXZT1F9fZGpGnXBOoD
a3OOzyF+JPXd+RyEfB7LP8NjuPyNwkkUhwdmYEcVO7PS1v1Ig45PLcF+/PiUTY4F
ROVa2NCF9/iUv0y6ShIuOs5U5MgLVgx3CJ6x9iNFLK6piWwE7brbyUYT6hwigJfT
XGBeRcFNtqkonHkgj6NSG7i9erUVvj9bsNln7BDagUEJQdrJ3k7JEH4yDjsMFFA0
/dI7vi+aMG8V8Q8USmpaq371DfgUDd/+w94XBKk5znoE3fE47zDHrIsYk8yV6R5J
om2g7ZYvMW5KnGsn2nkXoOKuylTNxJsxpRPNMyNqnq2yCG/cJxxWQfG1DcEXks/f
u37nax0ylPZqpZkxBKbumhgQHmiL1nRAyBTm8tlEtSzDsEIO9MHwPYGBeluOtI3y
tYTg66c41jnGQidw194CQw/vyWeNfmPw64T/ULKKLLdO6RUkWWV3Xx0M5Pg/qbyB
f+7MMFSCsOlFEgkukUVA9ogPqBU+B4qldFo/mz7fI++OE5lUIRU19MJk78lLcSKw
X8/7I34pXgSRfCYxfqAJA6Eb9/Zxs/O6KSb9pP+K0jRKdD9h0jErEqqIJ9n9MyH1
uV56DTP1b9Z8FqDdgWc5VRkV3QVOFW+Srs8piihG8l92gy/t81IvHbQanmPN45Fe
D5bLdOHi5qyT1Ii22DX+EkVBnQ1hhPOxWo6Fpj+B5hgm5Xa5fZNwsfx/DsjJ9P7W
zW3JRc/EGQeAQQJg7l53WhoVK9fCd3DNXNBrmkJGNb8O15vzRJlFfZaF3oALER09
H7aYsnl7oLh7QHPAgASeAqRUeNQSUS2wbrxYtsbg7PHtYSFEJVRPeOmMjYAq/6xM
q+wWqGJdzA9/wlNb/kRGIoryJqnpKJmzGdLshWwLTeoPusgmY5/ABOjolVOuiHS8
BQctbIcQx1Bl5mC+MBNY4hqrpMYGw7VQUy5pxxp93xZWBXKpioUI684W2lsqwq2p
1tT3vX05jcfXGV00RPa9GKn74ypIGm301CmlB2iEYVjaVAhBt5d/QcUwKI6I84ru
a745IRIjQfwukW6AozoVPrSP71erS3TQmWWuvOgoSHYoiYCIv9rvh6+uKVc7XXW1
VweL1vRLpM4bAtuPOl/k75xWdGi4u88PgtS6Nx2w61tvo6jOY0jjHYHLOh/5cwgy
WiMFpnsWYlRwxlH0+PuOTOT89wbCjj78izZHvjlWfC0qY3gR6G4Mua8Wut75j7ba
JV27I/cBAUgol/sMY73nSUO//utpvYK/xR4kfYcV+zv4SmBjLk6uE6BUfq+/4fKE
F6S1VWdrHRTX8UfhR1QqwM8jPeEneUiyVszaSfpiwLH4qRwiVVCH3UmN0z3zmnLW
hQCRYF9UF9VVqhp/7xh901ezqzvon6v9BS/MVV/CNEEeHh8L+EEBL+fDkjG7jc8o
JE2GXpYywNW240kWugjXTe70PJ+z4WLisjWBeS3lrPsPDiyCs0tVD9TEBFLEnhN5
hL1sFzxRWMLQms4RkrtZUMvyUUDawL1sPPtkUMyTLJ1TGCiXM/9h83MSUXAddEUx
FmnEplL7MwagTEI7NXfTpDgJV74yVHGXdujKNW3k/nIOZBqY7ldSjjEATKjE67m+
ptsB3roCtebeeIdItF7/pmkN2bHuvDh6i/8lh94LBHsxEa8Ak5okAzmz+lObAZBh
sX3Cjvzn2dsCsF9cDgxMRQghy7EIvytyewrZYB8kVnwhAY5wIot22JovIWqerzA2
HZGTeESgFr6pGndQc6XD3UHHdVTkHao8zCjhCfCS/rT96sJqN4110bEciIGJYsmC
ObGUu8i+xv+lytA3DqW5Im3SXFobSWfn/l1+SFL3vQ+S4N9dfxwPheaiODvCwiXE
p4/Ts1tbBsJPuskUfE6LDSiL3W+Wn0HRQw6WVJjrzW/kx0QsWem/HfR+xRGIg61G
PF+ScaPxgZQn6B4s9i6jEPhniyIGEUaO3NWk/oK8YeIVbBYJFS4JtLy/WnN12EyP
iGwHMKl8/FmB+x/twqtWbZKs5YwPyV6f9G9AGDjxibyo4BmjdFScLZp7Q8QHh2ew
Af1smVrGSFmzPUrJkHLImoeivbXgtz92vIl2/876z7XglyiWgii1VichBDuKboqt
LnjOSA/yGTbS4j0TOIy66FwOenwnYaJqtsYxJmI2nl216jOH0/ycjrs4N5+/y5pm
yq0h0cJsdctPeE7cMiUUY7RUxWNOC58XKAw6leNPJEZma9eOxesg1VjNZeyvYGRs
aKdk/M1hv5JUpHwsXeO4ue+Gux3jE8zKrKbN8w4fe5FX7SEaL550uZZgwdMirpoQ
R5cZwosJbrpGYXxcGhcGBldAJSK60wytUnv76kXmnKv1Lwyrfkf+GUtP9qvEMJ+R
2XBdrJks3vLkc2M//vC5FiqadZy5b+Mk0RBvtxYTQARO1zyNM+cZ/GccPw03sM4b
z83aK3b2ABIAUAUvZ9ML9BQzj1nrKWVF5cbglFTETFZJqbwYvOGuU4hKJo9LDT3e
dLL5zdKm+T6CoQSFPrcfUcVr0ZpChRMvq9Ur7NxWe4IDSUCFp+QCfe8RrK0qiFRQ
86yf630i498vRboEttv6zzGagXx4BPUr3kw1ev9aP1cmUMghfwA2QzLwECP+m8+n
KlBRiwJ6AnPbSv8FoMyxrtr5dKq1ZnA4c1JZxoqzDoEQXeLnCkVyl7x9FU3BO8rV
mV1ofgSRZ6ZLN20bXfsG/2PlJiJqcWpWKMoOwFAHztpRDTrKIZUm3j3vbP/JfxkI
Mdr/Xg/2xqPS9yFJprhAsI/HN4MUGFHMrL6eVOSwteZ+ZJYBZYLVBpX94SST9PHS
tZREbwnXdVL3oZKBEMu84QzaUFsLcQPJmC+LZ7TY2WxMymuGVhX28BqPJWnptOnD
gu0CU2i2IMGl+4iW1ZPFH/CZ22eQ3axKAFeKE3fMXwU0v08h9CG2UFOR83qA9bbw
kJ5EQQRAnSb/rrChox0EURHxKRgdPq1bINU//K3veCCjDiiBjkaucgt4Xfe6Gd94
8ApAgBGD1hIzcC2SPfaNAlRBwJpRKT2b7+z3xF9DkneFZawiAjeBfA5Sxhb0+xz8
U6JqD3iNEM/g8LXnu6+3enosVNREAalv0Nggtj4zUBUIrZI6uo/MNzvVBkrLlBcK
2neM++5kSRdc3upFAGClRvVrgAu6znkF0WL0XBX7cWEc1PSkuKyM0tTdO448oG+L
agwvfhxhHPbtPcb78IijryTUW4SyVWrr8Lg9Rk375LSjXWZZUh0Z13xlTPag8sp0
6JuMDIazKEfssSHrwkTWhgePnHB89OIT1kN2okdoQ+cX7MY8dCEPjF3NXjmmBXUB
3y/nEuIkb2TkvZ+2kKv+Zr5I2yO+Ei+PeclxxHC4cjKYFwMJ7HXttXwpHgle5m8V
p585pczrz9JgubizXVEU8v8WoAdkzBIuyKHVkuaNYVGuoXEDiMwRlLNqtrX1cdjZ
Cnc9Vs9cfMOFQt15j2qhcYGaeV4wmbuMPwFuiztLfBK6u4IcoHI4IspZs6C5RNgm
18ptspvej3DbfkLuwOzhcWpYkQTCuYQe7npE33EL6Y8=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ldG7PcREl8BZIEUr9DxQQA/g1w21Hoh3T8dK2xt9W62zuO10NiV5LqT/CTyizVs8
bPddK1/uh4MgA8qlDZKVDS+MQlFa4vUn0ZC3x99m3jG+DSedHeRrZT5mCeGXhUGH
sqJb6F00Cm1eYjMVfxGscy7vjIVvdwx6ASCaG2TpS4ORC/TlyFNCTGj+uNaWW9P/
yFV1haLYhqr+uZz1w9IMS04u1tOCqveYyZ7LxcoCgnUT+2ffXcP4Aatt7XkQ58hJ
XGzvBg7iZe6x0d6n5LhoBIxZcf/laH37e5mrFqYcIl3Iw5sO5L/nSlNcgGZoNqGk
FNugAfWxX0EjFc6ESNAF3w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3440 )
`pragma protect data_block
JRzTbdkl3CTQgIBsJO8gxWl1XV0fJ4xD36dbQ9nRKLaTpXcf6o1iiYy6B09XBX/U
7cQq6zabTQ5f1nM6wYYpWa378wHZaIQzdR75ExBBGrhp91PudEAGHZwTVPIRlocC
JzOoI7cvsQ8jTvwr+wQrxh8D9YAk9kRzJaU8JW0J/eWIsqVUtxKwXX1+DQf6tmse
qVum2zZgkJyKJkTilUxOl1EKcuJZk9ehxHHv8dtu685DTfWGoZ83sQUGhUloMB9q
LNR72LAN2UIe8A565lk+c/gkWz9cwI3bI1NaIgqQ+AjPRZ3i4BHnGcDDesP1e6Nx
DY97+PoDuJMFlTySlyTp5eMVJhi+/67mMjUwwDaOB+OJOH9BJVKh1V2k6+0O2oLF
bQ5bFS/xs4yKo0Jq8sfIm3V2rQ2Q5X/WUVrcN+UsLFGBw1WUjjoP1CsoyhRwISiN
85+9yCZk6i5krteJUdKC3ont95mq+Ju30oKxj3FNXn/wH/jgqoqSMcn3tawexWYP
lSBzuTgFj4SmzL3O+riYJnMB5PnNMp4kOPks7qmE7YOY+OWi/c2fTs4nJbncKjmv
0wVyFKIlARb5WAUL9TpIL5yVjG5bF4oShRouHBx7BjZe8wO5LEhgalji1VvmoVue
3Cf5pw++ejtYQYMSavfJT9/eTxcfh7CkIuMjgdqt9OzbMPJjYPxuNNnhEyw8XJPR
XLfECRtPIVVJ3NTblUYlnyAbBm2XTO1n2IbYL7MQQ/6iV9qISe0jIQee2eEUtAsW
wIJl0QIenfx0TBgHviHpxoTBezpC5lWLDSNI54r9uW2jiqOHdwD0yPm4QES0rSXb
pFTt6R22r/TDIsMquDlAtgJ4EMPxu9Bmwz7AgvF0ucAdeCaVxTesMg6yconQaQU7
ZiLpLPa99KMF/pZDgidOMgkrFAW+wjrAZPc/eq53bUN4XGE77vsPU+PiNgTGl05V
/gBCI0FlI476s07op8USR9G9bnDsBDir9xpE3YtDGEKjGRu7TEBcPTDuXltiB5+J
O9i5B1SBZEXAKHDkQd+y6OKKT+Z24xY++PF3TOM56wX4mkhDePoZFtAQlruTBWYH
x+6+tThDIe9ELUNSjtRrS+Aw80FcNHSeLTFkkvmzNjM3NCjw/AjJaTVZ9FYR1t/d
+SdJPIn/vBAdJ4MUn0KGrxDp+C7U4FW9QcAe27q1gJTxCVgdc7TVHH6319MAFps4
xgMjwye06o1HMkAWmV7scEn1RTw3AE1GX//AbJOHdPgBlFDz6h1hIjDpNgAUs11u
L1DmSpIkkAycu6fo+jTjTio1W/vH3cQ9F+oXYlICU8BYZDs73vpIXBuUupU83JuE
ztcxj32trPsRlirfoHJwTqDxgombqu+KVs+RnP6AX3SrFNYzVuklyxzwHIXMsPj5
jNm+ByjAyAqvhI28iaT2yphxLLzbkKb4P2B8WMdKc4qYjjFlI4cuVS26KXanx2V6
/JNuwJ+of703Nmw6kAFS0dlOLhhTvYJ+CzOfZdoqOE8NpTudflQ5M+ZPJWUgrInd
dWLidCUO5/1mJdIt2KwNUhIrgCkMJM5YU8Gva4+Xek5AwPB/xpV9/ROQXE1pL1Rv
pI5nF6RZFgwWINXreFDOuMf/5XP/f3JZBN3uGLi/V+IzK9a+SxCZ82wHujtuTbdJ
/i5y69y/Rcj7nfijholDPtND0GOPno2UXEc4kkDhqp8NJqRU/1B6fTlBunmND4js
/zuciRt2l5jmdRP/VDy1TXqZJTANTkq9JTpcV50pDxqMI5qv8DOO9V+ncNDLRvXb
Ey2Gs8fqBMGJ/co4x/3NDjzY+J3il+POCA9//LUcAvu2eCuu0KNIMbJxDq6yM71M
EUeUq71Tbt2FpNRmoJYnOKYbXyxhHRoDAvNvD8yX7EovOh3sDy7fWCcGP1NUsvqF
wO8QLc2wsGkcTkVmXylbJHVC1S31EDkaujCOLiDsLiSka/4lz2qIrT4l22YvOblk
oinLZiq45fLOnq+h6FCrQbhaLHiuhGmBnEbpR+YictcWrc8OrbVN/oSo/3pROXFo
ICI3usoE6AJ74seSmPqHunimjuCMsRUj4axprx2do3eXvAtiDbw1D94QWZWVO40C
4i2mMPYD7f5Fmf26/xf3RNmS+pljfFtPtykD+gEu3ECkz3BnsiejnootmyQZ91yO
cT/Rt68IEqnyAMGBigZ6E9G/QBrUdp7mcb0XmzyYZXnPurjTmm2oIKDrDZGy+IZ9
CZbqaSZfjtk7nVTR8aHl/ajMnvU6SFcwDHWMYiFhz4ybgHpvVpFXz1spLdTRUYii
lyMlDEHhE90Kk4KOweT5X8GMn+uRXumLAaCKADyFuxbiT7irS05YfqbY8WzpMlOS
hNArlsvelm6+76DoaRqgBQE9yicKnRP3942WCh9oYa6ljuZ7F8l61fFBOCmaXSPL
JHtCj0NgXTQwKuHPMaIAO8fOKTShE0MS4KLcW7Zpst3kFOPoaLm6zgt+i5DsqdVh
5icmE4ku/f7oohMSk0b48lQxS+9JM2OgY7M3FfqjPU9IoOtqBebWyItlFFo21wdx
VilTOaCw6EYxn1YzIjFIno+Ay5fb3FYJb///G2KZnKMZHR0PcOTmff0o6uIU6nHg
PQv1jw2nZ3dYcFGcvo4dAQ1LdQo6jxpGsTn9e5RfztmrCWWYMWk2zXC0aGCv+5v9
oUeiXT1FTJaaO11rhM5hJVLrEPy9hnYo0eV5bIeScHQp8ddrFSHfKZFtQV0TUoHg
zHecKUKKBfv31uv0XcMuRB2CRIC9SM2ZjZobjMZ8YdJUTlZ+ee008JrEehmc2YDG
lp6noUVf5nadVm8ChuXxDs5yV4drWZRi6tKnhPvy4Elhv4QHselSleJoQhEDeCZ7
/GG1hLLWszB1aB+WgSxguY5VEqV8820wxW3ZZPMLren6E33nHARgZA8ArtPpa4UK
Fl48oIjgZt+/z9quS9AwZ/xb8sk2nQANakDV5lk73UtDmZZtqyAIRGR/FW6RW4tB
FFgbWIUAyD4+BLqv8yWrMT3JAgfV3CaAGNoEKc+wNj5y1RPh8N0q2oQ6yftlOPN7
E9gw0cdzcwcbqznUKB7Bt5lMM0iF7hIk9qDkxrF5Q/qzlmHQqML7z6XJF0Tfz5gK
GAYaHfz8Ue6F9NFRA+WZZMI3xLS8NfZHRZctfPau9J2wdVd04iZ6h3fhjv/K7Gl2
o43HNPOD7qNcesatIn7SK9o6786Educys+PP1V21XsXp975ftA/cZL0JnxoLsDyJ
OE5q8lt/24VlcT/XVfz8tF2ZdGce2GS9DOSdx5rx5YRY9LQpRUgRP0xBqwtCij1G
DcRaXqYu2OGgIZ8njLMrQL5rhuugrTKlk7fHe+DelACAadea8OMEd9j+c/bmyP0Z
pO/lz8Pkmms3ihyV62awDgNZKtPgZyAWKtnV7TOIlfvD8hCs5/Tg2VSSSdxKgPVz
KQOpEfMBFJxzYYTysl+Zl0rDEFN/t/8lSTK3EHmfb/FNFCEeT5WiNbOwsFtwz+MH
sXDXsjKq5VbzATzdNPSiBHvPG0g9WhlVpe5g9PVBYxA1QwDSNAeuCQ/M6Cnv8R4t
1Wf6EIQKGhD2veXfdVNIYJDZeRxporpL2BNalHW5Ay4xFlRqWCw69EbMNG/0F9uW
iADCOPA9+qoFeBm4PYzAfXxzqKbkvc0zKoiHJsD1kyRXzNjmDerKmRsqC1UD3+lK
ddRtD6BmBmhQuhZLghP2QnaySEUqPHSzlncSIYzW3EQjw1b3iP2f9FoPmYeGrrJo
gziPEtUm81PB2qsiHYq0y/vUyv5m8MufSAd5yW0p0Yykq1hNRvoOkrFonkuA53Jj
hHA0CvBZuZWkWC6/NMpMssRQ4kfGd3HvRkcbmwlaaq/qsLVPVshu8+ychu4rsg54
l5gg8a2xu+D91N8rla6FczYQoH0xgMoqU/PMii//w/JtcSMRWjluR/hoq+W0ssil
rKtQUV1CvSqZYbJEzFjAaEYLBipsa3BuJ4qwFKKkSC/VzJlPv6Zhp62DhCI/4xHr
LleqSqWoCUsCE4UV7MzFW5SIUuw1JU8sDTUCNZ0oW2UBCUUWJuGAdD26P6ETLu6w
5FF/XRJyVeJEgfeFNsI8GECBE/j9rmQu1BmGcN+FSmObC9KPiS8eqXYfkmcMizxZ
0DxIadNqI1pcDM4xyJ1uFaMQXVvGXk0q9zX2G/ARObCLHJ+oWb31nsjF53PLYt+m
Vs4MTRaU5hkkJ9uH3L6tyhlV/gJheeQB31F68jA/qrAFonvohEb1k7JqmOL3a6xv
sdkLE0If7JCKUToijBUnzcBX0wISXrgW0QG5VXuwEgEJd+DkKhgvChILAm0Dvs3N
SkLrbnS+D/h9FftvP3wb8Q9ZjeIQbnJ1LS0gD7q3mo7+Xg0ghYhJkiZHl5KtjkTx
l228DbiOXDT50OeCdx2NHIttii0VgPIHu6qVa/eNqYCRVAx+LVUNjZcLawG5m6Oe
Z4RgOdd91k0iK0UfmtpCy61hjYjGlvYlbz99i2GhAZBpYHLXzQjWM3WtQExALIsl
QY/OdekjibQK+RSaX9wxFOE7NgNaqR3/+TDcCWmSLr8=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BwABA/jDqBrBjT2B7WdECa/Xzyt5GX0a+miRYK/whIXXZDFhdQAo36QOauSyeuk+
LLB/k8aisJnOMOqBVCghigTBfuXygC3dDOdlqoG7X+93PReU6zTYW3D5U2pyEGzY
3x5RTMs6AgURQPExI/u/0JZTefvxvsbYBcG57oqCa8FcpJLtIce8J9+eJsIDxKkY
gKoraBtsrBzbA6LNx00/WyiIHMdDLN3kR7kRl0Cnw8G7kXrPJnfME47IGBLOlD2R
SeuPSnZw14tO0yVVTlVnXl+OJHjHgH33lfhvN2gvSAAf8CuZRaob4TlxySXuJunP
uJq+xHBo44eDEpKWhiCISA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2176 )
`pragma protect data_block
cufXpXy5l1OsxZpsa0xso/3n8H1Y844vnDqNGexoxxXpWWiHHMWqSnN4Ho4Mpd3G
/DboJZCr1QdMrYItM8W2rSF2Cdg6us63E38FNn2k/EZVGDqrgGtTQXeqN4jBAOKj
feS0bS13Xqj2Z1McRfYOr8SVeDSL48WzlZRjaAFy2XpV9559jfDfMDvt+CUaoloR
+CuBDx85VnYUlzIFCKUSStupVFjPn7+Ky/4N8tb4W/Kn/yl6H8mKuECCjkyVrc9v
PXVwwByUkZYhdnNF7gRb+pPKlUhOoRp8kQEeN3K6PinNquWXnM4hKzpDdJiZmM9j
zAyymhBFO3Xed3+NZsBO5A7+f2IilVYWcGnzEfe2+0FyT7xUq7C/bWi76cb2pzmr
dNwE+Id0lta30JEpUQQVrvZxFeRBA4rxCSZeVYgG1D2LVIMJq313pOpVWAjECgQc
Vr9gl9XFEPJirT/ki+PxnRLq5naDJZRmjEniFzztMls7ArUV1ootDOVZXZ8FhpW0
dhqrGKvKvfIA4+eGViuzCph2mDf+S2XECYIK3DIediXehyDLOQbQpdaCoeyAvwzm
70yN/QQ5Zxd0b7BbaBwD0Ig0+ZVi3X5BzbR6tnohUCosM2My9DhSKRkL7hyfreOa
sE5DHyToMrd9uSJafUYTDFhgtt5F+a8PhdH9oBQ/yPqNzejGmbYRd3tBfyvs0gnS
2P0lkV8Oc6cZZfKDgn5R0c/9Hd35w4tXDCUE7n5njdx+WOAjAy/1pp8/oxzIt0Tm
nT44+AMau67uFJajYT/zVkGKqIchybfdoN2glbnqdm+yiu3u+iuAdTcJ6qnaU1n9
zEfYiJMcJd0OE8lWtdc0n5PfQAvsLw2bEzCTfkonKDY6Dr+NA+CR315K0kMoblmY
yeEamJAW19E7a8Y3qBmNL+qDi0VoqHoNjSOL71DuEscUffnrQvqwgSltc4PAniwI
/BV1bHZ0ZlMhwCdLzoAdN9ZuOWCxPrNsexaucGe93kUear1C4/1UgBrKRkTXXEeN
SHH7JxOal5tZzE8XCyu4rU+hQ0rVlP1k3s3QHiGzcE+fdES5jY4CYr3CcXYslIYj
aMoQbgsofdJLBOmfDeizyLcilQ4gZCDNmEJNo5QJpK/th8+9iSvB4I5VHuYuFU7M
tqnGsmmUapr1rKO8EQGq6I59sTRoPsw0ppsSvsDUn9atV7M4CCCjlBml7L+aq5ri
mCL2NyIKK8Suo4ViARWt4m+EcjsmULT8NA5KXBcT/cIlYs2HqqE0KeQcrBzUsO2c
so32yjV3S3oMcvPceo9WOEyAQXStJFU5sy7/JyylTfeb58UQM1lFryCBhqHzVlgT
Hlr+gGrpftsVL/hL+WZtEgqXu3+N5sKckw0vkSxy1F5680d4f1Wu83hC3AiNdDUo
xVxBpCwlYBL71diohtm5AcZQ9piEHRLlkZ5VbIF58ybieaTWD2wJZutLdHV/mjXF
tvoiFOW1iXAPJvI6fg154QcY884MHf4QTLUAbDDXt6aKCuxIyzW5JqpjZq1yVR3Q
hrXZJVeXd1BDAVor5Mn84cxy4KAnnxpqfOKSR7iJcwaSSxG1fkLioQgAbqkacnN7
O0haGmvXSmz3n8jYrJjY9dazCZQwlvGU3UsYVwZKhczTjt799gYo7ug/xwHODHzi
ziJaoVW01MshxMWL3exY6AYrMOTGUGZH5ABQVrIYkAE6IMlrGB3MBbns5d3bW9Pu
/mMQCErJdPYWq4yUZwkWBvn6H78awRjKGS5DsMu1jG47zfYyltMg4sLfaoXqOoeg
aTskGTejtSSAVpPtiOp0uzgY+cBETqJR7jFhRcJK2Zgbx1BAi1SCjonS3x55WOjo
M6e1P1FniUpQAXUs1v/PUjg8HaXzIDo8KNbWSxOiQQ5/6CzueE6RkwRUOt+fHlV8
baw7OSfVgYDezhSe9+Oa61YXGOdBBseoop4K9aOnhkfL2WCYxzi1Ja+ZhDvMZJQl
Kul/oDXkGcvI6+6lTwFyTfLUGwA/PfqKzvD5OF2+xwcsHGzu9GnOcuKUz0qDSBYZ
eyiKU+tHcis4+Q4PrpWCWAON5Qrsj6FRl213X98V4WvOjYX/0jcLx5FHqgVREGNY
Hj3nY/v2t/c68lLOrZUhG6r7nRn4VRR3n/Q9Zt0+vd7X9yb5ulcolHG2GJgGNZj1
4VttULpdzW5PcH0iTXYO6ArVVhamk9lYmh2sw6lgBSTRI0HrYKgkmSdR3zIt8nIt
8KeX6H29hbEU8liHgSXybFIxd0IMCuIVT1z7P44uxxBZLldQVMGaa5+N+PdQ2XPR
Rp3pBZ8Xvn8J/AIgyK8LJ/zZd64nN678TOav7QOwAKdNwyLz1Q8q0UFij2BI3mEL
mxW02bPM8LsOwmbHA1iel8/gvbzk2J2lqrJX59OoF7Npb2fyRHBKxLDIsRMUCjHy
sdNKGeM01mAor5PLJKdLNdDRSqdXRfZisWo0GohVbrD47+9ZuLi4hQxmVnCgWhKu
+zUJY4WcCXZhLnXzQu9F1WT1UbrC9BB5j7Kv6G3PRHy8r3/bGdNk2XEN7Giu5H4p
woB+8iD+CHm4GttEfA+Rs3Z9KHcYlAm4F765WCxoe0MAH7SUIrSHwCIHR9KDJhyl
kXFXzCaExqejGUT36n8zxR3uGRxDrckXKONZaNL2D2zHhbiYMIxUHu7KWAh4Czub
5ln4xTggIrFzxzgivs0QKL9vpnZzP3znnEommGctbY4SBRSw9lN/wDBDHcxDl514
YWik7a4NrXyPs7yuRIhQ6ai4NYUTe1LAEjtc/GhBiBAWVBva4If6pOG/b4wygsct
rx25E38Jg4rEGK5ORKLOMMgqF1hh5TWl1aTFx83+oxcG5bAOG9GCi0ZSIYhgaYo0
09I8HArx4bHL8lwkJA/NkQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
F8YptNaGhyrgSnS3vd0tqsr/0/dwWU4AyQ0Zx7UYQukeCxflHtNiw0GwE+WReT6Y
vjwHM/3Lapx9Q1ZJC6dVKEF6B5gNxh/a4DglZ/IVAII3yFx1zhT7LmCzO080e/cW
JxmbO2tmhgBMRFM0bvcSLBUS5qp8NpjrxnoVImJ4MDvv7VC9ZCBVshILFoAO5rUr
7cWrnpHs8fb4spjZSo/OofzdFDvWNiN1kFAtT8eGosnnzmA+s+wphsKkmDgbsX5E
plLyV2Q+VPlXzBR6DWSYAvyylX2c49HloSD5GAOtzZZANbi8pdBxy4c6bAm5t2ec
HJ+n649jq6cK32SE9fiWvg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7072 )
`pragma protect data_block
YzFv2/ArsJK4912ASPFnL5eWElvQcuuonsWZ9KftFTUGuOH11hHrdLWVswkdQQBZ
/kmsewWPvdX6EHmKE2BvXHBE91M0rdpTnh4A+iDpVvv3GR+fZPbyz+e6YSiaPQNR
lzSNYdUV0eqXG72C0FdJF+i0c/1umCnDbh3L0IdvitpOGp9/PsrjsSiEyCI7ovUS
8Viy2eQ62Prb7bcqAuh5kUR2AP5yfJ+WUC20ImJdZzPRbgZN05V7Zl1RqGs4ZLkH
DEKNZdguTvbvrFnazodPOwQuA703QbHNqCOi0EECJhYImDWhsLjBXILmbqJMFahF
h5Ap4IRJRIM7DfzD4wDHgpBnGAx7GT3RHSBFHIta7URtTHEI9V8K7Kdwe5TcqPyd
fQXpsAsnSQXTxMBxeuwQKOa6KCDJU45eILg49Cwd/DkW2NN8PJzJLyDm/CNau5gX
kVwrSjNudtWyYgHdjjEQpmGTifC7vugqknSlZMr88J0kSSVwEhkUFfjP4xKE9voF
tzFqTCK8wDHoHmXfWEcUi33QxG/yZ793ZF+D2Ja37nLEu3AU+Wp/6bLUCTp0kiwX
axe2kAxSsEqwNUPMcf7RFq8J8pnD+I3ukTdfOjGMoeM5eQLoJ+fgC6elzh+ifkdk
KkBm7dfwwm2mnGBCkVxAPmqPCcT2NcCZKx6wTtKCzMQHNOjGR7Xa+kvfmP2nSRfk
FQkGVlpfK8uIeUvPVu8YoUPeGgDwk+Bwc8hH25dnm3mHC1E79FaXNaEC2ECyXZmt
a79dE88LK38cUelarbEfhKNeFyXz9pBG5t/Il6T+Nry70Jl7gSWLzdgJYab8LO2/
DJGndAwdw/XmeCtu4tnR2Wdn+gRUhlZ2Uc+S66pAP0qNB7TJjkK3xM7ESlAeGbHZ
5u021PqNMjwYd7wqoVB8dJENA7tej2Km8z2MNgnU0UzG9p/VuenRRHkKJVk0kHvf
BxJO/wdZm+ryb0M5M2B9xRKFiVdtu+cEYpR0p5hJd1f3ixvrvRCyvym3ocSirQVN
9kw1i3G+22GcHlD6nerZwIIbH+u/qyy4l31gVHehTb3GZz/jP1yxvHnC4mhO8i9F
hCNeJ1OQI/sGtvwqdekOF0jDZJxhmz2gM/tHrq6ldL66tyhBLsicbYJyDTq9w5mV
4wKTuNtihvGI0NmmZ9ZJ+hAYdQmFCHtwCgEKZjrPWzli3VMDsIL+F8T08w4TsFGa
jl6NVzw1FYH1D0gZF+7UjtjlrEymiGTYO7nNbcHBSlgVeoU6DJI7lMXCz4bqs2q3
7m+rigoT5FSaiLvwV5f1vu7bWNxb2FCJ+lRydp7HbSbpt0pPmjz0CX0cK9bx4BGn
r2LDRY0pL9/gV4u9KRf4/TeIJ8J0cUYiifuinz0bcKrMha96IsqKqiYSi0r+tVXA
9X7bJZgnm+3w6ZsPxqS8lHhKaQRxsczdzpcFzR0kmn8Itck+64DS18Vc15zXOB+u
jNH9jwUP88jr1QcQJkkyF4UrO503le+dTLLbYkpwLscVI6Xb+expk2edlv6R0WFi
xa78JGNz+uLjSTaWU9ygceNW30uWxhpJMK6cCNPdxZAuAC3hDWbvkBtwEzhdW/sO
K495W0jrF05afFduagXRD9x43B7/ORO3UbXk1nkRDIeSguMzL6uo0lkimJtJmduP
8/z9flqi98zR9MyT0RHUg8EmRtHJ/rbmJQJ06VFSfToCnCapFaFZjqM8iFfn8TSq
kvQM68IkeqikJ3/q4kPBhJM7imaVY7F2kB1MCYUj12H+2YIzaR6AB7+7/HyW4P60
vGp2VlDWGnkgO6DJ3wwn3HeHXRq8VRqslHgYNE5hoLO9cOlQbUWg++a51Ksdhw6D
29qynMPxE/JB77DjqBCCHfrzFE3vNpGU01t+qPmMb7cUQ6dVrV4NNyuko8vjxp9F
3LAdX4SrnvYqs+l8mKvZ18fIXKCfdi9YSYrd/K7NGq3YhuQ8gJphPkcnY2tVRoR0
b0c90L8+7Y6l/wWyPEQTzJ3IO6uGnRvEc4upkz4wlWZ7C2bhsfZJbzjzWv18G41H
yn4UOV4vWZW7e67C6Vswh4YuPewuIbioTr1/Eok6DwyolmqVW1jVMStYKWtPCZsG
Qs8wSi8Yi7vH1KtABaftjlDSyqQnoohbA7jo9ESNFQBs8JlfF0J8Mp5D6gDBPlsB
xmWg6EcMIVEziVDD9D8GzFOkOnVmxoAIXMrMoKtRY6dI7aG7cStECHbCrHgqxc22
VBhnr1nE47hcR3LnSJ0sXs6G3itHlNIL076C2pO9uj04PpgdEgqGlpmtHosCCB9a
3CqNBoz2EmYlyOdfMVuqQJDQal4Okz0DTRMJfC9oB+UiIDI90MyWgj8yydaFDBBQ
kqi4fxj5SuY9r4CuxjlKMi4l8+3TshlJsB/m5TNptt+dQwUqsY7Phg8QEWunsZjk
ygVlodN7XrD+7lrfF4o/hzei/rORjl3xSfNGQ/qAFgCntGtmERkSrLnmoKK1/wDS
VtMBXoH/smodhDYmH2Ewj8nE/9qv8NPF16JO04ORYMy/UhOOQqjl4eMysiR9TR2E
3//TYhOugLLJps9Fx4oIlihHxglgNXZiqEK1Q0H2OjA1bSmJMK+XF9iWmhunCxVc
ri/kslnSOMAgPwynwF9uLVhXdet+CuuuWcGG2/lt52729d6VEPHnMLZyZkwA/bj3
wsPXkrc3Xv/WPfl0KzGBwHgG0v9KZcb4pXSEKTm3sL0LhQLMGkmLqNWhQz0TSJGg
4I/MOaEjl0pMRKVu2AmW7IKNVf4Gzty8I/lAEcCaqwtv2bdeUALbLYA5+g96r8d4
Oi5HbWQNO6pMEwHxCZPlcElUQhv39pXLcU6qrwMOFAsuAur3s/2erjithNuGAGX6
e/580nORoiG1iqCXEP8uqseEc1x6a8adt9+Sp+8mkVatz6nvVNTLglNjD1ULMldD
7C+ROI0WJ64Um9eTfcFWsSVyeLQr2P2O8Pr5NqKaJdTWbyOJZni/Afa8ZuP1vNU0
ZfglE+xJnuZH9omKOjSG5jgLWKx+r5FTWDIMCItXRunzjce2M/aX928M3bdRdFHo
/UuWoLHqBoE6ErBNSpgo6ScEJ+aQSFlqBkEE+WOZnOlzY9EnNlCuYOal2y+nNsK1
sy7YrvIIow83N6n27yOu8GDKry0MRNlIjyAfR2w2uifUf71dFolVTgpSnXzu9xMI
kxn7RDpbzsbO3woaFzgV4rV5LaoEs49vRoTXP/os2PGweX1UjzNvU9anWLgOqvEP
vI/XtbWyPWYWXBgqqTIL2B4bRn08sIu6xxPr8iiPBcLGpuPZ61r6XhP6Y2RCPwgJ
NCPfitXa0zncxNu20lnXpt5aAGTG2aUjq5lWLniODdp0KnnMaOTHrAxoAv/1tQdP
CQhbiKaUL5uQzo/X/Sf/3olrjSpTbuM7sOUP8pQ9m4TXmr+L8ejXyLSRcH4u4J13
l+cwOEvCEn+cieulo9ti9/mEjURBogaQfqfNMwogjkJYSbO8/HtXK/KwrYRsJ34K
va4OhmK6noxgbJ/jUqvmDxFcgrh9A05uLrSO2rwtMByHIiRz1b+En82l0X3b94yF
wDu1iprWgiRHXX5c6htSs+TfNq18TVAKnb0YndksWFnnvnSOWmVQ1o/62qPqfPrS
gHJs12jN+LvW9OY0FJ9V3t6j9WrzSWRWhC8/PlC7ZhOTImIPKVY7j/Xfxp7m6giV
6NQFpviYVtrzIAPa+bMjK5MYFyBNNwQVBGyrBhaLBl1pCvWxQyx8gy/YprrwFDTV
401JiMqV8Z1KverX++f/2Hc3T90SwfFqEXJfWGHYK14TXO6AUgKcBJapg/9k9rgm
Srd2LylW31PHBstqX+F6urLYp9U9ko7S8WXSGnoEa/Zx6sFl53W59mrCSV5sZpsO
c1csyCE2tV/MBKVlAixiCO9eaJw9psbu9Dmdzcj1OrB1vQAZgZPyZ0T2w98G4dnX
g7MzQjh3wvD0qSwdcaAv39Xwh8w4L9Fa2o4i9P8dOKlc5O3mbvzpOlk3qU19C32A
4wbO5B2A6WOu7uyTEzrV68WnqON5B7uX/FliHRiOCKWwxy12eFagTApUGiACoEdR
LA5IR5DytrefzjmUcDU9MULyKs7smb437VpaqeIq5JBQnVAgO6vOfWuCd0Ayu6ZB
mFzwfygGRkX9a8CatpPdbCwXFrBnXTqL/553O7GRYCkfHE/9GUjcgSTff4HKXmwE
/CppU/CzrCeQJpQo2mmT/5tdbGOO5txJfmhAKbCc4nVsaTk8nC8zT4v3dkoHfDB2
fBCaTAUb0HX4fBEcouP2Tg7DG0LgcDNvrm0F5aS7BaHC7rBycz68+bduXwrqn7uR
Wn0YZfHqrCAOEqgkjg3fgXjIezxdekRf6S4h5LPQ3E3nnW0xEZXj3w+TlFcj1y2x
lcHg0J549I/Mw6zTVcP7M5sf6rweEInqG+z3aFQcvk1X+dKTiCiNvvrTSQR81lWx
ArnLsKGERJozE5z+XZZwh7oCvzMwxXsf2onUWizLWrq9qzq0jWdIYr/iDL8iE0Tv
G4WGNtkZxqZzQZmUh1nVqwh1tbx9Sosg0pLNxEkqrEgdAe1JrefU3LmpZvcGtjVm
fljyaPBuVcTjIjKcFYPFIMCJR69fGvpsout9mjfy21KbPTPrMauG8Dg5cz98Qib2
LmR7PnYPB5LWB3p0wJHVRgx+WQCy02i+5Iajb5iUG81jB5iPARKDRBe/lCoWiAYI
/Cc3ymYrgNaYXfI28KeuxiAOTrJ2Ok1QkEt+6mr8s/eDs/NldqqYe0G/zKluSMX2
srM996pZgupi0PeC06Ue7qGZI7Zt82zi0zH/sB0TcpqdwJ2YHVTgOKH8Ckh2goVg
e1OoPOfLDemrLu77U3YKSMN3ZSU83QJrHW+/wC4uWTLIaW8sQydXVHcJoECAXB18
bll1NAaor/oZgHpOlAsoqkndqnO9rlfjDlAJtkfocrqPp18P7aSNBVhwKbv/rojc
paTkgef84oa8/aK/smP1EV3a+4+QiKcUeFFJ4i1b4/Q62Wx7H1HXxfh1VNH4F4aQ
ActNv6Fm/Vqn0dzqsqNUC129uBkn9Z2i9WwtviWHY+GukuQKV49yGk3KMSaPRqMP
XAN7nS098DwkcZ75JLFh4hCVifTwcoZKFg5zqkaLz7wln+6naqMs0F3B5cHHj9TV
pGSDN1QjXvxlXiP+JLIx7R/4h0Bj8geWOqss0Ya8Oyg4tZLR6hiQfH1yDbgmZZUc
AvDLuPF/uu+KOwKaPUnmmlTJswVYDBekZxn0s8JXnKPAwnDiBzHBVRU0QZkw3t84
gZQU0Z2kWF8UT5SB3kLJf1AuONkPOQuq99DfcTkU/8yKwRFGcEr2kYgoBNrx5I+z
C6tphawx/jOyQZTd+bomcLIzhS0e9jALLhPsXtfmmIGUtG3aW9f2vQAT1sgnHT7M
EQsvu6ewnjMNnJ+k7jcFiDgL/v/upmTEATb1/akuvdNkLXWVnNyTk5IVC4Qk1nIx
dM3tXGt/bZPzwKyn3u1LCLNwopIGwEDhli/AyRahLjEsx96Mib7xx4zXsptN+qfM
kFBaTNHZKXZf94zNnM/wXCpLGjweweVMZK/CpB43LDniwoVQss/iFxpeTRZScRvG
nbvd32yRpVUettxCH8TAxU4PMIPZizokybSo7jI1ZPWIbZo6NanDWGdwlDtjhKyE
E63bjLqLmDegFRYU81AAhMiAUrqgIjw5tC5r50S8Tv4ticJfQxet+f3PWJpgq8vK
dw4CYFoPSZ/dtgDMNa37H9UsAmtlopYt4BZg5iu/QKfVLcVsaOKfXHRYogPlRrTs
iMGfJ8J2NhotRg6zSiJji/xnfgLLwwZx7pDtlVzfmdm5DvtOIgenH5MJqdTmlhEX
OIX9E7i5E1QziJsqwwjegu0YkwTFSFlzwHG2bjfUALwfMAuG/N3p7Kuu5gVcIvax
1zEYeycTRidArWKeB+vwGpV0+8TASQfgV6wyi5Nfr+vrSEqgoZFaxLfs7h1vgVvg
of6RIS1W1CjonnefTm0caKqOOK2RX/VVjUM9dlbQGVjnGyAaJueHlTne1Q85FnVA
M8yH2Z/xAjsKcdFnTWA/Y7dLRJ8QZF4ho1N+WhpPq6qClHv9fOJaS2BkEZokzZoh
979aGnlpTU9GRPPM1+JRueXoPwdPNev7IofwYit3poj+Tr11oxt74kjsv8hLDZRe
njM738glSaVwd7yo4V/8jbZ64i3wI5YGyWO2rUl+8JygQIY3eScZFY4LrghiGN70
PoW5Kt8WyBjS102B88kYA9HWxvCETY2SC16RpLNsVfbtbni1O7OEs6oV7AX+Or7I
KHdfic8Ne5bR+ee5B86lPUy95worE/jTo1siHm5lz+aKxdsi+IQEUOHS2AqKTffK
DhsOK8ZYy4e8iyoUdKjQQ7n1R8X9Nx0Os7Ad84CwfKll3RAJ5AnhUnf5wetdG+35
6TpZbNkbIjzP1SGjguykQWU1VzZYWN0meMO/wBlHQPZZDhHaygk6fBv8C/HlXkc5
LTBrPBywFBK5MX5gqMW6zsIWHe+WEuD7VwQY3nnuBl9iJgUJatXHmfaqeqagsXuJ
C3IFlUL6Fkrwfe5CPqHp1VUOWtDN/o9w2ZvRqst0l0SbJpBhg7q8JoQvqFvjuJ9q
hmQ1TheeGN+a94W7D4K5V+muHbQAXSYf/wU5ki1rcjlPbUy0R28iStZ3boXlx9Zm
Bt6AL5eLQZhlCWQI5SCi1aXDIK/85vgbkqiiesOv+1projYH5xNFJv/iX4QytvBC
TMfZGkosPs1wNraOGSqxnvrLigSNGDQlDVuiLJcBRtGZunjMZrp6n7/l/5kkeoXu
bYmTDRH7fX3orGRR8T6ZL7pSlDq1jLSAhUYIxKCF2mY9sTR8LExfp49xL5gpPWGp
hDWTOtV2iXrpkz7XCKcrP2qBt9oCgCxJDUN2m3HsU/aozblPiVyCxj19xC1cKb1n
Xd7JPt9BKjfXnV68FWqrlpw0xLZ/vfwhuTXTPZBAPuOL4eSwJKHCCVVAYU36egzQ
8lSCO7/Dnw3op9kvwQDeWIesF/OPAKUVqHn4V7FotqUAVU9Ovr1MCJ2Afks4U5Wb
JVFl+wvbzfHRFK+ki+OsFofA/h5uNE51ljQeru0ZHQ//VlvfKy4GRIq2KHxEgDNT
NyUGIpFSZxDvfh26vy+Tfkw/5qjfKWJKLIdtTQiRMe71Z5D5dpC+llpiXQaQsCY0
ojl+LXzM2h2WcG03VadsMOVYPtGHa7J9TgGqU9ar5MmriD73dQi0pGn80H+hZbLo
SvZuE659qdvB+fy5PQUtIfG0yL6L3c/0tORd3Ixa0G0SaCUzMZweFPeHcxp2/clJ
nhibtCBgQAIDesmu4ADruIN7fMx6yycDzLxw0H90ebGm3Esu5XUHKf4TyKU69aao
8BgFiMjDMt2yDZBfSaXH1lLjs2vA+KBgkdYxKX8VnMvtxMmNslNJ55gaYddOf90N
ilzefiA8JSKRBAAceG470fpPE33a7evoc6QCr5V2rF1pmtpnOoYHvNHtIeK8csAt
mbbbDzm65ONeA+wSXVpmtCYk6Zqe/NGC3GSHCXpKDMpuluaMczwIudt57wNeIh9h
7OU918ZQSYAjzzXlIBVyWOatJMd12jz6wSq6yiVBjr9I7Q+ux/fb8wAmmAQ3tzQF
TVe9NFLrd0CBOvnjFCJAUVXQ4hItT7lbeznlfcrze69Nnl8pzs9lNNUKfC/pInB8
AZ2nB3K94nj6yNHvoWd1zOpEid7+SJiAQRGiDUxmpBmbozz5OhWhr782Y1ouMKnG
pl0UXEmgnHWfvFxvog4PndQLKLDqd2rk8PNda0nuliNFY8B1I4NKALbP07/GTwRX
qtt3dfu7OJjOE6OCmQTd0wS4lw5ZAy0qI7M10/ZoVRTaEhGxy2Zs8f2KRCoRsrWh
cdurlHBFqpgJ7wa3avYjX9k2HC8WBIaW1hY8uw01Ps8dxlbadvNF0Sugud2Babwj
qJHvy0hNG2fp5TPsoKXtY4DGIczNk2ncApRmuvEiVSxbXDKWeFMN8x6mEzBEa1Sn
FaWukWZiQkwQjoORUykuI9oake2tA2ZXT0jqUb9Xwt4LLUDdF8QR0CmET6amv9Py
u+w1hssEmRbr26xukiip4zVhqOU4ECmdYguOhgpcsTaUpL8zZIl9poB++2U/KrpR
aJ5XGCbJPMqsV94+J8WVvwF1gz95C1sOKAq/yDcP4EG+c8nSQtRIby/moSA3slgP
WLAIVNEqSmUsMS3Gdn2DyraV/ef+Gf/RDQUND8MagwVmD4xf4XMQMmCz9ikItLv0
MubHxzKVw7MgNoJ0JnjYf9HZPGd9ngmUnkNLKM1VTQi3akNSdAkS6evcHd9ft/0v
oIkzB3Ws5mCnCFYE/VAZ8N7ybd/fuiO2NUlHSsr4lPcYYervZixrkO/8D8g2yZeU
xPSL3K03cZsRS9nVIBRtSIg8jo9hFHjP4CMZGz9ZwhOJxkgMIIT7TEAHimP/N17t
8p3ZxyYeXAsbnDyZ7JXlAmPbH7nz5LfDTzlPNL7W/pkv2rsxQ0O12SvhGjBvPApK
frtuox2JojzmfyLJyvPkKWiIVoMgFAXhndDJ+va6m666v1YtG9sjKq89WyjQDyqG
UfxS7rmViDsKp41+kyGAH8n5HXhCPV6eRxEjOTVb126d1X3nCz9e2afDwX3NfRB1
UNLmtxoUobl7DHoqw8fYAz+gT7asuSLtOXaoguf4Z188WpL3tK806BJXoWsXFVQA
y9cWGuzMLwiS69pgREkVXF4bfByDYMw2sD96nA0LT+Zp8mUdR/df78TxyYxVNGvW
x7h+qiPNwQ0gl4c6lGOJnHLtxUgGQnvYaIjzB9scd5aQcXxXmjWP5eI7/G2jCFaj
NVYaRjuckebCdxiATxDUO6MvstgM5HYNaXYyX8IVA9JeImIo6bnCFn65Pnt9hmck
UXcSFuK+knB0RF8zSAImLjWO+hdNEgLq2X1/KjCUvNRQ/QfeRP9tYefCpG0cjhF1
V8qJhoGXVgaAiKibi2hrU0dyewFdaOz7TlR3uPPEzXtJyyS71o3rL5IWlqIZAApN
yzaa7DWv+iGOY6JiHkH7ikZs7WIYOktwhmLsr7FKkD/2mn+jvm3WJDQGnEWLqDL4
9+rO70wSJHDkHxGvi3x1iyAetqly3E3ryXOoH/vYnaH5a1fE1my+PKcrM4d9pPb3
h7SzIBip5AQfg8Bhpq6M7bidq24vHTBnaTNrvpRbmuQJwkFAdv5JhDFqRdGvFCrC
FqoWDs/HYWJKk5SipG/SOwQRmwEw8utIwsjBkCdTnvze31TJ0PLc4ZRkpFvFKDX+
R0b0pOoWM0Fac2NN51o1WBBqGqutVxKOMkZKURT7AtVp5BO8efyTE4ceC9Hyx+N7
mBSFpmTw80WSC8If9+Xv/w==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
CUofiODC9iRVNA5X9iJLwX5HUWOu/4E4gfn70Pt4jDmxTxVSeNDh6QtWiTi74Pk/
MbGrj+EI5PFroqu1mtqHQhJT7313mXGGJiPZ2dyIoEcQCmY1p/3cgfE9GGn/E/Is
SYQa6be5sfGGBQKQLnIrBwj5i3rt1kLk1VqupFZS4GRsabg1CTUujqMdIoBBWHIo
rmnZwS/shIEbRNMnyx4v47C/wcFdsxD5eFKCRdtlNCXTsMd4gs4NDdQsjhdsd8oN
T5+PjBGHQSZrYbP3IZt4lYtjNwKlwXo7h38QoFxOED/YF8l6RZjkdn+4DDwAoOXl
v/rzp6/GCkdSEiEg/va5lg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5424 )
`pragma protect data_block
nQK82fw0ee5ekwVESU4Y8SatKyEqL9mZJE3xIJw8OdI4UDCSQcyAJv028a5JqP9d
g+hrbO7gTugi2l3EchrOwRqfq4tcO65d/X1ML16WSQKHtziQZEALGnbQwdhdGz4X
y0gtIKp4f+kcmejLrzp0N/NRVU5aSZdZHTVaQl6niaeLyFvR+K6Qzx070T3eWgfY
rUszPBW+ciWcLo7MdxnqRFgYDh913il7woKVQkXnVN+kyGvAKFDMrJym7/zRMPPV
V8o/TOXBxVJx3rgYvqkZGeZMvvNo/LVogpJEc02h3pHoETdDt/2O67F6TBC8asnY
naEW10NafspfkuzhrEJnVcCZZdnwFWC9meCV54+B7mNll7ItvBKn2WWRuZcwD5UC
fqWIP/uOmRdPfrDFkh9TgWTZmFo/hUitp1IY3pZ6x4yMj+/duwhFthCuh7hbxoQ7
2e5CGXN5Ele2PFeJ8nnx4Xx/tNUgXrk+1gj/f/94h2wrzl88qCHuSSEhFTCbuwwM
h9n8nN3OXHfHeaRXxdA7RgRnR4WEqiO8Ia42IWK272yyqiJ7TVL5DST1T0A02Dpt
liaQ7HAHtqwczQdLGbmEXgwfA6NFlo2MIRI6OVYG759tvoND6yfG1jdoKc2p2GH3
KexvSR84G3NH573IJxxFymBEiErqOhLOmPtkb2zl1mDFwAx3ip6iR7yZrVe+beVt
xJ/VFgaWeP4Pnp36TM60HfrTObahVALPwPtywwmyT/C6Ewfa4SXDWNGP+C+utehB
3gURee/CY1rSaYg20jiOuSDGKxFi5LGtgS0r/f2Qic/ZwlWA8ibfzWjd1DBeQm7G
a1UyXq5Cuuuhr8o+ZM70avna4tPfIG6VgF+unwDcZQFMmC1DDA19gLrlapWCK4Sz
y6OLtdKDJjITQ/RIxaP2BXMi4+jZvRp4UT+Rs/LHBu3hZzVyAHv1y+VzxjTCaauA
9RAOkBfJYrFp1ZAGSTCKNWXhQOuVmlO9DmGEiR5YlgGCYeY+hgCUciiXNLHEJSfd
aQ8hfXyZiym/W7LKar58qCjMeNDq6LZ/orWAioflMDYBYyUqgyuIt4w24d96TX0C
XuNrlRqtLE8P+lUWc3a/Nr7nMpyNyUJjT47Lg0ChIobhw1EGl2n6qdCiEsUjHUAw
UT302BVh5WLZveOkLvd+V6K8PoJwhrq85vwppneGMo3Wn5ntS/xgfLU5J7ztDcsC
4+17+NWCTPO1ID69NVJvSe9i8psahEcC2snvx+OMPw6IBUnCGE6ZJMi4Sb2xyXP6
27V8xbf8oOiD4udgM85oLtYCLukdtKfiJ0Cwhzk59yKxN79KG1AgkNOH11jCKUHb
Fk5Os/epZGci8Mlb+T9keoYimWP8LdS1XcDs/cZARHslHhomG+yMvoUThq7S6/CF
ZAelwmXGuWgNCDtipebnEg0hUAQW0BKBSnniRLk7YMyk/sp1cCH+aztGztHgEH1D
YBP5BsPjTnpLiGtxIpDMLDjCsFq39CS/Xh4R66C8yzhX/hIYcNzccIFF25m4YrXS
TMDT6LSVq1zVYLPDCLfKMxLs+j05/0Y6sZiJjDm7SGQeD1ZEZ0q+dq/mYgGpVxsx
89WHHIqaJU+9/W/V8SU6A2l0z3HNcqAqFPsn40L4hLp5YqUnK/DHClJIQibz3bWC
VTAHotMrroIRL5XZ5tU40iZNFOyRIppGH6lIvzyYeOCOe5tbAgATr+XbsyMhLDZM
JHIS/jSPLincLfll5b5DbifQn9piC9kYR8zrdngP/KNduPL7/z3tFGiwx5Sii5so
YUbft2n7NzFjciYP0rHLV7E22R1skaApY6p4YWN0zXr5e/EEkAMGKWc8C5ZO1unb
VMVI7zZhsg7NsU3ERypdfVDVSalPRLP4IhcZmXicK8awYvea6PaMSwflPzsBG3SX
TDtBUzEkeY5n5TwNWcBUm1KfG8G90ea0Vgt1QwvQZx9dqjYxVkVl88eIG405j2lI
bcDksIgG5kySOrSAMXc5trizmPbVGntXk4ItS1hc6xcyNHqW4Nu7ZveyAoGk5pmN
oo3Ei0h2GJoafEWpDS3Bqf7j9RAHcuyUnhiv5EiK/nu9ADt+w5OVhp+SJhyXWtSw
Buk2E7NeI5nJeZdoUaQ+keR+/Kgy5dF+/o8Jy7u/ACSQFlG07+gVHsJAn7x11Vu3
0kWbFWOi6Wz4S9qvvfFuuwaws67LFteF0aVWYgcfueMsYSScMzusqdKI+yjF68q1
j1nsgDoie4hA62R6Ly4d0Z2bTEhautaI6v+3ZAfhQ8xHos44+MkL3GaWyDvJTycB
Cmriz+x66Xot2hHLPw+3n60kAR4isPVBeLqE+QFjRsnY85Fzl6GSNuhI5oD5N5l0
JJBoe/H9mWct60IfWiCHTzkZyPzDKPmsqjbuzGNXFIqs9fbGdny0zA81xTSdgWJ9
oXlxwlvtPwG6oWqSfu4A8GzUzR8eb47xRGDbSKSerRuF63uVWMlzRP1wGXreMaXE
2q1DsFU8CSKUJ94o4LCZbp+vhcX9oiJkrEeM2oxwZTi4PLFuwj1bxBOauqEYIYCs
HDLWmy268ArRFHeLn4UVhyVg0b7qI9GgZ4O+g11Li7l5/+61iGpl8dE4q02cLYcU
g2vM1NyLWEoeuKZ2JnW0D/wYTGM7xhO8IdcQ7OcDNaq173ucOyi20ll3L9m1mkZK
yPnw8polkOfl77IXlR6l17aTIWUOegQ8LywWaAOli8w2Yb4EC4XJaanqRePVsX5E
Z3J3Dj9YO2AkX9+XXITpp3Bm2pYdBEijztjAhbG6/1A8bx8++eB8W0VrzdaxTFUY
MqGMSX38EnShFQ1N7FVszeyeTEvNATAGiqPL5aQHtrJlqDiSU7AOTi6OC2LLb+pW
3JMS4Pv3tdiXRs/7B1/do2xj5KijZCHok6QnRV4NcRch2aZeRBs4NIPLb7fytwFq
C+a6HN7dJjz46Uj5YAVcv//tPlB6ltdMUr3WUBFXd8X62by1ALnKW9pkXqhyG31d
NvE7HmqlEFBjYC0ZgIJynfP9FxaI77fKe6IbiYmUFmrPRkLR76FIzCCD619jOqUe
FBVQqEplIaPddDveRXhjRO2ByYdj5Z9eCACTfQErnnP9sE9+uZZSNJwoT3H16AWq
lc2qa6WqST7S7ViLL4xiKemnU/1HI0sy9hSSjoGrE+EgHbIYW27wr9Czh88u58Wg
ieSSeJPKNLyUXF0ycGGnsxDWzRpiyLxKwWnTPBvWV5lbRfnhqhAC7chXKeTPIP8I
iUhww/U5OrNZNO0L3A9Tg2bFMMwx4dlitgrX+5AxsaIlyto53y9lEukuFekbipGf
iXj3gucGZDjqaZJtbBXgqEA4tUtNAKriaGyX30nm2vogkE1dxYvcsBFtag/S40YP
RcgaeooelfHdQt3KONk8m5SosEYb3Ag8Gh301FxemISOgq5iR6txU1GviBrYG1sm
onL5hFJCyHMui3Hq9Mwn2r5qP2vJM9PQb7/hwt6Fuw1wktEFeWHX9wJCCZFgHBHy
6e1pOqvTcB85VK9q4x3a+OZGpHc+CoyEk6Ly0+om4UNMis3OuZ3I6V8zz++OMNJv
Wc9Gr8BEW9cmSax+512MT4RdvVFAW7vMO3x6/pfeFAbSkoA4O7zOHpb/KosItCVM
+AmRwIAtJzMBnn6kyYc5ygLKfBH8NHctA5P8OngmDv4f+8AarBEm2w00IjxKtRGv
UVQkEfz9HdqShayzfEGAgrltuMxenQvpBFN1FjxoDMaY+MvwHShA2zejf81bpor3
vWLCm7HuIn/6ZvliPEpQb5UaLUO0wTJkOsnkbwotoxOmwCn8AygwvRZxTDihTIMC
RMjDOa76fopN3dVS4jJ3LfzAa3bkGLJ/JeO2WmmXSv8H0S/SfLBMuK+6cQuC3gqA
TWNWpvGLFLe3MKYJ0a2iEhixdxzRs99d0g+ZCXc/79WBDctOOqMOMR6wP90kWD54
lZjgdpm6KKoN6ysKqi9PGxPEqiEvu5YOKMkCFZ2ACexL3YjKOaQshIwPRBv9zaVs
V6XA5lzfX/jJIoOwpCZ6n0DaZAQX2on1aThW5BEgHDLfjDjJbwR1ZHcwpwg9qgA/
R6XOf788zZlLoJg5bDIjLUJLFSoxoOdvlgZysOx/lUSZQse44U01JXsAtdPf8G1Z
jqxfNVfr9JplHGvSrSCxL1w/Gn85R8XV7bgoLptPapYO7dJxiAIIeQl0SUpZRZF9
A1crt/fHrcR8Uz2mMY17pfAaJ25bZ/XgMi1RI6ANXnXlURp6QZGBhjIDWpXG4KFC
voGbs3rKoP0ATQ5rj8l+GhlJHEosnc6QzvvCJMoG2tJqXincXNOtXuh2G/gxRlJR
Nb6YtUifF9iIh3lt2VkmlhEvdenoHjSNiJZC0SF25IpyCJQLk4A7H1G+hPXSWg5s
6Wy+chIjWC6IjQX3VYk71JarMWVsMzIP4XcDTQVYvRtxddzrclJzPFaZhMGiE875
/dcnIqk2lFsuxuRzMXXpSGRd2qFBR7mqm/BCYzmbCfxuoFydfbBcy5LmjKvd/qrb
GRSUokG7O2AOdJQUT+70vyUQw/ag+e222CMkRwuz2zVlKnoXK0e3eRREa7xz8F8C
kgp+36BiPPrqhffD/A9X/HaimQqpbEOfoZ+9AWR31OBF8Rldl01TSzpBfml09lzl
gpiRgXhheJyjquzqYmNpdwat6EYozyXTUFg6kywF01gabvAK31G4UxXAkWOHaiye
NaA/d/RYR3mQMPRU3E3zQy5zw8mYYg1A0HxgJTqArpMphIllt6Fkv1a/5UphpC7d
ezIXpuyd17+VLf7dq3lTGBSenAbEXn0m10KJdYyYZr2slA0rtep/fDiljgn+JnlI
SwzRHyaWI+cr1USii2pLOdzMZuoKh8FaighYYrDAp4cBEq1+PNWhWOQNBghVcOcZ
mrw1gBSoLTX3EgFr5FH/jpASWge/bJhBfKDk7bkIDMj+FnI1OiWTvWIYjduDm1RN
PtDq/DmXaCqXmcwtSgEPZQ/IJ1x2V/V9vKtbRpGXhV+vZB5sZt+qT8BtB2jv/RQ8
9Fu85jI9kCdJrZIHDlxH06srpJEUcPnsPaOMPvMPrCMCXTP+b8HZJFF1rAby00JV
HLtXSiumw8TQ6sZ7OrkVx2SLqgE6+Di8Vmm1LnR5ooZKFAD+PE/f/TS5RvM9Kaf6
62YTTlxgRdI27F5MVtAbgeizh13YY8lOGYDl8g71VqgUXGra7dpr2Blhr6ZdTZXt
og4/9bmNF7Y7qLfj1DZ0x6VlAew1+HLdlHSx2T1hijF1xjY6f3l+JcJ4/93nkPxx
VVroU+2PwFhI97wwPzFemfy5exLczvd+7ZsPNXX4yiD/KnCjO8E4ALlPwvMtQAwB
w6QHR+xUo6QWlB/5oTlEkZVmP2f5spZDYAXQA6cV7nXrTI5lWiCaxgH0O8L53ldu
E49I2HVwrh7UqODHepw7IZXIwzMz809sqMNGxmv8l9szo1NHWQDdlMblEsFz4eJn
/vYTtt3HPiSTTvCC1tAEqeuK2QAgoADSEdHj99AJPugez1kNFxI/DwvgyOf8lVGX
mtj4hVYPUgU0Qb8mXx++5CK6N6VBf/tXr8MFpBWx1fQMWC8kgRvgazRl2BFXmhxO
+VR84UkAgMok3NfcVGGBPW0KCQB8Yu8451d+GzP+ecDNMkptj3xErsku6TpySjVI
y6pQehlMcwTV3J90PgjQKlFYSBl8Gx7AsH25q6QnkSg6Grqpc4iZYMah/SbbDdox
6eIkpak+4gPWrzCUGAK8VbX+rDPiM1ebeocUaNruhiRtoL+iZA7eYVofhIc5LSuX
3iFV2SO7raMTzhLel4I87NXZC3RcIit70EOxG+AwNS1xA8zBymLcOtadvBvZp6Ij
P4utKqXY7/VgyVQD0tYuxBiujOPy84Au5e2/si/zjIw8QACfxgUeqL3xqMTYzOYw
Od6eVDQhpRFd0I1OfjnkBa7HcR0Jmj8MvBuVz83OsXFYsLZ405izRjVOoS5/c5fi
4VI8yxMd8nYxGQsVIGcQmrzExJVrvTIKIh/pqpRfooI98dF+deBNvhppE4jCdWeU
YfY+a+Ki8hHEVNnzfDCrdV1Ul0oXoSM3RHkKjT3+RzrRhp5rJrVizKUqbQWcnDl0
PLoFgZJI1MJuHcdpdnTwwYJ4iiOWifLQ1NOsClRLX3fYwIROA/EJNECAClPlrODL
kc/Xr5yWhMkC30MLURYsGbrAiK29j+3i88+01B+sa1BwZ5h1HTr556UKsSPVEwWS
LW1ERo7riucMf3iXhPbrQSvHIMCbtxhSLVXn/XaQ3FRgdeFZQDibxMDCai8Ktwto
LRPklDsmGXTe7+PrIVyYT72YbtYup1XhIdnY1Arl6dOGzAdaNHZqeggoFa4j6ibD
n/KDcgpDqTBcSHoIGkGroVLBecdOi5RrCD/JmZ7Gs4c800aVgdyTxipifO/Y+/pw
U1q5xmC1yG0myTKeFOTVs3Dul+m3e9LMMVHrjBjmozlK692E1MqihoMJp+VAKXcs
6Z7ddvK/ANgCTnMszCViY9wwz8RwV7pnYx5uIKSnr2ihWCByolgI3FurB/rEG6/9
06ucjLZy6F14iLB08KM5K0/k/o32E9nlNTn6yWG/D8h8jdubgWaqdmPkQ8wOfRC1
f4AITs2Id7ij7V5a+/XKydC1AMthMRI7xxXuf1R2DWdH/3O21xMH4l9tyvIJ9yB8
8WOSfuMKKpFtgh0/fQqENZTv2GyfbBO4QFoqppEBp5ObDc6F7/MUreFlLnHBKLQG
xXJ98xCAjcWq3YcpYHiVK87J7XgOlZJG/dpSptduqvwwrOjQiJ7zxlntFU5djnBu
5IjsljvCJd57bTDu/8MV23eYKKChNqcb8hMMAaOong8WQqDQ0s7PN/NHgwRp1GjE
h9chCoOX0FOAwTVX/BNWEXgsJhed71rt1RgWvwwT1z0KoELaIiB5ma3KYLAKV3DW
CbxVB46j8W+lhf0iP3A1nab/FtwbGQdT0ttuYx7nPy7haP/uYxCSZ7VAeyspvgiB
1htN3UuwptdGAZo6q5I6JlGXyQxrSHBNJpFuAa4vraDeT5nLa8Ih8cMLtNqJ/Xc1
AIdd1xnXACmVbxjyzxrAfYYeKp/JD3HxfCWAk4MGR+9Lk28GeQ8gTAHCec+3JoLo
fKevB30+DA8V8TpC9DP5Fc579lfcjI9eEnNDHR4MPUOO2GfyAR5fB18mDyfIIKq2
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
IWC3ZOk5chqZ2tS831XHzGHJ197Bslcs6Brua1Q+F8HkUnBT9aWkiyJajtEShZaj
58V9MCsi5ixLDgMkDBX9BpbYgCZdYkmdiT4EmE1hV/bECL0E33IvZLOs3FqOTszb
sNlYm6eq2CXqj9E7yqA/oUimlwkmqNKdEotELafIAaxI4EIpe11kZAHnqkcvCz2S
QMsSNv7xjZczic48p0Qxxc3UK5AtRsqjVnY6G8oZeSWJxC5xTaV+xTv79xIBiyt7
6KVo6jj9KjBpfgQhbJJi1h0y4TcY98ePU8C2VntAg3xIvNZNieXbQC+D3wkwsmgf
E85777RC0rsDWR9boVgnTA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6656 )
`pragma protect data_block
se6+zhmlcOkNxcZH17lQkJ6dURft8STU7O8QRToyxY3LwEq5osftCq9crLpo6oFK
7Ufhp8pt0sWfMqWB+O7ek80EJNGs576IzheGdA3piqEvltg5gCmegJaF/7WttPUT
+vXxNS0xsIg3q3w8mx2GJtCDa3621umqMtqfMvrTpSmMvp+A06Ll9kMavrwQhv3N
daGtNFbiJyJtUFMtY+HApQwD3magzoLTtXWuXMYtZak9LD93g4di1X5+oak1rQ6l
sHBNbKXW7UlOy49uTPFmW3CAxQxQCXEwGBxbfjmhPCiL7VIM7ctLH2rYrGeZJv1W
ApKWEDmwJZNEff6zKZ6ylXTChG60+SoZRy2bnDr9kJh79Xfyaw8blPK2jm0s1m3i
Y3uAVh+msWu3bE+C+v8epg/1qJRnryv+P92dO57BCZjKf8zOvSYk4etggGtelbRe
/QpYnlAV/lvKZBLwAlql4IpVn3TRYDZ67B5gHGXjiCP7v369rkgaISe2tl/MD071
TNuVJdXJxzIYyW6WMzL6iVCpqpNevNMGAegLKUwlWZ9zOu1N2cR6OUfuckghtDXq
Ihx5prRhbZOFA8eb4yXrLjLG6sIN6UkHo4zrohcKC0C2fDU6FXM6B18pK9/ABrno
JtdW4njba2TUxKwxe/R72tiXMPYNqWtRYErmj69emRBt0kiNGnhlFCe1b/Cjanxb
UyGNdgHMDYIQzWUM2rgZ7rwHj/78hUFwAxjlrUA6KxFDD+tbGG6AbRWNPyfZJbmA
84I/Vw2BHioxxRuprEVoKToSab+iPZnpAmY/XJ3XlZr1DGwb0dH5OsmTlmBLyEdp
L0KqqqJKx5S7rjAA5jdTCOG4xAioqB1bvGYzs7+zsLbT1xwjzev4Ju1yzl/o0SBY
EBFjK8lcGVHK86K6ZJplRR15XkOPEJ/vExvhEnCjnOd9LjKfDhDxDpJXsoiZPFaK
58DCwPBfDLq5kXaNJXm+bpzzKaIoXZ+VovE4vuTl8QnuRlOG/7JkONagYgpNpWb5
LO4KQOr3iUjzrhlHSfdZofarsccVJmtxhbNeEPLUqVNdw38b8PwHta+wFbjtGi4f
9fYJSPkzczH+izBlkdWZwlZJk50iD1hXWSid7K6ePixFz6EK39djaCXXub4tIoW/
XxxT4a2tDr2h5cxXa5vPoMRT5YfOy5UGPwXUHQMOqKC0qpfzTRfU/S2DJNAkS0Cm
z3wK+lXON/d4LO9LbiB4IA0bU5UCNp5ihIsfpnikRGtuIvDd3IOEA110K4oAq9VK
nrTyUAIijmPEOj3olI/SiD6lhN3sZfKkn3Pf0v1cITLpuUsnBp5FrO925iRLjnbL
AU0MObc4hNN+v8UdZZ7QuKh5TcIIiEfe3ov0fG+lpj3FSwGsH5QEe74KgbZl9X1n
1dDTyjHMGwJ0oTlKN4RoYuIp+JoMZkcnKdydOpAjcFzUcq6LtCDhP9KMvorbHGkQ
aT/7XMcsbV7xzp8xAbY4THFsNZgjQTdm8K6bOADGC97FbmZcqtOWeBzUujScFirf
ty+8kJGAUb1Xa7NTCosvoY8CxXc82csie+NMlpGgzpnRSYF5cBi2gPTFyfw4Xnu8
N4z1ivntANwwrUwaDtu3ZJNWILXiVvf3VJ301ShetDKUX7oSFoaUYXGBqoUbKVuw
v4nb0y6Vi0MiWxJvW5dUOtKs3hfcJ/VC0sq5ruISo8+PP5fMeBG7l0Bz+6fnyuF8
M/Y+tW7kw7EEjiX9rkStdLVtN9I4X0hOjUJbQSYVP/mke5q9xcRP4abkDCD69Nrw
oJygvXhCZUaNmFBRc9JeUXHuaLydCohpmaslOuwoQ12swnMrT48mHnQQtqrGvYUw
i5oQ6pkfgcYhnsv+qHo0o17KkyrhomXOIRDxYbQM3f00VXPcv5LRoGvyMagPCb0N
9FQHsxaYlOxhr2+Ou9l+8qXpVMAiDOywaP3aiBnBMNuA6VHlK50+FQvH9iUgK4Ai
J8MNUn8Q/kM9V91AVDeWmNzRDFyOra17DhsTeIsSK7Qc8aeQDDP+S0ioH6aHNBSv
owQq6urkp+JlhidQGicWFkxxfIRJanydILJTf6AIqLwJYGhc45UQ6jc/V3zv1Rzi
0Z/KYWevLodaUg0bS3jk/zveh14idsrAILmvEw91sZ9Emdqos4xSPPANVTgMhaYl
7Rp953jAf+CjgRyXac+HU3e0iJ3H5TWJ6a1DXR1bSYHT9VDKngZnmIXhNKAWmuxT
Ax713kn+d2ZuNxf7toJHRMRH80V8mq3g4157ntlQcZ6pX4RqN3d8nzOG5vXxII2y
gZDJNV0X7kfqOLMbLatJ2/q2aVhXKnAF2tyfCdfklfigVpGGzbulRjUJjOHlysEa
bwsOCJgK2DqYsrkML6fE/ktqBoCOEAo945II/ZEENH/wOJx3DoYecIW7d1dUpmLd
UV2D9bSM8e8fCkdFrVfLVK7X1a23beZvPem52WM0IuTKXHbxOhmGCPOqJ14i0BqD
MT/4V6CeRCWEyn6pAxwi9RzUSVSGo0gH1ynCNqfJopjUQ+dvhmrjqYeBRsoXv/3n
aTHfbnnEILy9O5dukqU5xMNbnSqBWMGAe7mFCkHq8YM3Pu28EJZt82wKJnVb6HyD
K1vnIUhBRqkysEXzerHQiff9zqMzVmM/q8e5N/7sFp84jUZVlHqlTCv1uMe8jkc1
JeBDuMb3QqYD0wtcCRULKdwPtpsliojyzEKBZ/UnfF8AgD8HpySgZhJ4+SzoOdPl
Qzb2PCeH5uYDuaHkwm8VJUa6qswWSov7vrZJd30xDD6XJG7hqvxOSrIRT3uVkzY0
F5U64qqtO5PaV1BdWQfW4O7uCkySayIcWgTFsEwiCX2XJC6Dz654Ri32O4yRS3Va
TaHB3TNVpuhPQp/eivH46MUn7uU1B4bgUmOyK+SoZAcQi3APn00WngyZYkMONGSX
Aq8r50O+pdBZRZBq6L+9ckA8dCP98dRb6+RED+qCJVk373v1QW+wVNWM8PBgTHhd
dRZqsUn+OxUhQtTgfQRr3x9eEmkRO7UQX3NZZJD5gMOzoBnJxE142eS7DVfA6gQd
afB1ky2+f7eBq8N58gQFrD8NTbYI5c/Xtu1lG38Rogtfs3xfI2M0MbqBXcGsLirw
W1255I+4epXOleN1SJoA+JabwlvMJyLJRnhiXs/TWH7P4k+lapQdmpVe/rvKS1/Z
owwI86UZJ6WhlKH80GTix2mqyGhFFqr8S4yqrzi+ZOyfC+besdhqtysiL78oV0bD
6UL5X7xS9ss8cE3rO49MZn/birY6cPpBg4bRd6LYLDMbSnr5fqei9AtH9/pLY6Dk
shX02GSfWSHGQuzUI2BKufdT7WUW6CJJG/bJyRhr8lvik+o8RYe+U/9in1bgi0CK
53w/V5lZfGmU4ahP//wuniiENStJYudZrN/a6NznyLwcHAwIR3og7yM1Y8qZNCq0
SdiWYLtPkRiwrCKRCnnvhJBswLwXZ5t15anrSRnGBIOMDO7m+MHZfwvLCgyn8gTV
MKU1UlimZncbdGSyrPHC9JggeseprVWBsfB+LBc0HEJsG/7J4PoYThmYDLbBBIkM
9abIWNVkyyJEdoBdkO2LQtUI5/8oHWS5Od85kSx42cD8n5NRJL+gyOKtXsrxujnj
hTA4yi5ohK+j0uwuX9lV3PuT/PNspBuMSvPV96KeT7rdLDs0dV9Zr2BCWOseyM89
R9G7xfxvDRLsE//QLdsb1njkqhU6gzSVmzNDNh3rDViH+UaKTdB8pZcLpevNomx/
l7TTdiYRc4fSrV1c9H3JMAH8ENqIV55z6zE7Y57QcRPlTA+0jwvvRRZ6Q/KPBEid
tPd8q4jzrXHayqnkIEs1ve0g6rgI6uR8aTSw5J3MHcqqLvmD2PZLHNw3UEnWKTGN
6FGa/g1CJf3Tkt21svo94eueKNZSxAMLFtYSntJZLHUKqzlMLKEteSSS6X48qcSy
grXTPtJnf/os05/q8sAEtvk6A80VmLaVmtk5cwCk+kK78rEXvARGFrU2sv14ZJDm
dNXFY+ndJe6t8cah843/dn4v9UcTFb0+kNiOo6icdXEka9ALlYPLfO0BZkUUqWBp
50c37rsSpFgJRShLN2Ksvw/7rce6k/AOhrE5kkXc9Xgs+MJPGZk8VN6jwQp/8LJM
Rdpd3DtklC50t8JV/QvVdTGmxrCa0BsaxE6xs3oFiiIJh3OL+9KgKfOa4dhKmHjX
flmuqziQDaGXXudyv7wfBZ+zdjwjMaq5D84J7UDaQp+O6cP30DjcdLwPrHzHeoPb
wsxAM5Xu3TKHYBDe7NDuQu2T+L9PfnPY26bEQhijisaQk+aC/pUIswcd5HnUfREe
GHOTd+GIunXqptwOUF66m6g1SjXTg/1cNSpqD3H9updXo8x8duPj3HVevJW0jgNS
0ZDZpDDLqVeIYobAjagos6ShmmuXpIYS+is351g8vJX33PDR1mtEn639KM6/86pH
0WlFRQV1VtbWOoM+bDCUxH5gXbgb0gK2xu3TbSO0NxDR4TKACw+3kYS6IyWJfczA
1h51Af2Uz7IgXn7tYWnbsHWEC63ULQljA9rILBJBzeqwYKYg8Kk/dGXYvDeBaGX8
4m5aeTShsxdORgqFyLKoSopFw0WE0dFJhAsvC9Z/7pEXlZ/RK4KvLcfgG3BvgG2h
jMH3iOyeQ8Ayup5tmtn1FSHccSFuGCSgo58NGX0YFoZm+5rtX7F+ZjvycaTOxtoQ
aqw/+LsVJRZUd+IbZnsnlF2bfvxkMu0z3dd77p0tDXqmO0xrb9mug02ktktgh8wj
cjbmQA3pG3PIpmaulQlRM2k6byd5OWoHtqgOP0p9F03/5CLlwTiSHozOY4h5lJ1R
W9XwoE6PB7ZJMd5ccuPs0/A2vYF8nQOLCJSns0+zo1ik5J0BlMf1LTdGmeXszOjG
a8mm9aeh/9pG5/ElO1KOUldehkZTwIRhtnHKqdXULuE5ZOSVg7zJ3AYAgpxi7ldJ
3iZV/ophpeIJcvaaugsAO8h+m8suHhw+eMyLZMLlAxCnLjNU+raO2TqQlPFn569Q
trIkzYrE1aQ6eJkjGUWT7Ag8fD1QJdMxoHWOt+drem5A+5v750g/Z0ei2CehjJUl
ZQZXE5QeReaoE4XMGMEgkPSF5nTv5wMTPc2oesQD/HozHA4gg3hmC+bFabUtI4yW
i7JKD/Sbz9XwVWlpnT1GvhU6gSOlQx/74RI/UspuT7fjD5uh+7RqDfH8pe1O4yhE
ripZ1IIlxM2ylxfJMdfNynKm1NsRzUQOxLOHLDZ5mt8bf8QQ4FY+VtiLS1kGFI9j
izE3fYy7DFbKmTz7GOqVtjQ69fV1UdjD3kvm0fPKJ86mjeIP8o0RULJjsuEK/wBa
2RCD1EKfcC0eA4d10ogq7GAEIe2Ekgip8mLDii8LnoRMl9DYn/+FiPliKUGOBgd3
YNlV1UHgFGlgmercVezh587mTcvZzVkKvHwjkwPgU1QZbMvWBNWnXX6aRonUFX9r
tGrMPPRKyVEqePe5ebQ95vz+hY86iEeIXpp9q/34Dg2TYdOaDjuo5wczEgStdInL
Rj0uv5o6OHV3tuO+BwGTLB48FQAoRftepURGjNmsyReFfrvhYA+GGtBqQ8TkQxg8
G1ParYyjxC0O6oyIXtDX/o/M56MVgOS16p87VEt0Nx1ZLo/Rixox9kD/RDWmrKLT
9xDkU0/JjiRB13C6Q7ZAsgpZW+b2jZSGD3Y2fJlD26YIThTOSOUv/qD0IaBafzZM
0zTaqXTjmhQf5AhLYMdWbNiitvDVQhh/0f28cgJtNzQm/km4MoU8r5Gzvaww9IA2
1jz/u4f5XFAzLTyPsHpjJ496FutRtnSgsQJfZ9Axu8H/o8M1DU2eHMfcZiuunI/H
lYYFxprBAMJiPf4c/NH6e3Chx1Jvm+UltfrRm9MmN0zR5nb1TZs2mb9ICyNGU++5
E3ukpOpDUQx7jaO6q1tVbl5edrNQKa1xpQc1Z+Ce3sgOCYmXN788EbnEOTDQCeeX
G+zt+ncbMssQYNBDeiIEOa9Ixfj9c7tNEPVq5PD2X4dUJCx0kvs0x8YE2FgMpD8G
WfON+nJfZaFenrTp3s3rrIGO4Y03Uep6tBiDKMKs2EDlOgv0aj3Z3AgP1Tp3BYUT
QFU6gm5DvpLyGYWImWihj75X78fgv4ZtG6j5XP5Dk3z3otOviTwyuZnBTiynLr7P
WHXDALB96BolMEUnNkLNkVLqjWr40LSJ/Q5saKfK8j/nfXKs1W6oNDbTaaOj5gmV
IqPZkURqyjMdGe23E/h2mFW0p9rp1FQl3U2A2Rnb2DCEr+s6vUeCIHhKrvWM35wp
Tn1bviDKT8zM9YIvtg8aW6US7r0J0LocyRp3qsKoz+SFoI8+19tC7GYibmP8Sj24
H1ZT8msd4uw8HEo2VQO37BXhWfmGB/LWcnQ0CLDvKDQByzDxxpS6t3alClD2zSSU
2YD0ajl65iHfzFyxBK0Kg6Ls1lWgZVl+aTR+IwDFyN8PqSLA1kFkEdLz8iEfvSkU
Vfspnrwkou52g+XPF0Z5vCmb9OFM7o4/9zyxX0bZs9ujH+gTkOH/mhTdL5DOS6be
fLycrX3YzFAMODwxcR+N6wSsBXy66cTwCjFo9NCH6ymInSaPo9rMqIb3K8QPRxk3
/WjtIfHL1VRDNpYaLJyDlT10UCGyHz7yWJmZc39LSpIBDJjS6ZQMtn1HlZ/gir53
vDHWWWpnn1TPsie9gVBITFi0W/hvGiWEgD15nt4UoDKyf88CFCYzAt2b80boOPn2
Hs34s1yIs5oS7cM4qlTRYySMmG929iAm3GcYJGpXxRMx8SiECdJ3qp13OUWcA53a
3RCDXE8sI4cvDqL+0mG9Go5CXaDqDwn3NVFOMWuOSsXhVB7ieALSTBC1vrJ46ufe
9scrMUnSoXRBuHkZ/4KNA+KBifBOxTaz59U1Mw24oaga2m8WzFEnNJKc+fTtlk2S
lWmXwLJfzmT/qCMsWmmtS1BgodT3SYIAzxbJtw6RtEJuCNW7kxlWKJeAD9foEQgx
xEjnLQnyIG9XUGpZwrllPwX5JAuqZfHkH+uyFVWf8sqQrltI0HcjBPNH2//ddKo+
Q+UjaMnprm5Izv1jNtg50aPNr8WTOEbnVZvZQnQzuZzgvNVqQtIdoEP5XGrLtyE7
hv0v1Hi7lzNDvBrBpNH32/MIVSt2iX1WMgCSF19WYbCcVYYa3W950Iu2bbjALspg
HobvM6QmuAjbyOQE36UddKviAbgHcCdT5MPdgCCUSNjkudtO3RE3VApms5jILEak
DOFcVOkpqiS0fQ5GUfJTENg4igrrCqsgCBRUiY9P//kYTKNvl/YPEfC+1RfwvljI
GVbfbDwaCP3LP7QEHvfNNX8PbxLIM8O93vTD/PJuE/cspxBYu+tzPHhoaC1Uayyz
NMl3RJnRLHRnATwZEOTe9Qb/A36IGWa+VmRxs32bHkHtkXQRUFTsAEpepzNWN7Fv
CbeLP+ZuCfhJEbRCuWQcR/B+mKjVKJcLh9Sbxs0zaYZCssovhD1eE2TGKcUn8zKH
v9IQ1uz7gvW/r05JuCl8PntG/GHN9YQwkrRmnDUp8uGBlax5VK6xWEwoo/DHBP8t
9QTEO/LXO86ewSLqMKkStBmA5J+I9O1MKCBiK6nbhgZddoShbfUlBMATLC3Uz6St
jnb5w8wSZmeqyre8dGXAbmtmrQueL7ise9Csbs+XmkIUr/+Fh3gY5XxfCZvcNqBA
hNwVh431BIT5yFRaKgtuqGkEK9w2sCB2W8a6EofpaH+uPBmEp8vkbIzFu0eBx65X
yuf05a95rQed7Yf/GNsFzNZIdEHEsMB9c/1LDi5HJ4FTjyQHeFh098DU2de3fQjq
wtTqqchzyA5VeomACkUiSgktj+JsYNTLR9v+BKExidCC/nE/ko1dzXJsIkktB7DS
wfU7DPmdi1loN2kJHt1V/D79ks1ohJGmAEYAyJ8J1Hv3Y1Ib3K+t93ahAW98pw1g
6Mg/2chpiDHi0xrv71hcFkcDHAR1KRgD0gTr1h753XN0wzS3JYZAyTsfT0HfJ5Ut
SbzbgHFpLY3tjuk7f/F//J4HIV33rX5dHbECHLj/Womz4xEl+PDHeZnklSz0hlgu
4Ig26m+67E+xIg5m5JectDATOt33ewNg4PM+cuEJrBX9HpEZPFXZy8q2UlqTAYZZ
sZLXZ1wMW0kGuu/OPjr78z9T3SsITIQXJQjVPEmozDmdL2ff7Z+9RORTPCuerYRQ
VgHj1ciXKdg8sdZSxh2XPd6axNuCowGeIf9fyODEZJ/1//E3pHy5PCUEn+TQl0oN
x3N8S8kWrkQnTNmSgYxMFeCM98ToWm6dPY1ZyjYSsNIF682PooCVJdhb8libLfTL
OBB4Sv6dntw/pPAaXhBT8cX48wcZ5a3zZAecTrD/lDrmf3jL2bUceEATvHvY9aig
3JDuibgTuxqcc/IyF15EzJd6g19iU0ts0HWF9omO0eOSp0FiH5q2xSc2jC/ffL7r
t6WKSMPYV3sLmEptRGKxXWvP+ecrdZIl7kNZjzGbmi5TfbSdr0VJu2CeJ00jBf7t
vJeagsno08y6BUxahu2/7Nxswp89rCWSsPKr2HVs0kDnA2nOk5W1t5iv+SOhsLVe
tCT5SXq7lPMNmhL8aAMUmTgnyffeG0P5D5i7LZvUwzBcgrmWMSmrBBTncHsnxG5E
rtzqQsAotConWWJk4PwO66kNwQsGgFkxggR2irXafmgDqySUcAzXPs948StmrWYt
rQSPxHxq4+Z6S+xIH8q9WzbjCYGt9kPvaljjlJyv88pfDWDF4vf8yUnLjuFNtSaZ
dYm9ANbOxat+SWrvGUI0IkWWh8UfNhKIOQvmfFU4sS4=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NR5/25JBpF93E6AvaTZcLv2ENbz1p3O7r0fpaf3ro7w4D4hMPOngeG+8uihff+gl
oUKyy6RBiF+rnZMBlDb9ax/e8CsUFV6AerDPppAqgOueooqNS4k0ayNjKoTTUYZE
FnG9hjYQQjfO80svqnjGTtw5oakMCisNpkRvdFaqnSLBs/ELklK8cH9sFL2nQhI3
XsXaO8VpvDPm3+PRVELuSJOSU2WzU3v7NxLa99/m5sqLIxi+lBaEA4haGTLLTo5P
gEEHwmrCP+Nd/XExYYflISB85wvuKxT/tUmXlAx2QdpjHTytwcpayzhKqnsEFG1b
3/2JC5s1bB00yz8Wy0aPAg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
3EHXiWogesYXEDCUCxRmtYZREybJe/l0cmRBgVCWk7FodH9vTYXuS4XBQ61cJ+ou
XvMjbCKm6Squzqa4xer5tJGaKgQzfoHz04cuTf21XB1FgnFdau7iu3+uqlQHQBJD
0QDjIKC8qdLgK2HJFWopDY2DRuckvkvKgk4ioK3oB+TFiMiVREqihrCWjwwNbNR3
c/24a6/8+vu/AC2HHuuvbzyD/zRoI/eyDSm6CefuUQaTdhGK95OcZdSRNQPlDjgD
RmpcTaT4yh4SgaFEk4OyGiOmay+XqadsbP0xSxa0ZpY5kJEnt42SNwP6VSIVdMCH
S2sktoyDJpngb4sewFnJqy2rbPG/jBOvBQEUNVdWcOxE98vf/hyHu7LpfxYhe/44
7GZSC7pvV0qvmTYm5Ntfba54VyLVBbHotBojp0bp3dOCsUBQ235/S3hbyqlJRAIA
d8mUNVWRT1QfSY6RxALL0cH3G1/Z26tbEjPG2q9CzKd9dQo4Ikm7kqfa5gGpaJOh
1Z+gPnyhvLQcpRJdiLxO+jlDzmA8N7wRCMBfkuVjAja8zZ9yyaczruTIuhhf5qWt
eVtaqroFq/+yC+ieEobxG/TCZpvgstvPJtBrb2k8zHcpkv/zbJ+4AxmBwmJlDHlC
cjLTqqL6Wh2OzHam9KQ4oapZgVdeeoD2w307+yPMF86LBpUPlH8YCuxm1ffNNd1h
/h/iqLYdt/daNHj5DvZv5PaifurR7iOiIc8oSpu9nHBskSZFO5MZ4NAOHSc2LJSY
7oAOjn2McTHeBNTtOUQKq4jDYDxXkn7jNadSFj5Rf2/IMQEOPNkN7GOIs/OwoRZy
PJzjuHAd60VPbLwCx6H2U4FbtHmjpU5CRRxFq5LCpxSTxTDloWa0dqWDJzHl2O4z
vDUH76SwiS9H3LhVc4wc/93vtVollAVpeqvZmZntv3euuuUiYbuPbdc+THh40MQj
7ufcThM/HDtg8c6C68ISW9/zncFBeNgCXyiFbfex3f34PNKeFQlGGafjRhvmYnTk
jgj0LH/irLiG6OYbMGbSjr7w2ocRj7unuYxMUATOqkvfasXvXVRvFxXT4QgDOJ+/
wdlR7xteLEs3nl7Qzo7j5eFkEtGqOYKdoWzc++vAa44LNzDON/Nl0oA19fIwUg9t
F+wZRc8eFWGpcIXYpUYXL6TqvN0Oxtjc6pY2QmLUzTCTX83ICbhxFMF7PHUjgdud
dr2LZuYjNI9Fa1/i3D3RMwg3yamDe8l8/o13MLjnojyNTVjGWOtYxsK7sbgF6urB
DuG4zc7hmsTr6tV9LW4V3NY5qTcHG2hW40FyjZtrjtRP8W219HxYYnWHPykJd+/b
vPSszejzGOwhCBAITG/gMDSnuOnmagt2HWB3rXowHas56fccLBfAbYhq0gACK0E2
8OpCR+RuUgU8O3i4UJPu+58ApJISNRQnhstlpUpfP3KAqkVI/1mTgbuRR8EzuZ06
bUyL7hjiXboozskXeFVimT2vovqfHry28NEeHY7hTKjsnTh6PbUk4xOO3vqLDfo2
5uP130+0E2sJioxZAfQ3p/HbTzU8rB9+wEf/N1nYsOuSl0yOwTKW3W0UzV86hBCn
EVLEBYZwRGD5M0m8u12lyd6gBg5bb7fCMh3JearKTO/IrAJ+vIyh5/Pi/QcNCXvC
djx8IM+yho1hC2hRjk0YmX8Zi+FUEXK/4dek/GFJUfhvTrNT7rkzWbIE9i6Hk8v3
3tKZTrWKMUBB2NgX/+Y1lRQ7HBCqaxXSCrdLXFAfev43cNVw6fpUK7p6N4R9a44e
boPMHNN6mtDzeOrZ661jpl/UEKR9Rt8xUbVL/1yf7xMexyLNa/nMNFxCANZEyde7
LK0OtiUB1lRTRY+BrLryA/ukIdI42PGhVANF8kzlgjH4dQAKwTRMQAcKPS9dd9Av
GHRVJQboMeyriIBb4j1mtMrNyRaBYM30wGG1ZmxUlKCKR/szN1BdX8BdRx5Ap9qw
If51ZCrzBo2ACDv18BFpM0FFwPMbcDwAyye8Gi/fa/zJvflrcAzKaFTO9ktOKKlb
TJse32L4px3oa5NYkEy6ve884wcgLO0kYSae5h0eOcuf2Ot3Ti627IHw6N1Bpq5C
1CYbriJTukBZ+cAupzeaSn9cYqKf8Ssmu6y0kSWhlGjdIfAqH6lZipJGyxq3rQwB
ONa/jrw5+QsQiGhQhaMaLYD8f/kfXnam4In3ozky7YQBscMC42ga71IISGTkTSkh
9JEqIxxMBNpgV0pR4AS0kOnF97c36ZvqmJ6sV7UadSxvZNX+tSxrQpT7h4pBkgbp
uLyLa2+gCf054JqzzAV5F8571LwoN+0fJDS4z69TOrnyknK0Ctjzh5cYP/SaUtF9
lHF/JFz8TedeQrzbvaAed2jCqh7eBSVrBUjFABfcvOutmruZYyEFgEZT6xYzCojf
nbIE4WCuLo0Eehi3lY0Bo6GcA4LcVKu3JO+5T892JFT8TY9a3A5NlPiqB/mRt7ZA
lSabgEreVyyB2uXFVYQ/gwPQJYoKY859Sd423sIpVan5hj7GLMGq3n4kTPEEL3pU
3LEiAmsnEhMTX48++Xh1I9+xELaxXYlhm4Mu7+GGOXQhF/8JzxqyWFqROKTgOYa1
Ao8UJr6VQsZ7zzAM6Q2xvp4hNYd5MO1/0TpEmFKTq3dfxQoVTrVihz6AEJg6XGDB
0yQaH7jVBQxyPQvbDopukIUjJ+mxzPuNUJLWEFMs02H5Ob9mANTAL0G1SttXKS6H
w+zMD5JBK9MBMSfVK1fHlPuFW1wGVWySSLZDM1fI3ab82WH/nSgJvUkL76tZIIua
r1uDyJ6qp1j2iPF+OqCqBZpQ60ilsgiUPBo5jHBJhj1BdhUC/PgVHnFNyH1zyx2I
7qYO07hnpaSe552YGmEQbk3EPCCA/5ZbNZ0EiAXkNBHRrhJfR70TEfUVf7p+vBtD
HyDsOL7WbJafu36i8oviPcZAgkvcIZq346wO2OGfJaA+Zw7CsGpiLjbMPB5OSW/F
SHPB63bM6ZYoNYkO3ECJA2VmBEXQbHntUTWebvzLsHZJpcJixnD+bwkaueYhaESQ
BLVCPSEm/Ys2kWtST7vqx/GtMLmWYWyAUWnsEyoHVvzjNGwtBe+sG95SSYajCj78
DRcF1F+y77vkVN47UEC85222UCFcsFUwQIQ0Q2V6PAzAZegl6HkhX9GwR4NTWC+e
8pg1y+T3t/00T2FivEKe+KJg09aQJvQh7Ozif0h8YXUiBzviNnwuYayOA2t76EFb
e6CN0nY2W23OacSmPhO4sPg8tNVi2oNvP5wPcDUz7WIDI2o2pvjvSsn3aQPOh7+T
rOeRRt22tDs98Vhn32996PfsJwr6bJ+qZbEGe/RsFt0tDCNHpwlWUb2MZgcZNVVW
5a0IDs2ohUz+e8i2523FXBUzcvoKKv4qrFSH7nLzqpWSzsKxtzeisWzT4yJ1e/j8
5IBtVXQvn/bMU8ARebU28oC8Ynj+OkbgpJo+viOQpKhZe+JNeeZXEsuQmm2m70L0
YVJG5L/A44lj5FplxRskGuDObO1DRCTBTTwZlSyKPSZE5D61p1CWXeltSe06+8GV
PRSBjIhz4Dx8kxPmhV24x11vjWoT0DC5qfdN2uNC/LTelmyy3sSs1eMnAIoK/gRV
sPdPBUx4f0Kkg/nejUb5KZEyY6KekHYCpELtM/TA7nFAtrGLOKiOYhPqtPfdWxly
O+oW9WcaVJIeIYElTgD38UWNjfpqvTA8THnqYx0Zh00JkSWD02ELwFyTCYj56VfU
c5PjsO5XAHHI4NXfVHCFIkpMunm0vi2ToL+Mb3RYu2hWWs13KXtV8mMZeCxgo8DU
gKDdfcAYiIL25ff/c6s+stuIHjgxtzyby0l4MW02OHOAAo6IyHATl551kLFSjC6w
uTd2V+i3idl3poKtjmExQpjUCEU/nzjirAYCil7eLr4+BvzURZ1DfJyDsWj8pHTh
Ol+xJ2tKNBnnqbT9mvr1rhBr8UFSS76Yq/kS3jiv8g/Vpy++KYEOl+vCSezhf2jl
icD4JaSwwVsWZ7oaCilVhfgKyhRiyjOzADTaNNo3NnR2KaCWA+guQkGhHLa55xKj
r83842YGgMsql0h1rgkqGjLbJd5S/qQiVxHk+L2NznCaz651drJQZ4qzc1hQW2ls
Kgm5NNtPyLhqh4H54E585Ru/VUo84qKqf7cIxQkYSAPTVpcoX7HqqTemCc8Tnq+x
5bPRgDuxUuiQRlyGOAu8vbIjIdgX6OLcO2SObvsQGKv62BBmY3b6mDLKpqXd4gm1
0KAXwM9tnZ3Qh3jXj0ZhdGxFMKN+6uxylghYMTls2zi1++F8kNSfFhUdkP9FkKuG
PphBwlUPq3+skWg+B+fEyS5PHa78kwWi28WIesXy5nwZrbu8twN0ZemGEGOGyPf1
b5wPwNiV9OjCYsTwTPsMSspSy5OhZ9x8zzVkrV9UyMYtN/PAo/aILSYglp/iUs43
MMdw5pAhkkGIIaZV9dGAA/HrPdnAf1kdMZ/t1jOcoXs6Q9aaJ92Aja+u2LRnE60v
ck9RktD+1dmC4fOuyyy1dnYvSxUFl+Pw1xGhRfXUtAVskQFGhwFfsz+7W3us49N7
ecNJrs9sfxKum0wzPoMHZWKTfNfrZ2cc1l+etkA3xsoye+IcLuDoESong7hLPKs1
Zsnz42DoKahbZ0rTGuntr7Jakz7W3CyL66bND2jehXyUWcuQ122FH21v+geVBJHk
ZajdfwhJGxSeGS+LqLmFDxrmYMNwCroC1EYvXZlwLCry9mqi6VuIwCbe11y4ulyY
ruJKUqZYUFcKPzqEUl8vodRln9l5V6tEwAY/OwcKRsbkAEWadnhcyXb044fnk2tl
6pYRUTT8g72b5G+/ogGz5pbCx4l4Ks/9CNA4vIpMQwN20OuPE4dzTVG9bpbOiMT+
Re4gbWodB8uhjixA/cfkD34f/Lmmr8oW2bioSdLYvQMgm+hTOnGiOngBLc7kgEs6
kqGHz9Pin/i2pNW57SOeYzjc8aVlkMYfocYyivjdY8cbylRRyGEzGnJkP+0/DsIr
3UKZwQ9/j8x9h7x4JJH8QtslPGru5Q1J41wo8iFRcblJrW2xn2oZ2kmkqrf3IbkW
BW8FmhfrsVx/nl1FpGAC2Xfzld6IyFQ+snAYQeEpYtBuc1Vyu9s4WUjUfuAFwnsF
P3IqG8NZqxQkfxiVt7PJK6xQ4DuThIzqWaZixTvoz4xTl8ru34a/W4B8Vea88poi
e/wDP3Hw1N6YKNiHIszFODamc8NQbSt1FXSbrYqTWV84bWURnbODWYLZysvEIiYe
D5QTS7kOpgJZCbW75xl/Xwagqs0nAElqgc0MJo9cVKi/Wx+cO0R+V13cq9zhp++L
Cf9EMSEre3mKTk2XLZ80vcE0XDVyiQjN87YuyYk5eFg1+BeIp9U4NF3NAnFzub2h
Q17afpdI3p9zSjNYs94rmgKCcl8cTC1hcR9oXFKXUzkwyeju0aEvFpXE/h0a/Xqf
PpjahbDXp9Mn3s8TERrEDEj8e/NT0ZlWroXWVXvO3RRF7IkaPKCi3D3Kv7JfAxBd
/3B66gQxTuQ7e8AEIykpZbfyTaD0PY/qLG7gPptU5nFp4RxSjYOcm+bd0Iqtry32
lLYuTHyoQbCdFS0pi4XCRgjb53KtKmZnpfMo7mhUM2KBGX9emYJna/6+O9oCpz0X
AOsCk1n3J+ZeYNgDWl4IVsRi4DT4wurQtaASvRXIq5gJAO09+VlbJEOZpkpMnIAL
ocdzOy5r/eeQsdd6nyrEXymAWe9tDUCdf0oINEdDSVSf08GrHyXJ53I9LcLNv52S
ONvpTOVDaAPJ8ifaD8SCNN+gRsP2NJ5XlY6KZY4TNdyXnXxJXtd2DBFbfARMz+H2
dYUUQ/U/uZUV2Q8bLxmdA64xaKfre9eeJK7aUTqkl+9G/hWyzspy2UQE1MR5i/X/
tq6zcOBkBozyk9uniXiKjDjjvMRhdopHbrsUDT1laODrczJll1e2+t6Gi3MSvy5R
oKubxEakxja6pugOFLQMSoE0kJbOwFIF+vDtS9sEXszuyRHQQljimykF1aJSX5Gc
fWIcDy9DneRUrb+7y67Uo8rM0Fve3M/ry0Ii6ufoQBAk+WYm1dIxSOq3INvoX7w+
Axe3hwHB6C7GXtbSE0LJfwZgoCxMqoCgDtNPH1ad9LNQ0+3lQEWzH7m0dyHwNhCV
JB1bzbOiDGcselCPhUfZxIUvhgiQUbxtmaGHQdQQ7ncp5W2FDWJOwSMICgiKRPW/
TdtQT0F8zUGS18dG66qtzEP378b3FsldfH/YMB518LMK/KbYSKSblbSIY2UxS3OO
kTS1+P3jbovxWYbtGqKkvFfR3x0F2/KBJYDplotNGEB/XFeqo69fCQXaolq6pLQ0
CfIlm1+mcUfVhvs5x2LFzoV4Uuj7ifhwPGICYbteWLNDhhOWx8sx7IfanfwZmCvI
pvAe2dOzoqalZxT8wpz3KbVWczgADmncpRRPabtHUD6con6KsF1d2nB4jpg2DZQa
KIOKDeIwtk6iR2d4P5DyOIeEStXzhfeTZWAUypMYvtanaf3SDWKt8iG7iE3PvDcS
yNUT0QJbRPf9I3n/H7UTtB3A06soFRSC+gRv/b6cdKiWrjGXCXSDiCyy8Lj9R1c1
yTnitFbWh+wxve+xMxsemhK1NJzjcs2nFG/mrg3ZHK/xUodq9ywrm5NQvLpi+fdR
s2+hASRWsk+t03h6uUuO7bTLviU3TNvgTpgCsX/Y6xDxBgedRjIMdEEiyqy9lBT2
6J71PdO71RoPNtilG9yF+FB/chkfKGD1JDs1auSNvAWufZR4qQ9p3vUbix1zGN0l
t+BEPwIDG+v9eyoC1XPr5HRBSvwNtNvS+OuJCfE0C9QHsIZlKn2Wb+DBqI+Y6GSf
xdW2FN4Ke0OKY9JtiEYBbopW+jwTbK/gZT4+8HfoDRbUUBn7D+aVyhmTr9YbmWj7
jyVESfVcZftp7VdMjangN2Q0yUdB2xhTiOohn+quVnWEHRJNvMApc83iyA98ICaF
wxG/ICFcmqOwfu9X2OTmoap440gy9BYz3g5O4EBHYoa94YnkCtrGpbbWJhWmgeR5
hMHtIwSiM1KS1rVgb1t4kJusN6g3XjpMgMlRB16X5pDgErvxAr2MLwuXhP9fMI8u
jVnf5vsoXT6QYZxBiD33ass1FB1UxyoD31ELrly1pN7BFIJ7JJi54zJKJrVSNcGW
HAFjQGAM/noYCyw+gG4nBHWSj+KdqtOaWTYMLaWI4gTVBW2MbRQIhHW6+eb9DtOK
JBfM1CuXBbQHvNPSXjXIW3WE4IaK76iHQKDi4MUX7hVVdVKixso49sK4+XD4MS2N
FlXOiFtzJai8H7/Hpzt17PtIrhw9jz4f5yS/uaHaF2Jn9F2B1RW8SsVrkY/fbmEV
/o3aUiO8oK5Nku9A0QTKmwo1gfCdF9RewRK9m7ZCDbpQVXj576J+eMZ4BPXqcLMJ
woyg2zVfb93XmQdEH+qJlR1iBUNQzcL7YfnsJf6+l8zrgYZkl6qRvmhY0+IHWeQA
jw2xFF7d2PhO0W1JhEYb1Ydf96O7xyDmC+75EXd6AN8ss3yJ4t3HpzBi/PtGtXrY
6v2pTE3MzIxjozwNojPyewjSVyKwcN7vLOFG13jXfRJuaa4toVbAb7ZpAUbk1sU5
J1VHsFtk30HrSPWx+KGRCAV/Im3NEZ/O/5WgKe6/L72HonKTbddi0L8B4TsTC7nK
5dwv+U4917VKUb21mXgodhuDtxntxs+/A8Dt09rzxibSL3Rsu0b4S461CC5dKCow
ovKlMeIOhQ1AlhMkzKM49+iHS7CRqyExEVK38jJe3Wun+tJLqJSOl3GMwXXv1/rw
+2wIkRLnzP1KIGZCdHelEGu9ILxjXxF/vhOL6pXW3+u1R/wFza8suSvcparC7O0z
Fsg1XC/TVmWiL7FFlGxsgYFrc2hq/hsBKB3QmXsR5apEtV/OdfvDfzNNkZ0W2TwX
vN+VOHqdVlTyHYh7OB3qwQ==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dlYs5DI11itv9ASNwPI80cvlWUxHA88ElGPK30aytJRSowqslYLuPM55Lc2hALlJ
QXUHjPt+r8wXt08infFlpkvRcexExVbMKxJTmaiydAij+d5jPbOXnwRasJn4UulO
epgoaB0rKzZRnM28M3grl54i/o5hyouF7kvfdednoyoc2j+NzWLpXqKzXUqh+tnV
41MuwvhI6rh8JHToCsYASFXhK8weicZH3w1tXt2956zdFXvgj4P4khUKS89TdLvQ
hLBw1QbMjd8iG7jghDoTP6GbLgof3UitRcan2OWbbfCciM6N4VgZO+oygoszGnfW
GPJ9nnWtLa0CIQzEc/fn0Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2224 )
`pragma protect data_block
zBASmvZ2l85Y4aIb8beTx7LuFAqfHCAm6k13yhQK8rofLtdtUuB8DW+BEFcd0Oef
gu00KiBHoqNtoOdX7FH3nioe6K+//Kyv15r2HEX70rY+jBa3R96sHxiLahbQR+jn
TdHYwws3u8QNOgenwB69+a15ju81tpUeTgFk62bj6y2Rsx6AoAKh9b2cIgdlAcYl
lsA18yp5mbjW8W43fYeqi/rvwygixA/AkGjiML+2kR3Btd98VdSK6V+5MOBDIkNO
iW4GzSWv5pmESn+payd6J4KYrzy25BZJ1M8+GXyxGkajAiGuTH5Bc225hVn9BwES
BXWIRIhs8GtVPcDmM/Zzmr4Hp50frS7mgV8VQyKvnGuf2l4XZAm53d9ybnjtcJal
vX4pTzxumByN8xg4+pDvPO42yn79Muy4rQPGTU3Wcye0fiiTArdqo6kRvMt8kBQj
7MaIMD59vn/r/zjivWNWvtF5jJ8aIqf8kVGWzh93jIXrsoNnqQnNQy/BfU9fbnQl
1cyY5nzQst/5AXYRuuiv/n19+M0osIrb2aSj2X9xctFtX3+QJPeAqfo+Op3eN2d+
MEG38j3Wy5+feOzaniC6dPuEcPGUKa2gq2aCfUrrIrdNc/lgJzkO8qMFUZIAW678
fw0J3EFFVxqp97Iz5jjhpiXqPNKG1MIdjFQ6bLOHPAQDQd4OoFyvDWk6hJ0BunFy
ICVp6MMwip6LZPn8q0Zr4tEJ2rwtaTYvPx0ifmofWWX+VYMTQ17nUfwFIDpOpp6M
wSpmzihIdDuFcoecPNGCgQTIH8Yj+pzuQWRVNCoxvYEsbBCxEOymaBcRyLEeUkBj
CaxjfGoz5x7M8M5s8hwipkBjjo7jvKah8epiVil/D14dSLyu/fiZCQk8N7+yu3+D
fwIE+9MkHZHbbe94azu5Bm0Qk2hK5KUTx898l+83YQMPB7vCEboiVcMUH1GaPkKX
kI+EE943rJMmt7drZeM8UTQrmTEEMc3Or3SIHtWKL7eHeYziBC3+C5YZYSnrkc9w
RMY5yODOr44axzdQo+7eLW+xkHy4n3YpdvUG907esGWQQNXUxG/5gtgWRMw7HJg3
UxaTZZL5gTWHWH4l+59XdfJqe9Z2yrKGb1TBJ1gUe8MScjONOSliDV8SUvnwVf3j
eaVH9gyeamyP+TWtQGDGug9jrmXyidqjxbw9YiPjK2/P8pmvoPIsrZxDcVTIrx7Q
SI+cVYsnZnXv5E8FSy3fg706cjkpWOW3ufHrz1cji6vo4QqFnfJwdMBEueWD0o5j
ViedBCeJ/LmxPyvn7RMjSlsQKzt35VoAP2hsPURtKJe+qFBYvOLeu1EtiOB6vHtr
QDxIKxHNblh0FNfi2y+8K+AtTeRGAJY+2W6KSDinWRf8ZhXXs8W6xIPUsW0e2Zlv
UW5ObsSi334SMfddIKc/vsKpBdqlvgGhoKJyWLO41b3GEzCj58cxW3HJP0vOuGE1
nTz+70NJHFgVhgzC12a2dHBK2hvOgkTz93u570xG/GabEHg82ost9mJXu8dc1JJs
ak5ktGgBG06HzNCggVrlCPp2qzXRKPYQRbniDL4Tr17EgXrZ6M+gM86D/8J7xEhY
5kNelDEOiomMCpaEeJ8ayLGHBPvbXkFS5kXTQy2aa3X3MH7VlGAjhK03YVXt4zU0
CjrUdEZTBf/r12tyEzma3yA6SVnYqmLpIrwqnPTMQQFWKOMrnDHgk+VMZdYtuM3J
jqthS0UeH1Oe6oJvXIzecUtgDrMDsycZCftQfEX8h5utFE2Y+KDjVp0icDfnH3P+
7vyOqzrcnwwkSpvkT07R4zCN/jEO4aif/6/8iCTRBoaHPdcuogpn01ih450Xbi/Y
BJlbjMuRr5MKKuEVHF0p+ZNXAhhthweLv/HmKlLtDUMEvAoqn57jTAYtzwg9k8C3
pCcg5zEIE7qiGtp1Lnax5VVYuD/huYHeJHlNlIgZjS+1OWrn9nc30L1P6BeA5kPU
Wlaw8QJViO9P5DfPKNlajMwkGJA73aA757MpQy8RHmTeLrhaK8O2WPPd32kzbaFU
OShdTubpx3cTqCYZEdJZVijvwyOd8Q4Qe3hD8G2KrGG0i4tqmd475S6yvtInvaYk
8SM1XBYjKJx7QDWUNbxFz0zJW40tCRGzohFKmK+gYnGOXoaIIGcst7dxGTg7awy6
pP9x5bEaGrz7J8Jx1w7bU5r0Kk8wziTblGDFEbxgNWb2j9TY3Zxk/yBCURWVv3Sc
rD07sXEzm08c/AUR2ESL6mk4QOUr+tO6g/676p7PFjqxHD+fdCcqdv5PZCwwFVwW
BJQILyVRDjyo/6Ag0xDm1TyDfzjM1aKSd2yCfRu4BzXk5+2g2hpKdSTyhm2KwtQd
qRL//4yiyKwszqEiTCLfsvpPKw76MICC0d1M48nInrM/wnUYXFIg+gnomOiaNt1S
Q+jEtgqP8DU98YddIkONvchrhLGqiXvhfzrW55L+B5Gux1nJp/gr8tFBMvzcKWQP
r4J5fwemaVzcVmefrIDVBdOjF9sd71zr4Sh0pgwoT0j4Lf2gw2wZd3WyxO7wsGeB
Tgyi23k/0cw72o2XzP0MXsNHjsJmB+BPs21d8Pbwu5ZRBvqsABZBkgNDfgvqlnNk
Q8XDyM4aqW+MXEwtYjBIg7uS2pM9fhrtqaU1JEz0JJnXJviLyXLCdH6kMuusoAj1
3Qp/g+wpq9sxsW86IxkWQtq+kcdOh6JmfSYnqu2TZfve4hFH77MG6uBge/1ygkU5
RVXzwYGFTqcEZ1TcegLuBov/UrMn9brIUqJRzSycy+IC+SXxTFd5tqCx6D6i6T82
7YCtFVCgDl7IizgY8Hu3pYzb1+5NDRLyJ4DXy2j4/h/9kna4Q1obxDKgnWOa58td
CmbsPLBuFKVbPwYITviizj0g1NelY9FJuLvh3oqaz8FK0VFiAG39mIUz0RzXF/4o
iu9p7EkMdOTKII7T7qIKug==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HrXWfDwjyEWi6M58matq4C29CKGb2Ifd/5kFi1WXGog7a9KM8HxNvPIm4Nzln8SF
pd42CorFL61DPpHjbCxOsBBBVrTOXb2RwNk3OOtC2Fdc28cxase6xmHHQikybzD0
BO5PuxFVu8Pnm7JnnJGlVLh8eSpFeivAYNbB/NQIAH/8L6qs9lGXVdxVrLpxvZM9
STYHvixS2Q2vqNej9t65wo+iU+/IBC3sMFEerSrDZI/ebN69xXxQSbk7v9NcmFYS
CNJZFDN4x94cOqp0s9EY3f6o0UW9NkBnhKAY7kinE5eRjPe79sYNUiWMjj1/I3JJ
5eFF8MzyF4Inr90JM1pcGw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9328 )
`pragma protect data_block
v+K5Ug2SlPrS8la92slX87KpYDAg5uYjgAbpjk5HY3MfBF3y898gU+lfCkKuho2f
iAcxts49Av6sRl9q91kjFu4ES4HPAuT5I9601EYKczjxWP6/tsNCfODMhUhKCPVj
6pt4t++st5WLIwgokcEeXI/I7Qzm8jFkJEEs7crYJx+J1St4zsAjfTkHtbWmi8Hj
zU1tdMCfpOxxaYixobxzGUGxLnrbu7AZIUYrFM3EOBLr9wct/+5yQ8KE7P7GNbUA
byxm1lLaHyw3Cy25ECmfqGTaMFatrC3wtI/67GG/v5H0+VXFExjoc0/1L1MshwOi
cE9htwNMdfoejD/Q1S+xh7GeOL0Tn6Zv1UfnuW8Ir0RShR+VUqwtK9zmaDBHTjAE
3gK8WGh6iZTf9mO3JwlvIFpG+RByDr160A8c9NM2DLr0TKY6x5ey1NvlaQK8FhAj
xpWpuAyNOtIheDtSoAyMXQvykGqwBFr86LwRojQiSwXfy5UjGHdpzDLjakIGQjIy
nlbeaJjcVi/OZ4r8p6my3gokPfdy0iOu2fgxSFe/gvwYh6Ol8I8W9H5nE6V/MvHj
Bl9wy9lc8Cntq0tvDA2Xm7VLmBtCbY5L/10SLsn3P/qNDRXvJJv5k+6dF+GdDAOX
6EQ1v14qMnQ/MNyvZ0OcJJu03Rc6Stmb8DtH7+HX7K7YIeGMmOTLCswQOihXzc1F
YjLTs1wZEg2K1CPSgXSEf/yKiQeQMis/t69EX79v26de1ksVLoqBFG7SAP+hqKYj
Zmj7qKsdY+dw6gyWHapBXsvIhGLrb0R2+mMHi1T5ioYSLZDDDIJappkTmKxL2BmX
fvuGFUKIR68IsgyKvPNgD5kNFtvcbShFBWrqiuFms8YITrfZgauz2kJBvUAzE3lW
Xa5rKY5qXxW/XVK08cb21soMW3iyKvK27wrsfjPTAHBV651KQyFHhzhbSyCKlFHO
4R8E41/dgx7MXBoLFjOjH2UQg6E2DcPLiZeyJa+rHn5AhRT2nkbH+QG87O0NIyAE
jZxM47u22crHCfyuKgfldeAZrlfmlEyUffQgXOLve5ItmCHhbZ2ewEErO4qbrkFH
n4EzX1kdNYdy3UO13ShG24BaA79n9wYLI5NIviRQ6epl2440qphbNZEkrtc36Wv+
LdsgtdG51CZjPWCRAFhp3Uf1rTCoxW4tDzelBIkwX4iTJst2ss01GczUm27V67ef
7VDKb9TOhDHmKlrjJQV0qb+w9evM7B6Ue3hzx7ZIS+FyS0/pKMR97AdvmRqvJ+Uj
ysSzUUsvDtsfI30OyVN6qKJr0m3nV4sXXLCbow5aNdkaqa1sOUquXxAx08QrfACH
L8A+tE0nFYsmPesQRKmxqwquFufeUvLqRePlqyJPHQDx/JYCMoQpi+3FQWCShFJX
EGBaTd8tsjEb0BaNOVqa5say5jaIt+kajxkjwmH4RHdSVffPcGFYcd938Azy2PUk
Iw+mlnsGr29xGnPnKqqEzkGV7jt9K58Iu8/gMWWymTk2AenUe3f2GjZZFhTZdls8
d/nimKPt3vPSuE9XpuH03869acV+4X0/nMpsjbHd/2p5VcFQGzxXMnJJyeBb+Nre
Q35PKuPkGI/SwYUlWCHMXAvddWHlO/j6ZX8ZIVBnm7yzwOvFbXYj6/3io2bNjH7A
/NjKznLrCm5EcnTijBHGuxGZecnHZiw0n54JUo4iHyQyaTOhIYh7fdGsWZ/cUiC9
/wCAOU5L53i95AmAlLwBcmmRCcpJ0UpyEvMSalhgnbw2G53+GWdbDbMwhs5CQ7zu
dlgzi8R7cRPxcVOS58/GI1WRJxT4P9KpyirnWlxPPaa7oCxmACkaVuvkzxpIMj8y
BPYR/KYAyZ6UL+agnOEYYN9rkOfzAnRJjebzsCiTC2JNgiXq4LCIV+0HrjyI5DKC
GXR62car8gby+IV/Luv64w9ILycY+5rQaeWxKOQkBui6wi89eb39Rvruu3LKhoJn
KctbnvK/WIk3rxcwUnGQtndcVxNUE4lpCGFtoKqFW5ukoBjnVNRMNETFbF+qq4iO
31wypGCwKuss1o1tUniuScSdl4OXuR/YHKDBSv/+RNDDRrBtTHspSJPmma/1LK36
Yu9Ap+8siPvNVCyQa87ad9Q2s2OuEoGoMhUMfV/z7gS7DRTOElD4KKrnd1CdeYS9
0fYFkFTzLD3bT7Wd3YeXf4sDjNzXQa1hbmjIBF3Gsfc5DXzRK9yzaIxIRV7Pp40D
n9PbPYv6MSi2jkOKckWrmbApO92WLHy/JBVr0GsY9ZgzaNHxSWChnF6kMylW48bw
zGRtXHVkTcfapTiXgqo1Ot5HOXOQiWNb+Uk6c0nbxTU/lnQhYp7LHXkPcKxI7qkA
weG67brXl9niZKxzEvaVjdLDew4DjCR/+zwaAfDRGl56JTvbeGInRWakFm+jwspf
lNMma/e6rF/61xe6Jk+VldPqegzQlXID2pRWFhAuWWzFEXg8IVgf0OHtGdURC4GW
QEE7tJ7SpC3w72+xOWOZgdRz7Ew4udKN3qM9FZafaLxdBCRSJ0Oyzq0gw9R80wLV
cCVaF0DaJC3nW+jxDkd5M6fUax82ekfLv1C+fST/fhiAnBh7KoyEtglD6r5mjHY5
cj0o5ViNsb4RqDxRcv5deuVtRmQznQdV6V7oxNSewORjZGToR6hmCB5uSqeicYeU
0pXOmpOFKGDSXJFVdtOma/bf9XLsa75KNxi9FRam+0NrjzQUvl2ISx3O2pz0xzew
XZBvcmf4SOsdMRwBrCYGokxK/ofMwXoFbv0vrLk0U0joeAix9Hu5uTWT5nAtPKLs
njzIM0UxaqkVDY99tKnFZBOMVPkuaay0GKqoBQHSGpp57Y20kPs0ebwR8wBA4Zjg
xajnBYZdN28nJbD7tG89YCLwk2Rq1Xqc3HRg/lA1OcgWZh/nfAtoayh+zoaT5Svg
ATQku8HRjFlV5oRfQ+Buz0/1guHkKcW0goiofjgLkScs2JqRtpKhRQlq1J0et/JJ
gWXG3+zO+FsqkVxJoBj0UMokxzadxK4XCy25TV/heXDnRcRYLe1BbTlsIWregEpn
3+ZzK9Hx50HMqBezpobQVapxp8ueHKad2KGx5yKpk+4teqvWLiwYdxp/APLZU6sE
IOzEjlOQgq0YA0PrctGNVtU6OurQAXCGuD/AuBNHB2Lxq/lLS25RvYQvzlwG23jD
vr0pFcT8cXSsozrHgVpivG7clYKuyw2h6bdhyv9MO4enczldr9Coaw1JXm1qrlM5
8DywJ5bYkcwkenUtjYCcaqtfNFG2EkqWlumT7THQhg65i8cztQgDqQeR0hCk/m0h
CmvwzsEhzCQm80GP5XAhlnnyrg4tL6nKEVEH/Eb/XyQYIKOPs1p6LGbzOwKrOYpQ
5NctCMlOEvxizswGEsmy9QtBAkXk0y1xAdCaT4YOwgzSTG3Su9C7vfXFzCAZj5dQ
O5eF2JmT7f5O2rQYuVCc561nILaAcuAIGY9k8W94sSeKWG0g91XVpiO5u2v8NQ/h
4GEFedb1KTbiD/p33TdrV9vtQpOz5RVCXBQJ+19BehB3xkeIyKkSHgVFnl/bsU1Y
eemboBObShj62iSZpLeZm928BB7Ya0PRHiJFaqFRg2x6o2gs841XpxEqZohCNFtJ
rsqS+6/ExbI4XCfR8P5f1EKK+qhYj9jHV2iQ5aNLw1VFjASO3RdWH7Y4dpcfT0v3
gWRmh706WkJafWmJd5lA86uUppUxv7PYYeYVFPq0P5S2hkouwy08Lt0bzzQz2Z2W
XXho8ZPNMV9U5xrOkE6zwM5xWW+7nvVrVn7lDYUnA1TNUqUIjzvaOvxmtFcUHhGf
yOF5lAfNTOmaW4+G+exqQdKFkQYfh34yoCnXLE/palfC09LtUqWu1+6ZBSej0kJC
URWMbjhyw8jTk9l3TCZCTzDa7B0gYWhENPBdTGaoK3BOnHOofaYfbShaZdnitlfH
5PSJiz0h1uOii+Z4gNBpDFFPgQEdV6z15mbLS95WfZkjXmIrJAlA8qKcSEoNsQnn
SROgVLgnBMc9GXL0RCtuGXBfXoyyeem6Ppl+8HT0JbWaSSuxSBIBouTdfNOo3FU9
7/UuscIUDjDX+zw1UKbGL9a1trXnoY+Vt/UJvSITFE+kWHQ+t9fVKX8lG/e8QOe6
gy7Ylp9LF4k2xqrelBwzKe44iHYghLJrbkPWtjSfq9vO7Rr4bwVF0vMk4DlqGee0
MTqDrggGx3jIWf+FmbQSvFxG+9Cdl0mNSGZjtWMLCriZsfJP6+ZJxQJkgg/BZjGp
MrOTU/0+qFynTkTJDf+j908CRJYXCcxPUhsdVl2TNjUKlWn+G5nkByPoAwK+FqHe
enqapDrG6g/cLYjn4oGvu5lumDpbBtQ8TTFSDqJRIUpVR5O9k4Y9gawELmJeqaek
FwsQH/yw0ZwzHUKmnZafnZvUBahyR3xlgnWRmQJ878FUNqGgbC0ORDihwTxvk7X/
MsQePnoRk9xS1zuQnHeHW66QdE8MwT4tDF+VW8BNQQvvWENbACTdCUyIoqbBD5Hf
3pCDmA88ZGPR2ik/Vr02hkuTGcw4r9DrNY1e3fO5Qe6WEJPIhIDIrEWwprjOgcJ3
KWQ6hpxmQGt5rnz7WRfMKHb1S5aqtMjiz5Rhg2aMV7SZUviQd5BBmaXai34SHF8f
VW492T2BYFDushXDjPaWjX9GeVCYbRi40/mMDuID1Zxl1qZslW+XStQUOcbPc7kQ
bx8Q5X4QO8le+JzbBpwYMkciC0AvC8L0U51e2+zpuVX+RntsVNkci7t7nn7F96lE
zAW3VyP0AJFIjTOXlmpQ5W+rnPEjg5UrXhincr3N9kDhWRf6c1ype6eMa4koHEZh
fBRIuzP+Hrxf/vramKv4PjuIGvF09eXOPfmkc8n+4X8/6TNiRwDWpmobJ2lbgBYv
rLehqHrfu0n6STdSX/BCJcf5amkfJ+SpUSVNtYqjyt8GOZgzecbu0udk8yt+b0vn
A0H4OgCgNx/d3+/okUUxCQRjH+G2wpkqyckjeQ6ERNSN8JjJZI8y175Xn35CHP2E
w/BMxtr3lZuT5AuJbKDl0e1mCLqwBqJxfhNwfU2PJEm/n2yMMuApfIbjfC03utoK
KJLlZAYydfmGWI9I3aYnM2bu7z8SeXpPlCL7VSLhVLOW89Z0I37S8/JMJf4DlumR
uEhgpyi9N0oGhiCXMT1qkEUnveom2TZbIGoTHEXuAEb6vxHT2/rbzcdWJvh7pGcc
b7g7b/tL1j9uBvO3fKWoWoK7vTuYb/DStiAXnyjfOTsVjWnW5hnB1izKGUgKTpDO
85EXvTMxHWIoAXvZE7cqSGHCvzxnd3yo365BfbB+c/pHGSh59jI+tTSwxm9p1ke0
ZY5nPoj1bu7RV5Sj2yW9oul79UWdwjHKM+hJWpuOIDxgy/CFG6u7UJkSMmgevL5c
vtGTNLaY9HLCtQcN3i7FaTex75foAPsH4h7Lsq7qTnJSxy7HQ1RQUMDDqDgVIilU
LrLhR8Cd/w7mtWcl3DA17yreLo9Gh8oi5WlwGhaNKyn7OXPSFZNdgGhiaq+O4WXp
aM5xXIt9zUmxhL2fJbexuYWfGgiM/qluvZSdRuMjI8wT9PVk1CKJrGdjgxcETJyh
euXhKwY8927J5sGt+4CdC/VOY1JTgdFiWpy2tiCE/Kd27w9GQzqZN8fnH4qBLakE
pwKB9NWc3HDg0oDAmBCvDRuPnIjgxhIOb6uvMtvGLWUYcQATp7kiEmIeJb+D0rIH
NqCwIAT/PIRXwz+G8obbDEGio4B/VUrYlNSfF/KpjY0Qt8gR/Hk/qu0Xzlsj9ZxS
gmwR4yJA2MHuECeeylKKCwfANPsN/n0/V/vGfboGKF1AiylvapXFb17n/I6pzPKm
hfTCzX96WZ/CFrIOqCJCcZdVZpr5mcuQCGFwRHBlADOes1O7LhaIv45p3skyflNo
Wyvd0fKW96ePEe+U93qVS1Thk0ctksew9zEJ7QFSQMltPkI1HBTZBWsogFQYDbAi
gzU4/MQCTm2wjnHc+pQET88VYSwolf22CFja/W6gpOT0hzdBWQ8j7Ar1nwRC/ctd
zuv4wnIGpVHUaimq9kOZMueaupj9kA3eKVRwBhICsiAGiJFDJDLhJd/NuiBmRzHu
LnpE2LTbjRRUEfiov2iVdZg4nP5eFAiwHzvHzgAvgLwciX0DHmffQP6eONvBPyaO
ZX8wuLd6NcWjOmvZe+WXKnLlCj2RUcOufAc/IEjBflYJCPJqjFUlUOVffMn8m51c
IZx6FjNgWCPt3WEUq6gX0vzqEk2N/2yOe9r2mUw7XBOeDrV/6FK29iu7p4G6WMow
wf7/JdTzQyed4w/HEVyEKuipPKcyyW2LNZOB0GEwZtfJmJVNRGg3UD/HzK4t6y3f
cCgzQFM9W/Q526M66+6U/XcMBUTgf3l8FIExK1bKrSJG0/cyArNw7yvnPY08ReXT
F8xUstZE8ITFcis7aritkOmn/9W+XkNAaXd6B385oAeh4F2DAV2Kpoe+BmMXLh/1
65YqoHfGrpyNaJCDvrMyFFROgZAFwaR4+3k+68DXw+3smSbPEIkP7wiPJZvnm/Zt
3CnR6lvZf/AGwe3NEozLfa3aygu/iSb6n2VoKsLPLNkVrf7OxqDjMTaXjBAZr8Sx
Kg0KZBc/GyGJvvWpkTBo5CXYvj9zSTYL6YWM5Ht9VhkCSRi9fWacH2+JRuRWRVin
so73TcFb5V33NL0ZQeddGrx3+HQaP9hbmvFpiyvvgqbChzX/op93CN/8Gi3Eg3Ao
Ym42Mtl9Zm5qGMe3HMLqwueXJGX2LTex6JyVIg4XUYH5lOo+KNLthfP9tuTDD57D
ocdEJNlLTI8v7XRBb8kjxmtt11myPYh+Fb6HGw9mxT/qdq6K3pXQMpy31uQrsD76
4ZOQGdh6Braus/ZAaVLzXizVDydNHafSjngzGuF0zRDEmS1jDmbO9H70qyjzhyOM
bAqz3FlOl0qnEpjOpEHwDuoUMUHG4iP1GcgZTov+aUo/3bETr/Wb85t7XUJIuTsp
rMRMPHge6cmQJhQoO/0VPGPpij7bRZCp/HxB1cRDJX4NEllzyKDLLkJC885AD7ly
BPgE2o+PId5Ttly0R8YlzoqZy1O+akhayOfXe1MsO9DgzUQpTILTtE1Ege4rLBpr
a3GpKABGeOV3x6fsKdMsyLcKOLNxoC6Mb+j5Dl0lgy/Rd/SZ89ll6B7y6p9MbjaL
1TDzlSTFjMaXVCPEBNQgxc4XUuO3kBfZdgeV1Qr6BO1ZIl0wV+W44bmnsb1fKxhG
u9KKCwHCBlGFRiK4gvGphCWZBRDM5LVaaBqaktR1QhCsZOt35TGDIBWeorcmHDnu
oVkjtFrXzrg4qxxCjMrOf8RsefCwrgCeFJG1FnYlNP58KSmk5TI5M0uPnWk9iAxR
uwVPfYhDUUrVw4UW7o3yC3ezHa9K+eZaHqNo/us4X0qPuEWHiYG5uYrK3P0mWuB0
IFQm+kvD7bQfulfSMiMdlOoFMp1Pu6/DyXcwcDL2gP1VQVNoLSPd/L43gQh3/pLJ
6XxxBwblotAbT9k6aHoBVZNMHhXUps6bPbc9y5YItaLg9GhkIoD8fE/qP/m/bZjp
lxZ6prnQmiY5ZPiBjbXtwVKDt+Q54KnytVV5ULqTOGkMRJ6FRw+8+CYYLRmm+miZ
fOAR28S6Es4YcxwozVuuwgy0gGl8WvheykhNELVFkoPs4j7TtxgfYAi++ZTro5M8
Be8yPqkNSF9IR2LgxLY7seZta449o11a9WiCUIe7gcksUG6Ra2KhzAoR173nOtkd
IcNFg5MQTDDBl0E6H5PlwJ8eSlsWHN0jIXkRMBWKm8EAJKCiBR1TTWiwED1wDLrm
4SFZOd2Iz6vJae8Chx3rbLvi3V7uXNntvP9U+KWiWm3PhDhZav7aoX7+7IiRO/No
tkuMTVy+qRWf1+CUeKA0vvo9IqrurxUJmxTWfAU92B7wXFnD1leGfRwF2TBLHf2X
esk6xSBqwawUMDZuXTe4ku/0sRVlz5RcQH+elypLqkUtP9+Txalj7Q5L1S+QVDQG
Dy9cmNL4xcf1NeaP/MGPargVVKealgJo4VdhHhLHmiJfI1OeAl3+w5br7Gw4/XKy
VZoib62lOnHaF1MKplsxUPMV7MeISvZF26qvyY+lwXRKl06nnZjq7MqFwzOoYppV
jz/AIAxO1ZT2VLvLzbRipryT2EiNyNv6QhGJfzT7agWxPP2w8TIwSo/+vFdoPNGc
nPcDZ+PY/1uy4CmopeD+bkwhSTyDCgWkviGDiFluiaik+gj9EqfyNoSAPH5l8boL
GZL9QlQ3vKlBRV8j+uzVzhKkMQav0Xm/KJlys6KQ7Zq3qHwskxg1QjfyI49AFFj1
+PGlX6nBwMrrZEfi9DH5APMGZ5YyD5bx+SuNfxQFwSYhYDmUEDPkjsCWtM/A3Y8D
GSNqxuWzkR3Fgy/NEt/GHQ+/IvXHlOXatsLsaGI7pdTOCWPuY6f6qLu2NQv2A+6K
oK7SPICvaXA54DfJqoPxJWQPqZzYIncKNc488/PmQD78PON9eRcGi3MTN0EAboNI
qfGKk0LKXBcJdeFbTL37jbWHceFVIEL9oVyFyAP1Wk9r4Vf4xN9ZoogupqKDt9R3
46HxzttV1HIiY5lz00kkAGIiRXaiK65AdPGAJSyaFa5OqfDdBV4LiTGqGFWIqnPs
JH09yVyArpOwdGbNf1vIPOy0UfWdHLagUPFBfI/3rxpSZzX2oqqDU5A561tzzxJ5
MRfZR/LQ+ZClICAOR2nKI+ALuZRRZ5PPskclFzoWRM1jI8iX12SpIpvhrLg7QS6n
one2jsZ/24mV6+tQhLHzNVPBVTroS6gGH8f/uXHd3oP0a2ZgjZkAsZtwvUGJaWqG
x8k3dr1PCXwC9vVDcm7Sgwl2o1+mCLeQp1ca1H/QIAipXPl1Klxfbn7QQqA3E6hb
R5v9wbiEX9pWSGISmdVAX8vJ0XxXIhfPq0fgfXrhPvsbGQhWOKcnqAMmgLePY9Vb
2Lx1JttuIUrUEKCctqo/C1ObPU+K+gtUEvTwnnY1ki1k2gzP8Yu4OlkJMWWkjKNt
Q5gMC1dA2Irx8F8jDptcZOV3qaNU9WDHHoxxofZ0fX1Aom53nKQaRLfR+kEbWYvl
vJaZiVmoTfj8vuN/pwWDJpN+Je4DAcI0Osr0GG6PvsOrspRWGT3sq2oFIhEnZCCg
egmXCUA7j92cnis01Um1izPFq7lSE606fVqBwcwXKg9wtfdMzmVUQUKo9+q6isZ5
EwUactr4hiHiIWK1M2zJ0QKm+UNSbDkjynCPcw1vDF2vODv1YRr5LhF7tdjB/TyG
Qnvogh9wYTDUY2bDYHmPhpcfq54yXilbWhWJo3Uj56pgTmI4CjgsJhCpETa4MfLI
AN4fC9/eAZjpjOF4CMX+JcbfVwgi2UPpcjpiF5z46DPgChykPpNZbuhsE6AJOVmV
j/xH71HwyYH7tAR8zXg6a5mKrsrRLcm+6q4B4+ePWZSHzp0a4LtmOB7MuQSrab5J
OsXs36VTiVvk9Cs+fFwu4XQjxuiSxmkSGg7Ff5OZMRMH+yMnQDYgW+LTG2IphfKc
4rUuo2/mzJwwSuD6LlIRf0tWGgDAjHkpznZSA+F7TaUIdIjxepo1aRvGmnhPepch
wfb2lBUw2oPSOMTDdr5/orXnKXLu/4CRGGA9mnB2drMYh4xwrctxPrMGtl/y5gf3
tKZ72+1SC0vBsAT1BPlF1Qe0CFcfoF9tBZGnEpQUEZN2zHax5nyv81uAfHJKHwcv
2S7si767ZLbiw6m4Zz1QIGDR3nheKL5auWbXn+7EImvhXIMghshVd7pefmHC5cQ1
3lHreFwA2JJ6GO84vZGBwAPFjTZ4yVatL7DS28xwg70lrB69dxYEFDVPsfYb4PoJ
N06r93D0Y75dr1qjsKpMhE5kEihOOviGiQz99BVyRmrJNSMDhlGS7+YGTzyIMnFb
CvZT72kyYIUicVHCOKJ2HVOibKf6U2FIml2brtC0o6FnUqSkry4p86jlI88K3pRb
zbx1dZUWgvzzW3VBO9v8IO679O4IRC4XZYjN9jdt1MvrihJdbLM4WDGh0d6Md+Oy
OHxbOO+FnydqgKX0aV28s/Uv5beH0P5hv42v3qgMrlFGzLkyQwhMrgTaNdENlPf3
HTGrS6wWW1ShOsfwuYseDWd0jWLii0Nu2WBIXKzRUpnsMThevl5YxBMD4Nt6XOrg
urXoLSB1VuT33B4O5aIRixxKYF+wXTASIVvtRWXaN1lDnrpOXgLACIlSa8nvP/8m
aDHSe87BZdZ4ylb6wseyR8oks6hkXYvmPMcwiLdRAahdFgnI4s2v5iWYeKh0uK9S
TLt2EhEb4vh4NEXpZIrxmtavcyjZENCOPSGjG7c06xLQa7mQEPaKgjL3uNgexghh
TYKkcc0lKyVhePRFPsIw+LfpcF+f46tc2RJSRTw8FTbs5rs5RXIPvp3wZdPFYZ1S
YDh2HLYVntAFBxt3BJGixIONNDtJ/O/CUjk7hNwNH/J/yLBvTVXRh0XWqPTe8pAJ
jkRzW+zgo2kDJ7KRYQ3L9x1vqt8aT9C0fPHWiS6ybX8gXkG0jXHSy6T/SQSUeRWe
B4wO1LFJOqDYAWV6/jk9ut3fRT99GHfW2TgtepCPt7pJ7bEAsQ/QL4Y0MB8NkRZ7
s0HKYJnbM4f+NBwrz0h+jHf+gdzAG6+4NpoVb1n9hmLGweeAabrvMdHzvbOHbhqY
Agyry+s1bmXBRdOGVkuFJqRbgbEnMOT7WNtuC5sF5DuVatZUNeQQJxZN2ZWRoXw5
bB7rQ4M03LQhlYQk4IW6zDBNM4EiPkTZQ9X1Xe/UJ/WuOi9/TFAZz+fthlg1q0TY
IieUF2YpxDBKN3yJgBrL/qU0ayKzgPtrbWYewprR1AZURtAVG8y/edSs+xIKOzWw
yNyMEVeAXDa8GY647SC8ulVcFlvWiLPS2KFmXuo1sR8OTN1VN/YUiKEd/slzEf8K
lUnorCxemLlWPAp5SvSf6qFUba4+i+5C6rwZcNEokOXaucKQklMsa4gKJAOd1gpO
Uja7w0eEMvH/pseu1CTpp/HzZSzeBiWqBs8YWPhDJLGhP9oaSp5i/7iyOvvaFX2I
lI02ruUeu8anjxla5DB9oL4cfiTEjnfa6qBEpDsdRRAWy0o5t4SHB+lK2/45pJr0
p6MMLnHdAM8a6G8BiINt/UqI4MeES47z5yugVO6Nkp6z85eUCsCtD0IX5dIOLH7g
h/3HbZ6GHZ0l0QxvtdLtFnknyH3yumzi4dtItqd2opwEk2u8AcUVBZAzNCyPDA58
sriIcVry2x0hpS2meZVPnPwc7A3MJtTX5klCH+XEiAIXYZ+iiE0PSH+Q9ygpFxQ5
j9TYemHxyCE5Ib0nYqHZL79fNU156XFHm5AsirlY2D9KjMAHfbiJLau+uIiwJ083
G2AEALj1tXH0EtYR9YV3YN3XS1LskuWnjVNTqzSquYjeQfBMQtFKwRQcYke/pynb
kW06xWO30MONKC3F33UPKppEPOtvgt9JNZirPArTL4J45HoLEEy2Ha6C6AlpLTDr
SxbQqcQ13LA+qZOImEcINU6wSn62iSMy5/ApBiO+EMpA79W53Mm/vzx5QIwv9fi/
OZ53+tu8BRYiG9X5QkxVlnc3Dlf/+l1yNPVnI5i4Y8LQWJWWPmg48ncMEuS6O6tT
WU7b9y7UMuGTaOKjIM4nO4fQE3vL941aD6EGSs2Bxqo1GuuB1ow7mGtsVbYRTblG
Nly9Z0WGf7MevwMcfkO1FiG5tYAORm8O0O02qfQZC3vESPV/Jl+b0bnKIn3yAVda
Svq/xJ/APP72e8hhBwTHEG2G+J2qOhK0KXFz0NXnXrZPhTLpmLR0GTAbuHvH5yw5
nnS/hI+0UtFfREwSE3v+ifl3U2cLSKZt9mZm4PlehhOjsvtF6X7vxmpkT/UotAAD
7pA4Tl39WTUu8SQmUOhVpr189NQsjMUTO8tNfX9FB3rmNB4XdqtzR40SanJ1pgEE
JFrf4U1AB5Lz2RMBDzg+l4zw7QcfEvEBrLVhXsUbOaY8A8kmGJkXV4TLX1OLx7CM
qJD9ouJTJEp+4wh1qO50t5zG4V5UDuj1w7chrXhbMkVZwir1Vcd9DHRCdhye1Z8u
jRu5sTs83/pxBZAcSWcEAlmIIwO14PjJz+gPgZ6cWJ9lEs20vQeepvx/FycWr+Zj
+4dRmHNg6FiVX7M6d/1nVBqgbGMrjUsYTF/kY8Z7z5vDGvjXasc/W9r6HJ7XD+mF
7LAlFZDwAbPbYXCwTzI8A+FT0IlbOmaF41h6ScyZxJeTKLDm2fNhbWHuuEvhoSiy
OsYB5jSmvAgc9Bd0HJlAIbrhwNUPXUFUbuZar8EqW6vS6fA3aSGceLym4OQY1yqk
sKSLnLfsziHMpxLIFoJirw==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Da2Lz0G/k8mOOKyhO2sdyt26XkPRGDVnXu1joEovcS1/MS+/2wGrjKwzU72Ctj9H
cQLr/sHVGtyPVY5NHb8Ev1rz4U1LgdjjSqQkdbzDVEbhwzWE/9lM+yFzzhWzAOCK
tylDmemgldIafS2E5GuhrBIzFeEDih3aYkQ6C1lLdi7AkfeBc++aNAQtHLOEHh1G
Oup0ysq0ciOQV7nqbL+G6Whv8KjOff9y5HPrqOsLNmXioRBsYob3v5iuwj5MITvW
fZoslvASblkMDs7AhJZVNmHoOdNBBAs3nhivbHvuQc2yg6mosFphoeZNQKZIUjgn
Ym7fVQrSk+mWUHUnsD2R+g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6800 )
`pragma protect data_block
vy+YpBwOIR/5zaYtaJuQ0aJnvmRoJ3f5+Q7AVBGKODjQKng7MvIbUUMpUBls6GHr
WVZxJP/vZcVBZUug8S93o1VFPygJSShjqTQJKsCPFfAO5ws445Avy5T1CmrzFRak
byp1qogtGl+bTCbz6W7onRPy+jHPzqhU3WVtOBBBdIzm+3/ovtF/STPQ0uUIfXqR
G9AAtI7+cN78q4gD3XRrL0Ri/48x97ZykK5Fum1fZQ0hMv3MwuCSmxQWzccrSOvi
OptwdudvGz/Rlh9ZgJ8G9BRl1IRiLhd2G3x+YBZVC5vG0svJlP1enTyLye9kcT4A
VOs8RofAW9SrVAGESShMAFIwDLUHOvW33amaCU72jGwb2lXoDWFcswkRqexbxD6C
cRVT4SOg5XBcZVPXJ3tt3HVkYGvYrQ4YdcUF7zutGjPybIgFMv6EnBq9nuKSyW0C
AIuwdFsCcR+VIFNSPMUaJxx/IJhBJh2NwzPkeX+Mv8FrLb7l1elucD9SMIMqU3Xp
ClXGPrl7msh7rroEzq39l2/0FY/Hba2kHI3tErcf1aDF0qxg/WcA9OY51Akx49KZ
7ciXj1Ur8FSWkMp29DDzmF9usZdgj2rcI1oMESb6OgTwANxtfpAV+5zQjTgKLRQT
iHIJGj7ZgL09oUgN+NoGtEo/eQoePd2C1hd3knf/NAEf6z5l55yvDmP7dWrbhjGD
XyWRtbeeSf9ELqNW9nkHZ415PwJyCS7/11I4j9wz+GAgvE/nv3fQMDmmzQDCeyID
b+Jru3ocepA/6CS/b/akYCDZqzRWm/dtdifkf3W/L3JKGPLNePNJX5nGkTPveyjw
MhSOdIkYIcezT+8m09v4BUgsGDJdFiLuwXjfrAcH/FVvpCdnUpBwrGKiwYKXk0l+
V2jNhtIzv+obdAgTXJb83fPGLTPjMrkcvHe7yG3fMmBuKMPQ+jD/ai0DysUyxDyc
DfR3PaweUNolOVwSOpuUyspadZF5jxw9V9ru96IJ2dV1lM61yO5kpGrsL24HVj+B
9VdzMKBDnruTFxCendw8mpwX5F3gef7jW2z5NT8jVMe84PR072Umtd4V1o4dvhKD
0gr5t9lKhlV2/2sSbERVv3CgGZk0SANfSDkGzlffzhBUS0OrMfTLG/+/x7LzcGjn
JHZnHi/0unCZ749rUMl9rwXqIVC9GT31IVSiuyxufB5f62kzzqADQ9aQ+qWWrdvh
LFI3iyppTGEULPeTyqxJFcZhpQXwOWtGdtmZMgnQX53B6LJ0w3hPbkpu3+Aa6ZD6
G2NUUwLp/OQ1TpALPau96iUGcTCX6R0TtToxi7jc6xsPnBlRdHvwTPqVF6YyybEI
+ym3HbekUZ052Hex09vabXZjA8mAgLdysc8FRvU8WEJ4L6pZWsL9M8QMob/jw/BT
4FIyrE1BCaBXYuswJVG5KJzyWfijBzGskwuVw+J+s1YvSvxZAbXYOf6delXpmoI+
IdAt15iTUdvdHWZuJinCZhTguYtal98hQnvCLRQoPWIkKoAD8XqjCv3B/vxFc1Od
+vHpyNdPHT1e8P4nUtqFgoeWF530Qkz/iUND5B+6e2Ur2cJxmjyUyMUhCByvFzl7
aWTiUvsrm2Qc5WykIONkZYWQshMzMagas2FdqDOhrtO2TWOzw6B3HAAVyXLrHsYh
ANUZIQ3rzZp0tlAqvFjaaZhRUOSVrHtnpMTcb1LVhd3MZ4iC1HY6S4jJfrpdwsMP
N08ccph3bjTbKC/Tw3AtPVeZhzUFkAT+1EOuQcUDZoQM4btYDSjsv76F0ABkau9/
nyodM57zoTUr0lxbiklGrmAvY+dxWriHJd3AQLthKwrofyRFiBZUi7sxSKNaXZrk
2JbpO7V20wMm9GNiXoNZQWJIUEh4BKBq66ye5fNRRVlAk5q7IQgOhdGcjhbbhUPn
9DackoaarWM+5uoNXZjOmlV/9uPv7AMzsH751GWHlyxFiMV17/+bf14WeU7gCkbS
VdZ/r8l7dOjqI1NSDJTj0Hkg711I7A+MqP95BhdErGVRZP0BsFkp6u3U1IXsOdnP
EqzszUC6htD0zArZ99Qs4zhKXwFRHGOPJPjUMQm+skQ4TifqGcPEtwE2bFtLsUKW
03SyhJXdcWxW7U6veaHnZA6YViku5cHmEq11Injb7FCvSpMP5ASFjx0PNPn5dS+Y
Sy4MDelfw2XceXjBwHa1yMeHL26s7aIsTB1RRxto5dUbejNPkOdSLvWW46qO6Wyz
A2EyKcx8fmcOjQQ6BYvxejVe93X4SU5Jk6HCckDcpmtl0JjW810nni8upwfy6gSK
tnyzl/9H6rBnxKeCFU3oVm0V8eR5y1eeFEYpGCAN0Kpr62j81Z3cJyV90uSCaFgW
XycUFVkGInhC5qVDpTxo8DYOgI7lYejR/5p7cXaqLHQWauJ4YBDPXcEgWuc5bKU5
DXapYHuIkmx0umMjAcrMzs9durtU+5KdcApi3wtPQYpkPCmpco0mpTRDqej/5oP1
QRSse/6rXyNqwraVlkAqHhPyWSWPyVPT9vuom4FTR2WJJ7NJd44rokg1SPaMnq6H
DQfxneFLLg8S+7UOaQ4f8agx1dfvDLv87/gWOquZsZl/W62I6OR8s1QPGMSf/BW+
2VqIgDpkhKwvqoR6TSPmA2wUItzhCWaODYZjg+D66AevZCC+b9d3w7KCnQv7DMaK
HFBIsNITQ3yvd4pmIkgqaVUn3WnmBXUxnbPPUT7/JIcI+WsaZv2OStZYcyPbFV6v
PVMC6/1pWAp8H3LVv23FwCOs+VCF21wc8Q7TfRso3RU0vbXqbKuKW9QWc99ILudD
RZXrZKV/iyKMPyRqiwoX3W7wQfMTgeB/x4jBrJowXD06wQrCxY13jc1dm3Csky3W
oOzfxKjvy/k+uUmpat1fwgv51lPiaWmopFXHzOIOtvwaZm5JaZvSRlDYXGA9DwUS
Xot+ACirBwEAM9KY6C1tEbyHQN5PcsCDTOIPKGL8sIhxdkfQrMmKKcBLyZl0MvCr
/fP31VFsQSxxAsKzevQg8UTRz73r16O4aKImTP0zk4fe1fe2kAfDkJmK49YLssam
tzqX7nMEqktrd9o0drrvwnEAQkaJRi/F2ZxmboYJcAlIWMJL/KcCIcfJPlcgmyGO
PYsTu+oLBYt1NtjLETwyKFK1bleAJccxGgs1u3LVsYJYL6E0hZ7sjsETcm85s1Z+
EluPpMDCrZvPR0bRjEJUrXym6upxhj0cYI1NfzxsrLJvKXXvM6oSBw9s0tqPHBCu
8ptqcr2ty9kZ8BW7jZogUdQe4CLs1qQDAd6JjX/G/w5WkBbYsZUeZjY8Y8YZ+Ikh
D1FgQmGICjhJHc8pnDxfthVM1MOEfeO/HYdfL5pX34xOkrFutp42+SYnu3XkaNc6
/eNnoTmCQ+O/bSSmpx5mXMfPKE5sNgnL7Y3JjhZCezolBMvf0U9u8wEaPtlAuoxj
wFbzQ71P9aZ2bO+aj5oE7yOg0eekIEBr97+TFTEDU4awoq0Mp7HGV+zsJafPkyX2
PNMRQRo5XfKvPUSowPDZZkTzcyQin0/T4AHyt4Ir2zNaTSRPTWqZmSGpnP3xmshO
129cvF/QtpQj0lzKQjPDY+x1XZUiUJDifesg1bT6fkx2JtwgR+bccv7+T3wlY1xF
+eh7qBesrD2SvAC2xqDsqn1rz4DkK+NwYA0oHNMQlYwdIBulfoFw7vV3B1ua68Cy
sgFsY64oFGIkFkJGqV78mjRjXZC0MqkckU0JwBek2Y6AIICEWDz/4befwpYBvp8q
tbXQd2s48GdgyiT3ZxhPLIU91QCMGEjtiWXOFimJMRO7yy9Pcs46+dsTBQ+3zKUT
8gEQ1Yobq529TAlnsXDIrUOj+uW26aIQ5EWxfhqRU4Sv7A5G9irl6ViIJ2IyCl9t
kfQAx8A+lSXoFQ0+o9j2abyIQnF/8abiQr6fwdybx9IbCaZRzSo6cqlXNzyy+NU/
oGqflq+VUYi5+MC7vhPtYlHrdDo4h8WNnmDWiuq3gx9xaAfJVxu7rNLdTQfGZcvv
eyNrAX1mBq322PMc1agw8aeOxZqO71hTgLnjqIRSCTgx/bcwS7hZUUwnv59yVf6j
wI8Ri/uUklZqLb8NQI7SGX5DVoYAvj+R9oE02uZ7ck3VtsOGwQdl6pPuNc7xeGhY
WtZUAGncbuQOAgOgN8G1EbD7KcwB6K1Od0Pa1+iHl9eE7kxHHK8umxXFl+9KbeFv
fuyPK9kocEmdU6XRliF/td8HwRh2GO513i3hBFT4182wFKEbG2ltx0HpCkiGizao
Y0mJBhxcwomk7NcFdkW5Yed1ffAnxsXC+JTTF1eozJkXi+hpKsGI+O7eE3lCf3Ca
6PGSOyN+vo1/AlUm520pkz9TWJqwveL2wp/+m0HVryo+RjFiZNS6C1LczR7Gm9Rq
n9HgamCKeWWQ7MOtyOHOKlFWMafjPzeeE5l7JHPeFRIgpRa64aBDnUyfnzzLeaM+
EgX3AJS/9J+825zi/TBtR38128ok2XbOaNVq9Ub/MZ4l42oG0W/iRjVliwrV0w9H
DHQEBdwcd7LIenp25hqyM4A5NcNKUGmXpzvi/HOOM+vEf9hWD+74cva+hP2tJvQn
DV1z139C0yECZo/I1slqs07HT6qza/CUb81b7VMET5CvCMBmUf2Jky9r0MjaTatm
b2PguJKzkaVSlWHI5sQofoZOqjNYrYAn+dN3xF6Y8h07OoNE4zkalz8hqoRljzJU
q5rye7aU+gWdgLVQByRNACjkRWHLgKXJEOSus5Z144pULsKh95UWemHg07ry2gJO
GKtAqRi7nZTYjfvuLzSNJl4MyUgILF2jVYiyRUp5Dc4kBavBTPmMSzyR2/qo0i7D
cBfBPAevvRQPNPnSAivnIATMOyMNAxiBSBZEwv5g/qXc7oOlTWRUFbsAzihBLBkm
F8EV/5XOJCxb6p2PKirgVmPoxeZYKbi4T9yebDc1W9YXhG1dKZQmZA0DQO0qpkXZ
rx+cg8n8lSHE/NQIPZH+CBr3j/k7qn23FPWyDlonMGAvoOZWZNc95C4xs7q0nMMX
zsK+2Vrwx3/a2+2gx7PlRFk0ZF/9B/CJBnKHsU3hoJ5elN6rfR59NvDe0KY5XiuX
+J1VEr/voiazcgayZWWafuYgRhJC/XdAwapFyeT6aHUdYoBJF9mLn6nOUKYrQl0a
7WH+iQlqencOWzxKtEry5QoTl64Hfozw2pIBBKv6gqJ0B+4rnv8dUAm/hi+GDPeW
D+WTbAQSpSj1AK5UEN+wU5Q5LCohvm6IYuNjce5IimQb1/4nT+1yA94Qft4yBKR6
eAsCZMN5BhnLE6ZLaRAwLn3lwP/W7NGkZ8Da/+LpWTU8jzEzYxSoezS/zlgAddzB
UvtFkrJ45d2JPSxotch3wALHtGlGZFy/0flT54cJh1tFQgor5/rfbMVHFfdYsGCm
EBb4a5IOqIITLbeYjxSDhjUKqQCEkdhut8JQcahks9fsQSeFWs66gMK7CmXUCqnf
BfQgVLSiRf4hSC/tZMhq6YB0qoODf5v1GVGal6CFNCaU7NFJIMK9yA0XMAPYIYmA
wHehBO4/MUfFm+/xZxd6sNzKodU58jeEr0yrMJBvvmoEbKKAdupjmUoCXUX2sd9F
o0OK6+AH5zTsqZQH5SUQ8JrIFESnBCheXeQgD7YOdktP0F+0o1P4hdJ+2MXjcD4K
vQ5qiQK31jrVzRLmnARk1EMohuSasWTEhlBdkylVT+ZcBDlpxQ2YMvR7q/cohpiM
ncGB0Di9EFxiz8/rb1WWrqlUmpiLobLI28ghj5RYZ83rpe7pwOvheAyUVIsAEFIu
5x+gBo8KujAdEfLOOf+2OP1RNlsXuakPAy9H3FCMeiRDZiqVzloVTKplHM18k603
4HdGALNv4mu+ov9BpceFmMlAhe18jZCnpf+6ehUzpZCNiPLPqv9/QvlWCBLwJLIP
+mjfFXY9dAjrnLylsQSr2tICrBQMyY8gyolUdp9SH3O79StgF2sUZmgRXDI68ZK3
m10v33LS9FGMYLWcNKbKFKhki/hO9lSelkVwSYITA8oqGsQ7f/761pf0wkn1g6bi
/74MrztAMcXjtxptbhIH6q3fjsC4ufNY0d2R1apPyKzcw/Y5bi4kU6RsMciKRvDb
AaPUfHstdP+XtRvMLiYIbGfAPSo7ZvfnWRjcmczdp/9xc3PfxFrSTJ3N9pE85zBU
RbDyMLrAV1l+GTlwld5+hqlb2eJQGe/QANMTk8NWrs3nfIkUapzATkTtZo4mpt17
XrekMLAecJ26IzuNTARGMF/ee2EAagvwEpGmuFBv8D9Geae+0nlTSEFIT4BIO6y3
QYgarmfHZSGVn92n5UmM2+Ewcdv2moYTBdt+Sf+nXKpeaus79x1nWdomma34cIza
IHhunlQP0PQBPi8BBfRhJEAwnpPi+13OaSHKCINdmG2VQDuIUr+DcsAJfRAVIJAv
1gyR8q1k8kcwpkxqyu9jvGDQp6HVH0rpGy250ag/8lge/+V18H1CexixJmmJk+C9
xDygilix7+ifnYNlW7WLi3tjv5hBMY3jzh3d21FahQi8z1x2/2vKKRaIcKq+NRJH
CXK8kllEHwST/FFSQIe3lfxJw9Umo+uAY7WxgYWeIgRaodnk/0hpFS7aG85AnslJ
c6aFFpUxvLkOPHRdNK5xEgVR/4d/OfB8bcdeDD2O9zFbJVoKCaixlt8EdS1gwgGP
YWtfRND+GUePSrEZAQtHxYuNPP5ckJahhemUG1c9+oAowcn9UoK8YWYICE6E+4Wy
sA5RzbUclOwd5xgRMNVqA3oAiwfyKwRrlFIEUniUu/hmV2LwhX5Gjlywk61HBdAH
Kylx4OCYtLZvvjPOS1wunNFx3PbTi3FFFPBU4KQrO4MdNoeF8Wikq3MfYNC22ENZ
neVraDxavJXL6ANH/DkW6CFPHxlrDI7+xN2o4XjK4wfXXzHFC+a79Wc8ztOvTTQU
XhzpcHFjZUj9r8AnI3QjcVja07uCKpA/zSA1iSUYVwTNGKMGnDPhJ42zxxb50see
a5Qz0P9RDz1wvQFY49P43OjnOA9sEhwjeQFRNZ+C2vshI5NVpmSx7Zq63+lmcZof
5E0cdj9XXWw7y5JyHpmx38lLVBXlG7Xa15F6MimO2jgsthaFStn7m9S7D/yM615u
au6/A2LfH8r3bqIF4Dfzm6UlP358sswjCMnQL6BoMQSiwS3S/35KEbWxVpI9hM+C
H4Y3qrmEIfRm9xeS5Y71UFmKLky5F2NFs67zwkN9/TU9gDbTjjkyXBcgS343yJdx
gOGvvcbkx8VSwit1LIFD9/bqNMdQD4ZqjnYGjjwXB1WAouFCLRXXNi4PArDx5rqD
7O2Qr28u9qXld1Eq/IKVxWYweECfw+iIBl4fqmZ2vSvH+t6UDomNeaBG2RZ/I0bP
Xm6T0QWAp6r1uIy0N70/gmTtklJmyVOrbzAhVut7trMrsOqN7jxxHRk9ZDZ2X3Mo
Gk/ot1frPpBu1SrAzu3nyokbKyRvEA2biTnKoI6K4+neZfJPCpFVQ9VRIxVuR/S5
EDIqbBDYUvNCRUjmEr3SEX5IOdRvBDbgHHzsydGYwIIciXfXIhAcyHYKu9FgRX4L
pBy++v5ZF0SV823kGtBFCjr8J8wLJke1meThh/0pG10apc9aGvBJs9LwUaFZXeg3
c5nBWQQCrVhkUXYGN/SYb+gmj9Z3sQL/O91fiTRu8vbmgAYqLyry5+sLHrEaCzkf
PERgUzyC6t0oanEJFXA0MeQZIOPnwaDBJqy1N/rRjLkHuN9ZpXc0240EnJvmNdDU
pmBHBnb8BiXrvAYGDoWYCiMa7Mc/1p062QaB9nUfzOBuUcGJQ3b0mhYFVMlr02iW
3Ec4ORIV0F6GZtKWvkC7V+SryEHx2NDlV+l8H5bBVTIRs50J8D7R1rnZc+U3WeJH
EILww0cFsVUm3kiFzuYVB6330WkawuiC6r88P87uY1Ni9dSnHylDb5dBp6IdK6JS
KzuD0G9TdMyKOAJfPa7pNF14m8SnfRNrbuZBwi7JiiUkLoo+cHYheX7B9SRLfiBJ
SfN6gWwFMK6No/BEduNGhrJC2GX4fpaFyFmQY6UEQwF7ikOn2VrteqdsL0K3QCe5
ibaFcK8zBm94DGIE94/uzOI+77eaa8GAwDo+VKsW7Fm6B2bRNcBNqUG9eGommjzX
AQwuuiNMXffPHHTb22miaxzl2gMe6Mf6Xq+/gExVeMmtANBBntwLvW69PIvPqVZX
vuyGSTRTudsXaH76a//e7c5gw+a5gYo9uaax8En7JDoWp1A/CcWj+Bk8KqQGuZvL
lX/OLI5bQZvlqfGSlzmAPa9mboc5Ima/25LCvYFV4UfkBcotk1WPdrT8QUmQOf45
HdoxvCS9McaxfiRb+jVlQUgHCI/bGPyyjdAuytyV3FazrHyNLlgrIN3z9w4dY579
cvhQtegllHW5REME7tdooAHh1gl5HbvsimYn/33muVhqumPgLCcOlqC61Kfz3ljD
9IWgLq4GMMub1AkdmO/jpxkVnl6oy++Ats/3tXpmo03mwEZRGGDPW4VKe1sF3XGZ
gK4WFLBJycjhqGdaGYJL9Lr14q1hiTYP1MrToJ0nf1cxoK8peFS+iWceTHi+RYcQ
rsrTYTqojniOrCdtD9lOkXzP8qojDV3S/FcVN6EGKKhBf9YrXjSgTV6N5Y7cQgU8
EoxcB91e4oP6sjTNOLPPiBSgSmm8QtliExW8CIqaoVISK6w5JTfVXv2usHy9H6a0
UMvD7QKfV3aKaIdsLd7iDQkw1vbSbyvMB176d1FWvDGK8CaQL8mOm8/8+9R1KvEv
eXa0nodJTdZxfeYveG+CBwV40td7TtgdN8q3ZYCRk7iy/ARoIRucPs3PTO9ruIrm
6Bhy/6U72dSZdypDpuTor4eqGZK3Nrq3shz0FpB0Eh5tmen56P54qXBKW/p82jvg
0g8g4b6WcAPvtacRpPxdP7N1f4EUw8mmosWgc9UdoTiR5rr2XwdvDxeRagS1ZlhR
hdxfHmiDp91qZZ2SNALOGPWRFbLcqPqXQPPXTbFJ3js=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ZK+Gm0FnyNTX/qiNgUs/WntBdmMRtFIkUcV2J7Wwage0wpCMacAQbRb9JIVLzaEL
PAUAH4QE/kQYyUvWrw1j+4WmGfAY+2zB1CL0l51MaL5lH8xn1ETQcbG/oFnpoN08
gD8kPnU57vtjQgBJEOWtIYqxCZAwwrC3AUYGmkWRYxr7OKkN78KZW6eH/+AWF5a2
W54o6t6uHSC2AyrEWHX+01+MshObUkKyM4c2Chi7JyZUdkefyKXq/BZR5Gnzir7w
ksUkxDzgfCRyYBieYwtUajadznaZrraPyFN3acTopeNvtF/RqDhjC/fuGy6Z4HFQ
8jq9PhYk/Mqg/LFzAOD7Aw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15408 )
`pragma protect data_block
BsYDaoqrunnmu2lUJxDq1VH127TCwMQExpLYzgsrn/MLRgJS+PNPoxG3dq3qS5oC
BIyUhOOnsCLr3Rasex9yPL9QKaJ9ObeoEbi5py5DeLdjZpCz7HM1peiGnx/foaXL
YgHGDGWGyRvpGTqr9gu+HPlP9L0R2ug2t2mvYfrZuqEosWmVAF0za+g6q3c72A5q
HjDvjlpl0/wwaeHzNtr/sJd6JYCGTvq3MzEJO+5EYm1T8lCIzFL//Ij/s/LkAFu2
FkL+N+200nWDjKZuB4onXRtMSLT2Kc0Aq1xQRlL2NrXSSey5Pc8b/cFPmd4rPXXG
++pZoqjq89B3uzs7D5OdRpxa49lCEu0zaWbXB3fknOkflkupclfau3Iir2gg/YyM
ZjpSf09ZXT+8wB8M8DbhT8ZzoxXHJES+tDcJRD8n9WuiKAm86kZ5ZmwMZigTtvYo
D/ID8ixA6FTMD6Z+OjArdoStPNZjKrljoDUIOSatyrwFLXTSZgKiKxrxw0XVWkEG
bQs5URXNfVWIRei8U4uu1xPDz9+DIKO6FaoJpBTe8UgEgs8+IJFUzpqNrpek3iT1
p0KnhMkmYkpyQiiR+tppnsPgbrqVq4sWGoInyecs0nAqBVaAW9cfKu5XS/gZrC36
tYfv9G74GjPBmY/c6XohrYQ6PU31Nxez0ZaiWKMajNiniim2fS2DsBpHULlEo/xO
H6CS9HT/mA7byYc+f1zlMKvLLEbIW4fM4fxElBrlV7aw+FWTs8PHz1pvwWKjSH2R
sTsgtOKgKgobTC7hN6l4TBrV/elaVtMDhXGKTHBPQc1WNVew0pJCsLjXCTZcREV3
yGPbqph6stQYuUWDQcOpHMJL1/96ppl4Cg5CDYgPSYjqMumwtSDTZ6HbQHZYGtlP
8kK5+lriBtmqtlvIAMqdZsed7nR/ZhWTRY00tfmgphzL5A4jWr+oztoq9vic/ke/
AsdzHW/cSfhvot1jSEAUWL6NSL67yt87qvOAoBF0gaepc7kkLTWI6OV7gd0hCDAF
vc5XVX95wVxRF2Asc1qmoKEPJBKHltc1uF8mppuyCxg72L9f+yhXF17rm/I98mIN
SPiAsN5QNlFEfypKpRxa9DqA+mq/Czx2MC1b03Pxz5/Qj/xjVqGN+kW0IMrHbxB9
CFeO0lM++tqUSJE8OTlpySnqxEeU34CaKK6B12dZbqi/q3yiG3T1m1/9UOD8dQeX
mq4maXh9dgocUcG5Q4xA45liHJmuteavhTBXQkzYNaOg5iF8/1IYvSdFM0IIk1io
Bw7aXVB5AHfP8OdCy8LcghjN6mtZALX1MEDlmsJ8ZoG2tfTvwPd5eWsFlG07+ant
Q6EE0a3l5zCs4NBXJQC5s+FwZ35RgcvLjvBlipQbaBf9ggF7FL0j++qam5+1InXT
eVchcHENE0wZuPv0EDIiWRtNMfficPRcnRobxiU/XF7TASH4VyAggU5EKeRJX4hu
wfMR3HVJPpKrqIj0zgDd35hwWDsEuGUwtLCS0TXDIDcfY66UhnvneOqta2e2ic3q
04Gsnc70l69aYsR9HTyPL3B13DqwGgtYuC6BCTRSalMehU5dLolhVCqOlQvfzi/p
Hwr1E7B/Fq09tWbx76ywGPds4qHSGd3HmNGQYxSBMfS+2H36q2qpiLe4SoL9vl7i
ByhreFvs20jsEku7s9fJ0qbHNxD/kBFJmwY47w8UVlXX0n+dko3xTpenVRYkB1n6
g4iNVNDDF9mS1oOtJ+dtWUcMFVFVQccZ9hfr9TXP2WJKtTADYUON03QgzR0oOFcp
PhtPjP0e/WcSEikOLKDD6OFmB8AJJSseOejr1jX2rqws7NiiU0QHgBZ+MTe14V9m
0/NA3OSSDYvJQI3KLNAvjpRn+0eCLmYKad/bBEhz7PMwWuWpFcRjqXHcjcsrMvMy
+oyw5DLEy+OCbslxtAZxS+4tyMpTgCl5/a/BajcQMjZZNNdhcj836epNYrrTUnwJ
JbnOjqv4wP1+DuZjcpyHoFUFHso3gvuoRRE/U2XPrNKaI0pPmCXLnIkS+eXiga04
bWeWHNP9y/3Z7+ccT73wePFN53XdOgq5OcnMgWsoBf8NDiAslahTQqCi5rLDcz8T
VfB6IK5gp7Bo13DbHZdxXDY8YuNNj9eK/iEiDrzIwOHNRRFjW1lFdGPUXxobpsVR
v2guViWGFl0Mmzx9hN+0B3FJ4e3EyOnFxhhkLVVrA848cdwrdefdcJnSGcYa+XqI
8CiXeOWKjppCmBtICmTQAtfaxgXIqIBsDdF8iznc/ntRu2I5pm1Y0/1A2uhkypK3
01Lfc749Jbly3Sq1P7L2xo80Jll9lTbjyVtuV8Ug14RMlMmI86ZtEnnHCjnUMtle
tNwsduIVyHh1K5x1PX+Y79ZuOXCuB24BQlS3r+B5fXbWsncUn/RKQDvMB+XCR9Vt
jQUJbjHICMhQlupAHXn6KJ6Hmb7cAGEvoE9VL3ua9dd5I6FSAMw1vofuqVZCEhmB
RgWejzSVB0UNQH06FtA7gIYFYi6uWcsEFB3/0ACM/wyOXJzTRy4Xgr5wniti/d0D
eHNyvAY+OAQoPDB1KUu5AayHc/OLljeDbYwKsS1c96eKAnssawa75VWeVlwTe3fW
b4XAaGOvWMWtwofuTolOObzJvwLPMg0PW6pQLLGiqWuc8iEzOG68c4KDUFatPKl4
UxqAGcZDbrfhmPTjLm5UbXW3vpyT3dxoUBv0mbb+mghkpFjkF/vJRuTBM0GhJLV2
FnhuI8ZdL79GRVbpkHuE0AHtbjELTJi3FwYRMo6Bc5PNJcohP5SLHkSXdGC25F7z
E1Xi7G1hKr2149lRTQoDjE6TwtvtJxikN5tQNXj5p2EpDNLE3ke47QJJPsnHaLOc
3etx+c/BnlMMbiwXMTTy6B8Il9UzKZMPYOtUfBpOyuAFL6vT8U8crksTSC0WUSrp
eQDwGkx7buJxQjDCMt6CcdUY0VP7pag9iIW/piVaKc+vU7ufs3mynyqXG6Un6HoI
2gN6mCkjIgTKomjEaCADF7zKYhu3KtCS0cqbiji2y8Ck9qRMxsl0H0PiBpkJtJuq
KYM3Mw5kHyYnqlQiSar/L9X8ej4Ytja6gvusUDESJ9oIg9elDXyaM7zFyUPlywuT
eeKWkVwvOgO0ImRSvn49FpoBfF/NxRu5gTbv7pKSs0mdFcoTInbw8MIOiXbu4tjY
9lOJqT68X2PifVEf33igQI8HjUf8J/7IAjSQFcAqL4HWjGrdnnXlMSsGmzq6jZm4
4iNBIcoEiImcBlk/NopLEUx8B/zRKVhxs2egT0zUnNJKmTqzZvVwnt7ufNuij2en
c0G6Y9vElBa+i3PZqFwPODmDhjvY8unqe5eNv/wgvLjbQSIGndk5aJSE+gBrjbsb
au20GhSWf+aAug4vPK7DrbtVnLmkf203Ef6/Jayj66PSNTeI+11TmjkF7lwYZ2iB
SyocnZPVEEJWVFRL7NrHn9hhmi9DX6muDomEY0imXSaGCa5ESu/S6kNycL7OGPCQ
eXSNxUO8v5QvQxVJlWwP2N6OsQm8eYY7BDDd9z4TjPZYGy/BS3mEAra3PUzKMBX/
wvYEgdRohNQ8nAk2HH9u/M9WERtqdXlxoeRwlN8J4G+dbS1R/gIMUJn3b2krzENv
wcMgPvFK89yoSWIa6opLSldz63ejLOLO4mMpd5l8fOW1vKX2kWBz0CGJ2lr/U5ka
dClX8h5U2qRtn4hsKdA+e1+DHgb/OdJuB2z848JuD/2gZM6urLjpfKCzeZbIk1QT
HYLvtneimQ3xqV65FCB28ZwDW3IA0e+z3QIkfPAWDgfscYbCz0UvdfX1y1E8gmQg
CN+aRkF90J448IRMk2oqWjNU4khdIQgRF42L2cFHfiUDGqDh9LkMMs8CQ36XRiHP
dXnbeDGopGqKmoXZ+UXqBt1j7By/YAW/O+T1J9jAs0DcDXnZHoEy88vK0rNpGaAw
auxEPQ4Ct1L5dgTG3aIQ4DZc4+VVXYYJ2eCfZVpk23FSehGo/g4nCE9UKqLd4Ejw
4H+Zl9tOvsL/ecba5unZEY3aAuDe0Qr0pQ8yN29tLEMnIoi8+8W0jztJYH4L7wUQ
YdoG3fnO1V47X5nIQ2M2WCtRkRKM20b2uQGLBeQWDwBL1dP8OpHkNAjQunB41UaL
CVugsiYt6WlL0lrTe7yzLwNAV/VMUnptyt8exuipbyXQEMvWTHOxYKEHhUgQ6ZfH
FpaSRCYPOattxF/laxA2bYo0Ky7o/eWfhWBGE3CxvGYgBpluBMkfR+sqq6qZOowL
VArIrt2cj2bA2rL4oZDczfw8b69XStlaTaiq2iqGY3yiRm/K5lpejlU05Dc6xISX
ZSNT4+Kn0L51lBEHdkK2Kd+UAsK7JAQO2EytQgTYhCkrvayjBKxhC7NP/56o2hKK
O8H/5TRxhmI1E91XunZ+tW5o4udSYJ+TJkNSghacs+nGNybnGAyepEJclYAU/qTQ
N4nQmss7wd7/r4ZBqDkZfsjgPOFOTkuWKhbvuQ5CKcQSXKoQvp1jdCITl/Le9AqQ
+FutQzVJbUITahaY4TYsSulWwHDXsFLAttx/YPN5VLnk2Oad4Wa1I4Q8fPkyRk2a
5mWHMgFskmKp+uhSG2mTXTBtySgXlNqx18WR4lD6dI/JmKsCc8A72d+1xy78j+CY
9t3KStR38OLM4o3OLGycZi+l3XgNtOXRq6d4nkkLn9TSFRlRGGvclgnTwWaTLTYB
xVtJrM/MePw1iN+N9x+3tmjQXm642HFUdJ2VtPx35drYL7dH4lD/PWGc5+gCH5Qs
Q1FpfL/RUGkkfWOwqwnhhLtpDqflbUCVvZplJcXDgZB0SkLrGexJc16rZBx3qb9z
whxdvWt5Q2w0Bjnxueg2/p5XVDXudSk8a+Go2ieqTIW5YoDkgtxLY3rX72q5YR5R
bBJKYg3hDUBKg51oV1iLtx9mzYksVN5Ith76Oa5dZLN18M3VIlPiw2TGJrK7rssW
kxQukV541QqnCWa8Wg77fvfq/jcMvYYm9bu1bOtlmjKYqfNjhk4eYgs1qxQpVQyT
3hAueO/MxQKInUfmkWnp1znGCsDWPY0Uj7NewDshhne0Dv8slIXbDqKLIGdR1l7A
iCXJttz7uPysnml9cxIXzfaUwiF0U1ejHPWBy4yNnesTtLMVlOr0bQSdl8rskX6w
uma9sPCYItLhJc8CMkjgKW0q0B3gyB/002PN4naVBfoCqlBd3H/cvTni/SKZ2yh5
L0uQDQPQ6NrXvQdtgW9AVfjbhdYTCBFngcflTDdJH8iyJAn2S1Gst+cUzZxIQYMU
pSDWX1nStFrFaaz+UWQUy0yFeVtP4vTF70t+QwAVqvpp3bkUOwTdZB2a0Y1EOL5w
e/TsWilWjbx92HtmWhVDra2XCASGYzhKfQ+078COpXd4CK6KYayu1WNtODQT/BUY
FXt1uw2vJ8Of4SIMKCIqm2pkyE07ruoqTjiHDzQMOPV7zEQ5qujI96WuSsd3Rcn/
PJb5Gd259D/LynwnjZwQm+7Y3ZTonciLhCXWT5RHKeSwutjZ7g/SiGq0QTjQaTyg
bAtFu/1cmNtq14SkWbwNIlXsja9zXUzQYER1APwiH2j6jR660QEEVnLMGjgdOowf
9B1C2spo6WB0kBrXMLC3ZBpDKM9fNDigJm5GM16hwmOchCn8l/0ia/NC22LR0JGe
QfEU6oKpWgyFrBuoFD9rZcM1cTmpsHra5hqDwdYEOlCq+s3061qxy/HiMaieG87G
0GV6YSwYoGmeMJvp8LUDbEIGGa/xige33oKOf/BrILnd681RJdmQXHHz8WfeEOR2
g3N3bITB6MFTfT//CqUBypAzuvVoBIFKcxUGne0vJ6zQgKXIezCwVyU0ZQJPDv8s
eoleRo6Jdh7iQ6TOVqcYhDbBxUNrE5AhdSrOPCovb34ng35jzQlYf8Y1m1RdEZV7
/Gew/Y6pdQYh4tUBHpIFET2zrD13W0qUN//K1xVjLYFcwKBWxYg44j3i/YDhn0QD
HE8q65DIccw+Hua1gPy5HuANjZGXI5aD4lmhFuCiM+OwjC5m7FUBy3/GJ0EA4v6S
fbyAPjjq36lLhpc5FZY5COHg/Hgx2TwkuWO87eae5rAw0xdmTMF7UPTBtQRWmTb/
/7X5XpbUG39ryXLp/U73AVzXUZNwDA4/p8PttwbsR/f0CrLqvgqYWjT+jI+cxj61
qojge2V+/hvWaGx5KTabitda2v/6mk6r2zf1LvFE/vPzXMBMdEStufmnOzWUJi1N
MZi1mMG1N5nweoEEjYCh+71WUaWRSvkZ91I1gawnizm7MK1fTqGhtgjU9RMyoMNL
SZENu87843Qb9L3b/X6xD+eYwhDmHV8DPD+YDnv5qgVAUt53PNC1AJ0LRgwX0aU3
YhZiowlz6yPbLycTPvP+xO1XgWYu+KMdek4wTOywLfe/pBPMKc11S+mxRXEfi8pV
0vlU64zCJfQ5ecxXtTx0nWeH9nIXP1fpuZ1cN5sKE9RrTLEhQbBC19VLM1E6204c
Nr3dux5CsUEVbWgxR6n3O18qHaTZ2jsHuYaLc/dYW6WL20XqQMeQ2mmiITr8VNE4
GtpOK+fW+QgCPA4UEsA1ut0XBJHi3zb40ocbPlTtZ58KjwdVAMmNnxkehZdo6dWK
ovoqVoRBYkY3smyYZcXgvapFau21jxUhX/et2rGUDoKWXbchMoJilaSFR42i9xnH
M85GepmkATj2YDqk0X+yb8vq3haI9VgPXG9yHhCRGtnW/GtqIADvGWgBqaIxulL9
XzsFBFCe3TMK/J+m3QCk8Z5yjdut215IXp0FUq4HTDQbQdfZmhLamR6L9iIXWJgz
KRKUsywU3NS48Dp6JfNg9IBvwybIV67hvFhtPIJifuQyMD2nzOI2z23ODxoQjEXa
UqlMeArF05Q158Ac19ltaw7ID81xIaMql0mDY0Me1LjyjmBorybD76r3E2Gp1qcO
LSVOXaW5Cq1Bd1nCJtoSr5xk+mo1kvNKf1JWPfvoRmETuQ75oHkxmIU1jXo4sBW8
zMndwN8467Z6p6HeKfZVnT4ghfVNB4iMvqZIhvWxeCgLkVpwyVW1E9PHuw4C7thi
9M2jAVGMfMRJpejJMLCmheRjh0NBSTsPyCeLTaLTfxD6KebwQ3lEej34i5y7nCyI
58Da2blQgL8evA+10EqFVlaRGyPdryXGBAgGnc68ZMJlR9YEuNS2rHvArtnRQ/h/
bQuyDLbvAsouiOK9kDR9Q+KhaP8xycHZv+Gcb6kCPePiVu9fB0b8e2KpSN6H09cz
Fch05kPerl7uv5n8eXI4XvKSkf3X4Qe04UGXt9bbyXlH4GcDI5umHqAnlocvOhK2
zgNBunjyuk1LhJsmv+rMMkbwTot4T9Uyb4xieIxcSbM3dcG31lKIFiufQEFj3iGy
7uAQ5TaW9qsjXbc/O+JHOt+GCgH5IpUIsCkIbyyJnKlkcMtJjR3aWihGvoy2vyEl
8tZPQNYU6zkT8ukKf1+mhfrk8EVGQJLlFKemGEDW4Wnc2BfD2UvOD9ldDDpFFHkF
XujiTrKxSRzLmX18tjGjwQLlbRAbHD2zkmhQHHFfL1Ocp2f3xMnKhjRgFVHRUrW8
JAAIuCYkpHsLOSe7pueIFGiwamjPLWx896pppwkZ3oX2Sj+TCOvtEKSH8egxp91m
ch09VhPUz4zPjewoeWj1H77llNAMy3lt8XgQwEwLkwdj/Pf3TuWhkMn+dPGqaHG6
GRjAWly4UBcujO339ZuqYEbIh6dNrlBu7SnL3+QH7+W04OUIODJPXJ4yqqQN/Epm
HMcr6476VNMH+nqo/llkBgpSs+VMEpHvdr+CCKUvWr2iqup77gxBHUBm78XQHRXx
grYTAuWyBNbTNO+emWHwASERegndFnA6iW3F94zqduPr/cL5KZzC1mvPmogSPCJL
+d/mLvB2siUA1sq2Im9yjU/ptDpxJhREnHJmRNM5wIMFpZTRiNSXYmoUoGL6/i6S
GywTRyV84Y2MaWs9/kaTYvv/yYZ9N5vOZ0y3JUCcOH8i3ErRLiJvTDlIUNDt5wgz
MAv1ff+XNPNh2pwjkJUdKo4iLCsF3DwVfwP2nEND4V+njxFcT76sZqlCdhz5VAZ2
i5Doehe1ez2VLShmotLyEdgTnuFMOR0uOhsUd0jfL5m2olYRO7/QYWWNE1DKX+tF
UEav0CS1rRlKA9fjKwW810XDYr4VBw0C8jHpThqvDPA/9Q3X9jO7hhBZQ+ghrJFL
cfgyObAQ9H9Iqsr/B8EM5SDgjrL0Tb3MXHXepx5eNj+p17i8wUpl1PkSbH3DssFY
gICPb8ZNqqKFxBpe4O7pP8lQ/dz7Bk1tXT8kywH1bhN79mrXgWf4EwMRuvfBPaYt
AQ97IyLFXDB2X9UfpyWnrwdre+0ebtQv72gryL8BqN9Ab2jLXZsLOSqHNz10UotI
A2VSEaSJLCmZ2gb+ak0AaMOCUCGwZUyLYnqN+f48WFS8ef7bQSC4I9WRnNG6qcIy
03aU4Yz8IIZjx44bj/fRC4zVGstjymb4xBY099s8mzZXzFtRd4dI+WwXtuqISnws
YNi+xcjvlb3telE15qdVArTsAbUqgB2ZPnKxUYRyuErHm7dD7kgY6PIWIx7AUNuN
CU8cns1vkJf91ZkJadZ/SuTN9LzgoO6CNwxYREGcjSaER28mW/BZwegfCoKyNk3K
tl4npczfK2tvEXgNunW5eS2Juu/L06+uU8kjF5vvT1wSOZxIcVCplaY3+1pGJUbj
14HLN3UZmiwHDjsxFlywR5aLMavsvc+EMp2nMMumqIpapkSCw6oBnOfl39nCW80c
OQeu1Iof4K3yzdb1k2NXM58YRNR8ilH51c4c4DR6THGWw8KcM6LUFs4hhWj94c0H
1QSeiI2D1IUEFH4x4VvqHG6+8wiRbbpgGIu1jHkFByTya23WX4vJPYsYW4X1y16N
+4CfmoLVbqpvTRfozmR6XflFAZgxKkpWpliZ2TBXXyIZTaluMO+TSs53Tnxa7aa+
tgfTmg3kMc+xX31lDzvy4lhe1wRTGJfUJqvpjno4RwL1rebySDF299gPVmaFE42m
yBAF5JyxNLNmOoVat8vofvUBvixLbESpQbakzdQyWgV0sXoQCJYp0txD8GIpOug5
a9LEuPwPnuIhX1FhHoSafKcf/AVIw8A06Jy1MrOnC5nizmzCWniUa0MlSxdIU1rJ
ex+CapxB9MNzILmN/WGNTfSEduSrCeHtHhftoSONX3mg+ntdXCSUXYNSpxU8H4VS
Xm9Y5v1oOYDWT061rGXtc62fDx/zoPt0ZmTtfY8j/L4rRsAg70Z7ubig+Q0wXwhU
w9IYFFthhcVfmgu4jIS9hLwaTaeorDlr/gZyUF3v3BcHWgO5NADYUnKceQ3wK5YM
3sxB8GOedNeyFapH+v3FzMq3KIVd6b69Szxnc4h6vswOFsKe0jbVL1Un++Hr7gZA
AULotdu42E+HY9ZDS+GwCwwd9D6RmZX74HOtuJgILZNJAkJACtoDGGE03k/4lt8X
HBUEl7tRsGE18cG75fos7c7UZIgmO7oLTt38f0llnPW9ybXKmT/1NH88QTCmURDQ
aPq89JFgkT2ylM5mhMWQ2VaeYDztMglFcYthfRWVn5/YF+ubn3CdyA1n0I8xJwnL
YqdmsoNORUJDFyC5bwL9NkFflhMWSsjp50XdgOXoVlBcXLMReLYIQ5OxyJasN8Mo
kaZC2CZuS4DkEPWImE+ODRoUSsgpzUSv5pn5wXvrrO2KZ5XbeBjgl754pYRWWRi6
rAmJzIYWrWc2MSb7CFvvpBvn7UQ6WDVAKkfm+QJezQdHjG9TkjPoQfzNKnUsWj4v
5forzsVDVn634GFoUWg+kFGsJfryzRZ/AFPZg2yAdF5Pi/jEE+FSuAoi3k0N6EVe
ZL2RUlrkXS8g+HHu/q7GDumjwmdaMqqfk1ZmG95RslyWXvvnANnhVL6K509PcXui
RA7CX06xCLYZOJyGI+S3K/CbJPvc6lpNACQbo3sw4r+X00HhwTVE+jH0CM7f73Vi
xzQEMVuhD/T2rZGtYe9wVyHdl+ITTHXujtGPtveIt79jvNTWSscK89T0KKzkjfus
saZQrA0r9AxAo9NNukkUR6Q9af9CFdUDBGnePzoheAbvrj+UnFP3mtst7Gp+fzxV
3DGEXPYDg1QKWrwvael9Zk+C5Dc5SvkqwlV2d8p/e7jRWCSxRencLPq7dxcR0zbB
ycqt9tnKzfy9AITNsyzcfkRJnv41AWTleVwCoQScv5FV2DPaQBOUxiOJDC92OjoQ
sFiMDJN8yCtOEwjb3tRFniuDy2HnLVSO0/Sbp++sWLtOrx54Z4sxVcWJAdsS4vW4
lGD76XMvWFsNe7iWtRG1LylL57dee106/bpne+7DhXXl7m0iDtQKTxVtlPZSbBzq
UlfOWsB+PT5tLpwQpVBcPZ4fEBz1U2qKRmcK964hjg60z435NRTVml/Uc8kXrO4T
qiDEmjEMuXmGE6MReS7OExwlUmmfQryLiRl+iUFIsG63dPnd0nKUSuLp2x2Zrmbj
OoXSKIkznFBfZwn4rWROkCNL2kgi1pzqX9+rQslzYL1jvPfoC7tvFa1feQ/FdSVQ
aJvNNyXXUpTAyoH7NDeMk3kgxSJ1D1P4JrR9tr3Pica0dKw/tPm6wgd74cWdYU14
LNezupGwqRxO/9Pa0X4FoVBGX1IYvST0RCWHw7iK8owodU5PUhUO3e/Aq61HUfU0
+MMLJ3ceE9PmBZufXiTVo6OS19PsBhJI5Mc1He/yszLv3RQZLvzXD9xyqOJzG6jn
+0pOoFDCph/XkM/52zC9IN6OQLk8su+g4izQO2K3FyJz9H8NQWg5F1Nqu/DrkYye
v8Bq0Cm84gra/M8d9TLm6ZcPtUNEuSDnuF/aqqom0OjOFSzSCRZ810a4T4fH8waP
JSNqeRHj+l+29kuyDgI0Pox+JrMLwBkWQwHxmbo6ZK/9sxU82eM0fyGOSG5jdx6g
Bv9fqALsOYT720x8N7+sTNzsWvOrY6X5xwg9+n9H/38qfFGGFuyzHFOKuklFsAho
g/6N/SsVtwaH4vGUAU+X5dC7fLXxdfJlZEvqX7e5djDk1C/nyllWkPnOtLeseZEB
5RIylTtbYDhRfpAD5X5f1AQ1YVm7b9ttVJVFXCOvpIc4vGo7FGeqX5b4fMlk0Cff
q9h5nr2SlD31MUvwGfKSVG1B2j/jo+QCSncdZ7d79HNwHdStzUZ4eMgF2W6MiPMv
yTxvHUAoOnUWACbfeqQza+jfaKTwNtgLNIGgvv0cxkgIV0FkPV0zY4F/NhldD+k6
w/lB6nyG9QRUyqSRDvn+UK9NdlD+BhckAe+pnYc8BEMZG6AVwqQrANZ/MOSxAwZh
J6i7UQxseNiJwXAjphbzlA9dEyxtU7TNWnC8t89QUsh1v1FVLgLUrvmQ+v1Qq0np
Bm3T1RAaGdFgIqH7ZLFJXsA3cbZHgkB03tI1Tf/Q9gDYAfyoXJuidVHJqhctCuAm
GuwcV0ekpZIcBPXRIKzuu3embpHYsxuaI4KxqMgCk0YXDcJn5Bm1WGDqtiCtIyvh
hfW/MPRDQhr1TTeiX2hWea9RqLVj1EuRhNWtLMkIHiawECfDDU0bCIZGlGepx6wY
fYc49UsJfzqgIkbHjXowDq+x0q0M+fNW8v3JuOx9DTtleySMAWHLPd8Hz8Bs1Sd+
aabVbR7jWbtyqB3s2Z9skfejD1U9CC7hkAD7sehLTVeH5zOywp8KNdLYGsGDOq88
oUK1HgImFt63upzovDf1/bpZ7NuLsDa8k5EVLUfUmp/WLCmPgJIH8k1HKPHubm6B
Q31ohBXVrMvzcfONL1TJ0LoVvk1iHaIr3dvCxdGBDskFonWhpHXjggLqn7lc6mxO
uAC2AKWihhNkx2iGXsC0NVOy/+zxvoIPSXxlTDZ/6kjfKWyuSckV4jTs2mRC+gYc
M3zJ5MD9wDoqR4ykfMvMc9uU2nHEa5lrWhDpM2DSVYyyRc8gt49+z6627JC00Mqi
094eL3+1Gn3m6hdD3utj/ZrBYZn0Ebv3ZfL0zSXAacM66RAjg7mWkmqT8ps9sHqV
fULB18p8yr7yQSAfhsE5P0nasTTavvJtWKcMaBogGyGM8UZKSsDo5Uxs2WaSuyF8
uwV2Va5oCmiz78hSXiSqQISmUZI8lVq8zclLRfg7x6k43GUtt5ogOLyi4mF3ZltC
YK3mTNB3/CtQInyusDz95uCd9DdddeDBKF1mUchTB8Yr6nBnC8djKpoUoQF4gQdX
yeMdLFYRoGA4aAnh3okx36X7ge/aXgcmugDHpOl1dyASYVAUP25/xdUvkmoPXeiW
H6nZXkkD8FKFKGpIdsDBrp1gkVBvi7LTkVo4w0qVLpjNdezGHM0b/6aKtn/NSLMj
AU3DUwNVOfSfP0HTQct84OLwnXbesW3orTPTJ0JdCSS3mqLpkWZvOYrIiTPwVPfx
pwaIFWDo1CMAqYAmzAu15GctEvF1hdlrBG9SsNk8GWMrs3oc7N3fAnrhD7CkDvhY
GIyspAG35TqIs2egTaxIXpd7tRaX2CVIl2+rl3Wzm6Uba4NNN5ag6p0121CyhgUr
BZXcaoLf58+3nYX6rgHZJ0H7t7YkE0s5d2mlLHStyc6LDbLdPJ8dgDGJc3x+8SRm
ZChuC7NfwOPcAMNH+UUD8RPwBS2SPetUick7aEhm90ZkeccTuhcdx7WqlllI22Lg
ZmbAt6DccQMwJvuw278svbOjLiS/aNjENsLswGqVI0UOHehvN8eIopces9fkqGDT
dD236PVeyKGsCHePOebOmEYpo+o5Q9NsFF4jJIQGf61Akueg/9goH79FrI4P8/tt
5R916bsxPZGpnFBGBUoc4p6POIWJYgGxjMSKff5rgXbhNoiiYBNu65OWEfiDs+Hd
MyrUEXsdni/ys43vN5yFcV22EqkWJl+g+zc984JCemZrw6ZTov2uclII/ZTYXFfu
i2+4obIDvf1n9F69gOnzgi0+U7dIx01R3M42LiW6jBG4nxIjbrQopWs1tWW1MAid
TxpCZtquNi5sSJxECy71LQw65Ogyqv+2N+UUz2hSTF+rK0+FyRSUv9qSR813eulj
YrhZyLL8bect9BUytJAJivwvfOy785IIzgfqtDuRE/1Fmv+KAC54OBETI86cgiJb
J1rVqpnYbcNyoHQakT48CoLpqVuzdcG3eefdShuRnOwFBIT0qJZZ1fyQaBWnjFB0
MVE0AaTC0WGSBLCDDY02KCFtKDfVPUQKXC5lJ8hORg1c5s1QONGW6os6CvNTRPaQ
vS3h+Y/iK9Hz13Rm8PKWymqsXFW2knFDQaswHE5otEjdi4R4o8WfzbrZ26B4TJma
rqVVgDc03AcYnn0yAWGcRLmYHC+GEYtXTtfKTw0jJsqCvSYzY3D0TgXIXo1FLc08
YMmKN3sTP7ty0CNADnBh3jImlJRsorIxFiBdJWXMYfTToOXaXESy2Dkgbph2PmSB
jvmIqSZeGILsqIG+fIfFe20Mmfa9oz8vZTwnMORiuRY1xL7BF4v3w3jM3pOAenBo
WH0xYUVqfuGOh3v93ybe2LHbrohUkzfd4iHRSw2r1RnJfTFX90hthgJm/Pac+5T0
PyC57ANsrIKEB9LtFOH0v8F9dqavMYyO7z2qpurfjS2Siv+mDKFqTw0UlblVgHY3
H0vG1NZiurfytbnVBu+MhtlISGeGJU1AiGqDHv/KwCIVtI4TvUpNYr5xhehLFOCv
vYi7uIZuwNnGHbHwZoDWIzkxLv2oW73XjR1dfKLAhnBaEAjwzqTD+QfEvfj8EZCN
NMrgFcPzr1uRHDFYLrjLGSQ9D0kv0Wllk/2USNbzk/q3S38U80DCdKN/6lqWrzAA
Pryb8SssPNuxIM7uewnX83L1cSuHxKk1yyfpyzvkyBS+5h8jRZekZRYyhvZOYxbY
xXYjl4EGk/kH7txCcMTpcNUu+7GODf2DzhTVYjOa0M/a5Miutnm75kUgx/GmKkWz
ozNosrCx8R6ujbaQauvBvllPcN7qJkhT4hu9jIVfXMhYoEd3CLz8NLpsWzQe9tIM
DnBSSGkPVWyShQNBwhznrkioDdJPRSB+6KvvYTollY1UnsyBsvQNj3EEmguXfvyE
uU/pcfObhDt9mJtzJdGFdrLV8OWc39acsat5Ri0gCTKWaQP65QCLvN8f6SLufKVQ
Xl1D7vun5QdTFjEtp+4X9m4xIBmE5qoS60IBdQ+8BzvKFhvr7Huqu/M5I0ggKV4s
t10wMg/7T77e8M22MRq99tVeAl2i0CK17SQJPBK7lQ4AOei47NzxfaqVUl/4DbOa
Gx6Emfne0RCQFkIdxilaTZll+06po6df7RoigZkLDc+VaLIBfO17CLNf4drfBSWf
7uVBCbaQ91S80WUmxqXMcOdtlZ/m7KEVzSDv3dU4vLeKW6KVFDj39Wafr1XOBU7E
0cFupVRIQy1Fo/Z181P2uTH5egwNOItc2YpgSLFyAtw+xiVl6vUAe2N+nVtQGBT7
+EKi49zptmszGRxU7L6piNgdbA+1Ry9oUbdSP/38JU48HFUWn7vwJdAeBPpbo3DY
swV7J6mZSBU0GSF8Newxk9FRF5PcUKXPWAUehPsNH50GTZegSNHPVqgsz66iGKaN
AmTpdJ8hyJfGGnoIk3SOiOLQrAr2gX0v5qZVn9oC/ZofCbyNquYmNyQo7Axob9+K
w9z++DLMzrPv8EiMDC4iR3ySe1fKE4Rr5nQ2eG4iPRZJCIaddYtr9aC9kEy4jiKX
3Nu0G72IZcmOW9mBeCNLiBboTXddUkvFzhs5+ygExFzEGC20k8InvYgcbhkBZ19z
I3VJosGifHNbxTtWq2isx5BwP3fUbwNJ+mT9Wq8K76DhTAuABShHgCFF7gXqXvpF
kiV6iBXaO7kg29RZ3wHvwqSYPTGf1gmr2f0K1D59DIKOqwO4Pu198OYwwRl9ZT4m
FjCq7qEVYZabSuqHdBh1cj4koU0EOX/ybBY1AalurJGCXy3eARlATC/7W14bxuDI
Jr7UYe5Ye1lGOrOJNO5gw0EiT0ex6VN9tDi9BXfd8Z+S4ay3ynlX58Sr+IgFTzK0
Eksj2QFqz5tMiVXIyuuCXWde8eU3SrU2QZW2FyX7ICRP52o3/ycciM22ExKglX7t
DJbX6TQ+QRLjpSO1bdTMBZWpnkXLp5b0sxGMErHV/ENGH5kw4WsJYthGl9m+XyAN
BK8fw0kgtgHkU5PQQGl5cGm3dQyEnF61MWKWX/zLR+/ANUycSXBmy4NXDDIwysGd
Q0Gp12GU8ivIvR+q3uKqYXO6frihhMv6XN6TQIjvykxNJXyCDgND/eUQ63wmBye3
pd0WIu9G/I0Bq4k3naZpbZmJHGKCwyCCTLYkfpT8LzoEwUaOxWwf5lV4xzHBU25X
wBkga7FStI3vKOc3VS8rjh/JRHNosOoTPdE/Aau55p5FKi5Kj8sZApMSIg5mlk0s
U4D9XTDD1Ss0pcv7kZbi9iONHkSWjIZ/D4tb4v5iFnOQkIqkqah2suUlIhAOjT3c
H+xNdSEmeUfZ1sRqr4vWdxrZB+UkDxqyud41tNb5W0dnQEAEz0qVWVmtYIp9tSl1
tUPhSaOLy23N5VlvbMxy69f7vzx7u3J1UjM2ayuzNtJNDnRG0Ppv7lIGsOowUs/s
yJAv/8vEaVsAl213twO94y2a/45zgkKzPwGZJ3vZDOhvUDan9wySNbuMn+8vvli9
cCFcBE+zlO1EP6LFOIx5ybI4RFBHAe9lizZf+ITCvDhK9B/gOq4X50AxF/Bf9R14
TUJcHZBQ5Q1uhIqFPFtytmeEs/DzgI8rf6HOM2sABoXEB1zzcPLyjNQQFaZEGmoK
tQhxx0MjrsmJJLQeEHQ/wmf39U7Zc4gvi0oX0PkL/Zka5fdzMXUjl+Gh0ng2H2S5
RLhMfGvPL3+WrS7VYIYo4wus617AYUhhCGOx7d78r12C+ABMGwi9yXZ4nTQY01HD
tsIgU/Wdjs7jGMLF0zSDbKBCu6NzGe1aUtQXSsU4DsSPp/LFGycylFJ0VXUrhE6D
84LpglWMbHYPt3VnFRq61+LvLsvtFjl/ZFPT4iRRV6kw8IuTz5JRxtzsbGtlSb5T
dATnEG4BwTCGESebdGLrgJUgEmG4JOzfcnRtPq8xErTjkGqd4SGmcJGF7dcmZVX3
MuSmyjSAekrrA5XyloE7r+3t9l7wcuBod16DmkAN480xKbrhTACqjGf9r0FPFK5k
/ZuXh8rpNa9f1s001r3IQY6wAyWx7y7b5j60k8hBkpQ0fQIHQPKM8U4LqCYSmjzr
5EPTHpHv/Ks/Gfkmm4AQSw+yiBfnwM128wN6OhnPzI/FLWN/azhAaSQb/tLfKHmw
t92rj9QYj/RDP1exrI8mKq8a0cfdnSXx6THKfP4Pwg010P6o2NxMsfHDegiXPCcn
oqQ6nboQ9F0H89I9fvNeFy/d5Rx4RkvLxfwMqblFXh1fxH9X3hKG+GKUBAPCkD5O
Vk3RYfEt+Z+1W64bpjxkihU5MzQFEiEcyOZN2nKSkg9DnCS80VqBwJqsXkfthSLC
hCzlysjIjKIT9a/85La7u9AvokvMtX69kTUyZu7AVeRl3Gi//ETrUWQx3bMvdlB7
3GgJwStSownICOvyTafTcUTCH4GOh2vzGqB4AKHlkSQWoIdSiHg1RRelGwJQfWFO
RhWocMvr/JyFRdxw/Vz9U0GyUAnBIEP+aJez7NSYAHO3OX4pCaz5A8O8iDK5jH9Z
8EIEoDCSr2yk2DANk5RChjAWuFA1VHnwyehJG/WCMxKYSBroJQ3nRFwIfBEXzdeU
X7r7K2V3m+T2RGGtyHgOoTUMOygOESMLhtFhNIR5xaAyd12ERnQsqBH/8YHZZIzX
fVn2Hrq+IB1kEtUncuyhM6eI5Z/wiZZgkyKGK29R3QpjmdyzWdf6Shmp63OVKf1Q
TF/yqQFtitE2jJcHO4InfouQ25qllEdCgIvJ5ZHHU0bqpmaLZOPs1Z9xJOrk7Kba
1hD1D4hi0Dbmd7VjcuPaawWMcwXgzxxKj5VC1McmKuFPVoepYcMmUHq4IbqJSm1v
gfJ+olP0RaqoTBOskLwd2+CRevr6xC9WsS7IsqYLE+CT5GXkcqssMEvC5vauSO7H
Glxc4Sl6xaA8XXYzb88a+su501w3H47o/tm0SuEVr5sRLOV8xnlfkHNXvvWH/wo+
OyKfRUZvRy0RF71Uv7tSGQ/N6ObNi03I44rZjHboQpMFg4PcUM1Sn0bGFdLk9l7R
KLouV/LjdWve+ZObA8hPRtEdsazeiGhBowDxGYV3KVPOpHfXKIQAhbRgSUkE098B
lorWqtWV9xH63QEp0PH24H3tie3Rzr7Ijla+ukBvubnnhDPXetwRcPOAjO3CNfAC
lW/ahUc+jTlvKBrFUjOWPa4dzuIxKIV7LDwHq0nV9x1sblMYrZ8NO7cTvqauxJOm
tGVh56xlcCcGflH1mYJX3HKOlUTADZfk2Co+Qd2mjeTSLy+lNNTUctsMH6p6RDV6
/0QtxN8w0RwwvVbE6dX9crp3anKS0TrOdPzvJpCn8IfSnrIZ9NOiT0LuIfgfVvzw
9em1LIFCAiE21Q7svrFQ4uS78NdE7PIfQHXWUMVIQ8J2Enw4aSEJRJJNuR4SSYmm
jq/oYO+vDwT3HAjGKzxL6XXrYEwDW6CqZ5U+OpXxfQPzG3S8jf6EaQ9D21nqFIwA
iEdCSe4nYOHifer2zaPktWHS0cK+r9qQ2ZuKEebug1hXh1QsfT8WWxXmrUEPdh2r
fYVoQiWOcajNKCXzpxWoIyojmAUMGJBsoxeNrGtkKAg6YVnfAmJdcUFkVVryyoqL
hbxnoyGpn0TK1TpEQf/vcCyAswQKvkvCR5b0TJ8LhCRvIF122EoYHaau5HWCDe5K
7pFrszjNKC3caiInTS0nJUtpAifWvLGc8h4s8DFyio3w85h+iQsvKzLXVLIT3dKT
yz+G9/Qmm9izcLjd/wuPGQjwlrrxZqMCEuVsoS4KMYK8GxbWXpFpRT3K6WduNmO6
S0CY0ilMBi5MybkDcbZ7VY++sv/f0+SaWwHKOkUxMczE5EMF8uAw3/1wTv0iKVZa
jiiwO1toIBOpCCffIHJo00MoXu1HfrhsbLCarWLKrGFai6KNWEfJG6m+C9LYeu4B
4ZbrndCf4/8fE7h2wVzhE4ZzODdFWxnp2MToiEBXchCUJOAmNfP9RoITlTJuE6rR
JbJYQoRUuhuQtO7i8kYY04cNsmT/b2zA0ch6+XXot+bTsm4HH5cWmNVg7ayh5/M/
1a5chxao4kVhCDUNQhj1t5oTgVRuutVskGxqPcOuCTo2R8PZBx5OvcTn5EygYPGU
RFiCrAY1X4UF09bqha/CWO1c87gbV65B6/ywh3pIDBdY1e7dowPlwWGslPnZlXQu
5rVjms9uk/8pDBcSLMSIINFop7DK3Spl7hgbfrxvuhRw9ifHr8w5d2RnpcnwjKnd
tljSkdeu8EJCOnmX1KIr1ZFIGUb/Qfi8X/VknT7P+px11pNQzMEKm547vaHfFJiW
/JF2ceV0mJ1deCF1fh0f7jENKSY8LCIgswa32d0lVjzzg3tnPXYqqO5EdfsgvIpc
c2Xp34UbP/0+pLlHFKfovJqhTUACdfbKxyPbxOdCPNuMsmOBjIoRpbqAHZvnE+fp
ABVMH22bW27+rVd6X9hoOOK3+rkR6NHQ71eypEumWfBBCRDkHP8pTbvslkt1jxi8
TFEvC0sfZo/2DyIFLEh5gKNz4hpyw4uBSIRwYYsadF2WXdry0DE+n/RVP2gGz0EY
MW/SLx2Z0KaGSp0ljXiBFl+/01Ai52rxXsC6SLXaJjp2a51xujZCcT4G5m+WV9uS
r4PBSJSYDDT81ezG5tnz+XpjlQW3buX8e9Dst6iLa0mZrIY6QMYhF13Hj2nWCLXT
+QTg9q+TPFaaAO2r5VlFY76buwOQBzSotplllrXAGfzN9JCgcnjKcv+0PyEDEV9l
GJkvd+ewXdLcFobWn7F2DI2qbYnacpz5g+dMZKaDcxNgAPerSnih9NpNbs+m7kj8
1Uqy36kWhLtx9dSz0F81PLPfq+WhWoUk26H2hZ4Nn2mIzLpYj6Hm45x61imOe0Sm
fl1i2b8ewBE/K2TT+MBsycnEQxuraJOwhzTCbQz4guHwbWSvA6gIUSDftN2c+rCP
poWQi+Cj03KraN54NqQ8d0ERpjt8sjek6ZJpig2ICrJ11vx1sAm9YUIMccLJnkX8
8hpdj7zuPllgAFQr6Bj642uymrMYGscy/G4OM1fO7+HDyxCJ6QhlQmRJQL34TuWM
cnKsRJSWIuP47X4MxGA3VM9OcTC07TBjp+XAId0budSjRqw2XlMskZVUMqITceKy
lzw7eQah649MrDHPFHJO0f/qXdmCG1MhW7c1o5rKIk+CdsaxKQz6M5598MXp1W4/
GmrTZYxVVWGxHHnKlLK+/a7DnADtW2V87tthHwskM0zHs9ECBCjysVbFcfCt6oh1
rffp6RVCETtVQJ3hNmYMDkNjOS4rdO72+QnSJEya9Mkjplt5/bqGqmbcGGjvLoTn
zlJap3Ez3epqcwlt+5ZUJkx1t1Jc9mgvVLDkPKcfyTx6bK3Qv3GL/PIC3tsknUga
oubgfBYrem4c2C3offR1cpqJ/JimJjdQTRZxhKWkBRbM4f0MTHw9kREo35dyrbxb
K3zsdFttvh+e/EILgjdCn2tNY+NYQOXlS4Np9JXvoL/MlfLBWAdfFAHG8v9JWm0F
Z7UKojpmWaAMLQPA1eNgKJegAoRYOwkvMOpmba7PLaug+AERunHt9HGKx5PdQ+GF
217UP/PtPlDCg7f33arAPDhd6EJMz+T7hLXbsim0HeeKjzOwz0JC4tKTNq/9EYhb
22uyvZ8H/HbUaRXGxbt5kTPLQtF4EStpnT9z6aP2eniLs5qWHjD7bJUohK4XNMm7
IxenGCf0GIfM/nfRnkMZmkN7DtfGiE6y/S4GkQ34yjeVIGyyiIE1sgMAzsLc+wsN
T/8tIsoxNpXbyUUEMH2UB/NeXExnM0oyDZTjBIY0co3ZBWSmTn0NP3R0fMilbQBN
+kE+wWv1p9N7lRQLNxxSS15MKP3jRBqVEGY2C8k1tJJ/a8SlZOlG6CkvKySDUmb2
NEFJRaxLTu2AxnFggDwN8HS2Sfp0hG0puBBd0RipGsAIZFo7DeLuvw8Wfi32NCfh
FTnSj9xuCUolxWzY1DEoK8SBJXuVtjn5ZYSX66S0pqH2h1h8HzrpdVEekmnnb5N3
x021wyOKshR+mjtuv3Hq/R7MHIJGZx51yrTo61gj3yjEcyprO6nREtMwIx4br0LS
IcYPUDzLuP/Yn+Xz+7TzXcRurXdMUz6pbliBESIXE8hsK4mtPaIvTJYuuZLZbXWb
ZhcyXKIH23NrNTkyuk1HRfz0/+68y/7UerNlkXIpcwXOTuUJ7EI2a7PyMO3xpg13
c+3qb+DvW/9fzOlsLWqMMt9jYlaRbxI72UjEgNq4t3ii9KVZcJ1lcINLxpq1JKRP
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
N5av81+9FGvTDhYS2U3ErO7VMMwwgD1YZXCQvzu9PreORXqEEi0+OUMnXkEHJv7v
dUIT69M8oC54lCRoieHnGx/d2aKbE5R8763xlRDHuwLM8zK/mR3b3XwrNf0Muj8/
m0JYCLET1nXeFOE4+tdvYdBfunFH5dJHlUnL+tZlNRINXd+N/Hysr6zQrQdssRPF
+KUZtwjTY+uVSA1Jjw9WtdLc+d1MiwyHaT/jK/qZdhwWVzPBzGnKDFkc7Y55nCXI
VZVKVEFQwnTa+LmoXUazM8ybKTEDdlV4571lq2K5i21b2HG7SS0M24B3hjt/cC1c
xb5HR00NCaIqC3Uapwxizw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11760 )
`pragma protect data_block
FA3SDJ6di/2YHIl7TH1JS/YTzkgDbiiFyhQDdX+E7a0kbDG1SILmdxDfoXdhB/Fi
T8TYFpvF1tpPQ05GSp5ASb6juQ2w+TAf5f6OUX1OkbOaIwq993zTb6dJwTJ71nxX
wm/jObRZlWoIzGn+wQdU2P6mJagPArZiwjMirJcG8piBsnJ+IF0F+EvIeHftYfb0
FEEPSrhn4UenbzBTMOWjG5sQVBsZQuGrhfbRQa3nnWJUFjqvllCb52fDJ90oGpfk
2p52UdhWzZvpiOrMrOy8uf2w1In3C7etS78HmAxGUJqEPU4IZMrWCx+6rZ53LSDh
4Lxi8nZX5DV1SmU7kw2ybMPdvzeK8p52Q2TPVLH2sExVYdfF3+xqks5EwacUNly5
Pv/gN+N3PrG6EnV5yQrj57K7hH9PuVnibjHqX2CxBzyPnChZLJBY3NRw6SEIckCg
XCN8/BHAm+w+qQpNyTj4EKojote1gvzVAWvrAYa5U+y2rUQZumrevapE6cXODO+g
87Q0oASReGO014vGL1/MdlCIZ5B8NhSJWv1x9V0k359wUigZptT64ND5VoYzYdhL
Ejwtrjegw/riEsHGqTJcWWDhpX4rdx4Y08hAMj/xrJd70bMVBMOga/Pd1ReZW6J8
OJeqMEdwMY4eL44YigHzktsLwI7BLDhqp6VClZo1yFT868v9qEni/GfS/qcdBco0
gfNPXa74idJse33eFDlULN7VnJ1USvkrYvt2t0y0w+KGc1TTfjKfsx416EdJ6dYl
0yjX1QVwF5OmnHgZ3BT426vJZsNeDFuS3CP23sqAR1a8GPUlzhliSF1FzCmSD26y
Fj8szw/Ps4OorZ4zVJi9/Liyi68B7r4CIz4Ff3dzK/VUl5UX4rx0/hd5rPofwKJ0
Mhyu+lwrgI71/yD52qybOUnEzp/Ks97rDBSq4WItLuHjj/gPSL+EfGRkcqV+hGo1
fd3cE5Mnwlwpba4jYsp/ESowGe7/Ot51ayIOQdoO4ShqzhfItGl+S+fgmSQFkk0N
opJVwyHXC4wbp2gJrgjwUUjmQyNYu5BvoVN0X1O5Trar6PVHN3BkUZ5m9MV/hQEg
QcIhtfL/8ufv0IizIZZ2oXTw9Si+qr7lPKKB7ikR6Np+xb4IIVFC8bs1uoT0S1kd
E8V9svjwFlK2joz6xilY6kjpDVKmw+IG3GC/R6kHQhqokJL2Bd1BSjHgeb5b74e+
oVZMHcxcjUfSUrEYqDxG/dtPmuaL9KaelrB1MLF3pKrXP1YVM1ZhMHarAMd3i+tr
U7nwr+Rbl3kOl4GrIkLvJp1qKa5hU54c0Qy0m2/DaJan2c0LLoIT3JbRJsT7gbYp
V4eDn1kajL8LKpe9HGd7TnuR5nnX9wbaZxrPPIAfRTK3yy0tOryPoK9nVv7aZGtB
sbEZjikdpIB0GdORedxX80NinK4J9eXxF3Gwu/PKdyZX6zOO0JRIIB0BnrsLAqNE
XKEHIAaubzppNL6H2Uo0FYVTXq4Am6jZxQ9T2292H5hIWKWvHnZy3xmQyf3EdvoO
pjh4Rkz7kgQaBhqdA+oFhdThIsgjs/6jSlTi2YWKXT0piKLNxD43OVfefc2NA2V4
6eAobq1EdPC/iIJu97qB4FVCZQIEkZoKA7jfwKOje8Wz1/VMtjVdWERCqYjlN/o7
UvRRqbFk2AO3npF+8ZUQtmcC209mrVCEbql0dR60fYdktIbik4ClJXdsDm8o3l+h
gT4+wc8tEZKiEt1SlkSgJwX4aXfXgGHZgJWArPwqwGEhQ+rTYF2JJAc3wAXphKGB
55whKB32gFBHNcg83r1iU50eSMmrMwu1gJ5gmxTCd7zhJSuVr9vpzVpDWoile5nQ
2NrSh6JDXsbUsnrnxvnohqIdhd+hXHLGsRcfnTZY7cjvIxyhhUEE6luqYKW+wlhK
dJTDiUupEAjIUlmmwzJ2pGbCEvfBbL6xaX6sGC9B/E8RQIR4pPRTHCuoVdXR6IRq
iTKR+bpE+qrJayTY0LNA6ySsm/SLaqZPQU2v9qMh4vKt+7eGN05GiAn4Hq9qQqRZ
6nzJAIMDHrkCKPaxVcxUp8tuS/6hpz/xthKB2FaLHqsBqGPm/bvdyQQnvDwQjMB7
W8w+6FpJ7qjMY7LqzOsuPlWYrKWYKQQLLax9a/bLlkOxK8wf1YLJ0zWwxC1XYV+y
Zh0XU0SFzfc9wCx5kEpPLsxKqHp8r0XSSltosz7mOYyHBneHc43U13jFnBPIwRIK
gJmlTwtLWb/hOtmy3XzRKDCqywt10ojWw+SbEIbBCLdip01o5RTZDRIUeNThEug9
uNeo73R6HcSQGRVoNa5edUkq2B2+joRh7RM5sn3MA98wlIqKrdkzf6EuS8lD6LnT
Ed3avZk2Xu49BI1DbkL/b5/Z6j+YEmE/HsletyDo1ri6x8jyldFAFrb0qXYJQ0wg
4z7cA42kFu9zaKIV9mfJQE37Ef2Nc9icGGnRAC+fv8axhtMe7/1ozGZb3YAXqjEd
B4PyU1oI+UYAQbLQrrPuDDkM9jRC3O8e0Ra9K65cVVCQnWjLhTZ+DVWo0HXdw2hc
wZsfHy7PiXkHbti5u6RtWc4D+B74xmnF7ecxxdFWV+K31F176A908QQlonGLKvxq
5AXKSZvwc/OBz1E4CScoQNq1rXtQYCoGnDzjqs+DVPM6g7SN2JqVwmzUyEaNXoRS
H+/LixecxaZsLXuugF4NGyB8MmMlYCQiWiH3Jha9Zq5bU+D+xNJOaZ2hmoIunF8o
kkVmsnNl+FIkihcIf1baxYYjMvLHfvIriYSs+q/eKeFqAErhn9X7zNrcrki4NW1F
AH8WpwaXpe/uRVZ/vKTr0idpP2PK3EmlJrO+O2bfkQlWvl4CQLcETEhh7+IgSEff
6JdZHIBubZxpM1KN78ALaFlYxmqNYooNTOFib4ucAy8M6ht3a/wTl5iQGBSc8mv5
0kEPU7nBMdg16jZPcYZHqsxDldqDVaVkQ4Jbwtt7X3DB40NPt777w7tgw+80hCme
rnCHE/FnMwuQJduG2Yo9cA0fNX5yIlFIDKdgBWNisTicafvj1XbP/l6WHYUG/4rU
QmkMvlZPx/NhAcK1cTcfAT0PNWS5AtrsjdDbgJIGucVgcX29ixg9lUjfhW5NK/4y
T9lzoVRuuxCh87EKlLJ55+EukliQ/m8cHG2dfTghcxR1nty+MZdR/oRPbKt5CPF4
W0d1nXO9aVDNNknG2LIlmkyjs1dGgoNWZhNOCFtiGrMRfeYnXY8oKZB3R2YdR5Hq
D5Ta8cFpAAb2ao/Ai+HztDLvSY8zHlhBW3gv+mRCNbUBZORzhaiGD4rvXWoF/4zP
9oXugN1ZBflcmNXWyodtaK8bYfhatroMCJiGw6o9Pg2nDfuP78534EkgFXVzvP1I
eGskERVcT28urkbyYPUWFI3OkJGsQBk5EZ5KDUHH9Ku5IOEVb1nYh11EFemcqKCZ
QR8zFXjl9DDZ1UGkfa+Al1Ca3Zxxi3GVTS3fd60BL0N8MjQ0r2jkk1WHIVeAWR9g
T+FSmW5jdnfh9ukgIqfvr263UUC7VKq8cvyL3Uq30yBuM9re7TpRCtkN4Ukm4IVD
zQeJs2QqKLSZgWxFs0SewDYgQg6KxFYmX6ukxra08sIAeUtnHMuygO6zCOyz9GBF
0UwIjmAMjOaO2VHPKoOKiS0lvHF2xpqzSRAyHEacrtQ91Kiv7WuvoDoKMt3fwk8B
Ghyfoh8rQ9Wf4vYos+qjs30e1YhJZC4UaXp3GksWAVpE5YxpOvALCofg8CIHoakX
ktAH5LZlHeJLBPCRc6XCB4HYmsF2rIaHcfk4E274RLvxrtsBPqDyYQsUhgno5t2N
ftT3FNuSY329vHcysYk2GmBfaHnAWqGedHJVwWIvJBVBVORs0Y2mAGGEBot3Voar
xipEvHm0CIbVa/RBSR7mTL648sOq0XYvZzi8XhIy//dVBzkhxpL9SfuCVRptMB2q
oxpeJMeKv4X7G/S2WeubNeUob0cQyVr264AadSja/GIFBU94XyEcKIY7K/rVPonQ
pgnPanL1YfJ9tjT8EP2U0wwF6dCNJLambYg4cHKt0KyhyuLgTa4K5WJZdbnOjCLQ
Xd6o7TE3KgbpOcok117ClQFyMEenFdNaXzfrUTQ7mTuU85c622AmcFyWRjjOJz8k
MZY9Or3QXr24l1iYbpX9d8N/AjMQoQcuSy12VJqEUxKgbi2IU2p1zyNop/lQokkK
BjcZ2Q9LbLzq2/+BoQtL7YLcabSCqu0LsroDqNmheSnnh49r/FXp0Ojwf7fqsiNT
L76eDBvyEOLFnlRgNRYDoPJ3downG+Syf9onzY9Ed4wX0fx0DRl2OL+kdWobWHuj
XK2elqEv83iFio4KI9OF+3eVei57I6FM2tR39qaBwP//oTtoEymdQQZan8SmgzJD
LH/x5QBRdyIPQX2vT5Ixj6nd5H+dH/DaSo4HnpZ9394Rl1/k679geOv7wN3eI2iQ
z2T3sL3VUhlnwzWBlwWb2bC6qNKX2MkNL9OysBLP+q2PDpwHVzyMncew5MdfAaXj
6qMWhvzJ0tOSI4RQYyeNFxelRcHbwwVfvknTMJ7r4lZGK4JT1LR843LA1rEzUH8f
bAI6YMF19+bs06SGxBgDoYZCwu/pcSkei2+jhi6QqXuTjcRb1qg9m5xhvqA2rBLt
25tw5qQOBQP7FWGvCslaOXQDyEleR77AoQ/b/L0A1/2RZXxQUTVzyNgsBH+kpGtd
Q7BkfOhIDtcKGDBbmIdXFm2i+mGFpmLzqqbj1bB46lQNSYYWJE4FRkIN5MtUp0SM
xfMCunGXtuXqZqTtDywfpmUxg0KxIsoG9m2uAEHN3iayId2jdrFhZUuPhAka3oLG
UA03SiyHVAKhIkmXxVXKgreOL7dfw26I6V9Hj1L5nETbq8z7Y1pF+BlCZpJ0/8Om
DasZOi6/0+1QcPFqa+wtlZpp80fPMhawlrqbHGENvZV7Q4bCPQLI6A1DQNP03ixX
AgVudVOwnSYSPVYB/19m3S+QG4MYl4ZNTu76Gb/NqyZ5DjWxWVV85vJTWiA7FM3r
o6sTMrwqP0FgX6yUNLdyFjBzauAKcr2O4F4L4LWCPmmap9jKkIweU31XpwSJf4X5
Z+6qqBAd+kNy8ejgt5mPr2ABPSKWp8TjoyaQFMI6hFSEW01R5mOWW8BggQlDloLJ
dPA1p1LaASFP0goUZVzvFPhf2SatFj80+UukqPGagAg3p2Uoyo5UDmBW2GsobfWU
PcJNRHh7ygoOp4BSwApfiu1NpqUWeAkdhJ5cuCcDSdlV02aM7BErYcIjLGXjk8I9
1HNkTQlv8zLeRUPJunSIvYhkrXViU6+jusrwDcbZHNEN3DYnnPMw2OMEiRpPa95A
Kuf9e/UbqpDEK0vKp34c2D467WPcRnQmzF2gOO7GDnIl9gWS+l+pqKWo99GRYgMc
da/wMPJzbZbdTbGANao3fWVLtmB9ZLETywhKQ0pZyVbROZ++mtkpIn54bYcinMYx
wPKvNwzblmO/II+M9KhD/0O8SnxPTfJO7LgkDQAaTTrLanFsInEE0NSxOvOhK5CY
tc5YcKR1eAfv9e3UWzvkCyzaj3x/Xry37jxDCmPmWARspQM3smDUX/+G4qPegQBT
hD1nwUaBOvO1ifYH6zB2oqm81sguDtGAC4hCXDeGAbZWnnODBaIyQhSMvjzAtglN
8AC2FryzcuFkzKTuCzlCE7wX/FMuNA3qbOjekrIz+F52PBX5wmIjMj06yxSCa9qf
71af3RNu0yxM2kPJYb1pemkFzpJGNd01MnBqgIUGiQvCX+hueqXqP68w5MQbIm4x
vC0xWf32SUcD/3OJ2AEyf3Am4/6BBt51VMBxT+sNrj5LhIc2kM0QpN3/yivWr4hi
RC4HjHQn4KkIiHm8MRTpHHG2hIun62EgTrP/ekzZmlFRD38aBadkfzqkJPk5Z/KP
uMkBUlEsTpQ511DFIpnfwgVd4QfamNDBUp4OvVcXrrUm0dZ9aehOJCgETyV5kham
yqFQEaw6DMl/S5EMwEqfQJnab8LOISC4tLONOdeFAMQKDI+7XOBZxAdAMMtcSjdZ
E5I7jtSijy9sLuzFEYstgVWIl1M4NS7pKqTtLYYgCVPwxV/9MpRC8T7SuC83nqwg
6SMCzgzF3p46QFZP0NAElpa5GLLLa/KHiFpEtv4g/JLxMtJMZWw7vJfKbiNPRxEm
L2xOt+WqOfhQGWdDpbEYKHjTIc4rZ3qxs/nznHAePElQmxGylFe3VlZbFJ3xix67
lY5lFkqcm6tKrAGAx1Gq/NYILg2EQYNFFR26/LSYdKs7Ki1+iDxpTrV92FqSm/NY
4ChX98YSeqkTo2z7CfzKZAHkIdpybAJKA9H5whzeWcAjmriBem9f0Jv2mhnY6Ew0
+526hvXYz0vmhVmLdUZit65rQAY62JAlKcMQeFTLzpdhTXmh6q8LvvDjWoBDtiPW
6YL6aV1SM+goHtvK+9DfFx5bKyTT7u8PQl/EyN3vq4QNvzojs4v+OULIec6m64xX
CiU7G+tpXP7cSKavNrntdAEQNfg1xzq6Zt13IzPFzPgiR9AgGlaqvw2arA8EZO3a
NqkFI56Qh48fddKGhWgQPt1iAibHwLMIGsE7TlChLcZcrTnMbwHnv55ovAR5nS0N
HrWXWmVwrdfS6Ow2OM7B0VrEmPbsarjSwXzoDEWcy/CqKuRXude6+Qbke20Wp273
swQvdqXltlLnY5CHbc+vSHfL0nkv8M4+lWJeME8PaJCqf0A+RlmZcOQEgWxfv0kQ
znXi95xUiIxttDpbpAcMirP5HOIi7dya1hyDt07Kix7hDwrA6aur+m2to7gb37wr
oZtmx8G8hfvqVV+mw1ydpuSuDEr0hXq0qCyudpgzNdvA9kYNWRmrJG1wiYV0j/X5
wA3DQs3SXnW/8/uxL0xiCTadggx9XgUSPNlb8+exkVewQKSUQ0n4OXoJWSrb5VOT
34B4ZMqSSkzSKnsNKSWmONznV5XEgwZqur84E0UQ/ABxc6+JkQYU7CzXHYsB6yL4
WAiFSa5MPx12fnN3WvJUugBU+Tc+/Q85Zs7uT6YRkWlRIPIc89xdv4Bj/ljSNFjh
+02klfXVxXbCo20Dr9e0xVnUvox3lQaS7idXgqWx0Uxhb7MRVEH4iKZ2hhRbgoy0
7AFeLujOeIbvd2z9NFyDpN29IO90o89VFA/pBp86BRWOXMx/SsCcxVAl/TdbCLzx
3lg1l8sana9m5xKzd7KAJ6HxMgqn2NBJaCuHMncQFnDAbBgt2zrEendlDhfVz322
s8RFBav6XHseDsR1Gz77zcl+ONyFjt3GHmpcO30SNGONEiauTXV5rwrsk1ONm9RF
gSqia/o5ZFYFA2Dooqa2KDX8cCvGV39ch71Ms5lOgUfkwbTYSjkcTEvf073YhVFz
OVhLQDZJV6DAuXyNVyh0iStXx28WFBydbaz8U/kTFs6M3Sn6QFMkEV3PHb/gKlks
trO5WbsTyVHzZfoGVOv6pRcMkRTc2QgW2zlLQlQVnXleh9le3Ry5zHFHzRPWTJSN
GA5CEjMsWk7bJqlCmDvdqB8asaQToqCuFd7vSuEGQ9DFmF8Y0SJr3m4bMOVb8CoI
9AebY1paT6CBeu9ofm0KZlnw8GwLECLYr9Ywi1p6oCScrCTkQTBkhcxVOd6iG02D
sF7+Cgje23dUpcMRbjlmsCRG6SZ3+7UbfhwfXFLRo8+Ppv5/e0KjAfd8qEMZbkhn
An0O4YiaNH/vm2memPECeZzYa1CU0uziJXFcjc79S/kyAeEL3RtsLIOQ4UhoH2vM
Bk7sXwQUiM/m3s/7/TxtXa0YqeFFGydcud05qcUZr89Iq4f8RYKns0ugUVgRfaiF
ZCSQw75lL4ioLO8FZx86TJ39me90vRKHwHMRbEzZ9EfKYhbOYTaA1Ze6TZMatDSW
lY5bgVBx/smebJK/nDe4UEchG7d8jR+knQvZfdVRpoMLAU1Dvue9LqcPNrJOz+jo
ARDTelHZa3pFDTqGtOD9dB5+B0/+sFO3Uwts+Us4wUOXCwZMtQFcAFsO++jMvoDe
+klrASuLLTwdF8B1sXb6kG5JMyZjlq7GaC7IHwKUZKZRFfT0OaOX0a3hH1GM4/Bq
AL9YG3+e3p8rJB/terF2JSbrK8ciG1dEE18J93LIdDN/yDiY5Z2EZU4/eYgmSyIx
lKEGbxgG/uv8gB7ZYMPlrOzlXVBRkM1WPu3uyjgpP3T9TyKEPXqEbHQm+RWisNJU
QeqEteLx1PpYiCM5UyQ5uvgTkPz9kn9qZ0lELq0VounN1IyHLC5+4JShuqkD14Vv
ajghLWpJ3j0PDFOUeIWIVqESfnBzX5LY0VOBi+YQPG+2NBDfyoGC0CGI7qn4UfZz
NdaPqz3utsfAd3Jy6D6lJ+dU/hqWCBFpmIIGceOJMVvb3v5zwhGkNc6NZu4U/MQU
bblqbIZs3FrW7UiMwDufPbxmiFqI0NRCxjA+pE4acfHRokjJHVwvdThLbpxMePcA
Ac8Jrw2Gew84a72S3oaRral5V3Vgv4JMNcw2R9Fo16bHz6Nr3OMEshtjvELgPrtI
lSr1rLkRSA+0p8NXX7V1Ms1xXMJMuv6vUhkfojsZub5NN7uE5rSuqQryKarnMwXH
60lNOOD+n0MBI53O9HImO4/+GIAtdL0LveqBvGmvuAGOrQjgOhkIZMAralD0Xcfd
BnDqoMyKpp6WoWLXaVkmTS0VA9Q+lRASFbUhp8sS9ZG4PbHFo49TMlKAU7cTNZh5
gMVRJCOHSIoN8f3MRv4Uu4CEp6SMXjKEP0+AxdBf9yscHLElRtqQCgxAwZKDild/
BokJqrNY58MDSQ9VTEAnPAPdf8ap7K94Dw+KuVP0la/Pntz6kOmAfdSCyp7biqCU
62zr/tJzndwin3PQB7DqagA+uzuGWrDCyDVVrC6sWgKfb0gigyD5rDWZQ6ohCgkk
tPdb46ITCwj5wmmZTD1a5fWbhEMI+HpqZUOfzgnCUhxiBoiwqqYs+v01vYV0/ldP
czoB5tjUhHzs9Xi8baw6SGR5UCQKdKIzCalTxFEyt3eaAQOk3YgSF2ZfHmLqp80b
UN+6mugzx5m4oAfELPrG2QOWeUeZBlVYV6P/bsT4vzpKfQDlmsts3/N8SsoR7w0/
yfBvZq6yXAS6hX7fCvyb7DOitGZ7h8qA4SWEMxonTItK/FnAM49d2/vTbTk/XX6y
GUSypX2n5nfS7odPZrsjRvbVJoELkzflFFpkBv7bO4Ezks4A/2b/Hk/XIF/+AwNH
3KJRKaR1l7JsQC1mQEVtm8hKRy4FqUkdz9P5FPpBtZGzIt+210jMDylhvFblHkUr
IHANYNgQw8m+vI95mHaDK9Tjsw8Cr4zF4SmC9sxcB3OrwxMy35QSNlTWR8Y7F/kn
1uYtDSsMnBF+0bg+HJ6eD3Q9DxVWvibXReYMnfjDCJgmurqGaq/w3yKo/KiXWIKd
MKug4mrPaPfs0t1IfRXwXfvQYUEoCI3rZIiXOjHjf/HB4IR8eIcdUguyqGQallgp
MGWwsOYk4b5RDbGFG63rjcPqyC7+FNJDgRWYfLCVp2SIsF0Jm7lkCD0fBDeZ2U/q
PFhU1Z25V6bg6WjAi5LXWivA8IEfw1tXyjRGXyd5q9PPkxXDtEEHCFscYbWkaQJH
07fMarrOeVQ6y0gt/e0BeqLpnOQEImjezy0oQGC071pf3WlGMXrOKCxDyqO6Poaq
wiy5/ZzsEmq3xhvCkN2ek05LqPmws1jNqQIsilLmYt5DK8z1Jge/qvVJrnJa1fan
yoxMkC2Ahjx/wBK7eh14Cp6fOh7lrdCBW9YrCN/gigCJd/GVoEFbt2QFfPH4Ot2p
JZk60ohd8L7soFTuJN2xEUj2BhwvzsGpV+b2g5EFXg7bvB7kD156ShzlYKuUnGWZ
zKLCNHeJEAn7kl131jlkzxtsek3ZF0B9pil2oMRKNHH53H6TPQj6D9ChmBo083y/
xVRrs6UW7UgOZmAwMGf8PR9OBsH7L2EwqCzGPXV19zgrkyJf/owRI7qqqhgkL/m2
th4Snk24UyY7W+K6f9GJmasd4MLPQY4dy0nTcM7ZYsOgW8gSL6WgjOLUfOL10ogc
FSHRwNpKC8OGcWE2OQ5Ch3/b8OEd5C/UoXAjl/ThX7ly7LKQNzttUFXI+aFkUkBo
UqYkbrtf8BmET9vS6XxJS1u7fYLZvMx0tccGGe4jRj1O7nSweJsHIAPfJaPPOF+J
Sk92QxRlLXMI1uYf5d/5Whc+e12FWSPuMPbzeJZuqkU5dIqbD1gCVq2dU/kDvZrw
k4s4WoxHeY03NixhBKRjr2zmmoy8dP+nmWB+M/Nhs+Rk+Th5eWpjmaZhSHzmZ3lG
baiYI69WFS5srLJyVv+s+QFq2xRsZC9GRq39zTgPJABh1SD0NvBpvNaVMdDAm0u6
EoeXVFnMoJ4IuDsq1ucyTuvKzKG+3Htqs5fgXJ51OVQPUL2b2tnhI6KNpfwcrEce
pRVqFuu7BNzjv43jhigY6NIN/sRhL4B3dH1Ch4QyUEVZVIIaxiFRwL7dRlTSs7+p
LVcBRyUwedntV8LyEqBLqxrHRsO2GnYJAlRwneUM2Lc29SdaWYLUWg4nu5DUTTeN
M1KbgEc70op0zsJhWbGMLou2vedZjJZvNNzXiXdXIuvjcm6+yxwDMYFA3bpgQUcr
5noMxTWQB5Z71gjSzvbex/79Oue58ZXRA5wD7vsRmLDBtub5CbS8loCHeDSj9DgR
heAbabIlgUgdPAp1VLFj6G8FbxUGDr8N+4mGAlHb4ulprSUReKMRTzjtG1HhiUk+
Uf0CKdSRUtVimGWjhfLfByxqlakRb/QZB0FEFYPf4LbScPpEHaHQGOI++xHIKuh0
HiSTbqPsCmCFb+h5m7PXgDX0rSmxxs1faeFwXgr3+Iec8NSetJFtN13jiK7mZpaW
f0le9iFkN4kJLm4BUYBiYDFMxaqQbPR18wiHrNJ9FyGjUuIGBgddAfR3bmpopNOz
Y+Sr1hApU0CuJDZ6IjXl1j/1rF/kXUjhPDszPnEno8qcaZ051LBE+05I8u3CirAu
yfOjA4jk+ATvqhEqhgEwmwK8qNsXk3VHS7bpcqb+oB2Dt7yyQGFqtgg9U1GKb2Xs
nYZLep10EzlpZHwFv6E8ps4TRbbjRqg7wB4uR4n1QwR2Sm8W6qIBg22i2cK2rjbx
3xexSxFrH75tOSpNYKJpmHo8F5RqwgFaryMZPn/KNyLc/f7OrIhO/oBI9LdS1/XI
h+eReafbsM6YWc+ll1qndedkGgzke+mabHCsNLZ/QaQdmwmrP0y8ZwzWcJMGb1Mz
nzqq7T2icGEJDJGh9a0xxX5pIHqDvIapGCOmh1whPchmT+nDu40+kpfeXPC6tnOR
HA4OrXp5OxfdWSg5gPoR6sEwi3rrUSwdyPJ3wlGzdELPEvyyAtvHyG1M+X4jYOQf
wbjA85/XmUEOObtZWWsrCKrnq7xLV5BzGYNSQEShnSuzs8oM0wVY67VttFdTuwpB
DUsQy0J07DI0uugWrGoo8J0Eg5kgqHWNT5H2Vhg4fm1YWmfeEjzjKXrTIpe5MMAe
dgWffUQfmYjiBJlffdNMQGcRbakTYMzpTvX2c19fZQEFE9UKD20hLrC96wW1b05P
dB2Fof5v3G6sevhKZ2X4xEkiq7n301bUq/RBNDt4YDmY0MNvqwNDA7JGKElWB89A
X8BcgdylebK/qbmxlryH8VFMTxzH00TQey/BZE/49LVyCOTPWnNfpWoCBSojuGpM
NCWDb2v3c0m/ttIle0b0UFAmi0dd6GH7RTLfJ76WJlGqC2YRMc6npAk1Q0xNewYw
JLb90zxIbl7e6hIr4PP1+qK0VqPLhC/JjK1ANITlsUiVTp5zRD2EmsS/I+GLEMTZ
sNoq6KC3juWHuRa9vO3T++tHOcvoNJo0K1swrOVjI2yvCmCfe8dtKtPhwmyLfusJ
/mYQQW+0eznEHN8iBGJL/AlI8ke3ilKFtzcMxobVYyqkLUQ82mKU4xI0eZa7E5KQ
uVMLElbLB0Fa1Kg4QOaMire8n6ZsGWnSnEZQuZr8s0hnyVIkElemAIIO+tkfegAq
tOKchU+/lQxycyGpjX/2sL/8MUSxB3uLjOYPueLQUQ3TDoM/OehtvWOHhsIUQNxL
9GT12px+4QQW9eWSoKR/PkfT58XG7QbPPd46AcSSR7E1i6vqvr6rZqwSnlZJapme
Mox2lShkNn8D8XYwCPOESh7HPdIvfFncPTWtyUi6Wmx5fciA9V5Fa96nAVFrI/qb
cy7DzqdTen2us3c/JXpblWzXuMZRl4bmleLCfaXxqee7O5AXzuBkXbHIqLgrm9xO
ilS/A6t80fVeI1G7zHf8OaXGfb+D+WsZdQI33FsSJyHH06acvlWQQgq7I1Kn4Eki
fKKkrvIxT2TqZlyMwaSjDl4R426RYgxZ15jTJ85CXpVb476fPoALdA2wTQLxnYrb
9QwGfK/fTJROu+hXtPReXnSbhPV9GTm0+wosMzvevrOwYzI/y1hVjAnx7YKiY6zf
dy1qywjptXWrhBxnPms3Wb47Sy+k1uYXMuedbz4HFi8sxk6mOmE2ba5gna9Okytl
MaAt1GYzgOkHQRXmjJkIi92NDIiXYt06UzdONqQkEQOsEqO4bQ7Cr66fjoWaRFkq
bRY9RSUM6VDQWWMs3aoWNg/xqo/d++A3DqkeB/2nhPmV6XwkfSYX2uj02iXKyQW8
0bAx97E6/c/q6iAjkmqPyHExQeEoZ5T/SuZKb7ZMqdJxnfNJgFf4BJNEsKjj4AE7
VvIPWCKJXHYFr89/+eFqkJNgQowdyloxE9SYF1M7hrfuOivVscb5Xzx+8/6TMfvY
8rYKbGZqe6Nl2+EwI/8USG+SS5bAqzY3qYqeFc4BhDRwC2036xf07aY4dW81kRNe
jeFB59YC4Ji9SG8mc0Gkgj5vntEmvMmtRVXUZpLNOo+wWc7hjpb+xuKlEtfakEeu
802vg6rPrHeeKh7Zw9MMO8rcPePcjQ06+lJp7pbqV0ZMKkXfZDOR9rN/PYbjzLxO
1wORwSJNOOjA3sKrAMmbcYEG8wEzf80g5CVChFIRW3LCSHdaRZBfdqwzSMU8+sts
VGnWhxOOitLP81YzdVfwD+D1BGZhuuZR9Fz/uHQhKtoxCoickkIjk1hds+y6CXOQ
LvSBA9g59WSLCv/Nl6lpEE5xpdxKNfrChPk4Q6lPSMpXcuvBW5xRyr3hy9i/AxeC
XW18SO5ab09zTRmFLp8E1Mbofr5dsQkYvZRfdfnkYCxtKAlA6DKNGJ7E2ZAcKw+T
3DJxTL1Z4wtynLAoYmySt3RuY4yHG7bqZR/5nIDko4tiG+Xw9l98HfOe0yhO2+Cd
PKIfl3S5N+zB/uJfJZJ50E723dzdaK2vCUoPFSgcEOPcVCaD5Yr/wNb5/KmDmrWM
FyPU1QxDurUE4/lTE+AFNn5C84I/18AXdjcFQJzvoBWweagGOkC9hq3aHDCsiG50
tCmj6CTaAoe3b542PEXodD7irYeZOlr0jncXsx6iFFdBp9uX2kNey8Ih5KspoYNI
Gv4wpNJAwE7GBKEN4rMfNOWzxffG1Cldt3UNfL8oINoxdFsGRGavFv7S/dh60ru1
QwrSqvWt/B5HOF6HanoBp6vu0K3J2/6t0Yn52/8Y+q4Op0GssQDWJ0Zxzo0V/iIR
/oE4OCWcR2JGmyy21Y7LxixmlLhLDkiVCzuKxuB6cdBHoemUzR/qefP78G+0fwfa
zyyJ1SOgfwXdIvgv6ayeujgj0xxotPHJ4cVr8vQznfrTqFbhO5SsTIkna1rmXQs2
ysU2T0pQuG7NVWGx/tR6s/4sSOJNZ9b+S/NDVimyND4AHZ98J2g4xcV7OYtx4uVk
C4bn8uqlhqK01IHEKvggubAUtvjCiF1asqr+rq70Oinsm0D9Wtp/cIyQ823iiMmH
UoC7eLRIM+KPSSVNG1VKcidB+raW/Z/t2KVUbPu/LTHintAjpOux36ydC2yY+M8j
wgB+95mnyRfq+rFKUxMkqmbxqpc13HaD99ouLuGG6cHDsqXOSAl6i1H5iiL0n9U0
e/F0lCbI6A15Kydc32mhRz29BeMij6NDvXXvod0ReJj6Ayd8DeEiRY2bAFPk63DM
l7cBrinl238xC6UezbicudQH6z8OwbtbYOx0ZCn5z+ilcdk4Vw1ocn9Apop7Zqkq
b1BdnCmiHHer25Uo2C+zUmA6KNPJKLW4htzEnXuBO0yJ5kIp9vLnluFVMnSu1+6h
9Zq3pJ8XxJKYxO71tLCGbmmRzCvZTr0nofGm2cj3sJwABxF7m7kUghQeTM6o1RdG
CMZm29dm2GgKk8VRfPbyCdvAF+a074EFgpQcPiiF4NW3NIfHQJDYmW57fx8jDJ4d
yr9jkfealJBhjXS3rFWqIflvcqRkczZQTYAKAi8hs9Q1txjE35eJAUz6CZ+VaVan
+GfHCeKK6iTIFZhH9T0PE5T0BPRGIUR+E/RSUdWwhoS82iNSUUbzqPLJx6u4bzVw
4QbnkD5QbeZdXxjw9D2ENEESnx5L8SjesHEjv1SW/OkSnrQDdZc+UcXkrHe+gqR/
+ZgBp443pFs91FZQOXxycriMfmJpERVjvbwfPHakfgf7Qc3A1i5ASrW9jAeK4HXg
fa8pTn5u0KtGuLDCixt+c0nOKkNwcgf5ZXVFnG4fafyLtMMKtPkDiSZ/gjQpeFQ6
g53qZ2P9fjBUQfevQEsZdYAXj3XDfmTWDHyiRDpsJoNYRZOuekjpYRC4uyYPvluh
Sjv1Te9TK+8oP0Smp2aZZOHbX+fvMlUtwUm/Kg0q0+AamXG03pA+yF3DWKz5JkwU
vqXHJpavNwhHwHB6LTkhzMsZyTIGg9HNsJNMBdu+rwv9kLUVPVC6sLnl69XUy+ZB
i7JX3Xuf2bm+U057TPayJhXTHH0+PPEpo94r4k2kjOHqdzKDRZlakmEXzykx1Zbf
tyZFg9hxt8DbDRQVk5CbbFi7eBvOSDkEMSXMUVMmj3OsyolbqZWlD+0v5Nlo5/TP
4UlwNWuITOzeTHFEZK75r9moBtxg2gPxvI4LL57jKR06pL82A91FG4KdMKav9QBO
LgleSkzdlo79rGWZt2ACfbCWVuE074mX0SDj5OuR5oTabYDgLjqC7bWF/sR2FFMh
CM00qsIWdexpbTIKBUNqdjP5Q0pT3msEYBiK0yisFv5kyR5NsnNgw6yAc08TefKg
9Me94+MjPLX+d+STIUWM/ndQXwwBelKoiHxxATcQHwajxEgPrD+eoVcxoA4oNw4a
VbW2soud7qhxEHosgcrXO4WJXVDi8sZ7W8oNziNSjT+WREtfpXxOwcPPxPdtu9FN
iRhb8lmTRuPvVhGm9p4jYU/yIst2jJ0eboL79bXcrphPmQXhf+NINT4ezSPF1adw
QQWE13YB2MACqPFsVrKbpIwbYvHJ8OY5Fmc+1ReJ5SoO50bfclVi1N7VxAajM/Iv
PaOTtW9syaavACQbpqZmFdYfzr6naBCfjd2cJ0ATEd5QNFOnLvTyOrzVN1vxIJfi
hL8Dvm7p3ATyO14ui+FclOKh5E7FglWYbNMrkRiQoHiO8M2pfJ3hhMpMgiatxunF
oNR66t2n+Hyed9v6VQMgnYv4E9vJcsFpC2H6UoCBzF++0oxUk1BhjZcNLvhla+uE
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
MlY8Sd+iZTBoanKer6qRN9+HWxheJ9oOrXKuS2uBp7IIDIe/TWuqH4Ml1rDHTKuG
x5v7znHs3fBalFqc2qyxmi/E39Dop78tFrYY5m/6mngvszXoX+ReXmbc3mncJFG3
nRPoMp06drc3PzT1rawZTPQcENEnQs+04sNG3/Kkr4F1ozYh88DDeE+1M8sMon9C
bVS5zqJWplJ0Ihull8mWL20z08/K5/froYTUBdxdqTjlLZrpE8zgM/6TYikTBvg6
yLXrtRDUMX/7OO2eILoqH0gJei6tF6rHt/1kzQtDOFZLrc2g6wdSiEQtISuXJcyG
OOUzPZuLBfaOHLZwz6U3Sg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7520 )
`pragma protect data_block
pEXSjXnhPgdAfCet0HUvrE1NClRHa7uW2Nmuja/BMR5KLVLJN+UXQDi1E8uKzGZc
LIAI8FutiJowcJo79dXa16rqpxUI3rQHDo0TXt03FF0fasgiz7CTadiFXTnhMody
NOn43zSKOZ9RIzlT5JrecdMeeHFDrVERY0Eip6jxMyHRdSCYpf1ONhE1vBP2F22V
3A9DP6w14APgTZIdfwll7BjaBa6YhmAw9GsTPi5hxo+/FqjJ7/Fe+bINC0CEvM3D
wIfJjByCn5AywKmSoLAxWnbZiVgx9WmhCat6NypRaVkbibx/3T34CEiPvWUPD4Tv
m4aLPeybc4HrsSqsoMhRra/vFrsNPIo6vaqQZdf1uVRc86WJVshdKpsvsUer8Z8w
qOoriuxl+m4OeZUjTAmVhho6kc+szBG9GeXcr9LPtIJ/gGkqqvUJl2d/bNqM4qTB
CSWK56YcAqmSJaxqbdCEvseOiyi6dpmYuOvl18FpIKdwKwN3W7TbetVgynng0psF
GeaejnlVCYAIZ+4EuTgeT4wvSd3Pf6DvARprW98RrE71pJLHXmTDGH5QapIsuD0j
Vtk10dpqPGjBPWpBxbXy5LKGpuM8QnFqfpcjJqAUUUngeGyMAu4PjoJkTIxc/9Qx
RW5+FJNPQi1qtADPzO/ggTJs4Hkf4oEQq46vcjOfzb9m1YUkuD0P79hR2NjKetMZ
mOPyQ+fJhf2zsS1xw4QuwLTpLfVzCtNEHUWn5ZfZ1OrGr8U3vbUyMt/oqMlfeqlR
odqHOoDKN/RHUWAzeAk0eGtC1gspMxpywgZ7RENReS6RbLe8zZKbfWeQGqxzLbCt
ODy7BspP5y2vsPe//jA8WkMqdrjf8UJMtYH0rehG619cQYxDOZ0v4P/NBFCYPhAN
39bxsqxUuBZKPPsJky4Uap4z5MuZuKEOtCX54eNh1YkVK1aNNfy54zIN9X8yZgbG
haZbXP6jB+olQH5uQ/lmILw2QmyEltAhoiL2/OeE7jxEtgyWr6DrBIWl3zdPAJzi
FGFPsCS1l6Q8a93sKs36R2O0ULW3EPdOx+uRBmEsCwkdbC2K5NHAhua90sxeKmGB
EDnakC8vm9iNM5kEHCUY+1wrWZSPRwY0JkGQJtuejZCq4GnK0wab4Zh6tnkrp9Mw
pgZa8b/7xVqxd71EhvqjM+0PLyIEeNLEPRVA8eeIMABaoThQCVTKMhxgLgvrtNLS
/yOv2aftX0Ara26qwd5+DDpSeSqz/bILUigPQR8x8FW55TuPR7JZcLQAoOyD+AAL
hW1f4TYH7vKHdNtnsWB/0no9G0FNmDQ1EUOKlRvsf5whv2pTIte3Pl3DpJ40houx
/AHHE/TLk6DocEqkAoN6K+het6lgQrjchYcffNykgu1zjPWXGP8UlSyDbPRCJiOU
LOw8dmqdSMwbK9mDxGh1sfUaeyRIPVohqb8TMCeWjy8krrIP3EjT4qpHu6aoal8X
p17FlH9eC2ME0xg8NimgpUlKbSw170D0y+6cR2GhdIJLMsvCxGavVSNkkfCmhHUQ
J1VNxYeabtFShLpADbW+qsps1cTvRPNFEga0WC1wiJQg529VItmOolAUT3P/QMJ5
+B/I5Lxwysavn8nS1A6GO6nelGCJXrG/0Crp+ncvW+XhxinExacP2Md03+krr4tu
i/ID9rP2jpwr1ESVKyPC0sBs823xsvIY5tBQLiNQy5P7g0VjCH8cuUeUxB44R40H
qJphQnkXro0n4Ym2biBKcFWG+YopyA/88f1dDim1atTJ3aYkDGrs/r4QfWL9ErB0
EipLRZFP/1lvsei1zcfogcxE/aMPbEoxeQ/DKXw18nx9EP3ITJk/vwepjR4ll7st
ncSnoZoB1jSMSmbXm83sfX39UIe2pxerGDCPUqwiz2vlH44kQXigOMLhUQ+nWBAA
JfzSjIsA29p2Q2IzZ06mhaJ6g0fSTJuEPmA4uWMdT+URkTfpuq1xoev/nTFb/zKu
hL/9MRPrMkXHoIYIaKVHMsp1VBEXdM0eKd0DVLIgn+zAwVDqQChM+yRKsVBBaNxk
e8BHMR9tb5WCpR3tDREjAuoM7ix7SGLhzAVHnBeOpCKmuvLFW+C5WPPRx/mDXzpa
D0Oid9A6nrXnVhYsORO6uf7TnOu+yZqrDtE+av7vfkkDhnw5Lqwg3Z8XSiGKgXha
pga/pK57jCB6DsTi8vu5KLTpizHCp/C3Xe4BX5bX4u0vMQlypSSHyliKphoBFpL9
8GUld0/HUssGOmA8D5xjFcab/h1zDGvLX3Lu9HDOWpTBLJpaHk2isBQIBVXasaNg
ExEz2CbJtWQ+o1iYALJG454qeHNVU76QGoafcH1qWfXNUroVOVI2lPZKzBX1UBUV
qvOhxC1rfkV5+/zVzi2a4jhObE9bJZj/ncqOZbux8wifuppHmudjVN6Q/it9dYcX
zKs0bU8Z01RtBPJLICtnOnadLDILxJgO1Zrr9GUcz54hjC6JqTr4Ydw0HG2I6rYe
bWjDTyk24Y1YToYoMxy8JGw0h13+TCxGMXDohOOQhHBIuR5FDxtWuHyDiKyu0cw/
FgfCR+U0X5C0FuX7gyGDTq8L3Dpnl57wYbwsC030pucKte7sytcQoCFdi6QtiYfo
ywpea/FQDfYejwnjtl9K7NWL6KVhJuef00+4PlYz/eFIGw1sIM9Ro1o5KBHE5thy
DISA2Pui5E59B692UwjAyygy4v15RG9EP9ZaBSbYH+s0LpoJqEzE4zfhyQKSolBZ
Om8cCKAQ4Y60ESz/Za9GZxfXWGbMazioxwYQUfsvqBsSXnjAr6+OgHfH6Bt3Olx8
+3DpLzHrXv0oNz/lBDLivOFPpjV9r1wGlgioZz+Ao/7c5ejUOrH81SY4aOU1AxIk
E/yYIHsuWzsJ5xFTAFI5PKDKI+ZYA61ppuW51KVX33JRardpWvts6fi/HSAIrczo
7i3DOWBD/LU6lMB3BBFYilB0g3wQx/YCjb2Ht+R4vrKRdeaYe/pk+o2gn57evwPm
bYYuL+/uY7YHH3PaQXecBL69HX3Wfvq4p6ZLCmucojQQx6pIKeyWXOzJD5QNNb6L
zGGX94znWFSsQDC77cSkF7EEuqwHqohva3zdkt0JlISwS1iQuWtNEWfdJe4Li69U
CPCpUN1fRJKLwGlQvyzWpxnIdTZqaMzREwg4VpW9rXPdJIzy/NDSZGMW9UpCZo2V
oTcxRCBxmWo1YLrgBXnqs6jhTAw2x1XkgCAZnAmvsWmedORa1f5Tj6b93TMyyOUv
cY7qdIw6f6RAQL0uC7pAfJACa+8l9aQsI7ezQSGv2eq/anfdlNdYrq4hAO8777HT
LDNQ9e93hHblDDAm3bMeCF1zBghSoDNsnoxP4ZCTfj/25nM3mN/GuhyhFTyrUA6u
ir3QTmaWNnj0KyQj5h7DK+UaE8sG7s3MoJ93Ysw1NX1c1AqE4pJmEJZuvcYOhZca
c3lLfRIvxpX5gJMugSxdZ0GLTJnMdJKP/ApBUns6Gy15ZicSeCU/HHtcAct6UbhT
MwhjumLLpUEe29lMBlPvnFQFYOUPAmR2WdMLttsA0LHpP6jIiHLwZi+otbmvlMcx
oveO765BdjKjaDEmbjMcpN7UTShtVO5nQ7NCnDFbfT2s5K/cDgo7UQo4+41MyjVX
nvFAm5qpb6U9HT+X+UZTDVOoJw7tfIkonXPC7CObuHSI9bpuxGMr30jFu3t77OAt
oobjBOA/h6yrgHqDoa0KOVwQ04eyYid1uogSoA3fXS5ceJrL1PNaBCsUoiM0nPpb
czpYUw6C4dbxPTufyQ/XRFkXGQzZ3zcLDqfcrl9se1gGe989Ps+1X50aQspNIztq
hQGh64bxh2KCwTA1v5XbSXAeO1h8pKV2kJwTy7uuKdRR7XkWwU4a+9gutUG7131v
4M9+V8/Q+fjmPnxvH2ZlwS/rG2Ls9ViW0CO/zxP9K7KAZ7WgfaEsXMaZLqTVLYy0
Rq78LWP0sm8uoglEaMSE+iXGVBhexYKtgWdNmUXJIJsry/K9e0C6CTJqF6MgeOQJ
gstOgmwLQQXLUQlxDGEIDKc8toClhw0R2UPFNyRt9i1OQHEj5ycajktX4806hEyK
Kp0xryeNcLEmv5ytJaIxnR9wsRM2SwrVryynRamF30I20BAGoJp46jcQEqYwYF28
Cux2LUXVN2BtplX9DE80WIB03U+rQegsDdG+sPZEAd8w2wtwSdupTjCMD/w3kkHw
Rhn/YGZ3Wryo1UX4Gp80ai1LFFTWm/Cw5zhoTxnmZZUrITuW29SG+3T+rfoaRxo6
SKMMZbcZfqES7R6VzTNCGzV/Rou4RY1wGfFSEDw5SpP+f/Ls4OGiGXapwTh5R+uA
kru5nwFNOMCf1Eo4eg85deNMrZP4ZuS2NZjw667JNX2eJxNbszMDv7jFXn2FiPrM
ku8g9/rgP5IZJgJvY81kf2t14ijEzYL1UJWALYgg6Q3J6Hx58ZB0804BE1zxrhKG
LMsQ7roLxxj6hkn4xTEuNqbTSSNH2vDYA3bSna7WS3CnXh6iX1bh77IyGo0f4oaT
vOFaWrsRxaxX6OHzpi3zFPFULu2E6hSpSuFjYWO+hVkgwFDVvpRyAe7TUMxaYeol
KFCN948rg3BrE6v+vEg707ZN9PQFUI6gFaqaSccgLU6VxEFsikfpqSiFv+F/NhDa
gP92TEH7jg5cL5XpBHpbpgN5MgKLWbr1qrctDVEnFK1KgczEUDz8VEO2nhTnz4SO
gHPu9uig11zlQFVmQQ6aIKPqSKbh9Gl3mQfjJwu4bUUQ+pDwNd4/r5xAhaA2Jr5U
W5zGVKqrbGJ+lR5ktOLGTM6PScpSKxvPUNsZMYTHkRDPmFtQuO5jXJRmO4V4EgAj
gm4vpsh3d4E9MMFvQNwXfzaJAyMGISD5D+NmX6+UHYEwvcwx4HkWLwxOAmiD/JLT
zcCmtmImSqFFXBqFn4HfBfdHzg2jDGmnihRtf2qtTwoqAJTTAcBidE1jahYrm7ws
J9ylQfnrQKXvdMAcu58mfx7zcCHPNCesYcsEGFv+qcY8ND/mpgzaofpN3mvmG33F
MesndCmFj534wfmdaAX5Lp3h0VyX8YXnxApzug4wQzQB1eeB5nCqGG7FRrwUZ6TG
fMwsjB3f5+WAl6tExBGQOp5mCsP8SrOzN/mUhDefHlondzLOzRvoOyK016tyS7Ju
JqKvQccYJiSu9bnLl+NMU/Nn6XcpDzOhTBa8vUto+zdu6m0HTaFOmy+f/mlH1iOU
08gAdhP82j5zOGVmuLkB9Z/+h9tefgSFL20ffkc4cGXelNN/IRf7DpdaWd6Mz3tA
PW/qa61k5SQfLK2AGElJpaCj0V5TPZh/k2xcKI2bdnFUx7lJtPcfBY4HHtElngJH
0y5wfuWOYafB+tWxsPMsMSOD3b1cnEP1sFbTd3PM3UsJ1s3t3/srTlP0g8n/sZLA
nj/mPnFsMi+B3iBFyQcsIgHyHfv3CeH6BdAyJ8D3xk3+m/P2SyZRJeLoNzJ7OOsm
B5edAub1mexq8S5aiuAUvH1/cCFAgNzlFKh0zxDdzR3ln0l6utLKi9xuZOd6dIai
0naSdaL0SgXyTcWqnB1tHFrb8DXHiuLj+Qzs8FykoqUpKId1DRt0E4Q5uWNBsb4M
Oy0t5/bhOnyZzOjqeKJ9vB+AKITacfN9Csz3Qsxe/a7XJbo9Wrr2qzqn/ByakPDq
lFFKBuFusAhqKcTCSTcBg11O9JMUzzibM5xPupN6Fr/5QKvFQeGIpoJFRu5ugK5U
xcOTASQ7hVma00SuPnTq9gSgRwUse1hbCV86H2cVV8FI9If2k/Pki/wkSXGK/AcK
zg2B8Qjb8InVaI1gv0l0wyimeE/Ne9lzuldJ6lLMGjpUITN/QPP0w5NZ4coZ2jMl
05JBzI8eVx1EhbgQ5avfSd5paiPpxRwDvtYvKIvE6aHZPVq9xYSwt+Uk23rQlPAS
J6hm45TvR/FPrzuxFFT5OLADVkIqqVBFOxjTW/Yt0a02Hz4J5Y+6kOZdhVuqLV5v
jIgjn8sSJzrTkjqvmaCR6KNdwrMOi2wT1FaQJZ4FbmiF1QoHSxywzDLaD+/ldVMA
rmqPx8B+JCqPBqjn/+JhE8ZuwCRGZJVqq2hiZXICcHynRyhr2UjWFetUTKG6jrQX
WPIZTXDu1EuGIhK+3ydalyKeDKSAmnbxBViUW/N3eBFQ29so1lHvAvTxKlzoF2BN
3E/8bjUIeS4bAi7RP0B0W6QXs+329Jhl8lDRmLo3RE6FEn96ZNhCADzMMkKhE5QN
cft1tNGTf4XjNxQyr4k2Vpmky7Sd4AnwevlawuwUxBqJzHM8gFpfv6Kc6XHVkYCd
4vsYnbSa3EbSkiLhJaIpDfzhIYA8MKXPH77wVaiBz7xTBS1gIOIrxq+/ESxHAvrB
2mpDkJZIOhcFgXQQnBZsGbJnd9R3IcXRCMAiIQMyLTP27tOlnqqNIVWV/RC4Npdp
Zgm/IEkKpH0NDMTm2F4/ISeqNYRDZZG8BIrLeiTnPte61Yyh3srjAmgaCvAmqL5L
rgX18d1yHpCzEzr96ykE7d/duN7bukxNoB+Qxm8kro5q0M8qlEbrCbAF47ErVfyl
YLux/oUv1fwG5Eh1mha1FrAo6rWhmLTNppwkmQg7X9SiUHFM+Qc+Ud2dWEGejqUe
WO5PRum89hk+wv4mrg021JYtbxzg2yQLyrGslZL9AOaXzPzw1n2Bnd3NQbbB33Sv
S9HRfOMnrsLgmQDtaHUYvUkynIal7NHrYDEE6ODk9dGiyMQ2p840I+pr8fSQ2Vpl
InlZjaLDakpTnahcfrA64X1tIFVu6udoaHmvGpYa6fGSVaN/OLTWnCq45RAVAU58
nJixpGXrRfzQNeolsIOjbpUKjFWruI2+7HrlbnUKmjQY1zNuVhWwAk1BsnsJ03Ag
QKJUeBB1O+Y8nAGCY6Hwq7GlPPElYh5R4FG0MRqpC9SddTIlZPmN76xfYR8ezSaR
5HxLYoL5d6QwG4AonrrXY4YNzpJJc9n09ZAa5CSqNar1vEE5YODm9YNSbvYseSUi
2IBGfMZQZTZxNVoXyYZ2j4MmEs+zEGXlCyCBRhChaYkoPfoXLRNRLTi5XKz+/mhQ
kVlmgQvEuYNoKD2zz5TNdVSARfDR0Xuc4tckA3o7NIHUUMAO64w52YV/TrIGj7IQ
v/uw3WNimIcsMZ6BVVB5FhVnCP5qluFjdNPLT7VfJX6A403JDctEnEaCIeLlfbhT
ppzp0vLkY/AkEJa7orzorp78LvkGnyr9rdmEkkC9PPjo2lB4e3zeMmZhk70mglW4
2/ywIgeUHHkFBWnfPbdX1TbioXGev6j7vhvoWl+CBIS7FMob1POcyOooNm/4pX9f
+108MHepDuzIXMEH3l0wSs/4sboGUJK+94wdK0pkslpf/Gd9W1bttbyLaQgw81Oc
0lw92fruttuiTtHdlqNZcBynGwKuzisbPgQO3GWtL8lcT+ELO0SOP6C+D+JZRA3J
CIejpzSFEJhpjYydcoYuW+4IjgM5cvp0yJA8c6XEB/9oTsMc46PwC1s/iQy8/HjF
FYd66lhaUkChACOa6ADFqnG1SXIchsA0rjn2vvPEHNNfUcFmR8nf7SK/ea53CkSg
9GAp7JVaLuR7srboCx6fejvxFDO+152udPqgVMXLdr3bquEpiYEXzdTc3Xnh1rs1
SqNyXbwexnn4i9XuerzZ+gXsDTbiBUJmaPj5aSZqVg7LUR8RrMPx8MouzBDuPY3y
JjfTr7diSrcOpXdkxdew3TrixjLskLEqs0vsaWn4WpfiVgZ8tbViGBHBRaacinDk
1JQUeufGI+ROB5Rw6+6g0wZaZ6e6MXQgHUKvUIrZEeln1qWvy3CiTff8zuRuWuVy
qNAKiXJwKCuBh2PZuGaNopEV1W+bNa3ljKVWdfIX+zHN36+enj2HCkIGZYRnbMap
CGuTkotdhiNFAjMY8LxPqByFUCm07ADg+j8MwuoSCC74mUrgFfhFNzVN9b69Yjkp
cPr2zvhlhIfxswOpg4PHH8dqXPn2v/kCDUSglaqIH4AyN0zePN7k9BKcbi04Ej68
wXhNr/j2xlH9jIo1d1023lpLeTBmUR1JsW1wgvshSc3rqdazVorcKBTEdTFJMlhc
xQwfeXE1d5CwjOr7EgJSPYkdd/OyDSWiL75p518iYc9J+ZoSKlH5zEiUCPU663RY
VQKcihfUvvNI8qnFLKNAD+vNeAcWbZNL7BMw8abifpwdlj+CtKXVlawLcerYLmzc
F9/dJCE9BdZ+7gIET0B+QSbnqdIyq1mGEtZfLkZ060O6jxWtGPb1JkiCZ3bNMxxJ
XGv+KvFol+w1sqrYrVjbtxH/hGWTsWuKmAt6bhTrqIF/1qPwByyf6qSA6XrzGaVA
to4NDsnvcUB14y9KjMs2iSz6wii1b/Bx33R0FvZsFMeDPEqe2SMw4o1LhxSOoARf
dY3h9hpvn1mOWVZVH8uBRm4TnnL6m16bUQF0bQQczMZbhZ7wpS1sx4i1ymSWcmNj
59wGgYTGSsO46SlzHjx+OZvzT0q6y+7XwKc8NO4Lwcr34INFKdcq3JkBKzkQo1eN
sxu1ks8ioA2rhM4MpvKC6eg+vWEZYU+QbacVsJX5LA8pXWdh+evG8WuJ0I7vyZhY
JRE2X/GcZ+5DhLxE+OXsc5QJ8V0TVeh2Fb7jTT/0XSuS6iIV/PGPmk9900Smii54
0dOntzERkEsLnCrIMq8WasvIxWVihD8en2RBjQrvgWd8rTuhw+IfvlZhKaSuyLrL
WVC3WuFZOKDdQuVwI6MVQa0cp3BEZmPH23PdvN4AWklQu7wkP7gDTRYDuMbbiu/b
akXboREudKDQTt9GZonRcFaM8PEIi5isPRVYT9X2RFpfxFP8eBu1vGT6kYwK9w8X
NzKxY3mcsi1hcBIzzALht6WucQ9miG086UWyvoe654o6ixTOa4AGf6PFIEKlm57x
PHfs7VCetBMDcDTwy4IpbFIiqF9Tab+4KXL9HmB55QNo5opBtSS1QS2EdknTV/Pd
q1XjKutZUNHmJdX7PqcvtG5xnylr05DvrQgySvf7YgzQ8wWOsfnLE2cBpmcxruR9
T5rtVTlZvx09fdory+T4JxZ/xBS06HGnqOikfWxJn4LOeCjnFe/Ug9OmKgIVSgd9
jdFTvuVhugPrreTgmmGusYvX+JSqJ9w1HR0285kgm7kScScPzEJSmHlnnIibRuHM
fTWruTdHJZR1UBbYAknEvBy8bp8Ye5+hm+h8u1C1DPnxWbYmephdQYyBJpdXwsGs
bhQCFdCfxBjcP3tHjGO02bSE+DuXfhhvOhUPpHASpwXGxFgyc5DL3/Hf3bGQ6wXq
ZfxuuoFv5F4ipbVXm4i5GyedCC0VLakXGEvcKhpUmsf5fikXcIuxHCOC3id9G5lG
YENkgW4DJRb3WpQmoxB7ckT6Rpfr1bqR3G+b1WA5DnlvjOtXwGf5H4WkoKm3q4ES
ESB0Pf0c549wN4dLWiO1j9EuPSxF4EJxrQ5MtO9KvxEUUXXp/hTIq4WZjr9UTMEu
4+SmVTo7fG0lYxCujs5ETFUEf+Qf41Hvjl79To59P41gic8DY3Y0nhvjXmKzgbQI
dg55+9cCYckD8J3TlG4t/80vKPJPWdKsNP+ZceMmsdu1XAlqSbOmsIrCpOwkdoZb
TXpahEbljHPABLGuIfHjaq67eP+9t4Xf9N+gBWYNsEcfVpMsjAZw5lbleqMuyBHX
TuPZDyqv8dR+dY+g8x3ZIwhbGQ1w8avbI3XwGEHoLak6btc8AbAq1kiYHjdhoEnw
lqdta+jNvuGwhJ+FSiV/sbZK5pwUGzhRmIAMJA3uSiqw56UGZq+hD87+dT4xXh8I
P9US3sYxAxJ4ZfH2/iHUKvP8bgoxx1IW80SpDesMICHdwsiCn1lRyOlyl2ZfxPtY
wYoYqt9G0cs0jO79lCvXQ9+uMM7xzcG6bqbzLyYMXQfDNOrwo3/klYRhlibZw64t
M7NRw6HjR8TcUGZzj3JjfAUX3CY4nxRihm2MbgSLa5g=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
U956RWYAGleJiinRg2YqEK9sM3etXQMXlRhgNM4Y9gmcBUkfsRgtuz2xsxmUoOzl
islNQPcFOUo0OEQidXVoO6QYyGiqenSRvLPFyHIknwNBi3YYY3xhcDC08JaqKy1g
qVT4phfkObENzrz1BcgFMi16pCSDAU1JqSZ4VoZgcTHrpuHJsg0SX06Jt6EsKEz4
fAZNVo5X2q0UIYGbaHLZK9VjQmwRy7apf0VY5clUQSqnQu31EG0UQCghgsK4ZQdR
9heW/OtryzXPT+Ao9cnjmMCcyKSgcpxquCGPHUVGt3zSkMSJvIv7To2iMh7nW7Gm
3fVFFdGtVkL9cP0bIUO7Qw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4192 )
`pragma protect data_block
nfIPvVfRUAoi71yQoLEE9DeIkihF6z7df4CbnB1ID+EmTFTwL9e74VK0nqJyKkk2
JfO645i7VwEkvgcPkYGy3XDa1ilDMEDmu86aLU6JoONwfRlZnQ0+e21eUOTyR6yI
aZ5DoxFwVcYUdOa1g5lDfjy5tYtz1hcDf0uk7z22KzI8q9brBSSRp946eiECvrZX
JChugpilXsNKLQoxkYtXQutQOUz2I0tBR2UDhxtI/uPF12EpZZ2jlDlILncWlr7q
ow30XbpaH3rUr99FUZLRoIOoD3e6R3m1e2uBHsK+CQRyjZP83po015l4xt4PoAxH
94KbB3mhajK4pMcJihbUm/Vp6lb3bquJJLuueuHSdmaAcCO11YeBFS6DQ9QkjBud
qs/PuLma7emddS2DvgwhUg5cZYCDRk565E8DnJk6fH1sKRgVIvUPU95v+mfArkQl
dsqy8nHbtHTAXGIeW4bgqnYL6hAZK0qOBtXtKchQN4mCU5kuSFe8hiUUMMMb3xEQ
Q/Qflt8yay5EOh8X+9H76hWzvAtLH1MX9wgtg8+spiEfBLpNt/NS5i28wOxvJIOk
HX7OSkiWcZdOl3/0iynU2LzWwBHiosYjaCpFjELp6WL4Y1GMZd7+w2NIpwoabSUS
zmalpxo6N2WfcFcL4JrA0CAgpfAQFYa1CW1GcUAsKEAd9EtHxPJVGXC5Uv4qjiXH
DNROMSIiFDAW1H8tybC1xaY+8G+SEm+ZVzInyRymTnp7LVdtc4cpnh/bsGglPMHZ
CxRDuFsNJtoDgWPodNrRh1QmBqRPI5vFNuymva8BegbOCuW+zTYyO+FA7+eu7o0r
12Wq/3qTHbc/07WIKRlincdaWJnhfYrnYhGW/qpBfRt67PF58BhDZIUTwFivofHE
GcetRftaXGlS0xAXegX4ZNHSUEoakzrA1d1RkGHrfySQ19UNli5MIrBz7+TkT1iR
5MleLTzmmscCT86EiwA8AYJ2CDIqfxF/nGgucRKu1aW6gp7IZVig6Aloi9+To6Ag
nX3KMozrGdGtOpnvinBHzDcmy/SzFlyPSopl1BYsNfFjuOQ4GmGAb0bEvyFgnAHS
IHzXvwqUSw0R5MJE6BLkqxWZ7o5kZ6Ne48FKLyHcQVwjYDwBU+a5/Ai8Dy0nYQQc
MvmsmA7l5Y/Vx8sDg6jMAF1ceDirz1k0Gcho4Htee6fw6olx+0D/fO3q2zGzvabG
MOS2xmsO2JRwWGAJo9lELKDn/SY2ADDlrirTnxmeFKcxDiKgWVDDx7DoITgzht50
YjTemmEAcxLvuRCzGh2n1xGdXxUeNjVeIiUL+vmL2ltWIdQD2iFJp6Jceef2bACX
zPZMtMMtdwXW/oFGKy1P6hx03DNd1wnjqqGPu0ZBWlXFVGJ/4dvJ/9889ugvNwGI
NVB6l5oLqL/sBmbFvqQTzRC1fa0UY2X7bT6uAdm1zNQyMwINpGIMZU8bHSxB9qHt
NWnWMOyjHer0ukohITuUb3mIbzaxWA44nUrN5Nl6mZoQRm0fu/53H34DeZCXyvxJ
C0NtFzoA4JqfY/N4IXoVQs1crDHZnK1TaanTDsC3S3JGQX2hXp08Xd/1k2hEwD/A
k0mPKglIKdyF71d0rmg9ubdWeHGrkRtuoZSovvhfr9xyT+qqTenVDkhr5jyd4cx9
dOw933byeI/E2fu2oRka3K5wop6/moj2Rt/+XHrrcubJwXsCKpiYdRPIae5gvIEz
SApIkZ+LGE87bP5ZEMY540TabwkorjIJ+vIK+x0/OrAk+ZSePNZe+Kl4fPMlnf1m
uTKzOc394LEIGOX+Nwz86KiPMsL6Uhq7kqnwBj42VGkWwvShpBwbmuy1LXCp5dxj
NAFlegfsy6UC/h3plb72Xzbl8fUeW6M9vIB07xqwx+Fn84L9ulBPbij59uePCdtn
58QepRLKgZ0LYtKn7p2sJbCNTMLeK4+Py85y7mAXbxWQ6320tcySO8vjk2VJ8h7k
kh4o+dGOFCKs/49NQ1sY1AwlT8dS+0I0R69GpIj//Y6ZXZCNFy3zvq6PUWvOkvWD
sIk55u5Pvf56FtUKFT69sQ0No+2e8wkrbJ5q8o+bhO6pkF6FMaLJbUXa2/ccqada
f+C4qII6iKVPFE8GqLfNl7TJ5gBK4PkOF7hM0JCxkMQ/1OCeCET/wmoRXD4B+pZf
VafxgPgxmRlzEnv//zhHnMHZEbiEkA6TTQjHjMSZyV/Jh7B13dnBcVnvzZeLo4Z4
shaY806mnKon8M+WaLhNXx5T01j9vOSmIO2Nh0DuF4pEDxaW3P2+FFMWq0FVDx3j
T83RhsbSWbkLoA8tM/Fc+LVWhBKnF2XSUHbajGdeMssEL73M+kXTn2i6HXSrnhtu
fsNwHUL1kejR2xcTcgEL9lI3bALQpqEfIzqVzQnFFjb+ZNgSj/KTV2ASTeI1olk+
OpBeeg2rUrkUiwTqvIrsdqm09g/ULqfxnVulD3BsRvzRSaHPG8dgd+4HwbeHqzP3
sy/nfUHuYF//PqRp67sjgTeNkd/pIJELzUGdvZltjRvBnnI/Q4LlnjTtX/mpTJMU
sXpVict8IJsNdKi9UHlyXbQjMlAG7iDPA824nYipMXp65yh9WxOX588qmWqaMCht
9OaH+OTmiy+X9Q6CNHCxo5ygk02A5EuNmdrOqCb+hP1vBsDmvdzwZgbtkjv+Yri0
vh40wgHwFrTPvUVQPdAFjBeBfqAmHaFOeQ9+hSPd0+zTu66IpBJteih4CLJIrTG8
mzMIJHny5Wm1eTIchFGaF79PrTkQuW1zuPydxmPfwjHDwkSdglN3yl0UOLgPSSNv
u9c+oDHRZsBivIo7KbfCvqvIGowsmcr/iKauYV7gcLXirtTiBMQFRp2NYX03EoEg
VttJdN+RCewOx6APlFl+3hgVs2usPf2HdCdTekUDjH7TZwxhnyRDWbtZ+6nLCYUw
6blwZwKq4ouQDok9R5mzsu+AN2HmSZiHvoWz5zaIWSo9w37YFPu2jc4rePQzal6F
gRVEcV5HNR5nN7lvFZM/7zwkkh2xCKCrXubmprcfuJ8InCXMK2Swc5g+lQEh3nTd
vGBRy8oz+3alkOqu3HoGEtXNJNqhhoxjckL1/A1OjKp1rAGFjyXoe7ANbp/Gkozi
5UuD0xv5RFvYmj0OrYzMMx23AVQwUJgnf4t9N8LtAQacV5ss8o9F/Ndj1b8bTlNM
tc+ix+C45cgNDvYruixFcU0FTxv+FPmuNDw0RNWo3rpS5KaGm4AbvTXqv48/EYLO
c5l+AjvscjaRMfay7R/+4d9qkZJ1YwhO1vnxd+PvxYhINCIjMr1NUfTWgJWk5VPg
lDvm1F7R0YOouP95WlL9Jymqra7sVpdD/ztcST77y38y3LhsmjfxyvXVt1acAh2f
WUXac696XSQ7jMvvm2dcQaGczh+t5wO74JfHWkIWxjeCa4x0xxQ6L7/K4VzG3s7c
0erd5skYTOe4b0YcdHAnF1qrpFhRxJntvLuipV1Ks49cvo3CvATVkj0FqeyLv2is
3Omq3xeP9Z5DjjQO1v3raI8fFGlsjnl3c03Ymx9INDYp/6UNHPuHDg/+UshfI6Ao
YB78TNvRU8NuO7EqmgL+Cpii4TM8Q8+nIgN8iWjt5s6jVZO8QNSeqbWabwL4YcuY
Hx8ckrpFzKJQKC9nd+9V/7PTAmeIaCUWE+4iemcEe5LyJ+cu62m0rJk5iKCrfA7+
Savfkhryz/tkKuJxqC9YMq/fVkMtEyzOEEM9O88bbUKUfxyDUmukauqqJC3PLVeR
gaDk8/s5L1LuaXMi6cElooTA6/ZSdA/3G3VcUoYrD8VM8wJGqiole9IjbqBoKNRZ
QcKhoT9EAGE4u9+7QehcAoS4i9IwWJTEk83w1OE03Xn6A9/YATgyMaYwxmirtXaz
BONtkskGGL42p++d+IwkjnD9tKSefvLGVqNwp6zkcJD1vw4VDBo+s/JHtiQ56xxC
GsbYD71/aOHfo6M9aHDpBjuG+/5U1dbJRSITyhHNXBdhvyfhV6OCmCWMkDoM7rzg
bYEMWSoSI1Ec7zn9PAjJ4O5KOmv68VG2cvMsNmTV0JjW8kINGCqafYm26l+8J3gI
zP5trpejICPkwcgpTeRKkPdO/aU/Dl2v64AOeEofKKrO4fpDbMqfgujyhyN2xDJy
f+jNu1j6RrTgyo+5T15RLav+/CKsUM6/VjgOzsOBQ6ISaQQdKgWZCN7fcFsj8MWI
w8SvLAYpHWpGUVX4lx7loEm/OLBSWYwAm6usYl9c2jp7msE0cUFIw2DCmf061sgz
obkMobzqeQoXqp0OROMAiODo8lRz+dJ5NHpKAL3RgViX3Af6plj+k7B2///564cp
JKck+vwksDcxTY4g/B/rAI7oi0r2fx6/WINV840py38usvejACHwmrSx/VXAMajG
cLf8/Vsm1lUCBpW11AYWi3ffz6iPhwloGY3P+PvoeiOvKfeAFaSG7CZ17bwQqnAZ
QIwLDYgDvM/GE8UPz/8dPd5l5evv0H2DAngC5nNmqBtekRkL5TyIDQDk0rNC9BQg
0EMcFVSLxf7z69sOM171Ey23VNcWIn/vzC6/pfzsYyKq04et1cRf8J40qYSCtvMJ
rnIacNRWTCcKrd8MYCp4Zetwk8khvWaTibt8TwtAu0/duTqTs4i2gNx43CUJf/C8
YLNlGkbnYYt3tdwTbZV9V/UwKZxr6EPIAH+elbOIW8uGvWOlCWG9OhMzOWC3dFgd
dFqW1PLfBL/TN6zcYChMytty2clSzIXUBMKchuimDjzAJYecynRBlUb+/GdLQsFJ
wWOTLPBcSrlRG1XZAfpFGua1MIB+OJHR1bRMzQQfUTwp8gBzbor2ODbj0uKjYH4a
kfhTm/qqsLm2BINE2VlcfLqu+VH4470M+9bhpEOj/R8bHs2ICEWOICCk0Kx6nWUl
dAbJUubQDIs9Dp5GEdoHzhtNMlN+EL7emDI/jVaKLfkkUaS2p/0XLUpOa8ycPzor
XvgXt0dH0D7kLuSZx4NPdMou/rtjcZnpsBeavTwNEsu/ou2HDrsuSoOa0uks4I+7
oSyOAIcpqZp2ZlGxT0qKi8ve361fgrXatkgJXBH7hJG/24om0i2tr/Qu82WVSGyX
3IUrNEwNTDWHIw0HzW2LSgPABNDl1tqMSqYmgumbsdFx65ckZQSzcgESBbFtZwRW
VOMQ8Kx+7zFyrCa2LfRGUHdsHsGIKGMSDj3N6Hrs4ltUAaHF5PrS5UmXRo/35+6f
P1XIULBpQw4J76oLRapG+lG1KM03Sd2NykQgUk56Neba3pQcZNWJHoEnFQfTWjEG
6RbwrQLopB2iMdClE1MMDlrOqLo50TsZxgEG+70ALMOjaHemSaOLtF+v7OCI0RS9
uq6IERfJX20htQN/MwZRqlW1LboYGQO34unWvt6wo1v+7Yhi3gchPUps7NEC8p7s
C+N4/7lfOj2J4kn/zVNMaweB8cNVBAUEV1RyxOfydbynlIHmIniRv8g/MpN7g8Tr
92NkVGtc0Z/ib7hlpETdmB3eWgww/JlDX4AOixGU616HYVpe1b5h9oxXoeOk/HVT
7prsEdCTz0g04PndCNYEvg==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BYLg3Pf1WUg8/GOiSwvENvm7TyxR454nTAwhVqpiMruor8gEI7rf1dux3yK1oZ7F
RwUGM3rrQwr7HmZBP+9yZHEtjmbrvCLR3LPce0PXJ787y1lZIAvq/56UHzV+gFMj
LleSK7m6AxAOF+hACEGXfuo/12acSiKiB7s8WFL5qXJFwFka6Ok/SEq52IkQWwMk
Vk/IO950/Mlap783HoG8kxHnHGDUOOCifNdoh02HbJKFNLwbE8RRS2Ye+DJsGBp3
6mLiP4KuzoctpLLPS39vuH7Rjtq14+zM+Wv+vPbENov2Hi7CRuqBWinTSJwi9R6h
oFehpW612Q0IlmTQMACUMw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
C/6Q4stsKuD29NeC2pMVWOFVhdtwUEpHHJtob0oMwccOBXJxAC8m8p0Y+0yYdV5b
e1s4uXxLPsyeDP198ifrBDEHf+FhEsxnmOTDTZrAGitVdiC4lHsrRN+QQwqIuzRF
gxY0ZRFgTEtvl6rrDZz0JCPhA2zC5mHBjDzHiNC5qBjT9X2o4IbNDw8dcgYq86TF
UihnN8sePE08eJEZXuCoRn0UgJEePHi/c9PVKO0wbmA3sP7VVB6+Yd1Ds3X04KfQ
B4i4RyWZvplBioULwkn0laMhsxaJhqswRFXNUGuVNwedtOaJuZaymBsbNNfjX2y8
AG3rFERHPcTTHG+csm6xUYqsojmUysYCBbMoFbktNl+u6yhJh3WFen3Athb7D0Eq
XlCHKt9CMcb8SqONi00IqSKeAKStfwAMyz32EzZBG8GxOgBVgTCYQ2cRi+TVpFwV
i3cQwYX+ECegkIefUAgZvjl82yU3UyBzfNeSm6Y9SrkvYYANkXm2p+o4MQ0E79Rd
GdpDI8TpFx7vqdhnJczgXN1gDhFQ9YBsI7slMDk1IE/GQRj+Z2I9FlpM0sCCBqry
YHVLqritqliZBAXRy9BPSO9nLEkY0w2Zgkr1dH9id1yNOd2c4/IsOe2Toq4fIbwK
no+/KL1Qati+hGhmxrRle3FlPvJVyABOjBooz7GgsA9Eoa1GkgJ/TmmC+LjzUnVc
1Up+zl0Kwmz/FelQjgNeNWJBBemEd15GkcVZHpYBsO7ksvqw6TgSvwlqrfHmD08u
bQlXnchSlFXnLOaXk/jcWV3EO4nVyQ1fQ2voS9W+A+zastQt6iij7mjKzFuJ8AhU
v319VOEk6Z5L08QJR1CQE6SRjY0ifpv5KneULcAh50MMfQzlV+35YZKsQu6jFacD
67FEzxeHbHq4v4Jx5T+QChB0bVIWma3mcXAEDsUXt5nwSckM4zffvS1WV4v/DJSl
utmlrP85Us13gVDyEW9UjvPt3hMia+CZUnSRurgTc13anYxxB8jvF53ynyXJaVrL
0hj6n5uoW0ZkdwRxlT+5y4+B6Z4IP+9vszztWXCwB2MKSiydVHuIGOifCkxvWj4K
N9nTI50k/byJuvduTB/b/uAGzGI4fxcbUf627BCJqXh0Q6x4gp8knPx6XmE6PLyf
BvIcuQAoGE/Z2hWXIixN/eBSs9SAFRDh+Fmqe6rsdfuh9Word6TlPRON+Yz4mE3a
GjCIyrRLvsStPK5+7ebMrJCEsKjppsWy6i6FsAu0DMb7T1UcyKq2L5WYGfqmr+6b
1MHt8eK1v8XRPIdl8ZfdvQ0Wg6qHUiaIoeoS4THxGdQDeF+g4FEwS9B/WiTb5PI4
XwQgAM3/Me+8JuWCdt+IpIhhjbXzZSda0vU0wy236X6/gm8iPJp8y5imxwJrdP8W
3Lq1FPkFJMA4X6swxT3Y5CB3+QK44ZNuICG+1ijt8218LkAKpzw9QVTxhU0zwSIM
hrgIPSnY3UDFNOFq4PGbKnzrHnJP3Fr1suj/qOskYMdnpsvkJ2s7sIqeP0Zgs6o7
D2VKAu8O+FW5zUizVmjOeTutLNkjvT+olSf2dTvtlyPakOtodVmtJVJy+aZ2srYC
FG4cWqTKoxst0NHWSpi5hd4pxe7RRaWEqvreNtzGo5P8ds4QZ48FQ4mAokFHn1QW
S8jlWE0YdplniQldZG6a+bKcisqd8znLXlrbM0FOk0lcezuDMbG1lT4GkeS7P8Nk
/PeHTj4uf9YNlTLr5I7TIAqjTPkPf3ygAi3TL18T7UpsM6xWD+b1Ao5vmkKkZdKL
0jpP5TsmAVHrtTe005wRzCNRDBnVse0kJS3lFZOeKB+n/ORJWADTSp8lazv8bUCF
3Gtvy3X8iklY6h9/1iEoDiegQvjUjoYMnX8G/d52SMJT1PWoiKew4Iafvjmv87Uu
Sj2MrFPzF1zMbS76+/HcZIuyIxqQspBw+VLzPtL1kE1bIGXrO8vrlkjZP0cX/XRS
TznYct5SoD2N+Y66y0akjrTPmLvsXN/7k1WhhYWgl0ktkdd6FArqFecgCd8awWRV
lP+v2SJptIbErcJ/D/unrBZzIPhSWTZNpgf+C5ZxKK6nWZsON3z2q+HNvDqqpOaH
Dzb2pf9E5K6cParO3cbSPiWkS3j5u17VwD0FVxhhxCgMV5N0dQ+IBQDOn8b3aWjX
kRwDPaQYv9pOj9vOIcaelOdHbgqYIP5B4o2GGtiKFI9pGxW4GEMzouKzygY51aJ2
DX/FclhbSMgXvNx1z1ZllQWBsMCt3iacmXs8ZeEiMj+4Irjs9p84EezPb0173IJJ
FICW+76tmS45DO/pI2zjPV/NhDXTAJf8tOtVAdhS2i7rFnmecCSGiYSi1P32flwH
HK4zALtOWpEqBQ3cLw1BolvkbOSuv+qC9wySIIox/oY4JRGGta5IGQHKWGSmjYdM
d275aKFGtU18skoN+j0Uub/YH8huATy4phxtPe859eX7Hmm9neuiDjm4ui00ex1k
yk/sJKZZtYY11XfH07r2Uoeb0OSYM4XTVXq6LxVakr1ZNci7Umoa/yCbvkyNiLCd
j/zIXOcB2y7VDSy77AqPjcYyjtVfDVLutfSdV8CvSP0A5BEB3IcUFgYOYUJI6BfQ
qyl3Qygb6VRFzht0pSt9MFYxTCGJQBLB4YTWzBikPOw9XJ625j8v+/dOgDpbd8vp
M9Fo4lUar76AHtkfvc0+QlbtmaVhJ9zlELA/cgniSVe3UDC58pkbn5bHgYNI/Bdu
TMNbCgQcyNOAGxdTZiXgSD5euBt8vR+OAkoQS2he6ogJLkogmV/jElqYDl+HbU2C
F+rC/F0N/A8z/BgMCITD3JDpdh3aFQUTsY1+b3rVEhTD+H2TUbYpYWkYacguIG0t
iDJXcos2FhfeWlXRuw/H5UEKopa7BJbxRdp0KrxQIzvoRucq5gdzMN28GlK678+z
zCez9ho7n+rRSbMCIR4sT79rDVr+sTnCg/LjfmUZ+oVRfaol8LQmSSK0JVeiNhNw
bTmGTduPpzURacRf53nJJLis9gPU0eAsigV337d+5cQGpnqSSEt3hqKFgwmhJvS6
9piSGR6w4jOmMHb6q3/jzL/Zg2H53J9dzA6edVuR9S83ax6+BNczJRNh5n1MCt/T
nlh8bk/NhoY058JDYKurPr1pUIvibuqWdAOALh8t8T3egu3G6IFsVHW1h4BLER3w
Obv2fY1i82Ski21vqyaDMvCmBfW/8tZdCqwg8KaG56efuA3ca8A3GR8ct3Mawmxz
gluSminSlGeMyTI3UY4VDbFJ8J9JYtiOf3x+7/lFFO93UY/6gU9oZ9kjK5M2iC8z
CZKzlYQNV2/zBzpbmYxtVeV0y7bC0h4z4wtoAUI6uCyl3uCBClm0SVFfRzXWa6CM
Php24uAV7iC9mlvXwnZeJX5Bp/gs1AFOeXGnzJMzhhh9SvkAfmRSss8E9Mx4JUD4
WozLtr73uw87qwOybuZaOgcwGzkYXQ8ZddSu3gd6p393wtG++HJWMgyUFkZZXXVs
Z8HULn7XpU5QpKqqSKnXdsEb0dKEkhGpUPIlLlzAEwBDYSj4l9YUcwhDUdgnrViP
uRgA5ok649mkRy5RMtZsDM/hcBwWYg7krm6nHJfHrRKAyp3BqbEU/vKj9OT79CRq
Fvfi63Tp5XlWVGvZvTWAefejWEqcJsyVsCuM2CrnYxvnrKm1Q2Wdj4fMuXss359p
LfZ8XdfbRMvlJ5KMscv12Qn6r0oCnbCY5u58FswhMnAyvepewZ3qwcoXZIi2XrtH
AOAW8xXV0HPM0xbmD9udPR4aLfROyF91jCJ1e/Y9Ug7CJkXPPExnVI4lhzrvmjR4
XHysY1/AFYAtRPwEd8Isjl4EOxpzCH42fILc0MtwaH28raf7Kq9Ig+RGrLStoNVb
f3nnCZ5r+FixRLz5SUeg+ALSpyR1T/xxtUYNUx2luB2bNlhxxyDTQKlTcvWmIuwI
biLUr1AJaPhz4utP5LbFwziAhWAxp2zPkmc3M3kZYXUQOpdwhiq/70vkbzk3j9Ni
+gcNGSpaJb4YbCFIa3vLi9GOKl2ryJYhBhoSOPQBOozNjhU+qP82eUkVwa7aXE+t
3S1cqY1KuTzgA7mTHMnGrXY8UK9RMr7jIOIdDQBzjvPyyCKk78JnvuZOsY3h3RfR
4BTriPmu3a0xNqbWHjJOkYR165jpvfKWyHLALzGb4TBZm6lcnmKrSQLJqvWVlgcz
w29vtJFhJQB1bVupXO7FuX7ErrJlURdtaJwwaII98G2KIjrftU11m5Yq4c5c9NgR
oXz7/CZDbpnIiWqyjrCLjwai7m/IOBv2sCjYsBIxattBZqYOk9A2JUvzOIQMgG1H
pdL8Cr3g+CDOChUJl9+hh7lRoZUhm9CgUl6vSMrZTSLn4JWeTNICuVlvvHCJ1dbA
9SdBmG9n2QPANIrY23jHMdYGtH/10wwJiUu/YDhP6EpNXjtqk3UHjsgvkTQB055d
FlBEpZHRfVodwOjF8q/BRRzx9kZpMdP8zvXf62exdGIvlqjXXneAsGyhY2VgX8yd
ufXeqzCHBG2O55x7DVUbOK4kjHDTkUI5CszUmse1GXzgTdf6foR5N+5LH9DcmkKx
/U93yvdNeOc8wiaY5ffHOACzvCFWsBUKE4e1krhVXNoSdRXsHHYxL/Em5o7xtlUb
PfnJvXXyXEnjDwwYEP99saFbIgwPtG4Beprwx8YmUwN86rf3hb7ZSLsaTHha2ms4
m4eT0wQSL051lvNGultfmpLbibPBxe6j+ILIKLuXcRvvG4PmUA09u0VlpeAm1iAw
uesMrvWalQJQ0O8+9cLVIUOorwwAAZ377eh8avCicdZuM38flZ8Say3Tedf3wivC
gxBkaW3O0DKW7zAk+2fuDx2H0XXqghzbCvOSamxkkNCQVZfVZcOlRz/MNsUtUYG4
mkZK6n61l99srIZ0iSwcE4kXILnVlWmlHbQahLQAWJ93kyRJnk9NrdNRaWRsfUmw
nz8B2XPRxz+KXW+xqVwvWYU9KSgqaVW14fySSu4gDFjPgBkCxA7LIEJn+BE9hLUX
snKxWORsSbYpzN4stjLa47iwd0L/8uggSTobo80owTx73Zk+6Ama5rhV+GxCVpm3
wzYSIy9tVNvZ1FVUnfYYu9T/xG3CIcuRAiyh7/l/W39ha7YwCq2W8cTZ5TsAkotW
uHbhTff+GD71c1symIbbetx0Jl10v0GNFknPGuUJuei+w67AzDanOZZFhNVyYIvu
mLT9B+Yth96WJ5GmLIHwD7/wJyEYKMZrpAUnWm8YcxsALvr89tRzT27tzews+cGA
3srPnqoLkjd6+tYX9udRwDM7qs1Y6VRBrPGB0hLwsgHSgAuTGzoyOQbdNys5Iz1l
7DBNwHKbFIKxgX53sYjg0/WUL86zZMGzB61cajTEQeV3l53lJ4NhRD5iPm2Q9lwT
r/fHyYPVyZQXnKr3IxQolBJSorf+fqM67+a2qocIcBHhDTkdDREBiIwpssJZVW49
Sk7fzyH/apS4FyOFAtuhEtAoKMJ1Cpin/Y2ztC8nh1DJftgg2CGcmO36Tp28J0uv
S0m2YU6mhTMCZTGi2dm5ErS8onBSutJOGGXB/77BFrnEje2vELW44tsyoqr6aUl+
SB1WFi+5TcrriniOmCHJ5KVojr0QYw0MI0Kc2pfzdrCvfzISy8coTGZgBCNtb9M3
+2ppUm3mQ4D1asFJgUcBw2Rbou/tsWz+r74YkYXgg8V6J2HDeFeKCX2CXy1H5vnj
lGgWk21bByNlB8KTlr7rNAWtXeLk/NmKf7vCweCZzdY+iHumZUnT1WW7iDv1Pfum
+FufC82f+GEShoiWJatK/j4SLPTBhKwzDapMgE42OF8n/5A9Mon5/TIc+D9ucEEu
NS8aZiVRqpvwQaXTncQ472L8Mw6jK1zk5gSP/Ak8I05Tsmu4NlZ+L9VkhhwpYff2
VT44hfPLVY/mVMegz3LVw7e6emem/MAJ0nK0Nbv/ZIoYieAC3xKs4ht/Ts5ETPyg
ZRcxI5oTZ+E9rvPKt6vkyanTmFe3zo1CUY7t5aBSdm+tk2jXl+mSfRAxspJJMkek
cX2lMZ6jW3kd5scGeJ3mA8UMcz5RTxXmthCniKdLyxbv/u+UjuUZ0FN3XDhF7vaZ
FMg0r8KPgDKXzbh10A4uqsi4BZNclBiKtqktJ4VcdXReg1rq7Hb3iVoXMpuU/dr7
1gL6GxQMTVMh3k1qD2ZbJDRS+bm7/i5UMqO3WcdpcysnCbCMWzJ50pRsDUpiCOOs
/LEM7X6LArXMqBAq5azdHR0ZNRAom72zrY7eN4XQbgHI1HjOuLRI6uBr4+pgtkUw
kfyeplNf/DDSG3TPP7LrK2FE5HGZyHVml66735jyix+zbGQ+jBEWcjCa4Djb9a0r
tpcNOUrAsX56tZ8abfWExEZtUrNcLIDCnyhGjHIUvaxURtyxP6Q6QHrncOKO+MeG
3/dSA/1pv/N/imLbVuBZvnOVx4B3vxzeRRXlR5XaY1gICjwFRLh0g0wdqeZiQTZB
u95gKhLFVxd2NcAzThUYaUNVN6E8IfZF+cOWrgWQezJYZZ2haCWvKjolhDg3VbKp
cMFtRvSCqfYEMIUd4g859DDlCpzEUHlW+wZQi/8rSlKB5Cpjia3cIdRmtxBtPk5t
Achv7hN+zqHzDUKR+m7oVigtIadzjU2tk/cFce6raO9GD8fz13cj+QgGqPhGXE7B
atoNhfMYlHAgMRPBWdFnTTe0uWb4k1g281SvdpRiOFpZG5tPWVADKsFRY/c5MAXy
uvWUQ28bmDlcucz8MD8O4AYNY+2MPlPgs1L88V1etUZgArOxNBQkUU3f8U6+FXWG
zX/jHuuf+RI4o0C4Sr7AHfxIiE/q5AUqAC//EMxGQS6FtzAdpNw2ll3emU4Rnr7J
+gaRAo8YNm5Zpxgc0Jm6IupOQkxmoz2vKyJil9wjYtz1b4QEH5tV8br47YR6hHH4
DRpCsxDgr0Cpvs53QpXMbCjlgoryiOTZaxX4Sbl49yWgAJrUz88r5kzxLo2374vH
FoGBdz2qkiLONmjuCxuKOkTIFYNnvH45H2RYDea2K6OXlF/tbi8AICxUzbQWUOFN
x9JyJKj4Zmy2Cqz1meK0gss0EKl53va4YXWL0qkgzWCpH0bbpCm6HOVSQo/GToPr
PG5Dqi/yCF69nL2pF68bBBtTsafxVpBkWULWetS9DLWtPVjM2BWBeQNugdS51X/y
5qhpMse+gjDFGKDLkDZTWGT6Sm6z0q+L8c7/5137XzSCGZ2ysytVOGv2hxs7Dlw0
XEDz8qH3J+By/UQyhavjnL7OS5tnlkgEkbubj70EU583GB/ezouEakOkXvr0px6/
OCXpEK+eM1ZfMsdnC0Ztrf5bcm+tj841KHCmOAU/SEtrtTp+Co4hkajYGDTw17ZO
8rhWway24dteOxfF9tWFE6m8/Ey4+U3M2csOiBrBTu/TrtV3eRRlMEZWopeA0pfe
h3IgHN9d4PUfKyHTZOjTzpAKQB6UZAd4l0wzdhLXjdlibNReuytj/4uE/xk+6C60
7yQI6VOG2SUGUTzVZOA7BEXjOVFDC01wuvPuQNw+eqUS+ztq+xO/nw6Ca+H7nUAN
ydLa8IPaw2IpTa2xAtg1uwJORQxNNT8aUKCecJOROHxRS1P5cn3uJodM8LuPetjp
U0FBtZPeYXEF0xecHd5+73Wqe1duYVd5h+mH22v2S+/Hot4BbMT6nEMIC4yOnmNB
9b93WJffOddLR/AhqaTpPKiqJyUJ8jVecJqQ8ze4cu+eznTq2szOYwrtbJ1V8l/P
yCGr0yQBkSu+3WKhgLaU73gNQ89Vfv7ElOcmTclNHiT5uZUTTu4HXlnhwsJwozpr
vOz24rIrt1bhi7z95551CQwofy8CWt9jvOasholYIgaY18EjjL0b5qh8I+ZjyUuV
qnJNblwCwdcEKMgjVsMYsDoCiAKUUxnVert8u5A1grrHOixgnDiynI54KjX4G/8/
2/3R16rSbOiSK27aofLQ7L7B22wxuXopoWLV/+Vx1KvNdl5XgwovwJ0jcc9Wr57i
GHZ3Ex/dDU8O351Claa1AfKBBotbDNEWrsTyxHa+rOypyci8G4kjjinSdqsk3mIt
fSojyrWTIx3cI5oMFW/d7dDiobUZD8PJL5tcBMxwAt8y4hhL+Wvm3Vp/QtL4p8iz
X7RSj1hTGgs9zjBm2ARxOHJb/JTaLup4rbDxPluTVxvqdQi8jVNkkqzD5dH2wv14
ikwcW7/tiVkrNqhZi3mF4wT2vDdskBCNGXLVlyraztbqmh65+P1FtW9//hbz9VhG
P4LeunXxex1kyJmKo0MLjbC0mTzqWm2qmRJbsQoLc42ywNaUpV9PdexV4uXjnMNQ
bJg9mdUnh8x6KguxtKVJSEP/faK2oGeGDdhQ9CRsFaudIL46k0hRwowIAyOD0o64
1lbkhqaunkX2OlPoU82Npc+rPjd2HIvJGjeFNH7RpjUPtE6w22ewnL6GVLskEK+y
hXANEiLfzF17CgNChg+D/e3b5VB1rshNeJwKq2/erpjA0NCa0mf0FlqqdkwvBhAi
ZChSfbUPXRLv5IzUtOU4WYMORDGkK2vQECy33DGti3ZnqNOjl1GAhqGR5SxuLRDz
i0uHE66Itpl1aGCY0MfeDt1eERCI5RWQOGQsXqm8UqjaqdYX5Hc/ib+I2f15BHll
jSqBZQwnjT8snasQCwu8s8cIC7VXxA4YmLPOGPEis6QOWUDe2sqJrmkqNVpVJPf8
qkBQmkNPHxNMzQHd3klhIiycnoYkIn0usWbdM4HUptqnCx8mrgZMC1Nzd+3pP+5a
E1IB3X5C+sc8wgjxFtvW7cC5NgB2o62YMzg/vaj3A3OvHAZ2LV58HXhYPivWYydm
VUcBQsbDCECbrxZ3Vr6jlJas67wmunGwW5g1a0suM8aLcphyoncbOAasDd7gdxE1
EKuSFVjrsFKsSsRLZToD9ZVlpVCfXCE/jMij1dEZdyzOGzKufyeaSp2AigkcRx4Q
5atBMAvy8aAK+lQepJ9S4vxINwaJwz/Ap4TiMJS+UhWKj9TKUSHduQgUptW+n/Pl
u4qByEHwZqY8DNcgFcR8GbLze9Q3nCf2/7Wh0R/nwR+RIRCS5xnwEmJRn5Q6cAYO
uZcBB8JYOgbobHShJ3KoLM5OfjfF1dtdTTXIdsqAkS4t4flOsHJVUS4OIIylWJaC
Ay9OXcgLNvx6Kkc8su6eB4UvdLf48k3t4InCoGWan8IPMzHBjoG7PEASRWKcHeX0
hvlvFrgA17Z+jrQTbQSbrapQAmErTGO7pqcqcyQUwMKZrArq+lWaRBHEbF9NTW5W
ash3gBX5SDjR1iQBt9HuvzO730mjJWlJ71QTTYhaUdu2qwjy7bZV5SJt7jK+Ad4D
d+DrbYMNO2kK0+XnvJz2cQsRY8etftqjNXO1B4TiIHrVbktfJ3IyPCCcWKNQOEDp
DwCFyOAjyn7Hkm2g5FDAbB68YaQQVUoE81mQzBKMypCEzyLVohNF0oA991sjUxYO
qnx/O4Z287nVkk0wqjYS7sS7BKLLZj7t8z2m1NbPQiWiObZG+yrPv/eHfPGfsce4
XSpEOb+a3upZeOW3r2bx5ZQMQkj3SHsALuO1V4F09KsR59TUz6oJXyNGLdUhrTqA
kcq4UKq62U9CJoyMjlVig27xR1EHr0HLBUyycuQfiTGQf3bMS2b1Y/+TgThZnpov
HKWFeyK4RDdTuPYv2Bd6NgvVSDBQPgZRr7r7ykiie2zXajHI3JKfSVbnGIE1CjfV
+p+L4MBbuMOeNyeFS5UplQ8FBslQCCVWwqS+xQt8pSvY+IJWuV8Ias4/Xk3D2PFS
EqBSzNpqk78CUAPaChwxReEWicV9h1MJZBYaPSCEImi9a/vraH7HaPpgri0/+MbW
+NwpvOv/PnpUurnjFMZ/C+DsrF8yO+VXaJuIr6cxx9PrLVdlhIwbf+r40J6hD49x
0Kb42heYSNic9iwkStLQjV6b0U2C51qnGmfZTpC/Omo27twmrUru131KUu5huPMZ
LgS1wtCMtOZg1OL3VFJ0RNSQXMrUaXBjuixj0IJY8AHLpgfw7JlUhEYbCMP8neCx
7vZ+px+ulSotlZQUVxx6BuGlEi1AjKxwV0b/XWiKgTsSpVhDNIhJGf+6cAvc3MJe
vBuD5g3xBMiaT54lfYySArtSwKePJ9XnBdYa8UhWXEZhJmVqduyYEuG28WBxkHOD
+gtrYZNGhrMbbkOCu26jbF65RAOCkVe9Blfq9oikCxNfGEoNPwWg1E7aeC5/u6n3
GlR1ixwpGo1l5486f27JjkI5ZbgWMTOpeBucafJdoR4c+TD5ClYx4si2P/J4Dm5X
WpenUbyYpHAlKdzIurJhUk74OwArk1Whw8j3GtQM7QJvWYJ2vN5rSrzyFIehzBPj
LfuazWmV/sb7qVErwgaOatCI7rKFqZ5cYiAqaXRXaWogyRD5BNzdoYOZCu1YThE9
Ou84XJFUIRX361Kn4z1o0ADoITrXFr3M+vmccx6EraJCVAXQhQmZ8NQxsnkRZmC4
vhVEV3b0/wO166auqU4pznwbOQxdacVZUIwmy3VYCL77Gmq+7TJB0NgtgIYDu6yg
lWXRVWR3J5CaLkliKSIlUwW1pNsxqXpLQxmSyeJ+xIIGufasa4q08nsmJcFzg2kU
ScszocuAgWGbEmMcpNNCumHXbBApYIfCZCDeBrS5p6u9O9Gl0Gn362Vd7aB/GQMz
tKh7WSIvW2zr9Ir1lGMtIx1KpxULvpgpXMuyYtVFZsysq248gUa7SBK8jZzfGGWX
YzP8wh0T9KGWJwxKOqRhtRbvUER65HKGQHkRVSiTaQV1qHGrBJLS2PvkNawv/+ea
GFionnxEaiU+y0lN+bPGQ/6rYFB4YaKlWYMkgV3WaErX49Vbcy29KfZZgW14jcGi
jdyLQWGJtVrmHw9eJ2kcJ36i1tubtJZVHQuMDSum+av+TtIZ4mwNkfRAf7+yMecM
rZjTCMx/1jfGYnPeHeWthtBbXBoV+pdlV2xaR/dOdfH2IucBA1axbaW1kSlGA3PS
6BbuVjOu97TKYnxqhLe7+kb93GRfedsh0nqrQm7OgIbSmNSrqZXrNxct/lIvQvUl
q4Khbifkq0JgVCKx/hcfIDi0xwnze/ToNc7CvuGfM9N3v6I5q4Vd6WzUH/NNeQE2
LEHX7bq/Odwiqu1i80R/tg==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Y58OTqXH+Mw8kTJYGOiJwUYicMS+F0MVyTQ7sKio0zO4KiMpP3NkBQnLg1weWJX1
nGMKJyG4r0kibklBVCtYCj/RBMqy3jf3T9IbgFJD+njW6haNKfxCAgGmUwptWwOL
PHp2hQ8SzUWbw32hz1MRw0YEaZexwmQRQ5fm+vHCczI8dHlBgf8iuI/jDZEQMcQF
73VBZZ7gqaTztw8T26Tc3bvLaYTe3r7ReHAUcX2LCyUbouTEFIgV4V6sdmkKpxjv
xtr6adonQWpXsqAYtlweMXgfFz5/dK8avEyR2OQeJ0TtOwzZiKnZzNVnnYOujffg
zZrFl8NRi1RC4lcHDX1SOw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4976 )
`pragma protect data_block
pQC0NX7OBzu0y+sqh+ycGX82Yqp6ls3RF5/K8XeWKHWXyYfspeX9FrEiky8/QJ07
KMk1utWjTITQsd/2SbXuNFWKlS+r7/xirRCPUH38BpvaTEpqeTGi6VkFuonmD+Tp
5RYsuJKaVkfJ+0bWgT18NzZjHVLNYGX1UrpIhhROiIfFaps6y9gI1jIs+cgMu2lN
MCtrKcEHDjVlFLMDDeN70h0Nxd/5u67RYbWs+KES7WsyvJxJ8YhjEexJBY7IVErE
StKIncHeuHQ7HVn0VJQtl9vUUpeqlcFPWaw1LFnrkilyldYpzhCMtSDz7tPQqvMe
UN1t94LVRCBYaAonKdrZVKSVH/etJ1Agu75ZPvTcGsMG2hnYjI2eWlB+otjXxVi1
75Nv1DW1U3PUo8PqcQ5AEiLD+M+yoNWnjv3MgWHdDyr/kDRvcWUtZLbgegf1owCO
GyNp2o/2JeSDYUG2lqzM6ckEuKSGYYBR+C8LL1EKZo+QDarPPLEDqOkk1NIJDxt7
8qv5d7jU3IAJXi8cMC2GC/MRCK3kj8gzJ/K1xswshoQTIPeR7OA7Bmetke7mWqoK
A9YgREJh6TYCn12z7NnU0fV5ZLtxw9eWVSo6Zlwt6NEJ3jjQ2CSuR4e4WJeXDbFi
pi+X0gOJWPi35IPAiW30PIW40dUpjWbV32cj8mQ5tENnfTrA5OBFQP3xXvCKtV/1
cUMdNGP2/KIPl7avCuTdQ3rivIP9UcyNgTpjj6uzVbIhDQPsUwjMaGBkmcBt8IkI
6dlQIWxSQF4ySaMwvt+kwIxNXnHw9R2NBmgacwGO+2LRSS4rFgxjBFpiIReejaYe
dRVhpR94eyCmJW/K2700gtA7dSaXOF7BMNUFadw9PYlvekh2GNZK6ZucJX13QDoQ
Vp9Z3002riGhWAKUK0oA/H9SJ4u7PsQhepGLtdChsymotWUCR2WGbOaYlbMdOrCh
qN827cjd2Tlb2QmE9Fu+f0w65GVa0n3TncFxGSiXWh5Slfx7ZrpNiDht+ot24Era
T04uRYRhqTQm9oJuzFT3b3gFBBuEJvWTlqwd8mOlOfq/vMq5oLfix4CGvGuRD+TE
I/tb3ehJJ/g44RnmNXWDsHie48xP3HD4mhWOIXc/+35J7v/nOTbDDIwtz7KNcAHJ
uNpduVjWTI5tzNgebEJcQBeKMMPIC2vi+euVgRNzLwaDwZcIEvJgRAuRC+NIlX7o
452mgOCHcxyNFjxiSlGoO7YL4EzMz0bNFSNKSN1G0Qccni0xh3UXtOQFukX3a8KI
bzyBdQIJLCK5zkUJqSQs7WruNY+IqqnAO6V5gKsGO+xo1gB2isg1JcgkeR0RjNft
vhTbJt2dznU/pSl0Tt5fAvpPb1CheQtrLtLw7YjoR9dgMFr6LG/EpAtxOh/Ql/ky
ZSiaB+ELEozHiB/oYQnkOO1EmWazBxyvgkrGx7qAaAlrRKpNr6VHo+XZHnAkX7cM
/FK/oBCrou0sRbffNzzlln3i5gyV++HKe5FJ9SddNy+SRMBea0Ml75XbZmTIqvy/
BMsOR6j1nw6vFPvlOElel3MVS9UnqhJtjXdsovY1796LYsgJXmVkiDlcF9YkrheD
kF+zJeN09+MBPkU1de9h2iiUmM4dgiSp++D+DXRqyNG7qCnNSWbsebrrAh7/5am5
C2RljFXTTB6ORyjU+5vPDZs1tIjcXtPICIPJnpaFJkfGiiKWw/BJLsujx9aGiZGq
Nbe2qCp05KR2b5Y7gAGZqM/YlCcgsWU6pD56Jo8rRSEg/ToPTqk1Crldoq8Tntei
yXLAu+xEOoKUVEYAUW374mxcPi/9Y16ex6MyNNLXspaQaVjCXQ0/rM2R5RAb/ufy
l2YacQqEe36wQY8KaXFQbRf//wpSN8Tl3lBEA0pQat+KmraQi7nDpSkeQVPnDwYr
PTLP9D7SGgNEGBDgtFT+bwK/D2rzJCWd6AmAPRWHdThxNXclhEyYgsZ7Cypuiqak
Yp5prXLMEs9L8ZOVKHMw1imRnpoutyYQ32AqLfk0j4epKsJBvL2kSDFcD78BsJ85
CVbgSRmpUrsR+2BwOJnWAy0HYfTni7P8NL36NfkUz10i9/bS1f9eqPn9TTXdlM/G
2ZSPEMTV9/w7rb6ZHlrW3XwhC1qgDiiP9C89vFkavBtINxaq6cJRV9obBRxbZ31a
Hm9Xumee6ldIKXCN2TVLrQb/yImcPriCv1QSUBtrzxxw4TjqPAfDdeBu8kxz2SYt
c56let9nwwrEcXVaxORHIKp+jvRRByZu4zimMqsTHg+dhParKMjpe39hdsy3CPXR
zKikHAqdAyWZBiDzznNnG87oVWDOi9+lAaO9Xapn9F4en5I2IvsJnpZdzpXygVhL
vPcyUQepec+6dsBcuKzuWtDRFnh5qpjbWebypk6+Ylc0SLiCj8yJdKCcZ6EB1/Ct
TAGqQtpov29zd72aLnnG4Z4DA4pUqZ464Oh95CFvkVMKhx43S7eUOCL0YAvkUgmc
ipdk73ZT5XDX0NZnFGwpwi0W0ZnFDYw1O/lg8DfdCUaXhl0t3ISyUO2HcWPL8bmb
r/KU/ITvKKwjhM5tiT2oaSfxTPjjVjsEyAhZWEOmX0oR5lU4xzw+mIqeQ4Uuf4dI
C2yekbr2LCjl/2+UmfPsxN0YATMqHyQWT0V1jRiAKIiePbgXYnnD9nA8XkVViRN0
A/8KtFo2+1BRFomT6QaxYc2BDJqgis64RAvyghEu712pX+zC9ND+bgWKvbV8tDCU
gELCCpDnyDZF07IZhmv4sjHhuJrDeMe5QAWk+oxOmXL3nBsCVIOt1rILfpEDyOQh
yvb+aEN305Fz28FV5ebMkgTJH1RLyFOesueoIpCdHrOoAozCnXZyu+C38AdAF2Mg
8j0hEOvm6D16SdbJgBEDUyaFgHquOBjaC9Y6vnQa8eMzE7lDSKIEb8KX1CbAamOB
Ghs9Wih+J64gTmeOJfZSvqHo5BZ1myWNRm+z/rf/Itqgv6XUv6A1uqHZU3cAVgBy
fkk80CjzaWQR6mVbRG9sk8Utwt8bK5hzoZbNzHfXH5L29E5oA8JrjpxtwsoicG7Y
qjh4vo3Vg8Tjd0msDrBa3FmoX0c9n+e9PHFxNN/5noIRXtK36fhB4aU1CJhm/vse
/U3j96TechwFQacKiA7imqJPplYYdKRt7y6EJqE1YnPprDe9Ek0WyX27fXAOH1yS
lsaL3RhTJRA+8nfE2CGYPHW3wRt4Dzn4FTFpOA0poBw3T/fzYdjIhik/ts8Lx3Pp
DX0V1KXicWx9/2As4APOEszXkR5PxUenxXWmgm+pmD7I3LNmisVg6DbdFPlODeSj
X7nU3q+sE+o72zyPAjGobAD19kOkZTEBmMzmoHh9wzAMGTYULbdJ/FuJhXwGsomJ
SgeBTSVXRltJcQeDBMIVJpzxoBAa6AeBSzk5QRWT49f9J0W7C369/dWiTHj3D3zq
pMeIfVkt8FKVrVtGa+Q9MsU1PAMcfxePClCcnjAnfAeA5kWc40Qstzv3onwQ6FXI
oseUoKdwxQMtPs2r7oRxQInxrL7VPEmW23k/8VsZa3aEsCsoBlkevru7BJghEtPP
j861W5/5FY71vHknzt1Tnz1pwVvxWMm63plGLr1fs5/6gVcmVNy0Q/3GCQbi//aq
xf2YgHGkyN1wfLlLw+31qjpOQ7JKVSghiqXm2MaE474A0GH8RGRi0sS87uXIahXC
hd7WWy2xuk66f26Q606iFJiIwx+Au73miGeLEnMZU1yeTTSfJFCcFGkom4sovny2
mnGr/yKS28oc9eOZIjxcOFZesFc8gJ7EfYV0uSgrK7TKX2Q/UgF7urwFEgoXjjjx
8VvKGxgM6z/jEKBT71CG0qGudxDXPpzjqJAh+50dvYadsODNwR7cO+joH64H6TAR
MP4q0i9TGKrmPesSRmXqvBN+xscUJFQDc10I7rxm5CyXABMiwg6qwfghkRO5bEYl
K9PRyLQiZ0HDVYTXNSedJcFQmRyOK+L/FBjRPbDeNvfyAlYsV7PGKz1VIDedBdh3
uo5arkglAGVsbSwMz8hI+J/JEnkWrrFT0VaUbSreEOHnOUW83fPzcH07R+g+Lf2+
A7gntjk3bYEDORuA62xqGYQykX9zjbrHn/RhSkzoXcL9IwzkwNCPEiUQa//PkcZ9
B67vfaf4wlnz6d+RU3dvxxitXBNrLlDYe5VwcYNAey9cR5YJCj+ts3/tbFVg5ciW
ABuQvaIiViTStB06CgC4calq3Xxz5k6T8/4p6nE/k+t73xPLonp83IZzgTh/R+EQ
Ds+65ppTyMs9rGCIAEsdEPAYDQsBgcYOGUdL8eXp1QqRqW2w9+zlDT8RBQJnCm4/
hn87iymhM+Dtnkby+q3+AnOdzxZq5XMahvHejUnohRCMNY6elD05BUGCuIHjRu96
6634UHtLbmTP7z07W/2rne/vw2YRCl/9+cNZechmZivTQDiWLxh4VR9+qRoSs0vz
aUwgAajTCqkbJ4QxOY6Ue6Nyc7oU/WCZDRZrLw5hlofcN7KqlMB8jHAL8aSQseUK
O51RC4bh4fYfBIymNG39pUP/tSf9E2vV6CRV/1fWHT/glCXKKZ29Wv9UaLgAKIdz
s00veUJ9BX6e+J2fwv76QB7d1JXATQm3c51WKbSHXomLiTLz5Uo8J2EUzmiaJVyF
1Kmpb6vXTGS1KMvQR3OF/9Upn/6siJaa+zg4bpa9BsPOL3+6uYX5F0/IFtr7xP4t
yNNgn+KqLiP/8FY7xzEvojcJGQJQBeG1Zw0S5KhYwVnFEmSN01eCQUPh8KBiUu3g
I3iIJhwlMqFvCn9PSMwxAT09O22GsaGrRfkNC9yuH1GW/KAkRyolS8Ez1evXchgs
6c8EPZ2pU66VHCMqbrmpUSXbflpJYMDfwBQzOY5VHal53PwG4XycaOHDElLiJ3lk
oFVsSL+F7YYZvArNY/mj5pV8lPPGX/dCWUNu0gy/NS2nHsvDQS0W0i99hGoAnU1v
I5wjmb0r38EqxBtlZpwHBsw6WaRIKeUuIiRhFBPFNXmXRFsS4PEsVl9QtTPGb/QY
DUv+rvR6SH6YupSHIYHIzE7tlBi6fGKpDnPAHHEPKhRRlFimB+KhtJx0+8c2ySiu
1LgDHPD6QyYfiTOhXhIdhXBp4XEKX03siG/P0fLIVH6wTjxZAL0BRgG+srlADucP
xB4s0fJYw8s7811EnKVAdy/beeJViKIUURzYtnMWWukcEpo+3guZtXAR+tKMnWNj
ni0xpOuY5jBwV/qUysI2eFSfqx95IQsdNVZKb14Who5CXCwfrUa54sGAfxGUOATr
j8uIhp7O0SauFxOiSP5f4v4xc6Mq4b0tMnb3Klu4vHz23fMK9JatxFKS8unZAgiE
Z1WqV67tYB9A9iCKbTnG/pJCrCfBWZKwFGEMK2xcT5y/LrTZ8NqcMKQPH3tzBC1N
RE1RozYr3keLCTmX4YWbVwSUTxK220C3HOGLqjwbDVfBoV8Q71VXV0JwNAgDqi6R
HVgOCifEyMTzviayavyu1Tb5+MU0RS+YpNSduYmCBUU7XqyzlV8eB0IuoLff2gss
oWci2dDmXgmyvR7w/rB4QSsqAcUMt3CJOLcg5+6D0cX8VS++z59mV1s+Y798QtOp
b3LjBo2/+lE2ZL4qsLZ5gMoPM8GyjA49L5F74A1W7nCWnoKuIMKH5HVjh/TmAtvV
ji6xG9Su0oBVliD+Foy5YBuVq2Etlk9bIKvD+aogoPck0q7bwgCyWEloCBOSC+CI
DaPgBXMj7j9KjKrpOXNFNaYufv6xItE6fRKYjdKqMxDN9THMeQKewTnK2miJNUwf
gBLM6MShWIY8H6JK8iTJR3+GuI6qoMmcE0mujvce3DWczTVSKI38ycMFv4LALUvQ
HQq20kKjoH5VFA8PjIWS7Xo64pZrnDPqOcVGBeQriGnOq31t3Os0GZM7nOU2MU4l
A/G27OsCOpsW6/h76v5R3yQ8NaZlWmc4nOkTJVkWgEdW/cZfZuOr23ocKTUQOu3B
qmLNJCaoa7e9T8WJr0cloDme+Nj7TYbeFtIcmTaJlYf9MC1yhJ7d1HOOOGj1MFHP
yu3aeB9lufsHI1m+HuyTx6fpcrn2SbJeY7sqIXnxtr4kx5qhriH12gnQDvhsR9N1
1AWPoeuXqMEWzw4RRI1ET6wy52o7xF1GWJUhNJVqzG7PBbdjSKCb7Y7VrnVYS6Lm
u9PB7iUxXSIWZoldxQINK5KS7JdWc/v5OoUyZmY7g0fXx02Fckq9q+yJQa88aOSz
ypJPBQVolwIhFpaAusy4GNLcS22OO9V6BcCe0kY/IJ45EHyecUh923BeahlCuAtN
N0AylZQCsQ21LdFfucVTO+hh2FQUjfiXcyYoOOfg/eaIOZcg15oMtUNajp8L4Uap
XTFmnqNqCRJYXgEmOxIrZ8LhKUbIYWQTdfYWr/qWmG0ETZpBoW/6Ce9ngSm6TtmE
q7wol4CSI68oUHLPNDrVwfhDfH7aJTiNFEGFP02qQ5B31/ss+tr9EODbcf/VyB26
VKqA2irKXfQT9P/zdjaILC2Xdlp1dHvT78UfoPaJKxNz+fJSCR0lgZTg3NnY5JGd
hrH6Nf8NcVWA9T4BlhKlrpXVnBwLK19WL20EZViDW/8=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Gif4UeRQHQ0ZKPxjFtn6KtwYvkEtO0AJ2WgR4yg5kfhDH3YGuj9tSs7o1Ox0vscw
M0G0qUZ4CGad+iDwjb2FeGLWVddrdjlA1sRZs1oeazKMeqLz7yp8avLeioA85ygV
md9PQvbQU44/Ns9vsFoTlUvAdA9c9L3CAVjP0aNlEIo8vs+En6YOWhms1kZCyEPo
fJV9mkTtyc4RnFnMLoxC35K86OboKus0hJtQ6VOzMMSmdIq5/KeD3Hgv16lc6TJj
Z4IFws2aS91Jmj/lUf+/JPRtE0C/3x1lEw2NZlJWzcp/5Gmfd3/Gp8OJlYB0MDEK
ioOb3ULG7am9RejYjcN1cw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5344 )
`pragma protect data_block
hgMoYjuBU9K1y5ewioRfkzgT8mO8M/riRSPBeVbroP93oxF1w0MAKU17b7b50gW/
T7aUK8hJUbPGUIXwMR8FeLsap/F8avEWzWaxtnKidgdSa1djtDNlU7FzRykLN/45
JW3ABfEk7+XuuPY8jAAECJs8N7YVi1hYhxPQJnMzHHtfOeqGKRpxJlTMoCDJE38K
eeIFtrHE0EhwivxSEZ9vR/fFy/e2XCkQ03sx95PfRb+gqzVrHGPKdKwq2B/DCYow
AwLfPccVIkvDydcYmeUo5CWYciwrGL909z2vO1WWIG2/jUEw6GL8d+uMTR7E/A1K
bToWI3UggILhiuQ42n6JOXyaGUDNzYlXUGFw1FaCSM6tdNhJzQgwpq4M6bV6D0Un
x9pVTKYFDU539I1JiywP0bQGojnN8YoRSp5RdBqWAcSMK+iOrGBlFOKey091xNa2
+1B7STvxzIDWOJfRGquFtdLQDkPBnT7lUrwR+RgLeUsvL8Mf81iJHKKFdpkEKTkt
Ea18GCq62f4DtkTQ6m/5/5+j2W/ZH4tS1PI/HJBeO5ljK9LrG1HpjAegxxj+dVRA
tABJsKFwP3yZ/4vrZDhDH/1C/3JC24hRQRE0TwMhVdzC8rO9XDH+4aHTM4eukiJd
ly0uN6xpTBDlQVtloW8KbME1OpKor2JVkDuJRCSvYpfBpSahvBWgvlAkm7omJZhh
cx/O8+7PN4badwXTahOYEkBpQjL6yKecmf8gfwdfa9UbL0hcbJU0Oil9vdSS8WDH
Rfl+DPUIJRJvxOpSxXB/cbZLn7jDIo62tnYOVl5AEyRb+WlBsZd4uAvMDY2lglhb
eeoDbAuDsUXlmEmPCJsP5IXiZeenkpgPuS7T53VcLJKge9yukwfVgzbfSIdl4FoI
ZrDwCjQw00AhQjrVFoVcgL+ca8kfOoIn7XO+40CHW6cZP3naXlmADHm2krs/DsQE
Hy3iEHRjSCl2I9yXro2XtX7NXKClr4Kk+N9IathGWsH67zxaxxB/slLg4zA5wEjf
g0z6qZqufGkeQHxfkMbm0XY36tVqRipZjqat2VPS2yJtxcl6pn10IefFiXm1pEnf
S9ozbD664CdS5pw7Ez8H1ZF84Qdpk81+mHcifndZaXN+K8MsNUCySKDc976KcVlf
KlZxvac4xwOMcbCQyTNSdVol78Szx1pWtTZLQxOtniP9c2uuMzdbe5fPmUGKRobu
fJa9zJZxm1Fk26LBmqiVyATfzMSCVQs9txaeOvQpxyF84A/RXbpG7pEBARegVfLc
8U5wKmyH5bgqMlmk9TOARGsU16V+vzFd+GWJQj3MAOfqaCS73GAQuvShAso+vLoD
L/uRBHqjHL81r8ZETJbN+inPOm3OGT8Pzz6bb3DYPvvOghzKKahrvxix7V8byKFz
4FIlRNTLkzwumnwhnhgtB7jPc1IbGC6QAgmNHJyes7iB4aYgr8lhLj32/6OuNz0N
hWiYLzp3ddFfBgjJYHa92aEGA4TnXrB/bhYop/BKevnAmd0fGVeRnYRyfp4OQyMJ
ayKbi6hbgvfldHl3nI/sQcY0Esu3vQK2HX3xp6pmaZGKTD56+igYgib7U13JD17z
tu8J0fSnzzKA0oiSF8zXBVXk3bOVVmwgOEpZYiefBxArN5soUlYZoQM0gEQfBBr5
gV+514J37X60D7uF3Eyi1DU7tFCP0klfZ2+1TpxHG/U/VWr9Y4D34jHlyDSDyilv
11DDxctksp1dZwC9Fb9QpM7z9wxHVRmNq+5EjT4CC+ByO3bxxhQ+XIKXhq3QMS7X
VANmV3EBot8hK0SsYxTf3vgyauc0Bjpjx84oWXVoZkmmm0geOQvcurknZ9SSfjv2
iE4EA1/fQpHJHAkhcAO/nLC4U1mVNPM7olI6+eLwHE7j9YMqAO65YiTYuC5t7sRd
zVGRER0112steQOAiwsqzE4FV9uQP+XwfRL/fP3KhwBWgI5O99eQuFX/U6H9ka58
QKG0pQUX1IfRuKxO1TkuyykDzhddNmTXhqcQG38PXRs4yANpHUVF+ZP5XuVAp5ox
ZOwtjf7QzEZlDp33zcD3d4gKo721Pmnq4aLs8iMATcBwWdzV5HQ7m4MXlfdmfO2R
vZuh/1FoFslQ4BGimXnMQhZsYNvyizQbkyyhI2UK46+NGpDgJbQyhg9ZSBwUMFBl
ew3lQpGbfiawMYuFE+IV96aRJl/IXZsbkEmnX2kpRne/Oxg2NM7EdZgkqsqhyxUW
8VS6ZNXTseOZKqY44OHSKJ1ZP9IKvA0SWg6XfZ5lAnM6vaYgvcdRfu7+wufCBnzE
iJt2XCmNH1PV3MyINbRHDe/Cp1kqbgQr7BDisvEeRal3HByyKN2Xgc/GPT3P+zwK
XCF0kORdMuzeVdxRD2E2rsYtTv0d/4ANZ/N09P6+N543sHYH7oe1uxKYBzlp+Dv5
oWRtF3YN4l8vqlTQYPisXoRYjLYnzy0k0T6fNNHHT+uP+aWCn+fthenA3mcfTjp/
ISms96SYc2ykjP57GOCo410H6vtsQ7z7fDFRG+C4GZGcZ6YpZkIhj7+0GyT+L9yk
aUmmV/EFH7i/7qjrrn2AiWVQ7Nq3Q51tfjr2alI3untc9eqJhKbZqKitABV+KzEx
SQIy4t8fQChadQIVaTlcSExOcfSJY/SSgemMiCf5HEetH4ZIHniBXfsbAzVVTLL3
ZAy7Jc04OBTO9UNc3H1QoN6/i0I6Q1S2tIET0RZLDb4bIWb/32bMo8UqAN+vljSU
mygswypPJ+D/R/iG1HwFXMnQCVFp5NWlj8wocQ3fPeB3M4NgfauOXUeYfWv2EQz9
hw271OOtIH8Je5OQbnUp9kJxieROO8wARdnxdFRYw5ENcRrPkKDMaKAQLJ4V/CQt
ExAd/qAd3wdADsZ93sZuSnRXYXnTg2S8FBR+cB+s5YzoIC39UIz9fJHNvxc1B1BW
kQudUppFHd3S63yxbHB1DcnUhACmB9YzOeOpb5BOy4oc2iJk31LhpFIn5vkF9yrr
yvH0J8zMBlDGF2O7qTCFqfvWo50o6hIBehHApFMUG9XG21Me/2Nz2iZSqvzhYNxK
2ypIkBs9oaGvDwCaz9cXyKwkJyO1YEZujaFCqyZyn++4yL7UfNd9BlZz0VN18HAZ
Hpl33q5lY+0aQ0E4rZu5KaN6eZ+ijRfAtlFxwm1dnD+gFu7ZCeodrlvW4wVkTllp
+/WMqI4dlg7ZhxvEAAlle3VPoDOPeDeLUVqXGuvpEzPm9WT2mVOxdWMH3g8TOnhL
f+fNfpZwjis+4QTSA0HmkstFlFu7L3XxjMMzgFhU9/t6GLShVdPC/C9sgy2QdOm2
VYoPSSwfF1GAqmAeQFlCCDeaaBIMZdldVQCrjDmfZRL6adCpbfNHwjzqqzazNkWl
a+zvyUG5XBysdbqCiuZTfDuvq0g6oC/02rSWLV6vXj2XqFy42hihYJSIALuQcwoO
80/7n7rjTjBhjX+iGdX0O1VbmlQvP1VXtkTx1baXTjAQUDGsn3cfEasCkHTJPpdv
yVUxAN/+IgTH4XLADU8Bri5Nt0REpG0AZPeBOj3Vva4boJj3o0V1cCODgIySv5r4
M6rDFlxF0vmlWNIakIqZ4bKOT+9RGg3BFiDZvmfAp1674yqeKBXIc1QK87uEYPM1
LJcnh06ZI9rs8he0YC/wiEvy8wYhmPpk9yxOTg4T7HlWSc5xtJ8Xmhp9OCRI520W
PWOV1fS/1gSsDOTBvWa8+7yOtIqg4B+ilFy3QIC4T5ZZek50lHmOp0fR5AMBoJu5
EeRjqnzZNMUUpEPC6NhyfwVgJMG5vId7iDM/V/paxxHL3sYon1XKPUuEky3OECgV
83XWoQ+OClETIIuhLLr89h4GnUpu07UeGjkHQ8F6lryiAsTIHwODhAaQ3yZEdOEJ
2cEv8hdoK8JFvfEIzdquBlrGgJGjtnKBnMbUjl+q/N6K2U6BMR40mFO3+fxb4X63
8bml12eXETQMiAvun+qf9O2d11iYTR05gSxeualKQm+Dte2Nly5yOIZGkSzHyv8i
bMCCGhwrRdMY1tubbzxSQ2Fo439h0QSA0o4NLGIYthIuWwxY4dHyqGjAfl2v05um
uTm0+kgbi8AA18VOY0FgzDSlSM17WjgE2X86cjsYSU1Tyu4/VMYw5hc6yUJ++GIN
cUJ9XNCx6A0Aip/0ki1GUqHyV2ftKTf8iAz5LQTH45ongb+14jhUcTx8yf9S9k8C
ftblEaaetAflESTqrja5wfK1e6yfUjRmtsmvhepG5yUCG2xvG+/QnKZuEBWNxcvi
odClpQBCPQV1oti7YdfaRtySEPR5sHlXxpoJta9Fv16kfMfTcVsePRPe+tYXHvCC
2hL3IWuWK9Dl6BMfVYAow9zEXckF5N9eDo1MXywl/a/cFv4lSNv6vs52nOsilJ8I
hwFDoyUm/BxjwQ+0C10OzWP5z29v8qjvG9nxdbRorhVhzxQtN7gZJ/tOyRGpj2er
PUP5RGApTr6Yz/LUIlHO6glFSe5Ggh4r0rdF7TwytXFVB4oKH2GOfzLXEnrrklU7
ygzcB7D4MXv3vdt2MO0jRZ+rsmGnExIn1so6j0gYwzQCqSmTCS8wHg5RmzE/DMbC
luY6s19HxuwC6hnD6DfCaKMgcwugKlxcMvl4FPSoUL6HKAbOwDO/zXQ1cDTsp/FZ
795+u2utyJdc+hX6X5H6N0Lcd2qSBGXJ7zoTNvrC5Zl+kHdxBQu56X3MAvzmQ8dr
JtCG/+kBSz0EJxhN/NeP5VA0fvB0ep4fLXOQh85EEm95dlhEVpX0hAlXvyLOj6Iu
NEyYxGDjSBFNcCTPvGFUyARvEpsWtMvbJlr/ySGJcugaTjXUGE+ngrdXV4iNAcwr
8RTO02WJpkNuXeZ2du8vQjV3G7g3+o/QoytVd+DsdPCysBHo6ROtsAxZvciVqgrA
lW98hEy18XRJJtz5BWej8GELr5x4v74KD0XfAOTDA1F0ysdDKKu4NrnFp5bHT/tp
sasLfx9YGRfpVye1qPuilQiptXYEmnJ89BOZ/0Aj5Lh/PqHe/HuMMsQnJ6jW1TQQ
Wi47bluyPKf0/POi9d61Fs+0vJt/W/B4JiS3FB/bp8Xx9FrHSYaSRMBlI69J/Y6S
DkMz5NK4a/tWpRmeOORKzGx4Oh3aTHtPHia3JzE4TwMpvVF2IQHzcUnFeDzeSZVc
zhHJG/ZK/pVptwLCYasLI/UhSS4bp2cCcaQNBP6lCOOWSYCK+sK6vOnU5eYh6Z/I
1SBK8j3euEW5iNNB3WQ+ChSmEO6rcdOluCQxlZTQJ+IXph3a/XtjPDlJL+b/jWxo
1He9chNdBmYoyTQDdpBXZcxYBw/apQD+AEEXjbhgNmOLcbw0eJqWs86Ef9HoVemP
SeE+qEPiye3TUIFL7PC6mQCQUWdlWAPHN9ljq6kpSXmZ9Kjq00yyQFqCs415hs8k
CV2dCys23wBanZozTrhS9SazQI6GZmT9KJRIlZo0HBd1ss72bveNDjY6M/GqEnjE
bBzExHcMRJ2X7/0NJMs08HCYsOnY4xfE22/dPbjhi8SNkfNZPRFSxjklodT0DmwO
ySz2oMfmJa9uCbjxEFGrE3E4hXpRt0dMYva5d8CzoUNebnHV32BOSgqk7L1Ml/cp
8HMiw2OUYwdFAKy5/ZPw98NxW4/mpXedTDIXrDkI5aC1eaPtbjQil2rn++DeVEsn
GL7KVxjY7zWScmeemfM1VvVLwmNQqDgSCpvziujsXE0WSBaXQuA0+ZLTL1c2upNe
wvVExCOiKAbuuOb/htNfp2w4BWpI3VSzww+MoEcM8pdJPeqBlak9JvGP8zIsDURX
VpCG+Un/AXCSyuvZq3q1sRG6AcUmm7AwcOMvtNmsFiU2p13o1CHftnS/NDLNFyc/
hwfA7J5WJQjsdlohRg9V3fm31/vQAJ2B9gvy1A1AoxHvVsUfBoM8HGtRf2W8LGbG
tANTYFKYgTh+/954jUE8HT47CSXiWk7KSNHCY/3zoBMS9RwyHppr+CBy3CHWWmTS
HyQgpVwk8SV2YRS3B6PCfB7q/opXEzFSJMe2kt/yYxgaZcTmX+hOj6Zj7VhdMlfL
Tn/9AjaBguieGavCKI/cLZx1omE4ssKd0n5dBbqAr6Ne5IOAadMx5eLbsr+fthrD
xlfh4wvF4iZbTPNWyVA1H4fXUIB2eLSWzWuQM6KGbWIxHDPy98g/lJqAkXFejDZQ
QlRqg3MNfEzqEZcV73CXJvAc0Whq+v87mUEBV5MKVEXtqxhpRwsWqccfEOy+V+Rs
kGpSx2/eEDDHAwZL7iBe4+DrmRVkSTD5mjWUDnmpvvGfcGZH0baQl0EkcpBMlV3u
IyMGN683c+0rXc3ts2iSMtUVF2shy8ul4T+EUC/mAlcZT9MzhMSUCbS3kRkEgMBq
0O5bTOZJ1W/gf3KXE8G9HdXe/mQgmi5jBhwEWe1/GE7d36j6ujRhftDnwwqjUS6l
DCQhCJgZcQbWsD169ZpeM+1i2U8FvSkiNWxKCmwas3H0mNi1AGKkhvauG7XVoW86
4KopprBDpSbf6JW3InCOrcPGsNsiW98zyXOvh6Yg04hRJwskASGw27UoyfCj+NcM
mIK5dxBM5RyQa3KLTZClGw82w0tL+M38eEbKw+pSisb9p8C7OmMr+9EaUo3OTeSv
SyFla7n0bLfvSIoeMowCgIN4w8Qn0EacgcSvrhYmTYxKMWA7nAXn4JOQ/igH7gXl
psdepav3jlAuWXePWEAWn2xAKZOTwI/ttTavH1/RrGu9O5n22qpuyEr8CCyyDCDv
ANDSJvw+x5YL8mUyKYvyKH8Ym6E9KmAZ7Mgw0iT/khb7u0Q46n7SXr6GfiW03Sua
kuO+WbM69Y/zwxM0N+B6WCuONuumIrOARHnqlUZQ37qm+7JEA2bupZBbgsvyYQmX
5vxYXYcJ7gtfmwzUih94W4G+CQ8emdAB+l8LKEKYVxOPSRecWpfcH83bXrHmKCn0
F+D/Oq9BD1mMJ97sZzMqHr+0o9tJ6/AQvXq/YbNSKT16NpQRIpyWndgS8NugYx6p
EJPFcShfDifCzQPcsESG7P6EMXvCsRlCku2gyqMoaKauqHx6xg/x/zEefsMkDrM5
R4EhPAMG7mKyzbyhf5+K4Q==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Nr5xxX8Pw6cbzguQfV5ndlW1nqlIRSCGuGfpkE9N9Z/Uoz+oR5BuxJfSHxPZIRdQ
nJW9fJMhK5ISQigHN2Zn+4BszaE0TlJ+x5QrskEXu0rh3CqMG1tUDd5qJvaeWl3r
+DXnDuq9wxf57JfUFn93mPWbegTPhL6Aznzzlk4Ez3GF9lX4vwUlz0JSHtoXDgcf
bWj6DEni8ZF9RIqmXgjLtrQALGpEr8Z1/yDsDNTZTN/W86vYZagSQtXxDCCJUmiQ
ojwl8256YQ9f6y77GL4HV5BXSg6pqUqwDJrpGbYZn+kjX0IFNyCdCpkwVxH8n267
MOYv5gm7+asDwFZCZ9c5mw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 13088 )
`pragma protect data_block
gCpheGXZYWmlYqg8Okj/6nyFbx49RomZdXBflw4+BPOiu53eWjRSn6HwndSY0VSA
YUmqzr0gMUlOLNwo+fQdR/FV0DQvFBu56DfZV0kfypIC5DllhJ9u/m2d8Byue117
sv2W40Xz7coguKaEZztuzarDZqToGu836oas57TBrFfpXvSd5l+Wn2wdI98QP+Iz
ygmW93qSRQefMoHoKC9M/EAc4XWK89cbVq4lr0l+jMnzD3NdbuRlBLl4jaaCovAm
/3X+GIPCd/TmZVmvGI+7+rLB4If6xshUBU986iXsaITgnQR4hq6s7UekFWKt8QyC
dc1DzTTWCyZiJaK7+0GZdpujVqs8LRBbgHUADYlb4JfVeoEMedan1U0s+MDdtmM/
t5gTKRl5zbLrvcl1lJehtI+Ui+AbM57fvmugLN87CZVkzNPlHqEhP3gZu3KYThse
wvkfr1TNgMikp0z6TbsXTlyxpHReUPcdTr4LaXXgqCxYQUV/NejqQmK1QuT9P6Ny
qYgOWZu3HooCrUafdP8I+Xx/W9VorQ9yJ1MCF/s/n4ZXo7OAJ3HynTFD8IIIT+g8
+2eSRuYy7rC61gL+yCFaI0a3xLLNhpjdDvQMMyLlGpPXL7d/Vns+NY3zinJSYddl
cYjLn7Zq09nQFOO+BbvG7WqRMW5WE8Ck1QHfFPao2ikXa7FpzxXcgHpkbEwm/z+h
BTnE/41ERFBOxzpvoYLwAOx4liwiqNNuKmV6EUW4TF3wrYepEvnuyr1LDeuRGduM
jsiF+TATBOIoAGNrxR2Jua2mkpV07MA+bw/mi155Iy8M7ih0rHjgkpC1rod4DrAU
Kf+p08oD25GhY0IUGvKBoD6e3dFR2Pc5m5jxWZ6UmUIOTltT/LHpliQZ2WT44PCF
2pMKkJvWiyb8y5LWFZsozmOKoLF+EJHEOH/Yxo5IJQ+2wFWGHascqkej/E7Drojz
c/4h9we+t0fdYctV7+hS0tmMjeew11x/9dv5Hvcci/4t9qHwHsUefL6ZawIjosaJ
IsoQRjED3CIbbOOfJj/9vnPpuqqKylf/LZxH1GQC9y3TujQKJxonHvW88FyqHrKH
yOHzFkfEUZjwC2eLXJc12zDIsFfK6/94BKIdE8oXhraNb55jjPEw74hfpE1UUPol
5GS5UIrrvGxVThC5/HNNRs+run7nEN7+anOq9mnxmfZCeDuByi8VWIx/djhBvM9y
1kcsvgKNQ4aj0Jt1tUkZgsDvaQDQj4HTPfkg2poO8uOzV3Fgp1/gM2SjbomkDUGC
tKLbziG6PwKizZ9UttkHPTevXOqkjK8aG56zWSMTjpTzgktYiA5CCfvNf2kK9qMP
Wr4URIm8zoKZ/NAJVNvr58/zs2X6XuP0kadU27XXpXChxCvWJA9bFbqqiLFkESw1
giARkPtkmEEJydrKExjkNOydVBHP1gIsaPFWScvR92c9Yss4MyaVy7YiTHbFb0wl
auAoIdo3e0BRL8agP/4D2xZPDyZQbwA+bzo8rJSOwQC89B0m8iOQThrsCCWzywgM
fYJV81CbdQPIGOFChnZ5tC0inkjUcZD9aX4CtQqoR8v3wHiGMRD7z+i95lzkVCfz
xHwL1D15LrDP+jcJIx8v6/Q/jPwgtknwwC1FYnOXZ6qNWdinkZvGVc99WpEFBmvC
AT+Wq34ps2hmYkXAoJ5K34ucyYq09Zb8dTL7l5HCvcmcY8oznO8WaPcFRwj+tiyK
ql2qC5qBoerpm41JY5oOND5utH8zQpRE+ENqTFwYm5UmPNS/0OH19uj4/GQU/jMv
00DP8r6cl/GO5xdtrTYw8Y5rrVpEuSIIxNHWt6Az9wPDDn9rUNe5MckVeRPFyEAq
Q+GQDQKyDpbgOshVn/xhCaO1BSfj04qWF+yA6eEfCClj/Y59RqsK/Aw5cBreyRJE
MKvANMlIKaxfYQQu49pICH6QUnEpu2MGBe+/6pJOAnSa8eYWj6WJZES2ruz8anQ9
eCOyXtOPeCEKlgf0kIehsZRLI+K4Cy4B2zDihQED14ShbKC+aCeIgOhh3WlIqQmc
bFHBIRhigQ3CA6PsjL406Y7NjDjdn0jRjHml0W/CPJoiob+FTJ4TUxOV8lY0u5r1
33QhdgYqXl+dAo61N6g935YKkYRYOfbjRRiwg98rV+UARuplueessbqOtk9/0P4v
eXW3UwNZXlf2a9njLW9AxLGy3E5uYYLPgRWH4CTPV8Hihh2Xxn3yBmfflwmTp22V
O1aWJ35L4AXhvlw2arD6G1x/ICsHLv85C0i8A2gKQUI1GR/g6nqjMRy1JvbiiD8N
GJWBGwwuBnKvGMefCy63qsSTNzzjXkYa3p8iuA9+0GTfxrutQNJ6HJ8fYJduAP1c
Wdvy2Yykz8NwzPvvroohu27+9vIE1SF+yBMWk2Njujc9DUBX4ee885yolg4+iDzN
lpPu2km+CR2DgiB6X9vPSpoeTmQVTFcvsGz75qp387hrqC2tRV42cUZUqJUdHZ4P
6ym2U2dv8jasuwyJuAvg61/JiClmDoF1sQXtgKP5+a0Vhl2XDbbNSqQlqrFHcBcf
QJRPdku6BFoF4/PIZ42eOgRbmTLdoOcCWfbMkI7W6QpAIEEWR9F2K1KifCAEmN/M
oaLmc0Xonwu1UUV0BAOR/hck5NFYPBkgxePrUuAeeso5roFu6n3WOoE4/lzuGRvK
aCCbfklnM7+NRm3ttgiN6w78CZEwY286Nd0kNaKXiyC5JIgKiZHPs+bv2NXc7quO
sVvjGbmkujHhieh2fIwu3ZRIdT2F3VXgtvEYRYsLKFNkCoceEVB0IhzbadONEM+S
vGH21h8WVor8v/592NqkRqv7FLr0qHztnV941Qvq8wW3fpx6LvCXeWo3nHYEiEST
j/lcHKnRZ4/iwg1NEL19dn7yWdXzq5oMKR/FkPd+A1LYsjoHjopDmSXLYDuH9stw
y3rYIpH70DAyrDiVmvOyf8/BDOT7Q7brGsigNTFjeafC1MDYi6rLHhTj3Qv2rdmR
oKyibs5uuP9Fj5O2CChAb9FPVptUY0aFMEm+tU70q6e+Kl5AVJsMKcuSP84D2/Mi
ufySyTuKf1IL6b7+VD90ybS3qoJ6LEanQ2cBqjvXB3A24pkRLjcYfOv5DZ6trBgC
pSrUgrluF2kZg56aqrXU9rlxlgUTuIBfkI38aI+RnXUBzWowXCJ6s3/U4cWJPVtT
S3G/+lJintUEmzT/OFVuW4JSvYUGseqtS+R5DlLC8tUwTGalwVlDsXdnoYtwX/TE
fa90in4T24KXA2b3KETvwc01Di28NyjS8gVV91Xr52fTtKGx/JOxigH0/c1T0hI0
DrRhIEMxk41yXZGlqyXsc3hznUXXU52ZetBOqpGoxIta74uHzJLC9kNufvMt/6o6
kCzXBxEmi0Kf/eHRm3pMLINpUuR0RIxXzS9J35wt/I0T4UtqM+sj2UdPw6X7jHLl
yqlCgTPNh733TPnsREDjQzMLZ/YWKHku6BhYD+W9UmAvW33dKJzEzcfm9xmedLXh
+aAasR2v6Je5geCEDFUZ5l5OTVhxhoJ3+fxSe/r2cKt+/9vHNAEPU7ETsquEHz01
tUMxa6UsGGM0hpfFOKvIZ4DhssZsnAu1WVgTTbjvLvp8WESv/fU5OVKIG/iMPctF
VMoIgjpDe3yDM+o4pHba6vocMlJSyLl9krKcEBIyepl1ojko4WGexkovwO8AuRQX
Lylle6GsYtM17BokzbX5VmApKG1bfTRlj3a/aCfRZfRUVPx07HmTysdxKXSGwaav
pl8twIXWM5ZItKGtrBOu7sZh8deqzmbcmomqcHDHdFkHQejgUs3MNvC3K84hXNT5
1YXP/bsguq7fiHBYbhworyv3bmVg1jak19037kQ/nLqwMM6KoIrQ2IU15SLdqEJq
SE+kC6L8WMlZ1w9271lDINYe40H0kgaLZqoZN8pb3gOuDCNV9TXCAw7vm4znf8ar
xMerGuK5Qcb5+LDU5Gl7j6GajIubkexqnKxv+wY2VMCVQCeEc8aWkgd3799AlN6s
uiu1iliyGM1BqBQDCD799a1P9rSKkc/HJX+E5DYT4nCpDYNIl9x2tjg+/96/nhyg
FtbPwq+hmbRU0BpuNg5+i0yL9IrX8cSVMiPtGH6oPN51ZPsJZnxB+3tJKX0YNn0/
KqncTfrP/BpCs3EGq0SNxm/CDySXt3WvYLUYxtNr/J0PnjrxEHhROsbp2OZ3ey8y
5IrYTrSbyL1nhj/OCmG/q2Cp8JeyL9eqq5o/1mxJVjqQ7yjDdvIBaJ9ySbLWibfD
5qufb0rXW/R/fplj0ap6wjTqDCwoCMSlirEWRaPMmZVJc/CEfUOkNYpIcvMZsY0u
5ofL7ZTCo0EgsWuo9iZ+px8DY3vbViUlas2BEQu5fv1jfqS5lijcekV7qHFdzMAC
p2DCPeQwZUyfiYYHyVRryX60PW89o2QRAAmevMVwAz7YHdnSSs2I6/aLxd6/CEmC
cOG2FLKtsOxqMeP1r26gbj+5hQBRqj+/1kWF3HBoLNnBxVrXIJ4/1CDNgtDCVzUa
GMtewdJBUsZdLm6xqdxJ+RdStE0GJJiu78w55lXjCptraYzN5fEoqbp0XswFHXIc
xPNTLDkFVk9nWeXkGnz+8a4HgLchsYwCxHj9AfC82Rf6yJB1zIEeOtxjwUeB56Jg
d4QQsTUMj6uLP/iV4VR4jz23D+rTGLuaFHCKUyWjj6v8NyhqNdWCiXl9ary0V+jp
iewjbVViHtSrZHAVN0zBHb26JNTT5Or/4yvqC4A9lgT+h0Z1WmWuQyX6vIu0Zbb+
sqn2pFsRILPD1nQ0/V632epbP9gSnjnhp1dZ7PXaRbVlRHiYFyfrcPHwH+goF2uB
jSWWhYXggmW7ZmzBoDKe0ikjUI8t41ShG4kVHXazr1O0so7xfPUfUMdT73z9WTHD
V7B64JGO6Y5WdFviXIUdkMRvtsMZST74ZzN7r6dOCvYlEJZTpM09aaNBXVvzLezs
WdHo5nsdUxQt0zkS92lDdctUNuRSdGnHOmToA13ekaQ5idjeRr/UY+LbKKRu8E6r
iAgYQP5gcHr46RR38cSuMIs9zHsl/cnME+5fw9PdKIUYcuypn7jF62CPBd/9dMPw
IUBatG515bNic9Ej+HoyULvoDvLem9Vb3enTrsNwVGlndeUg9x+FSFrTISp6Rdkc
aVbepHSDoT76umEXnMA/l14RjRHC6liwbG1VSGnn4J+ZMhi20WRe2mmd9EaT3vI0
izQzlY5umpzlQ92yiUpg/36US9AHpCWn6h5yozx03YtHlkTBV85Bt33NgOgcYrH2
gCdT6dnUcmmHdyhe2sz0EhQUjSAanTqno/J4FAiTWrrHggaRaRUoDryhtjQy1+EA
s5ylhUjfTOLv6hQvVKUt1mZZ32pZURRCav6hHHodnP5nYmhsspTl/t2oJi07ln8y
E08By702PcJanJwsYfeXqrEYqEeAbiMmoJXZAAcOvEc1DOAD21q38PEfxHEqxhbi
/dOIXD6nh2C8YBjynKWTw5azyy7rpZxM5gPKJVKFfm1HBlv6qSq+kKCY5uXN5qIW
Uy1SokSRVOdeZCkvKncbJZswgXZibzlNlksOzcOEpjj/8mMVCBrN2CPF0ciHsEgT
3/eQIZ9Gl1H35/DGnwKTKMTnPsMIU7F7iEsqWvug5fuyHn0CwS/EK9zVYcFt98Ot
k1DJzT1nGIdGv/knHHdH0r6sRb0DmvPRZNMn04wDbBnoVi/gfu1SvlQWRxnRoPJJ
59+op+v1wEm/5CkevSQVXOxgBGtdxob2sxVFJ2poqyZjxL+53w0wQPxn+LS54eD4
lV/T+natAFkhY0m35SCT4EMgPEJdMD47NDYXILu2JwL9cmxQoJKaeQaLTJMf9pxn
uwnkUJ6EQ6kMDOhd8xb5DDNYtZHb0oszc8cE3w5Q25RmvHhmlrEsz5Reje84x6a7
cXZTPKg5ZXdA9jQZTSh8mAA9M8lLWzcdHweou4wouLoFg7UaLQbYFIZ1wJXHj/1B
LMIW7YEG313IygQhyCa3xLFc2qLuASFb1ro6K0p7dV/22ybR+cvASP6QRgClHGLr
c3x9KsfuKUjkPaNBelxoAsF8nIWLYZb++B1hsfab1DMPNfcMIxMF+AxAO7f356Zv
LLDAbIS6FZulmYljqXH4MJzXyxQkKbbIQ9b+zEkxdNh8dN52vaaZ8LvWCtsd1/F8
GCwY61+CHwWIfgOxMsVEl4Hc2vW5XqA3b1HjoLF45JqUVW45EwVFvHMeDmDuJd7I
0idWd2vHZ95DFbwx0kpl7HfGP+/Omx2Cfes9AvVO4IqrwOZCV5KcxbXXF8y8+d2k
zBN0t13fRBIF4RqgLD/OXUnDAaHmRQ2/gU/t3GfvcrttvKz5PgRyak52W1uBMHm5
4PZwSJBJIL6aRYDRhSzgAMq8t8iPPMmZ/Jy/ul2EBkRBRAZOkZ9x+l+ch1Gek6sK
tjp8fHIPfP48MrKBVOQYJqmz4jZJACI99UT1db6aPvcVfT4W9/Y5D9m7MOv3Qqr4
0BY0SFNhsxEUfeAMdEi25/7W1ia+lmOmelByl0x3750Xjuq3SfYPH5jozUJrFyg+
CGhUThvMuNzP+zRIneu99D/p5zKUCkQvE20s2rWeTCtWARn9vrXg36wreqhuTuSK
xHGlGYE+dbtVl8nS4WY/2qiJtiOa3G6/ZhTVvf44JbmZ63N4d0ar39hKvTgH08SA
uSz7ZBfLO0pk67NdEZf+ocVsytYEHdPzg2XhjfmUvgmMwD6r/ivQRUIM9CwnX0gQ
3+BhajFqXcY7U1CnJuEKgH4g6cSb+55RMZOuprsL3ZI1dJwxcTmgI8Af/tu+5wBl
qOq33FpAoEG7RxFbT2Al4N94XNbw2YjwsZ1FINWtUkwgK5/1noKhRyX6Wm6u3de0
+6wg+hAiLTCVnccJgm3CcF0/jwfHr6T19sfw0h2DqTfYb3wo/uwgb5pFysl1QBab
521nAuKKLpiISjFXSLROeeV9GPK+ZRnTSeJCPvcqJ1ZhDvkavEntrU05RLvm8pR5
MfLq7AlJphlnvnh8SA13M/cZDmm+LmEGaJpskXPCUNfWmRA/uawDahE5FRM85EDX
y+bhHg+Cv+3ZtShj/7dYsku0h7MJH00FEAHwOCx2C7LRwWTUu1N/LZmcjUWIUh+h
wkYIWBBKeyXkJtBcyEKeq2QRfwSn1atR16NG+aEQRbYFtekjF2LTGN34AiHlJlTp
tbcJDpi27LBbMW75PahhsQhY8Mp+aZQT0aIjdE45td7Q50a9A3EFbx2twtLCPBUY
YeIikEjnUS38DsFjLOMSIwJa/TWaZsaWeG+xfWCqC+S2tA+Qgc3+mSg7iU9nuaL9
CNqgrXBSKPIZo/ZDbDhEoQ/vvZSrZglcYBK+aG/UyrUBkUe32q83dlQ02nkiXaGQ
ZF+5Txk4rgcUKHLrs+xP7gLt65FFM1u50aXrtyXKe9Bk2vi340fSkRy3vH/mTHU2
etxKp+aVkE58Kyuc987zDSlnqprdlr6u2WOjlSdWOxPttN+Wvn2oDeUlXGRQF1yK
d8u3Xx1bKdIwfeGJVRK+fF2HlCiF6cNLsrio1/oHmOJoqc5nH5x+8NdBffAT1OMQ
uVxm2lAamWVPDRFc+HrNc2hfPnAOn6WBwBv7eeBJWzNpKMxwdNSHOvnznUUBzYB9
F8YVALHKN2qDbuRR4EQ1BZaSdTJuCV6kVPL8fASUwHd0fbnsec7gCYz4OsUM6NcB
CeiqoKtx/UyFCaCNA2LkCQo4IwSvPWMIBY422xC3sVL8Dn+qSKD8wk/a7dHvCgch
0+Gmr7hty3GVAYlbomNDJTSTDfLE42AcSmAnfoGnSwNkVtdQtzq+f3ByDoKGsK2z
LADCsRV7PhwL2Q88o98P8KTYScT8VF9rAQNWqB98FB8Sh+7ZROu9NJEXESRwFUHw
8D9Zxvs/q75KHaH7krDQ7OE4s6x3AC87DTHP3iC6IjP9UhnSlHiXEdkURSNgdofM
A94gxkoW66WKIdBtRSGicILXU3k+M64ahPMKFQgOSvdFzjHh3FeNOYfYDhpoEg+C
DKYDebPTu208cQO8DhMICl5MFv6o2e0t1EdXLwmifsI/zAU2WCk+cZiJROYEmfO7
fmOqzyd2MvRMDG3CABYGNJeeuDFLZwJn/4bdQYLjhkNN7wTUZTjQ577/E0mwvBQ0
ttYNelQc2TzlJmcVSOGpT8m5vk4+DAqBrvb17g/a3hj/A9TPc6wF9zVsuoUkT7Gf
tRmJ5iL1B3ir0uK7gtLMI2KNxytOUQ9Q9OSHEGhYZpxJ68ju2PcGRe8qGO6aCCmi
VUk051T7Qna9b1Kv4cWTsUdPHxNdFDim0EpaWi5RsdwVNwk0fYuA2DPGWKKZT0sR
1SS/VXIGdZ5UDMhg95KVgPg9h7iuSjNQJdafmUJnco5oqddXX5UkjvEMHB2iW+Dh
vxn+pXh0RV3OeTMBCbvIbLGhtgqdGp/iHr6S4O5kqzTJ2rOrZgBTsIklzb4o7wtR
p/mSYqlZSMlEWYQW3mzIXO0V5cdHEZNFOP2Jo/eBMpUiHzVOar13bj7aBMDLsfTe
kBRDI8CCpx2+9peDk0vYTvly///IgbBle96dZSaqvlynw2XlHjh/79vC16zdBcAg
VRcXVYKGGWhYdXcjH1Io5EIWlEmMo6oLacU0MMtPwmYr41cvp2QGYGBNMaMLwqHW
CXaNdMs1wsFpvhdYmSKGjX8mDNbsGxj0ehV1IXEZ4sAgRvVZ4GDGftY3WHzTqk06
sxuLGjm1EFkcKVa6xWmbxy/tUZD8d3BHKlY5dPXS1oFrr0x4JSYm3bhK/J+JEV4T
4jetntPSOYH+BhhrtwN0mlomIM96MzbAThmEcskUMlLWu8kJ4xT+Oe9QbM+/W0gV
o+qoAwPzK8tVEzOpn4J9UUOpEaLrhDAPIgb7Wku+SPyBDhTXsSz75fW6B8bFSVMJ
kPwbmOdTZtbq++YOsghhhnWuD0Mz6GhDsY0qi2mPCpQDt2fpoempmwllJIHgDQ57
nLOPgFGYXH5Usrj+YmFiucv3Lju4XNUJG4oWRtyC8XaFn1Po9abwjqIeqjw3TeC2
StO4pFCN/GELUIJD7B9/eIt0sGUaG/H8M2TmA51rWWfrhUkAKpXy0OqxkCqhS44F
Ig8vQQAN+f4t3cXDTgs2vCnPxcM367xIDP/izswfbqNXKLBYZsZQ0pXmU3+kaYrV
w+GFsuF5tV7NKdFCyc/T4ri4ycCGWZrvIczNGWgqovBi1ortN6jiWdpCHH2M3J51
ZlvVM+x7C6oaL4BzRD3CurFB+U+9GxkE3TDtlqdA16kv+aIJQwOxbRX8e1ksRDa6
Kwwx19Fk5pEJhQI4IvuxYVSyrEdej4D4WJtcDcpeBny2YLXLZxJccd6ELgpKVrq5
u5uL6MMD5PgoHjP1CuZoXxTC86ssqiPAvL1oXXq3FFv+CYkwZoyKsDjaNmYLfsLZ
cNYCfkhoSpkz1A7e4Kb9eAhNwpigE08TPVHbK9sdKNPOs0CCBxTC9D3gB5ZjXK10
CPL9D9JIDq+nMIR4o5vP04yt169B+KqjFUL+O0k53L5LiOba1Mbi9PaWGVtvmSyU
y31hcY60MvLU/EI65LrX0/8Zx2ZgzYkhIgEVGwlEISGwfd8HRfo/KLr/C1EaCYWu
nDwDJTyWoSDss5mXm9Dbc+5rD7r9/7P9rl2v5o4AQnQoYDYKutfwxasDCm7lP/rz
E+9c5ey4qiUq0mc7g/7Lwgjzas3aHkJe7l/5H8RvUaD8sgB8GF45Bn4W8e28SzEd
2MauIpZd7Nw841p02NTNh+LAdO1lXGlrRFYE/P8JWDft7i2APS0xrZ5FneLjnhIW
C++RJPeyiToBJ2CmpmnQb6syQls0lzWVK0bMtXAIXKyFE368/sWeN/pNBFlJvKv4
GbsmKay/2c//x75dcFQLoJGwIgy7eCL/Cx9NBGNYKLfyS0e9HHrPKLVLTizlhjy3
EmNLuhR8R4EGqdkW9AkZzHKfSOplu6szROG78Lc7oquoq4VS1+y8mMRLZBpdL3UF
rH05dtgwvI6IMbyTb+kjNWvqYPw3piYCaQOm580ChvCpn1W55lIaWGX/NIy1/E3d
0OIW6U3Lx/11m68qrk8SbNBgYCEWRFEqaVIFkkYparpS0DFSaqgkYZwuysTFk9HJ
zIhFQRTsH71QLYq7dN5M4AwaF8SAX0Qsp/ac8zxBVuLKIi5RE/ueUMmmuETF6H4L
9MInOvBvKynfNRrPJMNMeTxelrjnwrURqPg8NnIn6BPLpWRYwYV5J3BEZnxAdH+m
LY7uv4fn5uYE2c5cexXHy7/4CEJpvBjX9J0NzedqctO4V6JvaNF1zUCfaA5nFq7l
ynIjbZzZt2i9v6u1v/hBkC1PuTrWVkI5UDLWEHi1pQQf70H8CWrhcYBXNrGNEJjz
2vsR8r5eSOMYyRJ9+iWqcQ3LdQQXD+RQSH/OYbTmX9L/zkmzAAhG+k8Y/B3sQxfI
Ks2i7bdgPe0QlGy8lHbZFD6EHWuhMYnrr/IlRnoLHQU11cq0NT5/v12Hj76ARXf1
T9lMQil+NWikuYysd+Q2nxHgyWZok3HDIw7lXGj7coDdl1LmQeGTZ3b9obi4kd8A
nxq4Ly9SrrdJ/Nr/i+E8fhHTIlTZY634xv7iJfWQTNP+fsdUbeg395Uf6jJCeMUB
KWIX4qFB5WLXH5cVQETgrt2gtToUaci0m0C+kVW1rDzSX2cdZH6jVi2OMmlqvrxM
NuReMfp2O+PzBv7PT1mzHqVLwQjHUt++OJvNlVXWKZ2ENX823mMCFVYUWIpy0I9w
0wGjMa8c71ZkBWyIZL9Ixj6/45CbYhy6fMzbwgKnzV55YfQa6UuBPTLMYrJ06NEc
Zw6cmNf4tZ2QjjU3jYZNUneVq6kKCehr0Yo4N3BDDrhy9i9TaKBBkHGNNZIlX7Pk
ILVFG5yoCDl9Iqp7jYqJjsCtCRkzEHySVwKISmq4nRmX7hJ/EOdbiOn2/B2QyoZh
l6z6XIpykBwHPc+HjqBsc9+HEnoFRS1/+awaUwXlelZIbV1zTD5EMB2lCBqb8KED
Uyn4WZJLTFtjBB2GflDMqPknftzre4Ueu9hvDUwC/Q6meqLplcYzIekj/u4DQltx
v6paFrkuj4D0dDQtD6Uc9YGGejhbkIERwW+exKV+opMfhauvDZ971U8wMEGwf+iN
OIbQtSw9KjLIDyMYDX0wqQ7OZB8KNB8cZaDOUDD08iNPQJInhf3A36LrOqZbhqM6
8v9qIl4Byoj5AAXIfMUFLAD+2Nfm0Id98Zt88x7xwQDFU49F+cnZmrJT9Fhok7W3
UShGghmWZVt2meMaEt075PrILHKc+b9Vs8VGgvsjzuwYN3x9XNU01G/D18Z+ZaaF
Urc4NhjNtpS4TFP6zuSm/LvI+6j4ndE5YovIHMNOJ3SWtVn1KHJOIy0KA9LUQ+Dv
omQvR7vBygWi9igMwtaWuMzzyvX7KtiRjPx1BIhizohUBdQe/5pGelEq2jLNesHT
l1tG+qf7qQc1fQ5HEZhDHso+rTzE++5SLnPWLHrkOTc+M6QHafXwqx7pR760yQdy
+sPn73sL1XnsTK28+3kPpR6bcIhLZkB8R7tLPxFmuQIa6IEz2ucexcEZieJE7XUf
SFlWCeSc8VsIQquUwh4cKVPaZyyywSihAf0jtEpUq+7/YAEXwxqhbd9nMxleonZ1
fDPW3uMxsMn4zgCaE19LFDkTVDrxPXRAxKChPcmfbh+0OZKGssocOSaTJ/wX9L4T
HI62xO3+7ww2RSV2XYeZxniSJSkqHOnhyOACHwH7E/TVEsveElL5KMyGsPXdRlzR
5/D9EoKC/ABgu9CFqJ0zFJFYaGV+FHZJfQPyT5KmVJ4351oHBdtTSop9gKl/pO5r
2LN8kywo+kLopV9gLlowigItHeip7ibiZgtF7Zu1pfcjqhez+YFoQ5Z9Z98hB1yQ
EhISOjaQVNv6HZpHxNjodPCyHksZOrosjxYXW1bG7gvJVWRmRDGFBM9VobT9g/1W
tsK79NiacVP0zY72UDW5+O4uAeNz/W8OZFtpz2yeFf90LuaWqiVYFgD8T8GVwquH
X7lJk/RCmyyNYlvMyUrf8osTVH9loeA9xDkeU3HtE2gnwcpLFQO8Y06Hc1KI5v0r
bwftNemPV3wVU/ICnOVhG6WclyPGG0EDoly7toCwU90h3THJgAFjdKv2rSr/TFMa
ymEdQinzSqv2f2O8vI081q8OBhDgRe4WxT86FRX9PtCEe4o4WEBEn5VPiYWheHSJ
SJjBjdrNF0dd/b9IPlEuWcpu/f2R44caZdz/O4WC8pJZWgHp+Kw+RbpgB/SqWOAU
CQWT2sL2Y54h/fcEsXKdFAcw5jxi/L7OK7ZPW86v+Pk6u+Zi6V3N/m3CfHg2TiPM
AwpLtVx6QaNWlnr5+QUQwHajsswdF0adZZ3YhaUbpBWHJWz3TCfBDJmtJt8Ce4OC
k0PZfWb448mreeAIGnA6KZ6GHlgiHqu6M2adDeVi1gIYflToa6DMpoz8NSdVHDdg
JmUKGGzPozgu15nJjX9wdioBP9VQ6vZgFKUXk6M2pEy+ijZ7Oa0Bx25UFUUh7hPq
y6aSZqzZhGHYakgKevlcNFUNMCUMbQEB9vhZDBxOJr4alSkNntPQYSPkQ6yryv3j
HRNV+6EB+J67vowEaOqbGAn+WuT8Ncc6st0+UjmdGhhoPDKRb8zUmCrFWVJ9joLq
Ye1IseC2ylxtI6XU8uRmgNVPzc4itad9h/Lv0eB6j7u+fJl8PNe7teBK1EUypfhR
u1UE9HYGnfi9z/DhfaS1dGQWqKz54eQ79KRT2tyHkvrUik7L/cNq5QzWe7hYS3eD
ffo6PPp4RftBAWSHNc7rEB4hgE/4d+3d5J3CHXCfVWyP2AVdhwXAHiezlJ/iG3U9
nVHEhFNsYaxpqfq5sMkYI/NyAvkrpQjo0MJ0wrskmh7UwDlj688PMDI8Mndwll3+
geNMq8FMRWjPuzY9tVJCw56CezKVWvuSn6SXwNz2k0BFwazEkC/fJsNl7i3JI24f
N+bKQ+RT0sSAtZ1rzh7/QaygZ/s00onQkK4f6ljfEDdGpicDJWNgQpwwn6HJKKc8
PW1PAieuCSGc7Kf1gyvxcSUUJ53tGy6wMwq2UIWnLNQll5mWmKdLKIZGb0F1zQvn
U+dZW/FkzGnpHJo4DIHd21H3yq3NRt+ftEZ05K8sjE8848tqiG8ja0Gv+3AvtTsW
SZbix3nFT3Dn0R0YcM6iwnEGSTBWHSKpQgIuxDDnuKNXvEkwkzpDIi0AJ4RYhny5
TukjzKwDZSP6Rljo8epgC4qrbho8YyCLeaTb1PUDufcswJs/ldA2h+O4QEK7g8uc
3DuWroqi5dS9IfJIWiocSB7QOohaRa7E4D8aQ2pOkP+uzueEzuRziEPs74v/aDNf
VdRAs2liL1UBcVuLkghSvjKIgSZlTcen9peDYgJ0bXjMtM7ymkkhCTKuW2yPqqwz
x41XrN88lJ8T30EOO8j0jUSDi6vBOtXddWPEAXV2YyMFhdnzm7DNPxclt32hShsx
ygFz2E+/39/9cDEMfJzaI0vvwHKQ+pSjNoEA6RYNFPsWnwxG6Fiu5Y6ujkBllnYo
TSyZZglTKXCKR6QBNAV4z2zW4kTXgqct0q/1a45lL7BkG65qW3Y/IdFFldkPNq5r
rXgxQzwJYitzLfHMJUkUp3UpXHZ626wgAKM60c8TJpnYww5NvDi6B/bDmCSCq/dM
7L2gFhYA7FiNolmFXfyyEXIlrLW7VmE8fZw6Lj9UL9yy/sE+/BC57l8lNuFdow4e
wWVLw1auGBZSHUwtnLLwHIIUn7D2rumlQ1K19n4pkZWoyNe1gvExwS4N5oLWlhUO
sCW5Z4S2DS6zmP2q5EsSkqOGngASABJyXv+DdnVEU6QKhc0NrfXGK4GxB1Roa5Kn
WuKNoSFluPG7oErGFDb2sqUKhOzSkg1o4buN6UCkFKJ9Gbd/pPoXDNQYpBnAz+RH
NbPd7qmDQS3VsU+D/0dfoc2XSEWtsr2IH+qYMMry9UYQuwffU4gvCAS8LN+ahHoX
1HlPIZhibGg4XLlQmOPuK+bHnrCzAZaOvDClvH0xjkob1UG3ultUF12c24LzUo6D
8j49GgUMpRH7xcsmk2VdrT9HIA4PFpTyknCHXJJNkFxtWL/C2X+3BuCHv9L+Ix71
CEFBqiQ4ASwMAfRc/abKK0fTuwLYhwMJYfZ5YqRRB9STeBNhRB4hO0WFAFPKzuYS
An33EoGt5581vd6w17bO699sRbwEX3R36wzk17WyBAY6arWGZEHD4k4UAwMe94hx
yEdeSn2x9ndsZ11B1UaBU6qhm8IYevBvdaiqCU2Gh2M+ZOiuGuBauaKoOGSElxmW
f7J37ItxZh1XA77M1YD1VpPQy0mNeAfF0/z9EcGoG5Afk3Z85oVRlBBzP3iPWlTA
8jrrLOpwlWioO3tP1Nq2U+HyheShsQGmsQ7vuRwqolyYxuX+ubHS6TjLz4ZO4TA5
fuliQK2irkT/kWJPHwZY6Y54KkC7c+aAtya0DKRnGjDV3W7vJc2b5yBnkb3AChBT
chyZ62zWfepaOQJwmOSoBUZVzhDjGggw6hKfKgW6PZmN4OpA+t2PBpObuKcgC6hr
fg7nEb/CLHe8FMYF6sTnOihimDGC/VaATVysc+03m2l3Roh5137i+Nq5N6nBwIrl
s8pP6S+B+4H4Noq6qAfDwiVvmwG2+zyRY0aoKz2WnOCpfTggOXHrLFtAWCH5kVey
gYbxVAXS2ILgOsRItLxZz/4muswLzmq2IHdxQM2jjiKEBzNG4dHzjucg6G0jns8k
zGBDGNFF3Lj38rt9XgkULj3a5g9pTEZ+3u8jmdr16iwkjnl8Nswc+d7d3Bup/XE8
NjFboE3MxPElsSUWr1mBGxhUCwsdDP9PpEaYtiDZahO2wwcWvIBejj8/sJnYIl+0
tncvjGfLNG5PhAkKtVNySwXUADFegRCyiczIAvmC/52EQCVjZohj2E95ky6kd84D
/8GiGYwZ+pcCvw2LYm0JcbDNpZtokdRVLp2GVhHEaSub87kvMqnkXknF8q/ZFRJX
eamOEyujmLBsOM1J4AZCSD7p5kDo2ZGYDRujxCMUKTN4GWPXicLZuFjNsPQAwkdl
fMEa/NraQFiR92ToOzBl6ozNLGhw+Mzdm9TGplyrOD6AHp9V0IjSizKpC6CUqgT/
PdHIATUU9F+6VU+9svaAvdGRYl12jaetP0NJc3YQFALPAEruV/3G1JaTEcMKTX9A
D7hCRIX4BVmZJPbTvlTrralg7Odpet4W+cMStR3Hu/fmEgw5pFYiZtD6IHpLBX+6
QDOqYUFoRTjjFpsNAjA9zY8eKNePCOoLLWyxV2RtUkyfD5QmliQxlJL2Bgv9R4Ro
St1k/vRZmkfxXJIj4XQzNJFL0vVBgM2f7ZzxYFehTJ1CCRSxGTwxJf15C62L0ufZ
oTqd6SA7e88Bw0G17W2OChwuc1WP/HWKG1yfxvN29TA2fzy70OJDyGQQdvpiApft
JQHEbeuBbTpaUQMNdk2lzl11+JWad7/w5RBBx4hfKAmCGmw6YrDeAJjkS+C2Jwq0
J03diRJAJN1OUoVM4oxI4cXNAJiDh1d643UBDOT0weSn4B3fXR/XMu9kBKkxAE2d
A8ybFK83rSC9pI0Tk+MDCLWeyDzZHN5mv/CkHjCTF3fW20tKXXvUXYHZlKsWY1B7
DJRttAbPcOQDRbfRyTVysOdFYSi+KuBPSFtl25MUyqY7SC6rrcBdhdBnIxeARWzS
C/nf7QqFSjiQkgwMSh/R3IipF7+HcMAXwVmVihFXFP5EUxC4O3lBLHF7yvNY6AcZ
SbtXUdMmw8bMC15TiGvL39C5LkL++/BAPlaluOxBH/ixGf0JWOFb3iwJN+eY5V2e
1+ytsaQIXPmytJlzmyOD2YS/WZQ07Jq5ZdOx0MtPY2pMnVJ7MaRBsD4JiOPVrz4W
EMCiUYMUUOlEjqJ+MG5OUjnFl/iJ/9oQMcYL3Keku+wIzAfTE8+FwgE8Atp9MwK9
hsW2g93eIBJSMiGZDVvHC5itxwVyaxo0CjIV1lF2hvISYFvmEE8ddHqyNHVt6MVM
iKiimoDvqCj604RpmPf1HEa207gGsRYqroCJP5UCPIx7BfiqBPJA4Y20dJ1bmMcn
vPAhXqEEtmEmpEnURttEhr3bnuM2+SBdOWzRVsgsfOE89Ono56fYAbHIoQ8bUZzr
hEHnvNKaI70bMq3A+ABLHGpzMuFzxa6/iJ3KwtPf9U5xNOjUkIjAxlb2A+JNfujz
ZVX7mvyYhhmdwIqiqXhXp81LkHEPD/iIGIiR5GZA3ofbXHRNgq5U2EZ8sIkZn2MW
ipgP/aQvTj3cote3GSEQ3kq9pps03PEUv8GnaNq/RkYhZVPwuUN8UNl3Hx2cTo6N
fLOG/CxnWxFbk/j2ffrNDCx2ryEGzNeagc4XB2Rjd876YxGaFNbYCnD4bpnYFDBv
cmIrVpl0c3gVIk1Hg15W3PWx/my//0A7FSd84JIqEQ33+jYbuYyrtM3tWcR8E9Hv
NG5CMeevBZrMbBksj2DR/E1VM+kFs9N6fdIqgYiglZhwezMvANrJqNSDI8+EZmpv
J/h4tNbAvLcLCh3BlkBI1b8KJTr8Iv2Pw1L9Us2X7lKwbnA+50hOkmAKTVePcP/r
8xvkBo/XcyLEcKcBSkrTTanrgNANxZiqSlgTUySyDsAlstNH4/bo1jt0AD4brepY
EbjqdVHcqvdLVtDH/HzQ6cl7LMwdM4S0sVo6MnqMQRzm7BmWjHvMsJ+cvd11YytW
XxuyqnnbIR/iMCw7m/t+6WOel4VlunJc3pVgSk6rgsDGFJXSU4ZhXOZZi9x4zCZo
MsHOyeRBN2tsxzWyKz2LhQ1mId5lkbPsja+SAPIvGgVKeN401tiE0scUcutkp+kE
NcxAKeFmg/nAOoRTYVskvRkTTfPRCLoGymnWuLQDmwtbVTsdDQAsS2gvklArF1pp
2JpO01fg10aOnt8WLXy4B82Q1OonhyUbdA94Y828UZkodUFfVKY0vyaZCSMRIArC
c7iv2znBGKbaijOcgJ3Qbt97/BTuzn5ho2Uhg87IJ2F1dtmDbhHKhMr0qdr3Jf7l
C4NrxouzlVyqknn/zs1GdgagopkfPg2zOjB3/+gIqTcrLv6821qCZ0lsSAfchc1W
stNNDqwUz8bKNDVMWvKLAHsddZFCagaCWL8CI8t4a9gfUFYzeCeB4RbUIOkM6Zf8
xn88hRTTWkeT7Bfu7sDaungosrPSGqDHXfRWhUdrCoZ3467ecwtDkThiOU8NnDfo
eemx5JXdrTddiqJ4sEjAo/UxW6u+RS6lxAI94w/FSNk1iLbnx+qTbDPcgD64OxlO
qK569r+5nOyUsHjw4xJ4sRVi1EQe1Lg3JVd0y6URUbI=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nWGbZoUFaKW7MuYbEliAdW+FRK/kzzA5MeX3012CwnrMT2z/m6Cw+604Zmsky2fF
yVGka9INURe/AmdjPI5qHnJkEEl0crNv1g3fphIM5DPYMLfgn4lmwmPS3tmxjZ48
l3iDxw3A5LQPP649eTmLNol3+GVaJuB60K9CRoBoNFuQzKdgwzhzXRaRzpoyevM7
W6hVyI7MFl+oxrYzXdYvLtpwjPln0R4KPLCs73vlGrEUqj/oMnN6Rp0ObShZhor3
ulU4aGIe+3HCp11iMP3lTCitewOojs2n+tt8ycYJBzopT3khg/ODKpgHf9gAGCp/
OW3y8g7iuUjJmEgONyHSag==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8272 )
`pragma protect data_block
OtXSwdAygPrf0CaQfiDh2k3LKccn5aMzHxFaUJoYW0xYLyg/zgY85ZMej7hf34Az
7C1bfUSUiJ5b72ZVNDls3J6d2MkuOWkpKjIP947c4YXN1bT1Xt+VR56j5We6aAiN
pRwPzauNRct88x7vcB/8PGM3sON0jlVPOr+iIX4EyBCEcajndcsmvy1jAcQWwCr9
gsI50VhhQRkqNSV+RHIjAj+N8JQNJxIf/M5PyDryC6oH2XjjZZMyueOOje8MGqFo
qWL3ozqSEKe4somG8e04WHI0wFJplQHvaNE4Xz44KdP0CD81pNNJkfkhTawfuVk3
IaIsSMD72W+mc0/UN9RZYU6KltIUtg1ecsQcuTrYEiBng5Nyqa3gdgWOX8hewXG8
ITS3sR868eOPSDnvIHg2s4qYBTxTsbE4Zupvnhn+AhmWhydbrk2ZqvAehJoJqJ4u
m+2H+b2tKefv9wv/N7ptDOQ2igLQP+HuB8Pv+eqG2fog3RzjUTH185NJGCvxVVxP
H7eOPl2fSb6op+of2/mSKXjAC9/o4a787uYJaqqg74fQiBgCjGncK7FaDIJz6GKg
yZERuiwVK1ePp7jG45pOWEVGnbWtYZemPeO2E+WCzmoi/UXmjZeaNCPIkqsPnklh
B3F+PLsWEAJ4k76UBFfPQUp59UMtwdCTPz8zAQlVuJOBg+qjcD9CpXTN7cEzVusa
HHqFra8ctUEkoC7TjuGNmsVWCpk8TpZVvG91m5QUFw819pEo8jMktDijskxTCZNw
Maan6nqZuF9ciE9VmWEGRaLeBnIUinmT3vHTbBR85CG0Gz6tHx407dIQmGmxaZ/f
TL9eWI/yhUdx8GALT4trPuUd71aJh1TFXRyFK3gp3tyzbGKh3LIc7UWVLOKrbpog
3zUNVbPeCzQlFswYEL6IruUdgDjC8mSPOR339fWdM9WDmARjeaoWDg7Te1Ds0J9h
vpq9YRnbWCpHJXj3P1KOkfjNHxliSZfCZRZdOSRBNM8IomYBt8LkHhZ4Cu3qJZ/o
tLhBIP+cx9UuO0cukFWwF4kCnYHHKE4cm7xM6O5VOC+I8Dpsy4OMewTUyFjqk1mO
EFkaqdTZfNaHFbIoD/HYS1QyQBwPFtvBUHUJHXqMheWdyLYQsQzEQMMTPZgdTYen
Z9bBqtmdGOe2bV5jDTjxC1KaEem8tato7nDDOYTRrAcvQF2L1VNhO4/XE1u4001v
dXLZ4QE36HH67dQk+zUUgCa6hnt1MxyrteqrQdbog5zcJHQ6Kr8gRhF2uX908FNA
nNMW/ztpd8F+BvF8Jv3lcxjuyNZFoL1YkilguhoMIyoGzAarE0+yAfBrjlob92gT
KGmFrVzj6gnv6ZNTckVHvDbhDSHu0qG0O58sH/ZAa/NSk0K/1GBwgHcaCHPFoAjQ
dT/seR0WlpCNHP0/VeASSvksLscMTXq44K+N4S+wLbQV0YN/Ns8Dd9qC4gZkhb6l
ysBlDcisUAT7CGtJJHLOp/9D8n1VoDtFGUdy33umwrOPjyPsibcl7rOMMfRa/rvv
EQthN29vCqgpIxena8CiTFP3VPCujinCQ5cjxEQBZVegYxi7ynC5q08ZaygJieYn
NJQllY/ggxQm/3rAxLETX1SvszBMmdmUODSv3NLjHvOLEh0u61gCDBf9+qbr8yVf
/QenTaYbya3TH0m0WGWuYsuIuk2xaU+cV5G3bnVKGA0XGU88fTisElz5WQhJD8zP
+AKuJqJpOlIWZI8j+7jkMbz37Y5GcGHaD2KrxA2zZZ3jnD5IWCEKjKlnmdKiHGyO
ynLJ+TCHXyMs1LETMBt1vhYjHI9N1KQnpcowqQlryNk3NqW5A5E1sK7nfQPaXKw8
eVDvyfD1u7biePv/Jo7mGnl/NudW04fmT/GSOLOm1gBX6dEpTLT82oBVi/4yh+Ih
3n8IuP+4BfDDBJwtc4Q8GE/rooX0uME1vYfteNk3zBO3HRkNYE/Qr2/YlNtvxbP8
SBrTHfsZvvIFoLG+EqW6xiT5kv77zw+BCO6soyipwM4ZdiykUMvlX0iDCR8Pexii
q9iELmxiEPh59782VzjUg72jGZYwPhMCmbzYDUXQys3qsUr8ACp4MtOD845RL3Ug
O81zBWokt4GnrTkofJRcA6aNWdhZleRb5i1X0iNEeSz722Am/zNgspuO3rNf6caI
ra+k20wd6451dAnfmC2KZ9K7a4rYYQwl1fKrjoyZNPADnfiiNrbJ05dGBY/AMAHs
3sw+absmAOBhZT+By4NKLuz0wUUsJ4h0nzHO0ngnNTT+84f1AUn0Fc4PxguihB6I
GrSgpoCXna2mXMWgJJqcokhl3GM9i/QPQY1FULUso6PmppNSKXMY4Fq81lGci+WJ
lWjaDfo4CfKEe46Crj3auwAKIMWzP6Emlzu3FW/Vg41jDxlOpy6h7m9UAvZrHWbk
etsQ9eID6Q3nsBYJgojzbjCau5ViStZW7baw6rnqE1K7roDKGaUIiOjaf+bifux4
jvav8pXCiiHKJ50FIuN5AP1Y6WKN6QXF6Htqi+BEUPdfRegLeSVOEI81io85M3S2
sscOJM0P6cIubtLsTYs/MePallAJM6qnPa0huRsSZ0eOVJRPMcmLBdaUZwWD7Ayn
UXWZXYzG1KMO8aeu+Vc5RXOiOKSD25zcFx/kcrmwk2NJxuAEtVdslFOgMRDq6Ln/
H0ctk83eUur4wqc/iV3u0dGxpOt4jKI6lkq7fuc3Z40E046k4WGvR0VaKxp7Xa6f
4JX09Fi/5RZiPs7fQEcif2SzDJMn963nXz8nu6e/xv4I94hRpuuTIf3UFOze6ibf
aJ8WaxBV7cR8B++9KSJIIhWRZ6JApILUDYokZKVKpZZhXBvkhbSH5UW7LZ6EXh19
Ufq8UD40qa8lM0RAOMPIKTyAKBZOzotYs0O8CChcs6W4w1IBa3vpBumsQ9laVfZR
CP1OOrRj3nmwkoWn+ycZ+EhooaSNCWfATvneg71Uh969OT7uazQ8dSkt8g8aexEN
7vVMG+peO72KIA9XwSawRPqzFJfFl499uYvDxzikM3paA/ZRX8UnI9mDDJWrwOdL
lCPTnHi6114CssK12zyvcyWwHLtWOyHwDDMaL2Lrxf4iAK6f90PpWSHQHxswthdu
a8dbeuyAlHesZjtyw4PcScuyFpvpEIuH5pjT9XxOCIQrNvytZYU7JXIqL48YQdRS
ievLs8JkSoRtj8pnYXPeRt/ts6AU3la6OTkqZdA8EemqZvMrROxcqkogNgrPD4RT
ZmZS0/KxXOs+daTGfGhC6hw29ZknA6YZipLAPPLHSrDV6TdIQfoxNTP/8NaYmzlz
GEV2ByuaGgtcT+LkkBW9OBhWlm/Rdg9gxhlWxTBBekAGGezcJ6xOTcr927MExc+m
xEmcPDwzT5S4nNwr8pxj/ybWb9lmLssZ12/0AWJAgCgOKotwxqAPBL09jmhdNIQ1
NxmYn48R7PXbiM0SRUyYPB1hOTbYLsiePZIC8XO3cNodjN/75j9kVymU6QrIzAEv
kzzZPkx4VAaJ6j6W4/5UUL86nNSqol1/MxMu5V6aAd2fRLiWCSrPuw02AfPdPA0C
BPjg7700Rm07WxRjDkgRgeCjf8mpCpLFhX58gmpSx2BmZq0+mYSggziCi5EMEn1U
TCY+wTKUuAy7WvVtvdyBukIBQIG5s2/vkw0w/ufHUCPcoCH9qpMHvR6tsC7IzLQE
AkZkKOR/el6AyW0y1ya7v7sqrFFiBZFzt6/1Rj8nLV8I58jEuCnemhu+9yyAFZui
XzYILK7h47x7Tyhqdv4Xv8e9o6sLZ76ipIHd+iWYccKJx7lu84dRJA+1MKW3PicD
Yz2btRY524KDZ3zxWf7/KNzkDtRvpJSQWYtDliorIJM5GiUNccZcz3bQMjXhigtR
fJv00PjfW4pQe6bx7Djx+Am6ViUwH3DwRz+3TY/v7b1J7C8CprkOOdHYxw/benNk
LSqhvtPC1QRX1LcH6JQ3ArVSSU8kOk43zb268LrqG4ZDHrt4MiZIZzc3V6i1ezJD
UpptCXOfQ7MkBubzfddVChI0EiSSMo3/F+K+PW6QPoazpPVWuJdRBGB/GMhzKXtD
maELth5RXOua/WDiSdnQ3Fwoas9Oi05jPcRstnQel/cRHurtcJ6/7UescDaG0LCR
ce+6T/jf5DnaFXd1DNVZHDq9LyXBFAoSKk1FbSyFB0/O5Uo0VOsz/tXABsadhxIH
tZJAhfRLJEwle723mdjEFdy7gyN0s0jpoiTQvSz3WyT336NPsu+JNtO5ZpCyeD7J
3FKU5vipEuwJVyyHjl9i2RMAUqxXMOtJkxEKDQlCGaQ3juF/GuoGvqrq3a/+vDcP
VVEXhbymMe2ZtY6YGyYxual6Skcr5NiD7qdR8DE8MZolvt8vMWPjcshwFnENKTql
8s6m2LHQcQmgpzoch0KebEpfew5ZVc24YizrStWsjQWXgLKqWfgctrOJWI7gqlS7
QS7s/37C4QGjNLDlbA6uj2JpFhVhOLfNouCfceHq8o9T+I9fX8EwsWSNXLUuvHal
TA2PrhIln1fylTsXdVXB6CHiPPkadzLWNbz8LwNQYBMxie8wj1QbslH7pjyQ6P6B
cZT5cg0HtIXUXk327BaMB9AXvaJG7f05H3qkZ7TqUmyObq+jQOS/a4/3y2dfunhv
0+1WxsddtPi9PXtIc569GCpgdprq5Rvbt2g5aP9ziWcW/5I3k1sld2cUPnuwyRAy
LhhKYdbSMFsyckoKdZRzpaDFgjj1/FauakM7TSmap6E9dutgxM28+FgT6iEV3Ieb
DYNm3p/xvYg3YRHCRj6e2RqZ3sJ7mJPW5lW9Ywrg+2pn/hs2p6XtADRLXCmD9KW/
OGF5yUpnLyh/P8XZdBVmiuSpeOymcJiTlMdIBGyEM9rVxJNaO7YXYeZiNwSKw2pR
g55VwVS8+SOAPKxx3qZ+XOAVs+BNAHKm6iH4NN2datCwS/leUIo3UBgQonGnt++7
03xLYTZpwo+wUZ9jW1oQqJ+c76QVEUmCM8MW4Q88a+qSnONYvCyJSc4cJinqYASh
YbK3xeD3b3xUHooX8XDT3f5p+11RzIPPFM8PEC0Bdq/kvLyYWjlmIXyDAz0VdsjT
HpZB0rYoY4LFPQMGF9XSQFuJBuTZrSOO0/Kq1J2aLeoxrGXpygQzXCsXAwQ/3k4T
7doHI+pomPcxJOPXD03/NGtHEJVBpyuVuXYJAsaRVY7+pPGEFeBYh7j7GAtltfdn
m8LdQrf+QQH073pIkw0SU7q9H0YnArt+6D3i4EEd7eRLeMzQFpgQItH6VVu8hynS
BRD3WnEfm870cey76Akg1ZN5mOqK9u3VrdeYWOeEL1WmC8bi5ArXVVx2X+rUBOIT
wAdIT5yZd1h4GrQYQrZOjIhzvLE6f9+BBH5B6FyMC/YgKEyXdYTIRyogHCq76zDA
YMuiRi41WBv2Z/YjblYNzxohqh2Jg6RRFjfC5eYftIQ5mL5xCToo+HCf5eoezuEV
LiCYU0tfJMquVum7zCw2PIET4XMhKy2lvkmFazv3879InR7/sg8NDexsaZMJZAU/
cD5b6+7ocfBqdsrUc+LK7MYwwCkuv51Nv8oUwXKyJoIkjfjsvt5vfdGLIS/XFPg3
WCwSjFVJb3SdpQiLnY7UXAUpigIU1rdrmJy8BzUYI4M1T9HwH9sJ2mUT/ad9CTxI
YjB1w2OwjJs6PGorwNFfVqpZCPqSrybKzSscTxT3muOqQquP91LDA7F9UIICvoAn
Jf6GJTRMNhx3qNEazqwUKVTD1raspjU5KUe7TaKeQ2OdRRzw89CzyrYPA7qtWWvr
gQzlcWJ197J9w/qd2UHLGAo2jGoe4TTISuf3Ur0KmwlrYOIZ3ukfLGB1ddTtOWWY
AGETudgkD7gbJytH33K+656/ITkegsrJJH8DVJAeMUtHXlf/SMFXHk4oK1aJrNe6
E37lTqrWzWCRws2l3c3RibRuOy87kXDCMak3SoOB6m0slr2s6K243N6/m8Twythw
LxRORQPU9bDA4e+Mxj/f2ctxSHG7RA+F2uzHQNEGlunU/DYDpRYWh/dPwqEQVNdI
RsRtaXQjbfltCVmaV4uB1ZzLwcmAU029uwi91FKmnFLUpcWes+WpB4KH6qy3L0TB
zc4Kt9YolbBbRQYCodrnAoPSN+HkuL/FTaxRHV6d01HaU7CQVYg59nSgx8oxyJCB
McZY/7lb9/H/6RkBCY7c/xzokkIbw3YEuUSjdgDt/sUXepZT3eRas6IvI14cqhm7
KR73rVzEvs595/BKBBshYXrLwTU5YDMkytXEAONmFqOkVcMcjBpkLU7zxKJ//y0o
6AvbmDnL+zPUMG1pr01qbej0Yh+efd7bw7gKzEf3G7YdnsxXSU8n7C/4qUmjE1pd
shi3GKjeEWxy+P1V1O22yo5FTTZ00CP9P1sNfBo36n4wXhf24f916VczH2QcbxZT
aAxR5EfY99FmAl5LOPvJV9ZddBNTObjEg5zqEL8albPxQmwhe1ifuRtr4qPfSDym
1rJaHrKCqMjdcpjyue8RWC1+smyBF/0ZHRDMls7ZGDhiS7A1gqzUfj1FJJUZwFUU
5SHiVORZ713gtz3eT3g2+bYsfXmSSB2iAvwGjiS52gENKoHVy4pjQ4FWmu6SfLES
xE6mlv0o0iQ12BRwvJCwqXKzQrhfPCpg3ml5/PGH/ax6HvkOf2+Rw6GOyhsVJfND
iy0vUvk9Hwc7/SnIQf6PsBSpOj1pEziFH73huAhKJeVqxsgGhp2FTnOrZHKTGb6d
8DBueeV5025xUGz6lTPsqKOccMrfC6vOpT00ipPC+2ZG8JjIl/hDwBZWt+gKXLPZ
YBRwxjKv5ZyowNAYkLSKse79oEim1UxTwF1qBIeBBr4vGRYlpqpeO2asPJuTi6aV
U4tNZwhhOD/ATAB1jzGRKrgv9L+XSVxxhjLsw50h2qn9HMdESQ28j41ZLv/A8vHh
WruNwLcouj9iTifMpqi6ryMMyMnVsLxo+IC0d8ok17p+Ij4LtVG+JUreLU3miHRD
bFfqipFRJUzCOIII7nR3camyuCXPHGMb0S/0xyL4V5y7U+MxQC13Yy0zRqw+/qQJ
J678io6ephvIZCVpS9lVNTgfJve+3meg3ijC906HDvFOBLPpgbgHHf0fluPPswGZ
tJcyhkkzG7fn9xt2B6Crwnh7pPQFZ+euAd0u2SYHHGOkr3TAF491aTARrpqpwQkQ
8lmR2+Egbwp8XtBiIoeVIqze3GrlhFa0+SRvHBBat4kgpp1xENESqkqfdrHv2rt0
2W/ezqhem+Vcb3KZNtAGllF8bEhGKOVwqGcTy/Ly9Ra82jzISjK5F9nnLFDm+s3R
8WOUjCuXPzX9T9wyLPNVGxhFQv5Awc8c1/uY2Z5PAhD/Eu/wdTQyX6kjSCP6LcmV
/x3Y0G4P7niIVBo64xvAFsFGIL7TNxTWeGIYXZC06fcJRY5m8I1ddKsT8cKIz1ci
4ojDkAFzQs4v3kSNzkkVV8cl14aF6fEkpMODP3GoTtFdrVr3JLEgdFitiXSCwvB4
gW2Rsd5KKoOKyU4PB2XCcIA2/beh4+EqbXxHjng8ZylQK0sfJCCVFr+HHcLCDS/9
e+LQqedrwiMY17ACEMldiETw2aKiFRSSB98KbAMLN68l2etdMPOlbJeAkSPM6RWU
h9gHTyPEYesNiez/OQHKMH+wybVqtjS+Ux+PrjZjAYsY5CzdsGI4xyONdP6Ev+z5
MIkxhPv/zMtlpjI8WBuXfnNY2nmW/cfHeeq5jeBDkMQqYINqQyO4I7+EE7Aud0eN
r0uIRNKiwN0BbCkESNp2Tw5uIgLXnVKTVproBSwGnd/uOjDTyXXFeMHHqN2Uv6Q2
ewielIIHNLzYvrFJXlJbPedy9LimItxK9g5a+xqMfwOXzlnxfIdk1ex3r8IfCreP
AGW68WwoYp/JwypHcP4CSL1wKZAhqSmBLpQ1Wm0tNefJ8Qg7a4DHwcpGIZWWfC8q
xN/yu85XhDSlVIn8h+EeXb3yGKoUYt7+95k8+muLmGl7hV2LHDd/Rr1M87nOjdEH
8rV81qIwPy2Z7nTaEI8IyZMq/Xt8nqhgeHPAhsgy3u8/qbHv8WKFiQNFYRkmIrmY
8A5hLDv4wVjqCsvZyLP7e6qnBXdHY0ZEI/zeWylStc32hsXvNkbGHeogp9gIWaHr
iTFe26TfVJ4hdncAdvEwZK4HDVJQwb+pZC2Qb0KPiGbXIE7E8bGG1bexhp8jhvP+
T3SFySn+dz7lmDsa+lCTCGsuvAUu0rKbVQytpVInKdTkRzRGIst3wSMAkGEoPcnt
iBQU9NYlnJ7aynnHnB2G9sc3/aeO0BoTUDg0vsgdbKTD9426AfwXuv3SHfb8RDBe
Bk08Cr2fHoNegU5XW2IvBkSxtemHAcwuLM8vUfNZHGtACQecrLa93elolGiIz5Ca
W2v28luDo84Q2raCADBfv1c+F8PugRII59opK9qMStXHaQK4jttpn3sKIczLXyTF
9KFB9+tJodoqO7N0tIfXDkU44PM90xPkwPyFaSv0wlTi0s1JJqSjilmkq0RdR1RV
i4lNyCz0ZzRn95Zx75F+Qs3wcUrT6I/W1pYjgblGxD05WbyFFgJIWEYMsu7KTQgQ
UEl6w/Ykl18ECMX4qZSHsZnNIhObb3Kw8LsI1IwMS17NVDl9J/SJyrPwLL3wgFYW
r4loqCOpQ/l/SBZsugSeEgCv+Z07rNigWfwmsrI6aa+4Ywmw5cmV2y2iiTP+RAhF
qKTNB4xd3rg2IhdT04n92KHai920dzScjRlHMRk6m0WyS86/HGSyn4B104PcLxrO
p0nZ1roBUwj0+zfOky/9Wz5DcrEdi0TJ9A2Edf4VqJBr5SBktcaEThNxvpI2BKnL
5ut2CpJXxas5mICMlDaJMHpEyqs5d/DJStVXc2aYB82yxIcfWZ25Vjfkm2kxe6D+
+cZKlEH5sUYUKN1CDseSeLJZmK2mGVuaRvsAPPftBuGJ8KMcvnPsPJ5A2CSKx+j3
TztA/0/mUNIgj/RzYrrslxedCME3qMSnsMFGf65vs054ju0tgEyfETeUbQxuajW1
BijtoiUHeOemocPdUiOx8vVSvL3lGsCITS7mtDqWxG4x2qLA6rVRmYNy2Tcj8zdI
UosDI5Ph6MTz61zAOXiKSJtiFyWEnQb5sJ1bWwuLXmg7WRt3kHYxD+Pr2UHCvrv9
cQuCFiX9QE6KJK4jZxrK/UUmBSF7FYBnt/Wq/gPBk6W/OdY2SEHrc339TWP3hJH1
QmBJeY/1eGN0AbkVaNBkrnefplfI6juzvVLaJrHaqK4qLeirJlD8OojQl+ey7jWO
zCr3MHFzqcyiZoL/jdZOtyyBjUUZLDeGYMUmSkcYDfD2QADr6A5214JMbPIm2e+A
BjxFjHua1AZJKJqSWqSm7GxZ8mquW3IvAPQ3v2YBjQ5vHLiA+HdPLKtuFL/m/1OG
N9+WHZxgv7DMT2LjPbstRx2AdOQ5PIBeDvRd0KVXydZhm7W8Zwqm3eZ47G702DRt
YnWBUPk4vN3iIwhQIRGT+s/GdGO/7ZLXNPxOgLALF4dGg4pY2mkWDzaZouC2uFT4
5fQ07viWbhjMg/uzejZ//ovANqNHNqyybDTKO2bjefzepz5ce5HySy0CeS6FLU0q
LUVlq6ZWioRw5k9W5nfvDhqdtRWtSNg5e9PjXayPOv/7mNjxL9L67D5PZ2nd6vv+
SBMaD9Gtg/d7pvK98OSaAquURK+ynf2aFtAacJz4u2unET/lRPbByxhqqSN9/Ssu
6HidMr6WN0v5FmE6XuTJCtoV+VSN3hZ8z/L0VHv5u7AqngwziTuVbSSVPA1e01lo
V32Zrbaf62Sh0lrA0EAFPYii5RpYMXySQGnReN+Q+Etco4997RpdfSzXjrlxZIEQ
M8yZMFiFwncHm0/84X4lltIE03l6QKE6TV/T1rgGefCl0dgD9d8Z95eB7j6toWy8
3Un95A5wMK3jLzTQuCgb53ZoV1GVARaHBLKHvAseuSOLWrCqYAC3FdQI+5afdQaH
xqpxRePtUPZ7zGDwEYnNerDMKCtjK/vBhByzoMzDayzgSiovkUYF5FEOEwGJbZKp
aNc99u9UY81WonPCwftnhKLRZ3nQDVSURhgdTUm1wzXErykMGtMjyIlOAbI3a9BY
kcBFC+Dmg3SXkqnqcv614DHYoTwHjtm3KGLeHouLCOcB37OcoMxPZRlypvWrCgx+
q2iivyovj5ZWoPqtD73O4xQGOzrtLgtlw9/N+7o1iUmP8z+qCzjNnL3vlUGcNnaU
JccpSuAeNFl8zHQxqHUZQBz8ThZn3rk9jsZvYT/zNnEmTiB5ppJW27pq+FLTpaGj
p+uCak0y0PYFcjDbFsR3abviPlqg9YSLAFF0vNCp6BQFNPiDfAzv7QDkVNcdMdVw
HiwqqlLNDXRPIauDi7qQitLJkP4YiJ7GqZVsk+9+B3xfFVAXoQ+PB/LJbqGCj5VL
sI5ikTF49C1W+8PVGqUF/m8PLPUSgKtrWQG7mVC/yFMSV0Uca881Sn4KiENMDffx
nJvVZ7eTgVLv+zerlCE/eIfT71xjGlzPQrRyxlkw0QoHaZKSWxOTUp7nsvxonotK
mUNmyUeooLcHJob22BPAyCUSHAB2iWyy9Hyhs4O27Mpu/bTr5Og0//4UW1f6tyXc
FpA64qrPqp9v29OhOVqOkZV57jegJIrSkBjSjM5e6UBE/84F4w5u7zAKyFtIQ6YM
MSAeaXtwRt87PQytttbjo5tr9KvPmPF2yMXoIiMIeyjsu/0ZrwYpFPUdXVpppN0z
l9l3Zmezx4lgDRQekrM4lKVi1dETPu8HBvyJ0Oo6nj0GoNoo22BwsF6e0Mvx8Frn
6VD00G2eJ4OjQY3fMunXaAOqkMAJoIv9ljGChwKpJIZ+Fwxl7nvZSpnyN60U3Inl
fwGRtpsbaJwR5p64NgapX3+dFqZTqMIlqwjIIYwlYHzzNpGjWjf8vjAY+0FS4Ie/
wLqwJ0qCJb3dQiiW4vuS0Q==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
c+s1Bk0lQl0Zob5+ndEUuHavWGHSpjg8NsJskMqdbz/K5heSg/pzc1enmorJbDKu
tnc20HtYpQ/4lstYpelK8B3YG7InjecpAtDrX1hJCjqdg8bgxXBs2XxNYdUXRucj
JLFiQ5/OlhX1UeL6wqEA5CV4n1/kAYaCoZenzM7pp9KNj5XKlSDyv47B+WFDI1fA
LyDg2uqjGCu1spZ69N05BK3xtEWVj5vz6oVNgskDCVlziDmMFArnnxyd5ZMfZjUF
OUlfDksRrX8g7igstDjZgfGScEFyySFie6Ebkzdi/OoUs0nQ0PS1jbsP4dfAKvaE
5u2V2tiOx3GKyUzh25jQ1g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 21232 )
`pragma protect data_block
oHLWCBAbpgcUJb3Pv0URRydqMfk4KbAHtQGJZGtnnNGa5K22dI7B+gbTVbTtBYVb
/6IrWfZxiU0C2Ksz5zbtly19fT2ENW1pyvjVq+u+Mi5eG7CLf/P+UC0dW2M2fkuR
VmXba41d/1pWeeeEPu35CJyQhoLjSpiZPIkR4GKPzE8LHscaz7AsaXPsZOVTqksH
vW9nqCX4i5ceslSaW9tQ79Zd1m6o+i/YOQcvXiDONPHQ4kFlqg+QSby5PcwNqnog
nSXV231h6fcH1Hf85GvJZ7CpQI/pASzI7o8eQcI0frlFZlS3HBqWJGCXWX8nS7de
7NSijX0TYF6tQa2xwIzaf0ggxC7AJxfcI7H2VWvWQymo6OuhL0X74jgBCVQXqcBB
okaLk8KaB/H+wX9bFnZUFMhHB6/8SshyC62ty9MdQj2EcITp0cn4jlKxykySSrlZ
nHEnV5bfGEf1fHuJ12/+x+XHBQ4IUh/4VySkWpN/SIhVjJoZtZs/NBappYvNHBUb
rFTlFB59d3T46gXQ5Y2JNusDlqmuvC1pHqNRtSPIUBk5ek2julC6nYMrsF1k9OxU
fpJs+ekjlsPIW8Dd8DgJtwfq6uEqDqJdpmn+F/scwRFfuT5PCI7rBb2zGQ/wwQ8V
aKiQCzgWM5aLNn5w79kUpqvjHrdRnsVaHH9CnsEIwB67BtlaRRQ4T57XsjWwW7Bs
zgWu9LyCAVJxpJ9S7y9fBTVOBEgkiTMzuXxXY+8nICdcsIQNDM1CMzWToGFT2Wzy
dsWgfDJPNjhFE9AGYJf9gMxD4KfxXycIF63nOg9FGefypW1gdM9WdMYXUi2+v2XM
R9prDgUSaiJk2ZJxOt0+31RyApxF9WWUdHcXpnU3WijeuNu2qnCcTKlvG4sPJEIM
tIYC7kBuBhPuVB086ZGBzW/zGWalTo/T5yeFJRyDUDb0z0zAR7tNY2YoAYriF+yU
Mwvoqz6q1SEgGeSm+bYYhw3fZsK+ucIvY8fzbXeSAvvxHuNPKDi9MCBOKeLibd6r
iAC+duqPAM4BiDJ8veHKglAXqhtrpX/R+1G1Ktl8I5eWjgsVPO2yccW1BYWpbAAQ
f+SJakzttEGss2h6YbCWF65ZHtStjPF1fuQfiQC4BpX/2tLB6VphgijHYu9XWIps
fX3bFP8q17ZhVJyvESlkTsO+ZzssAm10bt5yjh8v651mjrw7wiVhFXVF2+4Koex0
pWpzwp36OjWXbqg6gZZgde7j2b+bk7xg027tE8BPP2waemUb1DmluHHhd5IRLKgx
4opzEY8EnbTaVlcdd6WHZXNt93H9Pg4jeESJJxuwlWEOxOhIG3vvgSXmRcHL4A1r
IKEXsbVyjrVl+7udz+8IRS0YOIWWei5K8dqNBbz2scQMMZ6gu/P3DjvNyzBQcQH9
Z1eqwpKSeIbxjoVLx7q5C3oheQClKigLpwN2TUSwQvW3QoJN+FbosnUnIHC6pZx2
e2WQjbOvLpj2f2gTZ1Yj6tBaph1EgmRR5RE2kN07ZNlre7ttffwFoR85TJopRqJL
hS9hIdnrL2BcLGopymWxogqhvv6aZswH7CQyGqdTFN9YR2KokzDkRzItiAWbO7YK
YtfgyY+odRkjcABwH4UKJ/VCif85xnju3bMO4wDnjQqcqHOUJeXMHXTNImrQtYQ0
UPKZZr7vQ8ie/mIRHV5P2b1SyNtkwYOuMWMvOyg2jsvFv3P/IsvH1GPJ1vTzIYjw
E8eA+z9GgcNHyvP3an3o2qCUxIfRvH16Ivl2lVKtUMMXoUFNluvs/oXGE/DJpKd5
ozZ9MsKyYWkxApAAYCUVyh6nFhjfitGasEYZE/NcJa7U4bcRZ3e4RpiOoaSRu4zt
i8dJgKUBJ0gEDsztjlgIn1EOR9XuLkv8lB8dMlFHtKLOXiP9VyBBVWg6zCDd94Tt
01tv3+eBFryhX6X9P95SvWN21cSAFZ2st2mLlQEo2XyPOJEcKEJyDv89xtLe6+C8
+P32dCG/Pq0MJF/RoVQ9LJHqlEORrCrGWKdK57D2lYRzoGGcSZSdGgITiXZ4c5t8
WyQzionvrR7JbOHa0wETV3BPAMdpoLfbDpTAbxqMrH/pYHKvfO/SYCAIXhx6Dj1i
O6FntVe194n/hvVJUh7rcMG3HCgK5kt+fLainPiwwGuoXcCZ2aqUZSKKtFq8O9of
axSz/18WllFC/SPrmimKX70kN1kokOALW7XJqWteuZkIvzUs9RDjQESXsn8WXdEd
GV9FCak2sVLMZom+oGnRgEMXav4CVnc2Wp9f+HztDVXnoDi3sog/jtT6HGRCNImB
V3Ab2TSseEK9A2h3tqTxAyMJwVykw1MeQauRa+4h7Z6Vg82GvqSBvDtJhdtUpwE0
ldvqPGLBO0nh2WmTsgdLf27wX09GoP6Wrhe9t9VM+mL7QV+sToufeYkd8vX1pAKK
EIutmrsvtJ3tdrJ4AtG1U9mz4CVoOFolkfUQxEmvvHL0bSw3qcUlAXrmHKEbTu5V
7Mwd7UokNkmK8LN9DpFvOKk1x6GuzeEDaRbrkRMlkytVDaM+3Y5JO3+w5CqxZh5g
7VQN7c1nw1IaC0SoWjTiaOhJk2hk68Ki+Y+QVusiePudcopbDPB9Nfvmv1n7bQzj
kitsyovCLCroRjVSrO9FGabW2wQtoGrs+mmNAuQHTUSAcG5SpcxMnNTwptLjx9v+
sanHntnt1lpN+t6HBEBBqs8tLySaNzy6/dhJlwBfxQ+moztU4tEWe7l1YsroHbl/
n5dLR2uJfqb9M3yzKaavSxzJ5y5SqsVKDOy+R6mwE2aFScwVrj995/v2CUk/gCg3
zLroasCS4WqpOqU2DnAY8ZvaKSP+Adi4H89o4Pkq+QF5wLl/BJ6phnmH1YDSPMkd
Mr1So2rzOGP45FLyj00/veFLPstzfm+ofkVddmkoRGCBE650Jor9kO3hZ+/zpV71
Krb71te5MC+2/O262rIwSByTyoaytEAM8SH/MogVf5tp9kWg/Y7u1+4Xmz6BP44l
kA+Ryttn//VkxJXeioIz32mU3YCbD8Z4DYe3EMGjD/8lL5oUQullnViithlRtoe0
EpNOcZNstfEQ4wUCu6gQDq49naCVnFJQfO5o5sLEnWsxXysposGQkkb7cn98oKxL
OskZY356n3G9jkA5hAkjUfjUT6t+zVq3kHggXOcNkb6APUTc/RYRAqddfp2JnR50
fuXCFU0Wah+sD4zvTn+iiGzpNhIqMMu4+PHqNIrfrDZo8ta0MdQKBMEOCh9N+y2F
ZIcwvOE/XGYA3hUG8xhEPZSsZZE50Pi3oqrAapQflrJGN/p/3LONfXq5bfuOnU8s
74cDB/QLzRe75377q4ptq3C09SNo5PfDrTx+sNF3c+GDsIR/Sv1gXHAGdUyCHgcs
cAxh1w5GqgoMWyOrVXFBaMyzSD6yyCues56IB6M1qJN5Pu0bVXoBqbr2pkgEU3a5
RejDn791S0/qN9Uw1Yn0OwXpPrYUYMiMuVjMCjlR2NfBUd1gkwaw3P6eFi7dVBAd
WMrxBGvh1hUrKfd3F+vnxGefqqv+dt4ugSHQ5v2yusz4lTmnzTWTWj/CxD/EpZha
lQyQ6Rz5pOs2yh4FI0ZpPzkdj3UWh0ajCdFq5NDZyTGKTGh7xL5dSxvB9lU8/ObH
KxnTr8yoQQs/Bc3dNf8K68z57ICZDYyj7iB9+RALs6bflks1XOhmLt4MHYppiq+Q
3AHrVWNCPcjC8/MV0DeztVeVQmGiX9HJjUp95DOO5xOthEgvOWQzYfWDttc40bJv
7u2vlHWxfVqFxr9XM37YlqZ+Pk/bGwHeVX7zrzxprxZYAXKGzhHhOkdz45QkznFG
bdpz/lVp/zyQ+1QA+6ZHbXzaefFTnKi20Xy7qWlJfeV/5HbRHCF01Z3NCvyZ4q8o
7NX9wD+r5N12jZBfRyBtomBYrZ2URvIn7Fh9QjDN0gLZfsRZmuGN2OJzg0z8wjUF
lGwDvaKLr/khLts+xs+UVSbS/dHXMJtumsTbr0BE/5y9I5KnDEedk2RN1sQg+NSx
xyT5Zrs+r1kVloPKtbXMeYRKGyv85CFbgR2fPu10+CCLni+1TGPotXqz0fu1HL92
Cy/hq9+HWPZKGKpitHRf6lI/jXZKOg3/iGVVChwZ3+m9UIfUzi3Kc3kn6gfNV2Mq
KE8+ilUdnrp2+zN4G0ztULZ86VJQLtI3RSRg5pf00Ple4rcHSUFpZ+5sFae6SjWd
x/xJIOQwCOg7gj4Dj42mXYEujB6yxvCUxnDHF7Kq9Qipwl0Zq6tmy20Gr9IjXxNB
2IbLF5B8G9DBFhLS7TalftwS+2KlhwpZ7+5VQ03yzBa5rR3gfjF0ofZZ3NNVjiQl
bW1tcX1QQOlL8uCPDVSkxQI8FsQWoAsqxvm9PstyU/esyz3Y1aZ2eR5npXBaimJ+
dWuLuS1ADUv9pZH+EBX1069ivxRmjhfbHLGqEgf/P/JbWmO+g2vDFFDcMBlK0PEF
AI9LNlr0ge4GK90TyClOdAZc73w+4AuP8fSm4rpoNV53GhIYiWoC5z+u/a9S7png
xkz/grsLQLAS1Somd0OBuUCv0riPJgYYGvHRUxs8SLaoHpQG4ms2NaGb67X5agyc
8CUbzI4qgNTL4IVPKBj0ZPiqEqvAv6qRcrvPVQHc3LEEpdRg2oOp6EiE19aodNu3
9vqT3Zek7FB5MiOtz4dXgWMwRhj6Lun4NQoLNGO5XlAVoP/ylzwSimNHsifccObs
G+B6qjL1TLliEygGIGBMiOdapyIiXX3itGp7Ir8B7GwO0afzEs1dzvrMaDW5TMe5
b/TImrgxgbWqtbzo0oOwuZ+pkhPqfqltZB0fsf4ZBKSATn/asrAkUKMm2RB/vKzX
+5oMNo+JLUnlBGdd8mHUbVi+26V6OKZBklrwv5sl1GDSOPjhKY/NWdZMxhBD3HHJ
OT79cj1t/sjdogKgEWxjA8ePO2DMvv/EdjFH5+3lNPYu7sfR9yIQXpyV1B/IbRRY
zSvwSn/SFy6MQ13VEOdAVwyZvaH6+EZvTsN+XwYkpudu4jiASAOM2fhHOtTx0r9b
eQUUCMbDFBI0pg2znsrUvwCaDKk31QYMnakJ510oL4tLvkWdMQjVluKRWEP6cfZV
APPp6TPTwl/kT7z29OpxHRzRAvAVl9//qUGsZ0zdh7tm3+wbJ+wayDCtONcx9BJo
3Q/MiT8tNfrV4FLGrNSS20h6FfkyMHmyvmc4ffnvjpguAo4BtIcIHkJ0Qq4j+WHi
VfASPoGM8dBQ7pnjGLgz12++qtDrro0PQhhKwyIqkWOlBFxFujSsVoyOkmr56QVC
KRASuxl4Axcn5kW6pE1odoxdJEewiNxcb1MaYb1141qSLD3S+v5bjhJyVDO38xA2
scdLDu1zTmw1Kkw38GgK2l0snSFaw5OBZS4nP896FXAwd3gC46cpC5JS0IxE7ZhY
Ve9iSQDQfcoHsH3qNCHgdRmB8JxYsRxVAyPp2GT3nHGjgWVKEPIzXKRnzbXKKGBo
mmytINIuJXUoPp/NtzP0qGeKh1pHdixTlRZ1RPtugT4Ew18tYFtWdjtxQvBvon1u
AbfJHulNC3oXd/UQ+9wDvpSkSH8cffrzletb6Kl+0i+9sCN5ls24xQgRuJqiNL7n
gGU1XuG8wRoIXuRr922VOCHo73TDeZDANKOExE/OfVcp1dw8+Q/HYBJ8AeTAAE9u
rWa/70QIkRy5MKM1G56gV4fjh5pWiVLteBYyJlk/T950R8lGMOlMXnHBPQwrcETU
bYsd5adN1oCzoWZuSVoGSum35PZEg7SEEQIkBPLNl5too82zVqVE93v3LjjYnQZi
wiwDKY6kxMVTrwNK5MMOUCkUuwKg1xxACxu5bMmOOpgf//xDfDqXwGDVf4jYApDb
Ylq59BTUsy0F5LpLSQwlhyUILkoSN1/v6lH4Cd3cI4w0bOqgG0PxXLDOeeDuMZYe
2AloKa3VNFlibq/2RMvCZ36XpZ1U/IuiBKryEfWxlRHVUfg+jkOgoQ32dtKeJXNw
ZMydNQGTvLJC345sDshjT15HT4aTN03j0za3vlYsOIrVn6GeheBM4/Zn8JqFo6L9
qC/lRQ6MZEW4YR7fy6fBauq2mSCob5OhQoSBGL6HZ2ucYK/roXGFYe6cvdHcfNFa
59D7QZCtqB5kC5a3gtrtE2bq+PQi4qTwwosg+rv9CE4NzX8up/aPKCeSvNRqH8Bl
NZ9sLJXmZLfPxLE5zuZ3CHTvAouI93WnmTCR+kjh6MT7EfQnnhggD89diEuD1RNR
eZq6VOMqpQKyw2CyTpoE7foNfDzEZCB31s1I8vvOE283ZVle4uo8KGW2lK/c3z3u
VHLziGwxRLG3Sop+iRGlhGSYeSyo+1YpMvtyBzsugSAHY5uoqtLOPzsJDVxLOIuo
jDADMCksPQu1M8UAidEPn4xEjqUBT4TeD5Kho6I72QgLxNrvJZgZ/C31a2qT79P4
y2IZ3mzAtCMa+Cke5i22qLczNe/iJGNLUkJg9SK9NB1DhrcVgkJ13CC/uMoZ30L+
ob2CURQmmwrHEzsWChWLn0t92u8rruOttIDP1paZnkQGKg3ylxPCf9hLo5gnxJbr
F/KJO1212d23XQb/MB/YX06vCRLZWGXqEBSlPPjZqwCm3KwpcXk/QACeDNBCfYhs
SCxqWS+ZJWHnrcXU1JQqgq1APXupIchOB9euioFSkzt+xgsW0tufzbq99dLV+K2L
9x9riyVwnEN3U8HBgnukGRhTh5CZb8YMPsfPyXRL/sIrpmc6wN0b6xkHmBFsLR+U
DXXP/7AaBl3tWDSrSmqrIq5XE8myj6gQ1/M5n5OvaRWqEolzlsd8QdON9k7ZRQq2
FTHM6Pef2v1i1nHj/3yA2aSBSA4BBzjxQtBwjbw6KJu4/SXwuiPOf9z2ms5E62D8
qo4YTNtnCqhZmQxbnSW7dGRo7Wrb5LAga0HgB+Hv5UTLtUTfPwonVAnBgfLhffBQ
IxS7No0gxlgdG526RnhdtWPQ7MBi3apkqeADdv4CQgpwg4/cMrUEIMwsC+YQ95j4
RGjPwaRGDBJgGtnfK1ZLi/B+n3XpKwKw/Ioxd67Ewekg2AUp6odpp0c2BXFqJIjM
pWXxo8hTuGqaliTQ2YotwdT5ZX+CWd/liI/LmSX24xcnG1zPCKz6Is/CQLUrLU8W
rFP+mRbWuf3vVpAzuR17q+ax2jqV6W9u9GPs/QL4s5s+gIssl4O2reTYlss8xOsR
7tLDYwTq7xWbfU4MCszArsjc+YyXILbEHqQ0Zn1mvVfjE9Wqz0hXwyt9oKOCZXCa
+HzZGWsQi6ngkkznnmPybOAx90ZflzBsxqImTBUEwoIdLV9A3YWQoGPk/L/vs9qq
K9g44ihco4ThkD1dvbMxEuyr49U2+LSN6IaGLuf/+sqAdmTOii/9PB+yL9q4+jKQ
3sJlVB9XUdTpFLQr3OG6xF64pOATm74rVu/WCXqxLVr/uWpRG1SqZv+PIn/05bGq
mTApvh110P0exJz2EM/875ICjz3Xler57RoGAktbolmZ3eqqyZQoot+//tLnQPPC
Pa77XZaYBAesP6dW3V9/jrh5HIgJ2GWkSmci1FQzDn+4zWBy2AywZ4svQYl35nYn
F4jZRlVhed0O0bChG3gpihZ1kXZmF/GX666/h1AWKyrVwVdNAjqPeFLJEMWdgoAp
fNb1WD7LgSw3Cw0zKCvLDg18oB3kEI5Enz1m9UK5oI3j1kCdi8VXsGDIW/ehzfW7
11s/0LtdQwU8HVF4cQdJfRpKr+hdFXSpvaRmYecMtasXl8O6geI5k7xDLbIMtrmG
IPSny7lEKWBDGB1fbxfXP1Q3Whn6j5aSFygzHSGOUrh2+JRqsbRoBCPpiEbqsPET
99HeeuRGtGEFjOTxh+wFgv6fNqMxCeo9r4WbJsDpSa6wrAEouwn6g7WoUTZ92Mvv
7k7IMWdoI36RFv1OTMf3okf4xqEj03KCSZu8FbT6H9M4Sl+7hjTBsuzyUBrQ3FPj
ZOHCf0wVQU5Sq2h3fGNHiRwGxq9YEXFnobsvvyLdlaYvHIapkvw+dND0HC25g3BH
KIaa68ZDfdPzuRPqeaKfSZ/gIQH1HBPv06OlwsM1neiQz0Ng9E6CP/cFZWi60V9T
2eYiMYKLVjeE1cCSFYsqH3S3nqzM2g0Kjp2AYO7WWZiKN8E4ElZmx+UzMmv8sm6W
D4gGloB89rd+9yElXny/xQRCiYWNPjnHnZCcMTX+giD/LRc1XlTX6tqyInwr5ey2
jodUxMPXXM/ILkuKrblFjksyc8iWLlwSpFO+jKkybS4e3exJ/EuDXwTX2bodvCu9
MxQwIsUb5VmhxoQYYt5F18wsOArS7iNzSIPxrIBy9H/47hqM5JayyORD3Q+nNPxB
73+ODRur5UGkZbo/sLTepsszXc4PucQrRDNSIMHe9l7iQh4Y8eCX2SOfLRmyT7sl
3pfJTUFQPJvpCMSJLY/zObuIJzweH2mqtnv0j52lhb6asVMirJ86y6qrNt3SEL1U
guYF8euI/T14NtYEVMCIINmrBcKFd4OUbtc+UvSPsVQueSgY8ATV9ZhvR2dq9l8x
6kDL3H7BxAfirOXuJLtopjYO6aM1AMRkpmZLo/am55diAMNMAWVYSHkInVfkSs6A
OV15c6gqrN921a+j0I5+nkcHdcOtMBzhh9t7gDXQcvF6orIfPRJPH75gMPbhre0E
lt/AZxN52mGA1/1hvWBLjXZ0QSpeZyRy8Mz82yLjz0xxfbEUkD5es/wa0KovY66q
tUzuNls6vLVgfEIxiKxk34kAa7M4W5m15Vz4MZzt0xj/I5rX9EmoS5gE5NoYKgTJ
qlwnZ6qjJiOR/UBFsS0j7VpztrwViR7n5XwXqfeGnToXdkqXv2RitQ4wUcyRD8A8
a/WLV16jYxYBT/oaeDJV9yg/e0R717XqvdHSEHDUd39Emi2RvVS8s5pJzYdMKTMc
18rcVYBWtWgRWRDd1OkQwvknJY92qoF95XlXk7RDsvOjU5J2ZttLn9YZsXlHENgG
ml4IOL3Yz6S8lel7sLEU1RljH803aXHUSiagbPa1NNvmucCzjy5Ba+wjGb2l/xMv
PpMapEC55xnODAEx9jm0V3lSPerQFRzVBZ+RWq+E7XJT9haaF+vguLSMJo28YbFY
Jen3fjW4fGnG6Q2h49Xl2oKQQQsd18QukLbgfEU7nK9YhXkoBqGttEbf9oPyZPdZ
czNB8Du5yj7Z7UCOPobNXUFVzYbyUKPswZr7XKndgKr1HZyT0KZa13D7ThcvLTDB
emAFn97avH7F2IbSuWCBgJLGG0cnqWORmUgtSMS+vln5c9YZxjOpo7ED723hXMOg
qFQcAt4XSX8ZZTQfjJOXofsMHiTYQBUT9Qxj1GSSXkwpTd8GHFQmQPOITA16MOIu
SI068Bzf75I2ZSirCZpE4kSN9datP45C9zYpM9HFmh7jr2SYQGaWQHbEevwvVeal
5GvPuzxwSKpZ3AgrEqyRcCihwxr8zLpq5SoFjRYQz+oglhBGWcDIeO/AFbn4+1WW
OWXgNb2yGPa84ZT4kYing2dGE3CWFOf2Ai8xoEHTeJGQUFWeTT5memYV8cjpsgR4
alEhpoTH/Fm63anAXTUIesaCplQW0N+cTqyWreyuHEifBlKLtwErHg9z3DXOjYyM
R7hTdUnntbP02yKenWDMAiwDtgVhWj7+SV86A/sxHmCfg3rcvQO8xK/X8p08Nn+l
EHeOluei+MBbYMbpgwFzpScvIGHeAjOpSUMNSdKtUm9KFfZxmI8Bk/4P03fHHWUO
EoQI6ha4FUolfIrus/NGM7jjIl/Mw5Fg8bcSTRIH2R2BY6NDw607e/BT62gu3WI0
dZMdrkdVfKcv+n8uzNf+NSSBctWkwSuUE1VEF7OArat1zUJ1ojLVcj8pkfdsQW9T
tgtdxHDbVdmh+igILkxCykkoQ+H9NqY9pMu8iFthfBu9oKGpZJRTFPHbL0MiXTAV
mn+qrxajgHLrG5rsWEKBK/3NfMBgxcJZWdq+Rxb5MlhAflYQ2YUEUs7getm9Pj7f
i5sDWz9Z4eTx6LasCc3l8saj8L8IUHG8M/o0AK490Ogaa02k+itKe51JAy9nYkNm
XFpRAioNMlzdYQDw2VTmcIAMrGbGBeeSWyoj6tWvCBgBYA1KxSNuw2wFQXzZwhlC
hTdPfroxB6XUqQGyThtb+w2g65163MVND0MhGkDIwSY14Nu2BkwIbP/LbZ4kscnA
xWstE+64VCZOL+WkSxEObogScdP/nKs2jLrcOaddBz5w2KF4Jl2rKmBdwqlIm1Re
81HnGHgHpe1qzflxIO0wi40fUSSQTqpkTjuyQ3H/xjoyv4Dso80yfaRVIcHxlqXY
b0Cp+37CtEOic7qJFJA1Oe2MEfC6ojAxa2yBzCdSH1n9gT5Sr/ADBBE77T0MvCVM
T/t/4wk2f7/innySriB9waDWVIV29QltfwitbWOpGYwHVPOHLPhNgfwgNWpk8nx+
e+mXG8GZmDOUzT34zgsoxk0RSnTxuIXTHMzYsJLAcuk5N+oWsRtZOSIIXdcsx33S
9GKbiE57RR3xoLJQgU6fASt/vkSmMDbvupjXy4X2wXOt1rUNkBVk198g6n+8z9gY
+wBnV6wm3aBI1/yMxhZargYoVuZ24G1wLPfq5Fhm/mZUVzuVVa3VJX9jXFzqvYj7
EDy18eb7CixVvFd8fSGBb0GoC9ObWYqgQHbpGv5ZFZEgN8I8Q709nns6nOLNNbaW
I26U8z18ZiG2zmrFKvBdbRY3YKy0qUa8nHeWL2VpQ2VyyvdHjK66DRt4Qr5dsTqB
u63kWju1zAM3BjD5ylhcxM7TfGw32t3I7rDUwPENom0CDueU4Pu5gOMEj3fnkj2U
+9Zq7yEywkJzB4Cowt5UaQL/nuGRQKbdgPFU+qerGfm3mJPsl1dNdy+Powksefy4
BwoRKE0ya6OH53bDOmCJWzLqLefNENiOsTbCuiA4z2cLy1tNyHKI7UzcijcayFHh
IiVmfV+AJz11hwiugK0Z7WGEOcIk1eUpNYatjPjmyJV0L7K+G7DHBF0LW/l6HhDA
Xrq0oY5VNhax0fAwm1qvbNZct38QclmAnPf4dIvZTEHh8s6dcmTPC+qg1HTRc7Ae
17mbjjuhAh+O9sOKTIr3jyVcX65xz0Iaoasi7Tae9uggdqOJzmDGe+9vSoOsQ8bM
9ok9T0XxZWuPNxaFiQY1T8MaAeLenMdgzyXkqqxC/TiI5nBsRV2x8SGcb8T+E35W
3Z9TX5dZYxT6DBGeFOLibRQSvIaqFztdCM0PHSGmCQYaNafDQ5PVlYAIZMRZPbxZ
Oa0If1LGDFrrv4oQ2S9vClCrA5nZeiIhM46f3ZnUvONXBrkobHtDgltVYgXk7lhK
nV/cpLljRMBGHY/BeDqkpOu+Q3ZuMxhVIchea1G8cFcsdn6Ah2vGL2sBk9YA8Vw+
bWIPwt82qjQOxlGaljVa0XXmHhQELix+zX6/YoPiJ2Ucb6ChqNU8PzGi6K63ZktI
MUJPno/GUy/VW/B/0KUvTsl7LfuFMXGGZrSnLMlR4uHJ6KaZJhYQhT/Rd8tXOTfk
zsrgvVU+JdTk6Wven2oDDXewm6lqSS+OoQwawPki1Qwl3ykq0W4+y6CjfbLojtMF
NXuH01YZGQJ1EH9LOliD/3ROlBsxbhjAvAg8K+xJ7jCJMtNQPLGMcUwQMuNtrge/
z9mppxpCZigdDwkxrtoM8pH2xhCnmpv8IHNpRQDyKIag9YKkDSmMf5iyFvzQ1VF/
xnbiAdvZ922Z7JJ6sGvLGcX4Cu+32arWlBqMaz1jB/kKjqjJqK7RNHd5Nqx85Vnk
9FgtBP2MgiYCFOWuCaw4QsEpiTz6Vb6ds4t3WIRLob2NUeGsS/Nzdm2jz/tbRkSm
Ijsd/1e4Nn9pxmcIPvpi9rwK6+rUhUNmxEwlmfB4zolYFASprJSDOXCHle/DFoXu
oCriEHQo4ORvP5f/jOb+ZCWVybGWzrn7FC6KLPYbfTsI/Hu95EmPJDhyDW3mmnwA
r9wbe6HDm1+1w7RpdApDiLmRbNzgxI/4/TaxVb9vbZY1A9c0zhilLCIe+d8jKh5L
/qL4e7t/LZ2++zzu9hTLhjKqsN87M0ETqRORusW8KUA8oxgK973oz0YSnY1DAP8l
N6uzCXaWhEva75GLyB/Mb03HHpUGZaHtlb+M5KzNyC5bl6GysxoAHhb6VTQmF7s0
8GgmD89CQ7toJP2HTANWWeGz9xaGHoWkgr48TACMjcC3KxtrRMy1RzWfh2aV+xej
7EkxfKsc2b+RGqf0XUUOe6UY719MPJqxkeH5lZ2M4RTtFRFf4HdyOGJm+2m+JgOA
/Sw1zs54tjJgvimPv7DIAJHiCPstv1qUP+U9mHPeKS+TkwPluE2ZbqXu/IvjckH0
hkamuWnsW/Sk8u2aNtLO4QV2LyVYklIDOShAFYmyQtgw8RTx9+JyEEiJV/yrFeKT
aJUFV1VlT1hNt8VOsUxtgsxyuNKn9dFqv7JkMIcHGyKuK9Et19gmOo6T8t3T57BK
qEcrKe72BWPCDsWKYfz7ETdVKY5PzS8/JnNb+0ylP09s41E+gPUOWvFaqbnJAtec
YwdtJSUld2WtP5ru+Tnfrlxc2FhU2ZAkrZZ1Fp1Bu0pLHD7P9ccPXVTTcAITNCc6
FaO3nZKcWmRYwpJbj4USvuAM+TCenmaEOV7S8Jma1K6qnr5vU8oHIFhL4O7RdFnj
7ul6I9TqqGAeF1xz0c0F4Pv/hEdQ3VdUvpsrdyBeWUByxIzlieXg484xuMR6+4mL
Flx0H2FyvV/a/9ifMC+fdAkF3vBN98rt/qUNdKGUdSpgSA+knEjPvVcNcIYtOQZ/
N20hyvVSGkJZ5PKfu5MR9TviuO2epqVVefWhhnC6k4vaZw3tAPaO9P2aWxkhclHu
aLJVSzFZaPW0yXJ6/id0K2wfq6dB61XMeGRjKYu6CuCVakY4afEJ8e8d/UxUD9ua
Qmgqido0K2FIvTknTP6l+y6hlJJEfy27BcWi3F1SrCThryDM8Ur/aLHPQKy6xbMt
tb219OcJkyZhhKRKdPWBiaeZYwDSWdUxZ1zOCE+MCuM8mnucORIOq4OxdhyzytAs
6rnsA7648t5I2vMOxcZ35pMHtxVYBwbzsS+V6e06Bl+msqB6nUwCnkRNgC8JHJL7
gu0Mrnf+9Db8wrnV8F3m6J+OBKXC+E/ECLKOyjwVyS8cqoBMZYNXBtKZwtNW1eHC
A/n1EigSl5XSEmmqOT+Wl3dw4HwpisaLri7jPvrAKgyM5sZvQHbci7prxcv6UNCT
uzDu80JERigvEqTAioeuB1tvF6guDjFGu4yG7NGooJ2IZFqs9CbhZWDcW9ij5iSb
vKzTdOr/BpsugRrQwk+lULJREvBikci3XHgXtLWPWV7OxGiqtIQv3YQtY5E+vPex
JlcECLpTcse2JZu9KsS0lELd0iG5aM9WJrsnN2J/a2C24/3hWAX1eWIVwHxoczgP
C/yXPIQLvJexSutAS0hu45n/kpKBEabiQceaVFbKPs0n4OgUu2iMqCwOJiVKFv80
GKL4sLjHrDphR+Y4MqKd71Nlrh7E71KRbZkxZz0fw+9o2i6Z+x5pGZwrToY2vdjW
EYk0UYKYMyyvqdRT5Kg+433ruJURq+DollnQLnV/uhWOidb9yth4BYzGJpVhl6Se
CFkcSFdZ0D2lXT2ZlS7jFBdTFVKes+3r9dEpN69cy6hhTU3Ej9tbXVOSrTFQr/4R
1YVf4Sy9idxrjT09abFrRYRBUZey64z3kBbJNL1H2NqyMWEOqNKbYnUKkQvpQ9yM
yuTtALrcTroKwePRaXMUVsDn/P7S93NPLRMFKH6F27t7eSdkf5U8caNflbZmDckq
eU7tDYOQaBP6ulVbBGYZYnAtATr6zAvVbcAWXMOoirw9QKp7Nw4slvNtdpyA5rih
86jcmPhFqdgYw8CV/lhnTRYezmVdW/l2TvNXGiJH6qq6im0N461R0JYVQn0+0Ev4
ssoKPuI97zZnSKbe7HYjm9HB2s4ru6+Djh3hruAM5+eyCs3ZnvPKfeZLxLhgiOp/
7nLadQO1NfEBkRe4TBY450YINkpQUcX5zSca8bQi6aJYlOpKhRk1JlTu2NBdOCgc
7h1SexcT85JnJ83X3zH3MD6IhPLoBsSKoJLVqX0b2SSq/KIr2MF+BUmrjjND+KjK
kil4co1Yu6XNZKbfsyKzetYVEHsEy6JhZh8rpTLVLXEy8jBniRH4BhQumGKnnQAZ
1nOdeUSkbypAZAAMxUFU2Iodh53FtiyTY/o3p5MJ6lX9jVYhk8vkoxC75OyqfpHm
nQQ/5Px3UnSwR56wG3CMJKpZJn85773fi7H6nNBjbrogsOyS2IKva4MBHYwSqyIB
i+I1SZk2xWXZ5obbEabNNJn2EqvB1cbb0UaldciWH2LzXysUq64em7sRa74QrDPc
2joB5+yHtvzhFS8G6e2MMmn736raD7A42jDn/0lbxrdWQ/PzL1IeqVolBO9qIx8N
vqTNwztmJJohki95yoRx6XiilekjrMp49FGz5Hx6mkwujQQxDYChlru53GKzR+mc
SbxlRM6fHo3gfddkrgNq05JtHUc3HcFXYffuZSDOoRzoEjQMeoERJWPOhbTcoTuZ
9u4PtgYBcrDqPy0G4CIvbuBGWWGub69c2n8Tkw8FGEGLrtxcgMJUVB5lTDqxAN9G
b6fFFRhDfh7BAxnnNjn6sw5BxMrCFL+Ath9IxZ3oHHqRQWsvLyRH2wWeRSwl4dno
lk7ddYtjv+UC2yoMyyp6qozhlY8II/ZaUSAij68x2Gd9isne9Y/bLqSHtjBpCdEb
/kPbq/W9BCPPbSsqiC7T1H+6FXExqblOiDaVNEZdt1qwOJnaFdkLoLfaNkrSVRgD
0b8W4ybCaf2/ClL/7mvrQXAGfTDUDE3BncNB/0qKUJYVmSGaPK4NnjbeJzeebUBy
fvkO0N+SA0L6M5j1N65ELNP+DA0pGl0eHSmwJfihqtOeFavX2nwNcTvvjmhFh+8y
BL9gVuuzh8Ib7FYpmHlBtWdD8Ep3f4jihxMua1/mbBFsi1DZPU/Y+SPrSRPmg75a
lOSDsZ2ieULfpG5E0BE2jin3EvCaNIxXR2fOMGgtrF7eqq4dxwRkC+tuyaX6VRNj
sZ0Hg44JgASVMIKhNos3zGzWcrlpSJ7CTOAUwIpmijp2A/KmMQK+cdnuhqR/uYmj
ayL89fG7HhuaHCKaRJrtLv9LR+UnW2Jiil90QjlDGmOZigUtrovs7ZJcwa46c6kI
Rsd5P8iWZ0PW3uCZNjeQ8asd77BziB9AQpSUuzsRwBzzVDHIUyESrh8sNd3L2q0W
qbTmi18gZGZOqiGlQ6syII/dd6Omo3T+HEHEWTPX+/17BSKj+jHVvF+W1S/vMAU9
WTRLMubtG4FuZKkNi70Q72bEjqX6xi1u+C2vL6EaWWGrqEcoRbDenHdlM+3uWSS7
RLa/WZTHs31gZHHpLDCJVfD3Cr+ruHOMBY0aDlcRv6CSf3N8wGtFL3rsn18Nds5I
C1WIHsk5OyoEYi03xCsrfZAf0QRa3xh9v5QYf4IJIdHwyJP9rmjvHBOxqRiyBfyM
sA4tO7UaEoRbjbRMoZiuIh2vzmoloJL7X/jmnfvxcvl1aUgo9PP6+rZvSVR2kt7z
DQBXBuItHDXUDChWTKRXIZDhqyTFvBCBOMJU6XKya4u648RSOvZskODaXBSJKAua
HSN8/Ww/KeTjg45drH5ZFIbU+dsEpM/3mZY+l70zTy6OLDIW+4bttgRvBSinFB+p
nj+Tsfra4FYF4fBfdObZEPElrjPcHqc3YHgNT+VgGWaAcsYmozn9nobJWLa0ABpM
SlCYOEuTuTylRDt8yPEGP/hFhGuXigvkYJm7lczlNHX5/HC0QWZE/4q27G4y9313
T+RrN7Zpd4SkeMhcyXRHqFp5pOQBSEasCLOe8CdDnFVKamQt4TrI9RCu+f5jy9P1
2KE+OphAqMRYbt2F+9xusKPzIGlaQI2afOwvvQ0WXoX6vGnamQcNXQ7S0SQ3EasF
BjlA+wU1gLNdq2kMANkOgIDpkLuJy1bM1lUTpUJ01WOIlaeCN9Y6KX/FgehYZ0Af
lLSt0BLbKxgN2iVHo5r0+nOvSjocI3CN24WAbn28UjSmDW2w8NvBqgJ4+W/o9f4N
86/gXYL8U58ECpm2hdrSCb2cRn1f6GEZ2ZNrLIsrzOASXhVopU2wBFsyPeBJEz/1
AFsbaxNty1hIzJ8IdpsfYUxhY3WkWOVvLKjdSdcn113m6QCnTAwDI1RxWL9GaMId
w0uiKf69ur0Z5ISBnEQPkLq7XRU/DosStbIP+trPfxtb2VJ21uGFO7496JX1g6JC
NKhw6XQ/V3QpjuMB2VGAbK5FGu71vGjxXfrLRCu4B9myg6a0qBPvClcS1z8fZh2Z
4vaZgrq5QPCMX+RFk5BPhaplo1k4nyuLJWhd5SQq9uARDOFN4lIbTk9F5f3NdPzH
RNARpN2C8f7ShSof6GaqYS18v7vZAzfH1OPUBDbGAmYlGG/1op8MtQNx2ifz1bXx
HIDvhr0wPR1WLG97iHR5yHduSwvSGRZ3U8AogUJIJR80s+HU0olXvdUGSvkCdVjL
N17J1UNz+Zc9YEXdiWYOwenJjm3c27/QCrNItJrO6G0IJ6bh9xKMTgfxUBxbt2P5
npWh1JqkRkxGjRCL3fAhlYPRvq7XOeXvstabor1E9CZ/wFTQcX8CWP7BwHjs1LSX
HHgI7SabANLz9J4IxhFA9CRu8oW265OkEkGWmY2gRq8FC1mnzmE04EKQYu96+A07
zw82EqgVpMY9HcFLRdJAUCeJqZbxnHHo5ZLOPcCD2YptUIRx0KORtHxAuamAgfMn
EuJYJu+ZPmP3yCJPrG4h67X9cSkQEIr4hWbbEIy/jzzKkUqd6sPI7aTfZ+1Hd8BP
VB4GHqFmhuv73AfV0hoIq/EnXp5fRbVpInl19gSEGQKlVTn4qRsKAQAij17ZPB8o
CTPXRnNX3Yx7orQqz05+WlP3PO/4l1d0/Ad/rxM3N9XT8T+JlifxOdd+yN5WtAb3
DbJESK6fA7xMFGGCMXJCM1p3K/O2MvXDIYHlB8Ch0OQwSuu/1BMFtf7d7+wukwt0
2hE4Z4Q7STtaO7n4hnZRSDSVyWYD9wi+KekVnQkLw+zc5XbCnYdvyAAn8+K7NnrW
VTl0DPhu1EFihv54//191xlKWAen1R/BZ/Wr2wM1+vL6G/ensdmwBG/jl0guAuA6
DO/pOOfIh0fBEJP7/HllDLtyLsgkwPk/QjK3sFOVlDkN6hKwDCNZzeMTydHyyLfq
0+K+bIHDvjVIxP6yNd0/+Y2NRlOEToBm3UhP3+3L/scA5dQ5BmQRDSTDBFxK4sht
lvh2lzyL+oi1PLjTyllXxjPRz+uxq3I6frEJRNxBHowYyyitzoacPlFQQiP13j5L
Nvsbv2x9fKdzOOzrHnWvUMnMd5BL8LJeYDENZKBNJgWJ+OqFCwzpQXkBIKnFQWeW
GwtuQ9Xi5RvXj6AuC0rKojv4lrDNmcrHzkOdggH0787IQzxikenJOrj8b7ZSqYrn
X70fu2ouecz0nq4eAVx1xEpoxIGdKux/HMJIGPuF12a/lIWdGquVVRqpF/pHoHxW
SBKrjmkH5y+BxzYYdbSM5GOxhWwhS4TJdi3ouOgX5SP/pgsJGxP/3yNaG5bC7Q4m
SOurVBG8ZPJ4vAirxgFPuCE44T8998lQbrFEWu02vQlNLT96Ffn9P2n/6Zk2jdAk
O+yH8v3lRjuRAlAIc3AuMu0WFbtZtsyQ7Mis5rG8yrsKm4Rkv/yFozLx4FqtXKma
0v7KB8pg0S+U7vE3K2yTxlrque24dvhH4hRsNIrFN/D2ECXOA/XA+R3XOoZdldxg
H2kZzLTUmr6T+pUl2xn1I8C/tMCfq+ElYMC1943JnsOSghhgQJ0B42lR57Wc9Amp
OjTGfMJTT0gdfOkDMiSQRoqXJm8jaP1Gx8oD+Fxi8YA4eyT2Ojk0vGxKa1SK29gH
nzu4yI2k4sMYJJOpNCEpEi/U4nizrdNxX3iqZjFP+nK/4Ok5MPln7tM+72BHfySR
PUSMf2F7YnCGurMVRj4Ks6hlApueKyAhJkT/yqIvNe1pgVeKh4iPaMi6vKo2+TsL
sRe96mxC8/j8PbVFnTBM0BN28A9g25DGu4rT4RGVLkRwYp4BYwkWoq16sOE48JBY
wmStFVDJlwGw/3macBBK1CtC/ceHwmLschME1tFu1ox/357wp9qtdpAXXp2c2s9a
O835xDH3RkXVXk8Ypn70cpKbIGQRxjv6eu4tzDSRFyTlJt18ShsT9SxUwsEI4Oq1
9nmr088njYQkNT2F8f9k3uxgIugLKJAPgTh9LJvpdl5PUQhHpcK4F+dTNwKF0Foq
RyAW1YQLKJRCZQfWJvQ2zFGje2SN7FWZk7+qLEfyG+xghE7mixXMA367z2/usMG0
FW0mz4FGDifQPjv2hyT8A3bdES8J+xXOzJg4+C4mH4Jfonvi0xOBKO0gyqxQ+qQQ
0oiswZsegtCx/dMkAFTJdW7vlFDSwInqyHG52nqicXVmUnVPT2X/r3elGAf3xr8J
7AqCa9r2XvammmE7zmFbqBkQcVI73UuVnh3bi7ZsltGLUMclVxMsdjIAugoeZKMD
QzhJ3+fdpxuBj89AbbpaXLJBaKbIVEP5hxAYF2GqINsy5y84KYhhrvGDAYzwCSFY
MZf2oBMcCu9IEAlEBzw2gNrll5VzRaCai2rSoCu7pi2G6ukQrqmO7tkO0r9FJDQY
Busb47iAy0uVrNiEuNLnJHc+4hZJeqekVAsysAVRr9l4TGNyjff7EFptK23cr9sl
8xOk65I5A0FQqpS3mymz3d+XW5cAqMDLkmX0g9K1iuQghT4LP/1kvQcy17sM/U42
8equUbqz5dnd1AxNLWjMUjNVWhj4mmd02cs6VGxxbXhgbvDNSV3g3hQ8WykqNXmW
palC0TYLksBIlrqy7mRVpgNBvlFKXp55hF3udaCZtYqXe7c1BtG0KnIFNmP0E9Ao
g6340/c8GzAI+5PblVm0rTRJOA+wf+d5vZinlpZwIS/Lcp8kh8f7TfyVqIv7JUW3
rv9dyDctr44XppO9wMtycKM3CZnKwEi3zFA5mzo9vw282UvfUOjTQO/Bp8feLX4C
osK8uo2KomVQGt261Y9QhKrTcxBFg+BVG2LCg+fee00XD2oTz9XpabYtIy7vSJBl
bpyAEwrzVxCKQx3jb99M0CbcoPGaylMUMcFTayDyZgrHy+OzWQF8ZTXdeMdwYx89
Sts/G2or3o5lrvAQoFnswy7RZdr1bJv67mnds8LGS6YpMGv0ubN2OXMEBqcAzn2b
7mDiLFMLpHbSdmlPHKxPydURHlDE4tfsSXpuoi3xH3z9Wm7/5VjpgalNZnl/gLJ2
2dXyDHSu4NNaHd/xHZEIzRX3yFKnQE2rVRmDrID/fCgqJR1HjgpW0ktnEEGSjPnw
pm5lhzuTe5g+pwluqhftguz7BIu6hBNp+u4LtTfFfolQcBBMNwnYcCUd+myJYkza
R24WcFa7uX97YX1iUMpunDIttNkTCDApiUoUI/SB3XXNvmZVvcFzM+sXsaM7QkwM
QvqfH7VPtRWSY+aEyPuGCharF2jhbolLeF5zxiJuhVrmNiC1TFD6EE7RSpFlI/rG
L3XK0kB6vRmUXpETki1lz3U8hemlPTghi87gzRHXcz4ctk/kCgHB2FUu30I5Wek2
jY93qDtQdKpXfjS4swLfTCBoNYkH8tdnCjW+Gh1IYtt1xhDu59M2JvwZy0uV/bx1
wwHbCFAuNz37E3JU9xX+J2EnpC4F4hLFTy55VyN5w0gW3gIvhULBjktGP9cFeStQ
m7c36Ex3+Ffhra48GfKLfUKC3YOV07R+c8gJF19AmWaeIZ+A0SEaitA/K4wmb2Hk
UXdFsZ+Q8vNRS2M0fs2zG1DohNETupXQTqdxQ5+r0Q20vcFkgulfHpOBGnw/Rd4C
Z8QI/7AhjEddEhO+SCwstQVUZNO8JOHSqhclNQhpMaqAFyiFqHoaQt+SeN0JVtWj
JI71l80TcVyCZAlrRAoa7LV6vEYOTQmtPcynnkXhYeC9E3ncI6H94YhLb2X8vlLR
tN4LiBC4coud41OAmq9gjsGMHfshqJrKU04W0gretVEvGwB1a0/gCdRqr2p+O7Am
Rfe6Fp6Q8sEz6F+KtAfjxANMcDZM+sqK7ewHztiTMUcIBG3HK26HM9Ie0cJmTYWF
WSRHa5hbmXCLhaNOfSXDawGqt5q4YljEBM3+0R5DWR4qJqo0c8Mn6IcTn0hDjieM
6LJHHBs9Mr6apMqTPOW2yKp83Mw/gCHBa/+ZwQ1CjN+sJxPZcX0AlKhqILoU7tmH
NUZfwaH1PL8iyCZaCa5+lmOPH9Qx2zTHONpu8GF9P0vtj+UI0sKnXoriScrCdPAG
H1qNl06vKoyBlVcymX1+sxied0pHLkq8kcmb7ixBUAJdU0Brhr8pZFTbYIGigxD4
bqXwMpwYz7FHhNdd/l9YI7UBB9+9eVuVQGWXVmxCvKExSgoww7qA+sOjhGTLGT3h
TfPN/L41iJLcEjvdxa83g8uvJe90UdOu6UuNhKmtlIODn0POXSW3C7fA7ENNqia3
wW4UhhxVzGFWlrZEl6qRdWY/fU5Aho4nAmIjpICfUeazCjrov594NICqayfQeUgp
d3pAYvUYL7q8APt2k1rgIF6ujtpaE4Z6tscBckq0SIf+JyfiXdMk5cWlOSaIQf85
DGXeCKuj/RQ8SGpQL7IeAmNIt0rpnEMTx4U4kr88eBz2d5vw1lg++dY1lgsBQr7O
toohgJ08Yu7WtbkPb5r5JN9OCT1y8I2AgUMDJdJWAPkI0ogLZLpP5jNCZeb+g0qm
jdy+KsZV/+r7BWBFCzMpZdXDqcBLICxwchHjyyvtPVB2EtUJ3qW2eFUil1mPpVfW
3v+8yoBQB9Hjfru+7F8qToJ5GscXY82Yx6ZUpba2AVD5nn/HlwJ9DzDJUgJQcv9M
w2ks4iKUW7SmCyZwb50cNBixu5XI/lTDmk/rP2oehyI5ECFOGti0XyR3q6swFJpD
l+fSMl+G2yign0WaQwITI6A+90bnehubLrVeasixTMymmnfUJuvUbFd0aCZR9HG3
KkMtFsr9kAt+B8ebGzYQXQJ4fBlM/WEW5Ey+ChqNJbIk0kZhqalczMsdzRavGRA7
fm8BEumPotjCkS1Z/vps5E3FVcR39rLJL+p4UyDyTpyoxidfoww6vfnVXnRbHjXU
QmXT2QxpZpRXWODKudmOSuG9fP0PwDV9CNoVWzfnvWhPJhr1beYmaphQEASUr2df
DZRSQygLzrfchC+BdDRDRReZnCMNoPpmCbdaqcQqynsWmg5m/87kCZ7qGhLceDqj
0KLp3NcXOGkR8A0lE731dj7zPQsSWK6To80RyUZJqUCG1r3mY1HfZ/+xGfQZHo1R
0bUbdKYBUoeGK9tL7NR28d/nrDHk9ccWrArmDV8C1vcXEPqiev9uj2IMcPEswJJI
Mwus+ZbuCuh4NXpzNCpMvI4r7JKOYxZTw22gwMjRDBKlOwBNm9mjwmU0tsVYtUFB
DbWCWfVwZ+pW/azDlihSmzTWLslN4jLxZv2elxNINBMRFA4QTRdn1VU4/kK5J31q
ot87UvLYws5TnirHWXvJvTXJFMx3eLt1O646CaR/7RMI8sH34bQMMIwH3LkvHjc4
ha8Regj6Is7bpwoop9WcIsBK0Xovk56nwiBpTyftyjX1IyOQieijAz0gyChlRbuQ
xoBsP9Q91S8ntomLlfqQeMdki/Jrx7pIcwbpgYR24YGNzhoHnsYzOFtBg5G14R2t
TGNuiVMGhfliNQlU2dczSV1pqI6YwovpQfxMh7ozh5MWV8gJxtjsW4REnOmex/am
aZOin+uEAFdz1EJHQx1FJBDE2uvUi9ShgBApbSk5V1buNgq+PNwJToaCjRbVjc6M
H0MPMBdgyzoGTsKHN4e5Osk7dRMAS6GhaOErtJ+ldO4OGJfHHnys6RLdaFyW2fEI
10LOnEU5i40/uRIs8vSYtYTRc0/N58iqbDHmfhb0h1f9yGyDwxSgl+dcZUGbdSId
M0TjQAQrNPALUTNY9QcukvvSV3wk/yrOFZXXjSBQpcNgGNJk05u5JZYTsjnblSRB
sYl2CyMu3cYIAaPhODV0SibqPm8behwDTXNYnl3kfUL4sgP2Hfh6Qkq8iu4Qg1sq
TONEPctJLujNf+dTzCwep5YbVY+s50B79qRd4BmR4h1SMlYu6WF2laa3xrF7OqPL
Abig54zKIZ5Ji2XCpwCm8E+FTy03Ar97XU9tnCiP47JHfnd//gOnWe60z2sXQw/Z
gPSbmoRR+VQHet94m1Quz2xTF9yhrzRlrC+loi8rFd8mkif/ItLxtAITje/jHyY2
OVuj1SK4/VAHvW+VV13IM39qJ29qhVeSjboc9atOKu2hF+0aI8MUTx14yBADsX3Q
6Ucy065bIumfIdKUGiT2x9v2dxiiGZytCHjeLxI50cX4wQINmGTsTMSmWRzdVqDY
hWCTstd+N//QZ3OL1b9tuzxLUiDMR8gcFvvhpt6+rE6yMwvosGB5YtSahkBSXlGh
0PJ/u4vmbBdvDp7eVY8ZwVJV+kUnprfLR8Uy7iABtLHZPBp1QAL6pVR50oWAbkXo
gX0taLPDEsRT/P1jLHlInE8gfkPlsnfqj8vzBnct8UdPAbdo5SSflB4Hjp5aBQ9t
GDLL0KSuMAc9l3P4KzBADErnqbItYhGHAvv5vUrIOjh3qWJDwqee+0ihlfKwU426
EA5dl/w2fHhkDr9J0MCkY6ZJ/N8GUpcA+B/reZiUcK4QbC1lOiE2GdLasSb9dxOh
uSdLI12h/lBqLC/nsB6YD7ro31cWEOn/NaV/DsCsy1iNBfVWcg3KWYipkSxDPkEx
y0+733xuLs8dE4MRRzPtoOoUqOPg0CeGFUWKE+aQNnjPNMwu0k27KeBKI4ZxnUMM
1Qo7IGDNwl6q7qOlJzy9nr/6HcFprrGRVmfC0HaICm3EtDVgjFP0vwXP4HwQke8i
895aZdjcyeMjB73H28XLxY1uU5PirOlBQnO7ZxsLKyYbBl/qFLlc+NrCc40t86w9
NwWyf+siRXByihwyD8hcNiRBJqdKG1JmSK2IgnjZRY2dVnHwHbjXB7Wdg8b97/Uh
6E2fYeP0gtd6YZnu5MHpgUe6tjcEeAoRLE7NHav/RIZVF5IJwSjYHBOzapGuEPW6
yfev+LI3MqZWo4IFCOtSnObYQ39Z609qnGyEL/obyCMB2hAXkR9mLCWGXiLW/A+A
QcCTziN0zcpa+hyEtSxXtF0c+tsNX4P8iR1rFialDihvixFJFVpG2iZ75QGgn4jd
j9QP6Qq0PvqMGmV0kXwufI+TMylK0kVJTdSK94YhbZ+JLWfphFEbLa9WjOaacvM7
0U5ROUgz+fwTx04KhZDeLEQYgXnWt67FqgcRRghwrBgSfeQ3xeWNPQ+Fd2PvrUmU
aWDW4ZJWWcL9mzP4KPxYRyFMeHtAMBKJmrIrJ4sgkzyGgrHe9vUy7tgmDuZUd66A
eavsMP3kEnppwNCEi1F5Xmh4lgtI6kPBRW0d/R2AwqMskvvyZJMREmNGmHoIKqAO
hk4mFzA+u5VzenZyq/SWtr2j5L8oj0imIbbUKIKAX930tySZvdbpClUWImCnvBHF
mMG5KlxN9bThJ93bsRrTO3UJhrooXWQypnHVIz6OpTQDUf56/Nvyr3/WOXRM96eA
7oQ0DRR45dejJ7nu1nMmKm0LUh2f3dCkCr/IJ/4nzLFdQi5/NuajD3+UshC8anzo
47xH/XUI/XhCsdBesfEWQX9QnG1S5ac8eE+3sqh6+OgL5uA+P4qccT34fP/Z6O4W
nT31dev0PVI9mtfPPmuBgaPKZFLv17f56ske4l2PyxE0IwCB5IBlDXLuzJBNiu40
470PjFciaO/cU8iSYPRO6c0loZelPEfmht8rDO7c5gPxzwhr7NufiCFvcq6qLh/2
KEIJCECupvZsgM4b0TquBoULjd+axPM+oioFNWgigmEHYvpYQKQoyU0jEpuFpkYe
eRUpcrg4MlhxVGyJCJZZZHx74jYbF7tOBWB1Poi0YWI5vnUbQA3hnuslY8Fo9XuL
tOqZidyKynIwupJG5wM3uHYZqIKUcfEEqSumj+t5LOUC88LubjG4qV3VCj/9jAc9
1zS+xjrmoOCUr7apR2/A5W8aUWvv3hu71K7fdkAfxVUHnI8ZywRtCUYWzd5v5NV6
6kSLQgR11Leb0RftQm/LSVvIJas4OfBAMGBK/m52l0yvVPxHIOjK2NJG48Km378D
cNmjhz1E1ZV+YtDqBHB3yApL6x99phmYUU6a9vSS6zRLxElNMW4hgi2A8fpa0/dO
hdnJw0pSFZ0abiT39iJAI5CX+z9mpKFzm935ef+TGsIfwwsPxL7W099fm/HHqIqS
Ph4Ym4xaOOEacQS0Tbn21pNfCBaZguBKJGcNDKYSWoScggextuoPm19kLy3oeaxc
SMiEwublcVivhYRhzt+O3nRnr9ccjHaEfYlLlSsD8VUSEheu+ld32n1nu4ywDu+j
haNbzVXvSUbUrmg50OLH4KaeEZPOBuw7OhcMCAICgqkNsYyQqVWV3wsccYOl9Drn
7h85CHdvq51BNJSpnT+uv1KEF9W93/7XUN49F+zlXdDEXwK0ieA0pCygEmZKwEAy
p3DULkZfflkLE5xMg2G2ijtayRaMfKNwqSMMrrQCPuwKVGhEA2NFB/xpWKF6PxwA
oV2AEl1OcS5ldD/F5DCm3MeNHYK63ruHtY4MvCw1UYuqZMkQWilwuThSfhiK6/k+
5V2JAGWzQMfKnwQNxIPLA7AazNBj4xx6q8P3qnCq+qoWazGV3IcBXQm98Sa5Dips
TfiBEDmP3Y2D5YD1Oz1rIxoOHKNc7bbpKkAJiKaMQhBGnbbeLshAFr/Jsk+BulwX
iCKGj6IKUjW25Wy6fYdagF4+7fkR6wD83IHLxr78qtE7t8ZPrGRE5OMeUEkBPlhp
0kydWDOcjeitpPDgzOE50mtEkdWhWtrZ6EQTeujKDIRYu1mci/o3PWvE2kKH7WYy
B18ebReI0C4pj6SLKPohgFZgZeCVqW9nsMFc/VZNhvvJGlYXEoAW02rdFSDEhEJl
CaVxOJeCOlqex3xjGF3vyy0iixvgU1SnNoRKzt8pJr5B3btZUp+gWwh0loVnTChM
HzSak34Flj0zK58mFDzRop49Su+zEORRSP3vyM35cPNJV54Bgiwjcap60xdeGY8g
zeo2QUXhE9vzsM1/1QapmCxnVXMwIN35nsK+dbuvINq1rM46RiA29PZh3cVeCrVC
ycJdp4WamLZuEwAAlMc8GSbnGtk6QxfFGbxuZuSsHn1XSmC9sudvtT+erltoNq3T
ddZvHTX1JM4H+GAtxonktXcQPTwaseNse3qLl4ShvMd1z2EnWluPkpHuncvkMxSc
9IPuqzgj5n/lNIwMSqgeiAGAZdsAwcHMaa8C5+n98QwHeqszIcBALvUlPKOzdxd8
Hg0Emebc+FOHVPKuoh13jN/jalVncpOVyZg1p4ISh3Z12HLNgWMDlDWz8LPoDfZ3
xwqJdEDFWisDNh2KsVFqYdnIuEw1NQ6QI8EG9s0qypKK+Zmmkkn+YQlzCPpUWBcD
iq5jI0HgwQsAKNwxWPhM/qF07XfgC48A4P8OoMNFKDCHF7e6RuTBYEty41h3CtNA
fyCiib8KPkoCA/TU3N/7GOgUJ4uMNwlvXmOOwnKHWRN7DjB4wwk0R9zvQPP2CImQ
HO4lestyoBxKszp8DBriOxJoLxEgVICvz6b6259u1O/DurH0U12lHhKiJN4vyRUl
5DHPtbiv4J5zAzV1zJkyEZyvHVAuqF8F+/nZyGQh8LJ1kbIjz+hnV312QInyEpDI
ugK0JIiDoUV9w5GanWPE9vgmjgFoNmLgRKQke82gmil0eQ0Fgd3K/j5MBivrBuGU
A5U/7lr47sYcFqlH0sMzNI0dftUhQYYj5TLVQzEFWMwJLaBe1qrMVfmnCQhxcnvZ
z9xoa2O1qi1TVfw9Qa7Pi1zWKh8YvkF19k4kgeZU5i3d4k+icbwb3Ah4oMpJiCs9
fdj6j7WFzmuxD9sBwO3Oj3KZfiKdjKllNS6JDx2/YuJK+AeVFZC4n6Uhjg9AuFNQ
yvx0nYl4ywRSrlYD9lrnBCC0NxtrAyaCeUlyHm1K5ftXEpXaj0a4iaLA8610qG3W
8es5X3A+qeEeInsMEo76LiriAO8GnJ+El3YMS45tAbQJkZU4/V8Cfcto1M6t5AtZ
r7PuLsG7nC3oy9a1+ZuOmvqDMsHYxYMYCkWg2BdOXLnTD1CjB01+5llBiF/7FY69
XMWdJ/U7rR4CC6hXZuerHWVvQksr2RLDsF9xr0Q6UctWXNl1N/7Jbwto12NHMO98
HgkSx2sdhDma6KNhHdSpNufF+I+8HKZWU7Ngb/7Cz1BV3533KZ+V1aAnNsyiszzs
ifDLJxBgRYrLN4DJUiPcTb0cfyaOKv8NFLeAmkok82hzIA70Wd4CqDMAf3xp6Y+K
zdIheXUUZCfG9ukFa7S3SJJ6lmpPA0Uk3k1G8s2QzPTFLXUh8KmgY6zZ+CMRNJAB
xu9zS61vGVFrOUglLZb6gHb47wScSlI9pPAoxocAv7n/DbmApbpzCKDrmixCGhnD
P0TQ8WqKXzFTtIKs0/ZOaJ5A8ZBVPRXZpInjLsuugVPwzlPMzOHnyflGt/mvP5OM
w1n2UdG92dVI/9t4XLumyCxoqmV4Gzt+OYiVrhr8f/0p6ZeYhRTq7S3ABQ/i/AL6
GZgFvyGFxdyUbbuT4Kri2NTTrky5XTqQQSN80e9nT6Bj+pfCkN7GLCOR7XYpe+3l
ya1c0l+IQUpuHHWvRUz26bbBqHEUsJbJiu5wvgfhkrFPq0c1EhI2iFMxNB0ZPCkF
SJ83aFWoy+6W3uGV+Ro3QQWg7scdG+Q5KMY+HuPb0lTNAySys9sMjpq0me/MYU9m
56aR766XdDjPy6k4pjW4+FoiS9JcJ7cxDjjX4vHHnQWpHcdZXC/hhgHSuA9awAlO
r8moF3OIkCM5WZDPO8I7Vz2K1Y5g93+B074Zd+/qCZifqkCZNuZTI79zf1R8N4Oa
IRMmwZaM/4dZt1rBGDlT5dwiRksctLplcTkwlVGQCNr8tiOvA1wRYl4JJ9TopCOf
Q41yTujdbrkXPNTxqS6yo12uNthTjGXwP01oV8/LRzAShpPgGLzF6wOxtaaf/XoH
rmL9ElVrTJa2APmUJc5VnLdMDxtNWh6yTCqYhg8O/bnMRtsSLSWn34A1/2H1REBs
jF4otyMOfuJdZjRSdlDoPXw4WhOatwkffOqlRLippmuQ6tH7XtNs/xmBKwJpFNo2
y3kQ8jvO7PFjfnHuNSOXi2JVYtaMamUt7beVhXxMobO6orF70Cu8Krabc/gpGLOf
Kyz3tpRKZUNT/UdDKtmqYzIjN+aOfBvW788af12/bpSQeYDqSDBI8z6F7trYscS6
KHIiUPUJgQXCZEkhYvnUzcWl1cLnqy3t+0BbzpUBMwU82y8FA/DqV6aB1XmnW/ve
OG99mKE0gYzPxLbhc6687iGKiHZrrKgCPTrAPcf3zz04yxt/Yujpn4nxpGhQZGoh
z/Fy1DC9tzvkrq/Wib32bkBsW2PtIK33SzIsKz0V+zZPr0ZbuEDG4l8wyUTN/9hv
P0Zt05TZeJht2Gg+gGebQtuwDFMg8I75b97DtW64EKBUsBWhd7/w1fWQxxvO6unT
k6npHlsrz/0G56/byZe5XJzeraxNa/0UQOUCm/KisbzzQ5aJruAAoRYaQR+2dCvr
cbb8z0arzgN3rxCaBn0jAuPPRRmGg/WMR17N4SLrL9TRSvzoLo1/6XOVUt2BAxWf
9g5i+22WwDmjDdm+rYp3BlXfQoXvhuseehTyoKyaDIImnWLqiS57CQDtnamLoX1J
GLM/4rm08GFokQTtlI6uWMlA+db9rSiwflSz60yEW+acG6eCxv9Y0OzeVCTNhgUv
nNsGtyTM2s1kjLTcG1x1HXTOheqYVGy2U4oaF8uaa5Y4c09/xIaN6jpIHphAipqu
JEq7aCZvtfwqur0TvmuMqD3nqTwJ73huPkY3RsWR2SXlygpAstTEBnbJsAgAuJce
qjeoNNVQ2EGOjSgao715/M3LLxO+EiTzGtnHak5k9Tgiqi6wj1yHtEI9IgrpDRQv
tdgISki6dfba3DmX7fJ/wg==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NuVRoNVHSdZUJJRGjC4J3UI2IedkVVvPV1HAPwoZi7u+g8JsYCp7DLCYqXpcnb31
F1KIaviWaPiyfZKJJD5ZRSEX0NEDlEWsW4a1Jm+RU0haIVADyqcmq8VpXqLn+CuA
FEw9EeD/akVFmEaVvs55H4oLXBnzVj2N7LqTxtiiiq878CSFJ0U8ZkQrqRHMfDUg
e6XJsaprWdeNDA9kOGNFjUrb6XV4CVRWvL0kEE6oqja+tEXxU6Ovm+7GPNjq8oID
PwaTk3d4K3ggTUY5DgyzsleTv8ND5nK/PbrNLprSvwzTCOlB6KCiXcuSpZhxEHQs
O5ugzCEIJUVsLpRB4WcoBA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15856 )
`pragma protect data_block
AbTjSgYuSVLKNiWwiObbyYC6MlJMtzGcjILQjZ138G+NCdXPh2CvuQxmctIuEBvJ
LaOHp1+sl6yfIJKC+Eu4CKFqIPHrN35udpY+QdzcVvS9WZgJFfUiCdOQU1JO0P37
8QDshqCNSVX6J6aoOjvlpMJjqfx8erHJu9yoz1xUJ60Ul1608nPYiNdxR1XYA03P
gAEjGiHCITFLqttPA0yauCkjVrSiROvWgK7hzjatlVZghsYBzfNXLaHtJ9lw0vnP
yxkHVSFhtoH724jxN4CBqrJXkf3iN8qd4x77iLbyTJUiskGw30L893kQ/uG9MzKU
r1qlugEd6W/Cp83wMYgRJM463Hs//zhp7s443fy6AGRS6j2s+LSc7tMapOkJyHli
qdWFTAQ78QPidliSzG2EIxjb4u2f9v5qm3Ny6D19VHSIOCtNb0/JWSHsJwLnbe+s
JMqB5hLiJUSrCwQWxJTw7bqPpqINIZKbuvYQR4uVwGXvhEwOtJoVIy3v02xNVPoR
Pb7vEdGzc+jUGBEaxVgNBnR+pIScQqHpKCwOSAxPO3Vk8QYZZZWKapf+g+t5w+v2
aY2GfyId0Wx1Wz5DPNp0JIrTAOJpjnUmBsuyB9UOIbgG8+HhGraEIeNTLTpIstOw
/J7yT2NfxFlIqsC8pMpN1OtlO1166k+3BpIntZ+r5IZvbyNgrXNdq/pK5c1JjbA4
ngEHfuuuKx6PURi+XMzhez346euGYYT4Wq6bky3h1V9VMIrvamhNkLQRDbqMgzq0
zopU4AqPkkFg//nr+ZN/s+r9rToQPgnx7vf7Jhf4fo6+U/AiDiWrN2W97eTsyz6H
+xIr/u0w+6FPnt3Q/nKVEr5FL2+dVr/gBZYPRj4hhb5Mx0uOwbeGr9/4/KbuTY3d
0H99phqxh5B3ycNnUTdkVFs21OGGUmEeUmWh8Ny9HgVQsxoHFof9KEsT8eykGkRW
u9RmZP3Uq/pjmhA7sQ5CdiOVkpgnSm6hMJLTWsHC7ky1THJ9AC1dD1H+RexRTfPu
k3RWeuGewcy2EizGfG8ZdPTXFNQbbf3rUoDb4C5fb8+0vNFINufH15d6lsroF0Ie
9+vYU1pct5fdxz80UuozMOwwXUhB3VPA108TRgWV7V4OG3DHbaBaCZk7hAyeH+lR
7J/soEeMAezm7D54hMLrsBHNDRo0PmELkZUSCWC/v+RZfiR9dz3kZ0W57W5bq1+Q
ZX4l99buNSeS0bVZYTi6+Vok7m6LSmIaUpuhVf1iL9RN9seBo0MoE78x29v16wHC
FmBECPc1XiSGkoQg40fCvWoweobpZKqpKFTcUrA1o6LPiURJU9y5wAv+unUfoiZc
+uVcd337PEMmCmyIpr2XhN/cg9Z42TJkfOPTiD5as/gF8h0eP498UogYeGmTLxnr
CrphA7yrEgzXGBacaScR/g+df3J3ZDGOYkxDmt8XzXF29VWC/FOqyU3+aRq7A7Oc
+a2f9fMGzZIQaobBwVCo32SyMb6wu7t6vN+xNhBuKvDQoy/TFwhEh/gVVv4YXg3/
D9a04Zp3yaWpK21XkZrxtl0R05UY7Au1lASBHq0TKcJiHeo9wajpaHkoh/7fyDv1
+BsDwVPbrpAA+73l1XNryRqa4uh1pYZH3ZwuLwpXxw0NOU39h+dWjVNqgEBvylKM
FWo0sntOQKemJ62oLvijuuXvPU3oECSNV7PCbkYfKMU0BVPE4/rGs+uqAxERFEZC
9AxWbtlmhpaubi1b1VWVse47pzFcXvrNXFSik4XZMfT363HJIKY7mn6VUue513IM
C0i1Xh2pHtL7aoojOaeGN31DAi3MAFdsbvOkH0o+G0+qzmoRkBMiEuMF60/Gl5ws
UYB/Bl0JAHKULrwqlCl7j1T5UaUbY0ju8tw8sQJKOCnfRaqzawfqlGhT/WeNMhng
kOU2irzYWk0YMdv8Cf0rxl44MHV9NzgJ34/XeV9YFEyAVD1P69WRw0++F5rhjJ7m
JlbBCHBNEXrBZKmt6tN3lbuNRQAuBCwzePSKd4EDfs/xrmpsK8XuSnWJweOlKACO
9qK85thu8esOg7QjfVj6BKt/NzS5q3AdSv4aoF+kPM/rgYyvx6a8KYn0qfGYgD+X
otaURAQPvbWM+BCIJNSprS9f+abkLAF7GKZcQaK4Hs4ZuDeb9Fl1KBFHlR2HvjOb
tb9kxdEERhQwijIh64GTyRT7GQuBaxzP8fhD9Qi1G6Wyq5r1zTkWIDjgZPJVnIAq
CTpHeZFNNgXdCOCwzVsUgnm8ESonF5UyE02+Sll3wVF50ucoRxVziGwo0Y4qkrtP
VIH3IWiqgRMuspJtYHi+g34NipgHGxj3x1wf0vgy2s7ctHIPE6LbnUdOJf4EjUYu
mqivbSiWlvrv6QpLso9+x4m3GzYPiJ82b3+IhV/rlhL1n9zDOeFTwoV2aYZdtwMo
MyQ7zkGM9G+3c+FJnpT567Yi5Ftu8p16o6ylq7K1c2rJZZlahkdnAnH+VALcaP3h
6l4gMDWVQmtfBDcps/ORlpvBDdAKs2iu7p7FcnjoKMCZwf3T6ZY9xyfWWZogXv0o
fO8ndJ032Pegqi7fM0f1vskNepG1OScNWUlkh4nP5t8jnS8bwMbGzwILJ5qJzjL0
2mgWX5A1rF0wpvPKIWXQ7si/VZxUt88nDNa9aUrO/u3P96lA/LJV46h9iLyKQhRg
tep3fmvOEQJQ/zoA+aaJb+ek5qB9pqf+SKQzYK/U/MNwEOrVrLwDft7V8NBuCbbD
7i44Y9l3PkYWIGl/ZT9+8UvgQtDe2FDoowDXyPyahw0V6fFwVWEPRAbgwvDcMkw7
XsmFtG2Cnkh9RVYu6b0LkeJpA0YecQpaJK5nLjfJkNle1D2L2mXYizFCVdakM/UE
5zisBB+AkNPQ7GJz6njth3bwbFhjbFYVDKq/IsUMWqCRqDNeHvpRAQ236ALfsCxb
cr1E69E6dI302tODn03BE7qXDUtePGSeHh1HpUCoLgDkELDN0mnVzoVHSS3z5KhU
lij01GV0DRoQVQW+xxnFMsH/fPCYHYAAJFn6rEs/MIXFE54QGMJVkVslAtPS2GoN
dcFv7HvotduTGrlBPnJ6p+bFNO6aoATp/CJlhry3RHnbXM3CnaNQRCI7vTR3jsZO
0PMLRbuPMgaCF4cvcTS5ZIdNFyaBrM2RKjGgfU6Jr9Wel01IuuZYgBsPSp9NkXND
ZjSo6FOigq9xxW965lQb7fSbl8iwTbJTIfKTWO5TGWhBPCNSkB2W+y0bT0un6N4+
JohXhNdEb/7cTQ3Nem8tufIiV1YOjtATOJkG0uxDfYAbPRRGmiYSKmUFVWW4PMao
BCH88W8Aphm4tkkgK2ZEEXcoNcIkmijEZhq8vmXuFfPBS6Gg8roR5EBQnioxAv3U
5o2fZJeQUAGajlKnxxgRtaeh+Ofv5y5cJpHgHYjHwdKelT1hCjc33d6aC7EkpROO
zDae19sBcqo7/vzBUrZNli2QEtWDlyMnn4OmNMaln3JzehneYe/JjY8JaKb3+jXm
NQAppMDDeFDsW5qYoZpoO+fpZs+7WBJ0AGLQZrXk1mxJYoB5YTv1OKzXoDUQfuJJ
R3Cv5mU4a5oc+GzIAta+aPKOriV3HTxiU6lDWd71GnCouCYtgv4F6no1aLHcdK0+
dfbXbqXMwhj2kWZ7Xp+ANPROLpDtDShleYZdTXuRXDQaKFk7RpgXegu8qlVCsXg9
aGx2jTxUZ4acxFkgp2TosakPpmTZTU4RMvy+uOLHheTr04iRFISiCG12fyoV33z+
99LKzgDOEmbIO1LfkdmWKxs8CxVJ4bqCeAfNt1ZonRRa6OPH2iRxZBW8Nm/Qy0Fc
Wm2uEot1CjNEifgXibASRTNfVqxMQd3ikNu/9SfGsDH7xfoexx2N+3rpvmHZR9Kl
ugtkQHXYkqhUH6zPbn7+Sgq/yY0sxVLvxd6yBVf6gtvstSamHiz1kYaj2cJ0e/G0
KHLq0kzCWzH4F+bHROjELj/80DJmVYQafoi+MvA56mubJp7UnMHfYpxKdFrAW8hl
/dY5qU8sKdMLyTF9v6PL/26Ljds9HNtTplegyZKDcfSIw4Fsz+cXSuqC9leJ7iat
w0nidY5Jtr7Hes2yQrk9vQ3c1NqrV6INMk55q7jfpqOg5kz0PWo0VdRuGoc+K/1Q
CMpxW+pwDRww17CLHWonntkOa8FEAx3c0a1e5osHkBWIaDT9tk2Ul2so+pY0gAy1
i6D8jshFe+FAhYft9TNUeRKVEIVPYfmPhvwOXlVTFGCKtyDQwlZgG1Oa769BND+O
KMgfwxs5p8OnHyjmkD65J1aLbP3N0Lpz309qakIFdXHrJTfiu78ycWlJE8mKm8QU
NaY5Q36alYRXLmZqu/Feuxffhohy5e1rpXZzEInBOEqDfEuPC+vwo0OVMsB4SyHj
Z39tFKSslOrKAk6TmosnS1kISsRtp3+lh1oz931yjS6sTrMxXlqd49hsuAuiADYb
B7t4XfCRoCFp0GexBwOUOg/+oJtMrvFtICkHI49+l/834Ct1Br80YGS2SgOtt1sf
JBKQOr/Mp4Qi1pvgSKTOVgfPAR84aAErW5AWR55cDe78scuVQyiG+/M/3uU4ZziG
u750VJKIa9kKn0/cfH5IIsGCECkTdprKWs4Xy1wR2YIyx9TFH5MswX7DM+Xh3Pzm
xRAdinM9e3RladF0f6E+zQicG1ognqTdUUTbsAaRZWBrfcaEbQph+D7iF5dlSN7G
lTAYX2EvnAeTyCs+a0+12QelyosTpnN9KHvaDb6ZiQGcooP2OR/RlMOUSFUYKLoo
DahlJ9lq9sJE5H+yyQv6Sdk6m7wkDjEFjGxDw86IT4lkhJu9bvkmHVMA6DbWvLsu
x5fnD/ermm0lTk9YHSpE2cAsPWpzegBaQ9ycOEA4ly8pArWyqLc81aN6pKsqaVUT
NdZQHMHFLekM7WbOaGKHSIrOYFvVhKVY/uTu47fyg8Oe/mbpF/VpAiOAyDEueiRV
dWkfKmGpkmEx/ACysH4gtDfbdlMANqXo2kHHU2JiReydeRIweORDWLoQFve1+vOs
R94avMHBRhojnp+zdtF5x5UUlME4UP5upcOockfrJhymjVndn6VaO/Ftn3fr4o7A
UteXx3yW4Ffa2/uA4n/zSeIi1huL6XcxsZXgCBkVXQvE6vFj7AlUYBEADIyDsBnZ
CVhbo8fCpr4bPfTKdLun4Yeso9KD7PHL/S2roT4DwfRjdn6A81AU3OLGXD2LgN5X
k9QN0XS3NzhTptSvUXPJr/+Sl7s4TnEpprKpEpO0rCvQMcgDvD4Z7r3djlTAhJze
hDa7oLMtY6cHTh8h2BPHfmj3x6w1Lciz7Wwu8qrE/8OOXvCk+Thyc78gPmb2RDv5
hiG50FvMNYarCtXvr3TwwABrd+3cCt4gaISRaX9toQEoq13yazfxz7YuLUZT2fTh
VNahuxxxHSx3EyJcl90MbWox7AOH7ko77bIArf5Kwuwp0hymALKf1qEUkl12wv7E
x0AZkx4EIAejLWMUZrNC/QWFqj2/yJn873b5pmba355uKnxlgiDgAmYDrPMIzVR4
I3zBhYLNyA72jfjn6sKbT99PX4A0DbL9sGQUgrpvXJgmkb0f/06tdt4Afrhc795a
9DdJMLPIR3bVxWn9bBvdbGpI8DdiSof5go+GzZpJZ6Sy1G45KCAPcjPuYnAcarip
4j2S+CzuAkKljlW0huzGiet23dg2zOL/buN/msb19LpPWyoUtI2RCm1M0mvPLujb
hQKR3w9PL7lGxy01aVw0GCSU/itW4DvWOZ35kIz4vNWhR5x6mxmhJaw1HOak+H4S
GtjzFrOhqjMbVM5qvAkaeqtv5gr6OXhqt8xNiEoY6NgprlI2i/xFcP7TNVVv5ec4
9Y5GVGsD6qFyX/nrDl4f/dTjWENQeyMWwsnX5TIps4Zuo8ria5Tzisn0cCTspsm6
IRDu36LFVWoa3kub9ynIk1Scu4j43IuqLyK5STrsyUUNK/aAd/pkZY5g++hjKREo
SCDgOdd8UvPl2Y5JnVbIK3R1EDJWkmhCz82+wCBL8RnDzc4e8SUbz43r5D8ka3B1
+7AQzHd2fEG05dFIETk5IZoYrOqACL7L2zrOQYy9g0vbEFlk7ywY3Pv+Fbzjwn9U
xAiTTqlGzhzEb7DYVshQ6v46ol02zDP/Xv0ZvjBAMwDcu0/uoALBgB2/yUHw171Q
eQ4fX5Pg6iVyyB/jsvvJ8l0FgtpTj3KHYjfPNP2PeaLeCTxE7PsKIYp6QhSe5Ai0
c3ykcFSqTTpdlT14NX+lLn1QTLQ9XnQOARs/RBwdXjw9AmYKztwmzCLpjAej9DO3
AmuiprrUlZ3JOgiNFy0MQ0WSevL+C3UCcYc52hbJGLqOOIJB6eU5AnXYi7kh4eAt
n7tTFP6LTywO9YMvWMA4o3CdWFkhH45TUpGZ5zLAWRD1NEMEdhhzDEEgLnm92tTN
+gPkh5nBE1F4CblbZGg22WBGUVP98eEMg+1HcFHkiEF9TGghK+/VoBxluPkp0/CR
M9cXxCPqil33wbx2VtpSsFWpKSJdcvhMGC0PSeFhZ36YKNrCripd7JfTU+G1JYpG
58tQHqOEjCf1AATHU5dISBbjwEGXOPexJz8Ada5uNrttxHXm+Hiz9sxwa3FBU5FH
Ml5AWOwaxzQVU9Y642wMyGG2MIHivTXlClGpxB9ZLZPYuuBM6LLeLmJ7tOtih3IT
+5h43XeriZkxwYMWmQBTRqo1Hjw8+lhcF80XbWmNQrldrMfvRAk3xsaAvJ8HIjqL
MjmoEBbnhkA5eQ9cXZ1tIYXuJTk+NHvBoDn/w1NgcFE4+B5dNF7CrJZkQvW4QDOQ
GYEu68MLcN2123WvpRm4jDUP1IsnT8C3UYO00kDEN2crTnkCt2pfiDwW1zDZdN6n
rwK2OfMW7OsMsnZkK/9J86gqTPWqDBIhk/4D0cPBuIrDLLNmWFIrAQ9tH3h+2qZu
Rimc2LRyFZDVUU2kBP5fAU+98twXxGP1/TMzT7U0IuOQe9YlWtnIjSShZ0QU5KqG
xPgpIibKjiNxplqzThP5L7ET5zG+KluPP//0viBe2o0C34xjGHDxMdAsFI0AgLX/
uDlq8b55nlW4eSgo6Ydy8cZI4TyRjStVqjXNksbWmWAoEr931KN1WJRF7czPQGvn
Q2OMoKmWMJ5WZVEnETmQaO+QVeJ8J+HyGXUEyxze8RLoDCJT1+FtAPgFhglzLQ1Y
QbxLA92XfGX/qXPXQV70aOtxXLxH0BclXi+dbkedch/RmRtMg9bmXfBSqapRXEOH
y2p0k7XxmpZvq7X/O9gIX5Ca7KhUbWZpuEUnIa+ouaDNggUt/WBPJMbTf64rTcxw
8X/At4JsZiqO/CMRWz75FopZZIBIs5QwleWJofZXhkvz/cCGZ495veQAynI2yebI
qMMHmNjiw8NhAO1l0xv2rCsyGBdwmOYrckGmw2XuXzPRhv3GSq3nPqovs4RmRPre
6ncQMUiPSW4mcyk7PzUU+TBtm3TIuFhm3pMWCnXxec+/YROi2igxfJ57oqLOB2ya
7WvfBnK72j1j9Sxf9sk5n91T2ve2Rh24Fes8m4LljSKEaHzn1FH52asZQycYcLGG
dKTQ8Evv/+hE5ls12xQbW1d7zILZ7Y1UQ/oc9N9lPgjQhwCLv0ZQxJQEGdEzMLU1
Sl3q7TpZ7XjnR+WI7SKSAMLTXSqthcbsQyXW8Jo3QzcRRQTct22PAoL9KLsbZ/DO
x8T/1zddLCsNrxQPO/raQhrH0oojmm8u+HARt4cb/mgLfcHI4dY2fOqqJtZysyLB
G1xXcehWmZYtL3mkLB90OfqMqukW0X1MRLQVZJpoNb+G56i896Appd2Mhzae67O2
bXdosgiaCG3vf/AAvMqwXtGpSqov+sMW5r/6EwOdKFdEHlChV+DMlDHSWDVP5u3Z
uJbvaP0zWnMH52SwOja47n/CIXbcyAqCL8HNWEJaEjNXJyWIpXPG0Wk1i4FPPlj2
vt0Ylp03jvtOHt6ODI7TLz5aTzhfUpsFaSRousmOvRBJIXfE6zU3huKjP24WuioH
eRmwDAjJTugm9TcFPrVStpK8fSSEEy+3JPJLR2kyDi3I77L79W/bGaEj5lT7B4Xn
MFvygSxcspDSMxNa+nI5scf9mw4n0W2tntnhtkaesH4YqyLq86nXcsJcLkp1kgV/
VIoOP8I5xX4MjbMxgtGPS/61bPRG2cpYxYw4n/eZS7DvqOx7ziW8T2+ZG05Zrzl1
7YJXO377HEyjh+BjFRGLdG49MqBY7QHibtu5blL7ofjwBl5Gw6YZfaCUON5RagcT
1BorXDISmYd5u8UdBBNf9YBGWPhxBWyyGI10Z9ajtPY9XMVSPUBdCpGjKYvd+p3t
2Kq0fvncZF4S9xkoN+amSRVbvC7UogutYm2rPyF6g6tMnM2sfmnd56sw0m1pTTUs
ESW75C2JevI5YUDG7Tgr5g3RrnfhT6JOYP0BicRP2s1//ZiZS4SKSbzo61wdAvo8
+ecyG6JHwuruzHch5OD6G6IYlhMHk1lb6LS7Duyq3qeP07Sn6nuDcgkua9iikBws
x0/Hdu3VTWtxFlAjFWnmKLxPI79A4fWd22E0BIMK9zQ/09eqF4i5yU8EJ8k+M7P+
BnckH1KvZMvM5L/3v0dZ+pgxj+mPzv0cV2c11DMzlUpCDmd6V4z8QpmxWiF9z/eQ
04Ah+8cq88DmfRRmiFK963A+eH0F+PDfd1RPNT9u7V2wObJpUmzHVcWQi8hosIKu
vPjhfKS/UiNvxOeKrh6zAJM1mU0Qym3Ek30Vy8C7SrCGQxDWxq2IAVE5c5s980rx
rXdr3XlFsqyLsKnjf54doFcQYsmRWy7hfBjk5/CvriqrbMElxZGifcediOpnGzgL
zIcfG9WJYoj0w1KtW62PChh5jJ8hxx8xxS0u4jz4FEctzbDg0hufcZx0/54z/STC
2bAv9b3UGR0Plc+eIxM0VpyjB58C4xhfVvDshpKE3MK1YeGPDFl1u0N0Zn1bp4dY
SzeOVRNGoTPNIK3kuQsdUwl/rWvcmrG11BupO2GcCuEa8L1wFVogOzEMT2bNzP4S
sfSzCFrQ6fK26wcSd34yfQYYBlGVN5DVfoMw2WdsmxC/Z6sZi2bKVdOSL+fns0AT
Uo/kTpiARJvz7/boXm7ZLqScp3m7nuQdl92KBchweRS/M3fmBghG4O/BLtzwkvOU
AGRHcbs89BbId3nmqHk9dUZlae8Pow/nmYIrU7Mf2ZOtIHYHWQyiO6lpfWPKVPPr
FIqaLAOgf9MF57yWi9zkvf9viiwd34oo/6k27R4jmFv/vPg2J/SOLo/ibqU5uw6W
5lqan+M+jttx7EHXKBqJuDcsWiRmoTEcBW9IfqK6c1V3vk1wzMHShslGnhO/5RWx
ZL56NfKGfIlTShrtEXpXZgpxm842iomOaBVXPFc47AiYqQw0YiYHj4DvLkMWlDRP
4FDr6F+6HAiGz3dCm6R33tHp+30/55L9dENcyhqJOVAW7VjOL+0pzEnaoFeDTVIh
521tPChzFior8isIT08XZWmoCZMlHdRB4UM6DsKBUDw3kLcP141v+bMDRjrZWdW9
iV8yMEJPmFPWcAHcgEn4Xw0LGPEjG3LmqgErwEThdd99VfNf/8GVvMg86fHyg7MT
f5BBL4aA/alUFo/T5xO1+T7wRexxbLe1LKEw5ZhGbST3LeUfW8WFbYjML9fsfGx4
DjBfkoEexjUT7DmRjMlaHs4tfL15MC4C79pvPB1iabOVsIf/iuD6gsg+NTjC8xY7
+snQt9H4fKjbJT8nvU+BI0l43ZrJUndMQqjsuTiPW7+AJETSa8Uco48avnG6YSmE
do5gNhFcBKLCV/+IOBlQCmuLHm2bN+cdAHVhsdoo8WXjGyAAnJWxl8fSOr5uq4IL
0TeHUj2rK7ndPFHAkvuD5xfBDoMu1k1LBaGmKEYd7TlvQ8f52apglLxn4ZW9j1MP
ldcUSHbqWBhThFDIwz8R+WM4WnhutiZvdQrAocUsMyC+qG17k25MQzSWqyfwmQxS
HFhg+Aiz1xFKSU4noctUI4m+JfnjP831dsbZjGxi8lb1Ox9M4GPM6MKMkSZBh0i4
tLBKjaUTj6dydTrCcjE+UuQY/mCN+KdAGG/VJ7X0O018YNlqj35StCBXa2SuBXHe
FEVEDMhE6z0As/vDu7bNqtqs5MEWz5MYsraNdyoJfsd0SaymQdYoOZCCpmX3KzZa
dAlP/ms0RpisrqbpRAxD32DEcXam3r3KSipinG3tYtlG7qi4pBC9wytQR2fikeEs
FPk5ARj212e0Gao6vufsjYBzLLrBuic/Mve6+hA2Hnv4ZDa8A+syMg3d9ujUutRC
c/qIdF6zxh91JojLX8gyya/o+s5yFbUF8r6+Y+NvKmDite6nviygnd7StEwiiy7u
1l9+An/3J9E6XzrrHin/JrgGDu47J2Dj78Xim1qwrrAFZ/Ju4RAaEUNr/khXBzl3
nDK/lOSEvGqDed5tCn9zDf4sPKv2A2JEl8Ic4LJgtfSfkARQFVuhy9ArXCZ9lSu8
gJWiNcldrrYUGteaywU72+92rw2S2ex6cpvErgkd5NKlSVAom+cB+5dp89i2CK58
5sIHWWxNcCB+H1C7KBcbmOE5H0n46143YVkwmqVQGuMPnLsLUXdfdIAYKOtmo5RD
Kgvw/6S6kcmn7UP4sg9W7rEyf3EO+PsNdNQi1qn5+qq4J6kBj2113aorTjAVAKT2
xhdi6EmJ3yWUccZkHXeAyZZ+oFL2L3bfbkhyp5XX3xKEWaRaNp0srZkHo7DpAVWf
w7Lzkkfq6FAcJ6uo/BA8DnjbjTa/wFX86DjpJ7sEMeC0C2EWnMJAcZPlN3Tn8ZWv
mfNhqCENNpwQiamrgM7hkQBQUqnzXN1r0WLF2q0rflsQEmxyU7Y6lA7IrelYO1UW
eJRZ93kExDue7prdxrC604QRYpeSxBW1FHIbPfiqlifmwBsz4XFAAwlwi01wpFR3
6O1PmilPVASgvW8Twi14XNp2ClhEQzKK5WQ/D9cK27ooyP7vFVV74xhtVu/RUYmw
LE/JfYXvWEsq7GAcQy3pxAUdbC4n/OkWcb7aVn/ihb7a3I9Uaxpa9ox5M50eXNRb
uATxoEf8EfnxqCtpb89zw1q1NSZfnpUDpkp50MpVy/5wLmxnHnYe7gwUwOjJgueW
lPa+vfcd3YxLekaYVLsrL/nxKdHDD0el4Mrbp0IVnFVJ1ZT+kTDQpzxFxyamUkQh
Ujd/yiBzRT5FpxmXU4Vl5SGSqhzu/cwHyY//3AFr437KMNeNsSTDbElJwAZqZopg
LLqE1VS0lrgeatxxYouvZK1xY2cskuZ4+qsUDVlrOQo7FKl++c2ufeVFWJ8EmTBU
Nk5e7/yVfYoa2O/SrUoT+14TLTYNGwG8tm38/IMQA7OMYznEfp3DAbKbpGc6Er1E
k7CmuutMhFDX5XcCgLbCpkwkPRZi8LtzpMbS96ophAzUXifN/ENrPeVS6+ZR9IyY
EO1vXoFiiVdE5GSjrUfTmF8aVxxX1sdqy09zowHazaDBfrDQd9yDrQgktTcAgWDt
OgTJ0Lx8DGaFqK8mQSa9+qqfLyNtuiK4uwZE+g545W9cB0nYxfV9vnoFsCBR3av1
RXfLBZ8oLvc81jFAq5wvXdOAjC+c1zQ5Qj9Rw5TihDdWNk++rykZad1h/0vs+C8c
qh27qS/ysWuL0OuP6S6WK3pOGdoeqvbP2Zm4JZGZBJNT5jD/BSX000zhj2dkGJ9R
RvuRr3R/rn/iIGqGdU+B7RmVvw4BICWJYFrSszl4fjXh82dhu9a2NNNLD6r2+Akt
GWMMBdNlYTZu2vBfkRJUCIZUNSwQmX2xJeKDo4eEbYZGWeOKRiC+hLqJWRy/2+lg
FEwkv1obCtr/ld5GrA9rD1e/fY8zrkyEIAD8Lv5vCLyVR9s9fsvVbwVKP3/etSZg
A08TZSqgtC/U8IRW6oC/zmoMSABA/ekEsGvLT8ghVZgslA0tO4EE77MXBOL7jgPk
ttqypWZSxXTq5UrdVYVeBR2jhUqlI5tajmx5znUTZnpFDTyMCV7XwOg47R/i1RdT
Vfsfh19OtSeYVp+fpK2KoW/Xfs9WrCFNSQ8aN2LRL3Y9vSXfFtndbV2qsD0C/nhD
29eDd+Hc+idvy93yR7W4ZaoJFyXD/8cpyYtGmpCG/olw0xFm5o6Dl14qQ+ti2+Pj
4pJPNYudF1ImJvfCvvBqEKYRfRP/D38DG+P589n2gPXx1lIfP1bbhBdYFh7MhRvZ
/TiXjCA8bYezBx7WqvvTbdOKyypQBZcnx2+p7wWMcar+dIsj02iv66yGcWJchGol
BphnxM/Zge3BhzgO5zUDBvf0kh33dJOjzkzTRH9vEAEndN38ZhyMKWR2vs2gTCXb
noB9/CnfD1YO9D1p2dmzrpAUhCCpm98+LMr7dwiyooW9swd09otL4F5XBFJV8VoS
GJfHuTWzPNoopH/UVftVraB/oUcckJIMdmL7eiT4cTWya0iuS66b3li9ow+V8tyx
Mc6/mFlAakDkGB5NPsYaSYtsS6llxCcVaZTPM36t7D8WpCE2gtk0VJv4cXojvOVK
Zx9BRNELujP0kyQmHVjoHJeyRwZOK7qPcxYcOLpJcNDxpEXPKwPwpaTdP27c+YNE
eBdKcMX6ME5gHGtBtegzTcoIToEyTWSxOx0IELUjt77mDyAJIgpVzxVzO22TUCX7
k3jz8c1WuuIUvrfzy4OK88pammRF51jz69dLlFK/0AqiJHulgTuLiCNhOUX4TnOZ
v8tEHP6SxKaJZBSbt0CF75u2QPC7iZdGPSO9xkq3Ked6nrki1sWffrM5LzrVo7+8
/u61vDJbRymo5PigcZhuQ9wAL4WS2E6wWkUapaCdyTvuOU4IbczFM9LL/H8bfHEJ
WcTsk/WTZvEIfgiRWkHmbPovhloWV34hUfcwdB0eRo1JceNtXOcGyVu60Mz0oxZK
LatoNbmTRUL1wSjyv+N5fNdbpl2WnKo5AgEDwxRMxTYY4bKbivNBOzniO5HlRQdo
Vk3yLV3IOsOhNXOjKTApWeximWHLZojKkO+1e4mdEPLsTt1wmvCRH2xspt9nQzqx
2LPS6G3ObCqvptjp0ZGbvMUYIG+yeaCDQj+HphCKIodXVkL1DE5YNidKmYbl4OP7
o8FcgX8aVzs7arBVaWL39q6yYvKqm+ekRPKsjahLZDWPq0aLaybqkw0pomFNnerF
HRVF7/u5y8R+WJWFqPq+PU5MxFkzuxuL4DbWIk2KdobrqKQFgQgOI6+ndZGydOJ/
auiiGveBzlgQlSG4bUdtamxeJdAsopJjtk48nDp2B/S8VGt/alvl0iqrE9HU1k0g
dZEJCqVweeJnRiMgkQRe6NA3ojg1Hl5O9TzS1nflASZIPbdo8FbrwRtUTnJ3OfsQ
h+PIh/+GJmlZo9I9J5UnBOepDpPZAMTFUndN6HxWm8wuDx6KN5y8I60aQ3yNpu2/
NE47mYeCPrH+hppoqFLBfzaKBNRlAMfPovrBFAnoJZAVtAs8kqRTkpGCIAW4MoYk
PoN8v3d/SycNVm58paO8aBKE84VaU6lkpajjoG4WehRgVGPpHUF2dfEYXkjN4j6r
lA9gWCZUNiT2OxS3o4lD/heDGf3TwoajHa7U4LxYwNKN1eQFElxMR/VjQdLJWbGX
wLYzvcLdU8g05YSW5DW++HEfQXHg51mTCfivV/DSPDepIbVTt+N6Ze0I/lQzcQrY
kr3Q6XQwLQAXURGxtEcdKHVk2bA/lqWKxDhCjFx4UZQ3egcgi1sj/Ai2vc7yHUEx
Gy2THyDTmTSdNuCx5no+8nCp7Ivsye9Gwb3MxbKMBtHpNSwb/WQRbG28EZdOcwem
1gp4Nz6rQWlAJEZFnVeUzJmIjgWYWSPXkkv39gcsTr5Ni2g1ZeOB4x3Gx8pUkUQi
FcVrrK2wlEJOLyVxLCOZ0coWuktXNUjDttRXDkqyBakuwuoS78lylH5hCwWkRQMV
28L8zDzbI6Cxq6q3zlZXv6iN5rla1dSQXoxLrB7TbsfrLrfxiDzUQj4TgWqcjpax
u1JgaCrLgYpx7DcSydRqBAcnpF0pwejMW+kg7NY8r4BxrwFey6c/VjdFUiwk4qVh
un7QPN2lrK1IjRRZgd5MgqDUl39ot2pCRTqyxxHDAxVyzQlt+/H5gJ/RLD9IJvig
nY5AwSOWtSC3hLArBPrzyYyA7ba0YnG9hKFPN851wygQeRaqKpjH7zjW2A+qcgUN
4JF2bnl1Nlf2adt+TnXo4HgNkUGikSeLHwFsC+ScBlRxmBlPmlaCig3UwEEgNASA
bwsKOEoA3pNFGv50872idvZf7epEzb7dO099ZxJEoy1XYJOBQZBjhONsYcbr0a6M
IjCXJxZKpW8bt0Jqr9/vqDxCBqJwzbxJ8GiV9l2fDU30hWhUGq3Rz0zeq72Ljdcn
pUXL5RBlFfG2jWSrMAGGcJsAizNwvnXy6+h44knUxFkp+OqsNiKBl5yvoNIoPiqu
JlmNr73W5T/enUgOm518j++NV9doR8xFcP8oeyuiLquEFTR9vU8babMNuMJRjPQL
wIeN5dXTdLhy1TU2JM2fA2BW2X/Ngr5m9hsSTBwaOe6plwI0t7KzbVWiChBdd7Ej
kkwgLLUqoriNvdcoxiu12l51oWg/mbckqQRG/NjU7aP2Jc55mM5x9bJ+uiw+PIxu
mTEf16doO0nppcEW/HxamKM1D5FiWfL8ZesInVfnWs60RZcNpTIyruMAqbbzVd4N
LhAZc8EOjVqC2FGkHmh/qoQSLkt0zZ7QHVDNni765lObppLLnZSlmBopMPaNxYCH
7rVCYVZ5816HR1xBjT6OwpJhJs0orTaKV33hTpmFOqIuoKf8KIoDy+yLawFu0UzF
IiIrG1YGWjRsWm26KSCIC5t9noQ010JE6DV01M48Eq0ESbq3YeXCC7HnKKabddYr
PXwYOskCDCse7HAmt130V5c7u197bUiVdND3P2jqq08hhnimy30O4p9MuGeIPmOD
bz3Qb3S5Nzj/VAjmzn1xjzy4bumyf67Xyoz3QSLyqF2vnoCqqp/C0UDfXpzD7OSt
Rzi8gzpOjqvMXrjYaifKvkr9TTydTh/ufYSLQkck6RunAB9tN051GitBZ/7VC1st
rtXwgeJnayVaWNgtTAtgNSwzL5dMQ3tsFY4QPQ7vmuDggg2tdKfVJTSvq5rraSLA
SgVE+ROJUHUxU+q9XqKDz+1uNvua3L3X9ausN+57QyOmXQGCna14sIsUqy4kBNbC
nRQlThrGpNVLzk9gFE2QLnI0gcb01arXMbtgtju+gbEhP/hW5UZmWlhRIIDIMRva
Fb0bmCQxZ5nwG0tsb5FpdFnJr0HJQp2Oi4XGtTv3QTF+Wx9Kc+DoJhqHN3BWufrP
oCZ9VCrUtEeh8i+kxVYNW6lnLQxOee78LuKE3GlLdsrPX3fa2MZZlRZ0JqrcBsuR
xoHZ3OWBWlFjVb/Tv6oaLuwpzlA64lG11r239GDfpVm2aw+EHXTxoScu4XWaWMv2
+qnD5YXyMgFUhOyO0K2hE67on6lYtBk3j7JGJYhwxQcwLxAEZp5h3C0P7kBtrpd+
s9+pYz2N/BltuQsygDQaIJJcwVwE0cGRLoQsZWpaKVr5to5uOamDKt2hwKTdC1u1
zNzJmrXfaP3Ap5G4DrR6fCTF8xpvNwGB9dmiukSTrAoOxKd4jZjWuJE5MBH65qFi
HxMpTGHtHvTxPqhzj5H9iOVuy2gqpB9NIdAtB0q7rHyymT9vBAFseXlIN8oCxIaU
HiebMCKkKm1lNBsI8luFjCduyaNe8f+LRTf9OdoDnuCYu2S39w3CEwjmcZhvixPb
aOFrhBxZbeNyvKYxGvih3ALYFeIq9+x6YboN3K7GcjVtFdaHemocYFkRlbfU0TYN
jDhNSCjKxvJlxAYEhFnS5LXW1LOZS8b8+kNVvdM7agjHZh5pVcbZJHnMu4UxeRPj
/zw6smlImm10ZD8Us40EOleSQXEpYFAVqm8TGCvmQm8qE0b6nyOduw3y9zFkdflP
ViPCy6EDED0m1amJzM1bHqMZ/cA/fo8slJ7K89XEQgxoudcXPS1MI7SssP8aQb0O
OFEaycPyA2AVtsBekXJj3eHXbRJG+bMsosAc28bBwx/FId/Yi0Np1NQGDnH/z396
faypVBQgRN8Pd3kPi0G1Q4tV+Fkn/zRlZ0EkqSPvlF1S7J5/VXtVtZDYPTTEew3D
a/I8+7OQ2QrhNkUFnVxDx1N9LewYy8Jr/Wh5Se9aeFV5FpqoElIsy3XssXtd4wDs
2Mo0OSUq4Z3qgzDUY3/nuqy2ed3ztS9HCF233X/1g0zMcCNmLW+DsShHYVrXRJnc
aPgjIUfDcWxz4pcE5NiDAuqVWwfFAQ/w3N3xryq3bNjwhoZxQbyYKzSSBfDYFPwV
tvV5RU7Tuh2n6kgKHoj0lk11JTQfa0cueNPFyWE4+Sf1p6MjvWDBm0EKntDCTs7e
jNOIrAAMviKoxNYCWZRq13qehgSlSgPvbd/BhXf0qoP1rgvWeV//EkvDat9Rw/QP
JaG1nIS5PGM7vQZOyTmJjxYppvVhExPaTpdGgON3FfJtb4JlT7ObDQA/OlNqI7uA
pGMY1JHcP7FZOYYUdXLoPU3ER/9Q+r8G1qC+RF/eliBGhFe+WBoAnAFN4vwCDDFO
Y+HWt45mHucT6gtwqT5xO28LHxcYzqrLFpCBA0HJHXYITBwZJGvh8sZP2g3pQVNK
+YHFGx100BYhuVhVQltNA+rf5UXHK/6TIXcEjGA9dUGpjBslyJ3HIhbLurPBYoJf
+zSziDxgOwrauk8EiHeHrpBnCjh1IFweZ8oeCnaPkY3Sfp1gCwbKJhUzUuEPAsOt
wS+A0y4FxB0t/psdGyXSNtws8F3gDV1IqL5k1AnjIErQTYsVT2LbAw+dclBtuVYJ
PuWnaPxVREbnIAVT1PZV7PvnbiNvWCIPdiKd+G/jiRxOFoxwrWUokUY6GM95vYBL
eHUz4/xp8QWrZ5ny9H7ZT4N8ChAfVKQ2kN1sYKLzz9ArnKnj+tVIzgXBnHw4cgb6
589g6OYMG8JFfluHPeKB9KKZBkFtO5Wd4gCJyCpKlwohn0w/JfjYmyQ8DpnPA8uR
I10M89oRpyqTC8HNGHcYQ1uc/h/pMNGzV4JbFScRbOxTk9Llf6FYiH8dGA4wJ/Rb
Pw8Wex7ECULC5DXZlwa5wNCkjtJD/4uPsAtujHHNL4uXRlcvTxGqFzoF12uQTf2n
jcSif/dde1RSepEsjVsbOQz3GLpCehMzX5jNq+4wSEOZEnuY+m3y1+FLRbFtaOHQ
CIOvP8QxEZIjPXO6rtTR+mviXO5vJoZERIfuU3R+nIahnlC3RZWgDoRwoIvqBuFU
VYds5mXLBHvuOSYpqiebyH2xse29hBFuOcyaJZ/ABS5sD6iD4nkiUMi2f8sa4pHh
cHlP6YLUcxJRDTiQcV+UsRJk7ueGI5rMsR8Cl6JtPR+qqspCI/qWLfJJkkWNVyo+
25/dk7bJ2U5ROH4yYysFJowNGpS5/3XiugXpXz5b9i8B9DIGSEWun/9Yy6Mjm5BY
8KxVOLw4RFaNu3bitI/moyN4WALCmOl7F0L4EAi/MxBUSQrgaRaclcv4+NJH6Y66
DT6+ZRIMuEikyoGP2vMRnMt3mqz1g989f2wEF2r+e1U932agCijS5S4UMKrmVWgZ
zXMl8GgqTIBL6aUbKY3/e6yZBsljH2jRDFcyzzBWSLSd2CNRt7aOC9wKabGspez1
yP1OlM1KHJ18atqTBJ8wiZeaHqzjJWd/vTw4oR4w6+Asnfwb+MJU9UhNyYzUHT/t
GER0BoClpML3qm60tpxmSJNr0K3pV37/WpbaxlgBlZUdqhwIZ2IRJ/UZ+ZZkMaTX
jyCHTBH+54N1drpHziohtJwvRS5JIT4uK0JDirJoJkLb5VaTr9HAY6kSUVQpkqxh
QA9K1PbM3fNFccUZapt98WnMycOjxTk7AlJKzAes+V82WfA09BW8g0aQ7Dw5Rr/p
Kif+0HoJ7lDgiMOAnk7PpwPIGQtsM1LGLL3I3zoaYJEG4gMgWadvO6qiWw7akkqb
JPnacciBUG70Gv1cRL7sSC89KuhqKa2cYkMn4C6QhxQGeLbwSKdyy+81KV/IdFs9
Drg6F5CP5fWmlKlhqwsWyRVX1pNytB2LjpTA6EkTwc8SR4g5RIu2/5nwWqhHKQVb
s7bVjGetEW5wpvUZUhfvH7HxQ2naidCejXbZUSkMLZ5zQLTCMqHTT5KD8k1YdIvq
K6W0rM3TZbTx/IoF1BSoIP9WRjrGCTTTQd/yKfXLkrwE8Qq22yheuN3moHbC1t8D
qjLQ9k6QBrJqSGFptSp7m0y+NgDvVN5mDy14albRuMcTHtzxRBgJECYq7DxqhKRw
Sdp29ECr775/FUW3e0KzK6ii6yUqi+7klkHnm92LWOlTX5tBkFfMEYu+Zt+fF++h
u9vSdFylgHj61E1/Lh6Q9ePrFT+nvm6k2QgIMTu6v2kZM66Gt2d0MRI0UVHUaYPV
yIrTqCdA11i4dqmS4nWYwMI0bpS+Nw9TiVAJG794C/pw6H0MOt9ZqMjKmbsjrCKe
Qb3uvEpBhOdeivViW5+KGBOUGk/UVgwN31Fx5IcN81q+FXzYh96NfiKGReNu9Clh
lgOEep9MKBFGaE3IAcj+SphZNAhXkKVzq0zw/sd3p+Q59uqO1dwslk7qGBaWx7ci
MegVNXNy93sYnvVgvkGi19Vr8jrNY+DPGPyLT7EwJq0qNvFaDQcHp6gn3HMvybwB
DNiGWeDjojqCJdmZpVumvNQD+uW0BEvw1lVDCepi0S9qY0CMI7r00AfYYYyS535L
1zELhR8S8tl8xoEc0baw9T1VU+ZY9EgbN6dOO/RPJfNA3OcvD6NeI6s1VPEbgBr9
yRM3q9i93il/nYZhajP/6++vyB3LY1UIbUvCDMOSlulmkWcq1N+/v78dTfQj86VT
M0O3cEXncRsdxNVrZRO0vosxVMUkUB2d4NOAnGe4gyDhlBvVYgxFMmJCpR/Nq/Gi
VjuTDBZWjSpUQJhFbNvVUGcbry/z4Mte16SuyvhwqgnCHYng06fI4TkeSRgiA3/E
/ZuCKnTEZmx3tNJQQIwffujTHTFdnkYW1Kscyqji3edoOFakxSsGFE/G/JtjF+ck
XpUFSQ5ndHLQWhB3yMNInckKBl+lDe7TI5DV/yRFfOct8904U+er6FTdh9yOFqwB
2bLINmjOnx+F3qXgXEQXXYTt3R6cNvGFFf1XE3Cyizb71pAJKP1+xb6SeFM7vGoV
JDfHsA7D81H07MekyH+24Xy87309rzpo8In+P431frElYfnP5uRaj3zSwKi8S7/E
ywblriFYfc5ZL5DaDwHB3VHRYOiJ30Al2QGTygQK9MV4WCOW1eHYPH9qa6k96rqJ
DNiHGYsLlf4qpe2ae4sCsMmJrnzIt4QepSYfe9pnAc+h8ZiqFu6LMd7cICyh/nOE
9D7tNpo49XSB1rY70/R0SEMEj3m8TTWU6WYSOQTT0im0qb8vvEIFlrQtNrEAvU0D
yKOjk+XwhPRdNtYjaEIFOFHuoT8oiP3C1tn1nqGO/R5oPYuUV1yC74sRjc/98Wxq
eLsv6T8d4GkLiHKk2WobMPsg9ZMSJ199XPW8/KltKSYtE6w9Z8Q90/48+MC5GhvJ
d24CQlKrqw2BBOGB//708l81kuPKe0u9DtOiGBPKY2nZlG0Rty63Q3G3ZfJZnt5k
wWmfoSqA8UZczwaiqffOKswsCX73y9ylYD9NJTD+KR97Xk0PeOx7r3SJ1OMOmVVd
zCMIamDiaU15GOQZcTLwsKp3b9QNabMzsgQtdRxEQL9q+d2u+gwu5rrCawKGOmV8
rcF2y2OhKT9LI5ipGMiwmIn8dO6dU+Y5XIwctLPX8XbZH9VrAgrPzv0Y8O3+tH8u
iiseeIP6ZBmY69qobevTlItK9GqiPRN+fg+fC4syM4ChAOONqMkLeze0J/Cwphc2
t8gHMunqtQiill5qJoUER3ADrgcYdoRT2oxiJgrooS6lN5VqwwIUi9Pb9yrsvm0q
B8rVO84+YYNjkehRQBmlVH8qRe1qs3ESDgA7n6+XDocEeQZxDUSTPhZFAfRfUwdO
Z6JZe8vh8rxxZXqMvxfn6mLQRx+KCR8imP2nwBrhPI1qLHo9Y1EWq2VXJRGf4cXM
d37yj5FOZOqZvmXoNGHL+r4FkHicnFCFmED4xJnxux8NKiDZZhzjSnE/LFEucOMH
ucCa5GIYtj2XOrnJDoLka4l5RDGNv7zn6nEW72DcAqiOCpH7nBnD1dDCw00lRpzI
xHTEBJkqTqEXakhmCHcd4piPnccOJ+cqwpbt4JUREpykbu98iHfbshepKKFUmRWg
EfVK7nZP7fYC8WqZu+QhIbnRkssGpag3nC6ymFmaVZmIHhHF8hVu9c69+U833bvb
C7geSCiZec/yokva1Fd/rTq97d1EtI9aZaqomh9XU5iOP8dChFRjnzvcD9rv7wJm
xFSjSyK1UOqrGRCJYhWoXTDpPB5Xk6XnB0sUTRrQBR6Uf2/D+XbjA2j5CiNKq/Gw
PqJMOi0Oi6dqy4A8fGl8939kvrdXIYarC4Co2MRvrOrT/gqsZ/66Si2ICO7NQg+A
fZ42mMJoe6FIjy6nxHMF6yrhD3rkJY9cdLnontO+5WDoecF2yBnt+XmSNS59HG0o
J1OeCyR1adUlNo/17lrCkNq71Q0XZXBqTRXl15iVezDm5dPW8YYd0AxMcCel7xnE
9kRckrQWaKeInN+IKG8BOe5geaupSpg7bdPQLcKZKD2UmdUtfQBeDoVWUyyNt2Z4
jQQEBoi6oHcz5oPPFvP2jmT+GOM6OWQ5lOG15bd/TWk6NdflHjjiJs1p7AstRR6l
g8rgHYJQ5lP2dOn563J0DZUZPxLrHqVdOpigmJmtsQO+99sg3NORpEFb1+NOyzhH
WfvSEOyEZLrj/wR1qKmhcB9ET7+Ub6Rb3pA6h1i1aL+KcD2QN6W3fhUHtEkMHtcK
FHSaSk9wOSFoRyZB6b/Qjw1sSR6HOkaUSi6Cwn4vmye8EpoDrzx+uOLQJ8G799W1
QBb37arMVJSg63uLupuI/A==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lzSejjfcWyOfI8KfQLDIi2GalvHEyPBULZjbjIfhRRiivtjV67lsw3h0NqnqpoC+
h1nio8MZbfUr9OJi5MnrA173tgqNLel27T8c01QSuZXuFpxoMAjHcVzisTE6rTYe
m+AZc97H3bPgEXsiLIPcP7QOofEZGEWRSgRg16pk+GydRg1scyRkqtDf9P5ANKHl
gmbNOKBNj00jvYAWpEZr4Gfgq2tNnfLFN324HnkdwbCulMUYfpPsVq9vZ2WNw+VI
7QPKHot76OtDE0IKPOeFjknNhOfWTYHnJH1Ph8AEsQN6mq5CdHZzjtNFTHlG3LXZ
cYMB31Amh1mlzuw+jUXgBw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22144 )
`pragma protect data_block
PuQgrr8ipPfKzOEe8fDcUU2FmLrLa7WLFPYBUSVvAOTqUwUm05iUoIw+AMu8onMF
7PhOY+W2E9tSKCLV+YgUauOfqCk1DTncuoFL7bFtWTDGh2CCMH9nbFH3Lx+o/VxP
hUzXQL+5V+3/umfmF7/tDtl34kywH4nfnipCWeWdS3XZGHR81T7IrD1jEKrzFhKF
0kHTvDI9V3XIwjBrVCWij+P1oAaYXAcYyFw+qr0TelZc9jpTsGU+pgyIIxf8XS9u
11f3kGjOXwt0zx5KmIwv6eGh7jVcHzdf3fSC41u7+62IlQC5+D7lLWH/4leeP1ob
dsgwgRpIRjsvAmGmd+Be25NgeH2f3uhc9MKjn/q7TNAx5dGOyzFQFnvxdou/IIvK
c2lrx1G8yo8v0dbzfXAx8q2CA1cj2U4hYnCeUwdlmVrhD/lTRbAwAvNzzYDjm86E
Khn+WrF5KHBGAfVuSSiHvkzF+2cnB7AzlpMoh3+C1lqBzEORHY/xRNitkVDNdC0N
9tNHXZfiMuWZOen4VrPylhK8dV3m5MrEaxwtLTYxKu6NGR74mr8Qw95hs1oretL2
Y8Y2hJc2BSe148wMt0qibKMCCHa4cmo8SE3gLDo5huguGyw8j9Xk/U66kNipMEn2
p57W6VfXyLICxbEQow9Op6YqueRWwWV7OjEozJ27Led9IMfNAbAGUVqVc/KgPQeX
HHxEioz1xaxebXI+sOl2JHS236JkgU+j7ceWfVvPsw6efTb+DXLP04TWiCKvrLYJ
xZJ8pacBzmPQ+GznIqCCNAHQqihJl2XDExDUsIYq7JkqUUZnuP/JS1S/hEGSBnia
fgz6hiQ7PTmgGM6JLZufuFd+26+tTh5VHFlCiC0MiAlQHQCMaTWWdldYTJyKRiSk
83sOPGi8fFYMSTuhd3JKsd4XA8TAtzepe7mHn/gxos9Yv8IFgTmHB43ngspiZ1JU
CFeVxS7JVwACyti+nygYWtyvvbCFPNtTPxQBbnf2SiQdFcxuOsvOpinD94+K/Va7
BE0T9mUkaqRvPnXXSmFZqpezwy5NCaVBIr7vnJQG6MwwApb417jzBur/7SLnl/HM
HSxosibPWDOgV0l1QhVcuc1ncKfiUV1wuUYCUM/eJuUJTviuB6Bl8uAsxi+m7Nlv
dAeBl4A96M44m/DN4NND0W/tDyXwpzqN5nMlybXYilWv3QpIw4FgaT00rSwTk/c6
QmCZrR5XNjOZbgWyyJl5lxA2WeixY9ZhwSJG79euwtG9C1a/4H84EPIEsWp1nHnc
zGe2efvPVkRwTWdEGU8GO4hpNYVXIKxH6OSHOgpjoPMqjq/cUmbADBrQLgNgrBix
1tgbyWezMaqjRIVtHWyf+7hKkBD4PEPzrys78K6XD8HrvVvEJUAB5lxP6UV/ZCI0
cxZON2yWfOMExH2SIgfmhSx2t1EKn0kiANO/eQXJEi4wZfFcwl16A+ZcafAbzlMs
ea/SLL246NKMxgBcOouurfYvNEI/C4GvowksKu1dmSFg9Thzf6/RC9GmJp/ZREz1
/k7nsqCQQcXp5MWmxkZomKVRXXmGpVcz3bsvygQt8AUDIv/DZZVQan3A8Zddc5Zj
LitPt1uLQCeLmQCwPfTx5hArunFFKoYCDBchRjA2k4apm8g1K0IcK/C/fORfhfbW
hTq0hmKCgMeBQnSvA9Z8YDtbmknU8QW11MNVWI6HilKlIg4LwC6f+PpZAxeWZ4da
ntdoI2yrqOoD4Et47qlqLrwp0LjXDLceYC3AQeD14x/zozB/aZi9i/0+CPkqIo7k
/CcPmEh6g1oIUq6VWBJrkM4muNxZnrn6F9WVo+7jVzBXr+SRhNlKOF/4iLLfBxzw
x2teFQphHNAkd7xqtm4BfXcr4xsABfzGkZy3m44Bg0TfPQ/yb6WQP3vWAm3ke2cl
Y9Cnp5sZmq6cGACVJZdW16gXiYAR16qfXlp5nZCLCk37PS5kcgb96Ihpk71bwqTw
syrXbf5BPctKXcwOxIto+7M742WRnrMkhEKNptZngHeZV8Q2oGMRVjKXUN1Y74s7
2EC5BAvnVEvph3fp/yZxTLY/j3hz7zfwEdFyJ2ZnMY2zArkgDsxNGXe+YYnchH+B
ZNhYumg/n4A5bmFjyQr6gJrrWHD3Oy5tM5sHYjBnm1KTe6wsYPgDtkwZp2uYpSgS
Pt5TRZeH8kqqPxFFhq6xIwshinGJyW69wOegMjr+g2XiNn99q8URdv89lTDbUxWk
tOWdbUAmNtXoqeYvNQ4O9k0GEW7aVum+LwE4e0PQMLiqPdojlhefn+HEwh2jjG+5
/ctL4wpVFr90X22UN5/xMD/36k21ZEyMVv0z9XTip3HiKzWnBCDuI3QIznkeOp+7
DzU65OV1r7gvYkNd5ksOiRHCgA30l7tX1MGi2QbAAHMdHh+GvpHvN772gcBzVMX3
QY6jfsHeyTpD7FSACiGsY9BRjPpuzfRPzoEUOs4RIwxRyDBKSDDSbFKSAnW79wAV
MbkYUdCLndM3/vXDdC85sXp3dEyEYWqs9uiug+YbZUEAwbbuhCDsBgr6M4qo+hFI
Zj5U+rwFGaiqrn+QwrjhESNR/W8Xj9fPSrbZuu52H7OGbNGkKqjXYFIoyEuckR0F
uifOPhYQ127XU0e+J5XMmYr1xa2i5dnQf/qV9Pd56fzTPB4HThVm7hFtf9a0cw2f
9iapMNBbzE5yafDSF+DwiEJsUqVrf0s/Fj8pgnW+vYGB2DJTWH+UGsgSYaJ/7m66
ws9+l8+aLDxe5pGNsCTE1fQoHMcutBefg8aul0tZrWPyIu8OIWaP+r/ajvmIzaLv
KoegQY0byXlrdwk+gT18FBNnuTqLBm3OlPtCTTYuat+ycmtv3EjDuCETUlVO3V06
q6YgfL+VsNSableWnN0xoQE9zBopeWZhOnyejBjo7zBoI8mzfjPQknlHigreUiFB
bYQVfUKNOefubmQcEe7XCpKBIRH4lRa1UVdjC+bTGxOUW3bA3TLZJNSTxUvEbntx
HVDH3HuXYagQtP8zddgNFeqlc1tHEaw0fQSm1GHdGiMrrcrL9M8cxxBkOXFHJFcR
bwz7KeiQRUlkt7ju7qdOcVLvrSxwjvgPU0WNHCJlggU9/zcEScA3RjqC6IgZ8AJo
XwJ/SdSQpzX0ZN9KuaoOAwzZmv0KWGrCRT9bCRn9lfVwf+yMWyxGySp+7Wgltdsa
WQ0UMA9FltD7qH2GoKmouMBcbVoHxjsIM8u1jErdyBiXuGWG42IwZxnMWRgsg8GE
m9sX9mxjIYd3qw7lbdMqBkg/x5TLy3VtzzY+MNElQsjTAHvS1lymdX+ebQpkIA6h
fk4FG3Bhh8zCyNxwZakbazZ/YwODFd9Tcr06NAydPPHVI9m5SZSEUgJeq74hqZxC
ezPPzengVxfSD7zKGYoxVOgD4OhsjPyTH0Wso9bEwsWQf+R8K0ISyHhjaFxzuU22
p2AkJ3DeX/Vf1DT0G86t4e5+bvjcTPb/OReb119oX/wG/bBzba1eOhzARNMJJ63P
nzVJlfHxzr0/CCawpLTzk/K1W5NcAR4OdZk9wGaIOVEo9/4o97f3ANRQ9gtQc3nV
OpRI6uYkFkHyjx4H3vTQiNmspiL44B8HACmljqMbMThy32LG6Uj1idzYRJlbLazq
G552pd5gD6HbJ7hrstFbZIP8k43Xe+76f5djclU44mGo9IweISGehTjpQZjBVfwF
cgECKTPiOut393HPECU9ptTnZIKCX1twx+h4z2AHSG3AoRX+swCYPtUMZtnZcK6r
4bqicF3ug8WxwXW0vCQyY+OjwLZlW6DBQj6rDOUCetazG3UucAsn8X5iv2T52rNE
vBRufjytTsbjbn2SzfeRKgvXqybtdT4IeyeLJcooeLUta60+YySEYhNzMnDCDUHm
jJR8mBVy+OqReefbiQZPugKQ/G1yeVDoX68O4kY1iRYxZBeGvTKfJgPYdk8Svusn
WBgl4X+SViGXHYmCr8Aoa/qE+Fu0NV2Pxp3J6Fd6lmWrha1VaGxHS6iKPgNAn4Wo
NKp5k4tP75+5y0UodRMNXav+G//rIBvOzFPfw58XtuXtuauc3NZJL2Sw3SERGzBV
MUKcW42QQuQnn1TLxEvQhTrvWgfv013xzcOmWkOUMt38BJmVSWsuO+u5T46avV79
Fy76rPvFf6eV4zf8fSZsgJHiZrRGE0cWCVJ6eaUmhNBn1uxcbMHZqpK08zDDwQvM
35boBbOTCnhQtYVsOdbSbH6OZpxGWfimO0M+Wx3DqolClDH3xFyVcJjzo/bA0FSm
21qqu0jztUU2PeR84BRnRPLn4iUAON/fGpoFu0g/latM9xbY2tRTZh/1seCdmpNl
xoycgnyZCgBhw67fK4fpV0GNpa3tIcgo12O5cMJZ2TqBrgl2ohrPFF9xs4y6ww1N
/cIWaZY+sZCbZEht56Dd/GoEmQ4kWiSJducwwJTVrBKep8U+pDKAP9R13kD/KxvQ
es5LGu7t4+fGUDc/pOpK0qgVfXTw28ZB7KNB5Wdy6ozcwZO+ySDzz0I4cqQwr3zS
lGq2V3Q9jCrALKyA6xPAdxW0OsJD8fEHqAdfefviC13b8QBj9RDu3GLddko/gR9y
QVrunR6OsoQJwDO66cC1P9x5JYWuYzKw/jk0ErSeMiBnXm5+5VYw/0Q626SDFyUT
D6AFneJeb4wCbBX60W3crG1Y6sUmbAzEGd6hhxYqQ8bPug7iUwKSMe5jy9IOugiQ
GvoVkrFlnE5UmnxqhoNpnOhV9NLnFQDE1pwN0BZ1rbUnCbw2tJQRDlIGPHDdTc+Q
JNG9hJZg+cIB86402uz6hch5aS6wGdf7aLiz4AO8e32QbS55TGlvfCgh0GjMiBGX
yvAshUNZ+v06/28xrqKunu3l7AwkuYx+QxSuDLeUaMRkuFV5Esbo9Y30rl4hb8tD
IGlAGS6Ax+kaqMt3cxZf3UPnQMY7naqQFRCNOOiycd3UYyZOEFERYxzOTuna12Bs
PSimj+162b1RUivGjsqN9mdlvWbOs0A6XIrhBwxPiAQmCpkK/rLPBqNAzIVFTMcS
ob/A2LnjarmNTIFqNDPi27iXRJmEh+YI8Cg5v1JPEXuAHfxiHziHeVZkNuxeuU+D
0EZ2adZY0Cp0b1QkoYIBF2dfvtbYpxmp+QqnGAVjJr5j9gVs6WE11Dcn+DEyU1/J
dPbsGg+A8FME3xp3cQNET9XhZLW0mkVevDf/PxBO2yUhth51AMrcJR62EfbguMim
ekeHPPs5iX6R2eopAGFZXEwu5cUAvmzA6Q9QU/Pq94dD4k0sIhGWCo6UizAwGfOQ
TRMlwkUFPNk+IxBp5m47lZH/Ey3qL12EMNfwOC+EuGlEzQ8Yd0kEhXf7DruvCjFJ
v6RQl2Rhf0Bpqol29E4jNz0eST1QbZNjJiJROU8RjG4QUdWTLt+WIn/Er9K41cEg
v6C/lP4a2kskmCc7wivixqpZO3y7fX1QVpzXD4yQQLjOmzfg4uN5UZ6K9yXZ3ptQ
RgWmkMpAMBU9Y1l2rZvvpOMoiAticoWnES4ftuZvnQdBvyrTL+IEmU5PtVdF1dmO
QlOqRcbtLiWPLzmf5RJDViMU83dbn2Wc2WFePPeWptkZTqYK7nL1mvx1L2AQqpkQ
SndVOHnA/sni0759wL2rcqGRbBPpc3sUrpqgiQ+5To9bPmvgZZBeJY1x0npviDSM
oXl/R9kZG3DN9yQ7BevAeDLvLhxFmr6w56kcXXFZNF9esXqiyu1CsHudtUgzryvP
xz7Uy78LR4rKPcNlKVJeiGSlLXEnYuA2V8hKkWPs8MqJGVMMJ5nFZAaSR4ix7yy2
0XwilWyu6zAPD1402mkQJ8lJrQWUz4+pdQ67b6LLooKTwWOHS9feu+bxcWOZaDn6
E7QvLDI4CD2GGdVavJzx7SrgWVFzWXiahnTA6y2FJtlho0LG/8ddNUUroz0Bi1pg
GtE+GevWjwST8690SBIPPw8cA8yOwHUo9AL+Kyg39n9h0CNS7hhZvhFbyoqtYTmq
ioClvmJDxwz1Vt+ktbObTy83Bc0OTHmWdTCkFpagBk6m75oeIjH9Ngq3iPCSWmN+
R3+vn1uD/FlmuGcU95t3Z/UCdIqK+BoP3cUzbdi1BRmlir++MsXtFrrPOR7oP0lm
Dsp+mE8ypPJ1o5lddtpTMjr2DWTRh3S3YDuL+3ZnP6xM/I9oVWiFVD1fo+n4t3r3
N3gVTVRfQTva4kTn4rMlg5XWscSSkr0Ws2hYTJ0NO+7TpHQmBAP5SQh+RsWaKUpR
5Ss0UBCWy7nW07WHpLa8lJQ0SurRQGQEO4gQno+uUlnmR0yrkBfcxFgGMafhusIM
O6d+hQY6XUp8npB2PWJDbdkd8AoyYzPsotcp5ND2kJRunvv1ac86bK2o8S6pJo0h
6OCLecvBUXpho3IFPKm/Ae3eakh64XAZxOG6J2kx9YAR+Qasq5dWrycumzs5nM9f
otAJDs21jtJw2oPv3gdNDOpz/pSqmbO+81Q+pMaQ4D2djdWNYhAdDEMd6iPVofrR
VGQJJhQPJXbh+Y8McPh4SfqX+XP6liPgVz9dXsibPsYHi4Y9LZxgrSYgFGfynDEU
gx+f66FFyElgqhvRsy6DZYhAM86zAAQmLQWcaq4CPXLL6Nrz3tR3Zvid0WiEtHyC
wn4rcGI7CdDTK6y2qjEdWcAMoH+eQsWEVSYO2Zj8NYAkJwHKvnbyq8on112GmjN/
vGVqk6JO/nQk6OBDwSJEBiQFZ3THhFGGnPPrNVG34yisraOIOR/aAuNb4mX+V9bv
yFAP50cV+x39WkGDt7J48r9tvzTqA26VrY+oDACyVIOoeQ3qSzqHSjxlHYptbBRe
2/YGBpn7VxrYfxw61JliBnsQDLs5hmWbddvNxSyexuNi9253xSd1Vt3d8G9lK0uv
etpkPXMmyyYPhvA6A0u8Olq2G/v7nJj/8dLpa/6TEBLPPDPgIx2mH8uT0a0wRBm4
VByUJnxCkeJgFRVNE/i4mKybbArZp8Sr0/EmzKeZa/CvErMNM9rExBEo6gPqDtT8
UNxcTNwOtWmer5xCSVC1Is7aHzebRD2CHhSooevTybhVmY1RCifcbVg7zUXUWa2G
PE3bi5N/25mXZnEClYcX3bdpkHm5McR5ihV30lnlh/bFCRGofawHsvNxEKUsE43g
FagbQrkcskGR9uTUhZES/4qncNJwBRgiQ5CqiVi4Ygqfj7bQVV1oThGx2gcMDQ86
eobY6Fy9+RNZsbVQQMvJkNsYoLpMyclVt1wOLmMN0pKlxjzy5kHHDQI01aGsd90z
qD2OJmfstvB8bJgtx/hG1I1McGxsDUd/50q+ttFDO1DrLQVOMLsV4MAzduuN09CH
Yzd+YuyyJLILZtfk5VqyRXA6V2iEFsJDUo6E6Pp/3COLr5g1RMh/ak26WhLs2y75
mwn4WBwjA9pLTXFyTyShfeGrK8SogUWaiiazmwq5ihIdOXqREgickbygAlxLr9ig
dblA4ONY0IbENeV7h8g3H+TZpLSxi+1yssVR9if3ZChgcXDjai1HDID79ot6MJuk
5sDP8MWfb3s0aHxC5062WKI4oUIFt81w85c/jtpWXGaWCNp9py2ac8bxWIuP+hBd
vH3LrPqCV01BFhVdNYckW2WilfjV2JSrVvJNQXCiYfIGyRxpsHlpKWl3a1MRI9fe
FWfXaIZdS4d26k02xLwmLlXkVg2h65vBzaNsOknmYcZ4M7cBQG3TSsIgs6tLTK36
wLFr5c4xJPiAJ8nRbF3nsZ97nHJ1ifJo8tQ9dCkC0BPyQDwGFP9yRc16ueeJx9OB
y3pFyUa7fcbZ/v5rzJv3i4f1DtPDZgIGmZzclDpKSSMnqElXplBOWjc1wfuANW9x
K4XzNKslOgMceWhpLFAUK3BRgf7OhTkVYEc6pj7dqpaAG4xS9+0JWv8/RQt1japX
LnE9dfQPCBwqRtX982qboURry3bVY92Ddp7g/1FGQ+WJp7jeGj5l2yhcFO1QVEy9
ZpvjBzujAk6Im0ruxR3axudF4lkyXuPZcUO9fgz02qj49E8rImBx0nCNdXLteQFv
Vfgxip5YzKGiwy1dRMpmSFnquC4VQNgGQ4AJZBxcz3JDAdTROKM9QvRoSd/iBdeF
0jh0HNSRNtcs9CrG2/5tsH34dWoCAxciZf5cagH1+0Uw7nfNnI8ODiK7BCGwTVQD
nHYbS85Wv/PWeShEGJ9VmMRwm7LkoisSSpodbnPqTRbpk68N2S/DisAhS0+AOPXf
ihlAWDGxVGnK8oqvqsKf03EqI0CadmgZHpB4BfZ+tU1hj6nOGfnrOjXMDAu+jDfn
uNVTmOi8VMEMtjiEna2Wf8BUUzGBOmKAbGZh/AXEwi5otlg4bLp5pHKbsFYdHD9m
jizYo1if4mtH78G6nWZoZ5NUo+EmteptWZ9jzqwDQh+k/keYKkUZ3nwoCaNr2JD8
W7ODHBgg/hvFYYOzIExE6El85Ui2Jdz59KzlwzrkL+XlB0RhdnsR2zceVk98Lifp
pzt1H2bCDv2nQd8O/PJMJ49Qy8Duf9H/ClxxSgIP2pNLY9p+xmcYpuDOUOVw+39X
fRsn3p/+Arzojk9En9p0p1ey6bokQhQhF6TFj2O1o098v93ArxxDXvJd9ehNF+wc
TqVxQcNY0BWX+hR1h40yENX/Wy7X/D1C+XKg9Kas+tyrq9auF+vYWspHR6wVTues
fzJoASpvkxlSN7wgVgGfEqYiqlgvJgDDNnAuq3MQVVjszwOhrkNIXW7wQVsfnmhS
cULVzMwh9Ic08wDWyIBZXx6ATPYtfmE1hrFThvUpSojygVfH5RA+ufWetw7AkTtG
rI3aK0cWgzWGNt7zaMjHKeGAyKs4CRuo4dXcu9RSuYFhfWzFqGEmKXg9At7QNV9T
AukoD738jGBSvZh6ZzBow0fcbKeiB56S9R40xG7X3CIfpfZDJwNV6JtG0AIS7dn8
9OoZp9VzU7SXoCOU/L6OZZPVhp9GJJB2qQmjr4CGzouCuE4Ft1Oa8XPeXI4FTPma
GlWDB4vBDyQ+UzuxHI5FhD+2Te3zhIrcIY7Qfr1MlT+q8a25SInuBHSeNRaWcWbH
DH4MaTCUeCt1mfD+lTtVJn0/CDw60qha/r6XNmwOMnTF4KlQ2Wg9YXcMHca2wIdZ
H6jIaZASPE/m0TFr6YYxkNKhpKwjZ/xFsdEQhC5o0l139DHQtVwGGvmP+56r4VdR
lRQJqIlfq1jWMUXIB62Va4XGYPH8LWcqNTlBJ7nDr2UiyHmH0QO/pKi+yQ1ZY9cq
Q8nC0pXIgpmh57g+JB0HMKKLaZU/LW3hGB/3SlsQivs/qvkt5qusrivd7pmd0My5
1zaZff3X99jwrSw7L98zhumP9IgHZy5L3gaezx/ZNmlC15+RXOPBL56GTpGwrcV2
fC3exasWxThKjrh/1cQ6JcKxMfknopPC9mEoDIYa0kYxnMMc0lSywCat1Y6gjtbd
O5AnMaiPz/7wNbDwazMAF/URzuKRORLDy3BEfCktAMKaoin2Z1/ubprUfdFD54Wy
9EhNFObVnKjOnu5CUFMgaps2HM6rpMMx8b5rZcF7pKNWQCKXyn2DOwBd1Ji26mXL
IMf75Ab1V6DSQZtUsxugMG1j+3Axzv0YKOPVTxY+Dq9j5sLtjfqEKvNYypkkqpEy
ugzyh1L1N4FGzzckW/q25/OVwvEQTyGhx8LKdTtcz8ywV+8kKvDyniZTX/up3L8V
2gNKzVfIuuEhpKg/p2rQRSWSZnBf99mElMPng5L/RWkGr0Ar/iDlEc0+TKenh98S
5I+gBGQlJzW7RY46dbAJzqS9+ne3BD+EnxKFc8dM/t1IIyGiw2FupjJVrX0rWFoA
OpwIE/4YTSdWjNSjolNibUST3M8muI+RXlArrU/nb2YbRUK8+ejWDF0v22wPRJ/C
Kxj1wjSgyuCxstpgTs0NO6an5SgPA7NGMjClmMAURTkprU588wGpbybfM0hLSvVu
7TySjRndfZ6W+Cn/NR2gD5s/uQeAXpyJq8ZHLY7xRWYGhhU+f1HFCejDL1MS3oWn
ZwYEUMvDyCr9vqzziQ7opiiaTUqGZk8t5kJvSnteJ32Akz/5wcmx8fZexqeZS35o
PEKVaPXS8+IvC/y4LX35VGHp3NznlMRWt+6Keb5OOYVIVHkqDCsjIe+G9qP/ZUTA
eWMLRk1TT6Yw1wVdx6vBjixaat+NCsRwnIXh2xdWIXIc4s2do7gJg69It2HIDqzy
qPlaDarNbobfKHnt9SsiSJp0KxzySiRN7C4WfQp42lMhlzo96gQ9BP2kZp7txdJc
aj1qSW5HT5XX/zVTQKQwlSMOlOXKxvd543GNBjdqhKx8XK0ZDwpDJzNwcdgVx282
LNccvpk599jsExJhyk0YnrW3fo2ioU9ROsMsAhrd4d+1dK1+zUz0h2QiSKu4nCBB
UcKwOEi86GzYpowhcLu3qCwBgAudLUEDywFw8hf7tXvIpd9kayq6cyQiP3cxcgDj
W+ZmoJWAzOwrHqVffsxcfSCOfmt7/+tqoPKFLcoLyHYidx8CMiNyD34bsfQBBNVS
CrZhgZDZHZRRL1uMWGqIi/OpGoLqoDBMNE4HfAlWVusAI7jByfIDUCOMzQcBk8Xx
0sgR3OFWT1S8MmoyBRepM/cUvaH6gmI4mPg90w+PDxp6gHQQ0QwM1440abGS5epJ
FAArvmnr6WpJ9J88pss2HwZtyDCL9G+TgxmDGAWxtEwxeIJnM5v/LcGBBZpiHcr6
Q7TCamocJsbiwWktF0YJxHSzXS9cWS/gwtbc4k+WdwpUryZjtCd1SYEaxjTCSYYZ
jXbuPrU4Z71nyelmsWfCyiHcZdxZOpD3vUO0/C945RokQcFKE/YLrBXoj4qxmuvN
FclDXc/iBMIF6c/Vl4fc+14eOPS3Yi2Y/m07LUODC8+e5K+1s0Xm//xMi0cH81Zp
J1MFP3/ar0ShtIDmgA+hwoBT4N7tPy7Nuv7hK8V4LDsBz8trTMDAEP/6aKDkE0kP
3WKn6zkMtF77PZhEUbXkfKGpdHkVb90tVj5sbJYirtILjgovlZWSlj36w/dCxElc
TzK/N/C85o3bLTPFFNAUsYdmaeuLG3XM7EpsI9esuJuzUis0q42IxmZSxCHV4HXA
IGrvq2q1rCaTSo7aG1w21ynqutBi0Sv/mYR3+U0xFjUsgDxc59npvavPlBWKukZI
C7b+9i56dySTFM9+EcG/pl7alS1Oz4/gGZpEF7cE/voby1Kz0UElU2rAaipahkwX
Wde+iOGWPCPKMjMbpwLghem3CNHosv6QZoTWpP4FVB2X2B3xipTIR9aTktA8bIFt
ACMWVTdq9Ad4ylzMnDgGDwwXBQ4V3PUJ666TgrI2uuXcq/VlsSQGVFhwoLizKX8I
hr6z96vcnR3Aj4rMXo20cel+TRDRQP/rfp/JXJ9ugdYeeZnMGENsoZEeWOQNHU2T
ym5/giZSyF+wiIU7bi5zO6HaxBj/Fa9iDChdqrMmsnUff2XAagYqgjY04BUY1Ol0
TyruNPI82vjpaDU0gUCjplLkArSHixe3swWaJ/jx665s3QzSnNxW7KAzt02Rpa6J
Lif4wHnJT3ZpYX/wMRTBSZDIxKMd96IecAAIWZ7Okcvmj4mIhYPM8z0FM0E8EQde
liYdqvsKa3h9srKQY+FIxee3Lw8Awm+u4o80OUeBA4I27HXPyhGHwSbKipvllx/9
E+sFKl2Q2o9cpmU2zqqnyEogrNQ0pfBIrVOQ7BW67t8yjisCcKu0MoOChBoxp1xx
O5mApfS+JYdyZcO4f3sZhIoWeW55Yk/YaOh6Fcd11C6hLnxoN899A/HO8q2avnn6
grso7TMjkz0oOOSxcHejB7Gejy7Ahd6QN6Bh8N7q1OhGLWoSnSJMu1LUraCyGlMz
D2+Vs7yDKKa57yk758oAo9ZJcTSRGWQzCOn9E4f0pz47MwkbjCNY+y3dBwADxukE
W5vJgQ6SRQ720UjJENn2EeCeiGfLOq4AvLsxr5cqmjHhj8ADcJkGaGgL9uM9xlIn
YN2c6Y/uYZnkRrp4s6s17MJa3IL3/BK2KjW8jey2eVzLDhcMOrCG1T+n8BVBf/yr
AQgPGc3uks+gWYB29BUXjHOsghT1SSY8kSqC7Btnz7Wiof7N9XO5i2GqoRLot1Zk
Yn8PZ4Bt6y8lI6KcTZVOCdcDZjA57lrkTX/lwbHHNYlqCG0V4RqXrxHYxaIiDnWa
W/Z551hr0k6LRyRfOW6s+k81uFX4E0l4RdCQ0sdlxgIjLWHn7UkqgI5RQTalZbNO
DY2PtbTkAC3RpGqgzmDcRRLsxmo9M/DaUZiP8oGJKreFgrb7UhqTJasAUIF687Mb
MJNTwzDMKr0Zca/zdcB4jy4izYhEMljizhAvjEekWMQMoemIgXhdmmX6itqr/vVl
9WPUFBjj9ol7Wvey4QpNX4AYi6zxTRD0XDMcgeOA+5nlzjZc0jbqkqRb2Uv7v1ae
DLl2FSVj7JwqBbsGoYYGp08t3e2FiEBvYbQSIEERSgokPA7BPD3DUekHWNTtG5Tz
ZlNBUeHXlSOfysAXgrF0wg+iHedSNj7asG1KTKDb3ao1Dwx5g+k3g6yjcvYFug7/
BGRJy/WMcWAJJfookI1nAqsj/HIWgGeqXFAi5cYMDDZMCKEV0SKqM8EvH+3M94Na
enJpMLakO5NFnGauR8sb7xMYKQEWVRmq08y05MDiE6jfliaxHKa+UO0hD3zmBf9o
zZHzSMmHeUBLpLubNBN1IcwW/6HB5ktdnkRMLJ+4HMkBc5+p2emJijOuV+vSl7e0
IM4H7zxTyTqEbGxrOxDDwTMu+oOZvkX4LzhHhCDAV8yQy8L+GEAerfZDcDXqoAg1
wbtkSyXwcNJ79TvPzeWUW8Of1rGJ/YiPY6C+Y2jzSw+yuS+mYNlNrxaWduTFCmiX
5rFq2Bds2xaZsAeUebeOAe5tfVT8/IS4csYUvQvVmXS1WMuIIzOL8nx7NYsLswGG
YQJTHTXhy1LGLrAZeDsd0FoVagEGlyqmM4AoeQbwfZKCr4ElxQflv/Vgi9BTXdsq
y6qeKDScn8pZuDRnk6q+j/y7rp2e9CHcU3O7VBf5hyo9HKpXaJJBR64AyO0QXoX+
vkdr8eCFUxkICVJoexC53Gb26RITWyp45dLEzaNmtcls3XNkQ//hylgoHzU2aT1t
EJrbdYnt8GTkbuh6zbyv7+rga0AYlLhSmQ9CztA2fiHOLGeVnpJFCHrvDHrEdMZ4
9rksl+j292jVhq4eVvSTdlNYjAAxfw/rl9O7sNRlKmiL53pgMK629OOxlkEB5iE0
XrUGtg8NOOa5tQsz5l5AYTXBU3SeVc/ZXRy2TytQnAR0ip9zILuSPX47kYndnvig
oeEPntBfZMaPe2mwJW4VLrmdghiAIYrjZSDyrqI1t0MpLeMJZobx1QtF+XqHS3Pb
C/3+IlhNX1eE+NpLjBpEJp9iz6OtuZPoAuYEyMJmumpCg9241oPeuJifhkXCXfAN
SpkjjYTRqsGGazmXbvOHAmt1xmRdXVJ7ZJJNXXw0wtnkcmJOHBZiDBQ76LZfLG7l
kOOylwLn/43HjmiU31CA2+essb/UiW0bsCQuebSAaFP7qsUKowUI29FE81u/f+Pb
zAFHOu4yzNBywIUVxh0WMPPCxeCZYKCQtiodVEmK5F5roWMyQUoeEjB/kPKJQJPH
5v3y6cirb0HohFO3t4thJyz4TkDbNIB75rsLYpPiUj3KjBNvb0rmFrUFFvYgLOny
ym93Q8g1U9nEgGiJZrNz1gAc8HVOPf31YJRBQ9UVwjJy7mbn7sgCl+CqvqJWhifM
sCYsMGjpYr7zB4hyYfI6Fi6zfT37LPgHOCmxwEht0CpR2++aSBrMLqluVYZAFjPG
jEjGo3XC2oh6BvT7FXNTbs4tIQx+dJW7au7UnVMc9ay+TP7bJxRJTRmRCSzrykoq
1b1b7sqnhUpU7Nm0KeaCYS1/aygCage9H7IYc/hLfH2Z48sz9GaMPm0v5EuHx6St
8xT8QAs3HHEY1QwCocAe4JKGQEsG0IawtmPUE9nmlhjYKgxYlGOCJsk2sCHWOkMQ
iAvO/5dpp4EZjVuoSLIfUMQECEJH/3fJWuBNZ/7DhrVoCy+eM7RDONuBIbTuOiaW
FcoW+/XG/ObmiEbixLbK6d7RYC9joBsttIFHMdBca5kAUBaBNa42lN/s0UIkr9Cu
wuagI+ORCuOaJaJ9HU8OnVLuznwK38e+2N0MZQHya31oCgDWM3iWA8q6SCJxm16m
2K9xKOFrnPl5z0JkruLEyk7x+WWtYFx5e0FwrlUsDbxdoB2IOdNncvphvKuDqUMa
DMW9SGwImL5xW5JAmDJ+CXX1PTm2LL+YMgw9Utu+7asEm5mHNX2Ca/8Qj20pbgdw
DQcw4spr6Qle6uMeKCOcreaVaV0jXFZv1gxE07+4xelRusP0ZY9Q7FoS3uJ1vVDy
s3jOF0kMzTBLwoaJBln07ohuSrh3vNZF8yDh3H+KXeI1pXTI6YOqqIaMlDmfahn+
9cxX+rlP4KB5GleGR+ti0m6dzL/g913TmXOd3zLJCfYxSaqEt7n9NcSvgJsNtiZH
UnlDhK6Yb7j817SS9Fa55vFdaNmq5HWzNCKsYDCnzznwnM+Wmr0jAsijESSQEYFN
AJcj7UmYvj41STajCuM506tbTrWNsZa8Ox7uf+7Hxc58Aih4aH7XsoGnc+L0i8qf
lUlwBDeXU13aBx1d2YlJbnuiRpUBVzx2M2JLYgvMTqiTTG4Espebeh922rqzYw0G
u6ZYA83rSgFstBb5cAIZmSolgidbZvoAACZ412eew2IadXSAVe7bUb+OPR82ju0/
gzmcf3ZhIzC9TRuSQe4ff+50Yk3co/sWr/xxtSxiqzFyoOTUJXWPOXVHVN3DTuZ0
ILGEUr5DB0295o3RB4dOcwhlT3QRKpARYuLIL1K8sVs6WthOeFsWY7zThHO7iTHA
lShUmCsIw26BFLmgOBJtrPF0fB9nrd641WkhGJ9PA/KSo/Rg+ZOQ0c61HRhc4PTa
yzJ/tcBgD9uE6NHA8eXqsGgRkhmYNnsxbr20vVua05P8ZZnvhy9agkRnZTG2ZJYV
GzfsCum0uGPxeZev0fE57vZYDeUlJD+3B4yH3g7Fs6rRIIHsc5LVttpGkWdJuo59
Nzxaby2XDwQFbt/9OCRJynw9fvss/UIYOIaj6npaCnYPTfNRJpq9qSjfldN4UFC9
0w/7qHEG7YvAU6RWwDMe17NAmU2gZutDYwVdXQuCpwN4Owk2cet1jeawz7gOxIY3
L1Qd9BlAczjLLdgJxf9SL0gz/BYk39FLEMMOe4sq4h6oPJNYvgtqBhWbygxzMiKh
A1MqLLPvNirOqFlhs/DoJr1jNOQsRZD8/VVbRykbEtnhZXeuSxd9F03mG4kMrOGt
FKqzmJnb0UHQnBgwC1F+zsSXR/lZ/g1AJnQH4pAQZ/lSZCljTR/P3MN2tUxxuP7I
PSHdQoyCEyOhr3vChuk9JhJhDGh4kBvJ3pKMPWKUfwXaBUNYIHLq+zM7oZ61+ByM
a41XUPjRVCrZB42n4iK5Fee+WaVLfOv6fuLLFDcTCF7SRDcJQVOGTs8Z/S/LsMxO
BN7MIb3sN5QdULtLH7N8exhFw0GV1MpHwSJeF8Emnh+5Ht0f0ue3xUXRh68p8UQE
mcJDcdRvEr23BJeUgybujjV0kV6NJrtRLgeTg9iShO/hKgCMh/6+QPMUdSE3SNkr
lem9PlA1qmNuc6002AH9NdSvzV1gOmmes8/wsDzxasVLxDkbXRs2/wq9pRX6Aebb
oc0DmhozHUSQymcykLx5mcBUte+wqqfmWJQ7Bic1yY48r4pBX0VHXAuXBw7Iyu5c
3HbRaVJ0Mcxv9i/fjxAy9G68Cn5W1vDvCTo0c8dJrQmh61WC+uuAicZ27APeYrFz
TCWG2gQ+qFL5eMvnLVOMWoeF1qiLdYX3p+Ng+TDsFAglNpJ1PcIJb24C3mjnwkhP
enE+ZQf/D61uZott1/1QvdU8kA8mrg+58F8eg3u0ECdzLiBCX9yQN9yGzmnYM5+I
QU/eYO/4TpvqYa5Uq86hTCPTofr3zuqjlYcIM6Q5bgePlOrrEkWBiW+txYDagru8
5H/3Et3wqDIJrgez/GK7dCH84wekd2UOrIBrnL/20SRRy9CeNY4PVSAkVnNO+9JJ
qwilYBUT/0tQkiiORlTU9PLJswtkLz9JmXlO6Qo2RCjnpb1M3HacZC6OMUcEgSoR
1AoVnFLFgXGYq+FhsMZ6wWrB85TCYJA1QxiyWL0ZvnveP2gHSFZw6wKuNYTEGtcG
dJ8NQ0GTx0CkGQodlpXRmeRNuEzYFfHuUCZMrCdEkfUw9/uFpldMkW2yt1r56MAW
RXX71s6ji3Eq0mLD9CDkWNQERuVWchiQ0yUBeWYlsCVN8AznUasy4N+nblt+Vrt9
uq2pC7Iot3h1bzPfGB0OB9M4tetesDeshBawVrnc7FKgyKqkOZv5je94dEHW8RkI
Gab94MxZkL/dNlCwhkq7WLVA9u7EmjPh5D2zFmj+cgJp9MvYOcAKYnbpOOlGvdP3
lHZwgrTKVLUrT9BvXobAjt3htwzoaUrIpbGkR0YI8sqo/oYci0x1yYJLboTKWrU4
HzAJbSl8V+FL4Pw6d2xMi4h0hXSbPNeskHnSkqHS7zStClPerdaGRum3yC88SPhK
C5BM8eJtzynO+con0AoQZ3WFGjAJisw4HdbeqhD8emlMsYngEE9E8wlYcO7t/cL8
w4gmbY0XuhCEMT+gONW+zo6HALxILzfJBPTqmZxh7762DeM+Fp94MmuO6JC6HrRe
T1S155avqMRsQHpHTuq/cffZc7Dc3QeiPq41rzPTkx4K27yobssR9vJeFQSx9mew
4WYh0ZXf4HdkDixhw/FWaSagOLScXxcaUa0lX6g2plKCw3++UwrO804LZnzVKemd
Wb758p3qJtPwRCmoVSsBOxKgbAC4TEkGcN3Drt+o1fWMYY0Z96e5FPNBQu0sMoo4
xL3szvwJoJ7ZUpvWzwC/m3XJvx/NDM9xYGeMdESK4EUQKtMT54fFqTZ77F/qoby1
3TbN6+Yjh1ZD3gHIsKWaGiUMydJDldgQxwoTpQ1X8p3pnIwSEep5fPJJzKvnd+W5
2khC/OKvjSKyEr5PgQ4XSkygPvde2D8wUDMBrH22N7vlr7DtpwW/84l4oxCuhYOR
//04k4cxwSlV6Ojhqzf8r4XNus17r9eXgOo9bUVmwJa/RxEdEzyETgGWbQ9diYHx
L/wpeM6CYY8+CJGkoBqgkb6FKQMUh1kCQzHIgHTULPkjU+t8BF89nZhu4j3gTgyv
+704peCNFXPgadhiB4i5+MEDZSjhDzebo7FM0lXhLvPCGrMvF8iSeLh1zBfb3w8p
eo3ClvoX9MSUyDzhWPX5OMvIKst2884Ghnr5F3NVbpbsmgkchYV3keKqgEieLUzw
dF4UmY0TY3Jyfr2fVeoNZPM3ylKXWY8ERvxVb3Z5mkz4ayt6Z4/l8X1TJwPOixYC
+4tUWohzgq5CT1TBfEZhpdcvxQFHS9tRXb7h56LBS8Vnl/PKgBBGMV/6rGlIi+u/
djMsWQeesNJZ4UEglFaIiY68qYBEhPA3LjlMPp1oNTmpjjHLlH5WPuxdZ9nNaXLO
wOZ9EJ0q/Gsyb5TSl3ZgGxg5RHDIpllTEg7DXPSd8+UoX9l3dDiFmvJI+v+IsgKG
YWtSeMV7rce1zgM21K0mUP67dDayf5zbz+EaJKu1PbTAHORq0dkL7lZCUr2WCUEd
CUmObFxyOi5rmsDqjuZkR70bA28QMT2GukvpMRn6deMh1+zQU6yShLHu2cBpxy2h
jYYuj1dfHo5c0vynzIUmwT+0DYKcJK79DqgKeUwx1hAW3zGG+bCKjxM9f4B0aS1Z
FEXvHOGx+xsnEJXZYNAipaRcNGMidcmC4CTe9uiqmFxG+bxqbcICKnH2ZZKBFij7
DP9oF9fRs56/vkAraYw4AIsMYBwf16ov5sQapgDX4v3N1lkZcdIAPtcVGqTc+rDI
7tiNAFch3VcBSeZFvbRqbX8Qqnl0lZpO0SKLp1giwYJ7Ms02EEW3E4Dm2xElzPzf
gAFwrINybvnyxJkiz8bj8FczllBJrn8r0Wxit+2CsufPXWZlauiVYs68Y1vKK3HR
Oenv4543tP4t0hGjMZiXumB7Ap75vsjR3otOTRVt6Ih5Fhqf+VPAE+0khXs0mj3c
1TmQ1gIjxgieULPS54ewNYeq9MYgFci4FjIDPLlpbNBU5rv5BxC07fZB+56ZHuOt
i6ASCkgtI8B2L4W1dvYOqQPGfboHXGruS4UAQB4iBuvQclg9UroY7fa1s6V08JCK
zYLDSgtDxMojZ/dIymzlWL9ON7tJlaC72BDNmmdxcxV9ScNsCj7wM5UvGH7sro1I
ry3xhI7uk9oHPC7uyVcS0fiXg0Q7EWZbHjIP7D//ZDOamB3jwsnvE49FVMOMFvGG
h6wloSSSX/iPUbFTt9ZrwugzfEawfT+8MUNNnKOvNB3uVDa7/pszCHiQB0k/bTHe
kcWcEnFKLjvbfAlUzY+F2f3wBcCz+yu94o5PNYOJjt/XguDL0kcgO0GHzWCNwJbK
jTCjZbSfohq2bNwAF01cIHY0V92WTJMRetU2XmPQRVFpCHdb8sNA9wsjOyJFq7Ce
mIO2NR+GgHNEr3ljuAIbDtfvq3xKKwRqL1Pc05KhBuuo0DQ6bPSViBMIAx7P0elj
ULbSk6akE5zMtQi6Oi4mR2DRUfyE6bimifEpkiI/Z0wVNz4lrG1jVBYwCXHOXQ2a
0B+L0j2cEQAFHV+4Y8HRP+8ZPatv5BzFg2dK3KSEBi6o42M/fJN5RNv+zPIHh8R9
ZjDTCZPk+FTL6SpQJoURNPProZ2A3tUQYcpcfv8N3QZR53PMQNxg2FdJP7pFrTz9
QOGm2I2QQalAdJAE8xK1heZK9eriQYtPZ5swosW2MeV4WP9WDqPnVh9wxyfWWZm2
++VpJ+/kvpyHBbdveVHDWHkUy6fMBkxGO1ImIuuO6NKK9gHu+qAEyQcZcDttpJiQ
MMZb5B7hqhU5hHskpt4nkjZOdERc0B/wucpSScwqsBLXc1AncDACuSFyK08o5MX/
tpfN9BLbWdVWWdwnXzytVgDii1ItKrJtwZYNsZymkURdL27sKIUu0j3yEt0BdtoY
O+Qi2a+wAAbbz7LkArMns41BRZuH7bl4C/ePi0691YaEeQbVs50kTminXIgiZnji
45d+SsfOeFfMI7gImpLOPsSazdoLTS97UT/SZz2g31XIzUwb3A0tjdz0vchHSkEW
cynZcaGIGJKUhUAT/thAg26GQf2+OJ6/nvh9pakVpZ9wwxkvnZTG+L8agEcswjJ1
cVVoS3+Tub119aNFVnKO9zI9k2CdS/GTYm1DBS2vA563cMGQL3WMr+CLLwd5GExE
2Apzd0FAUnJOt1cyJUt/fqIoAbb0ruHqUsQ5TE7htSXqAakBh5rqDyuP/X8GDx/R
NoGpzlOfZh5+NBHS6+ALUQ98ODjWWVJh+jeEVgjFbWxSLZskpTvzLUff8Amsc0bz
tO0LDwk4fK8hA3NfLl1Nlf9U32+lMRijLNMinpFmgaOuGvbgi+XckYDGPa9x4m8r
uu06SeD2bAoK1OFEXvGiBOndVj3emzM+FHbfNUzXvx/fzuCI+XSNsTJcm8tHtpof
kqGuf2JQ0Wh6WoxxW0SXDxbswqKn2LyT6EouP19Z9vlS5gZy6riUQhpalMO5g6KN
U+ZxOQUeIEQ6eRrmHQT/cZXaHgLoVDMXoFCj4eyrOxf6H7qLbVv6E3cn2DumDsVf
GcPN0DIJ5iXs37sgcmahrfJqSpueSumwTOCBZwxA+33+yfLK3+SEiDtZRp/DHiFh
CDXjeb8ZtZK53u5Dj6PmYhuG7dEMWb1E8jEmOiLBgTvTA3aJkehh3vc1txfzZLla
m8VEQ+YphAJD7whthoAo1RQW5xDGf+95w1cVy7dM+egU97+b7bMrvKruKtUZ84r0
wgl+MJqF9r1KTXJvpzNJqbzatgT/XQhGwBUR4eUKUKpwqgg+3CWzpSVguvkKrNC5
aqV2JhL3RbMyKNXFXoQJWCFRFZj2fbbAb0VkUOVtM9oQTT9z6ALHfk0rSvrax7ee
+tm1QRRevIB6ub1WNAqtyneTBxrYF31xWNAeVTLS80c8cWjnr9KB83CdsIs+x1wP
1T/T4maKGYnqr6DyQgBFBVrf6JOcmumvTy/LF2dqijyr9docJx841EhznBrjZinX
KNwRRBLTIa6HVV7MOwrut+PibZ5bLE4X4VkT/Qt30yy72okNHuBReA4nxuwckYAg
WpGWJI2/fCcE09RD09xcW++RWECFqQ9qK00a5mLEJjG3nLHpEbPkOUD9fKQGGePJ
44OAPFNx1nj0IlX4xZbO9VfjfVtyJcUo53eMFsGjGWLl3QnRjaDxexfXpNrK6h/7
5Xe2fAjQH5JtdY1pMT7myVcJGWWeZOmuY+JBAj1SPWItmE28sZ2tZiH2qF9S9U2z
cMWQFY+eg3xYEo/wq5wnACwgRuim+H/peAKccOK+DQmLG8YIXBq/0kcrl4cC4AA+
G82QoiX3g1a+PsRnZEYLHEwDoYEpNjLVvmgTxJf+XkFtJPvctG1TP9sCWw8Sxa30
HX8KCXwMDDz9OW94MqX4ux+XRDiXy/EtjLd3TxHX8tryKcS9SrPSqqK7fGmoayX4
uWq4dD/lXgAk6zQ5QchFLUscVqhGpLAhfc2sRetR65jMZJ+LHMe00/E2vJ4whQLS
PMboFnsMXjzGNbL4H1uVS2PTxSDChQM9Ois3Ite/6MnRb8hFlV5jXl4tATJzdb48
ry/jnyCtSpR6C5YknUFi9TH0BowkXV/TNU7muBqYPEIZy48Hp98a8FqXlhF4l0cP
z3l/bUkf62PA1+chgecFiOq2oaWbFGBBdbfsZtFl1YIA9tkVCbMy83zGwbFi6i4k
26Lwmp8YbRSvWc52bSQh8Lt0Ny2LLTnTvgh/tSx2Z88CG3CeYwBXJL/apAqmp0Kh
HCYWIBUiHtLiGVRyrIRkhgGR45huJimKPkBDaoEi3UIqcKSQz+mj2ddjOVwzbVyn
ZG90LJ+iHQobKDZqUIE+m/9GFRi0ZKOBgMIFosZuMXznmcFXXP2YKNcItOG2bg+p
dLmP5e5+bptGlEt/w24cYNcJVRZFWnGZSUre9m/Xw51IbNMynbf/HgcDfYP+b19s
Tg13h0AgfJeSquL1NoSKRwoLvVFz4w6p4ZjHsdhSKgUkrYiMeGfIre3Uh01Lyru/
PnzChdtDcAJvYv7Dr394AzI3Q+lwSqyB1XEnnWWcZQ8vSZpq8LBYhIcdnHGl1k8q
u0DT1n5DB94SGi7lp9efcmcjXrMZtWS+vJtbOdbBtBN8wAQZgQ7BkiYuRw/POsvz
h8mSeFNTaEXdnRmd63G6L9V9dZt8YiKCvh/QDlMsY8k+5jsgoek0bUE0KxDSeOOo
sNOKlPgSJt8mw80ZNHAnjw1oh374oGduZjIsFGPemEMTRX1ifTz2Dxc962ONPPin
QZkqezq0N6jxVdz67hcQ1PgpbJsVjcvNXDCE7v2AAT8VxDR1fw1fRz5aOzQE67rn
Qa5JCb+gE+OkxcJlXmWY6C2N8VCkY1u/EaMAy86dhcWEUMcvymRvEE0lOs/3LTzf
qBTa6Oq6Wr93H0kSg3kG/FlmYwxumqS8mtiW1fiP/96XmC8cedT88bFZooBQKtAp
F2eDOHYaniGpn8quEO4DEp6ddztbrHV2McHfYZT/QZaSPbyHe2+cOT3PZy5BMBtz
BoPiv4nvTR94tPbbOIDA9Lks7aZxafOsiMrwiBUtrf1DOtMz+fHjFHrJLC3F99ku
ZtQYIIpjj4olpo5zoGXu5BSO3wYYqjSE1ASxYKFciW9akdWrTjXAGHNnUOY6Wxck
LVbQcQaKOzrS/j8gL82VGBt1ixWwoGfcnw9MJAeiJ9U04TXiKg8c3rHa5CQXZiF2
h9s5ocSeSNMGnM5tHKFO4Ez/X9z0In6kmmBSz8eZ3zVFhtZsz89TSlvJ8Mvq0zAo
Wf6+le78mjK0HSSORNeC3AdWiFwn1ekSWtXwE2OVZtzUV3Wk6JKP2kmUW0owRWnU
F8nCs9v7uBKChMPLaQGcqMxhuhUj+FFNLmns4ori1Gq2fvkk17Ptn8/ntR2jMz3r
7iqioY5SNWD5QdoleHfwHBLKKiQ7NgctSW94s0lGuTB4oYbyvgaz5UXyrf+ey76p
VnDKE1LN7l59sAFqKuCp8JLgoD2hBhfmq3H3l85ep1Qo2hF1zVnwIQ8nL6953SVb
1UH4SgQMk9eESj9GuD9iyscXCYSDfaXW6fIwhEbM5KYqBDHsqXY84hgON54xLYuO
EuQV9G+pVqIefyPep4/4Te7zULFg6u/U11upEl5LBDIqGyglR8znbg1jBkCuPYhK
sTLUKYuDJc0aWYsMhgdE+D8xRikgQzAbQsjJ4uKO6SSBjWimmx0rtgoxCjNzXa1c
WA6vEKWaAiqXHNfHqRNDL8lwqoBqcMJ9ucBS01c1BIte3Mfd/I9JQU3KYOj0rEbt
P/OrlsjoOzFp7NoMuTbNu6AFduiXaZFQyWKAj9jBZHhGyTD8TDXoPhEjMDRfNMyi
GXMATI7EcNiFluUlq3d/Wl7/1hD5nYnwlvVyjgzmV7q7WKh676CbcnzeAu6fJdmp
0CPE4XkYTpn6duuoHotgh9SYz+pb1+5jVvdPZfnRv0BUp4f+TbsvKu7zxSca+KbA
bIfZ8UOyg12LjHzvk/00IJAqwSkcvNpJ8ZfDB+nnlmUAKlwj9S585ig17hHlKvej
47STgxijQ4NHQ1yET8hor/9FPSovQPCKx0Tm7z2mdsPXM7gRjaEiLcozPfjh9D1d
Qe0oe84sh+JOCXByvvFneuypr7R+V27SzaBPI+mSAHzi+1wk+IX70feAdOQh7GiK
xMZgXecrJ5TdRpwhwvp/fDnbLTNXiiEvTS9MyrE0nVqpBJQ3PNHaCMCbI30M7+70
yYZ1WjUdfwLR9wSnqCKWIkQz/mwxFd76+h/VJJ2f0VcbjQr/NIXFdU+aM1iiSTay
vJALwCAKhfSVJlQ57jznqz34y9IGwJz01qNPTmXJaNlE0vWl2fZ9xjk2OrbVDi/8
poz+1UQjbcHAfQRLw0p2oc1A3AZo2Yo/S5gwUjUBMRIWcxgilJLA+dCLi0Z+vQ6k
Z0pfiPBX/Dc3VaT52EXHMFlj9nRVa4bovkXgvps1ZD4VO6BCVHTgXWOoYVBO8+uz
r4l4jX/S9Q74aU4NPa9KtbqAO4WUluW5gpBP1TEwoedB0PdOldhr+pwUDqxHLOzh
miZybNQj/F9IAVGY+6wnG3nXSt4UPYzoQjqsFTSxvG8mQJROWnP8NDVIz7k03tOv
CPcjL8/WA9pGTxI1PJPUYBZ9JHKzlj1feTEKXZgMUxANlG2Eg12ZofClzYih5xpM
d4YJ9SPxp7vH8glNznuoFk4h7KAlbOQjbTgb78R5tOM8iiGyQ3PE4gZgxRAgr2BM
OucXsAPGC746QDc/e7G+oKv02NgLGCZTdPIgcumFNJLrNX30vO23TbJoixLJzO/t
Z/CI28dLbpHnMPMQ07CAA8SVkgLmfj46WxUXBmaC7B7JcQGKqY6VtBfXlxmglEiW
NJ1wgsLO3zd9o1ks3Yvd4EeLsNQyMaaP8r2X9R2hSSKIj+FcH6aQKPTc+huxGqf8
n9gHDzRUiCZB6SXxDp1D1qanfb2DZ/k8m4ZJOYxa1NoC5wG047T7+U+K1TTEy7p8
gsLYGTpFd0E1Cy9Zh6+KDbbG5M42xb/wpYSlvZy6HBroLMkHE/pnEgh5xSOrlj6H
7l0xtqOFpILmcGlIIymL3HoylGzwTO2YwuGumolt8daheQB3IguZeNaj/4u/8j0P
k8fLVWfqDBoUZ84iU+3TbeNGJIOwW2M1ZW+I2xkehiPUQp2XTdbgcM7VZVdPMh7t
pCukA+8Fmei1oKgqcBZ3bt2iaAjnBnPlbaBZjc5trXfKhyCHshMaBpc36lptVdvM
daOaACUhja6+/032+C0dvu1piiVC05nM34gE4csPAe/dW2dpuQg0BSZ8SSuj/yYz
7YbmbkaZ/uCvOnR2NcxbeCziwUiYrGxwbmExymbWj8k9MYOuxJSQxR30fTfImxRw
Vf40NhaaKl+QXBUCxmziAT8aXTmxG4bXNU1Cdnzl+j+SmI3ZkjZE+807KYulRnDk
pRkZQ8+fIluryi/J7kNFYbsbFob1l/99F8VFHV1PAefXcSE8f+5Qpftf73oQHg32
2zIwHPQZeabOHz1wXZPi9EEXQQY5Bs0XzMWmrNpR0dO0lM+onf8RqoyVE5JTAfG7
bDvRIX3VxnEjhtLvHc2/WB/rG2LlIQ38v1ACyTaN1zVhA08CVFodUMkiF9KLQOEo
3alv3CxvD5WSXFQAJkqQKQ4IJtGpqlgDfkmVIGJIZ1Ps06zcsz/pKtuyGRos9mvb
Y7mpIgLxttO9ctVyEFacRNPQ+1Kuv4lVsIJu93Ps4yozd3wsSrkW5asRm50vvv7r
zgOqMj3eZnkEFilTj2lgZ846xso6nL0lwOzluOC0r3XMmAUSs8H/mS7ueJqiWaeF
15TtEU6XwJhUm2dcJ5HWOQxeufcBlAEx44VHjmMgE1IJ2Dj/2VOEM733ZfdNweRX
gPdOXM4Z4gUDMhsi0DpWxZU/ggojnnB4XkHqrdObpo+zmrw1YsNVeAk73v4D6/E9
omMS22TDDav3ZKVbMdlrUQ+Z26qAO/qgHuLYk3mNpMKB3mbo2katXLnlBt6Tzube
odB7AJXRTuwQbdJGhUGQ/Gc7H0sGajyxcrqlC6hTMzuC7MN9NMnTBqCqeZKFXaoY
w9IYq6zGyvhrgPPHLzw5I8k9xb8ypEBP3xLTqHiQmy2o44ffaoebNZhig1x/Jg+r
OpwqTnrKjD7ujsdJWOCJ9XvyLWWB3RWbWn6yYGkxYPTiYsrQgL+BKJD+ZfBPNX1Z
YQeIHV7SqJNa/e40Q9azUN/Y4f3ffyxTgmJt1/RBKn9rg0jejfhpB8rNFmfMDT+L
wdOR3PN7RwPtmZDbj1y5kvBQhE0PxlLE9v6WN4ku2H3a4OlHVz67mkcPVSDT1f4o
u3Sw/rIxifLVWIIye6BuhKKjfSVdqowYd4FmS3M/g1jQs6ZkrHJMxusrFOkc4vkG
H/GnZBbUyzzBZaMeBLdFHNlhm2DChFIL0K2u0bWIzrtIAvd7CQ4ZV1itVGOYXR8d
HUx2z/ZPJEVnAHn3F+fsnk60+O6wQ9e9Q1+71lBh4mzPSkhlFAKxUPUb1+UpQbaG
1BYyCNHCALxyoYzbwIXEFWG8u1wXQpEcVaVAuHEf9sLuMQaW8PRbuaRYgyyrCda6
Of33yQ0+3smr6XX2YbcQHbcqS6/McyIWmRMzCu66PLLBYsjy2dAxh+rGTXGTR6CW
D89yn0zMis+Mdo5001VuPWR57w6pHZpP589lPfnPeiZm0CuXetLtGeZMHfTSBKA8
ejdVBJR7qxp1Kc6Ti6XWd3HLmmyPQCpPLjhHo1Dflx6oA/9sMF94cS1sohS5Hupk
EOmQRnURcxs+OifC6hargwUmPUUz6Hq/bWa4ILaw9hDD51ilJQBSCIQa/y3eRXN4
rHznr0lkGKpguCxROVNYNCUwalYCIOuv3GM92C3TLgrVcc1rdLAQ1jP2k/KV/7Z5
gcRMcltK9tbadTZz1WN1gGmO9vYbv2Nk+uIcscwi1G17YvueIVAoe9GZ6WWk7Sym
rHEQ2sCAe+etwnEZc5kIXEcCKMXHjPqlQqRLMMVjAnJ1v9z3sDzp1If5aDkU3FTZ
fHsoGv9U4IvXHfXExCgzJQC4vR+f09fbMSLhGbP4xIpmzzp/TMyxuPOAqla3RM4D
tzzLGaFHTGrlxM3EX1qs90LwaM4JaJMxpADj8EwjV9i8aiQiVPQR5ahRGUXNeUgS
luK6yhR+nMuNBP/CHaLNQ/mpxV85tyVdhigjy9TPCdOtx4V6Oof54lGlsOQmvcxu
x4FbhZhTiQuYcoXXuJsLzWLB+JyrN6/SQlMM/hE0v5yaGPaJp+kFLknVSqY+NUly
lQ+39YSfb7Is2PG3Duzgg8fNTeREZoqEOS86+dZI4ekl15Db6SKQ6I3DixyqCUcq
avpqjy+h51FDazAcQQmX18lgc4/AAjlKkRbxCKLgZdBgln9WJwURA6RsFW73RBhi
rlw96PMbaXOJjURgs/nw46lNNl4QyHmTsX9jBVRL5fm0t7NSc4Ufgj7JNEurk0Y0
L0LrGGeqOeMA6Of6s3XQHt+eHSHWUkfb9/fbsAAMDuo8w6EoFRetOUv/cYzqWeZ5
s2XOaqjWKdZKyvM+8i77CeuPVGNDSgn5o4fuRqBGT2SA2RuD990UZTy/DL3govSL
3xZR9f+QQy7BaT8oIfkmjsW0uKfeRS4rDVUYugkHt50PreOZJK56S0tsCilbus89
UKTcwBP0r+8tffGdVuFvXTno1gdc2d+gBIm2KjQTCueyTJV3UNeaoKTIMMWEAx3v
HErAoU19dU24qXUFmig9/V9nrVNz6O6X+ruZLhw3bynZSUpnYKVS8MHVwKSy45Eb
gFW2GjQKUpEqa5AtIDPwJKUhMzTzuwgqr9YaeT2CeNHiPCJtRYS384/67lp2k8bR
znXfXW0em38BWurF+sbap55ib1Y9/ws/xEJBu5N9d2oCS8X9Ff+hUDJLA8ISQJ1U
t8XNboELyz9b6uS/hVjHcHiXsKJSIwt/g7dG9CtQZAtpGC8yBxzlUUV7d582HrLB
dLQzgvXhtSigjPKI2qv0YGHj9ykViwOutkidbq+pDMFDwjZ5VUMv8ILuk10l+Pyb
Bf+p2zRKqoojjjCg6kt4zalE8gFuRsgWJhdAmqoGnVj3IckSdyjmLVawzn0SzxBi
lPeYD/+sABIlxljCLES09BVBhLNH8LDNzAWEYdE5WGtsJ/+ZTAdNapAT5X+0cAty
W9if/xLXBp0KasdtrcyRTqutgu72KdHxrkyJXpPU3wrwzhQV+5fXcQSLohMymG4Y
bGCUfuQYRlivNSFVe6385Zsla6ip8XZ2yFswmCaQhffVdfnRwLS3wL4iQQmwH+LC
aI8Zqs1+m+1EYS5aWsBjlcEJVpPAOG1PSe5W+mJ5C2spF0OvwQSMm6FXd1n6AEhx
9PgSLYAQDOdoAcDB0BUOcygUs4FedRh+zjrlVM12dB+GeMJcYyJKve0+uK+Unby7
jNMpiyY16GTSaM7DJUJt40c5XL0FrDnPIcM6ZmkX4dsiJ5HkY+r9zmAs4KD7G3Jo
Gl8s53uAj6TqFrA6bx5shI7YSsxg4riS6ktQ8WZGoK+nH7MxjwgqlY1OQTYwwKp4
ZCrbGGwIAntkVDLtlObsaRlux+FqR/mIm+dXloHDH0bMrsIGSnGbKbckF/PWrK8y
GZfqSmu5jV5ex24DF1s8/r5i1p4/XXizkr+HROZoBvF+1cMMLyfAvJaTma+tMWlv
VTCsBLmSXcvWXvA/uvaiL//8b0SLbkrb4uYsKxaxHsgFo7Dfp6nAq8+4nB+gYcq7
JW5+3DmI1D/3M5XdbNWbD3bld/kIflcTUXJ9xzMSoy1yDQW7DuB5DFFo919vIQlf
BmkdaVyCcDU7mPA2WW49SdIDqTwkj2RtdE/+ZBFLEs3qrhAv+XDZJmyhKh6q2UKQ
yHd7ce4asJ8y5qE6WlsL3PdPdwLk+3ukH9viNQu7k8NObxdqqcBAFi87FXmadO6g
F3CiCa3WIoY9LoVLi/XivyfNgZlpBOfuis5NeFN8H1B9TX4+/gOgsH72HI47jKBE
UT6sTWpeOJxgNNvSgUY4H1vj4vc0H9az2xzeI+iduySveQeUo7xBScbFIG135lIv
BaVBFwJDGMU5gFOaJZFXxuAG1VNVFN00z2ugljan8Kmevg1gzJShBOXp4CPDdal0
PQM0rNXvnG6E9eHgxcwSS8Bee26VkVnCjJ6GmlDd002HMvD5Y1oKwcpeVvR8mKii
y1JJtTXcU6pCVfgRy2ARZH/IPvCyTCdJgzBasJ+zP9InhrkJJmlqlsSQEOi10qha
37Epg+qsnHqMKlsPzTUESVYZL0XdVLk+JbJsyyvvuqbsHgijst3ia43b4PvQViuG
wO0XxSk6jzxTrPVB5oc1AY2n2sAZ4L0FlnZ8bqM6DuPBAepx/Ay6Lgfd79uzqI4p
GMZmAt4j+kdp4zalU7mckvsKCUzduME+qfnNWoBuPM++bwoOBqoUg4dudthyjv8i
ddRSbHoGJkVfrKUVLEC8QoNYFrff8PzCa3YwoOqLihnVgPrfyVOwluWB0/cF9DSz
2pH/Q2jRnzrU+U/oZAayRdlovyzHOBZ/yyzUU+RPzmEDho7dOlxQYRvYz8fZw0RF
GILYsyaIBzbR6C8UT6/NJCZuz+AWEktD+7/OrbTs/EGRNqYAfO4s3O6BT90YsK+h
ozPFxIe8mxbnzf87N9LilL0A0cFM1VkJ/3E3cfG/Kws8h8jHO8IX89v1YejBS6xp
CfbJ12nSh4tAYVTumX6maTnH611YXdZWJ6XmJWeAwWHE0D4ArzzHG7Seeka/HRNy
8/0uVT1TUtLtF0aQ+X8mE2RnQ/aZNETyrwsy/u1FTYsbGgmW66+oYPNFqIrI0AUT
OV80xn+Zfh4mi8h9ib6S2RDqV6rjLqBh3ZmPFKIDhYg4g7HOn88XR6dwXw4SX87q
HRVT2xWKR4WJLguGNhHvkX2eh+fWt2SmgKzw31NfDJ7YsDMwje2UtMT5kyddeQ05
3gLvsMAalU+Vg5CJ9DVWHa3GidA23ZTG/4yXUFSqE2Q0xXYcwb8eLut6K9lyV/Rx
OmQH0XBggWlk2WUhSjGZVHrCFw7xHIwEzHO5cT1jcVlfmtX/zOjQIxxlJLTc3Jda
qnTTiFGlwLhhE2AK7oUImR3rECrxIwyLipkHuzc1kyddIULSQBtEPONU+GLbCXaR
1APuzvfovHyImmVdgLSiX3Q2BHTsxuoHcZ5kUH9HAjDtcPwEhSabGu1oSHa50V1R
CSohapCPS15es4Uqgm2kYUkvH71hH5A/5VqPcsrlB/dGa5kmpb6XUBQ49OFGlde1
mHa0uNozhSKqjtvQPovgGAlO6znoR6/kC3gNzbhC36Ycyd+yP7ZxeGxB4KAG20eV
nZab9o0wF9tzVb7EyJsoD7CnJessJGFhAPix3NSFUiixhNi/uwKupo7O77lKXkCE
gXGENNXRnUBlIpkNF+g6kbTwnFjL5wasi3/04DG5+MfyvKN4wSBN3GVZn2mPNJr0
g5nY9vYcNC287PC3SlNJ4YcwuEHU+CajR7Y9sn6EWEWDUO9T+KlSZlonNh8eTu0S
qLDnbGvoxynDBJE+lL2V/kbhOyFJxcZpk9I+8VQa751gMJyL8FUsU0573HQd5uYm
XvgyaVhSe88ImjQMb7y0NodPPlJzn8s+oPQhhqZPOMU2FqgQDkta5Az6pP7rkUOe
r7uXDiQJaTzupw/QQV5VEw==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
c0T7t+h2p2oJ/a7MZVDCbrRz0NKRiSZ1I4kLtQ0XZVMQoFRhNPeyYx9Uz276V+Sl
Uf7BUOsdC0P6bH8Zrg8aFVLF8PTiMFVNOUa6b1Au04YID0sS/axLcIuxx2K98ltG
+3reLfY8wFm5MpemuMgbjzXP0Pd3OZiCf83QB68SoXPuLKwvAFcd0DuUeG/D0oro
cQSbvT6uaMYzUy8uZCvWgcjnfsYUorLt4fc3LaD6z1XyGknIJVml9PDjw+nYL7+f
heKl7okO8Bh0j/MvyAcNiA9egXXA9G4E3K3aswAQyi/ahNEC0H6tqy0+vE8d9S8U
YB6ISVUpGiDos8DmSOtpAQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2016 )
`pragma protect data_block
hR11EAyICavsFx3jdajUhlQaGtDnrP4aiCAbWJU4lhDXHYNQOrwVHVF1UL8hVGOH
UNT3/Iz/5w3F37CJFF08fG0z4aSL94PNYjxGxwZV3v8/o4L3UZ3pGPGTy35aJwTp
pAEKwyorhxZKMcv+DCfoRDPvq0wWZqMrCmYIbd4y1HJao3ZrTS1mgeZt2ppPeTAm
HW03PagZ6A4/7RfdY0tFGbyoPkMxmhMQ2ytJV65OeS2yaPLKI+qvAyOOE1MCS8GV
2GbN7I07s3TFO6BwCJMi1acddivytGzNxuLEgCsWeFd1aKKkHN7D4f8tK8n3Yobv
EElb66MFfRm+2xhqY9m2pmi2qipGqq7Fxt9G+ps3aBA4rveBTVfYOjBGDub6Qghg
MoH8Zsl/VnQpnoemjj9kDQjgPwU+rRmWrHNd8Ha5MKltweOHbAx+gyw8Elip2Oci
xPbbPUDuOy/M0H+kghSztlmmXBPFh4b66mrt5HXkx99Dwk2fiMpKQ9HMVI9/G7Vg
UYH17Z2DaQT7Bhcg8ZtJyO7a+Yk2ZMF7ZbcZdXa2grTV8Jbr34j0ufpFaeFecy5z
MnpuQm7pRr+X8S8aN0y9P750sO7q5AoTe543L4PcnuDrfcavQpdTeOMwTt3weMhT
q74rxRebcS3NmPD0lQhDUtX4Zrwpti+OIK3TVLFlJuHf+nfbFr6DaeKs4aXsLhOT
2NmqC22b6LipTqbaO3ZI4xZJayz5Ed8A7gHvLaRzAGK87fygbLRYn4xGYBZCzsXp
qt0Be7/qrWALVV+2HGHpyq6D7uCdOtV8zhrCqFbR7N96Paw1J/evRpa95MClvYoN
xrJ5wt7iBjo95eeEJFgv3jua1lXy1grBhmHQ3r49YifcbI/DXXo622DtYoPxvWva
Hj9Gk/AA7ogK+fPlTjToPjiBKPIJHPEd+3FiG8m6T7+JuTFqmVy3VUbjYbQ4BSit
PfVU52jGLwW/wbGAIO1I3wGbZ0zQOOS7qWuPBxiJNdeKzvG86KRlGMiqWS6tXl62
V6kfUmfG6h6T1vUsIa4HnEnU/XHpLCf+75lAGlTc4xo2MdyO8pb5tw3RpxabiH3k
BrYheZwQN64yfiGygch6gSJ6Z9ooN38xtYvtuVEq+JBNqRxgG5gl9X9RNubKt2V0
y/Rim8Tf8/0g9PmsqA/9j8k10r6HdhZTNHklhGPN/pEpSlo3iwHTLfuV/DvNiNQQ
wHKY/NWgTIRp1r+EcGnQc0vwLbDZZAC+aCQPv1U6uWBfpKW+3IHOfc0uJWdlgL2D
ZLunnbFKkqvECO5wInDrLCphp+5ji9wg6vuhtDhjdseAdDLLpMKoIl49C2h7QBxF
bJRR1HxgP6u4eiwawjGSMF+KXEYx6bIJJqNqW9ahgjZ3LwdeWzkIvp++8r78X1+b
Z1FK74fu12aMP0lxhPeuaO33GP+UMOi2GfFybiMvu8zzzqdkOtVhh1wMikjH1UeO
SaEfhmOGe6Oy2iv/c0RoCuzegFg5krSWuENZX3dggVdfkMnP4C7YZsm/SkFbuh03
zNgOxHCbyZMR31tZAamam2xnmdwbsuGk6wyp6uhbd465K3ClU6jLHOs1zSUH5XMH
5w3gdAJRlMB5ctUXVl4QVdqwq0lmXds4/zFdEDsWZDZaCxMA8Cu9arFH9/cA1e8Z
xuZ4jsvHyg3BNUVWw6g0LVi23pZYSN5LlhSM0AvyljlGssOwXR0219dTOxE0tT0I
hAWKYwAWfKiYGoeRRT+DprdDj/dvQN2i3v5I73inPohJOah5G6BrjvJ8GHHUnMY6
8pkT7palG/pbbGtLSEHBh3utfkfEhYz/80Y62WatSawNz290GIewv4TJ0ziafosr
pGX01Bff6Il2888C2ViMwQ703KS2iInZZzjQQZHqFqWDBgsbagspsSg23fvVrzkU
txACmHnMOUOjnV68CQh+d2VUoSE9fV6e5sXu4Gt19ekBhNGuO0gkYcbWBNmkXjHx
/0PGHNR1cCbDnsYq0BRNWIL1eZBfBuurFqCSWEGdz56JCtABDFj9Sdz7B84emAsU
iD56i/GtmUnicD17gjOi6fINMKY9Uh6Y30tjfq6xH3cTyg4QW5nwpnwTwSmYV0uH
n57Z8VXVSiw0aZ62yZm6kWEhnLnJFaIZtGBFSXRWVv4+vYgrQ6skxi2qJVOKbv7H
WQjhzkSNoWrzcXyIQbrQgrjjOjaGQelDrRzV0qjvJzHa8DsGlMIFcHpw2MYcpWuP
2f2azQTmep8qqoYROaNNuNDelZ2djcCvtoiBRcwh0kWjA8WlwI8VXw00mejXd21g
Zb3Os5/zQjyHWNYN2KG61gV96X6YlVqkQTcyFDGP/fZV87iqZVBWJAZNmDS16hFz
+5Bf9+zspKIcvfG0FTWAYm/0DT3S3YzthrYVxy83/MW7XBBu8qlxtJg/r6bb2SA1
XOSi1HMAlrtcyvBAh4jMhccm2RFgFySsmMzm3SVvNxh/0VYTGMpT9nEDdecOe1nZ
2F6xaGhE9qx3K8HCd6iWnWqQ+Okgvsb/VhZZ1CygermLTuAvThFXpeySzsIs+YsO
oHJ1c0jn2Ccsq2Ax4+6cX2vKKY6I9OrqsFJd5eiD1Xs/DEtH6NWn4O15Q1WLMifp
7M6/EoH5g68sL1KT0DezqORfCCDWD7PqGGXVftaX4xeLM3t5FfT0TSZLW19Na+pB
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
n5KJ2mXoemm1nR/nvLacdxpeEKDpu3tkeTMY4s8sfYApAOL9RoQrMh7GDTFeinfO
bkTsjvjEy5Go+T97ZsI5+roKEXTjH0jOZzJhIPGxWQtpyXR9xfyjV5qopMu0ySUw
NSFScc83b30k6YXz6X0Ec1Z0kBmqlyIQ+CJ+mamO5WAgQSs07kKhytOaMGIJL9Hk
NcpjamFShpOCq6C17c+mPixEguA3HEsw5vW9QfhRdfTQZlTq2h8GB4IewYu4ie9D
UWjI+jJP1GwS3AUDdo+E7GlAdY2wcQycHrpH8xHgQqZeKx7fuOBVre5Om15gGl9V
No4PhPAoJTkO3TDLg3WX3Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10976 )
`pragma protect data_block
Hxddhy+BGdmIDkoBV+s7WWnQ3JuW4SelUEG0r2951V1eTpJcDiUNT4aQMJnUrSG0
Ru2e2euZFYMZLqp7LZNX8krL5pjiH8AL2mS5aCt3cQM2H9KMgRKLMQJJz5ApZZZK
5yZb0sObR0cnutByGIs7j/3u1giSaKRkD0FivyzowrZyynuzCofovPsskzj/plOg
s2VEGbaeB2qcH+EANoqbvKgsbs3xjv22O+3ARwLbiJyhscxJp6oEMBaMtrLUgwtz
jSvYYgLsGCszClDp7a/EgnFnHJVJz0EmHtzHiEtGM/QOU8NrhWFUAT8X4Eg53nQ9
ctxQzgRgsQeALYCEphNG22ckZoFk7uEdufxGihUfJZIE6xChSbLa+UD89XsD/VMZ
did826WxDKd4eIN0GbsBgH66TpVV9WEjOSHzcJdN25vHMtKhhn/8kWyad6QA6qDD
dO2ChPzhUOVceIhBIjx/08Yn13BM9nD+CsM3zwA6eGghOIVnNfs3GPzqqfSUG81t
aOQbPQ3XjZ4ldqqxbHrFA1TL2yMRYZ6N+eSv/5LK5lli0J76EjZXdbg4CBJwFtJd
WO71sUs9rKr34cUVZqUAJkT+MtGYFLW+cHMqTqC9xSVFC9JrSL/A0lYTcw6ZTRab
OBs32m/5yhX4ug0X4U+W4IxZ5X7o7AyO1bs70zBe076QWXxCFDL9yxGw+qqM6NS7
3+aqIkIi38dUzbuB58lTYJ86MPSOL9xwhDVFLUARUBuFs0p6Er3QaTGtbiJ8EmiG
DNP556JrDOzl2wIzgEN5xIWiqfYsDbji7/FRbcRo68SmqfYl6YnwLXdL1GSUNMC9
UBGnomuQm3AFNpJgvNxgR2SxY75DAnaCHv4KwkHC3ad3M45rmOjujPO1Gv7houla
IIyuzHcm+y2FqYpU+f0JIGaN5dQ7rNgT/WClrnp8IQ3WKJiCd+JXBR3Nhbwkfiqv
PBHuGQxwFrIdMMMlQc8taqfWLGkNI9y5Vpg1wWgEPyD0kPQk+homZV2jUwjMoll3
LnytETv108v/iHiRdlnph5+objyuUovOLfckCGQNbsEOXmjkxJAwIN+MwlMcrXTm
rFZxWe9OZnKUO7Iz0YwB3T7kSNd3sNVGaqqcIVJnHdmW9ffLWDL5aLB45ndpbi3W
ctq+MRJnrMVAU4v8y0UTub0qRSkSH8QxFpzOX1aHqg5mU2W6E3WSxpRg2WpydJLG
FmMy5x8YbyToCM1zP7LzIXOou5DsfEHd45orZRpuChtjeZCv1/A67vrMH7DRp+Rf
9ll+hyVoO6cVHLcnnoZye1Xc0yrJvrPev7UQOc6XIY72UgR2Ikc5qQ0Wsa8tRL41
QU/Lc1mRPxz60qbbVglrH1aT34d2Q10l4JyG5yhjqFxSOguxZg40TTu++pzNchst
JUElCr2RCrMRyQW2Rp8Afsd32MswXog/4kClGOZnAHqqsfEkcHJb/ZGnEv3o70jT
3IhZKT17wVUuQ8VNGD6tQId3pOjppZh8Zr6BSP76DKSHfc37TBEwgUxrzJTiQjRv
DDLXD1AD/Ll6WmLEU50dM0syGScHCZT4Bgwu4xDFrOHZbtHpVGPqyDQgCXim4YLz
T47x1FffTIPILKKWGxKsoGwj7Hn7sJ6rkB30MR38diXs2p58XIpH7FJ72lQNiyfa
SIS5zLPFdLNfmk5wRHsn/JOyJVGux1WXS0Fj9plWsocqY13QgrYEHMgXYiWudL7B
EBbXa1NastbRFn3V9QobT04KLxBvjmuvZW92MjCiRk0AGQNeS7Pva88npXTX70mu
sdGQRIf5cb5TjqmFTfAgf89AcNVMbcT9fvWW/DpNANCk8ucnu/hhH4R+0MEWxy4m
lUG9/ryO4DqQY95H0ZemheP0+6ULfTa0zT4e0HTBqyvgn9oJ3faxldEJzamYDEEz
4EaRMHJeknYsPCvx0xUDLTRqGxYVFJ15vJ14FyZvCrvV5Olx6X8Ek1DB7oqJDy3V
kCSB2LpZ0KePLm3oW1vK1LNai8Nu0jZUPkYF5qMWEpDzwMzN42AhxlsfUKZL+PYv
2DpmW8eK8topTZa44fC2Es5JpBdVpG7l+FAtTjJ4vztUodt6n60XCedxF0sMRD+X
dtT+Brw20oJ6w/GUC17o7g+IaYUm19qmocKXy4v4toqbhmc6Rck/oBqRzxUnvcNC
CmJAB9CImxhz6LHAum9omYn7Yt4+FgnaucFNt/b5VaPZ3kMOLqANMCEgUaJgkSYc
h74Z65WPoZ779NEW7YECN+ZyumwQw1SM7LU+paG2yj8/r2AC57gWRk2gFvS9SwZM
2JHT5mtt9KIMbJAiCyqm9bMIXWQHfPLhpvkNeTzCwRrXIgf7M8FhSjxhrWpnpUE/
IG1q01IVGUhSWcpu7Si/DkMs+zDYkyj1r80i6IRoyldeRXgQ4g1Tc4rA2kGjaq81
x0JRX7BKZY5Zb45ESfmLgzMQI5BpouN3mdiZmMrZrHWuU1ZZcWtRmzzjMvMXpKRY
qeeHbR6B71eKKpO/pld+AjeY39rAi4QAdVJmOf/B5NlSpEmaHcGsgvugRzbm6I6A
2tYnnB51yPF4++mWKdVS8RvsAB4922CtNYn41dEgfCWHHbuXe3xnHLUhDd6iysPw
qmVcAZBFMg0uYzRKGMUAPKwoLXKppkRxNysLXSrj/tv43m2RGMOO3PtXQd+2n+Q0
x/0ysJsruKlC4VrZ2nCPkDvrHpUIYpNLYcpAMDXLzQcO8kSHGrd1iYnj5RRRf/Y2
l4LM0W7FPMA1R+jtsrFPXQ+7Oa/si0v3gU9EDTKHpHV57B95ebyG2YRpPVJzrKjF
YVjMV/RBPAGQKe5XQn726Pur5rbxB8Qj64lhmzvTyuLA7gGFyGe0wOQIm0awD+p8
4C/19N1rKr4LImAGIwsDAuMY74QrI9F+dSuT0LkMO+9hWdHVPvzfoxUm6lND9tvX
S/NciT91EF2Y1+6rJz4R0og1O/e9x7KhFMAA06Pewwg5iF9EtYy9LICh3niCBAWY
xyx34WF6vQinBrw+92S15mTCjDeIjb95ZG5Ogo7bieNlhTy6TbrJM1vsR1rWi7R9
Q9is7Dh0cZHM2aVFrbhwHxG9FzrvsKHJ67Ym1gnesRVasY8jUDu01QY+BsJnuC/J
TjOjrWYqdroHIDQSfWVhD4M6z0kTSzPO6hgoyS1nDZsfpjCCb1HUuRzr2FElPAwG
f/bVwF5nQ2me91f6tCBDc1Dg0kuCfArvskVclQeb1YojAdTFAc8jaHr6FIFB3XX9
och22XJsgHBTS9hGoTyljlmGZEDXEgikyG7AeYIgSzycTQne41LvPQlVtrfaSYvv
HfOEAfvg28QBwNoZUJTsL+fBc99ReMxPlm7YYh/R/LJgKEccXjOaQYUpv0HaSAqq
WWKRxHxzdeuS38taVyYxXw3MEsEddvGnDGsz8ObqWZUIu4g2UAuRuG/dRYUrJZFt
8pjMV3x3GrH6sHPitd5znpMquFuiQwtzicayNbc8UNa/ForjikVTW3Si46oxtThe
3cUDFvGTy1trr/TmQaabY4j3JzHCE8W69eCpLi5D+xSasdV9ZwQG7qCq23RjjenX
TcK6ZBNgAeICjnKhrQuJdpW4KV8ujUZaoLsox9nkA+ZVQYUfWzAFzNBjPzfnk8Qz
IAHaJQwFGaYaYlC2YUkGOtgFUZ8veKaslO/vRyrPrv4SYBor2SlULVa6dXz7BPON
94E0IFBS2LA2BH/wIwdpHiAVKXfKU1MpsqwKX6sIHyAFRSrvP4Ehdo5IKk4DLe3w
Ct9PF0rmKlu2UP8Lt9iOxa5Z+660HYG7y+SvLiDMKVnBl6q2WGbOLoe6ndsVzTdL
KhuKMtE8rrlCSIicQdYEMhGS+8OhCBJ9pX9hKy8fvUgAUCPnTbC6GJcMjVuh6ScG
wQHYqx1TqsUNTlfPbeMfhjowkiQxnWeD6k06jFPM+BSnWkZkD1Dv4/JUk+tbsVO/
m1c6EVI5kuFdgsV1c7HPnxTbi+UMbvO2mWMIkAJl+SP/JvJUqIhGniKsRpVGu6mm
4htAo+AbVlAujDllnpU+BB5JX1paJ4KZIOqGExWEAgmLQlk7MJ1R3py/OkqjaxEw
Aomyn0iGiOL5G5wosNsvaE24WRo31kHBun8FjDpkn1JN9sduItvWZ+0wCL0cl0nf
9tdfT6NHE7AG3KecQGtcJW8akf8kELCcGFGjA1sMjws9u2R3J++uBqNqf70b2kVE
JiNBXKaI6xhQNE6Rl/LS9xRdgpOK1fanWAUODmxuCCBn7xO3qGxL8nbiezj5k+BP
yADSZ0+qu58PhTO93KvPQ3DcJvLUqiqnubKBqpSZ/fML0v0bkzmmpc1flDifgZT/
4rcC7Q+9e01w2MPI+Sapj04yD3vvuxuym8XAXqi9YwnekZcQ2lEP6PJA1Cc6pVBf
fc0RF8xcojUkDzct3Pu0OmBAmDUULP4LSVHpitMr4+vfqF3wNbpXHXmxDvzTGnD3
0dX52cn4e2R69dWOLwevn2ZYRXVGrs0txvPGp1XarR46jzYiu7GiiF40+jTkxrZK
ST5ikIZpR+GyhhRMyJwVq6QnhrqDkUM8hrH0WkrmkLZ924EbWptvPZJa+vQIGv3Z
LaVNVgJXsCgbyUk8VySZV+VqQZcEu6L4rayNyHo7oBZF/2UlgGNgREIeLOb0QTqt
fkSYc9rYRYqKcQSNLIqVT16joOtA+eSKbsUfRyqX1OoBukzAQuepiUUpb2aPcbjv
2CSGlxa7YyBpb4wIncisu6v7gGzT2kYjM2NMblUnz8nDnXfsDvy26GdTfzy5Yxgq
btkMXv9ln27qMg0lStmInBPq4rkv6LGSkYrqoM3sBk9klD5YKKDSLIkoDJ+BQ9H6
NqgF4sQWEG0/lx8jcJV053d01f+xBni4ehRoz2ulHyLww8d5drm3qGoy/LpSaUfJ
tzDNHfxr0uT3XqRaMmfp2M7KMMl3o22WYuPqA/XVRSys5+abRvY0A4F2l3qWyXkl
Rgco1xlrrx9c3fJzXui5KfJsLTziAuyvPIHBzJfrLFZorq1w9eLCcBSb/W+gkUOM
9Xq5UtfH94a2w95tw0/PYARcO56SEXRMH8pAZSrt2FEYE7M6+8cnM/IhP47H8Prz
qzW9x6hO7igmEpWuuqH26Wyq/oHNhjD1+4CLxYQ+ixn+ncwX/p0U62gah8YqD08n
TMx1+P6aaTqADIPJjoYASPM8qZNhYL0SfapnOQTkEzTSzfGPx5CQkQy/ug60l5UY
SbqoWff03tEasgfd/5uG+1xyvZMJSOOyVMmE7J/k7lSTVS5KJm+UCama6x72q8zj
S5jsZPAbOELvn/JgE4V1VnfE1KBdStt/qKSW2R83YIqignxqH8zs08LUo7nx42MG
60r8fRkuBe5cjyL7syhAZaLKAox4QoguDPQV532XBFHTwUiG2CFJ/ZTSKew4ZOTz
o3HtMLgI4DiSpiTyCMIgigXcNxVZRhwsNutc/FF5jxieizCJYlGEt3PqkvdUbHZq
ROmZmRain9gbrC3TcXTaq3VGebrmgEHkzVzvMOd6yv+QhVbZVvg3hZuxcHmQxfk0
jmAQT//gbMYw+rJ7amG3k9h3xh/moUbjK6HFKMMDRUDfV3EhHqthioHiZO5RVdqP
wviS+FaIrtyZvL2pEqHUVJ6nfsFzkZa4Otw508GDZ8njiugsNOvgVtORB1WR3vF3
OVyFkri+BtUlyJN3rvU71O6ZH1s2ERB+X0Vcin8J/aMXAWF6XTr3jmzllZf4vKgs
BORE8FvEIPDLBJ56NAXZIsq+MkZwAUhYt3cl0Yo1e4re1WEamBt+sQ8qgzkJcIFb
cWRbEwCFTjsX7HC81xIpzrkRLg+vTqnE84iQ8nzLNLYkmXTN6QIKD6WB5pvYWf8c
2UhFmv/EQp+ra1WZYQ9o6pYNH4w9UXJY5AOOZZeEhvtKRW02Po0k0dUeMeSb7y1F
vEstB28EHUInCaXtWfKk8/4XrHrRsimOOejbSw9uvcDlD2wBBplvCa45K9aqOBZm
PaptGWDECJOMuGSD0RsSIM3eWMXTlmY7f1zGtXdEAbNSIHT9xNxX732JcTmW/2iK
ugv5lYltrxd7+lHKf1CbZ7WR0Kji8/FuzEWdjvRWWzrIzaF/pu6+CntUjytCmiXA
gvlEchIqSF+GQFQEeZJ7Jf4MAmHgpjCeUmy2CBR3tONG+WPBTRIxCk2D3GissO4P
OYRQom4pq3vZ4JsUZcrFeYK34MxaH9sibdDYZthLeTIKg2WDBQNy0oCpUHTZf4Dq
zdM06YRDTlx3WcSv8Vfjn37hc91wkz5QoEMaB9BV+6sf0xA4NcM+bn/BOaooEIAK
si+CJPiL2Rtp9RQkYJy2F4ogHsiLiGUfQ0Y3tGgxzYA1YjDJAb6Jq/jORXDtrHFG
/OrxrV5IPEgXHBHzuACkXCDSCHC5/XcCLf4wOvOxvMIrPDkaRTW/Sli7T/XQA1AS
YQw6L6qX74ZGxAN/SgYvkzc6L9QkaFTE6dEmrhwEW//qcEpzjvwL1WCUTK/AKNq8
H3MAbRdnCx4OWwgLN1Io31r5MpPG5sMrWymHZ0yVbrXf//ZC7Pk6ovHdXhxqxvci
e74sFTWipYdTVOWyQromIAPYZtFrFTBzN+8EewW+RxlAgHO2nKBanT5rM5POaM7r
bGqAwejMDy1sxXMicTTBgdmiuxpvHnCSkzZ7pUxn9Hj7FTTO1rY1R6+bO8otbgy/
WAdYMSgZV4RZyl1BOXdW/LyIsNLyU6DsOhHE8d/4WZJC1+dyOVXd9N9jvOwcI3Rf
rCiQ0XvaCa5gNhlFX3jtunq0E5GXiBTNlpBfKQ8GqbQtzJKh5L7TETaKtMEKRCLP
zA8YNvkPxJcKalH4c7P5vkFmiUuMWTAztluIVqOgVVSTTbPc4nPL5Czr65xyzIxj
JZbE5d3pugEQ6N9a7hRyUKE2sO498Wekkn10/Bbk60FP4qyfjL4pR5mfcKSVcW6s
8xiFp8eS8GcWSJrAI4gjsiff0ho1O57utiMPOzVnmJC/4yTJ7TOEQ8ZQmdbEpFGN
MvWwVlS5ZXTIsvJVbkHFOnveQl0ULvVWTwmjH7XNzBT9rTm1ZmRYlCAdlDCZU8Mw
4/kpqd0OFl1d3T76eYF2pINFEZ+SD1h79XEaUUcw8s3BgYrMWb2lORKToYuyycFx
98qWqJNONs3Y3dmts9G1jRmjZ+5SUifI4u2y6UCD8xcyIgoypYxpwpQFudnm5gwa
SgvgQGrZrdGaDlgkwpzwrlq/3XA3nBkGbXj8SBdRNOM/8TyVOd50BIG/KJ/qcmBG
lNrmZMFgEywMCbChOlV2uiHCpc/Y30/GAN2xne3MfIvFP4owWBqKc8wjT21nhOAC
xtDp04vZ2JHQqESreSmOBfNGIu6lG6Knl9Q8nrlpYeHvTzFtMi0sj0JKwDEO+AV8
JBJCGhaNYxt5iyUsk/GsrWF9kums/oxfh4FcluNycPU6Ke0TksB/DG5Kl9j+ceaS
QE/fNAFyhn6LHa478DUPn8Znl1XdI9z6fBvA/l9PzKgGewlPoL2yCYPjzNXYPn/b
uJQRAmwMHhXoN04BbVx8w2IVhHJWqDY16MFhMiV2mw1fkDJfZi9b2t5BGEFGg6lj
Bwt3O3ZGfGh534XCO6NGs93MGa7iivGTkxaENDH4CLmtK4dBcX952GtWoesm2Q5O
s2LDbYJ1btDaAJ5l46ZtfLhzW91iOj8skT04A9ayneWrQD+bp3SSKrYo+tMDLM6V
NNB9q8SEJfDTC4gkdJrFAtprtbajoVy9xhTVOSlLGgls7pNahV2ENar6U3FLUcNd
eQ66ltkeoNqCVi4/C7aVMiyV4Z3zh0D6WqYwrwq8lfZgyoosOJCo7WGaGdQTVrU/
H1QeEgcE/l9+M9QE/oW48R2MOlK0o3M4EGvCNqyozDjNCAYgXFIDszMUuLJFIDcu
CZsONvBH5cuifTEsmYw3vPmfUq18i881tbEeyeFRXlTW+aiCP3yfzAInveojcmJa
jERq9DqxrRitygP+ZwKnrnjIL3+j6qkDJz9NikeW+nZ7YxIx3SBgdOer03vS9GLy
Mf4jbtizXTQfBGVSWpQzodeRNeUT1b1FHs+FL+eYaI5PZsXJdKgx/yUY8EKNk/UR
6MiSDsCcqNZDxDtedRYazJjfLGFlEslumXOrpqsDBuBdS5hvIfMwQ56trh05KHbm
70lAC8DUTIZkw2lGycG+2hGoMrli/Lrs0dtYiRWbBjnlXRQ5eXdk0kBWQG4iPYwS
BiG9Tk3aeSUlqk3vetXvgXErNtWPkPVTZUhLKXF6qrGAOYf1XiDeWIq8vPqxn6mq
bini10VlJRJwYcNfagnlbK2J81YR8j2N7N9nn81kq2Qu7o2qHKpRMkIlHso85bK3
EWsm4/mAA4QtNT/eNZcgfRBHGJaWscJl1RI7ow5q3c538nQd1i8xkPj5oqmpwWDx
AmCrZuRwJA6ZveGcXM0rODa9yAlP4jo76nkqZlWbM13+DMUrXjJVPyPjC6/ZmHHK
C87myPklxoMW93frs8rwEnNFljS88lHx06R+kG9GLqFJEGhDmoGvfgK+2anIckBf
zPJNJ51IBlRDU7hb8B0NAkOB9O5QmoeadQYY5hwRvtsM1Hp1fsP1zP3O0qgiOMo0
idSjbkFyuKErgdQ7k3Ajzu/CNjHBlezTnaFkkHRniQ6/vjrYRQ+wBYipLif4kUZ7
OZjnYuEwrht1iV7G72pbmlL8ixaK1570W64vyKIbHBDJMtji2DsUybC6ZFIfqfXj
twBsaZQSzOZlvhaMBerU/KU1D2D8CIV9D8XR68uPEnrvMjahUh9WMK+qOJ4Lv/1n
ToDH9o5ouKmgAHAYJB7YL/EPdG0h5gqGoSYrl+zvmpen89rW2oifbT4+k/MUoXz/
I14HcGku0EAiw1utxLn2q7xCvZnfVx4Trc0c4zcfekz/kkHglVw3zkQ32m4G9p2+
Z6Hm9KfiA63iZDFw7u2Krs0+e77sl6m30XLMPnGlBUGrxrotsoEALPBu1U97DscO
YhsiDNN9k4AJ52/79/1TWnQL1v++zWb6FaKO4q8IkMSRZLr3KKgcxB6EuMusP92Y
b7nNWK3YPEZtG8NAp1g0GsWFTDwhuVW/EdQT1gGZ2buxh93lywMVMGafx+S7RD09
tJZWfF+DOSAe537+uBJT8/WOPRGq7wnbU2S+ED5sZTtlSEGIxF9wCB+m5iYzQ2R6
ECgg0NjaUDe1KimME+rwS+SOTv0m+aRuNgkiP4MzYHrJO4KjZ2FC/0lfau1XXt95
Lz7mQCCku+FIOn+sXrdiu0CAwk2mLadtUUh1X9wAlLO21myXvTkui/YDOybmeJaf
iASAObtmH4ETdfpD6gp0rP2xgypBIL4XZaLeOJbtzHktjtPICYP4TRMrHik5/KIn
qUmn243+ZdTF5yFvfWL/Wddo9B04U7PQxrnowfI01OcVgseRWgAq19R1snw2IUEr
NWYQmda2f60H3RczvEBD1eDzL5jE6jYDXu5qDnhitu5cgDeb3w7eWCMYXQuLcWxK
Jg+M2Jc3/+BA00D2A7rkwGadbOun/ui3hUwGm/QNtHIDl4/ubPWTYiSdhe/os87I
y8K3cLO7HAjWXvAwjnWeYh3iOm7bcSa1D7OOqP9tcP3W/qAH/z7Dywp1afehUVrH
dfM1PNW00VOryyrlagr7Se2CseUKq0w0spq+tz22WxRg1mIiz/R8trYZL64s9Doo
zcQnfpHOzDBWKghAzRS8OddxBp2dFun8BjNG3qNlDQMHi2yAsBNhdL+EjxnomYUu
DQRX0btIyPOzUZwZqLZSeJV5TZ/lUVoibJzdj+xGtfXtk2r+g+QVbtPC6XtuFBHe
B3Pznhma5iotN28qlFYG8b9JnmiGC+DlMfnJDbohYHDSsRrmVD2BJZfCqzu9txFZ
PLo3CZqZAROJi4+t40iNsI4jGJ9loOGUnsXDmdSOHI8MOf/g2s4t9iynDGdmQ68K
IQzaTzlFDId0E4PPAQ6/jMLv5CD2Nvv38SWBJrcJW65jpVq59ajR0UQVlrzboJxK
RPLfYdYtmnNXxdKbtX1qQLyUkuOqtWKEjm7PgsHHEn53vEXFYXOIqir8qwsBZfli
jouK/l2gJ1nVeIFmY6l8yk2CarzRNB92+7kFYMMVXxCFu4YpqDOAjxG3gpNGFQPi
jFCzThRHqAY9kAEUFkseUZQ1BQ3nADL54IYPcjyfLZ1105O8ea/YMwSpk8oqtKKP
EYpiT4gHslXpA62ku+anzjLbkNqxgxUWhGBkgJTGqOtQIQCS5qttNWLf0PK8XvtR
h64FpklDyl4mVAac4/EbxRDk9tsGZxxFnU8iqbuwZ03U3OX6a5FGxKaJYWsAxHvN
096NDkjYpoRY/FVrbDKF9mN/04+iH2RGIezG6XMEjm+gDO/FiCtTpGW3BluEALLT
kOF151KT1937GeNMEqrFmkRIiLWi/ie1aNQDgXUZGo//e6P9EeoFLo3WoepZ+r1G
/g8ZOpFihKHXxFgW5ggN1nkSyJORRZR+bCMU0N++yim8UvYv7L1d/qeldFVL26u1
Dhryfthdc0nPEiytEB5uwmjWeDKqxC4QkEoBt+M62NcdaFrK1xfmAjpisDe+0i/F
3YqBV4ANWcrubnA5pmLnHPnLsrJAdzyarXSuM1DAQXVe0Pt4DbE1ZnBbQk2FEnxY
q1tc0nayKRzmG6sE7LtgdrAeBPL1Z9/8jgC2qvVKPoXQMfxn4rd3YaNhDf/8zUSw
CrSPwRtE+izDGuuE+M7FRQ05NUYAzCR/UdkIosAsYiUhm75ItpqpkqnqGEqzPjA0
sCTUhyy/p/RYFVaNJf8NZqLKxmqrCZ7KdUpjsDz0/n23FXu+pJXYXs2vqjU74AG0
k1BVjrQonCl2YbCKvSr3e1dxSp/UA8J21hUzXHCTVSe/8gyUKvjPXDny1XsflldN
W7wLQm+aq615YnKXYYQvOEerLfQFq3Bhzxp6iSY8EmAExOg3W3u/LNkfqhtNiOqq
v8H+rPDM9Z/QjNKJ99GzQZJe4KmH1TGTu50iP5lvz0uR2eJNZSArigTIjvCiCDEQ
IzIKwWfvXeb7kJiwG05PTeowfJ7p8A7+Sf46wRDJmE25uHnxJlDgopLIaUW5gwsm
u6/c1uJvbYRg2zfsgiP/gdAHgZEPt9kFmfS/FP4VtD6uzVV8D2o78JAlPe9z573o
cz/ywvPdRcC+kMqavWBdHxNIkuRAt8V3P0ZjH689mV+kIpedCWMpAfpC9LJmpbn7
qO9XtLc9ZtnShoRRLDrQ5ohu8XoDBRnO9kDpXt08kIYuJKVpK9K7WTvIF/bkVo7P
vRXNXN8mKF8jLULZdYuozzlqD2AvIG7WmL46cFDSQECgPs+ZUU5tYnjNgzgfoz7l
c3AoiTrutfoctMDpXuoIFCtkhUPV+bsXbJI4lOAN0LDemXIfIV2GhqszKYLb2Rd2
pvWfuuh5BMjNfXNKNKX5FyhO5cKIeI37/bOikqE8V2P66DieWof+68EIohhnliQ1
f+SF4lXXIRIgQNu7FTIJRApsunGsVGSM18Ez1hx+yHWAxvDq5FX8w3u9oARQSzZ/
ZSUYl9qNKlg24m1kjTZZWqDZxjU8OdGtGyOABa6dHw3vkzCTug9nKpdlTGRi0iCq
YAbDNINoXFtep7USuyRwL+7NaNA1xUZpE8Cv9JC5bnZdoyzHmYSXpdVcrN16rYL3
oPsT1cc71Yalh3qMRj83SB2NK7UWWUvF8NPOwfRvLzXDwojFjE3wZyCHBS8Utj8y
EVTRY61PrF4HWHjq4XgWDoQefiK6cSle6PM9aMBO39TSs6nBmPAk+jtKC58wJDbN
NFaCuP5HPgu2zqi63QWeNE8h5miFsmNPq1BweQxwC9BjhLVK2vQVYPlKMNS1tmoG
DKR7c1FG9CIpH0tHSbVT3vzQlPJabJUJVHkYzxNZxlF2HZZo95P8WG8KoiB0h0rJ
479+e8PuROVEicvf+aMMmljOGB32Vqpu0eoUPmTIeulx/W64a4qIyilW+IrU9gX/
loffP+0g08bNHAl1FOT37YT2zBXZ2LnQphTz1OALEVx7NcS/drOTYMcjxV+mj1Kt
llH2l9qGTbZtZssALjeIdk210w24eBtq+gZX4pDO1iurNH07k7IcV+gt71epnEbV
CjUkiO/AaVDeQ7mDWi6ay6cHwTtAS6O1DpNCcKfeWVOP8e9rBxpDzNDTlKU5Fixs
q6eE4pcPAHRqeQY9896lAyhX0hdwCgfYkQf/I7drPZr36W3lQj8RRzX8N8ey69+U
Wwfqq6Glc9Pp0TpFsQrxJ8C8SiPdP639K+ADPPAYExoGtZHtxmHJKQCfHt+rw7fV
7tzuEYbGoVP07SYfl/HhbarOW8rPFoR0jDgP3cBG9f+j5cxJ/Lbxeu6V76rM5PPO
VTxqL8dM/2V6EjE/4o49nXvRHqvaJkBzlHLUKSn7/jcILfDoJLLeGCaEmFv5BJuP
STQC639J9Id1zuN7kWBHaAGUDjvwXoZaC6HijRKCTty9irsrPlLlGvSMItDDd8OY
0/PkWZsbnHc72mCMptW6jXupluVRzUu3XQs9MNfm6DqMYUO0uvHckxn8B/xBFH8q
LzJzi9hHDlHib/B4gmIGtOtCa/gEohQng5RVCTHw3ylktnOwkwv2i2IGA6kRsBfX
eAgoy3xpF34KNxFizXO+uN1HkUNHafFwtZ9IoswjOFAGsFOC7rbTrXvHRoSmbYir
Ug0/NK76UyayWILraboFPVMfjq/WvZ4duuDV6CUHVDVq252a+lzvGWnlg4HFvVO+
y+WqzQWCgDPr9mEIuYDQFdcNK0WaqIpqReQ/bt589AcJmF+XLMD62uUiuro+wutg
UW/ZlDKIHvDc8akGw5z9o7AsC75XDZZm3UyFhI/1nIHdEX5fjexSU9HjY7B066eE
e6HEWqLmggwyvKFmhCs57n1P4466q+Wt++Z74uG9VKtlnDPS/bijmZlf29SJlEIe
om2xyRwGSL9p1w+Ojyng3xWwy+0dTNdRbQGmuUe9DYVAAWHQWH7yzY/FgNo0bc3p
Sbl2JP+csjO9X5L1QTRofNRULcsvJXOMl1PNXrazfwEyLltc8oPc/lL2DmV5hdNx
xqCTV1k1iHKpnujDuU8Mx+ClYUD6l3pwbAf9yc0HwJT+x22jdnsiRg4QYD63gzox
tbL3GkBK/XbYHCRi0WZwgmrWVjtefBr1nMxMY8IQdmR35KcAGHscz8yhrSk5oNIy
vx8w085wFThdjsSnJywUZyQ7sMT5nnKSJw52TrO2a3+BY81W42vcNMJbk0q1C2jX
r5livIzJf7b1Q4aHmPeT6WBfz0FNzxeoWXzam+UhpGJU6Qh15iOwMluyhq1eXTWu
fWxLKmOlpkuqy/zfznVtB+XDHWQTycK9bYe4Hsob3EqlKQ6zHxhqGO/6E1YISRUk
v1UUfDcCEzrjF5I2lmrhyV4ty1SOj9mvSZTipNU+elHg2yjdjy4Eyi3FgaaEViEh
cZbgZMac9N0OCf6eBqkziPOsibkEw1DiAcm4wvDYot4lTxaamaYPAxAxO0O+PcTZ
8mKSDTCiLdZInAeU5Ug7A6Kqs+7c7kShEjTnYPBPkcWLL4c+fm1Kb3eGSFHbBFk5
sXXVJX1J04QSTZTmzGOo6vUIqIDppEzkED6QsVtrhvGk6ZZVXB50oRDxi0LGPUwE
ZBPydnNY083wsEMMfb5obhmHZq4rx+hli6WDpdXLaREBF/1JK6xUNk27qsVL/uCp
foTkzY9fnQEG5AruG7neOwY+0PWMOLnIBu2n1DAbPkv99gr94yrfmEwsd0i/zTPm
t9APJEnqPv4Ark/bM0rvTa0nKTs13a4nrz+WwtPqrlJM69+TDXqOuDFUEA5B9PAb
9xuRxvsgwTGzdd5ziWbVhBBHJHobMlilxFrSifInlamqwdsXP1MIOd0oJ5mV1Wrz
dVn95++xwwmqPKVl3XGpWjFRNj1BKve04wEmaFHoV80BMNWLZ9jK3/gsPtS9y4ao
8ouKR3B/ZXiVPh0lqFWkKVXn5YwYsimb9otIMB9kbMs2TPziadFu6o6fr4nn2Xou
CkuKGe5c7ftMsHRhIwy3JzzR0I2qIM06XSPjNtQAKZZ3mtt6+s6OgROEOkXcGwVn
1RX69V/34arWK5lLaHIED7NCVJVa0j43Y8PYAheaYOFi7G1h6X+1bW9QuSZkmQDj
thUi8n7rG/7qnSIw1qQP2zccsdp2hcNot5JDbdjL7GN6xbMVN4VB9nesjl2ZhApD
u0ln+1QPJQlMP7aqvAjWw3JvT5h1NEesSn+2a4b91UpTbMf6rLWfY4JRXwVjiusc
Vu2gIi0iSJyutmRa0WYD/fe3WrBcZc5YE2G6zT2/mebqGCqgneBQC1dqRtuN8HeY
sCw50ps/0loNu7fryhtxXQx7E9NP+mGerjZRUo1Lple4QVJdVqJbB/2RFkKogi3m
nsL2xWRbjwIAzgkM/b/RWedfLjTfUqWTofRHfgqvRuMdXRJbWGnjgMxmk/OaAD18
uVjLRk+OqEoW039dZkb1j6xqQ1XMcqFtKc71AiI9iOItgy7HvPOFz8Vi6DzQUpt0
Nf8gRIpo4iBl+nwH7urPBqJuh1aCRIQF1qaa06oGYQs=
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jwdIkhUw6ejJEjwHqxbJ7RIN3tA7T0B9R4r9BkYqjMSD2/x0KRDBUhoVpVZN7HB9
jfgkPIxM1710RuQ4VuvBFTlmKMmILtYMlfscfNP9uf6DX+knW+ljpaaUajBmEwmx
FsIEb78lKtMqkTbb+lh3Zn5TGTEYOJYgc8cviNVN7pVep/HXV8rvclMy6C8swLy4
CJBmKOa8gumkpEXlisVt+LWzflIbJj09I/W+7J7hOOeuZuMXsIozFT/wZtx7q1BG
zeBu36VapyANhf+WlmzEXr/rXJOCaF36BCVNWzST+fNgMWUxBWhsWdtoTJWw3nf4
6sgMttBMWIdJlnF948pFbw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5040 )
`pragma protect data_block
I/LvWgAWlnG+3y7fVtJb4Jq6H453hY+t8gyXZEM9SaD+4oX6kLmfO59BnXkRPmSI
4T7EwRXTPuuNRzdd5nixKtYUNNNu/HHUb5Kltmv6orMsPS00RHs1ImxeZYoEqaHu
isyF7Mz3o/qOX9oYPQtLAAt+3J3QlY4UD+/exeFrTEnvKduS4rDkxFCvefm87X3f
w3VHs5Xr+ek1wj786w5RzLPSyIiDLgNZVKDQtOhSKFn12cYGpaOeNZGQVYodx9m9
/Tjx6v7f5H/pQkM/tSeowkguPni0kGnigWxCSjT5+mCFl3YfiyMZjsxuZqkHeeM8
UNMF276vlu7B5/4v4WhLWVX1gMtYsIoSxAmLL2K+39wH+1T5A6WfO/Ns5i8vnQZ5
YndSIMjrAo0WPzK1ixT5R+AqbGO/yNrSyAELUZL9UWGgvppZ6bJrMuc0puZ4DNsb
tsOA0eCTzs8MC1xAcxCwMH+IGTz/beP8WLhp1T7nTUgAdjRldrGftHzXD4ScDCvQ
RfMWCzCa2H6jDzbzTruuapN7cuZdgCiFJaLzSbq/Abc8fpj11VoR9CGNxlvcplcX
tCac+ilg7fTSDnbGV9Av3QX2s+PGcPUbMvADl+OqYS83swl4JvNMN4Ibb6WEPuTe
VJNdrrx4oeWBcaFldSNQfOUqLJD98Jmfw/ET9DqXvOpSfd9Li70VotCl6munxP8G
YU/6yGPDDU25VAPNRPAUHjFv31rc4eGQJHFdacWfAfRRu+riclZK3KYqW531HMP4
+XSjb5DtZYN13UfC5PirqnvoeQUI9G9MsmEJQqj01jyetGS175hgNAWNTDxcxWI7
aZKvrADbvolIBdH7PDQZXfJBeRaeM7MfFj/dzfsPmkpcxelq7fqApPFNaEDYG25d
PGyP8+zDopIdKi7Y+hAzqhwThdgTMDL156GXeUDRLUe725RPczqOPykLwZTTvGY9
U+4NBno6vj7oT+zMUNx3Ue0yLn9XE8/5AiQ7EpjS7VLbdKmiD8x9y1Gyk3zL5rMu
OLNm5MD62jaEG6mc+vDP5ACVpBKwS+J9x+fV/xgL0uSA2KwceSq30uXzHQ2gV/Hy
yBbcVF4nLfFLI3A4HSxvOirogn0TzTz0kgQOoIQivIY+Ptv1c3TthKAQQqTLIs97
22HnDQa4ugSVid6zkhThjWHE35R6CzFgLbgn/pWc2U6+/k4J6CseU/666ads+UCO
Fr7b/Bm+LHy2v8w25l60oOyShvI0d2G1ZOJPv7w3WngKAxxi7WBoIizwnV45wjKH
zFxiZBmloXhUyYU/uthIRWt1v0L4Bf3pjjmNJkgA3HD4V783M+K6jyPF2j2+pLji
m6oE8wHro4FGZJeKEY9rh+rflCrKCsUjb8Xy2lftkH2ctjcLqTo88exkKMizqEXV
UlAKPLsshyT+zFbyVnR68RE9GhAhmiJ3r9ersAEd3yYes/dNJnUuor8k5c5EifLh
uWZCIT0lY0s8dc4L7NpnM4a4Ve5zvZhPAsMwmtoQYmUk1kJuecOhZLZtm5CceyY9
sOp3dHo9D3wgnDoWTahKrHzrNMdg+KtdptJYwhJNleE8M6Fz9GV2qf0+px8GIxte
spXUyTjgrxhqXZO5H4S0AfJqBwqFzj4ahfVZu41+xqqKaCJDNeMBWN7Ui9+P2wrX
YHrycn7WUyoqh94w9/KlAjK8ykzw/KQEcWXprw3TGZfD9KdRSNVrb5faHDlwzU/f
8VEnXaAvGzMEDdTtVgqa5H2IlUkm2H1T4uDkT1XLis/k0X0zL7KVXoaHV/Mo9Nfv
DvxOoITdfZNBN2QICCQBF5FMFUpgus2CH9uKP7rZhylxhiOyksvVFJsE8WBnqTPz
8q9T5mUrUXpsAmUc+2WVxDYkv24Nh8tHgngrEUtoxBJjUnhlc3/BsO7h8l8nS+tW
MrNOUI27mp41Z40/P7JJ0mhmXLPCE+wL/dMp97J5QiNKCpN80UJeKGoU1H61egL2
AIrldMsV4+R/FADVjtz1Fvr2sA2UK1BWshXY9vA+BH6+KIWpHXYdnME3RD0vkQuG
bm1un8LEIWGBk1HdGMs5UWpTBABWAL/LSXXLS6xwUlCpQVnLb/o2UUZ8IoIxljsB
ApweTOf2QUkyjWW1hfd6R2lJW9zMu0IzyAicF5kSomonWU7uKEhnHbIbIZrzF/SQ
Cuy8Z44DV/lcKBSYe6r5j1bih4dXQaPW4E6Iiil9wV9aevZUa3cF07LUPk/JomzQ
LYQc9NQ6MTws1G6+VSRdeLu1LKnU4eb8f0JHpUtjHp8PAQUjYmSNYF+KClOHEtOY
XBN6XYwkpKRNyL3TOxAz6Q1U7H8qivYCjFJuEPMXrSsldGuENQ6ieThz+UlNibkb
ZEM0lmdr4+vixa/QVrfu7JTpiONtogE+3GXu2IJ6gjMd3wynoog7WKWtXYgnZKRe
2upfk0JqsQs7KvNqbVLIsGBjJMLIbLduDh6QpBoT5dxmDVGVe4rHoB0kMlJu3/ZN
GGlOtfVwzNqzYOBKrUxvxQznDXhmCtnDm2jsh+lWJUnroBv6Ficj9d2fouyMqRQS
FbO/Apx6RLNs6asa62+a3IRrzW/+S8bZE1enwqO/vHKHY2HdDvAnaodWT3tbb6Mq
HQIfZAQ/D0QN2ItMs11yu+rYVL9AMDlhs9f3N5cjR5wQEec+7btloKzT4QJ3P+Eg
tAmrfBscYT/R2RJO1Pp9LZHN2twtIBPYPaNuT9aUfEAtAyHMEUSTTxKy/knUQa3S
nv7WyNsknAp5oMns/5rJmIX12/FDl/Rhe6XxcpMCydw1BXWNpUL/YsOf/zX/kqny
lW+GgArbZla1wkuFrEmy6nCp3HpPaSznTTdVc723AXjlprl+MfzJHl0hKX6tO6W7
gJ3x0E72Dpb/neoHYE79C7by3EYpflBs5aA+w0Pjo7qS9O+PZ6hYGM6o4DrNCgSa
/STCV2VrBhNxDLakWy8uUSZaDxOpNcTQ1zM6KVwLFdB6bF9q9PRwfcws7i7/flGF
RsKLv5Ne1gsjmaxlx/93l4z5fOIO0un6zDIMDe3ho3Kf0o/2mW42oC/Pj5hd/qs0
iOtzE1oMafxc06ugLb8KSoDnmh0e3giS3G+nf8CBJJoOuT8A1Ryp72e1N4/OYJqU
YAf0eNB+xv9S9SeZv1T+WjstBsg/59255A5OyRc4H3SM7+es2qBiE+YTXfSSraq9
c/Pw9LTUho07gxB+XaT7at6av/+6LFj47N4S6+1gB88GKei0oHXysIUnFOKoLsiR
speZT3kIgEgnGlRkRymdvIoDNZ+krL5tWWqyAqlKx8UA/ih7mX7eAQbyLI69lwO+
bfueq6XU47U8bPVd9R4LTjwi6i5IzvVvYeHCZ33o1OrNYSQbT5Qb8DHf78NXFJy1
dnnRUpjQ7x+L71+EJd12AvFLJNYudnWyohTjOfs4dFpRRbyN6iJhRTqvN1sJdOkL
L31d1aFxMBnIk/T0z7POrr2QWyZaxIwjDWujb8qQXODVUH0nAJOEP6IzoSiGQ1tV
rW4fH4FMQ3BsAcMHGq/6KrAhLAj4akgP9ttnB7FMIiarFQzK/N76TFW6Q6MDKQUy
o147xFmFuMUTMo/BXQANiynn7w2tzEa5yuiGco6bg2zbU2QrHurze9XvGvVdY4fC
2E5fZko/g94GSeqJfPZDCTjcjn7WOtayDPzAm76aB3oFqvZhnu9MVkRzvrzr2y2J
+r2kawIT1rxduRIfT9HqGbtIRwFv9XjspBQ6qoC02gYV0NREwfTsyB2O95VrReec
06K+WjJasDEhNcpeuakp8BzLoxt6dbKjtoIufhGHmMDG459qHmEF84Xjv0yvyM1C
mcguW81bnHbsURUvzuM3EC99QZool0DxL6jOT105O8uL2QGAcL/OnMFJ9yXRdm0L
7VSNGT0NMAfvjnzTOk2B/yCv6EvEjj3Ll+BZ4BmoRJGt+Wuqcog8tDgMPPgbbBtH
7pDjzZy9HAzkr6sQxuyhzXj1wjPws39/zK197Y4x9FDlmH4xfEF9ypVnBo9aZYgV
dLWnezqWOQnqPuophDJyuRWBptKpb2zJvFjdNWKf4ENXC0gucd8luoDYyMBBP9UU
gxyNMF6HZsNqZqyIuH8n+X1Fm986M8vYZ8hx4EJuQel1cgeq1hcS1Dj1bmNZAnX1
TJ6IvqKxpj61sPaeVYOqL/pQUUgDwtv4HItc16oGqCkx3XFH0nW+/0Spl95Zodnj
pGl5hUrQn6IVVTDGaXdccO+uHoroyOsAz3DEtTpVzK/lJhABo2GPuJLkF/TnccOP
27bIwYhbJ44Q+KY59tCa2N9Gdn+3Vvejfgxh2c6D2JXZ0kyZMlibj8MS0IF2XJm0
TwlkPlO/o/x9R5dJh+8kB3Qm+HGKQlFH2KxvIW8ua7QMGthAl/UQksvB5KJkkLXp
r5hQseH2DP/NexxNQNaUioSs0GZuBqB23ZNP0txVjhn5WaveYchyJHXanCDKQnnu
bn7TrF3aJe+zD8Q0xITsQDWMIh5Rm+fJqHRobmvbXkQPlzcbSkXoa0atAfC80d2h
r9swVjAHDKbkMj+tTwy4sGc7xIrd0GlTspRhNcBvu84ZTKfYDBnLXHlt9sAFB+G0
gsN8O1a4vtrw59va8sQp3k06krOwNz59Vl6Dj2lsMyvs2hYaDWLMB3uk0VCkocFb
crivCDnKCSnBnGOSWW4f91qUceIMiI4EABYF2KltG60F/LXidNEshnfU9VwTHgiJ
rHgwb3bojcLgAO9NHXgsCIHlYiDqklZmLiFlc5puOs8IjRF1rB7qNv8Og+0VjXny
IELEazzfwfYYf4yzs5yFZz2WUkLZVOWnkX2tvOoQrFP9MpveFHmgFwBmaRQ3AazK
XSxmfDr1rE/fSyEB3l0mDrYByVnWqnQu/cMW/705mUrq9UAVwXpuxcjHbETyf6aH
trHcYZ+TzUoXCAxun4hMu9IHipij45aDRDlcVdUTD7qnBiAs3g8yz6I4YjnmF8/o
E9AGqBt5YcLRz3IiN9tlQYEhSm2flAPe9nNbVbgxkBz/m9NSgdsYR4ohyXxkaWDS
gdaOIyRd7SPUfbzVD/Q42HKNTyT16nWan+3s378yLRCqhLIFZsA2lIgbXK46vdkg
8ytU+ESCHtzxkuKpDmxqA+or2DPDOs0IJpkgeIgYwZj1EOzt6PMPsqqFAqh/6phs
AfmbDGApG5pl245AYJnRuEVNVugQjU2I6XvkvJ9GMAuA9U339Vp4HYhVBRAsgKEV
YC/Rhs1SRrPILjx9/bUWe8ArwR5g40pN64/jpHfVVJS2vJi5GF6eVEvO5ZRE/7wr
PS3rbYbf6h9tg6XEpNYax2RLsePU8pFbrSKk6SIARS3dSaP5Z7qEgwrHVN8EeHIv
wB3L3p9DTZIQGqFJUY5FVtXZ6D+OhuvtwAfmVPrkFmOjz/sAvnDeHBZDrkmGy8u4
AgrqeYSsouSLO6ikLNtO3jZ8IyyE0tu81p/9WetIEh+645mHtn99SiCQ9wUTI7oK
rbdIolXj0F6RKvO11/rFfm5psy9QsT2xviCYiE98JMzwol8VxQjE39qACaMCK52P
ejaFi/0u/kQKC/cQoB6NHS7hlc8GL2C8DQswuKXeovfU/zWtz0tQOLokmEBoTjf3
jc4HeWbFe7mXYgrhWvk4koBN8djnDzJXwQtm5Eo6oGb+G98mqOgYWnGGwqypNPSF
1nWnUDMGIRc+oXPqSCoQP4Wh9iUYfDOZivubq7yW8MqLJiny2sQGq87+WeqevkxP
C0M4mY8kuMCLMdviXuSzgODF/0DFSXCjFNizSR/NW7zXTB0TJuthvLev0aShbxtR
QbKykwbBFnvVxA5B6sTYlJzd/TaU/8pHSUcaBAjVImix6UZSvF4ZCDTjnmi9unrJ
Wk2FVNusqL70RfiwVLw0cgra/PXfo8P+pXFXLW2RUdkQQs+Ot8YhEd1XHYZ8C66o
EqzrNJc0CucfZcKVBXpS6txPRCXd0+ALLuBZLeF5RU5L2tFV9dEXK/ynSkwh+ZmY
YHyrX23qUpkmpIfTAsJu/E5hJKSK/1r6l1IuPn4JN2iZxrZ8/BBHz8TRaIMkkS9a
2GQEkLcuYTPOVbPnmO9sp7krY6Z79LPdo+gfNJ0385vuAvhf/tOifSDEyGQ4Jh2z
sgI7aVW/AaLRjoTSqXmz7cB6P3rJWl2qFhkIwhdrPq4OjAzdtTrPn0MMeny0KEfK
kjNYo9Spmkb9WODnauXDagmC4sJ4o1rOkVRb7Al59mPox95l7Fj/gazbINbJ4bWt
eSrsITc+q1Jg3CZ47qt8INllmGrShrVAhCAALvDZ9z2HAcdKCQUhwo25AME8/7kC
ggeU7dGU7uyWZbItk9u0ZDNa9KvykoygLPa7QH6b5z4t/Nyfp7HYho1YYuQzXVuh
k6DMG1tTQ1uwe+9drJp6be5Fr2A+G+M0l/cy/c4Bp1/tubnNJfLdTp1AiSz9te8T
vt3vHWXq/aBVGQj8o0QimsOlGrZsD0x7Am2xADsMKkLXqc/YsdFCipj+l4F4YiH2
fyiIvZpK6ar+2BLYx/hYxyw3LUDjn9ItAgYo5wXMtWmx6xL4sD1/DThLYC1ZP+WZ
00kb/Q5q292/ibHNDj7ByFiG5ey0KdFP69lH6Iv/hgq/KcAWPoy2+YcgVVkyOw/X
FHqeQ+GbMMb9h5/WTskVLc/B2UD3kC99IcZALjPqj46gEp7LgtbI19aoPoe0wuzK
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
O60yyHwrmVAXA6+XyOEeUvEhscUD5tyzq7H0ZhApW5PtrNJjZvHvphKv2lfpFj+Q
EEp+zTYzh6+DkIptVbpADmOk4JAvjc1YL+2qnbVrvq+14DMwBCe8PrtB6HWyFP1M
OG/lTrE70L8Z4wg5xWnUmScyqSo2FdnZTYUwcYn0zUaH0+NCUwEFFjT+9m9S4yXg
nKjwmLEoVyulqvkM2l9KaPzS1mOisdc/+xOD8q4AC8edOLHuxqFGBcSSV9gy9E+L
lkjheknMaeHxJb8rNV4kidh3/JpuPKBJOHpKMS2r4+wm8nwMnoYwOvkIDhx/zG8l
NvhjrLTJsnKWhyM0mwYhKA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1072 )
`pragma protect data_block
MDp/RR29XRdwp14ZaYI+50LM09avhRsN1ybiQkzCiYU+RiY8opZtuClKtDM7vgyc
FayfRc/pDv0HnJmc8KUYoBA64HfAxu8CKhJ2nMats9gZmUBIDs3hWeWLHGlov1nk
CQrL5cn2Kkg49XTctu7JXJOgA+BdiDCNjdxufVNOZkx7rh5i6KcViC5zUjmcW5+h
u5ASZXa56kHTom9SDZw8CgD6k8pJKa0Few9dp1YM2UGoYLjrJwk/eJc0/LYrC6sr
mb3V9dC2P7nGPFsFiU1c4PL05i+TZtdS/cP9UQvUV32vi+MrhwCW2HhtPSroUjvY
ucIk57KH5fW3zv7D8Vy+uDlU2wCqqLQ4OBrYRGa3+USwkbyZlZbfCnOqnKT2RxH3
x5sNbe/kWCdfEoxK2a4K/UgIMaPKCGM9vpIAoyO5tEQNQ2QrIDsoAHbNInBgrnQT
HcBvEGfnNnA7QkgTjOrwFbKFG9PNAlaYfvS1y6uJ8Oog1BL6jYHPAffQrSbyUJQC
hP8L6PgO5Qq7JO1Ts3EvC5LxGIgiHEBHxNTnf2GHi21Qm7ce5Z6sDKBlrfoHLhd3
HUkyziKIr+J3dff8/CDei8dRIwKpnWwvwm2st9boWtenmw9nadrWvr6O8IQe8JSg
7KDjiZf2hgiNA1nJX5dNJDPExLEtFRrAj2iP9fNOYDQKFNWBf2DNo6QrnLflbt2N
jucOLr2uC73xzZPS2PI6VkE2YNITLQ51egtU+oDlyXIwN9W2lIXDkJYha+ATb6Qi
ZF1VkhRh10WSBaNWnj4/vL9/jhtxbendN58r27jdijuz5x9n3zyTui1L8VVtjCNM
HkXZMJSDX1kdhHpJcI+rnBvVmF2PcECRoP81Xu2kMVf9xPw9aLYeg7u+iFA/Dgrt
DH9RdR/xj3+mAA4gtFTJnJsNOgYbdEfXU0iz62m4PxmAAouJgaZXxc1Hys2+gHLh
gRZ8nIhwLGFat5ZGHsPaJAAP92Gf2SbLa0hCaKcQzBW5hBM0KoUbImqrzqceWP1g
pU3cMr5ocUaR1E8qwjjWaut4RAWevCSbGogPT+Y9ivS/G38fZuRYe/0J33i+xeqx
LeeN+olFArB6zbvtC4ZVJZgWWpB9z13KSN89QyOl+YAUtzPyTl75jjpAZGas6ori
OnpHk2Bi2sdbFskgkcJEYEYtx50Tl4WhLiA9hsoOhweoHYjtS3yerMO+c9uIKTTf
ucEZiMQqntATGhF18Fi8kH7TfVT1qlORZbVdWZdJHIXfcZYvkMO85tF1tMMJg0G4
ccMzNKjD+DZzLfur7sYfgLeZO38ulDD4EdSyBGl2ryIDBqDOQEY2b9nas5gPjdyq
mXt1IYR7ic18t9BfZCkgGavWKRSA4giXZQEOFDuUNl4GeTBhkhExdlv3rTlvSwpU
d/j26GX47WTwSpXoaZ6Gpw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
M9TAj0+AoKdMrEeO7ZibOkuivJixTPfVz/aIuwPzKSpmZ1N7A04xjZhn9tkbWh9m
zpWNwk4IWHEYkCefn6XgkvX4Q44Exk7wkE8vKGafXMKfujG/vmvJy/N3oQSP1J2i
WtTXvEVIJyvz1tu/eAGc/2aB9R3IX4OwTdrR55kx8x3c8AntLDpl6dA7CUKmN/Q6
vmY2fRU3SYawP8V7kjUbsyhaIgn9HOnFlJDKDQ5LSiFAuzEpPqhtyVyMppmsnpN/
SuJgEMFLZxTQ+0Jm8r1RQ6c/doBf250sU8COr/ZMeUD377jsfjmZNztsiZjDxyXL
n8xm+XuarV7PYrF1fYkmTg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 784 )
`pragma protect data_block
4XbjvHFhqRpk3pJqjCwC/7E7fdoJdvb1coh4dsireIuBnkL5s+Hz2xXHO/oMQeqy
S8mJyX3R5uII5yF3KivxvIhTj1/yqO8feHyTLW8VhlV63d3YlON+j3SCpQjoLZpa
09w+vk7uIqVGQ2tQpN4vZB4gOBpCjGBOTnpGi2djXdzZCnukxLtrVqTvmuGzR0wY
kyHYlPLau5BEsTuX/1NLcbsNK/Le6gYsSF4dHOkKnwgnmTNiJEDC0oaex2akcrcP
lN0QphQtFbcXQVzDtbnqkFq0ujj3Wx+aErqhvUVTREIJCa6SVNQ04JTxnP+I65lB
Yap0IaeX26bh3uGlQGCt4OUaZAnzRn0Yg54RYfszjCDLjVOXRsfHDEsOEqpDch/l
wfvhX5EyhC+SlPvU70zv+61nqphpWyJL4S4a9DkRl7BCzp1175ImcXz5JTdQnh40
1nIGj+cnfhfby0FdKjXcmM8goXgWDD6Nko8WKFdlvYflQZm0KfZJ1aMb02ZpwoFw
aw+56fHuw704AP6iYhqTFYsUjtiZmpQ0sdUbCpyBI8QwSfyF0eM3H1XCJ3CxrvoJ
wpNSXE6YMRNLoHf1PZFCnfR01cDSPrPfkaY8Bm2Sa7Ag34R/NlwdRbHU2LItkt/A
YQESOyqoUUut5CgGUY9K724kPxOlGxhwl8naWJjf1kTX0+7XrJwP190cGNZ9p4AX
1uZwgEwzexgGntcftXCYobMCLQ5Uw/Th2B68AT7+BBSvC93GpW+vTBsN0FXu4Y/T
EjyVQNC3RA/YDZpDZHrMIGQ2N/hXdDmn2S2Ovgw32AascsDHTlArn47XL0d+6+TQ
575I3xNkScpdvJdXrb63m/IECYlmnMOK9ToBsBXEdiI0iAmwJYsL2adLQ0sGh6SR
rv9CUXH5AA7hOnwe+VMVmBAP6ECNMr6IfmkwP3flvjqsNrY3wczDFcBfOXOTWqde
yES9+/vNlDQ9sUHaxmk8kc8yfPZtcUzcr7IpqTtXzREVkqOFmLUJaKkn8OMJ3fvd
W+NNTpnYWBAATI5mAspxvA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
IYWBoNFklRr2r885u+gOqeo4zWsur9va9HhbVShBBfpDulOA6U6DALdRSGbfXYVa
wNiTj8WfykWmY0s99ProK+Llr6JdjuoWSs+kUU9RhY39tJGA5uUWvza/+0rJCDAZ
hplSooXl4msHwlryP3EqnxdaODqpMwe26AVD/rrwwY4BmNB4Yx3kwoRgwLyNIJpt
Qv4QKk5WkMYrmSUvCXSe1BzKBIV50xhnagexcLdlRWr/MflDKD39MoE0QVsud7+M
POSMPKKSSGop5LirrOjWArfWeYOUJtUOjPTqMuZ62OyQf9N73pF8XXv0ZhmkRuZU
HoiQ93EL1hXSIo0iauwVLw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
frT7CiYqH+pbHLhbNEfojGSD5q95YzjPAWTiYS92UInjff0CAUvPIP7eG3++JtUE
bqeZ+jX1NhDtwR7KUG/Q1GPtq8XqCrjGVboYWQUUMezM8EeDgwWcGStsA5v3Qt7r
cAKYZMsoVOHfKQ5Z0t2i6L3PIb+6sit3pwMlsBu09n/aBNsxpfjR9D9NZqn6gSw8
U1KYJvdGUVAQr63MirMOYEmF8cQzudQFnd+WSICLcvvsjXU9V0A7Q7gbiIrTDBIT
ZJLL1DdRhJetc7qXJZoiD55Bv0YavufxA7/cp0ejL7JBlEBCE2AJg9R5I3WgSesQ
D2FIkOXZLxOz1Q9VNkBIt7XJLTnXQ/jNxjv5ghe+pCURJ/lJBB7BYGEso189bz41
us2T+XjgL60R6Uo6k+pnOT7qUjsRcPzv/DrfQePrOKlpKrO7Y2NnWpG7YCcryg80
3iTFCOBAmCnYcnG6v2gAu0+B7AaVLYt1UWI2ad9uXge2SHlKOgYU6wHjj6oFSlyP
ca6UesZWpCQEstx2UrN5vEtdhNUHSPrJyJG0wz4y4eRPHWMOYi3jGN3mfzocsMPT
mhi0fWoWzY1zdho92cC5jULJ4WLDkT7LQmA5eKSiMPcT8A8AvjXsEr8rhJVSrVNP
dXvzZVVNLlwb3xUyU8KNOqxRpdQwNFrADftkYjMP0n//97U1ZnkHN5Jpj614TkZN
SOGpqeEcy5BHcRWamHYSpIl0DezLEeo2pOxpKDGGTeMN8/RV1L7un6FUhmCIp5Yi
Z6lJEs8OQun+JKlWp6XA96kDQu/gBGe944ta/84wfPQuuspIudv0lQv5ipBfuFZq
YeQg57FW0otWq1S6kR03XE0EyRbrbIaSMbH99v5AfJUqvp/GYvEZ1w9Q2ml33CFW
3cf10SuXwF7F3CuGoZPaGOM/CQPNwAHOIcMAKXPlgkg=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BiE4pFOYDRC7XCA2NSt8/GB/OLkLNGByzYe1Tof7NoU5a1es+uT87jwZpd0ZkJgH
Hec8UgJ4FDCMtII+7HQfYjzLzm5Z21tNiwvAPHFmiPno2e82S2rgo3+xzqGQMkAB
fW0A73iYLYgq5l1R6MaXoiT2iobaRDv7Nh6rCj+sBDxzmIJyZbYHiGHLupBAz1Y8
NN7jLI7PD6hY7of4uuB6Yl375MUzCCKCAGgQwueb56R4qHGSLOy6/H0kpTZrYzB+
SFjxt0QMr3XzjYyWYnEUVhgC+ASlljpk+3RN2azfEPRk6nUSQkEg7zKWSJr01FwF
O+l4xbRZ6W2YNUfbcvGj/w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1792 )
`pragma protect data_block
up7J5rxniGmK2l8ijeZhWD2qikxiHFOEbYXJhbSB5rSviCiX1ZlsFrrnGEtiP1Vq
CKc3nzO+ZE9R3awm76HHD4bE/zEr1V3H8HfvjjTJuawuDfFHgHybTEVypBoqXjSi
DlLDf7QgG+L09APIqkUSrvXVoCOtl508ho5dRX6231ceCq6xLWwk8KEJWa50PmSX
IWFBi1i5A+pdqciYN+6yqYgSPUFatqWbBTSpcIZi7QTJGLl2Jli3P2/KrSouyQg4
5fOQ5678HaOKjAZtZmVjgCfvdYbOdRm9zlxhRpFIQQhTGEAWsyWrDp/0MtzpWU8I
+53NFggmmXzTmWD6FlKM0EIVmIlrT87l0vZ7l+nGVSN/8KUIhyiyN1qLlJxR9Zqy
A5wO5YR1N2YnX0NBkOR0LZ3r5A28mdpKTUFpMiHD3MGCgL7El2wMAizidDm2f8zq
tZa4R/E1hzsagNhn0CS1fdnbkDFcePff2/YFDwrcBy4UQlde4rbBToPyIVKIrDRh
ld31rwUJU6hEqecX0TwxBPnhSzCpj0W0QbL9NZkgL18qw7FrjjAktUPXowZRGIlL
mhisRBgGfXYy13wg7uGJ9L3t75OaTRKmd4tFIKQ3I1+NGm0r/AfN0rXxLwtHOD9m
RsgC+CJXrqak46yNIrq545WEsTRT1tDRf6nYzxfsV232tOmV9CyWfvaQmXAiHSEo
xuHQuTz39xM3ZVu+XE4VlqbrivR0TjgFki1sEpHcPFKDU9HC7BVIcLqi26Tray7n
iBYbnuClTPeaajE25VKHbp6MA0m9cTTllgiWiDdOiwhtb/LWQ+sEJc3J8UaftNtB
MUKcE5HRHKPwipiMVv3bebGVKp1imfelBK0tz2bhZqH7scw5S9vatnBFi5xtgyM4
ClAryfYM5pm6tIZ7yx0PDzle7SXlSFetilel0DTKEDZ5kpFWIaIvT4v57cZ0iAMn
PQ37wbiNK5S6b60PbjRbEeN9IBt112IgzoC03T3xgE5wn0B8AtvNtD15DS1umaUr
VHI0x9qg3VfnQw4WLIib4953k/wT2Yj5iQtOudrFEkshNNO21m0YoeyPH4G9cWej
cXFKZls9Z9vZR1Wk9aFVfuKPhiJbq4Zk8NX9F7k93k/yUDYap9ngNEcN9bw0/4Bh
Nl7U1T9ZeBX8JBvD+bW9Ko5JIyw8BRyJ4OIQn7KPJKBzREvIVTxQM6o3Wbf5GcJc
Oxx4BUHkWLRyc9cxMs0Rs9Txy2rN62DEKVbmVDvTq1sYskuhOuB4q25Ff2QfupAA
Rxmgr2ZE4U/O0cXeils3oVJwRTWpp9UAd1+At1WIpfc++9X8QhosJhHjrJLsA/xU
4krj3EyqpaLxecoTAhpXJ3vZVRUt4Io5a4prbDE9dmke8KBK3vTcuzHdnUo8bXVp
DuIqaJZm/n/zM001SWoQE8EOaDu3mc9MIQTh+Q90vlYHuNF+KBrZpE61Uwkhs4yr
mIt+X+eEsWZz8YSgpXwEVHmyFbv/ktW9tXBZfFkxDqW6EaP5pR6JKHzA+dEmkUYg
icgHBcm55upq0Aqnpusgr+aPKqwuY5J1MXEjrI0cpVph4ds5VjsGEQiHfTxUO2Cn
zrPq6aE8DM3zyXC2rmpCSVz45ByEGqZPooCS7bpEA4bKP/BeloE5kbOIHnxuZqa4
hoID4aKhmtiO7kUSMs7Lle1PN2UvC03byEDMuC+8EF1+InbJzN9/LJU7FLNDT3/O
c+BqN5lbW6TZHzxMx04yfuRB0qdzren83ddI/kMGJMUVlz3dq0L/9nZoOGG5oG+s
ucasuAqUWkKdjBqs1k0OJabVaCjkVFzOOiYNartlh3DXegL44kl3y0JvWAV+PgAJ
jPfdi2PHt09z3tjcOh6mKEeOVBHpEtcdqLmtSo5OuTiEtS6CMwpZ4DbwNoao3uBq
YdLeXbDZhBn2uPXYXTAQF50nP9WtWn2kwXDeQNtnAGS2z+AJVNOaQnABNqFqnqUp
3Dy/PncLE7wYFlw2MHdaJGyT5bVmvqURmat1octpzSLQ+Jd6Wrhoqm1uNzj2eyyG
/M6I+Id2qboU1CoE/NS6CjYbEB260nO2cWo+sGxKUOeSuw+bURqyjhIgZ7Tpbtpa
yVXLjRdUB5s+EedgcfJzk9i16to/nHiVBZ25bRDWfgQt8Zcz4l/XDhcVhrX2pECd
tSe1xvAs5DLLkhDjOx7kl1Ir7F2Tr8rC+zw5vWxizhpLxB9CcsvX7yIKzg5xj8W/
KAIS1tdnpdjvzCSvVhkWggCkt5Jvsc3BuQnRPIxWRNTCOO+QzUqZym2IsM3ReYi1
a+7rI3+4xmZj30ERwze10FTcQpF7vGrcndd89CSPKJvUxuD3xOH0VwuzCvAPnOg1
OL+641x+0ZcJk7HhBl8xeg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
funn9R47A/b45Ne6SQ6Xxk3ju49JU9j9fwJQubOxk83aPpmEWNkcT20UJhhOmH24
9B05eRiXoFyTDEowx1NXdoYb0+WqmOks4DuOyJgdJZN+dQryPL+rlKpceLzMgDJG
M0EYJGDhp/Vg1q9KDG9fq/j30U53RoUbbP8NqF0DAsuK+/YdCWN1eZqd9tpKhb2o
rrgZrNnG0+ISRsx/n/RgINDkh7dtWnGIeLhOWMW5fEa+BoAC/KFSrG/s8IO0yXGw
Uq6uRo1CLAHnTdtHLiDJoVCYktKXq86UIej24Fu8UjJp0V8UN0Iuj7N+FtkBXQZw
NhYWsyPyaHNo15ki2p4UXw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 38464 )
`pragma protect data_block
YBb0tqt7V8fq/XSK2ZPHv10CHxoXhQ9Zdh4Sltdm4sc5haleqC3f+OO1+LcVmLyr
uxpI+vbS9zdhP+2ofhZnWWU5fr1aEee4GvQUlZ/w9l8bm5v3FgmCAN2n4TeY292i
GQctTL2HmvlL2tuWhflscD0MF7bkkmpgtlVno+f7Lq9j+kh5hxDk9mhi0L7RuKvM
ZdryoSv9OqVKXtfZz7xP1eziIas10NHGs8zsY75ok3fIuB9uO1bd5enWZ2vbgNIF
w/zYt92Gtd/uGNcKOCHKcTiRlqUf6hP5HXDhdrjO540mzW/iSHtpAaNh0N1/lQtr
PNxvMaTaneclLBRNZd3r8LKA6bm92SUqExq6M4Wa5jwI40QeVizNIu12d68dEaEa
3RFQ6DcIwnX0hqCh3PGvjj0KZdznGZU2JCusjpV3r8GFgi+ypGZzolObmB+cyNlo
vDk5IJ5Gae2IyJMTF4W75eA7nkivE8hnrGbir/XWbEW+8/OQVzmT2KtZ7tvN5coL
Tu7kUglH7n++4LnXwDdvyhBKLRZIKgC6r+OHg0XtIk6PPAbsH42vVP9F8KdCv7GB
4cCtgej+CnPmBXIUN+D4Wpgfq3NPrUE148G1LkA6jLsfdhYYn5M+lEEokzJA45aH
Dyt8UzPJhR4mWnU0BAceuyHnZofLRvpLMtQlipjFKnmRO5L1P7wj/U1y8iUomJ7N
f0jAh0fiU3++BOSushaE5ftC6jogNvHDtk16FFPIjojYtFWBHdWbpz+4pIfBjbPO
1o1IdcJUqV5uyPQRF8xPgGCzwVmFvoqDr74j+eSKgA15BINFNHF95j9Ra7CgYc6V
lU1nrNTLQAiB6mOLVGZx+ZmhKuQlWYJINj0MTJEkPGMMvxxVRu9cXqlXOk3/BuYE
BK7ADErVjWv0TkEEL6Om+pyBQQ+5J+iEM6MosF8r1oNHe+sZ21VbGOXxunqIgHKY
9yFBqsUKnTKOhKN79NEdu4lDI+b9horAYfeRnmFPoo7hhYKRf40k8ck65ZDxX53q
0SKD3Ib+RLPlxVQZN/j6K+IlUs4M2roC/02NtIwX1rVIvA5l8V4bZSOnwXIc/Frz
NAgetrSxMTDy8WzeoCQcwhh5DnCoCl5Yd8Y7pTANhdFTo29FjUk+Y3wAeWDe4Svo
rvoUFUnqvnXvXgajjWxQKJn7mqmWdmCFmbRHarlnf+FLL74wSAXuNlR+vWZ9FqMt
Tns1FDGtjzDJipSpVV6n1+x8TfsDYqn0LEjnnyj1foVFk5UtzrCq5pYTW/jpwABh
3qAZbB4vN6IEz59j+cQ4XPQne6atchYy9HwaWoIQM4/bnUO7rHik2MFIqI7ASLcW
o0bT2vQM6eEoIHrHyp+GgViOy1whuqLt2ioRWUVnsZYXHEhKJLE4niPsykbejSUZ
PKVSKaxp+hle4yZS9pyEFEI+2JOatocsDAxUZT2PGey7BrAponUKZQIo3UYgwcn+
DmCS4ovq7I9zfGLQxfVaCD44fGbDx1GqpDW5Z/CvM26Xlsy3AmaufLYWvxi7dHPA
3pbzrFAeIuS58BVtir8TBarA/J6m/qa3fvpEvYXUMLcLIZLq0XoVuzN/8DwIh2Jb
Lw8UJygGE7VbNuWXrou7nn5M/FzpTxUegZnTirLKQl8ycWR3qmxctQmd8gvw8ERL
AFXjWP2T3Idr+SuuROhBm6JOBZGiFXrcS0uW2mbbodRZno3ZvjNvGLxrxFhItCYz
5dcEYWssxKIq/Rq5tNnkd9FeSxw1YyegL/1VlqAP0F8M7dznmzpCFV1/r8haljWe
LP2VfM/MX8AqnJVfzI5IAiYzH9ysTx94i0CZ9u6GahA0Puh9TVC2rtosAKeBLBHW
6zDVDFWUR3b0ML8jn4RTPgwq6xkSHclt0/5Em7j3/rZqMqDLSBA4spv1l5APqbcM
Mt7YdA99ouMw2mPKVrserAqUXgEKCB/Q5gKIT+F0Ov0prOkDlJlXbwIsxtSM6BF/
E64CW2IJpq93yL3F8SKQYIK4crTh9lybJ5gb6kc4zTVDfVX85jnVtRvTaQkyyiHm
NGhZaf2BeU42UPAy7wyoVO0I2cnkq6dPmqwDdotlD7SBHJzr1sdDDPxodOmVxKGC
hlZCgIQhviMorotaw0bR5YpuAnvvobVVyrJXDZ73HKpFeheJJLLs7qO8GXS+FOgL
/WWZTFfpG4XgQWgUgsHEW01IVfN4+tb3CtkvzEUoz8MSwMWlUm/qNhmyj/p2r+Ll
hdvRF0wb8DpknX9MRL+7id5hUV4c+169RE2ZserzBvY/TsyZt+7OwqcYGtaaUft3
Lehfitva09gEXyzFgHRLMXtskmEI3svyZB1gQ6t5P5TOcMybr8E4xdQO94etlbCv
7oZIX7YzZURC1EunoSkdeEUV3G/6MjU0Q2as4H2weVydz6fkHKu6pFaaDrV7D3z8
y8YUPZh+1Ce0mJ+4jFXaWeZHCX8/rAUGmt6mmuDrK4JSwdMh7uuHeLyzdIa1gdUn
qprouBgdJRWWQJoIkLjEabkVtGYoBQE5JgpTtmpjWwFsCobjPSgaHTck4UveXsup
8nIOJ6r5jQp65qkI0vrG02o+jmg3c55qk8xScZq/bQiYxiBppkMFm0spVTvnDdku
GZPJiinHbbTS5+wkZrV8pRcwIayvJtqtf9TwT/XlKvl75Suz1VX1Q+9YL7cqbbBo
osZaaw1np39bwxiBcQrM3kMlY7jqZ1l96lTULO2uOYSm+u6nYoVgiATKXIxdFCUZ
8N8NgrJtydfmczlKRaC0K28NNHKo5bY89ifXWTX7qAfkMYoLHWFTqaPoUY6IuS6M
4jbeb4VvUPXw/p6ROrP2f+x8PiKo3YNx8R9jb7p1aioF1cQNOX+9y1DRYhNArJ6G
93I3esp/IwY8xPrPewt0YV4ybzY7Wdi4d0lwKKHat6xEJeN3a3y4zBd1o80N0gxf
EobIaBgDCU91G172aSv6ZT824DfY4WcKrSe3Y1ZoVptsEfWck+twEa4s5RY7k1Vu
iH3wP3zZNhoV4SoK3dpNdps1ITg4Px/jqzROFfrQ03hn/Y+K2I6UlttyQW9sFR3l
SKTLM04TwiF60ELujS4Yj2rJgsUC21d0RFnM38hZjB2kC78ZPg4aKEiVnBCCA742
i+K5VJ87VgeyUMI9rLhzPHbf5KwNu31iOIVGXvegMuW3YJT9Q2wCJjG4nbkbjfki
Mj+GdhSgJ/sp0FWAhXXDUwH6jWqrV4erCr2lhxMVd3j1imeiKOCE9uJ0+LaCiUwE
VdnJTIIyngM9Lh2QaIFmIk4V9L1BT7FA5K72fAp3HlN7MADbWDkV8GpEFAEfwwD/
J0uhvN10Vkw21+9l1NpD/3/OZqLa9sb4ALdvvBTCafBMoalM2kOUyntGbsk7kkNK
a0ltm79LpZQHD84FZkoLIZkLP/z2+Kt7EfPRvMAk8DwVGowW9j2FQ200dG7Tglt2
8tVvLkqVNMPUwkDVKBHhEKgy+GvjJd+G7R5r2CRfZIcZJRZ6wSh0SpHuUeMkK6x2
TeWguq6bmNMlhpfPWJFsFt5UxGxSFojlFdZ545saHE57kT+i+QYHl9AgtUR8zhqN
cdGLAp34yHnC5sSsFSibZOLs0k27IsbLaNk0MG1kTCWFcWsERrgJGBc5SVMu9ZmY
nA3nrb6TdJAjeGjc7oXdTS3qxsPFYDY0lDUcuplg0TnpMXInl7RJ+T5/aNSRki/p
xJI+FX6cF70EaBAEDy7V9AZ6KcUJRZecAs5GRR+wEBR7LizVbgBgz9NV8rwGcS9c
k1za7cJdowviJz66Et65KxCBAswIhH5/vb6l7E7C3XaU97Di04w4fJ2FDZDgu21L
pg6XSZdvib/fihD6tW++zw9rFUwLwsdnydxb7HNa0zvmnIUiPhOysajMkgjYtaGm
frAQRro1ahBQHQm2qkWC6mVfgzeVSrMnVKpjFVBeWcKfaziIcPGpapGtsEsAmNpz
9d6cgE+gWTRHyFRSbBiBthTva5Hm8RjLsV3opoLnX2I77rB43PDrQeYnKRErGUfm
5o2ZPr0cMqC2FE1zuUyxUV5kYwFsLkYTlxF3yMz0RUrzlEW78S1OnBMrw0fzVy59
jtZKQQOYG6p3XNIel2MmNVHmcEm/IBNyAGjOtLiUh99U5m6nOhwVE6y6ZyQCR9+L
gL7RblKjqKbdWBgEEkGvO9x4x1GEekmCjVGBNtRp3aIQch3OgSux0iRN54L6N3ZC
2jXoCLjckb5slnPp7UwPEzRjX9xoFML04I4mqYDiLVwyqhmhvKNHZWqBWE3MkwsH
6ZIVmsVR6daz+LDJjiuO27EtwyWzGDO1SZgaDJdHxJ7+sJnTU3Ayus5v03+LK/bi
+Vcv788hodaE/M5M5ZKCliVwEN+O3vzmPtTpWkkk6dbjoTlNZdKuAun4hQGllEPc
JbBHDihP9n2pOBvGF/M6I+fvDyhSyOh2vSAmE9bwbXU1EQ+mlvSRCRilpc8Y4bWh
OF/VpskX2Z6b0SswGVF2fkd8JwGfzfXibusATmvH1Q7hqpf1sFxqRZGcf7y23x4Y
PePjXsZxXzO6V+FXCtlKTooqKw0AWq5lnVb/zz5zEaJzKBxAvl6hgmnS3Sjh44fB
N3nnSygCt9OStF2N92EYdVlT/lKOWTVteFSkqOaaNsM64DTeave0iOjcA0Id7hiP
ZfcVZva505f8O9l4NkfjeRqEcdpy7vQajATwFcvMiprVlcWwDWl1RcrF1CPeK/Ls
zXsrQo+Ii0sYeub2si7H5+80XfxldtNOhO6oo+FLMXExjfl/Eri1SBvIiGKWkltr
MIYDloLGMRrw15KuuI/fuuOQnGZVJzl3vhXrbPaDg6YWm2NHXZL+pFUaimBexSMm
FH0q8UQMYs5pS08TQuJoiRTx2s9hk38vyO1b+lxvXwyMcRWTxzBt63QZSraGQcDx
iU/pSuJcgXcJfHS6SE/q/17UwaUNE2p4IZ5q36B90jqI80obZvWDdzwf59Jh2/MV
KKIE0r7wByl/zKDvb0Ueo0cfaM0WOt4r8TB1btZUVVQxL6G9Aq/XrNLlRg1LY8bC
lL2HhoYSKMkBqEzdQdrfl69lOtKfrgpxm+nactCHHkJOPjra+wLWgY8ILSdrX4TP
batoXB94pVGV4Tpz2M3rhsl+zdnYQdbnXemCOosRY4bjb/7UNnza7Myu/TnDRd24
QIYLwS1xDlQG2CuNCHi+KPkDUH3a7XFWWqrYUt76G4xLN7oKwXDo3/S3zedXJ4HA
Fw/RFQnvZxUCfI2tpZn3I+0ruPdWLto/apr6khACUu5ks6urL/MFt09OrMG2x9Jb
YktBerbfk5GRGWj9I08avTxOiQMbgYGHa7Sjj8DuzqfbUrn8REZG8NG/fOVrm2SH
tiRmuEAqya3jcbf1sl4xKBL6ygOG6gZOIcZQgfKvDBkAafIIzQuTB7+Ys4Smfmp1
e3m0n/XI3ejQkix8j/7WSKWd1gMhb/++7V33p9g3oFIxwKvFxW6KE6p51FQgDUdG
J1jymqyYbJo3il02WkkkF9jbdK32DGSKKmsgyiEOFNT5dmGRLhgnPg2kRc23nxIw
95DyuyfmYKopjx66q2Q5AYujLcKA130Q/ENN/Z49HKcRgEWteg94xI9zoN+22ZCq
YLaU79RVnCf0UaZ38JDwESuquXXujxyfhJ3P8XKt0n/RdqfsDUmLSU+gEr2j3cwW
Gb4raY83j00YmRRiTK3ZJ7lNWN6x9EN7OdFdWknkDqM36TZNvuKR46yfoLVnwYhe
rdUhf/yFvsWoMXKnBLkpVrcTvSHi447owSHrt/fs8mVUUa28QYxHk3YG4EI1eM1j
aoQXEnsxAnTNgmOrpIByRKMj9nNkg0WWY5HNXi5DjfY7gmikDq+S9I7tNtVsdUl0
dfMiXGpwtSMxbVL+W7cFyNOf+RYVIWdGz6FmBR53lnPkYcphNNHab7sId6ZqEcl/
R2WndykeEFIM+JsJjF48l0rdIPYOW9WK4nOu/MxbAgtowGhC5PglVr/ojfM4a/DI
rglBYhWAAecIpaBnsjIf2y1hjlPZiFwJrP2x2wBJRvUmbzZDflsHTK1dbpP+dt00
oDH9KozERFz11vwYYxrV55xz7ZRj5uJgJVZf5V0VCs88pxEBTgQ06GlqTDf4ltMk
Iq8+5TBEnWRZDtoibac7xhGZT9io2Pok8LsMOhTCoGnHzu5lvApPDv/hd2ThZ9Zr
L9qX7BvR78SNJ+hYIAdEQw8YfgjSAXxTrj65WQGStMjFxVdV0dgfrWe+Xysoc2cd
6HecDSP3S5W6neqBYIJzKibQz9KVUtJIC9LiCKurHKN09KBCO+5iF4ELjcJ+AN5X
PY0SylI5d5JigPGHsmAXaT4XvWFE0PGqDF41JsGwZacnG96zeFlhgJHIoakCnbXr
IMZa2di2FB4WngUz3rJKJcuUggZ4s2V1XK7LR3Dyo+/cQ8P5OQ4A6AabrUiCXblz
gN62Y+hXQxBt0DYGbZSPhQ017o+FV9sdWsetTsIbRc0P+A24Vjj4+NcoV6NPzG+H
n3IBBJhm6PjPNNtnag8rIdfDNBcTyhZsq5cbvrBEdHjvfssfTfXp9JdrmhcxhTQD
VMM95OibLYVSn3nZPYKRLPh7vaw/hfxho7nr0+LlUjDs022259/E7Nn027lR7yfr
2KnzwLQ7Vjp0XTlZXdh0AQlLg4cJMhASAN2BlnclbPli+TpwtBVhGpxyhes1B5pk
+lzmgMV+YB4NZg8wTqosVTaO/WpcO6Hb4ltW+dq6D0HeNmqZI8BBoNzgbAL7LJBR
pF7TDSZ2TzFx/Ry9/6GRCbNmiApb349+HiE5ERFAAu7+7G8Z4Yp3hQg7gWQcgxPu
DR3xM762BwfdNQ/byb7gLgeJnEWfw4797lAG4clTFc2bUcGLSrf9OY9z+cNGbE9M
wKruY0bRh/T4tQ5vbWF0m1jxqxH85CqMS5ylQeJ7kjzsS6ABG5k5HmDxkdUBqWnY
Bovm3c6MPz4lszuLDTuwgqNmYpOjUPg/BX8JKPQTNVa89e7bHemAoLlflwLomFOY
jUAXLDNwAJ9zIXa3BX9GpYUXSq8Shf6qGzr4qGdzqFj48j5iLzOv1WYDyZZ7uCUA
MeBpiWYIotZkNXWO8kLpeQ+aVOqEP4t1HxpVTguvw617tr4IC+8hydji0LDf/0s1
BUnXP29Q2gBwtkGWyBpkby6wWWfG3eX0leIqrEdyyiU4HIUaADydTXzb/Oh0/8iz
z3VMJ3/JSFd+lIrF53r3VSylwZ9SoPb1BU8cj3iFpsnt9LN4cI6BesgOsVLqAkQ2
C5NbNfvtzQNCgZDUmtklOQgn6giElSyX91NAdvby3ZpRhW/Ftr2mivIQMJlTEEsA
Ndi9wQVblrCoTUbiR+cWqU6lO36XjppDE6xzEYaY3+SmITcKs8qBBs2xKGQVKAmQ
uf0rk6FSAUhZft0CTNd71oGFT5VLRJuA2gqMkMKNhRxrpcZyJTF9GmgmjzQEW8f/
9TGPQpF+doFm0OwBrD2dIdKqUMiKAodnT4I7Mh658jgOyFuo35jeVEbS6Y6IDywE
AitIwE9gIg4q9ob/CuGj5prDNaJ28ramlriFnxx+wRhqaxk42kCSY2+/1yhqEQwW
Nq0SRRqkct7zu0pPWsvf563IQ6Q3R1PSll5Y5J8zG03ehAt/lWKJyTomVvOq5p3a
cg7SHcJMQ7DIoiP+1ktg1nj5qAXxr43XIu8JmM4V9hrPv9bUw3iT21SxXOaE93aP
cqENEsrcITX9hE3a06uJd3uY0em03Uby25GV53ckIXX0wILLz1tQIhUk5aQ2njWa
5jJKvP8byMePGXpinlVKzEeTcsgfM7G83jxSfKMOlfaDOV6ZWgQUdRVLAOcXg9qh
jW/SIxzXFPU7Rh87cvV60baRe1SwWI2EuBL4lIgOjjV3JfiXpYMal3Q1v2F3J8BW
3vwHyFduxfTVhIgwLdSbc8qJ+lpMTZZTBOYR+PZxwaTgldQgmH3LFq17xJvJ0RZ6
AN27PQhVHMv/c9oLN0pc7vUtVexFH5ycCfQ0iZUMobormyAG+FA8b2qYRjBZGgUt
FL79/Wwy1HytH5+SdLzL0CBmcMLdBcNLYH6WjBQXlicN4GkV5RiODNwEH9pH779z
jquxLgoZ7qN4tpvlDCg3swC/aGDnZzKTqoVcuhJGEPvOt2hsN5SNXmnsC85nEB9K
BYN6aswN9wpHEbFM3f0KA0y0fg/30hHEjxY0UzYNku4C4AmihuxTzNq125l3FzBu
h3k43R9rcIAUNr/+WUrLmNYXu05hKD6MfN4UGYO8z7kls/28LCjrNyGIcLS4t3kD
3rLYanrjk/uLPH1FfJjv6b/QLF0pL1qSahZaJWQYbVgsWTjYc1WvBoXsqwxcgIWh
yqTj0Rt68qwZFBLBLW/oIWI5ZtwYQblkG/sDhIR+buv8TE8Se675gYEjYA1hk6cy
yLiSWoQfCyQnAVnU0tf4yQhfhbGKsmbDEb4c/6c+m5If9umaEBO/vkee/Tou7W/L
LNQjYAai5DhYu7UHkzRAboFsZOjP+Ms4kISQIeHRkrqflxKNAtCTFJNB+Ha7i7fp
MGP7yOWJEJ3WQcAufyr8wT3CThYXE2DFIOW/7QvScpBdPbYzgeC5vdt9nZIR5pE3
DIvHEKnOOOvrLWpjrFJSry7CTDRoysNuE/c90XDDreJ22yWISM0HJZuhq9IgbhHD
i+VgMSRHezGlJT5DKmPEHnqjBGQR2fnIkYycGYXtVgpGwwPn7hwDKTbHGMunqCGA
WLYTGxgvM4ckUKSNGXQpoklvA4YxHr332j3l1uFgvgSx/UnmwVJiFxcpMiXj/99u
vWetIVI2XJOahgFeirTKXu8CgNtrCjSeMUXW8YbqXHBVO/O+nofMpT4Nq0wBkvQ8
m7hb2OFOQ4I+dbBPOa84/BaZKhI5Fa7Z3qqMW8ISXhwvqndJ/eWA7JYjBe/2QvEN
SeE105IG/wIYanJFcIT4ZoArv6wjzcUoh1QT/aE2wG7RJUFn3gJFn8sqpFktY25T
y16zWA59Ybw6MrUDbdGeZadOni/fWZBkAn9zyOudsbM0sVnYCkrH6Ibo78q62mw8
rDzp5jfsg4uNRtExaeDo70pC+C98ssZ0LS4xbv1Ynk1e0Zo8rjnxq+X/Xh7HC2QZ
5tQ48m+D5mcrSWddjd2n4rl9qTKj6q9ObckR1dMR3hfcYGEGKwOaasm8N5mimmwE
0eQnzzP8i9rMBcQUlvJkxIKFBWS6Y4j3FGiTnvTuo7o7wJbAL+H/Q3eVVFp1fo05
/x1qgzHLKGMfpyXhe4AqfExBSg0A5GwCANAHWHGW+wLWmdtFKqssudGGf6pkDYWP
zE4zk5hD4ZNNAch8e3MmnHp3Hyj/a/Ye/2IJlGfkJn/zP2CVWTO3u7NJq7ybNecw
ucJk0IMQrj/4rOSQumUEC3VjmYiPsSWwuSa/QdpmZMXgqRN76EYN5uzTqJQ8Ceo9
7vcU0L9ixD1U+j7DioM4ND4fcqVatEChVx6RwqE/MgQm7PHtYABX2JRSjCQ2jTsk
jrXzZklXpZMq4nQzgcK1FWIB+Jx02bDQPUfAjKC41jKZl7l2mJu3lPco1sZnFvrL
Qflo3dNX5+U98NOy5aAcJDa8Cqg7gZ3zvbO54ihdkGKTRlOHpuBbVYUuFuotT1y7
Fsc+mfPOBBm2vqzWt29afonbb0OgYQVFGLcsaAAIhKUPrVFZrOOrTBNbkCodq2om
+fi9tPteKOnhdgaOzSoFuJKt1XrRDAm4rTW93fHiFUQPCT6DL22r3eYa4U59M4Wn
zq7PMyLJMqhjqp0qJL4k1LhhUUq061+gRlGuNjMHAhOSWkhLFThodrc5o3ZW11+1
vnpmdSuYKqRPGM1m0wxPYNwpwwsMovGqbasp5iGeURgHGs0+xX7HSliQkE1sixzJ
MFEdn5t0M4g4RQThEoud9rOjDIBHE/laRPe8/i6hrD1LV6I0JErEdrj+imq2JBJI
SyBZCfAMptuEB0xc9Nytm+DEDuYT7Buv3uV/1v9QVmXhNb28Vt+YilUqc6ZfNjUu
W0eqwAPN58xQ4VLIZK/TooL7Jp7Qvv5Aor9NPvjyj18GfCBau8Ym+n4+u6UwaikT
TF3iYsAkT1YpY/DrUBzRA4BiHar1aD5/5i1ZGilLtr48bxz6i3udfxZhyasBGFxX
LvvoN7x4gUsF0/AVqNgxAL7xWwX6t3DT4r5OR/MwJ5FE+LWrgrmCK2zun8TW4TH6
iyt+pMFzrvoBos+8/FLBN230ruNIpALLWblVFjzZBQS645cE7i+rND+EPvhYu9C/
IAPLAvmlidB3xxW6dR2Wn+e5aSjutnanuJoOZJ+WBr6QvnMMFLNXtQMZSdf2D6nI
5dyEi3QrOYyPz5lm002csXw0y4OA4GQ/bGGNTKeZu5gSKFXRG01mWB4iJl+hDKlU
UJFOoza6QUk77HNOfU1boxnQLdTS9Tl1i+NRtll3fry9U8uIIrce7rDPjrWb7d9I
OwGKFTYTuEWxVdcbQf0xiraxo0WyRfKFuFu/eLSt7tkx12wq/6COqiUJQA2PxXs+
RulT6fk2lOh8YNRwcdFkxFKWQCXGc9VWy6tha4QY+J6H+rBaSwNwSApb1MR72SvN
erotE1tw09v29BcKE1AfABKOEOeFUVL8u3tFGE2W6oxBQWZI6ehLDoLNE91dfcF7
n6FfO2ghlS/HYdZiLADLPKPJBJSPY0fscDXBZf2DVBtMBA2TjVtQEF7b6mTWaDmT
uEtbkbdZq8pxbOs2U+iCPpab19yVm23RiYRoPQwKkAI++sIqClHWYJODRIgu91xk
Y/S7chr7/drflfSjgoQfVgePYk0ppL9J2RueRR/eE5hZVFP/VXEMZqZnS2Dg6D8v
kklL7i3qMoYFSK9bGmgPuW7pTxyODtQ4vpfDIksD+ogvA96MRCfUZrvWrlXaqAQL
OYoaNgOd7P+X/w/SqXsVcGyMJt1cIkp2OLhTFzRUzBadEOLJJsZUNdLD3fmiuODt
3hfdIsZ1DfgwzTgcSCysVecZ4fijjurhfvxd2gf/vJ0F7Yix3mfS3sK1e6qE8pii
NpD7NkGBkXF6aOhwTTT1pKC/x4LOiLvhRjrWdlq6b/IdSteqSRWGiyWzqCmiYVK9
YfceK4iWnOGFOX7Qd4ebbLtRsnCnmHjpqfQL0N+PsiuUo7PEvvKyKK9z+dqtyfQo
RovuHrv7EXcP7kX5GsbqnQSI9HP5aJNNHNtX05qU2TWVnGAUZastqsxmhIAqtTDP
MvkFSo4tJA9Sd4o0C3wCZmhU0Bb2fowxSSp3mhrui72zO7a1Eh9mkQFw6aE3xq6x
aKgZKKGSh/79X+m54MarMPC2SwpI6sfRcpmj3gqS9Sapn73AzKOYF7HoWe7v0jUJ
0eRYIz+jFfkEj3bSpwME9YEDJchSUvtv5KE1Ni8IYcvrj1cWHTC+Yhe/o3T7/O9/
hK47QpTOvRJqH8iNMI9awciViAVYGl9QZtNsRl6AD33QfDCdhF8haPOVUoq/F1gE
3RACA6gVK3m/NeiGyc9y3vZiNwpZ2Ieu2cjtlM8alQusx3aLm9LS06tWcpFqAW8p
aMKZJ5buRQb36jbVtGa838WqW683hlcNAmO0DGRRFv9ftRq+4gzQKwA9tFJkkzGj
Apw5nOYK+HaGlYcgLlBx8qumdm4cRAU269c5Ump0KQccDTd1HSdEv5+RF7O4Fzof
Yn77Q2COkNNNq0muHtcbg2g86R7X5snZpEE7Ig+6SsjiLarP1Dw2sgFQt3uejYdb
N0IDj1pqNcifdUGKEwq4P20Dfcqsmq0okGNnSs+uqL89uD79VeaLiwYsHVQmch5a
406oOKmSYIegprNyU86oyeDfXEFIJnVRGOBGbWNYd19PuDw2rupXI+a5vRdiuRNB
JhHpIJUGQpQ5q+LrRY0kcAN34aJImfivI0oTDWDU7lcHdvBLikRkKBDR2jacvT0T
UAfegjObwshTZJfd+5R/A2oqSLfaaNpYM6i9Pj+RYkfcxRMgOefq5bkZE2TW29J3
imvg81Q54IDROPzwXgC9+a2tbneN0Dy0fgPI3GO3qQ2J6/ZyfvEbcp+gBozMaGlB
oRARV6vxkUvrBOTnAkOnck6crxT9f8kvjOU9rKskwH74eDvvI99vKpbaPi/0mEs0
mykA5m8ZpfcTfF6g3QTOsFMgBfHRKRu94OUmlikXcx0pCSipGeTd4XzaLm8LGZ1P
eDVFOJuruRBGRuCP2VREX9B7uXFT/Pd/lO+SUa7KwD647Wi9O31tUBHEa1RzEcRb
U1dKU0HtCx9Qu62q95z/ark+h/rDRGjox8HfIa9hl9LdBAeVINbSVaLiUiGEYNmc
NhYZ1lTw0VdiD8h5rHIPx5Mptpqnw9bANpLLNCxWp5r7FvLjm04Jkd+N6RqPau7u
NItsPl/yi9EYKz0TZoIETVr8bkCuTqKV8iWUF4f1oqvAP9SjjPQ4NFNNSp/xvluq
YfVS3oW/fXv0aIsVKWHzNxHzpWO63gimSZSql2a17LbEz/ZHVs5lmmWkGXhT6LAd
z0TZ4Zi3nLnbzB5K/+ER6ZaZ38E21dv38E7OWx1HgdkEbP7vXu7nMI7KN4YVFRKu
J4nWvNqN/rRlbYHQOsbPzHVePZcJU/eJQbbslDDJtHloxa4/TfM9zy+xao4haOom
3tEYXF4Z1hXfcAsYmbosRbuVlDrKZKioA5JeTffdRNJXaaCDmt0mnUJJcNd8OLVf
QhYSvZ/ye1slfeVdVyIpfKOCRCNHv+F/NT2Vi0fm5aJcJ+HdQx7cQyQX25vR+j+O
3+488WgLz75uH+jl+xlf25K0T74PMhxOAYgL2om8s1c1DObV7qriJNz7mDnxSuAI
tis+RePtQUcAo54AjNv/vlxjztrLGu4i1qM0JoypBZeBTgPmVDEVzw65cJfbZ2y6
4hAdqPDO3fY9OP6hkLWonRj4mAwcPOAtgvqtRwhnj3tjzgISJoqixE35Q0oOqnjp
mcqKciYCNkfP9z7OX23BrAvieoLb0+Q0TfDuJ9UP8b4Qw8vL0hVmTQPJlxxMAkkv
ZgUciY3xOEir3Zx7NQkZVKDKwc8Ktopyp/FbL0g255Y/buW0RW45PYwD+GQF/x96
Nyz8naQhiTeyU2W6j+PdxpfNiz+SvqxT8lZGBf3MyOlo6Wr98UG/05Ufm/p6YUC7
o1Ig801YMMDeQTAStvXal96Pszna2XqmD/9h7SK3TdbkPhBxK7pJqe+uCBdG9aVQ
NUZY9HceTcdgQeIrJtlFgGpT+tGdbXfDYbYxSjH9JH3G90+3+uvzF1co9oV12x8N
cc9WVg2OaREq4127vlgQXOjvqCULuITY4YbMs9TOT3CaVnnHFnYA0WNZeEwluhFP
/Zz/9Eq4V5SzB14FozMF0J3d6hZF25dnSG2WytkKWnhe/8ZNlhGt2XvtRIv6qV+4
omamcs72bp0Qu2D7Bn8vDKyzlLcvjmrmWqUYAGyrJz5xPV5Z3gZ5NENDcoeebCla
o22IE8NvsbZ0oX5jRQicuhDzJR3TeCqMTRux6yqGsbyILEcGR9kTQo+cACmAOC+T
/Tn3otuDMvXKb1jxkHIerdAJQfQHMFrJij335Mbjk0buCTBFmOQwtBz7CAkFyAb0
97hjqHJhtvsSVWCoye0Y4Fb2oojiZtfs5euQgxc++mewTzRC8NnqVm0aHzJEwhg6
bziEs/5XrV327uv6kWGXfmo/ypzItD5fm0AuvNtpljetKcntLpepIfk47xP0VWc+
Yx8xcKyoEHMj51pkJ33NvRfObs2gL9+ndWFv2McoKsH0Fa29uPfCYR1yAy0pOVv9
LgrpzV/1BROiyZ5tbbtV09wLToG3YcPxe4hAqwt6N3+wvHjAGRRerwi84dDKtODA
2qi26aO1NBQhSGzHGDroh+fc6V4r3u6Oo8Bsh1uETAcvQF1sTPoDcOtuTeYxo2NK
sz2J8QAUEYNgW+YIFMumc17jRzHKKoXwSW7Cghs+QF0VOXnR0H86pG0Rh7KlYM/Z
+2s7BIVAmj9To1tWhP4QsFMXeXxBl76gDfvRoZCxwvaW9/XDNVog+R3WuSdNG0cP
NyXf0zGAYgMWdnOnUiCy4EInucLeyOTLlceEzH2rxsuGsd59gZmNOxsoSCAjdORk
9uKiAlNNRYCVwmnfscdsg/7NG5HzzOz+MT2E18ofHDhA83vkwKpIf7WDSpKfrn3x
l2tfWRkQsnGzGEUaxrBh8n5PfqhvclOBgcZQ7jvtY63UCbcP7VpWO2VtJ6NLCEi7
SHt/DDOUADDtGO+ZQU2M7Foy6OyrKsqhqFycX56bRydSZTXOoR5JxhGo1IdGUN/b
gdqeghdTfOPX01mJX6Q8BhaO/HugKJNImV3XQ5HArkqHKeazOY/7ZoC2ZG0ah4nZ
axt6PEDFWuwWZ/m7AAMqB2YTXlOTHUJXWd2jvxcHsYQ+17aXFP0nbm0Gu1zhahw8
OCijbURDQVkAlMc9MknbrG58+QDvXvfwmOTuqA1YUCMI/8BkRWNboQZYdYojBDHW
WT2F9O+UPzkdYeWRP74ce3pfqIT58Fmym+WfpMnKlQBKVC0MViW5uSvrucH9uGC6
Et/s5OjAgqo/Awp5IVjPCVHI3mLGGGoze79b+8s0HttG/yJTTkavBQdTHAaU774W
bEHOYGPCaHhQGHLGnyabBeGFvaOREWyo1HeKUXBSYUqs9dbpWQbiR9kP5VrYN3vm
Pkv8z/sUnnXrAmz0ldJhjJ/Fs7bNIS4vVNfo26JDE3Pyy8oxq51sJIDBpG9Hec9H
YQjyizOA7+AZmESLIcS/FItgLhOvvIpBIQ35vmyqh7VpiVs5+XSEtH8ifGQTPkm+
+GsFfnh1SHloVyVgHXO9zIo1JIe/mCji+brp+EZt529mrtEh9B1AUsvDz/mCnREu
Ail3i4l5NdsurFmkhTBW+21dJt/tNk2Bc7h3Rc2sY5n4CybRW2jzQBmg0j7IIyPJ
w+DmaiTvtcqFX+i+frNsqbn2szUnWRx+ENThAqTr0Ec6tHdhwcENEhJNTFTvItjG
NooORlM0WYjWQi9utRg+QCp60PTQPsB5HpqQUnROTIq/316dQCfEX+0hPf4A9zsG
I0lLm2JRNA0X/ZYwv3e8dqOGbAIrvVxbzRDVP+Vi1LAWGpxf/hDjv5pljZfqTja5
xJvptslYd3h4v539N4cMs+VqOFIYxcw07WgQu1rG/qer/2TbIA1enYaUNCfVocu4
i7fkc3QrT24sqKnDJiRG1IF2rsaGW/H60rSCCn9AkiMF1EzKsYyb1BfXX1/zupR1
F1RzvLvue5YoqgNULCl6r1xzdyWUGtERW0SfMTLa7UumrlhBxhDGGCe2NHN7T/CL
nWEYBhxWRylMhKRAB0btZxWEC4TBaXH7Oa2ktcKqWfqQDVCfw42d84r+rzaQvTQx
u0AG62C3cT/s3gxzKfzDIz9cM2J9o3a3JZYAKmmYxtIWJ3H0V0RWNDjr/M3a+DuY
GHt45EttI0+IF8VuCVgFoSXSi0Ha+dvmOcTegXLaTngKxGwHayKUwgXDFLfvEBnk
228QrhSbbV8OYPoOxB3ApHEL/JwLlFQTFKvm7OmKueQQhM4k+MPvemNBUTRBwWKA
u55Z0N/87/zNim84X0eJJBsCWoVnEzTKkIaboQoar1aN0rqJ77bzBRRorCPTZKWu
/KtuD+h+u9vcpJokwCC+dSUdZs6nuaavrcyIEcwd3rk737WHD8Jtb9X+nJzq4LQy
39JuwCEHlDNZnws2G0xz80T2v/WxvZE31YPzfZCqntJxu1vOl2qRyUjZZgGoQqar
2m1BXhS/zRwN4uHuXASHrcIdcYVR/o3MBDrQEbtA3KQqgfqtZqMSX2F2gut+PoHP
Y5dVcrtpxOmjpHXLwodVVReJu0xOcfSSJENtX6t03/ZqOQW/nfFw+bJ6A1MPnq0w
i2/U6F9UYLETVZn5Mn6VSZw4NwfhqZ4ldXjzja4MpctejAwGx3SMWRDPYx7pc85S
cvfVsevElOTrv5bZboE+YWHEZLx/kLz5m/aixLzy71CTJk1+jp3uX5J4HRuiP8jj
oJkFlrnX0OyfQF9VRdRuQJIXgsxcWa2juR9sCxkc5yhRT67CAuB4icSbrCOm/ZDa
u9dIfLDDRShHvSjnMaEzAHYxz4mSMVzDGb8nG45UlkZ92Za3Ci5b0siLt2mSqWwF
IkUTzaMlhPyitFdf9ouvHdNYDb3pl2HrYpHoVKyhIhjLYA3asrRjefXTa8zD1BRG
ZR1Aa/mxL0/0ewolzJsBVjBfSaMWBZ2rl435eHkczBTmzhDpUszbjZvP138pW1y9
g+QbG4SX+yh44lFh7VGcco9Bv/dZ/EmtBcBljT6gNkANEIFtc3ZRIBxpUJgEbFMw
nH3hAdFt6j3ceE6M27HtI7lVzBKuvfyjaEKwL1NaZ8sqqGUWUDnuDZcnqgNSYxWn
bdal6atbSLw69V/ZXlFwPOWqFWucdlD8byc7qnA8pn+1jrFYR0JQ47SUoNBi9EKG
08WVbfyc9RkUqj+or+UxxbC5JL6StA+X0EVVJBShwtpjMEVVOy6dkiyhTLUmjeZB
OHdPHWXC6e1qXqvupn9msAnlwFTSzRivg1LUtnrL/7Z+flHI8Pfd1I57UOndE78f
LqjfEKY6P32z4Y/9w7bQ8lWLFyNZG3h9b3q0rJjzCF01xC4CiQUr6QTaeW9eyvS9
5OnjfqSVFCryHo/OjLzPe1EAWknGSiRuq3UEWHUFi/1Wss7Etz2scx+aLZAFLg6q
n64o11D1Rq1TgCZX52R91foQ2q3HplpRyeMeJE3VrkOJXkJttatQ+P2/f45D6OOF
EH5QiC4xuFnF073Bk+NALA948CLRgMqKOat6I7c/axi5jS7F04coLt9RwKt9HMi9
wtN+18acxhNDR+QuDchCmux35bQI27aPJHMLvrvFxrbMQB9yrNHNxqf0RKSZq+Jt
E/rJMic6mgtY8h32UxQGPB6vWVSL2LR5EwM3/OXGg2QphMJBQxptLLR3W04p54Ca
e1bJjdi6YEFpq600KAe5XzNjUH4SHnKGElavvczMgoGNHA7goBvgvFxaTp28OCnJ
eH3Ok9CGhKWMVXqj6KDbsgOWA8C6E3+gZ/79xDNj15ipcCPhPCY0pKus9FJQWG/W
5HnXttD/nvvt4+kpgzl/DWX7LqJtrfMJ154DxmGO0RbVsygywuH4rDjSa01Of/oS
RP59vDp5Jc7hcuYeLxuGobpJubJ5ohIFW2NlHFBPvObn+af7rc33WEnhPRbq5aWQ
xxx+bcBGKaHNGfU8OOwmwbgo2IQ+mrvhzlkvQznwSzYsvTntRiwTVOZJL6IiYJrn
akftqYnpL8EeEQMtNqABoArSnedhVJ8EAZIR5kjmXExCKdmzjNeKIiZpxvEBAzL+
xTiXpFCwtG+qwq6xyB9Sf+OkKTDsDzApVbuxfrb4nZ6/6aWhrBTn8ZiyWYf5E1Xw
Tjw9F8oMcmEnAqowjM+qKzi0XqC+Fko0DEfcV5nWbDgqV0GxIU4dmzWaqJG1UJbJ
WEuAZAutUVPWsVSFaUYGOG1/kN+djfdFbhxcwse/5+0eT7lF+yOC78zww7csfgR1
VW9JDCMMCcT2XFHzmTgCZ8ZHE0CIswWVQ0BIbfYLFnL5iI/Xu6PKnNnQrZr1emiV
vc3l1xVEJyC1R2GbjKt7yzClo0mRZXV5GJZfBd5BmhVPPNQ0x/TLq465gw9oiEn9
spMCYeXA+09au08h7HLm7vU7ojiK4paURosRcQGYVQgn76kXYb5ARvb+GvnDXxlI
8ndffYhrCuznbXSmTuqaFGmE3NmxaWcFw19Zs/cfQTN+eI+Pcg3FNxnhddgNR8Jm
yNXFsnxxw0g0NPMmO7otAoMsM9VodCqSb0XQNDxITk+BEFxKXD7n99LmtoMC6mf/
UyqbyvMhsR61euyyNxGvE0qJcmBq0QiKjaBeaVepdi7DCqI247+42qzcsYA3qFyx
jiDLxA71f1mSFVQerZ9MqLRjXZvD3xCW591Rgtij9mhrjNbjwKKdzwIxwkgh4FV/
LjV9bV6SKKmTU6JVXH94cnQuPLWADB7Hb6RpiqwHVobulpBKQOzSsUIqRHKQJhgj
EizvcRk34UphBE3DcY2qpTBLWcUy4NoEtwrSe4ucMLbqFJFhzOKZlizJEiunWSoe
jQNQLggf+NLAJoFyV7saGwKQkLezme/4jfJTK2clpSFjODZ4Xih3uAxZ9K7gbKVR
sB/pMZt3IEQZnmuiMR/HD9he8c6v9QdKSHPtKuBv1zojs3O/bnCCh/Ew7w4H6Wi0
iV3v+leTwb+eeswFrDoZdjZQiY1WjQIH9guH2UWvbp0XKascJ8hTNfV9XmVTe1w7
mxS0pCJ2o9doWcW25aFVPeQr+dAHdNNaW2lW9+CbPps/tJDnNGlO3/BwrMFppXBC
CWAIbFdIWn+LFI9fU5aXt9X0+bQLKk/HLmrTkNGL/75iyPt+LvlHrYWPwfKmMpvr
UYGzRYO91coZIWc6hSDfdgkHDgrAP0hRuqmSlGpd1fwF/04oRlLr8lvz2LXcXcH3
O3Zs+OWr4EpuYkY6XLRE4Qt66YjLjOddIDYRfZ61hMnNmhAhlNrmamagHnRgwiKP
q+m5arVxC91mvHrifFeQKTuDXP+50KfK62WUD0fRq7YPoVdVtKQQakNJnaXzHIqx
iWtkgsBdCaLGJIWGh32VKC7u0HyWVPM44ltDflslhhr5yrA9ab3WgezcSoXPEEYW
gaULoCAXSY22yd9DgNM9ykn+1yO3V7WW3FF574oJilUokq7qS6XVPycmezaG6VgV
WnU9OQ5KfnRK4QLqo7DReQZNiUaZDUOo1CHbca2TKgB7AiQEacp9B80savtYWv0P
j8CIewHP0QlVScVtlImWYn7MD8X1vcvHC5tRKditvZF3NmvrYUs66RDLzejmlDq2
wnXjcgwGB8cfH2arFHSLC5JxdLhwevDdR4AmntMtMg5srYYjht92kT2vOTWYNp59
XxhXzc0llh52f9OwMNdOkNPh9gP4aWt5RsZFEdS4OsX9TR0UvzbW4VsuktsOj+1G
0LyEr4TBKJpFh8OyYlbLTJ3fLdJQeWhgxJXk9DiQL5zyKAw+q5ANFygweERDEaYd
mdHUikkAE1CvGiWN7r9rYs0CccaG/JTeF0+CqfifyU0O4S+MpO1D302ZJZWjEZVJ
AezCEBCSfUuhw3/1MalefO91MSIHio8VVHv5VAxeJAvDRw5gswdaNN++Uxwq1KQc
duTuMcwkTdL+hdDXO8wYSEJN+AIKR0cvS8LxgkFdWrxz5VPG6zLOTLG/hEvs+dRp
i6+smQVB9a+85aI7HcQR1D5cN33vR3EFPWVQlbA4zx1LQClHcd6NWK6/C44VlJ55
gNUwlZ+93fdp/CqZGoS6bQjVbXXl/bkx1qjGSRVjJlj6MuNkVZKL79LLAjkVMN0w
AYjtiu0KRQNqxuDNE+NFusoz/WPGUmTLnIjcDNI9DDVsnVgjYuGA5MFReu2qdwaF
6kVTM/bKApU2vZ+/pjCSJT6YD0kNmfb6D0iD+oxCofEIOYJFkc3SOXpaiygeZPJt
u2jJRGcE6rHpnsulRtQt/i/AwValsJp4THkmcDS+Cq8AXyCxH2al8X6VrOrLlNQu
9BwHI/y6dBpMNnaQEuAGGLGNsZO5fVGGQj78knQsqpUrgjRSfLmZF+xay6WW82gk
2+o5P9xgxf6dzfy+FriE1MFgLTLPuHOSt56bMVP5nShFPfOl6aj26sUjsrtRZqAV
OQ+SL+ZSj446KjVmwUHHZqKMXOtw9lMsIeKisOG2S5xH74xCm+2Eq95s3x/X1RK4
RBG19KDgJqsVfejBXQZOOOaDFjGy8pdDROvM9jnETpnmRzH6Uo95HSxN80vbApeI
Nf8yapo+xRVitNonihAzSqObVGfqOYNcuQsLP5U477w2FKX7DY+COOqYgCQIBSsq
4C3sZ7KJ0JcwCcxzlNpXf9cq8QdNR0n/fGlbcdXggp+mny0MvVQR61YVnDHv5Rwx
b/VEeSBgyrvpz0gaWbgKkhdFHC7frrtUdJInMQqjj6nI5Iuc4PfBuceK6YqVJDTx
yYD3/LqNSbvS6mIKkizDB659V9nbS9y3JLJDkP5lAkzudJ7YvoRD4VUF7szyIV7e
KxvwqOwc76TD9Whoy6W9pU690Zs1cLVCNTE9JleNfFVrtMNf8JL+RtVbKMTw8YET
VTmNb1vrgReOw0UqsePGvcWuUbejpC1fhOHY74SCgY/wdqGruWdYjOl0+6s2HiKo
T178Ac0XBKaKc+lrlKaqaPknaCyvCR78z8CE1sQWlRI65fu7bMBi0MLX4LthpAXx
lHoC3hyIVgHy9vB/ciyzWXoqzWLhW2UCUfALDSKmc2CFGY/jcNqF3E93Q+vYRes8
07uTws/FSQ7r6DUaqcvm2EZlW95fweERB/dKufFqLiNk6g5EonRAcBV0dPFC+h5Q
ftYy1PS6hgnHsDGNJ2FlFH0kFsBTB7t6SY1uuxDySzn5xpQAOfxOsXVdndsmP7Q4
pd21SuGFak2gPArVC6uAeGdwiTBDJ0aLCn1EIDVURFpdrBxqcpIgysCLBdGdxrat
uA9/2ucsOu279lCGWxcNdGRlCUtj9aZRCyjXT8/KdtEMDmI+9V9DnsiF/K+hLgyj
UhHmJOhKKR87w+HinoRXx0xAcEwQ1wSRazDdZUyNLtzQT6Ylvxv6j7F/CH42sdE1
IdtCKcDtMlYrTJjUt4HtHZbN76q6ZaRdObE6LTupjUgpKMw8jb+JiloAm+GigcKd
LH+SVaPRbcB+Avmmng+z+i0ahabvLw/wm2l21VveoqC+Alis4lOZoXsyW3grJHiU
OfRxZhhqQGfti8Wm2L1y/vIrlRV0qVUXtOZ+u/zs4wkKZjP8r4Dto5eWIdJkXfno
Io5oToL/gg489qv0YNH2y6SldBWNIR/6KJB04EvrJFiFcH/vfwDIXXrWr9C1Yhdk
+Fg93na+//1qEC12xWC2GRN7+E+6N7UidYBqe+0zhu7S0y1MVZn/x2GQhTv31HNu
HB86fJvdpZl6mIQFR8l3miTbUEk/lUh80qD6CeZgeCPVwkqUusfObVoB90MwEeSQ
TYPWQrQN4DOOLELVAq3YCkSSQM7eprklNrdmAOe3i3Et30NJzwh7u731T/M8q+nw
r1V3V0Bq7v975arifDLm6dNmLtTsA93+sX/1HHmMpizkNVE2SkwqPHfyOoc3JRI5
uW47zr6xscRn3NUSNG+mRl40ZJZzmD8loW0tGUaXQbDZCS9EdxEwd9wYVNFrXJIl
31KKPBk+Equh9APo3Ud/LmZ5XdGMeR4Nitab6x7JX7QCjgvxizFEJTHLM41F5dR+
Sobv37oXfOIjMmGpDl+dzEDPEdIGmyofDyt2NWqtgwflqa0TkEFUtRVmzVvd0JPl
/YgAt5zZXVQu4lqtYEuUaQ0CQPowk46MqyjPeiB9CDIBg0X/OoQfaScbIFnCWsOa
gLGnMwMBqh5P1pMi1ajvWezZhs3vJaRbf6GYRbb2ysyCPHndhDJ+a4xh4rIAOa/G
EuQS0HrF3kwFNMYTH43FxqkTNBAT3bfknF9ZWyGh/cdBJvB7ZWAPysepIK2Shpf2
cEyIgyFpQqeQOEZI97LiZn9y13Mx3K4NxKBsBPADCPTITbvCoWQNAI6EWu1SnlJ4
lEvqQ2+zqkwjk829HOr17zq5RwnwSBXfabb3xdmFSkwDxLT21z1z8u/tXYgFMvPk
7JMCsbamax6zrUmkOG96PtQpHwbTD9q/PfZXUbhZrxTDq/OEFDea3W4vvfRD9y95
DUu4/kc1pwAcZ6d91x+DQqMODn5jZqh6FUs5f03oplIWFQnwi9t45LESYoe/MRV0
tMssoVmlBwBc3XJ5s9CxN42jwArFRCFsXAVG/tUMQqBY9JfCUhg0SSMFeud1HOa6
caVHQWoPv/u9d7IAbqaSTDxSDdI/HLqSi6+/wfjSxzz5M3gN+/N6LUia7Yo4C0dN
EB7FYr8EOkib9itQBbJO3hgsyfWOmzp1u3bhWQERzhThsFZkxk2dKwUdijhW+GD5
SFzmZwFG0ZBEsBeJMfOmcMbtEIwbetse5FLxYLrYDHgEMpO/UeJqB9hXIxU+w3gx
pCknx4M4Dg5eXwMnR14oc5oha501OVbTrO0Ynig3JowgD9R6jDI5gAn25GSU/MX3
Z+bPsqfFJEl4U+BGha82913IG2ep2w/cYyzeVcckSEY0T8XBMP05jbRU87XWuLV9
6rYwBM374eEJS7vPq8KgKLKMCiWCTjuVSkhXhLmOnre3WjUMP/1Clv5gTBtVIFmX
gHxFjpBEcqMQ6ccJXR5lIJLSv/iEcWCQ33NdbdLVjiCf9kh961OC+LkaLkMqIEKZ
k3Rea9bGMr/9wMSZA3rriz6EhSKCpUjrnJS/0acteNEZ120HyoxsKOutDHHUpjNO
sdniidPGAY9m6g/SJS4hgHm01688+Mbc+w+QB/CFNDGIANvpCLDswThhRSmMIJRr
shDrDhpxxI0E65ggJ/4m5mdlu84QFXOE/eVeXkkaDRg+O/5ptn36gg/Y7FWrwFu2
k+MFD+n5UjHGmnXTX2PVrh/AdaKs5g846HgIu2SXDaxdXiy+Q6iE01Qp9N+eIy4Y
GctaYy11uEcxk9pQCwAj5Uc9eP/jvyj4fNAt7e//WbaD5xYvnhSzo2UltJvvmrXB
psqknp8ePwSMWpOXBkrx1aU8CvcbTl5CufqGGCBLKTRQ4IgJcbRrUCEzS2yOuXJ5
T4w53SeBWaF1XqDex1a9gIuSdFlSzuEgW/1OWSsUkbE5RWZGWDp8oG0OOjNJTTsX
oXvxs75HRi2a83Xn07hbte9Cu4QygSs+r9OuXSgMoi2RwrvpixmkcaArjE7co58R
QjsNxFbMLmTM7zQKP3JzWeOm0YCJUJ6zRR0B7x7JHHLc342ckFXVtcdp3LRIMabM
390eZTclP/NR6vTvuAAS+d6nJMEUhhnwr22XHGaE77Y5MYjcWK3THYBeEJ+Wzz2w
qqaouK3z9YVlQfACb9UdrSbPW4UiI8mmM0nk6057w1rOqJDF7OTC349iOg9YeRJU
3gw9bACSt6nU/k/j7jEJg0jF6Bv/rahXKTP8PIgedwBckYBHwLlpLr8rE3zN/xay
ew0/pjQAMW+uX5z+xP7iwzFSSZrpNy3H/Iyl6W4wiahEsX4MKcfsOgAF0mrE3r9H
E9uHVS8irwekO0TL9ooHQkX/kLwdOI6bremAA3gr/Ms3powUWEz/tfYzqn5JgTac
HYSTtFhKVHpAJ64jHB2nwk6V1uXR9d771dYdaFq3YYAytxYO307FEVqZb2yI61fj
SYC8Pmilu/Zt0t6OjjYvrHUA6ZMLICUvm+VMjZLU4GUXm0wMGhkwXxWSE2IN0iz8
zco935A7P9uGiWEZ72Cio5iAG/IwmooSDkuKYmI2veMu3GdKn+wVj1e5CLlzgCKz
9LuI5632CwCg90nE/dgSZijnZVzxdYW2/pOO0vlzRb++fh071vz2fctODDcUvbz+
C7IKVop07gCsJ3yVmQBve9GCezTB//NCIJ1MpF5su2Rg5TTAtDQm0Ifn26PjoVdS
A1gvV9XUULBmgpH5tweXp0ISRYQENwAXrx6eqHaIv26Vr/PdWsLpdWckcybZjDQ7
zs5xsK7BZhxLilCVqJBBIcCeULSmPZEV+A2GUaTDUp7VUUCHiBQQMskZRRVkRG4g
YSJ5MlZUIuGgWpYmXMM0rnSKsJvsADKmW+u85jYuk0ytzKO4T+q3SbQFwTjz8JaP
3URma3+0nQWei+ggb5m9FOOl3XugvsuplOs3J8LpIDtuzSY5aeVAuc5usEfvN0n+
gJboz8KFgDLa8RNAVvpYaRIRF2+OFrYore54prC2+cxRD0pQ0B4b4WJXaMrh0ff2
hJnaRaKdz/n1/li2039z3TSyjm5K6uqas+c9eIoS4lB/pt/QiznbypNp0MpZ32Hg
uCUtUc0iIMEFpqsj5l6Bg6BkZtVM3d8nADC5EWC8SabVgQ0Ak2lNnfy3uidsJFiQ
gqAHysbTKdr8U8Q84wTPmuTVshuXIlCirF0owzikIlU/WY/CENxpDPKFFGwTzjm0
1hFs5UkKKaVuSpJcTl3VbIONvIRkSLw3uYvQhADHnYmPd1X+VcZwLC244z3EflG3
ksKZ/r9i0SQuhsd+MY4VY5AQDOFRHVr/Ef8jJrXGKCsZly3K4XZt9r73izxbDTHy
I0qAyQAx7mbclbgFHw6CuK6QE0ChXMjvP89EOdu+SzEwwMJEewQSwlcjKTcb9xdr
QE8mcCPvHlLuwGpsFZAxINU6wE7d4RlAzAuof9GHFtuZCz4gBpU+6FpkRbV7nIkC
DEUx+kJ7M7+KlqUp+mAg/EOfH44RW8qSK0K0mKNJ5rCQ/HfSIRoIX0dsSs0mzvCM
k3jfdUeivV1DZya5f8rdA3EEUX2GISZc85hZR06kbhGVb2c1WmudLYdEboq4rGBz
utpDiZcujB1Jy+LkvsloCNjjpCjh1W/USCm8BXrDH5L+o5bpsOLAALyrQNXSFW56
sL9aU1V4JUfMDAL/Srsg9qNJBL1INLlcaiGqVFQR5vHOqwN4g0Jm8nQlNU0yHo3o
8J9SwpYOHNp1D8xeWTMvVtyYqL8JCb/HeWAu2/L/DiG20G5NlQoyuhYwg91v1nHn
nBIBB65Xgdn5XwrvFqd95hl+ma1Z4I1upUyShI+1lWily4lOVHCjyBwVbwcLiEm5
cGTq0+ME2n3A5SrDFsepzJBC9KbqLBrxeAF0mHFrcUBsxD4Qu7uG+o0KvDZmwI81
B3/zGTOANtJ6YlHGnraJdFI0BLxwb7cXM+26L7ytSd30b0qPRBtf2uQxZQTl1uyl
0tlbSmaMEOAsNUBAWkFN+z7I4nu5b+lIQjr0RGeoOL9lzSTinvS8BYaKrd0ncn1K
7tNUJcLmLersQ2rw1rIJzNY8HHa2ar2muD8cj8/AGLIQuqlQ6mb4O+yYnYLJANv6
WNwqPuiG5hgcsx9lM6ZqOGsSQHcHYnhUfI6dTZV7Wmv8WF5JlfHG3CgPdQA279N1
1Eu7CaqeiNIFMZXwb7rrggmTQegGYkTEvEDVFEiZhjFwlr85pRBsz5xUQR7OdIH5
huf24GBDbA7J25nck3tH1UvQ1LrNu0AiaAS/CLCCpZ8z9Hvu5xV7/rQMndR9ayiY
uXY8r0B9oKxi+hsk2eLDWzV5KjLoPjJ29qRGNKA8v56SgZ1G2u/7tvzOCLy6vEjH
2LjHIuEoljnnTz1MGvte2gQGpcVeG7aWjR+K+/Zbu3EpxadRG1J+voH/m/xOKNso
Ui7Cgyi5e9ukosezz2VqeynRrUHUkjhDOjlO8coilgUAiDZwEtv37UfO56TTa73n
tyx579S/5qm1fiNz36YYt2kgkLjc2N8GLZIv5+7chtbWy6KVvvfFpqdoABHWFnXB
WxPhEnenVKYAzisq6Yhpln+6v/YmqTQ8+AgLkE8YH9cLh1Se9W0AkeMO8JZ9Wwz+
j9bkfFkNW1Owj615kUFtHFpbyVeasiGeS5gx5whA2otO5IvYuWXysi+2LAJuig6h
oXbvnprz9NCnXq9D+yaZMkFqs8XDUu8OyIvg2yLtQvpjpVuO+U8jg4xTuVqOa1VT
id0Mr85lJqdMMwzErfcSVZR1rmqcas9oeEMQjPtzUj1M9ZTj2F2g1iF4DNBVHqLR
N62uRfq26LTPpCambXxxHCgPRPTRsicGNFyARSFa5JdDkMPc7cQpsuLqTBBy28xd
hxqGRuFrZGF7WbUY8HPriAXlsAXtAmhhyG4rWiqSrOZo3FxFQvguEXkpV9alLXfT
EJQpJ9r/66C6icWf34SpGkKDCxBKI6emxF/i4PyL60YquhWdMvncpSFVV/Rf/h9t
Yxpzfe1avJ4DBMpxu5jDbc4z/dZcb3qMhkOjEpVtKIicfyacDTYsElMnzOJuMHZx
WkqXjkpjcMAOT57GHrD+KOYcoGRVn0+cVHQYFAZNjHE0clOcQVf9L/9a1utThiPs
vuAOnUO1ti7inCGIdOntyw7tmPOuYYmTHh4S6wHr1kh210DSWrbbex1/J9eSHeKN
g+LsCvYhT0t0vfqMKZVltRAvMxPMUVc7RQ1c+T8NvdXqNT49GvRZmVKkVJkiEQOf
Rn4fQ4HUm7n+ZdVEJD5xqtiXtFuzeGKISu8V3F1W54puHuUAyxC5lx1fYtpxQ1S8
XnJHDTrkZIEU2onavOeDWXByG5l8+jEN8h0zG3kKEpgYLDapuDHxUBaGrgqFDEP+
KMwlm/oEjcK1VTYAT1Mqavi2wycbVlVBio9ugqXWHuUYDCezB6IAERYCdv76Wvbi
lwLZ0zQqinNEGsaDDiYOt2f9lKHB6cEL3pVBmGpGxHHTFTH5iGlMc3Fs/MUbVjYo
O1eew+3w4bHKRV4QnMWMRafyKPN7sWXCjy+x6W+Afb9PBHBMB1n70FbS9y9aIK6F
WIUFsxsv2drQvVbU96EDUyMq8U2TynreDa1yC5lYvDJx9CTnhlklcbPvOjxGY8NI
yTzllPpd8IQwSjGZ5wiYwho8gY1dhcNbMhZdfdC9fyVWD5G8W9xPizsqiXviuwp2
lNXdXRb3Rd6TPzuo3+079qoEZqmj2qJ3bboE24e0OsgBbulOSczNum/SKBuBhRQ3
9dbMD89rIPDY9AbnXhh1jDrDisQdVr9cr99tPnMZGze4S4xRPxe14xWVE7/xQvJ2
M0X56u7fuFtqgKPvhTXPbTuEihBLI1OTJJcCLQdUeWVQjueWhVWsHedNKIr3JU04
z9S22gBSgcWAHgIZcPFx4TzUU4X2qn+rlp/iIP/zO5UFdBwCr3rAm/p3S/nMErxz
9fDkfaxk84kBiPrtBvigpVSRJyLpRQnk/G3H5c84SsHRpeygE8WxFC82NoMXP+Fe
6MEbYqSEbtUuhTWyn+cSMKCClrZwnz7+hcIKsz03Hphr6Tz0ehmB78QCd7h0yBMr
ALrFzq4kk0TYELhf6NFj3MpRnwZslQ7SFCxydIHwOe6+vbrN3GuG11+myVRAxV4i
VJAU7AM/NehCiWOZqo5DQJvZiDIJKdLBPIJovzRk1DGFlqwYLgrql7YC3420mOvs
dOZ2TZRUJ4S/DYXbZTt15jRCJ7UEWgURRzPDGavHhR98DC3DGCE0G90NmOO+db1C
+2rZMR73ONh3cWHeTyJWYotmSDXVHfeZrUVcgJ+b8/gcD/kvTUbzWwHqp3dTbtRT
aIvgK0stouVtKUJNBC/d3tTVN+3t2L3gD2d70qBysrgJM385gRJTCG2gHGjLIFho
VAkK+YtxSVW4Dmg6TSwcpZwc9skIYkFqtiSNHYL0wandLMAVOMgY4cJmPkOXFBbl
2wrfuJLfIAyQmj1z52o5met86Qe5qdEs/9i+Jf5RZlJivQ5LAejfM0pZBXwk1+8B
JTvr43rMgzUvIWRMgkpJqV+8Gee4ENnelv4c9nC3phszGB/YPCNYkPuwI5bqVujI
inJSaL7zEqK2VNsf6L7lMupAPKQKrpEU983Y3odnvjvZGNCH9uIioPQ/GaBBNaVy
bwHzT2DCGk1bQyxph0tZXAiXqXLV6wg0L9dViYnv+AJluV0XgorTkx9F4gbjQOuP
KMk3g0tS9OCRiU+6I2/WU9VwkNiqGg6c/xa1kLjBdWEuJztoTQKm1PGqovDPbGLr
l0Ed9FlJX+gO6m0ZhMyRBbbqzjZXdCWV7WIm6agAb55nI45q4YwkcwcFYPYWnr1m
ys3b0oMq6czzC98V68ij5kn7vjK6M+uilNf5+Lo1b8fuk0kRfV1wwYzXTOis5P2B
cLSt3EE6FhGRzdYEXNxStj+XRqxszR+fxcQ5WNkJr34GxzAANlFrOo3h7H0Vbrwx
eFYaWaHOCI37QYPj7vCsQuEjTskS7Ma6HUWqdGyzzGpZfxEGfCEMYY32nozYVKFY
8Vrn09bW8Ej6FtRCnynOeHr70DAcOV00UmEaWXj53VnA8Pg0/72stERphkXIE6ou
ibTWBbgwBp7f/C9OB8IR5hujUKn0z521kMQlTvWZs9LUvdAl+BlcCczT+pCSMDQK
d6oAb3td+HUP49spMxZlxRPqQ61T53Rv0T1haHwxZGVwCVRh5/s1fh8DV50FpAIU
ytJNYBx/4YX6TpGLcFWJCctbB/ik6ZKfN0Oase3Gn8VL67n1nxnb6/KBv2/s7KEa
jiCqoPunLZ9r+s37S3GnXFGOdPlogOTFjyGmt3xVhj6f1wdhINqtCsZ2vHlXpE1t
KpgHWV5ThYFuJn4t0zoNpOCIC+/2vaUEuJmNcM9nV2zsBS6z7V5zSEN/N8p38v4t
qL9P0LKoMdcTZeSZW+ocjvbIInIF98+eYW11zQYtVHm+VBmyavTIPdoUd50zVwPz
xvy41AC55Frqd0SJMyK+XYij63njX4j4aCsRMiqV+8LvM8U1HdPjD+jiKAFZU+tD
DaDpwEAax+puffZQ73pG0+3z//AESVL4zYOQ1yVo/s6DGJwhGfBqNzKXG2AV4cxf
B+uTNIya9umHV90UzFKZULH94XXXGziZOmeA9X8/SyE1y7Uh/OodIHDUJEtsddkg
FP/xvpqBV/FmP4lUCyicr7Woimm64LhWtgSGn+Mftg0EWhhhSoRtP7N+0HADNFGs
lWSRr5MeFrZ1tGp4IsoW0yGKGzMrGAZ7Woz3RNphRcm3+l+KpdYc1kz0kfbly5bG
hK/BSrN2B7nuCfvRY/IG5VLinDJVT6RcOmQ3k7bJWluIY+5+HYfVz3GhGqVimM24
whbQvZq63w2Gzjo3yRGsgbYlhmJbyJ4xzI2ibjW6A17QICk+mmsSYT4Ya/6QZdL9
cFA2nTPknr4fmNBKTGpUIsH3Wc8ZJIBsBWE1TA2DwaRNPROzxDM0r5pbM7frilDL
ELH5ll+OmWGSwirl0RZuuE6g544n4urFsbN9p4W3AtDaTMKg+fdhk3lYMZ7gnsn1
Y0AlsBRG6OEzmZIH2Aox/pdFZ96LUzQthYDQE/rqV5phrMBLEp9b0/C+EZuPHtgK
ysnvgJjepQXF8evOFIo6BBqLxYvykRkefxO9Hp0BQwpFI1AjSGz9/7OpAUrQ1GtN
dlMLVXWLlmIgkz7sD3dS8EpmyRvB4irN+GxnSeRCz3ed/lOyKMG8RMU8DR9eTcZO
IZ1bHm9eiUJrbZcwcqsGJCc+ySYSLcFmBJcKXHXB9kIJxmrP+L6q0CoM1UQZd9d/
WHgsVVPGc1/e4pWaSttzkdzhxmLPVq6NVuxab9/ffSxBdTwHLIgDPE+MSAM+qNr6
nZMBykSmr/Sepj3FSglzps02bhoIvrgCWL+JrEDOjlSZ8GyVJlAUDIaOWbnFgFft
efgnL73cXpQYwqRhdLC4ZTO0OtpCA1JmC+Ttf+bfiHC1epIzTOdE1jfJ1a9C2zf1
p74AjfnFwkGdHoF5lhd1vztdy9QkM6W3ZBc5YBhWmELp/P+nXFwKxde5x4OTaieb
IgRm/Z//2Oqx2mDJ247HEVsX8H/iUDHsNkfw/GhTIqUU234cy0St61ZX9Z96r6Ii
EPocowhRFv2YAkXQHx7QTQgVjlVXdzAIRZhKA7cyM8K3e8LhoWFDRtnoH2bn/l++
Kf5SRY0kT+cfsKPynffHycwDEEzTITFU1IBuHMdA3NOV54KSH3QwwcxpO2KvR43Y
kfdNCRymgdHctML3Eb32Pfj4uWO2SFszfQebpY+U58C+9IG9NunjkI1bqD50DAap
ZImI0FgO9zrqcJSJvdBiCLA9CKfYlxfBacey33sLUd/bKmEVGCNEySXZqKPb5wyT
5+s8KATIX+GGayjkGWopQmQVyQvyuFpe5O9rpU20/fpo36yUP12L/vz4D8+pLffv
/z1/5F+R9+bVba5FRe5tU6UKaIgSERLYZxhJSpz4ErsdVqz4rUcQnUe0eXRdjJ1t
lviGjdfRDVS/49rWqxnusIHE4w8/vOKZ1BeElq+D0ZrAvLU+8fwHw6GV+hS2b8dN
wN58ojuZGe/lLI7uxI7IgxBIDlw7UtyC3Lc2U2iUcZeAIL5nml+PUzkidXLsEWp7
r5CWQ2UyhMyM5lUBLEqLAG0LkUWSqZ/KUP5v58XCiEcC/Z/foH+YYOwbUro/qgTM
lmxCTUjA6kNRGakGTixaxt4b4AgExbqLDZcWG5m+1Ni9iCS9Ls4Um4Uwt87nCZ3M
RFVJEJC+c60tP9eVsDgzs68eHFWclFXmhnwDUKE55znJnXxHiLphgoWejljN+7EH
3w1p3P+EQLb3CWftXYSr5BRKO4JT/3LW1vk/mj98xed9ULlv01+ih+ysB1kD0D1K
EOHCvofH1JQBSvfzuR0MP1ia35CQkmDmNT1eGmkO8z5U3Nu+0gxk+4Lbca+/z0DE
e8GRh0NA5NEND0EC8XoeMaPk5Co4kfIgztD9ECGMAUwJBHUOOjZlgtq/EcVzBhtg
+Sn15Qr2Mq4nOzC4iTG5JpqUBbeR4pnN7Ni4GXtJhyuJWtNBTqrTHUXI0louR1gf
PysFrnQ3ZIg+zfc4eYBdxuGYwhtMjRBaS0mTT3Qn0YL8e7/kWZRX74Ba7ioNG/he
FCMt6f03i3ZbuVH3RrwRz4Uzl9fIZ5v7OPRuBRjDvaw/y9aXvqQ0Zng5UDd5M4Be
eJpXV0ID4EQQpQdB/vVY/CXajcIOreqVfe7sH0L7zWPP/XvbjDyjwy3Iw5tOT12c
Z0l9EkHBNhj+n/K2Aq4J9jRFobJHUTQnKBDxnQrLMeopMBanb/VTBocQ4km0kxl3
n6acu69+3AGTqeaGhFovDyv28CHIz3CkSS4us5Ap2+CVaeZmoBq0eQC7C6y3eErC
3G7eV9OsgyFlJx4Jb3wniNE9ozTJ7bUXObHYcWR+Aoe5RK2dtVkW7YvmWIz+EtSt
1S6F98Qc0DAPDc6rmycr/d9VBdB77VoMU1miwRNYPyHKYg3/bLB4Fi9AzNbCAJ3f
KfLD69qJ9Unm5QGd5D3a8+IxcvelDVJdI2DvZUNBZz+NYuXMo33lXNj+CJixtBQu
f5iwsk2bPvboZshzxpO/tp/uumLHKFc+GAE5kSFec6pz1yrKsF9ehjKi8fGuGgIL
+Mj1qDOJ1G/zrosczvK0gc5WtCXsKFdvysKRWj0ZddtO3yaC+WtlD6IOcfoYF0Yq
oCaIDuQylU5PoAEw0lXoVz/hWIvjfBOZdr1JEpCQmO2Uc4lTuRgm+mb9GtJq1RR7
R+crzkAXct+BfO6UNouUqHJNEwVC2FtgJRyTqEUeMarLyx/HMNJvpSxE1GJBPsTm
EkQTPs4rVt8SE0JyGGGj5VtsSOMxaoW2vdPToADagArcxOaq33MCP8ExwE9/dYrr
6JBWesy4lHARyaK0omtDgcUaB5jdXl96V3YwyCy0IUXtLkLYtfyVR5Qid4emWSRR
GRp9JtwBL4VCyVLUzs99RUfgEht7npsVT8NTeXuZUllN9oP9pA9poyd/h1sMWTBo
uGUPKhuUcLZOpiZmsGaQsrympefq3WUtQtWYM+uDnD1f2mN0U0H5Zl2GZ7BUAto9
Mn2fa87J0JcC5Ofhuhf+UrnAd2Sjv86r5s7adwS6gn2f2x4rEoeRS7Nk8AcXsbRg
B7L2Uf/Sd+4qvdarLy2aACh12yvmLp6XXzrE7KXhtceKSnCeCTy+zzdgECK5PMWD
YhkY6FcAj5M5aws+CIRz/ABf7ymFvnF9jfIGPKYvWufhdGgyoySLOgmvzPykSMAd
rS4I75hHPNXoh3Q/aQl4Jq7sZXF9W/58ny60wVXIQcNd2IPet6i7JrHJ5PHbVw7A
hwla7SRuj2WzUhz1XdJrgW+UK6OjEaIJCvHoirQyBnT8xcvWFAvcQT7jRo8PBerp
msAKhGYyusONQNJhtHecP/FcpNYZIYRsJrS9wvbzgspxO6TaE4fE6qQOE1yL2zby
GfNqwZnIk0dI7Yk6nh0EfRojdj3cd1842Hh80d7yJzVmLN7YuMxo06ANTueHLlE6
C5F7a1SrTBBsSbluVlFOU/S/NP9Ym0DtVj9hdQ6vMz/M57C6A/qAM1Qjw2VCXvG1
skComeNLykpmdPR+iAG1I/v1xbrWpxmVZpvNU2bpW24IaaeRKoI/871nas8ER+Kp
6c9rUYhIoxxoYf6XTxYr5rcIR2qIbIaiP1C5d7WaHx2QEqBLb8yQkLkypUw9hgxG
Gdu5IE5EblwesoLWXZN8QpuK8NjDPRvf2E0pXQhsLyb9Yzk9xSW0+VUICqQtLoVd
Le+ci7ZxJZOn1AsCUsXvge6FxFSHoBkqKMkjbxf0AUW/LbYjZHLp6OJSRuE9RAoC
WaCbp05X3qKVLznGSeMD7ovG2rlf2QPVzaCP+PvF2j5UdmX/UseUTIKaxOK4AaFB
cDv6FTCFU8PafDUkG/8Mv2Mx/KBoWmBLpAeQWcHGlRMG6eo3YZ72xmyuTNwLP4V7
4NR97b1wEwoAEy3ElLhIG+io1hx1m0vVsbyE4T1ojYNAD1tQKbEkbC2P0nhUcIg3
Sd4M6y3Eompty02ygUIRYy6RnJ2ukoeNO2BKnj+EedrvFqUHSjLh0Jz2yxKZT/yg
6iZ/MXzVAwx0lHqcZyXMCrO+Z9giRuL+A2i4j9qVHLoCnLaP0VeDC/sHkWxufGUV
lRtjC/p1i0WFqQbS0EloVmLC/3Z/aDa6JJsX6K9OC3gxwkbCq1/tVuFFiT3vAW9J
Gui8BEcyOcGOx1Vay1xe0OShGD3Or+on1wpJrPSUjlfqrkjr4Fm7Ui6kKqv6tdtB
tQaorTpKuQmwQvPL4tkuHjo3MNaHIFw7S+dtCz4t/ZGNEUMLs5LfhNskyuprNfdz
0RnoKtg6BYuCwFNGa4T2gilH3cJybRea4so2yaS311GPHmz4AJVp+QWHTR3AbuLq
3ditNLJUvxidGcpvu+Hdq2qoj1nHTTqBicabrRBvrjQD9yf2sm+BqWyyqwrzq4cQ
MIXwj4Bi/8MQcdVHyAj2v845SVx2eoh8fVR1ggkO0Va4fGl+c4CHQfyNZGATVKyW
Ldj/yq8FuEo2k1d2wRuwjmMJ3UnqGAACsxPaig8+V7T/9Xr+P1tjBgDhgrgCw5H8
LfHSotHxzmdwSt3UIE+HkORtVs+ifb/rg3FGRkT/82zTrWGFB6RgS4+8V46Wva5P
cxt7/WuLgbWy21PmzNzJqAh8Bga5zsN+/cv/sA/8xK86u+htJ1OEdiaUjq8rdaxK
49i/6l2lmX1syL4ngB4SPZlE+HzSm0CrYJ6PIX/XG7HC+ZbfURshHKtPrjTd5yOE
cLkN9umeWbMwdoaXAD2Rh+CZRgo2/K4o/B/A4oSp9lDmVczWsSfyDAejW/8oZ2LC
ZXnSZFIE+mc/AqUgS5ZroMjDub16PVoWu8isO8BSrO5vEFuUkKKKQ0ELHXE6vAyM
rLEOhrANGCVl9Bv8yAcmGLiaFyypQ8SbNMDwWOQzWQ96Y3NtGCGFnD1BU82EvOvR
2/SXvvWJDrhYUroZH0SM82apZ5KEohqa83FL6KQCZcxWs73ENGo5Dz5nDVpZjh6S
2cgl89j8+JQns4nU2BFGyKkECVHWPJBVpZDc9G/vhBj3ZACCL9+p+QuRADlMHFYQ
YaZXZSymEEO0R88fPkvlfaNCPK+dWDN+5tocEWnmE0ML6ibKzjxk7defj6Eiw0j1
uCOvZHjWqnb1EU58QYOX9yjUZ16fLtGX94nPNAV7UzHom55tfyrBN0QGP1X7rzg1
Yge5+BD/ilfHbruF7WbVNLsChWFbf8v7Cs+gMCPu9qswr9fcZRrPfbY9yrTRfh9w
yvO0P4XtWLL53LppURfVA/baMU+vI6Dgiy7yBVinG9s82Fyw8hQMgtKnbbD1IKvH
HF5BaRfevGmxdcsL6sZ8vHrhLMWM8tgprnrss1zgP+J5Z93fLiPw+jnfWRVIleKM
z9MLw2HZ95sDhpRsn2M9JapLhDOoUsmcQ8oLIz+VBlYt2uCVXw+FauxnOIK97Do3
e4ZHG6CDH/4OKYFf+IhlhTgcV+S5gDU+rOAHHaG/NcMC9vI1bSU2bw6IwwKL6LaY
u1ThVxPr2rciU6PgxthLUa2fH9x/DI1uQJwSGH7HEg+vb1WC6rirtqPgQYVWzJ9n
XyneDbouri5+H9MyZ5fYe3UzEGlFPy7eWSOueDuuCANubwea2YjNfGvvOTtFipEL
GLfAiIfW1ORQx7BwAXFzbg5rwao0J3gPy3r6VPJpoQE+LeI2ZBfAQgy0D7+LOLYl
dWth4Bl4DC22PHO0mncIk8UgnBXupEdxAjQha6hhGdd9i0zDcBJMSFCSO6/e4rCp
/sQJrXqNsv4qUFhCBLzOEFDKvcUwO0ll7dJwEkGEWrd8TALWBgP/fR9UQY1LofZE
Th6Tzi9DTazKSxYXXpNP+/myZJld9FQJerk3zH04zXdBmZQxwzVEA23nafRDzvNc
DK8IbNSbUvToeBfT7QRxYfXXGK0wtJt0Ic+wLybLHi1UxyILOIE+l6+lQ+J7j9m9
ut0G+NIpoI+WTz8hD75/RBuS7lOE06lQIS8Ugoa830CgU6FbltNduFjqdEmDoAEq
WI7CilSH7H0W0UOSTa/IpzlTPIJHU9KIaOITt338Ytenc9W4DTDiCedFkLqrkDxz
BiWDGrp2JhpbgaRGUJwBlblxMxbyuwe8HBhCeTfotS/QAWve+9JXPX7ijqzrDwHz
+Ji0FFsMEMYBG4/U7maSM0M4tBi779pvBLa3f/DSFOW2Y+F5G45dVBUw/mv5DPHh
nsKsZn86x7cQ4F5bOGzH6sBB9RL4zS8Kf05GMmISALInSyloy1gB5PCN8tY0TOvQ
8BehsikUhOPlp+OC95etH7bn/Iok4ZFeqP4+jHnsDfVq6b7UDRcpHU6iU3Klvm33
CBdkcm5Oy46iQhP/77x2KsHBulEnmix7t4sCq5ORoa4ToyrrJYVJP/eqOQnxI6Qh
0pGqvqHyukSXEJ1zfsS7g3z4baroAdjqpK/c33x0F1P+eIdsn3LkUXwc/mtUPqgy
jIIMOwrpYcXz9dDcmE9mf2ed+7AFE0Nk+luROD+nQf/2BJrNVVf+wa3zJuN4L79t
09WIXnj4o9KlAIglSTKcscdQhNojg57IzRgxTi4Y0KAgGx1/r1cKLrDPVHlQo4C7
4xO4byfIwVXPLQD/aXIHR184ZzlGq4o6+BGUgLSJIUTtE5oqFBNZkWqBVnYDswo3
Djkq98w3LLVCHbxAWV0lp/+Uaxdw9jk03SVsI4ZpjNA9wRE/hds/Vo3mxhMi3UPV
ZVJdLHV+aUmgvDdN/JapIf1ahksMtrj2m2fygEC3H0WxfmGFKYRtDUjkUuPbIBfk
9Sc7Ldbvliv2pdBf6kHUOPAGMLWtLD+G5KgOkg9a/RqdAThxjpzBqlQAYRcixZKI
k93moVC+XkiY147pUa8wmj1d/IMPVOJ1VdrdEsQnFjv+VOUak19WtkjXDf+KijLa
HpmGrec2ZqlF7bZlG05Gs4h93et0fPERdZBhAHtDoKuFZJ7SJhrYCNK+hbcH8eAn
SsvwEB2K25No6hb1OH7nA95yeYvDVNdYtrFy8T4x29P9NQGgdAEgDzJsYsfSwZMk
wRMwv0SBz+tvSRg6xnJEb2Gk9fYULp/rM1RV2NmiR80P6tyGBWpT80l1Y2NCM5QD
DN/FwEhPBWLXMpPo/vqhxVDo0w2lL0iHqflD2scDOydgjqSpFP/m9SKQHiiBpU9S
AdPssGRmWiaSNT51tempuUGv+HU2J5hPuu+5caacuCO4I2GN4V2nynn/DyREQSWt
qUnN2+oeNuM1CkodLo86oBl/h5HC+mIDVkwIRMhubYqsFfC5AVb7okjS6d7Qjk7l
SpLm6j+ripkXVUcSVH91+Zi3bc79/1eyNoa611zU7xbPaBRm3d+2S5h3m3oJp6a4
GBGV+t9M9GeOZjZHwj1lzKZ7f9zpBQe02vGGD7L12IjlnydfByvJr4VH6a4XrRhs
hbY5YUkrhwHkhCNJbEQVNZZzebPmOqMbrw+NWBMU4nSGFPPpWxywSJJKKXpwcRiH
Wmh7EX2S66Ab8kVXo386D83fFZXFJAIxbX6K/PBZgIyJXA86IKT8sI4u+/uUI5vO
vdaKmVvA56h8yjW5taHE7jGXj7C1d/DledmfIDUnkUMupLan8ZN3NOFX+Cek2CQs
jva+x9rj+VCN563+dzImjhutcckk398j7xJNtNfLJJ3VWtOJ6z9Af8nRBPmQuknw
67dcvR0prV6U4Uvg3MRUlNBSaC5YWEkBQ5vvA0Hl2LFtyMVSjegbpDC4S6dz+xHD
4OdYvbFvthoExfhTcI5I0aLj2btWNflozK1VS1eJ1hQ17DpAGH6CjO/BO1znLr+A
gapRdmsFZmh7YWGuzxAwWeMOQ/vfpeHE6Vqqiki7Em6AiUmKA8OTQHSaTFOLIhtF
GrsVbD4S9K+T1FqiF2on/TXzOCeBwfv03ms109lDZUUyzgS8OmZxfLZrLmy3k4Cf
hugPCw9tZYtwW/D1+8iU9fkTzcU2nx51f6mqyRtkuf4wrjgr4NXCGOtp8Kdd4mK8
/O0gsCNGkehaBSH8dqj3NZZQKfGsr3C6GmMU4+4QMbCO7fidEZFTWt8c0zClEfAj
5UuLvtwjYiVEdUZGLy1Sv77KDVjvY7irNCFzLEc9gbojWYKZV6HUVT2lq2awDfA5
DjVPGZDe8gX5xqj4bnDeHQ0jDXnAXRTPpDHN43QY6h7846mM79ogSuDnlvXbCkLw
m+7t4P4T3m6pfZkTa1KD0r4kVYvcAEsogEzhvTFt39Az/Ix8+QlZcVotBIY5lvyH
GU0t2Pa1V2dvGHzUpogSm4s7E4nI4mesfajyGgaIMgGMWeBaGbqM4GGKJz2ZqPTl
uOfV/nvN0l03+kbqaogJcCqGVyhxUE5rWEPnqHdiTr2t23gHtijtNqe7jzubtQSr
4ZGXsSqMYZRoj1SYNSkXgfxNi/uJB0s+Pak9ZN5Qk6rZ1snRdMpTc42THPU6SEfF
Prt54nFlo0IZEqYJARSZgZUmSXiFnUKFrE9yH3VzFdBWBxKBb2WkaXudRosojVbW
8B1BgrRfcsMPrPE1v5Z8PtDhg8QJdQoJDTYFNXjESZLL6rqGIn4EgEeutmp/3Dsm
8zGd2Oi4KWWHvciCXqsUWAHUuOOk4ISWcpkw6hLx6Uf1gzcA69foq2iPBBRtHFF2
OyhNyh1IkM49ladTteNhMl7txukViHc3IiPE+56bXqpNCsn7tQX49z5xz0kcolYp
GxKWwcTnR+VG4djH0p617L64jOH4B0YZt2gCORsnSK3DhF8JNInZoATiF21+uS5j
6eZp3m0IvuAs3Us+eP61k2SHcTvx/M7klLpPjNsAij5V2p2ZAC6KWVLhQysBB9Ii
nPOSGyYemhxJR3etQo3QPxxPEWbI/QKy5NPGQ/5jE9jBOAWzsGHzUH5dpkkaFekS
XjTK20kL65alXlTX82jwtvu/3BNBqCEKIo2OXGMmCo1c/0yyTcisqzpHv/UvSWqd
p81bmzbRhRILOeo5bmZnkWEO2aitgQdPXiEpr5/tHXO1C2PPgJsWfEqQV08uDLek
PVc5jDo4EfB90ML7ndXbmVZvn0zzbtktUse+TEP5buht329BAPGs2fqY2PHHYGe7
snuIyNT1nfu7eWWgZT+ycubsNMyJlUDILknbcLD8DmNFd6BchRc5YIHntLt0X6ti
q31KzhHU796l6VLD1nGI158Ck4LUDjr0yIoiNJM0/KMpNPErBjDNBE+W+g3QTFxY
34xYN02ceqxKSnFjspEVbEr2YU/lIDCqSHxHlvI6AVbuSJKR8DTDfRwycS5Gn5Lf
DGhsxFcuS/kUmFEIIHQi2JxyrBUG2yzwGK0v936C7N1Q14iGU4WoxwbVRRyMR3Ls
wnh47pDzM+N0+tKJt55o8XByy3IyOKENCnCkSpxfirh/lG7YK2LsjX7PQ3s5ouau
mEXTZ5XyOtsc37YTY0SQOBIOY7cdb4tSdtuQtsGAJH6efkEkEPf+le/vfhXIcwDO
5Chgkls9rnKjuxMpyrmkC8nD7c4bbywXp5X0ipaggySGXfUFgTS1l9P5vkBpm8F9
Hk363FHd1cXbbxtunqZ402EUwlLzS148Iw64cEon7O7l1T2/5wplJmGVbkW+LlGP
ayc1322D1sfF9Rcmk+9grG6mD+a9KE9+ZC9I7lJdOLN43Yp8Y146J3yZNSoMB6sI
wO3tE+0baSVHeDy2msvDpp1ndfGcAx/IyFGfORrlA9ZwVB6j6/WFPuuTF/OlTQ1r
7JthafCAsOAFYX1EdPtrQHqipxALH3Wz8IzefCrVnxGyVNF/G66rmx0waUMAF6cC
N2uy4+MgOzebLc9O5VhafYd5E6/wS/27isin9t1HbcK4WImEZYcisX206jbxPOVM
ozw2yymPP0XhHH9d2xpNybG2LPQOU0DSFCoLq/XFU4LOFRIZ4/1LjW3OyKnO6YEm
xoNaX3RMW+hvLwPYrZVh7FqeRQhOCbaurwEe8WzUagclhg2N6+azH8aCMCbs8xKi
jK8s1MvAdrbpcrkAH034qRj9nke3Cgnckh4hqQi8AfG7+RDYKQsb2DMbSomXF+T6
NZ3bLVhIVBHbsjltK+P5t2sUI/4b+lQS4m4BFoflBcYVns/oAPIXZ+lEpmQCfvyK
YJacU+7qFbs9bRSyR3jzMb4m0LyFUYleWGkllyy9jy/HRmKGHK2u/ds+rff56LQl
GresJ248+0o5MXwhZQfnGN9Hd+WlE8VfDZGgwvtKlRRDWC/6jeZQFXAskL1cxCLn
+a9kUTn5ZgAwVDOOC0bkVffBmEb8N0tHLECUF4vUGF9GQuW+FRX/tyDFVAoYD8CI
jJOUhB/nxn97tSGPcCuuTUwbA/LmX9Ldb/w02hx+oQ/g1yN8NSahQ3FqpZ20HTx5
rpl6kt3Y8Wn35mS1hH2gFTHvWfGVQFwZ3Is40RPppAqgOCbZPi4IEwXq40fa2W3T
hijtzL2BcevNpPMGbXbQJGLc1syHayBl7INxpbjAfNPqsysl3GUYFy951HyRJGYf
oPmZnRVNor2mT3Z0E7dQ1roSevXdyXrhOQbIASQwc1hIVXIunE8ytwx+pdxE/VJs
BeAV+0fl43rn01bjrD1KXN5d6FerAKOHljaP6RpdNyn+1eQRM3LLrBZ/pO9IdKGd
E+4Yh599deJnGIEH+owHMnxk+MHnxSxsatUHM2jrNknfvhEcUajsPOAi7PmUbeJt
qihZvfhTjrvpvItyQpJd7dRkgJ4D/K1GhFBijlmhNAEy9P54IQ0Gg+SgHHCfZ/qm
/giUHV+46GDns7TH0V5IhT1f94dM0iXjFz7FU9zgxPlkS5xgcnb13ClKe1xKGGzc
jlpLqNX9QwwSFa5giuU1N0Ed2AlcD4itin3GMAtxXQrDl/47AoTr+4VzCzOSOuys
oJlKemRL9Z/YEvrH+Z2CmfAaRKxZ/aIHhLCXQOlQcet7njM+ZJc1E1ASmZcBgz3d
haKWQcakVnXmJ9v86DWXwyS8f0OlzpJqDvaqKan4mkabDx5MkS9PiTBlNfCWwIsS
4HthhtXPgfbdSTOMa/9q9yyxQv73qoGn3P5DjAdMJ7wgYOVo5cuG2rIG18OdKwnH
W3hkmGtUP/LQycSTOMaKlZv+nKEj8D3t2O81tV3KXlaO4n2ps6NVpNQ0VZovSWV2
Gl9kqgNQttX118LCnYQsjN4kMd7ECi4xzZI7k6ohRlamap0kkE6AmELYjQmVc4cQ
9aypA7ceSqsEoFLZQsT5Ys8d/m9q9Qtt1KaBZfAaJEAkb8IwQkTBxz+LOZw9OY/M
ZlJlFP3jIPAUJcdGRrfui3+pYh0WQWFQTkh8EFFcjGaXkLJs+4H4jTBOqCdPYvu9
r84MfpAQJ78c7sXl12y1o/WaxJFgITCX4vONWSUgQb7pJ5QhaooaLwBKXVVKK78O
jCvXaWLsTlXM/dRuxqMa3kLNJ75MfLlRGR3Ce5CAqmjY1VKxqLzGH/eNlDa8kmgA
0hGX9mSZXZM1JLW1/VN8KYBs2PtahLL2g2ouEeeNAp2WqUhnUuRLRHHQcUsh87Dc
hYobkBf7dQPIPfzWxVBL9IZwRhI3Y8UafHGg5ZYwY+gQSHFjov/utnINAbaWA4+G
UBYr5glrncHThOIgNnx0v/XxIbOFSOFj/D5cSlkLsy6piNdO7c8Wa0rb+w+r8Ns4
e8iIrHQT/MwD6IfkznG9KBh3XYz9PD7rnpYatepbtrNErfNjwCAicFhgp6jtBHWC
SztVS6jB/7Bux/QXNovto5YHirOALKEt+B6vYrE95c6cXVhUJNNH7sIEphsfnGuw
GwnJM8prML9cPjoxAp33tVlmGOYJk7qVcSE0jGUMTmm8nZzwqISImRvOa0rk6ynf
o4A31JBg23CykHO7ZxGbRZWfhsi+C53FeJi9EAJoBZ1PZPqQOpxYQVEjoruOuzm3
jXaizEZyLLh62suNHqArHr0sBaW3Uin8rVnC4bfvYkNj8Ugaz6Xx7cu8gvF3S8AT
fjHV+qtRF7V1UxYw7NNoEV65fgcqRT1fw8P7Hly2wtQym3PPsL929p9OvPJHsEBZ
vt6uIGsHpH3LnUm3gv+OfkihJbcfuVms6boizIMayt5v/aNki3D9RmcCP+VYTWts
QV+kwMOT3a7gQdD4iY7FpSOfUhAKd8IJt+5WaNz36QPDj/qWkegA24Dl6K9IOWNg
XakS8hTNdbDiSRwbEqK9ykqvdx6pis1/xlJOqwXi6FCm/xfFTFAwAZun2WnJZ+Vc
mAHB5cJ5AHuwJBIV2uYyt+4VrAInKWp0OiKxndRIVoQsxxqejqEDDF10DH6XOUpH
Aq5FMjMIsyB0wP3OQ5bFQ9PejkPF2qkpHPPkd6XPEHH8dlsuM5o6HtEtZE67qaXI
WuLabUtpMYcKOKyMSIdrzPuXJ3CTyWmvxPbKPB8Qasyt8/1qMSgT0sA6AEVaUL2R
QWskGrMNMS4AzC7QlzeaHKZ5jPu9Q75uEQNMIueibEeJDjumzpD6KVnkNj8Ala9f
0ryIZQ6SdTpqF4swgP1XgmVnYiAo2BdIuwpawjvhelPFfG/Ey35xHJbTwwBcaFIH
HVHmLBsGLBQpx2ot/PkJjePEEYkT/Jhzv/DE+pDyomIkJUDimUPOruuXYbXzLaxA
mJTyVevsuWtzDcLxqc+UqOHEoZ2azvDJlourotVLvYtUO7dm4RVBFHNd6CtN2thl
HUC2jUH5mafGatt02ALvzaG8kXcH8ShAaJ/vgZ/2b5G5ROOgwRpG7TcQVQL3h8Zf
YfgAUCozd+sAqRw3qQ7avhibUJPmnz8NZd+iof7DCvSKpml0XriCHgPLrbVSiSub
dINqNcSYap685cdbJTTqDrpHwq90o8P2YVrV3vpZwcwzFKs0ANIVLIZjsEAUBWht
8YDl6fOybvVyTAtfdGvmPRP551noicKATcuW6OjoCPdgN8tt966vlg5Hcl+Gpk9g
9ZYGUS8P24E0U/qFhrSkYZjCkh+HZ5Mcoax039U50wux3DVV/R5oUmFeSUu6JhNP
zHjbe6duMTRCaRMDRoPUI0U3dGBGLM4P7GCWGdLJ5RGzM3sFu1YkMQjEvVdTRdQs
IMxbD8VUT+6lQcISdewMo0TCD9x2BejSSMBe19mzrW9ogdYIdNBVADskwhr4f+zE
VKXFnp53Zov5TYKDeYdvuP9oyTfmDNAeKOqYso4ntNMyEBzqgz6x7rQK06Uwa6df
bNm8IFwQr3weBaskH73LhP+yQnBfeOcjqLnbRjYGVvqgVqRQN20gHdQQ/5uf9RVh
TRtBiUlLqN7myCmgzgcXA9kR3xEytPNct+OKo68elRO6n5Mllcj6aXRh+P25jy6i
0RsUkiUs2BP5FTawkkKYHRRAvmPUzx8YjEFeLA18vHO/qPXHv2oEANYz+aaI+MNQ
iiTBdrwV61+PSuC38cmWEDsmNdd0kWdDN9Yr2/+9G2pPDYq6shKq3EGwQX57+JuM
NyCeCmftt7mgZt62ji9fBVcfRMsmdpcRzj1L0gCMdOxoPh+6rGBhO15ylNuOZ3uh
CWtusSwPeFm7ftQ6AKFXVK+yAha2o+k7HEirJQMWUN1EzSP42ei21NfK/PEAFcTC
jtEOylImQ64Mh4cdA3p429risnMFgd/2t6A3ZcgmariGr2IuZKR1VskTwCaNW0pU
Xa4XRTt7ctAPYG/7X5TSEp7vd1WbOdLyY89mJSaObQVu9zL3cffalKnx991XKvcX
ReBGivQyYU/NSpF7ID3Xj3mEgDLmn5a7Nh4Yua4GimjyyeR6Pp4xabv7fIZhQ5IR
q2qC9LagDD0Xr6dDYOmNv89V2VAC6fioS4IjsdQL+hrH7Xwnf9czoJvdozYE4RTl
IdRQDNab5Py3YU7ABJ0jE8UZ4O+pPzkD+riz5eW9jNWraHIGn3DrU013BhMFqCPz
fHK2vdBByEOkvu330SRhb6BzkD7PgzXu3b0qaHgo8mHuOOl2rwkHHN5QD5GFFiZT
XrnJaOrdbDFHnvBElSbC0BrTaRIct/VjcXCuxcVyIDHbwYRtAS6rq+hgyin6+S7t
QTj/SGfjOQupOwjG924/OZLf84Ct68RcOzsP6Wcp3JXZaju0MO+3AKy8t8b6oA5d
zWtiMtTOEqFUPMXE7uMauoAncQtFJwnTWrveRdtPLAbNd8ml8DP93WZTjeI15R9D
fnfjCdq4ij3FAio19/nZbUJZM+JEuXYZwtiJU1HJvV2QpOJkW+FE0RnsbAYl4DR+
E9fNER0xuER1efU8LNBKpG3PE7+ahWPG4/NDbub6SLWgQ0zz5ja25yTQjTZI0cBr
R8y92obvbog/sOYGCqOzlJuC/pWLs3Z8miwhBpbtPAWT1AXomQbbZGqdvZopYF2z
nVSGbI1ulE5kUFV8ONQeX37ItPYe4RSZ4Ayjf/+SdL8ZyqnQqljRlr2ZKRZ5ln74
PIl8Ik7WqzSU5TCov04mL8OfjKiGNYIWqDO2cL3YV5t/EhMaAObjYYf64xeGivaX
9jxkPeXIJUbQ9/i+jZEVz0k1W5WCNNMbczt7imN4hiF1EzTshE6rd0JPvjW0Gm9E
zTNO3RgPut2OACelcT+nGyRHQNsIoMAZxk/Ys3YRujjPoxM1jDESFWnppZEVxqww
RVGcZBiXwszfOADrhjzLgLeQRCV0vJvpatmWF341cAXsd6IlNmnyfUCbcDUpd9il
hLyLO77T6bgqnh0jzzkShgpH6LA9IullFhiE46QEVei6IdUJUZskfFoaUMY/F+ng
DH1NLIzCDaTgXa6HSqBjFqqW6YDWvDbcLMzeYjgVYxc6V7/phOeLX+HG94X78jEm
wITNp12aqjMFViIVsuAcCWShPeXB6tdb5gdvJJcMOqYaqn8v3aY+j4yqGRneRN90
1viFRqJ8M9v27dNtEQNGEYTz/CkBrJbjq8gOC8yFjHVWdDKptoZUYZxd8jgnSY34
4pWS5IEwPPKHhIVvkb62CMiJWetdisWo0JWHENvyaG+d0VcAbSrCeDtyVtN3vda9
j4UWtLOQ66mpU2xG8y9JVDvCHsJds18cGRl6OrR6ZFCzNFQJd6AKdepModI2jiWX
/b1m1cBwOnb374//6/pUysxE2JDD38tL1Ee4Kglp8C5PS5QcjCRiA8wUomxpj/9x
lOgwI2DKZXhIP6WrNpew9IFjXS8Fdm4R3GpsbSP8wk0nTSTLDpfea9TwZO3FUzhU
0kHKzjNqMIdq7VZXnZarelIDfnZPF+iMJvIYii1KLSlJdEkBv1iuEDgq70nneZ8f
6/sZWPEZNEON7OA+oX9bTVbaIPfc4nxfdTHKKHxLjNmMcnKmF7vNz9kRJOg7RTzq
Zr6FdzhZykVj2fwpEAUA7ToTi8BDRqgbEaIg90vMhcvqyU/yOWWT3SXGsnuYgAfU
OkFx1I41TaR30heXVWhwuQ+tMTimjFXFl230Iw9Jb0wBa00Yq7plJiOueITmDOmj
RpvVm+n/0LZUYgJg/HhctiHB2pBWP+X4TlrImnUZJOvIS5HM9CSqYKORvKMcZ75Z
UBKsG8qazu5LyUmZ/67jXNqPxCAQy3N4Rylmm3ZZwyIboHvYa4ACz+56ERy/G3Ez
rOPkwqruUAjERkZ83xjdMziZ+6fYJwB+ll0qDkOBnH8ztSa2Vkfck/yoFV9gzpbW
WYEh6oaj1AIN55Q/sWMYyZ0fpU1WppsAkUPbmeNdrzbFatBaaT9r0TciajWdd6gR
v/a1CK4fZl5DltkKk7El8YcHkAugbWpoFJyLA6yA0Poj2BbTDymnCiKGch/YuGkt
nMh/zW7JD1hgZriJN4NMs8OQFzRg80NEzySE76AgmhQt1Wa5PeYKhCRVO+WUw3RC
CN1UIOUEE9hMal6ZeZ+cT6vazLZtNXO/pAFVC2Ey/cDGgLOj35RrM7NLlMdyr5qp
DysUOhimqjLX0xbYqsNnBt8S6kn2BPvi6eaEtedtta9amGm4/1hYt/5ZoSOJsbIe
kWz26qrEoXze76iP05LXCbXYuVBJqZD6qNd3VICgaTh7qKilsomk/MI8tucvD9ww
jlDom5a7KRPzUji1ccb0VH4tqmoCK2tWUgHk4dPJqVyc6Wlv2D0/a/+FrdkkL1UI
VG+vKKOLza5Ffa6I6fZTXbRrAAzYaqK1037fDxyONuS0QImojV3qvS1G8g1RDVM+
vvAe0WaciEgVQOwDIdZbVLXhFShFnpOCFQ1X5YDDP69vQTeng45dgNH9/6JZlpVA
iwt0xzguK3xyhnh83UK5jXejYbnL9TZ0U3wyi0I7pE7tkZGO6wTn4n1sYXcvA72K
m1SjDlN/rSn3nLjzWI4tScZjb8ULerxb9hVp+ZmJ+AYTMlhyT4l2G9YlT3J6Z/ul
8kqabbrVh9XMMwHuGtF5Q87IXx2mdgJarnp4Y8iQGuT7JCBsSIT1GJABRxPf+WUz
pH62TrZCj+VYQ9Rm1+9HKO21dWxqmKn/yZDqKVxDSGUJKa1liMMBhhSPnnSchJBv
geYdpZfjeItnmFnunw3bC0f2n+TWywjaM1Gb2hI5smQEot+76O+vemIDd9OjZ8m0
rL/E8OuqR8oHlQATbQGEGR5bABEcOkVZIP9OB37qzm92OQyZ0JEuAFjgHiBcFcKb
gF8vhzioQJES2lPmyOS2TJsJxrAVsVZwwoV933oomRSGVfT9pd1S4wu3caOIjiyK
MRTBe8pfRrMPKwdZ2sa4xXKLw3rEzLw8QGVM8AEv2JI3Vd+zt2Z67mT1VvVlLu7y
ibuFPJ3qpO+N9cOVxpaV3rI9RzJTdLhL+SRDtoJKNH1vmvF89cS7GV6v93w6tRAw
VN6T2o42jRfA60CfL7rc2mGrpynxqchWls7v35gdC6FS4WFYl6MrKOEpfnEHEPxK
ref/xGnQQ4iV1Df8J9i7sUadx5XdtAs45xzuCGpNcbz12tx5C4j4Gw/LL9YsRuuJ
KThAyMtSc9JXR+L9wj953jUbzufQlpSTOKpNbRLBXUeMAXmURqmX0Ero9uHAP3Po
ZNCMjkon0CvTmPUMkOJ5jvvBIRO5769nk9mdQAZcXrU/vm06EkTbHG679Ph/kDRf
nSCVRdXcVUytrmwwgQ5dvXN0CtsfX3l8B9LVKZwJBaW5aZjtsgBuwuUMXg/tlzBW
jKjnRtbjsp+wSA0xgjuneW40acZtZU/0nABHotqGamLO4jmrE1BGezKtCIWcl6KN
MNQ5Fk6dsl/wI4C6XgN8uJBIwlC//dr+dFgvOKZJ15VZYvNh/INryJtyYPFQ8W6H
1ne6DuGLocDdq3Lq/xSLyaVdo/DlvziS2O4J4lXt0rNc+7gPgzzA04OxxnAlFxiK
BID66yxFekzpkixuFBV1oRd1WYQPwHikpszQOg+QY+Rf6qLQtPfcjMJfcWzZB9/f
jWTPkz7OsFxjRsqnov3r0JPkc0Wu2FIzSC2vT7V35c3G8PYguUMmKyOOtk0Kq0kt
5fwwc/yEadXofEevneh+e35zCTr+aY+kJ7XU8+KjBH8oSCRTnR9ciDXzWYGk2XAk
e2sO0ZSBlQPuGOpqfEYaQeqZaPOxHuxmBn1RjN8JU9t0JBmIOsN0WnY6a0kaJEdA
8OMCvIlH0XpIpXzg2Lkt5S+GgnpQdSK15fGTFOkkwJjdEHslflPCsVBIUT/pyjJE
RceXptOA+QgibwCNP2uStMo0dKbjiCn6LMDgS+N2F9HsM/5gp01XEAQ1T+upXxkU
38lGlPvmQCBVh5nkc5T0hZ3PAi9+4HYe7wo4AVn3EqYkuOFUDETgsElLYrx8Imkx
NQfVK5UeUcH4nFV3wIIkuhm8X0Rj+1K1H3SZdfw5z50qv+NWsZmxW4e7QH+e+E+N
rtqZZSBWOmxth3VQ3aab69WgZfFUFnr/QI3vt56VV1HcqDaYnqqTb8ufOan5aTJz
29YYncvhhN9+eP4dR7wzWuNFKzXAqVq945oyTDQ+0OBETPeC2pxiysRCt1Aff7Oa
aajEgKWA0pIXflzizq7RhnCK7hGlygNnF4uPUJYW1WgWxZMWrdcy4QfD09mjL54z
sXCIPNHptXfv8GyfeMKkTowmqgTV91b1o5CTrgveGrLkWoqDc8qBFHJBct9Dtl4M
uADc+qj9NrEZhzyYyhWgrOrf6+fW5+DpMkG13rkikF1Sw6mlFMdHj2my/No/NLmH
ZKSu5HmRPM9rNSTljF3mJqqLsuZaa9RVvjWF1SNeCVyU6e4puhKn66JTzob1xi05
V2xt8u8JefWrcuk14kH8ejTkb5NoUJ7pXA/pCTuXkD6CERgo3ojq9hf0+avfuQNI
P2sCMuGEToyY9rDGLjJm5RVqOEnkn9abeZUTwRYbuOR09MeZIYZIqeu6ATLMRWCC
XINMYJRc5bIoR3erYQCPmcl4SX71yB/ru6V0791/A+iLSFgnnprsWl+imq/qvNAv
Oit6zSkgLj8N2e1iKr52ykuOfz55xX44YuLa7zb+xR7b0yKMLMPYzwryI2ECwwK7
K2TPG3qrHzUzQohckSH1dBZCpCchdUNWhRvnWhD3Rm342LxMDWRDSFV0VKvFXO2x
SwYWW2iJQN2zzdXf+YQ69GjmYwCRC0CzsXGps56dm/jG2IH33ni0PykpQOwBSTQS
773Z9XrrA8uBYxSYdgD3yDhLL3R/hUpm1P2YkSrMIf2h3qrhLHG/pI0vs7zCSdHY
i5Id9kiBDkABu0UE8V/jJgTO40KZ+ss6hTYCHSyc56Z0rJEAsbgagf4UCSg+9kfy
3A9/kVF+jO5R18u2+hVWlXor7gZAyNhXzqdxBmMmaF39J1Q28QaiWYFa1FCSCGED
cONYmZ7ZQG3pFW7L7gUC88NlgV7hhQPr2IbNhEng55aXBeZ73HeZG7dbkaYVKxBm
FBGHBM75uJuB4fgospWmZYWLOMjf5hrZHdwOSv8c6VWb63NqzTGCBp1D75bL5B+F
MNp8FQ5F41Ot3pse1Uz2IkVHJQUTtNixiXBDIbXuxhIZhTTCEiZSohb7zrzcwJ+f
EuM1/6ELoLqQV8FI7V8fvX9e4UINLx9CEZHymFBuOaBKLg8L3Itk1d2wDnhGwp1Y
GJYVLSf0iBfX9XH2ryPySI387AV4cOtoGXQWvyckr2oDadGeVhQI8gEyou/gxR75
T3zXXK8YubrCufkNdLQr3WQQXd0bHk20uphtOi0Gg6mxPMLySharVFspTB0GWlM8
uXuK8EcI4r8q04dbQpGOGZFZp3PX6tgMMD1VcLZqQ42MlF6l6nV14KeTEVO6Fx0C
Dppi+ERoHyVncKkgQG+i99QfXXYM/QyBFXaRHUAYu/OLRm476DBBBOWRbsEqBCTN
TY28A7c2BbAyVvOw3jpBWBE7l2m9H9YejlwCDQiaB564CsCiQSHECFHlQhg8clqo
6rv8ud5q1v8KzejoMiv8iTTFvxUkpHL87SLV0G5mh4UiZkf5tMiZ2slTlZblynf5
BBjZovGnJnVti/k/rRZVLyxFGGxRBmhIg0rRByN7uYbWm+InHQscF5soDuDUjTaO
TTezKWryksf2P62ezb4zVqJd0ooz4v6fMGVHrgFdTSYZKKDtHLz93STaB2ij1ESJ
qAtSismshEaVijNjYDf3eKWUkflr2k133xitM8vrstwqSBN0+Aa29jVo3yuwhu6C
r/O0DpKuR2m7RBP/jZNb1XlrpcMC9yPT5bRS7qGTLM6mly5i/cZ1Bm14aDmikfwI
dZSoIFGfWFVWmCwczC0yG+4/AtMtJ4Jh2IkmrhyS/ErFWvIjKi/EA0BnxxQrINi3
bjsAylRLzwkZCrfFyFswEC4BS09Na6RMQibRtrmDnFDTg8+9j5ZJW/siVRfsgfzi
vt8ZIlVPFiuRkxx9F0eSPMWnMtUezWUGq67v4hX3+40/U6gnpwXr6PlY6RKu9l8Z
4DYTZKNHvY/hLUQmYMRu9tuGO7/bDz3pSKYYKH9PUgcnmDRb7wqtvnrI/S/Kc6gs
44MFAb2/dBiN0lBZIrmGuKz5Bu9tw2IEycY17gofw7GQUxrqXecfYxejDXSjt/c5
PGUfplP/BEaLXWGQnF+FQr/opaD9leysQxtaYvUeMGdhhnPglifsgtGuMp4dcUjX
GjIqrHsayRY3ioY4r9J6qE6n675F6xRSzb1a03gqVTiHNp+CKV+ERdkRXC6Gym99
h5+bk+amfxZXFESRyGH1Q0fmH+q+GwmfCI81jQ3TLLFqxDx5bUaAK1c0q2FPjQ+0
ol1IWI6jkG9qmevoR0lNCyVa2NbekVQnnrceswf3Ze4ul8qo8tkTwA+4kWB54zvH
VPH8Xm2/eHSIgvzyOCT+/ibqP4ehb2Wt9drrnJR4m60kABawe8lIxBWdXIudETew
m/1F6f5I7BKsnDSRfB+f3ddpFF4zV7YDD73PhmRt+QjyYLXYCYRuu4oVmVK5VsmC
9rnMwk1D+ZionJ0wpdcymVDgdlvCPhZE15+9BcbGbZb8YwBf/UB9YrtIvwsrkiwq
ZQAPn0+JUgaPb8BRuU+TLYNUa0pDLqFHr2JVzEO+mwoxXPXO1+p6DHsiQN/Fti4r
NhIzhECpdLFSFQzOxfY43ddkf+C78cEq9lwgSejtDRiTvha2bhhLYPQ+J+WcPCU3
8QxatH3+XoQktBbHd22oSMdJ1cjp0nyRORpjZd4KnwBDeMf9jnqpa5J3i2phyFKR
nwlI0hlhP1Fns1sY6gHbgyAmo31Uxq7l+yxOJzOB75jEIkAfJyd77rTJzLbRl702
tBePbPy3/nHjx6A3Gb+VinSElH5IV/dTGr7H/AaE9Pbhalurpkv0FsH3Pc9p6uNI
O/Dk50o+NawxVU8bZehzwASELDWl5jaKPraWgblTGBxp85VVUKkl4jCwUNa9NBb5
qLRGjf+p1yuZUhnh6WJUEWltmMjap0Eas+qGQ44vlLEMyUS2iQDw2pRoUd2CjufI
qEXpNDeuo06w4CpjsuiLUiWhf4au8zT9n3LL7aWX9QjTQM0iB+taxA75l1eU4FIu
ThAcOwp0LX1yZLeN5RcOb8oEYPw4j4+Vlgj7bzjrFaTF7su6w/eapFaN2smWJ9br
Qol4D3tsnHWjqApyYvYlFoPjSpuMwk2e90CGbdoQJPxAxGHISOGIwsLT+vCupQ9n
yv9XAI1bI3SbKK0AJ3AIUFkV+ml58JK3md1/Tt52BY2UCz39JvP4YvhEiOlvFEHw
L0pct4D8Y+UH14HV1aJaXlh1QTNnBrd8k4wZUDu2EMsw0AG9cE3oCRkSMabte1EB
hqxo1ClSAjRjGt+JeKxkxsmiKJ0i+4HLXd7B0iIK89nhsYgmQMORSgv9sXP4Jr5I
RPMpvBMNax1xTEgKECN3k4HI+JHJS4ulKrBdaLEzjIb42/8muKIiHAwhtg9yHcoD
apadDet2TOpfF+SHTcI9PS2FiIe1a1t9M1t0FfAW+JtRDe7Gsay6vwME/gBb3zbF
lS4lRwR7QIWWFe+pjvkXDYVFPSLkJBUvmn0nrikMvlsoutH5+h6pVoAb03SZW8Ys
VaRPm9ioNL+tnJ4HD038Pc+6O0R6k0q1E3L7Ohh2/pnop9dqQYcKvqllST9Vv9v7
NrPGQog19tk1uGBfF64RPis9Hc6Dz0ui9TtpGleNhoweBLzveZi2HLPclhdHWKOi
Ftbn1JMhmKOTNy7Md3oApoPj/EWfbdWgEc3WDrEBnUIGIPaVNzPDRvHkS2Iyx6vU
a4Zpo8ORVAzEzaAcoSMRAYN8KcrSSLwSP57NVVlzto16/Wd6/XRl8vMETkmwPaX4
Q5OGnZN2Jw2oeqaZlGSIp3y7N67+oUKJ9nSqkuuiyGNs5yfJXxvyKCGdMwhTnWcG
NWNIeZtivxyYAnaqGJCFl7Q62oH0tiTPJPYo3iwXQBFiDwVxNbruPL5ouslNpRRO
/JNtCV+U2GkNbidmvoZSzlW1gBblC5OVHM/gbr/w4DaHIbEMm0hU1VDPoI8P1uV0
dHeR10i2GatEt4/qTtug/LcOhTw7CI8fpq5LcVTuAC6cBwpSitiHbbLu839J3BE4
rGw3GtadX7EPCbQwCNzL+UXvovLfONLm/blBxj0ZmMggq27EzRy15vTcGnOaFZK5
91wlMc2GPfdCrX0Y4ZNhsXafhOlJBLqUKNJyAB8V0yjwLsPsteCXaur5jxgk5Gzv
agDX6/LunWCz8dxNHU2zyUpox2UYO1Uc7PAMDZiKkcpU2UgnPr9qU1jrLMAJrx7G
InHEw90h9R+W5d6NSrKQcKT2XdJ/h5yi3NDjPMaSUEcbpT3Jdixb0ygneJrBO9A+
/HjW4/kRz8P7Tsu62epDqnQe9Z5LFFAoSR5rACc8UVnpP6JUon0nw+JAAxWsD4i2
csF7SBWdgyr/d5RGf5DrVP/Ug32Hm/u/QI3XbHXg5TdT+PMJxcikFDo9BbBnf8GC
bnUAs9HtPNALQKpG9Qzp8VH8Upy514ITjtNRPjhKpjUii54ozi67vnEHOZ63og50
iXJ7j4HOxSyG22NNU9DYq73IoN+O0gT3mMuZRbs6uKz7frhcUQKcr/o7FX98bPRx
pxwf+qK+9iSBZaID0RFkVgpw/W5MW6+il3Z7nvmKzcGI51RZnVakthZLsfrAs+Ka
5bBGIdFw/83R14m9UZCgxYQ3RjkbNC06MGA3T+/Sdyyo02VEiNTh6pNdVo2q+BL/
xhS01y36bTkUfZwS0lqo9uh3G9tdfy7nDVD/5pAM/47n8Pndyh7CGGjd651hzMPh
lW1qB7PS5dwvulXIuzgOP+bJMp5c4eEkAThTb6Fo2dtP82k6ODR5hUAxXiW0hlY6
MOQdJO9O0WRtq74LSvUrDA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
emCVbMmoPzBUBen1ql1ZaDy1dd1lLxttxvAaSVKJzcROWVCcgM4F5sGEj+jcX6Qt
l/S1tpVPW9a+XiYiLapmr+5gu1HzQh49RX23fegVs7+M6yCbwVIldSFHHxrLUhhA
M5LBoMDSoS593zUYjCPI5R1UPqIrQmi1/S0cUWCKlX7lABIPRAld8ek562CBmeRc
MoX9qWJEG54l/kTLJ+QqYzoLtRXch4bGeQDNIcpwnmhnwmel4aMJD1wS2mTdSyPL
6cfw4nhhxfjlaLMSD10Kcib16SRnEymLxetd0cP/mhBCTfuLeIHuwLndf1q8dCNj
3+/eX2JDDw0TMiLASkc+FA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2864 )
`pragma protect data_block
zN5ZDFSZ3Ro2UZmhMPGHDbxTGwP+HNlSNP8tb+hay6+qJFZ8dZibInkP3aVahaiD
AedQl/XXntwa+PWgfJJSsoF/z86zaIUUiVCfZcEwfPB9ZBq9sAGHBatO1Soq8J6z
r7djCHHoLyYHfOPoWtqfWCLvcS4aO20A+LY6y4Dci/cpyz+QStnCET6SiX13NiFL
2GZ/VYb+8z4mf9saq6d5BWzYeZJab+lklsn/4cMWs1y8LiwPDD9aV/KTHJWrCpT5
MIgnkfwId7rXPzazH21HSgrInRSDl9CIr7uubrEPc/39vUUNLtVT3eIewbfDbD1G
URxxxaYc0wt9xTX4gZIa2W/cDDQTp/RTEXipsFhKIM2uhwDtu14Gp5UI0/rSz5eZ
pHDMU8COlIoRmTnnVbnl+SCYOmT516p2E50XmpxkbFhwLcSd59hOlErocigwKp5g
NLiCHMyyXbdIkYlNcosx/y7e3+TQKBlFCYCynH820oire/c9VOOEHeYGJ69Wwtm/
ZQ8IOnZT8jfxB7+p5wGpE9JT4WZUtypX5rOlSWdasaropKYfVP5+hlC2Qln8h+9u
RGDS8nGjKJ8YQBicfKFfbkOl5kpAnQzVeantCuFXg33Rldv4OVPmArjeRRYuIODC
Tf0h1wIEDKEbpccRWt1/Epj40+MWD3W2vgAY1O0Lxk4zsWTLu4adjdUufIfMmGKi
0eyqkWVoY4YbwXaBABmyIR5MWY5CkvJ/xaqcKYNWWztvoD3D4CXVfdVR3jKxVwYf
r4HlUQhQqklBaKjBzC1lmFIHSg3gmW6gx4xgcickXnuiwcOdXZ/mMkNaGUrh3zCx
uwUYQXv19OsLvayhpq0u56iUNjx5qCbGFy36ZapDM+ztuYLkMGmh5bLehJOcX+ur
Zwcf8n9eWfSddHffaWJxdKSHjdVGU/KGeDYFGm0cU5OqB7HVS1nAWqw8KAPa4GTX
gKz3CkE5VPEVEU5cZe3EsisSQ00ZFVl8ZKLLAkEkie2fcpP6KEF1uvPWFRCXaeae
MEAS7g6pSkuxXfA0LTbe205I6+I6hi38D+v7S3o8MeyqtgoGUZ1c2TOqCqoYGa7j
AXOMz7FbOl9zDbN4c9suseDohN0Su3KDxjZBcgTaxdW4jILN6QYoeNIJ5VaFK1y3
oAwTQ1NMXSh4BGUyrXAPad2ppyEWZroFubh42nVbJhtF3AlHENSL3wRgfrfzZMDL
3hmsdtaF6Oesx/QZhP9GrSmjEn35hvQX5w7vI6VdJcl3kVM3siyYw6ol5WP5QVq7
EYetgrXJcaNpNgj4mZTJuFLIhiy6O3Hku61bnEn6ZUi8vuv/fHPQIq8f7ipGk3O2
CB7RwPaDFnETNYQOrrEO8TnrBvUkHC68UsbHXcwFazd4B5S0MW+rxYHvPoBCeuTZ
0h2ntqdf+OL99rMustfiwNdfUhCp/YOwDLX4/OnwoNg04PaltPq7BRsV/fB1gq1T
5u78oQUgdx8+xRSIsG42ZQHTUGwuXXz82N2m7IzPZiN0PQYwrfWKyBJup/8AC//r
t4AmYKEG3lG5lF1eA43ACGL26RIKkp5+VivIVFkbjMGT+HbhHFodqpnjhrClm7Xx
L8HNauYwUQql6oweczZqgltIHsJN43uYPKhcq3B6OgvVnG/vtgpe1Rf5qJUP6usb
kVEn1jh7cpV4NRXczbj2P584gggBh1k4hxnzLp6wurQ4VqtxIJSHnZg26HgkKcZM
UAPzTphVBXtwHXLxNj7YLVadYVpdkVuOrHq1NBqvzdIa1JgVBGubhnlWEAux7PEU
EFzJSgQd2j63rRGVI4GoOtymwTnt/ZXAoexlxyWmoqZM9TBuzpbUVnbyUDJPnnWz
O+eByN7D9Lu61a8uD2Dq+bTfU+LyaH05A3JSU2AXWhamauwP8O0QWtNTXE2rgYDs
bD3bM+l7O5sfw763w7m9CAxtfR946EKm2obz5bULiEuhIPlhc8qPkZYqeHyovSXR
dE4SIfeXDoLiZXrIJMAXz1jcuhrlyQyY5VGb/dTQPJLcjcjN+P/K6iO942PDVE5h
DmDxLi9vLRi4iMeumnyD6ULmXup3kfjWhKVOIyXBJ4XTa+ZpmmyUfAS2f9clDVmw
PlBgISkXndKmNIxmVCbtEt1YLgmQTc2XyxuHVyvrzA9AmGfQjhQ9UPzPbdrt7Kah
qrVyGBaSA/VFeq64TyEm0q/P0F5vHyf0ZeqmggFOZbL6M625GkgslqQsrCr1HFA+
anxKb9d2iWU/2J687dU0Y4cAkQWBCzQeaybDU3igZk2K1/YCiGkFBt/ximuEs4Z+
SjwFruc6Fm9octBkLo4EPiK/9aMcApghIZodETLU7xnzq0E5UCm80UuMuJuox9sd
mUPzDM6Lit5OVedCMMjlLYmy8CtBr2boQWndLW2iXJbQ9VkFaMxy8y09e3Hy4wAc
60roiipYOXEV/zfrBa8zaIq+5xiGxw5oKzZuYbs+ztozEJ/sLu7ZOMRdkn6XBpQU
PhwkvuOi3EyQrgVR1nILJ6TXh5pCyf7Qc+/7YsoPfjON7xygrTApWyMPOHqMmL05
pxuBWdOAvruo17gK7LAkbG6JaYXD/mW/c02EqWniWsL83QAbmf5Cp16spxzA4Owy
1nGYtHQdPFp2T/qbdFrQ3WlcjbnOw1T8LsJY4RXgthTdrKw8QPe43PU55v46QXwP
++Zm2W/aWS7cG5EauaeFNoGNy65jbNvWIhgFeAGJQ8hUBb+ud8rBDtqx0lcs93NP
c1LjqhtJ+LowKDHnvpnZht9l+XBAc7Qu+MQQGjUeneueJ6yiXCMeEZk4zV5SDYfU
/Wzf88G7fvIfctZ1hTL0012mdn0WPcaJ7dtfjHNCFr4RAhu0gQIMOayBmlCO9Bz0
xDZ3Mjb/CxaOwflOAcwMSD6qALmxmH/hBlfrt9qF9JkRqUkwuseLw09SmxMTcoaO
BIWwXXISagqQA8dhrr8oiE2rpvDo6BOPtZqDbR0zXlzuEPdfdOIl3qXTdCcQTI7D
drkE4486brlvrtjJGuBJRGKuCtuambFgrfNLK+vaDm1cRI/0mWG0zhVxL7lCZ+om
P74dp6ogPE8gN64lkCUzFGW8usSqPvpBoplsg5GC1Z3SaKm261eIciSPl/KXKXro
29/AAouVV38P7F8ygdaZVgMJyBYgHUFX0CRhpHoi76esiYa70iXhKAsiZeEv0iKd
NIt0LqClGrmssI+iulPWWotT77Q1e0zYYd7OhEo66LA04vFmHbq665ZmzU3bHLTl
Oh/BzmFt1eNPqoXbBJriYzzZbD3yIToprL2gGR4G5z+vgBlXtWKXiCIs4vwb2TAM
dnY7y3U4Eana0G4JMunkV7F4iBwjqccDf10NNr7CDbp6vpp53jDwJfWqIVClmjzs
F57c7QdDK2RTkN7gEpc3GLdSXCjmcZ3JMZhx0NXOvKDgsWW2FS6IX8LilfN/+VsJ
Z+f+zy6sD2phNL4gXQRI5ETLmbdzZ/BzPVOB05i0Qx9lCNPapgrqNL84XNiizTSv
ZCMjb5LVwUmWtiXbSCxfgvR0KoN7S5avx2T7HvoNiH4+xeWuCKqJIFYa0gBIGrvJ
uT435VGFQ/9tWoXWco4P7uOc/EDCHRIfKWF7zr6kRm6Eg/2IdywLzvrtJ0TA8UDY
2oHWbN/i8dmk26LYl1e8EHxzAZXBpBNhot4hdkhvdhDybKOxzUH5sLMP7IeFwzMy
mksoaKsfwv+N53/pQ/HnuPF32L3u51p21Mo/k36nv5IkugE7ToBFwqftrcPVXkLX
2xV1TighUlLG40B+5l3wRwBHcqA9NpN7sy/LykABRr0=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
QctDQiF7YRNyb6MTDEfgr/TzgQ6eclWKit/gFok+Vty2jWvJlVyRxW9nFUjN/nvv
BG27pgJsqx0e6iFs/6SMfWpncZOtAUQptjoP4gDyRssvD4q6B9ZKcNqss4ymZdni
7IYZGlTMS+Q7NCWmyy2VInNlq3m9yt3Z9K8B1S1TfQCeju5blLeJTrXolLuwIkgZ
yJEdrXKGGXyeVV2W9fjwongSJl7gcxGjp40HGSdkykYF8uYMUNYPC9SSZhe63YvX
psJWShdUQPh8AtjLgcLJ3Y9ZobTcyPCkO5QFqReVy/eZHE8o0I7fI/7gS75ATOJA
RCaM+hMfr0d0SsmR1tg06Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8720 )
`pragma protect data_block
Ejd7dZI+XjzJw3dDfmAHcogR50xJcFRumcnYanZPBfAAPC7/Sy/B3r19D9pWhyoA
gcxk13fO2uOFW7cQhf57ecgpGiXkU8XgLhCGIqSeKmpfXvJ6LY4xNxXYJTp8o17q
V/4Dsv5d/JXN6vblRO4Nn54HpnJZIgIE3lCnRpzUCkHW/6PS7qDM6pZXay9i4p3C
7xBTGJNQ2WINEuWnGFPOXQtOyMic4+0IBGC1JEZmDy9Tv0Nq+QAwhfnsbfn8uzBv
rhXxOgFjvpZkzKn78kzDepT4B0now8FfRCwMVj7GU4y5X4JTGMXJQH4ryDTDi+72
y5LNta3mfmg4AMyQnEHG/AKyq8S5gfYxm71s5GHeaM4DZt6dHLD9s6nsUTBQP6OP
ejCNasqqsHY5rzcLRVmilWWVYpNrWsVlB3dFui8C9MuOWiG7jcND6rdruAnFBeHL
FcGh1VO6DqWFrLODWJYzLT8ws4KUG/cRi1TQAbQQKCcEOi7e7QcAK2/mVEyY3Utl
QKt9t/9fDYWAydkgZMnDJDH6TpK9ZWzGeZpM6m/lRQ+959Y9FTY9b7sfLrzaIdSc
hgPBaxBh/tsl80zi8elleHhbF1Y7Cmw9iyF3TgkesdddrM88HgCjyF8V00tSC8T7
Mw/7itPEIUnRQIPWF+ex1SXifHYVemQv3O4c5BB5rF7WLfWtXN+wsjC28H16GY2e
qYZubysCuonkkiM24WNhakIOCKfuMqM0E+5OqKu402gGoUlU/wogWAE7yrCYKCUI
016w4/FyZcsB6C6E5ysgHMl3XO8EfWEJ7FY7on5L9WZ9amwG8P9XeuT7XBAdOyFq
LLT20xC9BQKCwZB4A/PkDzTUEwmXSC/gGbvNOxh0P2lJuuDYkq4lCfldT3lQtbCm
bQwHzVRd2s3WbSQ6TpbAhsN0sCuL9shCCVCS/1xsvOejQzQbJUuImTn4WHX3foEB
ZYcQ0N8h4Hss5OtTMHuInaQH0lQfe24cXY5fmYVzghPLt71FUFEo6cGLXvnoocxI
G9sNtj5T/4pg0zoXza+w80JBbfFD39RNc0TCUgjh/F3QlNwIaaf0hiuCp9XkjBxZ
PJ2WZ1sHBqWLejJYDxkQRVMoFZLGytEEtrMcohSGia9lfG4OW5n1RBvPrDjLHvv5
r+J2BouYLa2+7SZ2dxh8UpgdG20fSw/R3YrYDCelHoxSN4kfH+/7nBWPkqU7j+Ye
30QZuviDTCxAkJ644v+QGWulAFYZ+Y9rahY0HHs/f7gr9HJfNOPAyxQ0J96StyTd
WbXt1dnvpYIHCEilSQBsscFT23TwbDMAWWqT3wvP4GGBPDubONH0S6af0JrxyKBj
PW5XIlEHkJFBlfq4LVEsVJD2PTFBnWmj7XJeMz8Th+svTx52SDvyGtcxywpz3Xut
2x1LV3IhMrsVAWrRcwExb8cC1k8ee8NQIH4sFlgArlSMAZ5hN4pMhWeUznwg/2Wt
WbXYs2uWj1oRxKoak8kHHCdoxfjv7KJNJTWEQ18wNFAJwhuGRuIeRSilcONmhVm/
0JCvxkaAL5tM0/onU4mcoqqOcjkVx+IThjhuGVSZ8fa9QnDYjmpqBM/XgIBzQUNK
3piAE/i8OW35KSrxS3pgx+5iaumqJRq1mkxyftO0AFTtCddwhsCaGAs0eo0KVuRe
SBbR8EmZesXG5pKrKhs3Yo3Tm9hsEUjhrULm5gI5mHpi/fHzI3qlveI19TQCtxsd
2iijNRrryl/hAPpPgssW2a/q9rXfrrk60bA+JbEn/tWyilSqDHrM/YBQ6oIZBUfK
nRgTPMyLRXG1Nsw5c6ckVh+WLzGUim5zeC1pX4W2VWDH2qwn4F6GLyN4IMle28vO
vexUUpNPRmPtdN4Qdx1RVyrPJiZJ5hukQ9am4zt+hwCplOGjVq06OyDYbRMXb/k2
ql4cZ8L9ZoL6ynq0wW09+Wjz2Heofx7lLQSB6aXbPtcauugupAl+/6f+4dCeQ3ez
MT4WJNcYovfM9JQqiuEhtJcqaaMRTsjkoTFSUZpuWeCd9k7mmwin0xx9uRuAvoi3
o3M+zsly6u8JQH3l6tM+Kk+8hCXolOZPzS3ezJEdO7uXja70Ju9zjZvuV+Pc6G73
lpKqY2o1v4esy4KLipnzapEELJSqUtoMD67XWMVCT9+n+ZUtDSYy1vLXTC3ItDeg
FoXls7S1JLCE4RVz4l8C7sVOwNjMFt+ZU75oHX7wNL/K/0gWDES+C1APA2qXQeM4
JFIS8mSSK7JTyYLWdUA0k1dJTQNf751Nl8V7Raym3Al83g/kEEiDqn93Yi+zUdJu
x8CScVUakkEWaSu0kwlwoWwgAoXD2V631yAaQnfyyASC2pQwTQJeUGLWInW5BWhN
hnCtKEfIxlh4Nu9mxcPKGBj2dUTUyYN/97qv/lM4bA5rkUpPRAyLdC3dnI5x9yO0
VyT5R4FJFdcbtj/GsBq43MoZYO8uR1iaVz0FZ8/a0wg8SMz91lhMU5hK5LXpWtyf
NS9gN3eT4kAPx4UiLM2NEa0Q6+vgETUIOR7CyMtz0m8Qaqr2GZxZrRc0kqg5kXrU
2VAB2YOp6457Uy0inYhuSW7k+veRE8eP0cgXdoxA68/eZ3Rt4+c73bBmS4ZHTkpz
vfF+HRDwmBkK1PV3Wgu70fiiynwDRS5xPXWu5zI1V96TnbvcQQMuYRVNhovNYv6p
wMqmc06tO5o2SPPhEl75cRPSX3Kk11tNoXGdj+7l/CdRVppwy/GkYQ5yqWFWe0Bm
NvA5xHfi8NDrJmLqCYtYJ09d36nXiGG8c7sZd3r7xvd4cm1AIFtklPj3pX9T38WP
GZO9TD9izKp6OS82w7+lhfBHe8gXb7vI1TysbaZICltbGA3/1a7LV1xiJ0ULm3Fy
AJgxlm1tSArALdHDH3oDC2zgxNGOvOInat4zOaPz3Ie6s9na557sK2uTCvwB+67k
SAeWO9LSSrL9uzpmouuIfeYrmJWevUQBYNxjiBdcdJ7nlhU9yxsxjtcvB0dX98wT
d0+/Eqixlu2M6UzyMezugrXaTXcwQRX/RQmXFPO/jDX0vOZQo6WJGkI8nhKqKYC7
2Ri/sIrFqskdVF8JjFGC8R0WIewKEZWsdvBg+myK7+pSVN32XJpSxaUe7VCGk2PA
UG5rYjBetfDXsdddDGxwz1MDhwUIwsFb0W1UVeJTHaM8ydYJJy1z6d3SmzRB0Vp3
w4lJ2pgAEBFHuFiJpO17AoSEflZJ4lyWYWLnxM5tV2BrSqqZRaJ+fllhS96qtWpO
zrQk/U6nPIQmWoqUjSz8Af+wKQY/jNEZoNGEJZ4ByvhbqsOHaba2z8yIvIugcgkK
YRYPPxSDZHRY3QV+vSKTwYUkEYX10Dk63HaPFiRzxu9VXRSJUf+yeLUcwdFWF5oM
AqBRo3gg62EscbLpiiaswxzPLnMcEQNlWWWHhH0FaRhC0i7Lntko7yp+DgWqaMKK
xqi1L28DdDYcPwXqT0RaHbyCMrjfmx0i5WdluQk4cUzyjbDDrD74nQVp7mlT4Bia
nvHq5dY80/gMwQ3KGQglONykwDYJZkZtbne1E2ElO6KEOUC52IatW9Q+Oq2iZEDt
YXf+pz2A31T45h05zt7hD7l8FWHnFfr7+krUnYUmV8S/UKoapHpAsEE13tJG/fpc
4rPvY6YYRQBqA2uo8qWbwjMwbn3RLzoklj49khsf00LaqCOk8iG8fg2qjNzJt7XH
bXDSvvUTFEWrvB1Qz0vbaka61+qQyVx6DPHk8ju5EfevD1J7fLF3f5nESy2QIywK
haroiRU0UzNaiGPGuv6QGNFUdPpTRtsL/sgqfMUiVkjuk6mgjN1eTH+jX86wHKkB
9w120KXK/SZisRZ/i8UuoHwPq5byLzkgyWMGgmKE0oxm2ervULAgH2MaY+k/Kwfd
7VZGwDHe1O3msmHEngltEGrSeZiiu/F5t0d38yJxE+Bze0HLqYZ8qHxWhYHbgb+s
lMpsqQP0Oz3afrIuPgY24a7QEik/REpIjOaO1bMqSELs4eKe8nicWlGy+3+IRVxP
Kc6XHFOdDn5kK0d66i5voTdVQLniFhnUcppIvoCPS6h8ISRnsNQkI90RreGgTxvj
ykJqNFUivzEhd9fWcCUVJPSpQVyO8R9EC/yiavx7zj0vTXFPZrFJRcv8/NJg3s6F
XdnjHUgN/LRMqyoM6/UWkJ+/11V93fslWB1H6tfze9pez1rtmMnSWFKJY2xWbusi
OrY5iekuUPK3Rk4DfTdOGCudpP8Veh0HNrCRQNpYfBlUnPLXXSs4cqyeAxxvS+Ux
QGnC+GdCRRDPDEm8rCYiNe9wCFmHGUnfwoWwlewYJLVfhVDEd+XdF4/Cb7eNtxZP
1G9rsIbTa+VLOV6V9uaUhyPU12Bvs/wUyrqQNxpBDaJTqXuFu9Y5s8MYNvW0l9sk
sy0P7qYb2Ho1UB/dsYqf5DyX3yGYzok7xOmZNM40uC1nQUmDChplkzSANaXSuXs1
KF1hyFyOXRp4EwgIxlEfJb985QnqvohToJCzuPYyeS3bDrWtewvrypNLsoT2feW2
QMGlTJB4jM9FpdYV1TO+hXNo7r5v2ZI3QCKCTcx21QXcmhk2FVl9DT7O7tzpi9I4
vmWc3qjtGU6Ku4F9oLSBE0UAT47pY8R3XHGFNFA44r3dhwhiyXhCLJWFV8RGOifo
5XVwj6+wz3idZE1fORMAE79/I9azvBn22usnXF0cC7iG9ofP9CRnaJ+cmKIFSCcU
PCklESviiJeImtZnAxy1jvq5rO0C11f/YwEduQsHhz6PfdUX/nokraFOQ5iqVgkV
8QST1lMGxdO5LJeIw6Dm+ig4EWuf1pc8tIijY+TLKwqNuSIiT8DjyYD4A0jGrYLU
+STR8t+AhXWCzwsBjhLWqyjd35aevZutU0RJRT0iwR9bHWbJhVjILC7J11jkwr3w
UwT85N4sUHrCJISkptNU5vc1YTgkAqpHNbjhGpahUuC2gjaJNek8BXq7x8JquDPr
Uaiqx/MMhQ854EBLTeQZp+dK5caMXD51F+itAYZg8RMTCPOFo4RlPD/ZQUEMNXvl
1EhdQ+Y/INWCHgiUkcExFNx8Lq0iV4dguOCaov8sMbqoxS7CoNaNOXCNAliKNPOd
ZGFw7rkNIhYlouv2Qrfb9TG1YZnqeZDZlV6BTvOJ88YZcDjVNBbquhc48q+XAdn9
+hDacRMhdWY91OrK7Xy5I+BYMTx/in7hHeqDO24Ultx5GETsV/+vocaHDr90zqJC
FJphN0ySZRUlzAC4Fjw50Ddr3S8Bf+RKeMysrGjov7lyPfEMjQRLp27n8sNdDo3E
zvMJDsDlQ105Xrf9ZIG6tz0Mut3YUSzgNsSq8qSzr8ryr0ybfCd4MLanwV47I4f8
TrsJyKygyYdJqUnp5dllfRQ/fJNSLz3aIOPIH/0td3hUq0BsdFytCplIb4QZfwWg
Dg2LBjt6swhxgWIDsYQyPSlMP4ShBlybY/ibZ2FSIZmBhN9Lnbq0YrMe0h+wfG1s
yOyAHwkplvmI0K+1jiTk80AMGjq0KEru0JmUs1FlV1qXFb0Yc0Trcelr699N4OFk
erbD1iiXs/4n6AoWoac+zUBTJ8bTLK7fbJ//cipFY2wIi8HkrxSIwnetflWxjc/D
pbQ/VQx7HHEqlOR5pMgpgUo7fsHZwFDTPb3IL1PvNPhuP1o2960TY26RhICI+wwx
k+KBpY7OhzlyUUhCxJpA8YcZrgxYK/9yX/47T7LJCQyrBDbULyP/zAOPjEQ1E7pe
L5S+99J/LlI93voOCG96IGjEhcHK+WiI6Mhq9IBABXETXondgparnN7ZL3ogQtiv
AabS6vnk2aEwWCbKwLIGszYlfg/zaUJNEJnJN9tTFtDSMHGA47iWE45EZVABn12+
tVF4a3A/e+rSX1GMKLUVGW7wB43WEjrFA+2Mw6xa52Mnb8sS6JKl4lezQ6HowXlF
BBHrek45rMqdYR8/GMRmfpift4W2BJxcEqDCY9YyrSqqViTFTyCqLdiFzer4oVWk
Cw7s+9uXQOE9bEyZhM77a9GNCxe5OIpBWB+FDATfqECdnnmcrF9G6nFg1XDFcu6L
CA+b2HxgsZKl9A3hchmnKYVf025NX22xULWNVDYHfnB98lR+/zZ3VwUT/EC/ynUS
Fkq2+C3nAV5rdeoXmasoMhaNluqjsPixXRCv8ynCtHlyX2jxIElF1FvHNz9aMyZ5
Tvh+K00yVnE5oB4t3Y8tQOLhdD/I1ccMjuF+LTzdFWQJQ68k59XS5YQ5qdaFLutd
JbzSKyC2mDB0iKBF2TnBHtHWt3nyDFblkB+Uef61wdnKY6e7yUuujOYmjLCGriC4
TCCLfNOfG+vtsUwbvoTRCeDwVfAS5rLDFbC8sYbixkPPt6xODbRhl7xiPCTEnuMG
s+Zlk7t5djY0e3bJ2CpAYYD3EeNjay8h3BIKFyWuxpa864/BhK88y8mzgE8217MZ
o8eyKYbQUbDNGfgZm5OEJB6MPUF7Fmb+z4kHrASzZdC5ZKXY40C7ZiUsF2PseHQ2
TxqIIFgk28UfTvT0wXvtbeykk7MP2eF1hE0zM08lmkJpd61A/8+mHJKe+SDFF26F
kYL+e3ydJUy+PKGw+XS33iXVUQn6Lp8Q/jMCNs+h6li4ykt+XD6rfWco0riJbYGW
J7zqpmNLbtT7Ep1Rm0XZlVjASb+AfmgykZoEtDtI3fbpJJebXQ7qFNidn+MqOppB
ZfK9N0DIHIyz7lAE8ohju07TDXJKg6XG/MZtEo72dDCZuNW3GIJMhB1fXuRFB6kK
5TbhK7Sni4pj9b5rU5zhoa9gBLtNpWYcJkKZcI+yu6GixomHTx60UQQ6ZlTj3ktj
H4FG+7vz7iQAtC7cvy8+gLu3EflZhX/g1bJBXjkCwknUhR1sZeMfwBBEfcccO8sY
+C8nXw+rJsLEEWGYiwD0E1pnqOF3LsO1mvgC6B0wY9uh2epWkA/oBlchUzNR2094
vjETj1a2j1cuXYMiWDOrreoETJOdhV70+9jRaiACiuR8du/td/GW3iRZ4GYsSAQh
yE0Dz/qKgtxkotuUHkqB5Ewo58AYKEc8KPCuBu75juhXAxN4K3XLeSiqJrB912X+
Rt1WQ6ddbhvLOblEX/dMpfvnvp3VrdtauLi/zJyr2yWxE8XIYscLgopNfgbl/9T9
2qxsd1VjTP4uFjgtFrO/HWqTbXhxYaSbH3PjzSQV7MqMuDSAKsvOwWyjJl+qm6zW
rRPFeDUoQVpOjK6J2wHkz88CONZkv9B88zZExd9DX1qZbi3oN1uS1OmP8iAy9CdW
VWJs3IvJDeOO8eLETKn4ivxVceI4E9XTqdyiKyObYQKQ7NSEcshPdlCmK9DFZxiz
ouQXaIMbsCU7Tf+yGWsJI8ZcnRrzzJLGn8QatKbpTmdxRdk1s5R+usVK/Q36WtF6
lt3jV1EKpcn0znrHOkfgR8rvDeEO6o7FJsnvmsEdpntonuV8eToshbxuJvkUFzTm
oXEdnU5Zkpob+X5VMRgQhbCTKJQUxIzPREwl5Y6vZ+L91/nzXwpjFwhR00sN0A6B
b4Uvv2O5y6oaKV8L8Tc+xdoOwPJPvW4fwZ7CzMDu0i+S19aQkhDSN0Nds7bE+FfE
797r3Kt5aJKvJZARYi/6NW5HxSFhR6EiQyuHL0AZX1a4/4j9lTdt19yULUBVYORE
3hDxO16Xcyc/upSWNQ4zHG/fM4x4vz49l6LiwWYljiyuTMVug4C0kHBnoCkyn9/J
fc/uGmoYYl7Ix+nSL9z7zQ0sU6NumEGTfk6788hVGorNsJv3zq/p7nba8PA39xq6
ZoAQBkexqw7qSFpN/woQPtivtX1gOgVYLB91YqPauO5oOCkt4EueyYv0ChHTSekw
/l7rTqC8Rq15Dn2awKdmsSKXRDAV7EIDQUA/J+qO0/KEZH9XHZn+/U4wMMLhfzFw
sEq3pKMJJXJ6oxpnT5/FerAZuwQoNbVKPNGDrZ3y0kUnl42YJT9MzUMwgImKlTVv
XEXHS8UFfLq1Qk1XTHCfvaITyDrM4r35lVRZ9xGrQzTEqUW/juOzA58dfSRhgkZK
dJe3EfkmIJMMzOtaNAP7Dangh5AtLveSYTqvuNHC0g8dlAHjtS6LFS4pg4t7C8LJ
mq7RyYLKKZDs6E8P8KKOU9yFkszEMPmAgbXXEALQg1e0mMLfpQJ7Gw1v8tos2R7w
nlZeS1Ah1TZ6r2nYsIjh5BTLZndRheS06/HIjGCIvadX2X+SRFY1/eaVgaoX8klm
T5HtQZBbUu1y+WUaWpm1PKD721GVimkJ/dZKP8SPH7Eqrxehr7x3WcN2PB5u9+Bh
4T0Uf6yIfSS7aUvMJMc9zCRAsfEU65mxhAcfbvaEwyAVIPLNu2x+RV6XDBY8c8oG
G1b5MW/uVGy/8dX7uhAHiOxgrMjb/4B9/2/WG+Sqsrmtwr4IwSC9y5tB+GBkOYdx
0vJ7aMJy4O/hjcCb83x4PmZI06dNBOodfGZ+f0UPJGLKXPRduAzXVXDpUiAPeciU
l3erjIerRpeyfHCfHJC98OYWblVP52cGJx0VbhzTpMGwvHpNQAFLmz+ZprDiF2O4
O3e8QlQCLHd7Wmu99uKd1FEUKbge/0OJoZkpUGOY3+2prxtKML/UAgNJXr0uKVkG
jNk3Qv5TaXNsF6gAM1aoKbA5l4Vpu6de+qJFvoQC3uQ/evbsbKdrt/MmWa7PudvJ
FOpzj6u2zhHH+EeY4CuuI9Dq4pQAJWASdrSA2doq1oNXPetE7Rwz97HlQk/KYLuP
kVac14EhmbZI7iQ6835CJPXAZx+pGG+DUAzXIeF4CVyh6hOJLev+iuP6+wPBN0NJ
Uw6TXawfz50gU+dLMEI1mF0sZZQzZ6KN30TmFlSyAxezbiE5vg0+ALhRwXGcxib3
jNxUrZAxfx+cCPvtLxQ3R3MTEm8e9w0wQqXriHNAP0kwlE/Bm6b+NgzEGHUFvBBk
njmKEjmARBBOnIInv9IiYRMXTZGmoprgPZtGAHr9zPVGhe5szEqEVX96spWP8BFf
kd4LbmXldxhLnBgXgun84a1ehE89IIV5y2dgs6ZVzIXahUe8GEG0O7u/Vjl1mCBH
IxODDEtwlhxYHI6Pp0e69/BUBJaxFnomIyBlpipbicvQLp/PBwYxBv8SOoXvJtP+
i+FuS/rPSmBaXgXM9WjbHlBURJ1u//h8BwxZv1ghUtwTGRVGu6nmQbNVlYS4H8q1
EJbTajeuay+UlMSBeyE7jLd2axZVuJJn+gukZ/nh3WMzlVqSAjeLHoYy7a3WUiJa
80u3zhA+dG54RmEN+Q3hM5K3VIpPxwp8aCNdw+UO1/1tQIPILNA9AbD8VaQP39Oa
lBzxsOb+bNhjpl38YQR34to0UYOIJQDvj/AS9xhRrn5/cRoIN/lyOcIKLxpsTcjL
6C5XMfD8osnQFoeV4vMLrj6qonTBq+sity8uKeDElp007w4iecVVFuu6MabrjJUz
mV23RO/GxdL7azg+KoY5NYujo0z9ABZqMOONah2Y2Xs0f9DgnKxROzrqx14R7qsv
JP+xdbV2MfAae6SJTFhCBNDOovS1yv8nwC0/Vc1ZdX/qY0Q1ASORwSWy8hEIp9RK
2qNpVOFhdFmVjW7nVByzFslcfesCKL/Od1tEargXMHR/4jqD/dIB+8QEabYeqCxM
k5mDdxXS40RVtC75KFfm/5i3kCAXau8AsuJvBvPU5H6XaYA/8L74q1j3XuQ0AsYp
Nphh/KZOzFOOdSby6tYaGtkRU8JZPYCmSFoLRfI2YTwlX4ddEB3OezEq/XDoalag
r7O5HbIN7CjaeF+y8KiUc68t/auPGaZv+WsEfj8rRDqgSbGg6rlasCG0sEprt6Nr
0WCZYH9CjQVAZRllAAmGxgtL0e3pkTcRbGTYJot5e0cp7XrRXs0qxMGSl3XRvhzu
ghQNDNw/TIlyATt+stE81b5ygoShbpJP3uk1VCUqLe0d9H2p2KoxfBfVhYOkf9wB
m1PjXlWJQ2YeKvP3/Qgp4KNMKkhrLxbd7i0WtHDy6pg00D9JaQ0yXBIp03UFfTug
0oeoCJ8/45fNYh9KSpzKXzanl4IRCzFvLTaIBfffhWWEJ2SMz01dbagrfNGEm1Cs
yU5lTBkbrvMU+LhirG2Z5iLoVVxAbqUPTZfhvNlW85mJSly22puiR5a31d4LUTNa
oI40Tr5QbXFAjgrGHzCaMmD3lbZiBRWcdjph2cG7Unthm7pMfYjRLBzP21N1JINg
wv6gioL2hHugMksBiX9z3vr6dJdFxxMlpI+tBQMXSG1BbIRjnvXVkEMFYnVC6k5H
F/4A311H22Ov1sATi8kzX4v3MA8Is5sp8F/LtDpGU7YMkjHwgA6/bi0S5nldfm/p
yGfb+4gyt7erlLaI/J3UTX574Gn5CcXdnoqcT33w9qVCDtiZrIn8+CThHCKLtqlD
Str5K3dl0kmRdex+5dEQCGNL8CgRDVi2USzZmzn+rGLeKe9iEAGTDgCX+UTCpdMb
0gikmhzm1X3nM/OFWsb6bU280g8fCg1dP0BD+fVJn4L8RhEndoWM0uyTSCR5oNjK
1N4tRUIhChqopCgDf/GLK1oggHEuOlC0MLGgbu9BdIs6BaEy+q6G8z0+PTcBHDfu
q/lsb3BvQzBbQKFIobJbGhjnq0NDSwUqYRVCrlDnD0OAf1QNt00xcjT7vtDS8xQz
w3azvTbJufV1KOwrzPmTMrkykCuCPQMkg6uIcGrvBCEWS44ELnUYJr3d0E7mEJih
KHwbw+H4+1HdbTXmkFxTJ90MmWzQznyp6DtLhVPJU+IpuKRBsntzdkWyp0l4+oBh
TEYFQNYIwsPfpDrFqZ2Eomb7EAtk5xPigXaRqficrGw+kh3O2OUH0aMdNjHgtJ1x
KhjfeT2Nk0x89Jwj6J0miEyLDlSRFlw/c40lCnokBIBG3joSixBEiM+z93IGc0uU
Za+vUMdZPka5825R7K+bjD6E5+D4Fsk+yu8NP1cFhiE1wFSNwapj+gcIM5xz1PdC
Hj5Sn3uUez5U6cpBLmbO6YRFK0YPwYK0xjmjEVL3JJkc7bzp7mt4S/SYjk+qNprm
9sWPb6179npT6pKbp8GUNZFdIvp6Va5AYTaHASSo1fFhLhKeOAqV69P8jUzZN3iM
bh/FNMsI+kzZK1ytJi22rhA0gPfbJHOyjy6NUwIEwvXRWYiFvE0JHexSlXj1HJCp
fgwmHoWxAvkFAV5tz+qie5sK6svsjNGIovIFZv6dUrEKzE7TIHIAGCspFdgY18E2
MNvLRVe8vJo/bX98J/EuhoMQtq8EKEXlIgS5xQnnumBeMrpzAo1reqv1paRszXjm
MQcjP/5nPsBWAFHY927G6wWjUhjGLFNShNy80KonzgpFU8h0iOHGLtlebAaeOUBM
4NQTad1g81GMib3ZQLuqgFLsG2Xk0qSdxDVSZ6HS25RfB+pudQVC8M3MOPgiZfiO
WR0Od05A+5uAf7lfltvYo+CVYNPbopOFHSIWb6HMqUAJZOWRsoLKGwzApba/VI7Q
mP0ljntQw5Pj7O7iTIjypvE1CxWJD0GFksHj+KFslLWhYtWlTV/kJv+N6z2gE1M8
47A+bzc/dOhti43guI3AazJ2wyMSKa13UbHfFZoK5uM=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jkjFHbSEUarmPdvQkxC+DrskiCFTI9UR0OEX8DlscF+78O6l1OjKrIsVWkxqfo4K
OzywOAaEC7krunD/fw0C7HXETnloC2JCdiRd+yzbAKHLSeAlhXN3X5R7+Ce0l2Eo
yoMvpVD8Rdfjh/NnYBR2BD5tcMJG/t1a23T3NeuJuHQYrLAlUBD0XreaSs4JIh/D
unFK6kXnSY2GBxp815mLJ3qA7QPOLlsipgacJG7u3txECd3QGwpzx1nObHyPWPTz
fzyoajtsOWivxP6KoQtoo4ZACT+q7qy1KPWEUsKffSimCW9NNneMeajRAt1h36JL
/nq+8eyhTjc4pkUFwQgDFA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
qfOGrHoa0qlElsTrWihylT7j6HEoyYOH4fmkUfOz9edmN/pK0Qtv8PtBIP/lK9dN
TICcXsmH7sWdwcYoNSV9Tmy6XEv4Wz7ncxP9IehxNVueI/sDLON/+f4XEKJSQQaG
ovpXONHk/hAftrnBdYSRYw2knLowiDPbkIOlQeb2KyKEbob840yb7quX1DlqPxa9
UZEWS66nZOwllwTQHgHKM0glAVi71ls/51sCtJK29lEoZjcfc1jucFfrJR6TU/HM
X8KH2s+zC+9tOVxSSfx5mkfiVSFmRFHesL7Yt+7J57jE2clGEHz3RfQl7ZWqIQGg
bA5lZ4lIXxzeQOiImO1f+ZpGANDxOutq689ndBvSRyb3iCCFO+8iS3G3opvHDjhf
TBagteZSFCfgknZ/IuIDbTYnsHn4u3Tccsj3LselzmwT7Rf+bsT+xGw4fnrcIQm1
XDYwzpzaoLr/Dy9R2p+Wlf+QKS3Fwuje5/2nP/wnIq8wXWobQ/k0oCFLKSFBur6c
FN9FyZq64QCTgx01uD6YJ3mNBtbWNWSSgCMdS6okqsx1j16ryEC0zNWn/Z8bVigY
cbHcK5/qL5j7yt0Fvya7inPGmEu6gVWN/OJU5sFOe50dVXj4q46t4tU+Qa5KZ2ja
veAfPM/EYIOW6lRDwpoAuu2Z+2qAHVqVykGeX+62pZPwSMBnrzfVgkwfB2uxMHeI
tSUUzPNvSaFCrEVqVGeCLSkSqyMtTeS2GBk5gV2TIwoAvuuwDGnlXFMr6CA3kO78
b50u6J3i3i0wiO4yq1jNNysPFO+0JAtMAuHGvfV7MgGK+RopOW/RG4ZxWVhhCc1b
uMy68bTzrZRTwGwdvXrZ/Kag5/39PFuHuGUzqBPeUUtHwZQrrOIte35q8TuZXOFe
v2EAN0BYOXV4z4z0A0qpq0FJI2jkOh8pOi74LQ5nFLqK1ixiJK/cnbV/MfnP3xJo
RQ4Nr+raJrIhCXv+tQWDQODXHdWTdlvQBymZtNOc7zNLteH/jL/mfCRUqe4Ubz3I
FCjcRh1t/fAuGYdyQktQ5NJ9jLmrYGwneX4j+h3Rq9eynMsuqSvRokSErypqXEEF
5ykN4c94yGIBkCBC41no1KxDW+DY8kA9Dgzgm2z64uJjY7Yk2CeH5h5F4VkDZus0
CNHWqZ08xFifLM2E9qhWSm+NFwVtuRCG3KOMEupdgphdkXodtVim87C0yewUa0/Y
zEuMqO2cmPZvH15r07JZE60Z/0V9fx2IwLiEb8QsSk8RomWg/19H74cpcpUtSbcY
lIWUlAOzN64xuLaZq79kELgQH4FtLaZQpbS0tswEfmkGTdWuGsuchNfWIkR4yJXN
IIwo5zym9niU5mijXd5IeHcDLRC60MzAVGM1sX2waWHbbEvSk6LQALm01WqaVohJ
R8atViVfJXZVNcHSQuc97rOGdda3FT8xPGPV4G4inFS9xDnAm83/NN7E36FuAEBK
XlC34We/SW1MFTn4ZvwmOjXQjp2vbyq30Kd8oDqnm2ppuf1y5n/IW1CuUMbD2lfu
NiZlVZ/fWmfb2Mqlu82thSi9+BnoWjnVdRImdoE1eD7hZ5gQxXevspmONLYZ+Z/y
8bkHdN6jJMH/RXNU/aQRvDFpDjTC1k1Fc6B+Fl1wztDpfauMHVQQpKNyMAvVNorL
k8k5Sjcdl9xttVem588kf6nlAwX6hqRXHCBvwRiE7L4n+J2Pm1/iSed1oeK/EwJY
sAAgwH9wfBuavP9tVHMwhpXLCgkubWHJuSfOKF+sctd3ph6Qrnsk0OyAl74OTc9a
onMBFEDmg6X60Dtdcb0jrtiIEYRVnraK+fgGauM2+ZiojHDMGfVDMQGTm6xgFFIZ
h6tJVk1W09IYUWBIkUVIow3ACp+/jnx0hGpED4M/yrw5AorfGx3Cz75UT34ntWWA
Nz3xt/RrODZo9wNxLw4tf5CdwO172sCU4ZwmUYGM4zRNu40bN7vXE1WEFk+l/r4L
GH2gQH6SKP1Hk0fllsloUbLBXJmbmpGivMRtuuVC+JqAvxALZgx7L6eWSxcBKXBB
DbrUOwFpZnXjlDtuQpO+NaaeFpXxBwLXz4womCqCJ5MBTLgyyzMGh8uXKcxuwBFR
/P7HqOrzBe506rrBuMT328OXrGw4DgKmVm8m2gB2SAfHpeqUBJbuYXnK9O1V75rE
cSBrGEpecD+HdHCFFEJosnztUqAhq5VeD/cswTT1vH/ko61LOC5qU6jiD2aBwNeQ
sHn5Fry7hSl4kGUQLPgVRQ3XZqv51HNCFWtFgqmN+GUMPREv7L+tMt3yKMT2E3PS
KEeWjAwo5SH6uWinK7WW6G0urxCpW2PCj5f1Uop2Io1PdMMkEtsHLHvvmcUS/DI5
dr9FLc1S1/v9McHK0HMV8jvEGKQ5XFrnJftguR1bXybzfCNH0BgGyG4j7Dk38JTU
MOqw4Aphiy8hapxfuL5wsJBF43nomNiuGXwengvTg4xcCMApy3LqNv/d5sRTUw0r
Gzn0BXXK8/lO20UkIAabagBePN+wFYlm+DVvsrt5aejPM5GhiQ3FOqRYZBy2bQho
QZK+ZmB8daal3ncsMDG860whwHbWp6whhrvlKon0PmJIw2vsZkNxqFjfD3evUGu3
cZg8M6Elth7siigaYhvl0HiEGayr0tfZykhSW2PwqoYtt9YTBHbmD0inrWGyD2GQ
Yv+wkccOJIxvMn/KJYOUQ/85dv1YMFmxWd1uZwd5NPYRtVlvaaiNVb2GOOqEk+he
VNtTS9t3jPsP2xJCUh1NTfIhkm17SJuPw6d3TsIQOL/lk6fraRyhITbwPYLDzjBg
AuKI+yNFkfVbQPh63jnI7xtr8WdiKO4dWCv1PwCwuqCMLvy0PklKuVWQWNDBCmKW
3yahzkBsiXkjPiPV9Bo3LHtjY9r1yBNclc6J0o6vfTx6kdDqVtUD1cOLzvkHLeEO
x58U9OMCSQpLgazV207FBVWuvRiikPOqLDIR+u/j6lfK/hKmXMhubJT2wS7NRNdu
njzW99qPab395c/9rcmbuBBJ5qLhpnChq2mTlv6Qk6b4KMRz8zkTcGTlBUC19Dno
XftI5jeQ6Xn1PklvUdf+WyQpfsiGPLwlGE3uVN2lacnrm4vEsxM9AhCKOPONccds
/Jof0ZxkkIPK62iCgXVjeKGZbpOHp3GNAKvzM7X8tySKZxmnr8eWI19fg05+NW8H
i6Zunk2njqeeib5jgshgq7Ueilj6yBPO5FFLh6ujgiXmQwFKobzYCdYy7FRWin9C
lbwDwXRYyABEqqzAOPWV/4VD59C+nIC7JbrZz26d4Man2Bb0oeZwJodSNYz/ews+
W1eNxgwzAUm/HII1V37vh+wv/femzKA17KRF5MCTX8AWqBFyrUh6RpQF7wHd4Nc6
o3m7uEZY5v1+urM3HBauAUsBQTUsLW70+NfZuRbeF/bIc30Gg+f41mgPR+2vuSay
Wh7UoqsRCQztFkvqwR67lEM9kG0yqe4k+FwQrETlWCfP8+wFg9S9/oe8KnhbTMTq
yF6P9AqUQouERAMx7HoLgu0enCyJxlUKnlZNVGQY9UvDDe2bheMADXZgWWfACLRw
hZi3h0tPVPvYs+Ct67UCSkh7wswSM2W9Rb/hCnpQ+P5MdCx042Yrm/aJfJIXjMSZ
MUuHaqcW8LKycTDv9VPh4wNJYIeRmJ+O4OwDvtp0xeWThj6z7Apaq4QBFlLN2Ha4
CpaPeh+IXW7KDbIfz1TwEtvZt4KcSUzp0DNW9QulR4MutfGObhISw4bd+FwJ8hmB
ZSQ2cMijiCuk62nMzdenSW+NvB5I4jJxjlM9fZK6Ccg2+uHgYh/KmhZySIbGKDL7
eH3ddlJRrhFMJ528reN/g52BB9KvxgAoyCaaOTQ4qZCVEzi2ckhATm1fcbe/TmIL
SoN9JR5bo4Pd2xVr0cPPh2TUK2iiDOGmR2/sbgx2W+bAOLU1AucgI5pGrbdMst6a
bttZnGFgnQnX1KA9TGvZtrxeD13DRTG0FzWs0LNGA0p5cPE2Ij1QpXh5isuZhFwg
if9Gtqj4geaqzTGUH0PFRn5qvAlPDoD+SnFiR9Lb25lze2aY2u+OXEBSrMRkpWxT
Tz6gRMVvYCtlpPxiGl1B8ctm6kYvq8o2NLfZNkvT8E+WN0MO3Ot9R+Bd0uy5MNBW
PkwpPLnGxdmp9Aij3rC2n8iRp4FSeZgPbfBOq+IkZ7p1n2pz040ZP4tOjaUyGm62
Aflm6NNyV7blppYkzFk06Dc+5QUsb565aWu1cI8UF9Q0/9eZupPbUQjSzK90U/Cs
3ULvhbq5ctN47qNIIetSKB/qXom8vlHreEHs3+fM1Bo5H3SgRNZUxI5GnxMGCZuk
eR8ojqxDnzEgoaW3nw4fH90vvddd7I7RlzBfW5yKa1ABQIgJ6+JP1fA9//qiLTSH
/OD3WZg57g5Z/ppfiyHJDVNWvPtCZoOg4mWX9XQYE2VqCim6l9/2PUd8vPbgfZ5Z
57f8rBLENue4VxXAVnw/Jy5ZSppTyZfw/FqT3+GuQAyZFiJ9CRuP9LQFbOjWVkNa
Ra/7iIhnqDb1QQ8x44/U/w6ZXvcQo50ZF/h8Lyg/ndeT5hAS/vTbvqajXqOJULrc
y9WMih1tZ/EA8sNqclnvn9er70uuNcU8L2CjykbZbsWw9kB0lgToEtE6pAzkPFDx
INAhZnsuXlPWzRSBOAElmc3c3ngsFbsiCESnEYDsf04qi61NKZJjgCn/+OJXA/rR
mJsBc7hihNi7fK3+ESYcEIN84nJdJwqqpc2YFUTNNkXBwAG8+k6yyb7tyX8Ooxzd
rLPqkkJWakRecUskf/5IWI4hG5g2pW8wN5XJ8ACcEZPC/dVUevbLStupQB/2tODC
/f6cvtpxLhR8e1hfdSdloCo9m2QIRQ/EfCgQjuUXlD+cVctRxGvCfSy60G5VWQBp
ddTtc55WkgcI0Ny2MG2f9auAdjks1EpcTDnIamKIltEHHN54SvTo0FF3wRGEClvr
Pv3ei7NN61ui9MtZH2yPR1teq/u7Jl5OIQlz3buGcZOT4aM4KPuF703nYMcfAo9I
5qAPX/ulQT0IFdv9orfxsAExlai2VP9qb8L1Be4T3unOfEPKsudNKWBv2eLs5eTF
IZFvsOVT+gecZcWGISvF7y2EOfRmUHC/sB0o7lbfhpZQKtgiPZpActlomkPLQj6T
+BntfnKM5EI21vvGOBeqOwvdJ+/YE7hlVVfoZX9cThfyzGfg5mQVhzXztgxsti13
JvzRVp1GPONP6CxnN45GMrI7166c4r4usu9EBy5xY+YMVd4uvD4VU5zj6pLQbt0t
MvaegSv0+DoH58X8jdWUSBqvZxzfzM7cZkoPmp2zY1Fp/CInzgPKbw+Qzy/cNJGc
jJAPnKsJ5nh12jF3bDbKUcZUiDhXGIOoeKDLLZcXyMm0ia0qUwBNEi2fOE3bgaAp
fdnwmU2OsmZMjkuixEyA0VSnBu/t99I8sVEXBgrSXZN4Y6iLtY0p9pZ8sqz3Dv/c
qR+mkKP73UYiQ6q54cv2icx4qNf0Vxrf8w5qrfQcEWq/2/5ckHrldHUdGlq6B2Ja
M9ocZnDPw8KUPNm/RznuhnTMhqrUZvS3Rxv36RAgtFmIRWe8SRxMCymDM0myIt6s
PQ6V0p+9gv/JW1xByi9ZwIjtSvalsc4PHs3WuWq+SA6enFFo6XArBMSdIPfesM/U
En/9sc+qY8iZqi2CLSetJti3SfhOYY01KKvQzCOLNu2kGZyLbrxsitFXWhe6CluB
sQssszhCjXjlBATeX3/Mvt9dAG4XRdoWFBDyw9u2bu2bi3ng5tcFzmQ7rezrSroG
K8CLKWYF/gmY4VUaci8Df3Rk08iUhK3VsmnKAivOlWwokZ69VGG7L0eRcHH/f+zf
eKb0PJqIBUg4pPIv3n5Cv7xvtq/Eq3kDXGL0Fmdp9j+fftpQ0aepiCSDXMqkPdma
IFvnIwnUxlOkppbqXYpdUwKAoRqGIoNWh4WnZjl8rpcxiDjByef/Q9LH9fZG1z0w
sJkB8yn3PjLxx+9Hk3NxO54tUsOjvFRby0Kbm5v7zDdBdYhYu9RUJOmJ2I2WWQo7
PgnSZQ0IiMqZy5KWHAzlWvPoWCO2veEFvcejIWV3nHw2yDbSXbfxXGxe2x0QPxV8
ZafawDemBnTQNJQ+9Cp7kueo5nv9CwnPorJZgj5vaThe6M4NSWs1BAHIlJuqoqFz
IyOXGcRQGVETM7C2+mXSPrPrw8uB8vM16uhIKZ0Jtz6Mh19NEZKeD0QDFEURkQkn
OjCwe+2ABOYW+4CFfaQ7lU6XI4w74X0u52RSHX+d2sF/QY3fUBLzk7uojgHBJMwQ
cbydXIL1tiUmrza1pxIyKLXYZza9lrURsDk8Lap+SQvArPOnqFeH3Yegb3J9t9hk
5l0ZQJvgX10h1d5HBmq71dif0z/4M26fsOefAsoa0fyA7kr3/PRMIzDbd0Ih5e7C
FIfdBty6H+cMuvcZYAzySPlggjI94ugeW0XyWqxGDDroKrfj7YeWEbSWTwh5nMCO
VU62XYlXFi3j//oSrbZFoUjGMAVQyUFghIIi1/k96iZzf8R92dXbonH2/yVYrlVB
iCwIzHY1J5cnDS3Bqra9FYu/pEkD27nDu6lkFmGWql+69lBIBZfvNFNFFaUOT6dI
8UkpgYCamf676sGKKrEjGOjzqv3mqRWavChLHPSVp1dII73w+K9gAt+t1kUmN8db
ZU1pootrroLNNWammGmFb8ifDsZ24F1hri1CnZNZAWObvYonuv8a8pCJIwzDo22m
en2/B8JLLuH7mFlWvSBP4Gxc725WbHnpodJJ/tNsC6jpJ89VESHOvw4iiSR2RLU+
Ij50iLy3X1kr8W43DzI9DVwDWqygPkVdvOc3wNPKbekEBhJ5s1haowNajCP9+6xp
SXlNMcR78LWVMCMsZ319Fdpa9envn8qYJ388WW1z4Q9cw/2gtDpEZ+OeQD7NCSpj
eU3eWK/eNimGgiaYc7ZWVFIcRwRJO4YHqe3ghBJTkq942/caPGVTcegooVHx8w9y
ECvoNR37eF1JPn0WnOngeDCjNV0eKAL7CiU3ftmtMveM0mG79a2LzRpxyB//3mw0
7ihWXBV/qd7w8yXc4o4Dyu48zCMhSzgnvTSQmJtqBWOFdyb63otIIX+rpZbTazdi
GXhckcYJMj5PnLvCKjJYQOxDbLVRZpe43NXYj+2Lhv3fxT9UqQF2kvkF81GGjFP+
BR/Hzhr4O3Ng4W+7c6QqauzlHyACcvNMF9b/b+PzkMMUaDYIDh34sEqOLkcCT0fb
Vf0I/d6jZ5ZL88bPpvRDNQKAtJ/EJvPDLf/GWp5B6ydWstgC5X94pgCK1FYaQY55
LYYzfzkTVqDgcJR30nlImfVyTbMp0K0/aQmAvHdhXEPj8M3gyR6FKBYIQ0IxKbS0
s2xJsu6nudRjqJ+m8BmevhMsdoOlERkDmvHYIJpv6yxb4N8yeRUlCmYx6kD9ZdOr
69/Qrs/3q1ykgABFkJZjJFGL+R7MWxxaXvubOOptL8pdCVfCZvGC40PyxEEHJShx
KaNr90QlGAzhJf+2IlIcd3QmNDkQnM3QnN4JqHPTBUNQFDDBemnUNLF7AZb15K39
UwkJIN4eaq2ySC0ggTHqCAcbW70MWs2JogozAEc+6JEP6ruoDEJdBLfBVoZ8WwMQ
mhl6VoRVJ2oYA1qVFvDvtioIlXeLfvp8z39t4tD01+L5mcKtvtZEjFvBhla+7u6i
ZNkT5pV6MmddZ6rhm3CEntKCr1fB/nj02FFEKQevqxxPocGspifcdNHN9EewuGRb
B7BkBBV5/vZkndzLT09MRIBeQJjFevhvaErr8gK8LI2OqZB1/Jjq20dYHbSgl8SF
NsLeRpbAgmZLwSbzxntcVbF/06kiMqsNxIh6S0YSK9EyhRxWzYKS8nS0VC2vdfjM
ne/SvFwGwY4HcpH4L25+V7euKNPExJLk24P/okZmz8iKl4re9y9V399Pc3QDJbik
uZBdHgoxor9OpINCC4P3G4I2ZIGy3eWz4FeDcInehC9jTrLJJN1gMtzeK4lByaah
zqYEgHhsFnR65XEnE7JXOoHdirXq3FJbRtNNjeQwHG9iLBwq6NACPjyroucY7W53
8f8Oh1LX2bBF2zmyKk2vHuGkOO5oGuGBE5Vfbneq/KU8vWp+ieR1gI5y0GOmEOxD
DiYoRRaZXw/X3B7O/s/C29vgPmRlE8icm45xH9HLKMD38/rh6vpsycUP+7zGV+ue
eLc00wO/VHW0pV04kifVQdAh2zg5XyGWbXcuauDZ/X2YiCnFdDB0AD5wSmTIj7y3
LuMNOpdvrIcWUwH/yGpyUFItPgkwCn5pl3VcpeDmH3p9HXeQh6vD3iDdD8TNZG/E
VybvLoTwRmVu6sxe1Nnx1lXXesN8LNMHrDyt1/WksWXKDKGm5M9+7pUJgR6X9CkY
J2rzGiRk1uH5HGvBjabFX0xf+zsH5UtJZipUJh5zEwN1FSArETd7KlOQ3moSy6hy
mIsvRGxjRSX77gAqwxW7ZRcLZ5ROWPSmv5QJ3BjGgP/eP1xLJGM1Xv5Jo+nAssLV
tbgQM5Lf4KMwdGKMyFi/2xwvs5owS+nlRSjRVXfJaYMUeBG+BK/pLxUVQQniw0KY
WR1QAorgM5V/Z6V2ru9I/8oGNyJvzyDchKFJgG0nb7kJ94YJTYc0i6KAaN1MGWwf
8ZRkEvx6M8NA0iMe501dzyaHtf9wggnUmQXdnW/N/cCP8bHNtkqUYOXR8iedh2E1
8PsJsS8MrSZ0FQFLFBJezUzozaK5NfMaTOdcfdpseTLYlYyWHHocZB7BtmiBNcQE
7xmPh907HJQBr9Lj3sjz1qVK6BBVLNdNgkte0SzYcDr4nZMJyjSuGjJkOSzGb/4i
AfB+SrWE9ZQnOFJu1ZmPxP1pF5EBHOwot+qezF9raCPTtivv5aC7QoMVmGrsTHWL
8U/BsRhFM4fIWSbUtD6jJemFKjWyK8XGQhYNIHPPJK8VqFv5BKtHNB1XADWGTj0U
dldMhIFtnDGnTen4QzgEIbsauPmEqTBeLtHHjU/DwSXXyz4wZ6WI7PxdLuLpFSYR
C7vGg3XJ9EFN1P4VgEi3+ac+8E6zfQxV7armBYro+yNEkEtgY46Y7C6JX9YODRWB
tb2Ke7gsmDPRx3bhRk7fMVnbK3kTPBjLnGinN6CfakKYWjTc0VYWBnNRJ6txqmq8
Tr1SZPLtullMO6i98HKPYgzkYlPIibZJugahzr2NOwOMkEhuh857nKAMvddFAfKR
RUEhVDwcJizWsxu38faEgeM3UwOaHHZb4epDd81QyvAyHFF8WjVgl0sRtt+ttIc9
vc5GSB3tBOaWJ22yhZRlj4/8csrtzKT8qFGOK5HXLZDN1+LqqgAYRoQerbKdYN+m
eIIcWxdGB6OP822nswjcQ0Bsje3vVRu7+Wg3lrUcwE7tU9TnPLL+6WHmxII+Mx6R
1SpXD3+t0J2JbG7VEubXozqvmdH/W5dS4ZLgoa2qJlHsW1JQttkbacDfDoBllL0/
Ptf6YBS+eWCGWvkpZxs+HPwi+TSGS1qtwp8woRPaflFOA0Epod6th54h7ESj8WKi
VRKWv6DKIXp5Xi8xyZ0NA/ya3qoz62V2bz+zzvHakeFYD+wJxZuVPHajVZXgBMRT
1o5zPliZnhJuxqv6+umWgqXvNSi/Zn8TJkEAeilAO5ZfwKl3hAfrF4sF1xPecqNJ
MG+8ED2ouvmm3mM3RLp2acsFv2ldzOl0YEnOPqsdZxBpPtn2JyQhh/9Uk244Z4JR
5qc23bOuaslt83Jhb/kWIdNVeAG7+Ib2534dWrLEGqRHjELTBE/mOISva6jIH7qG
lXAaB6xB7gdr6iAiSRVcPS2nRH3z9U2QdbYQrw+4EyzbFmxTo/Aogs75NyyyAUk1
fb9Y61d98SSUiNSeSmW9Ig4nvBdez3HBTXKU0TAsc9QyUgcz1zYt58EbCMV9TucH
JDjBTsKlc2XTFvFuW3nQ8SNcbNrs8GrX+r/j/EWg9cMIDv5GBTrF/k8rNnxLjl9d
s5SEFSDUd6MzN/IylNOEY8rQ5g8fLAGAh0UKLDUeFx9AcOsxyNTOeqkMPP1FEd2z
0vPka0dvHMJNRTvytcYvwgIG6zEdv7Kf+r07kMMCNePg2zMQ7t9B2cIbFtD39ZvT
4eLCKkNw+xoyL3Lzct5NkiPgEle8OUt/VJmeNkJuwFIRNlhx+JPvW7C0Y/n8I1M7
JQ3EkSNR2IrQd06AdFGIwod4eBiECuRnv1unVvnt+kDe0mw5dWmPigHYrJ5FdRfK
zaOJH99rKGTIp6oMrSYNx4EfmALNCnWPhqCnWCvesSLylJh5ziOdePfZPeElnWXy
vE8aoXInt4c5aY4qlAixzCL7EJDdTneOnGQ5ENE1jMQA6bU3X0FVUTQCqC8ga7oC
F0KBFDClg8r63TyPvZW6SrlsQvPpYPILnGKiNXsDY3w2sGTDmYXQidIhmoYC0LfB
IoPQQGENpjM+Db8KEfGH/SA6ydRPKN0oNYh87DV8ed3Jx30ZvDEA2AU8FySfBS0t
JAe2wI64Bgji26ysy4lIQwIfhzpOmTR2bDQIlflA2KViK85oztWXc2TAFab78YBP
ECYT8JTtcoBJdUMXcF01JQKkovK5MyZ9Pv0FN0HNECH7LavPuxwvOzpo7w6lggvr
tUtBYqTt8D7tvTgjhw0G8+PKX08aW1xyuaDpvVN0Hq/84DNL58fLWRrgz5hzK76D
Yq01oJCBrO/rucynp9nWAwkWOH2N6JbSWEzj78+WQXyOyq+HoiJa8SiQ+TN6/G2t
GA+2p3vk17KYwbnGWtblSysC4c7GLPKTVeTB9qcxveUylFjcu147sOetkk/iUiDR
QGk2ZeloNo7DUvHkLufnObuioMETEj6taB5a1EiiwHwsEi/jTSdOueFeasRizPFT
zFZujSmsojfzG8cBEpkHUKVj1gckn3yFJLrMkmV+hBTkCIg4qYhx0KgsPV/cNoWB
RlnqZRkVjeup5FhVHYyY6dGMrmH/I1XjX0zXOhiNPQ2isxf7eXSRFllUNiRorcnI
05eWiJDlqNMWZDytbV1sJ1KNHvPA6EuLVXqCHPkUoag21nyrMhIvuq6XkUPMtinr
ogmrQyrJtrUxelNEnTtWC9qR6/PfmroagGg7enb85QYH7sVzDhQPdTyif1fWvJUr
Maer6ofpAwiFDsiCF28o+A==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VWlVio+6q9rpzRCBV0mM66Yqq9K0wyBG4huC2Q0IP/VvO3HSJtHod7wXkTNPbJve
D/e+HI1kmDl13lW+yZ/oCqfbEqM1pMTv1+bViQQL3zcX6iImZYU9aXqpepsdwJBv
L1rLh5PkzYMeOgPwiOP4a3vTSQo4IHG02oMlqQCk3EJQdk7AGamvf1EnCm8jbN+9
LWdzoHL9HqK8so5GbU9I2HYT9DOBkJWgEj++LAOxLsp9040ydsSroFsek+zNFWc5
w9zKtYOGCaqh9nh8RLQwfW7vBYOZ8TG/ibxkeZ9XAISGEJP2SYCNGNwurOBSgTuY
C71YeM92ehBJxy3WVVf9fw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9840 )
`pragma protect data_block
uKCegpyd2jM/MDaAyvt2UpMVxvLkN9ze4LNU/SaD10SfRMZ/RKre2pa9N1HOLnxr
f9ITyHtBHOPH7Jl4klUp+BXyWMg8AmTvdDCS6Dlbathvh3R8RY+gI7YHDkUXHllB
e2L8kOTKIhnkihkmZ5PehOnJPwuHI5Nz2KgotnhQdTAS+J3C9MUVb9HgwbJKxuOB
34iWWmbrk7+DbNZ62vw6Y807lO2ImNZLWnA6EGE6jLX6c7kWG5QNcTbIVduaruA9
Z61qVCNtxPy38MP/5w3SHWBGZia8LkGW+oFTW8Ei4sdQ+Qxiy4StOAF89S1PCVzP
pUotMBumMna2v6e+pmCQNvSJhWIU/GIAww3gXzJz4pKmH1o93vLeVu3YBCJ9qPUT
7iDG82hye1xnFDWUG9mfyclekBH0+yw2eyqFO4hd1pohI6is4y0FQJSJypo4uMkN
Q7ZuY75566TPiD2WS4PPsZTyqQgPafhtX0RGhWW00/b5xYJ0sgIHXWePArlgDPUV
GGJnTiICbZdHATiibMXPAlnHuH/gYkPxNIyijkitl2g/zejiG7cekc2uCArEl22p
BGdyP44jE9cleyh2NkoUP9HbUxXp/QRQ2FIbAfTHTGRcx0KIh6sd3bhO6M+oxF1b
Ev7Pru955dA8lT9AewTW+znL+9jurEPkFisnMntUcrk4Ad5t9XgKyTy/UcG/U3ov
eQoNFpPLxVTOnEJCRG41tz9EO9q0yZEPLDQ9KvvTVkBQBdsKAfuRU56EvaGWudTE
REfZqnX1XkpAjQgYk/pPMBiDOaBT5FC+5KA3R+u/JAJEyCZAruYX+VxwIKgiXWEd
gDyOEJF8pEhJHJezJLqI7UHhMbZf0x7BB1h+IYJ6JRbNaxQB7kxslbxYp7QMYW/q
i64Tkd4yM38DSBEHJW45iqyMvIDigT5XTMl8xNnBb5tteYrWsmSY6O8ddPyFzHJg
kQjGVXGI6ZqMTDqst3xJy9r1qHjycYSvNKT236bwX6/JhPnHYrdiRs8uVXYbNUt7
O5EmNf9mdgQVx7a7r88Wstprct8HHjC1y81FiYqiuh2K10pgL37JyID9R4BywUab
U/F5g0ysDMXFX8iXOqqLAzytw+4/AyCTaGlTYfkVmrJwwze8xE9o8iqAlonlcfmi
Ltv/f2RhzA5BfmqlynFON5/LfRo1GR44yzfDvsNjB9i1sQrQOVrMNd9JlVzmOBhi
Rh2woVL2JqYx0IgLKbyLEYt/I/Fw1Ij6nlJRoJ6t+ptWV+8x1haAr/zSlwPqn8X0
B9TxCc1sr7uUXd8SeLL0omsAexIJR4ePXO848cvnQBKEsO4wDAmjwtPzNbAiSdjh
WCiTw0ffVQQHTILArhtFTKWb8KC2bUGQG6w8FWB3VGYQAFP7zngCsGnjAb+tZUgh
8B3QHxiuBzqFAsQ9w0EarFkcueJFDChr/o4FLtz0Zklx1dvk2omnwBjQRa0bW3ao
gYQeDbVv9vJQ+ROWXTeHTfvOOYPSiD6jUT0jnmMfb0JlsXU6RokgVkw07YdzR2IF
HB8AEdlUKNnuVxDAK3P/z+l4JHE226JvUs7Nl5lxCH3THxtWHBlLglL7reMFrrJd
eznwn0e4/+f6gRes8w3AH1xIInbN4cjYVCS+i8UAnmld2vDhb3qhg/p3S7vlXfa9
XKeYZIBf1LkcgLVBNdnG2qfjHaj72T+iRUCE6wzpcX6YamhgSX58M37rUDyyDYLh
QPWbsxm/UvTyZ+/5K9caimEQCLxd6pYSzPGoUgKBnVQpm+rqzkwWXSsis86n2Pxo
rZvGg4pPPtuY/tqX+bb7G5/bekrWplOonuGN90lAmSJADsMC83wptex4kVR9ifL8
0+rWqWkBPA9LQ7YINoqHLMvTfFur2Q6rKfir7VL2UTM2XbuM1X8E3YgIAe+wKKqT
4NgxthcfZkxf1eFnB1bdd2XiZ2onPfHa0LzA78YNV54mo1f8UyeWMP/BViXuZh+8
72qmYRDmqKLNdhNbm07kv8WSDNqZuL9YXroIzRRY476pfYTQQNm61xe7Zr06s9Uj
7oLmOkIFNQOxLOXqsHzkjSMKbd/kAxQz/JCOsR3Y/SRq2d6To4Uv16Wl5fdxnCBE
B5qw/PbYRL8E4C0yBYUfH6j1Rx1t/dZ9JnXgUEbLftsPXlbJUwPWHkPRaagZiBgQ
z+aFh+/32wxA1DrT/WPaJrxZ+J2idS+gn3gS+lrYElIw8LTpivzVSMy87+ySq+SH
NAsHW0dSlpuCotAEszCpBMEPhfXhym+nKu1NmH8v8001vaLowjfk/2E2kTv8sJ2M
sRBCkBzCYVQ7ARU5IesJsfXjOkxYvUHDrY8M8GL7OEv4VDxlzefvpNQKraKxoxty
lxNfSERKJhyP3STNa4Q1rf4/BJvThi1gH9d4YuUekFrwAuhsvTRJDFhYhF73MGrA
a4/6MPzp85L4wixUsC94PCBJBU+yIkQLYuhm1qPvO4DbXRlpGYIagYKf8FJMbg6+
eukK76pYgq8GgJA/G1RUT9oO+/HuUV9/r2Uyk+o6H9Fq3CsmL/t73b+4NBETP7GP
cpkpbU69p3OJDvvITcEDwbH5O7ZI+3uOa3ieTRFT/QqrXNMZ8rcMEBpjADwYQRt1
sBSSPZoMCZfBj0QUt9EM2nSCAkmUWKd02TwZkEod9c91Be6WVpr+GZLAL/PoQ8B5
Ij1VJpkNUYJjGxPwPqmAQZvi81UGtnbJozSe/oPYkRKPaX1yuezUHIc4ngJHLWKb
mlRxtLyc7z8O6UpGY8KJkSGd4CoRgWPBA5UvKxnduawso8O8bn3eQblNXSTMK6wX
tPy5OwVHMtLpSSBuaySRyAcW+YGD4JkwsrXBpqq2KLZkD9FvF2ntiM7SeBzFsfQw
3zcHD9Pow3EsVUxaNiRza4CH4Mq3I3oMKFLEfp2SV5ZeSLIYuY3vXSv5OWCSlldn
H6dkN5uxJlW8ZHhVYl/Y3IoUNsRpui3YpvvGtZW7OXyAqkIO9HLEca4tRO6tvl8i
P1jBWpUY4Ulu3hd//5JYKhGVcG4OpR6pRW96mfCjkv8sEzbX6No/cxpTHMZgKeBX
tP+iTA+cXqfY4Q1I2pk2/3sj3cAb8PBLUjNlBpTZ0l9tkbOKqjSPareHscsWfDbk
4Yg47bzCaCIyEk1ac3X0eNtB6hOKNDEJlyIZ1QnI+ZW+pk/4JscZFR8/oU9U+2PT
3P6cVNabPZKlzFLUEc/brF0KXr05TxcgWC/RTKSzCEIPfatwQqiG3cRCaULWlESt
Nh22CypUhdx0ilQrNCg1SGPB2JDDiqcopVTWXU+MdAU7iEe5N6laFlf2Xl5QKa8S
6niHKF55g3LlhTgXZyRJJcbI2ldm+AxW8d3SMjSD9925FCkF5YYw2mDlbmdDfRxN
CC/ceM5v4VLz7y4hhgt7pyOP9N7VUQHfgFlyWB0Xto2Qu+iAjAcLhpkFgcbQfvND
Haau51IVabTy6QOGMDy2f2v49BM6bIQ3kxkGcaWVbRumxjFRIV+C++Wwi1opK11n
EK7SCK8TpvOqA94unnMqoieCfi4lAYa+5vc9X0M2E9SIRxmQ+64g/lnahuFVbBEp
owYpM1asRzNdXwd9eKz6rZmIMQybrnE55kEaAAmAoS1pgYZEQkizXjARdZ/fHo8V
3TaGrjrevnGSVQOqgWWUaA3fhfytV1kEVCadUjNv0CTLy9kiGirtQ/P0NlB9mvz4
Pav3Yjg9Mq8wDcmPdIdyrG4JT6VMxfTHtTxe9MxUg1jj3oKVZKTfsleCr4Fa40jO
gyAcR3euWUcA/yNr91AdLT6bJFdjKhlCeCwhvuIlTbQeR1d+MZBmoJHGzd4zXknH
CmO7pVXwkRzaA0HiU3s/gGH0yG3h/YtJzCSAbAAwuFcZdhaFupEVFGtiYZBaqErP
vf2ymu+y2cDkRtDTc+PvzS5NHCRNYp9+Oqi6xFoHnyIZZwFPiqjVq5zRzi3BgH11
R7SsHvGMYiPeTTeHIF9Mu8vDj7s5PB17VYBeVLRATGASkAlKcvkN51jBAl28WLuG
+eWk8DyoK44yJcWM+4UUGvUgjBluJYRoZq/QHVZKFGTBj5gK00woFlfn6Xkr6gUG
AB+dwtyxhMdp7Czsh2+1dp+Ly7ZtvSiaBFZFrzsgle4TLY53ieZ9YsbIlYq4rSnR
LdQNs63nqsq94rBFWHWNjKMXteytNvJTrz5wWdtyU1yMy42XaKe8Mh0NMdR1+LSu
pw9sXujvJzeZVTLro2m3JSv6zkB/Cv1Psx45e4hQmkuRjQBXkjwJPlSkwf+tE6M2
gZ1dyhQCHrMupsvYo5pCfo4SLRakXYSUx5bxk2KtgxBb4btMPgbR3tDhccjb9gii
p4Kfy0fBIGZaseFphAXUI/Xry+El82ZHJ8ZsNdJ8T831NYAaXiXwCW9eRUo2UhRa
l/0Sk72vpUSDMdOhtSx11Sp3mbwPLCidk7SgsKCYUSyOsfWyeDIMp/R+vQ7+4XTB
UNrYdanWEE2Fl5vF7rbTv0E4bLwBwkofeOPgy7yScj2DwoGxSq4rpI3yJ8BhkrIU
fW8cPDXgjzTRrjsn3WkuGryXDhNkIwJ+psiHcRxWUPf+ckYX7YXEJIrk57oodd/n
oUuWZEBXnLmLuOnB48X+BBMxeOPBlXwEudEc54Py5V9zxAekRnXglzPRQy6rsEh/
ffqAl916uBcLV619+D7KPAmbA3wHBClKJvnif+UXObcj7qNTAnlk+oGzkFaV8rTr
pLZfST7jUd/KQ/IIGcMMPwFrf19AhIbcxNWYHP8TMiwWl0jtOzIVSpPvYZHIQzRG
4H7tMuFV9V2Z+JcXYeCIZ+5Hz0M5huFrAANr/yJ6OiBHT86fGzHO5Q2DNOo3iHdZ
I/YL9e2wWhaScFk2dccxxsBVHMrIeqUQOn9NYqT5ElGqj5cEWmMwVf2NOQXX2prW
3AG3tqMXlyD2GsqS3L0TRrspYR+TS++cWrXm+hGCHhAgpz0hqjj2KTLbeuTl/n7I
17SAAT4gjWzNtOwWk8/9pDI4rGXq04Q4ySGxoPtc4n+Fhn08rClRQ+mVorITPmoa
y0zSvBYVxgQB9J4s2haoH2g+JZwtzVq6yxghwGkWN/3NhpAw5Ub3WhqhVUgN1Ub8
lMGBNa//xt/UyvrgdvcM7LhB3NLxVaxosqk9/RJws4t4ts3EKSNPqfkdOe2QNQD7
n7PA8+p5c455z3SY6hEk3JykV7veZnSbMOvOlPZ+8/BjyXwEfM2n74XaHjt/bGXq
oe+cQzxPBmoeQ5TyvUpvLuIsaFqSCG0RbIMOxZoYt1YU93qjSd9p73tpwmSU0Nt1
+So3EYXpwDFOXk19+MulTSsmt6rc/+selJ1c92v6rVaqw5tfvnBZwZOPJjP2aOwL
QXqySykcZZhjMLLzSoLtiUy5fY0tTAqNnlDXEMxr5a3/TeWc/7AFsyLIL2zjegY0
1g1GTn2fi8QQMUcYe0q3jerQgS1XPfULpPeJQ6AFYVfWvFRWHvEoq2jj18/qD98Z
RWlihAgqTL72wsOwHZRlaH1DP1W6RkCOnVnpehLD9QO8BtlxQBSImzpqPD7hEsP6
I1zD+S81bVOhPOJMGcvjMuL56e6GtzOPeFF9sKIR1q1L71OSD/8hbbONiGUhY7Bk
vlhlhGDXETvk9ikkADIkUVx+9HO6EGHk7R+SkB/ent1T9v2BDW3XgGCv93u8Hatd
URAx9UBz53fbnOOzhpzzhMRpDJZBEoMVUv+Z9GnjgFCA4dH/AuGEK+CDmr8pjZE9
XAgd5g/i6HCQ2XcZT2RbmP/JtpoWHxGPVHw7NoKhXjfkqkBHO6jH+1DNsuGXcAQB
T3kgOiDogAimW9ya1lkvnAK9VhIz/ZkZs80iYkP44tDQXkVXci6Wg8hUaaNG3Fjz
DYF3dxnZfcmEUJwGfNUR42td/p40v865OXhx6ZasDjoOm48KiocNKlGpx91DrzQL
Cl0cB9TZCBzXz6maJ50eq4TfsZ4/tEQeb1pD+pYvVH5NX2JDLrkr4FZ66P8/TOP+
fXrZiOeRBPGWVvCF0YZyP0PC+9YJjn9QEN82gLYrMbcXDCBVy6RpjIYeU67s8mbY
xblRk4cFNuB1+8lWtS3ISmJ1p4LMuMEnpAOunMn5PqPFwPQCQGrKehJSvVNNDEVD
08tXVVU2wXcmyU6ZIQxKB68Hk5raZf/q4xrGrZYV55Z1c5sAq+awpPkAn1niVahx
CC4MctN6/GVciAS9mnwn3e9VkJcUllM9dqizRsNbZh0JxjcB4WJBA7AfD1W/STV0
pcvChgPuIkSqdbweqNwhbeJJmjCyc7SfJQ6ciQKexzF1nE+Oz9ZhlFshmT3feHg3
T4pKnF7a2SVlH1h9T4G0sBP+1lOx4b+VobxdN0/R2K+mmeVtp6pEW1v6h4Crv5td
2781n7vgAj4YAxfHLz91GbmsGEODYAMxsO1NhC4pbGe0b8m7yIUrkllDYDmpUOhQ
AiXuUic1kT/abpkjt8NpiiNtXcErwXPU7mCs5HdWhgMs48Y/NDbSx6H8mDP1nLh5
jv2Nka5cUqp91Ehr+CP/BkvLzY+twuIYCF7ULKOLbFSVm8xuyOU65CGxdlxJ2jUY
1K1PCa4DgZAAtSHJsjdS29kNt8lls3NBd5diZf2XEgSoaGbrRiJ/eGOxhf/nfcyu
J+SDw27cjr1l9dyyeby4axlFbVyHhvoib51/R0uM508mOwPfO/6k33//uV5Vm9Vw
eJTEOR3rXkPleyoQmz7TyZlpK6oLUP6IAeF964bh8ez5fQG9KRjZA5HvWoG77dAS
m1/WUhPf/2+jSrnjGQZrhwP462M/MEAuFu3u//vRsN1EYBnxQ9SeQ8IGUvG6xYIY
gyz7GBP4txrI2G8nPewEy0moDPpgUMOvjbvgDAd8xrTDRyIAbvFpqc6A0CkngZnP
TXTK4+30KiYVGUooqaa3U7MxVil82IwCclshITgQ6fN27TFKmsFPjURymV2qcIyL
nhPvTnA4t8cEl/JisXRCJrUV0bsDjiIjzR580F6iLh/LQkX+U80ji1HOV13nHDA5
6j0VPdHOtNOK1SH9gktjlmdF/ZPxNj5+25L6xmnoVzIXr1oy/to5xRHofg76iVHl
g+0mIwCO+cY8q3taTlM9VnedNZcInj9FQMjz0ClHbts7BLWGsdz//rn+s21HD9h9
04nk9ZF+h/+egh1VVOTAwAJlOkWCSovsYG1JjAgAfAt/C94vN1YLymsG/Bi1f5LZ
Tx2Kzs7q5LvQdEMSNDc3J5L9yFSr7NkaDdZjz+PXRQa/8hu2Hcp4Dk3E+RYtxZet
B4SaenxFF8xvmqC+JdDJcSoD/z51PrRM59206UI4W2uBbBmdZFHKPDuedzKlWwyC
RS93PsdM8gzw9z0c94gl+YoKv5Q6Kk9qpHz5ytQeiSmhFyMk+ucbVfo6w1Rq1+Wv
dIiI+2tKAE+zXmFpotcivER/CDptFnEafh1nyvOKY5Nt2cbrnAfi+RvvDGF3SlML
+P7ndGVyFc3B79i9UthV7UWW5Zy1xdU7mX4td8NcucJeI3AgbxQwN5ePGOM2Fisc
fSfxrmjx9fZwQ4nmMGs2H/hVdQfXdb50UlZIdVUu/zr/w71FTu88Y/NrfTLnulq/
jmGqvdkG9smSUbtLTzSUz4azZoeA62ljcFL6rI0kdmcK7AA8QbkZHE4VS1IdJTav
SEIE2JvOx+uqzGkHvZkpklAh411qxvV1yxQDUeqrsFh4TieEhNpzmLutWR6hctiL
anh9N0lPPgCdY4LMnrRE20V89/DeMmLR7Ep7TwZ+1BMnFutQSzT2AcobP72szgYH
9HVQdQ78tp+J1YaiUjF36RZeKzx7AjUtdYLGsC2V9EaiUO+TJ8OOCZ/VFtwh5Gi9
HqOaik68upcR90xb9SiOKhMgSrLe4oNVbex1e9TmjYm0HUvyukYTN6EWmRdQuxcr
J6yoksshcHw1Xb+A/aNeUiZfyLsTuje4Z4OJR6HA4Al/06q7Cx9HYExsMUwA9hy9
BgaSsKO4X8bJe7PzuWeTg1Zopm0lkgzJAyz/2+mliB7JtMJTfGWONWaGtQr8aeoy
6+VP1bX4smlaXgOReQVGbzTE6QiPKdb8Cz5GgIMJ9Z34xHPVC5KzNmrWGkU6+pT4
IL5w+19fMYuQqE2SnC8kQYkZLoDjofnteUTuyHDy4wkqCiN+rytFO9PhBvXvD40l
bo9t4ZArV55yLl7hF48KDohCZVm8v7SMORmMVZ1fVM6XZpYzdX22bwWwdg2gX1ay
OVMZdELYZSEdt9U8SGTgBqqiSz6vXLqAWXeA9UTfijoZuMcNQBtcjGrkCv0DpXcv
z86WviPLwoLYEzJ+D8l9pnE2W3ddwfTF+2Yn7FjFeFWc5xda9YqR82bD8XMauuN4
5W9PDfcc3+xV25w91fACX3Kgcq3jLmEyOYlonCu8gpbv6qJz9AeQwqt+Jfj2sUuf
Z855AtGXjwn2gz+X6VKjy1cSdYs9Z7QQ817wRKBjErjM+fNveqzCPnAU0mI0GtZv
dAMyL9NNOWCHJq96o/l78RK/2TOMsoz5ufbN4xlri1Z6ph35vPoLzBFzgbMYTJ72
VRxobh6Ebq5IGozjnu2we22w1fFDHdy9iqrG5ZC2cn9HMkRCopog0JJntIz0SyMA
CtvBd2LDawxrhaRUCtHrZ4zXqdpF3IOGQrLyZrIlYCtxRisDVdeoDjQa9Oo7BIvu
8wjjrgT1xvTGV9NrdAhTDtjAm0EsNv+XQ0lQtZ1aAuizpXkmgBZb6pX2XC+t7yte
iEKcogCGOIj8fCENvy+4l8Ry6QH8dMS3kL7CqFUpj3DOxFwqC6yzZ0279cF2vxPA
utGXykYueG8qsUrY81E5omjWfYLE1OWL7Tcal5tN9LaYmEpW6jiK0CfayFNcJyfl
DyXFWmTS28XLbPUF0TDg/CqHiXkHjHiFbTyRHU19YRw7DqZfZR8XifpesiNo6Alm
ITZpxHEKxcxlYxrMvMm+yr7cGIkopDaMrXCesdXYL5AnThqDCVsZMF935Vaxq7BR
9b3BUuzM6k2o8ZeHGWcemmuVrzYrvXaHzq9eLk6apFzUzzQQcQX0uMCo8Kw6Y1iK
YDhkErOMLbiaGoGEiYev2U/SXms11NMpKKCob4kM74q/w0ydpT4qpSaIxw5lE0J/
1OSOEbmHUZ8mQ4ea8gy+Aahe1Bsop42Cf7TkPq0GwcoEUr0CLVOdKeTThFcKOEA2
4/T1qnwSm/gng21xX3iKnvsi2bW/hVA/I6B/8z6Y0HQtg9+fqRqUsbiu1wJCMEW/
+2dDdaBkSS/I1AFt0LsI1ebguRmekf6bz9nE+f/AqKREe6YBVx2dR012IHnmpnoP
nZ9u8Y8To8SDvjpVyxvSWFvcWmc6fNSFDgLKa6hWXW2l1+ZU6/io3IZD8kR/cvFB
oLUuTJt/dw9y5EyT/DZ7TrY51kiUBDmJWWFhhOYCROQamZCk1E3wKFwv9JQSWD32
A5G/4GjTUzaRizrvFfv5vz1IKGC/QrvpY3V3FLejEShhguP01gTqjWkHhpsTq50b
lWE8xFbDUJkeAyzPf/d9M4L2umsak0bgaDhek0ucpu/rPEdLeU8o535WXpjjy4Ta
//nz/vkpvfg7cyyGJfloO//kVhrSIZ5j6mLN/PxoaPFExzxTu7dXRlb2/v6hnx/c
knsMD2LPFdfFmTaFIgqv8cgGTX4yUq1xTNn/7SSYEtPk2qi90RblJ7v7s2RHE/jo
DmW9E+nF+hcuTI6TWVcmytzdXeDBpy9/4zuftPRflO8W8ab54a4m2pp8LKzckGwC
c2ewgyi6jHZXea4SiqPAKAiADFEkTXsweFUpb/gGz7lxQPAnMvXGUja7NxwGyCeo
JZwPDN+aArcq+pVPTA1nfRtiR9+VSbbuJCAhcpo9RaxIyHXKCTHyX1SEUqI9w3w3
HH1h6ik5KHIvPeQLoJY4YaeqP09fED0iuSorvZuEyB9nc/hlM3cQMTscQWa8i+Qr
OdnpSyiqT5QAA+jgNpnXmHEnbeFB2v1dzrxxpNx/ZBqJb2vot031fzOSa8/7/lvI
PNtlDPU9nfsqVTcAjjI3uRrlVBTB5PxFjXeMkasEvjBLphVzOWgmKm97qXjLqO8W
3FNSXtsQY8lENBGBocePMoJxTvaEa7dbFkAqHhEBvHt/V/2jpaAo2BDCarn9YrFc
dIZ7LxsZFRo9bMow3JjP2xrs7xfGcI8efZkfwnL01o8Zuz9oQLBJuqCyXTrdbg/V
+bhhKrNschjjHP3s7Iqtjj8WaV/b3WpeO1iNuPEx5PE5BPqb425CRK1p1zBkQ4B+
/JnAY+7zf4F65xBRPGqP/702dStyqKLJNg90k3K4mU5vh6Rm1GmHUK7RJtPSXBeN
VRfXsQ5X0N/xOe1a5I7h/FHVcHelNmXyjaWAfe+xpooTEmWPBMR3Dqq1BbU9n+s9
/Ft4PAMvJrZlMtF8PLq4P9EKvwwjvTjpoLowVyUFkWIfFeZdD43JsZGtOPsu3NaC
FDTpCb5W4n6ufMHS8hnzUCdab0XUnzLKrVn7ZN87GQxJciCIgsl2yy9+VxOgIqUu
O2TsJMk6WbCFADTTxNXtv2eVQrKFwHrzQlPAxslQId86eEEvLK2iGsAE6n/iryQq
V47Uqyl3cCiVQmYoJXxNv6sRx3HK9By2zHtwNK0pSorr1fr0bvQkii+p/GERBVX4
0IlmnLSCnAi/UCuBj66l0yOgxpbhj0km5ejNThoTLZVgiTv0TPTmHd02ED8+tRpu
wF+L5JWZ4W3IKFTBzV6cKOe2ZY/9GmDhUbj1oWlfetFUZwIf46pAUmuHmnUg0O8p
DHF0mkishmqWNhr6bwNSh7uKY/8GZsCji95FdJDv742TGNWtpUZwOrXNPJ9Z3+hz
RUADSErYY6BoE3e+DBzOIz0tNZIxRZ/gvU8tqHtJUwPDsljg85LuKAssxHe/C65Y
44ndZjEA/bHraObKu4ocZm+8gjPCMHzNN/rzhiiNkWEH/JHh4v1bHjjaBptLcWmN
WLqXKUGqly6T3Q3eiO+/KXy9z3kSH+3u2qQGsbSVTWFZYwcnb23TtspLfUGoJKzf
6J+b+14kW8+jRytyhD9KbWMmUEtX15TAQJ+ePwXc87q4Vqk2L8o0XirDGGfF1nPT
+eOwEbAZBzLPsrLETyt2PaeAz9Zgv+R4XqQXQfr9vg0Ayoj8bBvsIQchYfK7Sf+O
yFBLGH3yhDQ11Ch8DyMRUzIfXDmuw6z1XavDmzLsuO4A7Sbw7p7sGUUWrwBqIa+D
VtOVIhpSPrTAUV2/wrQwD025BTO+IDTztP3aa9ZxBdKk7EX9gr32vqTjv/iEVh+S
3kegcErQ2nDCRrtrj5M92xWt+aw1B13pifQ9puHxA8WwVLflLDO7diHr3Hy40L14
Jt/fn33jtTuydRlsSPtpmcXFXzMIjnodJtcB7Y/3pZuaXdReODht7ybl9Hg0Flfh
COPoW/q4qYzIZpDmEBaKdboKt5AyZLwF0YtIiGS/uuwWIJxIavQ2NryjkVxO12dl
vIXSsmTedTCOw8OVQRZiyOAdNV9BuagQya3BzjINUJxPB3V7U8wQODVT1fCtsMNH
AlXJk0KxMxhEEBeNCPuw0i7kOJrmsWu6LCrKyJDwIHdHrqV9O8hLBrb9QqVmGIFb
IpKqqE/ek/rfH+yMJXk7DmOiuZK9LPRjQ1isG1Nc4JWQNMqexpB5aHd1m8jbvKKy
u5AQKiP3nOEqlE/0VYzco9vNqNh17z80/U5VrNvDiN2/iWsnCsdnl5AInr96mBrD
LSAqPXF2oReb+deAQJFHJrR6yWFhCUZsY+NrtMXlEyY1n6vFWQ1BBquus/lV8rTA
8u1owiTirKK9RfHjPWwFJLDhVhvoJNusqSqekpuJviA89LeaKH5gDXUrWsih0GCD
/LwkQJujVMGWKH2aCAHgi2tKLMr4jlDk9mWX/FSbq2DRk22sfKWxNy0vuGIg0RO9
MFdSC5KH7Dl2vtZKnZZKqVlrGBuVOlPRNItCIQ88oHJqZma1ett22KnJiD67QNcK
bOKtK/ILjzivj/zATZlanXnVy6hIereXFxVRua0vo0krQoUd1UVBq5htIhLulN2q
k+hFmQ31rKE9J7KAlSGaDxS4nVSgMj6wsauQiTy8VSoZ9CTqIaFpaTiYSuW2wzfy
onzF2hhTV+D7uv64QXbJ6yuGr+LkNVgD6bgs/Vsi4d3NKcg7ZyRmE7x4zSYGKLYS
cvpBKKX00+PbG2rSD8J8xislpTK5uzWMGs7/c9jbKnC5TiIz4IpS8b1yTBJ1mu6f
eER/1tBZVLVnLdb2TmHSUZ0ojXgf/UV4uYBfOjn+OnwaNcTBFeP2pHVkNKZMtxju
4SRXFintXNjigY8Wpyh742g69vZJZ2vFwbBcHb0JTo8MzkGkrYoJBYt0sbZ5XbzJ
LCEzRI8QhPBaT1qEYsSfCiGgAMHJYEixG9XMRIoXaxah80wGhpjoaoiYGgKXidFw
hTa2KvlJNfe5cC9+0PdbTPXY0NnCVFQ0aQsziLNR5hut79cxq6j8nPyClB9lPt/o
g2KZ0hARrnuHpv63TRQtKw/a6vmtrvb42KiMNrI07Jbui6es47Ov3FGQPHD9ZG29
OmJ74r89/FTB9CdKAzl5R58JKYylssB1fcV3rncpb6Fnsv5k5bNI0/0whlmRgZ1G
xAGMEWfvRAIXVadO4iYcErLuE5oCvutDKKyDqswg/1a+iCdkEUYTY3MR5Xta/eXq
y1bpaMSmftlP8ra8m/jvdH4R7X4es0t2WKh0jc1+Rq4bFqzf1xcOQEFpwZHp99BR
9do/iTbEQDA153p0A3QUXJCLUCNrHrEa0yHnpTOkGNmf3hkugyHnPCY4h9DXxXi6
ZgY8VfdSMqrBl6bYlE9hclcrPTZyriSA7aWrboZ+Ty8JwIbncx1R2YLIhRYuYi1K
6Uupfoj3gDCvOAZX5ubwmJ9oiqWN6A44yNln7lqVnXkAcPJFIe/Xzf3S9vennylr
ieXxKDQ9iTAzdnRMORmr/O1TwGsE/l9J2mGQ6fwqaBYQUSwed2YXDNggFfBB6Njk
7Su5Nx2J0zSDVqSPOVbQp+6qYoLq3F3RVURhU1yOZLTh2xl8gg7BkGWgY1hqxjES
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
d5PMWC9vOTaRvpZviei2eWdhViX5DY4Ew8IzRy2P+3A/JVGmf5iCwOVQRthYnFOO
nwXshfNwaRyD1IkDB4NId9vSjnRpfrv+NNa0JSQVJhaNXtZxlYlebBUS5pSLAvM0
DSUOl5U+ti30RFdcUGLFvtNxBQZ/vnsrLbELSfVQEHbZUVgPpe9O8m6nrIbLXfDQ
YZZ9UdN7Xj6XN+YZr1DCtITvwpvUKx1MmLqbUR3OerduRt62W/y7mLHaaPoAg/1E
T2buigu4gViKzAHaTD9eoMZzjrXUpYuPs6VdiMBnjRcqHuoQlslcqtumIplimzwe
IpsbaPxPIETOWQ1SR+aJIw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8608 )
`pragma protect data_block
t2XMh7+HkZREkMTQGbf8+/kZ93RcawX9b+TGZvh9BkfLqLriJTXoTqJxIXC5rXPJ
BjnxBOabtld374G2Ynq/C+yfdwT0xyQfaVROc+XVQa8CO/eYom9wq7Y5X78dHF6N
+6WikoYU7LuGGJTVauvdUcioLCUpZc7st/BBRRotm3L0qluu48JWdyx4OvDHNLdU
qdwIra91Y/VCVF1YZVmiGbCW3lS0aO0P0Lp75RgWfY7TLTxfDoOaHRK/Z3/S1Zfb
YflCkicBMzNMjwatefdDhkxmxfbkDkK0qaNb2FOa/VySLB32d+wDX+uz7gRC9P/T
5JXEyI8k2N0OiIPD0g6yaoe+62T2hIy9TMF7yH+QKz0wE+4aZqZPQ226Qazkicz7
EKon4q1TCxRxJqrGjYkswqSKZHrFyZtAS34N0f5fm4J3SaH/qgS/Bba2YfkgLGun
TwMeHLoK6YQtIXCQLZlYGXVtFBls3CjyYGUKV3u9lTDmrIxsAInkwQ8SaQR8FmWS
fC5WkHZmxV+FZqb7rcAAtH+q5eiVn8i7sN6q3tyUDTBe2Vr7GBTewwYwlUbIx2H3
bPa2EaedRXfRnYTvXYxJFmnzxI7QxqMv+bjZG3rCCZnnDWioNpAMf6KJHM4V3p8O
7OCPHe8W5BSNJt6AHvcmO5PpTZgmlM9XNgnu1VpwjK6qGyMazJeAxmHFUyXows9F
Mobl9K28aPg9IT92egvX55PrTKGIoN56yqyd8IgsetDRcw6o2GEHWsq329WzsGEN
FdOvP7R5BSzYoJNULSc2hCYG81Hz/pMfiyKCqbgwDvvlFyuP+fcXvUEEYeDFVdtE
GkyK/jWyQOlYSkwlOdKpd5Ty1Lowe8T8R8pNfq0SYIe6uA58C4zoBsm87KdOWbSu
YPZDVOE4mbjMeOfogW7LvKcYPWKMCluiglRKyA2TyT+3IEdn8gpl7XjQJi19UBfE
2fCqsyvs5PFTE9AlhQ0yzhFaiTi8/1hU0spZyM5kwQqFR1JL39BnNlZvD2T4zZhD
EOnaRwdpkkLwxZKdt59gmgNJo4ADFmbZUup3WZ6fEJsNd6Qj/6cR1slysw5XPNzQ
kEkuGaHzIB9DGIBM774r4AcusWkV7xFVNnaA1vTTsTeOnMQLGZbcBPJjI1HmmfqD
O1LAiDzY4KBteSsvp05egO5FK06wJvXJJJ7BMu3VFxdZRV3oXZNPvWXto8FJ+IiP
ReRDRppHE6iSrLMBWwqItwW3eG0DvX31Rd8SlMm6YUldLt5++kmaZ6droAQyfy4N
RtB5g/RIx2JMy8GZTlFXUuWlHLqrHkw3E1RdVUOPkL/NCfa7ps75gpIBknioMq3U
V/UwWXjgJmWfky8yg5LsQRhRzPt3W02T+Ou58SsFAp7JerPQqXFc1r19jGxoQuPL
zvIdkC0ecRNDPodu4E+lg4uop2k9GvIztiPTV5foC++Mskf2XTQbQKemvYJkkjjj
jg3mrnE03CDKWKI8rdlfvnHgwdzGhlVtgS4OM1vw6/cGL1y5JB9eKyQ5ZTDAb8YB
VePLKOzhBFFk/I63OjadHW46CXSiyXt2S8pp2V+/UkdsQ1V4wRu5mscvMii4s5A9
ztcHV5x+BojFO5g7c6WMR1ZX1DE1F2mE6boHjs+mjzAhMYB8+gkKnlotzTkfYVdC
l0VzLogqhq1c0wx/NKjIkMUDCtICjY/MV9gBf2gyi7LQL2QKZUiH9l1gEgaZBa5+
trS7/qZzG8tYzTbQBxYqnHGKVTJ+OoglV7zvyqnVu2KZgVXmTNfc3WYXZv4XjQ2a
8oB+f+ATOfHQbUsA4O8DJgPZk+RHQsqOdDaPtcmT+WeM4o11cwGfXk3mucvLcYBY
rX0fptu3Tlj69eeVCAQo/QDwqoTw50BnlK+/pHCSOtYCHGFrZSOPya3jkAGpC/kX
AayTnn4PGB+wMFXlhV9pdfVrpwyEwm5oVx2oBJogR5YifmdJvbiteWjy5m18VoJ+
+VXlVfYEqe6kXWaUtKq8sSlA0NbnTJcDVvEFjM9ZA2fOliYpahVyxVA0ncqRNs32
bAiPQOc4/e/LTcn2El1Iqc4bB9BXaCDAMqUzVDfo+BSNd8IP/9dGWQpycPdvcYjS
bXZVR7w52/STbMesKxPQfwRTvydAggL2vywyAxNQJxfm92R/n9/BjihGnmzYUjzj
SZjr+T7buZOnvPSmX8NpVScRCUlImgPfi+hBpDaQv4pzk4iBYrUtYbD9TnMk1cR5
h3NLd2fhGqlbDj4NjfXWI5tdqx6kFehIYsh8B+5ic/bUQLE71YvRZgeLa2E1lkh7
4n4FmNZEh88CuVm3zad7Dt9rouRywyEnN4fg2eAIjQOe5uD0swwlX4wkvy1fKPLr
17d40Q6soIEHpx35czBrEP+9g5WdkIBAkASsjcrKHxKYy2cUVAiZad0YYgow9vX0
0gjNHkk13f3kWWht592754M9AAW8quA9oxew2RpOcDzX5iFohSporC6ZPL3sLdnN
Gij6gRnjj9SaeWTDWYbBCzEN21wn9llj96s9OmxjYSeVkeKJ6IqVxV2k/AUaLKPU
CjeqqwTMHFj6ghkryaF9FYomPovf1jHEqC+QWS8jsY4/70CB1CuMK7TLGtMxPAkR
4XRtfjH05PzG2kuvlxfO9GD7JPBiv4MgV8M+U8LuK+oFvwXUaBU9S+ZatvVmNvgz
/fSGFMCAqJXgjGPCHVNkW4ia6ILw6FYWhlTSSlCO+lyO+0SzC7OgXKyjmyowu7i6
X1gBCRIVTcvMj2aAhjaj+CHnn8B9SV2tZRYt+1AIRujYAbQL4iRrw3U53jzJkbBl
nhlUihJ/UwBCpqMySdxcS0E6BMexhIOxr1uGRoLlCMYnRelMV7IE6dj+pVRJPCD9
7OBVDyN+rgbZRCjzIFQbApvgrCR4LFYHDntfn/W+jV55ERXMPj0GzI526a/oJy5d
GhU3RIiV/e4oO8cKGJoyJiqn3wqQSXJWJ3lANjXI3X+0il7qEOAdXC9uOHNa3Rec
PleEO2ssMPKuWP0xx1N2QWu4c0xGWuP73fyyn/TRNjLygqPPQA2LmlseXeIsDJuO
6jWaCQ2CnDG52SZC5U5TxehKI3TwEAAwwHB+DIc8q9DaNZfhRZi9yEbP5+oSAutC
xoRvZ8n9Dynck7FHTHOnod0bSmqJfKn8B7RDnRRSZmfC1vkfrtnmYnxCi0UhGKo5
l4lJXPA0SirtQvMKwMBA+efw8dxNQhZcr7DTE6IWd7c1Lz8j2s9eqxokmpYPBiuQ
ltxoSw5RyhtgokrevSKB58WS2dJFDe8xM8iywcG2peCeX00gncOEiEJDRVRSd+A8
wRYcp3gJ1yAVqqLz1lPNAXM0V+77/8nsbxjiH1gs3PiavvCFFx2WtmGufROs80+y
PNXC20CtHBclEQmltvJINUv1Om0PQ0f5/JVX4kvhlyfVQOdBeFSCSdvMILDuCFtM
WgQf/WEk5V+UKCmskzlPYlRiIJa44ReUH1GUG/P5dMsBhpH9BMBwpnzKJbJItXOF
rn+Yq981mErAujoujDG4s1IweXDWa3xqS4dDxdJEFu6/2jZWTN3K2HBuCsWNofV+
GqLNQQ0uXVLgas4jA0TVyn1S2orRxudFQI3waXDcz+LbPZaOLo+dGO8Jpu0P9Aog
iNioWpDHuFFWDaV+Sk/Sh1x+ntTM8RQ7cvLjqn7Ja5E4o0qutv2PaIYzUhHXjdIC
gYrp4IsK5hBCciYb3ySb4Y5TIgYkyW6KTTw6M4TNnvFFhq6+WPvnBifcA0DkcTxX
1PfihOn5aQf8oop1o2TFnfRJNseF19NBYHhbkI8W76CD8XKTF/ed9rtM6PRVK/yj
AHGeZpMr13Ggwy0J7rUwrYrxO7LAfFWgihZLtKXPv3XG0MPTitO4WFSXD4bwel3D
WeH/UtUJZEqvUhD5ujUfgzWL+6IgIj2j0cEJjmPHOHalbHbcIixh5eYUZ2mi2lVL
ym8vTA7VKokjUZroMOwk1wdLJwWzI7JUjBu9Q+ur9TESOKPgTgRtjeMwAn+HgwLc
QGlybzLutn/Tt+3hemDmTEKGzS9UFiBgnLyLAFeOfE2bYfhykcHzoTZ22iu9EoAl
zTMi1xVtnlfUFXxz3FpJlszPs2/p3JvuEIU3Q4WhbvhYyV2wXqnL7aDxAs7o+vwM
e9IR5wewoyTFOcNiP405T11MJ05eTC26UkHIMfB4i4/tgNQ4ZPcLoefVpOI0MB6V
HIFghN/0dfY/rtN+BvU4mO/DKr0HhFvS/OjaCy68FwkGH+7RB/ZcJiSh2iYdEsvJ
2ALWUwkQN08X/dMpF9f057JKSIJL08ogiVm9s/ovKGbKZPXPWjtpOvMTihuYdK+q
Dt7mqB5kQPTPGn4ex9E8iptPBDX3Bi6Od96JLACxd6H+ebHC/qtvGCLdntZNzCsR
6ugqA6fGrYF2f7ASYuukGgRqY1qHPLqkta4LItTarLntGmCI3LDvjG0eFFsUzA+r
FDT4q2KuFFcdVP8r6UewkXzTWep7yjLg93KRhdbXRjBd50sjeOtlGURHJmaRIlz6
Cl4b93YmTLeFmD29Lft9KvFJv5qV8YQL1pnwvSPYwzUW4jGccIiMtAKOCMv07uOt
8lMWRtjwRufU5ABgveIAKTM1Y+Hg/ZhniuSgLbrD0Qebd9Y73RQuh93fqHz0qP8a
TXBnwJVkKYtAbXJ16sM3HxO9sitl6bnmTSzTjgmk/adVWj1U2rYR22fXW0b60mny
nb96qk8SUJsklKJOlNASaYFAYNFkNUxO9z7UuLixD/cSpvzmH0XYlm/L/0qQ67Kv
0m4UTqXnnNZWE/KUL80Be4Zva41bieLoE8bfqkP4w/8i56mAdwOsvbHaP3u2khw/
nEdgH9nhpnXExTGN2c5heQi8h/LPEQkNyJ7a/VoJGDEeqaUFgqDYrNoF4ulQ3OoP
CJqjzgvI6KF123nmqfaSShnSRBLlK05V8u1U2dHO0s9jIushQfL+zju7PJylfqE+
a6MOVll0aqV91zUfFn7qTT2ozCxsWDOudlWoDTaBDVWxLjW76Cxox8uPbF/J9bhb
zq6LIBVZ5cF0LZmyN76AQ6ec1UhyvPSuyLD4Hix5MLnlYse66CDh0buXNaYZUixX
MpDQamRY29NxpQy4cI8/nRVT88j6Z5878uChjURaFfadkoGHuMKQAMAsZmnGkWdy
g53bSDnSaKIYSk1myzqHqbpnoy0ZqzlzY+t8e5iO34aQdbLSCkzAGpmC1DF8RnlC
JQ0jly6UV7KaryNto39dG9kHEGVUJV9Du86xRBHgNl3nS6wIze3+Eqa/2lWdj/O7
8TWeuHtnrA9oqIG5JzOurO9ZWzEcEOUr+e3bhft06dcpksuWv1qfAisU4l3v/+/q
geHdjLz+Bf0x9PdIEux44XLLE/citDwcGz2Qmq6onVO4rAYYzjvoTbAX3IrN1D/g
a//VQNuDLoMXN2Y2sZz0qoSWyT0+aU7sF0zRB2ufKKJY3eXsAkKhjBNnkIeeKCCo
0CsSHMtShJsi7zN9XLJjfT1a9edjYHmUVmsh8hmXrdRcuyf6I37lPyoN/dx8MMTm
JU/LbVUHvs8aQ93i5R6XMyX0P7iT0cCy4msMa/2wdEgfy3+4ApM1+gGbX7YzFrXC
69xBtR9kYRg8lJTyD5zCMBAIVQj3ZY8o+JGzxdhdH/s562PVag7NryLwB0nrDzx1
2cdCZscXaKlyY0xNxzZntDB8i+IsfUi2vNqoUM85sE7Ll6IwtyMXATy1wR51B09u
mcwJpqo/h+WhEesQdQXxOr7cutJhMN7R6BKYu8cGqMoPqxMclvnPCd8CDj3o0FYk
P4t2nz8ILklB6vQFgsBLvPSb+kgDjampUf9xIrgPqNd0SlQ9efQJrYPmMiYaq/D6
rEVtNd9CWUA/f6iTfw8Yjo/0hvk3M18oIvQKU3/RaccW8MOhe55mP8WDyFFZIT1j
4ZFtZvT2JAqL2Wr5/aXidi35aqIPS3KMRfBhZa/2i3RpqEvJljmgKThoDfGBrak4
Q5MIM5JX7xmBVkvqA83eK38kaxiIdfrLzUdme0hTQ0xFWRBt4bRIJA45z1dN2KkI
YAX/JTn9H4COMrQRooL3yu6Nrlt7ewDW3KEGcgcYMzgl8c0diphOi5bRa7iWnCBq
3/43KjSRkIE3ON08dEamL1+0fCcE7caXW91JcsW9pYZz/Z104cXhju+xwFiufAXB
FVwiGVx07250EYbIE4FR+w/DKUgFuV6gJHDq+QLATAhxzTau5gWUI+HjUnpypzJ6
Qr4MSETtsAsceATUuPt/9mWBKSXnUww/ZEO6S51KkQjvgoNSlVIU21wIKRqNiXcI
agRKk/4jS5IegZniOBJ9mfyTOec2iSCXRUDb1LnAeInMDnrsyAYJe5J0M021VpJX
gvOZlV/jnC4Z7ijV7BDJnLuErXelXIexlgQ0/dpCMj2rPsrW2ym3qqpVg1bk3F4T
QdjvONZvHczlQ1ZVg2pNOqxBYSm7/o3e+M/ZBWya+W98jXlUccLG5WKAbVb2s9km
L/Oavazs6hgctvNzkROGSfo9yP8YSEaS6elh2TjiELPNAK87ivQipvlmcEUE0OB/
66oyrWMY8dd1UDra9SBFN+qHcsNuvvq4YV/bOZQQk7fWepNDg4tcf5yFztPRHmWZ
tGmA63JimTyNca+Sr+BZMBOHumMtrr7FMEzmlmP8J9YHqJWpf9HexEJd/f/RgGM1
8sHY13NoL1GzP5HsC3QTneNZUZWa+GwHqPWjIcMS+5EAv8wbHNSo3zH2KrsXUx37
4b7J+ZOmiNHiC+Nd3wif17/7hWFrbrpGMsIq17f/ACDKaafdL2435aRsKAN6L0jr
qmT5WyNuqQTO01lhj7NbOBqvHDkdBFRorDDqFdtO2l2OvkwRD/KhDtXA9J6ScT3x
dFnQS0buloA53CjdFQeXqwicaGiY73zV1B2uj6hZyf6Q8XYFfc1z31hmD5tN1UPx
yT1kakNEVUNCYNMZG8LnAMVGUWLLlH3fDP9zOsOMvwDEB37Sj0q7hCDdLG9GK3ZN
FkUEraBUK/rQpqWQBpx7LsNAIBtsrHj2Pua6eL511w9/Gxo3c+U7aXsD793pLSX7
k2S5QM2x4Rn1z1++W8xUNkm2/tFTX6A7+LWosgn5oa0vvtKe5MejH7+jTfqoT/YV
0iNFPw6Jdmesool77V5dyyS6FiPjEARHtYtRi2H4HkjXYH2wnTTiwYgLdBGIUZPe
3m1E1Ue5h9xd0REV0VCNtNQVjgjl6IDOC8Jg/mTeOKgtuzVpwAV0ZuWCQHGoN/BL
GuHc+vUtCND1BmBdi95Rrz73ETMKXJv6A3k043RIDQnPsJzqnVGgA867vEDW5KNC
D9m4DlPVs4qgknmBcMM0lPcpmggPOj5gR/aq9ZM9/G9NHwtTsmpRkGgKrlqGQaoC
24WRzXIKYpionSnV93zMJiQiCm3YBxJQfzkdPuI1Uv1vbuYo69BYFnodyAWwXpAk
ou2xvFJFEVOZgR6d0qZsRMuOa69QGn/Is/n6Y3xUmDsX0jDzbf+ekUHjhPgQSyme
pz7RMH4VxhXt1EIwgsdToKAR8Kd5cs8h2SQU7eM29LFJTV1iUPTHqPZR1JXHpYPG
uXUjQRyqbtAxs2BjE19wMTsNAIxWCRub8RriwjfgfAHKxW6oy/27Zd94Qnulu1vF
l4pOdOmtpkHD+YU/6owCKK/TK/TluzGDjoe4NYNXGn5U9WeD8n6jHOb8RUw6Yc5J
h162NbRC2o6EOIhX0kNY1TlN158qTfRn/jaSkeIOfl3ykQure5s92O3XAgBr8+V1
PKgNB9KMXoObZ9oV9Gk8Ci2Lm/DgLbaIecotkTsczIlM5uDqwk7mxTH3aYK1Lj7C
Xq6WSEelTViT5Wu+9+4L/PrM6wfvouvE8j5yHa+0jUD3XS1yjOK56DlzohJAv5/z
2G6BrXQNNrmb1jfaNIiGmOHmgTtSmUN4GM74Iva3GN2s7DON/kJGoeS3g38xZtG0
BtWhTEcYjiNAM1xTTLCG5v85wG9UmQVwlmSR37J3tS3l8C91WQLDhthDTq3u2Z58
AG622ayUWyxPJUEPgxo16z+ABZt/I64cnbdmZwRpKisttdt8vIrkEUtHMUMm9p0e
AtJsKKETQvCjtzhiLYKu0S++XFC/F8YlQHsM4bh0twWWcP6MdvIt43C8tzoMeRg9
S/R02BPFrAvzDTiyZntO5OeIMm1QEyd8OanTeMZTqJk5VRHZ4AVCyMfQ/6JZvBMx
40dehRokT/j2pO5rnzzlsjU+cUwgwdE9wVkN+Liv6vyU5qkg4MAoEKADaiGgWUCG
oLL1oU1uW/IlQIcaTHI8cZyE4t+8w+vrbnkWzjqbQ5hMfZlzz13plc/NZddwdWJ4
R6xLVz6paOQ0XdO22iAxVcNPA37pmLJPBmAul9ydgslGQed4czuWgrhLKQOd1NLh
1WOdw3/8yKv5vPcavre4+htg3K9rB0e95qLZWKzirDzKcKUg2bjdWuvbNxWhmeNg
gnj55QflnHk63ey+PV5bsfi9o1gMW88VH6bkKiezmuCuIV/0C+9510ovA5zSQyTO
yJRK3XsQDFIMcey4VQ2IZPn9rH0JqSM2WKErjEebIMuaGNyH3bNfta2QhIGECYtp
UUaqU3JjSZMuJ2Pl2Eaa/oFOJ0OJoRm9m5/pi6+q/lfXok+R7XQe+b1YLBfeARXw
iWRhzpSfIJ8HNDK5Shq3ockr2J+NCuUWaOqICQTQTtPy6sLdfSFng9xKVxkvmWCO
jsUpfKhKrCXLs02JZWARPBlf+dte9uNo5w7WxQ6Yy4Sx7/rXOfRHUYoEtX1ey1HA
QOLCzvadrASaoAIweOX6LWcxVmgQVmjEUa+in4w+YU73T1NOA4/K1Z4HXZR7UB0I
vtzjTehfEhDlelzL5IBzxNqf92cw/jp4gNvr672eW7OfwJCOWn9DENNCMrIGl3g6
+tNIiZUkLn8pEyw2dStR+oFBAU6RcfK45YMA+sbncWzql3pSe10KR7q2JP658w2s
zkd+LZMwUySsVF6h/co8CuZ1ca2oZy3RfbsCQ25Umeb6zgrqiySjUDU7caZdN63o
OHmNTNG+DuQj65Cf2N3KhbZRtZdKML/mKIb6cR9oT5OVPqLRK+pdRsV8NcuyBdEP
cy4H+yBx07K3s/pwZN7NoN/gnmy6DjYtWqAdumrGITEG9mztW5o7YcvC/8kIxr8V
8287NHEv+ILF3PxJUI3BFkYRidTR38EoztCVb2NeP4UcVXUfo/x2uh5t79KOoxse
/emcyaVvPwgLU6d2nJJrZSJP2Jqgv8bcLvX4oplRXKnskLUkIkRuKxFpvYisCXFR
NoseFo1IZQLT9OTdH5WIRWkYgcLfCHmjqPadN+IuJCV3FjsHroDaRxIeJGU9BBSD
cjm+eAIyFh5sElBOr8CdXaLcV9oAMeooj1Sh3J5d7600pqnJZTIzlNeD8voY6OTB
ls1BpBWzeuO6ZfYvAqZs9aGOGuTiZl8MTOt8IWdIwuHinEdg3TVNr8JG9zQN+1+u
PwEWTMudV24u15IlO2d8VTJPN/8re1HJERfSjZ7IE6HC7zILlnte/ENa0yE4vBRe
aGYhoi/JDhfesfMelaOFSeXazrZmiBDodxUvJP0XqFIV76jjXnAv8yKheTBikSE9
/MNELoiZTKXg4fyJ8mRkfOdXUempCPjKSFrGxl/bg00GHy+FXlb47VxbQjHxFz9F
RpYT0XK5t9Z6xeR/7goDt1PXwsp2vXdEW3LfTWOwnRbTw8NbzHUuwGgxzwT7FAhd
mCaYnHYuC//kDwE5UIskUjPbnXmRWl1isFTj/+e9wcMtvpGTd8kGpR6Uh8AGYE+I
KSfRM1W3KBRbwugbh2ileBmOGm8r+61ml8Cn47xP8E3CPsAN2FXCFeYo6Sr2yiNp
emnYUw+wNrlRbhmGeAUmU0q+Z23mU6K9F9Yaf++H58/Ne6VA5vbfgYOXd9IyQEp9
O0CYMJa970hJG9g2dYo3ZHFkWWcVuLiU5N/gh1gBxSe5NmkzMkBgpnz+xAhdUihi
//d1ME862gxZNoTGEmgVrRnFHNHMHlWXC//nTzNutTsr0oBn2KcEJNykAwuNwkV7
Z/KovYoJ0XGRfaE98zKA0k1rQkoNfmTI027H4DqrRXOkCy5Iq17RwyEVRUqfHG8r
PtlvEufVPd9/KtP6kTpA55splNP5VSYZ1rhj6rWwulwWVEzxiI87QGSZKXwHvPNt
g64T51d1Mk7SJfuxwxmRCYNWzihp3g6PYIbcN9loahAISkeUR+9U6YGr6aLgWTJ4
M53EpYIBQ3e0OdgE6UdtWYumVGGtR3dKz877Gs6qRb2+YLmwelJt+tNAReZ84vpb
DS2uOBZJDJSL9AtbxKKo0WS6d4uKqn/2yh2UDnD20D2qVQI81hP135GFZo+YpH8S
bGjw3AnjNM74AijJRX/qkIM5Wgr9svlsGAb5gOL0AM6ugidpE9VdbARjlr1yqk8z
FPYLmqPL6thbS1a38cPctHwLoPgM9lbFSY/MQ48liZwCegNiafCOlc60SPexWuvV
kn4gda7byMTP5OncopaNsBR0qXuLzVPoZDMOZNJ7JkVNlftsX+Odld0xwCpe2y8u
6NeIZ+YvfTdm1cLk8pjU1WQAukwy8OcFcvaT4vbgSK8g9dr9fNtDGI/a/gPb/65d
Xh9Lq9jbE3KmBripuoR7Ubb7sD7qKGIlHz+mrZ4DLqclZ2EczgzuwSwS/p4weprQ
trJhvrfqggVTEzaZWuDsR8lNysFxGG5qxHqeLUAVx2z7QvATZ7BeSza4bQV0qjxg
cNEeaWCLtSVRQ4hMvgfyg4HiKVmfTkov359Fy7XA8JEv+fdR+qoHuuPzQ3Lhl4bp
Nh8m9n49xXwNIY5Fe3R1zlPV2DwxJMKhQR/jY90I+n1sxuWO0Whe/M7YBJkXmT2r
WVofw5SCzTN5aD0BzDqH7ak20lrKxtPY6E1OJk2HF2ouQ4o43aAYiGONHMYoSJHt
QqougjNDx7Wo6oSTe5sT/g/jEhpTGOkwIsexuENSLbzcWyjoJdICw1LUfLh8AxIs
2jdE/GnRO1DyVddAu7Vjq79nEp/S4riN91Enl8UBP+vO9sPvdDu8QCFUeRNbDLUw
DK0tV5hlkUXyCpssdZ6KYFiQDAiM80kJDvf3wqbxbOkc62egzZhYhGbUYlBR8S3F
wvA4FBcHji22TVtde37dGLL8prikETexXATitjBG8+bhfzAzX6yywQH1VyXL1+B/
IgapoPjxYyzn+nlZuNcPGOKXBIjC9BYEh4FY9ZCkJR0mn9IjP2qXhFGsKoq3/4Ee
asftu3hf4JomBgoFGizOwXt7vquetYRBfeiavIRbjzhsCMY3S27t63tI48PEL3T6
k7b72+CxmxNp7qcxEC6Y5Nf61O8NzzqCOaPcyGwCe2NdnkEUwNW4B58qdumDWKk1
IubbU1ilClrLxd88Kfvk+Q==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
c0IQrTzgreTGFNCAnZj1/wXehwJjHk7Rh3kNIzT5eoenS54P1kItUAP6Q16kHNWf
xzlKSljqSxmcjn4/Ui/SMHghNHpo30ex1q3PNMZBpbRWCim1oGDw0AIdVBAT0d0j
1qstenObcmlp35he4bVuTo0wChfoj6GLWepaA7qKLc9E0AHbualN0Nt6znrPa8YM
A9CS5hhWd0ouLC2AAHfpgOsY5O3nCrTgFIcR3yD/79MBiH6MeubJmuHaGnLznHTH
Z5da1tybQLfvLAEpLEVsA1ONSsRPuZsH+FVNNMqkpcMUjGKXLkTYWynLcq5gcXh9
ldh3sMD7epUPHuqXqDZfPQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 29120 )
`pragma protect data_block
95SXCBR/GCOJltp4pUqZQhuZqo6qLaZq1OTSeN7UN/aHTxp/qC7gprsVjKMEkNnp
PCJDOIT4RU6zuSdtUyAC+UrrijMTNNe/Xh4tavK6P3h8tv/A6bzwnsLu+oIksc4K
Kd+9Mka/lvK0nRd0eXkhCIMsbZ2+/KFK+8rR3kjvLfgLAW5uYLnQ/vE2bHKz4u5R
au1J6QpJHo+3XVk6AtAsbAxth2Buk6MGrf09bK9aA9aliKlyRx+QRMC9NN1/irx3
LMVCofy1F9ypDxUCONi4ULhQkVYKgPjio+T9EchZgkgAWBxMLRJUCB2LKXKH8Qi0
eZa2ls0b3mmj7aJgguJv0FVzuQ58OKUCD8LjeDq8T5cUd5Kma9ioaE0aSJbt392g
q1ENNCL1dcUG06vARQszaZr1vVDhDMZf2uC43rmOqWRV3mvuOxTxpTILqGCM/WTf
Cp5xItsAXAyZKbrp1zq+L083B1YZO3+pddjeb5Ny82pyZy04QI0/A5/kNng/9Toc
D294cw9zSOjM/ZETle0UR9mAduqo4SgBoU8eMrYxbCJvHjoZADf30j//VXRQOrhW
Rac9Hbldd7FH+8OzOY6ekXdyQd5G7bNklwpbF1Yf/itJYp/Euw3X4alWWrGFUVlC
DFS4ax0nqXb1YA2QnvQOJBBBpzBbq9HWFyJH69+PNA4byu9rFGmSl3KzWD+CLfgd
3zUYDs1a3QlTWVOO5h2deFhsbykih3ugQlQaz/kDfjnnPv5fXAhmKwbdtVpFMF8I
CzSvDfQJ8vScnhZwQlnyiUVXw8wvIPC09peb1ae67MAuF1dIMKD1jj3wq760lw7u
q8lRNzxYpOz7477aC/ThK/OMSP7PauWIsDMKIYEEtQ2bdLvB+/MzuaC7Cq5pdC1m
rWx7TRZpBFAPP0szZOL05QfI6isV1feDFuo1YIjZM3KYPHpcztKM3yFLeGUOpJgu
tASSd6idkT5V2TlMDUdT0QfIBV93Mp0NBz1rRzsgWipXZegfE5Lw0dt0whbHmCn2
RxnG3uFHEV9reAPhb0WoyipyYozH8XJ3Hx41vNMnMknuOLiZ73p+GKj97cDlkmyC
c1aq0s7Y46vuUuzVPVUgBCfM8dGJLVWnR64syR3rE3APRcMv/xoVjwRQjU49ffte
WImHn9lORrwXjqqJhS5Fbd6wzpKYTqcV+qvqm/X75LGDl/lHv3KgjqbPzbC6y6BM
Z5KiRujjO20n+bY49kjaL9XlxCZfqvF7AOxVCEginHCHjR2DuJaGGI89yYa/z46o
A8uER/NQk516C/YCHh+q+XvGVNK10dm0bT3tMQMg9kexjHcLyZiV/8AvV22Gh/JH
ujp9j1F4IecZlSNNXOzl0G5QxFCm6ZYmvo8ENP8Ybd8AO3OJf+G6oNwwPVJd6CVf
t2jvCylh+DBEHfmzHGLbhT6DhGbJkoflwNdHQyACacX5fVlLNkES0iMauZnIl/OE
fbU/QHTIyW4ZtBhenL76tojThHDVxlMvXCI6uVfQ0oVYJAga1/TAP0aWQqdI4nGL
w5I1b/p36JcwrEf4W7dskER3XsPYt8eFmzP47mxvj11XiJwyAHNjLFYrWP63oV9y
lz6TMBPXpTL0quB+nTbVwSIAd3tMFB/yBpHnWArxROBmyIKvilMzJRh7Cv7NIwX4
O6XMY4J1VFMT069V7PZWArOztX4xf8Cehp9ukeGLViyUOa40vrUJDaJbdVPeUfAv
keeT4DGnqYX3T2p+Rseduq0Gm3gNjTMTH0u8UHnKQ6YbaTaIvTr8swifGOpSYm4K
5ly/3r2YU6t4BvZPWaaCykD5Ja87SOK8IXRaRCZKZ/qz6nrShe9Vk0dTzy6VoqH9
qCPLCn6Oz3DUfFCHNMGs65Rexx7gK05dE2ZWJQm8nl9Vjl3M8b87hMpdYwrEnJPa
LgbqAnaEjaWe5csu5jAH8pfwYIGM6YIN73rmMzcZnFS8et0NUGhrkJB8Sbs+e5xd
W6U+qXyGoN4LgN4+Yq3ZKdXzxZNzL5u2602gaquLhwS6rxjgTHk4C1nFesBFmgXE
pq1sQWwncQV+YfIWLCXPW8r5aTfAGNEcrqu0x7NABFY7CbN8YDZ8/3H7HmrkTUIv
M9Y7dcZL5xpzrl/JAZvCP013ZlJw7y3gq4gEeAnuygE596CkuDlru6comFd8y2Rg
qdkV5SPjjJTSu1UTH65QjZpK404mcdGYMfU0qMUNDzf9z0wfqKs87ZKrZibBCBzC
XDFOT0BMt/3ymGoJRO7MqlPEIm99TzoOtcEpnInEzqCbrmrQ0hS7DFCbQDoLcgTd
+qvDrO5EGPsralM1Jh44xMQ8kBvC4ki5U+i+SR9qra3SdJUAgHAqe/EaUzXtjKEb
PzDaXsUwXTenaX0wAIo17cKQsNGwhw/RPCUbFfeTP5g7DrLX/oJ5ATvOy/XzGhvn
4uzvZReSI9vuYfS9njKWENn0+8gZMHPzTIjdBdzZjSKKCiJNEn4DbYMmngPI7xzN
9/ggiT1+Rqgk+/VbQF+CdBEjcOW46/orAJ0iyhmzjE34BySEqHK+tA3qsTDnODV7
ftit0wRaIidtsVWmCxaTpZas3kgiNulhszIHJeTLTzO9JJNmTUHoHqPFpJU4FV/D
70Zn+mwdr1gzZux4nPOuvTnHicklexWkjKO/Bhk2m6RN1c3HBqpi+ku13uUvh4Jx
khVSEBSyl1APNvA+sS0v2OA2eyYaLU551ByMBqLc9gMOMJvtVGxSgcBV9ZEsBu+1
5o782vd2nZHZ4zSvPVKG7uN/bwRNjNpFSVM2UPMgjJcB9n8QDfSRXcPrVzlxE8a3
kSA9YkpZqlHW6gV3BVHRgnRi+um3vhgYyb2MRXa62sgk+DUj4K4RLo/IQe0JtpOe
HBHA5Z9IilQ4TUkHt6uT+Ndqra+PJkzlMQOjYdlCUqb/2ipK5THmT2ux4UsH2BtB
d3ipdAJoCQCsXEmgPd6fzWi6IAf4Y2E6weKEuzcMKaQYfc4TqOtpNV6VZluStU7M
54Zp3iFg8UD9tzLGqK66cHEAtP7rSHVZ8m0RmyavMVbb56o364aRDR8rqk/cmhli
XHyNQvForB+pCkUrK3MJYjYKjpfMfc+5mHSM7aGP0KJriTApwM8MReQSKwwq0tv3
wXxFHJGvKKyofRTm33vGPRtGG6IGzRe/b/pm7o07rHfUrrne+igR/+bTPNvvJLY4
jXnp1BydSRmvfIMNl9a4cpoRfo1r2bzcxMGmyF2ZjXOaly56zab1PcgXwhFn5cfh
IFGRAVDuj/2wE+Q1fRsCnZ0/QPwmF4G/C/QscXO1MnKf6zlpHMFC5MdXvUGOobmq
rrJfejheQ6Cu5UB2ISx4dvZbSYWtL+JRYLIaQrfuzNIoJFfk5uHLxN5/+Hc5i3rb
HehCythcSMd8St0QsjEw8gcgpoF7gR/dcHC7mz6VTWjbOgjxc60KCbqLfndOyFaj
14T5m4KrPdR2tFd9RILmhpK1tdIOcrH9Vx+RkPOy6hiBtiAD2C0dPiQKfXRAyvGP
wei/YN2Wo4fjte+SkbsTW0SIrWDS+C1Y0BozezXoHT+5Jo0SktOSYEnnPFhOWkAL
f778jwWPvDfkMrMVAiGAsE4IPgItR2xUxC018d6Y86ng30/GC2eA/gSOzoMNvzsH
RZntm2UejRaClmZmCUdSYNwTjhH/UKjS9Z0vbO3sZORKaBjgfC7FJlJU3OGNh58g
kVeriKXQlbGZLqPX8j0vIeSl2Okrf9HgnJZg7lKQdj7wQBByutnFLdIyBLVraNM8
EKmN7qKuIruFsePPPWYaBQ2LPtIQj+GQ7fvvjy8g7DcPS8DbeN4qy9llgaohHq+9
PD56M6Bt8LY0cUHihJZ3UsNOsYf1w1emdA5zmVAnGClapKB7bCWP4DwlGCNY6/Ze
hc7eadoyBJ421i2zpsE+CKgs3gL5P+bJQ7P+ql5WFtUytcDvwxsTjgSB0cJJLicm
qOFYdaEUFnCVMy+6Lfhd46D6LS8ZMdo0gNPL+zSeIlU/M9Wm/nlFwtkmZ6Yejl3q
nzlnqjfveSm3bnPgKUlRgCdKfkhZwpDD8XSttKItChpD4jTe2LGBL4z5plCylL9F
BILj1Dd4cAAs96yAgwhFNj3vOuGNoUwp0fW2gJO+uP5wcoMAgtaOll2lmARVoZBC
F2/qxW+wuby5NELs4J2qLZftOMFE0DA+GCaMTiuvpB1lAOyQiDi/nwT9tdBoNJKL
orkGsqoA1tSZOVsWuESvPoVY6ivapB+y8E6oseG5bi6zTg/P4ieIdPcgbJoygDgE
gOFKCVbOiZM8cxQ3ZCaZsaEGyJxChqpNfKHaxAgKsA8yj34FE2IzDCwPm1Ge12IX
uIKIUo1ZFdaJooCFdXoyXPiISoSwQmdCcbgD3X4s1yE5s6jGix/seuhOxrZuyih6
N7TXA56Aw9ZuUaR/SdLAvagA7wyFpzZqfkaAx1Tv9F+yJIll/VKUFQL4U5RAW8Fb
wW+5oMTy/t00p44L6lUwdFGTQBpYM9HAO5zKjErs+NZEP0pmr0Vgkw8bQEAEtbnT
EbikZFTISW+iTky8MCQth5N1BHaaHuo9xZ3Mh56QQzW0Lj+hNVPPnRo174QNvpTv
5G58itJmi6Jeh8iEeFJIsRSxGm25rG4aVvA1vlP6JGTisnm1sjnthTaHDQmLf08L
jrspZJCO6mYZGKuodpn5kJeHXfShQDafW5+rmSSm90u4W8CFY7BKvz5YT3jRhxcQ
/8wCz+eZI97SP1N6HT/PWsHG6nXPuanL7ZI+bbmMig/yA1BhZcY4V6/HgqNvEfFW
DkNvJa9ToVHDc4oawIbLXsQ2oMD0ZI3BTyFbuzwb9093ViFT2JG0ssXAUiqj4VmV
kVERi5p5dN5+nSOLHoCJX6XEDia+nBFTATjKKq2H7YFswKUgoLgUBbAQJ2wEL1dv
9PpTNXqb7VY2LFK8oZfdH7Oh+X/2Q8baFSuJb15ZR/EDssz+FAxlVjYoz7VmAzLz
Cg2vFlu22GhXawgZqf/z1yexKqGnODwnmHgFHtTHulGIw1OMwNeE7s6+LZ7/dBrK
4GYm5YiQjadgkzW2bsDJNZW+4/gtY33j4nlgVf2NQVZ5m4K75fjXMrXpuDXtyT16
FLX+EX7GNpPeiQypRtUnSfz69Aq3vqS04rFBk5bghUtgBMXHA6E6WR62zhR5dGNy
Hk6E2XIabiUHEJGk5vJIoSfqDrbJ1QxhkWZQj6rGrHLyS6T1tE5CRaSr8jylzr9o
mLb8eZBCdroHkKkSMWQ/1CJ78Gc4WqGjzvaSviQXXwJBTITRLrOeZjZkMjWjJdBM
2EXyc8KXy4Bk57ZYkRdn7yOTbPGBfYBsEhdlIjGSQ4+XBeuDCjUgWP3G3eZpiD6f
KaZuSMzUehDZ2BSspTuTv3Mbm9BWiVIP42WvMyyiUYQzt7xl28UBEwQLt/p6tzwg
WUxDjrpOsMwiR4n1kO+RFWLJ+QJGCmrIOBFwiyY2lXVhmwf4gDonXeSWttF3mzw3
AI2si3wvLpNbrUlQHVz7bR+VFZWcZVJgDboKGyQQN3hVC7oiZwrV/r0zbgD8lCFf
mbPbZs9CA82lsa31h94y7ZQmuFNZtDNWvNo99SWR5LJaox/ux5i3YrpaBQxIMh/z
HcOyF9XhEcShQLFNaTni4dIgnRw3Ti9qglaJqtFsJlzVtp6R0BcoEKT/RVjrbDXT
WsSh37wUH8+omV1U73FJVd2cwd/N1TEvvLpdlXAAOkCJ13nWQOikQAU1BQEBghIo
nln0DAkUESd32S6o3LC4ISkR3DXVJA08Ct/OEnBQTeNa2DlC969h5eiUhsswudSb
25HWJVIQcyy3pnNS/5zf/F1uQm2dlsnyFahu/l12XJY938mUbLQUFrsbDeqZwh99
TsdkePvzbnMs3mMY/lxzykL5mEz7QFRV1dCuOdtXPByf1/J99L/T+a5iljIF9tLf
+SyjqVtksOybXGz9uHhqlfNpM9cJcaFYScauWx5ems2tqvRolt4GyPPPdqDp4crn
GBItcIQmnyK/8Xp0zh9ryo6YUzY/GPUgLIZTfmnklH+n8342bZKQ8uFc2CKTac40
zNR8xPCn/LP2j2vnd3K8R6/lXGRSit4tjPHiwDL6fMHpJzTBJN0vpl0PqsxT4seq
cUz+/ABKr6d+F60+6pS64cIH665SHhj5bqHsQPUTg3a/J9j6Y8BAKJ1Ovls5y7b9
c88N0PwbvMexizCCwFfouu/Vs9VIgyDYLDouHMyEDhvFqzr1jp0OsdLREZh/I1l1
K0lT6QKWmUANqvcVFOxwPPeoq4faDf4kQHsv7Xdzy2qxN59dmo3dIotdTYF3thm1
2khHrZGNbOfmgoJs2ljbf6ZppGoo4YwLdg3eNOm5Eg+oI65s5fJ7IQMhZz0UTS8N
oXpHDzvzEqU/n/1b0lqmZSggxu2CVup0gQI5LsMru3yrMIlHJq5OpKtMm6yLTJ8v
Lu/PxzY/JMR+VqL1ZK+ypWa8AcvX4z4pvgbgYmWxJm1KExxmobvJY0UQRmZL+JwP
c4GI5mrW80hX9kqULERJRPqMpf0oW9VHylFqpZMFWNC+rWZt/QL9OX7pQe2Jx7YL
89dqQv7APs9eGKTxFaQ99KUcE8Rcc/wmIfA/jCaMnVrM7HraIfcj9RUdwo8nnzHz
LrVZYhw0z5kdT1yWus2uqISGn7X4uOT01iip71kYlNcs6SkxXi469ZnxbblgMosQ
c7nvV2uN0P+hqH91mVJ9XnDtCgxQjqP5Qz6EG4lszdW3rzXbZd5HOTK6NqjUyj0S
PDOOzDay/XNUn2LS3OCiwkyZFL5cg/AKOvLTKTtqeH9+dDOhZpAS/K5MfaX/pMAT
Kf1+Bbroe6/B9CMe2odFthynPu633suTHA9R21Z88TwnKTJQLMPlNpFD5P9ZFVHZ
DAUvsw/u1E5SNNLT7toe2xz0OuPdLSY2bnOayTtRwhws6oT6TX/Z6qyxLILJ8IIq
CgUPAxpDbt6xqUeyleZ/n3No69Y7dkrIybQII1vm58hltv5LXCY7ldy2kLUndn5p
6SHy7vq4fRm1oApJ+/SLKEA61DowbSgFCk3Yc+fW2+34JmDB7CXygRicWaWwKWyT
4pzulJ2/CuC94Omv7IPQy1I/RnSTknZw1vzIo+/wcsuNHmdDzieRsAkld6L1//EB
SC/6BDbPzha+bd625VG53z6RR5pYhJ2RWAQFBoIG90KKOaOq73RsBo4Z5i9rHUIz
1GEuIhRJCDuDlvb9XBxck4FPx5S3TgYiTcsIVwxbOiK0WMLQCU58efNYtDBb/WxK
r+zZB+R6nht7gEaKfXBALPJzHK4w44bl9AL0j43FZI9v1occMdGv8wybs9QJOoqA
k70ULHt2mbngtxUQjMTVWM99hmodaU+F677Vsk3Mfuid5vnDX4Gf06MMIkOlVkTp
d2Dy3GygHzpYMyfuFpGOPB5QUB+CFOuBIpUvY/oGoTIcNp9tFG90tsSskwTNvFvQ
GHSQjFLqnAQjEc7ntO9xD9XlSTZSXQHNCckPnUO5+TCTyg9DiTpGcWz7gyZH+t19
YpRyN/f1ci+2v1ddzHWDkGP3Co35m9u1XOUkXICVFXAlUIL/quug7naMos1QIj59
z07ORT+07xWdFfWUnDmgPBI8GeQm9uVNslt1DgFCjjRAq02EjwfzuQiqEgGBKFZx
vF7/LW+VseDvKH8WGrJvENklshyWH0n+AzynytnpgVnlRVpo16+0tS4rQ2EvIfrx
iGTyEf975yKMMYub2Efk63MTui02n2eYck7GVRy5IfiA6sL5KGfM3CkBnm6Owfwn
0DUFROgiUudmNSe170U1fgBNyv3JWJ3Llpnc3dHU/CmIkD+QNrDfx58VddCNKmp2
2H6NECDq7gKnfsqVapIYR46XGb855qEUI3niV1Apcy9xWK/0DkG6k02STisXyDNp
mi1KCQn9E62GTxwtn6iJn/2a8sgu+zaL7ASsmPrfzsy5zA+aCDAXa4RaVnlh+7hL
Mww0Fm5uvDhE0hw+8qCj1LqxfWA8ZouLIEAeHsZAur+/ce8fgoKNqVNtHwHoqzW1
z0uBZh+PMlFs09rkCeWET32Yc7cX/EFge+xm0cLckbdXn1M0VMncHnvsSq8yoB2n
690hL/Nu88eeUIpPcfYl+csw/xEgKy8X8T+WwyUh6FRgajdVFR/7qayZ15Sv5bJh
99NFrvkg9FMbgTH+YGxL/PxiBAfDD1k5goRVBkSfJyuND1TwCfx3z8Fci7EBQrhg
jTkj2A5ghAwja5AxJ8iMXA69k+C3oPjFdT9a1OY9czwzUt0ybnTBhfQmj7yBF+PD
nYgbCO6mzOmgXQTmdSvxFnBFGMWB8a1rW52ScOIxEeVvNlwdYrC1MaTh5JFtle52
Ry1Kka7XlL6Mm1NmazRpejJVYxxFLHqUwckL5Xrdu9ycGrFpOjy6wKxSAzhhLdN9
YzJf7PF0q8oUK29pIMmwd0cZiWGlFmnXntXH/uJIV3TnZ/FCTc1v8l87YfAUtXgf
wr73c3gJUNoNLamjYWTpoChEB/6vs6t7bJ/ScScMfNMQIT14+vVkg7Xu1RgWfaSD
fuJ76HjoI6ZgHzkgYB7LAn28B28msTai5Go3OHxHFqjBBrdC0MKP+sFxTcyCSHZI
nZjcIlapfLnjLJJNoRdmhOg/DxM82utDevIYJKi8RZCIzRIilkMrb8JXBXI4HBNg
KVRYX5q3TLa0rbc6vXH7pSAzQEknupA8qk3oipU0+T6JELFpvD5qGajSxDHou+as
/Y9YNRjzZ7wei4MAn74TA7Z4Rw8Gh+FKPQbf0NVNE7MSck8qVDpAgi4QPEqQBeFx
Iw+mTmBr0id4PhtGF/qvJFKeTHuYjUkZD7xLo4WCJxFLf+iP4bU/pZf3JD1FLu18
/TZDXdtTiN39/eXA8jMwT2FDtQ8Kmpv2tARBYo6EoBYuz1ZQqSuDNL+p0GdoNwrd
PxKMRO7IOwduCQA3h6YQJzr71ScyL/Lk94EHAlX7/cWXA7H5Zr1yt2MESc5Pd+a8
34EYkklmvAvK4bBnD1UiEavIRyIzXoiHNmzZ3S69XvHpNOu7ciP1yeX2oVgCWR68
zNM9If0t75wQyNMinZx2p061aah6rakiOTFqYEOYlYo4NhUkz16jI/f720cXTLzo
IlchKZXrFNEPw5vfoN2E6RnKQQ3gK0wC82f9bM5vlo4bL7zArXSq4B6+avVkUvi4
qFw6Rn8s6rYU8JXlzlXfe/Iwc/Cye1YIeq7bChfZW1wRXzjZi3froSrNqD9qnMpZ
9n4V5N/GWf/tVrXSTtFTMDCoFcLzhlWNsreqBCpx3Rf9hCnx87zZFrdSvoMATu4H
1WZxdysXfQ2RvOjQb7eJvqYCexBAleFZqcd2hz+XG8YTIXNBJiU9VnMDzeI0fIH+
S31tm7HETOW4c/HkYF8Ao1W2vB81lJXLp83ElYifmjgBU+bbSCq5TMTKeaheclmX
1wms9RLkiQ70Nn4FHF6cup7nAFnMn3p3pSQ9y2qOYPaPbNqqJTFJx1ZrcGp8clNO
1b+94doRmMVwHxQpbX7MRPeB1tHoIiBoAT5Iyb3lF3LNdV8TLA6EO26F6tYbP7Gx
gg8jvLUsF+Xx+PER43TCPqdDgWcwXDz7nSBJAfUDzcsU5Vs2nS1J1A3zmz6YobrK
O0ttlzMO2iP6tlzgMwzPl3Y7Qt/TBMEFp5O2WtctNntNLP/JMApQwQEaL3CqEB3o
LMfjhwLIRvvP2+iN3fs2gO9gLUuyWZ8YMi6VavEKK+clkqWJcIp7dEXxymzgOAjT
IuTkhH7sUbWQu7LDr0stnwhW5o5/9rU5ve+QQKubhpQSnzv4x3U6VyhKJdJez9Ls
ozKN6xxF9uZ7Gaz3ZIH14QhFNkJ08FcZUCTddpml1tVgMD5ABYgrCWowBInuWTAH
gVkfmJEKH+tTmC0FwQanLkPGKwCtDdTo6kgoCCCHS6X9wKce58hKjP92Uqc45WkQ
6SSP/mSk0gdZLPYLBLDv2P/driDvZ8YhbXlAftNO9sxNYWyMkBRrZc2Og5HhJG7t
vL/79jxXav/mR+ylXixIKDxApLTIFQM45gLGlK8qNUsYOWZphSWKQwDPd15mznby
b8Pi/xkbkLAvM9J04GGRDavv2RioNvt36ySoWmVJTA/pULg2IEm8go1PBpHgg/16
pWKRJMnLkheMimgsyHNgm74nyQhl9JprhX+kauDW5PrY98YzOK/MKe14VtgrgPFi
sadlA3030P8PQzOhMHvFSIaCgki7Oiy0ntttaMfjOrZDGLLWWZ0Gh2hnsmhBacab
BQviSQ4iZnMI0ElsKeW/fd4QV+LEGdDhMEKNch/f5NGBQzj5b7En1AR5L4AViM1s
lRG6dMxRTNf48Fwz9BBrns4fQ+D6Ff0XWaC/lL/KUwCZ30Vg7yWKYBThLtWP9TEA
YMmvVLhFCucl9KAZLM5rmvu4t27KJeru81lbJOc17kJC7MpMR8b6ylusq0vY1JzO
zWNnDo3mzdrs1UppUvClAV7qDr4hnthm9yxkIYr67MxaOk+hQLAGaYpb8nbR6xEa
Gmg6RB7fj3BBzN0o+SeFQCEcpG3sMoxeQjlgDqXAUkl4kcCrnuvz3OkTX7YLb9II
CaeDBGVwgkbEm1OrP/o3q3RkEPOi6F993Tb/GutlS3l9pBHf7tD6E6DzfMwS9pWC
0bvpKupm6Vb0K/wh5KyypmS0U2n8d8o4qzKtbx++PiQlbTcxp6CGiNku6Z94Fm6a
2/k9p7vPHkKkoNJVMh4XMKijUaYDMuHlPd495clEuNAaGaDf+PVUfQ8DYBFs5ID4
bZecq9IkxHfNvLXlboKfKUv+VU0rV20NIeUsbozvtszrczQEkkBc/rB3P0DASJ0E
lK/Lok84h0uPS8XMoPwfNqnhq/RU6u4sqdbIwov2faKPxtbu94K1lRkuaZqtob6Y
fw5MEsY2sm73IPFLGkTBQWldc7YibjykoqLKmK4LbaoSNQVm1QjUSAtnpusnbKtX
aXUm0ausZmrY1L644JFQzLwGw9aRo3Y6XWRT624k4J2JoNaSQg6XwfI5edspHPZe
irYSs8jM51bpISebOwD98OQPs4fdEy3BwM8UoKt3G05EgDM0e7WYATqx9iQqrsay
WWt+vbnAbzqdL/eZWzAayZIgWwNO6bKmsOhBEb0M8ujcmkpgPcSPPlOjkxJ9EpRf
6ymmrQmWN1BqPIHjcplXTYLTfUdL8XDh7D2iKUMb/7apYpTOPiPZ3bJyWKk2TX+a
9TUMtVazoowq4KAxstpJVtf9E1M0uHrkPQx0aObG5ZOxB/Vyv+8aLnrErAw+4BAN
cNPPJni7R/v53KGUBujYrQ6jGvz7N298EfbkU6L0zVksneDng4wwh+zEu2AocdDd
4SB6wsgRUohGmgDo9BwzkvWe4HglIjSChkNBlnD8s012homKlCRpTQGqsW02iULv
slOjEAVxTGGlTl4ocw95l7btTsluMMv8Jk7jALu8sPYrbDonWMNBNERazfofkFBC
8MXuNIbIbuoJr6lPLkPj154//1jTO8+LTAyZ/6SZmS3IG0tkODUYJ5f3Ks42YTtl
f3IQWCZlPyMq/fQ5b4rwGwaspqZBwWyl7nJdi1IX3DDNvNRA+NZmW9eNUwCDZlx6
RMNeeMaS8gUm0el1PUWj2etewCJsVcrCLM4K/zuR2bJi+vGUQPvkWi89mHG9r5hf
T1y7bYFoVnrf5uGJxaMJwrrnL8Y2kY8XSsKJIt1DiYeH6VXEo8IRjIptCDC0429Z
dHEganQUIQdZmrXFfgpWG2ymdGwlYJzWxdPtFuk46zYeny1nJHn6o00Hsu6qDB8u
ckkBF8OiOsZqlssqZsShh8wP8jbmvF4TxUqrIFXAHtuHZfmOxYllgfcsG7tgSdrs
c+EHC3H53rzHCjhz1SVd6xtS69DRxTaGZkzsDYUqMJ0hwhXlaSto3dGcYpULBDpD
By7CRjyZX2p7EgmRzXAz910UvBdKYZh0xJKWU0rReFKAfKcxbKH7UCVxR6B2Dc9K
2q2EUMVhDXEqV92rMwV6ibSMI/GXG21iqTOD1coJKtztj+XuY3rqGGUYAzT+Set4
3K/KWHkqISQpWZ38/Jcf7AOM+x9h6L9rZcGL/FCWlW6pW7OxyRCD9W89Zt8CPrWh
EROHvZHQqWZtqcOgDoFVEWQ+WcZP9BIMs63MAEdnMOtOjG/qc+/rhyTOPlShBxwN
RDokeC3YkK6mMoqW+wbvSPJVsxY/NEBaEEvFjCbfvrATR4pCcHPjf0NX/M6HuBbx
/l04ocA5suw/m3nqsKrNkyQ/lzGJ/YGoDxCNEVQA/01wZvI2qmpA16K1GU6Ug2OZ
YqdDIb3gAplSX5Q5MZzrOlsO4QXckx2bjk6Bd1t1DkfFppcBCRD8uxkB5iACbr/f
Zb1oBUkAKLXrzHE7UKKCcu3a/qBooxkD8utfj3dDd03nPkLJuHi3Nxlau4WtW5uJ
UYYOkNtuRUQ2XaNo7BrJFfLrCDjDlSJdmZewslxhBDS8vL/CwIbvV/I7Zoy6Qj+j
Kyhh4Abe6jgrvUbXai34UWcuA+loO6Z1SV8MByOcykzP6YC5ghSgdz9WNkkg8z2I
d25PZARItGszpSuwLPYXyOWY/JInqQ2Bb1NY9B6B6s+6ngz/7S2CVgabL1UIwo1M
2Z3SVR9VgZF4WgyfINvWOP31VoUs/AvaY9WEmkUG4ghtfk2nGPTcgNfFixW3iEAR
ztT/zs35N/ljFBrBR7U+6Sxt73hxfJhDlZgVQP78NCDfPXcRVUPyRQl0RFcZnyk5
Q5l+zOQ/7wPuVCeArZp2a15h9/Qk+hEA+I4j2IQiE/NwxDLDHG895XPSNT+zX9Ha
G6V3qS0WBngODquB7y9Y+58wMOa7Kw5zDxyaZiKdVjWmlTqUJbaCyDaB2yB053kP
5gLJuXW0QsNOKJyp3GjvDZo7uAxFaQCv8KPFJwFahQIT9++drHPLrvloqdFZ+K3h
r87sCbChH3Ar5xNv1rUfj5V5uU67KtPJchaABPYk//x5WN6SlTRyKn7cwq6dD6mc
DjjsbLMDTBJDLA/Qi+Ut7JU//T+BDoxSAknGDtiJAk2KRipAfy8FTGAkSmCssF8p
pI80OWmvel2/VqyVr973d5gaHqjuvmpc35ylCT3BUUXv0pj4Jl1moJnws1XgL3wP
s1OP+DNeF7oYf9tJWYe70ZkK+GQQgOCIIOd0vpsJt+WBBh0qYE5/KSZDF885Qjqq
Hcgu2HmQbhXy/umia/l0cScfjK4TrQY6kSccLLhUqnfIVTETzndJDB8pZdkQ4pxJ
64Bpn868LkWKv/afW6+pGUY2hPZGB32tCntRXe+WcgYeLXP7oGmp0v7rR5eZ4E4C
Ls/icp/caTt8S0Fg5M4wWEHVlS7FHNdPejS0vgedTAlRJi5tB76nkEps+iV082vf
1cAg9M0XeRjkFxcsmcikpq84xSbHcqNP9pdBMjEdRIjZkBwM+epZthiOqRysVZYO
65r4DsjbJNygMNZV94mOGkPlCgpWFG/pWAu318TE6hpmu6Yzd9Y5At5bk+6u7Q5v
j9AUbr3M7P8fbGXabMUbO3n2NJbuW1OQiwn4Nzp3mYd88KHVRnY606vMbwWILicR
sxxcwPV3bEjQHrZOTqw5wKLSxmmo8SL+WhVMfN6JlxtyEG8Fb4geXuleLSMTIZos
/BrQbfoWBrOF32lIBO7FyomtludHN9tQ6s05nasnCSU/cc+l3KS6P9Okq0ttqnSl
b/PKcCXR3uELd89mQPTpx3epmMn2gBIomClG+/RbQeH3M6JZPkWORtU3WqD/tBZG
hZb5+w3GnUcvB1gur8V7FC7PnB2qE7/uWHWkxSfQVNtVcCdraarvTRjhPlV2JRoe
OfICeRst9nquJTX6E3wJlzQ7KpLdNl3YDIMApA89CupuofySjsfhcbk8SS6DW024
HQGLZPHPbDvAhNcqmtpnMhuh/gjOXVaGXgjeun6qayqxDOo5Z++pJhJSAoqUb2I+
rzsTH5ygSWzL3L+3kzAFLRKOkWQRDM4gVCtoW7IPh0kjboQBECy7zWUNd3WsUcec
zCsO7mLyWSzgYjJZQSns0nJUj3puJ7UaSpmtKB8+BGtS1ABMWi5kpFurU0mofTZJ
kifQLuaTFndftjyU3B/InwM9WqGyDGc34j+iHNVDNnswYU0oHFGct2JRma/gUa5f
sXR+dXctAjSeNHFyQGr4hQzLpg4UyZTpNiW9LgwS4nxpfvluE/Hjm1Qy7+LYfo8a
7MT4BMBKO0D7zWDsN1iWl65T/PgBRJ5ecxp3vxEgOmTuIZsIs1mAy+htYtzVcvtc
+zh0kjahKa6GUWAUIcOG7dMMVttlMaqIKqhS6kE+nz6va7coqhd+SMm+rYHiXITR
NYVRBr7SlFL8ozogqKnmeZ2utWDKQ8WWh43aUX/q1YOZQjw3Nv6vgXCk2A3hZTkD
WlOzfglfneybVxZ0fxy2BIfawc3TznW1qKYqeD/SSGzG5k53x7+09v0B/mRfoHov
L/8NMIvvT4kS3j7RYrhtv/PxiASb9lSMlPDvmR6iV2zoTW9Mpg7QKDlv/wrE/+Di
8Q4o2TbKxvoZLKbxyYJwtnbfZVQpGyFa3PoiPPlq62ED9UesTpAfkNQeWa13Abpz
AwG19r6A9qt0rWlLJmVK7aDKp2ppVhmerMYY6wh5u5VF1lZDp44GcI5jRKBcWxie
FfFFpbv2WTi+PLAdg0SKmsmnUTZPtDea9T4b470zgZ7pNAOccpzOOYIfnKTy8R9g
q6qE9yCjzkD2Sh60TJvI2vmhTgcLYPUup0ZZFEtEAqKNfgsZL2VOir/mIhO4SLuZ
O0GgBHsbnrfhXc4bUboZBziMAx3aW7+ZCbIzDRfzBIrIjFQbsl8ywrVZzK8YqWrx
6ofgFgdp5yDT9TKnDcYVCOx+cI7tw6HIPp2EP5aX627tZIP8yix5ac9yK1juH3p4
Ay1pH4tik5M8gNLduThgMjZyMYppJatK8/mwbeJo427+IEQcSmGYkWr8XYP2UKhu
h6CVl3pXDLXfJM2ii6wIWDaQmX6GUJ7mO4oS8B1kLJ+pxVz7NJV4P5Xxp2eYaVNB
B/Fc7Pg+1I+vtVp/HT4MwzgsFa+Np22P+5pdt6NQagjZ5vo2ymFTzqTj/xauRnb7
p3DlZXYQyRXO5sz3UWINrw9R/i7rSj3B88wQXEYZssvde6GarVFOqaPrhgISUJP9
aQPcp9GC5ADmvT+8bZetQTvD6H6BfKyjMhZj0R5oTNjLn1gFe7JCAdQ37nDvh25F
V2Vk9ssRwBSf5joDc+ub6ZHQ7RZ1HA0Evwda3lI4BoPCsdTMKBGT66Rwnlhm4s/k
DL2CH84fL+PEfPdWEmKmOFjEpmB3EL2Fpbq6Bv+BD41qT6aufkRLmozdEmIVkXuo
wmVF0BVLWfWYXIyvz4Q3q4gqOFC2/KuZtRIE6Aqc8HJ0FK8do5bISOJjljWeUgDZ
I0NMgYCODzlPiAjF7aKGA8favIW/BqJ8XtsbcZ5x+4/YiV4qth7mUJnQvRqbuzxn
uRoNABvyU2SKxh4vc6H6HmGGMfQlStU9fAzbenKL9OYVBiVT3uqOX4uR4b1P3Vl6
K70uVgmM6JXgAcbHixanQQCB7AUAQaoCTqY7jCo5ilcozKn7a2oBFTJhGSbos65v
TGEp9T+NP+hImqOqYpoR5SqfiEiNhEshw7600WpDKpiePBoU0egL0uAETJA+9heN
BIn/sztborIuKlco+ieQq7ec4SAb6HyzzuAhT+q/D/deDEZbKophK1r4fDyr21eU
GcU/OiSTNo9f8EdFX+ih9fiVvOddTZy+O/5ZsSEb8osW7laRidENJGP3vYCmJTqh
3Wt13r29/iPh7QIJDQuCkxqSo0YE/Cz59JZYGdDD1+AxQE4fgcK/+k3fw+wDwy2B
5SwqIcoTKOvea19U1OMtJ11j9LKhNwMzJLt/+9sY4e1iCNfM90jo354BMkiskDMk
GscW/po721adzgDze2wvDUM5KH+r3fCuw6PwL7PRprZZJfM0J8ruG7grddZr5uUq
3qwqw1APe9fdm8ZMvA0+gS+pol1QOmmvSGLDPUT3o1gy0/qDQ8B91lJCEkGfifwG
z9bF1bg4UFCU0fNlwBQ/9lFEKHkfTKgrnuvPEcdMx5ZcGs8Tt2qtdrV4BCcoXzi5
rdwTsQCcrhq2qO+9TW7z6jU743Rg/3KMKeRWR1QtPtT28nLTYYyLnTRPGwc7t7b1
tKPcVVJz9X3KibjWad+iUBnZi6J/PrjtyXOAnGm2HX7DqTBln/Wsqc2RaeNIa+By
TaIZP8Yp4jzmIKTwhBmR4V87bWctKogqwNamXTfSYGsMLGSLxR6dMMrm8GLRhH0k
oAVRnnRKsP4EZc8ecuHtyVDbNUFk36CCKw1LtVxAklR4CJCiQ6UkEUUx77ZsgsbR
EaHoM9AvvcwZ6oqMdN+wYK2jr+TGYwIegTeyCisJfsv1D47tlRlyr1T8P1c+e6QN
vIViA/O6z3DlMz7P16owoYbFBS7TqdtJyu8mdUuZle2p9mywInIJ/CY1gAtmnKeK
wONtub2sLNafopJ/Uda2gG2YI1GrG3w8ZUAJnKzAA0qO9bemXYdyeEeEjFCXZpge
AH2sQpc/J5FY3odEGnGBt5xlMRuu2kKp946PRV1KL2q/TuaGjhVU+oE7U0VD7vj9
NjCECuG80Ig7D0kcNw/gVLVi525P6JRseoFrTBN0Sdh+tT4dbIfc9gqwD9l6N1r1
L6TD7j53CReLgPuw/U9u2QZGaISWmtmuTZMu63gBbO5RqQGBTMLSzIQtEB42o/eQ
JiEwBUW9t/pXR/JKqWjpi83rGkieZIfH9JcG0jlHOf62B3t+fDAexxAazoyeEOy8
HaIImZKIN1J4lgKT8OmyZn08Jj+ANHTkkKze6Ijs4spNNWUHO+NM8st2BzIoB9XO
o26vsC2pu9PGWQ35D3y2PY/IrNOn9sqnM+F1gVOyZzfHTj1+CMnHBfnW5L0o/O3o
QWvypxdyVKrXykuI0WWYG5gcrkuWb9lO98v9KdwQl8EHGK+Fi+Tfo5V47tBqkjry
796qDn0QUdKafDHIZIi4Gq9yQGQXuZX1f4O2iGJRU+Y9FLwIng1thULLuo2Z+5Qm
HWJARaO5JLzBacFCEmSX4wYtt2tYAuytrarJdgPCYqLNO1a04YFkIeZfvCVdd2bJ
eiAF+4r/PBfVkAsM+KGUKOz126xng45vi+jhuYT/dx7eXJ87evGPSUix20FfvTtE
x0L8rc5WOhE6/Ay96m+v6YAV06vPGfDc6PPNKDJFZbKHH37Tsu3BsDEMsloRN3pp
Pj0oxxbYKkQIpSiSyfqrKWXrlP+fBE67/2H1QB3pKwBP9+9wfQFBcmk78+3cAHg6
wtdM5KhbfzxJAl3kI9ESH27YZAMkqRLI2fYF84P3VL8SSaOTtMutKIE8HsOLljq5
OlQ7QacUYdZiGxqFG6R9XbzwhCU0LpEAKXb57ekFrC9SyjiPl+QQdj5LNJ5VTQ5H
c3PsISYwGHzsMSYhnanckvcupfpgzitzyJ0/IlGU0gGd1j8Jg4CprYP197AydeVY
IGAp5TVoAKDtAnBmtynLfhDrcXFD1uwCrIQyQvoaeG4cLLNImlN3BMb0n5A2A09l
fyaaH/3O80EpYzzQMz02Ow+u4ZeXyXc67P2HuPMmbuvS+TEKkYAszP1ptO5nkOHF
pGNMK1bPHuxZzDJxDp+v12D8dExxyK55A3zYkmZqkWFMcjDckiv3KUziDq78VLCc
6DHEAZOjkuAA2mG0fNwILvBCnBUVrxF9EIfAGHc/lq2KrGi9V3UYqwPGRsPP6r4X
jEVCEFytL+UVLFdtCDI789BuEMovplGBh1x/2d7AUQ61yK5kzu2puQeuiMwHHumJ
LwfzFtISidVgKxPsRnQiqZQBdXdAw4sCFyeJHRNPB141scmmESiE5u0U1Nl65bCI
iHwTYBc7t04t1LnapMDhvoVYNWhmaF8M6PDhvcDGFXRhuJ2GfdBaZ9S5K9HmseKG
aGKohSHx1jN7ZKYxpbaUFsZ7vw8/BieVmHMuLlk6GeZVTHPXDngyI4VEm1/r3DSi
nB/WUSJsYI9akkfAdHnIOrHaUbtDZp+AY5vGDl8cCW/bMbNnv/EwA8p+m0aOQnXk
mXsH9UNR0XY9hSdxn1uwYtr5ZeXNItmAXdkBwlFSYdgicEbk3qOKyda/naAb20+q
SMSFXBgcDNIx2bEq6J7198cRPx0PWQV1IXjR4xGOBrzzgDJ2mmdRNwnR6MpaBrqm
69wfgYhUiaUoLyl55zhlyb4OGsrHnAvD60ms1JCV31eLT7sa/Y/2VK02mnrtfBbb
mVDqehqvMBg+8H0TUo0lFdvTsi3SrLnsJiiGY07+mdEIWnUm5eibLKxzieB7+tDG
jD1//hgx4BqXeZy0nloREgGC0bFRsucxnTiYwc2NQaCoj9yZhFI/AMeBrh7L+WcB
WJQqrwzNSu6yZs4R4FiqTs7EpYSngLqQGyc88H+/7HzQ3ET5gbcMkp6nbmV9ZKFZ
7b61VgI8LyLl1fe0vY+lkzN1KjHL5Xu64lkeh7l3agx06Kod9MtQ0yKM8DiYbm7d
G2epfihM8FAHfpMb+gRxsy331Qz70+MVIHmfj3S8rwEZ73vJGR0CiMtbelaaNvUH
P2q2AESJvRIF6Ka1ltibiDFi8lTqtGNc+7gb+HxGkLuH+SR3zTtXzeyqAVxb70Mb
8fLNTmBxA8Sh1U1APKsLUZtl03WcPuPWlkAncXcSEHPrjy0yC19dx1tk140b3qJX
HwTz7GwWk/bjGxDNdqvoLREH7y/0iEkOhd77ITf1rsbi3SXpQgc6rxFwSqMz3MOk
k7lh4m3EWUa4NVO524dfVBBzfzG/VphQhPwcTgekPbxHnCuREWGPDfiH340ZLpyr
r89ifjlL/kdasE5mOJw/H2NXwEhzr7FJvs8yTbioQaX/CvNmJJXy9vr6wLCFrcy/
w2eXIgLCclcATJ5xf0AZnH516X40qjOq1QA7d0TU5M96WreF+mJ5a+H8usWcoaC1
uaRCDS6Wca8owW0nFTaIO3Hjb1dfLQdzd3Dd5rLMD21YD7rd7kAv1zHfvbWvaX/f
8a17N1gpN/qCxfNiauWbzyfFV9EVhOAmQxgCRb+vdUhkdZFKvm+ctziajReJnRSw
gsb9GSNELeekAvEJdmM/fzRoWTQ/af+7FLGkKOs3DgsyWsOs2IQP81aRcome2w+0
ubTZZj4MWx5zLuezNYdK6eMzAwcXCE7E5iyQa6JjhXvI67l0GGGRhi3OXwnj0n4f
X4RybFyeNK18xQJgzYj7nEg6L57TTO80+Zc4dlm41tLJ3oPDqvc4MIp1awBydP1Q
S8007LOh7rUD+9jxezdCy44K8W9vCwVbEJvGgUM3NhSEWi9AOlcz2BJu0XCKOOPP
dzmGeF91J7K8ArQOPxhgJZPQD0rILnX3H2vjYtQ5B6739etkpI1zNJwHuMyc1GTW
relS+LzeMe9pa5/Ua0qHQHzkXk2CTOcMci3TiguI1T5qbk9eaJUD6jw+davAg/2j
FlV6dtZWPKF6xTMFEXJtY8uI4c3f3JeV6BNA26/Jcdzo62q0jL3eVktg8KOdJmv6
74UY184cNspkP1bhtxRFdWNdG3iKITo7TXlh+/OPh4herlvQxJ48Grz/2kO+Qrff
m4/Rffsj5RkLlSCc6UPB/boVc29jRwtzEIBbGuUF6bDhglQdWL/TcxLIjJ0cccyA
s1BgxLJGAzjhndq7pLgX0IEOHQYW0wWU/V+WY5MuGVL0bzF1cC4wgMKPMYJ0D3ij
+FBATwbKK1lUG/NHc0hxHvbQfcL2f9exRk1Ctxnhu84L6kVWWkwLJCdCX68A8CId
0FifUSobfRkV5fMCaqadA3t7i0zFkHU7emaR7ofJqIdec+EQCtzXD+3iiyb4TnAB
ZTrujFt/ZQaB7fRMKejL24MglHmsowUsS56eHa5UjxJpxLWE3X8DwEcd6asRSjRm
umpYctO5849LZu1xatMOAlKjCHi/kL/bEZw8US/IfbwxQzBrBX1ettZ4A5hv/N8U
8H3lyRnHgwMkK5spch/fHJHVkzVE5V0M1t+aVVBf/KSXPSgqbl5a6TPYQG8+A2Ny
ni2Uf/B+LQNdnEXB8kkIb7s8phldnFYavkJVHjYd4NRRqAU+CzQNQV998kd5k3Vs
9jJXH3TgDVhlGFchbvZfioi+tLpjhqPnb2cqgQMg102rkxHbhmOoy2lQWCQizUAb
r4qDsbwSkntXBqCzrnd090ldrgo4mxtITm0J2VspzkPRLzbXboolp8RC/lZKadI1
Dz74KSc9BfKeaczg2KnZzz0CjnxulFMk9HxF7gNyOxvnYHiu2+P2IY1LXzaVimgo
EqQhsSnwtDeC4cIGyTG9+L3sNS7GhiMfcRlYS7B2gwxVHKwC/nJpZ60pGJgOlK8o
mX0bhWIRrQUK4K+rWLy+2iavNLi2+rbQ+Rjks5I3Rv64InukSWnMR8KLb8nl5FoU
TY5PIGkBxJ5rxD74+ylTjHFdlTNMtktqft8eaRGVWFT7VomXZyGoQhfwVQv7Rnwp
UT4fGAiNxsVD0GyBG88sOGSe91ZgTetzyg8EndgZETDiigRD4gfH6ciHciGmgavy
NtmAiIPXx8WfYCaXHSOkc2icf2ZOWqd89TELFGF8Y08DblnfFclz3kwWtQwzG9xm
gDoU/lfxvNNPvQMev+Jibek0f3VHAFYJozQcbotP+BaabF9/9d6UottPbf3dWvDv
zLqn/1vfquhfhxdn3dNyZrdXEUDzq1LdOx+CNSuhYfcMWm7tSnLPldnCLj/YMEaX
kB1NLSLIJFf9wxSwE3zCsFebL+DVUnvIOVelw3zLkVGCE5po1YjMyaimviEoWguj
t8DEmdpwGYtoYT4i+F7TC29HXl9psRdeRbbcUISa0dCH2EIKE/TCkA+2fzyJ3UZR
Ew1VRd7uz3P8I7TOeqdgdTARnUXwvwtYb3C+I3wainmfTfaob4nCMgedqfu4/o3a
HkmExty4Cy8w70LTiOK45LGZzROBY84zSsW81B27iB8F/1rDyzFKIfB9raKlbfpP
UaLDwHu9i4dXHeAQ6uNv5KTHxarcLodSl5tjMoJ4w3ZT8CM4Ez/fFCsQj7lnrfD/
XE5NE+oSNVjkH1N+EnDDxtuxAO5fPND1z2vKnMS2R1jr4JGAe6mBwup9B1y/6OG0
Qqz9Dwr8BwBy8iG03xRlGuk/dNt8bgkYKHKAjPRj9UdyT/6V5eYpEibYpyKT/gjQ
r7FIozBZW9Ql3/Er9Fnlnt3tyz3p69nU14464VHbopwlGM9lRwtjBhCdP5YQ+EYE
T78JYu50/DyIqWusum8kvpSu8j3Hc4lHTjmgUuTm3x+U1Vm99uUxA+ZUUOaKbv8B
qG3qeL7f5tkNccYyZ0QXhDosFReicO3mE/bifSeUrghAVptXXg6mwogU6t2DFRHF
aFuKWr0pHKOkjuO0C4w08C4zsIYsnfJPe6kdJuGS0jSBc0X/kWfIIJ4eeV7GLEv8
nfnUxd1KbWhwTXBeO/6GCVUTGwaT3fW85rEx9avMCZyK5OZBpEQ/xXVcUdiJ+AwC
gD7m29xBsrqe6NFq1imEU+zmqyK/Y3fR3FbOL50qW5fDkXMVNTM2bOr/blNh05gN
8K4F+PEt6iPPgI7emtDnyjmnQnPrej54tXb5IZUrMwPMc+c00he0Ub8hH2gaE9cL
8HxMppvR62bVkB6zcm+L9CvzI4qbZ4zZlIDtkRRRdpKeTWGUqzwrXaBJWmibsyW9
oA3J8IZLphk/MBxMxRYQpFfgRHE3VrWPJF/iR+pbGWPs3kMY66rw+v/J+MKSYp2d
XcXlfbPUw5/rnEe5dW/dVc4STSkf16iiK6uN5jPiAv38USBttVWt5a8tQef0QlQE
xREHAXhffkitc/QZXkBYpYJ1JV1XP3aBg94aYlTXT/hxt9/++5/Wlj+KH25p99ov
FHNpkbgt5BmP3qWdyfTVVVWGlJywGaN5kTj2gHAhzGFrr3vZAx4ml1duCMe/2ML8
SuY/C7kr7DGIDNqbM0wkK6G9j+DFA1DE06VrPX9QajvmMLdRN8uoX8B+b/Bh/4QI
mmgbCShTXc8mnIRqGeBUOwqVaMA8EXXQTFowIYhfyVleZOhRIMDaIgRnqHR4AabX
4CYg/TeclqviJvzflSQlRo8hV43zyZK2VUYYk5oIBdaor63GjopntDVPsQM3n6Du
niFiAXPgnUabIDYJflMeSbWcnN8bLKS85yiM4h+1Rl0+DvBt+49KdFNS/PH+AbDL
z4UNFXRs9x4UA8bjY5vYIeZlo8xW9FIsx7ftaJeKfnqaAKKEL2tLVd+elUt/SZGa
DVZ+BOxTgAwqjX5NTuTho9iSFV83k7PTypm1L9tczIavmWvACL8IG//c1ECZ3F/z
mhkkitN7QLmKc1KPsmX0sgfeAFyd8q/r3p7UBiLB2AZi+przsX/qtxPgGUcbjq/c
9PEJzxqU+nc8DPY8objYHmSbU/ouxHIuMpwKkpFZ+GrsaF5SoVDawbXnq845vlWM
RuZhyNC8Li6rNYudklVLpBCR2baFxguZjfIKgQeIjNxJOElpOcodZCAmRtn6kOgB
VD6xfhFDwLSuImDdU3CdBhTrobU2BRp0Xpu75eHu0P1TxDUvIGalSCKrVuaPu0qs
Bhiyf6zQeCW4MhPAhW9I5FXRDon+62Z1s/wuAXBEXPkOrW7zxyxsr1QO52228lIb
KBTMRTTXd6Gel3/eKoOXRnpfN74z9fVV2+U0uf1Wtdvumf65VavLolDCaI0II1AE
BK7eTkFoMwkbLEImZoztNdf9CQLtDOTRRlzyiwGN0+fAp5gJ8OGI7jFeK5UtH6g1
Cfp1fgGSw8F8Mpb5QBgUgVIowFMZveJ/bhlpUOjlrSp87wTcCBzI+1QtNuaPr0S0
xroGDw0gjTfx4jjvEFuRFQRANZzS3v4bNOQVxYSRDhHXkMKFP9vnddJnE+LX0WnF
Ct5PLmeh0BPpINO/y8BDG25UYU1ApkHKoLvk5njfHOMlEdSTeoYeTMWtm7KrX1hv
/y7caWGVltN5DwM8ueB4nAToWRKQu5+fcL0VNCodiMkUKFtdMepJnifCaIm/hx7q
8mXkNUPJxI4EzEskpInYfKBbG8vQj0BJ7sncQDmORbzDMYMIMPTu5sQtTSt1A/QS
SS1+986FxVunSIGx1vtCktHo6cj+SSEaaW7vdE/evfAtTDew1e9S7H1WSotyDvws
Auhh7SWzHxCYcZWcdRy8NT8/EEEKy/BGAhcPIV8qjgzj/mMwv8QdnTOGOrTNa9j7
9EAgXLDhXl7O/UsFC+KplVTxEiycGuQayTh7MrqiaGRBV03Rj0ZPkm6NQzeWhhIG
YbqhY0LUtdzbzhF7kSI+vX56pDz3iIm2z+5+YNVT60i9NkWY8ApBs+6Qj8Q6C3Tw
/9nxjcOQTsAa8T6OXuTEl94xM6ysb2HgcFkDAxflw3JYDKecZvgtMmoD4u89ie/O
VJIG4vqXkOiRRf1IKNNQ1C6Ky3myVipS610u1Gbnyp0sQrdDMDswRbfkstHfPNJe
o/BGNIZbLDK7tZqDOXxtOd38uFxBTRmGxgbs+z6ZQ0VELY09YHCXknU9/zRGu1xA
E9FxOcINNzH176KvzrsRGPuTzOg2eSfTj6v7IjpVHIycRCY1hwlS4kaE8R27GJ5V
L7TECPlfLa2tnjkY/Lk19Qn3oasmoeikfCnQ2FI49GPkLmwqNEi7OjjFz1PgkiFH
47vPzGP+DqPqNwNKN9K5oBWXvxyFDKWTnliQnrtFe7JzM6EHlMIaxh3Xd3Pv0B56
FvZ7W4Wgd515FMbsfD8E4I3QdCzExOZIIqQZ7sYi8433woR4ynZQg8bmu6dbvTW4
/f06+e5Miyd+XEEeWnoRUI39I5w1En+yYhrDKJji8wZmxqadUszQe0zbT9sn6io/
/NQ7shgdhQCt15oOaFGb4nubkrkBdjhVjI38sYjsnvXVkoOZS9ZRYltsmN9ROuqw
wNZqY9PiTqmd/g88iNwe+ghCVxrW3YRuohZj2jpO4rJz/ThqBFpPGsAi+FRGAk6e
8BpRyKBne5lB+pSodeagqBrxzIQnPuRXX8xXlABvbJuZbV30Dne/Rdi2WsSAXRIJ
bt50fhPepY9jakOPzGh3up+eBAnxpRU/CAaHA6YKyDylDg9RQec8+Rp1me4bvsln
OqUMes/BKB/2FXh8fA2pY6iLUzKVHpHDozgJMvxgT7rRh+Gsr6m68LTIT81Xcsm1
1xcBIYjlNAaHjN4LbVzAyhwl7IhNQylogSF7TTgC77RfSDoz3UUj5roZu8zQHUHN
vLcdb2ewS3hLAlBURebznr6WKqzTufkyq2UQng8OjS3FoMWmAJX044X86icL0KQ+
Srr8qDU/EM77FtiD/K5dAgoLEL0ohwy+F0onS+tXKitBwWNSTnDAiFU7TBPLiDfD
sYeywSr5WRGehJ3enpgk9UznpTREGtJmeRTJA3KvOPorPdH1oTuuxBbaWl1WOOTA
F5qtAYO3inMRydosA8Nht9lEVAAELQ9gwuojwawT86fJrxx3ViYZKCm+yhzJwcSK
2JO3QUaeKIIMuYME6Rn78GVAiCKUU85b+uuyJWar0ndSqZyCwNTJ86o/atNFZLZA
dQo9H8XFCY1GLIIxQvLGnMdNn2Tb0UYn8MaF4F5vwp17ITfRoDS0BGB0e+Tsk9Kk
eAaEGxzNuWmN/UCgKOAg1sVu0bHe6NDfMEzv4WG/TY2qUKTcVwNALNdG75DwWsI3
UNtOMM2i0wuw9br+8lIsWFEP8snyMKL8rBQFigE+6VsBDDF70l229neFd3FsIZPC
4QfUO7G/gHeyIW1Bb94nkkSCMm543qBW6VXKTibWsZrFN9V3f3FalOVWDChoYK6c
GS0CjCHSf1Dz8qYJLquy7cDZh+yLjj8cftULdvwOYAJiBFdX+KynxZoEDsxl3rC8
xHRrquwOvVGyRL0l/z11em5CBiyQIut/i5+g2A8t/HJIDUEPxZIc2NBnpjOu05k2
eeQ9a6v3SrZdTpsG96qTqCrU5OzprQvrqLMGSgePWqZk+ObaCBUGEgdH+V98Wdq/
/paf6N+g1Cdo3uua1H29VEyAQViHh3+ZC/GWbIo8Ui6p3PxkRjrMt8PVV/p2YSzo
Ux6DOk7JbzpqzkeJK5WoRylCsGnzeBcsKqUHD/cNL6egBE3q5nt5W7VX7L6KN4Zg
/3bJ6wrb0Rly4SIqrsVmyE9qS4sNbZAdxlHbnYT0zNztetrNDU0/bRJeSZz5nX/S
sN0itKPXika7rq58hq7I2KFQPHe3UDjJt6VzuWd0/GRLITBkl8/aiXSh/5/q7FL9
N3EnMUivt1GjZ3Lobt7ukdIx8GHDbyDdLLiSSX4MeerXH02WMEoaSuQtpsnH12Zd
yKUbnuBCkokTwANWgihKK+s6URG17YVtlMIhUoHSewC6mEvw4uVrF+IgDvwBHEw1
qNbAIe/grEdOOcvxynBTUihcQSbIlrY6sLUaA8m9FFq8o1CeGbu/w0pvV3iEA+p9
Ti2Z+x7tcCq9pLz7xmTUF760O3CBWNK4KluOGQMrgU3Yowj00R1WzR3+3zcgsVpq
QYZnH+oM9O2286RAHDdwCxPdape8xHoBh32601UfLj+YNu5b2KqkfoB9M45zaAHs
G/UxOuxRTzzQQtSHzaXq/ogGerwHRc++S8gdyGJNuEK6Ohc+JFi12QGO9gbiM/UJ
zh4j1G2kbOmWzf/Fg/rMQiWywTH6ET0QU39/VFnXaoJr0a1Yjrh8fzKSYPPw8Ftr
/J/lfMXMkpxYfFC+5FwDXl58XQCrzXWlcbOO/gPb4JWI/D2t+NXRchhsMDGjKXMV
plI1YNsRv5JSXS0tiSY930C5zAIkw6GoK+K6Y5yNKKm5RzgMBmMsw13HPw6lC0b7
c7kNIm/rW8zo5BNbcXr1hWJfvBZVRZ/NvFabxPTLGDj6l/TA3V5cfet6/axulo+U
zDl7yDmctZESNHQDAkWEyjTU0NTkuE43x3G6YQs5XYMa8dfbdtf6u0RgURBBg6PE
x3fj8HuBeHqtYSkQ0NU1x22mXIvMKEhosGWq9dLU9W3DVuMJgVseqhPrf5CGh88K
DT1dekX44ZQANUq1dx8fcYxXkstohS+DataNIuG+u7XuQ9bjvuMWIiL6M9DLv/gI
qqq1ZMTsJ6t5STU6aYFLrW4TfPEpfL/E5cJ9xVf40cZtrhtywidZlkimmvJN9sSl
41JW25iFZeHNTZHfSi853PYfhJeO1cL1IgYjF1ntgQ95e31g979TE5mW8QHif2mC
AFg/OhyaTxNkbtvMYFArHueggdue+but/cStQ9R79pQCpT+vq1YLwo9vZtet1aoi
jD58DpJLzY0EFz36tILJu+dnab7yJTEJGaz6qulv3iwNYYStojqOTAKJOCNhxJgo
sd75YAx1Q018vhBOTBxugBlyJ8+0cv1BHMXuCEiRGbqvcCQYN3cicBnceoD5mxc0
aJXC+Dzubp1/V5s86grYn7v7D+PUnbL1P3P5Gf1O1+3aVzRmsHvTEQzDZVXsDWZT
okG70vljKqzIVb0ZvQQEzt1JbIruqNxZQkyjnUWfoUPDUrJTQ+JLOJGnSpV5V+YC
8W029rQ7Er0zZLYLUCWbUBVwAH4FIEcJ5E3CE+of7HV8L1nZ6Rl3DHy+mFPXr3u1
Xsqd7g/9R5weIu6diVvWiXPIxCt+1Y/1CP5Ko6rTr2mAEnJGFsq6lgBHzew8/CiT
nlPIdhUnZS7jYFsMSP3Qsak2aqxnNiyKuP2KoU6nq+F8mdbIfnTgifXr7BOvapHD
rTM8TyRU0KHWo41ZQ8vVAgsB+sXNShvKAHqxAYiOHwj9n0GszmF0X5VCwSB+Q+ew
3Ug83Nr/fJ/9+N0ebtTFhromqMKpA+x4Vtud8OxmYL/EZ7EvJgXVdGcjuOD4nfQi
8HmPQIi/kTOtMEaMj1iVzBisQ9nEz+U8JQ86BRs/6vMXnNRs/jrBw5oJMhDcnq3c
1K/BI97W2FZ5qerDOaCt8P8NecJyE66TObyPL0UdHuB1WAcbRphqIBgLXHeKXTw3
gStr+OgVaFJPIlSxJQCqDpjAcpTM5qBS7rErt+MHmtDKQpVx7INCk392UL79sxj0
1ZfcMfwbKOc28aT2ZmA/Gb/5fPSfuAaiTtYPmc3/EaIEPk0C0n8JbCZ4LVSpQ3fL
nVwLBpwKoFosMUwPNM8ogmaiLIxHHPp/ptjOoiLLLGZFh3HjdUkmU0gxUwqG+gGI
bdFLXwatCwZPoI58A+0rpnTNm40axpIadO/j8iRLwAcb3JlK9hYkjsodbFPjHECy
kZiHiZYIWNqXWC2XUMF5im0foQ/imSFV9XmltkGf+XqMXVHSEtCq97Q7mzLENVnN
bccIdxX3SbGPWRewzawsKLxMieVhWy3Bus2C9Gw7fdPpYaraRPYJS0MyyYqAbfDE
lUrtq75a2cHtGhKZeHZPXUhWjBM4ptIZHk9EOcTqiCH+9jDT0NvEZ+ybhqFjB6X0
roPgv8eUeRMXKm2imsjSyEsMot8Mb/2ml2Ol1OLmdvS8l0Hq55fMc+bwddnoSUwv
UXgXqojzRVeZ9m/rXKR/eokdUY7oAnAbFY4DHyT757b9FVe8Xi9+ry2fgK++jfZP
6+vuzeLvkll2TgFJ1sAAv1xYxV6bv3EI4wEVXlF6g0UyN2wVvPndteYQ6nA1DYAo
ccVH+MDS65I4TUby2vaqv74Sgc05UJv3vRDCEiq38JDJwX7Yy7LyMOyl3kos9RW1
XxrWiVViP+RMXHKMyQO/xa5x3CuOkN+qTYcTcKGQxNpLpi9mZDSe6ldSKScHgVgQ
AYalAp/4DEG9Ia0Bs3oX1Rp3eqvyUB5ueKht1alQvASWYDp+XGTRxTeC73esDbAj
1KB+/h+ZTwGJwy43dSt1npbaRJ74K1I/yBej2Nmj8tu946MtdndbSfc3jBSi8neP
Kt3xQfdY/kii2tQbo4civtCvHFQkcarRQ8qizqYFqFoDISQ4hlqAS18qE5kvMERv
1rwR5bRO4gVWqDTMjwV3UPBbCewK/9wmfCSpMoresqpEb4YI0Q+oLSis93vmjFKV
qnAa2tOIG68dbRqW0RQvftHKccKPUTxzWs2/d2mFGp+DZFawRUD9U+qlxIIN4VaB
oIFm6Y2WCox8buAugDaO8V/12SLOlBbCxC4RtBeNYd8yL4iuWLbBDrJLvZeiZnCf
jluohg5kv8kC5i/lqRX67PQNKZW9rpmnOBLRS1nNtOPeRrkqfTU+2RVJmNKJPF5m
G2jttdHsuvyfEI/kkb8jAHQs2zz5asPwSBCnLXr6LNIIWxRud+OmXFr4VFclgKQY
/NJ0MIONciXNwt+rCxC6LZ0LAPM8qG8mt9nc2laxBjBMwj8XvrFyn22DK5J8KPRR
7tstsEZj4BYnDqs+WtB3n9vii0WHEhmmyh5y2RxW4qzfwcE5EaTxXGi5hbUIJXH1
GdrAj/rbfTnNYmUIDQSoBfhQhTk1uJ86rRZMiriwevEdog5FZvnv+DQKGHHR5Qep
u4fWc/TBHsnYKOXfRNeq9JEWKN+1d0KsIIwtAAWwiueoeT93uoGMaLUF8Ry99mcT
0xxkfiMhhWldqSet04cEf++ezFVd7rscTvSxWmzGAk0jbB99h4x43AIiaCB4y85i
wxgEgsdnVXYsWHIJ3pN1tlkrRmMgpvyGa3oBtghupQoiATz1A/4XVWUYnZVJYVgY
ek8IQ12PcQAKHmf0faTkikwllLcTsd6s1/2PhdMbf2+zmf8ehk/Vev/laJ7JCtTN
VQ2dqF6N0k3I2WtYzy8+pvXT7bJqZv2j9kpCboMDfdmdytODUvLffdDpK9XJViMr
mS+6Wkx4NnMW8Hk9Ng0N0euRTriyr+1nj0XQvCSRAMvr1B1B+WV4VEdi8LtiGj0p
affSMOrfNbbEe3OkXFxsyfeeElQGjP47zhf+HX7396WJHFPYrfurlq1hw8oqx6/H
mDV/9uFg7Unq2coEOVxBH85XVMCxIh6FBlZ3C3nYoFoEuV7igFtWE14etP/aWnnd
B6Nhgp/1T8DzKOEu9dyKu1r5OtAdn+MUBftl/zX+6mCPCqwlvhgvAIuycmPQjgSe
gTjy7PveVm9IWL6gFUvu6zkVet63smx2xbKh15c66P+KhZyUmIZxCA0WFeq3QtRY
V2Em8bzUcd1qRG6Y1GBhrzOhHRzrclhq40YZTWaYmGS2k13KHOasKP0UchzVJuNI
Mly5WtuXE/oR5ST14WozSeTltAS1cAZwbnT7fAFuT1tBaBpO6zhx44dcxOJESoxI
noMOHqgLZ5n0mxfAc/3NTXEDIpomejj7Tujil5ozi5S/tSHk/n7Bta1xq07PUsUd
DSLr9m2DQwCSUyLfzbXlMtaGvBlu/3NCJb5KBEAxXTQOg1bpTmCrjMV/coA9Qc4f
mODDJsB3jjSzidXNxjHKzsOQL//mDsllW+F4mhA2v/bfCm6QZJLmOJP9WXgEF1+C
MxgX1R3Dp5Q4UqVe5WmaR1H8haHPx14gGE96KCxD4zmlMaANmbgDPgT7aXUtSCNs
54YK0j3MRgNw08TrWjT6xPxI+Fp1s1rFYI/+WAjKIWTHM7Qeymm84Ro1DzgwuyE4
ynoYeG+pfye5qnrnWR2+RLatGu1VJ53qiNzi3NS26bF840aQ9r/pudVKu5D67asI
SU4eJlkXb0niOHzSsADJ/5A9SKqb+d2lB9vIE3pF/kCwkUgeuWCc5TX9QGgPXqIi
1ebUPkweWRIgdXXG7A2eS38El/Lu4mcwWjLTtVVy881xiwJdDa7twUhQAvb0XUq8
MFSo9CwCghYsCW8ko9oh6y4hLRsG1OPHnmhu4gv1F0vdd9DL3AXUwxpTLzvIo4in
HW7SKhJDNNqmyzOA6NgEOngGgKslAwfeS/Bdqjll00++bn4iLgj7vahM+U6TddCD
m9YMHc13uDZ7cQvc6DmBzK63vPhREEfy67+7ZFbCouRmG9K8lVYSk1a/fdPxK3Wp
1edeTkAAp8F1ksfJSyqzKK6Zn81vt4z32/iBaSvAVFP+1GzD6X4OWJNtPjnZgyk4
7IwYWFSNTeDjHJG/wowyh3rijiteuamN2/qS/H3XfI0rG12zFazwHvRUhFVjI1lS
UrLePPIj8+NCNJ4sqyUL2UJ49PCTBepw+FkibnGRRhuKbNYSTWiB8CXY2WLEUH0B
rs1Xl6T88jzdG8sZgSBM0TxAGYwbC5RbyZHcywJhupuU/pFeC426eDeaitRKbtxE
DV6TZmY2hWaSwCbiqIk8WXXRp9LjjP6KLL5JsdJhMMm8bUzKpdjhUmc8ylviH2E3
JBtb1NODjTCNmQBt5iIJhzsTRACt+bs7VpCrFiI/bjVjL+UaK7719btP2NWADmGK
7nVPyryRJD87ZNf56DC8ebaxcdz2HwkXiY+PmvSubGqlLmgm+bIQ94IO5EqhGPNM
9xtMjJq2qaxwtHJQPmrdlDOe6Z6yF39BRZI11OsPELH1hvPuBqiSg7CjmplcMDm1
1Dx+HlIp4Ril8SsLSbjjtYm8uFm+2G4Ore4ya/GBiB0QVuPVUqgIqmyDPlxP+ZPH
1/NhsdksOP0Gj3zqdye84/hSlEQHE4W9hLKDHdUs0RcMFcnFgeNf/eLEVEsMajWa
edbcZg4/YIZDTZBQxrzX2hke3QfP8VEt2m1dO+gclZleKOLExDxgQDTX0Mfxicgp
6ZQS+5yUNPU3N5WMDQgTzKmiS/64vIM/sRVu4ajx8KHUbXzmcr91lyoO9CEPJFWg
VmmBesY9nzahRCZEH9AKOpNcxH4EmPh8A48oB1WFkZU0/LR8bQeVt28nLGF53xA4
1lGlTA6/l4B0yEELFLYJh5sWRZHqLS6U+eZx9hvBmHZeOTXs+Qflz1bxa9M6SYOA
PBkHdG17BsMoCG57vEPWj54waIzbFpRrcGeq4qqO20VCaNW5w2Cj2AJzutSSQC6z
gnsi1d4no9GvScakllXWk/WeP1wpHwvWtlBkABrZaNC2UyLHh2wiRSIf8HVx7lgM
92t8cHMCqd3uiQn8ZuPgnwcGqo0WA5ljp9syy7KuVaRSobCRvL9nqsFDdfXOlt0n
EXcoUw0Jk9Tk/q3fZe+NbevRVE4XECeZ/lJEeeYaOPY0ZbuMGRX9rtvlwSMIio6T
ogB/Y5sysLbrXJmaZGeRBz/nbpFurx9YherKJFG5T60OU2K2LpTkRcMgzGFoCkXY
V+p4kx9ECCuqqg1n8AhgypKp5dlpFatMsuf3M3wR4VfHu2kZj2u5zJXQYQMgydu3
B8h8C9/UrDq2x3LeIetdsYVr74kn8cw0FQxsA+TzqeB9MqOPsXWja8QiXAT/HGhd
iy67KeapUuUazRibtze0QNV8DCIjMGCG/l2V6CKXTZsB4+j62cICigYMyU56hRHL
lavLwARgRaXJR9I1TSA8wGCwBBK1eUs35fAP2ne2pjqAoGOXHPZVxokXEj95/OeA
fuINF1ZjTY5Pv94VM2zOscXLys+UeYKHQ+UZ/tKjz2Xl+Ax5IUdB+brM5OUlqQJz
WE2ZC0bY/2RUvUuI+RzfM4OqX/sE9F3oPWSyBmeoVTQCpJoImE3QBrV2sjcNPhBS
AzPQHA8vEZJU5vS7Q3b/4dUhdrcl44zoBKO65yq1BtqjaJAS0lMejm+4xt55pBsM
fn2xi4ED9XLYRJfPQG530xNmab8kUVZxtOeZItGgVNZGspFbZd0s0Z93svDhgWW6
TRcJZhju998O4nAVqzpXwMavRloNk4kygKjm6xhrOI3D/ey4uZveSq1CXKNY0ai3
4bs2K9Gqn1gCR7TM64JU0gv4GJroaSgdo5iGF5Ym9SF37Ee1vdhM874CuEzfxyZq
bNYDVrRGmY2Q4dThKk839vLf9RhX1zjy6rdKJZrd8z1Zxq26HPtQuvuV+gyz6FU3
EiuJx15RqLDFz9HGWstvHd2KZ+3ZH8aL0gP3jUEqyocSoN+g244j/OEFzA1nYsPM
e/2IlP8ryTOxaaRKNukyHgvvlDx60fXYvoEUq62Plua/vARh0/Lo9Wtq1+i3zJuT
/+HiuJ/tleOAY9WXwc5ew6uJ+rSaCzcd9hrUVZDVgraKYQA8TMZuL+0/Z6SV/YIR
9ylZQlDCx6KVXnWHEZ4wxR24wt6ZYz0gP1enZdSl+DFVgLNb6jgC1l8QjBFoDyJV
v4HtoyDoVt25edTMPiHYL5Px33NvR0Z9HTCAHmLNlYwg7KtOffLMTY717nsGH99G
lZy/zDEEK+wqkjL+wJjqWS6M30nk+nmC0bibkSetcIBpYe5ygxXtRz4bWjFpnCXL
epD9K07FrHvnT3/KmATbuSwy9cUUrlo1LGJLmIpUHYCFAW5a64uJj+Iajqi+oO52
dx0c22Zk9qzJmeLuzrGxWXolGkZhBTk0gE4ZuvR1W1CtiIyYgvXk4WntluSCrOzt
H6lnamEELTVfd+z7t+q42NaLpT5m3ToDZCBXNmr2MRjRb6wvcKVJ4uYTBEzjlF2j
O4IWsdWHkBu+mkWKH2V1dmxfqeWSihLZHUUiSRSAsYt47AqzX8cpm2TGUNl3VIG0
MhSWvOv4dlMTx4O58OGLYpolH49KcP6SHhfFrrvWl/YPDyUXZeAzUi0tOdIFgIJQ
OyQgcpn7FE6iwP0duQFtLm4PCWHnDHGqQ2yojukHPoK14IyGSq6x+XWDh5MdmTzR
cd4w6Aa8AxF4BxG8n9ElIYiwTuVd9on1jaeGazpfSGQJ0GWzeFwEbFhjJOmS37LL
KZwSMsa8X6vwcn3c3LE/e4jkCye0c8KjsanuWIF7/rjIfOlv7K/i4ftj44CghaeR
uh3XYYqSyCYJrd6kQdcqsOqGzTX1q/err5SPDzvpnHg77MpuET7czVC8z7bagI58
QM/91iTOSY196tJjVGxFM2ksuJ3T3PoLTlp8mnJbwfIapUBzdLoLupzKO7mHHTwY
ASwlFiTi+1+cTrt66AUFKvStUri333TOli99chDfYXvFrpY182wkUgfzlkw5OGxH
Drq3XOkV27QrZOwpwyswTD5STjptAhpZuzi47NqHSVVoSfr7td9nt7ZPCMq5Fyzj
/tSIs8FHcZWHfO7hQa9aHD0GHG7UF6v8TQBcPUJZAy8h9eJWr5fKc8WD/hcXZiPG
Im62kCBww0YVOXv8b+S/y88ac96+hWxwnX5QS26HyDU9c5y61gXDhHm1RQuKPYFy
q2mdmYlqbRHXiIpBitAQHsyge323E/YHmPv4+bMguh0rASuqdV4TsAROdUvq9/yh
3mkv/0gEB/gbv6Vi3Aem73gs+WGkt+4F1sSTgu8DfctYdZDznRkOeCnQsrTwRFaw
9fCpCdLMazVd3PQjNiHrZPd3Q41PP7tQcuNgRQIpgUXbKYIbTLsFilrOKppNhDx5
Qbx39CGR8YbX9Kmm44RADFHdPcj9Gm7fhcdPu+JDcjprWShlYOq6QwfjffiKsLMH
WTXDWGdkt4IIE5e5WpDorbaKcayxS+IfjJi+5WNi/zA5FuVj5g/iB1IA+vbYt1yS
cgFfJtYGZSYxA87LBMQ2avzSzIF+IsG0IuDlDoWPPHC6BjQ+ZiS327r7hZoTGFxl
Gk+QbD4gAMXT1uYzP34UOGdDdbxXuZj/HWIAIjm9eCtEHKXSMEyy0KPOTfIEIHGC
wg/GGpX61bQ5ODjNm45Bmki+i1iBFQ9FLz97GHya68x2HMf09RBEeMLlVhWm6sML
o6+m7C6bCZmuMxDrNABT//+Zd5vzI8qAMBlvexHnOIfp0A1Q6M6SljWR+CakkBq7
GLZom5ErX5GXrIXyepZbDgW/eensGKpWA7z5zAX9SiCMph3AO754AWCLNs4k5fG+
MOq9QPbq8h//mYvTbpdxYhb13TbuRLqTh64IAll9L8BVy2iOy/HRp/60NKihFIcs
4yuLMjUPpuYHYetXhLNVWTvLJyFjtqaNSaPtm4uk2CrwHixJc7F4r++G1rNumJ+N
XOfIYsod0kaz9bDCyjzOkmSPCrhF7ikZsFup2vuK1mSNrec6H9XyKX6ZegQfWlys
Bnk/rZmqlTbzZkG/UWcfBJhdmLGP3o57rof8h3/pya7Eoqw5+A65avNmpPyRtnDX
sBvgO+LwmBEEz3NtmZ6N9xgGpKGuiN4E3RCLvs15n+4XPbVbVcMHXluf+dUMBfxt
6ZmC4CLVo9WdzJZRR7C4aSBsff+Nd1e5EMf9K5WF1TDAfRdBpHvcwQVQKrs4rwrk
fBsGK1KKGY+R2GxET414W0sDUYLY6qo3iZ65ZoOeSd1Shx+0mAhflfkzvCml607z
TcQpVhXUvz6e9nMD70ErByThBx+E3g0SWbiF1TRFjeCu+qdNbPWA/0VEsohjFKhm
TP9TrAO7HM6VZe8Tk6fP9fHEa9VSCqmjel5llNyS4xUxxS+HZ75o2Gbq3CxZuJ8f
rLUq/sppRv+AVyvx4z69X5q/V0AkVQauH2NtGUYB/FWgI44k9SYccUGWsEWkZtVN
L3abx9oAsw75iUz7jGF7dBHiDICoATtbyrkj3XihWZvOtJmxn9PPY14CPo/YyyRP
o3jkHNptIJ7ZmrWcV6hEcYYP+WXMpRZeYoyNF8+M7uxvNFj6Rh6YWHi/YX73uh4M
Ta8Wv1PmPTDXcHUkA8n0uqF0PNhlaB/T4utHlLNJ35kzEdbLoY0uS0VioLGXebLM
EwLkIFb08mlegcZ3yV2PJrdjCjvRKBgQV6mIUpC1O9a2FhRR28Af+MJtbRbm1WC3
uwkM6A0rPV+bpr59grmkOxuB3pf5WcZNyqMYYbMO5vSNPDdM6HYxyhba2wfH9bSL
tf10VfvlxrmBvaSdmI6vTck0yrAPIKwmNT/vlboIpc4Xg4siZurfRT19De/QOmmL
KuEVoPYjqJLwJUg3kk3fQK9PDWVs/ohhWMvOCzt7Iaygv/LBWGX/OnPDYEgl8I/U
JkS8C/8Jon26eCiqENdPjgtjs2J8g7eMGQFSnMfIYLhG+CshI9Yv7A5PyjLLJjix
xMcl9lXd8thk5yiM3mhG0H06Bne7WHwl8JAjdyaJxDKm0yonQ94rSppiquyU+k96
wGYVIeqrX+tth+jhp7p93CsKOKjY2StaAhuGKS8kP31Ijgnr5N8K1qgsGbkRVfrC
q954MTGcDM3qTcrC0i7nKFowUp2PUhe649EqPP7GQxvmjcdOAkpEoyw6zhLGIiVY
5daPaQxKS2oJFwE8hz22m+2Z1O7KA0DPEfk2HxYNsXTZ8o99SGn5jiz6PovMU2hQ
RefUzlBSazlktAGp4pFJBkUFRKiLiH/PliN5G4Dg7ELQZUnHDGewgIpqIAVuDnAQ
minbzWg9bVVADl4kV8Ok0BjXeZERIIK5MEPwG+ZZE+kDGVPDkZct914zDENDbKeU
3d67TjjaDJA2+m9wNb0oCrec0RZjJk7DqnJCeSLh2AjA69/1rjuA0H/5pJcjKc6a
7abkKRj3EdsqQN1/iyIxIOpw9/fJ7Z3Bai8NFvE/SXhja1S2ZT96cMAjWZV6Dy5m
WEAUk+M3IoVq28Z/NFpxNOBjEsxAcq5RC7vkwRFbzDPToQR10hKTC8fmy9h3jLxX
SjTDB+rVBFWIxEN9/iVJAZ6qQSdOLR6tgG+ON+X5m2JBTtyQ21qxAPRsHeJewYUC
g2MSfl1Vs27FlatVCRFWRd7SPfEXVldPpyGOVuIdNle0r3pOLHnarzcAch0llE0C
MPJ6mv3+TWflfUa4AyuUWSOdMEfit1NmvRZfOtUlOxMlYMBupynNEhwWFtqZjLKP
YhK6TZmIlyD0opLOkWdQp38fE/h3KJ0OaEzS4JBQjk3nXuXORHkspd6cV3NTnvzx
ztLks0t2IK22ErXFd4tClPKe/9Xuq2zWvmoN7vMUYrETO002QOA9aOkbtKF35cOP
B7CoWLycIAWyvu2gnYSWWoQi8X8oMnGwSSXyGzN9A38SdddkJwEonuiIGERcT0He
aWUoMQePJ3Q9hP7IlbOzfJ6KHRQoqmHyT0V+sgltZ0HRkZB+VKHLDFS4Q6Zyueb5
WXDC2ZvrRY1y5N0jdw9pu4BS/avG6oD7j2kjq7A5f1yPRuBtKT+DhkdC2yBTldHs
mL6XePqWyTKci/tk2qQKx/vpogOft2c8TJKKN762H2aiRZRqaUI63/zOG6eXIGBH
r5TFTCtD2AK9rIngxRB9Z5gGXdXx5v5rnxdPq22zwr9Z73qKWn0D+cPsNqCiuGp7
KscPU+J3UDId8du6hU5QIXZ2kpQPfgtx5BZ4FZo3AZ8fSCi2xM2dwBSGgbwjJb/D
p00pd5EzP8zRSWtHaRovKKH9RHiMp5x2lgF+QRDwPXYJxn9EjFloZF+T1cRgoukV
n03WD7RY/zUSwksK9Vnc2kMKX/CgQlj0bxcTAjuZ/m6BLBz816FhQHZK4bMBhItt
yfoeNmS0Zi20Pg6qt05FQnP8YDtyKRzBMYBVpVd8qT9A2h2kRGgdUXqCEwAIPYot
P1JUCAwm4AdngJa19vqbEYy+d8dI+S2Da49zUFAVX7DFGX12b9EPk2k4iVB6z6Hj
fc1hsEUd3VZYOMtXgNbg5p0rsKRgT8kHk2lMPXfIKb3jfORRsztAuq5d10Gh83ld
IWqoCzj+7J8ZkZyx41MykTj6FWNgB2a4sOnmZrgSzCvStU6mU/M1taXzSEqaRwx1
Bz8wMaR6ZFDw8RA4EuBkEHR5Axk2FggolrEHBAFewHopDd046cDlu1nIl/i+WnIb
FB0lvHGAGryJb1IhsASX72GVVA4dRcPUzXCIeZOSIhy+snL5n+8jqsMcH4AmfJ5P
y8qmQ2PdoFzwTBW05p456vz8efYYH8M51YpbaH9n7Zfy4BipuuUpozsZUTtNnJqD
XifITgXFz2h1azqTN9GVhVB/YSHr30wET/axeHU3mK67TZuti8OmH+9piAht/CiI
1FWv/BDvI4+M/MopE9bOPpJP51M11UPMoz+Vd4vi0SMmrxXeVJRT7cZECpRlywCQ
1vH9/EfSCebn29V7X/WNaVG0lw7MATEUlW+7XwcO4hvsdwuR6aaXsIjgwrMYqu8v
HlGbpHhBfy5V5LC77CRhTPjaJGM41XRGvKyi7hrusMaW5S5UrhYHyYfYznbphImM
IdT97us+5NZfSsGxw/dUdQ96zq8dg8nR0F7NXegUzDUPxYkQB8mF/XSpaMhAn85D
GLPQ4uS55nKusJ6Y5Xkb3sCU5ExrERGM+T/Q8cWQTgFSmzUoVlYNzaGDGMDn3llj
unLsj5+BM8hIfG9O4x1L7URukoPSFdy6DpUPG2fOpoM9piRAh87ZvLiRPszXr9Nr
CK33/f0ZvaRHiesiZ4JYygWjXSafXRN/mvO+GOzMWbjYt95xj7x2OdZzwSJLNILF
v6qE40tZA6p9zHckR4Qn2obLVbLSz/4bBn6biY8dU6RzIUgvb8f+HHiTc7HskPKJ
VWpqOYVxvAZghSLByOn4LT+p5U6Y0BckhrgsHKVbniAGAHNmq6QFtWjNHhlD0cqL
iRpDhy3k090d6hY8x05rcMOCGSjCRw98HAAOr5euJ158R1VkWG+UFbqvvGAKJ+ip
CxGRlJwRU9gA0KXCEPeAXCakRlRqI+RkiIabrJrQLWjNFec77vUyrinDIbVBySt3
1I/KAcawX6Ktq2DRoe0ZnTRZUx5qCXHEFojPON+ATJMAt3uD//6+cpkOwrW5Fpsg
uoxLo0GCz4pmtEfp7ji/RAcB1IukvxL1swVoCA6zDPJJESD41SwKEh8CKQJuUL9h
AkUk1Vz/66Mc5mhqGvmEorKszFf6iXAUS0bEb5Hj+EpYQ1pdhnPyPJB+Ji0rNADg
2ZHOCOryyhbmZ/V85NTYBErYCo6IUQKlDQ6be2YMtv3nrxNRBgehTBTjcpw8+UHS
oPJCJ6LodAo6PRxsM+uvS8Hzon+mLX3HICUn01QJurQys14BrHEn119X4jJPk5yO
BhsQ5H/soL0IGTdfCjE5mDuw4/qrcq2Di7Nlh8BaTno6AQI97jX1sHDGkOzooT5j
JHNjEwQFzVIbO8+J/Rp5mh/klH5lVKBIwWd8EKMn5wEWkXcr4W3GrRv/ymWlCfoV
C30FcLT3bu6t9mZzzCPL+X2dkOpk9g4xUS5DwSvpOgoUP9ZFr213qpzB90vSc9qV
N8q5GGbozYPRPox4unHtvLifvAaIKXpTg6liGOIzrpJbzVpVD3NSwYO742v57aG0
EocUr4GAeEgpyJ3pUfXo7F8ATGRPY8Sm4qP5/DvQjDgynlbzi7r3kJx+8bwG0FZx
oGBCaYs58csdyedzBF/yfh3YgpJsHfJgJrZDBRSp9MJ7+k0Bdime3l/l6RO8dWNh
23z7UFMAFUwB7jAC9PNQ/wI8cNnTDwAWv/SmQHsTC6uHWIVy9Oy1aT9+6bPRt80/
xRmBm77ePmTkBKULLP7p5oVDYibUTMqALRH0oZDKSAoKITBTK7feoC0o4MDh57MF
KLdEJBMgO23OIUu9wWz0zpTXVY/mD0suA17+4miiIEk175H4O9kCOHm0rjHsupC+
RankRGF21Ea0yVDZqZmscYewMmZO4ocjf3/2q7I/Qo+lXyBeR5xaExi3mzobP8ij
tAGv8YooXuyD9GbumFUfxG33OLvgboiSh+sfUJTtOfnhXOeVvmvBB4zJEyEoB8bR
esBpuNb8mPbFc3IZFZ/w1Awibg1ZFi7dCsL4SBND1M6MpeKPEprHT2COx9edrNEI
4obslJTfnA7VjQrXsib7+nMwNJegY8pXWbWTbpsoO4E=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
OafN+vtFfM7aIELtjS3xbZBb36zZ3sZfQS6hFbHVQHpVPCNbT6Ozv0UD4pJNUAr5
kLjkxkP08NbYlupz4hCSbcF9EiHCe5FlRiq23eg9G8fhyip9Ek7b0aMqYik741lX
FKPWd6yCydArKys2EqByx8ODYJSm/ULYHLOC11I3Wxqe9Zc/RsMu56TfzhhE5LvV
OgqVhr7sExoljqta4sz96KwBexppl/PZ72meORSSOSr9r65sfOppi5GbejBYuv5E
R2nDj6OesdKDPJ1KndpER1gGuU+jnaeM5HIHe4FJtBbALg3zaDmhv2ZuOwnLcE7w
lF5PKetOvRv5hXYgSIxOTQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9232 )
`pragma protect data_block
iwpFNcwrKwX/qBwcW00F3aJIKOKEmSHU9qc3bWezOQMpZpUpfeKU6t75scu3wETB
23PblsyfWWJ7L1x3RLiSy+P3tbXvDrRmavzDEoWq90RVlf7+z5TrVjwyLt0DN+/o
k4oBxk+SkwpiTRy5KJI7/gr4dtWtIEgG2kwMN3B5p6F4AdykSiY3SOMcyj4fBQCj
s5ux9Bcqctv4jp3/TD5YOGHf/c7D/UtathKvWncxl0VAcWcaviVahuNhMiUl+8Qw
rgrHanGIfhZ5I9+P0thI7EZAeNyXYP1guEcYtzZGEhgQMQN6v4KMjzomLbYuEd/n
xvjnBB3zxF5HOXDn6GW1I2FOGrWE98nuaQJ+bSQZnaSBOBoanCnOA3MjLX94ieI6
kEYQDc+0qZkxVJwH2tyu79dxMHo2pBUjeV1QuGNROe+K9Mneg+z1WeLADtZohWMI
eD76+LdqnID8Fo8TeWZ4Pj2dYgQe9KmR8XnL1l9ofEtTMb3fuf/tRNjE3Z2bZiiH
iXySYvTlFAc01dZr1p+0ow2QXa9XzYZiozIp+N3ha/i8oYQ4zfz2Mc5kherNKpmj
KCkhb5xg16QN6VwcDgyV4WKwpPbpTM/6pGd7bZau2in0TY1Gioq5QUCUo+3/lYEU
+GSWg9yDd0ta+uOWsXFvP3Np0dj0rN6IOtVV3ZhAPrZVwy5XdNdMJ+D99M3ODUcx
uE5XhJtGbJHNxmyoPvbKDq+q72CeFeFdmpQ1Hm1+l4S7x2w/tQT3nDDT+pm3zN7I
bkxS84HnqV4hbCQBIlpqXGO5+ViiEeUFXPNheBlPKgKZVBsKV3N0ADviohKqN+hW
FCmohjjhE8tAndm0hTkJcq950CpNTFbzMLwOfABP5SVSgzGtudjGdXVCWtGDWMpd
umoTvFPxVMKwnF3igL2F8uLcq4YRZhiPuc5gl2n1zOh8QgiVAWUSOltxFi7QZHmb
1i+0sAmYmGeDR/hSM9Mx4T2roAEUqsrOhPgbAYkHXjmtJGFkbAoGJiYQm5GgUxVO
OlOP95vFkFtbf9ljuFMUzj/OdjH4zjm36+lFin/H/J1FHEHu7kgb4kdgxo/mwWR+
N5Dic1NvL40BT9pqhvwZpj56pQjNrqFnbsV5OggC4VMvCemG7x1/qWuCkslt51ur
NPz5NDY9Q22CYez/svzIQEAPyGkZ0pVckQx6UHNgpiqmUNbtouYBpAGz5815od/U
ZHz3FsNYisWal6MPXr2uxQmIpaswlkjpUasduJNPo8EuCKcJxsCqU9wtez9cJeEr
vQGipo2mdCap7kueEadLGmdHTEx896PGXeW1gr8OGyvHWUZQt9PdyEXao6fR0gUq
DyUiA/1mvWj3IsmXifjut+vp4yKR3KTDI+a6CfFc99+U4hOamOSyLYWKQwI2vqAU
ymwDxPY2ODBWHyiYPhuaWcOm/Ve0QMzN6XcBMXw2jsd72PPTR1SDIbPm2TYYKTaN
NNCUJAWjgJUUofknOcoG5++wfNd7qzpxK3nAnglLXAH1HFtRPSZsAC/+qsy7KIIb
m+fpvetTdrO7WgD+BDBum3aNQRIKLq/XyvLqceqovXpoXXtPc//Q7hBR2/LMBX0N
LhT1NQe9r88DsTKNWuadVUGCbxEYwDv1+8rg4REsOR5NK9th3Up39N/4GKY4DHpO
ErUcznml7AsfOVjUs2paw9K2t7S19XrQO2eSYVfuEDI02sOzV31FhDr8mo0/LIH8
4x1Iaq2mMeFuQH/zluQnEvyJnvNb23rR2hTfi95fO2n2epwJBj4DARN4K41rk6JS
4V0YdagCSJZr0qQCAJG5Jj6PtClRDXn+Z05CGL8GFSlJOqxyP6bVq4quxi6YyPV0
Hb4dxsQjiIIbyW/dbqmQewxv7+qJrVmZuQStAnTHn96+uX6qXqOO1v8Ws9DIIn0V
VIKRei5tBCf8YyKuseARCeZSdAwntxx7VXDW5hh3+05lN1NyJF8ChT9xmlRDSMAV
NG5CPVJDiiqTbOOFkWF9FDLywlTrm8yKjrd3BUDQB+dwxO9g0plthl8PWFhuNI4z
eUTlmjzhttqKTJyO+m4AdIGvNw7fsADri61crvqasTfXIu+cgog2KFOYFGK6vHNE
8+P9JDFxxm+PyteYK+1WdEfy5Pd34eX53pyWdFCLo7ApslPY3keSyBAh4MT0AMEr
n1CEg6IhItN5duzq+RZkaY14vSr5gkzHymrH5Bb3/TMkSbTXeh0G23PNsGY5o4He
hCjiZAux2yQNcyUjjQPoC6CT9qWQaDWQpnMKC72hVTXJ6uEG50KBgWEEOHx/v2Ac
EDfQw2jRTbp8aGQYO7ndfes8Kl9aUw4XobtRN1SZZ+JJLYwf7zu+n7ZpJSYuWxVz
bSboKC2AYG+JzLXIehpPWvvbbU78CjM69TcLYucbSNoy9na5KEJJE48calVkXMfZ
za4U8voLZEZT+dKljTlfInOgKecnNA68WyLB8Gbz+6nocz7CW/Pp2W1zytT5qye2
GThT3H5aRkVshrxB3WsOsRg1RuCemPLNCE+WnSSBTEEKPrTWFCYKFb57fbXQxCYF
X4x0klcy0rwCWjmvWfAbkkbPko9Lnl5MwlQFhqQWiTcxdWbzpzd+p/PBySqgV8OL
fXlJimrKmBqLogAwi5fYO+CPDCw045EXYEwNwTLH0OMDKffl0bfgpfC9cuBZOfuv
xVQWnelQzkniO1TyWjobmxzTN4/3igWSc2bFTHspLeXYfjmypR7gejw+tvyCv2vL
/01LLGlxzyNjVPw7ul1zYHGKK2ZH4DYe42HG8KF+l4n6SHm+gTzXC74f6jc6crRf
NdZSMjQGj43dd4ajrn+2p2o51VrnfHLEp4WiyThLx8QH+69tSoMoTh3iq2EhWI7z
v1S3REQ2le9vq5dDm0AHOOjEDbk6YKoe17PzSjeJQa1RXbLo/ehEyu4yKK5nSG1e
Ph6iDYsm9Rr5r1ok5Cw5ujGPSnpoqejgiF9HualbbvHu/x5L4Yjzb9dEjVrvuBPo
mGEF7lQpTI8leGswBQa2VnBVHReUyZqSY7IwlGBaLg5Wqekb/iTVyxePxNcV9CJc
O/8JMF2x6Azpa/iI1l1ENgnZ2mw37FbBtchz4gpX5WVMZWmwR/3rBpBN5BOOAG99
oztjcHNUaUKitZsXXaOVU2WgXhf2zpLpY0cDTwcpFb/itBSynnua/OXEtLrZ/SnU
j5FChPEb4Qo1EDgcfHOUkaWwPaUvh+gb/bjCalFTIOpKSsqiskC6pmhfDNPkBWsE
lmBhiFLgGdo+lt6Z+8n6uXJMdn3eIykv6ZvfiuLGXGAGoao2N4GdfcHCOSC6M2s3
QSX2l8qp6b0IOC0Uk0upEu4gdv6SPAUGjB4sw/K6ab0r1PDI5g9B0/2Isu0X0+mM
kP//klEiu3FmhTK22cji11Gl31+Z9KBguqJc56Pr4F6IU+KXGZ1llR1xXsUDTmj9
snXGAHMD382+pJiJKhHTiOTxMihmvcY8pUI0I/TABG5ugraA/npGUqlq12hbMiH2
Wxvo+MSQzHKDTuC59gMmubnROOgM8NSOTYQgML89Grq+CPgaXdXLrmYmDY045TJa
sdY03MRJqJjnZ0W0LQaEE6jplcF5bVSbu0MFYANwyEJi6ZSQEl72UMCew6d7bwLc
6E0M6JQD0DYwZukMVwbTidNp3sstNbSxo0ncv/HXYhGbwdvkKs584QAsnw6F6hqo
IdMsK64gQK/qzrTzmmV2zEyhKQNvsFvp1Mr587oCz+vzYHYTh4yv4Iv2ZcwnW+ci
U4t9iEelT5pEWxr3wlI49bZV3a6onXLtbzmJfjmNnch7WTeJ11KXANMqdNwnfZH3
YYrf0a69QVJRbo7piZlwde8kpe5UL6KhDrXsHYIlqejYHnsnuC30VdberWfoGl3r
mX5U6HCs1f3tN5VOQnbVWBAEBBhpGfCneRlt5OVtOB+f/vwEM9Hs5yy0CuXz7yCe
JzO4vSjo8S2ZxfyseZtufPSXsFdkud0VLpnJCZfQfoZPUKJoRulPseNF1htm8gjb
C+mi1wX9ue3asBP7a8mbWNT5HeXmng2e5YxZ+H1DOpBLrEjWrnu69ujXofMjXhhG
2i5HJYYQTRZh6FcVjuxkkOKh4Q4P1VzBOvYvlDt9i1zFSuC4GDNOmhryVDddaFyE
0aIe256W1BinMNVbUl+MQTcnjHjB/FFyZgsYroBPqgabRmYY00zcCdPCSZyI5PoT
w4gV/fhh9+UTzjAwtGuzjY9xrI9lMbphddY96da/7gwDEol9pc1d654jsv90CWGt
mqywYCoaikqsFhlkEOCznbM6pZbaZYX6zvwYERvLc3JrUNKMneotnNpjASEN4oOa
EYNNBh/mKob9NOh54kyQFyVmKh76ADiYVruK4uj5jlef/MJJc2yqpG3Vx9mZKTjo
895br++ic7E+HQL6oq8MH3iU8oTxNRe1qKFalbguM3aAO1kD1vCqmL76Qtx+jy6C
j00zJB9X42VIt3AiVj7RDK2njZnSz1y46afdq3LBoOBosuJdd/JEIORuS/Fp8OaQ
RSjmHZ/A74GDM1pQaaDNRHXGtMOGE0qb/qV76oUDl0RohQXxwl5XQsDIS9YQWHOH
XqcuUq7AoHm73BCJYEkBCNsBaLiw41dlAUSWRZVr6PRzgmlnZigCFhUo5MSHYxB5
ZtrFiclwQi2kF+wWyWtc9tCpJi056PppCAdTmFey43wIsGl3BxjF7wR3+6L3+wcg
35j9IJbXaT67NO9jbu//H15hu/+deiwbDHjqfw828etBiX3C5+A8jXo6qdYWB3Vr
B+0nL0rzNtTBm0ko18RYk2El/F/YNi5wJRsINkW231t1NlnxDkADXn2F+rO5WJhE
i5bkGWyyWJdbHJeujQv7yq4AWlMBLG8azwgORgOg6upgqui02s4qrUQPfZhPoI3n
TR0QAi/rDv1VStu3S/kHzaYdape4a2PenOjgc1xRRQCS+C9Hm0l5anpE9rkzdfI8
NUUSzRa9WjKbhm2sCy6IJV2IFCRGddMUtg4SJ9hbiA2PZvXKKUW+9twAfNRkIRc/
NBsnfAsgxOydVe57P15Qpvv/2/89sSnHVvzOpmpWE5IZXqdfdhJo5NCY+KUD/KBs
IwK+VYRh2q4QKGQyGLUdh9ZNqSGfytQqOLkhlPapctEw1mLBwtIcdPm8d8jDdDN0
+8D3CvZsA20XXcDQd5wleTz2YKTG36MSsEBdT+VrWTC1X4hDRsPxHd8+/VEGbUKE
XcKo2wfksXzOOlR/vybHDHV82nM2OS7pmrDRIRLykJpDo4vSWttf9NlIYvwGY/wf
VQCNmRlkv/AdJi6XBK3EAsu6eqKg+xsrq2wZECdyYGx2DbQieQPiBW+65EBXJ933
WTLd7W/o7Rhazsf7lThYQpmnpAILF1ubEgMySBr3wPQ5SW3e2DSOSXpBou6QHgeQ
5r10cXZ7km+GFyDC5gFQ2Avq4689o4pBhIrJqsI6uiWDvz6H9mnqs+EH5yFXllSj
Duzj4spInjfu3yB0atnUHft4FQR3RH1baTuNpip2H708AGs1Yx0uS5wokG7HLoJ/
5jgTuecx52CGZG9/vsJhYV8fZXIold3Lpf4PvglXb4n2EW+NeHnQ0vBpe8IJlnQj
D6auh1h/IUpYEDuKTZ0iff5eWLni/S7/Xp5bw4/GVPPMVsqGpDX+EIsT9Y8wlrKt
qUl11kOt+bBFgUw4JBfZHr247eW7Q3Al/2dDUj+9gxl6VeCTuyN4SvEMe9oTshIS
aIdehD86LZfEBhPOy4zsDpwqQ5+40/OZy5d41C5miK1LZQrEsd064ilx53Ubc5rL
XnKfwi3JksV6NyQmYMEpuC9cH2TJtl5KXpUZuFBL89NptRC/yaa7ao24uHhFgiJP
obzOksI9UzHP/jf2wpKgEd7htxtG4i/u2NDZdeD9v7R24zspA96YTTUBdAjs9qqU
a+b5iexFBExdJjqOWgUx7uou/TcWiTsHcOUSaAap26UuBqGioKKzYvm9y73gTr/L
0p+PUqh+gCXZE1HYZDUt5zB3bn7QkrwjYpGe7ufKmBiSNPvitluDOI2KQaT0bJM0
mwEqSf+CLpQpdbssLEzz5Rywu+IzezWWFirH8NQMdfE2YJb4LcbQrdosgrE75997
XOiDbfmtvGmCvxskWWbppUebUJ9hQ1LPQ0Nth2bjoDLbJSYE3OdzbZ3P9FVaUFQZ
y0/rrTdj1qxFZXn3JnkP7H+6+FOrYd/6YWQ84b5AdFYD8jgucCfDf/v4Geeqcc3N
QxF+cX/SUEKapiGxBsX6Cbry0PLBR+rW6hWPR+pQHGCpm5HZZp8AdTUIc03ICVhx
R2zuk0FgzLATnA7W4NNF7RrSrScqv1E8czbHWyvN5BSVGkHHYv+eynrZmBo162hd
R1ok3rdiA/sv217zKY//Grp1ipCw9A54o9ojCYuWPKyuDXDNtr6MGokUWYYm+jC0
/tJkzopN/98aCDjMBt6UzA7t7G+b2kauQVZ5NTNrAgbhmpfqEJ0nFq0SZya7RZTC
y/OOkSV82r77y1qMeNsZspEkmM1gjxuw36DaRn3XmIu5qEBreHnSBgN8WxBy00vp
Myfkfsd6Y0xPx4NKI/6TR+2d78DO6UWex8ygwUeHdP3Y/kl+cRoK11SZHG33fiHA
eup6e9KobeJ3QpdxNK0cOrFWEZrkxTYIBlT2dodSLhaut+1oO//So65Ly2+CWGkN
ck//uHeHDxB48D2tosSmzaLXhLdBiOQA8oIeG8bjI0DfLsOeUt8TYpi+YXcIJAGZ
SPQE3FkU9ZcQeJg3mBz6Vx7h/C/ir0gRU0H7+fn3R3lTdslyoz+xnOlKgjt0ISoE
cve4iwz7rJCUpTaIi+CBhu3CZWt/h2QaSov0aitnzGMxVnA6eXpxYjiL4hHJ46PQ
ub0KkRZoskKtGxgcLT7KgUQRSlxOHZq7LmafklMJsfANthAtofUrxIla1i2x0ins
ByT5z7rX9Yhf2HkowFQ/C/uvbPi3qQwJP9TmBSILzYPnt8OsC3tjo7rv6wadHYUE
8YzZd0BwSeiHdeSnNL2HO6nfZHPO/U2V4A0nC9yZKa8q3QiSWytvbh2R7WZq+G0k
RZZBO0P4R/BjS/x/5Sz8Y/+cZXWySdKj2eRRM3ut9jEKXtz12dsSRTtf3YXp69PG
DzDwBfPa069IPSEstJBncy5xTyfbrSZG2rvomhBxJZc+mS3TdLcEumIryB2kcEw7
f9FipTevuL3KmtK7wgpSTmKTlG9hMKH+GH+c+sHXBNGIPJprd2MoaZdriPu6Jj76
eHkJn+hUl3DYrA+ZQ2xJn6wpTtyMEM5R8hLn01/uAD9ks/wrWuvmXTMfmLR9P2UI
Kpp/f4Ve+4CQMG/Flgmoa27Tp1I8QqvPs5kuFauft2RCBGQ62WETqdvgFcnCdQE9
dvYcgWaynK4fYEeb73GtUFUXa8GTzN/azofRxYaZqqFtdIOUJF4FMlak2jd7CkR+
dd2pyvJL6gC1vTAqFOSmCjbshzWMFcreHK7G0B995Mm/lZzr7dlK6JVK0gwA7PZe
lcJcavGi+nWolzZYvJIXbVmJ9M4hfx/51+NMrQNZTYgO3+QrJA6aXI9++RrG43N/
qvr7TQ6zp9opgIf3pGojZu0r+t1uLvaSSffKpDvaWxWCxQQ5a5ALeD3NiebkTsea
YQfe5YF/LCjdROWfAcR8TYjseSghvGqWBtJfWeqfIOFQKPPwitJHoEEnrtqPJ9vC
KanIj0Yb3UMkW9+PUj7A1PDpAmeXHDsMzi0XFOjcUI+XoHDcEhrHaoafQ13yUY6n
6E20oDkCKVfK5nmTkaHBbAVTZ/4uwjyB7nBboMqzxpDnqHYDNzWVLxnrX0CBBVYX
4U/vIryXaIVYBG2O7Vyo1tQIVgKIII1duVM6y1ShziSIKadB84u1DO7DPAtcwp4L
YWCWOoMsrGUDfpA7L/h4aU1KKld9rOdGScobNgqlgfO+H/5IpMj+BcZNghsWZaRW
cNagi+I0P+KcNg8Fm7q69vM4geYLHdQF+ubr4e00wLvO2qWnt62bVdquhNlnqBv6
fvSi76ttL0qSR0KQpp3HwNoiXe/eZQmmn1pTqGw8Cy+V515bK7ccJokiRVNZHveX
YjTB1+oGFzlcumIVLO055HVoyM7BP5+SrgC3ywg20q4H5bMtC5tFfL0gEWwFFzXR
w1eEVJk0DJXL4XT8HRROkk9KGGFmbgTwLHVC0t1REeBSm3x8zwqFYgigCqp55DrE
wJGN+rG3bqLweVymkThYK2VjUE28Oh3AGFX2QX22Ey5JH49AKOqyua+oM2q+DbMq
Gkl+hEAPC0VihMw99TzVIFy6nyUTtHmlZ+T5iHhtlm/nHP5y0cmLDUkkmtdwdAat
t0X3aaSnSgw+3GqmDlIy0m94Ps0cILGs6a0esjTtkeVtgbH3aAU8I6EGT2gEVIhF
kFpI8Pn9Z7ImrT6ZdypN8AkMssEw5222PlN3LI+OXjiBNEBQ/wbx8FYlhPqpQMcD
M0SOzrpPgNtSmxHSK7OQ3zuG30HcKUupgzdMToqFyGFzRRlN0KBzw0O7xptHxt8C
KisnaboXZ5YhEPVT5DT++WevuVCJV5j4dhqxGPMJEvo2Ud5cux0pMJ3tvs7gFMVW
uR4gYaidAk920a8RnlRNMMpsK4QcBbEJOPPeuN2vI5WIIlLBZkyZkZ+QXpX7vkgC
G4HYmCCU38lOAi1mzFPfh7EeYv+jqi12yw4siGgNUOIUDQmOUJ59Hg9uKCdYAhxV
VMaXDnmiZL9pqrPqCzo6ldxWZ/XJcZDSmmZmVQo1NqLfsVlUciIPoCTkIg+gkF6O
a2HxKZEUFCJ2RA0wxe+ba1LiqL6vQSnbQdy6Qq3Oo6kfB0GZ7wah0ZoyBIULSrTS
DCDE0tIPr+SNi4BHjJ+LlP3/0MesnUw8L6iBPLlLg4Q+rSrC5mZHeOdjIxJQzCQR
2RALwALym8ey19ri6Eng5SnOJln4qGmlOs/8hIjPeU0sXGeCnQZSmdcJ5ojiF1bQ
0o2fmBkaztyidxkdOmdKymt9UIHCqxFLhrLKMe/mJGWV7bHMuoCXeZ0kO8QP1XbG
Qol7tCTyVBMb3SW6yjhDujdZzBImiRkCpipHUZ0NPsTM/lyTA8p9aI2FPEjngiG6
Dhab0N8LPop1sJkDCaRvu/ZSPE5Mm8sZEOS7pZAt9nZcIFWZxQh6665UxwS40BQQ
3ZW+J811kAAU9ROmjz4J3iNLkQnmkVAyxiNCr3qu9e/dB7Byll4Pt3GrYzhh74Ha
zj7I44zpdjMEbQNIM+Hm0w93VH0hB0qzGHzndw+1plgJgIr5mDgBcrRLBSQThHOb
UYlCESCS3xjYT320WgUc+HmZZiZWj90gbU+YLHad8OhhdQj8M4Wobr0FscdifWhj
j7mtrZPrTqvjKLPSx3mK5dA+JmtlVu5xVMXmZrFwLs2PR4plwnHIKszwBvCq6fXE
7ApMU0lTizW4qXol4cc60Cswd+8WEuxdPxbby9TPyN6LMSFvz0IgZTEYbKRpFd0k
6iPGkG6ERp1OzYpkhxMTvHOVT1psGzuMggmL6T5gp3XFiH57pzku1G9eRIIpMALA
rS7GK0MsOcu0sZRFeeI87qmFD5090iYNAjPnjhMlDXm8Pq0vvFj/0w1M5xp/QvjS
nWCF4RSLHXp4uPX6AugG2mKhxzQ5S2jEGgmIzhmTG+pPpbppkVW472RkFGS1YqQ4
c05LJKAix8nr4QfzFAFdbKAFEBX359vZsLNZaPTelxvbQQ/z3NBQ8MFXH+IGDsyF
m0F47wUgEYUNSK1EsRcKEcdkiTV4bpLlwx1NVN32rTaPsxLyQnMj3LtfRXhZKkWt
C7KNUikQsHp3B4be4Y9T+joVfx6QPF6eWrBY9y/nyZnU4w2e6NdrEUxoeT+OpFaU
hdUp+8BJwCdg6t0Eu/42+TMuFGcXoYSQ+fqU7pI+ZKBFcDYZ6dsvGWg1fvB1MB5u
FmEoFUzLtY6uEI8Ks7YfFg06JObOmP6mRkSAKo4x/aQRp3Xd+xM300GrUg4OpErY
0qHOsWbbrFL8wnyJQnR4j7AhM6KAdjjogFj0wkpJLoVOSVFyMFDoVtszdengZ4U9
UNIYrdDSfwU7KUPYY5JQO1yiNKYnOumZg4ZUfcrwdVOHxyrZMMRlrbmgdEwm1qgO
87/72ly88umWE2UveOTbxMdhR7CKpDEGnt6ahHF9h2v6nI7sRAwm4R/ffZqDH6yr
1dWGXpnB+KwdFSLgO4S/LHXjdF1tFm8KGQrYEiYrjFRBzycg8ZFwXGhug/j6Pvap
IE3Mj8Z64VzF6nTtITMs0/ACvZy3JpUTKWstROFXzKfUNybTIFhsQcE1xif5WJzx
Lza0cryR4bWNYJG2t8p9CGUVT4b7yhB3uFx8yD+498P7MG5Yy+LPGLWUtR+GjR+d
8FVKJp99v1fUpBgpdKphyAfOBi8ExelgFVNy3rWXNzKugzYcosa0lScsi1xxEG67
yRNP7ADsd/Ssp6n3IcWG8sjmaZBweTV5dFydHqi2O/pWYbsaFURNxFhjkpBgWU+W
CuTQ4kcsaT+77A9+dkcBxt9H9IUJM21A5h8m8WGQNyiN6B33xKDpz9LNd7tyR8Zk
t6I8jIIikDr+mGw7MlIYLMQrac7MbaTvmCKIOxvKTw3zPuWIHJqqPTXogED1fIos
xSOUNohDtP08yYfMnyiZwf7yE3JrGeJZhhByU+Fr48j13UnKOFxvF0GEj28VgohK
eXGa/GxL9fw3R9tMxzyxtP/VBSwSwbL8yMk7Nugn++gioUA68kbBd4aKQ/+69JCa
Inb1sc8W9BK9bq/jVCyHx8OvP+4DZr1gUH3NPfLBk7C8Dx2DEPZkns57w2MZayNz
DdDjUxtOJsgCfll0lOhcpPJZBqFclIxbBit+c0zwO2DdAuduVpGvj04ACcQNgG+0
YP4NEoBqvQM2OxRbAb+CGZaQMZ8D8QArjU5fYGULKiJ1vL5/Rah+BXMd1uUuaGWT
1jQ7M5amlKX3DiXbFihBS6PK4ft5nx6PirJu9n6KGcFbm8R3p8lUevyyMdQqQEoh
fs0LSfahXDEKPQqABV81fM+Mnmjr+Gs7tErqPci4r/rbD0fsZawTOwuoDIiTIhQv
S86WyYN046yAev/uJim/rBFY4wsejAR/2pLSNPmqtdNI/QONWM8cudqP8i1WkZso
t4lABzZcFM+TeTTAhbO72zys2sNnmrpl+5nAnxa3k3ac0MCgK4ktzoM4+c+iyP9b
Gec00F3T3JQdv3RrxuQdBVOBPDJRkZuQcld4B+BLyEd6SDJvOnUdYNoWRUunsPir
LoQee2P56MWZQJe3uUWIxEpttP0geA5TnTpv0X4T72JxD8xWD3cWmlOoNfBURGDn
mLG/ona+/5jG8uzVPMpLYBNW5aiuLdGijXn1WMcXux2OCMnRQNhPywC+UA3rZL0j
gMW+39JN3R8brkad5GrlNqmq6HyA6ZewyildcMMT0N+rxiNSh9cHULwZPlWFX8+j
ESzp+mQHkZMJf+cYih85xA3SLC8oLwZ2p1iOHD/rv/XX0CW98K+8vOhrshI35K5j
2eIVB4V89rIzi5qYIQO1I/Gk6YepA7G71L1HtQ28T2LD6BPzvGFBLbamKurkFP6E
5IZAxkoTT8RBrOu7T7l6NMKJfT6GAfcG1NIhO8d2oLFULWvj168kiht9pqdSQkr7
AhR1l3a5e/PMxqhaVu8IFG92LYi+wbqkdwxRT5hrpTfWm/BdtBdNJOx2g1rbOb6h
ngXJTZBAO4b+sjn/LsO2CsGam3iYAK38w7VCNpk4u1JxAi+0uqfHEaAfCr8i5Q1y
aWZAft7ZBygGNiZ6z6AsavmUm/6+CCeLDBjSdakls4ieOkPqJZXLTt6z0j/x9Xyd
0pmhvI7XCHfVMlFloo/LKh5YzT7UsuXOHuF8vfZN/WjmyEKTsdEaZshzhCLpu4Rs
4dIZ/jg8zrzKcWAi+6gmVe2u/CjmGU9YCLjv3GuOwAFMYidwVtv/ptw+beS2vG0b
7y/SU9FARHFF/Y6WK52CZvgR4ajYSMC8kiPsY9/YiPs+YcIzUn+c1gJT1zb0KRur
CR3qiP0nM3MRyoRmaEAYPqRh845ShUpLIVsh+pXaSfTZQHl2CMJXS0Moe3f7vRHe
QKOV0Ycf79e+ruToFRDiloxGLUEzqxIkn6HSXtEdQ+SL2pob6tO0z27fW4gprvDQ
fS75rGrPZ4qWTg1iyxEhKvN6gYUZhXGr+URlTSra3gqPn0PUVws1qfLqWErbPtSo
j8hXwn2+iSqPEewk4T+znw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
mmOarmrnz2F3Z2HBT83pvg0DDZ05cufpPo2tROvEfvDJq4AlugWm2sdQFko9ll+X
whChLDOvHXjUkf5yDbejckbw4agqN4txc9YZbPB8fZJJxbE33IatVJHiK2JXUoJh
n6w8LayzOQaeUsdyp/JmLAVPfis91DSvxsI7YHlfM6vHLclwOsbz8voibJyYyn2H
euzeeVWf8E4DRGG8UJ2ab0GsOSk+R+CSiK3ge0uzA7xO2pSXIIwMFijhi4NBCU+Q
mc6Wk30mArnhiLkbXGXOoN+LNleHgVI/asbQPXqlzd4yhwcWtQmttFrJFmx3G7Q9
5nqIndFHbJNfrk9iE3bEDA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15408 )
`pragma protect data_block
UXpHECDTTXSlAYyMwpBpBtSlfq6v9kjasX4CV3E03gAddnZsV0q6moEpQZ7Swi+k
MWFx9eDN4k6e0+8VHdqXWBNtGXdt5Qa+q18VJtHaOefU1QHT7BusGcLSI/QVd2IT
u6cuInbXvZqVPWcYnTAHI18L/VGxbIaiPJlL8TDpXYF4g0RWm3pPEEMm5YZyeloK
+Kfnspnkn+GfD67gYO0hFHrJD6bZt6J/t3WSjGW2VMG3n+zsNrM3rvcWIjlY40CJ
7Sc3b7zuMIbPK1KqOemaQP3hPNP7FTX/bFc5NMVCZ6eT8lp4HQu7xMEobRtB735R
nQ3k9OlcUPg5d72kCypO7hyoQoD+AWAsYFFbs0oooIk7XqDmEpV0q9lNEP5GUW9E
yi0yD/Wg3LLwuL0yCPpPIlZkz1qk7eGraztQcdr20okC0py1tecyY535rnPRAaIP
rgxo+N687ekvBAimBLZSmB0Y/OlQmbhCzXds9E5Sl/DtkGztSBwoZNcM30uqn+1q
nwvXwSF5y8gFq+1iWk+2qOQa1hp3VIz6dGVt9FNfAvw/N4CcW8nFqABcTu5q5w6m
LRW0PDDpXhuZ5XtPCOwqPw2eH49oEfrX46Jzy+rr18enOeo23DpWC5h31HBpSxXI
zrmwVhrBfyoc4M0h2ZLwW/ugD36XQZbwZ7HysFQYHqxW1xzRkv0GbW/yx75MHPJi
/SoipJ87q1iQ/7R3kp7rllg665ZOUfPo5hRLxAgatVfFvWEA0ZANBD9JDVgG3NSW
QCCKJ47t2zD6NSUHRC69egeTR55FBUp9rQkRC2P8FTPCTOOoRLUUfHJCj1+7aQNO
+kzr1cclKeCaRx50bS/9cxJmJzFcy+MIbXUvfHZZvJzkC+alPiAXiPi3k2cWA82M
klGZgtB8Lm7aRNFAM3jG0bZzPHtFQcuKVnyDZgUFbhp6Gjn7lC0BAFW4P01ucAan
uq25P69h24EEGKAHvgdZuRxELWY/JHcK+SHI34zjr5KR4SHXXYLBmGbUoKzsfgYz
/mNE1ezYmDPjUmdptFzRAgq8JtJYMK/ECoGGfCWCe9PIgFuOURexrIFW6UMKg01k
03o3UigM3cpVo+bDgFqme3dFkS3GVDoEW2QWFaiLQaHbQE8cs5llFlDJQZw4lIJh
UvFw9b2VSHzuoIkR9QsHwX4hkwAj24cLU+E4bVV9fFQ6+psnxxzM6cfNUZsfJtNw
fOz1LAbbxeezNN3ZCHdF+bfvFR1TBEF6PlLQn5ecz3S9n8xicAFtYnKm7WVEvFfS
6odxrxTStSRuN7MPEJEW46M2wEXSx5Ze5skQMc4R8Fds8B8WbCjQS5XXdyfLxDwS
PdE+vwVtfEgkJnxodKM9Px1ogK7tFWcT2dBnsRhpMDzxNABzGnwqXvkpNTj2MdOK
sEHASel9RTtr2/hikbvxdoRofkhtGtUxucm5GHECMiqomXN70qIAPZ214snPqldc
ehJsZTRTEGF55jzKSbAbT1thwAqcg+RukKjBsI3OPk9h0OeoKQEsQ12S8HVD+uYM
tn5wSHVwNqXIrX7T6eScDORCtFoKvN+8U3W0ExrJTZB5YMQjOwigjN2LgjyW/ufs
C/1SJ0VVUhsk7ex75OBEqw56pSYO8fvbWJbo0kxWUGRE2uRiQvziiQJd+qe6Oq0D
TC5uKJD4VDlLB4i5Vro0sCxIARI6rrzg8thF3raM84kS0r2ow8t3gNhXCBHK+J2C
VmrfyNUVKsJQkKgo2MByIOCD7siYI1C1lVIwC7olwxEZgwQVTqVL3HawNKpK/H1F
Bst49jArM8ijGxifQVjfqqIzZnByvyORvlpuAMHeILDE3sIodJZ6xQeIBC+GK2pT
XpYL0nOd16ekCNzc3I60tdIdhFGyXtUsH1BqSTaErZTTHBxEzr001jdkQeCMNr66
Gfm9BCaGis2IioTWehlLK0EDk/l8+Svk48cDfGesToj1pl55eg4V983G/h5F5IIg
7vxJEcRby+cNCL4twPSBEZCCnw221DinpAVHZsyHeiyfkgHWn1NIQ8O8L7GQM4J6
gdh7LBqsyzjN3IIp93P1E0IR9tToH4LFAYhnksnScsfFMF5iIy6Mn8sejdo2ppW7
TcBwByKd/BGzep50UBYBspEKqskNEypnJJEr1Lq27hwShLOBKgyrurhNqc/gA8GS
+j0bcAO+bq3drMzziqmpkCH3OgMOqUq1GWKYMc7BTTGrdlxBzudHWEIZ4QiSy+8n
vtWVxeM88Xp6qek58uvmuteJdlPi3JZra3OmTS2MjHzkYxzNizwPx1dojD1Pvsla
8M4l0sZM83x5shWxOJlR0Z1qp/EZINrdGiizjAMYlNrDYkwBvreb9prT+F7yJKku
T0oLhveqfhDwftK6+J2q6pyenalJUpudp2alc7Z3VevqFmlp9S8Dl5prDck9F4fb
lwbnr1qQue5ayj3e6rO932ih6SxW9bOw1GxjgJRO70KcC+aNDemYpr8GKe8YJZ/t
tu+NhUxmix5NmpWnVZzHrpikX7dDcCB5dq/EHToxG4jXM6aT2Z0J6p+3iAguUVNE
l680tu0NwZGk5Jo/2U8835knVl+kwsx92EgcvGidKOD6w+8I25zHiNkwmvK+j64y
8cw5+lyESldQMddFzjM8uPG9nv8ahN2OJcHyED/VvxPvLtCmCuZXdJNqRKQYom+E
4TII6sXz9XFvqFpIkJ84wrh7ROLpmXBzFEVaOd8Pz47Lwty5WJv4v1Zy0oa11SMr
UKLr2tqo8cLQjK3V8/jickNlfjQ+w5kpdCuTmNyioJO0UD4gbeHFpMT8MNOTx1bN
nEOor5FjaBPUTXkDzW2yIzl2R3Vwug/PBupjBKRNJ5x0suyDC+TlDGlKcEncdEb/
pFW7qEqwB0hdMidko1lbS4+wEgC68wqgMUsNUMk0mk1/P8YtQazHbTJ13yGczW/V
1T+WEHGpmeWeRhcluvNu1uZu4mAr5k+fS08VWiWa0MzrRfaFBtyE8b5xYbr1pYIv
yRncgHSZeLHmImMDfDdOFfN7lQdzNuYKPzsx30vTKjOCVNVQrRKbwoV/BnQjmhvi
d6ahC2udsLixgeR3eo2qyB/cnIwZB9kZqB1wCQCw2lDfit1LKzxST/08fm0KERNY
FJPnWb9bb01bBJwdd3CYAKtWVkGsfkDKLhL4suD9cH3mDyuUmP1yzZQZH6Mlc5og
K86nH9lckI0exljaDoXo4dCZ9AqvXwBHrdSnTVn6dOX0f/uFkTYgccuR2WvG8Trk
GFmB28Uy74Rvg1i2l+v3KjQuwcoNZpTcZHA18/cuMQmI6imb2LLQ1uvuHDgkCN4/
lpmwwPCjMh1pLclDtIJzouDjpRK2FL1U1bb1DwRPFd8QVKa6H0IQyHOfJeg55f/Q
de1Hv1mpoawlyAweRXe+77MwipFwouzQdfSu/Ub+FUH4AJFROfmanS/DovfnqFQS
2v7c44dmsKtZ/6/Se7XPuNjesL3ucA8/cm79/rFzP0z4ZqfcQLiukhPXY3Ngi60B
e4WPEymfH857N+WLjWxvipj6HkEE4iTzVdOwF/WonxyFdqUtC9L8BGFSF9MkrTBL
DuwP88f2hh7fjv7f47tQvZm400II2f4Bp8IY7ajAXIh3O9+pVNC93UWQuaJSpgEs
8u+O7VWUbpo+Wga9+Y4Dt+sxw9QQadXm9o8zqL+5al5TYKeJrSHnH5JxXZY5CV7/
mWsCR3T9XjzTffwiJc6Zr0qN0Z91ZGYffUXJ18qeO5Yd0TqnYyT9lnwdA/2E84v/
eZP+YTngg0diBLaDvHveX0wuo5lUJqY00oGfiVHlsvUVIfh9CFp7fGBmmyrGQc1K
/0zStQBSrKjt3NDzdhk5touWZeX98X4ZsdQXTbho3AyqmpnLrxQURoSmSrk3y+Lh
iQZZzwyO8ZK3FqjjetfnLAqBoAOaaujzak8qzbJmhjEFZBb/tpl57B0Ej0TFuYcv
K49C0mcgr2poMlygBVMfX+Tuj9rOcjww5beJVrkb145joq4OUKcmPZGjjR98f9ov
GKg7n7VADlITGAfV2ublJN8sF8W54/bz9fikvHQC9iKrMKdL96vottzu5Xj21DVD
owLu0VrfQBA+v2deCAOBNmGCngkdeskeJEVYZK9zcTJykDwKn2e1ce1hbc6A68XI
T/ZFRuFKI6h1XE7n1aCswMyeKD5RyIVD39E+QEyZjaTu1+GYMawH4Wfpn6wf50zX
oiUOH2UDGbDdwVH4i5UJd7bgjIFHBitbHAhC87VpvuGU5L/hc2J3eFmDUmTpKPGs
HDBIRyoiwPyPas0S+rPbl+F58NW93az+hbocz6Fh1M7p8RRYQydItUqUn5QmpXGX
gIpJoW0+L7tNts0BYSLDY379RAtTsma+nOHgrh8cHoXrk22WTzYUY7UO0ON6iivz
HOCz77RPBY8BetRQUdswzUE3yEZAKaEyZno84LVL7S9BKz/IpPHPPDU0zoyaq0Of
Ennhe8hj3rc8wb8MrCP2JMq0mwlKD5J1aYzAkcgXufxoUbi/Ly+uNjrl/qC2Ttq1
9Or/STciA6Kuh7lSci9mYmRcSGHDFwMJGbyenNjMAAiNxaifUYIZ9CvNMtz3cJ4U
60XnFeGYu9E907SXlPeVBOrVaKkG4vrEJbAclYQudT45TFbcoPsK+O6tadmwUmcK
1zc8sNG6CFhNfuYWk4nWTVmZxR9DnR5Wr3OH8CozYZQ+R/C5GcdwL7R7ljfrfMiO
Zqu+DdF+v3N4YQJeZ7SsxMNxte0lC2gQntrr1jOn4QRQhKVw/ozEo/JkkEo3ag/q
caorcaec2PFCZLNJNo0y0zcpeYVaUfRewvLpdprn8d9k3UIfumlYEbXjHsnnc1yf
NgF3Dv23GvqEspt3efYbsRosFOYiR5I9ALQ9ARrBWb0whqa8A3moK7wRycH1rps3
IHQSC9/+jN5uTsA8LQmLaGB1cFVWDvyled/w466rX+ji3B4yI1AqtHQnskHv5RNz
Yls+cxsr7ls7sIFbWUjg2C2GUznHe7a5eSzx9ZcfxIt/WnBszHP82+IhG+Uj5mg6
TwpiZMwPDdph4V7Ljq9tyGPgKcbMIGdCir7XQpCNJlgAmJwX2v2pDs5cdYfonbqB
HVP4W83k6rDApH/j8dLxyLlafEfAP2Ks8jTGCJ6Uy1BUcpLzaFDNfa4pi2ohz3lf
VzAPk/EtCyEyeR4Pv5WUyzPf+BXS8SHKjmWNhGV1rvSLcN3eY+9d8JJ91BkzlUsw
bE2FYUDxxlSIz0iTMzx+fxYdSyjK50UDiV6aB5eINKFz1t3YbilRQa/HF1FQY8FK
LYUaKpzisH7ykG9Rr3wAdBcH7UYCgpU9Ssvf8mwLZE8WqbXfUoKsvaEB8dmJmLck
fui7BapkK+Ty7Wx8pdJi17YRdQzml+0YFfcqNVf573aEukVboN0SfzbOReyBWXuc
CpzWrqxgrzuo0ordLe+b8rGqlVProhJOqTV03wzb+WdM9TXedSxwZKQMaArp3LPU
wkpag7A8S+4WB6+sgFxYCxL3f13M0NupWfrigPslZtj28mxHoW1eu5dfxkteOcSu
3cpquQnkHe4H2jIbdjom2tjoMN9wYYyxcjp4ucS4pE4SCevWsEASCiscPi0cIRWZ
u4UgrbXAED3m8eZ6yWwHaeark2XD66V3bmUjS+P/KqZG4pq2+Yww0ITkl7Iohp97
7QdrkSxxmNcc6qF0guCLZUzjsAEvwYORv5lGe2HVwOPc+YuDJ3zYwlibwkJCJYxk
yVI4h63pia+CWt8B20J2p/bx4xXQm1axO/5kJcWOaZgggMxHHnbvWxSfftGkK+n1
IlmE53n7MVLCWFajwOY6yNzr9PaVI/jefNWQtVICqczSWN5OwpU7kk+0j+xoROCn
ETROHl1UFBcFsjBQwCsagiUSoYyQZtu9Ey7+pSbYllZzwJ4dWdcxo1GiwgyXB/D9
OtSgA4PfWKn7dF89VgNISRHm6vMqi3lt6mquYpO/MKnojmc9Y1JdyxfX1vBICa8t
Qb7mfgsKydofz6H5ThT3zoO+05nzMCuSEZPrekP/YPhraMKcJ5KxE54Fvza6R2aj
f1j3Qp1FITG5qUEvnAEQDVJ4553n7xChSLJG2Q797odOWiNpEK5dYHCwh4lI7ohx
/PJVenNxroq7mU2fUVVGbdKYKQif3xlQBnVF0jbeUoRVvTojSRpOII1Gc4Howr3Z
DxdVr0HDBK/uufSycSlk0mQJQtywjg4RcAM0GRHawDE6gfL+CFq4gvTnJR4ctuzl
yImPkx2x+AeQ+fSyeXBtTJHILlUzZ2PHBe231wyg16Opd4Vl3Pm9fcNZxfANM5oj
ROvDjPSwx025LLZGhtHX8eFIXRtaCEuUlj/JhfUWyuL64X5k3dz/AgEBC0iiMNyF
FH6ESOyi/77hz7vdrsm7UpHeWhVZKcGAX47j8yPc0fN4ANIHThlzAlRi8muSrS+7
HCz6Ozp4+OdeWK0OGF2ZCWBARJUKh05nJuVAF7y5L9JrzhEnduavhtLf2S4cVjA1
Zgblje1QLShTPvY3JUSRHaPpVh5L1aL3SCPB5xoHWGK3LBemz9iTF2XfOcY63tD5
rYcsYUisbsIAb4C6ONmHCqzI+lQSzB57aM9go0fZfJwUBVv94O+RH8wCwd5hA25I
S15sza8QMy9BD+SE8Zjp5TvGOkDRA+yG4ja5bxS5HAE4St3XQL0GnbcJqoco0W7g
mb6tF97BwVXBFLbTfQyf9xzDHKyjH5eWG1kkGahcU3wO7g8kNDSsPp++Nl+DcYoV
DmIeASSNX/LTGxGJbnoZFSXFbaP7YEAPMeYlIkHbg6tGeaNYCfbrXiQs5ovvrKdN
HLikIJ19zh9FeFeoD+N6OoQt+ugIpSEujd1/+BOppNb+X++dsDtzfLC2nJQiS3le
MewnygyTu2GB60N0JMQ5KOcJbNSHqm2wROcwALperHcaYZUJZX3PQjbJMICYxijZ
ux5Wtn29N4squjQW84YEcfl3Vj36y8zJqWOIi/0d1s478qdALBjZt/HgjKmksDbs
Wt2Jfu/eCH3JI2BIXg67ooLB/8pl+ap9YQ5l6CIZhx7JFklrqL8PBtzluBy81Ibc
wrBzqZ4B29OCJg/DNrBT+Hif0UFGEHEBrnl8zvNRDX8XlXOkjfTp6dJ+gJOrnWxb
Afl599XaSbtzGDxDCrCOaU9lbLK+m/MBrHEUVta6Dgn1W4mh6LRIz4qzrJ4a5Qe2
dcv0YISxqsgqJYcJ4f/QNJOW2nAWidklzD00KY0VqO/mCh2E8OL2beZ6l+AypkYv
2Fnt1FSKo0sKN8dJnvr0em4LKZ5gZbSYmyjxs9lJQpk6WYidrPUzvqASR4HWkP/D
bAOKb9RjP8XTDGsuBn4LzW9jF+cFaAt8igLOP7R4Qis7OoafXW/uT7XwbSfF4+/R
HBMxLzx7LHgqyMnpc2X34UjoLR9Q7iL3ERI4jfO3jDBmPmnifP80S9GFWhJfm2Gi
a0VVATLVIzcs3BEUTTI+xmYdP4SHxblaFOSZDjEYUt79trHLeT4mbNXqa8MjjJeV
eGdAgnJvoGDJg3G+6EO2dwTkHVyg4IabCGrvfMNsaZW0+TByRSRvXq2irLjfrpQe
CXRPVowXEVyffIfIrDI2gFZAYTALGI7swjJAzoy/wHP2UvnsLA3ICLh1B1DniOju
6n9RcDCfwWtZDrgMYnwIMNacv0yt+OOuTjStPKuNcLO+QpmKUdTfuMyFViUlLg/p
R8s+pNh6GFV8m96Ld79NtEmUh3+uEjY2A/6RugNOSAalfO/lQssuU7qyI1eSMKiN
cFcZ0SkzQbJVgw6spvghX7MkXN1kF4SsOFMY7R08b9lqaGutibIIhsa3efnsj9yU
n0xh/DfXLXnCbypwpBNJigkeeux/1awfEAhaxEkgeUDvBJKF7J9W9O1PQAyZzygn
KYAd737ArM7iUeXQdc780NkVbeefWBiQWFMIpOHOYpkEjoYKzttRCdWV8OQL/y3m
wHlOwYNk6HX02jPbqID4StzcS3rFce2sp6vZ0J/ina84URDS5IIM+V35BCqq8kt4
a6EZzWMMA/fzc0xwITYcy7AlEnRNiVTK0srOMlY8W8SK3tDePgwYdMrs/AFvkM26
uK4PCVdLluFklKUX5MqJghXmEol3tbqAuaLkOHUerZprC3G7fV9+RuSlWQjEJh9A
TT/1layVkEE4dDdc8kfLM2nr9k+K16IdtAIe82H3Nus7FRKvY6mtx92Xz2fvUyTU
GO+ZDmYpP81eHlcVhD8vG8DozWDOiMEcVhYFJocN/h7N4W3EfK8uXOXRJB6vplAg
UQTQuoycBdtLc312LI/d4ziLKpwr4TkNfp2XTvxhXs5YssCLul9m9ujQtJFXUjiB
fECNHugXO4Krkah4fZB+p/cHDQg+NMRtXz5b7anfL11zdzJJL6WUkEjbKg4r+x71
LkoXVHXi5oFHYrzdPrn8i4nA2vTHxu1h5KIjU0lD6z9yxqAlOT0y+O+1XS7+D6Za
/7J+f3LppfeKugeveklPapc+rUOpXkl6b36mzBkjGold4yIgMqKeeBRazuzyF2sW
Tqu4lg89v9fezIL5KxSht7JRLUBsq3Q8hYxtE7TJEFikjWgKeGWVbKwavvtYPJEg
PSkLpGs59ji+PuCEli2OTDM4k/T8iqIapB/CD/MzbybnRHV4fZ2i/X98j8wMC0qI
1untf3IhartW2YdNwRmd1FJE0IBnNyg3vqLoJ6C1tNDnDIwkjBOvnq9WvWKM/WpQ
oXP+Fv3y88xXeD14g8yWSiP9hG9pYPFhuFaa8GSBJz92AMh3PdqZAXS4vykY+TKe
AH7NFvR6s3PyKIzSCo0NH29vbYoaqTPdZZa1kPi/hSyZroNnm8Pe+7BGUzAmXJBY
rHb4JJd4k/ynzeEWsDVOCWYq1XkvGQVnYyU17imbzGcS6eio+D03CSmcrfQ3o8jA
Nqm+QBcnQPNXH1Sl6WBcPpU0sO8GYhlVloS+9HIEId9Lfx8wBwCr+RMqaKpdakPy
qUxjRej+O40yaEa+d7fgx3WQRCAoxeyOaN+S6TOw2pQgH2Uy5m5Ixl0Lwya4XRlR
IK02oM++abqHYcMlxCnJdq26PpIn8FFnM3PCIcN6IhvJ+F18u1A2PhRWaSOEbiCF
fjN4UnKMgrS5ggMrEEj7oqm97YniSdGtQG1kwWIFHe4NpDfihYp/dczG9ao2iMQL
jtGPir4OjsUoqzCxFM45qeYOW2qHWdhSN3SGWlM7BUm34rIQcQO4E79DCw4V1KPp
w1tRpm1+D7UfTWNftD1pVsz29hXNa5j+TRYWckeXduqiQ0WQtRY+Bt/ZfOcxlxGp
6gmiHhkwNb70rnYuK86P5ti6oEhSTeZVaMaeCq8w6fkushGt0UiiQ64bAj62CRXC
G1OhNA4sbgYUtNkDYvG3DKY56ERdBsqHd/WleW8MFb1nkkPyG4Xxaovebcnvkh9t
y+6+ZFJ6SljwYC5rncamHGqxjVV53xVAB8wXu/QZ3iotX0QhDUX90luLjELLLFJJ
n78up2QipMHPElBF3dFBhEA5rXy8OR1+yWBZXUR0U+qd6nB0GDA1U9NwLUMcYxuQ
t6Hgf7JkdVdCaWbAzunJmc8B/mrHqOPqXtsJQdZbfqIUEcumCHsVI0Rzlt7JbXdn
WDe7ILXGN6kdNQameLQOLw4StC/8tX51cl9FhfVlsdpUHtLojjCHV5EuAyRfmB3r
7dBG0wKy98Rwc6J6Ud2hIDduUIrkkMuou0IVcMdS+c8ZLsgWKuw/iSSr3Mo6qEUK
ahhOaN/Pwg+GX35hXXPWDUGO48q+RVm0j6nIVMyaUAWU39AENTJfgjRLOJgEEZtV
bdm1E+tKu9uhwurQ8cFrU6i/DCKUVY62/c6d5yHqQTloAnAJgyJ+FUbV8A2/S2Ck
FVmCBupoxrB1AAPgQgL2TV2ZrX54J9efc9t2OgSalMIsdMnI6UJjgfGSbrwYivC3
VG7tBmIGkOZf1jyuLV5ccED2XWGV8upy9Ym7XKdpr7pPztsGKSqjFJ4RgRplZp2K
fH8GPvgL9y8/dczs9CfK1QKQbnqNCftoATwmNQufsefbBVxhmCZXVISYeI0guZcV
iwZlVDSyDq4w+SB6rDADcrIHFpO9e/CR5jScxaaoiLyI0FVcSNi7bpWrh0myqRSR
K/Uw8Ds+4/MwxKoJkDsGFs0VzNH+jICEg/Pep5GRQs5XUlXTVrY7a5rHLO93gWL2
9G8EB1LwrGJZwLMpKC1wDBrtNLnUNi4BOOK2w0iA1b7qYux0AB9CpNjBi9luyVGn
OWKppQpwE3yPBEoxQs19uzsYUixo2kZXIEGN0WtbsQrg2A5DWnQqOpg0UcirvjV+
pBQxXYFBUYQxnWU7Nd5lOuZuv7s50ikU2LCYMupzJTpPQVnrb3duV2Nvm0luaRCG
ZD+gQjjZKRbRoCfz5b65YwSlmu8dM/6x+dxMDaP9aRkAn8H8hW7bMBSmqUKi9jy4
kXt5Ag/NyUxQqLZzLBHsxq0yXrtAp8DzysTMOCSWHH5U8apBOXRsbZFmFnTGKsgw
CrUNeY6Cbz1i+ZpibsxGbgzvuUpc0WnJMV5v1mQeLWzSVHw4vObhPuOj09rDePoX
PfBiJEN9UQXx2K+jvqvXbM8W52iiHYvgXkvjJtxVETEyPkZk7LSLODAh+HspWVf5
ZhSJLaPg+froDcrhRjuqi33qw7xTpXcvyApNKeGTxVkzhoGmBPCtvNGktq+phkDV
F25tbk7axXs2THY5c7Zsfc1guRhHiUH7YmLHlIyorv5icpMRrR0jr5cM+FviD8z7
7D9OYmOknl1wQX8T2C6A9D4mM2AHCVIwGQdmCbpwLUj1DlaGMM6R3UMJsiVkOWXd
XfW3TAy46ymdRg7cOOZXvYhZB1kHRmiNnAmjWz4DDhJqlRL5d2yj6p0bIzeyB/RE
HdPlEpzsqBtTuZM6+L51ZPzB8YK1HAwt+whVmjmccU6cVa2I5ZXrbUzPtadIdHS8
XWGu3J9Ba1HmHYQRGwctRBEopx36+6oew6jI3HLNMph9wpOMzAdMGD9nXsgZAZvE
XQ4MwcOW9p8W9AvoQjM2nnmrtBSd3+kkNn5YRteXxZWmNIzNg1WMQS8V1/425WSl
wLKNgGXNG5pg5hCHwsaMRk0kJlXkx3kVQo8zz8hHjYNlk92TkEOYcjECjkjBXU34
XGVEJC0IznsuvLPCss8S21SyzpkLvLd83dXZXOYcYyb9YDNRCPvOiedxcg63iNem
oKAETxhR3Q/7j79zOnU49Uwjy/pyshvc0xN1A5dpw8q1ABH35iLdCWx4/dCKO8A2
zGbWJfypXVNogiH49M4Tyd+sBln3SZDsbpO2en9xzhknZBxempI+RiAtn0tW8ieN
AlI0tXDXoq9v2PJ4n+aqT0UrpkzzSiRJCYBtfbUdtdmlDUs1Hy/IBUT8HxF5I1+W
V0f7gM78yMxRgXw68UJ3Bu0OW1mh3fWrv1aRLmBVQQmz5aN4npknE3LqMuXPZJjV
c37ePfYm/8CvDKyMJk2ZWTOPkwD0FPS1Ga5Bkkr+22LNvZchXikeHi0rUoXGmGWg
P7wVZsu3geqRU7Yf/rME0N0p8Cz1vhs7FQcwf8xWN14mb2udmZO369Jk0+5xLheV
zOJqQMKftkVxv/IBgO3Mz+RQO4qWUl/bE5MW2L7G4Aj8FTV7XQmG24V5ibcFcWKr
+fg3ltFFIoGUaPjkGWpAg7rpFlfPfi9wBKW4VhWzDUOpHHkBjycGmH2qtn7xMYap
PgHU0bgGDADN6g7jOycxP8dcIzhu5amcDbspbX1FGZA0Kcys/IwAjzbRVH6V0skk
nqcWprQZMZ4TSWLveiVOerAtCLy5t62osMIWA40ED4gCO7vejWB0RZnzxTUwvCpr
S+TvlmsIkQfTsfAHYh1gt4rE6O1YoZsFcypU39eg5JxQUKbx27/GrFXsWujfuxVM
AyAwgly1QJXrSy6dnAHM6ICnR8e+CKJXqrsJg48Xi972DQxbnn+SJGbEPQ/BGUlT
Yi+DeCDGEENzos4GCSQZoJb4ekrwHhfUg5wBpPQ/ACgL8uTLcDtP88ihNhpZIebE
80weNPh/ADNwMllPPesMcDe+diwbIbnjGwT33PAY9MBCAkix60Si8q8VNNXUU0zT
jPyCJwzqRYIs0t5DhZ4ihKnUBd6ZG80BQcHEgNvYMPvyMerOYT82o5PbyDnqSGsO
4q64W7WUk2LXVdONX5fVBUEX7Ysx6H3rI2QEANQf9KCbyjk1VIwj8ZpTTiCkIKZV
GYMmEtmKp6s0uqaTDrJqkTcAPI6+P8VdAE+34eEZSkh7JKCVrcruu82+34s/caKL
aEON0X3yLr2yzYZzfYgj0Vm5s9MzMeduPeHhaaPSUFYbfQqWERTh9+Mdk/zrv1k9
e41I8vZEhtx3Uvw9M/vuNqL7mnyj3c+xNZllW7A7K7/lji5B5uAGx9+8NZ2ZWM2T
X/A2FRWhRyc4OPiqGoFTcI0cXUHPew6WI4Wfy31xh1WDcASu38b4jPV5QAkd1D1E
MFzIk0Nh562aGv3hbGBl9nx5+RlCYQxgMc2dUOJQvmYZcOVnyM2DfIxlfZSSGekC
3aQMJYy5Q7M22qTd8iidOZf+UGuDC9S85s3/V91yUSY0pwPaKcV33zkNaOz9EEDn
SFK8LYeKu8bU6pXg11hAe0j1+Z3575n2HjKWelFoykeEQgYlZlg7vJOuIxbMrPao
rnGJCVRMm/708MS0rInfFBkuXo9kAE2+1lAnQ+MMYedm1YO9EhIOEfCzhyckxQoM
zG+HyovARjB/pZdV06eoeyXksw14IL1HGClYyoWOBKehy3j/0YvXki0iuXhrgwuU
HPt1RWqLotKje3tKPAiUTu/af64OKbUqZmTmkl+tDcPDrFUUdlm40f628qdpEhgF
uxkrzJeVPI1cUSNesj1Qsexb0rhUgShWMSNhV3EGOKtdBPwzmvJElceREIjbyfxt
1Lr7Cs1YJELAa8EUrG4h2QUw9FaWuXRKWPDfNsosyv5MukNVusuz9aBXxjMUFPXx
0g6mABj5lmsse/9DAoVQu0AUzsKlno+AtoEawr/6rHEY1ARHdnUca5UpAkchHDxZ
qVkaaeWuyW4L4o++YuhaZi1g6GrAxgO/55j91PL8PpLUJsQOjm9BI+/qe/oH+FR5
6FOZaomiai4jCUe3wfSsxo3KlVAvIGqxNxqQ6EAFQYteQzwTnji5yJVgTiCU+Aj9
r08JzkKYPmndoUrSJloujenGKIDU6FVOTgGifN1sOow9FYDMvOXOJrwrDHh/Hhzh
cuKS2vDGl0U12CYoRIv2DLlVBBypiw1NQi5fKo7o2J+R1GVRmUpgdPKKZCzHyPcM
d3zkVEaEktTX/rG7ftC3ZkARmMOscSS73c72vMf7XCS4XA6jYaXW7dZUile1LDo6
DCz0xmlEu3H3WvZXOK6EwKumVejTTijraGU7k/rey4TgMJ8f7dq+mDj/58fC9x2G
chWUrGEEOPAeWR0Ru3h69SAEJEkkA4WbS6WGtzQzYcfho5jHc1YZdTCyJqpFhLgS
C37sgwtY50vHYvKTItp0mZ7VavsQqicGS1J/U27IZC1frgHlgTdkMXVTfe4LZrFB
RLcQ+Hpg0OQ2gxHmaCKxXfOIaT6o/ReErovw48Vxzpu2bSpP29hBBesj/o06iCvJ
bgFcnYlZPpNPw6hjoxzSRiiT1Z7lVs9lxLgxur4KATa3dujYa/BzQ7HWOpEvFS8C
HKxTHhQdkhnL+PZlULrtaM5OoPD+HYDK01msikovHuNV5ROOV3Y4pjQX8i4i6Tcw
6dVzVEgdrYqzj8d7mNiiZXLUwM/bsBNT0534//n/tWfmmJPBGFsNQme2eoIwMGKu
CRFphsaUX+b//VY+iSgTNlhvivMyEltk5PQafjGU5i95d1WrVxV6ljqhmLvVor04
ehLfapgh8/Ky3ypdrqBIlczgl8JVwCqoSHK2IH7YsHoyri8/oux3TZaXbSM/gvFh
OTn0w6ZaNrP70ZhJfTWVfCoEBkq0VdK+HRUkpArQvaSiikJ+LkPZ2AWy1JSfMVOz
DV1ABze5x8Th0FdeJc97fprvAv0CDI/EdiAub+HwZUxVfsFGtNET+YrrfHXyzral
Mv3qg5nLw6mbz4ynyuiJoeZBPZjXdV6gc1fu2UMLZ9wd9Ngw1gQG9V3J13CL+n3a
axzl3CCUGrh/9HHnsvZEw+yTqgIXRZvVTfsz58KEN3vMMjSbLVlIKmr6FGW3Sj2U
UHhWvdwf6LDPbSzKWT7MNAgz5AXSDzhbbshPP6z8kp0DnOud2ZjXla0xaIqXotzd
60tBGtk6/wlqXGw33qQsPxyQN6F8cgL6i3c9XR75SHNHb01jg2olLO+4x+KAolfG
Jf78OIPb+8yw4L/YVbJA8bJOHRuyPxbgbsCccPb0oGfAKJunUs0gnCLHhp/edKB+
Qk9ErxvJLz1mGlcxPRRYP8pdwNSIlLnH1MGPDlvF1xOZCMn6USZum5sdpi3YOTdE
pSZNhSmhdlH6A4vCwQjM+aw/a+MksxM5T9jPqwWza/VzYJl8UOyoH8B2Sd+/njH7
gxVJekVewlLi5D3yuN2CTQQWlM3zCb/xDPpML/utHgMERPEbXFZbhoEIegRmGcL5
jONlCEBtPudIxDrX9446ZVduLunD75APXMIiLHVa86D8XFjWE6u41NUEyvtoVxHj
wHdXeo/7B+L5Kpq0GzQMfyiSSIVMdqRIsa8Dfsofr+KQHtkymPrO7WnJbmlaUdBz
GcBvT9vnrMu9Ed2fu4ZBwf4la99OVi3qi2dgYY9dsEwY6Mk6CMjLVzyoSVH2BuV3
utv2U+wbln2MzL1xTlO4LUeGXHgzGNWWSKRZcLyQhoHAx0YeONf8lG30F74aGgdl
xSeQwyehC4gR+0Oqhgyx0/SG75D9wKWio98eKZTtoyE5sNfiQdcTlcr+GfRkvjly
T5TPANqRaMmJpMaVl/AspZ6XF4BtlOF43+HXFWTNmIU+uAolrxehYjGrs8sHLla2
jvNJjEGu3a9xgukqxJSaxCWsEM/sfcivjRDjRmK/2qII4Y2vKXhcN7UdAz1ruoy2
q+VWAVpz8ldha42XDqAlUSoUmmD11HU8MPM2Wt46D2Y4ZE8/Zlov7WQDKFn+CEDL
WZAxt3AoeGcg1+6IaR89IxXP0Do6w0A6+/5SLHlRBQRHXz2CbUJQd4j1u4l0jwgb
fq/0stMX4mGb9J8STlYZ3vZduC0PriLCIrYE+sgxf4EE+lnWkBxXA1eK6bBWRhvf
ylMKARvgIWXlhgcEQ5LkkxuUgsqgx5B2Bkhz1zhy1dDA6jFkc3Efj1ySNrrtLlJ8
NZUNAVxZnKVswi8Az5tu2+In1ui/mPaIFTXME8FCNKmJ2r561iwMsFBiI6krkO63
X9HT60pOyEchS5ZMH5gKjnRisCf7gdNCEDpcO3bapp3Nzk4t3IzWGB3uJ6NEj9R7
UdSACAtjwNSwHZbMxJeKIdiv5YTnnu8hcHAVo5gii1SGPEZ7cDLNo7MMJjQlTIPx
yveraqhDVuCI5PBW3nXzhZjn1Meo3MnOM+chemx4kvXfo+dNyykuPCLyIBHTBFpM
JbdBKlqvCH+SNRk+lgsqxxlDaNEKPnuXQLpZtAA8tomc6nraezyK6qBo3S1EFCNC
I7dIIFgUwU5GRpbS+IYD0LV0eJpLBzCOmsBvigcFjUDtyTV6R1AqoMtqmpKolmwJ
ecxHOCVvOa44w4jOjBQnYB1DSbxacvtSNPzYfvr0aZu5URVMWwT5rDZIIjGmwrGG
lIq9xRgCypKUCKWGx7hiGsRRklQLr7FcKFsn+qjSLhgTocyFUbiAUb9KBEJAxOKR
0WJvLMa2wCWrxqlpUOyjupA0tK4R2Bty15v9m0Q7fWAgrdMPN0B0l6EixEQG2tPf
PPS1meCcgdNDFLGvyfuAoeuYr/LtFcmA7k5/f4HmQ4wArX+J0vl0PjVrZwP2J767
gbQPyiYhqOAatXPIT643f2UfgixRmdxbyyzt2GUMFDNmQOvZDmiUvQxetBZJjjGb
A1oc/bX8lTqJJj18OQIIIaAaLdqb/qTWZGCiVFj7Qp9aID8etfxnqmD7cUoC+i1W
dJeYhJuaEnsZHtHn5tSWScnp7QA6jVMOiyGtXW0tgqOqS/7vChnlpTJDAi5U55Qg
0BkjLt+qQ8cjG1Fs6RgvJqT5SI0abXtVcij3WB05XP4RkXABx+SGRRX7zJlRNc2w
iVilKrny1F2qsLtX0dg7Y6dKthEhGynwsHU0YeUlYJsMr3ygsHMuvaHMtyaQsxOk
d/sQsk77u3LH7udWgM93d2Vmi20Nfg5x36GdyZUDDAhoqWNycwKzzmHlAgu5IRI1
IjSQh2RQsT4YP0NZEuycYcSCv9Dura6qDq3RuzOxqKICU6XU86Km4Z+3NUHyKXHj
lqHrpNuXZPsCi961rQyjBFvHuNgydJoQ/wT9ffKrsdM9T3hO/ZSakWRfcTzbWNSX
Z6q1Z7ALWWEavZCPMSMpzl/cLJGfrzgsvmJzIqvbQ+4UTWxv5FkzQRqwtTWvPwgM
X2pQ+ayvR4Vz6j2RpctFokmqhZ5jx+Fo6bpYmRAxPcUffDdUuUrS/JiH//Dstk9m
fCJt3Ahp+9BlV4Bp/E+QTtmjd9XdFUwW2iRDFWc+/00+xtzpeix4/n73A+5riAlA
V+tvCA0jBYxXyZiytYkrjQylPq0qrYMf3/7eXPwAkIXVB3iYcNGacXAESayThUL1
OHAQvA9w3j4TH2Btycqw8DnMCixWM5HKFCIWHxMFcpxjld0MYIBK2gorvKaD4kTy
OkaDrVmJ0Umy572JGYOKZvDGk8/imzKsndic27Sr+HuCh/+FLNyDyOrIsrEeTB7q
vE3GYZwtKfoGDf9E5TtoavVi1U1Dn4qs7GChneFiFgs/3YyrLQ4j39kebJm9Pi/i
IgErR35ZsbZhaJBRKyAzhMlk5FffvsijEN3oMrtnQg84Fh2/9/0lLwRa4z+qQxeP
RhmgwCccv3E/A14vdyRx50Lxa6L5Q4vNzm0GP1a5vItCQwBEq1wykuAs/6IdhlR0
O+iSUcnYLooBskp32CwntGANH9cTCXzduMK42Iykllla0ZcjTiS+LMTY9cQRykO+
IA+Nd6DCcOeot5v1+P8ZfvaMVkGdkIYVeqx65Wh99/QrGxFzb9L3VY805D7Q6tR7
Bxeb73j8511P5Pj/r0gLx64lB9tTyzk4QFbAtTJ0+Azn+TbC1tYOKUz9D+M6y6N3
qfEPvXyxM8pwwn0DMV2IJB9MLKd17lKkKgjpIPjLWBl3jEZq6alMV5aPj+GgklR4
hVfPqiDF5+42RUJj2lWUCnTYH9LPgbuYWDt4MB3kIfQhlg/LsxjoDzPGkV1iR/Gj
Z6DekrKggq4O+AWHctOi13lag5zuwXkcf1/odQoqVrUEFwbvK+94nffroXN8T7eb
nsOAG3XbmHHBj03oNgqbXvILn6alVOk6Vr+Up1uUyKMHMtG94++J+1tvZdF/1QDQ
H3WsB1jqxTQ7x7dr+3Dw0qICsQMXkkeQqidh4jEnZ296Ll3AQE9/wolVu3F/D6Hj
gthYWJ3iH3nG3bZE2zZIiVes0IHexT7GlJe0pGWCECoUmYpolPvuVykHnpuSF7u0
uJlY/oceLKCm1/LNH5UuBsc7SlJEkVNzrxjL9Hk6XVjh5nmbbO6LGn0PrRkowZ8G
QAxk8aw9fnhVs90oHbHXKPwOPJE7SoHuIW4BNqF9hd6yPjXqJgtrVePGlZkN6uXE
+jmUZHoxADrtbZwIkg7sOQrju3GVVWTRdLhMMHznSm/KLv9rR/ydY26G+ojVeFo4
NtEdXBZz+D0ddd9NykhZf7Gw1/0YceRrfHFJ1fG7G3GEmj/v4lFmfZrpGh+3hjoY
BLc8mnmMvk+wZI42FL9K/mp1+txS41dvh6bldAcSMKuqd8Vge7N90yfMvl4+g/wl
4IOQMKW9vfYuhEQ36m7UkBc74AMHmEgasrlL5NOkBeUy0guMiyPkr3tBfJttoCK6
kDj6wSHuR04vG+CBsHqkbVNMgyrBioe77hZziEW5579B/EePelEXtvPdYPY6NG7c
Pm4Hmo3owlnc3fIqNz2NztlZns4+w7G5SisZ02iQmEmb+DNgNxGMPmRuqugC5azB
9GZzd7emJ15Mrh78s1vsx5dr1KPtK3sJUgyBLPpRx6GuJodQzyw86lZWGBThlF5k
SX+hnn/NRDQeGJhm02oo/NNZ+MkeB6/8QXCGchrJmZ3WTKJmR8/fZ8Uycu7HDOPz
oSYKienhjei228FQnnNy7eMXqZpI/y0y4Zwe9conrFAGKgTncBiJ93C9ODxxpdnE
y6X8nyD6TaWIHLre7EAeqBBd/27kVrgdIJQT0Mq2OGcFJVx6oqmtEjPIn8oprxOL
kOLIwnc9JiqlG0ePz/r3E1jpxM2ns7ehRnBPemlAcjXJ2n2STZKsuDizBaxALTup
f/TIZT/Sb8sDmMpOl0nw8KTpfKIMJmmqrZ/BMvnqbuUieODW0ZY4kBKwLwm14NxC
TEJrHLw9e6Q5a/HecEmuWt9rf9xRy662l1P9IhsfMU13JlDws9NTClMx6UQx996V
IzZI0RLeh3Lc75QSlekpUYbzaIlaqoHiur95vZa0T9eT8FAYlJI8uGRiphCNSNuj
vL9KhKxgwVHedlhpYfcejcxl7NpDmsC/ABDdMtjM+6gDXwcKdlwbfOgrmq6RdvVL
gl/aCizOF8SHbXH8CBdb3XG49yg0/ACjrjc1hV28Gkh/5WOJvLKac0Bul4IaZgQy
4yQeB0GAW0PAz/47RFcupauk5UHkhFdFo0WxcBdKAtWA0UROxxDFhCtgux8otwH7
CWDQysl8i0MFfDghQeiWhpw95CygPl6RRJpYAObBJnrorURFBL3i1iaB6JtoF3uE
VFb7lK4/9O+6FtwUCd1EFuSgG9gtBsbp9+ZBQORQcraDvQGqrZHsIL8uF9elh2j9
uDrX4AWo9ONxB5zWFZQiKDv7WUcCEBzijjj8oqKunNCb0KtDU/hO2M3UBGHvQ78J
u+vM8KkYMIdfLeTqMeJfdr2VRbXaskq+J1q/GU0sD7TuwLD4TTuodg7L7SlJs5QG
JzqBYFmdVN6u6VdoQLpSVYiXMdFvsV0tH8KvmIobjQf40NRipiGq2vZ29C9V780d
yFTqa/f2HKUqL5dG7huNHD1QEz0MURi4ynmaJO2seJ1uSYd11RL0A13yHDOmYeCF
Bhtd8lBWTtF1w+Jfpv5WRdnhlJNaIsIuej8pwDUfSPRt5kvZObY0WohwS05oktGb
rfiLXvBJ9fq/heYSwhg2CRnAnNYVdV5EmJCczxAIUq4hgBbtjGtEIw2WIQBdbUAu
7Bci38h9q4che60a45sCxaUm8C6Mu8puw0JFVmFnSag0EXRbihUQEFA2AFXTN4e6
EghBaZ/llwxsoNb029mIeNfyRqA/xvIefmrMVtBPAgOr0z+i7z3m3hsU2tEYMwfr
/8Yc77oZBPCdqC8rbFxUREKdtKZ16x6YsTXY3PRdwJ2NzqTiQqlZepUTNfrqP3zl
CrKUXau29dE3ZBj8MNfPO+aVeynsHV9myyqk2B57DdJW2F0P4R4r6G58fHuScRkh
KNAr/g+lHpHEFbK6hxX9ybFhC3ry1ns/PLytYmnVWFqkt3mrORSp01xGoDHBkmI+
t75a7kcI4WeVyaANKNgYYvQL/M/LkX9Prmn7Bn4OKFcD4Nl5gLmw7S2T8Gfjz6QH
cAE8finIyssKIrPscKnT5fA1woEtWjBgSYpu9pnu3erwcRrtWknjRIkoB8PLyn61
5ed9K3ZWHSI/zVb9sCnSKnn47ey4yL8EwA6QZQiAvMKyRRQLk0Hskx3yOCI5ML1z
E1fDdisV8dUpjCK7HbBegMlcrGHWqMVy3Bca0lvbKjQezzAG40bdpOOk8wyYFF2l
mGm2ZHsFY4QuQ8wpuzdKq/qNwgX97Ld9xip5Rl+iSCV3/F6uaqszxbHcNLp2l107
9UU6Ij6LUP5l+FLlKSjs/ZXOqbidJwPYsvsNuA3VBz/CmUTyK5COsWa426gP/4YN
4qqZTlqwdE3ZEQlnjRLEfcoVNUlkFi03Lb6abMJOGixs39Fcygf6cPE1PdXbOzPS
ij8o0NBUqkPhG29FMym3Zq0uTnpYjTOcc6AB5BUdK4uqHu6FhTCiszHF2ycco+cl
kwF8c5mmNbrSn/HnXnXNZGuF8UyJLzL/mUwGGE+ZlMZ5ZxY1hCsL3acpK7k2c6eo
xlHjdKYIFjPwItvbdHWkq55lW3HcHEosqRi8VXNrCY/fV2zx3VhF/l/nu/d/8Evl
aDk/rM3ZZ7wXsFne26BKdnrHW2TNr7nKHvAu0QQcelSS4wgJe/5a0EoTLCND0/je
fGDxMSsvC+H1hUMxefbbFlLj2JhZU/NqzdlXMErNrjkwlic2tWQ/zF1R3lvq8lnd
qgXbdxWqsS1/RF9er0fSzzZYLyxJ4TFnBHQjb9bUYboExhg5AGg0k39afPQ0Uce5
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ARm5xTXmLv5qUl2gMxGNqghsDSlm/fAZ/evtIhYtIDGVJ5YYNuSNASDIqOpfMBiF
EEExc7LfFgVFfjwB7YohyjtosyvAa5i7F22zXrhtWxoVSikRWCdu5Xgy5E7QrL6D
lkRqx8mkudMvBMfUd6VA8SVY0pnKmCIt5xrFh8aM76KEpJBM25kpRPQa3cauJUck
BvE95CQdPS6FBEsnqk+83YWzu2JbmzHKWi3IiCOtOXWqyFQgLWLGOwRhxZ+Ps09y
zStj/hq/kkaNjHHEEGPFxbluDksshGYLdf6sW7hnvSCYtRVR4ebfV1+Q3UIkUmfk
RWfswIxYzj6yyk3Fz2fV+w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22576 )
`pragma protect data_block
+0mg59s534dAdT72GUj5izpySnOQB3wJwjD3hudwWEawnx2jAvJlw89jlErzDdE9
RaY+vJMbFN93T2SHBz0nNbex63fzFz0WrTpXoWnkEkGH1eAOaa4GyvGLJq3PfFKP
PrPphag2PXEgZVskatzKvFFgY4YrMBBS38zSfmZ1FwUlSD7WtVsKyqhHBxxXuGn5
wHxdBI9PWLXN8fNHPza0Osaa5xUWGiHeqztopK6GUWKNZSPGAlU9kr7Wml8R8XeF
Jvj1//C34ggm2e2xvEln/of/8fvDH9ra31a+gW0UYJUXOUvC8TDzChEa3Gq5B/N8
bzwh2KrVDwYkyOv43qrwu7y3o6SVoKs+pNIrfEpV2t2leD2F7LQnqB+ytOx5MRpX
ginmSQrk6YVOlWxj+EBOoa3uwg40jIIANIoNoWLHni/2YElqLvsvcl0juaOiSezv
nfteFt8K9GnObip3ksGS98MKGOsNYnlE6tL/v4kYnkrFyUU6dD6mC5sWhr5KFHb4
EZGzbSIS3dAB7SvrKygHs/5m1pzsgH1wCQBYwscuFXgAo+18ma10kBLXdWHgTWkS
ROUTxxftym6mPgr1hY24dBWDY66F58Buu3v5/tomh39peB9utEYKveSGNZy5FTAm
rySfSJllpk2Pi+pgIQu7K/JyVX19FZZsG8nUQ0Zcd18lY+P6nWgwaPr8U5LiX0+P
m0mM9q7vT0GNQFIqM4WcBcbw08nBVkBkV2cOwKKoCWIdHULcLbuuZtOsnE3NbRXD
gXVd78ZsvsIllb+e0zrWZsSVWuaNi7xnJARky3ryDdmuV2JbK2wzqV1iQdjW1H4S
1hp4MVYlOAor6gpxpfeZK0mCU/p58tRSoZ3+6cWs4Iadiw+pUjRfFbXyaPpz7HGn
Wo92F2BM9SYtv1UgNmvjvwVg6zYiA0lkiDM5oxY1/8kzaNwc5yWU3ueQn1tvmYKA
bgRKq4p9rBaehyWqqSQYvUrpnxl7qN/pZb2vuJ1DqXcFjGCuJ1ykmOHXainKn5pa
dLiMo59h1kKGKrwhhxMSX0w1sJn1VCtD6MB5uCeDWVUOeNx+JAOAXntQQmJlGSHN
vPHDIW1KN2OOdhwptFqDr4ITnV+UXhPsuur2ugl5s7Z/ztUX0QeY02vMI35c31zT
cowE++O64okYEMdY4VbAT6JaODn/yTjkycGZHkdihPfa38IdKNbdJFVQDJU+jscN
PfE6NQgTgDs+JEKxyAKfhzW6oYokrt4uGf2zU6f3m3euynqVMb/v5h8/kfdiFwY+
opyzA4PHHK5Bp7mG3ghqznKqgw0tI0dkeL/FzhBMBbfN35HFFUPtF5yLhcTkrLAT
RDCxVzgAYgGqpOolo9Vv7bDRN6qJNVcJeNmlQqjWLgoyxbQLESWHWATxvAjTfQJ8
5Re13iduM66o0nY1geT7rPP4fvgtH5o7AvvFE8QeJNL9SjV1pFRXiWJ/gWca+zml
cz97UA1w8TtQqQf3beh/W0Pf9j0EW3RumD1Gyg+fpy/GoyiUPapgzOmAbGboY9k4
k3S07ZT6wW0RcH1LFeThwLOuQkTwvR+Unn8pWVZ57Rzc+tfR8IUTvhVOzlOAaIMo
Ah3fCcPyp1YDKQtsQyfnpTLQK8l94r6xiwdNm3qEFrrQeW5RymU0Moa9B17o+hiM
b/w/xZS8WNlrnQmlzcCxZVfbAmewJ+ItKcAZKuPSHaL4mkSy2BhMmaceis45Vp6+
dkGgWPre/QEfdc+HeYugRuaQAgM2IAMCYsxKHUvQyR77n3ufJ8iFEV5TZRa/TxRb
kiHT+JP7tQgct8C8VrFX8R9a/sylosGhyVP8B2zEYHsihKQcRJahXAkFzCRANXic
Xvwzd1LCWdZNGedgwN5fMQWMQdi1A3HdLjVQpmQB3sLXS7suhOqUGAzEl0jtyWYd
V2MREl1O0CoMO1FDP+RUwn+A2Btk6I1MkASC5X+e4wi/0B+JP1CxlwA1kwHUEgYV
qqLqghn/tdWpueGPRSr4sC2xC1k4Keu5vCjaEC4zsqSpQrYNCYAdXtVTK8aXUN+x
DGCnLRSmKbh3KAyxquSCec82ao0xQJNjwuZF6OgZb7oc87pzjF8rUaUu07VdO6UC
n38uEIQXA7pzAuVpCxqN4K6QlQ0dANSj3d7thAGW6Ls9Faa+Fx1LLXZHp58pLnCE
U7DPbbCUwRcqtBo4UEohMod7b3QFoaugAYhBK5EeCvRFnnCuHEitSwAZQ5Tq79Es
yD/BpbRIng15w8WPH0JZAupEj2SD/dEWOsxyzwQTLDEZ7kZs50xXXes3FutlBS2u
hM1XfoD4Wn6eT23PJYinYiMJc4ENKxpf8Ak97AYDvNJjclQG6VmaeEGT8pNMUgcd
XiFmIFGkjLrtLmu+Rqp5Wcu7742Kpde8T8oI4ADKmaFq/M+sJtAu8x2LFXfvHXzK
tNlSdyMW7eQYWIToa95oqdVX+0GE1DLJ6/y75FQRkhw+/VAMp+k1nhsjU1WFo6OQ
Hy8fmMsScY/GcZ851OFVMCC/loTomPi/TvdfdJXtCq+8HraxKy3bLM0bLpMOK6vL
ZV9fya1//yTzz1b3NQLaiBGKRy678ftGtXsb7Qd0u8NaOcQB8y5xsPR3fu8gWnV/
DpyJDfxxd+13RHBqWaUo5gJYYxYXY5tcHd0AKzkx5sFl2WHDEg1cgUxm8n+tqGPW
o2+ypFaMoH5mQKoLPIIgrTVOoS6UO6BIruBESb0Dolf2F3uDrGrGMtTp8ehSpmRA
EyUNb0Ga3tmklYvQKNkZGClFDxZZ1VLWmQiKi+IPfbOamaOJCCngWqcTMOsotKmF
kKLcQYIY2uWI7bMIvZC0GzS2v6NLFsj2BMehhoPAvamg0wKi9yiLyKMo9YM+6xC1
l4W+UE4vI7sH6hP7UUtCrLAnkk4/Hgjgz6fu5vR3MVEB/hUq9TUpupe+G7TFhTV2
IyWxdvpziXk3Vurnmb7GBhKDzUc8uyDo39mrivIRdRTYAPUqXipDHex0GLpBXWye
V1XhqAmS7LNht8JbfnTN7+T9bj58im/Ke4XHDO4xSg2wQ6lf8+57VQj2xG6AMl3N
S06Vy5Js4IQgj5uS3y1HKkm7MnLR5eHPnbEGbTeevFOdJ/eAObZ1HROJMIMKlNzI
5+az0K+IsqVWFeaxB5Z2jQKcFRrL0SMIw/Zip2Nr2hjwQzno4o1x8PK96paVMXCS
hWKCEuoApZKcvaX6RxRxd7iahl/4/9iwOt1UnYceex57MRbzDrlX5kb83efYE6Kg
SdEdBDE7HDkUwraqVpu5uv+HfEV8kiuFCXPlvd/XwAuKHePeSRRL8+dMkWQeX/BA
nqlYpdDCkaQokm+LDx/cFX+sBkueFhHEP40zUZmHl8u6/Ns34PJwy+r02h2jGPCc
2X0Ww7N1uGoC8Fgbb85FmrI0e4HBgonOV0hNaWFGvcR3zslGR/T3xRN1ALZFq21q
yv714HEkQbMxpiJptHP6CUSOAqD18UEr1trf+lqvn02ik+Ei3LU6zmsKJDxRExbF
fwUnSv16J49P+T8sRRXyIViin93ypXZfDX9jTp/qA8vg43BNn61w3jBH3pIMTEaC
MtMGWSHBbjCpLw+cwybg9MPKMz5Nlnm87o+BOTqtekyLvdRBXyaS1cqp9n18SqTj
GJSq/f+R9bzAE/oXBwffrpn2cHbEnvXk4krJLNg1SuvbCpS+Fb7jLqMvUs8NjjBa
kzEVwm0/1YGIEma0xNsk5TjHOy0gJS6rPv+EyDMmPLMrjRdL2ZYfTfIL9v8u8njO
DzcEwSvfgTKjFeU7HE9AoOAV30/kMJ6yfAkbShJDjJIDvkKa0KHVCqee1krD0w5B
dj4ChykdR3H4e+bok7YdQhDueB+ce+celPE6tglzsXRCG40gcPT6V9DhN1P44xhX
DaRF2/j82E72YYTmHzBmJmotT2KjDHaCQxWt/tTEcpWuc+y2OwMhWGGmk8UBSCAi
iQ7MozRKuGbgUxXCKTCOjbqAxAivCi5ggqyeNxPFECw/HOjzDxsEQXg8/W67hFd6
A9nce+Uk4j7h4No/uG8m5oQBqi11BQPZkYfU17Zy2PikuFAKXZ9NVdm2gGqSMx0Y
woj/E3ODiPOR5SRvUOf/a7By4u5zG9qNrQlLV7L9jc+bRCwtCRq2RoW+dA99tuUJ
aeDGnOED8DT+/KjrpGfypPqmH+A/qQItbPThz+Z2NrGRfoSvI3bvJLdL80jwJ5LU
qiAf7cfFzeszO1s7/wk8JR/mDA/wCaGpGbTPCYK2kcsvP+QveIC9Te8QCAW102BE
Ox2CFVR0ISMg2saOH1Fg5ZgVwKJ9HrrGDUnN7bLR/TT2tfI29VzlQhDYX4uybBV0
kaSI2qaZNaTAceqNLMk1qcfKeepcbNmmOyNhsVlz4xgr9cBTguVuYD44m6H4hjlj
wkDZoQc8rXKInaYjGSMs6/9a+0/XOYb8bu+eRwhsmg4ibbyI8ToN3SnkZ2yFIdaE
W7wYUKAzXxElgRsgJJwLvAtyF3oSnLtoEd5eGv+Pik7vPpg2Xh0ZuWQrZaSGTYAN
S4hl2Mf+UoUmLugaZywlj+aLtBh0VvqBcR1X/xYfp1XCsxqPmZwAJM3lst1/X3Wj
L1kqUyAyVMpQZGKz9UXPt1it8gpwxCESEibWobnni+b6HC/cOs6GpUIvq7vOA/UG
/QPQshVSLAGi1l7wmnh/lk+bO7Pf4I6Qg5QW4M8KjUXBI5tWbzkZEHMd241nfrrm
KkY69HPf6W0r1JjpP1HIm3uSH7o6NLdfkto5XM3IeFrF+hUzj5GPPrF37qQ0wWJj
6bhSzyuXnt3ECm2NmneSunVTmM8Hor7pMGbvMLIPB8H2XBJ/o295jizwBQxS0HUm
LmUZTlbFX21qxcYo+OCmKv4o3lyEH4bgjXC/KZr8T3ejU3nDBL71hQRg7fquYKPA
gsu43h5VjhVg3q05jMjo6iVu8cAxULmdljpZFiQCZAKUPUr9bC3W9j3CO3+Uw9If
SjQ5Uy5wKcipwx93lyrPFRCdGEmYs+JX8N/kK7Ge8/drT+iYeAsX2EIODG5U2V3T
K8q3+WFeLN3SVkzALoPnl6C4iIyYjhXuIjSUqtwpqY6ouWabzXvaST9Fy054Rlpi
ShemmWbUJTQ0UteXxfLRUGzOvTwDFi27CTcTivSr+eABqRa1wrgDUBM4Jxk2b7lH
FlbBNoe2XRUGX2eZ2XcLLNdg77Kq8eK1gpwQU5bYR9GJWSkVMLy+uHl1sufLTLEh
4zPSgoqRo5MsgrWNez1o9G605dJrWaaq5JVv8Zo0pUD1S29EgES7HcRI0ogYZVTh
c8ohzRMFzTaO/hMxKwqIOHekJBQ6j+Yr8t6jfdwOJgIHO1b2RTbiij4YTXzaUxLI
ca8Z4iEKYWk7McmgOUzgT1gyspeuQCVGokHrgiUx7t9tOGh81HYlXV0vRu/sNxZN
UUJAKW0HSigI1fWNvAhKhQ+ljWGPHQw6BF0XARYJQ5v0Pyeqp1VfE0nwcOZQZsqz
yKsAoZm3nshoahLmpbuvFi3G5L1fzXaW+e6tZBKozcBNB4akfRSCZAkkHAxmPRs3
OhmgAI0bbqBJDfIs400oCniIMcWmKuzYNt4q83T5/AA9kCf5JTgbOXnZLAZcIBRW
dI9Yp0lYmd05tgI62fGbhNcAPIOQ/Qa90fYI86MAqbL1vBAz60x+7QISedRl5AxX
bhk7W0bzB8IubcUgDGAZDsRtYjrRwkCJ48OpJTgKGp6IvzBx00up8AznB11N8Tta
r88j25xu9fAvXPi1BFOF4wbyoUqwM3egm+zBwgEyEOjktSdQi2tf3g+nfpUst1gU
Zio24Ox8LlOLfCAtI285Xx/VESNpWF1KRiJ5h85psMyHN4kp46+fJSheAMZ7bnMI
CbwjA2uqNadhbKWE0Bj7Te/EDKKMMn9TEhjlmxd/w9HEkDNoTTpuKcH8JXcwYoDr
Li3LT9PZcdkyd3N4fJSn691ylkTc21Jrx8o4zvqbTcbMukF3Cw9B/LfxiaXEDzGq
J4VcfQWCUdouqVWjw4WRr7n9rltJ/ts/+EN5P21bn9XB98UMpG9qgJxB5EFVayee
+bbhX4YvbGX0GkLACZLsX9Vi1rXWOkPmz7kbd72XYKC6u907iwrjGQTIO8C4o+KM
wlUkfXSLPaHx3h0Ir7dmCik0i9w0qEJORemTPvyKmAtbsiWGLGm+apD2PH9lxli9
MUL2BF71wc1wrbHtW4YF7oPPplEN23rkauA1XzNx+amSlk1njFtP0aDLNLsIrJYr
AhSC2NGgOzNEJWbnxpPdjbSf9Hv6N0hAueBtcEsFWiuW3K3HGnXI1EP/1YkM0B0Q
MuruF5kFhXHwEwujA72gm1gQFWREFenq/WJBI7qgiR53BIYsk/L+87z9b6p62m9n
pPnOmxrTcCKRhrp0jQa4TaYjwLrvQHFtqNYygKGvrllGtqGlsMIEIOetM37nrZvF
gfhxXHQftqMTD9yvsu94HjF+v0o3RVRy0d3UIEb9edy4BqdTV0u8qMxXeMaKr1Vf
YmdyDyf4yNQnie8fkhl6dlZjR5s45TBfxAdxxvpKB7KEs5PkHz2Gv9yUQT8EHRtH
zQntmyFBkWxY4QfRz8x42y5gFCZFC+0mmJI5zUKizZnq6Y1z+LEcurCmgz1qN1v0
M7UFf+b2j4jjbbKwGJ2M9sjxjI2LHDChChsT1QyqwDABxtnU9xzBlVo39ATTYw5X
tWnCFk6I+q5kZnEHS8Kufu2BrKnDOXAVFVrh0IRUst+y3B41CSHdKaFIsUcv4nna
G8LQi+3xx+MC+2nyHSmdI/2WmcnwKxEj3J2m1ts1G0YI9akWhkgXsM+eylajhbw6
KmuwTIw45ezvRQ9wZlHe7vqvsWJpml+vx9j4mEBD37Z5EY8J5NVl5xO/GjtvILjb
QpXGUkVPctbRNH79sCvJuVAY4v5T3/kb/j9tuRamQNeRhq7EYxSc3H8z9vx8+HU9
lh6xq06YlLU+LXaq7kHADF5HRf1R32cTgC29mcrYZ+o66eFfp76BrfErhC1GhC8S
VNtHEXU+xPsuca+jI4fEkCAg84SoxVYZLbcBHJZz7eel24gMnDrHJlK0lEwaMPel
4+pGSMBvyxrcfaFqzOO6Rm+HJpu91JPDm4u2epsi5unATOZt9yH1B+361rsWPPWT
/ANJ46J/2l/HY8opywnLfOz8nhgl2SImzFYTQdmxgG704RpPJWngOqayUqIhs/Ap
Ar7ddaw4sYrp5Vrlv6mqgqjAvR75q4u3o44Zf7VTpEQKAfXwaZr8FWXUwXU0xYv5
/c5aFviYEBlrTzAgqv08wA4ZwdvahCykpNQECX0y/F1ZDrTE0gn0yBHH1wDikUiE
eIecnZK9choo0yS/xgAlxBP3P/Hn+9icwvJTS5NTu468LOWVbq9t2TCp8RkT1cRr
Gh8KlkrvhG5WeArBs83X57Pn2RpJAPbYeOGkNYfq0D0E8PJBaiReRauQRphzpZDX
mSAB3o4Zr+7pG7BQq9Xjyam7iBD+Bie2J2JXALFzx4OKZFNPBaqBsRmjQyvw7T8G
if3qbuyktY5gAMmWCDJatea0WVoO5VLHvUyxNLRjORofn7893dMN7aZWL94QwBna
E7ohvB3ND4Kg0ynMcPaASOqQ3biWpNskLdBI1hWa6zDA3kyFp7sLCePABdapCl7b
RbrAjn44AIBAv/l7EkYBVCZMZLFjmGV6QJXCPdg94nwsKuHz9Isb+ewKhrBHzI27
0HtfWRSdKMP+8CSajVn5vdT4Ra+kZfUHPRYS5cPHG9P3BeniTZ0izyaX5F33kYd4
yPgZnNV10bPKU2ZKICDbGcuYdbBCShjY4ZTyI5yHd6lKluxxZ1Tme5YwpAGiMgqp
AYHeW+0YzTFhwG9zAf+Gj+/O3ydMXitlm1KLjrq+eFU/gUGPzdTzsH7V2HKYkfDl
wyJGQTgWDfS3tpce6O4ML/jfXuf7Tp35YaWFR5bYP2rlAi1N9u7TE+bgZzytfGQL
1M4uIrWaU1hYTMo2PfhfyViCtC+FU0jCiDqYsAFN2usyyrQcQsaqoXs+ikxT/7m9
rVBepLrCQk1uvshELLF12Bt9X8b6Bzx+KTHv9EaCAb75PQBkaFAzYy2BXck7lrr1
Z1ZFuxdtQgYtGJarcfQHn4D1+miT2VTPFtTF5rfp5PMuhErxgFPkrIoFVl8HAtUt
MTC24ynR8TaCuD9jHQp6t7bY4r/MU9/RMsDqNE18QZjbsYDOWRQLsWipqkX0xzyY
elxu3gvxFEaUezfrXn/a3FQbDsuk5OQr5cyeghDCbSMSbyNfftvceSRhINZFNOUr
z9mOxrWMBcZfXg7A7tClFSEWe7hIsU5SseM74V5w8efkC55SmKiSVh/SGUeDVppK
cAND5X57q4/rt0NBnOxlpfLTDu7yaNITlktjDW27b1vZp8rPTDfJ2SwDoMvdX/pY
LJBIbgH+mXg02q1zhNVrvpiVg8eda0OX46rtLtyVOkjfeQ5tZQhRQa6wlyqAF4gM
UU8bM3AO7AqxAiTUjbTqFrOS21Ri2EwIbo4GqQ8XfFnqF0pAO/H+kBVOKvMj0+Rd
0cuan2lOvQM1N7gxP8xyv1Joy9b+SMJNEC6W+Jorl4GaOYgOnU9+PB5GTUvvqLJp
gYY3bnJONcb/inlsOmZHQCpmfGIbwIaKlRnymE3DIbZ8jDLF0mPRpZpiYgnTAfJC
HMgOS6EpsQQ0hR3qYR93YMGk03l+/IE6vWLJ31PZ6i1iFIaw4UkbMpyZwgCAWVTp
Y81f6yN5TZ7ABzqjR3czQMdgLyfmJXvPwr2bw0bkWkTn/EBC8rGhBzCjbzEPzRte
wh0iMt8KRKykld4T0rZI2sWLbx1syI9nEXw2PiX2Uq8sbuSdT8paXZYuiy3cvnha
cQr0Xd3tY37x6LIdBfvDa2Wxlr5wwPjcmUMZ3YnlldPD6/JlhWWmE9rbHwdpdkZx
FJG/OqTOvpDWbX+s6w9je+hAOLEhuu2WeoJOie6ywyrVtla/94HMlcXFTb3LA/WN
ptUtldVdFfpucLLKl87UbB4H2H44T08yiM4HESZ/Srnw248zKZFvhD5u53wbouFL
G8lt4gtd4cvJQ9mv1JEhe4T4XhEKjh2x9srX9A8pZDqPdFqr7A6zsfBdiiKmR3CC
y4NIoQFz10O6ZYRRP/gSw8+tpLdzu2J5Bw1X6+MbL0uHhGQ0vckr7IMzCZ5R9S8s
dJ5FgHR1o9+pRHQnK9Bpe+htN4tbljk+IYOg+GO/0e7iV8cwgtgvplqlip/DCqea
oSN+7TmHzSTiLugHUCBM1/v43m0Bvgc0kA6WOR2EY5pr8zJDcMfHVG3pLLURs/i+
fS+B9xqspzuPlzCjmFrbs93MKHCVh2fk+1GuHlrrPKcbw9ugOyXHC2FrhWuysaEP
CEvN/yxmmS6DjpIW+jZ0EJmTHiLZIaLal/eZJGJd+jtZ5sELvE+4ctC6eTCZnl+k
/cB+ZZfOvSHg7WNMjAsoSZDC7UC6uOUA5DwdfTiJGybmj/LOBKdd73AzYh+gy5zc
Vg6GWybuu6Gxu4RkF76D4yM2UQDmgXEhb+SqeDJcKdtyeX03W1TChO7HnxnbdQ2y
R0dxLKsMHiOYcIbsCfmodlHQU8x1W8Q7sDbHAZG3A/2x4YT8tfJdoNcyju/GBbpF
+K3eyMbbPrVZnV0sMxxQy8QybfpMzYavPw9mAxyqsrc5WvzyPSfxelY3hTOuGeGw
pN6nsdST4UmyyFG8LECKAZPNxCj7w5w5DpLhpmyh9sfpTEwzYN2gtZsZ7PQXgzKg
OaNWQeMveExZ2wCJz+e54K24e09aTHblknxwMhXhi8WCs+YIWkBiNHEma3QaPlIC
wjTgLyc6FM61vWP3t1pPAqaYVIWFy8QFnc9Qoo09DqhUecMVjfmI5rM/ppK6LjUD
LgXXVg1TG2YbZtoSyKD4jgnzbdyLUTIPb6DN/AKeo+7cZERXfrQtsTFkJ6PKTgk5
Sd46BMHP5bMI4Mi/CKzZxeStPyAncb7TDErwkxk+Xks7YZ7G9J1l2folQTd/TclG
ogyte/Vq0edd9HIEmZgyE6MHFDGAchuP4PCouC046TawIcZLERC86Zir8Rvx+2zU
Cn5KPa0+TsA4W27lr6SZIKdnuJ7TKtx6AYqzUrR5pStl3Tj0IrZDVSapmI6BJ7Gy
kk4wkpErrHKr7oSH5a1nftv1sZ4MxznSE8Pjeyv2N4R+wuofawLQvSzr0CAWAERJ
WH9hyqN+0Vvn2pgBGRkPCTIcV65k5AhYH+9mgw2jk463eiUHnWp0IE1s9S8+Yeoi
dyYZUdzPF5YcWaJT3wDpK+gT8jasNfTTLfIu3SERn3sRDcJv7/x7bRkrQK7o57aD
1Fb8CVAXapCHkgOLEv+InjqLxLe/uPvyr+SbGop3MFUYUnumaiJkAcEOBcWwv+mW
k37LUEr62cbnyn1PUmzfmeoG18VpcUXDwYlmhOHy7KuKYLA1r5E+IZjzKmjmWF2V
X974PtKogStJmItV+hoWfeviLIirDKtQZOZH7I/xPw1Irc2PFbj8fN+5w3QY546t
EyrqauI4p8Bd66c51UzUa6IQFSLv1Opg2TdfSontatwQ8Qhw55dFwq7MXqTd84Ld
rCyotK3foTQqulYiTgZJuMvntyfAUj9QjQg+QlQq+hWz48mSHUmgfc9w7LdcbMvt
RRNhznd9oaF+ndxVKN52A+f9ACnz9k5zk6HKlvgD5qRvDyBxJVKrojWmiTQRLMNU
Yemo09hTgGk78XladDQHl+pQ90VmO0vLxhTE+KmIjqfGxyUBDsatZsp8KwGs7dOw
sg8z/GXEraPTIxQREUUy5pW23qUYR6WEXAqg079hABbkatmQJh5Cwpdqghtj3hIa
aWxb79pJuYmYqoBMn3IvTYl3ONaBZS/WPUCySUtOiOdRPhOZVng8woHV4uAycTyt
UNtBy4kX3X7sCHBpOHSEZeU4zU/qD4UlNYtc7sfnoKJAWeezJ47druhDBx+oL/zs
XCmZ+dVNBqNR9vpQkwaG+jvYCINjEzt/tD9P+tZckOip1Tf0sfidoPrs/Fe4ZKwE
in5zUcGhLlzeEgnGB5hTnMQyyFGp37gYej2RltN7y4aqnHkg9eSf/+zHSXPUtyps
I2th2F3trzMS2rR0XS+KfJ/ENaEwWqqWRsdoKnkhzRM4XRlOIMKsUHd33kvOoLoe
DiIpKmn/x4avTS78/n6BHCwqAmm92CAfiVE+aNaXOYSUeNrIACO47z6RLcs1JTfY
k+Il/k30L+mkp7QXt0UaSGm5BL/E8dTVcB+mK5MwoR0LxVPIqUVLsxxJH/7L0XIk
sYZflB9dUEKhYnBHh4yYt1u1VxlAIpJT/3Rfl1oCW8xAeCB/9Mb1pWvCUZLbsz1M
48tC8dRLK42vIDItdkkLAXDKusUQ6jzXeEOQjpCUNoEHa2odf40pMtql/dC2TzUI
h04XsANTIFUlgOcpxdGNekyTMbuWW3eL7aQmaTPqP4LhlN8QxJeamUBzjIZjPXRG
1ptCN1MnVq4V3vhcmiT65CC676TjNtevf6/EzbOJRXm+QSSXhU4TXsCnQuc00Xkd
gwQvTXwQoqagK0OMz5s1c1PfW7bOnLSOdXIqe8BFx10eaRga6dgVagH+pTcQe/L7
Jh9/SsSBsMw995cPBv6MKvylPmf35zLS6zJIS6pyR7TL715qCRYHPvcMWoO9gsRI
fqFosirL1w3ZPmR3thAsCPmTPb0GAfURPU96XYEqV2jcxhGHnJr4509oI/kSbV7i
ydyZqCwup0KQ5Ku7ebCGscgBLyP7wAmaClwkkR8kR8vhDluuwCd0/Myo8X5AZKVg
3sAKTwoUh7oOUDVpm0NFFwhyERLsZ657jDeTpobmkCnq1uRgPkoOcLlozRYDefaW
4UR/+WLfJp3dpgJtPh/+5jrnHB+RNt5cHuogAqu0i8VEyjRzMLOVrx0xTrqStn4m
0HwDQBPnCE9OZaQ02uU2HymMfbU0BWF9i46t54H0QA+FAxSKwXodhGk8KRwb0dab
Ou1CjDQzSiUXZ05FrUUkiotjILm2o/fCfuzKRvqtsvw/AddQfFhEEGjvD8r9EbCe
5ANmkR4PxbKYttKeSMRoIvSaN6ueyy3Icz98EKIaQXR3jJ6RwNXz14hDkg83gHYr
ulsXMlatHhWsQJih8HTaz+cdgLcJ9IwA1vhKyPpmF8uo7ZIMmuVFwHvLRniroYVU
zUHNUedoaAX+z4pCd8servDEE3hpcSmZ7eBCvivaaSDOSn5VC5bY0JAQrrYZAycB
5GYWD/s/ecCis7etU5ro26Fi9Rg4inSx5aAX0Pk0TDYpcT1zJxaPm+2V3/5r1BQg
OjrTarWlHfXHNvHo5nHsLOCTWtQ1jPbHDxAILwY7PGEEaY9aOvRI2rZLW65d1MVU
1K//my53TmVOScW3k4cfEApBeHJIplwGBcXnUV2TtTN/CZNeAsalXr/Xlvwv/20w
b+dq7XfUKAnS7C1WS3yrtryjELYX6uXRDZjcxMylAeariqSft8ZD8/KZhywa05i5
NVyQEvnlF+UdtdV2YsH/CP3mRIZ03gkF9tFc+tZe0y09ccoMZD3vUxT0JZyD+a3I
nuQEYGfolWdICl0+6//kc5n6s5wRZ3ZEA7j7ke9ZciYYZ8TylFs9e723iO5nqPds
rc1HJjE3QrwJ11R8doCwPYSnnniujPwG7UoMj3NUVdWYr4kMjsA3W1v7PqX1kIsU
FJY/kGIPQ3Uh7AZiwHwsgIpJdSWymuLzv/sMNXmfT4zdXxce3cihOpKt2EO92JSK
sWun3aFLKwmX1LoLgyYxh2+yeL5xgEk/oPEs1eOTFCy26vvdJrkbDaX+VfNYWI12
yLBLULo9mU6a4vfDoAbeU3TdYzqReq+LxpVWUJTE862y3j0q6DyM8aqZNH+njMVO
X5B2oGgMZkMJCId0fxxiM9zW1xnwBtFqoiD5Q+f19SQGAjzatAJWUzcJqEIKOXYL
ZiztDe14wPDzrsuJX7yisP767ZL58QleETwNmBFxJjZ45J0L6nmPMR6WKor0dO73
yWJhYLApqSYKV/A8jdRLa3Gp8meabqNisUKXmf9H/P/rgOrG2dc5r9Q6Fu5dsdXi
gsaL6cwj9XeUQ+bzmbbcR29i8Hoa4Xuwa5Fx6z7Qp24PV10eH6kulXgPkSBQE4Sz
61I1LLI+/FfbCs0oDm7C5xjPeMyjddctnRn30Yy+al+863MQPNxqJ5EJgXZDxjqv
JDhG/UpNek1AiZIx0eKE3KLH+ss6sx7ZxTpBcM07/tvZbZMV+4o7PGEZe/gcVy6i
ehseJlLwS3tyY9vGBB0d2WqtbJuMTwoa0yPj3u817he98wYivcfIRFP9lpVmX+OZ
VbRF2yBvlv01gQdRv6xWqUBX4/R0NpUEmER+CarHM1gAEeKwMMj8kbyIb39X3988
HeB5Z4J9LD3YCd/sQpMZDjb1NjX1VptLadmVJxu/irIsVp+hNV9ZjjHRybWMtGmq
cllD6ENu6nxnazLFSxwl9V6m9LZPeZXhe/g1y4QCeBFFaiK7gqftGzTPG/kQEDpB
Z9Jm9yJ/7CmGveIVy8SqXc08VS4TTn4a3gEg/B2yjEes6MJffmGBxH4exWjQ4RZB
LfSzePggf/Sm4QEo57FbqH/8Sn5f1o1IBLN4xdYjUJF9UccQBwCg6bfHWBP1Pf48
90cYvE/51ZHxlanWEZMKm5migEjWM3hX3b1phB7zJp5GwBOL8HymjNuS8ovyAzlu
3FZZzfh+hiC57klWKwWyxR3x017VUHcX4NOvjsYPHq/2n70felSEGjwnDpOYSyX7
IBhTcQugugTdiV5CUThMiSl76k3v6iNcDFYHdmQUNJ/vRn2vlov7fdOULIExZCKY
+4Ia4bglcJQzkXWHWVLVytuDaw8uNPGG93kqtBX3c8PvhrVoOSGEcjzIjXxOJ9uu
3dHZlj+/pmns8E9uiMse+atFsaY5obWUtu2y7ePx6zk7tsWpb3TXhBM5Cx3IFGxs
POyA5d7H0yivo5m808OvxrtMEnRqyCo6JRV0qaE80pAXXJsNqRJ66ytfgwk+ZyuR
itvM9QmqZ8CDJIzz9Rh3sy5rdAVc0DHjH2J6u3itoXOXXDt7hRBB7X4NXddq/Spy
gcvXnfBDnF4IeFUAxOy4YjPvabSMVwS/T6TNIZMyD3mJJlakG8RQG8KaH2BFxmS2
PJvvTNapxXL0yhypMuV45iJ7woaUfdrElKd2iOSUtS859kv+q+aBoz2JXAijzy3B
U6noWPZ96bzpZ5P4v3u/TLF9JHEYdu6yfe+rFXaNKCl0fOKcR9x3GwXku/LP0RoB
VN8uBxnSQSbq/X+tIU9hD+e/uVRpPSlQwJ02S/3ZeX4B7DN+MURCZyMCyXzTvu1s
6cpUCNPI4wSoC09GZfQDYgBnvKUp/WWBsn38vGrsupxQlL99AVSw4vCPH9Uq394P
G3c7Q2HpVBFVE5+rx8dcrDNtpqpWSbFzk3pYWz2aHl/5UN8PJLMppjsmQO7YjxGi
Ly0TSklaZNMGVU14jJ6P/chMjvHZA3bMc7Y9lM49fHF9wM1ewI8B2sXPQp9gwVIx
7pOVVH7qGw9kB+1mjCkk8h1C82mDi17r3wOdvtTdrxgJ805d6hjblOC4XxWYFdGy
+X8cw0CIkp6dTxe5vPgmB+643NkZceiGnQLdw857B7pn8kAam0xC4dt0k/HjqGaH
2A8JlyZi40GoVWag2MFGXhpPR7388bo5NU79oJ56HTRc+xrF0y6Aho1y2+nj0+bi
0QP2YcBxflYWTwPT45b0oy6kf3yQgmsEqub/pjCVLdmb36MTrY38Assg3NFRnuT2
kSHgjmKg6tQzUv87UqyzB5QmWOgUv8CyndgLrxPXLP5hEZxhJeJoX0n+XU6jUhfg
9TWt/1QzxbwBsciK55jp3rcmix1rjgvdoon00iWu6IMCeNc7oeDsdiGjCKNTN2x2
+OhuptQsvXiBXTJjz765f0l4VV/Eu8ftOPQ4uGFYP8K8q+q7xJSrv3Ng8Hy6Nypg
yjrBhlQz7JUB6eOE6zMzbznuRpMEQnbtxAI+1ZCxoKohi0kL1zp6fq6/0rXIKEzt
9cKrFoIS+HEN6ezaFbVLYD9f4sKTPETvcCZUrft6U5DpK15e8eae2Pvr4KPski4F
92UulMF3T8OfZArlnzTUDLKswbLUK3I0Zr7oZ3rdp5m9ysC/00D0uohK0245526E
tP7MOSlhLzJxC+KwHVYKHf5Dhh5JeefpzcwChhPrJGwA39EioXVbW50bO+jg1SfD
XDfy9MX3T69JL45P0AITp84FwHFzTO9uCcJyTm6oVNszIGNFqvCUuAyesHxDY/6e
TDHCRN2NdiDaFvbWkiaXMPa8ZEzwcY/BR+GNh8wQSHWn7uJeWLZiH9M7fS80CORw
2+ZgdP70sFsTev1DcaTDE+JqfXIBFnB7qrdrSCt+gHue2YenhmbsRRDujYDC6vv8
AEZyk/us5LJJ2rtPHJd4Tc4dfpHVYxjHqn3+XSMZxQtwlymoib0ngkuirg6HaR2i
Yt70KIdiVPabKIedfFppdU3lzV8hi5Z6EYwKn+8OpSMSgZWuXyjLqfQNEtjRisRE
FIiLHS9FqQ2TK9reYI2AYb6RSZueLMsMgTba+JfdSnUB88iBt7BoW4vAqiT0TTlu
uh8Xa776uq4SRd19rWKcWvTCbDF+1woE/QXRDgQkkR8N4SoS/BxWQLqRl7goqW1k
0x/3TJLpjI5Ocj1bem9iCG/lv2nKo1o7H4ZfD2lKCcaiH5Dcyrsm1ME0o3d56FCV
H13PaEFzFgmnzP10jq4ULEs9BbzpySpQKV0+z/lojfSmwPlFdurf8LWWdKeJXtJj
5Vdg4wlvx/hu1zHJhbJDWdGD9jHkaYZls2+gOcaMCmRhHypq6RFUtIOPDb2RGaRU
d2nGbd+sBySgDZYOC12wvyhMiNBjrXmz6Y4rPtRpGBBqNGpBXbggpgdkcwcrVyVY
rVqzGXP8Vb5AZD7rwlRH239BMed5OgnmvmAVECeSkA8PPj6DcBAdyOQIFCEsUeqX
O0M1i3PrcIaNzxSKCneu+vEbHABF+GvCvnoDPqdoUU3jRLIGJqx7y0HL3CVsz3R7
VdknN46vLrErpLxXuke1iy7Uz2T6MuDFzxcZte7+U027d+Cg6RwC+lQ/Z9X+SCg3
DXgmy8Ne+OENkeuv06UmwCM+y3bk0UCgwp2FDRzmWgxw55kN5uXL/L6VIhxtDkqE
1wEtBxg0Gbkm2o0HwlhcJsysatSBSHzh9LPAZxa7q9dPyj9yRdjkUK4yMwMc92O+
n0JI/d8ySxlkPN/CUKNrGUgQUjUuZWSHPLi5tRjRcqbsAwIlnAAFTRAZCphAbn6p
CHuf5Thq9H3qLl3shjU86dElS0HAEcBlnwrbLE+mxDf2Qg8fArjDdWCOh8uXHU6y
XzS7DCHznMI1bhGO/Eb7yLUQTOkcAPY06Mpk8EXDPvEvREBsAUw6SjGs0MYLWZ4n
5E9G0C3ULLN5ducu3egQG1kqhOFr9qXPJ53wK78lAnmYpQcAiD8+c1IiRa0BOC1Q
peXkDUAuaME5TmmxWetUDRhbx9wS3wKToy9mlRx3A3n6rtNlx9u7MMqF57O4YEfl
TznR8rVnQTmPGjqdA858AcLUUqb880tn5KLFt5wunTw/Rn0wbJpZ/ARuano2Zfmc
zTxM44oQNQEXqEBF4XBMrHm4BFb4z3mEsCR9VbBcVcsXm1Qu3Iu8Qp3oBjFxit4k
tIQk1f9qIB0JeosITRCcIP4ME2zZhehI4mWE2ddxUw26wwtJU1Y6ZFs3Jhi1C5RN
wGqhsNIaYG42o71hARzeyvouO0H0Ic7YIVkgjHxWLAprYG8KIroj9mcYWW3+Qm2x
h1b0nen3XvaV8EpNhXvR4YoBCY10cKn9wr6LgsFEF1TuQpjFIgT75XIpVrPQNu1t
Oh/3BfSfw10DfW/PBEDsOkFHtA57OvJj3d701hpbfqADiTe8W1AG5VwtsgFhZWvq
X47X5HZKHp7lPUoCtGHjrIsNaCtrXVTpcp4UFzIr/XbzabfVBzVMwJeuX3yMRdAc
xPBwynIaYUF9vDMYBdHNO72Hm3UJFwDyHdcaIDelb3Eg7TPpn2iR867ewvEV3VGS
SJcpRjx7Lz73WvyXI/bBjZZHV1NZdh6iLkiBSbdc0HKqhQIbDiiWJokzdfR2hTzb
2TBj/zEqh/YL7dzuVRx8m7LyNgyaV/Y64JnxJe9aMuyTNWnees+/+Ad/PnpZawbS
M2ahDBRQKS1AAYnI0jF05LhnnksPTiiIbP/KAcLrMgTR+9tL7/oCBNz+MQ3PlFpe
Ddm9RuiJ1+McpZHTIYn/rPrHub4yBGSYOvxSkmXSVc9MSG32DpQ3nuY02eSNQy1s
k5KBOox0gHHhB5k03mwOKU1i5ueoyhXfiD/c3M4zmVYfJvnsZ1GX9VziP0S0LDQ4
GtL7wxGh4L8aapchKJ1Awjj1BzuRuT05svOTbrAnL8I7mxvLuHryk+alTB4B5793
HFPfD7qoIVwySRsOVSesndG0zFxqSi+bYzJZw8clum4/TekY2EdQAuKFnXKeTnRp
syHhvI1q7xj7+JyOzPjvaAB94G84JaWSbPKeAD0IkLzKoZcD7pEdPfK1XbQc8AFY
ShLO6gsNQoJZdP9kXLhzR90dmRJqikrYnMQg7laxaO8Y9Tz/j8YhBpbowhmwXq2a
PddnijnbfA6NUJnMmNKkvSu8/kFBCRCCyd2LPVTuEwmY5pDzxKiBiJCfdb1dT2ow
MqsndY41iXHpXKiY6K0IxYS1epXHs8ICX+NA5nG3S6DHjigwuWuyV9kUpzjY5hUG
Q1gxOSC06TyNWtrr/6ChIlMS7XbWHJcANMNFGuknv/JREMCbuS2/cnZMtbAFIN/D
zqpkAel8L5cLleX0GF7sqNSiGD6BHfjPo3qxglkETwNxd/NnldJ1FpE089/pBiNi
f5HZVgn8SyGccIQsyMfTsfKb1Bj16MlZnvRiQsv6oVwknD1y47Ar0wD18rP5Dbm6
UaJRrJCJJ3AzzXQa2o3KGQQSdTNFS1T0bN7sVnfNidfRajbYs2DtGjvFaD9EimAs
Bh00nETI42qPJACadYdPiqL9aSVjfljezFUCuv9AMkIXWTLVr5z14FP3UtkDAMTt
Wu0f0lxh3dcw1VS58xqUD+CnqMjr5CNEke8AQ5zAIkpjvDvLy0cOkxKxrGcXtKcb
EnCgdoe0R8JCcczIVJp5NN342jvMuIAv4rcETJvyH1dAAiB5qqyRi4V+QfYM7yqb
u0SV9LXmQvhaMpjrpZOK4V3LOx8ZBi4O3WpkQEGSj0UvOgOE4p4opq7C7ohJPIpO
WVlOP9zWoaTvsttYa24pZg1XafCxf/z+14tbarYyis9EF3PJRl7F45sRBFpfMrey
U3KinutiJZbpwmzAwKJp8M9aFGaTRJvR/KVRkfoBLsCvbDcjBXiY3ktoUuDSCmZA
SKsBL/++L8u7kHcnfnr92u7KRIuxUwcxfYR9lmXvlnHIm1zCG/0SnzS9qeIG1wVO
fOByJVCd3OpYtUR8Yhlh6X1tATaZeIC5PYJ8VNeO+uoR2ad3LwMnpYgp/t4VotaD
/YP9YE/6gyzu8qyD95f2+niWdGW/RyepY9X6oi+TV1cKz58vQOogH7zYHryqGo7P
LkPhSNLJXQtKaj02o7mTAjENsa239rl52efHa8xb5EF32bH+YtvnC2/qGKMX2gc3
DFRAWlJQEbim+kySf/ePeMJVBpyN9Cq9nNv13nLuzyT/5zF5h/NQLrhxs/rnx9+2
jwINStCKBdl0E+sdlbgEisem7mr5jEW0sfu9PCf4oIdQPwfYTQ0kc0MBFS8dBe5a
LKh5dxNwyLzQ7JwEizyvM5fVXuatC0Ej9rGaAo2TpZ+ngwM4N3ZAcDOM1R3luGVS
GHrdbCUrLlVcjiX0KyXHVpY17dst6L28RPtmg8fB2kOHBNcYmWZRIp0GoqOBRD62
LWrKzm6txEEFe51gLqDeYT36LFCyKQ6dTkK+nUn369mjT4FwPH02UObZNyM7VuKm
dJgqS0gbUpH2zQ5VD8spShB6LkV4+6r82202M0YKcdfoobhBOn9AnI5ZG+gGqvu7
ixw9PF6WMCEQv8aQXu3POTKaZZcurqj/mAzNsXq6JQJhBl3LwK77zWLjRbvcyFF1
3W9ko66stYOKr3OG8NUH7t8p6/0vX4KH8UikNjzGu8XoUaQXGWKKIacDgxw0jHI+
xEb6mscv/5HGfR7qRQjGQms08z7t8/kTRPKyx1DPp01WKF5jb7RdjTtofl8RznT7
JB7THtwZ/Xw9GctL8g3qKUJZvv6u9hL+/vYfMCJAHCSdRnJ/E1vFlqcKMymnKE3M
wc5QE0EO+OwEH09M8+mDC/crbPk858lJOGAy1KEZieBNKJ+RKOaHkdbZCC4NMBIU
HynT+DPzFXjJlHs2qAhgfShZy5FvHEyYz+8kmZtCTHZfbSOwe6LM14e6RBvzhIK1
E0vSRHNrBael875Iur4q4KNxV/VujbnIbmmQE9epEPP6zLWafzHpQ++LgYSU1l1t
5ZjrDd3joHVZJA1ixwzaqGDDKuQ84ioGKj3s6utDYD0GLjexGJ6aMlZQQEmWOuPA
gpNJRA40VY6/o5dhCBAWwrtaD/9I3K/7Ko2nM/BKHFxKtZEYiODz9ctUcDwzDrX2
o3D9bhmT5YfMV8dDDPzbRw6N7b87xkeTHTX+lTHfa0Wq8/PuRvWnDmV0YjKknmzy
JbDHRvd0uslLrMPifwwwnGFQaa2hXUI0Wla1LNL3KhdzgnPspNBmMxc0x01LOqlB
bTrgzILqBcZfu0kem7w0M3zVPa7EHKKma8Rr3D1OYoEYKwexltkg/xSkqdbRSrMr
pVaX2noRIEFNrlji2rOvZnfyJNIQg4VN60LZt4LwhEekY4nrvCwo5SqgbnJTWHyv
G/oaQzuxPTmHAyjeW/K21iyVSDnjVKCO/rg16t/mb3ElEpDpsfx7fib06+qd/xbo
DXvIJo0Ma1w6HFjB6gXD6UwKw1dRoCMV6SVTepBdRMtSLkyScdTwRnvAEQxXuN9i
RMgOsjBoEUsXovMxyhwXlvtetqso8j5eJxlEWMgx1uPR392GVlAxK2+oG7JHjPKw
e4CAxcbM6p+OGq4sWYp1GwrvEHbU8HOzIOBnIgrhlRELhUlPbNFswvcO3niPBj6O
56Bx9+OfXLz9ykdQyOAGzWRy1ImXZYUJgWihxi4XwYQcYh8a5bEqPi3D87GW0n+S
pBR6dz+XzU45XHZE6iwaxjCW0V5p4ra+gyF62eKllT9FHLpdnP6YZDZh4SjfkYI0
ZghYLq5KImO+Z+KgFU48zhxNv4PSS02rAvmZPdBU5R12qfrVSpDW1bub0/14FPj5
GpaNVTZ0sEy+BnbIaF+hFiBw5q/oUlF7A6oJL4pjibkXaORU9Swr1u7GlcaQIJTg
pgKlloyBvy/auAo/PssMQ75i7a7pMeZDknKseZthiUJI820b52kZoR+ifWD5Rb1J
HQM8g8ictBYSwgLklJ1T2TwVtgy/KoayPj3NVJ2+DwKRv3G1LVJwXd4XonrW6yGc
u0IRW2I+4eB7MEYRhwh3tbuytmeu7HyE+0hMBJq0WXiFrItY3aNNA26waqIVNF46
FZ375pNxUo93p+w9FyZiEERqIprnvG96b0ERX0pPvN9vdqnh/y3VF6evoWKMBCf7
K+hlOtoWneAgmAA9oKrH/b5wL2uFM+c7QZ2bafi0mMdfI+DvOB//h7YoEwoO+cMi
u+cfwczEbXivrfXsaNrbFdDKWDbuPp/MBX+3+ttNju+TQ6VcMYbmuCymFnhIFk0u
7POnGBjl5gnMcdMRoajVzAQXy3Fr9WG/t1x9vh/Jw5Ognr8MiQi9qruI//D0ziAW
iovnYMmJG1a5oM7RqGQ9KevtSETR8xE7YqMZTz1ATcg7rnsJRENvg4oerIu12oNX
AdPSHdXRUHbW3uNe8rzh45fcZefZJJ3wZktQb6ipCpQPdCmwl1EIqKup8WaS/rct
R4LcKnq0y1ZHDDgvpbnubQzhaz6AZ9f34Mx0p3zlEPLzaeHfD4GEj/ieYsfYXjYr
ptI/1PrGhBa4+S95Hzz1H3siSrTLcDdlHcW3EySDkHwJidX6wsbshbwlgXtg2urn
arkYgLJxbKr3IEPoPWkRPDn5unre5Wk1VkXwBnCZX/hiquQV1cwUv9W/Qf1BCgmV
VovgPBfJ5yMyhWp8AANA3TWYHpTjDYcMKbB7zEtV6VkcJ64WI1W042kAsSannuPB
bJbmAfLp7KtI0sSEDHE+LpgSrhYgeVRdx2+f7ns3VfyH+lm3hbhPQosp6W/YGRR3
s3QEFSeZf8jJZrUAexR/hBG/YJHujWqCoAMIDopwkqTGr7LjR5UTm/ugs3G6PU/S
O6H5FhLjhXmcwD6hU8S5ciUK4uA14fXRCJ/ayXYuhdZgeqbNjeMLFKBiy/rw+/FU
0TugiSx5jqlJlqrJxaWXDvDg8RA9bVnVGn+BJpuCLt2xFLgFAhsDEZseu0mr/NtY
G5ki8MpH1Mj2FvHfg1ju+hE7b94aH4EpbD8g27ohUlw61AH85ELixOSXKtx3RJqX
nNsxF4OU/RnhBwFBC674cho4bxaiJTW/bu3axMPNna9bibQeLev/gkzTPE9zTZCg
jvXmC+FwmGWBj8qUbtJRe5tdE2k6J8YA6OWcjUgjxd4KhJq2hwvr/57Rx4efBots
V9s8RC9rzKUJygFHYc9ginlp5lG0Rwjq2Z2N6ESpLdadpRH9mW8ZGGvhIvpY1Eph
JncecgDYOAW/peg5IvfH/sdPCvR69ij1613yLMRmHhxyqfKkab5Vize7xjGbmJK6
pxEKqJJ1z/RySlwq0LgztGjEH9+OM/DcdAozSaR6LO63AWczZ0hneKc/r1BdQ8Xd
EX/f4fb3da3WyWIDIkDK+AluXNlEF7imFID7x5cWapS2AncUSTMRxZOtEX6Zk/mX
eLva26EfiplIqSZ902B0rYjEPQQwd08ximuQCGRgl/e90rfRDOcYH69Q+G2EzzOv
Op8a33mmn+kXUlsEGEX1C6B4YWtHWB+qyImE27VeuG1cMwZDJSxslRUzg09njuxZ
WWX23AQ0+1xcniOgsfrLvN7hiOz/xQfoPYV6wLcL9frKzt4pXGsRRcp5MU1QAnfv
2r14RumA9J6DqFun5Fagk0FDViTzB6kjc7twC3bFc8suv4C2DJReJ0XZErI9lsFb
xzTarTa5ZfWFwRZha9F4g5Hfulw3g08J+Db+T0HBeBNB54yZhL3aCbwF2tUmhFMA
47Krn5MFKfRDl6WrADrSdMWMkYQ26Y7Fdk1/kqorRUST9aOmYndWFUslw9beEOHU
6xyYIgppxsEKZe2hQIt/yHHeK6KY9zHgM4fUTxaLRUvwQHtr7lE9zi+wM5QxzmVT
GPekBURgjxK3ue7bdmubbCJYuOhwf1L1q5mQwTrQ9kEteF/3X7VWEBcEd5OStKZ7
Qv/sEQuR3eGvzGJ+DPEVBJjGm+k75NBWskvHwiYI8BSybMX179l3UPPc1nU4gMD+
js0Q4n1xSX/LsUyROJSx2kG6PMrB2PgQH4FIjK76pKr+lacjmvVhQsr9+v8PXGHX
mVMZWDADtiiWHsvmlC+lJXy1wCqoSoxMbVtXtoQ5YRuN2eEGeETL3BhOcI4RWvXt
fsRdsTZImo0TiyQluS+VkCDaD/ifOrmNBNENxWNkfTk4YuhlScfvC7IYMmpRy9n7
DOyNyDmvS5z7ROMvCiOzxBxzFkUdmYUAryHCFZJSI1xZwA4Wp39NAVViljgqBepD
UU1m9aCrebsn1P+7W7LZBxXHK4yfazk0ktO3SZxp5P6HEQ3W8syp3xNUQIIFt7L9
VeMHAzxF3NqusnGNyxvTJ4dZt1R5SYc9efuufMqmKnTp4qbQq9ky6IwzRP5HIa4w
7GC8mm4xfIwc0apyG6uSTsG1rMoVyhmiK3ej0+1U/jDtO7HHk8dMNLhtdvXlA0J/
5oD6iAfXvPhw7xTJbSFZW33ldZPSlPugUTWETERxkTUSRX3z7HMZch9zLlh1ghP3
IpWFDEeqRRkCTFWgn27EwE2INPd2LbNPIee7pmawtkfL+6KFisd23lbYgNUl1cPV
udg8P94DxepMtX3pDdbL+Zi7tD34QxZHLpjNYxelxUd+868grnZexSoWcFyUOjB+
gNKVmPNz8cDwcv4wPy0OPFg84Hc22AlPL7UTlJa7uGjh0hdBGt7IlZVQtQ5Rwear
Q7DbOE04StppHZcAugemtXRhmkBbl/ONmnVOv1E3nUHeRybyu0RibBnJPu/7pHc5
qfrFBv4Blh6qdsfqfWhL7iFoZdEbYIYR55DkshaIRrbEmSPQV6bUQCF2Mv9pA2mh
5uPHI1ef4rm4Jab/MC5goVQgVUGjSBBbTi/+eoC54oAIshyV4CEZDuYEBR9bNXFl
qGgkVf/13iBKYdHn19J6MCT9grwRS1AiP/bze8UJnmrcZPx3yaQpahaXtCFYsO9d
z/n4qQeUTyOMKYiWTI6zao/ABUBurS63exzCIQeEs9lBN20j0lhADiyYbWeInWX6
RApoAGw3dbE4HmPOifxVknWfHf3whSrMk1mx0uh9gJfVOej2A6trsDHZdSQkMYG7
NTBCfdg+EzSLQldGiEF130r8rHMK18Aag8eAkmQ151BewXGl0F2jSJBF9MWM9KoK
x2ozsva1EbytYq8RQtIu1+vQnMs/RC0RCxbvFswHVO8plkwieTux/IZ2vaLdA0UL
NaKpcpFQ2BJfhLsuI+K7zVZbemP4s+9hbUfb8n60AZw0C8z4CEv3E8AHgVEN6a1I
j7os9rN7ngBNuuvzzHukm+vx25Q92nCKOPd9ky9r9xeuqpVVNE+pkkiUCMuK+MA2
BjVKb8ERHQsM2GItle0CAiBsq3FPstkGNkgYjWEVSqGl4aiIPXfMhhSvF8yQFD5h
eN4Zssh3Trr9WdBC+Fm7NbLwHqI6JLJ+lKJt1QSaVaCrAHwNgahO3JkToSsiiYiD
pQZ9iiFNID46k2kTGb0YuDZvGfpQpIAXbQQXy5fsUDuFKCvwSvCF0k0xQSye8aDO
k5u5GcOc7uVXuOAvdtBc+sEqGqhsifxrrBhtWiDupInpbyAjEknWwZWwahCJBLRf
tRdu+56FNH9Klw+otLqLzbfzZ7KvqzKpR+W8qLuZLauG+JgQUv6MP280c0ea8t1T
QJd5D4SxicTpEUh5+OSaK4Tmh4XHliPGojOZ5bzIuRPY9/3+PGf6lmrPfQEIDhVa
6vzeE4hHa2MnL52jmOqRpBZ2waW7UEp9WyujpvgmlikmKa0dZzMDR8eJhFgXx6Oe
t3uF7Na/QJISfRF9Q8nmA3vt5Rz5K+LplvJMph77GjTIgEBqsbwh3ephccAzvILn
hH/oP653AYdsZqxKkZzS+a0edoUS3AYxk74R8KL9lajEQTjqgBEPeyxtUZ6cuBjp
b/874GYhnLowtV+mM65Q3ehJAHvBI2TLRb1JDigg6To3DWREkC7UTgQBkWs6+Ipg
h17HaT8FOichLtvaflbh9MdQ+pC7wVWaTBQSP0h86GY40gE3/cduVHHJCJ1Hsnm5
itRwMHtymX0xczExQNs/yuz3w8Jtfm46NmDI9OWAshrk7UjKAjMsleQs3wpTK0SK
tFt4a4ibox6dV+5q6FLaxhMbXvXcw91leeiPku0FDGiN6sJjKX49X5+W4bI7yvUV
vaG0xIWlD49GLCGlHdJhVdMo6w/exKXO4nXZvtk8IwRwAwLOnOLvzbQmwdC5adX4
HpnCqaTVLiNrPIWA4QY1IezfL5C1g4RULBAanjqBgViTWRaNodBnjaJr/UMxIJs9
bcOCkntF1DX508amJeA9V+6nXrZkZjGuvY+H/hjW47iGneDhsMmiZGY3AHiY2jbf
aN5wDufEzNxgPF0SOnjX9nSz0aJJimSB4zpp3VuF0UMh0ybIWPJAY4r2zzxaVAVA
qChxinjRFm2KYqTo93SELkXuSKH8SMZjzcq5RqVVeb9GmAAg1gQj67nZIWkbh3gP
7Boxig+OmcVyk/250zKIk0Mu2XYYImGaGaClFuYj7lc/OLrEj3m7jUwzQZpViUTt
uKwuoWkt7jqRWNNANU7GpQwdz/p+oh1p+62cvTzdLFGnEGeYP9cYrr5/ijFiTdrP
3grABUVs0NiD43gpx9zkgCktob0Tu1RBaKkSNioC/hXnUMFt+cBATqyF7U+VTMUr
IQvnrB8TAOdrT9dYRpLL+ascc+7INa/h14gUiFBiy2P/tR+3S4iGRJNfnXeetla8
8NEg92D82vHHD08xkXDDFYFU1fzXjeFSiE9D8WPboCIoZLT9Bjsd0vobEtH07oQO
mgNY6WyzTjGufTiHtBtFIb7//7138nen44mS6b27OUouX9k+qNK6FAbBf7unqmFH
vBsD5sOxY5GQL1V2ZREvYKKrMF5kdlhl+BSHc0SG5gtPZzXwBR6LOtsi3Obu4o4g
Fpy1NRxi00WRB9pUA93XZSH0IEtZ4EfO8yGwhL3H4te3HrF+jxYdNQb3P6ISSDCO
HH8PHfWgGTGnEq9+7Euu6x2K+xR8Usz7AYa/Ql0n7RWwJS4++THwkIGEMYduZQdg
W5jkjuPUInVbZf7JUR1+D3sabV4IErm9bZsYYiEHcMuhXokVhouFipsCe9hHAME8
5YaIOTutF1h3hDCswtI/bqxM8EWqKQVL2QzSXsGPheEF55Tq78Pk+aIcxksnZ2ux
fe4ZWjmrPE8LXD2Q+kK1ufHqSLxtRPuXNxjH8SXIsufZQ1AztJcKeYMuQcr7gYNT
km4nfHS3Bll1XDyYeMznjJYDgQPi+kf9ZlkrcZsSX7aThf3ZSjkhBs1hIBRmoAup
jz+ES2dt+lTBMQ6PRFfHXdoZmG+yglJdyksRGeMBS3S6wduAy/yEhXXxZlzDzJWC
QoRaDwHgiwOtPySwZ7chSFEHw8zjxnchURpbZCo2casXJp9p5FL0u4mX0MncDzZj
9H7F9ySkSUkD8XCgffgwKuuzFTk4kqN6GC6t3FbMzFUGzR28P3tfEg4QZP3VFY5h
0diy/IjnuWyaM5g8ip0PWV3tPks2HwO8U9Xzrl+jvp9kacGAsGxvM8uU6ZXmgvKJ
yj5aFzpULX9CGPsWzfRIxW/SUzp7LkYsVGEoQdPmQAuD/2F1cdWSXo8XTIf8uWsl
5vWSirl2l7L7mw/QWK+CmVy/u+uUhL23/ZtLUr1cphjsi9BWla/aLNctNR32S1fs
nORP92ADcLo8gSn8qC9xHdGrV4xouRk93JCWnu1wGR99Ir1hGzrndw3LS69iuZKK
pD1zI4zyZQntFroIU8YYnZVyd8CwW9Dv2ubjaFdX+Oeab1ySFMslZ2Sci1CA5UgR
YVcAyNKvtHWEynwwMq878nRKw+fG5F0qmCH5rfd/uonSYZK1lQHm22so6RbL29ia
31ukH2S9aBuB2W23iBxmqkq9lGypUdTlk3Ga+Fvt9rHgwEGhCpd+gVyLitsEdxkM
Rigj9TP3kVrLKNwQtoSx48Od7ShjlgvFqhV2/Z4TO8zq0PY4JWVVV+VbzF+VkIRS
ZXB/WOOHaCWYvCZUG7WhL5KpH04Qn8alcmLbIy38Q+R/XTYCna3unqFQb6SJzVsD
gGW04dgs9abixAw4dQmUV53rRliJs6Pxhllf9aJKfIZuCsJRWP3IW6se0nNjJ9Fa
vWB1lhnGm9XK8DdNnMWaJ6ZrqFgOtR96BRSVJ0G2ZPZtUD++LCMu7ydhZYwI6rhV
ZjxL5BV9+gCYqjzGxunulfJIItSEtqAmHK4H1IghvSAJnWSh5OwDlHTfxkJwV+B/
dM9MU5LFu+QZw9UCOSqZzGkMJ94BBXEO8lmM4pWUyM1MNEjglDV/BY5i/5Cs4jXU
Mf15qKV1jD6FgCuSskwQyyGJu9cnkSeCvLfeyDDLX064aZq3uPmdDL0wjh8hyWMV
zLgCDP74ikDw/R9B2TIuNccx1RAzLOBBA9lXlfAQDdx0cOENFXih9mM3oUKBa+13
3yfSKDJkNfrFAV6MJ2PjNuvpJ+UAVMASZUliBseC2O7DD+xzLHZxGWrKUqoeqLNM
PHK/MFltRdtGVFsDkMl9XYZMfd/1J+a4e/1PnFhWyaZY9C0zQ12bb3IKE5cScJ28
/cgVCx0ZssQNdNRUacpw6vKh5tvSnERajAhMai0iGO7o4csl8YABOpjEwG0r5BVe
5eYrYWAOuzGRtmYvOtc1tra29jgvU5KaoVpuxebp6AdQfr5EKDp2N4AKXf42VOWJ
CgDqbAxCC6rg2TeMaNJopQ4X/SDhzKGln3TrXyDvZn2+7C4AyAAhCHzJ+nv9NbLZ
bGpWU4wEbRXWpYgg8O42i5Qmlvk1SkON28dPii5iNJ/Thj3Gre17WNg0PhS0nZuK
RRq5bPD8cKAcUFRmTjyvq1v9bIAtLY2J5NuiYhaHBh3yvH034vS3sLNNqtswmhtU
bw9dBsajU3+MhgrOk1nfnN+Vg0Xbpk5RpiYleS8UHN9HhLS9z+RZpL1bc0GCZDtI
pWjpEDlUwPBWeokm8xscYLMufIYjY8eFFWGFDY8lwclrfmIHx6Q8wRUbk7kpThHa
t/O4j39u7O4HT2KUebM4qcsyNeNXqUnO5guBJM1jXVWOLNF67jWDWyeND0WFlLZy
87A/7WDYam8Gd1NA3IPPfylE3lP4Qx7oDNvhxcY3M8KmmrruQCt86ZpsNG0imbhh
2KS5jHzJSy+9d59BBjppTHNgPF3OjZbRskiUpKZoAx+i3L7siNDCAUxLq83UcGzx
RntRKbe0QbgbyOxxMEsW0lzH9ObBHwQwNfVxYc6NKDAwnATAjowbmCTrp+ZhsV8i
fJa1fD3HnHhsow+hdjdhUlDn35gYaNZ2U0FaWpuzPK47+oQKeqUH4FPSJTF3Pvyu
kBI7VQ8iu3hpjpoOqzmol4FGv4iZiv17EODVGY9Y8pbVEYmplIS9F2wySCF9H9ob
eyjR+31FVrwVn3mw/4JaLwlnEEYVPRBxhf1NXb1IhpsOwvhy1Syi2bcy/19RahYT
+XASgkgDMOvR+cxWDpYbilgRLINCh31H9ZtmwJOOcQzBJNHFsG+FyYyK/ODaIqT9
+C4v58v09oEONWwgK8V/igNMb2Iq37T0nU0sWnxEaqCpQtOWsgem56AP90u8WEak
iz+13tnSLSU/fNOyFl0u0vgB2etwG/9Tm2cm2RVIwtppp5eKhyNXRvCiK4V42and
oKjz/RBN4bK8jo8XcO6irV5aJQTbvZmPPEaMTlpfe9eg1MmjRNfZEh5CvXbHlap4
oMlb13l5lraOgwfrzpgdUdbEa9XYSwa73iJxpni6EfVyuZwEacVgjrJhzRuWetNh
DyNAvw/GHRjKAIH7nEMsfyF8CWs0RCF7e/ReZLFo3xg9zZ8SJeUaD25zFSdOocmj
JrRtFsyAp6O7b3Z8s4edREEGzMyTXkK58sQ5cFCfOQ/ltaIFYhtuho+aeVhWnE4J
hW7rBePaagcm8b450CQ6zu2Uj09bzP+nCIMiXFcjkdtTmx6Poj+aARMA5PJdu6vV
NjJQOyD5+D3TnduS8DrrK4ek6RZmdwkXIReOoNBvXd7rcyrlfBGLulIPlisYLHTG
irAqtrCRIC4Kri0qGO3OsalApFGC88j1MTkiDMhYv06RDVtNYWRymQudB0afy+2G
JHHvDc0lxaj7m0AyLJtv/NSDMJPb1C9Ivg9e8fQ2PuDdFGepP2QpRkcLYqIC1ei4
tMelHFHr3bmb/+1PcNiSXIcOaXIUZzpjV5hQX77Mpb1R7NY6Cgtb8lgFzCImYmLz
bddMgCiarVZcFhqkm9i+w13bfiyZn9aK3esiL+lhaQotkAK5TBKli+DK/9HK6Ha7
6buxLV/1sWfY3ga7Lyj3kUg4F6Qogfpo+9dW7HsJ/ZPVh2kA9tJXlS1Yabwt2SH9
BKJho4fxW+jS5pah9ekbGDCrxVM2Y49CaeuaaqjxEl2ZlMIhN3TTZw+oGR3tzSaw
OBRgAK0R0aF/oMRzVBZSqa/jSAikJcO0VDCRwCgJSBZZ0fIi9JtDr2SNgFZGrauB
Zi2kcsYNNmI/0xVQYE4HnZ30ceWXFlyRtJCC2/4LpCfXaehLEMbpgRVcvctib5vW
dwngnHnAJTBafR3gSFMKmNcfovuSc4Z01TUO+ReeyrKT94U61l6TyRt6Cn1TlJWT
iPQS18fhRRUs1RW11yI35Ebn5LytGA++iO8CxNnYiiPt2/q+YQrBQrqgSQfllOVo
DX8v4tVHVxwiyEnSBz7l18MQe5q9LFsTwqGKt8jM2UQl7qOypwepzl3aUxqFgjhe
mqHsDH6bOgA4W+/EbQrnnV6ClxoOT5dnzVpv2Mq8cfo2ft7MbtM8/SoVSPI5V7+9
sPdXnf93T3RLc6WeMTJMwCCABmkpbcLnBIRte7QClnYV0tnN3gs+Qidun6JjH1CP
ktd9vVDmzHEFi61EloQNlxP3gdkS9L04z99sUhJes7m+PtMkaNXWhho59h6bFt1i
dk2m0T9SDy2dVQhgcnyDwSR37txt+uAgC4zq8Hm/rvlKxzRpMxw8t7twHMLokvDP
FTS65JzSmdtrOEszKf/gRUWspa49t+9BNztiYGdcgQY9bFhMl+K104dKFomch65G
vq4Cq2nP4YA9vTZlTNjp+T8alxst0YakH+cjX1Vv3qpkQPGwcqFNWxGw8XkmxK/y
3fUVudPUy48aa6ofiXETcZl7prI+qQLU5uHXVOH1re5iEhFig0hlTDIa7fDRPNxC
M5VCG7pdlIfyP4GjfI0dF4OO42MVfVhExHG1aizXG0smoS7xGHfzkyBbSyv3fBzy
mWFyTAIK3njdx7ZViX0uySD4/dct0r7+rM17DujSYO66P+FNqXUJlQ2bQk1ft2WK
H19zdjNDj+yu2FYk28kerKCcNCl9zkc3L/6QICniicqK+Z2lmG8Ar0Q80NMSoLuf
WnsNFMKQsVbaCv43XxAZdjmsnn6kazvMv3zsOImNJ3v+qi2tzF/rbalSj1dn+qTM
k+XzdEUC3ou9wrmRrOufjw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
PdI3TWOzp7YhkAIglA0ZUNoKIC8E1ErXuM6zRLyzZzdjkL4vL65botsEGJ8QZ8aq
gWnZxON/sXZCdeARyoOHpQO+P55lqq1D0Mx3o8ULxTTX4Z/8Lx2fcsvY3Nxs12zP
OPuujdYVg0SyeJFDbR1uJKF7aSp37z0ke1TMkwWW/Yc84cLckM7feMLk4iLdDBh9
N9YQptdB9nQg15RzwMvZx7DjRp+7/RK+/hEw/qSGNwZA20yfjeNSkk/S+pGxvcNm
hywKvmwcA1hakVz63myD/RtkgjATZIaA03ck2bq0+3vr4PEPY07L3k8UYJZQfc4Y
ZJlZI560KSZcR8cpI7umnA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6496 )
`pragma protect data_block
PYLKenpJZZUO3ZALg+9rOJ/zP4xAaLYEiK7GBJIWJZMtkhMJSBxkE7pHdMl3+QN6
NPamHZvnW0Zhevvj77RHI13zGah4hyGIy3P8QN+42m0rvjwjoOFXMR5M2Vitg7a4
OQi7QTK+ghoYIR4Zn11uGxtYdu6zei1iM22v+N86G3NmpdF4FaIsfeVfqZsvDsu4
1oZllISyjA4qNPJcIYAzIVeuqL+FOh9FY15aSrgUBvbWSOyUQEkcvMEzILpUJN9x
EcjrjGX7ugz4Dz0r1XhJoOA42calRPIxWjfeBllLwvute5ixvWxwP3KubocwRy6x
jQzgQ27/UVg+gY/LBQbpWACVYSYMqWJUeH9/0VmRR7qTFn78TyFAcc7Joe531+dj
5FxEQPs2LlSOZ0k7+/n4D7IHp9Rhfn8qIxQQbidQ3EjfHXrff6TQlsklBuVIpnv/
BUuqEC1+P/m9MGBc2VBdnXAwinPDsAylqycPiV2f6fhtN/0LBIcfeCh80BiASxUE
9feIdDo00ZZOaB66wYvb2UnnDWZ4Bv2Ea3iNbK9+y+vyu0yOfohR7HAMp9LX755b
PSt6AJc4KZ3DH+GiCajBwQ28+ojwVOe/N0SxR8lfBz4XdvDHnYon/l7qcGkZj0Za
6gmKyLg5QN7nRqG/g//HxpqpNTzKMC+6CVSf5HpcTLmWuGGOFiMNUqm632gHSG5i
96djCz4SZ6u0e0F6guDu8cVVm1+O+1GCgWbnvs0DNhVKZc3YxPgXDwfpkRiNBfp2
3OeOd9Lh0lDcPkLd3XPbV/MO1gHDClB2pqDlkRriESl5U/4Rb0nzoev2OlJEeCcV
pNiBaD1RTuXAZFdjVciEHFz4aD9rGkO1x6t+B89F+VkbPXnixt4OS2jZqCFoigxx
GBXuRWY4u1CpL4zzhOyRSGFxGyXcwBNsUZ5zx4pwbVKL0JqzrFubzsf+PoOXsxVn
ZuA8AD+qFXvAfTZwPtGwSOZw5xfApnNCprsWaHneIVN9H8X6Nn4BLeya3Dv7BQPI
5S6RmUfPlp6pGQodfoF8M9FUcJqM8reK7iNlRQ5gcgfE+yfTdZy3EePQ7qhaHnBd
tPar+5BnNOB8gikdT5m+c+veXqIRL2RSIMMRSDkl/VxmKUtcctr8ED0NFCSICIEv
vu/s2KeyoQ04NK2eopRAyN0qao94EPYTZ5o5W6ftV9JJ+1xivT68cgc8SRKPIEur
YXSqC7TbBdFFK7dyDC/KlkcBY9tShBYN+6cqvSeko3H0Ty3ckjT5xaKR5orAqJDr
Zc21JVtpHV0JQWwGWbpt8FLHYQUV9q/1Fuj+UzYA27hqo8VHnDdCb6o4x5m6pkQH
GGLy1ISbZOsWtdJw0oRXLxLSUgrBF252Cqad3bsTt0SRfCi2zNfJXsJkYs2XDLHV
P86VlMSn/9Iv3jha06g3FSjuhWT7vkmB9Hzey5gHqQ8VvA8ejmG+8NRVDFB/adtQ
ex9ySCkO0kqzuvPfJ7JLLHfjnglrc61itu5+yLOEUEGxhYp0qfNf2YA5XoLIOLTR
mtZrdiZo00jy/1BIc+8cACr4h9Trbd4wy2cWJZt0guDGIQQ7HCqWecXTI9yIQFXI
1IOkgpW44ovQb/pZhc7rztbcmtkSyt+uBoQxUZKqcWOSMrJ4S6rtSdHX03KyknKH
N0gnTVy2L29FtjaAH/QWyynO0bwKATheeHuqHHn4QzQXzgWO8wNL8zbNYDrKnU9V
Rnk48inMcNBcu5vZOK1n/z5Eg3VsyzX9h6I+8IqxzMw3h23dqBWyWEr+cGEkCAPC
90tu587uasbge6L0YSeV832sI4sH9i41TwxP4LT3YYOOX+KGxzA6NWG29f3yn0ly
OJlKm8EbN/smyfMC4PAAFaR7f9y1RjUVHXsNtzvSiaX1y2GX25PPkSgeI+7lwjzn
XS75pH86UTyy9VGFzWXvrCr7UkuUs37Guzw6Hzr6bx8CsZGBvAYOQ9CQC1Q8doiy
6mTJSHLrYasYx2DtbATPcI911HN58OdMlME61oj5Anf3Om1qAADjLYKXb70fGcSJ
Ngk86KlDQzJjLi6V2w6JRGz2JwREBuHRn9mskAyqgSBhVYXPjf5Fn7lIGCQDAFPY
pNf7LL1lXNYuLN2NEHdDyrZqYu6T50ehI5O4OUmnLDs4qIQ6j5CHM8eDPPy5EL++
RkROvYzUX0JhlnjglCQAzGN82nAGJffYtCVgNfceL0gqMSW70YWvvu2lJH/p/Bnm
nTt8bqCc9DdUb2AMOWGznxAoviSj2ntrTAFKbnk9PkJou1oHEnOaV2n/1eTledq3
Z6DBGANEJthfjF3NAWveh5cb1WcJUcVeqA5kFQLYrHPPxXwemTv5ASgCztdZMYV2
/+BovAq7M4T1vu1VYuBcbHY/7cBO0VjwjIDOFhdmIvZgiPn8UZY8Gm7obXuYsMpu
1gIbDfX6DFgL3OMS+q66y2O75gA147fw8coIdNqWU4TOLHFgiweWTKn6MDPJryE6
eY2yE57TDJ2l0JRBPnpPj4H7GC+f5wxch4D7CtM7+WlFBw+YB+Uu6eT0Ej7RoZeC
XGba03Lbnxp1Uhtmhlk8nNTPuokrbqAOtRG370VKXKatzuBmOy5qQ5VHhnT1wo9B
0GduNylTeRT+5d3w+eOSX1diDedVpo/2PGp+VLJF5mPNfhhNThu28Xsw8zHCGE2V
KbScN+jsAvrX2TdTGh/cUtWQuYY/BY5fd0pYpgl1h+TIU7jbulQtS3Omj6mlB4lE
c9EPJKic3d1hhneT46c3+3AruJrsRv6P7BNfxJJRHGHUSfSpqDAU3+6WSxArbyOS
igcpuqQWg2EnU/CngwGxWYjQRQaETBCdTggitsbbqlPF7llSus9R4QtB3Ey9uTdZ
/JNBoHG3amLJcrZXC+h9abze3d/c7XpX7VbKkGykOPLhPSg7sQwU+2LJOTCFgeFl
8SFWtVKshqGnrslp/gbllKBx9Er8UASEYbhDUU/ca6seTyFJy+8T50ruKOOH4Hw5
rC3BQdjibxpylPhnjAhiJZmWVmiQ+vX8DnpqOo5GYrPmK53K9lvK5Z+EcAQnqB3m
OTBZkbrtANHp5l/szYcfmAUje1O57Sy1+Z/7oX3fbw9WZEfPqvepi3I8p0lJ+3pI
mPlg/SQPxuhBIe1HcJtv2jjv+uAoIklDn99TPW0o7Em4tclS7H/gqN8WnRr9CBQH
Lj7W2eb2qKRWRMpu8gteI5OzzlSULVGDGf4FEFnjM5eQKnNKJloWIeoXpFq/mu1+
NNa7NpSyPkkfYeEGbQ45IIXgnjutYYxLurFYq+PGzuX+Bsc8dsP4jgn/5TTZ1znU
0wB5kQNJtPus2AOT9Y0JJM6DPR9BDW0KrQxMVtPfhfpiqAWnr5Q02RwvBqUUa+H9
aFbrgVlXY+LBisyl2pA91qA9lavKwb90vF+8dMEco1rQvT31l3DyvQLjNGEVpMgC
i2uhoP3Ne8+bX92CaIOlYwgsmglEDdmosdm+LDbApeMrQiFA0mDxniyZTcfN7PcF
eaQIqLdM6sMyDeooI0y+oELB4P5hEf4hRUU3JhsariMdozFgmN4TGVkPzx5nqAuR
BR8ZSJ4DXFwwuW+KYGr5awS4xJcdDe8onLohGg8SC6aoK8WVgGb5aoyAoYr/GOTJ
1RMbYD2VYpngVHWZmLeCv1prQiP9MMUm6nnAGB4VzgjLsHN5D45j+mJ5AkNR0Sm4
XA9Icr1zsz6vhVPVzg+vhJtrreI/U+kn0ns1udMTEz9kQdljQTXLcZeKi3e9WPSG
6fVLGytCzUaW2yVVJX2MmDOu/fkqE2AfzLe571U+cawOknlqEmH32JtKV8utSXRt
zQDzNw8M2DdWy3eoV5ynBCtwL2pIqIrqabFEk8or+w/1HLYPdiYUIjtTNc8sqMb4
G9KbPIjEzqmzU5ZMI7PPUKbK/b3iN1d2otPqpTjGjqR8OqAXZgxCcof0NEkval3g
Lg3/9J65k80N3FhVQGmTmnzorqqqYL6Cxn3577zpr5VZxztQ0QytkLHlceek5GVw
yjcB5KS19vz+Z4SxkJ8Gw/QzsJh5BwmMJK1TQp07/bVvCVApxxUj+oRqq8pu2skI
VzVN2nE2yxNAbnqGICHGMhTa9xLQhB/5JKXq1/M4s3PcDoDGQLgjWSwrrYtPFV4P
Ij5An1YbT+zkgWWEGeE71npP3yvL/MJMYu6i4HCsVK0rNZfDVSNWrJqX8vnMbl4/
4gVh7zbssIox5ahMvLY2mDorWTk430RfNIBRsM0XaT9FV2u7HwV3ZNaSff7yEMQW
YjPuNcJryc3UBAAGt+4rNqRaTbR/rYbaDo94DOdPz6ZW1azO6jSiCmmvura9HwzL
97kibjnQD4mdt2ft2angionIX2kdcVJ08767dqWq9yz7af9ggJ51jkLNEqVR7JIl
kEdbB167UroFhxkPnOvxa3CMkCXQA0UklSXBpoHufOZ5MAkQ7PdAQa+D+WUDhIdA
JzOrfRjgAxE28ZGgPUP6wABvinLDrETzeG4TL3vR8/qa8Yjx3j1p7OXJH8ZPCqTL
LK2AM45H0vVkzZGFFSaCG5AZ+WH8jh/AsQFp4BJAknHWNkGCSDWD+scGVzHmSwNk
J/oPVfMfvq96WYhQrzZDqMSWEgSn09yvnIGQnxTSTtINdSXOh6oT8zCgWX0YttLZ
CtMyXME888lFaHGhkc2pljCFmLinJY/5NgHsSMS++xFMcMfiMASHEL4tUyYimiro
LJGlQB1H8RJ/pNYpajHolc1Ev3hXL+ZtzHp1w9fuk0NGqo7sVdi2vQXzwGpTv8fN
75Y214J+eqC3/9Nr2TSEt0lIdKPsaSw3VvqBdAejtD5Phzi/lxqYH44ZNbZ8cFBG
rFmcRtu4+2E2OZh0tDiJHaxB+muQZOE7ncuM79ztERBDwQOC/9l24PKrkykw3aow
FDYPBWA0z2JTQol8sZRPmz700V/6+7EGTCwYLybDYPjRgmsXTN14yst1KMrfYzI0
JP1JJG3XJUuNZ1hz5yTVUt0wzyD2rsaJ3QYrrNKnAaiLTfR6XZD6+7vgDWOOKVk0
r0/e4Z85RlfcvnbevHX9aNJHrOAHID70rr6FRyANL3rHLhaDkJDvdOGhmEej9pT4
Keq+lgR6V2fSsMHvJuAlE912sHd62R7n3gaa3vynrqS9xyVhLBdwzDKQojosQLlX
kFRFr8WPKpN9fRMjLyRCVQnvZp387AUPVBeIiGI/OBrCiE1gCCZ6KGKeHBSoKlvL
vClloF+UHRHBGQPcqHGn20fz30l4erGw3H2RuIgz9eKYXQnd6zwplYW+HCYbNZvI
Wuy1EBs5SBKv7BCKhd8+KzZiZTjr0zGtM8tctux7dabRVZhi1RliMOjFNBuR552r
6KVXgMGP1etK2tH36k0Rn3nRDs3xevSvhkg33++JbThDSp7HZrWcHwBBc9o8AvHt
AStnyb8BIElMl0GXd8bniled1l2vdpDBB8h+y9dutuO7t595K3XF/iVfbBo2ALc9
2Ewkcg9r/s1viuSJ7E71EBSj/ArBks/06FO/TQBXvPuXHcgSQEg0GKrjIxxKK/LA
mZSUBtbkKJK9CN2B5hngO3w23O0M3ukNPYRinjzNYI1r6GE0KxheKFC6AmyVARDL
0HonYULaih/jnnsYtQPFEhtTbm5ZlAy9Ehy8HB+YCpciUuFzYFKB2wyXEhA9SMpW
LWKGHTES1k4oqoopdC4SdeUp/asfrdbivBpLRhZJpRlVTwZf9UM2IBf1llRGMPq+
74JvRj8c4s2Y+tNdIDN42PvAtkhY9fF4mPqkdBumbwYF3rmxawaUM9o5bKX9A6s9
Lg6zaLFs1LiPJUgQsalDdAwIcC4N/wEHF50IRk52NS/lSpfsGlO6lkobLUp7Mqcn
9/iT7vzUW2VB06poGxCcbYTKKjKL8nHESRs/FKmPL98/o9Yefoh7sM2vL0mBd317
u5AdJELlmFCEsHdyN9PIBMn7i7NIHhsXa/xNsI7/d3WJFPeMcADd+lhPyOwyVk+p
Iqdr4Ud/o7VyzEWv33qwwLUv+pHaZaxST4eIgcuPlEnUU6m8OjbhYxitmjtsBENI
L5pQa7KvbbsZRApgsbaiN0HXhttL9oHk/qrMsBn+8FvyuOi3Qs+U70iUojoVpZt6
OzPlNpb1TCIb3ETHuPFRyvjT1AIMaGnsHbpyWfmwlYbyGTo2KvZYiRS86GwcmYc8
yp+HkV6o9HIAmWI8gWn20siH1PTNfLJ31Y60dYUIxrU6m1j2IAf6ZNRLQYwxo5kW
lEpLT3cJS3t/EyZhOZ7jVf6YRpmgOFCv++N/p4e14Grp/g3DmkjlpjxZ6M5J6jqH
xNIYwC74uJGdT1n8RCvv7dxiq7yGUwLPIBEmIkEynwpZM7oWCZXFqUqPk9KUONbe
9O8MrJM9Bbav+xK1iv23/MD1tl+ek4NfwPkisK3qubyuv1sSVqcxDix3UwhxOJy+
cIX751LsSCd6jQ2r9m9YJ0LT6WoP0a9uz2pX9wXYsmUH1T0httTDn5maVi1z1SMJ
r+ekdhgpiQt9VjOXwdU5mlBaA4skSWo2GT55pFWJoM8HvgW+KsE/nd5SU2FoPYZi
PnVFXzeI6vY/86mxbGrbceeAX8vlSNGLrGpGaELaJNJdhSi7FjkVnZs7XDVQoF0Y
k732f38veCeWo2UOQ9UCY3uhfz+HlL1WDq6ZHut78RqYYyt6NMw4WwtNWw6HTEur
uR+t8+C0OEeYhKAh1xvYsPYo8n7yjBRcmBHCNxLYCUTX4JZIFsq9T4evvrlNX4xW
jEBggqbxbuPs4ED/0HVhFCC5HTBhxonFR4/1b/O2+Wb8tpmLqQKeKR9kowoeslQs
adtlIYwepy6c1tBzHBXEay/acKd4Zp2N2w1gLeBORbOYzPqL+H8LK7x6zWF5cPpr
RfIjV18EOSvSAqyTzIvIsnldMpSCZ6qYGiBAxrtyTt52/oiZpF4+NpkUOT31t27D
Pf/NrK/6klWUn6Zw1L07txuPJIVtA+yyqqU1bXpMLsSKkMhrmElr9IwcosZDwIVF
lK/u2XET2qFiUuOV5WQRgHvu+TLEbGpLpwaSYHVEOdZsjhHKdFBGvcVWa6UIBtQa
pYoVd+AcfyR8/7fq38vOpfoEUqj+pDRdOBS4SRVtuJf5WC6fsPLnz+23NvsSUZ0z
DLL8DOGfIMJbawUhlNpflcAOzY8vlYxG3rP8m/9XSDxNZ7dSwhD73YA/mwe76aGy
OJG6osyNBlYmkPkVr4l879alBtl8cMr8P6ijOh+Fr9z3WlojBVHxu0u+yTXIjIRn
QoZfvl3QyZoTbBADwb441BxE5MAAGC6SC4sYT6zFNxD7RsotUjvPfzgDLkR/9+Ss
zMCp1dsIOOiP2sy27+1Ii0d76/g8a1BW6cehXCrp55B8+YT0ATklvUVmypNNeuDU
ChLOsGHxLuAz2l4zRXZCZqi+5FUK0AwQEQITek3COhtGxEBIFaHGGpCsipPoJJhe
10BQ0BXT3d7+gFFunMit+YUKJLvruHc3ZHRLixuQxStWR2AGA9pr4VLQzCPHwmbw
iyVVif5KggawGxMK9wg5Zte4QOgfVlIn5axZPPHRrUFBKLn9zUAXVXwICPZ5opcv
ISR1kXqruC/DJaKNgjy2ATmtKzIvQaxEqIiS3p6llcXlWbhrmGVhYPW10fGu2EUK
t25OXj2y5WlnupQkd593Jl+92mNV/+InT9sCzLcM1nl+00Tv9zspPw2G+WhT5w9k
P/5Rl03ewut7OAlZFE/SvN/zXK346PJtNjE9SlPtIVsgYe9QZ5fYh9QYfNoTPgTG
fYZmdfBq4w3QJcJD6SfgGnMz5ELGLAu/epFTlkHtAnH4efrfI3IeHfpKZUNdvbB0
r+gcQPeeAmEXrEaRow2Y8iz/udcBg8+7DB7rGwaUwSWThsopON61+npc5PlTT5LU
F0qQE4FFmY36rxG3mQib8DBsUl+UfBDcC6/9AAxgVuJm7EOMoIGZ7QKle4DeyBdJ
gbYqZtXAi+qUwYhAM67Hdd/EDt6STdP4eaRE9825ISUTngANkGgAtMAnoDTi7ejM
U2p5YDFkQ7ujanT7YDyFmOJSfXHmY3qmSnmZ6I2fS14Dv7D44CY8gchNv1/6Fksp
r8TeEBTg7QlMqAF3pMWAKBxKI3/m4s+58j0RTclVAPGJlfYhFs/s+zdQSzaw/pIN
tWpqxM9KeUjrmaFFyGmhGEGP6YCFqRL7+qKUNtfHyWtRGyknDGT0o2B1E/GbOIpn
zkCjgmcg+A/Fn0Wf/Uhf5d6ccLl4MmbjqLmK0TetzH35p18qD2lelrkp+Kpn71vx
RGdJt0WEMsTm869p3/kxEnIndCIi3I70K+lr6WqQ2PiXb7U20wKT6i1GmrJjKI7G
E02VgCs0xUMKsz0Y0qvUTtsda/+vjjYDJINNe0vpBNT36TYJ/oPx9epW7HNT2BKe
edrIH5Kzi0NxBiBAr9b/oZzHuskWYnjJUkYmUYkDFZqUwo170oAW5FYqn59H8yeX
UZvWfgPWaz1kXR0S6+nXelWXVSWUDouWb2gXTlewMqo3E2ofrL6Zq8zpZLmQT61n
XDzFp4YKV5niaKNE1rn9PU1nTm8Q7meHYWcfANPuTfaNeqy7URdm8ZiQImKVRB0u
XXeMbpXNpcF38qioY/MA5g==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
MV/B9WgASpfXtQOE7JBhKvu/6Ej5CnfVCBl97J8f/wpbLY7QsNrxrmC1relpKaYM
w4KGWQVaTrT+ZogjjF4pIr+B/blvOonF0wWtVCCnUjGUXf7Ff3JZpgZVafSspIpc
oIuBZChkPfmAGaDsbpH/eoAWoiHq8uDd9GJ/56s3TAISJhv9899VX2OiFu+Sr7GO
E5EnXuFk7MfwuRmRV/7LXVn9FgpnDyflHEwwp6I78pLmW+VW35h1XzLO5jHr5xcY
JO8xVSFnyJitjpS8o4C5aoGW9fYHz/LhdUKpM+QylDMXdYThezVmbLJuR9dHz6um
2gU5bL/859pDYcjfa/tDlw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 23728 )
`pragma protect data_block
kEpL8+1+rUgqAYVbb3i7oYziLQH6DyGC9riRwAjisNDCiq740ySHQxEmlEw29QWs
++5qZ/lDgLRK470fpoZj5hctpwaC9rMqIcf55w8ND88LofVZZHGQdhiukD4ZINSN
WgTJwqN3tIq8m8JnLT2hfsqVGAR4q5Mc0bIGN1rmwsT7opEIspRM7wlwwEGxPn2p
l1iR8zNivezZZ1bjlPS5kMe4P0M4joWwCffE1TdNtUoG70DS+dujWqdIN8Ef1Mvq
Mby1CPi/1a9pL7B0S1xtXWARq/E/UyJhv4+wolQQDcU5414DpyTyAX2wMb4IM4BD
oeO2n4WqHvcrM8Vd8VAP8lPSsm/s+M9/t+uM2XKBYe0zGEUx9yC5czWYBjOyD+Gl
kjYpFSKW1zSF/IKrUJE34Rjt1y1hy0I8PIZQ567ik0P0e/L3Dm6uSp55PgqBfowb
q0LtGs96yiJxmcDQLbq/+IhYn4naBZG3gsLdURVGzTnAxom3k1YPdeYs5n37NvJF
/wmzDj0MlWnnARVZDWOaxTAaFsNE/XgfPw5GX9JGakeD+6Ihrex8B+gPXygT1w5R
HKvInrDeVeMoopJxm57IQEFkJTzhacH3xpcqUWtzwCLUoPgHwZ1o/zSWnK+sYp1I
nRK1zf9+o27BVmD2HZeKMJI3Mh2zldCzYQO/UxaPhlR/hEjQ+lAGFkcKJxnUXcQQ
X9hL1jzUGFurGRrIUPbB2um0c7cDVIATM7HlmMn3XcAyErDzq96tY18HBkluX2Lz
lrfF3otEwqlNp9VNNLHvSOVklv7rpXdYLDLphe5w5OHxaQKBt5gXMAxyDAkw3REU
IOKyVn1YPeTcmkuIUzKNr+5BhmxGIXlNpNboRyXkhPIvWFUjzitk0Pr88LMMh5Ci
cnREKm5zO7N6MxJbX0JBN8DuVGk3VQ+TvPbpTzRHz1lwpNPaIEtFc5y5m/nnFxMx
iXUA5yScxp55Gr3l+uxGneZFRGd0SaRJ4T9RQlC8WKeEVIazvwJrAW7sQdzdc9TJ
btJohl3IG+RWs25vLUc2bYkTMUoWsnKtL/f8226aDncU1EZYcPtL/dzOrAvYBLFV
uJyFv9oZIkSrrlKIoG8WEPt7bfOzFN0c4eZQWUpGb4JiUeY9CEM7fs/HYt7qJ2gn
LHGouRmGl6IObk3ccUhVCfM8gimEjXf0I6b2G2xcuHei9iPvmjXBdXSqFyM3Laj8
hLG8d8WdOkybkEai3dSadsmQmCZawiZ2brNIa6OR+FP7mlk1nICEzxR6ZWFkAXp/
8Ad+HnJ7p8xKsAWgBgKauXMBQywwaUV7d+6xgSv3okE/DeoBsHgok6jFTEpJzw/a
RxngLU8kTATHtwBjD+PrZBkr6NAY4iqdyr7t+nPhCrFlqgbFtC70rjV55gDFCLKp
FN/fde1MhtFj2LiK2g+3YWXM+OBo8Y0SbL95xhgk84p6JKcSVTPkCszUBtpU2ntu
FCNpX/YDXFassnqIy/9maX100PZEae3YPX07eb7ItRwD3J9zztnpGzJ1XG/WuzXg
hAAfOYhZaCGaHQ7t6+zejPTvzQZqJR+fyY29I5onNjlnQ10Iozrcurc/lSLWPgSp
y/3nUHfql9tyqU/4i9XuTwsNsao1+2hhUEpurRA9waMNM4h0N6+6ugft5aU8A3bg
Fj5B7Ir+PlFsINGyAIeq/U/gQ+A5OTN3FoCXUPFzUnaxsFEqpHcZRTX5jKl7TYOb
HL3ZsdBbqboliXr7q+YX52+fCeELggwNOPbvObWqt8hUqAxlEH3MDkCF3DixVl5l
MK0gkojGh7/JEcj6VXTz/M+swGoWXV9i9j8jWhIsQ2EpyO3f5hmdRKqmZuRatMoh
xc/XCO5bXBMttCERG0VXJ31+XmQFmb+PCdR5MLvGqvLx7tiwG1OYVvRt6S1Q/z5F
PQ0XyX5w8AeYZvN29mpIEqc93bapbx8ovrDdGNJCJgsFZ46MUwrYryAnsHxyStq9
tpY34rltawniom3bzPWDvBdLxfueD2GjDH1bHU19Q1KbWtK3Sq4Vk/Rkz2bO3ADt
nHeEYKzHNyqvIlyj0XdV5hi1TD2xEZ4cPBraW0MLIXuSRrt/nZXcNRzLukUyvn8r
cPdiG4GudQiRLsVBozbrHi9GucVZLI8uV5YUvc0wP1TtOv20lDDVFZvcXe+Xfht9
UuNXm/x//cPVlTgf1SGRkaIYm1tVSLp8pqsAg3Bet/vxXYr+pzZ7DgvBlwixpZDC
K1J9jkhDO7sFbmDLz6ojU0vskOPCPYEmL/Tk4Xtzc85QpCbl4v+DXRhj3yzrkjSN
89pryJxbTXYrNWjaOWsqTnvUclMhGfBiyPoYnHO7/BuCGualKw1YxBuXENiAx/JR
Pys25BQBL9v39zMooF7tgiYV+CiUM0AjaX+bYyZyQ5lwSoORok9KrPweDHP0aRXy
MBGA4Iy8Fg4VRF0sr8mPF7NqxjL4VHYBaDRQelVlYAL7oqDiDk1N80yp3so040Mt
aksY1JqQTlpKkNKkseNIM1nrsAF03/LlfBD7Kwgfs4r/91I6qdpL8oyGGKUgA2hr
dhT9SmjWsL6/Bc5Hg8HPLEKAofQC2bjO/QzuO/Q39b1x7rKsUbN3rJNx0iNNnVGJ
BPxm9eLm9fyxdY3hLsN1JfjnGMJN8uIavEh//dLQKQgGZjIWuEPscJ6ZBFQzkGHg
gpJh4XUIva85zkpETbVFlGpmV1TxXjjpe6sKgTh8D06GmDrUOUunazjvQPavN6Fj
0H8YCHEcLuKQgylgww5ZFpOEtQtS/wz02ZGLvkQPpVkB6L0nFAlT34uZCRBTQm2Z
G4vBNFIsUzOCbqw92yFQhYzf8nj3EEKAzu84C1KeLbyE/D6Ozdceg92930mIeRGr
bmBAbuiszmH2e97H2eH/A3WmoLMfBGNvAqPRd++bRTM0enmWjoxbIjU7VOEcXQV3
+KeBHZm24MiimT4fWNdURg82mwyEzsSV8h/VX4JCCV11Bu7ke07hZGJ9G47DJ80c
clvTQXebm4D1tof1u6F4Agxc624EJdIN5pGH9RD6dzLhHBJZUNxXeeCklW+rLQfd
CaquC60/fUC/72o10qIUBVNTSsjDNeB+c33GOr20/ALKuDXuOJpU9KCuKamJaokW
hnMn4f1Ws1zu/mELMBhMziBrq8b3VnQwUjsHIhMCtnqEHrl6u+Cr0/XyszvBSs+/
F/oun28YuCx+jrLvaTTrUNzlgF898Rfwuhg87X0nRU18D4Yf3f0KTmDM73ha2VUu
DIwwcPfVnyuXNVCUHdey4st4koKkkrE/79JSvxKMQhSLqNE3tff77WTKXYdJcJGe
k4JMFgE0b4m0Ov2usudU/LdjqMY1kjg59T9G1PiRse7TEDscQ4uod9oEIXEsHw5r
WIwlkTyauroDNEX76ppohHnXhAv36n/v7xgZqyAQNZpnOeoQekccDAqmRdCdWbT/
ScVES5vokd/SCzQJaZjP77MBzbQ59NA6uOQSUWFswKBxLhQXc46HcDMwQojM9zj2
9yyC2tO5ngUND6FGBPucHG8o/UsrwQ8fbwEyg1pAst+Nlo404Fkayh0FjYMGXKQE
OEqyyAck6eHwf8P5Jp9AjzsYUvdmIZDJ1pjpg5LEzRFZyzbl5MWcE10EfoNfy2Ud
nMVX50pMnF5t90BFq+ZgbwDR1/NaHynuAhAtnWREbcssYlawYZTh9WnZyUz153pg
bBaO5a7btRbynJxCF3XdEiX6XRgB4iF8CoyfLsv5NnqvzRJqg8lWJmvvnGLPGU4r
zqPhhkLR6Zj/kDxlyebh4X4hTPFGEKNfN+EQCiJcG2rmvNSgSoeb9Vp+hLFAGYlL
f7hYoru9tel/YEZujQBD3ttPKMdsRoLV98sjjfseQuZMJ0fQ+SU1MC/Imu+++u1Y
bMMFNlrZ+ur8yGfQ601qfqTS72tEHyLCk3W5KPR6U45wMinLSihHWsV2iq6yoF9y
hJY2xi08X6T/C1y/y39iAF8drZxTPFhdXRlGN4cnSZ+sSJo1UFQYAVmdBg2aBmSW
tspcMLHYr0OBepqO+vRzU9rfQMCD3j/CbeCunA+PMlXRqRF0AElk73d0lufh/fic
LZpqE+rjfTtzrZoQM8ZA22gefevO3i/8VUZayhBNyLRDfFowJXmXZAA+dJ+110Om
jfhiJDEixigJ3L+vv1q9ti0fcBh0ubV+NbSWr844B25l+aq1N3lZNQGR9O8Fke0B
BpEiF3Q9URGBrAhs6FPiA1RDFdJhJTaOTRW6LINg/uApey2nsldB9zTTTlpaVXv9
NcGo+yQS+2/gCHdDQOlcA99Mqq4zzwLBiZyBKeYLTYhAcfp14dcPOO5geHnFP+kb
1PbpV/U+iQTCcoKktLkyO2sa36U01rIEEzPGY3xHWJXNQJeoC48v2y78l5Kxkm+z
MjAFpLurExh3SxKnOX3x9LS6CDfIDbdaMU5PurZ+q6yLFaGZTFqU6zqSiAJ0uot5
fjWDjidumXXYPJfz4nZlhex2Td/lhvmBH/f3RhwKhtTGolt0LPdCNytjXyowS4Ye
IabUOMW7yHqlJszIgkOKao4XjCfdivW5JhnVFtXRus59Bu4YwjcNBq3tNSMK7slC
Lk4fk8v05U/1jyvE8rXt1+vNl1uI3kep0a35S2Uzprk06uytTIb2zoPA65n4WCyK
wWrtqmcQR1ZTEF87n2zRLoR8LeMOlTavDmVP0qTMvFCISgSHk76oUHAZOMNyitiE
/2JSIxIR8GYQpeMVjCPT4Jd5bAIkzQ95LtpVpNw7ShDAk059gu+/efYGgGUsYaZ0
QHxo4ziuJommZzdVS0sicFB9ZuvvyI3uK+xJj7UQJI9Kv8bNpn/Qz7XLbjymOfxg
Kw7LmIAM7+UcnDmnhiloGqdJE1YWW1bR8VzzpGwovDsgTEgdkTPTsDjj5GF171Xg
0MnTEX61MLYrpxNgO+wPlKnQGR6mxWloAUEsuh0juedmX+ijqDiviJr7xn4R6Ykd
tAvxVVzU4eL/5HK1E1jJmsaJVXqkh9LLVePfsgGVhLH9DQsDmK7ZIXv+VU00K5wO
UheqTdjWIXBs53PKV6fV7QtDB1x2fA+4QX2IhDW65XXewv6yOfwFZ+iEltI5cHkP
zJUZhFzmC5Z5c/RVB2n4GtrwUucJY9gVS53L1SENlpNZ7hN8aHZHlkwy1Yi7xD+3
FWb3YV38Ugjnjgj8W7IlrWMHjuEPpRWmwRlTcmVzHEORIVsXBdBgkrA2vIhmuTRY
TVE2w4XEFspHFWpV6wVbYth7bGfEUBVgcMCejsGuCOB1pzdSqFEe4b1H2uWATETM
tu3bRDO8gQQj/6KbCrdQL4MjkHPuC2RVkJZOImOHry6MNuo2EfTmdNS58Aol8dfz
uAHOu/ifsYdBL/Dy83cq7qjN0zeK7ENZ0Jr6W6CNUn2wokg/3jo1bGlhVZ/FbbTe
gRSSKlZNaRQU0yv6kQuHxLUGW+yhVM7jQWsSq3VcHHKhCMbybeykkTPpAWs/1iQ5
4QiLiK/HkDdFHevxQK1Ejogqc9h0FcLXKf5RF3sUnoUX6CXC20rXjp7YF2Gx2pr8
UT0+qx8GqYOfSOwfZou0nM7SIIjTSmrrtDzvcIkc0jwJwBBLMPO/zs4q7QM+vMSX
PzhW7KM0QxaSHuGFN1TtL3BemVHJQCGzjgqbyfKnHDb78PfwHXikkxK960E/Qi3U
sXXklAfzGsXAealjHhVyL4FypEQgjLjfrVFP4ht75aJ7/Lb2SBoAXDT9qsEsaE+L
vFoC+azO3ccTeZFydBQwogUBarabqasey1WHyCu+VVXoE+TcQL/n1nJiLbCOLJ9d
uL/cJTUA+QxdwbBw9lucyl5XtG1CxpjVzB3iz9yKspDM5MZPDFsaRjcJNWVYoMeb
4dBrwwtNMuPs5uHKWbBeOl/CQu1a12BY4lD1v+1W0mGgMGXifb147EGK08tBwSxk
yNdNRtzhhlyXLLSaG49aRnl/F+PCO7qCnIIWsZFFijFUzlqSuGssLEsGPUBu5eKf
WbPDqr0An6NKY/0HByHALAm2yr4mZUiL3UyfBmnMguhFqUF6ibWsJw/sQv4O5WyN
QV28t+XGfexa3M2MET2rLHCeCH5hfN6l02Ul6FA3IhjXNX7zz50j3zWZT0wmwXYc
XDEHzUTwa+lqjztKXALt4Fi0q7BcsvD62kwnGtB3dsmy15MU6lAXmb532qeyyV1y
ABPaN4O7XSlUJzu9e2dJiJF1csak3585Wfud/iUO0GO3+92M4GZWsEFJJjtHd0vW
pXeuA1EsRtk/8oy3HgN/pUG/Js927C/q6sRoayo4tCpokekuJ8IlNsqgAVttEHFY
3bn2m2KS0FRJu8MCA0KaPqiBL12G4AS8EYBo8HH2aQcYDYRgILs2woqaearcvv61
+wAP59L9kHKSUB+pGPLv+ZBBMstG4ntkZrsKmmLLI+wXjqQ+MWyJi5usWBAbYude
hhuCqDyWpvNM9PMZ9ooRf9BClDNCandLSe2JWX69X1RZYrx7NoY6cB+5lP3fLup+
/9vUFIjbntdo08XYVxgilwnn3/Pw6+yI1NMki7hiZu+5/sWpXE4/CCNCFI6mMpWr
A8fRj7ufYn00VtQ+Gm4mfLXr/EpKpcCDeWcjeM/+y82p5Hn5TUWpp2jJAGIe8cD9
Zuw9kKpZneoLNk6SxcBFrkHXKB1oznhB2Js85lpODCgH7BPlGv7Bcb23WgVFbKM7
CHk3MMqQdedfASOB2mLFqEUN7d1fkAoj0gx85b7dZEQr5CljmrNvS1renFIHEaWU
VVLJTh7SyjLMYr5V8OkF27sdUnY+Toyd6dN6vksGXzwjwqfMm7mXQWJJzJR40Kjj
cGScQj+UYFuyxl2q32mt75ip9l/CrIe6DXhBQNdlBoaQado5JjqNbRA4pnGs6vLt
WZ2yJLfT7UmVvThSWP4jLJsT4DIMZq2VwpAwh+l8na2/r6S+Sim+jFR3GEPkxo+I
NkGRmmEk1uH7N7SqQn+h3G3FRLkuGR3DQhoBVNmIDbSq5hsWUdmILBFvOTQAsPWD
Mj1KD/WxIrFYRuhbYj6FQjG11J734G+6AzPntp8hH95VA+hhc71zymLsel6jqr1b
riv4/EN8vipaaNmPPk9Lva4Is3plzBt7IZAn8JB1RoGTeD1WSTYd2guVB3Z3Oofa
EpPqKNGaeaOa6fuZ7PxClb56iZJKHJGT77/ppJel3/R+axAjWd6hRqQ/03Ccmzyc
xFBRAtNPIQu05TgJutiYNbP8dc1WIg58PBgcTeqfgwp4ew9DCtEbbU+MYP9vzsHs
unKvIchku8lO8FoJwGYfeCqv6EYfYcp3yNID288E6STJIl2tPLjCIjKQg10aPsLa
aMcSQ6dFjWBN+X0B7imZzufJYK31qKgQLoa5+JCzxlmYM5QH/vSCPuW1RjUHSgsD
FpuamYP8BtL0gfb5w3hcwfFRp/Rj4+9kQCnFNvM1XxCcOHjMP2UJXSoZz8PzA1D7
Hta4y9KfnVJDm0blqeG4Zv1tfttp4A3BLCPvPwoIKb/bxSfxcVkM8VvPYUWXBlKg
6em7zr4ntCIlWVEBjXZ/yjSkXkzeMyVVqpDlx+j9WFbp2TzSD8YVobTVJe1xGqvj
E9P/qROk47m2PXGZ7FsxANPCddzl9zcrcGPNqEVIwM/p7DFxeLqMES0l4ZMOSkUE
xuGlMeC6hJj9bYOdpS9rbQH0dSpLhEJG+Utb3VSpkrm5+Mm8VsdZH/xUJtswNwQX
1LQjZEuAJ80CXNP1jKum88ARVoKPn6sCQ3pr6Gs9xp1NvSsODpOKc9Yua9H/AP0B
EcLuceTRIAQpq/EAxFNoUcK/7zNnyqd2QNpQUNaxpKAnqSdrjQVcaR44FQI0XpbY
LqvQ/US2v+kMTJRgsBZhKRbSHgiODpBEhtNjJW1Vyo8DK8Bpc40XusvOdVZJ1SbR
SUwe/Vja0HVHz9L5mE0MgWU6Bihdn7RmIj5qqlAHC5LEAYlZEyQ4HpdtcX4CMc4m
oouJSa4ONrloJQ5kugDET7GUooJpx6vDqEAQimbJThXPVzM4y1T8nfMO0aBMix+P
MnkK6rt0fOOFJ0XPXyI14sWZBbZFLmW4X0uzHfbTubVx0an/07KYidXE6NzCH07k
R8cnSlgpckQn6jPG1kvnRvvPYQyBTQZ5mQ47k7tsHlzXUTkLxHezGqc+cawXO2dl
YPQN8lu1URRTgaEpK5ltG3Eo4orKe4nIE9ieP2Q/G5qPG9YSoWDt+R7hpsVpT000
6qttruWqNJvBbmqm+CHTJM5a/m/I8iTcHtvTU4i4r3cKtEKjeZci6UA7RWx31Qi5
M8qiOFa+LGgvRrtahoLtZMYjjvqVriHlYnbaY1MuGKOdvyP8Uh+Z65kgOqVrizSf
vrKdwmusEkNurPpNL0VrZky+sHLD676tfSjmJXInNak8RNM4vzDeP34ipH6Svb7y
rBLc3UAgTobm6bgv52E9XFf+NEdvh/nABfPUDyRBuG63pDIxcg713/0WYf7Gfnz/
TQqQhnVVrP620A9bG9PyD1yE5z1aH+lZVdZxZ610Gi5OttfuIRzWqJpIeBDkknBI
VEuY3lY6pV+zbQf+IuRQrrl7zoMraeKbYei30CUC3G5XB6Z/vmzp9KHLp7XgVsH+
PW6d1rTuyAAnbuo6+deC60MO78P2bQ8WMp3quDBytpyK+O5m45wrjXqlebRc3Fn+
eP/TnZ8dXeSQVGn2s1tq4JrenA5iU8CmK8fE4pbA0dmGZeSJJ2NBI+k5qQXcMPkP
5MIN2kdnaJj8I14oigNfRHBq17xKoVz+B0AMp4+htE1De8wMH8aK+vUlbsBDSjdE
DY1f3alUOvkaADiJsm3y8SOpaVY5WUQNU1o22JNya2W2jx2/467I21iUm0NROdDI
B34FpFEGViyDhTtM84FMqJvEKL1rN18OEvTQHJbx7O+OAmso7gq1hFYMr+/Jo4/s
BQE+9bqwQNwcUlVy2shUS5uIRqyxMVU6677SODOo+W/olsDI9ts+3HRI1VmKlOC+
i166Ra+EIskoKiCymfNAkOetRqh4LN9Wm4SO5UkIyUBhRdh+tMravty2cyXwXESb
v/oOyw4W6bp0ksBKWXvxkjPA1FAIWVWPnYQYti0+DorDyDa5Or6lPG75hzwMSdWK
ZXmVgKkfELoKhF0xcLqL9EDEoPH6KtV1WngGbXQXK9nHR9CXQaAYjEg3VZfjbMZW
uJpq0wSIBea++OM35+IHA1I6bP02tf9bA1YavZAUQuQAG1PXRLfYvEl50mD8tMNv
uAgZ/+6gV0Fkv8bfQ1zt9ej5rXwCZsvgygI5+W4rCIMEznuTfQrFYNVjOn5m8ze3
e4A0SVquM68UD5Mv7RNIHq5MwE7pLh7LFK/Iua7q1sZIpo4e30eL9puO9Lij1UxG
GM+7ouVx5QY1N37h2RZz15OPv0m/4gZZ4cZw5MvMCo5SWRBhCv/n5r99RN5bBjU+
HAroUgtzEl2w8zQQTd+X+6dXRSYMAMy9/OOg0r1KyZ3v6NKtcP28XxhV1HTS9crW
WA9sLtM6aqI1Wqg5P8ci4ZEF1b03OXpJ/rbH9zqfoKJ+PMcjfpZYCYejdgsJAtiL
C4Nk0YLLpIYZyNdVLJuJAwk9rP4hdjNcq+amNupqqUu1fWkiI/kl8B8LMpGPr1Iu
CnS+nXEjaIukLGaJZJgAf8kuBuMLIt5uiE+VBsuSMr3IIJqFOi42tZtfJo3id+RT
jMkJE9MI5dFQoAgvjpG8gSB1U3ywD3tKPhiq9rJvQowtRQR99FDVDtaCzCzy+OhC
UeRIpfz+gclRTTWvXSqapEGg6orfngss+bTj6Y86EqP+rVkH+sgCqYF437+lTUIH
0vi8S6uVoNtxPIkC2DCMYV9yXW98CmcJ+Eu310hM3gcYd1U5N63PWh/sueljaQ8w
lj2jxKQYWxNb4SEe/5ojYXfVNNCH9HJUZQ6/4smeReU6z52VUhRjn/K0s5KJACsT
Yavg6TekCUM9aFbE2ZU1ot38Wfo8crdjgi10ZfGvrqtS51Ob1UvAk4Iy7Jc6UMUW
jJx4dmqKngylGGcocVtfhAAPXKuovTFyTRJy46g7qY9XW4rNC7PmLqeJWPQc1XQ6
VDl8VU961wgCo2+VGzExr121sih5wqX7cZY9lYpyEXDRSgr08wSFK0qMLnb0N+aG
MWwk1SE0g2kzlryUaoV6XhXp6Tg3owX1UxFnpSoD9gmv6yr+KryiCBZxk0nkV0l8
cktCC5fGAbdEsQGfhGBRUoZKYCZ9BV/pWNab55ZF0x6YO0uNzNaDA0ijb3a6TYHY
4dHRQLMGGUYiyXX9+Z8u/qes/qZLBK0euvMtG4dmYipYPZO3+1wYVShGvFpR882r
9vyamLUDNe9uKgK1I+y+WTbc7ybvKUPCUP5wXuiSN6jr30vqR8XrfC4yqhvni0yS
RmYIauNKU4tTVNCYpRi86BBnCxH3y2PY5vNpTRpwtYDT6w6bJRhjA20SnDuJAStG
aFEOhotvXvQ4ljRDZnKWgKbpCm/P8QMn5sQc7dMXL+DFU834369wWjiuTUbgaPix
2o4hLNBeW8ZiLozb9vXoxvqSRxpvwUf9fVNgvsQVgH+swzh4ve6qnOifhUDRG3nx
CUXB4LjoVBSwzy7PsxgmohDwOP8XyMfMuDBQMAy4ZDOw7m9ujhscFkskNzsq2cws
NFZCLHr+cveXrKKbTyl7dHYe9blJw+sYSYoASG0mGkXzIJm0IZ4OjDkzcr44AE6U
GUiv/VBZFSR7LG569sLQCFimjv9xJm5S/UtH0i3GjDWZKR6KMXr6xWP/cFiApNH4
Tcyq7HH7v8mAjP2mvmv3pOja/oqc9fYuoTZF0Xl2ii94wTUdnq4sumXqosgY6cOC
jVaSDLOgFYCTEnbE6U2nmXX6uTZ+0pYq4eaTBLSouDklc5iJiZuiKIKS45UWef/i
Zn1oJhqM+XKkQzi/ztZql7v9J+VyvSJfxN+uljoRY/FG0XndFpWr25cmcNgUcbWY
5Sc5N7nk7aNGaYPcU+RBjU2CeASVGCj75SEXS14XLRx0xHpatryOcCUpC7IjFIM0
Qz8XDlX1uwFYVMtK1FWN9v82InNVYMbodi9+XCSxOxauXQD5YILbq4egRHBAna25
bJJFda41ajzc277bqanZe44vv6RXbwF+G83r8CRSR+BdFo0PWto/9IowJlZe+ciR
l8cLu/Gh+ZFOaiMdF3aGFptSHZ8MfrQkeEh1oi/A4koohQG4vDOyQH7htQOdxa0e
zZDzzH8iPt6TRIWHKrQ1kjL+9nST5VOY9Xtq72Q8tnY4wNTucbhmUXx1rrga1Ov/
d49wRnD26OCZFOgFv4TDuPcFelBem+yu6dNXDNXv4FAUR0pjZvF/hK/q/vF8UMXc
qektxYg+kmKkBZAW/Vv/n3hIdgn6069y09nPZluIT3t9Gqj+vVE25VYRgHbbPzOQ
Y7CdDck6NPAxTR3+kX24PoR1XzOReHQ2TtMGtQTkarILJtrQHN0U7wbPp62XfoKI
OKKerHyAHek3xcAyZAJyvC8krE/dCUylD4DrQemF/D4L2yjua6LM5CLu481faEPW
A7iKEkGhIgsBgBly5zk4//6I5EDxqtnFAWyy+aPtH6ol7hMD5GLXcfYh6jKAtxLp
l65+eDETmEoA4coQZb3jSoN5pAI5Cw9YGKV49jMrhJyy+56FDpg+Q7nOYFKlE5kn
rNlIZq/O+nsZXlUZNnNJf7ml9fTbPWGXg6ect6nynPu9vI3eVp44osVeYa1rRugP
D1+mSaMdhZRSUTiqXGgO65uVIXdU0sBe69K4vKy5UnR0vKPRSjDr9kjzGIhrWssB
snfRVf51arMMeDQy3vAawpSmwTC9T9uG+c0s/GE0NjmYcqrz7A+UZMe7SWxjv0+h
EA6bctYxsV5noA3X/UP6EhtG0KxIxGCs8hcqe7LUURD4wN8YwtgXg7QjBjhMIF3F
ZT7q8tQooqSfiXDgHj+iOVbgjGStX/2bJ72r2NxOZL2IvEJlFDIzW6giHShkz/WM
inoWOGEfL+ZPZk9MDXUu4Wo0AVnYuO4bcO4Z/7uoscpaCroPYRUQg+gLS6RLyEqT
D7GX9kTpnTglg222RHbdG4KFmniL7s5WA2Y44Fb61Ctv21SHTPSuM09iGUIDINrj
BJHhaZ35Z3uU5qnZcy6blt5DrtAEItxEFIWLuz9acnz4hjqdkNLvzce8612Bb6vA
yltSQPCu0HmiRhPPSGpMjQXA2eVKzGdIGQKT3Y4XaPJWzjZslsTbRfm9mDZMXkQz
47GJzgWNDHmuLBLynO7XRUodYTBxnozn9BJws4t5AR2UpVKe4AjnVQ9JUyLbcWfD
NQL3gxvg8buTJ22yQ+DE/5Fn0rKDWY7DWVEJyn26bM54gFRO2zsVfLUeW8YNSvLp
QWnbxbzDcVLgZGaFHU7XkyAWWxvgs3MNGalFlVk1b4jCEYEdS96dLbwd4Li6W4GR
NF+7C4P5GPKKbTvVfH54vMJxsW+uLPbU7m0iCoKcpBCyhIqNwG+kZO2aDSOEqBhU
6p/GBulxLcM4BnZWXPbxLxIQIOVyvjxE2kChhguQl4MYsNWHkd3EYbIQw0J4L8vd
kWzyCHD5eOWje14e991FSSEx6o2u9bjhxRY5wQbKX5pyOA0c2rTNzI0phw2gpTc9
r7f3yFwHi9wgxpU+MX3YbaJrxNrpPug+gUNVXzRrM5fXprmkjoniz+ytGqnIOoBS
rIeMnIPBbVm6oqGxzVMkSw5kOrmLnopkKl595V/Zjv182SIP+hahpD483Z+Hm4TW
P74GaVTykRKTB0VM+bbU/yf5/5vHgk7xK4nWVdBaGP+fRnpNBp9bZTkYpLYVKle1
ioSn8I1SshZ2UZsMgOGCxBOVXdymoqvyCcKBMu27ZHgrzgqjCwa4OQVDqIhggeXS
ZdJnb/1b5sEcESD/fwpSdxRzQOxJGN1mDedXmY76aKpLBI//oCm6bm8HHhu9sas6
r+TTayJvPlolRkIV+DSqi95nBNlUBRSnvWxo3tXNa0Ky4KNBQeuoBe9G/t0vZqs4
xSksy8pT8Ir2H2XVCl8K+OB1x2OO78Ta6Mings/VDUvvl74GJyIEBezz0vMTo9SZ
ZKJGRXQDqiSvjfRlsy1yvWFbOE6jRkab/mUMWg5wEpUKEFuoNdQzjMv0SHdOKDfI
ZMQDgu70M+SnvJVUvQk0SiXb7ArQ+Y7zk4bS67WubOAUj1uWY79IwsYJfBW+6hHL
pBes/u2t1pMLMhQc8WkNYkSdwOd9Bop3H4eS0pCZ3ex5cSXC09AsJwe1BLvihmID
V75M+lHitR+ByC2Jun2fu1r0eCxS2sCw2uNcluhFV/HtszOM7Dd8M8wtX1hSR0qk
SJWt5OAr2m3SDLjgf5kZv4gCaHjJEFAzVKfuVC1Z5PAIgD+eHKrfL8/Re0C80kQU
jhWZ0O359O8pPDnB1TIidkjI0GWV22+3p8MYgRvEzoVpn5wHAcbjEDhy66GaJrnX
yHMSCZtfAyziysMtbFRReGDWdcmzMZet1swLlpbnE9vvuoVRhWDiXtRm3nPZRu9M
VSoGimYRLbGXRgQCcawSPzLR9D72qvF3balXiP6BbnfOZlpn9tTU8ZFii6PgY0R/
lYMcmeJs+FusKygnF8S0aO05pGgTg/t6G3hAS2V+J+OcIQkEJYrZmh6fGcrewbcp
i9BD1h5g31TvDBv6kSZ0+LSqsZfGetY6eAlmIgBDFALkMeUoPDBaIywjluzfoVib
wPLUeToJ8mYizAg0kCN0rvPqkjEI13dta0/WYVLeEP2FFtIb0M6Fs96/xunHoNv6
Jt4H+nkatdReVexIPuIdIZtSF9AIwPFgKzhmj7oxKxkfGrHlaRvtY/5JU04gvnt7
GcqPtlZhvBAkvGjhn7PGVRBcf+ouH0cI8d7pXCHKE5xgLny9ZKCz/d4FSfCPNxuF
Wls39LQ3LsitozIP0q8dRoI4+B6EqmzXf2Milog3W6/KgwTKPi23RhQSY5uQ0D+6
u6ZI7x6eSfHdiNVyhcJz9XFxCgxylNdZieJSfL74miz9dR+6kPbXu30i3K24Hx2b
PE8sohUDaoaF1NKG2ZvPo6mIbuDN8GKEnQnlLJO/QiJsTbRb7Kysbt0SYYP1gOnm
vkH1SuL2ZoZWorgFInDqYJMQWeudCxk+iODcuoamTXv+0G1pSVk45+TL6Y7oZJIO
RkXwZMXCXJzQVeunh8NBAKFizYEU6jZipkO139M9woSkoKEWYdAPHOHz2632eKyF
/gXw0543lUbqlO8f7eZuShlvBJ5QdP2xApdIU9X+WKio/WsoyIEE39hMFR+rp6sm
EuPKQU8DPiJ52MRm7dNIfZ+mV9yvaSkjpXPZXlBrQNM9AitfUmPLbBW3O8zjuEBY
E0bnF56VAUigXCvoy6lMGq8LSuHgm5OzE56QH9lU4HQSsepfnTPz1KlBRWJRMs/q
rXywep9vQl6wXNVlPkYBaGeVTNzkhp64SAKvJ6DRpyaNT2B7QMYZuF4MOaAl7qR/
ziedlAv07HM78M3VSGUcFf5LbbZT4c1ddJ5g0KCoSWaSF1XEnN/oYfFsxmThAylY
uF2acjpeDUVm9V2tIqmdcPZIxEKkjMb6ii8nQ3KavnFzqLJ+EzfEgBgd40t/7RLi
x5xB+/rE3eB6E3my+H6XSLcxE1LDV3fuak5AblJV8oe0t1n7sTyRMhTsuaOedDJH
NHWSbf6M8VhdoEONhfOcEhsz3FQfmxp3yKyCbPHB96yfXMrly6oWuz9mkNoy24YP
ymAp8RSViE4xMBVyirSg7oUQKWehrOGTbv7Bzmluiegcl5NkaA//Db4Os1PnUcfq
fzZNKVPvibhD3vghrDOKLj1xg+dcgZ/wbP/lPw92ORidMhqSop8J5fLszDKTOnBI
VCYFokYhsyjI08VHDCia5URSRpm7zW2WTu+kePBpZK8CDoymafKEuAxu9xLjmSEM
+1qKgZLhxDSlZVCF5VGkbY3Vt+zSLg/Netz9OjdX07lJ522Um404nFcMfsmYu1c7
l5hQAG+h8snPHmEwnKZ0YrkE1yqtZtjehD5IkCclhYcRiQQHaAiKhD/5NZCsHwyn
aaesajEjaNsQCeZvMbDAK4PrUrj6GrerMWNtDnxynXfNAmEuP8wDYJiiXXNPzlg9
DGca20kxqe1goB86e2gLfwCLR4FT2RMn1wZd/93qo+Xoclepho0d/rIRhmvMlGyb
xUs+hiJNdr54qFukWEp8ljAW6ge7saO2C3+OM/aECW7RXi7C+CTqnUCekk1yZOxc
2DphAomba0bqZ2pNBiGghV14/5wbrZCdDueei+QUxjcd37KptpSsmGE6kql6WosQ
nDXN8e7JDigHudVxypRwpgcGklYzquaoBK8XnSUjvMhb/99lNYu5fzZiyUZUMJQf
V5I2+S0tPGYwt5w6QTpLo5L4+kx7RDd+7cbRTgph1uM8F92dsCjpWgsWBC5s2NUq
kfiJEPcZaAjp8H2OMr+23uW1kqEKOoZCcVaxtUOPC3KeG7S0YRJkeDn+KI4xLFX4
GCIoceCCckSp3XtYHW7I6PnpyS9k9pZRibeBGTUzMSpNrhEIBwatMwVDrJgR7Xh7
YfAl0bqN+yt8LeXwEnArzrnqSSzHBrkYUFomqt207RNLObP6v30PquB5QbduS/6J
g5Qx0HYP9unuCSgQb+027LawaTCTrtwvJJqJtBkP1npjFQhw/PcNixFarvdjkSGf
mbwBkN41Lqm0wTKzWIStvuJISGxTHAWTBAk9040XASUvHzXj3Yc0dijNZu0I01Wy
8Hml0vdY6KlsANe1NpGqf5Lleo+Bqhh/TD918J0o6ZA83ghAAZrK6HXCCcdEHfg9
w2vXyAsTnzLzSN7o18xEkR62HvB+BeaYTIFi/ps2CGEW4zyiDtGjQcLie1vNZ1PR
qJfaPIK+ALT2o5aPcjcHAL+RCdoZDUui6gU7Tz2TVY3fLLMISqtVVuwPMzJ+N5KN
jamQIZw6CsSudQUdrHYV7FNAt6aV6P9nrGAgcdrUhb5Blhgv6VaG8qlG643jBNMi
OyZw+EboV6PPeKJyUUWVjVDPbY0x/X4NOwf4SSybbuo80yqbvULQKX9G9vYYsQvS
cF5jz3ljjZDQAuBK+iGmoQJ944RkCXbRSnVzbBgcF26Ue6BOVeRp7kGufjKzf7ig
WjUQ/kIZe0hpZymzYC+CUcHtsDB6ySAsKp9v5nUhSO7LUoZWNOe+q6UZATB0rNMv
4lhPK4bMjIxB6qYlSg7QZdtERi9Gradb/TTHjdh9rktme+sgZzLiTX67VB1mVn3f
eyIamB2REkzamcWqXyZVMB4PN6WaPc2oolegqh126XWDG5i1K8RBy1jA/DtvJ4fx
VKAuznIwtdgvSZAUFoH4bvw6Gp/N3HLVA1bcrffyWzEFAsG9wyfLJsJIRFx+LXUk
MaaGxd167VFY96IDegdwtjM1USdFD1s2mkMekn8sTmYBl7E6bI/3KYTAWhugalfL
qMGMHFUalkdh8+uAkfPQ+BaCokFS8Q2YfcMQuCAtObBKrpsiUcWnovHyTEAtT8QQ
EAUFxZFhq+7OM9CBVeH7UbAIEz44OMDidiqvvCYJxfs9QBahC9OoucyyvTXnQFZQ
Cu6PPksMf2S6CX2KfR3EgJUcHjHYWXG19ZqnZIZHIl8wzTJNH0+9xjYc8esfEF/1
NmVT9YAFTyW8dtBAq+Oi5quFbAw5eCFn/uIS4qRR7l1M2hAWrZvcBWLwxmigcple
hPs+NGz6WDNeRVMrSEJLINZxGzAQHwpyoEvp8Q3bcIHbDiQtVQ10Y1woPs6dtqwB
tnPK46OdeNO3zz4t+M2f1NP212s1A9Ff+nOdhUxl3jpX0klMZrqIQOJqnP4PMFpt
u9N3L8Mr8p6ucLFxWnbjPYsyLf33+L3x8S1mXwEigfoPth71V65VK6foN7eq35lw
EntQRPPF3/07OSwblQqtrQUSOQNMlggpYrcD392aAdT0cJD5sXpSCEWFkVNZrXye
TdQQfoJuH1VlajasWHxTU0OSBiOMbo6eVt25+A2XbF02R5wjcdC2eTBfwL+mnc6r
NrGs/+bJedj/+AX1iNpesKO1OKfDx/0GMWWn+zrfM4sg59yCE9psVnsX+obeXHEM
8WA3S7IFW5iqOAOLhiFP8KONnNhxXmMFX4fa9vd7lWryYz53D0Cf8ih8E5wI7by+
kqebAhBExEN706qcOz1TQFGD+vW0Xf3FR481krTKY07N2lKvNu41XtpGb5SXnmrv
7p+KFyYl/go1I8QzHgREEqd718HdeDXvlbMvY6Alk+uo/887twtDyQ9gNGRT0YsT
osu3D7lZ/x8DkrVisvRwy3pegL5FRZaVEFuBTeQuphTG3L7VlvgQ9rjfgnoaxalP
rmrvMEc8Mkn/T6K/EcmfkEZpsGz9MVn9EDxDGDALA7h1Zytj7u7D0xN4lncApUeH
0Cuq+ytUe1K+THr38FM4BIR8tW2/K8cv8HT41nFhvbsron9rTe4XuBRhdv3cvrtN
4L7bVuTC0wrmSeEy7qC+R+JiQUmQUr7Ury0gkH9GU3ek4xysVc/4nRCKTJ+OgQ0k
kqfY0j4+7JjAkEoycTutho6HS68shhO8zE2kAWf+WYkpRRv4an8tBvhy1DDzjWAv
/y2+KeirxOYuPAOJezNbnj/zwIMRP9EcPh8EFuANR7SU0OYJkvTSqbIcQceBL7OU
IgysL3UQgtsGcp09IjKWG21u/G9fEtzUSSQurvfgyr3Ig56wtZqHLlshBvZ5SfXQ
X7X3IZLDdfFnP55Mrujrssh0bbEYB7JQvKZGQL9cyI6ReICsokjmzvmhwOS0zHF8
r4CzXotCsgp1Xf6WTAwtXXgyhxVnirDbavK1KN6NusEZcaXEyDZ9SdrdN782wRuD
8tI68dnaeXbXJwKC6YCRVRW3P6uoUI8rJPC8YhjUkorukoHMxLFeDoXctgJsFkT1
e96lSmWQPTSQSEtTpVDrMTAmNVRsG/WVyK6PpSD3Xa6VWwWEGiZaXGatxqXgON7k
dStafHGT9f7rd/ZSIZnJVMxZk9WcUUxfEtsxrD8Tk0urW10eT5QxBJXMhM+NZIbs
euqgyBvgTbTv5MsQJ/V3rVw/7qgep+GD8S94sITcR+b2YXFVrl+4TsisSw6sa6BL
4L5kvGSFFt7Db3uoFDsx05ooPrmX+JQfmwG1YJc0yAOaSoEk+CGfGkhYi3hs30DP
efbWgjTsa7oeQ4IJ67mARUkZ0pkGFX5/EOPeX2IIydqEeW0hE0CWXbdvH798YTNf
E5zcouqclbJE4vLmUbhMookhDnR/1jcd1MDt+IBJr+hq/qtUK5a+3ia+1zO0hYVN
8hVTLGK5djc5yune2fS0ff1zW2wlcJ1KCv+G3ard8dkksV9n93bma0Am88kD/hl8
PpymbjYs/ZY8Xwb93l18/aqhURwwSw2IzcSRZ4Sxk+TwoZTLpf0JOpS574C7SRQx
jUPASeQF82JJ8LBARAurmYxppSi6lGcqUWMqmz3FTBZDnvOOr6Q5N8aR84knOeUL
drpLvz3VetIGdaxUMRQEkURh2rluV0xRxwC5dfugVAme/YqmRBvrxZoMJFQi7TTE
cu/fur+h2VcK+xlg2FHKLer/KuIvJm+Jz+c4sCN1hNClvNH+PSdfHKJCQ32l8gSd
b+ZgTnUV7HqegvtIS/BkVCWih2UIXZpGBv/0RLzdxrIoooTgKu2y9cTAaGX/QHd9
K+BObjts/8v2UT+u9qRxM676Fqkbj9OHmYR01gJPo11ujzTSZrX3eQUlxVlxNxsr
oNDHD6Tlz5RTwH8/QRhIE4e2O9c2aCZp5YPixOTaLP3fJVdttXjO/WJmjbKEp+6O
lVcHdB6LtRZ0gRN6syA7hnlTdu5ffUlr82GBkDsetLhAJZec10F6Jx9/pmTRmH5T
PArkH4VSJHff/CTiF9t7HYCswh1sbsw2b+QHfFNwdizn6XXEJHS3C53MM/2v8dVH
/3GX45GhSyeSzm2t5RVnybIp87oz0akAxVDN16Fm1tn327W0YQFSyg2AUObzNnEc
ascnPpmFXRQjg2l1PymwFyxA2f/hFshsXdlIxmYnoj3pDqmQreGdkrXkqNeXH/UG
Z0Sdw3IWGZnUkaXaLoeSytoXvXd24WTJFGHiwwTdjRS31X4f3ASGE0655WdT9oIX
T3BtzH9wD4LPpWX8CKR4AFa/SNXhrKC/MOJwH4BuigBIEeeH8XC+krFrT1cUIhy9
Fko/IE78Hje+NZxBdic4gcJgHhpsek9go7ob2WAMkIrWD4GB/EUj1sqhgUW8jobs
XtQBXivO1asy2fCACJTh+slztoixWX2+zNxSCO/WvgDV87bF6R0RAObPlttfBXLX
F8Hb0eqs6Zz6/rJugOU2b2/uiapCn8vDqPseEkaUOThwEqnxFdLoUpdRm3Y17hG7
TLZn9wY48yeZpCjQpC80Yhi/CaO6GwmZNUmIupwYRg+eAShvPhOlj8xEF94mlrrI
kjelGq9PIH2QlnvA8sKoB9f2FxJKOd+I0yhg0eMCHkFGfk10DMdOYWLHHFMk2Os1
fPrQqRpiZJgOOGJBsNTdTvEtVqyAbeE2yXFHLnRzlNi4zlT6IA/dYjmfASov8Old
EL8Xwi+ldC63XwnRrbu0siBf8Iu29uI9B8rjEkacdzyXzRHRM+4cFMP3HWNBVRnY
IGEf49CdOQwUeHudPBsUvY2oPtCezZ6809jYDz0Ir1uYpK8ws8j3+s4dJP6K2AEd
R8aTBlKeg86Klmgij2O73SHfR4/g5PnHFmEmEj0Cnk6qfec0R33NOBT/k+C+Kqqm
TuJ/3HOsh8oBIFgsaBZHT9SWcgstlsH6nsAlGlYL4PbVyR0SUNNMP7k9JzJXZG6Z
i/HZdfweqHN1WgU+8FkgfTffokL5D6gJu/8/BYckyhhB+L7P68P2ElkYJijnT6ks
eMHwhF8BNX/qhVM6cW4mMqn43C6UVhApvCSZiYbA2eQr110Fc3grzrU5kCmvbkf/
HpRsignPurSO5CEIm/A7t9lW48nqlkmcYp4LQR65gD6zYV16UTUB6VbC09nnfdFB
eMDudRe6ABBFiBeqlEoD48vsye3IgtV/MKGrTWYVextCJzYpJtq4x655du2TsOJH
itIpkJcP5tzNtCTLqF387MbGaQTCDBnAm18ieWLXYhHF16JxGNPlaDGX+bSrjZAQ
5e4DKw2H8DRTcmRXHKCvtyVG+0vyIOai7cCZq1+2OlyLkikWqs4Q08zagE/ic2Aa
AQxYLzSsWuVddZhQB6zFCt2B4JqMDbFprWvnbOWXVD7DYYDMBFH/GhsQ8R2plwmO
Q0N8JMSn0B0/ZDydn/L22XLSWgOJFYfZKdzRkXw08mobP37CXnJdrKg3T0fPIgSi
jI+O5Rfsuin0bOoQfyUeE0UIoIajHmPpcFU0RTeiSTCIcvTx5haOYfZ2NvZtFQTR
fPRz0dKuzu9+qzL+P4loO1NvTfeCCiJfUawBe1oQN2RLA1de7lVDi5q+geEFjtYx
Sa3YFT///3GMulCROERcQhLcJ0LDoyVlhTXdAKKaos9H9DWRuJ2Smw3kNhOEy/h1
7W9ho5tOjmbp0eHqVyE2X//Sjcu3IsC+fwnohmb4UT6iR8E/z+OgcUkl/gfvnAIO
87gxJv2bfyn1xf3inTI55LF/ZuNgJTDVOKY32yYrfy97jOIsalcNP4AwiMi71yi7
K2p0LW7VV2ZzBQHyrL2vCSwv1JorvCRvUDom9rGnz2zRS1fe8CujfpghJeUhYWAh
3LxPSh0UI4MHOm2f4OGbgBtBMXuszz1Xm0ZAHPDnDLKH3WLxp88yfvx/KIv0SLJP
YmUq7c6G7kbZXKgm/W8zvl+C38aN/zbsZ2iKk5W4iPBfuIXtISkX7aEOTCUmiHuJ
PJVX29QLwiFJ5EZPnwzUWTEULZh5t6Ijmz8Q4TdSnElVFTiNB44sw39e3yL2eCzw
WCfVkNYjuit73UiolvCos+4HXmoXP8LayQjdu04FKLHxu4qWr9K7H6eoHVXXf5oe
njrm6FdC39bB/FSgXwHe1WM5USiwluVWWVMLBcUCcog/4KnxczGtEFld16cHUhCq
v0Ic8x0Nu/EPwX0b0i18PafHDwG0tIb6zoatSq86FI7UtzFV7vdyDJe3aKThCPG3
916UIO+zNbr7oJDfGZeFurljkOaaE0NIIVIdt80NFqc2w2Elc2w+AAGbKTplb67y
qnRXl7BMXt6KG0d4ZKZAAqPefaIukRLRdvksNwe2Lrnzp5A7f3M2n2BGY9X+ziTP
pyldndo8xJ8rSthE5RACn/McIscCSqdGVTpy9SWergARdYPQ0gM55WO3IINAa5zO
imWzfHZ2UKTMgIbN8MAJZx9dNuTx6y6hyyyxTXCNFMOIWD1RpOFy6cIAdzloRP2b
1MDx+jeZrS9c+/IWibOi/ovw1g/rxJgfsmwt8cEIA7FiE6E8G+D5/qVBOeol+1ka
xer9WJBWQ5rvsvqw+ZVXeOMSEf5BnhL9CyasZG8YD9pDEnte0CsBspniZqP97Vme
91pKepGkiuywjrSnqVZeS46A+1dmg3OnV9aZX8GMDW7/TQNJOCQ52/u27/+J7tIL
zC2MSedsizqr/jg2Dt7FKxPYZ5Ak63yRYRQwvHLoXpBSpmnKkI4m7XYDpu80Yz+g
5ebcFGj7XuVfs57Iy/nJAFRvpdOuQJXLwQZZZVV9sWvK5auwk2zrCjBtYcAom1HP
QiE9r+XaR+a2qMqik5stZxWl+5UvAUAA7TYPzIwiZ/UM1DdQRWFy9qFzMIpXOAq3
+LWIeKAnTJcuSHvlWkWYBMNQ1W9ose9Z/6fn0ucy/UDKGoFFt7ICUz3lcU2bGTGS
Nhq08RxTok62kEni0SiMmHzI9MITNXXxV5q8KN+zG64Xq2x+Z7TgP56PQAQZu+0i
21Yu9EdGUTTArG9VAQX5TWdNTFBJX7vRlpPvNJR1W7QBTNVCTJCGwFER8LOL3KW+
8B0IfJlqspRT5RDCvcdYJEjqUtLvptN2+uexf9F6G8F+aufLeQ/j1pgVOqtHOjHE
Rgww4YKiq5VVHnIxnR9d0KROxbwJPNFnJvxmASsYa/vsdd7CewWXF7EGFpOXQK4c
CxQNsECf44sYQenX2un8tTF8LAU4KBv1ZTP/SSi2Go5kTlJlBDEgZ9TMius432nT
+Fx2XM3c16Y5lv9ThQxbVIkQSOfURq3sy4cVoNf0qYUpB8amePIljGnEU/loIE1q
R0iC1YzXZcmEvgQhSBID5G8FKzxX29T1BDHCEAYj7YzoavGW8h6P7kJVnJRFFU7V
0cjlBdUR2YLHP8CEWAM3RwKTqi8eBCP48FRVDqMH0nr1eV2+jJML0TRL/sBHCm0v
v+gc5ZcnhN5XyMEcnaktiJZxXxYttuNjq5MtdpoMzALdvkRNJLrl1MeG46MRoPry
AM2FR8d0QU/PywIFB7bxmUYsc7w6Fl4AP9CCeAGWU1QQnMSuQp6WNIePyhAB3kT/
EJtipcVZW8vF2Vg1ovJkLgvz6EOXgjU9H/gxEN6HXNH4J3zxYvzkXRnKcuKkV1Is
V1oSKsT+pwMpJDZrWYVEFA6be4ZrPzvoHu0JxnGdf9jgF7U90oSVVDWXmCABopdx
P5x2JFxWHILPHR3Rf0Rq0XoCVixL99v1JFIIE2IrDikYIC2jsoBsscVhBu3dBq4l
CLWA+JGlhrB1xvSUIKCm/VmsHW+c73Q5kiH3Cbsgqi0UvYMYky4gM3ICdqbEZ1SW
NqL5rtBXETlJvO3SJo+Jn1/9TVSeriLQBjkAixL9JB977QmfKaY7esM8QMhHRNsW
5LoFQ/UPD6vkjp9vvsCA5AGPJLg5LkG63vG7y+hVFXd+UzTYwa04/YMhMGTGeIjL
Y3JYC+RCiyi8mdBS00Yk9O5AzmjIfWYGl9FXLYtfbPoPY/bCinm2KunYknpSp+rF
PRmypY7LMjPbMN4akXPtBevmWPqSKCcEFK+U2dmrLNztHJsDkRBJWb2NRFGAvmAT
dvG+H6hvBNhsDZf2rVmByoQRX2LzzgcJQ00QNbxeQTT9YH3YB8rOX2W8VRg3PvMe
5/MZ6aRZERsJhZuZwt5GHjgWEmRFXeQEHqRxyuknRuwKRd8XJZv6uSvp/bqjWIdl
a257x0Avn3asGEqB6pl92DGmsYzjnzyD+YfgmqqNYVxrVUNd+37yifSlN9DzDrte
DhSAFXHcf2/V+82MWEe7DXps3/jQo+w+d0aTNWK/tj8xdE7kjNlguGvAUMNCSsYR
VJqj+zWQ9ECWIfDdLoITVZD+w1zzFXfrrxGTdMTfxV/9hw529KtV5mG638RHYR6b
CgwCdcdJ4IcoNL+XxSG37n8OIYq8H6koAcrYY5nXFdOnptSnL/2+NdTykYq+Yc7y
T6tzMs79/p34WK6/6KLusN9pc+8qw20lGkAd9He+BXJrgDhRf2m8GXoIjKSwItw/
PyOlJWJQggxC5iAjKTmUiORHg0wo921rigLxSvvTYp6MgZ/zYhH4j2RGN7BE7V43
zp8VkN4cPE4fuzVc7zE4IHg4cZU1y4F7l68saNBwki8BJ3weJyzSUwhcFhBti9Qu
qLwkIeRIi9r7Bmz4KMdWd4b8RAzfIMtduJKbp8/d3xTb5szlfvwEaWoXdi28mJev
jBphoUbx6AkO4bnpPnIIjQqFS3L2LgfTvXPxyPLPvGc10/hJAsq5X4QQaW4RdpOi
iZgB8TMfHBW4Tfuayy5h097jjVWiwGF0IRBGCuNMjVvKzGgToH5owUD1qnLjnO/4
y7MLbHy+o2v8OxRwqM3XfbVloVktG7tmm0JcrjDlBjsK/a6n7cY3vDjfdDCbbnQD
bpAucdVYGSqzsgEC1ArDjtY2hklMet+XqMk+vGu2N5ruBwmmVBUsU3pucN42PTFI
7TFGnSL1UEwFJHKN5r43Jj1ZYlsaBvHf0ZJo/7U1i2A+GZ2FyO/+whWaGIzlMExH
bB/jIWXshWCdty/OUAY5mXmbWVkCJO3sbNmTGogInRC5tkPr1hcWQiJREDPivavs
wOuhmM2+k1Zs/WkIq9E7+08gVB+CqMa5r2FyW7LxhtBTXdq2k3FNkIP+ol0Lnw+i
P9ZlDNdR52MoTKkbe4n5x4tCXAClMM1gM86Y8pdaZNsMqHFHmuzL0P4Gi3yuL99G
T4n06uyCzQN4IiqbrmtWCPoObKg9CmAXNGe1MGvHsK6/amSynv3U1kBerEC3Nsk8
SPQkEFGaIkNTCh3ZdliTziOQs1AWY79S3E3R1/pB7dSdsY7C4VjLmxctUVTfFB6O
5IV4O/Yb5DIsGGNQLn+4nUrpLKkUrsovge26cMp5+d3iZrJDk7VdJNwpHCWM3k2m
UNzRAgQ7uiHWMLh2JKA8NQ+GyllP0j4tQ9k/rPr114n4rPiyKbb80Q40w4mcG4Gu
G/qGei9lKr5uyfq82IOJS5TkGZN27NPZIo5K3Rg+XaE0eSCSARycGB3RfB+qmyNk
rlt8NSpWGTpjLHv4n1QQpxQ+DvmZuvg+QbHGLXV8xuz7G3vCw4LyXMGj/y1JFqt8
G64wO4/puWuGgGgYX8KLJ4vhUE/LVDuCgn55+5A4YsXA0FTFbpWc3lI/WtJ+4NKi
PHVUB/V2T3LAi+x6O5ur2Edp0WmtFmoAhhKvtIRMxz1pZEMV+DbZZS/maPAOIG32
GXyjgycxRzibhJjMQvoVLkd2KYKWGi8vEwk6S4yu3mErSJDoIYylndNikhkOn2kw
eg94aBgC9FeJpZ0mm+CVyvsqqq/S2s/8nEe6/W08xv+u3o9UexD/PHtaE1HktaLL
vIpy/T6H/oVgObUKLil+5LEcjDf571hjMI/HioITtbKied6h9KXB9CLR3nLapRt9
P8sGB6SI+0Cs67PrbHFLMOLQ2Q/N3iiZdhanR0bDOQsSF2LhMLdOb0r9LrXJ5ShC
GWzQz3s6Fsu2JTIAAVcFDpNH+AuL+w70fyQq1RGKLdE1ND2YG/eTuf/8ogUo4qRI
KYRptMHdYH9dYvOrN15rVOwp0BYRzLuL+WizdyQ5OOSVOi0gd1oYD3p2PyHLPAph
3dww2i1r+tTuMh66lF3XN7LD7rof/QpuWPIrNHsQloRs9EughOTB5Rn9ekFlGmFf
uhgzoqrt9Fwc0SmQDjTqfAPNl/dk+lm3xiQjjPNExdpcVRSsNW/yeVZaDBccDHYA
g4zjSCzJpnU79bLh074OiS/w8ipLot6E6hyn9ZXlnLyZalTE8o1Yxl06GRu9dUUV
j1SwSuIlJ2ntsdbuUg6Wz+56F8dimH88xHEM92WPwIld9sajPHM17+idRuZvzgbR
7Y1lYV5WJlYZoeUHrfHjiPaA87pS5NLts5LqTZevwEpQA9qojRlkVqrDN+n/Mq7d
p5K0di2jYLtXbdeInnubilC6j/tNp1LyfXGsIGjFB+aFUFOj9KN8ndnBLPwEpf5o
6+ZlNbua0yBO+dxwWe7Qfa1uLOtE5iYngsxzCEb/poVDgJwlhHpcUUCf+6TMp99q
XHzH0BGwcxlOfjQ6uQ1Xhh0CR47hwvkZbUSRwKBJnAG3LZoCzRmKqUKTyzrluss9
c0YySnLTVKZIFk3wU3rO8I5LOOL9Vo2vC11xPSM5oSEZKxEIWftwQ3EdtEeNEZe8
NvMIIPJsR3y2u8DRYEJ0Vg1AJmy4gPglt4leuXof3t6BMdIb2MeNI1NKSfMwfEu9
Ki2mHG2DbR6xiLKdH+gSxE+ugDCe66DatOrbwAWFtshRFwbm5fT/ySHVzhVFmSMJ
tZLG85sKk1TDcVkL32i2wRpMBz0pcRGuMZ+AyW1IJprb/Vj8iz4eUpfjT+JpSqcv
slWzJe0nMtz4MZ8S84S1xLdSrQrMKOU7Kc6yIm28JXIk2L39jNciJYa70+RfMc2P
4YlpIR6SuYkq2hxbZt61NTcE1IH+mAV877tgCtPGnkulhkGe/Bv4Bw4iraI3ojap
Z93LbiR4hXJXIk3aa7TsY9jKRvKLHKnD24l9LhpQa4/sd+jOWHznKIlHcOzcvQlC
Nrm2K0bpr9uax+mMK9cfNC1ZvJ3x8UvEoGNrthycLjunYflrZmQX6xJsQeyCAbKJ
r2iKmP2pcwiitmKOyv6dpjODHOGKisWnOaA4xlDc4qlwsccxruV1IQvoOWR5Yi+3
NAkuLrxBub2o1hwSLRo0c3AvBJEvRrM7uFWneHJyiw40k3jFUNSXTHD5+iYDZwWm
cY8V0JXtrSYIOWevQP3tn3di30Iik/frBxbkpl36eUIDPQlaJpQQFSZ3IZhMHlMV
J8lj0rjBOz9c0G3l6KqttRiDs+7fDnlHA9rlw5yp/rk/gdv5jP8ZFHwdE1R3Iynu
gWYBadzfDeOcASg87lyUtwrVddk+oG4H2xAGAt3mMS090hbFR58YWUNCoV0syUvY
TjQ1TA8jrWkVH3FZPkGrCLD8Dq9436P/Rqsbesj1jAO2tI7HO+idoCZivrHjTCEM
ooCC82B1y84eTmLpqMeUwvYihkHG/5XNTH5PQR5MwHcgPb4wP7Tzv1lsGa4NxaIM
KqTkHUH4H7G8Aq18yTo/KJy6/k29iSxLEr4zOEuekQlDPpa0e6Pg45/Zvx3CI60x
TcGmWsMZ/h5epJqYC3AwyN+jWKGAxWzaI1A1L7zuMHs2a6tP+GPATkCX58IaRul/
XbQQqHnf4a1J20YRnIYH0MlF8lX75kvEFGrgnWYcdFVWHokl/VUdUpL/C12RUD6v
cXsTUZyzjiNTf+ZkK7GNJe7oEWCGP/xDZMFSfxHU9mae0lftLoSYFLn7OoQqa2m8
5TvnyqQBSTObF19NbR9y5TjZzgJZhh6PkzZqG3Hy0J2VKPifeq/K5MltyJQOIGk/
Gvr5C+MDgTRr3Xjv8uGevNOReji+7UL5KmFps455saV3MRduXVitNWcqAQ4pKQ0Y
aJ7mxCK5E+ZtwIFx9kYHjWceXMaC4jqsSZj0xXMeVrevSSq07yr53ZtmrqWhp7UV
ICeMTYdo6VPjFB7OE6gg5K8ZDAFqZvlKkyel/aYuW2h8UZygoJh5/285Qh2qYWwT
FZtuhZ/ke6HqdqY6oLxMPzcUN/CiFP0pvklCBN7ApQ+lsQGbUoQ7AZgrTCGiEipH
pJVS5/SZIlZgtY7xWpMZv50TGI6sBIoLo7l4tchABffSJyoQNCKZIMrfxO0h4Bee
oj4W4GpdaARke7Oel3XXqtliIXCO6rnuz8pZ2KArGfEpX1kGn4DHbbfjsYc+vMU4
Q97v69uN5m8V6HCEgFXqFuD12Sek2s1rrD9jz9e/rYDnzC/d+JMnkB98Lh6WrO62
hEOVfHhIxTKTuWKsy/Hbsd7XJ4teANSLRJR3MSKW9hxJtVPkyqhlAegLFrWgMLIk
6Jw7cZRa3qKSJEyRNBAt6edLp43mYBClp8zeQSXYC8w9KQKDnfqC9kENXqIMpRr/
SGL2Bh5Vc0NLm5MjSZxc5imvPotcuSThZGcQHCZbBr/c/rRwHRyMfQet4hcxDI/5
602tJDpbJHr2z2hCcd1oiLOJUwSjtnJwrN7z+nPNLKcwXKq9r5mWvCH7ktU4gJ7G
fAvtgNgXcIAPfDeOEG4fUsDwkAD02/1ApsMtqKosfYFGFVNn2lUjMqnlP64srreF
RkO0DoEI7zGkH+ArFFz/xZ+RKFLCG0yI/stlsMPkccd3YfAAn6WlF50bYUTBkMOh
TzY4MDpeO5ODjfT9Ca+vWctSEwjl/U9+mLFAAmgcLJ576OtuRuTW69v75XOD7ypj
ZGLUoVtj66jXJK8OllJq1H7Juw2HLQ/WiAXIZbuZthW5r1OYvLaJXl8ejA+wpFGu
y4s3Gpd69ZUPt3srULHLwk/l7BayoA7VTjkdIFTscHmU8TRhVhUUPD38OpcigXD6
6UrpV/HRmjbB2Oz7Zj045ybsidrSrb3N5gYJcllzVCFwVpJ4phZP8AivLjUicn0q
VT7Vp/EqxXUXlcQHKPWXmHKc1a/eDQWos9JbK8AWupmlFxLhCbQLPBxO0JAH6Uq2
RYYIfYynDtoadEi741Pcer4Reh53yjfbDGO8fbLUO+ccVajEXQtV0w0f6qLRcT7n
OFLzrOcusAGaAhezFm9POq4XtxmOinSWKPUxoEhNz/AD2b6FxhaaxHKQucUBKQee
8WLUi/fMh+B2PXk9LYk7midrFe8j4rGELXjPZ/Jb6CGnh9mI1AFpeD2r5NvNPd7e
h3FxMg3FAbjNv8uY4Z3QCqgFtt3+jQeRTWD+4UNWZCN1WevetmtI3e8zCFKDH/vN
1V/7jw/d8aVAIeMozFZ6FwBnR/kLtVOfxHaJuWJFVg3BZzwutrOEUDJcLSu8PGdv
BlFquTiFODcVAl/YXAs8dk8kG6+eaGyTY28ylHqI9cVGWmItEDyrWjoxMXm/zCp8
u8+C7myKkCPKk85UxFN5RUPaUBid+P7fxKkd6zqLaUe8quS7llOyKZyqYaKdkrxN
y0pzUiYaE+3tIYXdI3pNBHiqJxJC1ib8z6I03CG6fkr4tdp/MceCUFbDj8dGHxjy
Yp58WDM7OnFrGc4ecjiWYrO14qhoodXC19hR2Nvt4PS/kjy7A1X0rACYQiYrP2ZU
XvaWpPF48M7zfAT9YJHPA129GeiwJcEQvV0HGZLLGFshbBhSJIgtiexhPf/yrOwu
DpZAN9cnAF9q7PWukvzc/6/U4oU5XZ71SbRgl1/w6IJuFh8mO9y9o1gjVCjNPm90
ei2FWvAt4NoKDPsh9dYW/YMXfeGGXmQb9HJkDFkLZXcYd18aqkcF62f2FNTpJ7z3
Q8DgmYXMQbM/oUBlv6ytiTwmiEZioUo40sZzjEDBJ4XjsRS96QgV3LuWr6zXgQKp
9iK4NvNJwBHXzQ6kbsUQhDpSuvCYdZEvknKJhepJLXHELxmOBqEXOgfgz4KDvXyd
v0Wa1DwxYDCcGndbogGViRDkkpjs2f2i6M4mTpVhshkOBMFBUQYb1hc0QO3eAj7X
0qe5YziueAZyLPgBpdSiSiSSJhufcFuRmOO0L/Qi9gXTK2LtacqRblFIcijFgYzI
dpxdG7tYzFD7KrNNwKHbWpTOyTI1SIfR8OgW5qYfFSN66t88f4U99JGus1NG/AFo
sTILQ9wqaD74XerKYLq9iL5fIcZGXo3xCpy96OZ/2psW/gizZKyDZV6AE2mkS1Xg
Recy8vC2HzkusXfoYGsrVAze9atK8SPj8bAxsinkh0GkCniIMzD2Mtf5fCJCy9wu
Whi4NejXpva9JEPtt7X7YF8YkKhIhrRsWpYn3cNnmZRUd6nsCnrePPxEVwWMG1Kt
CqwSlIX+EyzsYqM5/kogvjmNaO0pFAWLJv7Qs0kmg0vFKJljGKHj+JZ2kboD19A3
Ejg9kbABrvdbjZbgQzeRfrns0LrDY79FGDAjy2aMDrP3N4zB2fmK6nm2Mi9gn/kX
tRGCejT5uS9OZjgEUy0MZ7bBodAj7CKlU32x4A8tv6KOsGLcALrsrOBsSpmd4UQ4
YVz7WZW+p1l3WBfN+P45OhrdUfxHz6Q3IiC/sNc4oujFJ/JgSYysfo2qTQQIbUNA
zrTQ2ncXAIPCt4g7IlQoPsGVpb3+pWhNN6wzfj9I4iA6fcC82u4UOFYEnUTw41Je
PghmHPfeQG077hHVBwVODF0i/v6yeMVgu1GEFS6enVrTlgV9o3o899QNn2GCrUQd
fxOrtztm8MVT36eZfljHjlYttvVE9SLubPeGRZQixvUYHrrJytzh/rvJq8SvJB8E
xJjx2K169D89ReddRL0m8jir9d1B5+BwPxudLf7tcpRbH+Dk5RipIB4HEJBFvfpF
yPI0T3PNg1L6UU05X6vRYmYtlflaVIFS9JXmGYa5H1xBP6YAyljG6rKHCF8marz6
+Z1JSpRnr6USuctxdu2V21Ng8iD3MiDz5oPBq2X5CG9e+HEnYWqw7xiNo+WcqFCD
o4gNka7arVLA3jkakqDRmcRuhCjT6EbXYI+eqX24w0Iqr16lI67+dwue8ZZbHBwe
dcIV9Ism8UqfTkFmHkg+wBuEFvvOKOzaSoL6Xut7lSkHL5fu2i6aKifDXoG4171Y
vBJebhxy1fzSsKRyjoDkFyYYOhWD7gCx33mtmFP7viQrVf+AnWlKeLMt655aeb8b
pmD5jKIybVqakC7GtaAUNDnVAbaZAr2P2wOFHMA9HEhsheqEY9uTfH8nUF1l9MMK
wMVZcCL12nU4jzcpNxjnuHAiBFN77UQyNV42/yERM8a1QWJx9+YOU/5mX3wPu7jK
+igY99wmJUNuRamm4WU6BTkIPTNlzXKFB/Pgv2PBwbRWniCie1zdiidYIrPw/i1v
6MQXShGSYnc9FGkYiCXLJcgYvFLUVwz8Wi0N5safViOu//18ATouAHapRdXZri5g
LGWd2Pn1os9vkg9jYBSXpZN3UT5MyiKy7Gz34lM8jg4anZDE9mgu09VNOqv3K/Br
12NITSYXficn7hrnIQ/bDJ6oQMLmXNlyOYe4TJ6k08Fgt8EPFYC016ygLUU0pPxX
8EF7zda3XUXk9NwjygAJEr83HYbrIPKk7e8lf70CMBMwK5sesNloLyYd0BCIH5W7
rpakYBmziUUpiQC4vZZP/l41RExcxG9AL0QJsPBpPO59sYNOqR6JvONdCtfCI1ol
8x4b2XO3lLI38Sm+/DDDksKhMsi7xW5Kqm2JoY7xE1LfRftxBQbQ1uHSr9bZQQdy
QApTqoEx74yPl5LMr/Ho606HlMC1sCyfqKhKgJBQGzOKcmdMWfXsnOpiav0wk1QS
y4rCvq5ubid/hi7Bpq8zvShPt03tEKzPZGRofGVZ4VYar5IREV7cJ96yQ1uUdDBb
FjGydeysM+3VNQ1TpTt+36v7D6YFkGD8T/77e1zJ4yQbIo1sJhdkE/ZjzDXYcX3g
sGHvsW5m/YjrhLw0bdLqpa+goE0Y9lhHrTvY0IRs8sR4B4p3iVv5nQvfDYeNQ5GX
5OUu7TXtPJUcZ3tPDceKhV1SgP0hlD3Qj30UjOptsiDicKBMw1LYVpdYaE9HDT8G
JM9Rq/3zorNg2dYai3XNmOdeEcztCK1VPS0RCKUX8z3wN3VpgLsTYwot/ycbScBQ
mYoxILHg2b0JQNK2u8KO/zxjl8JX5UuE+V/zWDKkyCwy0kGHHRallFpqI13g0k6q
yB4z5QzCxQuXKz3pbOvDzGyLByE2fiuGUoa3HZAE4p5nGWbpi61uKumkYR5jGjkD
MxmguArZmg68G+U1eVqeYnGqnsMJTsec+V5iYyoZs0AHDS1j8gqXYrdA2we6tjC9
PtKRFUo/kDUlavZ223iNg0lGN+iCx8IeBAKxt+oF7zYqrJlMfRKHEPx3KHjaj5lR
7gb/qfjx8eY9MBFNYnH9FydbdaOKE+4D5uaJJ86exnH7gga4CbUsa9MGG9xNbOq9
UmIdgsI0bWeOgpltG/egVxtglzD+qJip4Xwg3GsgHXyifQ/+mq6BhDJkiEmZ6aEG
191MxN0dq9oomaguK76K6swKj3tXhtU0hO66xTSDsqijoAFd5OMzvn5D48RDWv8P
ju/vMwj+pcvUIy4J0f81f5K6rSjaYkOJi1hGunWv0d0NZit2eqH7NY+gctWmf+wW
9dmpb4ZY8n2YwY/5cldX2A==
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Lkf9Ox3P0R8BVIGAb+qEKEyIzMyZvegDuqewYfYWfZ9GWo1/OUHIV9DFpdAJAG5r
qI5tD5sbb1qwsjSC2lrt68WLX2qNziU6zEI5lJNKlkc1tTjiEQIBJH2zxt7s+2bK
F8OMfc9SxyOPQcglnW/9mvJXQhyJRb0r48oo73ggfq0GQjyA9C9DnRGDFsrw7cU9
bv0dUt8RT2VTfmxW2t18gqrCdNVPgD26fNVv0jQnSIhST5HPPKkyzfe5HQdZs1UO
OdrBkFYYT05QVkL9kbddDQ0W/bdzNSH7BOqWlbAjkcTcJfNiHoslkdD7D1tIuoaD
0h0lt5n09Rgrfxzwi3uTJA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5104 )
`pragma protect data_block
K1LYlSW37xpIeEp1srIfGhL/S63JgNKZngJWp6YLdqhWWt6kjf2sgB2UGeTjvPx6
LHY7m4EsVneWi0KoB0NR/xW+Bteg9U/Oec1DMLc9t9uH4ILRlyDTivcmgXN3DYeU
TTMbfdDsdGuElQ4VVsC/bfUf5cbHRhPhRgPBIfPoheVvTTTbNPXIvM1yEeQt9y+I
Eh2eR2wA3t/PFukvsiGyIXH3MaSwFoDrCAbw2wDWvrFIyzFW5kaoX6tl4Di3aAuL
OrhwvigLniz0Tr29aldzaPdUhVqt7I5p0LOBngjL767ETmDbJwBYW/bRj/U2RGoK
EJ19/sP9zxDnTNPyRK5qo50Msba8fMZUo/4SUKPjVJEIRx5IPmJj1EhGFUuAswUM
qpCGd3otRmLk12/t0W3hJa59bpZPUKQxQnlRgu55dxg0MZ3dfgNMN0DUMwPZI512
mADg1bnUsHyADQv/4mOdeMclbRf6ThB58eUwt+XVIZiQJFAtEz2EzAru4iFziLqI
VTDiCXXizHDUbEmYmJu06BxDI/I7h7juR91KQkWvRWge3dMdAbF34LMrNKkDSQt6
RtjVWAmOV7Zy2q16lfigctfiUcDb4dIWUfC/DgG786+bE0JbiSQ6jYkwH9BLUGVr
Bqm+acMcINLNi2qwHpVlH8MuP3Zv87gORsBP63ctgW4uz84d5LX53Kt8dWSr2vcV
g7luQoTFms1P2BROQ5VhU2Woq6aIOly0Wr5vdI24tUpyZX82cXOkOJ9BIGSlhHB5
PkGJkxls6xseBPxT5Ftm74QMvdsfxDn4W7jlpsW2g4XQZaGjam00eLaAhVaGmMno
B88mDkPdrrHzA4E/A/lpePQ40bEivWhrjJ6L9Xp8SIg/ouVYQPqzinZxmLk51IxS
yiG1z6newELyi7RUKxPre2RgoruuZA1k+B2JXzF6KAPFvzjIE2FPEK0e9UkJSzsv
Ne88II8vLZHXzpp7V2D4L6A/yBsQK9qjYmWi5VRkHcNx+k4ZCRG+grRQYIHtjN8+
ccz8hWAntCq1sFX9OuOQovGhZ+ovUIpJgTsGbO55F0kKZGG8dbf5Zmcn3y13pdU6
t2eZB5rCOGwkvSmzeaUHwizWS6wDbC5loW4SS1/rJL3u4qxl9nzyhez3fMPuyZfp
6sbZ5FwcdYaAYDkOuyFCwMikoRTdIDEofdGylmS2JFBrcWyOZWopINiDIeW+Mb5w
LHxnbm+UO+dPdx/dsVsj3+MjqEhuvWwLQfPWZsz1dyRn2VkQSuAYUHgAU6TeTt4Q
7bMLSkw+6a4zQrbA84x3i2sfi5K0f2/RnP7HAbwZMocvuEHsohhU/pp76XJ2JIXG
hZhyBb6/0R/GgcnDiOTmdKYT/iGu11zn7sm1GCt/lm0M909rOPPvLSISth5vXVEj
7DMPG20TrFSQuabGE5cS/g3oUkFHpbOHD/ah+XGEyu8flsbwUKupjacnd3nufZte
u/+zuEQvjR7wsTw1rC/Nsi36aTwinV5HBSA9SSeg96Dto5ZMeIvn9QQYWwe9sboJ
HJb/Jga/cjFBJiFFTiavCgLm7p2lR8VOyPRvV41e4jQHIISfXWZan04p3ucfEK6J
oI9TVICIi93Q/WQLhZIa2WgdnYFj1v15m9E4TLv2shu0gRWKod+nrR1dyr6Bh5U5
YHi6NfuMNINZ4pAb9i0pnzq0tz4kW2mC/x6n25XMEkIYLyn4sQDWCGFWwxbLic2h
vM6/RRHMAVfEiigEmyDNfPq8IsjezUN3XHc9wfhwgs2A5iyHczcmFzdGEGIQJCFI
cNjnNwX8Sc4oOdjuCSPAvvUEPKlep26LHAxjVgVoimffjFwS72SpHSuWxesxxPz7
YFwzlGgO0qwMMqJVSvEUnfl/tUddM7flSyZ0AH5AvWklAWIr+dTNtITkoDzG5fjk
i6MwB+1hoqiqvZ/xWpIuJlFi/GRd3R58chWpsOU5a6gyrUOrXGepU3NWEgaUHYLu
JT2ahdsrFhJ8VCSszp8cGcYMVHuOB83iTwdkqs5JLI9eupdDqrlhsvjT9M1CfSSy
N4ptg8QlmwdzL2M7tHG6PpNEVOjpXYQqHVvQF2IiPVX3AyJxbbJqKQ+h9WmnIcvb
Thy9dtQ7cLcV6MzfRkEAyQwrYpeO8vmcRwDNkv6OwUv6bBu7W+ueMLZK5z3Rx2Nw
MMbnxayQkiBUTF1ctqU8irDt9+m01q24MIwTsiWlyAnfPDGYWj+Ebcc691SuLe5E
Opo5XFB9dTizPZldkdXed8yTTzcaIqs4Ns52//EEtl3gu/3R1QIaMYQiDWJS5UpL
NtmJaWoHrSnFSczxNM073ahUgHOAZI92/j/iFYnron7fRNsRiyybB4VRVM39G1gE
1K8UqDOEOOnRsfsqJijxWr9VTZgEB6w4lKt/1XAQRNufKaI84hlvBN8OHpE3ouMl
n8Sar2xse7B6+CQ8pQGl6X8WBURtKB0iVFugg9hMmApR1n0jXnNpZ1xNS213gdfa
8mo1jaD17iT1nHXCi6EVtSIdF7JKCLBQsRCwdFRv6lZvi0HBQxTni5Poo5DqsJrC
xXi6LsKY1mvJCUIcmc0Jy9tMUIJLfQl4ZFZXuXR+z70Y+pw3Hi1MXtxEcNYLpIKv
EvrMHi4QppvoJ4y5gL5R50Hmd9eCbIVBX0nZ3r+mhoX/Sgceh3gOOzMjdWQazlnN
SBQYnAJq5FksDd+0dOOsyhg52HGfwLn7j1ytDGTA2+XPUn3CIP5fvjrQOSxOveXX
i8c2bJYhTe22LZh08CUtpEMhp3KbWE9tqKgDjzn+vbxmQT/67QL3gcluUrQp+Q9K
ulezz8YrpxiGXJiS2U6z2ydQDPi/e0v3AozgSwthrQgnl+07bY41/4Z2up08z2CR
ymomR7HPr60qJVHKSmg5py34xswaG3dIAceBZkvT7ikfFcn7+zpD3zc67bGQBbPM
zT8GtvkmhgOvrZFw3ctUNZakGk71Wz9NyOWsA2NfIfspTCRqmlVunhQuVApqhPzM
+cFTJ5f0wRGwZw7C/ILXFzE3gh0Ar7MXiVY7WuTM1DgYl5qT8qDo+g7ycggoM0fA
l3CYoRpNCZt2X+KE7FTRq8ShsNLhhEb2JbUNZSKJReASSmArowNSJRUZxCqPb22X
X5QOGi+ygNANEZA82UdWvzrXFqluDUMFxsn5o8aMDFlEaOTJJ9mlPGM5qKYROAK4
fS9rvKnOeMYFS+aeAE3KACROPcViFLIbANx3NvNweux0vmpbfL70M1QuSoFXCCcN
xUQ46ZcOEBlu/bc0Mofc9qFomOhGf5vhF7Kvxacbi4M8tX5qQAavFCj76wNL/g2I
pO0L5NBDeFhZtFSoLGv/3W0Kl41SX+ajorRiA6duabjB1lh670LO+oWGL5o8wYxr
v252yXY+gJs56+qbUuGXOcxJ78UBKMzq6YOMqvrjCfh19ZymYU61LSd3OYxpdiHw
1pivbqndy4S5m5I5emf44s8N488/UZ9aakhniQ26PtQsv3GPy1BkaF8wAoeKkpnL
rZKIvTjUS8X6QUEuP/ghtc0vilZv2UalflSjvut4hL17Z2bikPE3nTXSsEpbAALe
+vclEiN/VxPS4kC9LMc7KEerTb1zzlcw+PB1PagypPMOuMOtrUJ0N+qtZJlxx6nU
vaEWIKztpW8w/FbKbRKbiUEhk90oOx1qyYmV6j7IsBv/LkbVeHfkmmJo2rfWguUa
nhsi+gPrblgbOExXiWXE+L7b+W4j4aC8ZhwPyEWn1zGB/im0+RWNLR2bVAu1Ihkv
j9FnmfqNyrHrukSucbeBlWh0OhLdZUQrs/QPvthlMbvNdIhe9NrumMde5QV6is/E
0D1pctSUSG/vtjdzcndHzQqaxB2+M4TTJBn6MKPD2NpbvZ1EW9zFIp00BoYnOYbU
ogpiB4wKTcKwoQpO/st40Rbu1sHa7/J6ZTq1PBM+8FBnT0L+mXvj5vVdhx9f39U/
P7raTy2ZG7KIGoPiqTj4Blw0lEdf+Ttwfpjyld3zgLeuA76XH2Z5ILY9cwF9eZtR
RbedZUPl9MNMkjAkgy1XCQOvcAhoHVVGMqUDjf1+nL1r0kHrKSAj8R451w/tjGcN
wVGZUlfjPL8tBjH9KLT15+eSzGCuaqO6oaKxi0dgB/Gj4ccwweDcR8GyjIyOWv3w
4oA3ZiUWZSuU5a16OB9jK58DDv3LfBQFKrWB6PTknG6D7yW7WwKSq5XnuPkweg/A
v/JDdsFb97lb2bryMwKZnkkhxbasv6lcdY/OVx5wBw5wiBoLCvdyYzemiBdMrDsm
vGaohklD3HibwsgvC8YLAEpKgK+UBrvsNMLgv5biUTMhz+QJwEUyb5Gfbg3XvQkk
3Ah3MKzpCfx1sboIG/155agx9rYRYBhxrQ13dMh0bQGwzKK2b0ejWjUYKjqXnL8O
vBlNOTm3PJ3wtRA99AGukb89ppY+j9Ave1mprY6IJt39M3W05lhu3OkZUBPm45HQ
Y18+CEUU6+0xP7VksfQ2PFZZ4Ofm5GOGL7QWPJgGzvcoxxKI7TE7WP22Ekwh1wg3
WraMZKzLF71pJx7xofgfwnWxdwSF1nA6lzyURiLxniJJSh1+BQtO3G1qQWm7HBbZ
JSowskJu+zz6G+LA+AYPkcF6GHWAxHD7L6Z9xksKj0x7Sw9hR4a6Sq9kZAgXJv6f
QsdjUmsfzqPuKadDHSof3s9MME79HJWm2z8vT8eGTaTTv1FcMZ/xMtFRprVCqsGs
uH9FyTvCnT2V6B6VIw/aedIkz447OHmatHDdw6PMMCvSg2uppXfKfPJmcYRD/l3X
ViZpWeZazMN4X90HZjPQ5HKH2DrQgzMnd6wo107+LM0JSac8x3SCC9lR/dPmNSMy
aTtGHwVSUYSUOY20fDNUYDyHEdnvR7MYpwQa7mZA6h3QXqDNjfSVA96IF5X7Aykn
DZwcgtyaiJBhwHMY+MtMoU5nYQQP2/ItRB0l15SwL/MvG3mh9Sj9boeOunCQzfWg
2pJzDkgcncLiK3Ux+AWHNU61EaG2cSk6Uz8hFh22chkWopdp8LRU4iCYSrfovoEC
7DNdTpPDsD236fgJY10sLU0j64+4rEjqplsJj/L/4m1nLtHRYp21guOUNvNt32rO
C0awN9yr27GAcm517GHtAhiF4DuDph+167CAUAdQYc9l05ob4QctgAHkLTwpdxxF
eQgdyliOoUO4RnLWF6A45cadY7cZfpTAWVLwN93Fr9k64vYJOc4/7LF854JKgXSO
n73C8FLg9Ita7vusJn1tHFejfaKLdALuKQf9UHHwV5dStbMskAMdi0KgYGinwGKI
+FPdaOOBiWTgBVDooDDWdJWpn+mXiR7V2o1Vj4fmFrrPu97srOouvj1C3a9jGsmG
fpLY1pGMLvXJU95rHll8T4fjZc1oz3W4ZMfx7ToOU5faBex2BkQVSnMb4kDw2dpk
83nfqewsinhuh+FoL9tfoiPtOfRXwBnjcbKCYG2dRJAG6uXQyY7wXlaYlXO8m7OJ
ePXTSSREfiOZWH+vA+2wA8Me1IiCNJfdOPwd2wpgzoVarJFIuKtJp0xTJSgRgtEb
Q/760Q9qSNgA4axv4MvcZ2OrPjNP7Os60GxE3NjmTsCDTAJE3akTujmYvoICLFKf
KUywwLYCONbuEdGf0VG7t8wp6fLkR7Z14JNNlK7n8bAZj7+HoXff3qZpsndgZ61/
srd9YqDSx/psSU3yHHV4dBSiWLR2qyo3nJ4+zx+HKLRi4/gjLGOBv5C1nKk0vqEm
OrvRu0Km+SZ0iJJH05rtYafuYWhOjVHfhcKiq+ydv2dl6I+j3oU5BujE/YpeYlH1
9338k/mc6LtxK1p4H8zxDbkwVBVMjwqMj4z6VvqMVyJme9YWRTemCBHXOby+2ONB
0gM/XwP+xvXubOWFK79Qbqcn3e7ifDj323SKpwc/rdbcCZsKSBOXOeS5KjiXg1TZ
PANltVjuy/nhVstN7bjvjEyZVPG6fAWyo85CJa6r78azsWT/y69Fg+vmOpybjVRp
nz8P4kAB3H2x54exBdJPVTUycZ5dLC5oH3pte4qaY70a6B2KUwY96qvGTi536YNm
LQUe1UYDut1Y4fcHZgWoGophuugsUx4AJy7t7CFrH1oAUGLnKoz0TDuuq2PJHQaI
yJRjA0sqccKJvRjseoGcvADuLHtDhexIUlI2plZDL5LIe3Fn3Mc9U7SbGMrpw/Oz
XbYFL2jEfQHxTaZB7DZaxeq5rR4sd7TlNIY6ZbRbMVPuXl4XiE550zUsofng2ezN
6Jocgg0di8T7dw1dSPOTbm8CmltFIapszYqbx/795r3Hqy0YHQsU010RbOdE7znP
XPim1YWLkMrmz2PKQvOXLSGVPwjt1gIdpnAOjZdvt4fX2PxRNlKwAXDCJbeWfxgq
WHyDcTV0iC7pfhtoJhp3HrMbTWZoBLQahM48RrAWhQx4JZQLzO61T2EqiIovw+4f
+XIni4FlELEsPD9LmdgO+9cPpOa/1vV+VKCabKiX3K6BSzTVdCevC431lCSpgWxK
wSY2Z6HvXb9OOaiyADHdSW7hRhbYjvpuS/iFMTOb6e1SpGUdaXrJOnlmeETXBDLN
Vxu/6kEaWKIxzjelVLEc7NdxKp62EPORXj+Eth3V/0ybi32r/SBADr3G5VS2rB1P
4GWb5yAprjRhufr9TAMcGCGcaIYfKT/W5GLJLMEBSDM5aK8Ue3k5EYLU7jyxmgwh
KGcPicxRGLEzIANNNPghKeL/RAKpXkbwSE1EQbZCg9wHw/ilnogoIpFGitnrDGqK
d5DQaBO+EGY9iGl2djDe5Q==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
PCJeoXmWiem4/HyiQSkOG6w1k64VEJ8cysI4jQCiltU1ZmYyZbJRI/0hS2qwPK8v
HNbzZHVXeW65eiJkhtS60NhztajPa6P9LhxuDU0fWay6rrx1nntQRUl5U80kpsJy
Rgao2qygKeYS/vUTX7W6MkiX7Ksm89dGhARWt2QJ1d38B4xEnfuJSZ31KozjreyV
ykjRliW7QMFkOIO5/nwbsNkVv5trnU39Rc8aRqKMvmdJ1o7TGvPFMgVbaeVnlPxP
qQaBoSWkSF1J51hTzez8ImkimiUUAzxTsD/QoyvB9UJKh37R2pXoNCXVhgzZbPna
hhywXuh37TFlq3Pn/p2WSA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2624 )
`pragma protect data_block
sMo6Kid0OxyGrflsmGhWYnOahT83K8BFvNX23utNKB15fhF1SgfF02Tfv2usFDUA
CfxDeZyGDvu3wiV2vMxvbcw/56a3Tn7XvprZL24cY41pEZZMBG+OSbMdvpNL+ioh
HdVLpR/73FBtkGa8qJ5+BthpOILW45DEsPOHpM/6ic9he8YpAjd0tJ1glGttx7oX
Yh6WmTFPfh99kz5tdNxVp2/Iv6ewGv5Qa9FMeGjLY2mGA8M8UEgrRSFiGzNc6rA5
vBG8X+DWoOttfw4gh5o9TDLW7MOixudbHi61ALW04o23MTFdBx1SXqwI5AR0KrUR
RNBZgyhlhweSD3+IykCI5JjpIii0MRYdYJAci7VdwedCpfPbDGTaxYccjpgF7QBw
m34D6hLTgsyzkvmdZBd054H6SdWiUBIyCbgtIDHuDEYPS3obWqHSKV+oy0GyJYHN
dbV6RquXbwkqCw2HUScASS8pgXZ6A+698MPpWOGXdKScgHGfXn+rnUWnYBi5Z4h8
KxrrRQfmGxaO+GAPwcHaBAk02VHKrrtMAWjVncB+agm+vYWCRS+d1vdVLkde/M8q
8+YU8wmoRJholggHi/QA3YkDdojGAtkEAWhDT4YEfPs0olAlPyjMqkLTWMxGr95f
5PBSVxYiJHTvSoB8/NZzBKa+GfwuSzpbmrfMXowJcSyGLtAT/qR5U02bldSawcj1
aSrMsj7N9HWzMxM/VBuaImb5rdJQHjjfKizvaW0zdteNNILLgKmdtewLZg08Zk/t
o2GHYz0ofpVmxpRGjnevF4neWeqvsYKqp1hKEwDxrwuyVEMqzBrU5JI6E0VmtKPT
Jav9bxjGfmAEA27k7RcSO4htaFdIiS28hLQ6fdAYdWV32KePDxV2SpQRYyIt6kRZ
w0Cy1o95uBE5fAWTKcIcYdKxMpioRXMwfaAYmrnS81VdYUPALkTbE82qSMGS6MCu
arsC7cCzPgebXW+7txk9xYmIldQMpejsXx7WSGBrOKrkLd0nKDlxDumgB2YU2AnZ
hfntFYOvyZN5B/n/HmIttN5LKJyTHbCeT4I0MGOx4QGw5f3liXp4FoJ7sI2O4TFn
otD1aRf/fD8nxrDdpUItspkqfOkBTRGNhC89D7FERefhnFUSmAasr5Qel8+nmwk+
EHJk5XrYUTN7J1H/vO8WID6CSTVOvIHBYyJDRg/K/7cNiSW4EblxIdgiJFFQ1N2Z
D3PthcD9sZsZnqhmv3PhmXCTiJsHhh7U1zluEqEGf/xXoF8U+W5Qdk6N0Pig+u5V
2KYhXKqdSd3ivMj0JSuurG2JjO27nerZ6XYqsVGEKpXlti6MG3ReOrOrkdxIHnxN
ZQOYKdY96C91ku7oIuyf1tonTtSaKbnNnhn7etG/NZBblo7NJDXvrKaScGfl9KHR
smUyGXbpB7Xlx+GffO3qQ9pQiNY9nU2nMq6p7jl1p0pqwjevmyBcO1If9b53IVMe
zWO6sNF0p+QdJB4cWJUIE9SKOhHsnjFznYt8WSpUo6h1EyTQItAweJvt+FxbNNdO
26pWHpEXYkY7J6L4hSQsH8/bv/n9/ElqTsWmfW1UpvSMW1fUbUbiXyR0fZkldwa/
SygZqw3f0kKqjk+W88WvFSIw5SJN9/Hyv208xA9N4gYB6agYdIfaSyuWCqJkq3gl
gMPWn8Yw11SfeH821D+4Ro/Fs6oLqYcKDSDANXaUYflOE07hISyuK+4UZHbene8E
ojTCyLPrUZprVmy0TND0R5k6iY9zTuMMFPz/DPXthjgRdYXMTkPUMgyb0a14adxb
lWtQ0kdhI+VwjTFyW42Zkkj1eLrmHwbJIungECO8ihCMaVeq0pTjCQMADYNlnqZ6
bEq9LZC8HgXl7fvpeK2oN9sfcvHPA+5Av3duNsdfs4XmYnTvHa+okpmNlfTl04Hk
2fImdDB3bTxcFrEt53/C3JmTEyIZVpaIbcrOu1Tyxn2rA5K334UELiEIgkRYrEiN
l37peqWEPTXOWTVRm56+c9zMq6kbDm8wSujQM+N3ESqxvqzMfclsZnXCPtDAymqp
qA0TopvcFkhYXD50cZ8I9+cEzgZhXQ/fFHGwQ0uZLLKJWpz+Ny4RXaX7jFLWvobA
7fanUxa7U+rukMyRPw57uP7tB0sOk87OFRHsMTGEkDZ6YSC30h92tEksnmSv7PDp
aZkJcJW5a+AhZxpgR5/AeJkpJUbkO4yHWnJeIO7X74lXnBWjSgSPQJqQSoCUabEo
+7nPZcH13ne8ciuNJgsDSuWWTJcNIVJ773QSZTksTeVzPNpM/crzWUYvb27WGFr0
D5UC8DFo/QGyULROwC89rUc6ewlj2X61ajeJOXcBAxPGf8vpXs3GSjv/3kPh7b8v
XAnhN3l/t/yliqmRfuanDRKlLD8mAjiSHzt9SV/Xn0gGSDNqHvAohJpDQpinIZpW
6cAT8q6nWLgIPmvgS9tkzAfJ8vwAHJ391KFAhJyCw9fkt8UiWnQekvD0/LKRuFM2
MmFg1i7qUURAonaFHeES91u2WcV1Qm3Th+YG945BQTh5+8SzE4HYd5HMMUxlg+M5
tVvrL2LFsu3/8O4INIUuO9dcQMdF3rTnFwXJIUQd7aoSzSXcQpuif2lyUnssZz0n
Ey3q6Ey3946G3kB3Xlreo8TxbRj4eVCJwEaPra5SrGVbcIBxS1bTycjbW7P24bql
9o7hJBpxGai+fQ1hpTqXcecIr0LhJ/VU67ldPynBQjV465rNP/zOs9+T33ljpWQ/
uBUbOhcYm6LVxaxqSmaN0TaR7WZdReXEM1Fcv5Mty0pc2DYCQIbZggagrDDS7I+u
mLwKKUnk0uqFEP1pUdVJnwiOYT/dk4kSbWmRNLc8oEfXouw/oBrQ3N1gyLzWMU2z
w2XZa0sg3bjxmlqxU3vqpvSRbmVTN7RAHZl6P3/jDlKR8mWcFuJfkZqhvnc/a6jY
L572BhkDHLXeuKfxG1iN8fGavtUamHTaC0cPYdX3UyXQx93knNelxOE5XCPAULKU
NmsDyJlk8LqogeB1fZkkKEsatAKVIQkTSmnhN77C0lB6vGCd7+m29hhPpAGE9zHp
7odruoNUeChiBxe+Sd+YV9xtCiFlDPfhmFMRaWPyUdcPT9VcGHQhENKxwQ51JT94
yL3bCfpZT/NgRgoV9yVJ5/GMCGExj/2q+RNTJboBKCG48U3PelQOSYBWyq/5sn+j
4sgTKBQWZcwEmh8ZVA2tcar5+XDlgYnRnwnTk+aj/G5x38DGQlZBCsD30uhr/0j2
Vys/fqYBUEwHkZv++UFZyMBfu1aAKzqcvzutWbXlFD5T0ks8mZ4JVw8GulrZxNQv
OI4c8HgL0a5Ua7/wHCYCUBEhPjSxlay6JB+VVE5sEqr3qVeJMs7iRDZVDFSf9JK8
0W0Oonxf8puhK5rkKCW9tQcBSqYuVQVYG9BZEHs5HmdSJAHW5Dw/7r6RtFucl/jA
kLwwCOdcuumqdqWyocZkLs4xTS0HJS7YEga2UTNnNdE=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cgU9wnMXqrc0/dMnqO+xFxbg9WwHbb4v5CG47kaojin+j/D1ZLowE4zjjLr2SEge
x2+/nar1IIhUcj50KFVUTLOhicQKmYhcalvYRVEwlPAeuEQxhTPyjFizGVZC11Ys
kYLbBSnkLoeSSmpZxvNvaaFVlMOiQhYIjJpyj4yRDpf/baZ7PIjWE/LIk57CKEdm
eQXULmjnL2jmcIET7oCnwyyrP5nu1uYgfuTP5tJJLRhMqF0fVLFvPsnKrEzcLDOv
ScW5w6JI+F/6TRPwkCHZH/IR5Y/0gcANGCPpcMYW7qlW1QPeFltlv33UJyqVXG/U
SE5i/d9j8o3c+duwBRXzBg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 18528 )
`pragma protect data_block
Inm/afUDpCT+Hb18oLHhACG48lGdK5qogW9+DxB/Af15TjS+0UYWEcibXSXklQKd
fvMWq/bIWrmJv984Z9InP7nLvnfMCKEZQWOvP3xJBUzZC1MDEmIB7edSTdM+kxiZ
qlFlmZJuTkHMXWydLGO5XTS/L6CfUFiWsxAuKYCRjGs6IYk95pD06/TpRYIKYd4l
6p6zq18nwwCVQM4lWpKj4HQTPJ81kqADVEbG8GGxv14cGTJllxZk8dIRxcf82Asl
6K3b39jK2nrvdeg/yrR8DQvtZuTK64FJWKlPCjm5sF+QROmOSCmitBhJwM3Tpgcf
qhLNF4MY5MOuzURb8Qh5A75/2riyYNprWLMCL8IgjvAGzXLhEclR+c3jne80IQrW
c7GmU3fpoSPfs6tUosqLBL1MtToDd2wwgra3vgEro0DpQmow5a+hkzRFpY3eD98h
0coCNPWb7HbcYc/6dyhyADMI/jQIqWQHd/eZ6HX0s3zY9b6G/cSwr2WcRkMMX5bD
qaaDKHzC3nj0GK1vNPYSuIFWN17NJD+Gm0qDChqIcIeFlJ5hNI5hxr1j+v1TlXJy
lG2eThQlZ22XF+9Ad8uM5rCf2gp/XKMyeaNVhLQhVND0zCXyWXPhQhi9aeevZECt
NkMCM951gLxhgnfRKl132Q5mXq/LLgeQ/uqq5Iw1nOOvYZhPQqRaDZLZp+36pl3l
5VEUh9q6dqGbmJVQ3i++kZSXS8X3hZeV84vgkimfpyZi8Am85ZImTy/t5XJJVbSa
ejC3zPBEWwjFC3uYE8sneLxJrs2gWWdvtgOFhSf8cmjKVP0CxTi2Y3ldsgsH/ex9
oUH91n+dCGJ+1ke5e2WNHmF4EKZcHJ8db626TRNMyc7sD92EKpI0u891A9SnYx1b
UA26ZR3oV5jHUobJE5gLscG8lTxbTSbukzKHC5W8MVDfYVgKANcM5juLjKfNIHMj
eJ/vE6DnCyvvmSIi0kXZ/SARBCqUF6zhQ+ByzblM6E7dcDghsnshtSPz4Omg03jx
TxzfLd0MNviOCdrmxd3rVhp96d5Y5xRgezWlYZUFm/GEGCCNtIWZc0DBnw42m1o8
lsc1fecNvqA/8GIk3tKBEm8+WRmzK/01VzkfEEYQsx1XkRXGcn26AQ2zf7lqVT+9
bZ3SfWn+9xaC04LWcZHvRzEGWiL9vM88d89AmrPKUx3Ec464HwbwkbeC2CiKdcz8
5//xhfP8mNDdjsS1xeoHoQklP5zu6yJgpamaRh9A2Q90iYiVqEGiJZL2pNIFXMIv
XUBx53EBDEYQ0LOc/Th86AOiu49XEL8icV7zX/bvvDgCnMEJvRSQU6ePhsN9YG3C
BLVlMX2+07zMOCeDQRN/wJkQ9SEoMrus9ir8wrNoH8Ky4XPg80dBmvxqmF3jW9lg
TiVxSzw4hvnOK3dpQVueoWJmi2/LWKlb9eI1XKtn6vRwq8gKvdNwqnbyfNsVREUb
4EvLoFKK1QgVJVZJtAZ0TxGx8RmUyU4ftjmKjsMVyc06YLfilJhdaK3vilink8qN
U6gulp60GAeWxwTYYLghnh7LEmaaatFYNmYMC2P5ZlKSEpoxLemjPq0U1Fv0ieAz
JAU5ctg1I8QIOam2ksEubrltc+poCLDOkTtwpkep+/yJCZy1ZMymSHXG3wPnP3vQ
cfeHdgW9V3OqqfqGGHiLhvK6fbZlZMccMds5luNBoq2a1DSRDn5cxRQR62vMRQCo
MgQWmpoHk+g52PDxEwmGekCi1i2kT2HrvdDwbko2+rT9XYCpFLmR8qWMO5H74tTb
300+FQyhohuCko2aiLFzu/AOqLLpDF2ib9jifoQxjK0pL5vHmGjvUFIujCMx4eHj
GbuNcReWxrJK9xLWVYf6MEZanrNmSSbMQ8PhNTzRfwyvQQMSjWmSGB/AvqRaX+rt
tC5EgrJuN6Gs/cjOX4kC4u79RTAqwY7uGkOdnLRevceGFmOCNEYaAzMxh79aJzuZ
nHZCr+xMB4d7v8KFQa3NO2nwSg6CUOEUjX1/WFrV2iCIzzL0XnA6kEYHBEuVLcmK
un/g1X91a/b8+30GDxt++PgOx+6EKd2A58mV2mIlsPdZzpfX/QvSxGvAAUlikvCz
Rxx71lVH+HbvxUmxSGHQs3AWj4jFosRkjEbd08PzGrBTVsQIrv5NNGG3DYGLEEZW
h3lJjjcuDKEGbaVgKCARVHoJjlDc5MESGi4xbJpr7puWnBmL0C2zDkTDjGhlYAgb
/wkhtWDyl/o8Ty6nuE71BtR3yNiLFe2KKOkDoipp9r5mDRpZdlO/4uhOqlEqdDZR
GuJ/Jqw3FtnOlpK6m/k0Jhsg09HqDgopiF0VveMMj8cOGFYw3byz/wThSqf5dOEK
wgxhTWooLAPcejXCQQLnO7fijjZKSQp+rAYR2Uym2YgZNTZ4BAeheBoeHm6hT+HQ
SxuuGi0INfDmaw6T5hde6lkVU66RSArdPHE4WvBGvyQC6SjcmaaZFQmVoMaNn5I+
fLtv958D25OUw+FNy7wQ7k4lZb2GzIRVNOTk8+ucIaQq7zqYcJitjB/wmbYNYA0A
idGg3tAuqNzyH7WaYrwkW2bmHHBstkQThFcexTvCa/BXZSRan9BYXkWzab3czpLk
8crdwjPvRRTNsEHicfpANksWVDWMtMWefZomEkQExTKtujeKzz8YrK2aueE01jvf
QsYcscZPqGlhl6eYyNBe5xf99qmwpjln37VbpRruTPmj7J/9MiLhFGz8GAcgSB2T
DLis4hiQCoMSSvibF6aK7n/O0vo8MRzoWjziYj1niG7yJdl5r1V9USqJKdJiWNVM
Z1ZNKPGZoUrUy2K3R/wX6+HyKnR13VJ4O35OTbPQ7y51tVj1rybt+hYHRBRqUU+e
x1WQiX3zVt4Nw6UgKTNgFZrkPZmuq7IO92sSopaB7uQEv3IdeoxA8qX0B07ynAVw
dQPTl0Ql8atqrwEBnvjdH4PPNgme1P15cwP2VK/1NuDNrhufHeiB9hUKOC7ZFFb0
y3qnzKWrsCHiHjaITi6jRUgbzOoyn0EFS6tZ2lqBbE1CIgjHlr0pzRgYcYmwHTGR
kpCjQ7y8XPFXAYluXYyKR/l5ZVB6gLfV0s8QWny72eBfUXzV8MAJJ2DLYbU744X4
i2MNTqo3tdqYy/72Ejmr6boTkZBOGx/X7RFuBuuI2Nx7QEtAKs/+YybSrXk+vbtf
IST6gWJMCPM5b+0nTLg8WISVebFqeSr3Wf/Bp6OAVsWvfHCr8ChObhyGjVsOYtnv
kRimikmv/1G+cDY7+/Bg12oHKl9e++YvzH6LA7i4Hl69JHrDa5Cb78nnnoQbgp9s
yOcYOuoMNixL36GFl881VPgYYsFXcjm0qDMxSg7vLiuPzIzHsqwNdAwUvc9u+dRW
YcJedBJduvH0YwaYGIFh9CO6oXU0o9BobkpOO4WCkz51dKWtcIbRJsHp11r53QZj
O8S2Pr22S0m2CaMkiSwSEj/K1yES5J8Gn4YhtxvnV3Us6Y4OaNGzhLqYILY1AEAM
XWb5ifiHwRlSCx4XLLUTw4tZ9zu9OGFeeoAPfRfMj0ZxCxhw8gwnPkrGvZ4caX1v
seVjPpQWWsC6SeY1GOG1kqZkvuh21Cr8ZUMNyZTFdoCr+IYowCTwAE3hkrv8K3yx
Gj9vXgZ4D3qMiz1/EL5KpMQJkin4eIm9+gto6MX0QqmFZ1QFVlHL4o8Dn8+vO84b
LDjQTxmu1kL5GXLs3+JtNM6eYkQ+Ux1Y7V94vFviO2J5mGbenB5G6kW0rs4TTdvS
i4a2rtXEQ7K5OHXueLGXvpP357H8OhgBa24cUdEtTaytwRTWXk9zRsKgtDga6sHh
mHvDoixtw0PznUZBNi/i/TcXRC0+2yJianuLhVgKuihGFuTN4zd3PKejPKiKjXqP
jqNYr4F5jOKrT43vl3AoJFiZOd1DyDxiwi1QdpAclGq8IebWuihqy/QUK6lWxIY5
98e1hKCjf9rglzu2RgyOA75S/08iUv4uLzK0mH6jfSYskr83pYCoy4wq8b16NxPg
jxFVKqhMcLn6uFdK0NPi5c60yqCq3Aby1zlBLsP0KY4woweH4yfr1iDdCnL+cco1
WFLw0FE7uuwGSnmDLgzIM9lEnw/m+YgrYRTIW2VES6c2ne1HwagP4MHURZyO7npy
ztAWNSgjuyIexYqfZueSi6tsOw2UQ279n97O0Mm5ITh6um78bGTjP2ZELoDj0zUo
kVUdCwKs8MjGdfIebO68U2oQu4mqeEPVNGGMq6taJ/Bp4qKnBhLDMwW+w00SgAKe
8+BWVH3DgyxlmFgiOG/x9eILeAZ/usIZyM8hahJX7MZRNtd8M0atifaoClfaiLB/
AdEusFl0IISD/xXlk/MbY0I5kwJGB+J4bB42f274tEyPRlAiSmL3H33tn44ulRMc
XOhZ6M874RYxH6mHoTIr1sNrDIpNHSg4xh5YMXGLw+CEOcEBdKIr0vRe2a+6IJDV
BI/EZB3WMQQe3zve8jQZQ81wQ3wOhASfSgln4yXrDXURYZNh5FQsxNvAfnkCUZWu
m2xou77VuFLvd209QYn/L8EWB344aAg8w6xixcIMLzkQ65wTNGhSvuk5Wto8gvP6
ioiW5PJovw2CsFy0CoAP5aElz3bAA3gZxi6M0MiVIXtCuUhjGvpQaaxcTuAGwBeU
1asPZ5VkfAHvwEbJolSIt0x2zIMBTSZiOc+ktalktnGxi8sxg+sxFwHMrNe72Yle
HLpTpPWum86NnpibLl3U8FsJb9nXSeh16gWAS0axLk3mBLB8gvqs5drjiIqH9IEY
BLhw3XZ5PfMU2G4FgmFZXVg8cR8SwjNdxELRDhHY62MK47N91wf6/rJJnVfZSFNY
gsZvRDrPMsIpCTLRGWlFOsBVuZSE78wpO/fWdrwZNgxb8zH+5AW0MTUCoBifbpM6
QAoPMQYa9ExkR9JZhgec63lpVjRA1hmWGW9YLPPg3S9ZFjZtndsz+dC5F3BcA65I
V9t0YgEIp1YHvM6gfB6q6zHuOudfU3yjjOT7Mgyvj/ibV8AVZZxPv3ezb7exvo35
s00rsa3eFNOPBfzM5QzPhTevvj1stosi1TGpTuFoBsi/hlRmWjqW5UytXT2fd2UX
hlB3dcH8nHAygNXfWUDCGT1pJPuZbZcpQwURvvYjCXutofjkSbxkf80kZPQG049O
oVw3hSoFqcO8A0HVSE6IzpR5xXi4m346412A9D7mq9WvnGLgyTMufva6c41Rad+K
c5qWlTgU/hhaJXIvPuPrSJ7tuNPZt0Aj+T/UnuoNaRUzJzyxIpBloItV06iWpoyO
WVDJdhidPWxUPiPmRqq+H9ZyI/SeKQEqsMju2mw8WQoq+uotMQpYjF6tBZxtzdEl
ob8JzPenSr9qpMv2kL4tt9XWUebR32oJ7+bKltKgJIgGVB+Q8wHpD4E24n5HBjso
p3Pyh5DvgZUyLidyX6CES52cHkfGaX8rdj5gguhb35KNOXyEvwfyp3vf+OiHvY7F
BgYgV5CHQ2Zh5xaKzDvFvwGwaZQ1aJpcL0ceQmsGP2ZzhZu+YSUENtGsEw6kRn0H
7CCEIQezvrl5Xpw8kw/yRfEZ2dOfV11gNW3q6Qap+tEn8bsUsZfHQDUk9i3wTVyK
REh0PUymhE67vNWqABKUkc6GRARXrKFYw4mcGP/9mpqEhC4KjJ/zhGDZGqUonv0E
zX+ESCRx/y7LJQRlNfLM5TmMa2oIcmZKW66FWvNn/yXbvAE0mCskEbp1wfmcND4n
Zlp+6Z2ZbumetnIz3rCCCNAsEOH24iXWq1Huh29nZoln6T/UlskIPkWUbFJHyFr9
hjA2aOJz7fDheBzzQhzI2rxrBLqJ3afVchKfleugIVOHYumSG9JFgzTekMMz2DOV
G8wnszI/RLQkEX6agRmayF0nyWH6xTQgmKM3Su7pLBAYWlCnDZv3cT78QWXNEnSb
fgZYo8h9OJF6FAfrZ0TqS1mYLCFchmRd+Q2StBEkPOI77/xH/tFPSI0NOeeFN5oP
leJsQW0UAe5klOkp6KOAXxEFX+y1qy+WManMpVFAL6q4xtrW+OrbhKnZ9a6mYN6c
KUXLDSLr7+x/s7RmxBBKcoQKbN54SrfXKuMjomHmEnbj2luzNeW8efMQrMWZxJeu
n8vfnzddpWg4CTeldjZnqRrWcrSDKcJnAwzHS6ssdq3qJvXTM865OeA6EmUnSpGe
C/lNZXOj4digdaPt6hQKEURXxQ8srZCxxs8yUr6q4Ks2MWeKsvEm7oEdKTvJXW/q
DwfmkcvAI+Ty1jLv5ZoNCvzZxhz91MyptUQftRm5suAOiZEitLPgUCto/TRA7czn
3cPnQIoP50EB+t8PjHzvoupfb4mEV4myWitsKWXCDCBZZUp3mGYafCFsBDJjZNJL
UEYm/GYSPZSkssagJjr1d7zNrXQYv2nKf5Q4MBhbtePTdHxb5QwfFDu3Ow9yyspG
j7hfPbwyxqhXpSaTii5w2ISQV7dsLSah+RkKwAJEyl9qbxYRajDzSHdP7kuD4esh
WhDtW9BBaMacF42hgl441pO/4ACWG6j20vcks/+OIvbm5ZQbd2nz/H+korKj3LGC
V/TCHsp4oP4Uumml/lX579qAbv2ZPmoI8fplwnZQqjBbhboyYgYcJYUCaXC3oWpb
RM3Cf9SuI8US3juhjkr2qag3WaVmRNQr1xHG2IjQyahLolSQxFDU3RHeF7TLsyYp
FSX1Poisj1Y4NXQD7fvKFFXnrr64GV9YpWcwtVIfcDJjNr7kgCBQSrfmb3qdPNeE
yluNDlZgchNWTtJDYYHg0zMrySJ6LjIloOeH9A8yY6ckvNFJSZiuDv0JH/i2/vP8
zMdpLK8w/k6XI+C+chmkbxegoBvvG17MQXVCNFztqYOwGLJAY5ucV77+phV8OZ+/
fUMVkRsUWPJL9kVeKe2fWJIlxLoJpJ/kiumEcHGg8DGrd59eeOHiAsMTkmnuZWCM
MFCkTWuPYAK1vJ1VRmTfyEGj70T5sY2lO98WQRholqFoINaVOp05r4W/eWaN4oz8
hQ3M2bVuG93UTYnNh6S6P5VpNz1v3VX16aLsJFAoRYNyn5YFNIGI1TwZLGjC5qAZ
aOMNmUiwW1skrH06gPvGRFKziiQn93wUR5a0Sody4KsFilS0Oleqhmu+LnmKo7C5
jvE0cDskYFMgiM2bk+poEuloDP7zsUuage3mWC/mDP8IraG7ZhugTuokqNCTPauk
GJh1Jvz16cZmitMzMlutk7qM21KGD6vyxpFQCcxpyDAp6hkUHrhfvoa1468UXhep
9B2WkYQkucpebnvvElLLd/5Dq9KX3zVR4ycPwFYGzEShyiIxifIRlrmLRj5wI+Hq
XIWx1hMTR6c3GKdvwwBIM43mJ/j5ApHfKkyYU9EudbOgdNFWom6MCDRX5hz4Vnom
VdsjXQwiVctVzVu63D8ZrA3xncmp26chihsdcpJDYKvIj1YtW/hspV4x9dnHzbj5
DiERvIwsqjOsd4IPHx4Ha7lWxG4VaGARUS+qO3sbmHBKQQeEfJAw8e+jEHafpwDj
eTDlqOagAQRw4HtsdEYe4SBW3gIrAqvvnSim6mqA1s9on4LH6X87slNz5nknrGoa
Oskn48TyeaMpNg6+hZmOr1nmDes5yugV9vwiDJSpVh7H4+hBdTek36nC16TAghDe
X/Jl4cSwYX/dUaVSAUY+CWAJNehEQqMmXrZhl9zPg90ugmtjRxzVuX3FpPSRrRz6
Ai8if3iH7tDci2ETzvv/HXqYYBIEfH20NTuGKl0PJ0cSMLb4Dpsqtz1UBSFLm7UN
oTCM3cF9wRmhTU80iLKLWfV2taT2Xn97LKH8oTsfg6AhRKAKx1L244WCSKMpnCEv
Ebhk44Cgg3rcTF8WhXCliWWnccOle4zmGKpGH0aspain2U8Foh5siKXud6prhe4L
Rj4UfPupTt8RjcoxxDWMASC0lHY5cV8NAn5an2zkb9BSzCHJmxNpkVmYsoMraNXU
GvOUkUHmZgIIA2eC3eAjK3oj9XhYseBvnipYUMgk1TCIu9FwkfQVSB0iCvgQIAiD
TX9A77AmIXXpB6JQf81ArM5zn7K0yCFbUQQDaOgoIdAyF1r/+aWBXEaf4BcGgXPW
NnFCikNOepbEIIVZRct3+X7slKlz9YVjrj6gUeIYUUi4JzvCKJJWLc++VpWYckLb
U3Bs9tV4T20vrBFRlpwFTxv1Oju+lAwUc+fEetUkDGqdmtcC8LYly3qLCc3GhCfs
sZbftE88OMKBhTzKdtc0ZzZASCf1nrlxj1vbpchs1TmhEPKPY7+ijLnKT36nBkK2
fsORX+5WHUiZOP7uHWg2WrN+wDtH9sAhfTx6joBKZ7vV1NfQyJCNuV6EeTgNb3O8
8ObuE2hGtqhqV2UXEte7VJqi5E9HIIQUaYoMd3jbEtl7I5KA/Ty1eWqt9gshuB8C
PFRw/FDurOZlOMbAs/V24lqSDor2fQeIIdsifPcBq5PH/y5W9XYSwXcrNwpnvkmF
6YDWA0cCNhlRfcoqhaipcMmLM38A1/AJg2xO3rV8xS/5Fgdt5/nD4JwWatUhvuw5
dvj7WYhCb1BbO7Q+0daoNIpC9Yab62Yij2pBSgeOVMbKY2s0PrvgbpYSXdTmcqfj
2zTB+676YM0Mno+dibAFtpdSXRXbvBb82nPVy3y2Gdw/mplJ6s1VNadnYy66Xufw
KV4xyyWcDAZnHIA0UFTqRTocrP9AzEQUP/SrzaWWCbVfv+ERXYpdM3czdW3Ndc9L
qvBGBl38MjG4MLJN243ksronTDPrPdEhR/wHJ3FzLH3FXwYfObhPE8gr6mtmgjOW
H4RXT8bZ4vEYb4NeU2R4WG5u15f5XXCzZ0CLso30AKXdFXBBTUU11pty4mWJd4+4
qlP0wYyHi1kWzyVHNQBVYaK25v8sMyBjLsfjJiDJ1V8fJkIFrxkYWqEn/iTOhT0H
QUWoSXp7wAJ7xRnMU6ud2W1l5lUzfKFSfmgv/A+zvPmz60XXAlpYR6PZ6RYsHHwq
V3+VgAb1p0okQhCcXvj6IwXKI1whsvtIbaltgrM2ubtDUiKURI7wknoJnqevzOtS
5uMAUzkmb9OZ9d9MZi+K3vlXZKpGFGNIvTLWN0qqfQCdmM12Jype8/GjLjSF1eGT
Mfi+UHH+GTrmHeoZdAp57K2DH/bSyMBfXXjX5xd6fcJUPHx69sriyUwvkmogHTsk
yrGCQdJzU0TPjct58+R9Osfarc0i/NDlhfcwKzvvOIqfJwEiLLFopj4HH7odY1W9
aUqJ9o/ZqApbUh/L3+h066kzK12vNfzyQVt4BKZSE/5CvadEmx+73KnrEdXvdLKe
O7ppkNHaXyu473k1jKjy0r4FA1rwV+XtHKE0oX6HxeXIIGZFr7wFORWzAsTSo7lN
jhWAWFpsiYmbc8X+mqs7glueq4AB/wQr8P8HbvUn6aDAIN8UBeZfIdCfJNzJhjV3
akYLhh12HhJTjzX8okT0M6MjVQyy8IP0SuSAx6pLRjw0VPlNQBirrqkiUueTcte5
/KFVF9rBT5o0UWnsZSNVpVIWRz8gMrvLiGwS332OoTYcRc5DyuRbP0iSN8c06uJl
ZCZNdj2GctnOQV5kbn6dK3eW5lcwfXVtnmq1iK5PoiAtqfwsGYZmc2+nrZPEGvLs
iZxwXRIQZfgfPaNKs2AonxgyIwZLY6Q6zPmwayXOR3GJKa5C3jSj0lhwf6ZuwBqK
3pKP2go9kyanLMyc2D6zxV/jAvMHpbs26EWlxsfwvETG/W7pfTFsdYIxy5Kaj9V4
u7GnDJWUBBwu4kSRqMh/d+c+yTchiBXLC6LjaCuYX77nD2zQTuhEazkjLbCfFyNh
3ECeBFt3tnSS1repeTEvuMvN+Y+5LtnQ9kuCmQad4ySf45Y4By9igWkAd7wwSGkT
WgYe45+HVaoAwSIR0zyz5CRU5FThNC1bzf19TQSR/4jCYZSDpVpIVRc9al0C3OQ1
1Zie1DW2zo+D8RwHU+f1Rq6Lu/yqHMgYA2HfO0QNxPrnuv402ZFxp+KMthBKFTRT
jXlBnSYztHqhD/pDBDxAsB2vGxjEcTI4v1b4cJ2YMEPqGCjS2GOI5ltG1bf58c9i
D07/9gGb5DIeWL8twl6xNCvLeP/kBhn7KmWaxC0MuUuU1129QQhxes78vyLQQsr+
C77MIoZcj0jB5xkHdtysyV6/zYpIRDvUkcrSTF7O8oOSdg8E19TqFZNBqMCRdFFg
T2jpkC9Bo5XKZtmy77xweyOodFQj3uLZhITlY6k7guXXOr/laMTyfBhME7zjFiD/
WeFUtTJw/k9A9hXtxDzfCpUahdlwScDWuMsYZoF8Uy6uqTVM+IawVYYHfXrsncIo
TvRBtl5Ki6aT06gfc7ybdGbEw7HDKDyzZvMwNOw+GX9hemWB/7zy4h6eQlP0wgjX
weqMM/tbNuwCqiGmyBdlWvbM3SvBVT0EblJihlx3n3m3xrv7q09ImI/TWJa45+3V
w1x9/6l9UZkCypdW25fEeE9VrjzLQ8F0F8gVMKwDopOj0DuFHhtd1+w19G1vF7RO
TWoPXvMXJ5jF769vP7yvsTzRsI7PvXOeYtrBzGHN5N1Qagztzq1XLkyZ66h2R+Wr
wlXT9UdjzjcAN1Kvzy9ufq/Lk3wULrLdns7zsCsM+4Xu2VoZKs2rQ441yqkpU5a0
VbnwES/shPvZIq5BvUW+n4dqqy2+AxItN9JMXZP/H1Q6Xd3etC4XOqb5LvyyMQvr
35aEvawrMoFcN+EkbyMHd6CQBEqe6pwX0k1VDiasc+JDKN+tY1eDWcchrOFgvh24
yrhBpqNbi8Flbz5m6PDTKkM2jnXE5Phd6GqQA2eeBuMSXOv0ZQ8xPPB/Gyz6aqHp
FXXwCpafD2moHUF9A0whD+nB+qVSqaJN+TI8vKsG1NpLhScjklgg7jncKyh6AUys
HFbioWX91oXuQWITvCHAPnRy0URc4D6F4s27dWXo6MqziqfucoI025M6B82qGAHN
Rkr/0bOuFF2Frh90cOUky/kpCFBnSZsIQn/YHtT1zcQunzYWY/hY85RaGCyhyi18
SzGTvk+M2AUpKpW/QnT/RonQtDtD+qnA5YkltVVcU42vDghPlqqpEWj/J5FDAs38
DWLtyzX+76jFxsTRnKwykVwc2hglpuoPj85OR9KFCnhLERarUCzK0AO6HFxiZn6a
iqyziB8rjy0BvIbM0+juTeicSw3XWPCtv7im3jVQn4ICwyHf1fMo9dutuXSchBbC
EtDxjq1n78W24/RqY0omKCauxsK0hk9ELU6AHhVZBBV2LX/78lxG0ONQtXDOJR4g
edGbXcrXDwHOyLAC6jLRlB8ZWYO+3ZkndxP5KNWfU2Bf7jYAgv37FK/3SETy9M57
5hGZG7cWjWyS++SrPM0IEf6KXO+Jp7ZbOAo74rKdJ+B3Eo9SLgnA99lBQdAxwvoD
MjuPscqVYP+mwnR9Z3Pq1Yyc2ua1n7TaawL9hERlcGc3830szRGPo0NgHF6S6zk5
ttYJ9nuAEk7QVimJ+FCgSEjYJeFJirNUkW37J01vE9T16dmlAKM/grFj3Pw4j7TA
i2ufkjlEUqHTFDgAvaJACF/763PnznYM7vDqoj5jZ6N9gakVtQVRy7eg8I1kuO9v
o5WUVrnTbujhtVXdru7xLgx3PudFh40ePYARs7cfx83R3WFmhAfhBpqvXPYO9JfF
ibU/3twpVPU9DBevy+Ql1yN3j1pCSXyJ8xsqq8YTbCJFSzDV0rKtCHBL6vZCNQnq
OsD0abuvRvkIL7zobInOQjfM317mvmRVOODSXRC8pPnUPYWU5rCh8moYzPSwaEDC
YoUW7gARq38ilkAw3GC1b/Bu5ohaOrZsSZntvH9xwh+YVId5Jejq6QZIE6laOSoF
Q1msbOJ0QSb4bhZeVhno9bjGPZm4K1RR7qRkgmzfwNXYM3UNKb4UlCF7K/p4TU34
6V8dQhS8YXUjnzDOVdkpYl6eI9pTmNacggF++u8K+oLAilvvhr8OMEOl7Xqg2RlL
ToV4daLal0QKwRyZ+lVyE56Hlau6eQswbvgABzmDRdO+j/4PJV1HIFXsJ8r8UTmb
Kkaw9yxMmuin05/kL31zinJ7PWpI3ILs1GKogg9aahqcqlx1DVwvQJLVuLAsESuO
nUpsws5lUNvdWiT76HNba45pzrpvQveXYy7R5DbYnjkJB6S3y0EvW6jy/I7PxAGg
a5EmphJqUtD0LelX2oehDI/1ESEi+1s7x5Fq7JpdkgJsLfK63HkpLpQH+2EU/MtA
J11qHulWzGdrPnaMNNvGcmAZgVginmW8r5cns9m3Aly67rz5cULeYkrMZfTTsYkG
sWQiHlAEL5fXUtABAKxnXjX5Bz3dX0I06zpdl8O7ISrpd5y0gnrVxUFHM+EcCOdd
PTufekacFFquJUfV6vTerOcGEHva2118iGzER79SvD+TiXg7YOm6NSM/s+baDgvb
qnQZBfFdRzYwE/uppxZk/Ma7i4Q5I0ybKgG8lf3LzUtCVlIlOBujprzhUqvgQm6Q
T1gxQ395ZwOfAx1OqNKPFW0WxXxQoZmFOmrKbpJPxbndtZKG4wq0qR0rAHHSb9Fg
DdRIRO6jqM6Rdzm8E8ccyYF0/WwpyoFzoeOFu+J+wjFxAheLuSkCNJNVSAku3SbE
sxSiRp+2RQt0oxk2G9hs3IklaUL11NDhdR58yNuTc9+JHtAadmMLyfyfjUifhBRx
djeSm+CpF3+hjtQXVtGloMECPlMViIWL+p6g3RM9kWYEypPirZFfJS+xVTRw/aqe
1ofB4Ubxlab7p0Og6HLPpL7S0CAGjFodXHqFWdUECKKg/g82rlS+MmJAU85UZENd
tNP43Ml95+ms3RaBDQvmT3oq4bRV7PyX8422mMiJAH9XcOJ4i8ob2jaNWS6qhhIO
gebkG9JTYFTGWHnaNa2DOQjfssTKosG3/iqtas84XZJYaJEG/5HSauLWRhEtfn06
C37z/U7XNcObQV1HzAcrUraUUQQ/tSL9Oi+VNNc52f+xwS/LttO0aXFSMLcUZj9E
B8H0sU6ePPmrWgyaVPUsg5+vkXsT7HAWVL3re0YpDhvtKYdar+ifASEneKOwwDFl
tfL7ha82JsP+rN9CDDuQiLnHzaQSbM8EJLBJum8vsAMhMeXP/N20FCldseNoYLvN
vF8EjeJNFjJZSX5ErkjrnTnmbvxgRa2MJU3zDgrqWRCkTaFa1umJ+x+gudbfWB1a
SD3b5Mu1Bd+vc/hVsRKcPGd/KYOBqTVwE9Kyw05yrCKMhToB6eeLo6NTD1kAKxla
kwlMkyNn8OgTyOyfcR1AULNlfX57VXapCcY8ymc8lWLXFsXaTh+pR5yyRrhbBKhY
dFyw4gy7jI5aRlUJaNliAL3wpvmCnBY9ss7jvPlNxHn44OZt5sm36/1pVyN9MB2q
RXBpJZYTtZTVHm8eM1EuD5rUMerTauLwPA3oYoc8Mq4XSR5kOSsZFFf+rFDxNXB6
rEE8w2H5lspU+3Kkjd4T1dUpbz0wbPGOylAYtK+7yCMI9REWcYV9G9d8MiISbwnm
E5v0+pkMDBaS21OX8+Iqv3MzAxtFdqJjGZ6Z5vVouZ7c+Hy+0NrGJE1Sl2LUSfQh
dz7eU96qgKEa7ket7bkkgDUjWhAANjMWKUk/xEEDqayex+3dA1FBxEbGvqicuJ1Q
tbdfxcT4N5eysECfwHvDPCHe5bXrYUe63PTLNIboJPC9BU+bXe2eeXZT7gBbAYtd
1HFNyHeIrHqOmIN7PfOSuMDDHI/eYFHGpfRLwp4V7sEiPGECf2xvHjD6DPHjwMUG
gS+4HiyWMwxFSxKAzcmgLujfcycXaewQY8ukmVq+qgJxnMsQtHZSMeYcNQTsPLe/
GfNZQuPuHx+5ZpTnp6Td3OTj2qtmwuNz2hk5MH3ZgRPwhMerdWis74G9Fv53oM6F
uSxFoJ11jiilySBvmiQxFPfzlZ0A35q/ldZ3+ooolJI8PXCZppUeDTVtf2pG7L3G
0ChlGz751TaIm+CHNGQRjCq8/Gr2Y7JvQ86phecKA8XWuf6/YFyBVb4QanNAl61G
LVPnSbfaR0QU6oyVrCj4JPW2pAVMtfON/7CMHisjtXc52wuHYOVeRwlJWSkxFsXW
VFFj2Vj4AlqbcTCLjRHg7p66dlrVQS9zNNPMAtqK2M1G/C/QefGPwAw/SgOfdYRQ
dkS5ugVNeBu/YMshra+P7MwsTA95eA/4emnETeMOzimIGFtYHBGbDx5iMQxl02LJ
A0cbMMvT5K+uSvpMMEQwZb2cJUtKbgSTg3uplAPOP+Cm43jU7tCmpj00ezrvCb+G
YKMLBYUw4T+L77kG+Atg57ZYXw/thUviNGhX8gEsbmvPuMIJ8OTn9uweGvZy5jSh
6cO3f7b4Aw8bx6X2ZrZjJa5i8c95Jhe4N1F9ILwFTWJhYDvUS1ob6Sa4qdzPve/+
G/svyKmIY16VbkBQkAQhHu6S0grlD9NGe6nmHx57HXxTCfj+niEAwASA6f8lFzPc
pTVd3wFkhaKh6Y1FgGd47UA8F/e0iikRhRlQpz8NRiGxzielRJQlvO0IJe/2/uiu
ELcMwstdXsC4vQSQKXZTXA9J8Luoz24baifB0k9Y5uF9nYAHuaQWcprIn9LDCCjR
jl9WZIPOcL3K44k+aZe9sGEk4nc0xsWjMkpuNpKBElv9bIQKc+EjCYe3TBSPTU+O
YJ5ZIbp9gNgPLI6Jt2OOeyEDsNDTHSNYuZ0E99xDKZ17LipiRAHFtu9a7/0/rUXe
xu//Lctp01ZQpHmOz0sP5Q2fa7FewU66ewfCEbJRYKTSLhG/uxvEEzTrjrf0t4l5
1nb8JfYlh2gy7caITTGkuGm9356ojw/4ZX9ZTlZGV9cBh8Ok6/lWZrUCAoCSTR2i
JeG82Hcu0fYtiDWNJIU/EvOYHRPZNLq3A5UNEharuLMxfa1qQdmm/2CQqwzTEQKU
Pd9/tOf25WwOJUFzigQoNNSr+EiXgE4U6HS2HcqaIA+YLHwjFr8n0wVX3LLNUwHZ
DYfH+BXo1HfEnCV5H9jc7R0RqO0DV+O0MCuGGnyXc+8tCOgDVPSWP0F1u98ym5rJ
JPR6T9qe816pwDoy86dlw1vR6p/grNmvDSZK7Z18TqrbbMv1xp8grXLe4ENfkOQ8
w0O77b9kcQjfaqvKAzGSKYubR4mpfjuCN5dTo+spohikiuErdT8yAuKTEeYaPZVX
i1oW19ZIof/Ktj5orTgOlhfW1ckB8/qcre7rDvgD68yuGJmKcaHN+5HSXGm2JYES
v+0VGQBMFVUe01RDA5q+pRyKZvIBcZ8i7qUYrPVkb4k22UqA/BKaZg+DEoLmxfli
I+BLjkT/SgbQUE3nuqHu6O1bcLAR00Ma2i2Y5ixYuWgfU1KN4nPdZ3QF4H7gfQy+
Wm95J3VcBBxjPg+QmCnMeWjbiq1sqwyY/RjHBxHlNxfLHe4jJDYbhEYV7MtgxOAp
i3qgXWJqrNAKXFze0ZQjGUc/nBfML4isPkC7ISL7J71YiZS6PCGlFtZNr23zs0hN
d0cY4QB8hXdI/InRwemMjYDG4rn82VoYcYUyLoaRtmYElVOLjSeLiHZbdYx7D5mJ
46nRisu0SGXJfzwsSgx4G+8qL0fVSF8IuX5RbgXJIOQZRrhOjqzw2Mm5AH59fvEE
1+YEUAi6125smca1kjXXZ/9kTBJB4fRqR5GtTfeBAz+dKg4wc+wcmzgh7SOo7tKM
e1wc50cipxHUaPPiMW8tK8XXSund5bnp9gx+fCzR+3fOtvO+gJkZ2F96PfF71cL9
1og404ntaWRnhJtYvpza8VdzdyXyaP3puWsaAcyTDxauGL9bcWtdhcL2Dv7s78re
gS8zH/qSgYDVfFxFhC9MLt+7eidKexQmQgsnRlBbRIlj+/98dWgn6IJluwaLg1C9
DWJx28tpNBDJ5qC3BGqE1+l+YAwYtxLn+pZQxLAvUgsI1FteROlUS0di3oT5YEms
eZoZyfcshFh/09/E1PtSFG+bW+7QY2/MJCYxyamj01ZUFiZd9pkmsXnti530pYDH
iyn+57Y+1VwaxbFHy55cRqOxPzUIzDrawlC/3XeQ1n24SDQSVHAokZTrIomCwk9i
SqjemOyN+BH+ZIt0pp3dAom2pjnXVChADmhulXPCy6/hCB/lLd+NmDdMzEo3Fg76
nRzvg6vJV7yyLgwj3fDrVCSmWYlriv4y3bAp3i4bkwf0KEBV60M/cfKfBGjZkYpw
62PGT+sPzKzx4LHSFHbPHJnt8nwq2VMrdp4zoTNBI3nEYcALu9wPGtZ9+LYC5KfB
orXAt1NOWbyfU7+dj3MRkYT5ve/3M7oEsVp+giRpO2DbuB3A4Bd+EPwHIyv2Ck3B
eAwlzz7MPCXSEbI445DVrZ3+YUpdIrKMKPv/R7+bBoDr14xcjqWSW/I9NdskIAuq
NhBVZnW1biann3uCy4dktXdi7xaPloKpjuHvrTRlhXnYljiqzks5O1EuMNbxjkEF
hqdkPMpWC3Z+BuV663Mw+PDE47FssQsyTw+TB1o68D8LXTQmn4p06JzwYAx+WR5X
LluDzhfVrW5YCChl6E5Gx7G5mInPe/PboxopraW+v+Qz5B9S8D1qF5t7e4C7R50D
wDr9vUD5UtlkyD1BRsjmhSp1CbP+earC7Tsg2cinHDw7gEhaNN9p+voZRnIuVEIX
lopbn1W2hm1rvAteIJQ2PY2L5mwBr1hXNsGPm6qVGXQy5/BKcpsQCNpNxpGacOjD
x+CJYUHSrJe3wojUMuHICgD4ZHabuKykqz39s2EztYrSKYpb0S9MXFQFYQ03y6GQ
S9MKgMTDXaXHqbwDSEys50o7Jjs/T0WLbW3JWSUNPjBDqgslwGankVxMZrFEBmS1
DyjgolEJIHzjxNKRt3wFresZs2/X5DJN6oEfj+rjONo/pRh/BORLr7igvGzHJV7u
qgjNPJ8RJSw9i9zTk7I00lSRE7hcqRKvaYJsmgDDKBDCe1T/stp6WSGu+WyZRMzB
dKX2JNCyysUGuGE8OyMq8UDuCbl/adTQ57ZBDcJfDn34FOqcyEYEdFHLB2VDZcUA
NWHu5Q/XrD8k8OlX1rCbxo5joncV71HlQwGpFRnzYf1lLohHtO1hKo/DEJ8H2GqF
idk+aOtXPmOU1OZ9ZwvbNMbDljQDqD3gbWQvjDM+ZPGRdsLv2wVYqYc4q0LUiESy
lwp9POYiDmEpWRR3b3GBFQL5I67NfiBXOYIIzTidTwsufXOit5qvNEREeRG7Zc6b
qaOgm0oU/rGzQ0JrZvSDUaa1cTLG/xRd/0+OnpCJoWyUWIv/eMtn5+zQBHmbR4f0
Of97GmxZef4DwVltdIjnpW3YpLuySZ+JLpazR3evzj3EklZlnN5wT/zpi2os+Fvn
bupt6BollJPJtozAUDWKeXnkIfH2J9WeewdeeJfLJYHGI07JrRaOaLLA55iTBUR0
H3wsIxzbjD/HQT6RMtAaC2h/MmZauhlrZZGtCkyCITouBMxZI6aWl+EI4iEj+STR
+TstEDYhech9aZ9+OYOpyi19vfncaw8/5CFHFOiS2l/SXI0Z+dVBHqHCcq6KjTRd
N/k+xpSaWBLZfecPrA3qdb1QGnJtOTchfiT+uYdMFI+Nty5QdUeiqoeXjfmD7oGE
nKdDgIw5KdUEhrfz9bL2kTXNtb+DVJNz0n9/wV38PhEXFuZGtucftkP+FoSAnpDS
5V4KtcJCBJwF3d6Tmlf8o+RT6N4D+MD59QfFzNa1xViao4u9JmfptmFnWTH7Tcgp
2mEDoouXhMdbWeO8gU7CLtixcd4awyD4eBV7uzZyX7FyVxRY9DFw4Frm9Hg+B+8V
lFVxtSVwclv4V7RJGL/nnoxdbjULblK31TR6FCCiKVbsGRQLsbcxp6kydNGazCGD
lUBW0rJKHl4LR0iXw9KS0Px9GwuJfWG0dMvhUKDDK8YQ54iIG7vSpENDIaM2/Il5
lNh8AkMhHJttBUZp5DY+xjVb6GzAYmm14s7BG2cSppKo3dbz5PITpS25BbxQFjVI
notkJ3qnuYCeWP5pp48/iixi/0oyFXoIHB5WFaMPSNsTSnv4q1WiwbbiXe/twyPB
mohusPhXxVoGX2T9xFPZq2UShPmyxw+7N8b0xIogWX6dmKirSaT0+GnR/kCJfJio
gVysOK+yENOdwG7TDKn7aRpBep2mfo6N4rQgVTkRWeWnOq55VDLGRqa7TgSOzIsk
4y1IxA3GL5yir+6H5aCjCB0iWJjDLq4WvFXWUgan4H/qkCWZqgjW4hc4+fg5yy6X
S9dzEG4RQ+FBEA5SG1olXH4wvwhJr80r9Tt1crsteibjj2XkF03m5Mb0u7wQpsBI
5Ew/eSpez/B6kVL+MA/Gc0gyqzKSp8+KIid36yOnxjpC9/Ve5XLASgsS80EzskD9
zNx/KMn5Rc2Vh2ToXqeP7cwH8zs0rfT17D+M+1W0OkrOK6SfJQAhenoHsch+yaSk
I2qb0f2U0srt9ApmHejxLg4AY0PqP2OxrPCwe+lxTjqLxSyibtRKNkYtAOCFSZGq
qlKt3W5OUZZYs24s1+eukWrthH8/WU+FsPatV8/GLhOG9Ki3zM9sI32P4Wvz/wLv
9kjZCuG9r98iSwjbG+KNCEJVC0wkZmQIVeFm9lEgiJ5IGiepok4RKENYsj9y2ta9
7SZrepTdX1328v1en8k/AJe5moS8XEOAklsN2g9dS8V3bStSHiom40KOjMRXCYrk
T4u6zPjG1uTQt9HFL51+GCogwxaD79XTULZ9Wdex5EQ/dFa9DNj0DJ8b/XrUZG9k
8YbwtQp8CDID0SXb5MqkIQbWf3URFXc2Fj4jkWNwMufTcAzq2GkmDwDzAXhM9aCw
5800NciN3gwwiEzu8w+oMbbJ58oRgJvJmaLsvZAP+sy7EHLE556WJMBeYPU8y45M
GlVTJjcLkJvWMFH4o83jO9Rci0v3dnYsCJdXpZ8uSmB1S/3ceU8OeMuMZeFxPoEN
HvM4rOImxAlChIZzW+pIvRIASnctC/p6v10s6Yr2R6BXIwQRrNMPqObeGnQRzf25
IQpFudUSAxzm+VRw7Yb5bk8/UEV5ZAVutSF84JxOnRMpVRtW/3tJY4aVJmq5kjce
gayPSi0ZiEtLB9FyA+FOCkp68Sg731gZsH014WaEphE8CnzofoX5XYtITs8+WmlQ
rPTupWTYozlcQJ9+9JZIS+CCHwle379rw/mNuhfzPHEWfdIiytx3PTLLrUB1swfB
ORP72jXhnDHMwHi7e4F+OZvDH4dwllsQY/YbFytUHMcxMa57Imy9Z3gIKesIkK6W
A60w4YKLc/YJCwtsbxmJsrKMpp2s1F61T8jsiblF4QMPMzcFXKnvdRninh6TFwOv
FkXB9n1beh0N8skMREGcRbvJkZOv5eHxVJQgMter+u7rzScfKaQdxd2EFEuE90xF
E27D9VSVeDDidt12U+uwKboXlpJZf/vPwJAkKlIjonBEM92IEiosc3CbFRJZeWmc
AXdShOqcCy5FY1Vb9WHvi4cBJIyfj52mC+SC9jnm8or0o4e12NDoWNHmgH9onGHL
KitVYoutfPtfROoVl/7N68jnW971wDQJpEb5ifpw/kxO8OmoUojqA4xaxkw+rvKJ
Bu7043znQzJntbw8/ZzV+ODOi/CflZMbM9+yxHYJD5umAKaAlPyeJXXVJRNPMUxq
Tzv2m41eVZKDgVQh9Dsz4tu+4mFS7uNaBSKKqcLibtwAzH5dogUfa7vG4irTyfjy
glIqumah1d3fV28ooVUcLQ3eE8yli9/5XTU+gsrdaT7UuNJaGzrwCdYsXDRVJCXR
unNeGY5i+I/Nx9ZeGFQrzmdNJBGwJgFLhQE9Nv6XgOj1Z3CQ2aAU7IuZlVhj3zjy
FeKGlCWYkK7yrHMM7uIqAAfEfRVjI9tzhKs/Myg9uR0h4Et4ah5lhtz2sLHrcIAr
hThrHhr1FJQa0CMXvJIGmVLhDx55AYdiA5c2fzHCfF+rw0iaR76pn18vyhT5q4tO
yB+NB6GqipxVusdjHQfQvnuVA+0B06acXdDzaS1tw2pxY5Mahqj6IOYgzPyywdll
feyStFj+7hSLVadsm0y/mN69xtuaCJ6gLSJ3d2cUevz3B0gbnhqP7xAtnTLHIrB0
J0nyce5P1SHhH0wxmb6bnL/88YSE5Kc1TXO1k1fpKWCx4vfkXKmqd1m3eQX01Y3O
pb9tw+Z00Mfk+STIJFdqk/gKOh3HRGbvSazI515CkKUhxxkj5vbIsebO8S6+iH1t
LyQG7LqkLUXXhs4e1gBvYjpPTuxT6fMBYuWNYsZPQWMW5aaf7+2prYgsOOWUeemI
mqYyL7AN5GxPsysCYxvnFn9aombmim1j/rADGdDxVXFmfiJpV2c2csyUjPiUAlT9
M6qxXqyCbaCn7YGvjmDR8vhG6Zp7kc0NofOcLQTS6e390mmNKk80o8OzxGZWlbRU
pUf4jAAwpfPjVElCp6gHU1j4zEp/Ek+9XPYNxQ6jMHhkSZjrMg8R/2xF1iJeCJim
LGh/8Q/qVYBEXOcpErgMLjrj2M3HCjhvXSyvbX5gJD0mBfIF26QasHo03BKfwNJN
KHVKaU158/dA7iCX39MeZsWhIG6J9pEhki+1nM2bmBB99FxsC+U+jAIfMfj7F02Z
lKlhDQgUXufMP6Xb2d+QW+spxGqN6XoMhCg7vI32MenluqdLCBzgx7AoTJtnIoDp
g4/F/M1RSnwbHeBJqe3k7Yy24XAm8+v7t1c5DQFkQ8z7UTe7o3nZDInYQC7C11NT
aNA9BON8tDIbs95r/3iofkkucXn3rFKnDgMYn0l0OgPLTGDXAk0tFVqf+Sv5s02N
U20VSyptIrGDb/W6Lhzs3HTaw1TqAtShWzjoBei5AFSDVbMbbSBt7o6IsSAsaufD
y6ORVrQzronXh1higjQnw8bM/vBjMwKjTRld87jcknUYTQMZJ52OU48aiZbBMBPR
dJtI6DZJdUgXhpf//EL341QNf/4l4tWZLQHEB6AHqdTHaWQswYpDuLwiE9n23gtb
u5Ts8txKNJ0Lkhd/P4MUFbQDUybx6VF6ZyP431xYwEj4ykskJyyFJpGL9dWSot04
U3DodzDO/ZNxUZGKjmxE1SDx5Uh0pYaDirI+SmP66RUE0Q4LPDsZ8kGpTWoerDHA
EvObELg/dKx3AOpSArufd1JxmXJbT2ADZjWTF+nscDZqzDgmfAzvdbF6au+qjOcg
nwaKA/MssbF3hSAB9CqZaACrgXbJfvuXZSFoV5fb13lP2KVLq743XphstCf6m7c6
2ygbSd7IYKtEMUuyjgaV2OF7BcohtDMtI/ZB29yrmJPXqTzQpKRd/oRKwipjItYH
FxpnVCTE+dBW64IMgNgFA3ZB4gkvOIHzOc7xgaw2BgpJv9YTgjdeRhBpFiaxHOYj
tKZZe6RyzVkREumAR7BUz8Stx55LW0AfOSoo4izM3mG0TmP8IdptzrM0QO2H5gLi
9AZgcvNgcAXmwhYfz++gS5PdzE3EqRGPfsidfCyezjt6N+RXvNPukpy5Gffogf6M
OvE26aFTNhfQH7HtX+tDlKVGGDEe8gj9yjbHqD4bOydwCsLYWRUApyDEcNlNXG9s
soMZMGlNyKboJQlMyJbhdweNBm+1oesjP28ApDJxkf1jCv+44CYNvvY2iSsixmjq
VMaHxKUK4PemaI2Gc+flOTndievnfmxGkJvJsgMry95ZQqg3VQciWMemZA3rtFMI
jjvnJb5GsMXxRQqfgLq4ApKX64tvWBQmwDGXmOgLFlHgkoies5/kIvSka3y8/9xb
5fbsMy9ZnayzdzPTyWaQvqkRhx1QPPlwDkDKrTzjX3m3PReqpzPAZI+2q4igaNTE
PzWDclpLg4yDgkIXR++h38+WpqUbJ70YJF85lbaOPlO4B5MsXljkoRIP0Ys4jwGd
oiDb4n5M7jqWlV3lZjXbPr8yfVql2lJyWQBgQF29hklRFe/duMYri3RFEBLaO5d6
BOksbjq0bbr8PkF1trrGgW5m2C07X0CdnYEj/HfzyCt16qr65xFpOHmpOMnRhubH
gp/mB5uPug9NukO4aZYxRiArLQCObIuImqFX+Im9e0qXAbFNscMvlFKnTCDK6qvS
BNa0K2ip2ADE+9lCZcgiLZQeKEQH7X/NOOdZ/OshN+PDZ+PgR7vx+6H9boloWN1P
T8Auxb1HoFEThtiY+ucHLg00QoR3ykFTKRuNcq0A0JG6i0DlzMzZ0m/05GH5m59x
PPt8CIMyqCea6hliPvrylNRLn6OH0ZzQCRiRyct4t9ngmtKGrURY+8KL+v/FiFPb
9HutikSjqLVkUh1nmkEaTIiXhoptIK+fuluZOkz78zutGCNtyLdUlnHrMlaWbur3
46OD6YrhYVsRKXu2J3meFbs6N0z4bGVG2CTjHjPb/REEfguOjLZvozNKGgtiTOjG
fvvNPfZq8dI5S0W/vaq5KR6O/Sy4dZra/tOHCTHX3e8ZjVlMAP6EkTBQYDQKA5/s
mQez8IMMEm+ELQ3dv+B/yJXpWzrn6Kd2kATmfvYbR58v9aw3eBZfzM69NeZy1DoM
wxCVcCEiZFGDD+HLA6dXcKjMi+zKH0IG/fqhgATf5AYJj22657rnxKCKS+2I3VuI
Hq8cLD71hRCTi4+R41OE2OcnxxrM6rgTPpiWQ6v40CzuAicIVUawfteNGivJ4AcA
hd5P7633jeBQU+UBsGwm+WDoZa8qA+oUwRtEjohCcz9o/Cb2nrEC5dblo0Rb5P7j
9HsqJd6WxIJdnffO+WVEXn4teHTp3npRYNk2yPciD4IVn47c3fsFUvHJlgbs756x
nlLghhEg29SsgcPockDP3z/POBgPpiHUQNFGjyURGQAVds6kn/bkHoIzZZj4UC2d
lX1scS7Q/SFTFYW8Cr9HnJUdkv64ma14C5ThyM1Ty2Gf2pHd4SVqWf+52jGXANFs
WXNrfslThD6eiYrbL8OQXjnCwtL6KVGn4N48m1nbJfo+Rk0Bxb2fZGMuf12M1K1j
4M8r7Kyf9JdBYPEXE13Iwp29Dc9pVW79zRx7aKP75YoXAlpDNTJex1N8DaN7pJM3
Rzak6QkeXhX7zg6sFizCGzSO8tp54tqmbadyT6YodyzBMyKK7Ue8SiLcbTRyE+og
dCAXMop8OwDGUA2tjpjdCjntI47Sh1tsO1yvN+0lPVnJDURa/XlHSMil32aMpo+/
sQMZG6esef4JYaSJTFOUZ98Ph3tsC/Hcyn2Mxqs4QvXMQyBoSqsdsH5EShLEx4aX
YkJ2gZJQXOgnHqBWkBbXNqzD5M/+i30JFwUuQ5GdrMtfim2j6Vr+wcvYt1Q119Ge
H8dFuNNkhppLujyz6x2YAubDSupJ/LBCVX2cqTEfHaFVOy23mB2K7tsALq8roc5x
NuiLrCc5g9v50ru/xII6DswC6Kjbu0/lrkP/9cENxodiRaZS/S3iCKOFa86r7K2w
GLKZYrJDX/HP+9G8AeX9yCI2X8TW1LSe0FXr0LYn2WqonR2Fw/0//RbiyBrW33BE
hRauDsgrgMLt5Azn+guNFN7jIh2oVv+cPWSjjyAb4usBhEoo4Hp9UD8HEar1w3Mm
xAOoySNUpR8G57AE+EWutr0CiqEAeRHQ82qKQ6frmJjU7TXordVN/Nj/DDRWSzme
/4T3mbTKCQY9EhMk2Mrm63SZrmjdewnW6A4QuqwXKG9HD/bCFaBBujpTiW73iSQX
aqboMqgI8+ueBCYzeJsxvG3BTW2LTV1Ldtw2XFTIs2KA8y/nP63owvfJVOX7xXW7
K2Us4jPY3N202czudbkviV+faa2H/E9zV1jj/uhhlQT5m3uYdlwo3WxKdlayTKDM
YMsmi+xL1N9Vj6ueu2+2pp2vNGS+h3snJ8JGCg7VignVkYQrmrmXArhmYmnDPGBn
J2LkRGYF04kawK6TnnlcpoIgzRmfdBByy1N9Yg6xGsg3IY39GO8HUfReqImHYtav
TTUo33JRkXzhTZ77V30vrzoTYfErddO+FIN5Snzg/a2znO4IXHWegXzFSHVlW/UJ
wO/lZSh/y14Flg+CEcyTK5SZsOone27/eLO1SArcDAPU0S0/HNhLLd/zyRkvqHjY
voef1pHOfyvVgnMhnrVWDDmmwF+c12lSNNQnLlKS59iAeKSkpjZrJuJryRos8C4+
zoOvSUZuNNYRPYM9F3CMt8kndTvVZO3DBbmN4AA6gHa+qJiHoTXVarWfMCOXMJ95
PPcy3IRRcR9TrdQeuIlrUAw1O4lQ7UR1tVVevD8bLc+KgvIM4PWJ2z/lv9dYBxlg
moH4thhTWdsjtvHSDpgwZ1cfCBMxoluluSDkYbvgAas8JubqY+Quo5ad5OI/XvdJ
qRwsN8k0P9FCxjacsO3nLiqgRj8hORrJPka9QVk6rhkYSrNBW00Hg7fzh5FKjtx1
f0unxOJuUsXBtRAEz6tnLcSV4F1b63zYAjuV5Os6YbcEUSckkWWw/Yu1dt4bb5RW
oiO+UQ56Q4DmNrNQ/E/UZ2kIhUQoMtnKDq9MjeGXbpIPmMl+g01LWvfsTs0v5sIP
JU2k7Oz0XZM0NRPT9223DccbMB8tIxxMUFYUgF5dw2mKGaGlQDP81aL3yn/oMEGK
ZcAZDiJzxiWaVYP3362qQ/hOlEslWjAZn5zI+TFbKAQXO5CS3GOm4LYWFfy0cTI/
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bWjVFJwNV+cVTl2GszCGPsKRyL1IZVClXPOGnC1DD0LABc1dUn+VvLJuSbcX6IZu
fqGGnORxE2nUIobuRNV5EU/Vd9aGBqAn8COHaz1W5PlO0+6iJo933A84DoiF7onR
IyEHFwbZjVhUsRwycFZp1+JLDLqMUeQqvMhcefe95eOpClMAMIaS9eGCLEygI+PT
M+I5wQlqwVVdpw27Ly5jh80qPY2UirG+NFGpdlFbO+0uipYCdR/7j+8Y9EH+LJKT
3M0GAu5rfh27nV8V9fg+XbFEBxdKgDdNgOJdBJWH8Go/KDPuQjnI15AfNTLw25EE
JcKs6YB4WUzQF4My0t3OYw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10448 )
`pragma protect data_block
sqKqc9sO8YGpqSiIIavSxkyu8Ay27CajFSkHaXqCOOl4iH0QtSMeSAd2OE1x0pdS
pxw1Pe87hVoZ1tTbXEADZC0uIAaXbB+NljNgfaIRl/XZilgSUG01C3mdkcOFw3Ev
Ybw4x3MvqHiRNRpm3f66+KhB8K+XkClXbMuyRbdqqUoxP1XeQX84bhryaHxTdEhV
4ixNaZDZi5iMujLTJGO31P03LXW3xK2KZhHjg/lyrVuo1SrEwI9kZtpti2TFov9S
uJVYffl7nkX9G8QEqTl+VtoU2LBpm6MxiF2N77YCME86qoJTcjGH16lVVk/PuGt3
la6ULUdIpUfiGaClAKEoLfl+sEtqBEPxEKMEkVpg7roQX1Pmb/+6Jv5oHwVop/Ky
W5YOk4pucK5zDF+S2SddfrINarR9x1HS4xoLSe/yr6gerUxnx8mDXxj7ViRwwy3z
/S7dpx/KLc0HXBFOD2D49S7EymdNWdnHktQREkheRXvPQRS+SQeRbq+HTz7NeLV0
IvoeZE6wzdP3dDxDj2PQB9+avDSKpwP7UEs/oCqdkB1D1E/8ueAyWIyjcVUSJED0
4uLpxPwZ7+nQTARUUdGw1J3t0sOgfWUqXi0wIMQcdqSJLo/2BKA+YJa1HGbmbCoF
Fn+VivSC3gP7dXanNpDubj0TawCuFARBpj8gTs2Frgq99bg1aXvjgJVxKj7JY5A6
ylUUOhVZJgw44AXgbKLZyqsMbC4dVBs7TrKuieCCRcHSLAimtFv/Vh9dx9tVIncN
t3mxKWadj+0O4FIpj4db08miaJmw3NrXSafq8zbTmIm9f/gU8yGjmdcgOPmODhmk
ZgJUGevAEFbvG4We0YE/t/LcQLwNjIXHD6jTjJ2uYEHoMw5cLGmcWzSzpWjclBD3
7TfIuLq+0EZo3z5CXEBkdqQxYIhCKDa50qBnXo0oOMy75GTM863Uw0Uqoh5+WCa7
ytVSQNivxmExlU5rMAbwTo3yQLTe4FCOehKyEGppcTur+5CthcLiQAXxp0B90Qcw
bBe02L+p+usR29rJnS38EXLiIIuSwHMJzYWvHaY3q0czxZCFQdSgl630t0igBOEl
hNUHJzbKGQebRZacGFHcD36Zvuq9n3oLnJkBFBbWAtav45j1ENhMgOf6EzHaRz30
YJRdYgcHpAF+j3GvVrGNhySFe9NkqliAweFXAfUPqFSfHiaFvT4ugQB1rftLqcSa
XNdOSo7epRsIYB42mg4uG9jtRr6PO5c67BE10HF12TYBFZuA0RPEnjA9diqHFXBG
vjNfkt7QDwaXFHidY+Qa7KaignICYthVHbDNDu8UGsU+BhrFwj68aSQVo7FeLE8q
GJMrwJS9BDdrXeAKr7vgay0PcFfE3qIhDrav22ylgpetqlxoEfevSv1x7oLE2RA2
36kJlpAYFIY27XdnGbdjx2xWQAgE67n6iKcvFk/PNtXkpMu2TvOnSvvb78WaKLsY
jxZj8qGh8Bz1g94MyDZrBnXZltgnTBhOCNDDHdVrqwMQxaNQJSoQIAqkO1mrEyse
nt6bUFGntWrWj0CQ65VY2D+JdGwNHgxuQnOp/k6zJjRuELwzSyc3GrmYHSaphV+u
S4OhvQDfLTtgUOBLJHoHn4z6o8TKrV3mhKXzBqmhRs4jDphVa1tWrq96ysr+DWvf
q0QLxoZsF9RNH8kMhQJGzF5JSrgDBduFJHNzZIif+fKmXZcS0N37SSy9oadFjWP4
QFLH7ew6yef9NeI+WfJ5ZZUvJJVvs/H9kWgwUPwhbprONn8Qsigr+CV/TBcAKJb6
wKMtQ0CctG8cG27aRPd8Dqyynn3NV3UL65w+TY7YZbhBGs1t3/l3N+RbE038NrK1
hr1z2BSpvrZNPhO7BxoDcB64WM9s2r3hGmGkj2LOU+lCh8NstIuBuIHHPI0tzMjy
0bTW1wmF8h6UZ1SYKYg5s+pdJ6rC5Spq1tElFyyv8cSNP3Rxu6fBGHAIxhYAVwI4
oYAk78pbBrYS4njhQdcsRjg1AJWaAKPnrq3t+cWj2kPZYM2SPMfSUFoHNfcLlpDS
la9dqjv2OWgtyDVdVshNVH9HKnhDz7v0uCI0kZP4ftC/Fxj8yln9sXsgUND6gCj7
W+BDXT8cOs/IxFeQu+POjv8v0lYuRy0su0V0vKwvKnhK0ROd1Rq3h2QSkJ5PTGNy
bHzjGzdrcPqD1ygFgjctGlPbdxxnlc1Krj/A4gnGWFkOWkozQ3WE70+C6wecj9vp
8pTLHEuHGIbZkXfv/+0JL5tMck25anvtLcUcLRi/yo8E7tcU9TChCGfSmUdOCdoz
AwFa2OUsGDzWStOdAKU7aFxuA6Dc/iEz0WEWsaJRqcBHR7wovkT7epzGmX4Vat+h
6CIYjWyEUWvR2Pczs2A3nPYeQRXBChFla3CnQXg52DNuEdsQSxAjcqRzNvVJIlh1
4/Jw5+8cb3Y3gJYLyM5UYiZjpoDwg9vYhaEdHNXQyxsVFsLpyVYU9Y49xtKtcHj2
qhKTgR1prxf3/9tPzCyfWHkq1zIYUaZU6ho8VuguJiVjM/EW38j4hPvXF4oeQltB
iznJneu3wVcYAnxUd+smKL7yX2FeG0ZyloPrsRQMAc5ci+rsVYQWT9jfCryfkBUT
StzOYy2SjKPrETCSh3aJrZlHNr3VRLle66PFE23QllczDEB4+2EK9m5LMTbTwrER
jdccfdpfvF67UjVmeWkP58YzOJrVdJaQU+uA1Kv7VLZbvbKShBehN9eIMqwWolTz
zqIYMQxDoDTm1mu/udupSRoi4Pl6waqUwgy8N/atLm85okGIBnKsYk7cQcv7BGAy
yfR55hi+ks5K85aECmVsDW+MJIQ7RxEDyN9m7ZpYcIfHFMpzBoWHhkuOyTxJUspA
9ldvTNxqLHATYCJpPcWTeSer5mV5qAPHxQCGpnOe9pPzibgfdkwUroXwr81A+etG
fpE8bRAbHxiPUwj4a4wFOm5aJbxG2Eoxx9+mEXzVBmm0ZWs/9Be8DK6Nor4f9bzd
twlgmwNGj9SXfx0ap03Hl/+ZXfkmXdHnJw5HMYLP/gq1s9BmnPrhT+gx7eGYKn71
jbr+vyjgrL8YEazh22gvB/ayjWJ502E3TplrQ/8xlmbY/e9qO5AJOy3vXC6FvIA6
PxDXJ30nW+aN/Ud4MbsKddnCC+HM0a/f17iCtUj70YkpERzYx7qGGd/0pY59YH+w
u3iEBnjUNRJD+EnVoWILuV7YQorh0BKE5PUxIlW0E8LhbWMCxYwxeL9wN2e85r/r
h/H40cN863/tQ+csGvAjBifrH1ZyPmzAzLnHQ0dxnrbBJJfOHDWDK2tlGZDi5K5F
578o5aHyK5EA3Lnun5dEOFnZLfygBlLayyd4wLZqLsMMMexlMhTf7Z0zOQti8dN3
tl2zZDkIRnAzZtYGoH0ndXt9xoMohKbU6qbS3gAQhzckL41S1uMFqhrcqEhyLEeD
MZE3LqqGGWuIFkHOxF/ZemwUYF2MX8ojDVSGJNCzYRHTr3zG05IZ6ajqJYAk6b5e
iDw3yRJFpx/qBLM7bPz05xx9716r+tEGkSTnxGrvQZ9S6oGZaa9MPM0pbxzYkFbw
BYb9KdZ2qY/nFqGrTVKfGUMrEjQVS70cgK0cMZNqCQqZAcjgWUWcL85GWG5EAVBf
DgiCuyHkfSTsttHXGMSMD3741PUeHw2MsPN0Hk/iVQdmw+qJ6Vnn0cwakaAa5hyz
3uD+x/4Af6u3dKgJEAW1s6Kx7Da2HdxBCZOjzJF4Rg+thnsmu3Zu2FrFHeSUgN6P
UwuQzABDZWFvOrHmx1pDoJ3bHUV+GhWwJdXSy5h2Ui9pyQ6NrkTxooXOc4W1xCwR
5zWwrBRwPcEAbEvZkzm7Gf1h4eDsgNH/tXszsFFsY+U3JCuszjNJX/GWVnL6RefW
+YALfa7vV3/b9JuuRubOU1m7UeHlHERAWfHialhBktgdVxer6vngV/dQmLP8MSzz
v7Jsfwt4IuC91UEelN6sMSKDHKS4nP+n5aqzrX2YR3zfIGXNrI+fEVSMsH6QARLs
jPHEgbRIsgIWcyfTQqSVS/4g+8iRrg9/c3iUDd67ZZ+/ENw63SP6+x8JNnyeADFp
Q+eEDVijzJwbxLE9lHQJhV8xi7YOcM/TDiMGJstX8iMXU8PssWKqLMJXHa5zthPn
fHuF3hWGBJNJ55UGRUgX8PkbGTRB6wE1uG+pLR3JXsyhF6uq7Y9JSDs+652F5tHo
ha1iqo2jOfAJ+y4Xl1Nrz29fTwEzWeAKZpuAXCAl4XUd3Y6qaK+cpQ/wquwfkp8d
jtpz3AGtccy9lyyT3UqbGub4Ep0qZgcap5drZ+c0TLWUIaEX1nNJS3vic75VQ9zR
syBu2wzw/t3f2cVKpGovEf6giVQZg/9LkCDrj3hd2Y0/DCVIakk/eFLy9sDKtEtU
2JBenQAHyA0Ee74a7kCOWMX+rfD60MDvvN0NhFp6Q73q6yzrWQ2V+y3M9MBJfzJE
ll1DAwFmloyZOe7iZdp3gonppeTqKNLAIRkHN98pcwauNZkQ9jcoPCVcBATGPH8T
trMbnhrkNXgReYHmwmo2uxv0D0nKFA82BPLJrKxftai5GJp1Y2/flaVPQPDyMCju
GFTceVBLx1JMUyH7hanvWx6oLNSn4gbjZ+pwkiVarhHQJiqAfStn9fqlgDbmVAvf
spXRgZFhydNmxul8HeB/ZXLHaUP55WpMhyOSZ/jeSz7U+NSPnU6OnDs7ediltwKM
W7GUqiJEO2LvF6gzZgX80phRQwflUoRZOznS715gnQupfplO9Np9tf3DI+YbhAU3
1rWqgtQe90UUOlPJVEoc+EIV5DFL/wRf85Us7lUa1c4Qy6UGxTTYiHzYSOnGlRk2
Yv77/w9fzaNPDrzwL6DXOqM9WhcZTC8IaCVO0hk5hfi6LckBECCDlzbfwndHFsyp
7HUCQn4uE+bdU2Roo/5fOsrXwwzOMOdKKNoASKLZ2PaSjq/sZ6Htw3IX/8r4WIbs
1CWnh2GFg+DaRhYhC9VJXv1ndgPVuYyZj8TuglZRRkVyUesRJ8zFLOluEpDwJJy6
zzaCueS/N8n2PrvTybeEdbjWye7d29YJGA/KiY+CY8CCIPj3nQ74agrGc+BNtBG6
nCEs+meTqmWw2E3pe391sOP2atmFMOhpxal/j03+9DIffNt5PlJfKRjKJIYQxyFf
wacJ9QafAc3VzPCdBsSNyvzIgMpn8JqNgQF9F1zoQ8iCxteHlks5GpJ0U450yCxb
01fHrGOMSlujd2j8QM5wUfuEH1qEsq06KtUOxhLNTbuRQK91YSOGjiLzmatbhy7+
RcHsiYY1RU5RuJdQpZUrTLXeLIFpFGBV8m0uQs4J2Awh601ai3x5lE2iXFq77JXU
tQFNW1kodbM6jyMIsHGjN83wODXD2Rw+Te8AQ938nUEAzMa+PzexIPv/1wlblHmW
74ieNRlwQHS5LKOUEE+PW7A7lVgIxmJlml/m5t4ZRSVEI89ja9Kq+HHMcUHHWoIN
JuREAG88tiRgeZH+xO5o3rc6iQfVkB6uRiC8SWmKT2OrDD8XflO8tM+Ow9+fJFzQ
Wcgg2VecqLDn/TIdWsG3JoBdlA01zCTDfthu4wjZ8YZR2eTzbQ/pH667asfYkyvC
YHgROV/cgkd58e3xH6YNd9pXQ9rHaaBQLCW0LWHibfvMYnBcrqZoqF2crEIe2JGs
+uEHexkky3ennUJ4Yg4IVjZGhZ7tCTp4E9sqwv/TNJ8tLmYpX2q0TqhclmVOLNXD
/Hc4PiZquEgfuxi28CgmKHvDTTOv+mERCtOjLDAuhgtAwwVMfZ06c9EfVmC6ivL/
/FDojzcePJt8fqmBuqP0TMGHHycZnTDtUGdqsAu9sslTevYu0amjdwU1Cet/9eqZ
D94k7iYsxulHSUvBQjmpEZ5JYABO/vCCav4zRpJpRMx6dhge8XpHbjkmcMUAjuZ+
FC3v1YFwHlNIZD3/FiA3/OquHveOSxGFn35vZoSoI/Y3JA0eJnidgWlPW0k7S9yE
dUqtoBkEpbWzfhp95y2/HHd4+sgzyRFucvuyLy8orcPeEFrqhKJJM6tegVyBkVSE
wuW3QHMixM3unqKOZvicZX+VQE8lg8a7ztFf8QsVJ6Ye0UfVNWHHDfQZDDmQ8bEI
7jpdUgaSFK40GO0u9r1dPEXDHITVxPscQz/B/LXVDQBR+Q7az23vAfOpYTx3CwhJ
6c9EMXQbCxPBe6f23ufNljzRfeuWAY9SA5Qx1Npi4ycxSJeo1JcfjVRc12DMqReV
kCRlzTzWVMPEY/Hq6uSSv/GnPsvv9oF0J0XxaT0b/yy6zilh8nxuwGzwadMSYm6Y
Fe3aMb+y5kP8/rsogGNH4319AhrcHys2wotY6U7XqXxmsZI8Oy8Z/CGXntTpIYdp
HxOKYm4iI5Z933/URRvMzn9EbnSK5uaX1VvUa3wowCGhowmrFbAbpwEdhe8aa+Ba
Ax34M9YcbJV947hmwX9ToGEh58qUvdY1MWWrFVZbzTJvRhcHUjQtElaf4OT4KKvV
+QXQpYUMk+2H2QScMjuNTTVlrHOvVHqESZsXCuqJGivmcJ7DmGOjti38oNu6aINC
9zkjgNms0aZ05ZBGM33F2zwc+TxTOKKTObgmyMP2w3XfTb1zF3rQbXCSoB534/GR
TmmAuivBURyJBIFz3eGAlb2dgP6UsP/Al5SqAubZOKaI5Fo9RHC5r72X2TfGttFF
NMPHgcMIlxVYbGkyBZbg/ueqxOYkrMNZzw8a5QQ70Zc66Ap1ko/LmCDjhKe52JlY
9zhrOFKdBh18SjufBKTrpb2NZnjEF/NOrPcQp+Jdj1mGf++Muv5XN1Sx9zLUl+3j
+/rNxPEKbhMOpQraT3HR5f0SKDNca8UuKzaUsCQjUhlrjb5gBfie/ZWxvzmfZ3G/
e99r++UtslVW4E7KTlymmGnQaIhHRDyOgycp3T2DdHDszW4gwiv3ptgTB5RHQxv1
aE9rrEtDG5Wirhr3OaHxirYptbXezK1bmk3eQm545GtkEeub1Ytxl8hxE94TLWTF
D8ij/8yYODRcMri+CeYwbYMNpk4lZNLv2PSFCSTG+JbjZZUECj/e5mOeqDMXlNGv
lOt9nt+Josa7kCgP/5ewwsKaWJFRtWNvmU9ttr++D2xLW1qYA4ZCOncWltVgG25Z
qiAUIJrIMVaBAci1S0IQIL2LcGEphZ+j3YkIA2KZS6aBFcEb5LxvytsV+ZWNR8ee
CR2Xwj24NeOD2R1KF8T4KJBIRArxDKgkziPFwHrvpHyRXYesJDWi17k0FvUGn491
eScUxFbnOofqiMK/ONTMPm8aVvS78n+XteKRQwowO4ODeykAhIzLhKN1nvUx1peb
srhf6JTgdsU3fLfhHvZ2EIEzXlseBdA7r2GobaOhSAueLW0G4ZbGC5QAY+ejuQdK
uTBeg7Nk4x6JRMXfC8f7vMb0NgWtWR87da6Td5gzICZKuuLWf5WSPOr43d2ESmRL
kSt3MEFx7pZK+jMxZtDxh0KnBDO8bOwW7bMFqR4Eya9w4QO5GtJDoF9GaYdJNhKM
X1/8i7xcfIZaAgGj/iTyLXeHv/MuVIBBCjK727ek+Jw97kJ3MBAkiVRZfDOfTYlk
MBWf9wUUHN0PfqXyOvWieZgXyU2r1DmBySuBpfkEEy7+NxmFqN6Nln0zr+z4Yhcm
7Bkx9h5ATL6rkm+6c0WBygDOLKzHXbSWISIKKMg0Ch889PVmsRyzG12uosPXg6l7
VeH8HGgo+SJEkIlAGLsXntvz/Wt2zq47CpGOVkw6Y1/BYsymEMusf2DV0bkDHVKS
hCmcIz3r+XEB+slRca/ldlAZ69nTtutj3a2SONiCyIdbR+15YoEQepy9ho9P59As
y09AZy/2mBEbbuANBG5MZ7HaP/ZGk3orL/pjfsNqOfG5KYtLQe72E9Exj+QuWe+x
q8EJQSRvce4YrRwUa0iz0dq9DyhSDIekwUZZemDRvbYpeI37cMP4M3bAmXoP9wgU
L91CW4GFoncZknueV5+MrAJuftRW+tdIkmBd/AWuS8c/V0yYeacBiQNRBGYOkrxR
AVcLXBBdmAlxdft3oCZ7VbIXLaUdEXNPedhV7alQoQhX/8soGvbJmjuBZZJzkilY
97TPtW3s0+FB16TSFECqBJp+AIrHIg0BfhquurFJmEKpR9npAEp5HD5rZQ3nU810
X5DlwTSgjjTiumn4vHcp3bTBHYRlFbKDmqG8HQ6QWQn6HtnEYGHup55cih7D7YQN
yVkt9zlT09VF3Qo8EXtBFPtkQCDW/c0rSO9jBedwhc2zyRwbmqLUeC1Cridtd2n7
Mec3W44el44rLEMlys0ig0SGWcizbrWT0EXY92maKtVwYO/MRS38PKHAsjH5a6g+
G5qosUX3djPmZ4EDSMOJVelLR5Bmj1Mib4/mdM5YYBkeTSqxropipnr3DADVXGxV
GYROjFzNRoqDJP+UKs3dNcOfY2churwrkOU/71wqhBaPgE/FfYXG4uf2Q3t9NiPm
P8i1mTL7zv3SKfVzd0yHtGpvK+WJVs0oWPY6jdFS8HZYcYytFJ7a/DnYaZx19w/s
Qc3nCrrDc+HuQxG2SaJYbxZAGcHcvVldlGE74iPClq/QEDrR4Ll2+sEiucaRMH3N
3N90i2qs8vspxnd6VBbavn0lpOkGJvn3V2Fo80BMte5ITqJeyU+i6mvTJieX4gKO
gdacUf5bHsTltEZnIwJY7ulSTldPpmgqFPVlOAAoAs8mMRpeEOC0uQgrPGRBcSH9
rqebVuEaPiC890O5byv3HSpctFy6glsah0aamCGxnCUNEee5MqqZ8IMEWEIz7leZ
HJ0A+I5hD5zvrYIw55oTborvpZZkVpagiPTrAekIyR3fLSx85fN1UUg7dCE0fgjv
ZGkmDKXjFtqdRVUW0hY72S96LCWaZanpiSA1N914wJuPNvELi3OG6IQvSVqVksv4
MnIbvVMd8798XAfU7yPzItYk0YumSPKLM0zbr3AmYRHjtp4PyyEsqkvHOoErfoFg
5cBO9hb6t29pg7kkHozdWbkGNfUQtF1rqBZ5UDl/Ed+yRBPGrBGhvka05LG6UdwZ
3jo43PBIWHfPNYjb4YQqZmgdKuJFkP2wrxk0MQ8a3EdpkaLii1uFsofWigPHuXNd
ns3Wp7dItivNPLRd8p89gWrgAcD48PZ8RaXj3Zsx0i9skoZ79LCJ6aSlaW+pdnce
ZrgGMe1fDgK322IlGXVioag4hLJFsvThGPqDk7lweWBfokYJaXHPHIL7RyO8DCed
CUeWiJ9e2mFlPxWH6v694Hw6EoYxVia0eN7MP4CqjLkECVxkRkfG85+/++9QeURI
20U7BOgzV/nbsQQBEydZh8205iePyhNI65NGRdASa1aXoUwzeocM6GMRhTt7Q+FS
aLXmaFS8rUnxSTwUULxeJ/bw3Kuw1FHfKUar8sp4Sv644TppXkjWEe1k2Mmmi1Hh
kHY3lRywveKk/3IfjyGUPxyjFUqx7XcC659J69JKauV1f7sQMSSLEQN+iBAJANYk
Qvfq55qc++TQEuuzwkoS+QN0CDg4y82ihipRpkHuq2PZQlD6EexacljxCHOTIbj5
h02uJLUoqGUMf31UuL4bTqnL//y6JymNzXTVR3WvUPbb9P0w3v6ooQHBCBtdDxNc
PAnEZlxoF8Ef3B71xedaftcQPXewL2lJUym5ZXLU7wvW98p6VloeOLp97hM8Cp/E
MaQL3c6TpJtwE64/zHxNUSgkxqAeKZUAobUv0l5Od64OSpKhQ2ZM08c/hOMvcSa3
dZXip4A5i3PbzzKRMNSpv5RxpSEHZmIYv0Bp2i6cmHdtkXOZrnJh9HAi/D+XY6P6
clSuBfuB4wnPWLOSdXA1uh2/3PaugsWrWSbwMCy2QixEEQelLpYu39X3z+lkVPgz
T0d4oK1skhbGTvuFOyV/j2PAjQmbYvx+NDJeMy48/vHqPCOQmXfZYzoBTv2j11/C
ySC+sNrtJUHFuoaeC2ygiGIhFihOhFb+rbHoo00NRBUCNCFf7plFlGRvj6WlHy+m
7tIkSofqz3zgrHxNQEIcTYprHiQGyx7EledPaDjhiRLg4WgCbseknKw5ztvwL2RH
uYvzzyjy14toikfxHCHuPzeoPcMgrqjoAELIEOkMSj7jA07qDiuqxr4ilFqDicUv
2fNko+OQtF2CsOPReqKWqmhGuca7zLebYMqTWH22YImAVUKOBdRHjpmih6NigeZ1
3cfhLmpb/UC4RyGHfH01ZXzxIdiBcRuFV0/d1bsBYwoyINXv1De24H3X53bHSe3G
cC/K7CzCgRnaz3ZS4/DeYUzVodRsmByrIi9VV7PPzN+D4kw0H6gMnK/t/kNKBGXY
qCiFHoE7oLUxdA4/WPqzzp0UV6/7frPTWI8LO/IGSnwSDlq130vgJcPG2N4bwwdS
Hj14VDKhR6seTWABFA25ecJUL+QzsBVtY3rNZ4P1OjBBjpn2a8dyzja513+9hzPC
bn3Z4KX1l2mHk8r7dAfdiU7+mqW1aQaZqGIXDjjVvLRun+txZu5AonIBAtfaeJ1u
xMUfoLLtiQi1D1+bU3SXkVpETzxftMY2ST3FDcHzj9NqEusIEjb9zLTqSGdUf7bt
FE7NgLaQIe20sshthkNr0+Z/YQopPAA4PAz0hKinGDnu3TLpN6kB4PylAIgTN74x
1gf1/o7SWw2fEbpJ3FQFNgzVe3lXnjWpnnG6Gw9zan2hNRyt0PIer4KWXfztV8ZV
sQUk2PTmMhqP5jXOohIi4h0D6YyYFvVAZYoYOx5j2nwe3OYQFMcb0TaQxiMAjVmB
IXyqos4/JA6Wb67vPN9ZRttUvNug0h/iaRhtniL/1AZYqSvo3SzCNq3yxMg2O6YT
41c73L+uFBpvorv4bHjgiKpEmaOpCFtxtrstbiswPOgpLGrcNIq7kNBCiQ4F53+Y
q6ffawHPSvMbx6p5/pOdUjWmX3IWDMva1ceuP/I+hQ9RK2wQgGYZ7+WbbPXfxnC7
pVPGKbttfmbQS/28KzDcIys/d+DoqiTb0gDHOwKpYfEBV6W8r/AHzm1P3k3zDDkX
6fkgBGwRZA9EGQQLIfSjJFv4XmGjfaFHa9JGpT2R/TsTncrS5XalKMN+IGftYjGn
VaoKB1rbXxYuYkohTyHILVFuRuK82lZCYhahq10S0Inzu1/fW8dMxQGZT/gMMaP7
FLrjCB2FULy9JmTpm7d1QBWRbj1+Mx7/NBr3k8CYE72Zc/4m2gR98TuTfoT/wAKd
r/awkZDGrMUjjYBxBQcHY+hTgPGxzP2EuEEeOaqAOPN1CU42IOHXAfwFqyu7OJT7
l+ZuDSPS/7lK14pNx9jIhPn84Ke4Pw9kQxli0789Ntqi5v/45b3E9Diqb2MQbAa5
5FfVM0QvIrtL2UQAdfnX6Ud+KBzn5l/W/PAqxNtMwufd89mIZ6rDSTswEzvH5tAT
6Bdkw4T/AiSibVzhmv2Pm63omRoxCJXZmUGYj+AUxgtZUuyjKqW1Ato4Q+WGuHpK
5t/+ifKf9Xks+2dvpGJLF/amIXEUMP+XscxJuZRMNOmI9IQnHwqQiraVGyu+ARrG
6Z7xO/eUvSkL2iiPs//nFZ5v43R20K7E1e0LEPsytDtjD0VOCF8h06OmcTjAlsDq
/57vXNR7vrsSnIRUNvzMu81p0pKylHHFajGRbas9O7l1e6OfVTKbcAXUN87rliTU
9a9w18fZj8NDIkO2R/giV6H9eazp1vIG1QjW6vNTG8XEDLJCS0P4xiK1PCom4Vp/
e3KVq5I0uvOHJqHNPaPdHdET/z87siDyVkWOwBLWyAJYNvQEF51rHR/AF7fbnkQ5
ohTaHZEoWthfVgA57w0tp6RFXF6547dM12RkwITzNlbtLcxM1w9K0maTmoATbgYZ
mSmSBfVeaXaGzr/jq6TG+NyaO/tevErO9UJCXidIG6dQ8xMJmUu0r5A8uIGUBE+g
60is9O3tI5WIkymgNuceZJ8/Khla9S7QyLkM3VYmG8FRhyqQNeRLzaMYq2DqO4N1
x3U16otuQT4InT/zlKbStB29QB7MgrdTn/CT9tJzTX0/13rCHF+mcWFuEyEej5In
4ICcOEgZCB2yzvUhPyl7FJ50puBwdPga/+zBWAbT2+sqiWygLeOz9vDxm++M6TGc
zXKTcADVDSaVwjBtnl/U7snd0AiP3hpZHmW+hsOm8Yvpdifbiwamb/xK/3jPvfgP
vhqG4DJV+aPww+/n00788+/hFfKiTV0inS/K3/Stk1v6IrgP7YX2e5S5tSllOINU
LbXPDWqOON0XrdVX2EPHIPGe5GBSLOzoniLpqy6pCuZLXD+htGiemA6rTfChBT5s
8UJCi8dbYQGYJM0F9VgGNGZzrB2Iqfm7ekW97tPYYrIy06si8cVPokDE4ct+TPtr
HXlQotPzF0Er28xSy2RqKOpjQxkMhMUeM4TbtMkuZYYdgbmK2XKxKlxVU1Kjmef9
UOFXFqE676df+5E45QyqYaZYwSfjTB1C6x9h1hRNy23N9rbjeunXdrMiaj0qrDhq
41+oX9skdQDSZxYF71/1t+3zmHmdHkRBXM9Hd/MWmTgEstbwshFVMH3v/QpEhSjR
zuUDWQ6O+ALIlVZTAK6Ehq1t3nWijntkP7lR6qgszArp2rEjFlMIFIS9n5efutRr
2rz3XZAO/GHSMz1Xhh9CweRFu0gKLzox1vYdCDvYVcEY9B9PaT6ygeGsEVUJOcvM
2R0b+/+kUwK/ulOg0US6RA6wuhbe3rGDgngWL7vxG4F4e5Y6cO+8xAXxy7uVvcok
NhopuO1hGWwG6xcn5Y0LklvNmFwHGLkm6lKZNU0u9+5l8Znz6S27AyTbYviStt7w
BpMa80XyRcrnNhrhHPMuOSQnkAf7ILXHtxZi4dRU4vI7s6m94cMp4k6dX+LiD6EN
/Ocy4shXw2opvgQgtiKtWsa4Br+19Spwc2eXrWgG/5uosvHQHNaTA54r/TmLEnXL
UBlo2c+GJByRvwYksVITPyR3oXHGB4Ddwrs5Q1VW55NsWuVZR9RjOIobWV3R193b
gp7c6TjApL1ZnpxUSFmJo4Xazrj5+UeTWybOBFqL5XCB+T/VEXmkWC0zgghJDnIt
UT9WqsmqMvE1nPq/wPjUZVttt75J25VGKQ3H0BZKwmTZJdTQheAjNazRX0xBio/W
Wf4bnUh8Taxs5BvY5eHaiZibvfzktCXEIfqQH37U9y8ja8XrAqnKv1+kjJtAVN6v
7vHeADqgejelaGMxdqre+umt1CtQDEZ8oZ+8h0mzsirpT/gs70NQ80daBnJi2Tms
LdClh5Kq8xXu0BBrQr2CpmsiNJxlLJNM9Vfdrk0ntAs5jLJ0+Mo4QG9Fic7v3IKt
J3ZXKBk4q/u292rPGShw1yG3dSyUWHWXSG/e1NxIXN9R0gWY9T5Pf6XlSQunJdtx
3UMHb7yjRzTaTnM1enLRNqDrnoIys5YEGafo2GSlTih5ecxZ45+1AlA67gNfNleo
BGwcV0FPaWIw1Ng3vJkJW/BAW7Day89M+EuGD+CiXF8sZIIU9rU+0Gnwl+ss5Yfu
QaKwFZySzSKz2fSPP7xNDRaG38vdml9O+H5B4rquQural53QyE7zDvgTX/RlY8Hn
vfn6eEMufp1cxbBdoAxqmzJcZtd3MwLNxwZppJOGTAyqIzV+XJz9ycHWDiBcWxtA
pSTLdlzaQbZtP3hxsU3dZiwsMWpE4Q+c+vilgu+I58L2YUT09EXRXn9eW6LPy4qk
Y5jQtuOVLWUAUCLL6UhqPBzX1yYIziNTUMrEtA9rkK6bQ0nNlmNjyii9igejbqEL
k7QRolzHSd4kCy9kTVZUMekum+kF2bYwwz+RR6KzNgN4eQCYf1uHJRhc9fMGxYyh
ImaReEdxotOYjqiuMa+UpDqxb0G1BYbf6qPFv1K1OAU=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NpJIjpcMb5XWJfM7FUHjOCc/qJEmfZPbpCOm0xu+S3Sh5R92zYC7GiFYF7d0h0lg
jPSPGAMPY0bV8lBMeMqlEVCx0oLmNZghZrQMjNbUc/15Dj3mNdr4nGabLp9XiGdJ
PgiAC2+stZaAIg7hKQ8rn38WWwaOjpAGCM4gXg/BJfTEutu8QFXhUyWGl0gX9INu
Y+TxVTOeb1RpUR7BfJeAG/PgkoVb7TGWjvc2ntBpToZ+BYvF+e0MvLZoo35/Vqcn
rR2oLkiFVE+TqSx0HbhG8o/y/Xgjq5YkGadgdv4iVupgToZi2a1mqjao0YLKPUZf
prCVoc8Lk+RMJ5XkOxMkOw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
5D4M685NYWo3UaXWzrDDJab+ImQpttQA5qwbac/h8oghjMc273Xs1EX18qbBfs+7
XGhU4BUMVpmJq1n8fmJaKnBwDd3O2iL8BGHtjhzR9ELjJl8qAPZmp6VR8I7mgnG5
Dgxif1yTFDMJQT8GToQgCPgeb9d5G4NfWkXIK76wXOIOV88IOwgsXTJkKIXsCYTb
xoEfl7r+c7yFPpTE8eqM9x/87UNLBDgUgwl78CfTPyy1mSMFmyxkSbIq1B4zT4N6
nFD/mdxJ+Et8G9DjbzPiW8JTTsmiPFTIK4ab4VoywqpoDW2NHeqLJbvX4DxPLiJZ
aDw39UdtR5wmzmJMes1ac60NGVmkKSG2TZFLQHOz4BSmBkmGowzY+p+ErHh/EiPD
HNTxKvCd1EuH3wAk9sA36tQCLvUWqzbNv/ktkwZ/rxBTwePE2V1TR8bxypLv/5Pa
N2Evr5e++HwKLC6efmmt7FkaKqAYtrXQotZtmJgzyVq7e2JZNIJ6oL+r88i9Sba0
Wjv/+Mp+lBqbBuV+va60actSipCcY08PurvwmPZ67fvjlxXgXqg3Un44rZBo10Xn
RK418iM7M5P9zaxSmNG3Q3F6hLNb5ki6DLBKN7LJE1FS2EPNYvYERFMcCEJFyyyL
fPlUEE458ZMfZox+1w0V1ttwPpdJCQOcnAZ968roYlLKXYx1PIY+Q9nk74hdqiz0
whteI66QOUt2m8Y9mwNln97QIFtufYGJLGWTRWBe13ij2vjPCnoAsV6qjvlrj7YY
Fv1LC9ntXPBJVi9vRoUi+bHzNveC0+BRowcqaM5baEp7lzgkkJnQrJLh1ZDqaxgb
n8dvhMvONXmKeWhW4fbOvLXo+ebILqMfRo3sa5JxfSrgSN4j/73ww1TMLiNIhiuw
2VKlG56I9r1gRglMpg2G1JPo5z5UHMip5xDw7VaNIY74pQPVhH1IiYxVP/KvqPjB
FVnWkaODWj2CbxR984eKP/zPFic6nB16cBq3n2kSzd1cBFyGI4zT4TN525o0LoM7
Xjmxp7A6zIFtbx/utklSEx3gERys6pcX5m+XTJTdJB3XyyY2Zq+qh0IictxLhSI+
jZqXNiujx17ItLIuK6oMI3SYrhTZVUDk4+oynAdx9IIDT0KDZvBqeiy0AkTlQVa2
m/2rc6bNWYgFdxUSYsiq2U81VG3c5DiMl/Y3THYmtYWloouLwQepgsRSG/iYtP6F
U6sGo2r9HDX5sgFnJ5SVwp+KJNNBCG9UBtv1BHFSyonTdl7YBL5skCe4O4uzuYhm
hQ1oeagx1o0cBTr84Gb0fEiCgkBzFwSvEX8xEZAq2iNyholem7wfgL2NzCcyU5Qr
TywA9mHjmzMujKWj53xk3pFI+qj6XxDPut3Mlk1Vnr/DtDa3vDRmjaT5rMAsP2hJ
R4BX3OphK1ngSRj/vedw6ljRIzEHihnQi9prqblt3TfYOegf2OxFsx5qGcqBz91D
7wda9C3kq9Z0gjcnqoPr+r4KmCMPTu3Iq94exybrqdqXv4x2gg7997qcbX3BwXUA
ecz6a//r/kmK879t33sxC9rqiXqknTECZBegG6NUIr96HZTv+mMIZbGzQoYsXYkr
BWLuhqsk3uxc1q0U2OKbLaDsTb1RH262UULEYdlPo5rWzIGMb7N67XbjwQdEE08r
l9lsfsV/WKPAVnSFiNpaRWvL/3wI/waKj0l9bm3YqqKBQ1rE+OpPnV5xcvXY0Pva
h2z2LNg54PmcOxD5XEuDmTjmuvQ646k5wigLES1DC5W+DhCBls/iqGjdJlkFSt5S
IUmSvuvOGK0i4Ga72kmJhlOdTwrSeb6BGbPaxy3YJBFPwzpDcBMaceOkNzp84rTm
F1jq5GfxyLHwPqjimjXuc4xs1DoHMq38IzmcwbIlEtZBOowW77NZ7dYNARnuVNtF
dR6OMHiX1AL131h1DyLUAyyP8bkKaz6zXfFd3/Hxp3aPeVJLRsEzMCLfJZpNWKlR
9MrUIivtDHOukCs3TftpMA1kLlYlWFfZfNSmvarEYUK1j1Bfmhyj2B3t2aVK1uOs
Q6aJ5GQ+TFcVOXce4o/H+qlObPsOSUjrOXhI5zkOCZ4UPsupSeEQFX21KpZszQ1v
Yc84ItiFx5GL8JcjMbCwVF9DtpEKdjO0DmD/c0lhu+U7u9EQqJxfUyoPJUzgvt5s
hYkCW5UoiWrtf78+u43rPIrBe8cpyIdt+1EsBOUMNg9q6L44HabKFfESD+yPHtn0
ADZ4e86YanMJtLgNwQQvNTgd53hIt8uGex3Yo2VYhtooV8A2Y7SoXUHCOGqEKxqs
SNojCdGrb4SrIoMp4vW1ArBvv8P7Kyjm9KWfLfj4QmfmvuaqF2N9KRa5H9/YVgKe
J8ewAuvqjNSKI+SRHrxmuCIfLI3WmO1pAkaAPVDuZQ3TGXCGNFZLr9l9T8I9UU4l
ytDVq324naIkBNGhFvMiXiPvfkJTK6kHBNL2n99R4v4puGXUlR3kzXmrPwWReeJG
qLi5fr7Aj84oXHF0HhFV6ZSSUx4AK2z2Y1pM7t5dH8LJ+saXyoj9Rdni41yC5RBP
lAoFrhPJ6Ff8saErNZ6j0n4ATFn30BL+D+HUxWsBPp598+qSBXzdEW4HlT6okHjr
j8XfB/r7z1cjVZnqscTzavHjRvC3wFtledUZPti+lkA6ZH2REulEbguDja4sixns
SYQ2Xfz752zz1+9a/F4IvEcLZuxABEdwyOTuwWqGgA+QxiDaM84CwvdpNvajco5f
PHVuyLdftmeSez0d0kh+4g9d8gnC0Y2P6SEm6BI5U4Ayg5EiDNRqIFV3DJknl91v
+89zXVyqrzwbVQlPkO1Pr9m2jKPq150ZeVUoBZXz3l98wTKSEzCWtRh65GWd14JR
oa0tmk2vZkTE2CLBb8CtZdjY0ZCaPhRaujP/83+1mCwvk4HXctvw4ngrKQbm1EOG
quwIuJlhu+aBV3ExarDKfJVei4SQYydG4BSnipRkmo5fwUme0h235eTXyzaQiY6y
flWhRy/zGIv0UEPcNe76+itopJ72e+TNO/sn0Gb262rHOkY2Z5LLaU0UEnVZbQCG
or3bl0M2OKuES2jC+kWi4+6nZfinxKv2FKEFjqMFecuxHYuF12araupod+bF+V8s
cvLC/XHLJHCgr+gWT0cPkHu8Zxs/yjtqFX+Ukdzma5+mxnk9buELQlH214nfpbem
9jd6HSNOox45pMsVPY4ExsGwH3kYvfbHLR7jkmOsNI4MWc34OaOq7OnuoSDlDgVp
s7M9OeFYcIYBhMuRixZHf4FaPQQndLeurGM0WU/0/4NP/d6dVnQynELFbTtgdO2p
HgNXImGE6O69YfAEUuEKPJGfgzqMwjf/O5OzKWWA3VMFYe+aa8puXr9NPJNxyclE
/9kvdot1OP69WtutYYUPx5PT8GOyv9sOrZTH132CNW4h/qAifEV08/gY3rFXaNmG
+8W0Hh+usFnwsTaXGrBZI6rnUf1mRpZs8d50/tPiJkJjLGa2+1wKzFPLhGRBMkOY
4Rgv63JMkO/YT3ig7+b+A0/H94S435D5ngycPJAp0khoRL+AsqCLObqpjErIy4ZZ
UH3woPejDKQYECLBN4QAhw/qRGmeVocnIvv5VJnCJVopYvSXm3iU41UkUVsL3Yvi
hwQdRU1KAfceg7FvFrxIu1Q9kBbM9UDrnzfVcJAYHRLKvwSsNegPDmqQvnQ3S2mO
nHCp6zAx2hs8U2DrUveGbpwvdKSEszKdVHyLSfCbew5T+GCSVmOUMYgTQc1DP0VD
B/9/HzlIEhpgmXvEBPgA8TF1kZKlpHDIDwKCNS/OPuyAOZygN8Eg71JmW3yiabGk
f3tduJZoraqdqLjPfqw66MlMgMMSMSl4N2NEgTkLzKxw1HJGQ0x9odIYZAYal6os
Hlfy1lOi1Y0161WYEJ2XaM/Klir+3TWgXbLKhpNpshX8N7PLAvryLIBXaC4TssKZ
xUetRK9FNUSucfqydsFJKuxpy4Q+zBaTPsrta8zNHbRvtCxx31DSWmcP6S2kL61R
s7rvdnsG6WW+ksek2LcPh6LNA7Nb5lmgEymXZZuzjzZWDKy6PdPvwNV50oVFvXNF
Ois0NHIQIliXxH/u9aLhUz22vMrqOg7MO3j2e90TzBhK4Gy5WGdyrHNNESCWm2ld
fdiOuzOiBr2kCnB16bZd45TMMYpC8rGUozHiOT8W4rKD0Ou7rzPPBtU6VgeTro6f
dLU0Lm6+WoZdSvzfUAG/WpMUQDqP3u3qDkVaRa7gKMSHZoufLo9jy8U7oylWpHBO
pKKfVQsYLh+SxoIEI/wazOUbMNrryDAYH7qvqyu4yKzMaxSMjlkE9zpN8zzWW7jG
L/jZCb7ev/cUEq5BzjisGI+guOX7e6dSWJ2L1I6ZJ4JaCRe4y1UFT7WkbSM8rdKI
9uByNykJjOzok92blToiMd7//CJYihj0qaUYJJMfdBkLxCOrVz+xyrElrZjcOAH1
OCQeID8wCB7j9fRg5N9QyLd483BG1BilSKdcRT9JG7U9Y8Ax7euEaQqaxoixGf4B
v5uXBf2dzq6SvIurRdEeUKT/KOmr9J6Zqd1RSkFsiKZD6wgfKF/iJWd+q97tofC+
wFZaF4iXYX+8gvNAV+G0+0aPbmJdXMMqE9S5RC/tj8G/AUd7HjubL+jUQdHrwlnl
nWNdb8OcSj+PkeQi4B89MWk57uvKYJfqmL9JxO+C4RH56e6y+plpmrQ5hlFHAUzV
qZ0ZV5y453fROIp6qI/A+u5cZMZLmZ9yZIFfnQWLxNMZz1fCS0Xs8W/8To2ABaLz
pLY8eovqlHW0gB/jjvcBrfamc2xXI9ZFmgmW3G3i9iYADDE7A9+Ut59C+yimX26j
pD7lxoWQviq3Q4vp8StE5xmfByYvHoOd30IjfwETnPwhzCa/pP6fMjTp3R1eui0m
MMP3B6xvBWt/T9z5mA3FMK8Yd+3F5y45RznJk/5jP46is6ZotpG7iWxqycfiJFXG
NObiSsYnVVbm0o8j60ap9wjTx1oVINs1dEmHXuhS6gDhXFoOpBHhi40VUunByoVM
IqL4eEcgjsh/PlhVenN5QFyQq8eFkLpJXCtmeHYB8X7RJXlSmYEbGBK05lWXC1sC
nkz7gVNbutJYwD+kl6tBPyl4tzZll5S5o4py9jv6wCMvrtpLBI5wgV177Bfkn9V0
IeKW+s1saofMVxsMclvPw4i5twxnwi+HzS0EWd07KZ+9nnDQrHcpS9TrH4Rt6x/s
l0lNjMJ1A1q0KO1btKHXTTnckXO0aytaFLoKFu3vjCDmSDN28cK8SF/Xe41OhNSp
ea5vgKD0q3ZOsyOOWYt5VFvfPOMDoi/l5OoSG6ueOJo509dx+676hrqVX4es+iX+
nHrHC1RXgbEijH31Aw2gu7ToYz7sXna67hi8aoTa+brjNzJTMWD86U3CrpzEyQq/
+vBROpJhienoSU4BuaJdeTixcRHNv+vI29GJvLYe+/DjPuxIRqA8Iy/t6SSk/zVV
ThBy4wM6EjbWO9I0AoXaSnRn5AcMYxk650hg3auEsKRPQpPtVg8wb0ukBRYvjiUd
kr4LKC3unciuzjP+pdLnMGhboizRuKD0yjPrmfiPXMzvb87EAg+UZ/XAtB6WYt84
blVXMsdj/56pMFR6/cCnfA1uJyORud1OxlJ62Q0rQbU11HOhx9A7LYpGFPG0N0Zn
/3og4beYnoNdgAAry5uAFG7D32viihQihDEvvpF3lxn8GgvR1Ma6p0KCUAP2FS2L
ElbqZ910Sia9zPIpvHe8AML5phzHmdmksvPvSlM7h1j+IIrassJITim+ZBUgB4st
2fo4qiWM4qD5QF0y3VajEGjWOgRe6MMH1Nf0MgQutwE74895OFzoO/IiLmh83PCo
rjbGT0oI41g3HGM43lWbFhhRr92ra069gI95UeyfEd718L9CwIdXH0Ql4Mvp0Ji7
BMgUF6vScOwgK5vO3loq84Cmq2VkCyBKuTctSSm0OqPaz12LK/wYRgH0AnJaqwKW
MN5LFCVCpz3kvxUnk/k0l4Fd7MK0TPyaX+e4cFl9hp7Cy47u2uP6c0gzy0iQ7Nol
9JYDiqUff/jyZ2vVSPF0ck0HBfDdOygjwKW9cuwFobqOZxz8MdZLM4nDa0Bcwyq4
EtwvEbsj32wkKqD+B29uaEMUZh2Mh6f4QufuZbgxcleQAy6bz5IfHESwY/PIyZYd
YVbkK0j5SQHmsAF5GsmxothsRwe2KN/uvNqyOlLjrnLFlFzSwfHEzORfBDkp0mcM
zRAxRgnC+0u5okM2s/8CqTBayEC4hLhpQ3/RWPcnKTWNPAojfC4MzYmvpLDiGmzB
vXqOZnTocBRYqwRs8ebgNo9pzx37R4jnAYnYGnAbcdi4i6Xq83P70k/gYy/wtsR3
7AcDXPEITx8y2RHGDjfY1ds4lS75aenhFm3d8yAfvoL6Thh9JvHUQ4fTRjfSHwS5
ffM417djuN9k0MxD3DMaiyRcvBlSwy3D5lIHBrDZjuj+x36+lgMrRuSlkCenrqAg
9IqbnWu8SXghl0pbhgcikwKfkKh8AreoTLwIx5piUuFoCq6mJEy0S9Jg+xiuHKL6
gDIfdB82ThXTmWX1KhcO0YgpfaIFjSSJ1akqLFJTCBFc06dDSUMtYlJu4XJ/6UqO
2tvpL+j0M1o1Zz7VelO1kPY5lbyKab1CLsT+u4fP0UIBtQx3IIAPic4cCql9oCAA
E56Jue7HwSPB+X5swly93hoRUUeZDMG2wOiDqchyfZ4/7IWD8THu3HfdhdztSSHh
BhuwIG5ouzJ/cQlcQeF4C+j+e3akO0hZKBqSlOx5gUsdKlQyA8vQpwyeZzdws718
Wt9wnq8VOudOemf/rV1FOPHg4DdLmHrSeOPP00c/72REJTE3yZnnMI1loAfvPjEb
kxglHJqEYtEa9nDcHUi9cmchutrH6WOCRyqeDwf4vM4YI6bUTgoHJ6sitHeYLS6L
X7Q1ll7b3VjZ9e9DuWTEnrf672sHhfNsyztB6jwT/HpAZzOUxoBgsjpbDQTuAB5v
8FJXy3aE8WGPqFyciKGEZko+x7ks/DGcr5vuSrougqEoaBnut5mQJafednEbZvHL
onJOJ1WEKQBQXDaxpN2vz10lOoUWhKs4+YTeA/XZndpfy4J8LYt+QDRYMIZXVOw2
xF2RQALfUwg4uzjW48cHOd/c3e2uRH14lg+yu/pLCypv6B7emsdSNwVgdioU67h/
NPeyd/AxS3at0V2D0kGgSR2RalMvsgXBTE3z6bej3ME6laKyCstWekgyYaYfj2dM
2hs5d1jHd3RfRfMuEez5kOEcwiaYtMC4AhvayLYjbQ5tJEbX5IHIA4Ybwo7cmZK6
MFlsgy3GU1IUVRQKMmStjB9+odzutBDWye8XzPag/f1kn2VxGP4v7bzoZSQNX8fU
Jye6HZVLfSt8o6as8CsjBxM86JkJpyk7btWAw5UWNOlYaU1K8ugHogQVYgd8X2Jn
T9dyRZoei43axvsHNu0Lt5wzd413TGb/njK1JrTL+VGVv1CggIkg+xmclJE5e4tn
y3j9cxaRsbP8Y2SK7zP0JWPdgvJ9o+1lZ18bvPifjSbF8qlXRvkWfDAcdIAimsV2
Nni9FwO9NbKma41MDMNMaNm0eiVOJ23mJQTuTxoU9kDbVjsrlDJ+eaQsYpu9LZ8B
VaaorZhWjufavxp1haaXneWRLjxk3jaaMDkZYPubNbl2L203+MLV+0NG8orpgdbf
cKh8Q9Uwyuqasn6JhRwk3PKI+8DadNnWtI2EcLDGluB3RP/rbn0Mbw/bTbIWkjU+
CrbAG7kb9Cv/4CUznZBuUFnk0VpGaqCVlWofvGehyfdCClaN7P2rD54WqZJJ6jNt
JF+lmGBGqbdxcH8vlpxXNpHdW541vY8Ot5vDRDvt8Q5RjhYzDnpZ3/41uh9q2JeY
HjQa6wwWT1fs+087yLnolnC6ZQvlTetpi6ePxp0ZDOZcrAhR0g2jbWYlrBSoVFLv
l6tYKyRwHzGOpdUEGuk9kw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
d767t8CYeJvbrdJ/HMkv7PpQHNYVc4qgxn78eBhBCztcu0kjCsFP3xbH/TBYqKqH
DP7juUaWQ06Cr1QbGdWMWQHQp8V1gxzWZTN+Bbnwh64pdwvlA/FcwiCmQC8xiljn
MO2K5sA2QMxHfbcSRWZWl9ugqQUOdkTaH3MGEH1Udv9VHAl1xW5fM03pJj7p17D8
91Rxpdi8r9xB2GvjEGIFOhI86d22+oaCrTTyAbkYLtVrH5M6dctek/TKD6q2/A37
MbHz2Uiu3Nq6632sZORSGAlFcDbWdFSzmiAJ5Eq9aHjbQyNWS0nwWmxNxl1ObL8A
9AUzUOFUIFPBO1EeMqWb1A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14480 )
`pragma protect data_block
mSieEmPAOYu5QoRUOB2432kuo/+Yhg0I0l8jLIsFRr/SkTDCEb3mt9WHhZ5zj1iq
nizF1/nALF51E56ooiy4PNsCgkakgdLojIU4SyvGCABb+OUBw/pCsl73dO+RyIZg
RwiEqpjgU9b+0oaHKRpXoXPIlsKdhGPhTE7WA62TPH4Sc11AZmq0Av0iBSS9ONEP
9dkSJko1ypbqVNnCKSqx2HAB3vdyBQpBNybRHuAhQz68XndFJMOKFdX0QcwKAR6r
QicrWYTgMyMTsPFz1X7kvxL8dkRxezsoe09STp9NKbSmcnkSIWRgsiQvI8BESvC9
RMJK9RFdoVVN9gJoGhmsdZ1b1g4fiZh5Q+vpsu+A9EUDb047u5i/jmffaR6bn9hd
0kHFRU3RSo2Ilr9CRTLzhn1mxaIL0zZDiFYT1KLkR8tAAcDcaBCa28UmpsDoMYgw
tV1fMPaaURjbxHoolqQSfZ85NdEdJI/syf+L0S98r2qM+Bwf3RDdrFyadrdFAJXx
8xuLrzDwVPsq4wumDqEsHclCgiUPPNoLcSenTOSX9ne1Ch9JI18KDDtJFWvYR7Wh
3yYw1j3XOIm7JfsixlE0MrkMrFiQqj8GZu2TXDgN6g5cwdysTpwC/5QwLrXlKsZl
TAfrDNjkVWSATlTWoVJ34HoebwqB7HZV5D/sgJaswrEj3l3IbkHQl0lGnGhe7PVX
v03a0XB5RZjmqJodE/0zeNIgaY4/KS94s8AK8PgvZeN09BuvJIyuEaMx/lDBrRzg
ZcgL4yhai071X504csNcDyPOPmy/ZZgm0ff/jbAekDHxDhZML8481cHS15VHTyuV
8R+5OeW1UjZrIIj9tvBW/SfcWYx3QQzde0KoRxHBn8Z33LOV38qZu4gvZWd/zfop
dXYvlvvtTL0XUoBhwLQsVUp10umdQTLbmANmjUrpWYkBGk+mAr8dIshZ9gUosMPv
BMFctABLYAIOQSBcA3kK33YaTlbfePtCs5LSFoZlFMjiMksgFAwyMkSbPnhkHahs
IBMzptDQrGeMyTc/4DNpbeGGtgxR2Qt+9TPxWZL9LTlCIbW5UbeuDSVr1R6NAJtx
B4i2GxYsEKinSO3O8FBfcRmwh/5YzVvUyVtyKCmhgxt8VSiu6ff8wthqPfkq9bCt
QqELrPWeqY0zCbs96nGB6mIwSNnXKENq7kTi/UqPwIj5Mn6JFPL0ZWjttRB+tumy
C385WqHqn47T1bRjfJlmBl2C6JOT/ccgXEMgujYz6s9K2Av7XLqlwf8cT1DQaN8R
f8nY0UpB/HM61tcwXSRAIk+p2ZOZriIpbHI3aMkMy6JIEa8iYRRwVzNFkhGuQkxX
lyE9vG1FxdSEzybYmdGrk4LA1LBHMqmPlcBsMVyT8EC7LxO8qT/nTWwdHIzTS9cF
3Jkp/2A/BhMiHQyk6t11oYXDJcHxGN9VcMxyGVgHcAAJf9MONOaXzpuskyW9H1+D
RGm5NylaT/Isc4dwm7qdRb+/wmGEN+8tUKR9Zmby42XTbdhwp1Y35TMReoLT6II8
aBmcCxQLlFruRp2QBRB8LlCqQL6SDQr9DNsbw+BDqkxqF4qmuDn5IqEoVJ9FBWKY
fuM3EJsU2qsznHyITyXneli0m2wtxIg6by0HpL5IY3NNQ8LHPQJAevJVLmYj3aJm
O8zUyIefcvzwKkOCY3EoRadFibKy/2Hfsgzq83X5eJuUfWzXIuZ6iXCQ4dVh9dLD
VsImg1RJPXAXaMI7ihWe0WXiJ/IRbgOCJm1OPR/BMdwyNksEUlP32b4LF7pKpkgM
yLpTr45gqiOsYxQ6N9Js0L8yWUNleLR4FF4NPq9bO5W3Gp6Rw8/rwOw8CAeiDNpY
Hiv2qlNIud7fIBjZQKvbsDSDnsMcn4GZBKqZeWI9zhJESOTn+TmSuHmAts6RB+uf
23ctBqIEKfy29ntJ1gObcKi3rFvyVUdR0qTpFfeGkX70A+5dPOsVBrY9XTu4WDE/
zN+Z4xTVoNbccdLBzFfd48lIW35nOV55PMqBLP3suLvKf+KANY75+P+oMsUfMkoA
hLZ0utTGqmJ/8+XSNJ/obFvpoUkLRes+KUOZnAoxtOcaj2q6I1IRZ+4M4jkyWrzY
CRLcDexDMLdmVOiDkjQen39pr7JKjLLpc5slqZzZmXgy+zv/GqIlhMvl9HHlV+JV
h2AD2FYLHNdLhf2Mblwd+PMHFdBgmQ/dJAYDnCkFdyCQxHxnUOGTVFG02FcAaWAF
jK9ic8EzOXgnfN5h63xbd0/U8z1CcLK6GOqP30IRYjMs53NoknQ96ifr4zKTw6M4
XTyta96np2KoSvnsT5QEWKOPvdvdRRs6vmyc1vPaGTZsCwE8M7xLR2+by2NSp0Ws
pUvy8/4IzuLN7cEiGwhMxuaSW4Np9pMK4tAGDcu9CjAoHvCmmTW6OF+konpZkR20
2njD9L4WJpdf2S7tskeGgE7oo/iKzJiQ0T3GLFPEIogAtWunI3qjQwSO4cKnzRDk
6DNexgcIgU0D0jnG+darhtHSolIqLK93oUaiFqSSkG5Ytbiv/q7yVjf8lN8bY/l2
lkPWrvyr+jZbJSIPxODeNTktJr1+R+ibc0eBbhFkTsCKQC7qk6Re3fIxIYgkGEaJ
6jjooqkJhSR+JCxWeiRU3u2rWo5SCInIkF6nHs/hRijhpTxym1GpExGGf2bpXTtF
kqZV2ZfxZIPBEDTJKrZdbs7gM8Gb6Z+C2FNJ+8skIxadqDr8gq+/UcOZrVtjrmH/
NdVHmIpXykjP+1m2EwVfsJ56oVH2Nb/9OlQsRXR3hOp3WubvBYH/m/cZkywf91BY
L1P4b4JYINQ0LFcLzVTbLYfVAcORRFzKsYauWwvX0iWNbSaCR4NFJWZUEDslIYbV
hQUjOgr6/f2VwVtCCZHoT0V3EwOiKRzg7e7cp2ZOquSAzU9vogb4WdAKJk5Rhlrl
+VflU2SLBlnj7RccZldmo1qKD/g9gop0M+LW+l7Kctvoo0I+Y3l714j0sgl5S1QX
6lYfhbDmoe8+HeoYCO2baRjOKY5x90vdwc0omgiDqasOuYzZaOUuhfkS0DxM1vyO
1VsI9vqNNYMbO8pARe/vrDGbJcmx0WUuSKJg7iC6FCEL1x70lq1+Wfk8/oYCUW98
qsvy1xvtVaIORKzO8rF5YP3a2AKWzcItx6G8Dyudq61TJrmKf3dEzZVId3VPlubv
z+10s8ghHTW5p2+5I/E4QvpbLF2cZuOealTo5SN25Yc/tJayei+uV+Cj62U0od9Z
qXM4Z9azEogxu69fpx308/R6p7dm3fynxdt5UdzniUn39bbH6BJJlZWD+5K+ytwE
LlhwQ8q91g7piAr5iSmZGa2CuZTM4TDpMsv2z4nATE1a/SB/05lfVNtU2o/OwNyr
dNs396RdWt7Wd+1non6HEfTv+oSLTj0/ysb+6HKfTXaWjG7zbPWcM+F6HnyVuDro
CUEq8m5VMpJ6RmZ3Rulvr0FwbcIPvxaPTT6RCpapsx6KSnogZIWk+C301m/B03yk
Py554tfLe0ICWp5sEAf8Yar8y0AiXASfQa9WNsBpYhWhWAOLla1A4pRtLrBPntfl
zsmYsTp8Bc02ujEOwKOTT3Xovjx2u/fvDXripOX0Pjv3jfk/meqEzusfbk3dob3E
neoVch+xbgWm0S6YujGuOB/xnEUraCZ2+wbW5aUzXDfO8hEmsi6CE3E4S+vCQb++
umPZoFD8VdFXioB7cJY2NsGAKB9SeRatGMdAA9X8gfRABXbdBLJfL1dU1Ye0UgUf
qPurypK96OfKbm0GFBElXfL4iSkForBn2opmssoyA1oPEea4bsiH9wcgDhHCJNHA
lC/D7EuxSM2FXbZlPUJqn2EBlz7GAk1eqg+hpkC3CYKh0GMa+NvJQkM28oQCCs/A
d1FvT23V+C7yJYlk9XxSdlErZgVKdeMB7iL2MriO6tdA/VSh8qeCYV5SEyZEl2cu
TDWhK2t/+Zt3S982C+S7FFdd9AxIWOVsRW6fQ2l1Ee/NPz/uKknaid5k2AZ701o9
HBwC2mC47lUDRjpLeNCPEIkUY1ejdDn7OcsGDmiy/0poufpSl1eEgoodH8+8or9I
M3AeKHG0sfSzrLktCDgTrWGttYKfoUR2HSzu/I4/vdAQQQeWMnmUq+jEMqNAOzWn
+EiKi9Mis64QP43+j6G3pieZXcbbQRZ77KRjK2xl2BvNX1a01CGGxsdE+ZH1Ievg
T6GcQJ6XZSrmgNzsZdiaQ+faI3w/FPkZ2oyWDRHyDflh9s9flvHuzOEXh+Dbj7Dv
nUH84Ypop6WXJTXJRhiD7CkZC/gfvd0GMpkSs8JQ+QI9KcJgsZjagJZ0/lyvQ9ej
84G41Y23U+WjLW9ecrAmmTvsN2qJDwXUUysv/zVwRRH8wbSzHsqoj8oovj35eGDz
fzpGYM7eSCXilPYke7RvWgepxKJ7VZZ2xAoHQl3rO5HXIE93O2yxQvuO6jpsBmJj
HRr5KUUNXMFa4dM+xpnE9aWgiM50HuVgIxw04zCJZkFvm3eBAG5RI/BKDJulOykY
p1th3s5f9oFV3W2VOs4RXZhLhH5TOGEX+hrOu06i93/JMpWQ10zcfa72zCclAw02
NwoXzE6CuW3Z/5MhR0J8s0W6sColRTxv/RyS4/snOVvyV4YyeHG+7HaBherYp4g3
o2FV/VvM7hVLEGMilrKQtLJe0RV9mUjF3LyUx/MCn1vSvZnSwYT5rVGtmOnnQwmT
JIkJZZhRAOjpQPVUkT5AAG2JrmEaQ1foTZ2a2A2UJSV6KnoE9m8ji0O+EBEn9vk1
XVt7CnCad19Cpiv43YKm7gwp9U8odU+vopHlpEG7Q2lUArwGGHP8v/iKhcYatKNL
NwlcoClQaswPJZlZ/ah17Wi2iXZgTBE5kNdljgnbT2i9UKoZDqqpvE9WZvkSyEJF
ED2thPd+4R10farLWD7NO2eTnOVcjH+YsDkQR2rezyqgAUa80O88fr8tmVFAvffT
bI3BUbFggtxeEcsljFqsaacm+FRFGemaZl0cMW7oi55JQOHevoFZTOy8wZKU90ah
HQxs0Baj8yDt+8MobPij4y5YjdN4T3GnyCF5V2OcTvNTWm6bQzD+xragAG1LbhO7
lEHcxi5OsbgyquzKhLiMYBjbPoLXU17e2aJFBtTAXIZ2y/lngIS6i1xwl3BxTM5G
VuP+47LxEtFNW7MxXWIcd0Ent5BHDnrMvwGGgC4DP0ZYj7Jh97Vh6C/y8f6Pr6wJ
kRnbUl4pNP699uFXlo5nAS1rqerhopuMx0DyIYoqJ54l9eX/p1ZpSK6rMCP3MEsL
yKPLZ1HWVSLLYY2NX2L/DeOCXXgRJ/TAT379ZyAMlIGxgwyexfBH6bWVjsf3tvTz
5jzjsIFTX3pw+VWHAYXhMuN3JrgitZ0lcmlIGzqIYm1/Nk2Witf8bbDgaG93zUhn
QQBJnuv1OPzp494jdmQTrwuKrR4TxpZSXh/jGCaI6JshBKviKJw47Zuin/9g7Jhl
M6trGS8MATkWoiclFlcwf+QOx/t/9MEt2tYWrKEMIJZZPosCYE1inkiGgOjgTBnC
uFhfNQtaUqxzeGvg7J94YMKd72c3pEl1PBDppA+K7UFYj6EXADhl8/9d6q7ohdWp
o4M1QbLGZlAFIAY3x05uOSRFCs7ATTfCWJBJfGEbnw3Vu75gm6KZCmRa4u1x5DUY
vAYt9ekmvciwnpDV5p1VhYJCMQKyExmTapFYuw80gzUC37VshrdXK5ouS/mOu1yh
7S/1Trvq/NUFwb7sRGNwmecnfqhiTnaxULBGaYCcYWIBJGsb6bmPC1iBEfQ/co7c
v5FgzhT6vlrxyvEdXhvlrLsS3en++QAxua1ohHQn7EBFe8LOwUmpdDdtOvWq0qrk
rs3q7yFU6WKfd8NGTfWRyDlggkyVMbxWCWLSecm6C+WcRd+w+la5UXHGQu5f3i5a
z/kbd3ygNS3PRWamDkqy47Ejg0E1HD7PICW6WhTN+0p1VAPF9iCFmo1fQKT/ZYEK
E+6GbJX4L6rQWfuawXHwWVZhNNFDNp63J1RPLMOSIU75/qWOrxDtfhSgVeA5Lr3v
CYNcCjv+rKLBC1L0Fbpj3xxls18+nvskvsbxiQ3TxQoW2q9lrlwUrul9MTmDyits
xlvd7cfV2fPt3bgujj/gm5STqR6zEcVd2gp14HQomv+phYtK+hmOh1NW8xu9w9Qs
t3ygVXl3kIgmY2o1py6LRpMfoxIaOQRNQTtA5eKidWoeYC+M42LIIZgBLm3PSBbh
Fq6/WCjPBoaoc4DF95uawLVcxLWtCywZWDThnKZKm3vHRddCL+yzLjShwXG+AduD
wJ8HO6mM9POii1jqYx0DXYSXFTFKvjNmvBrGy8ucCpWe9MYvgBXh2HiosZFHf4Kr
+JnrhjqKugfDBbYWRu20kPqwcXZr/7yO5nBSPMAAd2HwXd2PSHUSwDX8PLouQ0yz
VLjbniPBEvoRdGE4EYYzY3uRIhDEQlJ+O165LRdx7fuZm8Mu21AW/Fz33smZmpGK
REcPz3ODSr6xBebiVuWYLaXD3rLOGhmDm9m+PF6NTYzgvp9X8fxEs3HDnSS4qoWQ
0UsoHSMsjwAoEamCxPr1ym2jfjqEKmAQnTLrIxlMthMdzD8RFGgW5cpuT8ZPQDoe
R687keR871zlklSpWilI2gFbxO/Dfly32X9lHFc3QO5UehbA1kxDvaRmebpLIw9D
Q0E8qEp553WE8pA8e86a9ZHHg+y6G4lZK5nRHV6OULbQbCBg/uaXgx8Kaxy/AfDR
erRBvEQqyUts3TZodPIoEwtqjBa/0+uZGAvBldj8V3E2/Zde5bS6ReFsObNNzwjf
F0AJYIHk14JWzqotd3t2AP07Q8mfxEwGnOcnyhpO6ONz+NUmzk0D47YWARzUWnTB
bJMyEmqcFu4tYLt/WCAKWJj6aCKZmbpu/6f5o1+NK6itxyRCBlKm96yWhQfwf1nO
CciMjo0ft+P857qI4W31UIU3qyC7prgivEhr0fBrsyq5WCPmDUdubavmHEy5/czy
OlE5t4eGRZB/+fRvTWqnMTMGYdsZ9Oa6IX/fssXdFZjZe4eVyutRlAiNmY9bfWSz
YI3HVm7rPw506ZJc5tO/apaEkVCa2hh5a/CY3q+gLqkdV787uOxeR32hJm3Dj4sL
+/eSV24ICeMaG13Yv4aduPXbwn5Zud73UWc1yGUHxNs3E7303tYb4ivhbY7pmkb6
psPn+EY4DJeZ+beSQbWvr0+0KsGMKuqCC4VUjOqUmrJXyN240sZe+vJEneINhGkd
jehD5kH0bFhbuY7eBhLm5eVu0DMAfF45Z/4G4Kgg6XLLSQcRu3k7pX1+Ls+iF1YA
yDY5NgXgNJyCFCkiSKdkB/WxptG/R+Sgr5hpssHDjnrrwoRtkOwLeYY2R6mQLNKW
AKoqEhg4LdufovSdKTReWr9r5LtYvLLH+0KDCWlp35xojlflDlnTR1BJdhs/cNZS
0cxcWF9hagqGoBsZWsKbacJBpHWMXl6xxnxlY+mL9hgOKGzQtnwZwd/YDBrVK7Aj
ZAvNtkWSGiDRxfqXagC6ggECOJpvtqP8U5ezkthTdE+dVVhnmHtnCADEgMAESnyn
1/UINm6Yhvi4lq25yC+slr5ZKZtdoxkT7k0pEAckTKh4XoLD9gDieAEJO2aXISwr
V+uwl5H6hXoecorLc6wUzhr3AeR1Zx0OM989BwRhQmKezSW9hFjUry8oSUCU2Kpm
axdJI2cqWroFWEwX7IhaLnLhIODTjdi+5HIgk7eLIGsSs8mIMR6Hn7+UizPfAAnr
1wEwbyWdIRjpggneUfF6k/7aFcftwnwO9lJdk2g0vZY/iGP6aEZDSk9FJhRG0xCZ
A/Gg5Nf2FjVXqGVFF9PqcmJwvZC4W3ZZEvKb+4w94oMW3A03wP8i3jw9ewOrBHBy
DhjcpuHtBkMjwVINyHmz3Jgrk7TIg8C88DXbZaCyxHIiY0/psuWoi1FDIHLmU2C7
t1JfCLE8eQudBaHPcAIlJoRz/Q2xJYWq/ZQdEypVrphuEoEZ7SiLYV53JBRbouGh
FvSEig2UenaAbVCexViAdQK+EAvA7NcXnHomoVEkC1UMVG0pSqKlaInlCaFp1gyO
xeD2dsk8stoqdxE/914GNv/vcsHfkpJpliQMTXSY1iU2/aIW3P1zguYmotnMZYV3
t33xyLgByHWU4DCc0fm5vwp1dBrbTsPFzOD8iX8EVQnEmXG9+Dob2yHpOnkcY7cC
cn7GB/HTopRDRQG0eVLIsxsD1gMLGXb6P9U+/dw8V663lR3GGu1ZpRQPYozaEw3I
NWA8zdJOUpwuDT8DGFJiT5l24GcxsfnTRy8dUsub6D/ntszPnZRmTC3M7WrDDafX
K3eH+08Isxq6LlJzIJsXDuGqzWhCCgnNAd4xjpkhU3caNjFU/VAbtBjplOaHdtDy
SLpSFkHeFU5DWEBZ8khc+3Jqu77/hxTuOZbmKzN+dswVKHowd32fkoTaLSJx6XXr
3AJVHF6iCXAOqOfdbqnyu2WTFLrZekyHjccTT6THO9N4tjIhIL04OrHfg2WCrzPe
UFwrI+9kvW/WFzx89B8XfLsgRJuWf8qIUpRYzJeyy/LwMxjWPwJVjznaLyfQZEzu
Wj6efMepT9lF8M6qm8H5ONEVlDZgGPiKbKQxwucnKa100G0mpJ8uYtmQ7Pzxf2hk
bNqUptIqdKmP1dbj3PnOaMc904J8yGKqgpOocue+r8HcRzZmLQqAY8kSxkb4Am+2
oVs7xIIwfiwGRFlKAlVFYTLxJ9mW3Bfa5Vji+MjMO7DVr6qaMEvxDv7sQXA+/8eA
9Ron/AhhwJzY0GT6Ec56BIZUPTn+7RbUaKXExBR6rSGOvbLwutoXH4n9CgvMm0xn
6LnjTCBrEllOlgQ7h6nkrkfju1Vc/hng2f3uE5eehc17E9turzkiAlqwtmhuoyUY
8hcCUVBd+oBSvsXxeqrvcPAKLoIUuz9+LpifzPVInEW5Eb2WKOoHW5WEuQg7II0+
2AKmHarjdmeLqHBiGC6sWzLLPKmHJuzwv5k6l9akGWSXzgEx5F7MgvnfXNU5S9sW
6kMaY7/1R1CrqEmabl6uLQjJ/pNjrBe10NaEqRyStu/LgGNRVnJh52J82nLWTq+C
zkz+Oft20V2R4mCFFP8tjkuUDEk6p5VKtXETaEEOp4HxYYBn1wPpPxiEPrjbHYSN
FbwNyBBoFl55C8fKI/fua8WV+SmekflSawuIuWFoSy4WeQAjTRd1lzILE/ZhPnk+
9BlfY3Z5IN7Hwicvy1xB/S5kg3GrInahZWJ1uTOEyZFOspFiJjBS7rORnQQM1eH2
mv2/KStPy38YcBq/VfzzNI2PfOP0XoA89KOBtI7UON0YlLnlMxsJfzyAHHXngqGn
302p1MekBND6QXvtMKECWxcjyW8eeynUBAnDz7p7TjKVPcpT+d0p3MjDX9hy8ZW5
dbmibL2VWa65UwPBB9calrUdJfLfpEaUl4YvpcfMC8ZZkrYQlCDnWzfkqENQavJ6
6mMwFDQbvaH4cbUt6L+F+tgkDQYpezo9thrK1VFFoU3aZqCNZD05QxzmsIA5nI8j
NL+T8d2wJVkfqnShiqAVfEeqT/Cj84Gok9eNDuIi/U4AzejxIRzybeMJIkhF0iB1
lWPLPFw3Abqkbxuty+g/07esZUSygbo8QcY6Ml6EvfzQlXmIaaQiNwr4c/GcavCY
wD+jQjBHgj/f6mZZd/JTgj2L/oDjwfXaOIisPl7pOMOfaM/fjO1PhcGoVireKpL7
OsqVqpKqu9tB7Sq9D/SGTt6lMjZAqG48GxW9aRAWs3/AwNJ/k86hKPUjtaivzdjT
yOBJ/KB+HoaORMnjpK0QiQshzX9VUmUhu+q0ABdszoSBZySHmghauhrpilfAyJ5K
0uQbNS4EHl3ZI1/YZ2ZWMgrObTB63qfVBlXGibsLMvVDMcs9g9LQENT6gEf3Pdlv
6QZenarIWvJ9hpsH5rSDCNWjhZWaocB0pntlHGye4rwZfLTymFMNn9z741qUL/at
U+xWLKKUAuqs9KCrFZvrvF7iOj0ikRWU0kR8JTIxybr/48cH5q2B9fYmz0kwHhLa
+ineCncmzMAaeefjBSqIMsoffe9jJJGiAjqwxwF1uMW2z6uNBGJzBnLGLRg+JWtC
VJXr0/k1KWSxURbf6Ri+moSYHa9s3DaemwL61DI1N3xGatZkNSgeaEJVgiUflTCs
P6CoxjO5gzSpaLvb4FUl9HlhfYsluxHf7EttRyHabNHk2pIU+04RCEDEYVr4ip9u
3N5NSgZLRCYtDewUoBhU91hkDO7AvL6sGxyP2aTYas20ngcQLm9NzO8oXRpf/GYG
RJg5bRW8fL16nCqXAE2+V8WnSUf0c06EFoFiuRXuGqqdzVb0i8tfUv1x9jcro8r0
/G7OxXHYLvm0T+z1R86XnFkOxanNz4W87GVdFuaoRXFqFlkUjUEwZkKRzGaj37tP
ZTK4n3zg4oJ5dxLbhS7cf5Fh0aqWmFiKKaEXQxXejZe9SlYItiSFVVFizxmjDjNJ
7lrZkvm6diFT3u6UEZj4Ch+B3Y6g6jr/iT42JqFY9So5V7lO3strZqB2R0kaWOCy
noHAUe6PGACKv7mBgNdgq0qJaIEZDX7kcAe+20GMxlKpel9H9cUpv09VPysgkznY
eV17ffhtxu4cQt5P3BfqgBtuSEbxsm//loUVuanigOBaXnX1V2IEzjeB/OtNHuiW
G8ftNwRDYcKgV3ppZO8ztGnWGUPUeYNafwQ6+RnVQyfXbkd3LP3D5mnk0Fo19Bi0
dvuaWZfuPkhTevch7EslISMVkdD2nMKDONNkPIL4zlCOBdqS+V68pra7EdN/Fhnq
+Bu7x1XAF9r8j5DDk0OSP0ILmDOPzjX+DYGmEMaOYEidCALV0uTVPpDXbRayIOsi
d910oHCDqOxGn1wEsSLnOQMBS54C0C5DqAK/FNxJsxJCgGc+oKyVIfwvNy0YJyj4
TmMuQlmQhCB0+XHl0Yawo9W5wyyAL/b39cuUmXaCv7U8Qkg6dc2RIKU62A3AS6L1
xvEnNTCfgYpfvAzQbeYryQSwi2tvPl1cW2DvEvE0yAK1SBrosl4OcArY2RtV70/I
y4C4/R2HexJobjweTscQ3WJASti/uBw2O/Z8mveKVLuhZyXHmrpOTBRmX4IyNNso
Ks59Qvzz3XXiHRGEDAopVWB/QAMYpogtRztOBUtrj+h+bD83g/eTCxoh5XcyzW6Y
TzVsl/0qE+G39gRFmQJs8J0wJhA8tDg2ZSC3gfQ+rDEySbarU9QqF+0K8l5gCtOH
ie9Li/6WgP15crurtJVPmp4LoXixKNN+PRIzVmtSfD7fjtCgIsO9E2RsIwd1esrt
QCLat9vOZ22N29Xbgq1uHvxVCeFt6o4TZG4nHtlioh3hD6e2kFJJyAsSEVT7x1n8
+XSiW/RxoNiDAhaAvCEjHHTVMJwwM7InQZFy9ZCg26taqzGhCnWMPyb+nQngg+Av
lQ6sz9ABXk74/95nf2ZOUka2BDPdpo4pgIvt3/X2ESFbrzzmiJLNxWrZ2hw5SToT
vEINgCYIYqT/bnx2iGEaVyKXhUKHC7D6ruKHNtXCil4OTxejkkvgCEjXw40/UDjA
eoB8NKyM6RifHF/nx16+yK27vJzJtLi/KQNgbA8rNLixMdeZEZYlQJOd8YC80mnS
3k8PILVnckja++tbGOBOxurOKxo1sG1O3+3FS9HW+qg/kS5FY32ixfam1Imneud1
IT3rQ7rGYdhebD/Lae5hRF7HC6vOXPSL538JuddyQ4q9EXcV1Z/DgaInh5+rq7gI
+ibabZI0GPtSWeDMNBwdCMAH1bROQr1bRkbIMUPajtBucOXJbQDdYknlASQabOPp
ASKYnb54clkg+Ql+nQjrEohDrkyMEVzQaZl/KofgeMUHs+Hrvpuj4G2SY12MJB41
XkN7f+9ZwUUt/5ADA9ejtooiLH7EZ8MPXlVghz7HTeBFmJsJO4annmzlzjmapE5/
yg+P5HfbJGt3QvNlzzbJap3pAhKDePYTakX5e//lCNgtRelIkDNJypRj17oWaJJM
X+Sd3PnY6739f/dion/uvlVDtQKfEDOf4aAPTPfWJxeOd7kh9Vozl0Htfhplk65W
WRZPv7frYbC1j60pAfAI7N+I7dytV40RwP0BfG/g1TRqx/stkpjk9cdsP5cFnAL7
qYCS9x0Mhi7xH1LdUeO4ES3VED4Q2gFC6bi9Vp+/GkawhLDtZYi9yIBs60ukcPzs
5GTuOSH5jc+HGD3Vzoil6JD8DQUTwFIynhQBiWXJNM5f03c9vJWGws+qTwLqsay3
gfr666o57oLZjXlQGwcAZ45cDSs5buOVysE/GGCDH4nEBra4whferXvZOjQKF8Tk
JhYQ9/jvCaMCzdd9iy8MD42oCw9DegilhuNvtMvmiJJgS/qW40GEq3w32XcBAONk
WQiFtqkFmaJTfr2XbnfIw/mpphKLDT4Rt8xvAvR9ImO6o9q/L2aSRLuR3Ke9eZBS
4KxXw849qPBBAJZMV9gJ4ZS/n1q/1pbwgund74fBfLiWLx3JV6lyxqD4PqCAYyDO
3WTtbdhp6L5fG57nHMZLIkjNZITvqXVpzCOAOXLueOdnvYy5NxRdS2go4uWTJYYO
r/dFV0DFDUl+mDpGhu1RQUhjB8dtOe4hgq8NbeRfU7wpnGFK+AdM6wh9phuZ2ull
IcCBl4Vihu+fjJbfNZzZ61z9cRC7fhGMvXc89k1uJXNfGf1JwEnFVQBLH6yvu2LB
GUYm6syZxzG/lPLvsIuaS4pWwkM0VtrfH7wUnq7DKQhFJrQ4Fstb6imLzZrWn9ZB
MxAEUEowsVGCAWahWVPayFSq71ZUz7oIWOOuvu2tsGhtBpTtFPTxGIRrf9GYn3cd
WGWW9FW8aSL7MfuDylDTGhAa+gp98Y2+BjLledIpg8nwFluBiBU+LEpsIzp1RBlI
K1KMLE/aq2rQjBgWmQ5oT8qpGIGXpgvlmoZKaTsBfeK+vWjWrVDUixDfbylFVG8/
GoONaZTLjL2BRnGdPH6xy33D3Q+dPAlaMGgbaJCEVVIQJDkLG0uTu+54/uKPHRQW
+QE/zPdo+HiHzkaq/OXPGAqJs4hCgcZ2bvduoBjbr1b9MI08AzqMKJP0VLowiTIi
EcYtyzSWYwo8oghz5qBzs4FDUkd2zHHa6oIl/P21TfSDPQMqGwqVyDwSW3pjjbk4
1+Xglbff80bvrD9WkGIpHSpJ8ZkBu0QY36OP1VjozlI/Hhn1BQyrTmO16Kzfj92d
M7qo/Q2S9334JQDEUakw5fbNcGQzT9U94yUcN6z/TwYa+MMP5hcYYTDtMjOzCuZJ
oNvUrwQZ3BL0JLm7DCZ4yayqkZG/U/oAZV3shIeLKofMw2skEdm/AzadzaLgH0sI
brTj89DDrbqst625QCip5jgNmJFt/5opM11fbZkYmI0sBEKN13wuiuaotEtLm3Ld
WFr2C9nFF4UhVwjsFcrhnXiWGULNFzFkGVato7cOAAfvIi8uDF1OCoDI+R+1Fg/o
oTFZcYP7J58ftxme9JwNKwrDj1m3kAd58/IHqVbT4tCa23IM7fNuKis7ZJlbK4bn
ldCICEPujIOQqg5cX+4VPG0BWPanGcqswIG+eG7jvSnq8lrIXPNUj07pSxLOAREQ
ASsP9OgdUb7tM5VF8kwZU9T6+GZZaWf6WuaZT1ZiyBDBuZRXVV6sn7JttOCNZ1Po
y0dH3UBX16At1d93Wl5iPN0/4tmD4A9UcEAHzcjri8h8o9fPLztZRwsrv6rOYGRC
iMwhMVOANi8Sz+CJ7y50bpPQUtB5IrMpr+74VlaaMEuBxDY082KTSGTWGtnz1eBc
o741qpvd9PRNDicTzs0ILwk1xVwEKl7kfJz8M4y/I7mwaDMnG6lYDcjnm1ofYzju
jajBYMu4/ghcd8TJP1s+j1L6ERHcV2fUweiOWEicdB5eGRGPjaMBm9/6E1So1gAI
6xhefi7AaS0Add1nkTPq6CPwsplmmtORKnV1TP9vdoy+QtztqcOT31W7GzBP4hw2
0A2euFlHwlyJezwzQAOS5teJb3gH8DHyborikvlwPprC9WLyeLAEE8cuMGqri2jO
ZEE8Uxl9B6V/GPSs6zZM9bWjOkTWYFm6YiF0He3ss/I9ull3teH0YopRUhFbSXRx
YiRQuAY8xl0IjBjzIRP4rJ/Cn4ClKXTc1kvbuGCOZXpA2+PA9tzkh6RQbrl7+GKL
aWdiAwTv0BaDlXFvhtThKoJY6Oan/7KS/IXUrV+/fvJBVXCVhUtNk2yeNvr9U8Uo
9NMxmm2puJan98tPRb8byHPyTIEnqr01p7kX+gHTDkmn21Y05Q/8g1A4WGW6g5+V
kiejrVaorMJbiwT8xRmRUIMKhODWZvWbkT28MjeaFdKQ68EsuGsE7As2XlYUZwHb
vkO25Htgkhf0Yn3yfWbs0zjp+DWUFeaNC0xSARqSP6MMgVGJOidSp6kn8QfE8XzW
tQe3+UOXnTH41kRIKXi54EHhmRdIa5tQUBYdbBzrbeDOP/CJmyw/9EFw6vy5ah8S
xAdD+/uTKyQ9hW8EuVq4Nx30zkJ9DPv/5GNUXzvLCQdhXwgBdJjt4UiU+GMc6665
C5WgOSdklResGwH/SyO8vKK7gy5r4Mf9WZWLToy7TZ6A4UMh2ky/M4rHK8PL1acZ
LyntjCJpDugAJ9a4r41jxzYv6Blqe0S0S5lIpqWqifR/Wgi8QKa+Df9V0qGVhaIu
1pYtF+LjZNua1DR9QYRsjSjV6Gc0XRaHaaHaFGdnmVk8feNDIeRED6lMFSQ2wpDo
kQE4YqcuY/z/+CbfWNkvhUKmojYJDetiMg2pz7SUw5KfU7CyoYzYgZpe/sQC3rO/
/9l6oT3j3sA1AK9bPT9EPHM9RMgyeT8/I+YYMnrumZLJuRVjqhHgP23B8NvbFSHQ
ebxD0fQH90hkXXVlD3+7NnvTYfqfuKkCep3WMjHeZHqCXCWscVdRtLmAktaor/0X
Q3Z8h9T7J1Q8OrxltwhCaFIPpkB2mPpNR2ZbMnoeqZ3itvF9KmCdM/TezJlRONsB
JZdY18xUWsbuYXKeasHVXrHPAYcPciOeaJSDafkv9PuN9G0yR1BkgdR6Pp2rm07s
gVNU64IWRy5oXMjCBm4llGXZy4pnE77wK2skl+Cvr4ktGsBx1qegLAGNX39lTzXh
paxg+UvASN6xe9VC/EUmW897jjbNy8yToPt9uqy38YX8xfBgBWDq91dU8ZJ55wWo
Xnck/wjPilJj2vgOcv7C4RBvluvBMtkUkgzjAbS+N2MPyhzBTIZIsdR0GK7EtV3L
g77aDA2c1iH8YJ8qzBxBmkKZsK6bPSBgKjvwemSqYCSJx84XAGptzNbLYKY85AEd
9ZeDDpo4DmrUitmh78cbTqrqYapHWBiF4s46+Ixnx896FmHKEEJIJ/yy05Sgxfmv
jJHCwhG0WZ7K6mOku0nkUlDR5G+w9FX4N/UMkzh7kzE6WRRz+a+DREDIEo/w9hpW
UBEP0TP46Z9cu2x02MdeU8oaWTrByB1WhKyWRTGn4tQkRvQ543+S7XWSAEB02c41
nr26DyPtlhIcBjD23z1455T0WuLuZawnXKiIAcr0bEWkk0s62HB9wyUWHe38mGmV
lYNRL+dqsiEGYe/oqKX/Ai3QVObayoLu48d/DkkbV7YHX6WnCO/tya9nEuDL0dRc
SQsh9zjq/8uV2mvFSwQoIP7jetLIKoEby4ShQHFPHkUgrSpsXYmo7u5qDF6+5h5F
ct1+HFZmqPbn/4b5XjteL/MsAdov8IfbMJv8REH0Ui+lC7YbHDXH9xDz9zEEL5Fw
o7ZW03HAbwGAcrJLa0o7gji55w47Mrsj4epZE01y8kc9gKBntj886keG/QuNHz4y
BtcmWFsYJxK4j+y/qdP/5X/PaK0oS6Ob+IzhtnY9ldq8I3cs3Zqnb6YqA3JZUbQw
DDxRmq/37BiXcEGlhjlY/9dj1F48+Y4nd3hqKPLV0UldOPe4oI4/LFd9lQzjnCL1
x9uKvoMEvzgSB5SAyodzZPS06/QrghfvfVccfb3riaxcRF/S8xJ4mGZKEklhSIOH
1ypdBwFoZ2igcUSXw9fts46RYLv1ekOeodMV2uLv6819oARqg6q2bW3f1UwULgf3
xJo6nL5xJ7YhqGM3t6kmY074ebLowZESfZ7pGcE9kElIVhmPUX5nesrFn65uR/5u
ybN7y9h2n4PulOjyjXGABVITWnAc6Cy3ztLLczNdwLY2eNwfV7/WdMIRRkCYbeur
ojh71aHDBIKf01eNDD57Y32JrxxvPSAey+aKAsLnoJLZaS0ZT6YO+JtKcJMbj0ya
CmJWPYqXSBpPtvFaMyr7Nj46Mcp5oqc3u3loEtG8+10gR9KkXIeFrM2xjSsWNy9o
2Se+0HICbrkQAqXrkEwlcHpvem/2J8rkE2jN7cAQMMAy9OPGDRUdrxlmONKDoDd4
3VyNeTuexGhwJfORwd+Y6aECbCK1pmFdU/LnN9F0DcQrrNkaCYCPCNyRkxdN3rvN
lzIN1QHS1WwN6m8vLBoZvuAgiUHDH4RpO++9sanGYf+ID2YjV1Xg98QQWsDAqnq1
eYfqLmq3jslGriW/3Tgm7720qYCWUVb86dg8TfNSWeP3LwiSwDB2Nzit/toJkHCF
y4Ft8pf7ZC3AGZLXLckkCNyFkZ+leoPWQBLn3UbViI6i5MSponzpH9dinmbRCOKM
htyVheFegv76Nj0+tA+lclaHK7BzKcqHHBq1/KeTE5fNryPSqhPf1mhOsarpUeEf
1DE7FfYMhO07MahX4j3Z78Mcdqutb+p8jFVmVl1DrHN6me6KJdZCq6Ee9R6/qO3X
HeJdIIJ6nxT/uxVg59px8EtQoa7ivBCFteG+GzXkmGHWRBloNquMYw2/CSts1kwq
MBH6ag5/dE0LjFztAQJ5UGuKsG0EEauhodOg1P8SB6sDtePKlAWcYe6JdM+Hl5kQ
LrvTwprrtcRwVBG21XbWkW4WefF2zh/tRMvFA/8eR3qvDJkWloyuc8YQ/nQZtzaC
FLy0ltf22acluQiyzjKd65J3074gvpE1GCTopPrPxWcMvZ6N9ZGHHMNv7FAqpcPX
aqqel+byabT07Z4zBaU5796wC+QU5u7eCSOm/XUGt+2MGO4hGbGVRpp5wSyyZMKe
XQvgz0oP5CMVzFOISzKVD3xWS+LxhxOOwAd/78I2eqWoByT5h/6DRu/orLnBBBiE
MIWHpunr1gGBayfDumg978FsPKf0tQG57+6Za2xE0qAYFUWWVKiVNtL1yT6L/zJo
EwU4zsPGrUmmf/Kx4ez7dtjgxTYnw90mr/5o/v+UWQbyYX0s5YsZmxjE48VX7JEZ
g7WgxGt3MvnA85QcBNkXgMYyx2jlwx8r4PAeWobIGt7pKDzUyB08MkQqH9CSyMVt
GfFjJXDIJAThumcSLKQEItFHQAM431UAGpwW3A6Y9OvwXyC/I6kDInWUQ5SGHqfZ
yfUTYM2ZcgCXJ7r8r6haXkOrWROhY4aA6z/E4NVZSHUCN0um9GN+JbJ9MbkEsS+K
0uz909ulnFXhIorfBfM4QoxS4nSTEoxpATuXARdp9/e4PIEf8i0QYVypPj/1mYZt
UpqdzLFFDCkmoh6AZ3E6l9Wa/jK/lBvi+96i6HXPTbkOwXgtXtYv5GiGIkO5aLDR
Eq0gPach0NqZTnH0KsYtPdYqroHihACJz90+Mg6xxxSE0P9rnXF54GCSveFXRolz
idKKCYwxpKq5MsBW4JWb4Q2SEyNP8xnxiQ/Rp67+gW0TQ+oZBrc/73W69E4Nfa2h
L1zPZOWJYDDlgsV9+3nbOv16UxsA1k6TX0JGFcy4NStb9awKkQPqCp3q6USmIbc8
AyFGnRqisITE4fnTWjEJqDbry3e8TBYOtOOZJ2lhHuY1Ezs32FhqV4GJwXa/WHMw
bL00LNQnq4zf9Ak2voDGaBeXT4uTpe7q6+KorzDTsm93ixzntsU+tDDSZs/kPsRW
Lf/ZAd1J/zuFHh+z2kxxdn1uxkkPnBvTt24TIHttO0Ps+NT0p8v9pkJbm/FwGO/0
wFuzJQYj3lA42nvdMmGboxMxLtTuc+ddvAYZ+praY/HZQDJv7bqSs7EDIXKV3dFH
1PCc3cb9KAdD8Byh+adVbUVYAaLZlPmQ/yyJcK6MqkBsXmQRru8oh+5OHD/pDJSF
IG7P25hnsw324pA2No+l70SPVpWFXtehlUPE6jUI5+E3o275462b+r9pOhT/N+rD
ik4DaQBVp3ZL3aj6SUiftPfJKLHP4KMFJbAiJcmesSP1IAPCDx9rjqUcUX25QPvc
5Ho7XKvOgJN+kzcHp7ekL0nuCmyNdxQAQ7Z1m4oAyUvTWEvOY5uqDPUQg45FZdJX
4SCX3zB0la+u3p85ik3ibj3lANph2Xkv9/GrXxa63ibJQ4ENlVeGj2OPLDfeEZSv
fTT1jJ17pe1S3rHAPxcpULx0AHKMRJxsZQ4M6vjMzvZu0C9uBEtqLB1sUTgv6CJE
1xYgNZ6gQEph5fcIqWIIKJZN5afj3oaoqz0uw2XUCeuP3LqyD9xot3SX+JFBipmb
TOSDpa6Yar9mxDDxfokjatORXhD9dVLEtL0Og8Asx7CyaLCPv9du3Utw2NAyh1NB
vWMeYb7yYLhdIT0TJlNWKZ4Lgbt+7xG5HmzcaW4wk+vT7AVNzpewPPmqF3ev78b6
PpZDOd+XOfAzfVGC40+grcuA2d0vANJ0Op+hZK0cWK5LKUrJdxt86EqissAm+nR7
otUNpTn5m5PFmuDfeffzBcWI8edVgvbXc7u/QgUpXfRjWJaMKSWPp4d9LAnztM9j
qiJNm/tciQoeMOV/60P37tQuqYerqEQCgrqmilH8ehOnmQd9onQBD61/uz4ciOOh
VgBEt3mlYub1BwTbmGa66CGVB/Zm6GK6MXt3//8j3BYYn3JDesaEBKHtpTj0X4MU
bClhNcZGwX/r2CrtVTh68WZE112deriqpBRHHLsFbcOqXXLy79w9A6GChuMIMtTN
ZDOQffj20sLgto2h+VVMIKLdxz44LvGfRY37yR+NKY2idHZ/j+riPzYsjfGIKJ37
ZU4c+komrPo23Ka+d+V2zAVeukplCui1Cv20oJHFPI8Qam++w4aSbqfZPA5+fzPh
AVpgIcRFZq0JVmI9XpeF/UX2KvWDk99/69ssY6eDPlbrWvUL61NPgLSQZz7+ZNWb
dUiertpRfjbCMmFo8/ekjKnLzuRHaEoC4W4a2kjozbI=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
d4KHFJuH6MLLFAslIPnEMW6u02aZo757w0Hzmgr+qDE/iE2+ueyEBFSBhGS+zumL
yiOzJPrXaHguUKQNcVCphDeQ8fRWPgk/UU0VViGPSsa2EeTFHfefVVJym2QjHPKr
hmeDyxcxM2hHBHjyWlkg7vDXy3sUJNZNvE9CFENlLL+KEaN6TgOGlGyxgwK6U3sy
u5sOBHWTCcjTAIUuDUJKHu4g5TrqpsyXdm56k3iggtrbgV954knSL1mullowQqAC
cMaWuxv7xJm66K60Oz2fjemc/8pan5yz8LLCL5mwgCBPcSQ5FzlFwJdZMO5Oe+AY
R8nwEkRnv+7oNiwTuOnmWw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7632 )
`pragma protect data_block
pSJG6dFg7sS1rqOcPMY9HQK8TZNnmDWcTXdNveAMONWQVPBbZJc/XaXI+SkPufqZ
0hxXiuMRGPADwCl+AIz+GT7fCtH9atG/eXHHxg/UKjbMe5vkYiXK8Ylzs5RgOU/W
xZ6PTE/1pAEXj14sIt8fiByQVoruGRfgI5NE+7I/a4mxRYRbqlw1QYt1fVI+QkTu
TYIcKCrVttrPOb4zKyGUG5+cgHCJxFm9DzkRwuEcM7NZN6xGsDe7w5Hs6MwyA6Un
A5yanjbIqTHDwjM+up35zP5hLz9q32qozogibL/NRysa6k5sl36vXp5KXFoKrEtQ
cpHwOPPjuAxZ7WRnl5C2JLntulPHMfRwZdV6ZTXk9Rvh3URbmX0Ro2AE60xUU1L2
WLpIetjp87CSl0T8sHbZIbIhRjAfsHEOHGfbCQuwAWgUKGCpcw38I4xIN2nhAoMi
7MA8AlaABeNttQyd9fSIPSH8sRikxfwJgfz6nmlAJ1r2chU+rL6Wlw0QnKUMk8CJ
rm0UPFUdBjXbRKSg7rKswlpRoyHMSJT2qtXqtfIzuEHgur+9vfrP0jtpN2bKHeyk
XRKyy5sL2bCnE5DZtiyz6DK3XAF+ZpJ/gDr5Li0IwRVTc/Q6coGGMFuBTf16F6og
abycoAGwLW8W3IvDp4yGM/L7N7ON80/boENSNjL8dnnogbaxGP3/Hsk9c6V5YqWP
duOz1Az04KmIa0foIafXy+zKKR/Apal7JbxnQNM/0pn/mOsWM+vRtl4ZNDYyeEX9
Ve4LmXkfO+Fc/pBNK29kdOtI4Prjvf9M2tRLl//SA+Vq5g0do6cS9lrumCeiFrHS
OE1amrhMFZLgPUn474TD+H3iQEx0sdQiwFOB2US/gK3vPw2TCftaYq+HvGMkT2UX
piUvi8nImHS56J6dtEQQUZFYh6qLENyJ1s7y+dY2WGUT916UzVBo2SkpGi2IanvF
PW/D5MHbYvT+Tz2Fe4qsL9sreFwSSmd02Pt8MEf+qPk11akJuEWLd6EXBPPp6PDZ
8ICVJPx4n+4HwxI1hk+kjZeDUMSedFl10GUCpCcEZlX4obp+y2RZbM0J+oB3TlTw
1raILmqiX1NDKZbHs+iTGXiNqk+5Fsy4531LuaOX0i9Y+zJm1R3c20JQoSD3q8sJ
PfuZvclx9QNN+NDJgtrY6gsRI9kBG4itfGwnzuBE1NAI+OepQhq1XXERhf7FGGid
jK2QfaLd2VAI3CCtxBSYnRmwjGgaY1AZClo4XMIUaghDzet+CmQfp9FlAtg/4vEH
cvn1TaQd39e3+KQhbg0siQu80pZuh6XjIgxZqBi41c02cQ8e7PdLKxvpx3JiMlBL
NdwdVUBosWG/ZoeEdlI0+2X/Iaspbt3IP6FDmwTTzwijUm5NTgS0vIU8hrIErwyA
ABhjDjhewZlmDcwPjKVR4T+FRbD3kfdRe+NxKVY9L0pD3ZPP+/99sL85CGeLB2j5
82TJ5/G8csvNtul381oejOOfWWr64EX1tBoogaV4jX93HoM1F6WkIbBBUWd+X3i8
ubq2q7xSBmIq4kBX1I4EZaOKP+uQYSQur0ssHDsUnFaXAegdCpr5Hfo5YKCUQLiB
NaJh1fAHGF2RUDNFABLrOEGY+3NlP/LU9mhkSabtgKO27f0aZUysLVmCI4ftDHKK
BpSRKqzOwShFdyPRnBcYvAxQy2e+gIRbFxusA5mcy9kwS6ktuyNOkgCZJlvVbO+E
+cslkgFjlfGf4sIxY6eCYKd9ymA/SnG/qRnpLI5v0aOBwlSkEhm3R40CDVBEzu1a
O/2gAM8yMrYO23WMbKenw8cLtp2V1qC3zj2XBeP38Jri6h499W0MakAaOiqRPvtX
Diw67n2aYjaH5+88m7Nl6Gig7/suTo0GTxi16wHdOb4z1CtDQwfm/dVswLd5dDqK
dW68wnCOdcgTM2hi7dc1QDNAEXG3JzeInDGpikwYvL62kBwd7efopfBBI28sTa0a
wIFTnhmQaApgPsWVmAO0SnOETK0BprBZCw4BNnRIKlrpCcieZUmn9I1QBDCQ9jUJ
5MZmFqqbB/NzBSL6HJtfiirYFaR4E2Z6/c5bWR3Ne7AZ+sU6zFNfTT0poodidyDK
daMQHyrzeLGS36fBucrsO36UdMyGRBNADpeQ716AKixm7XBkdJRLbnygmO/X76gU
vk8umltQ4o4L/iQdhTVoWIejLh5Ca/tIOxZG3Gky8x/b5K0VvO66erENTo+fDcl8
LeGjBhqGFzXwcs6249gH1ro3OogtyGlmU5Y4OLnmnaKr9m9ID4atJwQ8HOAI/S76
wSKiIEx2p1l7hR2GjVBl+k/K2nz+XzTAnjYyJLKw6ZuzbMObMQs/lTefdd0D28a2
By1wpW47hjEU0Bv8Kj9AoYucMSyOWrkMUuwV4jlzz+LPDreXR/UtuhdAv6HPhgxj
LV9O78o3EzFAqFTJRuJN13ZdLNfYRZa220Nwm27sDxN665hJ3fsfH9Eo2Q2lsBrx
4F7TuI8UXfhXfodxlPDraOA8tgcaRZ47DcYEkX0WWVEfws6DpFyUdzxgx8uy8yiq
ItZtBIIUlTxxqIlyVVgeA2w9aFHR9yAGoS/DFxhWJxiYJMNK0b2A/HEtMuK1ntOO
5I1dcaQHc2ZLgkuf4dB7BIfUeHRyFFsw8otUUmYpR8ox+cz/Gkbcp0hioQNTBIQe
aMIIMDXRwMTNXlTVTDkBVPGGX6t6sRY4pkdA+cF6WbvfkoFnxVdUWHP+zaW8DT3B
uuXkxsLeWcnpICx3SibNQtP00QogkkhfsDPsqpGoMHTDyMUACOrgoiYBqMLvTIUy
mvK+HO8kgT8cZOxeXAfoBOfkmS3Vrp90NFoTqnTaNCa9WaPPWLhOAiwherFMhUgj
fRcld2XS7butawMCFedCxOeSUh5MAgiDtS7OU0Ctp7gFqsnivPzbqsUWMGT79sNz
wdm2BmCHf1TlTsCusC6o6P8b1jlJvign8KrfLw4pE9fwWZ1WdNZgEr7OFDaQLIoL
x1VVJppeNhUYB5mIku3nP6AuOuVK7QGI5h5Brm8UNlWEik8z3HdN7SfF9tc/OJaC
GyrSTVqaegB2b44Q/7LVbBPynq/cf7lyXGS/qAw5+75hNRo2j9+5gHFqxzKTnpzO
DUURtSApBElORj619im23XLwk9uSH8xFyK07kmCnj6+crN4Co8b0tk5WIjoqnOGw
Pr4kZK/PotCy2G3Y+WIYe7BwvCTWFBltjD1q0WnHP0nY7mdj6Ut38NrXSFeairKU
HNP/E7+H0ILVNLgfKlSm7S4ZUK1ZPLtiDAQJxIMLIUQOFYEGuVCIOe4G94eW6IN4
k4wrcPZXASK1HXjOez6y8JaOfmksQDEY5SW5vgkAZNJSGRmOK/0dqOy7/i2wM2hR
QwfOZEG/KuCEl/nV63fjzTvesTofhWRYTrZ3a98kyb0noTuRYapWcuwrJPYelJHS
JsHW2mFyzOl3QxzKiCHs+J15BeXFtxNQ6qsoNyHpGgOxdwWPA0hRs+sQloxdnB3R
gNqPj/lmp51KUwrueQGZuefac29uEYaDm2y7ir0xqY1pALxsoowpIalMMIcGkn6y
AEx8FW8m805oQ6bymFWiSVfR8OC4Ahxk3F4yrmjm0CBkhdyKjhvwHxn1MlJn2LtS
C8YVRhVarLKIN81aLNJyvOIhCDJKMHCFUGegOTT02w+8mZq7Id6lsueW/3D94GSs
ByeLTfEbHy2lim+E/qPlyS3jztrEeCTEupMVlzH7g08Fb1ApqXzWBJkgxVeTkJah
EBrR4yF7obXrTq9TDNE1Y5Ljy7EpH02lrpDSG8wFib0jAlAYm1YwVBCDSvhf76XA
4oyZYwOfrQh+YmZsPf1H4Y2QB1eBQFHeG+sQWA+kOOrB+IcrTbonhjdHAFhEHNew
k6bwFHefrh5E8V5fvFhLvRDysNfs9Ls+lQ4Q60UzUS3Q7fprjaPMUR7miHos0zJi
EJRA7z0ToVV+kJ5jRddKomT7i5GrmW8tey3OMaA4BZ9UL+sd2gn1AR7Jb2iD3duW
heA6Njc9UEeACEss32zBMalkSoYzhBQo5Vu19LSOVVmttU7OeGqxMA/vLYxUvEfu
BJe70k6z3dEzBg53ats0zJW68RsT1okYRgWBP8/v4IDIFgobnkn3bliu3C6zywSo
53CP2dEUoTwVpzm3CNg6c8q3H+wZThLtmAXlgAozk+tPSUe4o4SZdWb1uxoPXy2V
Y8S5p+yUFI5c/4DE5znXy86etPjsP4Qsb1sfjSqfbFyv7Jj5RaK4bxGxIH5ce9Wd
J+SWbOcPl0TBCED3kdAYeYHQFpILRqMGN0nzpEUklCflMiuDfVKaSYBK5oQp3FAe
ctYJ0xCgK6F1G8TnP6iCkGGoMpvoQLrgIypqhpEhkw5qI1boV1aNpF4Fx1aznSV/
qMaz51HFToSWzQi2UnNDZP7wqnD4wHXRnapYU5JPnkr2Z4wZWJ8AY8889Z3AKkWz
g7YG4H7kfRzqiYp+mnf1kEQkHskJio8ufp2e7Zn/W4eD6KDfaL75C3cix9cgLhi+
dUehdAsHhSUEyWpXSO5kEyiefn/fYgIacpQVkWmSFIgMOVhZgZdAXronfNZKHZA7
UUEXO2/jRLSeOgJs9Tzk6w/1qw6fHdm/81jZRGw1xc08xwYaT6OIvp2KMPe9lhhz
nj5K1wNrmVGUEOiOmLpNJjv8uzcvTrw54n3Rddsecv0MhnWEpFDikHNSNUhsMAbp
Fmu91lke4Ar7YptJdP+Y1u5AUc2r2xcuB45bkUbUVmNWY/3D334VZwRbCkt3fI9C
poz9oUH704et2N8dePIk07eXUUJqlWH5EgsQlAwFMcA8BeSU7jPzi0rT1OJ+4bE4
Trw2iAvQ34M3etmwLpB5o5hs2HTwPTH1hoy/+CWgq9qpI8w0BRg6qL93Fo3pUXu/
T93RB4re3BuhYSh0qUQByD9qPSYV7z+vRn8gygemMNZyqQMVnIchxBg+1t4+U2xQ
Fhmwz4EiR0cyuraBX02ySm1J1yI2SNUUGrjj9nJGAt5xXvFlvbH0542ZZiVKEJQS
ZI5pPu4iZB4NXEWCOUMdvOBDmINFWxTwhVSiEWNf4jFI8cjdv0aA50+lwcXMWHYx
KSZusOgfD1XFznitAQESNcDPqAmNmJG049RbkRPx9TmUG9yjQTjD0U6UDQHKC5NY
8eg6X7cM0Fnu+JdBg4JpL9VERi+9BX8iZvYI1Cng2wsOwniXMaOLDhA4h+dStJJH
Pxqvu85dHblsNEYeMUnFbYAJg7tgT80n2JTlcbHtwajXmp1YJn6mOcSs7DpvTL8O
P6m7xdS7/E2ldsz/PsNBhENH5NOV8mgbAk/COI70IFKjH/4GvQ5UFcfE4s87f5n9
szRVdWBueop+a9Y/10gi6AldJw/inBIw6iRg/qfTfFA9pVLQqhoecQMsB19YquTR
elnIiPiY93ryx/uahRyBis3ywr8wFqyiud7pvO9uQKnN8xnjdr85E3B5eRDByuLc
tx/07OjrXXpqv5N+KgerKaOLnnAWuBLFqmCS1WxuTDMoXLt+M+ST5SZvjftvqGGl
gANViTcqwOFqebb+dGHbO3mR7NWu2mu8kAkTFxJ2A4V5lhZf+svdqfFBPpvIJ5zh
65Xa4hwHC5JJjXGi1vM5Cj1Vwj1W2zd+WBo4XjAI9KhvwVZ082cgIUu+MuHDWTn/
gQVhejDeEc6v2RS2jAsoYzYUiIbNfEzgAnLhZfOJRgx4VzSuWDAwug6Ki7OCueSb
f9cpubV3n1w7vKeQdFrk4lgcwkEHouMov//uy/itBAFoOJBb+3qNXdZTRgotxYkq
Z+cMz/eYCRF0VQsLZaurQ45DLMJX/BbeMUmP9uPu+mIT7PfTij1cFeDLN6+gggmn
+V5ZWbcMXPpvBYFjRze91yaW+RXKxg57uMZEX25owyp3OMdpEGYdyZxZDw30q4nZ
zvnRCILCLITJ2rhEi4pO3ZyV6mPCcUdHYD92oggGlBZO4yIVooXeiiMyQta76Lw6
gdDW3aKcdGnjc2CuAJbte1m1E+TURutK/KU1xDbBvmuaLAT8NZID0GDXc1kggWJT
zBiiYgWKKRFZ4SLuNXKjTOLKum6XQ19PTHfGKgQ2tW9cOxEJXA17waABngpUDk0P
coifxWnRRVPrRBpywSmbEG83yERsViTZpoAfNkgQdpuEVtv88drxXZg22uF9VnQr
veI+JRQNj6n2uI3gyuEm0Fu6yg4cY1Kv255uBapJqGUofnw1ScODishfD7PWCy+O
8mI+iiQ3e9O50taETJGUzzXuRD3y2eGr1BQgWGoQ/Un9O8sF4V/+yANT+7OTkNdN
bNSFgc45iIWHiijfZ6zZ6fWX5aDCCxz4GTQeO30ABA6xYDWP1r6/ovQHp443+JqU
ZhNABBeI8wRwzzOxDIcAsdhuQZEnIzr2sjGy71DzojsF0/kua/HJdf6FyzdPZPKI
Sipt+AKgaxJHjFkwn4q4j4Y0zOmcJkrLtEkSjSboLUc2HCKwsioGNc3ES/CDos7W
oYwPvDk6elU4pliwrfbNrx5Cf7O6gW58XHI+omxXXYnN9pcceuDhBJOg6Gt8ZkoR
g3I7Gn39jRyYmDVLDfR2y93Odgm6h5in3Fu/+JQ2xQTJ2iO860DWkZru8mP0rMAT
+MkpSneRbdZXDYt7G1nKUmFeUv+BU5HNfvZth7oan82GLsXftk2EQqHTiuNO1bzN
bbio7WF2+OQWM9z9a958CXZpoDbNM5qWnxHOKwTnBYwIJM/Cjug8JSFrHjVNl3zi
/qHbXxBraR/XYLuHK9B4sjU3qfa0rQdntEyG723T3N9hOuz69TqhN8spKTYxvMHl
/7FwXJud7320p6wdiZOILlrQ8aYA9GyC3G+14lxh3h1O6697Q4S/vj6QHdf61NRs
cAgOUKc12+6raBW9z/d68LfBrnkBfRcKtC/QAchC/NHDzAwu+rCwEc0n/w0mvhG6
64NQlSHjyOml40PHtfAhHkj9icSQsa3KP8hvntrk0J4DZJNaKXTGm+Pvp0FfqI6v
HbuSpEs06HQn7A3rvjedxy12yIZTfhLjWXBUrD89tNrlQIOxeLG7oY9vt/IdS2zG
6rFChAB1olUmwgE4XCxhT8OqJBXnYLRk4G6xFcOVksTt5TbL2P/KgpFFdBraUFjV
CwwffTm2q7Nt1rzQRsHKhOZFnKKv7j8c0wCd5RlonGG6rIUD1++jjttuw6Teqbc0
A8THMZnUAb34DSQPLPT48VvV6C2/5tnsyksQ7UaQUh/nrpIqUvKpe9cX8Y+jJV2y
xRTUTaTyZUMXH6oEgigoFREht7mJsgaSyh62wkjOWUPDjCEeEK2VloABc+lndBwj
e7YR7HcX4ziSblduOTDvS4yaESGVBK+xWF83jJuxTJUk5Zs5ZDCSD6WR51dB80QI
klYXFJy7ON2Dk1nLogFDSL74NIzBcwBqyi8cD4HTXFF1ttomnOcZvVQ3ntJPae4M
3rRInpE6Cdf6gx5RzQEaOmGBdGJK+CUuQKgcTcL028aQFth3Bb3/IsDRtVLcJsY3
AIDBL1e19WWmqk+fxH767NMzufC7jRbN+CtWNixt3KDgOLN7ahoySBe1p6ypDaal
nUW+kxa/ANTaae2gZ9Wa/0C8ShtygxQ91tu/CS5QIyZAEGgdcZen31zarAgEMnX5
IRNYoLyZWMTWDiMM3kV4zuA77KOv4NYyvHXbjWwj5rUT1BZa6N+EKphKat2zcuzq
jVJf6q8QoVhJhfhZvlz9z0uk4BWHTJNynWuQn700PrPAqIMfYvBZIjyRaSApQvh7
vIUuZHFeWheotGRdcLzvKJWDLuklyyH9XZtjNiLvqFjSW4IIgs0vDj6kRlM3SFWH
yu22F+II0q7avrse/pzee8zVLVi0kcYbUjqj45zCI3ue7GzgX6cf8BtCIoIeyAul
49bJZ+OwNfmpuHDVSQwXUoeBvEei3FZTGUwOIeE5lV8OL8Eoc9OA6NrBy7rPsQk9
VBLJO0PLkkwhG/CTltsLJwqZh110Xfky4s06N2bQz6Rmy2wkEG2lPuhHU0CJmRu7
mT3CrMf/K1I7MWmDuv72L1a0E36Fv9/yM7E8Ec9WII7lEyAohmTqngwHJHR/eJpB
BoFZ5Yyq7FlCJ4qsl871pvWZf7/z0duMJ66Zg48qXHSyZONDtQEVhLF7TBp9Qf8c
FOsAxq5Kv6KQ4GO5iUgV+T76CqHtDJA+E7uAbl9rlek4hHAJxwuyaoDs/9opvM1X
ShtNpeG4HyiKpFBNy9t9RkCE9qPBfSeny/QmgxqLoikjMt91mg6LMhFZWftP9X+d
Dw4HY58w0MsUWt4DT1Vj5Gvm6cZ3SMLjGYF1HlRVmfUqID8XeQk5Z1c/9FORcIFW
H7XbntDz9im8+XKB4l7rNZjjulMnBkzYY3s9ARf+xHxe5ECheJ+jEDif1oQXZjpS
iUawsv0lff4fSij9+sBYUAGrRKtJh7d4XJDCkQ06iXk2AENA10LHMCcAQb6kzPHt
h0bKhFcil/soBa73YMP9vsBsLCC5650kOQe0rF/o739Y0+5GqmJeBiazDIdcr9EJ
T8uejBRWI47hq2vD/38K821BP1oDp92Qx9f5VIbOtEEoh1T2fz+zQTCzBwViqXmm
53LbrtPoPz/cjRFQwhVCx5KUZSg8dp5TSTTGn7H7wLmHuCQnoQo8GHGZus/EAbaL
blQTnuv4GY1ELVZhLTqDe5oI7LoCCO7uWKdORv59YUQf8yvBh5rHYsVlcmz5WdUw
xTrv5kVbIuweI4QZ9ecVbj4U31gOo8zOAiEgy5DYMpVHQtmRYv0KvuaC2thVtEiJ
XAM7UN/qwh4tfEs8qHYhVoS8FZZmziIre8pnNvm8w4WTtTysh1kZ3rm0yleU4Iqq
sopy/pPTWKbZBrSud2FJxzmJSKj9gpJroMbCNpZmCrvzUHpKbDWZrc8ODQ1MDz1d
aMq5Bl9QYztr4JdFxliOKlJzl3MMJA88RWVGDp8zBcuTVwZGVxiou64GraXLLRk6
vTvaxpIek9AFXVLZgd88iu/Ad7/eOgBZ1HXYO9tJf1AtUP4ZhwofaEitmqUTWY8u
JmpZIGD4W9HY/0xziHQMk7FLB0+dqzhv2dJ5i0HajO780AekpHFm9wtCEtwE91II
qaxPEai87YtSKoRbHevnr+aYTwAphFmYUZ24KwnzF7cR6B6ebWhEXdOxAf4vbRar
a7LQ84WYwNAMCigm3pPtFEs7CY9FZXAAn84y6fsEOwSWvaxUfmHdUP089CL541jn
eOPtifrO0kSAAMurboWaOk1AmUd56tZU2jp99NA7gc0TgfwdcC7AmJ8H58/1R6OE
TNfBKCSW8OCmudGmul/cSiA3zFaB5qVadVcTbiT+pQz0SK9cv7zWGrh+NRCJSJGE
upwghTL6uMuapgv1SmSgwgAeUSHZCtLhlcN+oyxvs5+rnJXYOpqf3poTSd9O5RWb
BID28p6jees9EszeuH5Hg2G681K7U05C19Wa/DK7AAUSwnpU+SBqfnPHHHqXGPHW
Jz4mj0DR1tvaJNC6jWiHMAPlOkMAMZjc3YfKGOVln9E+ouf4kyagJHPqplz+vISu
a5BpFDj8KX+QvqiFqBpbykvCbAtPssnGu+gYWDdJh43R/Cr90kXRBy4ioZGgHhfO
ZLnquRVn055fWx7FdUd830eqgi7cW3z4lzCY7u/2z+Oh0uRiI2+q7PbPQYaP4Wau
o5eroliLmPdwBkj9aCqoXX/f6/BHgnRdqnWtNlDECnzLUfrK5LSmTauvIk2fG05P
QwNpUdkIYcGpVXyKY3Wn1C9/yH3viTZwIffSYCusPasPt42kLSMT8HLpJv1Ogag4
xPBeq12yYferhJsTt5cUAIkmK0U2kg6tHm1p6Y2hxl0QCJtgKqio5U0+1CrHyZxH
fdMwQKVibi0cWy/U+fxAtl7PzHInXPiHIoICn06Kdvj4LMoTdthV/GI/2lOgs6aq
MlkWiDWTcsudmPrikE/FyqaQ2CNIeCVWu0jREDxtDqncwVvzwiuTc2Ail1xpQesV
rWlF/VhFgcjWir9pbTwIZdvBig4HVLWGUZwFBl6mtPqGmifSUL0cltq7xSKDKeaI
sPIY1KVw+PVR+X/3vSv0jiC5K5hPptlyxxPYVUDkOHAqBR4bw3Z+bi6rSV9Q/Aa1
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
L57mnrL9pOb1JL8FXKdvKXVlLDKPUAZRJ1B4hGH72LqvZRZunJmCIKCpRbIjs2Bw
qaHfgqUD7mXnMKQ8n21DudeTEaigPmUDEIkebvrIsk1mg0jXHD6rVdUo0JWNU7ft
rVRKJrgefHd2oUszbWEq4lL67/ef3tk6XoXJXPNW/nf0O33giSrhDdc1oVyFR5MA
JT8Bolf9UwX0URHGcoEb+pxZF3ga+6VTawriHP69kJBUOwnqE08UZOKpm6cjPVgV
2EWBoFti5ay7Fo4S+Zy5huRlM9Uq9K1MLvv5bUWpPyg9SEWNT6qZSsvnOl0VPnaM
rzKdz7kjj5+kpqLHPBXUaw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4768 )
`pragma protect data_block
7A5niqs2r7VKZ1b3f3gGlwV5LezZ4ZdKjUDrdA7s5BynuulNgGts1EIJHmApnVp9
ILchUGaWb+LkHcLuzztsE85MTl79pqd5qnl7+WBAypc1JqUU8qcKlF55nMzwIL8A
o5B6K6X+zVG5mSI01aG1sFxCaOz47EXi+rHB9afil2yWU4cjJg6VxefQh3Jeovkv
X/A4OQO+2ziqi0eV5aduunimCM3Y8IhXetdL1xNV5qVXkpjjr7z7h22bPqMzK3yN
6/68VXiaTM1X1KdGlI1TjBSFJ2htSvTUTzJiaz0rSGjr6d467TrLMSILqSfS6p19
vOuBqPBTP76813FSf9mrLsj2IRVkJte2LluV6QhGamprM78iYsKSm3q70YCWNdrq
CNopBZRfTaq4a8P58Bko4paKXobVJj4fu6bgvxaCOLG9Zmz2TVMxX6Ui9ewu+UQx
Z8g/iyIwrlhwfmcWcgnfbasPhYFeyzN0DUEL9AgXoZe6BSI2Vm+R9p4cN+Cnz6wD
r8SEqPXq93x4fhnV3rcC1/RDRzq8mpREg6k6YsOQUMMVrZCnH71itAVxvv2eluqO
VbhjD1RGjmSCiyNnpIY87lukGwWZ6zMyDxanlOlF/YBw4KP90/50FgyER4cNCiGB
1gZM0FiwN8VHp+f+A6GvxL0DpUt5Msq/rhLDmRIymN31qRJ0PELOoGPA9nv+hPG6
qZ3RreAr7nsA7VuwBGsr+Bm27lbJ5ftSWg1Pqxms/EhNPjtxf2bv1lShfeeJklna
r4wejraZBQH+D6ynh4Aigw/v5CMWA3Lzuoz9mTwtX8kbuuWJ+5y4l60mDBIcCCHZ
iX2N6ap6INm9mjk5y2XfhUtLgLqyin+6vFyPkfRbeHbsmc+LkAlI9XBnsNVRW7SL
bNtxCLxnMDqRquH7uBx6iPWqPV0Enxfr/pw9IwIXqkDvvYd7f5zaPq6DCRbv5FGN
VNFqX7DpZ0SBDrHybP487ZFj3oqJ7MeXcDSWvn1heMwZspSrizl9v9IWLV4MsXca
YaqENh53/Zb82Fw/l87dfJr7orqsdFaGw7hB4E0riYuiT9TlhrMCRzRZ8gjQpc5n
jgamICoMruavOXCu5uaT5MedtXP9h7ps1eqbWaVAXrSYMyxnbnrXNHU8tGEMn2kC
uHcSUyp0LnkIk4MjqREHJ5UwzrszloYpYSh5zBmz9gEswzShjkR9EWYJL1gtela/
wpMcbChKgZQIbxHi+zmqSxIkK1eb6AAY+h7cCmvnWks0tWMe4xp/q2BnUXNj3aMG
RL5OSRuKNjW6ohL3iZxkU/9p0E8O7rmZjl0d13KGbySe0yij83OW2VAQyB7W6V0h
fIVCdebJTH7USo8PPbCD7JkMqq8g468fJtO6VFS5TQuoBkRqgkjhC5CLBilvY2G/
tpmlMIgIbE2VRSC0LnYs/LfjVLhTIv4UUmJ89hpa6lnEHlAi8/cWIX7O/OlKSLN7
NHCsyj9IYpCORhtdHaFBBKmfyM1cVrr83WnrMdIOGqiyToE3k3bGl8YDtSWvddUf
JLGCmRc0mhJXd0RrGRh/0WOljZ8BH2ErDxQrEFPCepny4X2s7Iqt7qlUm9y6PzLT
hRDDS2+iedZUfbyUU2+8vzqCLeZAKhdmlNljK2C9XjH4yEQ7IhXUCXwikYzze4FC
IndQWB9drm0BoQCGR0/jvdEUQyf+qSFxGGexSHscbARMHX380kdQAB6P2azCaAv3
tlAVenGVLSH9AgWtrtvYjcylpd/Kl46RsMr+Pc1MnmB2As0OSrVqwVcki2IiBB3P
kmMAp0K6746QULMb74dFdFdlWGbFYi8qJY5Bq6/oSR30qILAOOT7+fAcCBX26xSA
8nXz2glK1l4yEOarsOcj1hrVrEg+qeeV+scDIyG26IilHRG/OR5EB8wJ0L6WnV0W
UNYmVqPiKS3MNrV4q5nivtoZCAORGHsRwrPUdOsQ2yM3bnT/Kkyagyudc/tJbDpd
6cSvvvTbysBY8m7vwQ3efbx+t+ud+v9klmHGPCqow65ni7UjE6vGpk/qcUDNiotX
tzrB48SHhymyAbEKMLctO57I7ifnb6FCxouEOOLTkgcIioSJmn2osm8NUz2N+H8u
tO7Dxg3wmow9SUX7QWGJJNxuA+8WGwg3AsTLCAELMUt3i98znIAF30AWLOFd+1CB
GBbNQEfmK3FPRIsZPnXz5jKkS6rcawXbxQP77fWdK7kY9Yea0gCu/tuGpcRgZFgH
hdAk0ErO+pdXlkRo2YhWuDDFj9eGH8LEA1DbOOvJA8QeXk6x729+RF0xopjGZjtA
CWdNO+MfmbCYDNSv1AHrBEIRqK/XxfiUvLtNKa81jETAtNiBMDKl4lDtEXsUTlyg
APGY7LmMvYGb61LZWqqJgwP8hbY/VwnpqaHxIet2rnLnH3oYvX0w199E7mx/D8QY
Co09fxdA7Mq4U6szKw1TenToBjQQNReXbi2r9bMzC4vWEBfwrCIOL26Xnjt4x9Bn
DLnOPSKn7Gf+65T+tWgpx0I8/RsQNcI1bDuRhhMCbpEDDI/3Cl6216mhea+uUciY
4PtxpX7v6Puw4DhFyfzxH0P0LeMQA5uottk5i6d1PubkVCQk18vbC53LIHwykRit
nyHcJ2T4nFZKwrFQf2jDn6b75Su/IKjrpwoqPkR4vU9Re3kmauc8iynCnXlQ0r6i
k1oval8GUbhAq/VFW0Bk1xONd3/FEj1TNyi3aCcg5nY425PE4msXs/yYmb9GuLS6
QN7jaYEX+gzpaxP55eYl45Vp1aF76BETCYLHO59g+k3kmAPsr3xPmu0xqjKqCY7o
le7im7n4O2VHIZV64tS41p9olp+lURYcaiz44vSVqZ08rqOq6S/l9AJ+zZFn9t6m
V1xUZHAzCyF5IW2a8u0u6BQhbS01QsSvGjwaeKJz7I3AdVG2qLSNVW0q+eY6VCgz
ZMecWGs6tZDBheQkbryAmFkTGUeoDpQBmTJs7oZOkHj4lvjt8OAnKAkQOZm94OT8
b9/bLiDox8rIocUi7KbJHvbTAVnHA0as2DGjoB/9QKbGUfgfczcdEt54NItJOXf/
iGyrOdA56SEY0aaBr8jdl7XQ/K9iSf+hDyDzf9Ho1O4CIdhw12Z9s4yhfuQdYZYJ
LtF6p9mzBU/g6qH0jeW7R0tGMPoGxl1EUdZoOz0nztXZClM/xXaxpgLXpYQnQ2Wd
eUz295v08Jp4HqxpfZpGUqKh/lrulTP/Fp//2GvKbEzlEs8k7Y3HoJ094XBR8+BL
p199shPMa1sKgaXoLplddsHQjFvIuF8zmv7sBULlehQsjRsoTbwLP5n3pZS+DIKK
awJDygBpt6xAiOkoAFKtXkKfOV0V1HBuM5ittKUTOAb7Drf/mEAK9s2MfrzayoC8
p1vOHlP1RhqXRvTjJ27jTUzy9id9eTYy+U9UCbU0lJ3eAnRaxEZr7OSn1wvLOrA7
fIXqOLjrGOWGLs/vvnUY4NgY849UH70X5RVe0q4rKSLVrR6iW/eIrcdVmweuxPzL
ubpPRL9dpWTzQEtrhEgnDmTpjG89LDv+nz1qrYhxYWeY9akckVvCkIMkkrjDWyQb
iqaU6itt5aGNzJuIgeXHCl+B0oJYBxZvVVPt3gwajPbXHtQs4gBTLtf5VBm30CIs
McbshLu6pMlvPoMQzJqQHPJH3usNOYMzcG0Z5WbXtpYr8bMnCfGsZX7ruWfsJKrh
tUK0UCWnVGtVT0wDEuxsOUl6RcMN8ATVHvmasXAssdRk3/sv4h5SfWjsfUP8YlPQ
DMz+CZ1AsJ9NN6dDWVFKGUpJJfBUlEoqqas2FDWZpyC+zl9MuU69gK6e3bfv9jQn
pfm1t14RsXRFoeX6FUoXrQR70AtfpCYQE31o8GGsQZH/snyLl1bs13MdKj7tekrk
HE/Tsi5L2b+irJh17fmrPamK+55HIbHv3gCcLIDPC007fyrkWXJwPEj6X0+6VMFc
FLmK83/fxxy7Zy/crH9MGzzQJrRl3ZB5KDQ8y81MaDsSfDPMnKMwuaG6iAFoTsmb
CJ3ITu7tXTuxOWucB5oYTLIdravmYjQjwchrbpLg8DY2HT4bo0xqoaOYTmPj6VLR
NoFHHgyRXOfDk1TA1obyWwzdDgQaFz1NkAXNKEwviTMBNaVfKQ+dR2/IT7iwiMio
2kEe8QBxgZNfa014aKCUrY7apD00WdcrXdRjRlXFk7gUDJeYxfT/wqmJvbj5JqvM
dTYrgSN4Rjtmhl7bPUw78MmzvkpZf4WlSU0XOLKHTJlFeUDZozX7iD1+BM4uqN5a
4oXj3yNto79tQeoLjycOBia6YEc7xkBFcG4+HxSe8IeNwf9EBFNwQCOUVSLoexCa
rVumg/mlU0mVS7O3OpIc7ogZYNcf6sC6C+GbCljRxwt2nxwKjnjwI5UGQp87ltTy
ZPX2lgon5Pm+/v8ARav/2wOJYP19Il9WQKEdUoQAMmPMmxZsV4MzCu28Fz5+J1fq
UYMUOhpyigqgYoJksVBaiGc8QyM7K0y8NhC8Rxs0qJ+XbihA1iNvcZU65evlVUxK
b6yT9UTmHhnlj/2fHiWSLcu5aOYq+xUzsGyvHf0ks1qQMBgacBOIAd7dDic+jVLI
PgQmW9eaqvc9hUpeAJ3SO0HUyaouXISmcfvKOorplX4RHWYOE9Zh2wMNWt5YrJLn
qq06pTnPbJfa6n1zjXIGnsIlUR/vCMcD6T5CZsMLY3N6vuaD7sU1TiMy7NkOcZwS
iHxvaBsbzRwCz06RYdrnWVgZ5RrOCPPlCwNxqHKOu5osmH2Djqj50MMachbArg6K
QbtZTjnQIlJxPVa4qp+EJgK55fOQoMbfLsjJwTqgnHGIU36n//0rLh8FsFMsGdqw
z98I69Zm1lvGQ+Mk9sWHIsLmwIINN4jBsEwH0wd0eCqfeKWdt4WS8gERfuzhMR6l
0Olhe0sVnIxQg75tlb0i5eq/dcDEktR9aQ1pxspgx6O42lDsDGwoP+gaSJFkK3JX
fUtQ478DaiXZkIqHVF0CsKLa9F3joCp7JK/tHtUXglfP73946Ye0NuZz8XGZUa+Q
oS92rx/p/MfKhFk1Z/HTqpsVVKehAKiXRGyQTBdMiZncPTp8r5jlfTLFqMIHaTJq
r+N6M4EWS9EHu2tUptDOM2Zp0i/0bjw2jmlW2Ry0abOnwW3uGq/Seq7KHpONTy9L
ztXkr7ipQf5zd0AWqPk3G1CtQfK9hiZ6Lmp6fjqYAb8L14UVd5p18u4ntkXFuL02
nUq3wdZBwsJAzwWx98lTtUpKQLNK2G0mfd7RsB4jQR0Ff7oHmG1GT1feS3rdmumN
DabiYCl+RwARAsttoV8sOzL03yRLe3YVaYYfAnGdLkZMPtudHJMSX1dmeCF1v+Uv
OkqBf2tPXEMlluadSLEGU7/UEA6H/O4PhwelpvLMDWiMgvC3+AP7ApXTB5u7xqQ1
lkE2uVNyNf4b+rKCe62j7zGFnYtFzZ7BT4mhUKSWsUIk08WqVdUJf76ctLwhXLWD
TSn5RXtadO0dwHIE/cfrBE8hEPvu7qrUfpzp2+lClxKlZXdLkpi8bd6xBfUZ8Rlb
5lKda2x1JdDFs4fzdUhi2Tm2VnBPiMbyj0oNPl9gz+EyOK+l0ZMjah3SirYwvEB8
w4H7RHukjRoy8/Sp4O9SnzeImsCp3mW14iRTF0sL4q/bCxGHKUk2hr5KRooFvlgH
W6Q4aF7em8W0QJUfDL3amsAce/OgPDxeTSsUFCBJsO7SwEDS3TMvs8Sfbf58b7WJ
S+vGW1efOkxIpjPtAhIe+iWtEozGVibmEbrPD2hdECc5Pt01MABoIRKsZ76QHbK+
T2XFwFMoiroZgMJZ7yfJPVpW30CGoAPsKYmSU7Kd4u4RHYkTwDiJq8nOyAsJiN+c
78L1Oo+X3iQ6Wywd6ys7xikq9XJHty93etakEKZx5aKb28l62ONFb5+RpV4xRA1S
Alypt2b8AcXlc89HNZyA31IEn8usD7jZiPmXEGx8bm3tXqSXPEOH8tWCuKM5kbM4
xMzjlzAYByNWcX059HPATG+pTKmb2Gayv63Me8Tsrn/IMqsPMl7eTiZtPj4pIrB0
WJuJArXtK1zu0vl0TqBE7kttpmrz9lC1HOUvX0WThCnYrPyurzROiDDSPvZ7YeXu
ENOEXM3RkG7EE3re7DhnwrQeIL5kJs29U7u4gA0hDKv1zJUSzsbUzNm+JcFoJHL2
1lFCYO+EbDUFuH1LZDswt0f2e0foMt9FgZfoRz4qAOtlaYFdVz8Hf908U9RSCsrS
KzYm0HsbQI+2j6EihFRSIyGQESD9o3Ur5W6RKTMRQ306yENPBQkfI5PXcb7dmEtS
tEHTCrD1EIMuOrXFWiOihw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hw3AhxSuabDgyXX++4lpkmEQbSeSgi26QxXzSi6UsQQDpCMSQV+jlFkoNgw9/cmC
LXiyE6g2cUaU7NDB1s5rZtUajl+cVdJtaTtRpU6LGF26V5KZOjDbTk/6HO7g+bcS
kuD/GRHjq7VHJVLaAKdhTXMSkddTUGtIRXIPAPVMtIUSNHc2ic+OoHSemqlKP4ur
N5IqXBTcuFzdtnsg1n7r4yc6c2B/4s3UFpb4bK1RtpjvnBzF6O3psLkxNjlG8Z4L
b2kwQFiY+ucw42GGYcCH2++Sm966+5+CTwdyusMoXQAQLRmdU0j6udy1TA2YSUA7
Z6fBrB3DDcS20AbEQejarA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8720 )
`pragma protect data_block
w3AL+dlyrBZWtaYUSMzw1Hy+1weWLFLEcinoSBykmBcbIKbTLp585VspoaXJGXmJ
kPJBa0LOKYloXCZlukHAptNksVyRwvfRHtTYox4tSOIZWxPZGRJs8yQnGNd/nySK
pRYmtiEIyM6593wUB1HWRzgWP4Jb5ii4NIMObyGKn8cumnsQuujc5KUIr+4KVCmZ
4M7LYnvukYPoHHjxlm5HPEBSsB8sUkHHH2mY3Mce+8af6rBnYWcS01IFmeVsTAGH
fl/OYNFYZwzqzl0EuDFGR5Xi6ea0Da1HGpSdlxIiqcSUQe4/B2HnObNrbTNrb0zR
HMZQGuv2uz644tpclAdatIjETZQqt7oOxLPuEA8W+usHsBJc3c6TREuRGWMlgXM6
0Xtjru4G+psXBwj3dSnpz0BjCFLbkFL8RZjv2Y1beScWrwfTJjRXfF4TF648u2BX
cffRIV/57Q37vse9s836OEeu/attuqkFJIPDUA7MVyDqFAMDE2ehqR0gGno/CHmm
fBnaiFFBVGJdvEZsTar6pw+uJTdbOJuC06uB7xqoiIjI4Z/5AtaffIfAbgu4EYLk
UocKydzyuqGn3k+JCyGdaPL/1BlTzFLnE/3j063cSW1hk1h8UqTUf//lyO/iL63Z
PeF+ZFjCeZjTi4nhPdVGQmdKKEcQzRKCMghNfk/4uClF5tt6kuaf+DFTDcV/Y10p
chC8l2oE6AYhbGZ6utJ4PNeI5XcgYb3CSWda7yuWLvDM7i1RDl4GhLqffivd1L0R
d78Ei5iHY9IIgSM1EfLff8pB1paZCpNwvHuzktB57WdtlpXmFCQkmu3szHxBrFYO
kynxKy9R20SMfE914FAzhTpWf3KgxLjQ26z/7BeaZo8z7v7uHvlKH/z3guM6+IA7
YcK2aErWyvGYXUZoFlx9/1xYpmok5pklCO2/4GOWwz7FFRScEfPRDf9IT0qCsqvC
ZbMkgVYqjrLUcBdK88Vo2fWGwIHVsrYK/xNQNeDoxyE1DrwSKL8JO9ERq2aWh1Ox
BJ6RDEbsgK6+dQI7D191E+aK6wqBgKWxW4tBuke0jbb0tJtJqIbCm4OG/MLYMQOf
/HzgQVqVv85iM5tVeUmwwVUYcEgQwcQgKYzZexvt+iNO0Kc736kpYPxirLTmYd00
JdBqtKoBWDyzQ5ZZpNuOyFJAASYifcpcBgN/jY4e5L7sWSmeaKySQFmIvGar6T7o
K1o8VkG+e7oWxQjIIvVWPnZeDT3cpvxdp7lGtkb+G/Y6o4+kGAhUnfZ7ZnigspCG
KH2Wq8rQeuTeTrdvhIv65RoJ+pXzsMk3yPl3C5i58jSS+NE1b9cVtBenwsGJeMbw
Eco265FmSIQhNBd4yL5BvQmpt5JwANrnIE25P3MpCCEa+s+9d1ofA3V806VaVPQg
IFetkgFFbn/hiLoFwvZglGHCjasvzly5Tj2Ddqhi9iAkS8U86ICP58D3FsUSX3ny
f/N+sqWGKE9XscmwnLr4E+Uq3Lq7G6k+3Ku1SfbncKD3nb/WRt0LmzK+VS+g6HR3
ee6wz3SLl7Ly58DQYGzgSMWqh0UQpaJpFvS/4hwN7iYv6RU6SzqOPYKM7NM1tkWH
EZ0LRqTY96izouGQj4BFJETAnq+DAJIlAgpLsqAxGN5VU2/HHxPO65cuJeTiDn3p
636N1rIlS8vBnQJ/J4kaxpc00Pq7cx2rTJX6BUM//aR/bmaY2fsLknp6YDM1smjP
+TujRtG4wYqpArFj+vHFWKcJwibwdXoZbizOQisMf4ywvh1E/cYrSbjND67eEg08
g9NDVsJEcAQolS3LZgzop5oOd4l/8SoxgWHEa13tyfXxQvC4MbC3vfYyujjJlcHr
i7uw7RRuembmCnGtIHkp7zXPfQ9rO0pDkZ4tnomhRhKzGVM/NFGt/4b7oVEdE4zO
m65TlmHeaQpalxeoL1W1Zbvwu25Gut9+ofOLXbxn5hVyoylPFpdMCRwDjhwKVaOa
l+yjV0V8UuQQeJ5+ysbbPHMFtZBQynTXDdhTJxBi+/AX14kiK6obqpoT8IdDrIAx
AllJGbccNcrj7ZAA8hVQHQUwz2RxIfB61+dM75BDXWxOZEp2+NOS2Of8w2P4QspU
6zLD8PdErBGwQsE2RxIxwF4umqKrVROkECXTSYsoNDM7XgwnsKNU9UmN2rjLNRoJ
X6osQ/iYiae3OqWHTdObtYDy8kPuLTDIjTBm6QpHI1PpIZyPzw9GfvJNDcK7Ekoh
9dGjCO9Hp0QwVxJvinWzAqzdC17fH5131SHCCVV5mBaFAq5M/fa45CdPWkeuKOh9
o3zHPL3ujUwN3cmjQJgUWcMpJkThsbRrLsTP2/skBMjnE9c5ym7lYn94nqKVe9TD
5+tuAgsqVAmq8QyOMqQ+3r+tD0wiM7deBCVH05TF332HCN+WLNFqDQFqXo3NzN0s
fI/9V7KGqnccCXvi8W2OPAas4uE83R1w4jnkNIaHVo9EzhV1GcIS9GlZm+uo62BG
T4M28L9XiMe9ZpxiY77gR2TpdYpA8P3gxzDPiu3EmWCEP00Oj5uHWEUCjfBPmt5E
GHu68DWnuXNQp1yRbEEvNZxtojyCXIrWlL4jThzjNPueqG2vepO4n/9U3Jbp6RvM
kuWDajqjGHVsm/bT3xI3JRfxLr0n+nJ7hfr+FPn4CqmhyR8L7xv/4HUFtq8o/ZW9
I0UGE1lAjDrdPtCt4L69iyhSNzCd84myROiljLz8I5KmEJuYj7tvc/IK4mkLpish
p9P7e/1PWZd4vwpr3ZqDsV+HesTGC2Y2ta/EkmEhkRlQVxY118QHFMj2s1fY6G0H
vAksRYP1325DIgnRS0OvHX21VvTUHMJR47enWKBf4tG2Sm+PLgNjos2IosRSPH0s
lRMMJYd2sHU5hTeFFfX+km2TpDSiOTaoHv0E7oMcUSS4l4Hr2hJ6GIPNh5f48I9t
2Qc1JAUelO6hBWiFj/5AevwkaMdZlXgP+ESa5W5FppWRYWDqbp18Ig1LUKEhL0+y
d2ga/LYDovlp1FcptCcSErv2YWTUIQNk5cVbEc/hWSSEwX463q/8Dz3Lpkd0U0yk
e4ee1qYkHj7rLuitx4K184qXn8iyCEwPvJyOT/q1fs/3E0vj8uWHbxGlUn9iIdsl
4K/FoBquqLv/0qpkeRqlZN6AY8C5D5aEOlUlB8f4Ffd5fQRlhm0JBt3QSw6Pqpds
S1iZXvu+0NwsvxaaJMhbSy8roGvAJeqtz/n3XiVqNm3Yue0s48y6Ukmosv344iOv
WAf4xnz9IqILVee0fBoiBFjLKXEgQEx0AfhMqg+GUaoRVUY7OF9/UDLQIT26mr5V
gHVemkJdTULrTAnLZdmfNadOzLMBRy7Hyg6ekxglC96TUdoWn2v2f/YL/RxStlWU
UNoyVaveZQokeKAE3Z91Lsd0dSrwoFQB6+peKsjXWtfA74PjoeCxvsXJHqi2YZ1m
OK4JZSdeEFMl8B00XMx3ThZFAUAxqI0woK/TWHkzpKK920S9JbavXT//DbqqRVC5
moDLBMI+jAQhT1M1Z55pZIO42TDQl4ii9pjn1WXfqAlksRW8RNPhhfj6j3RUuDi0
J/kNFFzgE9bJvj/96BI/w3WpF98ulCIxvsL+rQ+o0RDPnRmTVrMAuL//Wqcy+HXX
QM63WhT+UuFP6SHbNs1CoY2sXz/+we/SS8lBrw2juAKqDuO70bgBltbvT8PoYTOW
ttfz2EEBsTRn7NM6LOHNush7LHWECCw1AxvtJJQi8s1vcvxw4viIINo81XFlczn2
+zgPxHUpDaJLg5GNCtZeWEFeTtmmi+lJobv988IdgCDxIq30Dz2u2WJWYZmJtqQR
wF9DbNpYgugHoQ7BxIg8yW7XKMGPQeUtUJSNBNnbs5di4KTeBhxarPy4gHyq2mv6
JhEB+vPSXXdCabSQEYbfKEHemKdtD8z8FZB5+x38MAGh0nYQaymH+H/ZfJF7hOII
8nUVgFzsTtjPXgck+mDVHwcjU6Cikpl94qwHbGXeIMHDGef6Z1M8ogSK9GcXrv8t
MjS8CuJ2OkOWXdo+8oGFoCzRcnmnlFB+yfv57/W3GDLS/Zglc9nACfsu18hlisCT
TZW+Gx5qzC4XZhK35owaosxWWkYqGuMyXuwBPRC2/j2zCxWB1Vbv7Wt0NnOE8dzd
mgs14fPiNdcvZMV2Rgas7a0WFixpMIkDmzpBiKwtB9rfDFTHJXB+CYzak1/p7ZPd
f7bb4HttX1o2QuU5YB7u7oBdRszjJWVScd2ZvcocPTypPCt2MllRueyUcfO6cJLh
Zzo8dy5rVXrMXtZRT0+xTEzR/i8LwPE2yDP81vvAIkT0Z1XGvdwCBbBz/ukmJzNB
mucvyKw4vmZNHBSaU6YAaaU1ocskLDm4c0tsBU+6jGxmj1/B/1n3Ab8Q7QSDKckV
yn2LqFn/2wu1eymkbE9AxGBMZMvGbr/kPm9/9mg8QV1J8ImO0GWOWZA2p8Esu0Ry
+KqQuRILRweKo+rtrW0tBbXehyngdE3mfCDW1VC/qAEgaiLjs2riie5Z9jTZjd/Z
qEfOxitkkxxIzo0F53B+bRvyTuv8eedJdwoRR478ajeBYe3IJVY+4rhBJ/aA6Rr8
tKOChmSmbEKcQnnb/PF6dkFJ41Gr0RuDWMJWy7vFQ5z/JsxhrueL28xK/uyg4k2l
yIj03KrFSByLXmMie5UPl6AHJZPDJg43fD9dFwAhb5ggYJpvljmTvZAgwli5KtvV
SOD2xViJvCQePHGkvf5XTa7UYVA101Pcj8EIez6oodTzO/5VXkgYQSVwQrUSLpla
bRL/AOje55iNK4PHfa0hskvkqH7TJExKdWpi/tJZ4VKFhiyWRBzLyX/5ZLwsG+2t
2HLXIsmzFeDMiWA2cLHNB3u3LdxGGKC+my4k3ujfmSTrJU/AuGvtFC6mtHGgxSkT
QlSyH68G9l7TJAP5zLzjili9jSxcEEsT9BaJiLHrL80AfgbV+1+xEhKlME+6soKV
Vq5cSdu32BUR5zuPoIj7T7KykGdbhIqtS59ODt1C+HyjkJE4za/YpFScXwqbbnOo
pkhPbKuF6IzrZ2zUXMZxv/elTmFz8F63iwdNXjEQ4o3wDDK0RJjbAetXQfUiBDAx
nYhAPuaS+c6QxhQwe1/FK0ke2GFNSy540rmAfxqwesGO9useJ9WrTRlV37qZW33q
KbAKmDdBIU+6iJupe/9a55OuTiwbB1PoTi49pFrvcK2i+Dyynu2ERXvxmsItU3GG
gXWTLP0Xz8xPfayiEOeGMBSTkWEc5sWhGQi/aVVVN/Jj02yl9msIOvJSDfoaL7iB
Y7uATVnEBg+UhFaV/eWlmnJ2Wn4YftLdt+p3e8ki01sKZAA9pvOXLb+FjUuve5qK
6FGQgUy3CQOvcU9atZNm/1cWifgxiQYiCysMcNQQSgB1CGW/gxT/lgaOrT8wiC0V
Y0sXevCuiEjzKB6EVn6MeEh2xtgdcbWT/V7yedJz60OVPK+JLZ4aU6SbrUokPV1W
RRuQATDeI9pugUKV/EijSbXGUEbeEVAxul8L0+8rr5hsMkIoEOR6S1GkDtaTFWPJ
VEqzgzC+pRvnzu/fvAYahIRGGgO3BRap6y0aeg8SHxRnA0JUdvwud56qb+jIcvVz
myzNk71xSJ+/DBfKzSjPxkLlVVNhED7+tnzuv8Mr9hJJPMZulUZYcUc8JVybd/Zi
PSNmCCdfrVByq77vfS5CYyPO7W/z6ywvFPIakUPmrlFEt60mEr5XY/V4pjOs/te7
LHt9dGvZmiNXMTuo9dp1SH4XDS8wrC9gEbT6AIS/0sdailM43v3qwW6tRPcZO94o
nq183yFM3kFoVamBWB9Jb+Iqxd85mhVcIsbW10rQ9mc2BV4N/JvCMxsK8XMrkbts
gZORrZSY/B9PVJE4q/V7JQSY0Lrmq9ny/QSIigTsOah5k1n4nVE3xkAXsuug6zsf
OP7zAQVmDEcstbr91VLTmu5lWgSP/c5rc89FuyEJNHXWjpJUpU5djF+IdVctTwzv
8MR49zpGXztKQJOEZxAjHE+NB9L7iVUZVVdG/iYYQWFi4IDxm6KN5MTHvNz4wkOQ
daW6mVrOgc/4eJsA4EpUNqiFnmqwKTPLAXbs8mo3RciYJpcGCZ3M0c39lG1dmE8y
/JG+bqxuaZCySGU+CCRfeile1IjldSQ3Ln2lsF5Bx5F/mvejJdve77GPXkH5sBUO
fzICRxL1lMBG/5N624qZ8jI/HuPRFz4DAfKAOJcSesoieUyBy4KsUmbVkhBZTNx5
ewoGL6mjT0eCn/Gs0X1YFOCkMbV7DpgmRW6BwgrzIFuQwjqn/3Hk2doShhvbJrPQ
9hkURyFCF6//Lanj+sk1wb96GUKji55xnAsM0+cehEFI0llfjbU/ZzzZGiAOjhZ7
t3X1G8ydEHquEeNQVhI8eD0ykxbxesTMP7BOIzMDo2Zpfbymoy9dnNsidRTbEaI8
xm3LDoJTFe3qfFzGUQmIkwi4/rjx2QlJO68Kp98SAf0eJSVdqAyPGsNEEd0J8w+z
z30ZFDufybvaldg+4wGAd1CUqScKHMO8qX4gtkpmVbuig7zjzKOcUHOhVbvwgMuz
xkXr/6WZNarTNZbkbWzdcTVq7Soxb/s4mo+EkUsJWfjlLj1Uor5Gf7wX6IOeZpa0
Ww5CqEO6+LKkOIYrmyga7gF0gG4j2eU+j+S93aOf7M/1cg5GBrSjExMTkpYFK+K9
zGgTpAOV0MskRUVA6JT2r1UIldTu0o6gnO4Br+oq6OV2ncP/m8XL87R9kpzmvJnZ
MehXhUUq4Y/1is7ugi8F6cgNP3MeEcllFzs9Ncyz4JkY0Y/vvcV2I32nwXZwHOIH
UuSiDzPkjmDMEXKcwLC4ZyVm8oM86nHFMSGRyeXqoEeJYMfzqJHi6PHsuz98Z5Wo
vJyjaXhTYAxd19LVd+eoYYoNoER2Rc1M7q8xrPKvD36O71DJhJGQ7nHlGSw78inG
39V80RrbvLS7W6heAbYHLeOenS+kMJrJ4Nbsn4+kTohhKZ89hXNuCPcGUrsdW0y6
WZKoC0Ok4EvDjo+UkdXF9qKKELIC07iS5vPLhgBR+jy3V7VyjmtM/n2OSEVWIUQ/
T/bQmF5QdAp3DPe6CZb5U/njWJ6yDApwUndHZFMjMDLTHb4+AVMyrKdiVHQoCLT4
sFoayMliEQSRedAPJAzqufhv7EsvNYy9A6MKhcNIhDrYGar3oRyHCHRZ9iVnIOUI
/VIHIcCG5xhy7se7+cq16dbvce5i6mHp3/AFSYjZwfsFho8Sv1PcGCZS/83xZjtU
3AM6cSjvQqQ7h6PHeVmgNUI22s/S4AQ5/FvtBBluYzd1MK04+0KwBpT5J2sUIt+X
oRTUI7UEDARN8xXQiFJ1qOvjQ5ZyGktYDg/syhOfuZDhu/tPeDut8G3TvqAZKv61
E9sCq90fz5rACwM/MXpgdas0L9Rmd14ox5CI9sVq+YexrbAwzvleSJAwQt0UWpgR
8+YG8kbI4Iby2vgPS8cXZgi38NYB/BHjxmN4HPVdq5IJ12mD/MTdONiCUjSD0EiW
zQScEiV6vGlyNxFlRfTEd4+MwSu8Mn1lhoLZMp0MjNX37gzOF8L2mujn7LacbZk/
05ntX7pzZQNdO0yauXonl+KtlS3MR89AyyI7UWPml9s4HqMXin/oL2g2IDGj3Yge
AbMvwTjLsbxzDIgUUCAtcUX4/CqDYV42h8kW2YKm+W8LhHEE0wqQZbk0qjdV1AT3
zdqbHIrmQ3CxKAgZWYd2CwnZoPJ9YBJUvelUL5hpPVBd+qMbruM9VXFPZAkshcKY
nhpdV3K6I4mf5Ek0SSflaw/6lz+aZhGaSusfIdkilfSIeB/MrR+mky+XsH1b10fw
WXo1lJC+8X4FiiDySH8I4KCwYiN/0kLIpmoUlNNead8tqyaHSXoPzxeLTwfGqs+G
JUuBVEUhsoTclk5iGbSoNfag1C2QfEj5IF+xT/1gy+IPxQ9okNuiVHycWtXLKzzb
qxgE5oNsRwxea3Z9lQQ6ytV0XygAyjvg8k+m/x6bVWmv1U4BE/Y2Y7XKTkrJs/C5
TPufVgmjlOy9hSV8bv2IrAis+t+qlhe4Yoc1rarmqbVmLT2/SSRZLAdW7k8fy/de
JCp0kwVH9sh2AlzdTIvRM7G3oneHXFrtyKkajLpAW9VjKFUmOWBkT9dEs8ZJqLOJ
1gc05I5VWMfHi9MuGFrp86syeYlhMVH6wiCgIyKmbgwKonQufB9Wlb5QaYiSSch0
q+PKgroN5ufO4zydiP+smnOTXSaKDSlx/T5XCpJ8j50jCUD/wmb6ZVnSSoBxyp2z
d4GObP3IYvoE7qVSMbcUajRo2/1Rt0tKV+ieDP2Za26iRhyloIld7Agjn805O5JH
z6buS+iap4y/Yk/6/l7DVpr74OdjISP0kFWqzltPLWUilAVeZGkfFFtElIqFigVX
ZoFgvywMa5gU/W+3iKW/nvWUi5I2BeMuwlL9ObEgEJU7tFJgqiWWXXb/nnEnT18i
sGp8yC13awM5zsZs1zfpoaF4PO/fgjiYUWcg7M5uuLZTnQWWSb8s6yVKSSzxwSWl
2xcAZ05K7exgtFBVYqYFZOPs53lQPmNDRTZIMMOluidBrxQkw8cXI+fguaiBxkLv
SAgVONTWkSIiPEAGvDL5xL6o/qI51bW4tCaWx/nM/0hPeOZsz5JwOFiOYOz4tkZ8
CVORu902+tqPHysiEn95vcYDv2jfJm5k+LjZzjH/Kz4CRRxpzEWS/JHnEsPfdXAq
2721aAPkw/ZZ0jwDZmsP5zqAHWIE92bdamBkVLwMfxwurBqTTZOMD9Qd5YmXmNTi
WUMXm8OgnA5UzLpHWw67Jx1Us/7CLKLIXgmxQkcoimf4NtlOtmjPFVwlSIF6EghN
T6PflQkSvIz9Fe6pxdZuJxh3gsbPLuq8pRNxwHAnerCdEdtkHl+bjx2bU2d4SPmi
5wLHbqdxhOXGcENhc5TtSBidN20HehJbMshwM1B3JgbL3m9SvVgbkVLuU1ei2udn
9WQQDmVOQh3d2FV61uHStASV1vBJA/GVB8oCXUqfWz6AxAx412EfLNm7DY6l5vdZ
7EyFGZZdNIEOFGi0Vpv9jRFyVup79t7FV8u3gyecF703+e8MRejGr2FTt/+5cY/+
eXR+SYc1aVgx5XBGkplJFxitWTbXyKRtVU00YlN/+gyMtGxNi5iLg90Xc3pwuJyF
c3EomVOzaCIzJo3zJGv4toJiZTV70pxY4dsxw1wKZTJVO8+yH+sf56uV4eXPCY3i
XtwcCVcc/VriemS6HWcQSp0xcGuCZockU6zSks1q4OsBjEUCs6F1WakPr+zXK9WZ
mtu1iloyneIaQb5/wns4l6L0ReB+oZbp7jb4LiAXAKqUglM8cFV0cxLx35AcVU1h
yJOLvNY6q6T46y8/4+F9FndJtluGJlNGC3UzroJ64s1Bp6nOl7PS+HBk7sCVtzkF
guGsGDgmDdrNxjOiOwwy7l1aeauX44KpDk/JN7cuxlp68Ed7fHygZOc4pQ8zzs8Q
t6HeadzZZ8XrKtCV9PIHy1bexX9ez8gipu96m8xzJBJjWPIAXANOaFvJLE9x3FfH
FwROJZNM7KBFGPiy0XHjbOiXXO3JAxtDciSsJ0h9YGvHrIcf5Flpz45KBzDFq0k1
9JJKcn8Ju0miALKcLak05RWf4AdKS5lj/eOHWnVLC+pZ/dZDxaZvTMxUmhEckgQj
kUojug5lrjJllw/fvL4z0xkV0Rb45/HB1h9hSeZnFg120ei0p7QK4m92aXCRm6sC
az2YPL42711eGpQHkhg/L2hNowWdDBzDvh4zfgTwZb5/eA6tUPxMz1lmDXRW3OCX
/VJZ+LjOqtF3Ir3+UdXbIYOubMJdvrnUPle1in4syYL5WX5/vdkvpJVpMggJooaF
4fjf2ZrdcbXcbdwmuRydlBP+zBUu25FhbrD8mcGcb0XyGZ9Oksp7jNz0gApyM5uN
7fbpAfi0lvsi7dY4g2u8SLjLx5wmnMbell3A3T1rnBOe/M+G6aBNpwr5+HjNeCKJ
R/c1WXMgRZw3T4jgQVriZ/eLx+Y/OUuAoIL61Hn281PNM1H/mS9DXrigY8EtG31m
odp/1dbia8gE3J4395t6c9WdmbOBHUbYa4l8GY9etRnipF1J5vnHcO9J47F16q0E
9kZJIKpvXlL4FWQTGaoqhosylYcqxElLzOHE82eBlGgKHj2Q9QIy909h2P5IJb7B
iwWrZo0V4f62Ti4WhBjTfGNCLVc72vjskY5OpVT94zxKflq2kUkIMJwYOlZRKXO1
q0FSBE39LuOHY6I3xa2zZG2c5BjPWD38ZPL3unCJbL8aDxN/20oGJJfwJJR+Vd5h
uJY/Lbmg6UADUCjsFcinEALXeU9g3bTET5ecYgVGWaAut2Vt48bwPzbKihqGj3qf
xFi0y0J3KnuXqe+tUOtsQDAX+5FHXgaSvA2TbSv7UANFbqheftryLakogn+S4E6G
gpXGJCTj7ThLb0Y9rk69ntZqSZHDfalc5ecE2j9cfNkJO7bwSjfovu74biOW1E8m
eU3+MNvIVfuckiGz/p2zZnd1pm+j3wE2WglOl1U8IMAefYhq4rS+UUfAOl6lL+pP
KfrrM6Zzziv2nscKn89gsHcfNUYWL2w2dGuceg5qoj1OfPkUJ3Io0DtSTKRQs3Wb
bFeW4p2uYPd5xiQWR64Bx3953DSz6z+SF0jex35/beeNKpXMFOZTV9nCti0eZJBH
vh464faH4dXYBx2S54cG0z8Mx88buHd3Fb79mVUl+U1YVEUJbUv7/sGHDmpkoQsv
OrBqVoP9ItF8AFSEGbVivWm46GlwujJNR6MTONl1YVkZTln22N9dKI0gyt2HxfFW
3nQX56urLoOKatVGo+JtWQ8iPvnYC1zthD9lOW3trUmoVXJNe3bB0bsD3BQOrf5n
7lnxfSEBc/jupO4f5kXzUL+igLMtcTgE/lKRv+a0Ijt0lLQ1VgOPT0Y1dp21XE9S
iS9IQ29TRJrlZyQ2YIzvlP8TEys5bFrDno/lK3UgWs3yBcHibGIgIx7IBuW7whmv
mJsi2vswbbCaR9tIEv0qlrJBYSI+nsXfDk8wyOjHCsyoD6cPxxQyPBh4GOMrtV3V
Xserp/FOY8Y5yp2erbrbKiE5NvmBBXnltD+ShHN82fqq+KiSRDif+SJGTbvwedJi
iTdP1w+QsZqRBd1tdgmpSvF4WdJjIyzAbFNlXtn3inVRlZDCt6smtlT4/w2rygeJ
xOSTWz0Sxd89Zd8SGNd22WDr/3M3r7QjGeGHXtJHAzGe/83erLyV/YF0GzUtoR/7
NtBjjSQiZr88EOAlibt3hAMJIkcgxyb2iLy7C8NTpIooAB0UKZ5aNwn5n15XI3cc
PB0BM8AKJ7EoQrL7yKcgCZeaalh8lTRcQuy2fIBhU0i8EAh0W6EgtKhup1hlzsi9
5iEEwYtzZHBCtUt97z+oN26tc0U+R/atIC+kDmpPvnAfT+W8fjES/x1thpQbi+5x
3iNnrCad+TK16C8ZIadTvylVvN855TcZmBaIKf11NMloRiwRBujsaPjFyUABYG32
he7GhvA81QbOD3vjJCWLMqU+dtCuro6I66RMVBQcm8Q=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EzmzxCjWY9PkX/diE+zEs9dJcPwrEucFhDuX5m0zNgezts3lF9Posso9VMlN0+JY
TA8AUzCn701Db50o8sbzoLaQYg3i146pwWUKL9TeLRHR0ztJa8DSklELQESuwy3n
qn5XufhEzZo6MF0IquZ88VgSa4DXd5tGTIkseIP+2KnuIP2RXUGYmNZflopol3Op
eK2+tfybssuYN7wxaLWTHBFSXTKsiLC/sX7d47qUPo4poTZpx071u/Cts3o9CA3S
8iGAk+6mvoftO+AjEAmyTq4gVKaCOXEUxecsohIKYn2kbp+lXhRMu0WM3Xz/eaOB
DgPlRnP7pXJQ/EuaACx7Sw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4336 )
`pragma protect data_block
hHBYLdZ8zrg2VJaXHaL9ekyfwh3LGYXM3ezBVndVWHRFrZI+mN//lBAMQGZYVzhy
gTcz2ODf6ECNSWBwkk6tK0Ulms2Q1sExW3t1UJkpV/MJGoaNF0TZ0RShcafvBm8B
1qSe635S4EG2fa519QfV9iFKz/Y/Jvg90rgLfft96gqG8/WdyquRPfVkABXs3mey
Kbp8DF7mDBczK+FhGkB/uVOoWyl+NFET34wJ5/aT9Dl9hBgfRc92NGMzScePQknb
qOTJ9YVn3mOnuXQFT4sOTqv7WLT2mSUqXQz0OsrNhPCBGGIAogD+urCPX9tSOJTX
LCaibmBipeVOlHhdoasqqzpsMSJ1sk0KalK7LQXc1BWX+Byz1Xor20E3maRWyLn7
PVBJBRSZ8WIn1GzshCDRyXWzrw5x3iLpue2uhdxJRxT6IjbG8G3wYMKizT/ek3pv
4r/smKxyonVz/qdxUYYy9Rgh1didOnxTaK6hgPBct/3JIZsbHW+3hDRqWYs7RGyk
m2ucd8Yh5SskS5ZYMg6dZWzYZ+2Ah/NuhY9LC2DlZQ82J0AWpbijo/OLuH95pGMj
x4HetGpVR/AUIoEIJC3YZaqhy3Tbhgp55S5dbaKjU3urSImrqRZHifnQqFubQrvi
8HGaJayhYnNhyG4+kfv0ZGELiVrpsOroW+Sn1I8+o4RTRT19JXSK1Y36y1tFRehC
PFvBLqdQSyhIhM6oI+Zgp10pfNcqvFJ9vFDakzW4FbKnUsMPjl03jRwNIb8rRB7r
I8W2fLNLb+F3MdDJUxRhgp21IGHOFgFY1kbbmfzmwHDs26VCZKamWx8iTVnNLCQT
EzGgA+ef94xinY3FkzCjGuiGOtUeX/ZTlswQF1LebsBXSE5DU6+Z/8LWcpUjQr9I
gDhEO1hSugXM/I7AwkEw4ifGlnsAjtPxW8Szelw7RGCxJP5L2tqIuTG2RDQyOt0d
f/EpHGkG7SRtDTC0to0gMRaTOKXYNBdTF82TBK2UF/lOqZJqjJs8/4qJtLQbg0I6
3wqXCc8xBQI2X3kkqs6c9gxWQ4rd5dfLoSuHNe1XUYeas4knEfXUknibw6lvVZx1
PHLjoLJB2sXv9uJDCVAT25n7Ff74mjYc84lFhcpOSUXkCEluC4YdMfHoYqbSN5lM
hogtb3WSUPZl+f12w95zBiwI6nbCmZB+wQdr4vJXLwUfF0nBdSXkmrZniROybmt3
D7gZfIQfLVFBnZ1wA4c708Ag3Z1eA0pwWLTmwlB98p/qEZx22jVLY52TqPPSk2tb
uR70xDykS603bx+q/1SKg9c6GA3lbZXCr4sxRoDkt0RvZhfZ6ZP7+xpr1abwN/Yg
Oh54H4DIfaeAztYNEC5/wEsXaH/fyg1Vo373UhsQal8MEojWe0Oa2RofF0zYhrXR
P+yKDsTezzV+P/p3RbZwYj1JMYs1t7aRprw2npn5AyoijhhLz58mdZSsciSb+ZJH
Io6FOXD7s/lI5pTkW8VnJ9D/UlfgXnbfmK6j9C9MscieZxB0HL0fTk/89twpKrsM
Y0V/y8bMF3D+gmfQZE6+PVOHB0oIlHaq2gM3QtlTJPt5QGzuWMppY+mCVLCLkAdr
Zv/42ro/xRwJ4iy8oyXhiUXa5zVKQbNZT7CdHE45dMNMmExBnxx090i8qzzhkpjX
39/qzOux0VnuULqAfLnEhzitDmEQ+djZocyN8bq3bH3SYYCFfCk+3dsKxR96nOHi
xfibYLTTDipMq9vZbNqSgrCJxH36KOBbPpRDtK+omXn5oKdvDQaH6kiuWD8Z0Cmr
t7rmsSk8ei35oulUI06B6a/HWoV1V8dMYqkw4Vt+UqIbECjvkyjMv2H64Rxc533n
EjPxnnVbdXOzkYbWTmbyQOLHjAHLqJRSl1K4jJmhke9gPPVLgDwGEuMn+4OSgO63
VrnZ6vpPcT8oEdCOsStCj38o2oAIRRgglGBAwcFhP8lRqs2P5fCRi+5WGE0uTofC
W3UVDUV8KfQpsfPre24ne0K3SKdygZFonXF6INOOpH5qlq0S5+CIHIfuRw2M/8UL
yItV70LfQLmMTnd63eq8PoCWca43clS6hr2VvMdmMqPXkr2z2y9rICnKVGKC2/nM
9SIjOoI76JpBAxy3jvh1KAwtWkGDZIdkeMb+rReTNM3kWEsOuxUXGheJSvVjqhms
vLaU0YQVw+6qS3OgKujA9lFliYBBewcn528RaAhuhc+ExsJ9GhoCToHrJCi64PLh
XkPn65Q4VhxgX02IGqRywg+BCeU+82S0vz3iX37tlFrpRSo9O2S8FwApK0HJnCQ+
CNgt7A/HgYARkVmE7KjjPRuFsVeqOOT+HMb556QqUR/RRIMMHnmIKtS0x2P7Xkuo
auE9AzS/uvXNCr/PFeBCVrbZieIsScVv6OgPM5WUTUoZHihin+CEN2fqfhm6LJE2
LZuShwvN/KcRfqNanDIj/rRZw3ZWetmpS/gQsps5RKbyS3vQkF/CNBHURp9NLhVQ
CSZ/74BsTVirMhG7djzR9Me6fDY077IMZ3Dg03hKuhYL0pJSm0yy60R8XNhBH8KL
+1ZEuZUkddne6BrY4qFGuZjBVcIU8NG1EEy9h/s/7XjE+/EPza/ixr7tPhX50K+f
onTGhITdbQdhZGOcp3xRjezSvK9VqEinEsbKO0VKW6R4dC/hwNKP2YQYswolv00B
5tLOFD/90WX2/0GAGyOlQVvk4c0EHcBNpeGg2ExLKKYdy6HLMl0JuOGCbStVVdYr
s9vMF1DuxVjL8YHZFBRFksvia/iajVImDiXQFgnVOe5O/I48SKHU8CQRW4G2gFKy
gatVfH7eCBejsczJ00ZVkh9oyeBSZc8pPfrSxHlr+DitkV9P67XrT3qJMaUBp1Ka
a+nMMBOzFQJwXjJRM+o7hj3JhrxT5NH7MfMyKHLlZyh2LeDJ1FWqVKfyW37AwtP3
u44ve1W2qcJfxB1C3iz3OMc7tFnV6Xfhb00EXCcocyWMOYBCFP//7uNB8TWwvxCV
3E6KGR2wHhvGTBmBJ87twUEkDymHs14FAnHen61Fz2/T0N8vKoIfU06KCNsN6Gz4
xor7ORxzf2VAFQvuzY+GzxGsJ4XWA9r97TiOZ4Hkyj9u7SZrNSdWunocMm9zR3Wz
IbuYnMoInwT63EfBpenUqN2vPMuGPbVwoObkd6+WNJ70Dt+t6Xa1qIBRyPWAWX1P
QVvHdOsQydFG6JVy+xGIhu1giSX59F4HJicIhqyQbKUulp6Enyt73nBt7SI3NPBb
9/Gt6CklZpqQYgeP6RmdX5j/Zww3iAPjNemy+TYF2nXCQK9x+rZsb4qSVXlb9MKf
1tZ5WDqkllCjlUBendqVQ5If0qQKubAZWIcAkvPPlmQ2s0hR0twdliitKH5p5a2J
fPubHa11yKFO/p/IH8TKiaBrco2Sq6IW18QJNs+M8nU6wFu44S1d5SJPKwflUUqp
9LPe+2NFRRdO51HDoC5TMa7y5XdUtC/8UPPYnZladifEZNRsWqaM9XiJ9fIMQEy8
d+drv6PGL25vIxUSbudN9hBw1k/W9eXC07s7mD/+5bntP9oHsV4LQmFaOCW3aXgc
jWdjV13xJI6T0LWpkz84ZvuBEt0PKe+6pluvf2H5ENxg4MU0HfDzr9BOimWhcotl
1VRdC0dTp1EW0kYWaI0ZV4mUc1BIfbJXDQYp+mV4Fl++ycgpg/iOmMgD6ZCBSF2z
10V36qUlo8/xjhZO3byOD2CtO/cXTKqdxuJUGqOzrGY2XdMDybTU11KoB1vbpBIL
wSfUz8/KGOhiCVtsfXILJp0YG/DtZFKIoxEoBMoQs2lVhlW0WugOTDj4VLk7pN9a
MV0al+EjKq7NSMpUO/wiB7jkEOi0XDdkGKpQZQaW2bXfEq2AESWvhs3pSc0uytjP
AdzdZRBtasv495qdNEC2gd/A1B66aOmtUsg3khT4qJajtqp6y9ZVeYveXnAEVIBw
p53IJdHfTYW9Ar7XQQMBgiekEbho5hkqS1PsHE+NgV7CjIlF/W2N91BykTtngwjG
B31Elb3GfI/UqM0zuTXZtyku1vuFvW4ukH/zkhnF4K3WK2JiwepSlHVTXI1eOA3K
dzx84utLFZKVnCRNdI9JcfyeBKwnMtNb7kQ39Zvdng3iVd/y8NEBcm1Z6LbuQDOO
mLPOXxuBpEcLWlG/nW4FGUWitYZOqRZdvcBtB1tnS/vecW8k0C+oOc3eXZ3NdvRB
XWeA153V2OYr6GXigSIvsmL7M3YOeG9esFwfGe2iFvzUbO1UOyNPN55F70GI2o3s
fNqfRfKHtfIHz68f9qOlMjswZokuMbAF6mrnedfy2x771+N1xojAejqlr/zC2l6q
rT61OoeYrKzSMRkxujg7WREBp1cONGUnAWOuXR3VyJ+KNbtnxMgNqpZLntnW6bZo
Q/6spXQTpSmr+Fs571EUaON/H+h9Hdl9VEGnHZTMBLDVVg0zTvXlNkpr5vCNS8Vk
7lbPW5wtUGvxeozbEKmOX2NObvUGCD/wko8XPeYqkIXZ0R+RBTrYia7wX0uvvsJx
TCaOoPzTkUrXsaOcakTmyIfI2kscxYdN5RN6CjNbyR63KmOMpzXAbG03fggetdaD
4A7bULZ7vfjxSij0DeYzlPJkps9Dd4KveT7mnfBj8zNmSHJPpR8r3hA4g4itkaVk
p1HBtPtWn11mSu9Z3yWQ9bQ+uoMqPMIsqGYjrjuU1ZQforNFNXBwfZV1eVXlJ8t+
8hARTGAhDI4SwmT2A/jAwL/pop9+OJlqkfnhY6tOFRQG/iMGKxfQUzGjFLYIr7Jx
s4WRGFhxqddHijER6QcYybbaGclkx7H0Dekkl39FnvDzLBDBNS7JfTIr2ekPIR9k
a7OJaNvCPn7xl1DTInAf2APNOg3s8hUU/qo4s1+Lj07UmWNsswLelPhuKmxl4S5N
N72U6qmhhVuCOV4Ci7pipROwxbJNPHxTY+wtgPVG4A9aT910ANGOP/jUP1vfZyuk
H9nu/tY9VN//NEW/U+FcnIM1wAhrQppeM8cthRJkUD4O9FiqXi0dFQSm6KoQJp+e
T4EJ7FEPKaOh9PuJq3xD/d76NYXJXvKI7dPNNRHI5CmGAER4ue/5OdicBChtTEEv
aQn+NmfLnl7RsDgdilLGEfPCpmHoaUz1b2g9V5vWrqVtr57vSV9MViBPw7/PBkO8
3lJCjCHMFQbRhpDNaDj2keWBLQkiTn6sJvYOS38og+JxRuKF7wyJVWidNduORfAr
/sZDaYlpWyKt+Gj9YblJ8R4/bs9ZYS/5ks21S9eJE6gFQe3rwo/MDriT1+fwO87f
QiN6iUkwfkjRdASh/LPyQILXb9Fen8f7AczI4k1C+WV6x4aoPHREslk5yxrYxIx/
VeyBtFhYcSiG/WXEjoOfVGnFBWTBOmXw5Ue9IQKDFz8qLEbLH6LxMr/ModhZ+JUH
Q3pCh+iC+RREL75aJr+rvVquERv8gBr8cQZ8MvtnOx3f0uz2VsQ1c8drqkjNArfA
GVMF32IO53yq/3yStJGyhkhJ6qvsTmTnuMuMqI63B1aNn5+wajH2SeLtSR2lzglq
oaKQx3td9G3GRsKmQY6kiRGJDxVkwAzDYkPRopk0SkuS09krsXvKY0EXICGx7XxX
sxLaQFur710wIqlgmcP2HqpUPkjB3k7GsBCzBou4sjLcR6u0iaVa/aMidx+A723G
2NdAaT3YbXvsbYbc6iTine0GjxFuyl/EAncM6TsjUqhcr9SkqGVwF/hpbYLoQKGV
yvdBsKlLbxk3Ci/2dK6tmw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
OJmKll0KOxHRb6kLzeR9YcybM0yutybZJBIw91s43rkNOwIAfYrlzw7dHUBpROVG
NmwGXAcWITaufdYQzmfRzWCBkdjns4Q3NumjRRFobM5JgHu1PwfcvnFtbtcQt7jU
b+JP8Rsb+TDX38ck66wIJ5Uh5XgWqH3SbDTqNXYT4nDfWZznnO7O85X+RpRqRpMr
uE/1C27DGv5BQ7y6xpmwp3qykLsDccSi69Cvz4iv8SuChxtO2xcQORHXJYI4bERh
WqlABf0R1pv/FMZdVRyCFEtegRi3RAEq1Xi26BbWf3JJLpdxTbudJE+h03iVrvXD
sPY2cuimdkiMzD/8GWAKIw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6560 )
`pragma protect data_block
iLEEdvOq0GizvTfuLz3niQRDwbTdWYjZ/hHdDgdP9niHCFdsfbWiJVbLlNg03IbZ
Ah/WeBjh1WslM3ywPEv5+XYcHlFkalXP9lnZ5L7E9clJYcF91L1DMDaysBE8ZMUX
hVVkt/qFgrMTgkYaMq1Wzt+qTUX6ndxa2DFVpvsZ91kXmq7t8XIEOYRx0Oh0mERG
x8zOJc/SaJkpMs4ivEmWcD4p0L/SZZ2H6BC429P/X4Cqomm8cFpN0aGWBGlZmHFS
ity6PihBiVcVHJsn+wYV+tov9iWh+MiBTUnvAMevcMMl51Ps2sO/xUwZjX2qU9bF
gTtWFLOB/+0yWwx3IaKTcT1m4Dd14UtddVcpmP0j/eMtrfhObNkB5xrAmo60/Kq9
JtoWPQFj9Z4TJ24p67H4zUgh2aUCF24WHsQgeYl41t2xNUqZcJyOR4hBsfD2QxDR
b8JfflnxkZH86k0V9sgZj/aw8K3eFnYZwxUZIr7WQGmeEmi9JDXJX1D4YjCE0u1k
JvAhGf2+3saLNjw5PXk/xba0dX+STHHLJouLidaDBf9k1LwCJnJDFlKMnodxh+rG
4eeov2Uqc97zL3MlLwdCPGUu+GYjcli5VC8RJh9M4t8zirjBmwlqcfevy5PqzkqZ
ceSLzBfJnmd0bLexvgFZ9DTZ78xlejGN9KwOw3PU0XX24KzujR+V1OWO/1RpBNBf
087E+j1c79OvWpHhZKT1C1iMm4tSgMH3IkD0fHSC7WSTMeVszfudmJgxmrz+lQbh
KMQ3Q4RfQycyupgtgQ3GXK+jVg7tYYTuLijpUch3reXF/mp2Fqoi2nIG9h7wZguL
4ikiR8UKgRQiWCbRKl7QfMd1uKVYaxrOXadgogBXIQehOYA4Xkmu6xIiLj4FNMAm
aIhI9wgICn0wyuONmcNYb8gbgCJH+B7ti+4wgEeAQmg6htd2xDVbNWsKIP7oBPAn
Uaj+/V4eMo6S1fvqYg238IxkUNg4W/QdOKUQfw2VoXn9ul0bmcURjT3MJ+9Rj8gB
JeN1KYIQSJMsbfCpCodT7SipEAspzSa649KujOJ+9gStljiDwDOz/Yy8YZN/omA/
XBzzm2ltxxgo7xfddyQn6RzkyahrrIuXdmhTHyRrsg7b8t/q4VN3VF2CyPwFH/vQ
Ine7tzd6Q9yl6G8KHER/S44wtr2OQSbLtcfX7uz6IAdsLmS9iRoLU3vl3U7m822y
9Bq3rtSPzWQYX2n0bvDl88s+3hoQoR9UOADIv00znqLrhLZd1gREciihnLV252fR
B9pIQJhm/3ByWxaV8gOydoxTy9lSccLEpMlsH7Cix/l9h70l7paHMRrZztsFm5sP
lHbMhAhfyTuO+LnzcbQhgE0qTnXpfQZlVBie4B/v6dCJ94ggZJagMknQj1yw5C7Z
lHfZTKNqbVx7dRJ/KF0pXxMlXQE1cGNW1p36U3u2CjqOZyZSMPpch9pbVxlxCHJD
T5tbcFQO5bgUaFUrHImrmxXVdg8Vrb6l+nOzYFf8cnvxv3aIMhFc5C+QTGB2F/69
H3yNy0HO3sziNUEkivCK2V4ekz+G3l+imF+j1swqRMVBMw46sL2If9wYLI9DL5cw
Zi58XhFc/S8WzS6qCILQ3tjzdtzpVzppJ03yt7VrK41GMaWLEfwM8B81p3v9LboK
gKytIS44oRABcg32AKGGf/rsQ2a/MyReY3jwrWOGaVwvxgRk5UrYh32oLvINB3He
JEZF/4djH/LhaLpK8A/GXbS8hyOg4kCr9bXH/dFaRSfAgmIUIfE6wGGwI470+syV
9twEuOhJN8UENivg6ioNKR8BwiM/MPDlMD0gTZfF8wefWXxioyVQCy1m4HKc3vNJ
UZlqF0ccD2otI+710tKtMywjZThNDbolvvpk2oAqGubnh5k/1gUsfuZ+G9ikb7k1
p8wlSbsfbZ44SEoV7ix5I1fS45b9ko0ex6bqwn/AlxZwftoHNX6eLqYuvnGU8c7X
YnnsqQa80cbnqn0KSPy8YGaai2fvicAtVYiHRwBSIE6F0+reIrzlbtcrK8MXvkEy
PHTLI5fNaBicNvUUWcoMKhO2cxSzj9PPdvQqL/efOQsMaX1qLWM0n21rS2gFWAH0
0N/FHauDjfNNz55FCmUc6s7JIVwcXqkLgPLA1Am/lQGr27BWsqQ7h1HakuV8HW0c
MAkdzNiNtbpEXcKHVqe91Cjbj6tF2DCEqOSz1le4nYGybY79hYw/GdAOi94gZL3Q
RC5POz3E85bV7zOwfYfX2iYka10LEU3+eOhf69IcDqC5SCkCrLqpG0oGQiEovpm5
enBSOSqOIw27X3yhjWQhg1porwjHaPVHigWlmMRVVE3XPNxFREgAxD28TKFjK4qb
OnJf7SqjBoK+Zx7/LRyxEOd+UULUv5iYeCJHKuQ7EbrKAb5/87JTz3OAZ7O/pQa3
nKsn1FaAwbnMpy09q9OS/fnYL0a30KMqM7Fuq2YCpS1+UhV4ioLPtV9WIrr8RAym
HccJ7S3oN/CcByYXpfLAD0TbLg3azjyvL7SGWyJ1pgz0D6vHae0iAXAxB1dfcb42
ytHjxBs97SbkTAOkJmiyx+GMhgqUUw6udUqV4MN/XuWYUYuvbS1brU8zl+1KdqZR
XMbPG2gaYZL6wlWz2BeEyyaBkZ7p7pkz8gKafSktgCyOPpaugfRpUOolg7AxUm3U
schvyrLVrEkV30FONd7XrCRS2+cWcHqQLuNrDREC6gsuk18rXLR/yI/mIfRBU2Wv
t/2zW/vSO8Pbnndb+ksd+3T18Y6RlfaEi8iS0C5K8tIWESEp4rrLn5BPW/5GBOj5
9C6qrQq1L7rFU6si6oHZyzogbZu8wSl6RrJJETE+TwheYIVZLiuQ5MA0Gemo3UHl
GlhbDbgF1u6wc78iVULU6b2PYzmk4m5DoiM9V6GS4u0y8hV2XTaimksjvz1M5KD9
Cw2MhE7HakM0nepk5UYVqwzH3sU+X1DukNSRiL6tnjuwqIxLEHege0STSbTu6iJY
Poaf/Rpuv1K9c+4B29/GR0e05jBmiNOCN7yeglYz2/rlpSSdcOT9CSQfSTCWDO9w
wLDOpIaHpoTsxvN153xNNnDzt6nV/6JiDLdTU5eIjSVQVe6Nj5HilkUVz2rLR3I1
DGVXsyirU4QNsFiYiqhcESRAFA976jvrDDmmb57K0LuA/cMjLztJ4+kYfc/FTJwu
7h88zavNzIoYG2iIYfLEBcbL/+nQn8W2cUrmPn7ync80N1yy3bAgnDIrFe7SGTRV
/8e4pkCWt/e7mdNCe1qz16VMW211bsjSiB/NgH5Cp2UClvT/eutzuubr0qBDRwAf
sG3fH9vZiTWWpzZhM0L1AIcP7JF2Tf7YqPtx9HydIbNphqG2bTSnvW4+wKXUNkD/
iv34fynZXpoKvS+AmY4krywBdYaWcrs4YYaj2gBE6ZwOmnuYENBatrxpz70pZYSm
3LzwvQjZTICtIGudYTEvnQGPL6gq5mizWJhIh0q/YDtmceYk5HSh627r3ffpLgm+
wcTXFEAbn81qeQDmsGruTyMStVvHg2bFDYjczpVnfMi1hISAKqjnNVqITeFmTIJ3
3zlXQohTzT4RSTqeeAB/EbR5sn7usLp6l1eBh25SYIF0oXMrp6tRNLN0FL4T2IQO
mzu5k5UB4p9dufB1PWtCRO0rCWUp932w8z7vUtyjubGowHG1js3Gl3dQfWr5yH0f
1rNaEE6bsStVLDqoMHrqF4mZptVHx6Dd4Tk7BLKbTr5hs7m2yInIJ72ex2T6ilAc
XgJyYmZTRr7DQpcbWAFdQeUUdhrWaxMqwgSjOWlsCAX4AMkr+PwK565fwlPFcM8R
1A4d8KOHrBRoW8rmmULlVw1CMtPiIRujX6yilCFiRjr/j5puAbiMOXT+EMClIx7/
TLDzwfKEFl7U0eZP/a42aKEBa7+O5yrY4DfIRMZkwG0rd95Qw1YVQfAmv39L+Z0F
Bvd/2SPfMU1A+YrhGDwua4qpXM/CZejgEMS5dRRUBRf1S+wSzD+T7QRsqI2kL1IH
/KagWa66oWajsJMWM8K1MtFDmHUkKD9itzv7FxZTOQEWIbYPFGVQArXfXbvDt1m1
r9n2K9i7TbIMCArwiGdfT3NsWu7Uc9SQTWLv//WPECmxrhIY7NIW7VihmjZdHdqU
8GRIxM9Z/AnEOqf2NaJWZpDxBUgMVRwpwkouMjqfZTWtCTjykawPyi+qOzXWX2t7
vkB/Mf89nbgxCreyzBYmM3ODx+XwZUWq0aSnQwFIXRaL/fQK99dhiInLNq6Wdfpa
93U4qnd8jql7QgtdIONPOwLj/yckPLek7DFI5/PhuoMZ8x3Km+jj3zn6DFuA4Vp6
DABgFcNnQSN63qjqo83Zd+79CSjKTAMuSB8PfaE6BlQgP55R59w89n3AmIkhxqAO
0T2n9+IJrVF9A3pWJKFOuP6TfwsBSQYz7PTFXjrRZrnWTIdBor299vim6RqCoZ3L
ox0fPdS+o77laUj3iV8Ohsshq4LcfZH1aIFzw3YSE3YwyOSn4owhcUHkM+MFO4St
0A2MvMqqRRLNpgmtfQJCSx9rfinxnogzCIQRRif9Hh+WXvZ/1FeP/2nBetZbHh16
6he1ApsCL+F0YLIgdraOEskXQT3HpDH04FRYO1Kc3PfrtniZrqgCi5OUc3CCZ7ev
n3EWjh9fPYzKDnUNy6mrh4XQqU1GowzRCRW8rIbxKT6EKu3s3yDzzmk28ibhIlyd
+AELVX37GCUmpTB77Gi+EVUNm1iTYC876hwFbMlLBgqOO/6yAjJfR/NhizFMRlQK
qM4BQJW6/n8iiChw4nIGN/EtJkvcjrC39iW72H8Tt/Ff4KfQZL/dOzR1M4cTQHUw
8i+1eBYSlbSOYOslqZ6SPbFG4dQP6lKCXVQ2zAu/8ltStwAUT/vzVByvuMYtG4cf
XlD5o1Wetmtok5VZZVJcKoYfVsEbUBaNew1InluZC4ckJvbZI53A7NQBheXDCdyn
Zf/Qa9eZQx3vt9jqW2meRGLG7ZAWpHdEeJYD5tXC+2bsWEq9v87oWlQ8dmCalDaZ
dkuS1RO6ihKKtcoA2Ow+oRjpPExhjoIjerjtAn+8CuFPsJsn1tiTlx3uz7Zq3iCU
xbO/VsAyNlgKnSBInZu0Dl5SvgDLb17unFuhDDK4ZTl7fXSWxS/wIudTkXU4NDWi
p0EhdP2i8T7+WxQn/vhrzJs19l8yQ6TENXrmb+ejH66lYeQE8CzOQL0CdbGsXDjQ
Z6bmnlAjevcKxa2rdky9ZSeqh8OtNwMIEZIhhvW19hj35dGHWjGozv5CbxkKbDZA
NySbA5X02Fav2gLJvc3YuSuj0FMxS7+doT9pUGpS1A8SadtVrD4vqEfCfIGkY+id
vg5Ppv2A2ui0ri5nER/rXU8JXCvBFnTEJVm9Hqs8Z5Guqzq0MgMfHQyQDGbuTO2d
1fviRcBBREyPs008KIhgr7HBPZMZ2qZY8I4cs7Uze19ayAxvi/exSGH98yruI+Bx
TzI8A5PzHSCgw+aLPiM0FjLuvqU9D8qjcIWdPbNFNZc4xwACRfUMSnoOo1imSp/w
9VRFeGdfu/6jVTfu37pT26JElMvyGiGqOsvGF2cHRIZiCMv+3IZtebwD+yJGHXDf
Ez+EYOGUsGAZrTOGqnwJQFl1mOHUVn5AwqQSmYzvpv9tXyXbNcs38bInKllU2i08
6iaPDv5nPw2f2RTbIlTaiUs1FWS46Pn0DFrsRdmm6ni2n4tDDfLnz2STi2cPn3bv
KgDRu0UqqYRKqgArMc3kKpEkGYWndt/3R07sQrhZ01ExGi7ISuEomREvhSV9/oWs
VpPyVMPtXx23XuSQZ2rnLfzYF38rtlFRhJhzGBUcNhlL+Ag/7MEhNXezlMADaarT
G7cApRLpuMDCWRAg8H1eggymJ38HD/T66lu0PClt5YN+4RK48eCgQLsiwnXRetcv
1WkS+W7+6xMlHTSJRPh1tav98FxTcZTlqcO8apMSbVXJSht1hioylmG3TsnhpX4F
8AXHNPIsjlE43PqkRqO+E208nRYItkOa0nGMlVPM4ZwLRZE1Bzk9GmbSFTS0E0Xt
xBOvN7J8Xacihw5QKb8DQQd6oAfs6KxsIzltfCf3KHVU8SdR8gANvPwBhhH0WNih
47geTQBcQ+zKE+PNeouaOeoq7DLZFGduBi1YPlLAwjw3Wn1xlqHJX6EPWzCNWg8h
NFU96EwaYdQ113EaJRU5fF78BU/Fs0AzE7W4Zh3+CyTn2E3H9tjXtdMLZNrWDeVb
Cxfi0wi1NV8IvZO9RWbuYMn5EMtY5uOumsOOSZEKCMlSweCjKiEDRFZ5WBG9RI4P
XI5YJ960AyU8lal5zXBSWmioj2/0wxb6fJiLsrQs14M0J1u0c6dt7YOorugJxp6f
Mwq6cRoONjxjgf0pHFmxgl8Im2a4sOPP6KpwXVdvXpvERz7fIf76KrT8foDp2N6m
7sSvNIdcroEMbrVwJucfX87888PdFozngFxdDysRo9HMTO1/hP4jr/X+XS30tcOy
sahmjuF9a0bYe1jQIDxXp00cPiS62y+uebofP+IHjkM9kWIob6gKDd4nuJgDVV+w
No3IKpDg/DbaQ6cXT2zJjEK4lQXoSJZvk7y2d9UZgnLo+8pARLRmiPTIkC98Cay5
L2ioBjb0txKvc7GdnyDJo5gQdjvniUh7HqLoJuIAxsdQjvLzbeQZQBm484Onz4hu
TvC0jxAj9HyAdzOiPOVmu7wIkCJpYx6K/pP/RRHUEDJWvKgTKM3yzh/flTSgFEvN
+q94M7j7mv58dJcTBDTBErz1bBhRGDzqBJ5frzVt28x7IeyIZxLTVIS5UMlpvGw8
1uvXynbAOdNzRA5M0Uj3ZbpN8/hBOWArmlNDm1jmkCCLyD0mswgXdL/3CvlwVM+b
9/IlHMs9rfeUJAHHc5fuj7Y15cUsXM+OHgg9/6nAN3WXscDq4vOzAwZ/BhCvn8E4
k/ZQZBcHyowoJRaF1jQvDgSVZIZMnjd9bnnwx6/LD0MoKMCWmNe7aJVYAEwiJCMl
CgDEV7MvawGcZstrhgfWYc+pXLkHXn5+lX2FHz6i68bgYQoUPPnoIKhp62WFuPDd
TlxtfKLp9oB3UWNCdz+y2PN0oajv+5/tLQHi0zdQHa9CDrfazzgUGEh8f93Lnwy3
HEFoWtgbEUj1lbINHPRjD6Fe3t5+COmSwJA+sdmIkqhAn72uXkqpMdZbiG+AW5/0
CbqskxZZhSbdc7GorBbj35VnxFjKcLX9PwCnxBiGkEsrxuRaN1HvZbjHHViPThXs
mMNvKVaZYPi+fW5lEdPnKtrm0lV71+sx9SOTwz7Z0oDF8eaixecUgizPVSshe1WR
e6pSGFMGl0aRQo9qKkcmGwBVKkEDGetfGyA0a3TkcJRETot9z/kQqoRZei/DsnDz
V62YriOTkU0nXlh597XOXWnL88eWulMk1rgJ/QLr0Ag+8YmilyFsjbaY36Q/bnOk
Ci/GvXFPt7qV/NrZjCWbB54wQMLSbOhA0uQ8Vmr97OvkpyQyOYSjs4t8H+wqJafF
Onup9rkfc3VXQCuBTdHpk4KgW2z9y0Y3rDJpoIepMKmXyYi08cc7rgCfw98PjDMW
OLL+kKwUZ2Zmf3w2dAzwrS5kHs+LU5VQibQ21DiIjzdc8YjkiHy6JlAjQZgNtSDE
nshoDhhJwEjVDB2y1Cq8r95bAslS0AOKiqkz3Yd4/l2YcQm19UpeZHEE+3aGs7Ct
E8QczqbIc/rG6a8j/KvmukFkaq2oKS6PBMmgOHe60sf6j9dd8jPLkXKXUWsfiFYA
86JDs65pCALDFOlPQHO14kX31hY7piJyU0qR/YeQGL1hvQS24n7DjcZWJNtOSwFu
YIrAce9exGdP2aFgU7gnWXpGRwuyuiQ9K644CVgww0nV63zpMoC0wn+KPAgCbjj9
u95C7CdhWuxfvYLVUH3/bpvVagNRqP4KH9o6/HKDpbORx1iJfaESuzCZnSuZEHqN
FgOVawEgAlB0iFMTxQGX2aQQNyWO4JxmY4926cqxfX8K42PS6BQZiD3B9omsHUgw
tgdSDZjUSksP/IAN6Nis+UFn9zC+1hR1izolShpzEOkzRdvXynr8RgduxbtLTf+z
W3+VAjAtXZQhEx05VXJR/X2T9s1j+9+Z0d66TCfJpbfJkP9US+2wM6nOVG3+WV15
enMnbKCF/DpukJ/r6S6bF29qnWrOfH3xNp5cxG6Bf51NBPYPv4xiMpHW2HWUH/td
vECYuXHb/MIlv4fJYbzUZC8mId9J9uBjlQTaz4d9Nhzq2V2xm2A2pS5IT9WqRcuy
y752syVLjyTjt0fD+ZBTYo71eNXAXQtwTXVqCHFDWEaxpnfYsKE322vtlIHgxIiL
+884YkwDbwxABE1psliPP1qOzbsmyyh9VANaJ7Qk2GDWbaVeXPcP2FklFYQeq3PC
aCKHsi3OtWks/N1H3d0vnz6sOtn/KpMdSK8Ek7WFpML7rhmAVAVTxZIY8Iqx4Jqb
BpNQOBvPaE/Sob48Yc40F0eIj9/Z4kz+puwdR0vR/qAuCcHsifdbd/tZZholUcF8
1d/Skr6is4BHhSmUsV60ElSFAjsdTi6aadHARYl2RBeCVxnMdpAQuv86fZUTCPK/
e5DmrJnSm8ARXBKekbawe9U4wXhAu/FjtP2YpcJaptnLig5Hj4PZGqlqfAzhlgM8
mEq/tF6iI6fLtcQdeY4bQoKh6LH0aqjKUExMYYvISxo=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
CuNOITGoSgxg9llbY18NNJFNeE0yP+3ubX0ZNIr6yD3jSy3Lv6yQVwVpWecv35NR
nvMr0RGoyrTnu4v+1vNyk5Q3c0TuorGk/yuUsg4ZAHC6zZZUv93RFmuMUVgXnKE4
3wfQqo9bLLSMOU/SFBPOgIf1OnyHLladU1LLfkRahIpJpORSWGjDLx4VZYkVjelj
t/lLok8/w9TQ50LsO+bvuHCpgkuBByd1uQDVgfJnYq0OAhQQT2Wo6eGhtkEJFmFr
Hvhw5Qj1QLZBItE872z8+iG3vJT6MQckbHkDwO2on9YuVuhQBNFd4wvkixIblcG9
kYi4qxmvUthWA/lGdwqmiQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8928 )
`pragma protect data_block
cMlHevBFxwK7es9HHMEyrF/OKG3WfsdyICAoWE3XtRB+YfNfVzcllrPUwpCOm0kQ
cnU66FgpwEZAxe0mngu0qRo/C3tTTNOatjktcASr0j4pL99UXFW28jZZVJOq075l
ARlryxUXYDKWUAyAYdQ+7IW6bSC4ovt8vjrhFY5rpQSDqxF68JDAVQKW8v+dwQu9
9sdSbQ54egXb39YA59hBuRl+K+KIgPnxlfzwMbZj+Pn7DUOycFLZXmr9AwFAkGt0
QdHeHArqyAKn9V9/OAwg8m6NNY5X42acZl/RLFMJLwtFy9TC3sq3FyJo/AsEU5Kh
XLLQx2bllvFWgyNq+tXVFSziVquJZPKWe5RkCXST1CkROlQ1Gi9j8YF74OkY8ahV
Peo3DUMI6CHuyJlavj0BHQ88Cy+Jwwq0Hz/Y5OsOO+XC499q/V3IQTJ9M5CGcbPq
7UT6Wrhk4xWvQer52E9Lq79C0OOLryB4ie3mHh4lCh+VoSc1QGLzMsfwenzkCFcN
X06upxc/tNJCYE6Pu9rUZxsLXy83+ie/jXUKiNVajcTpGVnQqOqnFjgBtRlTHFWJ
PdEqBfdPZceMQzQEV+X44LcmU8OwHQgx4ZdUQgk0PtnfLhUXcx86Dy20Z9Bo/a2r
f05+Qwn6hJBQhasiSz6R9BdMx8qDmNx8VCN3bKudXpz85HP8te9P3gngh2PSUs0f
OU5KWMcw3mONgZHAxqR0GahNCcZzhOmTsbPEYm265ddzb7YvqvA/82zTfyiqQeir
WsL1R5J0uWj0MZ2uyRIUYcqkjG0yUfJ+NGs9iwAg4/UKVJLYQFb7P+9fhWGFGcrI
FeVDtGsKLs9qS1WoZQiCCMJ42DRKlg/aSHgui/L9G7z4GzDiL7+oD1PxiTLdEgdP
+TxRjdMS5WhXZnQhlqURKDybg0TCx1oGG13aBBF1POVZggNt6coxlS0OcO8dOg9B
HOgABXZoBle2qoz819eh1hoCNe71CH5xe1ZENOKLw4mL76cd6X2Xsi4knem3YzWc
4wV1MJtIk0jlhwNjF6/MOST5YAjWmrzndGhbZjOA2ZG9jWHRhnJcEnesbCOG30vy
LwN/3HdS7f0ppa+DYvrmy+7LkVBlGFhUR1I0n1orf1W4KOF9pvqo471t2hcJOIKN
3QiSVU45LCbzzqUdiUPiMB6mxvd5VMSPiiEUiwLTJcon/h04fMGXCigxiOPm+Kt5
Hf3vC9gA6+xXvZRVOn1B0JP0/VtHwT7i8Yj1TbugiDrjSCib6FkOH/UsZ9R0+3jk
ppNT/khasm5UiXFANHQwjETCXbjMqYUafgY9qwZWWU52K782TmfBuggOcJaFhKU2
EKuzm45YD8NI27Bkf6zbEaj+BBR3BG2L6VXD3NMWY17BBeCWTCV19bLgXaNSbceK
YE57dVhhPQC16g1cdGs6dtpQyK+kf6qNXt2Ud5zrjzCVAaq6spc8XHvkSeP4TdPv
z9uMl1Bhit2jEwJAPdhRka2eogC8+oTV1m1auP/Ye9ep13juMRBzlCoxaZ23QvX3
KYaxN5JkEYnQMtZIKe3WZcmDZHVyexG1scBzAE+61Tu9UqvGjZju3NrMiYT8fzEQ
1XbRZyJUaMOCzNQlZuCuKu4pKp99rS1VQY14+H3Xzm2ehvSLSiIiwMOoxKX4rZ/l
yy8O2N4rB8pG/Cd3/w1poK9IijUwC9eUsuyIpSBKBVB4IhcbqzEej77JuQrfc0vo
M7x46/wMIQNlj2h8lTIjOO49R79flWc8TTFNb9BlNcFX/FAIMSO5/DWHT+mDfZqe
D4utX7Tfnj/EbOP1kGSL3T7JNlYvjUq1hCmTdouGgqMfRPWDLzbk5O0NQm/4xKe0
qXUUO1JpyI0zVZdym8GVD9tO3DVVd9T3tJYipTVVa/8DQ7nGdAONbGfA3w7GhVQ6
MGlawNTJDFl/tHZQColQpTGo2dpOKYTWHRjh69UrRta7n/5vE0ayZoxCYta7KUno
hjIlx/Y5AVlyGhxQRLPbcoCToYpddj5o7xQGSaZB5/Hsray8f5i2C4EC9qiD67ze
5Ft8q/x72WUNKewZhYvI7hd+bgsFp8Uxg9As0ZHtkVSuilUj/ZKo4Dwk7i1niwz7
3etJ7KDlVW91dzyxpkhELqGYDolQcV2jRZADBs7ux5DHz6uxs2SC8XHFSFVCE3Sm
klKZWKW9f4WFwFsG+KI7luaJzUZD270qdf53WFWI3Ugr20+RLQOiqx7vQ6j3Fgav
jdFm17V+h23sNjM4lb1KCata5jlwSfixTgCZu6ACJbB0zsmWiM+r4C7tMEeZf1yN
7+XGp+QsWiFTk1YvKPm4br+8aE82ctmIWP/BeNDCo0iG796hUc03iXKi2tirV9Ra
oGFE9a6w23EGOxIXpzNcuORY86irAQZ94lCv59sTWf3dcXDO/lfqtnv0cM8rOyAI
B+QE7Xs3HoQldbqhXfv78RYYj5BQFTC1OMU108GGEwu/GaWZKHf+nJzTDkmMzNhV
75uw2lC4qvHadefOIt9i79jci9gAmI928JU8Gf+V+3PJwF6JO5F61dwoqx1f0F7M
japXPeIWorR5IOgEhDY9aE+P6sF4fOZNe13zgIB5WOQTY239JZm2JOnVdgHP1gNL
xfEHpNpGhFeKguALHC5x33MHNnGm/V/lOz8JNnKow7UBkeiUSoVOcZ6oyEdC9pSw
AzuvLbe0K3Kn+9olAYaQxGzg+1OFZC3dWsRQQcVuijF5e6rsNu4hgXiBWwAGomL/
UhqVrCM8gXnN+pyKdoNjXYQRBjWNoxQuGZEDr9pgg7JZWX3jTopeRokm+Kr6M3oh
qoRYan3Bfo+yjQOtVI0RnpMaVqo60FQaY/Lr9Og41sgUdHiHfWDQQUVAjwtP3iE4
TUdD/d+n0dyH7JcfM+fwGCrcZiowfBYe3J9JVyOQpaR5uwmhk8nexJftzGMWYMje
D6se/DyGeEiYNWTCCeBw2QJbxfYqxyEtjwiV0VqDBtvYmBL2JF3ncXuKIXuR9/SJ
UBHiz4J6I2jzEKUP/dhwb+qiL3MJ0q6DfgjUjeWO8bB5XA2Cs04XGOcf7wX+HDSQ
+9GDIt1NU0uEk2Lp6717VlpEf32rbqm46nlEiEqjlwfM0LtfyCLj/kM9EMTvHhBL
nP4DcPIyLAXCOQOiirC2iQyym2BUDdi5k4LOzCNfKKUXrnMxdpd+tSSpXNl2OOv9
Gqjbe4Zt+a7s0muar3TJTfgPYsmlyVVSDr9DiIZl1FsCGFo6vjy0FFIApCDPzFWO
JNY1IX+pKLarj2oDavtE3gFd1i/a7GayrCu0dBKz6tOi66Wz4GXqKGA+i6QSxWnh
FvW+xCt0WZDTJP7le1SdMVGRU7ZUo4v2kPeXIhif6Ai9JLu87rVTXuxaZm+7Yf5r
uXfJIDKa1vibeZOAfSSz9RaYeXwL6RDwGDtPj/2wxoX/S0hB1qCQ23wrclKTw/bs
PbQXLHWI9oy3Gqct1cW5Z4wDyqX1QrHPBqT4+Z0z0P5GXmEh+//SZbYC9zvh3B4e
MVF2s7N0QQEmPBLJXETSQAwiPNYDo+g3x3I7kDvPjvi2HG0Uo2ZN/wIAmuoum5No
UcEJNrwXQ50U6OI40K+8/qZUZ1p8oMKJDZ+Xfo29mrTzFB/qDMjDzDI3d3hmMY6m
4iGdLxcvmVdd2lQPCf3+Cs5iiODhxzq6ttZKslZHfE9MzQoE6JiV/5JKrx6JQeuJ
EvsHdFtQkjOFRF5vuk3fKPcvD19fmbj+uofLZ7dEa4XOm78O+UUzET4bedpgbOy+
LhVkL8gk+OVmFFDmA8FvYO7fXEQk77KvVhsnhR8SkMGd2yudcLG5tsvMfQ72MR4T
6iVG4vzvhZlugKmWdCmEY2bvLwvBzj3JHHgusw7SSKkhiJlELECohT0nGrOCGXFk
ypeQVqLcxXEBataYN0tq69RIkGJ5Q3wgJtFZyFAYcVlTsUxmLeb06mesOusWnWfh
X2sJElRB88clMY0pfkynq9jZAQBDEDM3ZtBR/3ZUh7VxicPyvcbN9ozxLtk7Rzin
SY7YKssWZFzG4vZ+AUzfxcWyoiLYl4gZ+u3mb9+Rgvucv0zqJNuk/NtKctPzhAqz
CcGj/Leyqf5G5ILARPSLebw3C6xNCnClvz7MgFrZMLly9s9zzOYnsRlGxH6A324F
JAkWGJUSb5M0K31Df2zwGpSnHtw5epsDmeTtqHJXbyCe30SlQaJqDfBXgmFTxivw
eeyeSpRry4BWiTj1DUkvZ/u847HmzSw0D/Ha7H4BRTdTDd/jh6LiZg+8lrTnd25I
T5Icsz2K99xas9CU6geCgc49KEr5ggVYjBtOHhPasKsUlCjkuEsinftN9K2ExgGV
kArbXuwwf2crWUNtWYJSWkrrGOLxDHc/imxVR6tWdaOJfE+1vHv+stoVhB6/ROZo
+86+UrKQ3++INfq7Efp/Fm+eYImV35GGAaamznL8ggZphvaKyvK9SrDcVzVqFf5h
n6EGgkLXVq3WYyI7vBa/KKtf8oAp1PZVUScyWZ6QHheOiPDckgV0yVWHpqITRx8t
SfhshmeMKztedET/Agn8MW2f7g4nCsnJ5ahLv+tJSWvq0zd6+81RtJPnRqUaamF4
fXZyfsoC9l3WA9LMiHVLLwloTWaKKYicUqTEHAALptEppVI6BiGVv87Obn00qZQA
m1P2TbaluQ4AXCyqfTe18mmXwKVYmsoEednGu2HeLO8vwsvkr0bYGXuUxIsXOeQi
YQFDseHQy1VfFh53gZOO87vi0g3oEwsT85jJswwCGOVCxz5zVVJpHbxjCOmIBKmM
FkDR/7w0YhqAlBO8F+TyCVuFHwe7MtWit6RwpYIFZ8zAt+gfY7IrxgpeLC/W9nD/
laBZJjDAWpdl2oJ0gD+0MsbmMkMao0wBj/1hbon8yx0NZ5niMuRQ6vH8JG8sLt/0
5uymKGEkXTbwAhT1YGLO/8tD1SWAnrcVGV68GhHOrUffNCDEr+GUo4DQnZexwnJ4
D9DYK7RsdOj0gZwsf9NhMLri5m80cOjtYxnnrRx5c06YtN337XfTjjp8chpD1z44
Q8TP+VvnqjtdJaU5X2gk55eELvH3uVz+R6YuuJK0zzbza+PMUBZcA5W/u048RQTz
MbbufdpOxNw1HKQ5AFp3OX9xZFW/ffUm609gaUeuMQS8K/XLI7B6MteyuOeVPQy8
WdCgozUdjTmOCdZm46QliaM+ym/Mm3LBulsPi3T9n8DVeyHzf00oSCnEMnRA5hyh
Y8gkGfPHpSaUuBdylJEvgP7O3KoeEofXgdTlx3IbZw4++kjD7jBRWkLqneUSLXRm
PNPTdtR2JvaTCAbr6v6ekAz5TFXW8m3Mpez4lwl9JQe7xk83T4JQNKtjlmu3LWq2
8NlZT84moTynfENJETEDNkH622nupmrtmgpckaSDLfo54jk4ZzzCBu6BlSZUxLbL
+/B/d593zv6d036iqaCtqo3s41HcUKNsG7m75Z8xAOdYbmfO4+cftRG86gTRAed7
GCyVt5Zn50AUXVbZG88kevTxZPwYnpsWGZDB0PWwL2UFTMrA1TMMZWIezjJ6tFso
xayuRSLbyubiy6YImguCpboqCbV1xfm1KIuBLdzNYQ8/7YeBeQFY6+lIIcK4t6q4
R3mdY33zzr/vBXe++c7eARNJtaMDnh73dY7HLfuZzbsSHRfpIso0uwuIi8rPp0dD
+3qpLtGu99DbG/Q+ahm0kw10O5TBi10FGiQTLFtnVVpxsJROhnlF4CqqxM/nLyVI
cZ36ccZo/de2Wz6H02KyPQ+e+jkw/JG+lFlNB0dKbFpyGCT/SDUa3ebbTe3Hd1KS
/k+1ABH3+4AOUVIBVSGLbjRD1+uWB2IXD6pxeaTA2mX2+AwUNpFUKB7yODojxxwr
TfAloK+uubpmSMbqtZr9ojb64447cqJW8kLb+x2d786f7TCBlOm7mVM808ymd/q8
Kf/jJK3hpAHfd1W07MsKqKDSxkIvY7inA9fm6UJVqwOBOMAWixjIP1y7gRwvEsi1
MmkKbERQfK4u5ehNTv1TZxB2RjrIsHgSoSfPkp+PiFinWXGWQo9NbFxj9iYC+fj9
458bHADq8shQcNMgz3wmYyd85uiTYQzkDReBMcXCpt5ZKfPqwpGrolMtb58Zdcng
wT0WMIxLZLR8dJx223ozvo8MMEIpl8ZJ9xeMpDEyK+FdDsilabiG7s/VO4h4+ELB
25WT+XEuAa013q4k9j0bLSav9gstje7QvIJl6CmkSpwAABJK/F4vetQhJlmrSVwo
1H+G8ddEuuJ2DdcJiaZO1U2gI+UQy/2HOwWpyxzYe9aYR2BKajkI+rGJfcaPF6kH
FxrJ0O/DHSPW7PFWXERSxbHe+qvLJJp5k2eQ3LwdyRGL0gZEVcBVpHDbRmnJcZqj
7sKs7DbDDHYPld88ic122vfKUYQ6PyPMRR13iCBpS+gwGE6eq9VTFSXll4dPdEqH
Y4KghSPTbJH3u4BdryceG9Qtiu5z9PTAoSUKz+PHkJqyydaHwMkmpeM+y+pHnQK5
ikMMnLXb/xkksXqlrqrP3lZzutlhYavyJg3BT9tRtx52pxoJ7hdbU4+ZtQPvGb8y
AzGl4STo+OnoApdinYi2k32QNunodpFo3w00RJE4Up71eJUtDOBKEM9Rd+QjN4rn
lzc2yZlpUm0jdtrN9ujEwQaW0qCPjNAJbt70/HIf81niLi2qljUwYPpEBwDpURJ3
BRsG/40SxzZK6Vril8cjJa0UAI7av06eA2AwKHEJR1HsUddD0AjJQj4/uYChqigr
895ym8cF0oh01qhTVu+mWFEq8Wdr2lVmuW5AjJp22D2BqYiD/jus92CRxTU2azEd
Z7N0RYCPRsmsUhX8g8XRvbYx/Lva/aixscKXud9Ee0pF8xMGPHxH50tBAHoLa3Xi
DZP63ceIz6ShGNmAaR4T3N66gDopvncnXIiIiR4Ny5W517IxBjYyNZVW1Zed/q1I
5sjaYnjqKVMOr7VKFUwBeJN7ORtEvUIcs/yG5CnTaIW22qMzBCC3ZggHMPAT2im/
UTBvbpQw8vmUg5IzW8cHKoKRPFPkeVY+TMEnjaoj4MOU0wa0KS0DIzwnkIP/Oa6K
gL/jhBI30b7154pstrYqUpNzh8d5O3pmraX32fUJlz7cllWJNa1W/jgGgPQRU6pL
XVpqofIKqYBLLV+rQ5Z+fhblG62GpQjKsyZPBJueMyp1jyhfscj5Ix5QlgkoVhrH
SlJBi2ir/NlgYi5SLvnv4RLGGXGBhTTxGuHNRZgzbD5MnRcwmA0O5Lgq7WapEAbu
0btAvSAisVYp3Zh8+Uvza14u/mNaMNnSWKLIZa0SERSTwOhtAKb+r50osD9RH28R
iQmn3chk6okZRDl7y4Wlw0g9KuoiympGscYX5AMaRqOPh7uNeDicZv1lp2jf3t0e
CZ7vEzKNZHxnGa5Nv3nCWrLIavSCMjw5CXS8RmwgNdiE5FVOp3ekngTOfwowN3Oq
TV5pLHhb7+ZWflKv5+IpzyqkzCab5d8yWYU6ysIPYQvLuI1i3j4GuZ2zn+msU9er
k6wYnzjHAqefHMsSwCF5+d3/mY6P2/zwIFVshEbjo7T3zjpVs30SCYbdXn8V0DZt
FZCOHPMFfwswyNsdmY4LRvInKlOBcFygn5lSry5kxHCUtbcMyPbgddEYB8A+svNA
qSxN0UT2QFlibg/KsY7QVr53n5QOzLlIyEqUh+Fnbje0rtMzKMp8KBhZXKiILW1U
H6vXpZKR12SRzRDK2ocdAfQ3UPphM+v9PIcDA/ZGXzWcAyI1zkbESChPSmut012R
0Ir8Fi744Zo6HfqGJedXggigJbLJXFS+WHuiWishbsFSd9sHrJSWtIUkCHeutn/R
kXhQcXaiv0PcLoD1Jr7oJJP74kGvG6md2Uia4QjkBLliikh2XQ06Q/ImiJMat8CE
3QHfVSw2EbYqLJaWFAP4PaB/a+cASFhwDqQ28FR1CKausRHAgOFaN5Dvus5lzJxp
jNPIt0Jjsqxs7jH81sFnE0Fh1Rg1de/e1TdxwLqLNhLwMGfW7miRaq9m0EftYUP6
DdplbWaxNOV0CW2SVvdvfN12gYcbvUVrZvGZtxyhB0UwkjDttGQ4iNwcnRdd3F0Y
SvxRVnekSpm5m/I9MiA6m+YjBXy79JR3IuGsTlIEp5qIQaR28rynmn+FYDzhsox/
eZ/cYC3HqZSg4GgfWrxOoyJHpQTwCp6YoUzu9OIeoghz8tEwYTlNgQsr1QHmjCLI
sUznbQhORg6lkdiVafPQsNN1+CKL1LOKa+ExFhP2TE07XSn710U++KHF5rDwgN+T
k6nS3S8PAVBZIdhintlDv8lyz/k6PZbiJ1SSkZAPHJ0qeT7XdS+CTgUAD+yALv/V
w/ANgEnWhxORg1//pRkGItz1vtR2OBsfxdhT0SA/NzctXf58jspXrTY+G+T3qPfg
bm6WDzSKpEyqKAiCictccaINg+Tb4nrdcMMUc6B6HVlGvwDL/TJEwn95erhKeb7X
LNWOazfUSG/l6bZ8toVL+o7DtynZr3ZCLH1Nkcq8W7JrxJzdaSaZGPCjwyoUyG6R
5+s5uieKTIeIFjnkacHdzfX/vaAynHNeMPfra2YHMiZ86Q9k+JDsCexpcfiSG0Rk
sZa9dcHJ9EdvZ/C71Rb9RXA8cAo+zd33w7Ms4Ak/LFieRvJdhlT3d12w+Gzucnys
qe5V3+wgbcKzctR77b9uR26tuOC1bKaaKc9qYJWssigcI6KukfjeMNcJ3T3QD7Es
6fyqDbblT91+xvE7z/dGy1cq7/Jb25LZlwR9USYc96qxpRi9LsyEHt/h8Fj93Tfw
it19/bYLkVei9KlVjVRz/Z63Y25jUtC+LvMq2UXs+U7goocVBpaapWK745rEHy1m
GlEOJirArz2ALgP/z+1rELD6dU5txxKjGgzoB0iQND3Ei35eRWdZ3/MRGVgoelaJ
XSoqjEr+6REmhWyZNWbkDIJJfA+zaU4HAlUSlGbBodftCcL27GcFrzOsBVR/xUye
EjTNvnwNzQ8eUUW5NqZd11cT6+KlbPV2Mev5RQvH6VX1Pdxmlvbn1hxoSRwKdoOG
pse8gxHgrfo2T3DXqbz8J9WpaHMfSfESVH7XivH78eyb2ghMnKwg5VhCI4nYty7E
sXPCSu1FlnNcPYxAs8nyj2vrBxBTOeseGwKpUtv+Hg4fy7q5yqp3db9sMOjntpmD
d4Boc4KQQP76FFBmAfyguX8WaQnPkKVmTeF3ZWJcdS24eLmwWivSryX2mYHeVrR9
xED4P8pKAlOISvFVZblfDmsqNPG4ay9hcLAx1Dq4rjZpnFeZUQncuXq4ZsXrhug3
3ut6e5a+F7wtQ54Jytvu7UHXA+FpNCEzw7GLVEYQFLfZ3aL3OdlCwURUQCrN6dl1
Vg7dh6GxZwXN1asQ4MmI2WneQtfGAfu8mVZRHJymYs+AFLrQTXDLtF3ze4fnCOPE
/MaZ8lb5X7wZ7aCYdjF0M9LdiPr2Y7Bu0Rl1vlykL2JWL9YOeAo0rBKmZXN9lMbq
0FFOOTPFeKQQ4aMGCDE7uDwKhpIzRep0GYaIoXUV175glEehbZWagC2PcmN7jHqk
4rKJL2d/g4VcyEGhyGuGRVETV1n/QY2ueL3CckIrFIploQZCvS6V9fCmRegL8Au8
/RG7HLicSAKExVhhhw6S7pD7nxcPdnrPq9jusFVkV1uCxZxVjDSPqtz8yz3qbIaS
uFwumjr0tTICiKem8xOq8rWutqSw0Va6SX2mrLOB7QYNcCee/H+CuG7nGDERrhp8
LHbaEtk3DCd7vYUdhB5SgZmoIdj7MRjODwgcYPgtGPwmAoQ8B/VpVNkh2/zSXYD5
9Sbv5xklKuYeFILOhWjC39YFcMZ4ReasbY1x5p03u8UEij7j2jY+kIhgqBKyWcT/
nh945pVf54+Ui+xBTDtkL/pSPUzWke+s9Qf+woa85jUyYsfNie753XTe5JYnF3m4
kSeNjlqdRj0RC5mkZb8iUHzVPCXynGuw5pi8C2IPoDGb58i31QIkzm1OMhw4w4gT
JNk+/0FXK9N2Qr7CGfUwR40fPEoGaZADRKmzh6NPmtA5u1eoxl5840kg1WSjxVpw
vnNWKOBG2blTzqbYkZIXxtro93fVSMFt8NDe4gUKOXkbQeMAd3hws5lfFuKn8+xU
1vOBGHskEThGHJeaPfbVoe/nulTyaLjU1kzuP3b8f8LJ2O7VNRzAQ3cW3UZtLwpm
dK+u44uqwUT64mwScHnrHky+zfvfwxxux++ccCykVFimF3FH+lIqV3agHTXHIlg5
/bM0Ilgp4NJjIXoNqeQgnDzwagaaHVwyp8tQWlC7pwoJw81inUqj6x7q9WPTRIzj
QOAWj8kQ9soZ9PQfoghqqSf9/G2JaQr1QQXEF0vod8Kau+2Yk/jy3PK5yS8Oh8sS
eVRIY/OeNum2GNmOLrQmIDEGNWX9hTrGlyWoe1nVBXedH3JfxrkpJhCgqgYiR3v8
SYWD868rXpecwpdsZ+g2SY5+rAf+Gus9ThNQuY3/Vre3Db6Tz6S+SMCifbt9Pv0H
c/syLJxw3sBnVmY+vxkDHgzbKFEh8xCdnoa0x8na/rKBOgGvjIw7OSsj2MZn+VjG
kPYJ2JrT+ItXalOPZYE/xTjH0GZbRd+3HuEPDmjqHAJikGHNhAuclu6QbgjAD1zk
0jv1o4A3r5GQQU3d/fDFxlVVFL2mPJztkwaCXweqTA4AzglMX42H5+siFBwH0Xw7
7OZf1WxplRWtVhG0FNvQlR8ksyyNj5ob6VbpDjmHPNPiQ8UhNwOgE6XVB5GdVSaS
w3M5d9Jbncd1ftaggMZDvJohXNM2m7fYRhyOuNEzzUEFI8WfmOt2HXabm7hHnDTi
c0LuQcw6js1EaTEV4zhpti36lDohaes52TyNFoLy4nYTn95rHnmxeQtVYmAyK6al
TN3mgLXKsanK7BM5QY7hpDgq56Vk+7qyMUwvBqpqvxaUol5q4I2HimpO+HmzRqd2
ruZktbGVZ1aJV6mqt5gPm+EHzoLOPAyVrFaDsQtAM/WR5lj2SY/PcrVBcAwz9Q3N
j1AGfGRde4b6ygd3YNFDWVfyBnlGHP2Px3TvodaCuoJc0ZAkhrfC2Go3ikAitIxV
er1oq4NkwbyHmfKgW4GIcSDytkH+ij5Hy8AgLn+sOVGUwIiGybV63C5mIdwQYBkd
ojxVvzOp2CMxj1j5GBY5IPLOhlwzIkmR3JaNQMohpAerhWsS2HtvF5Z/Y+TPRYPa
/gAQQRb4qx72VjpT/e3x6qsMDxN8qNYkn0BU9HUFjpW5qDD2oYjsM++j9L4rSNGo
WEt1JX1sxx2IN5VpQO3rSVm1wVOmW3NahBnjXx2wdxJtSYSRF/GzJfdaMPFEU5+W
3P/iUdA6twqsGS/aLI29hGnsJnh61A7yg+mn/vt/PzmPXBwLT1VOOnWZEEM74KhI
rmVY/zcMMCqpdTMzFPctlHXNyGtcBY6n657/V2kKTcUAtYnEfDWwv/KZ1h91B3FR
+hmNF2YAdXC237//AKvbH/5zv9C2aRC4M1JdtPhtKVSOP81NtM4cRwJTHLUYp/Ot
QNdfrBlj0RSTIoOo/f+KC+mVCVMnLv5ySJ/oy1rNlh2hpYGtCGVE/sECbOXpiIC7
+eRFxvOX7q90GnY403ZaQVbb53492FtyHne8uyBIrczwpzdRSegPKR1MlJdK+M5U
sOhIJzdsCdKsxGab8WoKP7yQN+RLcMr6wDS3evpLtQKi8vC2Gd1EZCuAc0syURat
fg9rdpnxvBW6AiHPzj75r38BquDUNJ4OjJr+97UoAYyrwmLoj+1YBNo6ZNyky8zZ
P3oWgYfDTGV7Mh8Dezo5GR3eVHFfg8HBrT1NzN5EFgbqnC1m9xfHid0YrHW8pUy/
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
F2CAQ6qaMzXC6ErrVcHkHqkNTI9SI5gpffxR7MXgFxiNoMTThz1sqA2sTdGQDHwy
PgkDsoSKuhS5uQd0r8Qli/kKSOe/r9FsJM8TMHWXk+xf3sFDClWjKJrLbET4ZKI7
VMwmg+TwcOk/NktWcqBPpcQWR5+vXKKwzEMh8JNQg9e1BOgldzBrFahOXJz7Jaxd
q0cy0fIBKtKTF1SvZVtEe8al2vvXo45Xj1XHE+ef9DDxxbSvVzCyZYxGZFflF8SU
0rZV6l3xQ6tXgYvHd/SoY/jkQ/omnkLMFUOvR6dNATD75g8ehYEV1f33v4ZH73US
WBpWVj/jOK6eRYD1mz+5cg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2912 )
`pragma protect data_block
DHekktwyczN4AsYeVZU4DgZALiwzwyNDRrUciM9CPObp8/EO720OAAPwpgRXK3e/
FtH2AFx2zousw+5mnW6dNoKqyUeTQGp8PtRHJQE7xt+P2Bb45mpW6uJNUIDw5R4N
vZ7C/0hPndlSDPNmCywLBkGK9+3I8CO2t2ohnZCbevLWQBbzRAzCjQl+7eNHskL/
ccSVcL3lFsT5tsuBbqY6S+RqYdpeporJzG6V+jCfc6qUTyr+LCnpI95N0L7+aDOM
KPWUOjy0++4uNmgzd6wUYGmS5MaeHGZd2dtZqmAjv7pIuG/ItAuyVvu0nNm23VVz
D1M7ZYwlTGfLmCpXKOs7NZ488nZzxnlLUh4Ngau2Eqo7uM1et1ZjG0O5GQdzD480
LxVmQD2ObP7zegwG/73jNY4127jBOZkKCGWslPJ/B0/coyGJhQAuhvdqnoH9xuD6
/BiWSTf6hpjK3gY73p23a6vaI2D2ZkX1Ag9ByYxrbiuanLRf9w6T/Vlu35VUfKGE
SsnfSc9oZU1iqA2gEgDJZRcyu57jMAc+jm+/mwZLsq/xP95vtrRb1RgPvOVchmGV
nsWUmKbgXHhBjj+aY+SUip7ZwzTexGQWg6hmv+HHWkE1mykMi4JvVznU5cSGHsT6
DGCd0uDdphngftzc0TGfJ0r+21SAlRVuipkkzJMCjtg2SPp7LpQXLNwJW21pGpzV
ehcB/FIeOgaqpdb+Ti2ZzX0bCzFnQD7rij04k4UPcoJP++DpQD8wUwwRkqQMPXQg
6jepZvfvGhli2suGe0jOWNGXbzDITDXYEU4Z+2YSKXj1UqA/nZeLkG63NyTIpDfO
+S+ysgy2Kl/JpGEP7znwgq2ElwHZgjpEZNl9tDqy/gUWAFStBQeGk7XaOLOPKNPP
PFI2/R1rB+tNnhgMJ7trZHTDQgGkuSDqQ8hcJ6GZkhHLvEyldsFtpU05RskdYIqw
w09Ae8rudlz5SaWbBV0ZM8vnKqA7sIKvMOfgSmcOYfCWPYoah0KEVjjximWMHdqo
0c4Pju0ET1Ou+88LLQ5lA5lwqkk6Ihypp4s6NqUtEscvZ2g+abSRKWIcHmaCUB8y
Osndl+o4os1q60R/QwNlU9wXbeORRVUcD3e/Utacaky9ye0L/RIIIWWQeP/D2vAL
Etv7AmYSdXrYhquxlo/LuNgv3ndwXlRB7vi3+OBoSYM0ea6e6h/IARylox8Ysep+
hQo4WmMlISuLv6FfsnwbxeWAQXXnEj6uq1vuh/pHvizK2FZr8T1whY2ZA3w3cZJu
CAIbg4xORdm0D4pmwDlw89qYxqCiyPf5UrqRkVE2UzycoIP6jGxiKqM94uv0n5uD
R6IzM3MGhe+EqlGgiElrn/hr+8DRocSyhyJ9YHuH4ssZ5O3EtKTeHUNE0+ugLha0
rUYPoGBkEYRpJaHUfB8RUwxo7BLUifzdhP2VT8lTDpk1NXtHQUb2h5L1AnEK7Xys
AgG0hGxgp0IAXH+BxmROT1byZvhBME74syjg6MbXVTMtZxHBMp8VsQAln9pyj4Pv
4PSSStxDS2QBgkWZ2B50HO4NztxQQYFv01sDjRwCC0Fxdox/VPxBqXltLfFqZy79
v7sAeJNpGKiSDaHZ+gv0NrvFS+WqyG6KWFqTh4uk1CwsAoGqxYAwIb4w9z+uu3gv
b5SELjMyrmYK9jCV5k588uY1XL+5n5zNlqP+fAgBHDPzwclj5JKLsmvihvgKYKlU
L1vJNdwcwb1FWtH9VPn+UGUqs+WCG5+DrJC/Ki276ZnCl0R4I4GNZxcbmvK1SvCg
VzGiikJKof7D8PzV7I9mhOs9OiC9vOLrozZxIlTeoZ2hoc/rHcHKBDIa8iMub9Ag
K7KTgBXwVVdbgTAJ1ezO4rzmpTCyJLSodUzp/Hd4sMgdFj0oDFF74Pu0+VrXU8m4
nANtU9pV1U4INY2AxgFIrhaIpJHIpdWSaK294z2B/05M/NI3ddgmlb0AE9X3lhSg
9l61adqq6cEAP0p3fI1RGZaY9awbW0kJmT6nUfkvE5L/hJqwvxzkJDtUaK/6WNWb
YLg01ehqpgaU+z6a2/21ALrSvpL+lD+WRgWotOq05pUwAdhPYv50f6BqLMgWl4DV
ElRWJJY6OjSSNroSUs+iFwadhNqqzGx+u2nHTNrue7+B2Ve0wzPMmA+XMsTW1fV4
nyuWfT9CMh31kjwrUu60GRlPXmhR9wC12FoOACUEcOSOd4jTygorfUysez/DfHnT
p6wLef/ghsMrFmAZUxdTNwSDIhHRxbuRx4wVCWfl7/hjno8BN1MxR3lVMvz8DvZ/
VkVV5HIAEHZY6pVtKm9BkerJKHzgetINAX6SyDxdKxgIdJHLBq7DnAehrkp1Moub
5EqkwgWmNP2v96Sg4frVNdxf7wbuItDRRtbmtg6qxgUD8jPjVBi1cU+RLBITWgAW
QOBRhX+6/53W6mxfiM7tHkOSo06+R+QyedyU5+pJtC23zpj6wxGR9eDoLjkPta/t
u+nRTMahbjG+/zAjJtPBYK/IvV6Pko9eThwCLUPB7/fqqVCa1BTReLuBTi+CFo/p
4tF3kTexAeGfPm/Ydfpz7IsTAIGjAKgg9L2D8wQFrHTGwg3QJPrO8NE3ImXZbYJD
shsWbrC4JvMoUDFcT6MtzF1TxfvyzwUK4i/shl/aPzgy645cshbUBO7UhZWY4oTT
UveGHyPXHd5IOifRH3vX+OdauPAt77sHcQ/WvFKSxPecxnh0uTFHfIvA368mnadT
uzjLozUMXnAumP/hF5uDqxS320OQigA9ufxWVBOcti/QQ5EAVMZ+fS3Rs2AqW3DF
SJVeBc6ANaD0TNRfD7vjBfo/99BgQlVMMlVntIG6ogd8BEOcFmrQ5PUjKrZJGm2o
/ZTrrk6XL2zv1wVje0b5YRgbBY4wv26p7PJqJrp9bbIieWc39NNq3wiA9g5PJc8s
ptOYHcG63QJ7RXQZoRSjV7B8fX6oE1Z+KMdS1iHdlZLF10cN+3yWZ+zdeANg0E9M
Sx9UXUEmoyOgxcSt5H8SJ71e30h4238+9mcMoCZdza1TGW36DlPvLbaNwrhwkOE/
e8w0QbgyoI9eVsB+Z4E1M+pfYurgWWcJGQ+HQ9tRg8ioMS43aR7J0G10P4emaGaX
oAw5n78SG/ChG0HASMl4zPV+1XmQuZXZXAVGFAVcLbSEZMOSKAZ/PrT3iRnit4rA
+sheCulOl8GGb5tVkPoUGdTYlLmH11BUJq4Cpg9wGCL8XZ8LTGl4N3m8f04eFyTu
S2xtre1+NXoTT8tPWxWHam63nWWtWjw2za4rP/OcJZ0jfiKn1YhMNju/fYRbfzHe
1RFQCUKjmJgS6d9BjDEikGjnHDljDj6YKLfQb+g6Rwk4YLoQRBW25S2qFgjbYfHq
SfHtTps8UepYhZBgma+V93i9aNO5qmvNNlf2YG8Mceg8r49rLVD2UCuR0jPW/BZo
mkUy+bWZ3cWlbDJtgu9gSA2H0ZdSXH+wXjZYeIKAu6PchSIZOVAyW5f32hPK6VEo
XhwvGor4TWx+MxA8kyXtLxQEVGx7G5c9E2cnL0YXL8320I/gu8+VR9SFl+jrrg3w
HrGZBqvF8U6QzaBZqWKnCLKtLabokPl5Oh/cxOHa3RlaqyEf0vMEYn6yFdr9xhyB
dt9enzDcT1vjMhd0bXEDbvsk/AATZu+MXNOWB4BP9f0qyhKBno4pdl+qcVUobDJB
rHSd+EOLM3Xxmop3NLXGJ1YFvXVar1lqGb1SRp6g+DS41vpjTUJgqcDWBiO9lgng
Z8RWZdnlDItWseLlX95alaZXzSn/dc++npZ2MnpPr7lPRxrYyaffzh8vz+jM117e
Ryp6ULFgC8gzGARfF3jbUenYMnWu/Q/cf58e6wBk2jY=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
mUy8fTXm1g+woPJrqJjFGVH13eW8377Ss2GqcfIyT1VHiR9Q8/yh1ijcuWsyk279
7X8VB8IUKHZCPJcDhZscydXYPZ+J2y8b7b7bsKEsipeiVhrX5LIbr2gzd6gq58Po
AehoiSkRj3eG2+X7/vVgwh75c+lIXay8BdB52Nv3vf+UobMdl4KZDQY7Vy16KgZu
Mlc7k8mKuOTQXKU0Ib6dhtl4UH8neCavtCQeQ+RfvvIu2kdZ9kQMRHGoXNVWpfqA
BQ2sFHQ1OjTmEsO4X5k9/PmB07CQ0lyGMcGfls6LDbQ4zn0xV3kVU4JxtS3rhVz+
t8crpW5J3eIYDUIjdLIvlA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8016 )
`pragma protect data_block
ygVUNJn405bx0Vm2wUZji8YsChlI0k2F4fEjcM5GzjZ9tiBzi4nQLtz87qhJEbx5
w9WVcUVfqlirnnlCKG7TZEU6p6c1tWO2ldL3n1cAhcCz7Lgi05BrxHK9xSHibFIQ
MsieO55KRyG6+l433N496cjo/iBtpV+edsVQOE9zyCy7BgLYHSOC2B0b/sesGIHn
t/0TIO+tSpxsVdwVS+qgPnogsgKJy/sm8RQtTLOl8xn7ey4hgCmXBXIWCgNW5m5/
I02bf3/nJ/GgWRfTaQ21733H/vBVDYbBIhc9fps6+LxDTdGl6xcomcuE+3KDG3ee
TBVbq5HF8kDaMzXeqdKcvdDDemAX7HFgRenZMFE9g7ndt4P1tZeOuxX/IObNCbsp
Kr3+vpwoqIppTEA9ifSNj0rQ+aF3wCen2Ywk+5dKc1yBvpsFflAwSHKAgGA3m/Go
LncYKlcNBeHs8SUXj/JmETqJEIBCra1uIOu5/Bm2Id20Pf1GN97q1NuMI96ncH4v
0sM5SXFdAzDW8/BHa27ZNyPylk01qGWq+TWYb3IDx0dLFBltifaMJBo3blU4gWmz
F3Wdaw5urf61QqC3mm4G/uWwMCsWDAy8WC3MQzaaZo4zSY7fkuTMsMzzHTc7U0eG
BviegFIyqQ70+YTTnEnFEhlXppuv3PzCa0fWmDaG6NFDggk4CI4OLNN4RN2/Vizr
gVs5wryj5GtO57fcghZ2FMgZe00Xb6Vol/k8OqnE3qQBRLz3QZizTgXA7SsYxwrC
S5l7koC73N3hAqfr8ckbkhunkMq9oVkwIE7uYIpIgahXYIafFHOn7C2qoMYi4qDG
yWHf+u8fB83gW2uapTlbqenjCVrHgJnBpIUCSMnrz+b9//QJEj6AQzoLHa2Fu1JW
cFeEcV6aLR4KxeFYa9ld8AN79fFXWHrE8k6ZmTsIrE6FizNbqqn5r5ZZebO0sTS2
6lVEu3kZTL0FZ7/RJn4CNYLNQ14UEZN6lNEL4O6dACAqQk7YvGrZVj+uXW6edkjf
NSvEeEaRZTmnSGUdXC83TAYgBm5iSdOGDytLCBqoff77nMkoL8FD1W4VjsNwhmPV
DEZljS3k7Lc5tlAiqN/ROszxMdj9SfEZsdyDiW6xmy919q00ADr+osyN/Mnvth8D
WkIigdTkZ8JpwgR/ea2OnvpkBKDhIbaR+bJGV8Omctrsb6s2XI6Wc4+DXoUgdfTZ
8cZnJ1tHrX7njndjaT8yF8AOeMADTi3YMe+vKlEji7KaJCcR5Ej/Y/rDbOvAcxEl
xfgtLo6ffIpAH3nuJvjo4SzSGIrldEkPF3dwHEVc8gGbF4h+BEVxLnPEMcEtM+JS
zHTI4gA8Tp+RTEKUQrFNfqjSbyylJjrKWl1Lm+x3jxtvnEAfrWVAEZ3Au7urH2JS
VwvyQgCO49aTFCIVjkzfbf8EdGzs/ESBpv8buIVwkrKqvANsDIGjSmLNrVw5Ibha
3pEIITHHxC+9fgwlQXW8B38xgumRYCKtFrPe3CTL+KDK7J8meuptqSidabrMMODV
eFDMBp2H7c+YPH90pLMFtqpoxkZNORgOByaHgZN5xAvJUjLldj9sP6Gf1xOVzULA
sUkLFSb4qOww7vHuWzVxtjEWe4VmowHMVD75yb93lTlXqMDtJPCodyQeIY8HS4Hc
3Zhpwwc1JSKxtxNokXJSaRA1kso4OCllDu3LIbbYGvloj4ljU29gyWmOTzXoMbab
RxIyaHGKoAvg8l1N7M4+Ch2b5rFjWWmCVZCAppe2FvgijZQuhdVdMEElBpHlBkSa
pk+lupADsUx7O92bmCnaZoT6+hDpZscIwLAu6z53dN/p/VkRXyFuT078U0g3y+rA
UsF4tRbyp2+QmluvaZRMQfXKaIOeEP7S7xp9oOJ2KHcZ+vx8RiH4YBkwGu3kDXwr
rJQOKEFm4NcsKnpUwV0KdUHtlZc1uanguJImeEQBhg1VSEFJ3hTSQnSrRkC5gl0z
4vD1dQvpy8Nbo22p+G94/leySzKjJNPRCawlkJqOPr/hD/HU6VAqj/GXRyY6t8b1
5rY1TrA078Qji1Z6Aq2P6j96FAodTus+l6jHz8JNsI7Qnu27WEJ2veLFwFyHiba+
KVp3wxvMQvFMBFEMqcWoa02QuU+oYag62Zv1uY1vAA2LdtNZW3fzPEEbJTH6AwRl
96HfwgchytIJCxfxlUFHZrlOfQCki3GGLDcZ8aHj0U2THN5InfcYeI1vpP3g6UG+
BEngY1GfyPcxpDbivbuaK9zK3sB+lZ4ReUUQRRb4gldU56CHelgivoaILU0THgQq
NZvzoALE885gz5h842K11L1V2BPW0axs+02Ausoho7WiMFBM8Kaay5dv0nrV9Q7J
FzIQ6xdMquEf7oAY8on0j/q4pCiH3lYdPZNA89wAzwsAViULlVSzqj24sHbBuALR
H6fRJJJZwHvZU1viSZVdYiIORXrXZyZFpf/pSFnw8wC9T30iqalh5bfdqjvZ7E5W
NUfWcIkn2iGJsGnpPPvomI/JK8cxESERVIG58dDQjeYolDhXOFPPff5eMLgQcewh
sJCST3rIoh2Fa6XT3x7tzzHrYu/8AkrwgcOPoldsLG0MNagbZ6o896BCDOe8uT1O
tu56JqeN+oQrJW0TxRGrZyGx6vZYJulvhS5x+LOci2jLXIGUbkSJI71BQ3SodgP7
bWqzcY820+QG/K2y1flNO8/vw+/7ToMuKV0yX5vCIsb58tDxU/PtPZ1rh3aRXB6U
xFFKB8RefFawwkcKlo2Dgi5pbpzeAWBppKuHIuIxeEfc1QZ5mUlzkLtjsadNLy/E
8MraKsi/TCK3vhMgdicJ8UFxBwPPfTl+bw7gFLB9UiCcJuEhPTbYp58Gj1ngv1pK
d+D6upwtV3U5LnjldORFWepvZEC/a1gnTdOhIC2pM94R1NmJvluIYOOn6T0As3HS
5Kh7fMlKD2Z0Zyqt9WP2VcyrwDzr6s1aWE4rmjZpqGVvnyl8x+n/zBNfksRRQJAS
j0bGmDgXoEQQeOCIDraeHF4TBdFC5C25Q4HSbEKLOA6ogXAbCWL2Cs+iRlp+4/eb
UFnhjz+WrYynR3KRumI+lGZFJYN82GnZLetfb8VmL4emLNSxSBDh9QpuGtTLpLcf
wGyCh76lL2+aboeFNPz1leRFjVL4ZXAR9h/YkJ3xSHDvv7riImvpdAZavnCGHUDU
a44nxQ75LCKMXSZKV0Jibc2mGOEdNTaWjFReJwRf/kMXO8d1pALAGU8FvwojRTux
GmT4EQkF8W+fFDh8Nwxsj7xKpXYeocAcfMaChOifg9HOCkVspcXiZ3LwJzbt2GGE
K34yshQQxm2adwlv9bR3Qnqf0he5KD+lrzhzWUX2dHToISlYL0Z2NOo8lLg3i07K
3HWns721zZQ7J+pHWcvc6Ves0+Tr+khy2Yg8jjDmcrV12f6wlrqgxpTijq9WoLjQ
QnK8KkF3EPnOwVnkCms0avdqJKizALI8YchJ5XvTrXaRx9pzu0dO9nYh6qNf/kkf
UfZeL5R8UGxFwSJ7t50C1qZrhsMPvJ/fCVtflbf2ddFJ3iE9KSecgjib0ECUwwjt
AU+yE9RnfIRIZYwMVieiDnSulVVqvgZCFenMFdqQ5zg95E7ZLL/pbVEIDcDJWxFL
v51mbWdWp+wIvgW15rtmpPGHpbArFcfSjuDiMxikIfP0iOJVfJ11Wq9nwbySHoF9
nFVqGNGdV0YP4J81k9E4Nn7/2pc3yuK1zOJ0RBSeg3AQtMZhTiPr/HdtMSXs0Wit
LiMS2jzw+55hTK1q5QD9+qcalGPxaIaS/LJ+GW7NcbbV/gxxzD+GURUBkTtGlciE
GUKwlnQGxoupjgqsheKCaDHKbcyxcUBYrX3m819tsR+ArdSyr7SN8aVDJebSRgSu
0RbkZsFCvT250jqkJ9XB7LsaNNbfJdfsk1KzHW0YDPJDJ5Ujgk3sMlMOLFqKMPQs
+0kW/AGHNnxRFzY+SMI8l0ccFNvivNv2RGeNWXwhQVCv32i60YV4PwncFk2dDeyc
MLVUt6T9SYhJlAhBZ7sLeuKWbU3hgpfoG7YSW+JJO9IKUI6rlOESmhY/txmu3BQR
8AAEkEH0z9RzAzADxq9tBn689oBzM50zbsvOBvKiegiJF2u8Kc3RqfHg9ZycoQMF
4Z+4zl8yQ3FNVKkd33bcYPPUD/2kiLMgJQzakB977CU9EiqZ/O3mEGQT/LpOSPEP
1/LMRCHOTKIHSDeaZ5SaXDwnIVKGhtfT/wX/BcU9VyylOZCwV+8/FKGTZ0Od4dWZ
Rgl01NlUCO3HKmn7kHoc1TSbVeRMNwc/3cqfvRenOPL9VIK4hGUkZs+pYHmUZfbt
nEz9YJfSHCEEMl71YtZUjuDnAGMfd/CjE9BikxRNvchFA/NBMxQFobeuI0i+w59/
rISR8csyIdRW8r4N71NavvqAgwYoL91fSX57ChV9CjzWya32KO5S/tdPM/Lw4kYW
ymVQQLquibGAOvvuJBcVL/DbRXV8LaJjezqvD+LSftjGku6/oCrnYk+iMmHnls3n
KXBZPxJHGAlvgNcAArpsNrbELi3sks/cBLDTSrdiemUS++AaCdeAxTZ0P0vRVfji
Y/lWlmjvbmVkv5+QSe6dpQPIh4vl+y7noeXOpEEDef8TzdkdLhJm3gRUVVfK0pxC
6CUA5yFy+CEw6x4R/n3rPX7GalpXrmlElfR6+NxNbRKPJzzPhyIIYbAX90pwKW5o
i1u+XLgfC0hhUfAAP56aDb2nCeWG5EkiPFvNUdgBV0balWKIkgSYCQa8D5OqCGXJ
pbDdBHRCApoQqlHjkQexXGnpkxoWkfoMGYpQS7cQGIjZN29sg46Y5xTWzjx+Jd3z
sQ7/pHp+N0XEFKjJyq0zeYeiH4VjQNWmrOBjJCFWvWKqbnv5vjjKLcPweT9ZuYlm
TddXxH7zLD6AeRSGhREGQHfIXdnuBR+o2dh5tLR/haJYcGQ2zYzr2/hwvnlqOqsA
pYc+Ll4S6Rkb/TgRzu4emNxXjOIhMHb7yHmD5sFBm1rPfGnF4r5B+dbqduRXWufW
eaEAd7HdPNNgRcig4gxj8LU5PC05SxktKcrM2GxO6JLB8UgKtcYo2BoUHfye6FyS
rC5zEUByXogwOZdMQR0AaPqfA4SpNh2NeuspWtuZMYfwH52HQxsm+JsmgZO0bDrK
bnJEuZuzaKMgCKCK5bQHEwBmB8Es4tbH5z1gD2InG8hPuFGeM/4PzEOtQlkyl9zN
FSG4JuItxWI7RY1KKXl/9V1kvFkLm9Er7ybKP2YSFgDy/x6NeL8fdfs0mg0d+C1z
rgXaRBU/txkat6VlXZ8wadQ69KH7hS6tOLT6KsdA9xhZYeUkAIqe7LiRaQa/1xZ0
c2ZCz05heXnUeK7C7m6jw6bZ/L4v4+cZgwmXzVSKi2CCBgSxu3pqyn2lNbhwdTOn
GSzsTeYqasKjW2JqLzY3CCms4owY5aZKLqim6WhnuGaAs4wr61Ei+FnzfViBriS7
+0iLM+7WrI8YT7SUfEH62nBoAsMkmmY/4rV9VR0FhIbvu4/zepR1xsIGVWlfFx9s
axY11m6XUBXT1yZAberBeyLbEdVdGt0ViqUpy7eLWdtd8Q7v79BjHO+bMg8Y05ja
/V9IU8hFl69jFJ4YKPAm3r+46kwUBY+bkv+W5jSd/Mi2No7Qp+0I45XWDb2NdgBP
QDKnD887zMIcAQ59zQZysiVctrGJk6OozC3a1AXgklMOd/AnpYJa0dGcLxoAf44+
DU2JE9sJ9pcwgo2qs70SsMZphncfSJ4f61VeE1yYKeodti8C3PBVkpBM3kOR94Xg
862FfsmkYy4UGeDDW2+PUj5saGDM6841HdGPEj5e+hnZ/NpV8WLmaBz8KtzAgqAS
+L+zTJDw1sMVK9ryIwulfc9y28Wt5KYVeVz2JU8GBv/X2tSkhuPdm9AOZBr5rcf9
KviIIkWiP624Vj4cv5m6gPxjeSMTv5xP09bxiRSl6YPQh31r12PfLi2ktBV+yN6O
6l9ZRxBJkpmbmip1Ywpk8yuAp2jSMx/xBNPgXvLCfG1F6D5VGJHLMU8/324dCGcq
V5dzyLQ6exDnrNU2JwUwu105jSglMbUI3TcUJv8v7uhbHjSG3a+7705f1b2EJ6yx
AUa19FpDZnprL7W/axMczAOF4Gl2g4LyTrhQYyS2FTb26gBSk/qDdK60o7gVmP1J
lOWGtvajjUUbL9gGnevDo7/apk6TrcMDBGk0w/ogZpRJONyc1RnScCyb2lYu8Rbq
ajFTycDIJ6++jrXgBjSO4QYDROrJTLC9YtRKC8dITFBBNA7ddTvJkCMhndL1Wqdl
AgyucnFulFNzgL5DL+4d2ZIl2S4QTQ6qa2BlKjvnh7iOF+k/VuzeRKR2v2IW0Hhb
bKUpejSt08S347uhnaCghp4kDBReeARtqqyj6aeULTUjKZV94EFqlM7Mg9D60Sjg
4sSf+kp04M2FdyxpDwGiewwrx4Th1vTQWSvICvLUoNKkRlf1F2LuKUiIfer1T+2c
sCzOntAnj+VSZGxIAcs8vRE2yqIGz58N/in2UuJ1QW0m/J3pcIFmY8WdCjJmWzgD
qK+ChsbJlfDXj9Mavw/3U80GGNqMC9fsUwrGeXey8y5v/LcK2uE/Se29aKdePudN
lD4uKau7J0YSIBXj8jvSirdp2G+eBfgbHunxI6LuvSWAYZr4sCfmVMks5Vc5mvnx
jiWiywXruBfBC5UcxJo90ek0eEIfih0bHdy1mtq3jDf21cv5O/pw3M5QoXk5AAba
jo4jGvTstNfoQ5DRMO4XcwVj4WayCVDKCWnfSFQFf+oznPZ8XUHaBKIketfRbSne
1LpYV8KbgqzsaXC740EM1/RK3cOh35ROcYfoNYo03bajqiFtyh3pCltEBxXT43/+
NzL/bzHHJHm+41kTe8nofXIwrcSSDIqsu0lphAQW6/sOD0HzXhxIB8oK6WUrDoRr
DHnZLI+s9krWEj6eg6d86YVQv7fSeEWzpitxnRbLaCqFozTwqrYKqY3glYlwwgLl
VuQDfr1DMQPTGdul4GpdyjTYFK9i2MiS7NLWBE5+vcVeBKXeYNm1xjsXhDfwm+nK
ImanRKdhZ42AbocLelQNANesucvhccHM/p+XqaeI60yVtzvjq2GyPoHNRgngY+Sq
b8hIdOepYNrjIl6DcDiU6t5Sl/gAsbBDqqpQq5VlbGfC1UNclLuEPmbQSfHirglf
ar3FvPZmmrQbBsBnUN42j49S8Y/EiwuUvbvU7vtbbg4F2U6RwDGR3oEANYyody8y
K6JgdYTzrMKcTfMjkIpaqXi23fQDbOh81fhlO2jopFf+WsIay0G0HGq0PsQBMXpB
fOtQkkRnMmzcQZph+0WFF2jfP6iEUUTFyO5cxMDHlwQbm3nWm78fgzxeWUr0drBq
4YMRL3CwL+r0v8QB6q5CdDB/5hyZLvULyfAwfeBZ5lT4BX88U8DpDp6fHuwgRHmR
sDwIwjIOzUqyYbQ77DmLiLmw6XQan3CMVbRZZ+Nhwk/Y/KVOS23fiblTrSMumxRy
gIumRB8NIGqdxzFhSFv6zuug8+yhKEGO9Ub9MdEiN6Cro3ubhla8TYCMd3a4ET19
ygJdTEYXcd6uoGezQW/jpfdNazjSb5VpysQcRTfQm6qzZ77R/FP9vJzfrJBd6gV3
I7WxXWD53O4KEwDFbCt6uJS7Ie9bCos4RtSvZpcH1aEOpXgBdTAWx7ly//ZSdVtd
aFw3KWkiwSsCi7VOt0bsxki/Rh/MqC40cCsgAzqQ6RHpMLD8IlN6ePw58XjwABH0
zvcZTeO3ppPPCx0vBFqAYpHHeHwvJx0h9nzjbHeVAH0At1srxqTousxoyQR5KXWg
oC1pbhk1/XTKhDE0w8HcSH76IezZXk1cZZlEfz3CxR2sjhh9baUtLZid0qpOiVHI
bfZ7nHoZY8Z+/2WD3ONUM1LdVJQvhdcs/x8t7Wxjif/JALxU6nn+pQMTEWtcb7ut
oQFWrc7TRgzEeurEnaAXVGCknFo4otf2LhiN+pm+AVN5tVc7g5026ZWtAgFSP/4Q
y3rdsaS8pcd6MhY3YRtncD703fmswXSDMEuQTRjYHs5V8/ScXKmh+J9Ua/5E98pU
Cg/7eLbUS3R924zSu+7E8Nk6U6p0R2ESsg8IyEi2QoV1zCuoMp6IkUt2qqlgt3MH
b8yuT5O9K8NX90XaClX44+JCIWZUjUyEGr4Tbje/V/ua4ZWDzlsXgnmPJbFp2oZa
5bELc8pRd/NYvG1DFOakr/LsICGJtCYkNd6bG4BYnJnizVJPSG1A0jea/D+xwZYu
8tunaKvRygGxAqJW6to9uoyMMo8erv+xPkNCOP6meJ4A33YnltlrXnxTffErFNkf
GWH2KUz5ogrSAEo5Orxf+pFs2eFJQaQBcCuJXqeDhdXT9sYfybnuTQ+9+k/58SVW
2stFZdMmdyQiHbI6mCBOCikLv8PhPWG9eCUp7R1QiCNKIr1YkSrq86UXmEBIuElW
AqmHtaL4R3PnpzpbPulnghscBcaxHFeNtQVeGJOyR1XXeCx8LxvQEg+oBo7jomwB
W/UJZyJ17exCP0cI9fOQsuLI5UiMIabKhJODDwWLndKVHZjVsPYmGnEPxCLxUjpN
dMAifgeAK9jgObwRiGB36Yw24A31X6FsOqV9kdj4UJYd9XEJwOgtMXfXuB4SaVTq
e1WgKAV0NvVMW+kkMH1+t048NqTxe/E465KJoHH9MXc7cp/CKsaLBeG4S+ikGER8
7A06NvRHvnHOxc+fvCyi5BLKItqKeh4i42U4QyPX903MLt13jLVUqy8yEM83Pc6K
fyy5LaPaPgLXHY2j0+b84FUynrdwzK7BwgWzrNTft97W3Ie2h0jC/4IGfUhcXca+
yoInh5xljZEDDCjtx1vH7QtJWeT/PDbQUQVNYHEuhQ+I6AFbPZOdmnVGkI9vOhC9
675fDL7ARR7xoZ2t66IKbLmJKdPJwbvAzo9uHjS8Lhe6O5/dCDCp9vLP5wczyYTd
hU8RA5DK2BvWQCXfJLNFd5xcW9B5mdncHGc0LkMFnIKB/1Yx2Jn6oV+gxpNz5fP5
sHo6RPBqiY6QSB1LbmUrFoOywaFYlPtgl690rM6YvLmlI8gknRRp99vY0CwpivMJ
cBA0FbWFHTotzWBk2Y1CBjGm0pf7A/F77FimxKjEZbjWmYqMkcXRXodNjQijW2w1
QG8BmmR9RQnPSW2htEQNWT9MRCfQTG62NTGyJbG4/EiDLSamDO37ewt/68Z38RWL
GkPCJ68hDbQ+xaIr3z0KKrCo2B6pu1Lo4wc8phNUNRnWkkc9r9BBzjY6bBIr4IcT
bHO7w2MA/Jgy5Wk1tt+VEhLATcmWthqu/AjRrVFwyqaEeoqMkpNAXdJc6KXyO5Le
QqZZm5yxLibbuMkmmBxxES6AJQmvhgj5b1d+Iu4CuWyo45RDILOcxJii1bmbr1hj
x1bE+hArdqsR6vImk9Hkp6aJQzApM3berg1IoZHf88Sl6gYd49mOWtgr4bi9OK4m
3ON5z3y3rFK6htsPTAg5TEc+eMf14vs3l7DqPid/OBwyT1y+ZHc6fuQRW5M59b5C
n6joavf9y40qb2XmupZAMmJ6qGyvWBAghf4/26OwkOT6t8y2BDdhTdvEyiSw7hSV
sw4SLbtYyTscDJit+dXg78eQElzVF/kiphvAJCJH1/kwYz2djKEb0Xwxn2OxsqgJ
PGJXjXxXPidD8niLYUNetfWzpaqjajxNYwnsVPKmXMfeXSzXSMT7DNgvr+TOEMnd
qnCZplmIcXbQnbGWA9qxUxYQ9XflvkXZbQ7VB3a8riXhz17w9dph1sBiNv8VpBxM
5MS5Qy8yfhLKTlXs66YKa9/nVswAjSN7ejfs6E19ieoNipyQtVK/zMqBJHv94lFJ
Un/bA4JgdTNgB9iLVdnkGhkH6s1j0TNz+cpoH2YItEnvMUu9aYFu/Z4Y2anDheFJ
oeiOVU7JRLshH1IJPsmseljTQmWQ/6qpuPzE2I9Ab0F77EjwWJxPzNGakWDm2Ozd
pZev9Dq7SHAXLL6UM8/w7ryNZsQSRu/7trJUiy7UU5DOQVn+T5MXPxyDEb9NThzZ
G7vJF9ouNaD445HumbpAvppugGerAN0eW+KsOqrK6lRC6VKY0xbFQGbclPGfGg6/
JPrplggO5E/ML3QUWOqxejja4oQXN+6XJtUKzzgp91pKE1+KnYmlI/sm3ZGQoQBj
K9NWMCzXqyyePoNxlTPdm+5MGoISWNl83a8kiWfFrvvpjEhWPg316zzxI5r1KgZy
RYOTWA+r9AHGOgp5SatpwzCOlATEduGJZ5CPlKOyOS9BdXyt94JW10yjVIdMyG0x
pht1M2N44xQVqSymIRX/VanO5x2rX+v00+QuMYOP+AtJI9Oo0Nher4GOFu/7qnx6
a9BPoebqiSEvYnXm2tOxaJkFzbteBjnAuwE47yZM/f6HNOIywagsP1Peoglbhpru
cePD23KekrMTlBAU7IxdXKDn7SF4GyLeXMC6qckHA5VrWxdSZgOmrw2JtrsOdfNU
xg0HyJVdPd2WQJh6vRjtaxM9yglM/qg76Eubc/i6NP5M2otaiQ92qRFkznkV7sjs
OPpxniFUrVJD1+OQmNS8z68PyxVLsYT/Ta2oOK5MMlBdZjCvccaUUJJkRbt8oYz1
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cMmcPmWstrYpd7uGZ8GVHldh/7Mzv6QmjX4s7msnWlst4y8LHHDFd/er9HQcArou
mlLqXvSA2R7UsPhc39DVg72/97VgvbY/f0AruyIOC+PpX/rtdCG5tc0KmSvniFpG
n1rbCYG8y+1FJ2v6N+bfgCLn/gGp+mHZjqOlZIyDaa3mY3MGJNtbB9FfAO4ulFel
GMWRoptR610X4hdZI3K8jQYDmlur16daPkZxXI0PTLYy6JbxdG0EwgDk8bDwoSYo
16ipUDtPg+m3B6/aszGcSv80uiaEsxuXg1dYXDTovhdBKJTjzw8vfA4WVt2CC5e0
MiLf4pQ75cz/ap5apafzFQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5392 )
`pragma protect data_block
DDffiDQYlTfqtA/+ZywaMyYLQDosFXxAXWloTDWUPwMcbipvaKJwbMBR8yADduWv
OWJyC0u5+7rArabJEwmAj2U2/4osmYCOwTf12rFnSk4dU9if3UUyt5FBG/oAEnvy
2vJMX9aCO/cK0UhqlaeuyuDU8YxmxrZH1J3dF51MLD+rLrIwP7yjTK/n1NcTUf3G
YZNeHkKkhPuaYjRAMQcFkxt5XPdUkmR/k7UvpoZvO3SoW73NzZYv/3hq4dLs9fwa
g9LTLJpW6qPN8HWavyknfXIn8hkV+zWvT8zErBzuATyryjTcCDAJTerwEjucZARe
GCL1PvoaEdCjJ1oalXuGTUxtcLP1k1LqBo40VC7LqdGgTzULqLrmTd1v0JsnHt8G
BesGt8RBTGWBPfsTeRyzx+09RxZA4meQL+qoqYp+6LA+eFzzK8N8W+eQgQk+b2qZ
F5h9lNXZlF7plgfiZrD0H57Ys95s7JS8XgH28DicnZXHzEMc2OswwVoj3K0BDpU1
fRyE81JFk77DUrkHTry9IURZa7VDef/+mO1fT8kBFBO0MZDAO593qXCPHO4nc04Z
m4ZxgxcIixsY7zxIlOE3b4PVfFavD94deo13boIIuXKl9D9bK02Ghj/19Hz5KKA0
HLhn3Sgfy3myZAdWlnjbLdu6Il5FrCZPRo47M+ldfPv/7fmApuWBlmmysxhZ3fKI
jdqgCMPiuuZpDhp7NrW42wkSzz8qTdr5U7ttqprZjv2gCEng7P25RKe4leci68Lm
mljb+qtTsaF/sz9QHpey3DUux5hEcm4e5/fjgKhtqwd90zBk+pE4PvaLzgtC3eyF
+tsIQ2JXYF8TWR/ZSJ1FHmpOBifTMv47S6YPtto9EjJ6Vw9DnzkcLpc3BnPqed7z
NhvABr8tw4tpE+hrQw9PXLmiGso8USvzgwVg4BTqcbluVjW2XRjWXageXIhEHHoI
cWk+d46knOYF0wba576cLDjCuAFCpSVj9FsHBTbGqqPt/NGyt5kNQfNGQRyqzaLm
9lu+5tUFXGx1FaNhqm5ujn0VWfsMrjE5ulvjgVMljkMYeW79371M7I32A3b5RqRM
xyUA6pp+AJ+UrKDlaoQWA7cL62DSa+hcHac/nfcskRcRok2It8DrdML9UMF1Krvg
4wTuyfLgMOrjlCP885etyla0Rbiez1MQk1ZZog5vOT62KbelS0CM7rrHZjtRRhSM
73zECKHU0ubxV1plJS+s/W8DDa2/NYw8+e84XgVDurIkrF3Me7NiccmjXJOudjm0
W7cHMbkHP+lty/WJ+LKx9Q+m9fJ6dydnPPew2r+MBcSO7/XxwYTSq/6XxXuZa0C/
fJIGHTerywDvRilHu5jb4p/PwRe9bZ/g8IVEEltEq17Cmkj8Q3wzod4wH7ho/J+7
YEl239QumSn7AJNfghsKn4dQrfBWPLuwUx0FFxUe/NfY/n8PjixUVKlnA5pKY2aN
ij5bwY+79IRzNjmbCskkG8Cql7InvDaKgsRp1lmKta1EQA/aHNXXi7yzTIS5SAwr
6iMzyxuVdo1o37zuKGb14AMBwLO2Ko9TM6Csrrg2s/5nXYjBHGhpPiDVyl/vcRc7
JqR4pE2iZMj+ZMm8zDEzfjHqp/66+boTC47VMM/J2rwhZfU2QkY7x/t4TUN+SgU8
FKqBKctHEPnS7046dt3b7gmFbPdp3c+Y5DDJLDXycX6dU+AfzWwJaE6/2PpbUCv6
L/ZRy/4o+A7AjKJfBk5PrSKIwnO7DQosSbsqLmGNUCM5yFjzb+xBll+1hnFnOSQ3
G1epYx8/VWTeLSuyYwZSlw9htyfiNiLIRmAi62H4Csa2YqlmK/zjtEUPn78hNFwK
XIr8DoxSGPiN/qiLHevGZpK04uUlsuFv3vbxp4vOG3/7Ly9tukcORSIlnD8d34n7
tSAPs0hpT8npoiHFB+D6coC16KmiI76Lpun0DxceR1MuGT6NiZm4stiDfMEV7PeD
MCpfnu/vndBC0TJ5H+p6F3AqikPxE/e8iRkhdjXLGLQOOZbTQiUo8qqmH/P1xfif
WPGqZNQKeXDo72r1KnMu9pboL4vOXzKdEefbT2uJzwB0kbwyZSWXBC9SJgLcDsL0
4MmiN39V6B/MpLxf2MtNQyTqOHu6VwGaNG/4nNf+1/4U8veWhsh9IXHnVMZStMDO
wMpsqCX8Vga7++jTO9m4SCHGizLPFmBeqopMoHaZF31+pxyywS6K/24Jl5Z1Qs6h
hwMcd1v/9ZjRWQsSQTPrcAHcEZoM4R7jFf6Wx0Lk8QuLLnRlFXWzmARYWNCT1Eim
88aGpAAHr7q1gh5Ql8QUrIDIxGwY77R/BWvCsAiQ0hnaKWrcAouL7Vv3gf+KD4qE
3pbkwfp4zRNIO2TbUnbURCq9hRBUQg5+s7aYgJ40wyp0jt04xjZkWCkrMGshqpu+
wVP+kXhJjp2+AJtogO4YSgCo2mwQQDA3zhz3068hR/CmTgstVTPVHE73t9joXx/5
3VENesisEridHdAi56udafqowG0e3GFI5F2tuQhreVyLJbzVB0kOR0ADnvMlvlEd
A5yiLfst6OzT/fPSCgBTyId0tJW6+oCS3SFIk6gmwrzGHGilLX6kSvuwa/32H+TN
+Y2thXC45xWJtP+pUEXUqpVwyaJX8xb6qF1BVmq4WP3GNcKsMZhaQL4c9gCDQSQW
qJl0h+oGMFs0Tw/sSRToJO0rbve7GiLN34biwsYLMT/5FSumebIoJDt7z8cTIuUV
SGNWO+Hm6gG0g8KBFDa5xBVDUxguiXOBZRcIJAnLumGzBAtyFVeCgyIGvIvyWgA0
t6icQ/4tTuXqFRufpTQnqTmA0akNgADdMerBW8vCd0f0MPOUZQV+85moM/N57mrV
osmY851PCvLO2UrbHEoyC0YeJzKZdlgD4iy7EZ9AI0rvTr/mKp+7M4cJlp2cFg6L
sWbyN3WbvRHtVj/vwgsVljgmWndc3GnW2dt9lj51FTqT937dmQF3CiwrBvJKdZGH
A8Hzz2htOshhauiKsyvh9VwXwzmQNbMTrW2EWc8T0zpocAjjgAJ1FKMnZYipVLVn
PTiWmD5z6QQ0b7VtfhgMX/m40PcM765gQzKkhQEunNzZJz3rJWRFAxZBdQoNpM/O
fDW4oO3vc64a3sRfGk0Vhs4QTnmxDlgYqZLKJopsatWUvacTlV6j9It24gJgAZ8x
k/DGC9TA9US0fAjGsVVvmtB1blRmi5Uba1/xq6RLsGcFa6jk97EIdS64hweXNooq
Z8bXI0N2vo0AqaSuYxnp+i2+m0wjxdJv9KRV5R1/zFiXFu/0uo76W53iu/QseSgh
e9R9hOF2d5EMLMpjWLwbqShmjEDYKzndKmewlhysk4A2Uo7y6glt+OcoXEnVRaZ0
Vd9mLsysS1Y4mKhQwwBV8sMtlGPgdBaNRR1HVbkO/MroW+yx/+E2bYLsMxRzLri0
HSQNfw8CdqNUnvRCn+N0IU/Msx1nElkFZv9s+py0bOUgaXMxGOhQXS1hEYTg/bUS
u39kZYE26QyP9EomQ3mjwaFIQD4Y8hgYmcIbf04sBYvE5g2MdB82bAdx9Htj5DtS
9PRrSyzgsHgapzGhJ2L1EqnomP1Bake+l3Bwv6Dt2/OlhvWwheGoED7FKIcFihV/
77t9gmLSjchyDy+snb1EUVu/5SCNKXiESU7Mk6eWTfIlRATZUYLvlPqT4aCEbBFv
9drstVPNTx52f6xkco9zUkmQ0Qk+9pB95jArs0z79R2nb4E7nMMS3Aotx56VYD+2
wejBstlX078fQ2hEXPuoXxymBrLl4unO3BWoJ0lO5E/kx3gO1LXIGVhaYc0kbb/X
Ee1/bFt8ph9OkzioJdwESHvidMwbKtijTSUMgerrsbz4/tWbsC+KZ3FdkD9GpDf6
v754O2kWiiWJ057k+6Y/424uccH0cjzlpB0fQRlGV8ii50TgMNuaiOxcOaIS9ie1
DcifnueD5XdI33g+V6cwy8bnMCDdgdwEBZW2tTILDgnBeNO/yHnx5L5KqL0b6oh2
wyLIQhGu4ZXEqbFHLkdRzG4g8waR0YbwM8441hXuOFW7NYNwIQik0pYcBcaol2AD
mFQtJwYcbQozJ0ZdnPtlzwEkgDRvgpRLNGEerSN5+Lc8VHfQy7vf5SmVeA15yhPm
smZLAclqpsHnJKYS8I8y4GdT2X22vroR+2DmA+p4a2KR953fxIsf1YIl3yPEj61W
WS9EBOYiXbEBmpWskqC0n3uOb/f0Lo3b1LW5FiqzfKGuTqWDeRQOOYhzZ40Oc3+5
nUG5iJtlwV1opxQF0+FG7aRgy4s+pwO9con6qEPvEeJQi0njFsK8cTIONSTAwkWk
oADp+/AHXdrsdLs+V/E/y3duEUUx1FxEhcbfNpxFizb7AyCEzu9a3lyObUumJcaW
IBhI/P8u8YpMTB3LTmlaNyXRqpAVytjloS/rIJ5X+wj1KGapMWzowTI2lUtSdrwf
wxyNkIlOo5sXHj2zj1i4OpodtD2Yw61Pkw0KAkXhoLwfQyWYPQGB6KGaubL5d+Mt
fpcK8nVhpOrRyd+4Hs96w9qcYLRlS8G6VXYwYcCnkdzUL5GEIXfdfDgSKV0blfNg
7MUyH0yIS7BUZ7T7+ZRC39k2QS58OQLrLzXQnc7altnzss4X/Hyhz1e+Sedpj5Vt
qySZQUaqjibeikzGJv1amADCqZVqn/p2Baui9M576ChokFGK2HoSUy96lPNepT4a
l6BhhXOhUkgof+UHuh+btkvIs5VorS4c7qS0EPuNFu5g2Wahk8iJiP8KWtqghJtA
Y0PfgFxysN3QaNtPU0czr5wsisx3Ax4KeDPUD0VkwVmcmsJPxoOqT93fojA7Y8kZ
8isJMJFM3qtH5BR+St3FsofVYlPAkbHZP+uW8ugRCzNwg0K8YlR0DGoJC2sQG1n1
G9uHkDFaRVKvpYHXHmdSmBute1uwywu4nMQ6a+xFqGAYW3jl8zMNK3Uc8rAGV3lJ
ZBJi1N3dyI6gGcrR1uudTjg5hO8fWXNspKD3huay7bEntt2QUARdXNzB+TryV4E8
l2Wgcu1seTVqaMWojIwH/2qHhPB4UtlERjntzzKisqf4dhDLIX1aL6TfPQEJLsz9
wqJbGOWAsREUIO+5VuakLeelABq+m8VBLQDkzDq6IC5vBGN3MnsZVnt4+6MKifPS
BwPGfnTYHlqCYFqwnP+TMRL1U+JLRG9cCYhOoLIr+JPcyKeBVWfx9g1r8eOeMNIw
lJuSWoiCBSeaM8IU0xIfLyeU2PwCAAbxcYfUBPN1pl5pzfaKdM0XSek3k/rIzwMy
qr3DrsdE+oN8ZIN6Jhn1pUGSkkKX6/GPby7J0TEvkAqpKBCBWYZJAeSeeJPmwPBi
QqsEa0gqK+Pl+4TwPkcmJ8g9rIx1iX+RMCpAlGPVOr6/jG9o0e0oUyn8AaEJa8zD
CUcyRHmE0ONk9GLkWwqFO4i80bQToaNQKsjiEd4hdeBa5lveYuRpQmTrm/fyBrsj
rAdXaAtM2kzTIEa9Np0opvTfYOc5vIvN/NdXT32/PfhETff6NmKtdfTE5+mSAndV
1sZLxfF5lJkzLbXr6sjSTmaEbRse60z0vPDe+GdWt2xKY+213sVsFNlHBwd5S8L2
b0XWGc6EpAVfgO+SevPCDYDyrLFwfzVDMLUZFBAnOLDXWNm91vZihzcR8dYcT6ZV
gz312ENKQ69svEg5qhGR/yUGR28RT5WzYcMV2NolBTsX0FN8uObCw//9gaKk50wb
yZWx1ABIEON3zUXADihkI+lA7iYxPrC9ivrai1GIJEXSfMwLQ47fnkcfJcFbPs8E
tU10zRDwoOcw5kr70k4qXFqfqtiZm7cQ3giaWn9ua4Qxt1w+eODciJSQcL5a2CUz
WDl+fPJqmQ917M+HZP6ge2kpDKxjKZkK5IVQdBWLB+lyQx4Qn8mL8/LMG+XO2d2X
VpZqlZ9LkwdXxI4pW9beUaJ5W9hjOzxN3714Pb3/c4yuk9UHQrCFiiE5KR/4m1Ey
QnTEHbdZHUvYvPMgHrDtOGQ1hm8G9jVC/RNGQmxEs2CfAugpKOAAWLfku4/Ht0if
sc8n3i5i83h0JdXZyvlY2hdoRiKgP+jd33MSlyj8HfzkJ1U/LDwaXpspGNOUlC6j
PE6+KzuwMzrlGIJprMRPKEUaManucKcq3Bycoys9ShXSoIvk7HXRUJCMLDqD6tsF
fV2TDAy+pPgvCYbTVLD3q9tCVHkt3GGbdsD4aN9x73wlHFS+IBeEe82pDeGs1NdS
C2uXejfYUlobFojPZE0Mafse71FuP/G8oieccUSJwzsBGCKIEvou9nL4TPayiXRG
M5L+dtGYRq9HVeFBW60yljwBWH2IEh+QN1J5oNKd7ha5PtaSQxpDEIpUfa3ssASO
5/j5eJ5GrqNYD87Wj5SrcPCPVK69anVsXsTFQEi9bAphNP4/jKmSTI8eODErKKNT
FU5c1oIHLNUFQcE25EWzsKaZ7hN3Vo/o4zEJ3uYhJfEqA6zVqxQZcfD/+rqvp6nZ
8iTSBAMKf5ZHGDPuenbc9Isxh97ikTNGJinZR0tUzn7T3+NmEjKsyJoQTBWSbj3p
69LJaIpC7fIQ+YGVBKWQYGZyQw9pdgv3mUQdAZVP+ve9BqX0LTt5LOhNCjwCpQIf
MyOb3T8R0A25rKKBUR7qxFMQurK4R6FhuH82CME5NMcDfrKbj/CSWaVxUiLQC0zC
+mrp0G/DVC/2Cm98rfgLRPPpKiYdYD2l019NIKK7Km4zGAham9InRkDvKdp7MtnD
DwxLIs2dFT/wwe66qtai+6gO6cvJnQPw/ULFZISnCutJqZSoSjzF1CTSxZsgmhGa
UQhxtqjWQ3/ZHzAN0fBV/GKXHNE600rCC8NI1dXPhjXABOb4/3uemJ3uNpFtVmX0
OP0lsKv+BvI2vh99ZnUUYGPhum4BJarsPZZ/d4JdJLMp3WwanPsSOFGGqmdKzJNP
ZDB7h/cC49xSqMQPiSV13LfhUQinR8k2kk5nPL/yansOhfpGKF8Odo6E1SCenqVn
a/A0vqkIszsg/k+TljBziWSGZqbNUC7Kt7LnZfpkwMLWIcp+tqlVkLHSmlTwRhft
ZEVc0sjj2BIQRb9G3NJTHjSlxtc7Gz4SOxNhTip8yiQy8Sk0jxiCyha7hY5Vzodg
Au7DVSNasktRDQSFIPzwMA==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
kQ+pf9fMgMMqEzYzcnOnNxSgCOKflN1QMNi42j1O6bqXeIFCrv55Z2sgsobWdD4s
8YsSxFeyM6v5N6nyL4lBFXLxOv/b0b6GMbpbb2iU5e6HiLbSNkHw7sliRKYi+Nr9
CbWks65H593MhntwgjOQ1cIZIrnf5aVxNc6xAydeeUPi8AApQmtMndv2thDDp4G9
hVoilvDFjiIQ5GgFb94SQRTu5MAObxvi3r0kEyaPAcjsEcDd0u3l9qrht/rxf+eh
cfjPeC8o6/q9v8/ajWx2qp1LJSqfvkn5UBgmExeK/ZZBCfW7o1T5Sxnf9bzyO5V8
gQLgkf9Kl8DBf8L6nZKeaA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8864 )
`pragma protect data_block
AtR7TjVjBqdmhqA2u72SjCoBVrRO79aTuLC50QVbAjmMFIr277ewrjhc0l5Lcj/Q
OiEbYK1P9FkMB0TW6vkxQydwVLx2TgYulT771cUIZCCuZ4zJQV7NRNjTgz8eW5KM
d+wUrx9UiMjwM6s874eA0wbv+kWwv660tQygbmDJ+SXCdxIP8wZurUn8i8nHKIhk
SRSMK9t4dtCcM/scjF9Gm9R12Q3RK6LG2Grjscav0ktPvzNXvPsLVMclo2PR3YDi
6BDWOgnTOuf5hRy9EEofOBnYbDzd2VpvaOmkUIWFrnboAv+3tqQhEzh4B7wdspVA
gIW40xv3lUCYxie4PUPuNhRrDR/DQ7nrZw8fvWhE/AMqyhxrf+14bI2YxpfVKY/b
ndS2xMiFFj/cu+RnfcnMNo+xJ19N0m0iVtAIVEBavzgDaOIfaMQfx8Crr68E4qN1
OfL2X40ibTRZF4UciVMj+IMqLwiDK+jhl2W4o88y3zvpYgwvW5TJNrhuNiDUmKU0
wJQ/Jt3aS008ERMASxnNmd2VejFfB1C173nu37tj7oSlkk4dt95CWZfvaVpcehTZ
NB//MS2BAgY+2zwhJUqdOVHcfXfEqGEaMgJorAxVEnTlmEU9/ihxOLuSICiUM6q2
0z9J584J3+cufzx41AMwNyKb7YDHXMgBzz+rPCJGR6MlokUoySX1FF5pkBz3G947
ec1r4Cvq84G8MQqCqibVhVr/zB+Quty6HHvBpFrwhrb3R3J0+vaLBD1X2FrThXdJ
TY2UwOmielSgJoMUfRFKKEV6CB4I+yrbAWda7Db8c+9U+PqI6/F8RqYULMfztahI
JwtWHUK8bi95OPEI11eblUd3QuHZRxI6xquD3JPpgZWf9953SQ2++erMzl75N1NV
uiI4WrWINLcUFX3DRSUGLXpJLnTg70JdCRpjGrH4bqKtB8OePmsdsqsV7liDzR3b
TI5DLbyhG7D3U1QLcckTa2Km4BVOGqdW54I6dAMvA5Mh/bPOAwMLKgexxe/1hptc
6MnVwpi4azIqGIXnYj8P4K5t1Df5nHv33fvX9gzmHPnkv/wa832sZf7mQehNh5JO
JCExpa1Fc8C2xT8LgP4f2W15bmo69ZZdJryt0yN85i3rXNRAmpiV/EgobrCcgLSe
7EmYd0P5LlnuO1/o+cqwpHUHUnf9Ggc5yZAYeeeoQLtbSzfN6gfLA83jgunrSDrd
+z5r7+/PL8DHgN40cHqNGrhtUC7FSBbdP0ek6Oj+X86BJ/T4eEC+q52Yj6ODMAnz
R28/J6dT9g31lLVgh9m6mmMXjrnxJ2zA+wFuoOGKjd7m9bC1GduoG4TIz8rRG2Ev
5IfrC2g+EZyBwZyrYDbhZLdzqe4p11kricEyYAvOlZ2U1g/0NWPLwl01hApAwVVQ
5q/uOYLR69/E5NEvRdWU3CXaAWNFE7CoaOqo8YYz9NL6xI85avubEmVNV9HkTSkP
4DHeOw0fjO+HSGRq6VMlCOHX3Z69nqfCyo1OD48KGydeVmiIK/hz3ywYS39QUpgu
C6jsEerHlc7tQe+a2jAp6inBhZya12yJE8bMxfepLmYAIz8OeRoNMDckcLXWFqok
JbqEXAuWsEchQ7ElaY4SBxu65GMxj7Cn/O8YdB1xpCv//00jcQ+CACkxMPezPnpE
RJRYpi48B0qltQZeQ8mjRXSpuHfySFfPPHjHse5o0DmWYIooWCUF4V9z2/plZhAb
yD2FpoG/bqyPUlYKQJJTC+zzgb/WooipvuYdrbjsvrl8gaEKFvh67sNO58a7htf5
UMosgcmpML5IEInbq81DVOT/zpvLSt/YjQLlfpF4T5sGHSy3PbCdLEAS6xlaVKzG
qZeucirePEg4UjjF4A1KJcBBgQeB8N0NbSBkO/sHsVFDU3s/QDMf7wSBd9/61OMB
csUC6LEN71kWjId8IFztXG1ZD20i+7TkM/JsurceMawsOebHgyASYzbi0pSR/Ila
hK1FNybU5SF8FbA8ZgL/WTXC9TcgvKsREM6YB62WsCZvJnfUFR7mxuMiP2zOxD38
PhCdDtkZ0vnDI1NNHItupFnYWV6yPOl2xRydgfxWzLQxz+SbcUjW29GX/lH546yP
Te9UQ/TsBKbVioDbz3riKrHe0kYtxy77nT4X6BVYsZtuE1DaHcn19wk4C1Z4PzvQ
Asl8ETZQixtRoDL6eHstvp2HRIGvtScXtsA/QFTY4ol6r2158QSRfFfVd7vYJ129
P1U8CTXDSb0wDFRZKwbgSQennSjy5CDh0OYa6+ltq74NaNTcptbaOQDvQ+FGapIU
JJwI8TJidTiJgxH3MVzvhVoJMEfRFgCsiTP6pmDGxHoVIs6ydo35Hvk8J7pYXzdP
+0qh0d9dPk79JbaWOjZo4dMOmrOJiHJdtWt80jqUhWIusO0OTJDiAZav7WaR+b88
5p7uSK61EWXUSNQMfIhbz8z1uPZCOgBMOa4RpwmM/HUGfijjyYRnNhpwOAdeQcQN
bgVQgm1AiNlOq+8xPxOa0/MUtv9JWyAnvCqA0eNrEmCcdaYf8Jp3Ubv0Qd4QS5JX
sceXJXbLRBn1Iplt3RgfeA02a0EBAfsGpB1vPCCK8x2yCDrA8JSM8csInOiXHwKi
UaV+LBmR0A4CQ5GEnyoap6+/NSaKJPDuKtIb8gLYrWzeunktD4ZZOO3j1+aHP8pf
jNJ+N3DglS/K9ZI5idCmUJ08BSCB/nxMZQJeefgFbncp+Q2njUSltb3CfgGqldWs
6YEsX7BCR0BI2A4xpK2wQmuMvvL2bk8eIRdzRp7DQabBFJqKmWoIBfnYLD2agDvo
E+7rvJCWV8GQoienPPnp30YriAXB8CT3hFLUcuZGPaf7fh2P+BZZK1CPGhC0xhFR
4Tjho2DwIBHQzAuujVCwIy1Oo3+IYht4xqq3iVhUct9oKCC5/i4dkuT59aWICO6t
H5cb+BQtAeqEMtTgy+lPD3DiJtr8I3sk4wUmNRw7Q+RrkkjMHVyFJrhsnYyx5VEZ
oyn8id+hmDiiYZ/XyFUBOYW4c3vyTjHXZwst3QOY+C4Tu8aNZP0O2KflMG7KcJA6
k9ugqYNuqEe4lFwVB93ev4btwI0jWZQjIcPN7+7Dc9AYdXL6fIyv4z9oS/noGtMq
kdUCjWpaHku9iyiKvTiOewN4NcFStf7xLk3LuXGIVIN+sEgUodgxEhz6HGyOYtDL
7Sa3NZrVTVCGXsNG0LWBjZMc4hot/Hr6RxiTU+KhNaKH/wSJCuq9zeBKBtgzrr4B
1/3G/QF4b5dSmVWr6dwBqbe2hyvYSeXJNqVnFDa6Ml7QYHs169SOl0NHSQsI4YPi
cQZUqCX2g3FtD6MiSBPKnGp8lptBCBFg7l3KCoZPaj5VK04xipjKHUMLiC5BngXh
AFrHamFDIvxRBJR1yNRFyACVhBojJUqYhun26mkh1WQmNibyJ898u6TQxo340qPi
KW7uc1wo+rFLnRfbpxtmFMAxzgRa9TZIU3JxF/o4HKoIsvASJRw7VAJB9T3lyZaL
EbQBzm83XecZ92HuNpPcTW7NQ//pyaoRNbV3xWeBI4+R463FDYep8VWMHbKdy1u9
A+lpvJurdurWZ42fegbSEwKdHkWh9FeLrUm39MfSmnYij6fC9wTGPgG/T5tJ9/8Y
w3zAZB27XM14AoymAS9rbBpuwkEKEg7gO4jofeFpPcjY4jKVnNAxDY4q7MADT3yK
No0/C6RoHE9QHEy7Rn3+qB8DXSzo/ILxWBdZLUf8rN7UPS6jNfm+9zGGm7INFH9P
65bjFULthsM6qvgtkIXCoi35qiFwC8iVBDYpwbYx8LfzPxcNpEey/0Y8yC2Wh0kb
z4nVkBv1c/ojabn1G4BP3Bd7dUOe87OMD0LK1/Jr/7SDWDRyTUGlMdiwr78qTADC
chYnZqRRjR81rq84CyN1u97WmvVjKsLaQJfF/qXmI75SizYVkCJzhs456O3zv2WZ
LBR6KArxDpNIMi/2t9migEKdm/idh1k5pYC7K2wYcraQBtab9G4Ofh4EIrz3zDJ/
3uuWLNatx8MyLNc0AmSUpTKKJpZjbuzKzhY10C76e0phyr29CQm6RaDEwVwEKRXU
KXXqlYq5iueyRWmxbomdbY1y3+/tQtjCHOomNEEXN+HajHLzy7vK5P4WbCT1YxeB
R9+Ne4H2zEV13JmBk7UqU8e2EK3AWT6eltghTCfwyvdfG8HsG993D0UpRrm/L/kD
A5c0aH74bIuCgU9MGW/YiCLgsm6luYavf+gEx4Cf9QznJ+QbwRZJX/65tM8jBB4a
1w9fXeo6pKqivZemw6IIqYMAsbbZubwe7TrbQ2hg/dLpJYIUfBWhDZfS6UEOqhUA
/Hyq9mwT3U5REpmmXwkbMXFBY+iWfojKKAmzIebrd6eyO1Q8HxrNGGzOr1miphSO
/1696xzh0YZuBJ0tYycAqXUtTiJkK3QbojTgQlrHpS6HHHa18sqQNiC6CxtWBdTa
+hrojlQB523dK629rHAFsUa5kLheh2A2tfVotu6yiilc3ykjhW5HVSJHrN/R+Dl8
wftmOooly0heCpYAcUhz5Iyg3gdWoy7vDcD+zrlN7sVmltWK7tS6V9hz8KFI0zgn
kDGdRGiIXwK9ScQwvXAhES6qn3lF95sWFI506sFhjpc2k315PTggErhFoaeGHyWI
mYLS5dSbuawfls12luxxeqGUshGa+iIouPXnVIo8DL2RUG5rIbLOIvAOUcKa2wW3
owtXEqAnSJvHixOWb/SgYdOt9aut5iRkIx0Q3A3PXLgaMGOyqz2HC+rHkip8L4RS
6XV72lug9T3rGSA4N118oVHO14nyHUYhvhXaa2fK7H02FwWgWLlJ574sHFVDr6sZ
G0ozFBWUXsuTB2KSFmRjDZn3WiczjEejaCqEyeWDUOKwMGZa6Bi0vaF0iWraBkT3
VVvURYnRqrb9BJrpVFl/67drotLR2n+uT9IXTSUHzLf4QJCvYnGzZqhrowfnuuY8
acVa3WcE3nNo6LC9UHQ1GLhFNTcvLidVmoz3HkCdVbrREaHw2qU3ZARCvMdByoAd
MSwOn3fiKmVdnjPxZF/3it4A01OpicGU965p0cbS4BvGAB+0bU4YQdzqSTBSS/WL
5WmewIJO10Mj81AXO/m3r+4Vlknb6vyslaAdqEtAA59f//VzCJZnJKinpRXf8e7G
r+wSEe8w53shHjOiClZzPpWKmcdGCpi5N3LGx0rKb+GgyY7XmC0jonvP7zKN1oi3
KOKab/iA+23kNA4DvZK594ZaLuhxXvobdbCjc66COe1euboKRscs/dFBAFF5Jucv
MsVzaMOAYNkvWvenlPu3awCtQh+tkHm7YQwE1A75Qy0QF2a6xkKcw390qzaGe+CK
vsJMMLHcqf5MDORCDs4vgEoa3guK21NlJ5pPF4QQvnmUbclDSTv8tVRyAa0KcFa3
HAzIb58jeEUsvmp0tobLJfkRvIe0xdj8QUPG9ifyLi8VAggQjWT1MpMsN8k+qo/e
KVf0o4QummWAJvteI1FEsTRW08b2gobPBk4o44mKDJ/x+n8rJ28ufEZUkE+1JcDq
3srNsjm2WETL9olbwxpPj1HAumKGOcGffWj89THzfyFr5A8BrnGjqOvVUKOXt2Mo
tqpOMtiCYjMfk1IAqXYkP6sGgdYlooP5PPf2Xrt7K63GMG6KO89/Hd5ZVOaVFKaJ
JndyufqHhrafxfqxFS39IGAnx0TtrV+KVAmmvXo8IpyCRe+1FD9GsVUBhoZjU2H0
6DNH8BSv0XYge22PapSiimR8caKM4dOt/OLIN31wiuicG7Rt3aA7CFX3Kyon0pA2
AbRs0HWStyvhkWGCVqDNx3xF+5hjPAwPpB5RVuGPoP7gTyVM1WOwGczQBEVwy5C0
gz7/KqJG914bpzRD5HqbZULEMEmGd2I4M9CeAwOMvJGZBlM/tGVWTwMS1nEDgn5A
S18eTU2GwOiB9nL1yzij+BlMkPEM1ROsAHn0U8nn9jblsCVCodm+mqxdPK/HKpnR
bsbS0nHnH0+7DL1xyYHeMJabJgylQ4uKpRT5OnLR4WcjdYfEe6VLyR6YqCA0BWKZ
+O+pfs1CPj2tImtFKInIo40ove/tePVAiZkiG3cKYYl01uc5o9yQn8FES2s6C8/R
LqXNepWG55JmqR4wNhPSlV83NEiRuprb7V40YAUtecYfTbm096mggnjQMo6JQXks
U2J57hJOzx1Z5gfJr6CZ8N7sCiR4DCpU47MGGErCmufZly0plVCJiNJLhTpK8iVf
cpcwH+7F6pmA2qeO1pTZKvFvBBpaB92nLU2fwSi/yQGacAujyz/Yijjy00A35fIY
EdMp6T8RB/O2D+OvE57tTkj1eb+JdMyestlOadZllXEgZySwWL2kRqOZn/A62kVI
0X77DM+syQcQ9Dn6RQ+vtSd+J/DEHNPFsstepAcmD+xN42bARKT0EXZwvODzuyIl
fdfeFpTldtrp2UT6DiClNkpcqM6AF610ZKjOvKk8X9b/m8L7in+f/KyVHz7eVJ9C
EXcU8fFQMYvMamPNJSe4ETU2KsngIgVJ/9CJMa3DjdrYf0gaTkAAJ2eCh1I1EYVg
seu8YiBbFsF9BdNJtcfMqj5XyT9Rwe1TA22ET3L7cw3qZ98LSkhqFaPf2Hq3NHEs
zX/E9XHYpYH4E5nvfgwIIDYqiuWvOE7ImfCeJN45F7+KV0YerF8c0iAO+RqyXXtF
Xdki4cNxlYTjxmMmsZuCeEg+sV36ZGuTLiIse5h1RCOXnq8Z9dHPfy9O3/4WHV8d
+VtkFm+udWCl6dMCzFroJatpR7Q5rRpIg1XHSWBTiZ6ajViiut3xQAv7+E+SsmTd
zJVNPftIb4QqzsUBTVTKk25qPKwqN9OQYnVzA4kpANxXqFvoLFTYeFmtPhzG5Ikx
LS/L1/3SJgYxjZqK8DDmjTI/1LnPUAJ3gvc/3yPeRrUEXgms/bVAmumChOClglgz
rLAUxyRJalf1Q/B3Atf0+tOJHYZnL6hoY7rJlpFV2nGG9JkvBYfxQ7zttaSqkEme
TbmyvmXLSP+Vr8z25rp07bMEUHq28oVh2bXt3I1+xL6gsaclOZamBOQ5p4kWyl+4
GBEMDos64I+SUrE8IwojXYH5qUgWc80fINsNgyUG7ZJ9hK9JMujOoQrLtzhTuaPs
k6Hjw309frLICeizNYX2gZt2qbGPYNNjKeZosHhL0PmwlKAacITVTfoK92YtIPIg
lx8HkEm1AtrVWd/9IBLM38DPosra+XkbDxq/HcadTlEV9gOE5WPEtxErH9loPvMs
geLRRY1TRDeoVruwjXJSt6/jATYgWcBt+9IAP1HLRbRjnq9NKS5HH/MVO+Zu3e1Q
USrS07g+ESXO80rZaLvKTMjVfgelNATiz4H4D1OiXZpDGT3M+4LH1FKaWHWfKLbe
Jm4ehvHigJuEgCzKFHiRuANcB3DgGzB7ikRjxxH7usnslykVJNFeWE9E+TstN30I
O4XTSfyq0v6zPPYgG5JJ7S/PWDzwWQyTrMtNCpyJ29o+/kmkGsoYs0DCLR3PnOkX
OHOlYG+x8agpSoLBNLRrsfUu9F0xTn5VYvNvnjgUHqwP78rtsU7t8B0FnoHcTzYs
sYGhg5lmuenYgEVudvfxXdnph3u0KzOMPvcCqiqYfySstjMZTUiEv37jNJ7NEk3i
EDoCmw3pDTsAR7ZLQe+30Ilt5J/F70Hbp1JePEYf/dmMF4qzLbjlBR8lGIbs/gPt
QighJKnt2VFLWanrRvc6pchqQiDuEq2UTv5whRIEFKeC7x8vioieiSy0HQmoki3b
toBUSGKCfgaSJCU7CDU3xtPj81cN0oe/1hpHO2bXCDu79WIdVU8Xb/Sc7aidV1lE
oBl1qh/lE2LvQS+J+4SYBLAWjZ9wivrrZL2TzYiONtSbc1XLBOXxwkjRjsPd+0Z4
RMsZonLylojmKosnt2G13E+3E+kflrHh/gqnovP2T6t7tFAimNwG54STtl/xGmev
wLZg1V8dI8EHMI2i5CiS2I759feSZawbI7fbZMiN3F0kZxBcH84UfFVbCIqdVKtE
rS+bKf4pU8EIi7HFKRxr8c69C2QVHE7Yrb9GpegnmecwOgi/vVr9awf9xVkyapSW
nrtPYMtdD/KDzaIMUwG9G0hAQ7paj7PoQ2CPBAA8pHDd5D3HpQK6DTcrmGveJxtr
IGxlqncvfe3V407TNYnFIwWDoYSQGpz6oqZQinMcR308H6FfrhO8Sno6wODeHEhy
gWTWN+15wIUGcfHAv5viq0gj4ExaEU65HdSJbBPaiWlTI9qgq/5OelGD3vol3xg2
he9H3PxSUVCNRlhCY8mmUy2Gqr7rC9HpHoGe/I4Emhd3pxYJk0X2mCS50gymGDTl
e0SCV52ChxlTY6jju5KrqLXaoaQsXhXooSC3ijysWwAWdNSkbvX5HLNafiaEWLhV
xVAwyA+REid95aa499KiVoDXMcrwyLOPU9Vn0vFFDpDnXBurM6CEHd9/IDSi68GT
/SfbW5+4IDkKc6eQf9iBxezlU5mAfMUwr/tSkBIXbLZmosPwecsicYJSEcTjSd45
DIXybhvNnDU4S+axsPksc2cbXWKKK5SXwUfFVg2Dg0saNgy1n9iFcPT6Se7z5nAf
+IyGiRKr1mcpxUXrGSuMsXzuMwD6pEaWDOebCya7nKGD7jkfKuspUxXuqI/vSFm1
lbCO5azZzFy5h0gTEVYXMR0XB1NL1gcnXc5ShE5ierU9E3+tFoky/H5c8FPqsVZT
eiaN4BISUUr18ZQ68gEItUiIPGng4lAiQl/aCwW76c6UFq0pBu95MU4xAVt/BlVN
1Rnjt+Vos26hTqfRT9uTGdEZbZdBn8NjOqEz98WhGmtAT/utt+REA3K5JCq8pX4J
YX2KIWyTGHcHim7zdZNC2q6pSd/rYXyzf+0WC1QleUXF06SThO/DluXNTBPAqyLR
qhBZJ+DY/wsm/8stVvkj5x9n9F5GuFgGpwQWSZTuGlWjl9WNcT1oLvdta4F4Afup
ZxpvOiScEaayyme1LYwlLjlxmxlJbs6jAT6dqo2fup54UxCDMCBEalDOm8P5z35U
wvYnDKpHK+LWzepQW/n6EQMsVW1bXBZU+5EayxtQpGaIT/Gd1mp6/jlrWKQ7Cgvy
PuWLPpmyafFznGh339hLE7Sf6WEmBGVnpxSGEWjll3urmPT0S+2XRPxdhepjkupF
zHOwXH1JWd8nCCRwY5G9JKSUu+CQTnZEFIk9chHhe2oV187oTFsbWSUjnoial5nO
9yCA4Kz0o9an02oG2Yvh6rWXrOb6J/N++OFpd/1DwOp94El8b1fhJWbrLLnNLMQm
POjz15CuWJTgB3um71vzi0HVUfJIbHH5VheR9rBSH2FEMAV72UPn3SJfPCZAT8Sc
0JwFIjqpGYgm7XrZldGnk21l3Sy+HcGN2j3Wzh3XRbsb8Y528q4Y9Sv9GKPUnlbP
GKprp37lpntMSgL2PXeT2GnoGDQDCEDxCxQruBR3Bj23gdJVGcU5V2YGncOHgyhp
HzywydlXyKb4bUyZLNJEB2avpmn+gmJpiWgn7Xc1GBxUtA3StU20A0s8R06Xo1mu
fMaksB3Y8sjJj3XFXYIa321x6ViQacdq5j1LLi4KpYkanZjkPUj7m4fDSXRfsX9R
kooOo9X8vCkCyQOxftNp6bcEviCJr0bTj/uAeC5iGVb461jyHhRzshkTKRbrjMq7
takUcj1R8uC2m8+adbRbyvz0P4PRD8lCUKtU8NeSQqWkbN9WHYba/E+dQ0rjBRmU
BnZxJpX7W7IlaWY4w/tZ+DHzgh3mgkDoE32IER/PEJche0tpo/mgwlRugNnl8AEy
M2DYIcs83l3AmCbyOch1Wl+RYruXnuucLESFfGhbgSlPGgWX75yXn0io9g5sKDBT
TLK4bxh2DpZYyKlY8qe3ZRl4CPBonXqg2lRvYYjb1tNGxmDUQkEQ5VceHIEdCSQg
eK/aE+WktZME62gaeIqmRh69nelEb+9lXuAufRn772xv6HbKjgmDSUY+Mii/Zoth
3dPaAc12WkbNeAMg+uBlNEsKdme2YxzwfjRRyb2VZMOOpPU15r2rT083l0o5jDE8
hmWqGJjMW0oN1v7R6L83sKtKCc7gzacP5vF7VBdufyqUDPZNRMCs0EZUMxNFm6Dm
p0e8AOu0E4PfOjAFM01JkPehDwST45jBG2k+ZVgAWwu9LvOine840TRBd8jrDfm1
3rqXIOphVLLi1OKo0Nw8a+3BMhlCh4VKK2gT4zWZP4xh+l2H7Efm82STnQaE0Vsv
y9Hv6WYyL3Wh4jK+JehP+o9DFlEC+r6+/+TGRPYvBUX7BsKIFzpvn2u2ppP6La/M
7rFy2wJpRobC2kDgeuHta7IdwRPlalDNKWTAsADnv4WBvGr91Y+ptwldORBxc5eJ
YylCmHWQdC39PzT1yDayocNmvEEHOMZPlGIobsPaXb69GYlnCo+3Yzpusg2FJO86
Ilk4dTCoECQpjBXDZJFiCo3dGSPtxbGqZbp/dLz9kNgCzfLoEwvuemOYuGD0HNt5
8SoOQlC6HgSYON8zFFHA3rKimpmy9RgLD8SJZ7ly+6/gN+P+vR1OrwZP64V2Pyvj
paAsZpcxE5zDyvZ6MI4N/45xT/++M7hQTmGXTTsfztPgV5VPCXs6lrpd11mB6lks
hzm/ClznBdovJhZpscEUiI+xTX3ftW/w1lHGhB6lmFAKyh2qOdjGzEOv7yboRbp8
J5gOM8jSTV3p6UAAPIJVS0HqA5eF0udaOEpCQHAL+hLEdt1nZTf3+qlYN+39rk8X
7lJ+zkPGlghDHage58f36djI2fRD+JjTqPTjXmfgFGoa2Ned5aiipZmQeZwrbKdo
eBJ16UasWS9m0MM4sl3DCOyl9nzOU91nn2T5FUfjQU3yqe07OKsImrF4ru71T6Df
X2YHaTyOlsDTg3dH4Ffm1aLOMnTehGTrSZRHJsrFk1z4GXX61KLXCcSZKKnTxjuY
+nJan1klgKQU7K4KH+uT4ecQzmBgZvrMgXO1BNzXFFM32BxABRl7LtjAT6YOft7r
V/Z+QPeNiELMSZkKIllQbT6twjhTAkqUzGFPm1FN9i5rnq0X3SCt0i3wnxW53W9A
r6tdckYinK6FW7fmaEar4ls0WaNPWOGwFxJcW1tYmgBLSHXuAOm9li1n7D5JH3B8
AdqFVivhnBa4av/Xm+i1gdlvIugRpMs3hUr0ezzq7nhAUBvBPwxz6wj1Dy9zMOsl
/4Cdo+uMIdovQpzI/6+H9+MQq1ieuYPswOb8KNMH0epwbbN6J7KOz5abfD2S2ZdO
2TnINPS17wXYXCvF49elXec81aH18X8/KQP7aKpbfq96HpV4S1Kkl7R/BlVl/fwN
cNDf3Te7swoNwhXsPMCvPqpopYRGbfoLV8idxdQ31csO28jlbNurmUy7u7baDqQ6
aqmwtKZ7qEJaduGdrUXQmQB7Skn/dgpwRq9zSQoe7W3hAV+zudIKr2ljtPlk0NCn
HqGQScmAsBrAz3XCS4ZCejOGbx2MQQ9j1BhQGZAzFdXTW7HouRT7fWRtmI7+nTY2
X1T6yS2wPZgkcGBQ7gMnwfvkS3hAoHiCa5j9SKizPxVudRMkw1csCd4CltV5mTi1
YXkYhYRJNTauEr7Lk6cdFVoBkSbudzcewUPsRhZGo8+S1sB/76zhREhB3wFCk/CE
sMf01xrnJKxP/nMRiq+R0qfOKeVaJBAomcMj6Ssv9vmcuwZjgsHEU35Zm/rUJFPt
qU+Qn3KQ7uRg23xKDorlNWBCCAZf4uhBHbPVhtgc7F8=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EiMh6Us+5jGqV458ZVglP2ARcVKBa7Q8aUbrqWsZ4gblI+otmveuDGgriCEqH9iB
Jj9dKqZ9wVY7tAUE8VvOPxG8765s5Y/ON5fmVsQGWUEJlMeLAg4jPKaMZCIQfPcV
UENTDuEpyjBUUx8oOYIWXt6abgNPEN0D5tMs1LppqwceJtvZ2psYzLIT+tDe/Rdc
tmOnFoYYlr7Rt0acwbDHNF1HLZMjp3XS+VxHWMspCYi0Zm/28Rl8M8Vo1YuTwM2F
glLvueQ+ee+FY08eqjXrviKtmzQr+F3oQZ6j77KsHblihdoVHiwXwJwUi2yC/51+
nodfNMWgBLfOyYkDQUR/cw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6272 )
`pragma protect data_block
PKcHi2DUZPt92ybn2Qa6k3YtCzHBY9swjXv1GXop776M5Pz6NWDDfhgWafOcuzva
iT/Ur6Dm2ogHFglPtp4kL6LGSgLEEU/OHRX5qVGWo0kio5QMAtjekRpbNIP6uQSu
HHeuZkfxiuCX/X3mFxQoLDq3Gkm10PsjjsqtCEkO6kcKHZhjLYqDUiMcBt0HH3cD
42lH6cE9EtucALqpuWemMw8aDO9jDHL8ZnHsO9Ph8AMJpIItLpGAh4Zli4+B8jen
t82mHnHe9FIsS5lrZ54m1CgxilsR92111WkhL99g7tKYIAkAx06nGQZ6BhIcbQqM
qkB9moWVJ6+CNjbi5gSayFDSObm690Rc2soDhqLlXoiIJ5mcO1dXMsHpFrM29O1p
mgEU+nKS1IfGRAkL/OB8SCVLq46qdF32wlCxzhZEDcVcs+u1kCVfdbB30p1bk/rz
Ka69tKJIRNbq+1x0EZ+yyboXfAvk896V92tW8/xoXLu0dMvIADZFS7q/xmXCE16D
gyfQK8ZC/PDqEMuZWlLRymHPRVlGmsZCDLVqpBbrf0F2ftH2oweEhf7s4upkE3z3
n9r4suytedadyC9cwNpbaqpOY4V5mr6j/6vUMi6+XjH/E57JAOA2eBLWakSALUML
07GlTdEPk356TIVqYXclDlhwhrMfAy3Odj6Nx1+ArEBO9MPKLx+IpHHcQ1ju8L3e
SG97N9DKtvjxNWx30ihF6NfbRNJxMaLP6ann8mJQy1f5VEQpkDlL2SxFN3x0ha5c
Z8LrrM0a2oi3u+BESpq/7+6w+bmPNx5lJCC0FfYND0bdBS8SBuELj8o42bT6VOS6
d4pDmo2Lbao4PmfWnGrzp4VdMsUhJP/gJdJh2OSVWxaBLbRKzEvzRkUIfR94VQja
HcAYEIXNFxXLmmXMD9aZL5gYNndLYcK4MTEkL/g4nGpKeB5gHB34bynC6yeTqEED
CJ11VDEXvhwpFC/2F7VP1IdxQjOfEytDvmUR22dWKAJvLzv8exI60zX2rmKcdKCt
ukz0m8Ja9Rgq9HnbJWExmfW0JroIYHj2lKv7GfuGk7lsAzWvPR2jjFGe8yr1TUVl
M3SLTi7VE2cbdalgc1nZ3Kv7VOLZJw4rFjpy7ni4prNf7IUrTB02mQpXJJP83kPG
2Ps7g+f041HOrQf1R7eukbQoIaPcGq11jSBEDQ7+P3KeYpEXrZZK0wFthUlcrgHW
f0IQz78/z3qijaQFvOn5pMYLNGH40elOr806cAfNOOzbBF1trkmiVWAQE8k6FxfJ
IrnpPyAoEgcWoeWUEXPb+zumwLvgLk+5jE8bczfWr61SbhvAj3AVpNwNxoDoKwvL
iFF6PXrou4Q2dCrUcHcvpKvx2OI9SW6/otOW71vzTjCzIybGOhDmVlEHRClH7XPL
1F6s0WttSOwtbdWcX79rCRBfrVx25KaEZZX2Syi1EGZ/asCujva/na7O3Ssqz5N/
hLYED2qMk9D8tccqR/23rU7AbL7IrGUdl2l8KBaMgF+qxFmqXm4v1y5NtytHz2jP
f7NdtqXkn5lB1vbi9VeV+RsCNDOnVSEy5OK7+Zgy9yI7/X0xv5iK29hkRG+7OkK1
U2p4EG/+7RZfA7cXUOan942PLqTqiabM3k7CC30VEHAsNGf1k6rY8RCbgprKEbSs
am1os+Rl3moiXX53KiJYnHbdihmjfclcUqHUMePfR2Li0ib/E8Hmzn+WzwfOGkP3
brQR7A9FU9akClQ0qImf5yO7px6yAqF1ik98D9pFHMnW8uC4kXwBZAJWojqWWLZJ
ZeRrO5GN/8jn8EJwHGQQMJZNyzK2x+iqLMyQJi83btot416olxiqxCZx34Jb/qcd
lLU033ZekwJHVYBCMmuElXM7bp5kacA2hGc+Dddw9cw5GewKJRTyyCDIV0ShYsZH
GbBbjMzH2562lM6t8oGMI7/QHC05LvxbglvOLJKIN+LXLwMDZwbGTv3lCUeGn7Lv
bXdpIqEgVgdckg0JBi147tSlnLCX4S+Ois2grVgLcWhYHMD6e2g1Pro5HGP9m+sf
7BpIcaBCJeOvxDcuthjxem+dx0cG4EXeJCAQ5MH6wyNx4D/eN5poe4WQlmPtooq8
B0MNHBEh4DxbpI1jyOPTJ9h9WE2SjCx63dBUFhWTR1Murwr0DU9PqykBZml5UOIL
I5vPX8z9QPk8C+LQ26B9CuO+GuQgpjuvNaQapTQHHMFv4D1fhFdYY+E0w+mUguMk
nTVyZrDEeL2vjSeZlggDHAGeCbMbyjcVxZpNqQrsT8MP+Z2Ke6Tn4o63I1LLHL5D
Q+e2bgk30E20Z0QRHoOJFd3xZfcL8OegIfA6Ma4zydm2zqyW5kKteQqCewzHsfFz
2WNBsSJyCaakHWvhcPU2yBzRFs0EQ7lKAz2EULb16X9hptkm4xLYbBiKvwjkP3eM
ecJvnAZwtqBacCnnB0cyTlQcVH90GDeOE/bNXGi7plFzj4ElW3LpLfCy+i1wmUkz
Nw1cQZoRKouJ2p+bOsgxI/6z5WGgBNv6XH6P7qI28CfGRFPBA7qhRObRqW3vI6J9
ZmhAJ89cb0CYg9ECcT8tTU0rvJp+DgXG2FUMRgZPNDSaV5wjXeSdX5GDJ4UcKWqH
yeyQK3rY5CGbbjAZ1rF9PwNuJmYTQLH6HrDQBh6Evtgx+QsfV7vkSTVE4LiRf6JP
ZwLTW+lM+qXPHoz6Ef+v3HNpNGY6292SgcOhF9tZ67XwagAps4bpUFY/mUI/xfdf
WoxrzVzPVT5WAX/vmLRY7dbaTG+Qmc/869nG/qjfFBOVw0z7hXoyeJkwlbmoNtBR
Gv56+xCKqNtPi1U5imU8ZhwOIABe4Kiafw+WbkM1q6DnpAZmM91lcgTf0A2UVx9j
JeDYDI2lMXxS3cAALSZmblZrM6MYzTNXsV3aek2+wh1TIcQ4kWU8SLKa8uaIZCp9
WYtvZxFKjboPNRcc8KzYeLREvP7nVQhCwCHLRI0YuZoIABWDlf2yWuY2GJMwRvhE
hqCOpc754Svvu7ulClU+9Dxlj8UOtALLUsnC0Oq2wKXeXU2ZjNvkis2FVBfSegYD
S7VJiIMWjTkyyTPzVhx3vM8VNOyvUVP652hEdLcvF4Vzj9JtAe1MHnWsL4lnkgHg
7bs/p1vxVPjusRjmVWVohvfenyx8L+WdJSOihvJh0IVmIoYa9kgjJRh1vfit6KJz
AriskMtBWKp2AdHnOQtEOGNxcvVYYpkWgKkU7UApdXdnywchzkh9FEePBDgjO4Ay
y9hQDwn2r+33hNF2On3MN363QFSGfSJZhhyxctxomyFlFthgbPSsel4/lEz2sYGa
LUyj/z15bWAyh08aGy8zc1kVG0u52ILmwur7mtL9OM8/nFtqMsyTPTxTRZIv/W2u
Nb4Kg7RXHQArbMFlLgIYTPO5e0vImLUafEkTYWw30LsG/b9nIoavQW6XGtEwP26/
x1mE6vzxNhoTkEfkVspNVuQs7rkWrgE/QteB9zQUc0DkHCBi2V3hjxD9peSE2Css
nyRGJ7xnbhRZ8ZBTVFATdMPtTTVvYpleI7Ki62UNekML4qzu41rbrOsGH2qBKkTd
Piwpcs6JBFKPIK1IKaTLoMmFDbW8BXaZ89RwW335gLJ7kaQbHrngtjr563fNB+oX
ygcbxGnEf+IuyCkZwEqZq1c58YWo9emVdcu0SY3z8LQLsVnXvGULvUp60TKeRTTM
F32Qr4ZduC4KxJY82n2BpaThQsMysYa7+nlILHvPGUmpkY4D0yAORmtuckKR/sWl
zxG3mtofaN0C1F17GdZj4kbV3zf3fElIj27PdHrPtMof1PMeOKGvX7MEaTgBQziz
2VSYmPgXqqhteXC/9EktBZxM+yjTzHXwqeX/nJKLKQotSe+ukQVwg2Ss+BLsf5/k
dxMSa6XEQFdCbQxj/e7G8I2QzIAbRHVBfObbmCwA+4v+0+h4LcWBY3+QNP5wPntA
nLrIlvawsB8sx7ZtvkF5b0BjBNm2AHvnw+S8J3al5Qjef19H9jepRZcuLo+igPw5
7cFR+/zDRKtWtryu4jhVRZlusy/9IbEh4/6ZPNNbCHLaw3gNSaKI8YkRT9irt4I5
sH52jRSZ9BQ2fUFJ1DWwbFEX+JwLVIvyUcc40phLe+HSdCknMfjR0G0U3Vt+sNmS
ddEO8jYjcp4OVGwtprm6TR6oIRmISBKynHVdQSBu/iXF5CXB+X+JINq8VdhQSjgx
dwoQ08+F/CW7gTaEanfAOQFzA7X0JLnRA/4DxE6H5Z8RGjMWIuRlo+S5ttVfcwEc
U1kE6fvyvdiit3pyLWU5wruTAwIpCGEFO7ZoC7S8brfP3aKIoy4kfnTLbufM3S1c
P0xAgmIPhzBeAzOEDvxPVa73TN1Cy2gnqb+vBMJ/MvvOk2ef/t2t9NKum0E80uCG
nNfYm8UbUGoqIaVliBZm/Sy18mnhHEnaPUxEax0nJCqJ5NYy/L5wAQYBcij4N8cR
+pSZCeE36f2Haaz1+m7jeP6psKO508HLay+mA3ytdY+OAAoTheEZkat+I6WMNzH2
3bNoGQ6ogW2YkFANIjy2SL3JDM9Zy4cMP0CaMD+/XcLMMxfYyoES91s5b+gK6+pB
NWlfZAeykN+ngdHq3C4G+KsD5SbuRUVe04+iCt/cRJj7aN6Zgxgm+vaSnhDVgFZ6
OEhYYk/NQtR6b3yyuqwFREmy1Rp1IUlXMvmPIwPozsghCVTNSJOgWn7vKvhcoxJG
zZNHIvhuqdLuXaJ+ZBD4d+0PmPTeGo5OL4p5+VVVuJr/1sEC7cRAee8j5mWuLr5+
m+835Ky1Ok2oEupkqUhBXOsilkQMDE8esGbwBO347vAkWbGqbjK5uinepFP7Pwph
oewLFQiOlfIp7m4a0hgl85COBGUWGPubTIYPIeXe0VO23AvWcUa3RNZFdyGzz6rH
LhclTQEWcWjWw/8Es+pVN135alXbCrj/v5mkvVT14Q5TVWJNKx9K0cD64p1YZx0U
pgJDOZ6/FcwboLy5wOy33eh9ggXGaoEAKgSGc8kh2hh4FmoinddnswcRRSx6uSgO
UwC+nwL8Sg1q6WOiKwJMytTg75S/44IoOstvnp7CDYaFmv6Rdf/eafQ8SiufuaQA
/loch1TnfCn8o2OeKvBEefn6z/c4AG+UWaUSVMPh0P2c3N8xow6FnG13Bri6VIsY
ECcsexWs1dbGk4i68K77naIDDrLlVc+LSKajf5IUDt9zV0luRq2rppJhTZt0wlRT
bBHpqbs8Ocko+0ej3YOZxQKYo/723EYlomBhq5vl3fFcx8QO9NsXM2tfL3G2wNHv
ZdJQrh+XVPVV/jCP1uyg4lwj+bdKem9sH8BhXuztinZZ/ohAzwYMo/ucOdi4k/rx
0NgW1r/BjHrqo1j+mgmVG+Kr0JBi/WVgSZ6gC+hMzkbBgLfCjg8o0hK3ex/uTaN0
1vBicO5ch/rREdWRSZMKM5QKL3HGPmGUUMKCn1bF/LqIKYOdWm1AeYYE01lDMarZ
p7dso1JQr3eWpb6pyv3k8D5X5gZuO17SNYo7eFAa7eKpbe9biLPWn/8sP2wOwGqj
kddePEG/kuV04/YF3lcTIt0YfzlavD3XwpZti5uuBm0MNbqBfVCtuEWvzzvKugBA
Yy4LowM/U1AVbyFSanFmJLK4iFCjsBdaoNTLw5Cd+sYlXnHfF02hWtWNSwFXQ8XU
GUszbRQsIGX79DySBq7gejki0X/H+/wUoi+7ZljCDtVbhojqw/xbowlruKvmMdTE
vJNzqkAXX1bzznVwjE3Kw1nShLMoMEHozkXQsT6Jlxu0JcEE6iuEj2a6XhvWeEHu
isbEMB5tgTBHE8iGS6XKSrJnfkIT+tdGnMultlFKDqNKP7PkPhXyKNd3kH9WuAHY
iFIk4QnqpTppLxZeU2x93vZcpJnLNN/0BpWRR+fbNuTS6dGN1QlYMoNUmGMGMwvW
k8o3ts1dJ+sbxQ4YEfGJ535XQFJikQEbWeLltFyxItYFQIs9Zy0DIUVq9kw6L6py
0NWgwqOziMLuhe1ZyIJFOsP8Tggv8rhywciodHgBEIZO5hZLIF2IXYZBoli/FX5I
FFvhFLkYbehGQbX2f61AlAmbYqZfT+mmDeUJHRxZSDawvGKdj2Y9wS+GHlsDO9a/
iMnlK+gUNWDikyHV+9EVf5wbIr4z5OOpQjXMrFyhqEsw99aCXRheDd1PPdD/eBmt
ZW8OawHRiUefAZccauJGILXNMqw7vM/h2tQ4WAaJkUnuVmcWjKJOOX8TBNF/B+h5
lSo4/P+dQQXHwmclpmTv8DG0Qf0SjZH4Gw0lQV2SVl3il9zE7JU0M+4XsFE/yuB+
9j1r76RFeRAIO5r+V9/RzD2TOQ2R5wsj9ygQtIBNYmKnCdDPziSYH9VyrU1zEU8D
oKJYzW2GLG/nCZqKz7rlqeGiRLZS60M3m1qiBUsELBbAxW+Z3xS/wJ08b5dA3hT3
XXQKxd0J2fG4ekrM+TkISFDMH7Pve59Jy5yqb7L3HQDCpznJqndlCXZx2aXb8tKv
ETwdF+fSo6oYfDlVfwV9xPpuPwDOrAwuRh6N/wjZs2uXdalvkN8UdRKAaMypjoMS
sqgLvjixbj7HI0e7np43XNV58N1ZfR78DRd3p2DrhJigykz+bODykA/gC11GO318
Wac85NZf8qfqRwXFrOkPrxEsZMc75wPflu0ob8t2S5upibx2eTd4tEdNe0Lj+lp/
4u01jOziyxLRxlcd/NESuKiBv2aCiBaLdxZR6IX06ix1hgRPfWlPJ1LBUs6d5Nhd
dt8HWt+8QHxio0cLQRMMTVhm+X8nx13duTmQpJMlSOmvajKJ2Ow2sjUE5vuXhzR5
uohE6r7SbD60LGowVwijosBw0LR6L2MbpK9cx+oKJFe3MhN8bPnRnZrAkjVA05rj
yfPR35BghH6Pk4YKBa0uf0TDxRbORScbPN9AohY8ej+Q5byYhkbIc1jsi7T4+E3N
43HX+7ttiIo/W6QeqmdxdmwWL7uRPuTeRH0vfpJ6OGUJEbhmKk1Hb0wL2aHkEWgm
gnMswWu7EWyf/ji6190y9L+ffLPIVFMjH6vbFqYipUuJ3TC3qF/LBwpEVfnt1iAG
66CxuBauiODgAnAOubJICOBsImB4LhjR5U6jwvKaoM7uwnZSifhaDDZfOo5Z/s3v
SnhJvrembpdRFCl095+Mo48n7b9nW/bCTx36egkTFx4Nv+BJDAjUWjlBbiv/UeeD
80vTv8J6cFLISRg6JMpnwXaxVnaaeH8+yrYTI4P604RFepSlH6qY1CfL85g0RHor
1RSDtAV1Ddy4bXfSHg+c+5AoZtaICR9ZTv6YVwkjkDHEDwFx69u0FkzdduKV13Nb
UCVBz+gF134IhEowxLvpKr8Wpu62gATW6x4OXieWYz1qbbRgT/3v4Z4hapvAnGY8
5WYBhHB+QEEJVEAVj4oHYFWoMCFLUWV1CON+glHWm06FVC52/UqTEnbB1eLxAA4J
v2oZZMddqJ59DlOE6vHQ3n7zjCVH3YsEXowzm8HrjBgiNWWPn1POjGE8BVRtGvsd
Gm6nyy5t7oS4N+urnEQ+qXpnv37Kn+zXnPu084V8maK+2mcL5aUMDKhfH90R1V7K
5xNE3ZH5z07qa+K2Xd8eqqk1UIoFOqrMxr4dKEVHw6FaKx5Ae3m+D2hU2Je50PIj
H40K8f6Hy9mArTsY89impN48FbMW7paImOqqdm7tnR6p+p5PQXAzDsQww6zcgErA
H4NqqwCmc/+CFzsFSh2Wme1yDsIQ28OlZALt+5ia5RGIz09W4xAcpxEw5FHg40sp
a4cjZ1TQJDWC7MAQJXCfBRWtMQkEFLzbKrz4zqd3DzHFFm57uvk0UWTnkPjnZnvz
HHGY3C5/BUtZ65QNX4ZGyq1W47AfqohyulfsACDzzp0X5ceZfWNZ57KCZH1G7bA/
yf9rO5F18A79md1048oj7GQMl/skzzVOd6iDWFjtt3rHvfy9z7zwgTMoMuKKrfvT
XQ38AxtLJJEMOLzsCSze40HS3GwOzYlYfOXa362kEHfHdeEzML2/LNoM4rA2NTbg
GiHvETkXwtdj1vvU+uGoT+uyQPOLXiEhl1mbqjbMr4vMH3+al1hhZRjx5id3klUo
UOnsZKdKn3NKtKeYg2Ieq6wAanVXtB/kUbZ4Ib6rG2UXp+CmFUHASmDC6XlbLPm9
ztj0IQKT2IwBPTslwCS4KyPgB2BkXIK76dkSzRATQkrzJaF8VNj3/GzFptcIYLn9
pYGqNsxazt5fXLb3jM+DHAIsN0l1XGQUJIeH1+lrWRDnAiwgDM9jmzXKv/rLxAcq
wRHztMh2zF0nLZDjYSqgAJAene9T9AXFUQ8EOBS3cck=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
MNiyUzyyCT6EvZdYEt2MSmI+Euw9jfZEkwOx1IHT0onkXEs3nnq9IkW6xZKvKtZR
eKL5T6bFCkEw7BD/DQ08dDGPBvMWVirTBhPvHIz0L+SLKykLuYpHgbxyqC0hX3jF
bFJAoie2YuKL1SNRFbkDEODuSqFqegTZm0+SpKtjw4RWyqUmn1BIsMjO2fnPfRbA
zAw4PZG0JcsHrnvtNmBr42wBzOzWgKQ/tnEGR70v1z4kQmL3CcwFIt54zpOjm+M9
eZA+SQRI6vKv+ufdnMSsTC9X1Av7uNSmqrBSGibTw4sOkceVCn0NN384wQY6yQeS
if/TCRQCRrlE5tiqAFhsUQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5424 )
`pragma protect data_block
W60QMb+8jqrgLbwSKvZekQuS9+YqtsIlnojWYlfEVujMIvrB+CzHnmEPTx72BFmM
cyMVrgX+/WKhSEwzCxGCq/vt2l9rAWv1JOMQ1XmQhS9ye5Fr+Wf1gn0wNduUgVCW
kn/ny+CiHqx0U3Btnp+R1i2Xx4qAWNcc9Ln74T7rrkZ7NJZyUf+D43cR4LYpDWKr
RZA8Jdp2t7IMT1s6nRgDB6TRXQ8bv93OwujoS/cuNorhcrOvqjWxWyY1XQvXMTYw
W4rtLu84j18VqvZfzeHeVnpF+57Yeuz0Cmjt3LFUBU2jt129MHrMe718SFC3lOm6
E8pSlJ2E03XGXEKFrWCLMCnNiLgWmBVDFxNKgZG4jlJYm1zjY8ihU6uMddreNn9j
L4NvXi+yvWazhFdIXtHQlQpHNlDVY8FYVPCePuyrCeciYByfiJy10nM+3lA0pWM8
XmwSKmEjwhj7F8yRFewKdZ9wJtcdnTe4FkOmRITP+1XYeXu+vJAFqYUE6aG9DZvB
/jCkXC2nmrQUZ8LX9oYn5wpbnIMLyLJI7J10JfiSUKCy+Hs0beUcxeX7Y4SmW7Md
LadUdEQUqCC0lROg7IWJP3ohhhxUR61nZTpb3par0K/cEcQeiqkF2l2mQPv4mofT
uGi3OU8BoQBLtljPasIE1sWlrdjZVZKKZIBbmTg1vJyDUyVjC+ld+KdmHBH6XhT4
Z59YUA6WSwYw+VZXbFaXp/d7Xi6UljBZP8MEpC5WHLNrVRlcPhylqptCVVrmsFWn
OGIAZDCiW5hXfD5TXAsCfWt9ReThRCKQFWwPVcVEKsr5Q8Q3O0GZm/+45SSlYym4
rfdJOb4M2w+ez7aVMz0xPqwVkegcQGZc0vVYcu2G7nBV4sEYSCbkB9AB0Bbun3CM
DZtwhUVVCmgtSGCRrDcngNV7rjlp/hQnOMYcrKb4CstYWZRxdfZ3y9j7e4ukiZLS
WUvSFztGNnkb27mB0eBsQdt+ROE4VXck6LSkoQZgq3nYfe+xDtEOesCjtAKr6YuC
emZ/9hVO1IZ/7YN7puUdyCylthvSsNy/DND5bJ/rS62rrxEiwT/nqE9sxnHHPWtb
z/aZ4XO7G53FP6xs9sFIGQ8IiPm7KlmJeoDJKCB9Y4vTcDtB5+0onKhaU9QTRvGZ
jXQpNkcWStmgIIMyFkA7eN6kR637Xos6NU1319aPU43H+qNb5/WcHKDz4/cbz5hF
sPUFXuoBOxCsZzJc7eJ7zb08iDJ65vNzjeGTdJqz01iDv1rt7jsKg+yGYCoh3xk5
g4BxcI/KalMMwzm7iZ0HZl47krVImM9DW7djzpaGT2QnJkWCt1qXmRs39UWKlSGH
Z83yDDs9W+swtoPoiR07vfxZzz68IgTeFAHAS65N7aBja7yAevfLhLtnOKYguEfQ
crHx0qw0JY+7qlBXaq6ONIejHTk/w7TA8G1MyHwrUB0CH2SkKTQ9OaPrM8ud+2JD
5NWqRt33C83M7jBM4hwi84+vul+3iMiKDXKznUTO1lA6DkOF1HVvUtrRi1KIptyu
fE8U9aXvg4MMxOwAd/LtAuAPghr8ch7j32TavkRgQaHkmuj1FfkVDfhvfScArXup
7gRwA93/z/nHZTO1jaLYKlBsLnXbqnf5BbEcmW6G8DTirtMxwpRxNQvju0Ew72W1
I0YwfHWj8l+BPvLuWaBwsEy4djEP+k764rjCbmzU6LsXzOYXPVicWG7wC7UPq1Mf
vmQ6+e7Dp1Vg1WBDeOjT//0I+Y4diEHgI1PUZr9OQ03X6rFhXKoWA0Cj8jxi9L2g
Cq4dN+27ROR6Sm98DsjY/y2QLEJNwRSHfQs5ULNsEMTMB+i3JlnXav2Vwsu6KjjT
zCzvI+GCoOXw+N4sZU3HshC/g9+4S6NJEU1+cFDHFGZDVGMemv8XK+3K1bsnqgju
4IPqp95r1BoOXQG9W3IJclMaLNzKmGLXZlEnEywIL2C+WkXMjkEaqHCqBy8KpGVf
PDeFxBpqIPRfQBRFXGOxwf9X9JPfGzU7J34PRiES6GXOgXebSr0pNOHZUTBaSSsn
3o/3U5B05Zi2vZQpGnfAYT589GcsAgrfFC/RVfhKphd1ZtsMtlLK4CglMnN2FTfW
rECFhQpDM3b38N0dOqSRqOxHPERcRAwOAtXoR/fhaL5/d1tX4eLEsfzEilyOab/L
AlJVpwFgrybSMBEApWGLBJzwDdDn6I3Di/u4Y+NkoCyVzqQQV2wL/JdvlxB29td4
f+Zh43WoZzTuRtfXQwU3BcffaodAvvPU7zTa/PkYBQEiTAiYh9Wt7HG0sK2WVKtp
GRApKp+tSifNYmnO28nEWem3VszL653/nA0dDOhLdGGed//wO+QSpDMmtlM7iu8U
RefoGD8FGT4CcJND1rxlcpILaokC6PyUMbXAJNH9Ufh3bkJwyEz9GgPGKzh/KQNB
EIAvIdXecubeqKP5fRfn/BjDPKR7ML3vNmOERNfFF5KsL/28VK7rrlCJaf7e4Veq
as5b4+wRZ1GUjKBHGoO8kY/xD1itW+rvZnFknstnLObnIDIsFyMq9UIYAbPKwPzq
nVkLzSg5o1RCoZfyeH0XjR6HsruX1Lv+VTapmSGf9Z7fFLzwGMqzcVa41/3qhFdY
7wsi1wTdRW/fUwbR9aoFWFz96xxOz1IXPwBIPfHuE8L3iwOAwHyx+n98SV6iQfmP
Se7gJPL7ZlR/Fa8Rw4YQi95Mahq1bOaNiSzUL/O0Rfr74w4QnyVN+wjT5bVpJm5B
sQFNnA01BICuQCme1lie6N6A5BAGcBL9PWoxW6SScDkUvLuS9sJtTq8A99yb2Jdv
0jROXeDDJ3xacxr9uUELmDJYiO6ILMx0hP4vpFWqDEGmkDbx89Asj0qDdWNPrJW2
Tf0eHwmi8Z0Z4Swhtm+W2UF6rE61yCnbnpz7xoDtxHSAUofTp5ZTDSEVYGfoWuZz
vPplYS6r/6Tpd8N/LUJieOsJQBgiV+nROjyLhhAoLFn6HioZ7gHJxQVnjB2ZULjL
ZadMchus4Z5nRD3P+csaaZoTkY/aAMviAD5gMnC+K5003TzOu3eLPMp85bSmYavJ
/mHlUpsf64esuT6Dcd0hG+ETNXQrCiaXDlcwg5mS0u/kPjsMxPsKBculJrIK1QsX
QsCVwc+IQ15I2AE2UgqalUqKE8KsqZXw5My3JVRoa5zS1A/XALNCyX4MgTeJk9zi
YtwSPt6U/mlQjN+p0s/tnfQGVTLm5klycQKOB71Kxr+Et775m17MRL5QBMgJHJ4z
2TWGET8v7hh0uMeg+nPYoHABrDID0KVQv0IRGV7JWWhKzuticdHojCe5/J/IlJMJ
75GCE4u0sow4J+w22gM7RhYHFlob9kranuB0/U88t6AvQizzlkjsuc/gdCrPX8o3
d/DtK44WLNFNQsXuaIMfDonIP0mpRAGzejRhck17MKc7wHeW0TXr6fdhfltQogXq
F4EP5ktCpSIjyeJ88lQUGgrcCi0ttUNQPeK5saxPmjMva8tf7pWxY3aNXzqlzTUB
HlyUrPMfFGAZdxeaFmDezHZSiB6ccZsPncmCMxtMVd/2VMxSevwfEg26+gH1u5I+
B9Jo7Yd5RiqVl6SxjbyGFhNj+mSX24t3ZKjVdRPbhoREtHcurk929jY4jHsNOWmG
YmZmiAaOrk2UThgQMOviz2U/xHGP8UJ2k+FXdeet070ezUlLP08TrN/tQV+xC9Qb
epsBnhsZslpk1Ut+KJ33ydpk+tSBNm3t/m26oROuC/qAo0QPH1f3NFhYVRaHtODZ
5V9Vioizzg7nfWHTWRNttF5psPFT7tWaIiU32ihH3fgh8InMCw3og58SMLsqeIAd
zhU6w+3zkqWcMTBLssEGk/6FGrYZ5dk2zaJetdgJmER0YVqcuUWtPZCjZJy5MZqm
DlJzqMe115iLKxI09kHJ+hhsRUqUnOo8rV4lGUPnAUxmuXXEJsDtJv4K485FDm6B
lHOk5/n6surChK0upSRTshsmRtom9PYCudM/hXZ2z2SCw4p4aQiaM5obWnJJfmRf
sqi/4zvo7ZV8LDwrnTxYryI8FPblPEKkh4ul6BCEeEimWu6C/5vZ32qhYDdSnK2D
TE1/96gSXZUYqaOQ163290zurw9nfnq2+5Ex52hS12theqnMeB9tC4772DsyJ/O+
g1KzU4lrQ8nu++1Sp8I2IAPdY+w/u+2i5Kc/ErRqyAdfoagkFEw/9/Wqjajarh3R
nyEJnDCfg+hsMW9jXOQh2DATHcbd1Lu2BtVoeQkxGqDxA0ikASPBFWf6pCbwNTEm
TwmEXCAy3Raj6+MWl4HCEORHTbYmk8AnyheXUbcDo/s9PUCYWkxxdWNEDttbXm0n
DSSCp89NZCaO7lo6YsTLjn8t9SB3z9MD7q48BmabA6Ri1/sfnGmnohMEIE3dMstK
QOay5Hg770Nx2y/3+0tT0WnTs8lfwh9w1DGdr2BPsEBjCzOG4FnJamQEk9FfGRWr
h9IBsz60N/hi5bCSe6MYN9TuZ5HZHwwyhJyoPd4qyzGnD10RDdG9t+8u75dWlmOA
qVHNUtE0Ztn2rcl8Ttl//KJTnVMGlPX6TSm0HR+KMSy9DV9AvttKqQ4sIdgKfYqc
23R6demmQ29KTFt5DuNXmonkZ3vtPEP1qqkk9iBBWlzc6/aHqsv/0cdKeXKQ9UVR
fRCEjxBlApduycrX+qUxn2KZklnOJXvB8G01XPTnLVA6opEh9/tDmaYFhHWSL2Na
3C8qtDXKCTNWNjtFKoiyBOnp+NviMPfy14wV/EGRUtshQEDAIo+rbKGXuNebAJ01
p9C+N/Vtb8BanJ3ZtI100GgBxQfDGYP7NEhfn/vcxT/g5zG8ek1Jm2YCEKrM8PTm
h7m9aQFG3Gs8BaRNZHYgbDkCbAIE1Pi6G6j3moMtq89CDkAaOKFa38+n12OkELjk
AIdvLwWMQL/nQ8YVutCYmPORlEKNo9u6WrVyGRw9gOsvpyUORtrk7aUc0nIHihqr
nxLj9OOWHpYQUbNa7wm+XxR/ctxhjDozfXlFd3idNdRoyhNnwM9L/W4Eon99GV5Z
bMIL3vaTgWpJZWrZ/3x1Hnzg4AlHW7dXbg13ia7FpB/gkd/miNctFF/J0z5z+Kjb
L8zlVQor7gdXZBf5iJeYlBTaNuhOooERgI6O9hLED+LE9jg06WbnN7Z0MUtPYGTB
RD7ZYrEQ7BPRxemOQaFrOtLeseiB2ad0kd4Rht1GHW5EeVOXyp2nFYAd+gsiuGfP
IEwtRI25K1/n9ULZytTp5fHxyJSeqMNFVfiHHtBfPqxdvIBgE5Zy9yw96qkCk1bO
SBX6l7/jFgiAfpyjaI5rwpVVv4OqtB8N8w6AqtN+SacopzX5mQy1CvBGJegQMGtu
mmd/VcLGdO52zh2GbqK7EL4BQga5W2cW8/ysJLHDkBwsyPCGAeBtlvFFt+jvYpcE
sRFb4BgGd4NshTBJ3Wl+e8GMBa588qHWC5741zjoy9nQQJcl02srr19RDZISfm/A
PQi8+h9eLzoBX7BPvKB3eWqUTjoI4m1UxaDpOVd+18JuQmKHBzHWDo6SuAkEw+x9
/0Bec9my6E9Ss3VZndM9VWiW8WdAIW8Ji8nl7ZbGK2WhuaTomG2F+bNa0E+N4Vmb
5E9J9LGyhZD7tKCHl9YKJlaToqku9rg4fli3I49n8TjBjIL76vT6lu1rSPzKf+up
WfhgPra2cADIKAiZaN+ChYrzZWTgqfa3OXpZl/fKq1l8QIhowAvsd6MeXTClukEj
gIRcqcxHB6wM7rb/V9dHkmOar64/g3OjrxMWhZ3V2bHdX6LscBsfOX0eXifyy3lU
Pl9MuK8Kxr073KtPKd9LLdqA1VSnY27ye48lKFtrg1KbLBuu0nMHEzkGFLuT3RGl
+BKzQsgbeyLI4i1Ysopv1pkM6YJVYBsYJ+DDkRp7k88nIfobjVKzjPspBAelBZSc
fu4fn7CVbEwlXJQXiASFxPRE4yf9uzZXopmBkkQVyrYapa9zT0QxXaVFLOkfIBKM
0sy226Z1ve97ZmrncJwi9PLmt47XPQ27Tze0hEvAVObOusiLvhzSkPV17olQb/96
VH0bYPSm+7Lkl0F0RERQJoGSFZBSEyZWAJZ74IdfKV3b1mnnyQiF+kpqJOykyD7r
kUDWufPhHcLTSoXyJjkmIEOEoZ4NvYrPwG78hig1wOdacY+3x25zJY0h2EJKeTEt
gzdVPU7L2NGscC4nBSh7Pl/yC+5L6edBl3FH/v5Yt+QjhtR1fyoWr3bC1c2H7YOK
H09cFu7pyCOjv72FtrRae+uhdXj40nOnPA1IW3YuImNZcEB55mNDXgJc+zSwIs5M
3mN4/VTx5G9YGdz4AhTjoVfy2oFpJGaYK8EOpBIrAPTDktOUzMUuKorc6ljvOH1t
R5TAMhPnj47jXxlyMJvqmDaifStawFgnCy9iON5ve/If1seh2fK3dPBaJxI9TQqD
d9WOnaWbOrZwA6DHOcr4vGrmETCh0Bkt3qJBkcgl2cILG6Kf6Ijwq6Rnnj98XcBy
D6D/n3JMtTzuz/JMQjOVPf7j1fasxgCTpXtG7t6K02lu0JjqU2Kx5La09Ujbwavw
ZCXWJSXowURWU+bp1/9CRSNKakcn+5TTClchXPAGmEpM0yrULIrmlVH7MF11JLED
ZROj3fcwPEnKx8xdTAhP19yo579WvAO2XcF/cL6/Bw5tc3GvnXogZkeoiroadhsc
Hv459N8x8ls22GUwLDr2KRdIbbH0sVBgiRFN1zi/3VFZYqqdHJliX8XurzNLy5RD
emh55pbWpwgD9tg8HESAgb+jJXTWyeA6P3ryW/sMnw9eoUn/krvsrsJ7iexMOFi0
uHZxkkR67yB8iNRZbpnUrO62UYgm5L46c270njuhiFfFd9XNVBZeYyUbBOm1/2KZ
rEz8xsmCZtpB75tcKNnoCrU6ARZDqsRn6Gkz+O5RxamFL24ASNnYyONgHB0JSO7P
mjMAOZOPkcH8mX4pr0r+y+f6mm2GWnBBQ/LKL4Xg3Gggo+Ho2Al0Ddl2qgIb2m42
0juOZsqiunWA3jCC/OpwY9ucfQ7hgk/JtDnvGvD4ahVdNBJmdDu1LnLE9bPQn6Mn
4IMjBoFf2zDbpqvZJUVJ9JrI3bzAWsrhAj8w2xSw8we3hXIQdNpy1Y0GfHvRYqTt
8y7+9erXHGwPJzFq0fsaSw7QHi7bMUN5zsJKS8/We1vN1806FlbtfAangbDaZLKG
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cZIMhNN+uFfjSLYMi9PYwnbEM6Mnpj3DrCUv3SIVKuYXpVY4zIYojojDv3FHa9GD
dBwy2EdR3EXdHx2mVPQqJC/KiWt+Jnu+z1fZns/l7C2jiLjsvO2Kkg01QNOvajsG
66JtJWs3LAZjtt8urp9ZTnkX0S78xRW23XnV3He9FfLdIlMdBv08Yjqf9QA54fUc
qHujs3v3r6vHH8pVIJJb1DtsjJgnBu+wuSHF9yhGuhE3goW2L6KlvrRbtboxj0vu
xFQ/wuMJ+fv+bIwoBri8NMhcYMl2BXrkkPB7kmcYXIUpSB48vrZs5flPUnuxXYQW
jGNXvWj0Z+DCaoacD84zXQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5664 )
`pragma protect data_block
CjxPcnGKKHswukttjcq3dOMxwX8c7d4/fZnuNp1nfITXWt5GrSp9dWIWGNSjFEBj
xpdXnnGPoNlaoA8Y5aH0FqEg5Jj+yxqQuIioEnb5XmiEDK7krZHKBQeM/Xx6PWg6
zSVgdEbvmRP6ML5a4tb344PmaLYveO30yYDBPVJqbAcjBlvdhYBoggHNIzLh5KRs
/+8U5f8gSLxtlMGlVqfjgQ1pZ564O8JGI4YZhV/JRph1pn0A0PLvaG2eR6/D60Ha
L1whlrUWEEhE5Pxsrf1vBNyA++iFpBQLXxGKS1jHotlNBoU+ovtmGwV8jhnreGlK
MK/XZUf5qXNO5MbA3NrjwlmX5dL/BMe8uko+k71oBEFJGwX1c1VMjqR5Bk44elqn
bhOO8k+OCXURTDg4QYPe55E6P/sfQg3tnS51gHD2L20Tp77gtY+9ZSpk4ZoRthkl
/QILE9J2krCdzq0O8FMOBsQYRFBMKOXKMEbUJBZpNfYRbB+TlXeWOExL0pr2uKmm
IHU32+XC20RcYqWAPqUd6P3lFQZp5/KQ/n1bkeLZ+Dhzy3TFtTrcTKojeqZcRhOQ
F7hblgX4+/20fc77ppMN/rk0mUgxhIWo/+yFPe7rXjbS3DJVjt1yJJImXftGVl0E
IPzUJUCEmiAF+rsXMQJVf/8PApotsTU0M2zIAUu+ViGYREutVCUahX6slrWAgHq/
pPjdicHLm4XHC/po5Rc3Zm48vnuBbD50ykdLGYHkAxBY1hBeF2rO7CBUfGSWFy7L
QK87+dmxd+lfG58gJRuq2LQLcEhWxBHWlIgYqX7pXDGvz7ZmCJV5LJXuVCUwQXyG
QQ40OkLiPSjMEIh7+egwQ3qAZepjtHjrTHbDFBDiLF9H2bTaqKh/ZMuNrPhl7kG+
MH2kLb4cwoWs1ElvtWBnm0c7QjnnEQ2WtqjQDRRcEmnQH96boqpwRJPiQu3pqHRQ
McleTNzePQiwcDh1nIO/SfvDogoyqZ9gSV2SXXEsuRR+lXkPlP0ZKBUWmZcVURfJ
nL1sZIkH6v1/DotX0H8ITm2DAz2HJgIb06ktxz4pPe+8seGMRRP6deyblx/UcO5V
J8lUGBk2OL82t+Ns3Qta5iGi+5qRvgg75iyJ/6me40XCBZiMOLhWdA5btnj0DLfb
ocs/h49voTXfGAlM6BvK3q0Bi34wQvu1zL6FA1nBKX25uJIr6UdrIBZTL69gpMMn
UtRVo+JUE8OeyF2Mb+REx8KWcng+rcXZhYx0SFnCZgBKVNlaUPNJMFVGQu3rSlh0
dwD4lfiYeu6ql0BX6pIHikkNrpQ2QPqktOzfA2AgRWJ8L20mHNlhRJm0MUbvFO5A
KRQLTz+I9k8kp3KEVDtnPssOe5/cQh2lpFEf6PPuHheDl28eHS/tJWdi1UKlrwqw
V9t45kYSUnXx1hqcb7UHMcIqyh2/Fx1QqBam/yClpB4Uwj+3YwPAtKWqbd9Sx2pY
T6b8TUucYm50+GQ9TWoYuk96+EURvfxsUU7Xcbrk97U10V55nHD3vWMU8wO4ASAH
7Gx4ADe+Bb7JmvbrmDmrzmFpeAYK1WgCCEqsrtEqX3mwnNzvGKMr1GZvXt97etUB
hBUm9lsgWFk5mDEaSkTOQ9JtmsEkOiQmPNPBTXBpo3YnRJPlouoYKGKI3uT5ZwDo
ofShUVw5UXCOfrIwPuJbB66JcOosnkMbKUZv4vDR7gEakRAg8UV9TeRmWTOsxyW1
D0u0iT8ygdeTZM+t1+tt6RvmCMSR6j5C7328gmnx6YnRPG/eUl4TeRKT/C4GGFA4
k2aQJQ/BLF9Q7JpW/NCFswiuA5W4gjZEPX8lPrMWE2jo9IIFh91e7m9wIMu3TmU5
8U21Mn1z4VMr2BxiMA8DcZhKJsyqkw2m36kOHwABS8GBnltzVOpAckXv+oa4ek9z
ABwpyXMFqWR/19LULH72wKpiVovL7VPArpKCJO9DW6pHGISkV+NJvgDsJi9M0yas
1PLvczPyrzZgK5qIQrh7dn0H9G8PbDgAV3AD7Yjg/838GBxY/2BnHsPv5Z6++AWf
wyd3KTncYyAhIYGxmFCDa5BlPfc8FsUAkMCXDnkFD7ig+CmhBKvPqw7NmC+OMhF7
oXspoYET+/sPrZxEupIAZRo55L/cAD+/6sdIwVtTzEXd7qpiPZUfWOg0FY7l8PtH
3pUK3jYavCq0tdc3F61Q0WaVcryKU7xFSj6QxezSO7OalAHUItEeHeCijum10Rkd
xIzHw6q8ipTiHP5FyEgGlxVIKhV8rypyDnfcBiIROSToQxIOzzYIknb+hnkhJDTF
wIhzNNd5oOvc4OxmRAtsS6R8MuLS3GJYXhtKUEqiQcVcz+JI7tq+uUTlx7wieaM4
tyGONUSK5v/0ozg+WkpP3StfDXzH2+lB0twfiUf1T/DujglyCJCxsc5uEJmSYNIW
Fis8Uts4RpJvLDKa1nHJNH7wRTG54ueFOUVNqXOK8l2N4bCET0UyUW52BrDkcnU6
hktlSU+D4V/n0NIBkh2SWs7FG8vS8p4gF0ct05yBxQ3jKF6BS9hufCJX2Pudmsoc
ZIPZxAA7N50WLib2ZIJeCC3C16cH9uf2USM8bY4oHgfyf4UtPDN4gLO9jEzaEz2n
vTCYp3IOSX2S7OClG68NN1bbiCVhA0hztkP9xJkehpvDMNg7wIRtcSHggDiPvhL3
bFXrkDJBNNtsiR97o9DnGS25cG025aKufD30eP8+g/sIp8qO8bZrcoux8h5d6izu
em5qi8yNg3UsOGaRZB9LwD3bOzABqjP9uNRiNvMmbwQQJ+9kq/9HfBpIxfxTQSXF
drgpbLOiu0IpvybdeO4qRGg+R79YRU9xBV6ZqYTKNgclM+AllEz/yhmYGu6OyyW1
joYhbj2DZFvJ4Rd3UfNwrWJ1gR5uNvU8H3vr9/ALNhDRWH4FVegUaoWrZJT7PH4o
N2zCSRhNAP5uVSMfomHbB7eteKEDsUf2UGigpjBGIJ8oUPGHILI9KXPshlOKAfBP
XpWpKmHIrKtXYg7lLASFPcwWQjnhrXhtahzs5AeQG2+CmvE82kmUi4kpYTn+D8kN
OU6VGYtPAHMMJH/1o8voVJ61XWcSXN0/pX9Cv2Sd69WAOjZdwoaDQG6Y9gjluQvi
uC9J01gEjHSIP0X2Ibj0ah4KZ2jNGc15pqA1ji0MPpyU/YEOzm/2AEqKQ1BWAiWy
EKUTXv11tu8QZAZaeX3FxQm2Abk6FhjBUlfgt9+Kr/MLDjrjz89SjWzqi73hvxhy
xlYKiE8YOuebm6IMewIBJd/j4yUFpq25G492Vd1gncI5WlOlHT5ONg2csUTULFXO
ONVqvfU8Gc99N0aeY370ECJsZVKOX01GMBKP6BP1doq0+GQxxPYKHbArVzCmZLet
j1OyZQ5ZIBf10t/z7pqetATCh/UcplaZLu4XCeimxmKvZN+RYGMXz8IKcAlR9Ao3
GY9hRIXoCXY3ySI0VpqCJOWi+amIVHClBvyvG12QY1iwBX7YswNUHaynE6x2DIiz
qB5280moLaj+nBGCAO0DrHeXL6hEcMso4Ni8xa4aZMcU5WVrJ7ClgoJ7EAQBA0I+
g59KUTKqqMMAJmkAp77FSnb6DseTumeT0HFzYL9aM6lsLxXdA+6JYQY1lkdyPy77
ncE/QKNx7zu6E0aqDLlQ5Iip6wgWEOtNArJUS3kOP20y2vJBi8tDlc2DOcA5FOMF
NxElLY/fyAzbU263n+Yag/kG25AZEUGSnM0SzOzZgEuqbxPfl9QxYW2U5UQzSGcd
VIE54fKOQVZ/v5X0oZvY88+YsfzrwY9V88814atj4Ni+0LWV+rXHKmdY7pPhkQAy
hYY0+R5jRfFoSJjsXSDVVMd7zjh6Za7frxtpxjyuNUdrb2LFwQU4KWb/j3s2KCcI
nmkJwOhem7OBNDxbVYKyVb+q0X/S/5m1DtoceFwM/JpAayjjwFzd+60Q4+R9nyYn
spv/wri+GdEZk7vdidih8kkiXSmpqCOEJZAHrcr25CWs207B1IvkutsqvJ5dYaGz
sHEll+qJWBDfZEepQYMEzJlA1Y4js1cQmeCe8Si8WAuawRhkDuSKUQtIWmulqEgN
7i0LsBCVjZFEWugGYgU1ikc65CkeyAf40do5uxF54ibmoHdlfmWsVKxO6Bp9v1Sm
jd6RAGJsAErOndexk2xnnewnqx/J2ipb40IVe315MDmXDTCJSro7DOjM2kIxtBMx
zMaAf5mU707GJ+XJL8mzOnaap2D8gV+WBzJa2q19+E0sv1PWIf1RGJoHAWFcqcZj
pHFGIBn2XyuY9S8G8fFqucVYVLMaP4+DUtWE5al5bvVSML2x2HDDbAtnByO4M4Rv
fUXAQBxg6PyKSNfh9JJRK4GGjGrGeJNAHqfM1sedobs+6D6nJ3sgD6njM5fAT75M
k7yliUyj/Vo1NQoHye0ew1pDUJHW7qGAVaVT5S9ZOXX/K/O24R1DYinxW6ZQy1Cy
M+4NYmNAje6AGYIoyUOZQE0+GpxsPDDHFJtK6qZaVnq72HsHlppPJCPvXx2/tFbN
qbKYE5eUkwnERTz2TaNWTnFBVh+twMhvClXSh/3DWW+t3MmxdT02F5w2wK4cf3go
y2wXzXjNHI+ukjYDnZqEtahiwHLPgPdcmMlTUkxwarBFRrfPe/TkzlliFsE0XViM
osEvcFFgcVkmS0S0h6uH3bhm5PN2xloUWTQH+p0UF/ki/Zw461EDKT9QwNjtn3eS
HiDZgwXobjpBGJwT4qtY3qmm8Z9WsxDOsRxG0d0d0EdRO0KqiVN/Gt9XPBTs57jp
SHh4V0VWZ35AjILcsv4As1534of6uIuneOXlDHA0NtLMmpWtXqf84LJg3lQNV1jX
Z4wqxXuR83xtwv8pyBCrPuXfchI/8HLiReg/ahCZCGWlWhtEvaozV8xyh/M+me6n
tGXVddHBDq+REQwWb4zq/r4xovfuf1+60aQxSLk47/js03261E1sBcCzF8s8+FLA
dTI7jMalt7iUhwqAjvYGtVMTPE4BqVF+UBr76W3rqkROfFRP3N8nwKSYsOXByZe3
Gr/nEOY6PhN3PNGN+nsEoNAfRw11TU/zBnHmkHvxtv2I59XEYp8zMSFGJ+dokeny
b9jZ8rsonKBOUXqetPOFr5iO+d2GgITp1w3+ffPhIuavr3Jtd48oLjtYn5e8K8q0
xxPXeTPtXQH54HcCDCRZcfW+mmZPyeAmnhqHkyD7fAe9GD5moJTnLMNu4aOPmY5L
wWJIfQPu2nMyqktBVisHsGF+8LinyFE86s5yZx+yQvKqFeoIzwIcOy53vl478cls
TYNQaavRH3YZwl6e4tr5fisOR3GC49hzWqsWodGOZJ3kKgAP8UQPqcCJwjRjacRD
7C9UOH9Z2I95bOtcvRAgQJcA9owMQPiT7QlyI1JdqjKvyyE2KfF+2FYS7WX9xDON
Antbi8KxvSoSV+pkuMvfUdvmq0RN5l8ovAHMqLD4m0HRUKyWAlJ1jaxM9ttqLFDB
RruYtb3BtMaglNocf7m3zPjltdt7ApwrquMlein2g93qHNaVANlUP0Hu13LcPdP+
8Km5qEviivlLT+MQOm/OF7PMSMi63adD+vK6qtJK40BtNInK5SjLZctGg3cFixN7
hrt50ew7jJ0DraiOsp1wAHQ6biAhs8lT8BBLvImuCju+TId4QLaAsrubevYEUb8M
662MdNG6fHQ3BL/ZSnOPG0dSSlLLPweqE3gn/Utuwz0EQ3C/XKPQ/zTl6u6q2Z/4
CNyPCjDzRlRSMuhOgryHs+x3eoy4UdjZ9qXtgcB8eAuw/gjZvtQT8uDyDO80UpW6
xUJFaNysTxS7MZ+jF2PpMtjqvYlAn62wT4KndiPqxKynxSkl6dHPHzr4fF55a3WO
3Arjxl+cyoZDt3d6/xgX6DP533LZhoLU+ksG7Sp7T3r+y4rQtO+psqYVvnk9UrOS
N+bRblKF1AkVa08dmVY4oapbwEGJ38e0ciaVoQA8VOMjZlin17oK1eeq9S/sQ+I7
XIF0ScBZ/hAnp6UlIXapPinBJqIdD2t+9Wh086UV16ypEdw0Ye4yDUnpZtISzSMl
Os1REEs6J37aMe3HmpFfCxjHXqIg2YTebMw7X6qpsAMbi2a5Tuikkak4MSPaU+fm
26zBq4xmj0N2WuLA3GwkflQbu75mB5jacllT0uXD2OjsZMIdR6CyQAdWoKrST5H3
7XDvs0I5e7s86hI/ivLJTf/Jo+iJFL2Zw0FW/bkSgi4/1mbIwsDsi9xA9k0mVR/W
+oD7oThpSZ7LjK637x73nfRKUk7HzhYG6IHQEbGCp8iq3G1e/m2qVe3eS81eb3Fh
p6PHYj43ZtkOfpvejQlaFeuYqde/RfLwO6nfMoNUdhidR29KdKeeWCQlUMSod/vg
rKc9C5crWwWe5aIEFZnoaAZKERt/OcHEPgBjvCYDura0hfshbWJZrDJLDRT/l+T2
B17dCjazgZA1Eq9hPhcCmMkx7VoCSP4iWofFZHcl4ySendKgPdaISF2HMMxx7Irz
SLEZK7OGOi5Sb0mQ1YugAcbCYmWVgQU1lsmjZtgSIive4Fxt7jmj8Td4tkaj98hy
mJPcPjpqjKf020xEXcXpp+o2GSU2q3P/Xf+Az+upIwWCe3eOY9ehsHIfkFicmB9k
wVOeS7JMFqPWWpk3gqj4pJOJxvWo0cgysEMfXqn+lPMyPuK5DIxKLAYpPpCu9UtD
S21zlx/mTXorjIlfTvDykJTSsD40wSZcBt9y2CDg8kAshu6l1TUfcapi7y29/EvB
0sIxokMScnqVnTNLdWpKsyWc/CKIe1EJSHkx86/Dh3V/t8V4y9xqBRDieBgCSVwV
bOcErdJemjLC8W6gOTVQZ6vvBZ1O4PF2T73dUsdX4BDadbfiSVdE1Q3OPgD2b8Tt
ireAwK7xuXb5gTOAJGuKGmv8qd+eldvrwPXAqLzlyHbysbVrGIxvBSPCijZVnKio
IMaN4UMf31t4Aruy2QhrnhmMPucmZIL81sSc1prWPcF0MhdxcYf/Z2CembCo5j7Z
TVmm/ml0kfsMp1FxvAMZQHONdzUeaIrmefhInew6hr+A97kckpHrB9e5MmDg2JqA
D/IHfFQQeQis3pcLWvHrM//ojpjvtaqQu/e3H7UP9rfF9eLWumUrtcc3I2p14xZ9
JhG53Oh7qpoI33FiBjGV1obK/Ea3IzdicbsRVnVdKdTbqVeRHlr1Iy/hLQSn8+1l
zlC0AW8guO6JSZ+3vI3A6mCnyglU+OGFk8CtTMDUuFYHihphHtFzkNoV0gsvZ4Pz
qKhvTZvSG/cO5OIEVV4mIHW3XCzq6wBOvS0KMvHQtqz1KSDdb3u91KO2ax39Q2cL
8Swg/0n+5Brz+qDwuSaN0paYywyqQdz7s8jdluXsYHNtoYL6oZ0ybSzYKrXiBQIg
tScIC5F/Mm5g0pza+MG8AUtZlhUi8sWDhtSAPB/mr6B77a1bYZKlAd7G/sCttnB2
QIryDdhY2iNeIvfJdVAO6oVJdksL1FZ4KFOD2lYrp9Tn92YRYymI5EFZApbxKSxc
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GydtFHT1GkAG5jAtz83uEh3JPK9+0uYaKnBEcUizkQtbrSrpJxHt6UJVirWj9v5O
85BR74uD11paClQY++CzxJPB8Wk2V4JjDCHsc+RTZOaK2MDBqck26rToY6oFvXIJ
fDaayVz4/L/tvUnVTwBVgtcfIWBbUG9FK8iC21udW28gPNEqfNdesG5xjzmOuMvB
78+z9FLPBEZ6ACNSAb3CuMnQvhTyRzxglFrSUggVOaF1hmAvRQQDgDDKzXuAaLp8
EK0afjsDwVRxKVyQtHyXLYh32gu6/NNDtbor7uzjpl81iS6vxUZSy2mRhWmk4Fdc
HOL0aDKTADg038ZmzmbfJA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4720 )
`pragma protect data_block
BsDJoK1qEDOpsJGTw5UjLhsrlYw8GBdvDehQCDfCd8o2CnrgZNe0jDTZ7WwaQ5b5
yUxs6vKvCWcLfNMdCF6FUhNXPADufuTRR0Lt3Q/euRZ+KNRRIq3PiLcbc/eXbRTg
Htha6t8OPtdWppV45VbU+HFRlu193cPKXEPibK4CzjK6UPO3EBm1Vko19fVwG2+f
YYoVq/+MpjT5VG8fBOZ/Ltq42nD9Bpv6u6Yw9+pyhE0/ICQK2ViyIjBN1WgKXSOI
D7rJfBNym2et5SWBBM4H9wg9h/L899vN2Dfbq9NVL13zOH+Jo0hoOfHZ+nm/9H2e
z0Iec+s/L2xYwYbzGY9raSRHgzfaxf7kK559cQ1hZ2zyP8DelxKhfKL8+nKhq9B1
5lgIU7ZD+t8weaOO7Q5HE1nma9qGch5YxIFO/M3lHc5biRoqqbtVebv82ygB6YcG
PwqT2D9kBk4wN8gl2oYmqMbK62JozHvrkU3ijAIEM6yvSDmRsxYg1FkNjo3R5aZU
F0r2L3370vfM2BIrOWDplso+z6DXrEYNrxXIissGepn8IKUSif5v/aDrilbYNvM2
tVqBLUyvgcg7WbnzLGUPw1HYKsAhrQI+4kORX3sywZ0ha7AicfMd2HQlv8QM8YuV
PAmRo3uutNE9jTHeQWFVWqVnQXGWoaYIMm4EBSfhA4H3Y3VV2QLD2zR1z/sq55o3
cdV6kF72j+KlIf3I4v7EHCoD1bAfNczGSimj3uDSfiKX0MFLlZAhhll9Wuol4RTi
glC79rK1XPMddUdBZXI4lZwMFjsIaR41EsVFneGwz46rbprK89GTwTVu7og6Np9o
O05M7g4IbOiN+sNcIDptM5g06Vsi+JudCWvzjnojL6O0yDCHxdaytzpdKQdid6DR
qz9oGORfgwbc3JirfgxrzkmOLHOaG7iZRspRGcCpXLf3h+N8RD8dhjlfBa3cOzK3
iEQZJvDI7lj2/5+Hf7TKYzVrIPOqXNz8nGvsCHttHlrYW1s3ngeatV2cv/rfU+FS
cYDq4pkrzltJW+ZXzVW6so1JEWhw+pccwFuZ3ElaoTnrj9fFyVacNP2CdBvqev6X
fRYNZzhhY1Y1uFiM11b+U6MWe0wICxQbHiifht1yNcP/dxhk8ACV4dr+eMg2JNHH
8yHimVDEliEQKEc3FkKNOHQf0FLsLrOdrP20ePhEGhQTw3f7nPEnAsxC8Y623MWo
7ZUgSykXUBMgrF2dgIP5PBEbiPDzF7JFML4MXYq/jphAa6ToGuXPpepnCWP4eKGC
rae2MUC3YJLcFvnNisiG+qcVMFt+pGjtCKOdnnfmfQcvd6FTwKpLWiBEUH2Q0PEQ
8K5lRe0h/ITohLR23lEEPlTkwXlv0wLlx12yiWHYe9lnTaOxpByKSj/cA7C2+bpc
Xw7Tjr1nC6XylSGtBpVbyA2f1OETQ9RKmEPgAkekaISd7DrRE70rxFaSNdDL3Tug
JYsX6PM2B9ipuPcSasTQJBFdLzsvhhtzNd20tJuJF3EyD+qY9NLWSyjh9LVAevv+
U7CR+jectrNLtCPoakh80f8I4MiMEAiSgTwEJ0O5IBm78xXJdx+eOsM+SqMnHFyz
dVw+58E9U89MwRR2rfuPtF6lcqGYfxX79R8RbDBJ7rMYqHH76kgu/xiE4a6/oQ4Q
cXeEocHs/cKz7w36ygSh+v2LOCJIk2A4Y8mvsVE5MmcC80cah2ufp93lB9XZGF2E
QWDqcjyawmZdG5SVQKqKFIe9MJLe8kCXjHBHlwHhyGAfr0fi61Z8PbLR8B+6np90
I83s15wFsboDJcF3yjusmd+0+Urmi1TQAHTvIA9ixmWR0dURPdD8AcicNnWRJCS4
xAcqv3KBan3Gghi5hFSwR6WvPtE2oSKP2WxIh1UXCXlxBZp3A9owFM/8kKkQIVOh
eBprg0ez3H/yRiAVOkcReV9s0PeRG+LPptDJivNJTtFBD4D+5f0oh7EjPO05v2ve
oKHf3Tfoqz+pm9HntsWQts+gBhqVa5XEibD7ca6dbF1tz1lYnkFAWu2BznwmPggd
GgKgzH8QkMzf5ICkO2lP3gVzn7/tL2a6f9/DatOB3xqPFzUyBHgG/q1YDmzVKK9C
7RDuLsJT9gcIWy6aVYl8hQ7Oyp5BB/L/UCb5Uom/ZxIR5OWFQpIIdbdFIfJ6jamu
8vdxbuXkw0fPZUoib2neGzRjypUr2f3JhhcYRez7g9qHgdzLH0nvy1uj5Fz/INP4
HKMs0av/IdQZJOp7z7yZ2aGdAl9ebZ/fRRnTI90+5xqIAuFO53SGPrHplQZnA8fc
O5EOF2R9OLpPCppEc03wq1CGEpSjnqcPAyFeh0XkcfAtDlNf6Pmp7nvYpKwnOsUe
F1Aer737TmeiW077ObvKxf3IObyojYu3BsmmREjS3/QPQhgrW97fKI0rzu2lapI6
u4IoeTN6LUCnKHQeYMWAAG5hlv/a5AtbVKHrm39p53x16xZMimaTib8QCUm6c+AU
yp7dw0CPdsElPvxMtl8JO7A+F0uhu0SfoSTqUjs2UcF22TFuXjJzimpB4gFFauKr
91g9Vi2dwQV+kEpAaQ/QR8zschfEGHYSAp9nIOWwZp2suj9NX3Sssepw4x1vQg6w
7YKPxc32JH4AsaWDJ0YY/Y32Vi76CPHK6/r7s59hnREkA46UCwBPtphBOLNNLfO5
EsGD30hExGW7Iv582xhEioNcVerANoilJHRZS8QbIWl9BxflE3vDTm35OUiZkJ2L
DCUG/aQAT2m2tChED8gQvBUmS2V5OC75Kj+g+ttksaZtnjEWoN8FNeATGQQgZK7h
BAYTBZTdk38ZLkows87lEPP6slwuEaE6iyT/KkAQx8BhacabC57Qs05k/IDur7dD
kv05R1/d7Q5vZEWnpGMQ3H6aZ5sLOgMG1xAczlZdDL3vw++cCpcRpONlKuF+T7Qg
mZ5Bxl91DLgU33qGng7uAXCs2Qy+iCH/wA7XcgfQSA0NTnWrrI3zD+djAtRFEfIY
OVmlRPCD8Oncz+y8td0CN0aSiA9UAQ002ivt5EuPqZBqXSxnTkzHgsi965I9KWDz
f9tfj8ZB1sUpFmLG/CjRJ08KfqlYKNBO4MVyhf0pKU4yOWStWEAwWBJL9D3NWnAD
TnWUs+wO9Z6i7G8oXycE3OAf8UNdB1tWTTB1vNJvuHB1xUsjorsgyWXvjSqRah2b
7uYNlCNYiliIOFdJ83b2fe3Zo5xXSZI7F1xGloCSV26C6f7pMSETewxTIvTJBYMo
7Ajj+0tc3t64psvTAEs3bJQFugdqTdcnXow/XJ6tduLBm836YMZHXoSHgFoz+pds
pKZeigeVSmFO4oqYY9j8BqYGKxOY3wwjNWE++E9TYFhmWxM1MThGqf5wIrAtiwle
QlRIMhTLi7kFSi/8kpdPEPCg7iyZVRP4aj3oEL/BgTxBQEBsg/LbcXiN/KjRyXSt
X1pe7YyF8/n1JGO0nTF9r/+e/THueI1C5ed8oI25dfaKNY7WXkMGEJFrkV2bhahC
CFz4LJoXBZIUCafI/5EBe+f14QMzqtw+BWqCphZVk/bv6pq68xiijv1Z5OcB1bDp
HXMAMguhnZY5Utb7lDaiXoDWFEPyrCQpMusFxoJSZrONqeISp5QnaVnVPJ/cOQZi
RDlaMySrZ6+dGliQcdzcEY+F0PG0UAQRIMzbODEHhYl9lJM28tdCl/IAZ3EReejY
KWhJPYwfOAJFGJYk9g21eX9zcQ4g6eP6doIiP02KJJclngi0ieYfc8fkRjSptyP7
udlfiHirgStmNAlryTpstUaKkdoTMuuMkRuqPLHUq7BMXXHUQ12NagxPMQsBP1ru
WiAJVYwgcnkFZhJ8AfHDRyi8fkYg8Al8PxWt4ynpVV1On1AYWfuNWGrXuoADxSz2
0ssJsL4XPb1EsSd76SL6QVepOCk1E3N6dtaEjIC28unLqPKx6TmU9yxgmCNB60Xg
R+jBAkDGZNgxwZxJJ99VNwhRsP2vDGo4YszsqBenW0SvMkGQPAgNBQtmhpVi2lX9
Mt9Ec5393Uewa7mWvzusSyIRvTVIul9MQ5Rir8aj8igTUrU2v/N3YCHZVCMRxZ5t
4oofOX1ncmyNzv2BRnZPutv3EVz2mlXsGTbSl9okEeJrunZmQ/zjfmDpJE5ggK/R
XQPLOIcrZxjEEye86KlfDrfrnN6Me3QLDBiFUHGye4i+6+oO6zEamcYdU12gPWoT
cLmkHN1/3H6A5lFa9Sqk0Wek5ajKVGybI8t7XZKgS8F7Lo/B7iezD94vjHtI93q/
d3IgkCXGpPWbfrjfFSu89ybcJp2EmB1fsPX/WEjz3iryvkztvDrtgvhZ0ikMzPqS
YZ9DlaoQGxUawKwJ2wFhKZlMnhZKFgXHRGjs2GXNpCRcFIgRsslIp4S1OiFiehnD
rQQUBT2/qYDzqSOi3Z1nnSlH6hnJLBncOwrB3J/X7/RW/4FDAwQBOjmt+PAfJ0dE
deLgyRi5wdL7HMu0Rn62ROm11CDVZCnjy8yxm/bVzkAls4cjqdoDJOKguKayerAs
cDBCYomQwUkmp7/qzLjvdb+kh9QHuTPey4rq2NYDVkOOFy80eTLXUWfiAN9eYLy+
kU7p2MElu/t28jA/GLPaI4/6gviIUSoAJp0t2nfLaIAn1Cv/eEMiOfr6EvDAaxap
uWK64EaRy1W5lXXhz6G6cmr4WZMemPu/KVDEK2GW3uatg36EojIk/PGGzfJkO42l
LyGBw8ln3TUx6i4eUSBHuURv8sGtj1cSfERgc59x9b1or37VxFPUJElLmCejtrNG
wpyqVE5I/nuzBiUkqiAW3TX5luZKDA8LFHAQwrLRPyDQgdYNZeuzrW1lJ3SWgyDD
y6ZI45Hr6rorx7C9QxtdabcvLKCx/q6ze2Sf8CarM2u6XD3S9WufCqRezSQEmrT0
QA2lNEtLBdPc8EF59mvAn/7iQ7FCaWXw0DbkzuDSvWxU21RX0PjVUa2fjKES2qKd
zxKHfY2yRRjdzeZGlZ46PVj1g6PDTMuwkK/sBGTHxDLtEjbJ4tLHymxQ1qs2WUvK
Rc2mJ72hSQZDv7psOYNEYl6fLyd2DVelFs9oL421cEo/XfIEsbkt1hIfBocX9XDB
09gsfBWj6qYcgpUkQtkbFVKOBskBbZDGQzsWEVwkZRVtrIlkaL4/1fhrsbRR1AYG
m+NdJKE+dsefFHVrDjng5iuGccDiVEOoqprK67p8zDo00qh03UNpZ5cajiynJYWa
xKRHY8clCXNMzWqwAnTwpmuZzg3kF+pS3MCdo92ANce35LjAn+X8PW0VOut4r5FI
Y1ZV7gthJ0LzeLdwjSm+9ZR7KwAUpKvUw3Ddja8GGZgbkn8eJFzOHqAcWCaRdUyv
MWyTav/Uq30Ht8AWIGR+6uVAOoNNedljzeBA3bAaQHhXkiywuFowwv6zsmZzJxnY
n+rQ4e7+Uv298pp51u+v1w4Sh71Ln0+3TrrrdbixzMM4BeTGMIrivglnU/l+tbfw
Rl3H94XeszFxcfQzZv6/maFd9wTMY5rSwKbRbPd6lKP4DEs6IKRmymNQW+lfnqUv
wKk+iAwXyxP1qQ3oJSwS4D4/+8qJbQfxTPCvR4G6M3D6XMVdC3/eBqBNTNP4qFij
Hq/bPNPijTOY8guFcsKu/hHmRDKat8/ejKBkR9ijiMg28UezZwqd2EMSPNYRfRPm
Nx+/n+DXzuZOGtx3wLQMrnOJPpFGGMiZ12d98QwBW9DzY1df2FoOdIwphKs5uaTa
ccY4K/Yd5Y3uQIIbfnLBs5kJebMmubusXJr11nSm/KKW+NOYjGXGcWJpYhb4N4Uj
v+u2tJtRZvrMld5D+1VW5M4blznnayvr8ek0RgNmhXQOwWmq6Hpe1pOnUpQJXbvj
ov/ZNB1Z+qUVj4vd4weWz6E3XBc2Zhcc4rTgSTUINMJvv0GWw+t5CDu9eWNo+Sjq
/z4PItKv0Ssc3lSKFv2qUbHEZmXDwvVvOp73mwHhD17HwC9zckctoVqj0bDOJbns
oYUCOHhgwsUj2tTHaTp9Uy08xuQhg+GOLxMUJRHarKPIGD0f1g9gSyIuUb5kxgK/
6bjUNvQsNj8OJ1dhgiXeHOJ3r7859zQRLheNiArFB5C4ib7vSaSiL9lOMsPJx76t
Y4FpUqWPkBTFofpFFsyJWZcxohZHhzhLAL5l2ILsoYVb2eSCujgtdUp7MY3bZF7w
Mc7awQCnusgIANNWp11USmsaXP32pwpY/d4FIiDji9RppbcgwyobViZpVyPFwrZF
jLeKLTri8P4bQMSongO+lg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dKpcnnhgesCnhr9IxjHvEEtCZU3fpAxXK60xamk1OwCxZDQSFRqTiLZs5xBrOIdC
HXg9UyqXXMhK+asbETzY4v/yx9qZmrIXo89/v1UBQwGVidJQRzoTfyFG4aSeIuRP
gJmPMPHphz8A/JQhkGXNV5LCsPErbd06E0WOtZb0KwQrLdQ2ffwZJ3iefej6Iyxv
Ld702MAArvCfNtM25+PeHs8k3NoTOdGbqPTEH1nIZDswPYmBDp6/sW9xobfN+dLs
YbAt26FMtOyy8hbNS73zVnsg2p311zs4KwIpOB2pIfPlAvsG0FBLFvGTgYPnlfvP
6+4VOFh/SyfxH5FFwfwwmQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4288 )
`pragma protect data_block
G3Pb4/tvWluCo2omPxHZ9mZDd5Udpb5AHS1/gU6im0sT5dOram6Eb6QnyBSy/GZL
bKypu0GwTkby18SZsu9sbiycJdJmxf6YQh9Fx+OY3/u2OHfDSPM7/xa5NbSa1e0K
2mStnP2f4R2Of6cTUg74HlYnOip+f14qXdiE94m4t94ai8PMcfst1NZ2iIDtpCxI
f0HWE9XRfiriHNFXfxzo77cKuaAo4a0zrpfHa+yiGAPSKK6CRzDmtRGV9uE+Q2Ob
yZW8RODgbTpt1tiGkS6MzwMa4LC5q4jBxdach0xiGP+puSD7SSPtKGyciv9AX/XN
0xo2mBU4fBetAM3Q+hr4Kl3ssiGQG8dYODvn7R7P72qdx0KXKFaufe+V1gEhOmnT
84BAsukHoBIYRe8pmEpu4CsVzZ69PQV4GyBXpJOcUD5Fe2dKuEjrkD6LlIS9PTAv
IIl++487mQZUqWTGLeO7vNlXY9l7cpMl7QIlO+1K04pVlsDT628o1GhjXGX7Ox4o
8bCnLRS4MQgzil1w1/hwNpkYHHv5j3gE93hUKI2/07+S9gNtIuaAObFrxki/NP4Z
ZZC2HN+Len8iL+5Ge/bbh349sdStspSRWu9nZGKUGpjGG9dcaGBtzuQ9/Y8z/B8M
TVEDeRKua3n1mtD4oNtpNQizXKfxA6RL9R2PoxFUYwsME03LX/lI433yk2o/3cyH
PQEXsrHtUgC0cs/wlPt0eha3/JRsUcjdKzfBCsxNlYaQH2HBRW7erHQGldIMZCj9
aaToLac9SaJhPDJ4ZRB0VVWmDMht6v1LNuJ2BRzxENw58an5PC6jtgOSJ8nw6hsz
OInTI7/kYzPG6rWUudAK31tcI1J4S+5gOdyN2CztfqxthdMD/F/fPzmIkJmr+i4M
OZSNs9kco8TrpaRM2enNrUBA8wiFeqJQVmOEqQC9DlFC23RPqy1fOBh90ZM1jsGb
0nsx/qIp7rIiPrRFdHTQvQ4Vw+KR/I99nHmckUSKYoTkvUkbiF/UwXAA/k17wEf5
ISREy82yxPo9oUmEtVBriysCPr+L3ff9NV4jtUeOB0GD2BbRqL3nEPiLH5Vktmlr
2ANaznyJQnjZxhB0q9zPBwTGxlzm4M5pPbKy9bu7a5ERSMET13ksuOP3rtlOl0zO
UQCpArsQOiAqPF7QoavevnsN3wi+E3AjsT/QcCiqiwogoxtPszwUbyuPQheAsdh/
7YZIuqicafjGkJggPCJ+2XmxqKrIUjPiL1cIE756NmXDjDPf5g512tA0ysD7mmk0
DU7WHLSXjDCIZ7l4f/mXP7qxJMwruQbS0nYXhdJpZ4D8mY1i4MJlor5vwYbOovVl
/CyOVmqcPKgFXh89wo3n++0gF0L35xWuS1Nt0PXVEeY1XATgmdYXJBKaoV4+jNBE
nnKTMsO+pyTH798umXsged0pYwN2HdDpFUHMWDFsAN7MFu9dGa0C8LcBa4clzSKS
WXYR6OgT7N0FSKiSd/ITzaYhbQAWqkh7HoEjd6kViFZaO9qPtzkN4yYelZ3NzoAa
pyfTGb5h5QZ+8vIfJeYqdQ43MmuA5felzQKArLPqq26hNrKfWsPEKdj/u4ac4pYP
ofoDOtOdTEFOB1cJ0w/kJkg2ozpnDNv4OfcziF0p0CN2lqXP3dRhVJNDyb5yT8Bn
33mAb9OzEwKxGtha0zUlvn6jxTsmdWkpZy9Axud3qGPFEggfxs5DuFEfqXXgrMyJ
hWhfpV0fL16bzHqFpVhyoNZXxo8xeuxqQK0dh8Ne5MWfgVWuarUX3Hyw26cmIqSU
TJa+4gB/xGUMv4wOE7FOtgZQeKcUta5MAiXjFPIqP3LTbEmtp3se1CdR20HncHJH
aiW4eRrgiQ0DeHwsdFdJkCx2co93CrpuJX1BStStv89kqB9x3f33R59JhSgDQHfv
4f9X7ryAGOqfW9J3Ge95ZZPd38Hi/Bv0iXNhx5EDQUMvXyyruJLMRQsNt69Mhcwy
NBeMEEh+8jqj3DMaoDg9TlGpv+lUsnYmNv8DMLsjqku9QKiW51tJRnERjfYcMDpi
WN/OgNoAl6xujEkr1s8+Ei+D9xNrAK+1w4Q4x9U8Tf8HkMao3lPA0zY8doO+WZou
9pcaasL5rdfvfXZAS4pZECb2K1J19ZYBrjiH5T+f+yEXEM6mS3M28zOatpWx10uZ
x2a12sQYA8dASxrjL4pMY/QtVWsdOc+y4012M6QqZ5wwlOeFRJTcFoYGEh2vZO/N
z/p7ihsM3PNN5xW7cXHwF4ZOP0KFXOeefX28Yjls4bYjD3G9A1Yu75x42dJXrGpz
B2C9FCJGyQrvzZo0dUBOHprEccW1E8kD1EZIObiOpHJgOTueZa2rh2SfnatGdV0K
oJbzCstTP2SmtqryTp/4oNp5t/vTuG+5LV6ppMbFOKor43KkxPzuiHAKm2FB+ktX
BsyPatWMsIizn4p08levaNAXr+5klrNj+RE2kwyW2Z9UOIpTb7p7i66v3Yo6jggK
qSczY1I0jemfFcTdS0dlcRK7cia9/5tssvNU2RAoT+O/GCXn7t/IC2DwAc5M+9vi
F6SU75hX5z4CQC6IHmei5+Jy6FxOY6Y3DwP/N/aPQq/9Ng5GDqOoW6yEYzj21nQ5
aTcokTq0FEhcdWIImrFZr6cQycETXXo3DOQ/OKueTZ7ffPBGyTziBVrdzPY9tGLH
K8O7UOsMmOtsBP5aOuYKCcsfd7EPMcT0ZXcds9PMr/w0CyNzJvMc7aF1u0d6MO5I
NPAJB1HS1sNHTd9v3RUY13d93fv++cnVXvbAHyQZog/iZX3pp0BTOt6Bhw8TtR8i
xb2lVWURRpmTr36A0Q7VVd+NjSyrzNj9vIE/dTIDmaRZBel1TlWdOIGzzVZ2ZITU
N1rK6OLzYh4uq/jy1HjbKGGXqNoto044whFGYjSWAv3732H7i86pM7m4ZCFFdKHX
uxN+Uk0VV+nxVndbpSxLHBtqyAvizMY08kzRtmRnn44FBVNEjip2jcZlUzJlqSTj
RcnWWGxU1uBA+0oG8bQYo2NyWBsVmSrRpSMvfkSZh1A07AQfPDZpUVT8FY0+8ruv
qFBCvpOfrU7y0HRAmX6od4j2QgljxfKWir3DuT6Wm7SHmmF73HHYQSuPWw9KHmPd
gyBnJXZUVbRmN+xq6y6PL8okROYR/pmMHt9MjZ9+16MIxYxl28MLPrgnszIyIXMH
vGqJ2WdibFdcsQewsLci2LNdqPf40fZusLKacF1D8twFGTtX2Ztrp5yqqJ+cXMgL
UGPdWsH8zMq6Mvv6knVgD7z3S+W9TT1HUSmIGds7v6AbOIilAqM2/6dg4L18aFkQ
WbZE33OtrJGsSm6ktiuLeqfxk95ZDskSLzQNfo4NCuKAxVLc2VBJhSS1XtZ6x3/h
P/NmwxfeC+oiOyoRSJppZeBGK+/nQWwUZXnze6L2LMsGJvY/HpGGCF5+BnyyEUWq
ikfo+mHbLjoLTMAC9NGIV7fcB4JcDcaevVHcq009Q0yvupFzMAPYdg8ApOS8iwwW
UG5rBsxLwz0pCGjUcZ9AN5vnh5u38ML4d0UDNiKZBc946/dW0h7AiVy7uQvQBMMW
gehQ7alIGCt5HDz+7oaEieTfxoJjMZW2tu0enC2TSBKu0tNdkpyjDHVc6sxPSoXt
T8UerArf8YFwzvUfPVKhwRM2mucX3BEdLhbB/VHUZB4PZckoGEtRupQgKznpCpXy
c/+4zCzt7dhqekk55F/riEh/bajYJ1qiri2MU0sl8LHM8eupacDn2XyYD3zQ4HGn
qVlzFxqR+zrj3LGD1QzqalSc1gPsB2X1sYqfDfalTBdSMCVMCx6Zk2jEnB8NGO5O
Ob8byapPFbKCxMBlzaDj6RC6zk4y8wrROxvnSjS7CmgYWBA46GiqkSV5Zs/7SOoe
DVLRDqhvutz7BTUckqcDIoZpvLuPth61ly+kUxu7GBSONooyuYIinjuakZStRJ1b
vjlT70f0BJby1Lf7rrQ9bYs0a1elsNvD41Ja83Zsr/Ra6/QBKWE1WAS8WDXsGhiK
DyBFM1YDwpGw5wLzDwWGgo3hDn7N70Z+Mad6SLKqYv4gycI56vjkbFE47PjRF+iv
jIwgmrYZEpDzLce1tO0OLMVmY2BxsxY1jvBusfRlAsbG0Ft9wHHpFr63xPmSnTDE
TQp4M8xtFieM59hlKjqLdKFHemXFpsoMF97fgrQ05NjZ5cu7if0njW3AmyoNo4+j
yM8QZzR4IwUgla6pSH1vBdMJ4gTneCgPBRfasLrq4xmG94Uvsy9MUz1uJUEFNVVE
CEz0lfMjXtZJqLjmgsjTEtP2/5UvpjWvR95pU4bvn0zmUVWnvXOHEqfHD7LcLpJh
6GYIbyWLr9e1toDxTcCRLpXVjLwuxNBMLskpXysq3J9gbt7bOUbZYDTuzd7Np41z
vNJqNRg5OBS5iFTTRBFt+Q5/7x7ug0/Rskuy6Z+TBl4H52/xGxpyyJR+perMsj18
IXb43bL6PXQdWZnLr4Ac8ivcYqSFBVlVi+kMHBF3w2jnW5dvzciJpX3BKjqUMvPw
8QcFkoF+77tuzGUHo2xoik//l4qcMO3s+WJA5XybrW57M5yMhui+doj7hcmJ9XpQ
0ghXPAvr5AQY8FGK/yrjJdS6vuogMMjIe0a26Eto/dIFJaRv1a2CJadAfhGX6jtn
PiqpSqn9QfwGfWq4eqq1UIbxymhWXvGI+qOgX3dVdzA5cWFHuigN+BbIGcYgkXZr
uh7NuDv0tiJWyvrUgk8socj8EsVRCq8BxW+9peTuONQyvdLLYDY4zPAovPRbBADp
UKmH9lq7seTeTNPJ2LuNg5GBQoSIihmiw+c/VcP9Q4JBDR2e57CFoL3vrEB5PIk/
Vyw8gTrCplpkOZg91RSvsOEPF81N4rmGTY4M7/JJiqoTtWeFHvHdd6ct11pJqy46
WcFLb6LT7IGkIwA7oyhAwle6Fp1XxVoDXSQGFNYaoCiuk5AaahBNIWv5e7w3KmG4
W65UQS2SiHMdA85BXpjnPksrD1I5/R4o7ri2siLDqD8u7dWeWwrkYs4mRACJ+mM1
8+WLK+ywjj0kaq6Y4rhJtJ/x22+nzckKqnZJ6xp7wzHlk8jSZV/lvlptj6quI5JJ
1w5jRblr4PiWNf4JK6pTZUWQXmJ12rp7yNEpJRhCJKNBca9ZSLgdE5iIvlbybNl7
NfUeoAjsvUMkNO8WeRY9bZ6oVsr+pijDjEBlVu/NbzQiq//62hhopTgYwiHSnFgA
x46QqXjHdwKIQuVlVf0IBCfqzKmXHJcH5ddvacQrlRj8faA9ZcIag0Q4JEfuS3oR
Cj9a1f46yfZC6WSQnLaoAzAO1GD0IkFhJIkgda8nIPXSo8H/DeZRSm9edbZ0ukVZ
3kZukpo8jcE42vS+H9S4HBniWQtTAmLe9nft1xXzz7udcAaigNoWg6Zy/Z+01OfG
wcCu95PHkpGojj5ILwHnteZNNNHpsM47yFYpIJl7RrQBTyl8roJo1atFLiR+fYBq
B++IXhVLU9m9ZjVexausIVHfQ2gH/p2qgfl+TBOMZhba810PFDpxJRLz6H6d75TU
JHgBskdm0UZ8WkAyMkPtjREt7EATFN5A4HacohaBbCZw8vmB4CRmdkq1mIKNNcTF
Cs43fcDMs+br/JiVbI56JEN0dnlxHLPDzZchG1JzUmoMD4dFQNq9FWNGtIjlUUnR
BgUj8TPLLKRGzHNGYpRoEA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
N4GOveMNwzH+hSdTVBUFGOBpWwQhOLmgf7L9F0Uh+gFKiT8G2Fj61NgofyOzQm0D
b9rJ0fFAfab3C/yLhFBxkVx04K0xrEShutbSA7FwnrNCviGKvdy45hHNdlCmIbQk
f8CGAOjaez0T+rgZ8e5PrvfZiSnAXHCUYU9gdMfEilwQeoouQL4cep3A0tXBeut/
8hwZgb8RNB+LNPWRu9vZZ2LPmFQeICkxfiDPe+yNj+GqMb4KlQFa9n9Lfx8Xknnt
tz3soVq3oWGbICFDKeWkAhCFJCzs5sjcd5f1zBgZP8SwlZ7eRh+Zbf6T/mmWnH3c
j9ulkR+UnEcZSTM6HDLJKw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
gy48xJooNTa4x/uQl+ZUiv5wg+tHlWBYcnHoAN83sCdXsi+MGUqxu7MPPBwQL6IJ
e6B78VRkkNfRFP6ZXa8RD/lLVQox33DBtGxY0FxnKbiBGm+/PHCIDumWuW4eCkK/
iLQZLgb11Yrgfoya0ZOYnIC4rYeSqzjdkR1JzPF9GWqiDHOyLRfsC/keKbXGo+7E
9aCQOH6wMrgEFrUKvwX75B5HLptnNTNmgS65hpj6DIKElUiwsw63ceypNspiZDOL
iYFakbdNENMYDYQiF/CsgpR6XP6QwPuarfPnkQLOFO+K7VuJRmRLzT3X/LofkKfI
UxZp5LdT+o7EnEenVXA4CZ3fZa2HG+OOrtgEg5HByBXFOiyhEg2d5lIo/GM4K9mw
5sqTY58lf7O3rWm9xMODK+sXW3VwLBUZw9B1cKOji2o0aI6DUgK02el3T43qSJL7
SSQqKT2u0CY1aRVAlOW+bTmlrat8GaQ7l9S96vgI3RTK23S5kzH9hvrbWtQBArWK
Cfz8AlhkRcdnnSDDkAIodp/Ewhi4g5QkULuvHHy+XSveyIiTwEVAWAU+vkSegtyE
bGhGQK+PfpcCaDzbwHRplSv6Qcz9Xyrvi19e1c1PXQ5Q1p5276aYlX6v1TOPOV3G
ieuY1JBZmmDXXEwXlKyM0YfIP8T7rHoNmEKrFDEcz8R+7CoE8H57yZHNonupGP9L
iUPiOazI6JtMEYqtt8fa+79uu9COBgT6Tsnc8FFGYReULsq+LwIOvrJuUt0gc9VN
vSwTY/9pVI4YkpUvcmqmQIi8rin4g4y0hksMeDQnhJDTHAM31mx5x8zmKETgPdRc
42q9DwiVxFRfC/VRYkwF/DWsaomQU/LojBCOf9Dz4eUeOSl3Yqaw7EwM5sTm1bG8
JBoYLBbb8qGqv+s7jrUAmoEdrOuRwmrSQO4LH+1zEPg+6CaW6l47ZTgZWNgvwkJM
tnrJB2aM+7Z5D4jEflqkiT4GiKX2kDBA9yfCgaUQbyNbUCzXX6h8Jbo8q3xdxqmQ
VvJvtGhl0g2SNZ3jHkJr9ZccFk51lAjIsIXkDl2FPhq0eACd2xkAbXtUYdRX1fq3
Qo3Cy35GZ50ZaXY3JTMTw5ve7BJ+RSgnHHT4ZplDDY83dbhod2+Sn5idEN97tX9r
sZP2MnDgAoD3jjaFazJaOfWBn+ktMqEjbUy7gA1UHyUTdsdgYggwCRo3MBc/sD3m
k97Z/iXZ/9gSBOYAh8Ncl81I2m9lE/XDrY159UPN7zKuhlxNKzwqRWXeNT8lz2I7
RE0KJl8kfAx7uwMrJBdZF/hm7M00gvTjDjoXUHujPI2vqU5CAAmgEsdCPxRDHlTr
rF4Hunb+PrNxmciQNTdiUBLlr9kewCwUSgTLmEb8gdZYVG4YdpBvC565Z+Xr2j3y
l+fiTmp9MVOMEOViFZPicSPQkwIiCfERAMN9j9NLQYw/2AN68lx+TNTbk/j0qF6y
hHcuRAFpKTGOqS9SPzv1QX4MWgDTznqGnqUgwCNcEFMsSD+7Juz0IbOjq8OHP196
LhSlpfE6QmWHhjQtxTS6NigdkDI8uDTGhIZndD3NnlRWEawtsjJecAFzoBF0OgxY
qR1dpEBpkJnAjAyB3UJW+0RJXSbou8twJAmQF2FpXi0FTXBhO8PumQZL4iO9Z2sm
5mCgdbcrTjGzmI3ESPWoDBZJC9NtfdZpzyDgxFHmDeZF5HaTusfX3Xem1OGeXErA
o+wI8Ha+ajjc8q6IuXWyz4oD0+jwSHb28ajV5cx+JIe2K8GQffOBwJooGplWsFaL
TUn4g0opGwJ5KvHoprZMvRh+JCRfKmXX4UOZABva+BZIj3kAPFDtRnaZXsA0WOAc
j/S8ymOkeHdmhNmaR62vLSW7C3OWb9cRRZs4tMcz6QZqle8ZPTLF7Wk7rL9JYNix
9uspQG1LVlC5nCjJ9vV/+dqYFLaEqsrUwlPKU7JFXj7oujl0319OzH2OU/i3kQc/
ag9g0PBYzWeARSxN7edss1b8DLHBFxCheyFRog9rgNi/qXIR2SsDiA4GNo/bgiLD
kSWA732FFClB1zcgYwa1jz0HGAYPiDpFj41RWn+YWYRaAgwtd9if6UEbRFn63gl5
JYTHZqgUZb5gz868CDv4f0eJ+LyZzTorIWtQFfd/XAvsYDKy3aUTcizN3rK/dy/c
uc246jdFSmmqXQsQX62T/y/mt3FqSS7I57gay0i30vUwISwh4B+yK3q15qvcpLys
QgndLPeOHFWHA2ON+c9QI6tD9VFSIjh/obA/IcZcTY2dvxNVmHp6hdhJMrCBjHps
6cBPcmHha++UZG1ENHWUVc0QPaHs2R9egdcfh1qTflv41dGPJOPliVvQQoF9l3/y
f0osy5wfY5PvMlWAsqaRySSEUKoNRf2Ws49ubZ+xXkgDWlMJHU2ek5iEDStXx/Gs
D8zAQG+mD1tuW/Hw7H1ILkAcXJNQYD2vL3dh5XfNcCh+4oqFkimE+WoAwne0Kd2e
59k3f0ryVl+4SfvueSQRojarwUYweaXk4u4Kb/lfDGr9qBQMC1uGaMY4BrwGD0v0
9tDm5jsdXmveVtqiXfCb9rFxotH52wcII4iV6ELKRxbq9W7tQUwkBFXnl/cjmPbT
5y1Z0gAj1vKCQ4oMZ5cZD6uBWtlEN217Mu+b1Msrf3WA751Rfbf+S+zzNc/331Ng
PtaJ3DL7ICrl0Up6M90dgmDZXyX9qgjS1u1Sl1ULRKQmcmW5J5RGJQJ8r7ab4WZs
ostu8wkFMx2brqMuISMZbS8+vd3HviVhfFmHrkUS7v6pS+NwSe3f5UWIxHxu7RGk
BAzs4NJjVQH7wIGFTxUWEfeIpmgs1UOd1Y1P320tt5M6gbJjHgZQJcli6N0O0MJ+
uHHEzKk6X9EfMzLaWkBkoeqU49Zb+z65EyB/45PcafwoficSZV44i/HAhugqQ5RO
RNcE9SUGWj2Ti2yQ6wAVWziGTmYHwl8qog+8Y4ux9rToGNVPHc4bHU7qLf3EwCLW
AjQXMAJ6jARTt38FZ3jD9CKsfokkcPPS1+MYKK8YVX21NVfYzwMzvYoWKWkJTnK4
tFa3ZrjeJTCddikAo2g83hG0B+qbuwIoN3clxBDSOQVTS7IZQSzPT8+v3MOJsSpb
hWipGvwMaVrkT5e3pkjph5Tk+Z6/o8/GGNFVZuNXQUQ9Gi45u5YwXZ0qfOR/7tMG
cvZPjyToG0xgqHZeb+Prdyz0dOegxqBut5NdwvnUwRonz0QF0H4zr34/yH/Qg8jk
2eJONWbErOJlQWD4awDXK+hUYRRVk0JG08Q7eI97YDlPvvqfzG717BJK/eze0U5X
9pkdm8VmOdSJ81Rb66Jax9YjMSxS+vC9raIqoc8ez7RE14k6lu5mdgr8YEPw/XYN
eneJkRIfTtW/3her4sAzmsTeB00736boLKOtMq4XXi21OPNu0QOZz+lk4s9PE3xb
SKYVXJqynrnJkOiYHVYntuSoFIW9MChxFkrtEU5p2PCLtvoQunLVYNjC6CKxFdzB
+qVoePwjJjaS8CxoEarha3nxUVZ/SLIEf8x//7AGQ+EQmji3vsEl4RXjZmgXZrwZ
sivNW3KCTQgU7iaVVhPhogwytnLbefGcmj+44iSLidgeHUHVDEHFKCehbOicAmjD
m1s7LyhUoKU+G0z4AY1uLetgbUdL31YbTWybpO8D7KCqtsNeRto4gLNPSBlUS5oz
v2iG2tACJ53/dEMDPeCVdwKT0pzxeMSOzMwnAJ8DPp1dShD39hBbojGur1jNYNed
x9dOfTVzDaFHe6Jufxe7MXLZ8VPyrrSwFsVZOaXE04KQh/N0x1tcdzav/+9TMgZh
zR0BehUtswsK4r9iRM2fx3UVXRC+6JP96chxgXpTpVn+nm7GTtfePChMalwv8L4s
fBsXko2S4bTQYGnZ8DWAICFqmwstfBZnDqpHXf/0hv8dAH0+Sux/PrLQ9pSyA4XL
ALbSTbsxCN10NPV95ogvP+7iBmHawG/jUTl8fERJWh3Mm8nehJx6NOgx42NWO9HF
Kn2x053jyEVgd6G5IASx12CJOJsS+uovGA41sd3NdD7atEBIbyUA8iIhDlYQo2W+
Wc2qgDl1ddAp92h2n0Mq8K0+IzamD6xlOMbYppUW0iUbzKZvR2O51FvXEtVDP5Rr
HzJAKFFHZUuh0a3F0hNJiOadb2Z1+IBnDZr0S5YmffwuwplEA2wnGpbYi4sQHRd/
yndFsXRcCPWaQO0Gq58gPL7EhJbs69bp0XdVEpG3zNzTf+U+JAhaO/VadbFN+CIE
vsR+no6/3BINSnEiub8ZDGPPNDR79s4XQxzsh7WJRsZwzdRqB80o39RG6HgthaqM
0qThPKyKD6XvHq5cPuFf/wwv3DKGfDZ+jA4C6BTscL39OJ0kJf3AE0TMxfdk3y6y
LCBqIeh3Lk0FlANuJ74rUQY9abHElUJS/LsuovIX+XzhjjkXmEuIS/1jysi1abhb
oHPXHafdSjdkjcO0JyP+pDMEgcrXeOEuGIXoPsrcF4Sk1NCXZjRNVvL64FF+suIR
QAvZZ+7gopeFQfhbz0CMSqEthj4XpGjwENoqGt8EGCGskNHVXvRBRZS+PcfAGVGw
7NaczegWFbxyaIwGQPFE4qwZC1u3WRY+/HsRXreLfEbX6TopbvT0aPmKI2RN37pj
T9/aed8waPQ8zwNd7kV9f2sJnBaX2EYngvoYU32RilR2cqy3MuP2l9ZVixxFK/W/
k2Rp5WTx5y/NM54XOpyb+hKuGyKcs4k7GHsUUt+DiHaXxYsVgzXcF0B/2EwobuoT
f/3djLryLEh0XVtVb6rVbuGqZ9+QhNjfTg6vEQjDdzI7Bcpl8X8zYQYZjD5Lnlts
9S8tECpQOqLsOquF6WCtHR9v/l5mqynUEcPGvKrvWtR/IZzxkjomd9U1lyJgbRH0
txPbwohPgRl9a4QUptHTYrScyWRAdXN7cZofuJ78oRnv/yn9sgD6HVwixSwCTD58
mDh02ZVmSOwSPY/tetgaFLvIAhbBT8ga0NLS3pnM7wpl77FxMJCqXkqKj8nZoexK
3clR9n8uVjbdeg1vOYXpTmBsCCC2QEy4x6acq2PomI6hGPdj26GD99B5ZHZCTO6a
zZ2uJq6gNQa4oGI27OMyTDpzcVfqMvR4gek1ynPC1Ss=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
fjfpZveSl22bpM2+CZA4SGhEQwPAuyvyyklIG2Zy52yutdoFvVO0Jva9Ujdhe/ue
Ay8zpnj+q6csfkNaR+dzjocnDjrYvwmqbafp2z02ioB6Y7X6iZbHTVqfPq3d/vVl
NojV5/cmsijUr5MFZvMvb9Uo7M1sNsUUBchRUTjYZmO/mIN9LHQs95gOtD3460KC
NxlWiZ8IKDiMvtSrBqH8Xi6JCyTy6mEn9+FVtyzaOk77FW01qhT6kE8Y3Nb17Zjw
j6AxsBrKDguWikr10ysb8dGU3hSxnkgthZgi6x3N8j5iBjSCjmdnJhtkgntafE+J
E+BW6ozBts/VhyUQAr6aAg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6880 )
`pragma protect data_block
K+8KAG+wpD7Pr7VFV1TAc1Ty2MsKZQxnvrRk+uUo4jpHnEjK5MGB1J79LIkIGlDO
kgsrnXPa0CRS1Ej5O03SVNwVn4ySA5rplAD8ObV6NSRIHgjpFNj4JHG627PLybuV
CiboTI3DpnoSFYM8vXQFNg3dSm1Z7AhZda7bPM26bQvKjw1quuRjDEWzg63IF1iG
tz6fxp13RuazfKrfYMNaOXQI3iQihN4YOtjPDSyp4aGbmoIZfrI66R+d4IMGhbE5
uYhB+6R+Ru7UUqrtfkS9/Wf7ilJK+A8ra+1U4ZNafdFIu6pgiPD41c+i9TX5U8xx
TYUTph2lUs2fAoYwo8vk3RMBo8rbc8qwdLNMhmVsAUrKYpzHt4wXdG91zi9WiOaW
jpn1Gk4J/vjTO/ShG7rohYBbBCsWC1h5kVj3UtJe3grIzFsu2puWFob9j/4+z1uf
8u+mpAXoS4K186EdbO/1yv7cx8sw32MejgAi+pC5r2H6G6MMmiLeiAGQaJhykocG
kNOHNV78+X8uQO7XCjLu8e0Pcfq3RHtmNOK5HNUHWJB7ckB63XLwEN44R/FJnJZt
WCEyXO9p7G2+foZ7euxN5//eJNUr16RkbcL/hsAHmC75ZdzEnEodOaStE3Ty0JlE
EXCRnD4HqSxQJNa3mnXoE1ya+ThIRaf+bYUVzFfdpPLIJQBpAtYJ0+h9wndCM/UE
Y19QQvgSMid6HV6ZgA+vgGrunXTjenVTH5bfLVVeBfejthxMUDgbamYPENcm+xIB
n/cICNgT2KsQ5cWBPJM90C9UlI7nHuZAzpyMnIu+4UjQAvQhekQf1MWV3+RhC1ZI
BW3Iy4js0efnfK4O4c16ZuhGCl3LQEjbsEDDeddfIDILUeVkFkJWMTR8/oPtDMBV
ZMuqn13IRaVh5Wktdnl7kvaW19zfvuvsMcRV/DkOQP0Ede3rk2GT7RfK5X69v+oZ
V/7/n6PfXQ4+Rol+JjJxuarSQ9HsbwLuv3CpR4d3uv4iI7zVEJGwQPfQTzafw3zA
k8vqrSW/nGgi+vr3/QvHUqjIlxbP1U+KafwOp8EfJXxtVFJzK+EAxqZyxDgKLhMj
Al5cPrgR1VYmTOeuFN7SbC8QowBaqR6u4zu2IzHeziluCHTW5IRa0tmfm5I3yky/
bEyNoeexzuKVbE8zjA6FOrb1igdghmHaTainPYh0Qb2qhhscMCt7TM61GvImoFkn
T1/FqWZ/gHcEMJWKH0m5bhBsd6voMxcJ6TXs+fgkSSsgdUWv1PqJRDL0gTQRNoLS
B4DClqcp2kfTE4SDdtkYiFruglFhlCTwsvJjFr8Os2drStT72P2BfKoCs0gaRCpl
iSimUQRPOXpRJkXhI6hX/NWGZEwsSr57hBdoPqvDwgfmyP1qcvVo16H+vifDQWiG
7wGkL03JRBdi7nk5Jfar181uPNCcwRHupvedqOhkYdWJVUdC3iirZodUXiUaC4yC
7xcLJeLgjglNOefFb3rcTbeWjMOIBaxGhAkz7WY7Sy2zpZ4sapbuqUu/EiDeMYy8
Xy8vhcZv/r+L2fXpCHwEIpT10YpE9ZzvCCQefKqpt94c5OsyiS+MWtvIOcZX4j+I
fkcDgvhxZcY7jRFA8ZcdgY3IDojnlQrm2+lvseoEpkA8x6NhvPKX0n+AAiHQG0hT
Ns7pbQY48LtscBy5ySIYRYlp4J4Ob5o47GrpJrHztJ88CAiAINQ4oFYZxrwxTaxh
1Ya/7ArJ3TSr9G1BJpblMhaopb+5y1/NsSTDxYPY6hFs2XdiuT69gIyKUvK0BdQM
eYV/8F+izHvHQ6Cfs2fBoW/Gr7ZIKnatIYC/X/Y1VM0roKoeXPmsDhWvfivWZzsT
zJVp5GJJrUvhMYTbZH7BvANs/H6VHuMig0MpL+Klw+Ktg2pz06wQDumzEU78JM7d
7hTpE0jJ40F8A1cnHnZwWQ4T52xHDSSWe3IKQb+4hPn1BkzzKTvBZ/O+0CwAWKoG
m6jJ0IFMOKCmQxwMlUijJYpJ3e74pXdVtEJeIvlfdjFfCtk7s5ONjcUg4WQ6uozQ
NFl3w8NFcltBBrH2oWzHeRPVZzn0B0a93x6vHK2YsDmuUZ11rGbwMXHv81I1miAD
GpdRq9mzGFlhEImnjkaUmI8xzrHUsFEuevO6oioo0mWxFpm+I5gdGvioJ2bR3ube
caQOdyf9hV1gBMtXQ870mrQo0qkyi34UOPwmVGPZbHsB2AqeqTNof3h3a9vW93j/
ynvabFASGK8TaSn4ydSFyTgLc9oImfare2NSHCioeiBDXM81sdryOxIEqFQp/OKL
12yfZyU+J42SrbN/UcVDRj3N13sRBeSTqkNxFqoT6x8XHsqlY8ftHmFQtgmXFM7X
bZT1SRJl076rG7vD7tIvZcXVYzs/kksDcdgcj78IIERLJJ5O+NvhhJLgyYVeFVxN
N+yXd+ohDeuP30A46E0D6lmTG2Dh7A56Y87oWAoAEvXUXIkTwMHotbn5mxBU2aNo
eHTgkEfjxmCx/V7AXWxV1m+QPpZnUNUngQjSpD0Iza8nDnGekh2AWmi7e93lSgDm
U+OAEByjurEOezhdJw7yZSJzDukBDJ7/AsHpPBSFoq3QPY50t3Zn56ZknZC70nFs
d7g5vZArq9RL/BRYOTqXV3Ywds7+PAZVax8Ec3fN5YxqrPJnnt+RTfUDi/BlBtT+
OZKpAUMiVDDcHD5Xw/dBZ01zHH/pG4TDjbsjJdDMTBNtIqJg39EAo/H7ZwklIm6d
J/ZBecr+1p3GjVmLAQVVAlAc7YLhKWnaUz2NfwbloWFDrKZFv5a9spOYa+BaAU8Y
xpvGJ+3vjyUdU6dKs92LI74sV/BnbugzTYgje1k21Su0LQq2LRqPHSx7PWJ6ZXjc
g1W5xjt9xuSIeld9VGebo3hJ8mSE+42nJezGhqvAQ1SHe2LvA7SZWdnZlsQkM5Yp
8lQ/QVNYBSwDIqQfFUxGzFmckgUjl4meuf5XXQhMD5eyY4K2pyhdnPZNb5EHnp+F
3vhDwM3oAUeNgECTi2/VvTz5FX+PRC8QbSV6eIM4YuxDvkw9/FHJNVeHKOJNZW+y
+Y2i4r/64aHBZ4jYM5h96mxBAgRROB795igKgVLSxIyNYXkpXSq7pbg48G+j318a
lb2fCI81om14NFP6wa95IYTmSC2shkZ45kpr6HRvexDNJkS1oMFmUYJMKj/cO5wN
7tZ/5tpHgmxu7j1DbSLitH3r3lrSY6hGONxb1eaBPzun2AItG6ogFduKIZch+/JE
1f1GvqrQWS5GGxUX5ZMUcUQKPV0wD87HHy/JzKPo3tArgwvpGqlopTs6csLFF5sA
gX9pf+p/nCj6og6ziGlG7xKHZ/ljXWl1PFHyt1+ihSqEcC4B0GYKdpfeJBohHEUe
bBcAGuOkR6cORJwsSyk1pkLeJst4sWHwanAbzDIOnT+7gPdoPLCwrBX6psXKZqiC
7gR0DUVGAIT7YXmXvAR25qTj8bnqYen/a1OmAPWG+26ejbPROrCn5ou14gZsAWyx
5UcU7BeDh4PG/5L43iI6bnLfp72w29PlaEcAZSXBO4zcdslAPMWQAKtD2I38dU4/
Gv4XDov6FsXHpumWgaA+o89B6jeRmY3Gd4snoEyzpuGveV7cJuKK2vFio6RKBSaK
H5B0BOFK3TK1jahmVni9PtRGOkFvLfDeDfSeFaVWPfHR/qNcOsf7DZs5TV1fI58o
aBOkJDndSvRdDJ2Q4zrjB+muT5oYApkpfNCdc+hj5fvPPpJgcd8sYKG4AF6s4Vfw
N5qf3UwWk5sYovc+ciZmLiokqQHiqTB0On5vbcoozm2I0WDmQsH1lj0U/Xx8YdkI
wJnP8VwlPdvlU8D+X55DWKxRN0g/CqepdcIVg26BYIFGjtRNLaiGdQEuaQYe5rxH
xZAdYXLlUNOU1CtKLY5k0myMDhuwPRrZLBQcwnvLasIZ9srjVvnoHa6T1ZlCI0H7
VGASUfkxjbJ1Fg1a2hE02xJ3ZwBnskV/YR7qeJVjbP5xQF5GXMh+8RXeCGg2PAmz
ULnujebf/DuOotGfwMsfHk+pE4MXQfP4iSVmkQcAMJi5YdV6TyABsCA+U2EYzm/M
jykB68jpMTYAGCrONDkSp2iUz1sQnWvBYmVHOxujAC2pW8WYgtKhx8JkP5qQrtgP
wG7qqyBB+S7xdV1ZwFvlzwVm6L1zXatXKz/CSTkoIlpd/jxMX20kaUaGyWddKKjQ
Jyy8wdXIjx95Vxve95vIgInOdt+8SNQZcxliQS9V6aLy3kxA35bqSLXUolDFpSaD
+IR5xt8LU6GOyM9RziWxnRRJ6hEjz8/hPJyM7QLBEtGsawl5zTX1KWo9MKAS7vgl
pn3Y8qKumhTJiUEVkapxghAA+sPqYXnoHFbFlH8U2hQ/XGzs3OEFL/zA4bZ6aWFd
OM420kS79SBHAj3AjMtUbqS143tVC63fbjKBDCHK4iF5LQiIOKU5hW0qPL55cliW
8kKHbHZ/04hKKV4udp3U+c1NtZlz/+4z+l7CouNWxppj584+EKjm8i8Hhxzde4el
Q5KWTXj7A10nuKIcG3QIxsifjf88LE2Ub7nN9Kheqnb9/XniExoTEP8dG+4cCXFO
UBnW/1+mnfYcGhn1hTjmFtzokDWPEIdO3T3BSC3cvVD2eAxCwrYp0nwuUicOgGAG
kbStYnePGlG4zgD9pqAEtZ8NaxmD+gJEgjHHoXK5WgbVyXpVBExzVMNmVtt+19Ez
mqCkkyIx0+w4YKWIQZYgN2Bf5xDoataNwm3i5uQ5gpshXTo/QsjNyDwXoHH4JC/m
wqsxruAbnvLoMUGgnzTzbKEBXkJNI0zyBByF0hEU9Jb3tfh8mzo9ZsRueZllelkp
2rO4svKvpJ19bYOL98DJa4iYaNmYBKvuUIIeNCq5lStBFea+Pc842vpbVlEwIlDg
DvbE1hkSsuzYLqwZRfTyRO+Nhh/leqKJByrJP3XaEAGOkgcGnbwTxBsz1Joa1XU1
e9Bv8xdXyFhALOhULOzTFctcLhvKG7r2WJZuYHVMKY6xIbpMw7mxsxEwhJsTCQ0G
siqW0HaA+RYGLrno4EgtURmR9ROS7CdW0PQlFxwR18jtYwD+1Hoe5dPttmoX0JnU
jACVjwTKczGHB8UiBsmHVzGRv3IzeAPhGQuUyD1gwY4RMukAsQG3OaTOAHjTKw+J
g0wgl9Pquc2iSSbXP/CLmNBB0MnE43jOUJU41mWj7aj/f49RQul14vJleh1fHSvw
hQwbTlLEjQYyAPmVmLtSiKWO3lVvRP0JdEGpilNdFPhmpoEPst5OTdqPSDgq595F
dPSmNW27CSyheMUT8uqpC04XQiw9zNbUn36Yzte4VaKLxh1vhvudj0m4gnpiHIqU
z0Swe151CBXwQmp3eN1/RWBtsGTPeD6HJngzKY+mpKy1fBWfAIF4KKO2NWbP3Y44
73q2SVdzD5+JTAWfZujJDgRELlxLFWaGtrUcAIz2C54GifpjefvjMxx6x6kdwNpD
9UlH7objxJe4e7CNmVREtXwqIkZzofj7XHmL2VwjWoijXKv1QrHY0GgdrWw8zm7i
U62EPEoKCmUXSoxV+n+tL/ZSdlf8ILz94HKoUbi3tW2ncpRiNIuhCa9F8cjSUlEJ
5hhkt7dbVALfzIdTG7W6weqgFvWQqnCDYg34+bvGfpU/SucxK6ttpUevF0T2VNOb
JntpTZzorzEcts2AlIUYBRbNdszJ0ETKPFkYEk/y2K/v43vkNpoi3ygRq7cAPIlz
oJIOIATj0fI2UVlsNuF5nmhYyyRhpfHm45zmlSSWEYf3/Ki4+fbUytZ8QU66fow7
pYN6jiXpNl6Pdq7yA+zG0EXPVon5ruV7V98BCgkM2Hgs68Es8OnQ8w8r6AavTGYp
aVwk7oMdvanNAgl3XysyYRQVU8njjP5CObmHgnpoJpH8vU3RXjmPZd+bSkvBN22Y
C3e4L7uuW/LU2XKgyseIHE3Qdtv5CWeXo5tutzBInIdGsgMVlechZWDRGVMkMNuV
anKRQJhSrI/iKKJfx+zROHmoWUxGKxHAqCfG5ripH882N38wQSV1hz7RCwyXXt+H
jImxcmqhrpa44gIyRvrCf5+hj4ecTNQFc/Y+zk71IVv/Mcs6YzeCD+uLAlitt7l3
t846euHg0kWinPqXZJ+boW8oHnG+GD3DHfEJXAABOGzJyZwdliyZi0PVn3RHH6Uu
+MRjPECReoKfHGVt8QjvwgqOZZybOARTVfAjMVaxKdbN2FGxl7spmtYwhUNw4NIl
Kp4/LhPYn9PSgubaUucDwIIFj1JUx3YNawAYmRp1dPEJA/voeTg34EiTAlSIjQqd
g8YR9FYJFZHy01IZReCXdkRvwk3df62Veghl1U006WbORIqGXbXAGieHxk5tQEVx
cN33Py9ECXD3OiBdRSTP9fntbYCgKOmaqJxeFvXEKrW0ezhse9yGj7FUBFK5LqxD
ENfwJ6dhAhnqipknbXRqMjCKLiefpjB9cV8Ha1WeJhZEftY+/vxrikS0TXzYmNTj
IyZ9PQSSFK8VL8nd7wRdlzRh8eRrP+F1tPuoL7PaB3bRLIZ+t2SDbrXz3HpdIsrn
H477rB9gRM980iF8IUEvIPgRZXkJv7VQ0xNgeWlWAFL1UInWSZiR3GLn/maWdvcm
oetn6VU9+ugetrYl7VF9r2xHMKv/sUdUEDt1VFg07uXjDXhj0YmULuZ3dhBvnXdr
4xh8EzRIGL4ha7v4J33mQ5KiVAZkQWcC7AsREYD+t8w2S1ZlPjEutxHgaGNZObVm
eEoNZS9XQIZlCLHf+MNhbZg+A5BolaVH3GlNKo/TyXBBPIQ3pgnmnkmibgCANCS9
QuNjd7PpcAacq8e/uebfLqcBE8VlEZsm72fiAhHDzR5VULm8NPaf4qBAvPtoBEyk
Px6ZaruV6yNOuTu2GjoX0icUE69qBFhcpLs6PzEGZZvvGsXYf5fNXlc6l9kKNAW6
xCcNgTeduQTRsQDdxQYKR4+tzn5KtXWe3dcsCfsiwjkC9RsWjaH4Dbm1T44kv9QI
R/LuFVfpedJg/0zPTptuvw3QEKTfH9uTmjVx5Q2MUvegyI5mWiiTRA3m5ipwBDR6
RHwTI89a94R60O7QWLeMT1Y+9K4IAvTAxF6nLRAR+2MJW96oRpzHo2m0ca7YuDFs
6Qf1D0jdPUafYyna/fd7oItkXCASSFEn8yHudokPzx6PcNN5IapW2dOdm6yfTHgF
CdaObP3OSFZn6QvTam6S+uG6Sz3xOfdGYLljLmgwDYV5sApJl+mnN8VrEI8v4A6o
mrnS8nDyH2q+I9UlrqqHk1q3jacO/Q0XvY4k5OEEDTWc/KL3K4sNgOBFtCdK4O9I
yWQgsNzSesphVweVJT3+O+VZ+hS9qpECbv3XLVwx5f/AtyY8nbFMxhwGxgR7uWQm
t9x8Jc3DjendNChAldG5LklyraLl1BrvRNdQ8mdFj0zR0SNPTOoodtNy0s6ib2DB
8qKOGMpKytJvx2w00kCeGskMMf4ErA4c7z/lxIGJD5ARBYlnloB6kf0+wWo0f3DW
DktrJGL7RerLJzdMN0lemYn1R5s2ma4u7bB1YgUU+UxXA9rGMBzl7OMk7Q4nYOA0
2rP7DZ/mWEkfRyyGHBpvnS7Z4S0n7y9paxlOZ2K/Uz3GBsFIAPdUS63QWKeQUvw+
L2N9X49WHhkniYAtCB07w15yRKa77oq5QR8+u9+yWc7H4O/TFU8wrwYsKX+rS14u
8rPMtgvAuudfWVZmqrJhUYEpM5XW2HN6U+YA3HMXEK3OvDhPHuKkgcHgsIBAoWgN
UwtXMjLFwjIFXlIaFVosXg2D/+270ymPLRgCH02IzHBJn6UAbn1R20DGp0m3Eoz2
V4xRSuPgMM+VwCY7pCj71cn23SA8DuS8zNVcZiEFOvQm30l9iSa/cuvMhUEok+fX
kQIDde67WZrl6M92B6/faeDllAfaMeJScFvxihdPKY4ZhZtUfoS5Ieb4AB+14ghh
HPT4Gjb8W5UDKYsXXyOP8kCuvLx9QCsmdOJwHmGcY5G9QyQTIU6O/rP2Up3PZdMA
N9Z8RpKP73FoVwY4WD2TpMI9KL6Q9uBnwYoZ8FWD6wIBvOyYYUsr1WYp/T8sOJg3
s7XHixlvAGxOnxt3aqXlB/WawevE9Wta2SrsmEtUjOUl4fiSnkKumwq/a3qAo+m/
/yP3bCgX7QHD3A2mbyQXkR43jd+HLye/mUuNvNw/djcG8An8+MZFwLMKIXTalguA
mG/EDfRhYxq7w8sS7hd59zzmrKJG6xgqOuAE5NUOcWmW+uHlSVUphqEwv/X01QMO
G9PPwFE2mJwSZkX+uUHakCsB1F5PJDjOjf7bwMQbWZeRrUIsoOVSPLs/4zh1G8Qj
GnoOaQQLmoS+MVv8LDQBSBcwflMPvtRZ3h11vMgxkZ/aoo5g2/vRHVJzowqNdUUp
WgG/+QcD5ZkvhFsjeVBHP3PsqdEN3GBEIUqwsaFNflpm61FHPGUuciaFQQ0U27Wc
MDw1/MmTwga9wwKKbgJn5kmEUmv5EvFb/w1ncNx3rv/mlpGX/Z5w5JZORSa5U0nC
wJB3Kl0pOWabAf2ZgVzlCiz6W4vi7UrqSM/EkbIKvNjv7vhcmFK6HJePxp029YGc
EaGcq3APvX4TkxltBLKuCQBgqsnDPut9p+cIvk4CVQdnZHIn+QKIOS9Pgin3mPF/
9qkgQgWJREqwQ9Sni62L8KnhAS3l7iC9JFjutu8nkAcnXyoP0VB3jae1C4bqQ9OJ
XLuhsy4tPGTruq1J/3tfUMrh2H1fXCXjREUKjseNSWdCtJknpWVF1e6x+KHhK4C3
XojMxM6ec+1BWoJ9jRHumYmdvNXTYEWv3JH1ExXJzvzyjfSWFQukvrw42gxp+XxN
6DBmG6cwu+scWrBz8Tkm9VVUPf4q+f7hIfJvjVsvs9zH4GkA63WlXwikaGlsQsrf
62ZVh6eN+9R7AMUDoptvVoa5js+SKwh1DaW9V4p3Kyr2zvELifYLW/qs7Yo2MtUN
g3u9WXTyQL5bT83617zEM3R5uwIrMkJNLg+MlifzChTtr2jW5Mo7Ly9eXy5ur2Gl
4FmhwsjevsLzbZhsiAjVkHwl3EYI/wbmNFT0VVE9BC04voy4VGQU+/i+I+do1OKf
gCDWa3Xq/kXBvcKzizQupw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
R+moTEEYNLesgM2+g4Fdh0RCLx7+ToUJO7OAuHtKBodcqvg6HMVx31gmvfD2CUGZ
OIXm0pF1vK7D9kZm9i4bX8G8HQXzqfdvBEQBFDluVdItkna3hYA8xsVzKX9+9TIo
klzX/DI1vw475RBlZdM7I52Dd/8XR8FAQsPJx44Xt9XKI6aASXadtDxZy2U4cudx
AqVUfHw1klbWx6YuJ+VWvpG6eFolmjpGhP0hQ1yw9HtqrcWcWVZuYyI3XH+rOIft
GdqawWedl3lvmE4whYV7gA/uE5p4e7clZ9On6aE7ejkjF8H23k4ULnoVylEV8jt3
g4sFzYSaYgWifF4pv3Qd+w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4880 )
`pragma protect data_block
Xb3NWJ5HD4r0RYeqGa1gBVWOP/7IiGDlD/+mPJwv/e38nsmSgHXWCO77DwnH/Rw3
+ZcNM7KoHAys+tG8vtusXnmX0x5By8Y8iyPgsQz8ijzzMb3UbEENY38Pq6ds8uaw
zTte3yQItVsGEn20jv48bTg7quuAQvtIxw0zMlsh5m5WBYhJ1ksPi/bqQQFVS+8W
jQwT3MF5a8PybrKQJtrua7D1UTSNddup6t/GjN9PPgOIKVv1A6XEqE/AlrqFnNq0
81AJqHANOgFMzX6BlTG6r6pm2MjhUT7NHWCEyTs1B5hC/Ft2r18noMDg5VQOJ4gG
dFLtB8CKZPEWyixFGzLZFGb1lsU0j70sP2TJlAbW6i/0yqyAYiQQTIxQjOhXxdU8
qX52YE8kry0Av/YF5fw4wgo3AZDwV3o+S2TWqJkoER9hiDd+IpF+4qbagXWY6hLc
w/hF3qp3rbsmSD66m0mdF/UuUqYBz67GcXuKLT55gxgfGfzvAQUrNavbWRKrymPq
Elykh61ephd2mNIVsn4sm/Uot78aCmO0cPkmWVjRYS2Wja0reolY9FzNe4SaEy34
4EYT9kJJm0kqXuc+iqPO3JsRVJ53Lkkeo2jdrcbkzRdwT58gccIiO/KDxM4dbN0I
K/jhekwkqECfdEsQE6nkVAiNgqZLcH/Z3Qy789DUUY5YWSIWFq/2Y3b6ovhfAA1a
UE0/t8Eadj9CdoeofDi+1IVuuqoepYx9x9v2GCDkQqjfdpCcFL40qNnGLlfXq1BG
mUw+Z03zwbErxYkwWHnjt5sv3QvO64lAR0a/WBJnoey9u1P2aTK1PnxiEI0D3lS/
Vo7yCDQQqZDs75NECzI5kY7cq4mdJUZh7QWPwL1GbTz7l2AsweW+X7NPfc/UOF0W
1BtTHPiPW3vn3xYHXYgOTggpLmv/3O3rKZWI/N0MHYsEzW2qhI8BtPzq0kWtg6oe
cRa+NQ1eDJxXzyb4F3sDcr1y6RJtHgEBnq4fzYALo/Nnkux14JMEd87gqrLH3Pyi
4xdkESUeeRJaFDM5l3XGuOuP5OJCqgLLZrJgUCBlbODeo8kX5Z6AKqTVCjG0/tXc
bBSSxv+HPF4cg8/PXwscRUkjQROHTGDI2Zekesr9wJHlIYw5qLInRvhf5fOYiQw3
aacHINixqIHaGv5GY3XEbfm1gEz2/JW+zC5wnFd3vQR9g4q/AQnEAeohWZS6BKyf
MDnVM5dJTBeRSsNdKNjJCclVXHMN86Y7GVnE/kedLZod6H0kgPpbYU6pG4n5Y4U4
OaN4MCigsedQ2369Z6klU7KvqP9hMN9lATUWxUxDtwBxBWYhecVE54Fl0qQzo1LX
DIRckI3VXQpgxExmGOnC0pgNVegSwHOuXQudqSXwaxoecDGQBOfHex+6NwyCn5IV
EHMkI3DgsnnQ6I3Yd0Nmwq2uxywcosdpDjydU/QodK8oZotux68UT9BFqa3FQTuF
dH9jDCLAw1mGtkOSG0j7ab5WPV+vd3rgy81IAdyAN0vlO2//rHBD6tUm3BpruZsV
yIOTdv+AAuonkxhluIYrzQOD/PaamMHYDF9nC9+U7Cnf2+dFcwvhvuZ4m2DMfVE0
/rfptD0CaHberrkBmOPk4VNRPB/j18MxCgE0pls74swctMWm+umaLttCVCQj0BaJ
zFq2X9jUN5jlBecHUSbq5PT1XUjeA3UQfIVLFaeWiRinZ14MsUgBpiUVh61Q83+C
D/KQBCR47IWIsNT928f7UMjyeU17h4bJkNqQ8G9WcpLCfz1lvEPNrSC2dxzzh66m
s+oUS4XUtnrAHHfpaUgA31sjrRDyqojfsNobOG7T007Y1ILB1vzzufnsrmB/7787
7Fi6BM4vpAmtHbKaNcMsJLtNABauKxbktpadzWukqNWWyFdbudF8JnT18QDJZEvs
it0NWqH+nTkWbzhnXstRv9EgzBMJ7WMmfWF01kYePjkmbLpYSdUCfv+Q+NMTPIHK
04Dmf5yfDSWGJySFMlPAOk+92KVdnOewXsvg9iDPAvfav9JjaSWmzBC5D5TwARgS
PsWaPVYDb8wzi3eANPqq/0Rl0F4ucJpzuRORYnXYv5mC9KggMrLkCa4/uDOX7EGe
aqPe8Q/o/U7XV2ffbfdYIMsXA0JIj4+4Dkf46ma5mpNPi4ysJ8lyGEYP5Bs4mss9
WSC3Tk/tOFKP5FdOFBVCG6pW3ryylc7FKTkvuMkY15syjduauqgT73uAKDGDnM/0
AZ4WYn+zawtPLZK1IlmkkZpbJV+mXy2rWDCHJYpgIPSoJ1QnWuz4qC4Vt4S5py10
cZRriioTww+MTlWAc/uadGI99WFyCVkrzn3O9/bLwjVCvAb6f3bGDNgxclovv2Qt
V0r7NVccQ4Mvmyqk63sTZKgXIH2rXzD4x4ecFPV+GPxZvzjZ06Otv5JXJZfg+22/
TUbCPgkd9/txN2B4nR0nf44sopBsi1b0TB1wssv/+LPPlPBnxAcYcAh41zavv5N1
a7KcCtJElxVJm1dEJuBEQdyQVUsg3Z5tj/ZfirmwzCXkudifmbpFvSiLm5lYj7Ux
bjGstv9f5VMz3cPbycoo8CQaPj2mR79A3Qdk3hqoPFujg7mqL4Pyo5rhkiP4qoOC
uf4pByiIdWcVZpgTZFNo0q57PEpwthKoONp3LbRM9YGOG/z93Xnmn0SCkcNZq0jb
UjXkLLCUbD0RGWhKAI7LC99/8RbwlcyKrdYruY41TpEqpB5O0BA1qIgyohomxSm9
eos/7e1tXTzzdodwbdh/wJt32QVy3uxiBAtKe4CqB0Q2pk7pbHF7on2m05cHYU9g
Ld0nM83e8n7utSxjeRDMHXTGcx/zru91evcvcgD905KC0p82yTTG4RI+fgj306BN
Y1MWLDNHhrG5h+bdBfPxsC/R6hCGqG0ZGkNE0ylzqvkkgaarWsSTpMeLYSKYv+EW
SILjltelYDjM5CFyFVs3NsThkTZjFL+5Mj4sl05XaqRf0VfF1N6IB9wTuTigRq4M
hUuTniOqFVDM9q4jei94B86cNAKjw1NQI+90z4IWXuV9LhXhzsdNwBxwRTgJOPkI
k47VnpiJwha2zD2keBCgMWhbpE6RY/ziFeXQogBOM/EDNFwgMs8fOVxOgHVHm8Vg
IzKNANopikGsAK9JQDq0onY9bbWTvvR5CpO2yPN7CojEeYwGvpQcKi2MLCga7zXB
1oOJ3djzikwEfukJ5vo8YvEwZ+QJp+dKM8rGYXbDgD3JI5Tei4w+H8UksBgqAGzT
xFnr1m9bJ21SyrHBlCPHD2JQvVdcEZop4Ye7JzChtjF0EzLFaivilDH3KJdwKjiD
lDg06h6J79+y9pxfiRZI+FjotQv9uVITASkMIZQnly4zPki0b6kpJlF2dynOMIvF
bwllIwOklr8IdidxUC/s/vchepMRC9B93dzaRXQB0yOe2hAxUq01c6wDVenkqg0s
HaQ/WYfmGyPHJ+7zum7O5BNv4mj03BFk6YFdMuroefLxHFLtB6gNXFIPCchL67SD
/bnTCmWUfBZC38Xw1XS0Dwm2usg8ty16CSu7RZzaTeknQLXCoLtNOuovr9s6PtRT
8EoIEwHsqE5lCe9yj95gX/Bj71+JMm/FVOJLncyqTfiEwHHrQdD7N/exrvOptIe5
wL/wqDM8fYBrsHqls8gCrnvQUYH5CzpIb16yd4MYExNLrAiNgET9JpwcwxdkTIi/
oWbzTcRzILfaiN08g2v/PR/MXWVDQs0ETuYgWiCFT63peRDKe2myXef0k0XxbDDb
w211pPKD9Q9Rzvhkwh31Agk29AxpfD9SUTnuMKM5xXaK3jmfsLRYR4UAPX/mqf4C
CnTrrnPWs9ximQcldyUfg9ZK0Ly16iAsL/DM3r2rt2vzK1VEC+JF6UiLolOYzlqj
gEsSEiZMMt9QtyLZqDnVB7kJvWIXhHv67UVG7qtvD1A/bDQYAWr2BYmkte3psaQR
LPn3wcKeAdZ8RL5Na6H8ncDLkdfzALX4zb6xiZ1XaoHA5UIuTnDNNBydGrNiOG5Q
tzl5nZ8MrAnfA5zac4SSNSsNp51I20cPtB5hmllkR0PAAn5toQP4A2S2OUkF3iGw
YVbxTUwpspRWNbXv3nDBNn5MBttSbiupiQFnRxHhQfM3WFBQSGNsdB+ewUePM9VH
f5gsQK1Ln2uIMZfFxB+mrobuIa3cY9n4lXkfmvcBHBYryj2HvOZ7ssSmW69y+wtV
0+riO/TqaC4ZtqKI2R47CCZQpN6ZIsbSkDL1Q52mk4jkGb4B+0LdZIlL7Ar63ZO9
wcpb6r0w/o6vhTGKQwTrsD8mVBRTC6VJ9KmD8lZLca1cb7A7hfDKCX/2B7E6LLOj
1sNMYf4uF1gB7sbXCK6Nlyn2jS+cJpaDV4c4w8TTL/+lGVkk+uQyCRwQd7+jpv+1
Gw7IojT5kESEmKrvF6UCy8J6zy/DTWXP3kOj6yc2pBofQiBFxxbe9adXNeX3ogrH
oKm31O6cFUSIF5vxW6LRy+36/vwiyyNvIrZOGhnfRuZNOgKuPm55JNSWlJJb4Uhm
5crMUY6zWiN4icwhAuR0J3RfxYfrpqCEJWUBOYLylmYOnhStqgYPy4aaw/BhPCZa
gxCtWrBl5/5AcWuFRqvgGREdf6T7BM5yq7+nJanVHjB0Il83bbS/0WznLsNIu+KZ
pFCywcgzssyI/5gXb6buM8M8NZ5bPN/aclaQzD4oroxlp3fSyxoR3fJCX1otDO8/
8vDJly6azEQRUrl1abTgbryBd6r9sPB1WlFVRjGrWQ+kAkRH0g/bD6xXhmeeKoiQ
T/FcorJZviZBX0bjzmC1r0dlx0KT5rAL+Q4Fa4kdyVAxFYnjFivtR0Bv0rz9d/04
C1afdlNIiRndZ+upB40N+Bs+ujKuu7WvBKuUlnNN6FJqskUGtPYgFtd1NxCOlZAC
VHw57YpVX1oqDrncGGEQJLoK9ULw1rDTbz2nM1M/5d7Hv4NvTsWNqXzVvvZxa7aC
SBnEiILgvVHdCe19BTldXhqhnGHjaUuq0vJHnKAN7xuiMt33TEDBR2hWTjM7ZBGI
pFpnRxUt/xlmk+VXB8hEUjS3Q+5yw0yadCuBTK0WpBb0J+Qt5ITJCE5p+GegoVuq
0a7fPIjtnC2uGG7bGLhQTbicvSISldcAHiH9q+Km3e4wLx5IRZ79EzbqWQ8xNIm0
HdOriqGAP3OsvqMByiW/4I5lVML2zT5OCSx1l2pwumcYHj/OcQ1mAvMkqTRU8O+I
sZNwilKweJ5C7FwWdBZSx3KB/PHihem9XughSgDq+dqYQli7JeLP6zugl0t4SIbe
HE8m3NHl9DvvbQRm84AMQaHTLA+2KOIKVPSyopnoC07rTMz1h0TA6j5oFXtydm7e
7A6q8nYmk2YTMhwP6VpUX6MsolPf4zPBmL8ZzBdx1GRqvBQKxbrzCVp00lImOq4h
J6hlr+iL6H7broHv/oqgMsvPyr0cO8otv+aXl8BZQa7uWRnhViA50j30eP6Sv5lp
rdOqIj2VmL2wTUpcONmS+MoYpGYRvVofdr2AL7tFTQszPD4begLDtApum+Y35iO5
oBSw66tqQEa2yJYm+mjJjWLbAi88gVDD5WC2/QgvxJXpz4tAdAOEbo74oLmr+5lL
DsBxWIFLIVPUQ+d/IjGGycpUc6mmch+GmbnNHFY9SFDOlU9fevles2v3w13WrvQS
JMsSw3GRk+lYAf7eHwT/i+SY9EOdVqsPvaa0YGu0/GCVzAVFMCjlVLYFfi4MWeBr
BER89s+GK+SZcJ6ljQ35+PgzjFZjnSOhe7yaDq98gJ248DboR4NGJNtj5GOVMvCC
MvRuHZEGuHb6CNFTOgVAbf91IlX4ZumOjg72yHfoQJtFVkXKBlVJQLSqSButL3EC
YgKXAPoJTSsc8LOyKE7/IC3t4WgOFvB0YDtN7IDszLbCIP1yNwe0yI1jD/5u+Qm+
MTaIr21Edo4BH2sQ0sChzPU/HXhxJzWT/1NkHjReKdsxzNCtvXbuKbDlmn4j312H
/5sPhXNkXy8j45DnJLCRzD9GQEey8PRgH8TWcImT0TDunmebzBC9ls/Uw97+ZETH
4iu8V2xAuO8PxwugVftjrlTWH5FWgzctkyWZGba+FdpeBRkqlmqPigzIDQ/BtKa/
6AArKIxmb8pi1vmIsmL7ei7KiMmQfhulDgW5zIuf5yBrSmwjnItmF18xNyuY256z
VRKbAeljXp7qHexIoYOWB2+HyCx8yL1lm8gtfFWmPcdJ1BqZQRz/Sj4c/7v43RdC
L2dw+d7uBnihFEQVdzomc39USKkXtCvkxoNtieck/E2q/XQ8rJ/EsMiJVkopxe13
Wlo3u+5Y81PEZpOMdzz5TO4zNfkAuFKoNx+F9Co1w1TDUe9pQMPDfTambOS0jbKG
EMVvEXIsapl0m7B0QwPlcm6BZP0qeEppr3nreLBqCedwf4ZRS7Rnuq+wWB8rSDb+
yJXkAUsexllUGpjh9K909bDBKwMY2G80LCCVbU/lhN8=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BEOZdpRYKcJgtvfvS0P7VfZxVpHYn7lrwnUCsw+CjHRCkx7XmZGaoA7nfpELc1MP
dKJQtvM9NQr2SG81vNvXjYwu0yDTq4zzjIyu0c4avnheh6HQrRYqHd6LakQKfQdy
Ha69epLoiY9y6WT8CeUtw/E4QC9n6Tr34IglVenI/4ZpqUb56ec7SgKpQg+UmHos
joW/jSuOL70YwZYjj3yifWF5Jf6eiDAKHPw1gHJ6j+/9/0pM+pb0t4JzvHiSgPzq
ioecpUjBL7MvGEJBds+Zb+DVGO9AnPn+p0EbnxrdsE6jRRUfYGdNvDIokYR9JzNL
n32I9SJAbqBKti+JkiKJqA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8992 )
`pragma protect data_block
I7lRxEbjRdtup7F4rJHobYMqJ/kp9JIxKKFco1lEAz5pDL2HTJ/biFD89HGZPbRz
KU7crW8YJNfgT1NuGR7VPOey9Py7h3u8TTTn5E2qIuxAHdGYP7oK4HEwOI7d7K2S
4QQVtEraYOC/cI41AaKKYHB3K8spqaeg+vW+WQEt0IZcZ0g8Wz8oU8KlkhPb8zJD
BzPOUoryPqGnVCJGLd0NLLRciwtHILmi1pRRQUIMJEOcgOZiXNNLydQUC2zulQwN
wYCAAclCh5ry1u9wC6rgrziyuhEnlvsowH/RO3AeaW4OnqvdVET+AoD1Rd+kjPJb
7ZaPZ9PpCX3A43TaCxQtt8xuo3Ci6goPJm3U3ZbwHgZI/n+r2Nr6xqGityrZoKnV
4hDUrqPYR+J59fEuwLP4flASuLMMivSTQnDWvsfMyKhHvInovHWNMKoprW2LBHb7
ndZHZIYpoaji359AVGoutJIlwtQra2dD/QiTHsGTSnHgQEp8DF+vbjBp2pTuIzA9
qA37sPFeAViqotA8CqbftCYbhOIvCp7ForcAuOAy0ZU/VwYrtUjjLKd+MlXIAL2m
PLBpKD2HC1nqr/A3jJMyQdcHsabnksffK39vUahl1LXoJaShLoSkq8zVhOZEqbhc
tjcBiB+akeFg3nrumZKQL3U9ddRVAaJkYMMoieObOSv7pbkI2ZqNmncQoTSad9WD
jvoxS/g/CgxznE1sfCwRhyDVjBo31GwE3kuLUPP2JTEyGq5SQonVZaLExeuz5XTb
EtJPvANB7/StoI83pyS/2VojjtlFlAl3V8PxSDRvqeVSf7Kg3D+HSueQFbcvTrU3
CmjT/uZeLfUVNe4D06mCtCR4jGgPbpKzfikeOvBg9/j3xPxj8/KZ5P68heTZT8Ob
k7NyonCRxShTSWzKCH/LkWyZENPowkNqx1aItKvU/BYXhUihep64YUSOdIhor04W
DsaNXCJWSnZRJMiPxLcEcqxxlpeB2mLCzwq2bRI7fNW9abVrTYFcLWVFr64KRQ0G
M1VIATJ4iXGCWAaofSYBlYZSEiobIHOYZTbjJa6SjxjwCWHHi4g6lAAy3uRa5A07
icOd3voUivK01E7SW4XJd1rW+mzulAny26JvhEwogW3PvTZ7YX1AKC4Upvzjg2Ga
H+pGXDpiEDv9VCX/HtXQGZ+/9/SCWG5Zx7jom1gArLAQ1ktT1TIZQqeDNnk7Sjak
la69uerXcukfnscWTRhT1bL/8ahZgJpCtAd7CbaTRWLCt+73QbUVi27w/OpiBh70
FVjpeflzQlzhoHEBTU7x9ViB/5GxfKfZ1jW/AhZ7YDfeqWc3AXq5+G1e9d36X20l
9vGFabuJWHXza8rg1WDR7jkGY9fwA/EpwrQR7LnuK98Xt7yfsXCGA6qft6BH2mQC
+QIOjMVZFL3szzxEAZcagefM565oTcJgJBTXdGdPkQ5tbYCD6RE33OLNQNBQ4j4k
crgdVqRhk2kw/KwVntAiIQVr5lpWdptd4nSi8Ywb1Fz/gEG1QyR6d8Y1cHPrwupw
k7RbLhaFKEsdG7G+xL7OrTgwi+lJoQL3g+8wNx60XsZLsRusx/gdbv1DV6ict3xJ
o62vy05rVds+OPS4U7oKvIwPMbUAQzwi0aRORmGeNLAOtwmtW9tXXK5OiW64zJvm
i0He1JB37I+uRYE0z3/6IUflW4hN6vAbKJd69/ulZAECwZb987Fs7BG9bL2jj82E
ug/kvMsdO84v9uott71kJwJCLAxd3QDSoh4bWQSzFFJGG8/xowgwLddOkS7h8WgI
bzTiK5kQbhxDEVMu8hdJXqYTphq9lrO7DGECi2G7sgBsAPRUrtMF9ox2ezLbLOge
ccYf3lHIDxkBH5s0LKdlzX9nIR1RCrPsDRhjsbm1AvggBfCLvVoA6Vff1ZfXNqhL
AmNA/UKfp8doXNcTgWX1VJi0tLtruIlD5MohQyW9r2DaVC7/HboUoMQPWhO1HcLr
2sjexITTMFuzRW4qzXFpwg0hj4TyMNMn8iEvmC1+6misPwK1DQcy8YqAzkyJBNWM
XWUXA6OsjxMb7NQTJwVPMgEWdhYr9chid/BAZ4CGZWF+1JSOXihWAQVbpMmXXujS
OJFP7Yjhot8GyHZSHtQ24ZkRQQ+5XatDzqUPOQDsr09eTzQSECXfeEg4GFK6oyup
phzXUGtRZCJahbybSGKGNKc2EmIWbEkIUS9VFmC2ikdWz4xDn9vvS0MA3je5Upi0
2j9jvkSTukyODiu09PjMBro+7LgispLexZn/nKEHrbTwNRHfA8mKn48s2LCYNhJF
c/N6cgEfhWjwy8FFUheQ5vSxX4VnwJTjuX0WFsz75fbZQkgd3LZNDBWxBCy7dBOc
DjFasoGxTxEcB6EMG3nEB02Zo7AOGSs6HtvDRg1jbG+6+mMqg37mENst+JSly4PR
zmhldVbKx7UF05vv3qr9nVB+4t6clv2Fd98kZQmg4lxzc3q4psh3/lHmrHxTZ/XG
BQ+7gRXfqN12WRXwouOR5JuA5XadcHnDgKzYYbGJRzXmO/SFAaTkN0/juMSUsJRa
ZbxIYfcO8B7IYwkOOnr+Gj3oRRA8OC2EuRxRU29QHGZ6jmfzkWqkNxqZFjkZpb5C
BaJrNmj4s69tK/fz1GETRQdzibKtRnIevun0oUB1HIJU9aEybPhFKCsM2p/GRevB
GFwxLMt7lhIj3IArlSoCE6aIpRKPjDNy413A4go0kSbjFWeXdKXky9wY2OULFBKI
uOK+Cu8d5hM7/ReqKGbzXOCu4GRi6ooZAO52wJaVp9XQIf0aObOd9fb7LKBYpUGj
8ex1MVP7/uz4jfqNxCCf9Nwc1rXVTEtjtC8QQ2nqETbxiK+oyOkFtHKENz3l2J24
7PydNJudKesPZ5haM0nrYjHEjzwjjJV+vC1KFSRkbdTvxVP34i3mjsfU++fXjEyU
Ypmaphb4VrDSLKDS/2/43XExwXzgtAMXSi6MZNuOq9h1JAoRpBmNIbZHWZhFIDLM
XmvUDYAZuE4dMkW2G9ieVNN+JYN0CX5l3Cu+wZ4fi67BHxrxztd1DSjB/xxnXCnQ
HbEhVzKuodIUvPsYhb3fOYK9HBWtlqTNpxrAbUy1vbfiSpzo9mUhqvAW1yyx5VYG
oXxFUxhgB1BMhZYNP7vnpZzus+FJv1FnMYzFOczbGTzSFOd9Xj/a0THyNvjebywu
32zbq6/LMFZAli5/lUEs5B/N0y+/nWQvsgJ8CJGxWWmEGikW9CkrH+telcMwYiu/
Eg0rV8zR5uxMNIDgdX/pyM0sR7ieJi/zWcyyI9OR8e/pObod2S7yZjl1g8p0TPLH
yIw0Igm6BV82mDtQt2slLFUm64Sth5oAwc2nD7Nf8NBAvgBa/JtnRJjH2givZ8sT
pdWTHIzHTY7PChkktEH/PA3MIllN+ypLbHpkjk5dYMRMgLJJ+RRhTe+NBQCbu/QV
PKh21wCvs7K5XM11Huu+Ned1jBt+NRuu87Lu8OC6NNbk7w9351LBQI/mw5A11TnI
7QCacPEKNVZ9dQ2Fwc0JXSb7pLULBWvkaSXMEDJzU7txf3C1XBCp2AHbiv+Qp/zb
2ogtz+NiUFrIj6HJNyZxktZ5CHr25mETaIfcLmTBQHdn4vv4PSgmg/cK+43pUhjk
rR5F+ubkavTmKotTlj4+FugO9L/kzTb3gHgAs9COEVU5hKIpNJwYkaY1PpcZq5XO
64rvzsZ+z27Gw+U25YQyGVEMXGNfWLMlpIubafzC8fnFdmfCc2LxVVH3rGUsNOjC
AtRRwQt29TTKDbTx+yI0v7IqCz4uc7kSsM2BQR0kh/xypJ+JAOLHIF4I/zuTiX5j
p+mX3qez+ENd0oC4LMh6GjkmRMtd8pNrcsFFmZSqb95mzmxiDY6aMBLe3LTKEprj
TNbVmLIcgrSG3mCSCO9utcVGwpf1m37heND1aQUjLYeb/mame6R0nqRyqIUWjg8S
+/zqCwGpVueAUBZp6WOmGtHpcKPK4XsGnsMY5joC6CizNh4CNZcyARc6ATIpiENR
eSqOHKxpHMFl6C17vHRIFJKJOg9FiQQm4NoY+/K/s55sEM1M8iW61uMTxS1aGB3J
3Hf3Po3N495evI1yxsvtZpq3PHarL/gjnTwzOPUa3aM57rO7QDDJwDcFCCH+qkaw
LBFIBNZzwHpiBKbxXnX+YJy/fyyaiS5bqccNgDq6l+d9HIu61hYEAa3SEuc78s9y
iP6NBwsFYUelUEOvo/bpfdlxEpbEcmflUB0LjvA0OzXjr/XahTNyJD24cBmCA/bW
jwT3iHjyv6ql0XFwUS51cGf+bGpsrdE4Re5kdlNUr66lwIcs5UMaF6UgjCOBZ8I7
Up4Da2LutHF5fuyfZ7HV6xIbIzSbu5CAV4hwceuXn0Wx9YFjdkQzSes0wLacnh08
9Hs3R5EOS7/WKao/x/iRb+t7yuoo/MT4o6ndLklAEEmKiN8lhxdGFqKggBXG2GwO
uTgv8hOruv1TZLgsRySylXKPX7XSiq4q7oQYQkVgbVr2C34q871EKOvgQj9eivwF
5K7U1hnvf26evaGAKwwK0WoiO0e8VbkP/O0k6HgI1w937yWf3RVK4SUF3Nsh6vQC
7gdOZ8TezjsY8iPnmW0jSdIecAS6CnSHBJrF+hdhTHKH6w+j8Y6O08iUU06qSRoA
2bMlUrw9PA8ioy7VO6RpnXS9kvDQF9eGjMvH4BG8nd868gCrjLlKUCNdHcu4w2c7
eyQbez6bbcyJrwydzpNl+Nf8pArM6lCrtnOndylgb+3njd1GMlu5KNwFKFMV0icw
OUypOORNdsuVJSjLJiTp4uyNinwxu3d2FR4uYeS1XGzFiezeBhtTfaqJyxVovMTr
cDICG3+I6cK1TCwajB6b+1GP47gsGbq5fcEi60AqCYbG6tB4F14TXVcccFegUGJw
S3SuI4yrr2Nt/SjdsCu7wmzvzHKRVLlCQmsaX1wsR41lQesWM5CbX5U+an9WH6gr
nlagnLzaLbYfTZRsCtKgd9qRgcPe2TzZFR5jOh/XCdBYN2ZkIMhpCf9pFjDZ35wG
9tS0KIodwhXPzW4GOmO+/PGVgg2KHuZp1fj3IJ2CKxi71rrBiJ8zM4FNO90zRirF
veLADyGMOuNJNJEdBkB4K1BvKsE0er3Kgki9rHCvtzBS8EaQRJjXMAhwGzx3fwA3
+88lwggVs7T/xsNxXWSQoARFvSd02Q9op72X0eXHNRCS7TmlvoL6gh4+t3bAjPHu
j9bO9TYBigMpqRViIVXHF+yI20uFKIN8zbQ9KKY+fbQzD3hKf08xibQZ/D8TL4dD
Nunn0FwHUEg7RaKHbN61zd/SBC2dHIcG0zQr9cbnq9tXoJqoQXh9sff3nY5RIW1b
t9IESYRXGg9D5ciLVqczqw343nAyPPAp6THPzFVJgtj4bAyVswlp0C1kMEzn/aeL
kcOkPfCYj2Ub/jFG30FZRjB1p5mKGrioypL069f3YyQUpMXkdsdq97Ih3YwsLBir
ZM95I2va8kC+qKyXp1A2jiVt6hIv5UbhMu7soOdnJKhUQON+ivGlZNy+KwdKl+Db
eKvb85xgVfRaTx4PG0jz198lTCLfcEOwpKPyuETsZq4kBnh8eO/QZ9Lkx1Fc5k3I
QzkboiE5j0LGFynItVlB2sMpJhF+tUhtAlBw9r9Q5JJr3gEoAjoJ8KfLG2zvbTFR
h+7DkT2M8QoaSgoUt+RFg0h59f6VIlvtZp9F3CY7DQOLf3cqEx3iGG7joIB6xAMI
sekCKb+cQYTLTxPEZoa6KXVZq7Xnq+afLbsHNqTqdRBozJ8143w31dmGqWeZXfU4
NrfPWGGlghD0oPtxgVnx/eDeXdPthNESly8LgajizNxPvHTbWom+Dn9HJ+UNuH6u
ZMriwcQYzoozyG6+bHJaoZO3vhJUFDz0CYjPCR3ga0XmPY9yrzetYTheMG75QdwH
u2YUivUUCtIgZCNyVgRyIFY2w3SXPnP9DdpUShPMB/4UXINbjzqvMrUiwhN7Z6sC
sIdj7WeCUcoMNTt0dMGOzTRexE6rT2+FfnAyVpQnjX9gqCNzaRWQosbth6wNeumb
HSyO0tzjhgBxOROYcT8t4JYEKx14ZU3QyKBHSGX6uPCP/UwaTlngkXMEJCEdvRt5
B089TQtB3szaBqhsYlXEk90EApx0fXpzc2hrZ46uTTtZQdWuI88aZdsrOXDG9BXP
TWrats1DNvmz7A4LlpxGNtwr5o7EPo6pmEfVGUmQiP837yMDzcX0W4UQXfBS3+xZ
DQuJ/Y8zBN4eoYAC7MTMeNosaHEgXJlHhZ7sESOaWdtGf1LE7fIPiQKRs0xzJ4VN
WN7bj0PCT+R3lRbtV0sBvnGPbKnFinPSCKCyx+ztJcEHHhXC+shLDcNGM2S+5eBH
iPBszB/ZVtuGGyEiSIURA/89ZQIOwk0QPbamWPqQM3IeNGZM4Why3YbBjLooD6lC
l9JX0XskQ4LLTw/8NA9NtUEwaIFl+vv4CrgWWu8zocgvU5/2H32Ev7/KPR59dMJ1
321icTLf4UbEjTUkrkRQvxrclm1fY6rwBklPielooCTtZiyTvQ2vYw8JtkFy1RQf
f10X05A8dXKYwj5y+yMaV+k4W8rONbxjE0HRQxegDWMVZCCQn9AZpcLJPRAnd7Jg
SC8YSz3hk7R3yYLf4nqhCpcTmYHyHXuX/VH9HIkNz6TM2ee3zr3EPunOkTO9viUg
6JySUGmFxFps2i4xT3w8cSx7YW6cuByHpkEZ3XbNyYqpNNtkOocm5QNY/IXPhpSn
Kn9i9V2JaYf5o5xX/Q2Drz5VUB1VEiPEBhxrB+rve3yTbTn7XxcEmXHFRKLPG1VR
H/5bhZGwS8WtosDFi/r9VW06A0zkdHrFredtRqTTfMx9/IOlOHnblCXvbBpbYm92
Ep8y3BzK0PS+cEEPDxjLxjiatzxXPPFTd3x4EJZfK5DLf9Z+9u8+GCNDeTn9kqS2
yFI143Cv+Hi/b6sXkvNDi/xDvacVo2MQ9koVUwGetPKHIB6Uppj0Y0+3Db6nmJ4z
1V0L5J5YtTmPMZPIIcbAzhWK1USRL1FnGyOwMLBWy30N2xWe8m3HDgkqVVJHD9iw
BSH4LB63WL4WpTpGd5fUqsfwBP24LhYtoFKdliiY8JSmSBeHGYNqT5SJvl4d/8jM
Qxp0BONa02Xs5/4D16ouRVkxHOIdhqGZ9CnHiPYRAP5FLV6bHmpI//hq0vXXo380
a7WJHvZjSEReTDklR7y53bVbO2/Ml8w2XG/ktdR1VoKUzkO625MdZ/9QYJZsx/Qj
peP2xBEV9XAK1NsVEjB4nD0b64cTTdHyshd+ZDoUtBD4iFEsK7vZ+sClUJHQpp1T
2Ppt2r78oCoQlmNwFkIMsFF8/YMZwOIlggLVd5kdkuPhV0UilhmMUCYtNuXudE30
hBUx2Wbd02V9pibuPJTwtzbYghY6hZY1vlDoyOpiwNVtjTiKc6zya35yWlQoWSLe
8589VJbU+FtmYwJzfM7PRqfn92n8NyxmgfggFueKz87HIpHj9SlseqWhxfmclbq5
wYDNITluoloDT3Uv6DU2vYKYM9/RvFlMuL8S3D/KOpMZEOphyUQySyl43fT9hrp4
7yqPJKvZBRsf17UNro4CkU8l92aRFyAulqgftPufm4s+s8BsC4LG5e1R65c8k1ow
ScNaKtGR3br5t71aoI38jnYQsTAKl06LYzTynotxpYoXJhcKhZDllGCvt5WBiRW0
vQ6FnhSQlmRMkHv8/3FlGUGgSdOjxCnYG8BHDcnJmpq1O7IceoTmXMP7MCH9Xsbc
Ea4QlFpBDBh6Q/mUkOiSMawfe7FNx0nfe+TZXyw6EhwFsed3APLjs4XsyAOCbrqZ
tmIbUSu35nTwIPGc9FmMRBxGIKSRJzwx738Y7Nv01PQek6Y2WGNgUMf2NgOJqJnt
Zz2P4oAghH6zxiMK+8vSPH8tPwuCU/KAG8IA0AmGKy8/CXkNDfDakqClO0rXHnt9
GegRb5guB4LgB9d/l1Hi0rRK1r9PMIQGU2j/3TwEj0y5tLXfuFFSACSjgpncE3T7
57iv4kKiupZGZNYcwmWj6Flp44HxMvhG5UZE13KkYHyksqUC1dke9jJCtORw8McL
OrJ81V6xJksvYarWa/aP8wpsw/AdPo0Ogq1XZ+6v5N7JuXaC7sqK8Ah8SIy4Uf0E
mevHuWBo2Od6tWybeBqEXtk5e4N+xqJZhf4D0shqyVL9fPL885iDsTV1nm2tUUD8
Wh/7nB3fKqpcBoissxrCSLvm0q+LWcKPRXpNtMSNcWK26ACJUE/Cdl0NZOzA/7L6
duBoDkgNQveKm2bFNKibelt3lb7fJ5fgCix35yDcDt3+09nPsOcyKMCV1sER5fS7
8f+cp5nqT8NV/DdNKnFJEXfI7pF4ZcCZoZGnKyyWFmn1FrbM15ibBjN0IaRgpJRR
Uc4KUfRfXBYAd8iWouAME/AyNzc85JxTwOsc+muWOCo6fxLEhtYQQi/M6a1kyskp
kWn0BJcXPNeu/t83/nb2s6WN07Y5b4PT+4IWah0oRJy0zLzCiyp6WE/00VW3UGdr
4X28X+8sJPlKSnwa9DmHR97W/lsfISpccPvRyhpBqRMErYsb2uqQZVyql0lpW0l3
+IpEGvOTtPtzW+aYZwzEYqTuPpuSlj39yQ/of65gbXBJn7UzUluo+y3zDLO5fj7J
bXvCYzxTsDVBdK88IUOakSgIT60A02MBSOFR+BBtc6TW/Yzn6/hcHk1O4WTzM5nt
qk3Swj8Jsy5JOjXy1vC8aEXegSDA+2qhaqEyKBzOpAkvJAtS5jjFG7OrFBS/CT7I
tBovECrVnmCImjtcI0kh5kuLg4F/MHa0kWo/Ko78oITKOzH0e9EZJevP15GJYTDs
tJpqWLwdoTFJ8ZODbt95ogYeDah6InzHZ/DXO/mEzoNhdVzS9vNduckBjJOuffh6
V31j4ao0UG2ffxkUe4i59UsShDMNvkyQvaIZPqP4Q8PP3F3SO+8UwBUpLkufEg91
ZAbuEn5pRR2fVm/uiy4Q4YkwgrFKddQ5K8BAUAIde+nioSldfjFWXBEAucfuyOoI
UeO8WsnRs7cxHKnJLjJrstqI6GDNRhVg5eHEgJm/e2i/KoVlQS0pAr+lje+9yQFK
ocOc3V5bmBRhaJAC0Vemfa60bqd2TxiX5c0HH2xHiSqzPFPKRL5+q0d8BspL6qQn
pntRGYIF132zUQonjqzQPqr4ahovKgB+L4nw7Mq/S7g3tQNhfpqSoqy9VytosA3J
xXkeWOmKbR6cV4JkABprYWIpmsJJCs3tGAaBAh1rIbKmYTZoJUUnJMTf0GuhbKtb
LPWodrH3I80MB1b6qp+F7jobLr/asnvln0fsJlbqE5R9PyHvRIUDau82bd8/mWQc
o7hRSep6cj9fdSVYuv/ipnYfBUSf6js+kXHv/C08eMc2dvMSjUS4qf++AWrCmFh9
+8EhPVEs26J9lyJx8/9YiGT5tDkoANDDHauppLj9GnWPPwmTfreIAku9+LRk2M4d
+TrRuUkA0ooOlib3cVLxjfISOYrPI1J8C4ddT9y4WwltSDn37NB9axNBwn7DNHoG
h658xgpT5VaAjeTF8ashIYx3ZnW/iy0SRSOnoYVmBqCkabA9aLa976PnZ71RUczs
0bIHo/Bal9SFK824l3JvnzfhH31P+ExXOghi8cWNLUNWUzEq1bIDYo/7IsHIvwF8
mpy4cuzD2+UvVHnFbalsxaJMgJ8gfZsKWFQr1L8sxzueJ5r52MPLgAMpanZUqF28
kdAWMMf10deUZDSpi/jWT/EVWm0BnDK2dbXdVS1U8loD9IzUjAeAPV/Ptjqeu0l8
RgXKlqtrcSKzQrTLRgDvuLn4nMhTzmAPPq0t8nE4nfuIHNTdgJVEd5Eo0WoV6tOm
h28dzszbbS87Rnqd8pR9tnMji1QKbDRCiyR/A9eJEjZ3+1Y7NauK8EikNJuVilpq
rm4PDMq+px97yCET9k2ibV2xfJsN03vh+A8MkiYxKLndgyFO7s6cszBL8KijW7up
9PWAdlvsShvP/qYEww7pKxTHdPGTn/HrU7TfhdCjcL//sYa13l9N2IdSj+3PTNSY
TJ7aNmBDuMmHh20vVUR7Awq95wxfx7zV3vYYBBaqnbai+JbSY0W2Y/fVZU+qADrQ
GU+psXGduziXhqE9Gkk4glw4aQeO60GK1YF4QYVnVfzzWF0Dmlafw82budXXvTZB
AWaWH9vbJ+ImjKHbNIjd78jj+jiP+xmw91bKuPZ30V32DXKsT7ZwnLRcIrXhK21Z
+PiazSJgYeXx/bNC9mFXrCtyuf5ZCY2Q7ujVdzeK6ye7kSNfPACXZi5XCxdoEbvq
xs7rIPlHRPjBhRJgG93WxhTaZdzyopOAP5lj6GB+bSMUgO1n/Z0PzAPAEpRJp6V1
J5yh0C8UhbJCTQn7Iszmwz3yKx6daKRhu/xS9ldpNmz+QcmALlilgZp1zDPa7bVz
BrSNAgT7YYwjACC1AnqNscxqqNkvnzNr5Y+r5oiMzQ3ZPBO1ureBJB3rrk5soI4K
f77ZiyW/363Eb6nXas1EFc/Bah5u/9GYM6XwQALLu1l/dtLEMUesCPt0AYzqDyRS
PH/54saVEqMNhISn5tm4XtMxNyAzyL1JD1xhSueHuqPR2rFpJOzhCtOajQh+rycG
T8NWReVGCSF6crxOEzxvHdhZwTfv5X/AciPcy0n1QcJxceG6ZDYx5ooZEJd311L1
r4y+sBz++qBDdbNxGIj7jxPAH1A8DC6Amp97Eh2bASE0t6Qid3YxjVHXRxjOWKTg
4P2rc7YIbPqA7nORA1MCkWEHefHLEMW4fZG1uOQT7uphAJsMWTGS6p0u8gMQELWI
hbX8tL8/ZtkmephHNLSp/BN3oI2cEmnrw9qmaVZfaDS9DIgRhyU9Ep4c+NdJ9eUa
Knw6HusAO3xF6r57Gyc6GtTOBMSB5mo4x0fcdpF3b3HG7rWmKs+Ho1JkPr22iMXt
anXDxyjcYdgE+yTr0bgjVk9ed6nGNOY26k1aEAF2DUlp+c65XtuwIg6TVKacwZHT
Ez6x/OStnfEY1+LjCxTYe24tZBMQHEMWhdH0fvIZNF2mWGyjw51J/F1ETVZ7vcT0
3Z3LN7rKYmUqLsOm6wSY7YQ4h7epCJaPTKeEEzO2ppzUXlfDZh8FUbqnKxFgYSdz
PtwQKAWC4MYwORRUVFMLb7SKgjpqDaz8f59bXqsPFSVZOXbM1FbVWlGHP5QWxEyB
EX0uorgQUnRWf8CBonW4NDGpWmtnju6j3FhZudAzTznGwwl6+EWgENcfCnVHD4mb
1j2BdKoakUBwkLjACSnuV/hE6JnPwjwU0bCS2yUA3s3KV1MCb1y5Tf2QOytR+D+U
Fynv6oj4LmunM1sapB5zGf6I3eWkGE6ODJLawfZ7KIUAvIRb47Nn2GQfuAhdNmnw
pnrSKhuCV8qaiXF+5XrjsA/zlQgqy7/w0R1eslhjHaJIR5o02hJnsVaLq1NJw/Xt
uscuQVcIH7eqU3YGQxnlwcMTcs79pE3yJl6XwpHTzorVoTQv+llmoLGOCGd7K2tR
1c3wzQRD1Z4hq0UzPR6R4v46iptJYT5/WqI7rJdP1M5k1BdI1hxd24HWhfx2Bk9G
VYD7UBFYUVh4MXU43mux6lK1bk34oeq33eFcbwjiRzabfc34jhcZRPqhjzhUruPn
rpMBnJ1C9mmHCqZQJDurSbiPZsINNUg+sODYe9TRlpqSo1loFWDa4zk3zsp3pLqK
mdVZrpt/FA7HbHWRuYGzBOTAYYluAUr22alW400Ni3rfZMFDF1gGD8mJ9oE6PhHu
xkkbOOMqRQ5PalpdJeavCQX3auMbGGJR5H+8YXIIALkeqiBGRAhDYGT/tG46q5i2
bsFLwBhsmBUF0PVid1DCIfz84+7WHny6GDN47fSlxK7P0ywvZ3S9oWsgwujJMfyJ
utpcZXT6FB9mkfg1Po2svw==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hEA+V5AHOCDdD9c28h2iGuNZQruTtBLPEIniZ5jumjRsucm8EZaSLcozz2Kk+NFv
g/KKYsAeVW2eQ8FpeKPUnsw2ftdpYEKwOWRxbiqBjcZWUao29zzbcRgSqGtDEoUu
iQY/phd5oJ7qUcFCiXGPuIKKWh5seVXjJZ0QSyjEcHR99NlJa8XZMezP9759dD1v
xax+UyWuJAqcczaRpmNGdBzyxCG5tLEQp/NBQpdL4XjwWIqn150V1J+NUnivpTgJ
OCmOSUXT8C8L2yzfeCeKoTGH5gWBU2SJApldIJeXajsHqViTZF5vMho2abOCX62o
XK5Nah7x5hKZY6tnXwLP+w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
wtqblU2hUNvdank9RIUsKP6rB+bnsz7TA+xvT0xcVozKda9NcBwcDSxEzVyiO8+B
lkf1707rB8Mt0ki0olVaj/kJFNFoCJFLrI+noWRnVUl0MjzKAnanf0gqT5WzEDMU
gGjcbrTHuj1eNvpAzAP3K2gOWIB4SNeiL3YZsppdq0Vbfcm/8NuaKvm/HSf2DYI8
5h2nDrbF8dvULog32R+jp99hBcvF8BL4R0H57jpzWKWa92EHLWEfONvj66LvxPXm
VwVe5gRPn30/jqoFtjcVExGQCIk1AtMexZXVTefOubDmBD7EjJvDPuUoCCkaKB0V
Iy5ek2bY2KcfkJHPuppovbSyvEGgnJJW2v2Oc+jl2JqUkApkNygUgS9LfmQ5YLSr
JWPFmf4JxqrtEZQ8qkFnjJbhIvlJoksI0Imn3QEltOSIydJCHAIPSbmLIIG6lz3+
n0FyZZNHuzjR0Yqun2aRUGdJjNt619EFZ7JFpdmFVGhGP/AfbmWn7YQcIRcXVnk8
QWEAxsRO1ypsOep5zTNeAULJSH/jIf7XPXWdKGtpRhwp+xjmRz+YrJk59SbNcUZJ
e6RpgE/YMbT5xjtSayJlsn8INK5sreToeUuvqAmBTqLxfkoJgLQ4KhzF0etdgiZt
n2+OYLhkq/htkoVTgl1aLGwUceb3nV/+LsPCmSSRfC9IEXRqVSol7SUtZUfqwnPC
0Hue7l2C037qhM2L36he/is3gY4zb5l3Y+Lk430mCvap3mOTbqtHaqpPiuXKpnQ9
d/9LFYu27ilL4ve6vH3t8pov6qGVPhc5F0FqQyIBV60lsPCzx312KNCg6qvNvSpL
46kWE1oowlghW4m8NkOmNoMDDZ4fCe2VLaAeE+1LBMbe5k1ZS1s+jHp5Z9auiVSW
QUoJXz40u+UGOIwjmjvAGXfTeFpoDjWwjAuZK0T0DOab/d0/3ZDTWs5hgZHhHCBY
w3rWo4VeyMvFfrvyulgTw/tzQV8Cc+OdXL2X0dn0adqmTsFJ0mL67c7FlANjFjnx
WCkvLdW4kT6NLFfErfGqrXeq5KRgynDo+BH+E0gZvlF9QBycbCekl6fy93ZkcUvK
p0ER6SQuCCB5BONSKJkWPRSmTfUKZ6l3ffnNiDWuk5YTzZmTfLwCN/Zq4m/Q4xwG
K8H5l9rOg0aevutrTTZ6s7AjXYw24Yo2zXRle4ni70iP9yP+y8LJhxHSkhBYmAtB
V5Q/Jpsr3zhugn3pOxA9scMe82ii9IiYOaDL9NU11W1rRIzol+vjuETx3Cq41NEb
u7pczvP6RPloqkXRrUZjGkARDdJU0JERfUeMpPmXzQS2JYp49hEOkXnfg9SKsb0u
WsB4UHRN9Ip7gbxb16ZX79zFzi2yGMhPbtUCdI87NFx8WAJX7B2T1e0NFxCFA2fN
G9rO341QBXiVsEbxnpD1b18n6r3sXP8YKsKqgXkNOowS3jgB5zeUTAM/im4/Ut2+
qCQ4hzxKbTx/gJjeZJU8qKGXB84fhaMjfXq2vsiCi9xSV/m3705SIowF0giqsEj6
I+6NXrEtjVPGjlyrUgR7ZmypfCbWdqu+OzK4qhPfSKFYMkOzes/+wAqTw6jVAknk
j72jnowzuZYO512LrcbA+Z6mQw5kLwiiRiqrU9TRct7Kd5ggAoEm+yn3Y8Euqedj
Ri9MxtTt6HTh3peweWzfIBQHCd6Pdrgw5M5wfIXXv8bkIHgBDSeWMBm59qeYnvgF
s4FQtF0GN0UuAUB7c0qCxfr+0tVA0CjrA5Xv6lkCm++jPQ3VToA4Ry9K/BKtDooB
uFZveCYAt5EM0Rm4070B6b6PN6dS+tO2tHpBcZbjMJAxqoNC/Z0ms1NFn4i0VvsN
KY7JdQUrPzxPsZ49HEEc4O1vCyJlCBKSVcPztX1yWQ3+XLH4fUDSsOZy8mdw6WXN
LH8GfENDK0C4ELDGDR5lX1J324RXbd6cD1+CgOPFYbQ+bk1+Oj9EgWtWDNz3tDpL
8DIS1kPgk4gtgeMf6Cbh8k4T7LEix6yuYMhqbLhoCG8KwNiNEYcwdt707aoWaiDa
pfVCsquAEAXqN1qUcZ0ltcziTrLYt26fkfEk5XuHhtRU1J/WoknnnIlcqTr4b04t
jHozoVub7hwvejdQ8x+Lv7WgMOKAB21Zda8Md6bsV7YuArymdzIODYmFzKiXvSxD
47Y4+PrvbjUdSvK2KepPiszbmN1adl8n2DfSzXrd4rnGP9RXoPaoXiIdjXLMXEZt
vlqc4FxcuqTGqXsx5PxI/ei59SciwLIpXV7N7WDLSGW/By4cqcu6f1IFHA81owaz
Gj9oWhCbVqawxZkcN6E115vf4ZiwQth8GMS9syaZZ6lENuYjc2Q5i22I65KyL8Re
q0SkUJUw1+9t1CfX+NnTL03lJ6UIDnPBKOKtmgfm9F2IDFP2NyGmxhMNRoQ2WuGR
3Y+qpljoiXqbOJ2vh66sg/8muKKIT30nCRkJrEHs/PvNzKMy5f+oF1QzFP4h+2Xa
BWTLmTh0oKT89S5fGcfN5b4A10TjkTdL0fuVSaXhzIptsI+CvZm78jPoQkyb3oJv
XnI/Ozbd4H1I6vWZBj5fdLCiGdAModT+dXnXBKkoghjI9R/7BJ1IxmFHlRXNwtqA
TA0y6fMTA7V2R3npYtT75JPvyAAtAbB2BGkH/5EEyBNRSeJduAbE0uORqREQbIGS
RiLYOKFvTMhTVaAvPVe5LksPr0DX7vJ83a5YDhn2ClXlYqeXRbRvJXnDx2rUoG/n
QXNa9Ua8hlHC2d4ID+xPxBCCFQfBbK5QOJtd0zOEyM+8YzdOnR4aeKcTkZlKRoxn
PloyJ0A88OLur52m/YPZw6gs2F66BOv9lAq/5+/2vK7NJMN8qf0dl0ds9E90/ASR
eFvaa3SRSXJGhlLvJGw5IsnmnlibRY5keaWz7CxqfvXa/6rrlnlvtyqB/+DSi0hA
Nz6kLlI0ftf8EuelMGKtEydoUmyCi7JdKzXy+OdRdZXtn/VQlNKlWJa3uq4G+2ks
uWlZBCCRepQyaVe/xIRfC3HG9tS4Grz3HAJm6PnvvRJW1j9mjIFBFOIJ6Mk4TbAT
gAJsM/4fhN7knNuyMZJororsDODQKMq5WTjEkaEXYzcv0w2pPHlS3EoAUPLyQBO1
Li7CRYus+iqRTRL4CKu8FwLvMZogCTyfAqfMabM9M3ERagQyrUYL7P7tBI6sl4Ua
medswJDcdaqqTOEvDWq7vmw4jDxf17l893a0lr5mq427kJuGh590ES80vf4BoOPX
iYWiOAqugKqnG3AFkXa3wBHrWtScNJNrnEzA2ylmDPNDPYxJWWoo1NDIMyOQuojw
9UZowxipia7/RjInoB2O9DKl2mAb+4CYqdP29SDIjfDfh2zuD4ENfm0lL6ktInQv
9G+7XKtGJnBXqDgLH2qLhF2qJ+3MKYKYvAS4NarbbdiHh+hkgij7GkKR/vtI9zhb
KdP/daF+p7SSLociWREsG3Fx8UpqdSYu8KKJ+5yHk6gJ6X0X3xoj1dfyM8fhgO+O
YFYXInV9OYZIIQoeGeBgSclcnAczHsUZuddEjwsKXvNh6XAO1GOc5aY38Oj99CDa
ToZE5Nk98pJT3+hB5Fr+VYZNsgj3KAw92qBBtSaYOJRk9SRX1q3FH6R69rKAM+3R
5BoG3A0wRtUNuV+3P3DIcSFcDvfutUsni4q6BNfLsaRWURA7N+x84oxsbNXU3XlJ
BVWJfwQ5FF7Ak/owRNiuVGEPw9tiBg4UlMgbLYRRrAkE3Ny+ZeVuBihH4HgD3N4e
/gQxU+4vOzm8Ybsp/jt7/1O9gM/K7V/fbRl9miGhiDHnhu3v5J4p4XeDRgwlD0o/
iJZcpb/D/9LQP/5+hhUpiBveXodma+GK+iCH9DclfmELa6MIqtrDQXRkgAIlpvux
/2Skx7NPsHVeotnTpej6m/2QWcK0VCN4nfuLsJ1ZSx6ay6bcvUJyTovkurZCqGXt
npYvTgcduE0mgL1ghCM6jQl6rAtEaHIB5lJQlxbyrn1xOr+5nuvJasQHJ4bCqHVL
XALImp/sVFyUH0oMkWKUZKwwcskFyuJP+q33/kUC5rl+gDkSkndAh6z/Ts2uzk47
u2sDfsnIsJdPCPRZlLZ2VLIOpN8QmhEVxgJ7zKt4jLbvwLWJcxE3hvTUO8NS47IE
p1aJ6QCdK6tEM/+AjtK5NMzq0CUECByDnhy5s58eN5abKW3rjT9856ayGfpBzgyo
R94jCtqKnLztg9jkFnYcfQe7gZ6Eb7PTMB4Fx0zhJw9fpJJ4qQWwuzqzISxLXRml
SXRb6WVKwiIMzcZkBJ+O3xYUWvwpmpylrngisyRHdRajgohFAG9fHtSO8Ajm2ssy
RsiKAhoedYXVKTj+pOlStbuQjP/NjZ7tcWzcckE8Zp1rlXx7MoH4vfjRmsfjNIwZ
k9ZNlpyHIieJJgqQhvkd2NkjdixhWj8agdjgwS71DS64u9/YrlMOZgAC8j6PGf/K
TSq7HjN+v+P9UwNujjcxvSNCHqbJAXZndFN/J7GTwKgiPEfYLwZ2mCAnWtrUEMw9
jmItaawKEMG9NXCwkE6A1gXIhkxBIgidZjOV3nD9JHbqrPiSAuReXraXgTLJRwuv
HmAjb6UmJD6hUpIIgRsqB7EjAY8QTSgmshPpEu7DZfSCPng2oqdPbgX3yZzxML2u
oej+106m3+khTGHFt65AGxAwqtoFd7WMCxeo+trCEwo80AtJuBcRNfj1zxgcNTTq
mvvB7MD+2muqvfT2ogji4wvpiUcQ5ShtIbF3HIZw9UsUDMWvRX/TbZtL45DlnKd0
uhBGzPKDORttc9fr3oaSkcxE2CU5gb47xZTTOVNwOfi1pl0mYPfTN2r7QNsJCR2l
DHfYE4JPh19JmY2gZ1RzBvZv/eHCfxvfojYPybVTfq+qzteasTwlioPaxDi8sP4X
WwAxhfiZot09aY3w04nUPiC2C8afhMdCCFM0hi9GFn+/OaLNROStKRcTXYYMKUX8
gPT+qg2Gyl2YI43mhKTVdI9gKIEghT9g+lyp8/slIsxzmVSeT7I44MVdt388cllZ
uXopdgkSnyQWPCiAa6qBjg88fcnqoUbYB/PRc4MLvCAZALB5T53wXm0hYPWrToN5
AhkSci0K3mstct+LiRuQ9p3eHNjthEJy97Lmp9xDUo8=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EIConqsysKsb1eeRracDplTe4m4FWLSxtd7wzKYM28bhy8ckfxfvK6l1OvGB4xK1
P4YmXFcTsHzGdknGwX8gPF7FjF2pm8ixXdvPNyWwvhFE+Sg2/FdevVeWsO8vUAxM
eKdG3Eq/hxlAzmp9wR7ZPMkXL05mCKOQpkLiUNpdhyDsGJxc2mX9DQLo5d36Kj5H
uq1cjHhanKTEYCNuGyOYY1iY3C8H9RuG67eSRkUPqhWkLSof1Z7L1wINWdErAWib
b9nY2QaPJgGjH/iRj09GVagWOZQ14UYzwqffghqh+X01r5F4s8jbKuxfXZcjDE5P
q5/8DZOny14fEson1lnB4A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
FuRyGK1eFiitQOafEc6kyDy+Mb26ognwfmE6sGrX+/bMF1bNlDHMfV+pE8zc9+Mo
xQj3W7qsx2P85eIE5+29jCgi0QV+BnGwWFt3Y1PNeaWbe4SCfXHBeCGOO1WB1Jz8
cemLavrZP6YJCq4wMVRzRk4hRxvums9UAxa7FwUvNiQrPoEr9pgks3MHHAk61neF
HJpY9yKY+/lyGWxTpN9vVMVU8TaVyFW6F5cQaSiUsbYwYMX/AuM57XkGAHSmw5/I
OGnP0hoJvUdOlNbCm/g6nubMnDS3xg7eneFO28wAgvcJDmG16OTVoJd9OqC2ok8f
fCX1h+3ufCOo8EbejUk1R2nrVPrZJ2JMYHTCpobhMj0eeHMun4whyoozHEtSxz87
YJjig2aLuZP59oOPQ7zIz4tnZjm2BG5FQ9SB1TSS/hyOYDGBx5LfpD58Ad2O5+Qf
B5NcEc2Tu9o46kEWwxrk5w8f4dCNaZ4PBXXRRTT7mpMVlnwUPbCSfhZBmxdeqUEU
8P8dKPQS/iZdyO0UhbdG2jK+WEjisG9lglyIXesHcJ3CHC0XFZyFIG3yEQNRk2e5
4wErxUCErLzgeOGenjZeJXOXqYCFMUtKcWYcsb9PAZ+yyBKWe+gkwMIM8adzwtsN
iGf4h0uRNKgPm8ybp4ZzUDBQl/9NyANxRyntx6kOWCE2xTkoBLjYKNHEa3N4B63N
HRwL0CrpsAJg1ceSqNvMhgBmW6fxcaHeojNKrlRXdSFf/qfUZXBu5488Gmn9xEIo
uRPEpb72+Y4+mwFe+19O1NXbaE++uC2eMWhv5p9eOkK+oAYWq5YQb85s1z3YewTv
f2aqMUJjCGauPW/Y+MAhq9N503rPd1iezJSQFiwuuDvTlBrvGqyO+qq7/7TBPVqS
VMHpL3/2d6WBLRIB8QTeszGHlansoSDDAdF8GBIo5u4JSmiUF7WmmKTH5CO5qCsj
7pDccelDUzbPDrUXhBTZTdAkBZjEDVlFhOyLVYQGSqBxRBL0f6T7ww2Mve+CoAoi
P9eWrr90oi+foq6XN9IzQ4pJ5lOm+Ir/unL3GMpOVSNh4HBWwTUsUtee00PdjJYt
hn/T+7KtHgNyPS8K06mP4891y7xxSRkqSSxRrBsN/9TK/ZRWMpbPoa5m7nvtc+Zt
zh6LKx6EJf913NLKZ6163xpRLBpyCQg/EmwEgzfAvuWW3YEibnlQBmdJBtVXUTLo
j736Nf9bndV+9z6+RnU/Q4qSMf5MGxHzbFT+UWHVkdsq0XbgsW3kuMcynGLcuoDo
VKtGLKBFGlqbySjFkznfXv6uPIgfjDbPLIx02JMaGC6vxkzcwG41M9cKbAkJazUM
UX5Rs67kTngFAXXMcOX4UDDIZwx2Zg2g6WwLrJBfISTioTuvVLfIwtlvS+1WZpCZ
LXMB2CHqXe/i1KzTAxnq9yx9dRxFIXla6vhkfx8gJef3JpRTX0S3Y8UbyjJCYIDG
CNVCuf6HSGA+L90jvhCc8hyAmcT6C6D06C9fHQW8uuUVQA6t0MNOT6I4CHBfDQ/Y
eJYjtu7Vycx1hiatwTIexrDNuVexmFnDrEX/PWEhheipSUeUNi8R1KiNOh4NGpQ7
Ax+BaHM3AxuEhfFH/mvguFoqQFHP8qzi2jp804o63eqHm5nHqRQh1AMABBhWF3OC
gCpj0lnOxGt+FWKTtvgniOWROWByPALFlpGo0mi35sDx33HxZbaq6YTV8Lz3P+3P
rv+ZMnRferSCBboUbsu0shU9QZjbS4ie3wZGjKV/qQA99Yzaj1D6sR4MQWA2RV7v
LzN8D2Sjj3ep57gun1T/OM3LgWi97kyJ0FQ0kc1WkVlrTC9R/3Ba8t8FWPLi+H2V
1bh+sRP60fRpjyQo0iCHdmAkaP3HWhKtlcpZLY7qmOz7+Sbb+sNmPbikhqRWDx2W
ByPrLU2plqTku+4UR2s4gOtA6BLwhmgi4wCANXn1WNhDVhbhSZuY9nStPSSvPfQl
uIuwC+77AHF7LJVbbOTsZvsYnXhJrGKjvk+xyEFcWKLDmvSX4JfnNdDy7sCxdeny
XP+fnFrfVzZd0juVv00pv/ZBsgCJ9OBL4C0MnaBVLcGzJban0BtXHCEg5DxJ0yqm
N3/Zq0rP0offiMWbCw4cDubbdmsBl0Cs1DPYz7hu6ms/iH1gdb8wXl/4PcmCb0Gw
XkrOZdRbkUPRq0RD9ctsBreQvvrYI9AoquQEfx87h3+HzE2nqfXltoCoqp7K2+SL
yAQbChot6bI8iG1cOvAx5T2T9MTTQ73NoA16IWCwdie92jecT+SAZ0dOsBr/4XC5
k9C886oFVXEcUW8339qo92+r9Exl8ULXjCbACWkzRwV2x4/7J4p2Kb4LyXq2EMDS
JLAKtlZ8bTIBbQuPxyfoqrBTCifxQDgegA/VOJye/0yKSnhB7ynMe8gA9OVcmnFX
+JV00l/HkPPLBc6SC756dMVP8GGrrjJ4IJXMLDMjRcVE/MJ62jl8o2Y/UodthR+4
XsNy+2s6zJv5GZ3oZrBrZ7Vyi4/3acL7dHBn377p9P7164EJG6PzMami2mjxhg2p
4idzWP/eHF/OQeVUFwlD1wd+AhqjQJzCGGclEOCcHHYNoZA6/S2coforoljAbnHI
U0ImkIGK5KTWkU0HJM1OvnDIX4lD9RTFoFqZP23+LpFjxk86kpIiDPI+L1QJEx4v
Oi/vffL+B5R+QijaTovmnUYmkZvn2CYx+m8wxtgBmtpWFG4BKc2n3UVKZfs9tFid
fNKVVcX2rLUsnoi7Vmg5NONjT/TpMi8c95o8fsljc2IX5w/kj+j7pCTk3aI68J+w
eNarCPFtLEgh4fi/4tMpSEon12vtp+xmPNXz9eaDPwBSPI7VzAMw3MmX+UAedkm7
4V2j2urm9QJ7Y3UQDs94F6o42UeIifgfJocQHa747mowt19NQj5oHdaiC+5YnUGX
n+BTwW5p8A/Lam/IhHWFppX7UYPp6NnRVMKg/6+4+yrbrQB4QKz7NKjSstAGnTg8
mvirdmCZKgwITCm82vLuQ1nIqHbtX6slJXUmjd2erVaHltZ0lsmjTBBA50bFPn3J
37fYM2v8qKKPveEG/hUn3ASgSh522lCejqoRywWZRmiqTUKZ5tRSAR9UBgeT9q0e
gVh05bnQWRihh4Nd3tFyaTcIU+tgzssjwz5E+fZUK392GiU17eDpbKjNGP7hLOlv
3tk52qoZvl2ja1iI0HHep3EbxzBhUvQASDmgK9Y91ffo31jTuf6nDaweCr1p2vsj
Y9O+sW6LD1G55Cnes+cHHdrWAyu+/0Tz3dYeoMj3Buc5Y16LwPiBv41GcgW9KgF1
e0qKLESHWDUsis0dlCj0z0G56zbP0EMF678n2aZYJGycA6ixsNPidiMH1g857hmz
YAZBUzZpFSbIj7teuDRYsi5lnjLwXpKGjbQkh6VdEuD7phCMCTzHHFkxg5BMknIG
Ke3vQNynwSUEFbsg8O3630F0YxHeaBODUsSr7e7PV7HUNQaR765wmfnk6sDawUPF
oy0JQaXheumokxpdQLzXAo2RGs0M5G1NJvGRq2hZX3kqEiohu0hcCXNYC5fjopUz
HSoe6aTRB1FMeAm0NKWqrxIJ52Z5uBzphkHXWC3MgTfM93fBfH7U9qJVVuOhDZHO
HFbWZXV8b0VkMs9F+QD3Gyhi2mMhcxpSzYk6Lrks9eNYGqUxoQvHJkyJP+Oxxukg
qdH8V9CXL3GTnZ7ICyyu3aBc1IPoCCgCbdaiSODv4GZqbvFJ6xDNfZbCJ3ngQrxE
Jcf01tNFVYyMR0G+ZDeoGaIX3QPhSKL9dibPmYhYeS4i84F8SV3eKOAQxigXHUPh
bFDboEn+d4EsjI3c6albSU6t4M29sVINx8qZ3wCWBXLHGPX+KyngSscjlMWJMB8e
SQDzCyftTNGAJMAP8LF7P4YGK81EkNwU9tra84//J+PnwjPwDx6iYiWaH2mWGt4I
OBfPzvNiKhGyYDQzpsvV9IWlc1YaC+HXmyqQobbAPXq3OFulvkpyhz6tmommjfZM
/9/cVuSlYPKZqorDJ8GNyIBtJR1DwroNlZlOiHgFulQwfjffftAT6WyF8/yzIpUF
fIEAx5rRBmTLxcCQd0pwl5eS5Pkx3A1pNtMfz0RmRxSYQbp4TKHZcWvAzLQXJ22H
TL/1S7PcYzPEohINCbVgpk7fgPye/RK7QkBY0ethQC+RW0gRtQLAIc3rebwO24R2
eSX8EbFIotAU6pKzEIl06Zr6fDXJZCfrE+rCNL76tuw/OusHhV3rQoHNQYpKEeaM
rOAiBrzi3fWo1kXjKodlMM98Btritark3sKGuLuAN+OiNJNd92BXivdT6XHTbwnh
36eWhmeCnv9OhF8cMAe6xV80gUNk95RzScN7rX+2QvN9EAJ8FJsJW30WLkcNGn/B
5Y21tj4oyIFe9U6hkxWRgTkNsTNXzpxFU1r3p0Al7hDQG9ZEhE4nIbo+AlnZK8Bh
GII0OmHQw6JWBjBd3JdZxowZcDUSA+FclP1Kn9WwwAMEoZzbC4O3IqYQT94zFCOp
e76GLg/wLbYG5WUemNFPaGJ0+UOXdJfo46NFw139WnRlhnJ1zNDfMVQFMAxEBiG0
eLKX7OAgV3mLkwndM1A9ZwhWM789cgAvfj4IeHy+QgWo2jZaEX+itbESVrAH7owU
6KNWNK+N2D8jmMQSOjqOTB4DDHwrNVOUDBhnmwibHot2T9XSAM0m45+UNXc/zLfS
qW+ldfD4Od1C5jPDuokYQiRuRMT9jS69Cchz9paHOv97NAKOskSATb+FUAFr9WuB
EhDw3kj5BwiilvYGcRGstGqzDikp/SaIB7CMyJVkqq/ZUf6yt5m7hSkGpQJyUt6m
ueQeq0e4lCrIPTuzAsCRI9m9vL2soKhre3T8N3/ENJ6yiV3VuvERYOTvPuHwVK7l
byz/Te3wZ7vT1a1Fs0iin0wHeqWhH3mmeayVNVVhwtW/vLOcV0E8mG46DeQQ2uWZ
DEZhkDOWqvMTWmUtcxa9sTZZT5A7O5R+JRKi78prqgyAEolrN5l/Z8LBh0ySDaB7
sd1C7CUcpb6SymQE/PzPzGfkZobm1arp+LKG5+tXzaieCdD+i8cP8x6+SZCOZQiH
nO/fjrb2whwYW8eW2tZHEXRGqsOxKqUkJISpW8KW7r9IXVNjn2O/+vZ2gr1zidfm
teiy21VR/oVcQA40gHx1A/8trvYDRZ+SO49yxJv8bJltSy0KfHvcOW0JZ2m57Azs
r0f1eEX4hIe8Wwhg4rHoap8vkLinSLFXoOr+DdqUtt/PSMjTzCq04/TvQJ7fal8y
BoZKWK6mXLwk0Kt69RHh4gX57ZKpS5xoDhvxv+7jPqN5MixjqhJ/II7m9qbqIRmP
sHy6jcDlbjwKr2M6pUGP5Lsm1NqJSQ47yagR7SzFGFW2UaK1mc04SmGeM3T9hvP2
EhxSavDlagWxHkbJTjQM0ptL+ICMmO7Y+GnLsWty47UVrnlecQpy8V0k1orFArg4
ANi86UkxPwOw7/f+OXTaapI0LOhPKu6AihTZ7/j0MLcybBbnSfSr1SmJ+PolyEeN
qjbzr26cP9OTEnkasX05n8R9PpAE4C296NTc+Wd45ZcRVED4GOdOJrdMTSSvQLQb
7EP1d38f4zL8DHpq5yUy1MjJYjNeu7gNtYX0C4FaQirDOllGgaVVxmmScUwDp2q8
HQBa7ZNDJA1365byO9KUTwKJFrlBHb6r0ulgWDexPKso4+dRLrUAOoHprfI0+EZZ
kqP6l0RlEfRtF1lePl3grTO5TpQFEZxctULxUEz9fYbDvtE2Tq4L241K6WYgaZ8s
n0PKWG9jEwSMpAkI7R9pqDqxXVK70WghKlqmm/Sfzd0Uh0y3TzA+B9AA9FaYJruT
kScBR228X9Sy/EPmen8eQZlBReaRAcqHRvaQbIevwcY3tKqchj3cE+xR8MkxlAII
ASKEB86XtEs6q9N/sfK+FW62Cn0DFCld9atPy917ym5mcjOJWsiLf7xKUjma9rXg
O9J8ggfliLth6AMB0ad/YgueNDDkLi6lsY5YnHNCCjsQwZBANJXBfe3s9U5wm59K
6EjroWVLsC9PFX7URznOkcyGvsg4Ly94V+d/fEbuKMc/W4rtglWwJYu0VqFcfTfS
40VRhvHIwjZweQuJIX9HifCQqxFxR1zWEzkPZEqEqh7t4YkzBqGFbS0eWZ3tCIki
GNh/OplNea7fi0dcn7j643/u1R/ywRob32bKHhCGb4YFt5YZBmzpkNaVxYY7+qjg
pikS6reyQpvNBSsdtt2TSMlvZ4gmsYUPPfT0zK8Zth5MA5G6cWc049hqxIXTzlSK
+5TgLpNxFka9IUYRSa4rTIIar2X3abx42upMatT0arzooWlFEpKmap9ih06kh2oU
LBDZfXYyiqDeA7VAyhGvKHlyKa5JXP6WO20RLDaDrWVYhxGrTqcv5b0ksVqkcFxm
2Efd0pvNmgYzGYTZa5cPJ9tSKOMxgw2HcnaD7Rgf9fqlzQd+lTsXCt06tHBoq6jm
4LyyFv2ipUIF+jc6rVXVEU1nYaB6EMHKJyZhktZdwSTdtAf7PE83Dr0pK4YxmSd5
2cAkXOiv3KViH2V4r5CvzBST+iJCBNX2abciZuhci3j0xzYcXDJxXG9pCBPG21LA
UudFqpvKqx3S9D0Z4WKACJO+KT6Ni5S4EHAgFQ8boDADIBJfCskLpJ7fucsdlpmc
VfgVPOIax6+f6rX6+ntPUf6cv83Kb8DU0jeeur4MGm8PUhPS/Y2KkD6FYrdc9YkY
WxBtYU5SFsLjmaVc/d04SdwUeHOZmjH17TrUDZ+22QCQYlmE9YVkoNLINQET2ASq
eerprePVYyGX0OSLDuv0hMN+tr0NoJ0qHuVnMEfTEs1spt6ncx42vJU6b79h+x/t
lLG6/CVAxBiclWSBrPOENgbs5u+Gvqi2dOao4LoGidZ+N7WNphKHlyvYlSAC9rHM
ZiTg22QcmQJuR2XxLN5O3hPQv3//SCzppsJaCsmdwBzmzdoH05qQwZRHvXbyu5RM
sET5mlypI0Ev8nHQF/jUn0wLfxYW0lz0guppLNYBnAJGdbHu7Vj0ADW3M/ypr28t
Ke2OQzMPYnbeCAONHMTSFh0kNzanUTvlufc93AH6+gK2RGVPWl9nVscPn3ktz3iq
XOzmbgxpQQ9qeAJiBXwbSMbWXF3I2/By7Ry2PzL7jLgJ/NYzipWzDppxskP3BPOZ
2E9ImPDDSP3YY64r0ANsEcun+ZiajwTjoUvT5pEc1wo/LiUeGQH9TwSejlOJ38EU
7FiEMXMBqlDwXK6mVvKJCcBWVUr9Lbo7SrpFxjgEOYhHmvbPMfVmfYx1BBkVHnLY
lsjL2qofV2KtcR8dPEGt6x4IV38ritDJ/FBzyB/T2ySgvkmYSVj1RpT8jEHyGMd+
kJ7mIhuThqWicsq6NXF8HBZMSAfgGPpTazE6hjLnOMWcXtKBpxJ9FnQOuViBpayS
YTHq2dG5SSy0y8kixI1PiQqr7gMjs1Cw/kpWChC4i0LTB/bOM2xMf5MPvFdP5y4b
aGHvISkJ+8j2yiF3pTgIQX2QFC+G/ZJLVGcs+HI2RP/kDEHCudlFPOhB5s6DxpKu
XSg8Hl7gnW7xv22jjyTt1wdiaClFZu0onhx5A0J78r1ZPk2Km8kT+jzHpffGKmRo
o0behzb+nDPL0eYY0RV9sYSEM3C1RP9OxQ8AHkbhiK70JxFM87GBra+RZTebcjpW
VHDXKeyPA3FlhBRKd8ZNHBbulK1J+2Tos+gLcWtIpfwUXChjMkzFAKBRorDZfzD8
LNfgAHMH73rubpA0eEQX5aattHeWcTekYklIN4n7siVCqa3e/7ipzd1wzncEzifs
NFQdhrAQRD31G1cvUJ5XBlcAZ0DJblDIOjfaf7G28e/3C0Sb4Oe5Qi0OGIh7/dWQ
+At+uqxmuAUs46/2BUWV6KkMCKKzLblwLY5wOpbYbGzE/NrbyVjud0y3CWAKLvRl
z5u3yKIyrp+2cC4gh2D6cO5/aBZZcjST+99TEoZ/SfzXxtBNuK+jxfW4A06uvEI9
hhy9z7ta5lepgddkB7izV4EpIT7RRPD4x34/tpi6w0Nx7wfggNy2ACTcgUMWuze+
EBdKlPH4pAVP4INFK0Oh3ee/sqdHVSec/mYKf/fzTbUAJky2V6JF56e/iy0sylIe
Hm+0G96WagScHhMecyca6B8Bvc/kCH2SdoYeIMMTmfZFZiryCTGOnQGL6U7h87Fd
DYYvlMwG/9mgNHUDPIalm1LjZHilZtJS/bpYNh83NbsCWMSbt+UkDVYpOYTczfvl
pxVfBNCCE0Sx7e9tnbNWfxwiVTmDnIzN8DLGOhTlQ5wErZDTgUSI2JC+f+8bi3IF
Kx9jTE0qGf/vYe+A3QZqQSTGnqtRkUI+0IvJAqsu/Hun52MWs2E9Hw/V4UVuLF4r
TXkTQb5a/b1Xe1WsxpgN8EqWkLL3HUmtGia6+ILn3d35tVtRClR9XCTOX28BrnYY
YGO8kyMuYUI20ZrvGlBeh9VoYpi/x2hqvqg4R5vYgG4J+zDJ5HJ0HUgjf6Q6+NRU
BKRmCIaooyL4X1c3gd6pj9JoMG8vvnYon49c0KQPyKbEfw/b3ig3FeQ+xDj2U+R5
CcAscEYKWak3sfyITbVUKJ8dscX4w3gpL7dJ/8c5RLd66rFay8CI8x5+VRh+IecE
+VP2z2/diELQCJnsmkJNKlTKE8EKoTAEQVHLYetT/V9tN4ssucwapC7ukVZQjCHO
H9+LvXiFyqve/6bt3NuqoAHFGI1C6wCgSO4AQuYtt01yhHPjwoO4dKITufRMiHDC
sO0PtptM4mB7Qbt/B3bIhdDPpTM5d1EREgiqOszcyeoP6tpC8Gl1DuNazL3/IZ/5
X4MuOVy+DHG6wLO7KMwVoqR04HgzsOQ67Q5Nc/qkn5X+DLNiHL/oIygk8ihCNGV4
DkCsIG28oNoBCtqimHKc0WZeo/EsF5fC+V8usC+OyHVh5g2VPccbcSijfWltgmRF
d7JyB2ZiIV8LW2LmDHypA/S8/uzUz8q5LXzclHN+Ww8iIbtg/SlYzbq+ynqWoV0c
DGnRw9s3coBBFSsSuuPEMcaxkS8C3yV7DAVgtW/gl2cmsqdeht/6XZRNrRcejswd
oe23jrXkJhfQG1rAPW6q50F2Bpp0ra6JBNfbhXB1RmHcQzTil1wtli8ebbum2Hn9
dF2Paz/VR9oEzMqTrlWeBd5xRCiijTX7rUMZsVJox03spg7uJjegIQsUR/jezjG0
1KEDfOdGeij6er7G0PHT7Cj9/DixvcsA6le90Z6bckMWVpF4snEVvY86ZMVYoKd1
a9iaKwxQ3SsLaNdnX9Z+6lyNZe1awSrbs/lw68IN1wNNYsAvy+dNvo4sPIudvus/
5hVl1sXxon0xvWpaIUTCTJhrMthaa0t1V7CUMsRt9ZCSetGWd+vklE+S+S7sv4Ni
TLmfmm68yk4egoJzKD6tNvpRK1F0SHuP5N/SSfLC5be4N6WsjgKrZRVbwBnSJSpX
zDFFipIPSC9r3asoGjRYyJAWfvbgu0c2HE9lWM05gqnl6i4OsMFyaRJw8cNQRpyf
66na9W9+5QxZc9twMvcquBeCRRJl/+nVs+dnAT/4wKioSoAVUJvkmJASQoHMgdgN
nhruCJakBri8VEeSQXHqu43BtKyU/VMUaH/jv2slnU2kyUUuSuX/5Yzj6MUixVjH
RyA6IRbYdE3I+r1bhQBJHNq0F4ZCVNSzEGqU5UomaTlUA7WFmS987sO9rxtX9fTR
MdBybBUs2ipXxjNyIg1+ONRmuc985BrVABLXR2VXFooCRFRw5Bt2JjrW2xe3KsTD
a2M0+iJQfg9/y7dkVQ4OBfXeOzSUDKuuiDU4KyQ542huzMVB+TPr+5XGtUvB/0sj
Joxej7K1ei3Sz8pI8eraoFMtTSpuA9YWFSapHWo5wNHyBVqPlGSUmS4Z8N2kpk3P
yByyD+fzWn7lbYoZdjqLT2+a4ORToU5DXDaKlvF7G/sj5hFSLFcCx3ik0h6K6R5S
Fh+Q8BA5vhSy57lgWXI4jd5UdpCeb9vMY4pR8NK6LQcP8fG0Xm+CBDLuFiGbOw+8
cR1TZ4KT1VFJILu75lOSXZh/dwgoVw0TO/utBZsWqnfmaQVZ3uCK6VKelrSHQTgH
qQG1LBHmn3vngODcovyzLidNDfJ5H0Q5YOUZ5tD1p/jp9ny09qfgS5iWUe/HOtZe
zDTXlxSap423kw2F1RroNWjSfV1fu/+PbDhvYN92kFUpeUhjU1FjTXbsfT2UG2vE
W5h0SbVxGHHpCHkeX9JdQm72nGDjwSDAz7EO/zdYKYW/mhdAXdjmleYlBC7UCcZO
8aO4unG/tFSC7Kw5ResaPVsRpXIuMs133bH/NC8//FxOA3O+45Yb6M2Pb/ySlNtJ
AGNOomxU6/okGC3u5XSv1EsfX7A/yXYWkRPgYL8JmhMegwwD7HwokfxsjwkqsxB6
z4M4VLzaJlSpmGUBAxalxB4AwEp/cAJOhWLTPvbI8OU9dobrFJ2jCBzbE6SZVBUx
Tm8WS0aXYNtFU87XIiofQsAaCKebloyiwbE4S8e/ye/2SwaJ/p381XtFRVbTMVm5
oIFRcIv9KKdqFZ9VpExtRCfz+Wi7/tyOaMaKyzWbmoIzTndj+rBjg5OptemZQleu
XmjSb6xLYzsCow7COV2eACOqO1jysd59WgwgnsYR9gR+a5QaEQYpHafJZ0AQzVCz
FkumombQxMUTCJIANooM9s4FglVHveKjDo+5Mda1T+YvkSuTNpVpccdWKu8L180y
dfuAagIMIOeVQyFTbWkqq/4Z5ReFcRyWcVkG3NqG4Ab7HOhw+0tKwNrsExG2OJFj
ROrZKgEUiJ2BJ7SbxJgim4nu4rbJ8OAS1O7k5Ej36WbIrRzNfx4fQjcxynOmddQY
8v2kiTB+1UGN3+hxto4wFkdKDn/q+SEyhicax/sqQqEBZliSRiUOcTTOTjJuZp3P
87a90kBnSK0CE94vDzU5bkWLJAciDTtx9Dz7XHgHllQEfdg9TH42cvEXg8QdldjV
SiTlegBGSF+P2r5bQg8/y956xU/ruD9O6JVwGS3s51c2KI9z3O/fMVbZEUAnmDZF
uT/2WzGZ/CBiqdhDrGFMqA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nIbpsTIn5hrNmlpeArDAZn/BWsq1RANRCEjklLBAQUUvISlVEE9ITdRj6mazY1ox
PD1ulVwY07Rh3IFtOZRH8SEtXbmCW2YkjUEsnWhD61YsuWz6aqWBFtM3VJt5CY6+
iGOuYX3g+LB2AhEKOF6srpbAKundbSRnAxyeZDBh8yP1yM/QB2KvNH5sJTUbAZlg
Hi0OUgc42Zhd67ILfTOedre6uvboPRicPIOGFLcJ+0Nl1QkovDbYNGDPsBH0TyMr
nf8A8NN3JSq8iDaa3aV/pLLRiinJ5s3yHGaN84BNwB+IchIo44ifMxDnYX0Dm8FC
47wk6wxLq1b29TyUQvUHUg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10640 )
`pragma protect data_block
hshfky10W0/RP5Y43vvcfMdyQ0vHNPtb+jDUNd6fGlWtdQLR2rUlj2ja/lCUKj/n
8ni99VvrvUSdWvE7gbz53BMwxLfhYTurfzG5Lh1DImINFGHJFVSdnFrDGv/4adv5
ZiNs+fSznn+haSzdgl6FnbkCSdunITI3j3NFghYAFXIDNeQg+c9FnV6LVwe18Oxc
C22Lfw0ki0449zlqRpiVA2hNUkmqfR5kxc32fcTgLq3ISTBU9mAXe3JU7bIr63ZV
4Y3MTTwBuj4hqpx98PW52u9+/4G1JsUTu47latqobGQFVGUaRiZNu6Q5dMHAgFKt
Xzo5gIHps/dCkKZRlQ9ThwJj98wDMfI+FpQgGc5MfcXhQTSwUsrQ+GOHtDeFVfIo
Bwm5X8OgtSt0Dojf7IQKb/AK9v2T4eVIhufdb/2SDjLop8OsGD8S8v7gEpHcf5RW
pa/6Nvjxdzhxqg6fN//4skFZLRbBtJ1dzWjQxYcgtvEo7ZT+sgJY9qq905XhY3C4
fouo/NUYTUV8S/6OoHSpJHYRt9LrCWSFwwZsNc8Yl3WNK49f1FNgjI4Sp2Yi4l5x
SQ2gBsUYTGpZnAH1m5i4tf68zamQjnINK2uJ5NW+voTMswPJrc8sNctajRSc9+32
vaG2lLDcBbiZmwDRowp+0jOlP5WyJxY82dI2VD/ZGuugnVzEQcu/1KKRZyY60YKz
NagyKt3NalnCanHzqBbW5nDBMDvuiZHxgssRYB6aEtAzjZe1+F0wt7ng+TzMov4V
20RNXMRJouoxLaOONHsE/ZR47XhX8k1IpL/xVmKnTs+IhYrZeACOcdffJbpyWFyz
dJdOxMUzIUBpvypGjEquTJAQhJPPq+Oqn/H1dmQKW45IFXmF0ODVIK6OFPxqdN9T
A8JvwFZMNvIW0UjEl/haCKur1/nBw3dyrsbyScYFvwhHtXC5HNZ30SftX2/szWSf
7j+/hTDn08WXdg49qC3O5DGsCbzTdfsHrKQr52TTsRROeWsKix2Lk+nVlxrnsJ3o
VsRRAvn9J4f+dROSDe9Dw1qMhzylgGDCeFXBO2haoImsj/oF+Yy/pq3nldzMQzUw
JlH/ZedOH4b2SerZzHRpyHmYsdwg7xu2CxUGMEyMV4X57L84qWBcPSKcVLqA3QzN
mVawpRj+yqXr/iPvPITgk0blFprhuzd1XPiSkAWHhFuZ5L2KSg/xhlhy+iVaF7S3
oPz3Aqb8osBLr3JF9fLs7uCUrseHNHCEWdMCr1h2XYmL64snKKOpJ074lmh9UpoP
BAQ5++avYogyIha503pWetHmAdKFq+z4azKmGcKaOG5buMH0mTv3bTApHX3v1vac
bd6r1j9XW6GQaftXF/NhCLC3jdijM96o1HIvnCF8gvGLiH3N0FwCepcw81nYta22
dCOebPXMDgSgxv+Xqqmej7py3pNpbkW6R48zUlqdmxtilhe+VxSWfdkqS18uUJmF
SL7+pyQB+ndOqPSRj7sYyPcdBatHD1B4c2j8YWXA3KpYfOcg9JyNqeT2g9Xq3oDY
GrDmY1Btvnz9CNktelkY5v6Of+JEqFLtjYMjBxxYApBfsU1/Oju1mnUKqwB0wtDP
qZu3qFfQmbM7R0GjXIUSFCkFerggOpwnxpWWDKS3tMIl5vpmVdNfmyg6FETOCAIl
J4r4x0SSlBh3BzSUNmHtdDtHD9+2IqJJE4sMbP4Plzv6hWXLiLOGwa4a2evhOM0+
SGwc8CzLx1nOJlOkFRmoVa+Y9wL0Vm3ejnRFyS2IUpHcfSy2T5oUKM5p99+OGCCj
XtpPAMl8EdDccUwdyymG8Hqz0I99XkeWr78YrJ/gT9f7xG1TD1O3SsciiA/FcJ5Z
ePXe99kvtcttFFbbaJm2i1Q0I027YAmvEJm3QReYRS2oIwQCTfqbS56RocG721uY
/bc2vDg7D1igMje4KJwi0fK/gI+7rfnIpZnuaHUyZ+oFhtRwPNlscFr9/u7JWf7N
CZg17J5CeHZ98sZWQ1dg9vW/0KVE9UBQeyImX6mH7z08DGEPW/Fl81srsQ/qc9kJ
FlcO69UI6fZ07A+A+m4Z2O+voAwe3wkpZjf8AHF2FCGv5/5xZSHYv8rppKCx4gPp
/pW62VYCvXVjxpakwxsSyG8/o/ZfapeJKzugHDt1f/ldk+e8QTzJkujCCdPqXJe3
80+c7SIDNjOYGKXns1wN69sncueXmFUz/T42HIQ5bvi42ttufbYZCCRz4glBTfht
pBpv2kGt3Fo/3HxQWcMPT1o8wx0vBVRZSmK3y6CW3722k/HFtiyg6wGWPyxck2vp
UiH3ubW4Av5aOOEprIPqDsU4uaPkkknH+SK3rqcif0yWPUN+AY8XzjG7hHwae462
Oloic6EAZ4hIpfPyXK/BByn2gDMV9oOk0lHD0jw+5N6xI+D7h1z8z+OKwqvbd8iH
f/y86i26J3j9g9pJEKdZZT66XpZhGyamKoOsLqaa8rohAVRMkghd9dN6RL2ykSl+
6UmwhiHXBjBFY8DK0AsJrfr/mzIyuXjraU+mhAamZouJovYySD4tT0I9DKk2LpwZ
GrEi9vy0QjRxfhBroqUXbV9pGsvmb+kOyBPibeS9nzfNYrJwz+EQkVydzhVaQjl4
5fi/CiZ3BFBZjsNGug/9hx8sF608JNYq79NMsoRtmdsRiUKf1RBXEcB9krIFti/1
wEuYctKXaes4bKmyooGMtfs5G2Xzogq0+2j+m7Uazd6m16R1UBjPb+HyPPznStAm
V+gv5bASfcrpwkd516ruMNfa3oqmKCv/pEeZPBWRZZJSsU/HVuST33/ru2BvG/ln
ejY2wk4L2x3C3uuLhBUhgKsH572B51BLlF5ImjOuATGk2tLaHb00/HxIsBScqmFM
RoqwST3YytySGBlSRrx3Z64l/mOXENW3EB1iOAQ8Rc5Bh0scCXDgrmLmsFqlT99L
Guwkjwv2qrDNl8o4osCA4A5Kn2JH1Pnx/TaXxijGQoMwp0j7Uf+48wYPAMW+6QcP
TklWLGAoQqG8hdrL+cVVG1GQpF2UkZk5GpAVmfmqwV0YBne8Rzx4OM7Wl/wv5/sK
4p1Xy5Dt56Ig9pRCgv2VYB9HgcXEJV9nJc7NtzZnrjzrdeehtH8NGZIw2Ey4YJp+
k/7rnzXLn0ZUtdyTaxWfY+0YiGfofoiB9wDvghT+z0GwSmiF45Tf18CxAxKtPu2U
kJrHdvwcqvWJXk+fZvrVTG3d+vof3GK0G/BWQr1yqOwrmHERM/qczKOf7fnKpgdT
iJTe2bagOBexAPx6ShKCisbSX/4OyZ+A8oJMyvX7/dF995PXq3zVKYf6iwvDPVKk
1lCgoCTRWnxG5yeHaq9Pt8T604w2D2i/xvAsOkIwjjug4aPMVt0OBtDzkIDubowG
hJtRXqAIwLt/OLOgnS4x3shHQToZtos4PHbaXVAoJPzKtCAf8NjfIb8PJM2YIEF7
47ho78Oa81SYmHLubBQ5H7j9yXr7mQwdtwQAW06jPoVRXHccfsM1T4piiWCp//Br
71NO2t5ITfggJzVAVSS3AxAmvAIMulHqNjTAl9FbxW2r+m+a6+v04VVDUib/grs7
kGMU+u8D6iZu0jbOMo42jaSteiDFmv5UZrSjZhBcHTUr0ivQbof2lKGtz3h1Q0Cj
M4e/SJko1OpzAGhSdyHzkPsJR4IuklKDmZEAshtmdVqLHnnvGixdm+0MW4uwpLoH
LG/3Jv/7t7tly04gNHz73VZNeLYLIy4HjxulWMT1zFQflEdYBfiy2/B7slPDuqq5
RW/tXobt/SK/4IJ6uitoeOUT0uIKGr8eIM2eEXJ45Sa/e2PF3lEvLI1prYefzBz5
XyHQEL84b1XQEj21JMdFltX08W+BNf57gaZM4Go/AJmseDV21j2voqEv/oG8Hgak
IuZ5VxdVzAezRbsGayY0XO0heVKm1s9unVn9tskT8uc8sotJ62MfrSmYpsC90SCM
zriywABPkbOHdF7aO0U+hJ4Gp7CT/ZuYsCAXB9eKJJjedUfJgYMynuZEltzs1rtP
uivvnmYv5idiXjVXbU0EAyxhAxAvgVmrVzB7ZjldxDpIhoO3f1RKRsB6uWDaWRko
XJeVWY2NDhIP7ZvgodJxLdnyWyozDqXppHJBmDk9OyGSbnd0CWxK6JK1qbXj7B1M
vhnsU78erbwrEYWCuLhXzMDjEIo9YlqPbqe1VWTAQBLU2U/oJMyuv8TmZ+LLQu1U
/3phYLzevFbTEoY6ZBKSD+pa/QXatxtkGxQvTM2hkxun6s2UrlXEi1+Vk1VRspYo
+bWFXET/28cGXdl4H/tnR8285m9rHVIUnfPsvp7qtBWvXM9hG82V2CCi8tCXe3TJ
OfE4uTHO2vwxTuN5MbwB3nMXjCTBmmCIIBjswXv9uZw+XQIJ9Z9FPlqUlatKtgpZ
tt/tNNpJ1XMiZJooEppcBd2Bd4mbclp4sSHg5NZSvvOvPQFNrbW/EyYk28CMqo9u
fKGLcZF911dF++KLb/2bIaojNsRcWvdFaEHJ52GZLaVBtFwvdcyYQb1PLgTimqga
8IS+3REk/Ov2mLc8qHK3qw18oRjy7ugndXel2gLZbuh4SBfYcvksiv/3+KPNTp2j
2YNIUcXTgFFka7MEpSjyeaZQf1GfS/Aoq/iMjpbkZl0MyzGh/7X1mZoL7Iw3WjfJ
kauG9/id63hpMP4wIu5bwt8DQPwap+lsDDPP7CMa8UxU+J6NA8v9M6RhTRtx8933
qi1tGIL7+8rFxNBmQnA5q8N44vg3nIJI3DwdetwAHCRs+7DurRky/YAjpX1Qy9Gw
iD1gKAlIv6OdoWdFmc4KO/V3l+5uquQpt4lUE6RIgfPRNF1RcT41UD3N3x/JBUiJ
T7SIXzdR7jioZdQH8Er7jUSo8gQqJenClAbkPia2Ih0AkJ7RNjnIneCvvCOhUBSa
Fmyh5Tqn0LX3fLcESM3s/V6u97QTVZ1LW8KNYg9UC5KzvyYAJiK7VHLKVB7syjTO
tMAX2zjh1ybX/2pkitJNANaUGof1c7TGd2K39Y4erUSasY8wcDbrTV/aU4isCxs6
On0wBERRZ/CpXqLN33M2AaL0+5BYtqAwyEGIzq32e1H+YVeCidtYcAdoYxbq3twc
2fZj1hdSP/4f9LyD7WyDbZ543YBq8JyWO+31vog0YqhcsgNMO0RW+jAvLKny2vQh
eg3wjIcNMi4+rURRCGS/WzB4gR29z8VFVy9LgMSxRxVOsPKiKjJKsv0a+is8Mp0I
2Ovo1gHc8a7P93AxaaXlQtXzaizSPc7JTGcqK0HlkNtd5anWYHaiZl5NgVieZKJG
GWJZzNnjjUKJeksYE9OIGrhOCJlyIwdnuZ5Vei0jWkUvFu3c3kD+ZAlWEMAzJSXK
7BoPCYlwtFXT9/QXqqXT7+OgT18kse14u56HNnVgKcvF+hQ6mc3Q+mrVxI+HNEzJ
Y0XilImDr/fT2bzvDL9KzQii9E7LAO3Nz/PWRWomsr2HetJizyEg5sHWL2HEn8e3
3zoQeHpa/W9BoqDcSRXpu/s6Qot9eiVowyRc2OhE6gPYE3+pQ7+M16jBSnVvAnWv
nX86YMYX/PlDl+K5vPZybDxXRM9xgPT5G2wtNYgY/3/EhKP/QFrUdrFlL1HKBsSa
+H0qcwSyZz1jQQqEBuH2Hj1wvVshgb3D2T3sOR486++EoBOFWjoTMIhAd5Gnj2Y2
r3cI/DODdayJAG+6XoDG4HE2aPnFThcGA0Sf2ZMoETxjJOLv8x0VTAEA5FL2ozf6
2K5rbC4qFPYSNv5wAMCI6ne0XjUEjru6lsHQpnDGlcxUYPAuxmAl/mk9PLGbxujh
zilp02YLtxgDDJAcmhm6S18fF7ikHGG18YqWdcCWL8r5SAOHOpMiVkh1QCjoqIEG
ww9VTzCTEMghYp0f5NctIqd71jplQuUOqw1zpHudGTIz7h0RTzJq6B4SXqguzJJD
zXEeO/nbp8qcdYGO4zprOkTNi0pCaFf1XWAYRsc5rTy5/SDSYXbFT8u+JGBvRpfx
ajJHftigZWKqdwXF2sPGyb3rYGFYyDavFK8U9rfi/aYShMrwWQG5w2j1gDoKTbtZ
Uj7SGHcivjvGIEjt7GPxp+DeZ5mP3rRrQmeefcZFsiUA5R2z53OWABi8ppZCmT0k
NNeraejmC5QYtdCuxVjz26kbK1CgtopB6AT9Z64gZTdgXgOANqkFRwwwTwaKF3GH
C9seE3aCGA23oe6Nf3GGKKjozb3BfeR5zOrxWy6n4UxY0mRBwuetTxWEuTSVhLCD
vEBI7ad7zahoHY7scEBL/fvzGKGyOeTkBNlc5xzjzPO6qP8hgoftYrRpTVMt1v6j
5q3cWOACaJB6r1Sz5J8qQoBVmkstAOYj/Z+CG2gOdz3njMWiz3pp6QEfT3QvWN0F
i0Qv6d/sZmYgrk0+4grfxqZlbjt7uMv55jItX+SZggvDMM7k94Wn2A/FEEV2TKPL
J0ICB6gmdEEIzQVIUgPZg50DbJe2J0v5wD8xBNdtBHp08Kiw2DCiJbSuXQ0/bDjp
nh85a9mdt8PjYF8Q6kYVMs1DdANvu9LUyOMoU92OWNe57mEAgGd27zSIyChiGdHp
mEazPZhFgfb0SNgIEbALbe/M8O1LgENR1IeM+nNDkfY1oUD28vCDdgmlwdpEo0N1
lWt7HUTci+WLOCobSadTzrhpeNkTzsIPdG9gRvzygAwRLKlxRF3V0ZyKfW4S3dwq
Az+5j9iQKhJ85NSFc4TCzj8L7lxc7j1WX+oqoU6EFbX4zX8x8RTUXXbn15sxOEcE
NJk6d5yUYZa3+92gocifRLjYGdRUJh/R/lvsY56NlvCQfnt2Wfj91eDOrqi69rAO
fJI6KJrGVZqOHCTdmOc1U/ahz3pam2mgyhRhJZgOVwwA/H+6FsWlsTygdY6MM6Tt
Av8ndillhmstlpUTgb+Tgfs5xKOlDqyA7S1S0XvY02du8ph8i4aRuoNWg6rWCtkN
cRWeyOz4atqVQuLPz12nSRXNerfXJ17yrJLPEM/kyefJ+YZB1pnwDZkcBpWtef1H
4zEfYBsIgPOG1jClfDotlD07l5WFMKONtEplsW1TfAQITUHdwD87HOcm+KAuijx/
B1BD62/eEImXLBs6DVKaMGNx8wN6P4/wibUV9qDwCBfGyFycykjc7LFQvxbNrXxa
SEp7koxaT+SDs/hPJMOEsnzHbuaCSFTf4LVXfO9zFwroLWetUXvRb0HN/imKsn9a
/060R8ZmgbmBiZn8fTK30IwFjtJXYc0vpL6K1Z6GXz0pJ0OErsMRb8ozm/+9bNlg
5f8XP2vvkF0e4wwVXcsUebziGsD3sR8wQAXBngiRZ56woN+tT9kq3JXU6EsxYqy3
8LxvhOztqZGgdxsCUw9oyLmKCYG7jcTi3wG8wBdCF6QR4xN4tbBClg6T+QLVRcLs
ZyCDKsVgl1Meq33P1/t/MqiKjLAZtgLCy5z4LUQDMV/tNcrPOzqMRCq3CJJh2AC1
pIiCFKyWafCADDNe62OJQRx4PamimUutJrwEErKGptzUrYMysKArHtx/PCgRCUTg
bljXuVYfzmsVUu0hOWJuR1bza5x1W+V+ItGZsO77DlGlwETJrNVlzQKyUd7x3gDJ
dWQKZT1y+frF2WRSs7fFbzwIOdtAETV+1S/eeP+jlrxtNEZ6al/Q3547jNakVb9e
Oy5G5EfIY9RR/N6v+HVt98M+M0+0vkov7CB+dcvAi5xukPx9KB0Q/nXdIy5WVy6g
xbVZArT+564SLM6MIeTdRQtCXX2cf40NV3xV+OmpEFBgHW6DPskSFVhCq9Mj2uHN
ARx9ZY+1Qt3xP3jNJxqdIUoxCWzzgQVBkXkikJ2kvQ99OBJUvp5uxA6UjjO3yBYF
Lvx0ZzUmosTfk4q/h6ItyqjKqCxuGZgq0y/pdZ3/QleXFf5osxCs/ICCLpg2G4Vb
bL8Gd9Km46Jn1LQ602KLGagEGlyQFGugBy9KojWrIAMvHZmvcv6ALxhHrl0PmzHG
v9NPcA5yw8CD8I58Tan7xKEP61cGkAMGSZqE4xF3OTdShhYyAtqHrCJd4/jO2vJL
SSRFLWH2vluWfoxWRWfJgSsA+IThQL9+2CqiljI33ZaBhfe2gbU0f22bmymT3o8v
RUGRjQKYw4YzFPj3yf/uT3k3doyymRWwgWdOnABvdLj066eBmFzu4QKQbTeGHapi
NSuYfCRfTDunTANTpqQh0CpA59S0leQRaC7I2fsZ6Q7CZq53p0WcsUre318ptxF7
bTVtPUtDtTmgv1bvxc8gHaSQSnc8sQkXO6S/pJU+rkZ5PrXY8KwXM9Fw+1YEXguP
mk2tgdoCC9ycAACwTk67I65i1kuK/MsR2oUFVBxHSyGQuvXCPZ1V3FSHq2REF2qM
kJsaFDMn+Sc5ll0Eg4j7n6Bw0wrTPqaNWlvAplTw3MMvxyocGbl7lZK0+Gj4Ywke
anG3IMffElMG++Fc3BJVCrqwPmJCZ1F8LKwRpwTTGuEtZig3fJ9TnFrAxBA9GWf/
lYahabjD1YhLuHI/Ho0RQ+wsrTOutjMhRjFz2LYMUuNMNxa23ZOR8i7/JMYUPw1n
SqxR0nJ3fVqZi7FqPjK76ul1r04jU+w6yQuiXR+/tZTj+4dOD21kGQbSdq2eSkyO
lRAF6aCm8UeREAK86wCBkGaTR5MStWiOBhCs4r9Js1wXBWZhS3jzYiX7EDWT6ltd
E8yo9LCB9pQmQc3CXBTqdL7mLIyjLcX9cda5fP9zvxXozxh3GFCH+2gQZBSMBr1P
gAJHpj8cHuk+HanMjRNyGN7+Qr73tASREDXTNMNzcS+RhgTMQtIk+mgkHdYKapHi
4ojT44GouLlO/hk6HBGwIpEcvilokLvVuQfxxWxbMrGGW5CN0LKN33NKBvMwi+9h
f9h4EjjsReoFXG04L8Nk9z7LvzXOi5RzsDbn5OREXhuVjaf6QflwOrCX2FzJtRNN
6lnVyDpttAN+uzFoGO46ByxOzaZ4/J9Mj3q1Mbre2UBwYYRhk2fdcTQLOxmlQMOk
8hTIduR/zUyuakNdvFFrlJZ66S3Ctyaa0CLgKM94oxNodaHB4TIiNf7W/N4vdEvk
XdRMIMQCuqjcDD27Yn1Ibb8p0EHHsLn0QV0LBelNWgmZnzsiJP7VS0M7c4xSDIug
3z/7SzD20yLV2F7jkrwYNq3ljjhvnO7wnfHeoC3uBF4mGjSaNaYXLQU9Mjy/e0yS
bqiYgrX4DjDH6q7pcsid5rvpNSdtVzUXDaW58W5sd98uiYx0hgef8vKiHUu2cPcb
J580iZE5k+g8nl1wBGrQA8Uu1f8qSqTH5bTI1W4WO0WRSZrm8ARPeDOvNl2DPdii
FCu+GGOBky0Z1bDUm8oo6mcdLLYrEIj6ep2COR2sl9lotnlQb51Q9RXDKfs8zZAP
wPOkW/T3eUFiLqKPSue12Nh1TnrWuBh7ZHkIZJjI74ehAg/6jrOtz6mxvi3QkuGi
imM0rzv5eiqVfYC9caJoAgV1j+xy7Tuay0bezMdroXTJLMyNIe0KPoTx3ZJYByly
YPU53ZL3sPfRaSr8a4fRN2FZh624yfsrhvipk38BzjWk0bsWSz2xJuoz6y8aFxpE
wRXW4k3m4eGW9ovMPGLpqwqjaHuF+t/2t4sBUGpvKx3SE0YeJ71rN+4mgEygU/LY
s/CCpOxYFUFo4OOzRUUAO7NDAV4OWxrs+NFNqvM5v0bi+Nmff1/A0oGUdswnWAew
d3RhVu24l7sMYg3Txm7364pg4orTKcjRx1GmBuqpGYCOv99Z4gWRwk8j3rCzJ6ey
isdfOnU/jUd2QPBhJBwOC3cGcV6bdl+XZCC7sWPjx3LAY5isDXYHXDUY+8uMulNr
BI16cdsKEvxsQLVJIHt/DldrMRofU5yt1fxTTtYnqkslYP7SrT4axptJBLEuK7Hq
HLDGhvkt5+cDitX99ES11yVMKaJYkRHbsC3rKoZEVkmxVzeuxtW/Z8W5tW6CwWtg
6pAnwE8JYwwB8wp6ubvFH/oTM2JkkjNGEP84w/LVX2t5sNGuR1oyn4CAcHemwNvq
3ry0w0kEXxQ2wzwsOtyXmpbymxHf0vsXK7//Xzrq2h8OJgCB//nk0aZrk5PhpDGS
5qZ3m/IUk5PO4oMB6CpLqxnAG1Ko23IVF+SUqCqa8EqX6w0ArDe2nURNZGkp1/zD
BY9gIn0tlpNkqL0c4hdBQHN05fPchzPO69Q+s360DiaR6GJCRQwNOEyZaRMWCIwJ
0y6h2uhUgeXVuAFqN9hG2o8QfdS1ElMqoLKTfDwFiuKKgNcCAtwEMJB75F07P+6I
/EsNipq/xjfATyF/xKnnB4pV1FF1h4p8fq3dyaUz3fgP+9d6HMxtDlJ2YC28xBLX
X7M/01slEKN9F+w7igOfHkpMn8boa4TZaIaL5ACuKACb9t0ANJ58vrxu8Ygxcs50
M0d3Gd4dsbvQKJShFOtr1HC+oIYHLK21dQLb4460ltevrjkJLloaeHJxiJSAeob9
Ehg6JZldn3SSTvKcVM9LL/+gMwVOYuRy7Ui+bh1GCx1ILAAJjp9up+CWpUy8G5Hu
Z8T+nx+1qrjIoqR7abnbiWbPsPgzbPcsDIlkpuqTwAeeHoydNER7r8dtdxS7/y7d
vtJSrCI8XQ1U47tlc9Cu20nfiSSyTi+uoZCowtvtuRmQZkHCFF4Pm70AzCJ6ZHJ5
pinxoaEe5vrvcLSjFidE2t9BUXD6iwlrXZDrbvZLqLP70ndDCnfr+QLISzU7HaoU
vui62pFD8c8Jo612pWNr8x/Rw3NA+95VWedTAwo25Mc8SWZebj0WHPZz5rX6avcX
Z6eN4D6F+rTOXKY3zDFwxBJzJRl3rNzJ6Qoy7LJKT65taCQI6ARj2dSxq2beS67y
WwiICo86f8oaYiNcOtntt6afTyFz6i+cpcmR2AiwsYDKtwXtN+dMt330y8LZo0a/
ejhLR1pdvRgofEsL5ChbtK3WXmzKy54/Y03Zs4r/IfZKs76p8gFN0POLFOBXl8xQ
AIlrjaLLbQhDMqUiyB4Ls3Sx1HZFWjGNHjSYh2I1Q08A8q7tCLdwlgpm/UH8p3X9
neDG4AAe3FAzv2lHzdes4JOuYZbu5cHHTeunQ86WTxEX4xJD9kQwho/u4Ofb8bB/
QfmpW9nJGe/MnJvxBg1vCFbjJbVPC6V0J8rSFMpgcu9BCge7DAn6bfovSPSltazY
BCWcZimI5gRzCz4BjhEFUzpzQOB/bmxHJpP3HtsMqPlYSoWF+aAOGf694Uks5Oju
Xh3D6Ay7/xJlGFQ3SJ63CoPiDuoO5y9ZoHx6Hfl2TJQ9/moBXxY/mmO2Yz29Mh9p
8wNYzQdu4uHzJO3MMns/9fMN5ib6bgFjD+jw3TCElb2dRBvO8EB5QnFq65Gt3voA
z3eV8fNEjVSUvUtEMwZcVU4dMYGps0KVR0iPS4D8/TqqTtWEfelEU8o+pZ/bQZ32
F6t/nAargl0dwCvRKYBqPRukIq9BVYvADLmnmBzVkfVsFD0yvlmZiPH9tfQojv/4
vUO8n/W0gzygEm4jC4YK3OL4c7+SR+wVabdbNs9Dn1pmGD84M41WTxKlBpsKeTA0
B5yzg8jkT9eKW9UhmfYCEx5TMYbyF6EjI10mkCGltUUKq2SKOf1x/IQxCaeHiWCb
EEQq0mx4iAL3QS1ELKhPbyKXQYx4dpPouPoVWZIWvHfUNhWpTASnkXCZl4zNuu+S
hVBl1uzmOXIjZavU8LhXYH5IZE8x/20zOBrvfrApdV1kEdPUG8sVJ28MZTpLcsKl
Rm4YO3ZnG3ZPumq1OgcaMOW9impPGWgtxV43hy0ajYsHPFHzvEGhgnpVvPQiyN33
V4iOsalvaYvverxA7tDucH+VDDMhZWWEzfiISjrSXvzyODhhdp/oqrixymiOMp+B
ZxFXjIDWnw9/gdQayD7pFXClmGRi1VIIKO94EkqHS2yFWLZgUqtrLvkiUl5YaKo5
XZMxBpVpAnxYHY1QCRqZ28DxLwqnmOHQCKRru1iLG20K/i1Ho2vSQoXHNSBkMzOd
0tsmqLPD/hLBsRzwZ5ps5eeIXmjoxTzW9SaPX+kfADXVPzbzWpb4Qkp4LfLWYn1E
TuYhtGXyd3b746ggxFJORGSCXQbQmAHGk3bx1U13AMAJW/Tks7xy2nc/AMfapi5W
tEv5M9cxno2MpEvoD2vhGhFyLTqpfXfD2E1XI3qpllHNaWnkp/XC2Ooc4PlUCdS5
JyKX5wG1f8VFA2ZqPpFXSHy2P/rMj5EQ5JZpuf4+VBzj4zdCao9tPPsLputULoxP
jIWU8Z/zdS9fsGrolAQWaDPcAlEkqAPRva8+DEHeFvJ6cJfuzZrXwsfoXyJb/iLd
yiXwKfmDCQKW2mPzcZc7n+yh94c0xWLwM1ZtzdEADf32k6c3XJTok/8F5lLJ0yF/
GjMHN0sM6NQWO/kr7VeGvYff49gLco8F1kKuU/F1eY2697CM096gDpKJW/JaYN6K
jSsrwAc39RqQuR7c7YR7nTgG9HbZzoHA787eDXM1kNFiXshBS7XoNo+cC3rfLowE
9up4SCn+Hp99Z+H4kS9EZkYOQA5L+q15wq8WBDxerIy/UlyWPpMs9ddMwbci8agp
Tx4aNLjGIGooqanzJeRD2M4X1IAjrC7Vgf3453QPqPL5cGEmQT1fGbF7ynQDReLZ
XqlzAUrOGZ2PFd2O1UM0BCVwZV/QXgFNe2ZkPd8YQCupuUSGzUjid4kf4svbGrdt
I2uQk+E8s0OHXhiuS+dYl2A4mmAj41CHG3hltxPLoQ6dji0tOLyBjrdd8OXn6zGw
FlauMxrRP/M0HEgijfXQi9Nlz0yUYCqMyu32R4oO0eUEfrT4lA3izz6d9IIj0plF
9bhSmoBohMg6yyDsXbVX5vi68a4f+X1NDO6hTgsIIrCJg1pGju15g+sB1rFvt6/S
DHp+REpIxWrI8KPRuzvZ/lCKtbShxEPoaUc9zZlUip0M+s+AnzwE9tRMPE1aIQxR
ZApAO2AA98BHzc0/Qu5gA61pN1Td3K2AFsMw68wzfP781kTyKCKgu0u2To0Pl/5s
lMkGPZr7ym7GA5/8GCQ132HwR8dTxAXnzFl/894/KmgcZlcMISzm4l0falMn6Yvh
HAb94uNMoRp8LzeYusb2ZyAQ2c5wSEfIusU1OK1PeyDcqx/Fv9WVYmkYZANHYmyp
boUen6CM7YucxvuJl7FbuObNR/RTtaRzMIYdU0BpKQl95PM3k95HwIMj1qUG0yX+
MGUnFqguiBNbPI1uFlsKh6fHLDKmr4pT7z/7o2GFe/bRMIGzn6QXhDvfV1DClzGe
mcQBGR8i0uWlDdeiXBfOCcl/wpELYeE1JjWpdYrlxmaBgfaRmmEaYj4aL14179VY
TenpzDXxX28hX8vpYmng506lKqLhVAMe9n1YmlWeZ4DLtALtOGcN7ZBxbqk4YVfU
KfB+bVqKCDNld0UyaNK0ij8rD3CJ12qXxS1OhDUTQjsUqXn1oYPKczWnBPlRZ0/g
yD+G4/MmHfk2pQ752EX1FrSgYb4GGtj+oSliOWbUHGdFxkGnZ3bef6t+mQkNtk5v
zvMOqaOJV97JWWdbI3SzWKtafLHF0NyvARA57xfA21Km3CZ0IbcWoSDs+3bFtr7W
FtaRmn7ZrGboQv1N8Gp2OeCzAHumvayA9y2So0SwF8d/LMGiEhd7fLyTIUfy0Yft
DoZwzQIw4ynBtVirAebl7vCwMAqJZfkvvHwy0v+h3mH3WbV4gn/U6K7iUCUUoXII
uw3aExaRjwdM3VOkvRXzsFigV/7DH+fnJKHG9bsf5ubKJkRh74zkGLq9muoccM3B
XLMCbKrDtkDA++Jr+ABk0LAMZpnSYCXPVIhPjv6GIexTKjkOb7UZPuB7J4AGea3/
IV3isswOKKUUW3hUetnUA8MczxY9WFdFOguko1iSr7MWhoGrwSTG16A/3dyimgzW
rdzPOELrgS0uIcOSjlRa6TJBkAmKZYDbypCdhYITYVoS76cf/3wEuPxtSf8h+x3g
tSelWl1aoR0b+vNEc6h+YiITtZnDF2RIm2Aqy7QtMAPPc1nf/QzBp8lq8yvspQNj
roBBcwVr/fFdZS3mxTDkSg6PiKr+amcIVOTkObKnEJsetRQWV+lSJis8t4DOUNQg
il2Apzhd7TexQqZKVE5Aa6iw1WPbdRrNy3HB9J+O/AY=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
G9cULIXhBwd/NEEe2jQYg2Q7fZsTHHmIhbsJ9cKa8p4V9xUhnPow010E/9H7NV1k
dMaRFjwvk4exWb/nQnUh5/UZ1JI3bD+GzuyJoCP5Xr8ZM9Wj5eJwOsVQiOVXF5Pq
BY8W/kJyWGs78c/cqVMg7uxe8nHMT3cu24RS8nQmD9f41JdpspR7nJQ/Cxupl7Y+
8jw7HO1AXAzjyW7Ve5f6S4A3+7q2a1qpGnksEDilcoHfmhEBEP2hQ/2yHpTSQ89I
6MoucVs5F7glHwqGIen+68h5joaZaorxyBxquOsHsgFmKYPh8zIDPpcEXwU5fuW5
I+WTvpFfpOleQb9fFSb1lg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2704 )
`pragma protect data_block
Fb6FCFPeijYdjiZq5Qg9E48M2spzH7s/3gdRZ1DMcNoJ3Eys/++ktY5KqU2RwG2Q
7Y3hvjbvB6emakB3CBZ3Z3CMSbWdj0TUVOqlFCQRfXQLqjIfhJvY5RGnF6m98s+Q
B77TgKD/vBFLTjrxLnvdHB7XNyC3nNus96u34H/xYoXPhwRGyNlsTI3igNiK/eYR
mi/ud0WI3vX5jZsIOXR1d7X3z6l1IjhtXJpx1NtPc8/gBqFkEfFykGBUtJE7F1vg
UkHq53Afw8k4bf7ej6vtQyHgvxfsSewLndjkHia3Dfm82gKYRWqahlDCllUqXTa2
WWqaUskMQ87RabBPGM4l1NytXbkqA/KonnKryGa3vfgqYGSc15mP6GHqDZtxJ4yG
ue77jd6JDqyht70iSfvaaK3zvtuukr6GUtMwGnitzRp70bGtCWxM8Ahr5zTBfSgJ
Pvs3gkqZWwBACm05F+vkyqBUIflRxA4+DsXh4Jm+dHmnYHLDO3LnnJVVufMCcT4m
gU8Y1CDJBb1e6WML/jPgl5OXzxyXE4zszRJWufeGdkWcIKrxAhwBmbqdyB05IF4Z
971i1Nf8loJSi1rj2WUXnBMeGwdNCGnheyQr99f3AqfxO2nyAfOzOg6ai2/TDyyK
u7QOQgzdwhNtLJmPECF/tub6O9ivuSYoYcc+gIl4f04yG++9U3mf28+/5tqOe/l7
E8BUGwI+GaG3VMa6zdjwA2tAD/30SY0guJxdNEnpkdwLqCKtKAPW8awEEnAqIGhv
kfA9IcZFlYQrh5DJ9bz/yoJbQpHMFc7CXxTv6lvXrL1WGS4v8kQhGs9f4iN7JtSr
59vH5x/mmP/KNB9R+f9SjI6NJb+ES0hsR/+SBwsiEGZ78gzBJ6cJbs3wfT0sguuq
dONTizOV3grij0Z3KlV6j1HldBoMeFUQtllLAWl+horgfy5O4THfr0xLXE/hJ6P4
5C61N4ZuH1NqGPRYDz99vTBdEGDoljbEWAnr1mixXYS1YYiqR4SKN8XIF58kuyZ/
vAIuqbzbMeZwWz22RLq6UTjBCrfguC7nHxa7FGAOEqePQevQ9CAcI+6TG+12hv0c
uHbA3esNIPBCPZTJiZF6UTOMw+2CG2k4aK6GWtiWKbFziKSptFWTTYeUztLZ4cxr
T1vyBthf6d/tqaOEHpDA0w9+H1ser6lBQtgNXB2J/b+Zpg9huqmPbrmNmyewxkrf
nJIBsjRDOV00dyvGqZbXIwgWeht6E06lIlLAE2AfaeywMj73aOYUOYvRkYCXrycn
wzdyK3ViSFou/Z7GFv2NfAFfZXulCQwquxXUcBT0xiQA33fTEi0syzJe2749DJuc
5qOM0SlIkxvMb6zQWaJORLiMC6SgabhxaRzHsZPMBl9LAumhXsUXOwnHL4lO9KGN
2hqfY2IgTUKFjgbpsBSBAwJ1nYK/CKtBGE0eKV7+r5hw/AjAw5OSFRlR84DGRjPT
aJWmpdyhNMOrWLvaMVAogqJ4G9OLRWtyIa/JBBsNd2IVL3V89KoTmBwkFN9qBIui
i9wOnq9fs6w09ypsA33bSM3QyixNLJIJYgdZrvRL+J7Tgxi2wKQIOSECuhcb7cid
+EEHBKBkn/UPptcUYOEzv6IuCKHSNp377Y6+R67T69rTHoDnQLSUm+HjV3tsoHlW
clqGM8bLeLnP++3WGpbxI7SmeiyCccTPvKr7/nn0U+R6vAQmmkwJm0HK7aq2BLwV
djAVtmf+drSVZpKAPhaCDFUjo52cYTPnUnd3zdyASeESa+p6ZUH579xoDQUVZeNs
18GwqnBbEs365sdPT2U0C1/FIIsQQKMH1mdpKPHW28ely4hAGhLxl/i4/RZM3fKQ
8BxgrkxMVm3edxk169c712h8oTb8ez/IxyrE7u5Fu1yqfgDvCVtgVD+jmMXgvh2f
dnSuAfA8ofPo1qAMYPhH2TSOvW4rpeBKQuzDFKe1mXrVtha3RAIAD0jntCjN9GBk
u6pXPB/DUc2+QE5lH5xWbIe7HQ6eO5LBmUn0V4wrubPtE5imNwvkyYE0Uu4ITwC9
b3BtkpDqCmjpqxc+38vBmD9cPunV/rBmOWv1GOvMwjRmQAnxsMCT92W9+E+ZZQqY
j72RI7ZCxm+qDWjCCRUrU0wMkpDuZXmjEM2fqoo0JkmK8imKFQzf+4HTYHpt/uJ1
CBA0U/TRRg5Tm6b77xlotJpyv7SjUTeUEgjht2nGjxCZcvb0KNjJ2KjGp/OdTjK9
0DYVrw/MiL6JlyMRp6K0KYYDf5m+cQ99zfvZQDZCJQ082oXXym8jhpDm5uOvqkoa
iPIp83ghRDytcP/2FvcJHJvtmxFhFtsYzkOXvfzZVlafV3P9qFaHuoOaA2W0lsAm
Bmkx2z3Eq7gtrjxNggqlnqFBisrMwFDbuckwf0oV5j5A0L1dJ8O5CEc4GGFQkn/d
/qArvzNT9KQRBT+P44fwhgQRUV/MyUgdXnSoykhU2U+Qi9z0tz5L0yIEw2wlHJcA
54fSGvTqwtTA+hgC8cNMq+iUyrhTEC3B/xS0RcghkXMsysRbi0XlO7GZWog2rwK8
yawxt5SdC+G77kt+MfgcTnESM4qWAyS6gXPc57F9tYWcV+KSx/0UWMtGggMGWysa
/eaB9S69qKqi53PUTgvZtzMjRfLcLOQlX+2Xvrrf0BEFQxPKJth8VB7FlcVYaC2s
hl7RNxMtca6+LFuByduW4kEsoqDe2D69uBXpgV71112a7WVDXhZR01gUh/piVdx6
F3RurGiua3gaXypw+fhW8Ax8tHEoeex5GK3fCqPtk3p3uC6KS2rZ/llzBLAasVuw
ovkStdmad7mj8biCm15GMMbQXpO9lplvO7jZ/SwQmuJRYnKQ6wRCEkL0WmzrYzku
oHXT6DCPTmRLFnE9vvQ10ZLe6x/4fLYX4E+2DpuDVdne+QhTyKrGmXhoGuUoCBNZ
9oJzUX52B5cD/J0eDYgSpF/vh/056GKdQOfQrq01gnwGAuUbeboxTWK6ApJ9J/x4
u25i49EJJ/ZEiaHdHRH6AOBoRfkh3B2P5p2mEH7T6ircxlStFj9+sRtGl9/seYzL
nSBDGnGSdgGslayWqW5xKZ2L59M0cGDmCJ7Kf14nkqNsQ8vaiiWarW+vhbUCtTDA
dJaFAzkXeUw1OFk4zkQu3QacKx0GPRaYVEtG8NcO1vPorFD/hrz2PeAQPfVef1wC
kirjItaMunrciUez/iPZtpv86ZdiUrL2igP4+scZDMhiIAXXcOUgkETd8JGS5ktG
rWKws8dTBfajhBndq6YnmtbwDQQb4rVDk19nJPTGNOcqU0P6JDXIpvm1z10jWunH
to+ARpLxO7YnpI/uszhn+UEUufRF7rU1YphzV1hxXC7KaoqOz9zVFo20tnnWn9OP
iOFUzC0ovUXD3tkDxh+084928llHjgy7nIPvmPQBiT0yTWQpa8ZlIgmnOucNT7yX
4vvKr8c/N1qnSP0oUE6o6q/rUH5+AJ/i2kduZfu7FuqS3qVbh00Acj/QpKZk5jXK
fA0xA5lVGkviV5AxYhbVrSKmCD0grBkHKIFCXq3LoJ9pYmICQpUrlR9FJlGgr3xn
GaLMk59ITNeQLlcxKyBzog==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TMJAtUbbNYSylW9FP4EZkVx/kB+ACapwGoOwgEaLrW5LxahqNUqlB0QDomrRaGaI
2fa6n4wq0K/1e/0+BUlkLvFbIDi7Jra5bqKarMfgFOlbsWDOsp9L4K1LP6FrC+dC
iZSM/mXjUfVRT72A8XHX7mFT5Wu2lEydiRh04fXojMA4fJY5hJ0jGNJfm2PtATl9
YmE0vq0UdGrKhi/DQNL5CxuFRuKeYt0v0DQoCIv0GmZSItHmLtrl+jhTRewmZ7A+
9Yuh102wVl6l7YbzFXF7NdNcIqjv+qbfpJ+ByA2B3nnhi9ByIvfCkhsASiSIXJXk
+MJmG+YsLSJRUKHp1xJg3g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8048 )
`pragma protect data_block
MpgonWG3kac0AdH4zKe+dWc+OxJV9EqnRko2enqr/gNdRxVRPaD/RC+wEmOBuLQ+
o39tR6O+xFjB3pxNXSNWE02iwRVj6ZI3pq2/yHYJ2TMdviDeQEvFv9TZb1tnoGQX
Cujd1Cf+MjlAgFG+l/RHPXQ+RdmVn7CNxI6gXx8r5IELvzE8xWWg0hp/GBEPssbR
YTO3BbAGtglCKta5zxcXzoQGpDRYG7gnOTI8rkpNA1H+cSkNX4/ccWsMYUnRWbsR
HumiRw+KsBwg8apEzr8XLeDjktV0e4A/LVH3VDiGgISE+yjx7kIugZMlTjQGE6w+
CQTnCB2krp2e7CXHg3jAGU1oZZvxy3yvzH3p/g+xZrhfIocmxoz1Yg0pYwWXHrhv
UqiBSerdn5Uao29GR4tNjqG5rnpTfwq0qI6UFjx1yaw7UY0oSCgfkTjyeDQ6BCUJ
/RKB6RBtrMbbZPZrP/QRWPqMTHKa8d8gSoReXDUApTAi5pc2AeDbEhmcF8LWcsCz
5goNoS4lYjrSYYU4C2CrPotkIJCzoCVqTcqmAAJFlHGHLuIiA2JRxyHfgPSHEtAM
kij99q7gl6ehAA7BOQAK/Hed2QnqkxHWXz7qCCFWUU1bJ4jpoZ0OQgRAeiAgiJEb
yw31EyrlaCXSrfGzzjZTXInXttvQTs7BUxZ5RFuFm+E+ntsJV38ZuRP5+72v1API
kEoViTVg7s2WA9+1zLV1xVXSftBD2n7jHzfS32B6qFR6842BvDxoWT/EJq/y63iM
RD54RPoSBmtFbyknQF29lep16/xaw36EbkvMPZJ+p2UvodWQ96vAT4rRSGKf4OHG
v7pFTPKBD1zD3ZfzK2ggmDjgPK6MvrepFJOPhnNfZP4ZkUwRRlnzCn3EzDLHo1EA
FCbbzTOL3ljHs6NxF4deyWRM5YxGrns6a4ifs97T+P79v+1S9dSJi4iZKvv35y2k
Y4UXmOXGwCFEsCEWCe7RCgSZe5dpD3w0E1QcFk4mXta0yYFAIpvIngQXsMYxsOMS
aPfjlVbfHPaTIuFbrLG16lTzuHcPXNiLHhhFmEfduvwYJ0l5rNDb2WsLXDsq58qq
A+UOmc3s5lMPlYoxD+bMWQG8vCi65Ik4wfivyxd8PUyZ8XF2gwZa8A3iVgncuvJR
BVvDiU1nVAUUpZl6WmvDUTijIXr25wowZCAGIbHDFyYtovGOPv+6Qbnr4wLi9tfY
0LxRqtpjm9Pdb4xpNte4GtDESUM3+7fEjT8sMYJnnzRNjLKOWZAuXUC+H+XmY4Ue
0j9FCeeGZzT1H+LJCLu++WPq1mEfdYuogsmbJmWqCtZ/q4L963T4J7Xo4BBhT8Bx
q7lVLQCYmhF5fwVbJiHpVr8990H14INtfjn+R4ED1Hb+9JjGJt2UYV8MfXIhNK0C
3/bI4ukkqXWrZUu9osxZA1MzG1sr6h2Q02dZIvcfIeaMz+Dj486UJhWgEYUoP9Dj
Um7bGw9V1bKmuJ0KnzOquSn5v9rYFCJScoyX05pKxJGh66OX96Kr8q6A4b3YuhBO
fsR6CJaZ8/GDYeUwNiqSykgFemeWtbfo0kU0pHg+Fi0kHJWaKx75hvsrSm+Tsaoh
jrskeaVteID6xS2uzL2hMqEehRc1ILxcSU/2BB/snnq+0QnMUpM7Hw2jlK8bQmvC
YvfDYdSU6O8op2Nb0rS9DFLVu+kjK8LOemBoVY2YfMiPcBG1+nB4XqaYuZCDAgtj
E9M6TQsMPzN/iG8FgIj6GVApB2wjthqCJLRfx5kHMPSP2cfcdwLtW3D4pI22G2pQ
z/TQV1c4KaJCKVkc4Xdfwqh2P2g43ghxWSto7LvMW+a6/dFEbAQ8a9PX06mCx5pa
OFmBIVY2aBqzNfbSkQheOq61F7ops8XJW5MijImKxaDhqR+75lu3IRk5MHX9IoKi
RrU46gIv3daJrkaLptp+MMBLE4II9tIJ1r9TlMWt42R1O+zfgFPLfR5/CvY6nmQq
q0XkMhyWN6OrYq0D7KHQZkdj5KAPQP5Gnks/5QNFBLJ5WsV+q4pQnkaJpuMaH9KN
kRg7hjdi/T5xaYUs01KHu4+/+XXmlGZoMB0CuvllKrEBG1pYt02xPKGYrTbpulNT
oaq7nr6rGE/1n82jLQCCqpvtDLl6jqc4nFw+yyj46bzuxylPk8i5bCxuZDvD47bb
Y2XtLHpO3CovNC6+QtQ7iWKHCve4UZw3FmTmfOOFvV6acJY0ZhkWDn8zSPFiG5nL
3L1SXZ4pBF5I7apRTaMxn9feKYBHADD9wYvyvWdW8QXQYsgKnMHDNfuqNrjhAvKe
B7XVGysziGp7NcbWZDCE4MUjGeYiWv1smUrmBvp/0tVIgSDxa/2/H/QkDyqAsMdW
Sos2jx79p9u0661HUAc7QRMQ3Le4HI+X+ruzMTZdGd1yYAR3LtWIdI2a2okX5b+q
EEpaBK0GYlv+EIxh8W8aPiOemkESi64FB4nemKYrg+dLQDzCrnPl2ESWDwcR2wHG
9UZhKaD5p6KqdFpAJe4y7oQUKC4IN5oBwy4vf/Tv2P3Gn+pR1TVX2mPalZc7lgJl
Jc18U44c6zxE7wjrXamcUNY3zrmfblIz8WAieWN/tomNOhvnr8I439apHCQ2Po0G
RmNdsiqoMVhYLxQNDpNA9aG70M5NWoW3lgXhIKaBrNhKfqrJ+sRdzI2ah9S5xl+e
34VDVpQGa04CEkj17lGml3NdBIJe5+NUvsWIPJ71MaJxBjGf6dPXQBU/xMvNOFge
7tCJJ8rR9ydul/2+qiHg3hOYvbHOjjP/O2nnMlO9YM06OA2nfkXPlnvLWR4Qm/yv
5eBlKN88lqti5NK/G4l2OW1fTz5fwNRHMZ1Dd8sVqTtEddbT0ycBKYWN+x2pBwib
QDI51rdzqr5sIDBx4qI+t+4L5FO80pFW5qR/sOCPQrErO5QEMqI7R6f0FGkeX1B5
QklBKJLEy3ZReW6Ax0ii5bTZNpdTU1T6FEHuykh+HuMATTXOh2RpPJtHRFNAQk/K
ZdOORn2DBrkKdAT0+yXnAuRCQIbVe7VCaM/jsshGj/ZR1O60GBnxi50pnb/QB6Bm
IAyHyyaTRG30JugFUuxcLzZjHR+U++WjQ+FbzIPnuKyq9bqEfVa4xflC9WLbFZBT
f/cKQKP+iZiTcXOjHhM2FGOQb5Ll3oISPBiHmV2bbMQJewqvGKi1eboNpbQweqJ6
MCR5JrqdOs7LJyB0MkhARWjgbrgbqegHCiOiNvkzcO3WaJ8FmiJaJVAybC34weF5
vVNGe6TPQZSZk+iPAlIMmAdMtbTQ6jZtEdE4KheE8yPMoidJZrSjXf+GmNb7NPiz
OgTr8FRoqHt6I26KiWWA+JS9i3yd4QTdeFbr8XFKBCMaNCOojm/iChcrSjA2uaKR
AVEjQXSG3t/YpinKY/ruSwNCalXdQWkF9gCr/QEumUeX+ymrf3TOOZ873VYuwBiJ
jIkdnbZHsMrwiUowp8u5KJLbPYFQYaPhVO2+PzTyuRQKdNFCh5lQ3IHroHq8N6O+
TXLPG4vzArQCiqMAM8VTEvz2JHbb4wE3ouhXaOQet5CMtTwE9Ebt51QGThgd2KUU
UDbWGuYRMp2O2yjQo0exJ1o/KDR3TEgy5a77c32PKbMP3xV8ZR+ACSTjJGXI3Nt5
xPxqTJOoyFrUO6YhCllqrejPjh6Ql5xUEXjIUrRA3i9RvMCWQfWtyhwV8exdNYsJ
ztXIIJvUhJ9OXT/JQbfRRO3HJ6A/rYV+enz5RVl0fo8eP11rcd4OJXbQgBWyxvIi
tdCj0NWza3h+IlSFcEzUQIRx/LJ3ZTmQg2yWKKzGUKi5ACPrA20TWLTR+/kX0+1/
DwPTXPyWkWu8BI/dfNA3vKIPcI+Cv0qEsHGcJAbypK57DSb9HBa7+fisA+G76FBH
9CpbvqlCohVNkvsSvDo5g2kOI1lC+uccB+cl9V1to6eWw5IorHNjs5B9zfhM8Qh6
NV+JR/1M6V4TBEI56+TY28udd7ib3ONbR7qPNUvtuoxgoDUCAQ3IqSC8zyEaadyK
JT/Q76EG+njX+t44vctSdkYHN56DwuyNFUIjhWYfighFUpRAvTvOTmmDxgxxQGVc
gHK9vspZJSjsSBET8qqTPk1W8jrFCXx5+XGmADOTmmXLFC4f+Fh+Q6ul5TCTqQUt
p7NMGW1Mxu+yduutfbZw9AOXssR3qODUD6cEvd3CUxixpvtqPNlHl4A/XrMwoR+T
TSy2zcnRvufqSY9Ij9BUTTSd9Xd61MrdyCzpz1JBtf9IUkBlt697lVbWubQhncWx
6k1qAAgA3K9XhO+JXfDzs3XiNtouVwZgLHU3FJNjeXDC6Kh/97N8lE5tHiFzDj1O
zG8r6vpBpRzAshNDbEDk9iv9cJf/HzD1KRlP06TKjtHSURCJQWPkPzAXQSff8jv+
AkLMn+FeMHosXpyvfBG9ZWpEZ659vleA31ZSQ/RR5CD5hHx/PwxTJk2+LiWCBBc/
XDo/WtKbvCR3qNfkjECAEMFHGswmEG1AuEp7IiRb7BlL/o9T+j50sGFg4J27zWtK
chnUtaioidYALbOecr45teMAjR67WEAuHQbOjUTW39uVctS9wrlX/vaTe/Tqxq1J
Vn6F77y4iKMOH85a+6UUi+yoKNZkraJ3l2qevlKAMxFGyhPQaHdzPEILeU3JOLSQ
z/dbjNbzSzDiPAEMZuCVxMMhc21I0H7d7UYZHeyPoa9E515LW0fu0j8eBnLobxZy
u8prJqeoOC9f6yXPZsL7/Wii3e/I8IqNYdI97G8Ro9W5928wTGWivPeA/RqIHwE7
jCTkFt5sdm+MKwLZAquO/yWckLuhgnnH0YqCtARhRgVr3lZWjLth5vLchIWtWris
GVOdG50Bu/Ff9vJqKkLL1eOB63YHiVv6h8qHJOdMMqhNfj4p6HV1Ht0HrqZc2HOu
r5kNhjpMjoyg9slDhx75R9OQACMcgSNMJDrswqDjvRX/2EIeZlYiJcyY8UGZzl1s
weR7Vi5qB/buB0y7UCcuJp2ssqbbLMkBQ3LGiSXyV+4mX09+cBntZEe/78XXi0aC
uCKF9WUE/9myPLx38Ov94zIds/TvpsLAbUDNV8SstNj+0p3ojhsPfLsOK1+PYfVJ
TEtPM2oRSXnIw2zBtOTpIC6U28cWuE0XcEHCyd751biAk7Yd1uWPBu4x2AeFsgAM
hzR/u0EjsSrPEu+sUXKVhEQi3sSkob8hOK6H+eGmcuIIDTTRjGz4vu/3vutW3VAB
Sf/CKTqNJ9stIPDxwCkulNjPiqgmVhl9vQKPmytKT70do5az4VBLJQrMut0H0RxY
N9+ZwKQ47vZve1EGxKC9BCuwEwAA6WGJZ19wJeWLYzM5zZqnn+bZeRFPEbs7BQzX
VKkPyeM2ouoqad0WDatOsjedfgYntol0ysV5Vdj+SWyfpfmCtnNi8mqt1ivA3fpZ
CWcpSVtry5PbFqC4FyW9bc1YKzVLXQeKCslof6sYG3vxI9MK5b0K20OPDO6vn1qy
O6ziMHvd41eU2OVwPiaJO2QR6cR0Hiu5aCPh17DjacGvQpRFlRnd40/RjSyQU8tj
iAByzMls5L30t7TOfWL8kIqum0RYTEl9t4/f/1PWMX3RFIHApOte2cKmxyfv3App
7lPIQ80/LuJRvQ6PDyyTu6Dd4hPiLF0TpflKQNvHIX2BhxxFdk4m9NHxN/Fz3pbg
ZeDCYjXNkckIJrt//5z3uH0YS1Vzq979GZK/JzRRLvLomt3yWa0M0DCxjSCh6tWe
aU7z2rKT/2bcue6bAzvYBXFBxubRrP0tc4VI78HXM1ZGG2VHGHFXryAcTahorLRT
11uOF49dPHEm7HLEzSGc3D3Km0/n+CXWP4tSaem/Buv/jc9/0BDRzC9zvw67G5H3
C0IdctgxSJg/rPPbmTqtQ6ii1sQaR/08lX153syRdpJXt0dYiyx0HgggnpihpSTu
mR75mA7OLwk02r7iAQdyPX9a497Eo9xjmsVSrBPOboAqaLARW2gjvkIpnW9rsTYh
b5t/H6R+GUrnCQMWVKIAkGN2CZEyFjFf86Nx1TmrSHUIMzqZYEs5ez1lLJu4R4dC
HbCIuQ5x3N7ybARUxcaqX0DDQj4QPdOvu1yqu++kRJx++vYG0LpQLMyhRvZalMB4
M55/92o4/P0lfImHrlFf44S5eZUpI6bXoJFp/Fg320hFR3Hm3KdL811MP1v9kTw1
V+Qn1WTnW+N+WIW4CbMHpayEP00M+QaUBSJrWTUAh4xFHAH+X2FN9SRFz5+tng34
vJKKJEXDWvcemmUT2VNP8cpeFNuyKxOVlJ+HhJOBxCqCzWNAgcKlYvkMlxsbtVl7
7BLhqswEPnUtJW0NHITxsWpxwXXerV+lNY2oEpfKipGVQ3e1woaGrOqRzdaeh3TS
R1VTAEC+grHMj+uounJDEeL3edHxYsf1ujzORu1D4SuOnCdA1iofCFlqrZr5HUfs
45gQACq3ch4qgKFvj9eSG0ReAergrhT9iZU89yh8LV65Xj0CjVkl7843/hH6uCm4
ifru5ZjQ06MLykuKl4SfQVSjNXi/XSYC4Bc0IpHaIOpb0JPlJyjlPOa8bVSGO8ec
ZoQl8qzRRyLMeEHVyS8UImxL4duVsd8ivPacEE0lbjt45QlA2bR6QItMrzMpTRra
pQNW84/+hACR7i4ugASXaYQ1v/ufdUYFTmSUCLnYWA/crAlldQNaa2NwwnWXsvzV
eYUFSnqI70fwMYhGMhBctHDLQuGEb0YQaakdBbvfntB6AIvnPzKVDzeuipLGI10x
GV6bwFl4+gTgx3IWGVXFWLXqFyMpCcMVKbGmDmQJknkUS1wFBAO1IbRViHSfaLTW
nsY8bc6Ej4r4Ldkj8FXoUcTcUZrAYPx2Y81xbNct/unBszL1nlW74bF4ZiveHLD7
VaXfYydY3LyQxF1aJFhv04NCRP9knQBswuV0Hi4/TNtX3Mj5II7L3vxeuIKn6Nmd
WF5xoB1m56Jz9HPqCKZCYf4iNLhmk9Yl/VQxZyTHdo2W9h0aU9Kl5G9k2gf7CpgW
WcMPm8aF2aGqLJJKiFaO0pJ/D1QriyPIwC4JeQLiCo0rL6+MLjsuD6qeL8ujqRBW
KeZuAy9cnoW/P3H69I4q91kj2B3aqsiYpWmuOz9d5VQA/TbmMzN/jN/WywFr9F0+
eWoWwJWxntormfqHvTt7Qdc8AoVXnK8wwVP5qCgkEJZz8Bb41iTMKbmUlubH8EHO
BX9E3QWtVK7plTvBu89UYtFKz8Z2gmexsJgdSxbG7/dUTFULHWnyi8C0ayHc7jSf
MSGSv2AD1k5qxEtjsBUAKTP17/YufwVSkhmFPRATKyZ9VuPXnoWgK6XNyWEXQZah
A97Ko/hNWTkdyDzamJ2T8U3Hfftv8YhIzju7IpVaDFY9cmr9HLWEoUts4o/p4VgM
nGeGciP5UnxBM9DfqhfECTSvqB5BWQmEBy2wJnGhgKZaILWP5Sf3hNfySfyHT1I4
CGAywxHbTXg0r4jS8kAtXWkblalCcW9Y2DaTOgWeyOoyRxoJLe1/y+xtavvBaNGh
Dt/g2RaqPAuV5RmJcmAwk5AIW1Qhz6bwmWUY5JHDN+KlYGfAflPjgCygwFWBrQ3F
/5mdJ53IkHJa7xomqSFZHiYfbR4UPl0oE5eL+EflXMFrDV+LfbPFDmtde9nqTRMs
FeHzoQid8X4lWXgXfbt9ThAp0W14aLcdMfx+Dr1JiEGzEIFouQnS+BYAid984XXq
n3nxuo/t7ZT6ZFEHMdJvc8v5GDA/aQh3P7LhZW3WDOEDoVzdt4O45DECAPXN5D9l
Cvji0FAJTcm4w/eTnoPyD0DSXXHA3buES2+AtTxMYxM3g6CSwZ+Rke6uYmwQ5k+D
9nYQHMzQvLdGMBsahdbngVuaLCz5QykU/gTplfmc4AKVtrw4bwZsu+x4L7gJ2ANE
U0Jw7BtdailewYL9CkwHbSyktkRMdn2Nabc5C5SR/1/+oYzhavol9myOQUSoYHuw
/8okHKxm4GQEYHSIein15+UJcIBn0VYo8f3+TvflFzFwgKyjolyf5a9C4+7gkEGg
aH3V6JlbI2KnvTe5h5ViA5JLd9IyLUwAP9YO+vr5pqfw/3QEOAwRKfB5klC2ZxbF
Xlvc8JMLDMPcr+pgP6PR45lvVPrCc0O8GwKbdjw2ehvRDZBmNmtEIO8NXosyS2XP
9p67B0ZZ4y2YZecjkkNnOdJSfz/VrUDUkcokZO/dOGMqXqRPrftZhQmgtbQkQ1Wz
puqqa7B2yAlkPtX0bpVvE0Y9DF6kpLhxrgOKryDgrF2+nJq9t5aj85nMXJKrkXqe
9CIAvwMAnyA7T1+WHf2XvnQtFOvoZesWDJDl7pR5JLh7tagcskdWGu58+8xASPSN
lAlp+8ilzMfFnfYPqeBFnYUNfDzWzuG6BJ00t4V6BJjyvpUkMcy8G6FpZDqpFA61
pkzu4Dki7dE/HkPUw6MnB9toZgfOhvert9IdOhxIl1Ue3gV95pR274JUjHlFlTW0
BUTMfPU97HgQU1SFWld19BYnXuBfap45cnaMJGSZK+iUNLOMO7rCoD1WgMU34yPq
bzLUezK9Ea+xTl3yoblh+ftPe9cFTFcFZR7To8ou2LO1cmkctnKrHdsL+S9pSPAo
EH5bMCwFbjSs+ukfjH+xQAvicgKi/Z/U5KdstW2UenyRxiilNXMQq1zkuay0A1RO
/9px1rvfWdqSFx06737EuxzOzkqcw6w3UhYdGshEdS7YMg/ikZNked56e9bgU3CK
VGeha0Pdbw+B3dmvVAoryWGPCo5YgaxfNKzOnW1la4tUfKzaznn7OTR7CWvpby5Y
1Js2w0567HxP9T1bB6NE66bDb3RjTBevpi4lO7yMADkXLfmacvRZg3v5fkMF7San
KEVimdw6dm7CvjhAWAIHcbnYME2ZRDe4MwapwIguzsT7+xx3qXp2eIWVj4brWVp4
3fFUn4k/Mns78XAHE8V35aO/ugBiHcqrR3NCXyum11c9YbkshZWRP5V4A2Yg2ifQ
ppwuP5PY06FgmN3HtuWOBlmDapqFZUmWSK6ifqHDt4HUYN9MOlPM8FGYZ072Trxy
kSf+bvHtTHf5GRs2s0jSfKvED0/+ZmftBvcCjqMj9VdqT2qbxDUzBClcD8y8w0Jc
lmx02aRoaiiW2yaMFu2DLyw1LPhv7n+drJbiB8kk2yvbZvYgT03D0SSOfRWw7JZO
qtRbmqUymWL+tGOK/wziyaHgspGp6ptx9uk92m3x0sP15o/pyy0m5w//bLKSDllS
UdoN+l42k/N0bkPilcdwHdYl2ouSXprqltoVMxKSX1TC1JcBl05XjjuvRspRxmhl
/Nh4DtNfso5dY3DQgxDvdAYTwpGezcBEQUPfVjMpP8SLdkwHwcVyq3PXa6bnNKMC
yuyYDVKRWul3AurhM2vz1X6d+ZGOL96Yd/YNk8ROLVJjgniDPAWOJGMIEENwX5Ef
8yM6DNWafEdSC40VPXFKQlfrKefGw1EbKsKmI8v4KaoNYU8QXVJxjs5g/F5fFAgY
XOC07JWNVZCGwkm+0EzX0pKShqmiVk4+r1lqep77bzd2sAFcObzwM0RXCusKSQe3
HvsxeQAXbWaVn1XTGu6Ns6+leDEasncHBQVb40mtlJ2rEnBJChkc7SvmOSnGQhKk
OsGb0UQ0xJJTAbrljwpaTw24QVkpdDe19xk3jvux0MkxKG4QF+QEO6Jo816JpFtJ
SRUoE4jUo9Qs6PPziDNHvw5wDybfYP3nv3zivft10JUnXVWgcxLNtgheBHQHj2fp
Cizrkij6ihSRuptkuQVNiNIrwLqJtYrIrLu1OsqqiNjdPsOM7Fn+GqbNJcdF0wCe
2O4gtIfbFDr2mhnmpOIc43y1iU5XklZH8QVPaVdjqbaa9K2mDIxRsaddhWkrHy6i
VCDn2k1PkazGdHN+308UHSVzbf+eD3vFmsLGXXbrXq4+6p0sdVkW2p6GjmaJFQTd
XL3aD+Q0pW3GHrqKGCjASWtRZHbqr7K1NsmqUe6o22NKbBq89TpE4DjmKUQA30mz
7HhUDdYJ2nTij0ReUCaulqU49sLAlauRbGteIyoAvlkrZ7c1QhBUW7I2tglfUtYK
e6KaDGErHjz+rBuVSh6sgzyxcQYAMAey2yhu2LI+UcqcECMCm46d2EbvpvsxoPC8
kxDaFQvNsEyW5dTXn/O/iWfc0J9uMJn7pCugilPTtQmZpFZRYZkEK6cOZL7QTyiu
JgkT66lkAFijR4e20X9I/eCsI8HTnFA0YWPigS0D8gFCGd/NFqIjtnRJ7QWv2/gz
vSnuHvDOp/oJs+s57n3z5fTUmz4qaJIv9PqpvX4tq3P5bGKG2pK37KYz+sETJ5cg
SgzL/1oJiSTwewo9tg14XWCfRFoMf9TsYEec/2kIGgi0clvV8IYe0oIqOVad4cAL
Y9j7VWf7ssCwCd2NOLuNa3Yt//zuayOkphUgW7XJdERmzLYrK+gkfD2KIBFGhGOL
n0kJiphLJowMxTegVJRG9j1+vPt6AhB015EOkwMnn9HsbhIJK5Q7HVg6dIC7HR8y
kjz0Iq+XMcY66UusJ8Wz7JnsZWFeyqpxlsC1Dydp8nAMnBcytrspPJkWqm9W0Saj
c0jIjBeX/+zMWfJ6p2v8dF1iV960riSqEzEIAPCROTqTGkPZFRsJcACoPCXYUs4E
c7V+4JaJRxSRJqmXhupwwcgrBjX3iQDddX/4nSHKCPg=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WcAb7SKX60eu8UvqB5OMGhJLDE1EeK5YiJ8kIKGtSBO2uH+URJvhKqbeRf3esm4i
BLDZ+xsyTmofMPq4vMx5ZLK6ecBPrXdwB3dnFUvq5XPOe88CkiAvS0T+dlrr/mYj
rA7j2BS0hel9Y4HCkxVQMueBewB0z/DmGQ2zUJeIGf920OlXIKMfpUA0tsL1ktr8
fAnIsrSIwe0MTJMbygormADcREXpsFozD7NkXg9OgIidFfRUufAtRmxs+4/gv0IT
iH3bwBFIoiRnYPF8oEELR3K5OR6Whi2RONN695SXRidfllczHnMU0J+ilyzMqAhH
A0YeKaExf/1ihQZLMcNUdA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5360 )
`pragma protect data_block
IXeGFQl5kCzEDiwJBFq7p/ORvXtZJ+GCaETzvY7iAL7MTSFWfzbg8Fcfh5Wqwjjk
FCoqykPBYptvMDpKavkyeBMF2UcW9vOpTLr4llOM0XWx9+v0pDIRuszJJ5N+DkPA
OZdhNl/4xbrrAcbuQSLP+G0sq1YgxwndsQnKHxRMo2iVce7Tmy1+Hxr+zIgs+Gmh
8UhSqWcwL20dTIi3m7QMgnsIx7xrCT5Rn+q8ob4wrJu+GXLDViWKJwg8L7364E1U
4DEyKIFlbhuoTPajQ5tliYCEHn0ZvNawuzJMtc87OswwKlgqW0vPUyPF+AmnBKOv
yKd3VbtfPSdakg/kpf2FSifIkYWOMR2VRACOay92L7spKKvKU3JoAvb7Qgwm9KNE
Zyjy9pvtYD2WIkkmW7zTWfpdpVG+MXNbhmGjEbGHOzmBUf/m2Rg3KSiIl04ndYXu
WxfWjPGkkjIlvqB7DN3VRZ3xXPg4SmImb7Kwt9wIJ3alzcuKb2TN3wHO0tU5rJ/U
mJrp05ovjp2QrhWa2bJs3FsqsbXGovd9BnmiSo2XVHS9g9uJ2wEAa8JWeJWtlQrN
xCP6lYUrvB3jREUQTiP1h7AIg/FRj2looVC0YLHDuIMn/YYCwM1BtSt69PDJPjIH
w4stskjCqRu40mFzJEDjdbLctObKLGV5vzjtXbznUU3iwikN/L3JaAr5ga/Es2Sn
NhJkGcNDnAP5O3U/jJ+8nSYJxRFxbaJYWsq9WL4tfbOmiRc044YYTBCQ7xWnMWR6
nTODwnXiquqjKJwndwqCqR8Fmvvx0mCu39I4seb4vJHJhaHo/DK3HuxT6wwBQCDS
WykUIX4RlCmEUmGGIlELMyMw+p7LPUTgtuAN1ihjtnitJs0GG2TETqWHmL0osI7t
euzjMiL05aXragP12Dq4w0NzvEcI7sBUbGTKJyc1GXRRCUCC5A2diXsLOyxTqiFX
qsJqBV6MDdiVrv6Sz1wx5UKHCQnMTvR/Rf8ByKxs36MZbQph/eUzWLcombwJrTlI
Ioy7oY6tSP+F4/zeKrGjP1c/R4VuUcaGuSc3tVrzvpZs61vuPXw8mJX0YPlGZ2xx
dv+Qay27/btulU6mud6Xp/xYZJxSU/gP2N+1G8c3t5mbRw2i/l6+jdkToT4bd64W
GtG6UOPXmEeBrn+YAzr8VZrEWy2S0ZJwRb4izKd1paV9wNlyrESZTQEiiJz0xz6U
ZyDiturHh/Wm9lG2fF74GmlpcSiQXzjQx5ENtMK93z9bSNRfu1YZTd/p+Bom6Sm4
9TMrVtZ0LFUvjXels4iFMB00QON3UgkaiAz8GqA/iMv8zak4gX2IMkAK+7xLlqjB
SC0Hyiebq38FgFPgxtoKXJuFA9Izo1WpNK4z2rLUY5pVXdtaXzOzMm7B5EWLebQ/
0IU3Kvw1p79/5v5LDRIdKSVmJzgpzz8HbNveHsyB3MHNEMI8p1ZPclvKEDZMzxKl
HhNLLZUYoPy+Uo8tivRdaqHf15anvyNLR9gLDvhDfuPThYb5sDVHPTr1KSNoViqS
eykNhbS2c3+1OjL2JO4EFgCZQ1lecWlMvKw9SBXwjMP0niwQqcHbRf+L2PI11pfU
/cfV2/p+YxJd0QizEnyl6h9MbLvqwc7hj6UQMxXHqbHqPDT0VN03Aq0MzDo1uNcF
Y/qzN7swfrQxorNfVGVpEpjCzXtzzTGO7Zq2OPzSuleuhKySxITWtHCbl6soPGHI
1rGVjjwkA12GwExbQQ+2xf8yzbvScAhlV5kIIzUYTqfMsk1u7psx6xNkJarGNlzI
/45jQFpBsmM3Dby5rK8lR7S7ZQ5DKaDkXngT150QSHY8WlAWvn0PB+bhXPco0Ptw
9dXsLLosWcT715virojwhwTXA5GNEIxeRlNmF6kGJbqjJf488NEXD7HaruZl6Vot
GGNKZFXWvxiNfprPfs1R9ctqPlec1DwKHb81MLbvEADtRkHJz+ly3hzFhfk8ZmBj
EZGzVJnmdjljSU+zc8p8FzNG0SLT8AT/olh3S0/g1ETXat1uDxofjlbZ13Z2ML1S
+CryNOm+SC0vzjr5gUI/MOM1lMsCjhrtqtVMI8CUY68UH4ptiYo4vXat1R4N6MG/
uBojU3bchP2j+4mAJDmcmeV52HdiEzJK5yqu1T4iYkSj6tf9ZzReDA4+oQi8gMgu
H4P1VLytfK1iEJOGZLFs+0YOqXcPGhJY/evgezjtw/LQhTwVfQ3eJW1K0FoN9ges
wM60ny0PQQ9e9Sk4qlsrIjkBMzR3LC1Z38oMq+7r3dETbZmIUqRS5Hhc47b5zpYn
H4n05zS48XgScXZinxmwQ+MRYSyY0xkP2aNhHlWYSbEDVHxWLN6koHXGQtrtg+oO
FO3ITMRm0oS7hnLzTEpJSk77AGvcm0+mQMk3Lc1lw0Soev9REaE05LWofgtaUFnd
SVhh2UQ9oyMqG+SVL8TeLXOoxBuVRY8bCetn8IN07Y7tWJq+MnST66DjZ8UMb+6J
CA0y/breb8NUP4yJ9963av0fk7LIRSFtQ7Ga0j4kZ/aLwPjEoq/TZTRzqCcApOm9
4p37aUeieoFff/mncU9yEfZllEHKpErGODN6MlYUBfEmTQ1PaFKarf824rpg1nIM
STyseqL29qQz6BTl73kp23GKqt1HIyjfjAsvyBwgBtYWrbxxFC7Axtd4Oqr3I2ZH
GXhEyt0YFj8ne4YsPylVuZ/CjYomCqhc4vXIwnqQt8e1S0goGbB5feZPNQTTaC2h
DP0R1yclFTAY0OpfR5OutGgMAZYjqAeBmOlT5AXYzp0ifVxbeMKBcZodn8AUfCR4
Wkm0HHEUTNyp7XbD183bPlLzsz+UCQTsAgUwTgL0Vvg1fbHMAGidtTtXYZhHAHdX
/krKZmYFJN3/4YYyXVuy1xZvzwdbBzLUrHX9Hl91glvUYXBPkdJiliV060eSJ2wU
AbITJU05RNWKa6b+s7XqdzFtbSSc3UQ4X/6qVWboo8lfcv9ynWQVd2FOv3CeOtYJ
gYZA+09OxCgGQwlHdMVO3JUNO6ClCLgmiM7LnP7BwPGRVti10HTnocpkf1lANJPf
fdeg3L5HP8sdlmSgvFRGbsnOKlFtmw2rQl0GWjDFTX+gY51t+HkC3cRTJhriQkmt
b/1ObepIUtZ7cK71hgCD+38hm/c1L/qB0DRcdFzyMgNth8+5zxfxUTi4W3Mb9Fx4
6+Mn+YAFI+MMZWLufPGbDSGlwNpRZO4smFt9arqoEsLRvcGqtFi6+AWcworODw7B
fuVzKoT6yQCuZ36rT7li8jhWIUSgeFwbLsDzBj7Z7Q4kEGGPNsLer4RA55QIVdYe
AGoXWHyAF5x+8nilgKHF1ymRwIiR4CTMvAEtYaijhlI37xqIn4UCoaqL2QGKfznP
J/12UlWZN1n+h3CpO7bVSWjPCvjS3nrZRxwkAp4JMjwm84fciKy+gwnlJdNKRgFt
69qt/UCgSr/LCHlcyZAO91dWv6AdkH+m8xU+bkoFVvYs0V4/ebt6L0Jv7jWs5Kx2
NqgkfwJgL9ocqXJ3BNAkGEcLvGk6iLoyr+ox8bLb519pJM5FNqmrrQvzSEkSKw6V
s0hBD/dD7DuwdGNDPDrxjfEPmkYxxK+ndGTnzivDyHskAU1iRm+0UjBxNW0EYmL/
e0sJTZ4kg5bucyOlTo1u8sxhMxosaZ3cqHevD7XhrdrRuSEjMpSJHfV62cdxVRJj
z7kqLCU6n87p5Zz/0InZnzBanE0pQa6irm7nYMOlK1kbkFD2n1E6SsjpPlUn+rS9
g6j3o8OPjLdlOAmKrgqMKUxHh4yEWMyFH7QYg+bAZWm5/GWS3RhI3u9yAJf89wh6
cu/yut7XrvwcDg6B52SA0ET2bMcQqAmiRPTirpsmSQ1JWXZJuGDny5j1y9ia/LG4
nbLEo4D27I+AgpBEniIbo/0UiMcckaZY7TFYSbV8QhSRQteT7fVuFfYDTFUvZqzG
Fsc0MvdHPqAI0/I77V3k7whCsvuUqqWOhyJq1cdbjbU6CebrpMFla4pZL7kBuZCY
zwgyZG9ov8yXA1F2C4tXLr5gE4uVDTKDza7m7mmg1Fk2XVcHTlIc2MDlLCYjhZyd
BaeoRLr1U0XUl2iARFgPJuAVlv8Ysikjx2OWjd2CQ5KkVZ1esQrf0GtovlPhtU/a
Dg417hNhuEZTCptWxFqkd7yabxfs3X1Awqvaw19aa/gvubNGYRu4K5KEyZgYLlt0
uqDP8VptwAw67qwlwtQMXQEdzBBHri3GacUcPqTEY/C3TcuooiWD8tpf8IRhg+Lo
MYPs3e0WnLjLo889ovbmTfLolz/uuY+g5TeRT/aFVboeVsQEvveRzxuexgwan0Mi
kGt8CnM1aOx1UJVH6Si+PPKlaZLtI1ZN3Y1yjcDHip3TB5xVqcJMM+wCY3qUvFpS
kPiegOL83TJE5Gy2Vp5cTqHGwWmDbaEN8qzeVgo6wBID49dJf6OGyPzpZwXFQuEt
kNKm57H6oCXMBowGeXmp3BQ1Kdobg90ffGiEEZohewmmvd+ixqTIPdh6W+xAc3Ox
vFfkIiSapgZUBurlzyyLJMmLPO19JR8Vw9YcqZIDnS/3iqSYjg4F26u169EEjrl/
AWHe4nfbzm/2eL5CnkfBQyhUuW3KOW7M6K3auX7N7ZkozrmygkWW59gcHDIlKBkP
CrXknk4EJkEaB0FMlQ01/v19+gaHGLCqRwhTASdCXNhRr84PfIpObkmdxPRiRIfm
EW4axuMk0edZcwU8xwz8WCL2OJZaP4lKU6R5PO/VAQjofLMruWXh0q8tEqdD4WAX
MVdvhRZzE/GZePSaTyE9YDoAtXJsgpyGZNcpGuKubCNk1eFF+fdPg2h+cNgBO9FT
BTqNmUTJSA69HH23anEyCmWr9gx7OYJ2sRT88oJR//zjrFbMMmd1bpxSGL5RIER7
EdHZbR55r5A99EY1DqZd1GjE6L9RdlsZTTapIh0PrBU6Hl6iBGff+a2526TliXed
K2A7ZtT6pAQ1yQ54UadudQj3v6TPa5NCcru7h/ukABFxmIUFL2ff4AEAGxfsYoF4
UCskpSbMJjXOzpf7o2HtraKm8KjSEThPE7dxVsY0mOhURfSiFkDK3K9y1KAbB841
41SG/prlLllOoDPI8Viunmn+n951l0KTXboyurwwaWCbrcKplDQUPB4TqWP1HtJG
z4bee6LfOpN+e3tt+HWoG1kBLj5giTUoOvVOEUZ+DIrB5WAOAaA4OKSZZw1UOHTf
x2vjGXgsvB3NAO5rFIr3Z58xYnPhbi3cBkWuipMMc07vId5/9M1Cm8de+qgcVuow
9zqQGWBuUV8Qhyp5PkDgxUfxMD/3NIzH8rWNhQTtFQjqAGVomaGFfANFpBdHGTcl
Ed0yCjFot3RriVJhbjfAxqf9J9k18IWiS0Y6kvHdgnkij4U+Wmrq2Knx+1gJX4ae
3C9cp4tZMcazheDeGVtpsBzDGksbMjUqsPGqozEKbRCoiHkumvPZocawvcrMFCJg
02gz9tjTweMRKQ28SY+bA+wWJgJyufWAkxM6/oqmG4t97IAEvkNX+Tk/RiYWSlGM
M4pzUtiKEJG5E9nT0XfevHEha57mJkpb+VXPHm/cfqaRwH2zikWVhfAOiNXyKV35
XPPfbEDm3mZRTTL8B9yE3fEbwcSAMxjfn5tECmw68DEBXTqVQY/sr1tSGeRd93eG
Qb+8+V1pzN7f4IiCuqYn0Ey28bymy00Bj6EfpjizKz6/+rp/BbM20kvZPOSk0GD9
pho/FQ7de5z3KxT7cLBax2uAquIL0Sx5X+0aJdR5OEX//lDx8nxL3a32GjiKlMUY
AOrU7zzONf/xmWfw1n1MPli+/D6ftPZ4Wo/xJhjnGh4NSbNLIP0V3kyroXx0ho5c
AIh2Qol4bTQwb7udhP9PRT/mwjCqxGWC750J9uuFYLEh1DgPmp4rimp1mxkRrBHW
vqnzCz1mB/WW6+TF52e65DqTCXiEcafp/v8PSQTThOo5rDROBFOp/RTT7wq9otqo
qcACAUBa3fVoNJyl2RonVrz7lPChKEk4ah4ScygID+uHg9K8GIDyqY7e44y2yIG1
/E6n3bq3Ed92KP4TIDHmltFKiS/jbiRMOLiEue0jthmRO0/lbhvn+Aeh8SnvHRn/
5fnceDmjWt6TlDHghfBl/kK8U/Df1qIjA5sXvpITjyNq/PHtmsgo79bAKr/0p+mo
5oBp89IcoqjD5a+ydSlwneVp+e3tMZA8z3On1bx/GgrZVp9M+jD/yyg1tYTCdVfM
GVj/Yy7VU6S2x/6S7IM+jlIAw36b/snUvDBzLkLwG6JNJ0Pjko7a4x5rszzvo3h0
gysfXajjv0GTc1JjEKvOpiGKKrEiAc82ms9USXFtO7Vqhd644YZp4sOe+hKqj18l
P7kYFZ5cdeICddxF9XNXmoO8KasIBsX08GyNLyrRGkQOqpJ6Nf0wJeDSKMQsK1Vg
O9SiB4KxyM5TJbaZzKy3PEe6QU5PGFkLxozbhG1FsBqQy7toJyyw3KUO6bQHdG4M
cu5xQ2gjLbusL7HrANYoA9aqt2mFv0w2QJDk4nuXjI4dcfKSE2zx/LcrN11Lr9eq
89ELtsLk+1Ijh/UpxGFflhsMcnzEeGyxlRbGrEOIY0PJsbwh+WIr0dzEI1NBLOtP
VM2wsDtzBtj/ShZ1FkuQk+k2LiqwpnwDt3itWSd2E9VoPi++ecJHShz6vT3DZv+Z
sQu98gtTZ5liC3TXrv2V8ixrgqhoi/Xf1fZ8R4uUJpOYfRBjMn3EyLsuMPJ105yo
9Swj/79KRjH78QbLY4wn2w4P/ZYkHw4L5iZwHoSW40AvQViYQ6RoqaZIxD/PZv1W
tyzhYYc/1nii+U1HKTKelNMAsRocSQYsbuPELeS34dM5xiiFfovbf08WRbRMk2BI
9P/IrYTXNP6xGnIceQzEjCE4kBN/j4E1Vo+08HY4xsEUQXB1jlFdf4l1AuO0qly6
Z/3Gq4E+ZGAnI+RpHmH3n6zBCt9Eph+CCiaumf5brIQtwR/axPDg2rloY4rAa0GO
ak75gJmV/kEdghyNveUzdJTTQzsDClOrBTBU/QzDzlljYFfjbUbkluIMdJ1n4hEU
u9MTJO+NhfR0yFdRRuaWJmZSk8z5l5wAuWRL1RQPqEM=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NNi5tXy06g0Y5os16NmKbJE4luBY9s/q1zEIuDb8nGPx4ONgNqVPW1gfbsEPvLoO
3qrJmSTjOsH5ZmU9FmU49oT84ONDQIOIj4brIAxIbKdhUfMCNiubC2QYOdCrGK7k
p6y0xooCCLnIlD+DRaKO2iS51SIaQ8GmgShp8d/aw4Xp1VegLEiLTsEB8D9cnJi9
puYec+e5iiQEmmQ8CDDTzjf+iucws1+TcJSv57x6S4WQoH5cM4tuV5HC8hhXfPt+
EmCxbvx/MiXsuP8menNF3+QMocHccAw7Tt/pbBr+F8zARtgNUUn7iAiIbuvgcpxE
dJRHnWtG80nlEGAcLbtLuw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5904 )
`pragma protect data_block
lYo+uMq1f1vSL8Un8JTgdXJb7R+mmU4PWEa3xaAKNCfEI1GYA6F73a5rLgBIks5o
DoLNeAuswlKJ3xSvdvYAeQwjSSUBWPQPLHrMy1mxaE8pgs92JFvgAXYuPcWWeTsC
Qas8iHMgs883dfwUw2k2GuzQZfOdaJLZl020XT9Kf103dsMhMQhXWtV4G01IhRgQ
UCjdoMIju6GJBS/A24mWRtUDjQiXNMNb/XB2R3bgAroDavVIwpHKX6YucIYdw0sr
bSIOmf+aKNaz56t8JcL3wVbitGBsSFp2+fBrFrwYtQ7crU29QpI/Lzeq4W/dlxui
zsc2XQ7+hJUpVsYh3SdV+i9Z5HgcX4yaLqxZcNtgPl3BxDHuWXiHBz+lANALNzgi
pq9TiiM7lMJo4rJNEfYC6O8WfMXsKso3JXS89jLDfVOEeUT2lql5ZOt7+b+ZxHbV
9/c+HSNKbzVrPgJowBHUQT3ishMWzFuDkA5L7UIDVzlAi6yypfpAsYV9d05pR9TZ
CsQh2S2/FGVjMgmqljAHHrp1bo/00LFhJqiMyjH3eoVkr61fj7kAmUt/vzzFTJs0
0pETp+uY3cC7lVwUn98KZ8ECVKlPxJiLpkKJwvUNdmJCsyWDpnUasr/XbEqFJEGv
2KYf/7im86WbPxwXtsuPT8W1QmUO6YisyfdZMCzyxGa1+DoRIyCdJsV8UGqb8N9u
0OcFneYO4ewYDSEjmqLeSkSCjpVHR3f85CKSVofhfRql+LLTK+8SyRqUP2Q4dG1X
p5B5a4aTCI6yVBRqSOFt5k7xbrX0ZiezYwqEQq3ReY5hrjS5A7KGa0BSBng5C9XZ
NcrHBFHKcOfpICt/2gnGoxkV1lfWWppZN8UEge9bmGsvZw+tBKdxFfqQWQMPep2v
VodzjQgarzGye2r2Rek5sJ5IGaUd9EuKwFYRpnYet8g2WOApmlH4WrO1rBu1WgOA
cf8ocfuYde48UKu4QvWUuQOHnbznDBtEzrCq36n3Hh6lMNdYn51RUn2K1JXQy2fq
dacVLCwrBLAWLYUQ0xdAAflwObKeh6X4tDUZhBfhPnvEwf+WFK0y6Rbs27Otft65
8fxlaYyXVYw3I1ZMTDv2EBb/ZwSPUkCOYmiOHyGjWyXqDinrVJ/yN/N2vt/LG9eQ
rU/qn+vnXRy6lGCaat/zvVtiQadlzKDYIeGv+kpyaYb9+yPRMHi4e5QMtWaWcsN0
xe8qgXMOd3nr5H7bcusxiv385MdHQkySqNGzDezgxsaYTvaBogfWFQJDW8aqvh7f
F83CjO7bulBPFIJwddovesFdFKudJ6OitlU8dG6SK9f97iIwiqAnAIZHar0izgpD
g04z+24qL8zJAiM4SZUaro3O6rKdwzRTFuLMerQOI/pJeZ0DDr+PEkow7JEOKyxp
AJza6Yh6CarkzFhScN1QREvTMjXEHGdmAlDtNIfXf0MkjRgkcfJHk2yiWpyKlaVo
JnIcok20lxEiyHIUFgfztGIJiNKIgirWlpsjEGuXmADqMya8HyyhDEZkhO5cKpoD
vOMhJhKj6PPXKXoU6y2+gOJJlevhrn5ZzfJxpXFiOuK37fDCcMimOtqTwlvwAVWv
Sg1DhSGaPAqlxy7Aj7PZi4PNPuhLfaTezKHkaLPyCXCoP7EgW+zstNFkIDzar+/6
ip1Fk9eF5tnGrSX9YUA4RraBemIINdXzlCOaaYDlCPCRxH6NcTJDZOkP2v8ZFnKX
mZmbPTWFwgTQ3urY5amWpZ4/PKnWcSExwEWVoTqCWv6idQ4/9TRCRbM0+H8grUga
NFcwpI+CTD/LVyq1FN8YnsyzvDn9Hr8EJLjnQEDXsN5qWgqJYSnQ4AJHIDb0tGbH
r3x3hjyEHdfPe336OC/1XwmqoeliHc0JSgb95b8+M0FXhDzDkOHmPrkN4Ns9hZ9i
IHap2chkkej+tXKQqJ/wQzODEbm29bS3YS7arqePR1mGdohRIrof6fW05QJxWCKC
xtQaP55ydz2OdF3kYqy1nUHlKa+IOzIOChakq6vzTV6O/9HAxClJml3+t/Po/vvD
zvtNh3Cv6pQMjp0mfsmvToGD5lMtiBRoXiKZNYxKexhx5YKB7qVMfaepaYb0ysOo
BU+4/1Fzsc+3IAZ16T9tZU40bcXhC5hgY29hDf64GI6JohJwtL68bEEtro1y4KSV
RxO2/XZJk/HkvEpDsd+p+obtj6h2I9p4Nc8K1oZNoVr8ZkHckYoOHf5e+fQxtpmG
pSRpAGuwJAOTlZHJZx6r18kS2tuJEc5Xjs/lzpAAiJYkaB+D7nliqabQem0dN/d0
d88+eM7ZZPvymVH+AyNnK03NU3l/pAKEnQX8CdF5YZCyaUptuI/zCYVEY3ywMwbz
LTU2ZswuAI7TgscHN8NESu1u9Gy2n6xwloNYX8TqulrtfMkBjUVspvz3itgE8LPe
jbf0Kjc9TWNMDkzytN8chIAjwOnrfDd715uVd/VdM6ZPKQ8P6cMQhPitAzoEnLWa
VkGsdffR/IXa1H93qpg+3IRmzVZRVYMLfP9Lr2XndeG/eBZE6dFrNNanH2NwEo+D
EB1Hpy54Zcar81TdYFvbYq2tQfOmJGf0YuTbfI1H7E3ha05N3y410YILLkqeTi/C
ZhvxB/7+FVEg314sBqYVe2UMQxmaR/qXillKy5PNQQeKt/AYnf93WdDO468nzvcM
ultvz2K+DXNIm9gn7b8o1MA7BsXEYegN96/fCOTv1mIKYnswp6AfmrF951ikHNMV
9OTIpSYCL3CuzOIiVTYjo2YOT7HV+WNNqg2M6fCsO+H9hQq4EnxSzL0mPu5THn2j
oUyE5SoZdJqRucagwUYMEfO6vrOWf62ldgtjkxCKzuFBzmR96A8wxKCuJJI2OTHO
cm5ZHmGb2Gj99Hb+2Jo3dIgtONPbxQ8mGjYly2KOjA+xJfHXUCR4eZZcQ7fxNzNd
DBWGHgRnP/JehiodeNEsIkyRaSvbkIqXJA7Dh+6aqQpZTO9kfqKX0Le91nEwKoST
tTuawSQp5JBeOEUyomRNSzk9zfR60UcuvMTsQX+g18erQfS/SMDwrYfLW9MBWz1g
kDgi08amaOmJoBkDBukHZBamdMa8sfxVT6UcN7B0jNqSqaAqq77vhr/P3YY746A5
8x9ka4/MP4yZ3lKulF76SL6D3eiUodAIvriEYDM6Gt+edIERvGP6D04GhAM0D4wf
7u4SDEEG/JC+yULVY+AviE/MMSilqGTS+P0yg07ylc/5MLwl+DubaELsSSn4K3Iv
ctr/OJ11gZ4uFylp3wcfzPjSSMTyWQSiw+YaH88nKbarUbm2dn8BCd5vAk/3s71H
mCjN7tvXrjD7jzziPJcZrKrLRtZCHD24zjV7Nngs6l8msO+Pu+xvUzJWXGkKvjCN
8ij3RHsjJKoqdgy7gZi/U4Hsh7dLdjyWGSY8x+NuTWAqC95Dd6fvXZtioNgvyl9g
DrM8LHpInehSjF1l5J7VZ/7NE6MkPOfKoDvGmFcVgeRZpbIoFxF+Q9m92KVeQlS+
wxr2sS+/lYSEvvYogpbviu9RSjzdAmSQUwxpurAmms4F1S/dsCudxjWbZ7X0wHpS
+OD2UxId81P4UQquYxc8iXEVCZMRdBX57UeCnnFilPunBcgcbOtWz5Pti4CWo5Oz
4+6BnCW+57cAx2bxM5KGhTGGVXEOH6Mk/J1tiffEZ+vHtDsExkncVYjxYf/N+Scy
AJ2ZIKp1Ihg0FqAZaT1xqnpduIsSfY8KptiXMSev7Qfn3mWsdvGK4vgslFWvxZjP
3XY4D+Tw4WkHpCiEXbKRwM+5e/FjaNJUW+fz7bCHRfmNT1zpAk263gphvaIjj2Ds
9YFaW720Lvp8/iRLBSXda6zeUvknTZSl4ToRV/hPvF7bAtTPhYxekly3aIGRIYUW
/QTW2BUTmpWUqg3npD8wXgJpcscHGQxqRTcEYUGRFGzsXsYRGCIa77Z+nlgBjkAg
2mNb98ltweCOElcpyCkkNU5ImxhYlVjtB3Ietu4EUlHlbrKI086doVzIZxMdxj01
EhGWlEXlvDhzESllDWfP7aGxdT8MitAuiqoJ8Y4EPvmvi3rQUH/DNWXwYhBXMCcN
0/C1Yf1fEmzssMoCGAcy5RMERIrggR7XYfh3cU/uIOiTBffZTyRSebALy/60n8Ap
xwn55M0ru9sXZOjNuOHEpjfY1SY1NRN7Ea/RFRni8v0wxZL6FnGI05EdM2sEoN2y
mmFe/o5j9pmEtv+VqmRadyXEM/OnHxmfRuAj5m/xktV9zcLKUWkEUvqOBb+jtz9a
ZRIv6fF+10jrDCNBJN5NCvIRmyzDlcM35GdsFUSK4U806aAyKEoGKlB/hqkr0pW+
786zVoYEpwGdHoiJvWNaCY2XRSoZKO6pnSagv1jg5bnwO6daxMBPct4V1dpV4Et9
BMfNT+8/u11Wygt+4FBGNwv+T47yvGF5cgwqxQ3CPTnKN6VLVp3+calNc/pyjjEw
IOPVKpNxIFFTlsdDTQcPurYdcKZz0bpY2VGaIYVebFcFZm2B+lNMEdP5vh2kBYGs
myAYsBVqHl5u1/P/VSp3ohBme2djqi7tsS+KQcYuMm2Ykln4LIcnWWFex4p+7GcJ
L2OYyu4F0jtFu8jJs4DHZKUezjilPXj7c+64YDYR5D8VbzTCJitsvGnHbi4KY0mW
Rv4m+nIAlEzGhUp1VbvRIb3xRxaUUGERXVXdxyNpLCZuMW5Z94kP7PtGEbHASHRb
oXGhPrp5flUWkC3cTzbhEpNogVqdHKHgVOn2NMny75pBfPQe+ABGmqkF18BNCJss
tXJGdH7WHE2QsNChnAd//2K7xF6ps/9C5MDsxHtqJPyHJA/FVV+gZkLZl7U5mTHd
9u3bSnsId8jE2TP5KkirupEBRmfGopi6u4c5Q7Fru7pPmPsE5DVyLLkENA6IciHs
ddqxVYnVz43EzFEfx2pqcHNVYr8Txt9Bq/jsKeouzkG642bucyrNUaXPBAGoYzwa
EVJJjdTOlfDVbB13Rm3yFbn6NRrYypKZ4lVKo9lh09AL09j2QiUQy0gqKHEoPD8b
wVshFhg7HuQRsnFnbMArku0TCqhPFP9PWbncY0x7egs7D+Kq5dGzOb5r3rWVl93u
KddLvXDxSPY5mrvmdOl0ANxfR+ngvV/jQdAwBcHFOcMHoyIQrhc8w+f2LLWz4ZSb
HpNqPQ+aj/Dl9EjIurUGjmttfxyRUdQNyHIpfdWEFpRSoFI7ex7A0eEs6llTelXU
EDOXaJ0tUZPWGE6fsidrIzvsBKaPCz1WV8S5alb48k8EARScmZJJ5xNDrDuc7kec
i2ugjamezmJZFmnrLytW8/D3FS+fvo8MxBGdpTu8re9Wu3HL1HtriqkSjK/GzzIN
Z5RKl5RlbcTWey/JjhxG68CSJgb54h9xtqM3FFr6vPeasvjKgwQn1VfKq1sdssnP
5TXNiiVeoLjMBNThEAwJfuTUgL1s5nS3JFLFABcEz8olGLtVt6BwCrvGhVeSKC+Z
9hq52D4bDSKbcHmwPRgqE5xlrtaSpkuKTbaQpq0aUMGGanX17L2NOJ2wiOWlsOt3
FU6HvkxkfSPUpzUqFQC1ZkMae4hLCkrVQSV2g75DVqzj+yWjmVGsILIKniFIrFvi
YNJA04/n+qJqMI8KzfTezYI1O1JXf3RjycFmdQVNKqK3wiIwbFuAHTPfPFkHxycN
uFAqwIcdelpnkDeSnZUa2kvRLsMZcJzQQ0kpQGpj7AjEnuQapjRHH2cD16fpKKI1
SMb6o0SchzIhN5QZ+XDyL1EwNUh+SPLrrFqc25KWXq9HwUv8O+yWP5I9o+5nCi1f
02N6gIx2mg/DXnas4RP+nwgv0jMGyD4V454Ggi785WD08h0IWmX+D9SIyEM5hr5g
Xdq3Vy/a/Lj53krBKrU6V36j/Ys8snWdr7795PNwhSCaxLt8DbURm9DOsrMHuZva
gMm2OpJbyAhlS5cO+IV7rlqK/DeXR1kBFqG2T/DLJssHaS63E/Gkc2FDsjNBAqU+
KD6NxFRXuEgWkbblSgvMmijbjZ5QhgJG/GkqaHVFjy2LqfDjrRNUGnjEwylc60Cp
MCI2ga7r6szat8tuzq/xknFefLyChgJvzDI4Htnt0PJar7N27F3SjIP5jKoPiZ8x
z/NA6TJdJMyAHP2gCj8ydus32gfCuHns5jjfOowuWhE92/nxGYiTpAiqlE5gReKi
A3ivK1Oie+JraWJzyaDKmdoe4HTobrBTPacOa6PfrlcMBIQwmRdZP4oD3zMIQrwG
P+cxEuNv9MVODe8CiMTQ0DEY3ztM1nBWp97llPxVZ1zTC5x3NUUFhxt6def54dP5
Iqcb3T3IoHuNyBwvVhwLh9nIK0NTvbL0UikdU0Giv2LOux8zpw15ZIjXZd9lX64a
hRFl4HyDbE0BTco9EJH7mlHWYezwvM1vNIiszUi9994bmaN7uQ2gD/iQt7SMIRpL
+EtbGiqpFSr/0uv//mobgEkx/NzjWDH2+0AqNqeTaQg06LpqLrkuxnGG4+9ENH22
VKHwApndmqlnrvo/SwT3bEvMipXImZbhIrPgnkuzy25yoXdY8tHuYJvrBa/+Blsy
gjMYNujUrd8KijYy+xts3M44l5e0HypjyXJCgDvBd3tugbNCKJ2cwClqjwwgAlOj
sDJxvyGVrdfcP1MwGb3pAtYsy9FtzU4x3UNDr4tOJNFKkoMXVD4eS9s/fXZWgWaS
MQcHuRxMIq4AxleaPETKc/M3NE1HIDEHX+Ndi/Mxwo+51L6kzHNFes/ABUf8xEtm
z84B8XnKPoCGdy0y+m/Blf5eEHVli6Sv/5nYKqsto+BDvwbfoGRl7/GQ3jzq/ycX
nXtU8GN0XQ4LdljfZwEboaQwBdy+uDOSDky8Q/aCFhOYL24GoyPY6gcKG426fKOy
cjFxoC+uNO9Pxr6Aa8KVwXRyKVPTJ8nng63Db+FuyvM4kVRYaCvB1Qzx4PeZyCIJ
b1oBfHz4sPaeVst/nmMuzv1R0o6lR2GDuxRxEErot7W0eVgD9I9198/bXOcH6Zai
aSHQXo5SeE/1esO/b5YGKqjBmDAGReymwcCNSEyRttVM1KNRytMwXUJaQGHe1j87
hrfm5s7jva35Ck3yKL8SubagaHW2XKMvmYGAm/oKnYtChigTPbVQ2Qh89Hgjgpni
z9a/WyXbKuCw7q9kQ4ixzEGHrRBOhYbrn1kgHI19hHx39NJGo/Zt/pxjXuEUC7fL
tiP8/p1MS0Fyh4S0G0GHuOs1ka0PwOJFVOM/b7PTVoXz5OvMKFbk0JyEVgG3BoI1
XU/u9520TyLrUVIvFK1s7XnAHN19HoVNVGKNyAO7qwAzjHb9p6koiOLRSbSRlwjn
xTYJlKUI7/XRFvqdiXIX/Xm71FFHwPXP/VXBPQHR5PmcOW7Ct6Wqs2VbFB2ofSls
difNRSd5VAj3HOtGCVUScZWDUgpJ+iUaMTggg6vxDN1+q0eOYVMLCyqGhBKRsrtp
9r+80Zt12glGov+mwlhqYtWLigzwPDal34kU/PyF8MmC/egJ5erFD0Kho/Urmkv+
Af9IMnlsJ0FeQ9ygdeTkq3QLr4nCfnMBQ+3Ssxbdtijcj1jsnQMSEq8gkpAq/2wZ
NDXb7J4Xy0Nm6bXMVF25vYhieAUqA+mP2M7NMsEn9SeygxtIQajFZvGp3Srvkh3R
t2Ayu7ydGeUL02hRJk0xQiIfA+6P4cA3BPCMADSET2swjo45X/YlwDJ/D73Ol8Zq
alqD8D9P3a7cfrlpQoHVd9a2GMzPw3F7YPO/poZ76YUejU7wLKg35AAB40Dr/vmg
1pRdo+vyKhkdpd/WyZ5gCGZG/yVh8bdq9WWpwlJ1YeUjOnVAeVw+kki3jfimDwsa
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
g9GmXNoTTKtZX5aRww7aZ39cwGFxF/tG3DyyfuUKvFCl2vaZrBdraVyLfziWrc09
Tmg+uNB5DMUfl/YwlMztv9SZMkmHnNA2J8qhmEpYSny4zaYz4575LwdQyu/jQcoA
GAVNqcRSbz2CNBnX0NMr8WqsPNxRb4U7SZ6m5l0Q1kFq+GjInSb8MtyZG3CGoZPC
ma6eAUhueC2mLD1xsTO5wVxXaq1xvrk99b9zKm29VHPn5/F76F+V7GaBhlyxyWHd
EnZ4BtkmxK3LiHMwWZzGGCFXm7g0RqgNqUlNriflFZddXHPQ3jE+sUg4D+QgAWAX
brr/Ug3xjTgjuQ4ZNUPErA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7648 )
`pragma protect data_block
gmDSeKJCcEBIvd71Vme8TfUUHKzWp61nrul7zuVHVfZ++evADfxswO1dfEJ8S5+D
ffmK7ZI/2JV7uN4/UwkOGeC8/wpARUJMUh6lNVGlb7Q+eBJV50wjEIcqQmISRnxV
OH6srJiFw6nrMKbrhnp9RQwrWH91TtrMjMmTWEMweFb/eceMoE3NwwvxkKf8blHZ
v1nOhRgbJ6crv7frYl4ap4rnrnJAGbrXm6aUsYBygCh+BqnyFfCH4c3+SkySRyMs
CJs/k29D+QEqkHBgagkgNihXi8qrAvrUXbhSXexR5Ns11HeyW+4JDIdFK9g6J0va
agnhYOzle8WtuI3EgjQcNFWRST+fV+wqLkhUQbWpkR27CgX0fJj12Yc2dr/+hcIi
4zPei+aogpr2TAaPPn/1hPI7dO0l4pdKKqh4LoJ07Y/smAGp7YTvOIdMoWjMKOPa
ED0GuyyRoslAkAXtNCz0ZXYchwk8W+SFlfrUM3bEZQZOY9XzauCBAzi+XSLdjLin
znq45jw+HhofjGcdrGFL27gVlFwmL4qtKF5Wlw04n9X5fteXlHI4wQ4S5j/O1z5w
PV30PP/YXHWAmFAk/1g5CPGBIWGDtyHJvnu/2aJoBOBdMHucUGlRsCPzCOqwGlni
hwJSoCqbI9dKtzU6fworLIr3MpaebwDyVDrHV7/J+G52/q4ylwdKRrdfBZAwhdpU
qBAShbkLwlpKHGCaQqS6OmYkR+AS/dStDV8RUf7NdG4rnXg/hZsOjNclqUK86Tlg
W5fs6YcEKYmKgZUQg0AsBpQLN5SJfpj6LWE3i9o5WeG6tH257zMO53OVybYLeySh
QpK7N6LdobNV9OR7fc+8YfIOEMKm8i/lnmoC5JPfTHHWJBsWznYiNWsD0PfCPPFw
RcmqZS3wqG0KNCo6UPHKp3ptVDbKPxDo0DBXGTvKfojGI2GyXYc1gArJH/Z/3HNG
AZKcR3/giHu/J2byO8lW2Olp7YZ7fUDTI/HxEYvnSGbt48JYyHs5NkwtBM3pjdze
9D1Hn4IxnxbKfaldDOCZ8fRdAODSj6DqNZBtfxptYfWg4Bz4Lg6Oi3q5X66dA2n2
EsrmDGT91dgFYJhlhbvCZPYYfCYZIeRtQYXEHU5sJZJmVDSwqWGcQyO+i8l+VL3I
kuUBeB1s8dlkoJKaU7QVWX6asdFzUoCNpXLI2xfy+sVsnOg04qAq3nHW+kYqegYf
ibt/Jd6dQSWnjqx9Mc6ws34Nm6JZ/12LVKLKnOms8lDFaScDBQ3qbHr3oL9Q2M4k
Tq5Ij/35JdMX163RVa2NAa4btb2IQ9KZ3qFj9Ff+bQLTsxTDOE8Um9IEETXx4Jqi
S4DazIzpQAU08QTFbn5wyo7m1e/DwIJiDdveFzELFalATtu1bgQFCJ1OH/dzwv+u
0+LMyvv1pPO8I8egCgyT87ws6ox3knpwPSg3lvwDXi062qKbFEfkfK/Gl+M0WduQ
zd8anit9hzKOpmjrX0gOFBCUkjOECRK4gyE74t+BYrci91jA/dELwQSkeZd6y63j
2mff1Ka5RR2yk8+PzMK3+fg+AlkgQYnxLGndVK1jCuFgJm5uvj6RBEP/D+xN6K/z
c5GVJ7l78yPk0FASwGdkV20oo0em8srSBGeKagwYfZf9XRwm9sHMYY7fLz4zdme5
ceAg+nABS/2BnIefJepxZDxxkg/62ruBWXGqsVArV4hbffIXnu+zTaMfK/td8niU
wajsfHtF2tus8cDtdLRPSmWOJQSk0pnHtOntC6S/HBSB/+AShhM569f2ZTWGMuUu
7PvbBMX2t65txLtibVjQYTz8wGMBWvqXDyht2IlMFwYW8mxWVr3bulgmA+a9btf/
ketxTTNhcbkK8nswjkGF3ZeUTAr5QmNOp6osPArhyHqqzHquSWV+Tk401P8J8+hL
GRnc2txlmPLN7fg1joR0ae4yGUwtIzA1QOu2UOEc3hRM72nvxkq7nwy+aUqdsnS4
a0a+XScZU1wLoOG1zcbSMM3wVRAjhj+LDY06GciGe+MjkgaJbqHWDT+Fyy+opGDC
yVe4tmtLJNlizu410LVELEa+2Ey9skFz94RKicoIaAP/kBdZBZSo4SK3V7vnx84t
uG4oykIE5Q5EdgtcmJkZMP9AK7B9izqSkLS+a1xIOqNueTPlZHR47sm2wU4IzLij
MaggfP7n1xor1yApzSLgGWQYj+mjJ0bXf5iQpUC14TK+jt9BIHZluBowIwBuaLY9
Q6SrMOlScmxFyKlNqPhAtuKQjsICZEd26eCAeWpvEUYnD3mRIzm/38rJRYAyhhX9
fTXtmoctaJAOkSyrnTJnkW6SMoz+gSB806Wc89FR+mvQfibp8LepED6Kgpz2S3Jm
kPVhOGGP0uXjRz5d4eoYke5tmpar3Df6DCog9mWFp6mHQfufozXlHzKfrWix//Of
mc66fos/+Wxcj6MsTIAz4itYq5RwK+jVOGuxl8WZSUyKfPHZ3kpiU/jd++aooV69
YMTMfVpyYyvVKNZHl2Z0kuVJmaDeOnyBMvLaKpCSlOPRaKQWp2HAIm1B2+XOMF4E
ae4NsrB/Sg7QkLsa1DtxBXftU8Y4hjq4C93BfLEDPbFYhAV2AK8uu10ixoncPiGB
P8V96o9Kr8Rzz1hubGPZhB1mkofNWN0x6DggtVWLeYkHv3i9oQpMHQAxyp1TeDH/
YXGIT9Tmx0l8i2bHfhv9a46AhtOm0tfYXB6x5qoqbOFk520ecksh052KufWFAPcZ
NptT7g7dq/NPhPMbgBarqYHeP4+U4XesVIsuk7xNNfSBKKOoN37sy9ABDb8YaDmu
vSfnd4qnAF6SYmiB98SR6DIf1cuLaoLxDO7nGEnJPJh8P6rcVLU74bC5Dxz5tROt
ehE2yhFn4JORLRSIHq95hnd7lQvrbeAivwHuIZHYCc/n2OzbsNQZEQM7RSpP2Lg7
l9CvzZ3S921Rl15ha7KZK0xu1vLx7YZB8HZ49/FV6BfO7yf0TYqqqphJp/dkJ49P
0WshY5aw78g71wJoI+XBIDphwnv3rkrKd7AIkbLt8rpF5ebb3Z2hImdi3R5a/kZd
QevFyh4cl8rva3N/1iWNGrb3jZHB8GIjKatWKjc8GZNnS4J5H4jqTEIA5LR4Ixlv
FPMts+NhI7s8tbsyPXhvTTnV/x6UQO5WaFgDJAsJ6KwAy07wLVwwyz07GP/ELcV6
w7p+LY3/vQzbO0PjHcjxJsuwp1pEqGxH67YUA5krb88FbTbtY7VGAIPx1QrCUSeF
nJnKoXp03KRc39et+JauMo9s0zTm4Cp/QDzAa020VO1fhomIiZd/BYErKz7XNlrL
+USodLQiLKt4xDLN/6K5u4AX3VID52QQ0wz7VwimvGWKJpD0Laqo/96+jh6pTp55
nKaHyO1PE7A6PXPLWiWpwWgOqiJ2J6mDrHV6KvUx/Ufisz1MHzlO8A2ErDJsmziI
GG7buEtQNadR4xsdg4zso+R70kWip/3gQ+5VYhjWDGtVx3bI2NhiL+m5O5e62wwJ
raACVabfxFEDx684k4f/zIGFU998HfYjtm9yD5FdTFvATthr2rq0Y6s2v7K1kw4B
oMlCyrRjcoGge8CAczSYNv8rQB0CGoLvf59RlLNNBhPK/hYvdYtdi7k00A1hI8ng
g6C5l7xuwg5PMy8iUAefPh7ybn3yw6kpI+FVs8FCwWUKbJ59c7dHhD6KzMZgREG3
xb92E/LmrrDgdA6rwPVZ1DBjTmLKsMdOcqO4W2JrblzYdrLmvPvkCM4O1DzLc/yO
OXVLMRhXmUhrn3LRNw3e9faOzYfft/Ja+cmLIqm4IZaKX+Pb6xmA5e7tlUH0aSyO
5rg2GTybzWeJw0zTm0d7/5N578ukrB+OC3EW/xdty7LnLuZq+HdcuYxpQOaWMYeM
d5y4oEFJ0iJMypKs4+zfY/v4PtQ+d4FCN4bgfe2De5osmvZYs4NFnGarGEGT6n41
6gQNBrFL1bE/50LVgYboOU5zUiOAFBDCoYW3yXwASEF1aAx/+N26LifWz2EHdsL6
n2WRmEncb4HqdwxqdHsyXYjVreg09NQT7iBrHmUSfcvm/ktSOSON9i7E46gPRfZ9
puefTIWic7rk4kEYB/GftMD0VJqj/5PYs9Cx6MMWG12oNr2Bu3FGpW4gjavUrLT6
XzjOhvbZ9Jp7zOK3rYnKuer17Zg5e5L9BL8RsYWQfDCc/ccNPwGFNIG0cadIVD/8
78rkD1So0u3xyi1MkYyNwIwd7oktJDJjctx4FKzD6S13CxHw3n/bJ0cW/+vKspLZ
2MH0Vz1R3lkdncAibuVt8B/aBMZGg/oIe397Mj823ac8jAltvsea6r5VRRlum+Mb
B13MvrWxNp0D2qnGYJZMIRhheySIZ1SjcXh8BDs7zcARcQK5/J++R0S6IBKFOiA7
fxSq7TiZzSPLufZfCN3v//JdUPrhw9ucOh51R+I9RQnEtz9gXfwV5aqHXS2lHnHQ
AohVHcrI2zqcEXjPBmLoxNxknNhJ3tEyZMfxoKU1iKrd1SAzeJJpPry8xC6J0zDy
eBKEDMZXmKmrkhyID820DbK7KxKb3Jrgs7uHeuDrkd/9cYcEhzhlO9VteAy1/K2m
oeSALriieHeIJIIWmUnc0L0BUyYWnXcfMOBNOBqvuq4s9RcjKnzmQE9PV66Wkrks
CY6S4kfyOSXUXzV0x/jG0FYY2J5ihdfVwW4bRQ59VxtlrGd/jXsXTu4zvPzBkbAC
KmHACIT0ojgC5bPv1hy7gpPAbKpnva+cx4HO9wdL3xiy5Y+TA0IUS43+Xfj66NnM
Kxd2sjPkJcx2OzmWg6MTqAqj1VIQnznEzcvGERJP1rw17bAAFOuL8fEgJzN+yMJb
fK9mfVqJ6uhotR33a0jJKdPo/L5SijFSdbO8u/kiNR8+Vv0TpbjAupfixmZ4f6lf
k7d2BoCU/iRsKwzDs/q/xoEXp9hlDFUhNNp5jazI64t5sFTg90VqJGBayDntp2mk
8Gc3tIGC9sEFGe9OK+89N+vIa4a2LrDBqlexxgiv0zh/AgmWAt40LnycGksVdG5L
la2ZKj4H/ep9ccCvdlW00hODXzfl6GFVz3xmFv53x8x+8s9dBJ237uQi1aPRYN4w
OIaCIHeaS0hsKw7inLxBs4SD6eFm9LAEWrs9gerOxS37L5zPrOD5GDkR7Q1bPDhi
2cTVdmb61DNJZABrvF7JjqJ0rGfatGRQe4KlHA6cBs6Gs9c/0iexoAoxdsTLVtcb
E3uuE5O03Bx4UzTWpEHoBTSiBH+LU5a7BuckgDteTqnhv1CBTjvjsCfQg86lKTiq
9032/VRkUwcXEhZgJe8RNp924DSW4ZHG6brn1CsTrD3c8ZbDirWAN1EEKSKLfSUB
dgdlA5TeMOSWCHB+9w+0JjTVOFjsrKvlsv+DB9gCTdkcDoNsxnoko5C02hkTFyuN
kX37Vs9tsgVA01U2BMvz3tHZ4kSd5IKT1sdxP6AUXaryFLsnzn4D3k7m8AFYXvTa
ClnAV4dewhp4b8/w7sRTKHPyChRvdNva8mKr+Qo0pmX4rXDhtf6i8fsaAV5KMf8A
V4LLFo+8R98rddVVaR5LWO632sCgDOWmBjSP0alHzKFiVi3csgwjtqCzcrP7iI55
+xOzui8Q9rViI9+NwklbWH4px8rhCWT4vKLxq4mWQYo7qXI/TLPLeyEemWrOvA6e
e8CNxpSen4dSngmHfXb6FpQU2CBM5ElFWg3NoizA1UtD9FiHZ4q6gPQSXzmnxM32
0hv2WlCteXCIT5XZjier8Ux76Cuk6k0cEQBZKp+jUk9OAe6xICf/ihtunyc4E4WK
z6MYX5t/t4Iq6mEG8AH9UMZa+Oou8V/nWYndyYZflAeCCeqSCW/jWscsY94wIPG4
kC5ZSOYvp91TLTcI4aCd38Li+oqVlKMIm8+IWloQpX+RKm6dsyPTPcEMwroMswHg
Sn4T5A9nSrJUMC2NycsssPFOlyn8UPcFdQCw3ipURPajTrdF0GemCshlbklh5Mza
ouuM5d17drQ2J4uomBq7avsCkX8izCCTDHyMxzHOfr6XrvtVT2lbsa6CjYFnE3BR
xZiWLzGr20eiIEafZWylgmMhozHJKoRL6KkuMBNDigKyJbO3H/8cpcisCS7wq6ji
Uwlv9ss2F6dg8iNx4QaGEB2UxHxu1hEFELyXuqN+WzhT7FDDfHOT3B9Hr+qw7oWy
VCaT+vl0ezr+i+Q3ArA3N19Q7Oovmmhym7VJkokMvO2H9Ix/e1ir2PbpR5YpYGzG
7op9ahvGTaj+lCaYsDyciUXHrGw2VMQtG81K8qQN9dULP/GEEOKNBpV/rEnzeZAG
fig/zJNaO/lYg2q1hzcI3u6HJCPOL8VKiQNYCwMkOScWM5HGE5nwwbQIOfsKDjHz
fuv4Da1UevF6oqfKm0vDWvscAF8AwC87CqtAIY7QOHgxutSAtmqxRO3Lh7tOlonX
ySvVY/O4yjiItAEaeqghHj0yQ57pDH4ERElo+PT4CQ7W54gz/z5KX7FqgtZAwBnq
FuRRjcS5F0Rqe9A1+Q+WkrbtQ9SS27SncqQsePEGPmqMMEUN4KUH/RaY9HCFZJd8
MbJpcy8tCTXhGZ1wZu/KdCcWUcLgOXzCwWENI1GFPrsKn5b46TMQSt095PWfSsWi
WBMij/Vc1bWbviAC1aXqEkWcUnaw/x+1LVD59Jyyvq0vdpBJ3Z/Xtt9Q6+LF9bLg
ch6DCn+qYr85+nBOS+oGMTk7O2Bhk6fgnjLFo2HCzwtmNmd0TXZPCf+Zb42RCSRK
1EXSV4GIvR6N7NqKHUaUsRSfE5yS5IHYdU9ZCCCWBS/uPCLsI4rxe7hXkZ8d1m9Y
wq2wcZC7Jlu+dTDExu11csb6gvWnYppPDZUOYzrGucb66DpQxxwnsd7O29hXj1ZU
vknsEifNQNZw8PK4dbMQA9GOOBbXxXSqMv7zq6UdaXMVlWfs2RrgIMPWrg1C5QZg
iS5oHwIinlZhP/xfi/MVVSj/b8hFIgaay/3mSL9nCPd6O/kTnfeIioTGdcx9nS2b
dXwRwOLBGuBx7K3Z0YR7m5WX9ZANFPS/HnnWgSQma9HCJDe5SGLE5O0UJW248vcA
VBy412hNrcDakyY3kKI60k2Zyyfa+MCm7I9k88yLzGxLob9IwLPi30Tqsq1lnAZr
zn8axn3KmxHutZMW6Z+hDz4DjOhGeonklEgbSHacgKIUcfttHjDuyWQRrY4IH8vV
SLsLbGnkE0X+hAdI8BTvCdK7XMDTprrHjLaVVe6B+MS+e6NV1/l2RIyXClyTAYAE
qRa28gRRFbFletf3JtYsEOz61djiu0rTupeYdNVKAz+rcNpVW+q4weXB7Zqaxvc4
Wo7BNaN1IYMwHf+S5hX10vEIzwUg4S6uq5XnXsqEx/nmOFKUiSH8X7aXbiEK/u/j
LApyOR1JDT3XwaCJ0kZU2h8yvI6mSS77dhp3CFvWn3jkSnKOIa1kxn8togTQkzB7
LrAPT9x2uKYqadHeR0NV5gbcHOJnjfBclv45TJKHoD2RLLoI+XjVMrYpysTi95lE
N06l+YMlhr9NpZPNoIR/USGgmrJY8GVoZbCkXpNa0wEQkfF2xjn8yZe77j28NPWa
kAtu8D8dVZQCp1b9XGAYNOr1CTlg5y9Kod17CrlCASNeAmdsCGeydwE/WzoP4L8F
FSXG1TO9Tyn1FIDS4s6eelyZYNan5u1f+Kj+eHSoQ5b01ZCHQtN7waFu2R3H7a7c
qI915lDZq+3hGO0Be481BB7c1eY4c4NSudGs9oZtMunrqiWOYUqUJ/ZMnlQOxxG6
+WZFlNAe0qM3iHgN+iGbTNsO2ZuELu8DlvYVT3zDDsPJlZ2YwaLUTURQ/L8hQ/lA
nHCUJZ4SUxpDSQohIc5Y2QojKHZ1RWd56Cio6yOE4tNoA9UF1n3Knovs1/RLeiEF
HJ7GchXATcebTf72cb/YlyCdE8dBmIKygO52u1ttoLvsxoiyDpAeoct/uKIH23J1
tAag3dQ6N2HXbv3QNTBwSmNWXyeP1kZ1zJ1zBNI3PTt9EG3qd/Od1KnXVLPTLFP/
/c2ViZ7KGxcN0sJzTItcePc/edaf3nsfC78YwnE5e7fTb49uBKn6WKpkWT5s67vo
o1DL2A6iXDeuVqqeWIuuHk3lQjUm8w1IZ3qMbpn7mKJGl58bK1KaxhMPSm65JVL5
G8nAVWWHwzPtdRCvhPFRs2BY0IL203yNnfw8FzwmznjL/b11rED0ZL/bJ8V91Y6Q
XvITksUR1Cxce4O1i2qyl2F9qdYCrG3ctu6PqsCZgQ/+X4s00GN5YNo7meoUpYtp
JJpEEYzblkCnYER910ECLXQNwM1ws4P/vQZkIlg3yjohtBZi1l/gdgSKEIAibPUB
fHUTgC4NwdNzd/Veo0UDOcDBzb4DCyaxVy1Gu55RdWH5JjVLweUcKc4jvCzg5keq
I1oSkDMJWkqViorPNRJvVx068B7cFYGsVDjkIIIS88ZiW6dubSlhZV3IzM70Tm1y
2dEO8Paq/X0Gq6TV22U8J7iKNMp+ujNg/huQ5Fw7IRrJ1yxIa0lJGorbf3fccIZf
ILuWGLRia1uicxOh3mdL9fzMLJE4VtXbPvVLboD1tgwtr2UR8xGT+GRyAnlueeOA
EkDS0P1NEaZL5EDlWvJscvz6k1Kyskdtj4Scr8RFua08b9smoDAIzCT0qo6BhPWr
hTGeJoEUhhWduco79ctuRmErrf4ROyXz2Qqe1P+sJ5c4wWjnXU1QfSESZ9WVzvEk
3IvLRbX63kwVM6VRvap60N9qMNBr7a4QujLZkF6n4r6rMy7N0frozQBq247PTLcN
k0j3hv37Dz4lfTFcU4saPE/lau7WQJG1Q6W175QF1aQcOPzDbpItPcM1sibXQvAX
ychw4Er0yveXB7lLDoAqUExeJIJxKil2VgMwd3h57t9bXPUzPtHvs0a2nbPlH1kx
RO2SbyLWahBpCTMlFEsrBWXYOECxBTUJbz+jzl7S3mrsDhRLx+qU/zxgpmheQhqB
HcMztQ6aG9J7s9Wrqz7e2Jj/UqaFhQqiHxa4Vk6EZ8g6XEtcTEiJ5WFebypsFUIz
lRmTOsz4wBAEnCzGAAdpXoh8HzLyWZTjKNr+gxvCqRzT6pQgDidjCq/zA9k5uXwB
cJQJRz7fF1HBJp+QHhKI5jfGoGklVrItSr9pS4AHGRWUF/K0wZTj2snpxy1Lp85w
8qgFZd271LsVDjTZCZoTAfXQw9IMt2wO4lp5A63JymTysLERefzqAUqdTFhkuOSg
kutT5F03J+qRoz3r1+/sazowhrgoHGKGl6u9uscZpWBHSQAaF0YfebpqVHu8xGAn
ZzVPrnj+aujwv28m76/oQz+UE4Yv7JrmCeS8BYA6QYlgIuopufCY0Lz+8bqtFKG4
V6n9n2TtpPgGKSZpv/b3DDvX3UGsBKdswF1pDkAIbb8Auyxtt75dIGHK/9IO2BjX
l0BzJby5Qn8Ux30DruZY8hZ8KanZsEcBjCnji9/fHeMTuZHFPYismoKdSkg41/vZ
jZBxIaMBhzaxe0u590vDjSMhuqs1orxW92oGgCUoJwGnMEJRm63Xv7dWdFFRhvnc
xEUuGzxve6o0lHaa9K2CFe6ls1V7EsC10C8frXPZptOlWWJBHlVpuaGEJbmzVr/M
4JLKLRMFtj+7FqHHxKNw3aYydd2hOMKRhArCH1EUEAn1ANicA6YcnTqV6/h+CfBj
tp1ubmn93k40dnFvzZSK/pJPmIxD5hX6LPtt4wmfhCGHAFdGh9VI7dE8xJutnIIi
2LQW2TwDThCpqwsEjp1qHfW/mhL+swRQiu5M6JFmCQJL+TDJ4R94caxF5QWTAtc6
jNj0IlZziPrFcJYk4lpzB2XsfuOS2QcFrPNa5jS/MuA5oMo56j8Jts9443GG07/R
HxQmgJJbtAeqm+nQEAX5KPGwjvfrXfsbfNYkP4n2RHPxMGhwWD3ZazzN6Hoh3ZIs
JPGMnFTSiTo+XbuPzRVFPwjA0USIFrHxplXIcL3ji0n4J8k85e8RrpT7hcmmXGse
6fvpe41gh2g0xupph2RVuLkcg/fwAdCa9ZatwqgGm/n1WHgienhu/ZY1rMpdLqqT
fPFMYCXpuisSce6ml5u/T87jRUAa01sAj9CBIdfrdXzR2FrgDPHyLOkesb7L+ssN
N3N0zQ0Dl++fisETxBw5EQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Hszfgic3Up1hXJByuCj5hjz+szbF2f+aZiSCRLTaQJj36YbmKwYq2ZODTOwtOGwy
j2n7HtUxt7vhroUl2u9CotdnzrldU79ypH9ALu9xElfynIf4IEQKgVUqXlGjdAKM
mtmaLddezWHpJpf8vk+dILKeVinqkElolKqBlEch/fO6ESDLkoNw1PtsOaWLWhT2
57em6F8ZyCq1lofr3AuVnnzAgcMZ8w1JI7QDQCAcpHdKwppCmpqUjY0GZRrLrbqJ
mL3Ko8m5AsBUEop2a6gnhS3GAu1J8oFTOJ4XVP2jd0hWehkCGocegcQSwFVHxamB
3Zh/07qmOYUio0ukvoMrDA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5632 )
`pragma protect data_block
pzjgrFm7wUpWWoDsDqVY8XV3DtakMpXJZDGkE0TpUP8w5rEnFkMdaOCYEnVqvO7l
GCOLKSO3QOtyQ1f8kIze14bu1d3miQkP74BpxFdNxlLUbFE7PepuYtASqWD6Hq8T
R1JsvkpPSX/1j1w5Mm2R5vrJsTkGrVrQmMw62N9fuMlXBNLLRc/hD52LXZJ3PZ3R
3eWxHXMyHTjYkNmwLwrQs0PmSX/0qfjpCFS0BhdXKOJrj8V/xtRKJ4s0pjf4oYSR
S9GC2TzTG+NB21sWlorJIc3GPhhIsXJN20b5BP2jdRu9BTpGqQCEKkLX3dX1RCXi
eunic5bnnUjLlQ4LPMq6Xad3sm1gwfzLyiDILxD7Qj4kPnMWhbUGKYamz7kbEA9w
QjgHjsNe/g5VLUA1eAQC98p1YighTxsZHz1FXIbb1UevpvYvjSRqO+YPc9aaWS3S
CgJLlS8dVIBUBJdlpydKHIkNyIwOPp6qtjt248AsnNDg96AD+qbtfQlvHlFiaIqk
b8HRZYW9sud2Olw2OkwdgVblYKmzglncdnOyigZlVaBI0dw4ai/ruvMSukBIZrCJ
8fGjUix//IxRHB4/85yqGPiHmOmhI1r/ZJjruDWXw7Lb9Uynsxb/wwpHhgVVWl1S
Bj5RYy/ir2kNbBB2sCVmS2ANaYaLo4uKt1EEmDDQeTtlKlb+mwUsJi+TDMYvfZoB
HOpKv2DGL/DEKAIHmU2+2RSJ7M3NiVMTvQNFVU6GTnxoZ5BniuUuMNnfcPjd8f68
2Gj3z5uV0AUxGe4DpF1GdSBKVkLWH0YcqvlaqxRnE6TBlWvCIZlzII0fn74Ci43T
jFHms+JVDF/q/ZHSUv3lclc4xn5GVRy1gclv7BDQr7qvnAFQ/LiN14OdpIcoc2xR
+0ApvOhrsLsX55SFpTbJLjf9nxWz8fvC0DaU18hK1fSY3kNbMqZY7jQ8TJxw6i+Y
v+W0uE6Dl9rx6qDnfgQakExM6g8lfcmSlHxjyh/sVrjHp1rRg5gRefrEsfLo+bAo
HGAMX4tm13GRR9hs7QWkXlRxRjJ2dgahAiwa7aOWjj+Fy/LDc3t9lX6QRO+mzsvN
0ccymL6gKAiMGT4htY1QKNhUNyV65o4ompnxuuxjVGX7xYZK0plZ7DxLRy0EF5Lb
BQODR1c3Pcz5AtSLIzxzCPvDNhhlSNOyrdAXH4qJG2OOPSPTjMgEGWdKnU6UG6TM
doymEZN0eNNXLHtByZfZevMZFCk4psfk5ycA/pewq4XpgrhBse+SbxYFQyaU4goG
4TyPkQUH2I4Ss7Wtpq8YH5efumP4htEp4it0QbGJjCPppiJwJRr7cKiDJsbnrpLh
K/a+W6BRWBUh0Epolyfc8rmdwbniUBrAhE7vKbs4l/0BOWlOkn/hEHNt6pMjcDTR
6ea/sf7J17F6/n4n/P7zJ0+rjC7BMCK19rOZoR6M/IPs1JXV9jWOAMmBdxPYN/nB
jnHuIaxKu8spvejGJPLZifzhlSTiYt3Qt3HU7IvnH9RKrWIAD6mvPo0u1Al7rEMI
mqWoQYn9elnMgPvu/va1B1StPq80r9CXxXkA+N9BfndY4fV3+x6fxJHI6t/4nnPk
u6pNjie+BcIEHLfuGxP5mNZROy3KiqZnTUiUbUa0zBGymBsVkwxGhuVligXpJotR
iXM4my7jnOOBdQEpevOts1g8oEb9WSEyS8JMT0rXIX1eeSOFuQswwWoK4KE1Ocyz
mQyg66QBoQ4zuO7EYQJnILoVj/nHN063jd50YCdxN1eR2in1y8WhTOVSFxQQJT8B
fVL2QYwHvS/WNBvz6WUTQC3yGCoHvCnJriaWydB0eTlNVHVuOLnekGS/NdePhNqJ
PCsawR9hCSOIYYmN/tPmMhuquwuBmUGk0cBVCH2FhawOZhemSiQHZEn7DuK9Ogir
+r3KIbok2v9/SnbxVZZaC18g7j5Ncbl5+L1lBd8/nvFmOKkxCtxdp/MCvfHQCagL
vwA3DgIgFCS7JJELfNREWJk4w4QiBOInucQBt65bLCFG8oWHT+gUm6Cro8fKb3hc
Ku9bj4HNLfq1jkbWHa19fI1ZtGLZkZSkzMPfKgWDktd6Sm74WRPNUZfE7WY/CjHP
GiKIvxE91/wf7OlvLBCTkG0a5bW2z4ODLdEzBII8eKhPE1LnxeRLbYr6d2fvwci4
NHbdxW4PDJf+rkxbgr9643+b7YJlLwhdEFJo35ApHb3dgCvuzp4Q0mlII27YI42z
zJDWXu2RFM6eYazC5pM/4d2vkIwHd7eJF1NufVxalomwk5rsby5beWYkEV5IhB3k
NFlf4RkFuZb90vxa/BDTf0HzjyLh2XhiBpf0h0gtRGMQa83nTGxMA6oQq3IIHncz
VoK7cq2FEFjC/cvThUuvJaP/GubyKYPmXYwgDqsfCwA9CXfMblHj8ZG4fV21shYS
VMgFpBSC5bzPE+e+iYNqV4XzomdxHH4/aanM04u0VaBJOkJygjNXKEfytuZre966
EiNg++m2UZR4Z4OhxbheJhUSsEtO6bbBASd4e2wmK4MVNASRGWxj4/jFWl2kd8bx
mmPbkH4N3y8e6rbb6LNobwr4q5lsECu1yWLxHbNzrCStKOP3WXvLA3QboGdHu/D+
g3n885f7/YkOEYgVjoNtY8HEM50wVk/QXp2i1SCKi/Qd+IIRXozt7DlqAwndXPud
aPLHyE5c4u5JypJc7LhBU9Op7YbtVH2KxIZz1CeMCDe3H2JSuIndNnw0tKb7MvWr
eL7ur3pfimvSTyolXHbuUN+kLhSnbPjraqh6sd7tF+lwWgMmaBIh7Ao+5RQljTSW
0/Dw81QH9SYb6bT9n0eMXYvHopQpqBD++m9nvpgLKMkxeJ19+ia0OdNvydUANfEW
ovfBrUzrrQoCVDsnJIjSMxh8gKhxlKQsw9cTKrBNGlsQKkO0+2kmFvW7EzHcvmrP
uNyXSsoqwwl3SL3UGq+jamDaojume3MdFMXjVEnlVKShYNAYLqfciKTrkQDcwV3P
2QZg6J2m6wIENoNObcyduFKP9W5pT6bzcm9ltx5XyTcjCkvAwU5mf1aYnNY8BssS
EttgO0Wa1CzGtYbsnRckVpwWru3+CEzCt6qAFyGkUoWXDcnsgPxoOxx6K1ZGZBJu
SjcsbUSYADZ4aCk4SDsg61ydw4MwLham4kD2D3cOAFUoRjswtn4OU3uVLD9tDBIq
euvsX2vc34tN3IgJJ+HPR1M71S9x3iQ78KNSohyiXRZJrLoQxbcwiglMCTU0efXi
o8fPglnCzi1Bpqsf3f6R5icyRi4F3WR7KKSK1nvKOUArryR3Z+nz5rYGhi7iZSeU
GewEA/gRLPznhcOSL/9tchU+CfgxyvSKDK3w5Z92c1VgGpYEINBcdJdj6w9jcoPW
RZ/xm2G48vP8DZ5tR0mKekutEHJ7h4IWeMoPDsVznuoIk5OyuNkT9GgVfUdOBwl3
mG2H15VH3JGBvSZRhTSfjp5g1dborGAzkq3z0wM6oTdeTh9tsJdO3GXT2O+n7wZn
WoEqqyHpa/Sfq1gFTPGIrr6t3kuvVXT1Ed6zQOMmMq6Mvye78Ac7zaV7IbXrxP6d
KnQOEBRDY9SX/e2kNo3DBKjRmwJoULEH8rlI1joX+oL7TnTI5QiyGk0Nrns042zw
uAtar271RNSYmdBadF70IpYkOPS8sL3TJ810dLi4IDrfAWQgPeSD4DrewQlyatVX
7XcJT/NYIf8KqxoeC1t5hO+MZI77NyDb4Xi4FszcvZdTAbwaFPFbV0SvqNm9JFVM
jFrwUbmdVRaS1CbHbCI1whDTEz77+H9dXicTHGbajrespmDFaugKTms25aFC3mMG
j7d1g2x+RI6d4LHDX14u3IgyTf/Y+LiG3pJWE4q+75T3MDBJqIaenzh1nSSufwvo
GP/Y8n0ehmVM0dWIiLzklIw6rXNFV9yWWbD6Jhw6V91l4+QipLindyY4uSj67lQY
4kFpKFt3awva+xYs5lcWmjqbA754ley2aXtWx8hnUC83S1N4L50xFTJvZIGkF9Wk
Xkl5bw16vpGVsVipo12o+b8ki7ZmlARq2GS7t3GyGTJSDmJvCLOnz/AOgTKfDc8t
Kw9LVealoMX7zCaDe0gzx1MzRt5haZ7HgQQBdGPm9NdTkSsgvorhuZoCw/PsHTpv
VG8ovjzeV3ZmZpBw3GojAY9Dpt0amEc/hCJ1eIuM+LemoUo7vXQSXzbPVQTfDm0c
5+f2g5NjLl7edb4ppBRbWIeiTz4YA2dTcr7s3NS1ANRsZGzg1/cEgQnQp7y5oXf1
v+CxP+B7eeyd+GkQQsAO+E4Axm5DEfERiz7v7dnVS3+rLBcie/KislyZaHEGmAdT
9Mtw/CCeM8WTFMH0auHUZlqZsPIKo8tCmuwRDAEJODTsu0c6BcyF3xVL2lWxs18s
7LAgrPjhyzohNQC4L1fL1NVYuRQvFYaY4L+eon+psqf/RjLjX5pKC+NKmOX+skbd
ZfeZfHCccqFKQt2ID8QsipgPby9ZOj7B//eGDO/MupKgBosWiD3M94NxCigOTSH1
oq1ru7xPskFn4c4TLDXxR4p/s7WIl4Ap21Z9L4zJhVW0FOCsnbu/FJVYhRivngpC
E37zjZl0cAO2kY5o7UPABPU7yZnPfEtw9KZNlKSFAR3eA0mbe3znwQxEyADIZRkF
htlPCiqT43Ad4LPqsYm+H/+LWj5XoXsvdmarVPWpvoIZ589OyA/NkzCr65ysXJC3
F9js2cwNOuMPm1Kf76RiIPD3OvJuBCDySSLTotcG5nz4EIR4xlJFgonICC9zYbDi
xeSNpUjAA0oFLAnUEDfQUnOK3gNRqCkN1acSQRNbZ2RrMKqdTjmbcW/dovPDMdxt
TGElvidLStKBGLFrGymlAn6/e7GDh6ChcFCf1Hj3ErychE+B8lizjyD2/0YAym5i
vKrbZaG6HxfOJQOagDqAcGG4A/GmqBbW9RpgNEMUOimL0yBiW2evsDh1bQQxMBCm
9V/WfUG+TZVLTnDRW00LnmhGGWkX+MyjJzxIwq/tdRhbH2pOqbeah9ofZ6qlhEJc
LIjKUNFATfDacr4xZI55BgK72JBBn2CnZRs9HIu4PwwmMXTRBJUL6JESLcOBKyoO
X5eaTwyuyr2NVuYftaF/SDiJzjMspsbTOIzNT/ot3Dp+xSaEK3DQQuWD7ZNSYqWY
lFGyPhS30IA29mYUcjKHVhy+fIx0u5S8Kuay5mqn0T2tjpSSufx13KsRFxF5y3mL
TuW7cwsH9lrq3XhixdXVNNquqUWH9pGpNj0g3/a8USEPj554y5S3sAOqomrdiHL/
rjGAjVfFM49B6J3BuTGlthXgFB3vnVuvj+58PNy6wGk/cwOtepjYPYFGR39Rv6n6
Tvd44uNeluNDc/kcGz+un8fvuy7dDaEkXkT2k5YvbMSTlSYA4QLWgybwO2sg4Gvv
VE+DsFwGWxLDDYM/aqbjpPZRXZqWyoS+Sz/opzNEqfEQ2MsSsbxct/XgkI7OYRXC
eP8jYlAGx9hE1N17AOBpQPQRcwL9ufawRqEG9dlXadVBQeMxRLachPCXfJ5fjo5h
tiSt7pfg6g9StN9C48TCo/KcziNe7R8aemkOLDZ7I4/nvbon4PrYaYbMtgRVc2D9
i/ciqh8ZWdFRJJklh161SLMq/TKrd9nicWO4QlKuxHh9DmpusUfkVYO4LBJxpOT2
7K1xmHV3kB51JaKJxVTLdvuYOiUeiL85yd2B7W4vKxw5pERt1t3hA9PWP2gC+HQf
VCBFlowUKwEvTGvfL7ULCppSMCludGGwniUcG3MyXKKGzviE0xT0yjrFbpTEydy2
QA0lJbBLVRcAJmFFB5HfDyf0KzqkpJFGewyXoR4SZQfh5B7lOeNFfI17Ix4jX49j
RUJo5MSTWdqflPOqU752NbhpwTkxSfJjb4XiqWVKzCDH6WS8nXuESWDBILOXp9C/
vUtz5AP/zLxYJGF5TWgh3EIAg0zt9C4uuHG+yBLy+6GWV/YUCTptMajsBnBTOAdM
Rwl8LUU62i87eP43pXaiplYt+LrDyD/RwGG4vY9EJoV6kS8XV6VCkm9bwBh9mqlJ
4CvjzguUXUmF0LJo7qpcdpAtj/1ncsuNHE9+g2ypBqwKNqG6qvbbY/fApynrH2sq
1ZtFewwvFFFog0n727SjEBxzfTSKCzXOYKIUjq8TC89FOgmUOJ0zUrNFwguJTHy0
duisvrdfusc54fLpnVkfkNjp7GjyOQ6FIxrdtAmO+H5smIZf2tDk1qsMIvrXMtTb
8rdsyBM9BIQhF+XWLiP2V+isK6sSqFt9bSEjtWqwaY/QUlcY5LrCfivXnwkHwkr4
lJvouDhML6mOkztZ4TkHwDEonKocdBASvqFnvOvGrj8GUxevMfJ+mBl92wjlNeDD
YjyrVLkNhOZZT9YFz+lJMADGVnFyYs1Hf/sARWHT90aEsQAJ66VvQR3/4p3++ynG
E0RgAFB4SmO+r33y9icYBedB9nCc5Vq3H/npFoLZOXVgekby+I+3fHRtr9XguydJ
DbdDiWNryUlp0xjchi0S3TurVD5JY/zJ888OGWhlWhX8Jx3SEcQKvrAelXCnPFKw
fV4nrap+ac0l5aSrKZK+uzNO2Fpp9F+3xbxR0RWgEJXnwklXGk0iMoOvPtKwcnZj
VW90WOvzbV3E+VllqQ1Rnh5nr16OQcyqm6pMW2rUkx2ECLhouCokv7ynFn8j5wgI
/EsJU3Fn0T+cV0i5Qz3hY265zMip2UvmMMM2xg+2WqmqPhKSrhAYQIeSft4/JF3T
x25wjeKq2m1G317LmBRn1bDRVlobZCIk7nHw2HOYzJ5bL7IopvlHNfAS58cEBwJe
aki/LSKUXc/glCfwtiVTIAkeD3zrvc8UyV3cDzMQ5hvsvTIoQHnTtWIevO7bj+Kh
xRzwfQaQ7RdgXdDB+KZn3w+0hDdQgq+Zlj9/+yeRlIo8TonTwz261H+LaR6rmgET
T15G8dQ29pqcXYoh352DbdPpsAsOxXZYKLtgGhBmfSWeuQN1Fcl3UMasM1n6P8n5
JugW5/OLMJ4ZwCxZmJzfXjijeY5b5JVuXUbPEEm3ilhHOu724odDPWKKmB+LdKQM
VoN/C1QRoPDKE9mZuN/zwWZUbcnFzQZabyHLaEbunhLt1dvfxMQJLpZlhYaxOahn
w9z3GgZGGAC4a2DLudrc1UyI1z1Otm2yRtvKY88brmCVPnhigG1pBtrJL2nMO+eS
93dtrvzsQRl7MxbxwmHP4ia01L/s0tAm95FBE/+BZYGo5zhRpFrOk4gzgC6YSNH6
Q+kkpTbgwoPSROBFJwKfiI3P2ZofbwPD6ds0GLurqfM71xKEppx+SW4d05m9TlTI
2dgyH0PjmE6xj/oo2nA/aXrBlDszfI1aRyhe35FMcR9klon30r2CzSAv8TGXfhQz
uAq0YrRusN1DVe3eg2H4f41t/wqKKAwjijaw5n4Ewu9IQwBCJaLAS9Q5Nsa6pycE
H7re0yM/NcnNcbwO4kwY9A==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
T/iqCmdmaObK8ibSw8gvL0PdRJ5MtxLCk2rVRMOWNU7JB8CmsGbXXo8oBAOrSF8A
w0zYjnjLSmJW01PcaY4L3pjUyzNQeuT1GQXl5+In1khH/bm3HIHprUIoiMBAyJve
TkXadmuKgSWJi0Br3osE3+1+Dmi6b6WJXjkdvcPhUgd4NKaB/MRaKBsOVHVZCvTY
wXoVqklN1o3TdWd56TKX1lqj6UROvtD0bYOKHuCQrUadruXW+GOw1SvifkitJ4uh
6ECPaLXkOGtwCuyRPNvlpISvHu7wBa4qaEscqrpHHwW928UCvk8YlygCpedcNI63
EzKkQwVab1lgFadRZFNeTg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4928 )
`pragma protect data_block
vfHwfZuUuA3BzTaNq7z+gAoE5gBdFZv0mHmQA7PRkC5ve/YHtDyHvqY+KlYGWysj
LEqRRRTVFmdVeXVVYTjXwS7qLEcvEZ0ZPxkdIMRe9TkJTiyxG/4MtGpK9YYPLfih
O7yzeVzRDuQGpxGlKtYR3mLYL+b6WlCYLzQ9v2uCqfg4ReLsrIZh9+1CdCvz8q9w
4Q4ucWLbgrP0bHdcxGGjWNtmRXUYyVB07BoW1OCSOsrcA+L+XvmJ+14cEpKqxCFX
F5kJ8Q/sqbUvC8KlF9aHL6rzgZd/ZtbmpOp+bfC+YbzT2sHYVKjtSOFLVzdVpuHJ
pKDwzm5AfV60+0S0e0PgASIqlUCL9DWbJDSl4GunkO56K7OZ2obKCJlE8Fw+5ZBr
t7opa7QrBUk4wJEatmf4F9dpcC7bjlyq75x+UE0VKQD3Xhp6yPG2vZp6WXCOEPXO
zannhYdepvji1eAAWiWztwV6SWTFuYO/pKBZoSyBzRXPmTko7B8rT5RgpyAAKdvn
rbItH5vRK21uux5/zTxEcJpLKsqvd+9kRTejxv7XZJcG+zsvnFKIQO3jb0OuI8uW
iRvdlxhzzsbNwExbjrkMbmtqP6B/3eGEFY5sex8TYEaA3Xeq2kGuq+PLUgitbg35
Q4dvTV0DmUKvpgPPhzIyCYJdJlzi7L+SLrYCJ8Roy7p4aKj2g6YUuBhh99zxMWTf
JECpInmgkbXw7F3Fpl2a/HaZJbaaYlmNAGaF+ymugJDa6K0GikUtbbV0DodFpGss
moPpT3ErSW8E7sKCNOyvYwvW9cB39scWMqLy+fWhRh5rLgwg+No3It9iDAZCKRNI
HRtivfpGk42Q7soFHkHKThIavevoou2eMIVGfZv0Gk0CY/rx4JsKtpttzX2sBT6d
KuxCJQ9m5bdANU+jVN1X+73N/VqcLXEzXswcx1KMyGYTOqEivwROWE96rN7JHW2K
Skjid+61jORZyGdz5MMweJ8PXBvReEwfqBZeUI0mAtECHsMFEB2DS6G3S9OGNsvx
M7XIqKdYoZwg1nLcTxFrvi+gqCKX9fd2Ep41gcqeqvpZHsgROTGAtAAvtdVSVg0E
rgxXDDUGrFlD7nu0M7WxC0Xhrbgd6aLMtdYIutp8npg9z2HkXESdBs98ccd+9CxX
Gd9T1TJuxQBpxaKSSpSOcJE1Wu+4qgVyGQsA/7OJaKPhT+xWy4C1OYvV5noAL0rA
p98YXdDVBXGTOgBm3nE/ewVPfaUlyOkuZVHESXGoEgHTSwTVCaPyJx3GI/ShC8Yf
L7TedKWsNsZpHdZLWkOaD8d+5zsDkF6AbGumu8UmMx1Fo9UPRsctP18eZ3WxP1bP
nTK6CzvCimTaTcJqZVKIXhmhLfjaHwpY7fbBHZNnlRXr6z4YuAM9HJ2Oiu0AQnNA
HpgnbdKZ/9o/fAoYa7KFiaRFjKZCb5CRQzYA8L8PPBZAYcPwjo5D6uWUmJsvHly2
8p4AbyRByVMCZ0pKN4jxEIZXjOogtZmtFteN2MZDL50YJSUlxB1vQzkeBSdWtcPQ
2Ri0LmF2B1iUP2iV24ypFJsNutRQFq2sJvUbFegCBQXf5BWePnDeYIbq+/spcJOn
+RC8UdV3ZqQuLZAdQMdLniecZb6H+Jovy+cKSVZ3KhMdVCKKqopqJzX3t2/P2vvU
cY/dAOXWR38AFRoqLK6Sf1LdE3cADgenWxqozdc3cTG57RaomzMp5kmJpe3IopL7
TPprD7rYxKtOSkrA1XPKQe+El4AbA3oP4v7x6xtU+xyGEbI7CaIgvheXET1WOd7M
sGhzg9xfevaGbP3vAxTLvXPuk+fxPrZSI3jK3LPiZMs36s1xlW043sF4S9nssIXT
tw9a41hD/sK6jGjovPZayq/YqmZgt5+Y38DfsGkJqc5bFI1O6J7kKIOTqwkOMyrD
nANuOpqheSAwS/f5qPdXv++8BOy5QEhkfia6zMpVhsw5M1utIsxihXU1rFSddJZM
f0w5dixyhd/XkqldJs6hTj3hzRF9FhsI/z1h5mqBbAkgoeQFSyrnbD939qhSMXIQ
zP6Yx3UrPzq0MVEZ3iJA/ZR/arHlVOK/WeWMvm1jbhITERDCumHYQihxPLSK9JeB
k0OTKELzIxf3JqU1sqqmzl/RQ1vQ6UctBVVfm/XVCBg9qhq5J/Yqx4Pp5NTz5Vau
YjEpfWNUkGyxBoH9OcvqazH37ot8WLm3UVEticutF0iPq+WJNf0mowVTpj+SBzOd
dQltGoQU+EevPJrbK9eqiKxFsnWf7rIgyNmGg4muPA586s2cnFki6lZmThkQ22Cd
NjZrLT3tMwUDi59vjOHfIsn9qoQIAw+3EoRX4l8ToN52+uv1BN/YojYr6oiylkWr
/V/bYbH3dlnJebL5a05GkcJ9AmMGDm4igJX2PKZERuf4NJQLtjit3rAyNxAzAEfE
0DIX2H7VPHUsPPFZxS1bcc028iqUO8lcDwLg5HLBBMnyxLFyu89kaIHlLDZcsTNq
YfTSZzvQihbouekWr4Wfn/1K7pLYxXxGbpO+/XhNs3tKl6Bn2ggWgD02jpsa7uXJ
DZpdxvrailuQYaf7kxF9B8o8y1rZUNhT143HkQO0pFflWT4SMyjPApSiA/q1dU0X
tk2PMKzCmmwizmagRRd0zIBKpc7tTw7pfbX7DWmaRPREdVjSCux/RVijnJmCIWrQ
fwlNCYkHdwv7AQ90UjWI+L7VjaKoBeGlZt03g9oFL3GyNG/6U4Hs9MEinA2bVSjL
/hgS0juhmvsO66AQpLwGEcXfH086YBPLF9vjic6yZjlPfHSmbnIXXXKWwRn+JK+i
8ZyLEYiNfELYtHJRehDPOOsgwhmFpC7XXETFBr3VFUVrnUKFgkh8zBY1KDnA7U3f
Zqjyl+lp28CxXdaiNCAz70DChokTCyurebKoKUL4PNdGPtT8weIhCXsizN1ceUUn
qxthPj39s6s02ktN2fHVPx5abEf3Gkj/e8NXgyUuvyfcA7MuGc9uD34H6IvS3zcN
xqwjHO+PI3v+bNbO+Ka+rnNn5PErDSV0HJn1Ne1SzhK8jYY9n4Hs+3gGr/zV90zm
JLER+Kdik3kf7PC4VQ2DOxcDPWBzrblISb+pnvS+tDsr2wAdEmLUTR3QJOCaHvPZ
VnQsHYf1tTJxZjJGFBG3c/QlsSf3TH1azHzapVtBBBs8yryZh9/PYXCDoSHDawMc
91365zU6tH0wgxpQSclBkxkDbUforfctewAMUuKERsM2kIiFSOHGr5VwnpcUdb0i
GvYfrKx6JtzuNO3z2jZvgNm/Ov9UQwyJmqdMkhKCgSYOWNn14sFLTGR/Z6I8Wxfu
/cpXKsB5PAtHKTJ2UpYA8SuPuQOwAjfaj5ijvsUmkrXcxhLP3jUBpcFuHLHTplUF
gCPvEWRyLVuWIFpeddD8P9L0UTBBMN0WZpArGH8QhhYvSiz+ptrWID+GKeFuN/wf
3GQ+/3OPc1QfcPn+wezSwcAZQ2ThMM9Fz6AIpgGm8nZXJa9HZNjtHH3xesD58WNs
Y7hia9Wv5qq0ZQOObj1BNy1iisH/PrkJ20T2drFqxQmNYPqacUIzL+3ZaUrINJd6
zv90oqjsz5OGYRLTNOiM7AdlNSpOa9mQC3uJJDoajZlIRG3PrRmAtQEIPOYCulfz
hm45UMJ8HVKLC21LO47I9dh9e4mxyrjQUrCtHRx+0xHi0DsaZy5tL8WamYV+UqGl
LYSxzdXsYd0RBLYQgYRp4cp4ul5u6V0iKZwvfrhsOWTh56RpuEL+4CxwUPil8Pfw
+igpNuHrVWtg8zZzwt0h9Sfqb7s8BRwpKzi/b1iGxHyWiYScgaELG5sdSbSaeR6J
MLCwcQaoWaoWwK07li1xbqbyqtVzWlkHWzkwxjXQdtLgn5CKIw/UP4I74MvwlalM
66+78hGgUXrvKCEk2qhZBjUWYSAqekwSrGoSKiqNuUNsmHqOuU4KePVM5EWgZN0K
W7tV5Mu22K7OgUAnyRVsNt3dKD9GUMZCyLgJ6oSKe65h4iuxRo9nyHBEfoqPUdvm
sME29a3zTp/gUhT1q8xg2vgJ9J9zO7ImhZnrnfNrHQCt09KbIpnRW8MCUN0qoU0/
jzxqrq7mg5lm+AAy3qJ1qSzbjv365+q99cQH45JBcnDagCJwH0H7XVhPaywfe77o
ysYmdCo+G1PC5oSjQ4ocG4yWAZW++WhTkGu33otUpxSlKOZeGGQ4x7iV0HrQv/D1
RDGINwJmCTeCF+afmW+6FAaaOW0FEzSt1GvxhY+S988n4c8Li8aIRNPPSwlU88Sf
Jw8W+93cb5b7vUFpA7PbQHUcBpI8W0qxth1CNWE/oFIq0ipnYhJbCDKuV5sGROw/
zjHCvCFaozH+ATpsF3ZDmneigo/WTwGj7w5Uj6BQTTeSDhZm4Y8LuiJ0BbbAtvtx
jhBlG/rF0XL+wGkEtzysFBZaFuaFTE22JQ+gaK3f5BdtFuej9EbOszgmejLMswNh
dxtY0JL+DKoo52f6BtkZMZzsxkV21n4V2A9znOFRZ2Ia/Juk0HL8SdUrC53dKYOZ
xLSyE+uD/tnftW01FgwGkenoQveJnVHQfxmFEPtZSfXC5LzJpGP4WBVUfAaVBd8r
z1/b/QJAl481YKwu7eHHtF1DbpnsqLbFLJX05ja+FL1zMksfZdik2dWpObG9rE6M
3qdpwEFmjJEK5Wdr+3gTzuWMc2Y+hJzQ+95oo52wiuDawlZvyuUSsRqPZSjQF8CQ
62FJQ1VbFs4zk49cSduQlJQxhaosgQ35d+Duwt2I5oSzDJyDzU60wA2+7pFqE0Td
nV33pNopfwfWoPL5FC9dh1uleHQIGubckn72QtXvpvKhOplsUbo6OoAQrp9b+6IZ
zN39Bx9YkSqqsPLJyZ1lyFmLKZ6bkZQO93ijuFwEfSPnHAj4FjjJNGivVW24h2IK
JntaKnz8QNgQWu9b4lOmSYQPFdZPhVn2R2L5nHrkfxHFtIqvAcAAsViKZCqZqKxF
zEhEeFGpKfS+FQaQBdkPp9xOBB0ZuZ7Zm/vbP3SBiqoF9Qo9o7L01Kopk6Gz6HH/
VgpjYQO+Sg57NJk9UlmR61Aj6qREuO/iWZX+fWPBL6w9kg1NKYmCoguMnUcTv7qt
0SHC+7Dhbqjyk1b33DLQJuty9fVvB9yZ8jPGKEBjoFF+jgl2CNumA/UzFyra0GIV
WOXTP4qnGNoMEnYXXNHuJWmVYWeA1ONjTjZvDctNOPaX+3X1JlZSmyqz14AWoGqj
aAVUl4dLIuzG4PRANllgZeLJP4FZZcoCj53ewIJQkxQgcxsGUbc8AT11Kb+KDRBV
ftskKHSVlMx/cESjvnkEbJD5GOBdwfRHko5WW4xcOwxk2RTAa2ThSI/v+tLJtrxg
Gxs9u1+EDJQzY224PkCy0IbiGvaXM8t6BOi0pDe0heKTAPwliDOoKVsKH0ifzsOW
ILXaNvY2mXwBEBxm/ceppCGXpr/MfxD9koyR0o5Y93qMG635qAaiSMytClAXiCIB
P3AuMMofMQda8EuPVAZJiw/y1W3GrPxgSsNv2Ws1sy82nSaUq92/wuSDnC+VPpHv
D84drdyvzpmcHm+bwHuKZw/hwBtI27spwjrjAEQKkjrQy13RBHRDY6P4ZS7k/iS5
UryImrCoBzk9uS69rK4qom9vFZ3fcuhhXk3fZ1pC6Ru2WxVf1MupK/Ahs/i8t/1S
t0sdhGKcnhk+bMwwbuKbJc44YMHXA1QHbqXd1AINEYAwKfpFyxxJVZawQ/iZaO2X
dUJ3/DC0Q5IQoggHecBphu5Vvo+Fmp1Kmjao8bKpwYZggnVDE9gBIw9+NVt7iDvd
8yIdGOaRuaWEy5RfYCnZve5/vbIouTvW03VSu0WebinCtSUNIxAV2GkmAXx0Ad2d
wFQzkdEIgQpGcdQBUXnT1PtzAiVcgWVs4ovbi2O1fzDyZjWHmGFK8s2J9BNFkL8/
fyibliYv8PVjx5dH+0+qC9GJUeRbZBbVZDbFXJrzc+8nTgNstrekeHh8C20t/ZDy
ZTy1FkltUA3Oh71Gat7SZmubpLJfRhaRoewN9jRJNZMg/cnRQph3nokYEH4Wgawi
mgZwad9P+M6vmD/E4qs3DfKQ24cqRYnThS3W2U+8PzOT9aFj3iEiJ30pIE5ixJYN
D394TcgMnZZdG3mvM2PuT+29WDYlCd7P404zMHi7JLk20Ty32Fbr+5cOkOA9Qe9U
S+GP+IzWAUJoOyxw0KrV1B2yjKwV4yKr2U69aKcEwIG7U1zu5mSYXns1ER258+I/
RY702iFnum5pknFmnhSePLlVS/IUZnl8vroBIL5kjylHIOrM92w5pwpkJkc2hTeO
J3Fp4MExmpQkknUjhpLy4ClTlTmuxkWPvTA790pT8Y407qBhQ5vOtD10oLdo1m6p
HrdZTUw//QHSk0OkRfM7SYGPrha467Zat2hb9QBKgRXDSuXGo2muLrCoaPzx6T0O
T7rcV3c3/Ny8z7z70C1K6CO805IuxhxHW9HzMEkBqIx56HHvDe69JvClAnMPk5TH
COvMoc1z6r6hk7v/544FNiJupBStp+zIhHJDtj9egJs=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
mvdF8lbv+v3UoHuWhzFwopJAX11X9+W5EMFXpWM3YalPrjsuw7IjBlWAQZiBu5hw
iccVnsrS6MzuOA+A18H4wAWeyHkm4fNH/NHQGd1UXJD3VN1XTE6BDUAySJlAaWSu
kbbDBfQHdCjD0buJYiapv0uZkkyNxlvtDKXvhmDn7svXt764PR+GhIYpxXAeW7uN
iZvKVzTr44PaZzAWxMMH5ACyco53LTYjJhn5ZKy4un1/bvjhMserRItTR0cWXxCb
J4rh21+mDzbs4uA746Ey08ZDqJRhzzZTLCcQgi6ZJWt0F39bviRDZqaKfMhCNkd9
E0SPVkXHeS5ypIqJ55ScRA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9792 )
`pragma protect data_block
ZG8RlIPnfVBk1vryf/9PwY3z6kvTcIwtlCnRXzpqFvHraWQ4l0Psmc9SSsp/Ay7G
gILgQcneYUZXnhfPPX9lna+QLkXU6pA2S7EZkN4cBGAoRDd4GXQQ2qFLSmXxus+2
ryjOcQI7Y1iX2BSNCtoQJbauUFDBI5CKJuTcM+70EY5VceD9fJKjanoJ7E+dB2LI
2kThM/5ZYiGf0C1Co86dAt8TZtis4owUxW3SC2nSVQCVjbal49xBNLXB0qOkgOK/
xk2HFfcdQUUOcRtjDiDX6q0pYCJrqJXmNQgRcTm4/IufL8Vzh0W3v6lbJ4CQIuG4
TI2r/R9q7lOuKvcqpI1rLyRh8W64edR+Yd+O2DPpJD1F49ylwy10Xv56AvI2Gc/s
gGBpYdbkBG1qZV01fKHjThcuyOVXMCldV54YkLUZoIKa8E013oFR1E2ypkGjl3LS
FghQ1mMfX4Fvsz308vlJDooifJsu+ghH8yw/KMgKCC9Kry0u5UnERqwSCTau3j33
+Fb0OM0hL40FXWsL9ZOhSyKsE2vgIoP98D/bTJX0BhZDfjSKxKmqQA4qd+8efk2l
MdwOEOx3XM3FqhCI9CnJoByPKhg5iIAoazN84Z6CQkShA2WWM+AfTWY27/mFEA5S
v/tJp5BGiFy0UCWEDA248/4MsRmhqLRN53s6kav7pqPSHpQGM0IbdErtr7aRHgUQ
Udi5M1OMssIu2srLQjRX0ckHBhnZNR/x1e2ipei7Aj9ho1VH9oV5rxa/C+UlhMxg
a3/ohcW+xslJX1a4NWFrdMeXJXY6vQcwMCx89C7SAidvbLXWokc0e4fYFpuvzwnt
pbjqRMK+GIT46E4O3pH5Ib3263AQvdQay77pb3KFYNr71qyGUstJfE/FhbFRzjCc
m78dxMDFarJG7R1yXc/9j2H7toJeAKOylP68IRDOR7eCNSMMYKfIuletYZxbu+gi
wiJgsPgeIq2pZ+7VTTaHltzfwsAA3niqjjtzl9T5GHcnIR60ZXvAXlX9F0fM/PJq
10Dfw+EpVSg8oizystkKhgBp5S53l7ou3MrWTx1gs9dVROm9cB37j/TNoywjkqXL
0VAQt9+pZngclvjw/QHFW4W4EUmTEshI9igcckAqVqoH6C7LZW0hDndlbyLQv87d
J2teqdPeHYBxSvnrmxCX4UICCaoBothnn+udXJ+XDa2SYMQ7qQf+HFplS+IsZhXM
AIQI7C2x/kqKuUJVYP3EjdrnPEp+FTYz7gGm+a1dGanFHlrx4NntScjHOJ4zlG80
KATcFqRw0wdIvMfF95GATYf6SeyRGlMadGPKwrZrkz+Pjlj0/X12SgFiRuIaoPrI
jYx/FrRnbD5zC3+fIPbU5pfcNlIpiUO+EvLcwBw07ySNHK2/odDCChmYU4wmtpQd
npmSKJ76E3ih4BCwT1Yexd5zFORbrHY3/SEae9hMgkUDvkIK79tDilaXP7x1ifW7
qNHk7uDC+q+SnN9XWLuLeiq6kmOFWazCBvclNfRj++jTnp9gF8aN0oSJp5jFczXh
xiILN3IItsPuzvPssRBQKK72stY8dlbiW13NO7OI/1N/MJCDTMwrcqUrw3JQmaoO
CgpH4wZtGv23erZbb7mSzMRwl55JCoFRPMUDkkCzNpxIeDoKR8s0A+e0wvkZ/roC
+KNmW2bL7u/xuadk6W6HrXntjRMmF8JAjBO1Cl0s6HktknXL3+W9Wrh+CIoxVDnd
epI1/wjZ5F7HpCZ5UFa8OoTRSen2fnRYxYdB3ZYG1tY3NggWiA2psa4qjuB2Kil7
x3szlYRy+MrW9Prl4YPAaeqR/NdRyJM4lzVbav7C+7mPPvrutqIdkFx3sVgEEPz5
s27qWQlstePjyUd7GAqSIJVmIyisK40zlWxhe7HN4nlRHUq9cxMIRFSAKIyOGZv6
zdYe8F5HqpyDQCFAWxqYyws/3GLrGdX3/lnEMak00G4+Xm1ngP2Dv3t06jaGnoGG
W/5hzxnVKh+XcV722yK7h+C/uWHH7mL0UpJQNmNzMIg4P++j4D7apojeJbxmc9t4
9TFomQ4mEuYu/FkwbakVvi2kxRnQvZxOSsl2Hb+C32bud2KgLe25BWyVrMRm/wF9
UBwf7v+Ce9azcwqoSJFQye3cPFUKAkWVwCDa9GBB9rBvwQCxBoXlPDvmRuUIYKBo
rg+BrqNAgHxoOh/TOupHIQ1zxlIgnTNPCdLI6/kuBm4HrU8tlLx3isJ8YYUUCgZx
OvCpx2tw1zpPd9uZDAf9WFXCER9L7n/LzUFT2vCxfn9X8Bl6IvStmD+y36m2+upA
ubzvyK8kTEtaRk+UdoziqM8L+qsa2pkL4/Xy/yWTTdB47GfRyqqM+j+7u7t8idD3
z5prmmRd5MgFFc8fdIqVae8WO8Rv7YnIhEMrHNoUmqrw3Fha7sEErCFSS2KvMSg5
pMh187rUiRDJ3sqUeV3a5kRpgt7NUWZK6JkzaJCCewn5sWTeYdHIeMEa2Wddwvo7
Kfy/wufkmGXPGxgTaaS460JBXRV8956WmRkqR6AY4qjmnQZzKNfkSdbPwgni8jLm
rXC8duDIrWpNkxsS00arTP3B8rnQElj+ybk/MgqrhrgZIg+CefBfAlgx4fkKp/nk
mp83Mf2N+xeJ2Mer6bHQmMQwfSg9AXIRdyHCDHejbYZN9rTn60qbZ89ot2Zno4N8
dUZVG9kBLJDceYssXmEhc6/hkThQflJ5/1pBxBsdJVr8c2sVaVN1cXm9j0GwitNn
z+USIx+cWATkFNNopc7aO3njju6JeVRAgBXfLZRIjrafm+iyvY+LXvRjLPe/ui4O
OWWgVyVW/7K8HuIzVOHrgOPrTclIUjf2tqhXbm5YgRbQP4I29hD6CFkPFU8gl+vr
JKlIWkl6iaZOQcVHYYNmRA5jCndNNPoIuxuPrfA5uPhTv6wpuZow5Mu9PF0ZyxVD
r3d5QNLP16PSujJjpk9xavpBWRnD2GSRtQ2E4eAUvXfX8Ib3B5z7BB2wp1cEyNl0
QpFna0m2na6dO2AJow+3Dk2Js0n0p9I9EpUVqvMInfCtCEe4Pk2lTjirh9Vaiwg7
vZqeAQXwPdafyDPa7PhcewX9duEIZdyhkf/NEzOOsWNkwTKxyWn6q60+b6vLJlrt
eHm5N6xeD6X3PGypZd0/KryORIWUDVO9lEXlPw/jh2nTwiDnRkEIPdRt2i9zYnfs
T5pNLx/dsYH0nJQA4QHAdXS7SxpCuTQ5a0tEMUOrMm4mlRRJnew4LAVLEhicqyjm
NG0xbHzylxkEusqyJBMsat4wZNKe+T0nNVqbekTlgxOF8jM6IlPkSwJ1IGbFsmos
lQabnwNt+gNthSPfY58pcF4ZMa4hwGKS08ykc4JDHtUUPQ137TAWXSTT0ED9bBHZ
sBxIhkc9HLjeQUNjyV8YkOA6qgO9p/cgIOeuxwwFIjuMXDuaM7CWVvaFVW6BjERZ
uv2zEqkwSdkbkYDUDl8VOY5aEDW3DYaSfzkRcBM04mSus8rxARYttgHfUeO0cMiV
9J0W/VSPGc0iZp38sGYau2IAYyfPZVp/W+4NX2womWR6/KN5Bz+16wlrP23/4Fpz
TzV0Ypo7ovXXVXAEmLOcN2VIjrhYA2R+ncDI/LtaUzEHSjcDHy4jI1ZEE5iITrBm
rnVQDqKHY1MrWS28IMGmbzk/noiams60i+UQNL5f6scbDJuyz+PWZY7o8eQslzR5
8TiK6pXuC4Kep069X4xgloT/M3Wla0qzwjZeR8WpmaEltQ3q69kxQyGPvklNXP1r
2Ehpp7Qphu80GytFZ048n6yRD1/QimGURi4l9E34mgeV8vGuqtbzw+wj9en7GXCh
MkGPBlTZMKVu5NanQAJg8uRKM2SZTngKfTujuijHHCgx4CqV29VgVbPuNRqERglH
Z/ZFw0LGEoqk7vN04YJEQaUv/aaNtiu81wrq9EhQa+52YHGOq4FMWB/ZXzJSnUDg
pUmLCDSZaLn4aJh/vGb4h/Lx6Zq0w5hAGW+dULnm/PLhFXhjWT9x1sIiXKl0Xr9d
eFf4namNaUu0THqoVBtbRHaJ4gGONtD+XL757Q+6v3HW9dLmgr9edDIYQcly/yG9
UTQ/A4ZkdMP9+9v2Sa5ykLt6if6EY669j5h8v4a+VxwNbUkIdzGuUdRTnePNwbNu
hN0KXBJnVcEBLs2ytQS+6y0A9A9VIf25t+fWi5NkZRXPEOkDLed9B8D5NiWU3H41
w3X2ZiUFVLAzPELQTVWYy8cNYOn6vaH8SI2UojvTvUv6xgmY+fwQU9ExgjGRiBn3
h8P/oa8YLsTS6rTgengF0IhlsyI+ZeVOSQoufMzqJG1lWkFa6b0iW0vKOzeDR69/
41zcuQfstFHd/fe64zLUV8OzXPSRPVQriZR/hRoTmb30WH7wgzDj2db5puW8gAWA
yf5eTSdZHE9WsifISxjbJbt4k6xPt4LE9BcJJ7wTVLjfbm1OXeqoNBK7vafzD6GD
bstCHaFfvwZKQZqCJgw32XBTfQSkV5KnYjWKgmPs1P0QR4m1q3VoxZWx0vWKcP3Y
JEuTNcgiqlX5PuAacCEpB4lPQWt/J5qxO2E75g6TITjnZrzxLo2oD5Olhyw3slGB
LP1jfXc7N/4n+xUhbbQZp/WoAcQzmgIzj25peh75+/tRhaizXF/NSd2vRJlc6ZhP
jwn5G77MmcGpxrrvvgUreEjaVgxerdxhVJOw1y/cOAUCQ4e3W1FYhtALhwKKeOCV
xi7LA9Wl3dQ1moKHOz8Rc74hxEmiLJAbYyAS6oSDSqmuh76yfcZowPb11M6puFuI
E3UZ8dzy2NMkmZ4DkfIoEHaoolc+6Y1QVi87ZMVB0RKcKj1w1INRU0DMGWg8Thrm
jaKyehgu4Tb7MiFsA0pJRZJVSf9iZJmHby7THDRvQc0r8M9RyAHbvNFqZHuywvVW
VnZKtIxuWbky8o6sxeQ7r/qqHemvqVsRfW6CjTAPDqiHaXfllSmWy4MBGjSgEUvE
nsO84Sf4+swxsUs4ZedI08b7G7scLNTGBuwZSSmgR35+xV56GIg5c7vAvhRuv4jd
vcM6fy7kzhV4bvW0aSkHlY9JCzkWOXdies/CiGAXQeTUmUrDrv16iPcZ3vmifqqe
eyEptMKCVd2siDRKVVBmjF6WEGJ+DaoM4g7iy0IA45hFYn7S00tKEQJ6TFLuYb1Z
DNgnIxzqkWRFfQocOS86YVJFU/GoaMIibHMicVLOQSIUq3ZbifBfHQQnxrFzJTb2
Scs6qvHVaoMdlfr2OVcD9gYkBgq620WsbNz3P0nX25uBz3CR1viQch0g2wL4hFWg
29dJQX6KWjfpBAXsUR9Hmux/xEGVaQEvN7GI06spxp4ykK8PzVYtxt359s4lwylA
6UWWnMYZpuKDUbYGuT7/6IvTLuEHfN2uimCPVrdHOGgylMntOTUFsHwPsO3Y7Eqf
Uew740f5/JMpTK4LqZuUmxbVXaNFuRyEGK36LzyGciPiuAZgHmGfjKeMcPHu7vEf
rcuN3Wn50056UzG1jrAKD5qbwUv9u6xZx4Y9hiNkz0628ncEoGsB3XfzlMgI1EXK
6qCUNduKSAy9xXMmGd6BHUaatXjvQ+MGOrnAaDQIwjFRp8Xokw84jvIqkgEf/UM+
L1lTGv6cHZJrbqSJ2+sr44YIIhhPslyI85nqPpdZm+NcDqLchRpW0qDjK8bvwOnO
6f0Bs7wpdwBmi9TPBghJOf1m7Jmb/Xzsbn1cXV70HqcmVCdPhb88mf+qjHvsk4CE
7TFK39FYZ+bnMEmKC5/V+OPIjd9PvUnlWRkYHzzJdjtyjOTzaix93ped2/z7E9aB
rE7ZY/YulXOD03U4Yq2X9CzpydDDIHP3LTaj+db2N1vBY0imhSXGyCUYk5O4ZvGW
TBYxBRJz6AJYZzZjb+KwBaYW7KN+pmPk8VgO2PnKEP5w3WIrNbhWcD/ZkbeGRSpj
jQbBYt6ty8JfUXN/9EoGY1hXeFqLqVc5TnG6hxcoJ0CJQjoMuJdB7mm1hUf07SXz
YRSftKFm4xml1kamTjjUD8mf4wpM4ZR2xCcoS0KE1B8RXyTxeqSB0XGaSklNKPvI
o/6CJEQPP+Kurt8Y4BdSkx8fe1M6Q1yiS1uIa6WRViPWD77Ge0q7+LcwHxCzsV1V
DK5ROEV1dG9N5X7GJME3EuT4w4/M9cGfXhrxUXoJcT7Z0neW64oaojKqV/hdjERr
DN4/Ydj+HHUtIeaS1w+MkWNxq3k0eIIxRTMxwHee8IWOE3Fmg6zFGJJBMAw33nUb
PX/3jB98naiL6ltetwxNf1OgL1yN5Z34uME3u0n/AsN9ufL+Wu6JcXy/cs+j8ycE
nR6L9ZeJPro2QAHsFvzYWFu2lrHLoxjnTAjy8S8aDZDT8vhK1XnXE1/fxm249dmD
Qa9OnYwCFFm3l8Fv5Ivsw0yvslhMKZfI0LTpTzahuTwfOPBfGmVFoIVZ4TWoxP9y
xg1xwUtLS3puoLcKOG20rIY3fhbgUkgCgUpuf1Pl0zbTVVIXoBNFMDgA9umwQzoq
BtANZYE42773aynWoRHWkH3K6ZNK2Y26MWAk4udPRvbsOBYVH2jOQnFAT72B/wia
cScAFVJ16H59ioL8SXC81FY+Lm9E6v6t2rKZn+MZcB0YMvCcHd/RDU2qj4rRVPRJ
6Ooqpeaw53vHf+QyS5UomzsFYCocs4sXDBRqcyNF1UQCBKQGtMQ0iT4q2xR1EcKF
+tzPxaABwY5xFZIlBJXogVldbrIhgG8PbfAPhx5sNyFvbx3fJaWjCy4l8aCzPE/b
S5a9LENpr3AfsQUBj52YbVpz2bCLWn1cL/aNd/HC4YstgKo/7iLZasixvQm7NUEr
N6RT2RY/SPBIeJJvg+WfMaSfJtV0j8JUrBadNNagd+1QFJ1iYmarQdsjfPAlgqnp
j/Rzbe5Ua/hQYe8cRDI8kfdCh/Pwn07XDmT5M/E0JY4Q9GXEWWgtSfCcTiwDYekr
U8e7fhXyTZiBiaYkEOgyww0Md1Ng7wmG0k4R7nm6KPuU/86RXcEBIQrE9IJ4tFJY
yodOoSPsQP3iiczFRi7ONNNU+5wHe07dobT3xdGLsbQ+T1265AiV/4WfjFn1fZPF
VYWaXWHFN/uWQcce10/spwiJIjdbV/Ch6lPnhCLqbhMV3jP0mbamaRbhz3SdWR40
vNJfcqOhpZafIle5gDCVqUSjIKcrOorGak9T66qPHWVfnZKj5vIEkuuJFP4n6dNv
+9eN9APQ3f+RHDN/1GgKI5gnlMvuTFXZZs+6MMGsbC7z2VuW1BeN6S6YcEtjURq9
spjvDXgxAcCEIRMk+LkpwvdoOvakiDEp+oGAcD40s5rizEmWpqaAt21uynJ4nANN
MAQ4Kd+Y56fkWzB09XfLvHSNNPoaXYyseqXKdbcDjFloKQDp0RIH6/oc+CkTVosO
LQGPx+VfuOAelU9+XHEIBdcXhKmYvvK0FNTjTJl1E54PTV6sniy0NXvCXZgotLKo
nrF9ogtV26sHas2hZQP2jE/dhL1hGH7MO/bXaJ26QeRdBo/AO8M7qMuT4yR/SaLy
wLRL6S0wKQb4Ya0u151TTshPv0Hd75H+hfw2edqay4PM0je4grhyw5bU4IpcsULK
Y3+ila7BfCeNzHNDLz5yDdyzIJhZHzySaOYkKvKiyWOLp8T1yGamJ5f860vQQxCU
S516Q6+eKIg3ihLwxeaieSq7u0E+He/nmf/KTAv6LAju45trQecZgoEVvi/V4Ush
LFvYdbAOEjOzt5ROZZZa6WCRPUoT2Z3h4m/qVICaJ6E3VwT+GET7XF3pjWBe7vYc
vcdkxipRmJkhpL9uVT/fkXv9IWsgkMvAo52P6rG0sJEgXeix5JeFB0JYv88cCSrC
H3acBryclM5u6nfqr44qX76ae8zZfRvXlPKalR2RRCs9R6rxSCcokmznlZvOvgJr
Oim5huGN2W11haiaays9V3OeJP3BeSpe2M5UW7aRPj3nhPqL3Doxub6pYyxPWvzL
KR8EuvxnA6VzIV5aHp/7OKWosC/ZDQ+oVsidD09v6HisDla5wWhV/u6C+fslFl6L
cau1JuqXtMFb+oGsOrN/jRHe8hMa4ys+6J2m+1NM78ZkhUbwkUO29qhlQdFEVYk3
ZIBRhsy92PSJefyWFBnPoe6kw0CHYFDl5wLA4OBInVCKrSxAZq34WdxTWrAPWJmT
j/aw6UurstqKh1A15FlT8WqcFq89fuaQn4XWLiCj0U6GFyhcO9OeLw9PBl7lETrX
yVTDLL2yGl4r/62p5ppmkD4RZ40YHG7GECE9wgrNwAr5ph3fjPirGdzAuS6vogib
zLyBXZ83yJj3SRErJcDjzuvojV2mMUUdePOxWw9T/MRF5pmnZb+t+bG24XMutLb7
4xYrB5bail7zWjUbCfAYY1EKVPofT6tAxideMcUdZU0lyQqRl/k4H6a/A/fOMRSF
WQmwgQ8Ifh00J7q8jb2BEFJMRhHaU92a06nm/w6AHNpBVL7qoRDjSoOtGz96wKeB
bzHiKYvJQG5IFmc3QXGm4azD07H669IGTISB1Eips+XFDjU2eU3hWPpvvurPCG8N
unsExPQhDLbnBBjdIw6Ukgz2SGnhB5QW7wQO7xMU8Xkt+MXJ7PqgC7kMepS83h1Y
gcx/8pr+QHEDH04CsS/ftMgebiprv0liSztr/w36vo+o0aHzpTuGxEMPK35VTsSN
sIlawykFga6+mlMCOuY1hW1TZxuPtioDanAaK7XfBLWID02Wp0ffL4tXJZdFJQez
POqa0/dmvJaMIXtJuOaWvVvpgrPJahEdC6ZRxyMp06YQ0aDUOlsCEiS9t8QUMmMP
2nqvXpFYxStnt74wx7CvkRDFqwLFjUkNSDMsmPBajcNZY/lT6QW0abfK9spwGkAP
9yarNIEqXwFtSdhqEKi8p0IljknjB91+Y/6Zy1DrZjBqz1HMCdHKhtUGEAq0JzkB
YMq6BNAr1JeDVuHeXRB5/IeOayH4GyZQO47A0DF83nfTsZ0GNR+qPXgmwmkWSb0X
WRPYTVN1MXulhkGe0wXj6iwUzG44pYZI1OvQb+Kl82K4xlf4PlweKrpG/fSKYVtd
WuK3Y8LcwTxrhlTopw+rcHdfOTFJbptWFz6SDSaspD9Gq8PAaGFCgeCPdONaXaNl
/T1S83OTTqoRKVcGu/XFJIlmlBgSySi1k+eQiPkuoUMRLKhi/UrGtrm7I37iEqwy
tSlseirRFep5AjHnZ4BkmDHm4ejCTbAMAhTiRtPUFkCWqias4rZgC8FXbVm6WjR1
w/UZbxOn/PAd157qZ3UOCZpbSjD+eCevBQGeEGpa4vICLIWI3XDQTmksCEsPP3aF
HzuzIQB8rziy2sMUEH+E4brSv0JBeJHMZNudX7D9njNiN+FPJGO9AK6hY6ttHzqN
DwvQcWL52MgvYZs79gCL7oxrzOIVTjM3v5m1677SHkvvXhd1Ppd+/F4/tS1G1eOj
g0RLQw84juXddoUTY273ye7HDRAojdn11AgfSG0qLHHsZkQi9DAPSvi9DHwJRMI3
X4b/ZyNYqDK7K2sLsPPnX8ghS1PqgKlI9vHt3psWUQvoN8a5oMVw40vY1ZNxj2s2
s/rwggEjaYZm8WqNU23dlr87UqgmhLYFsGscmjVF4LJdVjvK0/qbyRb7BC7JqHNs
Ao1AQFFTl7LoE8/CNvOb4fHRx6fF3sscUajUQBRtlmH5wpVvWasi/yPrk3Jw1R3s
mMD6rtX9GPpT706RY6NBoR7PdXP2m9Nq3qRVb64mtkH+eYwO5ao97QjXkiSxwZVu
vjzdqcg6zsBQuKax3xBRhoYC4DjW9dmNeQpOwD2iXU2SZjZZO/hjSC+7qF5Jh10O
BnVbvSKergR7JlP8ayqb4zR20SSVvbzHA0L6bTzTbLoqnS2MyDIcscGb6IpE+RJa
kwqBIwqSwxqkIM+473hWGNw8rRRdQkMorfo0PQpsj3LqaqeZXCj3ATzGsbsesTtz
PjepeBPNQbObQbSKsu/gNsDnCds95S2SIX2QeMUGRel1x1e32bMAYhVsr82rpx1c
w03P9JJwL9rZd5R9H6nm4+5V9hcGwf1SeWtNfled6sOJ+cZQX+eX9cH10PlDAZXS
EHqaVfbYj3tOiAw0lAwHna/Q+HfdzATeqk0iWMn8xqdAEw9CQUdxlREsc4TkHAJH
RQCbm6tMVyTdY8UXM4k34oMHU/2m5Qh9CyDln+HbuzHfQxHjiVUxgWitWBxWh8lk
1qpdvi3NjBbIlhJYTdhIcRy6LFbzDuUh6Ab2b6CEBlUW62zTByR2U3DWWnIZaG7Z
RHRSwcG7gEtsKj6Bhz+tp1Xjcf/nL528WhmaD/wlfMSQsWfeMvRpW45DrR8kia6g
EyMOL+Gf+5XhhRE9OGFhk/lxCMatvA6tOYm5Zf4wz2OHbJtYsPEYaGnXP4OTw9A3
F+Nsb9iN5ozkA0wTlfFKQeude/ppAMuxwBUB+mLhUg6KXR4Lb7o+l3TzmTOaf0yt
mT20S7gzFoiwHIO+amtZrV6qk6mw7qXr89tqHkNAeh1OP75RBhmvDdcO0Ruoy3y5
Fk2A21SZVgl5/NnnvLsHQozB27CLc0Bb2JgLQrzreFqC3BchUxfuJwWbEdPAal3p
okuW4FVCClXeHnu22AorUj4iMhLwY3OPfpxx1v9KAxYIMeU0FOU64nlAmacUTVya
mqgNrPwZIBPruhovuxhO20XtMHQQtvNo6+9wodTtti69ENGdB1gjGHNn99WTQ4oN
FiPDGYgSO6mHtdaDJsEFuqki8QRo14j6onP9Pue5Lt2qN4S0utzMFVa2wWYGPyOu
LwZuCch3++wxt+NTpZOpF0wEC1zA7QrVgSoE9hd+lWgpaOis0+fLRExl9ke0UX9W
+WfMmUdMh1p/KdReA47qMG/yDBirAVKXT9V+/mdGiNYdBmN64NNNBNc2mIayd+uK
xnKpmzlD7C8d1hvtIiqQT6iNg9qW902RHUHgjB7h+6ihkuJr/QrJtQUgoPJOBAd0
uXL9l1VwcuXDzd9gmRGx1r/pCaq+RJRYJQguWBXSe8b+baD+8vakh3FZnQwfoK2x
N/k2HjySeXaswIIgjT7RvFADycyHzXmxR9CliqC4YqILik3RMnTw/Z7jd8TJE9/4
t6Lh0cu/8+iyX7rOsZPHqbqemjNp3oveYvdfLYV8T33D4VNXBvGUiwFzWIwjaWTL
+weTKWsxSbx/+FXWWqN9PWVIbjAxegXMcomTVU3OoWCQgD2NbF3EGQAjkNzMDWNk
+tQDZSEADPaUSHJRj8PL1Nac0L5uDPx+RY1dWMjhEuucmEMwaybCmBEYtPzBkabE
kMl6YzryMwCE7oMyNtRA07RtfihI1ZQenDJTZ21+uBTN+pDVOIM9GRLXiBrAJpmE
n/aanJ9M4aTGCRyaQOgZ2x4eWmeVWomJ/bawTsvSRazRzTfMfg+Upa5HhUU/3VvW
bFfxtTwfunBnAEHyXQ0QO/BY/ZKyXeLLwAHa9138frZ+llK3moYj3lwz2LixHK6/
6gRZhHDaURP5+U05YoRwEpDLglYhpuNUx+SSyjf4WjeNbKbnwWVfNIYO0PXD0KBc
HkwqILutkxkjLduBhUPcqc6bFjGlM4vOrgwZt5cJGygO3EDHLH8IzEJeaGC6UA2C
XS5nNUCitcZ930ARDcbXnz9ZT3BayF3GG4kPWOy2k6V07g5jpAEYnqFwQ3y8acQb
I6/kCx44Z85Cd8lknlYOA1Nyln5iTgilN2mYBdmjY31Xy2tekmttWG3lGGmtBhf5
UCjYKIx/tkRudfmCIfzzQAuciQoCphFrhW/nmUd4e4Tq15jQlZHGDruXV9rl3gU8
cxrlh1DJub+azR9vHksx9TncW50GJJl68PSnnwBtjYDM4ogczUt7Zd33ZdIaplob
r5bO6Zo2vM6B51UgNiebv6qcFrzkfH5XVZWgojyz/q4gNUENVhm4ysCD42cKT/e4
2xiOKIS2M35xCSpsOqsD56zdwC4zqRio9Jb3T2ICis8lewcv9hh2iJtS2xX9fJbR
lUOI950BjJ05byJzPY3Nxxg9k/jYNULEy6WAi4yNF0AeL8QYkMhS+ijGQ5dYZPUT
UdZuHna9uS75vVlDulHSba78hQL3IMSfthC7GBqbow7upm0qdzkA3q839/kEElWN
IAXGQNasFuvgBwzk229JDaTxKfMGLjtGJm4ixEY/iCLgRK3Z2XGEwsNKytvzU2Pu
zvX73WHk0tAiWLRcL9s8qtjITJ83YolNBKgtZ1Ua2zyhc1ggJLCYG88rgk1W7kHb
FFtAPEV52OcGwu5gQLLkecS+AF6CAKjCyEwQNlD6Sl4wKqN4A19UfLbPUB/PuaDx
NJC0tX06G1jBCbRh7UuYImaQlsnMyIDep3LwWiNv2kn50T5H3wXCkTaDjMSll414
CHcm57s/JCLdYT69DvoZzCTgmId2OnUH/BK6RiR49R5mwtjpeEQlTyyqePtNMelQ
xT1BB2tbHa707UGMAjLO2GwFVMIOx3snOPBJyTRIBaiGP1N65DsH+IknKO+OWFmE
dLzjKS55S2qsWKLiYNDv85mFGtQZWFdqstRkoS4C08rk1HnW1PpVC32Txd+ezSHX
+Zh0trhMXIUPeZEHWYdZ6872USWGD+4dPzHLY3rKyBPDfXN0/JFcHTBnY8BMGIJE
eod+JHX7MN+6squ3Yps7/Yly64CBRHlRqczLCltOOSNAxSjd42aAzcQHP8SBKnlb
0a/+h3S7VVkk84wCYA3ecK5LqG9tPGyvt7jo5ETpL3ljqWNyNKPkenI8Iq5l/ZtO
fAGRDEsIZMYlhOihG6P9i3VMpIMuaHG0ViQAnzX08xUpN91ASZdFhoEPQN/qDcQU
2+IfItwPpodhxQgEFObyGqT9xiinUsdjxzGQ6Qid+jGS0Dn6AaEKEU1JFaQUWZpp
0KLhCFp+3RaCb2Vsrxtwi6VME54lKBf9okpA+6eMhSbLivSnRKrfUYyH+lwBoLrQ
Bw4IjLxUvxOpq2g3GHYo1kxaDOE4avyYMBdgqOM4eBopHCcGwhxsAsY4fNx9mX3e
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
i+8YeI8XhzCmWNi+vi69KzFDjKbpEhLiWQkAbFP4DsuILCCK5aKRrO2vZ40jyQvr
qdgFzF92+MMg493mEK5RCeZTwPnWDli4BauDNVi7ITBjAavTJ1A/fBUZOUhTY9Ui
f/STwdCpafvYIIzdjqPB1/FG5fBglwGhfWQ+PS4ZCJyMRzW+ZV0J+FK4qT5JjDYl
WYREOlwJFwVbFKlJJo0THKrCJ8is/VinrS3wN92LpMfEW7zh5f+WI1WIC+mM8+Q+
zezUvtWkTF0DiF5DkjhWpO+KKmlcAPndVUCh+vO2TjdQslgM5rM2cwIidwj8O+xK
JpGZkh7+GzQ40PAYm8WIjg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6256 )
`pragma protect data_block
ST7+vVp7HiTG1BuDR4uU3IgR4jefS0rigZdy/aNKf5v1vExcqXghpl2JBU0XLeLQ
uzddNJ5f8Ep6kHeN9fJwWvEuLBz1bhRRjRJUHtgAz+rIxjfpN9KRcebbdD6s0M/K
m8SkzlqzZ7aTqKHawGE9gxSIkNeaakKIw15oe7oyjdohq3wUcPT5dKIIHmgYvTyE
Rr7bK/6nUDgeIEFDl/tQjL7xXTRlPO7EfHvHO//06FkbCTOZUrkho559hqTXNY0a
oqc0h7NqzLXwJAE0uWJSo/Az56wf3XWj2KUpg+6qR4JyTndEKNfhXuZwbRQZSf8o
KAooNtipbtGNAI9R9GY9LFCQmd0S/E+Sc3bSPedevUJUvyAfAhb6982yutK1CSmh
2JVkGqvkyLuDshjpNNZqq2wvl1Fb4ctvfTIgW0zyar+p0A2JeuOa4u9ik2RgwFHA
m2tJS0naLBIqGICNqZypHY/0FF56bF6/kPThfjJgq0UcwYClkGCJSA+9VjWxROoQ
PhPdmgkD7H8cDimvDVbgSyFmMlpGfkhbQ9wXJHP895zpBJsn7NfrzDiSnHq7C0LL
NwfRuZees+nJ6175kAEdkOVfuMj8IMt4s8aZSrur4zXzB0G9AAUPEx6cN37Tz3tU
Uk1mBQksD3Rf2MLmo+Xn9Fpxt5JeAgJps82ReRUGtLP15v7gQcrWgUHvwhPDq4AS
59NX1Bcwj6jiYN9W+Bj5wVw+tFSb9q9DVRzjcSxm9PHIlNXvh3DaPb1Iz6ga+BWS
2MaHYyJyyAqRFZtz7kOSWKHP3ztvUyDA6vMySdk8hSJYr6xlD8gMmVtyr6N81CEX
nN7Qs8F8u2e9pWXDsuWtXgVa99G4HuXiVFKqH/7veiZu6rSpjMZRCKYEABKaTdSG
8HcCfHEAMCtvSado8gBmgIqZeezWfdarJ9chuebG1tI403s6j0AVzvJOYwF+vek+
gnWAoYcLt8hA7uueinCzOclO5MBiNzVPzi8zoO31iETvOJTLQMj3NLBSsJWzqTh3
kHD+flbzeW5xAJNu9HKZWIxYFkl9tA460tJmEy5UEynPXgIWHEMXe7/dn6Ax4hUa
wlC4xIIZjf3lOt6c7ceFAFa3sE1duhp5kuqhbGIOKPT5eFr4FIcLTlcIBvbl49EK
t4seugVCFW65MwUWnTXhK3wvMPRAL1LL/c7rNZ43I1DlxbYVQAwDJMVBfzRxdUmg
lgMjint5AGgCkyElcQ1VfJebSjm2rPN8O1Q2mms3Qt7lseER8h4Sr8UokBfVug+0
mBs9cLUW4+l302088+9txrqtd3bhDfAU6hxCGj6kAvX/G754O4OzXv7Q4KHkkOHa
WejyPf7mZwCvffCpKizp8DaemoL8Orp21rpbeF0w7ozkkXJTg2EsjD5OBdmJjWCM
TZloIdpZ8KQFTsVIATDGYM1/cCU33usiWDOWFGGrqwia6k+QH4R8oqV9Buqk+OMN
uUkdDrGdAd0qaTw/bA1fN53ahnrnqo46ORfjvrYTIs90/whUDmgDHnr3LbTPSzAp
YG/OSUvzq0MBMcXOLXmwvTJJ1aocTuNsZevAblTqBvGJ+xhGyV4PnD+lrwPXp/Vb
1lGbLTQtjDsGtmUlQuXf6nsgOrSLTqfAl3/D5uX6lgQqUEYw3e03gUV0gUcsc4Zo
pZFIrjS17BL1BQy5yC9xfYCt4G6MAaSk3HUYUh6rq9hLl74WW3MubYCpAnpX7oYZ
9dbLw/9M/+FFwyPcxXRCd7eOm1Eqs66/8qGXE4OIVfxLD1YZHkjgv7GIhs+Wco7c
5fM78SdAfj+D7LXWifAp+FJk6Sh4OeH7zvjd/6Dv1sOebSZeKjlL5tOIIkZd1eFw
2TUwlSHbf87M6N80r6lNCeaNRVK+QtXhaCDbS5tZ/Xn4xYyVfnOgnhtfs9Cu3LnE
HSkTd/WkPRBicK+qnkiELhqiv2LfCqxsoiEOCJjd+keTyMyRiKw0SzMxGNEWWY04
hCs3vfWQz0ZS8IU561aJ+TdO3B4pj0boi6M0w0T5H6pSqFxiFs9PO1X7yj3Jvmxu
jcpyOWiizOAkIKJqIFoyDkpGTsrDTogVELkeQpsQpvDawBRBPQUpQvSLlVoioEdr
cVwKmWHRfsPd4vXmKf6dMKisQiUGBvzqHPSK8JyWqqIUOm7UAglv+N29kpeg1/cK
fyjV+X53P39GRd4+wT3v0EVEQL6aUu6E73Ap07bbTEmlwDoEaUEsXHQAy06WrRuv
wOZkKvG79DKMdqe/BrygxGWMJ55vnj+Fv3EgdfglkOuarIz1DP1omxuvVZmCmS6b
7vmoUmgFXBVc58ceypt7knBG/ECrupjhSkXv+PAlar1kX2J+j5lVuSgLVuWcmTzW
5GvMOTRiLdyiIa3ClM36gBL2UUXSdBn9PmrU0BYQFQT0f7PdX71iKaYpB6zceQoO
C4tdpgJCgC2Kw+tIMJ32PFLzy6/h1M4qDErQdQI/aiFhAs7uxuOeqGFWuFOUqXR+
kRDth7kLAnqTJRHivmGb/yd38vMoExFM0tQS9zwyRU+2Wi9w5HGlhI4SnlzinOcs
gr54w5a/LFR0VYRQG9Tz4VXkyiHg9rPDjrQjQkgsFxFQCCuyRbxg9u2vnxpwm640
TVjxlSv/xtgV1YomU6jzweC4c85yir7EzU8Kh18LCi4feG8mHa6s1Gehl7Huxnwu
2021bAMAIfIPun0vppArjw99qKsAqfw7uZfE6qZUfzMdD2B2HAPsliuXEdzPGla5
Ozioz0VXnkXYtCXON3jg5hjvnZuxivQ9M4M/p3irGgXoM6uwHdqnCYGiSTBnbblj
EmSgHJ/aieJeyuWlyajfa1XPdYKHIj4bMtbcT0JQ/NQCr19XFeihpui+aWlS337G
XJccyZUUrzAMLDWKDCjhVEhGEdZLNhjyEah7SaJaz5Xk7XxNev0hGuvTvrOc2X+T
Qwfj5WojHHl7yR18XdiEK59VBX5T2xvuqYjdlDZ6npULa4hBi/rWwKRQC6XAqo4k
UviaEIjFkOLAGUOiyOi6uxiU2qmz3WAVmBf8vSSqCZqdRVrHykqidre0H6e1/yHj
Kjw23OxaHNSNXG110ZN6rKjEsNdCag7qF1zbaNhd+2rWTPrJ3swll0oqJJQL6EC3
Zzdp1aDyUK1FA9ygeuReJbxKinYAzKmteRj+FctGVFhFObqZEOqpueT2OEokZ41h
+l7/G0Fgv1NS5Ilxiw0npBgNikqSaZvXwsQgRy7SiyU1Vl1ZQARCzRiKBUlLOLmr
EV4GkctaxwNC0yfr8lK/7AoRNCY4gc6m4lPE6i5a/e3J2M8Gcsb9Nf6+/JjpG4KM
an4FtPtBTOgdivUzPUgk3NYU4Y4jx4E176pHvVvrb6qNmxeWqe8WShEgSsf4IyVP
Dkgoem194E4iYzmU/FIioBc/mqdaEcpPFRoEZVO/uHmg1BSGCgQk7d0epeQL8KQh
u2mz4FLRRaza6iA+XDvOWO+RKON8NlJuP/A6AuO3LE3Rhbuk8j/VXEbDuikbh9VM
IHhJNPN+P5H0VDuk5tRjrDp3MgjlsU0Zn32J69SXIfx719yaAM58ad9U+lEE53tC
T92s1kjHP4VycZy5C0IQyPPvNkHgzhnpbF6jFso6aPBZqDmVNHMLdMONpAri0I4x
F7DTTl1yzK338D27lcEtrMi6/GriSNzAL0b9GCcUvrS402N2KKph9UZbk1YNZmFV
GGxTS/P9ghun8zsUnno6nyK03lrxZekjHI0JT6hISMmjwIqQkVOWKpKhgklBm6ru
DgbiVeb0zseC3Ywhv/qNklvgAwuZc0sqByfPlSVRy98xKdyDBX5Nd2bwftXvW3fP
JB0orfPLgSyFGkpU1PSq5z2pjca2Uu2t+nC+0TRawekRUY/YDCyL3rD5vm8hb45O
Quq0drNqzyojPaW3cJCqD6JyqP13BDxIrM0ZY28iscVOZFHIjh9DGodHQa2LZstT
asDaCNd3ba574tes3FmDIBWEk1yL3R7mEhZv4iTYFPcuAyU02ub4FUOcO650bypr
0wOXtq+8MkCas1J68o1XOCyvl384PZruGECnU2iASQhY+HEcDcy9Vy0ESUa0LQBD
GPNkwtGcH7sFOJ6/bhi8wdoPslGbkqH9sU6U/U0OFHnz6uciKscqgxSI0iKIheAD
HXSarBZDqQSQyMlh+UQnS9uATwhEyAzHk3A8Md8XO0u9dx7ia3IN4ZA1xsSCUmE+
TU+fg9kBSCXoHG6mVjpx/+Y5gyGRRJ/qfSDGkVmuhwfJnQnwH+rV2faS+Krr33rA
q8RJwvzrwqdaUC5nKu+z3pJa4Y/F6/mG8P9+tXppxcBJ4PpDM6cEp+Z0OY8GL2jp
oJ0YAZ06VkDYwh+LjhS9ctolc+wfyuBkVnH4bZ9wtM+oAUvegbk5dY1XhEQMKL9y
nbhW/2SavSdBh9f+E2MPWYcyI/Vffr4r/nTNgyif8ZfZHzRLG7j+CbnTH3QUe1XN
KKMRuQdWl9lx6vO8ge4qaFsElJQyYuTYBrO8ryaUIh8T4tPziiLBg/W3UNlR0UcZ
PlEAtld0Bz6vKoKzelEwly3MbJdnAwQHtsGxkZ8aYIskQbKl18w+vck4zyzhY7/F
AlBlOtuLD3T70M93hTSxKblxxlC1qqQ6zNZAMMRUTZbHFIZL2u9UUKRhp7YTvvuT
kplZOvjRDEVnjMFVqae38czL2Pd/RnjGn4fWUytNFeKdVSxgdyQnfOaPv9gLUgqQ
+lr4ciKjKKhWnpFKxh5ndLCOkXsyUNqu3882M+mS0dsb3UdDX/e/LlOL07cxpWU/
F0hTn3bYi08bwuPCAMQUZTLtS8h2UiB9SsC4nWc1wzsVlz+PaaBPd0Og7pN+4n0d
Ur2S1C/cpUbPSyEDiGvB53VCmyAlcLyeeMwngKVE6sz+tHkfEkmuqHpFtM9PXOx8
NsuSw+7dZhLRa8g7+n71SzB5bYuY9omlbW56u9zqZmAY2ft2X30NMd5rWYerS8XE
JaQLneSPmG1IGxgpmodaSo6qIn7cD0VZJ7TTT2uWumr607oik734SAOF6e62WpTI
z9SUYwEhSEELDJoIPHeQnOLXjQINiIyS2DYKc8d4XKX8Veme4K4GtiIQ0yrHzGTC
dfhSCLJU5sxAjncA3jgIQTfSBUsJUE/v09dFDzsajuLW5H/HfAmhDtlushp1O0OM
NOdkYWrLVbQsi+5ZqCum4ZX50fgSxIHP1p4rhFzxYFtjmeQDuHv4jCK9JCI7OhV8
M2B/oVV8OkT1Bl5CaMT5aurIQqL3GmdoEHlKP2mVk6k7+e8J1yD5YItf6Cvywt+W
PAQaM3WqQzOJhxrXrUchygJXykyCephCmlr272evRvV04RwDHfJlnacVBr+rVh0d
LMSFv5a22ZmurNPh4qu6NtSnQ2X3o9wmOypOiRmfsuMkrPR+fvfDuQmDBS8Br1+B
8tFCjhI/tP9HLcuHp6HdrtwRSRSDvpSFizxPoMpjdDvtxq+VsFS+0qg44qz9B4Xg
f2EQxG9CcoSM8ZE7atVrZJR7h3Qu4yL5WIVj8cCotUIuy05qObXa9WbSPp49jVWi
adv7W3xgtigtAoVT+Y3712wKkVpD1P/qU6LPjhkM/dNaPqlrfqQ8iyiPgtZm6C79
WCEBwdfEcB0260ty/1c1TtmirkM9ULpWz7H6JYaX+Tk4X1PyNmfRnL51A1FMx2hM
FIpOOAPlDnIUvBpLdpuZ2QcRk07H1kk1xjagpUQMmH823OMTLgkuCYMV5l5eVXVw
dVT8VVHwlHYOXTmU5a+vgyj7q83L+TmO3UVMEZtHS6S+CXTh4AjQuNbp7z4ZptmB
0KeI27CAEHfrUzDslqtXlcSDmoKlD8TFWPwYhWAf3ydVgkxfq+LbGO7+mnw5UWq2
lCCFsODbDmGjt+NZCB3K3UH0IX4R/ANtKQ8OaK7n27yye8zixjYL5gHeSTpyrTlE
IoDK/SPSed6MoxGSA4QOG4NjPiM4WeVIHzvY5JhnJqau3rUlbkMjv/wRbfa9ieni
NjamGRSpSaNYI+D9jrdzvFPwKFOC+w8oaELQk96djf7mZc1Ka0XHMBgsI4JD/XwB
Hi/M8KcGbb9pGjibghug3mhJ85JuXZayicozSfPjc9Zg1Ql8LDygq8X1F/Jfx2LX
zme3a8+8Estbxy/qrsrXU3ia/Vv0qwSHP+e13Mg5dTnksBWVF+QQXIYiO2wXf3jv
2lf3SnV6z4mGfXMDlDgxID4EicILYHqAXYBSKfEP2Rz64Pr4k74ON5zpi1p+cojp
P5xdxa/4haaZFVTdp8J8LpQQVXEJT/MXbaxEnqWvzo26fQ2Vzr7Hd1wB8kyV+ki6
O/DewAdsjVvuU6XDd19ZywJfqSV5oqcf+aznjkFS6B/aCCHf1CxmOPENr6UfFkEa
PsqRexKMffYIc+hRtE1Pk364TT7CteVp7zuIR0x4mGQ4Hbhy1mZljOe0E2to2eQr
Z57Bwp3IWlZnooWRC7XRDmWgymd7IEZrPIfASSwaQ8FCkYBNFLrNcdDwgYdJEFhy
Kur5eydiXbUoyJgf1sp+SFzcPqLMMeFtg26MEqQd5HRhtl51Cw3s6PoWf2VCY4Z5
62hdiJI9OlnTwx58VPqtkqcHI2FQgvjPMGBG5V1u9xmEgdXtFkYOuLgT9tR0IWrv
TeieFTSXZ+yMWG/i/a8LLSHrokllJ33RhY0SK/pxuWe1Hp5atBZ2g4zJ3aTpuTJ9
D6jdKuTFgUsCNYfEuy838zP/LrUhl+0bmNEzeHuoHqTIvVBbFRtGh4DOQeJwWvo+
PE46yeXLJX/Gg07dT+/5lZmd+0GkcXx2kjY2clc+OZq8Py6m+PJShbUe4IdfvAsW
F3H9qW1KrqVOVxtvlHIvblPI0sPlE8D97KRaWF2PxHJgsx0naz7Xw3jgw8Xy/Ovc
f4jFntE0Yx1ekdQzUEnNG8A6xv0TtkAjcp+ks3gKjghihYb7azoZ1Dxdy/QNCulD
TMJlIElrWKqCZFKVldAr20AcUiMCwq7nFOnS0UFK9T2Ti/SNWoe7LRPusmJtEYCD
X//4tVt0MoIduDzGNT9A98Nz6V7n6owBng9CsjKoE2wbi5REFf1qbpe6U/b1uIX2
zSWST2L3J9ppaMQ/aoMSrkWq2KtPz/NoK7lU/wWpUl0Jt0jCfMKtWse9JBK/J6cn
+VFsEIsLY6EU/mC+/Ghfvp+uiEgHb+gMhDO9IMhbrK98XlvAIdjWLteeeWJ3trye
gF4UkxUFAXBZ/MfHTDCWm0GwEzfReJ6vAu/xwagGgeTXuEEOMkZDHql50tIAG4uk
78gsla+LPwdmXI0xqKAR0hqc77JrMJqjfejbLZXF2q5o3OCp/2W68JwcqrwmrH8Y
uwEQAKlgbjH0j8WFV1bZKRYJE3LTPjJEq4QJAhWivkwDpiOf0gxYeObn9TMXnCVk
Y/tevDnOp/Vt9d2OObw9fWjftFBMZqI5qgbaVr6gb/BIj6ZFAnwgby7welvhB1iw
6R2Zzbk7hbEB5zrQ6InGTacbCDJ2w4J8ja1fpWSo7KGKI3SGrDtlVXqnNi6tVn/u
HwH7D0kVJQ464fI89OoNPoIdxhf7RkwNpjDMWc335PfA2zUAF8ujDSBjkhvKHQRh
74CA7HmOZ1mbH4Z3f7BW3RIWkSBhl4khrPXDmn5HOVThTDlyws9ChS0Zo+qvi95J
OycY3MTQ8F94WGVTkzDBZtQ0M3jp+neiej6335NX2MKDmyzWFd/0uwKjByJ9lmnr
kM+WxkbUysyaGKIzL8Mk3zblVdnJU96dHcg8z4fvW8jMgb+H56oaA0E7HHBfXZsi
f9jkKMALBkX8GJLjntzpDPbggS/ZzdEsumdL+fw6YuiBwbDqbomiL+f/fw1+deVu
amUM9UbyRnVxN67p6zc4Q5xOp9oqiL9ubNYoK8LQ3YSZUtzR8fC88dkDrgO0fxRD
eAMol5X1swOLWTIfAPziZE6x8d4W0xk2WjTUy1Q9Pnnlko8tsLSB4xaKP07GT1Tt
GB/9hV8FjzvW2LOwA9kS4/bq29R39UgFv4d1ql5IFwbmvTu/19qGYftQmi9fvGzI
2dq1DDJ55CmYRPXYSYzM+QIp6JyFMpE0xlfZ/7bWIeIpKGUSDKO9qzfDvE8lO0V9
AhFaVd1/kiii975/qGSruO7QHmQ9Kb//qwU3tnCht3/anmORai0QGilRljfFv5m1
dJuYKScITRXybYVJO+Dq4HNhkYSB+LYjmEH5+WIdtg62/Tdty+lDmaAeN9/bCp6T
rlzo3kWB9zIIir39qdwtxttKi/ZppvgZOr5OpPwx6QVOo2G3RvyMB2jr4XFM0uSm
RYI7GW0BdQ3J/89kh5yS5w==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UOJXKMNu077SZPiQtogyhE/P7Pp/IfleEmpvUGb7NCUdfTE8fndL1RpGF0PdzA2U
ZYNaGqEppqFuV6Fo0eWfwvuW8/q0F31SlYl00xeGkFRWHgulMeK2OsZ/bfw61IZF
UUted4uDgVa0JbuEPw3GZ7fj68k36wNuBxjfCI6PFhvbUxArpABi8kGEOW1bT49+
g8fQSRomkUujrMpKam2G1vTtqFhp3AyPoZPeeQEGG1qSJkkAI8TXUt7ZYZh1HrQV
aNeP9HuS5sv7EFHpLqcYQ0hLboJ5dRlZ109CmVaRsZj3+Z+it+h2iZ1rehroyzAg
JYJTAK1WNYV+MmaaK8anyg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9456 )
`pragma protect data_block
xAk8gWxZLFguCqOJ+qg2QvlZD2K1unPycafaMrgXCZzaPU2W0pXnhB0pS76K7eBL
yuyup7NRrmW0/hbURHnCatLZFlpSG/9EHuMJuo4yPtI1kIBIvr3CNIfMe0QcoOXU
hvOd6xq2fSXsnMi2q2RE5tTi048Sid6v7eqZ1LRYkxO6bINuNr0lBtUcZly6LjLL
VbTYHV1SCPbFYSqZJ9pHOlYFug2fBjqDlBdAFrztpqJKV9F8JXodpKpBo2xjelwN
WqJJp/a17GaAoob9vS5P2F+5KpW6rGQm/dWHHprSqUanGNzEhQe4reqQOjCqvnKQ
+vbItY8iZtY1p+ptIhrkSrAwiW7ef1BPR8o2Mit+sfyO9FeS0LrV4jqXXc3vTWHS
4AF75XqblCjrknNG+wpju6ejR0PUtZ/vTjjBJHqyFsDw70EwDIcI54Dy6D7PK6st
qMfCINcfrauFNYVy2U4dVEysq6BYZ8dtcaMqwwtQdGuXI7mIbV57JeOrFEbGKJ7T
SAQjX1U2/ZzDXIUiqQMntHKihR6Z9oKzyttVh3+eDMDqYOdjANBkwe/it/ImTiEJ
IM/x9E38PtmIEpI80uJAwkY1ND4dLXoNiY/dW4TTBACkgW96LcG0jWUI7ZdxCeXe
6B8FXUFC7VGjxWSA8WF2hLsLZCArqQdyBUFqMTGjpa9a56UDwO93FMvK14k71vj4
CfwKreJys5hMNrZN9Sdk//JQIUpMlwzNbie9K1FQgYWerDFa2Ta5FdGXxtiLqTlp
MEii5fyctEfZLtjsHS1hAfa/89o2HRiEm4e5okNIjkOtfZtf+lSmJnfGU6s88DwS
2Kyu7Aki+K8PvmOD10GR7uBR2Zgq0cOP8gVLZLt75eqhg//iNrbAwS4tip508Y8F
5dxhv2qnNseBlTGkwB96XpHbS8mK1Uz1c1AFQET+gKGV7fkI7sWkxXyEDPAh7dPy
5RSrCdz+0wYoB83Ul6TTGu/Zt5wXvCJjbrqh/9H/UZREnEI7hmhkwDK3UalwZ3D8
WFYh0KtDp/oiGXcOfkSyqSqjRHA0/4OOUpehZQ76PfUwsGVTl3HbKVT31BHl7DAS
8C1U5uI0cWDSP43ZHXuUV365+tKgzKlgNC/ineErH3WdBiQ0t0AIsoX/30I+PQMS
UtL5Kqe/NBb5afiLePFhLNv34FjInwx7fZHBfaSZwcfdGGzhwm6fOfX1ye7Ev29d
Gb9c+sEQP66LgzcU1vONSpCkL1MhAb+aiXGnsTZCyWrnm7mlldbnJ6N6Y8zD1IRK
V5miTqTpjmtEFUSRYWom7U/UwgDVEuWeTKUDxFwNUdbOliWfu3QtWafZFSYm1n8v
ZidcmCBJZDTL/DO58ygmEcgIw00t0NIagSJLBldeH2qv45mweOpsTLzLhBUggDUi
5Dt+8ZLllwdS23GoMz4XQ4m88X3h3qAvDc/rcRzpKSqbothjlUnX+1HcroNoWYbW
hKIjZzpdh/og05Sq+uYmScIoDw2Ys81LNFiRRkF9SyKhatkK0mn+KNw9wUfAF++l
8ZVdE8ShuuJOqbQShO7AaSZJnGD2ZCYIln0E2FDDVOlhV7+JuuQAlYlsQdaaMfd0
B6cVYpaDz6YPCXw8ahnXihuv2NqQixq+ZGIbAOTXhc9WoTPH3nqIzjFSw8XADImm
yX58NLEr47m2U+IugQeD2KkMDY4Spk8djEybRoIDkoKt1bel9fBFcCuFklbcgLRw
oHfVV0Je/IcjT2fYjIfG7SuknPoit3u0o9eiBv/o1klTqUOgNA8Mjwl7tHAsqVXB
Y6AXt7DK1sexFQ1chPybeGt0zdPKM5V07nZJHx86yE2hZtacODn6ltRyjmFdPyWV
mWzuVi3XYxQMvX33cOao7hc1fMP7c5TFZ83c5DCGQdaB+MFPLA3F57Z9AD4oxrQ7
Z7qMXokaL39Qgz5drCa/Tu15f+jGHqOrVxuyC3/Rmy1QfETUymFw3h1XAETWkSpP
GBtZgilTj2YYhzqdgr+c0NFWau+/lhFTHGlrq/hOfTtrF7/06geYkOJeitV25xLY
O1sxhs+HzFt70pucskUn+ZQvRLmcBKX6xHe1WFfMuBTU4wkzJiYEM1YCv9QnAJ00
rbe5l6OyDRY0x9ENbnVAAhAyso5Cy2XywzygZvuum7RaFiY6PfxmUdfy6c6YzhTF
hH6mHzokx1Pjxmj6eIHh0DllGq9J/2MVpLWYVQAKwV22N/h+Y4Es31mU55r0GQKC
2nRSq6MadtfXRDjd7+L0BGrnjiTZt56Xyeu46gqI74InzCcC9gx2pKgoWCvOA2z7
jgAXaPWCHKu0XBcWsKPm6vC7Rk0mVwgcyZiyLLlIV1b93O+G8kaHuM+dFavvisAh
KnwKTkmdbSuEQcGGlX2gYdMtzZAGCd1/ZIl3sM1kslZbCFEeL5laXhT3UXXvAIC0
v5YVmgCWi0QqxccygpjvacT17k39igID1j7jkpKhpYK7cv7exlj1VbRwoyf8Uu0Q
vhS46vI4XnbTATkKW+y2WCmjZGb986sOyWnRtiscCutcn6qdpvNUf6agcLcWXIvH
NXnmUVZT/rw4EKpTggt8mZn7zO2r+bkDFIxw9CwUGiHuBUH0H/lDvEuY3u7rWsh0
sqnaS+ftGLxIB0ShAumZ8HyjMsElb1xyGOHltyb/sfs4R+1EoNFqsDJlN7KfigJO
/zCXoHf0lIVtftSyiTidNmlH2GhNM3Jp1DjxV9JuUxk3UHPGinE8svcJUKuP/zgR
KdkdqckQjJoMyumcOOtWwoaY3ZQr7EAKcnNvD7zRYdA3Yq9oyNFxOs5w7WWeta6l
po/yxKiztr/7HK0cqP9Scrj6tJjYYHnnsIkxEQGfyX57o8ni/gg7D5unLT2rYIPH
4haFa6N53pareZKz/E0vMd8Dbhks8g9z2dsXoanqngsY6uIkeFf1cXU9CXufSf+k
cvmBHaawH+kVSmPW3Uq/8Zv9oCMwUc2rRp5+WM1ANkDkD+xeXVZmWVYd6Tsp9L+u
5Rx77BnbkS4428EfJ2WTqIWFmdtQ6ddwPlmBfbl5W+jvIh9mKmzDuSgEICzDg8Oh
XyUqZTZqkcVWYqq4rO7V17ohl5xQa5XsjysHwGdeCWdyddFe5oNzXVbTVYKyU/pR
9x+cYfsE1mLFUqli+H7IElkHMwKLh9QQH1HiPo9cW3nPyM6vtk9F+pQwMqAjq7g+
+7crjOu459O6EKzb4KVJxLmtYl3rlrN215z2MdI11SDCDBeCSYlxffJfuBmNfPpi
fk++3c/8aV+9G6qwaTs1V0syF04QcnSqW1Pdmfg9TbhKrhhs93XzsFgX5blxgeF3
t9f6fLMUQVjwEg9g0zjwP/KIWfn54vJ9MWSr5ncmHBFOWMH4QtmDsAFqIIuRAyBG
LanaEAOej3WOaEKvKI5WoS6Cd8kHs4imnhxCJWYLjoFrTpCbnK/qZr5Ao09vDZkY
5ctWvw8DzAXzIJLUwzW46EfNDEbKHd0Xnuqd7FMVEOcwTFTt72PbQH/Si328BPUe
AYb5dYknituXL4qqLXSrzGrT7GslwqqbdjUB/9z9FNfJOpRtlsDiW/lwKwU+Z88k
NKWQHLWO+9lqrImoFY4bF5Z7ZqdIUKYPav3KNhnesIl0Y6PZqDagFngPi0r3NdXr
/fC1gMk/4dudd/so0frJHnbE4Cle49f836MfNFsCV0F9A0RwWuVvotVdcb2VwLkJ
vK6LMYvEtu/Z6XGapwNGm0p9kH2BxOFkj/QYqrF/L1qVT3yr63Vvo8yIE7eqc49C
8BzkZ0FIPTgx7uoCeT0de2QtKGPRssB8x3kWow+SJUXqgZExTxqFkyWMk5L+jW0o
ITIG2SVRC27FvUln/AJw4rJnnOT7BhHTTQ6/LITnJv3wMw8+WOM6HGroNGDzZPoh
BtC/c+w3v3bQqNcndp2ne5s6RrvFUjesiBEGjpTs+hXSMGuZtxnG3bgANMS8FSaP
XAhQNY2JF2xH2jbfl2g6GDT4znkboe3dh4hr3U5ZYbBJcpI69h+p420pSWTuQv+s
/wI0En5V3QuIT8DJAMmGAP5OB1LMtdPSqeTeYgAC3kXbqY8Q0caKZCDs/mIywpme
O56tQYu/pmmERzetAQIRZNQPDdw1Jocr6BpyAa9Dn5nm7frVqTBpc7dB+axkInYf
XM7v5cC8cpZJCkl6jOrJ/3F5hFR3HO1EvvrOTQhUKv5sQAAr8KkkI99CDIBRhdrd
3rVbLYNOB31wfvF+bb7+zuIE8GtJcwb4wrzaWBq1ahMVxjl47rGsugkoMsXdsCl6
yXdpKPHNIwKDsXzDTJIKLIHVtOoaU091xoO1cMQ8vCTgkidvJT/ituDOWIoL+d+G
FefLWymhP38qdbTKuhFslbRhF4l+UQsfMogpm2rzbw8iUkj/WwEkjUsPWc1O27Ac
4YdoU17fTr3wuDLzmGy0VxDmNzRBstdQ41mmmar0l2hnCXCuHVs7kUyYuVAm3/qt
f0YS8wSFW/18bhKlihMMD+058CFDwEthUxbZqAW/xyuid/iFX+ZarS7r56oy24ke
aZ7Dfs7Wi9rLMTJLfI9xURZq08bE2XgzU4l74B3Wd2w62gbkHvfiq61G5vqVP6E3
Tna7WhryRmdGZYfCPEvTQLf0FSU67tYhu7sQMDWA5q5Va4U5W1G5mxsw+gi6Le/T
VJRDkJ5qjmkyPwnAaxi2SJ41iKF26SrbclcS6jSdvsbeHpuD9LKM/jJNP4PjbR9g
8S+Ir/fQO+G4ROJ3uCSczIX9HwW1WWiyJo03r4m7xp/fX36Mvr2Skhh0gRHaeaeg
il8e/aIoS6GbRKRXMLz8WDWyQFdN1sWB6D1Wnm/fIrxkTo95ZtqxV8aRVjQTf8cy
NjZ7GwV7of81vFDjgUzCcd6SBJ5ViPszERfS7fQZLZeRrCXsYAlmVglM8Tgu3XyG
laVrJAER7tcGaxEBnBGyl95g9K5z4HYq+N2HybqFhO6GjFYc/6dXS4tVNDCNDr9f
0hQINE6c0HalsYdrDtHiz50nWuUFe49VL7LYUVLUFtw/pTUE+vW8QptmhciEgxw0
Frf4GuaQ7cRm8dG744pPnEW0HNLxVT/abB14W3cnX+aPKu4XgVD71ivwB8vGMUCr
d/nwjbUH5aLQ0qBQUODBXZgZvykOSbzBIRL5Y687RMo3GoIFgXOQBmWOFdiEx/Io
Lwtnrmu509R/fkWxHmELgvN7OsklYhGDJ2L6+8AkbGweTeewQD6A/r8kbe7ULaDK
cOifKurL3bYBHWFzjVau+NsFJZv1EwTSkwqxngzxY8P5boYjRM90Gt3ilzUmDwmi
kxFNfpWfMK+Lofw7X478q+p0LPmHbfaAODjMQyhKzDUY1kE90vMlVDSV9XGIBia8
xveT3dWjhnjcBrAI7ck+XxqwwkMe3xSBSN+T/0pwJGGNol22DuNCxBu2/ZQVbmOX
kTqkhxZ1Zgs0/7O05KV/ki/aIKkAff4iMk5cJHS/TjiS+asj7QNPModrTF7T0V1m
vYrQEyzr4hvd7L5B3BZ6bNDxfekyfUDpJKaa4nSPiVGLijNlNt+p1infk7sW+Kww
mtJloAmI1IOuZLNEC85SXpPGQ08ERP7rjC13ZKIjC0Tltm9qde3sCUPAbOzpF6Qn
SAwURAVKLv4CfXt6NCyX/CSqFKAu0g2bDvlxUF6iJxDW6r7TiCd5KGFrRVmUYGLB
FIBYt6gX8XNTkMMwtSxZ/JDVcL9Imj0ZewligBwjffnAojLyILS3lo40zK0GLVEN
M8IavIter+KkzGYb2b/euQRRG14AXMm0Ys9LKlKU3qUxMIfDkekR6a24d9WLG4LN
aODoFUuHg6LZ1TBLzdbr5RTogOFlL6AszMNZ4dSwUGTAEFu08E5nDz2Fivhdhux5
5wc/c9VPa316PXWhoiuDuIh9x4X/SucuVo9XtYhID4DCA7VGaMdnmfBPcx0t+l4x
rbncT4WzgZHgIIRzPtIAe434ui8rDswvad6N5lRpgkhKi/pWNAust6Bu/v4h9Tuo
lT7kWCqwRP54XWVJ4ewn6Ur5Rq1VhxD0a99F4kPi8aNDckcKWp8t+TZHOY9qQTUK
DJwWvlUioFOO2l9ZD+zFsiiEhzRqNo+gQwD9C6t44X0vkRDCC/UkThmyovoWMd36
uqT2vLENOPzTsMZlyltgTM8mGxRloxsp3zVycPr8gtwMeyTB2Nd3UK98I8K24LNi
BDjR/7SwBKEwfcqwGOeml8he/iUwHKCho7fXyv3apvz9jF+6RJmN4COw+4+D1oHW
TS60MBvTYGkSlHqiOie0GsZXzh8zRLP8Q6zjZMmGQ2R2QD926lr+QrK8BTVZ23QW
ZYqqkjLfihhRKNLKSrpaAE/pgOM6ywPydRGKvYtxDm1pIniVJjFMYLLgejXzQO1a
Q5f2lL8uoj5Ih5QC2VXmpz1o6OPvnwXq0QcXe/ikq5giWQI3DrgDkyBIyAuCZvYV
c/12Zf7JpJ9vC9Ry7OFKn0Pzsw6TeqOqbf+FbMaPnfMBrJaBlhHT8h4wL2pBcKMa
LqAWD/r9Cx1N8i5Gt34RJJdO3QZlhE6rpz4M8LH9lgb2AU5q6HxEx39oio3wMXey
+Scm1nLElb+DSREigGPg48SjEi+DsfCeMVU4WEbfznhrgdah+wVNPcXbkvva4SgR
q5AzsVDJorofSZBP04KLfPRUVuMcaf8VkxwRydmG4/CRbEtPe9oCemq9SZ0S360O
Thx6VA2iXvXuegJl4MO1KnjX/X6o2u6vgdVHJ5oAjIjMuJLeqWxEfkVL7wVC2yJH
aGZ50fKiSbEl/i8iZODQ1d/pKoZoysTR3G3Yv0vMQKZbxO8a1chBk8lgpTBA88vg
W3bugXc1ytb9h3K4vEdFLWRky04YRnw9h1Xe8g89KHQvI9d5FKcxf0las9C78JHC
HG74PxYEyPadZ+LhIa6pmIoKDoJPB/uIylW9jsk077XZuPB2p1X6rfQrN7Vvd6OD
P5n/Zr9CmkLzYO6z7BL+sdJlY8ddfY4X2PbrprZENvPTAQCnSr8CYF3h0WMXriwS
gypH8WI8bNnofC/bNJE2lNhifdZ2tRS4pGscTmck5eNwOf54CdbBEOfhdFZ4ZhTd
9oPgFNqz6ungU61ziQD2XIffZ6suoyU67aAC3C4zjruA9tE9TC+h09tDy8eaPc87
y9gUYK6f1HwDMW3T7f0Cv5qx9LV2XZ9i2HcazioWbrIsgaTBxPCaCdmbt5Br3q52
IpBg5xscM1wIWU9qBHbfpWryuzc6h5gfu468oJqc+XCMRkL5GfKcS1YE3/D50K51
YqRgdPyR8L4DgmmgsOwyvd6Oq16AWVnJ4dOvbDnJXqDhit2d26e8k+rOaWDd+N7N
lifLuDImmRNz+w5JjDnaA/JFGoHSsB8N895NQarFTkso1J6J1ryt3aqIhbi8emoX
7L7dMQNTEbk59WbB9n1UJXIoEvqA/+WsGoesyx9DDZz51ux+/PnwaG01y+NQJD5/
WOv45MmC8dFIpMJLxTK1YbThjv322+71wE8m6XchJuRaOD3AGIgzx+ekagSDbtqF
mdXVuR58rp/7REj7Jvvq1Rmxx9I0LOqGPcyhG5x8VE6rQ3ShRmxAaJG8wvNM6PwR
U3CmD1cRO/05JSM2rQyVhDe8lhtPXXN3fBUfJJzFlGRVbZC4fvT+laj1hQIgVCj4
1AXY0PvAlVryu6im6MsXxJEE13ahvjEeh82rypLchHhCDtSCpvoOLz57WqVj86fc
ZTGvwele9/k+asAoY1naIsaC76RnVkhG2CPjMmIoeqmGRSbSjnbW1xvKFrHCpgqA
yQbdGjJEz4hEFtr/4b9oT91MX2XAA0EtXBN/hvkCJKyYK0vJ2CjqP6kgr5qByA2W
rERkoNh51ZRDNf2a9r7Ovp+LS0A6mlK+s3h/mbwCSZl73nwUNRyhd2lkEAqZpFO+
MwV54V6AePDaoK2ENOuElikFaL1Z3Qa9r6hCj6miINilmWdUglzLBsU43xm7qS4Y
Ry8pfEdNJL0RhU+V7hvEaInlH3+J1JNfT2WsIF8azbPCAUX92ECZ+Han+dK7a5Dq
JGxv54WMeSvquCPOqeXICjcrzvfYUfuHSeRqtkMJkXtgXsfOn2jjpcKCIqVYN7fP
YyAcjHZNSk5CqnnAH2djl3T4B6SHLzYYuMomau5e2bbGGR04YpFgPYV7AUFflt/m
SFKrGpuD13saErLTjtL1QmfllyzLaAg5jeOKj6dJI1aYHsgPTDUSnqP7JqpYEYIg
ELEfJkGOl/j4aNxUMXH9jx0pbE2zB3WV2vijCzbnchyPvTjHPsDTp+I9fGSoyKk4
bIreOFJ/LuV6OxJtXxl5yr9sK1h1U+h/nW+PUoZMhjXus8MaaZuuSWkJoF7SDOLl
mC7/0wyPe7nFvsKxviup0uOwjMvO4RVDF45KoFSqKSXX/BjFS10pOgQVuJzO8Ct/
N1c8XcRVb1s3qgSqhZ8EJYHaBCsSxS2fF0hCG6QlmWB10f4O8oK0FvwjLbJzAxe+
3RAx8n0ZaqHSMnhcI3a8/SHhNYvD9mPeWGHg1FiUotTEqNRYivGtQ3jtg3j93FUD
OpZhFwolJsfNMZe1QwW7FUgzMYeu3VaRTHU7vBz2tqA/tC06UStjnaTAf8899wWE
mnKBTipPwxHseUDKDH2ThD8ZpxHsumeut2czfQL6NO4DlvPjDbZS0lrpcy1oi0z1
eSlp9MoVTJeTNlRefWxSyFVfLNqhym+fsUqTI2rysAQhJ1xrLgbnivOsKZiq9t5u
m9KBlpjQPSbsr+qcvV6nPDaAEDXQeOmWtT/b47Ltqc9OLEHU3C7cgopOwNhFVcE6
tZRyw62HtlR8AlEa5uG2nXpN0np6JH5CBfR3Ge4WItHPc45NkRbB+OW0/FepqB4g
6zmnT4ZdgpnCRjBJkLUOAHdKbeF8ExY4Oilmkr2Rt0ukHO7D4jPAXOZ1jwbJGZfq
IM/EUdUn4x2yUH5KvMfChj6cxcb1/Jsli4mWV4BT9LsZ/6xCbsbfWNRWXH4dRrCf
H3/zyVsJFYFzo5r3z5HWSVhDfUwUPvwHk0tBqRrX+i7ZNATzUpbuNuB5l5sV55PK
P9wc9mKVlzjymZrZWB8DqoEUwOpQdKU0XTfqDp7YkZS1yM+1sh1tqo+U5sw3Stwc
QKxUbQIEFnBEPLis6NLfagWnPPe4dsuBsPH1P1rBLsx0rFPQYDYZLbe19AkrFUBW
oHWZLp9UuQBpZL37E5mnUXXcVlajfQAYMJKiAID+eclu3DbUs72ROcgB9UdsupzY
pkapK0oTVENsBNMo4wSuLUCDR8i2MnAzG6EsaUibwHj63m8tyzBjW8amd3x4K1TS
F5DLrpuYjCozXNH2YpF3dWIrZwuwghkMQaWAtQB/ux1/VsDFpYtTNu7+btn6AQny
LQ9ml9mbSL7mUOsAGNboGZQq6Ck61rrdU8duxHOSxUKnBIjwypSD9Vp4a5KPCG3B
tWdgeKVvPY4td/rmRT/dUHFHwuhAmTjenaOTA084qBsvd7p6VihhAbiUbqXKbZHR
VEtb3cBStMEefrrmu+RGluRLd3dgPE2ShutEXSTvPR6qCLy/z15fwKMDHy10lidu
GcWbIE0yEECjXTkYOWWhtTFdUegZXx1PMSBw/BOVq75ds44+mA/omqa71J23Ksw8
tSarmu5iH1MILOc3/B/ODEq1M4XhgeFa9MlCWseJ8tYRPc8NMJWHtg4zqjB8bbX0
kMoQSZ20aYQe/aMhzryF7OQQeBSgy7KHEEpQtmQ8M54XCiuiJSXo/fVkTTmRgsSs
nYW3an6tX782xTLd6VOl5p6SIxoCykRCSPNDwc6TmDFUPdx1EP5QW1ZLHJ8/1+h6
ErNZtvIU+o92N9TiHBpL72ARMUquH0J6R/4MRi588hUGzdMLlrNw0nKzssJhsh7R
pTvhRGm+JFi424YpmIkMVV1HtzBmUVyDmsxuE0VRDS1OjX4S5U1GXjiCoJqSY7/x
C+KkYqL8sY6GWR8sFtOn9rIYJ/OLVGB6b0+ZCmczdyC6O5V6hP0n44vuDO0cZ1WP
c/blDRzXUhLHDtibPEKn/yQ6THjxkhoUpdULZbd+1RjjVAN2yAewrfb8VTgZpFcj
CD7/qRvPznHAP14QCou9quWVdUD+CXQhRjAQRIC/F/9SX8/XAUiUh5dQP4SZSnB7
9017DuRI74YiVCYjPWxormk6Bquxt0ikBXz3+yRBV4/9471CXz1zP3hlL69iWZjj
YRZIReX5Zprfwyl8dRxIU1jWdCmCLhuwJ0lAY2EXPv7wr9ebCXIpGD7HrT6L6Hgy
AzKPnGuKSYVfw+fwDpEYAJuZLjogALr7UeHkPx2VfmCFBmHFm/meX4qVIl7xXXJr
tswcH8OLCodfPGqD5VSdFLfD+J+w7sHi9gLcerSFjq3NKQa5MRWY+N7XGW/wJEcs
iFfg09yeROQFGgKmM55yH5yCWWoAhw5dY25j+EP4SRHrPvx2KiheNoREtYevXqbb
hjE0bQLIOSSVYFDVP+L7bXUMyWVZ2OVRQfRP1ky0IerN7Ox5wdsW9sov3YyGI5M6
disVD6oSjg+WOqe6ktQBTAUDG/mDjtXLq5Yh+fHcqBZbDl3MMRAggeB2PUNsINHM
gx8pgHe0SLsUB0AkO7qSeMD/JjYA2wvRBvLMk2m8Ar8yKy15UI6eDYL0t1BHJr6y
tYIaLHqiUNlqgicA7+hiBAtNjEoBzHXtPVlep6SIRTmgAUOCUKoYNiaFOhFNAI4a
ezsxmedjks0A4YNILcPSEAmiONTxmRCyA7gj9AtEPk89slxo/r/xrSdwvdXYsRX3
/JZbBjkaAJeRZVb4wf6NM3wMhLchhzYPFPpPnlXlbAINMtq/Z4hxDhMNyJNIgZFZ
r1yk1ewKr/+6r4CJ2XC5Il4/3bKgMoqD3QHvGyzsiuExBFhTWme6uQpXW1ycDI8K
QvDPuwRuorCPS0VMIvdcthbmG2q5FItsYKub6rAJ7nCih9x6fogQ9oGs/hhk1+ve
AWUMfosHaGdxl154mY0t2Ly9XYcnww1xluEMhEJahzaTVI2jXr3SkxUsmcfbDtbV
59LGisysfk8CCmyZw8JGkKI1q/N/snyUmQDkKuscBPJUdeZMougVe18K9oUhNFrj
snQqFd88PdxGPTSpYDtGhMhdx/xSuj1WZTqrl1XupFmFFy7DKPpcb9V1/fPB4LWs
p5uao3EIJYMiyg+YtHGYU5ySmZ8n2RCVPtE2ADZcQ9wsQOdPs6wg5glkPaoPfLwr
rOs7X4GlBfYvivZsFRnCyLQwpGO3DFyQmaDgzrhUin3jAyHFXdTxuJ3+vauOeuoQ
1GbemNo0OTEgCOPLxP5HohdKNmYeImq542hgKFL98ZRYXJx8fVR0ePJe2baW32As
vVIR5/RRtsyFHtuDeqxs92HFXb5eqQlzveULm5dORO7duEgMp5G+vsTCVDhGJpsl
wgrGU8nfeUqqtFZZ6V553wZvRga/625fIIucJ+yspACjpmJA23YPaTgg7bWkonWr
ZjJBEI7zi4GZkb5jfhjxkrPvNNrFbsdotyiUnCSTQ7NM3sQv4pIdNu/4gecXGY8H
w415Osu4dALOaj98aoLSge3fXMujMEeStvDdoYUXuPdo9plb/oODuzjVmk9tR2JJ
91EtA+63uHvVHxvXlid2orT6iSoIzrZu93ikfOYaL0SOHEWqHu1kURXSct2lNITi
JYy/tEI0YR/XGKsVdg+MAL86fmz3SreaORyMTQEZA6NRxL2Lf8dNb+YIFTlfUomI
S8lPnaCefwtiIPBHhuLcM7NAn+gl4JTcvMSxvAzZA+V26esLt5nx01zu6WJUDxJb
QU47eg8GhJEbwkCy7LUX6tPH3CfyxO3JKXWOaXgmckMPNIqepqrLrAbKNeZGd29e
K3r/B9dXnSElseH+KD31TYGg2d0psj9f53RZyIrlm6bcH/KbSIQqwrTyzPFYkYgc
dQGoqAY6W2GBqNWCIj4s8A2ldsMI6ex99PhEFYjn8Wc96HGVP50jRf4juaJyvTIz
mfQHCCd8Ve/Va+D7OPAKwa0P+sZQ5Txp8ZM3L1878dmX/Lw+2Uqz/vNn+20n6aor
NdlH2CPFw1hnElu7dXLqYWcGdRJHtnJInTbFZwYMh4Z7T8fQBBlnWd5qpTiMH+rb
u8kGOhIaT8bjWTRVVleUnVtjuzbNU0RuJzjViC2K+A6h1tdYsyfT4iU9BY1u7CBd
A4lgmkgQ7mWmg4O3Q4OVdb0RYiwCdV4BC3kgDqheGBtoimxkFZILmAAE0kS9zt7J
Yvu9Rt0jWNjHwOxhUJDLw6Z4Zl6odfzsNt8dCBXT7eDPP9CTkvoKwpyrFSZR4WHc
BaqVN4as14pj1JO+cbVqfIajixSshiJKZMi06lkPWBELUl4rSlAMYobs3OBVXcpu
St6YfRZjzEEGYQJqsq8HgMXJwO8k4t3SkVWT3kscm3i3WkjFT4nQlap8+2CgJbXm
OgOQDNzmR0s4C1OYVOHOWhdSVfPGvKxI1WyacKCJeh4gI/LxTMmkipb1jgtTDAtN
q5EgP13iJClq+BBarQEm9MVv5YGvMrYcZR88E7wOUATzKVH7GMWunlAgKFaR6VgK
`pragma protect end_protected

//pragma protect end
`include "tinyml_core0_define.v"
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
J6cVhJE1teU1Hem/mVUCPxmy5Fgtj3Gtp/0bZPbl4s9SlntbjCD1lrajrf++uBvn
SR2FI+NxI/xxGT11xV1wAXaeZgIKJSB0k1ytt/lIlhgT60PalwKE6QC8b/Vv5m6H
3K1U0XGFnX9LdDX1TvtgYPIpDbtYRzSvwe0izNqtRSxAcfTEvY/TW0IpwI5RDDZS
VJJRwZyJSHnxt0UA+NL2ajsKwi2IwHhoPY0/mzN1fvYplZVD7cLO7m8a2ey/U0UT
5oG3ETgrxd0woGUqCdwOIw0M3zTPUmfYbWjWD33AEy7YQvhc+oyVRhALMwmlweKI
z/nedbm5BaVmKCACZcbigw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6400 )
`pragma protect data_block
L2ERj401YEA3qe1WRKc2b8kSKpySMPPyCsmUCOPmnjqT+TzClZUfZbbz+PQzPKZ7
O2FoTJTY/fy+IsbMelmHUrYfglkhahr8rNqWv3YcsHMrrLeb6v+Gb2DEW6Olf3io
oZPHiXGSKDyXff6u6kMphhFgl8+VAKRve82jOaRupljBBfPyuGQaRftX6NDCgxWI
ljD2Fh/6TQmL0n4V879ZLoDmzQ5g0PJihVNJWkmvxehYwGHbCgtYmTJLEkrOYlQE
xKYteQWA467YK2Twi3P6a1OjX7/7d6tQvE7cvZvqJg7nbWudHHrryPmpLxANWLNu
xbj2l60yfkKa4NrkwKU0lSZQWleym314DbeytHnWGfw3Kmg7I6z4osxmKtj3+lIj
RNO7SKSuLOeeDWSkV0qswlDdJmIJBij31aFiUxxU5czUi8BNABrNW9gZLmSfzAJ9
SrGTm/aSXoLiU9qg+CwmgN+fkZFeYL/+PjQm4ds4EPI6ABBTNW2+ePlHw5rDZTmm
7pVTUnlBjvr60jJd1ot4D+FZtgAlZOe9f4paQOVqhoH/gK2h+dxf1GWYtbBbY23S
5Gg99lZecyvI+WYD5CQT5BssuotljRFSVXxfHRhOhlJLJKn2jbKsZvQqR0h7TPLD
hMYlgyo6X348AZAXYO8Y26f2aFf5lWSmhHJYVdtj9OG1ahsp8DO2uvCPMWCIXADS
VXuHsURXLzMAou9EcdstnJSbGcG7WBeHbjNVoS4w3JjMSJxIzVvzu2CuZUmBgFJa
POVvnNb27bVfaiocLMwePiBwyBOgi3NHuRu+jJMq+tJR7Fu2BCeytLfeX+o3KJdQ
I2LhMstcJr8Ie3pGrjYVwYVwhKxrSLipy7NYU6C3sCHOF5X4Km7iyi6JG5Tk5kGr
Hmcwgxuy7a12n1h4B804GIKgfuaO+6YpVLm6wso2WgsJOVGYX09qt+QIz4e73LPL
hMKg/6apvrMIulQ0uZBG0O4QK0fwcXb8N1pCZMBytnJesZe+IgEg5/dyRPZtKUMq
E5mYRjELnJVw/FNQiqeV7seKOth6qXa7GBNH2NU3LGP7wmEyg31ryJHg47WWmlhG
Lpmh6kIFlbpawrvGWptOV52C/ZDZGgtST3bQ1oyS/hlCU+OiwTfEQ1JtEHist2ps
9tqPEH/iw+58dMPXhbi3KamBKBn20xc6+yyeM69/m4OWevMe86CfBnix2hd5Anx6
hWm5Bv5S2t32F27kZfDNHKUGEnaqO+y4zrne9wVpzJfDyYz+Ow0lobdtP86K4DrP
wZps1LiArrIhvYnyQEf2Nu7d7gtnnRO/XZ16xxO5MWEXRk0rGZyU1OV8U7NqxgbS
7/TcDGsZ9bGjrKjlD566cgEPFlZz7S5KZTs1hgUCz4v0fo8Jc8ynJBUx5CjMyNQn
5iCxc+UM+0GGxw4LVqwdQC07dt/cOfcNuOQc86MD7kTDWdW0hxVO9dYXTNsc2ei6
LlFf9b+1dJTv2XZeoRSFWYtX30nOJNgI7wO7rEHDCP0Tx/On+is7K8CFoMaoDBpT
hn5JoYruw6cXp4wdthlkgBZNiiBiiqd9k+/cI6YZ/J9y0fDZOWy3Dlnjlj/xUkDc
5oAuaYOj9sxMEucZzqMXvlkIShG002Z+3HaHe/FOb4ENwDwa0LNiVtwiaGyA/vtU
de6sG+b6KRqFL5vzFfXOhAto3J21h5gthpPEclPjyJ3fTd1XF1kugsB3AvVt1T0I
rwWlR5GKO6zcZAUzvscNhy07J3blHav7VAWT3c2likRqvmySdL4mO1ClS11xU/k/
43ViXAHYuclIxIjjfARCXNUdVRgZAryUYoWzzVXkmJJqHMKd5l3ZoiVljOkE+oVp
PIWg8AJqJsaRfpSEaUDOeWM5ospHJcQ8XPQisqx5eg5uRVE6oWokWsowlNwC9oJe
LppiSegs/undnMLtClzcKQ7fQep/89Mhb8Wh87fCbA3Wo8fVFuJZUG1f+OjUOFGB
BUkJBdv695cpBrl8OnEu681oPD0QkrNvFQZ5Zh4+PZ2iF1AJA/bDn1FW39BXfrYA
UrZhYJvKbkF3OrDTOpDkXxRwltmjzje6tVgoxZfGRPAPKDKea0WuK/tR3vgBflxy
tKyyrLJf12XUfycGPsmL5JAEod2zIimG4zabnh1Z8B/9ZUR7Vbh8jZRoFpNqS/VD
EtzoIbre6bu3tffjFR+3Qd5yd8IRQv6I5JViDij5DoHDQlzaxjrWCwSx2W6LNmHn
kCDkchWwJ2VL5va/H2kDmItidRRkEW2t53uJTCYkpVa2mPTredUNPgR25ZDFyKwj
h6VfBi06Ilru45Y4Th8wWx1FSjNqwgKcnTm/XkOcVcxTDMyT/lrCTYn4qfqa7LOO
Pomc3BW9FMPT1AAoVUxeB7xbDSfr5mmsbvMEnq7K3Ii3wB2ejSIOS7XKw54yqtp5
KIK87ZXntfNzTzeIYCzY8UHIxN5pl71fUN8nuqXrseUjy5sEzNW34hQnLQ12V0vG
vZwEr7ATe46gj5j1v6rVRul7sndRxys8Q4tWCMV6lPQdtiSHK+6cGzOF+1wlC3cE
85E01EHCVPNzO1FEPNGRqx8LHVud3UagocEMMRn5rAyg4CWC59ky11PwME9XShJ8
7re5TLtWosrEGHUMJxzO0dS+U39vST+ZmR4RxEtkh8N0Cd5yXUyjImDIRl3jcWlg
hjRUyxeOS2QoAU45Ik4rCCn1DSBwt2eLYSlr/5+/DUwZ9wKVbG69XY/p3V5zH6pL
yI6e/qwQYk8ijWQKqUBxAW105H0LSpg6W/N0J9f4iF0O6x1C8NjBt+ZUJiQs0+6G
Xde8xHkORNi/U5Pwm/4jdwUj5o26ln3MpEPTNCa9qzsHhShwWWMr2Sm/P4cyL9Vg
iWwO0T/iFm9490ulYpUoyTpi9Gce5F3kah22EThlYDgKuU63GQ+hkUry6pFU9Dxw
5Wz9MFPNS8CRiRnJy0Ni3eK7rZnEgcd5RoN5nHD88MDNxQU+VA1/bnb1EI7xpwkr
YQhFJrnc7tumH7ef1ouq6p3ceCbZFF7YLi62yE3JAGJ5UEQWAu5iLdWUpyT3FHj/
CQWvDiLFDu2/4VWSkrru7woXoz/4yOfwC+A7fQKKYhFhu/Ghw3Hb9cL6WZurlpL8
n9yXlQNWHZtvQJWvQFyxhxYJYDKu1eYhIC7dafCCr5LmpshC9Pub8h7VwsB/oWtC
w41v7fKXQnJBoFcQ9sladzxY2H0Z/zmYBoeXEkCFsd3R+2YjCiS5HH34JCziRUea
u7A8PdZu82QZ3SBG6uGBmNPWFgOpMErXcAvzHaVOBvy/rLtiUMWXHVgd3A7n148+
8ICP5+7W2eX5W1Wf9sTXbiYk3vNK3OkmY+4YWWKUzLgdg31v/opj2ifC8e2U5gEw
XKswvFT82it5EiS8mRAalWIT7f4zqCOe6A8QXxpgkg4nEayiy5x/FJsyEx3xQ4dk
MlckgCLl6ucUyJvjUxZfXOcIxtLjaoBUR2rZaBYVgUyXkXxVQ/xadQVFqAmkyLWs
81JwfSItqksJRuUjFdAQc/QRaiWr6sGCzHVclVmPtCgxqpgsMvNUXkY1Ir+Gb1sN
DCsjugBcpy8cZF9h3IYCL9GKa0UtruPihau636mrvJlRps61Nlh5qCjCgbwfA5ca
uvmiGY5ZigxMnaYL99QSetYKfixKKfiB7B/KbLimfkpCBr3snpLOuitA4AE5YL0F
ejuE0YNIQTyhqe8zZ3FBf3zF7bS9UZidAoHPjPkSM67qPkax69vjAGVPTPOq5YMp
+3tGPnN8lVI2LttoVHK2wDEOYjI20+QD89S1qmcqkpxyjvywaS0szlwQI2VKu+eP
dyidrgC+69Ic1LJq9ljecsTzdsrM8UX6jBXN6GV8xaHOVldwZfw2ijhICz5Su0JP
5MjEPxE54xv5AScLVniXjix+1ZqP1JqxHSGFQVh5ZrosbZBkKbJ3KnNqEyVP8g45
gRZgcyUMoJ7Oz3AxbiYZf4FJYjEc3zAp4t4t0/kPKlVEJ2jTMLNruB2QMlY5VN4W
IU89SfWiwvmSD8N/2LVyMLJRYLTHfCc56CPK9su/e51gd7dG0xXGQFLK+GUU2ZXP
/jWLv4sC/JcAhKhGaEkLadtWQuPqgo+MLFD7gksYNVJorArVBt7/3HRD6UARpcby
SSHgPO/Ris0z3Zjnqkazh3I3jvXSv3+/n8vkQ7u7g07N2pPCLOMgCVZ/fsfqa/O6
KR5oGboq/y+1UvyeQ8I+Z4hvg3nc0NyKsmjTj5sXfcffSCgL+YN0JUJvS5ZJozoy
J09a12bBlu0JFqWqY9vpb5RHgcENxBTWvJNNYC5dG6c7GLcB3MM9HZ0Tg1nCbnwM
9t9vG6yJnno/II37gTOx8dhD8Ixdjp5h2AZS2Rkapz6frzhmzhASJ52IokTZyKix
CqBsiG+RpEL+hVYeGiwkrG8mGHTHd+TTIwabddoCDzrHRC1/S0UKRagdoGa2XKZw
32doLvXoTGDBsQRY5No4JCwz+SYVdb/1cySVqhWiaRpw+XQZ/tZODQpJtYdb5wMY
fHSo/KxRVPk8Q4CHG/kZctCpCbh1j8MLdUogQZqD4npPrRyFCAW3jS18wdIqBe5Q
BfeXuUwD6V8fJocFxOadIo8UgeUs7A/9SslYz/LEOKU67cWR3C/qhAKX1aID4hGQ
aZpnoD+NsckCe9oW6GzDfRbfqVfFJckHsf4iO98Td7z6p76PIVF0oSjq79LyehzT
dX6/9vcRPpbxEZklVQsFzBiDUUMI2QdbeAhAEuRn8akCnKPSCvRcCbNAdvNLWS78
21+EIwjjCSQds5RYYvtme92UruNeJWWhroc7oRrYiPpIoW3SKGvI2rnoRGua2IcQ
+Vqk4YUHBJWoZwEYj4AZ/Pr3Eo0AxgTOTP9eLP5ZKyMS7UhWST19BcAwH5VdQKwB
iGk9lkV4+GaUGAj/sNiyk+hHEOUfAWGHcYVfMBn3P5LIuJjfzqulNBoxYD0tgckn
MQ30zb+5N1TP+AT8Ig3yOXPlxSqy9IlspLREBNYymq+tW/1um2QC0ERohsn9pi8F
99DTAjS0WLbLaeYXtfistN3VK1iPXi1ZiwJvyAgs/Y7sodZta2zaFzffT/H4ZbSA
MMpI1sDYYNiCYvzENahQy9EvGAS8Ulh3lASxC0qB3AIPipY1DJ5B/BvE8np1lfLj
AelAkc+Q/cRBqsKljFdzWCGAz2XfTxWLX2HtV7FO4h6Lj3xNER8pxBl8KE6DcMIn
/e4QgCLrehrZpSW1HN+/9RQnsgn2WPzOIsCZS8vRj7a/AkGVhuqqCKuQoaiTs5eJ
ZEtMjt3OYc+dtiuGaWIB7VMzdX1YBTSBnicspUZQ02Lv6In1PJRKDE4DSZufczkM
rRsXr5/BlNlIv2z4atcxLFn4LSgEBVM7XB2HBYFSrhImvgicgdfLKvHL4E0w3Dua
YUa1X48Q/mO4+lT2XP1PYF3lB2pT4fVOHiMj6IgsKDWoS+nz6NPp611oEc4aYwzU
8Nl0ukNLTl2ckES+1gFrNYQBUDqEC2UjvrI1aGn4MOFG+by5kmzWcN04ui+Ibnri
TIJbI3NOf0VcrLuqLs1ZEptYmUQHh3+Vx8hKGdDq7NDRs1hPuDSNj4Pw+ZtP1XFb
oOHy6itUc+NBMluYSZWC1xxhDEd2D6TYwJ4ojMEmI5tEFaLToHuJM5Jgx6RjHFcZ
OA8kGc6BBIkWQ2ATNy31c1R87w4Gd2dwDV4REOOFLZy507Poh2xd+B8AjiDcd7Vh
uOQHke0/cQCHiD55I+FM7BXTrZEutKzvmhz5Rt8mbtgpTeeZT1b0jxi9oWjTxC74
zhqj94ySCRaclw1eiz6vsKu3BtOQB7UV9T/cca38jjmGBhAUCwPIDCD83FS7LY8Q
Wi3AJ185LXMZHdV4u7QMiJHutimljsDrcCBEiUtwqYdiO3X6UXBP527fFZxBVWK/
MB2nY9sAuvSaAxtY+40okRzeN4VsV3P2H6ahM9KHLLaHr6SI/EPGeHMzF1iKHTxs
rVevMqn2eYjexvQ8avulD9FYMpeniACB+6nAkKu2Q0zst2984Qilg/JCkQDJiTEV
o2+lcOCtLBd1x3QjEpiOWtefNZIxxePttz87yKns1XUCumshg+BpoylyNlpCOo31
ir37Bt0VWKqVTkg1IxAMGRB7QgY6JpTtctfp/RvSmaa7gvC8E05ihxUtAWVjjZuK
uV2OEzvceC6UEAApEnNliThNgP51dLhbXAloowK8zWjVMrt4v5wVOvGXg2PE2zhR
EIQG49qJy5qiGes4cRHh2Aao2DwiK8hiZbbfR4yn0xPZN2CVA7eEnEMoMjvC1S6F
9dVp/ds6Ui/FMmOK6ZOol3Gurn8rSRxvQ6ltvf+r2TYIp88bzHpzmMqfhz/d5RmK
LWxdJXQfjtK0tL9HdhAZwRvnw/j96lhoAySnmrb2fWaqepQrcRo9t+QjPw+8MGbK
Ejg89L7pIW/UsC+ZkXXOwwKHtjM7RpL9CHvoVL+8eYdOpq0b+4OHrg6nLXcmRpVC
wQ6EoStB/45PoIL+i23NX151nXl5FFqx9Wzn6zf+tr8+LvmXtJikIOPYurq2MF3Y
oIQ95MhplTFJw2yppKW6rsjdm3Lz0HxhhQA6iX5+kApA8VWHonQOThZKslPtiUn2
8GhDCLodWM+23mCQKNxIkXCxxWJRfRVVosZLeKjFcjX+bQImUleMpmKCYC83VGRL
WYN2ueF6daxMsCQ1bpY2mvMiljo7ziRCoyfsCG0cUq9tgKbqSeAYlr95UQBdQlQI
vSBKR6gw1SPojwseaOLiEAeGH/DfvvS4z4Nb0C0J3+hvzdL62C32omvgned7TuET
/0WwcRneTEtjyS5I45tUGUxoiQ/qnwclOTbxJfJe2q1C+cXl6+IzRWYplTdQdXGv
rlOCIqGvch4HopuVFu3XfqVMIew3wtQn56bg88i76fTEnv5IXAQqYTW3xdlWzyOW
z0oRtc5/k9B0B9soDk5MDFffLA24XUCWrjI8Ec0bcSzvw4Y2EWEnPzCqWanu+qBq
jWmKHmAKYMGjqMR8a4rMnIA8XRhev0sMahscw7d+kDkL573H7Mic7sG0nfU2wasY
+mst6Zaz3OyHUgJIRqtAzeXEOlovexHGNJSc+jg/iC4VopvMoSP5ZasWuLmbari2
O6GOmCmIth0IKM+UeCcDYtLnasV2GysH/CukIOnZjIZ/Dp09BP1TaIFlLcQSe8Xx
dXZPdJXPvmrQOz+FB4AT2nDc8YJg2wCciQ57BDFwNzRPgg5qEKoBwMLWEnVnfpOX
4gm/XtgO0UTW9Y4LkvyhF58ewQOY0QcvgGcXRKXE+PoJuItQILg3b1XuqqtW3pW5
ZxUxp3DnQL3mESPW922Jc033MhVrZtbYep6Ct5zNcJmPtWiHWpxqR1Hwrtr1hY86
jI4mlZSttDp/B5qG9MaatCkvpvWm3DO8jZobtd7mszc5OX+xs3fH2z43GdGrrNeD
rVs9xcx/GezCsY0+rAaf/qVjJ5SC/rbCmY0k6gQeP3J4MwBp7Dp2FB09rg/Sy2DB
l9S/ldpJhpREdSUkL6enu4xrZfNekEBE0l5XmwRdynCknPIFi0gX4fNLe2qnA09A
6YvgutwELNwvniXI37c6QMiovsnmwmrFv7AcitL+Rhepx43mD7IPmQfcpCBDvqV2
OEr4TdXDv3r0yaWykpZnNSzFveIeiey+PGedxHgo1PCYGECZ/nDXxg6569m2pjJM
YLlWRLCED2w9FsmJXiBdDZlDXRAfGxzdvBiKaZOcF6uj3+aQT4KAQaTvRpuj98A6
RYfS//+Zry0opQUd3johCoWT7VAB9XpVkztJq3bIjmrP0uP8mwl/OFVU9YQ10SgL
9+xy6BxBkoCkneoCNpZ0XEb34ZvL6sesKPobpO3FV+lpy4ZmnTk/gPZKO5OSm5S8
HrWbREdeT21foyBUcZhrvjjzwkaGnJwQFurlxxHHPB4SSnP5TkV/rG5PlqcX3gAN
NFnKGwUION2pVnXBTGjjwaxuk/R/8sVLwUqpfVddRfTRB6Z989Hl3w0vophb0hTw
Mp4zMyBmTDXIIKyLCHTeBDCSICLQRTYjuuKksiuUcMztQLEjq+jmGfioDZkKbuML
zLFpgueiF/amqlB+s6SUbwWnJddtrpVABTREia7fpAeHCVIIrbgI/+DDSWBdAODV
BGJ6WvkMPxd3P+kRM0Pjs18nmn66KcSrZoz8YV/WilRxscilpwMaYO2X/joI9fgs
G1lsA6k3EdSXPKbujQB9CUqjc6kQbATaUMfom4qImd8qHfHpCOMIU+r4x+deEuW1
p/1YDJTYZG1k+S3fKH4vb9O4ucSFgPWCq/Wdl2eh2shd4rPi7EX/biqA856eYLd9
gWL7uWvUHX+I2SIIGvxNqT+RpgKg7Ty3MoLkESdXIEJNWjtMYp48HQJXxAvHuQuf
v6e1FP1EZoDVdtAdEZxYN+9ptonCpFgfV10qBEHmZK4/XSu9rvOi9MN/x+yuLmfD
YKA+1FYI1SPsKH5k7U7w2Q==
`pragma protect end_protected

//pragma protect end
