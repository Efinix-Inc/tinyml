//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2025 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = tinyml_accelerator
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Thu Jan  9 10:42:58 2025
// ***************************************************************************************

`define IP_UUID _3ff0f8ede71aca2c69dfe983eaa810b159723a3c
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)

`include "defines.v"

module tinyml_accelerator #(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 6,
    parameter                       ADD_MODE                        = `ADD_MODE,
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,
    parameter                       MUL_MODE                        = `MUL_MODE,
    parameter                       FC_MODE                         = `FC_MODE,
    parameter                       LR_MODE                         = `LR_MODE,
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    //Convolution & Depthwise Convolution OP Parameter          
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,        
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,        
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,        
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    //FC OP Parameter         
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,  
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE      
)
(
//Global Signals
input                           clk,
input                           rstn,
//Custom Instruction
//--Command Interface
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
//--Response Interface
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
//DMA Master AXI4 Bus Interface
input                           m_axi_clk,
input                           m_axi_rstn,
//DMA Master AXI4 Write Bus Interface
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
//DMA Master AXI4 Read Bus Interface
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);

`IP_MODULE_NAME(tinyml_accelerator_int) #(
    .AXI_DW                          (AXI_DW),
    .OP_CNT                          (OP_CNT),
    .ADD_MODE                        (ADD_MODE),
    .MIN_MAX_MODE                    (MIN_MAX_MODE),
    .MUL_MODE                        (MUL_MODE),
    .FC_MODE                         (FC_MODE),
    .LR_MODE                         (LR_MODE),
    .TINYML_CACHE                    (TINYML_CACHE),
    .CACHE_DEPTH                     (CACHE_DEPTH),
    .CONV_DEPTHW_MODE                (CONV_DEPTHW_MODE),
    .CONV_DEPTHW_LITE_PARALLEL       (CONV_DEPTHW_LITE_PARALLEL),
    .CONV_DEPTHW_LITE_AW             (CONV_DEPTHW_LITE_AW),
    .CONV_DEPTHW_STD_IN_PARALLEL     (CONV_DEPTHW_STD_IN_PARALLEL),
    .CONV_DEPTHW_STD_OUT_PARALLEL    (CONV_DEPTHW_STD_OUT_PARALLEL),
    .CONV_DEPTHW_STD_OUT_CH_FIFO_A   (CONV_DEPTHW_STD_OUT_CH_FIFO_A),
    .CONV_DEPTHW_STD_FILTER_FIFO_A   (CONV_DEPTHW_STD_FILTER_FIFO_A),
    .CONV_DEPTHW_STD_CNT_DTH         (CONV_DEPTHW_STD_CNT_DTH),
    .FC_MAX_IN_NODE                  (FC_MAX_IN_NODE),
    .FC_MAX_OUT_NODE                 (FC_MAX_OUT_NODE)
) u_tinyml_accelerator_int (
    .clk(clk),
    .rstn(rstn),
    .cmd_valid(cmd_valid),
    .cmd_function_id(cmd_function_id),
    .cmd_inputs_0(cmd_inputs_0),
    .cmd_inputs_1(cmd_inputs_1),
    .cmd_ready(cmd_ready),
    .cmd_int(cmd_int),
    .rsp_valid(rsp_valid),
    .rsp_outputs_0(rsp_outputs_0),
    .rsp_ready(rsp_ready),
    .m_axi_clk(m_axi_clk),
    .m_axi_rstn(m_axi_rstn),
    .m_axi_awvalid(m_axi_awvalid),
    .m_axi_awaddr(m_axi_awaddr),
    .m_axi_awlen(m_axi_awlen),
    .m_axi_awsize(m_axi_awsize),
    .m_axi_awburst(m_axi_awburst),
    .m_axi_awprot(m_axi_awprot),
    .m_axi_awlock(m_axi_awlock),
    .m_axi_awcache(m_axi_awcache),
    .m_axi_awready(m_axi_awready),
    .m_axi_wdata(m_axi_wdata),
    .m_axi_wstrb(m_axi_wstrb),
    .m_axi_wlast(m_axi_wlast),
    .m_axi_wvalid(m_axi_wvalid),
    .m_axi_wready(m_axi_wready),
    .m_axi_bresp(m_axi_bresp),
    .m_axi_bvalid(m_axi_bvalid),
    .m_axi_bready(m_axi_bready),
    .m_axi_arvalid(m_axi_arvalid),
    .m_axi_araddr(m_axi_araddr),
    .m_axi_arlen(m_axi_arlen),
    .m_axi_arsize(m_axi_arsize),
    .m_axi_arburst(m_axi_arburst),
    .m_axi_arprot(m_axi_arprot),
    .m_axi_arlock(m_axi_arlock),
    .m_axi_arcache(m_axi_arcache),
    .m_axi_arready(m_axi_arready),
    .m_axi_rvalid(m_axi_rvalid),
    .m_axi_rdata(m_axi_rdata),
    .m_axi_rlast(m_axi_rlast),
    .m_axi_rresp(m_axi_rresp),
    .m_axi_rready(m_axi_rready)
);

endmodule


`include "defines.v"
`timescale 1 ns / 1 ns
module `IP_MODULE_NAME(tinyml_accelerator_int)#(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 6,
    parameter                       ADD_MODE                        = `ADD_MODE,          
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,      
    parameter                       MUL_MODE                        = `MUL_MODE,         
    parameter                       FC_MODE                         = `FC_MODE,           
    parameter                       LR_MODE                         = `LR_MODE,           
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE
)
(
input                           clk,
input                           rstn,
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
input                           m_axi_clk,
input                           m_axi_rstn,
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
L9wwqiZPzq0uu0U+FWui7UQpf4EfY3AEvigG28kLynKuijunck/fN5Grqmm0dZ9r
lhdbp7tMHMgojGHlnSIC9GszKmvUNIoR+EPPduNeUIycjN00fYYHFyORi4RaDKX5
Hv0o92chWAOBAYdPDx6LGrHhdcdtr/iW4z1KhApHVzsVit2SMWepVUmBz+F8+4ZM
xJlsLtqRfPLsFMoe8HYBSsBmIFOxyisGsi9cfUt9lE6LWRh2EWGWkT6VBY+FzW8q
bqiiQ/p1VK1rw9ST11hsd+zlC1lGWZcsuYFEHEPUgyMb5xAi3lzsJxMO2uc/CUkN
HM7DH2bdrXRBCSirf71zIw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 59360 )
`pragma protect data_block
AQLS6jAjJqxeqASPVePfBhvYtHHyYrxSH7g2222xKLqz5wJKYtR5AfFDw+kW2JfD
L5nN9QC6V7D45jGZkFXrZNwUkhKNL7/e8oQn18iHf3PXOOYtp8TacD9UrU6wZMQD
u6ja5tjFDX3DDFjwvGVt9R88+qdG2PLylAZI/fyFrJqDYc0m0JhZeYoRzrIhWcPJ
h3nxoVPyhKnCCoxQSBZMpiX7rAXrA9WRccK2WlYPC64B8n0C28bo8VDBPZTnyLvJ
HC2UY+x6CF5//i2tNRYsFsqFsSRxGyOH7b/QQZCMBoWl13iYTkbu5B1yn3AxpSJ4
FgEew1mdl77qmQYaqvaMemUezdcqMHweUBfOBxv57H1Py1EafeV8KkD+w+FDf7jS
Byf/sn1JpAAEgZV7A1rJFo3WwWb3BCpXDsBsxOMSBUTnCsjZsrBo5FSD6UYZAn98
/j8zIt8BtciVBJAWJBc6IqrZlXvhdt+/fZkHIkKo+TB6UMUCqajm0p6QhHK6lbdD
UHQ+Utge/o0XNi6ywaUvDGzRBTtVE29wau2upy5YmkSlkC6hRveCpyqiWNW2i8XS
ULYLaWdSdwI/yr+sis4utd0SiZU5H+7EsdiW7w8v66qk+8avoT5Dv7JrFBTKpY3k
JhMiuLUeQ5W6BG+SeUHxA7JwgQ+fM8KPrdpXh9LjeZCrti1DjKFpRNOJDP7k/bno
BojftyLC1ukitgpeVB8znhX7Z5c8i1fKWAzBRllUe5CVBPmYsKES/jrceBIb7U6/
Kdfd3TkkAnePupldY2DhBBlmokxmvfJQ+Q2C9K9yivep+Clv8j0qFXNE/a68rTny
E6UcAqNzdcoDA33vSeERmDS25XZsNJHCnhvtV5s02mU8ArOfoxWyiz9iSgCGQNBF
pIJK9UBjC//McVau1AzI02of6PcWxMBe3cBkLIs9nhNAaL23DDCMbuwmwZzC4h63
BChHmRXg6gzsu8cf1JIdimrOHV9N3XJf08AYgNeA95WFmAMzY2UG3N2ZpE7zbgVE
S3awEslsjqK4VYB7FT9hdmnebQy9UgRaNaLly2rFfC+e9AEdYzkhijIjM4p+ddnF
118RoZm4NVEl9f4ijLFV2LPgDpWgwa/HIRj7BbkhqmvXIr9d1DrplKAwYbnkTkFv
Z3iB31G788pDQEpxtuyEZv68YEVqEXUK+WI2vNGuqnLlQnSflTbPSymeQSOnAl64
zhX30XSyRAQJaSwRly2c3dj5wKtXTO84KB9KN3DnLim9UODgYmhJcYMR1ExWEu6H
54P/udQPGe9SUPmlshW7tDPFHcP3kkE6AjSHVUB8cIdQd+HDUonhMWj+Qlwl9D1V
a5hd7SDwO7twm/4p3GEoP/UhrznfeKbnxMOvVkeQLdw+KOZTBEVOxtE0XpZrtoGj
+Rk9E0ifxZtPsAPUpyw7z/+x0fYYnpeaL46rTYuPLfkmecbIU/XZk3rOE88gNZbP
bKAZqPdexnL2dAIDlZUHpM8/9VlynnFP4H8+9CDWiMI6l9A+75gPn2nSAf5/NaFI
RBoEf9v/HLxeOlgkn7z0s1xfPwYnIG2IvHgg5nDxY4dPqBNOkWeaggbNjwQBBAMM
breO3Hhy8UJoafjDWI1Xczds9J4N025kHeLSElHPCqA2pyj1Eu/me2FEWMGi82q6
WvhM5vmtoQd5zGt3jmbF8kI+swQNmcx60L8hcOtScB3OVN9wEGuYWg3H2ZbWK8DH
Atal1ca6ZwyKUzAUYB8NN7zGEryK1/0NAuwr5dCwvg739X+qWZD2HHSnnquqsax3
emVwkaouvZEbbQ1KBp//zmQAfJVjKplUpSn5jbw6MTW6PBuvFbh7ldTCzlLJjhx+
Z2qosetNsDqUfZHgsDiSvBDSZQ/5z9wJKKqDN/XYEhzA+n1IFlS9K28SypFcn4/h
5ZCZ3ePW7OusAdX51Gf7dBciQidcgt60OtlXUU2cJZipk5OlNGevclx2i2cf1ZF9
fhJ+Om1b1bEWggXonS3k/WiURsMwfAfrwlgJsMeyuivH3hXl//65znEh6M9ILAHM
8Ikf6QHtz/2/DNSZcfIstuW+XzHRkBAcHODjQNbf/51lhZnwAQOONGiXY9hVkWte
iFcKqpwm/qaPfpyxCLSO1u69PtPORE8WPP+eWLrwOtZ5uBIDzusiwjlqn+4DFTj2
Bw23jeWb37W52DmyBL3HB+4nQTsG8kH8UfSyidN/fvSDeWzjz0MTq6s6ffkhY8M/
H6xWolCXqS+WWVJ6eQhfsFYUNqOhBf6Y+TC9p6eFWtsIpMiUOePHmU1ReQB33TJn
2wW9TNTZxw7cybtlVgMcwEq3XUhXfCStJnKfLbZRgsk+xdzYXmF1PujzvAfaiQaQ
4jsEZeDoknyLvGC4Wd9qmUApxg8U+grRFEkA6Zea5YOIyk7FmZaiQautwVWh4qiY
IKoOmlD1fN4zDDt6DSrSEBXVa8NP0wEE1tFqnE/k3HLIViprYQVWVdzH44j7F8Co
u4A5kcVCg467yKtT+/3gYzgWY/cVuBogTpVIKTuJ8FWgbDj1fFA15CaeL2zXnmnR
FqX4iNFCxESkRb7R2yAZ4PeqTpAZi8K9xm7muKNXFRDa0odUl06sGfViwi8LMas+
1ttyVPIUYN+ieJ+XWJ+x0RtS9a/N7c6bOwwJ1I3p2bm7IRXLsm2k2Akce13Fwlu6
TBW1kvIWrqqMIrZrVIgtR7sW3NvuncKu0lCu4iC5zNJW3yOSATPWJ/YtFCUEWQ/W
TGSp39/R9CGcCzhN8RTIC72xX8+BngX3DMjiYhdUe/CqI8FMzD9MnuvqEPxlXqGL
WIhoEnBISe5+Wrs5FVkJMtC9yzQBwo/Q9YXU3DerS4udN5eiZMbpOyDlYz7puZ1/
zz3H7TAG9ARVyRdK0oG7gjiq2AhTSDJfHxDXsMSwTLxCOPYAbMiugFlRPFw/Fx61
anwLWvX5xO6DiJGQhjyOKOld/hEIS6Ma9OWIcswvyUz401sU/zyPcNUBpEQ47lws
gGxxbfUZg7KKVXfqybt3JTD5ipUHuNNOJl+DHauPU3m98bRIFoBfE/1n0f9wNMuC
CtNtl9FqolgqBI92SYeIpAAz013rAy6NK+RxWA3VyjF/3pViGFSCci2iCgXlhcUO
JnGMcKGEpEYE1PqzUbGhqrUQ6ZpF4UVDwG9xCpjWPgXHRxsh0o4GSjje2S4DpOr5
NxBD1MSFydclqjf18IRQZNEMrp/nbpQDyYTqCALUnQXJvl+8VYlHDu1Zr+hd9mIB
0ypPLjSGRAPhOwalFLOEVv05/iqC8IjcYZWA6/SHf0DB7s6sDNGjNhxwejzyilxP
zPAaGtkDBhpK3SPV6aC9Q7NQwnHaMVzgBCuezCZ0VM0+/i+c5SvQ24YFzj2hUu3q
Qv4AkCbjNa85h19pIzIesOYlzm8ZZmJPI/G5aZOqvAtwQDuvZKjPTTEBPSzxQtj2
SA3xJdbugrBZFBI1yxYhQm8jUJViYTU1+CjdjqyCT3Mrb9PrpKU3Vh1mHqGV+0XV
+7ZAXtIZcMV8PVN8S/OZizUUGWC2OkJrKg5qO1mkhbl16rczOQu8JBgBrbllHg+2
uFufykonZoAMcOGAg8R7DtskAxY1fRq8NBKdYfopfgm+N14KzyN0s/ouv3vR/pvJ
vg1G2W4mmL261weZfnd47w6pOfx+i1dH7rNmdq7unML1kFSjbRpYKpfwrkHAjBrW
8qr4EdJy6/e7E80louiclD3tJdRgdnFH7AhhjN7P1CP+i5t4LCIshvZJONT7czql
3NyQopqComT/1Si4PNdLhajYzXO3uXrcVZfH/Dw2L/UscL7WZdAcr4hCgvKKtByn
M4ljGP2l+TsuB9T1IXVgTKYfCNvXbqY+Mm+lXgeo0qq3a//pOloey+ISoYdUZeC0
MKng/D2LtrrD7usZTcjXWofLgymL81Rc85bT1cEakHZ/ItceK8KXNzz+3OPu6wn4
4cBrbiEUN/DGxL8WGDhWyjgiKo/FV+oCl0UxnMHrZfijvuTOv3a73m1TypC1QuYf
CpqgxsD8nL13B/EiN10qECKYef1aFpxZLZw6yHtiG315YKP9BRzDK5ftffPpeDvp
+KVGDwAIoneR/wADT/ZnSMZ4h+hBHqNGBi2gz2ijWJdL2OrdJjj25E7a2BkVY4wJ
U8ZS5Y32djSwcAJVzJzt/nCXwzN/W18OJS9Gjzt2pWS0IoFX45k/V+hwQ2cbsKFx
B+ETMtm9VJ6QHSM7zt8Fuh/Kb5vVKYSCGcGIhVhoxwYmf8WJEEDxulMpxsZQ4tQH
FqVIjdGaBeFuT5492HOP/UGCdJUaIfrCQTtrO+XFX1FnNGECQZgu0Xg6WzdTYuEx
WXBGzEQHfcdhufdV71B9sFiQ+oTH6JtqNmOKY+6yzkDb3qL4slfRokzpcH41KrwU
2jg5Kvqemwnx6PGIWlnHIxqEyjCGzrmNgnqWn9MIAUAJ0tB28XgCtGDas+ola6R7
QDPRHU0ZiwjVufOmVqEI6AHryc1Xlwuzft1PKoBlU5JvUCNCpHrK1+gZTs/ADvDy
naAJylAAc3sNInBRicIsvzLP896AQ8p/73w24J60HTVeNysh6roFFjO0quSRGHrd
45hYmrv+X31kzhSLpkLO/SNdWoCv7+N/iEASViz7p2Npa1taD8ATBnLxDFk6Jp5E
ZMasVMVZCjYKdcoP/yvZ10wHZw9PCplx0Xw01CN9AJBW0L7LrrI/ubGJO+L16y79
uIvUoLf1s4wz/kwyq8fDoWRz9ZK7e1LlVl8ODhdc8/ywASkHvEqXSxfqZ5NUNTbt
3OCGk5/Wis8/ulwm4fv2gMTZNyEVN6765eK43GO+B4bHNRI0KHEIlzpC8v8HTaIu
0leK8rREjWV6rkebgYv4mtXt9wjiprTrNiLsrP+YSmZq3e0Gy4gK6Btoxl/Nby+X
A4nzgMJ4GPhQn+wr8bPUTOXWKP8QtgXf6tZYHK8UUJlBeXUbkP1AkKl414CUWdan
Por8mgt/g0lQz6rpmkearOc6O/nw/ov0QpaFzMVjponaKkhUmDh9G/yMly+1IVzr
oaA8stPNMJMa10S298qwsRXRqQSMrMOzkSaquHc+DzFVB3b1vsK30pcH7GB+r3ef
4Y7UP8Hl8Mt736YVEK4hF0V/UVLQx2z6dz+/CoO7NmaDq0UMMN67J4vbTNCVCZz8
xseYQNNxX9hHYSj1THxUfg9qleAYgdE4DN9tfpP3uAk9DGsxbAKT+mdJyfhnQzLa
JjLsgDel3kF9dOnM8wGuW67tHrcNBmJdZAyuILLf6ksc0uwbXNyxnHBg67AsrERv
0Vf2Q5cqlGXIsiBIsj9SlV6goo1NZ5RtDwvyP32INZ5/AcHYQpmfiS3523U8OVGd
870cXvng47CDGLk17K8KoEQCyheqd+n72dJ+C5Nm3+x5uU7PKvwlj0dRswA1UA3t
qLac4hIVIUxIFhRETSlITpxV5BQDRAD+cuN3xmij9NsQvvAcdYaXs1WQoo2OYHxZ
lWcbj7jWU0VL/F3Kye/nLj2tyNo5n986VY07840kbNtlRJ3dT1BiWzLcmWLjyljs
TWCNwA8U6ez0s7eMd9iQaBEYRuP7KziyWR+JOG5MGrjvsdKKZ8shBbF5cK7BnT3L
NoS51a2+EqRKNhFyOCPvuGy12EKEIKcSmCTgZu8YK8S0bGqJDSpl/8ZmbQBIdqal
y/Am/fAQ/g1W/YkZo6TRLamux6AZkTm6hkTx6L6eBywsPrwoN4N60pqbkdpkkzAl
sPtBGYEsJUL+zy+cDKFZDzGYc7UTE3OZ+KW8pBitWIxOKCQnvJA3chAkx9JDhpWe
fXucFDz9SsYR50fqItvFio2W35NLIGjg0XPnlDbGand3zQEYwtuq6/47zzCS5m01
iaDikIbjQSYwWD/WM5gdkzdPe0iUXbKtoVp60ThEY/cs7cWokOREZIe7zDXwuG45
VtsrpdHx7oxANBabyYY8OxYqnrU5Xgp3FLdJXhxoLsstxjqc7fmePg7ONlxE0ekU
ZAm/YM/BqxZx6D9rImTsbAsvlb7MHLN8P1ZLNcucciDxBkfngLbo8Z/dKdEW9Uhi
I+ctVxo89rdibOycSAzpyQ57IO2GUiK45nS1n96p34QQt6+VtPVdY5nrVfmyAWH3
hQOeacHySsW3WtlUl3YUOA9zyvX/SBxHTam+BbEHGSi1+tJ6L1nU9KGZWmbAponO
Ijwsmnv1Ar5agy6iVPF3E+e4Pqm8QtAxiqo/Ldtn1AURDf+jsSe3AVoXRtxd+6Gf
5Q8I36JKqwxAPDwr7QXQvE6q1Vd2WSfclkzZkh6IOAZug47zu0qLdvsLNgdiMFtO
/SofkPaYmp0iii0udx76LldY9rqSp1pRFdMjJV+LOJVajjGksI5eKTNekhZ5wgEW
aWgdcozfreOQ3Arefz/1H9GDMwvwhxRbFY4+e/eBT1aBtWEWJMybiw5kTssQSzRn
TQc3H80/YuWd33SXMp+ZfJEoZcHWDOh2rZLNn6hafw8YoZJUuSKZLOvav9LqfqwB
XT9aKG9JSXDM8HS7kKVuAKHWuZ0LMiVW6MeQR89yIjiao4Y+8o9vryziJKLlSK4e
7xOg5TCTUfrK8btLa2kMVtxwAgrKTZbAwBEsPrpF1IQIVn6IO9fL7rV42I73+dYR
rs6tiOqUBR657DEcOoCPhKLdnTMpO3Jh5kY8klEi9tcfL1ZYtUOWKtuqH1YIpi7H
wqXfRDLNlM1CjONFaailARR7Y29heHby+0ZlTbe4aFC0ri8S3yE9psQlDX1T0XIf
BM7cGVFEcJG47FgybU6GolnYjtfTPSKb60Op+H4R2tMBed8rQVuUvzL7zqoOsWqP
kv37sIgYjWjSmBGyx7S6pOQri8HzLW+613IEciIonN/6IOsyPLdekTwWz02mZgsr
pNOZPSJY9hEfc+GCzMlTWsO5HsBlxPptj/XkJavrJoqxCDQgBjW5xO0e7xvAJK83
WfhpHWMUuoX0pBwtzinx8Ny+/rmghEA1nxCZ3pOP9Sq8nR5QpCbLUfPS6/F+SoD7
wUe4xgdkMgrdcXeqOY5OzVMJeV1fH6vkZnch3nK3V3w8oBRi6TO2g6ZIfpqvUAMy
hHJThWdlI2CY3bAPgk0tZNcRAwzaCk+BTUBnjUavSJa95LQMZpkrcNClF0jLNIjC
GDzeV+GMq1XycBEebpNe82PvDFcS3Q2v+cgGCpzdi+ijesqwiM9DA5OkzSqS8te4
8Kirn96dKdz2kwhWanlaUdXOw+O48cgrXJlCeVvJ+QzFwLE0l35HrOJnyXVZ2X/j
baurLId5pvcEST/3ydaJbAaHCoZ8EmpFa0Gm8QO+WLzYvzYp6JIEjnJnmaVfcxUj
O3Ck/LqzrzCY8bM5hu2Hq1QjTK6WmI3aSEypSa3HrN97ipwEFyaciSxYlF9Y9Ti2
Stiw1GHiL4L9LjMMBfeFn3PuSq4dg4KR1yuZPgZxjcFT23ALOd8fZg1mk+H5utEF
WLZnBaCvSlB/aY3lFtpehPBAD3D8+zhXCPxbzHlxKxUJFllIxYqoMaKHQiy0Ra+X
9KWGH7Al1Ut9qGI9nYahF7Q3DSDYkplXeMvIy0ErEJv1tU0rR9uNT4SygPqx8J9W
IeYUrMXCQTwd0HCI6W/OFc24TYU2c6b++Kz6wAa27+9jI6pWD35owgl1mcKgE7xS
bTrjRkQg59VOj/y0zpXVW06OMPNXOBKaA/u0Y2vs7v8CYqGj+OWqCYSxy6OLQ8Ha
lxFbzaqEIJCcHeOcb8vnG1Yt/EJOa/Cs4dNBbvVuVLHzCaBjQK1pw3XfKjUYcEET
iKqiFrnQA3X/HdbNQOOV2HRS4LthunUccQDW4+tHzzM5UKQWeDgNLLAf+69Otc4F
+fMpXAjG1NDUeJHatsA0+v918LGzGd7eUBlFNeliGmRyHXU6HaGQK15Cao7oT+cv
NzA0UfNrkRfCYkwKjES9zSpwyI/fR/0MTYHQfsc31yi6x/q/pTKdKnq+B7E47Aru
CX0F9UU3muly3o4GelXBbV7v0kU1qigITD18xqGU7wdG8ozyJ0YMIdTGp3H2P+1C
odqgA/Ednc2JnyfeulmvV2LSmE7NVbHdSFjV7cXnr0pP9NM3R8/RMEyIscg1gPBb
I4UrfaeLrxDIWO5h1xcJpOoUSUTMQf/llQqRy2Go2Rb+KqnnWjehfidYMGpa8SeF
7z8/Ms2NxTHai6NLX/erlnm+obIfgNO5i/6QLSd5cKqhAuf0Qnny/SqrviZzx1iC
L92u+aWb6V7RkGtMQmMo17z8YEtDj4g9tEKwGLFdH4rK9UjvDSJraEHSbH5CFK53
s6G4bhoa4lyanbfFUHyeHr1vhq86DLQDGuPZdoqkRNtFS7CQ0cpQKuJrF25DVRsP
leVZ+Io2F2HbLOyZvysronXnF3cfjHJ3/0WuGOPA2K3CY/MrSiVkBTrcP236aSgD
PzEDF7ilFsBaOJTjUTMWyFCpRhRbV9wzjmqowtcd85yBxD/XLjxBuet0z5mFtAcm
v/q/h9/QJ+E75qXKUIecTykWdVUZpJ63qCq333+6b0kQ94DPcdbmjambn6Q/NsmL
gwrjP0xo/3auEKN7TJNb5U6fvjLx/zoxdfHBPw0uBdntzaogF6TfL+vdID8LSy3B
anHtBcoEXBuJZ24TlVARYNs79ihpkXyrW1hYEjDsml8VEOnuD9Ip5A9Ub67iz0dW
nJeU1FjIUZaNlsTy+5ncpZrtSOnXwf5vFgrNOByCzmA9fVvdGhcjrbiwBkhpNCKx
C+Yo0MdwxdQQ1O8P0Wl1sP8hHKTvK2zElSPoQ2K+6aRaPzC1Jq0ARD8RJ0k2drvM
QtlotNeYipUB6QW821YQVUfBnXKge8ZdibPWAlfJzJBsZTbmGCXxb73C/xnVbqGH
SIXP/6BC/kwJAmjyWJp8H7F3wASfKPF6xQYggVBMVyzUbNYyKhj78b7XqGpy6H+Q
9k3WMCj+j0hmoeha8fsKRRtDektWW4WI98d4556MDeY9lm8tOJJtjMaYLUk8Smm7
Up+psrUjBHpmUGn0p4Ub79JSPJsvytOy6kUJyCEnYNA0A2MuVowYuQo5zjiIEKKl
mnVVhhhYEl3n5ciEDeevKDmUkhV5iM3OVXWUrP7775aXOl21quUUpNA4bk3fTPx9
tJ92lU6+kzoEo3j+6++2bLucpsFguwOznzd0+HtubIEdN8YhDzO80OPF3yTsIpYj
dw51NrzI1j4eHCykuRGp+/838GJQ/jPYh4P4MQ0ffQi8t0xp+TuUbL80Fhv7qpIB
mRugQLjST/479I/1FkypO2tfyyI++uGGar235tod7FrLv/xVBgqMVnl1Te+exEzP
5LkEiWyBx1GM+fVmzc/Wv2pgyRTlqJgyEPDrXF2v1y4p00LNS/+ZPzZv+lkbUVya
NKCqfieRtPRkUA1aLZlLQUNFOHpHMpG/XtKsiPOhkkTt0wnij3cvOXt2Gvv9VVXu
RUWOv6LN5EOyiSpgDYA0FC44+soH8eh3RBXiGLVzog+HEL0gyA/XflxtJwPdn7vi
qTbOsdLG5X70crUHQwAqk//qoeZCSxpY2S5pOrFvlTV2XhTwVCfVIV7gGBL6HdHs
UVAAYXWndWSBYIPzJwJeYntLmdDtqq11uRDUiomueJ95vhaAhyxVLJQbivXpqfM6
ZX6k+nJ6wl2NX5rouFBgLt8GryrirnMJs+MpVG42rnjrEH1YFeRQmLdSc9r3eocC
UkGl4u5frmvWhnbzlobkIc58DjsQc1Hig2Fnu7x0Posh10vK/Ud0vThytZzmYl1M
Tb966DMYaxGToT9ij0Wf1C5Z+xqqy103sDCEvkcEzTlQHxKiUJEtuXfFFaAlcold
5OclkoaYuSGQJZRut9hgp6GCWmSu639RY2CvGX7IGc8rfULkHqbfVgZWOQMSgc0i
AlYEbQEl1il9l82c0YrREOyojwaqzVGnR4eIEPGFv7Wbm4VD2asahLn3R3fUaMTK
UELMnCz2Oi0rLKzwY1cCzZXyd9T6AOm8ESbtot2ckIstjVnH9zqwt3MBOJiymNZ8
ak/t+gjk/avKlea3jnrXh9KHlP8T39ENHEylaeOq5lSxtQMuYh3nR0+muBMj25t1
hlN6QELBIwcqgPvQNQsGgyN4gDZz0Ya2u/SSHjuqnRxODLdpL/y92KDMKCievv/K
o/tdAQriTLMmaZU9L1RGeLn5aHhjwjyvslfXrV8WTiOdBBME/Ahoi0y4QTr3n3Mx
XvJ8GbVyz1f8dqyQqkUEZWOX5UGtif5qJG/vFZF9IsvOPi6KqUwzEcxDScMeXztE
9JdrNHAYZ8Two7kAUTfhM0WDC58bZ2K/mOKWcmJiswspI0lahGQojwsOWnRIywox
iYJQBPILHRKKl00aJXDTpviKeRZvuZhTKLS1DT7ggrgjcqVhcnr3oTz5co6KVtYy
8sdI2nZrQ2O7vYv01yMndqM7pX3tK9L7JvkvN0KYyeuOWs/KUFh+epOxnInEnXNT
tWu8L34k47pXWOZBjgxdhynba/wXzFk90rCBseyD1SeIoWSMlg6yuBR9ytJfM2Hf
sh4DacRADRy4Kqt+YHjQ1ygX2h+2TFujUgCsQo2lbVES6aXa10syDDCAUnZdImWu
vTNw06p5F++W4eHNU7cS1exoNSTkA5YZKtc0GRUBzT5/5n5htqfW+AxTgEBqAJzm
wLAanlAWb+ktT661hrN6sNDIXkqkPt2RM72L0JC3uJbMfOyp0s/hjsG9bnJ+HZM+
0sA1OPw065ktlBsiyEQiGdUUzP1RxOoy5Swm1GK4eRAmkF+TV1KmeDh3yMeEbD7j
06yJhhVTMJVHrAq69E+cLhDM0sTt+hbxJjzcfgNIE88XIO95iUJMJeTpmkndERQc
lQffhgUv5F4VBAmihbq6Il5euN2GmRUFejKT5iGhiGAUjCTzpJPgMH83KuLPc4QZ
2eQIQixDKbJRsgCWjSiFpAGlqMpY8PNURdok5kVtmPTpxLbx8mR3JtO/81uAJnuy
flHhVkhKY+XZJmtV1x4rOOwPZ5ZR249paYTOL0xE5tdED//C/iBBXCzjtkq/0qQo
vilEZvU6S0oD2jA3PyL9HZpbREhpY6n3QSWuKX7ta7r3rwXwbljQzv6bB0BOJtJl
Xn1VuxoNVVAuebUZZzJLrgiWO7jS/ns79XkIIYTsQhSVhMq8wm2oStUfgTxqbk1A
RZb0CUjDjAzu2jE+CgUvXpcXEqZq2VBi7Anc9YuWA7rZWreZCIPcWmA+RKmxrRZe
JgZRVAZUPkW5jJlod0IS1fYW3D78rDvOKSBDBiH7q0jPWI13qZHtRPkmghOztO35
vpqaVvKx3EzhZKoQroI4qyY27La0jjz33tJ7ofToeZg+yRi2OKwykgp5f5dUJNIf
Eh527kdWJs0jvlWhVqL70bd+/Nz1rzw6+g2ajSW+JKYlsCTvgqM+Upvt7OCjFSrC
fQa1Q+4cxV1UMkvSUy9VnT7e4RuH8BO6rzDPCdIUNXKKm6EEcM9TtOOKOrARxxxh
7rBY9Uz0tO+xaWpZtPS3wAaLUCv6ZVPP0/Sqncyxo8J01vuXo/dn6V2hn7nKPjzk
sdcMN5VByL/svElfgwQlyk7a8/goZINbznM1JZh63/bIx4EsMt3uPnveMAKpdMyK
P/GDqdTMxfwq3817BH0KXj6YuokY7loJVUpIBHIRJARokcoLu8faxggY1GCalgmF
UFITRl7SUqBJ98q0lUrK815bG96BiGBC8tydGpAGH8jSWsAmxzK2Woc46cvEYoxn
hw3F7JOnrpAjKVK7J3lKrcS6yV+Y3sFvBF3vlIUt6uD7d+/XCfreXQx4Nyo3GxAk
75c/hFI+YzrmzLSEBlC32+9lYbJJqib3VJoS2U+eMqDiuns1fSlX6i9UNlFChixs
5uKRRYSivO+Mr5Ju2bLhkJ8M2uhyYz511MhFdK5iWv0RrFdvIoenasRnAsXF6Nqz
sYanoaXVYIK8zOaXKcQUcmePesazQlK5fkR8gRL+lzIzyCzbs3ri+DFrDGayU5Ef
rwCmGTiTkoXnlgeZxTEBpHzCKVXXvsvSP2pO9IjLEUewzNzO6iLQQVFWJXkEZoTC
yCUeq7l4RBpID2Im2sd+gfCdHaaCKIbeWnCp682JsKOgT8/Sn207fE7ElwBSK0Bo
pFuPRc8Xt8DquWZ+SGCbuOzMdm99hIm/O4DdkM8ZLLl/Z6bS1QQb2OU9ol02seyD
yY/9vnF57yM0WP54NmBHgAWZFIeYjdzg+Gx9EHVRNqtMPgE2bVMzn7ZRdNSlCbPK
VTzYTBedTc0IJRcYmbu58NpPhTGeiKqoxM0ksoqBRtEDiPUerz9bsEyBDPq6Pmnu
Ia8kKGRQauVhnhJmtBVqJ96CiU2+NsfldMlPm0pUJ165SW8T2jOpO1FH6onlv4no
7l6TijJh/pbXiDilxrjCjBl2U+d7/sKGVKhPzJZ+sFyQecnOpSBWh0XTYUYPWpnY
hC9WAH+1xyGOKGWIB5U/lTRh2J8Z+ebHZ2kvNoytp9FQ6Unvs4F5PcVMm4JmEsYQ
ZBt9bN/zyjULcpCariRfeU4rmYIBVkzfCJoj2IOpV7o070LNU3IFp6y4aXU3d7h2
nUojr81U1+OZjnVcm2vwBDLXuSZFkbUco9pdegQKyTrsBBLykYFzN1dqY1TCRGGw
HnpQEAscWJJmK9BU2E/mHp1OSuSGbTg1d+QwkMN8OVpOrEL5xoy/4P3Ewo6zjv1n
64H97pMSHHSK/iKL58GwLXmh5EXb+S8WiO6qcYFkpmyD5HxbllOzSR0Qajtfjwcc
blo/n550LmUl05j7LRSO+oS242KlQ1gUqlHV9W54wNuOSzQ/tX5dfrSFF69SoOy6
IfiA0KRrggV9BpW8X0qq9BuXRfskfR6+JNQwwZYO/zGMOUrR/VT7nZx+U9e9fONK
hcNWrnVlffKf9lv2Mgw8Vv8DN5JRYZbG6CE8vlMxUCfK0Cdfrs71Df2/sj7gs3l4
nikTCmcf5Vyp1x5bh/ezIesyRnyYQwQW9c7aKcF/Wu4DOIykNOz38hx/pRTAs5Gx
HxtLSun33KLfBRd1le2jzukGZXNd8KIREbCnomixuB96Q3a+JPP7Vw+wY8DkKqZ3
I6WR+T5o8oFdwR/87/NGnHpFIUmq5LnmdzO0noGwnJutBFq2lw2qwWiMJyJxl4Tx
UkYt1uj9v0VeIt41oO69K0Bi3ps/zp+GB3/s7S8OC51Q+HG+viGBQzaTcOFx1jiA
9h0EvrNyEvx5+1hb87oW2TB30iA/x4Iwri7rsqZPaPlAwqL//NGypCYLFYxPJt+A
Z/t6OckhBnwL3wzRqwZ0FRZiz6GDzH6+QZbMtTLInDHbbZDajn9TN6l2rmjAe3N8
9kI3qtT7WtUN/yB89V6KYG3ABWJ4tbeowww/q8hrwO3a4axZGKGKCZ9Raq4/iysi
penTm+eHAys1w8dTLmBEjr0eiMhUSVUrADVTRXv9UxzJyHvladR9g8M73sN38Lky
AoHJ1l/ocHFbCxxUUUuBnes6fjQM7NxMmyFVn24LyXtsrgYTgsrtzjOjzdbwP2/0
gyuHHDPt9Hj/7jpBmFyHhDgcoWsCZ7DqfBsw0G+2ew8vjtxFEXak2aZVNZaprc+7
PvAvET0vMGnboFvsDtCevM3ExQqjrc26IWw8vACaWmX68oqDP/XHygn7ngbpbqxD
L+Ek7sdBJsjJMz/siNagvOG7IEhEq59sH7Ks1hU1tP25y85tU2C3lxdbvYZZ2Ttk
dknR+NcJmkIX5vXvRFRR7SR+59EFwDxOjejcT3URvHI9KjIreWpuabZwkMqXk6bZ
9D2PjIwOPlDn1KrsvVSIo9CXPL+o9umEANP/OBPIfugT+VgpLs0lIZG/WdUQib0I
e9+ryl/QXBwbqJl4exlt7Jfe043AhAuhndmOXjhSD6x7QHriCYhIuSTpxg+GslMv
Ru6cQltt52iQUuL2ON6knf6UH20R7h2jWkH5TLRIjN5kxCUhIrJQkfBvMMMjYehz
we1Ghefe7WjhCqWURA/xbUCTt7MGSZ2+tJKEaoDh55s5nEGspJZXC9RbqWqK54Lx
XAhiOsto7nGPxYJPCqPaPReWotSVr/m1VqBqTwD64c3eAl13yVu/qyfzPBMiAyeT
c3ZOfk/Mucwvii/3YCyvB87VKG/ZMrkBDSaE7jjFdpighfeeHgJ43ltoz3cQ7aHs
vCZtCecXE/9KiW1/frW6bxgkCQPIaWKduQppT50JRdTyKLPO/FGSYiJG/i6tWJHt
TFcUKPjCngXx8GRrm4VzlKTMWQh6yLB3xpXRLQ87R9YYbpXRIF8oh2cO4Pk8wTIm
ZZWnh2qA/wTWSyZhtjlYLmfFgwr794TnZCgvNCyCL/Yrl8MCaEiwmu3ZQROlDgl2
wTMSO3HSSke+a7UGs+C/DMTCoZMV5Uz+iXdD3bDSJahKGvFzj0zWG6r6dxjF+R2J
sa+B8r4ATovxDOYvUk/7U/6Pb4i1jvD/bkrz32U4/fN/yPlGIxSbsof007EuwjhB
zV9/V1VkRlTAaCXlgm9z98duXKLfBu2LPLA/O6He/WV+ojWFPf2fDJ6b06Pl5FCe
ajtVqGXeJ/GvCaI5gRS2PWWCfuGmPhACfCe8zI33N0h0nF2QbfpxBmj0FDdWhi28
yVuzfOwIenqrxYL+GjeCKQb9Ous1gcdo4RfUJgWgjGyIsfsIP32QPntuaYzEdIgM
mlV5WFgmjyZd7kuVwrINDQvVqXAiBDgM8GEYOy5NvyYH71vCUbpCyVyxPKPZ3dJG
ZzgDMjHk3eoPY7deNE4SRhktI4WXKSiK/fkQjNa1/0lyuXYbB8y9BBE9wrNeZylg
R2FZAx0WVkDr/4O2RRuG2+s00rfc8avEqP7BMRR4PW0PGQALqmKBziVrWIt8gkM9
EKSgaeFyroCFPoLNssB7UOlT9fd5duvQmJMf0nFhV76WHv7LOqZxRajAeEG3E6AL
newiWmIxQEez2lNl6j002De68LvhsRmyZHrQoGBGbU8RYE286QDT8wqB85JP+xt3
v9AmkJAy8HzeXKWffSg2dcySNGjxLCLs7EwmKMYRAE43CrFP6j9Mk/fDb0rK1RRO
8LMTGX7HGXuG2Ev+UNUDl6dJpOezrRwWIHP5VpO7twVNQXRz4ZVwqYCADQFty2fS
EdryRnhLQ1U98hGn7SzHAzJ8zIxZ68vQwnHXcmPiX/JJii2+ipPJsfJ0wGl8l/8s
uf2cB14noQ2Lb1MQWITHvXntwI33ti7WHcsmi6u6BlcL/FRQvoKpGYyglE5pNBTT
VgiiqoeJODjpMBOhUlbakGuafO8rWWmpMZjD6n/6Doj7ySadK4ir44hkvmPjUbxR
OvQUKe7cCV6pY+7I7J0DXT5sfyjdBu1CKxmImjOobW5oRVgZi14/F/1COSflvCok
1t6GDDzBpwVWAoE4W5RBms1ETpUbGSuhgy6FKJy4QpFkSnJVjqwbJQnr6e6z1Gk5
3L+zCy3Ynz4ExTu0FQ1ENuC9kEuaD8VxgT09MRXHyEURx1t20e096e0JkfIAwYWa
EPusGKnuQQjffbUCrcS8qRdPNcwTRnDWbjVR/QBapMaCtawn1C3ESgnCnacmIMvQ
ymi6AtCTBjGnG3k8c+8U1NVWP8UBmMBcSnn+mjzrJUL7PFizRx8fow0REICq5QX1
9lJepkG0YtoZwTlNt/J3FJAXG0pNL6NBF/+9efez+0AYCxbFDrJLnQnDWUaFY8ON
Jh08z7q7H6s9cRnzNVy3k/pUZUNCuhxBNigqFzR5R9BR9GiPI5Y2aHt9fS4dIaZD
6+Ys7582yRetWPNQyPxqzwN4k56CRwi9o/zoPRnBTEKaZdYeKXVWUxv9LmBbUuKw
+/XjjC340Pd6xU0Fy9DUkhhEiYrYruTgn/VkLTbBJpeG7vpQMzu5edEdRjkbxIC6
mO2thgZp0Ld7dzZCYLKkjBt/wIAK1Km6K1dQQn0Ze62CF8pleMKjJ0jav3fMlTQM
wnCaFxUhUSyc2BHj5lJRnkZh5kWzCI2NMfcN+A8/eJ/EQW/2qKLUP6uZlYkGHTXJ
PopqoSpPRXnxuncM8+XihiAO+VQ6YftDvCL69kgyiyCAcpaMzmkU2AzIvbl/u/rT
xFl4+hdMr3tS94Dm7uVDIMCN7GsyjPyrTteTKe2yIHtKSzK+dfWmJlPSaNYuRFGv
6NQ5fs4v7ZFr0Ln5z+paeVnHgI1s66l0hee5aMnWtCo3KBnmUXUdOs5Wl3koze0V
cOO75yUBaZBZAcMj7z+0bCJeS1zjwRpf+XnvsXNjSite7sBIj+NuHKb8jYgdkWb4
sp6J69kjVCZVFG2KqpMVoaP5vbAk2mTc0wqztTdAKYWqKFKM2EVL0m/bYuWrafoZ
nfHyM5djfWoQO4JfNgjRVobZZ4x54lSEl9nECehGSqFxPfdFOo4q+X2zd+toq87f
SPh8lA5yGHY5P0Rp2k1artUFhlHKKzsF/PgtFZavzXb1VnroZTEzbPIL7Zti4A8F
M88NOY6trLxhn7ahO0Hxp9GrZ3GxyNcLOyLHfUWGQ65+Te02LN7xD+tWLhp41Ys+
P4GZXHYfr/yyo6O/yExHFBdVAlWagldqGN6VRXOEguJvbkTOhMYqg8cu1YuNedvd
hS02vT/gp5gJf5H87uDz3JVEJcraDrIgefV+x7rEDjiA6UtkpGPdPPHHO2wfVR9j
uFMyOSk/8qfA8EkO5o+PJr2xZ1vRVAkCbtOnfgRQLLQ3ogjzdoWP/F23K4ETnbba
R5FQPSNpAncCFAmPhfTJLMwC45TKNrlndhC026ToqD4SGlcUKgFYTfUoPL9x6HS/
fvJvQ+QjSV+dtejSeDtxWfqRysbJRLHZwV5Soajdr9K2m3A+V+OLCGeAuojxIXC/
Cn2O2Ehvf1XzpysGCjiuckdd043fj6aWCL8sMT0sNwEXNwOkAoqZwNxupVGP78V/
i7adsF23OLIBnkxXo88/3QhxlpD1xPtJc7nNNcNi3ED4RgKPnZEptJsI/uBF0+65
7R9lADVhsaph0+kNXFhBg7OBsM044pTWkhGZiSKXsIrSKU5SU5wLyh9tH7HRCyZ7
QATN7AwPdKhpLcxyHZzkHjEjI7fco+wgg0Kwwcvbp+6oIRPWfMgluCiT6MPaWOpo
owba0AK8ofZkhxX9/gDyYDX8Eb7cGYMz2Rj+9tgHUHGCbUciUg9DacJPyDMutEEj
AP+tOzJO4vBthpl+TCH+lseirO31mPjd3kJIGPs7kjQomR7mHSML5XExqb1wId0H
yazVpMM8FNQXvExZBiDgfuCFYR9XwWv7KbBWlPIsR+jXEtXhXG5DvIJiMwvgE+wk
oGPdwwrYTr60iYTR0CQJyi2RBA+G3Aas6mghGJRH5Z7IMXkEhwSmE51tGUnGHhzq
L5wGgSmzXbOnojpWN5TouIY7MLSmSCWg4ncIJQfvgKW6HOq5utulhW/m2+s3Yzv+
hy4smmv872+gLm/M76LvzsiFsIhuxoIhJcpov+ppSdmHtorEe0EdK1NmPvgRGp+D
hu7ofRN0X8ELuK91RyyRgl0cRntS510i8BKmG5nQYm1g1tz3P8KldDgkQCi71zQU
3txCaokxAcmLAkET+usUxKQyvJOy1VwQ/ow/vvRHethR887gs48/dU5qIsOOOogo
08hrbyBrAPsRS4HRzyItDNqufz25xokE66fge1aUnjOezbxFGQjjLgwjqHt/kbg7
PBrLhcKyOZKcV5FNsRPncy06/AQ0ku9WVbVuHyi7MyAsoEgzF4ZQXhl0TWZ66JaS
hxBo29g/ZASO2s820dscmWkv0VNvLSeiJshPFfmqmnsFp56tTMRZ8mjyTmjz3mvk
xrNgxnf+x1YfuupF3CNh6kbUwTeDrmfcuBw7skT2Aq0vUWiXI/OWCN9kvPZoohal
8G7J36d06s69sTvGESmJAK0+ZTsxh6w5RkiquAqYgkS3bqoio05B+xAHE7NkNgY7
JbgbOeC/8TwK4RpYK7tWuowEWc3uEuc+vEsw1dYPICB8nhtuO65Ywl2GRMkBQqWI
iuDg7DWZtd5ClxmRptYyFcacp4WxyeDLH0gWIyfQPJIZPImfI3ijzS42ZkfbPtga
6X+NqiZvd1NlpX0RknaKoq2FHiCs8CTtF4xGygYvkvY/dZtCsOFqUskmnLWAH0U7
ZRw5N/7xY8uvywwm+EMpziwYQmMTSRA9q7HKyQA8NM3fznVls+vwjjcZH6P9nz7I
r5fzCcA08olu9y+7rNHmTenayZJDj8aNk5i7v62BKqEiOk/sJ3yWZ4SJanweNgRR
+vY60DHPo461Gs3l4xqfR0e0V7+p1RSszI9AlZr71nMDESAHHNIe7LY0YNgbY9BR
GbY5sIwjeoJ1WHXGm/4VE1csKBmYG22WItyXDx50k97Ow7C+dVvOWoYxJe9gbchs
RM8alkhIIYgORVdZ60zLkT/4naN7++484vknXeTZ/b7W2naBfou1NIl9/REeDbFG
YTYtdn29Avp6mVR7BpXUEccH8altP4ccXZUZc8PJk3Z02tA/uqLpMkrsd2fw20sZ
7u5a+xvNHOxH3YKyM160HcMzX45TFCLoUuirTJv78MN5jLrrMe6SyLzVEevsITG7
6KA/GguPfRLQ2NVn2R+j6RcaVsaAMJR1LelKjiSs83JI7Msuu72y1uM0VLoDMnTK
Jw/rjE32wzQ1PgWyvuX8fzwhhTHteyc78c3XE0L/FsdwuudJpzpP53Q0dF2PWNLD
gYJ6lIhxoQpV3YrGZgsGIBUBNpMUbePWwYZCjrlRlVTVgq/cCL+IPIEE6WJoPT7K
eF79g7Hj2WJp47o/0Hs8PHbxl/qYVt/Zam+ktkXt7Mf60V48V+VSFp7h6lkdvZz8
7sqRVONGlOsZf6jPyguFjN/2Elj0FO5Jt2JhGaLOsmEcnsLBJjiY8DB7kEMWbWWj
aip8D9UQnlwKhEA5GHKmvWsDRJ+CKORGFxINAHL05eaV5cLdsJBe8TanJXUVO0sz
1oi31dJ7rpAHddyGx8u3xKaMSRam62DcoumVRyy1rVsWNUziHYKyhAsedJzMwJTx
TCsN2mjszVhwnvUkAOMwIYMMcXhN3L94IAhwEbt/7yiX6/hq7e2AZw8w7EdKon2L
Wx3Xj1iyDEhIIrNrqdRxDKKqQ9osra5ocUO4r17X3f5125nqcgL6eo0SUsfQyPpM
+y+Cj3Nj2EPCEOIPccodzmE3GL0Q7w0WIrCl9i79LJK6zMXx9Va2nOO7g50U2cQa
CIdxwgpur08CAkJxv1exGpeq9Ttzjt91glXNi1UJBbAlgNi2rF0QixaWnJ3bqQkP
AyOdvxaGzCM113TXp60WRwq9DhVv+3kdJC5TSgE8ThJjoC/jgckHemP2hmnky6bI
fKKBXaiLDAihSMx+Zvc+EMfZE842b86qMw9U5g0avzvxTslNO/Fh1T1prpLwI1Yc
JVzUH9At1+ROyvCRa4420FGAfIofcQmSEsNjXwi+BNOGlVOt/f/iff6LTRk2P4XI
rohQ4kkFLz0uG0AmZXmcRiQFJH2OjX9rfpJ/IvBpixydvUsJiF2GM3Pn7xio7xTo
RczTOHaLzVRIAufEsPzPNkKZ3tBX6cinoHKcTzg6fNvQBn5DnNIDgNCo6dyvomt/
dSzhhFuN9UPujN4gJfX/Jl45pEAUves8Fe9N906FkeFVWKpjlIlcArclEgSiViEg
+p8u/uLyHoldxBKlI5cbGG8HMkqSD2IE1yykBYfPANOr/p5J1J9LULEAqDY/9myq
7+EFxub0Toc7c5GXgLPFhvSf3zxdQI3IAuV8oZjXwHWtybjm+3LKPGq34CiSXXBi
59x82EqGE2f4zQHIgiM2AelzBquozE9cYJyfsCNWBawz0KJ8zd1AcjL87VMvmKAF
73y9PYvS2Rx/HxzRYgcHrFy6KOO5cRwIOqBdzY3DZ8IfhEQOa3xa2lUSH+2YXPb0
rb1IhYcPclV4YYV6v+MG5m2xFB/VSaBeD0cWmzGQK0J8ej4kHW/1MPv/ZlkAJs5U
bc9hUKTlru7HSZTZhOL3o90h84fkCwrn9+3Oa3f8uyY5zDDIglumka3bAnmh/465
4Mk3PyATrIEY/8Rn5IUXFcethtQbvWR7U8YyImi5tF1YDbommRUQjp+/iWX8X/Nt
CpbU160dsKREb/KCmxTsi2D9F8LvybwH/8ICs8smSwS8hRU4tI0+a54gD0hc6Go9
2xt8Yfbh3enSB5NN/p4eLbLVX0bmIHscDm2SqjVBa69+/M5EQZzKxGd0jLyVAlKh
s4YeLiUrVoknXpmqZ9yemvhsgRnXvnruvGLYCjpnSQ1Lh+9xesKrDYWEuEPUsnxb
bZYUv9Er6mXhmvGxNuOoKJyVIyX/HfMVlFbVXn3Ty0Ug35R6QUqjpu1P2DM93W/t
AcHXMknHy+U9JIFxExz3KKpqt1ZlT/UitNmOJ1hOTyVqtiiyW4vy4Pommqc/yYo6
0B7pIR0+ZE2p5nPF3qVfVvgj+ZbWxnsIcOcTwARnkRgyhDmaOgoXUhb4jZUc1kZH
6Cz1JUX5U/vcB9CQROvEH6jBy8gJowuFXo04Y8XAf5qzZE3Slwt9vVd9uJEgl6un
iKElZBHgvGAvYxlrok2T54MjG113eEApi7N2weq+uutSSrgU8yVbKdBbxwuku3/0
eLPFt/gYUIf6ZCTKu/ZeI62OfQhmMRFAnXOEZlA41AgFzgTm7DNAeg2Hf+8o8VK6
fPvnnPyLdh2fJ026ShH8llAbrPjDQwdgDA49LxjbjddoF0RKOZjRgZDDYMDEPoZH
ILjMB1lS/MiKAUP0ctRq1WPMj2Hclq2pBRyEWpwFkCzey4lqikiBE8lTI/QjhuB+
LVe3/Duw9SU8CBxamen3Cyk86dcS8EiTy055MBHPaAMB+MJ8yV4pp5rsFFH5j5dx
Ek1sRNIjibWgbHw++IcOOeTVPrVakD5VcVDBKo0Hked9RlavF8fKRrGwZgZTvP0Z
s9CZNTG02OdHcwSqQeN5dGQ0mG0gaHHnI+4JEavgGaFQGOR+HfOSbKg3c5SfmXcv
t6FTFRgDaT2Gc+egzNy83jrqCg3oJxUl4j+8HoSy8ClW/jMJkoLgEddXYjVLYysJ
5Ds2HXuj1PELUpnBQBvTLO05wRr4KfbMwExUNhFXX9FqzhHkCacoITq0l/K9ewwW
0shhv+0H690fIkrhC3+YGRIqrDJ8vf6DRSz2fV4JWo2d7VzfVb74+fS0dxwIO4tm
VdoeiprMbzcXZMWaSxtBe0UsXT8nIWeywl62d7N22G9Nt/WKAy2LEiu8B7ZqbI9z
u56Zq+95wYJBIJc4v4izJKObbS/2J1sqFln5yoBXnlVm/rcX6vjo+7r2CpS3iC6t
h71joEDULvw+OtpzoJWjWTNqkX85l1W+cwwNlI+zXPr8RoW18emosfa4Xv4c30bQ
DvswjOSZNOFWpUCqLATnnb60zyx7jFZ8wWpuNR45rOVOKjRFJr4GcXBuWKLFl0wE
kfy8cZ9GsLNd++NIG9BdII0k0vbBxfhjayKLVMY0kGMxd4kOcpTwDlnBCTG+Qjeb
1hdvCgYPRQW6zoxjm2JLoiaK54pTZ32UP5oD3WpzdPp6uRyu/KxKdo6pZ51cx0mi
Fl8t+Re5o4p1DFH4kELnQ5XHC0BZqgkB+GR5M7/7KamLT+kCARMfHBZaaSazHfOo
Q1FnztPVPyYy2o76ACsSHDRt/8ZlqrCt9lAFie62Cl6jjN89IgkC4Nmn+V33X2mn
JCngig6WtgWiTAGtmxDIDBCWSuh4kIIeiqAeQu5LBUe5g8oIXJRSG2apb87ircdD
nJMQyFndyMWkvlh4W1g6FWSSYCveUt70AFSG+0hegDjbYUFm9ZlFNUcnBivcsEwH
BwGNaor+k/MIcIvM2QRe0DJl8amUXz1MGQfBa70Z2xo7YQK79rAcFfRTkDjkZM+J
HyuAVvK86XQgeAOBy3y74tKxfR8vWdB9tc/oxMVhAdvxYALJznm44BFDm6cGEcba
AblkzQBn2rodKa4YMvy/iZs0ha1M9CFxElauBanXTypCrezPNOcTvAhM4Tv8kSCG
TMDy929kBNqtXqjt+PxpVNs5eygb3+IEeO3zTTqjB0M0H7NzK8O5ai/Ns+LQVhCK
+lbFLxfDfhLucyQ6bmlc7SYvyVR0xeiESuhGnh7Di9x2IEr0x7fKpfbhsaXF3rNQ
AfktkNF1la+/SkreZaJgZRk4JUH2BFrm2zXdoDt9WUirnv52+cT+bkcQI1gF6BiU
3s7yu2QSI+zuvjGCHF+nmHjCqHsC4vaQW8IEjtNJrCzTFPmDvVgulpovVpYeDreY
0TySZqv/d2Fr3KahhDReDk+6f05+V/y01DIJsdALJZwJk05OybL+ASy6uUmxYKwG
RhcSgaqSf+G7IIeknFvScC4F4i8/AJdCoCvQJLf87sjs3nOMVtm5zFUzERgJRvCl
43GNAjH2lZrZulPEfLj58dFaAWTITmBriIwczIKmNbPJkRI0KzlVdhumpH75+CUY
LCxMNIqN1LQrPVWLz9voqxf/6rDl04zUbgWxc59U/d8ewuyXK2rvnl9Ov9Xnbne4
yuVDsz2hgLndLZJY4K5kp4yqf4mSzszc/3oP/njyeoI5uA1bVuF3JiM+tOf1iOs1
qqPVCVHO79PIA+J9cf8g8sFsUbT1yzwhSyWUCdSFn86Q4XwZFbNVJqonVixYkj9T
xlzy2qHgbXwC1EdNw6gqXvCUVAYUOlpXSt3gHDshwyba/Ozn/OEWD3IYYeIGqdhR
+LSSIf0oJ0MthSdIwXfff5L3f1OHpvAfKM354tlIWtdSD6H7mZgo5biUorC2maXV
TKaEfq2e5hmpHBO/K/HPQF7wowKE2qi6Ay4TEHMh2+f9B8xoxibv93H4Jp64s5Cf
f06C8usw5Y6W9/x1OHa10S9ZkFhUCXz9oFmZ1Oog/bTVcjErwvKfmfyXuQwz2RH2
gM/4wfsVCu4lZEoPddpjlquXrpr9zZ+6/j/y+yytlWcglrTQF9xTgK1yIialXc2d
RsJMlixk0dIoGQTQV/WP8d9hkeMVZCgYDHONKIjtljhRjzj5ogNCXnOg/2Xi9ox/
KjubDevuABktar0Qjqq+2OlZReoHrvERwDA8v+HlwWkvp9Fs4hY4MQSBaOksBi67
jqWCA97ocVvOf4qa1/ChYMbGdarNT+2DwbsXIUzcF7uv57EEktpjg5oeNVK5W777
RZIGpFj1Jvh5Di9YfjJ82QwBRlU8lcmWclazLajwj+QL9P2I08Q9qjNl2NDggNb1
uYIdZKvKnzp++Y0r1zAwhYTrJ12ewc6dLZgwArJkcPX2lcgJyi7r3Ple1DzNl0ST
dbgK8mK37675wqqKm4JqlxC8gdCBItVXGbjnFoBu3+nQgVR8mQgeYNBQ4khHR0cw
4c0a5KqDF8IrIp4AYO3hK/psRdTh+Llq+2d8c3WtDu3yPM5z8PIQonBuuzFXGp+Q
JdqNbH5KGYSm4Eryx3Q+bGxhCAwR56ZxJ/Ci3/7Gd6mZaG6GocckfATKjUePf1io
V9MXMWP1aKqb7T8SyNscxFw+ZKh9P08fVJUlS9dupxciZPQpBOIWhrwTG3RYTiN9
QFLmGIZzxBKH07sqoRBgkhAHLk3/NHzhJwdV8gKysFMXiECpV56Xf7yIJ52J44ke
SyVjAkSMEIAQoDZJdrcExZIHwI2RJDaUWSD5rsIY0c3h9xfxulNSIhiLPdOioICy
AXMngd1SjnpTxY7Pe3Pgu2xSDcIw/4HObaOjkWHLZBEZ1jaNDcRuS2tWqx7SHRQ6
2Qd3W8adyktUo2VKIgOvmh04OrLFge/IAHHjrJ41+LNHTzASqVAUGZJn8vKPL7ot
8xxVn2wcp/flZLUatiza45+paN+0Te0SgBwFLiU/+70xSko2To7E+OPCPLTA/JJL
9HQuTqcQqxvQjDrnGcTID+2l7pv9U5mZiYRlsVdJFxvBDvd+8wChWBl/dj+j5wN2
+kBm7AScher0pPjVjLVZUPILZT6NbxtAo3WZDzr3cN0BZlb40YwlRPO4dv63E/Xl
rivEe8fySD7vaot1DD4jxcCzAMPMyDU2PazEJeIUd2IW37gJb1MV7SCavl+irCYO
KrG8bOW0FUS884vtZUlkPoePCTn/+a3r9y4waCzG5I0TUMCyg9BZ2LX0kQzERPnA
e1E7N81xthxxotWKPU/zqz650sC2Va2AetVLV0IxM1XwpriIAK6dqUel1lA9wBgH
L8l1Qlb0QtyAfNEiKJyBWRmdrKJ5LWor1F7Y7XknTBXqRYJjQLqtyjXT/JnB+13P
EX3udQq2w/7wxgckqxgGCRqJZ9e2ebTGKDLP1FVjyC4n/mKIZ/gdhqmMqROMCZ8E
pSKd/MTf6XtO2QHFSgOPRW+zidQmk3E5Ybxyrywsk8QEoc5RhSPLd1gkkz7j3bH/
uwNQclupvCMH0zVZ5h5PWnXcz3R2BqucI80lqt5arjbl8l6rEECFW7LP34IW0oIT
2JQhcRQkf0u1UxHaciCZcpwMpmA0k61YHeHL7m5isjBq6qxAc9xjlEnbOl6iBHX/
AZTBxLW5f//yuoawOEj8pEgtt3wNwH3zrZ4E65u9p5AJjgRQuVyG8whrgoI6veMK
YzkgUzTAE92wS8TegqPRAVpHUaHaaMKBsC6LCOOM4o5OA2QYBTa6Uynh/hONjHfy
RCAeBh+dH6o4P6WE3YIWUXvcXX/5igaSL4RhOokV7NaN/dRI8vg1YlVucumRLPA/
Ra83eN1coUOTO6Or3BlfbiXaT4iuucbp/Rn0Ft7DnwFztxzfhX19B9Cm0VAOzCxn
xHNeoM9p2K23HV4A16+Di5vJFHqfa0Lq/QNtNLsjHGbLMfDXEI0FfqFrqpTMQf4z
9gYqA3IqTNWWuLjPfZa8Ux/yZ7Clakp3+Qus5n2dtj4zR8PYnKMBVYqmDuz2fxBv
q7gSwyZS98qRf/bF8FsQe2QewU7nWJXayYJQSS0/hURvj/UlWfYRb07MZdtPo0VZ
+dAN24kJG7dV4gIRj2dGd4bJE2BSVTPa5HrhN0eBGJQxGMLAfpjDVH0kz1LjeZi9
SlPLBsY9tV+euORJSqOh+vdxbm5o8VjtTqlW7rn40YKkDPvTqpdKNmIWuZBQmRpA
30zz2db2VVCpVWqhrndzYNfZwUkZNT0r+RacL/MfcVeXtholUwqAB6qFhoTCgcuK
xmb2n3lyGW07kqCdkalqwnmiI4gCuEFciqOgTbV9Xq0BXpiyEiW6X3+JE4EpmSD1
V5GG52FB1aXto0zNN47omhutTMgnMFG3JDhpll9O90TgnUFOvYpObfD9xKlCYQbl
436ksNHUKpw8NBqJ6urtolSngSfK+3uTi/Bb4/eDPv83zRMlOQsr3BOERcrx8nrs
05zTbAY90R63H/6RlXpBfpvkQCVQy9bc72DKFWA9PXXZ68VQn9KFZySwU7B+HDad
NWGHbKlsniBjelA0vvUWG41T+mySzBe/lQ4/1OjtH61PXbdEFjbCYpcVRyWNTGnY
vv93tqlgWma9m9T8GqIx42BgywkBFoySeP0HbqRM9S2iLHWwCkSpegSvmwDzWRKc
zk4JJZKINA6Y8gXFOwqO/JXesYhJpMyXrxrWgU279AGzVsuzi6Hgf9nkInAd9ysx
2FDLaU5MouJtfhhMq7vpsPbqOCjFA6POquxzC++sjYsMXs8B8cgR/B2xuyeUiYyl
YQPhGBPsa4K+0T85rdxrrtZWxVQZJVQq8mj7fIXx4EVXpsFh/hMtd6Lgw4GppKTV
3QZBBm9WSaG55iAG4rhfFHarguFZ2DLyPTd6fW/IdCCHP6KUfJ9MrI6wTKOio7dF
rEisF98Gwqq2CsKVCn4PMcCkMQ2WiBkN7o4aQ4Q9mc/SkH0P2UMRqhF5nK4k3nKx
G6Acle+zW26OLQRA0bUoU15BhdWecW6RX28FWoS35kQqX4q+WCFDeR7NJkdHZDuJ
7CKHc4ULGG2rQzY/5UExsVWDxgmTjsY4c1GBBO0V8GvsMQE5CZbZ1EGcHCRiq2n4
8At298ix2FeQPTQbtV2tHbBUyHda7RdoYKPfaHoEAry3GauDYH66NgkiCkc4QgXc
L0Jma4kHkBQC0+jNgVqYWMYoMM2jwU+beF6NhdkKWNx8320hkY7RTjncKv/yJsMB
Q7Xct7dgaua03CryCNLX7Fz64y7SUCeIXpOzVPPXRP4BciFsHF0mTQaeu2X8xLGa
fUF+NuM/YJh/4TOwB94e8XSdQgKqihLb9FFKacGNLPuiq1X3Mdn4k2/CN6YyhGMy
JRWH6MNxBCVTN59Phsxp5fqTcGDwFe+60roihbTImMNvg1idYtjxozsQ1TWfaIE1
aOvUTXwvTyqGxTQgY6XCb5e1lo+IKVGcqWwX+ehkWt6R5/Pir1N902yD4E7EVscP
DIcv9tbVK8ioTpCjZgOML1cBg0TYLj80NWRmmcFmYykbmTpVwmUjALB2KpF7y2pV
Vhm0uKM8sjq6goBSnykerr5S6rm6+Yi39lUQmiJW8ki9nCXfz+I4mhCSuhmW19Rn
EpIwDUJPdntWzPQTJTFIfwnBTDQLC2lQqxh6pV2AJg0NvWCoV8o6rDnaNX+Cpmsn
nWyAGDHUufe2uvEzCnmXMkULoOnfqh91uYPZpyFHs29/gW5/BxD8JA4A/zGavuAQ
LDZTDKDJJGri6GESeZQGWZ99a/AphRMYhqgkiPVMuMilWlJxd7RQGr1SDUB5RX5w
2ldq8gjRlGizFMV6aGv+NDEJeAj9dhcYXNKY+iEJiJQQAJNd66d6BJjNEDO3XWEF
eNmm8VTVLc6YEIzNgexfsiP2ukw44PkJaqy61Ol1/DEh50+dM/qZ4EGjmoYWlhh+
xjLMqVGh1C7y0/YH+weALMI61/O0VB/wLwlbQe93BgXAj9XA0nojqROEObf7Cn8U
jnlJ7VBGUjh6lFgpeIZup/V1l5eo5lwGvRqcztJmZ8zZdo48zd6A77Dcza+gLqYj
MWq2q2HwPNPeoVEdUUP1TpFj8/eS5UEqUuu2bkg/2/+1vcgKj1PZMHQUQ9CQGM1/
ShlFReNacnU7jDphBonbo9TyiZJdNSUAeQY0T3Vzzsusi0jSoEirxL4laMFZg5lz
7R98qlvERVu36+cw3t3rEiQToFwz+FssvBWoc5NJ7IqjNtwF6WrQ4+JgVNZb9uYk
qs++Yc8Zz4cVSoHeFCiLdaIIxhA0wWe7o6jzExSoqacbD+THitfbYqFSPH4115sS
iSiHGAGh7Rm994BAvJ58Qk+v0fU7hGgLr/ZWbtYWW7avQghVzpPPY2KG8Ksm4F/t
e2XwGxXYWLT3HKQlSmRyz37abxeq1xJQuqHxBz3JDgwFEdH0jqOn3nyuyl+F7lLo
J1wirqEgMW+zjmVM9lAmA9QSEPoFn5bB0Zt8i3kTxKtK22yJ6fbj+Y+r20hEsxLN
DdLuNp7w0OuNC4usMdG/sn8mPGZsAms4U8huJ4WmPwOzhzcJw6V6hM3JI3tEDN5U
5DVK0QP+3hV2krgW2hY9h2ATFc5p69WMruiFue5jNMeFHLWgPLgwAChQtHOkYg7S
LgXDvRNRpcpLZ65BdpLS+Rl+zFq04+OgDj6XJdmm4V9RPxBYgEbM3+59epcJlsFm
iL0XMAgWTRdybBBqxvm6xC+OpYa6kr1/ac5nTkdzhyEm6ojEBHPC5LcisHxEXZlN
27XXiYQx0DLOD0g+//L2OQnkAhOi0PUHam7Y3ezLH4QYuslU5YRsEpclzwfckaTG
NvhDTWToZi1VWut9HbNsPxVikOh35Bh7WHZgeaxJyCIS9SLZ1t39qRUl/JPL9nhx
tlPbWxhO62ysTWLekYQ/nHMpqk5FmDwsbd6e6h6OXPXjCt6UPYBizrzobOR80SFq
xrpHHO5O5WfxZt23JG4fvvHzxz3xclgxvzN0F+Bf3JYDc0tIb5auXTH3Qe+RME6K
OG9Hhs1QRTzyS5tFT+bR8EjwCQubKCoHnA4C/yOq8jzc03Wr95LzDzppxjKO8PdZ
49Tp5xGoM85Roku/Kby2wixF3EIInm82uF75RYYpdteQDcmJnaDRxb0wth6HtXAh
uzDAj54MHSh91sFrVVxo4aOOfN2wBXkHREbqjD96zA//atT2wcu1rWuHn1HXXaZ3
pKhI9iXi2PgYDvM2/ZA76Ybj6gAmUxSNtzhWTaLH/zXvVcjLdPYMrZeM7mdd8dLS
JV8yPYM58Oexy6qKGgQ01MfJwcsXt1LIA5RswcAMsPzL/fUF8XaF8+sHws5j2S42
sALcPSrn/ZO1VdNrsYPdAsIv2Xzhc9SL/I7CjWMHRPEDWe8qDHRjQQnMa6Lab+Yc
CjKzmPA3fJvqa2b6yMn4vrp8VU66/9Lxe2ws+Il9fAMSaOhgjOGa722WC1HZ57Uk
cv2F/VoL7tPXb/nk61HaUbCgmqQcd+tWwzm7Y18kpzLDzsD7ZAx6Xfyc5EbHNgi8
ZtmraeMdRwXkZi2jEk3vVx1OKwqTW7yEqxSrJxGI/nieE7jUE7bbRKp83rCY7yuo
HL1E1aSEerKfSsdJzqKYTr9+8iS1C25OOrkuC6eYNVTFFKWZ3JL7GviWYs5pL+u3
OAIgLDwa+0/EHoAJonK/zTU0FFHNWM1TgifSb9rQw6Q1ImRbMpqUh168Mbrk8BXV
OrKI48ZSY/wjGPwwrkXXAag1KGdgALloAEWoiuWvmxmhIsmJ7UyBZRpNgBbH2HSo
jt65naYJnwJ73DX614Sx69aoJcQpXuVZ3B3ZBe6v9mHH4Z7kHZxJr1rXus2/Y9l0
jT95ucU9gMxkTmvzn0O5yUqdK2GRuuPDfBTMdQxrDu/FdS4vCMFfJYytspU3VNcA
J7rW1eLFilbRMzY7Xdq9iwGJt9GcUKZwi7Yi3EAZQGLLZ7UiCHt6xJElz++Ib42c
XUHIlrtwvANaO+R0+nM68rS+0rCo+RAgF8CeTmgTkR6HhNWnmZQVVSARAKuu85jO
XJdza/fNPdlUVQ1qLObR5L6Sdyq8unYthHJWwogvU7G5g4egxIa5N5o9kjSODxyP
5jr6E8LJ6c7ANm51kBw3P2DTRPao//GjZOpGsJsTh/dcHkzh7Id6YTNeVyFk1t7X
i4fZW9WJuU8xCOSbDtL3/GYn9byyCTSTy/OPJdO7VRYx0rK7dZumhyruq9JLKScK
0Dbr5tjZXdJ9VCd0+agDOqqaMkUfJdmmGBE3x+4zrvJ6mRFYpJUpGySWQuEaZAvO
IkCKJIdBnSlZfQnJafLM6We8DxWzDn9BacaMi5cZVIXWlZRqA2K+pWPeIXO40tFd
HwIxmvtjyZ3ZiPmPYJvBEiLFcLIge2BFlzA0Te77NZ1dda2+1YehHhwomSIFWIWK
eAnH2j2U13vvzKI/xIwMxijb1fhEY5r19jQw0YL3XC5KeE3V6idvlCZkWKh+C01o
q/sl96sDCOmRRObZnHMyb9e0lsLDtuw6+pQ+h3FBa7EEGKdKdU0m9AKrZKNdL8kG
kGMR0aEhUY+wSzivAbj5ia9arKrBdb4hSwJ4GondRWAHN/XPsOJ4d7ohi8ByviT0
Nb06MPVwagtq40ofOTmFmCLmoeD4dhloOjkwvcnPEc81kYVoTeMnnk3/3q+FXPZU
vChEy2XPUqDImVSZGaGMTAhV8jq4k5KFEDDXgkO/O3VL8mXjud42at3J/u/uUKzX
UlVTZ9AyK9nblziqA13FsoCQ8LThfcljtU2iLNK7QSRwVtuPE5u5KG0IWf2BGr/y
laS5C+G5sQS2d0tTX99GddacwSlShBk1gIP2J3JVGatT74/HFzj0i3Uwt9ulpWjL
cen084nJ3SgPXumDJ/e+3Bdyz1pFGtlmjWAEfL9RcQTX3tRiYAuX4RDMV2wZqQ53
mUraSu2Oj53ukklRZEKp42mm8zqLhkDk4k6kmaAJiyqB6xXzX1mpQQOCVW59Q/rR
EKHuJ9iCrirrN4voAm6jX6djgqhezc3OM3qzifpAyNgk9ZXPA/dyxR149yxPfrY1
G4UEAPZJM2aRlf+G1RY6NPeoRtnvO2r7lwhPlBstGqZrF4oFKUHB6dR+DKGR/cOz
+pkqgI6ZphUDDdyTFcOEBq1xdQfmLDjqHtjuR/u/mOeBc9Qd5OG+qVyPFXcY+uld
m8jBXx8qdQWnl1KZh091g97NG0X+eloLvumm8gG+G4jQyIJkpkd5DDuJW0RKjvd+
MbcTiR/WaZfMmnuehNcywg4M6bfHgfFvsL/Ls8Et3NtwFYSGzR1gwgoEjC7B70/j
hiRoTmz5IOirBfsEzfRYc3e2VJ5HCpyxYWAtC3KBVY5NO+PgZA63St6QSP3SSI98
hGHmrxsKZ1v5YLxlw5Sr7sn3Bqya2Ridigx8YbMXpXsZgBBNWSArKoKlVt5gMLDg
v2NpSCAPaNs+nqGloD7fxU3xithYTcxUWbDnIUj7B8KmqcxL4D5tW/MfOgVs+ohk
qVqr4fCdDPczR5MEagWHh6z3zHC6GZ2aZf/VtPRrAue6uMK5Pd6JYgmRdPea79vW
6B+weoVpekZUdTSRmtIqyX9lWvAfMcPuqyVYLFEyp+gJg3z2oYhS66mAgOkY6ESe
PMWWsLGrT+M00FIWpOvok3RwlbLfV2iLhJXJ6n7b6DXixd8Pjc+Q4fmwMJ7zf1gT
PDnZ8C3qmi1pwdbk2J2tjVVttTi+TZ/Ihmk0z0rpMOT9OSKUg47DXzdnIlXBvX+1
1G6Qv6z1i7WaKhKJni6tnAq/bG7Z3SqUCiBEii8jDRD7AFQ9jHJZPxqXRXlEq+6K
nGokMZhHpDVN0at1saPRmWxU635EO6NGkG8dR5yKi12wY+FVVrriLevZGPwQf7Jr
sd63/XndPX2h4E3MGvsPTpYodpc/yJ/iruHd6oQI2j88O3AWILSRNhlSeFfrM4XS
5M1vIMEFTr4JYDIzhrHwBGlscXx4pLiGAzzlQT6rCynv0fBpy/s8rP3GB1E3TLlS
PlCSkPz0kU750vpd/A47r+H/9uuiGzbsXVMuDSXjGk+gHTWuBsrgVC4CeBb513vg
JwlnFJmzx0LCJz8o38YvcYBUsBCQJBtoqR7dKqDnmD2hT7uzUhYP0GyhrXF/aID/
Co1lNp1APJozOhGBYMYSsD6HP4BsQF1Xl4fQH6eYgvm0eyBrarcB5Jr6Dxoev2BH
JsnjiH7fVj4VAyB7wM3eRk96k6VVny8/d4hvXNv2VXf2FgGlgrX0SuqrZLLGN4XB
SFqxgthbwZyxysknoioH+4h/6sru7aNnRnpEmZ287wSI/tHzxN9kS33V/MLaLXKD
EgtUymUdF/LoQjTLqgEGfeTOtR64Oq3va7o5Vi2W63NN2gUmXFl9Xn6zrRb0S+T0
2RVn1la1eooZ/77UTL42On8IpEf8xA2+B8Bu42wX7fM7oNDfe+cLvh52c0o5Js4c
bAi0dOhrK5FEtk1l8l4LOmNA6c1IZijreSQstGtw+Ht9JB8ZBGC9VVZSUDo28yXA
1hYiC+J1VSA0X21iFUIGmjIB530LH3KiuoWWNv90XcEwNBABF27P1X0DWE16xtM8
gGNXqSb/wOA1GnQ+bBQ3cJhCburZa7zAJTNhIH++c37YiMnOqFOa1DxEP3cVg4TJ
hVe2S/y+72xaL/UnRh9k6E0OI4LgZ/ZErhrtrEoI+DwwEp/MRXF1Y3rw+I60o01k
fp1sbvtKqXHt2ASZBViwyvtpul9YgdT56e8m+6Sx7y5Zj2FeoA4AhGQDvtpc6NMD
aaDkRR19p9VD7DZ1V1OV6AOR/GkOsQsX28NS4MemsGOX+h4OpmG8zDqmAjPQrYIl
rT+huolcnzvs09/XMLLD6kmsJWfGT0ZJ2d6y/77AGFnkjxdkEH5vkpIQ3nTLOHIe
7MwQWTKRF+ql0V+aYSyscoXAkckW1dWPOYwTPLJDhvFtBMB5Bg0cKo2KV6xeY79g
8lMcSPVpRijDWuZlNhY/I+qBVEYG/TnYkBJdlT2ghwgK/M3YeXrIvNqlmwFd81Gi
zaCxSBoMLAqPhaj0FxGuV1faSj7cfsMzgm2YL/IUOHAE4jjeHVH/0A5PJ2tbTyps
fJZBLi0nCtnFEwQpZK2R5tkJ8PLQ4mWnlYjvnbnVneu7GwVbzekmWsBD1418uZZx
+wVQStYVyGGwbFWTgc/sQBenOdDUDp+x1Gl/p7xwkNVEUU5hZ9XqWVt3cwIPQAhR
qyVY5SHDgI1tZMZViRrk2STKGhESiw93X1XHVIDsiopfK642drgp0eCvuZCNZ9Bq
ttdU89laDAkOe4J6tm6JxMC0/3gAal4z0D/bh+uQV2B+JWKm2YDKSw/65cIeCu8+
H4oQJJ8S98UsHA0wdaVhhAUOakki1cVfDlw2Pf81CzruoGGUkBGv/enqqBX9qANW
i/KcOy0mG/DXUDYXGN7kU964OMErQGTq36xDlIGZAtXtf1/D5w/wTWukv/Yb2kFy
ngitybHp+fesT7Ogb1SmDmkR8T21C/T96zWZSrsuQP0dna5qkMbvppCUGrfIGD7W
XCyO+XxWmDAci3kGCRlVnOh4cU8Xudk+P2aK2we/bkz+fBNlHXpDx0saPodybtef
X5xzqvKW30G1JwXwaUZqw/H64HSRWeMC0xVvhn4wjvCzM38Nf1iUfRr7A7d48VmB
i6B5LNsKYJAPgiIArD3ixevEA+Tet5j7dVaN+4Kaw4NLelYIqRnIcvMzdN9jzSDu
WN3B3VPrtwoZvAodatwDo1EfcYq8hasTR/xaGkkSdQIVzWnhZAkn8XVenO+xE9Uf
Zc4836VG8VRx5NcNLE3dd/1zuz+rP0n0CRllmAwaYvedJf7Q5E0LGUHtZ3QkndY4
GmTkmFg6deT4C2kR9zFHUYJlbjzZKypip6NzZCIBJamHfaDUIRKjj1eRehE1MeCq
cvMiML3VG6Ibfk90wsNT8+M8JtYABMMK5FTbrls4SwTjlt9Vm2gTBuMfsw43Zk4k
uvHvi9wClTT4MqUlEfQBvXqxHxd14K9NzoniE/IjQtxtiC19/WpfF70sf2fadirW
cvcP4NigiKqnEw4/n/gCgFO8yJVxJJzlOGxuYxkiUVmM+BOkUe5d+26iWWQm07Dt
FBh8NJFwxpRUcW4D0/fcDK2ipOm0hISohfDPILLqjhDCp35GmzyCPjwKCR0B0SZm
mYvu/rjZ3bJx3F7bWR5hTMGmuYtWSpz6LEE2epYS3GCNWtH3TpoUE18s9tq6P7N+
VhqwvdFE9jSJH7cnJi8iIv/QN1HAZzE1Kq89me+kuQRdVNJAi4qo4RPGkEpfMxb4
Z4bzB7F+RGwNNQhx+UaBm/em1e8TOZGCspUe1bEALUFOXc9QpHvnTZSlD7cMYqLk
HSjIejr95uXRSWMQmR3gppennAD4/Vc3rdh7HAjKxF6g65pELO118y28QkJ5Kdk6
LpWp0N5U4b6nHWU/Qod29lQojELjZ28vKKQDsFQNWwLHBvvF6HxwgCtRdLESzaZP
n3FQfQyTWRekMiS933+THBuZ+B6XxhdCcqJsawLeiB+40YzaPhOHgPz1veKmxYqa
QruE9JXTAyI3tSIph3rKOUWuUIATC4/7kBAq+6I+T1VzzDM6YC9tsTORtcrwD6mZ
l/YlIfsCCl1r9vor5eWGNQttqZKMz42EYjmA0jjcbIpch8IPYyfPmQJ1IjEgXWdW
RL6vhJV5t30a8q6b19LYAWvdsnpF6AidTBGB46YDrJRu5Cc9iD/LaYArXUdkmytU
gzDSO/XiD5S/8Pgba8h2kBa+qE76UwD7JCMntAck0tu4JN3VaJogM5/xgOsRUZux
TgSQcrwzf15HVnz3xPYijpGJxQHLNfj81hXILh2bhjEaRZolsEiMmGXagWsiXy1l
mLjoU1yyqxhGqSyDeDA6nkmr3RerKNqIQyMpqoHgLWnu6fvHpFqrjRzpRPoHpO0b
2eol6gXZ9mSz49MwToB3PzzNK2M78nvcl+yXJ3zbfvmnfLOFNZxphNLbcmvfqXct
Lnuv7GPl8J36qgGXW/0xKKYKA8ZBFCULwHtwUG9yV/oQI0kz+1EbNpOTL33F0o0k
g12GP9vFx17Tw3QU3Vm13npndzFFq/I0/CRXP87PzuU2x2hjmTDVDrL4NRqh1XcA
NK3CpPSTQXmBc9I8Xbi1TKUSX7l7pQIr7HNt84XvOjaWyuzY/vT/1HEw6OoZ4za2
jRrw/oirRuy1obqiE0cOkc05+MxV0DFVzqrKDSsRWbFZmJyUhSB2Tx0FhYSdOOxi
XohUsBURVR4kX+cQ9gNzoDDYHLZoxgyK6eB86XWsZoghzvbe8eMo80szvympJcFd
gjpHrZx/uPsGhZK3oPi9eM8Pqmd0Pq6eHQGsJM6DrtRSM7MH3jpP5SSocV94BQxo
QDuhYgLHHyMD2JlfvbGVrd0q1tEtrqOdHcD4cdCmwNjJ3knaEyAUJohizsegcLA8
sgWV6agPHcw1lm4o9ChZ/48XOa06yhUR2KnP1wcxZTe3rg8z9ySGj8PD+1fXVPoC
xnzCH8axUc8JDSkk2hB+X78ELtiqsd2YioEKxxDoJY4dlR8GhN/txRGCZeLUIDIG
ZyOaOH6H91v9Nu61nO831QoO7x9IMphTPMIo2yQm1fbxNB8sb6yCOWFLZMvi1Vdi
s1Ky0qGs7oFncoagh2R7YujaP6S9oR2iv2znwH65wjzakk1WQZX81GazvvOi9hjn
TQK9rxbmv7TnbdFp+ph9WQvyh9Dm+MrO40s8eyKHLqpkfp1YBlkZ9mSQq+Ig0KEf
KPvNJYVLpAovj+PeGQEp+cwkJIHChKEH3xx2xA2HGM264uu43Gb2T7Qmv2D/KsBG
sM1c+qlX6e99npd3mK5lk2xerCokWNHYcq2ABoYw/H7BNEsa91Z9fIROhx1vyW+L
1J8lY9ojq9UIcbhOh6M7kj1TYolO9v8w08yIY7nML5x/VTPkULHoVT+nIpa2omFf
QWvVY7h+SaWd2eUgq4zhaXatlToajqFTMMQhUJsigxUD0wQVccCERFFK9VaNdJ3p
ztn7lBEWuzjrRGPQFjtylgYgQEUdyrGFUAB2SmtXox0efsA3q1oriw8OA4MeL64t
HF0dxTcuNQdwsHxepE8htrVhg9hANAotnttGzMMhb9RA+0vFzSp2TLANXlAEiqCr
HHkwDJVcpIE0vk14Y4TkPjI/BR4iRgKBtCnempeEalo5hLt0H83UacULqsGVuV80
nyO/MDvXo+8oltN7m3/EKflUIBtzgi83hZUC5n3fkxtn4uQDe/JKNNH+FMBql1xb
tRNQZW+8w0/srnLDegR1QFTugxcb1p/v1EUgCi7tOMalKm6UR+SsrHprRqFRSsCT
woGzD35Klk/QyidVecdswi3f1M9b4KpmjeikdQhbIP68XC9ToprG62RYGEaWufVS
7lJ9CtgokdtiehqoF4yEnzCKP2JH2VYe5ky9N6i3Vz2ADLUNbofdoZlZlb3SCtp2
mIe/Jp9czhiV2cKbpCC/A9Rbq6LzMNlQcrF/I+27B4ZMl01SrLAiTdmbsWhiUuq+
Bn3TsE0PgzDHMEqavqo2k2al66Nn/yFJIHRZd5eoyMrDsTlIhLI9BJTmoCqduFGr
jVz/Pg2CicW8WN9iLjxwX8/ip6PapX46GWYPtyekSK3pODO/WYmQNVKlD4T0kALj
BZ4xDVUg0ClCwdUr19n1u0oL4866WUiHFoh634IiFIb6BE4Z2dS3gUsGpTu5M2Fk
dTS1seJBF+icZvqBMlQVimCBgIisw4oxBy1EvE4G6biLm4Ud6vZQA+UnHjnUdiqP
a5jewfvXWK4G4Rdkq4Mk2flMo0a8QNt5sJSiWl2fNIATxI/LlmQRvO1EPWAZUTGi
bv13+goMWN3gJZPCkpokaeff1Sjxp3aP89yKEkifNB1TxLZdKFPp8SSd6tjUFzpP
FxRr1J218WcwctUlXQ27UCXhWML1IBRHO1+ruMbTIQxg0o1TObKuwCGFWRJHQstl
sBh2el9913L76DrJEjfONlqVNtxx3+ZYnr+0jU0G/XM435P0pSNDTxQHkoe5zD2+
PseIf31Sl9A1fMQDk5uTlli6z7F250A1BGYLs+3ehvWLQLv7umdiiGpufNco6ByI
rZb/3p+4Z9oPidCl69mL5Xhn0v56/6JA7KV/KRHIfnfQVL9kLN+86ZXQsr+YwWfk
a1D2JXTYRvKqEUABMuk2x9EI52hda8mEtubIsJoBFMFOXWpnVQWRtSRuZXO4Bm/P
37i8yZU2RH54BoWe/VuCbnmD+O5odNLOwysmCiUtZaAz8KEVyBGNswOOM8A4hXR2
s1n5nQnXilMjhw3osNeYczhkmBY68dqlLvgZh9Dls57VFSCwcAWmaKQyo6LY0aTD
xdR61RgjuvjhHT/O7vPmzLyz7qX2CiDGjWuTTDHaRFKlIbRGsR1pPUW4zcgn8bG1
cDoD4cNa00i7BE+sVSdrGZiNExGipvzvrHE1N61S9Sq89XP7l5aCvJy+QrgYLNlb
v6mGCv7c/TzYu+qNMY07YS6vftQKp8XHt/T73Wt/nZHj58xrBQfF7k1jEwdaw9Rp
6uumsHEfxZtrgahvZJ3dfDpMVCXknCkMLdY9/R5AkP7s3n8sstw2LivDoVKW6Di9
O6DcZkuyM2QCbLYXYPnx0VqOvIqZ06vtIuEXXvvPYKNdeDvAClj7gGbuxsF2hW1o
UnzwNJ1SbL3y4ZZdzbjJBhQeOtT1Q+9dxjOxtpPnfc+PUg9weY5aN5T06ibHpoas
CsHqUYA55NH6jqsevZyBv0JD6EuygzjseUYcaAJ9FsXAwD4YD5lP8WNYsIldfvmX
g8SaIAj6xij73gLgl+0mNiWksDsGCymutXzvpnL8rrGa8+GDc6ricD8YjecA3RgA
Ga27iN0vbtEj8vQ3lMhXdTzinFV14ULE8CaGgZlinoWXQRC9TS7CUcNI4JRNuZpc
iRn3i6ew9CBQKTNhTf5JpIrRtj+aF6Qvvueb1USzPuJYOj+xhndLD9COU3hNrQAp
Ao36cFicH67T2qEYdEADXVgtM7VqxSU+/kg79FqS7ghLL62lc9HEi6UXqbuRHCq5
v2/3ya7i9s8JxqB/2rJ6qE/eukookdl0wfnuIByB6harmT1M38SPEc0ua/wgCk+F
tlyp6ILtNjrjZeY4UC+AtaPllMjea0VyRGQ6xGYaql4JixmigW2xkafaOSyuWAyi
JnSQPvzfSn0EAlTfVX/+HBJFW7SwsZUvacBvhHmO7rfTb8s712UVELu837SyHTj+
mZ69Oq92EJ1NQyTRVwnkvQqrT8/lTAy8X8BSV/63mEU5FRooGQ4wIEHKoYrjMtaa
tWqiiJyECdKdrDHI5gw1CzCEDMQ1qnJNIGRu8D6fBPUEr+K9h1zVaRxGXbJmyDFb
E2P+CLrBPyOT9znDm9ap27gIQUJ4BEr9mfNNt915KWJDspkb8xWI0/v0/IAyV8qc
n5LEJO6AqUYa6I/mgU5S2/Wtpsvj53Sh5VP3Ya5SYQas77GNpiAH5wYlZDeD7A0g
1SuzcQ4MRMS6QG0fbcAywiA1z2GJcSz6gIcETcHxLPvN/BmkyficTphC/lvNYQU4
30a62veCCnl/DB3E1trJsEsqnR6gz7E6orZZ6RCrNETF1KB+MIKVUR36U02iLE1g
Zd/RHEoNOq8ZkhjxNpB/jY6GU1+J2b33NGxmRTU+R36Js/LzbIiHk/fwVtWsxNgQ
v0D+PIA2Pd1iuiCHkaQhc5NUdN1k+KGcNHd62SuLLP5VA8nZU+J9+YkpiLs5xCxz
3CvyeVrIuHk2zoNniwjZUhbhuHlZXVP5raOYDh6Rx6UkSV0Mfk7/xJtK0gg/RBuh
TidK+mop5wUn0EOXlp53VGh4fRm01BzC7AQwOaKcVq5nauoWrY+nPk3DSXX7XdAY
qLYTj/8E6DpqWvkpVgTjRHKCw3Ni39g/MzHNkXf6BUJAnKSRHuQ82goMLTrr9bk1
pHml2OLaK5pNZIJl/vy4n/wjeSJVnEZaVJBkHU3ZnApxkCmKmUjujtHC48dT0fUe
x99g9BO94no8V+BCVCjgbnm/TIzycb7JcfwMe5kAfpF8pNw2R3UgReNgZ727F4gT
ueoDHtKiME1fq10axusmVpb4sgDDGNvqqXQhaw8FevZ12Q3+6udW431Ly/oIBEdy
IsVrAJD0SltAPRzwCXPThhQ15wLbP+0eUDrinqBROqGEiIYzJYL4BlxZpyRGjRNM
VuYCXS5nlsrMCaSPyJ84RIepiyw8fLduFlDgvuogwDAgIzS/I4kt2/U9/DkzfFc1
NzMTLQvf58aKew6evaCLwoicNCdA43Sdwrqy6IgN8yGhi8FUw1ztw3sJySeiHWTd
Kl35S0MiIMWRbzw/gBIY8DwHWts0YMiwkSTCgDLKI4mY9VjppikzT7zVfbk7ZzUu
Y9KblLxExXEV1FKLQuZm+L40LVYhCAOV6q8WNGZ85y+mjO9z0IGMMIK3j2r87KTR
nCNitUds+4TyCfoh27pIpMFfv8mIpkhn93+Ap5mJLMK6J2IoM1gEr0EpHdx/dHxn
8LT6D2o61aU1amTsCRbSmJJne6rd0Vf3ucczqM0RxgtxMOAMIixH9wGRQl72j2qU
JVJTEuWnFqugIV04dYdOHpiPgDzevKMzqsKoFKapbgFXr5I/gySvDWVIsy85C/B3
mkIgUMi6vbrEd75Jq1fkjmFsP5b8peeBu5UD6EictSX41D75CRZFA1JAwLVbu9OO
LgsBban8C6lReY7tLO8nMZrcL8nEzKjoBu01+ywPFs/t+qRfR4pLsCfwRuYsdvca
aZ85Nq8pOTbVwb57atwNSThUgz67iiOClCKZOJqo8xOgNpEA7xOyXY61DjTrbSTg
6/p5kGzR8ZAUvWhgYfIcvk05lW3rVM5nIC+56X/sJPiYa2Of5+Fo54PmCOzps5kL
DBNrVExGpf/mItJhaiva+XXbcyGzJNZXxmswuA6aZko883z3nGJAFxzqZYbsMz/o
d3tLFfwHItOzBco5NsZLZW1LkEYjhl8+EI3jfhjjDOdzVNbrMAr4jbjLD3BlEQEj
Qoxo26ZpgKdY8AKrF/QSY0waDbELl15roBN7dQT/zZW0Xpx0DELuEnRUbg4XhiAM
SpbSGnTOe78bsmuEGpIqZFWL7pUNrav39nmahHXgWWYTEONQnNXAxL4m0ujd+XI1
CsJEJtUSwBPXiseHJc9sR/NWGIWRAZImKBpHgeYMvtPBRZ+YY0Y779Km31os27JZ
PI+F+an8mocVx0SgEmqSEVjnGHr9EY+TXetaaC6JCN7uPOwZ1k0TZMKQKP5o+me1
PImdxzAiP6wzCgVX9K/XJPOeBPTCcxFLO3ORX6ptpAhXbqv865uzo5ByjavtdlQ8
0WQ54aS2ha4gP9FEtSV1p7lhvalYg6G4F6cNofYtQrPg2ZFfOpsz1L5XjzO3rY0G
qMbLeAz6XoCx+mNzV1bYiZOpI8BqtDOepxlq5fDstBOfaBoDOXVAAIve5lTPEntn
QQRq5uId5I3pMP4eddA7HHlL2oPVZLyXWfIOHIeQHzqNNIeiAIeJuq5+a9aQ3CIm
LL7zX4jU5n22uRoAaxklmhGC1zTGT6NSiLjuhy4SAPRfA4GUXbr9jDWQBFOncU4G
zhFRs6m6BsL6dXLeKkW4pY9Y+wIwPIWIkGzjqeSnTDLfQNzta4pkxLYrl+HQ6ebp
D/YRySheHGwiaTapR7PNhrUAVxgzbLlHHBUk0M+SEu8j7WibhujWWAJvDLNIv9Z/
UHVXIHs2bZ2qvQ1HK4tCYGDFQD3lMjqF9+60XPKdup7btW2FLAT8lQJk2SSPfDcr
llSWZCKJv7GAb5jUYyrbyg0z2F7wFKSoEE4Y7d7tnP1xGBcMDkDANQ2BLspsT9C8
K7q6iandO78kyJ1mL5zQMEDS4C1RoKG9QFDzd8YBVSkM7GVs7ZV+QgBoasqcvPIQ
CYfOzjXBhWSNPhOIS0S/srUCw5/idUf9E3r2BottoTG8NuJ783o+4dFqrNdBX3/U
ve1Y36pyeYEMxc30eRzfeAIZ9+D6O38CuBA0AcCW7WxPVZbo6dKBrhajuH/8Ca2k
VV6D74nlfhUetSfE0cujQdIhgt1Z88vFZZvzryGf0R8ZDDOZ97lt3Sp29j6SyOQs
b8k2sEeZY6Gmg+MukDOslrVZvSOVB01jwpJvQ68w1FJSLuVeJgr8a3HphwX67ZDW
lkpo6PAqCjIlM0r0bBosHVBcD2+rRgvLfkzuaRaeTCLqcoKT//B6VEMqbKnuanm5
KZE7pGzbu9NhQDfIReMboBs1VXwEzaSzinF2kFz17U1kMEzDEChjkIG2tMssKUkL
Ju5geXlMlhprgT0Uom7A7hdkiSHLmAgxQkNnH4/HlYb4VMw81pU/StI4RRprzRpW
TmFQh9i+ERe4uO60ksdc45BF4aztJmPIeXi76cWNmxToq8nNBijLgOiRc8ilN+G+
mYAo/+BWQruDJiWePN4AMNHSozR9DnqcFPDv6OofcemMXFVYlrXdVfJQGGV2n821
eILIDc4aXBSN6wF5M31UKHSZ8L/rNWGrGKYbDcBbEmoDjPVCsYOTjRiRHCkUTO+q
rXL6g5gtMzlztuSlj9AGN84GDXCrzkRuhkiJ0ZHSyOVGy15gpcgAFnybCFZCevRP
ZmdJid1liGtAkxMBwSIZMwZoErOK5M1U6t0eTnJW0lsQaXBWtc+obiLKWB+jJiXM
gqUumff0aGAdLOM38RD2wy59LdV3QPTcl2/1vEUqK4au4xzPu4uVLz/I0oibPknW
37Bkzn+CmyL+Z4W/g5aRsaF0mAnmVZHRzv9XMMVAUaG37n6kO6WFwAoIJg0UEsz3
Y0HJVr0GuXaw4Q2BUHTxeBqfh+0ve0U8EqYfNM6++rXzCMYdF/afVlLW3Dm02G/g
+ABc1aGi2bkuzYA7p75kdy0wFJ8xJkYUEZiuEqzZIBXbsXf27XNuaT8AK9DEEJ4t
vdOs2/ZnR5ytPhdKdj2XldMOv/xrIc6ADfO3ujIsdyqxP6khKsdre9zAWxCwHuEv
gQXCWmz+MivI5vgfXIVBm5YW0hBP/NuU15jz5dnsbFzDFormnASJexfu9WLoFk23
hqgPY1Y0hGHyd7c7ppkzTsNDsXiGRywcQM/XCbre7+zo0pSYtF+h2/V2ShAzATT1
PXv9+7f//ltC+hxz+llxeVNA+a/2/qO5nEDSibKMknqgZ70e3XevzaKrPJS+K9cc
S2YzJGXyarc2lX1ck4Q2oi8G33QGv1Rlp+IPhmDlRuBqRaKw9tEHWfje6tTFbGOf
Z0rPFM2lK14N7up4yuRk+6YsmiXUjmUnrazMnxJtdh2sp48sK6Hx+A0ydhbGzdCv
8y5Z0h+A59CzBDRMR9F4Dtcr6byjPKC8cuexcWKYR+0bkkqjJ6Foy624bVLlpbNI
5tETRKBJ77YNzGzdIGtsjlAX9Hk83kzxEpq8fODU9Lb0AQL9VELVWlZXsoFlQSfT
mJTtU0oSQSpVlTiXO2c7fBKoklonpGriI/BzNzkAx/6j7b8a2wdIQS2ZvmZ4I3GB
+z5i7tBk3M7g5DF4So1NDxemb7pr4zl61SfuOxdiMHVrDa2voY03FPIHmDHn/O4e
EYu3uY4d/4cPPVBLe5CzWdOzYWgOk2jZktKEoMOvowkCAs4PFVTBsZs9Ex60VQ1G
FB6Bb1H30UTRqJJ05Ka3jrcMrQMhS4rDHab8G/wbjYkjfGsFOb1TO89GQFjHckei
KMvaYdRWfpGyw7jtUQaFbbv6HqwKXpSY3x/BDIjAbg0H2HLIcGNgm/Est3IpGgg/
JVVCxy78A42NWXrv/2VKuWUTZMBEZZY9zVdruRkZ2p/kxhLJXszE3B5rm2KGfZhN
OTJeiJn6Ti0r3uBATP+v9QPQUaPqe7gXfAp3hxI6WdLJLAB3ZKvmvNIVc7+pocVK
J0zpmxbjPJfsmzS2PK7cyNUQvcOAag5KP6v9Z616Y4ng4BHBblFCXoCY0ps2ki0A
4jefJqWENKexSFiatnLGVJkZTug5bosnLu8n13BuBpP2xHYWGxoQX14zm07laKH0
EKMfO2IUFFRzIbRuh0Wqb1K+YryR/YaTfncvLm0QlT0ebza5Vtq75W9yJ9/tPlA8
Mmg+y03Jm6h39i0lMnflPZeFg+BaHzkytgyPJVaNotS+n74G/9+H7/BsugjBikrO
l/HEn2dOBfsyMWKu4It8qEh6YlE5W1T61FhD9zkiVcVuHYe8kkh+n1PvsBJPvpnM
lZ6ptDRyX6g4rV5+x9S1vD5B4onXUzDrvHwOn+IYX+hQsA6JQ3YG3yTc1abpXYxL
nMOjls0754lB8Fk2fIxxS5xebVSvVD4AOoFVJ5Xo9WePg76p52T/Ky/7+5LQsupO
6IT0TNE8cDJfib7cpl9PquKZcWq7ibOdq961i0Z0kb7Ez5hhBEPvdn4oWv72BzqL
tZYWdVIVgzNbrOY9ie5Xq3midWT1q6UtOI/+Co28Cc9J7zqHJSzjQg/WXJwfVHzM
GnsJF6n0myw4TEsIqI7eof6CNiaRuJt3dDQlTR6S8JMZflcfAryJTsaOURZzBioU
qthvwWCx02qoGQDLAZet39Mb2d3s4QzRtaH2P7/5MJ4YCJHYPMSD07jGJMYU8zas
c8Z6A7ojOEj8HyqzPxpFVWSRy/0DrIH8DtrYzrhlbHJDKIJwx9C0Xw9LrlfNwVL0
E1AsmHwV4sNqv+h6EA0xa+kKlF0x4kttBrIdvHUJhf/fJ6Qvp/Po5qsK3SPPxl26
28hu3u4H1TYtcYGwkHCWLfaAqVRkVTj9HttPRi5ykIShKS4XDi9/mNyBQ8T3ff6o
dbGEDYtjoYgBrupDz9dSI+fN2JLgt74AFPLAkYzLq4fjt+BuNO+NC1dYI77j0iUy
AnMtreKhfNb70Xqd7IasD9GZ3WTwO70zhfjSQ6/P/VHOizZrvD6loJFMsJi86OXd
PXrTYyGZNY1GiYKx8+lCtlKPu2RGVMULdADJ9i5h1tenaRx08s9Bp/+F0DBX3yvs
go2nvKh8cmbVSnp5Iri3BCqetZw8IjjnXXn5CsBNOVhLNvEBfM4WE7vuUdDqNN9I
t3z6yU8KwCXUbwBi9QDFFHtbvNBorTqOJCxf2PspoeKO/74BV3zpLst/8bRROICP
fgSN4tRnZhSs6Ib+5i8W7QUeXE5dq7KSrTSyPioyqSM0NihdQ/kzAmX5jj27Y02a
+L9j6TnNDBQERAw2tMAghr+GtAqugvaWcc2jjnKHCKvvNBR4xMbH3Qs30P3feIJm
YA3hZ+mndNtl4foyZz2Nmx6TsMs69aDxMEdXYIPpic2ioTXglGXsK5Ze9vSd128k
FyOVQG9XXKNg7VhUBqxfTfP820Ffzn7w6LeVkTVRwnqh3YkR95KNr38NRBWm9C4f
C4lhwr/noYCJ3sJ1svedHDUVYTW2kk8rsWRbX6l+SSUXQ6R+eroqMXvEuVPLQ6Rw
ryQSuBDg1TAUwZd54CIJ8cg8xwakS+PQFvezi7q+S+MABrNILO10T5hz6qeEoG3K
+DOcVh9hu/1IbgKmbjd+agoDVXpFOQRurNo5ewRnJXXDr7XvZW5Fm5NxPjQeZU6q
uH/hIuuXkwCQENHakPMucEncFIVEemAGTNHl1hL+SmkKF+GOacytDjVj8Uih/R3R
wbxrw+WF+9lC5UX+bPmtSdSYxstQnKikT9J2qp0zzSRftXQvYSKdrvC14WjmL61/
0ZoAzhiaTKq50VbU0CqLNBg9APwbjIXSpIMVa3Se4ExVni0WOj6QQWpkXeE06mPk
XivCJ4l0xhdpgRu5prwv1D6mvCY1969Rc7POrbV3Lp9hY/IHsCdaoa5qFtgsN222
RDRnqvPrpBBsGswPBNeC1UMWEMoxA0EbcXeU2ifFuVw/8AFGkIR9TIS7+7N6IpS/
LTBzPwKoBPxnc8HL4t8ZC3hA7L4Yh+xT3LCvyAA2F2CP4qyhWfX6kgs5zwBT4CVT
DG1WqlaRHfWydyrB1jooNShnP3IY/msayj7C7mnnvP09pzi+mfYYlDFNImPPB6V+
eg/oZ4ZnD79cBnuSEo2HlioYh2DDJ924bSViijAZ5OJdSTbvGPXVeKzVgJJth5om
9BoTusmfhpK84eHAwNmiDGQh/y0QpfVLjALughRJRKVgpMq1ZEkBEyIqJnI2+0NU
GkmdqW5YAhT8hc3NmRA63keqNEUQwlPHcrXR4V3nb2F7s7EOZ5o20hQfCveHyLn+
ugysEy7buB1lZTq2uStcafe5QGT+ePalItLSCBdW8hn7z0fwWoWqUAIHeIXwfY35
YMKyYXPcHBCs1G7OdHNx2xhWWq5M6xTszZcqyBDRB/f+cc7OWWvIK7ymBgeAQ6zh
OAVqbr5OAZVYg/18Op5OoTKtw07Vyw7RMRl3wPtZzHCWaVid2L1hd4MSL+oI7MrY
9iVEuoiOCQpZ8VIY7oExczf/liLyMH4OiUR+plm8aRh6Cc3YjU3h2hadB5hAPUoh
uCGmc3bc51SjtZwCGLQeyvE0TXNTPk8ae1eNR8RcNKjg+AbEDPYlGAH3jdxO8T+I
z1WG8siriJskpl5zY2i0YY2fJPZ7UXmKe318EmLOaePhuYefc6CtCOXT+iXMt0tb
bVPDkhkmrQECq4eyFwgL+E6mZseiai01OSbLlNksC1OnX2FzlvWzmLcTS5S3psue
MCDahogrV/SOhLyz24DNYBvzrKylrctTNIpcDIwFi0g3BTP1r1j6Bz8hzx/qfOYM
zK58ZzGg1IXzdrA+wGkK8MTJ2+8RtrrBbE0r/d22/HPEg2u/8kYMIvCIuJ74hv2C
EdKE6pmkRPnlBSaRRQVnwlZnG0WX4ipImFHpJJTAzmdlaF8bCHvA77xmUhw+tS/y
zfWLFbVUgfHgQUlXNyEF6ie7XNF2n+hZg66Fh3ePVvZeIHtO+cmZSig6HmidSY+G
eqAw6NBjJSCt7KkSnYWe0oYlKXHglx+wOifdcfSThITh7ACbTbYs49BzxVLbjdSa
tSWRumufhgBdeLf2UeBnHO7Mx8V1z0WhHQoY19RYAbPjurzcTZJE919xGMvl/P5k
tqImGZBJx1hEeDdms1g+Gd/8WrO4G6VdSdx7oUEJiuBKmbwyPkmla7osbZa5XqV/
94V+4A83/l7bQ4DYEXkIWvYjfy0zzoo3z72lCC4XSfHFbMGAzoUALMAZzUhRdbK1
besl9zqVpD4W60Z6RmLv9P8xNNxpLiXQc2LvyBfiPItG53DpOz3FCVTzTDsGjqfK
DDj6YMvsjFebPHsACPhC6TjTJusXTWWjUsguy0wdZ6xwUu0xx8EJ1VvYBCGJNDGM
jYdsnLexBZ6K8922TFkXKM8je1Z7DenSRUdsfdHAbMTztipiWd+39ac0KMUOI/QW
Olmr4e4xdSO4V3AF/DgSppZOnXTiw0gvz60n1CVRV/TK4MZxp8eEUSjpk/OzDJ0T
nRRgtpcmIdbcS4AwwU8q8cmDZY9g7Yg1lwXyW1BSCcAxoBdHenFoFp3bgfCzDRrn
2B5sTxCYpTywLXlJ1XAz/TIcQHLWQ5qzVcxyOhIgd4XtWDpoJvGwG9zqcCzfeJ+5
n7eLXrk3WPMlRH3sO7XN3uAy9dzWpqLjDz/yNpT7E0BpLnVIFchJx/iZvFfgSf0z
gYOkxWt/tIwycLFSbVsOgXNUObhnx443slltzIRy3z2cf/o+htAghEnWnnL16lJG
Eomzlk34DA74AJgYUPVTk8xMt+NydtyYP8PpJH7a0bn7AUvBve3NhgML3l8dnTrO
zpZwOgE4z9ABg4PW/g76/awOGUlX/uLCFwRl7WeD++hf4XbGSjSUF+aOCDYjzJ6o
eBpLYBP+T60Dm0qKGswDoEI9xFBiEI879NM+0uABb4dhspg+OcQ/Vld6hgsC/aI3
twwFMRBEh17C5JK0UHVMQ/1rUeBEivSwD2gJdXQDAyDC34c/7d694pm3evU/A0s1
o/m8xLmDh8ln8/wIU61muqmNhm8n/dccYsoqaOpi3O8A7nokWFkSYLjwuR32d8cf
+T6ifOmcxw2hLGTVvpXZb1yj2C7F82MkOmpv3EXcRwDK3zlkFv++EJPl4FMG9AKx
R0ZvFDwUM31la0ivGA9klEElQPJmURGksqYhkFX56bYa1rI4/+rxWsEHHNDvk6p1
TuGcZJ3ypwMj9vDNEJMveI4B9wKPnfIe1h54ITfz12oCiCyATsdCp9sO9mao9o5S
hhRpPJMI5O46udF+KijmdOlBit78FX8pOftMRBBMnd4GR1tun9VNgvMx1tMDQRyf
KZwDWv+vWUGDEV+Jhk32XvepHkCojj0vZh8nYLXz0YuNwRCJvp5OW9QflAK6q6u+
qcCnUNeAeUA9zTqO7LpJYMmcQvJGCJWq81MDbloNoxTQW6hP5SnO0FuMuLyg5DIr
hPuaBqiDKV1zX7NC+ZL9Bzp8wrrBrrzA9507f1sosK8Kz0L08yAdwWG522rxas88
uCDWVrQ3rqwZS3c3DCwe2SEzgG1KdckoM04MYeW+fyDukosJZfqc/lzvpamMhENj
DJuF6O4GnXOwONQQYo+m4d8L3jJc9URNH13D+k6haZ4RahJmqamlxatYYNTUOBvL
fh6xx0q761PiV26Y3gPHQX3XIIEN/0cmg4NTKDeN+W/NGA9Zjzat6C8glGUrLg+q
lzGTtxb3EqCpM5SdByjc6b2w2BjW8EK2XRXQw2xLHjFyNeT7za0ghUmsH5fSEC59
j6SK6V3eSro1Ln4/YQMElh1/daxDbIRFCgSZNLtMoThfo+6eZG/BejQsVvmniXZ4
kWrrLsDb0w7ajRWg4hai1bTKzFfRzBqRI7Jld37IiSMk2/e1ORXF+kXrHhwRvKQC
y+fzh5cUmkGe+7O6BE1hMQm8iGUKBLSzwOYw++qrMVDEwkfalw8DFGBm40QW4tSL
zlPa7q3Y8WXaxPZlJNhZHn2GMCyb3TLdw8ACiqVGo6ugSQOb5zo3SHcpwYpb0P2L
U6AlpCWnH/tFSWiqVDYrhGLCnVVx+YwF9CkjM4uVB7fv1MrV6/PnD330uRQLXwhR
eNdN6+p73Hg6KdEi7H00A2hKHA9Z0224afIqJaGGW7g8KDUYwHjUzts8Z6IXiyzR
euIXCLR45gc/9xBmlFIx/tGFX2ZK4U19antsOJ+FwRsICMg0o3OVGRWQEDcTN75W
T0NZfArJTBkE5+pcF33LYOdzDFya4tmnCmMm+t1q1EOTgluThf40AJZwkNseTGKs
0G5wgzg7lk3UAf5OJPlFYWdWfikQTqczwSmoD4ffxQKAvR/LnVFH6xvd3qT+pFxY
q7jKiZrJriOgEIw2QmbthYAaJU5VEhHTGQ+h83yBPL7MDR53REaDt1JhTKzT8Vib
w3gZtRpPBjWT+A9C2zxwZXmWDpEHatfvIGXhxSCPvkgRiACaIxfemCTpXmvO4xkh
RNM7nR9hGI5w8dMvt52v1djOQ7UkPu0StXEpAwMFusZlc7zT6hRAh9jOaD970u8I
qkX6zpmBKF/8NCEsOko50Nv6XwdBsEtpzw6nfZkY9ukXjmYE01Hh19D4iMPV0ffS
y/LqwpIPkpIEOYBlpE1GiA+fq6GRKvGCP6mwEWQ+lEITgG/XXDleWVok9go0hb+U
OYraUumuALLtHGCApNGSvPTlp/HVnnsE94qubaWW6qyU9pj6Rt+dn+fuu5P7t3vm
y5GLVSEO6k8ReEZC1+Kyv07XUruEBLB1dPKCOtHDFx812xUSWZJyQMoFMfi4cSiY
QcVTLWCs3ZxbAL62aJZwzuNNdfOcLeqAakTyvLSF+uQI1twhlfYURzyYw8Ql1RdB
bjlSXQ5MyUR4mVw9AxiK29CoqWthB+awAEDMSSV4SRvxbUcRdG25r12nTP+Sy16J
HjGHHH+vPDxuUZk0RMbQB93QHV9Xw3TaATUOn+u4/FgAdz6xCF/nCuq8dkW6GBGA
1mZpTaVKs85FrlC/HPo97Jy7Txc8CIpBKi/Fe28530j5tURJ/dWWdo+TLc7Zdc2A
7OYbPB4JpeGVCA9FEc7utA7mn7nI0LuojXqUPklgR16S/3TTw26MoHESMNk7VhEN
4NtZhfzIEIDenZ94kN8ufnWCJZBmNRnanpaxMGbW+SgynMjh63Lm+bivGUoCUsKd
xvEDHHAGJ1U0jrAL30pWiJPaDJ5DloyNfRnlrtWDyIUhFuNX0EkJ55ZlZzfA3Awf
z7aQYHs3NWrjEX07mgc1Xj/pTRCD6fwYCbAzZVug/rywidRhUYD+TQD4PwqOb88v
sIRzyt6myYWHi5QUdOFOknCc9BQ47E8XFx7JO/DU4CrXBzIo1FMUrwHaAfuWOm67
ECuwOzTwIZWDp5dL+nIx8QcLy/4ujSlMxo5KDDFciyp3aaMuFpzb6YBSOB14w0PH
GWpaePB1aAg5kRMO3wBKtTAnymGfb08NkHUXwUPh2piMpRHWzawOn9OdG6fncqKI
iLSIMMMkyENaRBn8JAXCsFo5QqCtfoZRY0zjgnZrfP+Nmd+cvnEg624onG54GYvj
4hI9TcHgdhcpl4Yg10MnAHSGia28lvZtumgwrsoJNSE3Tof4WXB8B55DNL4oLHgG
RgoqDi2ISBQ9R/ibCdADSo0l3Nx5RY+gecoWG0+Ac/kMKkO3zU//HEaJC7lPskcb
fDwI9SR2tHqXddpvVVHPH8/9Ok/djLTjkTbWT6EMQIm3UyRb8/DS/0CutkxG7sLT
pISOmbtpo5nlf+bRygRMHNMlRTfv7Stue3CJCvHDQ5FKM5NQdJjUwbjo9/heQtDY
jhJFN/rw2cYDN6cPT/mlUOCe5Qe90M4ssU5ZRBUIZq6BrS1kzWT+TvgJfINDIsgd
X4XqE0LDeEIm8t45Ne7y/1hcjPhLjIU3KP1uG17zlAISzVwy8xjLV9ti6aWBlQH9
NZt845yp/5GqgKOfS76jWOGMI5NPZNRN9utWsavlS5XEJ7jxyklMyRPrLRmuXAa0
9/+zRY4VFJZLyAp5LIaQ97aahBuD91RkG4UOBZDICtTiBt8ftFvAvzUkzpbBDG1n
JRU1rYmCY3M5ELH290I4/fHH6CqzWNwiA5Mls1eBFjs/bUjA/jjYteL19E1OmBFl
Jr+lurqRwGyoCSiFVrr8BaGudNh7n4ZQbj59SkzFI7/sIz3Z2Aux6Yn29htVE4HX
4u0kqqU8/5JC3dfmF3tuwjqt29W+ovR5kCgeYxwb11rI2XgZ6nXcB9NYdPq1VD+h
h+gdj9E7+VsPvGXye22WqPH/XvSnzRApwmSyOrPc/F2zLn0uAG9TWKaVa5Apj8OM
20INWSDPuOOy6XBayzclMtyl1rVkRTzYStEnyKI/sqh4MwEALL/InoJZt/wR0ZEC
yxhrGf9Xti7A+lbeHZDOU5gE+/nnT4UOqIdCklr7LHhTG1ORM4+HZ3XzF7yJcdPd
p/myQ+cq9uQ3J4SEiNxK3rcUVBFQa0Ol355C1qLGfKsYFvXY568qsp6b9xFF0qEL
5Nuo43XGLrH9LrO+1cuqrxpnJQgSyMwps2SFlQC2hlxY20wYW2gFFb8qvfbTjOsR
hRsgMdSQ3ix4MeHfF/1SxpJxKRuMCUeKmFgFJp4XzoHkk21rQrb0blr6k5pF9cAJ
WXdnK7iOPP/k9z4uISOV+mZXvdMyZoasSEqM02pDgCqCq04PGLnYwsLxA35BD3J9
tNgcpa/zyhvnHqB+7qillD/V2w7rztXWBafaqRH54M+kySAwc6FX3DB/iMmnPR95
XG7y3hFgNEwKjwdEo5f5YnufWyuYB1lZ1+YZFR+7VTsfEwH/j6f6ENqhc+8CW8OS
7r+9rQaLo/L3nPpNR4FReHS2xf6C0ek1i84rN/Ce1pp8z1QG6Zskfsf6DYg8CwQx
UihjB1bzyJUZ8MBoE6+TqO2pk18eWIDwzUdEjQj7bUoRZsx/uQcfzskp8S+WA7sQ
J5op/atqvdNMUBWMM9bj3ELxP/3uaKsd5BHG9RwGruk9cM96ql0SF8gXjLZw7CCe
nji7oedFRHLf46wFRxIuRwIneKEYRjcJ8hJFtvlS1dAwHQ/yg/TT1gSXIrCYAEWg
YymBufAHeBkOUISJrgr0Mzn8+vE+cNTJhivwxx4b8huAgfEGIIn5wNf1+aATHiVb
niDOIOu5qjKOrOb9s49mSqrx7fiDW5/aAe4YMh+Vd1VyPPoyBRL5f20XjuSxa+Ea
24IuuNiHfqE51fNwLB0rm3r1yIZ5HCIkrZjGXrlhBmg3szr5CC4Exe+7O52i2eVv
Jw53MyryyuBuVGEIOI+2+znN2lefLfKjEXADSUFurlV18Y/2ou0GnfuvtARxjXA5
69Uqfsb6UmgTyeG6r9s9u8yTcIssqaMp+J9MWIttmaGVpHAnielu/bovGr/A+Epl
OkzJjvHacVW3YoegXLc+/4t9UjO04Uv++UDL2T0bPi2WR8rwia110OMwJVgBJFN4
V68BtvBvyNLK4OgN2jEqkbcqMK64ZRUgGqGHjDrTm/eDd5aJaPbBSbJO0kUJhLE0
HiXVIBrF9mnzv8vCvoigu2hX9lC4qY0biF39yZJnJdAMmE4nX4jgzTeMZPLDoNRC
Qh0ui3bv7n3ocsY4LLRGB2EvSFvzNkaqcuWG9ir3jygOrMLCPP07y6E6KEU8Nr+4
9EO5jtGaQveUXJyRtw4jHL/QLi1SDDK8gLRgTNvk9RGq/B+Mw84dX//W3e/hFJbp
kGw53jX2jJpc7s8kTJ6/dYLqR2JWRnAUpfARsLSOWMVBLucBFR76keENN1s9UCyA
rJ5csycRPNjSpyd3L0cgsJiY5ByAOwRcJ+nz+UWsX8sAvgS2ei+5dkSAnFC+7UPh
oKuaQmkDxmKbAFh6HvMYqLNvXCVz1szdXMF9u1dG6f7EpdJvpV7NbjiAjVIYary0
8ol+8VpwBWzbls7mTq6ao7fhnpRLbGTvitCxl+6+on9Wod9mD24cuZweRhnH1cSV
3fm4YkmEhTMTDGnGSEGyVytXkFyzNMVcCpEJF9hGLIptm0Vt5oAg1R803hlhH9+g
NxwpKdFpZhuYoIygyf809pes+k5g0xA5lfdob9eOGEYmEf53QyzHLAYtUTk2XYLL
Puvh9UU43SzFmygeA8Q9ScXczWO9YbcZt/2A1JG7SFq7QOHgSBCT4WRqAOlnQYar
qtU4xc8nr+TNj9hgVuZcwkEXI2gWhpiMfamvKTihqOV53kja04iFTYoIS/4IKb0x
3szwvoqQf2LD/uDLqG7caQcFWRim2TDVpq7IffgRKKLmbOetqkMPiFJHP7kZ8sKx
zxQugsuBRI16eayNOtW+TUnETWcTIqgJIpaTBWO7vVlezIq2eMLwgqfxt+JNCSf9
rng36d1IU/WarI+3QlGrqh/HCbjcVa+5cWI/clQs15VSQY06Wihn8jLpdLF/Jem8
8q3WZsNxMtf8lDEwcCN+U/A9emrvO0Vf2zt/Gi/tqf9nrWUvflX/+5OHInPBosef
rnTegLKeR0qQH3T1zuQtEWJeKfYhNsO9IiWJiHfXeOp3bboOAwomywwc+PnQ91yi
yqyPkkRT+/3kBj4PSbCO4sI4g2s0ioVcm3BbYsNaJgvNki6pWuIhRocX5HY0QX9g
4CJdvb6/HGcCZ5SabBo/nwQJt0SH6lCeMVx/8M7uWqlZrT/u98ussmwnfpfxe70Q
9/YZWtakv0CAAuNuPuf1ivQHYiqN0ZomnYdcKIFhNWuRgrq3tdiygxq7R8ho+4m1
OOzT7C5ZSkkwp+YGzdkYZJvFq89b8lNBohT1eEvk2C/22rZCWLEw5ywfs6ZUlkIx
uuh2o0qqSvEebRgUHwjL608+yINQwC3nyoa4RNEN+ZgKPVxQHmC3Y/BqHjQ0Bc5O
xbaq/evj+X0DjJymSM10xZUc6tnCYeyskfQC7EfW11k4FHV1vCsFlq9ekgbZ0qO9
VCbdqV45ljzHPT7+ILbI/HAGyNpNd+JuAsX4UsY4OzSiXBzCqlC3reZVfY+sRadJ
cwkrXwpgdJDl7Md3sjq7tgy/osNxUTGh4HvXP1LjvcE2zuotIyMGa6ELiUOXe3S5
T4cL5rJJjjf7zPIxrR8TwIV5gKv5gq/kKMVtiRFkDliyvGyc78aSbAILriTESdFh
lQVs1gl7ayEOOMRVBlRsyf3WCWTfTJ8oxv7yqnHY9Xo3ODl2/9hFPfSfmkmhv7U/
gzVJ/od8Zd7WY/j+zgDxj7CNcqKVhkueQY8Psbwu2b1Fhxz+/7Mn5FQzRNripkBb
p0w6twQ8aj805qYrgu2hy89QWdYw+BFBwFBKLpwzMyFcuoIz7dhH7iVjbQjv5VNw
GLuS5dsqJevCCk9RqzpHSwNJURkM0BP4Ba3hGjvMLBE804zCQEZllU94Ni+5Y9xw
yx0ql43/Tn5038ZT73SCLJgG+oDgSFn1ogrv1NjvRhcuFaNvMf1abKYOb1OguWqi
1zhM1JEzEY0ryu/Fvo4d6tjatXUd3csTG3h7IsTZ1qOWhLmE9byQZjQAXc078Mtg
RYPWHnz8sHY3VvHWpHk3cHPJBTT0oIfIFfjJfizq0LTQQUpJIs6/lSEnP3imVq44
sq/QzlOmrLXrTfKAfYTcbUQ3Qp2F5h9FkT2Xe6qXBd9O3dhH3PWua6mYJwSP7EE9
/KaMVbbnXAN7dVR08dzdZNg2c3mh5cadNs9s2u+Y0e9AOujDbN6XniiyGXqJ05cA
1iyfxBEwgZm1x/aoKuisAs4yau5bHn2lwOxc2IMUVe1wYdAgId1JYfXcdwwXRUzW
IBucu2jcg+kI4zyqkIH2GIeToB3bwyV9ko/tCvprMFJ18h+M/bj5GhZEGNRWsiZP
SToSlvCRERqwOW/r4y1CRaL+pu81/p4Rm91qVYOeJA8UgftyRcvhZnBCaL9yCPrl
rMbT/dI6+QJi8MqXIm2RQj9Dcz4dblbRykCtKupVXS6JEtdu/YWPSGvGZxXhS/l7
eXIfslXSS2OIX6RMW8JKlrpo2uJ5oZsVlD+oRydISZUGqzcKgqs/L/na6rn0KEXz
CzwHsw/leQ24So/VC3FWMTZJRsNga1W+UySyNaf0hRHLRmoqkw8Bu29bbGkLAsPY
cwhYPhyani10QMZb4njZSKKLGCucQNQKpuOwmDXzvqdfMDSNtpSmven7cAnKYOWj
C9V/zvQ7O2OZs+vq11TSNj7majReOGHF0jFc1/HLtK/RqWln1CVgsU7i89pExRWc
jwz1v+okEwQQG3aPpQL4P+87izXEwqfcEJF4TY9Mktxto5UFo5pTbRUMHzuVy0Lz
xK7w65Rg3GtlW3xBEI9xO86NjfsQcYjHRiiqA4lFCbfyo4c2IdE717uZNm+CWMEr
aI48dlsB5oZtLmO8fo4A8+ZosCPO9TTQojOnOU6Vx6wA7r/Iw98DPmiji2Bh32aK
GVCyMRkHnhWILmNApnOUx5/OrkwXzsVsONx3vWGv7jW72L2DKA7t3TUPjQlvW5Fn
dY+pe5F6iqaupEhjIZnTHFrtE7xKZFDUpxKQq4dAifjbZmxpTBa+Oj5mN3ArPnws
Iy28wSZCjxQZovjyzUeVOn6Jg3hRuyE2qFlhg12fbuKWdGnRHuCuvj2UvFDjKSdp
Iw30sdj2KzsRFXTig6XDnzZNnq8SGIRa07tPt4fd7F30XbfWVJciUFIOqX1sG/nB
YUBC5Uuu8bvaA9FVQ6hgd+XutNyMVaXxlA5WQNGsGgugPBnJnMqW2HiRoYgtk2g4
NqgRJMpd3DnvJvE/ZDD1zlSxEqvY1o43w00tD3Z5WrxcIJmYf3owEf+OfXECGRwP
ywzyM5Z9GZYEpDzcbfDaiPtVZUpVcMzl2WKZk7gs07hGOgw3SIM5aDl/wXOHbgQt
+7IClOv2nFNdL5MYVXvDMDMD0jMvuCNebX1GZmH1KO5kLXlF3ifoC27KhgoYqeSf
S2utzYwiEPWo+8CH79c1pkPA6O/UOsatFEWMQ6742LzM6ZXRohQvZqmcfXrStN49
/wmo+8JWZOptp49QzYhHI8rBKRGGtk/9XPKd+OasQbD/TuYfzeWyA6t2e/S9yS9B
mpSTbcbJZZzGgqAZX3SoCQnyReipv7TpvdU4RuJC0yBSZdYNmU1pvS7bOG341KCt
8VTATflWxiMtgNb9MHt9Qa3/rjKm+tt2hXGgeJG998GGphsaN/wczkJGTC29CIUI
D4TsY8q+/V2sOBP4dWEG9+N4aABZK2G3hW/b+1uqVHWBTDRotR7BLyP6niWPE4s2
mdu2SJC4rwuIfKHb2BlJsUiSrtE8dPmMW89sRLASAgKJZ2s2oeRt/hR+Eovfvb8/
YdeVIDfpZyeLR03SaAtJ9jNFo33rz4crqvErCuG1C3wLK+W0d+9iCm2PhcVt2XD9
kwn1QYns33G4D4GA5mXV48vsop+IwblEnE8SJPOnaJfLzkwwidB8xeCKtvom1HI9
g1PKVxz46W/oibhMlYZ4uEq2Y5QDu89bYVCtnFRJvWsILQtKBhCikiKZq7pR+mkw
EoN+T5SyX+7sUf/wm1AtlS35l9UUP+wu/tykRZlhvltqCAerg0Ud9mdl7SJX6qiu
HBqnFYLp8bEYbg1Ej+1vTFJfISRVrAOl/LrT/o0L7KSBbC+vk1gqegAqSMav1xHF
BxVl6kjqfNVthPE2VBpSvu9imV7AuDKAZ17xE+rSaN6LOBEVFjg60ZDgppJqJiru
cgNXWxrb6VQ08cHdc7r4C0BFuHcmUpg14WVvmejZ4gvILVlQystccgb2ciwCp5yj
ZQf3SLiMX8CSBgZjSBkJpnYKinTe0Re/tjx6goYRQY8gmXbV/iXUjWlCwE42BJLv
0ixOpR3zvkeJxlknVj7q+WfJQp2PUAvXDhNZxirzQQ5CxyuB+XmaHcqRfYUwPuqI
legxYWyny+x8Ky2HljJvuMpYEWucFJ7OFa9BJDyj9KfIwcDZCWjzd4nqeFXd2yOr
/JK/q9G1TnDln61Xz5kSBDvtHVT8CRQ/h4hUVEbOu32YkAYsRDragxXgW66Rf9KD
lZATTREmB5ghOGnTZR0mVGN7ySvvljkY0AVWLDEA24tW1paF45oPGd0suxabwbIO
3cnz35INDTrBI/VJl5XzCKMn70lRYCVm1khDbPSutKqlWXIZewhg5GFp6KPyrNC1
bJpZynS3SlksAk3wGmR0VIEoHtyJLGagnpCSd+vx9BCEA1obYEsXazLj55cStZ+j
sbbniM/NHhyvvabXRN355GIdNRGPYvKuXhuW0RQfddur2l0j6vtxwO8YgGAwQs9d
UQk4wonyO9Ae0XIsAiqBZMrwPf6bwP4mPQJRLxwm0LtLCB15BdobjAVOO4y2E7AH
uGmACpDubbsOUBNEhd5xb+OM53Rq3hqj1VjVoQvHkCGF00A/Rb4VG7BDQY1cd8ct
nebAWgUClu/NT31Q8tXmgR2udrG5w3P7fm6fiBkSSlqbrsgPLrNrQ+gIuXSACPka
cVXaA0tisut7euz0QujUFP9mJo4TVbl+aNmr7xxajO199vVscN/Ghp8K0lk59fSK
EtXlaR99zLm2n9XvYmiAdmwVp/t6szpcFL0hwKKx+HbpGIlx+HlWfYqB8qQYPks1
+Zl9p5utgGnFRZ49xBv22WXjDCuyQhXu/x9tnu3Co1UR1JRIsW/2VurFMRtuoAWM
NOfFDqSwzmqWW0iEdge7OHoE8pn/ItjG7sqLl49FC75JSahRH/c5wM+p3+6x0s3h
sBMIeHKC2Ikq63z4059ifjMbNbX8r1JyCUxM6lH6trbhRvxEfcZPbObbykBC6B2V
7S4JRJM6z6cKkZ1Yofur+iZkCDrD2yQBxVZSNBdL8fsyz0s+3Qg9e2QmcZpoXg9M
EW7G8INByAAoOp1IOPWfXSH8x9ovg+NI97UeOhx2IVhoa6TzvbbJM/8Lx051hWzf
EriY1HFmgcf2jRjJn9ZrtzJ5dRXHAL/H5EXTnN/5lTwqBNDlldqLfUihVYF6iEIj
Spdx6dJkgRbeus5hZJ+zYcHWEK4BBrYXUbEd7orffPJiQnht/JrGdoqqM8TyH7ah
povqhfCqlRN0hkm4XewQtGDLp00yG3SVVHcuhrWGG4dxtb/wBtCCblgL3pU5lgsX
K5/H4Mnn7CaUCO/rNjSlVcJjzKBwGdA5W12wxqb9QlgHYikRouuEcdlM74xO019P
tsuYSb/cPv3dxg/QSMAJ+yG4hNg4F4/8R/RJeeyNa4YTxiLXHbwk6FCLmIVwNV7M
KTUH6xrPEBWpwcIZOSxXIRcn46MJR7RVoEagF1fZV6kvLAaruM6u04v/FmL5L8Id
QMH5UaQ0GaJoWrRbFfxQz+EWCcfqpscYN/gbn8iSbRE968LlfbzN7uJ71myPesRD
zkf88mjXD1tIUSKUr8nkZP9fVhNEabS2GmY7PcVm+ZaA+aZGeU1a//mv7q+z4UdJ
5JW2iUDsI2AsdRyCbNqR567RL7EDDq3nES5kFzbOc5vc68aGDGHSlNnfcl9R83On
OFG2OqDmxerHNZOCMjhW0u9HHNkW3BsJoZS4ilNbCB/gc27C9C/Kt/uRZ7fQbtRl
iSqOmlwuHwacba21AvdZxvdmapyTqCueB3CyVEhSFfOUvh4O/NdrtyVXNsIWyvwZ
pM3Qu7qifoLS6TaN/LUS7B2DRXQLSGNYrr8YcYZhBhVUScj1oGUumM4fp2Q2zEDS
KUUaH8jrW/Ki2p3wBX2H9RmRsbwu5tzvK1mPanDaib1mJ8kfUq/38RVGJH7nlyBw
wFVRJzrgJRbZipay84pV7ICwadPAEW4VEfgUkuohlooj1qdIoYnUKqDQuyfs1DNS
KK6iD2RZQEuX7TlvzhDqG/QHSVdv215/MNMt21712jAFGqur9KgBU/3nM9hGpYzK
I58VlXnp2NSDb0FnoSvPlzsJp/tdE+c42AhiG/JKGBTPWqZ5FZ3S56oSRD1SjO8k
gtCCH38T7BK5LtmpEuvSY5RgJlOZlsRSo7tEVlhrfPvZq1fcwuwxlFZ2tQFt9s4Z
ca4WZNXpLXGHiYi7b1gO8tIxTRM+nLcUlqtREx6/vDmjnzEgQUYJlNYsjYIa4por
T9Qk44FCk2kgYeUQd9ieBXAzS13FeGAz30xtwjhN5oXzOjt5UDEz0VoIGQ6ptmvh
83El2bAwhwgAOUqvvK6W2pn1uglUImZPXzU++E7CDQQPUt13UwIsJ5+w4j6kmNrk
utY6MvDqhcIxJl0gCT9v83Y8DeDvA7SHoMB0Z3Ni4EFHZLL7QSkPir0UnsPcwhcr
mKwLd09yu+Y48wGfYg5A1kQixgo13olca/+7ywcRCpFd7t2+a0xWMQZP2Un9a3K8
hXpvT4jsghByheNdk9BZLJhicbmklA64k/rCfxR+VlpX90BeT5Q0N/KT0lLQhQ6I
6tFxc62Z4vLJfvitmiddOKrxb3Sl/lcp/n+lLgKZSEEnyuJI2EkGrOzwGD6Brp4G
onRgyH8PWlFuNseEE7TvJfsUSqawLQKYlYdy/kFADeobxq53mMH8YEHTGthytnu3
WZGv+lHHEV94fNyx7zcB3JX/QEUjLZLSNPdAYm+cMSTiTJcnhDf4Z20iU+4dcZr+
Bthurz5iHxO7r/IAeRgfo3GVKwJqZP17ZbshaPJVCRSZdnMREAhPLznPCUxvWbeV
IxLupqKKfOT7HyyVwancFr6T03ZzF8DEU/VlXl84I6xMFBbqQupeR4kxrwAE7xQN
LJs6bgkBUsRsBfoXKSgjpiXOMSGKv3cqrcNvP9VDQCY2J/YN4Z6gjxI6oNY7D0Ag
6GRQKTgd+RVWs948vR5a+TyBfSrjglKb+Z5byT/kvpo7PA7d1YZwRcT8TRRcqIBv
WkOQRuW7uB7nLgMYUcsNd7bp/djYAqV7iUtuYumbGACUaRma8Rs5hdYIolG8EOuS
7Pnga0n81uKAFSunuvNQlWK5LQ2FvutwAJeupNASO2Kcowh/40RZGvG4C1SyOOSC
OKnDpj3iuKpse/bd0F16jmLpLpRrXPU2DVU60fV8tfWTQUMWhxCDcJ+p3iXLsjJk
t1SSE+vGa+jF2tonOOvQrfrjTzVkebhnL5PFg/SLghYNDiO8kNVmtpk6iJmTwH9z
6y8erqGoSWewEoSMbnTJktNTaEKqBqJ8rYazAGodxnmGZKO1d18uIxRiiXjJpRhd
OISEiTobrOmO7i68X6kZuJ+Ds7SEV48aofPQG8qL5d/zpNpy5QHujbrAaa9pos0v
EktenNcm66WRRjJVxxi9WKTwffmWqPFF3wQEAwiXlXwyPVeGfkyQWdXGF/0RxpDH
URfrtryxxsZPWWWQgufvT77SrpFJ0C8HjEw5uN7vU8uZEY0mP1fhZXo/EK1HcW8C
C83R0vQSJTIXBk9clJdU+TCKlv0ItwKeM8bDaCd3YcJNNVg5Ced0qa2DBXI6Zrxx
eyckGHq6ihw+xVzoHa1dmoYt4m6eZgHw7shnN9+krubGycbBMEm7jt/V34UAhUG4
vuuH4dTCoQdkrk+iJV285ORc1FLRccGs5e/rsytJMimnXRZAQVbMNhIanLbn9Hb6
UMVoD3vmMhawbBLgNS9s9kh0GGK08Da+BGtOPMv7pYXOAoF+RQDYZ0HeISbJ7asU
fATPTGscLGDxg6dMY8r8sBGglg45/EjtNwHGua0GklqGPyzxNp3nS3s+Ic0mp0xV
FppqBqCjJGfl2gKqnFg9dLpL2FpOdeetlD1gC2DgQB8Dq4AAgGX5K/LqnOhkWkVR
3Nu6M/V6W35c2o0SEwyJhSWDzxO1P2cuenGC8qvG4i9ezUgzUzREv81xOx/ygaIq
zyF9d1bbVO4ZqD90Y6DfKAwSA0iVxQkCXh0XeNdUU9DjQKBmeKvUW5pI9eCk1+a9
7TQgfgQL/j46bk/NeJKWDxYe/2ck/aaDvnbBvypNrG7qJwjn9ywKtshMxEompCz+
1rnDFmFDlnXimtWQdOOhzivj4uNlXUp8X5S1me/yyqoJc8+EfD65k8JLQyVwBQVV
00NrkWOPpETn/yfscvcQa4ZmGALEQ1KVZU+QmENtnKlcVmcrrhJMiBe6BRSZRnp5
XdQ7A6NzcWZMgi/TVE8YQaSlg2uEs5hMK/yvF8mSnCmsopBH+1l8w27SNd5TepX0
HOj15BcmKFaolVsnFZkp1skBWGP+BXiSuAYBbpI9MuzgjphQq7XZnhWcGApCxGnB
qzLr2+U252KpGaYuDJOLZHRS6As5rpOf3EOcF9szXVhuMD804a1+TEBxgOkRegPr
rHbRtug9CDMP70hla9cROQ5zrm/+P1WjU44uVejEAANHcjgitfYOTi5OsL5EnyN/
zKHnYqVpmwvgvOWuBXrmGVUy6EPO71/Yci2wrWkvRtqS+9FV+xM7W96QeWDeIa6+
3iPaTTRp/3RpS6qqwLsheG1yF+DUw/W401w8f1OkDZYRP1CfCDA1PHHjp9qpyX1z
6DtS46jAliSbQuBlfCknomNgt+TPu35roW3U7SbE42Dzxjqp04GIsSgDdzjo8NNj
H20yzf7sJHo3Csi/eZ5BSqEiVLw6J0TSA8TxvbpZLJ5/bDUIPvadTZibsvP1jcr3
OUVxH6lQqCt7sADmS9pzERCCn4KIwmfqbn2B5qF/n4fPUCutYG7ttv8jlutRwicy
A5GOYKUEHNDkdkw2tEJFjwRqXS55jVS2iEVggpmk10iQ7VJkktRfMfY3A3lNqBvl
rid1ZQu8PNugyyqYOicK8q/Qv9rX3dEd7WN2pd1wExpNotJGh9hNd7RSVfG9h1Hc
10neJVBaJFwohT6uxZ078vo+csC4QIRB0bzRsq6AuWx3+hRhXu2faxxccWOsehb0
ZbzXWkrtpYzg/EAEl2GFl5bKGNOulD+7ZeJzOpH+nLN1hN68pvsMODUVIEB4/waz
vNZfRv+5VNZb350tJEs9Ny6zfLQeZ+8OB2zbVdNZr9uWWR/SfeJ1zCJyr+vNOFN/
ftkhHAr2JNF6Wn0Vvr9cijunCaFEIkOYRI/IQ5MUx2noYgsA8DIZiZz7WCkCE4cY
waak/BsxO87WhgkKP+kTkuXIvuvzusfP6vERC1NRGOl1C8/UYT0fPKgZFWT0pPMv
1hwDzSjkWp+E9PUW/ftawMp/F8KYjiPtAur/lnwqy2ELC47zulxQ3AP9xllgZazV
mmIZo8USoVXtglknnX55UCZD0d7nNu9YPrGEsYby0J6IRH6Q6bntxI4oUzAtR1uL
KdzHuj0PadG0Wz2gnpANebcF8Z5YIDSyHq9wl8/DLxQDWt4RnwUQRNc++QUMLk45
hdglbhY+kYVEq8yQbFp81Hfi+DWurS+b74fbxaFX5bUD4j1MOK3WdbnCIgpdXP0r
umbQpQ97HucTgjmfbFINLA8oCcCNhoPvfSsOmRbqnmzy4fs9r5pbDrbJpMGzgLUx
z8kvuh4agrdFWMUbTKaOg91NDcjroGEiN71XOgMCM5szUQ9Zxy5xS85GwQD6UsSy
TQ4IzraMN7ESIlpVAoGcQu9asSv1aVPrUhYYeAO0A9y2u8n1ypRGXCcBnojgdAnL
H7+7ehO+jx/UWhmsT57eSLfToNhq9rACFR59n6DkoQ/6czOJc/rBOuEMBvZHL8+H
62oqdUw7asVjLL4S3j5gQJXCO7mzc5wkm0D3whiLXh5M00U8sCgAraOFcNPfgspG
qi+C/JntXskfEMXgeE8WKnV4SvNaCdyNZz2eXwDkiHMlH/G3Pwtmj47Kd52YFz+7
3aYjRIUrg8KzCn6+7SJ5qIhmWnnjOMK4nJw0WMYq0G2gdyMaVMwl5wF/VDgYDN/e
cvUXuQILxmxP6var1+gpSpsxqp+dhVHVZMLRrRseAeoPuD28g35FihcEHzGoROpi
XlXXcEJqvmt+omyTa7skRao4XLiS2uxspbzCsUmmr1RAHae3t3Qswb/Q7fJXAeLR
SxODz5/uooVwjLpRXlAvhF4hVmDRzCDBDFgpDKeBU24s7wOsbL/ltc7jWz4u3BlE
PTqbF9ywXDl3sSrIiUOuc3NDwol4SoCoVIk7xOIISPZsJTg+dwZ+XD5etxhbzuEW
N3di41eOBztG5BNMK15hVabDHaJK7ifuf+INa01Yu96UmJ3rYbciMj/e2v+hhI+A
RMggWuiY9z+j4c/hVd6OuGklge7o0QZ7jP28s0+JybW3e4TM+i/Q75MYXTyWf+I4
ydCfdZC5yDMDQ7QW3zmRq598qdEnwyIDpkVDkiINksfMUG7WksZn/Su08qnOG6h+
g+uhhbA3M5sCM1DdNX+wzAZ0LbAvQVsx5cuTFwlSDFE4WpP/3a03lp9PvObjQhiP
iMQsCqsfiQa2tRbF2wHn+U7YYDwLLjIFJgU7L72fpezgBe9B1rnBLmxZYKrLpMGA
kz0WVFfZhxlrmIYyhdkEuJae4+G/bFD2gLzpQvkcn5mcDVp/gZvQLFlxzz14C96z
jLD2VB/iJH8SYJw4mZfQe0EZCTeRr0dggiCCfkZ9X2tVXh1uKl7j+VubGyS9XqH3
UdtO7qgQArEkD4T3vj77dayHw5WzPC6cDxYvxQxFIA6WsO9yXQ2YkRybZyNJFFub
eIHdGDPbI4QNSXjTVE53EkoNWnvX8tYi/XC9+wUX1iVvEZP3zAb+90+V+SeCqxZN
jP14GjkRwNZgAlrjMx0XTE7SuqSLTIHzwdzdmviXda4p1kjXqyVmtgFggubm3mdc
TUGSO6+B8FoBt2x8OrIs6IspGFLPQjkjsgC5qM/RU4o1bRyWHrf/LmViAvSb9UY8
6XidHkyK5Go4S1cfbtPWqP7iLHcmeeDqIhV0REWMT11MyYjZkGRfk5jgmtaNKZRZ
Z+RXncUDnGQ+ICislKYQrVrCgmuy1zoZWZVSkJiHstXRKcH6oKOD9hUTjrTzmFGS
qyxYn0JmrS+oVuQhx4mZoF1/rGi1sT27O/Ey8O1wNzAVn6SMc2WEsPymyDFBiWxq
6Fo5GjU7Y87d8YKc/+0EGRSrZeirKJ9ieWAW6jk/Da3pY8+mmJZTmtytaiN+QnCd
29+5yuA7Ak1AjtLfJhMetAGWczkhT1o2gZqESp4TKBZqVvvFBFkRShaC5AA2+8C8
EtAvFzaQ688hgI8kY+By0W5kCf+Do/rbRkFGbIBRmjv0H64pijmP7xCqduOyUt4q
UQnG9nfIabb2XDT+dXpvala1Eeg6haCCf2RU5BCKfdC/hsVHc8Nb3srfLNRxrPi+
E3zgQj5vrhsiFKLxy4vrS/Ng5ukWP0o2If8H6Ov+CHUQ0rxn/XaTG9EjyrChKw8K
JGjRVe6gcvMXcqM/LX+h9CqDJitLXrhfmKwVDqWLXrn3u5JgM+ot4G3Rlx7WHzIf
wudmcbo/3d0aLqAostuUclyPaKsn4W0aD24/0c5l0wM1+p/UJAMfkLEFMkpSdHZY
wWzFrjF92P+JZbs7UHIxPjESJllLueHWH4LafxO3QIlCaJCbILswYW+QM7Y4oyT8
aENRzgNmwhXqa1LsUVEl01+Uz6jLS2mbHr0/eXYQCMST4sVfCB1+Tps0aNcEKS+y
zdJumj8WV557jbk8Sa72/TrTiY7CgEfaczyKfKilWvU9b5eFkBrKu8+C6Xk7Nplv
+rX3FqV67hJo8HMgVvxDHD4bHSiiBq1TQD/b1Sst3h8Yx7xRBNZaO2gLA3PS+7eH
GWb8H3jpTfSS+eP9pQ5yqnBiV8DVakOiWAp+5+Y267kReTxI6UpD7srrPLRlN+OS
66z5aA4WO7jZTlpWbGD1kyCvZtPi415tGjeucmHSUKkFk2cnL/4R51i1aIzObiiU
p09V1nU/3L+gaTB9qf+yL9YiJRTs2alRMxTHy6euNRqwy15mMAz4npcq/znCG2JI
jKjKPIRE0BpcohlN+4ce1QwK4uFsChWqlurtYRG2BlO7Ht/1L9v0jJg2kWvpwuly
YsBGZKnI3bC49tfv3ng9gwmLh6VZQKxS6QdtLeVLrp/ADnqNPODjEHEgbwOZJ70E
lK2dNj8EOncj1iotcwppnv0pQWhOCRjPrvXlq/6nz08Z1l5B2QH9JWBgA73JrlFf
4SHA3XgsuxzXyoW9McOn6rXfLE9/ON0GSxpgfIDYL9ES9k6a6KUQxnhmHdbbqV1S
KFUkrGIuWy7M9gMHThNo9BNwpY0+Hu5qOZ/xMTWnhl7jSSADc/3hf9zT7pejmFxZ
VVh/vOx2bLcxTpTQnolfh2CzOzZv2H6pZXOY4/xrzqQiKoO0SqvIVknUstM7N2kX
Kc0xHTRv6ED+wrzh6WkAWoPmXcjTV7p0uaOoqLt9lHo/acA5FmW+jz1HtfHPW+ER
jcS4FaX8SHXwjgh7BKheWK2WH8a+NJ5C3UamT0it71MKOkJ+UaKBOVfbqQMbCPcM
kJUV+WHC3FKEUKU2Hzu3/mtOqDfFh3UDTOQu4wR+T9XpzNJsPRtNFtODdZlaSiOO
ckFvK2FiXkMcGiFSjJhkfdJKxmOFsMNhnRzR9kzqFzF3r/lfuNJBfqLk21kqU5LI
FzgPuAP3N+XNCCQuUyuncBK3rbEqjlFSB9VuQzEmDzrHHmGl3Cv35LURaw5YD32i
Nyp7dG2jouhRw2Yaq0oSJIyZIUX2cIHFCfHuR8J9NjkIbdGRvpPO1Q+0BC7TZB1Y
C1YWU1pRKnWTIUcQA9bMAeHrof6pm7oWE12DVafqLeE//NpEF9rFyzCOy7DPkEcC
j6OeiE1j+QlDlbsX4oIIdxmQ3hxGq+KLM2aQu9TrWJDBPtF1TSijTFL0kfhRN/Pb
G4hMgOZN9xUm+1Lpl6eFVGVoQC4K/cbGqF0rSx8QaUp3FNPB31/oqme5JkA7OfCq
8uFu2VNCbKUnqP5nDAR7KV5dWunk+F1aozcxJEVoYJkh6prfY1DTEIJ5wOBtnsZc
zvc/LjNOj+3Zxj4C1vHpE+53C5FIpqcsiEqHkBUMW7OoK2bbdgyRXYzpvOUF+FUU
BtrTsOp6+gZdfjrn0Y9uis9TpQSByhFhwn6m1J1/X6g0OFG5JJBoIuzAECteDBL4
PiqvoVzSZqijbFzdmSJyndVZVqVjab/gWPUFCgCbFVjN8IrH31hjYl+zX9Ef/EmK
dn0OqVwOewwegIEE/ds1ZdVgObaRoY0J9zcol5/xjClHEucwQW7VRd/zvRYHX8eu
wa2mD7p/Xx9dEzzcINg9wtjV2q87PD2O3iLd+21UJx2xK1gdh/03rGLCX49k9kVs
0EUiSHxMMhD5FRsyoarw6hb/JX/itsbAx2xtkmQXucFd9YfxHa/9tld2CFTpyV/a
sX58OZjJSpbkbLpEMrmOikWDoi8eGwLesNuNLu4MdNlPeRAgMjyeLXX6yqsBL3ym
CI79Jqd/x3YnMvHrJgA4BtsQg08b0J1MdtX4wN6vK0GH/WH5usUgRrroeAmkchJC
f3vlYYKWV3Xlgc8FkNPfd5/+JRmff3qrsybERgzJ+MPhflghk6US4gVfXK8m8/nc
aGErvxSrGWFiuYtIhVlxtohZ75SBXtZdvIg3oNA75e66nk5ekDHyHkBy8RYDY34+
HLK7tGpEhdzfSRmgKAq+9NfntlvgxsfQgcTOuH9St+fjPdfJ1V/J7E3H0Cj9ZP/9
ObJ7zHdV2HrRIR1GenHZmDKtnBS2MmBNZewOPxq7mdAV3zWVcJq5zh3ciRTpoA3D
1NgMQt5VuH7ZnjK8mIrOOaODoXZioACXhVLWoZTe6Eerq/jdXVQ0H6s1Ypj+e7vu
BbHPnl09WOYCBw/4Bb6feCggcbYEgGGW7C5CwxEXuRUj/a/f9UKy3oKHIBax2fKW
ivCzq8zdE0RcPuOOaxvkunP6OQp1pAHsOnlCgr8lZksNScMW5Nl+Vje9ML7os52v
Pyb7tKkaFEL4z89xDlOz36regAVd5fWiKacXXYTEGCc5/mgw09XcHvixZ5aGgvzQ
5lLWZ6RHDmTWuzhnpZIZ37YkibmC+B/TlCF2wprNIJeEd1ZzgYSJKKXOSSBOCZLT
q2vdAwjCX8uRcoTq6zV01tiIJyT9E7hTQsibVjA4DeryHXAy8v89o3Nh/ybLzWOO
5sLtN1Xx53H1ZMjwfiOb30ccGaK7SmzxaLnaCGz/l8qQh/Lr7gp2k2oHzeWrgsJK
lLV0biaQjCC5iF53rqY0QCheLBOkSWCCR3wUWBR6BHEYNS/cXlaxME2BwCnE2z40
HKDiyKZ8LACZicJYV6fSlcmpOhnxjTmVjHOxZxfViSjn2s5K65o0qNFhFwbg51Cb
ypDwUGj89B05J+ZqUOjK+h/UsiGIkvy2D7WexMKNexjVHu+jNJaGyhX+PI7f0KfX
3VmzSvo3yi/4czmbCu6Omjl+bXI7+5CbtRlSTy789uhMpJN5GzFhVk/icNYkyDdI
//Iw3HfsAGnHPLJvSTyXbjbU0D8HMG6g7TgHE6GRE/gJ8A2v4Eumz0K/o7spgRY2
MetPIldv2ytHA6jswqE6gK+5EfitEimOfTcTI0z9+98WLIXWe7JcqfnnUleSv7uO
+N9PnE7KDScDR5gcVX02zAKhw7plAjs1TF4b+W7xHbA4XVp4ySewlKYrMgX5GmyU
PxDJo/xnK1hVXipfPg4OzOwv4lWlsS9AEZb0SqmmOq9K3RBh6S8zDr6JwRPWXyxT
7ckxvZq9Q+Nib9JfX9fyZsG4Llf6Quv87KpYO1F759DCkIutnNk/BkLSa+DDeFxD
6XAl9AhSV7DFVpYXmcT5zdUEcxVyY0TjGWXflsNI2pmnX6CiPIZPosZpQk2iwFoD
fIUciZQJ1YNiHq+h00NEMuogY0yA0comDqLmvlgFhfO3e4tQB2DWxM/AN2Ygdumi
I6BQ4Jv3ZyYd40U5RcnhG4fYzWUQHT5dsKpGZvZByKaR2s2EK0YAWt6gS5KsT0DQ
1R3lmW2WLyuG8s3UYNQoXKHeS9nOGXJ/qmmNiP3KC4C42IOAaGLmur+sEiVbR8tj
LjADGEuJ15LnoyD8dqcSj6W2/J5hPCqBR0lV5qNmVqogRP2ta8ZTHkuCeXnyZgkH
ytfCvpvhrQs2Lz8ktxN2tOOxAkn/YJLbgXIPG95054nzXlyI42Vf7PmLHu9uXKpJ
oOD6r3Tkls8iYmNYDEVugFihUHan4qq8WLo8/k6ii8CJdSc//sJSwl15+ahahS6z
2vPQwaibybp5WN4+KW59NdgNB9X34joO4hGGnSyiKpoguQ/ks5uU8wC8Sll+HgVr
jgMz0K2uFifAFGOICMyo5Z7VdJvxl7sDO/+UizwhuAEbsAr3cwud+SD0QsyPPfGm
QAqR5pJQluJ9t8kwDgGld/hoNNxPOVyn+7LaLMohdt+mOmOEi6qvTCr63KxwKYH0
wmCycbKzMjBu1+fn10EymGn2UXtE9OqP21/fonhvaCDOtw5LOjkdMKY2Hwf+zkOx
AMTXI7pMxOhzaCzH7KYwmJgTwoTvD824sag05OmgdJLGIRua4Ifyg4TSfr9/P7gp
xFXDLx4S9xvcmKe9n3KyDpiRHL4+wqiIRiTL33PR887r9C9NVZI9cO4DWdYqVoqj
J+nnvfLKpheDOyBewnq+KWoq4i/gPSmQIj2fQkD2MolIy4ZV5SAsXr682/0lTvGT
udzmxcWupES9poayOxSKungLY8iLSKPJgtpQdVct5XEOoe00BKclvMly58rcdRE0
uqvznMrJ2/TObFJHhTpVDQdJXmiX6HMgmvzMc/G89+n2Sk7kqzE5th+/OP5XiaLf
uD2YajHosYX9xBGG0n9q/EWeTuwImDl8cZGMqhlo+yDR+tmSgxr9Bv67DeDGDxi7
oxUGx1b0Ks1DyjfXIIc3qXRep6yF0/Wn0RVlywf6lz1CgGhbzkmX6xcE0FzKLujj
dv2eO/MEYd3joxh8hTMHY9sWa0S5atC1wPkX/yhflMt0CjbEqSAkSEojkQewHJyf
tDRieR5x/49x824uLYp1heImKrwNsXf9YMPwLbszC89JHBxtjZY6/71T0pqlX1zW
u4bTX3z+Qcq5HdBdykzQLngQfTiBiRFkt4Gzn/xHPoDw60FU+/reLnvMGUIp8hix
6MpPkoTL7QUSoc56nT2oI98pFAf0/j70S9q+jXEJhSyb2UgmAuF3kgiXPP3MIkzL
9fwlsaEh7xj3OBXCc+02w3AuaEkbrzf3HXxXdrKJZSkkHs5yBOYnRhzuZbMO0dIj
C53jRUMOTfcC92LIvi0h4Yn1EICbcIY14S7wShsgA2yNagXx66GENJe8ZKscGPue
OSX8i0OAUyG5bXY+kS7QVwo5stRnDBU4eaSwfcR4B+Y/d67tBcrKWwiLCv2dibxk
vk5mn+dPQkixt7CyoXh+qfP7eYb/ruZDoj0eGLomhM1FQoJdTCktY9bUt7a7VC5c
EFyPL4nICRqMw3JCnV2IanzIYAYzrIYGyWAki/RZtCnqowIS4ZF0Ysq+QEBB17mb
7hzqHbv5+ghzMBckXu2ke6QFdmcP4VFKlm2K45rcKEZD76dVMxv5WG7Iq9JMxeq2
lDKM7luKUQ4ENdN1BKwMIzXsdHQ/1HJj2OEPB5B0RP/rmEnIPwZdjCME+TWCUxQk
KZewparrSTb5GxWKDx7bB1sI56TrZ4yd+pnM8HVt1CzeXZq+R1KoA2AUTqA4OlqN
PBWG25ktdMRQOYPqj6HE2aSQ+9lopsXJroWk43zSnxQMqucdsw+b24yfzsYUNuBq
0jQWvg+iuntVGa8j4n10YN/j5nKB17FXfzG5MT5InX5bLaIDCRz8TXPVP9NiOf4B
x/Ihtpf3lN+R5SAwcnMU5E+FDM5EnlFBMbeR6mVxh3KFeCp5Ti+pOk0jSA23yMkO
PAN4M9+0Mf0PDjMI1W43QrQYcyJGEr2VA9XG4XRefwCbzuKKlwY3TeREqLgt3Qb9
kKAo3089KRvybtp4IfnV/JT8LvniZeJ2B1aez2IgmZ8GtA06l4KZ/u0xWPDE1VYw
1bnGtIYvCUMguYHp4h4JYQNjoDF5+Vhn822dPdVa6nKzgrv41anB4At7G7wMNAcl
9keOn8uSsokV5lAhrxhUl6hQckwQeDOWh+GwyDh6d7/Bn5bDubO3DGALegAdy1vY
jZYfq0uAE91MIh4wZhNH17C/qE+XDaTSV6hCqNCaQtgWU1/vDbWv3/V29VmJdlDm
Vi4Xj7HwrheTs9GL3CjLQsYTKluWiS10Bnv6sEH4OMn62oao97e+vdFtoMJkS6n8
lJGsKHgSptHjWI5LX000PwcuKhvd+qll4/F0PituMKO4igyIfxYIfTFf5NYUc8V4
WXuN3soetxXjah8NJeRcMLXFajFG2bF5V6jaUpO/L0c7UD7JhsIlaPDXeJ7oDDHY
kaRA0FwcYJ2L6TBleg0YGUmvnwhNaT/0njBr3+aDX/Grej7xffT/veNNb2slLSjm
akbtK/+wF7wTtz8W7VZfREgqnnAScFVhGQPluMqpkzFFsK5hg/GLI7xsQE+zxXdN
n18TP4DYoy00n2kJTNaQ/Rgm8c5J4xGiZ98X/R3LuNlUjOkrik41C+s/Hmt+uMfL
dFIUcrIRYZmo70roVmQW1VmBob+ksRFKd5q2YgNUMEQT371RSPr3ckqX0rQa0jZG
cL3NJKjAuFWhgPGTa7SzWLQ4Qqkk0/FvKskYCjShh4M8oAtxk4WRkarhBPk2eLfJ
HChHsbCduU1Ysdlg7k32DTjcmwvR4INsAhSOniuHQc9yTmXRQnjyD1AEhQDDnxz1
9m5bIqm0lIqIS0Emh5RWUb3kb7gRzv6CnE3NcpPFT3Hs4/r99ySiO0XpoWXcXFOj
ZtyEIHptlHqFvrxHgosQAB0KOsF0saAWOuk/5Hv/IuTaYaU5+ps2p587tT0KUf4d
vo8oXyIvZ+HZk+EcDJDyoHd+s0gwcJzZqXK9lCC+QK1S9SEiLs1oDv4yDAp5+qJX
4GyGqUww6ITQN5ti4TS7dWH5WXKpWhKRbAZRdrBga1hs6dCOsD2cHu4jexiQSFB6
TZ3g9qLxa3tkteM6FQeSLx772UZ28LMEB+oM3+aRF04t+sYRoG6Cap58mN2ckexJ
/UROQ7WmwCK8eyZOPpQNvqpsCfDFaeDAo0T8/UlcJ3MFpo7cTcLTSgE7Cct9of8g
+GmxY0YZZ7fGYhWUuJr5YNdRcHwOc4xbt6ZDHZ7TPn+uNkqSg8BluNv9mQz3EFAF
oI8hd5ZlVMPL4KpVaTf9IT/EAQ2SzFl8XbN+tiIj9/jBIAPmm3T2t9Ceas6BxEUj
oO1I7xuvAkvh/Z1+OUamBue+B+ruo3FTbDFzmICoJDJUb8r/WaX5oSsJDMO7b9Q2
WTBppNF2SaExr5xL3O2to6EB6iurpMv6sWOnOE69XkfoD0K2tUP237I/4mf/BrX0
jHOnrcexeH6531w2hIgr3Vti3aaq2/vvzwTnvwHZQyH2QtIzNKEbTtABO4rDz0EI
0FE4OUpxFObKQskJjwdZga4CzJ3Wg02294vBw4GREb0l93ueMzTlP6Oh/kwLZ2YN
Mxr9noeQbdBi6NkP9ayaSj01KgItP1tWzFbfj7+alhMorA2NrNmX+OGPzGBuLClO
4kTY4qGaodb9i/CzOSKYM7AEDmjIU/jGLbg53ybp3KBWb7xUQVvAMv5u1JP4pTft
ouD8GSLiB+cCrwgsr23blnz/m1YtF3f6aX1FfpNPATR2WHP/DaPkCD/o2qCwXLjr
n0IOousg7ETXti7174t17Cbn8Zqpnt2OEfq9ZHkMdQcpufEnJkWQxm3bxeQeM6GZ
8BeZ/nzIW7LZhWUr0gH/ftwj0wyGBXk7M5qU7YPuriXElPm9ZXR/QoohvYCEEyeD
fZadWhWJPw0AgPTP9b/+7Ya/XlxPVTZ7ZFkb4+6+sj5GQwGZjen4g5j0sOENC8si
4xnvVYEOUBIosHQAVMFCfCQ6cqRN9qpHP/1fRUFWqhtZFDQ1wYeWKZVDlfNqHRaq
g3E+irHSt2sHKxaQMrWkl8WbyeQh9yKvQ0rS9wpQaMyBXhoEDaCoaTei+Ij+CeLC
VG36LkH309pEMpNqF4eaf8zuNB+smBvAyy1z75Ojjw6ICNRZ1BzHiDVMtA2Ix79K
b8xL8CuetG28uNRE2jujaVejp5qdl3Us9SvvQuR+TH1D4r7IKqMMVVotCBEnCND3
7amjS5D2vBkBbgUDlo3Tj3AaaEf1nI1wIv29RvQMyh87ozImJ79r1Gfsg0HDUeDm
WzJedTTxPwJVF7ZDfOa7/yPERKCpdpqCk4LDE3dsCoNO84ekl8A+go8LcJ4HJ/Hq
vHzaA3j3DIV6yLsoNomNrEgFM+r//u2oFAY7MBvHJO+uctHnxsV+xB7CZTP94JsA
mbgzToMdI1QyWBBL41LBZLwtlFlbeuOXYtt8CPybd9Q0yA7G9Xfr0lkSJU+rT3bf
3cg9QkmyURGcgvsIK5OcgiJKT3bsvMHL14WZ54WF/w5fZiBtK7Mjnq42QLEu2Cnq
pyivjFOOjrl8shFTpghq1kaYWsf5fMuJkCSLPo4IJfEvm3sF/yGyip9j6MOW4I57
e+e6EJkhFpo7QbiU8gTdMwVKeKH9VO+PWp9ChB/zlu+9Jk2/st3gR5vTzh4N2PVp
V45CYufblhqjVmI3F5iec80+FcBeDzT8aLRBNCwrsGUiLnNWrjhXTu5FgXBE6GGi
9uoElV7UwJWXZ3SmVVxeW5RkKPMYYb54JtUy6t2rQvnkzluAx1PTRPki3DOwg6Zf
jBafGioMMIR7wWq5RKV8CkJJwqHQxyuzh1xHpqXXiXs4ZT/q/p8cyES9ipsOTM4A
vBMtsBiaZy6vWQxLUq+KoORMtqzHqt+LkxdUadOD+fy6VTK5Yg/f/ghsk5KoU4ZJ
lckRuPelHsQwdgwSSgZFI4GhKkeRsfO97xDz3u/ZBIO4VtHM4mfSsHBXUjDLIOpL
9FcxxMSeZtYmD+kswdQWQW7Ml+E4xMxzWsnSS6qzborkqd9YS826Y5LrnXj2C/CO
hsIyPGoi9l2NKr09NDvK45fiMbwUctls1Jd1tvbTTLtYMHYPxdkRLaVVTDjx4rAZ
s8YTAPb426RGZZ1/4h8C3E8iMoZF8k007talvrQBzGcaCiLxRIS/vWsKPMhSvZdk
Ru+Cow6gy93e5gE2PbK1KEVXO/kUTNIiX78ZRZfKflA0TfdsDHbqtQpC/OsU5GpP
RxymOfVwaI9mlS4KRf5+tJf4OsOzdbMwL+pK45RIW1GcOSeHOqi+U7YHN0DU0mnn
wZCWO7kMY0ldEfqxAC9mKMG2iAUDKDz3zvDVGQdS1pYq6z556Y8TAXe+BZRwCGbz
JKuFAQ2nfhyjjgmrklamDCdwbJ0xjXO9ojjC3k78fJJ9Ow1GOq13kzxtu5qPjgdU
2lxOiNUde7fk7kJjYKW/QUR9n+M7MOwH/BHqZ2zBtxb3ItsME1kLoDypIe0guGSa
HB4n8Pk+B0QBPdHp7W+yCJh9O9pOz2CQ8DgC44Mp2KP16/x5R6nL/FxVm/5Rn7xx
wYIyycBXSMIRtmXrY3oWzlx+gSFiqx8A2RJ2T20hnvAqTp6txkqjXhierprYrNbs
ffZ2kFVfVXlOLt/j/7f4SAMY4OfxQ6wnqrxT7NIPrNww1PO6exP3PxN4H/DQ66DJ
0NaijfBhx/k5HnNe5bdIvZL4aU5mIuw00MKP54J/AgdyosnstiI1NoJaHSVcEodt
KbdsQEcyNo+Y5z8CXVm1pIrpq3Xn4rQJVUeqAllR1LcAgc2Vf9zg1Z8UUHJrLKH/
PtbKTRfVmVcSE9GZuNmEVsuxRX26l0N2VjEw0B/qVjnxpgEM/LBQJja8TrSLS3WD
7MI9J3mF17PJXGjT+n1fa6uGjodoNu8knFJS26r7Da0HIzzuEiamn63wHSYk8t1J
K4nSTidSnVU/vDbez+17Dv4wIgWZFC9jn8XoI/1hbyybMe2pVwrdzjx38b1a/1cd
kkNvgw2G1sqY+Xnu4nPy3/cosOJNnku4BTjS9eRlHf8oy6X/zeRoXWfVXVz25Hpi
wd7IaTSBaipz6BgdJaRjnNG5syEbsiqJK/845yFBAPYTW0JREPwu2F/yDtJnNovc
bFqs5+0tGvnyAcBQOJntt/v+iRdzaeMXFC8bjuuOH8izmGAaXHhz9irYFSSqHKuW
FgnVntkwGTvrnB7oGtBbB+85QoGMK0YdBgbgRi5rQW5U9c2Eb3SLaVuKwqOGIpDD
8rG6GZ9Hm9sz2ovlOzWzgQ0bSfo4uomuj/heJ2N+VmC8aybpo7BnIKE36YzE5+zG
OllG4FfNUFF++fFqaXlpLoIcBNwDW0kCYQ4xStdWPl5X4JvY4Bu47gx/T02LLbIG
YRr2sIabGyn3CVGXtOvMnAzotQ61Z+1VGge48hpHC4RfRkIdR8WwF3zM+omaN1Ie
hI3Kex+69OINPNeUGm+050rWSqRoqmNDgBFlJvkgDWYd8wDo7FuqvkYppiSChOCs
A+E+dn0WHPyIUdzhZX8jgvTgYBeuxEKYtwFmY/jwgBZRXN07XXoVgUKlCKO4Oj4e
zLkWUF1VFTQjKtoYXP74U82WBj5DC7DOVkvQ5IR3PMhFvBsplYql7vh2hIq0vIx3
mG0sPyYBBtrHijBAuNnI0xdmy82/urpHkRQOXut7gz0xsqcADfXpwnHQSlgAzxD8
lZNlEaw3NyRirrklsz/IFBo53hfCbwXFlAteL4UUkeVrNFfdab5bRUdEgs3xwLyM
iGc53WJjwPE11Fhk+vlgz0c93LLXE40OA5IH+4VLB841E7NsxKfF/CclYg19g1Q9
1aAXskq1pbJdO3+bIh/8OpA3X/7UIco2h/e8zZCQtOk6G8XDBfNm4AqI/owzkZib
Ai83OO1U3Ewx2ZvVfElap79lnWJIZP+TCgvEq7lNoz3jr3r7S1ZkDlGqvEZ6LGaw
Wq/q6dFvd1/bYcV4I350QKct4Jy2J9/aj3+zF+RoZZTeASvWX/vJ9uvTGxW3E4ly
QKqrFGVa/Nr0W0/ewgvCyVSJlO4yxMZxf28cEQ51sHBNNivygmhTzTP+PmD7CeM7
hnHsrtaxq8Ez0rMnoYSRhVp3izTUS6AHiysOSOxMU4g+mCuuq3CqhsjbRziLxTpZ
0+dimRz8KprZf48M5h0thdzk0GYj7t4USriiyuoE/Fqe9QeOrGNpjXWxvrK2R3ES
rKP83l74jhFSjOgRn1JD/NnYt/+c1v2AcgkTBQGlP4WWMHBBHSdpz/EBvy09LDfC
6MQuX2DxrWjJP1bb3ZIl1g43sicTQwo8K0c6aagbysYGP6GPPKV3gUWij6JWgrls
XGXqUVi18LlsU5Fx23hl5AojWnkwMtxyo1rf+GpP5SMW+sgUS3gXFqWC5EJ+ci6l
Mj5WqEnvXR8NiLbxfNNS7hg2mFn4kmLhLaq+gm+8oPPNQRgBFZLnxo5vO3LlZViK
U9Sx6SmbrH4a5EY7qG1BPT8nnYllINhZkAO62vbNuel6fc/0Fx5Bvrp+vNGualRL
mupn1TlbsR00a3p70O0Py7atfC+FOBsq/L6JB8byABLPmtxlxpR4vS0JGLvgFBVq
Oo/2Mhm44AvKhh1MXfS7V1lg5T3IjxrRqpD9P4mIAY+5tJX6/IWlpM3NkOd6M95I
7QrfVtQpRdpAKF+o4zqoR2mwc1C8n5jsSPA3QhY/UMDQ+kGuTDfJUp7S6e4ThxmD
tqvwt8vRZZhNDqDAk1cXOBSx6Kh+P+I3T9s4TUwKA5j5PiJj/uBnrvvxYwdZq5xt
oVcQv2T0/VIDRDJsSihNX6heZY+2N2WVtUKuAoNMBL0Ap6XRbjVcxJPitRIRDWhn
q1hNs5pg8ERrhjY3qWERYxIuGhf8PuZydY1zHdcgm0NyUWuv0Feo98ZCIzBIHJ/X
zrAQaohSya8wrBooweQoH3xJVmc3XQVeOPg4JTziz8ujYqQKbfDzMdWFy5E2bRbc
xmNmJiahGG4qRneudlcOR5MphDaYM5sJVWuPuhr9V+ZI0IFRFNl1DWRiBN05ypJr
BjgzfSTVhqiAFZwoMctPqFFgM49KeuZdGV37JMY3JYuHoMLIDzxPx6RWze+oHWIN
2oPqG7I4qUbuyLS+uoqR4w8Gr0ExKEhLFpfx58UvhPWij+/pFrPvFY7iOp6F/AyC
RBhHcLxvUBSuhhtA6Cx7gRaBFpdB7z+EYuafIHpg8OHgiDbpEAf4wgA5j/Jn9ndh
w9cFv5CHJNJktbZmlpe+lUTBVcp7nUNxE6/1rEsqri7Fx4JPR7/4mAJcjlEYbELZ
Fup0uvMMA3h2tANojfUXJzzELZR8GngRi9RamUDHppwloT74BPfpeC2rj4PaAGIC
Hb2kPBv2BgqVzJuU0S8VDLBkq10dfFasyL49c4N79i8cL5wzuv6VIwHeIadaeqtT
Y3goANgw/G8zcHx8acZ0rB912M3GbjOR8yRvE/OAP5CxJRvxkwEdTkPVmGbuKOLN
+lMw+ND97xXI/TsnWargR+B5llVvM8ghy02IP7EhnpCP5lCqjkjpWOiXu/ds6Da1
5txSEMx7pTZqfcCxkWJ7nzXrS0ZIDQCN8u63F2lFFQh8VGGKEYycvW6rb/Zant2S
1O2suYMi+uXlwB5pcKlnEf0fFDJmg7O8LRzMqLgm39jndNsvlVJ6nHmPQYU68C8p
Bu7nzrPuuUQh8NuCYIH8ifBG0Gck/NF0zodgWYiw2tuuQDaHo+cMQaKxUI3yDoc2
1xSFfFTzJMChL5ijrl1RHWXtxb3ln+yFvv7cv9NAwdZ5+mRnev2M7xCwfPvpUBvO
YhFSntrzOO40+VJleSqbeTrD1V3xhWsVTyV87aShqTkIHqEOmH+kRF0iYyHJg3DE
Nt2SU1Yo0VpL18LXxqyDw0MmZzJkzeUfciiydfRhgz5+5BwwuGmsUbXMhxGquq9O
7AfihNqL0d6+Hco2sFKjRJK/FGnyChGWh6vzKNuQFbLGGTtG+qnr/VfOrWMlM9z/
0X5C8EZdwt8ARgc5FGA43/atGrPWkFTR3pC+K1WMaLMglcBDrKNG/Bev/UsvFsiX
k74zF3xgO+q2wZmKDtTx4ZE2hSRX8k8Dz4Leoo84Bf+dpJ4ZmmPf3LnsiUxOuH1z
4o7r0x1QYTtGdSIzGl+x96r3jOFLeQLgEM0Z0Jrb4M8MWV+Ybr2f02VawfBiADYy
lwWO5kBlJHStH9960ifeqTCPwmRt/+oH4OZXUKNJnDYq16q/g9X/1IWy8skRxm/y
nt0U6cCOI+j3uP8BhfH67IXGO/x9cq2jSUgTlx4Zz/RpGuuryiLBPbYGj6+H00WH
UUvkHAB4KgI/H6qH0psuwfIycJ2wmPNkbavd2/eqrx8gJdsXL8nBj8hQNQ9Oowfz
sm+pGvQV3rKBtkbmNCKQUEcrCJ8CSnGT0uJM+6zMFDLapPRn7cjR7xoJmrBpE0tL
reAyMS2BUWzv61SnnLqQEnldkFxq/DkcmoY9wYtr/ezn3orP0wWz4hc5ar/Dd1RL
eqNsjlq+TbbEW1Vc4nsFLjY1YId/UyoAeblOZLHsgCE76vbWdRlgOZOWtP5soAVJ
mVIMDxOnbgYqyKcun+we/or8r/9Dw9Kn5GYG6HYm8TO2kcagWGx8xBCZOQD1tizn
tJpqRmIejEQT1c4qTd1SJ5j7ppP4bnudoP1VlFPkaUcq1+CJ+G/ywc25xmr7T3x1
rIYEB9uyf0NAMESCn8xZmexQiN4AZIwnbv5eNZVzv6bijzzrZ6OiuflDhsOH7P01
Dfd+AHRNZXvKii424BZYS5jE15usoFMCpXzCF3hYrvd5SCaYx2wXM/ikcfFX3+iE
havLtDKdmmwhUGRLoKIbRJOtd2yhjDyF3jrZfizzg6i8NoNIJEIXEMew+gtr8mkf
9jEShDoVmVAPYMX8bWaRzQT+NFRzl+kt8vDq3pS814yd/Yei4usOvSVqk2JuYVny
k1YPuiTCycWbEu+nX3o0H/yuXWMLvSy3DPAb8zXcaHUnC+wEM5LJZSkyQoxoNvc4
pEjoQprgPjchRSUpTgZRk5HD6gUG3niYvN9ekQAaUhqKhO6l5aVl2ZPW51Nr1RkP
S3bkXx2Wfe7CT1TPnAodbxONOuglZbkRJuulh1UbBf4tePZ+1C7DzI1i5LLwFMrh
j42+gsk5VCzfbT7l051otkfJsMM5lgJkz8l5M5YAi4JssE6YAdBVp7ahI+BeoAwb
4YbHcwJ9trzMbyHz8hi4sQUVRdJ+MryXq4tkFZneo8tmACldR9gRxlVesvGoQYIw
fptQkEAnqTrGHbwIt0JRPG+Kkt/sDqL02PqCvcxwNVGCGsjJu2O8H6UndxKGe+aN
1KKp1hRrFC8EGWbAl4VQf9TdCMv7iSxIDCAyekqUGzuWqMvbyobYpJzG962eVPP1
y7G4sbRhytMZpoqV5D3rBBpVygiGgUloua9i+0dCsJ+iHwS9+QBo97rRgENVs5S6
VaVP6yQJWi22Uy7yYuwuXELsdcZakzVntaq2a6QEMR3i2kFHqoZ73gAdNUCWEIG4
GgZIs+UBBom3qc0dMkax4MDPd0eBQNSzMKbOLcPLponpVcWMPHgcVzGV1sV6qBep
fjn7Vy5RCgsGZeo9JM4KOhuyXEIyQ4skJapSfUV/6LNTwm2sv+ezKeokhNA46Ekf
DHLAJVLlRGBsFg+XxLo//hiFKkn6f7h7aJe0kYmUnR4rRPAjUHTHlBockVcoPNfm
qRKn9ErtlwdasxUgYm8AmqVOohW9M9mD66DiIBI1e7QE4CTsnF5T9laPzS/Ws7xA
g/i9rt67FU52tu7w1grgUChOLKZbaV5PisCZMkgV7Ru45rvItmbNEUef9ZnzB8ht
C8VIPK1VaSpf59ykRMO4MNXph5XJjOz0x83DixkRtUyQJKkH7jyO+lU1iD9kSOYh
OhGLBR85LCApaNSXFYShczg4bcsgVsIPUyAtTRys1zUwuG9g2ELg/WAuUOqpkiMK
bHbNh+Yw8EkJrMwlUqiffKwLA+UwIRcOLZ+9OTklNTBMrnhPhMdMki120J+1jIeW
HMabg2j/JMSsFhwee8ePfmYn9KhEuHEfg9WLfDgOf0KPXyRjUpcn7NbUbWecIFf0
uq4u+VPIMWmI1GEY+bPGcy26kdrlBopGGs44fHPsS4jtwXp7ePS0bGmires6ynXa
b7e9M8zTUkkLclpYeHxShM4oZdxgfsIyDlbatI0K+vYUbRrUtNXkiyZ1VF430QSd
tnyV99nz8Ksw1uDMs9c6JwCWLXrEEzeZqGprEgjVGR03GNProo35uVi6NnMB0TUR
TNpbcEg2A3ee6LFJUJmRDTXjA8289mP3HAoKQR5VcW7ZkNStri4mVzgGBqiFfRrR
vckC3Ky5bCqOAsyRMjYaEUJDnMUVMkVGU5Rqg7Cg5tP5bGxrOTsjI6WUqxDV4EDH
XYu1p/uJ2ykJpxZehh2j9xNknhoBVZN64lqXdRHJuQ+lFPS67VShDH85TfD1gXnQ
75/tA35jpnz1B1RFJS6hIkSiDXTl0NGmBSnbQliJX/ZOTrxIDgnVFX3/G2hBL4Sk
3l1m6uTrgCASkmkKPYi1a6IS54VkO28ZSPgxPujUVrPFOfz53AjfM774I7sCMjqE
l+VfxhLjVNGJhIW8vghfcXf9E5F34uLwLOi26cBroGnVuu/zGDgSmPElY21np7f4
EglqIPVSLdY0DbvjUZyhhhuxjfrOOLwqdTBTiQNL2LVGImhbzSoVvrv2XAyNKzW4
8EN9cW3puCa1G3OxVKsx270ak+D/jBpwMR5vVBh0YoDnohRJrokUt9s289Xabtkb
tRnuUK5FvnpNRBjTPSscVwDncqKzl51LRQXpX1DwzBhi8uBmQ+8Sgma3qEiJ/gYe
rZsgO58nSblQFl/HFa9+RpTnen9kDtDW2XM0WEH1OYGyMjpOVlhJP7mRhBmpcMlM
/tXriZmOqrviYV3nfCWfP2gnbNYYqXS9i3R4ZapMDYuJhgmK8sTluI+Wbk58eWAv
MyX9rWQ7jTba4z+dNAZVSbYN1DVjSkdRg9hH2hFVNYQ5umo70XGhFxtjeA7d9qzN
VZeM+tgG6hkkK1IDqRPghbWzvgOyps+njM94qju3w98XDmL80Fa+60Ah6cXw/gOp
loh86QRERR4zVdH3r7EXtiH5yGXbSOrbnggFCMUTWaddXHFyQ5MRHcd9jWeAgSO+
NesQob8yHdlErIfT7LHx5F+PXhS/jLc7cAecBUYUNXoXJxlVWiJ6oM00IUaM9qSV
/zFQq+n80oX6Z4VtN4l50wnHLUTOy2iJELclcchNvQ+IphDh6/r/cIM26slDI+mL
rOieiJV37Mr4FArmseDEVGvls/a0DuQ7XzzQBF00BP90LIOD9Sb05OoCKGTcis7J
DYY+ZTanpQBzcZEl5DnBn+RHM3nqvAa8W7apc/gvoE6xclwe19lM7va5wXSOKybL
LXdrtMghCQ0J1KLFJaX9WGmrCRNTTJxsdIyjtwAp7g+ORSyxQIhyeIz0UgckFiS6
2ChHBwWFEhtMDBk6DWLCEcdb2csJjhBXhDnVrJImzeMGbC3trmzL33i76akrkEs4
RgusOOGpZKScKCrA8t2GJPfVRcK9DEjtk6I9HyVII7//iW+oA5Hab0aeoMg1vEM/
ZfzgDesDvKg+GGCqQRjvw9/u5kt9h2kpjlhkBz5uMpDg69vh9bGr1PWOY2L7Ek9R
JIBlVUSGtFC+A4WUGLaE6CAhy1vYNtICnXvT9rS9NlCAPIaoBvHIasHGWEvg8zMC
w3EG1egEQpL9VQQnSZVAn0rIydZ7TnkHsMycMdtZEeSKXIDgEIX6yGB8eRkGzDMM
iRLEe2Ftl2lupPcOb9IlI4NLq/oITdaaunEZVNLozlbw03ASLqv18u8cgKFYRbNS
X4LBWs7yycxHr4T9SdLkNVWhbClhhRK7tFYQlxRyCTCrK/9af55uat98rR8QKoCa
F6Zw/rUSmqDgna6UEktFTYZWV6OLM0Uz9FzX04bRnb/rqZr9n9WGK6hW1bHaqhLt
UVkEztOGe5JcURL3nvoE+44s5V4BfWWcGVo0EKKr52ouvDI7vX2D6mekzJjTwpGF
02aE+6tAoQ0sK4k60EvD2UzZi8sb95y6HmP8YHhOy/HQ9UIoy+Fu7yYcbOQWTkfU
OWR0JOltx75tvjiM4ak3CjveyebNuXMyVyCRn7rQt9EBl5QWYxhmIaSvfdt/ol92
zPrO54IiJYDOOeh5WokZqEg+30tyiqXa3clEGT1ZcMFf6j7sYu6tXE/0Rrv1Ya/O
wEJ2iNEXBVFw9kMqt63V/AhJoqfQoy5YeKPv5n3EdWM=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ZuOYYHRjJ1LPpLOrzPoQfol2zC2yVEekbylgJ0MBUOEnm6dvZTGuSV6/I0ryIMXV
CTj/axbzCwtXVNbab/lx+KIoUsI9J9jIzNbhFILHJ0G4wXo2SctOq143040PvhuP
raQ1T6cb+kvcm3oJ6/N1XNuYs5FBscPLfsNR5UP+VjM9BskU1Feti74SPbLtAEWz
yDMQQRD5yxt6yA6Ez7apL7HJmHh41e9g0ynsw69iJtdBYUgkVVZNXYHgKWrKA/9g
xoDWndzgTnB3FGYJfTGEXULgZGsLtIgkTlaI8Nejl+eaW0SrH7j7M9cdcKUGo23W
vi5p5TfQ4mTD3++tf3VPSQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1200 )
`pragma protect data_block
IidXndJO5FXzvzw+YkAbrrDoORI4JNZspD7d3G7zmhl6Gb3ZY+g5SFbX1ksp+ia1
TLcwxoGPBnmW7gPHxoBhR73zMv+MW6V3d1reUnm9r4vrOKDwvfAYMBoWQ5XaWrmU
mKUnw70YxFK1MmdYp9tfL0BAI+3bz+luf/HIe6pUoaaejtyuEIrYXPaypz+Tm62k
sYkV27KB2UBfJKHvVjrIszUEzPEG6oxJunF6xVNtXp7/YOLGu7RpWFmj4iXM0xQe
tLb03rn+NlqBQ/y5BcyRMwHldWbLAeZ0tokzPpBbPVYCmBtupABUO6iwXUuTz9M/
+NSS0LGtiRkwQ7FsOzHurdyRnH6f8yN97fI2lmQ1A8caUP04fWR0YMRWdhL0bX/x
rmrSGZnuWjQAg2XcWiwFqdSRMOhmvL2RPX17RaRWXM7VjZXtcD12mP6fBQHywxb/
ZoCRbic8i4VKHlyDfvKyC97JLNZu5v8pAYRg8ugnhjgA/bpjzZBVGz+HgsyMOacN
k4Zi31LcOuUs0GZrB+7Rxq0Xwj+kP1wzWM9/brsWJnXmIGuVgjjhHGOqr1kL3t9V
MXBrR8R9MKOB9Eb32euRFCJN8irCPintmrPfaMj+s83yWs7skv8PiIDZJKRIWs1E
/gjgWGN9sOKUPIJ0tqXIo082jGiV4CKkzHslpyLu0ong5IhZua+nV94ecwzpwuQv
HccvGcbYu6NZ6XoK3em+kHqoXwXChJjE1EbBcZOBjrv1rYqXoMsrXwkBhqmFdFqf
uyfPsC0QpTcWxztgT8crcSrPEVQOs+76llrMCuyMy8SvfGhKewY48/xRTPGwu+UI
VJOrSOWJ9NT03a9MX/FqjawcEjxhYFiP9VK9NKdRVC3fALaoKDENC3Bt7YlA97q2
N70no96KAjDu6y7Gyo67BmsOFaXqrpoGE6qL7bh+18fLkE2DCk0wDsFPIpOGXhNI
zhMsPzo0Q3Ye6QEzZzq6wYD6u1QqHm1Wq8KfQlTmDSmpbAk197bpEqxXxIMKHy6V
WJKBWIt9vjbMeLyJIhhdkN92wQi1/ZwGgYfd/+Mv3F7h838prJ761IfNj6AWAhjJ
naaJjC+IMnNKo2Z70/QuYvf1BHYRkPd4YXFDL9FBtG4mj0h0dDd9V5B2LdRb62KN
oXtNOX5TumxN585wHuj/ppluE59VyLX/zPcdX5Wac9KXLtxSYDHTzdnzFIRqDG2Y
XhmI2nL5sHpJTst4qC7UvPpvj3iZpf3xJcK4koGk/JP+UoSmKE44yWialC5SIRNL
NcNb/b1KZ6yTBF1Kl2xbm8Udp5YJmR1sScTJfqsiERhGqNJiiT1aHcZo7eSvnlbN
CoKDflAmPbdkGV9+GeF5EI3ok6/Ht6AaUdMAzRqIKdPHYmxA0C8DEV9+D9sJKANv
a4925jCN26iX8R2KhU6Hbt+EHb36EytW3mrRETy33uhTKHRd6G/j1wmNeM7rxYHm
TUWhAGCdUjj8zwtUBSkiNdvWkHqV9tNaM7n4Ne3yJutQQV/FIplldzyiPYG6UlPi
dqjSFnQ7+IXdaSsvEdsKIsX4LK3/5gvoeEaD4LO7sBr+rYVLJOs9vX7HUk8jlEDu
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lrpoZ5ApT21aSauuSckerHOijdnBV9gTVQ7WDN3kE17VhDjX+BwI7TtwtKq8Uusa
IxlZ5cJuscMPuVdDB+QzloHzR9RN2oXowd1ckSa5iwKmoOuZClvRm12KuOPPeBfe
y+AHd0w83Ct8H/+mG3IvqASaCkThhgjuBq23DM2ITvl322YV3W5nfAGiYhcjEG8U
KBwsnlpLmtIHdqvTg8LhKcRmpGSL6uZODxVitDfLxMFB1Usm10HEnbJuoMB9Y3QL
JhIl9Hb9AgwRcwq+P9s8NcUJsjU5WzkUZuZzwJGMj2Gl0fCpOubiEYEyWLoAssF9
eVLXxnumWUBb3Pe5KSdcUg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4672 )
`pragma protect data_block
yIsE5xXLYLhil79vCCgCVLrhlIg56WIrmg38cjrK5lGhIscIpiSrnUys6zDibAUR
sOOosPe7lZevd1u5L7y0tQMjh/nqBE53OOoZidDqY4qSLTpklyjDvXZxWoa6s3ue
+iX0xBld/4Awq66yWmvyCSrrIDsYEsFtittEGp3UPkGiloHPqYYJ3UwdAzd7BS31
jrwucMtEZCpBp8QWed+Qb0b2zwbrlCISWnAtzy3UZ3GvVSzG1XdRuRxpMgHcLxVw
rxNMFgalZuyJNfC94Yml5Pj/J15QVtKYToFqd6yIh+zXdbUuHLbDPKu6Q1gmllZg
fxWXDvKCGffV92VslAyAi6jouNBylKxh7ZVklCmRyXsixCknrj1FCpGcT/axI4Gk
+EBOwyhn1nVmYhliZGLTywvdjx8vf2HrkKsvZ99TPAXx132NSa36ojZMT9cZ9f11
2pvIejY0cz0WpeDegG4qhkGUheKi17jLcquEemB4DcYwL9T3xXcX+7RL0pHg4wNR
qdjmmxWb7mICRwvrXviUdVqlr3NR/nWB5fVOTB2WvgWtjeSTDLGLyRvLlMZ1R5Zu
Qsqs92kqqY+C7cDCeV0lVe9BJCsSoGpgrOaPKklaw6jGX1+LhAiK7aQa59iWmjNu
uaMugwSp8df19El3O7yAtshMGoaTWu5UyXlKSIyUPY06u71UniSQ6WV41iFSIL8Z
PA3lNNyL6fmSlkdYwDiQ3tyn3T7QaTQRj571no/Kf+7Xs/Mp2V0wkgQy2qNuKL4m
ZYr2fVTt7F2jLdvxCapQPV1agfSlAKAMJSJfhFQuB1Tj82XxlMjCle89dPcehojT
mkuKoHZOmSbqWB6hJvhQlGI/xEbRkXFXFBUe6KfFI3hYj2rBzQ4hYUlYOFbnTTcf
0lZGdXd4jpUrNh+EYDF6sZR0Mj0M0GGtSmj31vWIMPrFy02oq/WAYott8oB8dBiQ
tAByFya13onNfRFVrYOopjS7715r+ZAP6fCszmblrhSwfPON5+FTB8WA/3ZLLaWu
Vr1HnSvlvZaIhNM7D5FyDwBB658+c/ThjaI2IA1fsCGZ9NwlsfZCUHqPSTW8Pmiq
VriHKALylzDSYBNiK5IaMc7hlJwyEo/DGc6n2zln/8Ktgf23kAaP4BiV3Rrl2UzH
Oq9B61XJBdVUc9bwrburQYYybpdJFKTqHlJbWRxSCVXkfKggB/eJhX1tePhikYGL
9GhalJE3r73w5mykhhibGN16uGRrBy1g0UtQb+Hgtn4J44lGCHYAcleDv+3lWUpq
g2KYrANhmeBBTaFJJiTtwA9bPPxwVZMn83suI+1XWi0fz0Haqc+kXbCnNdV0y9FI
r4WuYfD7AQGfssdYGX6ogWMCSxjlTqS2y6akTB/oZoXktFkQ5S2qoKIlQLVcXabK
JgMLu6r+6xR1oHKIWo1NBswKx6/cvDom6xyVZpaefgg5kj1SbXZ5vqIvircK9YDQ
AWavg8jYgA4SRY4AItfbj+IfDEaocojGjSgUMflx0CjI5sEgRlh+zvJouBtkq47n
lsDCSPVhi2sV6mQ7dxTnXYQkifzzdhISRgZw7GFAR9AOpCR65+p9LzGPq4DhqjzL
53sMd/em+MEL43Y8nOmUYipvOaxQ0KJjVrVsNSa0OyCIUozba5E56RVhzQar4/yI
bweSuvItQXXJpY1YvcOiyNGxfYEHjfc311RojDLBF4si6btMP33WNUA2kpvmHUGm
t6Ex0e9okRGsj0S2Ur9JZvnmLY+ZRo3qUq125/uUYpl19Uis+nJg3rRw4cDlaaOv
+CMw1bpxpUruG98Xs1XU4gJ+BR21yevlnHIAkwLH7h5QfWchpzNDkgTO8sR3CVca
zSPS5LFxSkiKK70iPVnSl8tNFYl+YCqiYDARLCBXQXsm1y1b12zi74KCn/YLB3xY
FKa8CnqCjeRXrcjaYIc1PWMNfrgk7nPorGXVLYuG2EgZ2oAGyVlPG4DS+iBstsA0
j5o+FFh/Qf4pZP9xg5DedXuOeax4VXr1LBPQLVJ5Hz5UE2X0Yw4y0NQjTT2z0TPD
3CHmTfRt+GBYZ1LzIPf5d/0qyNcgE65ifElhb0GXyH9a9BcsPH9g43OCKy0Wrt/c
KpIihHacYbMqcKyv/9TS0lYTAmedd9vwSMqCd94bSVxRKBx9ldRxNg2qUCiQJ+mH
xTxdsl0TvEB9crMHl0ZgiouLWijip2OY/P4rWDKmMosqCA2hIru0Ur++wCiv2C5X
EgPczIjF+V+5FIvvPGJ+l8fCpVYpcMYlI1JmByvSIKS1B5GaaLSd6koT9r7ql5cq
w+5fzxsX00DhsE+wVterlHz5rpMbJIHY84rPzhr1W5CttMjTbFgwvFvvDdsOwY8s
quYAeOl0kBcFKxiRmL7ujnDvTMHjEHxgS9p/dW143j+fbWgvhukhrI92ypNaiuCa
q8qQLKkl4osghOu5t13VXD/kNLltyzCMXbqNhKOzkO+jFCAPEZVu0/8/kLXHYY6j
k7JMQ8PAfG6jGTqdGNI8Ma1I8oZsXme9NTNzDaRSkDYivDf8n7LCVUo8ZQKNKTJC
cxJ0DrAdz5/bZwdx9uP9tYBEQGcuJJ62of5HtxtUF2yzO4h7R+gT0OeuNz0j2rmy
PxJspkN4n+iBIJfeAYoIKTOz/EjU5Q2c8x5Mw7RCmjwxcq6CAnhl7BVDRE36RXeo
c0c+x34OTwews1gc07PEEieRPzSz+9Lns9HSrIVclrXIgmVn/V09Mppm6D56o0EP
GUzPE6limGyAq6iDFM97gbnHXRkb6GEuMQ0NcSPHwp4ML3Y11HZXfGH4Xfhex/rB
vjY8JnvsH0w3Hwdxq2IY6soW5XqdzxDBUIBH+yRHhXvLN/LDAgDCitqmyYzuy3r8
ox5SHNtroKG9bPeATw+zNXPuJuEZ1ivoBDVp7hZy8ih33WTzg77I+uXo2JJOwZ8e
bk6xtzCZCitNQpnCOCvkswRVecFEXfhPfxgIIKUvROhZf8u1eQJPkYDCxqOUie3y
nCbk+FKF/8va4DozuRuxOvD7ZP6iy0cXuVta06CcrOkvDPsHZ6bhQYG4EPH4KTgr
8FHuBi+a40Xzu4H8ocMWrE+n1PU+4EYgMyW2FsH1o2ImKMMNpc4xRzWL19ofhzgL
qLRThOcPVLS4Ydu9HEMB0zI1hUawg55iA7xOEi+w0UsXFizogGCsexl8C8AOUKKL
KNEeWOWcKODG4YDFa/vKaJAs/Z2t4DfZ66xJJAyBEY2xrYFzwHEXpM4Qzlfd0Nxp
HKOaYEZXz8p4VAwCfbjmwbXyydymn5QCUeMVdG+shDzxxvFftt9BjdIjF8SIXOvo
0W7tC3wWLbwnCwJXVvK5mWGt+DCLsTBZU4RQLThyXrq0buDkcvHw2O/yb01sCNoJ
mKCevGGNfneJbmMJ5dGhZfUxjNM1K7AGHTtKZC0rmcEzy3TsJzrKQeoEb2okchD0
3MQXrqrGS6cvSZ8SIBF8zZDZ8qhv4to9bYL9eZx/6b1yAt5k8LNlq6Sj85Sh1F+a
/vDI8TPSPL3etcve+311bZICAPOkmqBnD64w/TpjDOuuDHK3nCRFTxm2SzodeUbs
ofFXKyWdNGxhKet+f4NHfssiyYqxtNhZ+WXrU/voDybQAFwnrYkADo0hJhFVwU5e
En3aKZO7gRfj0zCCyDbST1/QD/CY2akS5SgJoYcAYFHWMkN2H6QFh1qoJ7WAplnQ
gTIEqSUjaF+g72F9UEJFTGQiARHRUD5aCdDUoghGiGWRX6IEZ4oNYj+psyd+tRSv
DBcTZz+HYSOAECaj4D8D1pNKCBxLlssaaA8QoYtc8VHjIb0deQR6HFx3OKHHtsT2
y6sJusAnMiRycOwSAyo8g2dHhhpISnAxWXfJJ63C1FFINetKiW43Q/xLy8/PmAB1
IwqycnDsEwVdr50q9DsfR3DbGgtQRQxhsUvOyy2REo3my0cwXgvWgsWOhtklO4QX
3WEvN7gwAV5DjFDIM8Ym896ZNun7T5m9i+bG6nDRYzMIIQIC19TOTzObfZG1y3u5
MjXUB9aLdPkH02xWyDynE38iKXeL04lvpNZUPyGI6crRpDEBNUrw5ciMhAddQxLh
0RlpvKtX2skB/d5SBKyXDliz1CU5eJDykMtXc4pun4GqVZVEZ2YI8jf5JhnU5MdF
sgMk0Aah4gOr5gkGGy6QhUhY/6+mQVdsoUJsLKgMc0jBm7X0yEgoLz/yKIbVtI+E
oytY7tlyhkAO1PDzvft0QHEkIHP1R41jJaLcHy6CmEk8/2i8K3EE+0lP1C5kzbex
nk6aoqvNYg2y01I9ELSrZ4tGVWuEL+CVMD5wFZ1y+WycshbIpXFuhv9E/n0MZEAu
vszBAnlpEH8cpbB90U2ZMAQnwNcFUIG2g/zGc3JWTsemIjjOmcUsDTse9IoWZ0i9
QjuZCr+A7YB4P7kuFg6QVdh1Tx9FInLNnQTmpfzj10n7GzgTJxpCrgveEnE7/C5K
10gwxpH9iupcNCYjYaYuEDPhc9KNSw9hrSBo3tqzInITNZ5OaAry4OvHxvZcczSz
clczIOsRjb8V434NrVrFMImL5Zb0A/r1XE3jPsHIpygRhq17FCP3ro5qk8OCeloG
AquyBYtjZxEvlRQiXmrzag5BMjlpP/QICEdTRSZKBhvSDJWtjhtrQKq52AQwrzuH
soEFCY1hIKgtUb3oSShqqPoD3bsV6vyC+CXShGDFAfSySPl2vPXibp5Z+PBzHktz
BlLALkPkV8R/N61rznOmflNRwQS8PK+9YZ/VfpZ5hLe40hM4bxk4zwcAqzs/eId+
i17Yf6P7MF3m8+V7E3kdqviXK+eTJHri1Sp9Byk6MtIQhQXPQtuFmpH95WL9+jMo
FyefHLQU2CeLHO9JJ9D0tUPrts5q000S7hZyXPajb+u7mXmn4SAsdGlbrFYqIOWl
+WlBa77TA675zfo6nHX15H1/SnHhk/2NbD2tL3avzcBnUWFBq0YoxqDAehHG6Fhv
9zPiQ8aAqLlWtlYYygqNMqs9XAUbQXSB8e6Bnj9wWGWSxRcxAg6pxt1vxzlto8dy
QMF2nF5etRuho/8tKvmH0hRXwQuLuZF944BT+LiXn3jZ7oHbREYAKaBmAbQ138rS
n3P31Gzy7MM+nSzxiIaCynGMy+hKdekkBzuEidZiHGQS+q58qQ1abAbzozMpaKCU
ua6bXyzgM/GljjtJZamaQBY1KMe9O/KoBQ+4VibSI1/6t83zzQpM3rH0StEO3pd/
Lb1gI/qsv6FOLAeO5W8EpZ3EPpCKXmIJe1bj8LHOaGcX94qkK6JfUA6D9RRmRTuK
vVt18yGqKCbGgvM3zpy3muoMdg0swhv45jfCWDWhLagKCV1Q6QHLrbJzrqZVSOs5
l/Z0k8IbpvbKgEO0H2tuajtCOV9lzoiDOtFBgbAeA570MqoKDscvET6QhHsOckCw
pRly64YN+e1kpWT6NmxHIEEmS7bguRZlZbDrDwMS8qfUSNj3tUMnIjr0i3bPPIey
flSfib+Axm17WOUkx3TkiaXqsTp7v7K9ofQjk5CinfBSwh9vtHDYVIvbhoaLnxzb
AFsYnun2X8buV4RzfZSxT4AImnGyXuMR/WoxNYCH4JSWjDWDpZzhxKyVty0VBFyq
g+iXnAFTQgz46JIZQb2HKQxHmkGqB5fQiYrm74Y8NCbeI0bIBQbuhe8qz4fV3qm0
3BQe0jElklU4yTD2NeiNTgag+48YudWPkPmjUdoVb9aSr1sqHN7avGqOUHo+phz8
c8gOy2jnWK/EaWsZ7C2BJ18LhT7fKvDvRM8YqmrBQr/eQ3FIadqTMFtsbRY87ElP
1F03OXQUq2L75H1Brp9N8z6JizLEt6PrAQ24yuAkkkFaLI4g8b/YVjcmXkk8bp7C
DKUUQ0mKGS6GKSx0n8vtLx+aZOdGyfuNJfdNdQ3gbRoam/G/06a27DwoUSOsfNmq
8j87K8EIP2bSz9ppuRpVNQNwHDxRXZEA319dFornlgtd9DWbiPYbyGhLdF3yKePL
Z+c+3oB8MEyfVtcSnDv6CQlfAwsiyyXoJTc4/g5mgsXz4B3YXDF9I13w9upxObo4
zgaeqSIjnvrzdeaX+IafO5xJ79udN3hE6VSOYQvXPsSIvYTkLjLb+bCszekd9t3a
XIGETuGqa/AQJI92+Ow/V803hCIoBzVYfk4L3ubE+nydDZb39x7HpcjKx/VDsUr3
P80G2Kgw7rsutkXX0VzL3g==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lsVlJNUFw3ZlT1XEjpqZjGO4fmgoGu1EmzxH3aRDvSg+U/SvH18PUqpNub/5tODH
0pYZ1LbdTnycQn8j5IPDzMxpSb1fZa2jAWJVSEUEVmMxgCZj73WuWKxSU4rifW3j
wCm/7qqJeKNHOomToy4nXOSUwP7Mvz17ceA0lIr9RKHD3GnLsGf49iG+ldJ5SyPs
n2VMoqAlX86eUu7ghx2bI4A2eYZ0xd4zQnxHkImMKG0yZxsTvjeknKbM70bTYbl8
0pW9ph5QGpgJu9rQUkVG0kG9seYWiGvQC0vn+ezYpC98FbI2ChWGtcg5INh/sjng
TMlQepBkBm5tNwGmfPszqQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9344 )
`pragma protect data_block
M1SeQdNKS+D22GF9Ta2V2WBc+uvBi/8icig49PjmlgY0IX0Ce00Jom0g3afFtjyM
6fzBm/zw86RMkUy1NyZunze/qXkFYk548CJQ3/ossRrAID/BUU6AFPT9NK3/rxWG
U3BWKX9DWoK0kLcrsKaukh/+V7b2uPYkb1FX6aWrdY8E/Sje1GiZwarptUAp3BBw
NdMhRYLVmNdGFPT82FAo0DSgR3BoXpm7lWZ/LObbyAn7hf8Yi1CYzUEF5QyM7vWQ
s7bU/l8VEMHPhpfkHktAca/bxmi8q463/UcPe3BFsWqFW88W0EQOB0+eJbsdqXsj
kd0FA3gYdPru2DHGc/owXQJ3A1wfHyvcb8r4L+TG4qOy7uIecYqjPrDtms102Bmk
jouEmk1t0jgJXcd6Dpq0Xe9zQldCTO4F9PZKFDL5Hzxro75+0v7i2+oej9MxmRZG
clmF25LOYK2lUNuV5FrDPdIQeg2/p2fksYcGhvwrpbxfjuNlFBKYWDXTaDh2kj20
VTY2MFE/Dx75MW54Gw9aFbwFYsPp68c2PGWwiEL9NgI8Yb4Z/ctFHspNn+mOkRDQ
YwLuFwi1QEvN/6PD5chJsfxtoGoXb+WuoOGBCeQ0DHe4VH3rEcZe0/ZPUTis73TV
mtDDxOGcHPm60gukfdpwJAkJrDlbpxzN+K63lzVUypxxk5ByTHB1zrMc3gMdKX8L
Lw0cS4PVW0h/EduWviRTyyp/zEUnrddDTDeW+ITg3QGUQQHfFZ1XxOGwNPQPcnYW
AF8JGvjINYP1Iekpr+pdUII7ORCkAcodAS5rSslsjdQJdeXkBpB/3tYXfPoViddg
LspxfUB+IatGqVcph0cJ2ASrNve33UckknoswbaqynV7Qj6DWMuiMHMYyGW77h3J
FyZY+gatDsf5z+gGnVPCVWZ9qTzg4M2CHmKuWYLaKSnw8P8COAFU2UPDP2ipp1FV
sU4NjczYzZmQsiU3LIJh59BBlNUDPj+ojCnZjPf/ZuC4qwBuN/ARs5PRqyx6Qp3N
w3Qi/se6MLQ4mn3olHNZKJU0hNYp2lz8n8Y0m7g0r+kd/QQ5ySSP4kcRzuqoNRUt
n0fGOrevvkU8HffzwVGDOgxLNejfh59AU9/GmriVOiOt/Q5GixmLGG2VF+v97WjZ
BzIbIWGFcU21hAciEEHkX+LjngQln01L0f5Dk+e/kqy752JSxGxGo/dvhAfj/1N9
HektAEgny8IxcGkDncXgpjihVdpJdEH7zhlsKgj9KdStBmN7uuSG76bXJoughboQ
CV8omWuEYSUv0yE/XWhEkKSQruXLjnzrPXE6grCXzNymF8PNyAUFYpb7rhSCJ7Oc
awL2q4pNhxu4hLChB+KfNnBIOko1UpOzRmoGnWbH/p5Y1HpekLLgvt9JPN3e0Vk5
9B38JSXSSodVnzNl7LR44BejymFKsodFU1liugQ0mEdKFLGQElkUEJCApQmuH4Q5
dR3Aan2qHDNn3GZQDhhtK4/ZOhUNgr3TIj6gRzZFidV6c5B1JW8F3oKRE1kaUgG2
jhWd0tuBNO+HPkrZkiWXHYuJ3vmMK4X3Au0BdG+/3jsvM4jY8SDOOd4W6fkc784s
fA6lIgFg9iLme9WPBSjEEnsw3CpstJ8hrWPuYWzqyBeJSw5aEzmm9YXjycqNrDRb
KgjPAcwZ+2mYUK8htl1UyJVzDfhJZ9Dje48SB0vfzw00OUf8PDtyQKHIOFwTx8am
6DmITUzHwbNkNkGN4EXuBeCrXLdb+2n5Kj0xns6ar4I2Q/gD6O7YGEU9F+2jlVSM
21vkl1bAp54Z3nDfyKdTJli6WHsqGDrFOpSyAy/g8DZmeHG+h1BXiDGzETUPZWVy
4T/Q4W7Yj0WL0LdRRlIbprkzDBnGKcLiyV0hzK4tqHbuHKk7FvY7RdcJFKAMKXFO
ez6i437DJiJc5ERAetgXHbEW8uQj0IGNf8ofvNGjtEeNs67p4wD2/T3VT8byFfMy
GCjKF4YoTi5xHxqolyg8myRc+PW1XG9gth4BIKvTqtlGBQeY2BilAiK5WNRTFri/
xrFBrUNkbMFraSp3w1d57PyyhuaPP5/NFK2iERzu/otzhDfk78b0HYqgMaN29KtL
40QB5yvhRnWg/z5ndHp4O70vkAReMMsKWhLXY6Zyt6uqgNxWLB3EI0VUyXVMGA0n
qwjeMRGSRWNbKwiDvpljfp69LJIa1rDEByPFPF6Cs9qGVQ1VF1egx93Oo3ASRshM
BO67/qZNKQVDRItnkuFyZ/yXteAFn87JFhYuayJe1UFy0DF98Gkifg8Xh01bAoP1
aLlaPHR3CPiDKDt/XFzqqtMQsIO+3AnLElYH1qpqc/7n5w6PG1DtX7AAZ1vx2wxI
ms3GLcVIZk5aWyJiSkca/U5Ohm5i4sWUKUYWK7571TSkHBNIRxIgndXYXu/HzXtY
KMk/nL7se2ayakw9oG/L8X0JwFJS5sKTB9tss/ytf/M1mNtn1LR233ZNOSChXEQX
5QfeoAKQFKw6w3Xy9C98eNxiv4zqw38pI8r8BX4MrxzV7h9k65rFi6aYkbuchzMA
tfsesHNXEjXZrYWH8evvQ1qbaHyN48u3SwL1sioigtl4U3E2DLYkUHvAFV0iuJ8/
L+2K5Y204XMLE+YQfpvCiGemmvMV/vApgh8/A+FK0o+iKP0mXDmyHTNbsqstjRRq
OpLJXp5Qh6pp+QYQX6Ge2sFYvi4buTUGWNLfzFsXEajpFVDBCvALwSIVAm0fwCVn
Tx1pWIktU2XpbAYOMDQMp+7lCOoVXIHnH9CWRe5DRYApuP9Cg+hHADU4QPeDQb1U
dMqac3F0in8daL1rRV8k66d7gt2aJrTiPb1hDla5JtIUvULcet0VpZDhzkBaUq6V
xXl91V//FK3I87vyjbd2wMvx7+GzwFlW1hHOXPS/o3BBofip158Hw8ZR/+Q6jKQj
wLyc8jPLPn/9tuMq+Cz1h+Z5rk4CmdCbTDlgx/cFs4fKcU8bjUIGFhDQbMOTsj3B
vwSnoHVoTK7fKOX4apsLMONJs2njEzkEk5ypjsqEt7CBejnbToIeJpWNNPwy+BPO
SwAFE/vq0+Pr5eCL+j8aSBUjByzUOCA3RmARI91FhzyY1Iln8QPKNqrh7k0xhky0
jQk3VHqPV1dQlgkKAnsJS+DSAlnwUi+E8tmJG4NFKaOpY9rkViJ2UoTwjGj+Megn
FjJexd7R+nt/ODzfw0FnXEOlbtWzVdoWrNqjjcjTUWUIUz25bXJ1HVn2b5t0GhkS
M0rNf3n97dauJ93ss9LBrNrSwaOJ3TM1YiluAAJmsYSdVxQ0lvAk/Red2a4rFqhW
NH9E58OD0sNouyBb712IYza4d7beTMf68ftrglzXie1h3/8InOE7QqmHHd0kHCYV
B/N4YUNJipFw6YvxRnFzLT50RPDAKb5b8024xwuIw9SFg12+8K5jHEpzi5NBwwE3
cI34JoJzXkyifpkYzwNCLXqDeBxpCvXAljZMo9BwHTpnTNLPdYDviPdwrI2DCXDD
BhC5BvlBlTz1s9ANyxjpZxsFqRBaHDt5dQtzJVfsxfHnGwC/AQAbsLiSiQxGyeqn
5iGeC9cyEuU41fgaz9mU3or+Ld8ixkqIfQNcUsnzOxLRXsygmSM+WRpd9QDClRGL
JGiJj+6IWLEq2alpZ8WrvdhmHbXhtvfi/vAccH03sHJpZ4IWBMBusIfSfEnoku/p
OhCRXVKahmnVUhe1KwJ+W1Z3O3VCJjTlD1yDfQ3DnWCBVHta/INGflfcXRXn2zS4
YbIJColOoufAd4v06AqNRjnIG7YbvOUlUu7NdtMZgYqjk+Bhfu4dtT4zNnruB1xb
OrW56W1U8K92wZSFYTM5er7FMab2iU3kWt/f5BkXCFOf37Bl8SckTnO9ioTDZiwo
sWX21/7v8nqYt+hjcvtPpk/OXjyQP3TIOGrNAV386QpevvdCISQFBU1dB7+HNoTL
+EkWhaQD26iA+a+SlLcdn7wOZtunVjDD4deVUmC0e+xxT0rCWdD6qD5i5UlTah7A
RdGlZyMv+8/qXf6xT4W/CX86a/vcIbKfjRVQujAMP5NDARklQhXSPZXPoZrUu1d8
9NlaPXdrMFpxGDYfMUZ8p5WdNkvxid458b30VsUmiVywJ4DJthmsI2ZA9ZkDGgCk
D0/PMEDb82lAi7F1nYS+21GBVypUgLAQWnjPWt9nn/IpwosjOUf1cc0BRWoSw+mB
AR19wcussrKxQCUPNbmD+BCAVob2IqZ9kQXS8K2j5l2nGopySfFTXIpg6o3eofVg
1lqsPR16G++lHXo463lad5RkPj92FERtn4pSPRSeSjqaWJ2zAaSk4V6US3Pk6Syq
Xh0bHRy0wUqeseUHSB95o3WZXTafBae5UiecMOxGzRLkpne93V5d8YeywV7KxJEm
8PrLRUmZIYU6+j0RY80eW0JDhHqkZGIOeQtP0zN63BUFoSaeIyZbfQE69mwmZWeb
P5kOjQ6eT3yQoPO7ffzLEFlyj4UawjztLKcphM4Se9nddByPHa4UUMJyQXmIRnAb
B1yFYvq9c5ifJHzXCzkjN4BxpglCP7p+hNl8/vZbzl8ZpWzC7uWDK9zJpeEznlxo
VWnJbRiCxH1EQMwTZIO3dsWn+iFgsuGbTPAO6GqyuxEpuZXNE1mDIKRLuGZ3X0Qk
NQ+3dGwws/LDlhUU9Clie+UK3ZnHGeoEkoZE2eujX8giiwOQVp/KZ+8kmEWHrCZR
HbjGeyxdh/h5YbRBhoANDDWGLwYSj7lqCR+Y0wSkbEa5rq+ba1cCN+mg74b9tZ88
meFacvLPafUQ5A6siqeA4N3MW2G1gsYlizt8jDHvxW1DwnvEk2EyGX7YuEnO5n7h
x0/dWRGnMtizO8RYVkKFoEbNkmkfoxLnjM4ajv4wb5iCgBOb2w4Pn3Fop2PqML8J
K9NW7EAZm4IryqOr8BXT5eS9qnamg0dZVRr5REs/GcZ624dBRCecO3XlC1qQ9Lr+
weyNg7Dy4altXySJwJr1Al0xPpMaKNCTI+x9z3nR30aN6E3fr+uB0EmcvTq5xGw5
XAXjnnKO5GtOkRnSwJnwVB675o9WZpSjCc70+ETXtaB19yLUdFCzGY/z3uF65V0M
cu7hP3IQcCa5UaH6gYKMxm8uh4pllvRJ1DTohIN9yb34GDj/13lmF6H+cEdwuYlU
wabqdX+H3rbFNoLJ2yBBjiB2rEHPixwfE6ONLnjbzrPTgGaPmZXlp058bZlTzRsF
0tF7vc7vrIhB9CSsPGASJFAAdDrWsjyd7UgH9H2fKn+7p55blUnlrRKkPLlRJtmJ
sjflG3q0xnvTMkESNJQmlQCN0oxMjnyejQE6Ujh7pndTqqFsghDC7DpzCVz4MpX4
Ype+umLMeg71Y+gFc8b1al2DMDuABu2NUASdBG+eeyb6r3dIdvh6NpWCbzCs+4Ve
xMpBWCMLPL0ugCFiZQnMK6HDloyS8E571XZinheOYN6K9VAT7SCovFNNzKkTyb0o
H6UknDSdh8HACS4usKBcUCo13EAvoGYPNn/5w4I/Rn2EeG28h4jlx4PaaPzpZ0hY
C9gKGwLPawphiwCdCfzPH7JzUBXIBT0srArGLIuShdtNXCGKG0TKIcpGA0gH12AM
ZyDOIWwhzbb7eD1tYLShW6hlhkB6j2LOwZMiFIkUGRTTSEPVIxYM9cbobqoSt8Xd
iG9jeh67oItSILSUKUchv/GQ3n58nitVOYdmBznN9nJULyTwDmJWkq8Wk/yqpCLc
PmSE67mqVOPQMNytgVvRJNJr9spvhhvqwwMyXX99hVTMQFBgObBmHLMvsPbe0dUh
JbyoTLARAkTjfQdXxrHVGo9qBXtZ5PPNP3t1iAXVqA21Y/nKBKrwJV1HC2t74p67
GbvDhVQGGZADlfVbndZSqLIeWtFNauqTJJCnpPXJiScivRBjh4eYKXWEedkMF3r3
FVjG/TNiuKTVWl4f0EKbs2/WvgKJCM2oe8E5iKwg07vBiuJ/fNxyGsfvlmJsRUBx
1GnkMUvbfuU6VYZZdqvMaGHCdqFnWz2/nFjW/9e9ShJC85oLYfZW72alL0ClahNn
qZ3k8VTQOZRjsgfa1vAxGruowtevZXXEQyOk03RExZwtwz1cvUmUxuMFRKEcoKh+
ioWqRPn/5z+5b9Q60KwS6NqEOjedNm1gRo+uBKK0k36EzFO+hXMbpGgSnk2Wmuks
CbiNgw9s2/ndLuU+YfE5vyZJh7qpDQICx5RScpMxS2yaFk9rI2YIJBrI9NqEYsJZ
U5zEib3WYHI9gtNUgWfVj3WVtkD71yyWRodgTl3LPc8GODX+24Jt9ffW/fAn0BX3
pGLGGYlKaxEKDfvh4DWlhO7bF2YRZajN/4ln6i1hTL+n/g/NclsTjhfA6rk3GVRo
7tNeIE6Du9Ezj2s3H2CCvBO06WmUl91zEQbbVJF2fe/oy0RNaGr2S7s3Y70r6cMG
nprxvi2SQzjfSyKovY1hgG3hR5BNu+Iu1GsHe93CYjwZLLLQVDWKdUmCn3zjSSQd
oXQ7r7b5v3Ss+k09fhHKOiuWPPJsVBJruf47XpAh9vW3jMEEALUBoKRU+ASTQBKJ
7QvttDwKCbzVgP/ER099PujIe0qIsc50+4BZBFE/um1hrtcTQPhlvocZZu3CzsKk
jCX9Telnw2gs3w3umukobrkEGJi8euGfMfPn+1GHi3jz3h/ZTgQR7iGqlACUpKou
5yQnKDg7xherGGlbBVv7QKCIzKEUOJQiA/he4P3OtsYc0DPTE4a9pAs1OXy5QzhU
Z7XOYweJgHibM20eIZyH8I42IBlW6HnZR5abgDt6V4FfyH0FuSHGvdGcYmEyVr0Q
vp0w6u6KtB9Gv8w1yMNrfbj3bR2C8xov9XdXrkqlYtopKxHtwpXzcm+KJiEjwxi0
yOJt7mQ4tsiFIE8fGCLzBKVv4jkrlktmyjZzepevu73AtXOvo94Xzin9HX5eZIRu
8jNYKbqH5sXQlV+ItctH9a8WVVaXegNNlPtWL/84EWN5wAZvdgRbCFKTAhU9+yMI
B4cRs50dJq2PXEEyalCIe8iMJ6fk0TkEoSfXNTY0Symq2pCicpuFngO4rVzLyRX6
/NAkC6W5V/ZGhIuOfz+2Llc0IkxcrUyU4ECXEdkERQHOjdK7MYpJly98dnZJohZ6
fXFZKeJsfW2UDwFljqEdijR9YbhRnAScIO+5DL/MOLpO42tgGchIpAM96Il0v0RF
waZh8e0zPdAH+5B3+tyFX1BZ/1Yh/v7aAaHa+APjb6NAY6Lx3P8Pu+SZYEhVzGn6
nPANks5VNpEXxkDSIt7CEdfQVRU7Sqe8QgNMiRvJ1FoDhGxUXKQAxuPmPUhF8N8C
5uqkIpDlOtvuEcbsQgPRv0NF8HNbGTVMRSqmIpDE/Bpoht+Yq3gJb/7yFiz0eO/H
bdE9whZS9Z4O3qjI93RlaPNsqNBWQ4ykycGcQGnIHz7Tx8jgfY234zkqOEPWNaIU
YAjgCRInjPqI2HTU9GCppIbxq1EwnVuEq4JddQcrZDheAbl7t+THHoRJA4Cv3+Pr
ZtILFgri/LdDI7ZvFuAWOwYyR0oVD+IoD275BsC7/wtXSGY4HXwJKUYdutWWdlYS
G79SLELJAGiPfBlK24i4G3T3J2aabEFAdUBSnHY7vmdCt163rp/cZqwdSbd9kDTI
FygGhqkSAuYU7k4rA51F4KQq14gURiVIo2CiOpnuLLzO5m3FxzHEPJWkf+mbx+eB
LjLbTZ5NcEb2GHHkvbvMByRXlUtgtVIQFwNMkWMLQsk+BS4FI++1VVTHMqtocFS9
d0LtdxjSI4yN7Cle5EQXBbhIV046Ax2352MFF1DG/z12YFPu1P+I279avO+LRwtC
BOAuNRlnq0l2zOgHHw1bGQpul3MhFFgBIX4Ma+PWHGRCkbG9IjLTpHZGjHT7BD4d
gR2hK6BEjGYWHVjeBwGFm7wKR70QBeLkot1FJMHjZi/+JZkw/G+tLr2ySpV4gOmn
CtW7rkX9nbgeyc7S6HIZSHi/06S2IxBgvuQphNN8EiTJTJefIDu3K3ehhmmIn5Xu
/FesklFw4BMdjiYHk4Rbo8arkG9I3k4RN7wM2VmbgvL1n1frH0nZVXKRkTMnXi9K
l5b60tzKLDY5IB52Nu+elnbFIWQnlbndINDn0FlCon2baq4Ee8gF0+KfCvNC1BgQ
/kv2abDjMwOj7LmA+vLC3bH3SChgSP72TtG+4Q0Y//1o/J0gi/VBQEBZx/OKnzUz
FRrB9QTenaxYfD/aeee8dYVIyAH/4DQ0Shqt2gsrZQty8CMeA6COG+W8UyyXzjED
9vdGL+0CBco1K9t9JnZ5xaCgrP3FjRSbhnTXx68RSVwinSQuVB93wYPd5nChgFmZ
/JhUdOm/pa5Ki94evkif1HVLjjJ+JXvkn1wn3W1+e5vgtETAniB1YPo56xn0QagF
nhlQHxWutmjKfr/TGY6BgsX0fg+MvoXWYVfwxKQUOhkPxi4iU7xc8zaPr0NLEXVH
rSybslCKxLZtWSaza8n3PMQYx5x1Vr2VXFbTclcyCuZ8CoDjHf5juFkERWW2a4DB
Uxzc5Xh8cR4ZMB8Y7DMohiBOzkJecOy4FrT9CM0UEJRNUwXFFu/pIfV7MrZc+nRe
LDTvQ7Wa3pAU6Z22A8VBNY0fXgUwwMAgqhaEJYUnSd6fv77ztk8v7oow1l/jpn8B
sxUA2KEkyUiHE8mgzOBcYYAwo4niUoM+maejrwXTbiLq3u6vuEJiIxWTZAoH/LRV
OB/NRTMvlnOo+n5vNUaxeq5DCJ28K+z6GVd+AOHshvLAn6bvs3yAxotforf68xDn
mzHaSgU2D9tksFXAeDK66jRqfkLbNqCP5anQ74VYbHpswfwJ+DrNWQVbtZJnzXJK
H43CAPFM7DAyI1lu6Z37AQITBQaTXY4AvDMi+fxbfa0d1uMBwqu5sDiZBNyMlJEG
VsmEokJZP9e6WwfP/qhUkoQLaUf72S0O9Hl7S0mCHqBIqMhGG0g3nyEOqplNf/0a
HfWfA/zusO0RKP2orZtrxH4i/KvEIdYc23+8JvNbuqD/XId8nQhkPoUGoE50xTgM
eRz/NpEcjPYyFTmslFY10EXv5YCFKXVHaWv40bptxbP0XFj3JqHWG9CRujooEnk4
0gwvXOLjv6nJOb8CJWd4vBmqC9JqPNT/KThhVqMlaMF7mKqydgVIfjil6ZKCJNas
Oc90G0lQxJFDOTsGg52FFTq94LSWbJ1uqW3TL3k+eMTfaydj+pntm2CNWlDXLQv7
zISziq4ck/xYIzz1scGh/5nv97iB0P4iIJtM7WcZ5Rnr3ajKYB33IRgXuPh2099a
Hoxqaw2Kna4gkmJ0Zac4xvI56/6kKVfStMk4jKgNMRSdXy6qCMRJcwvBp70uh5Pe
RE3shUCtnTfQolK2kgUsZl6d3gRMUo6wLRR9dwk0wuhtxDIEtLF3wH/s4f/gkSGk
yChtguuCKFvygn1sR3G+ZShlwYm8i/wukgB7hSRvgh1x4POlk7pRMgs2uKdpUACK
aQZprU4VfCTuxraJbHzv4VmijMqC0S8W+5F/CFket8lP9vELUOYRnXUDE3te/WDA
Udz7NTaJhdvf6dEFB+7zkicluZW6IaNs7u8rITYpozENi5TQHzkvRjUhnQbOW9ao
i6UmowjWtHpBNssiROFneK8Lx/5v5/iXrshw8Yw1SZNIH7yfPmHBHoJEpTfr+UPe
zAOJRHV1ZoJTVJjjr0i3WKhmfHirfLftnzmVUqNFy11YugEjk/NpAPq9zUMyOFc/
g4qm7Cwb/DFJgzV2+JQSxo6p/SJUGFoku4KrLomeNt+8zDSrnBALBuy1/hkNnbYP
jhCeADEB6MBIurtLhTI30eeghUo9nuEfUdx9wavgUqFYjkkHmxIh/hNW1JGDgS72
/STR4ogDcrSrRq8uUP0PvvoquMpu5/g3syGUb2DUsUf0U8VHDCVu0KId+EM3wOF8
Unzs7quWLxrmksHOT6JyZ+ytUo1y/u6H04N0NYQbEoDNm5La/cJEpBVdHmjJkeqU
K8VAs8znVyb9+tKxneoqi9y6tlPY7q7UIRnGCzDwqmXoIuN9GRki2zpfMY9/wSBF
VbZp7lv6Prn0KTQ8dmo3Clmg8q7mRtnjqxECRQ4dqDUoudOwImlzEb24wHbJIfTe
ecOnUE+KjORPJYNAG5BLn+TqAm6MtYR2Pl6VSt4N2HeewWMgY3NRsbF72ObcfyZC
mrvI6JCY7j7w0yUfATzQ+A4sktFJxhvqvkHYod0JMhNVj/WaZx+nnO/K0k9urwGP
q9jlA9oWSWNFcNAyt8jA8qJ2OKzAFC/54za+nlbB8McwhEkPn2RD1CQaH7CUOowX
e/hFC07HDxK2Mx8djsnDPX2r1NzvC/6vQMZMj2RnBn6masSmUQg7T/Tl2MYiI9fb
Hx/2qm9ZWl9AM+UT7/hhghxrx5cYYPzr+POrvt8xQnn7WynZZhk0knUVg8JWxMhl
klcZD1t4TrHeCyzJ5cLYesjLNZS9jGm0r3HQM9N16PwWL140Aias7MDALw4cq4l7
kOYV3ySHVJrvNkvRgkSQ/L7xJe6t4XvvRI3+kSuPFNfe7KsdE3taQm5zYalbO+zv
SLhS0uP1BzqV/3FOqruhzIN1K8PUaZGzJJf6RA4sYMz+Yu/StkivDlw45g742evj
6PV8mVq83vPaVecEdbCdtJK6Ges8CAi91OMDfwAb+vWiAl9AtCfkRfioUuUejwNz
wnb/EeV3Ai7k2mJ8W8BgZHoNrdui+30VHwiqBRTMMK9Jb4qi+7X+yG0TVYdTiNAo
KbraGWTyAwKE+rtmi+1iTjYsiLce4AwYfBj5lSK3pOirVs6Sh513LovT+Olqy/ZC
Ou2wtZlsbSLf1AzjGsejiC+V8+NZviW3SDaBSGuCAGRSFRLNAQGp2oEZ2Uho2nOU
oKY9ffANRZ4hmGyKKCtQMj0VYW2NOCI1dW3xmdOfZJWpFKYxmB5Ef3nrwmkd5v4J
eOmBrV6eYxI63aO9x5uHaRdIeAQPlS3Eu2IrRhNBCzerXvDA78qCPNOmZiLXLlJI
n6UZEFAD+SIgkrBjdNLERyR66w7OwIzFNg3yyjq+YjytIShhdZ5CY9Slf6/guBSo
AxEk1mhgkT09SJop+qUbF1Y0A8zAgLfD82FTgc+cBIGx3EtM+97WsY0nHTOmSxlz
riOpCiiZSvsh5BJ2HoPkN2EkHSw9Z0ulTOCKM0ONnw26Xl3RvxITUKxN69HYNFUO
ZXZ7fJcWSHYnarB7epv2UnRaI1eZEeClzWNLl5mDJI5PHlV/JV354zzpvIDXeAxN
W0g4V4vieRrS78SgEzP36Q48z3DUrbczLMprcS9wHPmMJKVl9EOH5bwp5/WnrhmM
6dgIr65ta1lZRM5qxugqJXZRzOwNLwnMjCW9NbCZJq2YNGzeN1scQNaYPVsFW5iK
Q8qT3F1XPC7tI5ddToLjrFmfSjY+gDw0jibnVwMmo2mr/nyiTyYRJEflmu67hxWa
4FsR6qMoswnMSoGjHT2pqSxhijnewJ7AywCgEbtLtHASZD16QEj0TGnKh87LkuuB
cbEe1GECy4DFnVMS1QDEPJUwmi0MIVmPJYgtIaG8MppLfsPWJS3pLOaLe37kdmCU
xgzT5bSUyP+yw5duYgyIeEusj4uZzIL5koQGcJmD366EG/tdBpI43RRDJDZsRvGW
bM16BL8sEYKquy5SAHYw9xB9/znFfAkAYgvFqY06gT+xCT3ri/Di5XzMOxGLoSGJ
Z8Ub9uPbZogNj1PMpHWQsVHUEWuNHpa501upXVIu9aP7X8yzY/aR2c9L8cOhufnR
ebOJUulp6xQYKiquBvStIuNXjGvcdckxp7OpQb4648OeLb7fRa9DJNUUI2ZRjyES
iA+OFMzerFZglfEf8u8m0DR55fTMtT7iYu4bS8e+unkaCSicrd+hqe1Qy3+ldCzV
faFJj/+4kTbUyr8qhwbeTQgGTSep/r/9eqLksi6Nes83qRoW1wSU6qxNj45TV2oh
byzOZuzFAqcLQl/VKJKU7uowc6dKEIvfKY/sGa9UXkP7z99L1UfcpN8FHVTas8iq
bsjmVdErago8WPgEvZoqS5Np880kJLnQ5d8XC6q0ZgEMyyvTazpH9y+fk5zdlhtH
q0G3h4Kyu8NNF+PlJB7SoGipAaCDNVcF04zPDx08ERSpDxt1+OVa4nnBJsWmSc2S
xsLMNpn/JdsInJh8HZaaNGj+Wk2iROOLCV71VSAUfgtBvrnzh1+/vNKh19FU3txA
7g66vbPWNDQXwkKMecHlqErfbI/ENgJTESQg+fyiMMnArOQGK6JfUi+L3mRTEyoX
G87w//SXdUYKUzZVpXrLW9Z5Verfbi0YVMktGJRwAhV/4bDP8nGxmN3XK1OdUpPg
sPgKMo3UgHqjBdZzEFjJtOk/LRNlVKPm4er82BF5KFg=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ZJZukCFNaYZw8b+XeL0H3vLVeO42+znYtNKFb/pd0db5JBPFJZZ2cp4twzh8maa6
wdlg51mJA6E1OFQIx43nt9s59I0ZVLHH6klWOZ1kRalWIqhteJLZhMRvk+IsUNZX
Jq2u0ZiUolQkofWLSRbwZLxJFlm7W4vzWdcrTqh42N+ROVYuvGu1eb4vMV5SMc3L
Cw183KkxCrC2q1qDvoZ4b8BkPrH9+yCZdT/n+SAGpotkn9MWIS09nHbjz9+EclK5
yEVJX859xCfn4L1irFDCJ17k+mOeez/zAvgxMioQGP0rZgbZcMhhBFNXspHkln1o
ZIyjJ9YK4FChw+4CeunrwA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10304 )
`pragma protect data_block
EMQl6uW5ObZUHUQbnP8mrZq7qDaAlnFNyMUoC8uxxaZBBcZ0AtCAm089egkjF7jF
h5H3P98R251RqdRcj3Fxsvp02Fvl/u4QiFNIf924N7NhuhZYo6e9YDDC4s4dTiXg
JnRfZy72Xj1VZT4Ztdqs8wBH6kqWCcEaVCHZk28xWi3XjUCwzVmvWx1XwNnIeDwo
HJ4EoWKdutTPo5t/O+ljadKOnGeLHYyB1qd9ThrKUA+HQLIz7Thrfno2IgQnIJee
Jdvhm/RQKfwdx0PIp8Fj35DIss6oZ+HdkXhmsXssxUW5ENPIdPS48WPpiHdgIa2f
xdarcJY5gSmDVzrqgVfKE2MbgpLen4NbkKu38kvDsE/FILGYSAbyCURkt0VsSWHA
qIEaTMAAh27Zz3hsWe1oq0HtQ6HoHj5eMEfu9M3fgRdGcxIze2O1kJztH8BMKkJz
oD9YPyp9p/6iHG8rvhO37iVV1w8eH4FqyJZbtOQAjI/Pa8A/rD4SHsnyn2E37DXQ
tFvKIsJ1Y3GnnMg7t+V1t7GYF+fvyC8q7z0NpwNJUEjxj/hA+Rnq10XUzvmIa+Cj
NJE0QAPJtBlNlijoTB8g2QdrcQcKikOeFpMid79gNW5igNrc8I18aqEMY7js/non
zwAVmfHHQw4/xaqw4YsBSox664mi7VrOeq08UJIrNx0LA2dp5LAvpMaskTqLG0wW
4Qr7RLaCM/eEN9IqubqEByrYDAfbkg76g2yg2TftI3Z/DTEJKnnJxwjZ2ecatbnn
NDFmQRwogqNyBY8ohbSaP9GnqC4JLpx468MToq2NTkIp/pzu+523JhuwMahCSzqI
vMavxh6JhEdmvNmjHn7lTTDoe99Udh90Iyl/yM8naRauDzSVx2s24C4Zn4lIzVr4
MVctxmYYm+GJ7433knSkxmFEUCKxIXFO+OQOtjBUdXfjfGbKgByVAw7hZWBytYD3
i0leFo9QHqKVrx9S6eZk5ndwihP4ugAxrlBIoQwJnZCWhLSLOCGy6AWayL8cDzZh
p1nVVzyrfzDI0BbF5K36v30x2cul4yEuA58cBmMjtJt3+ilL4GglLgR1+6Krk4ah
psf/HCy6AI+fRXyo3VwsUfLeoJR49OqU6qQv57gZCAKOczqJ3oYT+24VtVm/XznC
MlfaiAimDDVXHHAT5aONSCV6HHUQ1yU/tp12Y1rKK/tdJO/epk+tI22ofUnbdF5D
v6OcCHmJVdFPThDOIXuKK3VRVTshjLeR0wDWzcIqJxIbk7p9FBIp4mseqykfci2O
UhuR1GHNMoDBkPDeBAUmCoGRsTgWbN76Iwf2g7Jhx/YgS5n2Il4VZwecOQpHtEyC
SkZG6UH1M4s/GM2j7Dq6ZODX2PlSxnjST6UXaJISaYKEwOWNMYeLYECbAZQft69v
k+IL5a5vqH1I+WRYIsS3GZTPfji/yd7osCAR5vz4QhTNrrZH7xO4Wy+fPZlkLdVU
P6bS+gcgJ6npvJUc16+coqRWTZMwzlA1ixIFaEfbtvKNaOia6cboVdSyEX718M+M
dcDv0Ihy5nfO7cJbbVI5LBD26SmdDXW7br/UrKGjCzQypQWLd/+Erj02IsTyBrO8
0IZ8U3ZZzl0+wSS4i5Stqhlimt1bpmi82/wj+tIF+S8kJIvU5rjjNUBU2qafhlMe
+sGIlXSjgW3Zvu2xkk5SqlUWv8MStVC04zEmsN34TSCoCtkKNbHjE/G/OLy8mGhV
QGZPKaF70Y5QDODapx7puMrerFDKDSb0ChyJBF+RKIRJib6vzU4twVZcBCMnFUHN
cPmFL9EI4PtadOFMoWM5vlYNCxBxbNz7KJurmgf+zKhkniTjJTKiCeI9kX5uukT5
2psMA/dUEZCZU1uZ9fH+elvm/xMBGvaRmxxFE4lAFfkOUYDg1GPcD6IE587fQGAS
KS+bk5nlzi1H4YZsZ+F5HO4IxH3QyTJdKyA8nZHllc/RJaoFNfV2ymZ6yT5jVp7Q
MKSWpwI5NhYu5p1jxOTakWlcYH3MLb7BguZEnABATPKIa/VmjEviAfwEce96aCBu
zcPdKFLz+SAHwGCWDaosFSWJ6PikSEQGG91XfLWuTfq/cEJUonzDTUwfZP1QzDLj
qamvI2UMRxXEMZFGWqaorbmi7vULoi4cDb+tkwjMKuWAi5DbquW7Z4w2DbnZpOAh
49sxgJdAOS5pm81i5odzJOnl1wsdw2wO/6u0wtGgIOdqlab1LyTocy0trVMf1ydO
nxUt6B0KcAS8RG8Z/k8u9JrJLt03hV382Qf+TYMruqtFNzthsEllmaGr5O6odcQH
zwmnBE10imH6D373C+7wLqsQhR0Pu4lDIko5iS2fWqGIVklrfbSIQ0sXuKcNv/6A
2+5g4KRbmYt6WcH32TEoCQWP5yGGwrgfYplsx7jzFcRe/ufn7TbJ/4j7cxB5ol1e
/EdpMFxWqtSboqXNrwo1ii9OHBFvlTqkvgTIM9GYP0PgC/8IEBFuCxQfvAaayEGf
HNSqEtJDWaIG85igA1CVoQo4mOjQ6sQ9NhAgwuGVRssjwt6m+Zo4iJWZQ17NssK9
XMnj+PNvMWWUbXmhnL7yjs9Kmw2WVRt2PVdZJZW8YyTnns1CP9+UKz8VVQnYTvRq
wiT/fHn5bnHpaFZlBPhNsVKOZ+E/QDQnHrBxEF8rRzHAu0tDcsX2CgoFOK9tGhZ/
A/KVajtMy6RC/J9gMvTZHwhpv/aDhZQSfvWdAjy4Sc0QbRP7GFSN7vKV90TOKxSj
WJ5sHwDpQyd15kKAaBAUB+6vMcGYDJYIN7Gz3Ui7/zA7fND+S5JIZ0nMGE4XIsVV
FEWUPdBK39i+Nv97YaMaeG0NF5aD3szBqjQWYq/VsN3jzAl4bgeo5Vt20LbE/Bjv
hf+I4WKQymH4NjAuX6LFsk9WlbM+VA9+W0ynhBH3zHowEew8YdgqhJo9tvy/UDCn
6xBSd/6eIQ/fJ64pvb9wUMdiF6IFOZ8HHNdK8gY0FaW2kwdCyiDFfUM3JitK+ZZ2
IsJLBPdYwNzzkJzs+8R4xhhmlu7lpQtp61v0b3zMHYbbISuVm+CD6mLsEX/Yrfrm
Kz/kPbI5ViFNWUDVwOP8veiloGvSROiZC4zFtTsGv0FhDYWwx2dzl9EzbcL4/rHg
gVTIJCS8Grjx75EaHWraY25S5BjCntFRNLm+6JuidC5Lbb4StV5lOeof+NCJvZin
Anu0sVmvZyrvD2ob3dZkeh7rYImGnoB9mPyqKhQcZ2n83YtnDJUBhP6o+lobpqfu
mwVw1Y+i3D+fhm1WjtDfM/j9FC6txU0cvKMc8YDb/D1Z6b04xj2NndzCgnNA+tT2
t12S/k/XLHJ7BRragNkPezM03scJOZhTGz5X2EGd8RRRFXSFxW3iDp6nNpsurr0L
W3P2xLvhPBxoQzNUOLiR06Y4yX3XU1qq9pv7MET3sx3bFmot9LJZ2Xbo/w1ywEE1
qC1vm9tLY2uR0EpjSO7FPhJ9rNI8av6gfjI+KGfexZLeISeQMmfpa806spudgxjl
q6GEqNQtEZc4MDRG1cSeSFsxg2/8MBRsV5f6L2OCugrq99ck02u1ou36lxXrgy8q
LRMQ6xuooTfnhtLfxu3rUSV5BrJ6UbEetUXRrYWUFm7vIy4kC2bjWch/liXJavxz
qajDYveaLDvRJsJUai1YgLcRxKUoigX7ATTB5e9wHbtLLu0CED/w0RZTR1SX8j0O
TQ/wRQcKYHg+1Ae1sEiXWKaW/jIYMIT0JFd4EFBKLOdzTEx9wsXyWrIL52RwNdJz
FCTGuYX7hH4z0ABW5roqjCDM5d80nO8CWO4ttQPr3kJIm3Ozxt/k0IIBD4snRE0S
Qtyp3VWBPYtqBhYvhjL1sixDsmo5XzjxqTmJ5UiP86wO6LuxOIwfrH04Q5VJplW1
wFqEpwQBVAs4fc+gSFsp4KrYD1KOYurTxfBl3wZfNhAJl0Am3u6LmzWCzlPRav5n
NTLKQjfiWN37wFWmpjcZTBEW1IGpyxJPcyKKmN4GDhlDu6406aPjrwfOmS95W8zf
bAbPNB15MAh/kD+1j+eeMIDs9LsttdsIYHq0Y8mW3/u/+NipIn7n87JrL7pwA2Op
cGk/rntQtBZNLRM3PXwU78R3lulrpP20WKW4EopHyo10k5uhcNCSkzRHMHxeNNyv
F9rJcQYc8HO5xALxGc83KNjKsfM48xzjEGrkxcPDIeiBoFWRdjfa2nL5Ue4rm9u8
8dIVbxPiEhIdn7vF+U/ey5rlqzkQ0OVQ6mIhbPU/Obai1J6FSMsX3Qcj/tjXtyPs
yXS6zr7HW9rTUIRpQ7fY4L5DX7ISUAFv8bBeJgIDfGDOXc410RNMq23Zar4ihfKX
IcOw2Qqh5Y4ax/HHKTP9fKzDKlAd0os+prbilsDeEapMWBScrhqzfbSVEVU0foz5
W4COAAtxLiAE7tVYkOChIqz3Kb0GyVhNSmUCdQRC0VSPBSbXVvB3Uo0L/y333wZ9
nB4vEVwfSr6GW9mP74294ba0Qi1WIr/rDfUCXVqnFToKQGViuo0CtLlivEQGC8g2
tXsP9Q1zwRJoaUHFu1XkIEGldXBPjZuLUtwSDKNwzVofDwAhu5jihDRONvjLejNK
582/uDtRy09OO2n0SVjbmmecppcd20+kD4KMwnIHXZktdmxGipgkXx7La4kM3WGH
S4DMYwXuWK/VVCHxaOTNVe5p8kgT25Vnjj6GL4PKnSH2qGkxltxKYbNv0ZpORhCG
gdVAKFt7/X1VaMYEQZ86S7bbHVy9Nw/dn1sX6K+oQg6BCA9fZsdiPXE8ikJ8Qc++
lImk6x5vgid2aR4J2G6HaTPjBmh40rBFT8QF0rcb5IVKxq82hhV9yiijayOf7ZZe
b6GriTS5oIcHlGqHDgBlUCPk0NpCZJv2KJ8swxD9SCvp6JNWWQhrXDj3IqalDr0i
SKQh2hLViqCFYPrNe9PuPVhxQyPtJ5VZ8izN2mMBCcpbpfmDztWmn5Y8nlu7KY9w
p41C4egTmNaCo3+sCM8DvU7DwfkwMTh8ivj60wywluBZ6l0c5U1Z39+npu3BEfyx
1LkAhC0Lg7AKGPr8t4DSvHMXxV+rmqx3qBUuXMIB9ys0OvBrHcf0TQwif3kNn966
Y5qDkBgHoyH99TuhVVGW9nkG9nzD1sQ/hj1hzg2j0Z1tsOgMbNSMH5Uw6QdOFmcN
R6FC5KOuPKlt9raTjcKz/pEFP9/QurQ1SPzkdZuHPJrPUl+RdfobaRcPzV/DEaTr
4Q7Kv5t6h6+Fwv7F29LAXJ8UPWi9a+RQDsvH/XNOzx9kfOOrkDcYE6k/sGszSPry
6dCNGhavcQ/aa+GCsULlR8AmdnbwbvJyY4/xJHjKXEvWuA9Q+eLpiuR3YkmoXSD8
2fTlIWmy68KGmu/LC+ACOEWVESHTz+SzqUoH8CNFTtlx8smtSFjFMXOPQnRu5Ywd
+cAzxWUSPjIXvRD1OkvPrhk6uilv6mgUbH8IK4Yio4kE26yDZZpMbZ1UaEETdZ5m
z0TyvTZqEbluwA7OL3S5uM2taSTsQXt0g54WdJQpgRaNp8jBvvlHlikBfZ4ZbWz4
ei7scQoXqunSHkN0BOen4mRjDDaXfNEv8o9qmn1AeiOXCN9X8dMN1rmVzlGKwIrN
htlBPsoZ1r5AL1svhcr0aXfTSiBx9eD8z2YjXYcBqvzSINXtLUyQCIvxhCVZOpRa
hHhqZnO1nOMZ2cz8lDYyWHnM4IVkJ+3Kp7MxRrzRwpe6AsrTxB90asspfgvr495e
eZsXl9kpI0a00A2xiRF8gUB0t82iBSkWwMDzqR77qnoIl8hrrQeJE6hAdiccJMo1
NkWctYfUNDQB1TOBQPVXcQ4vczyFE6Xwc9w5XRowRquv6PqsD+/2mHIiJkdpz0am
v/CVLsdpRt2bu1WmFOu94C+3ytyrXwmjS/t/X3cL5VgvjFiM7e2lAWmtLVG8jOQk
Lcp2V6IB98LReGax2ycZd20o7RfUjiGnBvj8OHhlaW2OGUn3mNFyonqnKqiePXQd
UZaLii18xAoIfOVX1qWI8G/zxetc1iw4lxYYbChNusGo051POpk3Q276KCbE/oXC
hi10XX9e75EwFXnd+mlNqkqHw0wUVgbjr5gNznuL2wTCqe6PnsVtx1ASBWL81//V
GnqyE85cHwoV4p9oEVW4EFyI0ALHAnGZZDkwdO9bdPwNrY9oFBAQsX+xs3lxd0q/
lzIC1MN/3OVF6MiouXy32GAfF4J+89Fyg6++SK+O+XHTuu3tTPvJRg3SQWD5vHZz
+f4Wq3edup/Uv5QthnXieUSdj5/4vvYF1vIBVHbHSOYzND6BhbbyUyvbOQJBm/WI
ZIV4pB6REDBX6USJ6XU763aayeP9m3PX1SDSTRtqOFFdRbhEo6Tezlv3PveSOIvK
k+gf2zh3ZlYdHLBSHhfsxSW61Kzuubse+sIjddyMTxeCUgBBIx+sSW0rNJS30Fin
2HayWLet/sJYEi82ml6B9nHHbDXO+U9is0IHdM7u4gj+XJY8zN5xqwxnldSpa3RJ
d5Mchy1jIyDuZfENqaJDSqY3l7mseTmefCaj7naTOWm15ry79jqZ3B+VyvUf1aYV
Yhenqnc6I7J5Qc0N1UOhjFwm8CXA/DWovStZD5BDbElvxgt0pRlH8H5ovHV0ST48
t7beRqqEqVqNSB0Qu4n/nqloHfoJPowlNn5MMQV/d9IBuws5Ldyw7W+YKL2ULjWS
FrIhBE7Bq7+uCgorgpAghcbog4Q3fHs9OVe753/u6ISbDhXcJWTipebGwO606tkd
Uqy787puiMMGPa2dB+AIug7hE7/M7uPYJNx1c42mROIQiZ7g17kvzKy+1Hbzyc8G
DnhV9O+PZJo0py5jfmem1E3JIZruC0hybyzT9zfMWRjgtQ/7txXFCIHo8gCoqCzu
bYXBi5/3+3Air/Fm0dq8XYnFN7ulWzeUOXkiDsu+ambHbel8JyC6jpOMZucBH6W/
4gaPGa94VVC2PD2BLDLcihDKSK34Ud2/UNt1QVkEp1ArJ+DLd+i+S1/i/WvAUQt5
QoQPsNCk4TAXEHEasB6qObaN478BIOGE5Awqok14jOBub9cvAeVujaT0kWN/sirG
+CtUuBUjGM8GaWiu++JuE7Lsjjic749PUJTwWvfyCDmuyd8VVm5xHaFo+l6e6oWi
uTlCNw96hEcZX0zE9irY7s10vP5qn+HCCQBPh+kLw7onceW9GTaJh14ZnmTBBy5f
ilQkHPKHRcxLfY/wpQLegkTcKH7veeqy9L3uFepxo50bRq+K9W1AL1gRPqxV8Ntc
RQHZPJrsuDukqmbpeM8PEQDyCLRr/r+P496FC2e4UdwTLBq+cgttUcL97as7tdeN
NAstHZhIL4tu38pxT7Iq2rVSY5ZZ2UkGpSUkX941LvA53r4hFRratrzA9G9CQPvx
17SL/sqt2BH0SjpDA27fX0hw8GNHg6gu9uIwM6PulverE/xXWFqNW8Wpa7tMCb49
v/H/p3hkHYwWvI0Ch06e6pErN51sjjffeFmJrWCLnUMd/NjuOWsD8s7OHfj1i1Xx
oShQn+WLXQ5fMFFUqInJAbKNoyCYuma5zsJeLw0gDHZxp3/rxIzW8yqK2MweR045
VmQbIVhl9xKmZBxDGh69uvyiG7nU/16SyVeLaQX+WFvheQ82POKZIrB9ILmIJ3Qy
AmN7aCK7RFNbDfnyYPfZcC+vhJpn91DxrbusFO6xoT91YomNXQ/4DlS8PH9z74Vl
lxbE7q7sMsfcBSlT9tr22iBa2+E7fEhBDk4J8KsGJSYM5qpr5drTnA3uWiAh/Xj7
p+6VEfFnrIpcNg4/wya+6OQttDhgptktXNdRxhRf5hqbauUPptWm4qKH9y+BvNuM
IBwOhBcXJ0ALWJg4e5yCD6rUNL5dyMibkgiOcP8AV3Uo3p6eSQSHjGLWPLKfaU5Y
XsXrvTuulrlAWo3KKXM66Yp9qj++dKU/MAeHLOnyDrhTWHT5e0ASC4xHb+GYnU3t
L/OwjGeFX4ORy0bLAaAdE2oZHPGQh7cLEJbPmWoVSMeXf7hQUWrKmCRmc6pVdP9U
tu4e1r2ZbD4qOU6xHxdPMVPaWBNzmY4COdEBHbdSdA2CFmj+BLRMIBVEc1ih6B9M
plBbGACYUuMAo9NG2kmOvvrEiLgkM/ccQPuDVl6HP3RW+VCyFuGaSRXq23R1dpNK
ivVM6r6Ef9eqmbR6H9WRJOXemSjt/S3Oxcbm9BGO0/Xq8KrJjf0Ff8B5ACIDtP7h
nHo3ha6yLVGJgysc/DRpzS8bHqNPQIUHmHT78CLyjsu2CIBId9oWssziYZ9TMhwe
AzdlCraXuUvUVWHOonDS5oXPH+WTtweunUM2UYWziyM8J3adUs4TSpKnSuePIW0g
ThJB6sy2xBkXAz+viJbuuKkPdGcQUqlW4k/AZ7xIyhOBpv+wfSB2FkQY2p3prndF
IX9Oo8/s+qdubNCkdc/ho18ht+g/e+7WLeT8ZN+Vj8Zqyq+pt4y32Tz5irJT/Y4L
NWhH9wmftTFyKUIqht/jpIzVk/8x4HqjMud9uzAld93YtaNgoj1PawEwaNDDuhVR
d77IYa5R17e7/M7ZL6MPV7VqOm17BUvvcItYXX2JwJCBt3MEkl4XvrbMXSuiVTan
CLBgTm39X2Tiq5D+FHcj8ukl6buX++VuZVa5AYhtQzoHJ7B/Nj6MVYmyVP9G7mt9
9zoouZz4BDdNwUk6yHOiRNxQ8mRzsGY/C0g6qy6VseamNRb5mt1tNMcfjcf15hmK
US46XfKUAJbwsuwqzjgrkdq5g12CIivoZEmJqvKQFigL0Exosg3/lEM32bVlWbbZ
daCaFeH3pSu1OSPzXw3HWinxAgWefGuVqDkF88/4n9RmSUw63Yv34AE9NccgyCNA
J/qpaipWVeqwN2rvawCM2p6vS3TQuAmNoyB+fM+/bl5FeTRNp3rOJuKTq+rJFAor
8FYzDK/Q6VI2o6qFcepBBBq90t/mywzqG9/gafMvL864i/d+7YZWCLz71YytCdh1
Ga6mQh0/xQxwqi70cfnQx7cCj1aplc39YfoW1sqkwFraKDxz7kd28SfLcdYsVh0n
aLrjkTL0W+yPEInYez5+Y8gvb57vFeTrxjQkh3MNdq9j3LDyCCPLRunNTaYxCDgy
jSXSvBjrt8GDvXi0gYie6igONIoLWWgHpmJmtFwoaw4j+eOqZ8j7PuX2zcVRqIRA
1bqirxobVC1xK+ie3kCPSxmZMrGo8Mo3An83Fpht4lhZWdMAorCckPufBRXFZSbK
cvf4h4v9tLz06Oi23GZ7P/61LOuLE9qyVfuM4TS6snU+pjqgzyx232l0d3xnByXq
hfPcx9KSXVAhl1a6fR/ea/lnBxfZlxkEkKlOxvkXx97TIbrnEufxyZ5g7n9YVW6F
9aNuv8MfGCbNn43Md+tBWQrbe2tWWL4LmuAXuVh8MkntZKBzROuBmHvSNILak5F0
g/a5UJhZT8byooFCI/50mHCQP5PDfYPpCU4kjr49fwYdaVVF45Z/dzJ6kvQH4w7y
UwAJS39l+GoLM60R2lD1MHasSO1TErdyOD1B96wsjsNbmgnQxaZbAY87yXW8Iq9i
WQI0SmSLXvL2RMKoJG4pKTa1XoM+uTrXPgGG8Mp4VmXfwMSt6+bx7otbc33kFxKA
8PkQ7cnWMMmbBCuvZCKc5ODHf5kBogny63G6pW1A+2a0zT0AAvMJhYGof9wtd2hf
FFzMgj58HLne+NVtvarjkc7AaO82lrDLBsJk0PR7b/rHmanQbQU5XXoOvSIv7lJy
4Y+V6HBT8oceCAYntj6UgRf3U6/a4mUBeqCK/ePfbCkaJMc0o3US1KYWZJ+7e6tx
nasIoh1Fbg7g6tNp4MAq8/3CWgRalrjvKUkPjRzsuR6cYjn4uy8RRdgzHb21nokl
V8TVu62FJ7qbkc+mWJfZv3t5l1HKhojYUitA/zSj6CoV6pc+Oyu5z4CR5SVjK3yo
eONr3U9QSKcOh9NuK57s3LjXzBgAFgJAfc50he7b2xbRz/J2nyVGWQwa9ca/XZ5U
zCJoNKgUF3DmqhpVrLfckVQl/zJ6WIOlppdKceUvDs8azezv4pNxnNJZkucbQZup
3sl+LyyhxPAK+olMTmwAPsVsx9Nj6Aiz0CNPq2WBnMFJ44ruu3s1DFUHQexp+BEP
Gfkkg/+obfL3xPGrfS3EeK7sGM/8y/cg27YAIeIinqiDw7wtYsFq8+AkZ04zxru+
ifkzEJrL5TWDbrWUATuR6ELHwGNNygmmLSHWmWVLIrEHSg32G++AxbxmSTHBPEOV
rqRhuHpH4CjHaX4dssf5B1UfNfzroV9LfTUhMHMi3IN/mm+hBQbrhgSP+8MZRbbl
/xKpArxfX65FkcXPTW68os/zgtnnhhS24YZ75Kvb9A1vVznuE015mTHKhgmNXilm
TK39iuHRUtpU8L3ZU54LyXwMZNzrSBh4wlbbhxIRo5bgO74N5HvCoFB2RgT0wHh2
sf728zwg9GG655SebOdClDEhIvOV+XYitLWjgQL8MJbQxSGT9LxTrNdfJO1hXPY3
2nA9IE2y4LQeRU54zMEgJ2GEj6NQ/C+oEtp4XO8hSh8JhW+bZlzRxNaXTaVQJcHG
Syk9V2goAa/Hw4V59Jp9hXVOX+agU4s5ofBMqb7jRSfOtiwCSJNL/+nb+Upvroen
xpOkQqQ8BTZyD7LjFyUPOliJh59Wn8etZkIXiskj2S9sr9qGi43Au7URIFwpxInz
dejAK2xkiLD0duRQNZwW1NXf66r44k248Sy3n1QfiLADRAUGSYFSUMMg88eEP3jU
kCowAMHgz8G+M67fIV3Br1DQq1wyfRzLxtf6GCnLqHelEsOTXCm3y1I603/BDSQt
adm32oGPyCRo1eYSAZKdg+D90+MhpIk1aY/16vRSOICaoc+ftEjhBoEJH/mAAsIb
swNZ1o2rL4zpGccx107EhBJelt54wScYbjkPm2ftgwYTvbQ0BEsirAIoTc/TCq1x
gQQ6X3QAjmv6lzYrDTYpj/04H7DCzlaq7YfCU0Eou3VFDq7ILLyzD+wLHEUCnqKt
KkAmzRob3q+023WB1MwGXjepBdKy2KLNKCBp1m69QC7zsPK8XtGKfxDn4ShBbyyZ
UQkI72slJNZfhHY2isCTRbqTp9HH4oQeH4oo/dmLcubYkb3uzBoX1Qb8kpiv13SK
+7QwB/ITq0SsIl7kGYSUQ4lfyKLhVczc7Lyt1Ub6pBjOzoAM2UtTiuJurjoQe0li
/6C47iAeETWbM1HBSk8A8f3m6MoENTEQB5igbHQ+U+9X6dff5qJ8nayGsJpwIz6K
kzx0/rQZBbNmyzBWSddqNbw8jWMA9S7gTsmBn39FG7BBy5fUTd54Tt0oZ4Kew490
Hcuzh5NJZKHuDNiSj5dFHRK2iclk4WCBNDO94zQzlfB1kyG3eRDijWecM1Vu8oMN
G4bBImjP54uy0Ro3G0kBH1Ki42s8gLpMFTw/NuCH2n6hZ1Uf68q6RKauKil27/h3
nT7zAN+rng4DVvqMqXy9G5XfYLugFXCNz3XsBNWdkJZLJXpX7acl6yvDcX45BkP9
wkgIqnEkZvRfh3MmWwiOryut2oaP2m0ugQxmmrCkfBlk3Ov29hgFbSJovi3lJv31
syiNKbeybOfZ0I8oO0kU2p2G6PilyYjk9oVqGWM+s9BisJnyuxMgu8tz+CRX69sM
X9ebHHW6LCfOaX1CvOXaLbyXsiyDTWzxClbxL2j0ADwVrPcj8SPe81g9hPVed0wG
+xOOGUkrfAYmI3BxgbEt8G69CgTCr/y1qg1hUW8/Pkl1Z6nEEs3p2W03byDruyne
6alA1b9Voyo6fRzQjNoe2jdkeckRQt2nfbizy1RXzChAWEAyXWfpmVOkJZwLsK/+
B9TVSbRbP5RH6yOMIk+63friPqcPqsCrAYR1Y/dzSGQObBQcvVUb42sBUVgpwcwb
w6Xa/F5zLN/g9nwSD6Hj5lLZxfcgUVwWmDTqLxt7sZqDXHIXyioH/icEFvOl58ak
XQ7KNgwxKuZ6GlmVRbKK+lpKFcJFoE5RFnmZthT0UFAMTGwue46fXS5KkjIEBTDX
h9QWglhCSfdS0ASBHV2bVSMazhgpAOWt4Ax258Sb6RqshQgX7Oo8NaIgAfYNuf1l
z5SOxpZILEFzoUJdOT3zlhGr8M+I3kxUl6e59St5Ch+egtx4kcsYSGe0cZZac7jx
nBFRK1BNQWb5l6MX3G1xW0WpWZdnI9beQcltVcBRgfLNBGycUznG31b4v4cuILsf
K5QvBzALiHO5jSeIPQ/TW//6sD5N1ZL6ZhH647SJZOnFOk7LWbXrKGLYr5qzaLe4
g7Yd8fK/3tqAbbN4dN7dJFNIHbkEhtctmgf7UdfuFAoeeP1vJ/elEiPqq1QfS3IR
vLdXDu8uqY0g/ajqGxYZKlcNf5qrdbzxmMoLNP0cspVoiB3lYNCAJbC4ej5o/66r
z6PaYBkaiWT+aNOT3zmzOIEqFWfB/XejMK19XmmthVyMJvrirGVDehYndiSBMqez
urCfrzgopbXBRWL8l1tm6E8pT8WKG/le0HAvTVzkH85udn75tIC6aU2+1a84aRos
pQe5DuRcGAOYsRnW4niAeWE+iZFh7csjjVxpJm+niTAh5EMdvue3iCqz6Uko2a1Q
16F57cKn9/pMfaqhUHykogWU5gideNkTl7VhGMkwGkbNCvcQk9koNLChs+qZuGEQ
v26P/ee1h2GO3le6Bpi/k1f9naLtB6ACjinVaPwUz+vfvy69jK9ldaP7CK4zHy/+
wDyBlQYuUnjvJchos+iYyQKq3j76S73ptyOdhqVv+Q6vT4opio7XP/CEARxO9khH
o9H9RXi4Lx5c5b7nbKroEOejKEU2xKa09ZpnP49ZO9GrkLh9Z5Yji3NKf7BOAwYx
74J4aAZrv3J5tAI1XNSDJBfXOnBkCCV21RMbwZRt92K3Vpshe7CmJ0Sy+6z9VxKK
EcorWwWbedkoYX6NrkCS9EmYmKG/SkdWeNO2U2aOeuCTnOICOBkgWSjBF1WxhTd2
vSrp6d0GYu+2xL15Rs8kz44j3MYhi5ec+BMU9VtGBZ9Ry9BYIQwYZDYHtFWzrMaL
fjoGRjFOzpZPJfhlPfb/NLAAWQTY4Ie91hY3WuO0efV9q6Kn2NKsG42wS651BWxR
JXeGKyfBhX01kXWyxByrE2A9TBtRKKfZ2FzbVrj+NIvOhA/thuGPqzDgs0RToA2O
ffElLKKVpFXwJuEpc35flObFxlXU0bc85UukLr9Cru55MMr3cqCN1JVwHG2E6cio
ZUO2rsSRDQzorQQwdK9GRZIvN3jWDIHFaz/t5iBYsjoCBDKKHEF7igo1yW9yiILx
4uA+VzyhKgqS3S4TCM+7h4H2R2nFnd6d2Oe/Nws7ZGl6SRaFd6SEXjtnGve7o/wn
8vAe/i49gNbhEQ4SmPny3vQuZ9anwItzPIt7UzT73yqmmCWqQhlGFEWHmUVaeXtR
Qc3joy+2mhyCbonZeBos9N2wvk44+KHX20tWcHbxs3WziOpenGOueRGXJl3Aq1PI
cTorlJ5o3G7q4ZVQVmqQ8c/uaVPm6jXAV8CT7c2ajRH8jRqAQ0MlBHweYDgoJa3s
mJi4Nck4atUTGtXbkerLmC0idlzt79DvKB6IPczbmD4cmeWaWfJphQ4D/LG46+cB
1xLy8OETReh1KH/5ZzkCVa5VeqU0K06ZqjE+khQKVYs=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nLPM+OupiZIdJ46QaD292ew9LyzQ4eqvRAySMViSEIr0HzBPy2jz9syvkq1FlpBk
rcn9RAC8h/2ICPVgIudsUokzEQtnGASY2uuaFxNMkwGWWdfw9bRjvq/hRnPaKXbv
m/i3SkbBrc0luK9oYVX1GOxkB00GGZl4b0oOhR3DdciKGRQsmMVoHuGu00+JIWq0
jGt0u7AFo1JnNBOZiJspwHWUJZzW1nJfIZ1t3wafYZ8Q47+meiPzbGsS9cJragek
Vs3Rq0ZYjhvUMDjjGpm62YI6U1hcUmCtZHXbfdVuQ4NdGUSOCpI7Pgk8eig7dhYF
GRhboScHp23Txu8r7M1/Sw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3440 )
`pragma protect data_block
iEb7+fawM7MJKrUagdcmpqQOp7Uy4+KlMmuIHQzaFB8HZ1GbfQu5FQFBX55v7Zi6
A6Jx/OgCvdGuICUK9Qgu4Yr5ljzQ+T+G2OkI2md0n4qoHf9fcydf/C8oGMO4saib
9WehKYqWR8xQEiUly8UoTJ6Jd3M95kRmtzaMbQ4/Z0wJ4J5nSDsqUvl+x5Ntb/dR
egk9wsa/R+9NXzT/RHSAPd01KQZtV/6CWuNlrWAyL6iND2PTDnwYlLaXv0Kk4p8n
zn0I0SBGlLqgo1gFUFtJYSyhWM+IeT+LBbY2p1XcTzzpG5fmlhJHqJ70XcgpByLd
WeploBn59Q0QRh6qQvHYujzUDkmGIg6b7YBNPC749gP5MOhAi057JtEljIVoiAGt
5At20unVAiju/UKlkogPilrDFMw4W3KPrXYHXAV+cN4Ic1ONKsDT52pi9TdFF1Xs
f/22MrpB579g3vyfl8Xmy8PmdO9QErWgBidgFLOWfXO6ywcqYEwyX3bGGDgw9Evl
5XYHPq+uz3psf7wxkHgzIcvisxLuFRF3XQ7H4x5KxR5bvi/EQ/RH8OH9ErA/Ylsk
y2x9ccgCI/PiLBsqG+gs6iNja4Ym6xUpvzdPvSjte7iWeS2p+/BBSAyav3ORYUsN
RYKiL4cOeCUx/zkiesduBTX902Q38oZCzao/2uAfQfZ2wme2URA9rDfOStdBmam9
MZW31CI56AeUWIABf8tXdWmYe+51MA32Le+qkqJwb/49JL64+p4l70N9D5sRu7n+
2pBv/tc+EM0HgvoyoYtU/PKERr/8JlhrBeQwIwEGNZqdo2ZEEWAUjjtPfmf+PWRw
y5CA5eSJxn9avDdezj0hKkUSStWt9XfuCmBhtlXJSR/jNkNIPiZP5WLG9M9SINMT
oOVJco8mDnSKg+ROcRfe9jZiWVIlLKwDUz9JAHZyFuBMyFf5BCzf8Kjguv+83VU8
Gk4dYNSQT2kzfvS2o+I9TwUYqRDfpYiDgRnAHQexW5Y1jZkgp3bhZoB59vBmwgRI
IF9kJzrqCZSDxS8W7b81eyAXJtCunIDE1BqTPSkJ513BbEnU43HRr9XS93VAMpcN
4vQvYf+EB0jPxSfHmpJPNYhpQ3FW5R72G1evljCa6eUdXv72hFp/j8L4Md1m8AGW
TlaF/egJaYHWEhjrhXY5+Ud8feYt72+1RhYLzBcJZht/kTybImCOTP9bfqNZpXlP
2etTTzKGZ3RCwaQMTmdHdEkD9EronZZGIBjC6orE2Yo97kYVzzhwACMWj8Swjqma
ZUYNQogFCkcgmqqLmYjFhqbFuXpIS34kJX2Ng0BOAVoVH7x8MA2A6Nigd7JO5jrk
iV2r4lPn0aCvIlTcWXlVlXQQ4cUX9zIsEz+7DfnpDP1sPYM/Dhi6iRU8WG9/yYy3
WbSoWDoiNOcB0+bqI5kS/YeeLcXKEErhaXB8jO1GazLOGwRFj77CkeTi84iL3u23
kcwjcq9myG5AgBOFTH9g0teWY9MGn5YZlIvJ4f2+/XaxjL9GerG/DtH0AoGUKEFn
PIxUKjWqpRMTXuBiBOXOGa+Kuiixem6FrnBW4d8Hs6AWbiEaX5n8kK1j6LJh6quo
zZK+PDCMRP1wmLP0LuZGSKLrzujDMvjJOMex3FcivAX7/qUsSjQAMs7q1O1cayxx
e2PoreoPXX2gx+NqxHDKigsXFhtmfCiAWKQDM4ip4XTGKJsiGoPENyBLaG+WfF6H
25ecfQzbFaOUkNP+s4WtHsf+PnrUmsFvoSULAGcGKW53OFZVkra/ZLmjimf+ne+K
hjav4tLPbmSBFNumWWI0F7OCk5saaSiTyG9GcBjR+vZP2Xanwxx5rtbnfDlgm2/1
vx+X5ebUqA/ilJ67Vzb9ChdMaUFdO3Scy7RQm1RhB87h1FX+2SSPeZNwXCAAMo0y
RYp0q8PQ7jpATeDu6ZPcIIfnafizgyTDAuO/x0s+uLrOa5nNS1ojIk5SNNQqeOtu
gxYRjeiRnFw8F/vlNl+WJqaaj0vROTtXthnzvVjNLW1hXdDHK8t2s8d/33s5Q0uj
CgfVPCrpa9oIi7ib0m5tM9uKROpJR4IkyIPGkIu14vWH8pk5xUHbJmtGSTWKzarL
3Bj9zJAmfVPbannpHuJN25aFTNoS+oVqJEEVD8UZHH6rjAto1Y4kbLiXum+mjv4v
VL/s/mzwBgCizDUwta09+Jvo3LbnxfMiqq4n1wX1Y3G3xayvYHJayDDksjyHgIPD
cWWx6bvizfOjzlJ3rJHPeGUWYuj5SUfADi2EYIH2ociIBsce+uj75K9bvLVCtTMF
YpyIlReCYXkYQdsdsIrRq4ixMKcJfiBvlm8sQC6eH2dJsjV5U0kucr3lo1ZGwax2
Oy0ZNHvp7GQGiD41S6UkTmli+Y8tnyeNWSwHdDxLSadtf+bi159wdoipyMpGhjWD
/ethlLtzytvwZOYqygRw6ac+xuH+lU8jjioDzN2j4HlBgs15M+F8IDiwl4+GU/IF
T159Ly+za9V9s3+VCxmGkCUJoq00sdwsR5v7eq+3Rw9TdETQOAZqBWC4oG1/mXmv
UUv0r9VUQfMrUE4yhTEfC4FlLBrSQTLUxeRARExR47OlL157py6NXzss3f7MsPgs
WpaUPbbmxelKIX1xu5yAh7ACebNda1yEwEXfDUfiwv5OY1UoL3EgYMDHaPPWB15r
fq7tKNGRhD6ZJ+5zvpkcpZg8CG+aKzuDaA1nGTfA5JQc95jRf1Lr3/K9uMVX19aX
vrl5GVmPBYWN69lttXJPiwQXOuj7QYd1dRH4xiK4a0T2kJxTFRUC0/QBUwh69uZz
U2Bpl1nMuKe6g4/ReaBQTDWJdtN7ugoRXDXa5iTmtA1zygxoDNkUz+ayuAXdQhgY
7wJouyBRXCk4IOaKMxcUBuzBCl3rj1jmrvpLYyqqY9x1m2RMp0ArTAb/tIv9dh4w
XzBpehhit5lPUOErAy8TE36mILU5kZ4wTvK5192lItaEpWsAXh7PrqAKncKqyZZu
+qLwr+M+17VBhqxihwcKMMHnyDOY1cmHNxPfS48786ryPc2lqPlnkskRNeWnqDjw
0/Z0/H66cxu+gTp2N9BCEnrvR0cAeRXNWy4nu+7uyWgI4mNfZKO+kU6Owwy5evzh
BtnZ5UDbgcrxioVC8+9IMx5Z3PBkHIraYnjs7IsPfIT6OZS/V0lTNqS+WGmM+h7L
N9I4zcrJQhfDuTWaD80ppKCq2ojewMHKal0mKpHWCKk5lXV5Ku7HwcI+UOKK7whq
+DyBazz55wIHhledV4p+vbYwFNZLTaBqnUgdfhL9bz4rylUGZkeJ/3zL1FSRKLNx
WsKrfGXZs1s5q7MTUuNUPN/OUjHiQGNpdEbgCIfWAOY6NkmLXf9VbPFv2CyGpU9q
bn5PkTYb9u4FpvyQNefC8rLQIs5IZHFpFpdPg1ofmzkVCzjvOusQ57Cy33AHiItq
RbfhXqAtH/0O5ihhlH1GVCiki5cZl71q0o4iGtoIC+GJybR9PbZ9RBuHM8PodiO+
C1lHQV0YohBvjz6Ng/qwZvwMut1t+8cL4/pYSx5/Y6iP9oo0a1iNs23wAA0JJZhA
JLrYNVVaiDcNm7/j9+REnDxDyzYsGxCOn1Nex64DW5CxoIvg0u2cec23zHziIPSS
DZUOmZ38qjFA2L+cR8oCfmzGK64Ix+sHvJ1FJm/1X1xchKUMK39nb+63rR5NVL7Y
OhABaOv5crUAmtMgSN4+mjD2V0qBeXsda9v+s3iIDVoLJ20wg3m1CnMKrJwY3GIm
X5bHx8sWYB6Zrqo+nbzgFkdKN5f6H/w2Ut8sk0qXE09508zgOwtTLuIM/XBOoArO
wTgZ/Qx7f2ndHs2kTekE9ZLWXZWremAJsPTrjEEzeyzTQEZ7OWX/7BYT8fD191dj
hELfaX9MMvI3AoYdutyTr8tqgMa1rDc0IUXtSe2ygxsl2E82MlaguszLfRm8nmog
yYMeAs850J8QI/xtuSGNeLZ2XDXiEZEHQ9KOXA1mB+6bPsVTnu7PVYPs83rAd/cz
cIRLklnOAJVC+ZpXxjW6dK2i8C/QST8OM5gA7MqCw9lI5PfdxVIq7U5T8wluhIQL
K2RrlCOtHsUM2oigC/lR4U0KLoGH/cUkjR9S8esA96u9Pb1FJv3G+N9AlpP0qP0M
9gpKH2AmAamlhgeBpo+lWFX2HsCbWl9GIR7b5bFedIacNdLsTRN8ZAXUxsSD39ad
n8u27CcKIbPKinWhjmIqYgNr821HP7BuYS5U7vgjXMV8OCW8sZ2hBB2SMKGozs1G
gyEcrBAAq9aupPadlDGF7x7UsUzLvAKdgpd0YxbzL1d4O5Uvsi2i9yZJCnKtstnl
6HoplAFaYxAb67j1ZcSrhJqiGDVulco3tWnIJaAY4bwnbrh5dwHKSpj6TzI54dUV
2AMBT/gVtGvJodpY6y4lXgbTv0t/aDcskvkQzJRaLrHIYssepJq/OZNatGS78jZo
EfS3WUEPi7OAufIVqWaSfi3ZxTuUBLxCawWS3+r0sKQ39bzNZZOgGknd2oE/gmM1
AiK0mJ5rb3sKGAM0cKhEr+vaspSmb1BHqqRFpxbapqs=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gJPFuEjC49yK4TRNAnwn4ezYcGci02h6ss2q4uKaHwSX8gTUCsGvB9zb3nJukVCa
motjP0M0b4TvwdbecY+V/Tk9EYPnUr/jxU4NUQP89bdLZ2zABnHtpVhQlkU9p5Rv
+cUiH8L5kO1/b311rGyh9DGf+GCTNfe5BQEeJEFUc/eDnkPorwuz5gOSSYbOvpAN
FP81ux7fpHmeKqrgMq51L7XF+sC6VAgQUIVuXr19oKcw5kEMvKFdUmy1WfY/2KyH
mPSn6hmw9z+SiHRxyeFJtH/gQPeN7Zc9PHUQUSfCxU0tyQBS1pOOol9YJ6WyyyMi
G/dyhCvUSHCjZoKUgYhhmQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2176 )
`pragma protect data_block
t/wSALKZTn/5Ji08MYIxKdlJtdsUoofPdtrlCfMCFh9X1ZduAO3M5dHuBqE3f3Xv
QpnHh3qV7Ahu1x36lLNyrbReNdTDKqtvt5Zo2n1mutviC/Qwi10OqE6Yo4sFBkt1
juydFsIMV5z3blLgLdseXLgKvr6akOpB6XbfEMtoo1zaN8BsqeNRegu6z56cXtrc
tnSHUphfjqBxTfxp1jWQGgdFcAwgxmDmNARDYP8TzL0C8/QbXr9RVa6z3kuUOcaV
6qJr7Yn2d+oAEGMGygYaA/hdMEh4MovUeyZ8Rgp68frrbPnLY4pqmh2hLZ0w+J1I
sbMZ2c+DIF3WWTFgKoeEvouenUlSW3uc+rgFKlkapUZ2plZtq+m+6CSZbnwXluL9
42V1+mrOIGZw9i4HIIbMDoKYc2eMflFgbFjRZSde+g1OCwBNrxPkgjlH/Dn13yM4
ggZtE+6HIc+/tSOwoJ0CFKiVzRMMioKnUY04ec2Q0kJi5KnfcRXy3n1MrtacEDYR
HcCU5VQFQ8AFd2igOulvgve8mXr5Sl3LQ/nd4pCWtOdvFmCQJuQ2Zu5wEWj47QSM
DIKJxJ4rXOM+9P5XBNa6g9Zod79QOqFaIrV/YjQgXh+bMa5JYQ//DNg4StQMxZy5
fRqTD1TOBH+H1Cz3XGFdlt5jjFDfoPAr/oON28MVfmXpYEsez8TnHEo/2FMC11Al
xrvZNimME8X4bfmHj9loZgfVI4FO2wLr+3pNZZ5lD+Y3p+o+kvukqIduj4jfyIC2
GG5C4OV21WiI1fn1+BHTqDKOY26m034Hu4qsw2FTf0KO8mnuxcdHXx2wnKRikGnZ
99AsKmB1Cgi8PoSzKsQuU1XSzRuNt8oE2ExPCERHqOASqJTWzKkj3wMU1jhuAkvK
zYy6llrQWcJbv/Lb60plYHP6mzhQBY6j31xTSGXbhvIi/PbbERV7IJtPXl3BHZzj
P9JPmaVh69vrMjcm1B1zoAuC6IRW12gyyIjEnDlZeUEss22h2TqoFi+4tz+a+Nqb
z0ltZLewAn+7MFT3yNYiuSTtooyblSKJPNCZnfbB6REMtgl4lB0k3e+50GSg5Ggv
wL3E7EptKv3VZeTEvr/cwsfEwqcgCjN6ChMwNfWjUYnGqXFcjw/+HXmlinGGA4ks
yW56hJYjzlHWcUtD+D9amIUNDD93qHFGEQQL3+20Ev8Oy2tVCGMp9vCbxkIfV0MN
SFJ+6Jtwrg1iVpROW0A/EBtJqKuYbt6na10CNdThT+grddRvYeM6+xMnHS4KGMYT
5luxzfwIKPZrfwUp2gGNyn6RJofm1CM30bLmoznxLQVF9ubi/Kdz7Uh1/0ZuiDNT
Mz5sEZtxrOs/p2oH8zxYSAtuim5A7q8j0Fx3eouWL6xfLbyfO9Fct3FU6U4Vnn+i
97uzncSB0Uu2IWd3bdzPh+VTMMa7lorO9L5ii2VizMo7mTrsGRxa0VA2zzaozx59
ZCL1v0nziQwqm3t25xayIWQqy6JFqIiZ00CEL6l/6+Bh/vgyqIqwTfTzxeKRAqNE
yCCpBBK9he/csoEFpwc3PsdvaKP0QzQTNoqLDRMyXD7IJt+zPtGh9XZp/9RSJaDF
rZKDRTKaohb15yySTocvuS9UZxKYk59CT+quWqDn5rm2dVtMyDJkTvZD99IX44MY
DIbIyQ+OmpC+PcfaX5TJtD21JFeF1z6+B5N2M4xFroW2jNkpcKhUt3w1zmi7t5SA
4Ll42aVrcgcDL9jmnRnHsLhYXDk7xvNGt8AM8A+TOWQW0SsBeep/bD2+UvVvjwzz
GJg3wFbxIS18fz8sYdBOGcqcm4OZ0nQn18Jowzv10M2f70TEP4y+XBTtdMkpOKQl
EKVhIHWyRwkazXlHAOUWRBh/xp7+mPJ2W9QubEXMEtKFSmsZGKFAPuIprOU5cbp/
bkndqizhiu9rWjZsJJ4jpCxRiniJixCi1iljLPL/ei8lUPwbNUSFeIhRQ+ZgYrXE
bJEmjl/WOtCCCgWJiWBn52Q0EYv3zGrXVENGkNPJtaPLr5XnkP8MMJ1tdFYonz0D
Bf5xmEyc/YPeBu7XWkzYnEHo9b3V7neQ8HY0LMjejSRDtmqEWSmMzoE+jDlcgvHW
qqOWgvo4BtqcEJBKoJMPuSCUcXGGOTmhWb+Q/PqUf8PGITj1koxvIDcqMBkBmwOG
df1IaX0S19GQaVBTGo1f6dv88sD5uhfi45nL7aXVgCnZrUGs51sjWzG0vXuwwJX2
H34NBxTG5vpQ0jRE6rYuaHUuGNSyr4pHFbxHxFZe/ixZoI3oC0cBMmnTJi4zKUcD
AXddFtL53elODyZYcQgGHGMHmXOSRplCei24Of5hGDBaIri6010D9UOv2BlcE3PS
0lHWAx80zLtq/lACvLG412TDzd/Ssk1KX1RUuhzzZBfZiXWyOb1AcPV+GQsHpNq3
lV7f9L13h3AYWXzH+z1EOU7uZRjG6my/QZbNdDhrqSC33kchdvJzfZ3EcpE/SApU
Lojy3UUziwsKkZnVLqh0RprdjI7uTte+3dAeRKwS8IKzs/w6IyrHzEClk0QeulzK
TLeK5P5lgmvFriPaycstsdKzM3PvN6vJiRnmfvkoY850wNggaSDGs1pgZwdvmlbd
/PgrT92cCLPKA3URmhbxOUY9QN9POdggW0cZdhPtRvHZoN89Be5VJSeNykTNPm/V
EIOAakTeKj+Eb0z8q8NBqRDf06X3aPGPFI0rVkMwhq64ZVwJo8XGk+Zmn8gGK8BZ
v+AoWZlsGfj9roijXSORnqY+os3ZAa6WSqJ1nQCUd705pLqOVZarknabsUIxoJvl
ktcnwiCPN1oFVOtm2CEXA8cYMyIPp9tXQHSuMPH1AS84Gb45UQdRUvTPxSMPdk0s
c+6pUxMcFpBu0Ihx4hec6Q==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LDyrmDWrOz2K2vjnIvTVsmasrGBWkxXWeUKgVfiNroerkuzUff4H/7Kx2UjcwUGY
gnwzfV/fsx4zw6HW25Q3pwV/uczXpuGF/g3M/hjXBqSeubn8GeEm81zygwXFUcFF
Dkden256obtv4T+K0svElXkGC/wuvpRdQL3+S8Og3hOJOgsKcApgEStr0ySlLkt8
dX86xAaLv24kN33P0G++oDY7QiUP4l1XB0eB21s4mM0UMObxCM4TdS1p9DvmF+6w
41T8oMOvKBNE0Le/ZVv4ZprR9YHPKJ/r1m3poRHArTATE6Ba6r9/C6vGIpEWoq0B
uWU8dI8GKMEqL655bmm7gg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7072 )
`pragma protect data_block
aahQOxCz3uPOcceGd+WsLKVyaKC+7cqQFAjki41JaXe0Asx16UY6Z65zcx6i7Kli
0PltHsB0+3XILY0DnmPI3tlT0zbpzRZZMJrWMY3Njsj88MHRiSN2/Gc6jWopIRHJ
/+5nsEuOxtHva6A0HLY77jywOAueAasfNUvutOKyu/cV/K9QqfAppFLJXh2HS6RH
HI2YBOtMgqHwkL2AwpGjnyv5NkgjU0P6G2BJSi22GyK3fyOa5dfakGBiS0yeR2uT
OSyrWKB92uDWcWAmrFq4LQxvv+0ewZrE9445inasg6kIGpc8K49/d93MTQZ3TJz0
YHpU2bFS47d5EkKOyUy2xDI9ZEa+LWByltOMvQOuCiIdvCj1u0LF46oVCwB9TRdj
rpBZdP2WGmE16pEGmpsH8nipVUCY0n0gcVFUtC3CKpa1Dfh3fp7xCndHlPaQITKM
FqOKoI7fxezlK8WfTm3D0rTQ0ch4fr/yuMEwXTor98d+qWB+aswsXu6as8clOt+/
kJO0WrAAd6nhu/lbICgPrtgrnigTymnLnulZV5DSx3Ysu8Jnoz6aW33yWOXp/9SG
I0MEwcPW+3eGbgxXdNSYpy5PW8Z+jUMwCPg0bTR7WkbMvRUBATrY3N2RgfVrXUYB
xOuAzNSoWPajUEttKrL2JWVtx4Q+rkpz3V3sXmpOGjhg6uhgIClUSd6RYfqC4pli
qIN8aAw7G/GV/4N5XO3nxsrQi9aaK0S2FEfq3/LBYmmO6M4pQwSwpgttrN9rXIzW
ChAo67DxFugYnFm9d8ceErb14Z2ThsNigIfXEQOAgSSxhzUKSCWGIDKxWO8mQfrH
mDuoW34SxgcRuJUVEZgCh/q0R2nkEB4DDHn4fNddSK90wOuiEtIUgNTM7Ptt7fhK
J79u8NDoQUICcj0Z6SAqektORcIRCyWqzKDUf+ad94ulr2uk1twIN7cmd1y/3RFj
gx0ZdHxzT0U2sRwyTjIl+2cZRSpI8qI9k7J+nGXPwVVyvByy0o9UDbqZ2GTqNlNK
nuOOkJPSIRW/eeq+5JkIbGJrIQcIayiJcNvzFe8xybbfiqAoC0ITagODDVq+8MDY
/tCWym67NkCtlPQmOvCjgaeBcuptS+4lqaLQkpmOscelrS/76t4rI9RWvCCfQ6af
qIE3JePoIvLIU9bpirg3zTXYWikpqeFd/smLXbbVARRK9yF7Ky8oIYwRLWUPWOND
NTZfqMfBshmNCDSSMUoEOzdvHe1kqR/WdU2v57+WSGUkYiTY035viyq0ZwTb9KJ3
uYsS8hbcXO2eF+e2w2QrsFXMNYWUU2wNeENtT6J9+Kp0tMkO4/h0PZfyksxZOFcf
Yrrj4wTspr0xP5R4HZ9O9pyo+aLAEKejieHuWcBqzmyFjSV0Arm8W+rgOGMiep43
t7HA+cRtBSdubZk8S71Wm2ZAxGdH27xZfHX+0qsdDHurRJ0hEaFZ09RGsr5bXIOb
SArhIU+M5SkfwoGG6qh7k3lfKV0r5Y5LBbkxiE4TmWw4y83bH+y8g3S5uLiHytuN
mX02Nsj0Szu7/h67/2sdl/vcvDLsdLJtwzfYsH/Oqic4tmTwKvFqokRC3yMJ54u6
E0PAysCMXDFrYv/0o1sNjcLvmChynWN5tsA3IhvkdzT8XMlHeOSnvh/OVCip/6eW
0Pd/Gu704B9JIV/oupPyqelSa13O5iFSTrUrWNMnd4KT8Z8hxWzL+rz4skFp0Rft
D8UzfBHOkgSwXL+oIqD2AoY5wTHnEHCGLbolKdVMsIyYNJJ6ay5WpREsRILJ+TJG
i13TLXo3j616lNlxBIPxjuoCusnB1sYAhBhHJoKm8APCOwZR9DDYibQ2PdFHl/ba
r5qfOO7cEUhIh94Kb0H/c9wMHgAyYpBNNpIAtoj08dCcnaQc+0fn+VwYQM6mBXnP
qz9GcgDDgsce0xafLWITdCZSD59d+pP14cdd6qaPOVWT4cTf2PYpbzbQWzQFFnh+
1xowjMdX9WdD7WJdy+jlL1B4UwVpwVbPQDz/LCF/bkVibINd1+J7QS4ZJsMrW/oJ
WJzyN8tyV5DSFkW8Tduv4GEGbwrFdjjQ/e5dpnEQEfdroPh+PYYbgyjfSFO7QUgH
MF24vZxH0MWb1popgY4pmcWkUR9mjAIIWHSEKMBGqVzav6pUrm1aWJjRpw1Li5aN
LFj8ivCqO07a8I54DvflWVxp6hblnweDBwvpJlLA1Ys+jJeuaCOfSEwZBVxZjVxF
byJwAiPj/6fZ4dUl2HcurhD5rBnqB7Vmw7GLjxP3/dpHBzokWKp5/DZSI+c1jstT
maYBXnH7AScxJwO1fwRN8aXCIxoApXqH7DZudQ3iam+zoO9jDkaCsBrQyAhIAdhC
dSXEGfOEAtI0AZphWP0fgtknT1iJyoGXZAnYR5egF6omInaV7UF/Y+4RUF+95YkG
bvmKz+pqH3Rk2tUICCu0Lfx0X6iV66FyryNqsUBmuXDq1NKi5pzqQwQjVbzuntQt
U9zqEV33hDAsNlshFyJAYyy1Z+9Y5nv38wS/Azb4Jd3YAK8Dlj9UJfHixL1NzSdZ
A1j/R7VQztFe95SdBhIpxx1+plTPvziXTugloYuXcTddg4W7duLtcVzdt33HYtwM
GHHZ54aM34ALo99hbrjb+GT5g38Ls1JHATOXiHYUyQ/yHGIjBzvcfRgtvV8d40zg
Il9STo/+bA8FulFaIQTAaiHfGJVZo7TNCF/Cd5anQjC5PN10gLVB2Js5ePzvJT/I
zn3gnOI89GDVPMDNZy0q3JY4xJ5iS3s/nTFrmGWKkrbaoqGBya02nmCgyNimDW0E
v1mBs4ttAtEZp/A5RlGAmjEtuAXmAxFWCQpbOo+l9VezT4qZNo25mgzxMZk5AU3w
3Twh5EO/Rj8ni9vi3E0j7ZvmFGbWcix5BUolSUddka5gSmdxQF14rv8wUcQLUqX4
kuk86x430AC+9DGMhlSqInQhPZsbGvGCLVq28jaNZlbiB6tdnyJqsckGqhuxresm
4LgD0MfcLePQ7wsm/TjiqFM/0pzRmWrvLy8Q/m4rRxTL+jJM+UZpzzN+wDiaKvZN
7kHFKeXBoVXA4IJihN10PIkQ2CAd320cU2lirc98FsSDznajUjo8b2zY+BVKhFN1
s7tgXGxjPHDyJlajoFPOw8gxV7xjPsagDaX46RuJ62+JXCQrB2rIR0T/uNB8E5IJ
hX3lZ7uHwX1ynCJ+g5hB+/kGIxNRBK7yYx9u7/rC0aRsschImSSDKzWm+OvlMrap
nxfkf9mGpl7nK4Cf5OAAlmPbvBKXUqOJJe1BKzMot5lzxhTqDRT2Z8xEmjPCyVjw
gBaW9/krARLBtm5rYcq9kf+5E0lf7KlJXlYyabnbAts7OWx2LR3IhxCyzqTM/z8r
segmSx/mVTBZy7ngmSj6re3JSxp++CzObhXukbn0zsw+ypAaVe2DL8QIXxwTiFrd
iT8o2NPUyvoQX9N0VbZvSrjj3qbarqpAwoh7+sVttwlvjNXkEbIyD8aFDr+bF2tO
mwk9ATHr4GyB4d1ercGpt8YL87vKIYKVhUPPauu/pSFQIlwUAA8zfSFv4/OkKe1f
NsVfMIxSvaMeKesOC5bxKGbS78vcwsY23n+QwjtZEO9RtIT5OejKX8p8OMIEpdtr
XpCBmoRg57Aj0crdmAqoDTorAB45Sc3jsy9LYYxhq/EdQPucVYG3ojKDTdW5h6gm
rR2qYepXW9Qh+cXxRFnORvooZaBJTb3aW1DYMNv/vT2WojYlwHv1awmHyVVR3ONE
fme1Mmjd8wQ5GatXEyHGg4ev3vOUAZTHs/lWo3+hZfFi21VvnaK64sDv3Q/qyp3d
KVExX9r3PMmqO9s8nAtU6FSmW0lwwscCJKJ5Fsu38s3STCryjkFdQLFViMAkjou8
U+kCyxYd6aMnP7udNMehC5Heivv3vRd8SRjWWpUEtx6Y5Ywv8VqwHtbVHQF7k4Kw
/8cLb+5IrErxGnzAI17UJD712cjwajEMoY5PDdkfaz4mm4um0X/yx2VGeXuEMkEL
3KyNsN9sJYsy0QhqiSsqsbJHRvsxpN3XE2JYVZVniu7QwEcnSfdkT+e/xW6p8og8
B3MV0PNAkkSgg+P01yxE6LdGchQCwagIpzYIzJPCapHta9UY1SV8ulX/C2pkerXt
jgd9Jery7ekK8oezDelQ7fseAlUIM6neNqSJFTRkrCujgJ5eMbN+LE+ynC4zS773
cEWRWgJ3FNqsfv9oA4O2f5SpVNv2ff6yLfJp9qPGxjFJ13S3eM8GI6tBttiClA/j
5u+eFx68QWoAOl9hAxA+o+ZyJ74H7q+Z++3oL4+IQ85V+8dU85UqzfUTWIvGiibl
6hz1mAXMuzbxorqYwqcVK4io334Xzq/W73sOg1H4LzInr2Dyvv6RA7V/K5DrRJlo
8scE9Pl9G5XtxWN1CnYwc3lVcIYoVktwOb03l94qChPloRqrGUiLwFsm1woFTa5R
uNwa49Xrm7SVWp8SSy+6sigoSEuL88aujJB2tWIdDdFss8N+eGq58zfr1urOmwrI
hsHvdpMd3eyYKBvjTidfIqLeSqSRmJ3E6LbkiLtUe68Om0l9hDtqpKCjQPQjZfAK
XLg1UTSppxs2ROyna3/zRhNHdCZmxNvL5Ej3JJZ4XO+8Q21g0R659AKBtfqnKuTJ
kMKVM+Zel3+usOeYbf4/Ugy08sE8iRZYQc5un66H3Zdf+8e/Opf6tQDR61rpBKy4
tqcV89sUF+IHMDUNdkhZCVA0r32h6UK+9fr0YPY0Fsby1nUb7epa1YuN0b7FTKOF
/RNhX964C3oYFJ9e2yhg6cai6wSBEO1lR8LcV0qRa0V3Deodb21pDBhJrG74PAnh
KCd3qPBueby5H0UedkBr79KWq3wmiWujXatakSzWT7F9jKPg/rrgFYFBRyoYRtXN
PBfJPnOSsKernLXaJuBC8BQ1PZIBC5O5bISyl012EE3kC9aYUbUb1+juhkNgf8Y8
0QUid38TKMytpRtkdCVxY56XF7BcwekX0WMWeV6OB3umVfiTWrlHspk1RrWW6DCz
E2ogAIX6P1I5Gr+V4rTbiS4GXHjTMigLp41CVlVLzIGVrpcUfJQjAfX8vilGTl73
KFTOlpOAn86/IJV0CD+DmUEUiyamWMfXWqIPpRIspLTHyEvGyAVp+e5U7gtBOMLf
IctEPsEC9whI2lZP1EIUmuSkRJkk0fcVPluFIrtDXoN0oQ8L9NCwM4idslyZUAC2
bxoXrenCrOxh+w8IKwn29x2CP+XjU1k4e1/87TgudmNEKC7HbDGsYckUD9H6zAX0
e496qGBdZKaAmJVMAr9qTYeLKZKaXW7GfezvgXDnhxnKNGt8ukIAcQgfjknr4YEj
KNUB3Y0A7unt0y0rjOdK5Y0TVV54lLOdv1XK8HAWYcLbBi+SEkTsfQ3XgO4TY/jM
RRIBW2h1jmQNN85ivx69dRvlAPyvzHpBpVvCCvy/eH9PAQA2ODCzSTXvoW/BFuNn
iou8pU+GhQyDogHlZ16g1FL8CtKrl55A0ypam1U5+JX0rniyB11iZ0RdRKDYdN0D
FckHjEd0PTHwBNWluu6pv33CpqtnEXgYUZpl15UGm1LE8X6sxX3OxyR1mlUavcg9
34pKIVe1hX0LtuboD0g81I3z1NeCun+iqtq+XxePNz63GLGORwEHyiZr3DqA4bpf
sS1qjUlb7X+kl8bdPjB5xHbl6558oHuBgui8NJHRyDwJbqJQO1G4Rfz71PLZ3uzb
OkcI0KFUUUZEpoeP1Fxs49r1VDCG/CCwnDAd08XQbgCdzYGvJY4M9eRJ0VtHKs/Y
qv5nHiHGe6TfVkaIejkNS1a8Z2TW/wT4KI/f6TJcRP0OIONHiAzCXQIxe8H0IaPZ
c6Mh40nqjrRLE7hieyeMpX+LngZJJzYGAp3WdzkiN7lsxIGlUxFHpxEmkhqBurQw
VcmedUoK2ru3a7rmt5HcCB29eRdMdS79VwrSZLU1dF6k6d13mJBmdnyc7Tx7vjcQ
XBIK2cOw4u7yx8gqyKrJlHcKT9Rd2hOCgpuyutTP2hsGxjCrYVoQphpS0v9X/GVY
vNTq7YWEmlVYHmgkzqgIOb0Amw37GYcotV8TKg5+kRj3gQQcOtCfzYt9/chXQ0cE
IdqjTE2WSjIf6DNUddGZw4xVuKIEq9NtvJN6HlWGXNF6BhZHLCh39CfDVq+cPw51
iKzZOVYhbBgMxSevvFIZxrdflUAT3u+jEddPU+RdB9gT9fvti9e6ecvo9e5RmAYd
VemcWonGhs9R3yCgCKZAb79EK9RsBzZNqUqCDr1Z3hAW6YC9ivh0XJFPpdp75ySj
0nmvl1DLedCNxGU9fxj6ruUmcnlbbH3qjRDLXI6Oxjo9zHs7hgHipTCVo4R2ekSM
QDOjrAQzVr9LH2lXtxgqCaxhGwBcKMKPQa6KQZfPeglkkJO9pVreOs0Y2Lye3/dm
B0CMI95VY7KOZ527mKiIT0x6dykasAMm62vSjoySXfFCQQVqRmGmcAH/xhcnCVh4
+sC2j8DwjGpezWUe1/1VIpdthHLG25u4JHn5wrRYMVIpag0uaXXrkh4SH8mbF4k2
6Ia56NbLoarmKJWC+bJZRwIEfulUYvnhhuiF8B2eCTi3K/xvIGh7asV/NuuyfIHp
vfizwnkfgmphqxtTR6PJ9CU+o9d14Stq2fCl0oP5x7KvbJg6RpujQNmQQFiV8mpr
/D7NE/NrkvF6tD9D7usD4LGOE7s6NbJCgw7Jyme8v87vLsioB0lvoGApwy/oQ0Tb
zDSWIsnuQUdyTWx9svZii6xZi3EoC6BCFPZ9GZMZ4gYUa80CMpsTpvARZ3z/F4Hc
hiMr+3mgCMUUmvEsO3VRD+JrGj2STWwq9keFqmr8xwkYbO5WwqP2pzz/yiK/I3ih
Kbu7FUwxo2GE3C6sqpx8PRB6TfsLdM7GvXZq5lZCuV+LOGl3Pet1VAnUoxmne5GI
DvorZ5aXLYW0zhkR+DjxdWVXXdLT53WR/sG4mrN8aFT+C+LmLqaTNUYbLGS7yNiI
aLPedPLBPiS19CKDu63hH7ILGESDQrPEZuGJ1TNDuzxFCZxkRSj505yYt98MyAh9
KXczFfIdXYpveAlBdNJbDReXYBQuZz2FwEuiCcDqHS46ckyu9r/Zalc3dgIdEaJI
BmX14rf0m+PxLc706qWeT8G5jdGb8wmeKA3eDPbuwpyMkBgJQF9Ul9GbJQkIvDSZ
fTrKmrx+58rZKCoQnXxitm2nthIyRd8N9tu7YWXgbBSKhj0UdBR0V4J6GRXxWfvE
lP93oTxrT3VH/wRWvfdJb0S4quZRHgIqCnHlkgkOOs8ayBc6LrfGV1UDIaxuUiSl
cuzVNbvzF9lArkIyyxlwZ2RQv1uZ32ziw4RxhbeeDlG1O3Aw7RkibfCtWHhcLGzn
RKuQF66bV9bp8Eht6t4VRFqWUS4Kd8FNUr1aHZ++X5nUhg370ZuAIe4kMnHAhXc2
7hSLUKbx1EDhiC4k/93HU5ECmxsRn+pOH0tf6+NDC/tKUSqxHyl3V2nQaxTBTJL0
nHZl2MbBXFyWU4Yvb7kVDkPbMGOPcYyM9XJeYMlqcFUqhoYByGr8AXgBTrn3ltKr
nzRIixnoqJr3SMHeqfXTq7vCbENGlTDngpgz3KxU0l2VAGlzHFuBns+FziIUgdrj
Et6pn8F2mlOokbRdnEn/yBIkUb4db0DDWJB8dUk5yezwxPjsNWICItca43DsxgwK
XqB8Uu0VhuvbAF4pwSlB2mi6Sbl9mEO0diMrajTgLZIclAxFcaXdUYEJOThbypkP
Ar6a0nwYpvRAmqbcGcyi6+DNiWku4hQfKri9EZ8WDEjF0ztpARODIu8xTeisU6Dt
6drN8yykwA/c+B0uPclRL+kYqjCOiw7pvovBP3CH0MF+COERHN+yS/fJk75MOXHD
b5LcnvgLdBGX8puoXVXggzWM2/jwPWczW3EaZgtP/TWSjQJoCDdP75FgN7ZHfDHh
NyzaawbkLBGvy77jh5Euvq5kWmD6+slvt0/dRki8O9GQosNDbW4V8OVKsKsK7kIZ
TO8LEktpHwqiOUar96+JXIzT6+T1mbe6kKm0WRT3eg1tnfUkuiBlL245GywMDFfw
MfUheMLgVK0VcdU0LRvTYZo0SgBI9b96HNrue/yE1B5jBtxfPsw0u+jG9Rjx5F/a
sq3aj55PXnGFJ/egc7846HfBpBZWjEuQTGsIxrzoQNoCiXbtE9dMXaNzG7v6r+No
+G0+oQhU38m46GasodHg9UH/UGBV/ThSAfdYObIIBsROpSvZY8/BvSjF6DJ7nCOD
1m7gcTVSOwHPic4kn+1e2Mwg2AU9G3DF3788/C4GVE1rS4P23qijbnMf4RdHFboR
0jUbOVSPV7JXp/gULq4ywVJ+j4+uFfIm6EmEH/20VOMOM73lgjnDXtYeBLk/OBy9
6rffYFTjwKeUDNKkoGw9xzyBVychsYxsXLgA0R8KV3+4b4Pe2CzOwvzB9sU9Ohxi
WT7fJbBtZ7MiTAXYX+gIPSBlL3HeK6+4E9Tqifqk2ULAeRnybFDZYp95ZTCpSV0X
v4G6F26yjiKifF2J/6SViYYtFHNSBF6oqDcgtUkVMna0w7YDkBXR7ZiO87bcHJF+
v4ymxwtD2JU0B2uNxuUlmOT+jQMk7eSlCGl6vpRArvZ33yqhlURXjUmCDtKbFKKw
TEi8+saC/GRU2UgegS2/wLtk2xMkBVNlGtfa0Jidpa/gQalxoh8pzRtPVmiApz5L
IktNBEh55QW5JXrcPPJviP6XRu0cxfCwMYV88tXujCY+R5Ea8cp7Z0NgnEgxI8aB
nTrmKnqJWjCbGM4jvoK6ZdhD+vWaDCKcNuUW9DSyL6RiTRyfs0gTiXrjGCC1flb5
LjOQbTOltWWpOfi2a3++zrCCWxQmu+MrJI3QkkMQMcqV0c8R9YJp5QBFUl9xK4A5
k1EiAcby/bR3tlBw0CARJZWq/6LkuTOP3nJalA6I0dFeAI4JieQ1Faj+TSElSIPd
12u7SI5bxlUcm+ddk5bd+xKEg9eNc2RBTmugLi+0IvIlQ9st/EFE/J2Pi/QfmNu1
JpOS1HHdZ5qUlDznDNJvPlvJtd0QXbLxZ7J59d7aHo9E0K2SUWZzZbnTBhT221vR
CMloaFuQ0QWGzIQ9JZUyX1BJeiqxCvpgUUplfzIwtnipyDlgqcxl1Y1/8nY0NS1/
9a65UTTUT/B9ZPCSmfbQUwb7qKTJV0EHtpamOJ1tRzGEQ0XS5ot0IRfe1iHtKY5t
yLm+4HlhzRu3gNBCiXx+a+Htfg+0nld8LhQVrTljz2wItT7XNCJauZlEYVSZlyqT
Ye1uLJMcUFM65P/DQw+zLHlDgX9PsFxg/NNUx3rxvBK985Hm57bVQkb2qjVKMuqH
NMtpDai0ny56KjmV0u7wbw==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nxgK7bm/YEXvikBhEURmGOFyi+6aFFDnoZ66YW8d1XBqQyHzqu0T1TIqFyJk5Gbr
ciVsXDM3MzTd9htYlPeTI2iXBYQu5y0pc6PUHLf4TcVhZjtbzP9IbUnYjF0zn946
xyIZ6KjAkZ5KUS1BYCrea+g04LcE77UcOaE4ImynwU7FGWGlNjcsZ4hAHLru9uQh
a+CJNrMdNnHEfWh1szT0XlISCzNOeL1m+BiopOk78ldaw8YJDdtMFBGRb8YtguVz
78JoEdZauh8Y4bsmbqtOo+sbLk+952HyaCZr47Sbz11s0PNO9CMl0eP/cxiR4AlS
N81P24jwCy3YU+OnE61oug==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5424 )
`pragma protect data_block
elhOc++EZPL35y1hsM2Ibv9HyErG/a+BTTlG8bEuJN3e5uAcjb5bagUbs/LDFAfp
465Xpgn+5CqEV6mODk7n+2eXCOfCBkHVtTVR6U8mN38O+1jV6wr583etdxFK16To
fxY6XU+j9wvt1+55Va0csTBQdemPRFSzyDB3xhP0eysQM5ay8mMz9CerDAQlbGEz
aXRrQiXo5zlWPI6xJX1qf/cTP05UQVzo/Jfq7/9Lune0xAD6oIhDpJ2576ppjaNf
7OAWQ85CITKvYKdS/H6XvhHd998Ez2A7uLJ8lO00+X63PPJ9vMhmdvZJl24L9rpW
KAZf0Gp0vu1teATCBZXLp3K5wIk6Vv5lLN9hRVxq9a9QLhoF7h5RxefxP7o8nVfZ
2O739yeNMlB2vPJd8i5zarTuUuKSa30SkM5KWvYNnjEHiWH1SqWC2Zpc6J7WgrDR
jiQW8hC+069ftESBFpw646XGqCtO3PvwfGwKeSVK2BN/2laqbimvVei4K/EqQh22
oMEDWwRSrqTQxU2J0eutLQTmVl+YeMLTaADViGAg7s+E+ZMLNK7mTAoqNYB1eU8j
eE/Q5zG9M/bEYb6ZHKmNUX5P8cWjtSxrrVi9/4Qlnj3oMBRnrUmC/lLmuF0MJCZG
g2xLcMB4qLP3Bgm3TkbkivkBglM4+8mcN3WheuVy1llq/Z7XNCIBKN+QOySigM9a
ch5K3DlLn6uNref580PZ7gkFLd5J74pTe+rzF2Vjgkf4gnhH4ng13UG6z0K0Ge13
wqeIopsCO/bgsz4NABKUB8JXhnWYOQxST7oEfi5TqRJRK74yk/tCuFYLF7Od8Fa+
FeR4rKNVw2QrcMBIxLWxrDnwHkZ0wii40TXLX+ijFE5FUduslKRdy5MTuTomwlhr
q+ciUisO3JP5+6bMUD0Akvvo6XV7ua7cAYeNAYxYCvTpNRnWmYXKQ6exaFXaqHoV
+F1JZrWd4652maszgVkGMoDtyjW2tmBYIgTxPL6ah2+hA7K9cTe6HQlvbrXfVr2H
OKGbxVUA/LhXCDMFhYAot9rHUfOIzo4z/dBHHF4rQefx9KQnrgtqwLunHCuMfX8i
sEJyPu2Zyqu9Zndk+z1eM6jl+c/VYMZOBIyJDyfWMSlEXYBpXPBrrj9Rk+IOQ2BK
sO5h4ftcrqM7ZRliEhJw+MBMNYuaUsz4yqz2/6gbhKSMH0g8piJd7PjTYROShevU
CYJhzIWcGY7LGHurZcKHmXz0td6NDMTWqLs16YO3GBFLBU59UqduNyexwQawGMyx
sAhTORlabkT8A7yawkG4Ku7jc5dF4qn+I8UCLn+2CBxESWN5TUoQz+1vaI5esDRk
vV5eyj/mdA8rQ6wGWTwjT8vxR6cNH4rTLy8kwdnvbMRBQGLBN60pySGCVBNT0T1A
i+Q2+a5bvRxsIfIVeuP8ta+dtfiLtteTUXxGzpLSxuKwS6/uajsrsq32zA6gMUlk
UXR1Gk1+AcWRe/8JbpH1n28Q3vrkgUyxewXNnxn/mGkQ2/SvHnhdVxbes1kCCsvw
Q15GVPftJKjf17pETRrsqu0FeQa80oIiM/BodyJiWUF3/Ntm8+7ygFG2UOJvsJBN
W0OsCZk3LhKks6+l0XTqCHM/uxb0qnidTK1fPfLwSvOhP6YJ2GvqFnw6/T1qJFRo
hM/HY0H0qrG0GtdXd2+urvoeyY33wF0RZ14Z24TOukGBL2ojilH0ffjcvGNSo+h+
gwuAScRbwawgdXjUjEoMXupE7EnQBhPs1qyN/m/jIEXJu31l0R1oe05JiELFt2iK
I9YlrHeoRcP7g0clsChVWBkJbFcy60r8Hm+4BDfNeQIGDpJ0saYO09nwGP2ywiA3
dVgee+PXox3uiWgAWJUSj6H0xStfGcrozaPl7oGz6GbKXu6JzR8ycFS1Qk9Wu70Z
TnfrkXMXorpS8g70crHqtVCl5+AsnLP0D2vXNARv4rRQTRCeOnpI7lpxMzcYaWeM
svdMTyCtrzLycSqnzlO8GpKACMt4v3X4afGl6CVYL2agUfDl0H4jka2/Tzgk7okq
D4Z5poovqO1Q7Ra+fHSxxFF9RYFF1ad/Ut6y57Ya83dFaRwlSUXvjfvQnMfvx79a
ACLdZaPNuRC4Lxa2KZUU0CHk/dm8L0GvmNRGphZ9qLgpn9pXjeJcGm2g5rqj2Wa2
1GJ415iPsaUlEErGUSRzf/vU0Oc0RGVA9qW0rgz0ekiQAT7Wh6/gxXwcJFKVeLvT
E73tcNYvxyR0a7a+d54aCEFLqu/Zz7wTZymrZqLc+i8OBiVk2B3OrPSQ451ab0NF
SX6+Y2+mDNlYYBiyB2DqSaYDBNMYq/dhd7Nnlsk4dz/KWl7HtZ7oiVaS1Qzvz4j3
2CZzXVzVn57PUYDL0+D3QSdvL9c5RYV759nFM1w7imLuVbRWaXjAOWkVyldvKw9d
FeELyRzuOJq1Jd218YJKdtdUtiONa/1co9ALhZ8oTDDodMgvgBYiq6O8uQdk006C
Tvo+lhXBlcmQrXRPv/nL3PpT6pqDqaVIblRmluonMP/ueLQFaWlADbqMDnht7g+z
pl3EVz1JBthY4tSN9HzaFgJ7dnL9yhvJqPqqYcfpi/vRaapuEyx6YRJi1/MP5a0k
epxZUL2J5ksmKjqijB1dY1VATgjEBJ6XjCwDYxLEMzIqHUzTztxF5MMcq7f681/2
BQdkWFcF3BZYSMDNVp/qI84cym1D/aABNwB3/cF0tVXoIxtJs9Z/zbKT6bByGMZK
hNTffKt8SbvSnhLdQ1TMtqLTzHCONNSBQtJmQ4jpbDbiK2g0qJogppvPyasv/P5+
+OifqS3REaY+3Hqk/78QOdqrLtWW2Ex5sBF5e8IV4Ng05Xkzhy21yzbJDlYuiwxY
ybBjqdaIE1QZVhUuL8bHkRL9IZGxRTJOJwLh5Sqiz34BH9bLMkeOxbrlZyX8rdZj
DB9ZvTToUHBdV3YPkP5KcSe0kSAnIpErUtai16cKH7zm+lzQOfhmWdrdXXHmqPwt
pfjpdOfH+C5z+odUyW3SAAA8sxiU/vuhNZ/mdaV/S47n1GlGImQ2HlPgSeNKtZmi
q8sI5/2efi5a9bgxiM1TdWpuhFwdwudWgP5m6iABFcOfO+LUaiDJJPeaxoaAAQme
DyVYPXEP6VAPI0Rhk0Okos7ZpqeudKowct8zUBUpeUCJvtyD7zka+L29E6yUGXe0
qgtwuKCZ3zB2GrQpiQBJq8qDEgeLswFI3BhmeUAe5zEGfHzLrmeAXau4wNiJSAHS
dBnjH+SSGGEbEupHinwzegZ3B43BML2NwSftOXB67ywraGGr5tQ5H4OwiI0Vxful
qP4H+PYLUD6gRGs8w22cdcgBjjjR0ie+ic8LsCM8umzauot8JL5MsR0yuMKgNTns
AploUWzX7fADug0JFIU3tK8WzGxHY7oqKnJifhxZREPvKxX57DzjZ64KrEsNXov3
Oa14DgSs9I0mcknrgQ1TJfXR9fdp0IVwCj3a/2SPq1sfXNPbjJ2pckahgna3J3O2
3EHWSWZvB6IxDzbvxeu9T+BLCrSZn1VGdEzZUiw5j1HheOJhuJ4HeybcoV3WCLZA
k0TM9YTs1Bq49FK/dJWTxd10ZerAQZt5NEeVyjX44pk957eWfpk+NUFO8tutga2Z
a2sLgqSk212hxKBoUbzagOdCprLXczIUDAJho5UbMQgAcZ0tKK/Akh7oOJpHrvil
AqWs+bfa2ZU9pHABP7bTgt6yBzWh7QT1oZc5eIR+H78NeBl05Q6aRUhUUuXbJ+IT
aIOslT1EVUHlTuy0YNtbTHYy7BcsAOS5Sg+JIjVU9pl9M9zREDAhUs9XC1SzuPe4
OwJ+bgoEeccxKWHvyzYgyT5OPhNIbOfO6nN4MjbwyYm1KUIBhp0k27OTEkQkHbv4
t5T5bAaFd2Z+/CpBPaamyHZcEtAk/SfftIBHmuhyFm/MyrmDjFPdQtQ2NL6YWvh8
NhUA6enKjBTfvbfyaMAEJcgzwg+Go6oaTDzvmiEYnkia1G/IIvp+g7mBCsS9IrSv
jibq9c3ayhdPqpILLP+rU+ZWcMqYg2NpSSgKap44bQLoJlR3UdMzQqt3lEn2QCvr
lw0rwMI9pcMbt5IDR/mgnlbUlVqM55rZU4x5ZgQmBCX7FnXLaczpCZvlKR79phy5
c5v3+fWrm0HcG4gfFep+/TLZyqPzH7C5VzqEVaHzTWknHxIGcbMQugUHJp1fZC8L
f3gCJa/8aNKOFrxLK6fFXKSO0qGunqHwBrTiB7R+LmO36CDcIyvijAZmFBTjtfrj
JzcIWJJs7fzJ5+9szZS6mS/KJKJ3iZs5mSLbIw4bsUM7tLino1j07kJaKdkXtczW
vC9IP0D2x+YGLBNM0LwvOGztfD0PZfhcBhfdRvVCjzGuATJUpQPaL/LzftUsXMSa
+edXkn9LxOxWILDgPpgRaUu4BiHkT0rmfPn2uzt8s2mU/xB9kjdDqUPFBpBrUHyP
KV2PnYWKfzuQnmHy4hA8TgpjT0kvbeA0856InMmeluXS6+C/qdanxA2VoFkrhC0G
Xsek+lagt0S5Mmo7fBfl1vBGLlcmmrmHmmjp2CORpAvxMv+02xHUmbAAgzQL2Qa2
BgOshMh9Iwn5r99dY4xtKKqVFqoahH7+hQtf40IkRWLvKVyOCJjycVCs14uL1QB5
G7fbe9wgvmh7v1i+jSrhmVxBxrdmdByMbJW91rP73dp9jR/EAullsGUgsptwvVdZ
cKgGFTTHEd51Wzs2FLe1i9ouiJ3xjYt3exI9BAiL0eGMOTWmX/7A03n9zgIcVSq0
+mgpUizm7ri7uQ98VT+Fc+eC/3giq9X9KZuDnh9MjM7aiO+6+j3NzEPNrGmWm03x
BPdjb8UHno2IspBVOhnV0rlSZEuomuKKZ2Kszx+hzzr0XhesqwLeoFad5NttxYPC
NrbCiyrjSx5yMIe+ZD+cPcYnELXxRIR5kWWpMeuU/B2fZbfAQhkZlROHSsLYQUGI
XsXKSDRdS5BDTsMOgyXEI5Z7eCPCJhZvxMISqOAvnTJuvRf1M30pllSTRADX5kFn
xAhtbeqmLTcHktmQZ/JrgiSoizBK5d7X+t2rZDpIab9IOLFG0IysLtgterdYWYh+
N+zYPWfFvmtqhqGr8lRvggsuEtjzzOBwGu4CIZgA3OtSm4myjV5LBYeWtbpShFfI
ioGY78bVbYYks/WWEGp3mebRbe+A8WaLLxoSi1EfBHINOMEjjxrwA4sbq9ibwW7x
AjeB0kftx3wn0sisg4XenfTnnbWfvGxh7v2ChYKaq0zOK4ZQ2hS1/77he9fss//E
ZCd4EyXr41KeroPQJIsamDH1mGnkw7unk9g2p4lrFM2qq96MhvO2HdkCF02KxEg1
xd3/WdDJ+L6NDCKAL9ZrUu3D583bJ8zh0zOTeaO4a192mM/uRbSb8TuHA6MF68GL
xOviIg1+3kWj9j/yW0hwl0myWqHqlAxjqs7wzv7S4C+bQ7JApADq4mu//rNR3EgV
8JzlpBEYiwFyNqr8rdz46JB+qkX/G19r7RQrQ1t3QzWfGCYWeZMY8nqpKMs67sTv
iVHA7HijBKlndSbd50q157bZNmJCHgeSFRXCBd3DCJf6VMNteDeYkP4XsLPJA9l3
OOJgPDmch8ZH7RCbrcx3k2FcL6mwRRH7Nl+93QC8J3pcNpzEBArTCtjynQq9PQOE
hcrC4uI3SfRJEU49NnGe5oCkEQa/CSw2MnrVZujxw87JRfxUO9pLUnue4dUcKRjy
hXP4aYUSyVGU0IAsEUuhb5xU8ri3zQGlZ0TuhKONr62ddBZ2wcNbu7xihztHl24+
/YAGljRdtMSvXSAA2IrTYZBcPBsl9QeLjSeG4kj6XwBVem6UbaL9FW9FmmV2HUnc
9VLspeciOjC+e6QIy+grbhsMJ1QwVYQpwUVtj3RhS9WY0le3nTpW+/akEdbzMS0V
BKz/b9YFqXbODNB8MOjmu6aLlxUe0it+Mg5aXU4hAbejNqZEY8AEA9RmI3o8pAYk
zYTBIux6Q3lsP/fO6ZVjmWG9u6jewTtO955rusuUjNTdXXGEMwN/VAsC87cDp1A7
IoLFLA2TAP/eJC3rj0n/fCwQO+zkSmfHzJKqde34nWVnKJSdnd4f6CdXYPjh0vZN
I0aPCq11MZmKNQbfYl/AYa9wBeqBY972yPV3/ySn2Gjy4Uu31xIZ3p+iaWodK8yA
tgnXYDFMW88xzSgDau8Uiu39dwouwDpvDjW+cbmJ+JMHFNlsEmsVf9J7tPDik/2i
RlbMdPGGG5El5Ow9DvBia7ltf7UHezMB66FLmBz+tuB329Xe6YPEStDpD8JPy6e7
q1fI48Ct/lYMviQCBPhovLGyVdyQVMGjh3upKtJm1/+icyfpvi8JJ4z2Y70Wkaf1
T4LWtiAKHeX4ZY0/VrxHb7P9NjSvlFIxbKvRfRc9a6v+LeG0EwnOtk6gFW0uRmTf
jhgtUOFnbRVRD8EKUhTl1c18EyeYodwL0jq4Ho6Vs9mB8eNA5oaCy6g5+rcq5Wrm
YKl0Z5PInMd8G/NPuShWvOb7Xcl0Km8Q2YRBt8YO7XaYOlVNK/wGMJiI/d7MxC8f
IpR4quAf+Any6dTnilz91oZJq8jZPVRyM5MhMmnH+0qyMEpHPiGRX65hfdiAjIkh
zf/QrVzjvl5BIlqC2dvxOs4vLF+HYNsCUzsczfOA9kgnCiYkwYO6LsyD+U7jzGJB
cuC4rzz+3Q60/yLvsewQGEx4N5FIk2nOMAYBbqlfkfTtqjSppWvtFfdrj0F6IFKX
DbDlnKbGH1i9ZwLSsE672In0lO83rX3JQlAIBEARhK/hHkIudQC18IbVaIre7YcR
yQMtUNLJ84nV78LEJY/LjcxiuWfUpAI3wuf9KGu8cAyuJD9NpX0emvKtn8Ni1qm+
Zfop7cEbJERW2yeJ25FfYHqu+iBpBnRo/BDzKIGx+8GZqhG3w6CBSDCfUg7wqhM9
8BC7ubVsJoEqH2pANJtr+TEuRUrWZJMzTEP51JVoNp6WmeQR8rS2EIyvYIReDp8/
UuvLXq6l+RkIVSD4Fgj+rsjwULJxS+3ImmbwzNF+qOh0KRf/TowI++YE07ercPfc
KrC+oYFmxRIS1sspwypAsI6BGAK/aOvHSlnVi08r97OwNLR1ZS5JwjWofEfkCu8F
lj5gdpSCKRyS5PmtYNIiDbd2XIcR7ZcltSgunTXyTsuiiVlDVpBKjr0ddplDERyI
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JuXmDg4Ai31cD5Z8RhQZWRSI+GDR1HFSGPoMMTpf6++MthB9iHjCizETe6FeWolF
dYXlXZtm1NO8phbOXFQrgpN69kU8rac6ZpXto2EKeRmVbxjjuLc2jpXVpF0wHM8u
O7z3ga9X+OY9Z97JMpJtO8H2jrlHZgiGZRygm4o5B0Pew8xWRQN8+aFZxGech8IQ
fzSeeE+qdgtaUp4V6AIKGmRLa5YqiHF+ZRzgsY48h4Huz3G6jqWMBoinx/P59/5T
h5KEIo62MFj5Z45OwndMm7M3LYBW3jR84HoWuLFR8a8SLU35FlUGx+AarHcwvHMN
w53DQ9w2feGTxe7l8DH07A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6656 )
`pragma protect data_block
kD3M8OQO2PzuG1NTjUBKt7Nz3BhFv0MX80FqxfAwXs2hpfXkB4Tr5oDbhvyliVKo
oOC0h3r35FbD2DGMg98ze2dVf7wCpiMmRKHgcVcPHvcaejUDBJNVLeEdbK1fSQTC
HlEVQkpTxCls0hXuHNzUUtoQ5Fq4NMFdeBdXssm2hmFyP4zs93nAgUP4ck2kDKKW
ls9TRtIfuqdC9fyEfexD8QWHue1SLzJYFi6DLCWRxjBjKTrJsPX60KjqM47vH7Ub
g0goEkfo8l1LfzwynMEX/qOajFcw2S1AWZ9blJqQTprNxNWg3oyzK72chC9QQ9aM
1iCqaqizzWB+JPseAHTYcS++bClipfTnESTK6ORmvRLkVlsmti8lsmoQqBrHUf9f
xOgvK6lObK5gNvyiwIp0rDm6f8xDxVpATSqLWrSLtIzVUgyq86Vp8TBKccGrUqhg
+gC0Nj47ksVRJLGgYn6K6z/QZQ9T53qSXHxtveMISpBGHaG1zXyd1qcRHcSqrNg3
b5dYjeNpmahQSxs3INKWD4vf+zmSo+Sw2BqJ0IHdht6kUqEdhOp4M0ktn9Xfjg8B
VXBkSRasuSyV6CgLcyyPdm5Cetd4VFS/p7haamqxOfmR832KQL2LhvFRXk/4WSYW
5t31AjOJTQd1YJrxhYInIBphEo0kGODAf9DpSJZdieX+SdbNWQGO2SAyx/OiZu5c
QeUMK8t5bxSMtEq3A3PeYFUxrENSvmLXv4W9L1mL+we8rW9Tl0FT67LOm8FyzPh+
c2HNHaHmjiMHylzuWz0RjqBMVsxycl6VYFnMFXj9kSWISrUsGv6Plse2VtV5nGEg
np9sDCO6zsq9A6JRytiPc+dW5skWCluxJCTKyzgkfTHlxUiWRgtA6HM14tG82RnA
7sESf0R8CzqhKGhniUylOL7Ho/QJC47TVnuljjiXYIXLgq2yvoKp3/bYm9UcUMhL
D1gqi2eRR7upjax4Gd/K2ViI7HbhRnXbjQY4lsxCgJergxeLawiIzkReTIq++t2U
EOCpEzzW9p3hPIjVE9wSRCWOFuqcXX3YwUNO/J7P/58gkQ/A9P7uvK1rD54XRUWh
cqTnX7HFO00ia7CEVMVnI7GGor3y+gvUFEdH7Pi40qdTGwm3dvm9aHetMlRURJ0t
siIKuaHehrSlIDnLw9iOJOpeWPiHD0KvURwfcNGJBGN52H99xi1mlkJDkiTyCgTi
6pRqgKTL/owMhEkAFnScWKeAelYoHCqguQdur4ybLn7Vbq4WdjCN1zrrGotPIHnk
/EMqweSxEg1xMHgeSKQANVxa9R/3PLVi+6daARmCadsbx5eHPE+RNL0Aa/DRuudz
wfzKWv27OLdrhvxDi/7G9mK2Re0Y4dEvh5I8NSnQZeUNvL8oSrZZoltqKgZl7x+D
W6DArsb8EGtz/VhMyMHaqnwWGvM0WXpnElO/8ER1KemMH9GYt8i90TUx5tPopLL0
YIckogMVzg6ABHFd4b34naOXgXUcCHnd/y+ei95BI1Oi3jYlCPH7P4zZ/rS5DYIS
SUY4xT1d3CsFQNBuAPNqfZT6RuBgA548m26Omi0dpgXBH7K6YLT4XFENYgjOemry
gGWypj3nEin/6rIjDGYeTbUp3ngKv3OkAQd9Etnp9ZB1jGhSg/GEyqxOqz8e2d8l
j7spcm2RNiJPAq9e3pUD84TALAam1mIWLTuKsPit9t3z83l0RMnq2WRfYWdDnUnM
dPWW6dp6QlOzxHJy3K6tUC3yoeFlieB8FQhzZljofiMOTac4s941hWYSTywqPsLn
Kh+LbFBmtaK7VPK8HI5IqfxrFPuFb3hWCvvUWTxmOP1T63SCZMhmUHDl60nC96bV
PgZzpytpZZlTUFFrHDfqDY+ooTiGNwJxLnl0XRn7fBvsGMsRjsAljGjDHGxHQZ72
2pvdROQV6Bu8LTgHubQ1JzNUJ8HB+szsKVrADnfJfYclV6JdTuDwHvlkA2b5qtkC
b3cr/La05WpuuNEc1vr4a6F2m725FnpYppade6L1Iayw83xPuYKwO1VXJmizHoF7
p+QtAmHi4jBF4DXlPCQdk/15gEhzFFfM5UD4eWYFhxyHFWUF33xXzbKC+4c1HKT3
MLWwO7yVGJHkZ7sG8CiYjE8w0pmmIp1kyU8Xymz8qsSHkry8yG/7d4mCO6dGwCQK
qJ/6yU8aMWefiHWuygP2cyEzfz1nPczfUcc11wGXF9aZtc/QSOLVV/fmH7nqD9EC
ekLC+0ADHu4VEj8W0PQ1THqZdNGOSvH1Iv75u1rz8eIxxjRrZNPc3eGDjqTuM+iX
uGb/6BRjXt3SEj7JyjQt/bTJqFWwDkO+qX3ZYEAOKVfunJsndzJNm1rvjKOD+Zth
Adj20p8vz/Pwep8AZMIBz3Fx7b3l+SvHkAUyyQBTrGjJqaZVZKR84x/OCD4aBF1v
pvmEPbmGsHCkOaK+rinOKBjFfRyjsytZjpIL8FAKLtSkAGw8WqbdyvZeNKdmYcza
nNOxTvE5I1GX3/lxA7dlVOmCFufVOrDGpLQd6AceHxyQEa5kgzOewnsUh/8NI8QO
dtUDNW13u5p1E6yIbccg26U9yeYcg0Y7odX763l9BVmcFvOMfwYz0mOXnXa4LJjC
3sfJ8KlVVg0qe89Vwm78SLonMo/1FgCLfBWuboVp6+JmcydUNttYJdr6jcNslcpH
puaDAKmgovX/hymr4C441ZwI9BUbs/ralGBl99vC4Ap3BpDWdJPW1qCnqYzJu8rl
wkaqwOe4Ft8vsaPtFF4IPquVjNyezsX81qULo9pgMPJOnvy/kHmpobIqTwP9F4O3
b2XH1Up44HUtC77wIRy4uGFzqxi4Yo1x7TB0ZszO8m7RGVMCo8eMtRlE+pbRt487
X36Za3TZqQUvpAT7EQ2Wr4HPICrSYWM5sLWc5dxH6apkBaeSSag+ee/iDpC7qJ/W
nUDud2dYW6yeRuuQwpJ2HMU98QPCqfEzdv3mDPjLe3CajdtLIiYD3+yzvb353XAT
HvQ+x4JTeuZEw8EIMbLmUC8QDz7lkJZsubs9Cjmw5g2ESuKWIEe+wKlpXpGHi9fD
3Z6scxVmCogjyXpSXK+VOUXVIL+GFI366FOlAE/C1hbK0lq8uufh/IZnK5ntpDUt
U/24hUrPOTJpT8g84YtmAgabTJn1uWb+gsj9TJT3Iii0N3Nib28hmroPDJNpWerR
ZJ0wYzBb7iONJhjdEKEQ0NttpUqiHB07Ce/jxsrBrcSA41tGS9mILOMFjrxANVNO
MHME5kTvrORYNQbR7cxNA3R0rbyn/1Epzow8oU+tmG25S2TLHSJhKIUdFVmt9UxH
eKhuudsFw1UAEEiUTJGcKj1Tt7ZCafRd7ozpIbgo94LLSMndOgY0JcZv00TDZeil
PpQPuNKpt9/lwUt6VxSWRuynhsjp3rY56R12zpIjAmkIVcP4nkRtYaP4IwF0MWnN
2ysBsgwFPu1WUUNxpbRoR4JCLT19zOeruBRNThCQXtZ7rkTqKOwESsky5LaXQdvx
9392563kQ5TWGnN4qHBpCDXvywi7d+F8e2N3JytUONADTLpm+Gwz9PmvSMBgQXLD
BvKv6UonSCIELs/s6qYJVKhbtSYs+pgyn/BrpLnA0/LI4Baa4kAqKthMsFBEhzRx
J2szgmtZd2juNF2kVP0QZryftiQ2xQkzZtR1P0FEQM+TUVCqBrErluV5qZ9tfFeu
5HmX3YU2c/naYX6w4DU0e+oK8VUpRjdKCWnRyQEj+H1jWZadG7DRL1aj9uUyTGHu
MSB4D2vqxxHQXZQTDKkEBubNrSrZDasMoxvb3aOR8ZBK5ekndVQkap+L/JEdofBR
S9xjdoqnE2FplN9Bztapq2hDYNZ2+28CdoNkLeE9oI0iiFOFTnmtNm2MChtaPzKF
mNDDmZKLicr9hx/OadMutisy+p5rnnuTKqBuG8MLpdGcjKnPWTkx5WhA0+BUyfgc
u5cXAYkW4xPDkxBbjNYR03BHd4dtJ87PSMAhh5IKQ47ECgNp5yuUNwGKPNHjtXzn
v5z+IZM6iwgWCst76TX9v7Kl1nf8M0wgzPk6cUNeXwesJo7MGubQjwLtC9UX+y8g
j/4Xg8DH9hBtwNbaK1nNCU637rmpWjZ9ng5w0az2kJw9JDtT4EivHXszZKV7/qjI
CiIyrx4UA32VAzajLNMnkBFGNre4OtO9FQyvKvfpKc6gc/FvpY3EAuSz2UwqcGtH
7CuYhAE641BdIyOZjioXZEf0ng70WLn6FwO4WEGBkmxFcpTIStPnrgeHioTe4Uj9
76qcKQMe0D3Hn2VsSZyds65s199NV4b92KB4jZYZpytX0TH/VjGnYR0YnkUfT0aU
XENNQkNkQnXxa9s690fz+6Dnxwuif+9R2YUleKlz0MTptzeIXC7NytOyFDR7Teo/
Ig0Y9FQYVaFgIHVGcoX8Zeh9YBFWhmaG/AmG76mzmf2F927Tr7nETxNdKaNbAfm/
REQve5pHThsBWvF/dj6+op7c6XRnjBYCLrkQdCQqnD4tcGuuNXIPBigxYXZem4Hx
HcFjhRcpZViXTGJnH23CMbLCv5xa5Cn0u4OX0rt04tjAwdCrP7hjh2u1LFjIAQ+w
n+zahLv1Mr/1rMCjIxrgV0QiLT6KOaW+NC/k6JOrgN6AqQ0TvFnLEA5x/Xqkmtbg
Q27iWhM8Yr21faes9CRdJhplokOUmVhxmiU2RcJvm9JiU0zyJZNqjkcinCFjrYgh
3A8MHwfnPzohE6yNaKRN8uQfM/FZ3PxjMwmatI14L8rNLjBvIOH+jhIb4U8d2psw
UU2FsC0CgSP0Q09+xfZXLrNB0ZSXnKIJZknruZ5q1TCBALWinyG3XqmYT3FpRX6K
yhQ7b16hL0P3e/5Xg+UNowOCfc9lvZUok8rmR7/qfnGCrnlxXnlv6H4vrPe4DAK4
Evu3pU2qNWTN9BmcwoHLEvV19jFnobPnTY+hb32lCOyf4UX6inD8zyzsLeJNg95Z
Cv4JA95GSYPwQ///XGonNYiIRZKfl7hqEqMSElFa7JiGggd+hJseft6uBERxpI0Q
rubURA6BZwC5eIymbLX6DEpWDjzA+cIy5cxffcpSsjID0dbkbT6DnckFtgcZvT0f
DAkIrlUdumfGt8AjlJ9O6JtQCq/9w8YEj/DOS+rvHAds1C0+H9fDte1jYZQm23Bx
sRbEaRzPNl5XcMVR8oOPNDtV7kGvav+B8ZK1qaYHLUf05FBFxGNQM4wXJJfBvGbV
fb5aCL7OSnQ2s5qcTp3m/lfTG0WurQtN/kk16lPvCjEwBYJTvN9Fa+p4E45x9SEN
YXw/P3+caGfWIXxEXwxEnlOs33la8Q0tUfSho1mJNEbasDm3uuZLYg5vbmWTHUno
X+6nELnrTdk7MH5MpGL0e+RIdDjJJPwAxHrqqT/955B9sGoZUEhqiqd9gpctwFgR
inFzoX4pndgMXEzBtVLwBP8YTieTFx+6oTe5iR5QuGD5hOQS047K0/OVo8pwumSk
Y1sOKuPckXBIkoMru62V27KOq61FvsXa2gzkDHMDseGnfK6Vvmmx3nkONoqmS1DU
sLzERUkGpy7SQjYKRIQEudRH3XkPtCsgz56SA3RjeaaYfJPF5xbx6eqjk/HEbnUh
YlWyw8IHaN3SlRIprVW+3+7QjNadz0NmqbDQ5MPEvU2g2jQn0wOXI/FsZ5jUk0xS
xrHloTGFXi4vTy7+BiVlzo+Qo/YeQE3ow3JXROpUfZ2Cguejco+p1v//DcdMUxWZ
WbQFdVYqPQu4TzYTHxIUh16MAUvdZ4V+AxPXrg1KN29UQ2uzgMkfhjFtejBBewnk
TMK9LL2VZQDuFkrSxZ9ASe7d2RMoJ9ThvDFp8vWEojiwZOqnxheh/sYs80utMmy4
NQXs6lOxbdyfwyNnnyD6c0IIx2x+q/d/WwH7O2Vdrj12063+V03YXqVIy0tfdG1/
i4kkgj7lD7P3/R5XrTcjh5LT0hXw5prXj6FJqLjGtgVTAqRiqdY5Y+fhx4uZJDfQ
XHTFkKbhXX2StHVwbgFFS8vGbb6+SVH5a6BuuAMUsLTYt5fUOGngJYJmVw2YeE3y
s2/Vx9onFtis6QQPPFfdotcW67c39SvVQjo1klropOZsToE4c3Q/6z/ghJt0EvfF
6nwFI+Hx0M7JqeZAqtpZUlaqFwMDydiLVBsZPLgQCfnr3wR72HdVta4z3tcaD1EF
KmqqgHidxjvSH2bMk4rg/zIXhRzETs8KwnJuGmkLQ5vdDfhE8i9yQ1qEyzpRw4sP
DkV2eKxgdjYmZIQW5YWfkEoe8qG8Tl+mA+rzTKKxVT3KFHu7yAUWQxyzihhTnQdT
9aPLmOMPHdiz5HKQ+h4uYMXJhhLvFA0Vrw1IQejOeNXzazGkkce6gp93tFJB8AKT
ouQmtY7oMc1Sw+H4AyZVLUTNSb6+dtYqPc8+rEarjQOLu1J2piJP/MNbW2DlLKGr
kw4ZJX0vIlRm+Bf2qplYc/HTkKLycfvxYa77msheCDgnJDv6ZnmkJzuBhfY3pfHl
sbGWca+YqiEx+DF3g+T20FIe6H1//k6u/qt0DRFmOGPgrpG80nLrvDpistW2ET/E
ilRcrMy89C8GK0bYnofVnBbr557f6ZVA6GZhxu1dGVpspUX8HTWsb1G5rZoRV3xR
ZM1TSso/rUXqCzWSO8e89ZS7elCAylq9hGk2ICYME4Fiwul7/MBz3FY6MKUQR1ZS
3ko85mtfouV/DWXQEOLT7wm34VfuRXRjnvAmnie01Bmm5ma9Zj13VqIxl585fKRS
UxR0b3oEh0H+6mK7e6zBa3veRVSDT+/amGmQ0KlLPFB8a75WVu3kj4FyNY7NlZ1t
e8EoIPLvkoHcCIPBxhyeunMpXewnFIVVk6f3x/UQPq6IDveox9mz5QbxvoYNuoye
IKormc9zNFu9L8x9w7oFxRld9yP7d4d2rG3pZrvfcg/WkB9pnKa5owK7WahtaHKB
86LD8dMb14CngK5K10SgNsGN/BAyU5Ej2vBaELLTPUIEnJ5euIFjDCfVDgzffaih
x+3X8d03xIOYy0B879oUAtf/yqUSg/F9ynMkjIbEbsnDspDZakqEV8kuM1tnmbMU
YYg5GK02vbCyZ7zbM4oaN+vhRd1dCmdx7kZhmE5RADxv4/2kTjnXWMVG/UNusnUP
bxXdcUdAP/sbvuh9TFnG3y767jY+dnhKqVwl6AFOBB9tUg11FT3ItZ1pVY86TDTD
v2gPuJ4SGidQPOJgLAF62/sbMs7eKS08vZCkJsSDldgr4uOcnqNm01drneKkYu51
m0fcQC2SwdJVNP3ftOtiF4FdZy3+5jZyJx1ZSv1GhCkOBj+FLvvDOwbrESOILbLr
cknXiB6kkfNfV+mFGoJkdzpGGDhiyb1C3CVesOM83O0um75VRhokhzl9tPd6HS2f
A/KKgx31nWZdSeCGuxJY35bt77a6/GJmnR6s41H6eljPQRLcbGfxNsEawHFil3Dh
VojZCuVp1aJ3KIwbTPRTLckiZxbn7ViEGKx83LhR5NDCCalyUrZG8HkGbioScUKt
cWbdLzbo/FiKvYKM5dltNt4snPzd+rXDT0cuhOKm8hChQuq0HnYJZWieCxgS1Uk9
WTG6fQeYCXSnKybZyvppQY20EEb29ciY0fEGJSzTm4xaqmovWgloy11SbMAXKOEn
Gx80G3VwLbtiWRbCjKLJY0h3GUL+KuY8l5Df2Aeh/mxcSxwLZB265mXsDeehoHdK
YZXekb3/Hqmr/nI9Fibzi9sV2IzELTzRdYH5gAQWStqkVDmHLL93nDT0EvXxiy/x
lR3DWnMXHEczcx83JC0vZyjNY5XrXzJhzVsqssZPKSAq5kcpLcsGSFnhIARwzpa4
LbNKcoJGlRcl6zy81rMrpOJRRxxKzty2JwkQcX2pUNb+2T92XRMRm7gvT03XeDCd
q83A2UMm0LEML4V4LlLfteRwoB7ddpyFN5sXOX3Sn8m0zXITI3monBNF+sYRV34r
baCflCv39uFkABaE+BkMJiib46ZlwjWwYkauyhAa+1dD9FCrWHTh02NbUUYHh3ke
5wJT8qBe33DTwH9ZYnPSZ3OnyI5kCGbi/f/2PG6NQKor1LD9I9ZP+eHcutqTlaCC
5pf3o2oxNe+CxkYCqFh9GOLPibkaMoyJPLXfB9exWatoIq2wpsOokiSBgHbzx5eW
kZ3CkzzslyEYyvkt2+tK2n7krgkXKNagH7MVGwJCqBD+FzeSp4zPPp+PRkwvxOVq
9tbmTHiuleq622Jlc8NY4gEJxRFbMSLzGYymVZILE8jr92owuNtGMwptTdmCtd/Q
KVgKmlSesY8CcVGDG4++G6TDU5nDy5pckJcvDGV7ed+UR2GwTtCIFOMRJAi4ztPQ
TOUCfgnVXVK+lJ4AqvuJIdiHDUZNTG6awFMNYRVDybUNK2X0glPdUuorCunXAE1n
NK/gT/WR0ThbjYV2q8j345+rBq7VhU6CseJe6qgSbZw8rzH6YqZ+PV9Yvc7ZgBu0
2q4vgGdz0i0sa1mo1bvCr++BoatrRZFZjvEPqG7eljqMlaPVs0Y3YsgwVrZjl2Bf
3LU8FLL8cQ4e4d5o0lKsoQERbik8mnShaeKAvLcfKAA7vBk3x1KNBu/2GKaYHqap
X4AcF5YGqUd0AOhC27b6j6LVrghMTGMS9FMVXmIki6A0pXfnwI3EzTg83rttaoxf
TiQ7EfoNU1Z0XvZr9bvqKHvCF+VORd6uDfyh8SQrqqXWV42cFSBE9lH3DZiSMRo9
qF3YSA7vvQLPG7uxd6od7VjubeDJxEbjfQmZOfJ+ieJv6XL2dCixaKs4O9fBuj7b
R1hDoEYtgGWACkEsepqpgoxzKMvJrYo9EXSaNuGgqVk=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WxBLzrDJeipYuilmC5y9d7JleqvpuircBeHPSPCsqvbzXwVmkDTxi+E1EVCoEilZ
3p7kVGSunpDLcPGNfPY6io1t+M2+/DVwwdOrsWgaUuVavMUs5oB5dIol1XyR50Hv
EyvJ1TiwQmkdvQP/kzJJ24nI5SmHcT3UfzlMvTbh9ZKvz66v824l7USd8t1dDOXf
HWltZKUei4axMjNuYGT5QNKx1lYJs2dhZJm0o2/B5Xexset3B1zcTphM9jvTCnED
KHZ4dIaZLy3geIqFLD4PuQnK2sZNqeadpxkbHl2cWyYIXprvD8jUiOCcscO4M1dh
s5jF1S9WJpSE9zYnuJtMDg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
rQc6OrdwxGxuGatmMJzqFWUAMZXfIxxdDbDrE0eDQ/yLQvYs+62om0tm2fv4Xet9
4UGUyop5s886jWp4J/h8ZoJEjRUCRioAUqg3JeHukXi5TIAeGPeqa7YllsHtU1Mf
qcrf6ByJkuwaEt9+Kw8CVfwDD+zmSqvCXomhvHLgTHmZO9Ra35CEWp/uTS1Sorf6
wSSdxxWsityQlAPI76jnYZz2oFphEnOqGDCGDwRd6UE6D9RDCeC6wXYgeeQman4C
ENtxDU8d8aKt0PiJy5ESw8+2wapc18SoHCKc/Zci6jjLMBneaaQh5X92JqBLV0jt
Gw/xKihDCAIo+raAWEeU7yzuNf/iHFBpssZc0brs2iAn9JI/ITCsZ9VWWPn1HDML
N9OUAGU0WQ+2pMPNrZWGmOcF6PMCzsYjiBlSyKkTd0AyivP5Op0z8fU2Ah/9TQqk
Di2k7077kWysWG3HJ521UnS5xMeqEcS86pqOyyP+Hn5y8lREE0vXCTX1f1Qe/vFD
2yi2YF9TnK//UECds6FgUCBuVuw1Da3rs0KQj5Bd97SYfKDHpuFrql0bOYhvxPFx
pDn6iNay3bR/z/OXW47Jf1NK/OLg25hYmPlIewqrB5i+/L1z8YxIvaDG8m/07gCh
Kie0X7WBCOb3CxhVVbNcUO6xlfZpcxfPgFyHdBNiueZMXhe55K0fRgGF9S1SzobI
r1v5IXzHY7GGS0fgn8ZqW3LSlJti0yE8k/ZO6otua1lpcaK7fKZxoX8dFdLh12DB
Kmi5uswRFU9ADmeLSMdkVRxQB4HCMrEXSeiKzdceUuquc93m87+LlzG7vhuz65Ro
xd/l2Sz0h8ApBTxpZicIRy0a4j7BA24NDHf492DirhaA/lQ1Hgs2yiDLHdPbJABT
IIYBtqDbdzTDlvEuTUAv3b8XGwyqMjaixi/+8uRn/qaTdr7deUvir62l2unmmKJf
eWaXfK1HpMRRJ6vecUI3ixOE20HX7eOZUhL5aifxbdL6+/Ob6QTXjCE3/aiU2UWT
VuP5WCB1uFMtEWajfuU0eq7VJ28qMLnMVHGe8YmDX35OHiQ+Wb+MAQ2TDxTiHzOm
RKgcqejwm/oi7LVilSX7+bFy8CCmQBcNnbg49ocHr6sntZQvTNAeAKCYb+vCEoZA
ZfOb6oSephZNpOIQVJLqBc9MIck+9+9OtYCRh7jyHXclMkS0zxnP8gXBQxOQvfTs
KMOPp4y7DrpBOYHLvhs27WX5R9nZ+yJYILXEK9xTYCs+Ylc+gkZGozrgJzaOV1TK
cc7/tnUTNSdcY53HWioaJ1c8SalcenKhwlNPsDnSv9nOi1wLR7x3bbeZq6tgmJyZ
Ff7yJd8NDG7NIUC+mxp/vKOpZ8o+Wl8/sZJEQUOdos3VIa4KamICXTtDPjwpJrB4
Q7GXGCnDyS9Lj6Mlcn9ssVYtkWwUQBD5CFLirXrwp3AOx3+cfcheWBgncdXjNdFC
B3G07KxMItCYzcNE3JV6S0N60FA87KeFXKsssZMR6TluYTzU15DIjYx8y64WqU3r
34IenDOiCxCxUvlmosfvqQkhfanfpUGCJgnMHkXkFS3CvdYf7e1NjlE6H1c46dyR
lhPLAmkh6g5j2w2KLx62ldy979Nhri4Tecs2icx/BAGV7b+LwNNiDLGYhAPm8NrU
4k/cAtKTdPS/r3TZMTPdy9JqLI+yfJR5X19OXA8uOK13tW0UUSSf484uJL6nEwvk
ViLjyFL3Fz77OvBFeYtR7yS/njgb0xEFnO/9axNVR+lJwwWOQgTi6GYXwKIHtZPk
LIFuOq1W/rttiSbRvsFIIK/Qk6GyGUamOMEK7FIRVSPUge9umpHzO/x1UTWaHc+3
jsNfnvIo03ngyoluuz2/W/Ox4HwoNroaQPshKs8wAXwF1J9egUXoYRz6aRKqHGKj
wpIGNUfFNE+bLMHUBSJ6B4zRZJrZJzI2+7gT2k4CfVV6Kml0NRRVushCE1UBb4NS
Hieno5vK3DeThA0yfn52TFCy01iGjocef2ZsLvWW2EafZ2UFG6t63iP21PhYx5Wr
124uAb73im2/5uVGAIDVujcQP5UGd3GvWhB8SIKO1biMIu8IhaUg0zGcstURLIkb
FYwLqorj7kJWsw1jPdh5WLeM2FuZQPv3YcdwMYJXrhdotLzguiCq2sdGODgJPys+
o4AqHcLuRgVvQYH6Vmus73CqB74v4o4wiSbxdu6ygGGxFHob2rI5LvZ844TclsEv
/017y8Pd6LuvLy80xkuofFVHQv92nYxJxGnhF/XSz6qQy7Oe4y1t+Z6n6hVGbDI4
AkGLUtX1UAC71o214V5t9hoRENtExFd2Xy4S+dYkZR+RD/LKm2S3+baH1Dn/1q4a
QRD4W/E0bhgereHC2eKAKvZ27Fd6zXeUymKpBxUbudnhzBzquLJ2K1ZBDURCMjQq
v5gJXdGBDrtHT/4Wrb1VMFMZ1KGoOwu4G0dT36S7fkCNWJjVlk7OoRLkGqzqlnKE
KSej4p2s9AbETkFEyQtHixQZ8CzDl0b3EnUNf6YooST4lAk3bU8sLOMwkb28QEdV
rWWTSZOzH8fFCRvgMHI3jbnqZvu2R79tr0fL3QfgvzkQLWYTl7BbmPdxN7axEmt9
JJJhYDyTHep419HI1RN90wGlkCpkfz5TuI4fHuLsyB/0Z72gkwA8dRsBIAJcfYCj
WslvQ2pi9z0R/JYuHCX5zDoO7hxfKP4iK+KqMISiORwoZcPdA/GJd/F6a7ot3I2n
H1UDRHAQt1lbhQcVLgheDFkm0n9pbR0bqLqSgI+iOJ65folTw4RMR9AjNQ1MXe3r
c19pkUxcLSyT36UiLW9icsqKRsueSySmsOT4hT0/sYUvGWTXJMhDDTVthRuA5h7o
Ro26rNJRr3Oh1jAX+n2pk3e4JSP3QMquDwXdIb7Js1OUndaKBMLKIMbhyg4cHABX
w9gLmOkeZ1hoesN5uTyiahh0fGxuy6kLhgDmdC7UgCzZZBdDbsxs5wiIt8IyQKqv
5K9DAheI6eyT2PPW0iiS6ABDR9HboSp4t0/uzShvWwn6XJjymZRZQmCo/Dc7HgMS
nT+8NpgrNQ9AoF1FV9t7T6W0FUTGggYCMGPddLFuzV3HXzADTRAWb1WJGMcnOiQc
O4HV2U1UF/0kCfTty3eEWGGVHxhHC7cTneYrK9Ip+mchwqyjRzUWxUE4Pc+uc/p4
AaQlvSqJxo7B7ja0NzmekEx6jSiphM3os55eL45ZZPpzw9VO8rCBubeXXlDC/SYj
ufAAz6a9HGaldoR08eHnBXZIbGzRVv6RQ+rhHm26/CZL/r5pbJ5JFjvoNHUd1TXM
6U9ShTSSRl2hPA44QTG3w0lz/mB1ra8iDGmLRY6IrR3DHo6XNgZyUMTEj2XMtdr9
1oH3Y/bGPpx/gP7zoHuDMXU5jiZXi/YLaS0czmLo3bJs236TjIfaU8yv4bX4Tajm
Hajag+eOwCuLUX/+MQqJ7zx4U3Yxv4EYs6QUR7aniJGMvD6/jMZE5i+eDWqp5hN6
bj8x21dTbTs/W6A8PAVF0W1l/2bWSy1nylNFsMLwrog70nf5UBqeNzOi0/xWBOGW
rU0F/omjDmqQR53ILsxafKI6ONefnlNUC8jrRsPZTXIB79GI/dRQ6D3y0WIe6mdw
KQHMXSASl0X1yHbU/MVhw2kVhhcqlD3hBRC22uf23sg0SLDCDLPS25mpZRWzOxIm
P6oSLhpdhMqJcINnb/OyLySzHDvEWzEOXIIEPjUtiODP7WU0qVYnWoXyDFRzrmW2
vZEBKBuPFNMt5vZ46z+ugC1E9F2317zlbJizXGdgLpoAl3Qx4DF9h7IuGQ14uv49
QAxHLY+/D6nn7qBbJK0hKx1xQIvWHxPr/Pjd26omgt6qTqBspqoOtCY9BwBapRPO
n8fDqzs8i4riaP4NBbQY0nQecx6kLjEEq7x/t3P94hNetRbKcZlsikzMNhh7HtS7
fUdIXELvjctKEGVPA/zaSwID1ABliM2d2YTC/UUQgXFAQtw7xTbJTxbtugR4y+GK
Ti07+6WMH6bXKXE7Yn/VbVHHYHIEnOT+P6Jax/ap8OC5Qj68kFYCYMKc5Wke++nt
Bc3abZn7IqClbtsTM91VTUfsQNVGHVSDG2b3G1BJhRvu6DZzAnfA4rbfdnz2Bqgn
wCccN/DJOeIQ2HHRllGK+NpkaRS0al7YO++96vDXumHsUTUC2IyJTsi5ZFz9tEJ+
kClq4SbOR5lDG9HF0R/0I9gCuMSb+hDsdwsRE3y98a8s2GJdBiCwe9/2wxkb+IXR
LAZdEKnaBaiUizG8OO7I/F85Dh6YI7644J9LVXnCLwIeKuVPVONKnHhrDlYcgnn9
4cqxTavPjj3RgTf6wQ94ZC0p7jQ15jvzRvmtj/4rghhEPYl0qE83u1I3iehILAbX
ewv7r2YTJTvGjGfdOkWCNVGbdU0vtISqvlDXn4qMrRFrBnsWF6cSI4BapNMI8vz6
2udKVQLK8UxSMEKlAofRRUK/XkVVaci3TauBNvt8IIviErm576gzUxpHjMrOI4rW
qZD1Doe/5c/HLT5wMlUugwKXQylO3/YLwZymU17g0DyYiGp8VFYZjEW5dHGlmPpF
NdEgrigqDrtbFg7Q9mwNfQfc7qP+lY5MTiT66RYuJkF4PXO7THJ5O0r3ND8ZqcC3
N4aeZzrrU03G44e3qgCcKWgG//frAt4nh+EBHGGYMW4xXRLrjDiWUtDlVxgDuIMw
3G0zHR/tJ1mkFx0Fe9SkDqINfPa41nquhoEn8Og4pCeIMXxepTj4PyiIL1zePjbA
U52SXO/C9noCnMHjau7msR2NQj+sndwW47Htghb4/0CmA0eRNn9z7fUiN3X4MerU
ThjtPy6gk4Sk6aNCQm1t/tw0OrRLLP5vpil5AU2XtC1GSNYbhRHDeURXk5LuHS1C
kgbc2avYvf2JdSpGv9cLu0LZtoLH0Xo81e3ZlEZZV7A4+M7LjaTNjrb7Jz9lY3pv
t4YE4kuiddvYNAtnQC0cAwA6VKh/d5tU9/hLzdbpDooJZPEB5EmI37tLmmdg0whZ
tX7zkR0HZAESz5tChnYhwWY5RU2yfLw/PLAe3cn44TOVcMyh45X8LgfVQKwzKCsO
yvC7gYxEQ0tLNghxWeTf/htgEm33PeE+c/2F0Mkz/GsQycXszOrlma3L5D0C2Iar
w98wFJFE2qLVPjkbLj/RSI8hHO9ObU2MDD49125LIZywIMVvU23zGsEw8fIsOU3D
ouPCwlNzgNv3FAdEoQsmrFSbutfIPvV9kt03pgCxmKLFXSC9FvxTKGmpMwGBN02H
sTPRPJ9QJgB5NE9saGCY15odG41X5JECcAFfe7sIix2F+Rs2ETCPQexp8wAzJufG
08WOgCuq/IvXlq33dtyI2ePlAyGmgi17jtgzUnQpda3hPVnJ+yfsobBIDlSKq1b5
9rfsAZHzZcwkXoBL7YTMeAtj13ry0kjIyhbbIF39OmJ+PynTf18hOmXp1RZCgUSa
36ypxDA03KbjgImLHfRtNo2x2rko4u91Ahu5MwDfIih9b1bzJefh3Ou0xA+dZHIi
P24+HW0zvBCGn9Ikf252NirFbMxBZ7Jkc1kEPEopUfQSZbZZjsroLSGjX8IVidof
w5IZ9BaEB2fSMP/OpUMbGcRaaxxtzkUwVybmoHyYzy+V7LBGyhvuJUN7fPqxvDll
Yh3GY+1pFJ3fgDkF02Y4ZBRD4M21RIgcOtV+uC+5c6bnKBI79bL58Yb3MEVcp6An
rz/SCQkl+nEugfMgaIb6pIbMqkRt/V5FawmympG/GYoJUGpK/UuYgU/8Kijq7OPR
xHgQzMviI+rPTQZgEV6JOPtIATR3cEeezKNbQjZOcpIkjypasj+zIBL98V7WW7q7
DdRrAwAzzupw8Y/WOqNweS3/mGK0LTUY+XiiiBJelWRmk2Q3HIMU4WehUVRTLd2m
SElR42OpFt9TXA3v0Llf0922u6y233BA2fF2BM20H0jY+TasDj+dKVDwJ367KxcH
/BaIKhTppwnDt3k8HYgKJM8bhg8UZvEjjuDaIWkepUqq5nC2Pg3kZyEh/YmKHxWK
wlF8N4ncc6k/WmQcQ0buPqa4vokGmeOIQ4C8Sh2LsALNJjDnQBkmV3E/AicLwDfP
ESBw4TyNezu2ZBJto49K3lzwaX2D9Zm4NjQL7HAa1ZnYUo/pbnxB7I2DYSNZJL/W
ohK/PDI/DIJLt3nZQI1gxCBthNYqsFlhfzqCUnXW9HDwKtyDoE9hPILbG9unOf8h
6RGjWApAWlxxqDyJn9q1I6Q2n24XCIHvJJbxR7Zn5Gd6v0df8q6L54iKYVcwQfu3
USUl714QjutYMKeIcyQGWIt0EZrP9sfQ6tgBLhRe2jFsB/wkU9/vk9ohM9YZmgIF
4weBr2QKePSW2L/LAbp69hlafYYjfJ7LdAq18gQaTXXMpYXduOVCrP2iDdsKfIEs
E+yufSUeTL1aYc/wcVBSCwBUneb7Y16x839tm2fUbWsomDd7fzaNu4dw8zk/whxT
wfpQZfjGc7rf3dW59PgG75MKBZWWUX9U+pHEdTPoA396LhRVfZNQwYitpvqc0xbT
Y04LxZ4EBRQZZ+s2cnwNfoTUJ3cCYGA9Kkt1NZb0DNiypYhPjTXv/wF4mHUJCAp/
vK5BfN+xR9ApKLW5+0bnGxyA/Ic8J9S5iRj5gU2lvdJggZOp0+udW0fbL6YEgSlR
wIRBr4mGlPPzlDkhCHaG7LTHwhJewWs33yGnQ0z3qYWsZEBtPHyihpEtzG6JC4e0
VGYo8OdMmmBhmN4BhpBMXwmeCpWvXq8EpmiBvuhOvsQ55tsadKbrvP6hNaNluB17
w61idGhcY9XH16vRZjr/ZycH432HPcwYhUTw3MPAHuD+1UYYu/dmZRtJmprCUpc1
7sTXfSeojbvXsvHP3fMEKoOv5zPMFahJMNXiFtTqVYbV6oBFR+MGLCe0mk7CTBQG
pqA32y2Kyn7wDBjTsnvOYg6qcU+D53v1XM2ea9nmyply7l1q2ydCbShYBDuV4lM6
eQCAHI3EseJtuTLg7Lv5RMIHsEa2FUmWzD46wNkGbtPQi+SAKkyeP8O7D4SltTaV
i6F4IP7pTAWqNs3FM0bYRamCW3+8xHzvAGSp/KYKP1RK72TLJtrtiteHkfgiJFlD
himfEtXXD3bCDudQe8CGpmMZrdA7cq8JexKT7qZuvDNb0T16HB8bTDhRhs57L9fo
9ZpjUhPFNMCfuvQD1rRTfF5pcoMW59b9GvBQ9lLLN24f9qtrGyZbobaAYOWQLvJn
HKeI7fgzSU8pNZcgzsS5S7FSWyn+4icD5/RnfKAsRKP8PBNWG/gMlXImnua5HOXM
vbPRQCGGvOdBDpw11FxCpTDH7Va5SlTGWh/KCCsQz69lRoxPZ621RuEQ45nhxdyK
oYzScOkhTC7oOXRCW0brEieljJ7ksGMi76YJmczq7sAYq6+NbEFGo3SdYZSc9Oz6
nnwuQHqSBJ5AvOnWDOtq5Jshvg01jyzML905l89I5cGbhSECyLJ0pPfDmGehtszM
6neeefXwSzxRWT7Dm8dvnRWO3ff3E4XWo5u/GDh9aczH58vxUeSzZyjce4WdF0UW
GZ7WtkWHSvbowVzbchDpDpW6/CyMPwq3GhLgYhG/3hCeIGCL8tYyNLgRgcMly65X
TOUNQeM/P9MRwX6ZcGqW1hFhUITIECRCL7LdzZWhN4QGmiUgWs5UQJnium+Jedca
L03M1gWCYWF7YMjAMv+2VY2OjANm4Ese7r4CVyaGi0qVrLmUIl1dvD4KhJ7w/Ptj
GqQsmRJ75s1FA0/6u3oboT9mWOr4pg2BDq7b1w3/O6uHhylv6JfltJ9M2FLmtM9d
JjTBvK7tBh9wwzj+qJI0DXeQJp1hLcg1tjCPngn/M7MSRu40k4t/HfVPLUHe2v00
rY20KW0edL+nsD2b5H37QzkYT4xsBPKzYnWYQEmjBtTiNdSHeg5GhIv+2AAnyVYL
mQkKYp5Z5ihZNaQMXrWbvw==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cNnvMG+cEZy+u2QJryu2oO1HIAI7n8f31CqfRb4Ve51pOkviAp0u0+twJMfCx2oT
OsbspcXj2eDUMg+pwoo1hWMiEqdL3Td6JkhPYFhd4WrykgPJw+LkYGLkq6NXq4cI
Tu6P8X6iq9+NCdrppaUbJdXNmBLkDKq0M+nDS3pLNxusAXrU4vV12BAAlYytNWBd
P/tnsqUELo7lbMz5AFPswDHhmu9fGWOiqFIc2Iwf3Y6olI3WoIdU66ht1NUV1GBF
7TIIHfMxdI7pNEa5HzCPS7dZWHOHWwUibi0FKWoRZyBg9su0fGSmDe48WGO7yH4j
zczL6vmIAuDvPmuervsWcA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2224 )
`pragma protect data_block
own7auQSntetEtLwbDu8In/hLCBwk3KIAp46X5CGjf8MooKcwHN/U0XFDjoT7adT
IpV7NMXmSHnlsOPBnuN+dtwbQQl5uzx56+lSKEmcMqGaVWFa9Yikz0+uNhiTWYWK
2LDkv3Nvtr6rZXx6wI4Asa+62N4TYjg+DguyZLYivNrmY+nUSjyvA4+B7PGdUjQ2
+bjxvSktL0PNP45WoVzOOGSsDvraAdSvah6cTugqsCo+/v2e4O+YMaqfe5fA512g
OyEWJFZftjaSjVUAGfZ7J2ni4Ld4F7/mlD3vTaZ/DjEinNL1UD8N9F3WEHcgPXvl
/ZDWdlRJrEVf3FNnvtWBE2cqbzT79hLRvaN9v2JLEpLGEhzn5Q6DC07aEK+itzJS
ua1Dc3p4dR/rxuZvj67tfskQ0ZNHoeNnvMiL02GwGHubBP6g/rpyR8TqHTRor1vb
NZ3+RTVs6/xomOBwYKirEMskeuNSkshs1BGH8jxtLXtdMrJbnThRS8Q7v3s0HJfr
gsVST+hTNE9FFwodVYfC9ls12hmt8eP7moSi4osEC6r0ZOH6KctARxPz46GGHhXW
Vbbqern23QSA9WlfUWhUx+5CIdCtTtMSCinyttGrKgnC0tDtUSMInP+0QT8WMQUO
AwVyGt2CWic/iVYXMEdVK3VgFM40ow2tY98eZ7hoTPaR6wFyUFR5ZgEuig1sSbFK
NFAWXk97eDDgdTbEeas6s5OuoY7QRKJ9cqv9EZMhT8ZKS8D739Yiok2O75J7iLU/
r/r0lCABre2vZb2a7VjoZKFmX1dGxCN5Hoawij8iX02yCUvkauvOiPGNudf0Kk/V
TxX0lyBe3KiMbwiBAFpPW2E2nn5wIsnGBTjlsh2baKqJd7R6tVTGpU++TIBtPURP
rMf9Sph9fkXaFnuQzpPthNc932wECga4RobQzjGc5VjM9j8jXQtBeNzxQ6f7Y2vR
+N0eNWBI2hLTA/n/TQrwd9Q/jew1Wnz2OB9KKnuiD+fjmAm8BU0hAtOmjFNuCORf
dy0Z6Egqk2p+gHd+p5ZvzgWZWIK5wPhU9w2SYSCUhZ9at/PZMk3rBvx1sR0rgouE
lkFRKnTafebcjCdEDxqDiSVDf1d5vCqJngHhbEX7R/2AOIVtkNQZEX8w7OZEyhkv
f2sMJx1wMX2Bq4HIhjnBi/ZqOG0jWzE6uGP2Zb2JASrqXTX92/T1CpBUKg9QNuIK
RI2Hz2RRpu2VyR7ToSxhohvAGRFg9QTHaVSjpdwE677KhQsZhb4uJaYrdy3BzQ8v
wMYohfjTnBJi3ptPDGbocAwtlr0I8zF21dkAnWWSa4esBZxc0+qx7hO+jyJfN4Nr
xietwFkcCA4bzXucRNryjW6A0odM/1pyydAE3yB5hn/gbaz9UTU8G5dZpKnG0gTF
YGTydsjxdrBXeQDKXR0Wh44ILCKCDEXOmstD5wYP5F9J3TWwqK+gebWfN7Wc4RCe
C4KlbXyEXLeFIcplGRE2BqlCpA6GsJ+vifOv74cP9bEOkvCb1AaJNBVkEAnDvuDO
NNy/U+MHX0vask9mgp8Ol3khiHSDCPCTuzUEBjxPWg3dEw1KEvAhcEfEiS1NGIIZ
npXTKcr6YlmjDxSWOBFiykSHwNiHEwZR2JCjAO2XuepS3HqDwOGdC3SP1Hd0Kq2K
u2hFpcsVjDBddt0tctCcN0emRVWaGyje1/qCsaz5x12BttI3PBshHkttXwvi9Ufo
8NEBwMO0J7/BPP9IR9LcfBqnSyYImxQyF/0jvtsJhbr4oDlAovLijj03pIj2DJ7+
oZ6Bi/EvPXiocgU5AbbcWo/x+JBy6fj4RO/yOsWNdRj+wzAX/j+wExZzOc95TeVE
DUD1Qger4LHzLEhaAF3aPiKOAY0q9rWC2fO7jTPYH6CK3YUlXPeBGMgSmRescP8q
+x9mJsnEqrnoFRLhpM9CnvS9NM0w2V4q1DkXbYWbbDKxNp8nG+q5OtZpOAeCIPsp
6rEJXAzyJ8n03sNpqWqT2511QUAotGWRnAu+OGp91bDooFZey82Q4WGLDhvw4+ck
YAuUtVftc032wPax3F1lh4iL1p/8n21/9pMrgeiEPbFbCd+G5RDxC0spOJ1hJ1Ec
I2yhCbh+sLuQdcjm4RqHvP819s3yy78jRQW9DsD443/gDcjL8mVOsK/F4qhvOEtn
5SJ8zRb4pa0xdvVGGxxgF8tp6tRkctpXOYV+awjdsNaBSzS/qEgCcx4XcfwEXBfo
FMkJj9p7ZDcQAa8xaL/mZ/+9Su0/H0mS7dNThBK/PRdEvb41M5Uyc7abv0wsb5RT
gLZFfZ5uhJ9CFay0Ox5l7nroqUn+Atwcm7rQc0U1tJtI1wl6IgFBb8/SQkacyWLc
HPMapgX8b19ssnQtEntiknfMCXf9H5gIet4ckh3BEDIvkWE2tx9854Zl8O/cqLof
GmGuDT1xgUOdaPR7vxZNdHgfcTvcH3kqDF+eXJH2CUqFjPI/DJdriXx6wkfAjftm
8R6ZResTypmhtH/A1haUq8vNI7PA7ulqmvsIqNXh0/3IpJPtA3BH7kCSgx9a9x3K
0ZhxZA6iwRZN/P0CCITLOoXPgRva+4bg6EYbm41I/bR3pO6aV8mNMlkTb1fRPRe/
w5BdQnQA7ODjf12ApCS4vC7z1SfOoYm8m5fsrMSBhWjwIuk+HOdkDPbRAR6mMx5U
hmLGzGTCfR80Vrgr5BOvUJxiDnIWWZw1Xo6Y3C3zrjIdj28bNDP9ftxZFRpqvpYu
AQ0IbMB+HBDvEGM6z0wQrHbM0bbb7oj0sT75yh8AuOLPpuf4IcuNKxKPOHbQzlfJ
r7ZqTGLGgYHDJ2x3Akn0MdMr4b5IPx+mWygI80gtiqmi2sG4/tiL/qV/1yAnUT5n
+jkkhiaEG4T/ltzF9C+KDFK0O6eVH39swpAz7FyU4jHi4KSEt1zS6wrbWOQ2PZtg
kn9luL2nyZ3ZtF6mhhLvcw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gHSohx61XG+m0ejvP1IXd+s9otheu9zsjfDSKckoyygNk+ivWYebgFnOKosYrtkv
NETy+q6AYcu9Te4zhcJEGKqXiMR9qAsFAxujyzifwQYD4ExbcsaJCTLI4dgfdYyf
gceIh1uDkigEXvSmSxiO6QAENwRXoqYrcdqm6mUm6Irr0a8pIfsLx1A05GEOTMrT
83QZTMmOGUhR06YmugG29piaUSESNq7EJZiO/krNm5OxHS9dyZ6aD+XpbAJz1KjY
K9xSKhWU2YFSf7pyX0H3eY/JV9FqjBDRzOQFoTk6Tq76UHxmRvVKCEN8TWctmEBI
SqlFLOjyObch1e9Hcu2oIw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9328 )
`pragma protect data_block
Zk46RrUQZY/dub7qdf34N/PTsLWRV9W94+JQhXYLm3JiHck/eaTY1+CIXO7MyipV
223zvwSinNyM/Mb+9plA5OWOU5YNPBL/DfO3PCNc3wo5Ro3Ooy/HZPg/58datH1p
5JITlBlDwOT9EfxXxGePEUiGXrdISz4TbTdVqf+YW6Z/Dp4JfMkoAiIsVedw+sfF
uKsfl6wFBROMA9SgcL/xhurN2WWzIlClU4qO4lQjJ5vEjfvLTLrFp/6BrHKyQKAm
PDcwQvwqS/foIIB7+ivk0yrUbBVgfFg1sqptmdUSSw57QhUYGTC1M01Xyzmnmiv/
3R0qSOG0/5t7C6pCTA1wBJDqtvWL8WobXN4QbEs5xL9QVtzXGdpmrTnahW/cl9E+
cL9zJpxSUti2ts2FUJTzBHCztJ1ZOtv11wXVR7/SeZB7mRqheVJu6Bh1odr7vGqI
QInK9okGSInhNAIlSWwow/beSIklGD1tvwCKupMxJO5DZEbUaQorbjyMgmCcX0xp
7SDMBjH6a4/BvG956UHgVS7tQEV9byWfU46QSY71Vhe6fWKD2ffwW1r1BcN4MMqP
WDJD5RuGHaBsyEciRrSmThWMhbLc4Jmq3uSrQTEYPtiJynV48o1Z2ef6IcXtQP04
9IAHYVpYR3JglsdqFAjHi9rOzAkm7L/a+xyfv7iMHIDy/vtbUhQYsubp130sce6z
DafEprt3o+xRwIUZvsEhR7LQSF3ErLEYaqU1shHgl0fld6kWYMyfxiNRU47kHJij
bpYxBS2tCjzGSsuRZGhPN8NjWZ9ozt941p5KZ35aOx9jNw5T2F7RSDGzlE33JO//
dldrTeVe/l+OKoaM3EMnr+gmay5xpeNIXIDd9jAX55kHK4doBm9An7is7kb6kcm7
1UyQJ+kISFY1PQaXKW7L2YFl0qEJwB64PunstT1/7bBvKa1No6F26pH90CuZBvV8
uFGt4PSysmPAF0mAtgxHKdICxIQvdo24BGFQ+ymSL5ggQRQhZF0pjAseyGSo2eRk
Kb2+WMuwBBZTVQmN3e0nH3eKIyKlda8ecoqSC2PZz4cfpe4C+ojItKaOSjLVvKDO
SI42WxepbjK+zHMJv5dYAgGLIOilNdnYKR7+hvUvCX+m//gedj4vWcBqw8Y4/YM1
NxBQzzK0ZwYz4pBdHa6PSwPDuOr/DstBWwOPosQwk2vHUrg1+Bzr4t8IC7QDtf1r
dGpQ67cs3z5TUeKgqHgqU1JrrqK4f1kCKSLMw0adUMIgR1UfrYVCe79WHYIbp3Vp
dMDaDw7k2OxZikJUvyhKzWY3LZ/bMFFenavJLCop4DxgClFhCQgnfbbVtowqO327
kDiRNfVm9Xu+4lQ50Kd0FBFercoPe6kN5iuMdb5o3Z8wRWT1VHopDbLZbiePnHyW
FPJxqfrheeKuF9PCI+TEmTF08Ngb9AdmoqBBnB320VxQnOpoKe7jlDY0a9bkxKEL
41c0JyhnikeYf26GaNsoJuxiLhw48eAPN3RK0FajyyeROBZGzf8ZgpRkwtNrrWrE
hnULke8YaEmDvDW3T1wqS+4UGM4+KrdD4L7nL/4yKoiCc/FnIkHmkv7aci94985P
j2H7G0+bYMZ1Ww/6dVruqmrmTbgOJEZgY3hfp0HATqn6/+pRrN3lSp10+wDIFEkJ
678AJiNYGC7POeaql4sc/NNyJnAASxcx9X1IpvS6BLfjYsHMACW6QbKIVQJ96Hqs
7jAuiYWdycdC3xM69ySrzVFgPz1Spi13pfM5SFnkAzBsqG9IE7iYEqej0z/8zkHV
z9jWey68wPp+N5uUaLfgO1KubuME7sg3YrD/v7i/6WaJXtlTqBND9aZU8q7DVnHi
kW5FOkKkw0lcbLBdacpVF86K+Qhj+w/Qkw4Soe5Oa0YOXKfHNl4djgNqD3axNCz1
yHs7LrR4a5lls9dASi3Pw8tCXzkwu47ZaVhrE3Vcr9SZK1wjUS1JPjZ7D4Y0XKTv
S6TM2mrW13knyO1K2S9gnq82aopzR9MAbPhLJgcLxDEZiFsoAfNqiLF4k2yKW8zo
qwX3epe7ppFoEyLSZF1LlvRCl5tEDBVowvdF/1i0EHMgzFju1p6UETLmU3wFO3PQ
c2LJd9Lv2u8qFOBepqfftil3dWi5/x5LAOt0jHvaDXnbnTMaX2AwOMdeeMbHQYbH
QONOaejwgCwrtJn6KC4FeZ1UyLKZYGx8AOggLjnNSAijPxXRTuPCfw7ZP7AE1FNL
ssH72vQAUYPbA7VlOtyHe5ym9mo8EoRJ5kCpeNCgtiqSpciIDxOB3SikjMynf1lh
70u6sbYOmuZAdTQWnDizcTO2oFiauCHP0UKkb8F2iEil3cS0Us6vbHAhbngycezq
O+bHYbi0U+DwFeBQGZAswv+VO8tqk/v5W8/yeWTmait58CztPOQZKsl03pQU9Q5q
pXK46PgqASlLG6LYBaR1fvwHtwy9j5329kV/FPVSpTzeWontlQfLoq+nX0FMD2rw
/1ClN0WlJMrR6A1ogh4IZhH1aYcTJV0Ty82FwjNcxVag+14caZaMhI2WDu0yRYGp
imzcuHBpG/VzpOUAatAiaI4fj0dKFOXISRT5kJxa4zvjJWMotD0eNdoUfX8JlxvS
qI/qBW7UzFYPT52hpvGzPnCDzXMMH3CEQ6pe10ErE5TL96zn71lcfmKHkhLr4f9o
Rl2nm4WTwH1EXh/W7tQ2kqjKNVRDHz3qH2kAMUHX+sWE4vXZKkqacfxI2J9XfW2R
8OgEnLXdjfrk7JE9SPlUWUEIS7E/HI939N4baDVDXZVelyMeUmmpzuBfkiPSrIT7
gNiEfBpKl75vc+BY54cdt8JxalEAgQfP2lt8CDs9KEfPt87CI6nSf62hcIA84wC4
3Ni1MvV/B4hu7vjTHIvWGRlXOFGkCPh+01DnBl7OcXY6AWXx40jGXI5S8UH6L6vZ
Mx56bw+Mi1lD53wDF6SlnQ9PLKsQxNCbPFN0ixzhr2KSAM7mjqjIYtZBEasuayZt
P3ei4ndaZuS00VMZAIkkBoLp4OGDbenuHgiML5P9vhpwGfAZ3OVx4f1xFMlmbh/W
kzBvemmd9uZ3n8vJD/Qh18G3vRCnifEAlH1MWH/XNKgtNgnT3duQCSo7U9I57ugR
IfnzdlgDigf2F0vhOeVbeEnFj/gqkSVggLiwSSfD9eyUvpTwLgUI1z9Ie5iYxEEp
DlMA5075m5RoYYJ2uyvlNOXQQdxuoqyk6KHSv8w2TS/ueV3FhjjIxfMYLCxZPpHJ
F3S843JfTTSPyaDgCB82B/8iflT8hx8tCl+xSNi2KA89LJlZJzb5d+mz+I3aaDjb
3ju538v0tgH3bY3yHbStgH+VnZub9sWgotsb+YTjvxfQz2lOFEDb1UfB8OX/gWmB
fL2e7qKicNjPHkLKvuz9oR3DBtUnLhKgiv4np7pQPkPkvieOkc3GLzn1AOB5gNL+
1KOh3PwBWOaqiwGQPoBfQarOu6sn1bUj4HitGPB5iGdQ+GtnzwX4b0zL0yvD/tx1
rtC6f8spjCrJnKPESZU7iT8PqSZtJLkC2u6GOKCpu21Egis2fM81U7b66qgpGR0z
sShar+bCclx6A9fCiUcAMjjs2GQpq71t9oCO8xEzINLHt7A5g+08cA/PP/Gmi95+
rBu7dcmD9agZoGA1vm+K/DA8CkNzJ8+iGHB7fBJ1JnkaHhUn4IEWtgXnVPCU83td
nJKLOs5GXWOW74XOHmtkBh0EtV548dTk7lqY7W4kkGdZqLBzyncwaDYRRNBt64wZ
dnVI7V6B/MEbooRMW+t+DG18yNJkOtaVEOqo3frH8Y76920PGctrU6Fk26e1tV0U
vXkp2fuch/wBBRipsLbRktgDQlAfeqBZxOr09OZdNgsXUcFufXgj1sApei1qwcom
HmNoLUvq/C7mvgwWU+i0MRnuZ8l1WZKSZNyeFoVlcoqgboO256B6l25oVIjPfKwB
KSYkT+YhR1ltWI2e820Esh3Dj0a22YoXmHMeHWTplNwjPq5rdXwD2AkUDd4uS1gW
FkRf/Y8yF+vbucRf5LXar7ZQRa12u4TU/P4hp/erz7xX8spg4lzsPRsR/jqqpPC9
Xkv1dtu39Np9MFZQRHqSTySfi8rhrBWd5KDmaca8Pi5GGxIIaHXkbmpzBhPzc/iU
iJWQvYSIuQhepqpzSDV4PQ5KAi3R8pBuZrITs917fllJKrvGhQPBeyxR6NMMF3Ot
UICXi+hr4gP4NxZKq2e5omVhT0oHg2IuAlv0PcJ8UgaBOdv2KgcKvSagT2+eBZlq
uTLAFE0t5ceZ24d9+h2C7Hx6fFpmG7FoWnf9+u0VB16E+PNd/f+5gEInocvLWXcP
4xvHmkbdNKf87miAvvGyYs8CtqryF0vnX9A0QgSCIBgp8IaQhTbDQuN0LbOLqqSf
oRngi44wWrK9UyrwS9hMZEdqVVZhJsuOowQ35UW5/6DBUd9t43fwyYSubrzMTPUN
LTaK3dgwTCJkPn3HeArmxye1fYGil04Nk3UAvLuj4CYgaVuf+ZtljnFExglOHkhA
CzxWErQcjJYNODC6bC/WaFyR/17Txz4Ksakvzy26jtULPUPuyu1Urej0qgHnwzf2
s/pSuVzGlr/xD5dSECU3I61k7/3y9GLEJ+LNmmdykMSdhwFxkka+GWYWGd7I1P7b
p8cvo4Th5EKkkYue+ZTvGYURDXsRtRx4ksxmtRFlhR8Sql0DWNsHANAEAyhRCHl6
zCW5vYjf+KlmB7S/APRizGFchJYBUTrx2CJ6/i10N6FUAv+PgUx/pBC0umspsmAU
YM2VXWNr9ZuHjnF4Nyjk7yAZ/B6ryFRvTKH4EgtZXbUu5bpHZe1HYxREoc6438AU
1Os+23MKTk/vUqRCWc2rWYuwJnmdC+0Ful5x1ThCob0LgcBgSRKV01ABwiviUj2z
NFmwUldYlR/ngSAbipb/umUwqgKxsOjMNoPVpg35IaG+inzWBh6cWvYAT/R7xZin
uT9fHClVjqm0T2S+aEQbLVm2mU8n1+YSRly7CY5qPIo4/ULIyausZSE3C9RdchJm
GiKCCJdkwtfGPdCm0wc944QOUnR3vpizdtNrQYLycQ2OWwfKkVf3OgNdJGGOndgr
TvK8c64VhAwA5LmcPOgXBuoVHq3qPCf3pmXdwkMypbzB7fXPspv/VtEKoNBOWJZj
6LM3SjK/iL29pVD5Q0gIvih+C7T2tcWBI3YwxLK9JXUD/TJbfoMkUt7/d0mS76aP
1h3X6MKxhY4zWnWoAsEbEIXLXO9jJEibqWXBljiqqij9Mbpupavi791MQeD36MBW
faF6FCcJw0fzqdkp5xbkKRmUxGHVwzKrhhc5l+Ls6K+hj6WveuuEffYQlzc2TWR+
917Q3lbbLmDgbppVLYCfb2DI7pqOoXvHV5nod81iuIbmzA2T6kZ/QWz7613aIw9a
uL0EY6SLGriNLGEpWc7pr52aNNXm4eVo/XOggqZw3X7hJFK9RC5RO+GxqavaiZhQ
pCWElnjDbsL3kAtI2u4lfIjJZ41qLy2esV/Ia4daD79cVeI7wntiZbttRJ9/+oHU
cxlx8Fgp/YVzJv0ASSHPd1HT7Blsh8l02275KSeCyT/jb7lfjvje4Din+ziMKcYL
yL8Ix+hKivSm86j0FBGVEkx1ruGssA3P157zpc/rbSlMYrC1dFaKR4XwCWBtTuom
oVTIzcVljNsTGAxQo3LVqItnWAG/MSr8cgTYLmzh6mWIh/JRjSohnNkYUsli6vKK
88QgxtzuA4gozB6vlAUGzM8a1KrW0085eRtd8Guk3RaYPqSbzSbdtZRfN/kLWe8J
6QV7Ejpx07GkMZrHsJ0O2b0CJ0gmrBu892ZLATrtvzuS9zMaPCzNV2lrTUhwVjTf
AbhWBq/MKNs/EsHavcKXrF1zTdd9ZYZHZOuOUX5X7wNvvDXLEJu6lQ0JVQrXVMx0
a+CRg01U4px+kFuH89ikUlBo2esO948NBgicXxAvh5JpzByd9t1RXOTVWyTjNgMr
QEBj5rWxQSgr5N66FrCeLFlzLTIgwdAldixPjVG0pzFE2O/EXknID9fqDIUkrZeA
RXlZVFlF7bJE2qOn7AxoBW6gFVASu0cwxsbJAVoS304GQi2KlRwpKKKbRVb79tBf
sz6zf/S7+/+GMQ7T3sFrwbxDhRf424YQUJ4r28R8JOZguHcS7sr7pSIaw0pkRAsM
mxpEgTBWLUilRpXPS7UsaAdVsx3JpHBZK/BJnVH5F1Mhw6TZKzut5MthEBbSdnbX
IxRLCpgwVb4kwvx3r54LO/ONEMNbRVlV7ewBKjcUNHBwNb0l7U0paOLZMlQY58/d
SIMOBAzvzsTYYzsjBZ+W/wCkVuOVzqdCzzRwVAb8FVqzj9iaJ1zbVChHO6c1cMZ0
ufiwaehTe175HXKiY7wm9c47cHieHb9+jPnVRi74E0CY9wqKiFtDpQd9ksIOOmYA
2ZC9NucRzoqGGq2l/PdE94FDUf7SmofLqKl54SA4SjSBU34GXyAxOm8M/NT5cxES
D8LqW+5YOojpnhC4CwedqS9y1sHcG/OHMlWreHz3D/dbNaXdo4fcY1PoihO/YbXY
kG88whiZTIBpS+LDv9AX86vWgCo9WP5Fy7eCeOpSAIQb359DGL/sIxfTEGAPRiGe
rUHeNv30MX0xgowJn41xOPCYcyeklIThr6QbgY74pKZMb8awFMThzrulxwJxmqYf
JmCjszdlst/oNfNLQX8K58WDwjsjLTAXI4ilwbln+4E43iqC11jox4RziNZTnxAp
gr/+CiLAMr9XQCVVOtYYXdnRteE7mY8iZEylTnao6kYI+4G0/0IizLTenZOmU4nM
cNIoWBqQG5JKvuDioj9VcGpQhJpb57McQz4Vs/3rZ26foR1uMzTn3y6DympxCrvI
/XdyJgxpt9XvJ57vBjKIMOthZRdn3rWyGOJ8aKtjH2AvmcQ+2+9iylnSc9+yrgDy
OYEvQVMHPeMDPXOm5v3u6a1xwkAxAS4f31B4lrkXE/TCPowmF+PgNyMmoRpB44nN
ZV+XwYlI88DehLYWRlesWEI2pvhnx/lwCvyfBiAv8UYxF+LOlu+aOcKHhlVqOEWt
S8rVbcyVhvWa3Pesv+kRagZA+4eV0B+daZBbFWqPtura0QRx6ciT1Pt3/FbRmlq8
FfNpUbo+ZOHOZjoe80Ghko8qBsxkSVHSRyGuzWzbMpAJEc/YCGOc7EalzxzHIwiG
aiFfO6vz+FLxTAgSubvJ/R1CJT44VA8UnehoiCX9L6VNzmf6Wye07ctu1n1vbdfl
5a9H6tuoqv+HNRE0633IvbNTbzEe1yJOBTZAZeOfYXQ6j2obIRAPn0EsfHAyXFRP
b0xG8plPewGykY2zo9vKhiR3Y2JUTrgcw5cLWpJ/dK7s5rtn2wP1ap5AKJqIdQmt
bMF+wk+/93o+MPeSZ4OBKg2sh/ELi/quG1+7TAp5siuTdHYSHHWgmMl1EyvBa0AE
ObVedX7wVU4PDOEwj0JLSftdz/Op7kmP2FNl/96j1EtDfl1q9v5hnTw+XgH/z0fK
zdl8o3B3evPdzllQ/E+7ubrirRYJBm6C7F4pszaMsnV53dcBK8hTO9zd/8/WgxeT
TPB/KooWXPdSHFoUdQHa4TUml1bPCq/QCcbjTdiqP50i+IaS1p58iTPWhPmCQBvI
Pymh508OeBJvjRP8znp2bYFhtKyCUzpHfZYozwqS5Lxm++PgOtrWpmFglO6TO8RB
PQKNASwNgSZnwOCYlOJEHZr4dP7emHDO4wafcUYkgCHHw6bCCLCtQS2XTUs7ODzO
EdXcLTZ2nzm78gZfy6V+D2q7XQYKG2KxIY6ADyhD5+Yy3ySfqcz7Rqb78CcEInaB
rNOV3lNgo+dO7paxiRqR4WOs6PN5q+5v82YFPF6FoYoFnHvs3qzuC390iN1+6shd
z0sEPPI/BZtxUvouPbwRjAc1b2rIIwhA/yPC2Jnr2PQrmiOL4WUdGPO9qzefP6yF
9lmC/OZETXoQr+f2Ff5NPnIZLQl/KoqIZ8hbO4Q88KEEYwk5cHIQWwBfF5uuW7qg
d2+p741KLiAeUB+mzSxpnsJGUFlYLmcu/NILl1aZYsIVgz0mLAku/eM4RUBwVUBb
JoFrs9zWgY/BDbRK109r0iTqTbvRhqvrWhwi0FikoW8u/YAiCeDP6LG/+kkm4LF6
VqUTo6VveoaoY+AErAfMTBxSayaC6to3l1DFb6FR9YphhHJH875NSxiZzU2YpYLB
8YE6HF10WawtyXZuuWxiGq5AKx4ricXvGluGDiPcsc8JQFLn/iT54UCe6TgI5YXJ
1wXmMuENuB0ZTtwgQaKLVysQvQMgJ567CiJ82E049H25P5eKeTe7M1cd3UwkkcaI
PA7CBj8PfplTNw8toU96R7NiESB/7yEJ1/VEqOBsQFckwK7/fjuaefvlWAW5ZG9j
AXxPBYms45w7gS7WwjDAFPUM7bl4i/+eAv1kFbFUq64H8/dCFy2CamFOJfcgCQJz
3Svb5wT7x1aTAG8FtXxQrHRK8n5SIMCU4SEc9f0eH/lls4PCWJhwOoDZs6cHR1eF
iV/hajg3HY8cIF6FjjSwD1pGX+Gonc5I9sHNLrPpX7XoW72aqH+QtB4MU/desjxS
1WgCBxAfQxptuW886afhEXw23bS2uXvJwhBlvdsMFqk7DG1ouErEKx+xgD/CWGKI
4W2G3yyrPkmPwrUw5lrTEnjcxo2bGcaYmKYD9pK3u2B8jVvYX6c3MvPxPFWDQYR6
CJYC831qI4MUjwGmhoV3Ot2rnZAnh2bk4GnmJ1EE5Vag1GNeWgh6j3fJcage3qBj
sFnlFkQ2glabTU4U9BfhLfMebdsDMfnEIM5KaTKAISsgKmCQzuylEKjiKmgX3l+x
q2NUvf5ScH8Rvsao4zKvYtgaw7OeVZqBc1CF4eECpJL70EZ7n9DKEpCETjurxGEn
a7p+tKzlPcomE1oPhUiXJVv5oo261rUiGEAIgvsdujk7cHx0PCKe9lw9nLJd9LJu
mr6C3C+fFmQ+E0uYNo4bOtcjvJp/um+mBhRofMh62RQ0fk7driy5Dnxf41QMHNAv
hvUgOmYgOw5sUhwl09uJ8Bvagh2niFLvi42IAVx1FybfiqivMTE9qD/i3jZiICPZ
r1rwNWtN/Fwz5G2wPXhOk1XDGROWE24dlwS9hiRrHQZ90Vo+2FQW9fW9f/xYNUJM
FfQFnujFSXtRrAlCXZuY5R7j2JBAw8OAr031lAHBRTnr99yOBlJyI6PYsNjCI2E3
M1/So/QYmHD2RJsinefK+mGzhYzt2htk7fslnXgmE7BkG9/KI5pSE6EC0e6bhWgL
nEhTpEz7tZXcK7UxM8CltV9E7y9LylExIYyVLejwQrtPK+3zXG03Y747Fn1MT92Z
J+uqCD8JYqAJmM0DFUXiPr3p1L8VWA+z8rATS9PkDUeFu6ODGlRmosHPUCM6dqG9
3rGdcx419dFiFMBFR4LK3CBQDKQeXKjukykqA1XcaHn1YnFPuHukxVhrBgCrjbRz
RWnZhy/bLd/sj+YL7bWztcEdi2xXckP7AWldG2PittRhjmyMxAByVqWDhkeOdtsJ
9ifOKFOOA3Bt6ELwH2bEN6k2W3Dph/0ar+qO19Vl2PIUGgkAhuy1pFtxqqv8KVbS
bEM7WFcB4f1AB50bI1EtOHYX4ruE9FRx2FyaK7qzeEgwLLutd08Nw4M6K0zOqfwM
ubGPYcTaPIVzYZS23mYRMDSfMTeZvDsRqgQgyEg5teRTZDorlBSJ7KSJTa3KWVju
O2JMeiTh6kz72r0tka9hBGBKuVb+Soiu6sduqwAHnLXB2qM4TewlM8roIEH7IDuZ
7QvBPG4zng8YM+4+3Uxev9VqChcgJYcpRPuh1ta3PA8JvDz38LpYfoLd/WnJZuWZ
/vSH0+cUBCD4KzMD7GrQhoufuu17SOaO0xzavDdVZy5yeh410yGwSaTRc9vy5zBi
0RZ7huTquDaNuViBeiXTcg74xuxbiJPOWbGjDu3Vxd1hk+3wo3pjiJIVu77aS+/g
Igyf+e8feOXRLrRCK48o540h9L2dRlxm0pN/+hJIcqEN+R8PTLKzvn5epMjSmA3N
G5Tmdd/N9cv/D0fqbGQXXj035iLxrimmHPtlHyoJEZYRJV9wCi907eylabPqyJCt
rPbIc8Z50pteq7bQOa1hnu1/s23BFnWIyMyhueNdS4dQqBTGU+DwF+Eeyc0GkLi7
B5MPtUhV6DQjXg3eJt4jgOCklu0z+8t+L0GSgrA021CgWHpERyNlyOyULmyCJ/I/
aoJD9HOFp8vSb0pZQy3fuHvewNmm2ARONkF2yum6zTG1wI9urAS6Gtrvz46Uw94V
VNdhop/hPT9KtmOqvxIz02RncA7udSH+h4lqQTLXjtVJem4FqtYFoAYZ8N+ViU94
es/eOmzhnEBFNGtYstI01Zop/peCc3eQ1lUWEQazPTpAnW8OSmj+LM2p1DVZLl9Z
j7k6OXoQmn45Y0Ok4AgyNEHSjTlD9dOmVyOxwgi/8Fzqd7DyNnz2g3lYbuZF5sxF
PzsWyrS67shL2vzaeMGB+tM6Sq3TxaylADyJmwns9/gQj3ZLsDFiqmlbYjld/tL2
9PpEOVFTZoIzfla5ccB8OB512XCBylehx9zECSmP9l8m5LmG4x9DksoRtUMjk1V8
EueC9an15B3g/AcVI5O8EatK20j1B1i9GADE4v17rnsVhy+fx23Tc0IeaeFzj5ZR
MfwHnElAoDoSr9jaB5kKxbJUl/CDSNdLNTP2zvkJJ9wwD2VPe1Y+W1BEfRpJKsbf
Jv0Fpz9dWmxFBgk1i3ZKw9jmDP8jk4qwv8+ThNozGgEdaQcBCRXh7cdEwBRkBqrm
d0K/suhSqragoTnpGyBv/DECnjcylFYR2itR4s4QC6JQqh/qwAJqS7BHBFWM1XXO
Y2qkGLcsVYQUYAUpfNhJ77Gy+FGL1Dxr3PrRxw+LKD3dauLwLADx5IYdgAYbKqI6
BLCJ9fVKTEne3T51fq8vtqCIg1X2Use0YeaOF/AaLxfEbb+7kqJc5YdCs7/PnlUx
7OiieVzK5TUhnQavqoAKrkXTAXjd6JlpTXtCtUU8V+UUQ9Cu2TdBtcAQAZm6Nyis
USYJ80XaMfVw4f/rsu23wGdnE4NIJpGMgrkkVoCAGInj0m3Szkrb0T5epktpvB3a
J00bZQYWI33WVQchwpWaBrCFyUOU8nk2dzQJl/Oh6eePbeBuXQ0MoippoxwtMpvQ
KuSobvg6LcMixwxhD3jZvgmHZtvOp6EIEJC6R3FKl5xxEGnPjy/W+gzgJnDR7hFo
3k6TxDTqkvNRT9OHFgsuJ1hs6Fp1/nrmHbbMrV6vK3BSqe8eSrWy1e9Twq4/sx+N
uP8uZyJjBXLEqbtGzxgB0fS4gfHXs6wis+nXw8Zckh5hXTsEsfcOoFcuaIhjoOrt
+YlT4+AoBygB+tjKQNixuCL6nFy9tr/JPXfu4GoYnSb6hD98LjzeDhIi3PAZ/vfF
ByD7CASjiwlY0fPH2lgTkZ8hQwOyjiSHIWnTXVBM5t4NI49HYTJVnNDatYpDYAXk
9zfkT+uMLMm7CFctBF4s4HuSmMtCTyj9RW7kbGASRwRjaE2Sr9Zxx8L9hVmiEWBb
Osjpxaep4Qufsl7SF51bKf+5VxBcaeCs1JqskePwwJA5r0+HkTiTQvwkfKW0K4Wb
VV3dUfYpPy7+DJcRcWzi7YJR++GUGb4hQFpC4EflE6/RHjASogrtd7fA9kojfQ+1
srVwFBHGfjG5qy5+kyYGjVd47yvjInbwT8G47zP5kNJC12MXX3+Kd2+Z7H9svfpN
TuaJWJmvDcBQg7Ud82NfBKhXaE9qFSzX23kmEMDiprdOSjHdH9/rH00iWcjmo/uH
IpjIyF5n6Ydoxf0VdwKwLiWkbO6JDiybSA9MsX1eGRyVpUbQP7w60yfmGmEIInP8
akEDuyAUwnKF+0WETTFg29lnQuZ+WvwK7lPQUAKeOpDk4MV9Sjl6Lt0d0xGBKq4O
oGc9yfpzJRR4+p/dmSmdBL8IhnU5T2/eQOo3LlgxZe/HHctQiCdcSLzciHI7epGz
M0XhF3I98InhT3bFS6Jy4ohbhiGsJu6f5J5mOWbKWtCe71bZ9uccu+xgwmvCYz02
NA+KPlyjz6wI319F8pg1aWmpLCd7EhYsBYpJC7rUD9Gyu4Z4K0V2Pc1sTB7PkD9z
rMxcefVoGuqvQI/mvcBKF+AeA8U9/UEnfFLCF+SXsWb5ksg/mxx46GyCoSghN+vG
U9WgUB19D0CzGZunRaffBQhJJgw0d5OvXOeNAxzmME9Zmdh+g4Th7tSPEUNDcw6v
oatqtgdQ2vP3ZhMa6oPOv1BNIVRwbTf2A26+zAQMINU7UjqTfVovWq6fbzEDcTT0
N1gb2HPrxoxVD+Ypu3UEwA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
i7tdJ3fmH0YtDZMUp45ffURTm5LiH6oivEs5ax5EaCe4k6Osazf18NxJ8PkM8ZCg
DxuV7v2ebA1fFM7WTkWZus+XdjtvUtGJJYeW+ux/BCgvxmHvyu8fSW84Gf1PE5g+
RE8EX28dUaxKIDoFbqc6xAKaOUHYK3jlJz8rgmV8UMXAS3KC91I3lPUqC48ehCaC
UNJUau1SOiGfvRnuu2k+0U+eIfAHyFNV9f1Wx6tIOX5Fx9hQpevThkgO/GdGkoaY
MBbpPPk59fQzW75MbtrfcyJuJ87vuHxOkqwcntNX45Luymvq9I/x51dZKYmAo6cw
wJH/1rA/c0LnUoDWBM/kbw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6800 )
`pragma protect data_block
W1tJ+mZPoFTyGasDrC9DKf4mYG7z0TUDPvLruvSMF463pZIoYwRvuSloXrMWwmte
zps5nC7rvLYvAsC/gCfkh910OeLJPR84pUhh9ka3KxxuKtFgCutlAVgyH9xXfwj1
7571GWAr/43XZBiSZWqJHsMKtaCDkg/8L6uGer9RXL0FXyn27H2YLCPM9hvkCkqG
CmlRolG1+pE/CtUyFAziPSCJoudKj0RHlAfBzL6kGUI7VEDzx8xdmdccaSq9pkD2
8UE3mr+PtdoW5BO73mXq3ThLBxBNMg4G4jSVOMob/vPcJJU7CthRbZiQbANXRFJT
ir5JZHfFksmx5mQ7drZEuOkR+M6idf+SpTucx1k+D5fCcwGryvco/gX4ZheokKeZ
O/OA887qKyyzCodygB6DFyfQRqXurWGChH+S5btIwhYyrCWY1AjA12cFjIXqcb5D
fmnMKrj1LEPG0e/t5HEwd8HBB6jdVNl7yyWzLGqKa4jXIdn/9sYuYJ8KSOcvyV/c
Qzwk7BtbOkaDq7yGHM5MRoHI8kYDRgCRSHNMDPNgolrvaKlTweKBAuc6uEKV7zFT
N0QSo6UXrTQqMAufSNy4/P/KmNfqEE32ueLs5WH0KZVaQDbmC4zoCH+kDfF3azCt
E3ZM5rp7t/Hg9ach2lzB5i4W0uY4Tgv/a/CYVd7Tf2lwdy6LEA5jY2HJjjFJRA59
b7mhwSaSqj3943lNdz7A2Q4n9cpAGxG2pFsYrBhxFN9TG4lCx7O+vVL18dBfhBu2
BrUv73JgRQWG547NOjeLu6zE2qh23a32FqmKxu9OdmCRzfJw8MRNQzGPeJtLg1BO
KxWSqOoY6q/4zVQCPExlZVS/DjcTi/O2kkAzSdjDVenmIG0EGzJYaLxAjYC81zoB
a5+QDQdx+TXIOrh0FaANyk4Oy16lDo79OGv3CoFKkN3zKi0OLDepbhhyRaonXzuK
DQrT4+9zAEsFWaHTyMCEOE3/D3OPQcdTBaD1vFjwOlK5FvKwTXAP6Pf1kqCS8wFl
uBFmCJ73Wx4mqk1VyLrAQFQMEWKSIYuzljTnwyAmoEb6tcmgrkX5T9l1Cy/yfCkZ
zWgw3ZtEXQcQ8cq54MtBbO87EAxsbWc06iB8j1mpEMH7GCjFZb9zNoNDBOxQf+o7
H0MDWLLZrSy8J5vV6qnItn19grbwCrs9evLnmCIcWETSPqcUXZrOYDA9E3jVTMbV
7HXp+7lzGdEX2EzJYQtuek8MpmcN5UQBzRXRd/YbDCYaqTGYa67gvurUYY4TeXZB
gScu2AhJlNlQ28TrlUZr78OVuZ1TYrjjJH29Cb8/SwVnbZRSESoKM5cNFwpsWumv
HNG1/IS9m1+AQeZgwmEqfyy7pCugWCIwK9/zzPrvzPf6+M2ofMu4mvYGgOm1B0iG
8bi34lIIIV4hQ0dLEq7MPFYbB3JvnebtMUxmPl2+9uJaWjNir7ReBJPzrTfcefEC
4rr8gQSiJj/eSUwUhg0pMvhLqRgO6kgdq0mYauaiwU+w+j39AHzSliK/9rx9qXcI
0ood/SA/Ltw+MmujsfT674TJnEOryLEHADfI/Zf+hX6SbOraInWwFJ6DmWbgiqWk
+tgtLOWcaDFeU2jqaG1iRGNWlSCwC1pPLgYfAjgCBk91+Hj+YROA7SeCPKubqv5D
xisJzHX3lYHuAUiOV1t0QPlewkS4NrhzOpiIOk2ImhnVMWoMu2/gYLHAbgKZK0AP
xsk1uwrPOg0AyDDBcsFk3oCbESBIQSlLrnvkONA8yO0UsUYaSWe+4ColrOVzSqHH
nXKg1bmF4B7SJXPMT8cwfpffC3ueiAQxKRKBTHJXNvw1zbuFd3LsuRMQnGUhcUau
1xdGleCF4ddoRZEfGczMIZlBJWyhUtvhZMKjunVx7kkxWIzHEQw9xN2sVDvZ2pJ1
ffiF7TGdWi90dvAlytcO9dQL7k/CtNeScSCWNc0wEIw+7q3K3E+ZdC5j6KRO5MCs
thyzb8qDB+EGdoEa9SH1zypN7ZeTkzncVL044GjnTcvvlr30Geh6/uUpml/ueW+z
AYRMoYLqxZug6v2Z75aeTLC7HZ7rbzD3nWa+mpgZ2JwJZWwP5UFujDzhgZaz2vOP
VP1WxsxakAOKjKgysJ4+3RMXKzYPNjy/Qt6pC3GIBC7e7bF6DWwcqKqF9q4Onb5g
C/AII1Wnd7P8m71NHL1ZLV1rdcYKUaWfXW/h08fOIV/nRho02EBlu5ZwafUhoUil
urbGbpT5kBBoQ7gJqCgJ5ltTPmw63GTmVsZLM7tk3Dg82PlOxl2kY+VZVfbQuaGn
j1vPk6E0wHQPl9TeP/RRm2iV+BLdnEbeCxXpU2iJWI62TrATSSm8zzEjhjaJL0n3
vQgkzrqAYL8eIDr0Id3+AOkvxbJkoy4xymubTAV4oPNzIjVJg0Yt3V1PjsmpujFK
qGhMQKR2oTQNNuiwSxoRrrnNqgss6zcHOQn5vDwgkyqR2PD3Ab++b2qsRZW1gVqK
Qot1bkmmhSI+oH7PXko/RtTH+F5MZ0c+41BliYiHnEhCwSJr9A25ylMEL0OWd2Ng
OXBMYWzzYxPrp8Eqkb3CFSYe9OOBt5gjuLiK8Pb/9ctvPnP+74X4WyMe/3qrL2oW
5LTsffvIzyy/Z8HDIPug82BNJUg+4IZ+/qjj2z9NLrj3O1TjBdx6F3Xeb6x0ZFU6
Xb4SJezlQ5UcbY7Epkej1vPV/csIKPXu4xUOjJHYJrLA2BTj1KhFWrXNcaIxzEkj
hLpDuQR3XSViyuDmnuO1/bFsMfFwXnDJ8gP0jxr2MhiB4GHsAVcAgmI5E2635z5T
mxAkyp6ZyV8ws1CVV5cSV7rM7LpqCtUk6IRuG8B01BFVZ98sJv8zczKivIJbpb34
c3EzRoGiASuzhiwUjj9/W1sNcKZeSHzo7iKDWsB+JS4h/TlTCWhmK139rFIadmDo
5FKRIcvcad96SoxLOeEzvdscB+fLUU6MAAfr9hWFLrE2vM1RSnFOBIAjf7N34KnA
5Cq6ZN2SSPCGNP1mfIhAWPX+0otLVc8GTvEUF9pfG/wIGcb3TAhdjLaP6a7g1KPs
EeA57tAQPJ3ZW6pFEDTmezL4z5VXC+WDxMrElESehKE4A2gJaw+1GRN504P37aja
iP56s9yBh2PRZE50GTmrQkNr30DVq9PuxRc7Ozf76B26MBpZHvrx5yeMz7rwN2bw
lwgr42es+AdAcfdiUFDuJ+uwHXgC69cLu0iNJFpqBzpR01Uj1lnUpv3iNsbmyZ1K
5suvcBiHsQTs/32lqjlcTMPf9KvYOskSirkdAaRc02+XztHb2lWNlKGq+4EyeviD
467gWN8qv+fG4ljpCUjY392iKkGkuf5/ABfVQo3DAvbYMQUkfwIPUMWpnn0XU+tx
orM447ASPR1Pvo0JRyIgHVtp5j/miI4mMh65u15ygIXe32lLqXjtD3gME7ov12QH
0wE51IaZnERxypUnNY979jI6Io1EnR+UUqStiR+Qq74NFqzNw0eH6OXdnizJ94bV
i85vLSA/a6PAERLEl2l3I7pHo+Y4XXnKAiraAevI8ADapsM5tVT5syJkeda6sqJC
vhg19xF+jYlQleUEuy4ipW4dAz+GBOc/LfEhHmknzOaUKbrZhBTf5lMFs6f/rOhi
6NuxrT8fZHkrTIOmaGlwyBt3wUtuX1BWUjn2P7m1jwiCmxJUTizbKP7h+Sr2Q3t7
tyzsTSjtnYeGb9T3f1BOhnT30ds71A+C2YM7fl1ACB1tC+rMAtNeukNlMefcvqeY
Y7lcerx5Hdl/1THiiixPpVH6RcDZRPkcLKgRa6kLhX29H64SsRawI+/Mbzq13VtL
F9loTrvWgF2XvuKkV/4ssHuFYyJGqzUtE4+jRyW0Hmiz3qmfuWpIJ5k6/2gDhQwg
j5bdlQHy9XDtyEebWKfDkK7AdP1d2b05r6zcpotcNiEnhy7zwnnpy/SYlkOR/N+d
3coJL6KYSMjg/gmS2IxZ0TrKGE/lIqr0m1mf0avzL3nwleHChu+OdeSGKV5AwNVS
XCq6xnR2wzn0fPZFLxwxIuu52Evm3MGjoTvB80UxE6MSwwxorOO7CuTpRUipQJ5I
f2zrQRLLzZXhheSLAolew6+4/6Wo+Lw7cIKu3S54gs4UGkyZI/HLNDOuI4LiJfBy
CUr661qaMZxW4ebPJlfuFGTseBTxy0JoQqrlb8ozysKkZ8unpo+sJjDlVrWK6z7X
fQ8oHA8qECX1Rensvs/Y4FsQzW/vbmCsvkDQJPAlOOUcP+vk7nP7mrwBRHjNXqxk
j1/iZhagYMx7GtjqCdQofokcFEslb4vv2fcxpaSd5kv7pJDiHtGgO96+eUJAbCV1
guCdKIRaGxu0A/lLZ2V76v9Co7/c3qOcFVgGuPWhp4UbdNsaTgw60sAo0wGhWzPm
I/fHixiNsglcAmOWNxiVTSzji8GuuDZbkGQ1bTyO4JX6ZTjR4GQBPUw6OynqL2mX
3BvPXKk9wi/r2FmFEAzn+9vYlj+2fAm/0DfJd3T6p0SUo9aniQVIG6al3w06zYBT
E0ksJEi1zjxSUncjVZlwVWoPUdAMVdsuVoP1vWRR+HTI3hFiGqu/5+R0yIVE5Cig
rv2dDIaEGc/XqTGE8iFkS7e+M0ekGPqc8qb7S2FnUqpWz7Kto0r7sMHTDKHEXFzU
twTsUiHOR/kdMo2OKxqydTj8C25EdGbDVUtgzjst5A/pFuqFO0f4Az3d4pTZRjW8
wCgHZ/G7pSv1HPnrbo7iD6m0l/AvvXWR6Ifg8k160zlDGY+VHlsTmGoAU2n9HDAs
mu2cuonGq9G4AedYMPY08/uHxxr85K0+hB9JQRxjFBclCkRoIbKOvB6IA+YJ2qN+
ocv1du3mZWI0G1iJr4jY6tSpRUyS13v7Xz57+SExGiK2GYsS8GzmGMuDzi6RueG9
Y1xz1xZ9oHlRw//4GIiQ3+ZOOWfK20KH1zeFWNg8HCtGjV+VQrH+058hiZEPQ/i+
zwkpZJOn92ma/70RihUGSEUJHyq/UON/mH6TBwSQvzNK0Q2uDWZSsE+YCPONQnji
sbVo0zQ5u2nEHHi5X0czLgkZx/bd9EYn2tyfSMBQj85TD5JiLP6/FtqtxzLnDFtO
dqhiQ+DHEGly7DWnkRzMgk54ESQ2B0XYmvgJ5Ze447UJ7nxY/zrQtXC+go7WCkSY
c0rhHXS349WMJ/ZC7AmlQ/V4Hg34g3XbIJughb51ms1fBjUfl7gJy20eLZpdYQKk
0kvJ0J0iRnIhGLef4CxWIOWnEzUZx+Wc5It9N/54eFten8idCOknUQuTmBd9NPGK
B2vFMLBb4hhuMfOnij8mx7Zigfv/xc+kv7X3SZbUYjvb+FwGqErAkwUcFfB+RwYP
fapGecfpTb+8uKTUS7XRAsb/J/pbpiP1s8xvAJW4dE3xh2P73GUtf9nL37K/pX/k
kqG74auPpA0jfmg3szL4KglIEW7IHBij/lgGle+UB3J3VEz72P2WT49/XVGFyS5D
+cFW8Jfk741h6wAw2UySBCxXjJ50bYIoDE4w0D1+KqZAoHUn8WS9Sc2p+naZubhe
7aYrmT6A3vBzATc5Y14vwbQGKcGuZNnKBRItM1Nhd7iYDTelGf/97Csjy1Ex9jVN
R5ie3wWZyw8TuVKghYwq3zZ/vtvemRLNzYg34u0+t6AzV30N9N5jG3FWrdPZM4aL
k5CIbVETMbhQRpPa+FiHG0CrMsr6L296E0DSP3CzbpaINLgsk1TAVuowls/ANFf6
12B1ocUnYZgiLMiOgc1iiBe6ttqWU0gCmBcaQPOI+k6VgWDhzb0HXFyPJ2xio8U8
zti/f1AkUCyUA87giafAAFKwrnd5p5ARq74JCuKNdvjMPMs6sDj20c4uiD1fkceh
GsZTOMk+dkmbRRYPAp/q2fpnXI1SYI7aCRdrkUNFvpXEY2QOuzsi1zN+qVMutXbX
YCm6GQgTYZ9y5tMdJbxkKi6OVhswmokkKE+SkNRHoQxGetJ/czf/oLFN5Kxl3AtP
o10XT8isdkbvp9DGMycDIM8R2qcV1NB6YF3oehHfvATuHl2t1q7lZUdlTD837Chs
uWGPjT347BC4rAomghLgJ1QWxQYph7dYJtkPayU/Xmanv0FCIR+IR+zSE6GkNkpO
pjYs+ZnIUkVwkPk+hSqH4n4z3XCdh7LfDjQhEhD9OJZSX+o5kpdz+AnSm4AqXRF3
tnKebtECv1MlWYwhF4zzfIRNivEA7CO9kkydVc2Q/3d8Jp4wTSV+85OgGcUapL7s
jDTViJpe/XiRf7mtVXquYKMGJar2Q3BoaCKGAbG5W9HvqJZ1OK1yE36CTrbEswlr
CopJApV0fjT/Ts/o8xmSLFZaCLU0Tc1C7LAjB+t/RBQIT7ZYZZnPu6HK4h1B7elz
h0gut2BdCXEeg8nKy5x5EbE8wq53yslFuiyuxjvAeqmW14Rz9z6Kc4dNrKpnprok
U9puCw9WG5NeEPLodvHRp4ZRgLSpSTSzaSUIGNDUjPF8f5we853/A+wZgRaPTBYe
HK56i6i1n180RxG0wvV7nKKvXQQcp8FQEOI5YZFvGGmc5SjcTP/atyuVu9uuffrC
ygvGZj29Yd/btfYVNSKB2FXShqQDoDB+oFhfWnobGVcJzYg+gu3YGL7CFRwCUj3m
meh9CMIJADqq/gvpoc9rUeypMtHpocpbOdhiObpolW3V3RXj+44YroBMpD047yGS
4pH5IfP8R8YvpR2otpirAVVHzFLCDYprtlIfhU4Y0odixIGhAWu3zDzgQtm3C7Xp
fbTsx7N68qtE1rrMmwiBHqPBWSJ3ZtecjMbDavp//MkPqgRgBVo6O5tEHIL7i5Wa
IdcILcrtxU+dd+4j4FSQabOrs9tXZYoUQRCatbujo5/pfVzAgMp92wYomnZnnYf0
y/33rTIZKMA1KvxLXxqpNUZ3AbEymzIZ2z3iaZHBtLBQQGNa3YWulaTF9uy0yXby
ktEx+2S40L8LC/WOGBr5WdH/QjDa0zoI3FdfWTkUv8HpUIKOo6nG8uL7bymjBN1Y
qNAJgs60SF63gtBUgIn8ccU3kqUxkm4BJ//DqkG62ZqnUlqcJd4VfJZZV0y7itza
kkx3RIdnu/AKaT3+1D61RTkSp47XGKZNoX9nPsOtpvWgJ7C4FRPD67SjTIbUagTh
6n8KL7uDNVPAVanS/3FodQbtRAn6/XwqH4ZQKO4sbQzQD3Ux2fk9fS1CfRcLstZn
ea8R7J9WgThhZPCjBZj7sJ20iee1w+A0K+R7sxaO0PKCO2oTdZbnE8NTYoPlLVsP
5FiDtLmQuMsHwGEVMoIAV/fpHJr3/qEu49u73+hYb5Fr7vEh5ns3ivzHx3/sMNls
mUmiqV4H3dW2Vb0PCGN1xcqKBity5dafERZMM79Ge2HBXbR2Ug1VvuTM5A+EGnAL
cJZQ3OCeX2tsjIFSsPI1S5X+Q7El77Gp7ievexg2Wy6A9gyiCGalpy8kGbzZ5FAu
ABPejHC2w6MtkA/jgyV4aPeI3vGscC6MWGq6bBgN56augjC+XVkrQ+m/zsqtDJnA
LL/nw0SrCHV1M68/yJRi/uy1SDjM2PNkUlhu0gEYBESMYgkivyvXZx5B/bth5jHn
sHww4xaUWAppqTJnYREYShMrihIgc+Bm4NkgN20i2Fput5wrRE+J3o03o1V02DFQ
ZTPuLmYHNgC/IxMqk1r+lI15bYKrx1LBRjgd4mKoDr+FUBd3O/jgZlHsS8RQyMMc
F+NO/bfWOzM4DdabDuij7iEnZX2qdlYGGxmYVvMxEM6O1YK3NNwZB+OBpJZgL8D1
sXOXV07rwZlQyCWoJaIZ/QJuSY9+KkLtGrjB9wi529FcIZMRhaP79COdAx6D9q26
mHSdBnFiJhEjt2+izOLyvnQS1x8G3b1goh42VC/CZ7zm72HGr6jHTFYnDZ6dWRv/
0o9SRdWtfu8NtQSXjQ00W4tnJWZBv4yJ9B55p7vuais12L7xZVtf9JEwO8tUOXt9
64Om3PIo/Ol/WxFMJ3hsFUT1ri9kBybfWdYab/VOS/XhXvDoDd/n6YbljxjDlE10
8UE/SxG4cLYSxqKJD+vXUpA2QbDw+dac9DgdbMY06ERO0ZXGEmU1yNmggPe37Gjb
MCN/ElmN/eI7f+3XlJfT6C2XxUWmRPFswJxZc16hKrZPxrtMbzttbEoSQQEpnAhh
0XwYZ351ikdTud2WahxOy+899KJ9P2gScBGLyJ38r84dMeE3hQKDdaJxv1sf5zTu
WbiXZhHPtW/pkL9Cchk88ocJhCJa+zCGDMQYF3wokC7i2UKKwlViK+bD3WLFaEZg
ZOBTRh+Q/LasTrXaHUxtmF9oJRRnHEESd4B+Ds9AwrKVVvgHcgA6KzS4YDWacVjR
KR8xe5WXtf7w3V1HPVhStkX4TLJd+OX7872DMdk0WgjipSLSlbaa2/bT65veGaRG
dMMcAkKwERt/m9SxDMMOXgdlyZCiFAXreh05Xfb5+Ho0YBUK3gincF3QX3siiXum
TgJ3q9AUfvXk+o24T5v8huajb/EJU+OVurWx/7rMdt8xcdECFaSmF9xfmTsJDxnd
BoUp/ou/1d3EG2p89KELX2kx/vLurETNYwW8bJYfV5tOln4tHfO2LfHNZloQU4O1
/TQK2jtxKQ50Tw5XKU98ZHyMmVkJOsXTA2eQ95R4Mf8rOSIfo8Sa12ywRoJ/V8IA
68/lHdURZ9X0Ih4LfhAZH3l0/K2qRsZfMCjkgLk54Vx9/fnL0g7jEZLeRAA9Btnt
jO5lRRF0ILAsESlHVXTG0l37gGa+MTLyjQd9wwLEVpcfuS56pz19LPvf5abE7kj4
IKnryXv7oRTVLt38O6SgSxH9DZ8jbqb7mXgGa8FpOLyF7YAnFCRXiqjaOlG6tbB1
sg6VjpiFYCTCTxVtr+PjcQXCTBGP9eOvwb0tnYjokJ/3reQ1Od4I8nvPRmnlqNlp
kFp2hAVSMXAyxrxentfQjcQmla+//gHSu5zqEyLUD43d60P/CJ9Ci9n2oMqpxLof
y21xRjm5X0SsMMqem3J45a/5ziiWx8h54A+UE3FUm4g=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
fQDwf1SLDql+Vi4k/VGTlCir9H191pg9MCar5w6yEXs6iEP7pfLSaMgv2BpmUelQ
3nVLFVP3R8Vd1HA6AnszK7VnRd4ngAne3RsgZrQKi2X2vQUqPoRqQQ8eAOpGw0pv
2QYYw04A+k/Hq2pRtoSbxP8lX1267pyu7QTFfq8sLOv7AltjP+rM2/CLb0VU++Pt
SaYaW4inGoS6gkO0FaaxMNNT3+tPw9jxUx0c5e/R4nuO02srhBo/W6tMis/35q7I
xVCK7z1A10qeWGiYhLNhDYVM6nM5ymvOuCMlbwUsSoUgzLrJmVXBe3KO7hZRbpQ8
16FGN4hahI3e3YJL3pyhjw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15408 )
`pragma protect data_block
8QKp8qCk34Mfn0eFRYRW6WgvnyqGS3PyCLhxAkvIg88Lv/i8b9Hl+rH7tvnVMqb5
XoPgwCkBoSzuTz1oyqwLYzAGCHZjeDlYBylnlY3MO3OYdt9MXzE7hJbRs2lTFE07
u0giQ8tXX+Jgl/JytTA08pjrUuI7sruX8g5rP4waUM1VwF0pb49qav3M75z/KFSG
Aofj58UXYgaZWpkFQOKFwFThDrZx0psKh+2j0qzdHk8JEbILbBJ4fQuazirA0RaG
y9VNBQqGU62i5JNl2JzO5hOYA+G4HR2/pp/mN5TRWmA8K0r++SynliTyNDhPYLLi
xz/D3Bgu8Yu9c6vrGzgC/42+dKmQIq5BE+WHHL5RJDKcAtxtCrZhg7/AozClAzCV
3KMAvbKTCDJNYFO8itT/IPZUSuaxXIUeSD2CsSJWJxrDm0YyhNZlo6rqmhBO+c9j
y4bZx+8qqSRIKvTPfEVEXcK++O635KlLD077G1fjNiBqh3KRwuksbRvYqyAfVR3t
2MlUK2qEI8y3IlAroT6cEmMLropwG30GSi2UKSwxe4a3PDxnu+pLcmfMwx+NBdOG
rTk2JaZwr/+V0cxDSdZ8V4lGISnItzDANAxKuuWdOK8mdIWSpSKxt8y765XDp8B/
OTHO714zLG6FpVn2vbneElrnaV2khdRiKwP8K6kYZxIs1At1QDEFcq7qpDiRkrms
iHB24GMPBfRmpBJfk/rUzflayGNBe9bi6lEaJgvWcOfaoKtlCJUUx9t+OiRkysw3
j8hfJQVmM1L5m6dREfDoe9LnNmdq2TLxcQBHNgLgEkxbuzub4k9NOJJyld1eQ+Ki
Tfb3yv1hFVQITQ9ljmu6eL2yHY+W0eb60gKxKTJDgiP8Fvyi0nadvnbiHU6jOrFs
l5LLB60rConBai1JMH9bPSffvvJjFeGFMnIJBCz2L+DPIPDwKSmifAFgwyrpI8Ct
8TuFk2NZOVUxPA0ZrSKcbjpqfAkJHHaBWy31cgW1BjE/yYNIgMZkZ+2c88cfY4WK
zRls3ZqYs3qkzoAAGRmxIITmDxfT9lxc9rrd/QdRhFfH+V8zH2NEM9c02o1coNlX
e9+c2kilOzCFl6vb6k/jDbk9vFF73EZv9O5WMDEQNZCy1OWhauMcT0pTrJjooULA
jbMnxyBHgxpau0aKz0KuEuhWvsuOIdOsPYgZC7p1umMLjR26AFGXEogXfBegHhgk
IVt/kCpEnusHrVIUTE+GUb9qnHNEogZ9T6ct5jJ79BnhrEhgkoYuAUFYcHo2Yv6c
tkNlhQqwWma7Q1YpHnYC5tdzjDZYp0bQ8D9dZ+L0JIIqShBnTumYxsUNGsiYZsKt
rN6okO4bjkaCDVGuZ/+9a1vj/UjOu+ZXczEe4Zewbz24KlBQJBaodBdUP6EcaJcH
rfM2hXAKXNh2NbcL7SGzVlBZoUAiKvg4p+tR6dlzG5XVgFqtaLegS2ZyiBUTD/QM
zSkLgu+Be1SNrM0fhWgAuVLuy5tPeVzYyvcJgmTtdIFAN18PWFjp9GnOyQ3faIsV
5uAdyB4S/tjxlUBMlm3IPWgCXTyfnRpEajPeUfQSsmfKsNaznq+YKNi/E1xiBye3
LSuIHD9WXhgUwXvVsFkOlKX5hdCiOWx6SmFmiLCXkYl/IKGEVVnKzSqTYfAaheQW
rIQUximmBotMCdW4dm9XJu5BNhMg7VQUn8UR6vtit6WlYX4RER2Z+3UAEF0Lgy/T
rkZgw1t7H75laMIGP7J9ffGqZSCPEJJHBKB+6mP6Uygg2h90KVKh0UqnK0YKHQov
ZYSpwmk5T/UlCd9S/yybbyciedIQ34yPLXmmfyFcqzHg2bd1Yd+WfyScvalYheWZ
FDswgrE/tpUVhj0FBMBuvWeUmwZGElagJZg6Wk3VvlnxGhrg6104Nchz2ZzpVLvH
KpfX6+R/9JnST1HYQqwxJ3KWiBMR4VhszqhYwa6q8HToKezAJDokDV2lTMme6Nqn
2CPq6/1DnsQ+SRi3QpNd4N+oBPB78uFsPGPSCrnYM22ec2J457694CdcUU3AVn2A
P6bxcRC2TdNNQGIeps0I62oaRs/ZcTWAJIQd4pwX0ufzNhmGqT0Ks/MCrqdhUiLc
DGdnIoFA56Oh2+iwSCUqvI5ODpDV1KXVIvr90+loLQYgLTrTmnBZKKI2GTxslzNC
JVvGLO8Z4wfirsZGO2je6Vk1A0pdi+uVlRrtnhqsUO4NGHvSuI14lURtAy0VOMqC
9eX9pM9YhANA9BOfvxn3kaUnx9ZkfZ8IY6yy73Dc9Ojgc1fdm0vFETE2nJtnth5i
+z5v7VHYTLmXqWSeEl8QCkzlLaLFa3TKDjZtmSNQaaQL+DbU+etc4OvGBH0HSQjp
5u+XncBvwQKsP2X/6gEZ81eKpgSWbt1Hrf0nx20Zt0UoDhzolTDB63yKLjWShyDD
1fvoQtT9RncqBADQgQNuzSzvF73roqh5ERNNEh1++qsQ3MrgOFmgiT0HC7XdXQiJ
1HyrWRHgzozpM3Ths0Vr3DAtbN+Vnv1UixM5gehFYY3Bm6eCOHdowrAsFU+rN1cs
lCpL38yEvnACEYhhwNtjepAG4VR/C4gWqKv2x7/XjqHyXV+4w+KQWNDKdsiaakqr
gbGTieNKkCc/EEHmP9bvmsCVLLvjMqSWP6MdzgId1V63s4Tkd4buze7eRWICmTzx
vYydVGlji1fd8Gw3S1VZU6lUzBJIpxaUwETQRbjX88jJ8JEKBWmgAFiywA3IAtx7
wu+JR9LHiTV9E0ZZjN9OuR7nVtsxe44Ho8J52MvsyN0oMxBaqfYmM8N/XfbtcTHh
FbvJW5txYlM5RnVNU8fZJVCBhrLO6p2W053XIQ5AtnL5alxpEeigoPeoloud2wzE
sNOZyAdRcyjZ9tx53HEkkelfSZO1VM4m7UYKDf6p642iyAHp+8KZxDlXClIi5qrZ
6xk5TnU65mAnjdHOD+PyIWZf9yszkw1QaXVKmru/TomkX9RUDABDWQy/+CrgQqAA
yq2Jh3Iy2Ci7GXGPxU/q7LP6Ex16ZBh9jHvNOqAAWRNcCU2cRAWpndV0v+cV7XZT
Jc7L1TvzI9xtgcPxCgoiaSeVSDjl3RtXJNEzG0FrbHsxP9xJw+R1fimQh/U+MUwt
kXzjNWbKs+X/3nGme7ZaDBHACGLn+pq8CCTKZqUaQreesLwCay7U9kulwixaGZrs
s50fEpd8seSUaK9mX1Me0jkrgCsBT8QU06zumBqp6gXUbmF/s3TKCElr3bGvqQg9
By30iVwOYF7EwP7k/uau3ym9lD6NaG0OSB+tmEzmNq2gfKQbAsUsBdum40d5NFI3
Vb1Fvxg7tj3LPanHCEbr3ZrR/LctzlQ1+AuAx+3duY4o2HNnDP3RjzWXJvG/xfII
JOCLA5tTtLce14i8h3xv164+vlZRtwjBBct3GRAHIXnwo5RpPWQXH84n6fciMife
jTe2+4wHRl2UtAUPNardET2Z1jkHHuw4WT64m6PMFJB8P+dlpqs4RPF3ckMw/QUY
lsq0rUjn8lbhTHf3DIcgFzt8rEcsPYCIiy7LFiQq3uNgA99lH4oJyVGHFF/T1vc9
+1oWAxrvcC4ki7GBl1X7Ozepbs5h6wd+I4qc+pH3viSndbH6jsyzYVjf9LUGtJIt
1Y46JizEACog/62ndX7aZPrnAGUlakfwXFTiOw47SijadrbSfJ9ZBx4iRtrZsRZG
no8CY1IHF1Rw0P9qYoJR08ecj4zEo+9MSshPFZvmH0vKxDCoRRKZRotiRcXYWc9B
75IWnwrQUMKPYr6abAnHST014MIjoHH/hQqJStu5Gvzxin5nAZsY6KjpHfk6DGtT
UPKpc9KMDDMYe8shf4wREUyAwgHCa4Y1LaXBlRQrozTk/LJsij0eqTkPSIrU9gOL
E9P6BHjjjl02eVmiVsB15DcNMi/57S8BCkMrpT3+Hjndi5q+T9T7VDyg+fDW7G6e
No+6n9gNxG/VjJ5+R2/QD7eY+SQEsSzHuUgzk27UjJts1e5VRTz0PB/bwa2Yy5Xq
OsO0vbw7AQl/JFS1eHVtdXerRG0D3zdh1OEo32gVfGkE9l1edgekLSdTnsHRBF5F
FJc7bUvhNl2R113gvPoXjhDLsnY8zvO1Ael98ktTgekuyRBo4eym0H0r64yOZddB
kc/vqvxewg+E7/VH1qIxd+jKs1lvjAJcP8NDJK+0K4pFEOtGEYYQehJsaU3sLQJq
9096WXXc9NIUAybutm0hOoYjPzt0FeCTEgz6X8MowMz6UVhtpKo+MuS3+ybfMdWI
OHMEU6U8EH94C8jOnL08Df9oy08mAweaDfPqg8pvDv/whiClU+uKxwG7Oy4SzJ4U
iC+0lmlw0sIcWWvsI8g8NYgbfDIptqAVOEK28GVbyvTXR7KmiezbXMgkKaz9R9SH
PuRg+LUFI0BCDlLYTWDuwq86MVRu+BpgTOuazc6mJ3cczpDIbVoadVQTpB5kDk9i
+P3D+pyYD0dxDI3XKTd2LNpfjNecyjUtyEAt6yiYtt0IKnXR6HjA0lQzAQhdvJgO
ZJfhoYVV53WHxuB5o0rawRXKsBhsV7NaPx6gplaHgECkXSM/NViHuN0jZxsoA8RR
I37sZEN7okT3jAd3iBRxl1YZAT8Y0j+yT3OaZ/R0Cidt6kEbwEtK//Q5iF2rQatZ
JnnnsIhFmpYaR+EgV8MV6pb7WCe7YnItZypM9KEDVK+sAUdi2LCsaDSVEo+PFH0y
+gVXkD4uYApBw1+s846xOjYLsZBQHULY9641cAAOrRvi3PewvA0C9DiO1J5Esbic
mBlzbZo/tSEQerJkVpV6BOev8GCw/jCkVTGHs+H4YZ0E3FcnPmSFM4qAVrQS/bdY
RyW5gSQiNA06FWBtAD55dXPpxy7iwthxD9PZZDWot+5o8Pmdh4p3JtYtQq6K5p8J
QE1CC7Z98tGrtMHYFHs4moS2jHi/E1aML7Tz30Dv2+NAEGS3cZSU6WZZM5RRUkqq
viOCc3fYnSKQtMAm7yUhvpeCaTtDcAHgZv0s0Sw6btnNGkhuuT6ib6qC74XL5hCE
y+5Lyw7NxAfJcpMZjDVWOUqLczF+0qGIu715X9OrW7bhr6CJglNn9qNs0HGIl5qD
5WJD2pfOWpco7AHWmGBmOxPLDVD2EpMfCmI2ReAxj0nme/Y7nrU1kx9gdpWCkxHY
lgGLIpjyvzHZyaTAvrc/uH6SYWppcdatJkUYzaNAX0pHTLDp1jLBqeC0nQhwzCWZ
mPK3uUzq9UVkG9n0EfJVkLBN5wP0EmHNgDU+jiA1DOJOzBiRbvfuoC8K5ZhqUyvW
wSo+N3wjlfETx4yQKqxK+hLw/LFPdpoNtDRFCvH79jOZfy79MdbrPA6p4zYouvw4
qvbJ8fpTqvi8Sbs6XHc7S0P2L5/5oVWt1IjUtrj6/mDtLheU+GAQkQGjXaoelZOm
FJVQbRTBTPj1ruRdp93oJMyb5/5Uqch5OPRFGBd6cCksvFfzmNdTItboo7GCyltZ
qqNUQnlaCWd9baBwYrNyVUBe4HMAH5dGCJeyYGswU7ekqvl+4tRWLuiR1kyHn9oM
xQ8nmQJKM5iNkcKsw4CLjz6inYsbYY0JE5a/3TtFlr7m4HqKM675Aqyxwrc8bKr+
M1KBODsLGi3xZWexH7H4MbGiRx9yr15H1lIkkB+BsBxBRtrDrwTNu9cr9uF6Elg0
5HHSsR3p+V3zKxYNyiWxegOLwvqhW8qAlO6Qjn7OOC8cnKrYLOa0T2q18eZ7pPq4
9TC70di/FM6Girk7AKbck5trcRcZtI47L/ZoYlPbP/6W+LBVLIWFXvyy3AY3qkgs
rm+OLtzetiL5I3U0FeUCnMlYEDzanyRgyPWxYumjJY5zuq74jAoAWvhHtHK7eYrn
VdZtWx9lupW9QHitf3QhVCXpXibiOh5ogqgzx8ZqELoF6xEQaCXTuGjiCGZrwKW3
uQXQhDliAov74IdprO7Z9gwKS117KNUVMv0advNgEwjgBKO2aFqeD0G2sS+gDag1
Hwt2uPpwSEEwnTMKTxSfVEszKbQVsrJf3UKJBhg7qwGj6nnRTBj7wHBbPA1F568I
JzzCqH3+5NNsH1VSGCIG1lvDfzalLkQYyrHf/EJ/+1dgqJzik541nrJHr9HqEOr/
IoD+fntLLgpin4WToOtId24T6jRwYe4weulOElFcL62VewitIOYEav1EYthnJvw0
x1v8qSfuA45OKWcNlP+vG9Ap5HTV/6TA5oaBmLqBR6hW3elBCmpe3RQKfsVg2Ndg
42d7+wSSI7PA5GqOOrZsj+8T+V8tODwKwsAJxe6qT8GieD1vx78OsyTJn07Y6bbH
AekI7hyRXIjr617BMir2l1i8QVOJS5YJBBXHhU7jKzItBuuvq1ruJ/eNd6H/pysY
zsDLYLKLA0LgiGwMMSCp0l7i+VFvkbQtM6dNAJsZK33JTnxWtoZx9d7DkT2E586T
AAH+eASjBu0vdCSvAvcdb0j0/1GU/hsc9y8L2MUOtqgK48dHwg5peKODLDXDR8Wx
7piAh+rW+mdDIZTHbkOTKy5zdowHb65B9Dy9P2XHeYSjs5rlCBPh4aDUIukaHgHR
Zy1x0PUet092kIIYF/RIYAjF3ScaPLhMx6ANDneBqES6hiGg94LKwvQMxS2rdGSC
qBvcVCKrcKRYrzrje2VOKiENDXynJAWKeRvwBHIVneTTJLug17R417lLESv45Gmn
EVl4H1J7kM4DkZwPrMu9GYF1IgQA48SJtefrRANaP7AB4ClvsVgvf0tuDhNik/Hf
ciXv43PRSVaRwx8/3uyX70mVVCD/AVjpTb0eXmsf032vQ8s8pqct62uvvsfe6LOG
V8GFRsD6XobCpT1jXvzSxQkq5I+SUPnxXCZX/WcLiijcRYa0fLtQvlmF3fQmPaSW
4RWaXa/E+W12KmDpOgQvmZUWIXZ37xn/OJoBZzPHaLmlCPmPO8twsoHNgt6vNDvU
v6gWGyIf9bsIMpP/6DE1p0voMa0HdJRGiQr4iJpgbrmTEKhHswPKg2Q3MlvGgWQB
hyStL3wio81Xs2oIZCXDXFFevmKHc3pMUMnGaOq4JIz0CVcLWVaysfHBEoeoSYM6
ToZKX9C4TBGwBatreSXSmuhL0R7uctdKj9woj/I59YNgRoX09QZ5Q5HUYtzIgp42
Ku3oYhBhZCL3ajT2ZhDaJBCrQVtSbOBLO4Xef8fsL0vLPtzmCPsk/SLI0Ndhua3e
Zgj6Rrr/4bSdyBT6TNpTyn7A8Zmz1SedbWqXxBFnubDQTS3D0qKR9HzaMxsSB7g3
jnob8mklWyhYgYL718HXH8aqZaig6P16iXr6HURAVAlaGS1qRrVm44+6mIJoqffC
l2UC4kGB978FjmO7nQaykLeqbtY6jAz0WrnNeLdDR1vmEOQZTlKEfuRbSN0jKPh6
iJfhHHeALYBrCa9s6l9K4itFgnXxh3pVdHstMaxuPqAmIZYGw3PJPWADE9BzLg8t
sAb5mfmXvA3jz7hxw3kylqNsPqOITWtH7nVV2qt442rGAPtFt0uX/fhFC0Ua3MFI
kL6dPYEiLZuc2pSS0Wu1Ha0GX9E6a/rgmqu4PBZPDbB4RU0KdKGh/8hTQ5NJnxaY
cIsDYfDczIL8J1Jek38vL6S/br092VWU3AXvGZVSJ0Z3kmEGFnWMviT1owNTmthA
ODwlGsmSw80KPckBRwDki2Wexp5lX8XjXuS/ResgOaE85IeWLW2Dzyb8SZVFHoyI
BnnAeMiDCOyZPx2IoSAFMB1vKEyu7vBvPJabVcJjewC8tSSwpsMx/o/GaTmA36eb
oF3wKq7530PR6vHE48XWpuXX7jUbHS/brWQn1h29O+AW8cbYF9OQOlKgOncov1nI
U00Aw8zSAzrzS+UhqwMeWkg/ipo/ZpgqEznHfbO15SpLp6pSZFzIoE4coxyivco8
vUEiKfd7NyHLQmq2IzFiYNVx58DMJfYSyOhWM1N6vdhga91VkUqTYFxh84kSTNeN
I/MM+9GXn0RwT4+Qmre5c16SsArWLfrB2LRDbt8T3Z9Z/et63OPJihC+UV/D8T8C
QCNnjDIS3hiDw8c/dKwreNtgjHJYd1yDrAMZRjvQOmZArof+Va2Gcj+BooOQhWnT
kiVjbCKNG4bG3pfvjgE4d6g4+21JJENHfOBXUfnypHhZ63mRe8JA+G8erbWPeoLR
xuQ68Y5CEflmkbOIcW850kkHRHKoToqLNPQxSW5K2na2IoSTZM/bYYZgdFKCVoCU
y7+oWhQUxzTQnLbp2VXJEuEZew+wzl321QJ6SXXJYGU77ld9UXNPG5VcIPyV0gWJ
ITpZ3Ub38XlHvj6DM8dMFp249bItd220/SQlZsXrELwxFQgR8VQDJ+IIedOo2KiQ
zKfa7K69wuCwsU/LiXRQihy8X8T/BYWY+LnNqCcQa1Ws8me7gRh++CPdmN0m1Z8s
+wf0o9YhI4AHTCJU1UYy+aZ3YY6zSGr7H08j3DZycmetvDmXuhntbNphzQh0hFUa
oKLaAs6EuRQHdTrW2tWaXPjW5oIh/BwGdd5Wh5tTgNmLIeR3Pw0cb/+/Fa/pxRah
PyoBPVQgsBOaWHeu8G3JCtgfu937VQVAUBX2KkOLAn53SUq42WmdQyEWZLOVWGvD
mLyWTpiyEXkclp3FuXhr8QTcxe5HuDa8ENVIzjEDCBIlRJniS6WbGytz2iO4gx/j
hfgxcqB/BZ3YIAkOjN77Fgr0s/z2nDCPPB9BW7x7iQRNP5o9LcO7oQihINE7JDaM
r+sUFdE6XSWnPvw1NiKtbbEIQS9Ft/amZt2QquVcesnoThcEx2aNak60pBJt1eqI
ZaKdqXLn6H55D4+pYQM3ohhxO4zUSGGLQMcnULZJABCKjqYp58EVSatKxsffDApx
u2+V+nyEhiIur9hdPDV1syrcd6EHkVBsp2LqIywrjiFAOEZMUCqur4eCkxZNxWls
qjg3r4QW4dIWonrn3WOmfuT+jQiJTQC/t1e5cqzXWBJUbMEXBdnX2AfsSgH0MISQ
PAZgX98V/kYjbV08vtd/o/0IRUJFpaXIyKvPXyMD0BvpkSuX2LnXgopQH568ilWc
DMKMuITcYeKP0VGQc4rUrNI4yswqFKhqPwZzcOi3epJv5JCYchWiNEaXvmVx2D8l
RnrWdWYRFrpdzfteIkUoUHd1NQR0aq6/SiBAwDrs5rsT+uvw6h4veRrwnU1jVzG3
bW85wuk4PBcfAdOn7LjzfNBusHVqMWtgNzjOOuh4cnQBz5USVYQikOSQDEB6VWne
NBCjMCmIuGDzeDUmylwpUQPsmaA/jh8sa2SUbp56fMG0zKKwTKxviQhCbITk1fGw
rEqWxAjFogmw/Z1qRXVEU/ygBAUvjrK4Jwtycsknyy32y1DQ6cmFAS+onaP37+pu
AKxrOYpiSx6k40hBarjWEl5jAjhXvNudjyovediv3M42eox5RvZ+gcFDY4/AWl4C
di/eLdr0u8My40kX6NnVWu0Ws+FXd8NFnp3WfDXHiOaAxuN4lvgvcUTxSBCaMd0K
J+j+t7ocvAWUpyCcRyFW/YeTlY8HzUZVRUe2i8ILinWsNV9INvHzrJokwz1Tw1zB
nAowXLiXxVQdgRIR3RLhOxML7odyBvV+xU8KfCNp7Wv/VyvJEukKSjiUetTeEt4+
tKOrOWu233kiHr3vMvQBewWnbnNUYR1Xubxhh4vaqYtzaaQNjLHYHzgDO3SQcOfL
0VveuCMWqBj4uK64AKknN97Lvsidk+VG4XSCIMZgTfkxY4G30RLHFk2f6UaPbn8u
DVw/2vYL03S1Ulan7iPrwY6WiRxhf9fGgZlI6hGsbJKe5mZS5pfn9MVxAA9d9jX1
HLsJf4KrWMaRnAMgl+fHfeqF935Mld8lq8oEIj3HkpNRqyr440c/qEwQBiQ74YKk
J8T8iNZhdukZCmjcktmKJ4e/7QbHQE6G4B8+z/YTic5pScZvu94uwSZt2FCAKdI3
GuLA1kTgVjXHwOfpnlVmaE6gIBl6USZ8w4ySOIfkx7hSqZKHcG2KxU7upHIIxxgs
ytPLEaesPKlcQYd2FJpULZQmHpA+6dqo5Eua9vUvROy4QCCsgxxhmCuwWGtKI7qg
9RlZtylEXSPCwMlm4tRgnWQKrlxIbwvJ338Ivms9d6lJcJMfbQTcV70qyU01ugsc
CWyk9X6o0OYjdW6TC+nLZpyu0kd0eyTD4cSxNhN22x/49Jm65A7YKqcPGVgmOaOR
Bjfn6W/sJ2+7zwRXBaprZJWKKwsbK1W56EzKQAn2ACGKfx6w9wIAfcNERjdJRu4n
IzKQwo60/0jDyVFURvpsaVR/lTGxmi/j7d/r+/GFOGC8XQCXjEjIe+TDtteBfbvE
pqrO5TQDC4yqqjkhxSCpB4kr2WrARoxTf4LOLHj9LUBCS/2Jc/Q86srP8tBMa1I+
U+OxDXeZgaj3rmbArDkjwgdeBebcZ1JyjHJUrBR75IINtYumgEaWD0h4B/T2nBWU
wRsI8ZCWgbJaUbMz0MYmc+dnfyqVqOW3qu65xIl7ALgflEc2p/yQ7pYEG4cIewoC
Z/FSaqmJv4R+K5yMw90W0C5XGCMOT5+/eXC862tQRRxjhuySivZuIING1VSgKLos
k57ZLEUWXbykTqym81eiBIEEBEcfgQGG4shiIpUufN5fq3fMznIMskF59wh+8Okl
oJXivFBC+KQtn3kH0YYwKu/LtXrpqX95XMoYR1RKD803nNvUUoXvB0P+gakW0OND
31iXLsge0h/YPJGLHiIdu3VX2RJ4+WEHmwq0os1Klji4zEA6rO57AUL8QBUxbUfi
tStENhWjOJav181rUYX4TbvxcGjM8vswYq9jIIPmq2+RmQz4fRWrtZA2d0ozqcKq
RNB+0psYeU0zMtTinEKfee4da7EgQKojF38LunCegSBid9NZcwEIKch9Gli+yojc
/C+ULzhB8wygkTucHpwPYxXxcM9DJMzMOQyShIhe6IS9rY2VIym2O8lzK6tdu0ge
huKlIGb3B75Tbxyc8yjcxkGQy2ZhTRDLvZq73TXdHeftg7VaNtIFLjlcW1gcLpUH
qO6lOkqYWxC84ia6I72KcaguWoaWmAo0d/tfTNjqGDlUG09+GE3xId2P9riDrhg7
2Ly4kQPbyUnuLZG4YPanYLF/gmudj9jdIvnjLQeVh//BqLU+M8QDmkglypSLhYaF
MLEqq2XBlejI+zA/1rnBVmqhvYDEtKd3ogEmXnHpTnayLKN1EVv0f1V9Jw+YLPmW
NFKaUZNWImyr1UaqnDTEEdw324a34uDdCBABSATza4mROEjqkqRF3P/6P8aXXdbe
uY+wS3Oh5UstpDMPbcSllePiayAxMzvOCk13QmnbZF+FAwwepiIbgqH5STmlvujy
0J0ZDtl051HfrUpX7sQkCUC8EnXOpEdiVcTIgEktEc4IPId0ou9s9i3lyPP0YRB0
euGHPrUfugwhH6a/mGqF5fEPwqW4muIJqWKJNMJ+DHt/Eqm4dGkgxCD7xbRiNNea
XIhWTOjDPEhNz9P9/bQWKWimZlu6z4CxXT2qDYCTL9r//iUE44+hHmaZ3lstObHv
JRsofw+kQ1AMc21KZj502qrPdtC3IuoSxaSO7yku4teYJRKQ+dmn/xztKKsUiuEm
H9n7nhf9K6uv6Cvm2GO7zrkVZYEeVFWSDN5D3Y6AKsFh/YrzaXEZTWoe3WTXHqQd
xkbaVRapIDScEo86rC3o7tb6RIP48TIT3Z7hvuI11iJaNI0aRZq9oaSMp+0Zb3nf
8sBEqe0xATMGjGZZUmbnM1eV2hfL1gTkqM4SCkkZe2IAQgESfP2w+6eKlGkd9rn1
zq33FxNAelpqY85nkrHYBy06r0udpzeTkPy7qyhQ8DQ+oQszHlga73eK7Uz8cSZL
i5/5Vno+zYig5cTDn+zrmRSU2X/9o57qxxYubdn9XAOtWHfdpjJs/mApDgggoQa7
O40NTGUfZqXO1fkR+97Im9egGAqTY0gZyEsB6Kz5KpOhg+KngoVAoOEFQ22aBXuC
3iE9mu2AGeF7d9y5w0tkFnvq3ViNjViyJIZRMmgcBogItsQIQuaXC5qcp2MWSwYZ
N2EkYqiP0O6JKy56LtgU6fzjRiADlEXfNbX/WvmPuKnxx6h7PyFOigcktqzLeBPl
QUd2krXgOVjJwayWb+Br0K0sX9OW0OVRF5VZMqVkC6LLS7FVgS80efYFdUf19o9R
Pwl/ke+dxk8sguipLbD2AY3XPCdw+PM5ajvlwRpRyQG9FNou1Ecnq4Tj+7tVAtoA
cMJyhOBwtj/vBFIqqswbtFrmvNcUNKPrhZR0E08NVHgAkQLA6u93Kq0GhI0nUUH9
CovPkMzYwplcWrtapTJMRSPEwl+iZaztaywjV85bGSepp403wbEcdPnQ8zDyxg2b
thLKO6ogBPFwHQYAxLx6cTXAOmjiyGNy3jbo1kaCtTfCvXfGRUL4960y5lR+dvSE
4GoUXMOziCXLiKc7iKhs2HeFlfDSNaxFPzTYx24ISJ6vUuynd0xHa1x5Q5J2HyFG
jGYQBPxAGjUcp/ROYMEHAKCNLxJz50GvINbcIfGgIhzd30fTVRNN1Ndccn1v60O7
0cK6j1wdXihJEMFZa6yRVd97E1rnAFtsR4XfmyUVoD3+Hapr3UnCQrUUvd2osu88
Qg9/E2sTSky+6QsmkYZz9CoHtbkt0avBKRZQUcuwFw01+xpDcmZMT+val315B1c6
geh46dKM/O5FAQjYbQTVYHAag/CiVbvpA5Einx67j6rJ2qa/M49f7V0lktgWwB/r
ku904GGTqn559TSRzXP8vGpYpCySIZcOOkXOiR6fSlEp1UoiGKeR0rBBl8zfoEHO
X9NFEIQApubpVWlxevo34t/AVFpK/gvlpUc7kqGfLBwRymuUVRexty1VUtwzVBIt
qUixNJrCRp6daFFCZvztpyxtdUjAue+46XBsvra60pPQmkuQ4NMjx0se4WJxerZR
wqjxvMV50AaD2zDgBxDaaEmQRzicKKFtqOYmOQDmfHVlHSK/lhlqNBBQY7S9r8JY
HNZfniyHggPvJ9pGgZFEgkgx8FxklZ2Eo/YeWnbDNvY1hxK0LDWYHFDly/PuTArp
MTZz5zoLcwSk08MVxvLZL5nSeGqWapKqkrL1lJQ75arhdBdLEabrEjyRKV0pQUdt
yrzeTEyGJyr3SNi+6O7+YPQdxOB7Pn/D+z4jxaPPsIZwfY7z1nAvwn3qyIMHWA7y
kdA4Frvk2DiiZsmmw2qb5DpHjxEnPkFz+iI4YNKoKQuZfnI0APLG8k85TRojGRLD
vR/0RT4QTOStpiwXalB3H0rhxigAhV2+JNTms5mxM8hE7SRDbeyVygA0Qmb/2n96
sI3pAym+Gb+a0qX3evXZDtsmDGwkXN9zcAFKpvq6+mWZEbO3k2yGeCxesw+S68OV
nFHlz5riR0qRcp8GpErzSrfGlg0x383ovhBmZ/apG7lbU/u2w2rnTllmwVE7Mv5z
HPpANaAUINkBFqqxtdcOFU7gz92a1Yv7gK34doXNEfnsKpKUze5ps3ykKA9aehLb
ducHbb/xxnHKyre8a4LkM4S+tmBL32nsk8bbSkQ2qnqEy4lWgqnzF8wJUs1rBgIg
dnxX0MAbVPS4cCeTmrUjI6DVFJBtMSAMYS11icKv8w025orgNLWo3aGvZSdBmplO
BSNYlIfCXpzTP7hXFfVPAgAUDcUhUBu+jyo43sjiVTKds2/RK1vfBumEBLRJJTQu
DRxT/+0nxVqBPrFvykbySPV3plDwzkY7Hcz6IVVsU4oOC32aq7YRXfIYdwQnUFhW
w7j3lazX9KOarqZ57a6nGiRDEslMJIHTZ/H5LfK1uk8vN3SyFpAYv4DlK10lU5Gc
LUJ50HoAd8BOteqS4lBCJ13fQm3uPrNZaGq0qb92s0010rIx7x+hBy1p7ojAA2Mk
6Bz4mAnLNM4TBEVZPBLs0+2gXjZ5ji+0sIdARZttmFawiQVoZ0heMJg90UI5oRQY
B9Lru66cieB1YWgt66P8trkc+JhE33LjjdCWhjSTuFTyA3gsVN1luW+xr0+hNOcC
eQe/tqR6Q7Qit8QPEjjU5CnDmvFcYr14/25Diz51CD/1ZarV+y1AIMKQ01xKl5Hi
mluDrE5VSL6tIpFW1fPSb+9Aw1wAIKVm9QLJYqFcUkBgvQnDZvOswV6E/6WdpFvB
VMPt5h/ph+I1PIDER6nZoyyehgXtnr0u1x81QVhz0qUgiw6In8RDUBOr9m6KajdH
KT5iNC26+Dq2RcIqV3h0IPGhC0IY30/1E2Fh0FApTP69Moirt5vbKyziZDQkml8t
wQLPkJax9agnDk1KdAhfxiM8rgsniwojxJUdyPsn+mDgXSJV/GjHdD21B2VExnBC
dYCRYYYfCZW5t4M4YDfrk+0Rmj+6V61/Hty4wEXc8LbzJ767ZOd8UU9gfhhiBg66
uFXrfKD5nfZFA1FSUPG87DyuzSVt5CMBqtFjoFqwmghkWEehBNrCSIs+V0xnUfV5
qazQI92S4zPT65BlUzFSNn/MrVLbhqcVgTlbRjDYKTkgHwzSR1pz4qgFdISamrKJ
M77TmXfeIdkIQ+S9V39g6IYWAaUERUJLZ5/mf1oW7e72vMNSwA8M12kVSLKB8vc6
NGNjpqJotzEbmvxsWrluQdnta1BmvdSmO7dU3kISev/IGiSkz8WSAe564VuWzKrq
gHHosJ67mUw8Xbm+HW+KitHDhIFzacFm0pKMjEZDwjzPSx7Yb2YDNn/39/yAzFSN
BwNAkis4h5FdT9hyL8m0txXjxX+YokLMDc0wygpHukXeG8BKKj8LzSZP+V4XEnd0
6aDHCcmkyyivhLtIdm1QuQLiTvGawRmB0/CvbpAe30XlqlDj942QC4xeEBc8tpFk
d4APLu8lSwQvYb7DhnnJRQsmm6uGBuIGtS+waJ/43groSCr1u7VKfVoKOFIiUeJZ
zUpZd2RlixVVvsXvN83MkBhv8YhhzTDw7o+hGmWBpBWP2kl8BGeRVfaL/LbljRPx
25+jDPXSDyxB+apbWl738lcrJUwA309nKDICxD9GeVtD5fferMSURLAHsRHX+OJZ
lYZwq5QUiHYWGu0H933wlb7rIzxXHDgYZB7B6ac9FFDnuvhnrW8wgOAlsD94AYTw
9eSs4CA1ZZEXsN3WvZp+Mj/F71iPtn8EzlTJd7ZZVA4+VMAkMHezKDMSXeA09VMO
fpqfNRtptnRliup/4PrY0j/0/VVqLIVIL6eVYB4xgd13h/ZDP0ecK6+aRPUG3eRA
W53g4PmwELPPIqX0+6qyQR/QEt0ky10Q9y0sOTpcjrGtV2L3hD6eK++YuDIETgL3
abGjyJrd3GKSoQXlOm9DAlYWUCs4tEbDqIm+ITsXbsZW/45AsiWRQxftxHaKFIsm
AGxZmTr0vNus4EobwWZJw653IO73eJC5eGid5luNmU3Q1FGvovUP5S31KdWXQR3Z
jEZlZD5U9c1J/vb7tBinFj5FXbBu8bss8Ed9YOW3sbLJy8Nzvjho+TeauEeNJoGJ
Vq1CJ9+wQGhNTAFZn2I2Jb8vurOY40JHZHVmvWlWCgNUJf0K7d2yWgIoRfH8tFDF
W1RB49EqfrEdpfbxN+G4b674L62tiZx9rnbwEjURxpUJK6b93lwKg40bZkm1qc4H
Cbe1ek0bFITOhawy7s9f1MzXTVuzUA8SuxKIyyb+XPUa9F5o6aZZr/9sC9xoYV4s
Z5T6UgK7kHPT/jYUVXqaWLbzpVh4/KLb7Lv7e1KK31YLCmOFfV/fkZgw8HRctPXF
PCZXkClrksOoqR5Nh59U4gxIqw8A45ZRqvqW0lXrSeq0HW0vIgubnaSj6xVMULMj
0ht85Ayp64VlW+JZkHPitoCitfMsbWykQuCUNtDJIVVSS54MizkDJWbhHtDGHFB4
Civbi6nekMeY814wGS29Mx46zQxxsPpaFwlecNWuubjPsA1fjSqoG/Sepy0EeWdT
kau2rPkLvG3CeTwREC5r3BsDXZgxIiaPFlft7I4zWsMP91sGKrWr1eJz2ERNmOPf
HcggOb+WUQTxLzYsjDlx3UmKqTUALYgKjE+t7uakNvA4X40+wfLaCToBgkV7IvY8
Kso7Q1tx0d06uAXI0/hODhidijPjDFP8EUecLUUOl6dUzboKLTnvLBPcguaVl4he
d+8Dg8owh9UnD6EAoZqk0/sOA6BrIxFWadaZ4RMertg0Ukj4IA4XvRQhWuy4HVKN
2X4odEwl4JaDUB9eYo0qSua2p5VJij5SIbXzP2A+6EZeAUXYQctt2tyhVt9chtsi
7etcS9BxdyLplJb/G++3SawV+bWUmH0m50o6aM+xfSTfpBjdkBzh+DPjpetbqeKv
UpehmawX5j+hfjOIG6dgJWcq4zVEWKEQi//T0MuLNIE90OWhVrWF5A6cuOyaAtYN
kucR0a2ekHiiVafd5CA6zXMXR4UEfsmDj2LR2ZJpz38oxznUBXE1FRBhe5fSg8S7
IJgdUQIfdZEuk3nx4itpshFUYexN88mn8OcjDmjbMjN8zMW5hGi5BM4zCDCh+CD/
MpOg30nIJ+OGA8KN090il4kGbK3APwV1L+YdivmAOjnzW3VlAjLzaSDd3PclFh9C
jLNtrCcRKdhCzpiD11NdjIVmN15OX3y9RK2mmy/K4KXXffKkHJsAyYLmQp0FzaE6
s02jbBuYcQbp/2UlJ5bFAHAwGTVELB1jKhXxfH4RPe/TNvktXEBmBttjsP+dgXgp
X+oH4QxGkpKdCBijKWL/p2rXmyBReJB85VIFt2sWJGNKed2xUVQrZw/xDG28qCHb
AxNl+iVAPJUP0KpJZ8S6NugKBjrDxFWlOrkAVkZXopySpYCFxL7uU7Lo+IdU2EGV
OFgoEOledklmVEbUrY2cHcqbrQlu3g6N+EH/qexqWwS5siorXa8IqDXg4uFT+bo1
t0SOcj21TabudXT8xbUjNx6O/gQNPbTKCss6SR/lcAAsirMbECEtG9Vn+WuDhzmr
Vb6xgBgER9vUzwtq2BggeiY3lxUzjOdm+lkZXRYRg0hgR5tHrFxqQHoX11I5CsiL
j5UUBRaPSY1siRwDsXd5WEjeREytGNBVtlsnAfDZn7+hO7wPQ2pYJVFyjr7urkom
lDmdlAQvuAwmehmF/k/a5m5rt3gZs/YIYCzVJdzwVERZICDWHZdIJPKg3vqOIdBO
vLkunMZuD1IU1U6wkz830vyJzg0DoRq2TycTiBjsC3DpQTXY8+KSUiTALU6itKbV
ibF9jnWuudO3dlnj7fFO0rwVhBAn4oHuMxkbqvb1viLeVrs9qWnHwdm/9onfiAEC
lA/YvB69VGwRRkM2CKiMCnMJwECEOWbSa5PUSG0PB7dTu7pGM6P5RwwSfqeW/4a7
uhSKMQq2mkvBvy01405lTxtnKDSEl+5BGtVBqzVoMdswtTM4pkuKB8OdsA/V/oEg
/ONOA9aQAbyiJXVMYYiAmaO2j81Qe7kZKM/sGU+q3PjaVgz51j8iMHScUSAWcefX
o1jRdPwpYK0e6su5YWrGP+T2Xu5gvO+ONsZlAPJdArux1nrv9lPVo/GMGmlUSSDy
50WmHEjuXpSrDW+Ec84o9YOp24gZJ2/JSUth6PWM4mJm4ByyjdyK5p/acyjw+rMX
Q4iUzIJVGKqC7UIXyNmvIXy3VHhjnu5A/ZSv/2jAGOI1Zsw3jiO4E9Ef0nPBaY/m
poHAPZyefLbKL+IduBuJCwxsjSTM9qMBPHriLcAr1TNgKQJR4eNLG8dDbtnHKJBX
vG4/fw7zCKtCvU+EkCI5QRCRmj9agost2EIlQJpwysu2ICPlLzSSAF1zNNnXwL2B
D4Y6uL9/rBTDUojKGavRbrpviS8SB7ZU73p3NOga7cJw2cvUyI0Z95Mhpv0E9yiF
NzClZ/X7fwlrs7tT33csmGOQLXWmj+BXQzRJvWx9kmXanZ2vxYZ1ak4TphR4+ijM
SqHAeo0GPmv9B/kDBJPlvuBkqcBA7RgrCWWbu4OkLH9r3s5Y4l4EPStLeg8VH8OC
vQvZVuql+WYRI+fcbNhfrm2/qF2KrTMXGLbP6fiyVpdCub+ttAD8OEKIHqtFlyOA
kk6HZBuIpur5+mApqVmKzKX7M9wlNcoQr0PkjFEwaGNp5mbw8RAtsLv+aFtz5dLe
AIo/ZjzC48GhxxChotb3PPqRyOqr2M3w9A+IdhztxWgfimSUPKERoXYSUu9KsXCD
+fB9q8kv62GcLuG1G0/X191ZaSRAM7dA+DA8JLPDsp6aP8tWAN9E7zUDP6/uoGmg
JSwOT3rj3quurgHy6Wt1nBULsqhV9zMmN216yX/WdMj414Oy8NwsmijSsFnmxBeg
sRMeaTMDF2X3HLH9756Csfcj0IpV1tCKGhKAwGrcr3wRVnwptR2hzxidrfQzbDli
qeUE3r0Vc5OA2DJAUMHTHkEnHXCxdGpjK5D54C+L6FNbRrLih5BI5dti3H+z2/J6
RmhmH79TLwzbqJt8mIwTHCwlqbdq6h2tr0gS5uz31YbW8hT+JyDNSnPXjl9/8ckE
YUdSAfeNQu2wrUcAH6OEoK7qsTjCX7+G7xPSILDfy8wbSF1rNL5opENYBRETJc+8
VoBXlL0RgF81SBrT2zy4cjxVMIqXlqagoWPvgI01fboB2G38s172WXu04QUwIfIZ
+j5DF9m6KjKoxXhU3RLrRUqHzWGiV/I26OivH9Cw9pQBiwR0xZk3wMsI0yNPd0wM
SHfeXkdv4TYWahbI7TJdjVZZlrmb9xHpKtkrN4OP/GUfXTeqBpoZ64PXwNd44H2A
aaszNdxldPwrD+z3hDb2f778vHbWl091rIJ9V0wgAxow+5fnKv95YIH1F19JZRlr
Jc8GOn+6my3C8DQaG0hF67autYcMcHoxKLwfT/RW5GdH9cEiHBEFOBMAAVF/sdCH
YngMzIyXpFs9+GWQXVrcWeSASN6R9sPXQW3m24p/Smzu0E9a3lQ9Sfa0fhIsDFyI
cmeBYnPI0OmUr2+h1gIwQYPhxEumVxB/JIZuqcyHWreg0ko+vaWALFj73hu442h9
HiZfWfOT1zPLLOC/PcjgIvXGYGBJllGZT5ZMc7Q3Xwaql7ROf4PIL2q6xH7yDpMG
isNYmKVYy7Dehv/l0g4leakNP4lx8m3UhYUa3LOpVbZ09s4G1J4sbK/249YidNPR
H8bLzWjdYyQW+T5+yoU5I/xHeR1JsWYfXqSY/zoSxFL64FHV16Pl4skdbt5zLXTN
g+xq/J7LbZU/CN0eoIoY9mCFUHWY55lMNChaT9npwYDrHcY/Ko81WDT4yxSwKL00
5Xq4QF/B+9ITfh8UQGE4PYOPDANxyLVnufv4zxtxPcQm3QinLHIky7cxD9T0CV7a
x2G/JBU/u7hKdhPJJ4nKIJT/0ENJ9ZItCJNLq+asaxoFCC4jUFzsRtGtJjO6rJD8
ve1Y+75VtW/cLF81RZEzxLNhCUsb1YwWAi2xqdnkbJysvVz11PLHeaHYaXaCbbyr
5YM9eCIwuwXJpd1Pnm+x+yv+EkgEDCgn/lQUlxCYh0/q0xlV8ypvJl+XJkrqqdCh
UZJxGbJeJUY1SLuQVdnsDDz7nRIxZKir/NbmfhS/ZdTuKBxySsu/7caadtEZJmMw
JQfp5oZ3loo0E0k6Ff3D/FtOWE14kQqBu88zV9VG94nQufZU3ZdM2IG8R23ylfUk
Z3cdicDHNjosKO18ENPlFWN6DJRZCs6nkuJr9QkAt6NfAxSA3HVUwSkb1gJeFzu/
ZWxfU1IwWnGVPwAgNtV4b1+QPHiv/nkv3zW9BN7VimSbLABr5vuhA3F/Io5CUnVM
Th6pV7FxAFbF0Um2gfTPXCq6ydir8BcYYo4L0TepvrW8awVrwSb1Yv+f5aHwhbsl
8EiVcswpnaq+8eBk/saTW34wIQyIvr37GplAvT3M9e0vB0nl1qp4ZMeLAC/pvLJU
rtCtEoogtns1coZFYZhkL+T7nucn7oTR137te5vNssR5I0vhy5iY2F5s+2D35Ndh
BwUSs6WuYeCzJIctf5VHJexLdoxnoISYpNFV/4VZS79Y+Tw3DOJHj/udCPQhsJdv
h2ItC6wPRdMiQOWF1m1ZszQvlQAJKbFLx6ijCzHCFSGJoKFjcv1Ge1hjoFZbH8bj
3TBbM/i8SqIkFZkeEgCOwjkkUVnVz3L4kuNqlWr1Y4nHSML+0FFXAG8rmi95CJYE
y6ShDzp+A6GzorDFKc3Jf3Uh//9tV6xpV6G6hyT50uCthwUCetZcnNCJFmOkdPMx
Zbur3Uh0tGnq7khERtMa+rIwsLm15gydiCBESxQMDZDenMlKrvTv/6Yn2IOFcV6z
JjlFqNNU9d74diUeqlL+l7BuD/wH/YJvCbH4qnWpMBrm36ct4QuLX891y1g+kwZl
o3RylJfPMN2B9RRlFrNUyro90KUP7/Y1D6VtonPde1K67iPQPnMlkztS8D0k0RY+
D+K0tXTjyY+AUyID7g0ZvzXmvbflDuYYpubGguo1HgmlQONn6IZmr4usA5C0sDfQ
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lBKRJlTq8P0PabSfpaXFHjSyD8fIBx/cSGptpLiU0q0xbNUodnqrFvZGVhFo5/xR
y6y8LzojGbPLeQZLDddeNrtBqp25JxFzXR7BxmgX4B83huR/l5xHVyr6SvrHPeTI
wmr5RW0Czl9NSAt4n0rl2wdFVe4wTfy20ACb9x0e3Ab0xb8SO1PeLB8VBtZqt3mp
p6mtJSHL7R3jYThXGJ0Wm24BS5tVjsovlywPvte5NsJv+aXnmHCkUJVlY5KwpPhC
rbpQywYtwumcIzvHHAfz9ZGGbrR9B7MTepLTDtS4SccpashwGXRk76dbyqMGJcNu
HcajsP/1AWGLArkLNDHP/w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11760 )
`pragma protect data_block
TjtIYGCETLoRAw4gB86NdVNOXRcNkRnWFqp/LIc9T4nGCeznzQz+d+UP0kddYY5m
BhfkQHjPIUVoDZ7vIQdjH5uS+IFEbh4x4XmTsmSOIqA4Fz4SptsSGIqHL3leYsNj
O6z2g99OJ71axAsdSPaNd5mDxEhGQZSEri8i7NHrzCZuK8xT+t+b9dqnSZ2V+siQ
8W8YbcLDjwKpa4+NwZObea+vVH6TTxIqK7IelY8icTnhjatT6ZPnjjsxw+RL3z2t
qAu+XhzSpzz7PvqpbxRlOWgDTd+3GpmIQtOQD0WNVTS4Ss1y11Rzv1L8T7Efel31
S2Wm1nRMbipKode+nRdJnczqegg/Qot9v4e+wtu+vfR/R0wZzIrbWwTHMK0KatZ4
NzEdyq+523186+duHr/gXqKepXpRSlYhSH0gjHnZr2/6+n370X4nuNGmDROCena5
x8LlHHgjbThIC4fm1u1+V1SQtvu+pwe+nlMo42Fjco3tiNPJe18Y169cqDIdZizn
im6A9LFUiRxOygxM4FQkIwEHZdsZ/Q3MMFKJabN+36EQmwCq9zhXA0FdHJiE6rVo
Wg4RWlTj1ITTXRrNI4ta9vcLxFBAzksQTS3w2w3OhN8lvJS+JjhhcQoHdCkmL/ti
+2FABJajcqqmtGc3GnuLuO+youVaCnQqchQw5jK249dtkcn+ugKyvZNQArfXhnFN
Wab8qLKWJ/4q45+d6PfFmtPdeZER4lXDJgN6XH6TRwZycb3wRb8UhN2XhU4BnXug
xyk+RVJkyZN7PhtNXjx4mrDrP8bqrSMWBNqE9YKR0XSpwTTUhHBwdluZ88FDsZG4
xJCejOU+613iXa9EXppuv63cIEC8bvOA2onP7hg+fTeNuzdL46dAFmT8lFCDxTia
FblGiSkNP8ATw1HyJzD4Th5buTjamgRZK1VFRDDHFiLqMpjCdSKkkimVhhJqLcqT
1qr2IP9/gNdwu4cdEwbPM699tXBR0C2zQGQYxFMuz/JTRl+2CIM5iab+zR65Dc46
Z6wyHbiMwtvCHGXRLvq43rHe7lZ3FokXQjJ663QI5M7ghmnSvS/sPkXb14q5C5Oz
cX2wfKKei+bZTKC3dWrTCGqFmBxo7WjtM4e4UYZN5dJNzm37OrroiaTRaf0Cb1bc
drOYBAPgZU+GvZ3tIh/eE5C6Uqzwtbbt4gzoGyGtOnO0JniRtg0yZyQonTswp6oM
FsshcnJaNiAhuB+FHXskdPDxSbG5fJz3DJHhi/Na9POWPCqI25q/XstwiMsrx0jm
ztzA8MmxGGdMH+i0gUW115345psagEHCMTxq8lj6UyW/ceUBZYoHkFGhDjaKxkIX
74DeH4tBg0GRLKAfLjLRqTh84Fu+XbWgbHbh7JrpJa+RLKyeeNmhghY3jIKDnbF4
IRe9tkUGQStJG4DdXDYaJMlzSUI7e+HXT0Vk7cO5WY/gt+VBE6+ixlqpI5Ecvdp2
uZgZ2VoFZgWSX+LdtwJfTTOp+CVr7IDZun1CUcqaRvjRs3KIPD4TNp0hbK2tHEhD
LObuTr989+VQOuA6PrmX23kA62HZ7JKuWmw9qGXhLn4AbCTM59ck0eUWMreXogiy
oMZxESxYBeIbvCY5WlmVrhwYyfaq0VTgHnyidSyW2AdUiNWO1bufPsMW1nh60jIh
XgFCdi2pLlOtyZJPYNuU84NzGfhe2ZS9RTKKekaYKry24BSbprkUMSqrF2nw2lft
mPnVEHv06B2GZ1OQjZy/ssQfmdi15KXVUjRlQm7m2ePRrjqtvUxC0sIH66KtieWL
BJUX/dZmR1Hig5Rr//QKkfiIuX/MeUsAi5fuamKWmrsEPNVFkSwicGOLr0vQR11p
nJNLu1KkZijViZAg02kxniP9RVg8k8zUP1YmIYmOygzAF40M5qaaNKTSyBW+Z4Z4
YbTazAMGxXAFOKt3xp2rR67v3ZP6tJs5PfYlRjZydC2umhiKss3GgnwKgNh2LYlI
i63WJpr6hPyBqUWphjqlcPO7wSCdkhvhXh4spgcm+dG/suN8OKshvxxCWLRGmUTi
ziHDz2FbK5hW3x5zGZa6VEpdydQf7qb24AKfM1FGQdzdFfmaLYzRaaGE7xe83uhQ
bUtCf0i/eJ+zch/Oro/yD3u+CAm8N2m75yYrrZiwuFUyjLVYlPs6GltjFb8M+DoL
uE0nZqO72aevKGq7XmV9PfL4vqDLjfTbZyzuNue24jjhyw7BcR3TBZCVMm8rbVxJ
0ODIZwxUPVbrHy4azuHG02uZoGgNsBm1UZFWSLr1A9MjjOThKoSH31RgF3FdTMhD
BFufLF51G9GwflE9vHDS8mthVkLB8lELJhNeP0eU/lF375+adcaIPJj0PC9J+DTO
qH9yw9O8NJnKx4CphNbimx6zcB0OcbBWT6TW0UxY2bQTzQmhR9BkvmZ47YE0/1wp
3nAWLqvsyK6hmxZJK5jjt9jPA/bv9GPxo9R13BsNqSd/qni+kToK+MyWQyN9cjTE
NCHUdXxsOvpqa//JcQf4XDSPNS0d6RA4jpqsEN+Bj+SnbS3XMQw/bl7Uq6kPF6H3
HEN/ref5QEn/neWzmzUzjFvgL8Q1IqLNKIeXKRA6EXP0chXUeA4rD0dACqqHLUlX
e5kIrBg7/XUZrSLtdV1Fgu6iM2NGLi/xmIbNHYXhD7PWNX6OFKJi1Zpi1cdsPLWC
j/ctUWkPQEcg1kLLOUIPyKapuGwbhFAr+Tzxm7UlrelrTzyG6K3N6JLoTsRgVVTs
Ged9tmDxwE7jF9P9KENma/YlmD3mwaVp+lP8918UHg6RupZMWp+9jxPvYoz+/O8L
QqzjwzHEfZGRhkazGZfmwrvkw7T51x5cqVK945LzJVs97xt8fhNW7KkhF+DJWfrR
0Kh0HW9nc+9NSyuxrs6goV/Yv1Cyq0wQZYNJ0y4molVSRSx1D95CUCXT85azgKlk
r65rHYF7j+TvZxA3bZMRvqm0wfkRGCdStPtBBqcwKom8XwJmo4iKSfMmqTcVy0lh
O1d0kGz+3Om/ogLEdOmyPFePL9XV7s53S7AOZshXOEdRarOXmWzsqmMCYz6sScS+
28ue9wba9R1xaNgE4hgtsdntWkjhFvdwq9nKeAEltBogM5Yv+CWOZGMO3T1h147w
3khllXBiuZ2iRo1dXXmKYGDZt0aa10t4bgo7VRMc7gAjffB1S8GEAqspqtvRdHu6
J/zJ0Ab8lfNjHPubnfygha1GlQdJC/FWL1/RkRSCCNudtcIZ7Mh3JiftqWj6SI8y
MnaZJqWqbkalyOxbESuqEqQiTTxwgy1AuFaCREEZk/tGbOSXqLqgg3sitbPZkGlc
k1hoEv2ljnIbjXsNL6O3bKuc2gbNSiuHOTjwE3RNtDciTp+eT/+llVi0vXbsBd9H
YkE9uB3AczmtPCOAoIy7okPUpQpS/62LHSLEx59DoqLxD2q0SiUfjzo7DTn+UZ0k
DjzX7pc4q0nbPO+321JHn+8bk2xFl/zi+vrJoEbHzKuNhbj4R3Zz8bKTzaHlpIX8
MT0iv6tFeSFy5ODjKDnMNFM7zodT2foXMtkQzjRnCdetVTkyy4idak1gXarA/ucd
2MVd799bfLdaJva1+ek8/3mjx0rmVIrDzWHqN9YX7CnVwf4d2PI1UMNPYKswRxEF
Km6M4Of5sLIWDox5emcYh5chfDqg/zWdxxIypG+48iUmaZ1lqWerzELsMaxjdz7B
hmMlfJF3icQRmoaMen60OAE3gq6LRePpfj5WLxVwbrLctTrI4OCnpeFoG+N8oYs6
tdF0G1Mf3RFs7ivgYquzMdN6/uFvQ+qPB3MgxHuG7WvEZK8cngFfvm1HhPXx1u1U
XLu3ULttvuo9Eh6JFEhSVuJopTQRIQ1gv6N1ObG4B0VWGc5pRXQyvCU0kS5PkIXj
n17qxXhDJHTva6BjRlE7owGdJN6+YJEVb58ZBvffcvyFyF/lmv00S65qMsam7Yhj
BePM2WW47lUp50o8r4RNQ2X6FNj3kjEGOoduhI/Ku7rg9/7pBF9Kh1g23q+yDC/f
COkSb859F3vKgLNerLOAE4F40zs4gSo10QKvK/aUm60y2m7dPEJC/D9Q2hLTNyr9
yaC5ObH1x8FrSsQdt+fugq+oLo1NqHKiT5XFK8QEEz5uWAK+cmh4QKWg42gf+1Mi
w1GrxVDNWQfo9EOdnREGULzGsze9AtRWoxFZh0cWdDJ+ITFZLcrUI8F/uXfOfbV3
TFHSVIPVYr8JZJuvcenX2+mHDwuVSSnhfHd6vlT2YC747exzWHG0I0ekoYlQXRCS
lkRtk/7MBIk6clJfQpM/Bg18WB3DmqeByfPuBqPpJVh2ORcOFOWQ0KeGZmmHvLVB
5Tcas8lXfDhEpv/faNApdu90TYLEQHAFY+qYI5XztdXnQbrRdhChH0h2qqjyVPpX
qeJcm1XBAp11jES/aPLl4D9t2yA2dtacd5G3jFmYKsHFRzFP7tvAC6o8euDvyKbH
V9ZhtvAYmM7NpcLKQ/uY7DMTv9qv3WcfOmOmSs5HJpLeBFO1O/ep1HZ7+v3zXHNN
tOPUjsq63HYZngqOFXLVjrG5m17NOoLJLllusgDlpsTPC/gi1N0IqDzLIHIXFxhd
omNdvdxlCenoYvHjLvHbOj2HtkQ1EpuHBd3Lcd/K+YfVepMXyv+zKEU5ebCBNXHf
VCgw9vhu6mqTw5gWqy8BeGSM6C3ZWaPyVjelRRh1X9ZKK32viYMLljM7XSxHgHV9
uQ/TOIQI0pANPGPpORahuFcPZpAB5/mAxfLRxKA+h+Bs1tbHH6J4dbSQwqPZ+e+Q
Qt9Te1PDNEfmRU4/GUMQZkPEhEnzrHAysi6eUqChmXQmd0OkgwXJteqJNjHmBqDc
yKPabzzo3wizqDsyq6pcIZI4prPzxRM4S8oKD4fasdCcgQSf/bfywq02zJWaqo1A
vB4yHG5c6Dt3plRPz2VKxT0WK3mlHV8XWZFL1a1/GvAedZ3JiQPGfzX7iP/ZGunT
nlkqeVj/9ALNoqtnTTsS/Vr2jbc6ALuIe/U6lSxhirA9b0PArrF77MRUdGKQ3+Jr
LwbEMj/WWtHuOeFHrjhG5N2SzHYoKXuFylszgjOCcTPiauhVAiFSDnesdAoUCu5L
A2/qQs6yAJaqaJAJlEAQgzkQg2FS+Q6hJsOK9IjqksBFgB4vYDLhSGZBwswSx0+j
eZjbKKzLHyeVED2Y/8+GeHzeVZqBmNP1avrtP/eWeqbV6omS9HH2Aha39quzNZQN
/MD1iEZ8RxHwJ3ycS05KML2iChlSJ911M1o3oyXyKbMKwwj0BVkV1zTy8QKirjYZ
65KopTHGrViSgnrA2kNiphf4ZgOMUtYn0LMmGitcGFjS0zQyHUNlM5lgPwyEEp1m
ExgYkR0u6/ofVyP8XufPBXsebj46GwsBIDtfx+QULV0GrSVwZCS41QN3nq54QfUj
Pnh2BvfPyeuNPiGwgXsSIRdRvxlA3Tm2WQkV2YsneQCuey0XgGdWoDQmDrRBEA/7
eBhfZW/8XTk3uM59uvbwJFDL/2lJFT1IoZMmpU9ASGmMiiElp1dvPlresEBMmBsA
SEZ92JgEREkjppacejuNB7pKJxBSGP9Ks+elTq8FVKerU9golDVA+n61dlJzoUEh
vb2StW3pdDLngptcEcoYoVgVidckc4nusNtdfK0ng5c7P34J6A/UQ9dCJpkN4NdK
dcpsfBrzQPY8jnxkqGzufclXHvUd4Y2Md7/aOjPspi9bB1QuVivwO/jTVj1j5Gv2
oQVQU+q0+A1Am1Id092G6xy0+JpkhdOk3VbrmHqAHUF60KRHkWTbwv+bZWePbl2S
V7kyxGNJFoNBT2pGx4Asj7ZVVGejamHHll/GfD07RByc6s4qqygrsCh46/ebHlbF
/NRheZbSz2ZZVOcb6fIFFx5IUAVawji47mbEa1J/sh2uS8FrVut23HJyKoT4QjD9
gCX77IO5ggzz/k5CK6BpzWi9g3850r/frO8qk9rfotw2/LEqsvuDzESELtZS4N1S
DLb3ZKGLQMBIsYqOvPGZoS9gEAAfJsftyZBm5OBh+O78FhGzC6cpjn1hvSCdp1us
f6qOyJOOsUa1RGhReu7Atgqa3II7YPU8je5pEQ1jyOBcWRXqWGTjN8ATSEXsNoEo
jfkOfNrAT397OL9wKXkZyqGMKeWb1rS1j/uYgkn1ZyoujzV0q1C5zs69KycokX+1
ssk/er9+a6Lt95TEog4+SJI0ECDZQ6vzTAUCmK0B86TK+oJrBGC6LRL32Cek872I
T8x4YetTj7pQNA36GW+UtEx5RI7TjIkfGmHA3qZGZp5F1MQTkkEm8pZiPc+2mE+Z
PVkZo3PcSIP6KUnlj8d6Q1wpQ1PC6CWrwWPBkq3xDWDEQOZfPvVJs/0qv2aXbHgp
BS4/P8Ux/zSsiaazyCzfPsxZqRw17wMBV40WLBQPsupksEzmBYpdphZPG82szOWa
jhA0g1xlDEHy2s2FCrIG9fOrLdbdSqINX2Z7Ox700E4J9/aeBVWHBWhpsTg66jrY
G5JqNhKr/0koduSIYIh04DsHvwdL9TcQMA3ZkgerVwtKSCqcZVr4Yq+Gn42NhlIO
2oeG94kUe6dqfQdYnZX1NjBEC/4CMjTRHgn041CFbJb0VPSMT10XgGytR2kAWCHj
CywwFZkOu8k57ts7hktgfvY11V2Hxuhhl4rTjVhCxPvOKN/NFENIv1Jf4RDeEL+K
BXZ4CAut7P3XAZNA6uyP08uUwIJ3KWdxgq9uK7GA+M1qEklvZiJwUaEMvLqly6gq
xgRUXnnnh07c4bWl8xr7UUd5K82CmmcH1BarT5p0qbmcFJGyiMwHmzQFN3Se4NBv
Ck0QITItJM04VFvC0g9Bfg5RdqhAfsM/6jBo/I9WQCaG1XuuzoHAmJ3JRCu9NWGK
OGCz6IYtZnrun57uLnqktUksSrq95p0fWH2lRC31gQR8g0wfs/Mgo0x8BPjyohPH
rytKLg1qgrtizSpnFzrQ+hdRJ2RENpwm472N7G6MZ0PgcMUhJ+ECtF671Xvju3vW
IPGTFNFIJZ7eQt3mWib0WecZ5bcvVMVZLl/GdY50cqCZ5hc8N0WS9OeBztOsUMC2
huL8FgkGR6Ou7a9VuN1aUDs+3RCAe2Pmr5LiTeVy85X4dgQZIHgIM2Kp/UbAhMMp
MrFLSUTkHUOOK5JHfsLCAQMfgdrXq10DJ/tOAf2KgMkxvRxYlf4Od1poCyjs8JFP
Yd4r+2mc/8A9tpg9raajc0iXuGYx+M/m8wNqMG97PXtEE29ljrdSG34gvzBpGJjO
hgT8J4GSu5EdhMJ8rQhugA+v5XCaWONZskjLFAPDkAbm9wUF3dQVqUp9cC5e07lk
A+CecoJoGf9U4xNyL46LDvDielbPhyOAwJDexmBDyU7F/2D0gWhI6VEJy4n2/nts
2lU4Cgi8iuC/LQEjPLZx2WT0fxXHDYs5M7HAmiy/Ohz49ycohvMciOwTjcFLz09W
4+Q3tkP7P4AtB7toCCRENwJRbkICayNJraJr2kQR2HedNaKX0Dgn5HrW1Qs0vnoU
cLErhuIEwEUNyxNuY6WhBe/zMorRC61tgQpQPVdqL/o/Uz/vIC2KrsqC5WykWL7N
W85a6XKhh2VZKnsxtdH9uf6CSVI/Q19LblK8mmg62vtcK8hea+ZimSVpBNDIGA8Y
g46JO0jl7r+oxAco1NgXzEJobs2rCFBxC3Ef3bm0NlYhBU62HJGRQqapYlaOLBbI
QH9oGf3QKGvA8+xMQfN/wM5IwVAYJ2QMuIW/vcGplDrRb3TVxdtbnECoUGCOoAaM
NY4g7ypUxkevMHhmEG+1g+XmmPCC9EJa2GPMQLcAYNkuOHIX/QjwofEm8vbFQXaR
lrhdKBBAKnY6maMCAk261fd3kCGrIxe4PngJzBJCgBLCOuNftnAFoOE6aVL2EG4E
LA+MqSIyAhVWEgHYtRQlf74p5UEKFaRFtwEgKoBS8UhHmTOiFbpktAKfdJ2OcKbW
c36zYoisFDwEksBximF4gChYhDQqJqTpBhD5YgThqS0Hwm/WvzwJzGdmVOr1SLwU
HG0wBlfqv5IynJBgAM0sO1M5TXataCE9uWIlblqop83J8dsLWEeISi6NeJ0Hd+Af
E+tgtLjRLbbAzbmwrVn4G/euCV0AFsVTUbBH9/3YRLmbRCjAwD6wANnu1+X2NUEr
K3ai31c2R+MMEVWI2EmXdWcD+GwrX4EXa1qHhhyShE4dEytgb6fbyyg4wIZSbgTq
faHIWW5IjGJqCX+RkPtDK4NK/punqIVudGXVN5zyW6e32nLiV8okB8PfR0Hvkkw1
LPN84x+SnKiBrBDQM+T4/p9/7+g3BdZOL8bucDZM8uNi+pJPde32QD8VDhqY/C35
DEbRPNdBrHZ7TSLxIRcXrdx4clNWhX75RnuqlCZ8DQ5fjjQB0fvZH0zWJopC07q6
QwDpkgxOsw7qtrq4gG44G+engMaE1B9BCbwK8V2KgWhYBO0GuaV0mUcPB0hQBqZ7
ylvuT/4ZlWQjsdQcPdXyNiDYaV3R6zcnNeny8bDbEMfIAgUEKun5dBuSWWlygRox
qnM+flb3kL5Q7QVjTVluJZZUYy6UplA5ZvLTv/CWWj23AWUHtdVWlfJscp9tl3TL
D4EsFFXtN4fK4nL/G8Xc+gy8rNiORLhg52cVgT4cEw8akIWf9esz3Q9lStH08szK
S9r7GD34zPa4xeFMhwhvCV1BihPzM/oYei4agiVJPUnK36txQIzZDt2BkRJqYq9i
8vgpH/ILvUZGBS+fZp82bc5MplqmAIPec2QHKne4Wk/AHftPcFi3vD97V7FF/Fgn
HhtcNHZM1xjYlbTBY2nr19zSduR5KEAJe6Ajtl/sIMZuFlI3xTk2wKombBoYvqz3
uYOVhfBtEvNFdsbNr2/++yoAd+trXY2PrhdhV062KfANFnuVJzx5w1vt/ZA53MWX
uTa0C8N6bkEPPIl61pz/YtVvY1s/l7wcISVF+J3ZBAQgHiZM7K6kG+lPvFN5v+QQ
exOwF9i/lOf8bphR9LIJQNrXSUe+abMc6+jfMQawtNR4HTxlfP/8AWQK7yhsGdyz
0cNF0jg5AXNeiszq6ny0J7gvwLaZbAKaysNczsYjx/pavKugljc4Avq9N6ab2ghP
G73/gnIHTdcYnlp/Bkzv7pYWsvyh8lGQ+iWoW8Nk1hMsqLoBK7slS6Dhk6gGwfyp
VHXJKV/HE0bA/7mTLiLmTM8bWnK96L05Er2PVLH3MZbklE33Eqm5K95F5cc4ZW3x
FHPhDJFKS8aL5QHZX3MtEiaPIVLS+zBP+s3SEDQnEkuh23KhMDDNl0qlnyJPlyce
lqJMEV7ceoanSjeNgARPGR5Ypt1WyggQJdZA+4d6LWbGjviQUkAUd8tunrN/1Rby
DZVx1E0nnqbDBbVT0FILaUIhU43q1cYungFTYATvuKjIQPUEYx7e42RJkKFY5kg5
AoA6M6okz+Lx//HmHVty58nwJv9RpbKdgwY4HK4wAyixm3alfVekguxzCAz6H4VO
afyEuOyhuhN+o85Bpre79mjSKII35uykt1qwbXNHv75P3XnglThOPN3qH/E+I7Qx
V+TZtarCe+1pNNE4dNVKi6YuLnn+DcGVReCfMBPcFNMMFs0CTPZatm0WCXWt3fLy
bjpztSwFzuPmreTG+hSWZ8QR3iiUU+jFGdIOZt0SdD7Voc4DkDt+p6DqUx3p0Sbq
zl+z3M0fx6/I2T0y09pQZ2Sqr2d/rX+pZKtenwWWznVRWlfb45DqYjiX8LKdNe/I
B5IMSGdsbzbqogsHYeQFQaLQGfl7quPJRFzU1BJ91dLBmXGbx248DVUalM1LREzF
mGsRaLOiG29F0jUcE8z0sRSqqAwIVTyBxi1rydWdjY0jmzQx4w8X2PrDKlrrfLLM
j/QKrObt8k/D2+F+j5fTAyZQzMJJSEoTHm1hkRzOPDs76T2vmkkaiDPe1L+Q1sZF
3qXFt7U0YqWI0vlm6EY13Kk7xZUp0kTD78nEAWE2WEyJnr2SZe9I0hmvHL90BG8l
C1W4hcaaj3ZMelgMFVESpX4Fm0QWCsu8PTfPHgWPQ/TNB9Ep5K0kK+O6bWLSA7wQ
IKZlSKM09qGYhz78fJ6BWhY5F++Z/kddo33iQzzAvulLfGEtjc6lP7u9tI3HPXhP
q8589Q6m0T2G0xkFzfhJhdl5mprhxYWw0QlJ30I8fD/QEDDwHskmTHbdHLM4YvJF
XhT9eeJd0wRcPheeq+3HGKqKGc4jHX+f7sWk2MOHl8PWO36aqu4MMsO8twixk7+n
3qxBbCjCDxDaVSY6gMPpbY5WGfFIhKIvgddbaZZNwZsm5fFK4f/zw+4165fHWxJk
YcVI2rOxZ6J5qzwziYpZUSKKq+vhonEfmPp7DasSNTscFBmIsDO3AAuiIUVmvu0s
O1PPCLIMtwiZpbK8WLuKHwiHSgXvnu6U4xu5HyTDQeO9+CxqDSxB1Z9XhpD9nCuq
V+HaKo0St/lL5SHkWG05IiYRD+w4UopN73iEPRwUpgncNZ3nrjuVwLGSjrj85h4q
F4zGFZmyeJKYObC6dpGdOJ6QK3700GtdDLwUL2YFZGzQh2usJy0dUgtwogCAXxM+
BIIP/dQ2aXxvuc6LLFzLuIciDL4pysQ7nJt4hkr82RweYyhVYz5H3CVy6sr2tajb
TBbI9Zo0PbxJ/QfFr/6Y7Eb82OdF0yiEFqbxArTPAK/IfVxEBCzI8jH0JcaDosA5
xWy8zYO0CQzSW68q4+OEZf8Cpht7L2YpblUjB9KDX+krpD8rlQIvUODrQtCWa8Qa
YoiiYYHfcppKGXbwTA6GQNt0z37FcXiRFNDCMa1sFsRbhu3wDssqafVOjFsrCUet
p2FJW9A0FjAqyBDwZ/+rAqZsCYW2nMQgzQ2oDQ7rCC5s0xxnWXDs6gwyN/tX8htl
gVAMXti86QOM/fuQecTxUw+K9RcoXDwymxDcuR/Xt87pN4YnFmuHyaqpnWd6ZV05
NZkiNpNlby0c18L/Uc3/MzhmB1SRsjDpLMAGeItlKGyn1IjX+F1muCjQmRH4wG61
a6aMDiDirqP6JjQ455ew4SuKEOnUPukf3NIWR60cTP/Ui13VQeNRF1uEHvDtl0zk
+XArYeMiEqEsuogMbveJCIvYmJczZuCEuTzE6EUam4PrQEQp9kfmF7jxaX7u6vdh
Jdy+7cmEFgyPD6m45cD2GAigh/QG9HucDznsyl09sr9C5KBnJ8N4NKrnyRAjlrLf
DPtHKEqzzgD9tsNni46Y1yt8t6Nr7xTvd19q+jXGD3EkzVQ4uBHHIPGpkptptiwX
CBsmFeRjtOXFddUVruTVgnFTEZfGYp+pVUp1h1CZReJpaPu08xNFUz1BFBl2Cl/W
xYhCVrKHA8gVzAfyR/TtHOKYoPw6GoBs7COUYG4w8W1RV/8i1Tzj5cpoqAwUTcWU
HAaY1xo74N6dWWAol6QT9WkVazrvJ8XSevE5owgW19PhQ0R7AvpjIr294B1kaDnY
I2eeLkNAhHv/sDFCvzV2RSf0nmEKG/cTjUIV5YHR2JfgjnKfMMTN/1DmQF8ie6Q9
1/2NRg+3uvixVynGYfPuTeqCLWjE2ISU1gtEWzQVQjmvf10OjQC62K8MzXtAf98o
Vvjup5fnPfaG0xLEHFTBXBWv7fjDY50uKwHd4vSfsn3TWN4LzADsYdedUqw3n9+5
KCErciZhMr03XzJE7zMzHpg1tn4yBBSs8aSqQRv3zFW8YLTBQFYwcX2mU+lpLtPr
tPTyZrtL/d2EW+aWcHw2vWVXAZ5Me02ZIU05hYNvcoA2oHw6TyaOmDGdgS72sM7T
dIpsxb84OQvG2KsRMpDFuoJHhn1uM9542J6RtkXPCpaq+Vx125Y4lnOLdsXsdD24
pGMnOrrFRYMq8eUbTqrxP7FEvaRdFOWpJOF+iCWQyuVpQIiPastPrQgucwe0zwj2
IEB2mvQsykFFU5qZonI39TihxuM8LaUvtyu2UQj7LMYK8pVhnWKfvJZe5ptyIQ0g
WkIxVDMjI/vkLDKov6MisyQU/cbLeliYSK97Vu7qEgs1xE+a66spGNbQqxcdG/qN
RxnR89GXuEFZXRw7E/XBet3iV7aSjZHCNBunZcU1N0ra3yHHAb5w5cpOnr35PErD
hpU7hTNmdJCog3x0V05xc5nF5qvZloLAjwtQU5NmgVZkYdru+0Pcweu6OHa6MwU5
tjQDhJYirg7t0BxCEkK2fu9uXqIIAlwFIfta+9pk/bOnl9PsC7CEtJlY03Nh9HNw
6mqVo3uQpXqyy5DOdKWU1B6P05OIT7Q6zib+olB+eULDhT6lYUVjiCdGWOuZHcuk
NN400vUjhebl4cMxFQ/Bc9JZ9lsGg2whbZqrxpeKPrelQUmZ2rxOBq9UtkRzZia1
BTSCjlifhJLqDtxBrU2VC7UV+YkUIyDbr2wFIe6kcwKAufT3j8dYJD+adFzFvIrk
ipu4O0CzD4xFL1UqyLY4M9KCi8STaLJzwhPUikmPrHCBZ0q5V/k+Xm3UbPm6wF/N
8d/pfFuZSlpj/ZO8wrxxgK3XxTYZf7ZLKwxpw4hIew4N4QUDSBpoVMpUhS3GAMgx
0JnRrJkpPP1UBnpnsqHWF2JWAbs0oY0aH8EHDU1TNkXGESUl67ZXR2iHDW6mSDt9
VoCL5ZPJTlsBZtXkqIP+9LIu//kC5Hr/NRNvWxYIw5roovSTcxIqvzaRhM2KWGUx
mfHXLljg+HJOkgw4xJ2AZmjs3Zw69cf72h+VYnz0nqJ9PEttrrgVW3+/esnG/Oyn
UmsfY8Xq+8Z5kabjZWO2a+3C9lUbVErhf+zkIr7dSIpwBWU02BoGxfFgX4vLKoXT
QcWBgTsxb4lbgQ9UdpCthINaz+BTHI31DFg4GVq91PpO4G2SiDUkw/1qt67370pw
QKCPDbeIhtEhvgB1CC3HUvuMQR8c53xDavXEIzOYfNwEERR3G2gTjwsRPqTIZab1
aVxj0oH5u0wc7FaRTmzU/EMGjC2+oTAh7STtzTOOtOrZbfMWQSEETtalO4ablU66
2Fh6z45UUQd01mjc0Q+K0BdPoC21CSPkWWJwIhIcfOBPL19HyLzKgzTMVShO+10Z
WnWadYBMJbTIOuztA/UmX33VxyB+A5ESz2R+WJzS3MO6pmBAkYQuYWACVNiQQ7fW
qPjHkTW2vo/48KonRx6YCjUtM88Ax4ii5eD0HrYcYXhhK4oNsH6BWLk72Ralm1Ah
7etjpGcGN9xzYkxGAEQqVFhzhKTf7KIkus7/IF9kKHmKvMkEb/wvAGAH4zwfsger
ZxPIA6M9qhADjzVculbtsukKiGB2KNrYGX3EsttdC3RlaQ/rzSqKuXgKGgLKeZyR
gZnXQm1xJNK9zKywvR31AMe7r+S98cK9YW7STd8nX4v5yRNimG3piuJyUgODvdmp
U1P4urPs3pkYM+NIsUdCCCD0sNl41PpCIy+Qwh2+Wqhz8eKBame2SuZgGQ+SZI6Z
J6Crmq1/4Y0pLtLMeEMtAQYk9bRFvEuSwLcMlJhRrpiZSOPsRJ3GpIcN+qYakrZW
JPh08krHznHnPnOJ+1WsuHtTb3Y/C8aRh7buCY+UXPidK9sfpbTkyoPcnkrComE5
VmOK/IbTz3a+8R+zkbWnX0AST3IyqHnkEtfCQRJkzR/er2qhdqNgP/EOFlEt8DRm
qH258F7FTEDxW1rs8F6mM5yRgblbC9qItNKbr1rajT7YQ8tYvxDXXCbG2X7uDmZ0
ay/qTHPi7ybJzExk50M6noeoxkmWgER5w6Kxp9lFUCg9/a+vnvfgif8fXCD0TbI+
on+88TKfqiwULSRX17zX+JYbhbYAyhGkBjP9N3gaWiNZvHp1fXlAUpV6OkdnqfCq
RK0nDvK0lmp0wypCJIkgk51YIBUVb7zZ/uTFoQhtFb+6LaCjirvO4GoQHre86qRk
i6DQUeC09h7tQLTCOuOrMIVY65ZqxZkqME1XGRQe1jpfdoPAdn3TMX9w+nYohftA
VfujpODRHDInyuddgW0XYhWbUr8yKA4jBKP3e2GMvoFcSoqlLLLgCPzUSJo6hC8u
Byw1kpjn1OhLRrwR4UQtbOQSsxFAUPV7gss05oj8+306lszqZlEVyqDkA6jzgrgI
7C8HdetRbAqWzPQWOJh44rNdaDmSLUGiPtiqb49zJsdToOfm7+nXJofvXslvaW0T
wPOmTM0FdNei0YiRPDn0ElZAkf6QrpAV+Z0WdNp2H07bysPvN5wnpeycNoH8iMMe
Y524dpHfajqX7UjiUyxIu+f5oVZg9wr6ij4/E0VjrxN8maZ73j5tqTarFw1Z/6or
hJW0oHfIUlvxBQSGrclN7DN0Vp3oKoSw8NLshd0+QL7q3LEruzA6+HafosbsKRJz
66xLltnNK80EshULx7wWaCaC8vaMTm3hjx2G+zA21RcMA4EFsfjvATSjqIVfpmk0
aCpYwI3hcgpqdboNcO1w8D7nAlciTeuJfkHCNxCmCt6UlmbDx7ef7JRF4PbUEjDw
0FQV9IsWYNAefyjELGQ9nAFGvuzPS8wATgstXWeBGGQxfQXI3fFOtRX3nLmmnDsD
mqteSTO9d/aZ6y13qaU4bcHlk9oXgcqgagev/rOcc8rbmACrNgf+9hF4e5UVqowJ
TtBndLaEoMSZWZd6mbWU1aO+YZdweq/g0vhO+fSNxA8aX8jl79ee5bOVRQB/3oFg
J/4zknxv8kEOBL6w0Lr0lHJLsWYxCnYtdisX3r6Rbl/4NFcYt0B24soNkwJRhxku
5XYm+1MdlMqi7+I5pPgLmlatKiyjjGyhntWhEJghLUBk+umibGeMWKZUhy/bjPQY
3YUMluPHGreEfbA1+WWmIqO3EIl3wjVARdkpGAYlzwB1P6X6y6Qgwq2uE2WypnCd
Q50w8fzXJp+tWXR3aU0N9G6v1/RXmEqLk3sLAcmBSbMWV892+JTLlHvjrPuhdFj4
g34L50NLkljtbj5IjSpLm6fMOv4rG7+pZi8Ryqn08SueFCeCuzzkKCGZ9jY7y0Y8
S5WHjKh0U0bxg2veQXxVtPwbvh/8fCWbordctNPrpUgGYhMUW/0zmgw72lQxeaze
oEGm/eXPLB7BV1jMAZpJT2AS3o+E+WifyAQKVPRFjPvOoEgd3fGNS/KSazmPi14a
f4FGPHTMwTjDp/U/j9h9250EG65m85e62IvHR0fEwkBdbL2TToxvxw/SJCj3L4Iw
3e4xF4T+TeROMcX8b/vTIZwoDvr/yvCOck+mpIoLWt4HeybHn05p+Y1xZQwvKK+2
742Mrzz6LRCOrC2Y3bgyVtSTQDHuvXPCZEBHXcHmZ/yMyyOTp1STwKqqK7O20rye
6NExyrWt5yBKf/ZGnUDTn/ShPuL2CdjPlJySw3J74rYTFCds5jSHtzJkXOsanQnj
FlJiX/ohYIUsfVky+L+7Wp2/utIU1j3hfA95A3IWg9q8bdOeawdg8XJh0UZaqKDm
K4xP37bv3scAbTl7apyUbcFx3UtmQ5nqzjTXcw9GYvAzcCYmlUwoiQu9d4sWnVXr
eGLxrgpk403OhXBjV4bpWwenmlg9uW8ggZAY1fDQVQnjtljEqlNUMvXrJHbIbkJ7
Ygxb/2pwOhA+6QHZN3AG9R45W24tnkOlCUTl4h1HNBryTusF5EAE634m8jsxu26m
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
N0N7PXiKHiW5Ha8FrZYaewUFWGA0DfQwPy1vGATioKhu8mp+nt7Os9+sty0mynrn
N8avGnx9CuOKNyR+Ugfol9bH0DNrK/8YwY870YjZ/CjEmzizhiSwdI4eb7CAkiW1
XsmlsIkeiENUTyOyLyNJc/acRS21ptS5msSacwBTWBWGqMXA7iFIYikflpPHl+uQ
NCqrHQP3DWSzfMgHRVzH8NUYQXNUnKQlWw0MlqPCyQADXBMKuwlTZqD7fAQml8W+
/xN4qi3sy4ioWQc+yqxZDwjZyhToe299noz9aWy0aUycXydEDHmL9qYnZtceutmm
lCqQF2zL0h0JEnU7Xf4q/Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7520 )
`pragma protect data_block
w/z2FTZmFALXxvUeDgxnlXUShSpg8rF7da9D5GEvC5SVHmTAmnpPhpqnlz0sTaKH
/xF9uHmzrtse9gs2wRlDK6UsA2M+2vccqNVQLETR9m1QNZZGvNILg95AZ2YdeGd0
8cW7fQctkvzaZDVR9Qe50lnyZckRv1QVq2ZT+eLwTkZRoCzpggdHlty6jBckMhLa
MkrpBhq2laCYp1dJBTVWNDpqxInOSXhW1Q6Mh5Zt9bzK7YXIwhAU88aGYwSIh6IB
I3LbtIAb6zm1U+XPGOEe7kPiIq2UsYgXoxpBctOQ37NdGfHviKZfheqicxOsyhRx
dbv2MTSrlYEf8VnZkO2XQDKOXMetHubOh76+xT70yWLlNCUTL/g6sotastAAngb9
qA4Vk8RLBgOKSZcA84+h0639+QcBFS61lFqTjETv3zh7hwF20UqZk762Ccy2HeNr
BB3S0CzEd01EUCytwPprUQJXclGVoNZxI09kKeesNpXiKxUbgMo9WOe2oR+4clCZ
56hjCBFrxATvYjIfcz/JGMvnwrOimAVqmzq2rGDfxWTknxDG6SIRXc5kz+rE7DY5
v2iPjEbJcIV3IRVullgVzkuQcXwDaWnlJGDwA7/fwFucuCOMkSUD9fQSzSKy1jCj
eq26kSTcjZcde5hLSpKJbDBnbxnlP1r9g0BSEkpeaznlk1deJXUBAgZXeU9nPmwf
gTZBpCieeEQU4tI6/yXnt+cIg2zXj8mj/qt0V3gSEnq5Z5YGgJD0DIcCZ7On04IX
yNibIKuVP2u/7YZGUqXPEvHNAmqGbpribdA3vbso19DAFQTGyiuzeiUfVhNc6s7u
QmmJyCDuHqGjbS87e6+S/YmAcwbZCuNzEWqnAVeUKnTDFNG1NwPbKyuDdXYKaFum
ausqJnGHONdvt205i5od8fFKQcyHDuJrLxEVfYJyqK7QfQaMb+v8ZZaP1CdoTgWA
UpI2Lhm58TTyqDSiz42x6rK/DfnSVJCiBYocP46pakj556oSsAVIP0avM+jxag/D
aiKlRYHSpH2SUHu1Gp4rRYEU0PJhKvJ5DkwjmtaxvatVK1la8H5sGN2Tk1u/BlnK
EqG0EnSIqy5l1/QQGb3V9n9rqdGv1Zq56L37I/Q3A7MptrdCEaNYtF6fFgoTg7Ub
P2miPJoWgs4oDNv9vir3jD9HqE5MLKqOqcVjrRwtwSw1Wo23tZkijd1zygv5NCcz
I14Bzmf6mVSYENm/7U8a+3Yu7Wt9v8nLibBj/5GOafJ04366ZjNexSB7twAj0xcI
2hg2J2wLDPlxboKTj7kesIt4qNoi05gpTF2oJm5xjeYQ306PWLNnhmX8sC+lGWsw
J6cgr4j54g7VNlRJ2HyOSvROfkdJV/8auPsVcClVLN0SYA/J4ZGE0Lu2BmskNC4D
kWg3ik8wYn8Mg7hcqid/hrec8wpVkrDPs7Nt1Ao/k1wStCqW3/y6+9c+sx9rYXGR
KfovoimusRGbxtEfkamVl595XuoUf253eNY8YqDT10p8rVWw1Y/LLkCMRUpZy8wE
YboLkrMVGV11nMEHdDGI52nxSADoGMkMSTVluHgGlb5JuA8Lf1VvnpHUs7hCCwp/
sMExLcvHDses1o+gWQ6YMjh3YZTOhZaLRVZ4mGGv79xRrrI2Mw0Ww3nve8lRxB3F
CZcPZ0vKbuQFIQL6CDloLLPytXZy5v5lBrzVxuuZjKFmv5KmvgFtx2I/SSR0ewT2
uoPhavfDje9W+gnLLqGOYdJSVHO5qP2Yq8BSjBBadiVBuimeZ0wRPHovBd3hleBX
IFH72Z8C6JCh23Fl73JfC7CnAqwM6x4ST4pzC9aiiluL45nKHg+YbT/uPBNT9AGC
kfGmI4hKiCTNaXlPU+ISIBufNa2SoUDx9dkU6WbwbzhN09ZfRL4Uy7UE0XqlXEAk
3Cr+Ru59pQqkbJYGutStH/H0Mzek1IeWGzWq6pc7/xT4na/BeTeclvQpDsc6c5Ra
VFZqOrrIUzGDQ/TgWlK8Zu7+mNEvqMY+k3DH9YefYL2BPfsE9SL7Nd92jZfboywR
j7l1FB21y7qonKfc94RWaaDE1/EBaZjC3OI3PyQ68IHOHf07wiVaWVzCTBgL/zqg
L3xr2RJLC+k1nlbCu5J6er+KjKhe0qSRkDH35dAB5uTTMblrwVEfoB6uxayhmWRZ
da5MzkRNLbY+ATthbvi+kvoGhpVZbJeL57O4iwGaTeZZHl90R591FzbDwEbWbhHd
k1bXEFpAYR8tn0i9tLZ0SwGZa2RgyKO6G2u6gnIMA7lPO5HoGLMtCvirwRdEchJl
WHF2TmeNpC4v5LKD1pOPhaNB88XPOaGEO2oUSKDygggIlbvVNh2Z0Hs7r9GQx2ED
tM/OzAmRDn7sSakwTapmYBmR1aFNBnHJJGudRCvkll3U13gF/KQHow2Q7Tvvz0vw
U9qVKXYfvmLWJEWQ8pFdZjcmd4e+tZk/QSPiofO3YPuHBNUEDqJmRLUNMRW0Iv9P
HIoWbvdALl3BsW1m81RcqwNd2SapYgyNJzzvjtsg69vN2H9AAeOCmpzVM1/ec6Cu
V3oTeKU+RCGG4yfmtVy7xuFdRO494AJ7I3C5VFq4s2E3OCHQG4cy+mJ5tkX3jaVo
tRm2WSz+U5+PZaJrI1yB2gLI7oXbkBi8SQ1zeznhhErnP86kJuRlC1ZkOnUdEukH
m9iT67n0fcrVKR6uugio5UQ41Sj7CfmYWFGf0qrY+BGAHi7BhpG8+zbyGeLfA7uZ
R2DqAlHbeavfcHs0VbZXz3s7KiL8Sr67TrUq/xkQhp55/rirZx0mPqrlEh++wTb/
2Dnwd38rhWYwXjUl/ja1o+TE8aHekk6H9w5poe0PrlMUz9FdR5Weo7JtVcdAt8nm
4zILnUfBQv4HV5pSCIxdpaA0D+bBq7DO2oM/j4DkR6YvXJvAVoNEWVp5xMRDv6FJ
rKx/jjXsHNLD1XqA5e69MHC4StNqPAUvg00eEWDWERnbAFoiJnQ6unaXKwn6TDIC
5IVOQS0B4rxmZCtCm+YUphSpmRskiPcP2D+mtbmPFSCCd/C47VkcV4iynZrv1WU4
n6IPGKxaHe0LKhaljaJBsQhE/R2eM0UXQxUfDv7C52f9LRLAd9XBMUbTWG2C06aL
pPTC39Q2xVlTJh7++RUlA9gB6uzIhZfbW70KGtbGTfs1efzIt/pFMRqYBabGnowD
nvrri/e22BjKyI0vYpmKKSb7I2pwKJprSJ3cthb2ReqULdDmCCk6PLJmbMB9MNxG
xYQrBx+eCW281uQgcHmqurPTOSNuf/iG9r4jpeH69H5SQTtTIi0tdWQu+NdZ+3s3
TQoU6d9zAo/ffv4aPKOug5V7oZA+pxf9JezbBpx048ujxzWchLzRqkdoBdhzSlfA
48vb3mImGQrIbUFwITtCNnoOol2iRLfZVIp7PFzEbweno1w7ROc3G+05ajFRA1Da
rehwuWv3ZIMjByN9RXv7NptOyp568pknJeIfs0tjS5yAHOIwffErUcGpaIrR+Lgo
N86pZARA2OmyzX2GfYPsjgR3Zp9OrI1IiOE0gCvr90KsN6wbBWBymPMDZM+iQg9o
TMGiioyldlrhWh3K+9wmQ9R5U6hZvwHOXSWSSErHhudnMdUkMuVel5GtfvvSwqoK
na8paiRiuThoxzHkjw0tIb4GotTnyKNpTqAQ+6M7bNxYvNJLujPnDjMsxtqoPq8S
yTLYkxoClEEHvWOmmjB1AO5PX+gMZZ2QgfsSBjD6aMJ4RL4FJeIa8erfgwbIntVL
VjynIL5Z1PXS2pLhO2fdNzsswN1jqNusm1D5Ij6CtUw8Bgj0u/uP99w9sGH7CIhj
OJy1CJNlYyzdLKkVyw7aVzoDqUXI/6Oslw/TrjkLSasHj0EYDtPg83FvirTZs1Hj
sk2v+sP7rngXsduJiV58zd6++I7dWHMlb/0JwsuK1feF9rjG+u7DFpXEEijuuphf
CiW6Yl1FF+0cTlNmLcgY06qWi1SHRUkI4vow4Pd4fOr3g/++c3z59EXyho2j+Vcc
XeHXirAP7aLBLlE48/pEVSVJHF9T12cnIAFcbFBwWNuhBIB2AMOaCK324ZoPwwZS
BDWvphqEMBrKvnVX6UFX/LJ31o1q8OzpJ2jOB+fyP7h3ZDPNmB/TpZx9ikajNijt
QfKT2OvlH/FiTWxOysUrR/0Fucyt7yq51kYjXJ0YdLuwY8cqz+8HZr0Tx4fXoVuV
dkILry7+eBKslevXiol5w5swsCJRTqxwIXOFP5tfJB6RgYgplqyh2F77P1Fm/REX
at/VdDYe8i2pqY0MNUnmedmfpLN/uLoOAfA8P9phIBPD5TcMxaZkdBObDvd30SO1
GlMLahSWphrtETbU3gFtmz3fvYn+rcl7gAJgSz766LdRpWxK4l5d8Ti+NnTqV2BM
8QeCyXp+9bpdHaoO1pLRcHmdFRGpjM/K+rRH0mTlWGIBvbrFkJJO96h6ZCrbf0BX
qa37/H62g6uShCmuhJYWWe2YkBaOW1Y3498qY+YJIEj6dOuz54MYqcM9yHF6CbeA
7LWRPey0cISlAcWd5gAz4gKdIZAEpkW3CUE+3QVV3S4qfPUwljgE0SmeWW6KTbd7
ykAAISyfdyNjgtFEUDX4ef663UFKVb2g6RmdsSM4VQEt3wx6b/2ErRFDyE043mUt
snmqVhb2FBRijF/NM6j+BdRDlokt2MVEmQ7kEeDcVNLLZBu3XbyXup6aXEKkGzkI
tp4Vlwn4hv/Bwe3M/oVFSD2BaILwJigGpgp4t2W9QzRQ/TMIKd8qetXGpwYtQNxk
dGlKSoPd0tIFPx1QRvMshZfwZl3OpTpBaG8AFRlnt2ERBWtCWF5BzJIdp/SaH5dq
DneEWZJJTcCwPt7vir4ogbD1TYJUjbaZItIUBgVWmosVS7oRypgOL+qs38RirbWa
afGPBIqCAUOsSFrSUxaUn9I+10JjOlR5uSCEhq/Zr9dZeXW/ohRF1jy0dpLmOhO6
g3B7gVqyOh4w0vFI6C6Y772ji2Pc0ymxFYViD9ETxHpHnJupHfBMI6VpNBbvvKgH
bvP7S+fbtn+AZgIfb0DlBjp7nNZUM+CfTW5ldgrtz2QLo1fjE4z63h37X++NnN1u
LsbwdmBxv0m4oXKf6uJkseOKDz/wKabyM3FIeWZAoPEZqHy7EDft3UCBxZzWGevg
J1eMUSV04Dq+crjt4pWLTzRh6CZwuTQy02ZZaXqyss+LuOyx1Rn7s7nKYuuFad9U
CyE+SGE3hcTRMgj/d1S3u9rMbx/IjpTan0A9nKr/SQTlc1XUwcmZulIRWZRvFgLS
T86dUQE5/8wAKc6II32nMkscT1pP4QDCJX5pv/J5F+QlyZOZSec+Nrx+tTWWsr3F
+SyJ7eHp1Z2LoCzecSEB6tzg00xkxyLomj2KGfm9T79ARa3qhLUL4JX6/hiNsHUq
rGUqb+kmN72ePhylalhDwtO0QpML/c0dZ5YGKchu8lQLoYLXg2GyNRbgaqlRPR9F
VxhKRk0QqejNNZJ0YeqO8OJ5VO9qj/FWc+Sq/zmy0rCs8fGaB6l1bQh9HNkYiqWu
X5y8NWFwhMox3tUac2uJ6y05gqXm3CTJD9fQPU+k0Jtak7MIpADTNevxhvl/Xnyl
5Cy3wawvU3alDyEKa8qHIXcAZnzaXMA4nwKxHPlbPjCkcd9SLFd+QAfdSzIb3X4j
f2VLJA5A4fXpDNijxrPp3Q5k2Z33BXmcqGAtjBEUcdQQAhTdzXXmsza19FpMPH9J
2msaZztVzKIKNf57vZbb0UuOZDgY8U67yGZ8PG+vnZ3ZPPQJ5IEUeyZ7mhvnBf+x
HZgOP3i1QOqCq7oJIS+ZdlN67wKSvZA9vYSbIab1+mnPBfMI4rNdiG+Bk7qxUnlb
fQOZ/YptNvFL/ohiJsbCpt1WFKhgjt1I6a0izrDHZ/LqpHrSob8dCxg44+JDi5k4
lnFW8GLSBpUPaMpApPFy882Kqa6DBdmZN4v6ylQ0Xq+0JVoykEmWunROovFVb/1L
VC/robAR1YyPiSJ9tdUA/ZcCXccX8kM2qysyzXSJTLmIEVyBP+Rq+YvqEJzeUY/9
NcYA0AhdaEJcKOoL6bh1M2td4sJ+gHsD5Tm1fUDkRoI0XBmB9+v9kD+U/imrO/R9
ZOU1aV+G+lVf6Ag/yTdFJTSoSvldvAFCAOMkeU0DoHFf4bJLHetNTqnwEtXLEpg3
8LwiycImpb9H9wGRr/iSoMplnyqtSiVlhJO/P+9TBQq2prR0u5W/QE4X/osbuqoA
wRF2sYUuywb4svM/E3ZqkX0t2bmHvV+xIC0uMCE+ubSkaCbzv+yOWa0WfIIkXs0H
n/JjvoYXjaIe86uSTCfpbQqJi3bvEjGypqCKBmeoHfSlIZauKH/9Kvbx4Z0ZMHV+
eFYdSlFZeHpwP887Hk4FHtuO1cJZtjmuByOJUfVAejC7wrtHUgU5LzUIFaSPCKxU
7DdfLvSU6k+I5xeZXQHCGwyuj6Pf5TEWopyl7WzThrCraE9Yi3NehQ8NjJOqVWKS
7RfwJFS9mmN4Pa4DtFdBkUwDgjQ//kb4btVwSxp1/oOZBnllesdM9OYp23/oKjHN
TR/WXL9Wa1bH8JSRHe7hmDIXM0/qjfKcprno4KoLidYtuud60gxFSCbs9uv6yuAT
N2850hWXYjU8ODytqhdb3gmoEiesKxUJDv8XY3Dx0mXRz4uoduMRifFwYiyx5gZb
vQIb8b6xP0TkSvCQ5CUhXEYlxAqScxb6IiFKkReQLQ3syYDT6/KNViijqazCh+lH
DJM0SdNXpqiDsQ35dsru5GXHFiitLccppx6gaekbw1HacFyMDapDp12Nf3SCkEDr
LOv5PrDAi6hLltzVRoDVg/RtyG4PwCH5E1nst7AK6FJ/dNSo/luG7UMp5vjgPhTU
IWRo2OjwI+/tKpMDgwu9+tWDOZ7srDkXEprNA9o7rTnYlIwK3szynDbR7fr7AOhA
fcW5kFpxOhcpKUprkN2avVLUtjuH1yUvl001AeQi5BPj5vgaeCnMG+tGOxx4QhS2
oPB5xQLGRQhSn7XfjlHbZA0QSeXYPRhUQ66UkfGQ1VQ5sn9hryfEQiC7T4yhdjNY
Df1y+h7oQg8D7dXvjAfws/L5fgKi8Uyf864BR6OqkYcDtJjqsQ+Kfq12tqNSmvGM
e/dyGnIYWeFa5x6uLpIcu9HOGlIpEw4K5ZNNy/bwIOEQbUHEOVLkSA7w2kFJV4cv
1fi30lDziZlZBcUb10rIyngbbcT/ZK0fHjy86QnBhjNQn4JgAbXR7kBcMjI8TwLd
aJ7JENlHe7UA2dqTHiLpXZhGW5WzQAIvfib9ue8++N/mYHc2evM0h6pjseUnsqzK
xs4opfwBRSa0tGj77U+pfvaH+gkvHic/ep+kBKbAimG9iOBWdjAQ7rcLB2dXLTQW
TSHMnfj+YnczFNnuTRb5atH32n6rlMRHA2iY2luDhFHFySK9k1kWnCwQ3CYtCvwF
gyzboqLI7rRINRqHxmt34UUMpbY2WuRNf1DzL+0uwG4zIbZ8imfPmaKh3SI2lmp3
/8Cm6mjBHSBqGk8NxfJmjmkBw0VZRz9nST+TSHWKP0udL5yRJmQMNlTRNtRuS5AD
Z8BqVmJjhPHRPHX0OheIPg1xaMY6S2Z+DXG6uIbpVKte18zg3yaOPQjWfILZcJBF
6mrOX5ZgfCP3ZXAhi9huWNOEN9x0yBkX86fPoX4zV3HUL4wGQRSxkmJEvxeqMZfK
uk4CHPSlBW56ovTmZqg8ujdtdRoInypq9xCHxg2PVza2uQflLrDKAVrZ14HLEs0H
D6IuWQr6YWj3J0K9IcpK338Y/rSNFx45dKSXGUd8Ku/P2FL12LhOhzqjx5351DMj
OYHPEKOs/Yn+BApzdMRrw3ZYgUtB0CCQG+PppGmTDYVvLs82qAmud1mFFQ1tzZgn
xT5M+Z37tzB5Vp9MOibhhnAiCTsQbqUGGB9jLw6WwpWfKIP1OMebFkjfHf4M+SzS
d/Lty6BOyd+1NWaGynNMmtl/Gdaa3wB5+d0UKXjhcBSL1MHNmEgvhcBe5kBlTTRb
DxAlUlQwo+AjAvduPSLf9Ha0hJLiEmOecqQ4NIEMIFXY7bs3MRDxIHrRX4TLUp0e
ECC4ww+sxsDia/EA0+brYC0UMj0dwkgxITYbiJGWHn9adjNaM2KGu1gcXGednEL5
OqrqdtX5gZiyDaVhWaHft1h0AmhBlL1bP3aufzHY2E/+GbixxBU+SI9C0/9ynupb
HYjnCEltRTHey2Ol1iD3F21iBJG35/xKnVgWjbkfUIWCknDBc3zOBtyBAoH1+Phq
3JEtJY0nAOl5rlgJcoSEZVMDSESfk7Q8co8IMmF21Tyo0ptkPYuNLqjmNbXGNC8D
gl8px54u6La/ZRmK/Da6rJAa7WtP+Q8u4KDgChoqsOh3mTt8BlQHuM6lNckqgRhr
BnOUqBnf/GosDrMZ5I8Aq6tF7sn1v6uFG0NV1VNG9lHfzuHSng3InOK4rfiYOjfA
H28AA0/chNiJbGqD2bAcioYU8TRJxQsRLldf7XQMfDGjSs9XrUlX4qdU8gdJRWmg
HjJKfv/wdS/Uho8ChmjDSVFJLtD9QWIHljZeDlK3owjcCbsFTyMkJ5a2JxSOmgz1
be07HcbG9qLR5aooBE1g5/fiJGMt1SIexa+qYHvj7N7grXnEI+mAZfOuFJO374pd
piUWDegdWNpNI01BPmAHvB/CnvDqWTCCYcW1etloPo+dyeJTA1/uJJG0S4vBI7Nh
XVMSzsqdQbmfGUK/RoZr82ZlG9EmNDm8qLn8ucAjvKg739BQm/Yld59wX1wAwpmJ
idlsbIRObQlsrPqHLhGgZ7mO88m7ff0V/k9OVaKy9uisZRas+GvFfS+G+nkbuLrJ
cJ3ST+jVzx0MmELSjznlxp0Z1CUZQKmfYucOtIYv0iPbSxcQpnU7VtXr4EZFwZ30
99FODWXHciFfygFYILJBZA9V00t1WpLT3hpVvhKKZPQw9/oVfTwdkroQ9wmvbbyp
N2iyOoBToy6aigGnm4eyjlWLYxHdwGgWYfnSlkF0zlixe0pL8Y7+H/y8p6l9Dhf1
O2CA10vb+O1JBbtBJOpd7P8UGQGqqmmouovIRVwGAJ2vp2CX2HmJ4YjhHo2Y5MrR
ACZMFDZZ07jbRWCRa74vliVIewthA1/a7FmKWwquMutG8rg1DMzuI4Ue6aWtX5LU
Sc1SF3x8EhUoqqCu0cSP2qrzdyxBbSqVpk4f+vKH0/eLalMUS2CuWX+dG7LXL2G3
CvEtAIbmCqI/FEgAOR9Bf2k0R1BHmGvKxdJbER0Rj/zhFWy0QOfoMqw/JWsxmTSn
wjxw2xOQC4/DNTdoTZnp2+KOr8KrC82zcXa/4Df5xL5NE58mLWnH3ps7hlTWn3s0
6va8tTK01curJmhdWYVRGbD0Bjm5TH2EIta2wt1COBLOA9mIkeYIEs3fCATGDpPc
LBfVoKDV/OmGe2m5im5MLMUdJyZUngImxbM+aPjxFliOvQq41UOn/KdIoW4Iu0NS
LdzJhNDfYyCaeikRJTgwEUlEN5+Yx3IbZUuJOueW6tNkJwQqDt2arCghFT4M8odd
QNDptSLsQjRav50y1hAhnt7Nw+hKNcUZRK/X9CCebVMF9OhiqdxDBUft96sKwsIY
NYu/c/C22Dp/vRaBme7SOtHN2mTxcE8kWMqOb0XTA2I2ebqyf5MHDeKX59bexl6S
mnF7KtjNIvg4qPIeG7cRcYqZ2hdGc0im9yPuMKUzHnS8ArT1W0w+3C+WmMG73xjt
bFI9mWhrxthus6N/B0Vb/bXFahE9wd1Zxrln9lwRjUZejuYBsualc5+CJ+H+NLl9
G9gsY0IT5l9fllhskKFKmSUx4ezD3FK0I0iJf620JMZ6YLknGQY+4rXnrDpDM5b2
VHfmtMH4NDN98GHwnFl7CJ1p0finb/Rq8zmm+14ONSSFbuP6ar2snJ5AjmDMFPuT
sXBKAmxbeMw4nPxAOY60IP0Ugxhr1q2tLqRKeys1AB8=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jyAzdg3fssBFG/qwpKHHORo2U6QIZFZ8UrhKgx02N6sfk//CI3+ZP9fECNcH+oMV
UzgaZm3k8qbDqHjrdaqAgdrThWGFM4xBHBeBU3bGo1t1LKVEtFcVDqPCtdRCXqgW
UOm2l80pslfhJCtpEbpr59RIV1IkDqYSEcycL+LQG5sKOF7e9/ikMLoWsa8a283V
oWGlPgVGIW+V4YDQpBwPomAvAkl920NgymqSo9CkoL6GSI2F4ot8xVh9J7tF2ANu
4fBieKx9rnZ+jm2VYuVdxSEbMAJOcVve1BUPcwKlYsGsVjd9X4zUFzrya36KLat3
/dkUyR9FqqMcFYMFvL9adw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4192 )
`pragma protect data_block
t/dmxMrNiHRtfK0RfR6G4YLQI2fHZETTH/AWrFZL8y97/+pcguL0d3qTJRGwSMgM
AR9X61IUwlWu75nfwehUKW/obdENrUN8W8gGYaTkWgAGXb9/usJwJNSogI8/WJpW
Zv6CIMvtq+IlXi84JQvIsrNLBT9mEKJ/GCITjDlylogjO6WeHGKD08GsR+N6HZIy
k0iW0QWg3P+IwQqcsmxn5iknjiyRLtujkyz1uwPdwBhfjJ3AbYGVbof+qTam7ybx
HvV/5P5Fv6jeFKHWxUjO+8k2WrpD9uj/deFMeoNoVSjqF25Za3GCojZl7WGW7HwN
M7ifOBAfhEip4XkEarg0m0SzCb/krRO74yFW2bHS4QNk0T8XVS5cRJ0cY6caFRph
Mx2Ut6w2uRq4fEafKGFueYpd9aJLjECTh1POrtNNZr0hP/uzuCIttgm1kkAIcIne
NAW48Qw8jckinl+uYYKDhQp4GvkfqpElYhsxLlr6IsurRx16mXUkrqHYHFDwPKCr
Ygucv9JnUZzGG5uLinOlL9D+3zGCQ0hD2fo4QU2DyhIwqZKs4wK+m4mkMkGgqTwi
Y2BGfEt4KlWsQhhr6Wi7l3J8MunORp6jyAo2pWxPXUK43TF8BT+lNMLOj11ptCE6
uBlDvMKwD/5RuiWqGAyZu2F8+Y7Coqa4hje9SzudV2rzk3PgmmYrOsbFCQwDx8eo
5PCr1e2yzgKGI78KO2eHTe7Z6jOGoMGoUhiPTNPAy6j5F7G6bZPQ22IXL5OC1BOD
W1yYDF76ajfY37PhEukakBN+6WADtaa3T8DNxuBN1o2wlNIxVDv+vUSmjvqq99mu
/HNFthAJyp4IYwaIuX6mjcAIj34Q0b61Ge3SX7LPFZ7c3VUnpa1fmJb4PhXBrRhs
6O2xGTXma2cGmmRQmZXthlmmqOaLsvmGqANqCeRysD5XYg35unDhe8hc8PqpkF4x
TW1sPhsb7dz4YSy33BunSjw75a4Cf4+WouMhNFEpSJ/0PUQzHKai/Br6RF5EAII4
pYsn3esm/9cEn/k9Ful/r4SNlPgpgnp5zqnHmYdW/B8prVetc8gkrp7iSf+2Sl+b
+Kvj2fQsqouI2FQ7ER3WgIOdbBUtKqPvxBZt4f1Xun4z8ea0P6Q9gMzn9PzkWfXZ
MnUkZkVIFPNgjEXw2jvLCk64xTSVk09cVu+eeu99e/r+2XHyuU1xCegnXLkUrVKq
wlDgcK34J9PlZvSuXub+LlZCqGKWhhYN8ORqGbF/nAFEjl7vbhv6En9BH5cGrLO0
I5FnBNuhnHVGAhyrPHW7RocXrvbhckrpyMFLFEJ7QFMjHwM6njYN3fsdJBkKX1v+
A6dWQypI8xJyGoDgEecC9Bdvd9B1H/wzmGux4G/p624bSSeUKh0fpgmSkbL3jwLw
Mv+fgglYSk6YEgwrssUKs7prXcW6lRob+odUOfQ6FfzH//c8/juSMbpHtHvJDTzJ
NQ/aI+BKVycocKBqs5R+ZtsMyODJURXl18n08uqegfKSC9UwpP+2AF/sT1tPiK4K
Djkl9rXwxqsX2p1SYqVNV+nVesCkb796q/VBQqM++Ao+Qqjj5RNYrxhIA0Vn77CL
u0zZt5xOC3SCV7HkwrtMq+59NIf19CrfWfUSRnkJbxfOx83YjzHWNRVkWqAs/xRP
DWWr91w1D/e4hEBf31zeLP04ElyJimVlrjdrNNfm1OEjVW2KVTNI2YSHl/OUd8tm
RHrI51a/4d9mVB9h/O587q/uSlDOfNxoWlOqG0cvMZz5Xiq5Vrncm4GtGHb/jnFO
xH/ttTyqAlFiKfZ0dd8x54Gbtj4jPhSq5QAh4/S/B0ZOIj0rMLx8ySl98Ha8I+Ij
Q05fHmWvU+PZ3rxkCd5YsTs3+93daHQFSnBJs+tRpuoAXw+5EGpygUc+CrL22JVu
7Sf1yaP3UP+tnH0MVoRQeNqsGMb+1w3Frsh49XjCp2RdjziL+hSuwdYmpJ+djT29
acT+eyg1hnXVD44k98NaFxmQQ6dOv+YtIZ6adNma5bdBBvcwKW4Uov0jNpPw6XUd
ky7uWFUhr+l1iv+ZBUs4HtyDfMhaDs1Jb+xhs8Nh+hTTTYNfF706Ll45Fv8pF6HB
t/K0mPqZ5ZBCr5ZldE8iBXSsfNV0cStBnPOU13bHEE7jxYqzFtYaoG01NzO8Nrzp
nENsKa3y/G5HKXS1hYHya5CSSo8ERIUXcgTpJ0S5xpT/wIeHPRanSAy/JlNp1g2k
LSql7w2mANojkxDjYUwyl5OUcCtOPzfe/aPpU2QvO2NZ94s3NFt51OOTDrdJXExT
+Ck2sRPXpzfyvZw97qNsf/0wfAFG/vsTUAAuI3c+IgDi+IE0+lJeZHdVzuUHdiQu
o6ewsd6pg/Vg4wjc5g+XTmAhkfTjXDaNRJsJm7wWbOd72kD6YIe4c9PYGXstzLS0
aoTkeeUI6Qp/88wwqYYvHp/riY5w0r7NLLQBHXC6C3KDLiRo1A5ccCw4Mf2APEL6
Ri7D38iAbOk6M9Gh58ypKCSCdDBxa4ZcWYi+5696cUjVosQOf5yYoZrTNkleRrSu
yinA0Ta6sh5BHVjQS2dwK1kCFo4PM8VLGWBpostFhiWdhKlV0eyuGZ1KqWqvAipR
cZVypTJt7YtYQBZ5lW/QMFgrXmG7Atk+Lj7AKv2FU2Q4wJsAcVc2pasR6Av8aiGw
VyQc+/w5CrzA+Ezj3jO+bVLFOWNMAPscUcaTEHUxLXyVIEbQZaqKJUh0c7t+BU65
2doUcuTb+CuviKRIR45wUxMcmXs6EMFQb3hDgpT4dFP6OSRlxB+JQc98P8FDnCzH
t+eFc7KkNVcvPPBvfoP8n4yvArQ7iVY6CBjUNmcI+Q7QUQpNE1T7rDHKBrmnRpWM
IwY3GiugwjwIAPmcY7xjo1KvtV63l7zgQkSK/lG+RtVW+BfCbJvf5tIBlLBYa/2F
4041MAsvU9W3Abns1a8Tm6gepn83PhzMVgsLjdMDFV5mDMYTkYY94AI+0xnb6Hv9
R3gFeKsIaJqgflKCopooyzN1H4v/lStWG1Cwyo2O+prrkncYuKUH2eT9Kh4NnHHG
mlrfZ9D7PIV29JFseh7ZRV21hl8glkAM3wnEdqn5Yur+azdvGDCGh6cgh5rQOjTq
43WyoUSS87BdyhjF0PRTI+3AZYio/8zTMLdDtTQWecj2pmJ2v9/HN6HuHzvDoMDm
2waxpksZrd6jX0zz5LPKU4FdKEQgl8IjbJma6LXFy1A7XEzgT8c53lMvuZPYzsIJ
eCQcNzDott8CSsH+kWTZbSzJ7lj+wM5aRR7nYEugdbKIT9W0tpSy0iMlwnldAxab
hZWS6G92DYNsrthCjKJDLBoI+yod/R8NElfGW+rgCeu8pk0F/WLhRoLatHgLG5KY
qlEH5iK+xOxIpnvZ6U8mgpJQaIQmDlAt+wM5X5HzH0eTLs4TKy8lTmqVokja4uAf
yvu/reYqpzeNyoAJRVwkAfaCOHniVJyB/6R24fKt0QaZ44Wi93nZKAmEqk2rFRGj
cjy9xWVWBKh4NEsu98ryNUzmUV1V51wkt0OEeYZY4v78oEE/SvePvcC2ZLq3C64M
GDk/L9/tqS/Shz/qSuRMxBdcYVGwyzEAsSon/GWd1Luj0weSIT0imPGS93EjX02f
uptysKWdvm1+nD2QVVwPi4/ZLAh8ywfHJap3H34C/PZqGs8v/WVfScsIE1zAfjyD
Sjhq/C8ScgXX2cuPTSzIXtxCFWArcdbeRhCNj7zd4ZWVjOMBQ4xklLEAwv6EN70a
P21lWhmw66tThFs8dmFv8He0bHZDD/RnDlPLEJLB0DA8BAgZVNiVLcl2qlLvXidx
Hmf7WXYoo7uOjlwLbAUfy3MQ8vkKhkncNSXTDmgMFKOXLuR0inEG3MwKmBBV2aKM
5zQ79Jfov0OPGQvheUj7qe39+NhM8XVPxlDN2Vo+14qbaZ+Q2hR0XYoWmDM6Kpbb
ZTZ/M7PHZquxonZBC7Is+UbdTk1omAxuVeqsNY9TGewiboU2PvvJHdf92n6G48Po
R9389FSxiU0gi9z7RLt7Ix55y5E4E1qmaT5cCGXKnC5sahtgFGPefDmFGaLb1LHK
s06p4pyK9MTn/1tK7CjSOU9LB9eEGFHqGUx3m5ggWUP3pAfuHlzMgOC8V0q8UhPX
3ethl5rne4vY56A7ehCBOip5xeAAsKYOV3Gr6ExuqLixDpfd6NQZKDDeLu0bm0sM
9QmoTsdlRTR9vQxvIB2FDaawPa9hJRpkc9Y8SxCMLEeaUwBnIDTPA5YW1angoJEd
u/IRsFXhD29KRcCoJoeH9aEZenJOmx7G+kbQ8BHLwaW4PjToR9hqcTCkF0O5yK7S
CBNDxBBGE02Zs/A4Kun1BnR/c6QFhzmk7LPh3wxyWoQYeHLpvm0QeHAmmaAYhcyY
9n/5HZxMSXV60SmTN7awTZ0ndQyG8Mbtz8Ckg+a0YDlc2ziqpyOR3GgNg7vVQKny
DcTMRQETLNHbihzak0kf8Xqf4zc8zQ+DEepVNfJNXSubPk6gFUcF/twcsl4iVBZd
7FA30/j5OGIw1IK6Xn/OfxN6r+2fqYPyFZus3KmWsWs2r2gwQOecrhamWeIGiEmr
MZY7VgugDtdwvQkmrjfDnXQWzUkiX81jbEvFAtczNOTZHgWmRBEVOEWLdmIC4XFb
g1GQDouwcLDIw/kK0d2QPiHCGf4eK89bbZCXZJQ7uMA0W0cZaY7tt1eoFbStfogY
awLI1cgAK+AlEwNt2qPBM/68L7gFMYJiPmb5pF95Q2r5LJKH8QaP7+hdsLXkJC2q
/Q2lhZIIuqQFgZH1a7SJgtq6M+XZOw4rIFA3nkymIYCE7kIy0/2eyDd0kXOkogDj
Wbu85r5nR4Pz07NRRSeOPxlf/eBjoW6VduFbQtocJVJE1X9OZG6oMXKG3vuNzgxJ
5Cr1tsr25152kfMD3v1KtPYHB7uyEc3w5jWBpHxuVdk4kjIyBS1xnMfeoCUcR6io
3+oXk/yUnm5y366FAnJkv5pFNeaGcn1Q/Vl/sn9LGDfEE2uZhy+0tR/BHTHTgMp6
At6gHTTaLnJNCrly7J9+Tk5NWCcnHVcjbPU/1g8GPIM4r+wMdy5KnttARl/IMm9B
4nstboy/QRhgleIX3rueDHnns8+5k90h0nUrgQIBWLufKi9CHDW8XEHAhRO53kAk
iSyx1Ke3T0/LR0LapC2vEPBVCDdjIdYEoni/5cEmkyKmHsfM1m5UnSjkyWyfDbDC
hMPEVczQvG7ipov5KMiq5DrLCUXmhOklq5pMWDQjgyEXa1vzBP/bWv3ZeCos8w5J
shwtpK4nZCcfyaJiNKQ1shRR3Os+3Bwf4ADsXEUwpDcR+KdD+ycRvzQHNf4Z2fzs
P6j2qWr1KKJ/loaRUF6QJbel3wxdENySomlvYU/h0xqSnkgwjlOe5zIJu1L1N59j
7BTI+qU+2/vuIGFFqYCrVpmPt6jmJhAxkRVXWs/aXKynYl26zlD+EOpo0Ok2U6tv
J+O2LwHT7iAex2B98BNmU8aZ9VQvpSoBXCAMiO8CaESnFFWTqMX5te0HMEGate+G
IoPh9v2lcWg2zB+ipdEBtw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jmslWujGP5eBcLhn6MVkNRJoXjCk1G8PJnOzASA+SxMHAZiJOj2uHMXziDtTjalr
7fn+tVSE3EJfuTGnjjHuKrmc09JTZyv2Grb3aaqExvKgCzwBDnXZi/OvvJV7EkWR
n+e3SW4T66alNB50PAnhQHP/pqd/3jAa+Mok0MA1Hi1DZfjUrm+dwp4E0Ssf2w+f
vxdNyIgyFTWNGfKhfakO6rL6tWTccu4NZNqmRfWgu/jV5/ksU95wlHlMnGa6Wg28
N0sj4CWuPhPDJF/wyE9AM3EAf1RxR/aPhzt/8Gv0GnOilvCdRban7T/ztS/qSowX
J9VWJinEK9GJjAhhQaTm2A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
OsDV2tQAEWkPJC5s/5vMmDwbmOF6QsbeAyswcq12Ve41uBLlTVamGHzk4kXLdEAJ
ZPFiweFQOaifHWTkbllQBzevxuMshknH7aldBHgZFqbX6zuHXIt+mctiPb1vRppG
XFaV5rS37SJtGqxvTm0EbSd9xy1oSYriQRvwolV46XsSfUuehatifan4qYbsIaBr
dejoFW0cG3+gvDiw6qPIGwcFd1tfmEmAnsqHa6/nDz9EdE4umeDP32KUZ+090TtX
bM3BOTOSvWb9ArnhE38xTjLTkxqISrPgF+l1oHWw0ATolVlxbheJdPRPrf2Cno24
+yHseseHdkcH65Cm6UM7xEDrjlfmVQXxnYZY0hGW7bym7Qm/hoBJ5+xUICucuU1t
YNtSXgXq3HdgefXjVox3bHg82uKutjKg6jzkiA/iGHpE9Us2brqbQRib2KxSpK2t
zDhKmFTDiPaYe/+Cw5wLXIiLTwhmBj8SBoMUmlmKLitYOPcEivODICdWoQGkyarN
8fP64vVDij7stv/yBpdlJ07yGyBo/EhnND5yZtoAs+L49MofvYUDHo6nAr/s8Hbu
+Tie7A/Aom5RVzKb3QznLFyhR8tw9LWSj65/FQ6Iw7B2EtqzJvXPbCe4BNazS5CU
q6p/ASvQPqPx+HL7KI3Q0vVwP1DOW6HD+XfYtsYeWXe6skTHPhFAXyoQLZcKOb5i
b0wIqI4yEC4JG9FrspMd5tSzw7eL81AKl0YPXRcTMO4hJOoVyS7tTe2u6xTUX3cZ
yYBSPBOp9wzMJD3W9LSxP3vWEGCHiT3/6P+n2ir6XMmwrxy+lzJ1FjaZX+lQgM29
HqG3sEAMRoR0LMKNkrvCZ7BIRZiG4OvSndgiE0Stb5eCag/Q1qA6cpIPFLMA9ekZ
QuKOIMcVJpanOuIl9croY2My1fWOssNdSvq5ihEHhEfq6pHI7N4fOvwO+zxHMtrR
k005UDqcijMfnjiVBF0oAXTshaj2QIMwjJ1wywNu2S4l1Kx7MU1TYdBRFHCD204I
kdRAbR0gmENoBaIrtZFLg+tGMnCj/1BrXJgHKSt8uA4cKAa3SKu3Gan1C9e+k9dz
CtYL/ESyvjrrjquB+BmH88bUMhGz2C4WGN2+mhrwidMcVJaeX40LtIkg5D9v2iG+
MkVCa7pdI3WdvesNUfjldZefvIFgQk5ffYrlcRQWr0kvz+iVaDVsPALqhPCs7Apz
03Wv2yBsU3K7aDY/MX3/ZlL3LTMgsIRPu1fHJEouEQLudYzIQAQpiChaqlfxVmH3
IunJ4eJW0+EIvH55lmfINOqA4GsQELl2iOlHfg/GOntZSVxp2e/Ed199bRh3lUrp
jY1BgEhyYbQRl06z4IUutA8uiH5Ni0NIpnPYGuIGOiq2B7lt5H4qLMtfitTWLgxJ
P1MqXMfbCdMBO6fiSR0RWzAf6gLnfWHrc0tZFa0fWmt5UVUPJXLCt+gN0PO2uDC7
uMgdjxYWe/OZoTH26mxLKALQXn8ZRi79MK2eSxx0QGgH5+Emj9rujtOLTgQllfwN
PGGwgRK3EJuy4qZByhmxUReN1iwdI3cNhUwgazC8Y8znKmkKeNasyzUA47lGNkFH
FeB5m3skQREEfXORwfjtL5ELCS63kzSH9JamLbfbsyZVHE+LFx+zBsiiQo5YxlAm
0pe+OWUCI8j3Z0SopmloDBGUv/wTwN9nOBeq+gqu1m0A+zAcMF5Vpmd1NnulMwOr
yabrU0gtFUmVFxIabHxIgRW/dZnJm7rYywNBS0O4qTAoN2qsd1ph4S1/gFzG7UPK
12WoNz2JO0X/mRFSAi/TAYmKep8vOfh7UFrMgYmf8vNLRat1XhCQKKSkE2CGXnCv
qD/NX0Wdxk96CA5ds2JlhBpBhlzvSQ50nMG0hLnE68Zy4vbo6kIlfPIo1kpn/5+T
6S/GnQYnarfHNQne1rkNGe/Ix/ll6T67m7t52wRTgTtskNkuw4g1nNA92Ksyagil
1q5t8lM6gFuPksZchym1U74ooWhFxTfuoQJWHxW6+9BBKG8tF5rSBDHYTgQyZxzI
SM1wBL28YBTqnqu0fJpHES3pfBTpXw7Okwh9HExMs+ZlJPM735oOsQazz8r3308A
5eD4Wj3a61pAM8EeG+xgYitA/z03UpKAGkqxEO+z8DXpINXJ5IWPxv/g61vQ1l7b
zmHU4cnAiZsCqyrfueWnzCHrUpX1Zt4W6LERBLWcyPMpEf0p/L1hCeU3fzvdrOOj
COBBI434Uv08DBRI52jsz36/0x0EA0C27WvJSfKchNx1KbmhPh/lqzSd3CABxoxC
7qyge4B0uaX+I9hg21k0GnVuY96VPt+N0eX2CNJs43EMskSOJOI4xCDFpI7+htY0
PWQL/27mIJjA05qCHbusPO6xa4in1Ku0W9o+UW+bYGkM5Mw/oqJgYx6NXHFopcAk
Nyg4Slc4eRgCQM4Xuq7MUeODF9RI+kbhplh+Bdc0Gqo/xhk6mHDLRt1MBP67vXYW
I/80LHRBjZB5HGWWd6d0kuyddlyKIYRdosHvrJN4n2T0fOPzt/aRiaPu9X+M3kVu
x6k2HKjcTC2Mmz0U8zwtBT/T2K4oxOPWHpDUq8bDt81WBqyt8YIiIysWfX22BfaF
buexbc8YDMUTjVo7OLQdJ7DRum6tHb7/VDTizhc2LHLFvAzbiROsn/lbhxkSS0B6
L+K6v6I244u4XCb894RO32cMiggOp5PNptdE1cNUNadDd8ppi40z5czIsR99/1uT
Xs/3XrkMGPL0ZnrD8i6jAWx2uRtvK4+2zcyXKfYUdWeZ/7v02RIK5xP8lpJsW9Dx
MkYJZeCpkMYNQrdb+rq7snHR8iSGB4OSFZFYcJlk1Cr0hnsZX6LftpH8r+jy5Jty
DJ8Yh+l5hvKfwdd3QiyO4AJCvNmhCAXeVFiIjhdyOP/R2ohjxXGtdqtGmsuNKSet
IejApQLO+M7xLR89Vx3om4vIkbmJ0hWkzl8777yarSl38KqD2fYi8H0LjenQFkae
T0Z1wjXjaIVQk6MZ0LgHY38+kN5ya6FHqs/m0Jzto2vBjA1JVRXgx4v1OfYnFPnl
5D7B1gD1cE++r7VD5kQHcOFlPSV77oYWfYidDxs8XMLWasDBrhY9bqKYk0vbK6bG
mAA8A4p4wTzZVd6o+62FfoOFTyS/fMGeD12qcby6Rt4jeNSxuGkSk/LWOqor9Owj
n6OZIqbM3iGrqQoD65NEXSoc0zl0QZj2e7LHFHgew+FYwDgMj/nL/avAsmQHMLPD
xMMlTL7kYCTu/BZNYyizEVdPAyMoHSAwBPBzgmScV5YcxWVLYVGWOHHaVzpwGCc7
tMJMbKK5EqFSprzS49wifPCg5lZIg/bJ7AHdrDmWd07Yc/Z+Zta2NCMjrH+3gMTR
vBzPezXh50UAmT+jdGuk/4lyZg6Zc6RxtUiXJ1N8KFical0fiq2VVodBlPNwXFvo
RLpTXYrnoAuE0Dwb/0vkD+XF6YKj9dC7UJdTjIK7Owgxl669ek95StFLAcP+K1pH
BesWUD4iWraFDxDWqQ8ApraVAeX22t5ZQVIsQXac25MO4xJp8k8n2ZLnCdJ7xPQQ
UGx+l5b8qJWwa2a5/5DzxawJ+Ng1qwj/4cOAjaFhoqt2evDcQvCZ/Y46kL5t0lO/
nkOmmQEqWnDuqlHpc8x0Fpd/ZQ7qtRPcUabUev/XhGJfqUFklwQ4a+octs/n3hq1
3yPQMMsGl5QIU/WN+bM2mNOY9OJ97zoDTaYqU1oHABMzu5o+VXcRC0iKnFJYGcA8
DnQ0Rc8Px3nMzBhFhMjobwN7HoiuDi3ayob4ilfYJ8k8MOIV+7mepVgXEbhu+oKc
lUdjYPTRA9VGKBW3wGO8vhQKogbnqrPx9dekr8hajPnECNGkWo+tS9xNWI1oLPJY
ui8Tnr8yfwYJUfBwRWmZYm03xps4nWqdBrtCtfbp9Ue93xBnF1alVdr+RowYhIIU
06TpyvJAcghdltw3ty1l2Wnaha8Azywjc4tF/fjurrTSVS7mNndFaGOFJtH413ds
krWGs35IzLPyDAH/S2r+PPod2/W9GBJuYHB5gxlYJPz/dPMelwDyVUWyaPOoYQqN
ZwgTfAjEVudCgv2rhLoXZw89kmvGjc//vsM3Q8wbde1NxFU+YLbDimddX+H1ItWe
6SuOq9arHZKMZQivIowPTBi7eoBKAYO79NORPhtfUaNsqKqwlIMpX0bnxWYpzLQW
did6tFQ91edSG8QSQBKmuJMyrKRgKvitR34lsFdjY5A/JP4l7S1mewXwBUJygYCq
f5oMuFJfP9wZmrSWNdDCGHZv1gCwtIb77IH6F78digHO2dp44UToKHT0mX6iLRrP
+0p92lH6FIvU5eA/HoEHGFwdtqUKQpOYlN+WpaCUuqnFpIOdb90y6xY7Q/oM9OHn
+BXP3upps/qdkIPJAudnDt2DMiNjF+DQh+Ax0PIgDOIhtfsbGuB6eG8Ru6SjI0H6
g1sg0GdJhpHwRLMOvZfAsNCOoa1YcXCd/3vx+iXuwXzGHnB1XOziP34kfCFdzIij
1J4/F1pXBXdP/gn4JDX1XN9gQDFJciiWv6uFJb7m7SFiDrz/iPWoKPcLBJapqdlu
ISauw6ZLwzn7grLS+o8wzVQZSxii80Jk7aKeSd4tb7yIKsEWKTsw7yce1YwMffL5
nB3DWSv39nFEjSpfqGQ+18UnYM4PG+gnAIrDh+DeB/FXhSGIIA0CmwSjvg/o8SSr
28T9Qy5VhblUVzsHWJF/mM+WFzSrSW3hDCnDCSlfNywI8IREdgwuS6TkN1bh+EV1
uX06Dg8ZZsexKWjEYW08QjWNV3E6X2sJY8sZJGha/eyb8aCA67Y/hqhIBvt9naMG
au70yJ7edsz5zbvvYdZhGcn+ZeC4agwG8WkJmu8mNU2XtVlISCFdo6q8AZUUwP7r
sr5tJZfktAiQXXu3/VNF+xB91HUsMJJyf6S2nCtSueb1jAZNi3RJzoZzKATt1gFG
xcy0Ut1/f4iS1UV0ehJPuVGRihB2fTbp1H+HBgrFidVvTf6LF754VRuunRsDwsab
DFWeuLlA8FUp8nVyOCcfEsQbKjIIsSZdXqX1DpLdfSBWRJFEEys/qj4ohkIPLUQj
iePibsHEl/2clW2WlQlvXhuhhA/B5ySyMl3/BQfCJvZN4s1joFxAEJiX37ObR/SX
YlOqMNnH/x+DXYa8w0Kaztx1KznPxNu9txNf8IdgR4prBKuuH8I4q1E5vtwHIaTr
DLWMwzYk/cluFdYWgsTELfJoW7mnPpyyl+pVkLIYjmt/r+actoZ4QnOKKqjDcH0t
NfHmon36xTEtpkd5MKAkPOGGxjyXK62nkGIdFQq3dTERMegQgMjRUo+c8qdSJP1g
zRjXGizNUnsc7lPtEfr4zuGOY08dYf12w2eR+er1WREHFX3Epl6rEaellPPDnO2D
0YMXR8QgB3FzCuHaTcPRByonzMtPtFn8Vuotalst3IexHtYypLz1a772JIA2Sldg
uw2pVTobRa5WH0peH7G6M/XfnYorjjsucFjEbrhZcb9VKTSeUt8JMFc5nrBhTj2B
GX7rfjlNkodOK+0LEJUANrqTAJ1diOCyTvWsR7gXE1yKJ5ACVi/r7wuePmpO8Dxb
OJWye5oaLr86f4nJ1qajUwiA0T7uIZm+AQkEN2ASqI0B9JGOkf1oI6LEVw3robH1
r8NBSY33ZR2dbv8RCmshhKOSbbL1+EkhCdnK21H4DBGPARqBZLwf0dAmpwf0P3Ic
OIsbzekvf5n8JE9AVaH+LgnZ9hb3SV9+O09cU2sQw1+RNJN+oacEVpDpHFhkWQg8
uTJP+6ITnVXifbq+CcGYeee0FYbeCb5iuYB8yHYIrXwiCKM8wq28sl1e9RXnnwEG
dYjBFdyBcDAtB+lh/KUAw9PpEj3uOHQQBeenkBi08bypOsO69Ts5GOxe1dcSx6BX
IejbFtnow5/kJLeQVYtkRNnD10U1wU0LM8U1zMyCW2hPruqCK/OvF/Gx4nddEp5t
rWX9lKZD7y/nSgP4vDHAZI9zFFnRWBaCxE+lzNFgXa9u/lXDwOE1jAktV4Nkv1OZ
4re9jssV2JAotrr4G3aiAHDIvvoO03Kpmq8YwVaylC/1hWwkA3j0JXInXktSsixO
XhGZEj4Er8dE3ERRnqduj4w9Erjm42K+DhW7NFH8+w6GTG89IklTUPxD1/GREBsD
ulp/ykWXNT3sLMG1OK6FlR7PDBYgnSe5eXmBWiYjj+nOPWLsB1eJt5LgKvaj8WWr
JblrYYbdBzI8oLb4s+5pXqk/gtwgV5ccy33AxV6QtjJKUL++QdNOWBfAfyg9WHLh
hYOVzCYrB09yafuWKvhZuFHbIml7P04g02Q1DLzR3Yrs14upMzUDgLAURyyxv+Le
BXa4uSlNQ7kY/V6qi70u3siuHa+e6Uc3qvrK62GJqD1NMYfKhGlW6thAcy/gF6uF
IW7oMUR0V9DX/9Ql4qsY+ZqKXhKTsv18jfe38ZcYZSWgN1Pjm2VmaaBSPqjk/wxx
3sUTon+0RH2pLFVk6kiS7jWYFQxy/W7vJt2oXTVeLqRb3vRvP/GwowOsPg+oY18H
tKWGxoDuE9Pcw4nNCofTiezGi5VDSfgog+25Y46D29URrxtQpAginkohTbJq8emA
jnxrtAXrnnyZS8btMjh/Ti4+RLhlog5a6WzGD3CEZ/T6xLzLWGztR86bCATAGCzd
CCydp4qFgyrUtwuSsnukprtqK5PYNtXsjMuTZiWfkPC3I3jKrur9Ys5nePFaLbjs
b2cg9RNO5CgeNwvqitlyC3kc00WKmqhJbZ1AUh7nlpprTuayQ1h+Jw9U59uc2HbQ
D0qCUIU83Z/OHZLZNAHJs+hK+0OVB2BL3rIv62g7GkuWzLQVtKLlc7GwineFWLKh
YlpDWlzz3/qC588SxaL2VXtRvt8p8aR80OzR5G7u7E7TavgifT4HL7dRoWEtF6tK
FAdbM+kb2yZO7W/w8jEzImoNMcXgl1WbK2OV5DCGVmqL8FcW+B3ZV1eqOfOKrfKR
asLbVs0Kvcv6Dn8orYq8LedecZ4whd86Brpc9Pll07LURZ5vjjUXSpzsmecM4E0K
vveBYx4DsVBmPXowKBptW6daZUD4vB67Y+qt2d8170/wZBUABrECRt7srckrcrT9
sdxyqEq0L3qm+lSvApFF/PxYEE+K+HIJQ7NysmkVNu6v5JAAe/NSpY/x0y2XIfpp
vR8hMlmGsmCn+5iimVNn+UBkkcF6snxcn8nNkZesckb5fPXHAefWlm1QzUK07rY1
Zt9lz3By1d/nY6nWAuFufYLX9OOvzyMiDjF4RjsnvLQL1+c1bsw2FZKdoT0tQLBU
iKDYwiw70PXC8MYBjDY7p+WMl49+DEAjDnTmeo2ysLj0kNdd+5qyZIhkrLsaFI9P
uBJDfBpYNmEL69HKUe9JfWD+NB5OC+U/ePK4pFCUz6FNafy/Pvd5EYEYf55vAQWT
CKNlXphzTV5ML6jfYTCL2OPUN1ovIwVEoRCZF+OkzdRnKTHH5XM5wsCKGIhHbAsI
uThMTRfYspStzb9QNgfhTj2BqY+JDi2aNLVeoZ+TQ0sbiHcfGBFycU3JOUldu5Ko
X2ty81mfjkbTWvmi8FZCYkeE3bWxfRHaBIFqylAgHjOwD0O0NidHZz6uAnBeVISW
CpJisNIMi9SrORgngNwwNdYBFjkQRcpxPJQvMoVcy6Q6UZkIsQQdBM+onNOw7QGo
bAPruWxXL64uBLY6yLDZck6fdqN/V7wHKOwwEDxLieiEZ2mXAOJlwGUiUDkptxlb
GKFeEYiqaAxt5loVJp1bou7xytNsif5NoFL/JQBq8SnrUz3U3ZBVAiprXYbG8fHw
21i0MmZkdR5yxq+w9XQ8IKZy6/VxgglKnTaXJhR2Ts3G9k1WvnF6pekDtUM9ZxDh
bOc+tELU8qQO7UfM8cX04BdiZBSenpbF6ZQSDu07PZJaR/X763BO9Qz0xoTkmP9I
23wdGY9oAXd9fmXrJwzK0K3ECBQRBj1VX2NiiekgBgMXRYdWOhGvjkbcP3cfmnFg
J4X+YIFduIQFoNE8BwTiMpvO5MFPgvJ+q2PjwtSuje6oYEYQEVp7pQoYsy/WP1IB
HmfnBAcUbv7My3pfxAhI0DS4LD6iNminN4pd+i8Hcd2v3IP+EHLtD4NhTeK3e1a8
9aOFDz6cnBiLci0dMpyvodvuDXSTa2gDL+uVRR++6M9S47jy9P9g42REqsYFT0ex
anj6mp4HOMKvcwBqtQH8qSj7laXa+5QtDWwL3ZjHORecBEExd/xsQ6gtS0gVetQY
pZ6B4FDKy8d/PlwBedtXXFkvGrwz6r4awHkbVL1jZ4x47ex48XS+t3AdTuwDjwNw
659cWEwaxmn7wvOnWuhjRI+fzQlGJ7fD5Sjy5NTKnZYJqsPVUks6dl+nTbl/aFCM
l7ueOGuP0A3r5uiUhoDI3Cx0YZKyjc4EAyXC2ebFcACw6qpgSahjAc5GIwa9QPGA
0X9P2TMIPA07RAp990CEkDb1xC/TxcL7Nn/0zVJHWhmGzTYzewQbmHQ2bNLm1mkY
GS7zUde2tPdhCR0BfCu0Gkkd/GqnKhaeizeBGhE3nb+UfZD2OPQvzCHuc4UnWj0y
gVp6KJv7dvUdBetm4PJ/yutzUoRTByuAlWPJ5cIUwZla5ALiH6mqvnUoy2GvTZKD
aie9YyCB9gAWPzs9eB7kz7Q1M3FcE11mhIIU6Jy04IbjN1Ei7soXexWDFK75gFfB
eV+Dr0WX+1FP9EY3iTVEPZt9Sn6nqziVkFL1BwYJr1/NN1pe0Gro0euc2Oci9hmp
yIW/riygyM7/q/mLFiR4tBueWXVLU+JYffGKyhSqlp1xYsrbCrDMrwg2PB5AxvLS
aeh95dv+CMqHZROFo31rcaQaYmQYgtbDpNHFd7hWUP1bFw27LJFR6k02VPh+Q0Yo
LnJST/wMIKQJXAbAraui3JKQ7L/fKxaFKdyS3HjndNxOt2CshegULT39/vthklna
v94okkSnGyCMhWsLYYs+WcyS0G0u7B1/o6oKd/Tp3S/tsslY/MwzkZZu2r1kT3TA
4Dy1oOtxZiOPmbkqdXZfjoxjtN5V3TSq09+T3SQmyPx0Lc7SQtSDWPW9gaoX7pvf
HvaYK0nFKVGF3VHtPrAcAoxCyq4hVmx5MVdBvtTqLaTEkcNCJfJKUr92FjPjklNG
jnAXqBvPfVza2vn10GfRxakmf/OdfaB/wDLaRPcqgJEOKfIt9nIsuojTIyq7UT1k
o5KydsY/Mmf+O7syAK7yrFGCLj121WtzC1+EENiMcvND4muYP3tOz8F45TJQzrPn
ZcorivpLWFnMPHeU9n6eoGfGTaCxxyXnBIL3P8iJ9WGI4MipR5rLP9kEHNwwhxXR
NY/Yvskt/CPFmQHtK/7WFdKtnxUpOuPqJilcDIfe14gbwJ6ZYW0Tjfpx5P8eZIDw
JMOFJ8SgvxOi7wulNTD7P9ByO4U16T0VuL1IEPVEbWoUvg1ez/SVrMEJHIGi5Fi+
ON8lt4wREqcl7t8PhKoU5tpANWtJC4khRtZnQqq2EniiNDiail8wEb+egV59FmPI
lRYo03bsMGze9jav7CgC/93KoafrxZmd/Iv4OHPIY1exbIuSfu84GUslCmyRDaod
VVdGe/E1UmUI+SK8xKULHFcAgK5hzB+WwpSfTfLoKx6CDhxtdiPCgUXmoCWJryEU
DZGo3m8WeWTSkGvceN2eQfTAxiLu0wTX7HK121vupwiFEbf4vJPmUDRl2kfA+Gv5
9dybrriYw8b38AVhOC3vghEEkXfJav36OJgdovvExOZrAmRkUUyCVF/lau7priEB
8DfeOX2XS97EsWKHzd8AvYobp5XVyxYmJxsUC2ZPXMQqEbpu/uLk5xbORsuQHG+P
HyXc/2QxXyEa+ho8BxFep+rGLzcmgb7Jyn2I6hkh6oNfDxWMOOqlOIy35sH/zs3y
kmhOocWImbN0Uh1jIClVbQdeBNPplK9OJqk43OFS/TwSS4EGZXdJmEzLo+06gGr3
Y0MT+yTYcihP00+BoKObVqmru6L/KPDxIz7IRhg+1QworTZr312WIvBYO6rTWL0R
A1jbJFw/XrEb4a0Nve5e838/ZwqQ3AM2BrhfgCCcwkveTlpbC6ga4MrJHYHhJ9c+
XcX11Lc/fhNCBH08RHUb4fQebEOp1nN7UfGRfuLo6+zBDU28hmcCcu+CrXP8UBTB
26MD5I9GDxcqHH8quDGPnin/ZoGcx0upLXwTUaDi91tmnfFQ5AAoXAGEK9dmgJTB
q19FQsW0/IROphcOJOOPJCywV2zlUO+HKqC/0APrzwkBjZL56nS9hvEleXwqmddi
l2KzeLzn17c/CnE9ioq8JimL69MmB2F0VJMp6Ye77cMujE5GIci9TjC9Gmo6v0Qt
Y+BvwC6ejJrt5vkMslQX/2PEq7ZjkjpvAgZSl3BJr4V4q6y5kogE1am/sZaP2mvR
9+uC6sV6ww6Bj2pM5+dFxAri2msYF0b3m9EOklfeEAO5y6Cg08iuuemQSQsyEo93
4Iy9nCc7pxYxWwZi5QlRw4OCapQznZNo2sQtuA0Qimf0rMDiOuwN8FiKr3azlk3V
mmG5/IGt9lEuWfvQz/UbOXzLODjmb+i0rRgHebGTZSoJh8HjMfCCQ9/rEVsYaZgp
TI2TOuSHWbWSLYBt149Q1cPdvPEcxQfg3hLO+97sX0sIdORAe8jBk+HfV9hjh2l5
ZqmX1YKV2FFgPkcRc75cfyNSIKI837Gs2azWW2d13zQ1Dx2O+NIsmuDb4ix0iuqU
xJRXATfZWUVmse5xjbX56FXFzzBBr/LrXz1DprjPPG5PuCE9WnH7lfa5OBI0PcyF
Iy9aw+NkQVsHVqZ/yejJuYLxWpW9h0NZ+Hh5C8wEKTb+B7kVKKw02IcHYLwJCmAv
8fxRL0GqJx1vRhJycN2BqxolrPoYbsCFEmFE9qi5LV6FrPneT7CiB5GWib7Do+GO
fRwZjHDEFDvebhj+5Bw6rrCdFhmE4a3zKkkUO6NfkP+tPVeuuHTF4+WDPwW8AUkb
aFf1BRTl89om8eylgsLGsKtExmdEwQ8o7NLZKOhPAu6E6ZaEb9X8/K79axTmI8Er
OsLmUCpo136etO4hSci8eSani1vlvEmIX3kxzSKiQuAPh+vUqzmf6LX4euUFGCet
M/xNmitE6ypIuMLTEokWIw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
PLB1foTbT2e/2U1LPvOT+sPTIxOlk6iYxK/G17tdZZN0FovFJrnnwNmq8257k+p6
+WOkxTtExgdUGZVfumB5gQomHemtiIB9e75savTTafg5IsGr+pop0ehLAAzxrqsl
jtBW2sIO6Nntmgz7HpxFTkEWWAppoUXEo9/quld2Dm73GQ1G8EC0Y1oXFETMJIve
ukP7vqy+O/Lw98p9CV91urDhXpYC5K0sCedKgBaz9vlWY+QsLMKFq5tV0T3Pjv4f
5yIwqrTcS+MGqPkzJn8n4V3YvaSVSaDV6S7imqDGpGfZ2/TQdBV8AxfqghOJqEgu
tjHmdtZKrqtueXYHmNugsQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4976 )
`pragma protect data_block
ZWbt7HTGc8Btt7EjtJhVlnxDNtfOQCw61Yw7lzt6rqalMKtlqWtWJDIBpPEpGaSA
Gy83CsQ8HSGLNE2CRIOnUeRtuVU5DALPF3YdkxWoW9qWl5i2Ze9fiWtoTXF/HOhQ
7Z1cs0DxCObtke+dMYlG3PUuKjbBSWFOqCHJdU7ry5jR9vGE0tNgzD1bozhuDaLH
KSDVQuTuXHEFpp98iwMoQm3rODuYgDjAI9BEjgd9YCKB3qq9B4RiZkIYtb0k3KeT
Pvk36uxEnHOpqILE45DV+UU4L4f+ZM6kJJF4/grHJ7x5eeveAbUjEZo8DukNsfP3
JVhGxqUdeCdRTqfmwvjn81tqRnWvlcE+JMnnRLt2EXXuPPDrfzR2sjeSODYQUCLK
rwLnfwMDyTAlIUAyumrI85Vx6ZaBXPxqUFgbKc2OsYZ50+2t4M8Ap/J27sOWh9QL
b3A+mTPNA2btUDOfJcL1Aa6SKlY73fQtm/OrOWd6Dn9Ui2BaH1HdYxu9JQqyWoWE
BiOHyTEqk0/wu2dYRfODhgcsaZlRiDc3D0I5Kouzvd7CQ26JwdjTd5JMLICyEKZy
7yX9Oxft230JDGc89RTLov6JFZUdIUcFGBL6awiXyFuB3E4aBNtiiU3RaQJtWHYG
TjCvziCdglFs6OfZNkj8ziw4uWv/qK8biV3arY/URBsK+7H2Aia1/x9qQM75A75Q
KS3oIkqwSeaWBlXhIWm1j004QmtBXAtwT/nj9WKgdiWu22ufpDVYBdxe4C+OVh4z
xruZ0P0Y5iajRPb5Ef2kfB4mKqhPrdaZ2D79oc01xlyNNwU9QLx+eCYITL9BiTCv
Te2GyxPxp5C6DTVw1+qHi/5+RSbSKttLN52WGIW2/TLUqKLfPAZ+JtHyc1blnXQA
ShQDre6LivtbgdZmdacXlj5CawogPwD6YjHdhWHkqjnRd3D1QhXy1WOSN/gjW0Nz
AouQlq4pVH8THQweLf/Zbs3f5vhSCDceg8FZJqr2as8TRlzbRnouIgqG4/ijNvXH
ql7QkD0vJH/LqDtaOHq3Z0a1uOVQa8F6wZXdwzZCb9wqgTJpipjrxYhMNpK6rLxS
D75462RrxR5wx2+XNzykyPWY7RWIwVnmkUsywhluYRSu7zBZY3RECTzMxm826w/g
au5htQuF9ms4w++IGGZAZduDR3PlFvCgXX3/oi6m89wiklIdwKKSFevzEREoL4MR
VBVoBuN7RqRsTrZe7js7jQ6cWdFfwUTyt/rAEDzZIBdZeUtyS2+kQDST+Z+GgPu6
8efs9g0zRbIQvQDNibib8JH2Jbn5xtOvIRvbNzD2aSasaE5Z4U13Xpj9TL5ZywvE
1/QEA1wx0l7SbE9TM/fKx149PH8Nd92dEFh4F7NoY93tlY9SAlrxEbGNn/C0lH5c
BdDczoNMv9BDZkPM68LhYpeoQn4vcyO+c96206a4fPklsCZxn0RcYYEU7l7VLU9F
M+gYEALvFyArLDRl80dchwhsmCDARUCWJknsSfM3Mvkg2Wh7xCLEhEzhjDnOSBBE
9pGnQ9v5gq/s95OoHRA+7aG0fp5D3Q2QJ0ZBA7asw1FKxmYjFzMFoWGxcBQ4Yk7w
6BWmjatOlmtkdpgsTGBvoIvezQIWexgxN7MXjdl62zEFxQFf6dcpZqUpwLx/NRFG
+jI7uhZl1khGWaBwrnGKlpAjIEsN1FNn1iP1wxgB3RegwqMeZ6yY5R4tgtVkxoGM
MMS8gQm79jaOgK9PKiJvFiNAe1XRS6amQx0WXHG4o+IBMvpVa3dlLJ/OFyHXjbl1
0o98GVSeQ7Obd7ZTGSSkpFpY/CCOyMMUSglkvlMkFoslgZA8zQaQA4CiSKETGAEy
mlFTv4+gjKQ5/gG3cPZI7adf7z8dOwvxG+xFn2CZ3Z5JmLthTwatYkMvoCQO8EQa
YUaj3As7w/vap5xJ5b/j2lIe1dDtwIth/UBZkLiMCk0WHfqvUSlPvf9O13Ty0RxS
fmOU75pGsyGJkgU9KZV8s4Qw3bcs7KKxRAC4Is1/5/Y/ti9YUGqqGGiDijiOIO5i
vj5+64KRXQCo7M1pBN4HXm7OxI32ocRoelOSRiabaX4ml3hfA0aT2KpQ4WO67KZm
SLn1jFF/WSTsTEG7ul4GI7it3iBkmhG1Xxyc0cEyxb2E8URYnzl1AkxyGjYz/jN5
Udhsqh7C77ejObw2PwQFzBsUClbyFknPcWR0j04lQM77QTJfz7O5GEvjtTVbAZI0
g7GMntemgB1AzPssxATs5Vw9fRTpSEBliJQff6Ylv96JpMJwyK5Mq3bTiwelc78z
bvIQd1WI+nkysxVYXhoLWrRYoGQMsF/e4rl8X9B9B/+zc8v+FfBxY6YffSt+pJbP
QSC+FNA+6A1kWJAMgILeXFjPUsV0IyW/W/+oANCUH8T5Nfu0S72JiX9mIAvHDJ8O
IyVyutSSG7RVj+ZEjyyuvwE7xiUSYmqyyDLzTAFbBikaFl8qA7xD/7bQ2LW00GuI
GYcyTOs9ZwB8K4d5DMlse1kgeQBK9W9esu8uDg5icxEdcUVlB3hEZ2zLYuJM5zZO
8cYLFGhKdU7FdS9W6M8gEj3zrTLemRjKKIp0dImfaCb5lFmoUPsnzpENhDPcytFR
AZN5/MzGUtSCk1XM6qG0S8lPTLPIpUxXbFwAvByjiAJfljzo+ELOKzAQDYAyjsfl
ed9/2z72bdYCgGUWqqqqPUbvVkJQYv7bYswDfivkgY+z2IcoZvn+R6gEp94lL8oJ
HJKRjNkW+rzOm58m2q6mwKNMj6r1Mq61e+5cFJq5UKaRWaVjfo0FodLw9pyDtm6/
ROeuXJ3PglqP/qWjSTeSWYhCXdWY/FxxlApWk0kovH+Lbs8zveaxA436za+0eENe
Y+7ZUG5vZ1fKDvjMxPUHXUg7MPr84PLCPtxATZmiRt1a0QFWO0E2qFMqPc/FZFyc
9QroO+85rS+yex0LYGBmKI29JrHCAA1fN9ipa10QMjUUWgfbONnsYKW2sL+JPwgP
RNulabZkuc3nkDfHmveqFeaJK/XvM+rN4XAigLYnsPox+Z3SmOuEnLOl7Pon528I
1epXayUOYclckFPKZE/XuzW3iPV2h+/Ng/w3CpgoX1QnCO8SKuKbQRJGwxZo+ml+
D1fSFOaVBIoJI7w0kXv+mpaV4hv94huARe8NWdUTh2dtBjDNbY8BTPe06NnA7FsE
F6BzbxgVFMJOrDl9fuykN4UFZP5EhaZArHGKJmPRM5COA381IV1lQ+4fhVIvlMI6
hIRNxS/z62GlLfv/hyts0/uJjGzLbhIvIrPDADLMV3iJZtJgFTVMT/E1fcymTncY
HMctTeKsmEDLYdgwChquVFpBgwFjOt+CC5fM9pHzKABnPL8g3qeHhye8U6TDN7BL
X7AWyqxwLO3R8fsGONyb0ErxY/7JMetdD+zhtu6Cdl552gKa5se/v4A5HfVrR3Zd
hJT8r0caxbepOyXs91xxyvOsv7Vb8j1zzeKYad6/pZTuwvHQUHugRGB0Eyrfg7ja
z1oRowjRKplGWf+XveCXp74SW97PakTEs5kJl0/6+GywMtMgET7TOZCWfy7/IhQE
9CNd/ppZDYP/hQyYEA/n/HzoDLKScP2SWXJztva8LzfwaoWNml+CMPigCfknzWuA
CkqRGxkxc3eQu6KnjpWrr07GeIahV/D86tyVxyXk+S92eiEY8mq5OLhpGlDLa52x
r9DsKurrrCv+kQDKMWorzvyIBmjE2Db3ol+zndP6dbw0BD/a5F2Qo/MuHTP+wolh
39USRgygnBYApXy1UFo50GSqUTJyCxW5LkzZ96EiD26+Lm8ERKEPyGAJ/TGvkACO
kOAMg0OHrPdskDQ/4lFAANxQOEY9xUzF/WVMsz57telRG/SaxiN/Sc8wx4rTiQtc
FtTMpBQhOR6why+50dv2ihRY0vnZOY6Fgtmmd/rao/YZzHZ5IMl98czGt04r9Dct
AOyxJAkGTE16vhec16igTHbf6mLHmeTnf8vcq9xJYN0WYklbLt/7yjphDqJ8s9Vq
PRlW/kHGvPOww7fJTzcwp2fZTWYEJR8lm+rg+EANLoxTLbhPj9KE0vatZKyNEdX1
UKPzGtOx7Lb4agl4HE4pLkPbH3Yglyu40D5ksssNaQYOoYxDY7uxfoOHplNI2EmH
F0vUpNEx0rqy8h4Hs24KwRv2gBB7vZRDJtTWtMUw5RMA5FKf0Kud6L2wLws6m4n7
R/1y18H0l4vM6aWEefKQPKhZBd3xbg17nYExRJ11T27Mu7V2oI2Sqvnl5jkPbuM/
J/B20seiQssvxfjyA2dt/V6VZ7WWst+z++jVy/HfHflAZiLVIxtqJDHgGnbWXs4L
sFqQPkTCoQrsODKEgUt7m6/VY7X4zzClFiagSNQj1Q3c17zbt3VaLavNrUtqNOaS
PV8y+bQOvyF0dhn7KbN0kz1q0QPfA7++PZ9Qf4dJB1ofNeNnNwOqCT5Vi+Zwb8pt
o6tZF4ckOdUkdR4BQJ9b9tlhK7NVsvnekYPb5hR2MVvB9mL+6V/M0Kje07evVvwe
sELmcwaXL+AgnT9z1cfBDmm17uK+peL69HD6rWJElAP2nnAKobJmU6jN7B3TqTJI
HoI146LZWPhIW07C1pXbMmo3RiS271QzSBE1ysu1MslRydlJdFO0MJ5GGW3rrAw8
W0G0gdN2zjlXc0hAl1IMyeVAioyHNWHYEl1fzuZZpGlgGlqDycma7hV47Q7yTyZt
PbrDLom9bkhYzsQB6/zbXkLt3qTcsNuUWWT0TMd3tWqZ7JwlcHBBJyePgMVtX1o5
FrlXAEIZLN5N/wsU6Ij8AAJuNNqlFWdedl47HVadOFR7OCmdQxtVl1kNr2z3q+l1
Mb/DS2UnvCYHg1JFnRjDTxAYv1WCtGQSEaOyRayhxQhp0xihN++CAEjk54IymkMI
kX9C+DBT1FlM2AVrlGcFMULcfWeDs05Ao39sOJ8cyY1/qRt8vezNvBU5yrFjvvFo
XQQzLjG5YdAIq0WSM7jd7r2XnTK4dT8SpDLGIggcS7DuW2kWbR9WRr3xvnZ5vL9O
RthucU66OkeS8/5Y9DOi1xwl+OHVNcist00fEYLYJtCgLgBGslt7/r6GixaLrY7K
QKILY2GXe4i7vh1fpYngUluj+CaTHUlJaKoAgU/A/Kv5oXb/V/Joy1qXOHX41o78
e7r6nez7JbvPhYl5cjnFvXrFQDM+PTVSStBUimwCZCc3hZIpkmaBPrdrea19K7Uh
PaCMYbQJDj4sADhklAxmX7JOX/IQ9EYtQjj1QTqaFRnEgFUOOmheIaOM5HuZ4XEV
5iAYkpO7uy3QqX0MfLtYWVCbexWHyoG2DUtzmAfIJKlkEk5pr2d65Lt6rIl7xrdX
+ndN04ffjYx5LJQJ7QDBO8eloPhMepfDVjTEGVR0WR40eJv4DTdsobK1xhC6l4gL
bfQMWj88ur6+H1Nbw+pmv+6ECJJMAVoRf5DoZ/2yvVPPWPTufGLJw1I45lanKi7j
G5TanTW3mWj5vr2975lcjLz0+jDy8bOBbvI8aNhaKKRMsSya8bIDtDJisiPufOqK
AVxWV5BlKjYziGMPUKPbhcIJ79V7HB0UUkfz5ZLG5j8Vw6kaLcgPQ4gFmvJWGbPl
IPJQxCecVzQ6ylI4wB+qS5JbG3wox9JXBnNs0dWwjDmMpr1LFKLkASgshi+AJo6b
ZM+5ON92BKgwKzwIcm3bxlYGt/WipM5AkFP4ERmng5U2Kiqx+yjmPoSYWT/WUYGS
Eif5Ln/vhv4HKA9B0M8gBg/qNhT3QllrIDk+jg9zsaGc4zThn+foDoket4sGgKLS
UugfDH7pEuwQ4ke01YGKxQWkBFPobZYsQXnhRA8oObcaZqcm3Ih9GI0KZJ9ymEqj
J1jG88wS4TDsJnruobIrRvTHZ49R0rT1LANtX2cPXDpKBZ21SvVZkOPEqBk9a/kC
ZOSwucpVQogH8/Wk7sx3wvUHPqAxA6pTFI9c3xD4P02DQUQPOoShBJV/FfYrsOxD
Hlt3TYCY2Nc3uQAmLsftrIPPLH/k8KRjeK1OwcBwwBtANTcrIOOclZWg1Z8ICEhK
eR7I5+rUD5Nk3Y8/23O/GthQuxioWK//r6ar5QIb7rT1XThVVBM6/htF2vCl7dpw
dqKSWebkLvDUKg1tXXQCTzCRVB9gZQaIwYqX1qG29cvCVd9PdY4tFJ0tHgPi7cc/
zhMlFP0oYULnACfgrfpajg/nfFh3zCFJxPClfJFzpKLnvSCqQlgjGwuSJQ+4g6lI
pK+aNcJzMQeH7UMT/+7n376t6A1JchfCcFvBw9fWSejD46jUcPZQpSSjO8H0r8Io
JHpUBxbqNJNoepFU2GernvUGPPUX1YJkm3Ta8GCt+4qkqLBlBVzwqgrfGAvzAJzj
ihSdYxCZ9CgISY5bSD14NY3bKDTZLbjGMx9UGU8KJAey8UmaXFpkHA/d5Ck/aHHR
factYbBqcxT7Sf84GpO1nXZ53dLtwLO1iGft3+eiMLd9DJKCuvoM/vbhOJ1UmQP6
2fxJ08RniBjvPuxatCHDMtOdkY4ubf0L+Ux/2elmX7zsa5ELc4wmi7d+x386AxYb
MWTJ1E6F4m7m7B9cACtuubBudIWAVVsDRUxJcte5+gU=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
fI4Gkpk8OA+wksTVV5NfqAdKdLadkEL+bBVMGCb4nLFanAL0E7YnEXDB/NQSXs3A
/k0QsvvhnjTmoGBT/uYicpY3SFxQTCftFainQ+u50jShrAik0Q06UrBno9AXx2VH
1Q5RQIy3hPnvM8L8P2HuUYbWviyhrf5YU2/9MkaeGqDRu4GiYnKhRXx9rkaRXGWZ
0G3xXNotukYDKJa7Md3KQbmJuiIgUa5NsC5YOwcZRBifA/YyjlrYnmaH/Wd4Bm0e
heGAtzV54bLCYJiSMAok27MT9a8ta2OsNvPf04H9o/W6oaUj7myi7xa2Fq2oNRQb
5ywxJ/Ust9b0waaw/F8Xyg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5344 )
`pragma protect data_block
WkNESu7CGEIexSi1tqMnnoaInOTcUccBWabnUwlSXfUBuVg+AImDLN08XzVoVDO2
US0wqY4Bf9lpmFBfYDDxaGlgJZYyG3yKoXWZkJ5zNgGqRFSLZGYWKoeQDgV6ehjx
7DgJLh3vbswMW125sS8rlFwsKW5WL9WQ1eAUZOkFs4T06fPqvjimxbCw/ETQgMI8
e1PthMYJIylJAW1G91Z6dN9J2OFSVpvWu4oc4wGNnvzVraPwypubFWo+nTcMxJnF
BlxtiutuF3+on8uo3ohgU2yRtkSKhkzaMJpT3mhxlpwYYDvQkOFy/UVoNZejuIW+
s3TKUXvD3UXv6kp8MDYFHUVx9zEb2xTlgCVqlKVv8YdhCaAAQVIW0YXn2yhXa2hG
SGAtzxPTPgawTXL8FDOK9/zUaOOrBW5HxfP5zF8ncmv7SzhoBXvG1CrZPfNatuq0
v7iSpFurfTISY3CeQZt1n0xE0RlAZbUzB+/Kb+1pGSa5feUvEaiozK16twbvDUe3
EqmQ6cufvO1bzg+cBc3TWm3XMqCurg1JasFf0l6qOKtaYWGJoUiQjAMccLxHGELb
guFAl23rTrgLCyhnaQu5AfDp+a/sDKXFN7dAE8pNqugP9mXuGAzMHAHZxAH4qSGw
nzRbfqMFJOfMhGYqOq8bOp0qVk2WpDHQGD4y3aMEOFM9XsjY2aWxcwRdKXd2L/O6
zvbX6gQ9f4yupKbAy82S7Q6FoiDgJ2tvq7kdwnOj71z3U/cdLOz/iY6mGUTtYJ/W
1HvdxUNk+bXNpEvAi2m12fzwqREWTscjfvuEWej4smCZwapizeBf2a6MW/1Xv45r
5Tr6NfEYQe/SSK39CX2AA6YSrh3CVvInq8sxGdhIij+eY1guu425khyZ7tNUc0GC
RemSPjY08pKzx/MP01RiuTK/QzrlZoaKFDxyGeSIzsHv2xAMKWOWnq1d007Wldfx
/8QDPfPjf5nuM2sSzWryy+1BOh81KQc7Pq1ZyPE8AAbXRaPBEMaHnPJJOtCEFnA8
SI+C7eDbYjZfM4bwabKG/xjP0Unh20GiXyd20RO3iRSBQQjrv1eXqZ5sWVRQHyRZ
oNl4w0OUPz8lw5on491rDl2AF8zEzofXvCS7jP+BcpPw8YNGhxIxzvl+hpEmcCAa
lD+6chorKYpwy3H6v+6BSNO6W/31PS2vWAuBUQ3F9Khy7pA/IyBmo2lTgnty/UuK
35c2yiEcsILQRelMku9VRmDsGu6tI+Fqgk+zH3HZ+f3K4BxlKMIlWwLL15iMwyeT
06QfG+yQMqH8K8BDShcssDNInO8/x+AlOJbmSn2+Kx8SuaL3IchxqwpzMJlTs3zk
cnZqclhDRw0RlTTvjTwygSvwA4dsRbi0tD5CkZ0j2eo4xN5iJAwx4siVf+YojUYe
0LsVmZMiL2WmLvlnfC9078tnQwk+7Idly7pXxZAKvnn6E0rgGgvLmySKiK/gRZJN
5gRDMvVRgan39IsHXs+gYRI5uv60UBzmlnoBUdeyPPdjN3n07nMNauTuVtqE8g3N
zFUftxPYcyNi+cInJFckGwjGtdMLXPN6VCWch+QOh47/VhM9M9vt4pZo3Phnhc73
cJNpXHzac/+GxrdRiZIug4cAtjxKTG+3++hWhrN/ka10LiKMvCwN+xaFkiisknjU
F85NpH9KtpDASQcLxJkutiPn2K3Im/gKgda5TahO0v+ku49tMDE0JVUkhk+/J4WW
DuBQkTpxmOiyQapJP75vbjgyReEmoCBw/KSrMFEWyTbe1AYEx2UrLxH0BkqdiHRT
fa4yrllKcpqzeQNEvJHLN8HPb59cAiPpoeakj94uTn7TrWvz9Sup/1M0vA828ade
TtxY8ZWYSVD7MqRtG8Xr1d56CyrBOodZXVJdJ0HRnIsJMOBW23lHgtpz4oed61ID
V1W8SIf4x/Gd0HxMSzYWEYho08nE8ahQOyxZ2c6RIFsT8ToNmEciHfkkm7aG81CD
8qjCGV225Qyg2jJbycWKJF4/SRWeB22a88Gq41KIwrFh4bG6+ltgulWQLQiwJAZt
MXdMgx7ZWM1IvDYqr/ZK9+52dpBx8Qy5fi+bPx1jVRP//TMK2vwAPeewEQme69Ds
17Jrvvu4c079egdX/uxIOFJr8EPTs61d72Nk5ZJc6inZd5B5ULyFmY5uBbGcdpPg
phAZJU4DalYaqmLNM5kxVV6MwGSQtN9grFEkNmGBm1Tr1pkgfP0nzQTBvpmp+JSg
TEb9GHiJUYPo6VPkp6HoSk/qCGqXlGvopuQ5hsTmyykZXoT4ZkZgqcHBOfJ57LFW
pXPI+opMnM7RJk3/acoWjibmLIXpVQe6xRS7A7NVvjYzSjrRBUzloF7gAWjaVZs+
dmeS9r2dM/G4yRXSx7z5Y55JHgxQesKbesRwu1mWSkrLINoCKOMce0eizH7pwVgB
6HMx7ueWG3HiZwPNGhNjuz/jy5xooFIv15kaVxbhgAExIfaNivnSUw09mIrtl5CA
CziGJFvteSKZ4/Zp9Mu0wTruvBgNOPZ9vkPThNqz7gDu+Ktmhrj/aLF8SeabGfpS
XYl6KIvCAO0AY7L79mT1x5EfVeramG1BaDzVPw4hYVo317/BV74EiTc32DflMaCs
cwmyUZHSmaDJ3qShRMbVO7rS5RF5zJyClDIjpZ86aLbfg7k9alX3qmT9lE+wYFe8
J7Sx+NhEk8CjpB4C1lXMlfnl55C7v8v72g1aUQzpyLUehDAjAJDa/+IlFQ0I07HX
lT6PwfINbghepHEXWEVP48PoJanLcq/RJ6F7jjACPZy0pxvMMkbh1g7Bc5o05Zj6
Y6l+BfdIN/XODyQtwkDfPReLSihFECr46Vt8N85MtIbOvQgOXUQIKiinYFLQygvc
O6v+onqA2USI8nYoEu0Sh3yOx6MwbvYdy5vGAawsQocnKJhLuQrcFYtDgEFr36VO
1FR7dy57CJouXpQ/J7otD6e5gaSfxEpOXFwT9RV6h6VOoqFhMmQxUS7F/TmyOXlP
5iWKu3vPJCvLkx5FpMl5/j2mNguyoZ6etYHgh714SWk9tjcupGBoXRCHMnV/XOZE
CR2zNowWYdxZHYf0j7RpUhi1FbJoshSd85dxloqZwGPpzMGFtdwodFLn3Kq7sD4V
lAFuzUvriXc/8v9FJkiYTFUluXkqrZLUArhVT5IgZksNjVCBWLq8UKEFPKAP4zCw
YaF/+OOagKHGFr6DkAcaZnwDrGViiMZ2SyLOYoyviVEIs3aA+FM1dqwbkg4vTxHT
YZvSAt2obCH2jz0O6+f2MLbZeYKF+CdhvInw1HLU16ErSOKLQ5KHsJl+NqQnNSXG
kLBy/0UC0Oy5rx0HdeRIGH33ya4KeUJEtR9THSJ6o93MCZNlriYJaDfWWkbNN4R3
lPyk+JVeFjL7m8o9ydMfQKLwyvDXLVpJYM4MaUgDuTuK//7amBEY8p/EUZKrgE70
vL21Cnk8POb9Feb2JXc1cBq6DRQD9plaXPuUy6VteKndcjoa0khBiKX5ldIZuq/C
sxv9T/TWY2Mm2RDoxIO2jDoZuPWo67k6CM0raEgBC6OALBYfbeQZ/RkQFARmrD5S
sdX4dgXdcxmNj54VjiKINDDfIAHpAzcU/Hm+VbKF6O9pi7QPeexUNQCrZhv+cBx+
zuxdyZRv7kcEFcWCQtxU1f3aup0JHF/cY7giACQT3uVVyfxcPLRq8xmf1+33kwl+
nWwpt5vWoNrSHySfnL4RezRvMH3Rvjol7cVfnCXuLRDNfltMb7aojP+2w0ogZYsd
MIKrWrvplNLRG8PsczgVIfKL7TDvPndIGpTqi2AjKgmrdP3k51g6dKM21jpP19DK
AF3XN+rU40E5yBEzq3Dt+nJ+/g/+UQU/S9H553M92FFJDK/WfwIGOf5FrdDUL5pe
AXIg5PaC4+axlkNok1GhEmVWrCmzazUx64R76X1pSDj/zhW9oiEgnq1itNqbK0QN
p6Ok7D6l2nHs2dg0kgkdxn7OadOV47bEjVL7eOrZ7Iecbn9WazfLqj+VRxoshIOr
Dd7Zwq4HibOpDmjKc+IjLhGmBkfb7b8fX/5t8AfLb0o36HzeuRpA985tnCPQ+Zdk
G+ZjEw80elz11XCzbbfqmBrsKrVCuCG4Ac5G8Brs1gnMCrKe35KXTLCB6mQx9QRY
xUr5TutyHyYFTDiNP6lH6s+oY0g32Qz6ZPm7BOBKtVW/Otodq2gEoSjpPnGD8bFs
2053HsmsvvN32N4wDAr4Dn7VNqkXGOT3WSUXuNQZUM1gdjv0JyRvuk84oKkAfgmB
rEJ43vovkEwaecrk9vAjd7Kqo6kTt5nbCtAxj04w5Z+wLPggCN0bqoidM4zA1tlp
jx3nF6u8OZOkfMnffMYgAlRWFWQfEIuhecvwBBselsQOc+fpSgCK95oo5bBH0kOs
9eO/igUxbLBOoSKOKKjY8L/P07yzs3TCH+bHMrCu4Cd8ETJxSp7IcpHQc/slbzmn
wajZ0FUlvh/tEXQhuMq6iUUxEJ48g/a1ZE1RvjqUUFX6hxBBfbvQD0/gcEftD08g
TtkM1FhCA/Pl/qUdBAkN996XXLWnm7zKCBVFsbc8px0et9vOos0Rk1jCdgH23HJC
7p7GBrtWYPeCqMACvET9RjlKHH0mkHY/LtfSkZ/GiMj1DILnxmkoiZCnzl7vFNay
FibZ9ZtKHTMYPkvhopegeyNIijI1sgtb7FanxMJI1oNrjvz5SCC9Uj60yEkFxHts
3LPQ/edlvLA1Iv4jMoJqUqEyCZKLPzuEAtDvqfzWq10OPmP+gI10Fm+A4Dd9z4vB
AUyh9+WqNmiZ6hrZEgQE37hlHhWzNfomFzyv0+wHKt4Gg2KZXFHOAUDVc9eA4Q1p
2HXCCIS2nhjH2hh4sQ+lQCN5OX+uQgYFCrmn137kuELjUDrsGEIRJ9uPcPT0bB5M
qv9NLKGvM50R2j8wGaFhNjLIIviegiXcZNYmLPwyw6CAGZwaH5zNIMM5nkTlWZWY
DkDb3g7jSsPOh+gUWTnXVc19vDyPwrKdT1WPpHHwT4Z5Fz94TRl3Yts+ndjKMinT
T/pxPH9lyyMKXFyROP9W24HnMVICAVbR6W7riKzPq9i5ROZGSQ7wOiBkjXVctP+U
56CTTI0O9HxoTiNEptZQXqT8W052pYw1cL2RzZt4noqroBJYoit7a1xIE6MLb59o
HaWPSvXuwXbVh5RPVTC+/wOtUPKYb2IWh9Dle1UB9Dpq6B4TlSNyqi60+1JtHNd5
3zYmRlH6x3jRBlP1vxY9lg+QvQV8geeXEQW6GSnegoercp3drGG30WSp9Ryk173q
M3SXTxHL8MDWwyH/29mFMD39W+ggukgA1i4m0Xbm7EIEMH6ghIhAfJYqL7nf3jEB
f5cBtso0MJ721XaF2zXjoqgCKIyHjhmHLwZ2kww5boMiw+hgLxqNigaKVyRyEn1H
momulJIyoUm6LUFtRRNcdITnLidPufgi1qCYqYQCK4Q5KcPirIBtvXASaJp3c2cE
DC5yehMu1n/X7hJTa1/IN17iFNjP3Qyc5p59HENcAbZ4FXFaiTdZ9Ss2YTd3QDqb
4ve7OPxdomg7n6SVWy7zlyfx4kL5CJX0MU9TknDe7UcLDaEUG63eEyzB/QldkTSY
AuMF3feWXZXSuYLtMdwet8CD8Yh/hfoo5LjJtdA3flJ3vNCA47xfrjAXh6lxFH0o
ub/lRlsqf13kpvCRs+acHg/uTYM6m8k/uLmAxR5M1dEi9RGJ3Nap9OUASJogwRzS
oIKl9et8f7EPVWvLEltGWdB8OV/Id0mkkyeBPiFFnSzJBXnb10OGv6YfTbwwDexO
YZ9B4TI4F4NujfXP8NHPCN7RBF6g7EjZAff6Cg8Go43wCPOmKqiC8dLFVNd8Sze3
OC3UFYmhawdYoVigfOADSO5tx44VPjF+P/cxU2okcxpW0AUvoqNqnVzAayzZ/IaJ
tCcCSnXs5pq2W2/dQq4sCI/nleba/IBUh5ZUujJJbscf/FXjlaG7HZ1GYugwGrL3
VWvfAMhPLl7n48NnUwy/qUf6c3R+2MKYFnOVQv5OzkPmXFCPzpKZWhJS+s1G4/eD
2n5LuY2nSN2NwfcH4EbyrPWqelnIR/6/T+wKzIe+NpzkpjnWJEGU87rz62L76r0j
xa9yM4DAlVmLgOziwNgPqeiw2MyBRltzGtLF2m8ZrRSbtg2Yxs3HusLztQ2tAA81
LsPOZH8BpoN/930lHG1uJJiaIOX4j7a/1YZVMH77ebAZnnC8/ki+Idi3Vhw3paeS
cAYYH6cT2hRuHMSmE2dHsXFJsPMOaPAS/qm7LXy9/+dTtxio/MRWHWvcJeGykzkK
PXxsOl0mNCziRIi4TgyPstnHAscJxuuNB8zMmKJjLD9VVDy7fw2o11Uj+DA57nQ5
c/UZ8/iCpq7XiXNn9AIdn7RX8otXYLxRBx9yYN8ZSHvdWHeTDd+2aW1ANtjxzZnc
bD6W3bgvYIlDVf98NVIGx1C0c0S9WVpRMyo+jQWNYrF3RdGIsJwsjlKD4RSIBsHt
8bZFEI4wK7bZAFwd8A40cBz+ZCVF+b8/91mhWpgz5UEFXcwFUFa53aT5gexWZGlN
y9ED43yb3HMvTtElACF0Auh5HloYom2UknMPnZ0PXGAc3gVskw7WXLXmeYlVl9Iz
069gGxM8ZZXvAUZqJqLCBHMUp/NIusx8nllf+l/qjdq5z2ZIsovu1f4sUPzJb8Bp
G9R0UIY853wxxDpDDG4OKtyG1ZCUFyZA9tYwiemtrLlAviWqGi+mLuMwN2IwohDz
BprQUPtIwQmCMEOU5mlBGR6ftwI+VSQphOrFS00jShpeeKUeIHUHjlxStO2Ex1Fr
pEr9/6Rl92mhT5MdaAZHTPwwrXf1AiE1Air3NPU2mLCztV9h4beg5fDPd+y4yk9F
T1WMYYnHfBijeVNt7CSSW6Zo27oS3EGdH6/AfdpOE8y0ZmgfcN2ETvEaH1aVpNB3
3sVmsDj9MEJrB2u3Btc0oUnvqxsYeMaiapW3j9HuDisMldDWHJ/3oWAN40g6zUxO
kuPvmF0Cs/FLtCUzTJ67B7BQF7nfXrOUc3hiEHEpKuwnFG3mmFk3ZKslg68N6Kqd
n70mPvvl5h2anP0304mPxw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bxk7N7EEf7tfuLeOSLmAz8A4mW1au/Ps7mpyCyQ3tWyMHC6ZJQxvvSbSGuL3djbc
O4aPQMFsxaCrodIIlejEhzXKeYeRdxccWcqUzNrAPWxUmxNIyeYIPb6jA8n3luRS
U5szZeqaT6v6172yOvHgv2Ims3O4ENdB1Ev/RWDqea1Eesy6JA5O2/REBVfNSzup
4me9pgOp3GZkJZbsboexWRcLO1D4EjnN+6Ofaurmn9rfOx8iBGWKtaPQWJG5hmOB
p2J+cDJujJ17C1kNNiAf65paXcbESxL89dOR7TMrZ/eKnYyHMWqB2tR35rI8Y20R
ln0TwEaUU+KvPsoedFatYw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 13088 )
`pragma protect data_block
zeLCQeTvDA2FMRCHeS2QNT3kwU3El4q66OL5lKL9WK+MtaRWgv3U2Coi/T3XYfMa
DJKUGr3Nll8opwX+9C8I7Xm754KLujUFUES9el6ZyA6WuEdypN7a/W/D6jB8nM5j
48kdpycAm/5lHV1ZkzsC/raXUVFzjIq0qktHfwpZwmZgIp+X3CxBR0tTb1qZVrLJ
yIz62vYmEOfiaX6PGy43cmzNjPA8E1QlodTvPglx7zFeW4JSP0iicEO1g+OLn5dq
aboV8LlxL54pwfwfF5waeX/L/Xoa8V4e07oOTNpVTaxW00K8zGpL3YuGqyQAkTJS
XkuykDUt8foJ46MadQCUsL5/CQTVTYRNNMzg5/bqusynpxkScEibObEa7WolNjcq
RelKzSmE650jkY2q9Z934LucT83mZlky/Sy2dPUT5kgH//RKJ3MrJ1WKtk0nXSqB
7VlFfFHjWrBvkTuuvTt+WPy4k2UkuJ8UWCpdGI9v1YRLadcrEmElbmpNbqY0FxYE
prUN/MivphaNMcthUoDSWvQANhaYmmuwMQsUv/6CqEJKaaCX1l9z2wlHiHKrAAHn
Ei7Z4p5Mor0qpgymJ+aiE7pGQOFQvr4e7DJ2Hr1CLNX8wmhNuqnFRHgxfDTUbP1D
hf1pV6pAOzjaxw6bjW6X+WuXts5TBylOJpK6Yn2uAiaq3E413R+4EY32HMT0RpDJ
1xaw/7XWsUNsovLLPxnLlVoLua0ibSLTVEwkCbbxxI3b5P1QJm0frp9LvcoE8Wm4
niCwp7ScQBrnYsM6y+8KHyZBFOsKbmZsu4axWWyjsfEI2zL33Hb01RXWnBt2fUmH
CFthz4R/5AymDJWuwTkz7IDhK1CRyfS/XqFaIWAfWdQXVwnuRI8r8bsI8FB4Iy/B
cCyMO69QktGv7wyBvSIQKB5bXmdAEWaBcZRC+8fkv5QVUTdx9D/ojva5YqoStGvd
z2ahA5hJxg06FybRqUJrf19v1XphTAGyb1FoMktB0iAeYajv5ULNa/pCX0qKecKX
qbA/leP4NIlwMe0m8lQt77kkTT16Lb5rE6BAaVSgbm7O2N4LcA/rkWVlQaYy7LdX
Recbwtdg8c1lHHod9NYxNGNEuR4wCHmcatI0zbt+3CzXkpfr5J0ifNKk3yPjv6RZ
dTa0rpYGHOpg1Apcs4sqmlNlypn2WVPfiw2RP9u4qT7DqHNZakh88CrINLWK+TGR
Jv4Rg3tQZ4gaIBTGlNPNAPtW09I2c05Z8Q17WUvJbDqtFUUL4a7U0EouRrWpBi1Q
c/AjDJyP6yvyGBtxqZDqJDdg8TDZxJulX0kKjHcRnlo5MSu4nxhrE8S/ob5rdL6I
MuBxo0QNfdXnwFFl+Tki1rjWfpshwKqtNpv+gOSV7XcjEKLc0JDJGTflD13NR228
dLdZkQFY7AQ/Y0Bocw9Hef8SQ9KUiZLPMY3K/kBRqa+jHB5XrMJ6W84RZT+MjdPs
QfeXelFcLqMzKqwMTeYVyBQHzCHv+bhGrcC+sTOdavNAZKSlpIoLeLLKbs6UBmMA
iXXNdDz87hUdCL/Tq21lxKm6TO5dQCGLATC6L3MwjgX1D2c3Z3GbIsYqtOfizjHP
MIUCRoII0+nKauQ/gXsod6tEmH5vbo+mpzvk8F6FwiR18D+2jq+7+2Cyv9aiiwic
VZryjSerSytrCKgJ5gfHWf2HeFIOR93QIgR9dXn4C492RFOYfiwLcnvWw57+sKQz
aOnqUyWPpW8EidaZ4khM5R6oaF51HkVkpebMsE1ozZpAEDwwxcixOAQWwfVBGM4w
2SEwFPPJ4TPWOulcmdn9NDmWS9DJjyQ8GLPDPmzG2/Um4s7yvTpf2e2q7HQnbAA6
VEZ0i5Bm6eFw1rfFbj6Dx08aJ01cJ/w/ncRUrIIaeZ7kCJ4gy+WPNjVSYABbUEWB
ZtG3XgXH16IU1Qq/WrIeqeMgJN7Ln6uEWNVK/uGFDxLLubWX0rNnWbOFXZ8pQffd
43ZtbMI8EG/3ExSVi16WWtokusJXVgSH/S3cN1CaYD0vUogFLZ5Jl1OMHa7tgyt/
H5LISGQm2ULI/NYcRiNWNXxi4Ansc97iZ1S8QXb9t14qvuHlOXrArl1Ngz0GsJuj
srSXI6299nWFAtWVqqWM+/cy2rZcNMmiX5zwC8Oi1990OoYXdE4TvoQCVlby2385
lNCld6lZzt91JvFSRBBHG+hueWktBTCTydnFdU6lUT74UjvDImnNHLqxunk2rXOc
glvn6xBA5xWMD+OIrVtcQ2fomH7KWlxCPBZI5ok9GD5wLVDItCgTIS5ekYcW1x1N
aM9HbOoEAZ02Ho16upxKAG0Us5vYj8jKbT0re9M9atVZMlms6eLsjsrO0rasOuYF
QJlYYVDA4lW8oxD86WW/T0CNWzzZhi2aKgeao6LNkDGbe7J/FuwSLCzmNm/5PlpU
LMwB4RTMvCat2Wbk/Utz1ZKyVs4Tt/2TwryiZ5JW1eG72FGp/qNaGXzXlUiZUPqd
qosV4HYJVtqpxZZ48mNUugWJFYb3M1OLD6nphN0W4wOMQWopUE6acIuBBNCdgke1
V237I2gc0LchMsSenC66okcGflAN1G0jNqff3n1FxWtFlM4Dayom0XE7CnfYyvgJ
UxwjxXe3fKNtvO7a1/c72rGigIT72LU1FzOn95OWNQI3fuPOj7flA6avz4mwqj6i
buTpSNepYhZXVWcYV8PEJho0GcSXMdvpXilmcMgwKnd6V9+ZY4pCN6YfeIa3j3Xv
RL5ZbAQPV89lvvX/fCZGK9RLQpkr6IZYLDSLAEFFQxSauPQLoYAX6K8KjqymS4w6
x+84xnSJ9647qNYBSg3+657E+BHhrf+rl3CX9gghFeM/Qt9iDEAalBaq7v98tR8V
5DSFfqWZzkYTiMb6sCaDLJw3s4NvDnbQGssoH3+0ZER/DbM/ttffbzabNgMe2d0Y
ztmEvDn8vnyXJXl8d/KG5J4dFLgDhnI9UNplmEDyZp6BtnqFhykfbtFjNvRcyRPN
oj7M7axQAscYIdDLzsFXOoFbxsU1jeM3xcmDJcXafiMD6lPkm4OE0MoqpYVGWY3A
mo5wFilLzSzw0YzciAWZ/PPwVbG44JNUGz/bgmGUaUBoIOpKwqfWYNNenHpgYBA+
AcX65Oglh8mP3fQgL1/vwVRYehWw7dmLOsmy0dIsJk4WGW1KyWf/HyW+JKZniy2z
PhYcHaCFpgZwVJ+EJCTvkR/uHZga+NWWDEhr1UluNz6E+0Pn8FR5HhzCLcZUJr5E
6zJhK04r9Pdfv0mZ5tIFx5YMbUPHQI3Y0sGYfh0TTiEzVMO0Xj9NeZ/FB7RoilKQ
DNwQDywRW91Q0QRiOjwB260aX/Sz0ktAwqIYeeSBD1l6zn40apDmmy1JomIQulO/
FuCsrd2v7D2Ccffg1aAI7rk9NSrfMN8XFkDSVcA6qi5MJZ3UKXzXIZvxITS3bpbP
SgpAwPjmQby4iUOYjEr6om/7xJ3W8D4rptp98J9cKnKizE6PaVKZhdUxAVtCB27h
UQde8wxEiwy9LtMLUaqmq7uK/eMIir79hm48Ks6OvyLmAaAmuFpx54kteTZlMlyT
P9oZdzod3WYBXgwcs+g9l6P0SX77OIvuDU/Hb1MxVO4blkQmrx7JV3sAQnIOjDDT
IpQsZADJ1qM+5dK2n3EOQK2VdvHThJ5UFo3bi9XGwjUF46CnvJ3/qWMCR3/Uw03j
Ms+EZwI6uciwFxpZDJwyBe9Mpg9MYQAL+NI9LTsFckuLKuX5/0nRNxR7a6EvrCJU
cuSM+DfNoyxl6IvwW0LOgLQOW37C/QGFHpjccjHvNVtxeO4cjeg2v2YSQNP+VOqB
SwivZ2glMuC5tk2o1b1hpGZ9IcpN6nm/y5R0necIbifbxSpy0e+N4mIN5KmGws/L
9iaApnIH991mHC6qns1sYe7xlv00WuVXeB1XEhsErmN9ZtMR1kHQc2bLRAGxOSZy
BPboWw50m742q7iSCfnSHyKvr8nz6jxzH0C+OI6F81FR6fZpEqG+2pUMzRgBLbSw
DwctUH4ITJECyMgIi87ncHCaHYmBBskDItUn65wp03gkjFzVe+/3lov/qi3UHJDt
jpVN7V0K4eOxJSJC537tWkzeGXiOI1Qq7uBhH1c+0HfW5yh3w5aXshDzs+sDwiDE
q3GR6TzBcsAcZiayvtCxW+mCWHidsD8VEpLsV3vlGZTRu/P66F1UZOEsu4lj8uA0
VXTXHGvA/xM04av4mMQPz8/hag8zm0E4duEVUaLQU6a4q3trR/S+kHPrN1GxXjsp
sJcG15pNqTvwPAttwO12aL2QPVg9wU0BNKtHdrBIwddrNhYyBmBlTke59ggSJ4iv
jiHeXXr6sgnQTyYNi3LI6FAlKfW1kCb15FyPvMzoXANtBQots7AHd35vNL3rUKv1
/CQQl95KxtHdeMgBZZLUUwDDvdKUUDtikjITrUECHZgO6if6vZY9mt2pAHCb0lph
9hTFpjSjT7dcY8U5W/Ls3zpsZcdjyzZ5ff2SbD8Gtkwll5j9wvDZb0ViqoK3VAbD
2HOoJwV7/RVgT0kEfebxYNKDvg+CHuCX31vllTCOIRKnLER+683KIBT/XX70H7wK
M3TIA/L7b/uTiqtyWW6e1OHaP7SkCfJ4m1Ca9khLo9/N4vOSnijv9OuhUjA629x0
9XQ5aSRv9bXm3/utDF4q903wgfxB+E6J286BNjjxWhFUvPlZLnOGXWPNfbPJHydn
FsGqTNv5VsAUNvt9iNB2yED2+mS2/6SoxKcZHUlnQwWOD+emjZdCfl5fku+6vbA6
l00cCNVk+2x2bMlBSFweeExBZ6rA4pkEnxYvCEQOBO2QmJCaGkQcD6rY8mcij6Vx
RCOu0MiJpIblQxLNX97pftojtrPKhkTtvxcXA+wNW+icj0Pjce3x+Gx+YDw6Lz33
KP/cXD+fnKzrxYRsEBO2Og9t8Ts7+8803YjwUa14qJPOFtP73JDsQn/Scc+bbgfk
AfuqG+nla9lZ6qQHSGlKTqW0LFh4XvD/zVj7aFtC3c5nkcf4iSjGB9K7JCukuo0k
kUZyaJSUqxjJAyf02A3c0gi+sfF27xDEb1a+gdr6DGqKlsJXDO/95nPoEo0uUHrj
j+U1H9vpj287VicXUnUiRiPNC532D15lM3ioI5UP5GPpOPfudK1HO51X3igd8CtR
fk+9Nlvp7XMx0dQqEQEx3XbE8bN/k8YwrWSdd7y2CXq6HKk5ncyvc933iitwOaRq
2Oil/PjrqKa3CmGmxpYdpr04phou2oYpiytVSi9OvG7XRKPEKb14sf2GqGjd/qoq
GI6KVWUwGPHpOVU6b9zkSFAGnbf6ID1h9zBGIJ5eWlzAWERoiuRvmQjpusfl5KCt
zhs0AUUj5tvDGKYVOnuQTT1BnyLlt4HT4UsGrI3LQ0AtsoqCbxDaoA2yk8vnZKGz
uzFNuzRr3E1k9u8EGugjCA7FdMQKPWCmuBezcG3H+C4om/VWQViEW4eVuLVpEtsz
6c6XxTniRasa8dEDib3b/+1VP5pz3hl7SiHxrNyBpl9cu8eyaAc8IpHICv8ZwMO+
7H6HMgY4CMGlTObOf+Jf8JrfEKPrvOvIz6DRg/ZEqoN/Vmr4+bNiSAyuRBE2JYLL
wa6x8eR8+/F/5Iqd/0w1JsltheJXbllY+UTeLTS82fhEtY/W004g3cCbBtfcgeIZ
unV4dg+wsEPTY6/aznaySACwVrGDzHofyTXuPx79MMmadgpb5kV3DWyWweJMCPMx
Y44uUhxVcoQSssTIrOiuwQZXKSIELbEYUkZEDOT0K+tGAxR/aMum/abSHsfw2pqW
gE7biU9nyntV7iy+1g2aM3skgxW4RyG/p0g2HlGWzG3P730OGQJbR2JyV+ezvKXO
1YbX0w96kv48A29Z5rVpdY3iGrZLHc5gScfguJOClu9EayXzOVZ47aHs8baLZOcj
sxE2eZNUlCDIjnJvAjjl1txppt8eU+/OHaHNyp6L4X01midBr1mVSYp9qTBhrdQy
7gPbDhwz6Z7N70PWQLXPv0pJ5p7hA4pQWejHYwWiWF+7D7Rwphdi2vawCivkiWi4
Dswcqq37ebjblylu8YfnhEBzYw/3BqOCsyVCsdoYdkQv0N72AaKcxRlGgsc+nFKk
S/bTzo6SH6oXbzlBvH46emPjAdPMN6pixcDFsBC8qHIvCNde5HGPJvqRiZIq9IGs
j9ZS+qwllh51biktZiv1GTr3++fIUV6GwGBcDM+MdKSIvR+Lq67mLxfBEXBo1iqo
GeloAWqQStWt4jYV4ZnRA7WGgxePypPBKcl57GXRAYvpxoA1G0rNvchBVq6nLR48
LJCTZvOmwrcOGujcYCc+PfasQlEcCFsRkno1xYLWJZTVcnAbq/L3OM3gIgopEtFi
ZxlJ5RH3ldzZG1xpOACUGIhm6wfeZmAd8xCNj4nhy00ATZ2qjCczgSBvnAi0RD+m
ATxi/4a8MuXjbDpyUopkOu4CIg3WYsT+h7wWUjVXnUxY0HF4v7XSiZjtDOgDsb9o
QMK4OESnpAE3M9ZUeHHXCJi5kp1KdnIpS/JHnV3OyWPc+s/APt47YX+5ajrHVrhV
nYeqmq821qTTyzMrmmym1napbaKwtVgHVMsY+65OSHErY/wnX1O4SjzCAlvSGjYz
HfavSOgjQIz/+RACMObac9SnmKgh+ATLjeT3Z4sJb9APXBS9VCILLzKmwhQGmGEp
SDEbAlVMNllysBKqSqQOlTEurZH84otNi/3wyEtD+ddAGx5sBwXYBI1Gb1obJyg1
0qfvNH3CZwTypVSbuWayTCDNczf5OIpZ32Oi7OG8O/sT0/qRbYYm+MrCtusDvmzI
YDotk4ch+C9dXLO7TMxztH5gjH6vA7eTLF3X/azT1FTqeqSpzq7YrLQ7bcGLV2NY
HZSfOPuf7/mmS2EOb4/dJqCaSWp7Fwf9R9HYYRltcZkbNY6/s3eALcQAhrNcUcCt
LfUMRexiqVuHDWGBXdaxVvhCl2aiZq7jt6HjuvqlhR1O6pZAc8PXEOfx1uaNzmRm
+HDFwvGPXEYcoUomkghIiIYKX5tS8ecAJzQmmJmKCDCxOx6POsQHqpo7Hz9TTcZU
tCTHHzftpou3stVrNzh64BN9RJmnrL8+aUf03XpSZF54jZkOdPGVGwxe3UpXU97S
S0E6pyANaxXyX5YxVmDm8jLyb0eZcuDJN4kKKXH9qV7L5w3I3ZVn9UMtn3bJjG4b
gtiWwpM6KVY5MW7bWz173rfUYroXUZGMwCz9Jc817JGn+tiYiCao56ZcG8OoHhgr
WlElct9f2Njco7ZKQFR4LThUHUz0AB9Mx7mp3p7b2huoWxeZxLx+UknwbFX/XtIF
u8yfKp7PMZvtUmZe+Hf3iE6E97IPc36DfDmeoNTLmvzVIstnHt9vCcnu90nNsoYl
XgZrTyR5uwvkDonJTsYEXGad0VhkmlFERT97l+5c2N5ho5PfdnTTxwDvnWmJFejI
tAKpVupE+c72O+XgDIjqiXRyZ5ou6Gg2uW5jy0Jf8yHo7N0IBVJKB0TpvtGkAAN4
L8vRVhU93lgFuV7Zv75YQP4OfFOvDz2IhRHvGSbHsr2Bkl8Qe6zz+03oJNgk6EXR
vljDqYDYydBIOXTp9ru8l7LNlFkmnIbETlWGUaLRF2NxL1nMBw0zDzEqyNYetkW6
dEilmTXOM0KE37pcuAORCG8rY8jNuqnLwdAHy9+52iZ1tf9B18rgzFfB05yKQdxn
SKP3UXmBuaMbPHeY7CQPcOGpT+eXKjfxZHQQLimMt2lhRtrecQ1oczDq1SbxOwI+
kaoVsCOEXpf7/pPyZxUtIj23rAitNg+6NkPfWH8cth2Wg80L1lhethrq8LhItwtK
5T8I3bg/0ophaesnXAeIBdLYS4B5xHf4XGm9a5m0FCaY9JZW8ltLnPVuXfoB9G7p
rquUE4COD0eEAfhmySKfib1+u2Pxl8O35v4F+vjPQ/way/m6AanSdOf5p9L2uAJq
L5xYd7SkjyhTZeZT9nQLn4M52utu7ZGqjmpYvxTwyQvtHMMpOkSzDXCligEXqcgO
2K/ju03dCzp+yia+enf5QwxdL3RYN1lQNRBTpOUPc4OU9azrba2AxlHY/nKVXnyi
0vj92qSbTsExlGYTUp5bjKNhv9uzIPQLv6PLln3CpKHevIw3Jcgk3Y4RQ2cqILKK
ZFV2GEfzKOByzWzHTPpC7Kg79pRA7YKOKSXd+opBrdPzK9dAae+D2UGljgHg7xzF
p6odH5kc5eIVG3V0tEvUdHJqAAZ1lmH6wDR+UXPH5zqT0cDSuvnAsxosW2Az46wk
LeTAtZ9xm3Fa0of1yj80OhbZBuonm8dfYB726NBjV1unXW7Y1h3cZsdlqD689k3x
bOBlig5kSfjn2cxebw5DO2vLXnXlWx4QvecSt+eDCF0NHvWHm4HhC8a/8DBheM7o
MSJwwSJ3JKYHK22qcxuHuENETrcTS4LJ+wTkSCN92JvYCeNevupSL83Pf7nOBMsG
SFzJPf0DaE09wXskGue4grni6A8IqSS1K7kPZEoXhNaJi/1cq/Z4hYrkZCK/iNG8
nZ22c9kWZQDe/y00bnvij6Cc8F+RF95SZDnM8hPgdi5nh60OJZ4pueesfS6N1xgk
rwW8gEsIj2AueD70FFZpOEcSOgnAbhwPhB1VMQHM/Cyai3R5qVR4rC1NdiYvj/hO
CtlsVy3pXe+uTbn7WpJceUraJoUMxCUV1J4C4WQy+6Ronlw6QyZKM06MNBi5skKn
78wNhex4QF0LDeRpx8Q/8stkt/v5pgj7kpWOiEe6Jqt4v4dRq3Cc9buUGefMqSbQ
fW1WnohCWbOymF7GTPyD/HjVUEZoZxT3Uc5mzJFWacCM2NtmdTDxGAAlEW/CQxZU
fpUySyupHQyo5GsUkf1iIh1riNrKBVzzSuW6MXEgDFA8ljGntwuA2CwryIVYkiAa
/yn2f2TPeskDuPQ6yd+4T/imK5OXk8Z/rROq23tqxzg4NdJ/8n5FRIPhHl814x1b
mrKduScYrUYJbeM3YwZQAUVxfYS+E2nZSjE/mxRX31ZhcDRaIin52I4g2NpE9XJs
OLUNns1e/wbDyCTzfjuX4aw9Bn+UrfDTPjy7dX2rXZJpO52JkSxGJCgWPAXJeP0O
uKcH80NTpx/xI79u964tUQKHs3DwI/X+UwdUuC+GASqQWWk8VtNYYcqMfhQbpsud
jEf9fx6iF4xGV3AcWeAkl0ffCMrVZKRAqTO9LvwrRz4OO+DMh3AmUibrS2/xRtTg
AOwxYgIENNDBqitS1SVu4yFAYsS+s+SylafWAGDPq1X3W7Rx+f5bsZvNuuSoG2pd
k/Dk94poCZe5v7P8OD2B9JamMOu+o6FRqBejvVdrkMPFmubv9cx55CpEmTLpxiq+
nyjR3+WN6PNBetBX9I0H6kYVp3qJvsKPO6V+R0nf+A7alL5eKRQ5B5MvDodTfc5Z
dRQh5y7RF5cHokJ7IlvX1yCJSn4Iydo1ztEWe1pL7H2WBb7jsiXsfw2+E+ZoREvr
siqLleO72snjxXuyDfqv0lMoz0rNq6grJ6xTgfSSDYlXZ5luaTIJJXchFC9elWog
II3O9gYxz/NjfQxiflvXkv5CZpyJ+TpyOJD0E43nttyxy4hXpOKuNpfVnFN1ULD5
jzGz0B6K/pXzT/aNWKJjUB5EZZ9z5WDQmPS1Bql0E4e3SrL7tdSM1EQooYnGKyqb
Y4rPkgA4IXrw69Tx6apRTCtxiK4Ue/scz4dK0txHu+D15+Eypbed9BhQok/K25K/
13lPHOTGcoPRfLTQeabv94EEU0TKczUs8ZQVBnmHsnR53N7Tw9qWAEgVD2NIhHl0
t6UXm/I4FcKivMaiWtieSrj8dCdJQO9SeBvVSMHy5V3Nfz8nMW1emC1/5GoX/t8S
Em+vhfLNc0SEZEdoID68LXIdirW83OqRhw628QYzOZzxguPmjOkFl4KGk4sZJpRS
t+5+xkr2DoqxlqusMFyMjBoSuqXMQ12xQFmkpX0iqXpQ7pqZQm34K72P0A0Kos3K
KgKDdkEXSbcvjVDMA4rp+CjSWZ6NxE2u4Hoy7r9O7fMhV/n++kdXeKwSHc0fk3+n
BP4YVx9ixNMypZM9qch3ruky6XM4EbSVtmT5vu6/9ivImInEUAEHKCYlSe58AIJO
6Thi8IzlSQQAOo7SuwhBgxFMd3Bf9ecb//EsoC8mUTWRn3KCxM0aYzPcnVFoRVgQ
Eznhin7aHdrWOEoRUgGcu/7wOswKwtH+oAj1upeljvKH8kmRW9P1NiarBXLLTH1b
/DOI4Kh7AOxrOtGkGTQRRWsfPzv3Z2XmShy/QIfCBQitlUGxN+IbvtSGdZDdcWqL
3MSigNY4VnNwTl6IP91UVNsIScPGUCBelj96MPDDoGO9tXMHPPsI6PkSfhOKDFag
Zb0VMkYc1Yr5UpHpFBrZrPJAq/U0CnBZoJkrGXObTYSbUN1la5ICTjHyj+ya+VaA
uNmtLFiOYZbceMtOyeeTEL21bcqQDo3gZrDk0UDs0BP/Dk5VxaJ2gJz6f8ZPNk00
R0lnsV7+vbzdXEy7HUGIJWCfwOJOJQb4t+fm4jkYrsEuFjp/Ou9DXTpcER+fSqyw
4O2j0ghOnfpw1fEJCo/lbl3jFNExJ1t4HwgZLfXza8dx+qwJ2LwBbbnIfEqH/41l
ruYQgpBvNIk7CCYPkedxnu3zFYSrKxKD726uEfzLYO83kqP8trlM4lfpn2igGXOS
WcKpmmx7r8DcPXcuL2TW7nJTSdU6j1I5q5UN+9P+18lpnfzErsfhsB9R6E4VU0en
hKTlIFqfr08ysMWdAhzhXBLFqctyI8bwChpuykU4jrnEwyV1VznQzCpDJHzanHts
0LcYkqSEvMnDWk6rufJFkJdcMJtcEYZkcnzqM2VCg6PHyXZGmG3D07d0w8K/Qx2l
EzRYqqXHLwDrXKBMxovaiSOl4aHHx0Y4fYJFaqoQOsHRBxkBMKiR4kSufaudQauK
uenD8ncNFnF8QT4u9pfpJmiiwWx6DbV66g+BkF427PcoEx7Yc7zVbv2mUdm6AcAf
oJslwEZf+zpklTriCIcppkZd7whYW9lLYAJjQyALqzyVBdrwC/oPSMBgpahgWeQ5
TsT5oVuj5fYkYJ1v24z5BtvlrEu+avIE5wfnW0tRw1X/kJq6kTXJzd19HtTuSnGj
Y0iQep2AmX2j+DiVI9drPxTDtuCh9wc4QR79tMuMWebka1X0quFUf6BlVXESexlE
zXHxysysrIZ7mDAD2S/EfV74+PEY5DGSRxlvPOWJouiVtMUzhqrooAL4++yAl2+V
fvoEYJGSEdqJ1AkTDyDPyhSqKHeeqVYr04htomLGVo7oR/PNDSsU65e/8gqs52rE
zP0P5D+u9Gp8F1R4B/5Q0TQRAfCAm0Mc2WoPFVpUMqKF7jiLxtxxQ60r2h2+JvrM
OXEB935jA9MP7mTQVZ5F6pr5tP/oOoYpkbs+rhCnQlafNl0PpAsFf8roljtW9jOf
x5WdiGjDSswhfd9vWSxkw+2HQaRWHfBM572tuOjmnaI753oL8a1yS/qEREmO1uPL
ld9zFPIOQzQ6YdZ+LvsSnLbTMzdBvObKGzhIg4wHquAqKC6B0KB+nJvmb3wBJ0SL
iXAwx8qeXhiDZXehOqbU7t2cwl/ULyqfl5LxfuRExsVjMjWoKBWb4wQYVR60qoV0
O7n2SAs1mrDbcH9Y8ldRRFn5uDNDEjrwaC7lihzQ7qoiG3fGAYT73KXObxYVH9F5
BfLJpFOiF/Ec9/GMa00Vc3/bcjxWGMueTuxL1LFO9Xg30O1izt8PIrHgwHRutyI2
izr+u09gmJp9eM9lIIG4MeHt8VJ3oZ1Ewths7KOGvyM+nXSyF9tAnh6kK09wag29
sQGUqxZlxk+A3hisQL83Mzt/pmeha9Pj6Is7GO7QZHh4Eqj3oD8gYfPC2aytqBQu
XY+k3slgSoi2QFc+QoO+0vIN70HM3zu361CrnzP/a2y04JveYEJhPJgpKOqVlJvq
VnO7QF4Xppf91K+SHwtMLKE5082zB7fEWKwz4AT9VWxXA/XqpQPBaUDnGIZQdfLj
o5o1zRSUukEmSSVtX0xcDC0IQQMGsQkGAspNke3ZLRcIa7VY91K7QJgk71JYblei
6IAUoIQQN/CC6blgEcShbPe0zMGnT3f2ecfN3bHRzDMiM5957YMZJsXu1M37B1Zy
D7KBTF/oT7Kh38BpPNgYxYjzfPPOMg15xPdc33SPb1fC+ZiyMi0eUzXVuQztzbuf
1I3L9HoF8hC8JIPZfrWytdl0Pjxp7dhYRx+pex+Gzh+UPWckkLzRKstyurjw13UY
ZmImbxLpdULNhLHunb5RS7KOK65eJUZOwnmsAxtevWalzOSrQmex1VlsFOl3bUGH
MFWLKaYWslEfDCbJfDToUJvAwU+pwf/PjcTgG/SxMJaXV74kWvVpYI1ntPU7Lqob
uE7Ef8qexI6OjnB8yMsXmzLyuOtjER6lCofcSP7QtQmIFToLxtqfZjaQkFCiGoW/
39BL23BQhXTuf/wAU3m1el1qN08TrcbcPiTsx08y3gSC8zK4GNRJ/D+vV5h1ezgW
U8X/5UpFM/JG2dkSb/kyMgVX59YCFrDOsDajEcBtSj6hhqcRwmQEXDM3mNuiu2MX
55E5E+pU3NfiuNZp3ty3RBC4tL7OwVjFQfE3A4ESIVg3fvERh1UHNJuGJRq8Y3GR
mbPPzz/kpmJvwqh/bQV4wLk5Ly0MWAd/hHa8GoGPnQUaIVvF5MUhoH8eeiHF9Cug
yC1hqDioL93SEA4qjzWlNbm370v+SwnQhPc3rZSpMtbvIWtXzOGJ7JoxgZrPRkow
Rq7txKPMAiNLHeguf/ViWMRJHZoW+aPD1kUA7+FG9S89TuGM0xbzLkWAo5OLKMj+
+gcMHJn0V/KPhYpE0XGEJRkSpD3qdo7My9scYsBNqSLC+TcR/6uppE0Ezb12mXNU
ycPGKA9F9HQsXc4jYvZYlMDxEkR99e/r7EdsZN6KeCIcesdLDfqTob198If2tL3U
ahzIIGWmL2q9SOEf0/b2pPTcWYk3wFUVkJfswKF5qBVmZoqklqAWFWU7znOe6eRV
R1wj7qTcU28oHeOP830Voo4Qg0K1bsDYCoiYCKuJilrcbOQJCJPjNRwLroU7k46z
CkXoIwLJ3aJVLnk8n6CV8CdzqL8doZWE30GkP335SkLTRtPzOXv3zZTG0+xZcMfe
5SzUYqjEui7FGebibQambs39fpQhcjgmp6uPLz+z3Hv1CJl1yHNk3hIuyflD0o26
fT4XUn9h1D/fw02G9QAW+2YXeJDtsUtKJtloDxWq8foZo7WFT5vS28Fz0bXWofMl
m2aIrwKwO/9yORTP9ghAcIUO7QU7Q4E8qAmejvBfzFY/mV4AIardK6jjPPPK2Ifu
4M7duXL6PP3/1j/Z+HeCQ02SzTBn/R+jY/pus5JlZGh+1QGILhIWMQK9leOH6e5k
ub8sAJb1/J9WHQZNxcJE+z5FBwGn5YAAvNKbHQDny53zUxVjeHa9wRFro5PRwuYV
fMfMF+NIG0WpALCEev91m65fvYIA0lflnNU+3Qh98uEQ/fTA5S16B4Qj3QY6iOal
dWHMT24bim3VrHv+6NoXVlLbs7tm0jByfmJAMO6xIDIDmqOpW2GUaCHS8Zn92Tgh
kIkQVNQereNkpLpXjMKRyqUS/g1Nlj11/NpC+ClmXNelnC3q1AuS674Y60oWHRe2
/6Aw0wSKe5zFZjkccl7kf61N+8LuaRACWMGg+HDNnPkaV9R6Z17vXPpwpsLoBVhs
Id2SjbrDq6s7h15IFV5FWJLlIaF50QAhKxf/mi/ikgcg0dIcg6zoASpbCy4i6Ysg
ChwPEXMktzdgq/iRA8V4zntVbhHxDgHC6/f9gYsmAfDkHkCIOjc3WoVmW/KQwZeg
9JFa/eBNVgTcg10o1QY0Ifubb8BRplw0thVQ88s95N8r6mmdN7tZ0Lq1jQDweMkJ
rvW29ujFSAtv1+VGPybU1STFuWu1G/vAivoMeDUitqPkKgwE2h/Lu6UBw1GiEKSo
imZNhRpC3Szs3Tt1NVU4gD9nAC6pJBhPvbVdo+QbVGadD4w4haCD4LuEAlv9KiP+
0TLdfLdpK8Lr7plVnH+5yhMIIX5j7leqQPGA6I6Wm/dxF3+nBDJ6ZWT5oeSmnjd1
KqtYyu/ryYREhJ5U4q/EBe471OIEei9lq7PaxumOq8stYFqdsmxbvKKoKaTjB6Iz
HKGsRxKKW/ij+33iiq1HG8mzcsGi3vluU7Jvb7iuflaDyvh8wWJMdoAKS2qw0EY4
qbJROT+Au91Dwv2VwJBXpKSZ+AHCrXsgyB4No123x4uQ92dt/cFILnQHVCWkISjb
9eid4t+lb6r2VZEdgSczBvTJWWUmUDrDDdlmfewCucHiPO+08KKUbnMk4/rtyiC7
4pQk8j2WzeR5HWZXw3QG509QBPRleNpcIByz84W73sgDbkmiHKtXHu5CF2rNGJFt
ieOGxEWgg9xGQ6ikfiIFwxPyyWwUZL1g5gJ16J1ci1RSVWb8aZESfJtoCCXSJgZf
VVuGt3qYKb3S4IgUdYa2ZcHO+/W5/SGk27T1VeFBz5ybH3M4IoEQ4Gaw+xhrBBR8
0JWpIJAZVXjHJ4P9gk9ToNg8jUulPAOkNoAIooPyV9yOEZQzrPuBqtwLZ8PJLhGn
4vUKeC0AMavdLpbOlvVEOlQaG5LAUEGwtGJ7YU6b3x7FF36hFWZfc37WW395uTN3
2cERAvSFzz0vXG17OND2E/snbWmbVhb+DsO0wAPuxPpkEM6YGeX6425918x0p2B5
QlUe9hUvemtDJAhweFEMR+QX4re27CjEBlFFZmmJp3bNcfwTcAd/BAoy03a6jfxz
s+GLzHshd6yedvSw1iHYDbZuulkVEgSKS5mDwjIpV5b8OGLMV9MzXWcKCIclb11L
Bq9aMq88FJMhwPmsIsmCrtFr80Eylk4OGht3I3O20s8CIq45Xs5myy2kVUptAxIi
FDyzxQeZUiIe8f38InUDf7my2R+3H0wTQYUSM2X5FaX8I6kPW5eVPNmJiYVJ9NK6
rf/HlAHEUmaNqy4et2KM3JsGmPGDL6IXFJ+ux31zWjAVLU9SxXmd9ksmQjYgv5Xt
SUaf9MFBtstzKoD8yVNeKx15bTptjI7/rnDAVo32AIbVFF9b/Q/5Pz9YaeFNsQOP
QCE1kPdWtr9haP2ywZrM3mECMs+v6kptJRVvhIc2irfgWT1X4Oh2I29c4jpb/W4q
s2TiK12gRUiCbSjvRjrHGmyZkI5qOXQLGzWrNUFxpbERyHdtEhJc4DdWx83Xq7i2
hAsFVKLtqXwGYmU6sIcM1pLaD0ICdMHqK3vTOo+k87tOD02iXcGvnYFqBePfxMzp
MKoLjZpqHCTFH1Uw314RccRv/BRHAUdnssQ8Xl0IUujuSRe4i6iHdSlCV/kAP3QJ
/WUfnfpPTBaT7B226DMCUT87EPmDEO7+r/VWLdQ7J7JF9TmeyCfeZfF5HJLuXNvQ
Vbcu4qUa6istL31asIzyp0yTP2DmkTt+7Gaz2a5DJUOEIFT8L5M3dEj7GnzFRxAA
Xj0JsYts/l32z4EtMiAtYpeyh/FLob6VrAnglbsSwxl7KTGYMrlSOv2pRmyx+psu
D/fiziy0NXAC4tS+6tlJixPdQKXDMy6cajmP3ovc9x0/UpCxeS3zDqQKF+pm7kPQ
g171CQtm/XXiGYUFMQPRybByT1YghFwThMMhLpK4tU81UZHpveCFKZFc6TWXG71A
IQUaHElEXlksDVU+M0QbvhraoG1c0GzCF99+bJnWNeiiDU4262D6dcY9AP0bGXZn
rgeKiNittC8CswX9eqx+KCLBbKrjwN7VRclSipPF4yuHziJR+Xzs6/pbagYmboRZ
+yOH7pVSN4Sy8xL+o6yzb3QXcUnGuhLObEXyO+Qrya7pi8BJu4L01zkraUFWZ+QX
BP5qSOcp2w3KH286U8TM6Ybg7jnX3M9rVpCz450I7AX9cc2SVDWMS/XWhSkSpD1e
r6Zx3wn9ygarMIjElwnd2uutnpfU4rBOjp7fQ12M1wjX676BZj7/s7xlRkuvc3Ow
r0x8696608yvfvgI3PwGV5NI/bcU4Cv1Bjff9jP4fmMsuxVcpg+JXtp6mnFA1hDP
aFDWf02hlA1m/YOnPj9Oq0DecsYLNqaKR/aowYksyfKy8HhJ9mAaRVqNFIliphDU
yG4qs+bxdu7Q8LQHlK/+kwucfSBUWoBFAaegOW0oATLO+/PzOrgSaPqxck66XuZS
JGtXeWYzCFGEtgEsHFm/yUNVDyHq5qkQJ1hBzEjdDZ4qRySgtMlfBtU2VnehhC7H
iie4eti/ORpAcAPuU1qypQjK5zP1LjoRM3f71+Px8H51CRz64gEfeCgOH9FEeSAL
0PE4k6OXOnHd1WmtZYXLG4vpXVtnK2moq1AnaKBLb3GRb8z/Ov3z7FydAYvMWtaR
37B64+1FUpnEKI3h4Pkc+A4TO83z9luio7BYVAtLERPvRXVIL7btij66jGjS3oqU
uP8E4RvKj6kGHU69dZE9GcKOG8+q5TcZvSTyPqaumsCxMT7osiQnfmM3BUmkdjbc
47R2CITyZklcOYVQIrXFEccCixx6G95gMvxjydqBCrJG+EbleUF20YODvzxt3rqC
LMbuelAzi+ehFXj4YzUzkAtwW1Hbsc8yb5Y0voAKEy8UTgQxb+vcuS5/x5ou+TxV
Xv93xcObKZ+y5nrQ10yp4EwvlBw4oCFsHZaDUrLk5cE9A3XAfihPciJfVLGG8xcX
qX7vOdfq97CCp2P1RlcCwKi9qeBfvfOZI8/sDR/sDcz8Ph/0aoGIzzEJoVutU1jO
/OScjR1j1lVcrdQyeLZnRbRuzqTARp6XRrcLvGqhPFuezw7gDe7PP7TWpxSuXF/X
Mhy+WElsaDhqjP0mDL6XE1iQ1dQX55RUYyxM7VvuYUfrev5KfufJqibMtmJ6GdOZ
EXb0+GVG3z8C5GR5AWuyAd/K11maTq2UeQiEHkeZrirJhYUMNqzrg+wfw+/tv6rd
zeCfQPvR4pP8WwT+G9FUfEF7MHfWviob9QgVS29nVveBxNJroNfFnNeKXVB+Xv16
o82qLHnCAhuK1pHhnuiyrt1WIrFDJFubUeo5Vs5oz66vhgh+dQKJt31mlupXL3aY
RCfUKn+U40x3mTYXTNMTn9uRe6Z8rRzOuu3ihY1BAPPmdf64/43Rt49yE2h6cvm7
AhJIT/+lIkwVF2m8tJwPIHnw4oI8AgKT2CJkqUK67+bBKB7ZS80rk1iWMjkSQ1am
/VHIh6uJty/yCLjzXEn4KhSBtWktK2xYAVzbaXXyT+N5zn0s4wdqc2vuMspOvRZ/
Js2s4dTa/yb6Z4610agity1qRcRvk+N3xIFUWV8yZwA=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dOAxHclqvKBC0avYLJZMFcpsvmj7IJbCayq1wSy8YWXIUS8G7bF85c6ng9yorAGL
hCL3Q4w1rE39R/pB3rAB54xj+/4k1BiuUKswpueG/blpkgSPL+s2nlhc7Yja1nlk
e1s+lF4jvVxQe5xepvmYYD7RXN5OQHN2JBiKv+snNpviF5jqXhhqjgVAE2VN+320
PFgPmTCXfLXy7Y2ARrTl8vwddoLX1lWZkvlgBUkyvwcUOcMNRGKXpM7ZgCXUkIjJ
Mql44TMFK9rpHFQBsMlwHg3/f1AewDhIvVToYnmoNXocRGRmS/GA3KbB7uWtVv/7
gUXaWFRuM4RPX5z5U9i27Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8272 )
`pragma protect data_block
+3Mt7p3oRCWRB5KCgoqvAtwOnUsUrE0n5zxJb3dSxAPRfUEkk8yQamA/m1+fWzER
qvfG9vnLkRgeqCU8pv0LGXuaVRBqH7Mul5ijWWeoa7KlFBsjw4B03Fzyr9/EC14L
E5WObkEKLuOvfFVdTaFqimnptDKoUveD0+DF/1rvJiwAU0F+4/ADJnzBuIXJkeMA
a0FVxEuFzjoCFnvfGBqSHqLi9Jzy8j+6DSkAfkE/xrWRUgdZTNnGQjeJCni9ZUGT
8nWq11liZaOZED+plglWzj55n/r2YfnbAI28Q0ocqUiNlhlpxiUwBg+bXeAHSIIi
h9BgD6tgA+8Oqq5V3BnIxscWmv6nRRtZciCnbQCzrH/h8OdT03ehLabLf7PwPH2Z
8KStoGiOoZlj/Ih6Gl95XzEJ41omjs2AmdyFlH8dCpEuQOXFCYeUyDkN5z+7Og+M
n6qCFDTZL7gzMcWDz5TjDX78DUgLlD8cesWYiGP6C9XfjL1WCbkLFnAjQc8qRvUx
+ykq+8gG4LGjazywmKPbDkGk9N05qXa6NtzgHaXqMhbph0gw6cpjHPa3dH9nZ+lz
LFOK9WQe9sZMUxNo6rp/WrFBdc3+vrRSycF4b9S9Jmo5pCtZuoiN52MLAK0hTsQp
yizFyfZIkc31tEi25cvpZSr9nrMAzn0T3irNC/JyxXb+opGSXC1AhlGcKGKTKXGL
PMMX/bT3lCgE1ad2v+Aq9VqB5TQ7Ni9+S11uXmVjuOaVLosLCvNCA5oFD8BBU4yT
2x/p4xiWTKWgYkZw5CvQ0BF9xOCSNxW37QHUS4CNbnjtBtEb9WKTvpR+Ce26B4MO
vmCKHrTY7AVxLLUZS7H3GelH5sIkxcuH/I74XY3koAtjJjkYF6R52j03mtyOeeXs
V/yEMeaTKosTIfeOWmkUVddT0t9oUyb+MhRTQeJ2UV+MjuVPWKR5VipKzYYhBcMY
OTBrCJnX5Np7xbns1CTfhnxIJuOyCDXvPflQ0KXFrjbp0N4ZKHCFCBywdbn+Xehq
c5UA0Olj06OtCQKZs4wCVp8x3ax9xPKmzN3gENYJLiJmGP7L/gtHIreJgbEHf5FR
YxctHlGFfrD/JLHwB3BriPB2paS4tDZEYdLqIsBluWsBh2/I9LWgL4u2l7nFwYVO
5XEUTX075Se8dI+KIr8FOzoHLsZ1/DOFtNj8Y87NV4lWQZVLNJTE0d6fy4W9ebRe
pNxflhi6tseF3MemhwmFCw9L3CadTlqDgdzf7++hzh+hUCfnPJnBhcRTW/oxs071
MrQHV0u/Po3ZipX9D3tAoSzkuUIkZKUeVK7HhR/C7VvUynxJA8Ej12KwMnwx0Sag
fA3+XEd9vh26tiQA+bmzsteizMR5Kz+b6tolqOd327BUiVkCW0hWDrBVVxeTitMa
vmVc515nUL5uC0B5EvMEZpEY1kGxi/dHpPMUTPh24EQFUxOMoNLa0ozU/zXfC0T2
uGY0aze8mJCqDXk5WVeq63uB4/YphfPP12GHVwumm4vcSOuBA2SKWe0YglGsqpDN
DPjaIkvM5WSUrWFS2z8IQuIOhgk3FmyzP3PTeIIUkX3ZOD8kkOOt2iivBIEKOk+7
xMbrwsBUCZeLNILQL6psJGduE+8rjSft9AHp9LqXoyzpBNb50lUdNWQCJ1vGzEAq
QPehx0WHFQwZ3jsuFD8fQYZ2D1UjWFziE3UNykeZJGLyCnQ6IZwwRF6NYmB856Pc
FZmC5hXwYamvh00EzIwn6WfQZitXzR15WQSG8Ovfo/Ox5yXX5hlGEe4Nc7KTCcua
qA3rTEdxli125VCF1YiORp4dDXwfBpQmYag0+hb8FblLjugw79/34nens4neJa/w
/caaFMS7//22NRE3WD7t2lQ2yCNA2+sLeQmjCa3+/OfKsmuZ9m72plXBctRxN4xb
AUM1BY1tSa4XBWR8B82HAmFtUiAOuty2E7VFcdDSS7prBKKNic1uQOb21Hfgc9DK
9n9LCR/JhrjI/ifDbXShtSCTigi/pK03aweVX8H34ZQPeHMbOtReIbBzi8qo7HSj
BLGLOhY1j3LpBSossiO1YA6I38CDRt/AWczt4t3fPknb1d0DCGO3tBm/XD3RSLSQ
BrZmmoaUY4gaWOfdVB7Y0kpCkeZEB23cSuL6WvK0YLY963uaLZxJXsuaEeC29jJM
0I1AwLKobWwOnxIYqlJ6Y9CZcp3kDEc96JrzK7rEKlBZccII4OuXfZC4O8OAnk8+
S+qQrCy4auRQ1sgYmQsUjj6bVeDFsWhP3wC8RvhMpq6rzilymTx35iJrwkeQDE9V
RvuWePbS77RNqw0rIl3/6QuJDCJG2fV7TiL3khHcLegmUWR/dtM3psTLoGZk9eLP
f+Qw4mHA80kiyXBkketIanAdhquhser2TLhtSXajFoepcUQZctuWO3rkj4pz7d+b
VRSReMfkI0FD9U4fnut5xUHzik/fS8MkpTwhEwudRhS1BL8g9N7yXCykgaaijxSD
7TQHLBDuPLdRgSIn3v+ItFXXWRFF2FNOUkJiYlgl6wdhZCJGhRvz4352V7bXIpkH
TRj9eJWdsuvDjsm758gWsjJ7ZZ6s+5xrdz7pYJcW2S2UFbhs9QSMlTGIkX2AYcVP
71C7+Kkkp+hyDxGnD+kCM4iKw3zVI2PFydbCGcjE9Xt9YblW25uvYsx8QPC2svF0
G2N9c9kH6PLG3t3+IVCNb9ajs/E+FNvg+TbDLfTr6AA8UAviYF7tdLAZFN+Fdudc
mlv0uTxknCdc0B8dDgXANV0pdhwd7DtDSFsPNotqA9DKbrZsG91XNvHq8QBHo7YV
UoQhtclr+MMYULBZabl/7ts/ic/PXaWt3nfiXq/A0gYA6HW7S3MXB0VBn/tQ7HQI
AU777riNcpVX0N2So0XR3XGKBEcyolYCfOAlouoUvFXJ2Nqy1OHQKdFwe697lMqP
zizcVp6CnJdnRiKp50MFjLfedBW/4rdRGUKXTKe+VIFBYm7SddFtgSM/gp+PdevR
9NqteCrUweP//boazM+CtzF/Vm6sscKq9hV9wLM84pCeFKSs34JJEnGkGqKuZ9od
jEnFB4UXAX8cQfxgjGfZTdsy5aWzDa4/qplUEYPBdbL4E6aTKFE+QToRCTLKw2r7
5BVwRbGC5jmOCFqStxTuxQRApJ2kkEuxsW4BgwtF3QHN3FXc6LHNFweeTrc7CiZK
CeBd7HdfUONksd0gpemrraTKgql7HDSlVIN6+JH3GJ2VtFYmX/QbsOz/4Td0m6wt
D8cDHSJVsndxYmhKc54VSSvxkSIGZDnqj+Rl09bRV0676DwFkaZwZ2Wyq81aOMW4
H+wV3PlpeJVKkEfIaPtnSr55n++JBlQHsfzX5t7L4zw14kaF0aDazFznzYiy5Onu
gbqzmgm9DDEIdIip6CqSjtGZePMGSuUFF4vnEwLMMOJuJXzuteyO0XjvNqMmfXKV
xoECBoVyaPaQOTCDu2i90GNs1PRDtHEFMlefcLAkHtsijRm8PArIvWPfpsdAfghi
W0JYsvLRLsDCRaNpQQ/kZsHndbg9xQKqaSwB1oo/vg9qi/taraMAPZXhVieXqkCI
AK3G0TFb1GSPAOavtbHpnptxjDeOuAa8YJGpQ+1tCe8yuEXq2L2rDliCAit+4wwv
Z9bN2ZiTe7sxVBUqqKTGU82UkBBHQadKaqnEKlMVmssEd3hnLPf3LpqUx15XUwXL
dnDW/Y5cPYzp0VkTt9RyYHFr/WninKIo5bedzafuXVLNGgHGH4iU8j4zOgRmMir8
BzOcJgrMl1GpejnCzWnLZNSR04KKFZtti6MAVXHXLyWwaZ/iWkpcGBrnAdCDQO7x
qI7GhqpkLNgf/Z1PPmQiifG1C9ghq0bs92h+txA9If3lZH4iv9hJwlI0Xi45jWm5
yiHoYeYrnk/WDn6wb/CaxhGtowYmFFi+y2Xj+SH8UAK42WhFqitAqAXb8nThAdGO
7YWo5c3DI/g6rMZerQgltovP9KXDkOtC9hCfiNZFykUQ/c09xO5j/SyTgXNHDbtk
Az6mZNWISL+yjNOhraMqhMi1l3+/8Ew97J2MW8GKUZ6nVFKFsz0GAjZtVTSN1H0o
/hYc/i4AOE1wIFiIKNzWcxV2mC92lEi3xWTWshHox4Zw/PmtDyT/48pmOU8IypE9
Rsjfb1CDwRu6oCjsqnSxeZGZghGCMxOF6G2FJD5M6Htmm/Fvut1RRlBU+HXDuTUj
5KQLPigz7Jhtf2efWT9cHArHN9V6hiDdn7jpb84Qw1i3jU9jfNeusuvG3i09J9DP
Hi8Xowwz6QkknWnpNZ++JOqWcGtNvdiocUDw8oljoN7rtWgc8LodWnpDxB74Geua
BpLtbpA5SbXrzxGWdwh82FPNXblhped63liwPqdXy6b0Vbspdm3Ss8bajisfZzw5
FR/noWueQ1ncbOquNm2Xk+IbQ2LLYKqvY8yALJA5raqEivrXdNdC3HTp21xhQ9CA
8fObrIzcy1fDimMrq925nAB8pPfOkjCFJ+91djXXCiXjKg8UAO341aKLCWdQFjkV
E9aruRuFC7IhhHm95r8iqKod86+CphhQO0Wcz1viVMi6BUTR8LnPUjG8m5DoAv6Q
Lw+SUSJsk31mnJoBJ/k7342HkSifT2ObSSBiX1u0aH6QGDPmOScImKtk0THbaGeL
5olGr5CIUWk8MxMAicp10NxhqA4XqALS1Qixi4AGXkyZgrnpRC+RwDq9GlexFWto
fVmjGMagr7fQujKHgGNmhLrCjzht00d5pg9Zr+nuq71P55+SZ6fQYkRDnD2ZMj5u
NEX1FwxXJHTPW8gyXUhMuxr+b+JV/g4sDG5wi6ig1Kw7oxxiiMRII+aSr2sV5Wl1
BA5vP4mWqX2tqq805MbqgScsCaMGdVMfq79Auhe1bllkgNnsyl/uqPeIzCh1hZQN
/nvTbz1dEiPq/Mhdm7ZmRnVXvRIxNx2y4OX+rNMbXVMrAoN9ig6D1FEJX9E8twt6
opLzU0liQMbt+1c4HUY7nP/r/IQDXNGH8n6rDfMTB/mTBX3IAr0S4YmoAMiMEDo1
CkViJ5nGMxgnyehCDigtHkARj+t3Sd8xzlytUVA7WnjjRpCmeuRHuAvO7U59WWFW
xCgYKEcKPiPyZ8qPtC/gBqTCVQ7CuV8RpPjqJvfsaABh/9DbVVOS7ZADzZj7fvNi
0xgXxlO1Qt0f+OvCjcZZLT2r58GqeXgLrskQRAYjfx6QYPM0MlwWcxei0wu7NKWt
n6Dnu4oAKERJEeo7rRhlf1ujsgcyPRidcbnyVXlyo+zCfFG/AzVeehL56AKsvdhQ
som/UWxUlU9e3OCF8PYnnFfdXu31KHZH13MwTyCJmmd5ncz0TxBWr+h00hSykaWj
7apMK9mYY/7A4uCbNc6+u13b4MrTO8x0m9Chi4YrtzGEXdXFDg3BzMpyd2QodW+V
H38LMEHpN646/p7Iu+xvyXFPQegFBEe6z4dy9vYn7pwR8B61ggwMtz7S/5NvnnXM
KJVne5rMpg3IVsbznFI8joYc2fvQtBnpfLzrO9HTILbIOW02ND2Wmd1O5JogNEov
8BpDs7uo0MNh4opHthzwLlVFLIzinf/j40Q4e0a5WSSbL0gTeyyw6MJNhdddrDiK
xx20txlJdi/s4GYUA2OMa2S85rz9DZfs8xtMMfnhWHe9yAGM6tyJW8pVrIizLfzh
IuR4oYtu2GIkUpWrtqfB3c2wmpBf7ZgSKyRKnMZXJoTFH/OK3Y1QF61Ii9L9mCE5
XH/PpYI3xbqADEcPkiIPpHTti1pqtklCWhkCLWSWwyuudk7mNzo75D9oCm2eUi3W
XhXpYV9X6PTXtvLZqwDvl728XkBsHlqY82mMwn2q0fFiimdVQO+iTDElHrsURGIH
V9I6C4nQ/nAOVRfL+W3Zk1pcI3ChQxYCx/M18wRCPhriV/u+MsOpJpUYQpF4ljE8
7GpOa+oi+Yxq5vMB26M+bGgGfoviWYSzrje3VTDAzMXqUkw/GUMgHDuvVJGo5CLg
JtF2ETZYNuEMARyRiFdEov4+U3S4u1BRhtVddcf8m5hhNW0oB9f9peZR2TLwG6cI
5JjfWq9Dkg4XaZqQskr6G09k7iXQlebDoNSs/UGunWrKR+clq8TSUH+SCTKhZ4nC
9gHDddJuoHLY7pXEFWddYjNHWnCvuNz/VZqA+o58y4boVjiAlxKtc1qcHbZfgbx+
4q6e5H5TW37rZGq4izwMGWev5T3uhn92erdqeQSXieI+ji7M5nRKc6fWwVpiVX4B
f3M035NOwAYhKzDA+kyONrzK0r8Imyo9hRQA+v9/P2gH53BEAqi/72ns9B+AOZ73
p972KCJak1FlIOSRn2jaoIaPfbavnSSPRYYgQo6tbWzWNXjEiABx8NWIYc0RqUON
Oqsm0DV/6Hx8/37ZK+CNVIhd/8NYhkyjsmPQ/YYVfu3DxBln4Hm450fblFNvjivW
eUkYTlYnXIhcNOjMZe9jtN1TOH5HBwOdEiGinbT07KFPZR9+0ocIWJDNI0soAaql
18VOwGfxanvgqYEHbYmMkSuWj7x0Kd0Iye2TyA+Au0+uWybpu0sWB3TImlI9x2j2
OLlJGStaL8xTSxpgX+8fSr0NlcOFw0AQTil05CF6p7beHfQ9LxJdsDJ3brEbuVG1
nK2W4DDAzNT+OM9CMXRZfFt+zlZcnpaBAsPYYvtElx6YU/nkgXEG+np1v9v7qOf8
66JbwgzbB7hhTTrXukMUGe4wn4PKxziv408xm2R1zMIiih9ELktNrccOZNfjHBsN
exABJs/xRgz+lIf9LgZJOMz/D1i2UiHOvhyR7bo3hr++ggfEkTOWDiGIPuHoUi9T
irPKI5I/ZwZHrHCEiNDlxxIDWiLaa1OyNwNqpf0bz7CKPoAssfu9OFnAWqr7CWy2
+YNJs3u+NTCmhgrIhgIruiOq9w/pfa/X1wGdAP4LYc/Z2/NZMMbHJLjqcIBfBnaS
CCH+ZHvJMRa4ONJp9Ys/yL8qNgLbQycYAkfAqs9u1jiDDulk+n6gsXU8vAtnUu6t
E6JX3I2YPY7Hl4cnOFSTZ5uAlX495scQPDrNNwszROIMJS9WJpc77r5Xk8d97ScS
nhSEwTrv8JFc8Z29clY48vio/trKvk4KheGkA+RCvn5qHO7E3gaSVgvkK41tRY2B
bBSIe9MOe8LFr5uXyQAzLe8xXrOrgxVSJhEmRjs13wBK6o3eHGBmuuUwXcs8imgu
TjryBUlo39PxVGNsnWJobttlWA43i0GJblw4JbiJq4sMFitrA3BAJzoyb23XJLgV
S1A/y5GP6J+g6oVyKvlfVR6fNVwe4n5b91PgnEuBRthJeRY3vaix4xtjahZ1ZsQ7
Lg4zcvOK5VQmqPczXgD8cqJDC6FgqH3GEeH30dC3weB5CdQqZg93sqA0uFL+SUS0
BGrFMTOHSeRwOilLFVQZ4Ent2y8RHZrPfdr7auJVLxBOlsYkMBhpgCWbN7Du9Df/
Yzb+T+Yq6/RCcogmGshqIlQUkgGx8mS57S+ZHcCVYT3g9SATZXB4jEGVY4NWyJrF
TjwS/iZfVI4s2yAtkya2ZRB8kpvKH6low60VUPueXXeaEtVR5w5HDzW9bastPFZs
cJnhRQSqHrnmnPBzNlVRdKaIVgG2wnKi/ooWNExHYIzc8oTQCF8nKP10szWqNpov
aDGavWckn52lSDyxPm9ZjiycPHiKTIe1VMi/iPr35TYynLB9RoPyQJXKdf+7a7YQ
Q9ScNuMhbzGk/m9MI+dq9KNSD5K9+pflxYku+ghg+StItw4GAVWivAxnrFjYkmOJ
banszH5+ahlDxDdTP0bJNVe/NV6KKdj40gndKf9TwK4rZ5nuYD/mfkgZ5aYdoE26
7oEvv2u7fOrXfddX/guTixOyoRf9/DEFm8OaX6LculbLdsUHP3hgIduJopYG2jrF
FYBJr8TXTpjIunlRMpaFiLeY1hzKUaftDI3BbFnyAx1mdu25aO7Dv+SVfm3zcfVe
2MB5oDaX5QPxDbhgGKT6QR3QVTnZjmGh2h7FEtAkNsEfWjvUJecbsWCzgo4sdLYL
QcdcnEBSKyy3wQAoU7G9bHTWr4FBOzkeHqCapGBbtgbkfqoxK+c6oKWFN3kdnV5D
XEYMBmHhdsZF5b7tuUPAxe43ey/owyNBXX2nWPdWG1G/h+5X9cu1jHblHNau1dfG
OT8XzaGovlRQUzsI33hiH57Y0n5HD5F/Sh3CwVTkmieyez0Y6o8dLqdEGDTZh9NH
KhUIxlz18NXsx3IkZz5q08HnKPbwCKrg8Op4fIsqaOAf/FOJ9o4n2GzF4C7ewKMd
GpvG18PloGfcl0gBAc5EtyYuXCF6ofk+HFUIBstc5M20M8ZjNTxylqLIjrHjHOLx
XT6eEKRTmJM3YXjjX6MPaJzT2K+7hRENk6XJssHm5ApXH80+hzUVX0j5F/iDO3Z1
VaholBeap82rNNro3aUYZy7IUhmqmAPZ4DzwuxHjv4bLcP50clg9O2oZnYzndopd
L1TQ2rtcZkaZz+wOZEho/NbEUdNqTPGF2z7DSEjiJD8VqceP3wW6qtCrYDko4G1Q
eYqz2eZAuzQLNQK+b0cZmfB9R8z1yc/KqiU37pZpCr5bWdk6tThW1FeY5EP9wQb9
Tpro95X/kq+WZMYAZgbngwcIJf5aehUwjLiIqOgMZPRq6l/gSbCgOc4K7sS8BrE+
VF/FCH5eU330EMCuzCzOoc2/+oV2tRJU1pTSYZ0n1hdyx8viAlezTXGqsm9i1cG4
pBu8uwJqtQfSerBZmYJ5Tz0DrUwCox/4ri7tupb8ouZel+F29TjXrxY1gGGZHR3N
UTlYzUNCsAS7x/Yc/nWsguMJGk80CFZllhawWFdQZTh9wG7Aaj4UqHNDLzVZCDxQ
cPympD+2PzcJZyOxVLe/h4gIx9KB74wgf/L62NsQyrk9SlLY1zbAXrg64hqB5PUR
UxjgMYpZhJbySMQOOcWy/EGWqKN/AjnkifaoJLFy/ftW0th9Dj+xK3XR/u4yCp8f
b9IRQtF/Z8xtvu695tPajP+GKYNLTgujAm4/1wdlFidNfhlKNTq7ozAUF1Yn96rR
T+bu3wMFOqSMsVYGCn/90cdh1e8NhvA4rZDL352BOdCBhTWG0ncl/+7Q4keX2CWf
hCsESwzlBIxiJ4fn0tfBF3YiDAFLtobJAtJycfiLfr+trY8HF4/XHkQyV84AxTQK
wkzW1sROJHya+uSni6zIQDY2WljzWOzri2wfgerCcoz7g4yCeMDs4rUz1lMd/UsE
O7O8QUCg97cQHu8tPSt4rf1RgG0GBtqFiy4D2W8wG+8UqEpziZCPyDtn9HSmrqIX
NpsleIiebyXJ3sbmruFzxSEQvF31ba6ZTGg/SEa0RfSnAhKfnLNIWVAnzyFY1Pj+
OFTi85VezGlU2XVSsIjCxAUdsneazONXGiIaqPQsnUTbBwNFF0DC/bUF7AdruZIj
h0wdqA62yR+BDoT9up3zFAPD5ni79YMscDELIUruUAb2exJvQeQ5a0gi0/w4Pztt
9Ujfnj/ufTIO8iN+vGdgv92igHVpL7zuutyLuHrpuvbBRWM9HUZJvO6I7hV22q48
1hHO0AthMQXmZWl7yr6xOqm0x0JX3HmProVYXfOWYpEFuO5KdiyquE0YoeNmOnAh
VRhnkP9JD115EaV+atdbg2+izp11n0SJpGcUgudUElwD+U1Lexu8oggyG00OtIIO
fplrQX7+I85/ZPRU79GYduuBXfCGpCajjZRvswVgwa+2I6+G7icnX0p7bQMOmiFM
ZnD5GkPBG1rNr58yzu5u5Xl5wqEaut2fLi9ckqYw0pS0t3s1qrTLoa3UX5yHoUQ7
DuMaoeHLvCLsNvtTTN1Znrz1N0fnjTZv9XFcfDJD0sV+1TMFbGxwGiRap75RN8Sv
46RdRoQaSCv585drceYNLXtapT5Nw/sbfRWeAet6gLd+Z0YVXzOo0+QJp0DO5rjc
ezd+ExnfhJqUOY+nNb122tJ9fNd8eAr3OlLUnse1S7cJ9EchXxkC+oeCk+iR79nO
Iq//LrgW/UpT+O02bDr8bGD8/d4R2MwPDF0EPc1lPn47qCRmacGsR7xirpsO4ee5
AMFaKJUygq2xbxkRb1y1jIi/vCntbZ4kQ2tDBM4Wr66bUzQJjTAaUw6iyeQHntvE
uyNVUx48UmjUxi/akfB95/JlgioS6fkQJpVIWRcamtUFRbgU617nQHjxegcmggPD
ysFpZ8vtFMzRfCEj6owlhNc75XiheKY9xJOdnDegVWVYzhBKvUwqKV7vk9f8pw/w
OkOcv3hRJq8OwoZkQ6jSx0hsMguZUrDAfN/135aSoln1Sm9NrJJHH3YobazdpAGz
bnOZWxji9yhsxr9UZ3CThEgItYFxpNj+jl9laJUcgFbTKoG09MB68ya8S7A7hIPh
lVKFLXL99OZYETpfRDqd0bpcVL1kzi2l0Cp4Q3YPQJ+t1yl4qkS6aq2r/Tqiv5lb
IAVBiwcP+nNLud5Zz3l7JThdPnBoqpAfnRg5guc1wfs05I0QX/Og3/clvPgDk9Tf
LzgaGBubVtZyynXOW06RrQdRmpERSHk3LWRmDsWUBHX5HjQ3HnNPnMqH/1zcogTV
v7fSVwzUbMqSo22vkQxcXTodsIhy9o5juFwvZ9q6X1y90Xi+8mjSMjBheCKbaV0i
Z8sKDOv50CB8viHSnu1ghCyNZon37C1X7EBqsNJNn+vUOG63GeFzVdGmI9gmdOys
Du3V8wiBfm+v3Y6xM8md8HIsMZUUR1/L5E1mGOS7pl+nlewgJigLAOfLZdRAx5AO
7/AkkhfrDTfdfxJ4hDEg3zwsv6atMdZpsD/nda8PK7V63hN4iBAWiXuIn1aB5tUy
x3nUa26LfK8n1c1nkQA3CylKr091uVkfrhBrlKprLJSKcuzi4TV5iWTp81sSqTtf
bxhX44H7LT/zQXjAwLQw/Na9tN+XY44XH/3WUvWsaVy9+YoIR0ZanQbvqbKJuU89
PCOrZ3ltpDxfSgaseWPe4Q==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ABqr+3Dg77IIQCmfcS7T2UKqRWR2AyIDeN4w1tsg5h3Qfj4IW3BH2likl/ijgUV0
Mby3XisKMblwSq0VGYVMUOh/qQMYT/cG8SJfsTiSqE5qmPh+e8rNE7FpBYSqS10/
vb//tlwjggEt/ZjmA3kPQRkJH1nZhkFkXimApbAUKX4yzkloNZQsJYZ1UbmG3RNh
eF+9cogtoZlVvSWFqdQvAp+bS049c+HZ4EMOlYlt5NA0YwezUzb6enFR/qBAzReg
42y8sqixjNEHNS6IXsXScqBn1wwr+tFexzQC+1vrHCRzM9xvSkSiY6fljK6Um6ke
0c/72VS+LXToPek2GGna3Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 21232 )
`pragma protect data_block
tHn8tnUWgpLlOACEng/ujg05o+K/DbYJBk+0x04xwIG1EwdKpHgKDeMs6Ezt7QbG
1JQna8mkop8hylkyNLnEN+/FZgcYFB8Civf9eJC2rM7IQ8aQbQ7a2pYa/xQln6nl
AxBFD9GWh3UcAC00wXjp/cJN1ksoFR6VXs4ys1lu9bZoFqpvpcb1y6oIKodBkolz
r+lYMrqrPxrgv55GF5iQWcxNwXfExkYS6JvHEan9rlvHQtv3IeHycI1xTAkmdYvn
59vaGyZyk+pWCdJKfNV3rctySzY+ufpFhdh+5E04sTYDpzN97TPm5OA1clgdii/B
/0rVQ2lsa3HxjqBHtFgn44PpLF5Y+O1eSZQ8yZuub5uMQ96G8UXaURx68ajmOs/Y
UcKwpHo1VLRyjgO5/MSSqLx7YY49iSYfgWCiJGxgq+IyJxDUW4o+r3J6Za8mQ0Cs
5DMJ505JkCCHJlU+NlOtJR1puNVS0Pud3DXt1usXtUmQFFLHq7V6PrhWoa0opaWa
KzphY8nMBsZwWqGSYUtXio85wbbKqGj9luaaatIElxwj+l3xvLmzYhVAUVj5A0yT
mQnwLHuTZe0TjRTCTAOnElU05rSbqN2XStY2KCWT6uD8DROvZiyU5EZmgyycJXBB
mlmptKGSJv5yNLqGtH158V+wQgjv/Jx1iPNc3AFyNUh1pdUld9Hu7KyYvMJnWzTU
aG+qa8Bg9r4/ZebRmyBQTPCW3AfTCyrlLVT2LgB7thpUPPNki/BuN65sB0oFGvKI
sZ3fNn7HUFJrxJqMsuA7GjnwLq1ywQ3Yj8yv1Lt6B4clJy1gwcNvqsBoF67YUu/w
nhD0kkhaaVTPi6rxdr8JYllXZzH7xVleCcs/XiYGqb/2C9FqbQFDqMK+Ux0+v6XM
/42PZE9ZakL7qxk0iOvMMSemyHld0TEP7dSBf/7uQL7XmGXM47KARQvsPJRe8U1q
ocrpnnHOLfS9F7nrTwlzmZBI6sOe6lysznZ65uXSJdN6xTWon4thLNEftGcJYfWl
WzKPKFvl40GJt8SH+dWjtdOK2qxzq6HbG/jrJR6B8npK4Oyerf2m2u7d5lgfqePS
HtUMfWTtrjyZ0sjaugm6B9eBZNynabYXqH1RT05jPlKT3y1+7D48SZXVwRm0AXOI
Bj8DXPV8Z1A973yvd1lwzQ3dNXsDq8UZZdwdoBTRiYXCsEi4B6T3r6V+WzERHrn6
N7fLiykisVKGV7H9IpnWvwRZEfmd7pIqLQt8ARfxRBvrD8+5t9da91txxRZQwoBR
3l+rCx04P5jXS/pj4Xq03AhypJsA7Pd4Xly/sV/XeKFiLjktJtSP4RAJJXaVhBOR
VgBAUVkvQcEkGyqktRkVKh1vPcXU79nzWurJGyhDU2CKgRvyH7vdFwx6DLV7VWhw
2NFJdhcSa9bcW2zs2zidk8Zyaw7eoE9YzEu11f7PdOddOT74Umrq9eqIFFyfrLm1
0QGSKktV5AzH5DdwrbGdZ/lW6NaT/yTyostl5uta4nDwjsBXaGi6dtVwkqWaGwUT
asxBAY+4MWvXOWFvBF/wkkjagzXbIS7BRzEiezYD4dxvmqc/4JoO1fGmEnFt9JoH
OgZVZEo6AaoOE4hEYzJ7Fkp1Ob5JIhaOmNPZ+q0sFy0J1DtOXdIhVtAjVmsvT7om
cT31SFXX1lBT+rRJ1YZuGlkTl0hmEaHTwR9K5DJprVQwmOrETD3OkvbyAjFK/f9j
HVIjYSa+S2tSQEVZvWkHC0sieOdVYTZOqr8y137OS/TAXfDZ/drAZQyg6nBF9uVj
1CtUzZqwKBH/+vdi1xxdiAhk6QcIGa4895xe0+AqA55w6BQPaXRppVFlPrdPRfoy
mZjj0aZyuhYqKTEBgdyToHUqV4cx6iIgs9GQMmO4VajReHqMgIQEJfVe9+G5+s8z
3Dq9X2jv3RR5B+UFNSYIN5F0O4qUX66gv+wliiDmqVcIjAdYkHLmJhZkuTNkCUBJ
8X1/yTtmyVtnOURnwY0wDGzBypVLVlfZHY34pys1BBxtY5N4RX7Y2xOvGkeZvXAk
C3Nk62LWoPdoXMRHduVGOYfy3l8fC0e41KKoQ9wy3rOi56mUXKnUbIJPRg4guidu
1qTbF24BOSOqHF89aGWEVw5xLNnrRvLBCEwicBqJlthtSujJNoaRxlzgGXQGyFAK
QiJhXBsCocGZYcnagD/eA9V5kKpKY7R1nPIOrVgVogwX5scylwNJCcNIvlXeVpI8
XBRRC2jNHJaTKvbnUvtk0Cn273nyqhuiHFNa0YfZzcl6J8zHA9LgwsZXEmfqGx+j
2wsYy4sBavVyCgVOxBnLp+DsZDeTtTMWGhLZMuoHOz5zJtjxHkMHzzON8nDwCQEu
iTP87BHXlGo5/gcbZuiY99oj0z740oOxu/fxLBOp7gWMkbwA7dYWXfnAAtHAbdl1
4Q/iItpTwVy0yq6s3Eh89jeAtvr116Qo/tMVqbKJlg7og293MHxphO2yYDZKVnv8
SSNQjAiox59ppic62Qwu+tM0vpR2G6ANqiLFy+ArX+6hdrR7oYh2AEx1QvxcWvv8
Ntt7Z56GYLvj+p1W3w/NDYQ6uFHFbpNP17AEaO1zVWv+Qcd/dFJuTdNzEOFwZyI0
bsam8YktDsaF2Ija13h8V7QnJPS7AYBoyM7oenfXcBxLsKVg0DyqIog7lw8Frzbo
fZwhAHfy1lzQx9d09CX36tRv+TqsyhxGGCn+7Jcqsa2WkzJdALrbUiMbyzUTQ0+k
WD9+PMB9QLx8Iizgz1jqDln8UcgdhQs9JNqdTPDzufB3xZubpZtghfGmYRMLbzaI
1Cq9zPQ9OU61BvuSP8zqFBGHJg21uUQUBFywxrWopmaNDQw746FusiOdq3dISijI
U5KaMPHzW8VeZIEF9GrwuCC9ofjLAK+noA/JJdNdDyQHMz6tCGIfE8L9G5xkagYX
hNn0rV5yKWGntucRXOjT544tOZG1l/yj6GTHs59oHsKhtbMmGvWnIlnNt6wFRhxX
vWd8wp83lk6c3xv3dOKw9MgJRK70pngYkFS/bY47TSLwXLkkHgFqQDWPOimcHQg0
JRJrBXRW4loAEi7lX23nTfLn+N5VE4srtrKxuAk9V1XPJRRBBIE2WaNI0RnDZ7HO
BFEq4HPPU/ioAmP4EE5wcpM03JEOXAp9qg4cXI53lglszmtHWadlpKzLhJh9EI7q
tHZGhoKbwtthPqxZ6n/g0suFQtDwuwGZ7y8SlWJrax7UK4Tyf74XUl2lYrTpbYw8
WdU8peIC2/xoKmstNt+XUvvqNzxGJMwsgYum2j22BNN2AiawwJYxGOJd5QUH/aZc
cdlSCtfu4EnrUa/6NNENNA5EwJJEECMmoYjYhAO9oO7dlni5OO10uJMc5ZZg2vq/
JUXkZH/Lwrg5+Xz0tEMqTNsAK7aaWael70cuC2XujcMMLnSS/U1PaJvejZ7c9N//
bRcIi23PxwMswz4u+ydYpFjGHNGt3oM/trmSB66VK6Q4Mh+uVtFWaa0KXhFq76K5
CLilfIhjO2Wr5m06UUsMqKx+OuBKCehlGJbKa8r6AhgM0fG6XkIW5HkgdTAsNFBu
lq8DWMeFSIgtbXtr7+7IHgAuwLLKnB8kkpK1zELrG5s8pzaKWXNFZJQDpIP/GvJi
NYvIrBqcWRBVMm3gtJipV1yqNEfWHubGyCjP//4S1Cxpz0LlFLYF1aMFLoyB0NnO
YrpqMb0yT64aGk923PSl1GxLm5vTO+shC/3ILNWKKNLoZMjFJIiWlUgm0AEIOxou
Rh71pEjd8Vpe5+5FLSVepHTNb6O1ZBuWzw68etXWkoIHh4Lwj1U8hs2H3AvZREEb
ldULAqHC3oEd27XCAAQJ/9LJqgaVUuZJ1jzuwf8+JnwZSNd4NEUAUlj0nys2Ci6D
dKUjc/keDJUIN8hBPDXveSRgitbmFQvx2wwjzCNzuyDwZv5NyvGXcmSxiAmlzakU
xzCMVuNPJrIrZxKoA8InOTFwHMMGtttp7EdWMr3KWXJyl+klz+Bl3ELQsmFyoQ9v
fcuTXzyYewWV0NO7vUh0ujWnLxQHjvwnahPC5vKd1yWhYz8HTUMSEXBx8NoShmz1
hmE3kzEgdGVowmozAcNagMf/jTtB2VngCy25afrlqONLoHZhA4zfo2+dA7S3/NJB
+Kqw1C2vA4i0wfs4W+jksx2z3TTPi2idi/ReVJqnj/dFJwP6yYEyeougOJnHwEaf
u2zmtTMu+qvhXcqkxQb7ocllxQUGPmMFHc8MHSMiHzaiEQ2yh3PNvuCdWFzKOS4n
eCWvvUR5mDuTZFnmyztrekfngSill+MwASkTv1+pmzr4TmpA+tZW3D0PxL4q75xo
yWKaRpBRTY/4V5godG7H3tzwiyTKcJKrFaga9YfogpZbCrmilxVyLojejIzpuugL
7Frfpq9/hU0ZpqgFZ0xlg8/w9yPGjrzLXq5YN0a8J1qbhcfuPTrsh3VmAvOMbiCu
NOp23FwMmqtbn0tG3PwOzc2T0ftos4LLSSYxiyZwA4QcPMJ0nCKf72YQBQfNBWkU
nNKCcJl21t+3TVLpdxiMXMUBkdYwzbo6fM5inLNdwcrIA9cRoAn40dgZQPq0M0mU
l4a9hlahrw31umuvI1CSMfKF4RR1aL+EoS9t135kelNgsybz4ClYDDnHlXIJ3ynz
zTxWlR4tGuB7ZzTatyyE8Otx7EgnZ8CfNd3sTM7HW+Wiw0O72A2hTZtVEbYzXbxa
OhyTOFeEpJqUbp0zh+vssZtrKQOimiarBx8ahJWM5LhzgyUt6GH5iVELB/yZTWgm
8aLTARmtF78BK4f4bx4EVWCXOtBA7J0EF4/lIBH5Qqwgh7gKLoO7oTheyscjoEZA
rmhwqNRNoxzA1R8NTWq/0Qd+ygV2xhEfUHpUZB06e0jEgyUwiAGHA9AQ5fzwcFjJ
vrooAgeuhdBX8XQUe5E12IqnpFYOxKFm0FdsIqbNvsgLwrlvk2Tv1fnhL7IEgbOY
ByzsWu3qAYn/pdlMPPHqEnPfbLaPzqRvtoRAWqKWRouTLjdmURNedIZnSsnfYJBg
ZG5i0DUGyY3WDx1t8Fuye53hU7tG/gvv5Lc59hs5Vbemoi/1Z1BxGXFw8c3Joe+m
MJW0hf4SIe1tLXhWeVJ1OqTt824CeD8dwi6UrDTwZ/j1EuhUYx5bDggGmAoNg1dm
AHhpaeGeJgO7ZLwuEsoNeIW8hFTP3AbPGLKsB0TFmkciFpghE8NaI9YzxGdFmbpZ
NUQJFZ4IIbNo/MsXBBS21rn+dSakTj56ul+IweS2M6VjwiHPKPm9pybaSnZTZcl4
y/yN86KNQEHa4uyLiABkEFs2WOytQMv9A6ccycjnOgkaMssFhuogC/sdb81yhE0X
gKamgu7BNZquDfmLMrwZemlhIL4WzxMgmZyQ9mCwyn0BEl5yV/kXayZsO6De159b
zr8Shl7Wi4EUCZGnp8H3iKsI2eML9O7ZzIeuRDGkYEwHvmp7wQeuM5239Rnc92lq
7XfrmyBrmfjdSe47Xa0Ns7T30EJ66i6rX+GEyxW+05gvu9TvZwmLzrjZjrqXNjde
QONlFT+Owg7Z6m5eLOn33OfihxoVy9pWxkxLo+qOB0L5cK9q1Wm0Us0ac8HbtM/x
6va+1WmmttKDIaCtSRiq4B9ceZMcq6COLjXATp7Nj6nJ/2f1YYtJ2FAtLwXj2Nsp
10f7sdhWR/2OqCi06KFNO3PF0ajnLQWTIs0DMj94xillYRiAsLtPgXd6iKQ4e2bx
j1ToWmIYI3Y1QntkbsQZ0mUw1G0zQ8O/uTmJRT3t9dmwtcK/2VjrY+Hd8whfF2sU
WdBFh5j5nwjlRqrPgyX6YZQ6q66FjxL+wA44kBLNP3mmWGx7onpv8Pd/1GJRkuTF
j75tfoftXg3jLikfBlut5rC14R9QGkGHDfRBIlRY+f5tuWC/Hc5GteQOjJBGYSua
+BTpE6Y8uoEqSV3a2rNZQINcVrRh8u0kU6JSnDiFAUk9tFBW6C9TMmt2+OYqeizD
5nbfHYNcElim1TVr//5aIAfRBGpCzZlGjFraV3ykUhT/rW2F5Mnad6YGUPPuvxFu
YMjtRRjejsR7qKe3IMrO11uV0R+xuzhiEw1ZL4Z1PQCVGnrpYmvNAFCM/cdk8B1g
s13jcjSW2AWLUCSp2BeNMIETpnKpUsCAbAmSUNFrb7PS5GJjzSa9JHEunLMFh96l
NZz56EIFyuzVklMQ7MbOfvOXd0RlepBFb6UaC3VJIPUN8W+7Mcndcc9GYSyabkeC
Vgn7ePJcPDI4mh+ltCxVcpFH3PjWif+n96FqtnbMweQYfcf0UJIfN1Z6b1XJF680
ah+h/UUbZ59ZRSn3/P4uflac4/4SQY6xNvzwqHrgiT4m4YQkNXqKWeAI4bgBrv0o
KT9WrzHsCJDMQ72Wh/bGlsRiYvLFQ/dRSCyHdCZDyjSKnd8VuxmME0U8oO+Lvw7g
n2wBO1OKLYWus2/SBj2hMpfZywv6IXUG1yzzDKD5VklvX3ZMOsmztkV9Vl03qQ3q
kMHEQATKivPcqnTVhCJ0CUORTC3HuIEKU2xtj2hkUAMd4HaTQDrASgjYIFtKVxnC
oS0X6FAjHttx9Z68bgFRJf4/tno8Nm/yEnJMCrPKY/xw6HELfGCT2An3zdIXfDUE
o/tKX8RBRHK66EqzpGhbO0vh15JfCPm1RORZfxjUBivI3rTd0sY0JOFTX8yVcUm8
gyg4qH7J21O5TLyfQ6YWHlPXFWKjSB0xX6gC+3CVvDEbOaY3obSJrUrk/1WBnaQO
JPFtGQEfVuIcHGgB4xvx8aXUR4329Cls3iWUFHbDPabupfF8OTZ2C/EfLddwulLa
Fx9thg+h7L7ahAkwGMI3HC8qywEC7GUukM02+vOpa1YFbF8Mgzb0XXeCcdXUYX7k
1Hpp1FUwxTf5yQI91TFpzUpBW5nAyxsVV+ipRz+hvepmvIctEg/g542+wMgpGpF3
uu+Ti7kg04jtypBa4Vbrxwkpx+3zIF5SHNBJSPKh6l+EtSQ0GkoEy626CBj5Io2R
COTtxQhgnl6hXiVx2byOyFDcZ1halLnOArIJWk3qluJSscmJg/Toyv3FY/0kJZyG
j+inqEKHzU84yR3hvC98aC3UR6hULaEFAt86HFBnbmfqsbE5N5yJMNA588A0/+Kv
pJxWq/LdO5Ehoj3XMY2/FXw+gf9YfNLV8AAkvzfI7nnJNvW6pOLvF5VhlxkAhJk7
v2qUo6y9KkmjwfEO9xk/TTesJECXmNuAJAiF/tMkelHVBMmHZoskNTPDuFUjI/sn
w2gfbBLiCld4560eH/D02F99W3+g91HTaQWSB5EvrFpgDhW6tmRilM8DNfagEggL
UX3nme2cfrjlSto8PDKa/3V1VDgxRRKuUPjqdETRrvZQLhVZSs7+Z0ybFAYMDkXl
ZLC5W7XB0+1ths++GQQXHYD5MCektBlnOtjs4z6IAHB4GXFOGb2j1dKMPlDo/P/d
3f89hxft9q3FnbPXtcD23dhaoCgaeaOZjuQYgX8EELCKIeARY2Qeara9FIA4axpC
roQ4j0MZXXF2VnhRYgL2w5urIkhPzltJkl7uakf9k0MDH4EQSNQA5DTBQFHjnipw
hz7hBe2/6nIyR5swivM178AWmKVGIQAod3Oyp20qxm6pVvAY+GmDqmFnqnK8+JTF
alOQMMIzlS0jN7rJGj5Z9C/DWNG472KantqQehDY3xCnTYd4HG9nJ23dWSGgCgWJ
vLK9qVmTxguNpozylQbHQuAWBOV5rxBuSV5lyzzpfVJ63mGXmaf9QJrvYEMvBoXF
fgjEhmRNoMzAU2CDEOmXICM35iUHoZi8LJEbmj1hsgUheBqBbdegumq9Xp26TtGp
cJQmhqmjHsSgoaF1DD2eqzFAOT1AGVQmfBMMtoUGZ2pmJfbbVNOKoQjYQvo2CLQ2
xfO9dj3IaKkfOBtsFSJnx8jDHkbQJOb2CueZSFegaFRBjOcfUIYP/qaongUedMYU
Q9wW9RoTMgy1fQCkTPPP2BQD//gkpgS3V8Agfd9TyqIb5JdzoBvqyPV2bT6RZtoI
EyWqN23XL2KtOJtIYq9rFkT/rrun9j5o+vdkzXiJRSUk9jG4TLO0mXvyhyJinokR
xo+apsWKS/yHaH9kDdaUgKa/mfjnk7+J8nznsNyXHhncls+94+evBi1XUmrpF9AH
nOhWK32lZkkoBmz4VQD1D4/f0Iaw4sFg1LhdjDDji5Sfb5XcxpICNYJA6ouv86kQ
HHa6qz30jg56jTk/tqvKnnU+VjCiV7fMOJFBLIk1fl7NMsnHHUsPaLv+HT9uasAF
m4WMuHfVTN03zJphO4MnWBMbj3ORjQPel99W8/6RYTk5mDRXgl2GcMsb0eM+gKlq
aPziP8k5FOG//Xu5yp2bF65H3Pu5d1o4LzoLW8u8lE9erl0+aCh5BWvu2CDH9JJr
xDITlio0djH3vnxIWZO1YeeFZjR50vrD114Ns0aRPCcY9ZFHGWPUo/zWXj4lTj11
njuUwkYsB+uWt+5HKIX0Cvv24HaKwghmANUnau/fndoKxL9pVdCD3vhYf5tInSoF
nAvL6Zhy4UGJ589dMyOsqXd5lkOaeefoTLKhVIJL3OG9J6uQ7bXjxOEHytVVL3d+
g7C6vOeSf39jtMWwHQm5+iqCobIkEPvzw92P5UiwbLb9frQMyXElxfw4TuvhG/bg
PcZmeC/5I8l8GUvEzPwSl7rCLLjCWQVE/UuSLnp9g87jqpXBUqZHmJcz38CxJ9Fn
S+xW7BTB3oQqd1K/3wQuK9gmJFj2JliRTZ2eBEJmP9HN71UCDJtAmadIrhG8Ik4Z
8oBJ7z3OmyoCx4YKp7MQEao6FYcjNXiyl1tzlBZZAPmntc2ZZIibAhNknUJ5suC/
PTw42GVvdxNPHwwNZeFiCvMvbd/Nwz3vmwP7qg0CcPXBvJ4m2+rcd7RIvni4obV3
NZ1pf78jR346TrFAQwh5lUhGEb+XG0dzz9j560btlSY5Uz+BWQCNhq+lITag3YsH
FX97iqAacrrYUmL6wsZf8F8sN0Fp5ZRO39OQqWiHuy34JcZOCp0Q/t3xlp3oBBKx
YA7bvSfP+7WBz0TU/6v5rhumCw74OWV03T9BySb2ubOYsisufeYtozHxyMHNbNno
C0yPSS4doq6BQOUZQi+6He+V1pCNiRcKB2ZP9aUi2jQGtEb15UCtDCsDZ+sZZLDD
g+eM1bFq9Y14GIhdGj31BLL3auTPyWkP9ZidKfLf5UmWziKsWj3/d4BuHAsw45No
M6U3RnggJdmgh+R4mIizDs7gnoXIiSZHRYGV/m0Y7m4C1issRwsxUHfXFkYR5vrB
vcLAmizXrxMkg6iwb3FYgx1AW37jt7HkHHSsp9owXFOKvqGx92P9egr7FqfWZHa9
aO5JEhuYHE8V4DDM3L4wi0kl5HMAhxWjIxV6E77yk+jfJYSmQ5vrcZ8fsvM2jUso
F3uQOWbuHzbY/3+gC+t9NTvKC/3AGp766DqZfyKK+iWiHKZxPvvqx+8ONwc1RFwg
USd6r9n6I/yxmAJr+n+sCljsN3vNV7We4Jx6NFmJ54W7p5ij66TyP7KTWwBW9wmH
MovLXptkw4fIX7JWu+iOs6NSPEiW7Gw7aSUoQ3tNEa3IPv1P4GFrNlo73crGCZkT
SRPpdCVAA/TlfvgVNnZb7U0GtjXJpczW/RkDkJv7GE+b2nFnBDKXsGIdExYEFlpB
rPNbaqDgbOF4QnLI4OFrEYJy6YqsuOq7T5UA+87OwvSAs+Nkb3OxgB+8Ee9JCSmp
sUPvOTOzOkTv5jUp/LU2zCp+1L532ER+yI1CXTwnompb/poga0PXorDzEHI9za5s
YTVtRF3HSTds+j22s+HH0DC3jAB+nVF4tyxYeJ0NnOZfVDEbDrckNaW3+BLAfRrC
mqduOomJsaJudhFqWZAhquqvkU6oyscDss84C1y6tCi1LlZjGZjA6mor8vi7fk3c
J08hHYSocnq2JCaSW2fQDCrrwvnDmAUD35rrN0JI61EO+l7UGPLTGHKKTzY3gH5s
G+58LChn+r0w/RhN6tZ6xWZS+qoPEA0E25L+TrJdeaSKMwKKwrpKjGgCVj5UDRzN
eTCXPjHA8VAQgZJpI41XTKhSyfWQIF2DRJ2X928GpTCQ2SyiRy/KwqOo7sy/sdkV
g87eInYzjDgfXdof/oaQ94HHuIQvD+2S/ygJBnbcJIh72aubB25qZW1R7PHQVvEP
W+X4YTZ/V4ZgT2XaKNLWh3bVwM4PK4aRp0RkI/SDbjGB3RG4jhFfu8LrON5mtxSW
q8TPINNzbakLIkTBUAgA0g0bnc9XZZ0tzYAM/iSoV4PWcpSzTRagGnrwNzwzNuXU
nm8z21nv7LYx1QR3diWkvkERybL+Erm99irk3Fa0BCK/RS2Ydvfrz3L8RZJoK8qM
Hw4amGFt1mdJ5R0CM9PXbwt9CR/HQx6oX4z5qmyimpB+BcWXCDcHHiiYtiUGmpZR
woUsHANkheCjYBfa5UeJCk4j/SdwplLKjmHgThxdiJPf5+k0F1b++NhzUA+PE8rX
qqavXvJS7IgPYvxuQNaHa5ue4gEQAvoCxeXhiY8gkrVhCP/QmywCr2eqn6Q5Sc1C
AI+hv9opAWueNc9vRBOtxSGSU/x8OP/Tsm/YW6GO/JETcq3KWRZs3I2AjiSyjkKa
O+lB86fHSDIwZNMMzSpdNdDufTL/fcVIOHswQqjTDr3o1ZgO7li21BRbVRDf37+j
pKEdzyYZKSEhPw5BmPmr2FkOlBvYoDQsP4U8YN7TJWvTxtjMnVNlh12gRVhS6HNw
lt+hspBzDUJYrPXi0LcRu//j3UWezFZETZ05HtiK3UD3lrUN4F17v69kFtoy0LZO
VAT20QB2mLDk2ekVyVxTRFCJy4mIOFz2Cmf4ZRDMoRasOlz430jiPiWcHyRMl8+r
+DR1jfV+Fjrk2uBtrKURwkIPRNuDUvaCEAFKjH0Js5SN1o7gKdYBUYElLSwG8t9f
3mXKH7tqzysofoaP8nFMWCOoxiejyQo6ICKfBv/xPJNcsyQIJcgdvve6z/+VnZWv
hNWfY8KsIo4017QedPJSOrKKu+UMo5qymniIoNY7ETFKuG6NWwcL6uSr5tYhmNe8
qgB2aZ4sI4PxKeCknWKmtw4b+vJ/BE/zMn29qcZAsCEks7P1f9qy3UuchSCvN6SR
stgnLOzJ/7U+ZoqRo7tY6qN4vpiIjN6yb2xiWGvvI9JDo1B1hkIee9cUvonhygxh
/D8LouppByYHulagen9pLD6enLk8M56OSNAqNIv4cXVY9ihnM27iTTz5ljTB2tiv
B8L31Q2URPJDAHTzaec2m3R4o6HrCK6PDzraKF+Mr8GNF28RP0bd2izBErcUrH3J
bJvmWz0UtBQrIQA1nXhM/uD/PVBKGQLnxnjJ/GwoyqavM1Fwdb8NYqmFA5G0ahFO
EG+wXlfzQhWVrYyQ2P+RL2lD8ifsjaotXyEdhAb1Tjad/Nfg9Deweyuw9MG1pMsr
fcSbDegQ9hH+rXE4KgMIYdgIen+Us4CZ1exDK6um5CwUEuY+aTAKePrnKW9dXiKi
0w4Tr5uC9tY5epDoQQJ9aM1xqUrd3U7qtD7vh/LJxQdsPfKou3EYwUDwe4sAkWR6
B3dU0405vyagwZ43nw8Sb1P8aj/RLAwZ4lc1+VPn0KpqiQgaTCMvm/ZKSed2Ijj/
CCgZ5U/vrIdsTOYiaI/SP2USZUzl6uashtRHw/O/DE9cd6FkkjoAEWgDM6K83Q0T
jZFKjQF3K+RTrifrxLoTfum/T0+RCDYcZOVw1eIvbAJ5oiN7H9rcncnmc0yrtX/p
PcOdmgbIOyVv0ISAVByL0wNFjPB2SksZxapjRqQufNfXVTbchbJrGnyuiBu6AMqo
XaSswCad3ONypfvEQiEiV4ryyyA8Sgu2TAP1AZCMcZSUhsDf5+hz10F1M7C7nZW5
zj+flg6vGh8MyTvMCjIoZxuMAmiDJR84u7CBiIakJUruNqpRycSW1//2yly+5QKS
cC6CePfGuKkoT2k6C1WpRzl1qihlemPShvZ9CAgnIaegYlfDD8fEIpB4h/BaxLMV
4WTLQGU9mA45xXmihgmPFn1cYjKBKer/gt7mHSnGZ8/i2gP3qNYdjBr9y6HYS31U
1jB39krc+CGvEVY2gMlVkjRdjBNgU1oYf6ZeNAaW/1J7cjJTO9WMdKePw1KkxIHT
Y3zqw4bfeyB0x6s06kOHZyGiNqe0pLPOT47nxs71Sd4ESlD7vIsXOTP1D63a3Snf
4Ex4YnzScJdP2iwKT1OFApAR/eWz+AoykoVNwvWrVzoKYCpXJUNUS6kE9+ZwOl6z
CL1zbJyIRQhwpyIrVJrkKRAXFCG6faYAJbTo065MuhcqXswLvuoRLm3pZivp9s6/
RfDsiK2yLcA4FF6l2xs5/kLdH/p/59DVb7QwuXgiy0aDdC8Z2t4FPS/kXHORvb7W
nZFGD5xpv8LLK77FXlXc0v60ZI08iXSj99mkmaBn3goRW7MZz//PaFMQ5IdrjX3w
viSlzQxFu6i2RRMm9lyFytyYloYaWS2tONZgAI2ARFqQIDydYeU6Ydx10Rr3JCaL
WMpAXNvnOK8TwQDl9xCzWo6amDSSZ193lf1sObC66K2eRzf/Tl1wc4D/MtK/+fYZ
WBrZGsTV15XtF09zdOfUk2UblUi2hUQFhNtQDa4H2yJZy6EoHfn3vzpx+LJpgZt5
cKmeyzlsm+xUp+APlJlhyXhKTc6myyEyLhN/VNeVBo9njODqK/Nkvp3hY9s/azwP
zDtkIFplHm8Xwel01xhn044RNa2EWM7d5H5jzDi7EgbvKYOYC+7a9Cc/jzIbLoXv
tlP4OgUc2gOjdTDGnNRSe7F9mHIyvf5xUi3v6syBidTUIV1aNDHrLg98U6sqArUm
P91ewtUUADvLfXT4szzH+P16yBoQflUd2H759aqap3Gid79abKBvsjssdMMTe2XR
qETqlGqsaUKsZ9Fd+pkrzLz6wYC+S0prLdUQgAiWNBukw2aCGcENkBZ6q9v0VXUO
WQ6TnMZxIe203LYOnEDDf/06NakRlQU2lZrnDaXVg8V9JSUxcYzMQeCbsqeA6jG2
qZD+3o+Eoeuwyeqgkb6gIStyR0ddI2Yl2o4N/CtNja2yxXjaccBN7Ji4pMm0EBI3
y1Jp9NmfYsUV6xwF7Lnxfmk8MLq6U7sqn1EJhbGnYm5M4i8U3Um+idZg4Q4fk+I8
XwXW+fhvMAcJ5vwTk98dvr25zIjHMh7D5DXpakO+qXk5QNR1j6IAdwbNtjqAzqG9
M65x+5at+P82jUDgyT4B8UmuGxcFO5OmCQrnMTte4CVKB0dLZpAa/IlTBILJBU3Y
yR2P7SzPBbSFEivsTwTf0gVbi+X/GuZ87Ml5x27J2H1aI5YWYLfXuFFlUsE+NixQ
zvyki4bMJgiiP8tS+8wx1OBtgOSzDwj7LCOccmbZMGiCi01S1+AvExoQ4oaYiKhU
sMhwNfS6rQRUcbxBq3iCj9++wwPkMJwLTsghGwpZ8SfacclgnoOpL8peVl5pCM99
HKnuW7OaV8guk906mNzzAX6xL7MKvP6Jg2Hf8MrODSSSSpYCk5K57rFk4nlfR1fZ
nca0EP8oXiimal8SZMUdrQ9llmCPCxmU5wJJOSaA7LKHAoO1CzocY6PsuAVyzAov
YWG51/RP9D7uKbbS07/XgDwvZDD8fu1sYACwyAdinzZ7k77WoNaqlgSvSJko5mg8
F4MK4Z9zJvJGkcYRwPX1E2Bu+tV3eSA7II64kSeVDUasftXczvlVF7qDgGaxsw0f
nCBdsvHSXsphFd9gCfEqh5iOKI7E6pZK1U7wwNC4qYfFm87g6TqAEfH91KCrffID
SSiRuDgqmDh4XIlWdnGx0BbW2dCGumACNpr6mu+XMDxLRXHD5hue3LfR7flG5NNK
QTWVTfUDAszCg/W41cZc4Fi3uQIMq2YvALtVfmZPKnd2a/ATsd5rxhapQPDeCPgG
0nNNNQJqED0QFJFJkyulKTc82N0NJdHqDY9hQ6LyVXlOVJINZZfgi9Xraz2iQsLz
Ug2JpyGmggKVveApKZvGX60avbd5SZK/hhdirCJmde1KqxXkFvEweewW8SLo6+Xs
UkJwsnKfWk5FXyaZN+cLPR53igbnbPlDp7JHKigjI9ehg62jBy9Oss9CJrLaXVnv
d19/Z83QDjQG3WYwkQ/8qBXs/GOaO5xt6yN4hAX7a+43FN3Mh//nUZgSwLgtRv1y
sDWMG8rdg1i+90K2ZLreO2KQIR6We3/AL7hQ90vImOimRf0jT3EI9jjDMHZPcX4c
6ckaXB5VdAVlKscAuEFvrig/qwHsX1YtKEDNmwUGU5Omnc0HtYN1wHAF5q6snPAC
DAfQGxof+lP4X5Wj4Ey+F6aJ9FtdRVJkw82JnZR8Lgz65jbBH/ZsghMltTbLAakY
gSpKJ6lt/V94PivO1mXWibSMVe8LBi+UT7W8SITl0Y67PfCAr253oSvYLjwk+MKE
HIpMuYp9qY39BKWIhgs9zxM3kiKcdZ/N+jEOprzKq4/9QKtjvPVDgRnDyOYgePiQ
RU6KlKp/Rrl9qNl/8eXrp/OqM9v6GCBWHXWIjz42eLCDkUiZYVVipd1579chz9vC
MwkyC2DyfrLjvmpsblbuVKzxWrHFhnt9FvcRbexfQ9V+1RG4fQ4yuQYDu80CdwGN
fmm0uyzUGV3hDXZtEQFU/eoU9JelXA53neqwtI8hfu63FyxfdFyRbMKgobnHtuIT
DACtsGzaQS+GxwGFhyuoNWohczAUypMcqDNmzXvUBAdtT2tUeqJ9pno22IhkpZps
ic3JOF0s0m/GaKesjysY9Qj2qEkJJ5D8EeuNMC8bKAlKI8pvQCMaxOYLNBvDv8Wo
XMqm8IBak39Nw5Xv0PvJSbzxzEJbuMp7dCsNrQLnZTlrhj/i8n4YFIPgltJmSPeI
OEu0vCWiokAeWm+qrI9nL9oJZzTeAq3VRdAWBDcAyzqGyhaD8ayLzOoM5y6yzgql
ytww2B+AcjfCJd55Gz70vv/X/XlwBNk5+FzFncZu8V2m4+DSqrMoT1EJMstTZtGC
oI4ipp0O3Iw+WefJv49xrH25LNC60vaANEcc6hmBzFp+KKN2GxVg58xvrtiuBcKR
GzCj4DxfE4EtwfHRtacIMnWDeXAo2CjFcDAqO8oOLMX0bUSDga+/KZhHs/aG9P0q
1CJqTCtjszjz93IllASuvFgJbpMTrCg1H4tVOe0PL48cJzc2XPd3jrch4TMpzCC6
d1wXZKPd+qJh+9mBwUNpw+QYDYtFf5yYJHy/0mbH9uCIjlc2fy+MIHCgdrTmKiWI
GKUqaE6OiPzMOSZ0goFcfexCpNT0H5OTmNYV55S927taBix+3U/E3W5/LzB8ww74
hJzVvwhan8JNEycQEKKC23VnI4UzE2JXRL3uH6ekAiyTKKRzuQxHAbEFWRR8Itfa
Fk7hUuBeojTFOgyYZV+bArip+q11vmboO/UZ5fT+FR2NtPKr5L9BuxP5egoF7wAE
EUifqZGCg7Y9W1mmpPay7RcSXnPKNl0SoDhbiew2ZTuzVF5RtdH0RIzPNw9YNpbN
esQVIVIzsi65pG/rusKJsGPEkmIo5gBz71qoDzPEsBtEC3cpNMGn/6KpMuwqwE9x
f6eZNN2hEYEkRRMLzgJFf0l5ttwisnkYQX4ZKNeu9K04n6jVpofQzsGuIJPhZ+g5
vtWrn5LV1rf8qgmDN0vLvb+XvdvnSFM+RYvjIHwnVusTZnEARRjvVXS771ed4ZOy
pEpwPDm5AQzAzCVj38FbykFLJC7+ttCHXZJ60lx1p1VWGV1k68wN9NkuMe7i0cXq
cWY800OhY0UBkxL1ylERUxfSH6T6ysWgTXWPb6yBgNcj9Oa1Egw0BKJ3AGaYV/eI
x5zjmt7qp+x/34SenZLqu9eXxDj2kTwnxBGyz/+amq9HGmWfd3JbPzXWd5KWHmKe
mdtWqZVY7q6R/W84PyWCRQ4PxlbgRIcb8YAhMGNgmy3/huFizfW9SiGX5Mbt53qw
94MCL/MQjAObz0nDqNihEDxZV6O40cNuEJCoNxB0LfA4H/Km9siSdiYFzuIk7WPV
E9Gj5eQvz+BXF8Zzwml2fLNkEuczdIi6ep9P77fTWrR3vuJOoCHhN/GopxGkxQAU
aorkdjb68Wo+bXyiF2QRKsUJnTKMi7aEJfDSDmWx2oS++IoxXBq9/HCYpIlRHIrs
zWJht+GP4ZeM0AL1LF6Yi9EwRt/Rdh3duMOnxQBGUjvTkwTNdRfeRGTbs8hGnUVT
WauEO9eSpXQl+ttu+rpbgOh5jFbgFelfgGcQLCWwKelnWUCQXeknIBrhg22n2SfE
m3l82cUpgqDqBCdEpfiZWe3YkceAYdQJBPdCnmLoOQNwtP/wq6YsQOJcZm4vWrYW
1YJftZo4tMCPDrTkLrxSoT4PXhTqdpEUCKG/4mY1fMHEAYUc1KGzwII5sVpTQeIz
idfKUcWc91SiT+nnVMpfP3DMZqSlPAAVN1Ntw8MuZjLaT7XElbE0sdiRoyKaDqMr
pCBX/fxUSKs8epOPRqZZnO0uGRrB9M+Yb2FotODvx13lkRQMrM1C/Q2pA6m2Br2N
arh6XlUYFwKUbQYmw0siD1s3fSLoHq5umPx1oznKFEhG9YIK0yZ0Kl5/WJ52dt+t
l0xTNO1+xOCQXEU7ZxQ64vaF0+fFdpY/9PV+Fxp56zLhSEV2Bi5RfzyLu2N9TT3H
rabzCotv13iqllK6vdqhw99ElKpTtFijR7tPuFS5DY4P4fJX3DLW1pAcWNgOtSfw
0jtb2KKZc5fAsNczTrM9s6M17rG16KQ3cpBoclxfo9PFx39hwv3roHNqMcTVbPCX
8e38zce0yJ89/38djxvMClFejW6YHtwQveMVTEQRtqLwqeGvyD/KuLJhkBz45fmk
bp+stOGmHd+7Th7f/ThfZYELAKm5wxE2jp62XVS9Mx1gUU3yPNeAh/ocDeRSp4zt
UuYJ8t83LOkAXglc5Auh8rzBNGAfg0F7crDu42AweMsWyjhxhTEES2djQV9/7Ts3
03mQW21q4HL+lfMGuT2EDT5szPwU/+yDUNO2hxKom/fx0uYz0py0jYI+ZPbyWCNY
RNGoOv6igbmfnGWX+ydKxOqDR/wdZqH1BGgK3fdcFNhtt03pDwxqnQNZ+1yK+huT
EKjhIfPjViy9E7PJl7sQFsYyzUg4hq1EkMvTJrj1CMzFbtTeUjkuk6UEFzGdVElR
v51Idao2VvcC1K+23UrtvSfXeZnFCABhXBWjoZGAninl0CE+OndgQTA4WxMuCGfY
7hYJR1vSGDd/3E/9oFz4FJCPVuF4y+lUuTr3h2jE7AZDjSUXisHj/ZCMMeXyWdqt
YOAOq57lRBMyIeDO+aNQRy2QGio5PVNWwsZIsi4KAOe0vQHhr3IkHYHLop2WN8MZ
CpYVGSiYKxUcx+EKI9YxsZGttzqBJeAp5/tZhc5G1Z4Qs8KBg6P3HOv/5EDxuMMD
Ic+YJTXwEi5Fm8DYzOb+wB7hdXKWf/+RHY5LRhnaaBW47IBxBQWpZfBztgcnWjkZ
OkB0YQqP2NTSbv16FdtFFpXzxkkUqZoSjZWQHFGkU/h1qOy6/cMO05FWf9Hnny9W
Wf97v5oA5LhX7p60NHzNXiyQM2U1UdvsTM8f1P7itNhxE9as+mm7U4BlFm8OhGiz
urNuIrGowJ5lZ56Jf7IOs/jgz7fvIaz0zPaBRpjqJcH0L1X9YdDyzQmtrFyAYETM
9Xe6hGsxvr/8KL3W9PjxnAwhjjVYDOlkQ1f1TK99PA8ots2gmqb2405Amm1fRbir
TUWp4n9++pfx7HyBD3RDafiv6xF90fKSRGqAHW/XL4MwrGZt8LU+Wm4wK4ylz9LW
mxxt7J1cCUBGyT/XY+R0QwmvwNrYDS3IHF8DZ9gk5/c8fk5cTNgf8y8ZI2ihWdYP
bY/cmd0DeMHDnWIn5TAGoOivzfliyVmQx4pFCuJS7Q7UaaHkvj+RvQ/av5f+AuCc
8lqSQ87Wm7i9jqkyUC7b/XLjksvMcRJGLzfrf5qhKBYFwcwty/4SDD+k/gYSGRKY
pfjZtE6wQc+qyog3kzPat1LAhHJOPJSy0HmtUOcfUNuo7Ue2F4X7YCQkYeCgBuWT
U1GvRUTLh/rClJqyOtt5eyK7ZpR3+/DgoDrsDy2qs+UHDOxskU6tR+nv1hMnAx7q
JTsO1vL0PxHMnnLNakHqrxk88H0Q1ZuuJIiTdGaMCy7pIQNm6KaB98Q8o2RKS2Ur
z8/4cRA9ZLcnuSYrTkDUakjI+TEHiH+3GctTsIEAhEII8XOcU3YtmZi3BEaJj6PX
X8HiHOqGWiwhqMU35go1GerZtRfOlVC8h9b/pW9QVxtR6uto1cC9/aVrIADlvWlH
SHUrLNCZUWQcUK8NqO4kLwduZ6CGf0MVS/bppGilPuECQp/xhxOMZV0pVshsNjZi
OE+PVScG2mhNb+o3Vxc5Yx5txSVT6vJIUrT3Fw+OoXgkYpnHrVFCQRi39CkPogNf
V/gIeFJUPwfNTm+rbyDaJin4sSRfGq8IQNKYhH1lwOpugybjhdPVzZwINl2YYB24
1/TsdeiGCs2aFRonqSMQhrgwJEo7uCA05Gdcb4lcwySjbeXbNwipL8E+brHlrqMY
QQtlW2y0vBvyiF8kOHYmaNlVroLKeJ9hmjHOp7Q+auFZpkE1FF/Hl7ahOxy3sGIy
Gn9dQ0sOALWh0dVjsSRFDrAQ/1HwLf8UdHMJ6mKD9W9kkH65y9ma5JIU909srjT3
/C2+gLgywA8NOnUeVKuLuriqnEJGCdEP66EpKxWV2Ys9TjAX/r+r1SZyIzURLfBV
pPdagARwkUieJTHb46oedEnRzMKDlh9k8JdcvX7HeaVY1BZS5YUeBl5Ba/d0uTz2
HKFsOlclTWYP+NYuTM1KuVE6l+lGa7cGUZyMA2/Xqk3K5ilc562M5/ZVqsIqdaH9
DGXsX13FRVVJ7Tq3AExAHixROdfUdWnMMV65CHDZCmbem0CborVmO56uvd9dLCMX
5NDazXra0umG2eBhbLkh6QG/anBECPxkkyKjB/RVjHjBft/RUK6ZxZhjMbsPUrEE
aijdwa3zEdyTTnVuv2WlFcjzM4v/unfwr0k1/lBjJqBSsoBnYhrW/4PjxeAohvnL
K54kDyM/boSnCWcqkJryCysVuoqWq85KX1y28aKc2yi7DS+PMC/Sjo8lBDxJwYim
RGmhPqlPHwkh8pn8eFMI7ykxyTtvKGKRgDzaKVTVbVZflqThbQyOIbbyuDCePkNM
QvnNMK4DOaKxDPwbA50SDbLZCKH6JDMvKHMmKRB6FOkwZ0QAp9pUOd+Y8w78bHM7
LOkaJtGDBwkyWv1ZKBBhuYJj+O9xXsEg2E7Smbr7i0cCkgAT9p2YCfEANz9pnLNw
BaGTBYqHF5ViFcI/o2tq9PCsYj0twluRv73K3qmfQ26T3DTLZ/JeIQTyO3xHy/WE
cYoj/OVmJf0VfGz7jnJNzqzbTw3Y/G70WARBFfb1Fg+VzH8FpLrhkN0K9CY8fyrW
QHEFXFOCZJdaRsLIKRPUHTxesrZJobaXPdyX+AzyqnGnVpToGBTQ0g7MkjVdg/p6
axJPqdBC0+UCSuh8QbYZQxZno10BsRPZdrh42lf801QSEgJlnsCFlNkhFSxNP70R
7YaWVsqghox59oFhf0KbZNq6D3zWFB7JGhERe6nkFuot7JBaPxzR2jBsTnjWHwXk
+jhE3zbe444VuAy3AqmM6ckjfqcZxh1nbhyux2q8VlU2KMHGNvsloXapB6z0+8FX
AR5EMbiLaDWQqYZAK+PsUck7jPY1Vq9duVf8bscf02q7f7O3nzM1K8hmTXAtS/pA
tnLYY7tSw6P0lQ42VQLXbWTnVHIQcwuizkumwTtO+OSHFTj2Hjlrr1Z2pqhZKw9T
NiOhqH2foK4ted3u1SAERWfuxqaKL+3x6XhlcGxFEnY7dNenDyx8n3E00M2Yg+vr
JDB5RnjyfZ5+y6wSKaDU6UCEO3xmysp1X6WIc/oRzCgvK4WKHdzdKAJaEgQn8/wX
s9rq7XfumI0JSYQJs+A3dPn84EWBH5I1ORDg3A9yItFc7wBFX7UKfuoaaatYijqY
C1/G6rhfw2OQLUrLy2BSNWPf2Yor/liFv9oWoyOTx8YQgGHT4dBB2DHmeuLb5JiC
RwFIoXT8VTQAUqj/3oHTuA5dHrafAxZbo+i2r01JVoouEBDatNWF8Ontbl7h6h5P
R7iFOWVgFvm6amOmIl3LNrUxbxMvn/Z0wLvW7qhxKIMtS5jiEoeYxyc82XDVIcCO
C9CMxlHOcRAZwl3mW8TZWzP7NsRpWKmV7dzUyqq+FKZMIBOMrpdpxLkKrMm/oXko
5a+EAIVJHm78akuEo3bIFitT1AHaidwAkeIikN6FECze5TT+ONUQFa7qOJ/T0LCf
+lLZ5ZSn0Ylxzo6w1M+VHOniSsVFUb6Y57x/79whZdH2azzFghZydyYTOYPFXCZd
csoAdCj9w7ymglSay/NNGgrSvUP/jsXNBn/yeC9zMJ1l2oavHF+DzSXVDrhy7/KG
VlndoZX5HVYxWgB8hHWa1Tp3byRpURe6OGWGZ0+ltPj4dRJG0TvZMXNwnzOanQXF
m4N9cBhxcNiApi6HFYecqd4myGos1VxJ9OP9ohBIhPFnGDtt/E+1xzzJa+c0h5bi
vtw1F8V0k93vd3UJOwozhPGiX76Ga1AI4o0lh+cVSECwUUJrk6j0JxKqj3kKlNIM
v1vMHqxrYzHM9xyUS9wisgz9E9SCEfco0mcr9SkTe8GCf6Cvkl7nj4ldLemVhlR5
cFhLUGYwuml3c8pAlOK//Juq2qeYFwrT6OCLKftGv9KJ26ti2OZQ56DEjUeXlsZY
fJIVAnSP4SYWaOCiuvHsdrhjplWg5YWAdIR3uUUGHn0D1patHDwII2W0SV7vQJOj
MXLY6ivkYiUUAzFN9zDQ6RvsMaYFal/Byo4l/4lCU6nF6pzT20L2fjAw/IoPMR9C
l/q/KGbIeQxbjLIqxfJu/hTzYGAnD+E1IR2KOcru+j9cyVj8UBAoh4u70jtK3RXX
h43zhlNqZLJ6x//+J0BVexxdw/fWE/5jM4kWaBGNYdNudEIgba5OW16aLHapoRRb
LV0tO8W2MoAPu2IdnmUcoCji7LpyftJGbfSJ9J4q31s9RhFK3AjAopDcRGBGwNTR
stVLDiLtVg1qXeCj0pUy1dIChxD08dZ7WpTucyJ2WTwJ+Ctr85uTRW9XsV3baiCd
Afk3dU8SKjnMGqbkmS/V5GTblTiZFeIJ3cV8Begnxx9Rs/CKU6y9ay5/0BraO2U9
/amvkRYFKLZq2o4wlsVNrGa2s86dtq6kUCSk3da91ML1FmLy1r2VNm17+b06VWKi
OunMzuFSeikIgrG87BHyy5qPltCf+afcHgXWq/ypRioZOf5Rtyjb8gwL27cqqB0s
8iopZOplFsVFbd2GlDoCiOuHcvJZ3/7AWfVVqN5byRZjlUavIrNLPZKJS7N+6lbI
xj43i1LxJCfWTacjKneCozyg4S3BFh+p23KybLq8FuKydo5D6DbzWzlNY0LGEYdu
1ZriiSsQMbuM8rHMwlKEV24lf4R7HPvTcc8MDoxlHFQyEo3e7IhWd8krGY7x9J5k
Ci9UF7zjsgURMR3TynxYf4AqNHK6ZR/nSaXOJj4g4iGmwpgB32n1mLw3BupFubsD
kywjUKiXgKxMRM5dx/BAz6UkadFaSbpG9aqhOwHCX6ybTFYYmO0Kll377RhgTEJc
LENnLab5uFdBiBQYKQolzh5G8itNz09Uo91bkMZTd6Uqn63iVTlphv4N2jQAaq4f
UOx8ymyW6wkXk7IVE3MQaXCum58JVH8jLK5Bktg8GMTd/VC38Zevbs2Ws4eNNpYp
ly8bpM7hIaTytrptzOMJ3wMoqAXGqOCv7M7f5kXvMZz0JxJrNEEs1N8AYeynFMyz
OKuKLdfsDuLJzhhWo8rfs4wXy+bl7iOpJt6BxZ4cqKhE2MU2Dyw504vsbfSy3Ykg
d8lJuG8skR5F1C6xPRLp5ooMI7SSN1j7Mdit0WJdirsYs+a5SBebF7jYhO+YqQ8u
FzGKSvOU2OAWVQEY0sgykbrwaYONdI/296IyFEuHsc8qAI61Tx6+o+HdDon85nRg
jm5EYDSqKMZIQJPotUU71H8JiZ/CBU3v7Ci1TgWRxS2o9kHmYWgOLVGBefTRAIuG
GfkHTX1DSbm3ktQVlL5M90l6EteUIumRU9gUnoVYwbXxzSNa4/gwHHrQhpCro+4U
xVkRrv7uM1Q0jL2qf7SPONst0e4PmWzCQGXj4bwYQYV4VWNkeyjXT9//nvOKts90
nsReL+iypui/1+bwko8P68ueC6mhHwVL45tvbdqnKgI9EgvHv0p3rEHsgaN7bKch
5xXOvaAkGTFI/z3YxVRGUeja6cS91/EggrkZhWQA82vw8bsOrbAxH4mFreJZADJB
aaRQu+ETfdqb1u5k6sv3yxI4mjC5dQ1amcDFAtcyKdW6lFmxGUttquRgZ4os2DMb
k0N4C/0ajDesZTkpY2BbPn3wD1qYIdRkhgdxqsyq9SQf/JCMH02RHa3e4isoLb0c
ztccZceZwdZsYR7bKqbJEUlRbZxjUFwoL+i/OQEnb+52IZ9k76xj2U5l9fM6B2tU
Djuqhb8Q7yq1HODSP6/PRPkjNqSk6lNWe48pNMkACvROzMDbFdjw+8deq2Q+F61E
IaWR37ruQqxTuiTkSvA3YObw4u4g/bdDtynGY5LCc6WkB8e8WwHP7Egk2CQlrRTz
W2TiVvBcDDeV/PKo5XhP2PMz098G5KyW82BCs+elmJZbpsZNYSPMjMFuSx2raMA+
uGAPsz0RSW9dOO4gx8Dq2Yu+NxOa1LjNLPe6LuYDVJkxJOfzKkS9D7WfABx8adfX
ZI/DLl85VkWpMlCejegfptLR8h9OHoDtcblERKn7fxwJrb6I30VltQqwtXCMCS/I
u5OhAwwgqHicbf8FBiuPvijgvdwdlSaUvuqyeJs4JDChiau7hd9DBTbj//mYC7jr
h52yP7DNUf1Fshk2uR8I8LxiA/XgLnm6Jmhu0/nYLPo/rAH9sLZOZXABvH02WXgZ
f+4HrVw9myt9dLGnafA4x0+NDaXCzQqikMPL3dE3MzcS3uSHlI75VSWqdIJ5ly0H
8K/x6h5+DPO30l0ePyUQ3luBi7ntk21a+kGYqAfkX+RjomDMznKKB1deZRwCwlZh
RgCt/tGm5Usu8RBh01B4SAKA4/fVnmDVvdb982pLygMIHhmEAqQ4ngbZ+fiiBqk3
g73+rcOwKrRg8TdlHp8zgB7Lfta4gJyRlY2Jjzd9J/JMj8iiRBHSxjXMnLhA1hpt
lbjKsu41rmP3KKy/xkLw5iwEhGo4fXXearRktvoICRW37aotNLQFhe3+ZTbi8IFh
d/aWFwmX+CFREEbxtK5bU53xW0WiFIEklt3Up7erw0zqUfQ4vhrPHDDG10Mc/fAL
PrnOTCQ8fPK+Ccr6FWxnmdbAYgkMEBUVYt9RD7rgl8WVR4RlRc/FvIaIWlaJizEW
36G8JCXFf0uThS8gMwC0a1TPGgCk7XznzUK8DcgnXnWNKfVH2vkJ2GXjnHNGmY/m
xjDMjPCwbodfzF8dANDYKiE0RfqMAxHn95wth5UkL212ks6TJZOAbYQ2TTVwUOHt
bnCrtodA9PddHvEs5NEq1XONWrgiMGdj21atzmXHq1achisTr5cGuLL4FAydPSsZ
wLPiQbDigpS+XTf3B2FG976vZyY87fDv4buWDH+ByAKDFxGHhEX4KPVbg/IWTuhV
eRpyAvpPpRZOtXBstpkdzKfsnbV0/361vgY+VB4Gkn1mKbfncSyr3snCNT0zXDKx
iS4G4UdDRn+LCoNpgeyz/0pdhQpUXto5H0IvbWtPHP70uHn9DFGmqKrhfIRTc1o6
rYDJ/GjHk6YEOJ+AJP0FUb2J9B1vCnOu2cHY4Mp7s7C+CgMbEyi7mCNkAnTRtQTK
jkDK2l3hWGz8yo+AmZp0c5r9OBRSU0xnngCpczyG2VirWGk1xmzgTjbozk/rRJti
Gm71MREtZU+IAHPeD6g4ZUMUpVXJC2oJcR8oZB/0Pb5UkaWgtYw9mgBSNpJWG1o7
NCWum6ynqgpPxM8tdQZJumkH7MfHNEC0trrz+rJoFIUsl45e4hsAXe5fa34oKRTZ
JD0o1PwAeQdO6SCtUlCexzajbpc4phrNozruP9UCm0aE95d1J4+2VFvHNLQqK+Yq
t541kYNrZrIhm/bT2RFvDGTvogFRY2bJzd5t7RXMKZt/pQu9O2iOeJE1YQ4J4m83
E8U1qSdv8quK+V6E7IDWnOUi+KcwH5Ef1rRzPKATNFly0dDV7up9/Wj3kQ/S6diy
2pasnQeVD6K42Zk0BLrKwUOaTBEKbv3cTclaYClTvoORBFirR/hMQzwrhG73V9sg
osEP8QH++vHCa8qdUrPrVU4thJmP370rRqnAp3kwA172w61XvxuC+B6kFkeFxt09
XnrLdu8dIoY0ZpH4PVgeaG4nxF4cGBiiANzyZCL1Me4tPXLZiVfXhGKRfgom3pNK
7K48NCSmIr6f0EGU8wnpV0W8KKMtsCuZ1Sbhyf1SyX2WntZ9R89rEqydQ3Jrd385
1Rg2LSlkX3mCc40HcgIqRMTMwaaLcMLxE7ZZZKRSr6pavqpXmeMymg63mcRnX+Cz
+Fm8wDbyp/RlKI/c4AYq/sGxNYK8LdCye5eqGvJ8C6SAhWzrQB2mm912qJOHGR/5
lQiXStVKzZwN1q6vHYnkuHdVbkDpP8cuvlWtejChsgO5LXDeJXlOUr3CF0gNChdk
x9wdN4LdqtjXhZQ/cb/Zu5hE/r1WwJVPJ/MLDghBhHMC5xhVY3HOgzAJgE8HT/0S
zTlqkvb2Q9wt1dgv6F0y5uTBKFOLJ4NCvvMbYMzxnb/mJXWdz6wWv8sUGzxK0hM2
XzrdM7dZVlnpAoywx1PXg8g3GLBviUxduob3zAK16C33zlWmn2wtQHpnd76KyIcN
unwvMFW9Mj4cPgvxwzuCowN9+g3OFTnXbybJ/jhFa4vMlm2qrO43IWVewLVHQE1t
ADHP/qgLE2l3buEw7eeHaca8/mw1fWKRBAZob/085CWvAp86MMDniHxoZKcugQ4V
WO6HpKXRtqcF6tJEMiUhzqNJEVPl9eFm2Mc8zhpGfTVdVJ8LdjXQdAe9awwLwtRk
vfERwH7WeuTwiZpnDNycaPS18MizLzjCfXsI3VySAKBzPU4Cgrg25qjrOrtZ62p2
AXZQAKkO64AcIO4ixU8Pe2RuHfGJqPmfZq0ZoHqf5hP7eCHQ6MI03Ex1ThW9VxBV
erhB4GscNGoE1AnHHjtehuOgg0XpYcy1e01beMkIrc7TbAixYz61qu+HK8DgINE3
3yztP+B7uIJgWV/qzOJsVKRU9S3yu3iPcC1gsP7hs931L82w4vG7v+k+J4wi+qy1
FLs0oUEjNtjN33ll0KWkAbE0NRduhB/QlJsYY/I0n5/hEwokPYmTZ6LLCD7pYcyy
iRqDF1+xLW9y4xia1h+6DG+UXtGfHFjYZyQRNieNFVB/aOMmULy5xer5nYzbKh5c
H09j2V7iFO4T7qistO3csofY0khd2LF53rWpvYwMwn/hju6O7BY7TV6f+cA9WZtx
b8YNIKUghuKuqnaxbGJKL+9PDS0WLctP0K9JhGq575TIC/K/HCjyeBO2l0bj1laR
OOuTlJoOXWGQFL39e9vdjN2w0crzDhUvVbeUBitmEc0ZjEg1No5PPN785ZEjhZlp
Ln7DWHQYSl47dAqZWw0Mt/WSJCUQWa8cYSv5DO/GqeixveUYrJwn5osiois7P1Of
IR8rdSmliDysQePvyg8kWvlgVCkX7jHluZE9Gx3CZ2R0gJ3EJzC40t+XQlLBF3u+
8z0aGOxETIUl0Op72MFWKkxzJxKYvuHWtEZuvN7cdSVBxvQEE3B69ypjXXfwZ0od
bIS1zvLJ0jjrBrdYZMtRtQDWYS5x1uZUXYIzrzQiSe/h5BDL95U4fRoV8LDb7vP/
d/ltrrj2ovF5h7fS5OnsjGcIFXl3G572s0tUi+gAHeV8+80VHsO9TxO/be3lHYgC
bYAR/kV8piXvKdOQH8zbv2GBQBn/vX/aLMqTdUqu/up2Bs1Qr8Nwztl8ADZSx8Z3
FS34IjB1xp04v0kjelekDNthEYyLkvVVS339Jl7g2vsXXbDVTAB6qSaO7SD1UEAX
ttXx0jU8zimNNx2kwslUKYa1rTjXJBfa7SN5kcqD87fZh1Ldy5pfp7uuLQM9UUUV
irb3u8YhHOcOMo1IL2704hpGn3TuojqSnzohR+99bQIgudfyhtB6vmVw8uyo9N4E
QqDWPD2IMEaornC7oNs4YSbyu6wEBIvK4buyEItENPD0EYIxbQNxcYnZ3zNogE8Q
8QUMOcZqRTptzBPiZpIqs/XO3iMJmwg/MAKesN/ZHivim346/rY3mPaollvxWDvX
OyYSmigHl5eNgXUJsLtmPUpXNGpykaD0T2nc4W80nF3vF79auQA3uvCiqkWEsZPu
wrZx3rxFhuuC1ty+5WYBkycvUYvg6FwDBrXOlmuVmU5cn7gOAZgR53messI77VYh
y1m1EPMSmhkl7PpWksTrtIp9VDrqrPnEzIvAH/eXhsMcFfEO1BGUvTc0h96SndYU
D2BUwra9MvUgmzOA1OW6h9gIi4VHiSJlHuwfttOfhmYtwABcTC2ErtSa8YHwIu8y
F7foYrNrfvvWFVHNFTyvP7085B6fp8QUTbIxjIaueOS1ZkaPxcHBekbwjmBnWKFg
L3LNq8cW6PaIFFVM+R6gPqHJGbtYRCiNmqFHLlPoK5hfkeJGRWktwYHQZ+KBTiVj
29apyRr21bYpnIF3fjJkzztvsYjq5OPSiPWxWygevRagw2uKU6Z9n/nRpKq8EueP
Efg1MXf+7W1MfBnjqTfPIkLV8O+sKH7uKld12KfmCTr8oyVDZZBsQ2nm+vGL3qhr
ARPJlCFJCayBwS40sdiqFcD7+q3yrDLBnmQPUbtR2eL47U71T6mBT5X+IwhG6cVx
3yjd7s3zLnA0y7bIHpbQ/pQCyue6muqTsOOwxUCyElAFHwxXnLf2a89WSlf6y/rx
6sASaMToSD1/aTISqGlfYePlaw9Rv4mWDV5CEgpSv6Xjc4otbJinr1e+VOcfYzmz
ZlzsP9xrM9MeG9ySjlo4eOoEI6joMcXItxbKLXjmKf7Hw9Q+9JtPa2ygFtJONkYm
ck2TG5tPiN/q/X+/LXxAkw3vqOJnniZm8z8mRqoC8jrEIkwGpEI4nfjXR/eeJlWt
4t5I4xi+n8p7tLVaqvr11kENvmidV4oWUJAOmipSarpIztA+0h7zTvjzK9mJSj7T
cZtFpdiWf2d+C3OZtNvBYEY+5NWP8aRMSTL5FjPIz1PW6k92/yhp+PB4CVwDhoq7
fKguxZ6yo+Zwo0fe/rY94k3vC+5eyb2NIaSVB72nlALe/3HSU81aLXZlSEYLC7AP
zb5kW8aAJzuTKSfdrVbPP7VrXeLnxgsIZu9qCqqj2HQcNlNucwcmsa/1XjQyOqiz
qOzjTnbOK3vaDOHIvDgvnHqrl0Bhe7XNSkm3S0Otyt+dYIpTTQYdSl6SqSc/4Wry
VC3uoXVvcv7bHo0CEw+SQnTZnBIiGfztiOXfXq/ufSy+3OQaBakDA2SJ/N0EdwHg
m7SbOyPyWsQdgdQBjkz82ZhVJMTli/BZn+ZXR72nGNK3AmSptqBeAj6ZNUlNlb3e
mg7oj7VWJ9sttakCcQlizFzPdiJsOLI/EWSWyH5Lz/TFX0JWIZ3Oh98ESafI+s42
tRUs7u0387fC3BR0pMYtngB2M8bQTp8MJyZJZLsXelXdq3N8yNZ+Nffc8jALT16O
bewJwP/sfSaWv/T1s0emBv71PUar8aCXZh81A41qlxYp+1qoSAFvTzLAnJpypj2E
tMxaeUIsp/iTc9vGUzSVwu6XLB2GrWNIHnxFuW/6dW/XSxg1j09iWvvyQS9VRa49
sbIe2+8joPbWQo7FzPIKxLOf7YzBufZNuMMyv3/Tjf1YBC5V0Zk/njKg4JOenpFD
66rLrDWXCxleZ/1tCjH2Mb9haBE7hhfR5nyZbkrgy3Sv/7By1xC0Ng+sHrA/19zk
MAjZeqCnKTHTd2vCcPEGTeeQHj0i6L+g34Eoips/m9z/2CDcQcMiA9Bct5dCHlSy
fG0AGFAqdUDVk5cX+eYHQQ==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FPxlUY7isgLcu7g/B36Z1rOOpeXvz2UriP+aVh9WigVOmE9/F9eGCqNIq/NtEPai
CloZFaK7WwA460QHt9L4iA3c+90WE4/5yzv8ldmn0FekPWpOrri5N0o0DGD4uLYm
vETWwSZhEKMsHG/yinOZBMviwkLHxTbh90CKcDNYdRruLNNg1o4z3/o0YwpguQBc
e//JU6+Ctpxj+/LlROvW78i0+uB3tENbGkXzW2IcLXfCBLtQEw52MQiIiBH6tU5N
C5mDB6BIQ7VrKerPQa4RJtiYo6nUviaaJz7NvGCTG07QpbWphHDC9NhKvKAeCs+g
ivyxbVz609EklbbGtY24Kw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15856 )
`pragma protect data_block
YGi1fiIZpHBzB+MDAb3/90MHqirkxNitzrNCAB5SMfMVyR7iGVpSTe+MvijFIHf3
NSv2XHLq4wO0/89mKu9YQv+BGuTiuQYgKVzfm66ZrPC6VXRtDVmkfNfoeebtfMHR
ZzWalHfrUA3P8BEi3pswrwitmGcGpMx0fPO6Ys6oHGmxy3RtfBPewtQJs+QFhC8i
7+a6sli3L9VAySEKCKF8rS9hcAun2EKLTncJlJBYSL8ct9lnB9iXAxRLARkNvyLB
AdAWvCpr4ugGwrEIQROm3xVI+AaWa23xGiHhEs+uH4eOQVqbx4wmYcIMOM6r9vKY
E0V7zL327J5HYUFqbIZfr9iJnTk97GWzvuowF0X57W0hk/5wMmOJSHkMLKyWhYci
WquF0Ll9FXWAqecFLyicnxTUijsr76b4iTaZBmQKgO8dD41B+UfAKmrZYs97+2uR
4DldyoQoxr0yE3AqQsmLdJSFeXeD/gbkFhKanDizC6e+yFaqWGixtoijDM1mUIpa
Nf2KWa0XoNFegCpcFb0NjBC/YCCd6c5LmZ++AwKf+r+nKEcaEq8dVU6MEuxcB0Rw
+F/TrNaAGaB7oqB6Sp1ph8DR3frDULtdC39Nely52syy7wdM+IK5GVWzHCm4cXmZ
OsOOgOLc4K0beiHDADK8diAiyh8X1Pkmnli/1N1vyNr8HBlVffl6ibX7u/CfZzdV
NAJz6qSFUKxKr61fp4HeJIpKG4zlsVaGwEyqtBcp0LphhtWC9MPHj9JYw/c8SsQ3
DiPJxgHCpzL5cFdcP9aZodltTOhcw6FZ8L0AdKh249112rPKrQYXHbfnrpePcU3b
keAViqNqxDNIbAg3dPkCUNKnNnQuYTfEm75tZEDO6mgRzfkRi3q4ls32U1HDVFvX
HGpTyKLRmLxE985X2bBhBHm4NAGjQzjYEkOlhfwixSec/DqxOVkpUPkgnU0dRciJ
lS6nbItbA60fk/Apl1FM9/11uns5l1AXEkHMo6MctKY/D9QkjkJcMytt4ho024Va
zVWVEvLK+wVTENupyPidDhlY7qrWLmpt+eUOjD7r8mioj+QGaGnYRA4C5/8lHs0b
Zs7KPFfSFqf4UjO2QgGrYtnKELuFipsjlrYbe6RH5pBVKSN6mz4xVMTBxYDuq4WQ
rF/AyPHL09f5vtT8jZUKEVPsVqkjIqPrtgmAbA9tCRl3U+/27jPngoAaBuo5SA3/
bgsiqU+oa7LQId3SwhmAAr1OyzzlWxx+D5A8nHcqKMe0BZcT+A8pFYChkJ3z4hWf
99iHgBjSg+MU/6ZqqDbMkaNmafHWX0/SfuJVihvRj4ysS93oM8U4uPGn92EYbEOu
iQViW24polHLYfGL68Sb+G4yBFC1OgV0DkNXAWQyJogUszNO3GVvPJ1b3u8yfX2R
E9RSZF59zeTjECwMJedklhjyAKLaBqEYidP0r+juaSi+0DQVOWkJuDV/CP/9s++6
lR1Nt6j7w/ssr5IIi5uS44CTHLb7DCpERAvLugC92Pi0SfGJwGiBoBojL3ppUy26
ac7Z4+9P+OUbXiC2gIkK1OWBVhxvmYlM+Z4jVSCz/hMCr2NupHRBfCjmiS1iNO3J
GuNIjvtrG1rsKdcwYLkL+gSLfHPYiBKXBIq8sIM0S0PSX0XYH9fuCG7W5vff0sCW
RyjYSrr9P9kCb4EwaIPF+0RJlgi6KrUMgNBfFMmj5/KKsMheDOisWu8lwg1PDg54
Zs28PSukqKUTFl1QkUYnzZiUt36GNL63g0JQWlz6JyOUqkQzqqi+yw3tbKtmpPTA
bu6rwdjBUSLB23HptCTJDrcEatzaRDPNxs/S0C2VeBeARiagHg+7jZNkEDTV3rkM
tA75uYBNg5WOoZTrCE1Z6pJ5e9pHLOqefzOzcYJKhlQc/lNV4k9HGb7vvry2DU04
QGVJ2wEZUHwBq3JkOiy+exMJC4rb4JSkwCvbytAGd87bDpeP78LO/Jjt70ZLsxZW
nrD+I6uVyd/ZVchGH+mi+RdkwKryArjArSXozaaRvQtfoYzIRRhz3ZjinDfvf3tK
07IGkSUHJgX3e/wCTM61lCsEvHQ5yb2WSaOsObHAWlASltqYkYaqnGfarjuIH9Lm
sbkqvyat7JYMht6zzrZ+kCF5vd6wHLOXYEUaRPxIBDzdhw742x6c/lveoRmxY8pC
Ol3RNQEIbTtm7R2HcXyg1I+HgQxpd7/12TvgDuHtiWRWg1vqi4J9V7iTuwrGkKzs
wgsVUp0uiLJc0kBErHQVEw1XnSiNcP6MfpEcYh89EFWu6+fg6x5DrkAgAzhr/4TF
QugOsfbczklE/fLQWLAy6yubnq+a2DJP9alr3CQUGXOvyrtpnmx+oprbC0XXXRjO
1+bemw6hYxdtYg+7gsxcQUHbQ0fw2eeIli2jitee/oe/gw/ZzIKwD35VFXfB8ESn
3Kg7I2DuZp6J7iaKuCqmOdXRnwiQJ9nolQph7SdFUsIJgD3S7Vcu4f17LmP4/vVK
n150AJ+CT2Z5TtpqT87/MVGZa9KOTEuVWpy6lvd4Xw3ezc+OBE8JGvSJ4gJHOeNS
UJcBvFw+OWwdOu7usG0HSNTPL9Fl/vyCinelKZ3dSKwkSv1yhMek9GASiLa1SuyB
Wio1COnAiVVOxM6Y2j+Y37mQ+7f2V+tml80QdBLXhyLJ/XOAlsLVyc2dYKv1Fvdw
Z1sxVwPFplGw+EsT0aCYNaSZnrF4AYWLVoO2vpSKinybbNUgBSxai+wp6Nid20Zj
ZRy4vl/adT4eLg+sAPxZiO6UOh/P2b/C4lbdtUMmKWz2LoHfhbAGZ8LAXaML2Au4
w3Ao9GVeTAfCznQ6MtSoLnJbZKJamdha9Pp67WgAux7e3c35UUBkXX0l8YUXYvyq
MCm3gJuveL1SeYuvNGoBOl15R+0tLibJaAwDD/vaJfAyQACvqITYMUk2z/GjSKf8
qB7WsluKMdzANsBDWomCIEQBP8Ud6JndDWZiX/D/G6U4A6N2dpv0xMnWDlGswVsu
UhC2DF5VB9qBgymCZ/kLVUES6xpO6fHy9qhHf0QiiqxTHzkPBfNCnRwyJSij0X1U
CEdZ2L1XTKAwJTa44/y9BIdVnyCPxWu9t14H4oy26crz5mD71oMYFTY+JE1ozWI+
2tyFZm3P+64aNkjqcMEu/x7dslTbTbHL4PBO7G1xYzuJa0Ld7prU+NFJF4J2Tjhe
AfbDWzKm2tcZq144/tO5d8P3esaLcom6KPglq5aeaF0XykrJPUaucopIyJJ82cKl
1KKggk86zpQ+5f2WCyNbk9H8dp92ENrkwAWQEMVh4jFWnRSZHX6+VPLH2ltfONp0
j8as4CPf4ouz3EH3bJlqo16DzuGEr2bWd4/hPbVAK1BL9KEJgqdxZC8o3qWg8lqf
UYQI7VeVLkfuNPfdQnYokOGF8ikFNdAj1sQgFKiY+EGbwnXmuk0tk2FCFEkJvWEw
ntkkXoRZcsE0v6qHbWrlqxdA9I7XyhZlEk/cU4K7TM5URhdkKjxcYyGAyaZbZ/W1
mbsIIUjhP5+pMDEpxDXcI5137rQK4+CdvH1OrDzZAuhDiYucLKT+irvRy4uqHwMU
Q8jikL5BC+8QZw4NBe6T/AwarQI2ZqoWED35DixQkjq92pmAVQ5blleXmnd8+5BZ
ZNqzRr/POBIejT5b/68teBf8w4Newo5KMLxU8Oxbt3oBfIxcJrzPXcqFXO55aifQ
Z/sKKggBlFsgG+dIAYTWCbb5qwheQ+5RRVyiexa6CE06xS+R6ZvmX0M7H3N1w2bw
O9/0wTozI7/ze2M3GGA/VpZq7EjGgaOQmLyxXSfoDcjA6jvUl1F6FoPXkSnMVVAE
FJsZYpu55KEtV1nAYeklS2OTigto565WPquTJEBvDSBTmBvxe/XHlm3LqKcas/ct
DGD85QAAtyq5kBOUdE+fYORVNe5gwL2+idOESaBk28heRZveaFTIv/elOmnZ3hLz
1NISRCcH8onoBnMsqFTQlFXsfnfU6wiEYdChVfphUWMdXxUHecLgtHnXORpacAfz
E6yPiqLv06RVt5LsoW3Lpjn2zxV+5Z2kiwGpe7JpGM440p12IU4wtuY75Ak5KWkZ
QvsXv1OxV3knlizz0CoybEc6dmPmWyo/Gwg1fQjI0Ng/TAUzjd55anuy89AOebd4
hdwkexfrWasiV0L3XxXGmexReQFlGqraG+u4eI7nFKIMRJEcwWkzr5sgpPO5UCB9
uZDeNhMkV8evjTfpd9MNUI2hzNM+iKbVRy1K7dAhjXa9Hwff4LTJWlUDKP/k7XmW
DqI4wZCW9O5VPowXwnFu3MWro2L4oplmw6wuONmxm/w7FhDH1JIDiCFw24p5m9WB
+WiCbqH4RcXQdYEpdKy97T4PcO3DCJuK4ihR6XtUQvAH7QZjWq9MnfqsP2ro0H8Q
WFlWsmYei9LqLC+RdgIvRwweCmNDswPJNRu1NilElxCip9zFPeMvuchceFISN3U7
VqIhuG/EOAg9pydMlLAFzKjbikrQMJ6pIrfpTfK2gh2Za9gU75a7L5ckh8Xmqj8O
/6OSc0ZmnymIpEDc894vOm8Ng+fnZfCIUV0MZJ+6Ng+OL2qur6nT86nQeCdHhpjT
JUGJR79EL8ryhqagL0dqoni6oosMrp8esCCqWSttpxGcRXofRj3gImWjVAZhCq8w
TB8EaDnPvbV4PiSFqcK87uR8+Ncy5NDQ3f8JvtvSGNAoQileJ11cTG6AkPdY157q
ZfMkat6KHNjUPP6IJfl8WrxPvG6MTLttbhKgulL22Eh+/O9ESDaVw08jmZQmqThz
QSzbGDEDuPYcCk/IAK/RelcHYdTVYVS3NvaqBQ2u6QTv8Ou2U2oV6NpU08p3lrfd
/BXBaTWhItlNVWT/oQGLD6JhvIYsrG3yb+wXR0rCZo07g70tsqy9LNL911knSvtd
B9RB9viY53YLB8jRfcobPu8TTNXL20VCPYYtvCjVlvIXcDVko6sLHkVCC6DS+iYp
di5XxSQDC0dlBn0aTHs4ULyS0oadXn08uLpFLWqmmwLrYmJeft5iOGmzHp+jpRi7
wn4lmtDHk6xCmtJSpnJV1dZUOV/VRFSJmyjrCfi27aBLWAyY4ZFLuPYrKQfTK7EN
lsU+nfeMv6MbpycKpkaHd92PhyK/7lD+yg5TL1OXMYj34EhA57ZBQqamf7w4hFmD
iMn8QwRo21Kt+tvzp+HrkM/YoB7r0sTfLGwpApb8MLr87BYxSsUTMEhOVPk8KDNc
Q14PROAKnV4bynWSpDPGU7TsbzCtuiAczrVJgRfmQihiOwfF2M7HaoyTIr/fokNI
u2PMLLxroqPcDhe2evktk095nZ9pZsLHbkUQj6fx4KhFqmNrtrwX0YDyMNyhUJhl
nPWVh5gXHIAL2G5ROtaDKwKrbAV7qu2NY2x2X6LrsotQVh7GgMB9T1yKQceZQC//
9JTw/gNBLJddFfeNysDR2y7GfZczAd03RMpSXvDsjS7RVJayW9VaN09neo+9vXGb
7fKcuRYoO+vYK6hq678meGXmS0HvhlLKGqtQUK9C0tNF/yD8/xaNx9L6m0dKtDVJ
sNuefju79iROt8iAQoCDn7pQYDcyPnfN3VXe469guKKfKJ1MWZmWrEAF9vEI/kqc
lXFBVxeWaUj5aACFikB02K1ekFuqG3ursYO4q5+eHgfqXMGXrZ9lgx8whxDVSHSz
Rk2R9m469a99c8c6CZTgOYRDORdql8TQ3lpOQ5dwg8yv0UO2CIIp3RjS6XBtM61Z
50s2QWn4hmLLiMq/LtUm6aIRTYW56/7COmgDos/tIgrGQIafc9c41uX+bXEXZ8vl
eaBmaxXV09HX+GkxDq6Zoa4tjIYbadKi8Rpi4zz3BfSwDpTG92QO6DlbAP/PmX+O
xfzu5dRuNvVYWpK6GqAYZYxENbj1bKtxP1ei1AB5dfZaRd+MCc92a/OgBgiIuSBJ
oPC7RT6MkY8wgMm7ZefJYGg3+dZ1QvNP6R+4fFHHr1nTSAcvr8XelM17iKB0tKHk
2OdpNDczSn0J5DGEBl1lXAr7Yg6HBFWesGiWlZUjx5qwOW/+SIKbWmTwD4F5YgyR
cqj3BmEL6mAizu8sY66YvfQQfcMbuQYCslmWzvsUx0Mz96mndurGOz1xV39QMfPK
79OV/m7X3ZuHYFY/+8pdUkC5UipHCkkGPp6/ikYQxTbv0rPMQUfKr+xsk5N1MR3X
+V9HRkLH6gxK86VvIydElAoX3839zhf3vmVhnZdeB3x8yfjYmxsp1azcARdCCtDQ
/Z/2VG6kNzTZOtNkM/M2PHeIdGhb+Fe05kzFlDf6tNJ4vm2N4TbyUNpQgYY6zwyw
Jg6XB89FMo7JbBp/q9e7YlFSLYoYCgSwjMRUKaIr+FW+Dmjp/mEeeOyE96rn8PXL
IhLVCNTRTwa5LEGVCtKTQyH68ZcecT1QYt0RHDH6okdvkVbXL3B71NQAqOs4+I7f
0IrTHJVFCyD0rSlBZJOWAMo7mdnxKFTJw5Dcr2lSWB8gfpXrjl4a/KdxL9omeHEt
6dyP9LYqNGWSpvxziLjSsZmPcCnge9nSrerotRn7ZOe37YmK2sybTJuy0ujdLIFX
McsCin0y69I69BQKP3ceuy7PFgxHV2BTeWjX4QU4kySxw1XjCeBdYyHDtpL9dTQZ
O+kMfVIWVTDKLxhR+CB6XBzS+JwQgALezDlUZoVY47C5/OGbJCkCGy+CajFdiE6T
xM8tZCSUugTI2wyrdwO9VBXkFmQt1dH0XQGyecFKKv9Nz9tqUSWP1ZWSVuJAef2d
z6Bl3twInHmpkyq0SIliN5Z4/PEXyELq7O1gd/EHYIwhtqJXsl/6xUEeAyncezld
lhT7OqzgPPZ0gWFqXxiOyWnnGLeBmBjF9fJqjnnTgya4i2mxOoXNHZXWyiqJmZts
5e4aY/TH+Aq+0qo4RVaiuTHXW7OyHUDUeRWpuyBpBnzpCU7qm1QzFkpNYdyxQHdx
o77gOrrzXx3k6qn+BR8Ny8XnYPR5vuU++4FoV311Hx5mHqwnlUF2PTY+0FheYuHo
3PxYKbr8eX4nu2PEZACLMaOAWkHfeuZPDm54Wngcl4TzGgz3eTY/Ek6SROXaSiAq
vBECmYFSHnZbdTtU3Z1mTuAXZXBvH8FHozDvEY++uMhvrRydm0gx6rrykZTFpDt2
d86P5QNVgjqe7DvJJ/5GwjgP29p9jKa2Vco7vgfpNsfcbzca/pFhQFp6Bxq8SKD6
i2VrgyqIu4Pq4YubuB6gXLFEBnYTooXlh5XLszMt1nN8o7VML+/3Fe0mAyX6a2ab
8eXObiFQ14Q4En2BvgvEEn6dtAasIvUIScSu1zsnFn+gk4ie6/ZEGzKWhX1gg9Kl
ClyXIpTiZqUFP+ZgQhizspgZRrp4/CWWV0LoGOJxfnU8EV069NHoPbFDV9ivUCaP
jMt8nUYNEFeHL5LxYg1G33Tutf1R0t8nRjaltwmWotCQnJMVhCzBFkFWyULJQV20
YgtCD/VCfRH5NdHRKuEpkXPDUkR7zGS9K+ScvYc2sKx19dNn16r7QX66e6Jw085/
cF/hn/2MzWMetKpwIspE+948M7qL7QmpZFXQAiN0mYJWhPOYqfZdXzgesKgJ+Lau
LJudxBfxLoJGMXBsIDVSWw9GoA2y6j7Xkw/H2PB0KEkU53USOGTCPdkQIX35KUZR
3NiSBCVkcvB0CbQOGKAhcn8Ivx8JhGIQCuRdEb9G2APJ4avDLih3omd7PGicWnl9
ZhOIdpsqloKxbSdrGj3IoUFh+AW8zZUdSaDRGI1d4Ft7RKxYAPpgzG5OA6mnJuuC
o2guK76LIMAuKqmIXlkPY2/tbylEhXHWmXt0OvNhGfxfN3z0ab8KA1I6RduRw8lv
RqaUgPIJsabSXXJCaC3GVNQGub9awPV6T5zXRhv4HVrcXDgwxEkaS59AXMWs8tbX
SS6icbEr54hovAKlYpUbI1A82qvhFZKjC3BCn4fyaNKg/YTvi8UYpVIC/QF8M4At
t1bEJizfeUjTgAqkOzRZclHzSmKzTR6ZXJCVyB4UPyDeuSt2WA5jiUzSOsiwRyd6
010qS+x+oi1P6Wsq5NM/fzsdEMzOjNYXvkaOgMTuA81l+gs9v/JRfS4sSTPkGuvw
npuBOPUvHdHe2v7LMfEMCPCNuAd7LOuO7QnP1XfiYZOwTxRG558lSAeojswlodJV
vmCHwa8LGs9pWufxn2tO9RtvbUU5QqHzAZaHooYTM86/YRJHe4m2cyL6sclFtHOg
/kxEgBsmJak/0I0jHc2D5MUd9ekXsqfbwqOfz9V0YBspNJu71KDI6uk19A/HIYi/
m3it9j/P8eLZe3fRo4XcOpnTvhol+fXMCRZSz3C9KdduHZIdDjGgKj+OtKhIbZ+A
aG0qYwAVaYUjZZjUH1lUxX9WJqckHI9d0HlMqKHozVfgxa5iPLBQRjjUuK4A6EiE
Vnd5o1hBwxPOUvdp9JXo+KeFNA73y1IkFQlIDPr+mnMwju6Xf7Je7YWbJ0ifulnY
TxF7sPHPLrEhf1uYw2ZfYcUvNwoDpDFMHj8qi2gze/JgqmXvfiRZQxtp9XyjvkLX
5NDZ2O0/2k0K1U1eUihvPKUO+Nubn5d9EXwr3Bg+xWvp0CzHqiHB5VWJFNkdb85x
C8BdlFmOiPytdVokkwQLnexOsZZ17rWW+lyegNocnE+RXNI9MZY6I2WFOqLAjhfp
5dXQJ1/U7lJ9acq6gI+USNz2rvq9iVsAjTxU8sp2B/UDtvxsMk7eljYxfQL6v86/
ZWCcPadfU9fhPEJF7msA467RODuuIGwxDygLHt9OXvbkCy4EqhCxgFScxZ0C2EgO
lTx5jVT8zl3cviB6gkswxbsYjPTaz8vR8p8Qi7OZnE7Xl2M6tiIoDrmRhL2tgkA7
3INPdDe2aouaGm255QGCG4Qw9grjdr+ukPMmeiv1Lx57fusZpz7HoeoBiM5Ug73C
LeOxlKa3mhdYovTBhMgKhqwDbulxjgQ2Yd/T9JSB/k0CfiQWjDnmZF7xCjYk9QS+
kFv9nXqU3FFg55MvzHj64zl6dcOcITEpmG5wdBwU7ZG0eLRp9r8S/+0HoNCB9ioC
4/Z2j0noM7UlycStVOHxMQHP5YvBf3ujC3MdWLwqZdIzz5zcxhuGi18X+J9v5TJ7
IfSg0TrcM10IIylgxH7fcYK0FQs7gDndcg9z2Ai52yWx0Cbs8pM3nkMAk7XLu7Ja
sLnlYUwSvEiCeDQWZpjgHOnY8zdNrkf7xnYGDsTSI01oR62vo++DHDFCjRIwfkqY
HAnZpKrtnvFZ/0ooMxVmBxIgJ4uUG1rzZGS5vdFm33R+1dVhudsbdhWykEuYGpj2
ADNyx6cqLFDeF7FtV1tBKrFXx4hhLzRQSPuA4JiV7aCkJusttSFt6c0ABmRZUfFt
OHykN7aRjBAH1ByzMVWTVVgJ4O72rT7BHCyjKG7FWOXt0KG+eQ/D7T4+sY/dKk3s
SCqI1rpqGyMMCQEqqJ32Oq3OSvgTPVt2namHS6ZifzmtGLev41D2wfyDq8corynJ
J9QrYS4yaYlL65EFmjErRr2nnFOtbATqeZ8KdWBfzyNs8+159DqcRn9bc+Lj2mz0
58JXbWWhaZHsAKj+PsOG75qOhCSZvjhpkY3oM3uHVqdqqdnNbU9JCn1OtICqZqMg
ZjWlYLP4bkcYzEMQW2nlFWmWR9okUeUZdY7UPggf7s5bs7n1LR5GwLUuAHxB5IX6
nrMyLZzwrEN/Dm9sxMzIb6cs4U3xeRGQ99FoZ7GGYW6zI3dgQdAmK7ulr+agCvt5
ItvQTEeDla569VoQhm7CRfgbWyhvk/akOYberCfk4N/JoHScgDL6RmNQRY2QMaZu
7jL+hnhVnw0JFr6gHSMofWmEm+ylDrBbYJbNtwiIhQ+pAZshHcYk0nNsXvoAyCpG
ESDsvX/slAYq6OZ/xaUrbb+A2h2+p4TBVK7Fk5K3ndR0TUqH49ClmYJ2RV06TZLE
BI0/loZ5SyCXEEB2D8e4oZj/7Z36mbwn826JjGMshCbl1b56MPuNvN3kZmKqWMkV
fSCCO2HErFEnwcqP+DAgJlYIsSztahDpwlD5MXYIVPj5MnSy/Dsg1126H+HQGPC/
ZES+z0hNsSDgUm/4h1fLoC5E538ekGHzrGKXY7pK6ytr7AmketySAE7HRzPuoKVt
1FCgOUlgSCquPWZ+PoxvGwkXq5IgLHC4TaUTemoClkGB8vpUJUrf6EqpEgiGHfjF
WGSx/JlCcVX1XYHs7bc7oduXs5pgZOkKlslIZnJtPWLWNYUNA8Yi55Kl6f5yNeqs
gXQVtpXlrnuQJPdDgXAnNNM1wufEVMTTFTYnOfL9JXtosnlrdK2j6urYJDEecR/C
C/GP7xhQnRXG9elmiSayuRMCsyTT4oiTON8BtTHPe/UJvMn69nWU4pbBjycFsAjg
40C0gUf24NzvZrSPF+dQa3fq40vN331YoFDSYKSpKDOb4xk5pRMkukbQNZvcoS9M
uKSfZAv7VHFa0npnXcvZnFIoX24qZ6FjTQ0x1UZ5ujqju3y85UdV9yULz71sHfmz
Xu+sEEHVVdghOOBErysslCRhnmHf7Bph52X3QNv1hyhqELIKcCbhDtLOjuM4MPkr
Wz/0NFgAUrRv7UNoGbYxPz5rtk1ovdZG6K5siEcHVU4S3tVU8t4cjIW8VqpgiYg6
y2sX+vRkbkcppkmlRdzZifYFkBBgJ8COT/a+yZY8DfLaeAHlBIWSJAZKo3wRaNm+
/Libzz49o8eA2yYthv3rVrC6cbYv7LRgqBDbd+1OCMEoM/HkL7COUgx6X8qKNS4Z
Zg0EfwAcTqYO12r9XqBik0H4cO77qqQzdRRL4dNKtup8Hz4xWPdcl+R2DWvuN6Eb
M27g1cunmGC3pba021i2DjgvAcvALnOziM0EU6wjDhTNLAVBGsiDo7r4UqEAddYv
OrWZbJTcW8VdxWAuy+qTRnHxXBOsta86JnkOlUa58H2DBfTY1BLL27FEKbw7Ugjh
JZLBYn1HrXt2dGNOYTs/2tigSeWGy/6TL25OPMME+t/R0X+Xd0ocblD2Ph/aPv4B
7Ca3o7SOP3NkLMhi2ByygxOIak2qoZs7Yct0gcUq31+I2fUc6/I3oNNU9QfkofJw
WhI/wYAvgwDltMu9U0iNLA0Ry7XS4jPLAvNah3lHVSNXt2se5Y8oeDophy3Vx4Jb
xv+HAVx5+aDU6HURWoK/fW9UL/okegc4+RDVnHPq0IRvKE1zSsxknHwBxnlz5aov
VU8LPcPfsCbBsJLyfxhH92Nuq9gLQkDUg4QD9FmwfxebLLZiZIZ6SKlfUbOC6BEk
+wa1Ac5Vy4QBveVUNSVIo0Qw1WdP8G1XrIUtKgxbCNldCQZlG2vK75YUe8BAOkNV
cc5QoM+uVWGCWeKKbhyXC0CAL83tAFybEPJUWq7e6ZC6AwnTNM4NopTXNMabYV4r
VoWd5DMYfio/80ExgTr8DU6AZHPxat3XWuwUgcIcNLh2CBLDkhuPhVvx4ncJ2HiB
tHwoPNlWtmV8BRCIOif2wvzLnjVGIW4DJER/p0rL1Imn+rjm6gMW3UkcfzNYUxw/
8rGjoxPmfKEqO6FE02tgtFupMPsI9lEu5MLw1mdIQudlwrxxfxp9Nq0q4WsfdN3d
GwTXBR8LLRyhycLEFVcdii1h08WFbIvE9AiRqc7dfXwFDavqXuFWTTe/A7Svk1sR
iK1qqeKi7y9JdEyEmAjjrEP9fqWtLOQkYbCW2+oPcFjfOSaLyqbTb2Uefw2o5DRT
jYdJpLU8FdO1QzJ+uyGd496SDaKQ6y8u21jqsZ+i3PdrnJSgsIsNbVLF8LEiTNbG
sIG7mxPnJaCEIhDBf0HtPGjgKjJaU1JxGvqOAy3h/lKXg53Dfy7+hhTtqCcPaF0q
DsrLnilo1Fg+7SMNm+Mmlop1Ea4WF3O9j6w3GB4HVe3qodMbStFZNFPXGkOk4EQm
Mff9cOSRXLDtF/Da/bBZGMdxXYKm8+/ZHJ56Id7Vp80z/S76lBpAOBUx76bAGdRe
GCOOPtHHDaArkClbjNmbEMZhYlDOKJfY/wcD9Vyi8f8aHXIlSaLnFtoD8WAvUuwZ
aZHhFvFKbGXE4n3CpqI1Pc0pPhYgAo3fhMP9S+FC/DIiHLm3Mt0ZcZgXTgTpcG4A
HwMTkuDWCjRFmHt29rY2uqhjxPHlfyCxrNAAvUA4Iwq2G4ErDiO82so9rlZSf6NG
0NnoR8tQQrQY7FlVKd8FIQBxrBIxn+L89fR5tOw9GG6FbF0F/l72WdJybBFzNapY
KzExdHv2XxzmY13VtzUO2wYWIXPr3yc4bx+WmyD7I6/tZo7kQvprfrUeTI34ZUjB
JgQo8KkbVqa/mtqWPgaUb4ip4ZC8P8fnHcI4aNDm50hct66d6fn15nVkN6V6HGn3
zBGf64Wn+6ai3bHAkqmpg+P1vsuMaU4f4Bh5pmL88d/KOVR/bqlAIOhGL5dr2DYr
6dm/dIil2PWHlTJGidbPnWCyn1MYKIUWm7Fvh0jIDn/lYUjIciMV7CHGbhrds8zJ
n44mx2nU1XjWc4kN+lrOTUmNfGnP/YULFI5eP5ogcxGJn8a+K1kzTLy7m9r+qS51
X/vKyiKcNsMeLXlENxh5WIpfu+N/0wl2btPPoEkOGTA1/6oKRjc7w1jJr8ptnt7p
lTwWm7jpFvVB1Eu54dzHqhrvXSefF9T1fVolPXfmDqfkmqKFcY2CxLUeW6crof6Z
Eti2FiAFPaWvxgxnbQewI1KXvXTP0xgD4STToSCp8oEDXgdh8hnEnGAG6319E0pO
RLljB47itX3Y9PQtOWVgsnglya0GZI43BbF0+qHl6vK2JczIyBMZrSOEMBrDNqV5
9YG+PqMtOiMv5z7kMonqW7h3nxrVFqo9jt8Fl+dYm1+fPDonDecnYreBy4asMWDk
V+/17Na/NOvDO/3Wn08H5bPPXGgQHrQ1xFUB02+fBCtHsIKqHNhj1qeMiMZira1R
4+Ep0wPa6GWzDLygn0P63lKuwC5HUSLQGCXNjkWVeaprTcIzJ5S26LTUmJ9spkQE
LJLEBgpj7UnrjANE4QvrJlirj65lokDSnPv8wKqmwWidQ7xQp+RZ/uy9JF9hCdiQ
1zcU51zhlR5x4UgUx+WmwDzRvITTReKt8eyx/Y68tlV2xKXYmEUG2HC1QRA9g8k/
YOHBhuHHVP3ecOjmPhc42pG8GWImanSz2umSczi5kweYqocRHtxWeBdwLzf7yF1h
3+5Mc1GzvNNJhpqOEu332YT4V+fliqJIH8bdS4ATyN7sK0UG2BNNZL2aGr/3/pRu
bVzUWgWDJm8DT17QU3JqMuoRawGmRhhDX0qMEe+Q5kckJOgVX4/VMR3ZMnVuTnVL
c54vKl5COnWufwYAbzDsrqyb0us+y5Tui471YEIW7vkrR44S+N8w0RKfOIlwp2c/
z/m/VNhjEtaykidVdfRNs3sxp1COKCgquvDXg3LDwUYv0+8kdVm7XiI+AgK+0Vk4
4a1y2F7Z8xw3Oohhg7sE+lNW9p3/jBAoRWM5U0b7Wa6JT494oGD7uPngLLbTorH6
hWMAi3R90rvowmeAOkY6AtZcBhh3n8xbHdEfTRPfdKsQvCjZMWtiFiCDvVqcKfV3
wQJDojMj8FWGXne4FdC7M2YXupGeE8pGbTYC3UaIE+f/GCyaPMf//NFe8RXh5/Q5
mDm6HH6OBWsH0Jo0qDvxPhKc8MkdOonvyA5TB0YCuKhs9QXCSD7rPmvTawhrbs2U
PhUR4m/uKxnkZRBJvBa1U5QFF477TMCBKOZMqnYy7FeEjYcEpgE27hrTIWlrwV7l
QVbsTNP4uP2RHzjnJ9k4ikxdhOcQUH2I7WvX25awT4Mqir2zt129gs4NU5z/k/iV
7JDxf0t+KuVhp+dmCgMwv14sQ52UIQtPhBiychTWhj9NsIcmeneJ6FYvX5vk3t6V
jnxK4Y85/u4/9LuqTE0qJBvPk4JW2cEKe3e940O3BfoggNB50oGuzwMICgnBBJQ1
z5l+Qrt+4iNzOf+xkLU9rkCRUqnsXr04zUjozdHASAP2Jfunt518XsCNZlaItxtE
2ojVYmvlb7g932LDY5rbPsCPv8IJDPcf73z+HFHF3zqxkzsCZWglPHA3F/Ic9Cqj
qXPtN7vlY6HxfsvmDcgHn0T9VyllkUwimNY0MWLyZ37lPE6qlVkJhyTs8ZHOa1Ck
5XqLuXfV69EmSxJ5k+VZ7m+dtm6Z6bWbTj9xSSElZqU911ychQNujKAcAQ5GRTYN
YzwtggQEsMHgcwTYn/405ezUQHrqguTcnDcMzoB02Svj8fzLeBneKnP68+sdfwHl
ZIUbGHJ+xlpYn6SL+35bWd1uJlWBIG+Q84Aoirv6gVRqXJJeoEq7GmUqkdvu7AI1
8SVci1qdSX0cmihIvr62dYAjKbsLf17lQfOqwOIRwhJzV3iXQ+KYDNCwJWr/labt
HGfDp8st48+MXtxd35kGUWHIdhjHnJ5fDJqHCBS9NKPgaya3+7l+lbNEiAP31pIn
DY2DKAd6LivLHJGTOl+plWeQ2XdVDOXb+W1rDU5QaMjGbR/hIRhipPz378QQ0VvR
CwmcDlDYtktBikbAUIT5KNl45p/sEIr5n53u9O9iee3kW/oT9JRM32mXjJ2YaArX
NQWpav0kWNXSlNBKLio5TEt+Fv5ziupTBTrum/l3/6VJFGp6kXTEfpjspuou4AGF
2tdwHs2d8T9AzBQcYH7/5TFRYXMcgNIJUMveCXZcm4Y0uv8AUY/iadXhhvLbnYOM
/iirq/A6NtoLU8pVoGHgt62RnACWZb9yzKcq/pTNZ1jsDfdRJcnSfnxHadtrbKEb
BvJ0JWS0ckIJ5eRu2VJFKxadSAIrVzIVdGBPdTStm25ZF+EBhjVhXiPAxf+vWhwf
5nCQIQOnPDPohK9M6Bu9G4WDJz8pHLha1qgQyIQocObnrgPhdEY+c6S7L53x7/Y7
o8UjBMgIKfL/ELe7ByxPUya0BwUqde1qx98TP6KlJEoulvbx0r8eTziB2jR1RG6X
dFHDG9nPxe7TPxnrUGX7d5cwUyNtaNipEi9fkmaCRQSiz1PzksMCRtaelAxwcr/3
/ZqWu5HHfie1CCfQCvt0AWrD5R5FLvzMQj5b7qvrYisZUiv2szOD7qWXivZOuIqg
eKV4PClfVny8G+KJQuAMAuGLgND3clsDZBV/QEVMm2HzedGBLw0Ij0q66e3YPc9o
yLElsSzEOTY44Stnm2op5rfVKou4L4O0vJSTYI8fnzzFGOKP4+d/k840H0z/MBUY
1DkOUfkX4TSJ255uxiRB7PaP7PvHBCejeHY9JcrBp4AVNHHAoMdroJVNjU4sjOLl
Wi2h2BfRe9GtZwobikEFjC1X34bv2ql6Gd25WSbUoz2tNfgzq56mGE0MvqSjnGJV
fF9wnnA3k+TlQC+8A/xj6tPsJnnV29xSc5pURnqpxeu/j7e8HjGmRyICzAqXla9K
Y86ywIsIXKYAA05KzY4ymFiXWsS+pGKLC3XErFtx6bJYQijTD+XA977Od+nmms5l
NX7WJLAjFHZms8+3R0hlZbybyglpyFRFWRDznKmg8l1cqr2Wjg23StkF5aTrDLkX
DdhqhWwT+8hmkDpjAxpTF14226EHjFxNlnzxYPCqkoPzcYXjFP3vG8bfEQAUj4pW
p3w6VBs3ZWtKH9wwVikZ5mDhLrTVZdWmL0cpETaCQjDuCRAmWAx+xek8Y80etMnP
SOa9Hvbg5RvV488tzuLZtNMUT9yJm4QKldYaycZNOsy0Y+HbU0bjb9V/b3/vFnu7
NfZ0Ji3Plclj+rQrI8Qi+gysqmo1SHxMtKU4Tphim02e7twP9tlaPVXIcDUlBJ/6
8Zi6Tx8PSmYlaboNPMQiVdbLl3wdkcrAmg5Bp31wbYLCrefE1pcMxAu5dfYwMLPv
zwAZnjUwJOehb7hcLhTGyHaLGPkk6ShnznQNA1IrsAbmU/fEZqPxGOXyQ7SNckoc
iaa8PmK4Hp0+nldbxjrATK68s6cNht1wgnx4yTrxokX7jtNSo6z/umXMWNbhcwcQ
9VA1AH8pHLRDYHm5wjdvg6lxnb79SAlBcezsITGun0nGjBhSH/qOttjIjI1GkStm
GmJVdsZog+j+KKKEn3xeXAFYu5wrfY6UjLjtPjZ2KALoAuBv0NSp2xNSuXGOTgRl
NiDaJPuPL3/TG79GVt6fwsQdfHSwsoT+9mFvzPmBmL7RzCc5nHeD6TpCn5LbUCdp
Efs5i8ujmicr8gycsAJeOXv+uJAk3X5pvv0az5cpCBmCmD8JGxpVha6/udK7Blu5
tfK+eQfy9g2wjKSv5jrKBtC7ODYpzUDH42kzQrk8xVfBIJRgecPb8KJ4xevcfoxN
AMrawo/3ykBVBqw0FnhwhuJ+vz2sQWm9SooEW5zBRlymVoJqAzAknupiF42vj11O
LNt9hrq4LklnwbayTC9eGw244DRS0/1z5yR6AZQgGQnVQUxQXtFU/jd69fKyz7p7
3qT2Xnl9TBjL/dXly1hocB1cpMEUTInbwTNemYk79BZfHE9gRMh/rc9r2fGXFw81
jCMvXVae5JMSasEcnkctClSzRKOmayyKj6BgVatlqfFNPHzjuHq0FB3BJ21ppDMK
SMFzPfCfeMXHgrGAC19F1k90/o6nvwACSEdbdr/uCmRw5iWQ5t6eDuYNh/DuBfM7
46h0sd9hWSY/ofzzDhya0n7bGqup9bFiOcEo4fwMZov4PQjBt1nQbLVGgYh8yoH4
htz+Q7NYis1AeNTRwVrP+MtdFsQGPF4UhXcFdYDOBQKWKEftYAnoaPYUQxT4m4v/
8z1SvNpIPHPqQNX4vUWPArJun/CSdiuRk4qYA8C5rCoroNptbuEc/8W1tHhju5dQ
ZTLo2BDQgU0MEKVdXe2gfU3anHJnP4lnZrkaQ7kSR2wXVcEFcOxnqE7m4Vi36yia
joL7x5vhQQq0COT9/+hlFAphYETnd4BcCuhqRy2CZeuVs9glo/hcW40RKdATF2Vo
20kyURguAyjeBxnz5cRCoHBM30SYzvQ3/RjG2v7EYjGE90IH0WAEuPE7fr56DLh1
ihCHq23gMbug6PCAMHh/LrlryLcMprEmZmiAb39DFgHihidtQKAAcjaqjAn1fuxz
Nq8XznJgyY0abrs6+2UmPMcYe7qKXn1hxxAL5+X+c2XPwznrjh6pEcyI0bGLhpe1
sX9GkMFqhMrpv92sBAoD0mSSRxxVyZw30Ami6MsZy4TPUhHa9y4jnLLVy+pPI86n
30abbxeSWYDwvbHkfhbkF/4v/y6Oq+2W31HrokmcbKkCml7F7lnFsY3DoVQUe5g7
exv1U8k6r2LktOqOPoahbPUcz0JpYUanYovCoHORHRYNFsX3NvL27+5D+XNOSzjV
bxJz5M7+fp434bW1wxv6haq4tCVCpf2ntFjHqqt8Bs2IoXyJVhIpZeb9M7jOwvKT
qQ/263R2dBxExX3Qh9yAvHaXgZtW4MmMm9acwZqHIhtD5Mov3Q9KN6T2t0vo18nL
XreS6pqiuS2wuP/o+g3KWNDmkvLotCWM/HrtOpb72m5aRBjYDKHl+UmoysoADmSx
qNgR6EhyYO9H+QZeKp7QwiAsRWHsvmsdqCNwZYm6V26STt0BDOvZkwhbtA+RL9Hh
UFTcA4erM7I4jbSNUGfH3IpRsf70X1A02hscxOfGvYrNuNltC0tiK6PODW689eKC
jSn5XdbTCeo7sDLSouKVqQgzdp5l1nsJI1nlwOFZwmJcuS2t4qXNwFmaVDy/17dV
eGXERFbUQf4qXA4hxeVdw6L9rTU3OAm3A/gnrFVlwMjzRQ5hTTsY2EatMBM5HSnt
kJGhLKQr7JzzNMvVmDLvjc+fftoRJivqaTVqC6Sn+rCqd19pu5tnctSmkpAfH+FB
eHpdFD1r6ZBdEYwhDbGM0KBqx9D2JvhZPGlh2SwlIZN4A0b0RSb6Pj7rUXnbOMhK
urfbIyPOaPOSsA+3sNQrEfYncdhOTh5/7rYlfinPF0mkqkd5/gpnqdFOu01c8JVx
i6jHfbVcpdjDrr2C1Cc1/u3T4W3M91ywu3e3+ZwMHls8BLxLKd9FHHWt6woZbsQm
U5S2BKSsveQ6QQTd0k991fcdvB7rPxPin5oD6BY0HGt2D9HafGYqWgI+/d2po9Wd
cuGZJiW3HFAPIsj8YAqKgRItnUu3W0Q1M4XXaxHUqE160IWk9XK7DF++fZQSmI50
BNEX91vpSQkI4wlzbB+EmHdgeD7sQjiPapU+FDAB7ZUHy34KMLoKEe+Ha1stLKpf
udMnAmDXHDgbdMs5oTPrMFholdmqYNwSk6telEpLoZkAG+M8qtRpKLySVZXaLJjP
q4nWWrIBT8OHfWh3MJAPfDSxTKUJjZpfIq4rE2gH8UAI6gad4uAbkt6WQucXd09p
9S0pvQWB9lqgo8S0/AgxxgGyGHd9hAAQ6V7FgHYltbtC4vdgDDQ2bGNGi1DL+Po6
CNLTwGuqRjBXMAFrK1XkxDycBiDPURDIsyPqul3EgOtwXJI2s95Sj4O6bHZemgF4
k05Y7M2XnqYl6V0a0KhgCNpUZW4DkybeIIfO6HC64/BH1flYVQw45oazNW4YtSA0
JI1hZNoJXObq100KLoSBhoqgxxPNBTV2i56TK8TKuuyP1f7Irn/OGkuH3IksLA4N
WLLBny5h2zK1qh5ObnnENyNZkB1HVTmovj+SXzXMW8FiJ7DZ971eHME6FKPBp+29
1PE4L/LLUkisPQj0dihyCzlQqu+4W/0VuuIm0AfehwA9zXqIJjD86HOhUr8QgX32
onRcbd1P5rLu5lZE/DvnfKcskjn9l+7FhCUy2eYI//gNUKdBQzUuyvxGG6iCJoaB
uu32H5+PPsXwsRMlwnthQ8RbwQSiEBP7DtUWHP+2PVTp7g4quacATD0/okac6cya
jtBQV/kDCg8DUPtsUKI35PnFUXEBSyXbuovU2StJwk7jSpWwpusndWCRpk8TJHWb
885Y81UAsdONflo/eyOMM6QI7mbo6i+AVKU9E7uut6EgPKXQBs7w8FAPXLJY311V
L7nszFQPgBBd8p3ng0czGhXndDyzk/Of1TltIhWowW+TRBk3/cxcwfK7Hobkothv
GOCPwMgkvEbIRyornnauTew4Gqcay7bm6D60yzuKfZGbYdjKj+KZ3JeOSbUUax3h
HIVzBE/rpOHa3yhifE/YLEe1qQ9T+Hh2SshxoZ+3SE7R1cYpR9MM34f6hoLGijFL
kua66Pzkyos/WeHFRwmpk2tttQnkbtW+O6n8HUKMvO3DbHc4rJ0BeVsybMcvuuWh
/5TmORCiRGAMFpBGazyhNKuR0hdGXz8ztJz7zRMom58XWiDYWMd+weMORpNK1XBy
84XJtT79fnx+5F7zZ5knJdhM+Z3d1BtyeLT68Hxy7VTZdFDDAI7hj5CKd79+yJGK
I5PH7SIscAl44n6qgBhAVMr3Copsq7UJ06rU03XZwJlWKjhv2eR8oF+t/2PNhpOt
gof9HnPAp8bADkqtT88W33wz8psN0nnXAfI11Wfyj2u8kJvZ+5+03b66vRs7JYU9
iaJFcwzOtxUM6q9ediX0UWnVcBJXp2yiezK7tHSCQ7NVKM5DuHa5sWoX/nY7mt+0
lIIZMy5rGTINog/2w0Kr0OgChmmeLlEVY5jCojYnVbAumx2mlQpBJ19gDbtgmDtK
nWjnkJr3HfjBFOm4wqLfQ8qZoFc+8UOraa5dpuwanJvMhGHidvhXKEa5HPo/TBm9
KW7EHxOMoEy5egkteUh3eZm/mSma+kgzj/g4hgLPHw6tfptjkDR6fJNVI14UVSSW
Ly/yMvd8MV9HSeO6ZCVeS2aS30UR5iD39BYCaLJe0S7ohGSLM/AOtH0xVchRHyi0
Q0W4TwonyMS9Mp/u1p5gejFrZSzz3eA5yinar9q1EzPbpsEecAzmWCCqnHpPtiG6
p87+PFT5DI8IWCD2+yo9GU5X3poFjVxw3MzDncBAC0FIc60qbjqyynoe7Nj82ANi
SdQtQ9qs8YJCjS/vqM4R7o1HvuL3LlZ7JegtZcPtQwnH815DQdgHwZ06u+s5wyQn
wCtD58dFFhw408Shef6CvytyeVqcQ0rlueIt6ztuWin+7zIokbq+klGdEf8D6aBK
T0XjU4loOQZWfrcRpFkNdz/Li+pFnzhiepL1JSSrhCubOBw9ZjWUhcQfCbip45xM
3UEvZgjc9zMnTW9j+HhoBgAuXEOyaeWCXXQfDLsT0x3VEdyHaWkQSMIT1y8y2XBh
/ShAUDs8h74dZw70xDSpC3xa0aCrEBgRS9BExcny8MP6+AlHB8QyQQB4/uh1NpG3
i3v+z3lA1aDHI1TOaM2dj9bn5cbacDra1uVFwllJ5kWMGpzbSW4LnWUOblifcvIL
BSssJLvtL/bQQQjKn5xSizoLYUbpixjB857YtZZKwFQLeAs1UxBfIhVt/ydOu2KG
ueIS3IidVFV/Oxh3+qlWFgnDx7HAZLED2BIBMg5V2J1DjY6wnWoPobDzIpgNOgYo
Xn+92Pc/d2ocIC8plJ8aZldlnD0SIzMx2SuijjZIKkTp6xewHX3WZuQxiRW+s62w
/MQ8YcypAOniQOebnyHsmRPl0eHAcQXn39yPN5ExZDy752sNe6RwMld3QuNUCN9s
tAILSxBWRMhzSV7HZQLf7nY57axDrngmHfiQ/lHXiWqTo2jqpBvxKPstmTgu3cJ+
dtN5Ympcjswyp9QKr8xXmJ4rz8py2g7CxbYww6OaoOrkKdZcMYypnMIYMqSpDGi1
fVhrOiGCoSC9roj05O/qGf9o5d7ED5dBexKvO5S3WG3jgj8GwApkbt4zRKtr6wTA
pfVC/7BAqbGcLU7kmLvhMfbFnwy4ZUweV7UtmhYwPE25UsLRdVARBWHl7P1UgayA
WOjCkO6ctrSBbWRWKRkSoBVWcZRPEW98+zLH5qNfI19mHY5vMNVgwvN10bfKXcQI
KJLTkJHlchv+1WTuQ4KA8Raa1WxO8R/ytqwZbBjOm/icIDsk2506IAAwM4cxyg4l
vgWYIJndSbY5HkHWbxPqq527ir785GOVBCy98BdThKMy9yrCJId9I74v1GMUSyaI
dzUljolXc/pB7KgFSgGSiQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hpxZTQSnuQd6LHBLL7QRdT8vgy7Gr58E15Um70qCUBFpTdOJhEKZ73p3ZFvwaxK1
L+O6BRHT3/qT0C4J7WZ4AtqM+2c5sjq4MORE/zdR0ryLu4mJnIWZk10BM2jtGKG+
5CyVdxul3p5PZQkjyVRx4K6J9SrqbCoQrvmq6Ia2oT+ERJI3IsV15SZog4xzxMeW
ZKTugeBuPj8LS40zwrOy9c/ui0L/symcs8IYrtKk42Lp/BlQYkH5ibwx5c33aTIX
CPFv/ZXdcE8yhhaCDmCxOth36WSRN/bt4f3d1KHs2Zjoi/wwIkE85ncCe7lQL6Rm
SqlpsQ7OvJiatmkcK+y2HQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22144 )
`pragma protect data_block
ceAOzE5HFst9+f0K5hpha1hhuyOPgDZ9NgZlXCvXKz7jm0vT093EaG2lZjI9mCb8
VOeVEMMr6wmTA4/e6/4RJBr08bk/PPJ3TLfuCqFKWOmjQ3N6mRzCtvK7eaRLNSHs
OI23Bsc/vwctmfOWtGBh1nNbvHToRPZ7G9R4ZTsr+IBvIK97aRUpS8uHlS4wEfQL
3ce/o8f9FWNXfqDiLKtulL53BZye+ifkm2gcBeEwQQf9JEpq97sCnsZPPbuOmKGv
reZSXA8EsKItx/I2C/Mhm5kYmQGyF2pZxNt5V5cgvTz8PEbEfTvbUidDRI23vBCL
lax93sJV76LQZs8CSRGA9ea1op5r+eZCaMOBxHZpbpg4WygDIaTrhj0rPL7CNOU3
LikGnrjvdO1IEgBK1lRvyStDSdd0hf2y2wHTTtfC7R8cihWZHLlw3aGkZxpJ5Mah
ZMZe8qz/qUaz4iZt90hnp1sf1oO9WAjg5v4qJYe8sba0jEyP/cnuYhm2QRAlNnXc
ywNwVHQ6Dop4RU+T8RWdYUYtPfK2wWCGDGc7wN9fMRdQu+6lYq5u1mkafnObfcqb
4/xvyg7pzQ0QV1zAAllAWF0QuzLWEq5D20dlvWHpgG0wNgLuNWiuVLFYGFdr6Rdu
WMTHw6aMAStFLC35jJKLuO473mpKzxRVsvy7nwLRnTlvUGxMe8+TWmxivcXLIZAY
kWBujix0Yyz4awek0sFNUh32i+MX3uXhsSsBd/NA3LK6mOzyS7j2SQFyJW7rEE9J
SiUw534YgrzrGRrcwAZEZrefi2COfuD4yiIOM3BNxCp8uwbt3/wOx1L8g4YvBRt3
0QTuyKoeJyNnNoZNQBXpw6BQ4conY7JhGeP9tEM5DgmQ9czKEv0LEcEOv5ipH8i9
aSrRFzICTIiY4D88+lvzoi7neANz/JSNBQZf8zfI3inZT5EkqoNH/XcBO6nSv2sB
96LgePuy85i5DgJUtRauj4aR9pvYqooy5amcqzfTj4oWLOtt1KadO+Wxc/1TmyMx
Rm2Mh1k5ZfHiqKSVPG1X4jKifNNTsksxIGGFqiHw8M0ND4jnWpNU2aBHnhuaWNgx
ASQ3xzytGOpisoX7FU4aZ0pXbhQOK3OPxBfVWG3Od2QsE1kalsENyD9HqFBbfeEq
8bns++1WK9v3fJTzHE2wgAgFGmNAxwhhviYZFT8++a/smICLe3ouF5sBzZcvJNdW
GGBURUYCI0TYn87/9duIYhatbU2vx99xdb5//ijbpDxcdeoe45FK0m2e4m2jbP17
T8UMZTBlXhIYa/ULyDre229oTrsZfRu2HN6SPZN45EvwFd/oUttQ/DgDbycmVwdC
LAF1BQAQCsqL3jAek8lhpnhlrVVagYkjkxikVeG6A2u9Br3JaZQ5w84aqGAvVkFv
IJ4dzeDdat6j/HI6NNqZ2BAOiz0cJ52FE9xGVKru2qlSAlJIJpLJgoRQmQ28xZrH
kqhDUa8YNWs5lHfx5HXS6X3LInzDH96FrJdNRIA6pD7j7V8MQLFuIot+S9fGg4aO
A9dj85VmqwtsW7VW22SBkIC4fmv+5rtNwrzWQ9z376aU1gprKZxyzz4I7tRfjI8U
/RMUwKlfl5OFqcBLdLPb5DXfsBeytRmPXJHRVhs38EK/myeJPrudsQ6WCjZ7X54Q
UzZD4Hhpoqm1isMQ0e+lvIysizx87v4t4YpLxvaQyvSWPgAcuRTPvgByT9lDJDsB
9W6RsBn6y/1ViSb7iHHlwwnh7/FZJLt/BdaIgV+sezHW3fcSs6plYEJbNng+APlq
mqHIJILBuiqWsfCDlT/QsACZINXIimMqesPgGig4A0qvlc0n8Xx1z9/INL+To0Fx
6FYDpvOxn4BA2Fxy71ZfwnExzHJqOrgWIipa88hCGBxvRsJS2JdQDr5TlHLMwj9b
JtJoBeztM4xGOPVuqYLMf8L94i3Wzk6ZRv+aFsQgYKeh9Dh6jnWNpJAr7t6nSjRX
Vk0xo+ytNR2bOq+mWK6IITDlJFcf5JtkFFjTWCbQUDH+EUuY2RIHzfs/Kmpk2n1D
kVomgFHkRRX8sHSuRXTkGwcojiGxwvi0Mff8znk9Bt8YSQSRVzeVKPPG7sM6CNsK
NXScggcSlefYxwxm4lG6pbE0xmd0iGNdl7SdqtwI6sgH2+lz9+JIMcVo38fcXJpG
U2FJz+PGMHD1FN2QDFQbNYGdsrOL0zuaJpbSQE9wZXn3FNi36qD6NM4y2cuvYXFl
z2bWiAOV6rwDzA2ncPtSb0GMytNlq7lMlWVqBNikiqWobi9Zz+MJs2TC8vg08+x0
HyWY9sphCETjOxOLGeVRFgqAHYQUO7hErPYRd8bdXVUNqr8UfbpS/IDazzcYmw3I
JhVsUQ7dQ7uH/ycE9yTW519xL6q0W0vS7YobCXYRcI46BcxOxRAMEVHV/ehU9ixZ
ewAAY2Nwwd3DAsjB/aCGoldw2FZjdqk/g7Oo0NoIZw53mNQG2pI9aH10w1dMnAV8
E5OlswS6Mk7ZXbtQwAT+0QR88aXMPLxtEJhYvbjgN8Ntm1yOJcR1mC3Kw8N6cDgQ
IsOyD1Lta5B2VncoBrDM5nhx5E3xRmRufKUbWZgnwQ5GsXZG3SEQJKEfwTe1ebvB
/38iHmIrb1nWAIG3JmWatPsCdEzVyJt1d6H98YG78RJO3WEkjCCtoduz/BC3H9Sb
BNzDEe7FMtHH1IkxY8LPEkrZmaOfHLNzshHdL6O3HaV1uR2Q2MtNpFZXAIZ+Xkvr
+EwY4r/HUD1LrrO1G+kshrmGfI2OhjYwEIlAR7ktthDQgDsZk5B8ouwUgUeqGMLC
VuLQ/WlXQqtY/weAwQXxriSBG6v4nrpiRsvlEUp5zYUazRqRYtFjzRGa3oEyrn7X
GOACnxwjxvgTKeA0h9cUP2Gay7CyTtp+D5JcxphSayyF+VuLpC2e3Cb3ZD+LY7hS
IelHUmrnmEbkGFayH7mtZBVokxIme8t6MJbID1EiySMQNhWQggcCXHWyswfBaCBX
mKFc5kcGsxfpIxOAsPL0NcTqhFauMYpuk2MiyxzQax0civcKy//m1f1qHOWFkmB6
3atFDUYWttvxsgMYDWZ0xGiyBvxXu0Ykz4O6IWDI3imem0Wr1bPTEI9uTm/QKgrm
2X068M0H/6ULsbl52yarEuCSdW5ul1yXfqiR9N4fNyYfhxmORACswghg0p5X3t71
m3RhDKtrg862AG1aP675I4Ue6NyTJnRzStdH6SaRn8mAuYNTomI2F4NEMMdNAPMq
Gq8/Uc92C8uPt5IyvKO4f5jBYGRupi86Zqrx/rY/mwMcS4w2POPoO/Ukp5N1HNpS
AsRfAAtKuXxIJFxy8GhjvgA8y7EpZk1r97EaTqfwbhw0ZoZnsJE5x73N5hTvweVL
qdtIG1Udh7D8HJdWhj+Cb+uXRiLIupOTMwGmjCYYmYWV8OjtqE88u+mtHWL/Hw8U
PaiPKUNkoWUVeFoZtkyZKlKgrfO1ecPTwMTvRReUviIjbREysYcoPUD4AHMK/q5R
+9Aj2XrhJosyPJbZmyw+l6eamNbWPu3YcoU9Tx+nSd9KDxWnz6Vg5idiCXG1KAmR
Jxr5PnPSo8mOAgmhQ9wJkC4r/XSxIOpFY/Ts+WrSSsWrYkqtd5qq6mMR1qEpvRFg
nUJBTOj0mP9nf1MoNgEHTuPD89fEfHLSaKrSzZU7SSTu4PDgkDkBUO9pdtcL16RC
Ix7BkbzxhomGVoj65euaAH47A0fcaPn0c4wV7tWHVUN9AQv2OFOWL8sX9yvlPZ/t
krxkIxKN3UKA8j9+FrQgmBOJ6xx3iwxeblmQjn5BhxxKyOc+guYgi9VLHqzpNvy5
vujdaGCiyGHrtCKAqwdAhIcMdkiV9oA1EtnkBqrF0StilIMpcvI6DYJsct6BXOFz
/oaMw4oUnoGeMELcpizm/BfZrLAYi+SiUGUH/ySLdJbO7817AIuA3FRR68CdZPyX
hhWS9bDLgC72taEzSY0K+4gMKVbZxKC7rK5y5T/46AoeyUjKLmIkrAk4XWpj0n88
hMaGWtR+rlNCTcm+TBTPfPfTi8NwaeVETakEaS6BeZd9C6FcAY/Qls4oQmBPAvPP
8MuTI+VxLWyYoviw53Q6osHrXzVdygSKEz9u8cu3m7xNwb8f1wMOHvVPvhb9R9XK
UpHkBD/iYaI5iZy83lOILJGF3VqB8gFfnWZDr4tSEfl91d1JMGGdL/L1aJFl5zuH
kWYHKY4m3pOCud8ng/a3knfhlOqoC0ps2h5vRLdX5+gUAVxisj8VTb+6TtPpKSnX
uaT9lQSGpX9m4VzlN9jk3t6RgZKSg005i+l9g4XxErHTjYBuAxm4uIlkqjcT22sE
5mo4eQsROtM7SDGzstKi8sFEduLg8+sq4cybQxYSdB1EczDdmbxI62WPe+TkgKoF
9v2uYw3qJ3LusrUT0e0k5M++chkyuu2u6xNF4HQGFUEpmPJR0AjssV2cPLF4KmAA
Ywcef4L6lE3+uoF5LIH345AnsC4scEJpNQHd0IQjgCo2T4G801DaTMe/VD7CGJSV
vfeSYrN514iqkEGqqpyKgNDQ08ptFekYbQy54lfWkKTuDAbOxaUZ/tDbkJ/qC2RB
QoYqRdSOWN4gU4gSNI387fNnKsGEOpz1EjNS6b2xWx+83V2uwQ7WxNRhyvd+fP+p
FiWgIeTMEYDskjJIBsrFwz2UOYNLBOSufycZ3/1bo8Lnq4oXCU03g/kiEifAjcd4
wVVVi6gi5ztlk8mwUKhlgGjaH96IyQ2c22TFmMnQzAD+1jXnzW/7l6qAH/1IRHzw
8sr3y9ckMzX/hLsZTLhzDifeQSH94tR/AkLpJYa/qFsH15+bB5fUUjQpxWWcBn3A
xzj2hBfsYKYWOmrkj8K5vuYWt6GGnuo1c0mIL2IVJrhFhIsvSfu1Ly+gM8hHqgLb
pkmN4PZXESb7mozbZUsu80jrKrRHinEE5hbmvMmghdMOozORSy8NLwLp3013CnjD
fIUAUC/yzrrEYXrjfOVKFX4Y+7IBzf+Iu+182AdXNT5ZYCyQcoexaiKHd/ELUCyp
YFEaikq+2dbyhPG06l7LAXRSZXbg9vWxRVm1WHQYPxRA1b6XnLjdcOarhIHrgxtr
FY4ngiDMlqpF87zTbEiNmxcjw0R7gpncCSOi0ZXMewSVDyOHesXz+SBVUnOxH8WC
qWAfS/C+CutpjbjDvGcViRYAOBhfVjAZj/rGSacQdy/Dj5S5kvXhLC3pDxGMqJjc
TEBIrQjdx/1h1DAQI6U3e1vFoz18lckhtvSxc2819ywYhGEFZuCv6F7iKG2365L6
xgX3g68ODI33OYOGeyetrskd8lGR4SFHSzxfQiR6hC/3jjpDBdQnvnqrJZLZQ2vt
gUuCXgF0/wBMe53IkMkmKMRPuLBuLn5+RDslHNkC/nEj7g1jYttx1rkZh3WU8S7G
9EQFqv5109L6SZcmG3ZfcuzKrejhQLFw4nDW4RfvuX5YwjeQ32T5uOkeu2SBA8Ii
GSxYQshb52vRbDFZL8c2GF7zs5mgqdYEeIbjA6IZ24lfzuLs28F6ciCEDKevA7n8
RTwjzVfZl2axGzuJEGvFwBnp5U5tujdv/DjO3fzfcoL6Iqm/z2LlvX5zRnAwmvy6
iBpqpPu34FmEfJRfAa7PAqcMHvOOfAMBQ7L2PAvVGnSB0NP7k8rVXrtlR3tmyrHr
QZ4V9GI4qE07HJM+BG5f/qJkR6geleh6ECRAMeoXgJx7paip0UKX/n51XBSm/Ljv
eNhUPn9MHeRLAKFUZBFQsEaz08rTx1HvMJzR1FNHxFLfb8fTd7CxcclCsQDljfFn
G2uTDuYAQt/VuMpRgeKoSwCH0SjPMmyYk64kAjMXzTLh+4NjaDIFryOhwICiek20
59nLJ7gPn6o9dS90llabYlNJzvFXV23uM1dfG9fAWrAuD7HiT37B4vRRy3NPOhcd
3crP1u55hl8BsvXnx1C4PgMWJ+1lXSZZyFHs+i+Up2uoDoT9AKUmSNkXqMh9idPC
4RgAE+05xoOH891s22yNmk9QQqJ9HRFnzGyT+urXJt+wt63Ss+8K8w05hSsg65VF
IWtReoesBYjaCxA/1cVPJSlfwdAmKL4mf8FihmpKV1HnGF+2I6X1PqWUe/VW8KxU
m1FS+6y7uJ5qPfgAC55lmRdNfQKns4k7s2m5+b0G30E0ZAJs+XzOe24IT0gASKyU
HIZ3ebCFJgOz75trkvUXof+aFq/u9FPHamUJ9DOWyK/IQ1H2Fw/gLB+thKgviE7K
B998YfXpuBWOWZvm4svfciSH9c2lu04hUebf9Pi+2U2LO2iWYg++1npEurK2fxDk
slIhfqR+Qom7HX+DXitQMKA5S8qItIa+ljnZ6Iyq+9zz9b1RgquFinFzKCf3e6rR
TlHXJ1sXXLpoKmCePtvv4auhGyaqlRr/NLSFN6E9sObkXVkQmbBYcLZVnM70rV0c
xkGSvOd/OkYVQZaxdIOyGog237sq94Blk7m4uzDxqutdTxxzhfqn+E3qWkY2Zjts
XwbxukXC4jP9gyI0Zm/wjR+Wf3wE7azQecjxE6TNGgcnjZfa5d6m6MD+v9YwtdvB
2kBZ4ZN4lUF7okLq27/Xb/BZ5Sgj/lHhEWxIR4OfXIrvQWFM9b23t7h334SwOfLp
Zrl0dt4HSSXTFmI5Mkw9HLzA1jtxWwCeLA6M4k7YvvfGHQEyRKEtxl1w+UosFNdg
D7vhnPF3CYT6XcUzZXk0g0Aok8EJlDZie3iReUGnUL9KWrjgraWxZQQ4ma/ed5td
Ly5HiMx1Gzvr08UV6kTlm4GukE9b8Dk77WuqI8q5TIoNQmqs4hN6Dw8A9DTTNZ4n
LR7XZ5Ot/0QaKYDy5Y/5riAsE8rgPF/T9kZ6hJcq/R0g2QGrBYtqwoBtcu1EozAO
44j/6xyia/1YzBMlqRCO21+AYVZ2Q9DUBazYYKv+HvykO3DhNV6XSff/I1XPLM6i
bulDMfOGwTnWxAUpCFeOWS+7moRpMpG3nuF6r2yeDhMXzcr+Jo4ACwmEv88iYryC
di37tjsqQ3piP3GaFZ89GUwJwzl2LmGOZo6TZcJf3ym67CmaFcZsEqBmpCJVhWOm
RdegT28Vs3I59jX8v6N2O+sT9V/dt8k4UCVJ94P4cH82HDDr5O2WRIz7UZhU/DlM
6qETQJpvmkvR4jcBw9/3bOTAoNMI6eWgowSM0BR+ED6OMw1gmn97SHoqrQipwg3Q
ncAW0ERknGes4claNM3vmMBpOZE64+GymTW4sxUEMEApyD/HD8uUd9IlUwPsyZ+9
4s5or888GABfamKUPWNEuKSlX57r3r0ML8iutIv6EWXdZsKMk6BKh6EEtpUtT9Cg
LvLXiR0QnUL6fgVD589QChE9n1isrjpayVq7ridIOTON2egcOAbTA6wCZ31Fjtn0
YxoyvJFPv2mZ/L/20eLu/a7U4u8vx5A1Su5dlb1FdrcvV26TYZLfTGok1xXu7drn
qse/J7ti2toFlDH/jFDUlhRbRnADFgYI+xDoSVI/7fZyt04AuXuZ01cwTFhGvBkI
GupgMjqNpG81sbCAq34++q8EiwUP/G8OaGRBhIYbQ+UAscWK/WHOMJ1qS46idl08
Fs/Atnj4ydTqis3pDsd8uBkLK0LA9LCr3a3ZMOcl8wff613wFwotvMGBU+2YNNdv
fk4aLunRMAwZGZTun49VhgDLClhbWWnctp9ozuPqAzssJn8o86kngfRmmSgiArNQ
fSlM2NiZIvnpEuFs5sbmLIsEwHQDXjcf9WDG0732slFQgNf4cbngjq/CPouT7PXY
goWN65Zc/BmYVtCGgGgo/RoLTr0hJqFv4N80k/EgyR6wh8mN5WAs2UprBL4RYwA1
sVbrOPNB6yj8HAC/A6+h23Skr/MVzqW4/hAxf3sP8zJyqg4XzVlXzLPtbOstgjY1
oXbIR4ao8VZp149/l3iTR6Vr56tHFnKOXVpzQ+qtwcN9eHknEJM2Ndu1VsV2vph0
R+8rri81k4WZK42NdH7ZNMwP4HLGh7VavKc0FreBKwGH3Wr+xQtqPDafl289wLhF
du1Vdk2WRvuAagYuRrVE9KmstKYCLT9pO1Brh+/VGw6vbgo8HMlNvoJX9zsGcSCc
zJvJn5iZH04XHmHBz9zoj/xcequMO3d3aCqX8k6keCEjw6gXDneCX9z3PO0xAKxp
JHK4QKZ3AKtRs8KN1v2MSbLNS0z0lArPDuGckcxnSSKAG9dxpF3ubxlZdBsYBR7e
+Ql8bYU5D4QeCSc7P1jg4ZyRVdq3QDp1yPGXo4JWPBPgTWLS8WxTPRpSXUZWyZ3a
usCGg+DWbF5rdNrd0+zSqlwjBnZy4KmdbyGLraW3k3EM8kCQ4iwX/YwsI1awzfpj
wWBkGgX+zj2XtWBit7o6c0qMhon+XkGMt1AYBepJL6ra7IRBowruAzHqcy4a2AtB
pjJ1vVMYB/XqmIONFUSIVaZNSfoUb/rZ4zXtMQwPgG2kSAh0CsFZXAFCgCX81Yen
1Ag6QMNkjFIyAXFb8GgNDpVFTs4u5zny083Ysd0Bh6fJuayE0yLEy3ZR2GokOe0y
Jy1+FsgZrOVnKH07EBqqO4JLz11iDyzcOnm2hjvGCr5ICAHroCt2TdICiJATrjx5
PaEnZTSlfBNBiog7BcODmIi7MT8zc5l3M+shzLChPDDU1yMU3x3EH1fFXEedHswe
frOsqoBv+uFfH2C+NeSxe8ZJzE68DSwq3GPbdLBy8UpNPE9oGiOTqHkYHQVu4X4/
1sHXKZoYvK8SwpiI/s5veTRGz2LzY1X0SqV8yWpe5EBpPYBUoiMSkf3F0yHnz6p2
PcAF0PKziJJhf7SgQwBaGsWpKP7Rsvu1gSkPpib3D88fYBBGg+YKgFjAXENq+S75
WiXt6S2+AKlbC9Twg4cV8SC0rKBOm1hegPC/i3aqDLwgyCOKRyVydhaYgJyaoqgE
uPbtxLgKkhX2trTSo4RV5+A+YOIXD5PdmZl3/HgjtHNnDZruUIo4oLgZlFQrYhuI
pIwJCD+VNChOQ8RmXDr2KLuBLbU5WcliJM2DYMIlMDPDwAVxhuquKUMdscEYNzD9
VWCG3NThHkxei0jPbK+VsgoWfjYipjN5I8Fo7yh8M4pbmE26N8KVwoFFtlEBPSmu
pnLvDsgD1ygMLgykPyrZqZZHRPol+p2YwQ4N+ZZptdUhdVmdTOj9YlJQSfGI4ViO
Okojg1l5SyHpjWsPAuKwS78DwtiYZkdoJ9Yukk6YJJwKXN7vzscLljaKwIbJ5RO5
11g1DPRSeGl08gT0gGdn2axDum0MTLGZAXCDQTfHQOwK1EOj3blL/WMsOwLyq0VB
BCik8UFrkYxpD6654fMrHSohrsnZwawY+asZXk1Ck+cXqgG8xX2Wsw48eD6VqLQn
a3BctvJ9iy+5AAd1IbdrawMWLNYLAMoYQyyGx7bIlbGb3Q6mdYM1fMi0hFHcSNeR
vqYWMPzzc8bvR7CZGh4mrZXoj+zI7UwxPzTuf6XeApKGRlw+9eym1Rknn3Z6sB0A
5T4VO7goT3XWkpWacn3KUfwNZ1IjbBq0aEC3khNeyGzvFdEvNagZzelC1huWrRLz
Xl6FHjtnEXyME5zRjdsbnXc8Y4jRcm7GDY3bqrOELaGEwWomdxr0sY4OouYqDIBo
zYlfAJaqIriIpd+UVNj5xq82XTWiIIcAAgF1BmfDnpkafW6lrVOfMoSiGEo51pvc
kxUMoFDL9x8NN2e1uSN+n/IVtjQPicIueknS0Ca1eEGlpR3pnt+SRMC9xxoFY7gZ
r3ZrtuLp5Y8R8I5DPdWyigvTPG25E4p4NIpX8m1fcvQGHLCwim26Hp2fu2gVckRD
29xE5a6GbDoLedqLNkGHIbFzuxZyrIIGVMqQfKa9u2CW99jfWyO8oXcHqW1fNi6u
Y35lD7wU0D1RpNHWT7IMUeQ1kWBUbahoIwstJ8j9K8pjbHUda3ZMmXf2KTRvZYd5
lu+E91Qz9tsRowlfgxN33Izf1YQl0a14s4E3WgMDEs9QF4fPEH8qWDzWLZO2FJdZ
tN0Clxu+tF8jNk1ky4DF36MCqCXGm5WmvPraBqEYimQE/gFVyAieHMO6qoNtzdDC
WEJCFBDUVSKPsrLLzHUgL3HSpCfX8GFYvwA5XQlULdzEGJuJw3lT6K99WkuI8Uaq
E0cpFTfcWtxWJ4cgTDuvILqZgVOCgIGQcGCoqu7t0RSX9Ddu0tiiPO39pI5DTXw3
ld4X6wMwAIPYpIk9HWNw5k4LnZnf7ephyTXMr59M2P49OdeCbv/3W5/xUX3u5VQL
obmE/D80Is1CH3efpPGOKzz/aoNavhhyLubeXRZKdPmyP+nBxBzU1tCf+nfrrfcF
1i7voiwV3RXFtvL1xlNGUIrdmM/GBzkmRaHsEhayDFd7De0AMo27p3fQnABN6ch7
0s+rB7Zi62EILB6hjsk+r2rtKWnFvIjG+3YeKunNBtDP0jEvxKDL3IBf66si6S49
1j2VjoKSQqzRMQr/lUUFCtC/9GF/6SkdpmoIYEsn6IhFoPrnB0kZ8xiguaIWRFDf
giEdWkk3HaYDFGfAHwqHwG1u4TM0ju66xga6RDFwgKjkokp1JS/Eq1w4jHlPoh9e
2Z+Pf3dJl4VEiQYT9fSItCjL9KaAKccCT7I+LqDFa+xCsToYwpyCm/S6F7itk8Cv
VPhmAgXlAwdLWnHDzw8rGBH70WiF9VWgnXO0mTVwyqXArPZDYyaT0hdPil74RXCu
717aYlrxmlcnBkb2XZOsojopwSELFdfquizrcKr1IiGCpe2NDkN5JgD3zqs+k9yk
kLNH6hUD1Ucz0Rmy+Bys25pQ3oWcrambTZmR/jfskpMhOwkXxR9+/fW8BdmUJ3qC
7X7RmV7m9e3ETkIE6EeirL992Y5WrTYm89qj2plm14ltNSGX8p0GqNrve5okRde/
h2jfXBCgrVOH/1uH3JjVIQ+WQI66yEzEjflNGYNazxgzDESzgyNIhuVQtOGk0X4x
BC91hv/xWjq9HBdQAZytALnonKBmOeM5ftn53PqVo59LVKlsMyIphocniBxauWZA
iag3YDIxBgxG00YFb8WYB/G7G0Pt1++JeraRmiih4lFagPMr+u2DT4uyb+Z/GGx+
KQb/1GMWTQTQfLdsaatB756xkX5vsl821Vs6/Bs2WcHrC/ka/mZSg9rnmVuhP/Yo
CN0T8t8A5Smlsb1VfLSZDWfvXVvgRK+DDVVrDVSinuPCoyBbynSaMk8lhS8SaoS6
rPZtzprROPhq0iQGnk2tX9rOVoYRNsQLAtKNSQJuGIGQYLzhOv7bLnJfJkVaqn+E
z4atq8hFln+jYJckEc2PS6VU/Zcz+9X7U9gyr35UFPOXfzbix9Kn9UngyPQ8NbgH
3yPtgasx5L3WwFm/LN84VJbEfGHYTCT8ZKdYoFf07oQ4NYfbTJkzd8UZNQ2iCOuo
ET2IJlKgLXIFXfYaH1WjGB4bOjTRrA5W5LOBCSTVaoc5E29keXISvybsmGxf+IQ8
uMbwXLO7HK4PxRpi29AhV+Ki08FnEuZydpCOiiBMyBp93n/Hc+mV/HI6GYz9sxFh
PG0hovAi6JbFVYvCNjWes1lDO7j4xwuDkP7ZIVPO0b64lrtaC7oFkkZFQIyhuMKF
A90kYBxIiCfByx7BUKZFyUMStKxzkBF7FcePtTUNohh0hlBkvZNtaR0aNXbLrDx7
sLh2VHQTKYzyubw9h6UyUv6MrN9Edt8fYdKsckPehP6EF+021F/EfPZwTjpjFgkj
vGq5oqV7PgeeE8AgdT2de9QOwdarZ0uDrieEnfhEaL6OcH4NEVNVzwM+mHe7++8u
/obcULxX/rMImLzIdtAVwfOil2by6w8WiaHI4pVhy9AeQjRP3gEnpoHrrWsY0umt
dPmRXz22tOwFCXjFkAu0eaONUugaZe9mUeOoTByxVqyZT3fPuYF3joi2bt+FFLMh
peI7Q0fUaTBYsEh2NHzDAnGW38ry7z98caXt0E1Jg0SuwG6kS7t2US7Z+qQr6Vac
lNKESZxhp+Qo/h6RZCrUH/6VDQPAbXFSCOAQGKeXUJvTCW1HSg+at29s5YS1qbFu
kykHcDhgT1r5/9Rd98pSfyRjZDowOP1Tk5f3ljT+4Ghqdk3/34mau3/iPfTeeCBy
wC0brCaDw8Z+dT8+THCskyhjKD7KO6UKqS04RvMfYS1OMbEVAU77SkIPs+17JjIB
hlbs+Ci+2ifPL4KZpcCJmi4kuBMC/oEzsOY8y0+FEaqMipFvgu7zVgZ5g3XfDTfR
at3azbf2noPBuIF/UzWce/SeKFEH7Pst38qTQhi279NgdjrWTG5vMpwkI0UggAaa
8fx2NlWba0BSlBxLPnRcI9ACruy+Mw4J5E7f2F2cQfSQj+6j/U8G4S1C8IIqhr5h
HHMTU0W3ceQOx2qSz4iAsIJ0FkbQPw7Yd28QK14rsqEOt8t8wbj8w30FWeOVl5Lr
OrjS/d81w9oHqem2fVnEd4n8oKaoMaBRzcOpw3RswTKDqWDkmVb/Bj/x5F3cKBmH
0LUmP4psnLC+THL3IFisgePQHpqy9duiBFJonLvl3maqwXYrLd/xrRWn8rJTPPdw
AD6VZ9c+qVVH8u2bLT60dDWJYdmB9faaWmhd74kOOTzsn83fwsTC4lEY1IMURy73
L49Rt/6wbF3DCa8AMGXZwA6r6/+u2dgzbJWF7Uv9SMjDkrQG6IGYBxUROmb+jeWE
lxtxGZhb4KCixRN9XfZZ/wciIK3qI/nzvZZxKsByq+qkSUtdBfy0hqx3mLCpK3Ya
lSoByLnJCz1sAuEmO/xkKGWxvVobFfWZNhakFFY7TnKKC8gjGvfVRq/qDYU2FiJh
Egv7q4X7fPMLdyDGAWzqosb3s5XknFNrO7mwA9HyUA+0js875nN+1Cpwbj3XzLdz
qm30hD4qB9xHjO9m9NUdtPTDA71LHSxaVGlj+8i/NBvDPjGmhrkuDRkBB5nPDVx9
tqUIv3augXSE6hs0S5s4N65p+5IP8uD1CrLUPvoQ0zmSWypXBtjFiODqHhrj5yip
6SBpiVYbipOglsl0GuMoK0Pki3S+AV3bJFBVtVyH3BV2qFMCf2zpci10lE80Tdjn
B/ymhsFdf0Fi1NJxy5PEnRd0XF7dYHkuTboiSF3l3scKAiKQ8vgaPir5ndHKlXmU
pbVIia9YApDfHcReX8UX7/pJF0WjJgusGS5UfAihewcfoH4NetDqRZSKhGVV/UFs
aTuP8MS3ffR34ec4yanG1fmWZ7dxVlL5wmNvKZ9Yla6iF5HXHldf6HtYoukXqckV
TbZsBWPqDXgMwjtLxWZSuui7aXzLOQ6kQxyW0hMbuQZdp3SRH5GhfvOuykj7Ra8O
FW+dPXfEV/jeLrBlwg+9nb5rqgqKWQiXAWZnoXhn89eHYgy/PBZ3b5nnkdUy9sVI
Xif9qSGPoG5nAMmzaFA+NUXtcNL9ZQD96WEZbyvebhTJXBKTF5OGzOOfzSMDQSjF
sH9v8+rm530ayuv9S6ZArPH2kmrlVbNG5VAOWIg2RWLIpFPjKUCO0jHUVNkuEPNa
dyCLXtKJiQSK8QFPuCHT+Mj3aZepRysYrc9haEQcbpFUCVhnUnAcRjwFaPa3bF1M
Fljnb/8bx7Uk37oVzaZxSG5SSoM8O41VtFJR9TowHc0hfR5ymaC+kXjqZFwAnOHM
KAZfFmUoGA3LPv4cD79uZWx3NOOV12Eb4V59/mIjlbFEwFR7zq76ssxDNT9FRZMr
kq9y6tracMadqICxwUdITt+q7sNTBCyec0mEGsPN8pmDleO6HGNdshDKNPyoBGaj
bu4dgNSB9JwZV1BiEDd6zP6PP/TQr2aY2DQrKC2ddwCEPzn0zRO2j2zwNSnAZB8y
gsey4BzCuMDY5gbLYJLLJoxsQL72e7fDTKAh1g31VeZuiCpuH4O3U859EHKz8dcT
vuXpVckVv8clx/HaNi6skSJzG9vunnebuOYJcPX30km6ilPY5tpoxTrnctSePbU8
ehhLoBgbZ17xgfYXYQtf8f1AZpFqo8PsSqm7S/a/iBhcYcIGcgF+juMFbbZMvyF0
sx403VYGgUI9rDQA7P/2TwQM+zMPHGXP+rsd8r3nX7ybLSXmy8ldzXDlq/N4by5R
X0MRuOLzSM52qa8rIxmT0/e0VdJnVd9hhbiGKRm9n5Qe+ZmLieA+DMlY/JaQuRVl
O3oJyc09VtpsVxZh6hcS/wiO49na4QLYtl/JDPDr0wzqNOd9IIgnUZtPOZRW3QeD
HIr0JRCpzjFUFDcmv4W2xEG9b/Hle4u7yLeog1Yy23LXlY6tklEK4gXwmw3gfH2u
nt41IMjPbGYmnHCNH/QDvOqzE+q5EUR0oiPEUTaXYnojdIxHHyj73xbC8OLudqBN
cy3pYOGZecbF3Fagx8iG3Pl0ExcdiDISLv2aM9Ny6h9aT+kdsGUIL0ZUe7f6KI2G
A0oqp9qXI43YhoV7EA1ej+OqvklSWgJ6zApcvSaDYRzZ8HQ6WhXh3/mzjRYHwWe/
3fbj5vk4ARbE12KofVj7WSJNLTkjstFliJyCKsUk3R+WyqbnFDZIPMTIOKJTzdT7
gQTKW8oQXNbEd7ee035RypTz3RKYyX7da2bRHmgWawQCmrFw0g3+HvkSkePbi0ch
C46ZhwMZjX8E5DuqyAL18rNHLlGdvMCGtphIiKJrVGgG2lwdQUPN6GhzHXY2wLYZ
lrzI+QozwkCZz2+qQs60H/wVmbpj6DDa3JkpBACQwfS8RaB5gLNfxoWhZkgMRuxH
uQ9jxy0PFE8wwOYIH/4s0MhS5hn8rHMREWhNMUF5H/SW5GM4/a/8UrRaeOgaQX8i
nCcs6VqMb/Bl546vzpQwGIiZIfsaV6/PdIHHdlKIZXttpyeVT+LQBoJ9fEQ+bQXp
a81mDd18iae3w0eZxDGCItAng6WNrKUwll9nIvdTbMmswJoAi10nleBeYd19uA4H
/raRH/SClyTNQXW7ws4me3mi+BUNgdEOfX+b3I4IAuAKl+k/JzpWJFsp9hOM/0R1
wIN+vHd4tgmSE5AqIkq3/hqodc5RphlfpdMn1xujIggKhVkpREtgxVRuZxaLaVwm
5qQc3A5k6iizJoX7XfxZiYJ3yPuI1LhqXro9PeQ77pPNHKVkUkpuKXf+ZYmtfqW3
Qtmcme+mvZOcJ05j2sd2VAf1pa/x872mvBtxbIFZ8PNg28t8O2KSWurjcwA7aFxZ
BvHfpuyvLEvhSNAEjazKh2ZurpNa6fDWidUWdxv96eM+jEepJlLLs3ZZqh02D+wu
aG8TLz2dm08j2aBnpXFf54uZ68sgSqyLM9loudY9zu8Yx9Q/+O3O0/8/0Ehu/tzn
i7I14ObkXHsIVQ6GJiLYEvlZ9enNzl/HooLcP6SKqogCPWmXFFquPJ9SZ2trK5hQ
D6nPbFooTFYu8NuO7DklRaEMVmtZ+K5sgVJ/9mVD/QlMpzuU7yAAG8pnee49hFNM
1I4F+2Xe7ja0lI3AIiXOhxoTyPkPWM+pJYS4nEY4eHo0PBQ7kUgWiSLmXyMH98qd
Mb9EJo3zfej9WCiYAspqXlZ8LUgMc+8nhbyyU6h9+yG9Nyp9G3HjNCfaxRkkniF/
WkvSwUA6ni73F2rMONT65fEcyk7VeCuypS+J7v5qF7fXNAx7BayHOxIlRGWW6JIx
kzX7Wz47xYnrged8FSvHHsLP0YaLK3RRKAc4SyqBxNlN3rj8vjKbaZhPOzlZYyw1
nTF8WceagTr9I5dCU5zSaQpgAZPvuKOnHgt0dsP/AV4SIKwm6eASQ1K202hJNja9
I3MnXZeZ4IM5DnsrMzfXdknyyho02iVcqigyux8eXtHpFb2r4kiZ8hAFmP4auoqc
YOUnUkLhDaArtv66zGmdhodgLgzYuYmtGl15KKHRnpgAKBDoUAoomcAeZqbcpmJf
lO5E9/oHfRZvfC7ySvo6GWYUKx9XJdQjOIq5WmEUMWaq9sy8OpnLOjyEps5oP55T
HFFbehT5l+MHnlgD7+qI45Y9KHhQ2udIyrs8NeKPfuT4n23V3+jsJLkt8/FtmETq
Jqk5PPBXDJbGnMlpZPUhas+Xo55/1wbrpRsDI05bbIQW1qiFl+1EsHweplmSzykF
6lm65SbWzcWQjOC4Vl1gy00QD/4ahpa2QgCLQbE9ZJIVVEipfrvD5o3xVwSVw0ev
6/a7f568AG5Fuoxx9RHUYMYW+q8DmgDQURb+K/oztQNjC487XoY1p3wv8veCYmlo
S5pGl6HrzhY/87PH99UPYWJYFioOCCT292yXgCWC32JLAnvjuL++ZM6dtSi53ZdK
Jwq77Zn/NLfpt6osxdPORjAP5duhg4NTw3k6bVrGBZ/Tf8q3QHzeeIdeZnJ756mL
iRBkSxGl5IN6cdibNyKv5HFmbLOQQ9FJiZj7IDvBANq2hl+aC0gxarwGzp8Woc9R
qe6Jr9uI7vpjWwK0vGCrbTH3DE5SGHtTR55EhGbEE/wFv1wQGS1Vuxvx9qjGugT7
04G7HwH2utCBG4ktrXS+DnvTeN/q6EmxWByOGPKWzmLJZCL/xuweHCCqwNRC3EKy
rXnCfzibW4QqRgubGR+Qbnr0eESgKxpIrjaeQ/SIz1Ge0f/VTqKKqaIBTF8mkchY
UZEvXMkKaQzHJ6xGUeziNR5yYa0dX7q+dw57aGsnciw2A8BnT0GucYDZPWNwB88a
1zjygWYnXRIwcqFFp8jTDQkBq5LOC5R0es0I3UIXN6h0YgoBH7+N0nk3aklyRMdK
3HuQ4vHCYyrywJnC1UV8YaUV7snuf0c/a6s1sF7RhrJ2+3oTv2RWMtgUrnXKtX7+
xaCUaGR3VWm7aP/5QHvhrvIPZyLe9InKwQDvrPukoIhLMjp3lKPQCRtw1/Z6BiDy
ua+QVKQNis6piEYILsoN0FeG7Is5imaPZ9ZrNu1/83ngpt6NChwLlCMnpVCfCRYv
Tv/I2/zXSqtCaOLEGJ739YZwd46h/4AeGwJnrFtIMJj6bXy/gGWpuyDHdUDLvekn
ftaML7q+1eWvJcoYxSXrl+/3CpAO8ub1NeuTev//7LKbS5uc+dd00wsWOFzBLKSq
aeaVcA118KdSKLf/aYBEZgMtLBfZCjBZ393ju6D+0ehvQF5iuM90jA/7qL4zjma8
qde8APh43DnufsFpaUGQ+ZOnbUM6LNCQTKZGtGn1FsmPDTFdeDIZwhR5aOK69XOD
hBMMcViA+qF0NHH6ad0rYQLXGT+JE+mZl8LfHJYvcmHjfS91pPJ6Jj/JNSVgmayM
1yDq3kDAl7ZHd6vrQwX8tX2BRIfkQOTqRg4/VV29RSYPQCAapNqQ8SIP3cbjYoaK
SJ7M89yvEmBioxZQ81m7jH8l7yYUP/b0h2qu9tAMIT9HLbWnDnqPkyXtJm7PRJ/k
C3FXozFMJ5hJNorfVJILNggTBc4ORWRK8SeCE5WPmeucPyMprFaWfVJvjpyRE06S
+QsgY0UE4tOLerTtOog0qfI8+VdLjGJ0oNBg7CYaHKw+H7CB1aCEg6RZr0kznjpm
X2ruOSbpq4+cghUz7/1yyQWHzbzPMbyteQrtKBHlXmbQD0lnZB8hDE5+eH7Px9BT
icyBOwGikoxEWbD77yd+3WeNLa7E3kyFSG4FlQP6C2TrH8K3jmY2ffcoNfaluP07
AgBJbaJDzDxqaXfsEsja6Hy5tGL7P6nJST7gCDyDzFskcfL+yilOx6nNSZKYGJhv
8i8wNQSMcYjBRFMga+ATSez1RB67M8tgPvaS7JrQuTB1lgbwC8cUuN21+8sM5Crp
grLiPfTSy6vnw3j3NTB93A8ZYQRA/bbr1jtGFcO3b5PGi3EXGWf/TjlmU/njyJjy
CWhmdtKwQwxZdzeFlKzvRM3n+FNK/ZtT5XrrWbQsKOVUdVtt8i3bxhIbpf8W2CmY
ikJJd5mTLsnS0IQ7LmqI9X2a0KWYgBVYXv9byyL9ectVrdWTVISHC8+tcE2U764Z
6fYXdT8wiRnI5Vlc7DBiiV2rwi+Cxrf5FUAsIQDvThTCXMwxbNMY6zYFDCrYDFNo
84uqVsA4ICK8cB6gNYFz/img+JldZA/6BxHgu4JDBRglnNGKdAUmzFWwwdDI0Hg9
+aqZe4Rm89MV4OlatKu3faswSVX4uijVuovMm8orwsF0u0g7nxdmYUrzYtyymjcE
n7DXD54vQmbDLt+424rMD0NNPh/qDmva5a/86nJs9ocku0qWjJCwtakzJu0w02PS
2WexVKAvMAUsdDdSMZPayCAoAeogC8Uk8TrvS5yiTm8tvENY08dd9ayhSLYSnjGg
StyMyVvaxj18M5YuihDgJEmqjrbIFudAdBg8UQZgU70ZT/Ti8TFnWQHf3ToXGNXx
QjrOsI2kytd/zYGevnEYjyk+1LfA/FuJhYBdwFVgsvH2Fcu/WXP5V75wg23NrUcR
Jiw5QxLgZK2E4h2Ve3cR4WleYZm31A/xsaV52tM/X64c7HMn8mC3gRP01+dNEvMJ
V2OTl4kyTiB0QnJcifQlfhFzKR4BZiaTvIqRkP7UNR+Wv895fJ5Ilb8dnfGzYN/s
hjgZEc+/UQNiRQOXxtBAbw8SlqEOWCY6MlcAKD1hJfXj73JG5Rc/tekotwoagJPA
aDXs4L+PVyB4hDfO3wnf2AT90b23Zn6qncT5xB/darbHtZ0gXu5oPeD7BRaNEIbv
FIsGJLU4Lbs4XZoj84ZTTlyECjp9vL0D11AbzdQL9/o4gcSE2SfTaRDuWrHFvWMo
Mhh1Zls56eMq0vsOoOOpILXMhR54oPPsKzyIw61FRNXXtgH3mgjfVWWHV3VGFxyf
Bw95I2dYFO7khvXiz1dXC7JQvz+madOZHTrR1jIooEf9k39HbJKyP+I8kzjRAaNC
mR1o4eoFGBOuDm9r3Wf+wr0CR9hkIjb8T67amjurO/Y5kacPUYjvZH6+LWlqpUFs
P9J0HUKjytABitX8NQwVvBQP4CDLDj1AJop4dtaHoIdcxo/FCzOgjsn3nUi6PhVM
rXSAsBRy5El5zNRfMZ5gc3+yzUqiGhHSGVr7mtohBxx7+QJAKSvoBK98T5F0QjV0
QTzDS0jBjJrun26185gupDu9hvAp9KhCZJcSBOplei601bVxqyZqDFHul/lgSlte
Gv13OIUurCTRFkO9Kb+4V3G9MoIj8cPcf8H29KVGG74k/wirGTLUAu3NuueXwg65
1aSYLUYdymuf7ejfjRHv/7mtNy1cQoskNAXf9ZHNNg372fL1zshi3WpsGbCnxbFc
I6G8cINQwxmrVGRgbWtgZYyXHzVYSLOtqbw5zzHP48tlMcnyhdxHNVxlLalL7C5z
fJL18o58zle1XZEAx8UGSFsXCupjsCkyf4eISt5sbOVDPjzZY9y/JtppmFxVg0gq
i2/am51dF6cFi1Aqrn1uw749NkGoubn3c0Ji3H+SbSsD7edbFAlFhOGSYjjN1CKr
AJ5F0quwmtibpdZMFjcNCacCHZdGN7ZNdOXbgJc6r125HFyTKjJISBZRUHhh3nFb
/YKFRXh0RBQy7jU1n4vm3Fw5oobOoUXDBiQnrdwQfW1Yoy1/Cn5uYFV7R+/6bRas
u2Stb2YtLGwPdvEHUHrLfNZ4EC9OgjYskONsu0owM9L118EiUaNA+3xn1k1lo5jO
GFbZj+AqN0gIBs+Yaoy4uR/sqzn6S9nyUo5mdRP0qZRi8TfPwGjtpGYJ2E7e4+2C
exxdnIRst2Mcw5iOtPiwF2U4RkswDUqHMfbGm8cPpoa4qis01t8Y2Ztop+3dAqOB
qORHxE1VuJq73g1FUgDYVYuIk7TxwgXxnQZ5i+ZtUkMY2+ik3xfyD9omu8QaG8ZV
P+tGSeI5xIsQ5BYBQg7dQDKxpPg+T0w0kILlU5gqC2clyOVb0DzYZUUsC/lz7Yka
zt3wtOsWOxrn4RiGpFSzDsZPmC1vkhS1pPWPg2N5yfxpYMiGpEGULxRaedjIqUFD
A6qH8AdXvz5hPN45J1LnroCX0KXzEAeFfhvhwgJ2nGuYeANDM0tml/4yURG24LzJ
RluywNuDgA87CtkaBB4xlmU+i2yoVDHjROO1hhVWygUzIVN7gp/OxYHhhXgugwgm
DwJFXfe879C7zngmF7q4hASJMY5Kr8edT0KiWi/QffRYDf2kYhjvvTCaf6fba2CN
40Le2iIx6pfanK1XADBDKWubUDiLZiLkbIPB45C8NhXVpRjeEM7C5mrouwmGQip+
uSUmP3DofiHAfmcjcbMJeHgPnsUlsRtGDzXFKzCFBeV9Kla6HQYIugq3+q8RF79r
iQyCeHwP/XXqgdd3CT13+EbgYQXDLiVhoynSjxkXiYps6PFeh0tdqKWClysHfbU0
6/vXhMspynwgDEQpSBcFSyMKt0J8rIiYyP93kqxJDFwL9L/wAcj9xYbuMHozmfhJ
LGh/SAIkfWVW+nmjmyKamKGcZE/ZmlRgO60fFCGu4fWRBelEq0b/cgAYLEzFN2ap
8jMccEKwAZXfdYIch6KNMZWqAVHQ1MrS0bM/UDNHePsKfTe7ADud6/kotvTfVPnw
Sy9Ork7PtZMj6oqjAynffKDS38pOqd3bhtMVbc/pgQpoJ5q4xqCOMuMPPvX2GMCF
JGmiDdhf7EjurcgZT0Wm3trEsM5Kw6qHJDq1JSvkNFqHGgIT3HCv/TEHT0EWXRyU
31NwQr0JzO4vPBHg0YpBz28Cpe9jrFPJ6Ijb8Avq6Ia7rtaIPwzOSmAndZ69HICL
M4JmUj6/a7YqlOqPV/MHZpFT4vpjOXXrgDl2ySl+77U3rq/p3+rElVGDqJYUGYmD
i7vdOABNs/A5wHeHQB2auuP3/47fBOnw0/jlIW1X4Eo5dNmqpJfg15sH01CauCKS
BfWit6Hn6Pi11Au278s9rzgyEh2teYgHDsnZYZVWO6qSr2r8lTrmIzSMVeC+oFao
ECkfsPZKF+OLHo1d8G64qwIeG1UJvhdcZ08mIIZN/npG6fOKQOFG+Q7MjV+svdgf
Aqd9M9Aj9HJT9sZw/06pb74au2l8Y9i9CkGT4tw510WvZCwsxzdImG7XYEnI+k5i
7xRmlTM85Xv7sOKkAvsKDD0jPa6OPNSCGyPYUJID03gRLCzesmBvyWjJCdOo4bcK
hWZjJ3sqKhi0oO8hYrc4U67+ezDA46aYPSK7cu8yXeZVr3xJtOP1JacuU64QIazk
jxR1TedBCr8KQeSmrWqJ6frq7/M2OSCVDwsuYUXfnw3UNRG5U0FI5Q9kw6amJ6Va
8VdmTO7eFvcdixnn3kJHoWhcAvAe0OJHpiuM3t3eljlxqnmCojj/0qQyUIxQ54tz
tcJFHiJbToV97cVwQSgCg5K7d2NTW5PQYfbqnm6nKfzhb18bt/y0zGfNXtJSXJEI
lc89AHPrur01XfSIccS6PV5Sn8IVSVt5JpHRtE73qOd13Ioly8KVlijqjWoCtpLA
C8N/WhA+kw726hTFB9+R95gvhNJUMk3CQ8rIjnJ1YpVWzL5gto0tTTANCXHEtBAn
BieC/QH2g3lmNp0RmV+q5DvDZzrnqge1e/rTgy8CzyBjZ2VO6pDRUFsQaZmjJNr5
UDuWEq/r7JxCSPAp7XEH8jozSThsRmb7NPHFOVvHMS2FFrKoMPxr5jTu4EDWj4tw
EA8ICf3N6a4Z5L6FWeCS5UEnTexFmvaER9oEA0xd/b5Uo9dXMCAKTWhf7+o/1iKh
Ek1NyKADpw3kKVfti0d5q2PgE6WuDidrhzfrf97N1W9yum+0esM2bBtOaBrtmd3i
sYTVQKYDs96NP65tLk0KgKkrHA1GoejTJA9zgAfk46p88Ylau/+9EoJuRq84CrDs
uJxoWJzPu2HQUxDAZqKu9wh0vqAdtWypBy9sl49P3uIa3ez3w5XkHI9XUeXT9TXl
qpzbeCYT2JSN9SVeoX55KJXXXMXhoeh15LH1Tj+ydoifE/AHlANTChEs+wJ+QBKq
5ImxKT0At8Vv3n0mvW7P1pPmHVoz4D/tV9EBpIHUtS33iNNiLKICyusJSEZI5cgQ
NpeaFMthZxf3XWu3MjhoGx3bZzD2Kw0C8vZvwIr+WxQ1pI8NsfFwXVj4g0EAMhGt
bMyV30xN2WNn4NntaWRE5Dy7uyxSjK5ecDdMuGbGRt1Z1B8vld1SdU6uL9Au7RHj
YFqWUogvElhpqurTSnkRtY3OLCCddoFoBaBaT1nizBvjyi4apZRti3OxYyT6vopf
Cu3tcSi7Vd5aQG6wSdN142Q2n1HrXsofDwdSRuFZQ8imGxy7uyuowm/iKyIhoXiK
yQWUgwuI5pcE97iL1/unX3EMxIzzttmn/ftz+alOPnHAa4d3fydKC8W0Ov8RoCI5
G09EdMU4RqWmbV42AbjmiH4xgj5yE3eTc18AqoRd5omMRek4maLhS7YElEdLpa/j
bYekzLjUXrcyAE7v5AZwb77FrMvp8QiE4rpFztJ1XOeHR9+kMBNz6ZSaUHEjQIzQ
SMGtwSuW7UqVl49mLf+Gu6IM3YgrRuA0uekznjoPk4u6JJDMtxt7Ty+6rVLbF2e3
g2MkJc2mpN4cZUMwDsR3/77P5pqJzDIc6+oTEUUCqe6EA9BgirhY4o4Q5UURxl2i
JYROFJkrMRp3w31/lm+pnCofItJCtTMKHdhA/jXVqr2S7hxKHF/lpdIdJSl+ERoM
GpM88NgUdGy/JV9680kAMXg7xW2jQVZKwhtfQtgcVlhFm4NQw6GrkooR4ZE1ITKM
HJ1k/0eisviS43S8Wqt8qpkSIKMApZP2EemeyW2in/xPE6a3iF3L7AEKJzxOwBpg
pdaTjR7ZRX0udCyjerbj37obSpaC7Kn759ymoLYsOufkhDPQiEQ9A7miLRN7uTja
dGe0p+jJJE1js5eSO//gn9xNU49krlmDm9lq8P2Tn+6C8ABo4d1BbANoyDpoif7A
fJkplfJ7WCxzvh73Lg0ghtB6V2ItAXtqFGbbOrBQELdHw6VFFk6/bHOpbF0izsO3
tLZGoHEyGO9GWqLlEyWrxT1w/BZy4xLf5DPY/ct1mOn98vYM40EAqGhiiajsG6US
cmWy2qKiuA6ige9EuCOeUfWIKc5GO4l6CInZlOUADXfKrhm2u/yQAb/B2VEt+U9Q
TdN1PXb5oL7t7fjpJvW/taszbjYcxxi0n+0XjdQfWqRtcr32D3glzYnxfa4M/rsH
rXMbtY/RlCcXXG/uMJhRnJ5YL3xQF3iJSjX9EEBVWsqVx4RUpjOiXWXjKbIE5BYS
MuLAJu04HD5dedHhI1fhNrVJbIS3M8bNZOwsYoxXFYL89i5qqTNlet2ErV4BytiH
T0/96OsZKvVWvY+754rXUNlBRLUzIFt4z1OZwf2BoCEoEJwQrft0M4pOZpwhgOR2
4KPw4OLqGP2AqFsTIGlzj73OQGiFioFP8Z+13tOr2OC6HpVO++7m3d90a/KceW9F
Jm+blx4ZBPdUM3rvIIvb0GNG9v5l8vVJKeO/yu6shwsaji5ymmiMIVVkydkLMTjZ
m2kn1cxW2LsFgR7/sESz4xLlirY/Fnfu8tVgPCfjxrkcL06qPwIzJhUlTF6PUVlz
JKSDmn+LHUwS1T4jRPj0IqFM7FqqZVxXfzDDPNaFqPhWA4CgltNQrvVR/SIwmgW4
CH6LBTovld1y7dybNZk357mT+G0D9bDAGEd3VDa18YacfAWLS9/zFOsPOBbZjgeq
94+vPiANJK4Io/P2wvHPMZC2G5JoQAzROSakDu/BSjrO7bPAHqAIv7WkMxLIuZNa
5Q7G0/CUUtdbJbIrjOzglf3FaCUAJ3rPfiCKhE9ahbzVl+u3Lg5LWTu68rFxNUgE
1XH9WVTsL/IwF+LSKK1hQZBIMaJFsQTxSO/5lVcrXWq9vDmmySLyiyZeLQBFcR53
URaR2PtK1rr3iU6Eq8NknWFvLBpg6s4CCfUR62oshAs4/0OQocOvHUDIKookgZu9
fXRMCdnKhKJ0Fsz89fnwdqWvcE+h31MfdtIJZPbRVXuvHCOiCKvYNZ0BsJiPz6Pv
90F1CUVyhSLRtlDPOIYT5rf4WrqHUkfeCBGrup5XHn0guo4Chria94jRwyAAMxqx
9VwnuqDV5FYst8xfB0mIcOrCdKipvIKjkwy+k6wujqv+0y4mqt6//0CYC9T8qEAl
dz4BLdZBIxBOfRrRmhYVWwDT41Fxsm7ftL/u/tt7Q0mWWFrJpUNAH9Qi0w9fJupE
GKEK2P1waerQ0NWqxuEKssjJug5CX38/IRubpI6fVg6VLdXQnIWXDuiFpycdQRsK
wV/Ll/64+NRl3O83/uJmyqqlN6Nx+mdsl0Hpkxry6ay+rgmO/X1DwXSsPly21onR
VRkNb1e023qIW62G2h9alq+qX4KIAOaHK6KNFnD65kia+9uWhwc5RJPzKc5lSHPV
G/BuwnJOKMQOLBbSY/KXOPHuTpdHp1TwpvW+9KyRIpk8XSqRaYvoB+1HyDonCIaG
I+uMJKG3Fjy0OJqa78/jbG3U9gEH9+qlRrg3BOJpdrjgFreDBFTVuiiI45D9O6IJ
npOYtP5UGt0ylTPuiJGORixjGxliaSqXXX+md7F4nWQsPmDGcchG9Z1yc2wUVaNn
6UepCTBnzWf5LKQboc0064goI8oWKbFyzb+4AS+qzvSqiF+fHMHEw1YJSRUNJK8Q
dkvuesXW0xKAYS9RCI1tRugR3XYE8qXQJ6eCWKwUxjX5OQ4b1DWFPjp1WYgSFLVv
ytYNiFT29ZD6WXcZE6pm2N/3kODGH/lq7PSSy/kjHfDJ9rNlfl1UjfP7zRqhTZmA
FiYCxjuQMk5wA3xTYNqjnyexnLgtyNVzqPAw3lCt41eSFl3VITZk/cWWw3j55A/j
nsf6lyQeVxGULX3MwcHTRuq1Ahkgi9ammpHNVk48X749CZejTXJbJfTbHJer/yWx
yI4pmCwbRz3vFxl24hcnW7SN7SdgHGJmpHbYSiFZxFikhTQZgpNhuwiOYItvSd6/
UK03IBjMX4B2bE1LkjtDXrFPLkwfL3bEsn/5sSYZfp8H9xDXgPMNkaXeHE6SP0o5
l0RJ0w6MB1W+FbV0xj+67BnntOyWlhMI486JXzIlV3kyd9KJBEjA47C0OXC9qK3f
FUY8S/cSWGdFkYD212wNTrFYUzqsfe8e8RsWg4bUqrkMmYv7DO7GURl0JZesj4Uq
ozrcij7j4AXeJdXZVUxXlNB7ClpFq/m6s8CvBAIZRU8z8ZuH1K3d6U7xSNiYBBO7
sZFZbOeBVwggRKvSRR8wxBAA9sytTMJrF9LjAvU22efr7LrZum6C/odjgctliEnR
inYTUjCJj62J7xWEPR6JL8WO92tmu3M0s145ZEOgOcab8J4PIOnma5D8f7WQbihn
ziyyTRsPK3YKpmpA84hnvp7ApmpVupqTSNjIw4h0Hshges13iuXmk0JOlPp5KtyR
b3filjgQO3He7x8Gucv7m/G1nI1i7zrK9WHBuH37AEaGKIHCkP5lV07e95jFKeHK
Jasq0JgRUOjYiV2Fm/Zem3JTx/VSuEqlRou2L4FF8t49GsjfKIolfP5J9tcYzYcN
liM21G6hJ9RXS5D6Bgsxo3vvcqpPru0E8VjCXbBFTzVRmdbdkXlXG9iNhQwIozV/
LHUWR3RR7QlT/d3dm7sBjFcmQCP6oq2+ivjAzXKKM+1QHSmYRozJhUpOs7tQRe+m
GaEF50slc65vkmQxwBhJEanzUivoaeOp+2oFxHoq/GoxwdGt24OL8+ZldFWiX5dw
3LFzNRzvB6TGmXmp6bm6wKMDoQZyb+l8WtN6FsBbVgFJzwT+HyQtR0tHhevYppAK
b3s9oHbWiRoBoeEVu4oBi3liXzwlXrbzg3LcE8/BKis7KffBAW679W3olM0qNvJg
MbVcxiD3CP2Bgo+QqelWIl+WHUlpo49k+aXX0oW2MaCkVWpsz+Wq9nq6EX0YBkNi
6QEpOYoVZAjK1waBRKchr/0pUVq6i8Qr2V8jG+11ZcwxiQC3dGBDCXZ3rqC1yG37
MThIB1vxzJ25d+el2FSBMMGvV9ERkZx5GBC/gYRgSFNIAVWLPxedG7eHvznjWhra
R/ljTlMw/t5hl2hlcNh/fsMksL3M3y6bT1LUEIB6Y0g7+0HrW8Q90iBcXsf9sXeW
RGZ1I1TAEiWwXIFCsfeURVxe3yiDVhois58cJNWwStlc7fuoWy0xylh1LDj/8Mtj
EtBY+dZxhktQlCF6Lj6qqKJ3L1KivVwu07fnScL+GoYQJNPO4ZIu0ynJGLyNFA5Q
W4LsnaavQs1G+h4p88cSSXIT8AHO9XvJuFrYS1ziHuB8j4bh+7Yqhb3+LbB/QBiD
SFgrp9oAEbKEu49typCD64NCo2+ijRkl/9Um666jdHOhQ+WeXCyCco87mALwS2mE
aO3Mdp5T3vcMhNQvGtPzPO8qF+kZIzWcCFwzepJ1JAfVAN3WghArk2YTvaogmkCx
ivLz5jN0W0Z9c0If0F1AVyWhVr9UAV1FWRR1DE7NTvtu+MBcq+cJrKOqFNMlKZGJ
Qz1iPOf5xbpydbfngMmq4+bSQYE4h0dTKcm1ksxQBR1XDztQASdNv6siYHFiTzuI
2N+u93wB1arAi6CvYbubuQEiW6xzimN2gNRWH0m1XHfQ32BjQc/A1QABIr/QM/xm
yxmTJYaPkgwcDZW9NQ5G/jNEcbI5Iw9sCWPthMnBzH8sTNQMfVgc4huicilDCjSu
wDlUj1V3cUlbqkrEKDTNnEeSB/G2aqlegPAAx+Ln589I888CuXjmitHGZZo3+lv6
+pxU/8EKpn1xdEr5NKBq2otayShbHTneWW+HCX1KvYuPPYualaJkboYpAelTYau0
CXEi7vEu9/VBjzYjkPMy5NnEh+CuBDyt6gwBitp6NpwA7j55Wj9UBoGHCf0KIJdc
rNvcGqSW0y0UzgSasSdChQPV29NLGMRT+KgfpkcvZHNI6zRcWvaf5q+uDLFNl2oJ
jnqBhwTnI2xxt/+zg6SoBmP7JDiJyvHWl+EuMHXbZPqFqpx8OWOydwZxYpl9b95W
wgVkoEIQrIPxxDNsI05H3uDIQF8Fz+l3tCCXmfKLqalC5w5Cz4PC3xMPWwdiafnf
E4seVQ7ELAZz4PGxALSdobga52eyV40sG5ndNxbHVYW/JcgTcniG5Zlck1uvFx5j
MCiEhlbUyILw3nxxBsybldkCTCy13VLxbJZtQ42eipcb8TEKXcQ3EYtCKexWJrQg
VKPAsByvCnOsG8kS0/bcAQCfvL9dGurp7vjrkLTeL0zabF3mPSvOvPNG7ppGQaD7
sa7kL1/G3KDf8YFEUcOzUEkvSrn3n3MxM+p0SWclPxR1cnSX4cXwvZGjn7Febh9j
7mpnXQWA06zVC0Gpy3BDO273F6giyvKVSgZ3Nyptj1VRdwEn0wGWYC84NggjfsDz
NHpI6s2k/YFdrAI/HgaaARo3AaZNZt4LzivIqrm/yvygas4NNOoDySdW2KuaK9q8
fM+klBsdL85V1akNNGV6k7oR8KjOoS0XWSb8FCjo6izvZpr7CZts+h/zn0K0Xwsx
FukFfXZWVl5XifzoNTOJYbDB7IREg6wrcvnh7JbkqHBKHgkowrn6RTU9h3X37+FN
D54pOzzPDQ8yBX2eJmdgfFlzC1zf+YNerEqGqz4QQnwAcCHb8RGx5/gVctFikg8u
J4lMUyK/vg3a/nswpl2h/KaZbPyFWS+7ljY6O1u78wAbQ9h4lWRxK5PmYvRmBF1F
mwJNC87CgjmGWJyPjHscph2M0KAp+I7ApO4xoHbSXcL9b6V0sOB4hmEz8sdnIhxN
X17v/XUCSABBLh+jLQfpqDj3H86hWvMUNLUUlJMkJ+0T+TbNX3dKJHZratLjxyVg
P6nlzf8jlWY+yWdjCnnQNTXtcSlfzQdBme2FK2Bc0AQyfNcCmMfJQTRBCAY/NYJ2
p/mQGiPFGv60SmkFbyLXOqUwP/C3aRoSmcWYxaAOdwXJlKTMDW4Ft9JZx1xCgvwQ
SuMepRk7X4NzWFBy9f5mvdBwajqWqLau5syNR3YSJAKZV7mTsmRrZ/rtDIF+pwTD
tG1GcwxkG9/7Kgvk1bZswPTeESG01LQ3w3mBYfrZ+7e/BPGTrW0I0gXQT053NCoG
sNr9/gG2f8g8bjTJhBEr62ocm76XtMn9atGnxWoiDJRXpaS/c8fomquQOBnq9Jcn
QFBNWJDaUgsmsXo15O/bW0Qd64SUo6J3paI7jUwkjtwR9uVu/bv30HAt0j5YbsWJ
the2vg/fFC48jeMSrqcDdcSGvlfGgiTeViQ1QW6iOzCz+45Y1VhhfZ0hnpbjm/PS
scTkROACtmcO4DBM+gvudD2dKkPZBC7+L1rwt31eDZXK25oDVSBk72U59ncJKykw
uDymcNOBWfQ7kOQJet8eadfVbRVlBVwBynaLuI9hMtqqNvKYfKXihp9XnCLlQJN6
NEWGuMmDp5DzJ4qnVcO7YmfR+zKR44HZ6YbO9J9lVVPztysKwSpPYVcLcKyOs992
diOLtM+USUAQ/O4aKMJIV1YVMe1SbnnItBOJvLw/NNyWx/CNFPn8ud5yk6Sf3Fii
s+DSKMNLrrKFhV4j2wuLp4FcLadLErGjobu7TZk0QYkZDkX/rOHA5IjlhAxCAns5
N7vT5L6Jgq3ldnrURg7dDuPOUUmJZd6bI4yZP/SMawpmdR56JEy/vC9E0f+/WrYu
XJhD7luEhsnz9B7P+PPI2PW79gZNCNTMnzCu6nxJihf1nQPMFpRyVC9jlusxc6Me
dzbH8xwiiK7Tr7Rz7LJqt3CVA4PmzzCDATwJHehKIkJRHiHLskbGo8pY4HZaPCAd
Qj6hjFglEJYynEid9wYFHYtiyAfrsvQhf/ltP02wAnfPnm9V4zU7NaI0hmeEWBFr
JF8h3p5+u3l0CC182Z8nTOEcZdJyOomzvLvsTEbwHrqc0b5vOayehZP41Z6aa9PP
cikqczYVW1jolPUjx2h8IZXUF4URqycHQJUyHLn2eWMIdmZX95XzT00KGni7eB7I
wcWiwfg8udBTJBr1YXCzQiKapwowjigj9zpstInKNXba2Er0+a7+pkSysTYPZil5
sa7v/r5zXxL9dpHNpIjGoDhpSA9c78GIsHXzacz2Jz5BXsJvylVd4joLsoItk3K8
+KjZDoRdMvggRdegtbkhmMOnzEn/eQArnw9fpR+64WDTzB9gtOc2vT0KZBliiN+e
LdQ1/YDQIweXxhMqSbFdBRLrOOzCdXHTzNzQj2/5WUWH6RmhSqiZ6f+5h8aStuJG
nluZPTVnnDVoquxdDBCVrclNA/U9CQhMxIRS5HFiVReG0GtNNP/Zbr2Rji9LeTqs
E7g4G1HNrBsyyVTpVtSE4yIZ+tRTzQ0Eg70IR10gf+fQGHrZdfuol1OBwn3BYzlp
mebbo/vWbPQTui2GoL9Ew5ogrx7/uvOSBqvmwKY55iU79Ugso2u/KqoBFQ5iZ3eC
O62XHudVxtsoREeyr8Xfc1hgRynYGoBfF53BMzGUz8trDp2qMxLt3TzWA6AMlCS7
MzNBIOArS7/aVxorF0F3qg==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bTtDKbRZVjr/tPR+ocbJ6CIf1ngJkuzO6cwwxEjCYlsphcDCxOCqF8pX7DTuM99z
HXNNnfecg8sL3WKZYmjP8Ur9rfwqmJaEDyBg6s/1nENdZL2s9eV+N/3pRfNSx00g
uIH4ERAp31CRdnefZHh3F0+lpPwNv6+lAXq1mjvfJ4XktYtAn+l+7HcO4WSZpUvd
jO+YJgqLhTK0XZDioPh+K9Ej0kxNb4SZhf8FyEACBelqo1KM/eJGUlVHmrtfN86B
bvMSvvoEezdK2z9fzA8vOtwpngody00Qe+6lwXlXeooLGsBIzxTD3Xbs352AuOHc
aeJ05oucO6VdmIkzoNLfOA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2016 )
`pragma protect data_block
qYNMqnBMvkARXUkTdYCJ8rG0KHAC4xH3ghPlX43lIyYXcFRAGuvw9hmchGJGUJcN
qNsImWDA+XPqm2QiQR1dcqgj7vBPMZadna4B3DWQa85ZZrrr1rxy3HRdA0Stz8h4
4Y6fH+/K5AMGNulFPf4zSfBpbOaitUu7GcpIjhVwQNOWFsG8Bc1sBRm4tn/J6EMQ
28NsJ0OdVTztw4v2HmwjqNe+kQvn9kIrJzPg+RFhCJOL4NczY5cO6PwQ4V4ZI/c7
Cu9wm1K0Nl+mUwx9qpsyl8GPkwTBiVYWi9pjX801hMGFAFSFW5kl4IO3KrLqbfpU
Pl4SzIB6Zf3SnUh4Jt9rLE+x2lZVDKjjeeFos6bR+pgkjCEnNzrhjy7/8MU05L/+
iXvv/w1PwMRP72l2cyZpDxMO4e1oAvgoIT4oD7FjeHINEiPT8m9hnjhMO0BbXh/A
TaQ4pAPwWZgtnX/QcowUtl4wi4ebmS83qOqCOI4SacCo/+dAEd8EumwnNny3bFnt
DD1bNCpo6CzznOzyMgid6i3VB7MMsxS76/U4JzhMK14iMJvWJ8hMayNSfDJpwIf7
yA2Z5Jmbe0pgh3mHTMb72iR0yqd30mUovKwBL6PNXXR8vB5tOM3KdGpACdgK/0ZH
vcKONv7UVNteCBEM03Rd8Q3ZKM/1ZHn7oGa1CAkQo2SIx2pX4EkBKdpkdCEyFgde
PD/t5jLBsCBohL3WxPivBepOCz1SzbfcsdKrPmWxzm+Ql5kp19BEngiOI8ZXrd6a
1HzWdbes2AtgRZyoc0GFI95Y9gKo6X4B8IAXdH7Tla8B78OWkJL/PLN8iOyD5BEH
kn+YEDCO281sdWbOy3dw1kIW+tv1m9PuypIWqgVGfYYw+7KGB5ii2tQQ0ejaRq2T
Sl6X68qPZR2W0dBFdKyu6+EdZGRuGsH62N8LfGKW8z6UEVO1/QbTNvQoF5sigAUB
18yTGLqB6IDOzcJx2cyXMsQfyr0dPAczwof1UUd+K6rrnZ8C5AmadvjmZe3GYQ4R
FwdwIbp90sHqsCoNnitqTAyUDuCavkIcZCfca0BixMiFsAkwA7u4NjbmI/5PHKo0
KUB6zey/W4X3QLmD+byFQrNkFpf7P8YNHH7QGQ69UyXdSE+6b2TMk1+BJruNep6h
tIhSn3pqQHma6QMLiwYOgdnw3EGPAiI9FZwU9idpQ3Yx1edYXKCicfeaPwKjeu+c
mFvp+ZXVjI3mIna49TFSHlYtuffWHCrz4LK48uo3LiNfqYn86Uxpb9W18kBCDgQF
8M4YRewXxpbUXutnFg+BDnSgD+wnRZJcFcJWyPqtVl//uVgXXOuemeIhunRatpUk
k/T7zAx+mpYJhblE7ccTaDM/Ll/9WySCW+aHoaEuYXBefjx1LT3PWbe4RZXyyS7K
z2KecW5UQJj8NpNhXirVNESn/e3LUCfNJ1KQgWG5JdA1G8K5x3OQC3kFcTgMh8py
ly+Qi3JBVRSjNeLEbaGOinKMp3h+UXhvG2rQSy2G3w++YIdBYhbpGzUWLF9nrB9C
fgPzU4wtibMzKFkvULqdT1BPAOXqpeH6iPsDXhu/AnsnVmwSpw6tWrTNkMHZdIr7
WTy8yH/e3NNXY+MTMghWhBlvMMkD4S+wrq76ZneZ3R7oLYWZfIN9C5+R62XDZrMi
j7tJLXKD944N1pn1plm0YeMF56M6J7dv0cp7PUaj+3ozOlw1Kcyyz5nrgUTxg+Hi
PFehbL9s60fFAaGmNvvQjctxQ4Cyvg6uXHocAMpaAGdx3VkBm54c50Ca3NeL6IEz
8AsmwrPtVDF6+XZrvIrXwx/DCqPh8HXtnSkQTwj/Ko2phVDNpjnwJLBZvYRPnU4R
tiqkJ/kfjpydjLhLiXC/VN9RwD6nlWxu5izYLhas7ZXP2l/JnAknhIboHJW/6r4D
a5L9ykupPr0XviAqv2FSaGavKYekGY41MSODtrr916J6x3NL4m3yxj+9d4Gj7GBE
NJwZI6IzlkHuf52tlMQFCw7Y5KXXl2fqXNBl9uU4Z0Mox35Xcsj8HGhLLb8xnOjI
8wZsynDFZ+PjWJw3vKAfXezjlGwSoV7Kirnb22G9bcd3o9CHi1DAy97yYeyowHF2
IeFFAhwddLHLd0tu9/lNmqQU7R4M4mRIuQeZskyg2NBvaWw16UL0AKURIiCBZK+O
VCyJ7NrmtLn1hGbCQoFqH9oiem88Pk1riXF/T1WYuz/dcwetL0y8m7va/eddvUe0
dBy2P5bHPPKn2d7ve3WRCGQlrKdEqFx4pQUBChlIvlvRj8NOdnsNuFun4dNdhXAu
5xF8NxTlNVqWv2EIViX9ibqL7VieovJVkCLYDvu/g3iDzVQiFHlPMOA6al2jKLou
Nt03/6vvMOE1kKRcoj7ftp0oSQzspu/XFS55TmB6TxLP8xGzfKmyC39keo9WQOTn
14d0+REx35XXjMhjR9A5fW+hFHFEPeZbCUx74cGlbfR62Xr+BQLeW+Jlw0jqJKez
rfPnZUA2RqmFXy2JVP9eMpmFSMxH2eFncy7oC0otGsWnFDWlQLaSA1ohyKBdOoIJ
4NXfuU7x5mFjcN9EcPlCXhEdk+BFcOsT3FK05lo94rHSiLII9U6ssne76CgXcpkD
DchhGsIVQdn5lyV39IpXVsoTp/sZH2za8q1eI9B2ReanWXNFxTvuuo2Q0kWu+joY
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SIddslL2qY0SdO0i1KAygOTsgNXYoB7vJ7CDav4t9LA3m/1T1nfSShaSg3WiKuDd
F14Wepybks/zfKksui72ubcMq8H4mxxydiOzwLKDgfWgBJK4LoSn5dRGlv++i8Po
N3cXTUNLOHDUwGiVspkLfy4+8foo58R6FhIY6qqW5swGmWXzLj3a/72vojfrptDR
KiiOhGxSChXCrCZ7V2yvA5sgzi3Vj3Vs6RZocORlcoBLb0suBwi5s4F8W0CWI/je
JrUZesufoyhQDc0tFdpPhM6VSj2Z8gKpAnafaMSu75N/P0rTzC26qgsioe9S5+zq
BHY9xCJyAAvOtHWmTmrErg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10976 )
`pragma protect data_block
UoOd6UEYBaAhx9IncwN+GSlvj/7BLqA9WZUwYi02WkhaKF4V40QznALrQhT5sxQU
itEpPwpodiPLej8daAb9Nb9esVHA+egE7LOYcOnywcJV5+Gh1EyhhQhxzTWhOHRG
nmusZtVzSpiEgc2l8AycbBx0cNFB8Sum955xyXaVxB9rMGTedOgBd/bunC/qw5+n
QBnzSVmnpj81y2uiCVXRQVcqA9DscknJ26SXOpLk5i7zoc1f5XjDIFxfo7ZB1wUo
4IB0PlbapUztgDFV7MWjQWEya7vbjPlLKa0ioj6oMDQfrboE9cfoKihaywC0ABwD
7jnLJpPPlIqDY4HZ9Ds9L+i1tIPxxon/wVlpuQpoju6oVkVNpofiSwO5zkdjBsxn
CAks3m8ApZCcyS2BiS3bHdY/FfffoOfz7LvYRXylIH2s6U9SedWOgb2XIrK9vmqD
Q1ulZMmcqolrYNGKN9ahKvsI4K2Qh3/mz1qSibxpUi5EtWqrUhi9zpg1Y6cXtRhE
yO62RV2mDvwuszZFaZmFjxwVgS1qqLwqib8w4ZliSQtTrORb9dyeb4Xz0ve2ckPy
UmNDqpyH5yypVnJyo4MNfRYRErtd/1Xa4gqPUTMBoC6CFwnueCVuoWIBltBrEGhi
n5fVHoxwfkHx5ct/VFqbrYET2PJkD+r1qYcwLbgU4wnEtRaZHtrlEcEbyrVvfYvt
Ju/Rc0NVKMC9SibZHQliYfXpLU86YglMwwU3KE1j6sZGj114/cUVtQv/tZPwJsIp
GDmo7TYEEjJXFEooKrazbuRLbmE7OEZTEZzw4WRcLFkHY5Gn8BEVsLKNgRJmu9/K
3YGwjbGqhHrZNlJlCN5x8tQ77UmEzHqVrPyHFuVEChGggWsJ+aNuOncI5aEDJGt0
ve37ipMIsj4ZWWFCitbUsPb7qBjfzKCRGMbng5ILR5XjwkfJbSDVmT7EKh1fOjuR
1N4rW4rwUi70n446ZzoOl/orLR8evClUKGDm8zSvrhtFcfqGpy1hBYS3jBMBz+v7
/FG+jHxVEkD3CnagYTKmvvP7p9usrmYYTxXGY9pHSXu6yrkQVIlkquthnPFxz1XA
9IllgR+uyjk+mAYBG+43bSIsAvU7LUaKK8rD/63qF9i9oaMTL7/NzjjaSHjOwNBV
97wk+ZpwCLI51iZjGlqoBN0Nfqlw1RjjHMIsF265hrLVtjm4H2DuNCeiip+/btlK
lQrs3znQYQtF5VxQZHU+JMlKs9OQRsuQZLF3fJf1lFMb3KDRRhkrl2MDgkQJuRZe
rFRXGkaZurFzBmwgl4BZa9aEpnY8uUmzDCi4fs4gBmI/rYvZzT/UpYBB3DANG2+P
3t7NvUWBQkAFSKxQ/PcqBO+onoLbFX6JLZ+pgACyV83F5be58gDxmDL+D+H2DIX1
D45m49s7wqBjnX5apRdhYdjPzZMSpYe9L8b+cuCkpyD27pFXueH7O1Xm21rDLGYn
SejppvHPqn36TATbMuoQWssa7eVjID967qJR9PLz1p+jSwuSu8Vy1fkjsbxn5/x9
tFc0/0zWFIA++x2J/UT9WSIOs0qeJU328b2dPGNUJ+Qfmd8A6aKTWd4RrqsuKGBw
iIlyEgJZTdEkgiWejAWFFGxnpN5dUYUzllJDSO+MJU6jLjDLn7rqQqjN6Km3IFJX
vJv0Y8LygoIDozUPEslD5Tegyp/ZazMNi9jS5JOrmliP2A1cJ6mXqrVDmThvd6zM
B0jeNxlSIOQ0gs55wvruVHJEfTqXtoJUrLntZ8dOBVHnvOfCeQQto2PLIxz5eb5f
qokBCjONrXYfAcWAjKgPjgS4i+UCU3CCz2P/IzTgqGHI9LThTSjoqUK/3pxEfYri
1lDw33FXV2IPgGnKuUi4WzBwSo9maiSaNSgxbvo74ne+QwGWR2DHbQYVfCNA7pOY
FfPuZWK2VlNa923B0ZfZy4AB9ufZFIANTmaBGaopQTBlVIhqLyK59hRZSIZ+NrOO
bxccU5iCliD+kJbB76h7YWgiWpqmqrM01ZKUk9qt+h28u5vuTkGACe+WXvSTgJ+9
gTCsJyrRh1/J2dLNyUB8eySmv5WNwQZSPbK9QT7+GzEtsN4AppmXP94zmNYHzLqp
G4HBcGT3NBXwOVio9Ml5u5KBTKKgFqgyzXJFBsnv/OTypGgZuMaHuG2hqfb7Lf8Q
cxirbZZJ+vcrhoqUz2p4uvn2ASBPxkHoeDDc1dS6bKMIUxMfN88K6TU3r0cWMsrP
oeDkaM890Mr87DnaTV4Ap4vfsUaLEdyDeGj1LH8ht9f/2NzlBxI5cUtOnQbrhCUX
D+GWx5PmDtb4ssmX7lhTzut/aSoJRsxspc5LiERDANSfNg0Rt5s5G0loYdO9gBNo
93IU0UvQi2inBM56sMLLdJLtHz9DxnGom3GazQKdQgUz3J3pK6MT9owIfHnorUHS
zH7OuGdrcm+LebjfffUfwhhlar/g1YociPkPlRrih1ceV4W3zQ2U56dYlHyRvj7l
khfI3QIVgXC/UT/XiiObjDEUX38LCTeaKVwOzpawywP5cmIbHLRfngB79TsZnZGQ
oswLEnfnYwH4xIFTbep+Xv71hSZhyzhWmILc8BLaoUFHIxehgOn5ydbXobPH4LCA
6nj/RqclQFnrN2s6AEa1WdQfN6dcIB1fp7iGPOjZ+Te9iPcF6iCvu/zD0wUJ4glE
1HrCz4WLV/5QqvUOOXxd9XIDUKIfmuOhDlqVZZVJprdVQW5f6h83g/1FbRDuVAoI
r7Iau4py3vK5CJy2MD5uBK/YK+hlzhpTwd0k3WTyNi03mf/rOmOUrgqMQXR1WIds
ywvvO101PQBnNPAN+hh0aR6HTW78IWn2WiESINp1i4SAwMR35W7NbkRNkyhyMvvQ
tT8+hcm+StG56ybI3Vypo7Ok+EyCbw9LQ5Jl7+hQRYam2Ifqpu03KDLgvr3qpMv+
k85mPrNgKhBWvTNUZef+ZyeHx6exC8HdvE//1WhdQ60ClN0KhzMK5YWkBaBTLyHt
TN0F59PzWHkSry6vbC5TbqwyME/kkqvt0ACoodaaatIjS/CULx23uNmtaT8LZxLe
nQ4yWjwylLl86Yvcmj72yuF7g37UMBw6ppLIagvSJWGPhZzxINgJaFxfeBu4+3kj
/tx2G6L9wGDzfQD0TVElNtar6wEssEy3Ej/CZ6e+eu4DoneFON9Mp6CWeW0jCCnG
grKQySBSUpxTI1QH8PkKHFas76WGhlCxr7T3RbcffEl37m3PVUUWMdGHu82Jn6wk
/wQ0l+co098vxbQfhbCpYrwBQFPzyy7vf6oOczQXJ0lRsMnEeEx1/+pSob3X5LUf
kWVLM350gFzIpxC2qOYI6pqTWAsAFJ4BjI2bPIJJMXcbBnUfhuw2vm8I7VhbQP85
Z6SQUkzDcEpG7jgwnSxSvuAKbphh0mBNWi8CVlTgXWJL0z2m3fq7K8jxpnLG6mef
Uj8EgFMy+XzKKnEmTynNEh9hk1e5cGxXcI1zQG+aXbotSuZBJh1mriOtj/4raXTe
qA7IAzRRyNyXWYKM/ak2oXJrqaXEnLvTUQhO5FJr/tiyr8WhNyDdpxIhqRptc5bq
sEcWNiAOGbQ8aoAqOotWWg7ZLKNBUtWfxMdgoNolUm4FBEcpXpikjPmj+s2fZm7J
/12xxkC4eqCDRpv6tfbqxQo6Vo0FDnC8NBDcHMa2uVxQvCg9UH30MKTCFUAJggN1
PVKqmsbSU9URB2AWWWdWfoIs2N0tnR3jFbAMV9i8Yi/5ssOMr2FJw4L+AW7TH4BJ
7y3J1mBxwusfZn42DJdb7iSZkrzSYB3dQ+9KDdPmPMQQQ9CuEPZSOnSZf/gQHEj7
2tNNwdJo8Upt9EkJHvvSTx9EJvxrqhR92eTu4zDsHTNo1fEnTO56e5S6d2MeFU1K
QkSf1pFltAdw9Y66J8JPN89hAE2bCtngYYq7BseuADnmHAzzlqQSY9aViIIqCNZR
dBSlcPwbsyxf/cokTuT5bNgRNvQ/79yoxrN6RJuB1UfExM1Eapb3+d1UvhhMzf5E
OtbUhoGnA17Zr7Gvc9hE5pgNMhLxv1cB+Z0mHi77E8l9DMZ7oo1oPiSVFYWmZxqo
t6N1QaUptCFsMC025Xipfg+rAErkYtoTTaWU8nCeJmoNitCTCZ9S67K3sVnr0R5v
xaATz3rnKVmZ5siQQ+bEmpUXU+/D+rIMv0tVe76OwQfBEJ7wQcaFdpxLMCWvtsi/
Xcm3ZawOdO4Lu8FUI8e248aya5ixmHwqDQKS3cL6ihsrHlRiFc6YUGFzPM7oQ0AM
2NfkaYfKeJVhlGUk/kKhtr7rmcZNOJ4jsMbu18K3bqWiDwmQgYQmnG7rpAfACazc
QzL8E9kA+EwwjeeAvvSKvWX4ip9o8WDNFGFboS7NSWb2UxypIuYceIsayUPit4im
klZFX0/ClHxkNOGpse0HB2Qpo6MhcS5wg+lSRkrdLDXk9plFFsuVlUXuPat9Inif
EEoQ962yMemSkpqqPr5DsGPHvFAcB+R/K9EzrB+ko0emrHOWS9TH/diaY0jt4SfZ
Mwf+mDjWJUnVjN5shTJKmv3fCh5SbEhgVx9kzXgBA42QlxJzT22UghhlDlXXEgcN
JDj2WlLjSltEWcghykXVfCJ3ckmgrNphHvSU171OwK44B9TewL2fBLcohPsfcAG4
DRD2tZBT8mf3mDS+WMfb7Ve6Pd2RbAvYAEFGKiYpM6BpT6ojQxd91Q/VE5G+WUpl
vZ1d1kbRoySroo74rgpMaIBjcnhkg/lCwg5pYjuVOtFBBLWDsc19qGOYWmI6NZLz
1D7kyJZAhrxiqJ5ifSpUTwZYSijHgAN0EhB18DX1HyPt2VEYTN6Xgd88f33B3yC8
Pf7kgPqVuuC56N6tVc/ZJuj27yAdQpVv3o/ruC/VZ9M81S6vn9lLyGiwB5dQ9Hm3
NMf6ia2DlDK5YRybWdk5bj80Ct8W/xQDCbjXgv6GIvlatSipjIzM1Ap0tyRfVmwM
Q6VBQMmLM0DL3kpS4d7+s+vFJxgHr7RfWgz/6P1avfXOiyghSmtoBkHiYPX+xBO1
vt4kENXLqkXYIHfjx2LvecgTlhV2el5SHdlB0jORcbg1dQUP19OdTj0b9ZvS5uXk
rBgzTQpt769BCLqzGWIy/8oum41zYVP3Celco+dEb863uYK/Vp5XjvA+xpsAUbcG
sqtbVvlwGWlTOiWYPNCUO9oB1GST9uY7VfUjzS+2cBnTHY6S61npe2ye9h6u763s
bAgNgBhx1hLZsLU+DSzrF6v9DnyKHcy/CxuBfksHi3EuyUx0NbDi4rT9Vo5x8m0R
jw3IEXU+VcimBnwvK6s668oqv1bIfbgTq/XY5bD6ZOV4ekvOWnqvuq/iUyVo+C32
olyfVfGiBu9s0pvhz2ojY2YXr9pC26JGACj1dMnXDCjzMC23LxIVJbWAENHvKLeb
0wid6mARdK8Bna8lDg21gUU8Z0uBT0QXI8Fp/uJvuD9gpEG5zQMyyIXpZ91ZeDwc
Y+gOezgxYCgKHH1gh2OUQeufYXafAc/vpvg/tKTEmsVmmao1yEIoD8P2yvnIb2xU
C0tzg021AfJUerpgf5sPYlWEYjzUULI7r/Q85QVh03Obur5YNisbfiTaHp6/SdEF
7rPXdWwYeAFz1kN3jWtIOa5bL7ovC5WUyAIIHFhgJMicApVcQ6i6kKCUwA1cEIw3
/QtywJhNCSYYToNuMiZJ5IJeAWMEjdnTOcqHg3JljWzlLrTviFZYcE9yZILqac9Q
CBlNhNwZ7lqoefmeARTG+HsbjC7skQrb3oWg1urdzh3PGX+/W9h36EpmAeq89s4+
PTdnTn5Xx7WnBvGNSAJ8fEf63WfDKQF2dRvLaTUhesh+1h6HzAcuwmO7+jU1WbsD
PNaCCLK6ZVjFOeycES7hTSZdWf5WdL+ehZA2ukGR5o44c4I/xYADcDGpEl3LXQ8U
2GtymfEsLtint+dU4gV1fZmP8yPWWolyd2B9IjQpbCxT8lStfHqbpfC2RqAd8h8D
AU3sofckqN3EMXBq+/GOgL7GQ7a/dJHQgmmngOYNMx3nMN3GrtEDKLt4CfUju3vA
SOTTQkYGOHvJGCgCDgq9ta7m9kAHSfmSyKfUL5BieMvmblhCT9Akkuo6Ix7DTiwx
trLASSX5MhkS9srGTAtcd5pKAxpbWIKZBkOrPS2AniMXDYYeCjxPOauLi2PB3iqH
FnM7cot4Ni93sAd18+iya3dnR0ITXuuEJQofxsMecBPaA4+Xh7cWYmKEz9MPnjK5
ZvaMxtD6+Hg3U4VxmcfV4KVQOcyBganQ3WdyTGvXsVqt047dFYy1PqUylOWXrpq2
2hfA5UK/JG6JWloTSaW/edVahbJh2H32U6oYnxY8XvuYPL1d2zeqiQxfBQrKYnvK
tg9CsypMur3dSfNtxu2KnnrXDtiYbXxAuMGOyjUnpPei5wiV0oTH2ARZ2pg8KuCy
2UA2m7IBQnHamVyREi5TKL/XBi9zjFdlFb7d/7MfjR3sA8gJezDUAMdGi2ZIR4JA
My/ggB0YT2WBHHhx2PlGSLvPaP/Y+4l2J7kbLE7Q9GQ2vqe6ZyMphycHjGWHlOtz
Jqgoi5CSKccaL92NhKxHB7mcK5TdTgX2gylCavQRG/WwMnErdT9oY26pflBhYhqN
vVbwe2at6qVblsUX+NvzVFLHx2O+VTwlRdrWtXLn/qPI2IuJf0jJRY+fxDh/9GzJ
QIH4jX7vhA4Oikv1PnQJd5LKrvnCwV/v/BFZarQHLlQuofuXT44nQkZWf/1EuEq1
RGyBb4YRGLmWBBBHwsdGv723/Y9wfLvk2Lj72szRdvTIhnFjCkjggyTI/q++0ghK
jeI16hdhHXfhAVVYVhB0yzQkSWH9BBHKb2lNHzwkDk5byphNNHJGNnRREYnOVZHj
nAI/rIaS3DHk1KkkKy2PDii09BEcmEkMJ4Wr52vHJAIpNwqCsaDDOkcr1GRhkfpd
9cQEFtl4Ij9n9Xlohz30JxsIQat8lYNLrUb62xZQNJ7iH1NmpRgeMHntQqYb6z72
8FxQ5EZ9REWZw83abFuED8YthJCBo/l4Iiw3BD2Zvvmi/LMkEXFqjC5lj5j19hHW
B8RQCfDUJnGOaN79sz+uUn0MxAo+oEpCBQBjMQrRyJqjTG08EDJavJVvYL3VHZJK
3BPILRzZHDL69/FnhWQ9bMTnsDZko9J+gkmcYnpApzdLYd9i8BE6T04hXenEeEUa
O+4y1uoPMzuVwVpmg0uq96gLeH8VWkVAcyyjeSk1J0FyYpKiMHryr21dPUwv6gH7
8fE4h4KHKaMEOWT7njThudph37eHOs8XAsDS2If/qo2pjn15bk8R9Y+6A8fTBT2s
A49cBIbs7SxatdTPDlHQ2koWfUsaNO3kbTVqTc8e7x5ItOMwuCgGpTgr8az4688A
k/KZjuAescm4rcTLPsRGsBYWd7R8KV5+tjblmkeV0NNwn+DwQ4OaFfFXKfkk7Ma/
Xmk3Z2T21sl35dusY8lFo53fxyBiQqkkJGRaApyHuDbx+qdnzPSiSxQrAPM5grsa
TJC/IM6SmjqUpsQcv0HV0fh46CFKqc5ebCD4Fdu4fMnTwUglI+rDpcOCm6iCMXaj
qKUKbW9PV4tfbGIjP2KmXeUGPocMgaN/ucm2HA1mYaQUGkiv0xc62aGVZo0oukri
MWJTZkJbj0kASQdMdxrBu7+NPJXwkBmCaGO4EViCBbIypjeVpWS19qwvEDG/SD0D
wY1iSeAY6ebTkb0obM8zU0UHzm8HRp7IAcaewv6pWZfTlivDxr1QGikUjAr+H5Do
v37cLKXPFNOo3IQLgRoPPDIQNjKUPBOHcPXFxzIEqIFQP2FfWTO4BwTqzl7pn43R
1SfaDMES4KLF7u4K6sHvD8jrUpJ5pSjDdx0ySwoRqSTWn7CS92KztzfFA04KpAy4
DRHSKO7lLEXhVadrS8h76tjVpOXkZCEpvbnoY6pQ0rZqbn7cH6TC/93bBt+x0GWI
/BVASIFW5tCCW8lC7Cdmk1flbuYKkHftHxXkCw4+/zLalVw4974Cgh/ctaZ5H2kW
V+EEW00U3EihkpK1bo2Wj8iH23gkYXSeM8w1l6U8FdynilOT4nxagv8TZG9O/zny
mMoGzWNK8JLbkBqYVhgq++wTKmKHt6atAmZ6JnUbSpaJSzvnT2R4hgyB2I9yfC87
kEwBS800+tpdviKRb+WUFfDLwIm+iYBSC6Hxfwvk/ildlqgU8c8PKVLxWtPLUFOH
PXNzpE2/jAEP9D6jAv9nz0Zp+C+zAmx3rj9TOmgZJmSBxTJ8iHS3R/tCJ8l+jyd/
/H0kcYwvYHdaNpbTy2YaMvuoU+jAhcmB2aFsCXH6GzZ/aBE3NWz8G7yP3n7A4ilX
y9bHZ2SgQU3ytavsGlbpw2/JrffbC5sh9q5/fmdZsAyc1qPYN5EN4UPT3cn4NxcQ
bYgNrbc+4VSR2gvDeA/OzXAi1JdQbFsR6P0N2uSxIVcX7JkM0XDmLPoAqw//L3M0
lqmpQIiSPgPCOmYcyAbgv5q24YFP2kuooqLS685YmyrwiMgJKK6YPYP7AdEsdnAM
m4Zg0Cr+StrSjNP96sE1hpa1XzljPQrzB2xYtjT18IWOR/qjcsXyYlUWJCMglHYD
6vFhSctaM21wTEt6r8voFr4bGgH4J12pgvXuAeBtLPvDj5dCsprj4UNxV+jBBdtW
i+WuXqudkMD478A3O+F/5NB1ytbT8jN3iyZv6rwHt48cycP6mxRzZ/ipx+0ph1Ox
neM0gYgIjectuwDBfQvapR6PMAn3ymXRQrxTE91GtuYaTbM6iISQCuX5CD5ShaMK
RA0pGkH9ntceQJfrD231ZgjRUZ1JxFpJ+Oi4iaQ6ZvqUaEHeiWK4Z4IU77OIe3DG
g8QfK1zJEYpPuejOEtAAFeRWY1tpyjQRyInX16/H5pUDA2DYrRgMAPnuD/lRbmgn
OBxZLjvkQPKbn6fcKWIZFu5lDfUdRrTxtgB75FCda66J1ix8uf9TWvqJNwm0ong6
Qk1JZUsWwEyxxe9uSsEXhJAzql+kxj/oSWt5+r/yY6fBA2bIcc+CONCxZPwi2ztM
/WNMkQg3QbQSGEMyk67lPrVzvovjNKbzLlDUKRpejY5OijQPhU225znuVHDluSsD
72OZLZEQt7n5foVRzcJtEwemDGvnnJdTTJRFMDDS3pEzMYgYpNIHMX/gMBheDe6+
+RaguLkL/8md7/4NqgjYEuVdaqLNa8dQPvz90DNfl0YRMUzKzo7a3Bg2Wx8Bs5DS
Nj8UrfHgFYWBGAdAxn6yC4zVU7CVfMsBoC5nVeUk9MUggRO9WitasD4lxezk/G6W
cLx8x21aV9JswOdgTYxxbLMlSFkgAXxMn9AxdJ5Ik+Pgj6KRC4pIzu4GMoYPhL+8
hCuUR9h8hInM+S8NsEBFD5jHONn6iNlUGoIBxNkHrvdKClfP69OvrZQPvbVDiZUZ
DJbdVuPj+CWXBXnaIbP4XnBjsskHJCYcSYCYplBqTI42zLsJK1VddavHGTKZorFB
b1Yvfws9Ghn6nJbTxTlwL01D8+rpzfKBjmYSa6tEdbsyZR7eLQaN0330yaEkqOhu
0h9xuJWTkv7+ifIJs2Qi/GzH44E5tcAyL79LGdZ7WYK2Y8PhfrqIbK6tKtI/ZWKc
9ptSvphkrFrleNycI+acf/+zX8EPt6JJNbGg3ZvTFEsb+lzHvFlIpAJ3X0AovTt1
/Vz5XYiv6kV0FevCUEvqLZbMOIU/bvY494DpZKsMvh7asD26D59Th6RD2YlBjw4h
QHl24IRZOIoP1vNTkUanISn0GGYt0ubZ8nn2MIbYbtYh9Irqndv8t2E8YPYjWBIR
cd6bwK8ILN41VG0huBq1eMO2Mk/o2NAb/DOYnJQ2cKkRuBoMLoCl3wW3IVhZAZgl
I3B6p4PZZs+cP97XZW/MaSYbTi0nqFvoAmKJAwziIzCQ8F3xXzG1ZH49PyefF4Wr
b2VBHlvqvbkHN8Umsr7IIS6e2NGELK0Tfaa9g5hBPXGWyqESmJJeVP3FvKPB/Z9/
lIEBDH+ZIOoWyJqkCpDT7mrUMuNg8fDgwyuxGXMVw/2SfMCGHzGI7Pxf8mIt7ElJ
W2vrD5iWf3nP961dYahrY97wvbh3gT0V2bKFNmA/r8sCcCAuCoVgaNgWKITYyyJA
EqeW1zCSXi93r6FLT0l11nXW4m90tKVFrMfuaEIdselI/WfPB7nv4zSqOnlfM32S
aW5TBIAQbiSXICXzXvJMQImvPLYxTvXIoDIRJ7uCQlO6zRrYx/+/DrcIzfBgFgTl
2gI5zD+40FTvgwLgO5tZrTk0J2IOqZPeyf9ktzCoezVSdqT8Oke1CaNOUhhNxOaj
1JeYWm6AKHO83yGx4bPkBTcy9RU0HpPKeCD6EmaRlKIt/+/zK3VciZKtARGvsj1t
Gb+909FmIfKdGdtpAuC6xilOcvf2/8CfQiUx84WLAAg7AJEfozXlyhYNGePCbq2o
NyWzlWmWfXAQAMyhi9GG6hRoQASzBuopqCZzTZiLe48G4jc4ZBrzmiZT4DclNTGx
en4/+4qOMaaLWw9bQT7ZnddAd4HigVGUvc3XbAh+LtUy+WDYThU7G7fquz8QCPE1
VvysSc6hvfNZD9OcDff6tUaGIX948gzVYCkxkz45ego3auaU2jGAJEQYDK6cjAly
ooUiMT+ppe9Z5ESPwIzjCZwT8Ag/DECzP1+PckzuAT6nUePaLF2fRd6BctCaq81u
pqAMAK7IQiNHCb4BVsUeePpdQSyg2xUMmGFvvPyvhx2DqxBsjzaiheD88kZjHmJM
jT6TQG54PgvbYQ+K7r6F0eAg+OuOlkxnteTbnma0BPeRI4MfI0GtSIZjoAEU1OSj
bDsLfobxP7NWtEIVm9exFeX1fvLlZiNpMhcJJ5j+rG968TpResUynsX7oKXn6Anq
OMutuqXVZTBLgHmwIAnDvw0rEN/MTdy5fbRhXt27qsG/iLrmXvNu7aqJo7RrHtug
e9gTmGHp5xCkpRZJ6oRnw+x2w9Ndg2BgbJLDWX+JDY1/GAyktwikLLudx7MYXE1E
2HtUEpVLnoZo0UjlLosyRLfnwzrrdr5FsFGj5nKHR9/floWTnWiKdSYxBfyw4rEQ
v5L7GkIpwkxzS5rjI1LeQ54Dhecgc0wNy7YdKZw9EsLam7eJC593QwAiezQ0Cugw
WvGEIB0EgfFOB9Wwjq2rBNVSa8/jtR6NOdvVhsM3G5lFV3MokfX1GpVeAtC3fKaF
J9V9Cu4h/IMg30kw5w8sTa/nEVsMsCmGU2U6f8xkEGbFdvM+BjBMVPLtZwDPOqIs
R4XEctFH1eg1wS85fEafCEhclqUnDedXtXKWyiV1KAWGixqh0b9+cChiJt93n2pR
IkdbsqnYgXq4e1RSfWfFgWzfmfQ+mlDnBeeGtr8tFS+w3pIgipmz1w6kyAUa8a08
97tZh+oFsl8II40FxvXOJrpRczsKdkP/pQgWvV4QNl+Y4zffWZHCdWLSFCJrUwu/
oAtdZBXSI6ewBS/1hqR8exrvWhEjn0K7AgyTWYXNaK1hZ7RUuxxkP1w8tIfUNxsK
s6LGJH2LQCJdxletLmfyZZSpj7FQrIi2pJmdfCytXtpzYU+DJWmd3HGXt+PIlvwk
TBoigV3f2Covq1qnBt98fp9/nbhyAuJBT3idbjfcOzYUSDUGd5rnw4ZPKm+f1xBC
dLBGzbpKR7BoEevv4hZXmq3ZLL9Gbz3e4yWOCbN4581B/1Id4covDMel87IVs2ef
K59KvYH2mYBmwT/lEDFcXvx9ZDDpk/mWYgIVKDrUTeCfKjZxxtNsCjpOg61EvIa9
jggizIpKGr/dZVNQ5dSvSscewX+LmxDhCWj/QcBahCIRosZESli6MivdVXBH3AoD
H15/XTtPJdNwLubPdszRi71kviXApUMXEqoA9tMZECXUqT8G55xNBJScapeqZ5T+
73uj3Pcp/G65zSUJkcwJFJjZg2Iu65gAdXuqf1IiDUDkmHP28kr4eFWc5cYmT/aq
TcUDk+5pv7ki/175Bwn99I+sWRyBm7A+BpPGG8bX5WVJn9kyHzEnOvJalk5hDiUs
eLFzwlSHXbIcg4tT2tX9rRa/joeIZWAd8GdtddG+IPy+jjYzocVGSDU02l4h2i27
RUGKt9IJgxW60CCwTomjc5CnOrlEtBKyV+ivcftI4Znlfp+utjIRBlRBNrNvgwdC
apQPmU1LKQ9HBMm7g5QXG+IMHkU+nXJPo8oOIDT4ukjNucLPY+/LrW2EkryVVyBl
B8nxYuMGKi8TKR5sS2QiedusZB/f71fVQFyKTi5rEobH3ilOQ6OUI02EXjvlSZmI
2e7jXahvu0MFNUOdVaUKu0ic9QBiPgZXrowGmDLopmo5URE0k38Qndzn3s27uGHG
uRZZgBErx/v6OmBHFmhiL6/O2tih73sPziJ0nkUXbwNicczO6J4yPuG9OYU5bu0i
m4SHOn4cpSl6cjqXqbOxP+7Td9RHpcOyg3IscdhAnirDQoNxR5xghZP1BfbaTdvT
X1XgNO8gjTLyNaa3omJ+Zbd+ZmK+9dbn9fmAq8I8yQNbm4E6i6YYAQsPw9iGDxNh
2wck1VO61sQLx6OMJJZfVEfsjP3VQG9wFYeyygt+bEzadPsgGA/9xWoV2cvVtiSM
Kj7GYhWPiazMPLhccr0ng44sLHPyw3KezsNtX16Jm6dZRRurWBis3+fI9e1XbaTQ
h++DatdKB+5beJBhgTMKgc/IAvfynB3JePImHv0soKjOLdndjywrDNfFhgAaQgt1
Ux+k9mcF0DPFoPw12JdzFLCgHK5kugFMEv+jbOLVQxTm/WVwZ+dlGPLu1VzQWTDs
o72XPn98uMVOBx68h7u4i41av+jwCrVpIO73Yis5d2yWNIQ/k5LUkKuhxyXM1FyU
f2kq2hd1JQTD0nZCD0Av1zTMnj73tfa3B7lx/DGCMGG4BDKQsS2uq4gtbYuCd5R8
n/JD1/oK3yz99CRKaZ8OxxsgC2GV8ifADwToXpGLHGBO7OftPFFa+2rHHsBzvCY7
x1Cm/6O+1+lDtjrbXu40Ho7CJc7lIwfR4UC2W5z8OPRTD2IJmlX98CZo6eBqFwHa
VjP8j7aImYP4FgmzZqMURyTla9jaIhnmvDy0TiSJ3i/1jX0vK7/umxromZtjDweD
WpNZ+XvbQ+iQ/r2JFbMl3fhmiirKrfr1W4+EmfsXbH8udXk7MCRZe3O7VcPNd0kr
y85fWVRAE5XLcXgoIOwHoSHYv/gm9sviHPVBmBAvJ0omXXrq1E5MD0/58/Ul3Lyp
y0N+ZMdY6zsIJq2snroQl4YWwQgnqUCOKlUuTgUd+Xcc88fnaC3PL48Ydi2dlq5u
JCZiekN+6u+WxwBdr9TRtW0WGMFPA0NVITkMhBZaAE4djGzh8t4k1GShnMJNR1pT
wwbyKG8EoiI0ptO2qJOMzewwDhCNTMglhjUj/7riHwe24m2idHgc4M2BfTapanIx
/3UtaRmYXHiLp0Il9vR3W+6kz18NMNQEc6RKr4a4IGEL3niGqv1/k8LpvAdphVnc
vHn78Q4NKDu46IweUulY/TyyBvnsaX+MBm2zPtoH7nxFHCtQf48sShJNyuMHrhfk
H/tdbC1QNUXaCRG3Nhjk9nmPGnuDbS3vISds9ZLcSaTQYHFy7mDHTkvnUMMNYDDz
vdm9bdf+RhV/Eu/y7QL4TlGBPh3vKBaWekYvqOrgHYv6n8j9WOPxLMXa0yUGSMvi
X04pjUEOIYy0TqEsEwb1Qf0I6tzrr6do25OcFp9XqjJolCmTK6cKt6CV15eddc0V
jwXHgTsBNd+PBe0n4gxh/IJbJkaIydZKBgOzH46uA6UHuNIGPEymQIkWsuOTOc9l
KOhL+wLr7QFKioQewKm4fMrXGh9uZwKUHafnatap9JkbkhJTMJHv308FOOX+29Ls
USm4sdlHgZEWviCWGrh0h4FHGgHLKlMWOusIWYHuTJKxUdUXNcfuexfTMZxIZF/v
tNPbG1k0F8Y9bWt2e6fJCkS5DpOftUFo15JwLxVC2Dld4TpueDyED3O4Cm49JXIv
m036BIOu9AQ8/r65+j03D+q3VGZ/pCLrNJBORsoH/h+fm6re1skBxhqSnEotdNbs
3b5q6UelD4HTZZ8y8qZECQ9ebDTiisFQoybk5g4sNQXNtUDHY9YrEJDSgqygV5ol
wmaGd7kz8Lm3jTABWJdFPaFO3ZI8DiAZguFsy08pRlJ//3pqMhib9YBmkgUw0Szs
w8Hyl9EPIBUy4+caR5ZM1OeKaEJ2v7LN9k+4zAOeh4UtLyxIwnFiKttlqfBaNeX5
C1mXakrDP+XPbPNjdnvOe6iurb0hWCBld2PCfmh+JBAd3akscTTkXh5vmBJ87evI
3R3P0pNyXf/XzjWrbSiktYub25kTYJxOZ9kXBq9/tr+5lIKMMOKe2ekNZHhSfrCE
Eab3hVsQ08kn2L0NMQBWkAsrMeuhgkhEMy85h5hlNAdSc7E38UA2Cjy9fpZBMJQb
/bDuahRzmG8RqRrQh6tM3jcTiaLvKSfBig79faiT7y8VU2R4AvdH2/g1KTUuxQ9L
uV7GBXaDGIXN4srp2vMQwT5qU3UL+nE/+QbkZQ3t4Ww=
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
QC1xdnWdmBBa3ogfYJYMPyHyv30uQwz+hae2WPtob8Zp3H+cB0cwoXM8tNr4UZfV
LsPhBMfw//3yhN5V/PiGV5V0p2aU66EO/35NEsz95Jri8ifwoohSOavKaHC3yJqN
CQhGHaUkMCWmZLKgTpnWiM01RDJxsJiasIgZaGhFYLQ/G7obBEv11BnpeXZj20RG
Sk6iMAzSmjI6TAfDJI9gSRvKaJpn0qlRPHYh89bP2PFn2BPoDp4QUUVb1ePBTyVv
ofIoPmn+jZMZrkTNmXg4r4phxKivJKza+NCj8urUls2mrkpheEOzYIsoeqCbFWgI
jUBMLKyLD63xNIm35RHQrg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5040 )
`pragma protect data_block
tLkD8m5kV5iv9EYc7Ywk3tnTiPmNxm4Wby2mTDvj9wnyGaBl+gKeNqXTCHGVdw63
vABwNs13AKLscYSVpa1Q3h61fM8kX+YfSGtC4OyBd7vZj029OgNjqVQjCQnTx+Hg
aukpUljzXWR6ibQctNIAHJjW50WnGW0n/yCwhldWEEN6uXU8+dGoyhffOmfD1hjA
Pyr0yl1HmbIEDGaseQd0tOkMQlbJIeDCGH/OX0CLbVWx2ESKarmmPCZIz3YJQilu
CI0bl7oIGns50FNBFKhhn0YQ1dJpbEloZt7LliMM2N8WuG6t5bHk4fJI3qRdXX1/
ySZ8yhOwNSvQDMV2weELIsNyVrq1DrkSpdVuUUh7j3WDxeCd2SBuBkxv6K7aNM8I
5IeEv0QeeWG8w77R2VYHNu642GZ3vLH3wTCLktkxRxeICkoP5q2DXKEojBg3s0if
AKaeiSxOhGRWaop2Rmwu7cngrjQS7mVchKa6eN3TrOCPiTv/ehQHHbFc+Ug6jkae
v9EP0RNQ6LXu9JqmgTwScLNsdnV7HpeZU/vPOP18ZbYPN3hikLO4SIQCDNFEcQyD
RmYB+exHvk4JYjN1bhtr9a5iWujwXSXOSgkw9bp2fzBnf/42UFiru4ow2OMGc2U2
46f0h4PC6R55BwviJhGlgZzF66S3HtVq+ygSwQZ/HfEmrOLiYXxGEC/XMwGY68GB
LjZZ76HYja+4LrgOEgJFtrjU3dKejWVN6n/2GmwpYpNRBFMp8Q+hnJaYfPo8NoIq
Sx/2558kaew8eS/lhtPcKE/bspUQ+e3dCydf1Q6byQM7p50/MPRbEzN3qpT2RRT0
HzidCgtF0AdsF/ZJRVRmhsq/2eM/2XRpP+Ulsyu3kDDBloOp6ud5WzOk39PLkZPf
BnlUZh8zRyU0WlAzbxkuK4QJ/c3oDXQnW2SRj3ASYzcrrryUUoXAupFifzOCrTPw
C0pEms6Ao3avazm0YFI9gaTDWV1F58UFrb5xb4vyuTdFQTpXk4kGVqja8qgFo937
4zkoGsIo5YRgocPCI4L/XKgbbbNfbcbZ01q3SWXnGVSMyfChvnEQdCrAMR9SQxcC
nFxSpDqRnq160HfC7XNPVHjTWgyDvjVOT0YV25blJ+IHG1dJ1mwg7IPB8NK3UrJW
DfMcdlyfJss0Wf3GIlI8uRtnIfCi3/RKTpvSp/YtbdFZMnkxBy/fxnQ601G4g9xh
+/0Mp77hjK5wFDoNTez7fuKeJpznnZnIFAnGL4k0VmIr0HP4I/4eoYrH7iidMXfJ
+5q+aVlWSEdjXoUaAYj+XUZqljoNesYGtjXIw3wBdto2igHDQK3dGt8ksY9IZuw/
D9XlJjJyrVojd6ZCDUdFGIUSHssNmXkCbOyWAoNeDoMygmu2PIgtzixhEoAT3WFf
JBu5wmTGe0r3Zp4Dv360G8y0oKbyMy97GlEY7EeMLpOSMa2OolGh9EejzYAxIWTm
JasS5XXbVvs3QFVN+ufl/2lc0yWUETE/gL0jQFOo8iaxcSjruoQLRM/dN78u+dTX
r36bLtQoSW3Ps33rGf+nINXrfa2AsgO87BLH83lawlghzanLW719RWZVMCIr84sM
ZMVw9lRmqRnHSTqqiQ76/lvrF/N0lDcfSMgyUo0sSQxjtp16+i/IVgze44pKBDvY
Naqy0y0uSNUHdLYksk2knCtAb4SmUbQ5RCuOfV4lSIPG813A9XmLCDE3UxoTaeF1
TQm3SRwWzAu47XFnVrERq4Je2igIawxseJcG5JFdOeW1S27WIMuSIBz26DyNcY7x
JVf1eIYREggektU5rmV5u+10U8GXzN6wST9kNKEo9mt5bJKF/lEMONqPwf98PCCn
O7EvtZXuMm4y2QNtytSWpEvSxrbnJ3E1S1Tg/zfz13PWiphN6DtRp7PUZ3h+8Oc/
nAybhYw5xT2IplAqugylpbeh2leYqYvsvpiTk/gY81zMMtaoGzBacFrg20KetgIu
Mbj4e6u8ZJ9H1trWAcZYrHJEn6MvWX+7hQFUahIgu6DOzDG4RhY6pFV4iIkljc8Y
p35/USdwlhW6WNx87a+NpwmUMLYbpNxrJoOpSkHFEdNvktGuLya6SF6A7fKUXNE6
EyOlNuYJ832LUAwPiV463I1iFzN5DYngCveVwrhKjB5PUF916xQO3BThnbdy4fXR
fY96d9rOrsMZJRKqnDqzFNluIkCFOnIIX8SQ4QoSs56bsdHe9Lx0A1DoyiihLUPO
ID0Y4DWsAclJOjBHo0s5BE0rf4YY3g9t72OwzjxUHqcwhzDtpzi1VKqQX16xcUCZ
MZ3rcX4SAjIHbVRI6geUnJBu9FanSrUnShRvYyrjYMiBpXcN3NWYF9Zr9Ad76WcB
IQgmLVW2aAHzM2W1ybFpFkK2gLIi+ch+1BfJI1MCuy3vQDKkgql5fCUy53NvrBKu
CYr7n6MWkAt1wId/xt1KA7nPGfCsi7wveK+TK+UKu7yg9o52tQWL22uBcPdIz4uu
GtMsSfEEcpEFaOGVXH7JJNdJa81yA6MOjGp/9Gd4vr87Hzvw5gHO/qRQlqXW1gfw
KfiN5Eb6dqL/wL0khcE2fxu7xfG2DXPys1Y00bJ/rhKQZIIws7S1KPp7CWpIT46N
m4xOf+y38np2r4WFb3obghX4ZR44toYLZs9b2+SGv3nvElMSE5tr+/xz/x86dw4T
66YYlwVAx0FrmsBZff86TxJce015QpaEPoh1uAgUklb+Fmhb+MWUOBIDxsZTnZz4
RD8JELT9G0Kvui3PYOI+CH/7pEn6NESQJrJdHOY+MQTaBpV8MYMtBHMOXqwki0y4
kkIDyhDC9NgXknnFKB0pKlYeRTO2TAeHwcK2Q2mUUQoimZvMSXDjH+JRDUTYjetz
y3ZdD/n1Etk/EpjcRDOCxBuk8Hr+BJ0cqRloNQuiMXpRHlQLIPa4KYo3NlGMXTEl
WwHRJS4gKMbXOQneEWyoY5FhCjYg+ltSOniVmvqCItTOSr3xjafCT0/84wPGTEWa
PZNClcSRNufpwHt67/mGXQVizOD5HdK5b0gE8HOxp1nOXYrOYd4Dk0goU4yprK/M
rZg7Bi+dzfY+bMbWjDp3YSzw09us0Bjv8k7KfQwA45gEMPcJv2SqZ0WuPD9nLL82
Ppht8tfz4qGYdVqhEJ4vkmARdZi9D4tinAJTH7R0RRP6VcrjqS1BYH/deFgZHJcs
tuMg+vhoE65DeKiBuUr8AEXUXFXqvo509hPlR8xwl3F4KLzyRVqGb6+5QkHrTGK7
I4NgvFgH3CKXchylnYZFXOSIDivbu4sV7cv3hPs0HTeP9iDicn2RCRPyMt50XcOS
7TCxgdSslnoYCVoxX2nUpf7NVC4sDkiRFfFpTPCwDJ67ezWPAvIpD0bFhmS/6mxH
QFlI5EBGLJXGUvZBGAwvL66qfGmLNH9edWGAXxXFcDawpIHbY8rH5L9QbQVCD8bm
NwbMg60jEgp7gGyrX4/1tUlYqnnZqUI0ylBLAAcKRdTvG+vojTz/DvkjK9PEe/9b
9SymAGF07ItotRwwsrDR9fi7xyQK7Vpx63qbWczvYxvC2e8Ob5N+vPdAMtF4Qail
V2AX1oT+CvVGUG/aZ5TqtBc/4AHe6/3Za6bTM49uiQlstPkqr6r+VfWF6G0D+V5y
YfSluduD08S9ikdI1MqCZwFhCNAXg0/3fVfdQZ033RNY2hlFaZoCRk6NQH1fJl78
Ql4KdWZl+IHQodrX1j8tiXdy8Nkk4xPNdnTn8/j75QiH5sZ8STsKzzd5vkM7PoOa
VAFY/YY5GjlwhURb7ux3W0q273OHefToNDH8TENFK2VtO4YouV3CHlfUGwd71ame
dfk/R/lW/qfLPKA0hz8H/ZlUJdMSO9i7CWpH1ALKOiG2da8AcF3yWu0glulkIHcr
t0GxTstjWl4vIeiOYWEJ7CBgpy/b0AiuB2QUHS8RjDtqAqfLlyJsGFcc0ORdlbmC
S7GaBZrbrCx2yNwiDXHyP95tWlYKE8pkOAMAI7nB7opwwzh/ZLOnxDDnRe5HriCm
6HTk3fl6Zatz5gpv8fZS3+keksOxLZCUm9qptInZX2QOIsKVcMcqpmyRKvY8cCib
adKTm3DDcsUZH2oW/pkqrGFdCXO5cJWHvidyuycR/eZa4uuEDFu/McOqOteXwX36
ZCVtPtKMTsMytskrG0v1XNtqj8c53EKBKgbQiiZT1dthJfO001G06+JpmMpm4RUK
7DiJyQx4FIdAl435Ci4TyUg+V0hCmgH11XUf7tl/FGI9TeGf4pkPH8TEsv81/w6Z
oGDsfScd9Zmq+OGGT2FUCRWqfWvPfDUlLovzRmckHoUHyNLkjJa38TM/yL7U9PBF
EVD62SJA1NVrx5oazYmA1oE5nghyxREfBVomUKdUA1eG+fao6ca+AKBKHaq/8yh/
X65A7GuQojfmmInf14LfMaQcIy4DRogkgJAmbvr1ZgPU/AnunbIq+IZKk4J/7aAn
gUSgbXB4cTZOLUkptzw+FH4XO3OBQLI/Ctt+qn7UyeCp9ZKexXaPy1wBuC415wRB
QXuRkEVIT0sGiqbmPXJLfxWwmGt522oM3JWP5f2c5gSNedsBX6LMzwGNxv1sanzX
cjrFMe5XHcccBQP1jAC5KWbC0mzFH7XBzLGaT/CjrxcPmMZKllxK+FneiYR5W12U
7jM/9MEXJyiZusBWcOOWgglyOOxQlv8NuPYRsCdT8FnMaFLudcLx7TR33679RZ1x
R80w9dsntA9AyQQK5VWpqnmfwy9EWrjP0dgrZ7BgmRqKDqTqwupDQ54Mcst3adsc
OEVFkzd9y/7SlVU667KuXGMv10VtBe2d7bNWinyjIBq41wLlARKQvuCFK/b6EfK/
EKae+PZinDhD1bo2DQAoc3KqUtIXn82zqePWgNiIKYNy9Pc0CnzTe6CVcyZI0mxO
GgBaTpIxG8r8BU5m7yO+f4DzqsANoM99/wU81tNtYmg4CV51XDzD+B1dXplM8wy1
AfClNFyyyPH6FCnwgvV6aXttri8smQckAW9mb4Ka6NI9LlWEMf6ucVURFjDf5r/C
19ed8PtLTFmieAS/ywcwH7GESBxELIwgcAM1nRSLjQZ3c8X055zWGahJL3MErWor
t3aPDwFeTqzKvAte7KskzZ8hoS/KXOCgG0J27DoVb0hGXjUEDlpowX+g51afZNRQ
55Y7KTZhzgOcZjA59hlWWnyYRynEbUPSUfc/Q20thFwUGLR8h7RRjDMP9pQGnol9
2jBiGWA/mRkPngCHOijl4dKyUyg/VidSFO41tUpUskc5qwWFe3LtC03Dzlv2WxLp
3KmiiQT9295LFt5mQF1dobLIjaohfDEkIVi0vq6qPUdv8yJ2ZWPnotJlU1dnzhxF
fKKmN8vtU+OD2HF5D80d3k3/j0695a2U7JZhtrKRwvScagNKETiOID5HYBH505Gv
odnFbKTkUtTcEJtg1ICw8Aw1CpvGchC94itbAfQZxjilc8MEYa62u1WOW2kLc7P7
Nlp5OmLoZMLD88jIBqtfTaqWKTuMXqqdMJeGr8noAWdF2VCYCW5M628muBijkOZO
p3KkmP8zj/JMuy0VZyKMJiV1JoFrTmRER6pbrFyYnqPbe/I/+5OJAvkqBcaRgV/5
Dtzd+4cf4bFUGRnTUI0UL9n6AaGFM3UfldOUmonzZU6PqE6YeRf26syo0XMkcgFN
Nbhd/dNjFCovQmOoplqVi6VA29YPIamD0mu/DQk8RUwpDM4a+JlshCUaX1T2/6IE
TNixOZHhoqWeNNFFovFVRsSLfqyJuB2bq5U7DmMvOP/j5e7PR04A0P4Kt/9Gum7/
bgGR6T6nYKkE8s38945NB0Ez4ssJDhxNn+KTk9idc1cLKiJT2PDt6KzxBf80bILy
2+PtjdRTyCSqHX73MT7qzMQLcoohaMRyQx0Vj7d7vY0P893N03zwSuRnziAwOMqJ
nPUZByX8PHIYF12cL9S1Ia8gGRG8pA2IXt0ExmUqXeOlZTOSLdfGNUoMEhjS6c50
VmtQH4csrotWUM28e1xxccHa57pbq2CYXz8gXmzE8A8rEeprnx2MvkVgUACoIRbn
BwMhWSeA7LC+ucPVwHWCLvIYCUDaN4r5hfwisPk2GOvwtmOf3QyCXJaWqPd0jB9e
B4drLNMn5frj77FxgaoZR5RLzpWjn11R0iQSqJHnkHpCfZala1Euxbh0hOGa5nDA
cWhwQPnaFoKlOzO8xMNy1LAHfu4T27rhLAzWB9pYnal1GE5FZfORvDAPP5ead/N7
33YXl4QDHOqYcW7k0kn6ejntxuy1mefoCjE5L/5FPBsmdCMOMEaQRX6xLxUXfD9K
iXr6lFMuQ91KjMSThbRmb+mHCdJ9ocCEOolKL94H8Y0LLRn9dqiCh9iNHM+aUDUU
bx/rxkR0MiXuAhsniNbeE4noLi+62z9tZHGccX+ncl2uySeIY3z3+5yWN0PLZ6Za
QGVoNgh1WF+COrz9YkDc+I4Y6HHAvL0+wcaoSIlDDkV+aYcF57tpI8XQr1/g8TVR
BhEaxjzpeDPljS58DDf2e+/bD7dHekRxm5PjmvfpJfaLQnzEAJyqbcsNowKOwXTj
IoUi3lbbjYv5qgziDeaJMpQzD05/j5M9VK4456FHEof555Bcke7SljCs8XFMGDu9
123/rXL7szAcluc/wF4/pSaGdPAxTLBFE+DCQBpaimBzk2osj5yAk9L5AV4qpwHa
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bLE4oUWSuJO29voDQW4AW9d7VCc7ne2Qa1En9e2V9LZvJYLHsBp1qt4PkEC+Gblq
lSpu/Lz44G9VZ4L6RYfmmtUH+HNHBBZ8cXQVO/iOAE0ZJRuSJVB0mlaeelGjFmSy
77FYHbehnVuq+jHQUJXHX7jbfuQIJZsrMUjEIkEhsDqtawQPCKYl7C3mN9CdmUNy
II4fpMl4hGKesov39Ym9BaqCvZ4eZ2AmDp0lM91+MBwq6CRNnLXICJlhx+hjxrl8
PYucgfWwukhw9jrfjwvams/Yv0JK3E3vF+Urkr34Daeg0OZ5ymCzamDqiqbVz1fA
6ixnuqbs+QGCOiVUP6r35g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1072 )
`pragma protect data_block
N8bdsN+B/8RywlzTJQa7+KvvDP4Md6FGymmKJve51vW8yX9dGWtdRecImSyiK+mr
rVtH9V1ccm6ReJQunXItwnSNDp6kmaAYAhPSBtmxas9e8iHA6S/3ly2GxjzSDLNu
ZqVMxb1L+R09UJoh0TasvkQPL4KJsuUfJPXR1FAEpT+3Z1x8l0aojXsnHINhisbY
pv6B7jQhDdHu9TtEgVfVi5shwiiPJo2UT9KLaBXNNj/t+Th+l+mMPYzx8QLsT0Bp
dQzIZdu+5fap4E5vQz1WI/TRlhu/HOXyBwOPWJh4nvsGZn1jW9Kcb/32Etm2tZLt
bOD7MUcANNMcwHF9SWvs4mw4TThluL5du5y6n7R244OPfJ5s28aR529y5kXaym2r
JCxmH4Fo8saTyntfgStEwiTDpYfS3B9QOpBbbkr0K03NbNGaMbTFniKudg7R+Uvb
4fmJd1ucNyOdGQrissscS9hoR06SP4YsUgRuxBx7kIzd9asOXc0UWdCqqMCFyZhs
EAhxI9lk7giEavQFK5YQMqb4AChHklQwBrQb4PfmohVRuhvtsQFGe0cpQ49s7hiF
grQrbQB84TUvoORQXfxZhVAIl1/EFhoQhcbQ87YRhqLbLr7/kHGiCW/UEsGlia0H
yYbgSPYAqs6UjY1f1VoAh+krVBrrZJRw4d+CpW6JrwC/CZyjcy0+eBRgUoyDJ03W
X8hgLHLbNwEvP+ctab3JdsqGEdKFGVyMImC9pFoRzg+pob3mlU+bxjRP+XLCO2sB
4sf/UxPLOoFaFGu26bBxpsCwMj9K4WeCziOUENBYsD0MrmzLORnV7ZnvXNSRa47e
dmoBDkqMqRaLcWbZExMBZXZUaGgxs8EeP/gcmyIgVd9iFRNWwLuZGSLi9mgyP2+8
EMi7uxDpUkE1dGanW2hYVgzVHqdeZnrT4GFAb/1hRsEStuuwgeKw6s7KUwAqOW18
3eZMcaGh3oLXBc9lYTBndCSNc+SLDxgZ5V1dtjmlwogOSQXWyrkw4iZUKTObEnCa
EjRfK4A0ad/1481OAz40xTY4g/nEUJKqIdVL77g8xOJ15aplMbNBy7kPmmQPaqbL
FupRc4SN5MagtAwiCa+PcDlTCSh63vM+4SaoO+o5Yjucbu8VYqPZwkRqERpaMRcB
5OeDny41Fq7DpvkmZKEHfI41QmNKRwCslE+MKn2tfF205coo/he9jMO/Ks8XsRAv
9OV7ai/l9mV+guqsh/da2KzIkEh0o2aMcx8kY8IzBkiBp2iFrFm6bqGopN77zu4J
W11x6bOSzy/mHP7lu81L0k23aJJVjzsYDpylEUQIiiMUD1QY2g9BdCJyHSsmha+l
CfCcDJ0uzubgsemXPO3AaNN0MONe36pD2teQhWNVqFKZLgdlPFJ+T2jGrXoIZTEW
QR5CunkH16HCWI7w+rgtCw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VCsbo2Kajss8mlA40Z394xG33mVQyZLZkoxjMyDIElAAJH5CJ+n9EedPYZ2PIB4Z
jFdnuKnBTv8C+fy7OV8BHeMVGxrtlUfi+fBTCXUaMoCzs1jZgPzZNObRMq3HgFMR
cOFFro5kan0w1wK7YMSuZFmU2dnoNhAP6rKbMjUyVZv1m/6KN3Csxaa/mN21zn43
kJV7vaurRiL1aEE2DLQ25K7Td9VTnZiKmwtAtDh+9UmJ87pA6uRzmAQ2JFzWdCN9
UV1+bJZoKhSCO7nEC+TKU4jLil11xcY4UmP2hpGy5pNaHqd5n0QtEWzqwhKanQLB
OyNEHu2rTd5ni8RWgZfEtw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 784 )
`pragma protect data_block
KbgpckERqn6qwqaMY5ULKxjnGm1gzSoCtbMW3un6oHtWvLj2QUPT8OJK9HgYKhYq
RyHPOyWZ6ypYul4lKvCYMkPpDwK2qqFdt4M0agnBQzfSEETGCXUQNRSaBWbogRz+
f8EkEkCL0KqNLMfC0jYp41mLoc5pM5rxSQAV3xIs/TthDgJCt6sawSo2KiTZPb+z
lVV4DDS8+5bZ/IXHgzDK+j/29E2BQy+v9rQEBVE1ke8Pyw4a38NXEo3EGRTLNXmf
JzxysBl0rMc+aRIRw4SU6RGyEAYUbf+DwcuO1Z/K9Q3ZEw14T4ngWB0H5b5aURjD
dpEM1WPeMpkPIxMRJGanWzSwevrxeGY/KjHjODt7PVlhDImZujuxnqXS6JY0DIVl
f8NwbHndv+sMrUwWcJJ7OjoPvt8gJrYNQU9zWN2JMNpuPSRw9EwTKO9srk7cEY7b
wGtIt/cnEp4qqPmsYT9F6mJx9YEcWTFVGsMEQ0kj9S1pLvMc+17Tg1VvtmksQ4vF
u8opwr/j2QfFn68dVM0dZv65dRcaAjNJlDSDxp3nCn6F6lNFx+6KU+GzWdB6zBBc
1OAdI1rk6KwfE0MggNCnPAMy1ssCMqnHnB3ifK+s4k9PmECPGOBP85vkiFOrSSg8
PgzoxN1988lBddDJ054q0kPkS6DL3gTqskWSf3ikC1hoOGOZ4BJy2rG/Q7t+QMMB
rHDxRF2r/EyjVVXL5wBLFMPmiQEhAU7yshKdFVzDMwJ3fkFQXypu+sHhLjbIKQeo
G2SRH/iv6zfwnj3cwNR2+65quBax7lD46b2TKdqYpCNm0xf8QI0OUwbQ0ekjgTph
H1LKmcQH1Dtm8tCyVOr/9jFHS/V29152QjCVUWzYu+E9yhAQ/g0SAvWjoUFUnoAD
EEVjQOM7Nd0zvxsQOEpTV95jBDDth/uu/dtKltLxtD0Qot4v9WCg3dAegRz1oV9m
rQlJBqcGFqtVrLKAkX/mpb0Jrv196/bjJXWmhBvz9xK0fIP8DMv6aPcgI44BFygB
It1sri4YfQuJ+lbdSBn8jA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
V7uqkfXZhZxXk2DkqEZrIaVNquSh01HsGijvHqnwhaej4uZPYJLCUUz1zS7/Z2Qw
DYWLS2KNrFuQ5HqlIyGaRH1VxNHr3r4Bw05HOUYivoW8e6FcHnWWQR6VBuoqT7uX
3DXo/EhQ/WQPfh66eC2VGGKFZIfxEJ/ug7Nc3VQ3Ei7z1PeNVQdm1xRcm+jZ9YgK
uglSTLHx+1pOBUXlavyha6ei7qm2m2RUsJs+dmZOjyR9zls4+QSj8pRxEqex1L+G
vT4126RU1DSu405lP7wqG9RQG8R/cpx7UpfPCP7AuuP01xyyFdxzO2Cp5n+j2q3P
sDV954b2AxA9W6IANFKm/g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
Q6aI0tjmBw5qFEiba2HUU8fDCE5uacXmmII5FP9IAa+JdLcVPspoiINoxppbudhW
xEfrwTIcEqthN8WFq69f0Cy9GLv9FrJPtxcDwJ74kyv2ik25Mzlp6kkBp309g6qH
0D0mhhIrKKzWrAXoviKpxKBmXbCn+l8kSYHPzWI+h6GpvJ+cG8uzUcHJ7WJKSqkx
rmdTamKX6vyJnhbH24me2YkUnEHEGuoXUc3rYXmyyyf7ruJPT4cML93PMJLC4Q63
hGIzj4a3yZ8ecivocsQm0Q4st3Kra+DNl2HNu/QyxU4lCUteSNfIfCvxkxGH+7yW
mrdTdfZ43syJcvy/qSJS+DDz3ntKivnZ0QNY3KAA5p4DvD8znKi11SQ6J6+UIkcr
SUB1136PTWxqb1ixSvGcOCu9EnnxiFk4jCUnahlMFfe/V/YT08gcBFUeahJfkWsn
kSZytVFuGr+PqsZDddq7e3sjSdua2rE+i9Z4965kCO6PS9FFUzRjoaITJM6VwCJd
ZfFiHA6M5iQEE4Yeuq5wnFFSjdCZ6ZLN8U4/iPrZ54DF08taA554IaXR8K1R6yAb
tm8fwSAVF5OOrGb0zuXifggNORMJ3KiRNB5W1jpafXsnMiIYJtLTVz2i4PVM1tf1
iveKLhpgPY7lvW58VOVaxq8fHLrk5X1a8EFyxBk/PxuQmTH4Qkw25E36ADKxF7j6
fQSBsIF8vCYGWBetVHUKF5SJCiit9YY/kokdmY+iHOsXYlgo8e07cLcn2NViCds6
+SU0AXNDjVGZ4uzMjEElP7B+RxFad4G89WZ7m5dvg80AfYBXR4cYCrOOHWRrwEZ9
4B/Fd80D8Xb1k42YtDDPjfgsFS+3fh3kanpVWiTOQBOuSyPAKrHzHjA/1Nh4q3AH
Ghpvxz3xBQ8cx2msaR+oTRGMH+w6zEb7MdrCiVGM4Bc=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Bit5m9YVBQr16yXC78xWPHY48nwzc6A2Bt0JvgPsl+s5Vq+OvCmFALzhfB/TPTUn
/ltZ8LWQdReIqR3IFR3Anmghaq5OwMnWBf7gln/U7ZXLsrNGv2JW0HsjfAwrWd5R
1Hgqfb1NoAQPcohK/HDko701+4QJ6yqeevxMod1VQojluO4iqbuD6tGAul/U2KtZ
UxVgQVoDxLRhCW4gjecwqYLN/JJIQUWt8ARj7lF3yTOQikLNIS4E+0s6lgKIGbBl
uUOZYrG6MLcNyPOLE8IbMuYmLdcgmDQqbt0kDYNOKbC/PXpxfwIbFwJFhqCR0Vbh
uBQcWt3IRLEMpDvmsh2WKw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1792 )
`pragma protect data_block
baU6fkibK3UIAtK6xnbPqNAuwOXOWuZCxb57zGk5qaDdWRoSUebcVi9O0b1C/jgO
WLxh7pU5s3To4EMCvXXJx+MsoG0f7YA8YNfWRqlGerSC9ivHWuO1e/G2i4scjlgd
v2UW3GggQIuYa/E6g2DcqE+ZUEwKL3Vs7AE5/0skkC4czzcOs2N7cMR0eTv/pvT/
gAPptHY5EhM6/an6ja3uCuRjCLD78O4Io00K+OIK+zn7ZkHYH7k3qb33OVm+7jHB
Shr7+KT0oVfrVR492TtoN3emwb247B/oDgaRmJZ1UC9aq46Zz09IdNlhW4Yk0Ruy
F/VuaOcR7UEbU3BZ3YkjbP2NMeo3qOetcJZ/njee1KrbMZYki4OFgW5/0rNHC/pO
4csQuWjI8n2L11JxeAy76PN2PAMqpiZ+v23NFnSdVnFqgMkn91y8H87zixvwivcs
A46OVLb3fdXXJutgvipjSiJ7N95rmb7zvYwbmmmTefNLa66IzP6zEnkH8pyE5ms/
dI6nR1EmkwBjssKfbpL0glI+hnHaLZeqIfmoffoVVLQdGuCpHoc4h3VWvrjYBkVv
FsXwKJwUCbpgg8R3R3KxnmPlKJqGkpyadg/0XoVv/UKDnkYCUKZ7//7h79TWYQ68
lrlTe3dbM2IzKCBeOVd4TS31z4qrjqahe49Pe8ozITCyFxI/n0/oNkaLKSe7tgof
3gzFcsKaY8U2XKfWbo2sVvQWxuwHUX97VjXIB4YOFd5hGMkt242BnxbSHukvuZCe
cxAk/PkC9je89jnmxwVBJr3ldgSfnsxnxBVY46bOoi/+mmqFeJec0KpZrLbQ1lnN
eCXJTxiyDFyS5TPTYLAEfO8cG6Zi/AcZQcO97rWWSsFFcFTsrGTSJRkCKOM2qF93
CDwbT3jk6uQRQXhUhTPaxdfA99KVi11kfoRPp+vebO0JlV9iB8vGPya3SJkifZrZ
n3iUCh2FBLV+7dmMTMFtDY5dtgm7S5s22fcUb41140zPJIO/NMH1vVpVZOPCNGZV
k/kyoTVhp6sMazcLe6rOtmwHkQWvrPeuo40gE0KKaWKYVl09IPpXy77qAzUmpIYG
SMbSAQXjKz8xpxrhCV9N3OdoCglzWnytejZ20SC8xNtOzJgYQItcHibnVj7T3T5Q
LbK9Li75lAqCxAi9YOWZsDDQ8EBB/wMrb830C4nPgplHN0tvgDMiHP6gj4rlbAZS
4DRCra1PRsc0yUGDMWr2/LQgXBob2n8M1ebafahH/9ncfj9jeNIgJI4CJqz8NQvH
WuquDOKQhSJ5pxl8kr+d+fQnFgi2Y/HnH5hvW1Frz0XFQKa/tcdxkz9GLfRwKD2B
MxPVwWK9oRPJBmQO2qBejAO5Sl5WFTSR6BLklhMBYmNQ0nFdupQPhVi+JUET4XTC
VcYXzisn/QC801I9woC6bDv4S7/+95ceuSDsr86/iYL8HzQTK1xgNaQMXrLqAZrG
/fmVYotzN8NX7U4vNZL0xaFYBqiOCo6xnSoFqUQl7BP1rS7OaOaP2e3Zr0rIL/8X
cW6JQI1jfuw3u4M60S+BK3xTeUiF2A1hPc4kLymLKaNnVSzh5qz5BITBI173foRp
4HXiNHChUypQ2bG65L8MDyb4aWBed5fxa8kgxH9OeIpMwuVDBJH94afxlLgXhu+D
5PEqAhp164c1eRIpO528Ow5Y1LNop9J/AGIYg553/652QuoI+kQKSa8Gd8Q65pqm
GhHYzZX/qaWDehRt8hqcq+LXIW4P2xc99qwdEqxDcED68zYcgcF8uAWNxgJpCKA7
gCXtfcuPxE+N14Ej172nYDFyk590vqxrE7x7wAHjgKbZgyFkzUSuuIwsxcyEWfFP
/rr0ATN2uD6Ld6sk2Fzpwau9R9kUq5mvrlezZy+sCLRy779cbqtTKR6kBisIDVqi
q/AkGWxCna4L4j0ejvbSKYnS0QD/NNoVL3hbnXZDzYuFoceakHmoFkVeq7pa/tCr
XcrpNYdsdpbvCE6ivSstjcHyMedg0Q986KeieKC5flLSBbAcDGP3TGiHKMUPMTUQ
DYXd0Jibn+dMynG/Z0/0vb5IWggyt8pEGLwHO9PvZcj9h3JtqMoavPe/FFXMPWcg
kxeUlFcpn4ozjKWTCsOYafjX6+Xj73YtIPEQRlvWKLmvFEuVXAoA0EeIyFXMD6aA
wpGjTpB99g0+CyMl+U6Dgu6gy4ZkhlPFwIfU2VCzIQA1tJ66yuWE4kZfrkpW7frC
23brje07MmuOZXU8MoFYRgVWEH/sZ2XqZMlz1zP4BlzDg3lCteDJuu29nhCFvQQE
MhQUpl28WGZ9N5AEHXJ+X8Fx7ff12TcVOCtyadffBiwT+pOotfmWkmWjqfXzzDkv
pUNeerbY6BPVRCgon/2KuA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TzzAT0kuEuPt9Uy9H6+KVyWCKisr4QxdUvLFKivIZfjYh5rWaR2nauxrmgrv5HJ0
IzZ4ZjIq8+OZFzJOSPOBEfGX2GYzU1+p9Iv0tjD+rkreq6G8qlER5tnkTC6bfqT8
S97Cf5K66fLTk0zI0jA+FUNZ/tMVnuPwBApZRYon3+FgDKl2b6RkGS5650a8gMHW
tyBZGpHgWnEWBzBWBxpl1PMeSq7OOCSALEXApJTi5JM1s68fLMVdY6doQY6/yBjx
/GXvMBXExCR5my3iGczhNXjRVzvjg91ifTsbyq8MGmzts3dF16KhhWkfCKszyVi9
XEaTzonH8wEUFUW9lvqYyA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 38464 )
`pragma protect data_block
vhcMMmP6WfJsJLEkXMqBj1heveBTwdFseDf8fkvVwK/VniGh75jIhmI2TNF9/Rfm
guYo3LMbA/1WRCV8Zt6L3Ga1swO8pp4b7W0ehgga+ShfhuvKpLjeHTs6ym/RdUVP
6Zz+sM7zDiXx5Zry8lxMY8wGDWeQfjE8x2ol0M56DLMQ5NWC27EjC/SmcNLS7c+Y
Rvf1N8Uxfw75sK2DocTV/roYa0EQnPrZeDvyk6qa8vwNTcUuV7ioxYPVBOeG7Eoa
S3nbwl1F9pSf1NYTNpFOI+dl5HJETlY7Y4y77V8Sh+JolpuMk7jvterA7Jx/QaBT
tOYcKfa0oNlRzkShUa433X6MEDf3mzd9Ore8ndmCdpRMKFKb4W55r04OvxQi5mDg
cwnVDX28L8qxRHpNAbUCn14C0f9iYo0z8Z6T6woeqKwsuZWososcQx7hbmnpSqXA
xCRxs80DmwdcFDxZcIynJdsxrFrYjXUZNw2Y+xMEqmt1OwjDLrdkHoiXTb1FK/fW
+yPT/YWWTzcw6kcAavtlVswZBzraEGLH79TL6rPTdwaBviqarlrdYHxvufDC0m2w
rFXBDBPWMVSBt1I5dWt/CpphUp4VEZX4x3AJpR/zVdpYjIafAPVRdYXRIB6sE5Wp
uNc7kU8BDwL+cfnIUryykVvj4trdjQiFx47zu4v48vBSz0+3/hYAGebVe3x/HJxE
cyMgVCe5yn34awUxErHaFbnd1Wk0lzibaO3b1jUCtTyY6/nySEhAX8oDbNkTaDJk
rUAAUYVs2+7I6cu/0FySxN4yJbzbil7lzS6fXntxLiSYCHuCkWvqFA+ZmONe2QAM
tMzqSRd5GQ7M5ETBZEC5RqmUxBEgVv9nKvmqkPJ02pQoOZdlyFXa697VD2tOd3sm
QshremjztvV7NiRPXu445mCFcTsM3Kci2Sk6MV2S4ppPZFh8y7sBycTwhJ0hhfkh
Sfogk7DjZJpbQQPVmFxFcA+D4Y/sAjK5Sd78XRl1lpuCffP6kEeixbX3IUoaiGWV
F81YKFCb26kVxPsmqI+qnhQ66s7XT5CP99ZqX2575GNRcxQwuriqQ8qVlWI+mYy/
ENFDArI8FkUsbcNNfNU+ywIjKziZuxwxYr656OasYY7HUIh4S+v+TiJTjNh3p7lf
AuD3nzOuPZnyNJlpBZlmIHLs8d6hGxll5vSjgyN8MYYMmFHZ1IuX9wxs76GFSbca
BYpsa71Nat2RsPQxpDTsNGpHVC+TvisrhS3OHI/yf+iqz5XLM1liRiWj0TLlJTaf
vfCYEwTHQ2lWtMoekV9t4dHB5a3CdQ9lv8kqBIK9oWyf24mhurQqVwuZkju+TxkY
HxQ1ekG/j4+623o4P/E8F4HuLiJ8ULI5wg2a7IcGlSBd4G+WI6sfwWC7tueE8diK
lZINBeCjGYavF3+RTCWfbBe0RiRp02JYGx3pSQgryMyN+pLQQFmqjTbalsRfDvn8
atxj/cHBRbNhuWrpoA/6E1cBq3cgcFX/dMPBeV19PKPNi80sLbPxBRsygzmnCvUU
WAmJFyx2QYWTe1C2SOFj1VpK8nucbE9PacTdqsuCD0yLhgsdpLDk1d7xr2jedJZk
GkzB+KwWK++SiKjbtjMd1UrCPIS+ULU6cc9T3nBR/gUusCpclB7y9ykFWuVSfQ55
hcLT86SQu2GmmGdoGbiYLOfMsoi571WtCRrZgxre1vTSBVvyrVfuatH0+9zm6NmF
EEu/jcEEqswZolcba5X7fBf9DjBYiWW9TUpl4eqxsFtPcCDYEhxC+V4JnJOfQh2G
y7CgvPtoyet9lpE6/e7V1xgG1JPH2qUBccHnUzm7CH8j/ErzeAEn5wbheaBedumy
DKV/URVw10PrjMyraZ9w1NLxdvSyID6AU0K0eyKX87o45FK0aHAavhh6sojq2aBV
1Nkha1rj+elg9ceNJl7MrisLW1ASs/dzGZdFxg/zax0Zs9tkVMbAK0IhFM6aeeMv
ylUuxCJE8BPEK0J3SjIy8PQ61alpqKFWDljDLUlXfN0HcPj6X+i4u37PRjoYEI0W
sa3YPKBBlTPKb+fGUj6pNCN8stF48hKapIbSxYVPAJaGVh9vhWoTxfkd3IT0b43c
XuphdEzYSD3HYE2PHHxCBTOAX6WKidLpC70wqs768HaB7eBF9I9aAJYHZeqCfclq
uZhOkUykwmSPdgmypPD4mlzgMlPi7BxDAHiJP8Dls/XB0iSFTfO1M/jtyOgyjxZp
aA3lN2O6AffETAmFEJREUob6212Fv/dZgYPXKQpIqs3Xbl1/1ohznGWDfgjdfTdI
3ltQvAiPghobWqytYoyzacH9YhnN2an04iJm2XnAfue2rfn2nh6XUYfxL21eR2Y3
0OMafDT6/p+fu7a0EOCeh0BQkYIef6OpPgGo5Kcijwou4EKLOdPobTjd3YfiTraC
r5U5q5+iGafeC4oJDlBO5x8SgKMfsBAmWWqw6U3Asd6mOUnvBqRY6kT/bVKywgvj
8/CU/MKkT/K+eX8/p9UbYV88HcAiG7F6RVJZPLiERPQszlR87m5CF1/ukR+DfqUt
XcyHdYVpa8CnEjSZQy4swtmC/NWL6VkxO4ibEZsQgCn+w97H5Nhfqf+h+1WgC1I4
4O1k16XvWk20bbSENS48PnfdD2p+oTF5MahaUd3mOVcYL66M3gNSI4HKwHllItoE
id3iYnc0Dx/9pNOi+9g9z7z8FRsNbKEMdf7uloOtPtgLJeXAt8HpBg8v/xlwLaFm
Orxcu1DRFZDfBpV1DLI0TKdxWCJk5ydwCxEnSdcRkOxokXcZ7rCsZJb6KiOkcyqI
81urRq/i0jDEwUdrXWQgUC+VWcjvm1fxcS2aTgu5X17/AyM3VMHInMm7oeXrNIjI
ROZ+VpyxDzs4j3wI5TsYzo6PvcPGqMjeo2frYytHfD5W08Av2N9wiu1ZXkOwBhRm
toAOVnjt4Wwe9MSNFOGbwHeb0S2O3UiasGm6GvKsTu06F+uHUs9IcNAwXV+MGLmK
0tbZ8LkyP8b7SWbqy2u9Mfc2FXb0Vz9dsQd1M/gpbr138nhdlaWZCsN6pTFJA5l3
XNlagQuIbdrDK83BTGLduTWyYcyITtur9A/1//lDaEjwQgpEdu3THB+RUOPr2nrJ
UI+ajgENnlv6rvNUGEnBws2ht8G9SqhuIg4ZcomWNzlDfPKKU+BKaoPiG3M3wXc2
NkPzlLQGuzBHvi+5jaGC4jRTE7wCWNnx0HlYJfdFONR2XILHjJFqBIK26IaAM/MC
atXfHL0926v0JzIwSnxibT3td4dF7rVtjfTMCB/B0U9Zw9uWOepta7Yq/QEQksAb
8AvE0n/Jad/j+0mkN7udRepbq+HAuXJ8SqB7/2kZYEiF5LakXY/V6+wYPyKDaZdN
R32VbCFHHn6nMS5/gAs4Fd68M73IWWswEQwRr2eu8nM4gzTrcInHFpQv62vV10XV
I3ne+hME2AuWCQbO+0gG73ZFhcpfuNRlqG/5AwD1JZgzIDR4iSc8Uh9zoybzL3P5
mYWW6iVuQSy3gZxVAX4W64TgxE3n1+unShWldXiZYCixaWIFsF1pQpjGoWr8Z/9c
Ttf2wTIkVsMN+H3V7CCHs68TxF4C/rJQYZ6pALymwiJPr6rrpuuzLf2XUg2oPAvP
rV168fc2nYV4ewkXWDPJkAuxhgABLMokO0EepgxYv/bdBeZcC/Lhna/vxa+t3sEW
ezX2u7OjnMptGRF5To/cJWHJzb3c8BZKME6GHCmQjZOPiI01paUbFsK882gVl6xU
MiUMZlWpSlm+gob1Ug6YfJmymtUiyBwPeeansqsgWEAX6TCcCnj7jRmbI2OydgAk
IvQmGuHSriF2dOkRECqwlu280vd0PsgFQThoC+kVNoVggzyvKFIgk7QwWGQ+c1b1
p/jGdpLj4qRVlOLg1CVOGEtFcEhNjzA9Xd3nPOcP9r9Rn+O5FUc3HnHEaeFCNZxV
g9+eFjNgL4chQtCvP4OGQhFgBLj2dTXMsNUQtft//KduYp0q4Qn/j7REm6jpjOI3
1SQMNXOnKio3+oeHE7ia93eQ1/e/1CBlaYP4Kev3pzIEugEGq0n71bhZ0Yk/NCXZ
W8VtrHO8IfOI30PUvibT8mlZxsq2170RH7XDaECnYVA45zvpu9lZ8AMN+4WbBz+D
Dr/aEww3oJlFUDGKg0y8aLJOOijrxgUswzASVuMlhrw+lDDfk2T2lNnHS6F1HhBS
wAR4vwVIOTmV3q16oKdNlOD/CtZTv4ShpKgPPtUHL1Y34a0/jpFWT9FKI4MZh+Ix
FqKL2VespEjHGz6U6ch0b/tLk1egTacCBYJvKBTxwTl9Sbhpu+qgiEegyyC+P43k
e8v7ZJGW/5yyW47xPyMBkYEC8XxkHAbpTJ0XOyIgngyKWWcYfcdn7t5khoST6VIy
3Q0hrXopOvrrKHB5Xzc03sgeRHwTS6uRNJBT5z9GUJ18nLgJhFhga+nD6NRrvqak
rHhvw+j/IzOrvVftgRPgoR9uAIlXXmnZx8le5DfPZwWjIBwmI9Afy7mGb5wbfWVt
/JiLUYy02GT7wWqrLfbuLDIlAM12h7yyppGuqhRbA13VfxTIuKzeuEPeSjO5fkMu
SY0et7nqVKxZdfaj/E8eeqv1XxNrKkJwddtNdi31BA+E2flwHJlvV6LetQjx++kx
YaND+bVshH0pnduUKLvQAD78pP+W+jP/Jk4WXzhyVgIRIBPUN6VMIqL6EQB7REBC
wm+Xd4Jm64l9sK361W/5WE4L7tSDB4wpFoN3DGwVlLnPFqq7vf6gmhiBONWNYK6f
sbBnWECWnNOcSuNN/DLW9LfNrSvZCLGNvcJJxH2eERKpekmFmsNskNgG/wvVW4wj
vRbzgvhkziBjaeXp74vm6H08J1rI+SP7sK86zyq5OzECm1w5AvcTsI8GEE9Mrn/2
/rvuSA4lHHJCc4KLISsi1SC3bStltLgnAeVskB16mzYm+sW54z4SjdqHig94OAsR
iyewyW/RShTGL4O/o5DLczmSh9j8lxX1bFKUUSRmPp4uem2ReuGei1wTF+bnPqle
gq13VT0gi3TPmHPyoNY9btqQandMqq4zFFyw/gXBmDVEW/cUolx08Kse27UhrvdE
4EzHIaXB8gbOL5FMXrBzbwll442RuUZ8WSwzONnYsnbCcrg7SDkIXO6B6AR/E3ka
xqkxLaXz1p6Sx01zn5AzbiJL7VFySU09kKN/L4NOQvXH0PVCQPqJ2DGtN3KF5i7I
aZ+5OE/48+mKQjIH2KGP+IIQ/XLY1RA8jIAopOv8Svi69AvGs9DZJIcqcCbD/E75
U2sIEJ/3n/9X0tIMJtXjoHfMcroBN7TWLRMg+faXRLSU+M6/j55LuB2unJw+xjMR
EwT+XYYItDPp/+vCYj9JgnWYMBQeMmKXzb4ZOAoG+dug3n/UuyprIgqE+Sr25f/8
vh+7R2cbQ6j67tYKsOjyr1G/2qYXEKDn3TfVDBvfnbMJwqDMB5Q6jiZ5IkkYM4CC
arDHg3kzzrOXqgWfhCex+Iu3P5ZUhqyrYk94CgGsHuZn0h+hvSim68Yc0DA5DKgz
O7/cato4pqhUpD+UqcqHYU1QdzKpkBXAk5mbqvds2ylpV29xJ9V6xkIFV9VBYH7o
7dSlKUOYo6SbrmY2wnNvearrYSVtuDHHH0HEyXrnfbPEgYIoDjD7GSkg/cyjOaWQ
wCUGG0ApCy0SAKBgZerRD9u+0RwCBdfHXIRFT7DkkZDEGNYp0S6L0Cu9OWJpsxWN
om3thcSkl+pqXDI3EghW1uWZGwALTIbK2Uex5r+yyuPYJCpzgJsuu6Y4mobb2SA3
6/tRnk5NLN8Hqt44/REOXSm8GqT+H6Ugg8g1ThbidxCav3yk+ZFL2K0El2fwAnWW
6gMKptxGTDcQps0v1hp/UBHA8hU7Rc23p4g1uhaRhKmQv28lE4Mhm8TgvmwRzPVl
dMzKHftshKkAEWbgBg5CTIOjQLgIyy8Q6woT2lY313tI1Zkaq7cJ4+0GRzCWW44x
Cw+trU3zGOk+l7dZnQPCttm1JWV1H+qPFMmHJKsBijFXVYynDCPA005P9XUzw1fw
Zd5XBIPghxK8WlAC0Qg7hXY/E5D3+kMt8WhzO8GKZ5ee2flea7sFC6+z4BZulWpV
oDksTbieKBQRuD82aXWBhM4JtHpFTQyHV4Vi6YRjUaayvK991ElUKN+53VAtsZX1
uY5m4mK2DS3EmMSQN6EO/TLc/zsMggek/5WE9yMmIyCz8Pgcs79kP9T4AKGdFmKZ
8yANQFvANBFYgz/DqMsrmASJqcdhDf5ED8MzyCBFIygPUjWmAnVK0tJa8VUPKcft
JMHGPgCNFVKkvR/+tEgTpUVCNYWjEMWfdWfb1ouCmNyqitedzlyS0Zkai5uYMnqr
R1qxmg8RZccCMXLBZKv0y7U9GW2TcNkcjBsnonkjwxnUQyISRaTVPaIHNxJU2Xz2
g2hkLNfuc6NH4q3rzPOa9TXeIswzcWJ1ZdSboIOvJLKphFt89FVzlaMBMrNAv8CT
oFHSFPkua5xUlQoRYHqR1b5xDxxfFHGkNvBUrKJzf8MtYdX55j9TubbflybTfq9e
XDCp8RX5NlKJcpIG9PCcz2JClfSdVy9f29oQRKwr431v6TZo5skdJ25nCEAvsLZh
sd5l+6pThrExI8soDZjVIjZCfe6Nwoj6HUB3Y9OdHTJ1t1/RPE3wEF0Hksv+80Vm
1x/XOm9PqlOuQGhOY2hTH/jJsoP2wpGwGOBnvNnNHcABLVpwUKIUMgMZMwu/4EeV
yHhaTEzkeknjOTChYsoXQXbcAu5tWXVA1qD/mu9D9FwL/WeCWPAh5KlrQFS9Hirp
lTyOB6ibltrSfgkx+o3iXQRoPPAjbLMD1XCdcdPkFFXdad/9QUWCQFdB3xJD17UV
4YaDpT/ziFGmdwtiuA3npZDEkuKXs+FNBtejxJniDGY3ETcJFfWjXtmBEppGC0dE
HEuDip4HTxEfsn2xeuPSY+68fqyquKB1OZbYY8UQ/xnKoHWGRBrVCxHue/vAy3yi
tW2XIDRYYJSDcpk1SH2zLZiRC6PWsYYvDswU1QBGhIa6nufE7REee+sgecKeWdQb
BSZzkRqANUSN3ffikIdbLBnU+M+qfEWEsdnIniyUz4Pcts56zqsrsdJCZa5uFsvA
3jaxGl/kBITImwzsiKPNUNDDCPhRPh41XTbEq5jOrw8T3azkMIkzvHnxySm0TcFs
54iMzRTc5yAAmjxhFlRWpq4US0GzAGFlFLz09/LVSZ6a8BsdNZzt7A8JvciI+s+O
UQlxDpahqVru3RFURJELou+h/k6zkR2iiPSW88mZYGwF1uKIvj7HJaZRcMng07Gd
sXRyvnKK+x6cQl4fMav4SJEE4FCyYzkMUYVNcGFixZUS+95t5yJIigfPqYg63bWy
Q8IRmq6zKgYXQl7hhM+X3YuO8KaE5ZgUe2S18E/Gn8/7Ttixr8vt0iZGqEKi105v
O4sRC4gOcWJTvYc/Hs0NzyVL7zTDtQqXU3+jvnEfj8EHYewxRWFZVNVZGeozwP3d
ZKMOA8hwqjD9/n+p6ZqL8qbqf/WtbFRLb0Iq8ZGGf25P/2eA9xOEnOY4IujRGP2u
3SAYLtit+ZwKwZZwP4LTOi2Ez+VlFU0CeR/vmiH98n2qIJTfrkFk7JYP6BugDY5+
CnxLy2maDfxArs/txw1Ao+47cra2Zv5HwWTHSSF3mMivZEp9K9p/rI1Sjjq+jSOD
1m2+RZA3LB+dSS9DUO0pQX2ngRY8ypnulXWCTrGYLH/Lp5ZdXFIwzQV4xbiF1s1w
ipXSDNptrkfw76uLMEYGX5UaKUOgvPk1vYxrdoRb6htZcxOuEFZLz1VmZEx8nWwi
mA93sVYkIewhQolPh05yDnEVubG7PKQIU/bRqVJqVFwTQieTzfljqttLjWR8GY1/
GYN//GpPjiCexkrnQZ37GYkCUzURmwfUEVVX4YssOwINKWsWBY4U2hbZC0p5F6SK
bmDs+PNam2uy3PXbouvvlpr+X+m4BwzIXX9/94XhItMpLxcRB6FVrNiU+vFsQcLR
OnhgRiF2vnRwfhKkkJle3Z+7jk2L+yhYBuxMZN2EY4K2QdNA6Z3fueoVtRfvMkxY
+fDPMzeEqey5atfaHOHhmOkUNz4/6Qtm1i1tajgKyS2RzfvZ1W3OYx0A30hXHx8n
o04J2qwZWlkb5jC/0XdN435prujGJjJOMrn4Csb1kM8/hyeelEG0i8Z/do+RLGTV
6rCXk/6js66w36d9uknKzUEM0IcgAWtPCM562k6WdMqRugqWNd9TT7Au1ET5eDKz
+KFIDF0x3SEk6drbRgJVeTlfxCx1vUrgxBAIlekOwzQwX0BoVIuWN0e6dSSFQc82
S5y4TLY1Ck6rxzSr8vMEbpj0AvaqfbjPZBAd6IM9p4OueKzNS8sP//t12nMDiaqG
FXmixS1ExD7gydDjKxnX14BuxKB2ulp8GU9CP3o17hKZ4Jj8VmqB13ZpMjeFc280
6mX1N+iU9w2nu1RjrTtRlBWMuPjmKjUdKtBe8XKBQK/Xdnmh58sKxMUfOn5nvapn
9vhODvAA8orbVibdcZUcCOF7KJszlFGnDntlAFPSogCJG5tNzi6DydbE/s5Kvik/
VHm2NFFWNQOnTR1MjZqqX2OssqNAdXm67VFoikEEFDVuJvuLVL7hEMrii27wPCNg
oOLAYfUkeleRkK15YIX7PiS7uPIl+a6zEn6jxKS8sUZQN3N4ataVut4FYFpbqPfv
BZ0ja+CnrqYvCrxTRO5dBcXOwHmSTEGcxF2fvTBJqhhH5i/XRQi8AutrSd6zJZ1n
imOjcLC1G3YdM/lqIVh9KoPL6Mj+39rqsEtDd00upv6KV/b6LhLyWa8QWzPuHu5a
tWNTzQ708oZPzWnov6dioPK199nM5sai97wkhG77VhAHXPdS3TRMlEce9QZFJMgK
q8b2NdGPYHOpz3h4UmN7GFxZKuFvlpWCg1xKxBEZvlUzquMwDOyj4+a/HOnCpU2K
pggHKnG12u5SF7E07QuXZAHNGEQxSSGQG5SVJWCf2ybdoJBzjxVS5UgxlJryF1Ef
q5nFsLYoYEx88/mvaSOyDlI1k3NIsbyB1jK4YnSLsRV0Yxn7nn7SEW0hhc8A7EmC
ElR3/zn18egwYrYPU7HK4gasOOWJXgg3yRuQq3KhAE2+DWaIr63NrVrFvotfOQ/S
INscrpnmcGiLGEv9SKbAFtMVeYN6ols4jgVsuM+hn71fM5VG18wbvfYOkDwGRT9p
rtYTV7o6D33opcXjlP7q5Ncak0EW82vPvIlMeYlTDs5e08XuqInuv9HSEMJ2qwbG
D3jtDOQwXlcS5Il1Qh2nCE/1mypMs5fRNTZFv65pqFohZ3i9Torsm/WzXPqnG0p6
15M++1wPfXCnDvZpd6RfBCYhMnzRFzZLG0P8tQUT9Y0mo6Uw4IqD9IXvwMD9uqiD
kGR5KYpmq/FTltOIXWSMEWlVuDkQwy5oKc8ZaunZ+kldbYfmrccYAFVkWgwAqe22
CadhP9klZ5+UhQWCOZHokwf0BddRFrtdlzjr4CuPwJBcmwQTpy03zARLhhJfiE3r
erWi9tWCqP7JTyO6nkBB+xws7CcadkKIiePCYEPfEiteP9pwnkRzUZuCxjwcCjiT
aPOdB0tNl75lHOEz9GnOPkg4vPF1eWENwyHxuMuFL8TVNjz/Ricw91N7+rvaU+Eh
YJ+DwoQ5yZbAHgDklCzAayU6j+ZnRjRxCFtitESfcNJh0vccmxIfGjdxAhpi0FzR
N2AQzZnZE+FwvbYcgnQUfHa8quxVi9yJhlv1XbzVWkydfcfx9VK9smFJpMc8lF7s
KBD3DXwoxQrfOHDbhsmfsfTZ82zYfNwmhCVx72RaJzJov7EhOHIGMiW7yOfDw/Mh
f7/QZn+dzkDJxXOnCuBrPmsqx1yoIpjtSrAsRynIQqewAANKfy2tu03t4qdOQhWW
WSNAMyOKTW0TBw4wc6c30K06hI0BPJoCtbE174MC7DVTqu34eI85DQd24Ib2TZNA
T1BevcqxD69I1p/ghAD/F+s9qyZ66j7BMmpX7HmoJO4YuQbZegfIrlVWsWGUO8We
QKLELrjOb/7WF1VAker/OEJY2q2h5I/4ZlawlPm8bm/sf/2xLsTS0zqGEx/BI2fw
WUmqxgRewzKTYHrmRUwQOKW4C0X+dPo2n28KjBMNkcEhdmP960Iwdpfi0Xid/25J
PIu+bupeCUc1147fZx9QHhDiAo7jO+IUM94NrY1SVq5/I7plfirf97SBCKnmurNe
cHteXh4GeU86sLeZ92QGkh2xED1XiMqexTW1nJwiQuIVwN/XWx6q0gNZDDeiHiTV
hPqEatTyJd4gZca3/Z5BsRyF6OMPzB9EAUPlWswC7ukWflE+QBLAoxa+6lhzLJkl
wl+t2RKPySQhlp+reUdOMk5jXt8F2G3tafn0UDLhwWp//Sz70+/2fOtQoNZtMkue
PvaUh5HVPGWnl588t6ngyUkA81TP8IDWFYr6weZxHKsPYGjuBJZ/ieTLvHFlrHKf
E6NVFMXoop8mPq0aaQ6XZQCeqIQDC88Lu0JRL+IqRINySZ0OFr7w4RoJWdu6J3Hh
r3MENOD4MzGrSnlXQc1b43z9t2mrKyrWl8CF9I/Si+zmYR6MHZfXF/VsJuaEPNwx
WXoc7XSTsOomQh4n3uN4fBONxSZvfAWiay0EQnFfGSsIDHDNajHJyrb8dXfZVqiy
LIDWesH322kuIBbSyKlzuoPbE5Gv/E4GBFQZzN7TXzUmyWxQDWU0VzMszSFwtQHw
eLbeJG3hNlyGO0Tt6Rh8dvDAuwDwwtXNFwIjBoukOKh/uVpQRMH5dQtgMlBAgiY4
4NkLJO+TomxcK+j+OIbfij2obnowOpJv0koUKMNXD+hQ/SoEw+JhnoE8LEtojKRr
qMmeYiF/RD6v+0vZyeVbeYEeLzl4CPfnFUs6It8fNYEySHvoJ0o722x1WTQjtHFb
Xus8fZluuecjpFmLyw/vRCCsZKGOFXd6CA9PQsDER2PH7NxP+t+nAfB30RS4JlAJ
F2nabYRYmJo6xvKowHhTZL/XX4+SJWt3yVwXQPxmDnqa30As6i6W3N1vvkAObdsi
zG0YuL0W4OdOL7Q0AgH6OmFFiOdk9oZSP+5YIh0vY7r/Zak/4WcXoXAHRKS9RRFy
7OVrqO8KRwkA/ab+B/cGPQdeK4g4mmnjl0ncuL7TNrCS8NTrqTca0ovaaMdjFIVF
cXlVZM94uoIDji4ojSc6I5HskCT11FDs0mO/lgkgL/UrpPM9n9WnaC4MvBbCzhZB
f/kZvB6LvYcYMND7Bss2jZuNwpy7SELsvukdEX//WCTVk1XoipbbCn4zOii7jq+d
o7LdDzZKlckZ976yCKqheR65a5v4RI12r7BDgoGt6Kc7sMrLrJIyCUUQgn0fey/c
lcbhF6l9Eqe+cyzlDdpoHOcVsEDmPWjqQhcWVQnup53bKnG0/IKZbfw2uHlBE7by
w+aZecEZvSDawlKaObzQShEHFngtZ1zaUXiIAcayobgtQMNXdJt8zSprAPd9fjI4
aODcxoGHPKRMv6zThjf6e2IITgwZwBS1fFrMlGT6WnR3xQth+1XlWYQ/yRBPAli/
DAx3OqBIOUh1EPKlMIW8AeQ3vhsJkAqqhBgzS2GftS22A4JxjaTcBgXjFcz1cAQr
cc7gTX2LDibpF4q/We1A5yzq619EKySfUuV4f5BBMcHYOoppq2+T2Q9lHbnU1juu
rMh5xsFtQSCu0/zw3IMoABJaYzF3ikblxVWP6MyuYSX5f0wCyahwGUQH0AaSrkqO
3ooATwmYlVjVWNLFUwlQQj/DoBwXszAaVWxXFd0rPFM7Y31c5YhGjUm4pfNi5lQu
qTrAv6T1yyG0uB61MhKzhyEYVDMEKGsQxE3gKxoXuMSJrBFMq2sAMQNN8pH4sIBj
zWTgEl234b9cFess1LDVi1vpp4Nn8d26jfnTpXenLVHct9qBXmif/KiEqKBytLdl
+f2x9ZghpS5gezPvsXZPfYMYGe8e7Eu9VDShkq6kLDUV4IAMFQggY9yB2WKby1Cp
vHy3ay8kmpBlNvBebmBxRquLoGAKM4J/YgTk49V6iowbPXduVki62wmr+4JNzUgS
MkmndEtYcb1siohNNdz2pbJ/1r2MfPkL7sTsk8jVAscJZSWZqZO+7Ne3oGbp2/y5
akxL//z75ITRDPd+ZiPJVsIuyLRrFdG4HixGOfPPZ6QYRU50wVW9BPraZ3P4I/+E
IqrrmWJJeFvdP0H2EsfS655HcxtImOnvukUvf0DuXC2YlG8pFLEe8eyI/SZ6iAo0
wRpZEClG4UgMF3CbtAqr+Do7/4BAxNP7HzS5ousizqTKrapsz4gdT+EqFCjDF8Tr
P8nQPDGkKaaEnw26yo+Vb/RM8qyzDshF0kosBSXMg59Qx9rqwI8yyo1TTVAGLmrk
cMyyxp9bZwVxSFuR8vWFBcAOkrbrXXmM00KWFQ/u/OShHZdfUD0HPx6qicUrCwQ5
iC9UITjk5f3JM/7kNb6sVcjHi2/g01xu1tzLacpI3lVGWXE+5H3zY6kiU5ei02d8
2Dv80aeFtUTUouQRwKYEkfOl0lG55QZ3PHmg7k38QzdRqst+snd6W/kaGt+pjjwv
olk1QFF24dqjYFhHtKzUYXcJqbPo3rj6MzhvoEBuWOMk4cEGP8YosOFkilxoLmO0
lXm7oXXhXLR9QcPZb4CL34m9v+d8nM+wThH7YjoTy6ypZroLP84BSYP86tE7oi3k
PPWrxAgUjUbmADpne2KAU2OqeDV7jfNhRJcKjVpifjYqmN6ejx0ogHjU0NOVaXBV
GV2eae8hWcVQeRhVdFdBoFX1um92Kwpfhsf79x1dts61NDxj/YXrwiRaA6V3ead7
T0LlnRamOWCJGwmi5kHmXC4pjR9rQCWQLyX/AxfhTqaRTmBMwLqQwQX0wZZA9/AE
mSZBsxfFEFpnuUdy7QdHw/DUlJWWVew5YZk/JMI2R4Cn4MIg+lX1NHAdj/kGM8YY
mAwWWq17TRPaFnF0hiAycdMDRMIgmcyUH8qIpyT3J3lGkuDfrqp5Z7r4mVdo+fri
wQosmw0lHVE9dysAcJpFoTgZwkE5EmtHQWfdFRAJPIvJCB1uuawlJgRaEagfDBhS
YS8IzsllPj2vMu/qQjuhDgSlorA4NqvKiRSTUhX/Il9S/Q2Lf+mfZ+BpzZ6U+P2C
exXF7uZA+XYqoKt7xOi1QX+G1MbWMQNfCRoIw1phoPhqOWx9U6XdneDCaNLbXIgI
vMArvc0EAzOajmc0iBqeRC70iU6zN5lrw/IJhJS38OHBb8/YX62T/vVrFuK+XoBu
kQA/UtP335/Hle8pZc/KlBTGnKOjujZR7ynNiIxBDfn/e/aRcAbA2VX55ktiSQfw
Z6+CCWZVCkk/OSre42Nc+BsiiWlOZuWJYytVIbKUyQ2dkMIpH/mj2FHvEfV0MCwn
5aLkuQfP9m24Sy2kPgFqrIkPxREY07+cZJUXZHtV6UdqbRt7kzrOcIR1VySBMgyb
hCI9xHbgnbC8ZfaT0abwVEgV3LKK1dvGbezy45bShwz+sJseFxPYKhU5rL9FsNql
y5Ms7/jiZpSVIBbRdYFWmQC/LLfCZJd6NMmUnRQaXd4AhirRz2BD++9LOib3n6wC
/Ylc+/4MWydmfnpf6i8X4UNp0CzmoTcWXcO3Lv5a3SPoYOK1HFilRZuvpcVitTZq
p4Oca2cNkDOTd66W8ifKCIuFA5pkM6ILcN9V+6qzdk23fBk3qkgMOEXMbRoGRFjp
Fq9kQ0O92PW8yGYAA68a7eUMUiTv7j5ICjrmE6N5HZXurQWMkwl+PcKtDNhkfkba
KpNBi9xpIHwnkhCuL+itSXhRCaok7EayYf+PhFli8d5prBzjFMpcWdSaa7fu8BzF
tOAHKTyU/u4qizhSSwht6n3/lRDC2fkwsAnk6U1vPIFHajolzqihg3p3zrPCvZIB
bpSQryChPMLkmgzCfakrJ9ahnkmv0BBtNV0wcAX58V/zqjpW6/30z7KjrecoSrOg
+rcqYow1cTWsdnjUkhNqJGOeVQWVXdQYMulME/U45Mjy/OtBP/J5kelEq7OlY5E5
VKm/Bq9s+2oYqhDUCaZjcMElqBDQRrs22JbByV+3GX0dP88dcONINDtA6kcD4dYD
SIO7arslKqqfYWrhwoxtS2pou6NhzCIJGTHSPBekBvSk2c4fW9dI45wCkcsQwwNw
nnfuGe0E/R1qlHMcjr2pgVtQy7hA47vQrz4dzTfYmW29W3Gqm+ZRvXK/Rbzd7Mgq
S2yx5MY+lodO52anCjDZveSQ4hTldkRtMkNtbMgWSLB6+tF4FmHEt8VVvDma75Ik
UCyruYkg2jY8UcVk1DQmdasXwiUD7GLGJTfGX9sOh/rRyIsuWSk4vlS6JGJzydwh
IPgFsSleFFKLdmDp0GfjkgqWUn3Vt0+oyTfzH9LRXY1lRPdD3ejkqTXZ4PKUIiWc
g10U3F9ysXujPCDqEbpwZ6aM99MwdVKuqKgIPFr3mP8Gg56SOZQqHw0tRuIadUs1
7v2FUVhh6w+4VC38Tos0iJvoWpTQ7Gsg1yXXZDWF/2aNMgkmciFKRigTN8TjOvU+
tznyejeEX9oZFPETnPDL6jPdfZHwdQkxZ4hPMBmGH4o57pWpYXEb+8wCPUywh21u
imxnxS8OMHr8/EUR+kaC8xqcaz30oIuQcB79GecPEMc+cHEKh4mb+EXPeXe1T8v+
BJpz1T5QJ06/t5OYIi31p7pKh6IKiJuWe74Rh7Ht2fclmYdsyYtkioN6f9b/ZU56
AhpguelXWT7Cfzc2TcoLO7C07djtCXNn4pq9YTvm0vjjMRTSIOw/ZZjuEmy9o2Fc
Ehkf1y3ia4J0lvBTQg686WC4/GXhpDr7Sk5lP6lomu8oZhmcPrXJlZdEFcOfErxu
DBZW2KefRQ8HdE8qug9Ua8KI2FZz289rb88hspmjytx53wBhwtQrRmIMzgAQHos1
JxC92TzUdraD6s0fW7UUJWbwIu4A6N00YdNDRfSS2PtO54OGBYe82lXq7ZCDSe4i
svsUDTYOYlp8cuJQ0z9jyzsSMJmzTFOF4Bfz4hckSIqoSWZrGhEYxuei9kqQwZ5c
sYw0Yx/x0GPC8wnL8nxh2+owbeyDZS+SqRlaEptIRgd/qqF44fJBDVX1rCr046e4
dAC9CD9OapVaHV2ycRTyhBF81PKOf7Z4qlGA03F58hg/+FVGrJItAARnvssiIi4D
MCLVwNSSX0Iq6/uUprv5O5atN3IxTajKCZO6R2TKLftTwKpeoBJxZNoxOjml0XpX
gcNn3GLkT61WXgphoakNVax/bmkZaKGcf+L4yocY6kCdlkuvyPHZ1VDLsgDwJrsW
2FSrVX0E+cwX71i1BDx3gchQJQEVlXS7GclpidEfImBohS7LADG8QNOSKwJfIovG
o/rAiIjrTClNKA41mfN9jdNJtjKmbXykxxl8DPp+USRa81Rn7crgsn9lFqMIAhE1
UEvuJhHYvWP3nfdman4nP7g8yVfAGdLX9kuOzTtUOEeR15xemjDsr/wh5o+yn8AI
JLIsGT4SmRoAPU/0RXIROCkPVYVxlAigPX916BAil4IxMtuul8/K5dd/sSmTXzud
RvlJvoUPrIAmzm60Uzu1RhCK2DtgMnT5etRt8Q2BFwujBP8XfWaVUslizeF2YBOw
jqM/S+SnB93ExidEksOuqB0vhz3i8VK/n0IX9JsCn3PsSKKCDfxZ5n7C6NuyXQqR
sHjS7VSqTs5RGFy9bnxltgRTW0U2vw0qGA8MIoUgAlFdjP56eT5aAIfLK8pfoGXB
jeLmNW2hSKVE1wpIt0SY4VCZWIEmaLqwFuxdHhNjivy20//2/FldUwU3S6epEpbj
5kYUSl0C6+ylV4R4tB7h+C5yx8WDsgl6BFJhr0IOYHvGmaIT3XOzxovCmnbqp9Nh
jxuJUrs10Q4cicVqxn3B4OWv+7u52KG/yUWodc+2UIx33Um/vGF58729Yk7A+agM
k3q5ExjbPsQAjIb47wekyUVDi6GPJXBRX9ummoqskj8+Zg5Q++/Bq60XMqj071hS
awhWHxaTL5J78oiN6BDNguKMIyX9P2JvlrJl8eTxK/ijFaHDVYxUMgzCfYVn2CJ7
QEs5JQ+Yl89n5AyyttxdoBYUWwlyZuIHxiuhD5phHd7DzbzE6GJbYWLOuKpcZeuS
XQRFtr5hW79CQ/MmLQvWvGofN/NrApIRDAXE4KD7xu9tNoqRn9ILLMWizHfpiNFm
8Lyce7aPSi1Z0j8VC+rMjMW+/OlmkLmbim2wJjIcIvDbT/5gAJAWL9jIzP3+5y8Z
i3AeeOMvbAeLhGR/wZJVQPXTpAkSMspKq3/x+0n6RIYK2ewMB0yO3QG4beMgfdNS
Bi/SmlsMqA6DoAprElldZr9gPFmiHCEEnvRIozADVzjXcFVJE41jySWuKD5HJRUI
PHxsdFlycYxEd6muNcLrc651ZrKppbOLXmTiFDMfWDE7Az+SkTl+uNvvwc+/U0Qi
wDamowt+scQahlyvcd5vcTuCXnQ220YLyBwZEh417u5n7QMkYRbz/3TpG7rKq4Jj
oQDZACVby2WDE/SB7DIzYAPRu2aRS0dMQryDeJXFqIFkhYyUooWpKeapSjtYz/Jq
YqisFiNXGGRvAkrdxKKjRU6BSpClwefBLwTr7kA2+VG0zMcl/SDIbLC0czK72nh2
7wRClR+uikRznfBi72U/5myAFFSABHpwM8cF6cW5mRWHuZS6A2sePnOBZrjw9uy5
XufSf+rOcQb4Qf9DTWkWtKCWOuN3yctt6hr2M2gYnptCHwtWldDlnR30r8sayZAH
lsCsAUhkAHMan5hGHQnewHWNYycGMpG+RmffsLbDg/qQjHJNywUqJkQdpLheTI32
FfQHDto4fPRAWx7NwzdqJp6eCjGpGvtE3eVEH7/iLHDgI/OK/270YhwIK+5Ii6Oc
5Jfu5QmpgudPl0XFUMAYPT6V4zdz18iz460df5cRWU+plJbkE4QfJZYFcVuxRafq
jJv1tcLzTPd22f9CzIOOAWCr7PLyLxt+P9L6OUlSp3Ji9Vvk9ac7mkHbHOagogrT
Qn0Yoy9g64ET+svTS7tgUlFLZF0nbNidgS2OGYBIsUhP2y3nxxEnoyNWcipa41Ex
r+4UJF0htvzm7wlXehEDGbF2bh06wiLyaB7QGHJ+AQj3Sx+1ifBtsymvcS0Vg9sN
I5HrPXXUvCmihvR0wUzu6F0ChMAkmMC4E7OcruImOINuho/sVRwx6Y+7TwddwIem
k+NRrvWjXhcmxqdsAu3SdCuz+7IabhGtt7Au4qTubwuxQAQHTrWs8CXltSvPhcEG
JOKJPAlUlhDWXw5bb1Z2qAD3TkuIdagtBhJ7j5oMfk9tU51kPVLKFsW/EhJJX50L
JmrkhbaXrSdY9t2XalTxrwO57/vJ2XyRSPS2nDSTC/l4s3MldbPUm4kSnS2exgEC
KFPwkKysgzDpZPVwQwxDEZMEt4+0DGl6Co6pXpEsM8KXlp8GJ8BI6r+3ChzbD03I
0OjpFgCIgZRMx2arVFldUw3ZFUp/oC/DrbA+mzpEIctutbVumILFZAUC4Q+e7bm3
NfmvdwYxpQNI506P43Xv1oKe9v+LkU5ncUNHQzdORRwa1jgFOhnb3Idm8f4aOQCy
Bs/hpaIBDi+O/qsuP5DAJcTRS/8FnvSJjwXWKp0r5zsEdm3UB3MPrrBuLX3EY11x
opgoLpPmsW319NAsbVcDr4myiTKW5MVS+ME0MdJpoVCpN+b6mPl81o5Xlmoi1tCP
KBclEbQ079aCzWVje8dOcmSXQ0vMrhiUgWzcXYi+bOPNNI/cuh1wZXRcovkp/sPp
jKOrWqR4MZlVpKH6ksRvmuZS4PNIeT0+rnDcoM2AFv2cudrb/S0YrlF3laZ0FQv4
p2/0ajLBidLZSK9GIWV/DfAQ0yljmZcm2kfcv6JdL1nVfThHXBW3zfdGcpjPzkMH
Ry6YYLEG8RcJ33uUKLVpNbhRoEicVrED/88sCu/wJw83vpNrDZ/LXTf32CTexI93
vZqJPt50CHOX64iANFw2NFXjsvCAF4qKXbL5MdOvW2A/is4f3s0YgJVxYXkfzzu3
HM32pit7oE/cagnZ8FGkQbw5zOMewuT0X13gmEkaz0/h42psBI6OLLkyXdL2xwTB
Yjl8VTI4ry1ccHbaxkgtHXHZR5p3uY8aq8yAum9PHPcDoOq7iX5S6wxDR/M4LQB0
YzG4j3ijCnPERByHjztexDlJTqTagAnhorIbKC+vQu20Bi8BUneGuYNqJiUr66y/
BuILkwUgnPZPFwThErEkN5u0g6LoYewawDRKOuN1tLNGP/WQTHKEN0o6oTsKVc/S
aYKDiSpYKYNGQLW4zzrT/+3VsTHO7OxDG2LoQIZPJPf2wT2pBrBLmcTEzsFWYKtW
8De2CJbm04Ydx+qpay1zLjJD73xDYcFirygXP/G/KzesvINWba5xR1yznb3MPQFi
US3biVqhFcHCd7ybgHnIg99vagGDJnxLdtK8ZyfYJgz0h4M9/+/vhRoGJAclB0m1
LDd2TF4mskmzVjQukQT+7+Kp8Y1HUCni942KuhCWAIwNCk6Hf8xSGAt13uE6SIun
VhfnXDrDQsPsYD4ie3UX+SGW4ADhvROnkcms3pUTyo63Qx6NQoG5sy0uVtceT75R
JaT5O4sknoFi5wUqheLd1oDGiJSoNLUiDUuRBQioVMyrFI+OWIrNRHtUAZV+mpcy
vfk4yVIGRBl1wbRAY5yK03/BL6W/FqRSsb/yQ5ZXL7dNW4crxjaFC3JhfbQcFiAX
4IhJFpHWFkuRGQC631LGpOIjKMaK25OtHjJD7QMgTI9HPSTa0jL7jfi7bH38pxuv
I+WA7ZncYlGDIfSQ/vEzDtKRPRbGAoD6jbWY2hHr9ZRb0PPF8otsf2h3HkfY38cy
HiceA3AO9Ki4OJtVDVEGMy+z29qmfBsl9Sa2GZHGP5uCm+6wwj6fFYg8gsNc0uUq
hy6GP6bL4tmo5C0jkx55SI9ndLaunPfBPVM6FWj95hHPlXQgcf2bmOyFO9PzfLJY
Ldq9gNa5j2klSVXSwIg+0uZJln4cXNdgOynh7wJ486tSvSr9/VoqZoRr35oFtjyM
YJCaOZs3JQyZ9sYGQK7e3yovKxkrqF8bwKmMZkaFZ8qqdQc8UNiuf0eX3ahZmIGK
zD+L9J7EJ9o/zW/WF3JWo4z51HBWwA+ocg/yOfUlihamdytXNDvSU9ai7YU+UpZB
DcOMgfu9No8+xnvUaGvNCnobbjBlTcTssUHwaGFNgkZpm7AnVQZA6FF1B4rNH+zh
QO8+uSeUBvoXYQXr/Wf4VJojS5/Wbw07xZQdb2HLc7wBkL7xVjcaoDzgviJ2HvpW
5ZkxXoT6I6wb1eDgVKIyKTwspHm+hsAfgMk40uMYGGgFFcoxPzw+kFM+lovI0p2X
E95EOLD9XDZMPafCtdkHVaxoKqOeSHPpzGiNPurfblSp90wL2DdTltegw0ldzULD
/0RO7hSuKN11clcJ9DzZn+8X4ChsDSpE0CFZVdvNk6xbmXBq4AwitmV3z2px0txO
bXUmARWizzeTkKOSWO7TJ57MIjOHH921NgcFZN8O7wk0os29H5kExdu6v9m3mles
xz+MNDFVbf/sv/5/3G/hjVAfhmWDjoaChG7FxhIqakOUVEUWb7HH1ClEZRPvmFud
15SDfCcLKYSi+LRw8XaulAf5HBrClatwHCKWh+IzOpjW1n/yBgS09YZU29SOooK0
d7Ek2ghqOtvkrUYFa6rzSEGhsrtT7VlXC+1dshPR5UYKu8kPgoV9236GU5bc43Um
0b5DCV8KhiQfXY3ReOM6mRHNNn5xX9VIxF0eH6JlnikIBUwEqdwmPcQukcK0z+Z1
6FSfRe4n29aAoZSJ/luGXm8qxtGTYf9hk05dOoOQgdUp4M52fPwBPMSBp9iCy8Q1
dT0RSAfIJIkzmeDbXrxKUIHSaCIrmxZ5hwyDmq7Xqr2C7hvP3JYITlxXxmPNsirk
HJNOT2uFRF0Q38MAKUugENtLpLKjFhEHI71dryz51YRBEVp9Y07yeXi3asS9wfmq
ylgHRf9uJ/t3D2zevviDCXzza6abD+jkxHUflZilbsjIZFqyh8zIVz5QTpvzkqqU
AA0ia+4sU8bb2lP56FRV39Ka/i3sPB+zYFR7JqTb30wRAKjB5WLtt9pvqTvZa8kK
pKLuVQPUQ+rfl/13O4S86UoTOAfIVmMqiUqF2Gx8SjqedifzN+Qzh6WjZmthMR2t
CROQiq8M9IlasJkld/Ip7BR1DmfYDicqNnOyxT/DAnKfiu7IsfiyEoXJC/GtJKIL
FV8N2yuzkd5ZUqwjNXVjx9NvtEPaYAL5Bg4OFI+jQz4GbaJJA0W2R2f9rEqgHFpg
2OR0kCL2ZiXvI07kFdb3QqmpXtP27rN3WUDEjwRWRExseF1jMss9UtukhrbGcPfK
rbCUWMrq8d+FhgnQZSy837mhUo9dD3MNYrdznCBsMao9OUj993Z5uoW4fM8Kgw53
K8Hqkx/AyJdU6dEAQCuNu/3KJo7PYMrrr/myU33hf9J+8k+91toeZhrzlh6Ud7PU
pbUln6vUlpba4GiTrPPcWa1ajquDE0RY85N9BPU5tDAgRcLXoOriUiK+P240lmkj
+7l1ZO6podoh3k+dbpOJOvf6yHvUrCjHILCcNbZ3JOUpE3S7NUjhNyinJhiAmOm2
SyH+6UYWkjcszAe9PjALm+Y1Hg/V8c2tMt8Pu9gi7sFo1/PwH7dRQDJNP/RhHBM2
U4Xf8qX6sQpM10LjoLVeWfU/RXS/HFvoflQwT30FkKSbVtKob6S1tkRphTM9I+2U
Ad+5S3m1tcFTKsyI9THHqN+drYB2POU+ywqTifYrGH77RK0CMPueAuYkVCADN/M7
rR1RwWCUmTjWHka6oFn5W0LfOSvj+Xz2wFo3dKcOvUaHOYno4C2mRiclIwqV2fZ+
Ieouoz6OMB/RAxWUcabhE0plWqoYEyAOQT3G1gegiWw1EhhgokF3PnbDzoijJ7qs
q3Nsw37eQs+rZedlqjDjH3KGFgAfXdv/h7by83glc6B6bQenSnveQM6qXFKCfWlm
GQaNJ39EW0Pt0WsMzkAVXBLhjJZXix6bPbIwr4219eRl8RDRwwLKDsxzqt2zJTkH
0JpQ3J+VqFsH8is9I9i7kiuKkvy+u7H1mkcAUjSdmO3PI9jmuMx6NPsZvAW53ODd
hs1wSm9ltMG4o1h0UlaJMcrAUObTVSWg3gWx1Qzs7Af+5JXhmXWGTL806UJUSP0g
SGw+NbzXdstfFDzOlVAMUYL5L9Rd78+8Sgirks2P1OVEEvItcutP/eUnxR0F7db2
fkN8ygD8PCo9D1i++P/VTWiAVjFP2ZcGXU7hCrJien5KveFw1k0c+TrUVJ+oHOK4
2MyjAa5CtwOP1lulVhjmN7hVrOsOY82+MmQEu3cInW3DUZQi4uQHaGP7Gn0iGN1z
KlNyvCojP6ksIHrAyN374x6Jp5JyhzmjsFGglRscGDtXh+fKOVRo9Rnrn1C4cSZC
2bG2lS4ylbd19rKAamQmN1eyhOTA7quWbvAcJfZfCL3+upmGY8JbcchxRICzHEBg
n4zENNWJre/ev1LrHmMBuD2nGtny2NR0vSwasjxFfd5C53vDxSXQRtgfxlBYXFmX
akX6GNOHbm3xDXiDOZp4mFzDkgFmAYdvlcaSZPnGOnKplwZd9zWEPCjBire9hl2l
b6hEtkwADawIPHcEtNz0haEGZDdFHYeo0Qw+rZ2//pNIlCBXc4zWH2/cm2sBNoB8
8eg9rL54qFN2D9HDTzwKih7k5un39BLYj2uG8cKeyjSVeoI+HkxHemblHjmDgvLW
wePQfEOjWM4UoIKWjj+tQqWSV7hEkjy/21Gpu/8aWZpmlp3EndhhRlD1Mnn/nhdq
ZJzLrHXsPopomFsg0sraIai4GVuNYqbT97aKOsX1iJKfvx8ENbQtq0CiE8NVWfZK
R7xQjgx+71X4JpqguG2gb8AvC1DEa6JgmWVHtQY29PPLzQPIOYnvQ8GPlYCjnUTf
cfulmW7N0/BcldwyolMDv/GUTQxGTfeuHOxERVUECcG406C2c44hnwBvsJ+cW04W
5VBkmRyla9WNWV04a/yR504eEYxsXXyl1FGB5Nc7KaFBaG9de7TP7wwHl7F19TT/
VIfwiEXW48K4u5sqMcZmpUfksONTPBWRHfsvHQtrKFyWeCMSLPh+SmVGDXq+IC+/
b5wuklcclIadBYw2u9JxYMQKAUkMjeerx53NYCARVm3xlLE213CTXAT/FZFTJbGX
+gCRQc853OFy//wu1bOYnhgVV/ogRRJa9076ypU0iSWsaIXAUJV7gU227wtl8o0p
m1R45WOwbrjOYVbrfrkJ62wHNlGE30Z/DLvelwQ7HFT8okwNkSVNIoH71XbhjxTT
NXu3cDoFAnsgcgYLNJF2zwiww6F8rIfIkwIvD0fM/BBZprugW5i2E7u7xhNSE2ny
hPYS9S2jumj3LPUgiTuzTlBjNGWfgQ/raDFtXU3/PxFeeEZ3RSWafuK5hDMyujHF
6cWKoLDEzRf0wO/VZ2D6WajvFS49A7pmrwQHiIJeIRnz/zDyQ564rp9NPThF7iBQ
nKQghB+ouVivoWImO0OKN7jdUnWKdjSHyaTtKtW+91DicUI08cn8gcV9MFlEWNo/
X3LXnBYoKNkEBA9LN+Nw0C7JcE/MxAeUq+EYHRerXVsZmciAob3aGRF/4Pkg0wt/
e6ZyZzmEhfzkK9b299fSjNNziIX29QbA5/+SWhFoOWeGzaIE90drSnEj+wJ1xv+Z
dyezAVMNqHv5LgjY0Mt7aOJcGWtVU1XZkeOKYoM61V/OyuJDOvu00Xef2SFxAzYo
nBQ2vju5eGTnLeQJRD1nHedX7Dz/0BWrDOF0vuo/nwYZ1RH5PW2Vi8uLm9m6RkrW
j60vWJAz9UOLZsXwpudIcBbjOnBUb32J9MKBbpDhK4ppvBToY8dIk5Zts/TCilGU
rULkc3er71lvPB5iHR6E+scLJkO0+Xz+n01ZdoDpvP8h/oaQnBirwLRqQ3nwi3Tp
Up0cNY/2xhAKZd1LTg7kxb5wm8CYGjsc5uligaiKquPy3+L4+hoOgef6WZBX5zO3
sG30IwcVb+rr0gcfEGGeR5v3zSV97MwzBvlrPQUXCEgdBNC4Vb3o0l4uGTJHH2H6
BTtxRZHJdvFnAEG4HI6gehd5TG7m8SZnPDBQDwhXxXvsTmzzvOropB21ejwPh6Fn
WpHHxc38/DlnxcDVgpjIEhwyfXUWN5rkH8harxDpbzW1ZR+80Os3vL1kuvKUxxya
LlFw5n9AnS+/yE9ShmUQe9ZPIqXXR5F1F+t0yply7zyQtE8pSNjoeZJBc6s5GnXG
EhPbU1IQqqQ3QW0pEbrYKx11/5McI4YJYUCtTV7bjUtZdT2E1EVqabxIdOj9WWJs
hV0HqpXUzJy9XCtEXKWNpjV84XYUxDDMoPquq64LDddZX4NaaF4oz4vssrU/0e7d
Y19wW0WKsCApLhUh3Q8bjn/f3mnK4LlBl7Kx76Uwph4ouxvXXURLXBeZ0Vbwpc2P
fQQi0f13Tx11kZ1N7YcH0uWkoz6Dx3vK5IsuLnhiOGg8fI7pSRIBtc9KStHVq7/5
Hqb2UfdirV4onKW7jbDSxuygLZyqvhel6OFrX7Qw2U7RVLI5s5pNYg3R1OJAhVKw
2Nd38lhFZO67rqTDj2x7EZjzCDYgOZO5SKM+1P1eGK2XgSPb1wcUAdeHdQkyXxdN
VZEAztfasI80WVgvINqNebUTA5vxurVADTTZldTN8knStOhnhvpdRTV9cInC/dow
9aF+PvBWj+2OfbvCMW8Udu5h9QEMYhZwY5JujXzgKyANs2V/aRTpD+buSodgi3rB
0F4qsm/VVkmLVoEIiTYviOnOVel6+qFkFXqKYSXwP3Ld+luvgSOslImHQ5DGAW8s
W13Aa27n8rfaJmuKakgKfREEqeMW1DmgfGCebjJ9CPCfJR5fhIgpk2RoN1yY3Jn/
ALyt8H+8Pn/bjOW67UNFMrwP69SZOjfjmiNmeEQ+OdurksTwdKrv3MZ4DCBGTDot
Y372VM+DqOYvobwk98nsTuxBkC1xArFClgD4zG0G2uAtLpkecOZE5PMT/gsN3XTI
sMMgZMQNCuEUDV55b1rCyDW7GhTKK91k+4WYZ2TBhgF0hRNDI0LvN89IEqitDAaG
TDwQh8Uyfheh/sFML4NR7F118BbGY0mgUWOfZfo9pjqG265ZRHZlB+kDNEKRxrJf
85hSqm3iOCE96S6kDxRS2zakcZixoWvEgjjYfWujPT8r6zpDM9MRWXIf7Z1KJWbv
rDC0a+yKAd/CWUHz2Kn9dX175Tt72QgwTB8XvfbHTvnD7FTi8XZugoM6xrs14Qd+
k6ZV0F4wj44zWAFCaCqerI0NxF8DbpNgTrioSBY78x+Aiu0o4eAgzkD28Zv/gI55
dczFtnuWmDyXXg2mEOeulCwEMiZejFJNWYv6zR5LiVNrX2+lwcBMzb1o1kYv/6rP
iAN+Gk8gvaDuJJ1wNjhbzLxoz0bUWW/i4VAY7r1R3EsjrD9z7WF2uwSX2e8w+h61
74vpnF+Kj1uAIfgFlpsvQHZAceDDgStcd45NfX7uL0+VRhJKPfkHoLCjO2vZUvwl
uDBueBbvL8HhA/BDAGncVp1AskKlli+IQ+YVdEWOeiWeWGKyNp+uw9kYe45uy94p
XNozPIJvm/iELx6Z2MycbntAgCiLNRS0jA9gduxaKsGsFdrv0bKEVNY8o3+JjIzl
O3uavYE1UJAj/UanWDGRWLDqBsBpmz6HLmxcNECL31OkkRpjB46RsIB7ZqgWOJ+V
YnTA11qkYMjVeI2tDZEKKWo/px5PzXn4gVRfj2IkgI4yZLzlN38Ku/ouye6L/pZu
HSKEPTNDkTloQ1/H8a/Gg/UtmajeKWQOxX75aHR73aP2jxjk9R7xpgiolwUQWQi1
GF9v9+gmLWjLvnYdojUaES/bX7CIGObD6OeKLZkVpoRamImaxkiMqzBTp+4LeCE3
cmScyR/ofaAOb8VyKh4IT485JvmXz/dTf66rlMcDcCYVN5n+l4Zh4hh5qr0YzFi5
ByLLy+mTuv/VE5NxYAFQC65cF0HNvlGuUqkbKL/ITM4kODG5U1fJw53W/gN+ZTH4
mrQikjxDn4eXi67k6UrnNcX77JtuLbhNAUQzbp+Lo/b+8MM+geqKD7Cl5d8jOmZG
2l1i6ykoUIzRAV9W7LkxlUspO5RIoMxn4hjiWjJZaAoxj788r3t52AtW+93rhv+C
sxDLxmfgCb8cwfJ+zp44k2n5hk1ESwUxfxCfTtNfqxOeG5U7hgvcFVYdlcnVJsbP
m9Q++825AdrpZ2A5jAioq5XDhk+DyqI8xPPV9c/0pU9hsm6FT5gmEC2s6kstk8E3
WnYFffnlx5GTZyd4/a3dBuDxS35xobJwZugklAF2Z+Sc9fmE2og6HxSHmrdAbYkW
VfmjLmQk0kGljUZ3HbFWGmoAR553FkeOhzBIkdHfezvnKa2LGzgw1TRBw0W1Iw6V
lvEXKo2QM4iTYJk2f74WMbRegmgynyrWiDCIWXZY/o/K95zDSmJ0HTlMpA4mWdv0
XD9QtNEolvTtrRPNJqbE0CoL2l2WYLfJXU8t2AMnVXBCTlhHFpA5d+ZGdzNKwEy6
ht6tQx+YhFwNVMBMuJuCOT/Sn0ofciDkUWRynl54KtK/wnGXSOUE+TwvN1TmaNe0
KjrWeSzCf2fxS0TRxAexmkDoC6s4dXOcWQpxqTrGkCDkiXD32SyYVD8okYpt4k0j
QxdemeqRETAsG2U3CoKq9H+hCVpxWvo0KU/266UCcZSO2gecWohQoAZpo3rzccS6
kHTM0RWl1xLnc4ma28F/veXiIMjLyQYvPkr8kWoJmDF2KFhxrh17fsF1f8xV2rh4
36ht8GXgSW4YMEwz4mmkbG9OK+sKbSh1aA12vxYqJiH2zzrBMyxbSW6/Jy64FDnP
C4SbnuUWEqyM+Q+0UT9H5nCKmleD6y+IVjMEv09zjLPqYcMpZSlhaiJ0AWXCsIMh
2HidRGhEZ2qCtA4XG3m7tOSkvV4oqTzRkFd4PB3gW39+xYNYn5I+tKXJBAB079NM
ThhNlJ18CuV5WP7OnPoDL0oM+RgQH92nJClvCEokaN+ZEKhTaHsHJdUq8tUZtPJE
8RlKlUqYN30tiyKFy+ILrP/LAuKOmqnoz3ji39onRGfApz00H2Eylaj5+6dOdUTO
nJgiQSuoIp1/5VUgJKuX5zE1AR5LP/Ayxw6/T1+b+/Xnb28C+KzuHbmIa0wHAtLg
HDh2jZim7NH2H2g67exrsDxyKh+fIh6c6sCnBqLzC5+8BIn4b5LoL7j8H0R1LRnW
nmtP8cRNr+BS8jXOKyZK0+UC5oHV8ZcpD5iPeNs9wlLDulKRA/0EpKoj8IrzS2UG
ZKgnuLIAQsto9sJuMC2jPqhVXiwra+AkXdBTKv6qLn//7vrb1+ydnWy4wi7lrcW4
dwt+q2I+2obl2CkM80EKdaOsy3NVQjVsTPGT3jCpyEKAjQAbik6QYtwfrV+JPYmy
pAnQWGr2ca6A7NlX2bXFPgzbkfgXtBl/fo3g/V+6+eolqnzdjQ08zmLHomM5Pk6D
lMsJjydsH6aVKeuE1/a8I7sHLBFgWdJa3V3xklj0lTdCt3Y0W/FwVUQy5f86DAm8
urykkivT+slYEga97t3rH8wemiEtMKZ1dvvKLSmNooRUL2F/lJY/KrKv84Ppo9ef
SIxKNNSJ3rx6WPUQ6QWI4Ke02LcBK+OEdZshAiSEa/tGh9/Uxi+spDyUukOYqF4X
WDqhmgx7mawVfkv0q368/Xw48cF+f9u6WZmf9LLLs8U4HcLTj3mx4LfaanTueszg
6O2kJ0zGchQyEn0jEPbo+OIcsvZSr7ZO1kf6tl2t7CjzZC0gbIVZrS5SGknX8gzo
FmRy0zaWz860fSuiQ6dxfvE7/S6ELQ9TYiV0xxLW63QCFsg+tHyqLC2tIookU812
SphqQNWWTbt1/YokAto5ii1ERIst5IOpz7i3BRoSs5gpp2kD+hysg0R2xoLSgCzj
vYh9gjosm2Qr37MBq0fxh5Rn1PJLrbfjLOA0npqlSBAN6+kC7dFcnaVyM8bVEgOt
u2qyCcoOpfQlc2LvS8c18u/9KQvlIMHy7HPYps5x2N9o7xPYCvQdNS+9zOjWwy1X
4T6VdKVyI2GGT4spze9GqshsMWPwb3WZfUBtSetvF6EXPe+je5YWfaIRDtdjjxKT
7gzQ7jFFxvkns8PGdoY6obJvnQvISvXF8ujj3V5sgdyVNCDNglSjJGJifhRueSS+
UD0HpQ7ZuZ/a23+tYlgA/proUHZ/sd+YqqHG/PP2R4Z0Sp1CAIqaXxqOcepK1rr4
EKMCJwI+iZpSdODztla/CpCmD3ZhARY5n7wXv4I4eTpSl+KGRWV0Zi5efKxp03TQ
4JdjgE5yYfBbuDEbi7Vw71Q5G+GgyaP74RsirM2DbzDHKclan36Wp9JdxpCrJ1UC
mb6ap/nE7s1v33+UiJkEKct1dIDJcF0NxeIKmVNVpI2BtGp/RcSWT5UW43QsIHPg
pj/4zJrGq6hgzFnKeRn7uHnAbkmEXptnaiR9iroDRZtpfJ9v7V2cjBMObbb1SLXO
D3K3Wqtm/BYn5ZSsgLqglwRInInNWZ9kMGA/1CiQM9q6GG1luZ7aotktFCQVufhv
fCUP1jDP8QMOsffKEJG4eNbLPUxV3u1xGwXXcP6nVcoqn2WlKVuQo3oZnq/0+8O9
4NPK9OH/xfkG5i1gV7HGJ4tzcKjgs9qeoJPZ3URvlhLw7w7HtCWDFluSYa3eBJBX
OTImc1LnMVS7BTGEXjnC2q2m6NzhtPZYeAGWilKP8Vl/w+NuH0psB8Un0XLzUC2r
LQluId8apFKLjVpDKPFnF0m3N1e4lVYii0DvzQG8vW/UdocqPQoRv1ww+38UKltV
S0v92MkV9NbCEkyt0sd+S4BuIG01pcFQateUwZL723eI9d8U3sSPkoSzMnhxmwj3
1OU1PAlQi8hu8jG2LOMdTX2DiuaHDlIoWEz6wO/81vGYQYkmbGEAwZE04vdeTbgr
Uxt9of4532ZqTd4bhsGR05NYIUDawk51SIS75SCqLJDreHHRv3AEUQVdQeK7dWa9
Wa1M0KJrJrLw4vOfiwBx4FeZW0yy0u0+RswiloO73FQcqEx6cJKW9meMxqtjaNUx
poRxxiakGBLX9XxA9+AIpBMNyb/B/mXolhcEQLD16xoU7mtYF09IagQLAgypAe4V
acugeVXlu/+sTlzNMpyRLFiERd7bnb6w3IgXssF7YEa02pNv/K9zDCSYdNdmMlDk
0NCPvBltAv26Fa4gvO11QE3ozGdgatyYSSfL6sXna+MjOaNYPczO3I19uGIoDkpm
ef5uNqHHDXC3KmReeMY8qFwLR6/FZvM3Ecgs9CTa8et0NuxdKAyVJNfWzlu+t/Yl
QlGJel4ObDvFYoCx73tolYwNOwoha03+0Q+ZI9RpGBXBcpiYyJ0RIYfpVC2lncrc
A0K9XO1FolkJfWYW4FtxkpLRsjJKWhT1lqBmaXBrtpw57LQe9bmzWi/xx9wBheTy
VBOzdliuspgCpSnbC3ltH+Q5lOggVAsn8odnk5uKeEfH50N/kwWIDZ5oi0/swQpA
DvW+aTxMzYySLf+84GGAsknTJRBBDcYcKJ0XIajfvWUuX7o0ep1XxyQfsYYETI1b
2g1fBC/1vpCLClp5xaHJBzhKLg39VJ2HFkQiYbnp5cNN+KExZksEcPc6JzahVZEK
iSzCdOTJVOjQIQrsMV22rIYxrkEhrNG/6zXA1aAiXs4wak4stke1QGbqavk8C+Us
tPKnSmwUYKFL5f9lcMYO7qqL5P3uPiQES5N8/QeWRcpgqG8yW2/br6Y4kNXLA2D0
Vz8N3Og4KxhpFzhM116P+s57iMzlviTHEE53CcpkcqCLw6fllZR8sSPN6b8KrvCn
e8xonVz0g/yPGj0OV2BgTtk68b+MosEBCPgpaus2gUkHjWfhenxLSyY++fBWjtac
b8rvpwHhu1VHn0lWma0ERs/HQNXpESpjwLoOlqPMUMXWaihz8eAPbRwwQ58aEHrJ
F+PZqKX6LVIaltWiaLo30QQZ24fMN0u0PgQMQzKiho5oCgGg6kQ6Rn0AJEELtCQz
eCL1IOn/wWW/R5iFxRYj5qH2zd6NYHYM6t7IJW06/7H0ffjPk/oIhBkv12UEyHWg
ztDxhyIxAgPNkJtQ9AbeeojeI4uv7e1PdsXkXLJeRqr3QNB5kyzqMItLyKOOfiiN
L+k7p8BMoee6B1NAqD0rA9lVmKl8zgwk4dm+t+ffeT4MHxEyyCsU+CC2c61Ydswc
2dv6k0CfeEldD4yc4ekN/SaPHF0kIx80nGKSPyfUTM6Hnm4LAv4nw+3gllQ19sEM
CVZC2+7N1y7VlhAgoPJCihd2KsmlAWRJK/W2Thdh0o0od9lYoUk7/nBNWbRiK+k4
eAJWv7hhWIg6lWObHezghteirKcBgBboXyNE5ffaqnbPTdiX+YmV5mbCY/1B9BOr
5NC60WKFpZkKgrvSYffH7FXHl0bopXod1FQ/7i/CaDMtu6fHals9B0hq2LcwqqnA
HXOp00gOWl4pqX53Mzju7mwOWo8I1ZZj8taj7vgz1cNVJ3U0hYCk6rMV5oq9bE5O
HIm/SnlUWqjxN7GlUIsytEeEH+G9nY2TLyjO4LG1Zl0T9LDf9FuK7E8iQ3VYtXl6
oqCE4iiryf0AzHgyAMcWWdWpO4DUvzMI9F6FQ7xDDOYN/JIZ4UfttDp9ACQftsga
gT6ff4LZsDXr2gBrECjfhKykuvp8ZIlGqMk4ZFkh5wtuGuU8GEEtk4G2jKjHXfDB
v0xbLbbe+rOeX2iwVaxdj8VH3n38W8hdSLnQ862Iw5SacE/J3fJNijW6exneiXsK
p7Z85XFqm8pmUHBhPE96h/WbJLlpkgjENciDOn1HpuevrKCx6VZSNNBp/Q0xrjEs
fjOnTu5/NMI+pVhebgbLQcHTdrGwAGFc+asIxXRKMcNG/fPFFjqlZW+OUPMvX+o3
EzXOxfXePWvrCu3ySb7Loq1QRGgKOOr4LOIzGNd3CFrTclKgO2m/XFxWRI06+VUF
qjc8hqyxQljNkjfowEB+jwYMPyUlAUpeVpoQYyU+dVORDHb09MywIZ2enTZQ2cIO
DcKORtkNYRMcPk03tJbqgk198G2h+mJeJDq+BvwGL30ZJHVKzfeaiNq/HHcua8DS
eyvEPPzaAXiWwZGsUW/3hwRYDM8+i71KYvQlnUbuGukoj3erQiHoIwPGJJ7toee3
dOoSQzYzfoQBBfj8W1ti7k7kmklmBEjI7WqBiksv1l/yw8Bvu4IWVDjEEjga/isl
ozCUCyj83DSCQv2wti7tn6uMG5rc8qm/MCOLdcIE2PSKO8g0k+vtwDs5K9hEr0w1
rH8X/Giw86W7pAVIf+mk6Op8oHJmB6nGFI+gNa51oOVdzjYOKHsxcmC5XG6s9u6L
FH+N1JdKgweCm6TdZxDko67Yd97W44TNN3oTWbdjW+IIvbw8WnLAqKfiegotNfbB
RuIGSLOroROXNaVsLGHPb0G8/cjCL5LDR356Hi8UApCLdG7Rfs01FOZp250Yo/NR
mFHRhfFZH05ddhMXcCRwK/VGlegOS90rcq8f5lMB7NqTTWbDaL9azaheLz/mMlXc
R0vwRlXvtaBjNNj/GNsilya56Ki4HIVquDr7JN4Q81YTvKlFTzxBmjaKxivg6V3+
gw7Yz9oyq6jbg83kqgl6/+/TzZk8sI1kY9NJssAiVelPNZnLnvPU9W2IVnc+VeBl
16RHsKBsBgKAjbbMES9Ljo3SMCBpuGdyT56Hu1T/757SfRF9d2e7ewASOWqDojiz
XDHjXJoF7wgnSBUkI2sUVd4d/7XZ9dIf+J5U70n0otReY7ZevRFM7MgkUTw+kYFm
Fio1MQvLsqB2BOY0jDZMcjHOPloGAY3V2hmMryu6k/dgS5vDwEN/2qqh/28MJyDx
Vyl5lebjslELL5BzTn+y/6EmJrxVyA/XZOASTIJHJ9+hLL40XmJ2sKabpW9boHXA
YCBD04PtAqBOXnqCkO1T2JYEWIAuJme7ZkostD/CjjX7ELhEw1WiP1829BaqVUtI
h41pFxID9tK09ir/q0rUJR7xsGNeH1ozth/WQJ5CRTfPuS8Dl9bti4BmnNVBz4Ve
YgDmmt0PrVIw5Iy25fcoNd+DALi7i7LiAdSJqNKxOZte/mbSyirJiMG6FrS3y/zm
9XKgWNzBrtidamWa3J7MXRk3o00ANIcEYeWll9Rkc3srJ67PO1b3/18OX9wQHQ8a
kwU9WbCm8+8imRxhE810FkJ6oYIyMkgYM6NFPnH515TZYUG9Bo+3RmChjfaOICUz
Xpa/+72cSbH0Ut0NR32qsA1J+FgiR0/ZvVKtJW+6RrCs2SIERcLaziTeX95wGAWp
IEskTW5uDxJnZCiqTSN/zoHzwgQ/ifNqwCwOU+zcBm2bBSfZzmzIH2/08cOmNDc6
5nD8nwITtStxZNXlhWV0gRyJmM7MR0OtdnkEmVdXPaQGghAzU+pdKKKsMWS4dFKC
nvb5wUGCfrcM5RWME/jFwupkvkz+DBL9Ca7c2m5nfeUKnipEyxZ2gf9TyUuMyFD6
LPAhkfSPWuS2QXFKOMG8Um163OyC1GcmvKFzGUt5Ox9n8POtFmFymMCoqSNtPoyi
eoSzQFw8h2YGG5fg6UaQ0XXAqq7Saj+lxBjg7LN36aZCIMKoDiw/jiI+vsPtPeBy
aRGcDL8JBpgnmr7xiM1ph6JJCZMEX2YK1bNYDPUXYribK6ZORb0DUIWAFqU9v8Rg
FwpAI6ksDN1PuH7HsWBwt066i/MXveo8pV5Zzk47kuUn01S/vGFHpeQ80utap5Aa
r8cogSLrfE5idKWnPKAFJI16S0qlGsAPlyxTMiwNF+GNLUcaVKeYwPEmYTTv0znN
YRJsiwCNwAeJszc8YMxivxfRmSB9lI2B0fvmyb6N2iPP69dC0znxYWafS4xT7ofv
YhgtOinr8niWUyhA1gr6TgmLH0QBbJZI8NRssjIV3PT5y+SsOfD5V3TCmZH3wua5
H1uq2cFRCCYSrhWzHwT2wn6Pt0c+w8nYp13ND7VKlmJPaZ7ZTC9wrnJsNpy4HzPe
qY43FaqL2GTJ7NEKFHwYsUbmeGSoiCHhND0bBuxPoZPFPL6/0BQoc3Sateyz2Lz4
8NaVbjC64oBt+6l3cdfOYrUXwd40TVRysJWKVGMXXP9smjslUEUzXP2eV4UlBOE1
b2K4O/21iMSiZxX8HljskueFvpsbgOE0uozIsLMz7IcuWyQWjYbLS6XFFEcIeN5G
KG/ezON5N8aJSO1wSYXtbboxmPqJxC74cYGEbRacUg2wzfx9DWDWrbUGz4XDRt62
e55oBMSDkEAp4K2TnN+nJUEDXUK1PYfYOtfx3ZpZ1i3oK2TUzvDCpDFR5IUvVscU
q8pORIZUA7OC2DVnIzZG2a94FDLiY7TAuw/ehfRQdkO+Z9vTdgaM8jJjQFrhdmMr
or3c0RFaXrOSBi57Z2/7ZnWdnMfS05VJpdKY8RgGg9TcAiq6ZvuKbrnP6b2fnmFJ
Xv7eFo/oyLY6vb0DTTlYroSBmEPlmEjNgnCNoI312iZfx+aWF6K1Lb4dvq5QqCpc
hwVf0tJSOX+zJbhHLDOh+d1YlWMAHN2zqShw9TS9BrHTOvC8qwkEunz2Sp9+JYts
kk/uPge/TBezZJevP7OEkbO/uSakf3zCrLuYVdOG5M4j+ngiU7aNENQ0IPzkNh5a
hVyFmOal+cj28hhpgL1Gs+rmu9MmvkIRfwu6udKr8e06AJnJzqQZhfYEVcAvwfL5
ZPTCiDrQ8ylH3rntkvrCTYgul2jH51QtvQer4m3COY6yV94XeLUNVc+bYKe6pJDc
U8CjmyXE0q56pJl39S4UEaApeLNexrdcCbxgqtZklxi24S8l/txsUuRs/iLRoNeL
uXy0/0/PlFRybs8ZQKQS/Iz/ycYIIzzDfRHt17WLZdnzu7BnieH92QlhLaEU5GYE
/C0KlErYQajMs92dXLyigbwrUcgq2EKrymBUeWKsMk6eEjPS6a9kjw4F2Cle8eWJ
J0MrHfzVztSMoVAnFmW9ySvYG6Zs0TTqlGjzywlGDs6O4Qpp+OltrOypyW8c+oAt
MRJ6CS6JJheoqlu3EVvp3Vdk2Sj9+WPQr7+wKmu9oVpVNXB7I7zfDxc0Aw/W4dF7
YdUNqgDwkMydAZ956npHNmKA/CuWDi4VZmqvQZbT76afo47i/mbfe+sYgRH787qz
NMWs9ABosx0IBiMDjq7PrN1fr13bPy3dPWrr3LbHrm9xNU8QAdgfcqUT+x2mVPb8
vX/ISjYdE4laom/zI0pFmghGILCBTA3I9hTy5F7SF4hynAaM0GiFChVvngCt1qFY
cr8lTw7uX1YMr36Kpq4qq7ZGmoRtpHsGApn8mn6nz4f9H/i3Ew6Bd/uN/PQcWXjz
WiMp4712yuqyNwY+kTyX0IndXljdAlqFWtwZ/EusonKNYgLoPQ46KwS1ohEz09Bw
GYHocP52HghptLMUDhPYeDfSQkHkypdEDwsEVsnwlCIjGMCTrI4ZsW3loFVTM3mD
8p5LfAWjH3oF2thnIw5B04QOrA4GupUNE3IQiuOghHAJmjgYygF0n6dDqTAIPzMj
9ESiWaksaDUPVwXoqsmexLUlDyYeq97mIU5xTZOUJeBoCyTfmQtZDBojLB3PP3ki
SDzuBrllEYHi9gsgm6jX2ywiag8/wN0y6DWFA9La2ZZkpEJKg8tnaU8thDT7gE0M
l1jwYErJa11h0jH/Lp2Zs7FGDG1+qp/nfLVYLqxm/geJwXmdZkEqybT3gO13jaSU
7m6ZqREm3JE3gxmT2HXcdC39OzvBigQq8STYRtZ62kLQ52HMoKbt3OFiT1GKsY9M
8A9fuxj8Mb9DwlSHtupxGOIa4+n3WUnXFokvZNF3SpOWYFLT6YuVWHghv960vUq3
D8FVm/Txl8D3L9uofimuwGqHxJVi35D6pw927clS90Qpkek6+vjFCgmZpkO5dw2o
6PipWJ2Nvlnsy6SlmqEKzsC8kayDNrcqPt4euTbZClcU9KNs8zwhHMGtpa/7wNCO
IeHRWX4aG3QmRk8B4HIbs/vQkmVDnJ9UWfTXgNxXjbBe764MW8g1la9rlux5vJuO
wsHszHkp1hBI4OBEuTph3Ody2t3+wW5d2jzqhaRK2f9rh0kKM00ez6BxmHcn7eb/
d9U+RRv15UG+cOLgFI1R6AGSSUwbD4a94jjEF6SoZM55qlx01iggnNojObRNCfxo
PTVoIEMgnvGoLSFgUQa62IJk2jGMVPHjXL28MNUIKJYfoNL3WKKAooJOb/ds86Wy
ML0ibxxy7rhDoibt7UzM9D25QZCvtgOS+WhHfaKsP7lu0p8TBm2c5HHgvTdv7Sjw
SsTOhvsdFqeEgZoROEJ1r+fOcrKULyF/7IiIX4+NJSST0kO5+MbGKI4G+XgFEGFE
Kxaa0/K9p+JYhwEdATHusCvLMkZ4QDw7Oc3PovwdrzLXBYYuUulHpL/IrGiiLlHX
xWrLdhz6NvVWwAuG16LTYnSIW207vOn0UmVSjlVUbk9Dit3t0Or2SOBEnuvBvcXG
B6nN4dkVXJjcjFJWc+IUbftOddFeHHg4RkeKhMG8/eBZQ4JUOgqh9YvDBA964CIF
SRutbnBoXuAZw1Cku+cgzGdo74Q9Y4XQJimgksEfolAYzYHF8W9h6K3b4jK/mOoa
IOpRqvyr1l3xRuYRGEO0ySmdRzC+JuPNulSms+O6vZPvPORQISpbZtDFUpYEcDnQ
hsrku5c8557oUztXuQ9TqVqvHeXCuDKftXwCGFbJlO6e7Sgutgzqz+KE5zUBrL8P
Aq5Bqe/fGv9Cy2wfQkHbOVqtMYhHciDyME0rgBcDNbvky2VUanmGsZzIBccTIFN4
Z6nuDMd0uMp15jF2yUICQ9cbNivpVZ7zn6QwMgkm4fneFrle6Hz3UFrbJoLTuG3T
PI0Q40QpXeyzjFGv5K8mP44JiCRDvebsRIf2pkWyqRZqJ/tjSd6Sq5nkYMY9HT1J
yL9ro4rVPdBIdCTSV2mgiTz4aWsT3CFMAFN/uHXXS7Dh38lYzbGB8bJDN5PhK+Ya
xfirr3OHUESTvnD+U0d28BTVf2elaqbUFlpt372CTwEK58yS0wcvGAuEmmQItQjS
A2NJJ5XLAAbeiSqSOo6C6IiYIYLUFbpxnY7xJzpwkhUk5jJ7cz2lkMWNuIkinbRq
8wUwCUIcbCalWS46k4l5J0UnpMAABy/0GXYkmjvx1bLIy3IYhSxlpUtbLHMlQIUk
XAKMtN+7y6ZA1t3BnTTRL+gnFW/KoPYk5pSCd2wrNxfr/wzDOwzEwJ6pMjpwXFs0
s5bO53SIvoSakfe0JvPVNfMA43yp1xWbrjnZkRd2lL9+rpCG0/4UBUaYYMlb4iKP
36CVaD27PGvumqylW8lcwAmsQoIY5yKJE80Pdd9YwIFPP+3EavSE6Gym6GPsYfU+
FETYaIOGNRwFj0pZpIkN5zLBFQysJkRC2nZW9mx4NT8+BM88vJvxrid7vCFsIvb3
DZ0DQLI7rekxWoK9zFI1EDmrz5qLQ7pGlhDb8pNZpJdW5C60oH73X5W7NaaQ89JG
7XIiKfRXo9Lr9+RV6r1Zn3RskMAuGRkqly5dZn1UMDKtSnx4EHMN2J3EMqBuLK3g
PbEnRzsQ5MMmmB9DdxbwWDPwX8vbm+j4HCc2FmFZQHgqs+MWremT4rMPUgFt3Ty5
o1mQ9QdPMVV1CRVhPSe4Y7HdixFML56knVF13LPVQhzLUZArdSQZQCxmdBHuxdXQ
aXM6FeeNeGdCbns4EPfLrmhE20NOZQL0cx3Phgym/+XmmQZh0DekDA9hp0agG1rQ
Zbh8J+wPDS6mi024xzfOyijPFJJab9no4fVzr5r2B3KcR5m/oIg8S4eTZALEpuv3
y5MJ3jVu8+jmIA3vW7K9mSGGkodQTTtgeoQVxQfiMCzISUCSc4Ahyzs1ZvFUBuwB
2UuUDAqlnp45D7sG3p1O4T5HCIYV2Elk13fvi9YwdCBlkPCOzBCXg5GPJQXTxYg+
RDpP+0QbUw9tI1bJRh/sSZ7WN/aGvhO9jdBHSrdw5cpYyP7lNp/elJLCxGJRFKxT
hk13xo+64bcldjS6rAomztEHMrsAo+eLKfvmkW97yXEewEB4L5ksy4TX9oxWnk1w
L9F2Yf1WrdXTC3IGpoINRn5G1rxXSF+PaZ5AYzFlhJsBB/zSxL40Hyq5XOOJpgaB
0rbeMnFtk6/lC/eScX+jnvO0Qysmf8r2ZaYp5AfhpkRljd2TX+2nXqwUsefz3ThO
ccwMaZI6+p8TC9T6/JjJAlleXwGz/oKGvT/5oez92JUK8BMgxBcyUkKDDRaxPCsu
NnxZFEDALIzW4OvRR22bZrhl4+OCqsz1jHmENgYQtGaXv6SlW0wHu/ocsAaKfHMi
mGgp29bB+LsgnvDJduOGKjRfyhAPDA0YFKjo9XARdX79vuIJ6ISS4a/21ZSdZfck
58+Ac/ydQ2krPm5Bk7C8UNZbtA+SV/wlGSnX9bjq7JZdYsQHzHyHRKG/4dkE0jqP
MtsvA95PuKrE/8/FGMmNX++8cz1cJxdDGmcsTMkv3QLipBuqHwddEi1LezZYakQ2
m14gbyd7V1LMATAZDoSAONhIM7Kv5an7Z4opJZ7Aox2anG47vRXE+Spayncc+8aL
aUlD2HavI3NgJaSW31sSwJlEYGhydEjmbFXH8DAFRuvFMFZlRztOtm83Jre23L2W
69GmqgNXkOz86gsnlySjLQdX6DRzjGAYpBK907Oqtb1rdXoFA9ZIAHM7YV+0z6Jp
NWDJfrrMI+VIJRr6FjUvO1OzumQISsA+q5sUDp9lKhK0JW9rnnbTrAk00o+SZoDq
C+DZvDIuaCgiSlyr0FE+/zTiFPArqRfLkYkSF3vIsLHtIRlasVJXYJXgj+5rYj95
ew6eWaOOc2b9Ql8kHPKhveyAZnRspZi2Q9+O6d8NBSTKWcBoYObcfmsfkptavBSq
AhxgHAylir+PxWPs3oZGp//9vg/YN25tKSR3hp1WvUS96odtSoIB1uAAb4Tvn+jm
S34FzugC6daRIiZGIvJT/r7PVLwKSOAcq+yj4WO+ImAwwoYBsmYJvsvRYmAJ0oiF
/9kgAUQ8JC28wYOcGJLP4mlpaMtpeBXoVMZfMxUOuKkmV6NFGsTfOPKW7KeNDdQq
/WBHqUbo0bqDe/5w/ba3SrYM1G4kDHzH0NJ58IrBGPGpDiEGYmZ9CgAbrc80n00F
73YDVBNL1bkJetpuvF7rfN9t4Ylo/drGSzx3uk3TbskWUyyuWA4WyY7cCwbj3u4C
gr3QojhuZfdx49uSPhniYVgnbsAO7TgxvtnfA0rsMt5Rqh1vogLba6lcDgPM/7eU
VVdb1Q+FqcUBsWgX2GxVdYBkz3FI+ZzOiDoYyVM+YdOOBbG0L3r0yu4XwyfiixIF
oMhxKmj6K1sAH7dJK+VoPb+r46WXH6WuJaSP9NFVBU8OPILC0WEOn7GZyqGznYtl
O1SuDhaAAloIDlCpWz8rHkNISUj8sCu3KTX+Ja+1cIQ26v+2wQWODSnLyQY6Yymd
esAvemPAqQfP+B80YrWHBNWdhvundXPr2rgZogWKIwx6V4hBDtINdUBCXcrs9A6j
K883LmVFiF5QXPoWcoRj9akdZAlX1QDbZ/gKMIG5tn8jP/yrs9Qtm92yy6Vy15Eq
SkUq/7SwgKnECNlL5yfkN9RFitW82pC+7yJ06pRHkNi78tHIO1+Cv2JExclUUUxq
fCboMr/Joyp1Az9C8QXjqJuyL4c45ZeUN7AwTLIqHvuX/H/2RA+B1vZWeGOL1kpa
ikUQu2IhwHVxCQC+ex+9BXWVhcz42QfxLeGxRDxNg//a5OolXnrfR793tUVyuC3+
55LUNPrYySpchxo8kEaII4ZFpTAad8CfsnJMxZ6glytLcA7zKkHBaTWbuZaOaLq4
BQmEElvgCe5Gw/V329zcem/Brv57fNHxt15q+ey5uCOwGwtdQu39n27rdACjuBQ3
VUfkqOzeqSwyd3vIuufBRakxr/RPbwDypmhqHITHWMATeswkXAiKnXBZwh4SODCU
NEV8eUom93W1EBPuQuOrXMXM5vmt4aSZDiJSXzW/EOCTu4jwnD8oukppUWmnw4Th
xXkeGHKX0nXg+5q5pt/iHasoNTHs76lItyxMa5RfYmWZ4yyEvxIHuV5ZUWFIAPdB
qiiSTnwJVw4ztPezbwecveHKl0oFzNvbfzXayz6BzXwPkg+kQoJrd4RUetuSiq5+
jfJ2rHubnBzJ1EaNF2iA//A1t5K33ma721wBQa+xX+IvQEEJTarWGzRuO2rJHl20
xyIsXkZCOyAGyZy3WLUMYnJcFS6E9YzhTLrA7tJFpGun7P4GNDBwKXDsWqI4QJPk
Dm/79GsLqxVyJYqewH+E7d6EThjOR8HiJDmj8u+N2h6QFxuvijetamgau1lpg+RW
8+ZRzT7MIyjkwknMNqVONxY5M/+ob9q8OGZimRQrHMyaQbpdPan9+A/17+/+Y+XU
kG6Ag1l9gxkslBieCmtRS5Ha9K5ItAx8cnD46hcoGq/eOU3KDWa4N2i2inViIHeA
eJ+uqT4N88ssi0wwksxNnFBVPDdT5fOctseZqTMW2Vg5pgrkQup0xmvyLDr6Zb9f
5LZ8VO3mZHLTPOa4eeGMs5eGD/tWid19ZL4hcmYTUW7/L69uvSdxLNIOPlPn/sFY
1Axma/Dn8M0PbR3IktT9qOo5As+soEDsBrZBuKGKRQnrBhx0lGwBEY76OquhQPMo
c0O470hBdN+BmOUP+j/jQ2TOBUkUeAOFf1pPL5U++Qp8iahtqsEYwUMvxZyTx4oA
CwPIdol55dWBz0i4l8igYqb0tGrZ2y+nNlg6JPX+V2CZMTCqYEfMl6rzVb63gL9A
CW8kOfkbn1Z1hb61Na2bmW2GLCUM7ZCMZLwsteOh9hceGzsybhgKWLinvaRf2NRh
EXJByWP331PWrKMZoE/8RRnDcJ6grMGqttPqqfK1H38UR1IRB6053OVHkGg7y78y
/tsaUqQqwaeLt2l/UcBB+kedhxBEMFve0rsnEDIw+YlppYMAh/8zQN5IfbrMxFNC
YEGMQBaDDCauZ4Vz9mpfX+f97LdfSqN5sMUIgpJLXf2jLXjP28X/2GSVs4eGDQom
AeuE5iwOQujdqULVZR9kTVSxFLXsFJLOb+q0S777ded67BXgScmlmuqRj7Qlq51N
ixf8CEHAMnjO7qzqbs1b/IkIseEeS3P3syl8mXvOgXzaZPsKIBjA9KeZmP2LwUoR
811aqR/uVmwg5iw201ZdXFAMXzFWEh3W0nNpVM9UVcV6HMUjLGgnx4QlqMZ4CcXl
Vglthk5m+wC7m2zORx6VdAqEd/A4H6eAleHnOdyKiCrSroWXG5w++2/DirR8RqRD
cIXFEApzUtrmTRYSW2HMtUZD0J6amWQ9eBL6l15FrGR6KI/C/AJn/1EfCxZ9h5sB
BNWcoi6DaWXJNPSjliRjIIHzMKNEMo5mIwg/lqsrrIPEOa9ATNMV7WhRJTZCJoI4
Hpn4e22Q5TicnPFBD486wEiZCKGmjmwfRPQvA//IGz+xg5wbs2Tc7wFKZEP5ddyW
XJW2XRq8QUlrYHn6tXMQCm0z1WB7nW/vH0xmQWz4ZTzmhKoON8ton4MzwOSI1Jg/
mXi3aq8H0CBpW2GtyI3RRWaxcqmuF92Sw7IBL1SA3FLNmeM85TLKuzV2bRj5aNdP
ZEb3ASs3DGaGS+0nFZ1pJyBh/oh00f47DSXsoXahQQDLHZufuq9IntWB1aXIdABy
YKuwR99IF9Fypgr1lck5uinzBU9kYlTfYeHuH08wwHHtDMAo8mi5iuJtjQsUmRRg
rl0LGbmULEU7F7BQz2FgcO1VX5gxfQMaT5BK6+TJxx1QvG7RPECJtaZd0cIAi/X7
clhwYoplJ+Yau6KZ7n2tvw4cderIqiwJq3HCDEEt/ko097rINI73LRvq18l1ob61
xj9dwam4flT8Alth4zY3h2LVbYocHZh4TCFA/ZUw9X6m/GMt+JaytmgdZdXEJDSL
pBm9zRK1AtBQDVl6vN8KA46mujmauj9ShB5/s/PqCq8IOxR9SWYztZwkDBuS1hWM
J5qijnyTQPKN0jH3eZj7zxmj/HUApUPN6i/GyMFTaaiYDxkKaGEAsvK8FYy0K2ye
aIYFrSGxSi/LumjSHiH6mzfXa6B35znPL5Za/UFe1uvXw0AZgsx2/H/vXczRnAxT
nhd/RRXrjOqRYia0bOlrjFIV08mAWKxmoeyCMjX51NLRbLjhXXFzpROeuGo4Q9xs
++y8W/X+f5o0ZPteTQxtFlOdziuwxzegIMvhxfh+2vDGYiotVlOxlEw7N5s/3bgq
sa5eSS5qB+XbFer5eVXJZ/CBirWmACmfkiVpitM3nrQqHAjlGOB6Vs0fR/PRRMYf
5YWm/NO6g1neQMr/RBTEp1NnkHhMuuO+XxKcVw8ZFlWUWq4CQo9kfzU40VT7Pply
GEQYRPGddETWC3tcF4Rys7Run4jCOXlMn7FJXN6hoOdrMxhVZ7tMPiqW7lCfNnBc
/W1GSAhp3/QEIRqCQTp2QMlqEzt7dHQknt6mldlyc6Wd88xapI4uSzREoG0ZmTWI
Kdd+bJFkXgDW6sidYFroRJcgGNYcSBCIzCSuFATW5cOT6sVdf5HrCgFjc/O3y866
832Hhdmopynh0zzkAwO2vlcgsklN7iBzO5bznOmRWVrgOT79ix0cYb1Z98FiWkMg
S+SYUGiDz99/VtrGkIhqgp+ju/KNfPP0bIAxgeZZRQ2WbISNGAMhMBv+6zWtdlDo
QGE+99UF90ZfFWWiTn3IH1+eMprtGo9gUomVQa+/s3d8L7lmEgenq5UpKMxoGY1t
rT0D1pIgnP0Ut7Q/w25Vw+DnLA16RwTOmpzAS3GLu8LOqSTDcqrNgV+G/qjduGYU
U0mznWhyuB36U7Oq2EaYBbBsgbRkZ4kC37HhOXDj1+CZfKzq2Sooxy1yA/Vp3YbS
YZtwHCN+HNTn2wAn2IHiu/N9xXQc2UqH9u5pL5DfnRpeni/M0N8RXY/21udzwkrB
SsfnBDMxy5PR4U39oAZb2eTp9p6yqiQ3KhAxsGJ9thfhu6xZ1tTGCXSw1VFO8b96
5tPIAdHwqFM8aWxu2P4o6diDvkC8wATPJmGBgN0EuQJ3urWOaVB6EJ5UJ5+ZgueM
JWJJz8Ca+oy8XMWrDmeYWVYZSj2lEd1i/5akraktK8vxZOnEhhXAXrI70Tf0SqM2
Eooape9pdqjqo5RBLL836VLGCQpcFh//uLm6otVeo7CnEiqhHMQK2v6JS0vmCJ2I
RhvNl8cN7zQgN42HoGW8onxeyrfwgjwyFu5AktuBIKeaBHhJdWoZZJY6aKA99OwK
y+GXXtiDnVlXoI1ZvvhLvtOw1xLdsConvovKUvM7VJC1B7qAUDtxxgRObmzDdMCr
w1JAsiC5HiuQtdvzrBRaRkyg86qlXKJ+cLWBHoGVXhKQyCTRSjJRy2OAHvOq2x8I
7MgFW5jPr/lZVAtOsWuHqIanM4eC9GPj5EQYkwbLLIgCI2MPOHlLmRqXvG1vzdhi
+aKwzSR8KAlnLCgE7RMbMKy1TaEwoKvN5aRUNtGy8lx+vmtmZwHBWlX2E+pnWHLy
Z+nhXH2hRf1724tCBCvPH6GEhAB7lBP7sX1/OarsDndYlSenoGKF/dqiavzr1qhy
/R7QhNhMyxiBOzAB7HaFKKMW5J7MTQCO77rbOmbbvDUJfR2iFyKsmAD04eb3JwMC
qh+Wn5qZkhwNBa1cTNPZ5p6Oxeiwg/rI0IvcFgtC1av2Q0uB/pZcJC/Z7HNzhGNL
6CSv2tg68HT++vj/SkxYLjVKvbWn3biEFa8uqRZ99yBG9nHTS9ebBqbwpoNQr+LF
u6kDgK6O1kojrj3399H+n9EvgFgz21ofc35JCC9ekq+99p8nBTpSFjoOTuekNIrQ
IRGFqtFw0TN7mEuPta0+qm609+u+0b9dLLVRnQ7qlWI4yZwxwZrZs+HXsVNCjNkj
x4PYv06LpN1Ywb8vFk0NRBSs6ru142zZeHKHWiSpkEee2keQr2uzbzLs2onXI4vr
9qVN9TvpWKlug0ID/nc/QSjM1qZX/wGsWvttCX99GB21pSLQ0hazH80F8iaEIxtq
NIh+Ai7Dpap8rCy+D7AXiwut5k7ovDNYDcKMWOxzArh85sIRJsprGghv0qh/ZQWu
cjjclCBGhW3PKwV5fcjCIYK39WPMtfYK5ApvJT9fR6+RNyD+qQda4O6EN+uCn5ln
C8c65zaCnurIsN65xGjtfbmCKpKsANei6Gqdy1++WbZtaZ2TC9LlVomj1fxzYhdh
6lSbEwbxD4CAM1CsbxD11qPXl0XgpKpkecuBtfxr3kH4tG9rgJ1skpt0OinbU83l
pVadLwwG1ASX7T+SoPZaU6/yIO0tH/yTlIe5GFbrIXzyFjbaZVROGfQMQ9j628dx
5Z0PZDE+lhM9xVKzsBN5IXpH6GwC4CxS8MADdY6QSCEipZ5GiEMVuOMX8wfNKhgx
mYF0DfMQ88WqPuv3VJ26LvokVJinYlOAuJZNU5ITWiBUGyd+YruN8k4N9DuSD2+c
zjB0b0W7d10mryGxDoAB63FKc3JgtRKRERPn9oQQQDE8GR+xO8GRNZl3zy/cCn8U
/jtIxKdGc1jdtPZP8znr4ZF7pvUJ2pBW3O0fbKsc7g7HLRvSzdmHcFLN0H6GdJj0
2xAi68k84jgY/Y/7XrLPPxCS9vaCdCyVslGLzgLKl6Doimnzyh3n3muP+E/2MCP8
lu0akqAS+b+geg7TTmIfVR2XCYa2vbK2IojxT3Q5MVWzmrUNc0fzuwWGctgQHU1X
L6SGbgoEsa29x0q/oI7mHWgsIfGlEzPZPzWLblILxZYNkL+qmUSiOzrXe/+DKGFs
ImiHAy7mk8eAKc49jCwo6kwSvT5zG1vcGhuKSDmLz3x/nMmmah6+pP1dAFFtoapG
WQ4SCnsDqJ7oCjFEvCd3aNfqtNKBEvtMA1RhBOiRxdEr4sgHpQjKawL/paqOCJrh
lJrTn8e9mfR9RVGur3NxTLyf4A1WcmD6tNkNzQ4rC3ooZtM4aTVfbygTBZ5hLxlv
U1+MC1LkqGK12UaI+1gBkdpJ/VGExDg0lwePm/n0XRad4kSjIIL3g9xMmbdH0l9h
+DYV9wpFklrRCqVoAc3OxPh4DocQg0NHejjdoyGpV0+a3MR5m0j+SFS0idPK2r+P
2VtGPgjb9mXWvU9pnSPbLowfv+AWOT1he5Jm2sQdnJiTZPM00WDkcU4+57iR8Aae
my5m/xan22Pg0joiTMGXa31FYuN002/MMRr3fItSnoc7u84KIyPDiMdE20GJsQrt
Ja6R5r+2bgEFRlp5/wo3o08riwgWoZRz6SwGhu8Ejs6UL9gFCxaHmB6KPbyfA5BU
KBZ5dUibjQV4QRdGgtsEcOC+5lG4w4qch/vDrwIB/LKX4I5/F21hehHYZKY9kGy0
0FKiqqTbUbXXD/xYN4vU29XXitF4ikGHxbdKp6maY87Mdz/r6BOJgBIh3DaFM3sq
+P5A6HwLEfXprXV66lV+Bt66mOPheAfUg39Wtyf6bPXtMGKIwBbkQhcgX/R3x6ZD
FsA45//pkT6ePzspuy1KS3dVb2aAKHHmEFV/djbE+UemmEhVGpd2G8TczpA3cE6J
L5BnIAffPjiK52oCCj+9ujdcOBI+E/4cigCe9GCzAja1grW9Vq00Ui3SqTBftn+U
TO3XBQ66PT5gNi0g2dg2swU9Vw8Ll4pEfmyZLHZg7UCFTGZU7XF6X7PpSW9YBgLS
2VgEerxnaPblJtUJ5BLJX7MZ8EpvNBn5X8B34hY+rj/KmMVqk5Eoow5Uu55BHlke
93n4NWSqhp9aXq99YbTo2YX+0GfllK5d56LItD6XlfpWhhhMfWiOhH8KFQLDT8PO
4/qzrQxt8dp9jetmVo6QF5cKN5ImgpMKFrWke/+8/tGkPk8K+hdNDqCpZFD7Dmi+
OUL3D6NC7PjXfiTHc3/UeUsEy1kcwGBwYM2QhVa67UMU9lljSrKdwjNsODsecYmy
B3hnxzyvP1IDP/xxnCneqmK+2Y8YVJBtlUGikoEMT7piIpfBO48NQ4B187kvVj9U
DisgjzbxYlsa/jTP3kU9iME7iNaw9pjYwW13bu5l89oILbdXF3ta1ipup6iQ0upV
rIZp7zqu3ebfDBLEYRhb4nKywsZB/p/lTwmR2Feik37xovNPrS2s5igr0rdQ5viW
77v3DzYmwqzO7BTZ/Adp59nd0z2BvhPo+GRX6ZjySJGmQC1xISBLbtRi9KbTCT7f
7t2ogUhO5Cru2aoCPRPK0r8mkEYtqn5GpgtuEm4e7pMLXaUJE9506B1uytNP0luZ
4t0aIRx9KJ2EZSu/4IC+DEWeC5vh19FlR1QVH8inkh3CwRtmC1jKyJZ0dQ39LiHr
1Oo+frNPViFr6Fe+vIsPaFuHaiKoccdtb81Dhj/J2QlSdlaew//q9jN5lxWAIm6j
tRIuaY7xZRmkmNdjmh198dGQRt51odQ5wTioT6feVQJGmcLOIKGEmFleeNjDY5MR
gd1QullgWCFTt9oSJuNemGUNQRROx6o/i5ZEPYpHj2oS38gpAyUB2Lz0y5eBo2rD
m6QERtX5tmq4Nsm86QxdFri7P8dXdLkC62J8xdMPCxWhivDoVvUHBBvaDuQPxuzQ
eXb+SUCg/8chK2gGaBRKXd8vu1SjinOg7o9BfpShK5tMajQEjs7f0XSqc+t7rBYU
z1ldklz5qGriA0/amKBGYUWo4qcv/U5cHRdtm9Ibzt/y+MiD6+r3ZnBjq3HmlpeB
hn/DNBty1zvyjFNC6YTqw26Ny+/IIeDVE4a4E5RGQls9TvItQNRq/a3HQ0FgRpwb
U2eG9nVOvKbtSk10L5bwMHt0w3SMxzYCrOeI09Ez08uySWwwSQx6X9jF8EPHuIsq
VJku4I7DGGHL9o9QoYat83BP/V6B870IOvpi/UR6D/GwmWOkkCvrA0KRRYD8wy1s
rYoypt7czZzJ/vvS+Uo2R8qRfsXL6R8LZuxnt4V32knBMrIWmyyNYSNFjGPiIQUa
27attFjdqV/LUaUo6BEaz4u3kkfs+WFWNWUoUuMTNo5goIgXc9VITh0sDvQWlc/1
VufF6u2FoMJHjuzyDAejFerrqE05X/9Hk7X/qTGDGPbNG8ep+KryrS62r6ussyDM
GKRi8UjnmOvjZKAj+SO0K34H0AkTCet/EA3Y1hy08UFvZ60000RaxR18RVsEetz/
oIKF3iO1KJ+6/8N2Yyo6z6D0UgmFZkkwIncS/FilZ/9wwi78PncRRyonDFJx9EGd
FUrpB5XBvnPMoXrJNREt9vrURX1+AfUSD8yOfgU0580sY8KS1HYfWNa+c1Au/ham
lx04NCP6hHY12wzEcjWMo5YQ77/WlvMf4lsnYD+EUv37SEMr5baZFbbsEfP0ijyQ
hk/QAp9Y4LHd8QFflcKTdNediBgSg6QANLSMig7c/UAVn3wzEOZu0D0RfYjjjaSs
9J+YTVaoK3PdoMOjVz9wVG1q3UUhmRZllSJzo+0hgSZKb+UUdTEacJV3QSy6ygr8
+jcfFU9v1/aFWW62Tp0cLZG1fIxkI8M/LWcVVmU6mvj/MoBMccB9biKQd/5yVwPa
A3beChg5ldGiRUwiR3qwQKwQHWIZrDBnPodQVrVuKdBiszlBbw8YsdcIN/0S+gvD
uR94fZniJEuY30Aod2a6w1aU2Rmw3pY0rRQVdNObL6GgXYmwYq7Txq+L5RPXezMt
jtd9HuLuu/UwEeivOMewJbghTcuyxGNi76Js5wNcFdrCiFFWpDE+Qc5XPl8PhoDD
KYMERPYzolCpy108m5EiT3rzeH2VHoYKbXpV3tGG8VECJLIAT7GISBIpc0L3SU85
+7BJWt2KU5TG0DucTQMZ3FS7183y99MJt4EqeRL4l3AZPVtUPPMB3blNm2DURg9H
pU4gXI+DazZpBgJUZLy0fo7+1XuhY+6XY/PoXyN4F9i82qKlN54Df4hlDoHkJ7vx
qb21OKMc4+8VMaAVyT9X2CrDb9KcKSd0MmzGTXhuQpT6FJM7jatsIoe3Q5PYqk68
yE8s4iYjJP2GVlUATyWXNILZwXVt7PTZo/LTlBqz9+eZmnN2YndXw7brcnjWMP6H
Q4rokNXZy5ib2vuQ6L7+W6311ipOOEuZl4Dm20JFi/GlfarNpdI6R06sCZ3W/zxW
6r1bZrrCCMgToVX7DLS2fHS2Xsz11UGhFCTWTaUTwAELeSInUBkXczQzhlGtJMQR
1sGkss+nr31mjeOnIIORDkLBPhcyRToIVO0pGyRi+ay9zfCNoX59vF+2IvOVG6cP
vvJmqWrFqOdzRCg2DgddGf+WZfB1IF263ZND1xBliymFmr89R0ai5sWzNPhdZOpp
njEUNOE4+IKp4vNM2ICagjCZIGZNqO+dF0HpGRa5oKplCVDP1FHMC8ULtplUa0t8
w2rK7Z1c0tQKl39W0e0SHalE9LEZCNqghkKKFz9JnDNFvNgcm4V3SBsnSGG5SOGW
ViFxENSB/JTlvkInWkCJ8EHeVQyX/nIB5xt0zfxE4OYuCQZ7sUybaHh/e4wstUud
tFhHYPCZ0xVsVSGDgFDUfrGBBLPTwR/kpX9lMN7gzueiSddwKUuamRc7FIxmth2o
7bmut7XlFQSLzS+7DDQo2rDFc4HG66O3cDTCweu8VXibPIy8terfXNHR5TcIuYEA
qbQeJELz2dbCu9BRy25A+6AxTNJdypUs6PWvdOn3iltmy9/IuAuXyGX9GKSU04a/
YpXuvLMFa6ZTR8v/KqF/ytXmE79Rb5/PintlvqR+W/lwhs/54Tcj5P95rYvQRXWX
Q9u+5ZGm/+SfVn6JlCBag8jukVfwcpEvnJHHr2eVFYB71+xC8fE9vwE7WvfqRcaK
tsKLJzFTpHcfcHranI35XgoXIu8swdSJ6bO7Z7tAwVsbIZka1PuYgJ8kmXHMGpGF
19tWBbvwxEqccAaABqyYcKBojCJ5FSXtrnKN+2L00SFRok46Du1N7BX5f2zK22Zu
5LOBUGOzn5HZXJf1RzrfdWhOwTOvjdR0gmulR8V2jwgXIbLQyFX+edMnl4LWzDgt
yJHIozkD5wd22K45s62TfYz8HUfG2mMdOsD4fVpfEfJQJjyi/v+S8xuE6daROf2b
GIdmqRk/o73lPUAMKVX2XorK0UMFwmLOzck6fc8YiXrecm8Lvt9y57IkYdaxkKmL
eGk0Bkc4NiKJrxjzToBePu8de9x+Cv81OzZYy/JH1K1ksTp0HwtrPMfhExb2AA9b
rIDLkIILPoUD5cb3l/Bt4QF/8dBcYgo0kHbgXUDTeYhZ+nkN8TZx3i3dqprFJo5W
ARvkKQ4CpmPDU1NTNR2eR9FT/yvLc/2JKBqs3TuD3M0lONpTAQuMbF9eLOSwQzSM
dI52j/UdJ+05MedgHOPFk4yGzE7yvKkEu9yvC/53ngnoZVDVXVlRDDThg6yQoT++
GaQxZxt0A3g7mwqHxH4k24MkMnoI83T2M9YItXPC88imGW3yK9KCuzuISYn7lFEK
tv1W53Qqf2SmxR8Hpa9ZzZiX3BauuU0p0UpX7e440EJ1sJdwzQqviBHHO8AJh8oq
AJW9DUQqoSDg7q43TcdB33ur6K9mEd9GNfTDp6NsGafHeAw5ILKAHnZu9Ii4TJMl
z/cJCvqwxrdwj2cz/pFNqN3md6UYwbpx4Uk8+8K8CxpCYlQG46c0u+koKQ9+oVG6
AbjCnKyfLvfbQK84YWb8JDKchWGb8ajoRbA2SXxtQZwYm15IgG0ouNVAxpOhh166
PtjBuh9ojGrN9Veph2S/dw78RM91Hl65dy7rz4AnUx/c3G65olNvNadrXorcf4X6
GVARXyCwHFtYsBbuj15BIZqmGq2JsdfhydDeRRVahtQKJU9i03nzDVY+qdXQleMz
ULJWGPYJ7sR8QAaQKTYNC+Ks+6B2lXzW4qLpqys/5mHyGHm6DyMj++uUmml4nTPU
EBQOpu5nPYTm+zHL35EwzV+epIvNIXAk1fYe8CqVmUySA5p6sfVvDag+y3A+sWQy
ozepV1VkFd/i/hX0S+fj7qXQF843GmZPZhHcDa4MLhoOolPkFA2GM+qN3Yf+J0GK
VTODjAUjl2LGVq5fl9TR9mImb9jrw7YEPmixfzQuDGF5BELdYtArfHbyPu6Jm4N5
PzfHqTEUaTKXXqIRyUygn8mfNCLjI4SUZnqK1D6iCmLgMQkYM78KlPq6QWXqXizl
GTTKX5E9OuqxKY0nLuIiGuSo6GJADpoXzyRvn28I6nLrqVMFsu4PFpmmxQ3ssHZq
8mvHrpmVfcvVSfas6489+Urs5+DOzcONtNDCGMYK4N+bL7+rwmOjnivP7K0TDXJ5
6CbC+cKed0OG09aLxxmNTHQXuRf12Rhbo/yd9qMRthQ3Q6l7w4fRHAoT/NIgzbdx
Iz2lUvAxCixdRU9oiVbcFzYqn00ZdijekZ2+QO2xxpvMTVmP3btWGATAEMWd3VFe
qrqDBjNc+J6TvElSmUKTwINeq9dPVA3jd4oPGPY3PH9g9TVCP7koqCFZMlKzwFFC
AImR91rzvI0NQ4E1ZHpUxgRDUOis3QkmwLewEOn//YbEO3LLD3zSJqvVzEJeTOR6
l/Z1FqwJc9z+TYFlu5lDB3ydPoqa/OeFn19rmWl3inqlX/d9Bgout0FxBiG0glpE
ItjYaKR3x+OStRar4Gzn7TSFitZEQJ86p32wZdtN2Nqb5Bbw/OACrxwHn/OSMq4e
Q/VGLiG21KjXOUDc0lLyJfyE0MC7+sQGkI0cKS9lVvIl1rtsDxzOlfJVycupByzr
RX8RJGWrH5FiDSnw/9Lm4OspINht/NKLTAtN6aTdp/+qhVvfuxZmRf61/wwmX4hA
rrg18MSLUDg/JYRCr8a5uqoIjV71gsvrw/jyF/B7RJPnB/b2lCKLz6NQ4g4gTzvE
XjIP6oI4ZjnB7VORwbUMYxC22M0Q/qBOY/45AxinxeONMCjRj/+f7OLDICwmgXVT
YYAvfas1lH/BpPVhE9e9OpRGAejULvd/ou9gZZU1TyJntZjwOs90o7uHr/2M1Jj1
nMzHiD40P1uZ3MectqAZtq4Nir5y/bQPAcQBjcPBdhSwjHEiFFE8XsuMGWhUjqpv
DWJ3qOcHzX4Pu35j+6UwrmWlo2F4CQ3CKnjpOCOkOmc7LF+SfyDUeG5XnZRimS0E
8ew7OkY1VrkPYO0XNC9XwfNnJHrGnKQXZfOYzz1MZ38QHctSqN7IoS1T7xWvJ9iy
TUcT175JIhb5ijRxr9jCd8qqz822yUz3rpk56QwAwMio8TmN3ZrkknAQtQuAa1Sl
f8c+iZHmDvHrMOF024JOa6TUCcg9S50X5u/fOUgdh/xSvysoL16fQLS/gb8cxKRa
Q0DAP6DtE+yy/uU1eJDKu0+SdNGwAxRPbZbTbqw98SwB7ZT4sxEqOoQdKy1C3NMm
3I6L2ARrgWaeIwCH0lMYIBxHyKxKudy9W5gulHaBnGO2Zg8D+Q8TRNZaxSX6ljQ3
hcUeF+WIfTw29rMIBoCmJScdq+fqdcb5Yil1r4jkxJ+sMDfQvzaQy6g35in10pIN
azzCc/3IzeFkRNt6Ngoqdl3TinzVFZlnTEnM4rr3xcl2UuLRT1wAsZMX2e0C6xtP
S4QlKkD/NE41rscn3lx7YLEKY1zOiVi8mOnCXW+DW4oJLBcOsV7snh+zn8pQYb/F
1zFnhkfTKq2X4mX/QXY9HorSXCPcPFgWAbU5KPGxyUTrvG6tHxQd0Ts/xSqhXGv1
NlNbhQuDmuoo5rKMKne62oXDGs8g6K7UUtgZbJ4xAW55cuUTZ360EDnUaWYLklde
HX8JeSfJZfhX5cDJgcWwjrYrwYNDlHBmOkNtheJuk0gcQxraUGjT/jGW5zsLzBId
bpkE7/76FuCrLnL0lZhd2BkWe2RJkGMe2+Y1XhgYYWYkU37urXsI+Pcflv/n1JBX
PWVnhhjvjMNeo81hnjeqsrPN6f6td+DkM+bKN7F4ZM3bRTDjpTpmBUYri0kgQhLQ
TzW5SDn7fA7CYL5TRlLDicuWh0IRybOWJDAozK511JaE4VDqZZREV6qSI3o09M5b
AFfVzgEMqoJJHFZsqimAHv9F/sYS15QDQ/l54yPt+zkyXC+B2ZQZ5T45xzkyJKUy
RM9HasmF+DNL64PE3vaiCYRbQRZES4Xvyq2w6wyOSD+wLOMR1rtBwZvx93q6Ma9j
cC5ELYYCn33d5OlOWeaVjJuXS/l1DkTbdIzTDXZJO8mtC0EmfKIb3na0nqfRQZbj
WWzUsDNDJCUokSbAndTuaGI/cSpyZ9wi6Gp21ikKS7ZX7KBKNuf58VWd5dsNxm8q
Q7wT5gDzJTKmRi69q180ZDihF7vCrNtJxU7Q2wh79JyPUeUN/dvnsUOWBGvTqmYs
xrdbXG34le5AoLdA0VBQA3EnUyL35NkYWdPh1d0sjh4J53FrSTdvVLgUr2UeYoCw
kwyFMwI5G/d4cENFqWRUqyaFXvanE0VVbJZ1i9yCxYFDwvGHQXEmA+iSyCUvjZKm
FEF+vBrLeOMYJPcqBt/rBFTRf3+9I13EOWtjyZNTn2xlwAAp9C4UvqYl9KDh8hfQ
cfMVdCET7pmQ8WhWZl5qpH1KhQnZWpa/tGC5pllhr+SODhoGD+fL5pkmgNlTs+Of
oGEXe+vxjcjVtedBJL2TuHowDUz1q+oEk51itCRRIsuGuSgRqk4bFgt6YLMTE4Rb
eY97I6UP7k57GIr15bhzxorrbGSyGOPzJ+SPbsRSL9OorjQbhl0uNyx8aL8GackS
qU3xx1kFXvmniP1riGoQzFoV9BDRoyfVrLX5DRAKRJJBmZ4V4owokUHdIQ9ZTb4f
e+j5pj1KCRdQEOYMUuREigSJJLI8vdtWWFUklimWRUBU7SVu4mVqIMm2ijflEob2
I557gAdMbkFHWldVHkAmvw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
MFnENI3YEohd4L1CXMkSxxjOREwjJw9lGwXFOXW7pKnS6NBlb3gf3OhGxn3vzseU
TBi1TdlySYTq7HIeUZ5EaUpBaAzJOZQa0CY0BP0hDo0X7I6uXeYHWFWhKgyLtoSp
yI4e5VGYMzNuhpq8fT0meKaMXkl0ktjyGZp+B2kioUb85IPe8h7tFWDXGzzzi/OG
Ijk6h4JEH7uISYzOGzbyUCkknuD2AOJrMXXR7XnWyF+jjPgrw5gPRlbOHmdg9oTl
k7Vuvfjw6jj5kMm9c7uueI8Q74x08W7sZA2Zn1LZRPHwxyOXnvUO0fLyf0RhuB3M
Ushp+/Lx6Pxxga4GmQdsPw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2864 )
`pragma protect data_block
NI/vwzSR53wGa4MUBOxLBgQ4Vlc0gsHmaefg1EA50TrzR8cdOjefiNAyeFx8UjkB
6vs7k20S1nsnSPXLJOkp5/L4quqh6uR9Uti7Q+V3rqYgSITfakqG+sag/UGJDOUU
tI+7l4Z7ND+oCN4aUfMer61qwg8Ot06Jc5O8pUMvQm/OUfw3yo+DDlZqcRcbedGW
wKLb68X7j0FamhHdtOwtPaN5r1CU39iiiBRZD4cIbfOBSZRNYEYhBVWyGKJ6B6+n
MYTHrl3CMa1iFLNTdA2aIwF1EkkBZHtlUwqEGNSy69ByOalO6WVNohBTpv1F7SGg
YDcagWtddMEmseANEI7lyGZYg+btggcfo4G00/hY6WVG4Vw7hLvzdZEA9NmbMGDj
JrpGQ0dhNMwLSx6Dv/D/ijW8C4Edmq1R0JPdtosfV2C9AY4j7SGaXPXZUi7LqiEe
KwXmRDqk9tSYTh4lYsvC6eru0dw9Kyc+RQaqZXw4Tg2O+hoF1bYqIU0U5rpEGVqG
HbF5SWYlR3a1zQ3i+OZnhhBPVYBxtPzp5oXF6FBXhW8NFFJDTLL9pCgeQUNol3cb
QiLnggn8EAgChF/hl7uP3n/c+yFsxoFdagyzE5s6UIjcao7jtgZkokauiUONjhNz
xrmWscSgSk4E2ZUcfsk2EMeRb0ZmKttSaLxyBOVVQTsESLeVF3YdFvkilbSIfZYb
XkeIJ4wVZ+pTchI6k9RuLIyogPU+e9miQGKbr12U36kWL6IQLUT/QyDCq4HT76QN
aGPuCvSl0H7jdNKQ7rD3BkkpnsiZKf+quUbkWAIYkuvx1sFfCq8OX3t6u8XEaIup
0aFsqsShCxi7vqj82bEXeWiGY6rQCTKUeenrgwgrLc3UfPi/oiCZakRIKoauV4b0
RNAqLGpjFYMmnjpdpu+h9wCv89DDbrKq0dFBxo71o6ePtCeqrjdQ5k/nNDDc7rpX
ERgz++AWXXvFlieeS8KFkvtfmGa+QjgMDlEU5mqQDLjSrVsHbbGNLTsDlNdcl//e
s0+PfcHvdOvguVN6U+DPS3Da9Nvqo4HBJI4t+4ZTZDis5Vr6IfP0L3GBCfmBmkgR
t7bKxlqXHWHIPnRaD00O5SQSpKbg0PEYxT01I0eM2o/9z51fOJAxoojFqHKQ8fKF
O7s8Iz31itSzPd+mE5dAL0w6RZlCVNBf7rVc3sSQxOvjWXk0/XQJx4tiSEzcUfFq
dJCVoEqOpw1FTPVQgPAXcxu+viBHAhNGyswWdUopRx2G3pjSwz3WopLjZutYMayK
MrKN96r4gNZ89+JjQ0Qib7sLwfx8XI3fPa/Q/XYevlkjL2zm/RU94JJEjwdqwdch
rnmNnHbIYWweIW902JZ8//dEtxC3hJGokecXDg5i4Vvkxrv5CKvaMlDwULo9GRVn
iRyiDqjgFOZJjn+jDAvrzg78dRLU0X10J7jev5c3fD1qxNvFKycZ4z8Y4u5c9c2P
gWvku+9XVADbBnM6cV1zJkhDkXFwEyp3rf9xL4hhPFf9B0SlSqcAGZeJtjTJO52E
SAbDujb8wYI0xZPQfCYX8/tcBqZ+Le6SlNSq63o7DMr6Sm79Kz5cUcgedxvEXXjl
S5egAzf5oYI1V4uGqif7lBu+0FIToujCxnyfnIgRqIx/Y52cseecRR8Mz5uXciYh
bmVjO/rvQpX/ta4pMovdw/nFmQrU54rlQJDeuxmlx3x9fEGtLkrA2o6lBd1fRx5r
cN0GXZNElMDodY1RFNMtoEwtj+XWrzHc4m00/bAlAjwns7lGM1gZgfl2vQKsplvr
Q9TticitOtd7LNlg3WLfzhYAkouAUA9gxlCXeFVNAgnYBbc80DgIwh9XUb6HvD+h
k3spcgG6Ea+13wa0vYlq3WeGELMLT32a2cYNjrkJjKTBn6YLxwIRUO7yUyy04+h0
C4l4EK02r7usfTHxbjsJ9Jdgx4nkK5WSY76bpyusUj6zkVcJu8ZbIRcVlVdhfgrD
2LLymsFpY4UH+dfiZwhoFnv5uLq2fnE5NUxcgpw0V0ndO4UdWn13sazWeGvPRd8P
9zWh4uUUe/yE+mISFWGrvCknRzVk53vMXQK4JyNOkngEn1/sRaRF8r8UQrdjrz8Z
+UgNAY/iCuJLdyZFR+pHXcFmdFhQBidaUti8Rclv4dsE5yc7TCZyX7ywQzkAvbeX
niA/m/fNsisv9vrfjijkbOl6byPVPSj5BEilYpNtkDi4MoZhSC3ImZ3pznnqLFRZ
kXZexL2JGfI/3FM5uHsQrG3ue4FlQgpMH0gyxTr31U0R2aQWTicEtLkPNE/Bn3aO
XYkfJXm23NBiwM/gcx9ckRg1fNF8TTUhjH+LrQ+OOI5DbWXIXDj5LjAIuZjjzHde
ZkzgGZ+s0yRs4s2NQczHCvxDobzlXqBPahhTum/+rkrLrLL7Es5F5YwgWNMl5Nw4
F97xmNkWnBSOTnQxR3ZRHYna7GUUvB3q2izANxfgu8GlFoYio2AefxpUgciFwxXn
vusJZIq8PQ7L/yzSXmphJmjHzeA0lgur77IoXhRJZ8uV5flMNMx6ehrDcfH8WhzK
MFqwLyMPyBguWMYctnmLJG1B7QC8w5LlccHX+eBomUtYco2nc9foBSNuusZLVdjh
7eKjAPQrQVKexyXXotJMsWCs7oyk4rngHXNEeKsVH542mklVru8UlgtjFQZaMGS7
RXCUCBGRisxOKchnOuQ5KHjh53H7T/PhVLxtWlkhhNiGrAullMuK6/y1M4Vx9MaI
cUjTvvrm3b9ln5KAv6GmMt6Dj1Hs5GhqY3x+0evnanAX8tAAZqIGUamA7iwgarUJ
a86IqJAj0swucY1XSUEUg6NF/2PQ94/6zGE8uD/nJzpPsQqNdhzUlAZDEewXLRJA
6MDQ/C7EfmI4KO5s7ZvMqZBWcld8G/wVwcWcuEf1t4ro1rlrFHFZg3B0ixrnr6ha
PrtIGn1IGsaPlRNqxOiiFF6KYlJQXvfRO55iieuWSOjh3DU0ikL2WFocI0kgyfJX
K+bJg29jOzVvi8ZUFE1Ky8CK0fDREQcK+nFtW+RUy2f1M6GHGxPJULaoW0AToJyo
s7jOov/K4Zz7D1Sj5911JbB+FH5i+xbxXHnN0k6fbs8tKnyZqPQkaPr817mEHOP/
y6zmJZr+CfmLpFHZpQMtLtiM3m+6r7/kJElnuI4+LABPVXYK5cK848K6mfeNrsQ3
4vwpgpwQgHTlWzDrxsl63YuIsHExkRMxAzqsqIIlwDtSdDlm9//+b096ULznui3Q
jrxQSdWbRrHzw6Wy95/GmPs9+jwHnATN3YURBAJqt9wyZ7WkdOPbn3I3lgLHhBXw
Td1nn2O8UUBQ60kg1/aR4co7cfjJoCa/uO2oFqXKIIOlySa5lMOz00xZpc83rp57
4QmbE0WmIyhBCyCEYFXDfFM4qHMNfFFET3NVEL6+JvwsnTGj/B11wvNXbsXuGpAK
CLneJnbSq4cwULkNE11DLW1TDl9ZPOxgQpyHVtTPhicHYtl3vZss0jaKQzpIXxj4
YFe6x+ofyFs/q6ojIiU+BovBqr6bBxlAhuvgi3ynuaNxh025f/VbbOH8OGcBO+qv
f5XfVVfsRTdAKzKtwnP5RoDGk00T0y350OSCVxOypxDfy5I581I5UHnvMJKIkUS9
G3cLVS3ekiItnSZvdHqKs3NX/JmPmH+NCazcVgM0nLSwfj6NsZyfsvRI62hMaCNN
lHQwSLgqJL8cYrXeqktHO+mjmSMrFCQfMhHOWKhHAL5oz1qovuY/ldWgBKJKjGl8
0UTr2f50k/lbGlEQ/IIw+EBlifQj0fWHjyKc43/Q+WU=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dc27KO3yYG6ls9noKufyA8Ckuw4WO2at2tMzzdLNyyMYCqVTcfpCrhYC3TsEJtBW
FsUHNzUPmSrgTiQpknLWuvDBV5uOH9iWN4LW3gkuTrg2vJhnzdH5ai58hNg1VkFk
9xHwJQllYmYig9PNnRISEo4PDnPeosTEKLR/7y4C/VbnxzP9MUabaEUNWLBe6SAn
3QDye6mU1X41UCvStM1UwIuGpXyJMm2ru+BGznAxbYDqtmgW0OATPZv40O+f5Q7i
nfMSUDAV0OZLODywhZ4VDxfEvr+Hp7uBpSs7R5EGqrrxsIuSYwZcf/xGvjAqQ7oT
vABCc1Y8ArIaRjx7V9vGRQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8720 )
`pragma protect data_block
qSUY6cBtxD6WtsNHVuXvcKVCx+3uHVIqirhyzUDd+beVTrhr7GgDaPCS9mPPLeQE
fTXM7aNJKq9skp/FsiDtUuijPMpFc1Jz/mlFCKWj0CFlp3M3dHXAAETNxDVPpwXH
wbT5tXCLax3d8plUlXNzxWFSG7Z8cMtJhgS4tCgZ5noEG8AS418R4RHpNCcPfFq9
1CErwU9m5MwSBdJJpItk0o060rgEpa0dxeHQajphMVSoIN12AIh9/3nmCZTcktCc
bGAfxTvBSUxRCxzvuvyVUgf8ec3Ir/PqE2qqiVNQQe15ImIjRf4IQY61Nua/vue5
IYgy4ivBHDhmW5VjqEUqConVypJC7PpNcOjU0/yOR8lyno4iVhoyjXvuaG6nydXU
vx1NDXbFkSnnC2Mzbzvah/uJfY2DHBOZvkQoBESazjp7J4LWmYbt6FBHwdh5GqdT
zDdbnp+LOubG4Y0f3YT+a9pPZ8cFCD2R5D3gLMcPruruZ0ZR9zIBdTzThAqQWHlk
RFGJD0h8MmnKTtojl0c1u3u1J0ZbxKnCpdsL9yjvfmztm80l1ikZ9+M6RGtGHLQ+
wPHqHmkMqMw0sTLdV29yE9hTP4MwL9+1ZS0xuEuKqxWNbIddVdeRmYKkfIAWTCUk
WqCvtzwDytxy/w4Al34JhOFQyuW4BKMV1ZSuKytDUuffVGen2cM1d2razMQvwhaH
ArklfWY5f6v1v1B4Etf5u6QZ0e7wzQwu1IIV2HNLMBcWp4TdMKuRjwm7jKbqp9Fu
0mm+3u1tFfnSkv6TAU5vS40XdEDpwil6FjHxZg3CI0pq9M2cPmbdc9rYFwXZ8ztr
JUKh8Sartl/vwiHLd6O1VasH4L10BVPR7u0bVcg+A1lDws7f9fQVk2v7tNOveaKi
//IUF/uljEZFfQ4fa+csysoDbdy0jCFkVXoOZIC6k4QL1C63x9cLWIyFz/D0ws6S
FulKC56l1FVm25mxFxhuyWE4gSKbhdxx3M1JXgIgaGzFxqlr2Qj4ncE8pgPwSSM0
GJf26b3Oyno5uFYHFRRuo/2NOF9QnwChVHcj1d+0VNLxU8eBM9yB39owEA/whAH+
2fANNgOc2s3NSjVhZcRkA6Z0KA/A398+RIi5GrxQnlHPPJXmSDTTew9enWlUMB9Z
8U5x3IaFZPIoAcD6Ul6P3+qtMH0vYoD/q7dKfx1Au5ew7dtiHfa2fwkbdU7du7ho
eed4bAHo7ckAcUEchKNHUvKgIi6FM6KKVjK2ecu6ino1VWm3uePO/7xOgNXg//Qw
xsGQRN9MRnBOTiHtillmQak8X9jWPRhnjRYXkjhpWbLxTHCoMjxJkxUxrOtvRy0F
CC6KaxdFYosJYmC2jbHmGHVFA4YJq4rbjnb1ZP6pa5eKIUzR1Bg28MbEAbJ5UOfO
JGU2wX+Dg8EXd52KO/iHcyopIRba930E5OrXMRdR5rxwWxI5tzo4bkwqaJeXocn/
vadQkFVf9IMeSujlvsuZkrWucWk352nspeNFBx/bPO+5/cyZYIR4CXJ9gfnmJIK6
en/QKAN/P9pyL8ZyRBH95gzQgJdIvtlZO85RpP3r989PrOJ0hAu9DZcCYBUJ56nb
DAGkKQjg8EQSuM+n/2W2n5Wz16A4CYoBG7zZycai3PP4XJeANZ5kFM2lwhz/CzH4
MpSwe6QuGfGFSBfytpJGeq0QKsg5yB0fr2iandVWFdm1cbIVu1Lk+oXbzjmlEcDz
rNrgxobsbllFQ5Cr2kXk6hlzXPoV1IIAN20iVA+RlLPlKBuTYpSQbD28TnvxdxoD
aHtx0+aMnroGsL2ksGs0WCnAw19Yy9j48kpblhflywCcTVo8TzCnyr8kOaUGdbiQ
rwqQkWvdSXNSW6fnFKtcUqArxmhLcfYG/K/PjJU2PkT7aeBrNWDU+zTlgfnnJqLg
Pa5HbaVl/WEc+1L8YYxWnvapBzOwmsK+MoHJ6Pwd8smrsTHApN0tj0DoWXrSCPLc
5bOVXKfRuBez0mSYlixh1HXv3aO5orsjl2AYEPje1QgpwIVlRYxu85DejP3Ybkcc
dauVOsRqyYeJ2opu+yNkgJsmlBTHpuTzEgsm8dYkGl6KRTKE1Cr2NbINvTKqSiaX
r8m6026cMJsAp6VQ7BW5CP6pwfeyMak6alMRA+lmGgXoOA7XJzEftSOQedpyaXpE
SnFrJu82OdfIv4qODBfPsqueUYfhixP4UJN+5cEpKW4k3edwPRPu3z6mxskBAUZS
p7wIyMZnoIsZtgNxyYfVWG+Gy4h+lAppuex4tFKzAt++WCV96AEbui4jKDPkVidy
bBLAnXEtmX4JXOSxAvlL9bRQiwqXVF4gkAlLqee+qaku4hK58gI8apRTUxEftT5y
Axl+wPclEbvUzav5Z8Q52FTi87UAjxRNRnIAvBiuPT6k2aCLMXAFi4ObmdtBxhSu
NTqzi/rBobyBvhyz2Zat/UCwlKzyGhmDXfsXA6aYQSw0Uq7kJP04SFrx/Qs9gMNu
ByOCcIQWyB2oRIa8eUytXphXA+ODFF4zIl00iuDZjaA2vzulEohmHrwoCJxRxABB
4K/Zfc8HxcgDOzpsWrIb1Ker/Hv+Wsjw8tfmM/YNucixGKOKIWWEbMHlo73qRnRU
iP4oGvkyQMc/mFz44rDsN6OmaIl6Dc3JQbpOXUu/7iN8gJmbrS3/woy28gzjE7TS
dIMsmQwmKhHAW99ZoAjCMN4VAo0J8tAGICP7LiQJiaJIJZZiKi3S7QkfAScs6UuW
/EdxjoJSun24MfthNq38k8rPyf2TGDFTeCKBG6mPlHkdMQpJP5gkwNa+WZ06eS72
WkKj4pPvOpDB01sRHDGg+fxpOacutWdJIFLnfZFV/Tcck7wcOOhYaZXAPNAocy/m
xMC6wlQMlo/P4bCfegAtjgxXQ27EZ+otbcfVzORDfWQ7gEEEQluRXcN7I9QiKBSR
orykg9VrJSLiKvFMVNsE6t/bR91/PzVWc74v/VdNuyeij96HrswdsWUXO70A3aHX
PdsV/Ca4Te8QNFZlZ5gQTaz+3osCGgzJfSj55ytivKgKp7+M8n4rbRoiM/o+MX8b
aQtG8AMjR4B79fbgCPzBIjfI2QR4n7t+kEWlIs8w42NDh0Bje8QF22iEiCpZjIVo
zk97Tc7ryqwbrokYr2JmF2lEnccrlvrGSEPSuTGANihex8VgMpSasIp42qrpWiWB
7FptUiefroVapFnIldmOxcyeWTrk5LbhylrdlOSqwyBwGiqCmoROFjYRATpPQeEj
bi6GS9pMLo6ZCWm1AhNhyom6GldcMdXPtbPYSuJ4DfHdCYTW24xqkbQgsHA+VUXI
qIirQNvPBuMoJe+aZLJwxfJ+Svnl3FZxlgieQmW0FJgKzfapRxKq3VF5PdodQsMN
w6RSTKVDxSmNVUY3IevNJKnFqD9vbykKqKCdkZ7atGSjkJjyScelA8fbWDMwellE
0wdI7UnPC+fUnCeHryeNd81rmIFQXMDNQ+hKSRptYLNIN12e7Y6EQkgEx4qwptJv
DiGx8aWenq1TRaBfemvfmdieMXOeI525mAPHOUeB1pt2ykgnNaRdC2Gs/trxOLVL
68l7Brj/0pR/9IQjJ70BwLt2bu4ubAsscj4GxLXw57mk8Zo/lqZACLa4ZY1izR7i
LT5VC4U9CMzYzxRW4tgVVbVYIMGdOFq/zbAU67rFQps1XqHpaSk6o+jLVoZ0Y+AX
2/7iDQvs2kp2GzYP/SqgN49dzEN5+I9kDEyC6SxhOBzvOLOs4BTR6jarwAanMzWR
TbSKrOUxLkqu5T/px4qEuvJdwbXVc20tA8pkusHNx1sXoIcXTcETFO0niJlZMTS+
vFMEOypXcmXwoSywqz6lDcCo00qyaVTppmxphAhuzpM2PUfw3CXOYn/l1sZpFnFl
cDG5N0il//NL345/+7OCxzuHgYW8gEhOZqfKy0mqTTaE95FKbLTbXg0LHgComqeH
U3Z8oQbReGfWWU0hrygmO1eBbuJc8mrfVcw3kPodlyL8LhvR3IewNdeSWWUsyK62
I3uXJUNHKcJS8tlcy/MUZbRakf2nNpsXazbpVNeXmf1mcNiSvzJSMMjey0zAVuRq
Ubx/9JJkr0VMzcujBEUbFI9BvnaZIpjhoTn5NOsg72kserjrZeewScn/cyyKDNUN
JTg+z6HnBXvNthzpGYrWWWO+j1OG+FtIv1nWIHXSeVO8TwXwDYMC7k7y7IA4HK74
ICcPImqG4ugYOmzUrPxTVv8w+Vqe8Sq8qJukIDiPNn7RqWB9SAY4ZIvjoOXKpOMT
Zq730fDHee1Adv+JIYA8STMoQuNdoJ+E524JhvJio/h84v+UcEtBblSMtus+6sD/
M30VB1z5Z25DK9F0Vh3GqduT2LATKW9AMECapB95rz0BNDA4gjWQe9DumkWlXBLC
m4ldWxEmeH9q0CVi1nBdBd/23Xh7jGrFgLRl6U4HF/eWSZa6GxFA1WxxlhC1LzL6
sFjVpcS1w1jCdS4gK3dXiaHkjXHNzu5/9lFhT1yk1xC28W9A14ELYzhIFcIe82lM
nQkoXwSp/AqEYK3gKtidhRhkxZr3438zaE4GSRmZcaaIQqyg1/j/c5k+Kuj0WzGT
qJ+O6yeMU+mp7+bFq/DRtbO8VttoXSEFc6ztAtPowtd2jtH1XhyUz/cNzie0jAlb
zWEgq+6xu/IsMDITGql8bG9gMQ0u8h6ezqRjagTxEw+q88CLX4zbQd1AKufVcRmW
G1A5TJvNvak//DjatttvQZAaryqraL5Z84fq+Ak8zwJwtnKQ9tth/slsu35PQpgL
Y1cSaS2Jx22R/c34afnJz7AH5nGNXPSsKnYXYeq8ZVtU2AzhPLv401SogOo8OkT7
TOhdpyyDQEwGpZ0i5vNx9X3CC1tj6oHk2XYJdTrsLQgVqVqVyKq0cOZgs70cYSYc
iG0e4ZBc+Fa8FfbqiG+bVJox0+ghLZJl3dnz5Vzt6qIN2oPweqBEg20gYcQEWWg/
v73aVW/i5A0YI8y1UDphF0bj7z8ORifY6WIAdahO8RXVJcv9hnCbZw58B6aumG6L
xxlUphU9Cz7UdwC43WVq23qn20BFNSLyieXPrSt3rxrK0g2j7ODRYSXzBxJjuM7E
hEbGj7AANO4vSzw28bK9tMzVB8rK7hYMjAEuhE9PUn1DqWf9Si0NPbFo0T/UKp/l
ot55y2ed2ocezm/JHi0+EbCd0a6AmbXgT4JhCZRj94mhNql3YGW761MqWTZBKp1k
vxizs4E47IbwEn5bc/pfvzDCz0XtbFNEbK6ldZgNtwlYV12rZ9eESvMK2FHnkzTM
vIxh2rWnQrQqUdECXt+NVUeNKDhnVJypbQNVZZ1fIcxN9/MEc22M6YSGUSzpe+P5
lp9wxmV9FDum8Z+W8Qx4GtCtC4YO3GIwp3tfzj85VQ2vVMxF7oTOljkzzVD6taMf
d51u7bvkEgnzzk0xGDTgIM3eLR0skj011ZlAmglp5zA5MJwx3MQS4jzhYzSks/re
a7SgLjiZLp2TggUPFduFoHlmybbFbTQb+lGAYEWI8p6GNrxZRpc9AVm50nIRbrG/
WCxSdGXwkw86Pj0PwCC2mi2q9mfFO8L0Jt/hzNE8UTJyngsVNGnubNyRSRDF52LL
h1kuU9J4oFtdoEQDiCCeksMw3fgfNHr1KOVdUv5YFR3mneSZas/XbY9RHH6MdHwr
btLhQq+8RVViRiJoKUhSfBxROtUlxRfMgb65nfv8Aj0ZW/AEea9ngyIIW1tU7hri
KIYIMB3WtvYS/1tSpwgE5getm4lv0+W4mMoazk0+RoqpzIwkvrSlVHMZgsihWi4P
z0gm75FPUnA0Y5g2jDCP0iPYgwiVOoD2QoC/IwhU90or095zs0tEAUBFSQNA7RqH
gEQtskEXQlm0/QzEHkt+nLe58Xm+Df554F3K9BY0tjyO7fXEEphlA2tasYocYFQE
/T8uheA3BOWcM4e+9EC1+FK7BgxXutbpIvm1vfiXFisjeq2ojMlPqWWf7uzKYr5C
IXujoEgwYzjBFV1NRlPpoG6/14wJh43V1Lyf54TJOG3HEoj5oWrplwAkutKB9yn3
s9pNvhfRzPURS7eadtDQroF+vXSR30yEyoP8suG3QmrLMF4WFrcGtYlCkQ5iThCH
89mX6dB073ePhvPnftEVwNax6b7yjjiOOjk5lFuq39cscz3cAVrqjAQM9Y3myPbW
yaRv4XFFtP8C/O88QX/yxnSYhceKvupuHGDo/L5WG4cfZaRv58FZETjkSOnfSLIF
h03OeMbSgGr8k6gQxRdaAM1r/2voh+ZI/YdcRHz212+xTnFsv0o7JJn4J+LcXp+4
IXL2Vn3hLmphErbfzMa8DNCCXLT2onjPU/G8DUCLKoCDvZAckhg+hKKNDzMQMQQE
sgYPce/LBkSUY8/Ikh+wTf+IakPeFzo+mmhJE1X+eTXG6aL/8O6F4gwc5w6cSll6
36x1EGQjrXeLGnaV0Tr4bbnQoO9FBa9exk4bYhz9w7TMHJ0CnJt0kEInxqSJzpMX
lfWHkcOtgE4XXLZ1fSQ1CuL6JQfBnut/XBI66OCL5JTEUTuDjOjusfMTNzgVJfzz
WHyjL4f8X/TaPO5kAvlt2nS8oVwf7NC9IMiNeVhllr+mZnOGx30Avc11eYOsexue
RFfwv/D1zvb8pHYA8ShHyGcVLxyqbg3/KkprJm/b4XC7L5RSZxxM8IlXAfdh0Ph0
4leLiZVoX59stKuJgWpFep0BqP3fPwtXNnqLki/D6/4xm5C0kShlzCbIVMiyKaEG
ZS5+u13oZ3yTNK7ULdVbaEmkwas8O5NDrZ3wjrWBwAK/HuEGoghYpE0jIY5ow4M+
mq52icOANfw7We/c54qKhzXDQkRrv7PncDXsYVptnRJCnNRQ0qROqGTF0p6QxhVs
oj0tcdK5NR+IEyOKKzv9p90+F0np7JrZDLdlH3XHHzKx874q4zrIsmZ+8kcwniwk
IEfGYO/pmwuAMyWyhDeRTwgtDkZmcXqTkuw4e6vD3R1OmAIKUNHQFSgSKcsJNnpA
M8QYN2C+7Cpg1CnfxOuGKoh5GLJ2TsUUhV1HJS9bvxEHvgl+kEUJoUObNPNmGZok
fYF1XUy8grlJlvxnX3t2jF3LxvbK0sCn2FtGUAhLKrD+FWBv6BkTfYPM/56+MAi9
LLoQ+cfbyx61XAH+sOQ3oDjYZ3V2mA2hBe8ZOBchk1dcR8yvkeud8cRQm6YCGLCO
glFbqbEQwE3t8tDciLbTDHAzXzoJQEtGXcvm6PLeROWT5MLYUioN5IpgdgL4c6Cq
/YZppT/OU+8s/dH7s+Vmtg9yD4RSTSVO3ZEOguJUWpcXG4bkVOWpwECPV368Nbn/
2bzCtzmYbukcSEXUErae3deMY06lDA7jA4vpkWQ5KZUOYrV85V2rMfYMYFHON2JD
YQYDu5B3OWHAHRF/m/6vnBApbecZz4MfB3ukyuEM4zp8JFFlmKFMBx50H6X3lFMW
oS/BWYXYTaRfWWszKovdeeAKm1wE5nVDszgu10s77CmfQpMHav0DYc3VsRB6EwOT
hitubVyeRZ9TQ9sRnFyVwkvyIuSak8ml9gmQt/FtvaQ/fQHFfK0LpBaKJYl8nIAC
1y1kyzGvpwZRSi9tlLz/nc5SZle4D+MFuCEOrqJk8bSkuXteBvhRcLVVzpBdZZB8
hA22HlnNEZdG7rclYyy+gZypZE5Xmt2aUB83doqF1wuhhPkX1HZaLlSxiLkjMUu7
/y/GZvw9xt10m49FuWRJutG2wqlZNIbpL+gswZndKw+9MdFyT+fnF3ckXtW846db
RzOTBE6uHfe9IFNdJCNWH9N+1fbnA1PIvwEUq40jj8AOi/MuX+cvA8DS25cRRJ/1
yf7YOCsIXrBE0y/DJTCvKTNJABfXUwNZXdogY5DuF08HxyB63kJfyVifeb/5KP58
BRlAlaJCJf1LwRgPKd4ta4N+8xjtRBUClIHDU8WMe06nYzr1emXMr9iqpdFMq7GB
F7eqcgReUGYzhrGw6G5+CYk3w622yQfAkZEVuHcC5DqZ2fdL/nP+4fk+kAbGPl1T
zDiHJ95FzAO9P+o7/6slyHyQeL/4BOXPi+ZNyTKFOIHx6oW9pjVcE1tOv50l3lNE
ONezRjDRGLhjnCfi07H/DHpokgz+bG4A454862oEvRrth9sdAiOzZ3TlV3TPAq8+
IL7Bh+sde4/fygJIj+1FZSNwnqYuk6YrLp23tajkxsMzon8zZ2jbmwJDr8sWgQor
6DEtEwbrOPcePH6qUWMJF8xLOmhKGMmQQTrTOkyuENCW2l8N3ZriyFwHWu8p4JbH
yOCr4iVTrpB08jvGF4IjYFOsJdNOOtW/XLEuFSuxYjn8j2fD4mK+8eIjKEDGJGam
Esn/Tpfg1wIXUlEO8JZuDAWlOv/qxTU4V6wLoucBVuGYH8KmGy8ITz2UaBJrfL3R
ZDnotnQT6al6STnVJDg3MyJVYUFLHASOc2o5qz2yvteANM8NUbiR+K7pVQkihRTe
DlIbLvJ8o0usGLO2jm6aOFx3rv18dc9tpg80ALXffm91QL2/S+yILhqnfkeC90/a
/RVTS/EWiLBst9P9cSSKDMTA/IZt9dCsPzIKHJEX6t0fFP+r7kq1vYeruLZJ4/jO
lnonGOUsew+FbSS+O0b1LK/c8SzhPDtx5XAr8ZX6IPxpW5OWGq6BSUhWZIfyYMbZ
VHs5VWexoOrSDE3Wtbe/KCcWFUmBAZQr4OTRnbmR4IIiT66PcnbpqKbn/+MjuGTJ
r2PJelzapEcMJkoyJcuyyUEnl21EgFb2wYgFkmh4sYdTEjbNZssL2qjpA9Y2hISw
t1PbQUwmMfHFWayQij+sbCUwTyLchpf8k5sXBfeP7AY4JooZP/zwy5+AeV3/jz8S
vGdE7I2Sfi5z22vYNgllOPn3/7sTVCHw0Nnn1NhbmTiacYhqLpsfn619ptA+BRrv
3suAAbL0TtbtFidQuNwkiRPuywqr4c/2Es64szsem4wT1CkEAXqAo8dGoqvgESfs
ZCvSbcDH0adrBTbQPZb8ItYWk/hFdD83zNmHi7cj5JIdBZ4PL3BAGlbUJjRvdQX5
M9DecwXMTA8nH2VaSsx3a8NJqgXo2Usq1zfDvXHs0mwCrvrKyaKdXitVYdcpTrsF
MUyInuRsxNNDNpbsc+ztMbhpGLL18+LLswwXXACkf260l0WxGBTPLmZ6TUkvjNz7
d77aTrEuTLC7BsVIFY3TLHUmqM3kdNedvrmr8Egux4xuWk+oG/xl/4UxLMdJccui
95quKHy97X81nIM8BYeIpOzcPyvQLsmpznxutd3jb686LfALpLpeUdk4GkoLYUyv
HGjBOOI6QMdH3FI6Oetd2t6+4pupKosWtG4+rYQqrzbO/vxbkCLqNKapXGHbHzdF
fZssDz5TRtFXQYmN4YeVcO0iZ9/T8dQFhTNc3DAUmkXQDQE0EA7Qt8E03iHNVncP
mIj2fWbCDYLtbFTmPzntughD+Ez6Nm3IJwCs0YVoD69e7AWjyJAjpRk8MtT0BscJ
21qB/dKYNBjf7XnPv2VBz1y1F/cg0fBqNq2jE9bgYZPA4+o+SLMcY4pmlLu6WMXu
Xw1CJYL6H1jbMBjBm/PuV5rpMXnKCqvaBYCa+Kg8MY34JO5SO9aGBYreAMupyraS
FpCJbHIgMymxdwI49ge7SxLoppUyMKPVXpK9V4ltyxtbI2t+mQEX1Ntbdq3xyjOt
ZCe0Vpi5ANnnzje24d+zfQJYQqHWDMbh72hzAZ6VU2yWdCEfVaWH7akxGy5qhLTM
/pKnzR6idvM9bndO5GXwgD5hbVWaM7vsK9s1tPPGtSRuWtRkT8JFBfcx2qBdvgcN
eoSr2fOpy0Bx7VcWUqL1ivASLKWj4RLYVepMh9M0m5ewsWW1VSMjshyiVoVxSsKA
9rGJ1JWZU36kpopKjOAmmYzNsOWB1YoP65a/RhclR/2YDtq5BCVa0VkGA9gVcTNw
C2zU/ViW4UoKZ8pZVrhjkn0sZv8SqajELuH/O+MZ2HpEwQigKpWozuytRzPlf8TN
gXntE1Nz+goiODE8OW8ahpAI9IsyxlKnvGgbDlVizkRFOJookftzrulk0O5C3lp5
2fDsOU7kO8nkJSFJO0IgGUGBgdm+AQr+MWL2UmCUyrSshgUjEC4uhW1Tf15EKiRv
qUkPEHEnTZiCkS6cmU/g1mjC/TYpHNabKBOStWmuvfcP3sCCgwJ0SCmWTOI729F+
/LVOArf/i77JgEnVWMUDX6IEdGeUXrY/dKQHccuXZ37DZY5Un6jzY+w8mP2zpAdM
YjXLmvrcVdYADJOiC2gJmVz9FS7FPDoi7b0btB23MiJ3wjwPceGLTL49O9Yg9/+U
5hwCrvgBnERJBAsHUVVvdP2SbjHeURIiPE3iZvlGkdJr3KvQoqLTpOg8h3nqOI1a
RJ9VvWpsMHu5ltN03ZfB6+UJXAN0T8BCBO9kWajLlc3tOiLvUk7AZqHYDyZWjXRv
hBYCIqxhLKKlr9jZnpIFG5JEJRaFhNcpoLKVxP+ouWUr9JQtmOuNyLmO3E+BxUqw
dDIwjXXHVh/V0RVoISoa50VMUdMZQLPULhu1P80LHnu/HUkLDaZ7/b5YOVkZ3+ee
vhFHbibBa2JB8UwcvBwex47BncXk3q5rLjnV6RHTdBKwcQm1Vi6KeL2uSJZG2Bfi
gaxg7hC1lNjQWRAIy5t6NXEkbv4Uec+oThwbXmx2Raz+17julSh2Ox7FK/EAX2B9
Utdu8kVzDNsakElDWdGBj/iigYuORs4fl0/q2OqnRxjhGSkL8r5d7Z33k0YQ/Zsn
Hu/6MAQtQdabuniYABHJhmO4bRgEXJHHm9Wvg4q9HC0rMPTZdkohQqOEW5bbhAm0
IyD8bI4d9HJOTUgpkKuY/e7vzPViriaLydxbeIP+jCuH2V5nidlH4N+zDayliIb3
/Dba45QFRtWnuoXNinzIva/7jmDu+I4nxtZK9pNlQ2S++YbWvEk2x9FzjBqZ6toJ
RVvlcwmyicuPtxu4XhuaFdLC7HXLpD/mF8BJrjRNnQeDxeioSpGQl9XkwBJLaw5U
rs7+3MgkLUb7nr9zl+HKzW9aOQmtA42qFueMb/hiyVFS0+Qp+lf1brUzW9zGt9lX
+9WQhqjqlw1shnqmjybBos2659CmzjroBqgZe7y7NI7wNeeAtqxuU87QNQEiB2Ps
tOw+5WYrepwaBXVrfNZXF96TpybeWLWb/tS3lF5JLR9akvHP7UJJSXrg+CTrO9zJ
dTddVD+uZryNF6iXw6AAaOkoQIyPHFM172zfH2dEyYaGObqP0C+KaEH4CbdLxC9b
SskK9KBdJQ4LSuk3D4gVNzUBdKrws+Pl9W0o+hoUFO1vbU3aDtY0/bBnfI5yxf5/
brIxZphz9ADG2SJ6FJGH8OjSRRJZL5h50lbBMraXXVumg1LfUE/XkwZSrMJB7QKS
sEO8fvodumhsBvwprmoBVaYK7Vl+XoeMb/Fq7uhd7imPFw7UvOhxMfvRzXZ6ivRu
xXSrQW2PZgI9fBZWorLQQK6Q45oD3nxmIB0KTt8ywcOz+EUl384ppZ9Tss1vA8D4
OKfRbcwue3kKIWlpMPaiGWZTSWzkw3bg49TFB/d8Xz0=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
amEesv7rzRz7BD74gOn/1oIksgShA7UV8wnINPjYWLLBB3Y6vj2SrUmBNXwGLkJJ
JgwYbt67a+kTK1PSAThJsXGspuPRLgFy7vOkC4vXe1N8LNrOT5Ex8/k1IodQEl27
3emTpiSfHBqyM70wn6Gh0zCMZ+wdeKfDTIVJwb1OeRXF3510l+/aMxCZ8jx7/AFO
tGK9sqVRJKg6OfgyPQbNDl9En97luuJQ9qm5osZkCyby91wvcfRVRcgPriOjxB05
EBK+KO+ODTjXlRf6+eyinRUGD0Rc43/JtnlBv9En1WSs6RLzgOiWxFyJSpztSn2T
3swMW+Mj3Y5Xr8+nl+68mw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
Cv59BNIZa7jVG7uQrirfsdDfWpXhhoyNGTOxEcS9lLUTsskm3udkNhCgC9op3ShS
d5W4wyC0opznpmY6YUOQdTQ28s1NWvXRE/x7jsskIQJZ3r2Pr71O+Ci1sxM75MG3
Z9P6wxSZYf4ev5i3vDhG7XBT/ThGfqmjZiyicreJEXAcFbE3dBRSdymcXtbpcT8D
bLi2vZ76O3TrcajPMh3Es0bqAdWLvFXrxsfioKgNHTcVawa53XaFnHgeJaSLHoWu
XiBRn/PzVThzQ3RyXnRc5YrsSdANyFuzR0ejGWchqfzM5gemVl75HR39j+JgTKW/
RWcQUjNkbVP4YUAhbufUZcbW6/oU2wjW0bA2i7iSALB8LgIMNJH/Qx+HHixx7BsI
UicUSAKfSFG/GlvQKSX6johjGWmoGDST2SAgjD2LelwgiGI8WZMOVNxAG4dVupll
knFuDkwj/McDVDguYN4+FEd9sSFoX8hEL9CV2XSe3O8azHNdF4TAh86CkZgujfaG
OJS3nWTReBRFItGg+5qh8EFsDj/95VjW/jjjCjCI3e0fK8nAqVnMp2y/lGz+rPFB
VMZlC4ygSxN2OAygh0O7y8+SsBZc2pGVU4aUoNVA9uhDX18c3B2ST2iEA7TZBNR4
eLkrp1BIohISeXxs5Lv5G0TkTV2a4atw8L7olnU5ifzjDgABMW1TR/UWofQVJpuw
WsIxYB3YEJn1iBS3D1hl2oM41tRUT7tvdlxRHmFZHMtJtq+to1BHMnLl4U6iqZFu
ZCTl/F+NWRExqjbQPMjmIgRJp3RRaarzjccB9tcHWdXfpVZF5BpYBrFgMpm7rbHe
Q2jEebW79fYyB3EhjTsfAhumCYA1k9BsiLxn+M4+/gi3Ywm3LuKHtqjNJlGPfDC9
VifdrBmlEqZiknImMNr6Bjcrdsd02oxxOQjrffHBLBidvYoBC0VPRfWjxMXAun21
fr3SGnKFA0Ra5BAAv8BK63q12JrSK1xUC/EaN0Tonh+JrzRv3MjLB4IzjwOoF9oi
ydHeD7e6UD+QUaO1dVFnlijoXAkByuBI91+E4APsVMHwKpuM7po9nt8G3ZV1Q8gF
WL/5HLIRvt1t+t9ZIKXOVGl9b2n3/IsjPRgWWjj6Iwb6eaPCJA8s5FjYlDvxJiC6
Uki3j+KK+v9JKamcXU4TMhSOlCm3aNh5tB7LU0wWDsqAwx/IrpCBrqYJzf/60STP
tdn/x9DWru71wjFRzjQ2OcZE3hNraJGual0X2t3/HHVTUSu+d56+6F9I2tR5ii5+
552Y9kCXnFqxnixHAHqXTq0zht41nhXrlVVGojk2I/31UyOG+QGSOI5iLcBNsfwa
b9+f02zgylIBKevXsZJqmxPOpZE8f+RMlZoghBTrY9hyQsv1melVzdJ9ZrXFfu47
XISq7gHh7O5iFhdKzfcpC2ALx8BbsY5ckO+Fc2wjErderRezZRw810GWjVLA19B3
WjYRFD6qn8tGvyVDpsIIPgflmIu0LzWu0qlfyfMZnfOmLd57DO5wQ1C7SHqPDZjN
ecw0T3FE4aiagqFbVeXjftN6jBSPbgnLwmj8atx9t1QzCwjEPmBfjiTxOcikTuPD
BEsq1CgrQNEsVCiHNNw0juPGQtmTiyuRa/wxysQk+TvhT5NF3FT3vUzGT1CUCVaz
svaCkrE3LJQ9DROJSVZ4TYg3HrVpVjlYpGKqmgSNB1u2YreeERHzx7qovB+2VtvE
Y/W6V4HN7sbOherJ69NdevkLGuj+IR7IgM08J12P+xQv4m1aJB0o/6JkTUkRCIcZ
DJBifVHu4uUSyX6WH4ll6APkzzuE+1lW2Tk/IUKy2W/rvNwVWHpEznVt9qc28pq6
rzPVsMgmUaT9/gjbOmAoSJF5D6xG+yomqKNJsUodVUFF6zMlHYZ4jOC0oJ18Fiyx
2pExnkJo1FNPdAIAGBBoPql5dhFt2l13VFOjLUjMDI0ECKu0c/pNmo/21bi4jI28
JPSXDNCueIYJ7ZNy+OrUc2klS+nnMqnZHxzt5Nj7d6CQZAguN37zhKtoZbp6NjFK
KqUf7ysocR3yXQvZffQs/t2G+D6IznupCkmjbRvg1zz7XUISlmyzGYU6Zp4FXnPK
j6h9PyFjaIeqSL3ukvEoywksRmnb8uZxve+KqrZ7iXL0MKGJzGHUd1wAwLGuFpV9
F2yK+Wv9tEnwP6Kz1ZCY3lSlMIUia6GsBcCDadWOKV0q7pH7VIL1Hv4c3AJ19LKv
8sHuYQNV6CbpjMnGi8jR8sLAx/uz7w4TtEK1sFIB54JTtonve7bnq2iJo9z6JnCr
anSAb+6iUJLPzV+t95aeEMOR0fYcxHF2Brhg+fdJdFSUaL/9W/3g0WTV6ty0/pGS
RVFthtbJQQPrKN77qNRQMkC809EPAcuKn6n2o27RbB0rJC+3+LiAJpKDgLcv3P6y
y0abeLo0TewVpuRq5HHVaAQN02XTZF9xfH/hljFNi5ftQ/eGkew1HopqoMGRPH2N
E86UTT40c8I/ez/5lt8nGuxWbUw+g88esqgHDIzzmQpIm5UOj6CJLMVXKT6Sesl/
N/Nxio5nM7TuWs7VKJUudHmfztw4AyPZcsPu0JlzBX3BRNMFwxlzoH1ovbI/f0OH
inwULOdHFDYzs1qdW8Z5paQ/b8iQQsDxildBktbWZtYwmWB8YMRpRUiqoLO0u/A3
0HzXkuhGKIn7YAV403xXOwkpdkQJeSSNrVf5yyVFEuZvvCHCb3VjHdmyi+ynNr1z
FLw9XL83biRuzOMJ3QQS+mMl5hFn/pRErvrLmwQ5szO8u8i8j1SmTBk+dehP5RqN
pFSh7OZpvXXAYJbKn4JTpAwpOryH42jR2qC/dADBoJEwc4IeI84+1URUuE/pUjYX
bmOGrWyAR4fM6Vq+44kxesRlYeu24/FtxPw+SX+mQ3MGFiian9E10CEcmaDxBKhC
l6cp4FUOBIc818LkcdJPTJVcN0X7FJmfKFz4E/p3BfH0Bnp3VpphwVEPYaoJB0Cq
bcDQt3xGVBtCvWLcDfbgRove0aUsX6sP5h7o36QzM/FZ7ZOkNfPo+z7GmBA7Ijzy
BoKgAp0ELCShFVxi4KJfeYxtXH/6QBd82VIbsTOa3Nb5JPOAWoJeh7arFWBw9Gac
mDu5yNgofixkfvDmagN1XlIfRe+jGh52KPvzkKLZUqcdS2iXGxHIYomsJg3IIixW
jHXZLIpd56po5RweXZwa4tq8JHoPQMC1qkjGXGk7njuwVgLyIObs74wOBkXpf6VE
XzXswWVqkCR9Ez2URhQnVvIUJhlgeH/J7tkcR7MW8lpzj4JJlHTQdz9GhLA7o0Ri
fthPQle+fmlxjKmVYAmj4ife3sAD+ML1nJSlgh67asGlRy42rqIJberb8BoFtk7T
ZAELeZO15Ia/yScEcpxS3pW9/QUI/Z+TFsHn0kJxsgd+cHwxy8kfSV0JfQVdpsem
zeR6b2PgMsTE4tPQF51IeC6nwRr7vq4cwRSEeijh8KiKX4M9jFi9u3PvArqLo6/6
GkfgSz75xPlL8+MUIiuOikIlfHaNMi7c6UZzGQRjrBRM9qjFhXBqMKZvMS5h0vfI
/Xc3yJC/OqSxnDeBekl5pHpNBJdgUjG/M5OyYzK6Lzd2HQNXWGFBpEQp+PtBZgBP
a4GsOUyz82i46QzLlw0Qxt4PYH/ifYQqRaH+WyEGAH89LX8Naq4kY6nbct8e7NBD
zmEQnnrr5yFtNkFSqndJDOLRo9EkOfvQle6F81Imly341SmZm5XRErT02Aq2u6uH
V6lQHBSJRpqol6vJb5VKlURGro7JCk7eHYSiwhnzMlssH/p2r6j3oc4iz1xr+6q/
P0rIrIQylK3uKGXuRKRHL3grG+PF0udJT+IPskN/XOhkajtZQuxNvdHe3DnOQuu/
ey+lJ2JQjdtr5EavXMEhWG68NDS5OQrqa8MKVxvJ2UIkhXmJrA1+F7Zu302uJ5R3
UZGkjY37XZGPVnV7F2N25dDAPLSUyeXeJ7ok9vloxN6X+9FN7wofj3ZlVxlr8TDL
Getn12+7k2/tdb+WGSErN0u9jwWuVD5qwx4k+n7sqaF0AyrObOaDd2M5l1TrPnf8
Id2qw58re0wTpM20FfS1qpoTUhWE6HXZ4IZVKQFJMThmfYkCGD7mfLAS1h7oSCrx
76QKymFImaFFvvfKs8zEzb2V+9Jj7g5dtujAoEgZT1ka/fy9qrOugX/MGIHwtn0Y
Br0If9WHGPXbpXjBXnODypnRzxOIbcXeOHkcZ5r9TP2tj2wIAoC0JD66oebp4lW2
v1+xhCrgXnI6GxNr6FMn67zDwZf72GbOC7t0IxsNaptFknLtwSYz5VeF1/gSjYKX
I6zoNYDCpbOwsgK4yQ+djWU7qx7aaLlheCA+2la6+rxXhgjB7vN4KCWhWPDp47ZL
yxGN7+JYpmFcXMFfTdPt4TSdvyUD5Yxc0LaQIZ01xJSZxx1fszZawYqSEyRsQX1v
qnA99BdnhZTtawCx9/DWVXh9tGIOLhJnssPXs/EdGawkjGzoblr+T2hEstDHKaA9
si3olLIIJsdXCkbJFGUC02PluF8D7b8/QlSX+N5KAzdShWe4BeDoWCSXgAkArBQ3
+TasBxJvgGK/Wr89KmSqek2pz64JIhkpSWHI36yYVmrylWAwo/o6tw2udCdbuqWp
HLGRj3TwWPVTcuTR+Yq3RH4A/GEj3zBDLHZOwOAzF9MMp9xTAmtWsISOolE6fpQi
6AUPUxbPK0mTZx6mHGl8GBiCLHB/wm+ZMEzzFD4w/+24dKZNDxoICGnDCKhJQyub
zKfVrua2VkNiuMSlcqdj7447bVzbLbv/9BZt9VUFXqkaomVqh3WYgfET6mp+Mb/C
lkeel6hBoKOvCf9jHBTud7umQWPgVP4v785V5y6XF3V64xb8qlWvEeoLctOVl4j2
O0NpPK55AURob5MnnQigXX3J5fbHL8pPhoKGVcHvVfAnmzGgJIMZPiyA3YXd/SRC
muVZZA2/iEjXU+vbGycYgMdgICCHO6lqJpCkw69o0JJbfaMs0cRK2Oj3bB9CwCs+
SRB3T3/5eydRuaEgm5A4sqUxZCwRcVQEitFnPDMFXTVge0jZZjyordRhVa9s2aaG
g9IovL5pcV1DgjPmp3bA1wmFunAzke9Azdzmdm5CN2pWmAqFSLxu6sjK/IR6xgIW
4njI4i6kW6/DXlaMXlLo6ZzjL4t9L0ZnGWFuEm8ZgGzgvTRUIOtd/LDUJ+VsEV0g
9qVQNnxTUh4CnpmYRq44AM+8dQHJ1PvP8xVHMsP0slJxljCW4NaUBWbuYrWEoxUU
FPbrtgtV/nfYuGw6OFHvC1vdi6UB8fq9V10p9yQNd6fB9+QaFJDL1HLROc0MHrgr
VrjBMLsjPHg0W7hndjYZ9vG3hwWYlSSFXccgvAronRmVkuB8245C7QnhWOvogbcx
VFnEh1qZ6Z1q7hDhcraR3behdeXL4IZd+J22isFj4lKbRbubCYGYvBliI5Muh9M0
d4At8g4TYCRbVx1n9+iSzrwXuRLld0BtXZ270cmD1dmaiHbMrX1BfW2qubLamMxt
dS60DP5/+JImO/CqhEHe3HmG+XX9eVKrIsuCeivCfBdKecQ4wo/aFQqDsJK8BpHU
qtSTi/XodRnnbEgOGOMcx8FmzELC0wYmn4d16Iwe2feqMAMG3t7ZAULFT/SwaoN8
FeIQu6cuym1gZ236FwxrX7R+stbqadn/TW9mNO3jgpU/3/6jdQRWige2xUjTmtP4
KOky/j/IzsrZ1rPuQuAaGWP0zoJCq6I5o9GUhaHcpPrhU1kOT5pTB00s/UY4gLjv
EPf+PUtiqEFahOm0kyRBp6zlW5WzgwlLdAE3ofhqbhfdh53iRgJD9q+aDNxG+T96
HupbbfiFIM8PefYrTeMD8LxHB2gpaT1x7ujBF8xYjGsCUxDWX5l2+RUAGRheDZrj
h0m9fcUUC7un9fPdea6ihr5UWCeKN6rs3A5pE1hZRmNyKFzDZ7X8CURRt+H3aU0o
vku/uuWN7rJrzcJ1lynq0/YPBRSQWdEvQmMEcZyYfHMLA7uD250OpCr3qVM0nKRI
9h+2vk/XQ9+pJyMw/EsZUr5hGp1rjbSWNpEb5PfCk+tAVW4LOa+gLdeC0p8bcT8F
SWy1+DZ2PeOhmZWbfYRgbdbu+/mcQrmfjiLCQQN3+iluiNjdk680chbmoEcfodj1
iIq5NNH4qSRJ39Ii9xSlQ936T3wV98pbD6TPT4WZTFuQLrBx9INWk4oqvPLbkexB
SfuKWdsz/LZlPBB1Iwc1Mmw1gPYAk+1HZzf4H085Z5rwzNu072WcLj+CtC5lEJC+
rPMZ4bwACpCqIkgbFFx0gh4nKtC3g+MGejcFPjMWT3a5vt+Ia6Dvncg16bAojgHW
F/cMAdTr+OKXxH4WRkF840EQQtKcmdNlepnM9sjNNmr+O2S68TU/kfw325+KbBA6
W5O+dKurkpHcs5l4Q35vrEVDgJM8aWQZ1BN7tMpv7EKXdQ3MrVZHe+Behw+tp3SL
Yys3St1dHZ9aOsNqRptbGWa4KfpG8GERBPStkfT2vrwkYKKzXdPU/DTJrnamP9iF
vlEOLZtNmICWSNSrKVhUlvfZgBSwdWByzcGQOHJLpgVtZruyIXvsMhdSBhubg1WL
ISXju7lPSjg02f4XoJenGHNnJibMW/YTI2ZXoBhZ+ydbss5Fji3lMKZ4Rdaq5u6P
rnROgO3tO8eWHUpCq+0r6465VkwBRItWvngFG0zqQwYJKiaf4HGGaef5//OaB1cT
cwo6q175QT2CF+ACZeOeQu11K9JHG4kByPYTrhHEqGNW1PQPoXSlyAo/XDGdW8Yj
da9lgeEg608uKnvdci4kDjmTgaiqAlLSuK36bfj0+1GPGVz4ZiwaRIVnwwmaLO9W
L/rAd3SnbqZO5ATCaKqIO+QXFV+3iRUggTiRH+sesa/7+zNHT2uwDRRmihOMjcRg
q/uAdDX2LNIcUPSwu6J+rVzaOYwMoxOjPBh19kp1Aeg0PQujwLGC9hP/nDiVEuyV
fjQ40LEOB699mHHQEk1BBEsEW5hDwK9UkRVp2x52UoBUbyccKH9oaw9QXz5SgOzd
op5zE/8jjcjevVJ2ajbCoqyck8kHwrJ6vlL/xPlkKojbIoriA+alQOVflhfizUzG
AzAVHPtq5ygr93QDkWG1xcSj8gXBXa81SsdXTlQIkw068dEZtrYZv3pIdzx3kc6z
O24o4vYC/5r4bd1cYZRgq00K4RGxq5iJWd4tgmg6qFtceA2EYvwqcIZbYqv48DsA
QRqYAEOxfGKNNuUMv2SHpY8qOg13jOS8FboQthFTLJQSiwPPeUXzVf+hqyLt+Ire
YVfALZsFf5KPuV3Dpw+zFGraNb1/uDIlRVsZ7gQv9NWzcGNHMtT/jX6iisDG3iVi
Q0Ovsd9F8eDKXJpRj3zBmEbUNkrHvzKQ2uc9umLLNb6rvKT6PfbSRErrHu2Enrb/
5g2oeXEO0VGkO+LIxoTgxYKS1APx9bUMUYmujWgZovmEYhaMZ8dMZOJEfV2c96yH
I8QhVlx8Flf7HyYfqtyPISCCfkY/V5xIFHD+hvHvrND5YIw599+E5jv6fEVfWvQP
z9pZDCDJPhK9sPeFMEIVSSyFoDISEij8mK3pZqb+hdsC95XmvYhbpYo/iig+GkXe
dp/dETHkdlEEtTd+kuA82l633TvX0ADhmm38YQvTJW7uk4fG7ky+t/GkZigtW39p
7mE50g/HiJwtmPBRzEQbqgeuk1dpHHxO4uZz946/gGPOhaKxErs6Rjst/QfmUPpa
UGAMF+5TVnf4PPMYdP+6slf/yjKR0FGfHeb+u8bT77b/Lje1rh7cJeGzUFfNkCAG
rnvWsisYUdunFKlfkEFL4jHdtpMxoZw7dpRisZNI5paD0X1W3AIWp4YMiGsmwaYc
snnWTB0PjfJqtEYrZ8/vj8AufG7yg8IixQHbfPuaZagOAXzHVdL3EOagut8vaGZK
z7kNQ8LeGSzHsygIKOOWWlazTsA/xVj2B2d6zD6q9csApRupHPwNJzpeP5iC49nW
MX3Jdjx7GN3Hi32p9REl1DuKc1srJP9i1XzP2SH8Kp5hFNl2xApSS/OViubV3DLg
g6iGIIFzmnRbL/gWwiLf7PaHERVW4E6BS6V33wbAkCT04qHR/lBVRuhtkG99Udai
3tS4mA3+YrTgNYVJaszf84QEMAY5yPwnfvYkTR6mhEp44/cMkVid5zbUMxt0ypq3
JDd9tnM0NlDEof3LBrOrTsWQ4Uq7COo6f5Zb7LQbKblxS9/LaMTaXAN9IogNIC7V
kzPW26epIzS7v9CZeVGeD3KGOqUpQSSsb1owdHjdvUTr8UmygQtH7kwKJg/+LtdX
cVTWt2RsYzxtxJKGOahVGlr3rTfYTyAv+/PQN70YT303qfERqdN4MrjfMnwCgriz
AN8O+rcmQcVSjdnbQBZUV4u7GQw05EEjE2c4ivdYVfPJKcOFxwTXL1xKX60Jcqln
QrsXHKUMc3BBN1uxO1p/e+pHZCyKptr9VMyhFr+xNxiWUz8nS4I39txgk646/zgJ
cyOAbTC+nBP7cSGLI6nqsRLEeJ0hs4flMwcQc3pY+vjvHyZROeN9L2j9ABRTPN3f
bFreJiSqjdfAmIB38UQcrUSxPB/LIQ3Ho5XGfz3iQwq6Iwc5fdDlRDY6yEMg1P48
TrP08cBkObldrVRwXgfN0mpB9KTgE26qVlP3CQFsB9cyCI/kEfpfnMn55U4Eakjq
1gRKrz2TevskxxxTREUi8mYRsDYF2r7om9zXpzJ6PJ/9+XlI8EBas9BaY93HE+fw
1uLxpS/7QJ8fro+1OChZKX/Wn3QcYbk/ht/YPmJUrn4AkKhyI5GNODz4rsmDdDND
nnfuiDc28VxMoayDLpObWCAJb6yEm4B7LXfbtKpNlJVYC4dThcnVmKgNIu/F4m7C
tdBHjdCvXa0PXbi4myNxY2tn6a5BtL8J3aRrvzY1kz10Xe4BKZb0o1Su6VMzVLIZ
bHAG9ZGlmc5Pu805tkJj1tMPXM46r2IgfqxRpd28p0qzZkKiFvUAgj0sIBA+0bBx
mg4Ow2ODP0U1+dLKTVATXyMre71tDRipQDhEi7K2W6VXpurZrVgrGGe5/WTbkaD/
+ZmTUjQ5rEz86p74AaD1Dwpojhk/k/SqWqYbruy2VzIUhGH99T+KfLmEs/KIoCeZ
GltlN9RINmq4LG4rVKIecH1YVt1rGeiBJ9IpM9zaD8Ojp2s6NXvFt9RxzVReICLP
emaF8UOLWDQAGtbBxor9jdcfc4nFU5JVPrsGSv1mD6E0FeOOSXqayp+FH157DPPL
o2i5r4xdL1l8Zj1Q7GPGVnRszlaFmtj1WgOiBe5Dtgc+DIWm9SV4AhCm0H0Hg6Qn
vhVkkxAEzv/Y26T3uRQlX8GbZhLw6GRymQyB6SVmQqamALr02rYhSAgcqA29lyKM
6NWY9x10d8as6t2DZA0xAIdsVfQ042+pgXq85wZZWYUJwYTgSAWpnKHfIQxYKk8d
R53Vf9eb0vQhn0cwUgH+R5r+AN1oWAF2YthHkOQ63bCCkteeja0Ce/JArd7X01MH
2egH9j/inb/yXlr8K8Eox3SqqS5TCZlskFEzpdfwmGEi/pxbTn9Sw37sWGWFW8P0
cP6Vp5Im/Qk/c7iP+HVt4nRXLQbC6d1d7rtvruHm/nPaHDawjyZEjqbcOJPqAsCI
U9992ngXNZbq0J5Vkmw3t4YlEV4oFbCnyh9Y5eldABZj5DOZFlUnBAMXbAX6d0tD
Xux0f0RPvM5dUXp4HbTbmM2TMKuAEpJptKjTMA3vE3C2QzB+2HwODibbNNgiE6vO
lBonsFrnUGlkvE6TvSYRe/e+fKZ1ZbYzVBsvApnKUNpFSV1tc1FQ7KCCK7D4OQPr
gURY3pbdWOBCEvGuGwiLEUKGduVA5SM5i4y1XXDDfxv70IN5xdBwCAhldGMUOHot
xfiFfupVPNtVJJ5E9vmk1TwwakCI0TCOUMV0+swFc5o/XB1Gd63oHa2gNFbCHQwL
PwOEg9Zxc6ONKQZmz6gykcFfcDiM/wa5z+/ogwpCm4VJde+gWotbkMKa4M8bU1Nq
zjnrSlHrIXajLaiJ/iGk5R2wIH3ajZfrRd4UGjanKZsnq3II7QqbYEKMpQTMb1eI
yPSxnQ6uVvDKPpbgO5kO8VkGTLNjFS11P8tSf0n5f2WRthXafojdf4KPevob3A2Z
smFCnCvllBx8xFGTihnXYMQToFuTX4QBQJUkwik7qc639Coqa6pzO0NCIahXPvtM
aRcXRK+wGIS+p2Q+ahlUNPm+WU2Zp6XS2zvEZVCbzpebQDFYMOV7fOZWv7VpMIS7
rxSTeTiGNeipaT2s19lG1yec6AYfRf3dqInj5QK1LnpFEJx9oISWfSAuQ83ItufB
sHZQ1DZh4SOUOal/Qk5QnBcVFHX1m7m/mqPi6/nY6/RUTpmM8UcY86qpZ+5bfdDi
i3MznXTfEuBc1oKKn7kybOGKbRnOFnzz3ZKKv8/MXEQJzBFoOE4EAQkbFLTvemDY
r2FK0NNaBBvp52N0aQH7bbiX3KUIsS7ZQnharS6n6qa7ISs14Rv95ZWu1BOe+W1s
PttC3sq/kg8wvZCzHi17M2YuQFZfaDdb4mvykLinQoBPnyrSURURlpCPRBUdOwzY
DWod1SIL06hl1l4dMTZFDFnBQy1f9lVBOqeecZl30RxLU01rOwyuar0FIU6pwtgd
FbViAXic1j2KLBppPnfEkiKzWNIsTghpEeLbE8Y8sXySFfZ+FJp9EB4vNTkx1ALX
1QnaIseF6jZT3OqzNTtVRorN1aPL+VG9CQhndzOyIdRkl6zImNPFossX5CEJNDxh
aHm+TCmwmQty+IbDcJIxv65vubws/sfdHQMh1lzjcmn2WLrKD8LjmIGd+/3usLuF
ZBC4e1RxGHuYarG4xKOJi/GyAlxsR+Upa6QzQtgUpfQ9ga9j60ywdd46458RJ27R
JjI4XVi9Mh1xa1JsNb1WtStHLS1HWmDvNbSedj0rv0/H0GC8FiPFPLHVfTH6ikmZ
6lQhLjCrGjAywuO8PiYEXNCm2FsAPb4NUC2NrDn9JcsZX2hrtbrsQbFEhN7YYkUT
RrLscq9Heuc4SM1H1c9SImhQbMyB0Mz2AE2/iBTHmCnyPdAWkzhTq1FHj4uAyBaW
2V91DUzcd36lucSSshGUgg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Xv/AObL+AGf1KnPVbkE5P1Q/unvohzf6jQO/z+UB4ReovA2lx7frkQs9O+sz8hwj
R4UV3MosPUAn0LPKiB8nJKZoAAjufaVbpPakGdLSxILen9DPXzsdBNcynbJ21scu
FV3qXZZpdAZzyqq8aZ7zJBSiKSdk2kKuCVUACbP5UHK2AePDL7wDoI45wOey/MGx
dnI6J72AYDeAl6zD6aTFgEhq9f6dloydPyXBIa4sy9QHx4TamvVoa7s+AhkztC92
Ta4oOi/BID17uyl+J5QnFR/Z5RAvOIj3Su2kxZYzAWJU0h2WTtQe/EuoCaSyK3le
9yDjb7rRW39A+qViopnCnw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9840 )
`pragma protect data_block
OrKGnf5mlxL+FsG5ZW8DLQsmfEvlEecGAdJ1Ru8hbBDyX/sZkCKkd3fjz7MQJmkd
W5nKHRLOQ+no0CU9ScsGZRZq4iv+Pf7C6m82wkLj3mrev65BO5L4v7h5aD9qxOP6
yK9tcG54/nFWQiRCVQyYns2PcWqo2f7z7YecTBpKm8InJZWTJ3C5DOTMiqsD2jl4
6irLe4QQxv7jLFgb7x18EsRBqHUFPNN2/y5Gv5+vb/Egp6WK3QSF7oOt1IeigNjO
cacG29LgUqEZgCIDXQnzqlcsLvYoHN2mtuMo2hNyf770PNamQ30ktQ3btgQ5bUJ/
2ZfllZ77U0ASiLi3SN+XHDXeD8MbxmTNuMuGMV/SWJoIjlLkNRFqFjIF4FEvSxCy
mk7vtB57vIonGiB9EcA1N3GKLug7ns2C6CRp5nFUfM5OLp0vqhv3DdykR179uS7H
kO5diATjAwscsJBQ2PLM0EjXWiMaSxDe+yYpZAKTRWdWPpbuwqE8wLpokNI1acKn
LpmhDIYihK+hxp16s1wqXUMohPV7kVO/seIfbsTJUvmZZZ9Qb9pRoOxGffKAPrgH
wTUTtXCoqmsUgfCMubJaru5f5g9nHoj//Kd0bKlfbzeGRahlNH8Ms01svD3EOwa6
SroPxacHkmZcfoCWXEhzgXoIbCdXHJAUoMvxSPi8xz/fHYtGHTB6m+GPhO5LEJSi
tYVyN3a3iszBneNGvOW6ObQ8no9ESZFbAwUHXzqMs3fivwzoDfpVmCn8qSOk9KAA
AWpSTAuHhQV4DeJrNdc0o/ZtuPS3EecvXL89jX46zyIBD/9QNEVAudrh7dGKuLDq
8dri9CFPrOFg+GSpJM3O0xPAmH6qwEhtq1f/CBexoMomq9FJaSpZotltjdUY6Y47
dxxA2nFnw8HCRm621egk/jjUmK5P/W5cTSXr0wd9KgqzWQIAFZN9IVE7xMz4f0Ro
+h3TZrfFy5Inbmj3ap/uJzsO5hplMOwBdSNiBqS/ffL8gv78TCCriBPDLKNJNf19
nVaPoCMf7uUfhYD0kynvQfllCKG/vD6sT01XM9LBw62xSWFoTrH+Lk1vI6a85wPl
USRLDRBgCi7b5Ln6SRHRHLs6FaDc2aykciyiqkNAcwOhLLF3PbGvLesSVG+8AOaM
HYpk4OKFpbDA8VBpsrWw1o3fVy0Wn2NwklLa0PXRZIjVKHQ7I6CAZtYKRQQgJZy5
pxup4uQesesMilyYUsq5WNAaD+6vKtTstla2jQ3Ps7ZtRhMyurck9GEQhgC9SooI
HtN/q3b3zF+BHpaWR3WuXwGdEzNg/Ged+3I3xRKzrIY47ciMHnz6VwhKphnCtnOb
1XoFWr5g86DasDXAF0WzllG+JQeOvIA/xqYC3keobH7GXNMhAN6qAIy7VM5uLDJA
Dp96LNhTAJ8aKdzeQhPwpuf/edLn1m7ZDOaFd6/907xtNACxtmZzmf8tUNliPjvf
xjWi73rW0nhJ/yTY5K29FYF0RJ7A4cDGX7ozl4kPwTQ5Cg1iTlmBdiMYIGEJTG/i
G7OvY9tOPwZQCD/+oidG8kZ/uvaWWSWoLfZUT3YDqN8J0OZ2Wuc1pUnEpy1Tl/b+
ayMWAaGtW6avK3GLQNIbvp3iHgU34Q7TOUEwePc5v2qIE3ipyJyKH1KRQ/xjx1Rk
IK6ChCxhOn+WefpZqYWj9FZb8lnaYY2TEgmUrear1h/VwRZNi9a1cLs7/f+osCQt
qyWeMU+NYIzGXbGBM4dFpWLlmW4Ds15nQGU2+bFcr3dQTcwialBI7AhgXQ4jJXMy
MbwXozkmh9ylSEt7pfu3jGtmaTfGPDtIQvqdg53cBPGJt9tJBvi5DMGtA5qs8UBj
dRejUbQanMn0wq9Cp8PtmjXb6U7GZYGRDmgcsGd2c8Az0EvdJt7wukLKBg4stMh4
zD9mF82vlbVVixb7dfVdagf2VcsNC1nT1DuuJom3+K4gXBq8JlzaJrc2rNmr6FNY
cgWl2nV+KgFBaGNk/IclHArmZ9qEQCJ+jYTp3SwpYHZqC1/pRbpX5X6yYLRcj5lC
AjtXDBIs/eKNYqEje6lBRITJuFoY5s8AF1lYp4wV7TNSxhKTnPt59zKQwZNKp0TM
z7o+tt+cpCt3/EWpDF8pA43OCJHu5DBD0rCY4T2+273/PLQjr8BpSn7By1o5qGX1
hlMO72gsn0T/46UEBqv99a0X/6nbq5pW/HXBoSxWz+EhAWTuEw2SOnGzw+rjB1xG
uxotqNzpQXpiuWzog+df0ZrqXKqtAhIVBB+M/8YfCSuCg5GNv/ZmH0U7/0Gs5XH3
m/T52XL+Bgb8VjR9whayBIFh8YMekQwiqLM8gD8WU8KfUr5YGMSyfAYfF2Tq7VXl
khnVPLHNPSbbiygrVeffU8kuVAQqonmz78wGfm2T8jEpEFNhJwbCW47XIseH/6RS
4rBvn8DVqC0nXa+MZOlW+gZTLKSlJKQBZYHe5x9itzer4BwKm6h86+9FoyE63bx1
jcyB+zKMbZTRLVdgZ8Rst4r7YTpNvHmYRr0JU4yRqlIVk9VG5DgePrdELgj7kj5q
vFgxxXI9OfDNBTq3K3AMMlyi8irIoZxVrnim+HHpcSLopRbzq2v7CsKaViq8LULi
W/P462XEJiVhw+fwMnNeyfZvbWB3Qz6y5/tx3533P/ZxRhAdDcfff4m3SmgQFsWB
RTRxi3M4mpb6ej7uZTW8LtmOmMmp7HC3HG6iwcoO9LCDOtSWt8e5VmlubOykQTka
XD7/MIHzIuRVy67cEt3CNvFGz/lLZSa5lCAW45l12FLb1wAjBe3Dd8UwtPLkddGe
xZ5IfnB02JGUOs+PkvbndqPDGj9YcnMPPQOw/m9la3ypqo+W8kQLGnKM80IcrVdN
XFh5W0NMrOrSYnxxNIf56YhoPV93lCGFewvwCvMsJZYCglw6rBXz7Vlz/h+HvbHx
bunJvrWfryHdSR/pU7qNmbx5SFee+mm7lP0Vu1hnmPWbVBnmdn51JwZ4MFH0z0SC
lgV3T0szp/xVb5ZTD0+MBDoN9jh77r7BAni478H1/3/grpQGx8cdKGh7/81jGoBG
GCstLn1zM4c78RedJs3r3DHD51SCIMX/ro4/Ws1AT0zzWZQI/kCJWtYvYcF5Q/q9
BSXjT62gBn1Qsuxw6LSy7Q3+L5kOMUlGS7YaVm9WrUu8aOq0EOaEi0SL0eHRYrqc
ngMUH6DObZmSUYw2Zx5eRjtcbYgSKM+lPVQYd6PvLpvElrV1jIXGvHyYdn9Ppn3O
urv3o3kWL8VjH5BhGjU9sneUvE/n2D0gtVVApDwrB75mhyaQrWXATE8sEQ2KdRJg
uZ73OHQ5U0hF2iui+Xd+GiYiOEdm/hzysQUMHgACc8K32PDWg7tGv+dX0BKY3Kaw
MnfqL6pkICUkw56HfhGAAxhWvhMmt3ooDPu/D8MkuOQaonJOpiUsYS2vdEqrALtb
mjLyarMDzh98JB324+0LzhcgIVtOHB5QP6K+co7byqgoc5iC7qP8KTlw+YAFoyzM
vnGBpGfAaSn60u/a2BrsKT13xmy9Pg2V95HFLZwVomyKzgZ66o2C87CZeUG8grUc
JNhvHypBa9bPXaupuKSJR545vfFW3hCHgWc78sZFGOexpVL743/Yn5H+KnuYJPPb
D2v8we1HyLpzgVLVTAzfdAHxJyqyZBsBCEb994HcSTKAqlNPCZE4jwi9FONSvnQu
QenwAGd3MRes/pdQdDfK6pPr16Ro7ZnI4iMTgMzS4dAe//m3D4oCFxo7WkHknEN0
uRlRA7kCRNpITJKwGz1l+0IRWN8y4U1/is0vWAKq6Ekw+c9FLF0umsgRu/I2cBr2
8OBdeB8ibCevyaA5899G3awpfJAnHE+J5yF5S/kQu9aowhSX1pEy3uBXdJD9EviW
GEG/um/lY9jRIlpvLNEFfJdeZcmiuD78wUPo72K97tWNcXpMEuReXLcQ0wo5EKP1
ZfZJgyAwtY0pP2Ac5daj/lB18pQ4AO8EQqw16Dar3nIr8rwMW7MdFdbcihnn+2eW
GaXB/GpEuiKsQ7B7ZNpF7tBg5DodzKUTfuu51go/32IFzGoWaN6ZywvzH7zOMtBy
/KD4QcijSQzWRhkByJY1w/DW36zCI8gn+LYljtCqnJV0hqRojGytAi+4kXE6FtBk
MH7P1NmYExccv0D35ATnjefWGVmOMbdYaAd2FNEAgS/Mrb8MoJowPS2wzvoCVbcC
KDASFIhilNWWupzkQyxSa+9bPZXBg8qumuBbi711JNsOrLOZH/MvZ3A0TZXkiW+W
yChOC4b2tAtuAY2aDZw+Rd6QQNGOmpwCqu7jpVgnwrtL6RlK+z2pnB33orcvU1qA
KXraHY4etWk+UfCOQTpQpZW+7N01+4rf5/YjYf8TQmfjLqt/mGYyULNcq8Qzj46n
LHqcSNm+/rS3X9CRD6PZ5lp4fKvngx/yeucfKUiGxF1K9Duw+8YC7A7ewlb+lSH1
AfYGqefqQOtloEUB50Mr7w/wiKNl26LaSQswxgiM7AcGAIgT6SeVRhmV3MdGKt7T
Qdsx1XLgJEeh3XTBASBdhE9ODGzDv3LA/YSEzPIgRh0v1PVu5zzv44qO5GAmERdb
DWEbUscOi/cefjUk5dplfZuao50zxH5nB/0xP6u8tLcQLsIq/7CI0w/BxPeZ4BiC
/hxKqMWNErMbA9J9HtN/AQptMh5pRFzmgFjB3GgTNyIZNOBDBsvMN/ENFZ79XHQT
5sWeYFwqdCiOjc1q8rLgURoyU91pXyIJAtwGUtiZuM25QEfuQ+6UxlhyVJdKpe24
V1KNa8NrN8dEDRYjQgD1kFAhaB6HSFfrrIHKFAwmcFzkxyDJOxGc9d0VQ5ztm9RB
NSPpzdK5AI3oopp3DibYUykGT2rVYvrLw+FZ2rzBuPbS7qSqJDPFtNxrNnCpO1PY
NYHOz0OXDF7l4g0ImvXot1QtVBKQtCf0+zEUWG0hLdkr4MEK8lNze+leT2yZQobx
3x9b/7ijbzJAewrYGCWktoDB4fIMsYzchZ4/xHKEukb6LXnYeGKeUlNKnM31HRuN
jSSHqEXXuZ8OJ6owUb6qLjipNJQMyJY6eioRH1UVWQU4mW4YHD7naMP8j9zswKX8
p8NdbBEZxmuImQQLy6diUh7B5CyVpn2v1Kw28rFemOBtWiH6e7b77V6AIsmPC+pC
ihsB2LJ2XhFvLv9bn4OdtbCPDb3li1Lb/CZzUrTdQ3jTA+zdRQMDEBa1mFDMfOEq
67pMCohYsOEsdk6+3plslcwLvlmXYUIGezIyRn+YfMH+vL/piT40XR5zX916VeRS
jeTG/4ciNpr5FhzaVI5xMQtqVmeqmv1a7dBD68H82yK85EeMTwBDbE+/50NX3c83
fLjkM05tPiDcrYOAIFdeR4M5AcJUz+WC7QssRPt69nU8hMwImdbAaL9lOnUk9M8U
cb1xXcDWq2LE4iq5qx5R1TPpRxnz+fZFaC+5BPWescsefWVeK2ksULlVHJvxl6BF
LcFW+PYi6eNWe8sE6wccFa5yh1XwL7wFiGozeeFP+GgyitqFN2JCH59aAM8ScTXs
N9g/IBCOTfidtL4r7Le29Z+7HjgW0uO+N+kciAlJeXsX+HTELbpFIqngTN1vGiBk
p5TVEtWwQHJSGV9ilY+Ps7SZ4ZcZN27tb/oiKPAaAsLeFxlMvAwnQK5EG73N7rKd
JSTaJo9a7tZvQMiVVaWNWHfvZnSTeCUdYM+rKAGEsVVtw7s0hd+rd+AwHy4/BB5i
B0CEDddHVuPXtWiRtge2mcjbPo+TK/IlmDCqpDE04yGj1vG5AVJY56GFZ+9u/GBZ
MUrOK8hEc8T4Dm+wQ8aaqlXT+QrzBPFHX83b2teiirdw8ay3WpBfIRWrbZolQy67
95qkrKmB0j0qR2goRW17IHpdPkE8LUAajaHbprz8oRfpe5gHE2jatCRyZg9sYOnq
0fGI6hdqCsiaTBizHzCw0A+wG151JTi/NlrREkVDqAl4BV1jPhAx2hpSiZjPVDhK
U7UxX1BxtUJa58AZ0rKRmJkqh8WTYlg7TPytwAkeG7Yb2RwECy23GobhccOxt8PY
pEKbp/KvJr1Rr+O2Xz2wcpGwyWPtvn39fo+1LyE18Pou18ehH2+Z65xpzP7w7+yS
mcN4SbuQg6ZdFkCYug4Td7QL0jcPSBTcV9qc6AsicjX9bEqH3fh7CvYnP6+an5Pc
DyivyRXLHwZFBmVRUiI05Exnat35jAPWxm9ys3RM0Wh5cDFY988jm/T2S45hITYr
SKHi5B27kenI7bBw2ABHFwXCltdUKpaZaxkVz3QArU+YOZim3jXOA7f49C/Ni82B
BOYIrUYmmy01mmEj2qFwDuGzvZ2RkgEj1jyPoQEUO4B/eFtqNNYi6nSPhZ7NY0wy
oo45xE5uuE9YfRR/CytXdSuZdJuDvszz4XsJK82nHxgYQme7q7L54PedHAba1PA2
zx+F+m80vf0i7YDdqox+8OwGxbSbgKHRqrEYKU/YZfwsn1horkRUSCi/NG502+fK
lHd5URpNQWfCokxUrZ1N1/O4o3R8P1oevw/f8LPmZKQuI3aT3n2OMZh5fx0saLHE
UnvGREBeRaMJDf1De4RUrpq9la3mEKE44IP2CP57e3T4FZtbF3m3M7gX6pp/t+k4
ffglZjXw+IJf8LFmCGllvafALBfIx7dKcBTs8QP77FJM/rKnEy6rALfh5OBKfaB0
9TUgdtL3KFMk06+hr/k/I804WLAoSNiVclBFpOoceBGB+sNv0Ni1u8eVFIW4mr0b
s2jpvznxl6O0h02lfVc4c/OK+oRwH2iT6JO4ARt2XQCtvhpOia09oWBD6vGHDgA6
eOJHdOpYUkV0DHfMwk1dElg92jDFH7MlT8y1CkRGAdYkjuDrpV/H/r4vbnFZbplr
AWIGrB7mEJqbB/XZ7pQrYCRq9M7xvxHPQ52V+OJojcp6wGHZfrswuOpDSBy5pYQw
tD7BgXJZgBRBg/Pi9wXjcJ2U3i3M6vIAFiNsauReD+LxPqx75gARqtUm3uA3MGGi
I7lXbJVUtfU8NVzDduN9CLHgAMVhbV70BA3iKx5O8XUfZo65ClndjmiWZe0HHGze
kaVRrRLCfwc9VGpG1iG8UvTct8BbPjCIq+G3AkIa6LTdeOotroN2HsGtkk7DIV5Y
akxNrI3uz29LDZ4K1vZvoRwkEYL9v+PzoMJhqKoKEEVaDgALQb+cSoTCtJ1FZh0J
2UhHaXDsW2iraZRENIdGpafORUjL0ksoTd1cEcT1DmEMbkDurkaMuFcDSqBiQpHe
D6YdW8HMsh/Qb3ubZDJ6M/5VXDvY6LkRTiBRblrcTsU7YGYLm0tSWmN/fVQxQSYX
uOG3NU0oMddxa0gH/YbIB02lQOLcQvWU/rEprpDg349hQAcrehaibgSYff/0DRUN
wTstR1Qdga5OA3iRRrvil/iyTH59zFXKJHiw43BVUi/a8AlQtPOe25oTFAxm/2+J
3CzYdHF/qzTz5CGnMH3ws7REAF+USpx9AjQsFkYG2ixTSFWwqqRg+toVmpx0+HZn
Wz77HdFS8Qu+7ahDbjflfm9/UXlEdFvhD1CaCehdCEhHsOSePxQsyCItUEjtf0o0
UAziwJ5sKm3SfJxavwZmT/IeJIhVnq4xfwNnGL3mBZuewOfvC7dCseDi1Ok72xUk
7kIgIyLk6JcC94l6CzLyu3smuoKGDyNBzOzz/8mIQTKjHrfa+I2G6nFe6kZ0kfeX
ltQmB+JpYilNf0/uqUb//A0LV80D2kkjmpM2EjiG1Uqt/Hsb4uqD7dfDkNJZjfT7
6gF+ccrElIe70/WTlxcH+fKDyP0pg9l5imMgNtXLJ7KbEchvLXbORgN7agWaAp8x
9krDH8dWNsSk/AlXkvmvJ6AS7u44yVLkwanEfH3JphqmhAdA4lZU+rEm2fujtSPE
3UOLT1606CcEvQ40IIzpPzGWnvE2gAdgRuEnBGUCwpx75TqFvHguAxRJiv0Y+Xxo
gHxZwdd9LwqYzpBs4DdXaQflmUDzLSJFtLNGkzl01A1FDmLbdj514+yFUtQaOO67
BBY2tIwB1R6TCIJCuGV0e3LGHFH7cGJ4YQ3NFgdwTiuguiecHY89xaId/arxALEl
NmH3lcRf6vtisGtIWFXWR4UFcAjspZTgA5wUQHNoDVZr4S1Szc7xEPkGfVbk0RJq
1kEsbboGxtLibOZeAv+XO45qiL97kfL9l7L2nKFDh1sTCPLVbIu/6gOkzmjTQpAd
2WOsP/R77+yXD5cczEFnOd1kdGyrf1Bd0oU7AIw1CnTublEd1mSLs2QEZhXoh4Di
fJ+9cBKHnukmjonllLRnH3TBRkI0SMU3IHaWZUzuYQbBcItWXJce6iO/VE9v6Jkq
56aOnSfeWN0JxKPj+/fCIAb91ZHOZ2ttuGuOllLUS9vzAHMcPoHridxMQqHbR1B9
9fJUP+BVcnIu1W+fJxUIVLvmS8Wsz2y/vtsqfiU0mz2kggLPY9d3JgrZhK03mq9p
cMXCZP+nn+SovJPlFxpdthUty0mXeFzXACe5zHHxEnUGVXuynXhuT1eRe/HwVh36
z5Lu5208k+gXog158Zp2eOohJIghwNxZ/LZwW0V4vF1Kz7K3ti/oVyU1k8+qm01l
hL8SgZCrwCb1i1gKfXDLSSb1SG7QlPe45lUG5QUStE9J1irhKG1wnIprIJsF3OtV
h2PYvNKS2AgXkUwWQkHvxprN6sJ4EDyqqsFoEyJu2lJR7kiHh3G6lFB3UVTeGOVO
jNAq4A9lSPk4PbcHIZpzdtxXbzkiW9zOjrIB6bjXnZ6clslmGHalm2PtDiVMZQDc
0atuuc/aspCeAtdmEOUYnXYcWRlJlnbvAfiquqZ4fT9A7YEOPtI3zAaFoXGfjBwU
mC8Tzkf+8Ddli+MGL4R2tlV30cJIr2AVheSRtrcOxVzvKXzfutzRGntGY8HCDY2G
vYE1BFcu1eqQEWJkcoOJ6klcE8IrpBBlQf+e/6AuQ65CLsNEbey+W15WA3h0VoSL
YJGLOTztPiym0Ms2r/mdNDOTBnEQOv/tUb10y+mEgzQt2pO8HyKjRxJ0p8tZO5ro
mZofyKdeN/bCMQBZv5g6QPz+kDTH0j9pHSx7XGVV0cmrt2DujmFWsiiRof59wuCa
8xYmtmKFIbvHtkJgDEKjDHEPBmWVJf+Q+qKM+Njg7F8l6g3MY9l9BdM7jFrWqhwf
i0k8FoVBnd9QDl9ms/DDrOrW1NWx4dSv1DXM9sHidBxfUYYONGaXCrV33XWxtGCm
YO/z19Lu/ttvOek5y9EHbpZm0e0GNH6ShlS7ZitaOKkeXtNgmC7AHT51SD6wew+D
1iczuOOejQtva4uvWwkh6N7ucEdl6PVVKCweecCIMyAB4EaIENv2mTHZJ3xqUjaf
mOvDbJZZNNQTaXoAvpI5pMEYvUawQSeqYHRjR6hsOvc6YPxnsidLv5e1ahyrVbH7
TC+yTa056Rze98NQMr+7o8KwZrAi8vZlYISzX9uHVeWtygaGUFZTWI67pEHxjqeK
MLo0LhvPCT2uuCwiE1Hezad+JAX//NaqRfq3fo74D+iAB4a2UEeujih4gtUr6m0w
4yNMePZ6yqxSykx6dKmb80BlE6tTvs+O/F+akG1fCWXSNRYGyXH4B2ovDtmFpHVU
prC0YFqlUv+Zfs5JYbt+BLB96txrwMafwAY4p7mWA3I3CjbALQdfPsDHhBlJpBnZ
VbNWSQlFzRObhGMTGEjsxu3xod4odyHbsfIon8A4rWfPnfZpftzV8RhbSErfJv3O
qfZkgXuw3AU0lqclTUs7pM4MVtj2wrS24Hn7D6mZnP9dZAkaj2EVWOOWRherH97R
Vv+PqkakqhAMJ0/I3ZAARiuntW9TRiunk5ZCt9iDq9kvncqLO3k8G1Kc+MY+iViD
mCRipdlLYfwYX0f/mK4AWlZoFqNQC/lXY5xXkg7YwIkftQ5ffoOVbW1jqAkK01KT
Uk5k2/ZmzGV/qkdCBrWms8URbcy1TmFzngs1NjypwpH0DEbhIggXcCm42SzhHof0
HXTTeLvxe+OKkJwlGfRjjBRzqfR8yIlj4CcKGXHzOQqQa5o7IMgqJ+WbzEmmgQjH
8vDh6B7U4RgREsyyrYKpI7dGGlQHMsz7UsEYgsLXRlNmw+E5BAOF19hVXGgAU7vz
mcziN3/epbALZAVl7Eak3LwGpJ2z289X4JXBbJlO9JtTJ7ozhthilKDpHkyFJVRE
lbt60u3QerTz1n3JmLOMmw9mtKoTK7SMSr7Ff9t4owyOAsz20yDfEjO22xcDC6Oc
tPpY/2sstgFbjcNVMzpsTuKYlUxJnpnTek9th1kKdDqRhl4L6PQi92AMpRYUg09k
O30+ZKQyXX6DJ0hdewF54Nh5wexbDeGxkZQU59ErQA9O1oxRytC1o+G/vd9ODIPF
m9f3xXyU4uD19TZ4HY64wk6Kyp0MB6+Vdi8zrZpL0CXg7++lgLqHGpOVAIR62wYI
N6iVYCfz//Zp/7PYMPpkahEUPELzRNNN2MqcLI3ebhEnwTe+1qhMVsMUy/P33QOP
gvW8pE2J9fTgLuS+plwX2060Flrc7PEg2y9LYjQqorHDaytvw4aSRnBk45JSAZ14
a60l+8lwZ/Vnl0R2nENKbVDfCcHVD/agR2Ra9r78w7jot6kWX1aFOLFX8KW9Yt7+
IIRHZnFDOK4WHHeQqx42BssfTnZfMEcrr2x3k0fq1Uu/22cUZFgo+7aaabHciJMO
Kbbf9Gv1zGoj4ikyOiSuz/MhQqZ2AAHed01IoE1liIJqlm8bhBy4mpIjDIvUmtHy
ip998Qdy2WoQqwo/PprztMa25J3HSTWHmmbu4t+/ET77Bw7uTgw7HGZWg0MZ9ud9
qR5C0JhjLEDUxN1lRP/gHqYctw2EAWkJ8084MMH73CVKeWV58g/UrEtOU9jUAdHd
pe9WDrAdAK9f5Uo8PWvbT24mz0WYYdjVMhluzvgRgdML0jbCRPWZB4PC4tpb+BOW
ul7XG5ClsIWO9dcQMbcak5+C0p9wXNryx/6YnvKRg9HQVQRlck9Ks856wiF4Eyd/
bAuxhKtLJ1PydKfYezhNQVu1tyhqmwokoGvuR2a+E3FbRnR7rIQLEk01gnCOS2WE
dfuuAddcKkGom+kkmB3K02+XLY9XhMqLmOOmG8ZfLrEmE2WL40vh0LqtyTM8XaI1
9ch4h1j4FiX0rX8aa77gSJGinVYhJ5h0Ys50o0ynJKnwI4S2W5azFvDy1GnTiGgQ
R2CtSAHXhI6FcT+ow4qUvGuTnjhe+lCwLnBHd2cfga8qM9AJAUXQYoTiFFthx8UI
sPKkAj7th++WmXgJta0X4NHnj9DiWhsfl8svymKDCWh07YLOLDfYpsSEwpTmtinu
zF87zvKQkoCW+8XD7fyK+wCkah16lPgqdXTPXUA28a8h6W9ugG8F3RZOCrnUsZJL
D9UOjV1AI+S2ZvwY2+OOSQU+WIhkaUVtRZaNWd1h0jsGrHngKeA8ZFgYguN4E6df
iWi64y/LAxMf++d+cRAW07Tg4eJN/3my9KHV5zfeXJWacf1cm5Ur2YlsZPcRHRiM
Ie9KTgOt1UkSOtTr5ctgr+DJeDCHxzO3OjDFdLH/VHLfszXjODUaZI9uZdkDD+eR
diF6ZMjYMPZfBqjuTUCo9mKloDCzHa3D+zSQo1iVX9pOqVkBuUA7dGvsTaHq41q6
EKlhvPzY3DRoPJNCFT49fLFRGJFc9R23F4tUdrc0Y+T76BV+LKj+ad2yh7r472fu
NpdvhzjiweCVz351IsJ2q66w+K4xq5FcAIMiX+XyOZR+ASAWcfnkGFX5N+1vmp1N
JFyjoo8YYct09M96PNICcuxkLUhe9sGAzyXOSsMn2BFLTfUk/bvl5P2TYdEcVEpt
B04cVLrHvKTjiFWsL1jGCASRjY4Z3SZ5wJdpJ3t/naVjMUVPUhp99QLl0trxRlBI
8O10FmCM0ohmff6Rn7aVxsQNpXqSC69s4sdSIpG3G2g/y2KIY0KUzGinBYsKg5db
C+Rgr5dKrXjSTp8NpEWjo123huU/YS1nTJqSn54B4wX+APTzf4WzZqFc3EcDH4ck
E5XnpeOHGhueheWqHYdylrvLtYgUnvC9E7yYufHsTbCYNJ5+szqWYsVgFqOrh5N6
5g0jyBqkrfB/LO1pO1q7LpzNOD2emgGFCDDqOuN9r6dcUvty50j1rH8LarDIrLNA
fTZGKYMZyPh04KfJwwUGCT6rxOgCQKimeXZcsmm3SKUfexppVw2CqOr+t265cuIU
8wbvpX0QDr1l6tpUp2mVRkjPM3cfG1yvU1TDwlT7ZO+b9t4F0VWvcbRuCgis3iD2
ba+jBMoXBuBBWcNhTSf+epFH7d9c1wpV/pEkgV5429YwpcqgXxcAtGXT8A/OsFAP
bSFDCXEvFtvnAMeppepyMuPRgLeHRpzr1o70OI+mrueNKa2Z138N/ZxYxiCb8Ouy
B/n8MYlz1/TdTQrffV1Jkk+DFyroDkDATWdOIcm+c0m8SNK+4/Q5mc4tSXVlehb9
3WV4C55DgMTOio/Gl1k6pGp7zdkAfG106v0RCfNYt/b+mBxmznFvH++icvP5we/G
lyrQD8gskgYBUh9jZpCpHr7fHx81HqDtcgoyy8qLT++Sm9j/r+MCPRfpF7ThARy7
JMcti1RigezjvKBw/Dqm0WPMqVlpjlapUEKl7ltuk41FHjj0KOms8doAbhAKNPIR
5q95zwQ4ZBg7vSnuNOApPZjd1VylmcPElaMMHX7JkHrepVs0hnf7pXirpPDyu1WB
/FYN0Qgar0Iwf8jUSR5tOoGTeV0ahnadRdDgQrVwItjzpNcxUnrhAVRigpDIhHjS
rSrhjazsvflUeqylQlm/yXd2lj6l4qS3+4iRNMmETXwfjh20Ih43EJevcFSPdg7+
a/MXKDa6uU6HFrlR/dP3qoNqkR8fOcpci3MjgB3CyIEXYjq55jIph9683iZ2NkXi
tOmvzRSZFL34K9FOKKSHthpf8AeX48JyZD/frPTjMhu2H7xYH94iYTMYsdcnhlBK
CHSW9WMazwdsGs2y6UPaP6dV6ADNh1ccXNc3p+MFRqEfZ9F2hO644UkPmGGhbP7N
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LTiuiFdeU/hL6xpPYNNm5XNd6QNvzJLT7hBfBLargb++dyeUk9MEbo87ZJC5kDla
PnMAYmtpKp8LAXp6r4xuPMjYShTWf+UAiRHEIJDSs4p/34r9ucxO6GMk/oiu6q5h
02muowDnSrTLrcntt1eWEk/NrgRgtv7iYuCGK0YO974G9laeyyjIe8se8+8U4gku
bx56aOHhQI3A+EoaOx7zLQmZXtj8LO2b6NPrRqfiBXhz33+HQInHSfAaGcWKo2XT
xbqin5OAvzmMfwe5V8tirMIuBCSIHuAaqEXXucjsmqJUCDZ+mYLVHI2p3Y2bw8eh
C40SlmbACmTYkMbzFq7xng==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8608 )
`pragma protect data_block
zYo8yStJkUu5duzzlG9Ky+9vRc/nBAktf/a1z5m7SDUBVfpYHrjiWa2+HzWKKAN3
14becpyX7kJkbWb9t7DGfdhJ1tXmRRZ8eKWClvm9O06sE17idBev3VruJZWw+ZEw
Fj0uJg4trE434A4KBPH4wtibAe0j+PauplKvj+ZMyc094Fb1/9RmKdVfKfFFm2aB
mobRB5SZTW1ZjlK6gXTwiANXhJcnhL2LGoo9HAGtOP9TDpA8VICO/bTDHXKIamG8
eiXS4QVGLQpkRukjMKRb8JOZKvXaIXnz3FCbtUXlyQ71efjzoF+GzEBmSn4V8b9q
5HnnjgBtI6a10q+RJBvisqEOChQ55RxoZXWdMrnaOwRPLO/tlF4KGSUEdnBM+29h
XW/PbMVkAxv+S1O4SS/T9CHz9ilZgYaQ0VMjT/5W9q4NxLsnCUIa8bl3VllFGLLN
0DYZTD/6WpSKBRiOIpjw4JXfFTS/sy/j5qKQFw7CiaxRQPzixKfRDdQMJ2JiD8Ed
4ow7S3219h15ikQcbxJWrh/3FkB1x4LFySK0LfrzUAZ50eSqmwsoagZCjfAtVP1W
PRC3gpZKxMHw0n5pWW5Z9WYLhYL7oyr852xJe4pGy+UzuYrMcCcWD/0cWxJcSTy1
lUxIGotYtchakGvYAGoZfDcWqn3i1dKj2BpVYFP/z0UXcMcPjpIFWDrq+3sctwfD
f8V8icIEHlrFSrl0ihmmj33AQVG+d+wK7x6QvJqeidBszSMO8AFgJD6eFRKF1zQQ
qTRmu9G97FnAG3cJkaAUdHjmBXjcR9qYnLPKb/Z8tXDoxBjceaSr4iZW5PyNo/V/
BhUek+jYdJeSCgFQig8DTbbsnobdN1PDWGkdUmsSXOt9UqgufFHtJzwlsWUxgOCp
TeBwU7BY3k6kCb6P724I29O45+mz08M3TqAOU+DRnzbPe4ExTVXLisesN7ex2hhv
zm7Taz5We38AoKEn+64h6VA+KM4+nTP33EoLmCySVxt19U5+kPgfm/HU2lHnyQmX
pgA0o1op+9E746P4N8GqDFteP0q7y8BrGo/laYANtsN/CU2BpDc7HkgQH/DyY2YH
DEwIaP+S6HdnFm/RCfZimYNttKe/WgBJhBTLXlbremdtBbSFMCLIjuidRW4ljDs7
GNo8GAFe/YFX5gPfa5BAJsNux5DzaBnvErRgsuzMsFEkJj1GlQ1UGYVd5IwWnOGi
5jYNIF5B/hgBcL6o1l94/eLPLjIxIYvaGGHphV0POPgSXoATP5cbn2jPTdKoE/c+
x8oVEIVTpVAGE32vc10qnvh7iX7wbEN4E9DCmfQBWOf6TwFUL+KE6LVO45PhdUmn
Fpag2DQ3PQk3RYRBHbu8rnA9dYHcOHpwfcrK0A0XqF2WI/qeHD4o06LASs2xUkOj
3VWYr8J2LPdIO2iTSNfZy89HXiFMzaKZAjFwPdGyvtbz8tXn6ZZf4E8I8B741WbQ
/ncbJlYYy4W3rj4f6d8C57nyjd/Hq24k+DEaC5QJoINzVnsvwqeaBKWBIkcrxtay
RU4SAqQjjSPuTm9eqTnsQwBIE4oY8Fk2yQM+LUqzCG8nEzcYkxtGp3dI07efgsIn
mdbhGdmPYXQF/dI+frwPdNqaqZDZYPgRyE5v1iE1l5A5fMY9rKZQl0frBzhBxAAc
EFA+8GEisdU1a8wdDkwFq8TTD9NQOxWwWesO8cdy4N79wqcgRrSxnc/KdUI8eWlt
Dn4p6RL8Lz/IdEAUrXPaOYsmg/M4OZjxqjHI/eseG5KUlsUvSi3/4QEZq0V2wsmH
UqSbAdhdH0E4VMbwEGRhMfi8LMvA0bQDlbU7Fb8+ZvX0bQHh3sS9EVJ2f1dollVE
RZ+UXTNGK9I0C6wMsIL05JTHe2oI5iJgXA+Ps1GORUD5UFX+6hP5ts1j+BtlORxj
4xgq5W4/rfSh9BI3y1qIH7zDhLD1ZcXntJGCF49bn8xt9yl/IJUTFxCzFBd3d45E
C4E6LxEuXDt++hfw+k4vBk9TV0ivduSLWcBvIHDDxDZrNSESJBfmKnYXe6e+v9OQ
XXG8fxDjuq+NAXfFnQ6OXLmg7JmyQjLZnyubuUVQWrENFJf0LRyieui5WDx8KGuD
b1f73AFQAKLISUMMBfa3v290514F6g21+HwufiajMs7bChBZtAkmapluEXTOHM/x
IjI7I27U8WZ479KwozkwA5F5NVT4S/graHQyQNnhXc4r1Xkam9IBY3Lmn5UnIWKD
qZ430MpEakoVqKX2ytueCxDB47HZkvKbzXlwE5nY7EdllsrqUFye0pEbBgP4/fya
gQnKWOp7b/XTI+r3yyaAYLBg01IxoyLwlA/NIzgJQxucFldhoMR37bHCgADm5DTi
VeHrEDAa3d/87W8OM1VrbBwE9b+qgJxp8yq+/ZFxc3K1R0vNi4DRG6/U82eZln3j
zPSd2woKpLWZZLnFbNFjTCGC4XVDgroaToV+4zlxHLoxLRflOW0uWlf8ueLSbvaO
vNz/Pbxvvc7/MroInUVxh74/kEY6eWQsvlH7wECeFXhBNV+fvE/qGzACvyAw2G/3
J3tgwDphrbTv/exvZfkfJm063gp2WLll7+sJyC2YdNuQN+k1R0aYBoG3TWmW6IU+
Yt6akXfwzcUHTlI551l1bwQLrXX4UKzz5gNRYc3zc0cW0NX3186MB6a2512856/n
Zh2mcSU7zybsBEL6Yz8QLshkzUCVI0NO9699388H7YtlyPUvBvWvQiH6/yg517F1
V/Dnm3lqwD7YNtxY0WpypHGCLT125AY5DOborcCOUy/5d+l2GpMGQPtwhNmdj2Wb
1pfdx3VMtCSUydzCXpGQh6OZXpcc6l/nj2e/St00SB0ja38IdN13pnWkxygytgDv
9l3xYJAidq5bvv8EFPrMOklLrglUUTpbBIZin9kQQtIM7cEK9kGV27PbH6Yf5Ywf
0TlWMNg6LY9LFiKTVzEd1YnkoZSE7vGqK7Hr+ihH+dZIxq6fRksBYEMsDl+B0Bu0
DBrR4tbyBP23TDpoA1nmiIXJWULuK/h3FOBSR2AhhXwh/iAqSYMDGdQfeFF20Kmx
R1Ewt4iw/jOmy9LEt8tVemBA9GrBAClqITsODPQM6Lvf3gxkCvkJZi0G8QbB8Q0q
Xx24l3UOdDkSNYYEQPMq7K30rY8YNS/27FGEaXE3mUiwpgVWnMllp66rPwQLb9vP
q6b9G/lNTfca5ghW+/2yOIRJ6oEkbmPIIBjGN6Rp9z8yONLhxtINKSAiQNTFobRW
gCohtk7jkXIRq9/yFBwVNwDM+4HAJvNx8SVzje5MdTwS60ubgYFjQ+gaJzuny2Di
qVp2Jhj7LIm6vg7j0njMeGc55IER2tqmqk2+Jxtqxbqc8N726OIRAWWmMKw5h78X
uLTJsDmJ6Qd618iDYiblvN0IH5uBVirKk6vHI/jayJ2RqIbcQeelWA3hOxRjajyJ
wjbsTbkEtakFwIzFW6KwRBNY3Befd35GU08nnVoERlLQ4K1FBUvH1w2LdD6DGF/Y
9ksxjYZT41fEDbBmppGSr+lUwiuuSDeN+G/mJyDU43nQtpuvP6c2S3LRzmCy8UOz
zOyyzZHXpdjd+3WeKY7v2aBh97cyr9eh3gEty0hFleOLkhn0DXFgWPRWH8fwExpS
B/4+T1k1sXnHtVOTRMvWIycu7anNzB8305slQBw/KHX0MAk5Shm1pdaX51JvwBTN
bm1jBmypg8r4GPBTlSilFhbv3AIi3KK4c5CLcQ74lIPwWzL41+039mJCJ6nhtvn1
c1jnVVmt14cpzZPrF6maLSpfQrVSlJlQU09jc9z+hyE8fH8+1NDxi1HrWqTJltBk
b2SAw+MElG8+TMo/LkoiRnfLXpFym98EOSkDKSMVZ49zAYLdSDpTJw4MAGfPwZh3
TVCJqnD7aJNbbDGvhWfU0g/ZqZhn81d609IMmWitm/ODrhIb1DP2PArVQgTf5sYU
FyAW6uHMUcs/jDJriazEPt0ewItvHhWb+HrXrSW9LAU02yJECXPHzofm4o0KNkvd
nJq4zw2lkaAMK9bJzDrKD2thBnRu66I/MQKBfqLz22xoG/5bpgVMtrnZGLnsVrOx
C1+o6UgrVCxbKkhKtNP6Vdybt6AtWMmUUdkps/ehhoRLsqTn27KGxAnZwzKKZ4bj
8nWhSlPg3WVBijjeehZovWmNgklg6isGZ0QQL6LlxmdhaFg622blGg+LK7rhGVTA
M7k5vVwdRcxL1pgsg5e9Ci22uOQc1omGXQUOy5IGg+hMONoTWvj/yuiqEsJXvYvk
aTohzzRAlX6OTHokr+Jmfu7rL0RRNXuPtrzaLA36RMwzXAFBqOJTOSPlA/1vfVho
Z0TbLNZ5rw2nxUBVQomEm/YIwGbsKBgby7JMtgGCehXPQoD/9LrXoJQKuCvwQ2KI
Dc3UzWM0eGCXoFmhWyq3eJQV1oqIKDJo4Qt3otQwHgeUfnxfKn1LOR4AVjkJOTMU
9TSzxU7D+myMmp+zCaJib/Eji7Cfm3gihqNCHWNX73N/cKitd5VtjLbt/26n66Hn
IUFBH5OnXK8NSAehYGJcfq0ZliqKxRgnSAxsS90RRamHfbdMHySb4sI0Yln2EhlT
n5DEHsGUkaEiUuX4gV2doHngcBoP8Ec6GNFXXJDSzb7G7CkiLC8PJAFUE1HCZ8zP
2bUedkxXjuRrRHmibslZ7S/VuDBFVeSyn+o/DE9c9jgtrePG0tMnG7O7ynmsICtK
3+3t/dkdsNebIXc2zpremMt/FS+fHJACyImkO5WICPw5mF5Z8N4kv9aHtCmJAfmw
CKTTwCfjQUzvHF645fZZZeyzht4vORZNc1617kRRToTRLb0u6MJM9+zfc24HNOMA
9h8cEdTFKseBMD/rzsSSXtQZzzCCyZQ5bnZl7uFexW4mINr8Xae6vI7wOq88FPZH
8U0oHxhYYEZ7AQUUdMIJtK/xKJQYMVUIqAPEdXwd4qJYjmx2E4KSFmEBVy+ipO0T
pg9zFQk4ZSQd1a5EfGrGizeOrxwWxdkfKf8op1e5mWjAD0zgIRYI0EOxJcYpqf96
BAnexzV7b+No+a/dv7y9F1IrcLksI3/uip7jD3AER3cdJAeOf7HvMId3hOc0UqTG
EKgfSt8ElWoOqZ5DQ6yA1bElohyntaw9Ft56LcsGNtV7k7Jxyf98e3UXIq0loQ5D
9suCN4vLs3a5HLkMPGBF5SOnnnMnAuUOOsUIeq0DOCsvMNn2Kgp1+Qh4Ps/U9y8X
oi/HM5AsxD9JK/GRWQwxW5ZGEeN/ushWYiM+WPaM/INYTvpBtMd6SnKkG72BJwMW
rRC3/zNOCRzIWIgGyI8eX0+0fgRLSDAzAfLAYc0qBxhNtRgBRMqPX2KPCgX/gkWD
yzHAyuN7W3Z9SDvOQMAeaSezjVpZMq9fgfSqF1lQeHZEiSTJJoaxwLUG3m7x+JZM
FjMnK7GSiT6GxMim84Ppu0wFZpLOiUcElfzZh3U9EGsChfKfqOTgZGoF7C8xL1rH
BbAVs0vpuCWXuWRER4am6HIZ3hJyvmtXKi/i+zpWqURPTU/2dQWpWaO2ETpOvRbt
4tqHXD920/4aF/sN46+yD1GVIp7Pckk8iFVBwjiLATCwThTyDKPMR4F/z65MQGG+
p5x+Sz6d7ssTXfRoRpwVWoupwdefRbFb2Nhiryhtvl/lj9qZCMoP2/e+mgcBDD9+
jfJ/QnFtdg7Frk8HTDZPPK7QHy/5G4L0euHJi+xdsRss+ScN0+gDEeXat0w6SWSS
9oOv3f5SOVF4CfuS+fImAFhp9KW7ZOmhQUC4aO0g6y7REL/nN08y48EmMrAYe8hH
uhXNGu0CJaDbEWhyGcYawc2CsvE09uAU0K3kv2mLza14Taj797h06eAt1i25Z1t0
LVu7y0xciqbtIgFdntFuh6BidWRyi+YPh9ehHK8qODpWKXicCqqbPLr0NPOCT2+6
RQkeyX7YDOhcPvzc9UTa+LNh+k+tkRWxUYQSaJXWcKxUz8D5CFgvedBwem7SB6qz
bnd7fcvtNC6kevtmEC7tzPuepNCu2TroUs5qa3E1T529qcOvCyUBB1wvUHMe7M/I
nDD7ZMXlcF29gqMsMLbKSIx35PNX6fa+9SgEXzb4hobeuYXftqN3yXq1eYExW0+f
9wGkvzbj40xEaR/EvwG7EZQIEtTYJeKX39kVObXUMecgPPn66Q0Rw/RlLSjelp9J
9wFkUT+Vdr0OtTrxFeTpklyLYP1JAc+CyZFu45WACRqI4dDNAjzXWbUl9ojBI9PF
HNxj5Q47Mg+rhiZDWePnZqEK+k7740mWO6YQB7qpwBsrQk3EWkIm3gp9SKWuk2xn
y1c4Da4Dd6sG+eqGSmg8KCnMqR0p8CfZeX1fLutYhynVIyUQph6srlldVr3jDuE7
OsAOGc7ThU1z/1qrnXsbQepux9gHQGOVCJfYSdB7Xks8L3gvFW09CVkBrNwDOcTz
Np6zQNm2WUYAJ4V9HfTq3BjsnaJcX6xf+nVSZaXjdb4EYqQKbL3TdgiNgwcaF5l1
YFIapVwAZum4Y34A64ohbErMf+Y3PSf29lecDLt13WLTORIR9PixL0RWrazfkYn1
Yv3h9TNibx/pOaJImfXszmLzn9TQINq69RmoKE/cv0beHOOSO1Cm5YZP2/+xkfrD
h4AVZ/IV0FZu72iZw5AeMrXeNZgFo657zRmSSHEYMgNKmciOKx7wp8Qt+PrflTCe
dDB4SkDvkpJe764faAaM3Kxxvt7+A9OYM4twBIsThgtt7+0li4LPT+bOSl0JySe3
MaC4ZBOyr1SQqO83Zez/KEe4iEgRtONG3aCQTDlJZr36ZTvhVktcLcKUaeIVypuk
d51LpolWxvaEEnGQHmgNlx0jMn/v8IV7dVhJj3RodZGCgtlaoY13enj0UiZJPeVB
wunrhmn0PpsuDRcYz7jktMUPUCt3mdzVz5Aastw4LKlIRIlonjdD9+SowUkM7d8D
wPLJ3Ap1SHYSVhJROXzRJWNnwxpTdNTgNFxgS/CloPpvcj+xfMmxtExEytzzIZOO
snsFDdD9MuOW5XDfcr9nBNOvvCk/P420myAwSh1yVjG08RORLSvCqI2GcpR6lgs0
GolO4RBeWSGGyFglQ6DUHpn5uReQpapc5HZ40qTRt9Hlii4yHGdqCj5vnef2OWY6
F2oNH//IuuaQ8Z3SrQBWxzHwCsBJdTrpKolevoQSaUn7rp0q+dEpm254t8kghwfU
FOUDK+u5D+vjiKa/NPZU9InzH8iGiD051A75WGnozlF/Vm/4pQ2RSwiH79n3Uz+m
doYIxICxA9AyHQ/Vt9Q0i9W7YchMwqACo595jdcC++6rXOEKMb7Rux78iBmKXoqQ
C75q8k+pB0FduUdev73gbbbeFf6DwGny/Jahi/CBzymCtYFlFdM8U/UnlWpfojtu
4so7Llt6GCdS8b/FHUbL5E6RLXLFB9ZBDoW8RiTyQt6ZMkFLvmTyTLfFzmmVqNKm
1m3muP1O9/PfEMJrBclTHQH6O8lxM66kBkLvB6SyEg0m6plpAmFclAvxy8uyuq/z
dxnPHU7aAd0W2MlSDarBE1gIyElHb+b05OsDE4LW8Zg5xVjZmGQODO3peIjFTo8N
u/pgyPqBwquL6iWZmZi8AV3qVuY32VP+nnWueqUOgukJNwCUgrdvRZsZbnmO8VMx
BkuA/T5zrIL/xn3X0XsuTAlYDxq6UcP6kcP8tn6273JidD+2at/xqu51XMPkVC1L
VJ5Io3MOvwurgGT8Y3dhEtJveAOtGC8FJJpsZl8BRTQqhL1sYYjxvV/Qd19tSY4s
ktQUwhMi/DjrB0PUjdWDyjmYcZQmraAPkgSL+RiAvFkqByjv5VK7ifcnW/KMc8BS
NGu9fq9l8JPJ9i5qGH+YccCKOdqzuA5wSEAkD7ZVufTWHkbxpuh5fxg57zW6SiIv
Nnt7Hosg1JFr+it6awDwxgm6AZsZB7fjFVyU6fVjFAN5hxj5201NUVU2MoyAIB6Y
MDdDsTNq7AXsvIKh1XiTZeyz3t24mOUiIa9dVk0FBDQbvHFJoDu36TFnS41oNwp3
hhD21WE7itbtqE+wyduVlP+MQxTt8HWZFYK/NUaNeyh/xsuiMa99bEpTpowOWdg2
mvJvlkvQenTua+Llo2Z0B8/tNvnQeJnqyhJRFq+aqtMmEZIOSXCJVH1RGRBH+X0h
Bxcfk9+259mgqjqS2M9EeoonqcMfKFwXxk/dVn6k8S5b/87K1BBAMWGqdj+fTegX
vmieVrte6/WOfJ4XMjcDAsBFXt+bHStLbulecF6dZiEbNP7Iiqatl+0e5B12DptJ
pIeH9qZQfip65QdkeAxY5vlU4e8GrFVVKXnlhPZfWBjKZbGou6cDyX1nc9IdnWfh
0OiJXB6A4apMw8fthZvai4w6TLnHH6RxdVAxMGmBz97yyrGsTkfznGRVZoKGW4Qk
E61bN197KaiVOVPrEHGSIjZ5VrPFXi8dzqa9E5OU4Gc0LBFtmV1iy2JE9ILsAbDp
OJrukwrV413jrESLLQMMjuncFWmP0PMFvUomjpi+4mk1xJp3uTZDr1FBAxWymQho
IAnwQ3ePS7ncJKacafMUqurzVzmL0UB5edCFhrv2g85MORgXwykvUMJwlhvx22o6
20tnIAwVsw2ZmRbQyyuN6OGEVMBpQcuDgZ6tOD4gS46H+5bvLSIwrd1HRYKMV4dG
DmGaD9RhGnVqadLUY8MceqqKMnPQT9GflJD8QB5bwt/y72UX1L2MlIq0+gk20mrS
x2n/XZgOsBWimBPF6uMgYkD1/mWn+Z8x5ZhjZZRbtLDjmdntUl/fVzEnGwCzRmMy
e5Lx//NGWdhYlGLBUHqp7LXrxSMWm++ScGV5kgqaML7w5KtJdCgBZ+H2Pl7rnaBn
GvU2Ba4Kc2/XhvCO0Re51xN3ZTF6lEzefZDKFy9VCS3kjzZxeFCB/QaUwDj9oMnn
uIK3/Ghj54MuxHaLzMH77CcQQ7+4WjBHS/5n/NNCh1XOyOwggugEvLRBKkmhlCnE
2Y/iyNQ5FdyR9VA92iR8Up0Eh75IgGKYaYd2u8EaLdPwM5neE4VYEFL0UtONI91q
5dNQhIHU+cpelNiJ0f6AcA/zl04tHAPEdEkhZlTZCoUUCz8UXA9bm0+N9WJgxewj
kiI9fTZna8WV/n9EYy0woUrl5SIL+woVUBQD5IHQaiAMWCrL1R3AENusiiC1v0Dx
22ZLI1PU9DEc+G7uityCRikDBWwkUDE2iKtwCp49NoyB6HohF1DG8vfLSWRBEQ3z
xv9tku0Ost7zP+5sU1xeYnFLsx0X4fH4Iy2pri65ptpNMN8d8NyqEcadgI34K1lo
+FsaBXFASTnXq8/qfiZKtPAM4tc8L8WmsBBpF3koHTZsMZTFV/khnGvyhgUpC3dU
9W4ky8MvkbduGjPHbbUH8BnNg5me/+beY51em+RYiIjzlos+cZKE80nB+hAExkK+
Hm57KI9onVrWvLk8VTWz9EXcwhbQAk54xltucGVsP7EopA433p5zaT7ug4SNek5e
knRkFWMVPvV2V7LnYOq6Mxa1JzbXtZsTXHv0dYVuyXjP8HVrxA4uRxIk2AqIKa7g
wUUgFezABm4vFsWj9B6wML8jTtBGvndNYpRc1/Ov6xAwERv3rkz2jQSsVDZu+hfG
KhrzXIDMjKiGEnPGO1TYEjosr4Yyup/y5lSf/Hp5VdDmdanx6UUL7BKSsoqq4VeJ
BVF9JRwo5r5FWp0sz93xpFOsgViI4CtyXHAEex3jiTY7CnVzsgT4WMH8j5TAnfta
oLgA68X/fJhJioqOEqbS8mFiXhD88RDQnMjVmZDqCW8CiXt7BUnICuHweIWH68dS
6ZdyKzbNAtStrVoLg2QUvWREeFnKwWOCli2Ta1oyRhNjSwqslwXFra7Gz4LWg2vy
kPRDK1pToDq+6XaHf99B6FKpOgUFmfXzMlkvMkdhDuI7QMcuEBr8dbCV5OQeQOk+
jAwgxSXTJ4xMs+aSE/qxdmQQaozNpGi6hA2BtphGNQP1iypdFjABJCZ9zAs+dMVn
x1IQnt3dGMHusjDUnMe6EXlgx3dZQHaVStgFEGkWnIlSbSGhxltgPRkvh4UILYuB
JaKGaSzSXcrXZwzY4Atm2d9u4R88PGlwcyzdkqGl9th6tKW+zsPhtd2FxiRk5MGI
SmSJqOsPCc8A+lX7Q1JmlT8HWCZjBU4n6KVde7Vn4c/v9v2stj8F2j5SaqCcOMC6
elXCj05A0vhv/nnQD28YzEIcaC8jgSJJYX/athDiSJFzSksRaMbiA+DTf0LAJP0n
rOJDEWrEGFHir2mIDq3FQVE3l73ltiQnWEfWsns1UUJI8M++GciBJfUsjnNjX/dO
UcW+IYID8i6SASUfdH6Rgh2DPjZlklUzjs782EYoA1jEOgfozVkYLvp+h8nV9iB+
/gSNHHj+a4KJSe/wzzYNM3hPnD5jWVvAzynoVgJZXcvwG+KFV5OyNLJdUnuknVEU
1aEKGlum+QHcJK4ysVwjGpdNrEbp9zbfGLEHjrnlcz7nQ6MjXe4PZgFzmJxIHC85
jC6BXedfFHs2dfreDGVvn9Rf7kH49/jsWEColbmw97muw0+DlxhNCBi/CcPvyNEI
rCuOLyNnwzuTFeDEWXW2HhYQPWiWAPHYA+HU4TxnHMSZrpNJkJSwPeZa/w02Hf95
WdZc2EJhNpI4YvQah09+nSrPOZ57/c2JWST1uNJtMElIY6QMU5IkrlnewNR3UW5g
NBMHkJqWAayksZwroOCRZ4/duPoAT5uAt1jwqdy8hjDgA54cEJLFI/+O5+nJ7XIK
EK9HqHMHaSS4aIc1SDYZBI67IQKNsUfrRINtY64Ai9mo5dRaKW91s5+rgaJUP9Tw
mJfS/vJT5MzIkbcX2yMxU7mxeANZo4W8lI66cqmEipXXxwqIjB8Cmzs8I1DtMnpK
kkl+njOJq9S9HqNX9IRbzC/EtVAlo0DXIZoOS/s0WPUfrdSq7Tgs+hZV60+1bgD/
eaVIs0zT8tMMMuAbiOS2Dir2fcq00lVsWl8V56/ROiLhDcDdQEz3WfkY39sC2qW3
h7QSf5RgmYnHJuyNVF6Ws+xq30CasTQxDQd+lW2wY3PBrYif/pxTt9nWRmHufaKy
b/uWCficYnFv2EKlgL5Lmxr1H+lDRzkrfi8O8hcjnEcTMSjmzlpFErPorbFcguXO
rVUXFuVXDM63EKihDL6r/wOoLq1F6GJ4XYQ9eF7xodBXTm4MafvjcskDU6Y5Rdov
VucE+2QeWq51zZGnHmyNDgiHefv46/xYfgRu4AnyDwjnlkgiV+qA1oTj0i2nKF1y
axAMBAP1PhICh6ueb8QVw74K8E9CpXOScvB0R/FhPPJjpSrak3NwDpdUsU4nP/vP
v6q/GtapOdKZFe7cKr5/KoivtJiUPZWQRrwbUYgPLOz3pJiMUo9fCCy2kuWd7bSG
nhEvR59Brk1mT3XPQn9pag==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
XzI8avv5E4dtEzlQ7FAZPfyYghD8jLTJwMxJLxxg0ChaD6eGP09iCvp1TjHaqqwm
I0NtWOE910kFUFCp3bcDxvp2YsUDVNAaovrtibm5vfRgOvTVI3eO7rxQyTkHp6eS
xaSwVTIbX4cBsbNkkwgQIXVJBk5CB18QtdyS1szzhp4Uo7/NF3dDHmmENH74Rjrx
WC7afBtaWjKWw826z+s9B/NNyq2voIXCAcsAPMTGxskXahKgN0RaFvX4QTaSK0yl
uQJSUigSsxpCe2AcNddednIXKpbfk1Op5cE5S3aoxhR6tiAuPPHRRCfqqCpPet3K
+Vs1zTZYyLHAZYmhE98fLA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 29120 )
`pragma protect data_block
v3NI82WLDRngesFXVfzp/czXHQQP5B63fHe5mEsMHHug1eDtwpBGv8Pau1ntFl89
Sfh+4zdJ/TEDGXGBph3kYt55FKYTnI/IJezUREflz/2OO2qPpdSAha2UDFAGngaM
fGz3UWNdU1awK5kgRhOnQhc9xWx5mHDRymmzJzRp2t9lKfWBGSXCxjKWhT3PVlBj
O9N4++OoVITdlFTsygmQX9aZRlSKtXQt6BG5I+yQATeNnyRD2hI9wL9IKWflZmi+
XVhgJQSS5WHsPfjxWBCIZjQ9IwYEjj1mDT/s/mhw/UkXe5IlHIW44tGcN/nEMUy2
+LNSa/rbiqctrgZmeoPmGVEquDxHcWgC98m61A3p5CYf2MWzghNvzfmp7sTu+oiQ
+rwhH8VqEWva7hZqkMRRgLa0anIyl1AYC3cYmO+32WazNPuARJ8SKvjnpy1tKG4l
GlLOLTUJ4jGV2aVMXLYkzssJrTgVSFLZKEl0boDm7F++EwWCKKauLOfKzR6upHWZ
fljpuHLmAyuHR4/voEcKmutb9bu9nacUAwvyjOtqX4njlKmYnSGE4yntzc9285cC
Zf091ZeDfErtodXywiA8FOVHA50Xbl48aZv3+PqNJhyp1znPlwtishfQ/CJaEPj3
s3tuALVMoMXtQB6ry5SsEAFL+5nVABY0+7fAIo9NF5Ysh49DZORAaXGHfTmClUqc
Q8FqxsXd5Vx+wOgfQpFqgmp/vWx6t4DVUC2AbxHDYOVx8966jkLEwS+JyYBcWR8S
LKvhDChmICnmdZma9cCSQun1EvbXlLPwKdHE3EVxs08Jw1l8TAsMRtgex5JooXiK
+Z90wqYSylvxWuIE0SuPKxFGSr8rFbOn8473O4prHdia/k4erJ5bVcOXKN4zzmgq
lpn0RjvYiE1j9dMtbu10nZKqZ2jf/U2C+OCXCfXPx5D7nCkyj53gXXDyl4TkRDg6
hc36TChtf2xwhW7b9TQjGh3BOlJs2ofINNYx9Yd9gz0HmRLa64uunIFtJ7yMpAJj
WGWwzsEh5+6vQPS9XvDUwXqXlAyz2CzH+E2UaTPNja4J190O2/EkfIuL05veMyaB
3ZZwE33fAtdroXudxnSPkBOhCfPk77XM5NOvBKehkYLXqKPSi/S52MxGgqtRyXPF
XSHbXOJWR5TaWGOVFrhKAOCQV+5wH6ToKcaSTvIAQsomXoQW+NoGvuDOKXV78lIf
bzuoaWEm/5HTB2r2zw4nJ2VY6rzwUQvuZJ8Ewmo2CZCQkoyLTGDFWt5XTuTl8akf
ZX8KEr3tEZkUfPQHkvmUfT2CtT+XLrmujZZ34l1aFlKHeRNdgavHr9YrA0RYL+Qb
QE/GTrVcVvp6nu6TxZBF9+77DGuYHMKXSJPXb2cpYfxcE/SUTx0aVI2Zgq+rn94q
ky/0BhO0qUVDmINodmgAeSD3WoTSMvQSmS7NNrbWIDugom/tRXEr5VZ4czgaOdOw
b4k9+U/xuGj0voNwJTI02iT/uu2cZ9e9CJLqQbJjBq4K4VN8t1ww+ypiT/ufAoCI
PIDdplsWRKaEPffAjDllfdwY277z5nvxeoR5xikY3qanc1kCe7uLBeH8gqOy/PwT
RCdV3XvtD/cyWJva93SQ76L0DTitU+Gf3n5FyUUrXSZ+iYxjwsjsNizWkPcVhQG8
rmJQuFZePghM/8CuIFlJvj6hXiRFlQwoRYlCw27FeaHNQS7M2tK8E7ewH51Bifl0
NRlTt3tYmpuQOmWSV4BFiOuL5gHcJmk0RjSspblPg6ltiBgYf74AVPMEHHke6orl
hBGLHPfzVOaN1HRxEPldI9FG89V8GgsnWHirxNBRVJM0QNlanfF9ZqfxuZLz+xVb
T6NsdXbTFj4fmSGLjrzFQlQDVCWoiVvv/tvMUsjeQeEN30ypLvk0bE/o5aUg9ZL4
NCkaUKCJlc/HI5bJzJsLhb6tiPqn2JLeZquA4nI6sK41gRlQDuJSU4LmmZ6VUF3b
5Ls9kHLySJf4L9stPNEp7ktwFz+TO+7h71dnjfyL0XpJPTRmvOJDp82FJ4nSWyDm
rU7zqqRQIQ22TinY6f/5LZ4stziTjivxKRUBMdCqf+aDOIaQ3CQjnpHUFMuJXC52
fRTkZ0s0er+yTymcgG5EtUivTIAhjVOh+YN+e71M880iDpVuf5yZd60gqCXTlHqG
7P/g4NetUpYgUTmg75jBXuNE3YmrXRulmTgW3rWnhFjV2unYhPT66KKnOkySTsaS
svrJ4stRiftV5XaGJH/Qy3gWcbnr/RUx8EDlLX8qKRXThrmyVXq0OjIVLoZmFsUK
u1hfUfIsatzJn/93GdGdSYajAZtuhDXrr3jS9wRl4uNZNd9lhfXfx6rHi2jhrhjn
tt1D25KbTcOxLIh5xR3Hj5MKX4Qw8eP15IUC1qKZ6RtZHNw+W++O7q5RxHtV9vDp
CT9vm5fsQxXFx+r8Y9FQM/Yg2wpXHpiaxTsCh2r8pwal8L4ZsGr4Ammr2TDkGl7s
ZIilalZql1WD1ragq9MSCxL3tiS94G1Eb+9MNZOuJ7SHBmfCTgLmMuTN+iKPbdFx
gzIR8zMAeEpveAh1dBgkqUhNU2rMuYMfxWrII8o0m4b+yshhnGso2SLnQK3wTqlB
XK26kWy6t/UoZB1swRu3gdRfxGH26LAQXF0yVNu4HisS79hKHPsnCjG7MSeZA6Lq
21bG43ox91nLJwu8nQmq205gQCxnflU489LG+VYvWLXMoXJj7CzsJJa/UjPH77cu
Y0H0ucLuQ+Kco4niyTEO6yXJLr51WvBT1YUxOe4NOu1PplbsYBBTsB0Hi8i+WFmf
NOx1PY7wA6YjdyFoRbRffBsDhVap/mgb+fXSDStiJ6+qCwINwnyOT1jt2LLW1xuh
sXdnHbZfVaP38lGEHUMeRxSfcOFxoqrJhJMQkQZC7DU2eZc0yZLV9HvWE5i7brxr
QEWoQmOn9qhUCjPuWSS4ayEsR7lATSsDZi/dO+YhvcC2E4vP8w8b9wyEcPB7Bv+n
A5qN0FezTjbsKj/75mx83i3xbz2OqJso6EIQ2OkAtlOdcm2zXK6drpV+0v98rmRT
2m51WHh9YKuGeHOffUFaw0TzuURSsu9L/XtyP4ond6oR3ZRWks33DEKVeRAo0OZf
V9YZawbdrC4KV0FkP83P9AMmjN0UNx2ksFTAgnY/Kf3VfibxgE2sUva2tfZ6px01
HYWlAR1J6o478xnitWLpmBvgQ0c5euND1hCn6lra78HHxIfhPZvXR+Tc3kgXYmm3
n4yWXPCCia/h5Pg49kveWrt0o5VcwozoDioVOPJpUX04fZ5PRixuXsaT+YcFUP5D
vCV8UU5WPbxizphSfdUxbfpcYamkV3KreZUPkVkCd6CmNKmNpwfgOJRLbjgEd14H
tJYQHDOqAsOscjJ+4RB/s+LAcp8Z36QfZedLFYXnreBLIAIyaLzQr/VG0+0r+3Dy
bUuGw4xkO0IN4Cw1zmYJLSII2Wd/KAuQD3AMRZhcHtj6uzo1/HJXyRGwIIIqDkdw
ylvnoutCMNvYQIds56cC/zgdl6q7yxIYqCEcZrRQsZr1OwQYZgEfB6D8xmk72tHG
YzNXMW1yRej4x7XlWdKG9FfLnWe8cohSOORwB8v2H2x3APmwGKrqWI0hibVNc1K/
jIwJe5tBbPO9K4quxYxLaFSDfsmRDBmQ9MKfxvKP6X4bPSP974HrPqZ2nt2sk6qu
VEviDQk4dDOs6hMC2sA3GS0ccBlLTdmoSX+o5yCdjF9g2hWG0diDCTCVRJIQdt/b
mGeO3z1++8hmMXR+diZQpxWmYwyKn8X/9jTyoZWVvU6Kkia+iTD4ihzR4usyJCzD
AuWefoMe6IbnIsRSmZOXw3fIkientfEHVUOYTEiJa24dJmSkf8WOMsrB75QscB7Q
RkXP5GQv//JWLJTBFj7GIIcF3f6i4kIwEuVfH8uz8+UqyauEEe4vy5/T1AstpAL5
r54lgARH4Cmku07aJFF6rYy474NUoY2cKD5w0dnchX1T7CVpCWYi9l4AxpWsajDS
1k4uyuJOzyDj3opZyBe1qCfewHMtBCgo1w28rSu25HYsG0enc76N0gYeGz2iTWHl
2t9J0hSUdpE2YCH/JOSWBe/IQlHn7lo/J6uUYu+Cd0gTvOyjAm05Fp+eVZy8sdRR
piuYVKzAXXY5yjPc2iNVF41RN9HQ3F8FBd0XDoVtsImV+HaKlYWVUUvIMbuDh73A
5DB0CU5HU9AwpXoWreuZAC50KEwJ2uvNQP8hOQj/o8/CltzE595pKaH0ifZkYxqu
xeFin2kEW3zwe/YELiHJeInSwCGm5TYSGMIeKDCjZwZrLolAz1GHsgC5WG0+WUQ/
bjkKgDJasmYdRxJ3LkCWtZHM2qby1jWyEvi5f99tOo8QB3taaHNFRRzyepnljJgV
D6kWxFkCZiCLFXT7tCGvDMotWYN/0FTof4PdNJj1qGs4nnvXhNI2ViCq5JB4Fvuk
mM6mOXjV0bjEdLI6n7gzWaKtIoAOad//8QN1SryRK0q3QfsC91FsIkBZbtq2Gg8w
qTjvDs2qSFcr1YvUaXwxVQCUg2xkJ//034V9hVo3PW17CfMjC9trgs7TOXYDqBGS
rqI4Zb6o/JBv4x6HmeDTI/X79kw3WElwYcs4GRo6IW8xALzuZ++Sd4IhYXdbGUhp
DQ/2S00ng1uu0kQChImkDjUX99dQKB0eOCmpyAJWXeLopKI5W9MGo1zRp8+O6UzF
Iwm532dbGDQsX54ufzXZ2lafePdXTUpd+oGaefny1f2XdKB37o5KAkyqACVOapwl
sMhK0124mEclaIUo+pDG7uV0vBTyxx0t/QtOKKLT7/CPPe7vFf7hV1iZu3NvSfVc
herF5YjE0irBblPHBsvvDPKSuJvb6POQNxtq15zsdv3YH0ruc2yO5ObuJ4Ba5Ffq
PQ9m7V8XBP+4r1n9zXaSmGI5D7wkiPiEO4vTzS0TlDwTtG1w27JVcszHMxxuEjoN
oSwKTT7pTXrMrAEUTaEk76dKyl4Ok413tCsuAx1c0OKkHzkigDgUq/b91DyWxiTT
+64adGlTwJ9Kx+qMdwjb/vDdTRBX17rfdUTqW98HeWLzm8VTQ0wCqVayQU/0r/5p
LdNdKEoPuiZ4yQbgi0sexBaEdCkqod/JEZshS0BShUVHlfMArFw71mQS/+Y/zf4P
AEkHFrJg0hWJu007/3+2HyGjj1/E+YH7GU5lgMLmJhEVgnqXa9ft+DqM9TJ69bZg
Etn3ITDPyz6ZWx7PlzkccNmMOEr6fdB8DOv+Pj3DTK9KQCYFs6eRitnNOd+oopO1
TpYJScRQsQ8ikgDb2mPv9JmSRxdvwkrv0d6bipVSRJGPhW8fadP7ATMbHiCsdnev
CCSrVNeBkOPetSJHitnxlg+x0M7aflDPqi1/xywYwNCTNhQ6i/Y+lW9Uwu2wfQnU
TsDY7Kjb130FM6X0H8rbj23RXUUtJbJQiuPj7KvOFHLvk/nwz6pHvUnoSOSPFHN8
PFHSDKwxys8DvozhHTzkBmRdIgpOscRc58cOo1aHnarmmwYvVYzI1PpWy9F+gMax
lLP5ky1uT1DL7SENYKGeO993HPlFJY8asTGXq5GExnaqRVSnc2UJ66vjh2DfOinc
CZb9Bq/mNAjVuLU5yjNED7XYlvTpFZ9vkeg0vBi4CUQOFBL30T+UK3yT4gwX6K2B
j5yKXxEtKCo5iErD7LmIuoBbUrb9XuJDeOABaf1UeAZmtjelZuYuKEjdSSTKvMPO
o/yKYPlXTfBttUuEI4IDGtVlBLhGYMPvjOc8rrSIiZsMG8SEbG1ihEDmi331FkGK
FAX9ETnCajRS0Lj7VJJBvTB5gKz3rfSpaa5B+o7O6rzAAs/NkELk0dVTSoPvz5Dr
t7gjJu2ztTC/ik5MWoSveYKNM9Eqo8tBiWxrEtPAvfCcegaBodMWEzN8VcoDpTNj
MoKAeKJVGLT8kMWOr5uwQ+rgem167m2HnGd/oauNi+axIrMqW1kQ2K/XJFFAP4ac
x12wZ+xnUSHyWDdh3OgqPlL3rivGmNO45GIDHu0o1p2S90oRu6jfpoBYrcQzDi5k
Hn6V4JXTb96x8JbVl9qqx24WNF6n4e642AFaCevtFWg4mAEFc8Bs9l6DJqzTGH+u
z5+/sIT4lBXWhYxe1RU9LCytDvQVuYuY6mpc1si5YxHejX8n/ny3zVV6ojPfILtx
cGmvpTvw6BiTPL1v7IXtS3xrc+6C/JcU0kwjkja7XLAa4BRptemkIqm8IkXDlZ1m
hL5lrUPRVUWelBJ2roPq5vGeG1TO2/BuDgdRbWnexER9VG2UeGpudsgUk2WCkQ3w
AQnTM8oojUv+j/ewgmwU9RgwWD+I/+xhhlPSFKqWCfXgpCIwbIC8WQ3k042PBw+h
QRt9NYW1XqEuVpMj48efuUWrWVwgBrrVSSETDZhOrwc9VkwQY1mY8Ma6MApjFyn9
t1fffJDULXvwCOWd79ZB6VAJheMK2L5oYMnhma2yRRtTqDF2ogZpRJqwGzjgfzga
O4CbdHxLX6cuvuFSNGQN9S2b+LoVUrSjfby9EwXbty2E/gO7XnXB0Phsd/xOpjP3
Ub863n5iDAbOZ89ze9oEcY+kU+/BPlPks7WpIO4AZJjOsMs//fjJ5u1cfuEcxkVr
faXnV5Ngwxbu8sI/ZJ6ZuNGBrasv7uqFm95/Pewp5erzBNJFRsh7v6NwdBIu7DMR
3ufCSPj14pN4paLazG06CwS7VRblmuttJCrTDQNFfkgrqSNPnNlpRbCM3UTaMv0f
0YMs7oEfK8pXgVEKQTsDL3e+mXITVao5Dnkw3TPorYEfYelirzN/4jYrUujovL4m
t9LCohoL5Kgwk7wPM7fWDwYLvo7DU5Do8mwAnMpDFQDkmlgcvNxB0+Byz2BH7/x7
JkMeALtzZZ8pYwAKjrLHeJx8OZ09AKbC5CcRxuKBFg+QB3FxmCsi1j61ISCtjAqc
cxuEyjGt1Tf0bOImZJsY5FO/HBV3yOuRzWLV5onF/vKlVWmcYF6lmmMMJUDdmcUg
vozf33yIXGiIJy8YlZy6/Jv4NOBFpFYYcK9bg+sToJAdx2tal9ExY/ukdp8K+ahp
py0voR8yNQGdRq15Ul3ok7r7zgR7PIf2O41iSyzKa8/WkhobtsINPRPbLK9gB322
hjk9svI27t+FuGBinBZr4iahxt8Hcy678heJXionIMrX75h/3ZYxcS8OWk9KkVMm
kwEuQ9QW8Qrj+k34qNyTGLD/K9v8c4Bp+3UI1X60Fjsn2LbRRJ0bGlJAMtSEMZNv
18ZAtr6OHKZ4hQm/3H+2yeLwXPHKrcNEp8JLjYt6TV+4kHL+XW975m+EcPrBLP+p
hYNMmMvsdVb244LNL9o6LWaWJKRkKgQAGelt2ufAhDQXTpOnpns08Tn/kY/CrGT6
23csgphZR6xOIzqRmTkY7gNIG72ZZLlwfc5I0SSDHJkR03fKbVCvlqVtjgtxEtUU
vVIIL6HauDEk11HcVEzFxzvvje57c439IRKn6lf7K1hpRiBSuQrMRqwjwdYUEoyD
juEh/Tk/f4yoe/4JkPqU0wsu9kUKEuhpI5dvHkvgO9qYlPadhZd1Bk6NaPRI3Rff
laCMw7deNe51DWBXhFHTHaFnCvha+kqA/Dd7hioFFp59J2tyPM3OyC8BJbfkFdsh
vunCXIsDbUyYWVucMtjxYBV3zXM+JqcJtIjtv2fKNisfURQ6LdSGpM3+hNElwZQ+
lZ/03x9aFVEF9RrZPVDKaHAb8CcBoAlOFDVhK2Hiep32/NQWvJYyD3IFsG0c4HtQ
SBSKlp/HD34oUP/OhSr50tt3jclMpkOkRuuosMOXmbEsYnz3jBBTpRihlmsRpWO4
FqAZMwseYCoLXtdiCpas7MeQdB87ij3+L2LgsVw61imL2FkpEQ+wFOnApiC/ip4n
nkurePl8pmKuphi52BEk2EI3uqqL35PKjrpoU9Uh5pZUOsB9LGzp2VWpAd0/SIMc
qNmBVIE9E4R4WkSJabA5yIgRSFpPQ9JXDM4PMjFzRli9by5RQAO8yUoWYE2dZTK0
CduJTcL3kBX4A0dmnmZzGwSA3JoivM8suwhvFs5F2ArXC4C9/ObCjQvyEQw4JLmR
pLvRav25wmooHj3qUXMjetc108pbvsXK79BohGuTfpBViSf9pagoA3ERsl7bjs7a
jxwE9qVuxsGjju16xiWq/RUUabZdcbB16AMuhfImqDBlh/uMsoqSlVsG8MV5QnA4
oZeY0GQPrkVnz2MvR4KGGCo/xep4HcSAJA8hRM2qXEHURttq8I/CMkjEJ/skkbvW
hXwZ/hsZ0jCc+2VNHoqxmH9VinvAgPKc0h1Qv5W+fkyd9d1oKYzySZng/zVhU9HR
kEW4LAJmPiZmRuW2Xa0xdF0GNP/ETgV1w9UWRfz8oP5Br0cq3ZrS3791XTCPAK/q
mJ1KJF1h3HAZb+sUG1PDk29rx86ux1m9dM0CeOmwSeFxQbgsddai/N8uU8MBzzpo
yG7uiQTSqaCe/kyYDnWb1ZNRnP5DE6R8UiyohOiXWBtqaxAxTmVsY2cWpG+WKGAe
TLqzM0hXzCa6EeNoT5rhPPigzk+gYm4TqQu+FKJREq1ah1EmAVnZ1Wpp1LmpaOJR
HK2mveg34zqc+5iRBidYZDsKAHN32+33fXG6f7VTuvs8wZCOWhICIaRzE020CeZ6
xBvdHcTmKUHi6p0QWqKsg9DWtzFpYaPkUoIOUW+1oBvRDOkqckRRbgGv7jK0IoDB
Pd+5nUP3EHRem7QbVQLglVXVN0vEtFFQJsJXxs3tTThO85/N/58YemKFxO6YqQcr
tudfxP3Npe5SPh2T0RMUG7lQQ0fvjDCAIjnWeg6g/J/1pXGwabFfFfuUXVYNCgBU
hLWj4fWlySWdpqHjXDgfQRa+I1WNZyqN5Pk5ZjRo5KuXLMh8BKuxFaPTz0+0f7hh
KlepcSJVSzkAbEZE1AxIN03qk3dA7ehpVXm9O3pzh4xeMKu2yUubZBix1iClKSe9
E/4inJKZCTILxKEAyHiQETQcGn5IGP0fG+JdGh7LYvSXLXetQjZ39+FvBEd1bS6/
ymRJIdlvc50zxSH1PQYrf/u3CDql4G9xEt0Gt7gCfwG4u047zLvLu6HJ8RLaaWug
LzvZyLgbvEbXOVIY2xVREfk7lLpdZs8VFhOHbIKFumS8CpsvP6NtQxGrIibkg6Bi
XC7f+3jt08qkq2ZAPFi6RyU5UAd1V+OOoL9MAV8SUzHCc69tzlamtKFiULPLhhri
BMPgM+3q5XvElmJTYkojpCaS58kX0ICvokeVkccgggmlgPrm2BlsaUvWHMxNLjmT
+Auv7lCvH4TaauuE3s3xObzXhxTRx31jPZzI5TLD0YnCVWfwB03DZN12HvBCE2Vh
5ItAX+RTbwL8hd3q+VVYNlRhKWd2qRco/+1MLCeUIWNeYDIN543sZtjilfLXumdK
LikPIjbOjarcNxTIS/zQG9axQdOKxKWDkV6ukwXzKxZOdX4+sT+P4YYTcH2Iwm+z
WLvdbGDMnC2A9yEbgc4e7lJ061EvJRn8ywhKS6RUcp2nfRhwDhqRK9TlavOPQMQ/
V/RhpPCmVI7G73hpHGVNjdnD6B0o+jw1bNFCU2aIBXkjNlr/yoFW+tnRK519cYhb
tVQEee3cmdEjevvgZHtnzJVBM5vvtZNLVgNkHoKrUZ+Ee5u9Cd7D6WF0fYBI9xW4
5AFzHr+1qwvCvPHpiQWdeZcXwFalc88NAgzfEkGR3iOyf/VP//sc8Z7Z+oDG13Pr
4CrCZpk1BH0DfICn310zVCdBjEi0xUk3NjS5Fkm3P1nM7cR7NMpeZ0qBf3WJkQHD
idQkj60u/3/+PvzSxKAFES2AJhMS5GhM4/oEUATN3hvvBRDlsOf2M1fqXrzw7uq6
lCkUtZRSHKQ60OrBGJ9nYtL8/k576V++SK3VOqeoB7olJyQ/Te1CyZJihUnlOXDT
2D6EKd+Lfq0LKdS9FNOXGkFgncCP82L+3RwkLu9Bzg3ty1T+eVN4lD6FVpQB4WiR
b3n7qiYbE/XdnQA5JfDxfeeo6I4dnfhGCSD4piXMmKJY4NLYekP/swy1fsUrOZsj
/yPzyHtKX6DEFIvfY3hft6MbFmjs26cMbfhpI+aRWbE14t4AJStuQ4mHjskWnMeL
5QMtGiO+dBSswSMckCbCy9fqJlmi1Vhaos4kMzymSKPZ3RcBTIB8djGmoWHAu5Ci
Km/wIk9UgF1dlREbzZYXJ6M9Q4HXDYlalmQBUZBGHFr2mhkmTi/hpliSYYWPzYPC
2pq9AdlJSBbB8UuEgYK3y1MBjT5LzzIjjXI0w2tVDRjDT7AjpxrQjRxy/He+A3jp
TWZcm9HswYFNCVID21T4KQOCrdhfbt/aLIp7XatJkF+hTwm7T0A1ggGz3WaF5QIk
GDWSpV3TC1s7P/9CxdnYGcNMtMcwcT0g0DOFgWFRvh9WigkKN6lttG20Jz9TTdJX
3BWWMwRegcCPbpfsznsgT+9xCkwqGwfUtyVUk/S4aXa/HnVPVGbvCdYmuKk4s/es
1d95JSOgVI/vY6tCNGgMRvKWMldnfx/ow5UW8jFOMRNvpu5GjtT4no1EfgFJYfhp
0+HWlMy3WomHT8kTu0MrzDMCg3L35BBSyx6jMw1qswAers3nev6ZSLIkVCh0J8sL
/UhmqsobursbgQQ18BZrGA8YGVuLW8D1MxLgz6YW2eaOOTeDSzHYM/Bcfj9YU1we
hmUDFEkGi16gkqfU7KcuQ5rzvvMQtjoniay+Yb5HATD7sVFHQcPF8kwJD7673tL4
Easu7TQwmlDmOX34EIibXiDYNsgXRnmJVUgUFqWuigdqhWEY7swJtLd42vETP5R6
HP9vJ48Z5BNz+0ahr64prOFXT4FjSZPQav7tOsl6DoeQS2et0Jim3cklnywO/VDO
CKYkn/cb83oin1oByRJOpdQqzfx2LVqwUp1JA5ZoCwACRfU9flX0EhALEPPZLGUA
ZOA9syjudGE9Bs2rfTVAsD/gL/G+ekLfMGLvgOnn86KSmL5dQQ8DuajLVTpurueo
cXmHUgdqUUy7ckvmOif1CtQD6VRDeZdR2Jf6+G/BgJdK4V03d2FomP2i9hdjnDff
/4r6pmcfRa0m00uWItoJaBd2Lu2EVEyeconkg0K5x2OWqCls3+Cs7O/SOA1lz1xz
kUNIqY5diYTAIwOx6VatmLe4SFPv6vBtq8OYeTE5f4wHMvB1ku7J+qEN0Pdm9257
1M0awioVEx/9XQPxrfwDWBfe0m7Irflr+gHRfZn7pkRGMt0Bb71Lu8ht7HkBNIzl
5ODc5FKL20CpZ1ECXw8++Rx9KEIHvvNFsKxHI4rsNfVzPECZ8oiyUwwTiAwxB3GT
LKgxHUnxeEWKUXfbwctnkOQ7g8Mskpf7t2zHYu65e6dlWnRu46lnA0j+HhsCVMTM
re/aqkgG3QbSFcXOpP1TlFqTLZQYHlcUYgO70yaOHtm9IfVaYM7mKYW2VfNPIsdI
HdnjrYTFicG2o61Kd0XDjAZWZXu/NAupAws7/7JuyEE10waAY4agBS5soOwLR26P
xITzj2auJI4T5BZELA8u3hhMcHk2KYve/94mThWRM3ckX4siepAgbyVsHTeDwuzn
87LShTOcO/X2rhH5yl0uxl7NOAnajA7z42O4Z8MH5N+crWNOdJxmdFthPXCiNbXY
hpRjwG4hT705qTiz3LRtp5qZQBaGyzlP+lu+/JqUsK8MlwEuinNsNr8yxbjpzirF
TYnrUN5KrJJOhnnrt/OHtB28C7MHA6Wl9TzZ5MhqtjxIG0cMXmFgEUZZnCQA8Y46
W3zuXzs23wqMMMJu5tKX+MJfHBZPNXUpyQPrLFAI7Rwiem0HEkO8FdPvPckP7DXN
hq8z/bINjMHTAa70GRvIy3JBUAP6rDtstlPDjQFlUSa80ZSOMRuDoZQwOwOYyn6a
w48Y1uYaeJvnOHj6IKqJW7AtkS0XIT+nwOOjhwI71U/ewPDGZnzTxrzo3/tCBrW8
XIkDwe2D7pC3hm/fHPtZwzmfgqYvMEWkq9AOncS5EJx4L3HA/OCjh3QY9usABF90
EsW3vqmp1W6wtArRwPlksdn/TJmdarKL37S6S9spLO/TFIW9ETZQbOlKVuaRiJpb
ifib4EuAdtYo4Esh3cpccNs1MdiDNQa2/l8RtZC5zuJj1tLOnNyfCCjsmVXlgYPe
ihL13Bvtvyohqs3U4D2rytHyQgTQvj9/7Hciqylmhj3No+tSoH0UtKQ6B8QBTRW4
LxXbgo7ndYOmnBBVaYIM0RV8es8JMzNuBywmr2hZLZu/iSW2MMaJjwpXFBIsxtel
8qQvvSlYV5EZ4dcXUICcc5flHn/aLP3KUUbGwxDBDurLJTwWrGiRUEMVLS9fXJ7w
AOIK/tFV8IkuFF4DIGkSvtYQV+nXL656pL7/1+1yWh9tlqfFwE/B9c45rEunbGRC
kS+rqFquT6j+woJ9koZ5Jvm4Fq3VCHSbOLesBhBsosPqEv3RA3YeHh+RtT/ZviJm
WL1HFESFnJ4apBD9qLhgqAdGXSVjRim1EGVmWOMhY4vWLmNv5sTQMlXEtGlPJHSm
7zaC14zPk8CFj+I+/88WAE+Gp5CZczM87TJ6Vb+55ujBeblEVCPsCxjEQ84wfJPX
NnzVpWMAii5TUcylL0IGjojM1NecjtXR6rQdsHH1fVmU979NQx/hFZvoXBy9j4/4
qhRyL5WauY325zX8vFKP1GN1edxrwedZc4kvXs54/7X9QjDPVcK73x0LbXLVFSMk
OMBj05k99NbtP+YMb3MZIQPqI2Yx3btp29B4BoBbZwq7KackIe7V25iZUgSc9J9t
8uHphj1WOUhiHCt7BoNLAfZIhj3iCm9MoPNeyjjXvQzKx+PvI3s4et+rPcwQPc3X
oMznAgJ1KIHlJSDNj/uDFy3j8MqqjrHzu1P+MtQrx41IaRSbZN7eQmqB1UPBYcPl
bziGZhvyPRbyYu2nvT2SYRt0wGU9ctXgL066I3JI4Fqoir+monUhpAVqGsvY2u35
xKlhRnyzBn0b4TExxhxEiCwdC2WJKQq/M+If9it6KfMiMYgCtbUN7QXu2YWgTucz
H7PHE819y+0iXpucXOvYgX5M1UXw8x32/Qxa4y6eWZqAnguaUotRMgl+b1Wc5cis
28KlDF6ZDjX4/9fzc4yUxP1xwKKvKicvPLqETmSArrmPmltWPVvWFhs3N7Z27KQO
VG5aHP1i0Ao3yAcjYLRGaX+/zSGEZIfnXMGA++U/PsiEwLIdOKGVL8MUprMXqeJV
gL22VZscQ7DDcpiwJQhj8tPvnak6xF1NC1arUbsiDJhbAlrDkWj7R81bORRBe1h8
XpBEI3MnX/BfSKp8GXw/H1PMp22g8pK4tf9OdGOMxfHsPcAvbbAjeXado10nLuOD
DQFtBnRHfYJl4FR5nKuO1ica5fJs1o7Sv9XIg5xEsrKyObP28cJJNjgozDMtHQ1F
UXhUwMbJPApB6lpS7rvUa+7eRET4eHVqlZmQPCgdrayJnBOsMi/J99WMffPdF58q
5wlGVGCzZD/3wpXKzacP88q25pINJ7JHbTRYXjAx5m5TCu0JVy4aNegdu2oGq6UP
i4/z6Pdx3lGMOt+m5WlhA4s5GbWY3GRW78OjYWsLmsiR4OcK8+8B0Kxsws5OEXHv
3pVBSGprKpDricPIoQLoFH4E0tDrWOOLW1KXLRk4bHzjf1uft7uFiopQO8ZTW5JE
Vg16NISvzdGhZ4Bm5x5kjT1Fqf2H7F06HGNGVdw4kifN3ZOSucvnjyNxyTpgNQOM
f+L6Tzc6D6iHPKMoaIqrZ6AilMBVAOsDPcUTwiM+qDnaH65RbeZNw6t4Hl9kps1S
YJHkVwXHtQbgOsvJJmYUibAGSXzs+3e2phQDMBYnT550tiCm7NlG6A5R3e765Hk9
0snwGwiUHMIwciv74snOrzzIZvIRbUh5fhBmX4Lqx/gazFK6/utOBc5ifIp80JjR
2CYMb3VYqbB/UUvA6fLmONxdL4yGlf5tVXZRaTO4MzQPp/O/r3kionzet5WwqBXI
F2s6wnv81lJSOOSJgitjLs0wa57a8/BJkQ6h6fAgdqHwmQWLpc3uy8sAo26/uoFr
hc6XEvSUXJhpp5Pf40DgLocKPUOMZx7WXUiYCOxOsD3dPP2HmGNN5ght0SNjd2so
X3ZZwXkSxWu6yhDEbmErwsQvZ0MMmtBZTWsoa/xD5azn5CdDvYCMHcCwB19N5HOX
7s6AupylaWvK+qYNE7oYmIA3yVdhTlOJi+pFfK09peVDoa/Zxgxl0SvLVw3kaB00
ay4B9wh2xKAvOhxWMtetF/hHJ4DuZkmY/lttUHGsqQ24iP3FasR9PXeNCFTWvaGY
+oEFyC14Xb6+4YhD8w8MX/GCj/Jw5Vq/zdb0SnCOvTYZ1s/N0jlHc0/B7DLkMhJu
aSwU3ypCmaBc3/mC4T9k1y1pM2TSwquwuyHgPTGpDN8HoPd1PEAF3A/RtLIHiOdX
fpZasMgIUBoFm56I/8r+oIGSqAEOpNaMEdbDGhhQ7Z94+orW5klMyEiKPe3x3dRy
3aVPVrNumFhp1ihAhi3ZGnbppRPNVHYCmsRAXeUT5xsN3etDW86HtUQotk/mjyZ0
xA4yy59A4cTYSSZ9WIb29aXZkMvBDUpe31CZxhUYmKZkbFf1JXr6PsjKURXAt1vo
ZVLHQTI8Wu3TV+yZnuPqfFfFrRs81jXhGRfaEEqsKVm8YuEppoaUZZJbGWdfWgdu
DEFW2eYjnyPdWSS3li/TOiAmcUnJvxUK/3Mc7QU/9H8dycvWHiE+rX+wVnHw0Z3g
yitDxEDV+jFA/XTn/Ic+Jzz9zUAEpJMgQs5TrKElqM+Col4ogGG7hhF0mH4pkeho
pH6ixO2qLHzlPMtOYGToykoQWFEuXtatVh1wANgEhBFzx0hYgTsKZ+2K2JVs21TZ
9lIT/Lw8hELA7Dkto7k704mZvFnOKlOotrWh2oCGYRNLzoqjOA7+wW2rzKdUHHSQ
B8ZhX3nT2gcSTPw9VRoEZdJ5wpRwIQGK90KZPp8O/GjQDXAt0qSyLzk5xd+N0AMS
rnBDnWpxNtKoURS9+hAf8qBPTe+Lh4TlOd4glPJj+iiTG5dbYJDIzwmww0DnBG7i
uPAGcIZhVHHZWlX8HtVxfAvIAiJFJ/NgX/nPJkPRdSH+8wZr2PexAFVbCXcxlCG5
Ic5PfwceLSjZ+qKjvSNeRcWiNHBDrF4fKVXiAqiARpoaWxl3qiG+06P1GUzbf6pz
XJq3viul4eFsObiWV37d3wIEUWeGjwg7Ax+GcQ86GZa/AkcZNJh3cjgfr+eZJQzr
2CDSRzxbloyccy0oOJleSl2oHZTFQuOwjHPumeoY6QbS9UwujfGzXzis/HTZLHSY
5Kmkxe3JBwLztPkrB+XG9G/O+ayzSxjOk7KcunHgp703tYIkpipaJaXuNzhv0P/k
xbIJdAuFf4drVE/It/g6ilNmMDKHEhPHXaMuNRZJFyQDPM33XQuTUh7dIBQC+IcN
4kTcbi9PplFsahNmSFOlc/ANwwX4XlpYOcWHhR2NBjhqnHWlwlSk/kRWpqSfoOTb
ndVO+zkIgZ//POv1yT59WkXJFcpldTOqJWTpcaNYHpP8l4zk9iIKEDMkf0ZLYjPY
uNSYkCgKooFRv7IvRfOCDZs0WE6mpLhn5a6bjTxe8kOzeLQzKknQPArrcqUWRZLy
HpRfWztz7GohCZCHYRk6fWzpe8lO7gS2FykY0pY+2M8aF8vWRciw1mhX691Yo07v
LfcjZpCBubItgQbhamObrQY8nqzuUrAbUSJHIoLK67TGcLAdui0MolUvz0gZ7VFF
fGHPtwH026yTRjja5oYdZm7El2r+JUscq3GUXBH5iwOpVJkTtAaCS3AS2ZCFtAGS
I513A7prdGKI/QU92B0UVJGCF3PreA/ii0vtaXIqzz91pZyhY7wHK/kd6GW9EJDB
ShkewHRwHiiVyE3TP7jWXkD7/fHFkyaiq4rcEveVnW7fJT0BVu8B05hstQjrYlV/
YaoxRc9oSmEf9WLQ/svCHN+tEx0+OCTfHTzdXKgXDsNxrprsrUpxV2FH6ndjxfUX
wGnN3DW1HpM3tJ/P89EQZ2EyOGFkLR4hZB9oklxc33+EDPRNMELnB1/nTnvUT98W
SRWA7u84VltkNKr3fHgPFbVBeYKGtlHy9bByfcXhUy8U59S8l/rQ+XNKqVnx55iW
vTU9wIGcx4czSgBoGGNZVXcCj4hYYcfgFJ0gEC7DCF01iEx6Rrc3kWqxTOUy/7ym
t3MCFXW/IZ7uiwKYHclbNGRj92MClYdVXABpG6xvZMaMeJgUHEHCPQ/s/+aBY+xN
UYsY08viq+c4xfLFkDrFwNo31roQZbkTIwDYGLTvk2f0dHWPWaXj26befW4v6iAw
s5K4Ud/8FyuRuULTip40FG5iLgXQ4XTGCu4n4V7o9pDO2v3djKnQmE0dzACc5PNc
I7ZQGzdmRe5+pZejEU3ATvFtiZPmA81IsJMQEptvbF9qRlYhhP8BdsEt8yAeBZ3n
DVn/v/U9xX3CovQZz7oX44RNLyqej9aVbWtiC1fgWg3UFi2PofIE1Svijn6oaqYp
yh79Sq8KfbN3b8nCW5PWO9+iNVUfpXNqSzF1DepuCBLJ998thx/b7vW3G0NbHVMn
nfA/SkC6XnE/nxo2I1XprRiT6TkgieCItjhjJVkVlMNtJH+b4afXMPosry2aUsb3
QqVq6rDzwBy2vKR+vZwjtzLY2vPvTY11ELV0GQtKzruOsN4Cu7Hz6+jzT+1E6jz4
ebnlzHRRaXtz6lydHykvj/EgxkmLsDWhCGG2l4Tyb3FqypyjIY2Xb78g7sb+NWY+
LZWMpk2Qb1h0c6XhsjidjjJmT2MgVyjbLNtCh/Oxa95HhNuxXPP0f+2H+BA0UAkQ
oGWajqbIoZ3j1Ilxe3OAPvTEuHIQrgRZ9fnxpws5D5LPiAkTNstTnbqtlSDLCYXY
/KD/9U963l7wHalCDdIe0HC2WL454ZtbxCA+O58irtWAddyMhvbR+ruml4YGqrDv
q1bUfpzlv+QjdSw3pbYPbZyPHJVFBnlH5E3FYH50u8RuIIqIKjK48TN5lmDGqpnV
cprltkNzHvjx2+dbuHqW6YanA/FtUEIlrKF+nXB08hUbdH4zSqqnvaudLpKGcYqY
B310gTnFg/ngLbFPjpm9SCxnnjZnKnsKQVmVsdYrhdtfNfvdGw/shjxdTepQfKHH
UbMy0mjdMQNzbfRBmqtMYHATfv3MFlhqcZUfzK2E0TegVuGqiZRjlMMN4AU7+eqQ
tC/lMIIWz9ws3SYrayD6WSTuZL3w0gLfAvcaKLBkXuPRcU2Yps6oOOJY/yT3cX6p
Jp4IpTBUQ/b9rEcVzM3pFK7vEiovawL2ncESEHfzTrRWH8HcmAi7uqw1h6B676od
PsiBaH0JXIvrtFsdnmduK+VqoSxvNrwRzs3/xG54HYMOYCBR93UCLrFtuS5yCuK7
fssgTdXc449+HAvJqmIbeCgVOyRw9Og2Pt+zCVXR4YPtYG702PQXrmBoi/aPYanx
1bTbOLH3iY/juQzF5elotar4hQrTyehsBzA9h2FG4n8PHhlaEdDOoFaBx1tC0sN7
p1V715OSZWDCcTDnfkh2ItDbTXSb/jY1Kjv7tLww/K6XeE535Hn42RH4yIHMH8wb
P6UYbYqqoUg43n72PIFs0FjTZQ/CwEQzMVwggNVlXXdfpPDkbGvKN/fuBPh+YZP6
4hJEBVu3DE8kQ16R5eaY0mdnvpJdlttnTOyq1WtkRpivRHjplMZmKV3X4XUFWn5E
5oHC7y51eZODeo0k6B+scXWNzvoV5a8kyNNhnb497ZCy9Vj1/4lA+TtrwEHa5bpP
sq916dYyPZZ5L7pvK93vWPiOG/XTDTygDBEH8strQ6mEvTDwAMWivT7utoT57C1u
4Tz6xDZqpBppVHnK8o2pm8+ajCMKnlQSuRZtEGsb3azj1LLydG9OH2PmFEg3sjTQ
JM38U8xClzY2VhG2F9WSwmIvDkFx5acVZPXf03i1z9uqz83SA5RNtTnIdNuyVb+9
h5Ag7y1MNKP5mNzeAj4fZLc1lVbvNb93R3gvTCg/IWN54PEHLyC8SUgy4J8xp4Yw
XpsxWz2YVKaDoWa4mbeUg1Y5UW8TIsX92lqKYY1gcjzFxOeUwuY/BFZGR6F51zR4
KnsLwWZu4hS1YTRTP9XDZr2n+GwdgSHs6CyzJuzVnPvHMf0w6cDQ3ZMyiZP6YWJF
IW9MyQFk0c2B6TG3LzllHp3Lh0DBHg1EtPDoevEuNK0Be+p/xSRTawoMCS8hF8lV
EI8FIlGMEJkBIswXIsWRY2amtSaT/zXVvA8nSlrHxxLjwqXurvAcIeXAdJSSYlUe
EOkaQPWtuY7AJ2GIMEaUQ3dd7Yxx+2lASFkv/sb2dspdWofBUIWZOG1NeceS0OSg
0LjmcmUY9s/wr0WbGXrUQAY1eHSSGDNtt2C54UafvVao5gF5IgwZqdSfqBdVpVxq
M75qDQIHL3AJ/Mcv9Ohl5GNxoUImdGR2w1OCpHPj25zJsb6HJup/hnePzVrpBIJ3
MEa71RKk2yxW6gtmI4MHrnWEopRf751tIZkOdN2/DnCJ3P4dhd9nuII0WVWwWUMz
6Kws8X3KRBKjO5rEV1OaQCcd6T3qMVpwcM8i4sc3Pi7a2d8MnIccgRHlqIh5Gjko
AqTAV7/Wo30bxxWKTvZFrObfOkkwUssA2HYX8A2Imj+kjQX+oTkKuvosSDlE8g0k
Rz8Gxkgg/m7yt0NH64t8QgkV9mcBxjtERgqcCWNmC++IrbMBohYMONfJCn2GSOWa
PtxfF7v5miD0LKIvBfi7nlUbtSSOKdRazAwiac40/r2r8Ty8RkY6OuLRyrw20aAt
YwtSU9FvzvNX4OwgBeYzOU2OZjX+478BdvH/04Z0fNNNkSXV4rQlU1VN0eJU3XvC
rymkBqWV8F29H2IpaE11G9btrTehCyQgSVcnvD/CrMFvCsEeVKPB/TPDLwnDBawP
EOGaNTs7aA7m7mjangUvjO5H1lBgdmwhcsHEuZjmwximyXpWYgd4/6JMy0aLkx8J
+xsjG4yi0IEIqLapFE4Ps+Yvt+E9Mbh9SQ9HvE9K3mihy6dTB2MHvxKov6klPs/m
6Ht2sgWMuamyZZOXRwlc51zc2Ob+Q3OkrByyChs4Nkqv7rAawfUu+xzI3WaW8+dK
CvFCZlOh/FPxd3Ujph4eff5RA28Kc8Hiweb18c5CTDgymdaOz47GhVoKwMBnimS0
j5sE1YZyhphO2xswK4kUQRwyJImLs+aB88ld0jiX1HZvkBIIPzNVCWWHs/siqJEQ
VnQWbuIZ4QvcjFLoVGH2OAavfOu0PMoxdYJbodlgIajtNhrIQQZ6GaD/LDcmZoUe
BGw8GPn146KTUpUVcHtvQTsBJ++v3krjUX1A2PFI2tTSkKnMRG/d9tf/Axrr1+vm
zBOP5ZbLJwTE3hR1/wUXSGn6tMEqcU6vg3k/vwFoGFAKb4wOcssrTkNqWHMIsRho
Zxl9x+rTb55kyQGYKTxB5slTFuiCUPAn0uQIfu3rmVaCJD6pzFSRwLOxM6/9oIHx
kJvxPZu4zOfqYUHGkmGwZF5shYosud0oJlY07qoykVP//LfI2O00aKiqPo5q0sa6
u4LOM3auHzDS0QihOpZE1ac18Uv1WiGQUO6oYbRmmdcsYq5ucc9w+xMxRy+jl+jl
mOrfdufe13F2Rwz8yvBEZuzheXZnkKMDgUw4KtCEGPeoC1XbSt75CwCIzPewN2q0
DS230SIiziWD5+xv7FnwSMeq5PsXyqq/yT2jeIiU0j/HSnqRVdfkrF3XGG6TW78T
oJnsxB8Q6lb5x9buRCGzNx180nHGQMNjZTgBuVkfsWPlbpQjxkzoNrsOhM0SBIQG
qyvpli/xheSYe1L4noL0k1+weFiMcKumtm47TleXetGBkIOiomtg66NWW9Z6toRb
KRDtsOYQBy5sELQfctgQBxm+SXoHmIxNFGKIR+J2iQoMXYM1keSCoFL/htLv5wO5
lWr8r1r6qe13l8KemNzzz17Wh353IF8CC4VNiFkoG8p/2wwCX/7S7L0BcYrQLFPl
bFKTIiylOVNpOC7GakG6fuU4edwPgwuSZqN3pgxebzdH8cB1wllL251zASlBo1Zv
uzJ+iOHfvlplUVGGjtImWdy79kmZX/qqT85niJR61jrZtmxxPrgA3+sOyStF5RWf
7j5tp2Y2hnkHYavfuCLFnZvTta+k1C3LH6Ap0T2v5zjXLvlYUJVJgrjpTYUEEinI
RvWMPl4wWG10spAFfYsTMTV3d1LRDF8Ze7ctBzUmrXhWe94FbxN1x4vElKIDPDPh
/+E+/wlZNuu9DUHZFuUhGtrm1WTKfAUGyMO1GBJVexTCzokmY08AyzsdN6hMhR4U
Z4WyddUNYozjFEOTomrhQnhV4BDFKIy+dyzDmPHXXPAL+G3TNqNKVmBV7252ZMJ+
oFRtO60cxWh6laWtkWDZKw5rmGMvVgtv4eBk68ENimG/8rSDB9pMQjzEtjmYvShR
QEY6pGBUTnJHkVYIFCqA84A115VYo1W8U+TIm5YsqlUwzM6480+n9FdCeLTy/Q3L
roXvu6wECJmaDfy4XjzO1USFF5deo0refZMjR6+C736Pe/MwG0DWssh5xSDm/DBo
jskg73Ogc3fQWnMl+EbuGrex4lr5DXCYbKpJCj5zTXwOnrGWFFQHKKb47fw3nokK
JT0EDiRAAxM1Pdq8/J3/z2pzGEaTni8xd8RXrZjJkya0WhfVB47jUew+QQcyqvCp
3AbncRikORukBO8UagjhaCnjOmkJAag1M737t+szkub1+cKX+6ZghKYI33y3r5Ob
+H8dKGtdj0f3BcgwKhjML+0XvRqQ9i6z8FpltSWfTphIFqXPrPicnncTrYP4h2zz
23OBUJd3TTTaIq5zvWl7KTm8u1PHTPpikcJQfJ+WP5wiir8rVkfB3v6M/f8PPTKA
qMOR4aOcqNtQoYm2StZUemoAKGDj7jXFLGjaIeD7odGlnW5YSJyzfD6MxSbW/Xe+
t4d7XD58XVUm2xeUz0T54NahOcLs13MvdTwfPLsiNTgLhwaxISXgwxBZCx7rNrib
2aBxhtiGKz8J4roM1gG7YBGjypzrJbYGAI1gE3EHxDviDYg0YhiPzcf4lYWTQJHg
qfZUEtdJLhPtXKtxm5EFGEk0xFVG/CagyVcgfIortCz9fVpARM22PFLMqyF6aLy5
BMV6k1Vm7liZAideMgn4R/KB6IkARSZHJy2uZiBZmdv7Q7rXqAAYGDKRsLBbxV2v
o2J5uDz8aG9zNy1s8WZH991g9zbaR6ba3gyiGB2YEeAx3aUn1Njgn7w0cL5I1Ctk
EGzuZTHavNv5VWbN0IFJ/aEMLLPAfL05ifjfgorZzqscMoeT7VFfe/kXujQkMHno
iOZLawrzFs050mRl4SfAi2C6SkEMFzIWy5ZVc1xa+WAESKfykm/DbIN5+s0ABGDw
lnDPbZweQbAE/wH5E3Wf/3YcZtlwj7zRL/7E//UqATSHU5N4B5YuaWEeZNVEBbn8
fMTac1w79m1/TBHiPiWjlfUFocLic3TL4+W3QHjCYYjsKpcxFtn5M/cNB1a6QV5L
vDxXPIixorr/56jU0L09hjc6vYts6mBwV5U3VbIrRl3lehw07yzggbjxeUFwyHdI
Vcx35pOa0wp0soH2jggMQhRFUsyBrubByvGLmAIoXC0Y3IvCqozo/aRqdlfX4VHc
M7Ot/ThKZ6BhERFrI1G6dU+WdgfR5OVnc5yjURpub8nGyo4Rordsa/DBJXvF3PfG
Tb3qmebzHuDV0eXZBGkbca4ogVQPX6Zm91xIkEh1fopQpFYgKCWSTt7cfrIOD9iD
WUVm+Lplo6FERP9hQUjxlIZvpecEGV3bBMPac1sxJVkbxaNh0XuZ2iMXulYOhFNu
PuYVY6lVqnMFC3QPnZRGvJY9IZJG6KyfCeN31LiCl0nDz47TPXlx/MqEosTdu7pN
jz3uM+knLXhYgZqDElDouqlUBo+pYsbr6fo9SvrA+XUAXG1M3TuobLzPV7FbJVaI
rHiteCttQxxYplgIRf9MF+Uy4AxboBOn7hpkq8Th3IdSRrO0yX2G5kvFdbJOLaUU
eoWRUXBo64zxH5CenPyfhH40SUwtTxcw+jHaHr8yJveLVITrDitvIg6DckNjg3sF
F6L55C/8hvephRQZPCFBcoY0saiNkW3RyJBJUf/MJa3/ClTE6cTimQBKpHkCTbwj
ct7/RpdwHPRR1lO7P259PnMLEJUVjAT+CuRqSY0mfmQks+5RumLifeKZSF000i4N
lPY4JQaocVGgP6BWeug3T7IB/cjZL8FbMjn30OZ3YCIoolRLsjw21V+q9HQFzye0
Z61q3nq5S0JjK3gZk9gn5texi2N/l6Bt5ks1J05FN+Fz18IjnDl2KMcr2ibfgD8J
P1R2pnLer9kMOca84z8APZyDV6jSZAJccJ1Ps4hWcQaXxokczvJm61qUsnNv0Br9
dhhHc/VHi4wj00hwouDjGZ4GgGdlhkLmOmuaJwN+fP1AoWyyZlZqExsWJx5xdYJ3
+gMrs+JUbI5qTxX4h1KgGdpxRbbw2VtMKauSSURpf513yHCscgpAmf1FTnurBvu8
0Bvx77PSPHc/MCKcharl9SvqR7AFxIQJ2CY3nIiJCVAuhuk/VOTWZoegnludiQg9
7xhf1ePruOgv/pDuSxG0Bz/ckL42Dpl/CUGL0fMQgLCWy0zxwT2uoCsQRIvs24LA
o7QOu+MkKdBO0494JtDIasRqd86oZLZGnnZKQ4T+qoluFzP+x8s6T7+CafvWNdfp
0ggf1XCD7RZrN0A8i4dndgfNqVZb54W+OSQa+13DENkWXiMnBp31lZV/AtcWnMBk
GJQEX1msmNoYci8gxf7CGMzxBNYERHeXb2DZAXcmS5V/wFr3v7y1L9OJShXsS+QC
jcXUDyzAOBv5UaAjoLPuR21DMIM9WHfuLUCu5QJIf5T/8sPKOr2XMCI+XTRy8Zf/
YIXzaW8PW6NTWpZSYtwy78SBSfleMSppri4gHuJ5mWAQINTwB3p3qXKoCztEyRyf
FUdxPkm0ExuyeSxtWmJbcSI0M1bzP4gHxEdIsT1vhMWstyaC7g7IoTnjJGJx5ZcF
K5dFkV0mJJDJ8WQKCq6qcvQHSpqc0JzIFRexREbySJtqG0gStCfn77GSHozcTSqk
7jXAtCEDRpiZnXGI5ugcGoAewz68DIBxnlXOnTuVg+tClqcluJIWiNaNEaI0xPh3
cHVJpWllf3eup/Z1CEEnyjG807r0i8wqeqY/e73Qtvbr9Z/zB9EnfHfdUBM1KoDI
6z2jrYJ+7KHAVZXsjwIk2L4Z+7QSz83pFq5W5ecaI546LpOh0JhByyJ7kHP58c4f
CqB+/ns7IzYOXqS+hvm5x/ur8fmb+SkJqzuGmBIF6xQuRu5H7r7Bm306oiWh58Jj
kBifZyIJ6sBAz+Z0vsx2BcU7bgPXc4cVjiBwos2DTusoz3nAu/9pmJwDf12pjw+s
Bq3WxmmqrBDNJMbhnCa24o+JOsZJ/U3+9qFwM7rpY0lsnHSFYpc6MrRjffaxATtz
+x9iYy9BzNdoInIFCKOTNV4r9VEIBJ43g12abrsg6bK9PlTPjf/ZOKfAUEBozfY9
CXl7PHRf7zKTCeHHs+0kBwY2GFTfs5FWXEcRFqmoWrt3MQLDmNGQX+pi+YQFPi9y
jwB7FEwMA8xGz5+7AlYvTyRcUEccAQU0REAG90sRjreH8hon2bg5lU5mB96ontX1
p3jTAJaEs1Vfn1nW2EwbLWKB80JkL4DrUKvkgWsyLBucO/+MvyhxSyTc1c/hkc0K
INdcEfzXudfs/ZfUGgFskQ0YtwIeoD8k20a4sMidQyh9v0ET5Cz9TnHSomKdW2Y0
7m/ekoKoI5DRajtmLHinT5r4iQVhjIpExm0tAaa7RR0czd/ffBeSlUeaYDW8AZbQ
bsEX/z2m2svEaKYq5B0O8KYLMNQqS7LzFc0bR0pnbMVQF6mrOO9gfopJSCdinEtK
qSafTzKpxICShHBtz1PzQesbDOTIjXe+iROo+oA4kRn9sh/RcQTJaAFVdcimy09o
cOt1eNjSp3gKcUv7JpM5e68SIFZtS6z2Vs1fE04xoToHxQwQjkAgZWQUJmnkU5aX
Svu9M8scZzsaUa+cNzeRG2vpra0Nq5vcwvvL52sAQfsYzRNDltXj414IlehU4k3d
QUo9vItIMRa5r5VIahIrDUUg+1cH5hCpUe01vNDyyECkVzfB+WbF2rBeIrYCuZTp
mgX42A3blw2lo3WSq5aJlaBGD+7nTp+BYtqNa5cC6A1EHNJG+GBcqYGSUzx+qKOP
v376DAkKZwz+ipvd0TcKQzxf0d1cK5rWj+vlMP+nwfjKppkqJg8YvSk7w0gwHzTL
P63zwoSeqG9qWaBUX76yztc4qRQAGqxm4/cuKAEIG2KblaJknMlEFeTHJyhnHW1g
XWYplO8p93oBiPzhw+NSaIf7k2RMfbFBc6E8myecggrY+ljcTVr0iHXeiqptxD/e
Xn9vjgiznnFwVPZ6cWBoMoUG47sTd5r9rCdl/5ZlAd3yvaFZmgjLYdxKjdjbTTGZ
tSTOsnCxotX8ixk1Z7+Qymmm+NGaJSO5kCHbaHR8ym1bRaBWjS6/OvDo1qXNjeMe
sM306GWHdqW/bLHAxNxHKjHVKL6uV/7wOaF8duJnJk7CXMKrKMhM6VYLtUWSZlFu
FqGEMOQJUyOHYBaEqrT/N8eJqFNvw3lidmhfivNlf4WpQkaFTsmrCE/PDodp8R1N
JBRHH44oPqq1paGVm+juY/GuOfY+9o620+drINLiHeKLQpZmulPkxgt82IROWfE0
5t2qhq1JooXCr/npCx/VdhZmxDd84h2bhHwzMhk5V0v3cxGacUditmbwRbK8qvGw
zc620SwVdkqrNhA28ryznFe8L6q5/cRtIVMVD2lacyV24mwNoI3aPn66waGa2dCC
r3yyVDd8ae0zIbuXIuiG98lTJ/YMpRDaayJ2914KkQG9bcyuU+I5A+RaE3nQuQS/
JbEgKI9mewtx4nhH1A5CZsyKPonVQLqIBYg1xM4XSLpZkpW7VWZAwD6vfAjuD1XC
gMpQMst9lRPirfq1RlHKpsw7xsZMp8Rr6qPtOSueOUnSBw8NZykB6D6AVbhvVvis
9bgzn22eKWHQiYQWNVT5tiETL6SVC4mhj1F3qxsQD7ErT1UJmwqWanU3nzO7c6gd
Wd1TaJhzfGkqLF/isR+LC9sdZWu+8qn5+0n5ComWfLzeVFOWJD3YnhCq2aUUPkoC
xhVYKs2J2uRWgLQnBDxK/ua6B3ahL46Sj/V9CE6XUtdp6duvrC+CgTFi8q0wlplc
D6bcaSAht2oWFZLsDNe56NtXNx7SQ5rIIwQDwH98hX+pKT48s7s1NjRkxkGNJ74p
69faYG1R1tuqScXP+AkxNbOY+CLwHlYf8WhbMlecYqW3Rx4g3TbfUzksSk8yfVTO
KRODZcwdFa5d0Agbbab516s1yoVqSN70MBY0ysHBAEV+uP55lP/qfqvy3mKMCzJP
ZG5cujk1RP8xp5NAJJprK+Okz0jq34js2fvkctwy+SLl0vV3Xjfqo+Jv373D8vyt
G4lr4ABC9F+0rjoWvmV+bTApF/umqH/LfpNwaRKFwcMzSMxErulGg6hlErxRGRl/
LpLjrEd8Wkx4QhNzGkR8gvyEGFNqe4/CblHMEXcpSNDV0rtf5ntHFcoNJvh6f9uA
ov/Dol8qB5MNpF61tRhEshn+OwHI5pt5CJrDJ6vaUldVXCWSjtBBhfarW4zzuiOv
8VYNC7Tkr043q1BfvYv9CUxRR9eSvs/kiKP0j+VhrvMj/Oz70hGgXpcZUqQzwzEZ
0DO9YgYKdlDsAmlIyWvd0f701Ta2iEyMhQQA4bgY9JCEIngtO4HAKatQMkw+A2pg
VMcA+qFlyFFxRy3cu1fFPWSIO5P2+5BHJT1oPK0oazftDWZTWnKAyAxN4q1f6Byy
ivixjTCT6BnanPbpkelpLht3jY5cNf6Fo0Tj2cIb/GN+7DKAXLp5DWpZMHdnf1VK
B9rwGPZAIdHraZBBnEvzwH/kkqb9KBWm1vcRE6F/JV1lYeDINsANJU/yy9sMbqH4
SG5N1msNgaLdUwxzHfm2O7RkTH6T9zuhPXPBtwXKSi/uB0HAEbY20rC+1guT/ikW
nZosapxaZkHNqpsONJCnPyh7KQWF6cUMZ34OIKRYAkywhlxlH1SGUA+/obXR8HcH
ZxBg22Nq2e4Zk2N4qi8RSzWOd2JoIHI8eDwJdlUs+cpsGGC7IqsIxGBHjnWfJ7Or
vFZ5UvM4kn8RUmWElkRHZ8yX8sJVKaf6W03TPQVcf6Td2gxI38j9nFP3D71DnNtT
0MVy694SHza5254uqNT5Lcl7gZEXJVJ6d3iFLqBcBQ3RH6I/ydC1/zaXZGAxNtNH
d9hm0fVS14fJBs+WjbyYWjBxuNiR3RmUfTbhs5wuBHk5GlUOG7q2/R7th3fpGXEf
ABe4DAUXcs2xXUYmDA42MYuB5ghOfPb+vU72mf2ZKFQz0Lw6yCQR6OBLD3fuNNts
PPJmeHC3fRK6rB15WrR9uKLsUtgFvcUUk28rrVgXOW/6YAgDYDHH8xCxTdZf4RkA
jVGAYwooJV6q9XTjnHLDr8hLrbwFp6/EZ9ssHOjuKohbDvuDywhiAuCRmDZnKjB5
cxycmTzJTMuf5H/3otWS8Mn7r5a23zU+7lABvraYX3SnDWZjg686RZAAH0AXa4Ib
mSnP+AEINHUFKQsw9wk4f2u6FtCynkY28W4seW36SbsdTxsqEo4O391B3BBzchvy
bS0bxJnCRZSribF+GDn1HYOEmScnDJNeOPv9JvdeggnaXpwAmPEWI+jgqT8gBhGF
ET1mU3ZS4KpA0Lhq8iqtpBNSi0mopWmoAae6kadAG3rD4kOS71kQyWXZIzdqXSD/
SdX/mVaqQfjEIbcpfqFErESqvBjp+nNi8dEO4dkuz2byNcweN8cSuTMsUrqrV2kb
n71J4KeP/R8w1TN/cSxKO7RMWQQLmOMdXGj+c8ySbnSWq1wXDx4npkj0QSgjfcK+
su74PojMey72W5TYPCNYJWsIJi0+To+X1HaWvXOHH+BzI4uQZM63LTpFpvu6AFtJ
aHR6jxq8QBUWcd4cxXsGFzXc8d2VSjbg7/rPYbCcTIJptnJ6D8/T/QgLPpOkWY64
q/+k7Rj/jX80CietRE/44gMnVQ6CNLHeHaLzRKY1HSgdXUPN1bmUsNQBXXtYYPC6
5VblnsfEbGChlk/LrL262cjHwOmb7MFxfFNSJn3NexA1SpPyqHQqv/K6TxXR91j8
rGkcfoT2zQrjT4DjftBkui3L7ERePb7e3L3Esl4Cfosff6eY8HtZ9GAeGiwbvxo9
Wh3WfRhtKdAy2va6lqZuJTH1orvwPhuM+OlFX2eWtPvxvA3H1Ggx+hg9e1U2yT4V
n0VbsGY3ee2TgbeS6jq5twaueltHGE6ndBQZ6ISKKQlPeDzQj83dWGVuLUTkNIhw
cbVnrtcJsMeAa01F2lsPVE7tWlsKQXVNVrBSS6mFn7ohS4Jq4j7iuERbEJ+ao2pG
9+YrSLaDe4gF1bw9FKidwdfGVDcKW/5+b8itBhWrcVFcSCooxjxK2Fa4TZGAG9Mn
QZYkoaef+mVKc8By6M4O4eIWK1qxiw/wGB7SHYjTG2JQQNuCFdDlTuR8dP3AIXj9
bbMkfytjUed7cenQmQw29R85Cl6WoVcaZlnnG6ektH9+XQkuLCcvswXHGo1wOtKj
Gd5JeCriZeWFY+ZymkeQLsJ3PSq370F9xSv2+9LNb2pUpf3aJe2xp1WZx8pGW5Fe
0f5k6Qwb8srp5Vy+ynlp5w49GbBpi0PnlMJRvS3ujg743rgLiKTW8j4MMBlivZc4
LTsD0dJVUO7V2jv9q9Tjk8Mj6UZX2ADgzietyRZgdN8/QpGwIQiYl204WnBtpLNo
Z5QdMOijF0Rwpwrxer8jm8HWaKV28WTu1QqsZhAU/V6hIokYHTcRHxGvN+PsMeZe
DtnpQOMtYAfr9yDaVDdIhl2wdTltBFgEbzAIfS8BFiuUa5pwjR//Vzz+UmyWhizg
fCgBRLx73U99n7yLpkHSqFi7Ra+X0/SjvBEnvLfQ5kpFyZiIWQfA7JryY1Utr4vY
s0AUwLLQqzvl6alPWdazkXl6wHzQmwLBN1FKDzfkZwaZ/gy1BPYTL8W/KE1DfSPH
rdrvySff1jD/N2MAfxxCnLNU6b5Ssoo8GadGyzN6kU62QUwYS8u3H/sumvwntj0T
iMhvvlUMj5yollMMm9DLZY4lhN5676IyKj+DpU1wyaqsLoZQk5MBK3d94qFX4nJH
qL1ZtZY2rzQWtT/4p+3DrvOrF0HBpPjUqq8kh9IECSsUAI9LtuKFceqKNrDDDCA6
VaeGzpGUz9Z31BpLhdC5sBW5xEo6cl5z9jrMezj9peDWsw57PWM50ffvR9CyO+qG
9A4ocVEqNrcJ7OSNxWOdYRQJbqZu79LuFXT7+vmnv+vzciTwiEHHbNf9kc2/9Z1M
u9GSXDzbbnrZrvqOriax4Ctqd+Z5y3Zh9XzPRsSQ2+NMAA5Xh8y9rwVXJqRXi3wd
22JThiE015fbueeUJ1nhJv4Ae4O6yl3exLjhuZqMgB3SEPomt5qpJaRJOL0+pAWF
RnRiDErv6LFDRSB6Ev28dRP9qp0kGd5HyKZmUkGt2S5kxxxX3/mMeLueajl/MbRG
Er00B5zhyL9ewfANCjPAKg3fecy1R1/Um/FEM/JCcTIaqoG3LhguBTPEsSoMxE9d
7dJ1oinRkpD04vasGVLmjs3eUTUaEQjzX2q+w68r3nffZtA4NfxmPG7HQlKDUpoI
UzmWJvjIf658JDaHNvEMoqtvq5q0BVZfBiea+hhLYvVesoIPsf+cwVU5SmUztdTL
MbS2B3r9DBuneZoIw2wi/OobX83ujp1b7yA8N+3lY2kwSU7PcRRyfMeXIBAAstxT
T7RvRndWo/uPAw1+PjSpx0UnIgbSBdvytHOfIvjDM1HukW1H3Sb/HBKF9bm+vOaC
o0s9X3Os1FF4nuGcIqWLZt6S79Shm6/Ywv5CbxCqmDyDevaGwCBcEA9cTCthl9aq
iVjhxH3lXeGnvGkUlZkxn8wRGpH875vkUN/L0WvaQwy5tRkLwjQu5G6equjOAtjR
BxgBGLY5tOHiJ/vtwTsJ8Tchk55mm4slrPRdjeauSDpNKzjKeFMpQ+pGR01JMYuv
8Amz0uteUu8ElpaEKfWKV3YNZH7e82i0APfyfYFpgK69wyHchBZ7RhQTwmKK1ttg
c2ywMsZ8z6nQ1jsy2MLMbHtqpGOk+XaDaVBUE3ehKiPTAQVwW+cz7yAL/XW9xAir
8mVhk7VZxmNRSkul2ZOq1iKrZD1sNwRw/YwkqArXvAUMx0NOYEvPpWcmdZ23INmz
Vn+e/Y44j473fs79KfidK0Bjq+lRCKV8DfBpL0VZBTPHwSM4batuyn0fQ9wQfSgy
HOGrdgDUhj7Fpj21Z9dLzQBqt1Eh1m9NYsg26xRopiNgxkNknBwWe64BenhbtgQz
7GF3OeGNsNE5S+R2WWvHAQ7iOxJOoHfNvZcS/nrtangQDZSRbGELNd7FI+DLrPxi
TsqkGynJlRO7Jnz2ayitEF22vh92GjLybtMuA9juBs11eUVQMnrsPq5A6K4Bmglp
TqFhR+TPXzSRZ7NXzfn43gDjBkYi7U3q9K/KaUvDS6Q5NVJWEZxfYL8B92HmNRNH
od4mf8Z+UGzgtC0k2x8onlzfc42ZM92vbSmGwJhMNU2JsxAMkAPbcd3xI5hHRz34
rKU57zhrP+AcA9rLcb+qVuccpA7Msw1qmx4d+2bDCFvBeC3VBtiMePpFFOsdpVA/
/eoGB4gEgsarkVBIxb1Sg2L+Wqgr4Lzpv08GbnLl7YaNwEGKi9hGTHMJHqea5dhb
hQjhoYFs8vamOtb2RE1RyvB6oBiAJjqVe/n/UNcA+IlN1GzD1bs+rot8aP51mbwi
/dQnuUKzO5S/JTXZQmftpfQjmrCgxU9LNZHJd+unZHOrRSxMPJFHDvHajP5vgqL1
MbKLp0EW/dLSP4O+GwRjD9WOfH433RZy0iaRV4qCFOArBdhseetyC8QdHJ/CxDaL
uuqtNjQkfPhVN6M6mMnN8olzPtN9F30l+eBdoV2ZTcREvBk29qt1dejuhfp9eYDq
O2FTY14cjFV3WCBC81AqdUsOJMNelylem+ZGk2ka3N4rTi42u3z0GZS8EzO9eZg8
RjeR5609BpVlfHGCLiqtqguyt0oEHSEt1EtVp47GQKgEKVb+iJwBTtPdltF705EO
Js8Bwbfn0Wa/eZZ5K9zoSMIbwDQHrygzCT8FLkXwaBymn2EJQ5ROaGX7ByFcYtQI
o3beXvztpY0C8oTuY5c4NE/lF8+nl+hrJ30xpnmarcB8/2YKIOafT/Zq3yaN0SFF
WNHsCqGbz3K+e2OuIcPvr5abK5+HbznN98DECu2FG9O2C21z/KRCb9tfqnVL3UJF
iYNump+u/m+qB03KSQYwld2WXUKxgkEBxPDdKypSgCVp69F+AN0jpr7/J5ovLndS
gxqpMtZqsG56hecJESxUYDcLEoi0t2lRiKv2mKTXnkjgJyatr7LZBPdKpB55Ayjm
QqEf3bhqLOJV41RTbBMzO1JokeURe+OQZX5u9QjlXTZMq0BR8eAufFv8RPSdwmHL
j5JHeoHCd+GB9zhM45iQfn7ZtvX37+8GoptkYtHtAbNHGsRfTJTzXBDfxDowd6km
rEk2miLn58ZyxaoRpSBRbjivyRzGcRtSTg53gud5UDpWrC01GC0JseAK60sVkuK1
ilUGSTiX5hNYhQG7yP+hh0BJBlHBef4f6EoA/EJyj3k2aGAVhL2eqR48pRhxVnzh
NrWSujzaRJSrKka9ZRXcfuRxTt465VCb20c1cttCw2taY7w9bkDqHfafNKbJIFrz
4n4vIrZAwm9IiiijULHbLz0R0SzMxrSL8WK5J9zfQw3aTcLRjib34Rn6VWn7D5os
2aKc+exL358z9kKLVBeSRydMZeXk5Dy9BPNU8A5dRIjItt+fjvNjlRto+YtQNX2f
xpRh4H8IOtCeHhLZG35ika9eN9nX+s4GQoxP+6Hq8WFYQs3E4FPdDmwMWW0OZowH
AaeZZIH5mEvOwevQ/EojB/9sC0ZXNjp1IBSOMsEtiYAh+nfblPEMRJJCjnmCh805
37ZanAIDNXWXG76L5yxVV1ea1o+tdSHVwoTpGift3YgxBQQtjMej3pdjpLUOAatr
+PsTcUlDX94jtMOfhtdNcHXJncTW1P+Czh+z1pn7WEmz1Jl9JqVFXhFTKtO9avs3
pTcldL+H0sReS9tEstfN63Gy8GtpTpQU9ig3iTzWxKS1HxYismHmrA6Sioe05otU
W74Jar6poSEJD6yOkYsyannVkm6+FgBtTNQIN/CcirKWjP8/Ny1nPjcCguxVpLxl
PgcYehyLhSAdypVAylVnBKS+LyzTD2zbpWu/Ybp+LDByOMqSozX8E79uZdCFUk7i
KNdX8JXf5I1nyoZ1SpFWOib1ua6yCzbz8WadQbUraLgQdzmUPIy9Qp+tc5BdTbDc
+R2xcj2f/Lq4TLyRiFs5qxe37NEmweVU5YfW2gzJH9hbnOG9La03kO53nTanDWNf
qGSMdjSQ8xwWUvv/xNRQwKpdrUDi2W5NbR4oaCcy174xOZhTLdITN2qarkHxbSj0
CnGfOYH2iozx6faT8ngELyu5l28O1VOBlcQX9SDDo7aZzovyVsd08vLRyBv0rvz5
Fz1TBgN1OX7y9YRMUuBxAiRIPgTPi7kM08QZ/wfgWun1G8mrJrjBwJKTttpN/Zj2
g0td3FNZuq80GKreFCWGsXRk2RHtASskwPJ951YILw4vE5vXS5ZRx51AmXFwjPv2
bvsxNMLBFHp5RfgHasQExxTBFJu+SaPWsOgUdAGFlXucBLZ5TqUi/vrmwdGQ2aT5
vlvlGuAg7p1cxqrMihUj/VdReK4M1GnH7bvV/yiJL4K7hKaZZyyIdZDb51vaBpUb
CSZSx6ND4aqv5MaGrRHikIdI2n7F7iJflO9aVnjbF23ten9sInbYwMe9thT6KFiu
YFiMfezudf5EbDWvVHZfKrOWsc47T/u+HhTvzekeGsFIBRlPtN+bvP7sY3WnCwfZ
EYiCGRpq16zjCRxFnGmoPEuitzisFdk2QMJDl4+eUwMpVhenD/WjRSuWsSVNi/T7
ggHLhh5dY6YFPERZghWp/MywR2KjqhBP6I/yh669ZPCHAqPbhYU0nAzRM2hpRrWU
c/Jd5EOBW5xOIBMjYwYDHTShJzniXuX9eW+V48ZrN1XVtEarq+tW2ZK7Pong8dsy
vRPG6UpaUHdioOb3k8WBypt2k+lkw4Wn4+sNIsdtGvIiAoQZDGlf5xmAknZ/jMcM
xfxqzlWxG0hd6wTy/5yWR9B4yNhC7oL2wrKM2RGfoXhnW69PEZ62HGMpS1p18cL6
S4G+nCtJ8MQ+lc8/SDB8xv6OdkqLU+oZB8L1zD9K5/TY2NvJhHhw17qYMMkWE7u3
Iu0CP1WmLt6n+MBQZdIMdvJovpiqyGiIZvtsub2Bov1/gA2wQcN0+t6IvnyEZPql
KZfIQCF0Q4wGiXHtSkd/1svKHkZpoZsBfiuA8fDHhiJDsuE10bA/JIdNc/e4QNfn
Z9k5dSOe0pA5AYTUNrbROpQLfE+sx8dGMcqZ6TbEYO1SBUSHUV4Aq+WMdFl0x9+u
3shq7Gt9cj3mT4upJJuv81OYifHeSvWnfHi2fIiBrrq9Te4cINrM2BvEWza/RKU8
iBERlk+vJgv7GGA41FQhWUjkJJx2oQPm3Jf5fCYN61yQQJ/EeYmk2VK9bYmcZaoI
DdsGiMaoLxMqXShZHqhSqPaxfu4DYNq0rQtKaZrL/5RfGtcycX3twEuOwlZ5yujK
VK4zOaJ59l1nIkFWQpI/lLzcMgpJpI6SQ7rL26aW/s39Pr/k3jGrkIew+R69GlTO
dl1mKg2c65kTKfv0RxSgM16FiKdo69mwLEAlPe6yoOr0eTrtEFNhwaYPjdLERkvE
tFSiuqtq75EaPLfiYKqxKQz8jF2kDzYCPDCcGqjwQxqK1ll58OjBiJwimTNqFSy0
bHutb1XERt14LBVhCV+eeO5c0N78CGsLDkVizhNhLal6sQAhxLWvSh1qZ+T6myR2
A9LSk3e/R7FrWPycE8qbk5RrCvWBlzKeBqEQwH8YmMDe0+oXaAjeMKLMpbtzhftZ
01f8qv8R5gZbGqrdd1JJe4QVEzRRkzQrfvv9YBu7gEHkH+8f2KVW583HjzLwlnCu
H7/F22ctSS+mZdoYBjlOo6on9vqpNry1tH5+zNJJ50ozn1t7X5UgpbNkiu9yd2u+
rnS62HXpGvchfLpKYK8dS1O4K0YWrmznUDQNRL9Jy3hHrbvajL8xeVJyXDNPX5Jj
tYwYqaOD0C5u+2ONDmV1ACiKanQx02UabSngXPO7HjoJxS5U8d9n1M1vJxNjLMX6
AfeTRjd3kLhOnCHDQqnFt8TR5wIsC8y+79cHEoLXqkxtMqw0a0sX8rwBLVdgeSYm
eGXow4kkoy9pUTawM++VbspksU6WPTSF4dwaXG235iBMT9FfwkJXSfya7DN59dQw
kciL230btP9FoMoDsVlkaXG0DWQ610wQemkhl2B/SwhmTfPa6t9D+r8ummg1B0xa
uJA99oZI6B6z0p3zG/4HdBoUUP40Df5OJDAd0PMda2EL795G/wFrACdLCNpfF8wb
wW9lzbEL4GKg0hcY5E8h5ipiPZfb2pzQ+utH/iB+uDHyxy8hv7L6nNVYTD5bjZyx
4oT40YV0Dht/3inn9VX632UDtWe0aOaHzzgJ2L+5tGsKrqNAD+kj15d+t8GFjWHC
aHCfK6Uy7t0EwZ1YgaN4V6K5YgXr6Ysn6vf7rem6UCLbYtph/TxE3U0u2LZsInCI
hnLfdOxoNLyvH26MjG3zglqAK6vQwgwfhToeVsjhS+44mUtVoIE4Mmm56BlSLfMb
CDe7ND4z8ptg9mCfgiIjKWZYIZ0qy5n4ziiXrLuPTfXVfWnVgxeMRvlLzGqnm5tU
OR1wlDNnNNCF3m5piV1alKvZ/MPGZ8QJnyjUNOZ0K8AwqgO994PErxz3MLq5zoMw
x/uvBf0lo8WwL2mAdeYMViJ5p0jwRARUhP/iSczK4WzFJDbYDtJMZjEcpTnW0tGb
uCzw57NCYgXsln+HaGuYJN5VrP9b0gP7NMCbmJ7UAaDoltok6OBOYAZTt9XhEbk0
hknuJxKryc9hatI/rfthW9GWjaapUmQH1+Jzv6hGyJtgKuw/5fpQDjuZuXqMtVZ3
1d8q4fDY5p3du5LO0TTftU/Z6GAE1eQ4M6EKzbk+ChRZ624oYrQswlrQMkCL7k+4
wGY2et+bSDjDEAKfmsX8iDjHCvu+GvQw8tJtUe+qWyV1Q7s9QsNmV2O5NVF0cwBT
I8ChBhg+AWZutN/dAxFx9DIFPheXy8KEeZ67Q93dDQOoxKntlLsO5MWTylG/wqgD
IajXmRCee9nuf6XRICrH/oI8OlRPXoRKoZGFWwDmNd+gZNLZa3fFt+FeBIxmsMk6
jXWyQm5hldaqQ7gPVazTyKAhokdoLoCnNa8ovyQRXNkNn9sG5A9sG0xa0LFQ61w/
xjoqARkinlr7WzWgqXMbrAFK8CU9G3tYdjQH9C4yo4Afg0+o6tbHen72zt0D/vS5
3+lkd9iqdtqyBbqpZdd/k8bY29Y5iHV1myuiYw3NRHw+0eFW7AH83VVtRbivDIrD
zNoTMQHuBicRiCEvBdmZNdbB7m37ZBl3UtwOaLNWJ6swRr4FyzzS4lGNUL94SJXD
ioF2EwxfRknHgHHJjlBxK3qHPy+xzUwrF9hBZktcZ2VE85zi8r7u+7PgZzp0XjQV
GWNvjQnQn4BRKMdz7jkD46pMi3t5stLjjaazMVcTYafYgvmwoRV9IJCjxbbd6P8+
BSgxR5zQE/VcKCDggLGo0/QoIP0wH6yx019jj8EY0I6P1g5qnwsAaW3LMAZXRxzw
tTNFYfdirQvJ/XbmY0l/bHbA6q/Mtdnxk9TL9J5ppkYhIz6voe1Mmhh2nE3RlyvO
cndfELTl4L0jpJ0ccW6Nm4zJKvaeI7v4m9AMSP4YKBXhx60MPGc8NVJ78eorRxte
OEtEtvMjt/wEZ6u+JscZxtiwzXAnN8b+aazPgwpYr1AmuqAO1w9QHw/Spxyln4lq
haeFaOF3xlIU2AdfIkonySfP8wLfyyqMGz6oKXQOsL6JQOID5jJeAtMiwBZ94GEY
7Uq91npTXjZIxWFMbNJY2ETRaoY+WfOXjg9DubiU1/rJhsswtJsz0GQtNH8eGihh
SiDaqFfE3Z5hs+rwhwLSPw+SJoX/UIuGK8HXTALqWPB2pn6860xuUsMLGitigoPA
jWSzwLYDuahcKrq0c2omIAM+zhBFy0yy6n6VFLd8Q/UUySN63vZ4hYYfmlgdz8/Q
haeFsO7X9EG4iYBNGV2wC+TU97kHVDUqovpazwsz9qqS48wXpGPyma0XBkWz+Cg9
p/zT+MdCv4FZfKxLRuk9wbKLMDJK4ujm2mCCfv9uHcIrpwLcKOfQkXXadeH24+N/
dKlonmfmzgLa7L//mxltSbJeOhxVWJMSRLGUkX4NJ3oPWQAiIb/WZdgOqNARqjF5
ng83zCu3pNp2ZtjUrLhTp5GXE0CnxR4ntElauqDam6dVXS7Nq5Q0lNtDtSDbbpMC
deB/fB4st3wz4Ua+kd+5yZcW2UO8KND5EN3LEAeP6GqAPxcbRnzkOvbs4XO2gUGM
p3tWIqoiIoPEdEm88AqxaT02yWllUicc/BXaKAKY9wKiZsRl4Z3Rn/8eX5ydKzyu
GBU2c8DxLIfBOdFh0P3akcaBqKO+6ueYOwo1QYNl/FbUI7qK072EsWuDYsCGkV51
tdoQrRMCzgSA0WSdzXkh00SQh4iIW6dGREAkBHMqDQMkjHqabVRlsPq0n++HUxZj
4xPUfrAKt//N7X3qv8vaBT0GwDcOa/8EMFjpx6Axz2ncUAyw5eF1jA7MrBZY5xQk
QKv5gkkRXsMge05Lz2K+9VYaiFWgY6LtqpXT2VAKroy4mJtu3K73QwxpIp2Nzv1M
x1C6g0GN5IEVRdhpHBV2WX0ICviuWYTi2zgtv6iCG5RKtns3SONbhCVmP63g5lsJ
Bpf//cdF0P93qyCqwmuqC+VjWjBltzQytRa/f6nKSlew3u1n6Lx6qoDRXIKzKNuv
Ga4ayCDO0Eb+GnYCflEBmyl/NH9q2BTOhw7V5MeMfCgZ3l1DbZNWboOserLXQ256
4bocAFKvsGMuhU6k3+GS01mntddYiD31mANTICeYr4JYvZdCc+BxiL27gzr+kyVZ
f5pXS5Ip3ku098dwHONr0fPo2emCynBfrv7ymaArhq7FsftI6NyWwNmrCMg7RDOT
ah9dMgxD9oI/z2vCw1ENUgXyHfWvZ2cXhCiJaVjaxePTyGwZ4Ecbsfw3qSPm/Kyp
GRNax5Ga6V0bUMF+Nom0MdN2jp3hS/3HJRXDjxeDbnsB2aOZjv1vVMFaeiXmZT+p
H6LNY3h6ObaZFkIfhdU8w+JVmv9yBE/qwq6+HPeikHAdsa+MHebVfI3HZ+4uKggx
qNtEX+6um7SUuftUDiBbYm/+cV966Kwa7HoHaJZQH14upAjznGxi2BjTtT+GnbpR
MnKNjkR+pg/MkGGgJfvFmnM6SBEcBSoXWd7cUYc+GyNH7ghyL29Ckj3itlYxhGcV
twzW3ZppI3dRe/Ld2tgOi6CqurVUtvavMtoVXRJns0GWRnNxB20Q7Nv3/SaeFweG
aa7FgpFlOeH038y0WRt4raC0FRBHXV1J1Q0BSr/Egjcm0PNncaDpQW304POTH6at
eXsPzgWHOz2F4IWRyME7g7JAdHtvgQOeBe8JZt64EJJ9acnLcHFEvJXEVIoYI6xp
THLT3TPhtbliFSbFmwkVLEBgIxsl4pcDLROFlI43o9mBX+Pu/FUCZmvHGAPsLU2s
66EkdnskzrHM4Iybn1SO2knSQ5ReOqwncOgJz/Bt5sRUZYW5U6iGdVoWNupS+GMm
F+KIcS3WLS2BN3YXOVxnV+tpU9EbWJuZEDw4jq+0nJm5InQKqtRi9s73hYfDcL5z
EBnOFsWzxEcyOoozTvRHUlEBn15qWH9BSYla+Yg6pk0U81XJiizyVEM2MqelCrsh
+ULuphsb3xJq73rziRgWQfeNOy0M88za3af3QzrMSTNoHQZXJxV4Jd2IszV8/Nmt
KvUAldfDYIihbXA2NASQ2QFhVAi8HydVNbbsbfprS7HDsZ4QtsLJ/sVDF0RQ3sH5
6DXqYrfcL2XVIJ1JuvQAGw//1VVC8jihrwZi+L/HG+yRsYJsedYVxKauoHBUhDnK
nJvPTGyY+/nYtUELLK6YV8M8yWZnrlv9SsrIY0Bm8Tsq7FpsCLwu/v1CJakzvq37
DT8Rf4ompUGPBzbEb8eN8y+tcOk3Sd1wiw5tZBV9GJBG3KsYRy0MQvyYr2EZjEOU
0PonsMSz9zLsw25a6Pja7k1m4zLF+a5rAAXTWkw8Crl9WSI7dVI1KF9zf6CizxfN
O9w791awoOe0k+C5NjKG90z2+OWkqe14yCuTc+IMlNBVduNUE2qeFg6nXK2cV7V6
LNTf6Gh/jompw49bmt/Htjh+qMJcswsM4RAxG0SfyNfbtdJPRsnkzJP0TOS5zNih
Rjtce+JaGaVKdX48q/UO8mw7LYOH8cqyBzNdBfjRM8glPMUjIBriTeUbw1FecRaH
0nYx1VPetdBkDBDD66NbynZdSYCeYgYHq35SJOyWrIdHwEsvGIpgyAMylDlr6dDz
jcykd8b68SQ4rwjikY9CAD0HSWVFyBJKlKR1BSUiLralqW1XIdzQPQI1cC3G3WD7
6g6lPP49UUfoeiCr27tvzjtJ260E1XNONLP1YdlLTv025VTqnxXCaOO+xfxmCcbG
EbIcWB+NdpXyL3XsrkCc6PnPGNnhZh7Eeev7bJlHgsdVuYtPrNlgQuhcpAMMZ2+S
RIJGjvwaLQz9x6o7P7/nAvQ5ar+YN5elmdTK7fXPTFC5qa9TiD4qHwSkDp8JNf+4
gT7cHtRLxA6JlYcYGut39UZYsuXft3nmnh5LGuFK8Ck1mKLHcohTMuzaz8wv6Mvo
cRHo6tKaEBz8Em1YjtN4MmyoWrscPXsZxezMGb3oM1A+EGKY0/A1n4nWScL1ZI5/
X6W5EXgMKHeGL0uYjopbsG1H7zFI8oQx6au6tiK4Q5xFlzAZl3lfSMDnmMJHZHKI
2UVYBNIzh8YBgWp7zgRefG8YAgQ8x2sAQmCNbtxFyD3/UES+hQTDwgkwBzp5dlzR
XJ2VLLIjANOQvIPxBgvA4u4J3A9lbwMZhHamkoI8i3VSttYRZBPnzxTv2ngbY5WX
IZOpD36Pu9v4guAz1IBu+EbR1yHQU9wjs2yvAdRsNTE/ogl+6Wg7WsLuowwoVbV/
IsUhassNEeOUlXQ9eqCYvedzgCDAfhG3pv7/0DJi/qsqtLijia201PX3KEpDMT20
uTNhx8C8YI4CccvN1+PFcgeJw6S5oj1gdWdcxGGgqadwaWqrN2wemQClvoqRgcfM
Faj74GqlKogyvaklw4omGctwUlynsJ9OhcDCvQHcESI=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nahO9nwSuYfHz3Vgx7k8WZyqG3cJZbM9qVpdPE7KYFTZfJ6A9vdb55i4e8a1LECT
qLWDbZNrylgCIClNBTAdRxFVvk4CsAzi193PobXRMaWSMeN5AeSYJs4xqMRRJvT/
tn8nlcrFBSLekG6boUM5eq8HSgEvnlbTAMkCMm+0xmvSZKsCaJOQhZbDOnJ1WuNv
4PqmDwT+vyyUnPxyGzJB5az5O7BYkFENy7Sd3/pLB451hwgCxfEkxb07nxtqhRo3
WtrpLEobGy51DKFPwPTAflLqd2m/R+EW/l0JvDbDE8BWbuyTaoVrLB95kcUmkea0
cYB63NjvclpfBsNiUnQ5Xg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9232 )
`pragma protect data_block
UtEAhqa7EO9u3ex+9JZM3h5GXytZh43j5NSSvxnMrBXYN8mU3DUFpNs9vOyrDj9k
wh50WQ+KZ5CH2T0Gsf0MLPMD3sUyJ0V2fRSJ+f/t4QC8ZSPsg5cjINCqKBwgczQ4
Gqja1ZUnRNv43jx8jWdB4liUtvXlXba5SAW89ZXv774xOFviGsgZy65nMwEzn17G
r3stpd/UABcR4mF/se163fwaDInrZYVMuxrLSlpsPv0v/r3o6Kf7ybb0zjBlFjF0
XLRxQFJXmuj/KMRgCNU+3y6lsoHtrkGjl3l+6xlP+gFLA6e6FFXQGAxIP8njudY5
awZiAcUk6AaWbMwH7I5116ZmIsEGKFTKf+64OETAEaVh6djecPijWuQEj6sjV7wc
xRy7zfiYG7Nb4Jx1rpMgF6Dw/OLIW3uEXkkhw4Ve8+YUym+NluSwkWLPy1gqAvnc
olI+Sho2HQtHRfcBuCOpa7QQwtEmFNWJFuZd9xv5xzGeHLnPyYt8rCgEJBLc9iR4
HYcaE99bxpJIacGSTJYlhESGFxfhAiu3TMpHv+UKD12AqlGy7z8JZk3dgnmX8hXG
ELCG8iaBGg/Gype6xirYUPVh4Ba2d6dLiN1H3lS5nVi1RqGIjrENYQNKZQRVoTPe
BIlcqLavQ+l0HhQM5n5T0CfaqNSUtbBXMSEh3aS9GU0M+m4FIoMQN7akMt7r0FfQ
vxPIN7n4oH4KlV1mPRdQJnH8UB5HOae12uYjlcPopMhBsBg7ovxGG85Ihtb1hXd2
+a12Kj7WY2va78oGOt+0d17bjgJShQqKlJvIIKSQLr5TQWShTN0QyNJ88umCZpm2
tIVGarvkEN8gnL2o3eCCAKwAKZLSs1y9AOvXr5qITMAwHCLAz2OOs2Mu61AzKyz7
k9wHGOYK/eGhrk3PbIcTAYolZXtSUOcDLQaXgAiPq2KeOT8OGlATZ/7X5g2qPsyR
xwAx8ljZeqdLepIx7vu6/chLQDkLxQZk0jNipEyJK8au3RaAYsnW6TbFZaOPTrsu
a+kEMluqr5ZnZMcpxVvxqDFX+3xj8gZPEUj9+xRij805Z827IDcFK8BYq5xk/fn1
nXI/O1VJERGOsw0s7vt+dM/pU/r4APMvn/uFPKlIrqCjrZjbpueBatPArsbDX9Uk
z75sdUuJ/2x0w7pE+76rdil6a8GLqSKw20WDMnmnayeA8y5XhgOmaxOtIjMQpnJZ
WcKpi0NhPzhks4/7WZIKAKIAnsEM3aEtqSJ9BN9FX3dt/eXA1KEmL5VxV87p2WRm
zswDGKgfF++Ef7o7cKQRNk1wvoISuuw52TC3V6wxuN746mV8s0eKQmdiJNjOshjS
ZgqKW56SHsX8d5TUOrZ4tQ824PLYYS/0qQTO1Uytc+mbN7KphpwOBMn3G59Q/Ml2
07tlG4cI2aMTdWmmjqU8a/PF3vxMhmFNuy0lN1eGCMddv7DSlaTGuGcpvjDPMEb+
pjhCX3glvNmeNQ67OQ+c2xALS03olhNAUhJXWeEVI2+jTSNMu2EwLbVDMM6GGxur
MrLeQtw8JTrvzlkMKkyJQzE3Wj2XFDj+TM3Wbbdi0jlPR6OXRQNCfqtgZAh+NK6M
kQGl+6Ok/8eV9Jxr4P3N8CG6zEOsPxQ+s39b7jDE7qvIFQhuvAgHj4ZxnFm7nV8H
krqAlNb8J+UmaAR0aKI1OwI9xPAiLz3SRIMHdjpNItBD27DNzCUflG8gaym/Fjqi
2m8NyxLWjUdML4QsY9YnEXaHQ20bPMjpwCGZVyOW5rZCsJJ4I5gX7jIzjoEGJnOG
iTQu9nUqq/45KJ3LCgmT0o4xHWKKqW7D55dU99Tf0/ftfRzGLjs/cQwlZlr2LrWW
i+JQfGS7Ur0GUgtJE/+JG3eiYBrb8E//UEzkr4nM8WGlpfg7gLwNx9htTB3fwmNA
lROx0YJyYFI/NQ9eZxVd7hHF+EUny9lq1elRe+h+RWBDls5yvqdSwAVs0A4sNKSl
S1/NCYiLe8XZZR+hF3FChI92bJr9iO7l43kGJWe3DCgzE+JyCNtSRG7Q/Uw8enZy
pxesggNe8nFqKk4Fp04d1b75Fw3X8aGXQiNYfP76ptLs4nzSOfLKPzIzn6ejY8tX
uB52zUZVSF1vrcUKrC+a2/0gaGa8210UbEufrv+PmID1Ov5vVYHRxlg0YHlvDxZg
1G3m9XPMvc0OK9ona3Y8iSx1kqIT7RQp4d/3zPs1kCSlV9TCPgINk9k8LMQ9M/9k
gzbUge0MOxdXdljX+N2Oir3o3P0UWhEhzE6hoIM8XDBgxReqHnrIwyj2WWibSaSe
4osCyZkmVTLBrZXR5I6RB/Yd27cGc+RiO9XeU/Mv8xzgLyDccxRH390llXGCI5eU
asBuT1eTaJGFGirwV6kRY/4bjuFiVFJ36MJE/zeI4NUe2khfpEODsailBWZpnddZ
23SGPhzy83oC5OJASCb20i9r3zYeMwqwHt+EpyVCfzPRXlSS9TayreLmqqAw2Zx/
cUIi7seIQceLy48PWiA3PXBeFo37fvWDBtasp9GeOiwlLVDu9yjXMjNo4xrhNPFZ
NXvWEzyyJJt4gOSxYkxnB0r8D/Nt8JLgOxyuWv4iqjSC3c0ITM4KlXfZgiO7sjxo
R2XId/3bLFtuY2CmXJvTDQISlmAqri7CxeiH7CXTzL1tbf23U9Nxmhx6Bu+muq9c
46AkBEXSwRxaHkfF6VVNDaOqgKiaen3lG3dQkHBMbs6zEEc4szYz4cCRKYm8Tey2
Ws+u/OM4QqRz1+5eTf9z8u8VhLim0YNjnFeZ+uHaury/woS3dKyc2xTB+CuQeNgZ
CEQEFuuRWyIsUcuE5IEwibO9zRb67x4/xWtUN/IAZmGAwAauNcuGpRDuLZY98bQM
YB9Fzgxbdbn+IvZarjSP3WCOcTRkXOD07mjbTjQky2Gz+Ze7m1UrOu26EbqummeT
CYrhOc9uBQlp6GHOGycqW+Hb8N/cuP4Ik5NfF5nSFN5eP6Spakd59JfnreSEuegT
3wilmY+OlEPf2Yw4NZaacSt1n2fxvLhSktBOnKOQWSEOqDpL+hbORN87xvPY/ByN
JuWqr1FjEyXGQTUPOhcJapr7pvR4n2WC1s+nYn2gD+bL7xTDmhd8fxAYh2780Qmb
e4IxzYYe4YCH45MM0KriZkAQ7jlC47CStNWdPPXZ22NPGOMn40YvUCvShm30xTd3
w1S54mj9EeA/tRgWhFh+Gq4p6AtNPI/7ZBtm+0t0K1cqfosb4MjpR2bEGkGAQM7b
nTrSfe7fF/uXYbHsHFrQ8Lkrr5NaoKRauoEehFXMzXCnC4MnZsUSpin5hHEQuqH0
CK+J1eyLNFXW295cCx0djSA3vbMrZD9NWBEPxCa7PdjlGZAtOfJ01lTy/M493W+F
1UbDGsqSIg+zQgSeZKBDrZ94OrA+6Ub4AgVc3zHnj7aWxAuHZ4wA+9yOhi8CGNCn
86XnZxa07T0Q95xG5Wgp6O6y7KZf9kraYQrIo09nGf2HFH1s7mgLhxo8npPxVpcN
dMImnsL6VAlM6umKbVpqytwzZDXyWX03zB5ZK6lpFZBytqCOyDz2uQHekfxJiuWo
BIT6BN751Gz53tuYMwCdAFGrfEvIHfq4xV+MV0PFO3FqMuEC5lvR7iQ//mJo6KTv
4WGeq1lgVzWb2sTMySQxVTpodVMk+1pGtarVFVAROzINTsmWRtpbhQyGsIRYb6DM
vxEownbOsNBSv682lggZZsRzHNWUJ3FdplpGg3JeozKtOD1e7yi6pJ7weVk8sLd5
O0COFIotn3wDE34uXfNkLs4bmXqtaWhtOTuVXsTwQYdXZrnOjPYHvYY/ca80hBFV
/afZIdf6+SnvhYoZZG53fT/Hn4P2RDmSQZE2nhVfxQqmHEfuNM15Z92bU/WPY64d
lj4r6lBGKdewX85ywjEs+3kbPDEySKqqnIMFjaR0DMR3ufSQwHzC/htjF7wV/RIU
6EFSfy8STmyhBJgaXHdOeSSB0GThFPt2dh9MLkzXrFEb86BkTN2dhix0fpM7UQlf
iJVKiBnDE8gN/tvR+mxpZtLsObUlOESNou5Nx+cLDFJlTiY+1d6nshmjRtHKp7jN
1ZG5oM3688D4mRrBKe4P+ulhLRQpHh3GXsFBL4CWJOXhVRkDNHjkR2A1jICeClPU
KM1mcjRN1JFOXY8mC1JhAx0y/bCgwQfhXumcMNH1+SCOL3Pwjp2hUQX2Mstk/Eb6
owlawFLTAgGE6sa9bdWWJdePSHmvJHGXzV4Jn/QMpsjGFUGEOIbSTCUhNPooCyZk
h4+yB+c7S942KFgONBcaHUSFBFwcELo6h9cq2KexujyFBEDE5RfzsoTYL6uDhWsz
Sj0YyGt3VVwnKACNTfPCbX1tyhIBl/GDdaX87gZlsDwfCNj2N8tYTo81OX7BykQd
jIIjc0C0NjLMf+qlnJFUAFJVDj74ofjJ8VMyLvxPkLrmftkclapRvm7X7zJimMdW
/M+sWe8EGty5Y0HGJmK3+18Y9nwMKkGKxPJidH7HybhRThn9o13QdeUlHlo7xvb7
e+ARLHLEBdj31D26eI2WmcIeVUQv8o2cOzvkd6xgUQRsRVuz/1+DpFNI/+duWlBa
/IhBEIASQQBh8AKRU1SblJeDaa0J7VAFdCQ5KQvqsdaKSoTJ0IY8n8atd+GLNkrW
DJLz7EOYf6/qaZdDzQqsVHrqc0EGYDmViPY9xxQwH6ZkdIFrN9eZoZx83pX426Li
Ox42lzIEZo+VToMd+uCAuu0KV9E48Apt9xtak97IdqMkzkrS17+vHoYMnFQQsT3X
9AamsmGSSdDYmcYq8FpQzEmVVz/pnuxOYqWEP0BNeLlEteVCb4mYlnJdJA9OoZGV
jJeOjeSBhAf7pxr+hnbkFlKvWyqEMqqwwpp4N/Ts5xBF90nxFGQ2cNN1Y57z9ZPz
XSE2s3shWBUvtqal37f4Lo4ocV19kof0sOy+oyb7g2bCKD90gIR0vjEbO9lsvjpJ
G6f2Tw/t3XUuNoPWMKrCZvpN8qqcpk5HvroaLTJo1Y/hqgjrbN3WGn869dWfuM+t
i3fbMWyT9ubkPmIAqP1XlnFFmkkMXLs4TvsVwlEFSHaXjLW3UD39DTlauCaL1+j0
Y7BfMP31/MUEsQa2BcGqkNNOhUJ3+pjENY8SmjAVIEtaIoPliZwtxJAz34huCj7d
hBNbI4uODZO9fLGlJN48nZGQFm2JVBTblPB6GJOMC0kgPgPKDYMq63XZaJ8coJWk
jvq0MUx0/EpqXNWti1yZt08h6BPgm0B3Qf9pInZ/Cl20k6cxYKkuUeoIXYAMRwNx
dsap497AIjxoTYiWChjHDl2IxpuBSWkh86QyG6vSMVlcNNvTgvmOdYzN0AlxGfOl
O6tQR+bUrqifE4zOP5ZjBbrtCFuY5HRhQBbSTr+TkufrQa64Jc6bd6hEXL479Usr
r3rNElh2EMTrxyBexrOxCwOGlHGEIOZuuDa+po5Vu0JSr2EByOvWulnDaOXFbBWC
GyvLSjK3GQuhgxe5Gv0aR1BB1uB3B9zzIKlmg5lvo1gdwjGinyNDKOHkgjAaDONd
F1XwEB/WSxpr5maFrYhaBZDaBZGkSBUZkBtsGNsS5EdsT5vwhrt3VUlZ/XlUTuhQ
zPxwR9E/VOMHxyt3GYHhmZ55lZmr4ORisaV7EuGF9oxhdX9rR6vFq3BAxbgj2ZdT
VI/YEl7OzQS2DJ4j+o0/9FKFA1uGLFMA2xH8igGHr8unhF9mAOa9CYqQ9aC7jYsv
t3tFEZrEjfehQlDuKdwRkycEq+xpDfNoSV/7Jo5iJF3eZtWvdg0FTD/ZiTKy+pDD
3kDsDlpS7Ypi5D/kSNwpsqFTy9IFRFyzuv2ZJegoEMIu4nb4uTkdWmxUJaxjPnE2
bIUReIPKtV+ZKcZvR6lE2Bd1Dn5y6n+n0ZCjNgUkO5JgXPluLoKpx+T5zJQ/iygO
V6lXi+8GCSABoQXQkRAiQrbPwTh8qXUB0VVb9SxsFr8scNyJNHRcWIjrBTyQwdv7
EukqacuPfLoYMoSdKcxJfoMWxydEUWqWbx9DP6tSu3XlS+tshk7A9mZqQhPI51Ar
NomU5C14YeJoawF4IY3IE5is0e9Kj4FxN90M9WiwPK+O0SK6yE48yE7GtOO3o1IF
Sm0yK3fKXRSaVHyAHMJJ3zti8kuXoze4G123G8hv5eCj9IfdA8xS4DFqL39GmtyQ
ivUPFzkv0P8Pvjamr57z9Afr5c2E6nlcxewMIgCiSthe70cF2E1OqN8yjz6BJdcb
/fM59VqpL34vX2sPa6iOzK0M6MKPzK2lZeGcL50v70nLQtmc76TLrh4IEZj8rJiM
pcN94e5fmDM4w2OC+1f7xgcTdWhGQgXVyOfJAMr4dwWXIXTgV/ofsTbj6WI1g1wQ
ElgZbtzxP56lpJoKxbCFsXV83Pb9fTLxgRZHzicWQGo26AfSa6LfPm8AbUjO1aYY
HASD+H7E6ScHfAjuGv672JTp0V0gzotNITj5iKdpLzRLt8LABNLTRNZ7nIypzu8C
zPilgUhd/tk71T+VHX560AJC/n2aT9W9Quxcbgcq6awFY3pwUVqDWQTORYnoa1hZ
EZMh3dypXiIxwqqaIcP0byloKCevuA24WednQ8j4VYInH6+5rWrB1tUcLuL5cqTy
LblyOI1RYj7eFxL+RA4jQieOcpaQWzXHDbQlkAOiAJhudBX8b1qFHU2NHUTowWAb
LCVQBDRttvAoIMmzcpaFMN6ku39OYyGfi/oLnUJVH8j583KzHzxjoBawOBvgwlDD
PskzLNrNWrnmN8fsZvhj8xyOJKSIgun8UXQfiP/IjZeiopeeubzb+qVZCEIuOqFq
UE1uITXkWOfoqVtL36efjOP0G/xgVuMietqMGdyMm0wstz+wf1VSuIGo94sBiWLR
r8DzfyDp/yGtJxan2SZpp9JV3S52Wca43eW3nEzPClUNn5ROjsuIvBNEr44Mg6b7
JTcC9lUpcuhDtDMaYEYW11umxMeDi73PeOdttfIwzGAo4DAfawLj+OU/oh86urgQ
wAEFhX7T6uca3s6pFFIYpXhoUTHYaOzjS4vu4mtOank9s5tG0XXoiOxYDmRu4vDd
iPjfLRFysmCEez4Oet3anueSlTxHYb5ZPCH8cXLo//PORk3j4MKjHvz2q0nA8Hpu
bt7avpYt30H4l3iXx903Nvjbvld0HO71M3lMqJTpZeN2aIitjF/JLFZFs3RrZZqw
rjFHdPd7NbL8PI+vt2lqYcZBB6eJuNtn8JW7+8JyNoOaD78QxJDboDrDxuR0jg2T
G0cq5cY8xoP9rvCjVRM0NtEKr9vRLo4N9PhwAwQkaCBG8vTvYd3L+fLGJjO/vqM4
OJhs2f5E0KGVZwww6JCMl9eO99MJ7P639DlqI9Aij8vvsJTgGuXrxCPU5DBBGgwb
QftidYtGxrb6WyvuPN1+zuEAMzQjiNi5GsGPlOwN+7kjegGtj1p0yQPenX1xrJch
V5GnAG04r4koBOvai7cWSyRbcUintIxt319qPT7vV3xDiFPrGopOdCx5ul8TsJY6
VzkmowGgy1MUJ/VuTybvCvQ9Gb/YqzwBrw33+Pup0Gj+sb0Gr798PafMxEE6LyoU
KTwCSoiz4pT9Wb8jKZQXwFxMGOjdqWkjkoDPjDWCLGVhg3S5XEtbuBqWIsM0+0n7
1jC58LEjoO1aHa1iu2lZY/YVVoKWPNbHstQnNxwPY6uvkGtQy/tj3/jdDpO3dVZF
h5Lz7RohSZQWFTtqJhfDbovAFI/MLS/6Y2YX9Hz5bEd8t2jpaxGUy1xt0YJh7hAy
U1MxobivhnJBH0ThO0u5tQYUace/V7B0DnG+a++RCNL2ZV2A5/n6Z/vhAqr3Fate
Rj5GbCqQIi5j5u5yyrIrIT3cd7SAFEZV716TYNsV29/ZIL2HqEeoG24BlE4Yjdu5
APDUJv1JmdmaEWxJshqmSj2Vmi3d1zwpo1lElB5MtARTiTDpxjmcU0THPeOKoiRi
pPTaFy6mQJnj3P9IZpeOeGXC+T4DL3kUtEmQTcpfISLVzNwF7aDAfEXIPytEp+VK
cgKSBMyABB6vQcjTiYzryuEUwJAqj9zxbBsM/ZMBFHW0T4B82rZSFtMIjPFgp7s1
a1GJDvNVAOqV96cVqbJYmsBYQjfiuJQUTallsmbVFYi/S6A9ExFwg3/JSJkCCmbU
kmX+lI23NOSYnAvbgRb4OSN2R00dJxR2l9Cg4e1yeCq+wMwN/w22y4HbrDzc9OV3
OkITdRxKvWAB+iIiINKBdso+bC/5YiCN8Cie3Il1Ua+Bgft+m8RYWrBdbLZaDk0S
2LHOMB8TFnAfmHEhNFGu2gryDLnRRo2VGpZSu8mfQElO6KdsKM0gno71uy1FXeUf
ucM8SFO6TAZeIHFruZJ5vB682WzFgCRFy6z4gUqqnRGXnkBvxAPCU7Nr6YPKCoa5
FjPXxMyM80wAr0iopomPT7SGJe/0sV0QJCWASGHsVLwVXK1fU+3Glw1oPGzDDXP+
+POqlWf+Ez4bffN5ZiGiOR0E9tMwTJ5Pg5+g5AQn7C+y2AHaR02hmfmk8PUvQKdS
YuRtTrqEn/clqJiQkWK0NUcvagG2z+034BbSG+MNg3M66nAj46sjRfR0TUB5kwk9
bZLYHlC9Yn+TbNxs2dJqIi07HFkCa3dFTOIISDDnrIm3N0AZH6Jldi/vCdqWSYNc
nk9KhBFP3L0wIA4GYBr2KdXPy4ixO1WEibzu4Gi4xt9kyIPwzvvR80Mvo9otruqk
UbciQ/molPuNphM7ngZxDn5y0xPf2KPqbQgqN6vL3WQWoU/0w+FYwPjNpMHdl+dE
pxXuX1Aanm1KvzGVCWOw/Cei8clGWcVsLZuuLk7JP+TNe00VX90rQPqOxQRjAcxm
vd/0QbUlyPTFq7sDzmPfpanA73mVyiXfJm6bl7prg/8dVTfkGE1BbdIqYZfNR3fd
LwMByi0JBuH48dBE+pTrEa16CK//OtqtRJisc82oig+xb1XVebUCXwuhd8YgUc2j
lpGCw6MTKV9NxZiJHuhAkcg8XPl7mFlXTeCNPCwQPT+ZCAgtx5eRg+V8UCg+JlZP
jmQcH6fM0LWQAVQ09/w18a/LnB4q0F/M9ZKchXtOS8SNhovAq041I78vEh9E60tr
eIcTTyQKKlIQLK3iXj5TDCADAtKaJQufgjiMZFCyvD+Mmk8IdTBPxtA1do3+sCT5
1GBHi4GvzISGHayke5ukQrBWJr+zHcrlSqKYFGvqSwM7zBhigUVuVr4vIHhlInxk
X9XUlDjfORrjeMNFL0WX7Z3IqSpGkTsMfHKZOGCwsLlGhAT9bJ697bdRGjMtA87R
Kxfo7jAW0ge2tcH0nO2fvHAXFqnCAe4IsFGXihOZQ29sDdoh1zmWJlhLSozSzC0w
OD6+pakd0f7mQl7hJiMbSjVslFZQAQCWnseBck5GpNUUP3dML9KFQEeCbKGeV9Ab
rKTaND9lTkRF0atpj7rvOESftIEob/7UzAPM/dm6kPrVglxeYMIupBYQFj4cD4Mb
/3aEo0D3PhutujJ3tC/1FRnP3XVA06OB6qEcvsQjM4E8JPayZvWKvwWkIV3hVJNh
luhai8AMqbClGzEVghQD+6qH7tk2EFBL5U7lX4l/cUKzTkQyVAQjsgvmlnPB4Oti
MjH/vgjhlzl7i3FgGrScQPmMmaMJzH2EZeIBiUeKfdfgdKckglDQnuczTQXM/SKW
vDi8B4mxPv4pVc53wGFDo0BJGmHH/QJ2CLq59erRNS//7UH2CyWobN6hH6dM4J+v
8Re+8ifhJ9Wq2K7mb14pp5MlOZtjoT7zB5OZlLVK7rfouFYBJuv1prt23TbbC0e5
l0bDN4QuauXuKMsl8z1V4xEd7J/o20uE65x5JQV4kOGZDpFpHfwXZ6DdcMVv0hBS
nzxdsDk13+mmBK/JVOfzUQosa4xIYQZNbbUn4V/il+Mkr5aYgEqIRyy5sD6Vdnm8
YRhacKjzMtkDV50h9pSczJk4iLy04mSYVD7Nt0os1Kyl84CSK3WqcV4t0mZVd+XS
tJSqpzCkBXX8PfHlEt+3vp3uwE5WRj8mLijnOCOtUThn/WE3Es4NXTVF3Ez3JILx
TPs+PL2TJf6SyBhP62C5XfhcfgPb7ZtA34hkNbmEB491Nf3Hf4R4o+5nkk5Wlbx1
PJTeRC7VOtI7a2EiWW/udFKiM3sI2xKZku5F/K2dnvnwTA4j3/2chqbcCdfuTtdj
YwJ0JgP634dWI0fyeookVgu0PvNITR7v2V/CVWMgYw0hYpf+aCdzaW1tgs7L1MwE
WVIntT2mpuTsEvUYmCKmw3uxk2T3fLMyCIMpUY6j1nReDJXUL6eIk+MdMzmDLNrU
Yn26jOwucnLDpAI69JD0bLo/WF/tAUl6j5FO+CtjUTgV3E89dRv4ANPgqtOHU3Y3
ojXzDT18K2vKxo41ZfVK62wFyVnzdsAOR2DBwD/B6PpgpUU1ucSPcWBpCy27mYU9
2fOthYyqOvm8DquUHEAtecsLuqBDPpgQZ3DgstCHhgFRb6Lj1q1/ukEgPtwz3OvH
kRiGOxpCKNNlS2a/TaSL36VM2WERxvn+bnJBuCYKgvHDRnvR0MMEZ6trfWsPR1ub
6WDPLQ03BU4SOOqLOXezF8OYYbG4uvxGckeDV2prlFjmoq5z8ERVFSX4386+fyBC
zw8yvdMx9tDQTImv7/uK3RBuk5P/JKzPc3B0RPoJm8RCUp5dZxh3I4VMdqO9n+nd
oAF3fXmEUL3/I7uDm6Fk7GFOjrI3UUnxvzIhaGryoaw04Yk2x3xbQR5F9hEorFFa
MRjmwIP3DJ6NbnOVkgv/JmzoZEyoSURv2037Ygo/SNywuzfUVZzLjASn1sGgegAp
ZUw3g3wVuvYKQHOCEC2rAnfyIrYVxZBruWHBl68lLqr5+bnNAhfpHuUSxgqAcMLE
1F+PKZ6qIHAp/Zkac4BWANUx4p4o/dnt40RbZjyuX04+Cx4XOs9DeOL7hEeWhZil
EsryQ3ns6uSPRsouHBsiniyhKKMQSYkVO4EXFJCWMTrMgllXkMaa/gy97qFoaa4d
imFfxNJeElzlIreDoqp2YhanUnl1nIlsAVtTltUpuNimDKzjEutmv7TAzAIv+Vtm
ByeP5rgveUErmmMnm9cTyWPTaK0m7l9JxNZlLmnVBp+WnT7/iF79cCJveocHUeT4
F/nyXIoajNG6eYoCzbqlvLc5ZiQfvLWzNKWLEi60Yk5JcEOqEDUfTuju9tvUeJfE
pY7YTeDXxJryYzBcYboIjFwIsHQbgESbQZ8QY3JAFOF0sidZpx7nVOxKD/Cx6mB9
UdELIOG9tloi35pWgtB/JSDd07GpkTZAj5hVwnaZKtfzOr9ZEQq3agohSfbhZNnU
e3cNBsAy2mnp205e0X5cJWwjPKTMccTxJm/YyndsyOQQMkDd5DI+1nq99kKA7zk9
rpl4c+ckezWAwwsIRaP+e0O9pATO9+a0HbGLeOfPh7X8iK3nFkAkzaSxqzIGJ6Wr
Sr1oZ7LAPzjd2F5zzl+DDg2ByJgK1ORljXmcDuLWHchjLMQH55O5bb5QxVCxvuvW
3Etou6m3CWR2Rv7HZ7vrIFxHj2XBdaGsNU8k4ED2FZYyrJfJ/X1uCo93oJ/AcPlP
a/q+YR5K5nCzd7IP7QdaImdA4zxIo8tAW/9ltUxQDW4W4dJ7mARqaIYCDqAmw5u7
LlCCcogNj9y/Gb3kglX4JvzOpFX0UoT99lRM+Jt0CvdNKn/6tLHan50vBBuZwJxl
/tDdbGTfNVFlNLsJ/V+wN/gvRnsVomS5RCzjSBqtOESGufzdzfdbFwhuWk6X6u/r
cnhlY5pUWRsLTH6nWncAmZsIQN01o1aQVOPcDOqwuxRx5vwImzE3ZQ6vUJajRayg
qsohYVERfCycGLZ0BGcW1p5mR/g2YDTm+AXAa4I/ExC0WyTWKtt9I7YGNhMIf4bW
CgdHns2gmh5kJb8Z0hIY+4np5VYGqXrR+2Rxlk6uUUTSS1TC4KOfmsj2YBaIpnbX
SHYbyLkueCZ4sa7oee5tlHuDXYgszIN7JZrams6AYvAfKc1/tAeuzZojlajyIXlc
jNIHJcRCs4K3YER1BE7xxQY7cflnMQBB7ro9+a6H8H7Uv3nGW8QmvgQZeE2fSuZP
7iO+bFanZCNRvXCd9DRoTywgOIhhV6V0sgwhqrI2g6/xq3KU87oUN402PNOsvA6G
ki+kihuo7ojedLvqlQHUrQaAQlQ9B+RDlnklv3eV/fWXmc349oJMFdWwQzcyEwJ6
zy8R1JlfqlBoHfevJ+zrGg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
T0EcLJHqcgT/Pap78E0VyfWXCQUpBp2evhotuFGPARZD8xH35HbYaYPEN+SB0hRt
tIGKRKMtxHjSIzJ7Q3kfQhk6tNkykqfOEVU3yLgbhX9i2HCJxfi+se1u/pnVrdj9
gTGNYb2FzgxOSeRj8odmw6NaUPkOghKbw0amxHriunWio+QWF8MKpeLhTZMYGOEk
yFRqlWREkuD3E1Z2HaokotXOowWFoj12Mc5TaZbOUvVa4p/73hMZCMtp2uhglwvX
ss3Y8QpBZWborcykfvHbviNsV4W3hrIvg05QqNHJ/Tr7Sbft/a8A6IbvrAs/AFkg
Ix/A0GjONQY4lqhzlPaw9Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15408 )
`pragma protect data_block
qrCSBZYLCRdrXl+IXboeU6QpgeuHf6ekzm3BK1DaQKsQj06wJp7h/Up5D2c3kgsv
yN+eFmx/HMFIN34XJHDRHwscOUF44uGvfJtHVcr2ENJWtjkSOgR50mZJsqjX3P+w
p51S7YokvNw+0hIGQHEzgTLrC6hzEwTyB9YPXmUF73REvxkgtexoaUkFBMSoBzQn
3U4tqw250GFrrTIij/kYRbe811/U9fdEM9Icu18AkD5Ir/3TkCoUCuHWjFNS2BhZ
bbxwSvDN1OgPVOuksHGIRy6ANfEd/si//fI3iSJxho9n4WjtXOQLsx1w+sik+D1Y
42NMeGtwGw6wxiPFztCH7EEv+7bS1/AQOZDH5Dfo1BObvrGYdTe1BEBcn8dBXt3h
/04TGotmU2hmrrYW1KY16owa0D3bWX2bnRvSLoalqF7zKelTiqAIItZSgYfn46lq
S3fDdJQL9aTlwt4A4YsHoaOlMNa5cfACMfvU3EPpCoDACFd8YlkvTnEH3+7MOUOH
++R1eUnC8DvjnJm8wX/FFT+qYiDvd6ZIZcBQijYW1Dk5PDyxg5/hZPcvAIbN2jxS
jMkQRYnAJV8gdvdWh7sPcn+duivVsFX10B2Ef98+QyZS4RIZDqixvJth7yqgHr9M
jUFyp0z8l7/YgJB6ChYNRAuQlbI4BuIElxhJpxd10qc5HkPBCp5cNgnOOMS+cmZ7
8gJojzYiS49uTo5bldZ6QzHNelMjcw48uR/Mbt6shQZTFXW/suoSmipQs6uKpqtm
qlYhl0XhXx1CTAcPSpbvqiZPmG6PbgCu3B1xGUiK/jQtKzhcTmO+/v2NEW06q0JA
mORPMAgfAxrUqJ9VtLSPis+F/wLG4bDgcZvV2OmW1TZwJcPR4H4C2zBLYJqB0LS1
ACH6EAvA6LPkpcA+DRQL/fL4dBWxRK4WmBPN0NfQYR0/KNy8znXFhHUekGcWQJyU
VAmt95BVI3I7q1ZfilGHEtkk1TfxO6HFifmFPCzSpYeEl6dVc3A5s02nwSHd6ZG9
L4rtYAgtBB5C8sXuijo8vcJnHVAY0Vpb5xjgy8EAkgNBt5BeucqoM+ltxisWnf6d
1zVo8/vyC1JiLo/kjWb6SeWOH8PLSeG+x2r8UCwoRjCTQSzbQ4NvIL3Zmf3Of313
/SGpHrq584kiVwY9+MNplymn3Ivo7MS4IdmNS+Irbfhc4ZJdIOp2J0N+8Sb6yl55
bkWHEAJU/X0my8+X1s3dtvApG8XwFgjWq21UQclRe5P/WjRcBpxa2WiidFUuenx9
Cn7BBFKdvwBbdIBpQyLbDbXp2GdiL4J/PbcEe61LCNXXORe3nGefcwJUsARLxRAP
jfEN7NfWIYEneQUIYE3tAjlmAmO+vHM7Qebhe9gXMuoAjDI+u+iyUAGyqkr0CcM6
mZJ3/3lZlf0AUurVRLj9Ci5PiKndxOIvZ+oDHtGDAuGGNv+X/NWxzqd/+lUd2xqw
zrHSnlCUhw2l26GzUREDO2R9sLkb8dK+xoY1InpZpoT8LRZlQjM/Ahjz/l1Fl9KI
0xbDwJP0JXKii5KrlT8H5FK/mz5zqXKbdR64Fc9DErPr6Yw0C59/lWHpkc5y4Mut
1LT9l3RKgBk8tPZL2DGf2mx0eHpv6nYqbTr8ig/3YZKpvn24vIO9Pcfusmwm+64V
fHp7/GSxTlvXy8/z5U/IaH5r/+5zom2HazrSbhlkaAl4pGfZ1GB6ELx/YyaxhOOd
hOCdMbtsLmgsn7iMLaHTlI7u6pVP9EDbOwIbr2RZFF9hXPVo+PCfhqWo8PNflt9J
cpDs7rmwklbQvhRJ7ZLlXMpASqk0B7kuBnCBxISASUl9o1VvqgsN064L14WG6THU
K13G3Y1PKIcXRIbiUlshgZSC4az9f90Wz/Dskp1JI6b0xe/Hpg0Fe/g2vtSTd1KE
wUXN+qq4UUhDB1J/duM/JJwrXfkC7NZk+Dx2Av7OyUloujuPYxWGDdroqBJYEcGd
L7+74IP8ZMh6ycgWs+HsVgGVCrG7No66duinopv+vPxeXZW0D5WgeyeUojOjNJOD
LUDqxsd+VMIKPt83j3KIbB2z8Q8w2CAakL6JrprowThRbB0AV4elQ4h4EKqVbUoy
7thUr2l2u5Vanu5QU3bZPexmz+3Xexk9xg6NzwMBsfglcaDzOFKBtieP1tH8omqE
4WYh4D+9OWWVqMtxBCDFyJ67ltN4nbr0UAiwjfSSvXGWy7jxx+AUzdHitr4vK4m4
cC/WP5bkXGtvVMnH8K1mqZlTUZ/Iv9LQMIMauChenwsyDs2XZCUhhQ0w9qFkoSe+
ENOrc/LlgQNm4FQ0D8IYuuf8SA+mpxgWvu5AsiKsLMtJ+VDopZtE4eoQPxp9fPEh
4HJidJ3ESyzNA4JmJ/2tl5Kn7TCNZZ4GdmUPYIiTqTRDt9KlLexCQ076MQH+3Vyo
PSAqp+70wITmUnr/DN1THn94T6ndrmL2Ha8BYmZ0jgz991Rf4grPPOHPZzrzgqzM
hMk3YfsE54B3/xPPYI07YM4CAo88D3a+39PPvIr0YRa4JZWU3cZE3B7ZXGlwQa//
/QxNZRNHr7NCBqSOcmCOLGFvPVkgs9VMC6iJSWeNKzDigOvv9HDcB5D6VNkk6+/N
VS6Jti7ssPHrtDNAUZ+xcHehRhbIC0YthWJ9EyqukYDBhu8/c5IH72hG6rzbYNVa
2FZVR0h+DC/I5yBln5wMtzfcO7qdfnRWRJAY0myr1bNyDgKy7nZNrOanr8Qu8QPi
HP7MLe1AT8pDjG9L+P63KYPotUkrWlf0tAJXQKzyADsEZSKoqbGLfz6RNCeWH1n4
QQ+cGjrcZZN77XNlO5vFDdLdJQZuQiDUusjgLJDmeFDnkTiLIjrHau9YczxmkqFe
NHXSMaMOrjSBB2fx/n6tQcGaOJ1bDiFJXq6uOVV1yzUxn3+ferd9Xsqb9ahUINfQ
wPvkn7dt0gfV1tEnOs5/y6JlJrehDVJQWz09SCfSSYQoVx/Ccceg+/2t7tOCQ2R4
IPb964EEFaJP2fwg0tntrGxkiHzJ7SyCnBuusF0LbL66CBUmJ4H9D4Faz751Ater
ie1gyd6AfQpMlG2Nhn6h8mS53S6uJ5qudRtCsaUROv3XBMW6PczgZyx9pKm1NLsb
5bh04zhIrdlAKYtOLPRpJ9PFfk9RmL+Y2BaDswFt601nk0i1ZEXS08HPh48NdBtc
G390XZDJEbNWsINdPz1zfyRRpuSKFYBvXVLL7HNGlcgbYvCmYU3Ol9O9XpGBYL2l
qZt6m5P3ePL8rKyPJx/eBJ1wE5TRXADaJut9sI2KFRhXi3iWp3fsznF/C0+n3nNS
l7jEJQsTELdQkihWChw2XXkPEtjUMuKq08D4QWxhBm2XF+sVK2uuetcQ7KM2vxJl
BR+NrjF2QyVJJIlpUJjX1V8XxaNKni/yN2U9g01W/agVW1UFwFg/HnhUJXe7Rc4c
HZt152Dd0xZRqwPOZch5iYZJKfVdU2NA2kMIfFXSDWSZFgfUzpiZh5T8yaTe39iG
wYcLJ9pKHN+7GE6XRda+Mfav99gEDaGxmZ9ewROecxnD3FG9N9jIs7B5ub8cLilP
aCbm5fwDN625tTgaDp4FIvDRsyE9leICOhpDOZIwbQ9pgNhsvwe6ddHqmBYalAFi
7TaEl6o5TwP5J08zVmosdNzEuAR7NTHXDl7+6v9mV194G/VnZZPE9VZSkpjqN6X0
WOOrpdK17aBP27kcwIsEvdJIUpevCzW3qSofVVGzNaW08kDgWqhyU8Aabw6RjxUb
uYW0bTqNEEpYhmu0CmKsopWQKfIh2qKaGBqYdFE3dp+UMJb1Fo71ozekkRXm+LgA
5b7IBUmj6fnOhJzSm6YZHPK3kPO8Ch+XATe0VrUPkLKzhWRLZFLy4C4Yl+BoloOn
RCFnakA0FwzCc6mjcp9B44N37gMWZCqBVfuoE2bjAO96dQv4FdKZmzCiTNYRXIBb
gFfDiMU66WsD5pAwIKv0NPQrdHwCBgdhHj/AaDNAFlB2oOFHMYiGi8sKdEh8Rrnv
vf0vzTL7+EuSdowhCwQ1L9VBavbKa7kFYlKUqRqg3xIurpfmnITIDxeIUQWlgzvf
t0j8lHBBmI8Ul0VAX+mvu35XWrusWAeOICcbMQqglRx2DMHonGVjzLhHllfjzIlv
zGMh1gaMJXQRMM57HZWPVW0PVsAsZfMGd8JTINcfkkdErmln01kSAsVvqiOaYLWb
IWdPnAZakHV0bOnUFa1uGsq7DoFLNZKgD+m0bjyt7MCqtkvViwerUDRuD8cKoA0l
Q/mreZM28xx2MIJCKKnYOjpRQcMll25udjzJLwM/u2QQB/nV+cMPVGXR4b58JowL
XogNZ8eTi92VEKP6CV7kwbrCJCk6KTHwmhTL4pKYQ/yn7lkzFXIqz+wAq6BWe3NT
QE84AesCq0PbkYPaJOAYxNWw3niyrEg/0HquaL4AaO3Gp9yZRJ93HKFuM1GbvFiJ
k7xJkwuoohwcN+83tnxWMIZVzR6fFG1ZHOwOgNXXXD+OxEPVRr0kFOnpsFyc9nq3
wnVcIPFY9QiUqKwixlQ4C/wZHEFXc3311fbYBUWbmWs7kFr9PfMR4guq5giduH2L
MpS3LP8ydzuln1xFo7cngIx/Ai1IQ+uEKhnug6F11/DUJw11f/mZ/OwUYboGGwix
bmdBAKbYmZYYe+crtPiAavTIY85/dDv/fMNT/VH8uV0//TiUulRYDCxthTXH7aoS
/rAJXYody85hl3mEHZQtG44pJ9Wq3H5xZv/eeZ3BgifoBLeurB/+c6AMxfIY6G7r
g6JR40R6XMg/wQR8NVNAoGe4emURMyUrIIYLCe4lVBh751yUAiwLB1WBMdz19GkH
OSKYFMPKH560FqgisjwTvMz4MpfY9thsO7vbe2wcFz9rchVY6BXIKOTVn/HLmFPn
AV3PuXJN7c49P0YXZyWGAYNbTB2aAm7ECp93G5FyJAJRXz8AyxSaGKjunh7khG+j
lDAEdTGwmbij54ER6l64SDtve9X5S03Tpp62D6YdJ4mIxLNBtI88AkTuRUrrUO3P
JyQZhE08tXdyM7/zuI8GT/5/FXTaBJUm8CDfdXDJk4H3FSNyk1yIc2g5JF5eB8jl
Glz1WqBuLs8/hFCc+M9oF2ITJe9vDAv+lbHCR1QdBD8r7Jdn1q/df60uvDR/5PVd
gGR9sgLjq1EK87fz1MGDbNOjg88Ca3tYYCJgjT47uMo8qTtAZdq+tJzUxRwcSgEW
BKX6bGtb7yb60sqca/q0zHznyZFMiN9zHVI3M2NapIvxDR0lPxWH9iG3uYTkpSgi
y3Ts7Q7PblFPanBNdLSBVQl9z0drwA7fo4mmup1mMo+yKqcCvqhsjumOtBXYF96G
4w5nc3pbVgMF45NEf2dZFXF24rpnz0ZzK5eimXlnp1bRQ0x+vXYHmKKhmQWTxOIr
XBkSsKGPlJ0bWWR7FIhruPoA5GrmaYykCjKmZ67jWQ8Na6pMyzmh0J9hyhIxYxEu
KkB6nhozlKs3XiSuLTGEILt82SKMMxHQLW5oKlWEOrX4kBb1VwouDrYSs82SwqLf
OtvsaofomAco5iVA9wRp8tshovoSC6DlPMNVsXtKQO1X8OQkRxZXkrv/bsfSn6Zi
Ed/7RRM36OcmgnnYQAoAPCqEAI29DMb970KfQPT1lCaF6hDpBuNw1UEqI4Ex2YC0
Cq4KMaiO9iSwL2VXxwm4jX+J4lxsD8CJARPNX0jE2UQcaR3Bvo5ACcVw3LdSBJSH
7YiTQfD4wmlbuMdWoZyVe/H2xfMpKYznawwcXptWNdb3YPa7w1KkmQanHYHfRh9w
9VeKKsiHDEpRUnmnfDsS6PKNxFmrrBHUo4u2Ysu8t5Zpz4LaRzKTh5T+YZ5/QE6L
GxFH3w43KJgQwupUYakTzngoFDWW4ZSyR3OkQAuXABBKnPM3wvnwaaZ9mkVZmYnK
zC5qDyVuw3AfYAqWzwPb9EU73pkPA5Q3jsyt3m+SngrhmOI8bBttfG1Xi+qUQLxU
s1ALdhP8oCISx8uuph5pzAbqd1houG7rie5tWZJf40loTHpLjs1BxGnNb/S/PHp1
fTc/GBBfefiZGeWcXAp8WsxTbcq5Is7KA1BxD3QB5zAetoE13/7jnc9BFlH9DFkO
zGmnFjai95sBALUJn3ilbA3kSE25WGHPN3B7JnWE982KoGi8k2wSJD6BpP9yq26E
nGbXRRLob6i125XRyT4Kx+kiond7J8z96PHckJa9WumGZxvVr3AtItZ1TUMZ0CAx
htuivUMfCXnhw99obQuX2/muElaFZ6LYvrWg0lhQu1GHUCtquhll2k7qxardNIcY
9ZuFJlcs264FthwG3Ai4zM6US2krIbfZ9YsHwUrYK1Tqdkz6avaUPRR41QKTOLfU
mQh81saqArjzKh6OYhd0lTnzOELjpygijtkh/29Jw6/j2kuI8pXjEk4jM95uJgyf
kXAtEggkPida94O9wAMjz/WmoGWmJB8ba2AYIsuttLhm//u5TstTOBEKgsIO+Ork
8lsIihEnyFugKY7ZL+H3aZ9MlDTXSMx9aZ/0NrVV5Oo8RZ1gJf8G2LyaklwIncw/
5TYxl5/nabpJZ/SGEuh72FOtf6Dy9GP5606AYoYKgcjX6VS5544YTBjldX+x8yyZ
aN5GET87fWWG6QkqdJHBU9PphA7aEZy07K6t2c+2LZYRRWyWeBVfYIf1vfyA+IWZ
+Kv9T+lllI3DU/remY4YqFmL00DeAyxaj6CoUhFYPzCtnq2RkCRHBj0md3G8KByG
tOa9aE93ssV2+wHK96LVJoW7DgUbcV93quUaBJSKVAMrEF/+XiwIagcbicaCf6fi
2i4dHeGhWg1AMLAjEwG7WGm3SL7TKf1OMbVVx4QaxtjziIX/VFm6RvGktwkjAqV+
+wsWSw9E5HVuBI0UJCVB9HhbIdI/2+w6NM5+YP3IBTo1ERBKQSOXXsFmX/2ZyCJ9
NftyIqz8sTZEfhyvdZLl5h4S9AyCViqpFQJVkZWZ86MGGitzKKfzmIc4tBgXgcFu
+LChYRGaYhc81d9k87M9ukFwblQvQniluE2p4mLTo4oIAoNndg7JQeeZSyjrI6UJ
YucuJ7tpJairk9CgbxLCOOvQ3S3DeLpu6dMkvk8wR1a7G9Yi7fTDardqv5x3oieX
p6ounwiYUJrq9eOS2oLzaXtur1ge1G6gFW6sGGr8xPUHx6BWPu1L079MUtVGWNjd
i5oflbxx5A8fjY9QqfbxxptrdEZrc29S2Pgu+Xior6163Es7iNU7nmL6YBzoy2Vj
EaVPTGuXsFE4433wlZ94fwruFwem8KqobkC9idtvMoFn9jLb4aJrN9XwDY1niDDJ
MUL940dvlOKEY9aj0Cd/26RtOY6KX7Ml3loM7CKXk0A5HJ+LAQLFKbRmN/nGJwIi
Ct1j2bdTFH1udkBN4inG3s/fsm3Ox2t9j5Jq5TWftWrsroAjz60+kjzXe+VS93ei
TbgzVk/NCJ40jv27lrFQYfrVNTibnskUxjLuhYatTIqVUG/40/JxKNFc5BQNxBrL
Vg3ikLY5Sa1XK4XQKn37BRRARNYOhmRUZMiHb3yiqfo3/qlvTgzw6f9T+pcEkSDa
LTp/0XH8ekRZKc33nwtJfw+UMIigipYndKJXTJkbLe+eKEpA5mXy2xcJRU+SFgzb
mWAqyoVGCJQDw313nr18rvxgs/2xKxLpRriIwZ5pHpZTE8wlLiZh2JYkgSVkQXRr
f6KzMjJsKbQz65nHpWCHlbTBqhAV9hwB4337HdZv/MSiUYct+57KS6WYIx7JM4yK
/4azW9n1UdFu4WgXZkrzWMdfcN/Qtq5GnrbRe4tFuXnjKPM0FFcHtNZaTlX6U10E
UhzfCJB2g2UEhHj2ijh+cS85n0IwqA3O/VDUWTiiNkDtzHv3w0PsKTG1JEs2vMhE
0mG6iL/CR4DTOUHT2HEKAVHro4IwlauVaw7ICNSbBzZQPsQ49SuAWWS0Nd+y+iAp
CLZ1F0/FHomrMz27OJh0GccEOqVLMeyGinURstvSuJrc9SqK+qCq2G6es8vzWLT+
EqZX0Pk9jXYog02NKwtMCFHC3Mm6166QTqq4IAgGiM7JuQnpAGmtavtgr8jIJfD9
QHUV0wZroEDBi4GzFSe9w7+d4T0mdlxnkImhgMV+jmbiekcFtne+KcyY54GTZS23
te34e2RAwKrpqnRmfb390x/H3M1pFxTv9jtNAKC5VqSD6tqCgfOASo4+4ludw3nH
Uu4KWYsRRlc4R5SN8l+D8ekuJOdms0p8kBBpyEiiQjtHu5/kJoWIaByVo7DF2Gtv
nV+4RF/0QI8bnYNLDmlLPhnDNhLLkm0m/ltdfuKADJ+yCqRxMuudqYHPR000R/gk
ko0WR9x1qsM7/8GUOIuvhiIireD1n0bzhOH6E4ADRMHS5NwWUb+WJWpem7VLHzEM
SnuNbSLQB9BhBHoPS6FUwtgLlNWkcNW8mEFIKfFoSL+B3EceYYu3JVhIPeHQginU
S8ZUNCRcPDTtjDlB52jnmtMNqEPLRpjxgfMxgf5zRzp3r/OPnuSyHPV9zxsdkYDB
kUtBamz6IyJ9Idt1pdXyPn4PjEw6mZ2B47ruuOrbrrZ1DWYwRaksxYrxftgP9qf0
b7TXhZSROqeX0GNWREEfPW28PEg+auuoQgWjuMMYhsZP/zSvCmJsISKIBU7ZgKXn
B5UNVffb3rl7jkvbHm1jqIwgEovDAlSS6gvtoQsl6v+RpI2UQIYF2jivRfQgLqun
YmNnP+MFPy14NHGy+qORKfFiS4PfG9GK1DC842O+G9Sct/Pg/Nb3taTu/KIYZJ+9
FoFO61JIbBDSjfDQGio6WvYY1viR/FofJlwmrnXj34uFY7/b5ZP756sr+ajkakAY
3hC2WoZiulYd9QqC4v+DbvWSIdRo7eJnEMAfjO7x510WBM3t0TO8vDg4S3+GRtcM
/Q2KU9UMlE9lKPJ6AsXQ/MyQ/kNVtglC6cNq9si4kREwa2SQXtoWWYOhbsMTg+pT
D7Mw+kX8xveAv0NWGDM6wUhaMKTFw2PEZ6CK+ZxarM/jKWZmFOnsdqIKh0kyMJ/B
UtX9USAterwAGU644lFlHCiAA+DH0kTucQNtlTttU2N5cvv36liBxglZP/PAosTK
ASQWGmTBAUaSOnvQa0wLokDalsxl0NrvRX+6E5krSltqYvvUVHLcDUIjWC8h6OeC
0088SLyfhXgjL2W1MGFt+4Fo2JdT3StmhLUtStT2kHDo3UCUHxKkalL8u9ncJWgk
yfVKc/UOL9ByasZqUJrwQQ3UmF1f078Z15nE4DC/jFRzUAqkhMr2/IzSsNxRNLEe
Jb9QxSv1UBTB9mYCGNMQRB1O9YxBEVyaip81z5jJB1REn+thb9tm7hZnssOOLgrZ
b5mWOQ4zNRxsn446FxXdVzfbH9GEg8lc4mgAL8AF8Uj7Cjm6Lg4+tcyzQe4j729k
V/A6AZy3XV7cuVUhctg3s6jBdaendcXxDVKxzSmWBKWY5uUQl8VAl6gkhM320yNN
EJ//eKCXeukQFJ8PUPYYcupj+k766PGN3HNSSICdcXDbeRUhLG9KI7SdPUr7NZ/Y
0p4OFyvEA4pG25LWfz/7WOd3lTqrM9cG+gM07w7N5hLfofm9ku/J8XUndmZblt2y
P/XrzMo4rzL0L23510XvVfFavoDuQ1Wm8xV2JJ/TiCJ1Tp3SEGTwu4aG4kangLcp
3IubS85vVx1/F7juPksq/h/GrLtDIdXjXTRN9oZHybVxaJRnPGAQMmoSfD8U35G8
woZPG+DUg8Ldfxy7C478bsNKODP6fUoTdsxrFDMcdK7YhIx1RDTxdWFeVy2PItlY
ctAw3cYBWkda1Q/MNAaEyNNIY8zUOudI/lXbJ1nxy1CnhXr+GHrSag1jDKdT7Yeq
npsuc5iyeGuog80mjoNF5nTphrZ7rFPWZOu0rz+mk9iWkQ+a6SLgFDXX6fyrn1dO
mzK5wJhlwi44PyNAOZiVrEiiPqTpuz72vtDZ/wDMk9E2RtQypo+h9Sfj1DeBmRuk
mFdsDgAbnZ9pTRqtzu7skKR/UjJIVvFMRgoDfCy62/Bv69ZX6G+3XnuFCdJ6ovof
oaa657uN+e5n75gkxumO6rhpFTHblpdZH9ybidwrYZz5SNQ9lvKUEWUwW/Q+yadi
W88POQ1I4ZNCqBrUYFvNzUgomhpABEyAxVwz1Rw22yrsGujABS/autvJPG3bRk1U
dcsrcFXUqwD/5/Bahzo+c3iAAi0MFDIy/lQzKbD2mjC/EDwcRK85kpNznz3/82Ns
t0CEp6fo1frt42fL2+JiYFzTQF6SH/lmTYcpltKT816R2XIM9L4y/5maJt9xNZXU
WmbTHUlygtLX8G65LeB7X6F0ZbB8VKW8dZMBKQUPfMyx/KASm2rgHG1OcwbiaLhG
2Gnk140ElkLRzQV05/30y1pwGq59yOpIsMvHiQTjnhv20VWUP5Ojp1qE2siw462b
3ayeUtDRAE6H4Y3FGt/qBArRqZnvX2nmKcshDwoyJ5i855gBaYJhiyxLM4DRcEmF
85QH6E5p+Gv4ya8sB/s5f26bCPQkWLuaXokpokIXAS3vgbxbPjDxSTVALbjsJntT
1IqvUdol67wqRhwfa47lnT7eLguQTmZFQQ+QD3VYc4eRBqBoMLPfIZmQBHgSbt/m
9RTMzVbcF6kNLsHfpvlg9mYhIMx+P01n/p8vxLcwhrjC5XjKAqyKK0Nx7bP9hxUK
2GbJuJedFcLyrqkpJn8iInRB4KMIkBuB63xsaMCpd5INWIEiDmqMAPxTsdcXKUOb
CpGJ99uvNkaEcus9XiSoZAItjxka6fVllb/es6wuH61z/thKfsidLKCHOepHGSoi
X5ndMpssqFsNPy5WI9nv70W+x+Nes/yxlMF7zo7zsR2uijJ582UQNRDk4be7o0X7
bOP9wjbreQsSHUd0PtgfubqtIZF0eQwJ1Kqe4oPqjJQVFUTp3vrmcUe+Paj3D0n5
pxuXEKFg5pN4HIxclMh2Tv8pLslCsmtTJs9teEOQCV5uR5S+53vhISMcAiHSfNBU
q9JuvE5ItKcZnEkf0/2FMyScVZA9UbBsz/9SR1XUvSDThA9USZCbwdjqKmcFZ5em
MGadAJuvzol+T+Gv4aexHRyxljxChlb8HoeTSzNwlOThmhSWwi0vxj5sXSLy2hRP
/jbu+pKjkPznJU6GQA+FPh1HTkzA+CcS35LgzaIksWRTSieCxdLAf5Dmv+GeaPN9
jt5MtIOK+MudkK2zLoUJruD7Fnn602mlUzNieHuiiXdM+HgrWgm9j8+NB1jlFnYZ
uymPEEBtbqxok3Z1QcF1qWPii4eP/cIxu+xDyc3XuBWIprEGrD4hZr5g4bCn1Wr8
m3K6cu9JYlY2O3Eouc4dH0uT7h06zgd5IxOUOcnARU+JDHOdLYPcosHbdDhezKo0
Putb2QevKIWUwIv8ukeVCyNHZUiJqbMAnojmUtdGaQrdDjpJDOIR1+B7uh1txbTh
F3mUiBex4tGACVKBlwHFD4mfTQwmMuqbxIE2Ubkm+pGT+ttka1xYBpD6K7D7DGuH
nn21WbfCktj78s0cRxrDDiGBD9ReAlpL0aNPR+ixDwZ0/CZvDRGZDR9x4pw5Qp/A
VNj+/AODJGXxKdamifYYajG0vImh6b2DLOgCHfayW/z+EPkjGBgXzGh7lewrFBsf
hwdilntMSG1iDLhFSKAVXxricePF9Klk/7wxI5rJoApPDOeUS9SSSeR8ncftiWDR
2GjUxsPX0azwxcMuEw9tHiBYN6HIc/vqHIV1HwJ//xEE0QVa61KsFnRssHq4UNpF
iGE19wNXPMWvDoHBHfXvh4+7TyL0jZL1WA9WzFz/gT/WGx0iISK+jlSiyZK18CEC
TB/Tg1J8iEeE4D+dDF8NwfSfNA4tZVJtAULxcNXBSb+7lSUgAiZ4cTRtgG8WjqYD
S5d5TV4gv7dJPV+zE8wZRlrreoO2pgKsZ9STifuQYtEWKB7XDBGgjRpVPkCDeocW
ZZsoj3JcsvIesWqrufAk/Xr/V/W46+tc6PVK/tACuNm84bapN6BbgGGct3tzX6A/
fvEcx7Iypk7Dp7aNP3sCGUVeChrRe+Gx6VAaYXHolIcB1sarPd8ggz9E/F+7e2uI
NmvgBa/h+Nrv5R40VOjFae5WyT3K/Qw7kBNj0MNmIOg/6RhC8hLa6saOxHREOSeR
8pAQn6NtVsz03/DAvdCdXJfK0NLyl8a+d/2q/DVDJRYe+pE0KXJ0u4cTyR+2nLUL
vpONhZTmxh/Ljcu1a1TUPIZz/yNOAusqBrFQfauOnIOsr2IEHVMtdbIGM6bnMPO5
5WpnTmYDtil2K/5ydT51v9MP4bEZ+sUJyPvqGSwyYVMRSZUibGzfXUY3lDyHXVsJ
c9JVmhiKpt7NnclVxpbswRNf9xu0ziwrsW66du7t/mGh/jBZpTZp7ojNJcd+xvwY
BMPA0Ebh06oTgF1fBF+OTJB66fE+FHaQUqzMf0aKuyjsfUCSrDmTAN11k8JrS8Zy
/lzt/bYuWlJzJOLKCKfR6OxBHH3BiQAlxrM327sDnhwDEcfVY5H9Ahz9PJjCU83B
ZI9BElRK7BGzwmUzjnlVqmoblTjORV6T6tSO6rH2gGL37smAIY4KSdV1IkZ6Ngh2
uRHHsXH2o1hnlAL/Y51BYroQmvmGnf7Rd8+kVVBPBzZngAAFMwVGn5c4uZt588Yr
RyoyI8xZPl1ksdr6pOKzK4lMYir/Qk6MIEvMzHFQIBXYP5tSwlcYDze0FM+hJ1AX
w8ZuShFUYaA+U4Ee8lYqpYDznw0HDChawGPp6wBTlLPgw3oyPDIGFDSw2s2LgRYa
kFJOvMLN0t6lXFGkMRQAT+ngY096jUZVKfRlcdakEP480XvuNP0C3GcD1msQ35tt
7kiZYE9W7OkClv2IzwPv5VegXi2N66D1tVWDKdOqNGeWRCg/X7RNvDTiSYd7A12p
ipb7BaBKbyci8y9zqG2NO/oXbohjZWHXZSDL2uMfuywWIBQzKGVVtAtoqCGWWsIf
89jLCv1uXgL1vtZ2qjWkzVoY7AJcUrMmN3BOsTl9FNq94YiX4gbA5N5by3HSTDZv
0VMKbt3grDANEGE6WjKU4f820PJfN1QI1+gNMNAllBLGOQI9KV221GTmAQO3BpR4
zBwZe+8GK6gR8WyJJgZ3Emg/piBLw1PaRFi72Zf48jHgAY/Sl0Dn8ZV7vIBRXOLJ
4EfDJvM3KpGymTFEwmSxCN4zS6Hn6TotIscjGvKas5HEj6uUi2e9wzXhM56Ch0+W
07aqENDe+Gx7aDqQJ2PBMkPEHa1tWC9GIq+Yk+gZZyd5CB/nVkReio21xOOuhwqS
VGPFe2xnGNs0DMRXoFl+onkDXF/mvHrKiFSE4SegqZYpjJGqJ2UZFDKUjP/F7oMD
gmiDcyf0pk2ECKS1nwtfVDM1DhBHppqsiFfzpPTM/DCmLFmJO/nOYf4iWrV7Nsf1
L1enc/016cPWk3VlOwzQzKc2uggQi1PxuXPGqTkwJogXjdtv3VgdQIIXF2v7P3L3
UBzO9Jr6JwY1WC1moWyldX7BLScK8laXH0aPmX8DRW9v6mA2c4srqawUCW5j6Tal
opqOjOQrwdFIjzn8CEi0jP+g4Q1N8+GcGZKFezFOPPSU8sIf5k36pxTtchlWBxD9
pFHpv+17KupYg5A1IKKpQ33hMxm/pqu9qV7M2K8lSrWLIuq1iJyQGMgJ9G3l+hqo
1xTtQ84ZMVfm1jPyze2LaRn3TRU3QSqdr/+qRDbKykwli4vnnIVUsRk2wyYBwn+d
1SCztxKUFJF5jfwU3KqadmYfS1oL7OgcvQoZK/jxZbuGDL0hjk0Pz26s1hWPVV3F
rnaByab4HhvsDfgj9jqQ2Y4DPNFe1+2ertryDMb9I6r2JIUND99PoMib/OobCH2R
mLyZObHWCtOD5ZpLtYnWHhNd74H7Yl36nIy/l/4bzSTYl64dN+uB3tll79rEsKh5
iHLMu5tPHT0mzZbM/WW/E4WacWVYaeM1/pT+e500/IVyPJFxEJXM1RIXoqhnoQM5
0m9B8NYVxubuUn/QwrwkTn7faXDm63ecmINMqEwerdJF9qUWwiimGhF5PYCjrxzX
6UL0/Pfo5SSL9qCWbwskzBszW+l/Hq7OtsFONGQX4iQ0KDzHEumoR2KQKjXb70dg
wVbv4rUQhlV0ImmAiUcFMKaltiUJpECmfO1xM7qGWC7VV45acNlBgvkwv5+h9rfA
+IXOzzCCpi9zoPn2BXgHsZHXGCSzmnqIkPQZjeHtvBCPfd8W2ZELz5HU3FksVMls
mbIf5E0l+2DMsuQuidUpb+NN6GJdvGltWFx8sQYrOAwc3y4C6a8R9PMRh67tuBte
7vNT08ggZxym/BZSAGZNndiBIYW2PqeLytSbzEm+2uju2BpM1wqu0CCsmPa2TVMl
eZ9qJxubvy+ivy0PL0Rj/wsCJV+35DAnQNpjZXtH/gEC0gKfWKx8tiG4srJg5Fpz
dJxhgzQryTHzl5/icsi2uNYwnp86MARnIZOJ/xoJRCCzvIIxcsilAJd9hF+3/VUz
P62+xVYmnEdMXmYVLY4DjmEo08H1xITZ1U9mx42/Aa7L4Z3dc+CV7o+p2DeI2En7
N29o0cvwR5soDPcdHfWXcYJEs8cJaQS0kF4CeYA5WRZCGr3lDPGHHSrOz27LRCh4
7CddgrfFY22mGQ3MPfOrcGAFXg3pI09OGLyTi/v7gcbpLJZL/rr3vLyZctFA93Vb
vw3xAlailXOh2XZ1Q+9IT9LWY1h3/BoeETIYv4Oe7QaD5mAIQPaqc5il+UJ0PR0B
jJq4wfQ68Cwnv6g2G1ChkN2UmGWTE+I5seNsxnIRTTNJO7m0fbTmnpLpLr7e0wOq
nPl39juX96+OVGdzl5d+hpPNRpELrzZVVtCOEEa4NMFM3m5OApv5rpQ5ikM83URa
M1+49e6KoxM2rgnWGo5WWRXfBNIPs3/qhhtZxAvY6LSPTXe+h2hvISXXu6Se1Sbp
pjusbVsVfR+AoPS4ohhtVq7skQHaKmaYAMC7iZc6OyajrXzedWZQfaLc8RGGhWiF
w02hXnqzvVYlDZWXANIBJ9UasyCt4hjkJ8LMvefy3Llyd0XjgRZ9LwG9ytKeq3ph
BHPPfxmMIotzq1Vnkk6yAVU51GFVMk+dVOoIbYqdyP2UXk10A+7v2vEwgAAsHzAD
+zNXmwjHWI/vgdIgSiASnUxbvE8cvyksDFM2Zp0viAaxSGs7y3UdBsph3aTf46gn
nv9hGr2mamrgew7TEIefJ3BwkjcrWmMx8dmEoyQgsqqdPylPPHBF7/GqpMAM9tKX
N7PKSnUIL1Im/U13VnDOHDgaLuY89TsyEb7J36aEQRZTI2DO2tEhqyDQn8IoLQrR
+rCzZEtXRUE35VVld/Fb/9vXQdYGtHWKd71OPpA914nngis0zOw0rtRkRZWlvYK8
kYA6xVVaWtBN2DuesQrfQowjy5ZA0rnR8Brr907L/ailET2vA6TjjIe2EeVNFXPY
IF1CSn5tKbj6J6ekrGALdAspolhEvNcaXq8S0ybwF8ho7ABKozMCpA2pXtJXAUju
WxmFiTYeHkYJT9c/k4rinNezK85Bxi24D2cVnak0gvNczdtRDPNrC2ZeNFV//Y+N
WZ4UZDrx9iMw5WG+tXCpiqACk5XEgGITYONHjRnMbfoo1Q+f+r2jaEk4fWPmXNk5
14jEbkBCehSCjobXfdIQOBFim90EyAzfqe9gYBjjwGBWkW9J3ZeEopw/bJRi9S9V
OXYMS9zl0QkHRwjLBhXrlvyk5s6aPVFjG9KsrPt6pakswh6h+GH4zGTRHMmfrWhQ
Oj1pqO6PU/aQal9hM/dZC8o6CGRoGEA1J3zmCcC+V/cP1KK29opw9g538LuMOI9w
YD30Vuiyvj5ujolQTVsqOqyCBiJ74gcYcaCYPtp84F7zL3yEQkcYzQ3bC3cuNajQ
7xbL8su11/MngEqrxLhaoFv6fEy0yNrb6cDGi3XRiXpv4Q3p1KlQy2O5btTRAsCZ
W4KHRYyAP6dcyBftXt3Rja3FTGQKNrSRkCd2euz7grTmqFHpTJk7ZS53NbIzszI9
HHUGGtHLx220r6kNUwtpUnSozl9vZ0OjPzCJYl+KCKfPGnq+JlEdfNTEmPmLvmbY
ZtccR6XE+mCIPeGvb/25dtdNljsBdkkZQrxojjv9FgrpcH3cd+Q+TVDR9OnPahwF
BVYN7WonesENYo/YI4cfp2M/nT0FUlGccTVGxmHg71qNuPi4A3Z10ILXIOrZw/kf
LoD/ElTiU4cTsvvlcpvwQiKU+j0UbUlII3s6zp+8Qth83misDFKTXQ24wL2yXaUA
RKMF7LXV++1XBcwtzwSEooDwD7p8OFGPxfvbNvGWdWwqQz7y29ZLaRm4y/cVds9f
SXBmj171w0Ge/KMT1aAGMdov0KZ4e3iMZ5BQWmW7JxnkwaFl33ZFGEs74g1xu9rz
Ivq+6pS11FfOAQHJT4AIOmtSg6Pt/haX19hP4DHJkK8VS/Q28B4QOoklsvHkhqDJ
5eo7hGXXKnAc1tc8usKZEbD/oyHcrys1I8ni89fvuCJziR3pMVFJ/J3cgEJwlJtd
YgV3Ik1nnfqe7U2MLROqcUMf8y/+yJAnqA2HhgBCiryoSyskdtBnjJO4GvH+C7C8
HSAyzmzVHo8RHhS33LYyPgEafgYWQ2FxfwOQiSJ7tA/lpIw+OAGdeBegWU7s6GGg
AcwkMND/T2+x3N+Rk+df7BYeg7FcSMiV6oWDDEXzrecBIIbCTiLAFf1iA4UQY80D
jbxj5XzZyILoSx2Y6ljMsv3WcFQzO9gnq2w+4creoi05lgKedCamL7F5l/HsXkBl
TFvFj1RMsTFGElJrqaHThJyR83+lQSY5ZUkqa6CvLpSyrMc26l70pQubN9RSBWvK
7D9pz5sySFKPtkq4J6/yoVSEYV2UteDXoLMiWHRWAM3VpE/Ybe2kxeH4YVEHea8q
yIM0jAJUb274EOp77mrL1YqT8FAe1RmesITZfAQSMV3Wot+wB8bw14IIYMVjfaPt
Qsv8Ys9U5y2aMAXrwCyRTa/m7uYsTP+3IcKSJZgWvtCJD/+/osgYsUlDhBG3/5T9
Ev7d7G8rgl9yKwb/tskuMvJXwoVY04P5dBkWtj/piUskqGFgyYnQStSyccHlzD3B
4KP/iOS9yuwdkUae2a0IOyjUtAT6uuCALQOKhVXrJ5pXjrsvgqVAcE97YE2vBtGW
v3ylHJJWZv9HwQa3m8nH1VXG2CvdyZtXCTjpmH/j6CCQnxFBwYUxR2RL0XoUO7fz
XAco3RPYyFQwm2QTSZud7IDmqX62/JHzQmNQqfV7vFRLEm8KZRC3eLBF1kBojElP
pPc9Yy9haRGNZSWdyWTY2xvTObEw7Ar9v7aeUDhU44pOFtT3fzJoIfzD3ok1bjvL
FCDADe+OIucnY885KAXa6PJ02fhl33ca1QHi8PIHI1rOi4ncwOpNvwCCEZfW1uxf
ysnI93RgWDUIk5ohMtUXhpkmtmiESRQLv49+qP5BdMa3NoDenJ9P6n4a4+C9EHah
OEb9AvGBn011GT8B5Zn7pMZfEzBvcXj9RmT8XONeX4ETSEvmRZNJWeXBSGwtXHZb
C51nqdDRRM6uqIF3E/zt9OscZix8TckHjNAd0MHwdu33HMV06k0vLFF5hOqUm+BN
0np8BOHtkPLs57UvVmYz6/CprirFpcG6uHj9Vm8BS9JJHFPcBg9ktrb5MovbktsS
xJ+uEajhn3oalIXLTeywKHHXBbIbg/ccVM25xqDfcbBVNYY+baG8v4D/jKQqWFRh
RvSKlBFmz1bcEV9o79O02iAvntJ2YsRrPpEhUWweUlMAk/Ze95+dhWReDTY0eAVT
X/+MA0Yk5DQzZKVXQisVetkrIlYZHqpKEUcTI7uMEaEpZIVkl63WzDx5Olgy9MQS
gsF8kpHsAApYSGRE5rQOzX+l5nZYrjZNJe21mDiOJls29tzG94POw8VBJ+/yK/Uh
xQV2VPddEdPy1l3sGsvWy3Gjj49aNCoFDbXq7oL9bA3/nLo2QNc+EqLXgF3yXAL8
HA4iL7ORS//7G8vQh1755AIKJlohOMKJkkm/JBG4gRAFJZWuX7rHNDJH4wMBXVmx
JzAVh/2RLiPKr4kaZA8LKbmYQr/CUU0V1gBmpoxrDGmeZl4mecWnjqO9kp3XcZvd
mPazU4FSk7wOs5f4B5nAOV6eIJnQLBoWgcjtQh7TOT5Hli2xAmQuo+TKcp68cImj
9YauOBXs5bICANZ11QnyWNSWbvdg9N1lrQJ48ucovgRMnHEQ2KDQje9YibMIBG/m
cs4kOPTEME8H+yYRGF6jQNvOs/R49xSUM0g7jV3xfYyUzwDuxMO8Yje4Hki97/XG
x6kE3bM6bX6expBThy3ZV1LHWZnBPysU1vO0TEr7AYvJsNkdVa5A/ytRBi4Lvv2Y
HtYB8NVWeikh6MR3ZxK2DBmSChtD+g/loNqQmQcTwgOm8ZjhXcGxQT0gy+l8w6ZG
l4QBGiZVwDab0dCN1TMmh2LAK2aGLB//GvrmZbVl4xcqRqfUh3reMvZkq+MiDc3J
AGquAMAoBvqoiR1m5OZZUKLBUqmcNtnr4wLTLj8GfSZiI4b+UzLmPwcOxvqNhdz+
crV0UY2Oi/zgtngHObvC5BXFhOiyOHGerSz5w6qnYL4fesy51nZ6NMhp0lLASYz5
76B1fV790Tz0J+LnHImuhjOiw7Iq0l1ym0KltPLc/Ad8J397zEJ8vBrGRgMuSCLZ
Me7OWp/Gry0fWcibGoUBG6XuxUbA6xM5VrZaaxw577OUGVVEtHSg4WVghmGcUpA8
XcZQLtDdBVu3tc5tpI3QnA6yB0HfvwtyJhrmzfCvdzpGa5HLwAVRJ9l5dcNcs/xG
qLJnFlCHol0wGygb90dtI7dtruJ+G7gFh8BVdksBQ+sWBLCG84Q8NJFExT5CzFnL
hnKqox54GNyG7SpXkA3ohVQhLWe2evQbNLukkV7J2j84EuNLh1bh0fwA/xUAc+n7
dWU8tk/DV6Fq6RRT392B4PqH3y0ihzSmjY/NBle/aK+oF+89KxGeG8iRu+/zcyAA
OcmqmLWWcvk3U+/n+NbkGniMpydbJ5tRqgdgSa9BHRKjkBuooPB9FDiCAm1agmAS
GwPLk8KmIZUs3OM+cw2af2/HbkYIwRav+3d/+HIgJ2iJ2nkqa6DSWhirxB0U9THU
6wMQXZS/nis6KbQ8ENa+7XMhrhTMsM7zx72ybGC+kQlM6c5j6Mf+IbkTEwBgQoPf
DVBXbyBoGidoeiOA5A4p4LT4cSQrEr1ScjSTm2SBfmMsYJqOzIB35DxCQeHIvU8/
GE87igcJhmV03iYRurhX5d4fKjWnqzQdHpRFWkbtBbnrsde1V81M+Ce0Q9Zkotzv
wi4SjLolQkQKSZ7AH5f8tv7pO6Dr3vwCqDHEOQC6hZisafaBWqgVGHO3CzhUyKT8
qvIqOYhoomtmjnFd4vqv8Whq16GklOvRIpNaAcYUBkGOfz/W2Hlme4b39JRuL3GX
jkd0X5nti27AeweGNA+w/s6dat2qTQQUujjzS1RynmXmfj+aUR/fuEuOMIBYf6dj
QtZxwu7+NBRmmt5oml0ltTxGxCG6hwP0rbMMyIY2+RFNdeUXaoqPMeWxna4h9iZr
6gLQFa3c3AmxcDvl23xmhOa1cj+lhyPWlXCJ6hsPf1gfxr7tTyna3AYSKqde5kte
vnJKC45qmIklTpoHcfj+JCDTHOvby4vR2z//8UAOsNLHWa7OW5Rue/O7YIaWGBbq
PHcapytaLEd4kUsLcq9Bb2b6KkI6QTd9SzYZr+92iuPzX9TSeznEac632duQZ67p
nWCjgY2gqHgLCQJ829jLfZR34KLiAUeuFkWxAj0bvDMXxXRaUQu75g+ci/Yb+bPA
o7+r6pjo8VB1ZLeynApFJN9jugZqSmIfCsEOxWQy8b/vtIzAzsG5cKg5TIg2av/J
thNodIvitQdNe3QmmN3bLvuk2ASjSlW+Yo7qvKS0LNAG3/TE2l6AWvXnF26v8JgS
+t4J5QBUDhTHcrV4TJE5k1Xv1dSC7R5yH1r6zaIZ2nXw2cBH0yDb7bhdysK8GQyg
6smkhMp+8TQfAAqs3xtKVaWbocGLQWVjUilljsszcke23BPd9N8ZrHeMN9WaFeU4
MsX5aa+sY96p2D3rSn5N2t6sp8fIbYPWHEOr7Gk/GunvE3LTH04dQVT/6bbtMfxN
xBbiW7PqFH64TqbQCBVZOf6TtnmuQHEN3vlms0oBpTjaixJasqqxXre5JkMWuvxq
+rzOJcnULHz7CpNnMunCElsTKxj+nfZ8gDJl5hD4BcWys6dfFJObULdpbKmdGalC
x0gSDzliZ7/wq0Lv8ySPJUtM0x54jXsl+p0gzv0tP3PmQVQ0o2rzPdsvllGDuLeh
ut9hHPKyzHhg+LWMgjOH7KptZVfrcHIXfSjxi6CNLPu4LfltEHLbLqipMj7uePW3
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
b6orJUzQ6YrqwvBAFMdiqS16ySlg3MwSHlf2/YAkE1h8EyxR1JwSCnohtrqyv8Ro
FPKELPlFvJ5FvubfEds2H7gaRKGMaDw6VHZ6b7oRijZExTlYvtsgHXPUsDLHB4Xd
AVK3KXyv0E7SCNVuWzRWMZJflc7b69jbqd0szleDYn30K4a/rzmmsS22e1Ctxx0s
ms+Hsfh2t1E6j32ttf5YwuxZpyWnBB8HvKpNLOBgS8rB/HDkSi7XE3K88MXWFLBm
YysyXBSGvOLoTSUSbDC5kJW6n6h1VyCwWLu6PdicdQ53HWKfTkDXS7qxi90Lc5Ev
lMU7j/DeMBS3l1N1iv2Fnw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22576 )
`pragma protect data_block
Gu/xMgp4H2KpbTXVL+5uN1ViH37X1U59s9P35zLoFhfY2PBtZLW+clyOKnflIzYp
ftCDS+OPJAKkjNrOITzdS6bZhDfJ/5g4Lih8zq3XjTUhEobtWVOeAzNWW8CWk+jQ
VCIJHF9qIG1cfi1gDj/errOJzjqXvTqgDmF2jidaPkSZ5wjcI4l/MO4Cr1nwVKc/
PagS1b5i0CR2rUvovoKV8DsEZSQOSR7OioZvpm4xO2LmQ7TEp29gZaT4/LiqXpxf
ZZ8tctahBfAW0yQ982ZFR8z6mYcOnRI+9ANuXCfV+xLx0QZ1ttTK912oDXlYoABt
ILeiiSGZ2ItYqBYNXcLxLqvIsZHyg0o6vtQzwPM42pGnwNqSa7us/byyrENCDeKU
8sa/vvbP9O+zzsVQahN3fxJ5J7xOiJJV37J6cSI020YSyGDyMOA3gajiWetXbOUF
fL3dnr+XSCjqBKFep2hBkcO33J1fru/oMROQ5rifJJyRAjVx6RE1aJ56OlihbBHD
/ZPogwaZVES9+edqwijQJnrgOLUrlSzmnF/6L1K8WZ1qGdMQqU9K/zsBfHyjKij0
wpphesz/AsNrqh8SK2KsKwxWJei6SIQGquB9rlxH/pO/x/Ph0aSq3oOnewfLY4bb
tAWsm0ylUjoxIyoOd4ok8U+hpfDMPGZ0SmKMTdntKQVNNKT856waGbJqC0cy5VEn
kmeuAmW+fIae+24wzXVTY/WkTlLRrTfTsqhBNgB8+Ld3ZLfkKGnYr6S7GcavIM+Q
e6jS/hICodXs3N/U/8/JXG3XvUA9rxpiELXrxi6JtNxPFXeCbhC8sMhLktaA52zz
vmcG+HtbBI9ryDa3B838pXcYtUhpPqQBuDSbnQ8yzjJCxOxi+TUAjlQWQ4mqBx6n
mW0bjoDbQ+bGZbGrZfRusqAUK5tgNVpNCvygqskCpF8Gd/QL3uGW6YcpwtwrOXvD
2uDpWO2XbXgTtI5r+NrJXYO1y2F2QRa+Dt47WOqcAE2dWwIR82Z/6Ie7glMcFhae
Eb2Yo4UQC3XxIVVzeSwnI8egamURMaXIruw8e67j0/NWzxjZ8qwvQtxHwu/Xvtez
lQaiJK3Rp/ksIL4cbeAdxm5xjdrruq3csKofyVIGsGW7ANpFncaLt4PvQqM/9o6v
UaW2cdRwRulQ6+fnlJV6EYgq9A9uf/JK36syuzdQHsr/dLdgNPHKQNsN3yzlOpJM
DqwPXdANKubMTlWN2ahk0Ixpr+YS+pr6TyZmTG2uZdiFSinYnupZMCLWyJn6wuGA
hhwGmLAB0r64Cv2QwfQQb2/0uzrs9D2vlCZ4Cvi2mMGkA/KNIhoeQWHGbj9GOBg6
vdxOmYnQjtCFO3Zu8pzAfxMElUkWvPx+7AMHfjwW8Ri9Li7+YR51a2GmqxTw9EI5
fZrn+1W9OZMGd40K3vrEpjMZpxpNGOKHryi+/MC5AswjwaAsGpBbTyQZ/u1oAj7X
dmh0xBn5CPQSU2JZnP14C/X3A9FGBnWTCsjhi+s8IcFTfRzAjvMRk6nRXnoQvH6r
K0JMq7hSsq4JBr+ubFQH2iaABP1mtgj5dcD5u5/sHfKBdc6LYiNhhlzkFN5gqFiH
A0/Gd+VoPxB0ep7fVkxxr4/ahXvMuavPRYs0msrHj5CWWTOO0iMvvkuIFyw/PIXS
gpoWs8GfpIAHLmiIsU8fYg+qzn81OOf/UXHsnYZnwDn7LMJOo/Kppy6d2UNO3TCK
D0xpXyiDyR/Tkgn62cyRIBLJQXhuVKG5/zq38UV8hLZPsXVS1kUp2090hjMyky8e
3lHyPJPbMvWVZXe0vSThGECsRjYq0jp78nmH1NwQHfb0mKuVqiB5BOPG/JAstz+o
UDMt303p/oInZOylJVDxq4GswUie+AbZ95jdecv8BInDv2HN4yu9XnwHv6N7yIz+
jFCLzp4lsmyFdTylTLYQKeWZwcO1LrfSSRgGze7L2VNY8iZpYNQTpZSuCoVRrqYB
bYss3dCpJ8N4scuaSauzwIH7/KgxCD6AP2VRRbi+D78uqDRteexIyS2Q6qL0K3Z0
LGR2cD/Mw0BQgj/hkRSZzz5dAh1YA4H6RQYSj+wmopYqidXzkaOC9ByPcWUpmBiy
4fNLA0CL+NWHZq+lOYTRegsv9nRV+Q7tEsEj94VNekGPqxyqKaC3eVd/dsteZvhX
0Z0aMg0OuoBfx8H9zMyL8biFv2Yf5UTHYYNLbmoflNidcxJF71LZhKMrXjaeDo3f
VE/uixf5Lkpu3b5YgLZ5TcWmmtWmL3BgmxtULGr0VDfQltG2/ODvWisaMrN9kWT2
y2dz5YUoipZDiNIXjYEEIQNDTlt9JU97AgzyKrwGlZJAr960GKKiu27Q3MvWLhRi
whde3FT4V990JCCHmXP3Ekt4Ahz3+A758h1XFg8nbOrTrrW56enfDkD+9Go1lT4E
h6htUtITsXR3m8KwXVs89LvOBAYE6ExXKNX+TytK4litIL6m4YN72mpfzr4uBkbu
OfJSulaLOhDXFc0r4L683+r8EdIxEm7WLNUbM3PVMfai4Er1dLzTcgvwnbG7I5Hz
HyUIkcl88JZP4EJGTH3CjSBLoxgfLNz+8nIMSVgy5+0aouEITfkx6XHg6rSAQdNs
RWjk3wmI+J4wXv/6acOWK28aNPSVXGSyCTan6B+KQxNBUW2XeCYC2PuJu2SASiwN
xsj/imtIowlnVerxgaojq5HlLbYi2dm1ioPHmmIFBHq9ZyhtYZ6QOEniqWQ6DVeF
M/OMniv0wf2Weij3ZHjdNY2toIurrtgSFuniK2CoFQllL+KPMA6PCDf6gnzDyIpN
voGu5C/cb/zGh9jMmX76kURjx+qfTH1O81Q7etRN5fC9ZsCSidJWpuW9u6mEhR1U
QCqGIdDJMJoIBwj3XFziHhWVBdLYhWGRW44OBbjwQcfRMK2l8+eIQ9JB/KdlL0/z
Ts+TQz/OzkrW9uM9CxVzKKE51Jc49AXpFLgx5f9g//2sXvS4mVZGVCIzWezrQjsZ
e63ec7tX4ffueVDd/hI+spWk7s9mmcfzySxOvbwZmT1yqEnWKehWiMcbZAHd5WMz
fpUrczuG6VRNeWmmRRPkJuyziNfE7k76m9x+BCYW7wS+7EKt9F4iwBNpYaTirNbW
SBJ9HXoF4cKlscYKDZMa+psk3byRpFve9rAiqOakRmLZlrdC+an/1wTc5iXvKvjs
q+PyhOb8l5KU5lNGyJoBiawX3TzKjwQwwrmF23etyV0/N+9t5qwBiwqcbCiV9xWx
xcHjqbeZ/S/qONW6exlPzf7okLOTLzdRdL8wfo4NIaGaZL515WP6eKWL9rUWa0Vm
BikahbMIFWHVBiIvYhTtzH0RxewaCRREfimEM2yFUZ3/ky3tIPJiqixnXyEpZzlC
oQAyvxlgoxBbp0NVVg8pXrVieQ00gQtBPmi/UckB7rhner9ExB14s9Tns7Oa35Ek
rdC2x5G6N1zhXXbhPbyPC1sRwYRomEQ3qqp3mv6oNIePYIq/E4BaqD5hUoqxV1UW
yJCRVn+i9aqGpEMY/kaU2/YNkQ3NHYqh7TMDZtfqk17/7OMugiRSVmc822MnCm8H
PcwI8SbqMrP5j3M6LKuqL7CMLvM+qLCIm4JHsVH62HlCx3+453J5mnWUbCoQQ8PR
C0lwmdFFQX65lKxEiC+iBOcuWdL5MpfkDD0oYfcQYwSkn20STvRJF9/d/OBpzi+u
bZDXtHpfxOFORAT9n7sfRboZIrtsvQ3kD6iwV4Mqt2uI1CknpTppwRiVoeTjIrfE
AZLaGd6835mmW0oA2dA6aoBUJQVA0BDuvHnLTXwnMNM1q+QeK0P2QGfS+l/LRUXX
HmxYjrvkMqiRodspXprmbJFHiXPcZlQMvGv+yetv/IhoAt3oZGrxRSV4lLU2mGE7
PXRT7EQmc2nGMxtChhgsknGdGHg+8V6PEACeOC+2q64xkBL7Wilf4Oj857HY8WjK
AESIpyeA2cG8jrEIA3DRtjY2W7xnclLJVqpHbv9aYw7/5ARyJtJaG/1B7cHDTOQS
WNKD/nI6j/6rv8dBMiEUrEqNggIMQLu+YsK26aFO2zbYOd0BCgi3CZUetA22l0V+
vpBl0ST7V8yDlEr2kpeyOXGxrJ1ROfhD2Z5NnzxLbDxp+nCisDGe5mBl+vgnkxXQ
eSQlcG3Vy2FxoXA/LEoG0cdbYzauKp7UPvWVfDVPTecQqr8k2FOC88GIxNtB1zfp
rPExM3RAU+L1thXaP69LiM6FAcd5B4So767rr6k89y4W2FpLhU8dCVXLzMDv0Vsc
DmaSu9+KFAXj4ea7h1xBKNh5tYCKYlHXea/r8Ducvn1848qJTCCAGRdKCzE9wSBi
PE5i4j2RTKdQ4Kr2GK6pgKTNCJ0eWe4xy5RVrPFsAkphpyhs7/ttVXdax4m9PO7P
MeHStwohv3p8gbKPED7AiDbCgGN933MogMbqHpF6fqudpz7j8bNEpbtJ3oUudEsR
sBokbaPIizW//+adDPpjEQWAzS1FkbwHLQk1TqnND21YBg+PFOKhnfg7jW1xVbVo
DtorfHEQ4HCBMaSwlKL7/JMOxNt2kkcYiVStE4/aLlA+wqYUma04GLG5K1/JvRKj
0bPlp9V6gdqiyaHVGr5WHvqQTiS7ELSbSyhq/PKMn7OUfIz8it7KJvFitf7eYwub
wL2Bq6JA7v/YEPpvwYO0HU/RgGl/IFDLtz9GlL5kbpoSaTFSCPoAUFnDTn4xJFRN
RD4IRLwtaQ5w1ZLBI6sZOi/iUrMcHufWvD4OHcL4QAbF0caNSGHaQosEnV+NyK/K
yARDe0/ub4RdGpd3B+1UXrPRbnMzwBGEQV/HfSe2U/InBnc9DFhc2+C/YHw4uu4x
qlSBdy5e9VXZi3v3YdnWYMjezFJe0QaDrXdLbob13zXyZCVRSfLuAlsnTui1raCa
3DBvQp/EA/oC2rOnscucvkqq/X/pSnq6TKafMGdavZ7FO0425XAm16zTyUplNsMR
1x4WNS3jPOJq81oTmoTLhvU+fANESo8GkTNmMKcN2sbaSfTh9ATiSSnfYlG7lUFa
8Qurdr3LSDRfXmN9VBY8gC/g1bwW8bBz5MI5RgIRQ7VdU8PQZWwHndB2Suii/qD/
JK9nu4jIBG1VZLlwOtRiSizZW8I4hT6lOw2dCHa992uaZDPmE/lPdXoCgkezXSpb
AIeG8EKe2FBxwzl0u2BIcA8tOtVj4ILKCCiqb11PAzABkALwkiv0cihqQzBOTLqi
oIp9NEeq6YHr4NJ1nHjM/7EeqAfIeMej1ZDewwg4b/i3zwaVoyiT6U7E9ahev10C
UHw6eO24cLWsla9PhCy+uvnqXDe6HJgsLb4fxlaiLsLk0tMVsxvX2RZFKGt40NNF
doAtOPraZSbwyFOXrBxG6amX3Eg0OWDA1x3H6Kzx/h7XC68dCTtJ+BFOSInUEx1n
DsJ1XylKhNyfuspnlmkb2s/G1sXIGdU3kJgyR2g/56TYMujcrSjTlOGfqyfSXb0h
ATeiULp8DROhUsnK8uSXoDS19ADqaDa/ndF+vWkwaLsfvn+JoK4mPdwMN+mfMu1n
D+o/uTlnlxgy/9K+Wf6pQj0CBANlFelER/HT4C4u+JIR2rJjPJJpVkJS2/IvFv4T
poJuFJni5wcIDn76SBSBbSLo1tajx4e6GMLBmDdzGFU29OxBMKkPNeDr1AbMX9Nl
F13/8b443CDE3uSujhgcxSQyxdRmTxWX10jhIQYYqI9BWpMVewb+6i2qLPKyoRK0
NHY54jh3HpDumY8IVTl9EUaKa75lpizYfUqXKu7kV7A+gJz7ZvO/dS+JDGM1n1bk
vLdxyqBc6qbKT4nBlaXkkR3RpS4dCaUxLysnvbUAnQrADu2aQIAxMDh+7U265Gzy
gK0nI+v7HOw1myEn260XdYepjAemDywQHJjUOBCxDVoKsnRleZMLyGAzCc6TtlBo
b2hMHtahVHZ+a6ioxRrfkwyML1Y3tkHl4tCgry1EdUO/Bm40SaCH0ay4+/nPq5HC
/ZobN/9bwyRj8/Tfy7ZmOmxW4s21A2giO/0pjPLSE3nWtz4Is6ufsW5DeNNbfCsv
CljEi5NDUorQWxqEFoV7/cjzM7ssMtguyBnmEivyEeu6TeNuZfcX6w54k2iD3tZg
4KjTgG3/iP19F0wP/nBmSpSGPDIPQHygmHwjn3uwEtM9zsdzYnFT72R2qscWOxsl
UyJlsIM/RQmB8WdY3NvGECh3ajmmPweF4zWljCdkudxhIMpz4f7BCWq8JqwOyCXG
q9GlT0QxfPbaW7Ny1X8uMnl3mGirezc846zLUgt4btwx1VVlpG7/yLT6yfS0+pBP
C5XyEKrTu7pCLiCfSgaIeufc4nwKjvCBACkvTeCGbwnNvMwKZyGaXV+7Ivn2dnGv
N5vR1xkWQo6uqdZP4eOffpusTzmMA6uZWMGWktmRp8hJ3b34RSFkxE16o1VabU7k
igTwv4PmGOflmX6PI2bgeCDERi9d2aE5YxLhA9R3OZz9ab6QnldH0pzeYDGpUz52
WqBsr1XXoK8jFhVSph8MqDGpVMO+EEDTziQXfnG2HIVelFuCyWAEU6BPe1TYIXWZ
mh3xwfzp8mMdXcWDiYXFEm+kfbaAi1Yk17Z2RL1J0/yJY5kieMr6zAPIff1sFtJV
kvcYQ5Lfu+3kXh+RPjtiT/1EZgqOUpx1TTNS5ehnCccCd3KiTKll3CQvNhG5xif7
f3oMFpqyQ10LrcgHfnh/AYNPxpFISfFN9IDE2U89NmLKYpq/VWj5+Vi92YFQGt5e
5ka43zJ21JJp+1NiEsOfBMhDOWx+7NRsQ4csvYBms0jPtrfdlEZ1m/QrokHwCUIc
CB22VexiAfSSk7HdmoIkTUAQPUO/RUXJpV35866q8Z/KuucrsidnunvddyJlnIaZ
9zK+tsB2ELR+3aSGZ35lPHoNX8yJ0TfSORTApWeT5FraCG2aSLXPBVkwOuk+7HK9
DtrcbCpcecbthAr4zj5dYJoSxJ9GEcaT27agBBXBWgJHsVALw6rd9SCNnJ27zx3R
OdM4UTrmMA8qIEpWWNc+VUAt5GkCJW3NIEx3s2o9OGcy3meKdf2y73k+A6TR+y7v
ht9HWqH36O0CoZEjEJr/KYCZzH0iyW3tasKJFSf246mZpzrOdP1PSN4Pvrrf7XE4
4GyGFdqgumM5W4qdIHHB7PT9bdelNLwQZnQddokUGXSBx141NHRG+WFpoBArpJ+x
ezpmYqRlLMhqwbd5NWSJXjCxucCGZNbQlZuwlEV7Y/QC2NQt1qk6gA0+U+WN06mK
HkSh9bjnEJLjzhFkpCltI/Ll8BG31m+DGLnXVIltuZWusopXowCv6glBE176wX1k
jbuZGVFcg8uC5NdgcgHO9RMNeZsCN8yBoN4bQfdIVddxeJi6SS9ctab45PYGX9IG
ewnL0vljFf+i7IbvhLkqQ+zDpQW+T7em323QsbNoLe12l13DGb4hd+kK7xF6whNF
zH1W9fOX51EfH+trg58mewwn5F4wsEA4oCeLwo7iTN0o8BCW+VTazzYDUIy0B6fo
gt8JZrAyu3iIqg9VoiCIOK/mNuqaNKcVlqOc4kq7BJYGGhcIuKQ0Rl/2CA5fW8Bs
s+FJy9BpIUP+DfL3n5C2FYKgeqdY39toG1iqV3+L8oOJ0Ps3pb1evujTT9eSG/VW
0DTHvYcPwcOmAn3y25ZdBsTM38Y0owi/38PMJ5YRoiWtjFFPDzcgFQRMlRTHH86B
vRxC/6qeN7lNKpDA0lbxDgShANG3lN3BjzANez2/8rhqq/QH5qmjgQ4XNiWGcMyQ
RNarZ10ZouupJqxrv6Qj35H1gMiHHqWSM5s1uGPXpzbbOyhcgcE6MecjNIJPCm02
91Jpy5GvnyukiSCCSrxu0Vx/WerrOEQ9a01hJKO9Na9c1ykaufNy23nU/wiRTHWZ
vndavYAMF0K4M6FL3u8vSYMio/ejqdM9g3oKlYmJeSGw6A5bVjn6I/8AA9j6SVqk
a0bf69etJ9ViagxVxQTYdalqRy+4CJ8oOJAdCsPLRejDdwfgI0q6nl3tI1PKSj3I
8YeDcMON4rSAHU/hQDlf4vA+0n0Dy3iRkB03shlCqEzpL2b70QJUpjPa2fazzcMi
JCtG/kP3mHzWd6ITUHusQkexgjqsCWUD7yVrchwy80m1PtQgmR07rlwmszjx2xR4
H1+CkgMxgHJuBG/BXs+Mmbntoksoy9qKxkjz6oV+AGJvmoco950OPqo3+q2jjqDR
fj88cpJp8opKL+sOlO2cbOBH7jt1Qrf9YOWK5h89Jw8kZtydh1z5BzQgfB6o8EXC
gBsJF/SUsDIRufp0wtvcI2gArl592wg9lGD5UanQRNioGPp+hlXEH4Ks17t9UzHD
fM3uchBBuZqvZ32jXUsctXGycQRGBRkRqnrQYdBQliEN4ZK+RftFa4F6GgKsDdeF
9Ihd3rwMEyDSK3UG+UmfxZ3B044mz15EZQpidw+cGO2Ms9tfp0NvW9LGgASo1lZO
6Fcfg6SDm+FlL5pZnVEDkGVz8CdIa450493m10wLwJ72emFUnYQ/YQmtbaxVhRdA
OWhEeGnSSCpjPhn7TcVTeqD/RX9tbU/vyrAS1+aAirADEr25iH/GVJ0RiuPvxDi5
8Ymkv36JT4OlAKgJsHPxZS6I3tUMFw4cAxtf902Fes9tznt/q1Z9T5begOmaCAPZ
iXMEUMwHhEVSZpam3rYUdnd6s/8NGRT3F5WOc/j1HqNei45oiz8ohdFu3UQoVyEV
P3okmcDNs2W0gOAgq4qQdYX13coJLA0Q6d64cjfI+bjejOCPeK4R7SU9D55/JBoR
o2EaBrh4G7YPheU+EyhSWUivtc11zkhGz68Dr/hGmkpVW9hgfXL47120t3cIgIRa
OjFDJrIv2SLM3dcrxqZL62rVQa1vqQgI/W1vTYUAlmAAlJhS2LobnFwYZCwt0ONn
1n8BystER+kNa3ms3DLnWvy1i3zdtI5tvsEyb1eizCVP/9fTJTaMQCRW6DXIM2Jd
hBhpQgYqJcJ3pTw0n+ew4Nyrpp9B/IJF+ctO5z0p1KynlFCCy9/u+Oab2e4oK8SQ
RUBMOYOdK3Lk+8rzQtQLEmyQAW553f0s5Kzatx6bDayyfATkUa4+Ik6pWx34trfZ
IPB2ZJ6uJZ/38i674xzvJxtJR5xv3nNsvyWahb6delM00jftp6IzbA7KPHaiStwo
6e/XDBKyDf1st43gFVvzKo1pZjlJT8MaM0KjFc8nxfKXK8mOoReiPV65MppHY2tH
mUSSCbeosHQU2HwUxJYwqk/P4gYhK/FKbz1563GXj85nvW/jXX6bZ4NVSi2s5/FY
s/bH+Qfcj/G+dlutMSEUY7P7Ew0dmy9nNrfJModwGkj2B+i/uDRSmAxzU1MDDL7Y
392yZrR/hfmiaYO2nHoZa3/dK/9KS6wWhyO5YG7GammYivNk4Ws8vpfeK2Kc3zzW
/jX44kjA2hXh8lo6ApiE+tnZkoFov7t1/bY3LntPux6oQ1xXWA8wKgy08C2bp7ZG
4KjMTW2AMip8gsolQSyINUBradbLkVTyrSueXktmmmBbAY4p5ghXeyZJqpBoWNoQ
nXvD0RbZFcOpF/TC7yA/pw4/1mhWCUeb+iTX+Yv76NxmRswlJjoGEzFzeE8Opj7R
7tn7OqgSBrUWfZAg8N7f/dMufStFB4cuH1rz2/FJsTKkAdvwneLgnrPkbYLkGkV+
dSR1KcZQLwNYCeaOccaBnAVPJlW19O1N6FiW8PvLWW0dqg0Zs8H4PBPC1h1U7FpS
h1gFmTJeoDa/7fXnMtM/Risgpw5kdHSsUhSYnaeJ9PFOsTY531FRmBT+QvR30XHg
2YMGrCXBXkdOegQ1lo0kLPCUvmhnwXjXP7ActCljNy9NvISLQeQwzkoCf7veDwOe
KKe4Sy0enMBK0uV1g3DeBFhBRBvnfxbHtGM7woNuhE2OJ7VWEaflrMxMxfF3S3JT
fBioRBwhJVtzeY4PLqdMZ+VlKg8lDnDqTCGUyfP9+A11OQX6AyemqhcUThTX7Asy
IEc+FuBBT8kW3/y1U0aj4mhP825gDRZGlIU/iXj+Gwe/oOSkeTe9PWPFljx6o4Qm
y7ilOi12+k+ewWbL4L1UwvvTrg9s3pwwbUmE6t8VfMvQIYvbbv+HK3Lk2QimDobj
ykKoAUffjiXj7kBsccCO2rvYZVy7bJK4Thb1/QRedRFuSYaMJb7ohRvm/Ib5bZ+r
tQ3+/BQRNPPRzUA2Dm90it2AwsplPDio/MItr2aABIxf6Jsb3HjSjtVSKma0W3Gu
u9ctqZWfhB+RbiyDlfnDBFbwRf/l6d4tHUsYO9Dvi8qnmdiTlX2H1JMt/RBzdtt8
LuQmEXpYVnM5i3ckjNqfthAm9fWBHNLXYGe3O6GdoLk4IAzeMueQx3hZuJIpIfoX
TKZPRcSJAuTzIhrb7VBxpgj/1KL2CorO0UgWTRF+KOgv6+V1VPJQQxXb1wZU49tV
2GYgKGLAKw5BXVbgy7EPlDTT9cSjfi6Lu94tU21YDbMqwI2c8UBGf6AO6NLnQ9/b
1mhPSL6DgUcQ/SHo3R2M/PKhqjDgJ/5s+cARV9mJI0v8yV4Vft+vcitl5B85S5mM
pYDL3183UdeYT26NKgmDRfXgRsGvBw6x2GV9u9EUstoJStT/gwVuFqw/IYgA5i3m
RXho7X2/mQrXYgO2WmLsMBoh9MqHxz3CT41X54P/GKYuA/6bz8vmA60UuGeYvmcf
ETp7isMMb01Pk0Owkgw+kVscJwQwhFMeKocK3rBvmP7SD/7Vzq2pHqDjEOew3pcC
7vRHwQQDnwSdC6EFbhtlxcH5X10Q71TuW91qGCOrass/VAVILcih3Ur0rpXeENRy
SHLjfBBDMUtVB4H80hQJlWiZOx1D3m5DG3UbSx8YGeggDgHYpwoQsn7oHrxE4NEg
2RsxiADZ5b60SVazCFgIADcOwEMtshS3LYSU9X4e+1WG7Rl+BC1hFGffzUfAl9sE
i4y/mr7En8jLqgAJ778BFifEcyLmEBFqX8XIyaWJM0whokf5x6SkzWYzsGVLOC/A
svxeRDauTczvJw4OZ0wBxmEWm43GSL3yqO+sHAokg7D9KX46gzUHTEJ+B0OnlX5L
02T17nxyVzxQdbpxTyWKCtIrEO9jEBcHuLqGtouPeqA9RVgPXt5ftcSOi3SdU7m1
CgB5bHnFvK+Nw2z7pXX66xRlqZlDbJkxRLs3fmPbiA1wWEdHbggBGSN7FQuFZCO2
YYJ0KWOGMGMDNWt7H/EbQeFA8MJ7e+Z1eycrHIVMNCyAun1cDquplIlRwSYd984j
LgpU53vdZBsnLQv212EYz0g3IYVn45kU9vSfaCiOj9SlJRi0QC1KzGd+XYKYh7IU
6qYmlmaHL3En9diEA5wxHoa1vbF09Sy3Ud0opp3bC/D2lmsrFs6Bwd72JcwW+5x9
ilkOGErLSpe/kyhXyWUy33neAYR+yjkUPz+7dGvEEDVYoWmnxN7ZVyZox4T7goAj
tHL+nMfnvdQH7EHvqBBDK6iqzECrCV6hxhagoSFjtV58/zaTl6WDxSyhOZrYQakb
HkB67vVtneo6srjVHzZ17t2t8BcHO1VQ+/9xsAzONHwNYJOlYN2bsJiPgBH3nsQr
4sTdr2B3bRxQQQeyaMa9oFH8V2LXM0HDmB+EqZF2fqevS/iyUBGTxp1JbcVwfQJi
UOQTzhwEf/bp/Nt2VmNq7v1lmRlr5B5SO7UyBcxIRc9C+OAUgE4sKx0xIFtbUasI
wVs4tKMrR+zSXZFEr7kdff/+Wi1xgV9cBvfpFgqQUWUAHTMZUikh9Ca4SYzTLLte
CYsvWGCOm1KHvIT1Ta/F5ZSKzMkUpRUjQ21Qf0dTqyUTMaHqJ5dsd6SIDqWTEvkT
mmNFtx1da2Xf04uR1QI9BcLW2q71vl5d6iX3xzCfCbsIvkyBsGFBEkR0xrj8IZQV
t4Kej04fNCMW5DfJZMCbCJpEHxcNDDY7JkL9PL/Kbcik7kGNofs8qhbbNtdadoZz
0NT+ch19db1le3J4eAENbd+R/hwOA3uG+6GCxg3xkkojaGzEIbUMlZaLtc7eoyOI
21uTHEWMUhaI/7C5ngafaNGds10EPej26Vz1sOKTetun7HIWJeZ/TZWwLKuiRGBj
RmOsmI745OjmUfchm1nBHvW0mZ71geKcoOpdyh+ooO/IpHJsuDBoI3fiwRYzmJng
OoR2bVoRPDM8CcHEcGVGxPX4lUOAs0l2ASU9HsKHE4UCs3blt32RZ7ixf58eemVd
jo3a2twz4kZTyCJW6UwexdEc5uoxlgsEECS0smg2VDdeEyA5Y1UA+3I8HIi8ntc3
aU+ZVPbeI6D02Ro/7vtY6lpVywJHH7F8PiLPnG6TxJ+LB00tmuzm1LQWxieX7Ma5
KyHD0wbj3tZ2/tqG0bWVy+frLrhJcKecaZlezNknpxNZRVFKXIsuyvE1m/RqFXJ7
TT+1hHl5Qm2SYEck8oDEwdhJJFqNFmuN04LOEh2mqYj49+lkKtfR77NjjAPDcH6N
Tqzo+znbyVePh0PuSV/DJ6a7S4pOsKiNVxhmAIrX7IeuWor/eQckkv2hvy1moHdZ
KV+kyGux7kfeDEW1bvCV4C4HXVgq5rz0sQo3hkWm7s9HR+rCbeGlGd8wDxymymI6
3GSbPA9RgG9SVAO5Y6v+qqtb5uVSpseQ7dVX0IRcOlC8Lo+r8rg+ZyUgSqosRQjg
VIJeymgKPeOCjDzj/bDmWV7GiS4R45Dhn0ZQP4hmE1v3VzzVqDXIi0l+4gFsKkQE
7LxFjYHGvE/w4rRVoY/34cg2Eey4oH+L7F1eINvmpQN5Sjw3k/N3Y8RAKzjHXVSU
VbQ4lYqH9ZiqGNSY9JUQQsbG0wjyLhpPbaE63IAA40TNu/5EAHnKoqgJ+66mFOtu
eoZBlEvacL+GdfHfW1ZvWeLahnKkXFCYeDkayXtpCcQ5FuHEcWu5SNLIttAqfbSp
dFzbu+A+WSJEJgK4F4Bgf90bMSuv96VFKva8G4zUJ010oAHWAcnEACpkD7GAT1jG
TjzG7VQkwvLBwgSZyV1vmfUFATDHRM0cd90EfDA96RGho1FyKM9Q6qURjEVchTdv
VORaFlApRavyQIo5nkaaKnQBmNYVwDTRsPYhv2PuyjbLzgabiHx5pYyO0Nc/fF4R
r2S4f9f2oZgLjeQawSGutoZ7nLrPA3CP3rziEG3oyOaVxDSOf504fZugmkKAu5f2
6K/hDRpbCmBIP9Xhsoh8ryJXxYKjx4p4LLt2UC5H2m5wmAf644Ip0RsuUkWkLCM4
j2PaaTcFWILQUC/1du02S6gb9CzTbBlxjJfxAjuxF+tqKHMzYtrgiuZ+5oKjKQKG
YSlW6b+1EEVHE/6Df7nv1X9zRrZmV+hDNcUUJkzQOH7jHZaHv73aNxneUiFEv/uV
WJqK+EyLfI0koUZYi/o4JH7XpHpAd/D8eHmR/cP86avZG8+ED1rCAm81yDbTKCL2
77y4hNm8DCkp5JrsBtXaky2m4u+dyu2k3pN29K+gSMiA7hxgoXf0nElSIuigvX1p
TZqX3XC6kN3Hi6v0GEH9Ok37B6382FXxeqFGaiQugwXgnVRyLQY3lZqeGJx7Rd2c
TBT6GHw3GB6dP4JHXpMB1FNdKry/oDWw7dL/tzazU//uDb1YWSHla3c8xp7MTTzW
imxUdDTvxjLB8masImqkRx4u06Nost0V6rM7kHwgwItYq3yhOmot5iL7aU7VTbka
ZlYyVrjjBRRm53xeNRN6mpqy553XwA3ySF/Qf5V9JMtIG/5VxGPZY5K+3jH98PGk
W8aYavb99kgEdDQAGrHY4yXyBb9JVGJPILFCAGWVr6zju57j2jReuxr8z7IBajgn
bAgFUfD46XDmdYzAgAtSAlI+aX/KTarVWlNT0LCpvbCUnO1ju/TO+rZPBLFDWulY
G/Uh1WrHjluugEER736tRUpHt72Jwu9HjyuJwFu3QmGcjjnkBmd07qJSDdx3PBGg
H/Qia4+aAEN8vEzFw4jzj+7PifZ5ue5wXt6hFko5HxSFJwzt9GHGBagCQu1ptb0R
KojkyfE8I1n5QMpuL5rW36oo2QZtOdyHLnIrSt/mAIx3zUzijUSWW1cm/zte0D1T
XmsY/zFtoDUmSLQAVU94Xa2JIAzaLO/Espgox6sTCLRj70TxLwOvbnd1VGDckgoa
iJoUHN4VliSfvYaI6NVl6qH8HXdyuBjq8rFLfSjOxNNvo4wrW10pmpHmuU+nJ9QM
8O559IHahldRMi8dRsCSpgi0LFr7jaCdrfzprlZgVrw4kZ7BnNWZklaTrk/xjdyR
aNs7yTn13mlCYN3hr6N9vCel7ceIJZpwEDt33XcI59Q11bGi5rE9Qu2m2Tc/gQ/M
9YdwJ4hzzLRO6+EPwr6hTmvgNhea5wmfJ3S1PuNPAfx4j3biVviTbQRyNOcR+z+D
mjpwbXBQz3WKQyF82VnvBtwAblnMw+YDa6kst0ExMSOPw3JjMKv/s1ZW/IWqCfLw
Y1ouMz2Zst6B25JHDjq0RcNsrPub8MYyTdNiXOwBKELH0u1X3ew/TQmVNkzsvJRy
HumZujoiYEQEMeukEPnwbLfx3s+zKDYFdhkMeqQP7D9mcWvpWzcaZJWdXiAOgnwL
CFQ2dntBxVTjTm5S5lfH2dQHErRG3UjHaj0jvue4t4J1TLWKszq5CE1oGDr6ITF6
MPpGS9F1g9WJZcd+dP+wv2X7y/pejyaY6d8r8dBUTX6+6VGg6qJO6KFYy5fbHVBw
lIlssB+KnMe2d1Mp68Qp/iQEaAHwo35GCHGvoiGEt29bAYxreRvjx4kx/5y23YbB
GC5khX8hXLGmXdEdK7VlJvtbk85Ve6WMS52oUM9C73/1Z3Kegiads2Xa4m6FOAVc
4EjHVM6a/OwIUWfwXN1MHeC685A0u7UA9xIY9omyTNIUvoFvOjEcUlGoWhAjziH1
KxvfiKJ57yMOY92uLZs5Af2t/OxNBKmUmsxSRhwwTFDDuDmQ+dpCfkDwlJbcJ128
0jkrqvgk7XSO8VNcElUNTc5kIxzK1oWqdOMU9Z7P1+GhaInDER+7e4ht54hEcFnz
BcgJa/AkMCGoDHWowbkrebpLkW/1oa1nrq+KdtbtGy3BU41/yOPgMIjtiJlh36bI
ZtCwSysD+1RRUDd3M8iHw810wThU/nToBHPeHIyQ/FWiaXof0VghbohbIhPgeuUN
zzizV1kdiZQfNE7ySTTDQZj7HR1uVG91s7Ys4ZMJISdBY40cD3qcbD3Ybb5sEUCK
9r4EcGJ3x+bJPnupJk6o1o2+kjhpGUDbw5oF8zue8VUugf+EEA7VeFxFXMiAzUhq
s8PYiaic4fTVLg08jrMqzLE073M3bqyWjgfIpyMdHPSUw3tW0io9itYMbLbk5Iv3
QfoYYnPeJtl1856s+K64DcN7xL40cMHnC2UkOvKTuynvQRXkfm/y+Jfl3fxPdOIK
6tCxR5u0zQWsg1SLLpd18AimLQ/jwe5EoaRgF9oO4UPFh1ef5xBHE610aDnGwNfK
Jh8b+7e8vYeoz9KDapIPRYa15MD3was/w4zZncWRb2HAEmHjK2lEP19UhVdTp+Dc
YB4zR2f0qPTiDUgetXEHmPAg7bHS6yBBQ98n+b9LQQoQ5CTQsXrtRUXplVoDpK5d
kyUpTKcn7Rqvre6N8OqpdMKaF+vTkEwTc4XDme71qCqjS1IaLMEn8OmOJH3Isd2m
NrEVdE4ugBPg/I6YdVgA8hvLAv5sVZ6cbNjWnqrbEZnhC5gkzZRnnO8YfqWSVO8G
pnF27M1zdGyoF1sk5vHHrrKG8MSlLNNtuG86KwTe8O9kLoMyWOzK+4wbq3e4zIUc
REPtJuKT61W8Vwv0dh3NBk2T15vRjsZrWYXnj/QzAJtxmGf1lL1zR9yUHaJWfoNr
6R/+eASzMNNDv8nOvD4izhdGDyn8FiohjtZnkw41vq15zmMoUs4WjC+nFjdemiOb
GJ4XKJ9JTZfFYdEozVxKlofrJJTcTtMnuBtC3Wfr9XGyE59BaRzyU3anWz8qqV6T
GLd4BL2cyBE1PMOvbjWvR5I7PGJO5rT+SwR/MlOPd474p20FSjOAL+IHSkvqM71v
B0L6wZJ6cFyn/S4CYCh2HGHh0Zo2hHSxDNeN50LVZqaA4fPUg+CTigWqLuOLYnpc
TqTggvbFAsLZTCbGS9PeWug93jpAz5uk/I7nAVEq0CB5m9o+JmxPtaDXtpVhRWez
hpiOFpAUNKGBtKdF2NmkvJGqdbVdg+53F0BDNfBdphSgEP++gcEdrLJY2Jc+DSnl
5Yvl0LDIM1f2FTMYnafBXu5ouglTwvNJmt/sVZ7CDPzfeNhIAivvb9yjiCBZTNTD
IoG4vsPjg49ZMmfDf+GJNlPQ22eXRBOtIROWNWOXkjhpsnxqRS9vVRBKaZv+DEU0
mPWJANZh1RuC0e3OeeYslFoQhl9gVzlMxf/0vd4BLXZLcQ0mPScO0+1HXkJCjCne
NSbTNOkf7qkM91tXFhoobZbq+O7m5RCAjLrUNTQ5BSIH6XvhvCM1ZX6uX29fiDfO
119bAR9hVSiB6hvBozbYR8vStwPMX/T5GnwyFydWR4McWb6zHGmLUWTWkUaHLITH
LWqPMNuiBoBgWXfE2cMPnvrCFu1WmCRJz1DtkU8ATdSJxUZovfDq/3fROY73pQm3
KUnZ0BP6ucRwkObDqM1+ptrEyLDPVZGtgGn7DgmnpITYNq/u4GxDJd7USp0mVtge
v36gdir5zySs+JfM0lfzkOI+bEnU2NsMPfjDOhZ4ZnEd2mEmH50tvbMDy5wKXPM7
uhD2D3uBmSoyG6GnzXv8VwehmZasQ6ghP8ZkrVi4wwByG5uQP3KCE5iAVNuyQPU2
DIQhPV/NrVgIYX6UUHCdDM6nI+3GbGt0SSMoi6SjE0rxJveced946DznY29v7zYL
pF8dpOb26+J9CUqnSqDpXFOrJJpfD2PNZgPusfbUkoyvEIgonNiZt3bwTYuv8P5+
9nACTfE1UjW7nFIZa/TbGLP67lMU7wpecdM+r7Y4neG2L4pr+BVR8FxsmxxtkKG/
9s1ciAcjaDyQM9X2y1K1mfOm5zCrd3D9cVHfCKYEkp5RVal02+tQreLqkhAw83tT
yMyX39BHklGrM0N7S6dbGzm6ucy5jeGL8aONW2ZcIuZmrKF718YFZ5VpMQtO/uhF
6EzGIxXX3ajJsNsgN1Sr5kMDutKGHzxvxKId/qKlHq9s7BKpVbaCMDULv/sRBz2V
/kSr4Np0Yry+mujn+OkjFZeil69hlTfvpT1wEnAKQ0rQ6agko9ibIRcrx3HuzwNP
aWcdgK2QLYyMtsBtCQmLXZS6+4r2afkoBlD7FaF4qa/FMl5hUwCIUa8OF+GJkt9J
XNQGVqi2NlMPoaz+ZVEaAxqMD5hs8lfvtiH8uv3Xt4/ej2NlA/TcdvW5oRQ3BJ4l
4iFtiql9ujxDeF+/SNs8xe1coAF5yHEyP12/xonfEEZqT7QqGAx/WgU5m9Al0uLT
+vWp40HY2JxilSeC/NpUfzbzMO3TzYxqa4TSDh2Spsc6j/1X7l1w/0JesQQLoxrv
/2Z8e5fhpnnPGaqEhDztiElViLocabcAL0v/AYlKEViWSQLLgvIIpC6qLtspNV2R
nfCLxxejp0cVQBVpkOgDnYkTaL0pGNzEaGHyU4UdsUiESrZL/ti7r9axFaCtG0FS
r4drrXzfHPHO7uezB9OOlbs8jdo+9+7NseCv5wvcRPjU7hBf2/Y7xat2HT5SpJ48
5KqCbo5Nd9IEo+hXEY0yKgQ3k0FvQ7fGNM7wFMyzt3AlWG7bdbDDP+xBAJ0k9s4Y
XBBW0JcWdJJL8sp8R5fd2n/1FJOJMWSvdQ0l7zSDCO2uIY2b3oanwUIGh1BJ77Ay
crk+1+EzFXrwztTsmsm7gpVKm+DpJSIOdfozMLoBBCClz78E1cSxny6nzqDYTUWy
xfiwxPGwOW6I8hLN6Bgf297N7yN1BL+a0BuT/ahfgHnyvxg2D6t1b/UOTWq96pJE
5HwSsRet2BvudxdEiFIpAHcr/EVUK8P3RTYB6v1FhKkn+HyqbzXBH8QQvZ94QMRe
tmrKjShbeWJhpbmzFRNxuZHwaNVIjhx9eDyEfKxxSevLsIGyNyjynB4ZrcmL33Sw
vhAeRdrPvXua19+eBfD99c0aQdZgXsz1LdViFIDG8y88kLaTOygRljUaVsQUpZIe
UdvG7mGsR+UI0I0CzdIvGwfFWLxyvJDM2Ke1PSkSP1fcT/hh/Hk00qBVdBWlGSYs
ByFa5HIEQfRK4E5Bka8WrLErKI+LehVUxzB5mRSTl6a5hGDwf2VxmTOrcBdHQVY5
2NvclunM2g1myyjqBCB+1oF2vSCWGFAd459mlEJNzTu4NmLsPEXx/nmvEKVEuV91
uIIAB+x/vfTJRtwRnNisxL/LFWWyoGgrBFGE4ZfIPgWm07m2GEQqRVAkCdAGi/B4
+F0VCU1TO4/X4jwHBVXjpXFo2SwaoCpzLeqreYHn/V1rFSJ1/E/L+yHSV+x5FuHC
22Qsg/Dk4pdCBqnxB7ZLh32Ukd9FrQIu0rhdQ46vHCn6lpDZnrLEeQmF9OnB5r8t
xR9rgjCxs4+nwL1stJfv2MPVlP4dqnz1nX4xQ+tczagYJozS7RYDqDQte1frlaAQ
3DmQhy3vRNmoXHEnQWxwfFqrEU+ZLfadip5rlEg4ZCohlIx1+JB1ShDiOhilmUCp
DSY22LhXfZa5WJd1Ihc3/0ZtVrneDRKcTnQqVD6S0NBBHRcXVjAHS/3cMSTYzEOi
BIlOTaJ8cS/ru+LA09UebMcdcc7mpPWn9eIqsF03BBu/p8qMdzRtvWRGpoP7ZUf+
SKkZiB61tr/hChtdkurWke22vy8noGTQ4yssfr2RynP99Wb4mtEdLafhj7I2bl1f
xk/tdxna4Je6Y828PkenT9dWcGYyYLaAcOHTnPiy+7xd7tO489HkrhHNF/NMsCx+
jg1VLoat3IZv578Noc90B6WsqLIyPVR/cIyObf00+wAwA57RE6h1pqSofCguLG3h
gcFKQDAaYYRn6jlB8JBs3t01hM9sJQhFcI5rDWRHR/+clYdU2U18vvbeiK14Bi11
7QCFqzzLKPzxpOf1MHVe3GqMom8o1kB0cGuqWpN7SUaMAW5rwRvJI6SmvxNdOJTU
0o/HBd8/nQmXcve45bNJkeehCcCZgoNdGEXgKP7STanX3FUx7Yo1AZp0uB026RD4
6ZLJBbHDCv3frpuk0Hekq3VXkEcFiN0piyZS8NXa0AWwfw7eDtLOVgBDFLnSumyq
oDGPpENTaYTuTZc8wcS9gN7WuT1rzXdVmQrqeYw61I19baltp/wZem8/K+FCx8SU
ldPZHfyU9wpxaf2lHFQt4yiedtq/Gd8Ob6dCRWF//uWh+chpVmCgJdFL1f/VycKR
mj0tEeQrx52SP56W3gtEFa5v4LuKsAy9dK8akehuMGq9HjNR2y5/G5QURvy3eAyJ
cCBVKRO1I4ZgPGsjpDYF1pQSQ1uYZ+B6+spHzUtzL37yOG3XgM+Gf2D8wXrfp/Yq
mLu+CtKzjCpLM1AGEZHplkCS5qQi2CHdoHJb0LleGMnD9ZqB6Axf5AcH5cq6eE83
KLvpSNczDwtFAOtQq5ZMpxUuVNus9QbsPXoof+G1GLZOAAKhi8begmKzoiMl6r5X
p08VkRQMJf4ZrqCZHolvGGgvKRF9sqCzqyxjFgmKkJgemIuLfLip7RBsrECcNQD9
FuW3UXVP4BLQDvaPOprjQSS/lFYsLTaiKpJ6HK9ohlz1766HsW02Y3xS1U2T3J9W
G0K8Q/RAPmTmItGyuHkBm3mSaYqT8sdcNbuEJUXITf3eJ8iPKFksvkFpXZ9iDnIa
4Jepuitobtt3LRhK8YrBJc/NpfPanR5sGFk/a9e8CsCTKV7vFROgmZptzwSGNks4
tsGtQjM9qiJZeK3cohSSI3m//ciG242ybdFHq12ZCSvdABoUyXctwK9lIkNXxhfT
E4sb3Gmutt7533TQtuq4WLRWmE6pS+AV6IXFRDaP24RDstYCu/KSsdV5Eet/cABD
uUxyV8/zdvsb+UzddM/tfqrQ3FEMr1Ivsh7ucJKNA7Ob4UbUaUCgrPdW2ZyM3n0u
UnSFjY6EyceEtO+yWwC9tnalpaVS1r3IqrdOyKAtbAJOD9aH/bqyVuro7cfM27PL
60lG5MM3zAHKRxG5h33T6SDGso1JOiXKo92nut6AlQ42KukljZuZSa1EU4WoQFBG
8fZrs35XMgDjfDotHwDufqqePc5kcb4QkOz+Dgruix05JhI89oJss9wN7OQPpgCJ
UUFDXRh+gDs08lWwDv8bAR5byZW00Ss3g6bifXK1yRWkP3lw+ZKFi3nB7Y0Xm07F
AWdEBSEk5Q1SuxCvIntHvr/vpZvmwXIHDyk4LkVWj8Py3fBcQjyKhAew4regWBBu
0guhorxGqgyobt2VHKWRRthUTXhS49rbjRm49CDo4uXqr0wKTWRWpVCSWhbmDimZ
Bt+aXpZDH0AKoQ4rHFP3pDwmJbIRmA+xSFBBjxMJ9KIsiKNFglhN1kKw2VV+quOZ
hxwlRpAUYjVTn7oGiJBE7wk+PNlZ6gukXc23R9bGFBM/0X3l5gt3kU7JnN13ObMh
xN8FlPGHZE0rNGDSie2wYsy6nGO1qyo5Z3jCGxTMzeoPJbc6plNQH9sMGMfKRxQ5
xFVaFnRiZXIuEoP6S6d/BuybWOo3KptH6DCZLJwZ0NJFRlAH5sTjoOx/Avrn1GMr
8+lVDIKA9hrW5Pk3Vy6GnunbfvO4Bh0/amTto762XZFKeFUG9Ebxo5Jzvgo3KTHc
4EJoox/olS0OWWFaCOs1QpVUbjdTIkKfP5LS/mLfztiuUxqiR7XZgSXM+o6Gee20
6++aabGzIl8GBTvfq/mP2IFSrYuIP6uWji/R9jJDveR8p56uNDxWZA2+k/EppziL
ZN5Sz2OAlu5YIrl08sUdiOyEiFW3pljTxAm+jlPtVdVJGKfw9gxpWm1Zedzw56bT
aFkK4oBchUsOl3vJXO+rzu5WsHcbHKT4VUWJU/L7jIbn8Bs7dzlPk78vtRRoEVkn
+iVxmC7SywE4jdwvAB9pJUOXFm8z5Wu069FkZy0PeS7VO0gq2XtUhHeZ2JnYqWlP
3ZRrbAf20NSvNaee/fcERsr4H9jxV/UvgF358LVAJ6UACKaKuVC++w/KXbX1Vhvv
yeqtDoimPmFi0Qvi9E1oSvej0VaM4hxtOnY7YU4IX76FLe6HwLHvtIqH5xNWM0OS
gBM5Q9X/QUbjEUwK94UxU7SG9UW3dxYVSFahB+gLMT1ganpE4qgfSwQ5Rga7f20U
WFHFGCiY40jMGW6wPCDtZavCIT/Te1hpD6Tew/9dbpJe86E/DmVTkc+cFnI3kfeV
Ma1Azi3eTN9Vt3A9mva13lkVeRsbAIuYFI5GoxK1cZO+Li5YTGo8HYInHJYf9bgH
7adcki3k8L2JOEoWbvr2TiIEXBtTGNKhT5qIM/tGiqwafPcIgPnHRImPxWUuI+zD
DfzlsLS66sWUFB/blpEDJ4ng61h+T3CTi/SecRiRjZxuYLbfhpnmbSOzg8og1iHf
1yzU3Hh8IgxJCkGliUG0Wp10fujDy23awi1QiWL8p+HoLYFdpY2FHec5ICVTUeqK
Vsb4lDnAv9cJvjQ1fmQSstAAGNOVIle708l6jSbmjbP429teLjWzrEHkVBqrIXaR
FGjxPwAg9Y4MEXzcZ83/ityS8lLhcXMQTIPK2BpXbQ+0mzgIM9FpIJnAPiB41jQd
igcv5PPwwAqvicyqzMACim9S+WzOtjbsceUx5n6uTuWoj/o+tj0wakj1mJZY2651
en9BMDOijd27Op47OWO0OP92prFU5ArxIEp7+ufKySWKPpni1enht+SF5ALfgwa2
rvCSlAX83wmLPHO+UYUsLSFdNGtwx+2yXN30Z0xuVTFckm+wOKdkgp8Eu4wLoeof
nubLP/w6IBkQ+tRSD2ghwGqzoTRsudukxHEAer0KmMSGHY1loBJ0Z3MAeku140pw
nFroa7qZT2LqMlq2wZPGq260TgOHMp2wOEjV2wd1v7N6/NAWHGf+i+PdGHLsEp6l
urLsS/+Zo6+5Cnr7RkWNOqK4Y9/wOol0vyjlrq8JXMVYx+P0ygbusvrEuZWeAB1M
Dy5oDocD8gQ6mcsNOnqyhGMj2devjJPddvo9eM2ZcQD8Z/LhNebFK7fnQlJwJT9a
7s2c8OdxZueggJnQyD3677vJkyaIQrOuDvPk8sXO9kXv2ZSBRPENqLCVWjLfzKC3
UDh3t2eB91rvk8pvOlYw05uz3rFT4Y9NPVkTULq/7H2OBB8rsS5j+Lzez17GnIhJ
HcgwIzC60oQ3qTfi/i9N818c89tRyMdkokOtzccy3c3WxepwXgQQC1/hoilz7li/
DAmn7RULJ1StQDPcfMuzB7JzrPp2f2HKD381XWzBXrJUw4EgutfFszFhCNp6TzV6
/3Ms3XQerUqIaHbJI2iDbC01aeFcZMPax3quztTJTPqbSZA4AE9QU40AZv+QEKC7
gx9dlFouAz7/UEts0ZF7ywkFm0nlBNe/GwjoOammilLDnW94BJTc8Gb0fVf7v4yo
RH97dfy/nS/Y62IF/twQ+R3JOEZ4UbWMF6TXTUa+Wd6lDcyHuK/q4LORw48LV8eE
f+Lr9Jd488nrOm9a+BlbARCyUPsZwRrO5bfn0Dd+xlyuIS5uvNiCC9Q4Kb1NsYx9
Th2Q9rbKBAyDGhrd3aGfm5c/9+Hj8LlBe+n6w1LovEqxllmgWH3gVO+j37k1kOj3
lFSkQFUBmFuMp2wGh9n2B2Sy1rYIb/twl5kFLJiSAVdHLKfHUGUVt0UG340m0iMr
xekOgMC6SonNIpvnnrBnszwfizx2S71+7CUwUkDhAle6nT13ROdq0C0mHkXsHmG/
92KgkwYGZ3cdp22YtiKBHH+CFfnM3DzvJWUKS3yb8ngH2Vap3pg1pJtm9FQgQ4hW
bw1WMFoWwDPJ0lbd+ljkAhK2+3KLKcyIS1JEBOKTep/WoKPyOOea3/NvJtQwEPcB
TivRsIZoQShFOyqVkHpTa8p7cRTZ2haF9pzUakYwLE9SSgJa3gVMKl0oIxKoRAJO
lo5U5b2AiYRJ8xGD0BTSdFxUbe0HpedWNQMw3XbiVXFhBrbAhAgtVPXofTG1djg9
fwe+A0lqBzMyf7cyBdmZ09ddA/sFpLs53gB60ay8BHvS49OyfXfDmnI39PW0W8ir
RAfJfSoXgrmEr1/p00HKGf+dwdYSqlrcdEkBkjeYWqrvU6OaG0Boknoz3ktei52w
YXNNLFWqwzdC6hNvueG4C5/J+TpzFkAA+6P/oFCvg6zkxGJgqWggw64bsVTzqmeC
uAIyXOZhGfG/vtknqv3wc63NAkZTJ+MGV1w8LmMZAqZK88QPZeLtgETde7sOXAAx
E+5G+I3DLn44e9StAsJPa9xmEa7/+G8XDxHCSzu5dsjL58PktViLkblE3y7j5rJJ
lsdZqRfCbsOjcHrxoEJm60QBpKpceHnNIBKmLSjeqLDl89Uj6nvCG0lvU8RTcY/z
mBfgt8YvWriOm/WNU0DM6yEvfnybhOHB2kxDBfeW3ZoQ1fix7GmC9SrHy8Ifq70Z
hjmrxSjH7niNZn5cZPQVacHUpSxRZsi7/S0s2cwuuS+xld2uZUWnlWTcIbsEotCr
TU2G4O4QDf7RYmrWtneTSdT73pW92kjCtkFi2ZthJyZcyb0z0YOSk19d42cglLh/
Au/Chm8jTFVTXUBibI6zBzfEqOBSlWme7PyHHz8OTkUc15RX+sjTfAFiOOdQ4y+i
G6xlq0zHtT/EQXp6sY9Zl8dBEVn3gJSrfKT2wPHgjZl5Bei08h6JPVWjR6o6fi6L
b+8i9xJRfxlxmITB9yQBqlQ01eOlfKEpNGOZZSUJdys1LMD+Dmqg22AWCY4ijoo7
jdo2rhNYENoiHzt5HJZMellGP6cfRQUHbDB8DMeQ5CetZVkS47zgE4gm47kEI5Zz
Dwhg/bQietK/t8WpNHBHc2lij+xZhnlvLNtjx+t/0Wr8jWH9hm8EkMSvYHUIXTxt
JVFcdr8dgI3HIiG7padSsidtJJ9FyuIPTXQVS5MG34aQHRkNQPm4xMNe9Yt73S+K
XlAThyhh6xq2Jhkz7bXAnPjC/PgKNoeAZ2b87oCrkN+v0PQwE5wrAxR/K4Y3MMvh
rNjngO7YhudGnjZ5Qrc/b+FDtGHBkOkw3NfEh+gt37ojbNlAKzRMOL2LmPQcBI5J
S7SdXECnAUCbJF9AmKFiOrYCoDK2qCQYURlVCwD+c+MM8xxziZqD6XmttgYgpsZJ
5lbeXzKdOxyXa0tiTh0k0NmTsZgQ/tPzwBVCP98HDP+yIzGN65WnSTmiqLTQHQXH
8cRckYw0zigrCoWoNWI3XgMDtHsdjJdVqfvA+IAt153xiLp3ipB32HTKGUZ1TJI4
zFX4bklzvgXq7yOZI7uE1p6lrNk01/FSttR4HdE7dYzit0y5J5XI7ll4302OQqrr
dYbx805QcGxcmbnekzcdCQ+OGFiDj5bHBdHP0W1mjrak5sJq8Dcw61hAXLJpHQio
eBE2w/rMuTE6nRdX5hceA3ggDWRyxGar4dTz/neATZqeiWjLWPCFX5llF7b8HapI
lDwOHTwbiq8cOHFKSuXPL2eK6jfC1t5bG8rycq4DI+TBa3Rugayb7Vh/b7aAhZ/m
gdong3g36juxR/7Fu7Pk6xvZiYfUa3vGsUYo5Ld7PFSX+hMN+zUR1/2L+Thq+BVw
vUNFRNGD708lLLrgEA8MnwPbmN1CxYKYABG0RZn2vuP/QD2PC7+eJO52Dmn9qvzX
88xwPZa761yS5/GrpptDiCMmGVWZz5bsA5wvgvsOMEraT6sA1NaZA/+tjsfHen+n
FKBfBAmExrfZb/7NVebPkHlZF8p1WOGxzVAVNvZNIZYhPNXPL8dzVcu/rzWEz748
CdOejbvj7775PR22JnD93lR2+zVgqWrQj68Im4h9deQHjvaBl2AEeID+X301wMmz
4suwnlhdPeOavcn+kXJEbFwMrVfLekoBuRNY2cB/lPAIAwMrQ20iyn1/T89iS4ex
8TuZJZTKQisbjFi3XOfmObJ4UVHizLIptf5epT47kr30SOdowgIMjuMBkt5prCeX
9ZsTia3B2lY5DntKqPoyUG5Ssmt/vSJrfpj9dvAwWVFDEMX1XZC++5497pckr712
27exd8XsO7JHnhHLxbgpcyyU3eWHIuTM8kaHhvPPdCHQkJpqC/Q6OiUc639MxCgV
XpE0jVMB8ZPuBCxoxN1BmboejVCnSMpqS8t5Vol697G80KgmqCNupuqcGiJzCelK
Pl2lXnQL5Oqp0+AIPSJ6MeAetxsxXhvD5uAyAUFfp0V+SvKnj4XWbb3acGHF299o
vqnF6HSyWfkuhVTdGz9JZ9ydncXfm3lHCICnCnJvNV8kjrWkpWmkDjfCTPn6hYOc
1uG6NhkgTGGeg+/2dFa3N56C/r9fBsAv7nAKVq72gcQaxNk6vEjqwNFfRQB3uYcn
WELBBKIqneX3oYGh61rmwyTsc1x5BRGl2iDABEpfH6ZjI5Ov45z0Ao6bNwTodcYU
z8bKTppL4vb+GGgtA2lJsR7BnaZ6MVkgL0D5VL4uWeQQHNrGBtl+W7aeRQFgpE/S
jXc9vWe8pw6dWMIk81Syjh9IgGB/66Myuy7VDY27Z6Mx9LL/xvAP5JsL4HbNSEhz
2twZVbrCtAJE37GLn6tPe8WGGFx/soW7Sr93Z1Sr4dO+Ko5ad5S4/k6Crn58QWvv
HX5r/P01g4hLCV/oeYHqnI9DoArNqoh8uFlXvv3hE3SdcgNyKescOrtcITsI4oZJ
3e/3wZlel1GoC0qyHRTgh48UCUmxBOzVYijQPCsmPvyRSIBYvRgWjOb2yLfktImB
tFXN+ZBNw1jA9zHMJyS8tR2zgcUX9DsRm2lmAp95C40iRWfF05jeGQOFMFbfHXaq
UBB21N/0UuQykk98pgb6ywbuqOQ6r7FBu0wkGD5SZO52qwiwWPaOF3r0fL/PaZQT
K1e5XqWe0SEhhqcdGWE5lit9auYn4mayUYi19muKuEl7vwmNMlrBTN8Zn77wyvbl
lnsFJCRRoxMNY+FmZEeTHSqKwPRj5+0hIquR2iFgddNqG3uKSGW/CdtYxBAS4S0s
qJSznPYWp+C3/hJWmKmMePmm6dMyfDD6o6OgyJ3OMZfz9GMCMnbev9XW2DKxjibK
aI3h4jhSDvARmwEZYGBL3zoUbkISIluGFR0JGNXyBBglTRQ1oxkmLm+6Bx+8E/a2
BWnInXueRIwy7SsxTtCZ1koel8sA4gFD9+Hh5ygA0tnwVZiOqxBu6T8NzpsoHcN3
wT7evgpqNH/WTgfGKGB37XEbVdlkvDhS+y9j3guteXEZodXuKSOo5uw7y9U4cZLc
kvE+9ZPtnTKcyMfsjqnOHfvHm8xqtVN92iDTPU9Lq2v0bRpoD49HSQnq2Klw4XjL
0Qofgf92RsXUlyalWD3RnisUvEWAjzAMXbM4R9o2sKjyrM8S5XV4pzJZI1e3WsCp
r0fvBHO8864wXuM+kSFOahDFU4Lbk72fiECEtg0KZhXxlhCunf0thX0goDC6IL9w
HT8ZNPA1QXMYC/hwGewqajkZkZ8zL4qlFJfDcasDCxmFaBWZhSHLnr/ZvqXyNorv
heIYtF8NqsfsvCH/KHkL5UOhMcJAAKEohMIZL/CvOJo4Gl8WPV76/JLtvepvl+5q
l7TpSY5LjWX+kd/6tS26jWYHzz72CS8PAqO4pa0krJqQFxDOzrjAZGO60iJHUwG+
JPFxxlk4iR4cH+WsUQNTYHtQtcoeSpr9T3T/aTJW3hX2Kj1Tm69C8VqKbqgUIqYZ
BlUsNZODskD4ie9ENfFl3MdGRrPNKz+9XEdW9dMpGEIXr+uUrdCB49lVIXn2TPSs
ySvVxwucQwjNYMJjOCsu2RAsNvD4Q+cwA2Ln2OPdt3S1Rb59DUZxdNzvSRsj3pKu
ZOxAAFaE2a6n9YhCPVj2m5UnzFa+/aK1mJBGxcjxi89C/cCxqNjBbmowYfsPogn8
lcAsVYa8f/ck8fPf6C9fdLjui705rZwNwRRARRZ968Re9Exww/smtGFpuYAyNTY6
OMcXVzWinrF16V9bA+G9QbpOuwHoN1BuroqmXS1yTPQZnJ009ide2oKaUAEPKpiE
I1GQ4+L98OLCHWLh3G3+g+s29xHMw4BjcASPTbNBWJPmDgG/byaUp3KJLk68RmBZ
WZ6Yx8qZ5hiBi1Mv9qWtCMEzk7B9zeHMH1atssE96HQ9n+kC0c2YO+hsj1K2iwKi
rv+C8WHFbKXElVQPEFfyTi0FI1B7VM9dkMEDEhm0zQJSVK/PI74Wg1xObIZFUVx9
B1jpK4+dZlJ5HfBLqtgij7wt6BQu8bu6pBRt9P/PQ9rZae/EETSZgWdGndmmfLx4
uP8VlamCgxREm0KN4EbBfCtN8ahSWKzATYLXnFIckPgPxg3je0o3oPMPdfDpDD+z
lS2eG19NgP4tDwEQt56l65BmmrYHC5TFdoDkA1hHE3Nk0vtv8cB8k/sA6Fa4fMtz
bmLfqbdn6fZAVeNHE2mh/gRAC55J0Ad1jbehl76eSL7tUGqYAARcBHPqobLylIqx
cpBCKMH78Ps6mtHFJVoP+COhAWEM+DOEcKM4XlRpQ2w024DBceNM3wU3zv0Jxukw
cqHEt175L+d2EF68647hy1JQt5x0py9DeTPoEo/HtLjV/OPtVBDHNZLKExD9l29U
DoeY9zHaZH5DmMGYueMH/705gRrey1ywYQJWnPDLCJjFErj0jiM8BwxaJ7GB0Yyj
Y68ZcuFss0JjSI/5RolwHCf+fOQgj5dUCnRRWtEKidKTjkSmxamLNa+rddGxLIlf
1+RLCPd6CA8VLxWVjBvreBYbBXhvVj2wsxQ4UtQ7VH8P3uIXiqIJ2QnxUIVJZ1Mr
WLSXvI978mCClv9NZyoH8DgJF4S+4S6BRqUiRu3OFgjLD0iDEJUqGb+aAEBZLoEQ
dKcgTMRuXb9XJzLcTUp7VEgMv2v2ozv7w7w2S5Kgl88gBEbuVwjSvxg+CAIYV2lq
JLsVYcERbxnoonvKStDs1PdD21UMwZtvEhDczCwKRaZMi7ifmEZBjwfEY1OF79Im
ZxNKZHHrJqeyaG5n0JwK7TYsiiYOgUlxiM1AJKd0rcWFqe05dEsGeaunYrrsjWYC
PZDRyRqMDA3HpTpJKaok3AvSiu/wntYBxpSI5wdjwHZRNeq57gFui+BEFr+Iu6vt
+EQO2DC4Gi1nfvNQBeKoi/sIY+RIj9aeDBTI73qR0D+K7fmi9VpoECxiLAqm+pfM
kDFXDREF71fdLK2gb08XGfkJsx14+qOd7WxHeKQl+zCiKK+bAq2Lkjz6jHHYVrkV
HUFw56/lkfxnknbU986I5q6UxbJ2cyXRX5fs+Sw1Mx3mMMANz1O6StEzueYcwTAq
DKrddIUJsHDcW47iJFZSZEY1oA8afO8IcgD8CuveaDMD3ukciiaKlRGHz70oZlhS
dCrljTX8CAKU8RfO1IEnNNeUIX9ssnZIh4c/9NtyiU62VGg3V6b1HcxgyLypLaBt
tR+3bUCpCtMIq5zr+1EgFPnN6YjekwsOnxoqw6TVJmP1Q9bgrPCvW5NFR9ZJmn5D
C3qgucYoNkE8tjargyZx9e0xnaV1V5kGN60VF9p4ZCxjASPzvflDYsKd2GZwDdLI
jz8XSN0+lCSHFmGvzUU3asfiw7KsGcs3yh0yHMaKKAdtWQPj1aYb7d/wletRj9eu
BQdwArdAXrhcgfliph1mRG1d43ynGYLefWtrT/bQHW+dSaiCfrWlPuMl2opt6vDK
QdywW/46QIW+/WWJ9cL+azDDhDDz5YdPDSTuJtF0n++hAgnrqvYxaKPXRxEjHYwA
OID/NT38BxLyCxws5oBLX/3jmnk3vzrZWKfMP/AEkttmKafKpYqAVl/b6I2VP+Wn
sibrXdFtKvMkrUQmtztuIP0r/ZPCpjwWVHn2oYXzHxgIEyFwMMsF9zeLSV33Kkfu
zAkJfOCmxQItzptCXRdpsajatLcf2+K2QM30HXuui22V5BZhH2+bKIjHg4sHyTzu
KvaF0iBKfxSyEQlAW7SxP4fN2TCb0NBPO2e3WCc9YsD3sp0Hdo3qOdkmei5eScrW
zBieUFMV0VKliwmg9RRlfFLPLQTaRAkh3G8t8wgd3N04Iq/w0qPxzc0ifTQ4YYAT
GdClRFP4TSLR5k4J9SZ0RKckme89lMiUk9HhTuU37EVzJrKs+rTumzB/ddxMrwYG
hd6oJ9X0RvG1qmN4wZ4SXgCuiIekCUJD+5FwvBjT8TUE9OtLgWT2/59UiaL9Yj2w
aY7NGUOa0hm1UKyy9phqjo7nWx+mSuV86y6jn7l3QqQ56dAb4P+Kc2688ZmPhG+i
xRnVys8+nXexiaXMDQgX/VkQfp5zWuDQacTx33FrTTRbe3Q3ePKdeo3ji5Fj0kyG
imlOEPBvnLoH7r/4LKc+7ayRu6cLng+zRLkKPdbhPgEIBDBbp6Cb99I4ByNE6oSS
mJ9t9tlQJFPg4ss5xjip8Wvi0VG8mbtkKnN4qOb0Mf5hvtwhxzmxs9P1GiE2kZt2
MXPoTZ8uNwIQ3AJgta8SDcJVigwCHPuZtKPb6LbZoqWXnteU3H0bcF72tqDeSgjX
LCiTC/BWBYwZow6j4W0mdkfyd64+gO0f+B+oOd4vBZKOOdVhuB45nBl/3jsW3xpI
7ZG2u6KnxxtCDg7vXSS3Xrzx+5g1CRA5THqzqBtfOgeenN1ob+/g/bgsIY1z1uIp
ODEjNwE8qi6+d+pEY/db72czSC0sLdfxMm3yje5QKguzu/CItOvDlqMEb3NpPMCI
XYkPOjPA9G2dzVYNBp3niK3hSt3sLjk9De16T9d+St6046Gxjcvaj0tlnoy/y5a6
hpkjhXBzJElPrcKmdW421Vx+XZtjPzxJZ1wqTPrGL/F7NI2/hxPjqKNIJY0E1nVl
pCvnXqKEtO6fkM1K6PgaXw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
eaHFuaStTzimKHF3CctKIyIMpCOHY5uZeb6GNpw72FsjWbic6R/7CVFLFnvGgegw
dIeDIRnoBBdd2bTP01qSrOtxcFhoiwuNMvh2XoD6EL9Ai5kZMUEqhrExsD1SHF33
odgBe5xQ4DVcqZF+8F+BVmjP3BUqdIABI7jxlKWzylSjtt0mj5C+dYZKTMCTPLWT
zsRhswPnjvpa2STdPOjt1uE5tWCfhGQC8KIBHp1oPB5QmWVRe2I2mJeYvKECp6RU
b0HuNj44LOLRprE0VvNk7hSLYsa4qb+ax6dL41m36INzAQEHRwXdZWfaoQU31dSH
0VcIRurRktly3fGE15WW6Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6496 )
`pragma protect data_block
1tt0ef+OA1LxRpL/sd5IIOdwGNUfkjQs4YCWRQXE7rpylBfYYaxYEfSpYjLAX2pD
P5U9FmkECgmnK8cmlQBJJD8Lfk7l4YPhX7uR8i4x9vqyUpVhVAaiEfoWIYlo1MBj
8xaMd8xlDHTis/Ft3pbg3cA1Z6XuK/B8JCLZE1aM5tfqBR1sM55CtYwn0p/EhI8V
y0H/KPmN6g5zM7Yf8Y7jrjFxfuZR6kTHvu6A0umL64iPEwWkyqvkT1qx8liDjDvP
Mjp0INwUeFxmrlBhmEpW3CKwexu9GRANNvc58H4MJALJF2D31fpFKhkYGyuLDn7N
ykXoiDGyD49wrKcdBSrydyDheXIaQaXuXd6U6TgTDFi7BmRXUa1H/RMTA2+ldGop
CwnX9GeZreJc5YLvwhQQP3yPOoQklmyrW/srL7S65CdvDJ9yqIeDi0b5p7jlxR67
H6MybtG0m/8SDeqX0JKrS7+ghPzVum4omxA/nPhP18cfU8F0FaugcLOulk0r2GMf
xTXgeIR+d74w/Lb6toX4woLTeHtkerAXAG2bNETttvJ18ikq1McDCrou6/nC/xKN
tTAa7dm4zFWFBmg4cBw8ZPLCRHVT5aF4TLDPEF/7zixoX3refeh/3U1WHbZfzmq9
pc9CLvwS98NCpFcI7ybVqA7lMtaNGUn1swYGGK4bbeCY0Y8N9UTf/ZFDcoSXFQMb
ESJJ1XBb97YRxjrC53MJJ0ohV/iNwhPfp+7BWgEurFB/sxJH3jLQnhY141wELuYc
6bafecumkFom8ODoWQWGUKUAJB8BJ9ijXxAh3f1C6ofZOjUW1oyPEeboRUKwPmBA
zarU2Uccn+pXa9hIOHnpG4XlD59tF/Y+zSxXMioZdkx65FHoXLzRDkV79Y63iPPg
2Zrnq6lqOnO24YamXiCT4j1msNiI8mkYqXUvZWUt5QgGdyuuiWZy+THp9i5/TQ+N
ZYNQzOIrO/DwdHtRr8yHF6fSp1P3x8UlefhTTTtQIRTzU+qLw6tltEnKKV7H6drG
DaxfuhXNmqMFd+L+S5hPKt4UAuv5Xk3Cbb3gUKvYGoQwxnp29ECEHyVi6G4yifG+
yM6OyzATKVu5eGGsBqmM6C/07VWjfmTLpcoqj8zwn4hylGRAugJ/UlNfTdgE0eOH
RJ2Y1pOhPNKbaU4kayTwtHiTRLQh5+LaJl9+MJyho5lXDWbQ4Kvp0fuJB0gk9UOk
h0feQe8bGYDcbLib6E9x0lpT7HSS+Yc/wfundocJH6Djju5sK/+VCzKrkuvSa2xS
shBbhfd+woGTSjhbCrZm3zThYg79AE3UfAKk0Oz8GGFvtz+gj2SqaORKiPQPkSUx
KVi2OTtFaBGeplZqgDFj8vFjn4jIZbIh3xJ+CxyVuG05iF/p5E+wldg4TgYkYRjp
Qk6S6zG0NG0wg6rnySg8W62ut37Z+dvg4uX6ARAB4qAtO+MCxbBEgVQRHM3zq9XJ
d00YJ6a8FtwYhTg1ZjaYtwlrGf6oqe6nZUxBXWdKdhJJO5EyxUtcP1228w75gNG/
DtG1mJkaiLLUTSuha35TrO8D3Dzxvfza1XOEqd+XnB63ut/pSJK/36dOK/N8pThn
/1xIeGMcpJWZev6Pb7seogbrFfaQS8aZkChNlfQ0uM/7/Tc0CG1DgVhVv6+CJ8x3
JV67GbFOroBMU7tHPTj/c4Mz+i8bctwb3KJsjO24hzkT/U/MVlyeMDwbdr93MHKJ
R9H/hpWdEsuPm3Rwhsa7DStkYu2+9ikYvigCCy40EmRP+weVOYWIdKVT2X2rQSTK
i3xePq3jjwG9LtNjhfGJHFoxQXa4s/MuRWYv3+66+zPU3+Sl4yQHGSEc8ud8/Ucs
qY7Dmm6Ma7XMfaK5GepSiXWsHi1CwVaN8pI0U9SbT9wtfo4fYAuQSNa+/2NThth1
bE3qqIkJv++vWPYtOkccIW+ErUc0GZGLNR//mEQjYbFZ5b1qOkm1W7zgi9ruJ1sT
cFUQb9cmwCf48eCis/VSYOHClOfe79unv1BXkFdMXHQQ9Xm4nHEIMY15s52aiMGh
lRQb9Bm3LwelPrCtbRLMIJ6JtfLoLL2rNTA9aZM/Otodj2Wn2cV9jUCGLhvGaNBb
kXu2n/HdTwARkt+CQUi3W2Sx+4C69hlfR70twZ1YdINYjF3NuCRAZZNdNlbuWsNN
1LiAV2Ge0hBTBReVVkTHBH+8IKLMPPrb2r8+rTqZSusCYHQ+rmfL2v29qieZWwiT
rt68MjeLvW2VF7hWHOOBNMH88b1DCuekFWAKcj1XI916R3w9iLP/j771a9i8VgdM
DnEeOvnOqTzVeUb1GQPllMkYjgdMfFAwZsG5zJbDXks0JqwaRbuEb6pzHWc6xxu1
CoDogpLSbFUIKf+Jhv2Hse9kgAnPd7ZvqSxsGuce1EHgN0PQsPRuegzsZLdjMqkI
iYTJPI8ZaX+77GyeUuLolZBWZUi6AocOAXlePcTVQ8Izq9c0Bsbl1qGyIS7dYoji
z7VDHkq2P5gbeCmnnZMwkLiygQiY+nDoloW1gzBFMSFSkQ4hU6vGBA4GkRCd0P3l
IX6Jdmj+YqWw4FveyQqtEt3yYgvF6i1FWpwGK8CGKbWAeUIhNHAB6gD+dofzQo6c
uKAcR7hZlD5gs4/2IQLRzyF1Xy1Laudxi+wcGyBZt7VK1/svaPEIwVGd2Bd74YBH
iDVgnOf0Vk4lxSW3FrUZpjtAR632ZzjWpiIAx1vvqvEiiseJd+Z7BcZJStndXWw9
wWdIC4KATJxt88AMe8ZK7lHyHo4UanyW51h9XV1ByXDeNfhEhrZjl8/1H/b3HTOO
N64D13l/0fsmLGSx4D8Z787DYBB3UCYPs4yNQMKVle2vTg4W0ApVfylS69TTdYWE
WETdECWMsPUeVmDM6PzLz/7mSG9znLZm55QSpeK9HTd0aOXhJtvn/QBP4d5rCQHL
xtAEZTuyPG3I17IaEoXpa8/dRd2hnB2m7+LJi7VNPZo7urs18CdI8pbxMqlG4448
HgFBb825LoGHfiHPcOYcdBaIh0DV1RvSQKhHdDTPD34pYNXWE6oLb0qkCdYTWmCS
dWDMgXfoHQNyxtlBit+kgDOxM7jJzAD3I60ISMte2gGzIdS6lf6fmok+Q4ImQ/UE
8CP8ds8hsLryomPGPKmkuCnNTin/iQZaH4D2VeAuoDfp8UpAi+AaRL1A4Nuv/Vn+
Na0HBS5JsFwF+E3zEeKHiwjSpbDWA0Y8m9neqS1AlSi354PH6e4LCE3cMS55mnRs
0XInVgJB4zidR4g4zANy5tBacWkI1AMnG1xd4AP7BQw/VyoYvBFlu5mERXIYlWcq
w6Jyx0C7QhXMctN3BVdRDacPVIaDIg8eS96W//qTPZy1NvTA5GIDPsbMZxsGwNY8
knqmKZ7LxnsJq2CRsTErf5Z8uXC8Ewq2rGKpVZYyNrGn3Eg7o1kMcWIhSNL7fCXM
lVYMvC/hr7Qrczo50oCf4OnO+MZ8yIYj09JOTLNQJ+rSA7i9XeG4D+HfGK8/zhsh
KbtjdoaUssdW4x5kD9cQAOGXMHJZKgGeLCPbM+s/goa5sL0Zmb3qPELZU4qVyXa6
cgpRJ85V/H+rpflHQDhrXypdJ+azWJDgp5y7PwgPEy8rDx2AWQ77EjJO1T/QSaZB
RYIsMf0F3MXfw3eYJ6d6l3EzPvMmjqJ/rMYn8UpRrRdVqkuRxxwtuOhkN9srB8QC
8Q6+D/v6XxCzplAzki3VwQJHdBJTQhxgb4kc9Y6Dnk9ZYoD64p+ePfuH0/mnhDEZ
NOvEBkL+zgy8Xhpf22M/F2BPBKC6cu3JgS01/1iR9prdEjTz3WgROeUH9jshX/Mh
Y+Xm6Bfp6CooOviMLCRSF39DnSnxjgs15VospHcK05xq8hznSfSVSHIntZdjQYD5
BlNU3sfSZJ4fGUgaYcr8okmclG2P7qLOhimGc/QtDQ5D2Z/xsVBHk0Okkz0MGV3c
lCjKSHMMW2TDQQGnh5OW2gxczHadtMuQWTfv1ioiO+1xw/hCcQ/e+RVqw72RzrHP
Urz3BgtsPCj7PMEgT4KDumiXgcX3t5W6ta2Wf1DgfFOGTGKU+Bk2tmogdvQhmhDp
3Kjy7fCZ5mY7hS/PWmkgfY9iKtVo0AdIiI7kwPwQBnMkuU1+pqbGXmJx21R9pv2c
/xnfsU0902TEP74sGmSX5M+wuCE0dGMUZO6iG4aXn159+DrL18rIZXMECGRV+A/3
FeskEEy4qIy1Lshd1YZtWGQonv0+CxFqBO2EpqjEWBhR1PmMCrdTCRoVBUcTGs1K
V5wQe1CDcTnpMOwg+xswcrV+Lv+k8Br2xqf3PfO2Da1HswNI5Mu4bvwYzGhZ4JY0
6gKcFpj+9iFfHDCGEhamLDLt693vOjfe2ItEpAeDtjihXG3w6JIMlcMW6xJ1oF5r
G7VnWQJOBvvzc3VFTm+yPcIAF/3KxIPWIGj/pYAEJaDyTHiqwII9lnWDKddUogX1
BpQUU/MLyloOr5IbR10Bi4Xr7L+ofrVq7Mn3HYSXXUXViDxSLDH1kiQfZv+TUHGP
4s19JHWCEsKk9yw9+YPort2q0u3N5X5K3yWL2mPnHvoWXBgmblkW9XYt5XQrDbpH
s6al38c3DR/Flu6Lf1IMoIpaXIAyBLpFUNizfFEqN7Q1wSoeOeoOMlN+3/RGywJ1
6re3/BfbfpqIamO04T4TOB96SlUP8dwEwX3xrCYkTap+nQGSt82ZmVlH8lBm8AaC
mmHMM0DZH8Ija8tzEvhJcJDwL+LHiBbGKPWk2JSbOOz+gQXyGPyLlc5WU5Lgjc94
1sN92wX6b+lnQbkoatLfZY4zGtwO3OxJKsb0Q3Fyuu4YcgTV5jYyMhIgW5Z8OdiT
X4QqJBv8brkpQeUuwiIsLkID3Ilj8ugXaWz7RKptMki6NO16Z/qgUCWiWlI9zMtK
y2EY7CZNyQuUzewF4MTeV5/EOSy2/TnVbwK7cW1sHeb4bI9/dNjZfEDg6zzfl++f
SxcAdIBkOQ7SFgWLorlUCuBqoF7px0pmd8688KZAQkMOX0bOgQs3XBVXfzztYCKw
1rfd/rvqiz/a9BqCUM/pTb1AfsjIKwL9vsYqmsPM619gccrcBRO/ISKlAlIy7y1M
t5aXlg/v7IVX4tbn3RhdLIjDO1Msh+t7jof/bpj5g/ij3mfEGZ2cXMLTEsTuPTeY
1BQEIG69vkpJPGborbejug642nEcGWJKdEdAHlWnH1qvVpsAZKF5Tj+gK3247oZU
2DIrbcqnuZATPRNK/lkOgTxeemcXtpx3/MaeQf76gzLas1+5ATQXK3xKgjHIHTuu
mcQEtVXJX9rrkpBJrd/DX9dAUWmVWNmq/yGZ1Bgv/yHM04yAm9K+kj3/OoHAPpRk
q/7zOT6wNrwdho9eHkyx3yKK+KpvUspEy8T+w5gEYNaYIhSj3Z1Rr3AjMgI7cwwL
kYxbtBcldVRkt/F7xnDyi1GtT9QOAY8pTkkY41bewzKeqmqkd5aK3+erJ/PqTJEC
+Ri53WUbMVD5nDoRkisdMdTDuns0PqDimQL1rEhyo2nmFoQhqNFHnPaGvtRAyPNq
c/DikMYqGt0MtoxDTsGnkEiVOV168/GVU66MK1dRxHl2BRLF+nUflm5pEedqltht
jw2of67jAVGae7VAQpKozc02snG27WRKJW0HTqkTvrXr/CIO2BYnd58hVFF8panF
thuE+r/xkI4UXzQm7grIsu/44uaBvGxZtPoRf1YI/YR+gCYhW6YGBQOwuNrpzmJ7
9/KNYkwm3ne81yEyJXJkVpg1TsgPoPVQ2aV9iy9bSXYndfXI9N6v8n5jCIXY3A2W
x41EH6/00ihzC1XuOiB05NxEQvRbQnZo0MWxbI/BxMWij5ig4/pLvS/sm1/A5RJp
laG3YOcnEWka9lzfAg3TnpMxVSFL5wB0I5lFtqLiMbq3pfxwOAdhEEKbFygPG53n
bKyDSlN00SuyspvBH1sVbmDU+3e/QsKifa/jNKU8T+ku8u/+o5FJH/W9i2dF/vDk
+TjkyEz5LE9D6aVbSrNQ8KWQXmNV5TldmtpMojStSsgHK0CGFjqItyGyuPU6J598
7dc7Q0rDX3nVfIjeNVw/rZJiiA6C7Q3s9wSWlxys6OyTGy5xfl2tDgBO1tNtGx9l
pOVjtHgLmBwhfXDgNfUysS1LQww2HYP5icltSXGLJOPiisupMjPFCagCJ++AwG1p
Pp93BiEK4k+waBBSPueel1+6H4xBqYyCdaizzshoDTf61z7ODUAaaM/BrzpSM4yV
ThJAsZWnrWiWN3fJ4w/KAxUt92IjDQkyIPznyONSHt07n5ek3Z81syOWFA6tjEI/
dBziuB5lR/QJ1A+UdI+XN3fRU5oFb5tDgqvw8LzIOgzGpyOvkSRyVeK1O0406b5o
DRYbMb3zbKEqO3kSnhPuprw7K2T073uJcSOcuWgk3pA0oyJVOGUOU/Mc6EkhtrDb
GOejoyjyu7VbhEzqvbQDG3iaTDLtiU5XhIucVYK5IqGDufvV9GIadx0jif5QV0jr
HHPQSLZerYtGWNEnRTRTFHkdIZDX4V7mK0KZExWRQCbNso4UrKAFUeSrgp+ngSxj
tYf/GTLQimSU9kzZHZwcquvamm9FYEG0RTsL1K7To/2lnGEYlovFUI/rKEngzu9B
k11XIqCq1/vctzULQgUxNIUmW3h7qbkRstPCHi5ksQVdeljWnRxEq0nrDKeoca2N
Wmog4h7xAKj/cngvR7UGuQAxRVd7UzNosviqPsWPf/F8MFm/b6NXSpEfJbjY2o+D
7xxgiEgaASvIFAwmMRWjeD3kIh0UCmSlNSNAHI1zBirw9/WfmDhtj+Z583zlnP0+
Bl5Ve57m3aWwP35VluDgQQ6zNKhiw8ak2/tp8wlbG4fLsnCf+EIEHBi+RqAXFD2R
R5GVELNhmROLy+UrNuc6srDI4E3ZSvGk5i7e06mpq3Cic3aUpFkqoebPRgceE+Np
jL/Yx06P6Y1KSg6JR7XIDd5ktYqxznINaBuTIhj+2+CpCaxi/uR7xBp9j8MkSGvH
JaHH0raObJdly3h9ERHG47s3w/FC+nBYsnDvUyWkav7OWAnK4C/+KdB/7+Zoo5Ew
W3SKvcSgBYGd5YU1YQJT/eZh75AsihfkBhUtaTIsbQeHOwa5FTqo+9D7fPzWH69v
OmGeJmFzCVLysuAmWi1nUec8MUz8IKHxgmIVrf+XY5eBXltlPwpHqD0/oxpoqX4y
c242bT4D2JkC+t15HCFD6o2O090YecgCv6/2CNivExMKi1kN8yt8eOCjS8f1MM4s
tKXjH+gCiUrmG+hhrvtrp3j18sGwLbdUSTL5nWsZ+bthSyX+b/nnJurNctfaJ5iO
fPpjna9gtkCiQet1V1NQg19DuveEMgx21zEB3kSNiy21vXgXkBbpDv0Vh+9MbuFu
myQXWZhotdENe2wCK0R+hbjfc1gczDZcyXmh8R3Dijv0hD6ok57jgtYq0P2rmRWz
VA6Yo33VQY5NTQze4DKuf/Fn4JzZnkYcs5VZCztmcaxqDR4oFCd9sdrxCB2geBAQ
fL/ez/d5BZsxdocNGUBLwS4ImbU82Mem9TeJUjIOmFukcJubrvX6k5hqqZ21zNb2
j9Z0AG0ndC01jViRgeHRTvGGLuXXO/GCmWlMtnQOxu3PgfpDnblFbn56XzhEtKrT
pBwoc7FnaIHv0o+YE8lBc91yMsflEa4uALknabmaM8K4RA01DKHWy7Xfy+arYx5k
9JGDZ0pNyyVlFU5i9f62LUlYftwpnWhQFQeeffXRLk1g30UjO2ATYov4cPOh1rC1
5TmW/1roQ6ppF8tvuidVly87TWQJ1M4W3Ft0ytxDwzjnjrqLB2S3mBAv1Beoydlt
dxilUYvTDZIV571R1XvRXAnvLN5/fcsiQichh/eeVR0eMBop7ZPkYPAyKFbiGFcK
vyJRYOGf2IVK2cBYKa3ryNDkaNK2yU8oMupeUZXaiBBhjzGhh+0PcsGRVniHygKN
LoUiFMqwVXiOvZ3JVm/z3xVoCw12kb09lp+sre1xzlVFMkI3NOATdyiVIobOLTJU
qBH3mWUbP/vIVGfZ8ElvIIAH2+2Ij9UTFZsNklZtSzqJ6hquoAJe8wqmJKg5ADAz
ybnX9Zp3dmVtQNPXabo0+vO8Z8MGZNBC4ZN8NhfKicEIPW+AlPgCAw6PrbjCbKnD
nE6Nb5NTUkqmAcqAia9nXnRLn4ui3z6Ra0DiXao+nEUs4SoEG79xylFsFMpRkM6L
kGrezPZRQJwwC40mOXchGkomtcRWUwYz1OycwPystgi2B2Rtx48uUTZNn+TTj5XZ
V/2AhsVgUyo/EstEYAC/0o92zgWupuaP1kLgYwyaS8FoCxmaaq+PLq3VHhqI3JBf
fRbaLdxnZxbVG+NcRpiphJkDrA93wPV9dM4GuHlQJt7TNt1bzEGa5FV/yMPycbJI
Ucq7OTSXCV/xtw+jSzIT/CpVJgqFLq5e3ezLrULhK+S8t7ocZm7DKLjPUepUxJ8y
QW1Ofs6OmIjKwCrgwXfc8eOffnmZXdRNPyfOEe+GxnVJhJBpfQP2P9BpJMvZGUFP
/DNGqK0d14Q/MNXlOuOM3eXLxU1IRD56c9PAF2wvxbmM8Sb9L9euuBJZjuJZHSfW
urHToPTpyBiMqqrdQ7q4kw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
eJNsRztOvRA9wm0SAr1aBSuoQle1zZt1Kxgck4Ti+bxOKmKwMtlr6rgBI5ukzlVA
QByPGj9diX926ieL4UHzO6tNE0qFE4HmYXy8JIQDWmMVlqQ2QMBVJ9KRlJkaEUC2
rBfg1/UJXQWfw5NXM5P+uMWZAi+nZpRE8dImotFfCQM/dPfe2z0n5VHpPpjIA0ys
OoqOU2uQ1HDqCpIdsEFLI+CrHYvUaw4rWLvCR3TmoKoS1SRf/cJkeVz+MPQ40n5O
vASCJWNtS1oS9u6npFWaGNvibe54+Rrq0iDpdwrg6UYKN6I8tqfO+OOw1SfscGOg
dAikMnfSISNwOvQaauOs/w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 23728 )
`pragma protect data_block
3vtUpZrb6hFsGXnGhAvfLpVjlNjzFyQq8qleIX8T3qfp1D8ueKBkV2FVEJsFVdlh
zcty7czq+XGPEdl+KMhLcBD9Inmnh74/ntGLzypQ84N+/JAN9BXMwqb9q4SHAl8w
5UcdcB9jGYzgAU4XVcazjKEXMomfCNCzmlOu895lrcaHP3naMAB0EupK1VU39i+J
8GucFokuMXKBl6/O8BV/4mRIpPNrAxraA1BEBM1AWyUCgX/AhZgU3wM59y+iVTQ0
xlKVneXm5q78LU7CYDHbX5y1z4yFBOQBHrh0G72qPh71AVxia4l0f6QqxLnNdjwL
gzxI3Sd3nBXyD7DfkcOHAslhnlfuyyJMZGdPqVhka3xxhbd6MXdZgjFB4Gwf9IpT
F3eg/YzNkry37fBwfOS2PwkpEKDZo3aEv22cMbRPAf2J+wDk1nMBFfjVrRKMWjnE
q+hJReMjrPcUAKP45iISzD/hBIVmci50tLQGICXyIKo/sMTcpKLV76t68F+pM826
OHH9SHXYO9RFnV+z899Eeqm6vaKwUgph5s0fYqLGXYxjgBZy2SfnRat1PY0DKKjf
3xWbRN7cgNhf2bSBZYTXefjTe/ArepRdri6aRWC0//TZtqr8ooDVQqyMvQS6WWBO
fCyJQv+193NeRRNlwGyRU+OwE644j07AufhWjjCS1XD/QKmhF8ZSAzLp9XN0jG5O
PRbuOPJzCWpKs7HJ50y0CWFzS8lTcJDEaKKLv6yA8K27LfZxlA0OtbD6vCy9nfBk
VjwuS8gYx+PFqbgotlE9P0NYHAKwVhV7Zsh/RzyyZETGLlgJixQl6PU516NOjZFr
honA1z/YWkLA0SPDrDgaA70JoUQydxhJ61S47VVeOk0FSCiUfQXWAsx2inpaItCe
7dsYhIVtZKS1GOKhkQdNBZAZS1No+SXNE9A7qC2wDdhlneFBiJfsuZuyNpAWuVXZ
O96kz4SFzjGSpEBEFTMsFcmKej1WaPtITbpfGgmFw8PvSo1uWomDGT67gs8pXhEC
vCac3gQwomenLoWRg9SzFJUJvomLsDBWWXIIdzpU2TXGDAwOXXhlaK+Sp0jVDHVJ
jML7zFVv09+QrWHZPjIaNb57bgNho7aOdS0SII/YvIUWLIcjgmk1zgW7rmJu4Lsi
OnpVJV1YLQNtr1Gg6ZPt7qyLpe4zMPkME43qxJM7TKMsE3e6ljoLPKOhk7xqGvd2
PNJDsVDNIJt4crTsquClySGDJ1hkGGmTzxzKe3RwVqFfC93OP5DU7JO7eCij6Cvq
tdN5hb+ZUuRdWpuguZC1iFk6DYbozVX1FoMXKFaBVDuS0JAL71zyjVEpg/RST0Ay
Or5aJkkg8kQ0VvVpE0cxyukE/E8FxjNj7mKnF7JvIIK+JEjI/7ouOb12eHTvrEsQ
/7ht+axx+7j2GatUfmuELRPcsduxDIcTRPM+fy0KgB4QJvMlEwMnqiLZMPQrW0qA
ggIeeTPhJNcGia4PsYySEnAHeb4zaIvSqmfmuztlHLEhzRYg4tfkblitJ4HNae75
lPE1X4kt36Uw/CCDVKKtaOYJOuFFQKAsEd/SunHJUIarPQgCNjPLnH/nIbZ9LJC5
7acZo5ZVq5KuDoF4b9FB5z6h3PrbEywU67DbCGYzFLiOvmi5nVwL9Pe9DSpQ0Sga
QCrQ+0z+ilNbsCYyaG/vmH7XFINYJfr6PS+CtmPXm2JanSJSpd04t1NvBOjSqi9w
Y6UZBOuGClak5Ivf489jI+tGB6J45dNcZj3B6AY/OAF8z41vP3ECZwd5RMTCYCb4
DjS4yknDGhb3ghu0vpADKdFv9dApyk6QtDYM1dYKOa9Drw+89b0bJkfhYwU7KT8o
r6r/VpjJBH3FWjrdD5ZibRX11Z9dASjN+p6HxxEOEtmYuYsnJ+0zzgkDRKIXHDZ7
35kfIAKD7CfgVGsEm6YLOtxxaT1Q3eNtkVOwI4ZIcffkiRyqZdjK8nAcpR0yIWp7
c4AHnxoFaoynN0rTbYIMTDWMYfHWC1vkp1+XGFGk68r/smCz2mJ1b6whFhKIIsJc
H0ISl7Gy5YBEaXEp8l/Q1WYmhTwEUwZp7ogLMjn8cCycRlq4BrWJOGFFsPImXyJO
n1ymA/ofOteSCQ2oGeemb3DPcGKcvMglkrhCXN9mLBH2KN5T5Ahr97Z1FJhqjAbs
gyI7uZiFKH3YycjEnmHXYDEvIcy1Vx4FIyRiLOVgD7iL3+9liwBSOYaSwM4LoKJS
n7b3lT6+5Z7u0OKIj+FjIGBxaWNiw4QTjKr9+xOIVNwYOv/aeNpuLwDIhFFizOMD
1ww/Y6JI5GuAu1dvFH4Iz42RGWcW5ea55xyi/AknWQkQYXI7AYSX8JYA8j8QgUwm
3+vKFnrO+AGP5oP/pxP+6Zxw56pqMwFMZjB0ml4jYSQxBkWax1h2EBABqGJFwRrz
NIftvi/+rMlHuuWzAnqfXzlXIC7L/2JhttPnqQr+RuL4RUTUKSxMHTXPwiSlji36
NBIY5u9R7HDnfdzRRFzpa/ZcXHOlECBHxIZP5Gk78+m9huoXp8iBvEFeGcoEhHBd
PNCx1zJGhaIXhG4puzzdhnGwaxSFIiq4N+NPS089elO+gbodmo9OYaLIbiu1oUEz
uEUq+89JPGvJYoycFBMK/1RAz/hyREbfzeNNdXa5QcId5ZUPSg/3ucTs4lmn+Qts
9GH32hJePtQ61a9GwBMtU9ld7MdUKxt/yNseHITmAt+U7yzDiZ5V2ntRDvQibyHJ
YjftzXgjl6z0bHjJS4qcjz8A4KPdJBII3Gf4IMqV3YE1vd85jF0JWXonxRGqYAlS
vxJC8FeSmk+F5pLBT5IAd1p9CJ7j/BsMD0t7GNqaYJqHGR99b2xS/qxHe7nfKsVA
gRLyqnKqTQqtgrWtvMQJKt5II33XamgowVxitRMFt3+NEBp7tAde4OAb3hFpdj31
Y1lrmF5jEtEbbxDTn67JQnZ4ytY9TOnpHo6pV4BIrXlloGo8koUEKmHEnqDrRLSF
DvGfB+kLiKABayfcIVxzdLcbuacC4zj7nxHNxDLBOJG+WPsy5gjAWVqyIi10Rr9C
2HjFeU5WZpjIDJH0ZpKmW+Lrybe4ygO4/jaaaBlYvFh8BL7+mzW1hjv74GgrlZH1
cDexIdBCW4ltFhXoBwPvJSKdNF4bSv7zHTZx8kseoIHj/d6PoRRWnixDTeEEhBjw
UWz7nD0970Ol/SfQCn1OOgOIu7cION7pmehPdIyDGUvMDOEVvmNGfaEyHH9EJYSd
i/mnm26Ny6M7MUAvEtmsyiOB253LQr/2Xuemi3nQsYhitCLV2UgUaarfTHxLbxEd
LEwctpDkIVf+1EdiH0Lnxh9cS091S/BsFBE0C0IaRm+9XGBMLta8dFo0VROT/qSK
Npx7psLn2uheqM6i9fiODXJc4uAUYvvGq5nj1z9UQw4m80/uapJpHy+xDWR+3ai1
VOcInnVYc44mF5qTGevUPMFBKDy0/AFIdDw2+/pV7DTprQeWdaHAO2pIZAx9Z3nx
SujrW8OBVye33fHBbkAiDZVaBb/C6Eyt60EXU+s5fu/sJu6gJSWK0RxeX898EUYT
BFrCamKyfh2ymnHOmYTcIc4i6Nli0cQx9dqC12iaxbOOpeIcwg31/IT5EJ0do8Fz
bSZwOQbipNiq0q7W/OeSgtOgWajK3AK3C7NjWni/8E8ooh49yePae5dgZPK8Khbk
NM15Gi1B5vE7CvFHEFFb8rpKNekGkwb7Dgp+GCsvML6wE7/DBmgYjD3F9zgrUGeG
WMpCLNghPDCGXG434RwQH92gPmX+25iWFCEpeZfQlsm4UdZdbIW0p/6kYVK7blOV
tlbBIWdhft3cJGlGhcX/5g60JxGVqeK7thQj2R1MrE21GA985Yksz+2Ib/bkbeJh
P3f9E/sd2qkWSEQy4zpUg1QFq0Z8T8sa9Z3V8BIWMYeSV/dF0U2KQlso9F+dBu2x
KBASvAJzBIgPU1tvTy+AOMB3/oZ+l/IeRFAfVlw6SjMSTiqDi875nxj/hItdwjuv
fR7eNIHWuB+oraLaZRTocrNTXz9PLbvJlTG6LuBbakTPncorH34QZr2X+JDTCzsa
d9ch1WFoWNQRYx4RPu5aaabPa0QP6zSRSmPt2ckDQfY+O+tBDn0o3signNF2aBVa
jY3UWCuCgL9ZQHcssNEUZStzCCQh7tUH6Ly+f/LTaV5d6uc3gXfbm4f/ExsHyIIF
XCm9+Vr58hsDKkjFaKoyCUoW6beXcjuqCvIcnQeLQLueVX/X+d8k3Q4sAqMR2s73
+mK7zz9Xn8WfY9i7H9NwEATD5BpSepG7e+qhLCQOGaF1ve+IdsDIAnQRjU2+pCys
QJpRdsTzHAzxH0KiBQY9M099e52IWi2dgJ9qGCW0SS8hvxZ9TtyrB2SrSKu8WN3R
OU/cE+NmNKJ7tjLWwLzRoDZRa/MsUUoiYK0056fFYJB3oBVxFNyDMut3/LGGDQfH
7wABjQKpEDsQHFW92de5eYOdycnrA0RLXibHh8gccPXVBIG38ud+Sa0B9RsbTaNk
tPjtZnNzdFvUIYtichxkJFZRiMtGVqGbUpK6p3VpxVZm3za+A06Jzcbw0ApQPOqx
+lwgOrUFLebKfzOr28YtYca0sHAXiXnAHBXHpSFQFtzFYNqKOMTjybDyY83sl3OW
XCnXEVTIX16IpIxUFdQKaEq/oNDXvcezPUOERi/+9U/mKbHJT8audHr9mmaCdYnM
b9JMDxCO8QIMed+OHrGwGCSFYsA59PZ9w8QvXUvWGSz2AI/FbDAgp+OlNSmLOeNR
P1Hp20mq7g6NBP0azAtJdycaUlHAnO6dXgOgSaXXJtIXomhU3AduoMDxywqUmhdF
+mweiuKzWoBO/keYNy3WAszenCnkBIrN9nPDiDpA4WO7kOnXPc3UN9jZe1GDfC+t
k/HqnYBpeR3h7uWrBYvRLkkd4ObskfOVzzv4CrwVy9vhmcnV4YxYZYEWZS/CvGI1
kv7ZciS5J9oADsh8a+wF/3ewZyOa3hyvfgIGC7vfR1v+wkK9OwAyq5upfh0wtijO
bkTDl0uLD8ZFdTfo+4/L/8ghDcENZssQl9cqTmqOCRipLmLl3ffLRzXiUr+PF8Cd
c4EpsZZcCcvhz/k7oePQMRRmssJXILjzqrUb4irNxFvl4gKyY271CSCXRzhZJZxv
5FFMNGngWVGScjFhRA7vBf+Q/hzlheqKfm5bxwYjJ1WwggFZeZG/Rdb9Em3ihY2g
R8Xc4REX0INEzQaCx/BGXnnLftdaRBL64indHP+XVQb/pdfYKXQrl0EtZqKcFxAj
McLV9qVSuhkkzU1YZ30t0pL0kagibn3MNY4ZkmmACrIbmOP5CXVH3fPN8ej0emDs
4X9t1AfnyI899izdnN9AT8KrPLU5E1BwdFv4JfOrRE3ihiweWOWJDUiuH/87ESHB
YJ5W6vG4nR5e+6z+QRHDW9+LIWSHlUnnIFtm9j6IfaeMUD9dSmIQNwRx9KQuwmIt
rgHAzlAgjWZ89MyHO1cpT9sH2qxrSqv+ktQGWwAnhUmsMrY4e6bLg+rg9g1AloNm
IHzuQaRMk38W2Akchkw/Mp1dKCOQ5j0HaRxtULWWibPmpGCtR5tI7vu35xMbffUa
YIQnXcPFvYvKibfUC65A0N2yber9hYON4o+Z2XNwQXO7tQrhlScqB6UGXdwp1jvt
xBKwPu6KnKuncXoqQa9lCgHQSA8onpPheQcKbdgfa4pPxzgbT9j1wf61IJ6OwoQO
Io3ZV3iq3crqhh1vO1AT/mp+H363/NMUNqVIx4KVA12s9bv5TnjkSjoBv7vE8I23
W640i9A7HOJjCBGNwOUFdwmTV6nkTbgQWh3BX6lt2T4wrSIvEaLFR5pPq4VJqmT/
fcosOzZ5erv+rbl6bxwmfEP66fVdMUre+5cLdGnzh3HKRaiiRgJ6ygoXtwwelzGc
D4SzGXZ19V5VUUkFnfch8nDTVV7RkpepmBXoQepbIRmReaMI1P2Ud5Gjf9GJatE7
zwxW8lwpfSkW/Ydo2e5LEn7TudhdJP5zytOfmLwHCUpt/WZ651legwF6BU5uTfE3
8A+XDwEb+uL6RfJdjPqO+Ss9XuHGxKxEcDnA7AB28n5TwfNswdFhqYmr494dbC8X
6AlUyDyrDBiYqGsqger/2O6On8rnfVMjxKohvUb9Ih1tTNmB/faCe9qSIiiLx20v
7jUS3rUa3KP/JIp9hf1bkiHBWm2GomgVo4T5A9/GCRnAVBRcxb/CuA9z81ZWaLEC
+woGsu90Rh7ykr5EHkETmsrTh580v9YmBv88Y6grfDiFBITHaWAQOKl5MtvpUoqv
qUVONzuap6yrmuJiSgPlDtHDHqm7pcAZokrsfCYeorIgLD2RxUoG9/oe62lK4ofV
ikzVxlskxFO0TS7lj1dNez1yLOalbPOtSf6cLxzSRYCCmm2syf7cX6MWpRXDsNCz
OlZPLDNeNcGMqzQpwI0PaN5hnF8R/pLRa1FTmsNI4zoUHbtCqwVpuAYttX4FV4wb
rAtf2TbnDAO8ZQ1pVkMPiRk0ckcoqiNOiww8xZCQH9R1SftIghnwutbXZzxYyIGl
ZZriMr7mQZZJEpbwVKQv+zg2OCtzTKwq8ZJr0Qurh13FjhRLecyrA+NfuG/MFP6A
fxZioDY3dAfne621OfKhCHimFBvykziglfDuD2fM4FBJcNHyNWk63+sdAOTiJVO8
hPhwGZA8JTI71JWMi/HvVGpn1QAU0HVEJmllWqzQoblyU1pZ7eCMrWakHB6QRY9f
4QbFFPHbctLObAmgsc44JUQys0Cv027+CTFunmW/b0uFzHf0vwhDgdjMpOaltWJq
wmw3bqe+u2BdRRXuH2UdExwE/xmOerFbeo26X6ZuWvioikcBwnIxZMB+Iu/x4msY
LIsCnce6Zeu6waWELfPJf1wsH0jas015Fnz3s2h3SSHMiliS01IbofJMuKP/svfw
896brTHvRYsD9EV5gxHN/Ab7xDD5O96DqSudiOruH9Q+FkV2g1wDmeLWWDqtFt7x
RWnJH8nz2Ixd42TgIhqccziPh+fWxbiBo7ysqulnRZ5SeejH+k5QQbJinniMxHkl
m+NqgkHO/zGfjA1yuXi9maKm08Fjml1FMRXnsPgotnNmPELENSahsjgXX7HsQBHO
nEbmamHkV2/lRJEvpsMDRC6pbEofBbxrGttqF5N9ZPQ/0/8jFt2uFgV8VSXYom4t
azZzcFahntR/fdPl+oDJCZzz7dKkS7rCuxVYR2Vs7duLGSqOvypypb/MpDgrtP9r
IkDqgS2rcdqZ0S0Nc2vLruowx+MMUOE5iGr/TICdlGLWgtDJyiv4nRBjOTsRRXay
JyGhOnb4mFDWVFGHIGVlbSnKdjhhVTrFyBJW3NrbMzKRqlq4oQY8MVy0YTafNInN
nLODV0ynergGzHTjhjxmJ7ICqFqrwoXm5TDHW7HkoeMN8TmMq+2bNgPPSkf4unwv
vYyUIf2VVryRe8i2oOMUInFNxj+2tvA708d1mJZP9DYFwuplNvRXsT61JUIxV4Gt
DpwLv+F/jKwZc4c/hU1kTviLbvP2h02OXRK/qG1I2/krxSRQNNIlQPssz/kH76ki
UWbdGp/nYhaRobgK9MsIkFxJVxqPjA05GgfvfG2X8okfy4a7AtA0HiJDDkYbvV0l
pUEWk4EzQGdkviQSey5W7Ednge03ocwbnAvMvryOQRb1Ow6MdxAl6/F4qCv04EZV
BLDLynLqfqD2Sd5UaAh+QyRwTosZ9nPaVH6f4OMGqA4Xe/b3ZKnCXWmWVzabnyPF
Qbs/DHBoE131rozRuAqRCqv0k3evmlSvFvgEjGfGuiBKLKfk8aE/Y8WcqkQKRP1q
h9Dr8re19RYamzrzgc4shaXS7q8c+wwwy40gsgwBg/impHSqFvxkBGH9qjmWi13w
fHHldEuXHaq8kx2QpaadNh2zbbhSGEjLezSKDQtpLZKY5KMXAcKBbxdeJOGodll2
1eH9y1FGB9/21HdbYuedlUUjnkD2xTNyuX8FeXz1TSOkIr+53DsYeGG7QjztInxs
TouR/QykPahb/GVKB03WTHTBNg7D3QufC29RQBVjb1gRRYxaW7fDiBK14sQ9BIQ9
qIoX45EKg2v5zOTuPm+NUfwPdf4/O2EGj2F7UfEmsY+uXNsSMXkyRPEsQ2nNjV6A
lmU+lYNHyraopYiAm2cqYCTR+vhQtrcWrV4JoU/gfATOzJnjRMwtamoh5ybDRT/j
MY6ItfjPsTPfD1/zUKoNGiJLJXyFX6vTqCcpakfsR+veW9EqORoeJAmC5evUqin7
N8ypRFMeMUflCfso98dzWN/1JUfk8CpUh8q44jAiWHgoSCiYc6SSZpnNfYAZ21qs
facVnUVZRw22RGl8VwSmJ188ggQKpTSMtbwwd09sjCJ+v/mImEYBIf7T/9Iv8AFJ
mqlzUsifcYUrsplRLxXN2NpxF2BCZf9XsOzky3Ken++tEj9xPOMaX70fqp/NXwxZ
WHi017lqUtB2Mu1skW/fwAeU3F6LVvD8/Ecg9qjnIOrYv+7/wJGvCgfXYc59dIyF
8oms4Wz0TN5pDyknch1tJMo8Mjzh5WAG9RoFr+5lnwCJhipZexzAgXgkLmIgWUFZ
2HJljQCvVu/n4BpqFwbq+pAUyBS5/3WsX8mN3PvmttPHzwq3/SFwkwpBSNlm/BW3
Ma+D/F5GnSdT+IeenaRQa/1jxmnwnfyBREaXR6AObCFJhWWlD8mBKw6iKv29mt+O
fAMuVyxisIF58h1163g1tTqbFNzslPVbioXkGP9AnqfPGj9Hh4qq3o9992vcBGb+
4hHEDMUtcV/4QXZBq1PnzyFtkKA8+x8vCcipAdJ2Kw22Jj6VvVJGTr6WnuF5nwtI
EeiQcbRp6e7GCcOwZL4H56wYAig1VW2pyfGHXXc8pSKFIdbmtT+B1aa9sZ9KIh5C
5wk6c/ZKq6gIdI05II8+CgHmbO45U7bqad8sEmSZErYMOIK9J+foWN8LUsmJJ9Zv
Xyad57D6eX/UVNA25zrWIik7KC74VgVsMsapI4VM1qhgRUVhKtsGvYM5hBEZrKjc
ZV38tBk3OdXainYxAS1Oqj10RIpJ/RuHYr3oFZeOkEuaIfn0dKsBpePCgXPlJOdT
in/9DA92k+aH7nVGqKMamqMRqd0s5MCiONg01HB1xRDCCDfJoXLP2R6PaHz+kMBJ
4yfwOIxXQ12cpSVG9TUQKFkUQoLY7lgFtTlNkqE6BTi3aGD1fxq930L630rzbQaW
swX5p2vgVFmfMNWS8Pbb0TaAyKKBHMFliP4gOKoxFh88HYhY83gxsnfI065obSrg
eeuBkopfFsJ+/HhNQACsw6gYKY0MppOvzUxjK0Y+tNaIZQJ28K9SEfFTNELLElQn
F3wjatRLDwP6qZ2p/2hWEvnO7gKsDbNaRLXssmjc3M8FMY7LBYEaVjfb+EFQSOuN
C8NwjdLlsF7ACBHMmB3Gf84WH7o6eo3Q+2DDxPVOd6ufefbSGHsqkwCwNva7yERR
PLbbMAV/J8tniD2ZtIBm7BMkBsTo2IYb4bEpB30RBWSFBxaqtf4ky5KyVINGWtP6
mJ2hb7SOd5/FLZ1E9TFkGnzUiULoRa8xZhhWfoyXBMt96MZT+/AuYtaK7DZBy8ID
77vOGJmeVLfkASSpGCyTPgXKWQqAFpycVsdfXXyPkOunNRJIgtikJ5QBWXMLQKZK
8WcFJ/eKCP37knYLCR2/Apvap7klu4+4YQeLAGGYO5dTQCaxKyQSZq9F2LgiSLbV
u9dPYBTHLxBr5q6rSTd6G4QcvDyJcZWJcoyN9aDi2upq/QA7bSOPAlzpyIgyk8/u
73ziMWgtoLZaThK1o/VqmqqQZNFcJBcVYGwiUZ13FPVIO7Y3cxLHBEMXmG7ax4pf
9nGH3Fqjgv48QcpYgfIKf3DWEQ9xepKuqXZpqj48IfWh3MtFCj8uGu0nrCNUCoxA
JXeMD3xuUr4XlzKdz7Q1anpDTVd+ye4N7PT4qweQNfP9AGlrMntQdm+4uxXFrnrg
dSJzVbH0v/3sunTdtUfcN1/PqN207INL1O0P6AUKTd584RAkXCKdp6/dVtYqdguV
OblvoK115FswZHEFuE6ht3eO4n2njNK0F3C4YGKPYdq6HfO+74uzICKNw3U57VDG
ztZNOfGC9ktxhyK8t8nXrFYy/YuZeOjm5R1iNFORGwuoycymvHHs7dU8UKEc2GS2
nu2ToQoPSItUq4kPM3a91Qko7EPWhQs1mWqBEhQWVoXr8LHrnTW5EmGiqXx/wrNn
ygIB7g1IY5X7KWZx8lhcTkC7oFshnTnYk5pkmZzoMYDbrxnf52LjR8fnR3KvwoAL
JEpPjuaIYmYRN2eIV1/cy3Vr6JceXKb3IVCMNh6y4MIgwZiE2wbfsLQjInsPLi86
WFlT6U6FBvHtoL3inFsWAf6f1eJ0+9wn7jGpHYQ9oSbA28cQXL+/Lm3E7I/Z5VR7
4sWzpfPuHIBNH3OwPAgXtHGaGDB1Eg8EmA0l3Ii3Xeyq0bGDz0s3L6+QdfA58kT2
VC+XXbY9Qaao9sBupClkwiPUZl80pKzL3nkvU8YuilQB3KDK+D/qpsm5IOzvngMd
1CMgLYwd3kbw3MAG7YGm0VBHXNdsnqJ2f9cUaocY4QwOiT9UfWzEq5twVO5kXZF8
aDme6oGvu0OFq8o+0aDt92tVVwTH+kr12st23wJwZ0kO8dqTwPrSB0NRdzGAEmUl
jInmAkyg3sqh4kEUPqLQXZnQjwjVt04NyEBmtzzEeHZYwP4nercqSZahzJs5CLeA
5ZfyRh7ybZN3zKogBt8a6N7C7f2DJKv8JcIH+sJHmRp/HI6WeCu9iGMIuEejy5My
TzZGFCy+WpKiFNLYQCSa3Nj9e3ThJiFzvr3je3AQZqocP3AYNHF8SKwtN6N/px6Z
SgrJLxxzY38+B0D0w+8d4qp4fgCAzKyu3g3QgohFBrMM/mvBy2TcBN2spubBwMBq
om0Dqkzii0Ay1QGM8B0sEnbWod895kspBewIYnGXQEXKIGZRChBV7txILzNvDRsC
7DWg6eWmCqAZdH7tY+4jLAtnw1vuKB3HlaptKXJcLazcfq97ekTLUtNGe/XjG1R3
d4P3k/+8TRydD86EnzbGOffbiVeRlHxsP3tEHX7FRMbeCKEZ/rFZlWaXUFoWGdMN
+whIDLMZ9C426gal5bJDHKsKappjIqB/9cWdi31JfivRgJJ5fgF9q2+YEWDERsuz
wiPTwy3Ogakz5KP9QYr2tFaJh/CeMwhmIrYWpWYps6qZwpAf8+ASSM4TQRUm5itO
nF8hgaIDEBT0XJOU2U2vC6k5bUdLi6LJQPiaPHjGml5UxOgg/w+rOnXPU+I5MDe8
f7dIwtvtVJ7jyrIZrLa3ftUKl51Y1wlXhV7eCtQ6qydBpGjEoXyy8LWOcPL4PS70
Cp9jZCKK6uu7r3uYcDfjy5WSBbXLEdrkP6giG/DrapODyOE0qqYP2pGE8qrrTIn9
uqqw7DHCou+m+tV80H3vHyZ0QSdsNHYO29SUyVQVVmN+S3FA4eYqXwy5Ziu4jNw4
9D9EWFVwzycafTfieE0qVih0owc/B9gxC8tZZwtBEUsIo+N6GkXdjKSB9APfU1mG
yR2WVld5dy8kEMUrsVymTNoELymqg/n4TivPGGgbf13FgHRCu966ff97gTRRhl2H
zU/slSwyKEEEfehhPLbJMCqp7AE4sDdxJNHgh83rJzd9n+IvimxP+gUqiNQhYNN2
ubiSgIgfQfv/QOKbkxETq+TwzyjqPk/pwF85cOyUCJ1Uuyn8IvyQKmJAvLYhNi8w
OW5304mvz6V+JolqQNkrSg+b0J99uJvcGiRoKVcVVw0yfViz+BgX5h59bk6E6jPN
N1rlmR/X/e7RbHwYqI+/HiUuanE9mPf5NlNDBQkfZLZ7asGOs+DuKAO69kaf2qZk
0/m4e6VtlqLyewpHipwKs26S4FC+j+/w1uTYlBvSDsFzjQP89If87J/Hx1N/IFd5
ZN8mgCHqtlxp06e3JWJu6d/IzyxwImJXjP48rgleEWN7bxVtxInbnF9vvAcRU64k
EyRxfGLSImaJYJT0U8jHU/MLQW9h+7iD8ChC/SceRyS06iXe+wfqrFiDsVASGzZX
GcPey/qt253KAmW6+DUPGeFO//O7gXgZ3VLcDZiaEJzJwGqlYiCEPK/ka07lpMvi
4v8TCwC4hdQnJ2wD1d1YOf3L/YV72dgv4zwJd248jygFLDZ8zRtDz9pnJDt/WvcX
+FE1n7yNoNDEVj+orE2DrgGhX8xOlvvEU8u5BTl8IDZS9e5inCHymQzgLnXGUN9Y
LyfW3XB+Hhg6gIadAkpL3Y4wiaDmZBjhryxndvMgTBzJJ3/3w0ulkjxlQrMBzoig
UlWyTfSqDH+rauST1D5djQasL5veuBYh+Hm7Re2cxlO/G1tLHS+hvv8b+jqetpke
P4sZuHjKhVLv5OeDXr8mWTxN8V3H8FJabOzAq4h5mX3433WFYGfLVNI5cqufCsgU
cUvF19zcDvsJaOaCZ8d/l4Mpvn7usfro3qG5+EE0u99XveuXl0dyQ6SpMQxJjdQw
qEibGqBRp5FrAb2JfNO/qoUwHkVCZ0zR4wMNQgtlXmMhiLgRiv+Rli0B16bU4OO6
P6iXHxX3dtpfJDx2ECX1K22FsxUGU4fF94Bj6Hnnv6+HvQfkpPr34rU4cJBy5aSi
TdqGtotLg7KpgQ9Fj9mEONU4LSMKCuQ2SKh86gQ06eEGM5m3VpamkI7cvSOOjK/B
u4M6gzhUCxgXJDsTPiBjDTdJwcgYPHhc08vJpc8tD65ctRCdOijubttX5fbrVj9I
qdgdtVUuL3fmfUJprRt1+/o4oS+GQ8r4+x1EEvGceSInxNmN95+dee1jykLr6cHj
Jkt9ik474Pu5EBmtMWkLLvbxPvtM4BahZSUMuK5EefHWmO7w/yjwuEFrrBo2PIi0
B/8FTUZfppkvqj24RS2Xuxu9BE5GT/jgQ4DyKX6tCj0UeaJ9VAnlwRVZiaNiRx8E
m48dMVuoI+8OTkYxl4r13Gt8MYqtyCCQgYIf9/wQBbw3T+0/LdaHLRmblMfm9G68
Hi43ZKMeF9m3sxYdshl8NAq0ih5BObidfW1XT/f/FGwyeihYvM6u+195Bs98bJlb
IafjDVnflQ6Ed7YWjqyo9SD5KFiE5LKOlUJ1UA4JUSzcbhxhvSjGCzJK+6VnyXsy
optsfhaqfH8iofUwd6CIO3kPA7TS8yTgN0AtD4VdQ0vmZCDbga4P6Z0gLd9x6+dC
s/AYsHMpRF/TGxd3Lg2h5SOfADg23l0Z9+w9gLPp4yN6/6OHYG2cxGHqSZFu6SXF
g+K+vFX8usd2Uti/acmfbHZOMk0e41ZS5KG/6u7Rnx1Jm9G2aWU52VG9Wwwo0sc8
AiClGytR+DsXVADEckOK9O7clfwhaad0gaCEE3BgCtl+GVUoqRbQ+dgJI4oGtF44
tgl2d8hjy/TNwsQWI/vRZE5xSIhvceina1eM98imeQI4KUuwTBK9Tn43uZal/+JD
qpagFT5TI/rj3zgWX1NC0GoHa8S4+Evdel0mUAiLTOcI6yi7Cf6/lZJml79VCz/X
Ze69INQxScvZGu7oPgGn9pIheYLB0bVKbVqxQfUKx8lAIVGLy6Ol8GrfX0w5xGAW
xLKOkwRnewrSadpq8qTbT2YBFEE6uBldk3Lg4o98EmazG1jIPrZBDYTXaF00tKmC
Oz2M7bpinbykSlbGyFz9NhXrN7oL5TCI9r893ffEzPCvEjuG4niBOl2M0m4X+LO5
fCRRW0IsGW4oeIB6y6wMgciOxb8dRxh47RiGtKGFp637S6nDQICScvXorNx/pH/F
uhmPDPMf2oPBPZGVAeKNX4V51ynFVwtitAhU1smhN2c3lLnnjCbACQ79HhpjGNZk
kAS3lkwyQwXMRwKXdemcCDMhixyhCO6PJaz27Zlm+IgSg1mc+WxnITeEynnHehJQ
cmHeBTiq27OYs/eavqZa3nqlGfPaOZGDoUWtfWWhPON8EO7hlw3/tltFHOYsa50j
7JNuGe+fa6/Mw0CHp+t1Au5VWynaSdtwCaW8vF1rbvQRhZgeQeYFioxLTn1sGYwA
E6r/14MNTUuLjdNA1l2F6UXkemvSUu51S1LeBEm5bLDvhi5IZ0TQo1CHvtci5+ts
tFPz1CSQHJhee5zvHQKlLVJKqbGo2AkYvO3yDt8+Ey4Uz4BsPbd24oyGOCeONBJi
v+dvzfOkHr3XsydrMcL5QHxzXXbJ30EcDTV3VpsT69iffHYga6QHHN55klWgTaar
b4oWrzYVJJh26+t7Wb780N95jYDrp6KYLLBYPIEvky4OwQ7uMb2mhPv5FvCRH7Bn
OfcBeAHBraQVeqHfxZbparuIdc3YICmoWXCY1d8UhiIiHmyyHrqcNi4jh/zdsHpg
7qWgjXlbnCXEqKS1igTevMvZn6yxSZMcrcgkunZmOirLQVPmbmJPNxaaCzKAlrsz
JUDm7snsER2HdCqifdsXlS0ieyRz12BI5iTn4XRa43NyMe23icFnlLoJxnD4hEnb
/8JCQpRDXHWW8jzdPEnsCf1nokmgpkpcNxael2aEBFQzO9V0zjGj6HWYWRSXRNxd
v+bVvMh6l6sMC1otbUCilJgDXGWb9ZTQ9zc5Zk4XpBnqFElG+VJLRXBchNcfms5E
ZSPs9UrUBXyDWK9+n8kMNbN5vQa4KHGNYXJJOHU7CFS4J+Y0Nl9LWLpL3aJFrIy/
Wc8EBCYnk8npswG5mM5bp1FdwGFqX9g0t1fKpGLNJhfIYt1BhjvRef2KaCbp7VUW
BkgZmodq6uqzC9kB2XSTjuOl0P2Vu9ObkUlcX6cz+BRfgC9jTuYZ240PJCNPCVuB
EPyIZheH4qFmSnFfuHxJtCOJ5xBW+82l2vk4gdInRf5XWIEY56VFrRTfsNgXBpLl
9ttf4L9Ru1b3dTn+CqCSITs6/BBplNTsPM8TKspRQFBnJiC/pgQy3Utmbu6sGtCq
HY0hI9/a2H6oz/c+/p1hnDNq4hs1CXTDQHm2P/apGiHZc10lYyOXKuZD2Iuphlta
xaGvbAc5cqrE/oWaTBKpUuiJUnv+yTYRpKQPZ2ZkLKycl/pMEaH58CcSkoLol+bF
K6NFsHT8RtnHFdw+Pc5GgVK3ThhXM03Sn/S42DEVqs3ulcFGuNij6z+LiTQ9SLzG
GaxZpYVV3NpUh3QiEJDcllISt8Iui/VOO6OGjvc9HnssxeOWs7Cm6UnJKkqidOXG
jZ5PH6OrM58GiOG407vf8ZavMAAhnrILE7Gi7AOx8XzV/NTqSkRGJoT6+syZL8Kx
D5JsHlph8bSG6Wsm+jOmJ87+oENRS6eVqHeyTP8gHoRn4K2JsFjDAg9N902Am1nb
4rhmFJkGv+y2uy1JbLizqOwX4Bq+xFOx53ZygiuW13DC7Ss1N7xG2F1Fi3lF27bE
FEy97tZuYnBJMB538Ivo4AmEUNt8M46ymO3cCOiRsNM290cFKrrAYMzWykZPPQnw
VbkjXCQxk7gNDi6ZuqUa3mDjGIZAnUFZN3/mvFkuVHwkm6RH8ua3UcBUyxKv88nB
EbyR1YGuJyg7jqcWAe0FBU3JhRdaDIThJhf6HAednc2489jy/VmxiQtBPdGegCRN
V+ilccP00b/zTf5CMQqONUOUqiGKbP1ZjYFzOyI8+DHUN7ir+sYTHPntUmrETwnk
EZCl5BFfxHokEQT7IIkLmhT6KTAiM2DMvZX2rRFKyH28KAIDkjPv9wpMjiJAssd7
dSpa2qMWco+r2GLfz9P2VRfQTqlCCeiMq6C7GMQRpcq+baJq/OEtrYCvATQWi4gr
OMtipRUuZRN4U7uXpZ+WtI4Hp8yPARCT1MJUT6HMqpcKdXN9DpDjUkRpu7d+DlBN
DJOIxpJbauS6YvHp4yivop1aQOAmrLLMXaUvbtxntn6Goh/3iDH9DR1xp/jlqplq
TfTV1jIKTe85EPAHGAiQ+bmlq7JQ3s+ft1aftJ8iECZhRqmgw5mi9G/ykzXqjazD
Nq5R2qTxZARx8b0HD1s7DhBc/fR2huSbzPgA3xt79W7wIC9+rdodY2515moa3jHS
x13uMe/wc4EwrLFFYcb7moTqEcd7LutsVBbXKgyEW3F5TsvGX2Bq6MkNcLEAdVwp
HEbP7qMtaeanApA4X/eIWG5zmN8U0iWSqWBdODKtREcV7rHwUtJQccHDRKYnxLhv
i8JgqeIAdP1iqQl3bqTVf0nlu/KltiZHwr+xyO9Qj5qlfuG3gUJjugN8W7VC3I1w
z9bRcsMsQtCDez70yp7G4v4k1wmD8YYKs8E2l/WdCxqbUDaFtE0rvEmhmgRpcIjE
/0uSAfnStEHyX/DuuVKPue657wARCxexegKxsbkv4R6T/xJv5IMChD0GaRKNjXWH
ijdXsUCR8klrm1F48oHIqvDRmFUwNgrER6FPginaa6bjoApXF640Z2DTnFqDqqII
dJxnmfKmfgrApd1HZ0xRxtOlTqG7duXj+67VN/1e+2LWW1TZ8fXByQn0wvcAnSM9
/ygZ8NR0mApe/jJACgvzqGHih6T0Kid/PCBf4FC6Cq++IthER1y6ecAYtsC9fr/i
mJHVtQ0P4QWVx/iyAkzagaWFUPrDG3p6s6y0s4wZWukQNYpIVZLsu1z9Vo/++K/N
CGAJ2VuYKO8DvZC6MMOACMB43WnNx8TS1qO6s+gCT+tn7G58djCkHbo9snQdSR1J
mF9uHlX8eg3erdl9e7eAut6xlOMxTPM3ytla/VAqzCp/A/P5f+4vu5/03zUX2X9z
IRCQVk6Z4u2k+BYkTTxawFklryid02CGk6ySc3K4PCTDH6Fk5tCkcfsovBnjOpJW
vxhR/5ISakdaxQ/pHn5++UaL2EP7OxtB6ZbMMBr+Pu2D3NI8y6GvgOlVam5dRhNS
2GRYCFxC296llXUn68rl37/LVwoQWfnudsGi3dplFzqaC0Uqla4L7Ae6AOh6lbRZ
P1HagxZaMlIzceA2x7VCKUEoLAkjpip68lHYxNXX/xOjzamMm1KUHuBn01kR2wjf
COSnCJ58yZ4P5fs1K+aAAs97qFvl1UcjBu5Ix47ZfuHyEsr8llBriSL9DfO2p6RC
6FA62LEEl/rFTlv9187D2xUUOyIH9INUVLjme6BwbxzrNkhtwzMjCKPoOMDvA0ev
ACF3ewqL0wbJJYsXy2omrkjQAQfp2jA0iodKcLFQZsWUmv6oeoiS2U5s91wK9GOa
uvnU0DVSSYk/DX5va5HSD005QsfTb8IvUfdTnbsmJ4glSZ36FmIjAOcwNTgZ2SpM
CfyNMWgy/WWTTi8gAO9u5qox9D4djeN+8eaC9TA3khiRQ5WgoLsxncGRiyYULIr5
lJKjKf3J5Dqw/CRB3npYm4u5AWeC0oGX6NVi0v5gJHSzr8GxA4ITgJYNUuWAlR/L
+ZU77lS5rAgUFc43VxsDfskLL6MpIvcp1k+RBfhIeLIShEP/gkIp2XpOPh+dqSZM
8+PbGvqoTPUTmw3z9uZZp8N1txchNe7Kfcsz+O/fpIr5q0NqSRKHkY9Ejd/jagK2
t9HXHY7/ARpYyqD9jFFs3Hve9aULLIGKd1WLWlUhfmA7jXFOpueYqJziPyr7l0jU
f9+2PqlTRQys5PqnG64XpLcfs0zjXBM6+mHeu3xryYECi/Yy5qFUcjt6iQMRDeky
Q8dAdRw+ZdeBq/keuxX8gGxJbjzIdF2/7yvHwinzOhrQmQa2TOcy8onZotb1FE2b
RYgBjuQgptETsz3tBjzqR/qdM1tl6DLTyYdggiAaE3uJQxerWrmJD3e+pLv4CTf3
bKFW1/o02nzwt9xYaKL03aeDRyuyrO91oRtOJW1mABiaHMm3+1qtRg0qwF8qYG+w
H6Qa8ekNN9P/V4gQPcuW4fVCT2TqYOyorX9x4NZ2L+3gTL+OPLwGSkN7rYQeae0K
2ikwR9wzgP7CWSRHu8OqaFoG131U5kv0aCBCS/QkOoZmxEKbeYlIFfpzOSW49z49
2e4YxJnTJ9zAZfpSev4RYRF5thzXcIs801LGgPUpirHmSfRg2K29dqa8Lp0tPdVV
2LGXgVzEDeleZAYIchCTsHw4pX27MlpkNKX3kKz5aPU6p3r52Itxak0NwHDAqOS8
G8XvBPE4J3qgZROIGLtDv+OJGdqL0gJFD/9JytxKD7R3lPNeJBF9SoQBbgzYWRl9
6IoABrYzXjwb5+QripAqWeSKggPjKgow3HvB+xXTD0zajadd0wGHFfVNg2aqQxPj
+fvzSLEpNqXbcN7vTKb1mOyzo4CuZRimgeukGKbS6bFA0GB+C/AkyHXBDpe2qu+l
LuZXxQK4eZv5n3rGTk8uzyIu4/X3kK3pTbZbw+7YESqjoI7scJwaniqjq8sTPGx5
mmCWsrJA29qwndu62RGKfV10NEvbQbD2/ZBcqw1CCpTpdy2XVNViAIQn/CJ8lFWc
tJAs6caVq+KYODGkcfHdEJ/r7I8qS1BeupjY03N9jJYa6JxR6P83pPgrnhn/L0hC
Bxq5D8pmwesoupF+Q293ZVjF6iMzJ3SnQTwh+cjPmRe83A43LQXI6cNP4zUKxuDO
yGqW6ae6TxRzl9WMrkn7hnRdKi3B4w34QqEAAMXffxzBvDHIME8r6PGA8tNCDmMx
K49HTXXsjXRNPSgQP59bJcN2woSwSqvaFGhHEWqr2ha7KrsrZVRnhZikUaeFgH8n
d3U8fLV6jp751cfK21V8HrAKA1CrouIgULlKlT7E+2+lTfRq842iupXHS1c3aen3
/50noMEYt7Z3BspYtvXY9ha2+7Dd6Y2mndex3x3FGv1cnWS0ApJaLOJ59NhJ7Jza
h4GX6J4+X7VbK3AHDbZA+fu/pI0bJ/AhmQMO/ECiyDaweNtwRtsaIyxH/pitYz0q
YdLXqAeiITIlLIyxb7hm7SVg5212Dn5HL4dF3mBSUgi/GbI4six64jGooJtayeif
VdIfgWX7MQKRp1FnxHadFKwvIEeRHHrlf21I48rtc0ZganjsopVgEyyusxh6P69c
nWoMtVCFbl9QdytV9q1hp6nmuOxfO81oYvKP3Ym1mbHYphnAeP+51wmqHP9q8FTu
BlqsTpl8ZQvTXrCy2FNQg3Y1GWTH2GtcDrae/M2wFGw7X1+ewZllqnDSZiQF2ha6
rpn8EJGvhRLwN5UGqIfqruSyLj1yK5kHlrEG5vYss3MZjY/QhDJ36uaLQSLaxO3s
Ww6J0DxNZE75Q7AJ2haJ0MnAhzu0zhpe127NJ5keA9Mf4eXCkLuAdTwGbnP8NmWn
vQo8VG43Ny3BKANGL7C2e1kQtdDOhPwTw5xQql9JXhyxvRFAIdf1YKZbrYT4zkpW
tyFIqFQFqGyf30SSc688E8s4xQbhydfo/VoVpwGqwVKM/Q2C78mu5xFSsVpSMCM9
G+GH/jEVlVsk5avyBGT9aOOsBilzs7PajRLem4s6gxECH//QYmxC/Y6FyNqmvQPA
du4jL15k+Rl9wDi6eyP3gPY13khuw5OGe28xg4BoXW2iZO6HnvwrfEOYdMwjg/n/
7LFkjh2ZoeYupnwZZDclMj5i7IOpRDhQ2U61789EaLGomcUE+6OZpY3hfJWGOn44
c1CEYJY28qNwd5o5cptHC22IcLwHCGNLofDbwsLAaiDEkpGtVI6uvV1HIcFCVTpw
S/w+/LVjedFmsPpwcXs+ldCK2TRC/i5nyGvCvegbPWzsLU3CX388DFDArJCLu99S
1Ay5S7yW0h8zSt3/oCisqpXpLid0rOmDncOVLhgu7kyHT7gok2k50OBGcky300g5
igAjF7McK6ezXIeokzapJg7q2lWVsQfQWwhYPZEBWx1WCIZEE2WRnaO6II+sycgf
ttTc1bySyIEbT1L3ds3EWSce70Yo5rkPTQ9cszFm2By5c0FVpoC3UYAdHhORfJuO
Hu/+QdTvO8Aeh7iIMCr7FiZkrqLERY9LgEV2EoBqRe2daq47RgbInwiReMHMWa/i
MMYfA6fRYFJeW1dO5GQ1pVlSqxxYgILexBpDgt3jbEKy+efDbRMgu4QZ1/2fbq3V
//pICdOOEs2H1HLXv1dk70JMLkgaCsZn5UclPygamtfJH5+RKN9XovKbSFUVXRBN
nrRIz4P3CYGIldccHscI972J9f54n3zAx9PgOh7g0dIcpmFX6wnkARpohYOdHM1V
mdnesaa5PvuC3hbUP8tzyY/UDmoml7O3v6mM4KmJMH3wjlcwilsb5NfOGNzoA8Zr
Kpcly973JifnlwaH8eHSe8GB+5JmBvRekYD6GDpA3SwbeOhtsu8kmzkSnCCnh0ZR
3f6ddslx5MwBpyctsuKOo60wqp6Knyp42/rj0F6HCL0GEfGZ3sW6UhPyME+nnHTy
rL8J+zD/JXMvrzucc3Q80v5UYGxRjNIJof1UqaMJ56E4IkqlXnhPJ28xPsueR4iw
sDKrgrs0vOIaxBTr1Vv8tvrwW0ayIJIEbz4hs4fWCg2QmJ1ofsyC0hZGRPCJxyWt
VrRgIUINH9mSckmpqgvVXtX+zUyg0S2nOIjFHQozGAQtuixjc7skDdhfQPHOHMVN
xhhIdibl/Rg9lOiNeB6qFmpfwBpjaZRm6kGXSpTPd3jep0BQOXCJd6DXa5Mhtfi6
gC5ZSAhRAzylLZKbWlCHZaam5DQ6Q9JUtSu3HjF5fgMCvi1EArQRevZVBuY9rb49
vITyg0+bs39dN9+m1Si1i0KWWGqbp+NF4LiN7YXNvXTbdJJhUrhFhEUiy9ftQUjx
/OUyjeO8Opt+uL38PK4SzqNEehKZab0dIpxkAiJ5hAuDXUtb9qD5E80FcTGmZ+o0
ErV7q4oedDfH6Ct+FijfONbUJuyTjqPA6OHqcr11ciz7yuzEKjF09JPb5N+VfyVn
DlGvgw/L3+b8fMqhEl0dWCtyAi7FgAcRTpttF4KyyMv9lt+BB7LZOwGJ1qw86OLU
8n1VBmJm18MTGB0lzTRHfcfvMqpm07TM1EEzKnFyc8/2ZlMrhcqQEIYc4InhclXX
8atluQTuLs4FEYKHhBOBV2ifjxE9bxn7qfuD1i2L932VhpTV8j9tsAOjiknLJzEJ
ibpdipjqqiIQN6k3x+K9WVfeV08UukM6T8js/wI9gIEfqS5xppVezNsy0XSy5+lf
F32m7uyEc/ZknkQlGa9S3P1viuei3w0J4oHYg+FCV+xBfkNCM1kg0gOTpIakz1Rx
KtBp/AwIXCp+c6RzkzcGfTrTOS21GFVies2scLzf9AJL9oX/TFerDKgkNoYWvD2C
qMzYbldrlrMg0KWiTiBrjkt/2SXbqVubygmSnHUURsud/NyBKyYcCeuA3ITw4ono
fwOA7BnnQrClXqCB7pTNv158ManwPNH+pR8+3MY6w+SKsW80gov9H079g9CZ9Xeu
nYzgxAj/ygstY1kYYwGS9q/mjzhg62Iiw4i/g2dQOBKVL7bJeivtS8/BX9aXurs9
wRw77Ih8xWRZMrWohYfIp8U1rqic6KvHKr9v3HoW1mY3auaaENRg6EF+iINVJhMl
m/Ix2/3GA8bQHmS/zEKNROeCUdHlAm0t8cCgNSpcoFt/gIgBISFqCQ8k8I7x9RLt
CUhH4ZddYQXpW/5tkjxz/Df2wPX3jiNe6B+xahe01TnVvBPAji3UgdNmQ5aLxuQ8
o54DpxE5HbFgUeBXVBH9EZLaAMQuckhsPauf3/OGTMOltmFIv9y8wAUWGODzAS/4
eTjVGR9vRPjx3QL55zaLSbl3I66XGaiyetcdqVMotTvzDmGjZXeugzIAmJXdkFti
ERNwv3+MtJZmNFOlYn1JJIF45ElW2DJWSgSSDTNno/LaelrIR5Tz5bKIBN7UDMP4
8MHSe9mgfkt+3wcH+uIFXrtHw42xg7y8VzNeL8NK7VvVtwt71wZhgisnZEjRiyZq
sAVgnC9YX4Exxt8948o5k7ycrN3RMa6fO+Kubkypqt/CYqtAUBd/7t1E3RHSFVcH
aqQhue3rvO4eOiTIfGVCKDMbW+dZXTMDF78/dkLIt5kvs4Mw/WG2aX88OJzILsTi
rce+C5SmDmAYcAdXyJV+FwTsue2SDWGBO72cNcpp5DsM5WmkssToSBCMK/QeQPel
Ie3kkPLDRuaH2GqPFbCuVoqAsmXtOfjXqd+eMvTsHxDMxw/8DYCfrx7rXQ3Mj7jr
HpR9lSXgX+eJXCd17ToOU/hIsIDNayFV8ol3z6H3RPg3HN22lISn4mSMM/x8fho4
plyFk/Vx5dicNJ2kKASpHZqelDAEKMM+eI5xj306CU2FBFKLejnYuvJL23HbBF7k
Yx5F9/AR6iewqV3etER0/aIhykiB64pxF6wLfiE77WGrEJpuaGXz9DDTqUUGdedd
Urn0EhBUis9tRuzPnDxC7TVd9EI/Z2TVOJfGUMl6YF6x5vmudibNEfxQq3EtkAYf
IKNyF+PA+JZpZ1GWkfNHaR6QK8scr082nv6iSqc/il/somT3s1mhH1xIxv0hgoIi
lxd2JbU40/WObGgH1ZgilFnlEKXqK2utv9XmKN4FoYQurOtWxMJ4XlOa7kYRAXCz
JKO+ml4863hL3b5Uo3cmmlbLhoaHl1aXhGE1wjL74V7cLiemlU1DJeP3Zi/ME/Kz
hYYkyLlKjKqdYAjUU3xbDXa7oQ4zjDd+uOJilgehwN1nZSmV/AJraKu0oz4PHaaW
WIhnJpxC66HyJjXmLKvrB9RsiIgEPoxgXaRPjtlhFlO9qhssDyWZxk3TU7m5JGKj
wtcsUNPt4GKcerc9cmV9jjRcAMARdXCn8dbcZK4qUyjvzqogU/TImooQeFeVUEQc
FIJXwUpp2P0wfUQ5O4y5ziPHFCEU0IZYDF8dPmn9U0aIV/2wBCxH1U8ZNsns8Prz
3HgXgRQgFtpOtrnhiPz/0xbFGgCC7jLNQdDd4fAGxfLMyPkWALnXsY9mSlLFgojM
P35puMO4i0Gs6gRKinaMi8+Mx+m+MCHe+bj/xReTxxpal6hDjhfGuxBZZpuVIwMW
rjk8dP+dXPYnq258OSQflD7KmfTr508/AyZjt/AnvZSlByK+JeG/7W/0cQ8/XSyl
SnGwdkMHJEdX7853YmEBrZsnyZ0IR2IvNX8ARultepiqWEv2AQyGzMt0W7fGpcnY
c0/qYwZyL95kGQYUlS+mUZOsJr/a3Pjfa0VKi0NNnpYQHZwdUJedVGgNvjLHqXH1
LC5T7K13QHQV5QZHOqfZrYPvsNcUV2RjnlqlVW7cB5upSg7/tj4prsJU1xCydHc7
j8zg2CQurviTHmsKKLQvqtLUp/gmKxrLggVyyoVjK6TnHCUe7e5LZNeimX4PHdAa
eirgTJMGEvdcNAH0SlkiNaTF/C6LPeITS4Ng6TN3SkPVixOisB/+H+BpJVDkcYe3
azb7T1wUCbV5o6ylM44ufsb38SAuUgnArCNwvOc40d50G7HCbofWl75a5wUk6B0i
u0QV7XPZQDqwZcNHoJYy2wAaqYKVosmFXiIfON4DV93iVR2lGsyK0xGYcQG5nk5r
Nqj56K0XAik7W7IG5dVY8Sye3WNIPaSnkSCfHQpSnzTE35zLUp9S89qjbXRUket2
G9OXQG6mAkZsvn8pb0cgR91++Pr9spwEtXLfS5HOHZiXAE7CXqHkd0sfDwOaYN8S
QzSo+0ZIvT8VGQQbPnFmu1RK7dh/PFCcjYHIh9hs42gSwCa6o6HHt4SIt0DY3wC4
/txVQZPRXE1+6sHDLqW7fDkd+Fc9MRYANR+kmmyUL9oQNdysZ09yboH1SfKW6Rqb
jIonHXoZN/iREPEbvvZiXTDdCrpPsozMQR5tvHprn6cCcZ9jpwmUtsJfHT47xwJ5
aTKLZ6uAwHMmEDKE4ihMZNFqm5ebpxUfJfF0/BGZBzCfFAoZp8QPfcsKFUVGVHJd
a6VTH3i9t0581HAtpaRGze5ux8RwZAXYB3jKFuQCDcW3tJT4W7CLr1UW17pG051V
dZTFnUQw5P5tRQqE4HSKj2NbahMDYECQaAJko3MhFHv9HmbMmhT5kLsyIGU8ASY/
7D0h/EqnWyFLVipMYVRqfP//QrWv9KaIVRGDEOe3ntjFqS3ziHarWnKWRghCNwK5
LCbQ1LlMsatn9OR3J1188lxmisquuNVMnEhF+/RJqHzA70aJwgLaLXD5NW2P5QwN
yelIsS+8dAQ/e9VLsQVi6GB0U0BANG9aGXu3WvtOvNlOtstUELNPXJzd1SzbOdfm
Vy22XWhN1DkRYAVrJREToJeBaqpgX/L7KDgcNn8fo5RSsKPF6ShOII1v7PfntsG/
IP/1gM0yXasNPn10Oy6ngxNJhb3jlNlDgzQwdbxVyXkTVsjWGbzW4BOrB39g3fEA
HCzNq2y19YIZF08JYq+VNdBjFoJHcPcwOz4iPe1s7uFPnVpzBskFF1loC0xRHNgm
k+O89E/GwiePfeCkJPAJ9SAnJMwH6/gsoYmc/RoOveewBRDLud/WgKGIYOg42Yhv
FQF/yIhW3E4QiiZOiEJly3iVra/ZYDQs6UydKTq7x55zksL6JKf1kv+tZ5tWWx2R
unGhfMGZbA6uP+no5j5fyvfeQpOTrPZsNSTzP16SlPUjP838iJB79Ox0Zx0jWBM1
w+wkWGryh0z2jBLHHGk70Uo0zc/qhx5aN3+tcKQVoYBs6SLp38YCky6+8ESglOhz
OWGsd8rKJ0naQXirurQaoZT0FDxlGPkImYepZrzH5BukY6EpiMqAy/JOtyaa/h06
WrAVbdIAhlcpKIhPCdAiGsfDBSNZ0USA53YhEox9SShT/DeBbD/DTDsn5YYO3A3j
UM4DDJBvHKIo8bveSfRiBm4TXMrXf/xHHKuIpgcE6249KREM860R6iMLXNGLS3pd
gGB7BiujFEEc8Xufv32rapauuzVKn3O88CP7KrAHlgkHD5lPohR5nJElGO602DDL
ZnPP4O9idBoRnPS3QD2iWSzbn7v/OTEOwAiGyDSUWqa6a7Bjt7gHb10fDIRp5edL
bgYruYZo98XbPAhBTn+Rtw/M3U44GfFwSw5VmqKqX2gd7VdNLxnHnD4KWK3PSLaL
DlKFlCSdaKHa9rIQV5SiztkrU1MROoCz+HeM7gFGFFZ5mFoMoAXC5WNqWyw3bOyx
b2NdomC4w4YIrhyVALumaU0mPHE5ngGfZSGmQ5D9r6MPCw4uBz2w6a2ClaQETeVN
8XU/BQp03oQeVmUDTlEqf1epGMdmPin8simrFqQdFNo60kLb7rmN/s+zGeMAP/BO
H+VJxwPZrtWB7j9EoYAw48ewMWuRwQvB1zzoyzSRY8YZzzvmYePMBKndgozFk0wV
5Z/bhdnxo7ZgVyB3/NSHgqb4KPb2CYjW9Mhmr9iXraMSZcsnT5CjTaSTgnLFXLJ+
SrpDcTmxFhDrG2yTO+qWWsxn5YqOxyBXBwAyc71KWWSZ/rLX1iexMq5UesnDGuRD
ngwv0n3YkLxD7UgSoZwHfL/HK9KbleG8Oxdca9E8W/X9Qst7J9NvPAPUoXrVZB93
jf/Vbm/7ce5XiWmQt9hYiUMylq2EjDKoWXfr0qO+AyHkq+3rLXSRG1hY73JXrre1
OOj188vUWRp3Oy+hWJdC7DC3qqTUsVGPNCAGFF0L0hp/kjQjIEqFIsbm05b2w7xu
ZlECBo1U+Md2enQrQcpdUe0ZTZY4jdPzkEceQxUO0S0fxKsBZ9mb2Mf76UOP4IwH
kdh8ADxZnWmSBQrzb/ZCq5Bt0N0OOsbptd+MN9m4lpFzJ/l+sTC6EBbhdY31eSfA
9yoIVpPZditbmIP6X0GXcBEdYn90iDJNApxm66M8QyiSbDHVqNlj2ghCSDiYQKNG
zlts7+U8kxM9Qhf5niQaIdYUcc0E7nJQO0lTKRpUT4BYcPFzrxynx9WQVRNxp5t0
BthzEQhHWAMO2Hj7bBNI8mQT9osIaX48wvTs1SEGrjgxtB2363FXw2oEdAJyY9wL
SRK1YDjw+/ZDl3jmeKrf+KTFc97xUqfxo/3eDIvy7Eb5XNPj2l3Dxp0uyNHBqZR8
8da5O8HOlgb0aUOMOUo+Gvh1XJOa+Z21TSySYb15fqd5O3e3nEwTEKkjb1eGZ2Cr
mhTHWKs7S9Yu/K8VNMA0JrcHbez566OnAEL40qckh1FviaY4l+BtcEJWWMWs2kxV
IKTEEHg1mr+9pNLYV3wcZ3m+PnVFSqW5OoeN3VJWxdHBphbjLcI/V4rD6cP4lvNq
/qsRYRrE21IytXWAuzlHAJxkOv8rqK56rSrz09a1SBwkrJ8qxow+DVHPbZmD1oCL
Fp86RN7Idfkjiz1PwpFPU+YViEvRy5c8v/amzkxswanqRVRcMvk3JVYFh3aenY81
ydIll+kayVO2GGEjliiN/eyDKRTZlSyfNDA38696/HAeYI2B+FQT9j06tgLXWF1Y
lvmx43oahoz/FQc7QhJmR3iE/SvZCEnh+eqoW11WIjgq+WZwcCsLln/H2+t57h9p
K8VJF+Pehgg2H2UCWwO3wb86OsENQCaO/1kkv08eHbfqT6KcmyUUq1i5j4peUfpl
qQnrVzRZdP9RcyELKtaSqFHb6t5YOd9HdU6kO+cFqhEud3br3jHPK2mlQFH6P5/Q
8s+00VCggX9i+tE4Im3e50XrVEMUVVQp9U+U0N7qS3w3UP5NIH9qRSlFCAYqq0sF
P+GbvuuG66laL8iKf1rw4ILmH2Nx4I0kQcPsETKTl278Rwnw2Eduz9Z4L1FNg29k
MylnZ5DlNPcwZjDoq3lvGMAusVXOGOlImIemNuDoCucI3oloIiRDyo+LT9wer1Ai
DBxMIA9ygWrfNOTOoe7obvgCDD9BjnIlqAiOw23Uuf/nA8nkwYOPX5sxnaH5HSUo
+Un6iH/x7zy39Gmk3GJ5Yn0r4pomCfejZV0HtWPRlCOWaHY8gKt5P5zN+Ba1mZ2J
id+A1dHXE8OKZWDEJq8ad3LZ89ZW87iQ41E7vR428QgNjzC7NzQnwF1TZ7zlfaM3
0KDkXxlbEe58jhxlURMw7cYNpZVYcOBHuvu43d73gKkngB2nufNQ8Z3utQtwBbYu
OJKFDzvexieP0h+UP0flK1NciKumXxBBSiBssA21FlWbOQaXmrJZLx1+dkjlb2Yh
2wEMQW6EKDOy9NgoE9g5ziDr+d2nLWwowbyYyIJgLv4+pAcznnZ4JI/cW1gn8dCX
wsACSwUmHy+JjndjUYF54dzVVV/MKLhJ87NOcywgO25/0I56WTH/rrf+VU8fbYzm
Q0mr2SsIuIEHean96Qmc90RTtCfBqHt+KAsDAXuGk+8QXIcOAwCJ6oyU+Xbfu46+
ioA5yqHV0VdKK23z5KQ8PtDVssKv7jMtNx6IoF8P1nnuVuqSMup3ZeCDJ2CiOat1
5OQNjHj9+SuGW8DjkXoYwYbQU5SvzuzYrQFReoCkZ8/G66GUbP792BggkcDECO/x
ySj6cyeBogWsvnHvjRoFW1TCEyHmCtSxStsr9mnOAKsygTGZjrwLVc5LzMW2rPLc
T+QU5WhZADqNFq+HU7l3Lz7kkAfBv+mcA7PHa6+u97ESCe3lMPrKLZZHGXs3fW2J
OZWizo44oLYiiv8ZhSnAzxG5o4OW0BLJCOU7wDiqfYtU9PXiMwzajakGHFT8XZLZ
fksaPKp2cIpto5icmqSFwUIutIWlpvuSYIY+2g3NHFOWIipAMF/Wu2IJvxI74JhQ
Pxl/CA1jJTALGUZEH7YGnN+5iZZmJ6tZedbq618DXVsEaBUmAigDEtw780jABmhy
k2a7Ds2KKyV18LpGq5HhWg5S5qDmz8ihFd3YM9A+3LRuHGjqx7PiSKUE6AUvQG2E
0aM5L+BPIiG3E+x2wms1Fdk553/+hO93e3vjQV4VhZRtKG1SmJ8PKhTREZA5JmJG
NDhnMFORU15rgibFFFU4TV3mbYWcr275wL/AWACg415kYjFJcMiw2c7rX2lzeQoF
bNxQxMzE/1eItfphNyV+kW0AUpXZ8/wpdfYfwJYAf8rKPti4+H5ZSszGd609hjDr
/7yCmXYOB0GPKAPJxWU24RPtYW5BXtHtzpbRGkp0rabWO+NDblV/vIvXtLYCP8vC
q2aj/xEUuZ8W6xD5JWYPY0d/rHguwc8pfQNnpDFF4Edr8/IgWT0Lz/w2zA/+/w3n
cw8Us9TsANvROsoQs2Pytmpx2srxrq/+X/oRaL/5wbP3ywVZvMf/w3gPOoqHHBe2
vlIBwTEvcwyOYrdPjJNjczKHElPeHGNwTGKyVDy76DLfPwNV9VuKx737ovwnLRCW
a8XaFV0IMx1tQu5meTesvjyuNHtQEZNZOOaVF5Y/Xuf5D7fCh63n8SYcNQ2pjjkv
MKrJkt9adX8OPRPuXCgompi16MQMtxGDAC0kPq/S812fpjmZ6geRLue9+ZKWp+K/
iB3to11RWDXmaYnJd+paG7qdI0lTfHShCOzWFZcyR4913m+ELwSQwLbf613n8GYT
s88W/hQgbwRDkUfQbCvIJixxQU8cEz1xvk9n4PfPehiYOD/Ryl3c+K5KtEnxmKeV
6+DSbZEI8iZXtfxgStPxOYjP9eCtAhJUHfEPaAmKF/j5ftUa9WX0RZeFB2A6t7Yh
iXLoj1p+tkJ9jKWP5BwBioGdERombXqiUurNGw6J+Odhnugv+iLoVorrmQmCPiaw
xBxu6E3aMeVzSwq731/TNSKeHyUeq03UAl8b96Vx4pcOSlkPLTrAU4n+v0abPdms
byKqDK6LunrE6Bi3vgxFJ5Jzqfoly7wIqxDR+6j/MiYIUdtRIXEBxqeritmpYfRZ
VSiiQJaT36nkNUzBcEvNHTymDs+oV8CMZVnmZIqLt9JlOtyOtsdS6uL5Y2C21skO
Dy11FnO46OEteQxLKVB3IOScoP+vRM3B+IYC8uGjkMtjTofJRNhuyHA/0PbYnByz
Z10iW3VbUiauZDxOYI6wEtnj+moKboFcNnnv8MuIhOKWTIE3OwZ6JT7a1zcf8Yuu
I+cl7ubUK9jWKKwLpbElLWRPuByOn9GISTmreai0SBtVlSnbapQ9gcjzPrPvpKjH
t2XV4WRS9gxW7qFx6oBJkre/DUwtP1qBmafM9jplPyfKcDlVl/3WbmUsA9qUuG/+
ag332XCo2oaO8eawYIO3IeQ3PQYIWSGJ9KDcUYBVLNsc99IJ+TSZk/DpIblx97q9
M6No/vnzbvHTYqXbjq2+iGQDptCeKmDtdNu/IXtaLRYIdt927CHc8CGIJVE3TqjV
qCzBPHOiezzjFcwAhOFIYTbXa+o7hW3c/2TAeFPcrdIDgr3eIyGqqsxcgtqWX2sO
EUOemTehz6nX2sQNrleAXmjhJUR3NAi6A+dY2AnB+uksuKRzDcuza5shw7TJZAA7
fMoKQTBTvTHy0BDtdpc1MEvxdvnxvErOxSAsfdNp7Or7qmmS5C9CEDal037RqyO3
qTXYj9GJ2qLnTntXFvxMmOeXdFq0Whf1pGldJemIrTVVYmFvgAf3/a8REVCmolxQ
apVwehj6qcsfIJVAHzbhqiZ7grOMgQL3rRtrA0RCWorDTfbqmbtYc07BBjkGtXh7
aGKms2Vk2/xeo0/zQOycy9uBHEz3En8huFrm9JP1ixwY8xwJeOyLxJ035zNIhyO/
FpYiw2Cmmt3ZecjvHxtQNicSmFohbGUmNLmNe/6GeNSsHvtDCbPO7BCvKLBvJpEa
LH0u9+/WSc1tiT088oGesBFe57tKstMUJJIaEKLSAQG1dX9HoGTQB9MO6Q2MT+Fu
d/hxUfOhSbZF1jgnhZYOSuYrpe4LKM8PQn2OBmvPihsz45JY1dKOkEupiJfSwi0O
IRXQcqt9/R/1JQthVgso90q6opQSMTZqHlz863QkCvuteAQItFsS05Tdy8EmDGZK
ysXcbUmYxOHphp/GZS6NzSByNFiy36+pL4ruXa/uMacnU6ctdzDzl+jOY0/WrLpi
1d1gRbWWnZnAssUkXa/pnKuwS0ZrfFGCHzLNjlyLNh2YDy7NRYJpUq8BKL0iZzCT
O4U1BSrOMe6w3JvNcrL4K443ZAbqr24W9xwEtFl97lZVtna16s9AKxc79UFFc8tj
blv8SZuR0R/0EihKlG2MzRjEqjPuUAjUC15DykeMZH28VnXcqaa/zl65SZMZao+D
SzNSHrPbZbtgcBD1JevdIhaLsKsh9x34E4i7B5WQ1iK0If4OOL1xfjkkD3cN/62w
e1p76L1Hw88bw2cHl2vmvKzY6S26SaOI03C9+ou3GrqME4vwp2jNCd5hSdcfHg8l
q2hnNqytXO//XfYZkggVmrHOImkpdxB7jLrqFTSN2edGQLF/FJlkEIQqABLM1taz
w4Muj0InINvupc3xF38rqv96edE5CoYiC2uFK8vXrqU+F+eWzbH78Yz54WGkmKaw
8bS4DJPbqgMGjrgSMP9VCnXfKparfYPj9J/+dx1whDRPH9nO5S1jzT2T3jUkAlDn
OZa5FHd2ogNYiKvFV9UoEKaumZrUZ0gFyo5s07oDldnsU6DsqydPcoUg6crkvlMK
HSxkxpZNbbWJ+8AOevfP1Uw0WS5T5zRM7tG6ssV/4t3qG0gZ87NVKxl698kU8ep2
ggxDvPbLGmKJ+dkx4QHYgAJwKdd7qHVIynYtupqG11r4dYgNapV6gpUumkF5CPi9
zWks2Hu4lJ61DZ9E9EF7W31LRYztri86gelGjvVVl0pxEeYE3oFbgBSkZiZ7+Xol
Q93CdwvxLPc6Qbgt6ST0Bc73r5X5Z3G9xIcwUM1Ll/1njklq8NJeaSFilij5omjM
uQrb1V057/PdTuyoBts+Il6W8vjbqaz0/aT1CvMR7vvkUexhrS7h8QwHKp0e0+0A
C9InJmsd9rSaift30rz817XAxpQqazQ/ECkijfFGVhgSdCsvI/j5ytfv1J7uvzqo
wJz9g2K/cPN4czi+KHpyCf8fcp0rICuGYbEjlkIptYzHcSWXlfXWFef81uh9dSkA
lgwvUqVoohiWOgvEBWoNPPrtDFhjDgpgF+O0z/AyXMwmpSo6mP3umJuMFYUfzT9j
GHG16elTvOXfqHhOd/RMe1UArVGcj/y6rZ4TedacpqdWme2LGhCoQJaiOqQlrgH1
OwkN4zQyT9j9GazvfudIG6c0aBxKiCeFSr7aope6Y7vCY4W4blYvfy9HRnvGrbEC
PC+2DFpD1twl6cNbj5hchMbJW0oHovgzZ/z9AN3N6qIkzppXiiQBIstLYaJsQ3WM
8MUQoUICe3BxTtmC9xX13lg2r7v8dd6HJW7EJtZ350lChkRnkpvnX7/k1QaINFJX
ljS8DJjCpKDVanmzGoL7kWBoHHRDHYWNPfyldKYOgMps6eWa34SWDrVoSow5Tmix
wQRb7dv09YUF9yH/GxqJ4ebJDlVGR9+afUXoBQAfquhDj5FIqvIdj2UajFjNaHGU
ztBwcsnLUiAa7Aatewj+pkGEk+Phn9RrUR6lJaXSFl66hp9H32iObWcpNAhCArcR
aDrKqLqgM/T1ViH2LoAuwWazVT9CITkjCltwVr3v7cTFDpRBeXHbMzVOtWcyEW3e
H1KfuRfX6QyLZV4IvXvRd4gYBOABV7PCiQPAu07EzMXxivU28vbi4B4+00RAabYD
QvnQy54mi0Fu1EK0E3fPAA==
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
eWG5UCqZsnQTkY8nX7W8PvnY4RL6EXG7kV0lD6jwoE8WpKbrn3YSAKprZCN29LJ4
gsNIDCdYB7jNBYT8Ayw2ZO/xONyqyBuc6NZw1rPc93UGEi76tZ1dH1S69xXNNmrO
Oe940YkXMupYwr+EDuUvAWJgPjtFZ0TmtcojswfgQRtSqWgFdUlh6KAmahaus3ig
USOsnBPTLsKzOG4Qmk9zN3sPbMT+UXY5ru2baGzPITBBwStDlGCP/IH61WyGh/Vv
59Bt8ixw98KbzFEyEW7wM3O38oSWD3gRughk2Yu3+CdXCEJ2aXlIo2OGyoNAmL/V
PdyThslJsWclYXnC5sGBRA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5104 )
`pragma protect data_block
kN2rLh6yEm8uxKtcnlPu8X+ed9Cofj56BZ8IyQTI3f2ern8kwZ2i71TWfNF1hMZ3
Ve4Q8BQBxxEOoOyqoI5kT+kyvFQN6ce9m/xGGtPRJYhtNf7ErgO1jHbEEsSjUfBY
gzqHKxdg0jamopQi/hJXAoGHUnaqJq1S6a17W3cRqMTiTbroj51nTnJfHh8Hr+yN
7uoKtnYKnvdo8Tj5ll8M/6Q8KrQIwRtw6Z3SUVcno5sX0xglXJvMYSDWTscHbj9W
FXI3CxV7+kBKesUiU+pVJZv/B1NyqKFYXKFRvXq1A356edfPamLmtqaLxZQgGlAW
NPx9r65ykuDHV3dxzP6ASOspwLQj58MKo4+2/iclwPLw8IcVkeRZg4Un/QTCYTLD
Er1Z6ZTjsWUDGihEldXK90oDNKvEYYt7T8OIucWfCedNZd8epwtTRZ4evdPZjlDM
gb25dfCmXQDZmZ5B+u0yb/Ww558168azB7rbf5RWndxjrUTfheGXc0LXFCXdRXRF
MttN9jqkCJ7cJEiksQPFr+wBn4AcuzwZ9GXo6zcOaTnlTDOx8xFpZFqzRFhBImn6
5vCD+xW8K2rZsdEgyLevDGckQ3JftR3rQjDWkIY9n8Zx/Gt6NojLqckVObQZekpi
1jXSWYnT1Ngr0aAwkeLbuFfknoOzgGJGhqkO2g9aYGySfifw1PqpSc9zxPv6cbn1
lKPkM5P+YJ+ceHQhWgjuvWg4jzp6A1PzNDkdg5+Gt0k1QXS+HG5Em/uJkHHQHRc9
W0/YrKDofM6suNuAZ++UD5JYQYRqJXky6xZNtQDWulxg6XGvZ/FQTy4OmJ2DIWJ8
eA+1SB8UIZItQSRksQQQ4EGBRN7ibpuipvcSBZ+JbLnJUcIDOCc1IXaGzz/HeXW9
qmWzSpxxTfAcrsrxJ0FCHcALv4LIlP9+Q7/RVQdl1Kgl+9co1LRraXDEkJ5d48C4
4A1q0nLw46oO7WmZB12PkW26p7YWVM+GW+eDsfCLR3YYOimki7HD24kQzurugGEQ
0aFmhE0XgN3DcIPi0B/c11IvBJdRB7s/7Mus04ypahOKwo/KF+1A2dtTisqSYXSW
nYAYKnFxk7RMsFRu7yixP1ElAYfqMLd2lBqrXLVF3CW5D/ZkqQKTlwmgh01rK8aX
ay9cg81l6AhT25bV5fbNlLngPU+ISAT9RCQlrWa1EItS4HaKOyMqNqlU5oeexEs9
ywf0e4gyZBshLRNZnSXn+fO6F8+EOIPj9TTuAxMyuxPSU/BvsOKJdZ4FGwdjnrXx
5Sv/+Gi1Z2Gr5c086WIFUBGD1aOzvtG3wZVLZoxL2IO3WCeet6Y9DD9A4NqUJrl8
StjtRAphi8VNztioSbPSmWeBFSH1OPmBDFp/BA+MHgJw/yaKGHMwj1SGtUtv1QCS
D5Y/Dtj82CELwoeGJ8hmNOQBF+wLfw8CDgSZwHO+H9lqXJ1rvu2OqbHaVf3yqMv6
Jr2mSWAm5WFeHjlQTg++jGB6TVJS7R3LyftkZaqgZdK99b2U/m42NqDUgomn5Cwh
1Po8BblacN6Jlus7ACqQtzT12QgEhVkocJU7vnCGA+qTOOgUQHvHPC6nczYfTg8A
s1ZFkKCSzNskw7VrDg93faed1j3O6Dw9k7IkOOeTkOMkjAHNErCHMMefE2qoGGnL
I9DDJQZ88t2en+mpzivnmh1zBrDczB3com9Y7V8WwV2lhVpkRJ9lUq6TLv+RBdDD
cw2fxgdm8bf/2pU4y96gINvMuWW8S3uecCdySZ7/ptPB1ioVnTHrERIvxASbbO7w
L/gxkyTFlnm48OcFPKXvNEvZUlVJlQQnXzjJ7+1QCLdPU9yPrhEAS2opCUNjm95w
fJtvgnL6fIQwoy5Z8yIz4bQRKDiFWVdO/+nRO7boA0Qe3KKfgTkKe5704RogfL+R
5gDI5u1o9xPyf93Hbpm5pXz9ZSGr1xKRzJmbSfWopxnuliEDnXQHNWJziF0JKdlK
P9WuNvCXtwFp0u5eqAkFO9ZuGaN1hgT3UTWJDeD4o6r9o2uvRiQiS84JSADvx6jt
NUoHFa6Zre41RdZBVrnfl3FoX97WlCJtphkG2Kc+QOLeG5CBhkDZk+wVHhz4BlH8
x5oKz94sypuRK8c5Sg6+iiavRXNn+t1paUi+dwYo0VhCwKY5WRe8ERa5klkH1tLI
yIG7av1qhjbD79egbjJMrn7t39uVaCvoLnPYx8LIxeseJgwG9r+2LvlPazw8uUaj
msZTI/n5DCibee9osgK5iIgkSNFgLeiNUoavH/FxKuC5t0B5FwA/s4/pCN1UKn4K
6WXFyp6fkuU4vZp5jgxg3iCa49V+s7uR7Q/aj9/YWAG20aNQenM6Hut3/+5hm4pZ
exJM9NKHlhRMLeGlhano6Ryp11OO3dGHuHsLgPccUnR6bCWdiT8u8HhQSbeRjoMI
I06d8E8vtGm312Es06UeRxkGQncXecYulg7+CAxDLQNddxl5Obd+U2iePywlCZ52
jy01PbBne/Gd3wmw4DKj2/Ig6ya9fHSg8Y55SuxRdomk+E4i15rgMLpQiaKeoGN1
CI5QwpTESSamDiYagMHFkqzQ/DH7fjLrqaM+9Jqt8r3j7nEW594Pcn37scpFXpcT
KL9Semo7lWP65wvkb11MUPe9p0ADgNSNbB/YlMM+DuMr7J1/sfYtjCU5TREb3S19
mRH9tM+i117tIh7jXbKb2TyqcCLQvr9Rlr+KxD1XXZ6QWasIO32s5crU6Bkv9aGH
2Je/bfigcQX1IZCQk+hQy8l8SEoBcHALH3xEQYntCQMhB6mUMahOHpG4QNQSR77A
HOa0/RaZM/2a83z4hTPAt3S4KS7pCn1KqWJr/X6TCciWp/Z2GEzYiISnQ8RSPVda
JtFIxsSB8SYvFLVUfVQxnJQ8LH8d5Xwg9OaBJ9E+ipC2MfC24JB7hAy/dwhBPrwe
L7gUZVe22tn7XOFP5OIz5pkqCgubbbOrDdq8fpJMap4GCZok5maSDSrjKfh+f8vN
DhnP8Cwps4bzeeWJf+HZfYxPCYwbKKQ7cQOc5VoLf2VuL8h/5gu4AxFvbbu0vDdJ
CONrI89sLR7z3uxVAZyLtfLSD6gOLo6A6anrXKdgvwE7wl7q3zYHkltJfoyCs/YN
4fCQAGi8zSJoWJ/4Dhj3NQlUtC7pCUGDdr2CVH54VvUgSclHhGaj/KdkBl4PxvR8
DP34Q4NRUmXW7eCnXbJdNKOwOjtc0Ri5A6jY6zQoMN3U8GFblNz3IbIVuYZbFXF6
Fb3JUMyBHA0tn4hQ+Ok1wB7rKtPEMi5N6H/Rnnz4krynlNVZKuoa4Dxt3A4E+mBx
Fq3Oy8Q5puMRqwuySs2bxIi1fy2M3bBNY+kJvUJUCvh7rIEf93oBH1znjMCEvSG7
JHF3HgsRZQMEXwCDyaPdTOH3d73lsta/n/f/J2g22R8k3IimMPbhTRVsFNYOB1NG
m/YeOkDjFG/wHOdq+4XhOofDDpAdfBvfGjI3E9SlUSVCQt33DSKNGrC9h54svzo0
kCSF0o4X8znhuKYkkrGw+VusOOKhXiHHTvsEEHLZ1RY1ZCaSQihkEGZsSirqegN3
0hJjLA5yzOEI+1snUE/6Em8iM9xtV27YqqXpvjuOMUd/ayXjx1/rm7txyDi+/Opf
KWKPVfJcCCtFs+aXZYxoBN5jc6fD0cJj6M/OtXOtXMqtEbahGA9fz5YW/D3CmKda
T5fEA/irHSVuxyAMhKRAv/aOfwhYRRpaNEM/TzJLtXa9jBt/EFg+WB6u4v/lmMCU
bUiQFjjmypFG0lsNPtyQJ1M3p7BznCK0E+9HkE9bL7p6Q62rI/xQTDj96EuE5amh
sA3Ar8BSmXwSY4eeJdCAUnyA+3ktqhlstTfaacrSKcBTtwv7uDrO8plLJTIQorw5
mJCqd/fasTUJ9kg0xFrbosQ7iTNaNCvZBwwt9Dt+9SZe6cdBMv/GpTJblSMcchYY
8M+NdPYoJ/jQn3/QoevhEbAkHvE5CfXfxFWK9k4zdfm3Vxw3QWa6T4w6b3gFT2Xf
96AZRVNIcf7/6j9LmsHGPUwtjuw28a1eiaM/RraX4FdsGZ4Na5bHcD5M6am7EPsp
pjKsGjiYeFEiqSHDc7goj4CiHrE2FE1+TljQ43QRkJknNnWCNETTZ2QfrSsFrTpB
7e8k1btWl5wf0sQhzzwYdr0SOJfr7OnvOFYHoucPpOXB3Wei5U/oy7jz4lF7u5qo
MkuM+WD7QLvngNPt2Uhmvp0h0uPp1L/3169/WJuBbJPMR+LHZad/uUIeFAwHPUvn
ZJzChhDWh/+tXi6sgH1ijx5dLH+Ksw0eksRHrmnaBo4uGLaJsL4M7T/958nUr4xG
fCZvOwizBwFps+RpDvubulkgePS9D9GdFKC0Q1nIFFpvoHxhoxvATsvdemrfz46j
XxgyNwBTUwV1jW58+/pInlFia0zC+maWGNy/I6r3LeA53VcH+BhGl8zTInlZiJR4
t7C2ULrpdNWfkF+gmf3oeTyN3VIwUnuKBMxQb8a2AWUgi+s+9DNqslWJDwbp93RN
sAcd1QFnrEYyTLefPnNmRY19LPe57An+GWeVR7i4bzpnJQBDkGAsbkmg96rLzHOP
7doP4/nQczYs1VBKHZlhGLbMylcc5B+QiP3UpdM/baQQFAqoax0I0w1zjhCR9brx
g8U6gvK/rReqTCG29+HotssCq4j2ZUQTJ0CGuYwzOzFOpQOId+Zs38dZzIxDBoWN
L3d8Lq+JnSMxv0Sv5sMeCgMdfGFkuIrJ/0u3sieh1gjq7KBMeyyEMz1C5PevKYVV
C2aXPXuVmQC6vHiwxlNpwsuqcBG8ot9WykFWzXemshtftu5DBSP1nZCLePRP0bWz
H3hdnE2OX09z2cd1zYYLZmClyKiLE994Cq3dXLkhZ7hiqeKC8EqsDL2vIM/5ckYF
Z4NkObM4IemXOhXAYUfi2REHEgRuaj5biM2gABP4FpYM1tdUqHmk45bv3eN4VD5o
aSwqchXxlZ5Xk3Yi4usI9g9lLt3mzLpUXoM/w81Ge+xviK+uA+fQx0jsmPdjpXwF
Kk8PLMBzWAxdt7LYpodsKmlUkPLTwb7MPXQi6EA1w/Nm7+gqLCxsnV0ZwX9cqOt+
xFp1I4n9O+ajHVA0dn+Rinn7OtcVOY608tQk6KVdNsOV0c4eYaTu2855ZmJEP02o
ue2VfHRaogusgnAu84bWK1HEx/AqaurSJsk3h4+9nIf0dfI+S5HINgZg5xzImmP8
y8+a36luMchtJoWh2v56akA+9MwAtQebi/qMkZJWIgRkBeElPtgRhmohYQN98CSO
kN68o0rS/i+R+eie11EXihr+h+HWBRBF0hW4run7pl7qBkKPLirEcKcBcj6Vwr/T
7CHYcuqgyUID76ukvGfGoSkpZX5JRSGwtsWUa6BJy5gFe7wiEpFSdp/L76b5A/D8
fcyIAANJX3QVlLUZSk/6Kq9CdU6ItJPmsOGTmsBwApJMIDHICEqaiEzDpwD8O9DC
jnOvCXBNMVrFqKm2Rowld3T/lGBjg0DDXjXtALRj41mbDtuumMsc0wzuOqpxUTDH
PuEHLnzD6xO5KHHj6XHJemqCHgJcyfdapZWWu3rRJ6eaOUvwpG1nCD3UUB+8hG8I
SjsQP9GPjtehic+1EiKgJS9CGg+o+8n+FaB6sFkvUfR7ZWgfR6nb5ECslMfm0oMm
iL5bBjrBNitqcZ/C0mKZc03FpWcdcmArWYUlAccde9ERMp3INMtrEmde/Nlu4lLh
FAaRXSLx8f3Ue7gCJK5SVBK2z2Wu6gcbxsV79Bcsl/xy1HIkvONRK4LAu/roG4Zq
jKkE/KXa+bVwC/i5qn6mKAHvnR7RZA9HKuR4uwXFSRX+SmSc7idFMhhmoEtxuF9j
XzC/IPdvtHCMlTepTY2Ml7bqSTzTBXT2mD/aMnGZqXhaMw/h2crcenpVZSxiH5/j
1qIh70Cxi835AGSSCvPvDRoYGSKwGDr+0thEZngSF9vbPrIDJGBKg4T0q/cErG/9
9U2PguP0IdqhEKfwBFQ+MObZuw2SaEg21Ix25PAnJunotquqE3tuVsg1DfI9Zy6D
5warbjykAoIJa7CXa1euIVIJi3vOX4G5eQfe7FP6t4O0FTOFRbqqDLXHRoxPRBp6
hFlTrX58Yubq0T1TzIstdlOX8Tc4NchSQySrxmJd46VoqJEfSKpvQ7X1d/f0uZ6V
4CBPnhN1pGvH+2G6l67oFsv59lUgzt1ZOj9HE/sTIRvoGTSYLcVdyfPPSJIAuV2M
fXSaW6cuXS04d8e58+dTfEZ2kDaOn21EYkfVNji8rZ+ScbxWENyfpDoyDQ3CIfzT
oldMXTbinHHJ3VIAZg4mo3qigA+BU3QWrbHRqNIigsYXm5aXsg1oi/05tyLb79q+
F+Ao4Jav/adr8lTQCpBV/++tE/lAIeuEwSH0HQHw0Bndu7BjtOSg39oZQYamfYiW
GBaLOcVN8YH41Nqjr81lOlxgo/ABuJ7t4ycfc9jVG20Lj9XSxLwdgKpsaCCgdjAr
hGbhKY4rduMxjde81Bz86rC2sKdlQEsH/sBnkBiUrh6J+KyOnkWrvkHIUgz2mwYd
2L7+upYfKGzwh07YJioTjLB341Gh4eWNTf5CAAl5VUoEr640vN+iHCD6mcZBWnr9
JcldrDkbYlkMEGpC0eW8EDIcr2aGUNhO+JoEY9cswsZMinW27EoOOA+R5+VhNPU0
flUn7/EmAI9S0lOCutEyXq+unQjckzv1SYQiqNf2PY7eXBOwCqn5FGQoEuy7QdHp
yt8MjsfTtRL2KQETGzdpqw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WIVUlgHrrbEQlmSqUjYnBXJ945TGuU6V87GrMD+HowlFm9eBP1XWjUwG5MT5qRtY
RPPHOXAzn3VYDbFm6r8b0Hn4dhcu9+mhVUbzDj3uw1GIMHO13muT7qWK7o7jGXLd
UyihXXcKCPb+9eJioyyPKEiGlt4RrdFQF2ZNmIyEEzUXC0Ty85j12/5OW6D/BHS8
svP+qkSZsbr1RYuyONHYPn/D2nZRLAaxvkKA8vkS9DNjITw50QU3t2Vn5GZRxK75
PzUlxnhjLdZEB1W+gc1dN0zVUrxhmjoAoRuc/HcnR9MRvjyWbWuRJffHeCKcBipk
F5EqcN5Rl6H8FPDXwr66pw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2624 )
`pragma protect data_block
6zSLqFbtZQ2Bo9l9ejCjrd1FtKkSeLzwlWxYOjAsI4tBuV6IxECEv4zGfElL/BbR
k6ChZPcrC8Im0ZmhmtAUbgekt1PZ/BUjnwYrI2jJACTUV6eVyuiNQmtZ1swcAg17
MCnD+Aal8iDIU1Hgzl6VpXhPZ8ofALuyCzfNgk94yjepliuCmEneNOUjDPwdOtXd
/bSqMFjpFEKB0mpwbZI+13YvPveSDanD87GITve73SP77kVwlODN5CaF57+wx6i9
LMai4QVfrMyo6qBLBofRm5KjqHehz3tuknr6Ky+MltcaU3CfbJaAnH2cfba18RoH
GRDfY5yF1dYBdHWf7oht0j2Xi1i0/9L2Csd6T3gxCMxZNq698ODVU+vpfzMAIEDY
QPR0Tcioj68KRuPvVcc6W/WmO0aliV+z7BIFn4WnN5d96VvtS6uS0MpTszO/DivK
IomZNn5s+gWpx7l6oQK09OBa71//r7ka3osIlmypvbDnzDG9P82jrw8OXjhxp/1l
jHZ83a9er2kAeBLI8mhI6+sErcPOkjshFqOCsbKoBXxNca9X2i2k5GcIRq0Qv69c
1Q170ZTqTlJDBd1s/hBUsatnnNIEivKURPsantjE4Gv45gyqKfXS2bFK73COynKB
dSFkYT3n8mmS/rzILS/SNi/Fcb52HufCB+3E9AKfVliqdPQlNxFDeZdSllLIYvWj
La/4uqmF5ZaRqrznLhsr3o/GMW2WiCIEg3GJnu8hcckGvUCPJB0n7Kk5L6zCFefL
uWadQWsh3kfjz/KeF8OV71R5Mp6PRWlwZZLNOsVperWjkYxXb2i2vpQAJ4XRiRoC
5evfErJtWAw23//bpZ8lyTLXnkTsXelUyLJptGivQ/ylJprZ29XR8aSxZzG3kH3m
Zm4zQeiio9kpc/zfsYFiAdg6bUd5rC92G/LJL4tDaojYVFKhMAQG5iVYIbDqjSMx
uytIetI7TtXvyDwS+K+kHklfc/xALTLfr+wPHQp+15Bi7vvsl1rTozV5tomsKBWw
pTb/dea8ulNtXLw7jH2yFYBc3Azlgu7BymGcn4yh/3bhmYmonzuXtWEhAM/GI2+F
zhKa4HtaOhSopW4ccWLWFfZ+CuUO4cSFD6ftU+g9G5UEj2j21g1oaUeHzYOx5kEf
w0PaONfls74vkMP7Y8JRSF0t4A6YR31KaGyWGUTLon36WAS753+xtzN8/s5q5pdn
7C1IeWZPKGQcLf+FM95v0IDgfF2oFi4QZNB5LU5LyG4CUfHAFYMpJtK89O9Qus7c
aCjzxR5xwmrNJovVwQy3XF0hT+tw4GBZOfRTdcgQNOlvBZwFYEbTjRADUJjfCUOa
yV5M1/03bZvXa5qCpDjB57V7gsO7fJQ8l+xyE/Fq435t0CGRvsuqqO7gp4mT9iHI
PvjVITnOlVMB1/N+gYjHA9Aj1jZr2nD3uPMNueherYH1f52KGCNIvqiJ7TQefbsR
+LkL+Hx/+zBCp3FN/HdRtUsaR6u8hmpfAmaE/pQeLOaMIw6Enfdr6pDKYYe/j9ZY
rRdxCSx1yZ/jJsBc4r8U6/6tDEfHJCdVnf3eCpd9qqbw4qv+hM3ktb5398wbiyOf
XxIgd9+CiLQAolbAkwSlk/0JfiAqjLUqLnaZGeedHUnQKUwkdxBk0Sqt+kOFyPOF
L25UaEXb3DzWBE51EEvZ6bbSXu6e6eE11fMbsCy7xK0AGXuaeZuqCVVJq+v58ohz
3GLN57MoNsiWUrvf1JloYFuj220m56GKCWOFFqWIbIJf8kIvcrffPonPxLXr7BLE
fvtMjt7EESNnOuMZW9WLqL52qJHClpCmW+HYV43T8t4OqqvRHaiugwbuG9YQeQC2
tJAcpHUvfvDPxja+AzLeZiyCJloLp3VvHvJisLvPyN/e04wIBdVyT56tnYXWnrc0
AMWF5LnYnCTmYkyxDTv1a1YU8MZLJDzj3GtIE7ObOlwbe8md93c0ABD3o7m8Ajtj
LjknUqmB5wb8ZYVfQMK0AgYtQcBWTNzooTIVh3rkRH3Sro6nyRxzx+/d1PQfDLTM
pW2w6Vwg/a64WDofJAH7UweOeSYB1meBLxiyGYgm0d6oKG5aERKFhSMBrI4lc78K
43s9+h4ZjaWQsLMNWWyUZZqVIMGFK44k0qr5iL6uVOIb9vvmo+g/v2w0O0OUD2s/
RpHIZUjcFeRTRTScsoE+pEtpetiGoRusZknrl941bwyVdLh2FWlHkMkBBNKLjhKW
WnV2ReUJ7RCoFp0L18M4l2WUueDpBva+uzzVkqs/9SBKnahPLVn0MLrk2HThvG9r
+MvpHWmyDv+YM5pjZDC9FK0AcjNpDbJ1ue7J14KvW0NNcRexZew5XD5ht4HEZe+T
jk9ppZvIPrap2bIK1Sg9NLAjl3bmfkyUTjxTmfpKuXhH0Z4SthVQiJfPdg1RJn9F
RgFSHwQkdfUvO6ZCh7DlrbkoNZYHIEjjO4ZXcaPCbY/1KZD456tjV9zcUGMnnwrG
XwOdDtG9yBDu2MO7SUeB0xb4iKd7dxA/yyHga4vvMNQpWdstSPfCc/Vwgv10BkYz
7wsCByds/ZBZBvu5DkOb5rldeeAxUchz3NTOT8eGMys+KANv2gMnbBq89MOfQCTz
6vYbTR4bwRFNMf3pePXaTALpE03b9J5YMDDjaAIr0Qp/3o9XOzKvPkQIUfvKjIKg
IAYCWdnZD61o5P8uY4G9iVOjlBEnwc2A9RtEYR61iz1qDjZrtrzbMBxGS+57AIYJ
xhp6td74cJOuCeoF8rZ5ULvPxGH5CgwqQ57POHcoMOy3lKFpHMHM8mbEziEaFsPl
vXv0IeBCaLX8F4tpd7VX7GyD1NehcLLYWGqn0ZF3832wIhwVMOU9mS2UKQyf3gSf
457QdykTBXKnc4g9RRQ2QvKhpWYAHxzdJnNsFrCMsLF5CmaX/kCRxc3eXAHq9OwA
Q8aeQieQIWOhkkm3Tvu8Pm3kdPpBMtNXNRXJiileDcnB/4HhjhAZ4COhaTdj74qr
N5pgZiGG0eRTNax+BbAyCLIWjwleIJYv+5WpuGUEKMDmYlP2L7QSOvJeoXj9WZU3
TjQUpn8XZEy685Hf+3u3mV8ktEGd4IdmFgesXiY4Rtqd5RgwzCWOF6dJmrIxiUcZ
2iB/KOjAeQjWjdNP4sydZlKCbFlZJpxA6113pFoR+fRZTGuqIMuFGdk9Yof3Htpu
tPU8XpYomB4NR5XhjUZv88QaBotCjKVHcKZvog5o7wpjlIlsIvul5peG3+qTNIzB
z5SH4A6aypNkumQmG1TM7D6Nijet5qTfTpEXzkFxWP+EPr3xTnc2Xw0pQ/Le32sB
jQVBw61RuhU1MUXktlBups/7nqzIaRVekweZWAqry6lUHJQm67PEx7j9etbksRB7
qoWMDC6TyMpS0bU5k6TDIDv0xC2rSq43o6frrPE7DhpD7atg/gW7TG0f2BIUr12I
AR6bN1eN9gThZNqj9g9XYhj7qu1b6+PgOv+cxnBysUY=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WnZ842WMMTt4a2PwdF78iSeWsUjD9vM+yC2DIuUeguJ7P9Jk2sI8mc9ft5aYtdLF
zkvqrPPQsC+sOtAN6CaFkzCf1KyR5YX40Qlveeu4Vbm7oSSanMsA4LrkzJ0yCydu
CG/8GDUOTldRAMyxa0rRpRyr0koN8Ut6QYKIGI5OVAamdmzOSUL8s/kgauIRPQ92
Tl33fjbRXH8qIR6kbmcmAzto8kQV8qQ0oMLerzSTUVHlgDFdSZ+UEOzgaI0mGD7f
P3IV4CVQqUP2u5wCsU+XH31f5bSs8Y2QIdNekQ8CcC3gzppR5JLwbKcy1xUc+sgz
9G7y2Yu2kc+Svlhxo4WbFg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 18528 )
`pragma protect data_block
ft+im6/k0Tuj11IX06Kz7G4jAy1dvxAkazxXN/owKxLjapCyCHWJ2BWepmohqaXr
jmzTxBUqcJ/8WkMlyBQg/sgVHS2AKvfIu63iUrZq08eo0PIJfl3G1S8oSieiyIaA
l4l9yhpEIdd4sjP9rEBk5g9FMOYLsbi+AFVgA1dS+VD70tWHh5ktUQjS1Vywq+Y+
tKMfxOTKFsumjYhHnNUYwcWMFr1pER9RoFgFyFB82JV7gk1OdeQHJKXPeJ1Yx2AI
cCS4RcpAOaOeBecBgbcDAtLwLIbUOtBwqVKzP6IuqOamXLMon1aSNUklroYEePi7
PPu+BPEev96R35NPpp9z+NgfsLU0+yOqyiylRUWhomuN8a8MJN52gY4Pgj767hzW
r4Yvdk01OwKQUDQJbkR0wYdg6PwFCvojo7AlbF80tNexUVWg2EjQ3yr0mZxWDV8G
v91hf04pqsJp7QL5LkD1LzrTWVKPEeY8xO5fs+1VAT03LhKj/i5ZD6l8OViZ0lc9
+gMvpIbhEEZyIlQel6gNBOnGhpAU6QZV5xfF5XCjq4EFiZazUqUdC7ZCITkBeoTw
Uge9xV2rcZMhmMOPJf3RZlfYgcrmgzCJONkPRII4Eyp3+yUUNHd0b8llk3t0vMAe
AzBF/dH97v3zLBeqZ7BfJmJ7/SX/0B03C17NdMl7o2WT42iWW8FxxEF1z0NoBe31
tVRbDvy5sfvDLwwBRA1VDl44zeZ7d5+frTBhoc9HUKtA5eVLJ1DYdUlLDaBTM0ub
puWD2v+zZcGKSvilon00P92QK8RfNKNvWSgt3Ig/dVXBCcIw80JBVmAKzNG1xPKF
XGmrbGiV++HiY3Y+Fe9bxSlsAaVf+FjxnsyPndeuDk7BgQt0+igEEdjiEkgihEjp
ijyEXncWhnV+Pibtqf7RER2uyajuTOSNborG+I0ZfnUB+wSLkdOH3hXRw3zASIWG
EHi1Z+kSuTzJ9X9D2VrpizQaKcpiOMXIzHr0L1dy2ZZ7FwDVXAufN+L2vaY9Xakh
1EkdaytMF/69nqJ28eGHhh9lIajwc2ExPww4OCO+xj2dtW3SZVDBc3PK7X65daor
g5S5ysXBNE8YoNqc+0tcFchatJWzAhvkiQtRDligodpAY/4jQrqkV+Sz1FD9YHju
JgDbShe9hP9nH4kaSPEtRxjuQ4NOyVUtQVjV4hhdaLbv0loe1CuDgbCHJRWH7vGR
hZoURfdgjjtQAbL7GrQuI1ASXtmW+VQfIQJitJkNcmpnpy12hhD8zTTIMioqk3gA
zwtmGJHfwEb9QQegKCDrGlOi/xYWl33jayTNPNEDntYOixUlaO+WHp+1BTHL7HPF
0+uPfVqmLlTm62HnoOZ7G4oOI5vZnKY960QxmkBC+V00jMKCRwYqug9sp0HSSWPO
0mb0dxaZPUIs8TUohCu4BcLA0N1NV7JS3zcXOMiMipc9hScNUVum0nXTg/3J2Pom
Pj6AT8el6Bcmz3/FYhYic8jImMuAacEXCvEm+/xM7YoNW7eYWM6qU9AvnGe8g1uj
9Cfo5ZtB2POy3tH3KAfgty+miixoYx6apdQ1Crbfa+dkO0tlAhaUdBZr1PDUQaVN
+Zd9MW/x5XhnzlAVseG40gWp6wfU2JJ/ZYAv9+tg0bwYq8y1bUeItxf8wxTu9EKP
mkFA0jdKH2YZCCnE//IZXU452EVpF4I9O0tfP6U7lmY2g6/OElgpoOt9GQXIXZpx
CncekMiqanHu9ANPQkXml7KI/k6TnBRVkG3cN5aRgTa9e7+hyMyos5lurdVLQz2b
eacF12OJYZ4QI7UiUxjVFmh226OkN9mR8A1D3Eor47CNq8/2jpnrMmmlMwGl8n1X
lqYR4EwkbSCLogo4rW5FWjEfjrEJ+LWMKVw0mPoi+DYDJtchcUBN1S+j2rFdbAoC
WVIs7KdjUM22S7GYFPVtVpia0gksdcXGeBmbXWC+kSoAHuDL+b30McfW1cf843Bb
YqeyMnFu8E/WGHVkAHtSHEu1899sIRxCcmgonwloNVo8cEOcFPXTNmq+EugojOGT
ZR04BSktsq7xVcl/VY2yW1nw7pOnpQSW+Ndzvw6QnBXDmHivcHsd9pYodco/Tx1U
6TcC6Of9nXT4FvXWKOXLFiqfZZQyXH+wlsWTpPDdktZtZRQyNTHeM4vQddG6Hs9P
HAK5NbIzFX5AP1CWBmk6praZDtKkvLhJ7/1tO/Ji62HJ3+x4L2PXlxsNmIkVxPGy
V33DGWyeQmGgi6CiJq53reJFk4g+4Ny0adioDC9593FC9CG/D8gJcWRgQb8zi2gB
Grc9ldOhvGnbVnukbSQeYXBRcftsylAubSHJXJkbORyq++70m1O4ejqoTuV3JxiL
1f5UXwmH8cGdX2aK0r9++t/x3cX4j81FT+pAFyl+t3b/dl5oT5NSe3R7iDT8kDrX
Cc95L4koJoV/EIXZ1uYi8tqV5K+ms/ViVBrAHNxll8vK1wC4U7TJJpTd0QdU6hBp
ZEARe7uwKd2KxTARqi/S7oAG7RVS0mJ8FG4yO+bAby1G1fsQ6jFHqQttv0xflrca
Gs9+CorJP14Yum02bBmK1xKLjmmCN1588Kskn4r4RK8JX4iGjiRf29IjwoIUIzgG
AashClGyFCcEbYqqTwGM0cz0/XE9wHPcwFoIegdrswdHUH/ld3PkU/by+AFtHb/3
8rQ489PK289KcZ3X25TzxkAr1gozkmCpc8P3zifVabGcQEx1S4ViLt9cnxxJb3L9
6j30X2quwswUnlX6nF/JwJtRU8uqTqxXDqdsHiejKijl7CPG1pBORFn36NkIrcIK
h7m34R36Hfk3Iv0fVtz1qiJTdAcB4+ydC/bS7a0K2WI4t4nAFs2pzSDrcUXqJ876
aAA0EWPSH6Niv2d7X77QbQgN+UdKBHYBpWgPmPcpQmB0Vi8U2sx4KaQMY5x/Ck3S
w8Icegfm54kKD/7KSWUqWLNj8dOPb3qDsMi3EvLGkXtojTqc39rV9W5XSYQyztr+
v40WuGGG14G0/dvEJ6ts14BwlJxQpPmVS7tdVrOI7Q/2WWGM0mqJgLWTzSIL6kAi
7zMpyAOwvIdHotHWc+cMyhYFiFnaILVhov0/VtypMbupy3xwuJ00o+Kx7sz8KU6+
BgCG35SJ28THJB9b115s26x1u/8N8mLjr4VY6VxnhkXlg8Q3Qw7CACmyCVqT3KHJ
uE4HVPf7kt9usSUoyuLLzaGjO0br7DB0N6aFLgEohoUWFObXtYV5ZCQ0l4YJmyL4
WKUWMolkPGgbCQ+TpujED+BlKH3knYx/1HJI2yt9AwmXn8kooFHtQyvY9p6rCMur
zlryqxtsa2d6dkvRl4nBY1po17R+8n1GmBGunXjcbNuacypVQeO0wOo+p9Rg0zVd
8a6UvSswsJzMlD/IxC+eYG6/KVHScqydmQB8uVB/uoL33OO4JEgWH9uK8tWip1QX
UR+H+pp7uw2rmCfSsJRIzGziSxZkwQvl7k1iu26Zm51FBB8Zq/OLoGFXGxsXr60i
CaY9cVjLT9AJX1INP+J6tBtb1yKD+CKntatS13t+fx3bDjqNBueX6m5XUiS94fwl
sIvMhdLJ9xpVdcxYGTYzH3DVBiPQ4kKv7vYdZPwF3Smf12fhuxhhVsn5yA3eK/vr
MYrZWre9rBPne7ohPjveQlQqO3C30fROKuhK05rDtxcFtN3SjfQRjqDOgwV5/joy
lrx3g5t5ed7SK6tfOBvR6FDnIPvkmeByuf6vC9iMsV8pgdy8zID4kLf/A6igF0OC
UaTX3vSdMokFhU+KrbBiUmwoRddGpyXRjR7FqxwJtwuVpeNxT+1h4/BcqZTPVshM
zlZ7Mbu3GeX1UT3K4VRsP/41uhPob7goVOtKFYMeerYecXOmCiOwm/WtCsw667hZ
uGS6gV3PUDsd3AB788Y3L7AfyUCQ32aGUdwRfm5hh4Ss9JF+z55gUs8ItJ6pyI/C
an37ZvO61gwkmCqGv8Xym/hUkBTDIu3BNK/lDglN0DymO6swsv679aWGbsqC+wyT
3IIgWw/RN8xCYiiAWtJnXcw6V4Mjm0sdC9VmjUZSBkuUGCBmY8sXEk3NRt4oZclb
4nKT6QiW829BTCa0p45Rh5GikOUPvpLe524HzZ9OYCdTyboniMPBq7bLKQGM0pvn
s4pl2Np63ZTfXf/g8Xfm0K8k/lPpXyqnudcUYo1yvCkah/SdPlmE1GMH7h+iLSaF
1pGR81Bj3Xt6ef1WTCSUL4CxLo2ohx5ldadC0ECoXgwg0nPYYj5D9kG0g/nojYib
I3U2tooEo+mQfsTBmKriMahBnHvyx4epUzyXHcYWO5Am4EQBnP5tZkTw8QVzoSI3
jX0b+td6ZIDOzX9690vWdDRdqjHmlOiG4I5euTjCTNOcVEM5/avGnz/QjeAtJxWe
WQIwihI7Wx2ccLhzJvzgvd/putmy7wHWuMcMzeWkMIldOm2IeeuONToqi6gTv2v7
VVL9Mtya5zI0mvEJl0IRNkNQ2bCbZYZ8Y9xSrlwW/aEBodhN454ESixQAPBmCTZ3
YY4mtZuQxKikT59+BpfZOjhX4BDv7NBYAR2vU4BsU+BbKeZioQkytP9hObX2IHDP
Nkb4TCAw3FOSC5Zii0VdbK5Pfq4VhZYJbw2A7qYQTPiOW6sJTiA/FDz3u3sdq/AQ
4diys5AFsS/7rXzWYINrEDieuCsyhjU4OFl+wbha1mdNgW7w5ZaFXPqjHPRqV5cH
ctxiq31Upkx71vBhqGQspwEHAcWXTHSG3csBS04d+cIdF6L3kd+QoAExo1VkGBZk
P3juVUWJAmiztOmA7TR2eVPW2+iW+OeGePb7r6RRVVSN2HPaR3q9irXAXrLjby2+
AxCd5bI2HCkmvCZayUUTHGa2d1IHWhY6vfRWxq42ZVRY9azZFYhRTmOwlkmEwaAt
S3WSa/+2UsUYn/u4/Ir0mhNWClYt/4+BSyB18lRLewa4mNRUf2BEf2vmgPp13OjF
yRm8aQsDbVyJ+SbS8+5SD+Xo9Bk0Cx7nygWg0irOg3smgGMyiCpcO8L58aC8yCPi
tJsLnfyMAlgQOzYJ2r9RI1UNRu/8SkR9RzOd5wLwFPXk6ExIsMxCQ/p8mvy/oBX3
I2zbZJAWEMbukHvdPI00nG1byykWc8W73Z7CuMZv8mivhy9y8bvVPUdEP/KddiPZ
fzzZowN6F0PfuwIqOu3YmSd1Lct+2TV1qV39kz7WDqScqxWsb7DgcuWnok/67IMr
WjXmQ1hlAdjuCzY8j+gDX531euLLF9UdWSjvAXevjHtJ6HmnNOaktLqn0iNcJvFW
gA3jHPqodxpUd7PFeMUg7hStLd6GYNMdioQm2IIXNV9XwlzD1aYUce445L61UV7M
BSp+rMdnC5GoeNPaa9uclkqy7b4PrJ9MyELNPiF3h0mKAENCesXwzXNhHW2+SHKE
pgppsEgdibVDM+1Ox8zE8d98hVFoyl0COx+HtvV72TDm9oTYSREKNtQtGmZrGCpP
gR9D04bs9mRWRYuFaY58oELrpNmfB2A5Niuw7z4dVzOc3NTJ8lEfNbV8SmRBRtwc
RlUTpMOpgOyhIx41Jxmid4vhy3NUXZFfpyW899chBHL2zWItVNNW+0hWuxV+P/RA
d6HwGJam/6FF5ndOQZ3/9f8i0Wb/FvSxBX+7PxMtz50gHGLeGKJrrKHia7gvx0a6
ICLYMPTaa1zzgzF6FhVvfvLMxnN1g8/PsiBVUnKbjuUlW8HhxP1gkrZhbUT0YLqA
WhuR04A1dVi+o3rJuWi7C0gG0JbYu6AE8N208Mmi3T8Q8NSHKxyIR2xzCQ0dpvQD
70tTvVWOkQrUH8PArnNBqu9zD4Asx4ehsFmKJxcPn5X75D72D4W3DLVECuegllWh
UpU7Iul1TeF/1tsAfvD7yThqrXktPCn6rsM8/VmHpGZo4gDEmfL0l+bh85jz++fl
WcEOEzss2JbvXP8bs4pdDdL8fQr0dwTAI7XYj9gncDBopkwSBK073cAri0Xx4pKW
deZhN3x/l+aqWfUFu3gELQzknB0AMeLlCSq2gKQFeeyCFA5EHetbetPLUFG6GxT2
MIa1RO/XKn6ebC/OCEgoLGJARGKxAjo6afxvg/TzgX6Nha61wQfpi7f0vX2bL7XB
NDQuGgjmE6mWwwqJg/2sRnj/qq2Ai30oY7YU5vufEPAgsMCtn09HiA2dDgHQ+rbB
h4WSa6FfyMVZcd6n5d/wuk89AdW3NvOMiaPDjzAnXZs/GGpZmb2htgBhbQK6aSkh
+URsL1aoUPjrte5DtriIn8okvjmVfJV7Rbb4iN9GVRzW8iTb2GIkTq8Ukhq4g+n/
va16X1ebDStzrrJUhzB2DzFmlFslNlNq1jFni0FZ37xUt2ejmG1pIgJ9MzMNmq8T
CfkvvyYkk/n6QoYtBEmlm29iU4vXR1YZDStcQMLxo7ZCWnRWlh8oCH+gtSZfMeMq
YVxw2QaLqo753Z4P90uSaBGKiIKf94jZNxbEdk6Ti/v9H7MYjY6jQbmo/ktKok16
fOmsqTNnPsx+B0tdV2NFa32zbgIS3+T8JacWeX3PPw/scQbUKHrMVSew7IluT2x+
omDD7ydCK5jDkDgSTUYjibKluX/HqQdw/K+ATwKhG+2qAA3zNZlMjySDjZ31nrU8
JFtN2EtVHd8I3g7m6ju1rCe61UwpwuoOHLyfpeEF2UuPKQwocUoigY2Tr+bzlAnK
xQimO8ZKhd3Lomg80qWyKIUT/ewSUkHM7hCnW6DPvk6bn/BRWqKmknzbMyYBUjui
Tohz/+o3hj8NLs4WqAMZPCNx/L5yrx/dmkJR3yNurWVsjrxGyuvX6jk7JOMfi/X9
C/iGQJpkQ6IoLVNuxEoauhass2rLdH1abapkxNkn6m66C6abO51ZtgKPDNssHdMC
hU/uHZ/veNIsah3w0vXqjplj00m1j7+rup4SmjEavGIxmFg/Q+w0Fgok5d7I6QKH
koCGKVq2EslKIJYuUGs8Lh38jRaXEt1Vj+fcFAHDk1x0t6PTuQB0RrHfIgn1fr32
xu6zCiqoH1mgQnV8A9E7DIQ07SHC4bvTNEKptvmRktaQaMLd2SK08D+MVfeuO+Wp
I7l03xwmLitC+5Sc10VgOC0NVOrTPpaxLe5FccxyoafD+kfFlXkut5pYqdhBxvuv
fApSxGQXmNY3zCrkLMZvUB6IiVy/0/ooprg369b8aH0cg81q/LTILtSowKaOy06m
48DZY+cAABbkhMnusj6FXy6RBcAyUtpYNVrB/s4XkmFOmFEKbGTfYhitdPuaYy9a
kC6GvL5FIEwy4wj84B+DGU2LIDSEmXv4CEU9s861xcHbhED3LbwBvuBAabyQ7lzV
SvHDPgQAz5DmLDzhqEYZ5fqsa8ImSw8qdtQOLF/Y6RhTBQ/n5VjFyIexjC7T8DSu
e/QTQ68d/YX+91xz4CYqGCVuldWb5xerfrKwbo8EgV3amndgVaHRM6qh3FMh/dLJ
1O7kt3rfoCvlIqwpItZjEPN/DaqGGviQIUL007BSxkREoB8xddwwmWm/KKROHHdS
P7VuKJ60Qy7Q7CBvWrcuVrB+FEx3MtevHSiiUzAK7B/8ILgtSWFnL7E+qoWB0uBi
Rk2oOdDk8gZlTlMhj5n218OaEyJnB9HCvbOnvkz8ywGQSVwGOhcgbt51AQDZiiQ7
jKoWCSGYzVWg070MS0okTkBTUMSzAVL5errWxdBImwWsr6NbfuRYQojztMO9VWGP
xWfQnp/STjN2BrY0mqykUqHirommPQ064f/qw1NryoYaof3KunjYvNInFAu2gH6x
TPB02SN2S3Ucxyjf/u86MdqjOW2JeiCsKUbwgX+Oxy/N+IdilHfR52MeYg+30t4a
ufxq0+YkG2ftMbDR6+JP4J76ENaMSB8ECWbSfG1SskhwZlCQvf6sFDOedCKsmI8/
cjAinE5XyyT9RZ3YTuk16umbEvO6ZEaG+u1lmkAhoOI6UbwlFZB5qS94ZkaaC4Rp
+kQ4OG9xdLXuAsaMMpk9A7lYWYBZArw2CYCiJsv+beuPu4iedvPyw4ZlrZ7PJ9jy
tTxh7ia01+/yGAg14sx3gZfGqnnOfJSREnD9XqKGFuGce4bbztGkxegN8N8bMeek
8gySg+zll2wIAbsdplrI38uIKcDEUY+eeIf78B1kRDqMR9+XUMGysUqWYJrWrk42
r5dtNgseGLzksrKJCNh4cuDVw/1dcJrZ8HhF0qj1S0q54BVa09migBBEdcxfDpj4
pF+juR9QEg6fGSAcu1Ff4nUsxOmeXLjZUJq5A6KkTg62Uvv5HsYCJcXi76cmkZzT
Evx4dUFoC7AWr2Zk+A7KgTSHXxKdyBkwUFIHue8fYO7xvPdLb03dRQ69I112kG54
j+yjWijNjbmUSvdllUY10fdEKABofskULQiXym9ZX9h7Prz09ltValdI88LYvTBQ
FvADARZqv9QImJgylx1qzTxebS7VdQC9/V3j3xFsAYlaxuTTYRY8KJYZviFXk9mm
wpWzcWk/qbqBraHbaDOl8lfEsQbFEAlD0wGw2ZW3nVuTojOoLZQ8t5SMCVm21S10
3thWZyIparYw6At13CIHVI9iGjvCxJGlI1kUV7gYDltCNrQfAVx8qUkjvbH0GyIH
Wf8Qm46I57UX7iG6K8faAELrI5vRaBjpNKem70nS/YihsjanNY7JADugVbCY0C3L
1vW0eBauM/sr5lyEexe/5xHB/vSaNHDfAsJ7zVCdGZ0ysERwwZKO58FkVTucnlUT
spdS72C7HGmJ40RqzYNJuxibo15WZIfSL1WDH9GbQ7D8BRNRbvL8NKFK8K4saRvm
8PsE5+kk0czqr0CzSpt2yGcLIC+jr+wuEDWVp5cm9PSmUlYS276iOjZw4uqmJzoz
lgnZJ2232tQochIPmF34FVj1Mog9ii5j/mjpkhXaG19cM9252vNanVhpSlFURpiG
X5fu9xMLJ5LIxAEgEiG3Ha8aKH7Ssjp89TiP/bipdGacSInVX3VUBonC4MA7t4/c
/NEQijGR1zQ0zi7soWpQWcF5r1FhrTMlHLhlLlwg8aK+EVHifc5vkgwiG0Vg2HII
1D2zkJJm4yZG7DhPdLAq0QDCFzPjoeEDigNObzSdi08atqE8Y9GsiAVEB1U4FqE0
1QrCGAVjpIUvEPvgOv8G3AsBFLwkJKGNp0+rIvyf3Wra+trtIO065pekUtBud4Jy
bgp9G5Y5BptArXJgK7/56hY11jlPpu86TFJkUjuEhvERvmJHyrYTVN1P4IS/24Vz
o6oWsMsIL8tsQDcick+uIKbEkbxjGS9F0iaFl/Nm5cg+VrKbUF3Ss8RrTOBL5z1q
e3Xo66ev84mYhVEYF7isxqAXq6IJ8lQ6WWxRswDqJW+r7meZSqB8RtXPf4qwlH92
vdDicI3SeBkdxhRRW0ef5IVmtFcmflNB1qU8T6tlJsLSSaeC2v0xgk573F+VBYsd
vhpTr5ZOghfmOxHewYg3hXVQnb7xTOYi9qRf3ufdM/9p5abDTPHMhFpu3VA8Tszz
FuCzOUpX234JM/s/VUL8BwrpKW5a7RJhzGY7dv7ocUHcj2I2A67oCMIrB/V+bFDZ
rohdLZXj0Nr+RPqWdYFw4OBC8ttBtp28CGZo4U+zVDHopFZm0pq8MLw8y4HWB6JO
WgRGj6fyhE61ZEp5emVwl67GJmxsFaCnTAllsj0swZVGbcriRm5OvaKKFfMOw9L7
E259NctOsxaVo1Cl8tDGMNS+sFrrgAf8CuXwxB6maGNuRRXJOmBByInEc66fxIxw
Wq7WGLlKvfflz8tGbpBZEkt6jCwXrAfEBf3thbIHlH0QbJIuezCiqc2hCKDc8y20
8mqqG9aGL43wvEJrvfdQGm7h5Ks+irajv6/Zk8DmaMSl+xMIOoZrDjSsxDC0qnI+
t/0NJS7mfZAu1A90E23qLm66N+geP3XGBbcJGui1m16lMJhqrq9CxCJmmgeswksg
Ue3mNtgAAlsv/OumnnSetAj+WFbBqM7HyKW2PaiwE2cS4iuvY3dF5todhZULMfmw
rcF5suW/HGBft0Z9W+KQqLjyRtq/ZMgkh4CUqRUm9tzd1E0BahPQpPqIo5KDzv+Z
hnSrmTedJrnDcMWqdDpX2kJsB3MXStRef5GVmhUqr5LQvLiVtpofuySTpkBMoEv2
wDJsb+gUQbJ6FkoSCC5vPDX2WIJ5aWLLj8YFS7thjPI2NeQDR8txAnYTrbdemFtU
YzExjuVmT4N4zv9Ar6eeE/E0Wg2YR5QsnDLy608ZzklWhWGGQKbkUUr8RFVoVQAx
nz4FSvxnNf5mKAkVilRVytxb8DJ21g8BJe5+bO7nSX6kW5GFPEBDRZxRzaimEN1i
1ACfRMwHshjmBH+mrSNRvJZOkyCGiBiO7uz7vdU1hxWnj1lJKs34oozizU7b2/kb
rdsW7jJlTCoFitKggaSmGlOMtgOxlpe5/0AobAX0bpOexEGKKUAQkW2EsE/Ptxrc
YYB9YMf8ja7O115uV0D8e1sgV8aApxRAhqg6YSAsiGyWhh3YwU2I/SHM+eo8Jg4i
XU5qEwyP3fT2zPRiVDX9Dk0HWuAwZNvJKDZwTcWgFCw5eureyL8ePqIzB9M8CKyW
Xpoeh53HgbEtuuOai5fcxcHR5wpqnjDwvPg5ObUFob+SOClG9rFcJ9pimGtIMU94
Gpl59GW/bOsm7wTxUaNQWFRwWgpHDerlqeYHET1y+7hl3lm1qJ5XvFnBkhWrdXKS
U3cPaIcg1ssNKd3gqg174k91lKsc4LSv4ovtNaLG16jPSvnmhvmeGi7O8PwQ0UjP
/Qn0D2vrrWs591nnWBHPZrraFJ4otsSu6FW6jk9aXPsfQFbS0dGGp/DuboVB51ru
zLJ4LBp4tnQd9elA/J8HzggjgiMcZ7/79wcAB61hhpYjPWY4UzZ1LgLNi5eyVvbg
DOaTISF9OGtEhEXLfDY7vLxBD0B+B9SLYAIraqMoFx1teIIPC3hNWEbevnjjaNor
8CwNE42tkT1mC4WXtcUMY2F4RNZIKD0010CwsNjRVaGDcm0RmjaD/YmJ4fbjW+dH
jVbjIGfHZj2s8ZwrIFz/093EfjIzdWsmjm0slfXESrDuMJnG3WVZIzOIcf5EFBA7
J+MpSAVrH831sO5/huZKpvZW4crhXL+Kd3f763ql8EC/9S4v2+IC7p5fk+hww2il
fD45JaZBknpuwOBrw8AoroBZkSLmhZ0UTok9pMcjs8eu1URrDglUMinXeplrm++T
+OgAhYLQLLuYqSDdWxvzpMUk2Z9JSVLyJcv+jYNWC0sSL+52GrKNRlFU2a9pzFT1
Vubb2zFri+59U3ss1bf9blSjMxLWBZfwnUX2OgGXOjFRnSukEa8KmdLSGJy2HNrw
WReqQ1qfgsT0iuZKyo9JQJUedz2YVhKzUBvkKzSmNSULIVo9MveBPJkclvIbuyQ4
tduPOuZu4qjTn4mp6dRmtbHTxI58Q++ZHe/wjxqD49yAwrpmqxwiIAeo1OokSCy0
/gcUjD7aAO8H3x6Y8BOvNaodWWpBCr/5nJA1rnCyHwhRL2ANpHdWPDdVqE9n/5Yj
gCCnmIzm5FJxsIh+ptKqMIOx+CLCryUWJCbYm7kQMjK+U0E0snArAVsdpykGWxyE
o/p3A9jgmprOR0cRbfpXb/lrkTi1REeDoVwxdyuXRcE/0cQ0VVoLbDgAisK1j+wR
Uw/9pMPmO1Txg+xAp357gmMorpNF68+QN1iSYl+1msAsfxV77rz8oVM6T9/dpANc
o9sWcc8Gx8bLL8a4xhOaYvRJELA7+dufedLiy49q1N1NcagjAxvadpXHE/Pv6FHZ
N0ygw9WoaVADnOMLKXlJBkMRnHFxFS93DcfDvJJfEAejTXn1/S4UGUuHJkp6Ew6e
emkNlJeT38zAamanSrIIdEGOhHZWx7s+AY8iY2envKyO91+Rzsyjd6FPdSoodBc5
KSgOsFEjB06sFETLmr/HeEYkEMhedce1sl/XxCDhdrcDdbFrvZWKzR7FHhLVU9jW
CC3P9pORPgZL1dOc+8CbZFiteHTUIU1rt0tzGVCb+iNPfeYgGK14n029T20HadYF
ItfSrczyacXyz2iZF2wdJRQGZ80tKk5Ug8eY6yWWXi+C2JX7HVuPV+fHP2xaIw1s
BW5+mMUqClrwKqBbYSnBtKZAlKJfvHrxGBTHcNoiog/aUmYKsrFdEY025QN8CBkQ
WL7TDDZcqw+WMOmkTHABz7f54sTCjCHSGQTDhtEOnIw6ZpbYeUZKjnCehq0+Uxo3
CDEGt6/tAo2rhO2SI2Crz/YDFT2SVHyEExttakUn11e5wYtjInclxoDOGEkqG15w
uwN9R87aWwruKIHK7m7hLfo6YGJvzdBnVwvOLuf0eFYvFQG3CZRGdKnX9y6+wzjw
R2f5qEQhaxnLMZB8fCzU9qdXs5tvP+qf7HBsYXKN/FfkZvULXobT9yD5+LYtP8c1
oeaD16biCuUmuxJYiXD+LeTEvYYP1EyO9h3WelabjIRNxAmxkjl2cU+SJkvKKMvu
ORN8PEUNPQyoDJ9+HaiEt3XtVtcQHFBZPenmvLWMEHG5WLA7PZP0GYR8PKju2fWq
EbcU4xvlaPxU7dJQUnYFK8LEvu/PrwbPAScCohARCNMXplQr2zXMk4GJs7p/2f2r
zxo9LfqMZsi5gnAlvvEMRgZwrcFsaCnN/CydYLXP7gF3cfhCpBsKNerdpbgNMbmc
CpwR4pPIFM9Uuq1zdrir4LxC+tPSyD3iCvnz5W0fmHXHDMcXpiI74KwDql2JNhxh
BlNI2fkQmaeSYkPDASy0e3cTmcrXFtwpn5fbkcHTZ5vM/YlbMGesLDmXA0d2bw1S
C/Jn1C70/K+LA79s/FO67e+r9UnX1BTo75Pll94Icqktz17TnbwZBdWBqYfsft66
Qryv9AJPRGNK+b8Z4GlsP6nFu2XURc6sohkV0OW80wQ6UAyutQIlsFxsXF9G9m5N
zddRf+ib+igtnamBiOLyo9GqIEpGMGHRTgfJMrtO6lQ3LEdVn3iJ/xy58/P6ITPW
rfdKXAM3fpoDvy6PAzUgMH3rqlVf8QVY6FjMGxJghlDDpV3n2UeKJQghOrxaBJ2X
HCmTkC3OjONPi7ffiPq3mOe/R4mqyTVX4ly7aVfwku8B+CLjkoCPKeaKCVQ0aYXn
WduGEUFi5jB3I8z3cUtyvErBniGEYEKed/Sfbk/GNgdWRixb6Ooblrxf0d9exp6D
J2i7NIsf5He5dYccmDlnDsskYkmVXdjNIN/gBdwI1phFdhli3S2qXS5+hTCXSWuK
XsDKGLbFbSartymC744Fggwkbo7443mgyk0MVB48s2xLcddrNeC0byB4CfAOXfsM
kYvWWKmvNoKGkboBdLoBW31aMZC/s9H9pf1l5JM7P91MlPuJlM9sb2lGxp5wRpji
LjjqgFgkwYJdyRC8NsTDxsCIg0Ix1Bztx/Yo9XGEXWgf/spTrqa/s7x/QCWWMX0l
Z5nLcJZ/rB1+QqL//Igsa6abuZgB8FlIc7WZogrEPtTgtgtoMNwZiZ60lfsm+307
xzCSgkBiGSgXqWiVg/9elIuifFtoQ9S1Htamx+IaPYt/S+1V6xn7Xm3oUE6TJZrw
kQQFWTHQmueVYjQCba7aHBaC8uW+sHYXcEO2kEaRGfbPKKUocpaC88oIVKhO8p2n
8tGt/KE/7ca0wMnS8yml0Muo+1WgS+eJz8vEjcbM3nGSc3oFWQHpP1uoG64mjI3X
r/pf/My6QLt/HLGM/4NuXu590qeVC6q6fVVw2YfdRWURJveHbDo2KROl2BnsG7jy
HuzMNZZAjHIYG65aTiagHCLrolBmytbgoBUfWLR9FXLeExAqEHtXhvjo+3CcXMKF
ANDPBLlHSx3TjTbtd6Ggm/xR03CH6DXioV911PB3OLZ8rVp/1ozOwymcPVEe01U0
cg5tOGByUf3guHZODehnezQMBsQcH7tQ4l+2JQj/qDdObqWKfGsdK4BGnZqe8vgC
QCGlAxNho1Yh0Fiqg5vzZPpA6tbUrzywsYL06y0uylYKj5wvsP3WFIYGkn5Cah9E
b1ct7TaUP+zwrjs1WUZuM45VrBCn2BE32Maj1JTu48gth8b/kN/mcAB3OUC5GWOV
OPuBSa36lWxerjsSpZBo+4I7D2gyjEcZ3UChruPzHcitlutlwBtVicbPHUBz4n8u
kJTBPeoP0mlQPWcXQIci0xFU5EFDlnnGOKDtvVajPBSWfGx4UTU48ZbMcRz2x7d+
BRRYj7N4iVAWoMPKoTwcueS7kbSUJHjvUaSggaBuuRwx4IIj1VuJgvbJsKABHMpD
AB6ir3zj49b8IOOwDWZhkehTivWvCtUjN83JzBVOdc8B5eaS3aNu0V7zga3o0XNv
djA6SQSpT1R3hvGfl/hPak0rGMTcZyVVFCbVkhzVOifdHM5518qcHyjriT8RaKL8
ZrjEaGe1zGzALVw+AblR9sGTqJoxawBNJiRG6OVsQyUiyQCCiwPMG6rUZxlCsEqR
JudNOTn0cr7I0mxZEaKff5EWEhk0BX9Z2Wm3wmEWSL3OlH6G4E/Uqn4EVqV6dMZS
7WvcpG2swSdJ4/Kb8XsoFcTeeWvc5wwbsIXOc/tOlUZXVHMJik52TfOMe9T+ov05
Uc5q0Uei1wL+7qKAgnFjE/YlqFJSC/Wq6mEYnqACqyFzzHxE4Io9Yyr+viFrNR+m
Df+te7do6RQLvHmU/4/oSDrVrzSIMkahwWYzByTxxI+jxbSbWTYnbT3h0wuUHFyB
gP17tvFVlxp78qmSBTcBbvdjtw89V3kdukgQb+GOV+itCWX5uxt0KRzP09rMv3YG
HVDDBNC9dKgeksXbGC3250fd3mX1pUX2+vj9OGb+D8B2QV6xH/g2KGDQEZ2DjnHA
Eh0zPEfbYcRrpmFH4ivvSuY9USVhTD2GMhRJCaxXlcY2l27dJvO53NhRsSWvdJ88
3kKFvHj7e1MHXvvnorc93IGo0qYziAC64e0fcCIcoxz39xJ9n1fUtRXNlfvHUwHm
f1AdNBVgeQH70M6Qdtsy/a3LuF0DE10b2C87IbYWQtbmTK/9UFqQ9wFlJ47+kIMK
r+QTZNvSXB1D7dXJvaFpF60qGakKoIL9TlfyP/y6/RtdqVQhfv6jahsc4xZm87d9
ab3E2KmWxxoikzDxVzCwU6Ycdd4ASTG+u+PySMYbnUB1lXy47HmL0wd3zv1o0752
0pUqup5oiMwLrK77gB1JWr1KItUdta814fcaxUEBYWi+5jd9lQbw5rIapx/U8lPE
GN/K+/bUx5nofT4CK69UgGz9ZcwXeO3t4C0EbvQOA7LVLF3MHWWYPhH0CXoow9Ld
ficLwmDx0ErBSlAgUZku2xM+aMSymjyf8s15TUsp9B/p4B8fCrwtopp69PPU0IIP
AFSCwiuaeFnGqwWdWAkX4nfYaAqumFegu29q6TUF/cetiRi3vQIHmp3q45gZgQJW
pAx99O3egZioyCHP9PjOMsyrNREmw9c7BGiA2pJB8rqwrBWc0yPcCN1gBeLlllP4
Dn1JKKSFop5GMROjxJTtr1P5tG7qD0PyNta3u3zreL5I4WGx/9A8RWpwxQjoR+b6
Vx/m4mE4v8a7pm/GMQRdeUFwc5mi4k1KKJw7hb5xFar2EcDtEBdMIOROL0pgVZ+9
TAi9mcBxQOleOHBxv4niXEZTEMIyQZDevlhtbJjU+g/03qY/ktqqDGuqVIhnE2Lb
/UtZKuy5mEKdN1QNpLCHsH6VQB57ADFPNe5VfnXTBfhhK287OL29M2aHzNRyaj7U
cxdeFrB4TIj6oyT8xE/VYPwZiPWvjgiTjxg2pgbYrEvhKiv/sK4ndmZWNJ9m01Id
pbaIfHqrVCmCJEJArSeEUgM1tAX+tgfB8h7jtw3OZVxanwRA1eO5O4MxAI82gcrO
uGXOy9FOJ/fbZ9RoMmT35OnmFQvHgDv+9rYBhjQf6JGZidwPtW1JH7ESrj5RPWFh
laQQuEJIc6yV3TTnyREhfWXSCMDva73UDa618aim7sJ3PeUo6PLMyU+tiR2hp4fX
SEs1ajZS//oJR53llNPjZEMvrGWHVdIh/MqmpNEl6A14XJjbzlacA/sLGxeZ/kFQ
iwUjKi+6vyD08CLmIFkxSDulBtjRAef1IQo80pntKWZQt1thnj/6GPbco5NwMpvz
9CZdZmMe/KMTHwrwc/hAoa++NNSzwqHsEqIaeet3AiMWDhdi3pHQCxbsjwTZ+PPA
dKEKNkWJS8qVw25qsooFox4Mu1PR2ogr+0wFlGAAQ7dh20GTrG0XkLLNy5J/IgcJ
/WDGDp/i1rbuQXLj9cSQwm37h4mnye5cIU8yHNOuwBhhf/cUC/B7kqHqYt7SqUl1
dle9wU2N4ura4RcvH7BHBhyNXVaTzjqe95jFiH7ggumeDtaAbNHlDFH1yo0B7dYq
ZG/beQgz8CI3/BB1ZvWPCjNUC2hXf4SCADdRBZowNb39jfAVwE8xeE8xQSzNQ6Uc
fRPXQDeEXm3JvIRE5l5go+eX80TO0ieZHII8cum00fCqs6l9IlYm2rt+JhYfvs6v
Nre7OZ/n9rIfA2+Hp/y9v7ChRUlgWKmYbU/Omd1vOOYS7qtxsZferpDDn/jhBurQ
eZDncy0ySJ1Zxl/2IeqYTfaIPiT+plBx0qT1C8KYim75rxWbznudc2DBlqu06UY7
ht04P3QyqxepfUx9S7YsI4Qt3Z/Q+VMRUSAykuYF3KxbQ+BmxM/FZHbOd2dVecAH
MHeF7au/L5x+e1tCP1QCIP3H8ah8Yins7yq3Tc04vIJNgmypuerPthQZjTQHrib4
RKhhYvyjNhU2j8JqlcYrqU1LdL/Usi3i4TaP40fsMc7uKx+owNv/NP3nlditsdDl
mm8OuNB6IsXbUK1+cxP97vlwuz+1F7dZfapx/q+UMbVJktW8/VSnDo58Usg4HZUS
Vx6kCAMn8cVfSZ4/iHUcCfLUOymINQpHXZWg7jdvTbyK/Ml9Ro017bw6qhF22jSE
/MxKUa959/MZLSYwpbf+4jjYYYgBXLGFF8wTutMbFWxL8kLm4pKx072aw5gZd4dg
Pgp1wuEeEOUS7aHVxhWEo/mqIDjAHmL1p79CCLjW+p2o7RPNuiUVdnWP7dlwy8Qi
05JQAe0BCdzH55DVkMqcfNIRf14464xbc17emvhTay36c8o3PWy5QlqtaOhZzzL7
ZfmkcEAao8Z97Jacx6qUSf+CY6An65H2zdLc3wt725StKEoyLNs32Hwb72SBdfgw
ARlh3G/va8tZ44wQf18REPOUv0i4hlZFaW8QrpRBdlEKvwtpeHTRKqnsV7tFu/4H
d36VozyxuQPTAePIqKZgNs3OEKq8sShKBeri+dj/mW6jg5YuQmQY8n74mUUIZD0j
jvv075fSrDgKXffrBBNvYKocyKfNbpNFuTqz5jzb7hgL+lbOcVTspNMRpk99+WJc
dgOlDDlQRb0m+1Hx0fIBKufe6Q/9EVFxoErcIhO9pOqKJ1zPGh0cAxp3bjsLxQ9S
bqHKjn14bNYqEK8GSRe1JxSewtoX/p0qZgeFMytBC/vEI5P5vG2yzvWERppxH/e6
gX/LzUCehI63lAZyr+YPew1R3R8SLqf77fuu+LvwH6Fxch+dji17BPqKGxCcxqT4
GNnD0VTZNsFQqfXT/dVj7SrKp4TphDrp4RfZJWlUnBhs2WrsEbNFEautoxalN7Hi
AC42tR+oXKBTkOXKg+s5BAMqEMalnryIOv2jBOXC04co/uqOnifL3OlIf0ZgqqJg
+MSR9WIRyfdQNzyhtiMgeI8ZjiVDk37BZmMBcRZEIookn4NowfsiXTgdT/Jzg6n5
M64kqpVZswfySY3adPuHg71Ds7lY1AUfGwz+cJfHU5ZeX8DERuy8eGHvcvyB/2ea
wxFoitN0i36J1ZAXV7CoSlXQALSkBgJueOnf9C+i53XCqzH5xKqS+uh9fOr3HXH3
eq0l60Dv+KNox6yzc9q9JzmN83iB5m5Qt9xoxpb0a/YPTCaDEBp6LENN3vAQOX/5
vNZ2mQ9oyMtGYwWXi08ixwmvD4ueW3EK4iJLtMjqhBBS7TKES89rjQPqRMQBNtJE
zg946m+vI3crU7QR5l7/0aFrFBQxYHy9WXyzZxpvFoswegPNDcLJf0AvQQQDJr30
BizI0H+kxJpTTfHkyyY5xgBPwwxk7fFfd9YhXFKuYn7WrwNZ4h7284mVNz0p5cC0
GJ1erSUhDUw2UEyMpG42Kn+RyJjbqMxcckAn+Z1usq6jCHAPjQkWZHVISrqtXYoe
ODH/Em/maI2UJRLEQikhPMiokoLbGdQ0b24oNww1w3GxgIG+8ZJW/d3c/P7zbblr
JY/vUW343IHi7NICOYI5OBNWzZvXbJrBs6+8mYQPjD9rJpU7X7i+ZOyR20CpJLqQ
8Mm+nIx37NTDca0flkU2fvDMdjMbttfuZuDp7kbDu8GOD5v3OVGqEvmeoYfA6UR4
mQytQ1Z2W9PIk1TqLXrQq/D83hzKQswpL1yhg5yacMprnaZFu0GAdGrTXAl2P81t
4Sq1u4fVxCXLVQ9dARmZuvRo5ckoq9XCn/Id1YKmcqYdBPaXjlDpXEn6jSNANLgY
RrTpOLUJFeaeVOLBIo+ls8ADiGWOaHOeKVdu8p21Lnj/3KTMOqh9Kn8TR7tGIGwy
uDAE8m7/sD0fDvyVXGq885ZeyaI/Ni+UXUf4KVxu1IjooVo20bMekAZd3e/HHXew
APF8jqN3ZN3gg/UZ8qt3wCh1Pddf9aHReafbC3XPRabIpwKx0dN16peUTN6d4bQ+
xOytVPaPXjrpTyDWfvlvfyZT2uhqtYXHSK8rrXxv7XuF4k0Fd0iM0Gl9dihtpi4Q
mQu6YgsBLACYSvmdrNKu8/+q4Q8ZimXhokZQ0CVspswuk9zQbHigjaBAanMuMrQV
BneOKaKNM+8f089Oe4UQM+oi9xRE23adrdOL+cRyk6sT4fDvMaIFw2IddPvWeXvX
uzeN66ISAEdZXncsqU3nwkHQX/66wxTWx1zFCSl5WxlcHYncTiQ4dy81HjGnyYNe
9qQzZJjbTBW20n6Wc3JPqybbHNdqNWxMovSfMlwO6ZW64sU5YpErJwBplnsZ5v0Y
dstieMlXoLCT0B2JkuOU/ByXNQcX0VbbTQVjw5YuobItd3dT7G//Har9x/iHiVTI
ao4bLFT/F4xlbnnbGbJuf49QS30RmhCAr8q3zyb0nB7btX23rjAtI/nC00vtI6NP
tdX0J7C09A+hXnD/IfQNyDjk0FXBI+08OFFoRAdM94joyJjt45rHQRtSQSkI3t32
9HlXcWz1QogM0VtjdbRsF9X/WmR0/QK6UJ1jfTdzI9bG/1JIV+5rut/YdFBtIkgj
SERuXqk+3KLko7VNOBHH1K0nMJxuHl9zMJ7hlVeF3ZRHRBj5yxgyxK3L8bu7tWI8
u6CJwk6c11LRKlmK2eXdey8+vYJdqp45/qMxYHBgcVJ9+UQFyyKfWk9qFiMTBw6v
IEREuFVxAnG9XOrnt2BH2kKVM9lTsjVPmnThmZXELFbBfA+t/Knn8btSqV9Mvevo
9cPfJWAmw+NdONcrDAUNMslZ8MVo1v6W1DiLq5Bn7GrZ3WwdlckIzZ/FDsDUTfj9
uiH7V0uzqWwdAPGNsQIMtlxvmWwMasFfeSgWhYpJ/rIuj26s9LmavrsbeaoXiHdG
nKHyE+rwi1ctax9iOA0nYHUvqL7WUgew/XX1lR91jbX41Yb0qAua3hnI6GGasQ8G
IQI7msiEvzVVxU1Slc84nW0U9Q7Ou5QI4yvMu8OpVGoevywwBSz9W9Q5YH2ce9SX
hrCLKp80yDRzuS/dnJENwm3CxXjkRp86bHoWcuZ2gXvABmE3Fc94X86GXFc924Wn
+E8mnEmcBeMJvOPpRYn6YFhUA5KdaVWuZ5CuykOXZMYXUouy0ovf594MUdX61b+S
+j2kn+G2+5et++a1qxVHZQZ/ePJtB18tZCCs6DoaXkS28Vy+Ecrkx1QlH/mVRea2
fJNZQ/2llWzZ2RaB0WaNvDz9b5zXDcsOJnt1rcpxv6DUGXjZnQ8HSasIGBf5hp4C
9wBDp/+4fyhrjysUMtn8xBWW7KglCAIumYYTAa1ZetairvieFqBQtzyPa9P+Gbjs
R945swIDvMu6k5EQJYTQXG9rTvktuEWJoceuJZ2mI3W/BLmprN57KviSgjxz8e5p
GuBsSeKGnKnXj4LEQqQCRkrb8vn8KHibqFnUtdm+nkoWv+ecJ4YMEdyc3MxtnUK6
ro+NfFWq4tiTMCszuu+oXy+VQORS8CuyWneOETcMZU1ARd0HbzRPKxlFDw88SDUV
RmOMnakNauqVw7J0RnermOSJfwZWzvQ8Rc/PQ7cUTqBKL9Q0lnW4H3a3LG0XpEO7
ekTTzV28Bls2Taz99MAIaBtM/p7SFqpxCEF18igxfwHx0XkH3jeCvXDSz2CKGxPQ
SdrYtcW/+Vyr78Zu26YzV0ybVx30KRFhfB59iXxcbxVCV1XLZd/bdSsitdTp2OkF
XfrGQH+98m9cmjSgn33x58hw/pDYqBmpOcBaJwri5VPcigg5TIrlsC7biUZ2GB8Z
1wef/wOydo4N804yNtXIJPVGygfg6XZRQQ7SCp/TxACVR+RXxFeVGc+7vlwxqyJW
ZK0hQ3W0zw2+N+M4NFGVyLWEvGDFmzrz90RFagI9uvlC8SVSZHs4lYCop4tPtjyd
zAApSx1khtDQWNOAT+n0QHndUP5rQjCHXhFX/Xs2VwQFet4/5b3RhCRt4u0/i/UP
64T+MYztsJaOjJ7/MgCmkSq2cRAVFp18nGiS7WJHY0WSXXGwLE4KoJVhOHrpuvc0
dkDDTzbssTOE3wkLOShkHyGV98x6wEbIsEdwVZmKHsCjlNqy8ycBdJcqlhBpiE+i
mm/OcZ6UCeGkcHFP1rbgSNQvvR+Iy6bzFLMQkgiJgPMR5ryAMErdSi4kqhbR0hBK
WGAO1Y0do+O4Rb2W62ESbwFBGktzYsgb1hf+jKvHG1LMYBgrZhnGc1K2g8g53ABM
7U+EFIPFGyK/7m1tOXsHTiyVFyg4F3ya1/WpOVIXA5KhunVNEWOG90qgHR0ypk9Z
T8F6XbOibuGa1x80tcoeKQ8iSQZ8NAick8F7F6tCBTbqlhU5gmtdj5sKvGL7vcxy
wfcCHTOU8Pu+bjy1ZvUyC0Gz3k5IH5520JEMGK3/LTNdmHA34WsF8TqfzGLgtZB5
n2smb9rkqRUHJiBqLz1X6WKEh9u9czByoSl6zw4LC7l0MnOux6jUHBXlMnTqjoA7
a2E/Fd0tdjJOn1UKBvOhJoygbmBrU0a2HgrXcDc2gE/3v7sPcEEAqK6jZxsL20Jb
zPfYEuIBdASaFaFqS3jj08c+pb6SA/IqWodSa8SiqliX1Qh18H2svVsP8irzLmQR
X5bG6h72RO/R5NbYnb9QnflTUof0vFAzZRYi87tfPFdV6emWviS6hLhf0mH//sZF
abPCFjDhmZ6jzW9RpkwowTUlcbXG8g0KeUK/FViXHR5tWpQZ6HtCbr6vH5vBWwO4
GwVpb3QfwlwmT/+GPgCpUMyT94XfiupzHsLf35Pg7Fmg8NhhAtnHA3uoQtgRLZCG
Y1/GRf7fJpGq4rRpH1l3mNXLhqrL5z4CS95KzKKVj84828dDzxlU9vwE6Dze2nsx
IZNlBAixzhrBx77jtouuaMoHR2phmO+oDf1H4p9v0j6/rtsk/egHe8tR0v0GXctC
HEZecYVVGPw58xZlEGu/OSQTeVCC5tN3qg2ULB+JVQg0dfpGOBujOLkbPoV38v0Z
3Yti0J/XKCFPfp12CrRj/cDQFKrGJK0EWmxFg59gmvjx7SKnNg8jDOGZQfrDsF8j
8H1913rlnEuoSyuPC7wTCz+kktcrHxKjxWe8Q0pIz+hhydreqB/l6GmKXVIGjxpf
iOM4Yn7i7bcMehGaY53jmWX59+/4HEGRd8xBPUmo4uwPfyvJvhn8vvg3fIQZoYwR
bMNZ8KBV4myEUEwAJwLHfns5GjNo4bw90Knh9yDhrzQqyo3l5bJuPrzlZXS1ktvn
DnUXNVkkd3zlQYSWWE88xnQufr9Et2oKcKbyphSg8A1cuPCU/M/6p1b3SefD1Uh8
dYa1ZmTS3toreDtg+rTlWKqz+d7KySpG5vNxPPL2up88YdRXU2CZiveUg1B9BU8b
EKEpTzoYbz1J8REUkhDRARQvXW7RizHc4fvQf8YQ9ehcbgf41u+S3NWYW256aglW
0sXpzHws9Ik8ZCuvZFgkEoYDSp8OlVPwHEVGD/f/4ty+PbToq8VimD5HeWGICpUQ
iOZz1zISunIESap1s+gFjiCpDbubwXHdvnN8K5dBZiJV8APeTM7duFm417zTtCcJ
2kbbILYa9aofHhCw86Tr9ZhnTEhK1hLdWxy/mLTBgvM2hUr0d54jqLbpXqYyI3qP
FxBlYShaGmLfhToX0JymIuJu9oDFNQpAkrCC2HPqEhQgXIPtFwsiLdPEfYvcA1Mu
+y0noQyE96A7ngebe9FwsKl6wXKiwvMidbMqMQY3drnJM1xGeRnlDGDTg7tXH0zd
NcRIjoExMqY/dVA7o0IU04+YLO8XNepFKMACrYE7iWVRTs/spKgmuhBqHQ7d7OHJ
ri14eCajqpxjtbtvAL6exZegW502ijD2cCzKdHzne3kVxjGrbbdOsW8L2uKInYZv
5kYqNlve06Cwr2ooYeONdXq8mGrQtQL5NMhv0HeQmo69nnUAk9mPt5RzbwobvxHq
B30bAEx54fdJGon+VjvCX41PFch1jgcS4+MXf2TQ4LnwHozhM9kSsx/aoMvk8bNy
ZWQsl8zCMcOMByAD2M0WgYLBubJ+n8mcbbHcvZHQT43k36Bxx7HNMRrJ0LqYIVSh
SaIX2nW09WQwhT8sCvCPc6XwIp7DQfyUxmlibbQpEqMv47xRyjp4jPTBcWz4rKcx
wiGHA5f0owvVEUvn8Eqz5RPCbFxORrrL50/DrMavtqPWdmmOIm5A7zq3t1sr3T2e
NwdwAAZGpRdW4laww2QAfcIviA6PlYLTzu0kwpDaSpjEmiFgUtlcelSEb61wfLnV
/V4CFO7n4DivtqwQkeQQFo5NLShpjl0IrVMOFZ6hrRes3hN4PztQ9OujgJ6YGuXm
p9TPzTtdfdHLl+WYycoybpk6T5SSa8Al5/UgG2f7L/ib7mCM8S5nQ0y9ZgZ49Ovt
HE1uTMavsOU+VjzDY/S1YMIjIHhQXss4H7er+CeUuSw2kRgjZeWyGcWktxvwHBji
mu3CefLvxcYDvDpY0uy0E8pkFVVK97vdEVKrF/5ZeCzViQ/x80IMahhnO6oj+oq7
ZuO6zvOgT24AXaJGieSyTNoW+b3MZ4QiHS/xpzRONZa/e6y3lncEkBsE/d5mCAPS
XFj6GFr/0nNtO9uPhrbTOJqliDGi6q018KovO5gxGwHeKEra1KDYl9BmAnGXJnHO
8a4oLP+sNsdi6T7YReL+KV1Qbl/KTgELc4ajoj2A4ehThrFckOQj8W5i1LeCU9Rc
Re2E+VL6Tv6m4eVc+B/Fa3KwQGwCg/YDkXmlq88M2MLfef3wqkIGuqOFWypjGVZE
vuv4jj3jE7j3hiahbdkwjaccu+B8ypb0L6NzeleBSv6U3GOvBCTn72wSxqwW1TjY
SGtXZlrLbrF7EItSuhIv05SSQJ1pgl4zM2oRnjfov5HBc9mKIOPDp/xdaFXJqYeg
Oj4kcT1QewKkWdQjfskiFMpMeAxasH4J3gJPqMejQspHm9O8dgP/sZDTQV7axh1K
ripBhO9VD+UFtDlq6wD31JlrshLCre0YONsN1biHyZOXdSNkRVqdtFR+JS4voufF
qp8YmyGAv8CZptSdZVtsod+mPuIaeN5sULZn3UxKgmRn4Izg5FI4GpPdThNm1qKn
7agB0ptBBZI4sGTOkidVgxUVTES5RbYf78yhucrNPOAt6o0NNOhI16fHo4rcQMCy
Z2pIczITfkJpgWDcSByr5rwCo7eXOkCqZ8Q/TuBrFNeUA8dsXvT912ZiUXJdepIY
yvi1HrFJV/cck7xiX725+/vMV/ktOQgXsgJgiBjM21fDZqw0AlybWX8lliwmhdYi
ASFdpoW3U0/9qkF8e9w9p1x6YYPFfPxJLkmYkrRj+92bBQW/gDyh88fEAJGaZLqq
0+OGxuDXyzRGIXNM2DbkEMyfQXsZPsAIoJXeKexoExemWtcq3fXsZB4mwiZ3TIlk
Wgg64gdeZaYaJIZZzcrVx5WJ6OBG8CR+6osnSgfPv+wwcyq10wQnZrgbQW9/u3TV
XZc2vseFx3AKH0Mn7dEceZ/nP0Nx49zjpGAZhP6C5z05LxxPC1Y8Ea8mTZFS/QQF
yJX+sSmmJiz9RbJvkMxdT2Kebwn7A78zsItIZ6LrPHpiNkRvGZ22XLG4KKre5Op2
wf58uHE3MTcMAQnkN/Y/5WcHIX2dxea+uXWcJons/gWlq3kBS7ku4SS9K4NLJ1od
NshKIOtuvcGUAi9X9xCP22GFtIaEVIgGiAh1KLz5ku+B7/MM8aGBXBij14GojGQc
YYyeMSTuHHZxhPLV5RbP82IPGDq7unzpq8bzDWukupEwO5rXXBEsOOcuRFodTgoy
B28pogmcMr2CgnUDh7WqbZRQgU2xXGuwo6LYARNo1fT1+Dh+AnYsqwjloVwWEvSl
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bHZRsK3+7uWr79vL2w0Esg60sz+rE9jv+aAm4p4o7xcH44kG2X0K2/Hkoo+qSzBh
3yJIAnVUN2DICUswZuOLkVu74yu4qcArmAEkyFl+HAdedEkn08G6AfTB7Jc12ysF
s04iTPB2DFAhhb7VCFP4cPH4B3HtjaU8/BbyIwxYRnCIHmNaRbG4Vmca26Y1jBSh
heW4f98YBB0HInqi8doIAik/rTvzdIFd72J0vrXqz20+ZMPVd/3ZQZij5hboPI5z
njUDLbc62J3w0PXQBE7kEdtxjyegNISvR+c1HYzlyIq/+8ONsPttmpOWWs1X1gnw
8Na47BDxBkdnBU6vzm6Fzw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10448 )
`pragma protect data_block
pFMMYZASTz5B+roax34JCiyfM4tz1F8uuBeqm7yiOjxps6g3rF9DNtugtL6TJCUa
w5QaUv8YC36KtP5EU4Z2Y9yz3pIxyTPCQd7QAU/cRuStZ+hUX3jGqVgSaGGRfKy8
eaGlZ+j54VVoZTYiSZt/toTviQB4xV2IK4hoyyoD6nr+xckVBuxrVNMLoMcnIEQx
6l2PqYdPPqq4qdXjodHa/ezDJNhbXLEbL4Kd08PXiBA4PyhKzRNEpDGzGxepmQX4
c/VQOslTCprSCdYECFmjtCkFtVxfeRJK5SthC6VUwqcEDmDk3duoddK9wbRg7O4r
GyOcpT+DWjs7GTWx7WYG+c5wc9W2+mSGW4I1bknAq08sT9ds05/bhNtHuulyIXOR
f9/BkgjbaHxzb8aueyXLNtVTwxKyFGJa0A+CSqJAPUvZqtFqmQOKL9IM/Xup0naT
NWGeuBS/zw+ry61FWyLDoQkY/L0SpgoFc2QXu4Hi4L4eKU3hI4qdVSZD96L7JzfL
Zzl409jjy6rk9HjzLBVqvUAgptm7BMiPSDE6gvCskFIhQMtfw+M4vkQWMPGXVrAn
4Tef0bj23k2V3PRhmkimypj++nwds+sO+2BWlC2H28kA7ftq/m+b6qa3lT+Wj9PU
dIlT+sepoIG7dPTN9nMFu8RpGS0iE85D6xAkpXmj/3a4wZ2C1kdvXR+02kyBc6w0
LrPoZkwSgDi/3hvnu8ksw8nzjm6bI4AQeA6iTYlADn05yRsK9x1uyz8t/B19D2Nj
6+DAAN6XvkjUOBOq7pd08n0+AQVF4ngnhxfLdWh2KGvtepBUp9Laz2MWo3g1FXeL
OPGszZwpucfiIGkBQSzDsESy1n6MrlFo3vwgyfmj+H0QFlEGjGDULVulRvZvA5xY
3mCmVv8ccSYMmH2HBBuMOQ8BE8HWRdA2cIms1LGC9gnIV/47vtzI5w/8SYTMJsq2
5dcfBtJQ84wvO6xLrKx2SEsbSf2N10qfbyIX1IKbHRfHBkq5nJTxVaF8u6isOhoQ
GrD5fiOSDB4Rc9ShRr04/tENQDIBbufJSfb6UDcLsKfKpSxGLgbISjg1bQ6LfjbG
FL0StuNLjnSkzYLw1XGs73WPxcI+dcgtMUfjMMLu/RmjIrJ8eZrr2ZBCzvliGyyl
l34UOaDDW0596hy0vd6ILD7edkyglaRhfr+ljwMF+yh5m4sOANMZqp6F5mGa2w4x
rvbypeCNPgaLlXopmrpjaTaB9YqrazZqYarXCTDCaAhMtg2I01JnHVwK87E9molS
tkqoAShCjDhBdCbPeK5MjroZ/HBDMhfclHwS6lnh5eDZ/vUD3aMHSUYTOeKcLKDh
PlqX/pxz/+fC0vfWKMB7CQdHTAfVBdWvrbAAsdXvcWcyNBS2IspxabrbmIiVpnpB
osGLOWVE70MJuG66YqpqtLYoFS41trcuW+45oW4qfhCA3dqUPdQFKcXGjfugCpE7
HQ3JOKcfhmeiA0OY6Nu/AVeBxH3WBu+7DFVf8WCu7Cwqctq8PgVY884UIVMmSUgN
WLlQF1UhJ9h507Q9xDLkO1lF6wMgTW2NE0p4IXIBYjGxq9i5FF3Ej3pqo3BpaCgP
5zLDIRP7El2HTaZj3vFvnqcwgt21HWcr6BuUyXFxkp8xtgOcTqCGIi220qIy5tzI
Rxw/PKbkZ/ocAOpOxp3fAZZ1V/wIIKdHkUkhz6TnRwB0nWYivaxX6Ttmjl6MhPF+
qfzLsH2+wWHsmIse9HXlrgB+7M9pnKf/HTI647JeP2XpXicG0eh9JV0kGFLZvSXf
JtojsXGegQvpdSZQsA/sMwvGqRxr3UiGPbBC3u/xDdegMmwxe14+EFaV5NMOtObA
EoXs3bCeTh6K0xhd/ZBoBwtsV3d65SxpHgvwHjY24NhRSF6OwQQmHnD10Rn8J5R/
mSMVL2NvJEaNOwpukIhPqFsw5EIVFMeNr2Wo03uQJxy9ACW7FJN0Tm4jAHtsRryz
bXi+Yso6jfFO4anpxJYTbtJi4OatgP94GRPcmdtBni0w217G/gAoPCa1siRdS1WV
SjWWkVw/fS3uu2K0Vi2Xq3wbb5Kz9Ts91j3c4HBCFlCcl5cUNBSAQVAQxyZpN/ou
jw7ZrnsSk+HxHW+O0xvlAoJE8V0vULycy18qTd9CRs5YxCcCBIHxRZurzP9gQflP
TgQYHBFIRH838CM6oH3L7ZdhbXRPKB6APy8C5RMy7injX+dCe9ssxFequI6eBYgX
4XfE+KP7GTd5RKFCMN0TKiVm5zY8fEOj7gcTYVdl4adxX7KgWN0Fcs7tA0iBzLQ7
RsHTszutocSsbO9jlrp8FKBRRmlJJEFGW7PcqjZqDXVlAa+nDjsRQsj3NY3NSeYW
sYUL1ZVTqxuzOfxtme8OZHTSAPiMjzbRW3gesr80hbvn3jeaUTJFMNOPUlpaIsF2
F/GnKsAYp2tFDPr3qbDgT/VE24z7x8kmrWeYgU2Dc24xVag7VKgP67Lm/BOL75nw
CiiQrthtyBQKaVyzDWg381m3shTEGf1Wv4IubbkvyKvnWCepd1XuJZmb1nMFjUkT
gVYX0P5ryo8XfwYlbba0PnoDqbZ9GoI/A4pHobrzTVZuemwFrJVHmnqiEKmApcJM
eH4yMDDa16zLCs6jfe5htli6YXg53oAOic/34gCSTTKIFn6SK3ycXGL9Qf1hqGMw
oi8gOrErfezhZ4ngxilzbge9+zo/jrxB1yvBvGJjnXpPs4qjl6kxbdROpt4BVnHR
l2oHrO3q+D8uPeHsL3J/eq0g57799aLk+N0YYEIiS65QjmObsLiC+duV/VFpfcrp
zftTA8zDJdGTPZUavbTnwFL9sKJPkR3ElOhOMsjUQmxvKFOGHQiUBRhUsMEWtZxK
J7x3af5MEH4XhTlDdEozBxJ6XrgslzIu3W+kj2fgO0yYeOBMyE7nj01tCQflBF0p
04X3TJb1BpA5kmmXnZLsZ+bLJiHO0l4cE/VhPWojpHcZdF5ieGb++8GH/NRvM9vY
r1uWHfrMhKjY65J6R9u3uhNHhoebzuuBQNTKk9i77rc7xK3WG4Ydupn7d1w3wdXp
UUe0xxfoKR3JbpMpKijTIRclR1PMy8n3zydJESUtZMs7XLkeCOw6rHBPNmFpDuWL
w0znU2dzTDfffBXFdqtQaKVE1x2Bs2M8+Lh153Ey44cGt83+PZeR7IZi4CGH6Tf6
ppoILnumXGrbZNNsyRZeuMp6T5aa0sScAxJZS5LlsLBW6hWmW1AZzZR8cX2Gtz30
39bHPvj8y4cbfAbxguIv1qheqy2FqAZgI+/ojrlO8Iv7KBNQBSonNQkoohp6azl0
kuGWRpDVP45DIl1VYhQY/ZkPdCvqMD6HZjcw0ciQKnuDYVCS2QDgCPRHflO04s9J
ZROSeOr7S7TMnoET1J69Lq5Po4fLh3xWqEILhI4m+KS6jjtsZTrbiyaObLle9r4C
S6uL0Vb59LhFRjTMFHuR9zqmejj+ye4h7uPvDs5yDPpuYguqgCmGiT59sqM5Xkqe
jjnKZeb2FzlJO0UrOQyByltz0tcH8WZB6e40+XVH1g/1RyGMuRNGg24ystHgiagk
g6z7bAPrBVwTDUNECv0yJdgDJ0y8n2WefX1hADw80ndxxyFDOxhe8p6THqaEh8o8
gJWO8s8IGMsohuUx2cbRF6xHX2uerrdaD9fRMD92w6v6UiTKYJvc2BC/Y1t3oTPT
e6A/0aqzRp1TSsdGzZbB3jkxZVtpo/6N3UGumtmayCVoNnZ5t9FIM2E793Z6EdFs
JC1FuQRGAeyt11VOMRsa+69raTgXGturpnMV7/eo7WiQB+ikOQxqnHQF7U6Ot4Eb
opvMOG0eJNu000gGsdGeeuuKS2AWsb4grTPKv7M4hBZt7kCXDNgjeJVXz9fJ2pvt
rOFezZt53KlUwkgYV+TiCbtfrnP+3mzHpIEYDvtSJ1GuEugVaBRpbZSpLH+DH2bj
Ifwb0Daq8RbhoJxCXbxANnJz5qqGIdvFzCEGyvqUPl23K4WsC/9ukJy1463buSNW
1FZmx/pLi6ihUAZdsoTat5YaVDxnA6Y+hD5uB02Gb4oEuMwmORm0R/+waFfOEZdq
Y3XAICFybXJ/ayFqloCzzvuzQJzKQPldSwWtsLbg8iEY8ZnPr+bw/A70VrI5DBhc
s67o3UrWRAXosm6z7f4HanvbLTZSuvHTrQMeRO53JmdqDcKQHfCGKY6a4OBkdERC
MGklUrQOWF3KFzLnck8o0M+C0TnFQi5v32c/1sHNXilyGUM04n4wWbJG1XlUjW7w
ZaNTt/bRUK31A5SQcn5xRlfujyzx/SwkYiRAgUeOOXIGzvugr+DElcjyk5Ny1bDC
hgYZoHdyrZ1LaCDsKIzy8jBBsGarl8rvxzTtyUGWdysuVLqB1O4fvoTfYMZqhYuB
pAlk0hlj1QA0OFb8iKjmsA/LFjaC1QEwPR2b6YEOI3szoD83fpdoAsYr1yJRHhlM
8PZZ7K0jEwUL4OyMKwsURnVZjKo6l+BNZlpnf7LmFqbb3sh6U7smZQnh/lGPYFpy
dg8KKd4mEXBANdYtilVsBSt9+YEHY/RypAXyep/Jj8LkO+dRL0BHMW5aJ2M+6Q+t
8OPdWrnLO6kpqu/B5nGLOWHFQCUbsUM2T8sWJShuqA32uyL3SxXVdSVtImPI2Wdm
iD9WsCaRUjrjZA6Fya1XtXpgE5LVymqc8DPUpuSzDABo7hDx4WsPjdtTHGbJkmqU
BlSLD8f4A11U2NNxNUqpWndr5qJk905nRP6md1jNQOe7whTFB/fLk3BzSNTb+aLI
OsmWpx7KKBwJP35hFzRz1sYBtGm05t40jcNwiLfIiJC9WhpIhbL2oj3btW/jvgsF
IEe7DZKOPzVXnZtHI+tUbsg/fHlY1l4YjPPVmPGrnzjRpPmU27Q4ISaBXwK2krZS
WSJv7+9WqtcnNUFttcSyQuxsjJdy3MFEx4xO2Guuzns4RmqG0FeOGD1SqD8+QrIo
pSPIaMiQMvFwoYOVKfiwU1TcihFwykB45JjKkAybWYbuAC/7ZGY9HcnISD8PaTSz
0kSjg0m6/8IprLulpWeoI9JaP4jwo9RJM+kkaUXY5/vJ/t6v8tVVuJK/DNmCY2BA
Hwy+xNKh9mdJN5L0S82Vc8n6mV4G3avyIfIzbOyJKhToYvX8ucDmTCeEya36POcC
qgXOfRejt58Je3EsEQmslNUtyAUSmBtaU4W9BfcS8OXTD/bn0c8Hb5o5FdYXyL5K
qJD2mcyDlqnVI/I0mOKzDZ4NIvQXEALnZZENZ486f7b4W+Mz4L3xOZsNn6+mrvEZ
LCu6jTFO5goUAf35nZtBPYgK+71qWufc4UznDitSWD27LJW9e88wbnzf68sZ4Mrj
cZIGCvCwrc0Lrju+GWKiLp7V5zRXQRRZHQExD10diHmxhDW5/hBL08p+AxyTLis2
xap1gVrxFl1uHQLppyNXJHjIh83+Duro5TRPxUzG0QSxdrOcfbJUAp94YPqow3Df
n88Iyc8UfmJslu/SZWbHXWgd7YGZ6Oe1ZHD9VURtlMD32zLlQknLFnkV8zhSj/gm
CZcYtP9/pM/23n4/GBU+P77W2qBy8xm1jprvW/d80tpGqP27N1KgppHT09slZrzY
bgCWVBq1VN89Ekd+sCofckyKQIRI+8rJefWM+6TWANpzOOyt7Hge222xFXCc18Ec
2JQkTQ8OWd2knrv4h1ebafiOvJwAKrpRMA7UGbf8YLNakCmwvYzKol9Agx6SaEwc
iwfvuDoU66ZjINZa0bRKW0R42iOee6hS/XmA7yQUYHf1Mhwvsn2jzoA+UiHpEVds
qXyv+Fo8nSCjrn4Sv7i+6+M5gfdACSeCkEruMd+s+MYEHAKB60Rnu5ystH39UDjP
3XMT/SWmZkjEgMpTUnThZrMW3MJedFiNYvuF7x2M6f6xlpfx03/5fAvVjOZZJ5SJ
xTMaazFnV0XPLNrVr4DB821CO/9NM5rPrb/KLhN8bBfKGpVr/bXHr0ToWGkvAvWA
VpjS0P4pSKKB8GZfj9IWp9iEUA3eQ3DUvRQkaG3BjxH0R5taiFG5YcPcF1tiDbAo
dHkFsZ1HjLhexg/CRzOXfg6qk415rPp2cvm5R8p6xjLYjXtpUdDQ7VQupd4QOjyL
5oYZ6cXSatOMatCxRvM4jGyyE89qDMx2rCrxbXzq9XO5Xo+/Ozi/gfrdGaqXFTIo
xIUxI54//8AuVERwlAl5QMx9ybGaKoUmyVhICA9iJes/l3/Qy5ahdZIXDVgvP42p
y+ZWiYp2ReP3kvSPWOQX+37NZJkQMECwM1Ni6w63cTNDcvXYcu8N7kvMyE64fVkL
9tv+D09p5FqlIn8cZf1Qpa/wUdeqG/WI0zorUKQeqUJnQmTjnVdOFvTQzyD/sOUf
H0jWQcUpfZP49+J+eyE9pBVXKuwfWtggVDLtzTFt4ov0LYBa2HD57CZDurnAdSNo
+nEheoyHt/63hcPytfL8WiThYscjjlNfb68JjZmufkGot0VWHY6rjspxMFL5LGGW
QfGchv5oJccuRDJVh95we2isJRTzQJ1KtQ0aTidWwsj58k6pOrtDzMny4kZWDS5z
cVQEnyuANUyHkPFM1HW98vPHpo/I6ycmS6s5IL7s871WFFs7c2jRbNGqRZUeD9Fn
Z3V7+ke9YSTI02V2qSAF3eA3bsq4/clA47sx6l50wZ7tXKDmXDRsNnCsTJSuiVR4
GdB5W+fWtuh6br7iV3p+i+F0kY727vCOiKxlCvmffJUs99mBroOvvFserQjALZWD
Jl+yqJcXPeESJtXmx7+efecknkLKsn0KXyHNix6qixL2sVDLCW/uPmgVA4TlivfO
Tr+79zqKuxLPpuiAVDLvn5HpRo4soOx3RZRyRGr163UW0Wwcrj6xAwEUuLbsuYYR
NwTn4AFeVrqsYEd8x7lI45XqoeIeY0vyOaWowsaj+khYsPnvd/LBiowNsQPM7jXg
jrw5OLytn6WXVF5xDZx5NV97KRnoTUWAop3Bb5700fLPyrkZkgrMhNlYHvN4Q9fK
Hy96bxwtN+/cK5v4tldWxEPSYV5oIdTW73BujNfbRBvOhp0H/H/O8AVnU34sErhh
JpDDXDhnVu/Tgr657W1rQ1xAAabU03hjwmxvgUpBEafE7/QazySNBj1q6PpLDZaH
xiKQhqKaoQqSqhrqq5L/IH0H37LKmNdXL1Xwr4rxGieGUcRO99yMNv+Fhkkk+98D
tahPlO9gqJs4MmNClLvnEahqWOgNOAr/l2PIrdTQdO3LJ9y7p+/S9T5VMIhU/bl4
BtlYefdCocssLqqC2b5JcPtaQl0mfAzV9TkOYVliUFxiO75pdlHVGUBbyXS19ctE
5OkkI76guvw5jIC1Zsp+0pyyFAFQIqf1Ia0ZVlOerx+5koZHMdb21QipMSstV0hd
FSyIoSOtgrxOOabBedBfZ+jiARGYtKohvBHlmx3RVUYJNUsOY9PAd/h7OJGjHQv2
fHdjF6zG03C2bpI8obdLHZ689LElgMTx1kKFzwqaf4g7STcKRXZUh33RifaTfMGo
2/ecylpeFknGa93VXTsjg/H4blGmCOMC1dMIkMNmlDVvhO+4A+Hi4T/kKMWz6ACz
THz+dBs/X/Oe1wRiKX3FeYvoX6UjS6t1+88m/zKOR8oKSR5FYks4a5AVjlXo4JHG
OJ0UegaQbNCp8o2uqcu1I2P3an1rPP7kegKpzp3UaQqGc4T+M1kvvWpN6b8CMNDZ
dFN3TZ6izz2hjg/B2J8VwOKqL1poGkMLlxWttHTBUjSwaO1qnKD1IWUVnp1w+19C
70ovHIIVwMhCtxDyv9D5OgV49Ul2yL9tH0ojI5NRXztIDNTOARcfleZ+4Rakwku1
ZnUqQNtywCvPURxRrMM1B6Nag/Vk8XrUxw5XBgWWVwDUg1lzm2yiai80UkbogJy5
+1KRX7IsTBvAIK4YYQAdQIrz6psUdmSdWCVRk8JIpklhpxqLaU/JTO/WreFOvdvM
1fiKuBh7IFqWfu6KMWczeSLbtBdaa2+IECPMgqnEvFOt87NyJqLxD4lrnzaR+e7Y
Y/k4BBvllwdpJIui5pfhXtFjUWA/OAkgETryx7H1JHYDeMRRmIpcg3mo0+eGjVws
O5QQGQJbjsCqb5fTKpGQ5FWoq/w1+LWB1HhxkKuMQz5rqDYYedX7/7TgNjsAxoXV
tEBLYwSK2jEm3rA9eBLA7R0r3mwzJbSw/stlaK4KqlBCjDhZzJk5lkC1ND9dfAEd
d47YwYs+B0NlQit/Pmu6UG3mpiu0uhc+L2g/yWiUH3q5il/JLypylPudspxICkUF
hxFS9/3EkarQdBu9lHbgTTedG0k0WoGYxJwKt+it5ou23Tx05+oyfi7bFndSBX40
cvx+iUD5RkkW7nmBms+9MQ8MSJ3Y0TdmddBo3otTjy40ak2nsBg0DDwBU3PJue+g
axE2M7HLyq24bCFCVl6smT70LnQvW/vfLe4xPaSsvVM1kPk3Gg6HB9CzkwgnwT9Z
OU9AgZNQQ8AwPBdEICMVStku3cUeCwqVTSUaHxhwyTcFSotn/V+iil1frdoB16nh
j0zqeLcM1aAF2eBcW/H1W0zagIy2W8aIUZLrMkEbdsaRYuRYLfciM3YYlRwmqrOk
Tnhl9ypH6kUgXCDKYMeKdfFDn4FD/WPb4rACMU1sJL6B57+EYrFzYYKISjjrxx4h
tfGPRGKfymfDxkiSufBar2lL45owzK3kSY0e/zSAIklgjkr3o/oINDddiOLgQQYX
Hh+1igYXy613qZwTqegvE+F5uKIVAyNk2WZN3QxiPE8MrVLUGhYy2LpBCNaA5aVo
aIHcdB5mTFcBT0HQYw1FGSuUqXiIdc9s32WNKvHkNowA5g93a3xIBPgK1IY9M2/l
Y+ujd3yH99RORwvhtJyOR33hq3VsYcjGXRDzYNEykomzfPJYNy9ISVfOtgngqQRO
9nZGxlSk5skuFNpVdc+/tomw50wsGEV/0QNxaWc/8/jQhJwo7TihcTMQlWct+Aak
qzOnR1X0bGPRPFjbs29oHx+qT47yjnf7a3k33ITNdc6Sru+e8OXlvQG+bOZT91ef
0j8zBCO3NHKBFJhifgyKCCOkaqSy5mh0R8ffBNXKGZ8udzASIjl5/wH6ddwc3hsU
LmzmvVuIr8CPC5igmueYwFVFTLQWXh1AK99H84Ukq9w34t/h+Bf6QhuJBJ3DV2HS
/h3ag0EJi/zHFxuXpl/lc0SUoe32YXNQlYN+d5HJkbqGalIxYqBOV0b2rD4W38iF
oHPTQNAP6neZ1rsiapvnLS1NzKG3shH80aSsMeqxwKkkedxASIcYfnNE39cWOkwj
xVyNU4mFixePMbyg9xF9YSkVJoAtAmPZbFy+CJf3ImQlZtFMWYMHAc+2a9tDyNrN
ZeG9mf2l9eVvGiLhAFzPzMgfGRVgleYZSzsrTVZWtTNBME1JfLedA/hHlANoBVZz
feSURW0GhOHnyXO5Zb/S8bUAqEm1JXcyR1pKigaapr+JLRhOtd+ez6lBFx17ukgH
IIRLr8Ve8iOe3/Wx/6T3vVgUih+ADqmIhzmpI3q10Jg+FY9i595A9//Mib2v6Vxg
Fj2zTKPWOc6GoTf+eQgGbLYhdKR8tJMD7azNwe66LCNHwzOIUKLN7yyw1ZA9qD8G
yaElCkPGknp8XOA0SMiluWykodZsrNG7B5jyhH6HNMKcJDigQUCIYK+k9AiHlvQI
l8qsHLv+oQK1+MFSpD/0F59gTv4K6kpXq2HGpqrIqntpPJdindDAz/e+tTrgKzO0
ASvIqUQAdjFKMMGpKL8Zgy4jQr1FAbWRrb7iPySnT8lFrLNhKmC84kOi8BmbUf05
fXKeju48CzA8aFYSxSbzT8RuIjww0aObPXQ7EMtgAR8rJxNVy1MfBQlJ4Z2BZahq
MLhJk8yH8Fmd0OMT7RC6Ni3tQvtGZilyInknSunican82BxpYHb8YIg9dmlPL9D8
KziWxL2dZ5vXgtjaMdvjMq4AXGlXMqc5Fa6M3MRVnsFH05F9izz2GUMChM7OqPFg
Qqj6DClqCYjLFxBkJZ3mqRRPRHo2fURa7ajQbAL8YFlLLzXuLgzyTwL4MGtZzPFS
gWuvEMEjcY74FwaN8NR19SErCOzVZTFm4tCdyGIr0s0FA1X268bHToohIqqgitVs
5k1JFc/dcNpZbc1DMC/v1/WlifxoFmC3xM8m1F1H29NYMUrKJ8nUO/u4ezf3rscQ
q8zHv6xYMni/K4JVTl2E4YBrfj+rKr4bvlqrIaRs8qGr/S1M8TTLQun9TiLc97Cx
ltWTM3Lh0k4DAys9WaaJMTfMV0HAOWcqktf6o+jDTOI0dFY7nM6RcQRxfCuaL52S
0sLa4tGa97iUYbGA/MaVRwkX2zzY/mzZYdBvIpX5tc5pISLC8V0VPp3QQ9Q6Rm9G
eRp2Lv7IDWA3Q1/+CEmgoFtT7Jt5CeblL29JTBkBz1LIEDLLBm2VQOKPNHzBtw9F
yU33iKje0j4quN+e0Yq59a+lc0U9QzRM9quhMGi0MSc3vQFoF6wcGWEfKddd/a9E
6YJaYE20n9YsiwkEw+bLjlTuxDx98SYE6Pqf34C1HXGeaKSNsMKsGU0YM6NRO/Ld
ln5Nt5oc4UGqy/HOdI/sTb2cDo0VNYHIRkmpiQxhAsZvsfj6UGKEkaNsod3JbKXp
MdQbOVs+Gb87QmWDiiCY3Cs7bCkdezAqyFjrkiDQVtM5Cd+QaDZddcMA6zhSb8Hw
ohzhQltHHqGKVnmQpGjoULy/khn+PH7BBQAqAgJJ4ZtwrHT52Ij0TaOjaPykH1vD
DNSHzh/h+jJC2C50JR5ml84jcjfg5K1aNUMkFTk/bkTLrS0GaSbkilYzjPbXYKPi
/wiHMmdMYMTQcw5w9dU7eJiVoUQab3j6XIpl1AG0Yk79swjPBTUfWr6zV6fhbW/W
o8LLC8NEY5xm/2lwA8/sfCOFvNO3iEuCNGD+i8rugujkazEGAdXrXtal5LTmb8jT
8mTgAlyyKGjyUCWw7erfbnmZbUB4wLfB5AMEUTYH3Od66BqQdArzOwUvkEWWMq5F
HAoxzxqHLxNu7DW7Ux5IofUzNDbGNCi1kDp1U4kFZ10wb9zYNq9WdPAAykVtflvE
dy4wzSDpq8fxngumODJIEdMN+YeE9tzH71hU5c8bB4PUNUE9CO3PdRiN3ZAAFvWJ
Sv5kSJjd0e7DlvVC9/qCuC4fGitTqh0zwvD85J+wPH8fJ0DhANE960tkvv9wSN7h
SXE/BiS67kc47XnzsURWw3ySyK3YcrJ8cb/kqo76F07PMMGeuVzVt4SbCGcyL7k/
Ix8qZEHLQviAxYG/NP5DxgdsZqPXW112uKS+fL8yQLUDHhp1u4/2qPlY2P1S+eFO
B9NeGXMSiMOj26PKZH16W0Xr1krEQ9rOMSf/jS+2ovUZpcQRciZA5yU1RJeKKdod
sZh7Zgm2mnk0hFBe/mII166pB3f8OmeTCrFLNcp5/1fSkXXj6K/hP3UxeJysIJMU
S0WkqXMRg3s8LpiqPBn1cIR3TiWKff6pusi95rLzbGN6+aucUKbVziR0hiXhlkZq
TgLXdyXAOLlrUJgmWctFXOJwn7oXd+gMllt1bE4KQRUeBw9NaYunoxIo2txFo1NU
BliYDTZJYsGfexQJHKHcYmjAbpPWKbXzEM1DmKqMk4sfv5H/QoDK+6rErlM/1NN9
Ot1uRMd0R7deqQL2su5M8iM9c5f8uSQMcx9pkqTTRMYncMXOFflDZaf4Mf4Bwaef
T+rBxHNr9x//0fZTeTe0ZSJgpe1yHIVPeU4NMZXW+Fq7dd6JJXtFFEftaCMnDd5b
sdLkch65/XnZd3GZxR+cCLNhVUzt4mTtgLIVgAwDqKiRsJmRM6Phvd8DDeebO5ZZ
s0MH4DtBRuh4jhHOPvJEsmo0Z7EThrQG7phYfgOV7n8U2yW7kOKyf87ormmfOmrz
cpXUQM94ocUFjlcDBkrLOZ/e9rdWGcNd0/DbMg4M/orz49mNni9bYMfZguEX0hya
A8/SdwEtC7QAAIwDSUPkigOw7eLyXda96FNf4h8O71yBlwZd/XbC+sbsr20vQs4f
shh70RIKimXFttBdnIzzRT1/qcM+W6BqMIaYBHzByrEowmXg6xEy+siiHiDH/fyX
m+XSNixdCbmkgECUOpjkzUSW5WG3dU/qiahDydlxxi169KbVw6pm50xlpGNc4UrR
Hq08LGlWiDvnQ79/9kMMYawKBepVb4IXAO43U4taDbwE8lYnmxuLcOW9QR5REKkf
KUxyR4DYnXqc5msAXtrS16AuPG53bo1yxzyEky0XawnS31ZLgMzSV38sUTdMNDRU
LZQ62ztxjy1AohYB0/iCYvHE4VZTmtz4adp3Y5nP0Nw8RHc1uTHiG7BH5BiI7sB6
jAbNtqjNgsfAoHgv8/DfJX2kyHzYULteC6oWPvli1263OYf37zj/K/B9vh+Qrd8C
usjYZbeb8BIvahob11P1QX0LtE5FL8svo0ZRIlvnrAOubqryjrUXr4K/sYpcREdk
qCPzkBy9Q2vMoXmOczA5XvjMZ+zWYFE0JzITlE9tKbggaEK/ft2F7cPLxUD4R2dm
vtFsW/k5k0httBZOONt1PnHsOk6XT2fPGgByLuq6Ds7avyCas/+PVgSJhl2sRSvW
WcC4W9dSBXxgFAKFtJACqSVttjdhiHpxJRr7mgz7Z95IEdplH9o4U88nsVjOkIDO
bBjj+l4fV25FTm60d2hYRELI2EdZn8UbfVOvvam7muXcWECbAzqeLQK/o9xPPGwZ
nUWGlr+EwqlFDausuWeq57k4G8uYghK7/mOteojXae+uh7dRzEtzlvjwWSUD4FMr
mCBHLiDzeGgjggo2O/hGVIYt+wzGvvNyZPBGZWct2hSjG9WIk7jYoUp1VC0D4TsO
tuJ43IsGx5fn4AaBmzgenS/sGXeBWbB9NhuPmDb2M3wjVgN3Xelbn0GTxS2DvpSI
q+xwcvckabgJxHQDCN0zDJe5TJxZP7iNHtny+grl3C84kwIcBQ3/lyztRs3aQOx7
DsIRZHnA7JcR5hDUPar1XV817J5KSstWge510Pc2KkLg/+QO64/CPqq60v0ss4pZ
GM7VE+jOZ3XTFHRSvEmaXhoZf1wx9Awx67MWTK8WQBvDx57DVdF02c2IjMMOZZJp
TFN6/U5N/6skZr8g3OViuBN44Cm+I2kzfwy+6CT/MDJvUfDNzlP0GBPLtBK0ojUg
pkvEMtpJrM8/5PCJRTI6oTX7BGlidfdLmMcaLNax7pd3vSsn4rurzquD4G6+jugx
XC9OO66M5LM4FsbXB4Klk77QXGIeRDk2pMIEOJKbtS/jcWCxdDLMAyj9FvE3xYJ0
YUfGg1kfrQF6X32SV53st/wd13fKc84SUBkBkhXdz+IjTHQsew51jgrWImfSKfWU
eYUmO12wHnswZZ1ihHkALTnLwgeE2nlKqjOzeieUbmqSVauIqw9eOg6ZrZmueDzc
4ce9KDfNNDzE7yLMFarQxxLsbLPaD+LNfaKN2a5zNQdjKPM6dCL00oSwPK+1Ejbv
NSYOLtY4CE8AN0wDPdiZGZyelcH81hH3B8h4PDdfQQjAVCu5Sea8HEzLiScuyD+o
RUkxfEqATUo4S3Q+od/PdqanORnAf0yCZn4vzEUewfTzxqURRPw7lxd03Vm4yY09
JTHg6FCslwsOQV2yVFWCybhOoXgHTv3DdVL3HtRoaKp7bwITUZKfz7BNhanaCing
TcpEfthUrv7EG8KYXB/rzYbw3FqL/NG393IV+HP+LqvktaTT50+AbmFHMpIB4iBQ
YISUlR7irEKrLvQ3Fchsxi2HrfRzhQ5i5uwXB0bQ8cjOFVzKv9XmVmHxve0qUupE
kTpRAUq+5h7vac0u99tzkmwIF1zSXIQ7swKVCkNIxn4=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TjxqAsJ1GICwon2GKgg8j1d5Gn0K2BhaioS5583DyK2EYObce7H3JzUNAU8w5zcq
QrZPcvBpU5MLmK+PfN67wfbEuxWx1qtIT/kZ3Kis8E0fusVDM9w7BzjDrobTCqUH
rdFPtLZFpf77BsA77vLdAlVbL/1nmGLjmbyS+KjvbQ8xEbpYWg8foAI8XvaPYCla
RtSyrPBOQy2muAmXqL0jDkffdokgRGYPPUFMD+agTJvoQoP1mpGA+d8hJz1a2Ogq
bw9tt9aJIh2X9t9pkz0NjtGUgQl1ztYY0AvxzRWjRft3zrEnej72os/EbUUiHQQj
GRTnpm1ZAjQRXxZp5yL6/g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
ZR9nKtcVi+uwwngrqvh/yybM65IYknZt2NhoG+UYnrhj+9zAHPMcTlop8HIndP2I
rlDVBtDl1+Ca5h8SVP+TT5So0npjBjbXi1AkteJhOwf5s9fQ6DIsLQKNDoxVxN9E
64m+Vefl1DLsM3aA+qrZXN13T5+URsCEdQqBJjpI6eJ9sFLOuivqS3ksi1lWSItd
Bczea9HpZ9iuxsdYaxWWu7fCtfjxkyluTHiARwHx4zEEveX3S3oB+XT9QoWVmxHt
EPVzuI3s8UlD1PpvzI3WT2e8PbUjJesw3bEHzYIQaajTK4uEgp09FWR9wuVIShAI
n2BLLn+99pvY3PBbF3ZiyPIPdiCJhuhZqhj8uRbEAINuwiZ/R3aZfIsBTft6g+Bc
E1PEdUiT0eRMtmdxqvWeezZbg1e6w4PYmvq5W0qYV1/EEmmucRTAZCT+PC7mRIuN
AUwepbPzaUzPo6PqMLylYb0mP/saSlHNlmZwOfZfbeyZYM1Kg8QNt61JI+AZYrCj
xF1gl8m7TtXELW7XeNIg0Ks+o+XX77LFG2DtHFXg56lfSdDG9fDP+RAs6gdD+QEw
9QwTZGAkqKArCbuesitBi992jcQXXA5ZuBy2zJVwECr8se8nELsJ8L4yYUbBCp21
5l9eCnocNLfCwKIJcQvpZwjK+ZBGeNoOVRSdWiNXhfwaDEkb746quU0FIOomrbOJ
AdZyyghIqzu6m7qRob7s4KWUXFoxvDyD1gQni4eUqW5jSKMYXgCnifoxvunmtb2G
UclJLOZhIXoeUyqzxrVuU5HUtNcd1X+rtgvWiWvfpuF0cweHon8HXw/WoSChMiKI
TqfH1Dbb+rAWr8lQ332ZKTZGgZtC/k/m3anydLtc2eibezSiYp/JWM91q01AAbKL
tqMpWattU9VgTR+6mawrGNpsHNjyV9oCY8QFHtkQeZMlVR+5RbuprjNYNPSSywO4
LY81sd0H/drAmxstJ/cFyouSFL0m+Se7F0eYkiGUP15FFI71ZlDMrXT0RGa5mU+E
9vthp0NYk7+axOIvJucPbnFu9uj0PdVttWicnQ7piC79LemBhNV4scQha2Zjv/Fl
8edIGMU8T+4wfB+f05yvQtATFX9XbuDPOrIlBAo4Vk58dipMPNcNpK5afsDbGcbL
7lpg1334vEngA0sIWCH0Sg9g2Tea19B1AOlmq0zuVMgzQ5KsP109RpjsNmpXZxYw
9N49JdlN7hiYKBHnJyjjBaUTQQDgHIyTWQyUyFP7PYrHFqSXTQoAFNOhsT9R8ujP
qX+f1YNosxm8w+eifufSrvvd5jYMjYkL4YZ9TL75cDkb+QZzk4VWbcE4J+yKXI0M
LAX0KY7rIcRc7qPzDkfELML20gVB8j3lpgRuElc3EubPnVTedTgoE7v88q/fufRc
jWomgDz4Vbyf3n0smUcs4caUwpzCYsK7EOqwVUOCd2Vl9SpJXDId2n5+IIoAtCfp
b4TFxY5X4WN9EIrq2IIwutXPzoxSwY3a44uylJxiCDp1BrWZhGm/WqFLN0987khL
a8mmvmTE267LpdZ2dF/Yq+jAxsVdpxTbbjd3CCXsiteR/WJx+3sg38dakjM2Qpg4
BuIhrvpvfEKlBnqbEFODI/v0tPXby7QkD5vsDSHllnu9SuFn2Lh5d7/a4kxjYIhX
jQBAwD1tUJoyGQBpLTLq2D4e/DnEEQYIg2hdYE/fzl3LQvPtm4B41U3SjtrlimOP
etnWbfbRRVImMJaEA/MF4xZLJNlVfcJ6NbdmqOorySx/+Gm+tMgfVq3lSToE+GDJ
+X8e8JTGBWnnQe3qqOBe9eZRcy8o7yglG0eoWUZ83keZwjQBe+oi6aF0joQEcJjd
Jnsjty4uGpjPKeerttBIOWWAfUpblc/TWA3e9KzSRo1B7TWmgn6hF7o4YhIqkCZc
AZasvEv0iK71Z2ZzDCU33t0g9lKpHyt3MLQYPEIajk+aO46eAgDnkQbSmzYCMGUI
BTldM406Smd4jb3nplm50p2QXqWU1xoCUam4jNxi9gV0uYjXMSTg2Y1rb6OpSoZp
rim6kmzoDu8/WUqf2KOJYpdsKe/IKUhRR2ru2Ca/N4oiuz+NydnM1coiiV3E+tDL
eh6Rsq1MtUW01KtVZ3n9pf6Wvlcp1ReIzkbn5yeHBr8nEecRCYWCel39Q5CAaGp/
ZXwYiVIbu9rIdbdBnaJatGVDROKo3hECN0Nj14G33KGdwdWL0vTlkGiqROrGec2t
mOzuUsavD55DjPVklBJbe8Ny35jN8R1fSvNeA4I/AE+5yxtEuyATHqBbCFYdSHDe
+LlECcCpUkWp8TaMtqO9ia3bEr33UGl1d5P0b19SBKWm4SHfcsP2UdLvWh6HjrcJ
YtW224NyPF1ruqFOu3dyKZePhVTIsxcHC/zS3EZ4+hyILB51okYclzpL+DD+ABeL
WcPOAWXW+gRvTXq9LN3Qo0MvoUADTjtc6K2LijV3RZAqHaTN7KfCf0SCtKCIH+gN
UjgF+sHqB2y6LSLMjb3kQodUavviZAqCJnivXALkKsj941imD1cvAkHkxE19Cohg
SeqvgPT9s/nhp6QPSw3rX0e/laJ86gfErk1jJzndB0al8qJZ6+66zrzzqy6f38qY
urB9fvfZKiFLQUS9bxrBjGrq165ba+JrHBipdHsQMUuG6q9ZGYIoPDQdTmEiDaXQ
p6OsWS7kz8xmrLYcWR6Zz7HqiJO//A79B9A54GHjiy/8Ny602EYBoRcn4JN+So9g
mUDyHQXKaPozPvVr/wWL+zL6sCH/PzrGQeCpWVa7XpCVlUGsNxlhF8W0CEDBmq7o
JIqVU3duZqju6TgZls2nNAQofLg/8SulgsxpFyfDBNDLo50Q+QZc3SEJCNpItaZE
xgmFnKQ3/wgvndRDhOEvrNzbVGurp1u9ub1e7J7vRDthxnTm9ElfJtq0qxzAG+hR
Db2xMP+UCo8ye1HVQaqDvz6xw8wXO81yFbNHUVqkNw/8jSdSs+AxYUIxAGNupb6C
amB2ryfYp0FFL/ddffdTaKNASPgk8ghS4GnufISjgvexP5wt1spuL5dU9TtP7qfb
YmkUJJCvpqNLQN5xTxonYhBibcyM+AwI5vgXaFP1GFXU4YzMDQoYprNPhr7ucuwc
QjKwH7dcaIQY5JbsZr3YpfcM3U2wkYEG/kwd7yyAMUHTvw4vlQN7blerB57Wvd+2
VKyun0CLSsAX/TN6TpOObQwH8umZbIqB+GjwIUrk8CDYccyXqL9klPdjHZHD9EsI
yCMriqPIzXGhy/d1BDLLyMDBs6KeJRHF/7QsMpA7JsTJoIMD+Hbf3c0m5N3Clp2u
frt+kc/pSNzSs6QXBgENEny+RIC8hksYrXxb0+cPWJmnRwzeddgH9fN/2d78MxWW
AYkI0EuwXagnJA2dyT0Sq91/aEH6mCXcgAPS2KQvfu9uA6UEUKoBqSwv+iYdDpsH
IWO/rWL/HGp7KBFCXU4lh6kouNzCvurO2zqA2/nP3E3NCi81v3lj8QOyotJnsjX6
FoL2D/EUKORYl+LxKJTMHB2pgbPt4ctbw4neWxonCq0ld62xBdbEGevQBW6LBkA0
xbUcPqjAz2ktVkp2zj7+3/NxTBhNy18Tgjldh/OkZQUTRyxAq4JozW+l89NukCCe
2q/Y3vifux9kwsg4rlTNOmi7T1HsqqisVX/EnECWG9qzZ7mAf9CoFr5RRJdk34g4
dTk6AGQWyOuBVR4eqzu1E2wrTuUrQgkYW/iAcqQCHrKxaIILwW7Ch2zJKWgEW4P6
N3+xhUXFWqAV3zVoxAlcODyOx68zNmYWFhgqEP7Fq0PzVQ7FVq3jUvG+H9Icbq7f
AZMRSmtUhwVz8xTFBHRlLLXLzLgpwIA7K+USjsNnGChgA+A/MsB71XHu9AJojwM3
WEISHnBiy3hzD1GfHt9NpHwA/8iV3r94hhVNc1MGjQiSLKNhdJpPUuOSYz5JxcDG
uvDs1BsnIMUbIr3j29vaHpui/ZMGoC6p7Y///QwCWunGib1JA3nNFzAi9rQjBinF
OAtqUmsEEoCYHJ13BsXhm5yUfqeXexg0DQWZeiKUTkx5qVYU1MHoYZqezi5a44Mk
SpGsH+GeNHxfJUfxAstOGHPx5Gsw2uRbYowXmp7V0u7TfOeOtRN3V1kPVtcClFX/
iRWu9AQ2ariXAdoPrzXcPA9G+B2BKiAqy0VMjmnu7ReexNX36adyIaYL9S19CCFZ
1JnBJpon/oBAJeBrIAgZitaejpNj4d6qCBaG+/8nCaw6yWc+xSrKtNctDWhKyq6v
eVKdk43eDmRc83w8+KSgtSEaenhc2P+53s//0gMJs9WhHEGBCd65K+/hWCrzgZ9r
l++F6L53zNo1A16w4YU5HNQrchiGBW2myIKyWCbGSemBgUQmAW3BVbTjtCnjPOeg
qRx/nRcUv8dUEHfPv1meD3w0FwMw/bulUaZ4diZtOuYPBGG0oHc1Xz+2BLnDShfm
8/gofoen17w+BDH7C1w1IRst424U1Ph9CDG9rbGaw+8/9UYmkX1JuQjME+ocz156
8VUmYtmQVJrpRqqTtxzZDNVg/astmEYJW21dCCR7ymTvW9USG17nL9p9TV3a6Ark
z9mPzek22FmQnM67ezzouX2YHC67508FLdZWl2swv8yLHAFmeWFYBWe6dkvHUir2
yZiezt9/jfiLTehLzjEbaMV1GhvgXpmr5G7R7fKetMKCNbRP8MQS4b9T6ZHfcvZc
tXK1lFfdItMc3Rnt23PdIxs0KFFBqk+v9jqd/aDDQKrE38zzcDE+n5TzXH2Z3qdu
1ZJWDKy65RfjDRfyi666XYuBXi7NqWobOuyBNSLv7vnfcK2j4gl38iHPB/SVnm1O
5IdUZ8sgHiRSUZRW/Id4O/1FURTRyeyj3LDh3KKwKMtuvGOuIXaBlKMejxf2L/6A
42iTLHOI87oefDsmzPZn4c9sHsmifl7oYJm/VEPt+yi6RKrUo4YxPG5TpdrVz8L+
5FePKaS4D0Y6Mh9vtBo1Q2+oq2Ocyf6xsDsZjR9jQj8WD11Im6P9ouaji6ldiECW
hu9iiGM9ZS0KY8CnWu88A63P8BxrWj4Y9vG1aFkEvHDz4vpyPZmlGYukqk9vFH3A
LZD0zDtO3Wt60ZmaVyp8tKQBFuHJcvkKemlj3/IvNYLlJaClluLPOzoq1USGofEQ
quCOx+nEtWdtpH9ZPB9nQgQmld9+u/GoJ23IGpzzuhy+t5vryJcpg4enEwVoTrVP
Shz1Z6HY1AOHsE04KVdlFRqO4kutc5n6ge8mlveOtcl+kUb70dSlXnvTezhvBAKy
/L6TbRQBl7oBypBarGoRoKbSG7Iz2WywstvUnjb2jfdoYKleIs9Ftz3Hr/yvPLr2
FVI6fdp6a/qiTFBkwqktUwSmCa2qrLEcW37oNpcLklOFdvykeQ3V+gcgiOVDISb1
ORiXX0cBqMg8utGWHidtuDFgO3d5moS5SNIbe3U6MItjD/yC03r2KDnetUJDBEDf
W4OTclLHADS3PhkTAC9s8LNzD0R2VGGTtNOs3d4InTZgCrC7gKGQF2yqQ6Jpyh1b
/SQVbgbK4TqvlXzLe4mGO14OPYBwpP6hoptCtIaYXA6ybAR23DdfGStSjl02l5VM
/u6rkDkUC5hVsP9gmtqZXucZDedh4qwt4jsLGybJVFq1GQFe+dDOVyRoRPa1lrGU
kbb8qlNXBBRSdDVIh1WfwJetDWE+HQYn4MN5JzZkIbaCIzkr7KwLqNfx7Qfp1WG+
G64syhUpacSn4W/67fYarwkPKDCItXY4agYKVv9p0Np35TbXik00zb42q6OuAXZD
dhx67AOHXFx1ZLpR7PJnxkccHSk9Y/3UfGWoVbAKeZqBkZwA8iRA6riGMoHz0ggC
I8SADru9/KGCq0ekuzicCUi3uhjR8hvdZr7Gqk3Se1ZUOkcWB7BBdiIUL3VjntQP
RM//DWeD1IIlcqGaYnMlhXbG43HWIRwaPMnuT5eb78yRNu3XHTbATZTKDJpUeQbq
8m1WmA0PdCIDrSRKXC9bS/0/57lePXeqXsNZ54GzV1C0oV+4eNUQT3UnI5H54dXG
VCBYyyZFRRT+u8RAftsYucVTayaN/FSTSM4rd/MDM+soVlcdJogjqam/H1CvEqzM
/+LLXK4Rk2I6x/E4GJfU+WBDEX1gbpkrJdVTaT/PWdfOsadC4jcAYc5BUbgMpbSe
iOxUGmFiprC+5Zx26/Ka22pomYb/Du50KQ0FFvLfN9D7EHcpG6d3pUUxOtbmXofe
NzhzNOk5lkhNsXmdUwvlWvE1TNlF1Kg8XUNJhAzF4NUzDxowiKtcKQFOokmownTE
+/nlvgLAFa1LQYdGMbTgCr3uvwkov1wHHsgp2kB//uf9VOajua7xomfaogJPner/
I6qQRlxRjGvxZ1TcugmoTQD5OVN0sYLgqI8+wq3j0YxkMrQL/opqvfExBlsrtodJ
sDsjoxsglxt6IAYctjgbLy8hksZYO3JOEa7cZ00ghcN5jVe0Onei2YKBU7GjzZy3
kpSDsYP7RN5aJLzGwAZXY+h0ZPG/VeZPTb+/9vLpDg40kRbc3dK1c4s1qcO+InRk
MSc6c+NJu/Ut+zKJvq8uoChuXXL4YIg4pfySXVUGyU4pBjJT88HIEf7AZaQyY9Gw
n8Awu68d7frrS/z1KZ9ThANoUMcZeFRK7JQghT+YQOwmKFN5TtlSLM1EH+/B1YFY
Z+o1An8duTdBpW0r3EWGJtTT6i1U0YjrH23EH56TIlJR2twAi63WzWkoJsdNVLst
8w0UuVjihfd9QjIivd7pHQuWOJEvk8T+m6M2k1ifjaCUTHY4+nwL2XiYfhagup4w
6kcRsCmMZWZpgctSr1nm1fYPUmMAeXI1oalbTDQ8EUkwTZPJZwXkOZveDnGccRwL
RVYa9hs9HTMGYr99vAcbdG1BU1eLsXykhC4YxB0RcHjt5KdyYIvKMUDkgAy0M33j
LjJs2oLdAyPMkkotC7/Fbc4Eq9ppMoL86JUmWAFGfrh6qKdKyPkkTAiw+7fg9qDh
CZZTYfWJTUNh7a2Dm20uNM2I4H6exdE09y8ZjYe8nKMyZs4npEDclMKph0CCbxNY
G1lEY63HVXYLSdLbltgVRjlgwf/Y6iGcmefmDB7tjTnskPvk8dGMp1op6VnCjKfH
CDzSgX540R+xdpETdT1M/blGVSZs+KsU3vgmodFHjiqzcPqNSsucMoxzeIAn3Znl
4UfqVRr3x60kie3+caL/QRBRFWJ93YyMY1LLn0fzBbhEUnu+ZITHLiwl+9w9hiyX
mR8bQCETH85NAmbJ/4SdrRpq5Bz2rHDRylgQL0KiXqFeXi/n28uHz6Nh1ACyxDmz
AUq8UhMbqT+f48hQjbNQyeLQVWXGf18+TpPSL0Wdjazh6oco67v4kd351xx/L41c
FSLHDQGvG7qHU3Jn9mk4qki5taMvVxrOOmYjUmz6w/BaTAAUgsD15d13dhic44XH
BGvrj5H9sl1ZHXXW8ZPHJXr8MAtCJZvDB4ol2rDXbZgEok5msxXCPozesSQ28W9D
PuDHUWQNSMe3Jf/RUo3voYo9/XfsZLDat+WNVh7NgxrPgA8oRf8yIaLxd2Mf0752
xhQO5XYLaZON0h7115ZTWYBcVV0HlT/W6Qb3DSNk1z1LnWSfoz2GAs9VtnmJl8zd
tSw32HKOXFA9cLUsWHUekhi/t62bbQP8JR6gcc9/VoS8lpLICyiO5zZd0XGzESjr
4ETOfYO8qL65qRomGGTJHEV8exMtmRqR3g6ZrqVpq/idiFcQtOQJF9wVpMEaZTv8
2WGvRjQtUQFoZN+jwY+m1mAnvH+UdSoxJlX2nNk//AnOZlVTaZrGkQ6Z+TSHlIFd
MZGup0onQdkvvWd8xotm5ltO/R402fbXj3gxwJpApQcETNmcGy8QMrYmVeA+Z2z6
+An3T4CFSby5wPKdgNVD/Brhvnz7oxz+FiI8CRywPSe0fEPACtKRV3Fgl+ucE0pU
0upfi7ZJ5LslDLRkIA958g==
`pragma protect end_protected

//pragma protect end
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Atf0Jg/8xJszFVkoaJtcOuiXjvpcD2hSZzx+IopxcjPjra63t8RyFP+iTmszuATX
W3niCw/40ish9jr5BJbzYCWsVIkvjwd/beeeIOnVK3b2c4T2OPInOabMcNt1j2a2
qPC2bgSw4/4++yeuRUmKdDmEgYZqFXimFcHQUpBOIj043eMw8CvtJ4+exH0aVnDD
CqhUrNxS30kL8H+rpAwMVPdBCsnTBP6aNXfTZsN6D34TtU8erBO2aNuDXSfI5MWP
ZFV11ZLoZOVXHbK38+sv03KtSufj4S6hfbr5CN8zLc3ZZWdXgxa3kTvlw6mN9Mec
vNHB7dJpTIMvlJULRemKIQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14480 )
`pragma protect data_block
62HPZtrU1ME02SV9xFbt1S90Qiyo9d2ogpuz/b+gE/Z59ehrWlTK22KWn74JN4gJ
32xwPUhtY54MDVDAT9HECNM8eB8rWa7ljQg/YxyUy8Qtcp6sGBRUE7feq8fbQNcU
CteitVqzl85RQVfHpHPyUQFUCRIIOzlj4hUKhgIUh9vD+tncjZLjizEJ5hb1a6aU
2YyrTUVoD/r5nXzAdKLZuAlP9NHSgNR6w2Q/VkBfjC0Px7FwVVcU4uGys1R8floB
Ggmz5WlAlaqmKGl8bors8286iN9b/M08VAMVBJBjO6WX0AqKnh40oCg8P1zDjuQE
bKCB6MccNWcooOBNERhwyUbHzcx/8HcdO4VmyVL+isiIF0CbPnIY+ZtreqebXeZT
pZgx+DfXDFWzZeS4YrTincYz+M1pZntnOhkj17BCQan9XIRtsTGRjQXysl0T1oTC
tzYH57PlwdcLkAFUPZo+HgRtDM1B3nPUlbIK37GJand34jvN5fC3/wmTAn49SBo2
SajAhkFwS2+gL/Aq+VZop5SUafkvqUAKd1Sft8+5SaaeTj7OnfvyWjc6aov3P/vT
5YTovfL1ZJH3FmSzurGZRvw1p9UvK01vFd8uoxwvBU8XsYPkvwILI3iZDFqn/jTW
iAPiqgF+mHICo0YRJIrY7GHsMLKsyKcCNQG8Wr+nRc7TPsEJb8K64rYFmcVNkXN7
DKUqvfXGFRTDqrl02bNoo2Q85B8yPxrUazGLKX6wKCCuiMAZkpNh26lqAYA5M4A9
eYHSmo8Nx6Obtf68J6t3kYfT4YXiIdxqHtOt5EW3obcslPL5iEWTi1ua5TBKiOTS
iF1+PIbo0+kht3lzHUf0DeRHA98EZ7yKuoV2XvSb8InQ00QAMOFqIXhlyLl+Xtq5
C14gfT8vMLnDPCkGaAb4OzEy1RfdC4Lyh1NOp3E5yhxgEH9XoM0tgO1COaWt4+G8
II2bA7qJ8EdgNz/tj3h/nrvvvV/tr+Xxp+Ixr2DSaIBgRTpGOBMyWe02H2pw2y/w
+02vAlVTitzYM4e2vZ/GRzWberF6bHP6+UeM1snRGOhyQiZB2EBszcld/asOmcZ4
r7HU2ZgUW2YfNVy+V7I2VPsJcAXLDj5Bnc12saVVaYv6UAwGJYiGxFxuz4B4c4Zj
55zP81X2s9QEd6zuUcT35WMsQm1QLURh7MHegynQOWb9rwWakTzO9mLBXqPkQpG9
uTCvbbkA2VZRqHYR0OhzUYOPUtAYFAJdHWmZ4b6MrF8aYicRLIeiafyCVdOFI08o
wYaPlH/4SiLtfpZqwI5BqgW/xE8T6PF1nASdAs9EaLQYo5fzA42qlLmWIPCJPHzr
8Lh7sjNzfEv9QeQTbGd47UZrCixS8VGIdU9j0eO9QowU2PfRqE7atidKSsqn/hCD
F0X0uM7qg90/24pahl79/w6pzTUkSQEN1qEHxONwVrCsbDnty6T5JKH7QPrWQmKk
rBr63SUmZQlQYyH8hkoOjBGFIVYY+VmYiHv62EY9hKGAe9Je/wDl8gOyFDjgraVh
2ER+Sxk/6k6zhnT/gFoQS8o4KhfnPF+wmMEDAxSXS7Jt75S5bIW2sC55g2Tg87mC
trrs4VpFu1yRUa+L5qJg4HN0UCHN4IBaY3wOsoeej24LqbeTmDVogSvR6mm4eB8l
GjI0n6YbWkBWKJ8RPn6MWxStzEy6KRkTh6i9djdzBWz3Ml6U6oT2TxsPb1ojBEFT
H347YWtagKPeiKrM4FxFde9xzk1riPHZ6C/4XbNiRS5E8HlcI5e8HitBjobo4hJs
0p6Q1NKdP1lFZKSXnrAEmhnNkxsm5FVAGRAo0WG6vZMfzqTDiVcYUJbPzVJWn2yE
ljH8g0RvFaZxGNatDqkxTwUb8wHeYo61eBFcmFJkqwzbtvetOFYEYvrGYUeINM0z
G8YmySVzJvHJGdcusMi2ZicdzurM47KhfsSBkM0SFNuns+ftAlmTwa1uFZPzx4Nz
0xja0B6OUefELD3ap05SQLqwUaSAeGnHo9xEZBsxlK0QCBfXUCacPSWGJn956hnT
l64MBrGFBWwGoXeEx+g+1WHm9LvlMAlhdrxVOf081/2FXqH3KX5aSG6vJk1ewSMD
Az0e+hJS2KJsmSftYb5S8eLRdq0y85R7Cni+KXqisnmqSEhUFLn1x5M9EDmbrgzC
RJGWwmwvIn/vx2ZxNVn5eL9HvmL9sFAiwqSXIkWmLY5misp8I2DAij9IEETHDUC4
MbwsyR2Nzv93HWOWHT3iYucvLx910a+NRtzYRRBdXQd4PHOskCFRRP1P7NETHDdN
j976fxLDuir6OdOiTPoCXOmQoc9XuLNcrFzwFucgR3ockBa7z9K4Bfkfnv18heQS
vt0fcNV0Qx3zAC5N70k24tGjTueEWhIooL50OtAFZikde/5cQt5iDeLqnHHkbJ84
6pdGMUfc/7hKB0gdQpr8af/kxSzv61dYueZPNYlLWdXJydc/pIhQ3mFbgj6ZvWTj
KlSokS3DXzNlfomTO/ifBGVWevcx1YTicHKHRHnlHCQDMGhtvrU8G4JP5a02htG7
+ua39NjCPDLmKkSvwlSfrmR6xrTjTEap2DmHKXc9JqYa32aRdK7YHkGvAYwxjkFe
SRu0yI2rFwIp7LkgV+4fz0rk+3j9vF9x0ZsLJCJdLYEussT/0iuAg1uTmTbrXaoH
NXLzIIY3w72f8lN5BuoiyFZizjFW52VaNzlVCaC37xhw1UY3IjC0AD8Ei3dFopPc
MOOf3z/Ga8/iJx3wAJb2IWCEFpDrIZIIdWhZVzkJlt/TzyQ9FTXnSIu1eQ4Fa1PV
MAfMLfIlz4vbk05urlQKEQESl/gBIzlF43Y26DgXcW6P45PW2FZwW5DDh7SfDW9s
aWqG5OGdvWLQydpWogV/bi3eVOfhbdcvpIYfOSx2jN4PzyAgJUhjycmNtWbghpli
KxUZFfdHvTG9dHb3VMpOSU3NbBw2i6Q8TCFC0RZggL0mZaQc3356oHRNyV4Dkpvv
SStgqu2rX2QrfnVZH4AWG36yN7L9P6/zd/pDm63tOpE+Q368KTjJjHxhXv7Jx0NM
DOH0zP6QNCHvL3GmxPpMEDFeDRJx2iO0QwvZt+FPdy6V3asFCi78JkyUIk4657qe
wlEuIekF8Nl2gETF2h51Nf5C7NT5AnyMWESjZV+6u7ykQ4bBzje41Gh5Fo3ZFau/
QXLD19dnLHVNr9v1tYFxGuXij7Dqi9uNr0USrd312iUl55rKs4KSKHXw3+MN8oHF
mmq/a6kLmPpkEX+9uS2aKwwhuQva3VuVlQ1UNxtw0j519yNndTM+QEfslW3scSlt
l4U4JeDRiHK6x4i88wAFFFt0X1fC2bnfRQFkjuA+vxnTKMnUyIrp7T+RlgFfMtJE
C9PnX8Xr5vj2lErQfOYU6pcH5n4twrexQ5h33msU7vitSuuyRq2Wn/1+smA3w3x/
gr1q2uF/CiKg2iE239AKYTFN2Lws9cgPDBlewO2IGIGMEtLs9WjAeIrXabGwRtX3
J6XkSmxDGP8cwWTEupnXEwcZXjEPCKdKjPP7JZddwGE2EKRxn2vjhNDHAqnTyLaC
spbVirsDU4QVFMsE1R/CwNOOrW+Uxu5OTBNYQO3h8F+Rh4+3efFYIPzR3mbi1ZBL
zRWRDdLc8kVzD1Z5meBhmOAxI63UZpaggkxotV1s1qd37BJ92vsayEYjqxaml5qm
TY128YnFvW3W0x2FcAFHnpGvWMWTSGU9d0n/qCwa5322dF1RgguzQ/AAEul2r1LL
KGVx2V0okmfDFetPrh32xJ0EjQOBkmARGspXPS9OxgsMX8SJg7LEDC16nCpYLM2F
+M5rRY6xkJCl+R1NdgzW0vvKPmtYVHx3WjChXorEeszaOr7wB4iMfqEHJskPuqic
p5TRE1AxXkZ3Gv/OnTl8wAdMSE7wFX+TFWv+8B9ZhB9H+p+bBlangmcZ61WkQOZP
h/Bra8VER5xE/tYhIKP3/1fcgn4qEKdaALyt0udoXeibuaAsET94ML5+6rZBLCnX
5lTRWwC726BKNbOFLTvY91ra6yYwHdNmbNYflX9h23xjkYYB0BaWkwRzWVIWAgcI
Z1u8bCe5msCdyPERdX1RpMcVU+gDmPL++W3ucfPzUc4jwpW/KH2TVRCCYVvVTBdc
mJh2n2EoSJxVVhX5hf9grSFKDPj9QnkD0ol9APg2q7CYyvri4QDS76Vz+xCMbgD6
7N0x5UW7BTkh0d7ZbowrsRKAY5HWaaRMRSabKi0/k87o8k+KvaMGxI7djrynsZ6Z
pU+YtPqPZTVJKYnyxEUxrPISvmy98hDK51D8omw/vHNqssWKIog1Xa1pTgVL/6ya
AYByui0OKLztFaqJ3kl0OlT4orUSkmQYd6nc2d4mDsySkuPWiuHTj7i6ML5kGgnL
uIx7UXNnis91k00tY34imfJOb2IYB3/IAsxZU98FSVfxtVSKHcLRwJPLo4Ky40kP
02n8vP7R9LLSCAE3Tla/w2oXnVwMqPE+IdZ7pMqpb0PbAbTNRNTZSwniY/w+nMSA
Cvwqjf1Hz2VL8VutjQD6TIwlhenWrrDFxN68PkUO32BdO2QMgXj9UOex/6k0SQNw
NWYsosImvSL3Wx4Y4WcQzsUf2g90dXQPF14R/TBLjyvhJyS2z/KLKFD89TnHiZDw
qNwJdsy/jsNt4oZBYeySaUZBm/akY6AVo/Jv18q6v2KCwhNF86XxxPX7w5YiDOB5
vJmiSdeoomXdwh/xuG5ZtuisQ1YwY1yYBSl5x+3moRKRT6L2Tv+ri76ZBBjh76MI
AEtjIQhWp15SJtuQief+rhStWsP0wiS7k8y8YPRpw7cAw8NTsQaNmLsbLEGoEuID
vNbVOyum3WvpOYS+4RrFD5Y62S5+zB94RZVaj4DDWtQFwJ0zsSTXAVZfGB1zwL1K
ujBNplTVnmqTfD0c/mNN4jeRdf94zpqav/nKsTTPQ4heZQccunNIlungsFDwoyeh
XMjv4nJKcHTDicJso1QHCGWQ6ULR/ZmnLMcl6PMy2aV2jsaXcL4piMZdZISosq0H
hpd+MV4RuB8rb0QQL1MtKQpvs75/1Ps5ypy2jc5/+1/582hdX7T9GqIUsRdnBOOP
14ONMM7mZVmnFFoVw9tZGhlbFWd9FI8EDFP92tCPaogIPz/bYhZKTU6BZSuqCeqM
rq+GcdzoDBv6apFlu5B/KzERe/siQyME9NkgrBAQu5J2Ua1wxYEsPzwkQwbZELim
1J+VNatEHz9rCSeZVQe/SV6dW2Sa4f3CooDTt5AurAzBb6HwR3AVwsi8JUA0M/V+
TrbV4QJxDOW2Yma5CWbXupl9Fmxyc0nL3N4oi71piQB57Yq5E7OVk06q14KPwT0c
KP87wfwMKg4oesg5R0c+WsWzDPu0Rdvu3llOSUblQ4HXE7sQu0S9pvRbu582JDUL
dE5iDnktipS5P1aLVlTGZbHN9ONNnA8mzkLnvJdFmD27koOacu2hiMi5VBraJaJN
II5lIHGLOBwblfKe9zCf856jMY53zTdutmpRlozs/YvzE+w2DDXOe+yZuohWp4h0
GK6pvhJzvtfCfBV2GkVV1/b9/d3mGxTqjfppCCtBk8A4k/y6LyhPSOcO34wmyUYl
BKYxIyDj48zwVilJlKRQ6KnpfD9yjZhWkuZeqdr94nIIA63APMIJVjLb0SQG3cJY
iEg3nPDZvNz23MpG0nrAUvdVHJrNqCG8YPY2CobH/tFN8rYH/GnXkgatNNaGwvXW
feH42J/0UVid+q+yLWNALyi1bsWY/IIpyLjn0sgMYOQ4cSvH5IMBNVE6xbAtp4cM
0R+DnPJu8NJMUVEXywDyp6P5JKql1NcDcIPN586n0fL1nXv4vYCCxVKRr1eI/KMm
buupCb5FRfeB7/14n4QGbWAYcAOo66MaKyYxKpJYEJPyr0JXOSYwz3wBv5Z8IKWg
mfvtDO/73fyAC2YruJi7K40oymv95rUYLnXtSPayGlce7HBu4+4Xy/o8wnmGVP/k
3uA9lIy9hJJOEFW2ul0Lplb2RR2P2XMjIs+FOS6Rp4DQVzbLrrSrW6LT64/ozm8q
9BFvZyS5Et/WFSgQN5+96FAH7ArDn2O85GS+adu2jXiP4iI2Bswn5sXtUoDpjZAd
6B9SmZ9XzadjyIh6zP0uSHgMBGUk0+Fvxufz206IhVrrOKOUWRMFl+VrUJbOc4GD
TM0Bbjf4ldFgAWwdT0DHiyYS7OYjdhP3SCiCiA+SwF38vQevHOJ1uLBp0B9dVAk6
VaulTDk4QfnOAVnGlvNZS1cqOMbu7R3JOC0xEiK3InLg72+v4ZeYLKtqdg2hldk4
eCiyLofrgvRdn+Kxv2XFXHc3wdDAU1g76NVP/IdcCgO+3hb3+ZQpCIeB4GJ/m7GQ
nNb5cBMjwOGTiC/ny/XxHhgGfJ9Mz84ShnAGBN8vgoZjyuaRmItGe1QL5rQNz6bN
fXCEC5BAJKfg67sqd65gPhiFvwWxw0D3x84QK9KiAbj4f6I/ZdbHqWRw2YSy387d
4+4ndgPbQSO+7q6hLHagj+C4+tvYdmNVryQ/zwrb07aSvB1iLGMqjNP5gG7pvgTx
691b0Zj02xHhhp8sqppThgVplSZ+Mz+/hYUBCqOSrmp/77oFiJJb/gLVMn8zckhg
hOg2jM1PpeEsusZ4TBK7e9zM3N7VPy31pWLCJ3TxGJ0/wYgk7iawARUbMzUgARLr
aD7NZJ5Ff5N0xsV1WnwVswnSsLM30CZEL+qglATwly1tDMDsIkB3EBe9kBQ64D6H
iwI81P4vneUrnUSRtuQr0ienEvJcfKmlIrQPlvs9pJGMJVNAe+f48kWcfrciBe97
7L4cZTsdWif2IR9UhfhKy95o9n9d2fHn+2b3B0prCCZHYH6REe7iWnXZ2FmPW9aG
6UhH9vHqBYXraakwDRQU0A2vd+UrCooWF6RbpQ78oyTnamUkfB8qJHbifkaPRmqu
0DGgEVVGxAB+1NP9wsC00pS1OcLB/x5LViGcJVVIH8ryoOJ0cs/USsPcSWDDGj4A
lKZVnHMILBX9RTupnOU+KFt2crvK9KY9AsFNGcYJqiY7R0bey74uK42QmW3YeFGE
EMO4X11IT1kzMu0QE4JHw9+l5PkJgSjWHw2WcFgGXnkF+1U6OVPHqKrJjR6HTJnG
Q/VGYi/goeSHhWFhr4Apt9gN/0Tvag0awunyDb5YNj0HHF2KiEA/a9GfUbv5gz+N
RHc3QD3adErOEUeztYI0ni4SdFZFe4AsvjweDb1y0ooGDqR/NvmbcrGTWSC/IDm7
sygJTGmJ8p7XrkhDRZye9Op1akzqhFc/N3pDLCHW5BRgYQJM0XwoQVKZpaz8H1wX
MxWJNojxmEl8r0XTsypS86LG3DLX/n+rya93uv4fBDiWFeNGxZLoyGfPPES+Oikh
LAoUKthhbYEa9tM7b+S9jaqXrJRfN1nBenvZCF0SRJDE//B83/tDEQZI8HIkgQNS
vYej2JhBrAmp2tZJrgbN1/8hPt+0zzni1wChQaVafto2Jrn9wHu9iZZi1k18vmX6
h0N0JWE6oFGZ/sQt2Bw1TQFm6bNeuJC2gQDlIrOTo51fLyXkkmMz5Gzs4qK2j2XS
QioMvV2n5v0RBylAW1p9J2KVaHoMhg9BoQhcYbijr2BKJzVvdy4Qrg+g8/wCYTn7
2AVr9XYaQQ0TSNZfZb8YX5X2dtfDZwaMy1RiBPlQ1qP7jWlhvlK/ZJ42Ojy//nvl
AM6QkSGhkRs+DySYuMYqc6RANURU+GOu+6pZ89RgcdxOq+pQkq+tGdvt75sQs8A9
tjK2JDIIQ7ihZ3NUBlnDN50SjXPbGfcXR58HHbLZ+EyyAeLMowisfaHurKbTSXQf
ttkdf1SRTPQ/gkz1aS3eEo9vL2mSpmvhT1FdcC2WeXN8qlXJ1G7dLTobm1pCxcXL
glK/UbjOM82XBNRINwvOZU381cPsY/7hcLVI0YFWKJjv8PT0KOB3ZLLuGLiucWOi
e1/teciAREmIG/gW7KIepoVwM+CHig3aDjk3KCf7xOgGb7SQTA9en64d8z1QTPDo
t5qFFveZ/dmMm0+wsBGg9Bvt5Dl2d+AaaESF3/R8K7WXC9d4NXYbcnW3MrZNmD8Q
uaCtzyHyDtCsS6wo5mMi7dU4s+YxjeUC4Pye+Mh/HqRQ0dos3d/yA8X+Bp5JTb4g
t02Wbflp4LaIpZQnsFJXK4Zsx+/JVPlN3J5HxOA6N9nTCs0SSfZFdtlJF5rnN4HO
LbwIB/1OWyICijFRhXHlR5ZW6vEnM7/kitANEmKsvmi81Ngl+ueX285gvz+zTzSm
PnNu2EzUaJvwwyWKtXskx+1Pcx6JQMfHJ2FOCNekaXfMOLcK/ZJHbSfhDoT/N0h3
5RFX1Y4JfF+9lbgHPKhwxJ+as1eudgqtLfYPzPEP9DFPSPFWmU2bbS9lf8b2atcJ
LdZYTUOY54ESNOC6fRLLbEmYyrU6WtGnpL275o2f5kpohKCQd1p3r+DJ4Z/fRZkO
vDxS7+RYzazsIY9Cx7SW0MGBITUGyV1rKQOm50fQGCuqPjZRP+C2+GyIxjsdCaA6
jXESoTMz4dYepYOeqDWoj6v1adFhNNDaWVkPNY0bnztza6Zqyx70O79ESWFaTyYy
XV/+rM/IH0m/p7NYJ/1d1FBOKMvY+qQgdPcLxBabjNNtTXH0n1XR8FJ5JeWhHC1p
S8Lz0eW+T3ahT7B0iJUNBnXLmT666QsQ62UvJDiTej6X+wH+DCC5reCPVFg4gfad
iQFzCk9W4e/iAVtzvoYn5oI74rKGxOjSIzJ8vEDDzpIy6uIh/aDLFqIxu+7ko6fq
jr4yM8nmD8bV/DCDRG8zzhEqXKZ5ehs2ABdPJQyN04Tao5m5JuaSnCbFpTG1qBND
Xyj9Ob+S0vZrvvwP+9Kra53NJmWJ7E4jR4f+CA1d3OWValVfYitJT89JoZtOwSki
+RxTCOzK7wJIOqZmR8t+65THR+3jPOwqhSR6oQrMyyMfWtDp+6k2kw+9H+5u7aJP
x2M4edWK040xQWL+SF9HOSOcYWMYnwEfjlZgvRMcn2LTXCgi2DhG0Hx4ycJaC2jw
G2qiCXtE8wvTV7u7LavBHBiDhDFdUlo+Zq7U0Anr2qxgUGeZOakVx1uiVagpL0Pw
i2vqUmEzYnZ7RrOcBuW15TbOg17+RQL15HaoHCuYHdrPkQTin6mBn51R5T6148cW
4ffAgcQVxPfdr0ylBNzHw6PMC9Pd5719s4qaZrXSwx2BVtSAvfVgP0lTq5FRm2JZ
o+JupO322IM9kDpCWDjEJY3blLAMxekF6oaaXnl1U1YpQ9R9j6mhee1cn7oUyBL+
p3O/++iXPFW+aBggepUBvuyPhOLNsIhubQIQuw0WevLZQtraMANbGlOOUv97U/1L
XozaCCOVZMncCwg57wnvihdUUmu9UkKsXMzVfgYZQvNXzv8ODqhz8rxps2JuEW9v
8PCTW+TOgmN3TTt9zYuVvbm2b7emuOm08eY+nvazJAHtber7Z6UBZjl5dM65mOtM
qYZZWf1gPyO9lIopADamvCkdOHTIrUbRXGgusBx57wsro9QZK90Yvl/OwwDqHmw6
RvJ3UXzjVKRcXd2xy7cf2ANrvez5Uls5SGSvsl/yh6110rARQrXn7ifqL/8QuzMY
Tn4vKYV5pMJ+yFvSOa1OkPojw4B8vHoJnQ4DwNwmaSKJJ6oZmbZ9ZGGM8rMOaN8D
idZLkZNpcTpJ9U6u9FY/nBNlq2EcjV2IRd0Q5UiOPEOmLoFRsiTyFk63pBCSD2LD
cLITcQ2E19/PEpAlGDrhz1rZx1I1BnM+7pEdSCa+ITIkNnEgcLdnrygTnhWhTNnc
HOFYT7/wSv4FTnptr6qmSJvTMEt0+AcQUNaieVGHIYOLTGIhWZ7/JDKBmGtSLJKy
lsJci2v8s7dZ4NUjzUSj4FpZrO8WM+7hXWCTXZEcdnD77eawidZt/H8np5sd6lCm
E1hLI6nvuIbkhseeKqSyWkgCdVR00BwaLt9a+EN/Cbi+J4833zRpAbANs1/O727E
aOMQpjxS8TiSmIqukQdH5fy6vvLJGqXHsN3AKKn5dPrHD+JAUCIX5Qdls57ErAMN
QqCNOpfDWAx5Mmnpixl91yLoMT/Ot7M/o2iTK3yOew+Zjl34F4VDuk7bngRUxb7R
G5RCByDT3y+ubL4k5em0u+9MOL/grLdHT3DX7fbHCNgXQ4GLtxiioYN8I7cVlJmO
WiYeKh8pY7yvDdV+PZTRi0h4e6LmrlmTcH1ZOobuqOgy+R28NTXW9x5MSn+wASAn
tDanCr2wwTBqnXYhE4vGzW26IIRmlL7ffGfvf9QwYFxrFSZvl1fyQNM4FboK2LTX
85VMj6ifZZ7HM5nn4RLzAqhDebjDLIlFAXJrj3iND8SLP44nN1jj50zm7TK9uPR6
9YrdNyGKzBROtXY7QlNWetFN77i8DEARgT8jcZzvVbJZiplIEY32D1o7zZL55jeI
5ROPqfAnclVOEcu98k8zXq+QzwjPqsDbWXlVa0cJ5i2v81cYj82B+0SasX8zXlxu
UYZVwNdLe1bQaVm+ETl/9l4CfFsTZWJj6R6sUvQmtssJSMAzUSY5+b97o2iOaw8m
NWk/d3Byt8FdI0oR9Q/b9KxlG+JYO2BlaZHud3sIjwnHdnRpGuxQ4603h08UW0rA
lGetuAL5MAezWUSJ4ekTPbB71luCvJIThCNR6kaCkrFZAFK1xvvIF3a6tP6CMh3q
pmP/yg8GqmEYL7mBJ9NY3Kl9U/NHnBois8f+jAIn1HXKnnnI7ZdMbBa7STGorMEu
DwHuk0sGGpiq/NJZu70qK5cT4A75HgSfWUfZDJdRS3WD1XQBIYEFS2lANXJpC+Mh
6PaIpbjunMI5PH94GyUmdbA2HfPCmYv39jbQ9ZCIeYxsLcyHpHl+9F1s8qfClT3F
kmaPlWu0+jOFqVkk3UTgT1s0MCPAmxrjTBr9ztctMkDV5vYoREfFvBv152VXtXCo
48fIhv3b9bi17YMcyFTCzpSXvfL2a7cfO4+GJdPTYJ2cIBwLOMFjNrdX2S0isdJ/
v8NyWcbOW1LhdeEPdyZdmkeI65u2BgDIfydxV/Y1nJvwj8rCOYfx2of6m/e1b2/s
JuqOku9xCdUKxlZOxSCA4AAdKr0cKJrL8eZg5gXjLWvxCAS6uN69VJGZNRO06Qsi
dqDnN45MTpGD/A06BThn2Q6dI9Vnk5rKSWGnr/LVen+u8eclbNvOgHuloc977zD3
z4Lc/cWj/5sjJuptmMzP5vnLRCsfyC7TD4wfvcDX7zeb5l85z7qfjmnhX4buCu6o
S78qdkAvTRqoUl9qMlBjTNX7Tb1w/VWi5+XYyX0A7h09XQSYEhkAJ9E5mKfamgS7
6rAKCKM36JvCg8vhuhcapB6+loyhFl4G6DN+DGsHfnen3g4pBybHAJ1B8TKjHWuG
gDJhrtDVerlqXb2e3BQB41IOkTTMF7ZoolgBjRhr1q4dhcydzsjmJXxaSbC3028p
zWQmybnb9EyIwN1oYQzZeyMgNiqxrsD2hV4f2BYL5wmsGw4tQ7EKzdN0Uf4E2yWj
OD3gr8F6WXcx+HimCLy8Hmz2W6kAgQ39xkwsO84dHlSMpzcKxuB9p3zLtgv23G/0
YFtjUK5wbTGlDK+a3h3oVcrp7J+bc/WqH3d+o1SU8g4TL4YBj5jTQFiT8uD9Qi5Y
XGnFpgNJ+VrsPTh56Ee92fdDTuFVP9rR8QCyY9iOUzDavs7y8KSMwSugxEvyYZGf
gATmsUm+RRqdtFy1Xf9y+VSnd/V/I3eY/WYBXKT5/X7Ir15weRtcVJFpmDdcNEop
LpqiRxRdvE3gLb0T9S9PKRAhvxjWnsLLswVZ6zl+Xf+G7Jdc7u+023aDKSq06kg6
+UBCpk5eZnSWznDtPPeEO7GHYx/m8htahRbh5jcQdG5QVxolJuBq8qWuxO0c+AsV
LypA13WkzDfVrAPKHgXRHCVXVnh64LjCpFVc7JUumdP3Ifp4Vd7yLDXlXc4UBgp1
fB0EReXFbLAtsllC1NW0aBOvnGHQNKwNx+J4OUJA1LwVWIhOQUIkJvNHHYxpw4fL
PjiFG+mNEdoIajCd0xBHyEEOe2QvwCM7pRd5mPSl0lGSFFWoEZnjKplf5Eaf1irl
ah6GNOnZPN2OOVj0mTSIOXO7FZNRRU89iXWZrL//NhqV3Anw4OnCAusjyDtbQQi1
c/itYvVuT91BkxNQgycZ11x7PgGngDa2ME1wQdGfx3ya9Pi2V7m72tei1XvBUxxY
HzJhdPTwBK6jqeEQTvfw5Tme96XnnrON5aQHeE7ZHpZMISujHucZw+xR9pPddYDe
2sZDOt48IRuVxLt/5Hkro5iBkLEv1pDBNErlw7Fr9eUGuTNGe5HUehIGaNtWPLoN
IGQWgPnIWLpbBfmek6gt8QDLssZDAPZmF6XdWGZo7gEwqklzkTzsKEfYF7cXAmne
NQozYrtqGOFyErPgfODLNOJkFPF9XjMSmswVOkYA/qPEHyLopqjpb6Qx6fr3Ag7m
kYy/rG9Dj0DgPf38/zfjgBdMOEwqFyykVOEsDzQ1G4hY3O/N/yXy0EtcEc0E92Rm
3/qdj+PW7DYDOYYIDrGR+wemsMAniUjS0SuecNcy+GCXbEbiYhhzZOz85CCVE8uE
Iz5IiB91KGXRcejGPKCPfdRZGE5kJLtuRPrWLJI+tWMB/zfQGj6D7xw1jUs/FykA
PBCWoanjk4DSecFcIpkQInAf4TCn0ZrPGFd6HtLyuCtHhvSJcxogvtjGl5wZ5W40
o0e8igImICTo+K9N1anWr6Cu6z8Ab8tCE0lPrsqSRe4hz6lmqt197htiHyuzxA4n
UEqqbnE4Wxg3Gs3xmB+0XPsjf2vG+SnzNF8IXEseM/uYJI2wlTaOk1EZlcBp6zEn
hRzRbLx7xg/gmTnPh7uI2D+2HkjfO9wyD6QcjcxF9gxPSgm81QbMkiZWNl/aCnJN
EwBd8dLxnjVYWqYFjLhfaf6nfGFwC//SPpKzjjOfrH18T1CJoTkUnQi4oNQVsJPl
AiGVM+7BdMFwdwof/qidghOcAsxozPKvhxm29IrQ+VTrLEc4Z/p1UBJoqoXXWfya
gZ92hdEqsQY1hKatyVqhYcsJeKIAEVkEAoG5NJ4Uh6Ye9W3QfbXPAPPHXKm+AH7o
tDbmp7wB9KCbMyrrbmJxo5qqKv9APfeF12czQFL0RCzLkt7MI4jqndEuvhifgZE2
vjiXSJd/bOJ+lDJtgoqlHKbYgWNjTipajLILMwhH4kKXeoNN7uosGUILLDpNqR0q
olCBrUfuA3nSP1XrDK8DAND4wSzMhflDbj6FVyKiwFJ3NrQ5dn1r6KSU56MU6jqv
cB/wX59ksbvbf6RJsUTXhEA5+GuxjrA2ZOoSqIFGWHXNiIlrDdAZ8uwTHznOFPDP
zDinFJ3io6kwYhcB13+IfEXR/tfD9fn+spmkZ7lRwdk7zpeMIsO+dUCHc/3xkhZp
eXyT4GIF9YNFfD/r5olTeAUi1dMAgkPTJELcu/MTso1xEp9jqCgkdyqARjZnXJK+
Wk1cVfG14uzLgDawgEZEu5B7k/kt0ldtR/HI9FMNTmAiVurRS4dnDSDcD0sXaVSb
NrozvOS/qFKe9VsRcsxoniMUv2yoLFpjec2h5zlYpoW204NhWp+hrRt79Q08ma6E
63D5GMYg3YK7/8WALebZJEmo9hK5rE26GvYmCjhw5YlxJUK7ZAzAd73CpVfriy2D
SDRxxqgSbC7kUZDxcXg6imj34JuOuezUhEKIAd0kVBvzanhitwPXgfA/CIHBGSTY
bhbrURZXHsJoUmc3vKombhO5CAsj45qsL5tc8ldt+UolSZrF0ziVcXGIv3GXkHaO
o00umG7SgOwRtfteeT+tkO2YHJ7uAPB44u7OhBPXg9JuoREHwjm2ySngj6xUwuQq
4SMueO9rpxjvfvjJw0v0l5V8zw7Ke61Pt9+NRLqYVKNwm2ocY/nj5Ml1wB0BuVHa
9mURAboygAvonG43hiX/44kCg9OavvP0zJyA6Oh9l9wy2pA9zT477gYTCIdZ31nD
2q7FjojDJ+QkUP2vKnUEi66jpVrcko+zwoJ+HrDWefmJev4OCJmMNKfy8JZFvRXZ
tg2rc0EK0H8dnvqAfI40AFp2sK1xAjlOtMK6GqC/ZWbyscsMbSdL4/l+63/S9K7h
Tw4obvx58V3icdIR7YMjbMrc7W0sVNJCDr92io2Mb6ZQVftHQzIldT+OqDmX2viA
lQPfj6MbbkFLDwbi228rG+XOkJzRVFxrgYg4UrcuaKoVeLVJoERQb09SlfQ7geyn
H7hhc4X9j+wG2A+B/iXzdmzdhc11pVm36nlixdSzYET2pjjmjIGCtgFkmr9eWgkX
84ibA4p95QvXSrQJy1syxTAZdIyc3VFXOOJVTUOHX8OQZW9tSsUsqA5QcPCqSSQa
kdlnN3KykPf76f09L0rR4Xjh/I45oDefvFA7jF9F96DZlr3QS5XFrAqJtMUDNUJn
VJtNS3J6rZn4hXw6sKkP7aHrkVeaDYeExxj/OO9ewGRokxTG7vdomEKjF2pB7ocS
XF3vZvCsJLpIeT8wgdjiSpm7WUW0iJwNNUGbPhiyuVUwYjCQ6/3+e4MprjKfQf2z
BJx7B4evyMnbmmxx5U3LWZkB88ZPp9pdfwrB0eaDab0oKwRBePekje/wUs5Gyjpn
/zZOV29nM8Z5xcUQhP2zEBGrM2DxmlyZSz2zs5KpOY0vgiGKRzIt6dqHFvIu8SnR
ve3WT1wRFKR5RTxeoeYnu7Nl4i1OPe50fnTAKPzRqMFV8oy+oYTJEEo/hIOetQrm
LA90MUdPlYfCXvldJB9ofY74MeMDkJR6cnU1Cc7jIQY0xnzb6wq00M0WtfhOvt/P
7quO+1iUdKqzvccbCR7KdsqK5dDqH7NdnM/Yg6YUYwZsVlY0JFgMPIu8fIVi6Scc
0yDVJy7iEbiUhOXbHrGjJ12oeT5IN4DelmUqTnZWmvLpXyoETN6r95rojwOtyRxx
ue5a35rvpKtwwuUkANx35SnUWdOIVsgXKjjcoxEzPGfA8MD5Z1/LoJhrIMhzMhLP
so2LhuRvcjbJCxmF7+5pNDd+lOcuwo4CEZM8qwuT3HoH0jUo1qC9y85h+nbBDzha
KYnW3MFWH6+Wtefc8a+ArF2nQS9uLUoYZfCImRAOXsZpAAe+pM52ZvazD6KKnS1D
tMiJajc1V5z9yqztyjzVCEfh9Sp7rHpicjA7LDzeOkMryMd9Xjt9oJ7VIPc/me5P
wqZCLR4lmctvbHpf0DvUTkxfA01N5iXf/zoJZADCZGRbBXE7/MIdQnJVOanmBzuI
HGRS+DaDNcc6dXZWRd6IcC6bheJrNp9Tinq4JS1RghkBWTOoTJ/uA9GQJvxCVvjP
xVhsrcARsieEVdLnkAf/T9DYjVvhcIzwsHHwCE7IzOsZ/ekk6W/Gxh+1G5kyCads
+j1y56Jf8jWj99lVAcmsj4hfzdbqYjWRnLuqZUFuC2sUabSh+mJrCynBmKqy2FIL
zUb+qAQV/E8tfAyw0Ess9PCURDvc4DMJh71WcTu5RrchDefEDh1lHjf4JIa50OY0
7+Gf4QVtuNtbpG749bIlt8PeolUHHA2ONWFp//5qTSmub/52LDVD35vjjnn3UHyh
fbGIZFVpUzL+VGZbwZi7hdJM8lyCipPxjqPrOlWZiTQwoorGQUmqDJsGcGO50Vox
7I3aueikdA4oaxVu5YgFx0edP50cvXGAvHawfRTB6T249si1uXQXBkWc3NWybYSk
/yGl/MV3g7FDQvqq4lqZiCXszNF4dzwvY/O17D0vdtHoW+je4I5W4Y7+D3mpWd6q
KTf4Nyo5xeBRtmX/oCFTzXvt8spNqhOmdfqWX2bxIFM+DRE2Duzikvpmydrm90WV
3OJ5FTR4iFM2XnmPhck3LUHRy+dPOQ+i0MAYd92CBPF/CYAMX2/FXnppsWWO3Wg4
jXJ6bittz7nYFaAZ3zbx/J8xDGgjCXHp7pSAbYBiIZPwCFy3ed7U9EvDL5QRgVBg
oPU6Fr7euNfrs5rCBd7iWLoP//8UWyKALbUh9RCtPmsRKYTGhKKi6z4hYVpVQUzj
TvQdYExcTYqsY24LwKAxcbGDFd3GJLlRhZwH9U0lZOV6zvUoRGX2JWG3RFSyPolR
cQkXS6lHvMTyG/P0lCXSHnwjIK6W5yemgtetWf3WAHhdpgPnOjFJMs0AIUi9nIUE
eqlIEQp01Rl7FmaPhVKB/cXAnLUM0Zwv5hDXVVTo2A1+fy5Z1dQIXqcm041YQ6lb
CSdavMP6RW/fjHbxewTeEXR6eGK+Ce7sNF1yyAWxxcpyWLls5altFrBSzphm6F8F
dXZiGSKAilnwEsf6jU9yJe2vwWZkUjsdU5B9cuMGTnJ2E1WAOMSAinqvyvdajE9S
TMypCshMe5i6HlD3V1HBqBapXNx8zV3Bc3ZigC2f3Bsny6PoTgYzEMhdaNZyeWoe
YktVCnc0KwBPuc/3YhmknaOsWeB6WoOqh1+smTQvxT1kBScW9QwkN3Axq8EW0xPy
1k/t7j/VrwcIz2MlEht/Zw90jb2YUMjfMOPp15gHRAGhAWzPyrKSQSrf6DicACoW
jSU7tPCuEka60hxOPX06M+mCBuTRWuSjoWDnP/o0+Y9Euu+l/70SCQtMPf3L4uEQ
sAiTmOHcqNb8yA+5M7efj6/vcwJZdzomPNBawca+kq6AhAoJ6iwNZrkCh1N4Px+R
+aam+spuQsvC3KFZz5nGsBDx9+TAaB7q+vD/2kzzwnXw3f8osPbG9uNOTGv0aX3F
O3h6nYBFjI4z3xct1ewR4Nvu2Q2LChIXDsJQ13xjSpEwDYL15Meh7s4qnVxm8hP8
BeDheGNVrWcE52OKBHgoUbPuW4Lt5/z6pMQccWLEppCq6l5+ZwFWQ0ff8LMVD8rz
c+g3xB7Tqy3PhkhhSYF9nO9hLfULz/b3+sfJqpR0/qL71nnQHD5s0X8RuPNN+DTT
LAkTaSIQh7OZ3+3Hli4T+TumRZvUrf5gYBfW2zkopuNrgFgd24vL7iifY+MlHeBz
66jbKYUT0p6Z9qNx5hn0QSwGw/SG++LBcNWr+MtqLKBIzH35o74tl8cPHgQ2J+nI
Fxd/vpQrC6Wc5bdptjZ2LJLSrHcHWOKNzNlz3KwTh35KTS0UTKYS6pIiavnxb35k
ZfWkGHJN0bysr31A5tQ3X3lXbkptCFJE0yNFH/8AeSiXnAeaou+bXSPk3MTgUUin
WwJwYdkHYxgrR5hY/8odJmvK/l05AtglSUwzd+8edPfEXbH4KWnC1TkulY6xwMRq
6NyOpdBjw7sCVyTXUF8mGeCheSgAjI4OXQ+I1OOi7N9sSL/W3URWz3ElCkq4axk5
i4h9QGOvEIkQF8yNl6y5WlkjxSQB/w3DMwYBYRAUHmU57HLh8OmGY+rVc8ObuWK7
D6Pb92/fB/P/Tggkkwb2KMgZpzOFn3xSleCRrxtAgpLnWGkU/nYJNzaFlSyJ7HUl
OTHEg3U98QAHxPLn7XLaeDc9kVJ4BHV9Mxo7mp67QkEgBpsZed+X6Ukofo8Km7T2
lJWfMMRp/zd3PHQBIrWPieUhLDOXqccKH9yzB0ONysT7e9JUZ/naaPFlS7WVvbuU
CoenOPzpUg44p/NZLMrjMDlUuGy5GmGFXmemtvWD4HrLc3Ela0Hl5aCJ0QBhcMXd
CgZXvvP2WDWlrQW396z8r6gMXyD4z3pt/Sn4oVzHzjWX06o1ZpFjDkKuvOg0+v3e
CKkDTHKZCegNuIGgJMl5KXqm3b0cHrWFELUWuVhTAMN6ClKwN5hw9HmcOOjUSI47
uoXgUXgVdfPDz9QS1MiyE7FtZSgVcca2V8tMw+mykpbNEMpf5JOoaheUEJEoskLd
eLrIuzSJwZ2nd4yfamx7Q3V4NXMCVinlX+CXuBduVE2Hg6lzLThq8McVKUgRnZI+
8FlAuQzMY4ZbvjsAadyrgFPN1ET+BoC9B0h8VXVarWEEwXhcWvoc5WReGhD7YA8w
Ehgf6+VvK5B6rho0vNjO16jX6JBsgvitkJbK+IiUT7GODGBeWBLs3libteps/v0G
RIznlPps1TshnVwc1xjb/HMw9xX8hzcuoA6QbAxd61VXPCPC3a3ErmZy2Ty+tnlx
zbkZEoBmmfc7o2d3OgSM6mIx99EoCvGDUz9T5I92iqmur163vSvM/RSjR52Suzwq
c6ANf4h2sAbsoTdvQT/HyFSk2mYo4sdFu9LRKp3+OWd1JEzZChuF1fYVE9W85nTv
k9JilqJQQ7mklSZ3WQxkZyPBwiQCXUSY/uSWEY6jn36NziWj+zsM3yDYt/s34Qo4
pA4zg+FDgojhNJDB+NFdmOVXHBNibvbfyAmTiiJb7ZxUKaLyjPnkcLZPoIOASUzO
wNJXQn9gBGX7UfTqyRBxsViL03y9lQ/bQi+5KfjbTa+dGHGVBhO/LVV5QhigpJIK
IEci5rXV26swxSkH8T4yT6tz5NrDZxq/3tmgrTclMhktYJzACPxozQEATwnJJgw6
XllNIBGu7kbOkiBo+hrML3xJ+7JLbcB6seaodyt/ZlFUZBbNHTdPBCcc/oevIHMw
fYT5wASEIJy8z7HXJf6YYkae3rmJzJM2uC19ych5oGs1ElppBECUDKVDcPcRSpRP
GU97BjHf1Wp8InNm/Lclhh0OuZ9wSD5QhUerN686JPP3kl+n34p0mjbyb8ioZerd
ACPFteSDBvg7+YH2DEeegdUQuZ6bPWqZiEMWOjMmheTr1sD60aU8XWqTEfXipYLU
gkFP9agghTlb82lraDw4koyjdwfjSTMYFEZBHPXXIPhR9cYlx9gDnvvRYytLLygA
pFkCQEYtHSHV8oCsehVbC3a56+vi6z5XIjb0+ZvUUbV+BLzP+cVCVN8Qg/Q4jq8b
rt3QTefhVZagJvy6CAxQHgRVepNVsL9ckeS08W+LrTDu9DZdsQ0b7LXzBlgmGrqG
cQJNqJeEqrnrAOvLZmYcIb48nY0xZ5S9YzkXvaN/fcL93kk95TELICT91YjqanOw
1EJiEZ02TJ6csU10Cjq8QHuj6a8jU7nXQtBKTx4lvvpNCE1NkYGAhnfD4/7A1Cg4
iVL+gNK/LxgClsqg1DHc+B36kqC+p3CCq34QvbKZAbbBoUhtgaZIktNOc9W9IRL4
sBGhwNcZC0EI3O+fcNLIzxC02b4sO6WcFcvoOTijcwPn7yAhnqrxCIQi6NC5RDvd
h+GaXc+2uqplQGGKTI4dJkGAUggAq/KlWfjRSmwdFXM=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
QHmjfy6Lr2r3CgpASAFvlrhiAJt/Y2G4r/q89zMavfDGfIOMaBf+Q6KgUrHgO02m
GzcVwaFYHnN7mKd/DVkmupeRtPDPgvGNS75kUPZFDJRUhQ1PZFckLOM581Wxrq9T
t50UwFlo4l6eWb1rZR+bFG+wIxOKEegrhEOjfoG3OYQwFyb7WvUrxl+/jgEmsmxi
iIUa2gLw49KStLLQu4Bwb25aVtigp5XPIa3mgsglF1SXY3QowkRV2KMe1ei+taDQ
TlyxFZr+98p5Ud1iu7ZLVDECLsfjR5DOGXYiNfaU39eGznvKgT3NvgFoUGgSLp/7
wT2p8KwRMwpWHURaTDhoUQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7632 )
`pragma protect data_block
ukg/3+aC8OgtSV+t1LPKzLzwGHPuqbI25tRiwBx/YH+GJMYCMcJ+125qcKWlSLlK
1zAUul2RFqWInrkRlflCBQW1Rx6MYW6jp/a7LN11yUm66J8AhR/rE2XpuSIYLvPh
GWTrHr48ccIx3jGa5eXeYGqIaMDoVePmNuJTWeH/ivbjdWr5p6+OxBWw3rtJrIe+
VxKGYV+VN1rRq+unjHVWeAk3iCn9fzpSWjvDhSJrQxCKAuQqXMqTv9G92iOxhtJl
+n0XMT17e/flbwjGN49pfET0cLt7yWBO00f1778OtkrXo1XGimNQm41m3UXBdu4+
bXJSn9YZHMzffSBlWEBREGrNakmPmvQsioqRbk4VrDks5PYlCt0QV6zz/ljXODQh
MRXnKrlEtgk6vqMon6D4ysyF5AD95wf9cwpM9CIT9bk+g9kY/vDgcigJBWNxAgI4
PBj/TTuExaEfmCO/yCQuO5l3Y4dqTtoO62LWdDcjr3nmKBG+YnoHzg++gxsfDApE
bCkPviFjQ8xuUsTpi9zRanL+x+DDF+9qc81lL6KcCU86xA4rdLeOvuSwGFB8LJgE
l2DDnTG7AmL8BCbdGK0/B3CY7LvpmVtvXlSQX10IqC5GsRD064Fqccle/neyF66M
PLvXdsofjXRWImQzlKNdFRSQtTnw+IJYv1eSsH3f9Aa0EQeZIazWmJcQsd3QnqEI
71HoGC9zrF6Xg2Dd6lQPl4k2OOp8s0Q3Qj0bMLlgvGr/On+hqgR3ZwX3OpUUUcW8
PQ5hoiflUPh6+2w06iu3XYyIN2ji4ASNpWBKGFIngwyDpQ3ySVfUxbRkNdkV2uUo
7F6f1+CCQ+LVvd2BvtdoaBsM54TKIsWorRQpoM0Q3zApOAx6frqICUEApuToneTC
GbL3s3zBPO9m19d6152dqCQWeQ17uU4BlfCZr5ePd7RUuts2qJ9WB9kV40jQmy0N
A8NxvZaCIVgAfNFnalDEeyYxAHVuBJ2rQDVtN/XLMizq7d06HEYKQzNvuN+SFC5j
9wN61Chm2lmWVEpFJEPcIg1b+D1mmVj9Ir1dX7ZtYgh4cW96lOnj9GT6woiFue4e
tQ+4/3qSjBd/TqftA3fHlaT8AWIDyOzg2kY3C4+sYoWyU0/yhomLLgaFCPbRSEPl
+MTctv4d2Ieoz3ardsSV4rXEJ9iCjh8dARfd0hozFfHKsHNE9w7PAnP0Gv5Z5kxM
YtSk/stlHJ4H9UW/E0wgbGDhplUe3PXl6T6BVRp6GFQJ4MyDmDL8sNIS+oB4D4pw
QxjxTlSHdWn1L94PWxdH8cixUpsOK1GYj/9sK7YQKDfV6zT9MdC7S7mj9bYmMtlU
5sHViZQpqamI2aJkugTPmhV3AEQ8LP+Oz/4+x0byqvkz2gB5cr9JPXrdKAQ8MeVg
OJE2qoxBpXiCEwwsnGgNMjk6lnNoJBsmYgyMomZjgM3zG+HxXNintrkefFGA1llR
wBIhsbHNVv06izOMcSPqD1xIOV1p130q01Hnv+6TqA23iZ4e+4fwTKbaklyoSIw6
m7Yp3VPcNq5z4uQhtXKW/qagSHFF6Xcap/4qeWeTU+O6BVMCTkx1jhIOmlB4FgFq
hqLepZF5iJCbNkYIYlBvj9skUBtxjzbiG84yZXRl5JLBDpB7l4Vou+ziTWhWzXfY
I5BEA1KgCpkZ5heuxgy+h2QP6j4Hn8zapqWXqQWug/DGFtjBiNiwphvt5YKOXa1S
N2Dltabv5zEnUGEZlNpJO9mjqBK5LAsTO/o6ZErn1TvqQ0tWWWhlTvRhHboOVxln
diC/mukjoP93NyGXAFAOyeQmI3zxr2CcNpUbIIZK2grER3DxFW1U4DEIFYp2uLEz
Cvyb3WTq4kny4Y2Fv1yF9b5HZw7HdmEw1eOJCVMUK1sdK6xBdezBdpNre8eAC7M4
j2z64keK2a8JFsB1lhPw7n8jT/prL3XChIZB6WNp+m3bSKqDCWYgJAWmsp3Ey+EJ
HIixL9njmXC3eeDONmAG2jKdiWaWhY2vRyVujSwZHl7lfK87bbWjLmEe6hmz55UV
sKFn1aGe0MOQ6Y1Yj0jYdnQPq9zsB96lKLVf9TEokFYc7JjpYVkrsMNSk3j+m5tZ
2uYgkEeWZQtWUAbcqv66yWWNVfstag92NQMVMVBNUUMwPoi+yWi5bIreLHpftyy0
MOmW8G9i3fCisukpb2fBw47olkZ6FSY6eEiHLmq8Rnk6/ZLYLRgFEMv+oCGPpdWZ
+y2+MhB4ti07vSsGK76tcSJRCl0Tp82acEckR2gikWZwDapdfr4C6kUyfBwbyfnK
/I0AmiWKZBaFkGv5ljvNFcKWBhpuC+5+8nUS0+jIC+T3wJVx2893oUk/+B84WIpw
SOCYugex2W1+n7yGJXbHc1TzqJIuYA2LbKHCkNZCYFwUhFxlYEj4Af2SLWICGu0v
0T89XLXinCyvbjXshBPw1auKJOCWDbCRz8YARKabK8gU6XWadi5Vbzy/rmqX9s8b
38qv02S/e5rnNXJdwObqwENnkbzmSQCzTrS6EcIoSjle5JTAnauH/M2KQKab6ZDK
4Ytdxymk/wCNMIqzv3HL29it97nRNkyTOk6AWQUNJt9WmoO6MzRgtVHUw2L9UmGx
YePfM46/52AvW1aaewRcK7dACNoEkTAH+/Z104EnFeJoYE7gqhZpVfQ3Sn6+fdxY
qDytM6Jp5RKMUUBlJU+9iBHv8XSqqrDRQBu042AS4QK6VfqenbT0fiaVh2LdXQNf
XeQ81AEcr63z3m7/1LTsPQ/jjZENr8M5zC7Zm54QVeytcD+URCLgeGmJkjbyN8HC
8KTe+Ln8/hvqTIzOL0S9+eeTc6SUbVS7J/7Xq4crMU0NAMDdYiLH/5pDuYEP8Lcw
/NrG2l/o5s+xoyAt88qQtxCihpLpl1QVJV+sF7uQFDLbznGx66y/Minb9PUxytyt
7J8cjXZrCheN48SuTR5f9bua6PyrPYZuHLEc2x0KbprHxOd2jelS2xXW9vuIRyez
sS4Oo8023KddfHETZYTwGudQM2AQIrIf61A0rOLbx59qcZxKgHcTmT9N+wpAZpOg
5qLgEVn8geFHNLDHK8bgG3FE+laD7Y+DoiVO6GxDO4IsjZDLs0p5kXj6Nat+ahM7
D5WTP8XV/suVwqvGQH+Hov3V/W3seC22QzIU+Nml142oUt/Tor7bmRuCkMgUTg8S
sjvYWPQBdpQg3yd52IGOKhvy1Z92GsoDOfClroN5/c/PYbbm3G/e0FJwBipUkODk
rJ/ocFBBRrNFeJqdJe/WPzhg/z9R5Krxn3a2eM+fu1Jsu1sSmwCtE2pW855tX2oK
rg8BZq2QwTkef8KqQcK8xcImTDC9UyrULQPJOWgBWRQh16E5gW1wSUPDvha21E6b
FQAMlhH37rYjwGqRBQ98CNEcreYs5DS0bN4PeiIbCTuNB4SDVCq7fnphV9Vc9fWl
Y63YBY77pjxr5jKTuzSg4lxRw8JMOisz09LcMiQcj40pxUymHUKS7YFD4K48bSHz
/shgjs/i+PXEKWh/ETO/jSm7fbYyf7QxAnOoCvU1cT9cKgoynOZOmgpmQVCW+j8V
rGVsoTOq3sMGtQAke7tmOvI2XxRKDAx2iY2wo/NLyrshR9ZAtq7ogMX+Kg7MyGCs
AG3rshSiXFRAGUa6YmYFgj6Fn6OCExXgC4RcPXlu9lifQ+SxQSvxjCQa6VUOHWUK
XIhoE9he86evfOvRfEuRssTm0PCmtLsF7fs7xBcQbS9jbzmnFLXk7pPxebc6CvDC
WDr+SzVXn85NIvGLQ5x4tydRtKK8+zIX3RWh+ahe889J0tglwXIIpKCjDKwHeXUP
88ByEXUU6bTsBGBoAegUvjEWpyqVzRDme/i5vTeUelK3Mj5uAVUUbZaXBBG7oykZ
S90jm2qh6jWC1zYpdoiFfKEhcZLck6ZR9ac1osrunJZb5RS4qJnxwdm62xWYv9Gx
433rXnaP5kKe/KQYajqn9DBpShrDdJQR5Tvx5wsS9fIrBBx6D4sXLcONSmF9/TLD
RaZ69nBy2QIFMyqqGre/lP0V+pH0BJAYUi1M07xNIhg60bj4luYoftWsuitDA2Fy
3xAteETjyTUD4pJKAey2WcFaURsZPLrPOPzJ7sMMOxOUXBh4mlNZM0wSBOxUVXob
jwpStzQ82FlhP0wj338QtOBOsLSjEbuewZ3SsqTaKapLzL0stconlt81w9gozJm3
fVGhUCA0fvldaZbubUamEOPxu5dbpSDYuR5aY7IkLp6+V7RKhp/ImS+U9sdEdmVM
IKwwvJr9zHw5qgPw36tze9TqVgDrk1v/gQndKepFypuIebayy7zaDgR8GbpSsYZX
NJQFKkhlqWdRIObwgJ+/8KD/ErEhfsc+kYzNF21Snrh1oq40eLx+8Vkyp7HdTaVR
l5ZTiCg9XZjQTOCJobXLPm5P7U3sVJZJa4/985+I+Lvg7WAsn2jKUkMmAZNkGCVM
JaO0/KKuBrabbc2rGNmZwB/8oTjHHxwsdWp1j3kjQoTkzVHVP25GTuEj8ySd/v6e
0zyVFSK8T1o7KazpG7HajT7mMgoPG5BJHfn0lEe/arkVdbSvDDERLaPPbQp4eyT5
cF3h9m3s8NBSqYnZ7rFf5BreFYulW27en9YJ+UwnjFsQXuwa3konXvJntVPxs6pL
6+HuAMlG1pwLI48BQssMH2wCtYa9ZELBhcBU1SBZfnqEFEOK4HhDNXKeWvTWihG7
j7Lk8s/Zo5Kk7UYNFxw0uj4oYM++1NcTWD8it55ssZJL9hvw21AO/XyLbIMofn/G
VO6Wiro/1mbHR4qgk8Kdwg5hLc5Bj1m8IzukMweeKz9NDaP6a8H3+ar5bsmgvYhq
sqrB1ENyN46IUid93QFkwlFyiYOKxX0Z1pWWBcr7yLaBA1mMBgVagbWryf9cVdIf
BOxw4AykubSnCUx6KA8GbAF/H2zD9X74i2kOqp268xroldg3yI+rt/J0ygnh6Ypl
r7hyg9K0woGh+5HEM58xTpm7ryxK8nmWlF3/SXAMCbae7N3PPQ9F1AM9wTEaQ8ug
OcI7QaeeNBQBXtsZsKk+63/6nY5Ii6gDbdp5yUaenzXIB2QarnXVGs/L+kMeK+d/
16FruBL+8cdfaYY5AVJ1873mpNpJeKph6sv09k05USpXEtQBxPTw+1a476z71VUa
DsxqBZYNeg2bqXzLNOA95vsio3G4dmoBTgGkWzN1mohhhpoQsPLhjphtV8FJy33X
prJQlm47nJntOjCrTjDP2MgD3Ly//osNLCWsSmq6zX5l0qLgpQWt0VkQzPnYmU4U
x8Lrqf5g+UBH3DptoC/0L6QQGXSfvcft6gQfv/Eju7YCGMzKBKrcgQsUeZ/+cntK
nemwMvcSP+fKHvWncGynWk7hacVj5brLEwMK0B/B1q3NssRgqqhiD1HD9cZ23yf6
tcNwi2WItivdvsyuYBLmFmO4CVXQ6TLoDWvxXPF6NaSoz8tJaZDZlxPkTCPG0N8c
xHolmsiu61TwUtUaP5Mj4ubHFE+unRzyC+zkIwYc+UHNYyN0OIzK4JZCgnrXcQdo
DfXvi01icWBo+XiM51s5mTJQr6R6BwXzEjJM41TGyIH2DCzAV+hF01/4ugIog982
+5s0HepFQly/WpNA/QSJGo2QyV0mi0G+3BDrEhsUMADPhU3y60d18i8obHphc5xe
zu2q6Guh4rmdKpbqSJa/VLimnACMkVEsSc+akn+L3aZ4Iks2MHwGPSGt51KyJX+Y
7ByI4tkGTLUCJ0CeDHNz1Jbi86Wp1PaNXUxvlJP4hRnf0MTxJnviFvn17ryeSAf8
f2XboVnUoyM8aA8YXpPAY3W2GYQCp6japHJoSY92gzUj4QghINtRINzaHj1K8ocu
HO7x37KQh3Mgx0Jwv4MzQNlARiR3zSE22wqFqHQBp+dIwqxb/OCc2c1wKbhEZR9A
y1WU6yXoQoVXDJ1kih1C449Qi88NRwsBIWwuaGkT5D66Zfyhtc0jtwUq7by8xID5
UK1ODp8+ZqLkbthc5SP12nofTq/+vmTRDEfLtmCIdEzHvaZiBfoqDHeyQ8Z6Rn1/
LBtoLXUaFd6NXnpN9J4b91PhRIaVS8Bb3YhsNrdn74VfybSKZMroA4VLTiTf3/gx
YC7aEJNXx624Vcg0XqKoD3c2tLlYPrHO+q6VnnTCrF5ubj9viBi30UvZPGjYbcsn
4K/yDx69IZMbSwMcgKSvTM0bh9uZ+sQgCIZp5jjreGCbdzuEbbTR7tGKpvsEhBLq
/jJRmfcXoKc76Av9746VZSa4ft3bzHgPVpDXtT4wNcL830ZFeHr5nExSMmXP7tIw
XX3WuyOI9YcK1dG2K+pL1P/xbNf2E2MAmwh2h1g5BOg6xhrWrbDS/GepHOiItPSM
v02v2zpdz/Jn21/hJtTB/jwYWwVqmQ2A1j9meQpyeDnnyLWghrB18XKn55BBkc0C
7mGA4SSRQwEj+1YX8sHHC21mnlLZhpWCgkjrOxbydsfqK8mzM99MBSgRQE9Suu0k
RorTnnRLFc15IxAHH1kJ/gN5R+tnYW8/f+jnRBI9i9tNrRKTEu61ctSNKNolAeW6
/6oIyDkRYOziGojqzfivKyLvad0+QzihosaR5QcrF6sTkYD4Y9X6K06Ns5pSkbUf
ln+qoiTjEHErZKJ0+Ezp7knrnE+R9OyjtMNP/Ddsk09ubfkbcbskfwNPw35BcLRd
fnC6MpX2Ea0T53GUk5jHJBEzypRVeMNByj3QGPOxqadC7dQMtF5mLDUSCr+hH+Fg
ZkipthHpHSy1J/ew47Sg8wmO81jRT2qfiycEdnmrQYwNMMJLgLi9Xalk+IdGcMst
ve6RPYQh+OIEwQmVYjoDuZfs5Bdc4Enhaic9NwTkAYUk4fckCDph4E9eW/Op/m/Y
aaNL6vXqgO0uUCOzM6tAvwmqHB1bOFpDeVw6EDSTXQmScbahIQ0gHUekbWHILfZO
iDh5oHV1i5WitLCusbecVzMCh0wTl7nw7TAIne+7smxfwEc9QDZnXn5a+D2a6X/M
wlE3MF2RLlTBCy0ymlY0WU7aVeYicdQdpTWhz1Hj6LmSZVhKzAPZtnilQOrqH7jO
S1jlf1Cr23dKx70ilIDYb2wtDkf2GG6ElB6gYI6MM64sTymrc/d3z0HZCEvCdNGq
BjAmWs3f7p3xm2YcV2vTHetRDi+uvnHS41a5Ri/PaNRvsh40szX//VGasAtyK8ny
wclmqkvqjoSQR78GRHBXH5aOcokoZc13ExxCM5FXZxcZGli3TDi3DYRSPTrAJTQ7
GU4hd8jPhijDhjTuZy+rVMRzh9M+GXpS4Si6EV8XJGGmYa4900+Y+kPYFZMIZQRd
XP/B1ok3bg0Oxp+UFqweW4RrRJ4s6LpPfLAncp3lpIjmjAjW6eDYkQgYPJrr1xeu
V3XsRnZrH1Z4ceUlIPDfGlfKhHibmDvX5XXsE+bROTJpiOAGJgKF5cq+MG5xMgTr
oUvHo1DJNy9lUlSYxrrFl7efLC7V9U/NQYI+MZ/HkFa3CSrrkDpMfuJ8Y29fxLW+
5wOsvomk6OQU+vHz6Wn/E9/e3SaO6fiY1DMYNdWhd6Uy/n1Ml7NuCTGLNqSFbICe
lR3Rm5fakOqC7ZbF5A3xmrfVje1p9BfttRNkIt7rRZ+FwDL4gF3sNkf+xiRAEhOe
BUccyjMcIP1u6mzgU/sMsj6Q/9eFEpIB1TuBEaNWQXMUUt+qa4WsFHrtyYylmPMK
HJBG4MVXi9ywbZ41vpqvKEQC1+GHLDcYrCG0eXUZQil0uSFXLubGCyFJBnyTLP5s
sO+l2I7vGldIOlaPMzcKoE4ox36AfLx6zbEn40E/sEKvN9swmj5xAjvP/e0l/SHv
J5nEn4dwvlIqyEIFvgwjTpTr5N5+BiLqO0rrtzDCx/savvZtJWkz4efuwq0BlHHa
9xa8j8CvgBkikVu9bP/Cixe5QQixR4H+tDQkosL7RJepTXcvu43W+nRN4MLP9dV2
WDP+RIZEwshL33LFo9wSwk+oR6xyNlKGUW9F5wLHM5oUIFHon3t//rgFuo3Q02Tp
j0JfzPMlWpwbh89YBr0WE5UkXPKV1AM+81PNM7g6+G7aWsSMazAW7B1EW7J9xhBk
KxIU0rMhZ0WNzWLd3gp34PyPexTwJ93i54eNNbK3YbjQYO4MXwdOxtaeLURHUI/4
7FjcouG2S/lpvRTiJcZNZ+FXHp+TbPjOdj0q+LyOaO8kvv6RKu7tgnWfWHFIA5O/
6UZpmNNfiz3iJe8TFen/jPa3CedH1dH1KmXKhS0W1ot0Ytfc081DenGtU8Y0mpdY
+bBOveTHxigX0ekqX2NW5tMcWC7WGWdY9zADuZQlmbF/HaEbrseNyZ1c0bZdjPuz
Di9B/P7UUpp1+58HtrpH9oJJ0/TXG418xdGGsYsiKLnffJITGFu6xRs2FmukINZQ
VjIJLPIq87Sb6nqYhNKjYO5w5e9EwBz4yOWiIjMrdajff5EdiQdlP2u3mnAVpBs/
HeaTepu4WvofEXwYW2FURVmUlo6fKDT/DN16Z0hzz48VESsGVMaPDViRk8BGxDf/
0xenpwrd5GKO6KClrjOZ7vUNF7NdlZgrL303AOyS0NJ3DKsljMCyPzp2LHgcyOan
tf0vneKX5HwoLL9V11782HaAxy2STx/grukTnz57IxmB5Tk1XSCRphpwzS65isxd
jzX045Z4zgjhI8z7gDsMhdGalO21R7YMQQLqYmX37v/5VEfFiSn2EIo71QuSrWk3
+Z9EMpXXFWFxhCZyhbyrUmesHuM4CXiFX8SCWzMbr660d6fHSegSKFUt69Z9lfkM
n+WFANNmXO4YWWzRjp2+UV9hHmm8G3veq6lfARRph8EyWBixh9JdNxqhhQ6WykTb
Sg6jNFxlP1mkqvp8K9zbAMIiIE+JXWCHdn1usQCd5HfFIzPIcBiySr6Qvx1EJEqb
klxmnflfZZHDPAJ0Qnp7DxmdB/0BSAcDhnXXF0pWSAVgM6/NMXi4tlx+M6+nQSpo
eH8I+UiA51jPHpM2MlkM+qBGe2i/L/i11ryrrggIjgvBF4AhgN9UQ/bSMCpWcjIM
6SPV+Gcp3DBeeUHO6VVRxrCZb7J81RVGi58GZLE4kUbHbrpv5jPIBp5GZDE6Q4Fr
JaVMZf9djRvRKZDzC7c2oN09k9Xe3ETURJ8mHp2FeljIBhkN3wzlxKuPjqpjg8gA
gJ/NUsfA+2+hclI29qbD4EqRYpOya3kt9BYT9qw7TWl4psaQnyypwotjXhBPQ6tj
DxrZlFmv+RXL8OByNODFq5qsbkTMTizVt/copVQBEIIX8f68KKiWYmnO20hucOkx
HxCxZvvzUbTssFbUQY7kJXYPAEqX9CJpqSveDh7CoFBHWZC6ZcfJ3Z/THPsRShla
3XhhzuTdYKGRS/QPQhwFXs9YfohHMAm0zrjlhZmmRBWX6klIiqEEfkytJtKlUPid
IjcbleIoVoa9iFQeE5pKmdiWXlquIsMttb/8B2dNyq7BsQ65w+hnzVXtGMiiA0pG
AYwb56nYmWXmzTo7DbBIIZ43erh2UWMar7YO8Dfxz+qTaaDzoDm5V69AS03rrhCx
cTwq82EY9aE6Qq63bFhJlU5OPHBoFQvKAkM4gkwvjKKZHBYwzB2PBth8NV9uCK/l
nbcS19AUAyG8uZmDVUquttTztyklBlPbaqKr8MNRNkdcZCu/K7Wti9aeUw+y5eLO
GPaXcTTMBnrMsIK4Ai9ZEL6y9xAAmHg6av11gXE1TCOAwSkaUjTgJZ5KywrRHJyD
5xAyC9pwI96OEFi9H0oK68EzT5PLnKBIqzp6vEeqDeGB//HOjc4KBbHZ0MIGae+b
3Zu4HI3RDOuhvXTPsojzpMhktJgu7gkgTjADR7i1z1Tt5plkzrLO8AdPf+2Q1mES
N9LH69Uc6sbKE3Jsj07YatKJQ7WwCEHxzs772kU8XnTUELyxVTjLxmQEzYbA2u2C
+Kn0Eq46cdsfoRHH8q/34ahIyiI+i4Lpb3eqi7cudTVpgVfBxXMXABEWO4MnnYPk
qAz8e34C2sWbnh9QoTEUVl8X/oPXBZluwQqAo+nbDQq1zbd6cE2Q+tO/C4J4DX2k
NCL498isfuwnraZ1ectHfp9MjMNUMg3Ul6i2Qah87+kwSK4Tk5zwLwTkMcAlbPUZ
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
biEbQ4zY18iHRrgeMdN6wumszJKrcN5IBtyY8idlMMb0tTNZGWr4eJZDZ0KqfwKY
RBW0KfA+zzBnlI2KT8vqirwqY8SShO1KBYatwmtfqNvban3iEVGzFXct0L7qNwff
5QbBbJriGlO8CrMTHXcLgZ33Ek031vL+4YCoBxiuDczeYXJCSGzZvoRXko7YiqLx
5CuHzkqYqBZMKxlS6pGtBRnfayukRRsttF0h+rfh0bnRdSPeXgCMMpGyiCmfxB1X
3VKhCay8NBOtQhqAT4XIDI7iFhpmUwTj0DulAS2HhuOcOXfBAjDtf1A7OKgTqoY1
i0iRv6DFKrUdJzCLqo6PAg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4768 )
`pragma protect data_block
I0dIrLswVd5SimWoaJ3fdLBSsYek7b6vpZYIW1jD8d+vQ2BQPjNn7uNHzX8L5EkG
rHJmZfs9/zCRCUbFUgK7Fd3jyOKWxM7xrdv2tJ7WnEVbAqG5aKm/EY+iznVSbHrE
p3lkgu64tna6ApL8PQqxBikYswtQTlA45dOiyiEhXaxVUGEFbPtCvoN/8tGfoxSp
F07KBjFqVQFAqKV8/RX1KTbUrdOcWyEoYfx/DiDZ8lgOpVBBR5iPWrl/liNaOgxb
qCtgw2XjS0trliC6p7RxLoEC/m0oaI+Wj0yMUXU6F9D0j2QshmsPH6x/j5/Sh2Wg
kWsblwCuV+rf1oYtgQ+jJOxTC4cjgzBnkvdJaTHLfIfKU08O7zT44HFW3dEsPgcV
F9rilGysZIBRttp05UcXq3vatL7JeIwPPigutbLqckAw6heaTaerDWkdMyrLCs3m
/Lj1BJzYuKp+XIqz5/cg/GIopAh5Drg0SAXUM2Z2FiMdqJB0zGEkCHcZH9Zog7yV
NvLpz9k9RHnkcHAnsLRIPRkef4ocdKAOXhaIY5R8UVmkibRFaX/XtOeqf7Pqfscg
j43XWHSUJ+/rcG2ErzeRb962HP7QNpH4XG/d7wpDhIhxI2y1FmbUBHNSRUZaA0kk
udfdcb+8UCq9xND0lBhN7w/6tO64X4NUcleO4gnJk1pKoPtklCfpN6boe1t4T25/
msGv3Sd4UFUNLKFVJT/xYFuAqE/HHPI154Rqsl1BT197jeLCxyHBE3XlqA5SNiCF
r3sNGR30NnTiSlqqSO/kx6dFneweCrxxB+QrcFOZNV0RJtXdxCiZYbdWTsXUrfrh
2aif51nLvbelRQ3VAkRtibO+RqxMMwEbWItt/SL4zN1FsduZpMYZNsBi/DbrgjBk
U3jl1RjatRsrmtryn2VRABDxJbJHtWqabs056JEUcthF2kBjggRRqXh6WAdSKWV4
t66EPy51ZD4kt2WAqlARhiYmRIyiu2MbXy4hwcVEQCYgMazmZ7t8OKjcU67PZJ8f
10Ky2JUkZ9gZpUQaL3H64xDifmXTFXzLZ389riObSC6qz08DIz9ScvqvspwA54WA
w5ujpxwotsqkel1IEo5jHsP0/LHQ959nR3+IH2NgBivaDetcfl6cD/BlSB6ZTzHE
Y1ah06N3av44jVT9V3ChNX5gmdXj4BY9/IcWHL57bIsY2Y2oAXNgsTxkL5/Vtv6n
+qJIQ1w1uqL/QXKDRr+s9yqSe9lNYiqLcghBROgXyPl2wdMp+pIeqbD1EAgaBLUU
7xcZP65LsSynYs19dP8vsJiPbSSeDyogL2d93W1y8kKZR7/bQaKaX/Df/8TuVHV0
jN/8xL1scBibuVz4w40kvSlOe9KVXbZg81Y2g6QDyoWcibDOpK3Vy99LmFI47Jop
TDif90R6KqeJdf6X/AFFyvBS+I1zs0IvY13WmzywWsBNaFa4eY68djFPGp0NhCb0
Bwe95bjEzTKzzz320azH3SY9qH8DjkANUKuSAvWyUIYo8njNdDwq1RY5pfLaam2Y
xQKoaaBplnKW7PHv3LJTp+9H68b/tJpSVs8jGMLODCbKJC8FgvQFGbJDI1+K8Mba
WiuPfdSmydeZ6mYEbCEUb9lI8j9hd5DoFPr8fg4MgRsulWTC7fI2iG2ZhYcz6ex7
1RzeFlj44zo3Vb/w1nC7jeX+p/2DJCT9rPXKBsyOo9/BI1zWVDgsp+APTcO/sBnc
eEKJohFfNkPG6REXKZCVe1ConhqeFQrMCVPK8PW9wQAaZAz2R5mHDDAI2MOmurIF
TdPINN7ZFuoKUUwHjvWjw7qb95BjFk4D/l7U3sSzVOj3VndyJ/AudE6uJ/isF102
ubldCUn8A1/iIqa3xxF05q+9NmEF0LVj6bclXGYdDnBPa3SMIfwXwjz+8RrgdNvK
IkXK3ec79tjGaCUtr7yiZQdCI9ZUbL7X0iPrsymtqGs00dXRF6i4a/8j6nqt0zMq
sXNyUDUWOgOLT3OTCrjtqk9o3PvmOoa642n9CzCMXCQ5CNc513plRfWwDmvBNv45
DgR8EIFpPqABqxK34arT/iKlZiULLpikwjyVL74lquQDhHEfBT6d1s9Xd9O/oVU4
3YMJRhDeSvparusubTxqcKnLpM4DWQM/uZTxPEBN/aBDyvBIt9NiI9K+fEy8cAsr
MU/pVizT+GDBYe0ngV4qfVv4EZG/Vup8F58vyglhbMatkT6h0RQWCQmPB0PRIb6K
SvwLJ7GTiEontco3B3eeNJKg3KCSLeeUEKppKtbOrGS/GNFMPRy+XF11S51oEjdQ
pwinF2/uGtat/WgbnFhT2+EEsC4eRx5EaZNAzRhtsjQSiWEgjnLmHi9E8NULgFYX
cFpmhEKDqG0OIfwGlWbNm/ldIFo9JsyTNlnEy+OZatYwGGjIChpF2b3q7Vs4rkTk
cnmaQZnJboe37ZZP9Ri+bSMVqqpjXmvDV51qRRoYkTSH0RMmlHqjE7eGQyB/PGMl
QV367roal8Pz68Vm/DQR9Itu3eysUoUFOff66qSFmAB2/v1aBY2fNHowvZ/sXam6
DbofV+6KAiik/npLO7py8FWfiOxMGZKFY9qIwPyU4Mx6zjPHVIwlvU0+l5aQX5Z6
JoMZxAFVjlNcqM0W33ptD9LXTQeDzgq9Gqt4TQv2RaU/yTHVcKbIyYcpsrSkYUwL
qYYJe1++9i9MkOgCNh9Hmtxn0wWBeBbIa2Z24moMJgGeb7TOR10T2ubGtJ6en32L
EYUZtyYgYJFu1cL49x+i1HCjkmpACcpMRLt7gfQ6g5EPXpGzdBfdhXiXccZPmSPY
7g7bcCqUOxKycNS+HzqMC0wXw8GWG4coSr9duTfS58f4LLchasFWxwbxcYyJtg5x
1dn2yFzEBIIyTNkqCWkE+M7KcT1fvw+1eKUCm6IvqDIHK8jjhbKH+KsfkxHVCBHQ
3QU4I0KPQbemKanb+/Y/wnMj+1UQyIWZhznPIc0S9Py6BiRW3/TmyRbLb2MgV8Dk
msLs9fxex97W5BPWA7HqM1uevNwCDg5lC46IgODPL31VAiw3/oJh4yF2KSom2YaH
22H6TTi7udAagI7Q2LSYZGz66B/6fC3oBhFcHyjCkh/FKzrNSkUB/c1Rf9ilU3n5
FVXOM+DpEarWjWVcfEC6FAnpXTPX9ciSGQA1oPkF9Sz5k5ezpKls3aCsqVOoWzdp
tRaYvwGBEhGp5SkdYj8DykZqeT3Cvp/m+J0oevKU7T822y8x7Hxf1s13Ru44qAOP
V+BkQJajwckVIq69snT58U/jQmgy6eT+3umTkiRwQApMhz2we6d+hNcsRe++9BY7
kitli6kmu/DjtXr6c0H+rTusRSPNYM1DwjPZwuFZFTdjW021TZCSm+P1zj+yxg/X
jvCIRQmLcdRUvt2KgpELKmsJwXOa9VG/gEF5d4PO+p4swgZemFMRncWYSRYKe2IK
jdFWTlWJRXNSa2eZXLPNNFTbkvOKvSF3sfnm/0/qfTrL/wqK+9r3UaAWdYUK46vB
MqmYviM3G9nYxFr4UsWzHVHQd50UCAsSasar5G0NDjumbMpOWWukECLua1bpwtsf
22YN38xLpzVlCx5T/sc46nuU/bG46wg3m2fWAfQCDzs5FAMEyJAGmTUQNfuJWGPj
GB5AtGbgMriuCFuHcVr1tp2doWMb49BSSg/4tnIh8gFdCPMezp2KSPkNhbWk6rEL
9lgo1vccaL7W28mZpBBVD/2esXnAf4FhMTm0iHIF2cu+WKtEn1UXQ0FV8dbkQNVH
+r9N/rVrXcDTH3K4S4MInBllJCzyKBlpRssgqxX4wmqHqj7HXhACj9ObIwR1mdvg
0zXkg0aQ87nrc5IQfUqQ1dD3ymmFRjT9+A4AQeHp4GpTUFgnIvRH+C63GIcNbw3W
/0d1gc26Z4NarZLXVZT3zjl47erWlFUuREDScjigPPM7Kg1pcj32cGQeDUWOSqP8
fA4WN4YEZZn4+uFgPVLHPS+F334Odv1hWl3FvpvpZELlS/7WcKuck3NrzybZPw3/
LhFuJUcu25DhuorkK+on5aDS9amyKUb+BTmYRMktRCsjR+SI3ve4rFWTE/aY+0Xw
qLaRACTD2zGCH29V3rGu/LIU7CPcxXbtCxnceHLeZjgQEXpFeRlru6/sHSwjz+zm
YrQNw/bkgElIBfnK5SabMaofvGm/wOiZYI5HbHcn9mXrw2bgTW9TJIWwhvZP4XRS
EoTWRjypF9QEH9hqa7W8F9MrBUUgmPf38GUDM7WpHGFeLvcQjj1xrgKQXYWGCJwm
PeLw8oV/GzPUdwbQpgaH8grv2Bw1Z9MOQokCtEDZfBKifoJDQhlGt6jPz22w0Br9
lRsKVe66msTS8rCO+skDgy3+gOTrMEsAefegIcM1drDABDainrKccfaMnonw+UQh
DknUNnzebZRdxp2Vtv+/ubdsRmTGBbjDvQduE+TO6xdCQUz8+Vy67XM9Q2r1G1ly
dc2MiOXAhb1XR7cUqe09lcf0fy/GlQYzOa0MiFU26vVokenazVZeVRSHwjnnuQB/
qav9tGEcO9QSMNo+W0slhfGKcmc78wXwO+HoJUq7kS+qghyTeTMpszkuulaMEone
/FFAQa8+2+S9+11nO0vyxKN3+MobZZ5HMvNNtx2i4+54RW7A3T23Vmfm6yQH2ulo
9FQ6vgNj8ZvrqU8OKLKl/2t/ohg/dmo4jTBiD3kD7Z7egj8wCSBku0MphNiFofgt
8vEvjBfkZ2NFTDdX6en5U4vLLb2kfaBBV/Mbrpaos4nkpkwaQxgOu2/c/+kRaEeU
lPgqNoq36JZBgrwAejzZlH7h3GtSNZyVKtLy1oHDVcL4qf5nD17bv62R1M4CAmPR
osxOIb/togGi85mIU+A+FVdqGZDXwNYPbbEngf0wr4JaJj0dryH6wd/Pvfwpe/1o
4MLFFzZdsCtXCa8MgSMPlEEHlVotXGAh8kCFMitLEusazriQFWzNCobnDD3CFQyH
h3z44ME4D4N9FgTcPCzt3oq4D71LYKHGcyYVLhh58SEXX/RB4TBP3oe27vSUx9g8
smmLiDqWLDvZHEpVHRwnMJwiPd4P14MUJsAFdS8H0VZc0a9LvEOGJ9V8Zi6mYDOo
VyW5ehCaf4ocl8BJRjvOcfi00aKip+abtOBpw8rNxx0K1b8A93vTLdAnerAu0pzB
BbeCP4EpzJ4BTIqBl1v7IBjmCpk+UR/RuTjDi+SBxHW7SHoBs0SbM5WXYJCCfBKq
lPBCuK963TO15imOGXjifrvO9CP8KeKBQ5hK6bzJpIWA24MFCFmU8Sc3cPxE5/FQ
8BTDsWB0tTL1+p+N7aQfzwsJkis4/I6llDjVxLVFBWh8zC7iQZOCC7EcCvFz/k5N
tPDHxoGTfIJ4gkXk75eJyi4Rhjgk8KbiIPcLiUXCU0a42fii5LHeN5D2Eo67j5mN
B4ftpf6nUdI01d64IjOXNaMWgHx+bqPjumzcZXoDgkAlogZLQ6ZAITXNKuBPBWoU
4zoBZd35FIXvGOb4azid5tyqyFOTspofl7gphbhvG4bgMHsgpgB4QZO8Frb6WZgd
2ek2tl6n6tnXYGjz1IbsHruA7cmOiNwrGJqUe6b/zSI+TeElzsVWqVzuYgMTIRvD
r3UYDJyw3NS/ymdCV3oeDJmGML1xxpvvRVF1SFt86QinpGyegtVIA77uJN3GwBYA
23msr5SkN3oFdM/e4ZnMjfUqpMYehh0H5B/Fc0LTi7rFaHmAVmvWfyqV90hPP22b
fb+1nUS09h5L5kp04j6FiDlK7dpMvOvg3nmm19TeBLm9f0Pmv7IzWfS21aq366gG
dMbEWHem2+c4D+WCdiPFsy9adQwoR/NVhdg4PS+isoPEiTf2FhqeRyqMMurEFFBo
nfXmML3RYiXThYr4yjJy64AnkxzJu9aYtjZnLj5Kijq/hXN6F4dyAQZiJL7u0XMR
0U7bv+kko0uXVnj7jkkpVr7fI9Pkip67eQFhSab4ofBW45RbZJGtvg8X4nj++yL8
nx0Dkh9ky1n1hM4iAMZAuAZAueKeJ7PKAGTqPW/0bXLJSC88dfgb5K+ATGEbmQjk
kxuCuFGCs0BXKyGejAyhdW1aWigqrk3bO8jIR8boIwgEcRoU4VpE4eJ0B3rYYJWd
fg6py0o9+e9rAcKe0JOk9qi0Rsf6z7ztNWRn92t+HrHgpJ4zP9lmFi6w8AMmxoPQ
0AV0ZFSR6Yh01ck5VPlotQPeU6zRYYvdpiGOG20WoR0AKYWvCMm9fmYU/XCG3z7C
jcYwkxEpUD1PB5i1d5Lj63FmQ7tPz4DUSdcmwegkZ964xni0KMaTyPeHKuwG/l5k
SEjGoCLYP8sSeWu9KSulEg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
CJkHU8g1nc+Y+jxRVWWGdRN09cOeDCP+58FowrMOm4FV2WDFj957gJzH4PxaIH7r
RGupc9xDWtViHNXbAceCzB33RA/PCRLW131M5LtAU3/vfFKuvrCh1Zo7T/hIS5t6
C3c3Y5CKwIP8FlzBZMDOCOCXowkcNViyddNJyb7+OxGrQ13oY2Xo3MJVLc7EjcPP
LSsjyU3fihClqM7WEDkMEg5H0PD0DpHx4O+I4qY15PWnxfS5Z1Eh/gF1KsHxSnMt
3o2Ke9qrCarJraUWt8P0M3zoVA2Ki6OF1G7RLKWSObEXPLS/PtiNXInK2jTw7Cs7
lXRWkpf/f4WIQ2d/MNxy8Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8720 )
`pragma protect data_block
ZyMW9RMJvpKQXJ7Z9KGX7+S1WqH/AGT3wZXGXGc3DpIofVs3b3B3mqGy7v411gUd
oZitEaHG+QieJ/cwIt997fKxnaFIh2O0h34upZXzkIbxj5BDGir4hbFNPlsutUby
SV1fU0Gx/2X39STlElVotHfJnTTvTEeQoMzQOlkfk9fqVp7mFfZTDGrmXyQ2/Skv
Taavyd9SkjLK3VquIlsJf0N10ZYvxgI8h4Jzlq/QyMM5b9y1wa3TZtuYzB9t0SGP
RDLJTl8G1N2xv0goShbn9EFnpnAPMzweEPEPh42qi8RxEMz4uPPJSTbaKD9Q5sDT
0UcBRDh1v+qJX4rIHzufBq8JRgdt5/CIzmys8xbx7o++499I0mUUNzKXFsRQQUgl
3Ps9XKGksJ5BurWJ34MDJ1V0LqozAjtkP1HfZueJxFvba7Oed8ccN9xPir6W2Slb
tepX6kuvilT1S33LTYS68kcr1BWC69g+IALO7VkWchLIHfwq2w7O97jRWXJNOtJX
9zWrf1Vkj37yL2PvrOpb/59wlZRB7/Gf4/BjqzthSVMNUV3157+E6A+tLVHAwrL2
CK3ekWJUO/Qe2iPB5jXf41HLUQIuGUufmwWTHarXELol0z2dMxXTpvuBtxJfnNlb
9fT8vCoHM43+GxEAHSxj8fWklkFEGAaz63km6XaoVAm0YNwRhU1PAj4belWdUOE1
qERA1QV561LAYJpzE3YmbWS4oZ5+UDD9cyTOLggpZLqvAXBNQAO94++QCGbf2c4G
ms3JwF4UDO4f24wnWToA8iV9vjc7tWgV1Se4uTjWPb47Zn/45A3znVJ45vvMJ/yV
DtOzG+gCZE2KH7SUlo6qy/FCmBf8NACcf9wk1PFcIYEGzWTnzmggqjFzT5oIkBD1
CNKRFGCjWp3/6QpRQUjlsfaEDHNDgG65+WQjIbGbzFCPLD2vJmCeoer6zJA+VE1C
6+bkB5O4mV2Ows4LZtnIjWryJRx/IghWdsWSrMZh9Csrk75RHMZbdw8VVFvzfxbt
3DEPlt4j5pGVfOdUj2r1nLLUpB8VS0L7ZuTParai28C65Vf5tdAb61uyKQWbggFF
queFGhQjqij+yNuR+kQugqQk3ayOXgcQHYmdhZShQkHMAT/JoZGTjyREf0Xa+vSJ
Euj9gPjONeMRYfWMb4q0exFW0iDLa/hCk1vsJ48TegKtYNGf9ExAGilCW2G8xLaQ
RvpaH3ozzsOvAzf5RsqtPU8RXOjZVuZjY2YdHS/HTw3OMvzOFfqCJbm2rZmMQXr5
2md7S6NPdqMXePxDAyf3r+k2rx49iktzv2MCZ4kZEM2OHq3NbeRBTElpiKhL44Ml
41qknj9JdKx792dd5h0pnS5wGgEmtEVB4FAK5Ze8J/S+YdobhhoeGuIZVv3wfd3w
We54FoobrHhabHoWa/1pNz5U9agytlp5YhvQJo1ikstq0hP4H0AfD48G543H0zk1
y5AhHwkcDahUmn2KZHSVDMlHxe2j+SWrvNDOM3JkSP18jVDXsl7wfZAPPj0XycPM
rifB+oQmWbsArgViR2cHrbNlx09fo5ZVeBvzDPTXTQD5QuRJjqyflxEkSXMSt8X6
k+kOIk8V6Ps3un250G2A8i9Qx+ZE0lOd4WBJqfFCR/PdRNj2XlG2MD9V9oaXW0f2
PXveMl4SsOgXkSAS4Cwwxp3tP7reQHxSPqg9Dz1PPZ6NawYiWNZ1pSrW5RtBKwn8
CqBQwF3FE0fIUkg2GXQ3y8zjmWhnrY+xNqd2xhpf6mVG/jeJzrkJshgQOKNM2PnW
Y6jIA8zmxlNa1xApF71dCjDhjdfeW/i3htuaclleG+XpoDh0rE4kaZ8yS7plQOYL
fTLOhlBOm2IWVc0dLFby/kmERD92HFIxgOcFUhLs50YjpzlxWy/olrOMNycaYKe/
DMl2gRJQGZoAXYuv3I4r00HKHWifYOhm1pyo4sjA6KjFCoYu1a88xcld7aOfpM2h
iLzHdHfLCfcDcnOpBzottGtso43YLAceVjVXtWYnrFcLWDJAxJAoMaN5XCSg5NZJ
6pRYqIk0yPxqy4r4AOGToK/ItAqWEQHB2uP0nx/RU9BlygA3Zozs9WyIEtiDeUDF
uy89rK9TYWzg7b4LjEgKWtSy4oLs1iwz/ZQnbOfHrANWM36Hzrcin1VpDRC1o+AC
vd/LACbTAtUyhirRpRumRvo5M8Yv8iuPc6bBHW8+bywyW4iO/Pv+nQCmZ4NGX+J7
tjJJm5HR/h7nhAW8M0B1hiPWbWn55PWvgJ8I7PelbTXX3bRYp3aQXWWNMw+StTiC
T9cIlOGxpVlVenJUfmMpdU25Jcl5dHzxfeWnv7VUmi4avi3/wmh9CBiDdLYTegGg
TaVBSr5iwOollJuxZzNK+0robL64QtnUA4Y1LE1dfqHxPPe8J2BF+FV6QmRG6zFc
fmuuXOYG+UBiIVWs7UKRO+9DaT1ku8V74E2RYjbuA2453bC28BOSgJTvx6USBq0K
WGYoohZzQkk4p/SXzI/1U6iOHZmVwN7qYxfslYA+/UB7OLEsnG9CYy5fXwa0MqG+
UcSAU1K+RMH/0LdnQNEAiEXuBM192wOy/BLePYnizlNWt4+q67Vj723OtMIa11RB
kNKWEqnqWuJurdDAYusjHIgrXZL3MKJgkChOYX5dHiJPIsdF15DQ9jwGVjvvzvnL
RQoqEmrpVv+t8mDJkFY2rkswXH8iVrzPBRiBahfsoigI/zsQC0LGoC8qIs7xkzfC
22C/NmDOZcSjfuhOIaNYwdZecOEB3Mm7Vca3dbJtfzHosckzk3Mbqa01c81Oez1e
rJapOZ50xAtBAd+eYMKmatBIHgXRboaPc/IGluTPNDiQ/W5fjNrJi8DqfkqsBdm5
CBy5RXSrQiaqjFKCWMZlu/q3eumxvm5mEBPjRkWtUQNXUJ8oYPjFhEn/RGvlKZTW
xR+ls8RzkIXXGa2dIsSPMCXU4eEG1t8YC17hL8rZJA78E+9Pj0uSH2j0dVdX+3yt
yzr1lKsFPyXvNr1E9dlyEpRCXD4yq57es5TgepNsaQIRDr+7BZO76xNwlUrN4Z4x
2gv67O4Zd8aMf4lplMyqnJBeB8jdEE5yiUI5iJNiuvdNOwunDr41HRF2ynlvwaD2
N4OQYYoR4L7ic4gquZu3zevQAMshRY2f3ppLvRiOLyULTMPzSIAQmM5HMVBHDJR4
aJymBZ756Is4l12CD/S5vRqxHiyueC78zYe4m6ubpK/hjTogIiVxwYrWMbPZUXIU
JXZ06PFj0+Yw3TbDFr8dMwbXT6u+AIyIjti1A8mqoOOch4GMUtiB11fIivj1P+bv
12OpC8owVdFEGIQdcnKr/ZgunpmBMmjBGpjtx3SgojLVTpYQyACkvK2CWN/OGLzb
hzX0i8tdw0lUS+1VPNeEOvUhd5ZxJEgkumrIqtIB7r1XeUfqd6g01qvfWjT6kJTo
azMkqr1lUyAKX+/F3aFnqi6nZ8OjDk+/ZI0zn1SWU+RNmxf0ac57ZnRNEipdcgSQ
lG7vaOPXCyA9BWxtCxnI64PR4d/Y5fuKUtkTwXF4YMVj0AVgkxN+0DQD1yqz5RzB
LNX1p5XQqntVfqRaj8zITnUm0umJ+v9uVK11QvgT5kzJ1Wr9URl9BibQpm7hoNvH
2M+O9iWc6zt5Q8C+ti2VwugUp+fvvbVS1FHcCiXtPmDF6MQSyHc9e6KigjoWdg/m
PksuwfyinVHPeaMvbx+MfTMH0nT7UdXE/et+7EK+y84JFPJqk4bf2sDwlHR77a4x
5udHT0D7uEVZfyZizU+FiJ8c+6L0H7vmYbLs2iCEmAsXlARFxKkpSHZfyOr7eH4T
tH7tTbzVkO9lXdqqTNwiA2mleBmRNMasbVjQl5zqdAvWc4hVgiugWifQ7Mgtd6Ox
1eVKXHzyLAVXLtVvHzTvoFOZ9W/YJ6mqsJ/btPAhZv+Ftm37Al1eP19Ku7/z7Lti
BaoRztrAgUwsiJyjnWknDffCz1mndQYMTBk0ipixaa9qG8oXJwcR0OlLsYLbLR4r
kDBXXFspijPT6ok1b44dWeUwYVmhvq6b6aOUjAhsUGYdELc2v0eGadBRNaPT38N8
Khm6QPzM8IVw7cOInH0X2MrYPBYO7bVGcLAreBI36JvmxMj1zr5E6hYaUu9FZV/Q
aStnrPibDXLytnyY/0w/Um5ViQmsCnSoxWn72z4EjdLWR8Oy5xLwwEyboAsiwRP7
x5G7rVQ8ddT3V2Q+yLah6+8/Ia6Kgeh2q9Q6E8cU3QPJU3NXFGfprywqDpgPhOQC
VZo2rEU/FVbPGqR8ON9WM4YzGWgvSxFLLL2op32l0BTt/MjXewEbZIO8k487l1LU
nNxJY0A6Its8FO3THtDN4TmhLNLe5P1iClQJ9tf/Qr87Sq3GOElCAuIHxOeYLsFu
JVyfj3SUk+Tmc5ajll7GumZPEb/w1sklzkiPDKHANPTzVJHscUxc5G1j2oyxiBPI
AphsOpfJFFmUltDSQCXL2mEyFSIpKUbZHoX7HBvEGTzannZ19NHhJm62CAO9O5fN
Z2AjfDbs2VUqflRN29bKpy4PReoh88nzw0Zgjyf/NVAgUxTBW71Ir02JGWzNNkwU
Ocg0rH9KqllmIhvG2DgrxhZp7/5UYzPFFh3I+0sNx9k6tTUGzfGAkKAAAu1a24wA
nfY6rGy57kJObVO+AsZxBppZzD5D3CQsPTjR4ZnH/GAguLbgnZ6Lg2cPs1MRz9Pj
GuZ/c7DnIP97pkQCiX6NwbUec47CTKz5NQ7JTfKdvi2oOQFMeM0k6GsH2sQp1iQr
o8drh5++lrXUI2fgk2lyZ9WWeUumWQ+sBX27uThY+ZlkJk88S76zyqufTtGgmAQH
mIeJuip2dCioidDhU1kARjeec2BeV29t0Qs4twLRsy+5InmqS4H/ACHXwY55V00f
cAM0T0m1Ok+napRLwhIaVZt1T/EMN8Eyh2MmMqOOXnF8OGeMT5GT8RjK/v/Rf9co
72znWiD7stYTlfRIY94fqz4RxoG+TkmPp0ZVeod9f7TxD7js1pRvTcODHWZt7AZ6
YsjoMmlBCqwQ07km7JcTdXKov5Vp/9FqtdFZ8CqBzT9TI0brLD+7XgMvaoa0zpFG
jdR1AM1ARVZydSwleH2Lg6ZNSGFtboSaH+lWR+0XJAvHVB+o80ds9/OcXUAp9NRO
9qinuCWvCVTKwzXI0k505QmnH4T1iTyCQcTQvsQTKHfzBDz8alDGgIS0uwxe5rV/
kaSCLW/6K9A5MI+05o3hj5DKcWB7vBNSuQGN+wGbOuKJPLF+lVOe25pfaBeMP8gI
cyH2/yENXcozz8Is+we1CiUqGgclIseNykEDTSu9QEsQDvTDWhtQCbq68Y6aTx5J
EC5/50gyZwQidc+Y3/xB2Z3rzbjcUR1Nn6vQlxsy0sTH3yp8res8mgJDOThSNf3b
mZcDPGzHuyhhzrNQa5HHhE14Kla+K2P3UuHPtaYYMrIYqy/qbgnF2ADFFvLflHsu
t66qAsR41M4i1211fBdqg8km727CzB5D7u4YxxyROFhOQ0ubPDAzYUvMx/vwnq+G
g4qV6WUHulF2eO/kDpnwWeLOZtBOVqn2qr5yPhw5HZgSo8FbVHfwqpPRnXoMTn6q
ryRcqP+XsvjYpL3ai3ZVabe0FBe5gvtAs+2JBNh6tLMp4y9BIiy8l2EENYLQ9HRt
dWK+l9FbF/BlYhZ+UjezF6U9qjaeNGr+YA7be7FEdcKefeTjepd2i4Ru4dsIBhmK
YumzCH4cMGqaO57qulMogrBvC584TCUMAg7XmSoM4JgU+EnOlnVjZOnnzA776H2K
4rnof6QIvaG4SwRIF3pFWKPblMDl1QtfICL7PybydEZcj7PJTNYcc9K1LEbwhqof
oFRVsoqsAB9TOExh8/sEXYsJuXmazrKl3OjuHi/XXpCPCAldlxYevDaYOww3OdiN
+SC7cj/gXd7PoUNBjJpQp7MpPw3CD+tr2ImBVSO9RA08Bzg/3cuETl+SEMl2Rhwy
2VScq6WtUn+vxcLTFD78F1Ex13/8N/xqF88iTGO5O3XVIcLkwmBBZbYzSmN4jNPs
Oqw4CsjHhYtXCXpWC2I/h58RWA7akmvGXkQ1fAjpkEyEvUjctUsTSr/Z9MkCBe+1
QDjJdTMQASeLtnLnrfonKo2h2y5wN3CjslYjNBbwqLGJocc2OnM9dcT4HBfhwjxW
VkLpEvI0TthyBLxQ41sBRqNfito745tLIfl2D25HwwnZqJCJWtbFCS78prV1R+FN
xkpiH5wJaiW2narba/EFNxBl5iHRgfWDv8iHy1+8rFuOn8BUgQvEHBkWoudKmQVk
BMrQxR9Vj+6Yaz9/KQnDE0n1egIHmgdmQCbco/Kt1uL/jNLAlA8LD8LoIFimaLVz
/EIZFR4BdL5baPin8qTfYiz4RC8dbHzGnkVq54VJHvqa+wMtGUwUUZiutJjWaqwD
7qSp8rFYJprtLx/XqcWdBWj9Aswg0pvYkByfiZMG1EiXbSI0Fm6vkPewz2Jtq+Ee
e2NfDPFqLxqPiE/DLR+OZoTBIkiVB98ASfJarPgIPQonYNbZs4mIKv2Y3kczPFXd
XjYFXA2anSNQIktui7Y/5iieI4oA6CqPXpcVHPm8i1X1rlffvyfkdgJU7SaKHhPI
ilP50miYwDD8Z3jaDJB5YN7iHzolf5skIzAX0we8gquqgAPZpvtWriIlNj+o6tI3
qwmQ0XWI/tmpjMw7rWgBiQEpiynAhsRsHitezwvM4wyYXGrotP0Gdvn3I4GfpT91
YDpwUapFtw7U4uqN9TGlcg1Z/hti29vvR1XvLcFXlkcvPPp4x+IPJDRGSGc7ovkl
b+omS8cp5BDBEoDmQTfclQwqqd2HriopTu4zPakY19245QJ1k6vkEU4EhTOaCRYe
r04ZjSavTyipcDpG+Vax5g2UBTCURJzUQ8cdrcOMZmrSOzW31uIEuYUaK9dqLjxX
0j6fI3pFAcPCKTb7VoEU/Gl/KDiyIchMozUV3io2rB3sFtonBbPzMmY3sPeycJjj
JLwowClA7X/OSj7VuWfdZiuGE7fYgMGA5X0jatCzVI/FycOTonzt5RT6m7r/6voc
kPdZ1jEafEJuP4khSeUViEQY/1Vi2PTfapEq4E+X1vXcxHWGF9WHb7oZh+iUi2Dp
sg+SkrpDiFvA+ogiGMioGDdgAdhqGAWZUhdQ6bJ1rlw3izgtZVZQS0peIh6PnmIm
3rsQZVjjQi3P4fgs541N4uhshkKV8+ls6ETX9WTho420oPT1jlb5wh+05oSpsUvF
Ae1X6qYCe2FmrACLxamsOSk49oXtx7C6pLijAvzbuBIvtx3hbT5mZlJjC5Ia+BrN
ODuuxvghmM6p4v1YKl56TYZnneCf73NaJncsXesGff2Uv4bgIZ4OUGE8BSLNgXDo
7OBcGyGbtsGv6pNVvWoxaZ4unAzErenuedC2dzTiJsBfGux58YtuqS/Ta+/mPinw
Fnq8ACQtXooWo5i5Cy15OPKsLUtxUf0G03GGN0cArO/jgJQ9jIxaTFgf81YeVXSz
qZXgMAH+o0nyj57mzqxoCj/NxJ8rNoxmEHGychDMDAbINQVuMx+PPTgjsbQ2ppDv
DcCUxbgkTwLLyUFBJic5i0RLXT9ebv+t8yR2sJGU0vAIj3xG9Ekx7+l7vxha/Jkw
WVB0lcnaFp20O3jIZV3MlIK35IpiEZyJz9PwySwq6X8CnIv2hs5h2LvLdPvVRcxj
3OelqsErAKH0IXwhlIk9WuqINl5UCZJSjpybJgyblwlt61ZWymfreihFwt5IUQbU
n5SykYTsr/X5B8ZAeQx67JMPN0k+1/0SnenncZFhfjXRYSFi9M5jPv3jzr3PSfpP
1mn1p5hw0bA9XcoOyrRT6tHYHSW96LO+wBCQhuZo1r1csd/glVarIbo6kEk7bJ5W
hUYcJw4rtaD68I4SHyy6PhDO1xNt5DiB0qxXIk9vKLjjEwelM2ZBFEXTRvtvCwrS
lTBytpGbC9ZDNuSxZv+zPtlj7IA0uZUgfNy5l18w78qVdosLbILSWJsZ3R2XtJ/i
utEvW3K+2k7B+Q6dtzgUeyT4VkzuAIGLFNBHiKh5ZLbBal837nCaxz5Qiy827/cG
+7Qb/6yccPF82T6vkRTyEid4d565/E+gZE9dVSh64QEReas0XNWIK5iG9464m+EC
sw6G7TDeYdFWtlFcaHBtJWoxyQCZSH9bdabIaIuFSNpSEuEXHgOZvqzfqQbOj44/
esnV0VDWsOxnZaODKOFWCQSG+gsPrcBTeIplHA8BNcDPUm4p+D9D2e02TV+iqIfd
SSaEA4KCCkMY20wCdHkbgSPsWjaYxNU804Fr1+G6s+G9a0+OmAkVCWJnW4ybwEMD
8FmzwcNIwwoMlKmGnDa0JppqlG6cm1xlGhnQmGpbnFU2EvTalYNEFMWT2jFgjxZt
Q9c6yzL6AB++mm9PCmfWfgfK7hcivWTMv/PbcKtHLe8/pRXEwzX9rKIU1uxWhfRO
vsJy3+7COJcmjNoKAUchUM3N4exdnzDDF8mtc0e0iLSfr6MSGS98k7XIrgDQp9bq
dgnyvA+9brBIxX3lxo8nW15BkH2li8sN6g9dOIYpSzhc+4rXPjNXWYrQf8fcGmny
Y2jn95408Dg2HDin2aGUhZnIZUxJ/SdtJYQFEu+qoOnNYAm46yL6M83hjlWE06kw
fBbBSVcwZwVlVqcZVWJtbI+Ay9JOehssk2ui3P9KWrYa/InU1BTAH2WSmKTKhplX
SSMgGAFJ5u5LZ+atkg6qwM/pq1w6pTevCnaP0UQudVvgNFpNTeMBBuk8bxxcEcht
DuYTBoWJeY8Z3+8KCTDB3c9E6pkQxc/Xwbx4t3SwdaSOiF8sxzGojBgeXFygMpu2
3si9YVnCUbUvEtuwWr/4dC9h6gfKRAhRUresQ99VxrUG7MwVRMt8Be8p2xI0xwxR
b1XfsH0BtZed+e8qZush+7nVahOZPCCAZ+iQm74L1mmvB/BjLgNcpaAhgp10VqzS
rCJv/LCqf6FtAbqpg0O+T9jlxVL80sXNAlE3q/mhvQFFEORXcdvk8XbFz/egQHUl
RtBkSzFDjurGXiZ5emSTt5/BafrKn/wv65DS7Z7bMYHnLhGtFtRSwe4RU+XxfXX/
KT29mWTLQGX54OU+ciGA7X8cSNQdj/1KGyqwd/hzFp3hNLGXBQ732xx9+lmlhNiV
KO6QjqoTzwuUP1EQlK3Wk3MEHjwHt9WiT+gtUatdP6GGiEpL/8aSha9hFm5kAli0
YVRnBj7dWhdjmSGvu8tjQ6xTi3VEdQnBb5QjU3AQoxCGRbCfDtNGvcAn4vncIHOZ
4jzvpsNzz+i2Pzx++xm/6VzfU8JijQj0r2tDZ6mGYrcek7jjDP9s/PD/0PGGI0VE
UPlbhCfgy8BRU/JlyqjlBspBFtLuw7Igkmc3oPZtSOPMl4pOWoDg8LVc9iMNPZ7x
M9lBQE42fG6IzT/LJGd5FnidecbODDyqpX9gWDMBb25MeISEt1vHj0E9Gm3luNVz
qMTvEOW7kaMX9d4FvtJQbm6fqKe7oVSZwvEAmD8JUM061b4aIxNpK4xwgoNij1pv
SehF/Qx1XWjeAXCjssVHsVk9O+JyLywkxHwnaThgMSm26lHZACBYDTPrzaDgiPuL
mG7O+Wbkh6iQrylK+wfH5vIrDIP7BYPNOXkGdFRLoPrl9Fa1/4YetuSydgsZjAZh
/u52bC9Q34bcM4tdPUuD75MyKGDkNstLAvWHDSd0n2tPnsdH3CRg+gtTljA8nFZQ
eXuahG+VUi6Fqe+xXrS6E8hrQWVH4b8XmplYaqDsIX2TBZtGKUULFjjPIZE1zRKc
C1w/i3Erap8YfFF69UQ3gmnPvnk3kEMZzncPix1qdegeO1vQPsoohGi00/nBSbfE
irqaRIuBRknFF2KWn86ev8O0+7qhCJVSIaNGBBRR7tBdA9HqQSkTo+qkGQQoVCie
3B2rfhKKqZJvP2PeLnEhtUrQuccOpK9pSUPdR7naXiDvrMJldi71uM3HLvY3Gf7g
l4o/uGtJB+2Jnw2Rj67zMUH9SHcUIn2fMn25gQO4MiQZqI320IIPQ79rST6aIMok
cg3BEecqCKXlW6duamDiEHubKi2PUwzy1wRvQk0YeYeTNqtvbGzFKfa6eBYx0mjK
SNsYWZqJTBSsID5yAaY3QnrgaRj4engqswekCU6v2wtMTJAUWRSioCmkQJ0h2j4t
79rdybPf4Lo+PZGHoo2BM4r0WZ1jkMAXUrpqZqUkqbVvLmsbhhWwpRCTwU3ySIdv
yorQMWRbBCOFZ9+Q1CYmjhorjBAVZy58+9pylU0iTDohBC/2fH7PPXyq12uLmm+u
n3VDkM9b8sjk7sCxW4Akwlw9GZgZfnNq6hsDnBChu2QHPuoZU59k5u8QDLlbw8Rn
JCIxo3wVLAAQwSkrvGaWLVQKjNYKePZ5bd5MT47E1aJJeZtFFCeQ3kY7LMp1An8C
/R0NiD54bxzJsKg2BRrqfW4ESNwe5btbPocnBerN6pLYJkW8w3OyMLS+LqnR3pkr
HicO6TuuhPMLUE2J4NYIVjKV1wZm9qedXD8NyNyOfQv5JVt0DYy1cQczxo3+s08A
MJC/bP4J66dT9woXr4MTNKkK642OgHDsOSl4wPwIa6CLnCAVoc9j8XwhEjzEL+O2
0N/zaPSOUlw6MDERGtQj3BwvakYS4TR+UqbYGXY6BYlp855rM0/KR298CmPVh3P6
XxSNGWS/M0yda87DZA2Wkv+8oz71Zqjg/Cg7uuLBBggjohcbDbzFn5RvsJVF2enC
fKe9Mt3ljC7bu3lIaPiKoc4ge5WpPRCj0YJJryy5bflVH5YnWcUWlOrg1WsEnGjl
tzn7gJNLR9pvVPGpKc9kHS7wqMOFIcjb8tPtLJG61I9ZanFapxH5m8ndJfHs6LiD
GRMZPwPJZzdAMkoMwO4f1sSDb/7apWCJ/8A71OKbiteXzp+aJYyIzJZzbxPDasbY
FYxW6qhZnOnmnAxFZlQS8TxqrJeWdzFQl8JmcycE4wBWV4HdRUA42MDM67UOpZBY
/dHpBOUmQeyPUQCshhtf4hwrvlodUSPXe+lpYK6vL5A2bXB8ONa9Lv8TEIsRJXuU
6bm1Hw1A9y+dux2bOagcIF4vfXATBJCgZJnX3/ABGNku/yEs3M07n9GDVuFJUaKt
dL3J6VG7oCGMQJiallQCKRVW2aIJ4dQyPYpVtwg8xf8UnCJY1JBg+KJblNUKSEmg
vsnWjfAstXffrxIfE3k7d5kfh1kSH9JJOjQMXoC91vLvRjpFyhDRA6WlGNv7jOaP
/zExN3BfFNq8r6Ok3TJNJFCI0Fptlmod4a1pp2N+P2DdfZKc0jWgWt1uDZVSFkqi
mD/CMy9GG5WW4mt4JGuOrq2I3Bd1z6QNwtOLulZOacoXV4U6/aRvhCZwA/IFXhez
ZmbTkaAHO2NlNRLC3gi3vCn5/II6fxDgkM7u1ktHEZmbqruvA4/MAhHjjfZW0bCy
HrXhTz/S/0VMHdSDHHS7vCyttoruAx1FQqOfyJSGAWuCjpTCv8Hm0lSOQaeJvZrT
UDyz70smX1AfNQyvv+ujTqrF6WZCN/yecjoqa2NjYa0=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
D6qaPgx4MhFfEnaAIHZB2VjyoGvvV3ttuMkmSNrld2bLIUNJZnVbMbOypRmqCkZj
2BdQBipq2tbRX6PDJkt75fNRIze9GXvLsRq7D5s2fJ281RQqOEsIMcntp64fLHkc
bxPBYW8/K82dr50kqnDIwxXbYF0ohA9bEnVzf5NCZ7X/EB+O9WeIJmBiJHrOQBWk
u1lSeiQ8Pn4n7HHfX2qdaWKSGVkxaRr0RtMyWbB61Lx56IkrMXvh1t5SK1631tTe
3QlL08s7YqmJ4ZIFgo7YNPNxml8ewPpkyDv5nHdP16OQpk9wyHUDjJgEMoGx+i4i
/asa3hhCufdQ4OXsIu/zqQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4336 )
`pragma protect data_block
7PZcKnHuBDT7egyMnYNdoSknDr5inlHu6JI2K8kgHwTdEXkLOIQHdvNfrCO5KL4V
FFaFRstaxrHTE51OwRCPHNxlZ9la0GJhh+cuB/EkLwZkOPAaUlm9xoQNqwQo4w00
zYrfuNbbAHrogFeFhHnNPvuptPTONPlori38yYvTUHxYyr/IJIxGcxdKiYBbuCaN
Kjzofvyj4ATO7niN3Jh5xCAx/s8RyqaUsGH0zO5DBzrGM3K+viTU9SiW+qgkYXeG
DtN04DNgZ05e9INd/ewIkefS33EA/5MH3lmrx6nQQKCRMRKkCrvt421uHDOPESp6
d/uqh5+QUbng6483V0V9j4oqeX0ZxzrMyQ6ZV3YX3K6XIr3mARL+3MfjA0DHIduR
QvUyHQwoOcqxiSp0+dCg/gcZZQsAeKD4uNzETYnyTkjpIo985JRamlueOPHayvuo
zT+nNMpXdH8Rs2tUNcFWPnAnA+tsXVfymaYUmFLXw33STiWvn7Otw9N7f7bLt+ow
rpmDvQYL4tJKiYEslnLOoXNy5DW68lLF3Fb3QphWkG8bTJ6MtJNGa3IescHlTB0E
JVuyWD8IvQxXkd24OLXqT4GpbO385M4m0vfqMSK6rnQUUYg5SWaMAloJpMzxpzKz
0qMvgvCd9OV1kvVydXC4NBuvfeXeQEm1WzoAevvR3KArBumlqAy0ZVWTexKqlMGE
CMsAZ1uTSyGevzMsFKziMH6V28qhAhU6IskVhHrGWcU+P9r7EhbmGqCqaYNMDVdw
LLDIEkvBlfnXbWUPo21eI7HoGJwNvwqmxsoiKk8dmwcMTGqMRS8GiAOQ2G0wlxWD
iZuuNxOvbS2ITWM8x6qUI0dKh9aQXhHeFqz+OfJW7F3PMiM3YIM3Mkk7LPDv0UEg
vIfSvAOmzupWK3s2SX3f5N2jQ71gnlg8mHY8YQ3ZpoKheLbqiYy6/VtoYPDe12xm
8ysUxcmDFZjE5yV+7/gvR/7d2+UHhuigN2kjCbp8faN7aZafKRKsrBJV0f1kLFhA
z3hQVtbCBOCEnLVhZUEJfMgBoKPbVDIYTJXiELApJ+kZoJRqSrsnRBBReF7j5ZSs
d2EzduaX1SEDifkcmYsSyTFMBOL13T6GjVBHUW4xsn6Ov2XokfPPQiw/RbwpBG7T
gKe7feFcjJVC0RjtnG37YFttmlucgGiX0wwQoJcef6fUmEucFQKZYDNItIo2zq4/
cbRbB3TDbGYiiPxLZSTMab1QGcLnAgFRMae4cxldR7pO+8JCJ8JeqYgAncuM/C8G
AStOR7CZLuzQORTSCwVvDuF2DcooBbxVwlY9HIUz76ItxkQ3+oi00af/79QGHftZ
FfviCb3vPkqzVMGc7jJkvDMNvCh3ny+OEZ2Lrm2QxVVhvIGD3LFJAUc59fJqr9ek
zPJHEt9RwGRWq12LfO3K/o2ePSRGNyboMeNT+BpvYYB7xsR8+e6KAdOWkAOS4/CL
UzS3o3E63igrc2Wvzguvi8Widw3OVrkki4TC6Wvn51C4FFJWUj9l0CRY/VaPK2Ck
8VhWZdQ2MSQzz9aSFnl+uhDqfPtjUeaHSXXS6yAXrEqxluIL6j9wS50Mipk074J+
Df1xvKPuD6fKV4GGxZcOYuXHL0n0kqcwKlqZxjycve1LaO4gBseki43nfrmZ9Xoy
FqULAnlqNS/EpvafwuOb8G9PuDTqRDnQxj6GtMxu0+vSx3QBG20topblv+pKCbm7
QfVNyyMn3lQncTz/sDF5UI2FnNkOsseB0mxDL5S13mF0l2c0+KSSvz8KbO+6O1Oa
6I60nsQiZfQ0jEOQYZlV85h0njGjAJZUtp70j9ve2lA5CBUtfL6zmLFffwg12eOe
P8y/qKzpzIKIqwz2/bNBKxf90qoI2li5eQVtzsmV7Pil/gfwJ5W3WN1SwLaYSlRN
M9idms6B6S1FBlTo2cYkJxhyOWTDxQ7F5xbB5mbdaMXlSFJevg4ZGaplQIcIMKRk
/NPoAn3gLA1mAc1eR8vbnhg20FwQRR2XtSFI2QMwzpF15Ap5SXgQ4ORvPycSIEid
f6fdcDl3SDiVvcn0zCknxZ56dbLqEw7EJWIhriKaP+/QyLQtR+1cUkFBAXWVOQFY
PyVLoSMNeiWecZZQ9i2HKacQkT9/Ya4wq36TIx9Db/XssieQ5zv6ktgKWMiU9MY8
QowFwciODb09uT+sEo417ujpeXpH+cjugfiYfyZR2wkO0bjqdBehI3aKpS1sRtj0
24rIZSCmtS/3XeDcikillQP6nQ5PsV1qFG00Bu5JA09xBkeBk+7N7opWCeWt0lgK
sw0hUxACAs1xlvgB8M+3mU8m78YY2LVHor9qXhXxODXU6qhL8KxXv1d/DLOFnrp0
h947ER2ooEgAzqvVMTmQaphRHPXTqgdNt+yZTCA0jKhz8tLq4f+7rgyHOnSHWoPT
u1Z0scKm4P+1PATwhVUc5n7yOE7qSOy0u14qkgpuxvMY/6/yvEFNiG0muHxXPWT8
Kkw5tcLEzLK+eaN9S+17m+yUxkwy9uBCjVEvbx/v71H7QEcpUY9Zxus9+6AI4Tbt
L3v9ETM+HGaGRyViBiMd2dq63P3NRVQ1x1brh1pW+IgKWDHbMvpiUwuOB9CmRLjZ
o6vS/mY34b3FW97mN8p6MzcvY+A1edw4gIzISzZjkCHwTQkJaYRLXf5cSBm66Hap
BjEtJmmoCFEXhni8cUk4w94irUhccVOxv5uxBNA2lXcqSLoqrWl6PxBWRU5+aVIw
OLXVvVj1CTHEF19fuNKJ6QUENSpFgL2LnI3SvPinDG30MG7UEzAaEDfzcTcC3DJR
wRrWoep56oZfmwuQy/gr3joJrqpPZBwJD4jH2y3qTpG86Zrj26LxpgyuYnIDDbq4
pX7wwndSxYDlGKbGFKck90IfEJKqKqv15pJadZtVKgWbW65icyhD7PUSJI+beXLU
OhYANnAGEzGeBe5xkmb6DwE8CNAg2ESdBsVMrx2TJa08f5sAqOcoYpDYWJTud13C
dY1RfYhM56+UpzvCWnB072WhOSdRi2+sEad1UJogpTsm8tba7SHoA+ncZgOCFIkj
DSIRm58DZZ/SFJJaiARIr8e9J9FxdYit3ndhBuCknEZv9cVurkVeg9vbD7NPDjP4
eKqCG14W9KXejn+Djd9O6ja/F/I08bFvzJ43rz1IrhMqjNmOVaQWVUBs69ebhdsk
ntuRIMGFGqFAY75HqnB+UCpwutTawslRLGOhAS1xHwiaUYJGEG/BGVgXDbX6XBm/
v3AqnCMltq/LBhG+zkGaeXzTZi0NIL44WEtSDHnoPoUKNc9HbGe3pw5UqueoTVWH
x0/N71ngXq+YA7W5ry6GCmqyHPabrtTZKZ6sftmXLLaIfaLSoOKdr+AQqKd0SOJ0
ZrkTFUEFWvC2rUaMJBMWWXLjRompdR9pttp/A+hPkOCyyu6ZER0zBo5M3sXq63k6
CQc0CeTqlYbfyDTihQ35AV3rCnwcPABgwUaSyJDig8H/JJfmObOKByXsmpb04m1g
XDptq5d1jcbGm7e+TYkEk64WJM7XRu74GcXUIHjHk9vP1Hz3T6693Ap1OgYkQkQS
7E55PzcZKy6wavPfYXKeIYRT7Rb0KIe/uujO2xLgB2gZv5dcfuBdmtgOwxCcX4Dp
/w0zjj+Ju+YtdgEu76H4sWbAXw+MPRmKwID6n5GaBxAMhVbJM9EWrrQdcLYunf8z
y22SGTVpA1NnZdF/CISCtIm/IVxDnyS8fO5EwQ3nvtUidCWPNcS+QjXc7vRZvgXx
k5sg/ccxZVgpwFzjqwuh8e00g8jJws3C3iObUr9oixRLrQdJvCQrd3SpGtuztoFU
HMy0aiI9j+czrqcorab2PEtsiU2o/bLFG+KKlIQXPv6EaxVnyOxzBzIsxu9UVOV8
EEXPA7dWnnQrxcGhjdAJL96R6NhjTwLmNzSixRY9elbPQeAYFlf3i9jb7TLNpydJ
vjSEuIhCIRDEv0vGXmM3BXGz6PnP/o+g0JWo1NZ8feJbALGOlVzJ+89EhV7EveS5
w4G0wF5Afto+49czXUhDuh/7PkR6hBsNywuBCc9947OSyfv5ZRiyofiJZzQpcPiN
NLsgufxv3AORWPZMNDfYxI+CGaLqaMcycDhvhStaneotNcKcP822BD6wq6iuANX5
WgcYcD0usQZfGd7PfKTc7WMGwIbHwGbJBYb2NpJO59pNgwwyYwB13qaqziP1p3Ij
cUDRGGf4xgcxUUaVXMIM3uy/tvW+5wBX68QflN8dOHmUAQwcEEmL7MQf6hVrGMYR
gX4vbkyp4Ee00kwXs/QJHHSSiZbkkUC6uzhx2fncvdsUDZmrUzjCnCbnp2qqJMtG
WSz++Xl/z49qEve3CHrPuZXkXHk2iQC2ZQBeEupkrqAh8FqGNy33ddZAtnSUoA5a
C+qunMe5C+owaHzv4ADaguU72YdZnTMhMk5gSlD+mmxMZPH2efMrE8kmu73xd/Yr
7kkvL2B0YIA+VrQuCs6LsEHRLoBDnLy6Z23zCaT5DfOBWYHV7DX2lWd2DRDAHZav
VvArUyg/3q/HKCWTqxZSQoB6tl3JyHombriV+qerckgj8c0QFXiTft+7Hwfykzz+
luFnVLQ8BW+qpfXhvXGuD4Ow4opsEhWWBaCCxFHiY+i99VCyq+0qDrFT42udE931
aaBZDI6bPp86MITu8GkgNFRwTiAeClB0JwWcno8oQGMJWbFAJM3hANl96GJhMDKh
7JyodkRaMzIPBUqtMdeQqQAa1yPnN/sb+Fo9QVxzyBiOwPVRaPQSbtNmrdkOY+Rz
ekRv5CLr/+Kyxi0OnbSTRgP9bq6tGxQAm9cE+1qvQSjOw6JQd/ftqDN7nHzpq4CV
XzJ635y7N9W+qjZ5zQD2KYuQpLqk+P6SqjlHaUE5HqVHAPfVw/Xpfv0cPv5PNkLi
9vgxamImEfmPoyM2KTbg9pe3Wb2DN7ZaiEL2j68F2MNo4Iv2GVZ7SBMmGd1qmpv0
PzisWi8/TVbJIC7cijIY1ioT2ECqjW9Qfkhcu5uKeK1PgfwD0braG6IdT7Kn39yk
PSgPO3Z90XA6q8NZo3uGjB5gjPlLVTow83TPhnq1DNaXWNkit0YETmhXZT8yp3Lz
2Ap/w3AnJVvJHvBY7N4FxYwIGhwlGL+7mJIcfJxxK2HhZuQgOOGPRkOQAEd/sgkm
HBBC6C/Km9SewHAESQOeMwtYv4TtCyZZItkg/e5Xom1S89lawjZFKGq/r0c6SCDC
IAQ4g0Fez6enTBTzpTJasRkBkXJJqpd5P/aawNLaonWuT/68QS0FtDRqJ2Z+eX6R
I6EX8YyVyNo1VQoFeCeIoGeD3beiOPTolSsbPHt4Mfo5qV9wcEgaaNj1nLSMmWVM
D23gqGUaXSkLXjYeI52e1nCaWW7Qo2soZae/MPvg03rm5ErUVzcAkEXmxN9+9Wrr
Ce7ZAyWnSkPJKNvg2+t/wmAXiqO+4CHfMGYotG/4mJBHoMVconPHzep88+apKH7S
5QgJqjBwvtLbjTfNtFaGYdA+hBIN/PT3sQjSUDJdeyLdgMfcHmnbSZG+rV69ndv4
SUzrwJH6MhVDUcvxM51sip1qdykKvHyRUzssFisAFJ51byk1GpdDwTG6oWOJU67E
EyJk+G38yKEH6KEyquav5z37Nih4/QEa6ZhIqM1hXx9n886gRemIXUNzhylheEb1
ouMuUXaJ68kJ04oYkPAouwbt8zBq7sRhZsTG9QhwxgnBv7b43RA/Zs1R9IYudvim
84wCd0stmh0HTW8T6SnAbw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JD8M0ji0RvDrVZDxWw8TXntrEV41y2ERhAe9bNm1PL2yc6q7TRImaZcVQfpDWhvB
Xfg+sESqcScSzQAj5LPcxfW+1wS4nXoEkrRlScPY9TvOKdXIrrOLINIm9i3UJAdY
Zfrft9BuIjOugZHNA+FlhWEu4q9SxuY/SbFXg0mMks262tlP871kfThlF9cEsWbz
zP4RNeUBJNvRcSZh0llcetAfYUEtGAp4u53onH7LbvU2mWrXSredS1L1bb5Tg1Er
Y2H+BBfGdzM8jhlADKdG4QypWqZ4+oY2UxJ2OAZ8F3SZrukijQ+cGk6ikt3NfwjQ
tJXZrXEbQ0v0uK43qf9L5w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6560 )
`pragma protect data_block
1VeMh0VCUvpsHv48fYYxPHhAjA1tk/fQRFu49Pvi0OzmmE5lX/7KY6Jmf2YW4j3V
1SDTkqlaFcGJ/G7WetbIFxl+pzuBbn7WkpVWahI06VAa+IU8eWRn5ow79kFsbnGf
UmsDGg7JHmB/5s7WZxdCTspoA5l2v4cZfxLq4KOPWMW52RyCCp4PTE0sXp+2dseF
9TDThBgY/07rMyiw16tp34K8+vFlDy7jBPTWm7mbOIkXvqViLc85UGE8GakLCDGD
fczNu5EYmUNVzexAB4tWni1Crp4+TA9GJdt5gcrzjfFpn95At4vhl+i0RN4G7IiO
37StmkpJbl2robn9CCfxsT+G/smgq0NnwKaZg46FqG6N43EPZqFmXElaNeBHLnAv
x5fYC7oz/pZq9/CHSCuNgUzPa7dJaqR40aq1mPIXIsgWivSOyO4WNl33Zu3qRm2Z
KUtS6dTstgiy5pXrtT2amwVsj9HXdvpdNR3H5w2BAXAosx3ETUissFqNHFdFiUK3
k+zckTjIUSj0KYJUdwFVtL070X94lrT1pIneQf3kkXytydQvPVGaCtLE35rZ2OjK
YQoQZfveV1DeAuSd6HFLZ8DPHLBj/prWGF9sh/v+xpKWoZJcKegZL1ls+xMXc+Z+
zwB7acdCIISEhGUBve9wW7wM0kL3emIgusEROAZ1jtiHb7LFCX4n24W1gOiApcbo
Y0lIO61cW0g9b+P07Q7A5vUOHqccgzcJIW/O4gZLym2HENneSUjqpT7rAKdhzThm
i/InPN/epvYqJx8ApIItQZBUm7MI67EceN0rdRXR526xxlYxhkOjRZ5qQc2w4gL9
aZ9jXcqJeQXzlhSG4TuyYbXOSoYOJdYJocQxIEsk7GRwU7srPffKn9LFjb3iZ0bl
tYIaw0J3F7ENB0fUZ0zrcqpGtG2Tsj8AMePlDyaLOUx3X0WiCAsmDnmQ7KqNbMpT
CVMDysyQ4Mfxr1F1Xa0tK23PBMQHe5vKVWvlNgy1Cvalufbdw1YTHVSm/m91+uhE
usCA65RJto4nJvPwG26gXMkAchB15NZGYjq6Hzru8BrHOyB8fG8Sbp32urteV0L3
LEmTLNRazY9sYcQ3FMRaqRwrGs4wu11bkF+7hOVMWDLpFbbjBmJI1uXBpjiSl9Pf
QtB4ffBQmQkRU4OIIsRpwauaqZTpz3nCa87n/ITChriOmBz0ZNFc2yg1uUUwx3vi
uFrKLqqUyhO9wOM5FOIrobKe6m3vTvjcqafeiWZrLAk+vcYsqpaVHU1Bj+v2x5bp
KRyKWLoVrjXvlROFdm//LobsbVfkwUHewA1DaAsjB2QChd30KLY+MiRzh9ksGSUH
t7rGAXPY8ABy81vWfZbiUOxc3SkHu/BnT+wHH5PDS7qAR0yw61/Iv2dmiiWkP1wh
NKRVKAb0LS8SKE7Tyaq4tq548u3GU0Gws3RoThAhi/OMmHZpvxcGpnw0hEUd7Ege
k3GqtwhmW12XeRd9Vg8igz7eM/olbcVTn+1hZQJJToFtx/qmRVYoguragG9qI8Wo
WVQlvJlC4uu1YvfstoZmYbETWfMyCRU1UNXuhsMWMcWlm3DtzLjT1sFPzpflpv9u
5A/NAOIDQzIDm0x+mSoyDEimobg4gmseC6o/S5/rlBE6+xHnwOl8W5msO4Pc3mYe
YensJqNIPasfscJvCLLdtQ7D807F18fddcpH97p0fe0OftQ7AfEpDM78+EhaJw79
o+YR4jwgxPfxa3ZIruw4id70frMjRJhscY9YFt8K44v1J5f9Yn/yAlp+ekI5ytan
DjQ1OwM2ef3WA0eoUy8JCkOdn8d+o3mPcnWAUgs2oTg9ZQC6Z2qlkRdmsEfN4YQA
5k8FUDSGZVj4gyhnSJYoXYZ65LIYVJOZpMVOh/d8xVQDGriF+Wd03fYYl7tygXIC
bg0fexvGLQNh6tzR8jtLAxzdTYgz34SXhlCGTOwTwKbMempe6WT2hEOQmEK+GcX5
2b9EsXMLDEX8Pd4JPtHzv5xhsnizhVoSCNX1uCFc4n4+1trhyw9/f9Gs+3f4aMUV
k9Crnkkq4GFMMGnx1Lb6ey1Ng5t/1qPxd6Myp5fDm8Dp6nUO+eUzLQDM+enNr63c
si9+sq7/C+vD50VSXcZ09iRqoLR94jkB9vwtsKlgNnNosUlU2j5KVAvbMTqejAFs
XPjAuf8K9Oij5DNbaVY8KVMHyXCabD4lWMi+SaAAo/fNu20XEEoYHj7jsCT44GvE
P4tXfRVsV1Zi9ben3KRcPfMXe7JoCtudvBdCIyVlxcv43IiDYbMHWx5cc0GkXLQq
2AaE+IlypKorpO6fK3Z/y1CXR6AQGuLemIU8lmZ/J8jZeOjYztoqZhMCy4Ql2HMb
hvV0G7p1MIdcY8XyKLTaxxiXT+2w4PrwVgl9+nSPawCXE/DILGxM38vFy7zHjTTT
OvEUG9H1+Q+UPRbGIvr2VZ5Q1dQ+1jDvmzRfWAYJ3EUUZPdacf0o1+oXGD/H4ZCo
ybe+uDT31m2DtbACAzNa3F5O+ZyvSnpPnv7awNRDXqcyT/MLStxwEHPZwa8d6ej3
JcitXXmXixOz4lX9T6pg+u+h4Y62eur+6WZgL076Ap35Qj3MPPLAPO9+EXqH1tdn
eF5X/C3CAGPSxX2G+5NIYetcFSgYzYsT6ySX3cTPy5KNmgyGEVx68yNF6dBG1ysc
+BHSncyk57oX30tshBBUSoFoH2Wfo3qDtk/MeEzJk1JMkgAknaIu1eAOuPrd0zjS
X7lDYrwNNGBkqkw5TEbqw5en8sg7s2FXyWzzJV6yrUykzqNYC4TBnLYynZmMJ/li
K/f155dUaiGSly+peU0BCEFQ5cNdTUCRjFAN+mo52TgrWAhup9yW4DYD0xL9wn8U
cWI2vVvp/EIzdczobZ9KrTHc0hg4peTHhTRxVH7+lvaimBA4RaUvH1LG4buK1pgo
eNTe0BSfU7QurEp2uZjyYdFRwhEGKl5XOma1iDMVaYuxuEfRFZvU5vq9+hoJywkE
q4vKoyvHTV5P+9StxLnCtGYQjIY7DdUm6mQyJ0FqLenBhE2aLr6Fw6KJZbyknTJs
uMCfOeUjvfaQmZuEyYZjYVbpLpH6pmUlCE/GWreZuPn7fe1Qv8SdUOv70uqVnelX
LPqITklO9FtWjS4CJyZgqA6zkmgdhzqKEBAGr3GBipMzz679A2kSmrnsfUuOoXf2
2DbIgJHaZbohCaCH9qmIKEIZaRcxHOvAv9tEjeXeYNkwvmCAzgrP9Yg85hTGcI9F
4otCQf7Xi9MSvVqcfdGFdAaT1U3VvPQ5GmJZVcD0ga1w/rsTOX66K7VPh4gEHuWj
tlZCojveBnrxOU5GiFAFoq5D5eM1H0hFrZdBEc03m8onvEm1dfaF/Xg0IpSNEIgE
KF34i1QeVL7dgxHt+cwurn+OBYxLzSmOiLV022UYA7A2+e429tjEpSfEQn/GTZFg
ypwOlbMFguUA7eJBIqw1PuxkyEM7Sbo74Q8HizrQ230nnxIJ9cPAjK4XqEnJHtgr
Tf/WcDAR01AzdZqU9Z4L9LtLyWvwSv//zSRoNmDf+4nTa51DMtnZRPa1PGDjgpgd
S23CSnIwokludLXkyxlh9zKSF2EFzuivecqLcrvZtZxrRgjVjqq5RM172J98sXo6
3xXx15O702SYXmqEmoV9RzGAsxEjr2H9FEaLzVIfBg2QunNLio+gu0/RRM4Sxex5
hDo7yWvTfCJRo3YijxfV3XvZrR+ANM10o0eOJYTrJ7u+7kIJNAPoRGsFo23lDYYs
2ylmVWdYp0kQKIUCDHnjErpYhNOj9mbAvMGcVc4C5G9q7a/bH9BLIMg+k6NHhQGc
+Zr3d3blx9ucQ8hl23oZOqknnahbspvHEL55w+zP5TVVh9wOmNraK1j+O2Xoh4Xg
c03+p/t8S+PlMpPJRMNvpI6+gHtOkRe/HapXMlQ2AMxhTgGKcJAXipUI9IEGBZl9
5y9DC03+TFSvBugUTvB/FJUZTwhXknM53+n5vigjwOh3U64Q2mwllx22xHGFybds
s/6gtJxD5KGzx3+53GCjORLTinEjeCHTIyCTZeQZUvibx17MsoRSFMiIvUbPmxLA
s2x+312y7/h1EqgnESTfhJgLNFy32QqkrOlZz6RozveSgpLFBLjX/GY2AXQaKxln
VRd+Nt0vAmGEBYRZ7pkAzqPigUuMjlea7FkVUF2aSO67o5Y1HAIYAvzMvADvTFEv
6Rv4RrHAyn9OCrcrWXjZ3ffxCgYLM/B2X/h4tMEeimli2aEH6a6b3uDsPpWgJz2d
UlrOh/nkxCxSoJQ9DKY9tE70anHuCwDqrIGV4Vxa0ZGXX5z6/tgWWzLlhgfLaBQa
tGenM3X2y+4NEpoYk5myETMNqoYB1oRO8Off+xB8Es4KW/VXkKkG1XkDIiQAdDME
8ELgzlJnSFlsPIBwi2ShiCKZ28z8NQwsOmAPSb3IdJDEzRtcF+cFgm9QeIls0atk
6VZ797Hecmas99mVhz4K95mBMzw2a2+ibYDocjPTiQZ83RFT5MpvJha5qkPhtGc/
K4Nma+CXVluPWrSoZQ25/i486Exd6cNO2S4duxhipcIcYLKpX8lobmqQx2hu4ALr
7LGtPKUeqhlIHnmEBW57mloxZJ10H6lM2j7GhF6THMwytp9aP5n7ssHFUcBheQho
gwxlPJM+O+Rcb2bLmq71hqShjl+Upo9j6um1K9WQnISbHhQxagaeXbfm97tw8n9Y
xMZ843bAjdj4hBDGcSmPtrKdqFumpz47e6+s0O3Og6b1Y7T7vIx/DmMV8EpxT///
juaMVrbzGKWEaq5fVOxWSbyAn5TvgIzkIU9BXrPyK+McmgDh0Cu5ATvtSWJkRgPA
LbB6Lnl9yyqMiSIusOy7ZODhtqwnoeUT9+bZnk1ZlSefZcOR+g2FOxKA9Z7/Yqzx
+qgeK4gBdpROU8QxJVyeIVKZYjSmNv0emgi8S+Y0Fis3eRNDuv/cb1xfoxlGQ5m9
DiBNR/I2igS4zybV0qy1Yd5kXC2uBjV7HH/Ea63lg3eVR1XG1MmAhFIZkBgS/8zK
BuyECVwT5GHPPb5SAug3w23uGhFDOewF8RZKNvG3KvROUi5LmFGVi0vmUc37Rqjs
4e3zYgdHzDwP3hLtV9PYltb5PKWO1bDeO/ddIrDmfIR3qSajHIAl/npUSmdGDH4Z
ZeYgeIqEs4dqEVpp/X1mvo/51EE4PSkFIKKWMPHcLmcuzgiinX9MZaAFXYDTgOxr
74SJyXyD/bfNJ+AoiWWxykNFjPL1mLgDaKTIWff7hLZ5G96BzIlVfayccUEznA7f
mGQVESMvnq1rqQDOL20/YhQnIV706flg6S8I7uEhScLJ63ipgFT6ROTNnOhoVpuv
9dlpxYZvJElQ+JWBalnlBHkWaS8JoGfs8yFc22ho8ikbXF//vCMqjX4xVdK2dtF0
l5B5lVivRu1oZ/alJINR43RN62+c40Bn2iLOXXb4xLu5kDfGvq84HAfZoKsVxjNL
cI72Q/vHa1N3bAqxunK2xgd7ELlELx8wqpM53QaME5YWMqNMEg3XjYErA308NGue
LBOQMhHs6ucItly0yaiRfB8LKm6UhfnFZBXQq9KakDGk7Il2CXM1Rnp5EvQEhxu5
mDJQSbTBbDTGfzJgRXEt9qhNXpD3dSbepMtjCB1VBiMZnagWvsmU+t6F4bpnCPm5
LTJLic83/+7DGh5xeR/26DNZIzoTeDOPDQsQEmURppPW7VKzPD0bRy0d/zxjNENX
drhTARJ7TaBVgLUfR3YTcZgwrZ2B1jTo8YolYKVwDK/gCIxGHsBR+XCWbU75iQOW
PC5bmb6nfxFm0DlRDf1hEw9GcWLomzml8I9wrFsC+gvimkosXFmTVzUK31pF8fFM
buNmVfiAiBj3pEp3I0iyD7btU8L8IAsRndmRHX/gsob4KavQeTt/+js2lYINnqfT
06jaf3MCP8r36dwlzRaPn5lTfd6UmKC1FVyooiuEy+zrD9+Mu6Ljl7Hq2Pq/EpXi
Ejc9fXm73QvJjRRLh0NBFtve8v2B6rzzAShqxza4X0MR/QmYZlNX4e4+IWC/DTEl
ZbwALTjweEdUw+OagXd4BSG/QTbhZBshseEZI0hCn1b7vKqmLSajHNsdDkVx5wBI
7TvnZGmNY/+x9efqg5VuNGi0sQ7GpKSMyBbVjOg+do7oJ0uUe4CP3mHMLMdx5Awv
A9hjmlwoghQNvqc7Sn5eCOK8y/IkCM5rMr8Frh9WmPC0mI1PJRZ6vnjxItNTqc5o
XOvFORGXQLF3aU2m2uf+S4nHGTMkypc92+ADtXIdoTUnNTzufKTLCD739zSv7a/s
PMoR8MaRfu07odf0Hf6TaORGFb+XsY5lXVLgfjdgu7/dfY/mfTK/xK9ryTOOMYE3
eTQ68tYO661CucLgWoFHLt/zp2id7OT8EiizyamdhymT4meAE84Is8wFkRMcoHWY
ly2p3QiU5jifvKXMynG89cuvt4TUMmwcWrv3qQXS3AO35nw0Ba+b3zP4LZpkouQ8
G901Qg4X65VxGhUSoEtXF0brKI+plXh4BfOhbiQueuKKHGXJ4HkHOBfrYV3W03+j
1DdYSfkvP4sOjBJtfBr3c50yM+fsy1gA8R0Yo+uiKwUohQ5YmG+hhaV4oGRVfT39
tMansls2uftUNfe7Un+ILpx08EvR++45BxGARadwyjGOyd0+VvU5/YaR5pwBhjNe
k7cpdNeGYAcHgqdp6J3mofmiYK6mzwN2cdhsZBacg5cIPao02PbUngTKAHSKQSzX
a5SHF0CyEWdgNB06rTEkAw+gvY63RrP6AxlHfsqqSVKHgQ83ZKKIHbRbZqqgE052
QMPevMptm2f2MPlu+gIs1HUV66yVBkT/zv3ja2cqK4nIMMbm+yvER4DhUWLdfBo1
i3Wb/66w1AA2TwKuNcD8jURAyfclVCRC+4lMjyMH03dYe5SaBZB4S8VIV4fZCDF7
qYnQYc2Dyctkmnju8d4Yh2F8kL1+fFX3MzsV/o8L7ujrdPvdPQNE4rKDPNsjbt7m
7EFnXgVx7r6aReZQ9J8K4cpJXkMBFDdPvxkoTbYKii2Ye7oy5NBHEG6+qf+8dDhz
VqpQcXq2P1zlRdfvkGUjXfuUzPLLfd10PObYe0sPEqW6wmMW4zmybHsEYutiHE2T
TT6Q9jeOdQDOzv0n/djPu6BbHWie/zS5Y4UPjvix6cshVo46WcGJe/P9VQbBoA/k
dHz4xJcH1P6ivzb88PYPuKRDanU7uI9puHfn00KbZYav1bsBweLaFbj770kkGzGO
UklTkcGPhBMk9l+6gARlx0kVqzEbjJ63jaqXL7fhrpSvBy96BNlXlF9E9iXZuREl
U9y6WnIS7dIdceBRgHyjCuPvheaA1ACm3AqKJwJVqMyeLnPy6SrmHctsAaOTnbmN
RbUYZM+/9rznXML68Jw730n/nW3VCqANBlK8t+nhRqDek5PAMpYjxuUOIr/+byx5
OrhcYVz+BpcvuMPu5nH9YWIIl55xIF5PmKBt6/+VTC2x28N3ISgbyKauxssCVSt2
UKmbsPG+IlA4zEgEuJTKoVEKyHl9pK3VMJfQkymIqqyxJv1xzm9NjgK5ijFerZac
CJDOFm4sL3qy3qxUNe3vsXrncSZu/uSWGLJfCuxzVCTP/nQHVk2gyOsTzhCig9OS
IhMdA3rbqBiZm/eUzpAFHlUB6MjrerFHn7eX9KdRZaKcTvGAOCrrgCbPbDxqhexb
k5W/IYLOofEYnhNpK4MYsgL0RXsW+AbHl7TN+xTp3FfeqqStOAGRRLwgjMcWzaOF
3hxvcvydNnI0v4EfB2Rb8XK3JFvfDrYEy59HFDZ+6tYpgkC0mObc5gRunt++HVlQ
0cLjTTCoZdBlkuTCv5/ECGN3MypA6+ApS9bEVkC6xEL0xnWicJc+X3ZuQFA88M7A
7Ber91GKEksoBA8QwfAyonejLDw74lXOBmf1ZLeY0lLj78dzCUfnXB+/MGXurYki
VblZiUQDk2WtVQQbyKkK6Ibb+vxlGmHYjfuRfHHsMP91v+QkHrbuoG1N+jo7LpQH
DNENXhjV96hXCREaiTL3UA6EU595ExrG1Ufau4DdD8uCz7zYOVz0jH3q0Px5s3TB
UsaF3jlwIl4bxYU9OqR0tnR29OLcQon6Xm+qXd+Y+m1dyJ0hH0I9E9w3no8iSUie
tQJuarvIZQ7OJxeFeisa+mbENUPv7pJwpj7fCFymla/jX2RXneSIeipnsiihsFfs
vduPRDufuFPxikN77qXvsw0wXPzUex7wzydnvzamQbnQ80TQP7or+WRk66wAmHWb
HLWA9BUIQqslYfpFvZiEOERRRgDVrh9AC/l+0MLyFsZHmd8UAfkHT45mFQ3Kg1TG
NZ2ytn2U1MfR4Hg2tcyJjnqXy+7HB+AD4mX1d3QwEgvsN3NScUgxM+soUepz+iP9
3OY/QPit5fWXoU5Yjb4sVI20zATdhqohGu7mNR7TWfDxO3jN3iZL3yroIwUpWPKO
npWmu2eOwJ55xFBTSZ+017tuMxcbze0kurgeZXPhXmKMShya1s8HxRcVTfsZgUYA
jortsdeK7khV0+p5ZBLTbt357lvv1Eejfq5O8Q2IMvDtFXylahJ7GYzByBNO31Pc
TZjNz4SK24cciAg6uzNYPEpBkcHNvshlCYCpZzQ7vYwxHuR8NzKx2qVoWtv60ZMW
DhGKM8Ex0URYJJxw/2GxfcNHZlpngSZ3ttIHmbMLRGg=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
S8Gu5+SJFCNQS+KOk1pqWl1GiYOktAf28REiSfIKZNT79JiPtDmR9p5Jd1OPqCJm
6eoY7NbFczhmzGL53ImOhAv24rQk2fWdKRp5HYLfjA7n/P3BQtW3L4bMFTktg8sh
JcnaPNAMM+t2E+O5Zxzj2pPoxZmT3UAwAAQ+9aCE3FS1o5XYeYF88vOfga+O0Peu
lidJfKzLwJY4acIKB8NMw+j3nS90xHeljZooE8cAWJ90YAjelYbLDErnSAl3ZtH2
n0V6nOi4dAC7v94pu45cCS5q7wK/W4xbiEMjZRZh7yyyWsCahKavBHTMez+9WKtk
TPWqvnOLZ/PO8o1pQScFBg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8928 )
`pragma protect data_block
cNZPjgKU4V8gftS3iQotttl6bn1WSKThBRFm6/RWJ3UUHZPVAOD2m2kwaK+zPcRw
rLYBbgVdGwbH0qZ3lsi++1Hf+Ys9nNM51E1isiyBO6Qp0mlDTDyQP4KYBU0kjEgs
UoXVLxXcTJsGc4nopHAd29N55tobWMsY6y2FRw7rlbUMvk34GLw6perEbFG4EhrP
+F1/r+TKnFyYbv1aAEWnTCs9uRWb7fE8rcHLsRuifi6Z//tJD9pwtjsDo35S1VGO
Rg2stkdhqgD/Bv7ad4/NtvP6V0kPeVu3b+Ci6TPg/+jlDCelKMFVk2MOz8EThB4K
rU1eR9YqHAXSL1cILIsEZHA10McapZSKGNpf1nSYXIICHQp85rMFEkRyulrBq8un
O3s/Qluxt35XLmqjH4trY5L3hWoVxahOPaVWCc1ua7m0VI4KQSENmXei865gfRDe
9KICXNHC649brwK/8JnQHbMwWrPnGJv7q7aWwMzokHU6wPJFPEyrEN6hHv2CpQCk
ofbBihqfYKa7W48WNa7X8TM1VeLSsALGHzM4G6kgU4GRaTWScRtp1BBB51MTqi3k
lIaJACyfggaqHABCG6y6SdVl68rS6kqRe4TUHQfAoxZ/XiyzfXxq8khQjl8OneEZ
Gn7dryhqgigXWs/FDPBp4iQiejxuJB6VUOON7Pho5FPPXb/zVkkWQclaM1+qupR2
cWkex0JM5AqgxmQp9Ifi5UzlCTs5fya/eZTRZtFbvUJp/2iSDMbC0U7rTSz08NS7
+JPjQCUpdBBFrDXV3c1tinYPW8onskna+wH7qyMCIzqHj7uve/EbdtlREDKCu9Le
SRJ9R1zc2Ik6cugUw3QAwJSgmxUB9E3koEgDyM54omCWOTo5rdc1n9zxS8sC0QiX
2ugIclPk1KFDWJMfXaDzme6fktSr0MCCVkpEFLbCkiAckDkPG7GB2k608Edug6Hk
nf8tApmPKK9b35UbX2wX2Lt6VsKfBrahmxOwJvdcVUFz7zkFJh9k1ob/yW5a2tb3
4SpcnhYcYlI0khDS+JLcZbwtoSqZ9SOgk3JIJhe3gHV9cR4bkQK/uoP/brZSqQLY
Tphlv0PlQGFhEEInPZDnues4boQ59WG++gA6AhvWu2uOOV7mARgAuOW9CgQRzt6s
xTdxfoArviaM2QbRl3c2kgWBapBFKi/vWw0VOsOS8E7SJ8OqRUTegFaejIWnG+Xs
CVa8htYJ+//zPCqzgXKlHnWJ2OY89PiqIOK533xGe3qpLxPuQiWqUYc5wxk6BSef
VF7hlgj6Wv+esc90TXc4HNHww5fktnXR0kZaVl6i6ljtmUewXdRqxkR+JEiFab8d
Td5fQIR0yyj/mdeLu3S+MrmPQEjY4FhFk3JP0NEyG656vNAyeCSPc4sIwZkk+UZI
l6biBDqwHQx26gSREhhW0D3sbZN4IRJWNIhouXC5O2qS0xxsv0i9lnYXaI/dCNfp
tq1hPEOCd6TUevxmoEMfPL0yUs1Sl3BC+joChnJTx4opOUOoRQ7blTItRYXBjtB3
xvU0cJZVxndBmwHXP65ziFly7u7I2sG0/oxIOi6KudWT9+xV8e3xJw4SIVg2Jfaj
wWGOPPw60xofZumithGWLmQzVxx9XK850FkDWCyYq1KB0Iz45AU6II+vagC0T4un
KhZXfJzmzr0gNbH/0be6RYKG/qyj3UXfrnQYXevlTL3tpz4Z+n1eOk4D0IDYFoCG
3LcbgK8rifgGzaAvc+sgHL6caejFDXmGEcIYrVjkX3l2UE7PdaQLhYbLA6yIYCqI
+qw8XGXIa9VAE+UXIHXzPPZqNfCAwrUOEiSGjcB32WMsuzMR6UZ2LoQJoMXgRHg0
cVvSnlXFcjMVMqLnQWLQ3QHPZlzn1UZKaIQBDqkSHVLrCkoxbp/TAiwVQMQH65xA
iL6mq+op399kjqGQIqV5rHOuRMpCxrm/hQH/lq6OWEPVRgCOZtK/lK1gDDXUIho9
qNLcyZMFqncJJzQG5mgr9mBzOXqNPtqu4t8boJjuh+tE28o71hyVrMd5XZOM6QuR
BqBpd1gUG53o0r+1vd4Uw9Bxsq0VHTQpWI51hrJx5NCf8lss2WIStyRp152kaG5D
qmf9Aq1bMCGZaqbwzJmDLJcqUudDTmPrj6eS6oEyJtrndyzNFZhoh7GZsaXZeGr7
QrWcWsOQ1dNT3HkgI8m3qrMq6ZAWyu9eHa3AwnIjEmd+SbWqYGsM2X2MdBwST4VY
HL+op/ayfVAv+NUj7cf4nTwznVUGQigdgSPcfFFEMdjACi10hgzNkR72j6/tigMQ
/0IzTYz1JW+aETQN1D/H2o1XimFMiqYrMtkhV6H0uRdVDxY6z6dtL2Yt4Jg8Jepx
WlZ26A1irq6m7Vl8JH4O3gHfEqBXkWEi2pxdfo7GEwblYLlFdndtosLRZDwLNDjD
wghSvKeBhGQLAIqbiB92ZrN+guNqOPPpJuq47AqIdpCzcXddP+n5YpjDU0ztP3YX
yIM2erUNd/sVwU7bYCiYzesb8QgtxZ1Jlj5tvBXBXCiso3RFRK4U1ki/jpUn6vrV
sQY6jrp/cO5JxDRl0/OvdwMAmPe+bcHBTnt1P7e08QWAKUdRJurvMeyJhly97N2q
Ss4tzDWImxkQORd9PcimWnb0adRA6KY96Cc6lFrLigOxpxixs+YyKt2trzORtB30
1q463LOTF0fTc9LsHB9rrA2l5hQo3ueBNrqkGdj39u99X0d70xOx43hxwcpW5Mx9
MOKlaEiQwUYL0RAXaq2whSFO04saqtx1AgvRMcOcYoLgiFbFMCQt6i4VautXUZ77
SuMm5qiyjRP2Q5HlAxSdfVKJJZPv74RHmvVCjry6srmFcJZQCxgnH3hXyTZSw4od
Bv+cIFlcWkA4Oi0+RAwkPZpjetCoffJswEsrAY+9Fcjr9zzIEFUMMOA1JKsgQ0gs
d04708hjnOfNdQhHIOKGs8D3yt5kdXmp/KyAuroWSrBoX8izNQwjneTUhquNWnLD
q4+zGnY2/Woq8M0L/SyxqwM8uehTLADTxUXSD1VUSYQ6a6TGgN+vy0ST4Ly0Nggw
p2/7DZ2mS5pSRXepUp6fM69Vb2/CF7Vk1HcP+c0JFQSeKYTjOxauUbwxmji3pCqU
vHH7V0Ys68JjdICtqbKQ81EWe+g106lycAJtWU+n7QNE6PVstQSxXaae3hBDQz3t
lmnXX4U6iLT2Yck9MD3ofJ1vuP/F7FSpcU9mPiodBE4rlK+Lp0IV0u5XFlIR+LlW
O0gwIQSl+gxHZIL2zSjK6mnyvcqRfZ9f9RmfeGa+XK3dUR5OTNyfMXsruOtrPXVL
dleCnjnrbsTQqx5t9HOAJ70rR3c0oK1rb2AJHCh76Hxc5OY+RCwBNQb5vNkSef7i
3GTlU9lrjV1mcU/qwNE7bgv5bm0BvKPCJ9B/JDPV/SPur4jf+A25IvXU5D2q792h
AzGx5IpAXGDAssApn3JC9Cro6PdtfyLMliPpVlDWOo0W3tWdo5e8wUMWOGqsf4LX
OGwhbB19xFmPESgaZGgstTFYINHrQSjPmLXu8JyVqG4Zduom2RT3hzjvuKJpgKJX
0/m4JbHb0BnTy8iytgWYqcKgoRWhD37JlruRw6vKzlhQYQZaVqCaaHIwjzCf64D0
xbekBC1RH4TCQqNKlW1QxUQGWSU4lF2zCljx8bHRcv2fr8R4Y15VXrkBNlyCP9qv
6vmd197a+oJJq4wCwDANvhmWC9ZtgWeNewANz7Kdoz0OrDQrQNVqMT07SADin9sR
l23V/Ss+7R9hzDZ+/JLMkpNgznmP9arZMObdzO9Q4hv+M/FdA2vNZO2WqALf6Cbo
GIP8YKV9jBh+KCbSYKHShbxA156TMe/p7trFxk9Cf+G6vgr+ZF/KD3IgSXMVI2jV
pfy78G77fA3iT2d5YADcEyPCL2r/djY0QMzoBgKWt6psD0p9oxDjxKtQDRhjacUq
f7y3KTyacj0ZPncU+aNrkq9JMXmb+ZN3IAy1XYvw7BYtY074Mx0nWG4j9qrIsXF5
Tc1DNtwk6OeHxcaOB3aeKUIwanDX0dBz0xOegpjEWKaJ6u2eYtqOHJBC9G/tGAtB
+tPFVjZo0RgsxePurld1pxA/Heilcw/PqtWNd0VSork1TzKUsczqkPiDouC3M3fn
Clz07wcr1eBYrt76M3WEXNQsbV8H4KtvVNYaDAhkQEve2V/jt6GRdSvwsPZMqgUs
VrjbmcLHJwRjkMocYY2eUyiNa2hz+aV7yoGmF/6wGAbT8nYt87sTFBQ2dyjamKz/
k3rR0DmHsb9kgol0MxxUEZy+tu7ivRV/mX/neAUwKX3ziRO0tsbGz0pJXmzwDhQt
iBuK5ri8FfKOy7ARQr1RFXjLCXf8QqgIjbfcqagSRdGGv5/FUk0y41QwhBd7YSfh
g/zY3ydWhe9wMAKqu8S78vtYUuEsKdIOtJk4aN54MsPldJJUuz4md/wAcYYmMRrr
yzhU2ep28FF9hVTkZyMJqWboweYf+Uy8r0zNfJEYNKHlOGHbHqI5lMUsrivMbFcv
romq8dTEcOK5yNdMOul8FSe44PgpBfd0ss1JAdWLtKdSSw/GRttgQKdnS3uxmnZr
e62ktdVbIqcEMGOZ6CulIARFXJQse0I+fy6n6iFz6Wiwk0A7OVe/u0JaLpYHYGlQ
B45Gu6xvTu2M0O1jlgOukQvMhyxQHqO5ZPwGq1NZwZT0P/+hw+kzBx0010tfE+Db
JJXRLCsot1njWZTci16u4d1sEN1KfgY2dGnAvQdIx1xsSH4IFa0HllMYJ4kVVrTC
h8VhPouOyhh1Us4vot9ImXEMeOSVF/kNMwieOphuBbbQO6epP3b/Jz3sGAQsmPx1
v/odNiQOMX2eEZmQxFhi3d5cKxPvEnAguMSBOlCiuo63NMe9kUWQBAwZqg9KqFTy
a5jYXcasnxX4Y2ahzUizvfgD/UelfLb1ms1j8hKgTaWTAmvQsucx3r/Hb3TK5dJ2
ZAjyGfj2ykInnejb7k3Kja54THzQA3hRDFVawXf9d7d2OJgXoclGufutyC+N4gky
SIuJCguYUpgkI7CHi+8mKVugy/pAmXQF1E1AsuLdaV+Z0EJH8Fef98HWNkQ19fNT
LWBXGDqkbRqJcJJ1HDwkTnGpCgbcFIgAgr7wezZ48+aLcrM/auL4aU3+iMXqZoLB
GMfkx/zQqRIb0NaOUsdu94MCymB9HeD2Ah6hwOGjmtQeBgB53c+NnSOH7XhHgdT4
w2f/sNg8RkjksodPIpJQVlTlKG2W5wTMahNsH0lnC49pXXTI6J2nuCrkW/YM4Ffy
RW2rnBq3BF2qk7rbtiACSfgaUCuW31yfAx6Riiga3YHql3iZF0xXHcd7Fk58t0a/
ecr4mRDcDZ6tbDLXyDyOdzMBnFqhX9GbMS9tjkVrLuUcRilI9kSPltzPDbGNqKXV
/FyKdCWjuHV9aMAVMk0FDbpWqkuRRH7ZVAzBk0Uz2iNOAVTSd7/BFCQoRaIA5+JH
bsECEKdL2lrm077DP/qAKQwDZKIqoaSukI+L2/mOKuUvWNJrR7DaEEaIZ9J9yXc/
Qeo//09zmkjemxSf6t360oWd4K2ged2crbRoCwIVeMoWOxoAd1kJ2l01tgG6WxBK
tc2XEe46HNiWbfVOg2IdPOl75iGDp6Yfbxxhxgz8TnRvkJlxvsWPMotoMogL9FKq
Xj72pHJOWdSHZcvMRRUU62JdzOMX1qy+Fq9sGj2Vz7q+RGBvqiwpnVrZpwc/Md+F
Ojtui63sZB/VSqDuhQd+R/OMvY/ye3KcGzA01hMR6PAWznCVLgbmEYUG+/RUKYqG
ACMULD+40hVUcP0Wf3YRHnLV5ae3FWDNOTi5vrcpDiDkHBLk4t5jBVKbDGHRXSiA
j5OdE9PSvDSzR44a5MNBuf3mkbMMQktgnngMQdKi6Ff0FEyf5qrHaV3snCpBBR6A
nXWi752iYBeEjvvmhNTBxFBDj+fuQMmrHXwwQSFQsInnLYXCk1vnOz44iQoPrePa
BhTB8jFYkepf4+F1ZB02k2xnoT1b8x4KAMWKP79EcCNNZC43iy/pOpyEiVJk/ytS
SStdJ7LcIvvbLCNmdLbHMkC+1bVLvaI16Sh4Ngy17r4MZ50p5ek9QKskSC5wkaF4
W4GykwAEJlqqlD8LGR6GZqXHqk1GduiwPR9xNzUVPnL5Gr334NXMZhU2EVVScdT1
/nLFKxIBKQliX7KFm6DOCNZ39Fy2KMgN99wAEAOXLRY3bMA6t1LNcNKf/+vbjlWU
JN6eibiId8/qcj/W1/Am4sIp/WAKgqSWYFgVMtsFyxFLyyTwmApwsJwKJCtICrcF
o1ZnszM550/w8l0LdL6B7Tb5jm/koZm61+unV1ZUU7dTW7GEpHfiZeSHo3xvj0VI
SLbUsk5w2LpEWYX2qlogok5o49qbXyPnII3IQn1avj8V6hJ0oLzTJAB6gFwH5Dq5
lBZlYYxbxiUxWXWf+LN9oIqX3hNMt7fYDhr1XeDVFO79ARTbXKCUHNRT1/r+VFZq
O9frYGLGlfP0snE0mPeYxTnH+uV2hNXQIrsTFgD5m/ultju+9v/eYxyIWocUQAdQ
iIj5aLhjv9JJ0sjgD5YfYi8BP3z52hy7bjAfaY68R3e/4QVvG0+j2aFktDqD8lhy
DpO1AesLS1IReDHxYBnyOyHySpOTKWFclF5DFFpg+QcLZaF7a6APg/fj18uM2u1V
H86Ah8BU6rQ+HdUdOEpiSPN8LhML3n+4KhjdFSyT82QVAV1FclHIl9e9yfKtKxUU
orqMjQ0aNU7njlRNGxjX9DI36bLzE+yzlW+xQmsrvbUn7mT5y7mws+cM1XCeTrRr
0XttPJXhMe6rWEt3B7SyfEMYiASvpgIIz+18p5GqKBtVSf5LPEOztkOzCPRRw6Em
rnOV6VkvtKm8oZBdLC2FGkifBO8QgTnxAz+PM2tg3g38k/6y4P3++NW+8cQpJMt9
UocfJZVx2vVy8640pA9YGvCqfI+c64UEhFd0ZvzhTWrMkzQ+tC16U85s+6fGyLVM
0mjz1VDLYQ8y0WEI8AvIQkKHd3x8JuIKS9rmc3heellidSzcOTnMgPx54Ja63yEd
Q9Rn5qVDPhqTwaeAKqhQc7WvPzf2qP8QkNiZ9F6ezqQ7Xmu8jY+UXUtAUPNab7qn
1l7RyblX11lZR78VJ7eFgFV7DKlFGlGI3zDc1m5+PUJ61XFtSJvaNhXfRDGbYDM7
nqJ11Im5VjYohrpyQ6VVMyJaVAxezl80M42TAVt6jEP3hqB4VqiHGVYeW7ehoadu
MD+12yLARA7i9HB5hzfmcdVFOGGlQBLrMnKvnaf5FstXXj/5xCufZvvYvAq+GMWR
3aV2SUP+38xYsiZ62EnW/WLD4BkRVWq/g/SqkrRnAJsD/1FB1WAWzJpcSjYuc5zh
BdK/lhLhKDKVGetwJgf5IQ7EK9604yNgxQUiF4u+/G1c/4DcqeqewI8KUfO4/HfG
D1G3rzIWxIuQwdi5mPPTZhHAtkGUb24f/N/4jo5Fa9lTU2XZlieGW9XsYaa/El92
xihRIZMDBOmRUA9M+NKTEo+DHKuol/JbuzgK3f8xrWipbdmRgybHwiHIJiJnYI+0
4zGRv3JWzgjgnATwdxBrfy2G7OAr+6JyFECg2c5pSQfWwHtjQ3ThfyHhsw9HQguC
OC1YgavBmzcFwvKvvFkwvW7B67Lj4ADNO2Sd29MKBVH4W0SYUauIaWx5VbT3dgyq
5MN0akRxsOY4wtOeyn8PwgFnyIY5orxmF7axH+23/MrTib780vCVoasDBRJYXTA4
0QVKcIxeBGDytmIH4AAhdfm68O7y21RQF+yEYIEMQaDAwpf/xV4Eb4oAsipvX94R
BYqApWfx5NUDSfLOYNQNh33/162JOat4g3AMk6L8IEqhrbBcVXnTFbU19OsvCFiB
D+DPuXAgvkYJpFMQMyt3yajfXFPbIBffVFIV7giCYE/34331JPOQGCS5bLunkVxz
l2WlBbHrsR9qWupSKsTknzV75u1gREyEPW01JA7cwJ91sxOWyoW2MRiGZyu6WI3O
XjOdzRARONaMuBctH/fabvXg4I9Cp7nKmAbqVZNKn3T6oODGeAGxMM/BN/Db60oL
g3TpelnCR9zIpZ53AJ2K6OVI4XWBe1Vc18zfy9xFEm+/lFUFrDJ0Algp+jUvmlUQ
am2b9jR3/E1hpsPm2Hf8xPkBeexTeuM9lbt15BopUmOl67xFikxm1GlJpha94J77
TBlewBGBhKq/n9DNBCwbaiO3UdkTkuwbeUXELE4/MHhZ8ECqev0dRhNY4vizXVAf
MD7utE5sxaDTmHqCz3vbd2W/shDb/3whUwLEI+IPOn2lr3METHOvA3dMoSbO9rA2
I8SZm127bz8O03h3xHjgAsETl+Jl7KoMM+Yc0c2TChi7T+IvufiVsCqOvedZTHv9
iy1uCrlaE3eg94GCt/Q2O7YfqOB/fg5BvWmGn5ofvfdkka15ShqJ7hovugudtAuY
0temQhfWrzraL7vO31mAtHVwynMaROAHc0l1Qnae8IhSxLX6dY0AUOw/YKDIUjdZ
I1dkiC05ZGTAvkQ+t7hOOvpIEkgGdnrhdyWZvJCWPTl917hygSE6BoBG8TztOUhk
ZpvSPwGpODwhdkrISgQFSMoV7SFZuXOgPlUDHYV2IqAIg3bg1eke/7murwV6HZTj
bjOs+iLL4I2nUkoUC71m36fSx7y0Ac5ohK8+iaXP/AhAaSijs+5eZPNTZbWArvjX
5mSMOCCqjoxEVdbsNdiOFssmv1WNZKOk5lojks5lKMdjW74Pp3V7b4nuTeToKH8h
TFsRaBAowdZ42F8b4p5lWlaukoyqqDYFo1UfnZLZKzOtg06HtkoCZR16FLNZP5+D
+ziZEZ0wUaHQw9QnnsfbqX2IpIUu1wiq9jxPH9FdyupN3rreWqZcMhRxEYbAht7X
8X1tFwVYwQ5o4puNypbAVV5XXxJGLln3rzkYTWXN+G17PDsyMLTYzF/1cGuQiUcc
6QKIA2LMNn0NoaDYD4M5TP8t0YTHkHxX2islppPjPrc2zIhMcaMDoojn+ArbGbNu
jrkwDz2gEug9vZsysbKaRIvBhepJahw/4x7VCdUJoim9xeAkqE3SPKaNiDzkkUg+
hSXzjHN4Y3Ww5LT/JSQxiWKc5F9AhjClkWp/RIScs/hpd1pz90boYhitexsqsJQJ
5A6CSSk8RGeMHOvh4LgMiRgEGiBT1AO7x1g2zcCCTNG/Bb+h3q6IW3GF48uGYysz
1mXClgF5Ms5VpQmoPpGNkF46fA5ykDCR1zqJKuE3k7uVqzDnYR6s+n4U4YmEzUfE
OptjbzWB+e/SFXgfF/qnI2MhBloce0M8G43ED1i8cdN1PlWJ+9P2Hr30+bl+rXHJ
hrEBpJ5veob6efeXlXVnOsHU5Mp+oA/sggqvt11zgUgPPQ0borteOCBkSJRjQmfU
fG5dsbWsRlbDNwF7HGTBwLCGwYuTN8/99zGn0zEKwzJuQa/YsUK/UNTQDuCybd0V
/MLArdWp7as2pxTlaKHYngC3z1FVjB0CSGjKZKmOXTKuZERSzwtCq6P1inJQK/og
RdOfGrJ3oUCXCxPS+f4Ysbme0099XZoxIpVg+w7ctvMYrZDFn5RjTLgwu22vUhwf
xnGT/pgGPaZ9BV6KjBmOen0+SqBdtcDPLk4qoqzHTXlXSgRmjPGA5wcIF6VCSXkK
6XZ6x25L8qj6Fp7ro0BRuDoMD+W6b8vFruQaARCS6bAch0DzzCTjxPAahfszPaxH
2OyBZYKK32ME9SsnA6M8wJ4iu4Q0PUyvmGriqSARA+ZZKOH+GPuThl04r5rBmVs6
dqb1rlAWzHUv8l1VuxLiSnMfzTH2LKQXZ82HSQzIBel+RJpTWOzWwuQRd++xTmKV
e5j9vKZtgBO2TmrwEeoRcvgbGSLUcV70DXWg31y2N3P7yfZlyIuEweZCfTYGcLM3
xrXgVK6nRyLfqY74bge8S1sh7k8XZq3OGEN6PGkJUruSzxDWV7EC0N19zWrOrgGq
Y2a9gLClun3pb4wx3a+F/dwoTh9sVLqqPU1mdECc+ey9w9Ne0iHiFZI5AZz2iFfj
4QavLDqj12m+2eksD6CUvxtTESwSiWcr4RlDm5usYjQGJq6Y5jsXXCfJS1pzDN3m
xSjJxXuxMn7HytQ2NVd++IfGX5WEM+kXO5c0z8Bdxh1yTc1iDX8IX6zaU1vE+Kjz
Re+2qjjv4gCKgz8vmOR7nUxowlQ5PLjgBkZD4l2oG1xnGv2pIxuvGErtmtRYLKEL
rkNzkvyvngAnNKn2h7P9U9n3JmvEQF+RKRaef5as8Q2w7SQOXILdFjCEpac8T09t
EQR0xtkwi7sAh0o9f1anZeUN5boTZR0PS44hWpZY9qZ7JZ+d2Crg3xv+dQwW63GL
aIsiNW/qURaUW75TIOgmMJAVaeWWUNNwxi35NFCQ9plVjF0r6wVcH/etUc3wghxI
3QqEEybs6Mc3LrBCbyRh8h2sL+wwQ/JZzJ/mt2eMoxLara6fv0KiADGGmyZNzcEK
+a+JD3IOcHpjlcC15GESVz5Taqiz8AkFD0ksTEIOJaQz6ESlLqMk5tu5K23yYGTm
Wrh0wLNGSQsYljSObI6A8+AHlbdwr64LUonGOGp9D0dCY1fh6lJYcik7ewKV4j+J
lLFJnScAMZz/Gn2+n5TIOG0BDgDM9qJ90YwGgvTSuf810KnOoYdcQgahDW9RWd6k
ul9j9jW67HoV3zxqesDrhmAhRlBlBTI/KcNu0UTFe54iSpx31Ew9m8w5CPhl9vF7
9utNjmXDgfpaTDDtms9TWZuyYTRVhNGFGNmdlqUjJ1xutwSTi2lZfoOS9nB6NURX
07FFRuMrnZE8SqdhSTEdTuAqqQFCGJGIf6H7xM+S0gWEYBnzlHVgHRPSmTz9dauO
hJysbDm7EwllhY7nXoL8Nk+dZEpRP18jZZPKfWDFKjVvVQFF2j4jKv4px0wpLDfE
7uzYXRUalU1kVOTaonchyPMJReiad1AWoYxRYK4w9Y4syOGsXu2OwtKQYrxmGHKk
Rl0JpPzTqt08q7uAw9O9YwIJaH6jR5CcacbBkGDkdxiR+SIEOJbk2reFsZTcDOZL
n13Wnv8qXjtwuJfSTj/KR3n+yYnBInaGsrBMILhbUoZyRBC9bMBH/1FDZrpoH8gB
Urfk5xRhUSQbU4Thav9tooUdY1nS1ZdXUaUba4YCOTjbyRa5jw3IgJw22CILHYZ5
7jShWEt9zG/nEyVea8TVgmzqw7wf61kVV3ZJRQKALvjrIuWr5j+BG3nOGHjd5Tlo
7pDns/sypAwGpxGLgOIXH6YiXa0RJSor7x+XRrOM1kxb34zdEaLl0+Jjl/UfbjZB
PLwcU/Uj+Ah3HqCLko0uD3KtkILOZ2ImRssGt8HzgWl+aRPrWEYuFPXBgrDQdwEr
BOhJYsiyTQA9OBbH7GKUMCBf1nSTiVxb+YnEh0qs76srbdZ4ZVE9go+REPecErs0
hhsJH5Qnrus9OD6Su8zeR8gO8FLNvWSlhNF7PWNhhu26xOwiDnlGYinVWjwac5oZ
SyBjkueMCK+no8L8CAQLtombEo/afjajdgLihOc7qDO0unWRqszuXod5dP+f1NKx
/YbdlANATfNUXDRQ4u1HwMjL7ACamjz00AKfRs+DwoKLg/ixv/eQ7HayO5AKqD4N
P4H/sfsSvMS0S9nHSn50ExaNyi/Bl65VklprzQo62DSFCwZE/qhwGpLmu5JNGLTW
muAAy+c6DfPBnPeZss8bZ9/2kGgiZAqWmcpCPMTwqvqvA5m/BJtnzGGoKvOxXMMd
n98F6Rx5d6X1K06onx1snSr0ElvqHWp0Tigt2kcHEPnOTsJqt6Cd6lLIejPtI/Cj
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
fxSaKobJ+ochhGIaVVNZrB5c7WM3CPw0oc3dJyRpRZhS48VpSC9apAOOYq3ZxwUe
QIyGxhmEmxp4hgs9sgN+pXowpUU9/1WqS5jF5qw/UCtW8EBoDs3F6BH2wXKp5ABX
CtksPNBKYsy6t+VOMcmk9LbeszygDO16owVgandB6xBGy6mpDsowP8jNKoPpihpx
7/cFIArb1IL5e29E6HCnRlR9X3t6RhQdeMq3nRZ4PP7dzWe74Y7KbgbLohb6Oo3t
imjGwX5aU3DU67cWvqBfytQHHdSJKtLWNPNqE/O6BEO6a/0CMZe8D2L+Txow4k5K
rMci9CidQiU/yvYRhnuivQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2912 )
`pragma protect data_block
avNM9q4Fo+hbInEHkUqWUnqB3qQWCXmltSKQHEYy57GgOiigJplLkKD1iaSexuh1
GO7bp/uDUeY0CXCTK9IrmPTQkhBXgFjbHcUNgCpr4zF26iqy/6MQNheWQxwhJBoU
mPvrnHOGTbX9E87/lafTr2CbZyxXeEaYN8bd3Mc71hDTNhZrANybw4GymehEqI7a
6RInGjdfvIYDjsVV4iPebGO/3kGb8JXYKZaHVd62Ls8vWiAvLcx5TrPqD8a8DFTX
ACCB0EO0idgvOMy0Dyr2O2ipujdypC757xqOJ9kkEZG/bUVTCpBXroWmLnT5pais
1hQVb376nqatOPGWgKEbbPEtF8BulSG5wTUEW9bPCnzgPbjN4DYtF1TEjP778sf5
xlIX2rqWZ11wTmw+uF89aXm+sm9Ndcwa8CXoOqQvqllI7xh5KQJZuGu8xYO4BG1r
PIEKKygz/llmx9poHEeYCCfaSG5u07NwaeJsy+uMdXMNI7LY/vf3Se+slhT0iU6C
BPkI8/GCfA3L3senhogsEWTTRWPP5eu0Zx8dQwTRLOtzIvepM4pCuEDxaIC+YfL+
DZ+zrDfpKZ6c3mxqFR/13+SbrcrxF2T1esk3Rzxz81+WK4LGav/I8A9wiMVVzXpq
FfhAdwkvU0yOOB/Dq4kGIEnH0GEQOjBWeJ1AisraSqx/NCFxSTJ2BB2Iqj0ffg8d
nSazWLuZNLmeTc9MB5sV/MPcJsGnUaF0z8FdsxaqfiG8OLcFa/tf4TSo7Z3VrWcx
S1IWoh6kV0cdL+KWf1X484BoDgPt8JY6AXH6V+ZmYYAfDVjLuPnU8RBNSqGExQpK
dBYffePOrYjoKnDUgUr/0vKfC54Kv0sDM88PcmLf5KetGrSjXjBYZ0NPN3kF5Frb
2XM8WUTnvKHSVmiKGv7EhxXagK3AcNb4MgX6Ur5JfeNIvTb6vpaOp5849XJ4ar/H
iVv4ptu7UZCpYqt/HOhoy46xgJYoz/zCsPcy5QeNzV+jkLTXP0m5RSW4VM8Wk0GJ
T8xTtff0QWzFeL/5j8tqKxuGHCjKAm0BLBDRAppMdmv7IOu4nIZRUH+pHKtK40ys
/lpvsInIUvC1Iwq6QICt9rwM9aU2gzKaUbbbLQAr7HxNuPjDdmok8owX5mpBYVZM
wfmxZoSZX7HAEVNpGFN4KOHbaBc9WjOae7wlkQAbNuF1WRkb/qbW7lArNczaSVds
nuhsjOfuStUldr58pyOgn2a5gdb1xtWpF/QYEOLQ/amzNYOtMEZBrLmgqstcgrBi
+lkC/poZniLkPzx/bX/pwtj8f3d7kYmYxwnEAeyDhkmJpbQJxJ2tSkaQg/PZOsjj
2JBEzvEsd2zrbSHOBYzvicD8c55ZY7bs210bFqaSzgNI+ZeCYEKhZ+XCldORCIr0
APx6RPcdefviJQ8yU0e62GPOgNzGEi7Y/5XHR4M2HOSBqIB2ZGtBgVSLST2E+Fmb
v/gMGrb7Iu+zo+Z2mojaU1XOqq6DJSRiabpXyP/7vh0e5UQExq+Aq5Wy+rOcktDr
N4I4MjssFSQd/3Ez9hweVCYE3dj4+rQKzCM92APpyOo70kR0EPQZBoXSEButT0VH
aMjWWODjNwXDrA8zXxi5gIamBV0P77Bw9JYtCJPUirxMNTwmSIp67KdR0AcFX4tf
vSBJN/X0i/6KtTzHYayYoZEKyynapmu9JrPq26zAlCd8BMJTsiI0fYslOA++jk79
EwMEafWid6LXnOHyAF6fK7v6DYjdcwY80+mDDu32VE4/VPM4jg5m/A/H+TU+UEgy
/9kV9UTylEqLlaiG+8JXd8KKrUOltfsjKRQTuIePH62IRxnRF3+9amrtddY0FVUh
ODi2BAnZjVH0d/KizCBdpJulGMQgyqczFNdPp9BNPqGLxCD1NrHod9fRGjNupG3o
+gTLnShP4dHw12XfxmBWoGTf1zJVvFIIEB1YPl0mDGTbsllU3Ygh0yaeHQ4iWWKx
2m/zBCeBqWpGV+zgaMaBD6ozKSJLxwqfFh+iIwSiINJrPdgNxHMHMZMRdmTbcl3F
cL77Iuc0KLyKAA8IzVFsmh1Hl9xVHVv33LzTgnx9Vgp89XqhLnnnkOucoSF8sqYg
kVy8XdQ6JYK0oL8oRMq5RoJkbZbnlbEMnGDS5oloSn3Ns+wFJj5NKh4r8ndErVAo
phC2zHfIqm+PivMLialBiMrLABdLa4Yf081oFh0IHcbyuxw4e0o0mDAcis7qoZYN
69bK9VzZWTMtUyN/q5RRqqG9lnOpeqK6tFhFmViPhrohK2w1ypshC1mVAqEDP91d
3tBpCz5vd70YKQfexzHc7ndnIbj7d3gj908oP6ht0a/IBKlADVDDFamfOiARPnzy
x7ckOVOcIXPahVhrfuqb2cvIjeWS3ViL4jKiYMnkul3z/b90D7Oftbl0SIi7pvcO
rjlrWo80s65Fb+UDqFI7c5vlHNHTrSG1z6cQfC3vy9ekJ7GY5IJjd5ycvcoy6nJn
V5r8Bq45mhjj5ypmZ7n421JJ1WkOxaPNODg1ItjiJg/vdiRvFOMlY87xbHMKdHD+
JxVYoWCJVpirq8WX0FelcZXRTdkSPHYbCVjvtTtFEBAr6Ty4141vazqaLSygzIVT
ff+qYqvVBYJnSzUQyvUH0UvONYhDSSz0mwwY1tMGsg57527CLGMmeRQzIizYarTl
ovYhtEOm9Bx2IstehEVp/oh3xitKhf9ucS/+/4JCbRw/zA79IQoGTTftjywWb5VD
kqtEYgJ6rsWevKAYQLU/2YEeQyM3d88lJQ88W/HqyeF5UnML82UcXN7wT2g62wZC
GuEPVL0IDsOjCV10gWJZwOYq10kknd7Umw/yIuKEgIDXjWPx1SzjkeeTi/Du5NDN
WOlXzGY9Ag+UOArCyHP26Mq+TIiu2cXEATVB0HUGlXiGFgcdlj6E7zH6nLLzb5XB
Pbjm4Ifp+T088N/pibW8FbfKdzQNFZjMSPlWP+mxhT6OfI+CdFPmCNKiZ8/pShD5
CO8TYG+qVmMB+A0jf5PZGNmeb47bMj9ORehrhx4tTEZtw50g01FXKk+gklnzUCuF
3j1iulao6aA6bbmmgANeIb0acTiZ81iXtgr13ZZRspi8PQNk+Ql0rG7OYJ2cKf3C
7hALT91T4YzWOI/rdY1vQjHH9cHS06ch/cV29js/icWrM7mwl4fmJE8xYNgmuPLz
RW2HSCqgGRVCBzzFiJkwWZtwOmT10ualA7FpQuM+yLw90k48VlttODay49OgQXhS
10ElgUBiycVJFHmSD7VNn6iaOGloWgA4m7RKQ6uCyAwaJDR4ULeJm8erifTwRfJa
ZVCRE7ujQ2oerpyrHhz4GSxRFkNvQBEVse1nG3qo7C3ljp4GNGvFUip0ZzpFc1iS
SzHTooBKw4ZMjnnJH9dTr8CK1khocz9GePVeAiCNn1zNP2+Paz0dvBpTKs3K0B3X
iKq2+HlAO80bVS9W/a0icLRNpquwL1EPDdDrVTgyY/M294eUDD7dujZeKR0W9A4V
7J4bQxrfYmCGUWnkGpj/GItkGnh2AzqCbiIRb9MEqs+Eb3/lGkDGjK9NLS62Lqrh
YbQpp67NCZioDfc+s6np7BZdQgfXig/se5RneXu9Y4BAm7rJTWaq9jc35GCab00X
Hi7CHvHiAb4NS0NGWONZN2S9MngW3QE7ZxT/fWORpVPQZnQQvH8rf7Byj+ubsScB
X+EgcvzlrbHG5XQx5ysNnqgtv7Pl2E7VnGnHQBCN+gOHJ5CjT3qXyqswO0QwnvMm
oMbOk9CDOQG8OypQCodcRW7dAj+x+VGMlshzf+D7s0MQrRaKBOlUyYkedvmsd6y6
BXLNisrfFSRyfqvTHtGYRmHOqT/Nkg906zIA4sHcKm8=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nBPee3NySvLseUSYDrOuV8drGC3E5BMrVIJuehVwKJEy+nofmJIambbjo7EahM5X
06F1pQqEHwaZUgpNGpc8dW79yduduw9uZGpv5ePWHHTe5nzHxV5vcOO2bKBupWAW
MzYMUR/rIyjy+uLen4LT4WL5x0gPd+8ylIsb9NwX3LIdwPMmAOyJ7Pl3o4DKa/VL
XPi0mH7hJWkBsiYRIcONFMMd1iffw4JiH1wvzPP2khF730HN8cSRJkR7ybv9L32y
Hvyl34RvtBReJJ0UJ44Lr2enNs32cAWVgEjon6OOSVlZiUJphw0pF9Roq/0PCO54
AoFIIfja6RKxTD+cJfdpiA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8016 )
`pragma protect data_block
svda2NtEnh1fcUtNUmkscvS5qNScxkdg7GJrTb1xIVOdREbmFp6YIGcNRaMMUXIy
KT5MeI+XvnGAEuJWE+jYRpe5CDyFz8i1TJviWmTiNwxQMAGQdj1fDcelQjIUyrNR
wAjK1nAPl2R/gnaZ7oH9+Y6PznThnDWh9czfKyTbFCy5tqM/or9OWq0XQzTjethh
RYHlW6mqQS2Yk5qIe41++43mif/zEXFqAYGdgINzNWhZ/De6KRKZISKBITWhIJHQ
vYvJ6JfO+2m0X36PVlB4hH4HVTdV6XV9MDLweds2ZKFDFH3tE8TKFWcWPZp9jpzn
/UlDPOz6nyhUcxHQflFdNmOPmYJX7R7I1WQmeAEG5HzXiWLGwFwlnsQ4wdjny9BG
aREu6U+1epgyO/Axeok8HduZd3t5OIW9qRP/Rsy4n7E6/87W0buj3+KQawcYTEl3
2Ufb9e0NnDP81Qnw0cJZyDqwSFOmM1gKrD5RxQBKZi6iAqsvpzjLkurkNp25svi4
T1nDWpGtspiJYtelb0PjRy5elix12taNHRb2ncbon2ik7ZErgxo4BdwH5ARbnVSb
OO4O+EeN1uebQHFe3Pnr3GGw8KyRuP99cpb1E9qyObNmHXAvFIWJBeE8tXZvlLLr
htktFzznt3gIMgNWUelA6Yas9D49KfHKk8x7Qy20gCLkMsvTymu3thoY2PrfBO8V
0JcO2cZf/buf0KN0Km1khkjddd8x01OYsdT/JTzRgEeq7JovC7vyBzpRrdGwe8gc
Fp5Q4GmeWDbhaLaIrj0QNQc7GBtsOe4cj6mHj57BKGPNx6217nG4gHbzSuYV+NLp
C/FS8e4Ox/+XZofYrUWBqjKwLetL/KKjzvcMRPROIOcowhsJS/dUR+EWxU1cBAR0
0zQI2pwPu4PdakCF+ova/CrbnsRRsyAtWt/ASCYohQKic4uuG18ONdHTsO6h1eYg
U3iS4flcEh3LV43mj0a3fB0oMyiUV15cTwvQO83fFbOk4LupqLcuM6c/Y8elxo+V
P8QZzi8d5HhsliwYt17JJX/1kntaz6+GTqy3Pg42vwZ4dDXIaTvXZ9/9J79rkmjm
5wHFlUPLOiG8iVMq+khXrDpRIgU5vciTo68jvX8d4HpCo+OK/69SHmq/VN+LazQ5
zuy1M71MdvEO9ygdK1GR47pxaiOerqVmIeBh9yPap84dPA4xi17bcyXaV2zdDCGE
tprib7mgs0dmWUpb4CvnumcKtXpIlkoM1YgGbuqHHKyaVSEe5RVFF0bJi4QojBA2
CZ6MogcOV0Ks2dDWbsLk/w8tJY3EdmuImKbECIflzPLUm4awnx1Z7uQOagGSaaeI
cVx2NcPpDH4MOSoXHJGTa9WFWmkfmnAGcAtUZX8IBMFWLqhLO8onZVarXMMSPqOp
xSW5Bw/2CTiSghBFlK8zVILIaVON6/1o5udQJvto8vvvmsRVdAZvFkF4OWNIqm5Z
cK6OTpFpQ40XC1gyfkstQYhsA1aDVGIHCQUskckoMUheaadQmomg+WtsM9f3BE9e
ieQbR/qru4RNh710TALQJbb3eXG/JnPwE5uzZ4k5Ns7AxDp9GmrJXsLxm2UASWMo
08oQ1w8ugKArQ3/X19hmmg2lFtL5Ib91crezawPLk9hWQ9TdnhF+AiKdqwGyLil6
g5l0dRj77ECHkmey1YErdnFJCMU/XLY6Kp0/zCuEQKhbh/HKaZ95pXQ/OoyIJ4vw
vOCIPagI3ucLq93K5ZrGNm58WOMSW4nvNH/Cm45Nfxn6r5igB13A84ZhfpokccHQ
60s2R0+pZqV+o7zY0yAD/zh6vbuYHRjhrcZypkXv5ow1WsY5DgEr09hsjcDXwY3N
gpjZppnEerCUwrdOqEacQiP8+VIzw0O05Rca6AmxdpLNmAGQhwOwWVa2H08RMYwf
cJqvvG5PjZkvPKDxFY6n2U/PRJ/j0NpTkud6KlwP8FLtddnIGTgRMj6V93S+4SnT
DLyFMBQhkAMiJ6QRQoAhJyQDgAM3npZxwx2hFApbg4N+3DeN2TmrX+5SEmDf4J9v
eBFaILM6ew/b0W3A/1ulB2MN3DvYkO+sN/qZo8iHrWwhIwj5EmG7oxV2f0xCeO54
KzHyHxMmA4BxICZqx6QAQ3gI9G/KT8NUNQ5qqUHz82o+IKMJlZSKaG6krjat2T+d
hrEiNhDTtPp0J6ujry0+08CdEhl7dGO7SM3atCwB3kb81Ipu/OtejbH8jHQorN9c
16jG2GFIMPJ8eMA5abpTowf1KuPW6TvDUeZYncByPtgsfUlEO2ykvnPAchek6eft
UVV0e6eNVLH20nqinXgKFXR60wQ9HpJ4Z7tJuCPFDBuYfn1EKxbHyQi5o3c9z/EB
N2R9P6bltr8bQ2NUlthQTj2TFAEAXu5JFqxVhbvzGhgj1PtiGG1qZq8lCLoBRGw0
z6tvp9w1vGgeMw/1PUPBUwPaLKw2+BmG44wRf639g39T6tztbYgNC+G1Pyekp9Zr
QMKx2EJYFeQFkx1fRW0XqhAcbbUu0TZqyOSKZZ7Gr2+bKLAO3sfxKlQTgGEl7xTM
048Jc1OOmyKS+GdpLtygtPhaCq4yYFmRYMDpwNeDsdsnb3bfip3jks8eMWiSgtLe
9fdmPWsBzBxdtzp8ErEm0tGd2s5vii9bWjsdeSSuapQi3YTnNhU/JoFokebR+9lV
g96LpLifL7k2DeiiUQ5vRGLGqsPqBYUQCmnp5fdDihMfKXFzE0wUmcOTDMpCgDhF
LJsP9yzhTMutWkaccRcyXmWCSwbWJ1KJai2fi2T37KiRCRNuCOo4L1On/eYV9D10
MDKKMkRsVEBneG6BNjOZBWN/IjlGqyAxzm7hkAG89CdJCUULm5G/bWkkeXgaHmZJ
LLz4rU071L5zO+vPfxpSqGrv6oWHeO643vN1OirXvN6x6jFta3VPd6IkYnd3+hmP
UB5RQDXW1KA6byV/zLEtteeYVy3+SCs6ZKmxEqDWGcsTsshbxm1AFXOjOpBPIP6C
RafBBozJzPwpXAvw+U83gnzv00rXRrIxBHgcvGQf1SxezihUAEWxJgdFwNnKqv+y
VwnYX/QVxxcHKb3eOD8IhSdVRZ3LNFLpkwoeniPtVm6Q3sPxp2gSnO8cfCiAbEBK
TeCZNsVkgruG6WLW7ej0FAdo/UQBi+H7K/H6gfw1PjKwSiwX9ycuEILCquQhtged
4d/f7dFcB2ygFXnrIHw8j2vYIYXGiD5VBARFAnKrFBOEmJsX4IbNUjuI8QpHmaIb
RA/kz+BR6LP8Gvww05x2kVsa+MXDi21pl4QUuRVK3eTYh1mlbujjUKbNf1sewePy
VD6l2aRSuTk5WPgFDtr1j2L57c1mGpPc3A53XMhBtKRil/tMD3j8y+k8QgmLRdFo
q7FSJuoKDBvHvajvzdEy8RPhG2svEUlpB/uVD0b4og/u3jBmYmNWXnmrm8hEHF2K
zxGxMdnx2xdlZ7j8wCXo4AdMQoDBJVUE+RoG+Jk5KFb6KXYT51sG0bMkaiVefVt7
80Vz5NT7kzolWeyv1MKqKiM7lIPjnke2v6IcrKk/Bw1RdmUJJxFSxgLSqM0E/Lm9
mPj946oFL8kTgGLotwei5L8eQmZCbFiuRJQag7l3rz9lTFMU2HdTRER/b8wnYhh6
9OINUTvNE4Oyl6SNVGXMMkl/589NQ6xUPx+emNvf267GCoO6Rrfm9mua0WxERgxb
L/Ftz2d5/1Tlm69CZa4OUJu2YmTYwFTO4FvV0DtD8NFpvh4T3OBvR/UokkzpA/qd
D/woaaLp2CsMyh1IMqayGLeN9vxWkmuKHB8dEk8/5VWPrx23BVXoXasZLD8/N9zD
g9ZYDxDS0QcMMlxevsulBvMv0wB3G5bygC4Nj9af/UNApxf/YssC4MUfPQamjttG
3P+FWAjSGkEtA9x9B0OnYWhXVoQtzmL+LH9/cn9tayqWSoDaorKCNrWyvc30y6EL
j7lo7+LzTjcWEzP0IiYHUd2CeLPB32Z0+POCQhgxpiquL0PZxRCEMzsQfTvtvn4H
BJyxuAufaFBxG6/f9/ws6pcYgA17yQwy/y/mPTIFPcttOQ+4E+tknYaYBiV3Ld83
X9e1uQ/qKNeSUjSG+mHx0RQ07jVBznUAp9HRC6GFBAHytdOf47AezDFuArKE3FS4
+DFoVHDiXUAs7X6z9gkX7dPlrXbULdNCwCm42lZYTqseIYErwWb8JLsE7j/6oYpx
7KgOibWQGljVPLRDX8h/QASHMa/T228Bxu+VJRk9pijcIwo9adFbdjWLvsZDdEMh
1oWup14vrSztM+z6D6AdOwnHL+Cbcd4Rs+MB3f2Gv8P1xI5bwEXdtbu8CYj+i4Jw
UsOJ833bfsR3//0+ZmnrxVbF62AX6rnkoKbdR40k+JueAp5HgUY8HnBR7AI5WF+2
1681ac0PLtyVVMZ08P/+Pbbpeg5Ye68lMlB/7K2HNUj2basqpgRLZBbLB/ro3S/B
SM+4rIReaIAdFrR6DuTrAoHC/x/D/jN2salUk4Y7fhETeMHa+5AtbBhwl+uufXX5
WtmGiCn1aJNwTfvt3iYIiyGG32uNkGZwmnv0aaymeGUHFhUgMpi0aHop4ygCO1Mh
b0MJ6YE8K+Ajon8faV9kuw5x0I3zfwHhKReMwd/EuXCVY+wSfzSyeqhQUZRGxkQs
sXcpYSHG8IfF7nmYdWvRKccUkoUf9nZ/AnQOqd08DUBzc5lHC3Rh4FngnyjzpVTE
SaNl6xZ4f5k6LuPXkVxX8edemnM0wQd2Jm2dfnEYWcBBgvdSrfHvceBCF/ojvrpd
aQQBN0BOk05OLxBTPp04pxhNXVk4/tMQ+jP5WT1IURE3mq8d9kyDjOePMdnLpMkB
4JLjZZ5aotpCocLDm0axc2+OPwLbgFuGV0vSYrkKAtmCDw87/Sc7YCEYPc4YZu0y
zjg0wOtiFrBSPOUfwcWweRFGMyGjzMgpZ9X5juMQImm047j+Vbz4+LQ/qgUnIo3j
tbmST+veIvTfnhSkNfOfqMdrdSkqPZFR5DI5VgWbFjbaAm/tcMvNY4w4guaIk3VE
BA4tJo5qhNLydyal6ikc5/0RafMcZ8WnAksXLF+zx01V+qk01RB2R/oD9ybdH8kM
EIpV5sJmbVPbEFxjXZaeQ4lL2wNKxuuLQxopv4Nf2GwgFPuqXP2BvejDh0sVwUSB
XAW/1jDeAvm0IPJvlSSkL/7kKPm2qvy2/1VIG3svq5uiBJRBELJQZey6L9sHIIRR
VcaktChqTKjRhIKXiLrpbYG7WC/8L/NTiUNVMUYW9qQkpyb+TTFAqYwSYHcTyWGQ
zynw0OVEQZ2O8+TqhQeh+J4RFvzbm4CAhAg/668tKepreF6Ib4Vi/dbxbMI9Leio
0uUYvCmcs8LICQ86IInsSeSnZsK4D1fnnK6J31zT+fb6xRVdsHpBBldredlXdppY
4dmEITJJ7SSAbdR8pcJ13CJFgnpdETo72DYb2TeV6OnazyXC54lcpfoMv1tVT6pe
uAx8uxpH5xl7+YyAyFToTsTJ5V+u2eC4oFMFP/FQ4kEA1Lbn+LgWPAWo1IEHHbIF
EU50xnP5wMBpZLPx0VzN2wUw4UTyGuWXK8JqiwNfqY5kvuKJ5NwYiP3czIZIWXp0
19COto41JUXaZSwhUPW/tVtJpTjjFm5mn1mpkAwLWP0F5r/nZiIOs9H2Uyy6jOvY
OdSO6LBhoNl8XklmXAfjNRgj23VfI3ssrg+65ogUbbp4gMV1NMwxeiaVBg6zR1HN
QKAM4WUQMIIakMKFgMOE8EXL4xb38jr8F2/vhsIur+dyT1q3wvZUXOVauU577WkZ
s+mRHYbTXXKvB0lMqX5Y02psOOCEhvgP4DZcRC3tcqrco59yGeQ8xmqsm0/24KxQ
g8xMhddYHMxkFSpG4Nv9yYckzIgjtlM67YYMHOKiWuZi/z50T61uCUAEZe77xtJT
xp6tzMhzm6tk2G/z/U8K3s1JklMGmiVxBG9gFtBmPI4qhomDiqUIptzKlfzxObVw
6nZ0G3UmmdEf7AeXghhtImCWPbOIVUwR8b/c7SUjAydBlGWz07YH1oXw+sq2ca3l
EQWmITQA70LtUY8PPD1Qg1Gj1x7mT7GhIjaoktsLZycTraRshhgG3bQtK6GLbYGx
Baqg6Us4wb0pmBtKJJrT50S9MO4RzLy/TiFndldMNs+qbRVhZrg/dDSviE5WMR2O
Vmv/4SbZZeTfNW3i18zusnZT22UChA0HYV1WB/E1F8er9lw4n59DaDlsSGySO1sq
PuXO/WHfvOiheDSbS/se6XCQ589uZ0qO641AC60G0dRKOEgZd314Sa+9+Lr3bIQn
yuQOry4V4xGcUeyqyhIokX0zfiblqYPCN9g+osSPYQzW3qbmGCrGJCLcgzMYcxoK
mTc21sCsTlo5Ou5qM8iUB6Bg8S5ZZ6TMCmf6pphQQ5VD7KI64tCvv2+CdzsiP/GD
YMuWwjIrfULFXBUX5OJBf5x9quZ2ctHN0cr0quykY5SphcMoko5ZT5vLywYZFr3k
35LCLb3eeAqf7C+vX9EEDVWsV4xUd+agZAkWU1YtMNreLasQLdfOggyQmyKyw/Rf
tSS+rmIn8i1yS4CYmVNnF3NkejbtRG85Mb+7OXRDuYyv3yNg7F7cyp42Bf6u9AA7
EvqNqj3DZnT9teWNWXuJ2d3HZb1mEeF9I1mAPJ0Q5A66+S0ZRg49OV4LrxgszUt+
TK8qzPv+lq4zO8zDnouuG74JXekzLO6luXqBna9vrjhSQ4Z6NdUWLM9jFuWjLeHu
APpXqbL7USZZsEt6dR42MUsNlUhPNe1IeE55sFslgIJE0RRuQD232+l74ZivfmmW
XciaeGRUQOqJdpvcDEZRQ/tBJxECrNqLH8Zpbx/EWkA5YXAPIp8l/Pmjkf2kOGju
3MLNUuMMvobwKUQqDNLMxLyoRRq9+G6fyDkpkurfOdQcVtKcsNqMVqZhBgnqiBw4
YaBPav/pIYL/HIFzyevlyW+jD1Uc/tcRuLuwFLSnCLGs+a1SQVhNPlxGJc7T6XSb
cP3aDTgNN7xWtHxS7wO0eIbSpM06+1W19yaAlhq5GygCih2SPGU1GUSO6HDcfpYg
HB5g0SxLjc+JxLaEXt4zwHmph3gAb7ZZHulroBX8k/WxLN8nwX8CYwTfVTY6magN
vXOEAOvT+IU2Kz+5Bk3HuR+woZ0QGhZ4/4OE4R9rKMGTATLn5usEfVcRyFvlFG+S
mqfbykJ0KWdyKf7gQOHZyHPnu6bd/hDBkVJwD0sFsrJJdrpX2YhvoWqoRyuPHDjB
ft4yZAvMlEQQujamRsY0o6Ako2sKLy6pPa4YtrcfaOIKNct98UBQY9kZ/t4js29b
07XEvtpcsWMOl2mwwygzrRg1XFIAY9e8K3stZHg87i1xLyRqbms4Zep8xAfzSqyE
1vAL/kuf7NFWWIDui5NIPDvkD2B3tgQa6DcsalhHnTP0L8Nixv3P/nPPzo/v8WOW
NsN4zTl7ra5eo+Y/2t6fUOwl9R4Aagw/3Rk78ygHBFmo2qm0xfudPMd04PWrGauK
/hajvs3Zeyirn3HeNklq+KpudLmQpOnEDPPPIt1aWw4lIkWLGjyOvvikrlKCuJyB
+zSc/dE4NY7mPD+OZU0TRrttYnmobVxf0R8rvgqXqyns0IqeNnMEAjWXMduh/xHj
bOTU7rvbrZTkpQqMVOPPRcN/1+V7nFhLXV+ULjgU2/gbp/qtHscSkWUq82os8APr
k3tLK48X2BEZH50efbZuZW+GhQsv8ISNMnx1rdZDIUNEhsCmjO38dnWGovbNTuMU
ZOEOscGzIviHZ+JeKEaRceZdTgs75dUV6DZpZACVD0u9JDoEsK8kYRT9cGlRef9E
VZS+NKJOWOD6nDyOSafEaG8bH0QRrqsHRSX+2FMLGcpXtRSomMAibWlDG5tZurFc
CABAa2nigpanWus25Wy4PVj4uK4BnPXqAKoIMOOB5Q2WT76IBIZC6RLmjPx7S7JG
SdTHgon7C0eITcuOCiGR3VMH4Pkp6t48RUfsLLVE/ax7MRgZ3gQ+94alXeaF617D
UxD42tmjafWfqrlI9zosC7vkCIUt2qTHGgo304aEzAXlHeNGl539v10dNfaAmK2Y
6MsCgeWUceiEhppQRgXDn42KiEZ1/Jjm9YD6Cet2znoc4x5H72ex82QUt7t1SLJ8
uD9fhNrEmhjjqO80wqBbAkjqvuoW4Uv74GG3+hITJDVniT7FL6MmgWk6rN+GeaAt
TI8QKhCrowj3BTNiVnt/BMeSVUPxYgZw77fM6JCv09s+lNvbzJDVTk7KDO4S2ujk
cgeM1Y98Y6SRmeP2Em1Vwc+lML3VX/+3jnOdVP7Ke5VFucqoywxGtIxBEay/toRa
WhQmD3Dn9wLaoFrRZv+UVnhetJ/npHqc2DI0OkA+gshf5gyKF0eXQm2XNouv9SfR
/K3RxjSjl80dKJJ+gPnQg27r0eqE1f3OaniZELJSQ9O1kdm6UGE1u09cmbx3/vir
lpg6yRExRLKRgyhcgeQY27ZRdqdbsNS/qPgptdpJV+pq7nm1Lenrvy/pfolvc9Ib
NvshUFZj54l+yNWQLGuDUS8v8BKLQFJqcwbC/iN9fxWdtltr0DvuANykHf9fiW6v
CXBBIBu0YOGxMwuU5qV60WpY4p1SNd963L45VCqQyDVeDXEAs3wP27OIU0nU9ePP
Ig9UQitsv/e9n6xxxyx5l+al/x+Lur3i72uJwR8oIsJwnJfexwPF4apwZ9fL+aPJ
eX9wpC6EJ0SRwGG9ko6DbzymjwqOJkqGMhMVubYlCjKTQ+sVJZVnt0yo9pwDolVW
NoCvyOr7LHyNixBeVeXVV2gtdvbOnyvl3QdA7Di6tjlFDJ2MgtjQeLZWxYrzy5ih
c0sy14KXJcsT6G/kN1tJEYQe0j2B5HY0SmqaiAm+VTDMBRxgn6iJgZkFsjdYbz6d
chLnfuosG6BgeghFizQWe4lqlQdGKQy9kR4oBjsutF3okoWhv4AbOq962Y66JtuU
FY36T7afa9D1Qqm+a2ZL94Y+TUPP+tDRjqX9lePkoLRHudplrc4UiT8bpW3P2KdA
10MflErUpu8YbmZ+wd9rNr2F8c5kFm4x9G1ugvgiK4JA3CTfwnSS6hOyU8VEKCVv
smgKIIusNclzf3uREkTRT6HTxtKjKP36auOa2Ko2aqlqvFKTxGEYhZdeEOCFXSDq
2qklTJkQBLHr7CiZITUNGgWAA+q8KeDbGQIrhOxZtCNEEik7EJgYbkFOLE2BYDiK
6wgA5Cg41TzQZvWGRv5StDTIMhWF1jPjQzzbdYtHLVWUfuuuCtZhMk3HT+sT7dq3
jsVROo1xV3xNHovUkEAKl86jqtYNiczBnGF/IciLxkXByGt5xZCt5kUmFX4vYFKg
tYLi8lW7dHzj/eQ3QmwjpITBR4tKQGhpGchN+kzxd5W2AvjYEJf1L3FeTrsiulNO
HRzxBa8R7z90ca9HHhDs3JT7eMo900CiOJmdQ7WOs23TegcuK/1/q16NsQoE34UD
3wTsG6Z1aOd5E53SVsYk/63+YR+vUBh5nEYksBMHsAPJDLvlTK/Q0c7PyM9O2El+
EsS2f5DCK3ndcqq56mCTRQjvo1g1cxI2+O7Z+2CrvDCMVP19Lp9CzT19Vq8w5OvN
Sao+h2mkA6ttPgF1reEtt50L37te+w2KDfXp18z1vOms9kryFy1zl05UCoyBmzB5
irAtShWSUgzI599Th7hdtFUM88s9FRzGGGitMzQcUnuUN7eImvkmAHCeCUlOQak9
X59QktO8AIdM/yCai65kGCOVZ91GmCu/rmtmAH1MZjSZyLxB3ryO8btS6i+Vppa6
8QSmwQFrJCkar5pDNEDXEaDr3EKWwZQpzIsvZ83QuokUgfI32cwZDeOeJc6mfx43
GIV4/y9Y/mgvrPOXIasNLlix+REXBnyDVEv33mQa5pcwcdJqruC1H1MzT6CSTaJ9
zaEvOB9rrhFlrNsjNlqlLsWv0/0lKjLK2ByKml28xGHZUUqlFf+BXdjQ9JLvh4tZ
tI4bZAt/ZC86bx0FBx9/qsZwsHqVgKlouOVq/Ts6OSJ52ltZjkgqZuf4r0HBnLWl
2gXte7BaUJRJAAHkZFynC11xYdxOgw+hAHmZTSOFPMNsrwJqLxWjEJIgc0GmYwGr
8lti31S1xHtAF3Fl8/9bUOsRaWE3Pxq6jFWEDB22tAKP9xxPmX0YYoZASi5cLCYR
PNTAoZJuGY6fBZhzab9ce25dcwd+af0e5cB6yw78Z/o0QnebbT0Ufid0W5wDgVEE
CRQuArH8h6zWnSe2LOC0oAtWXpA6Fa/pcV2x6pgJ12mArXXLkU5fTkeHNubIN6oR
0Awm2AjTtPg9+dinvMnG9EfmkhR8/I4vu4ACdGQSnXee6/VkbZYKGP3+QKVyPj4D
EyLt0ThrTd7gxRwIgFNGu9mohhzoYL2Gs9UQek+w0pAz7ydF6dHsj2r3x55xGNtO
mEBojznMYb2iBNJ4U+5LEpGJwiEo65nrba1Bf+8cxEtILiyHugvEPTUtRA3Ewx4+
yas2nbxOTh/oZUeBBKpIFJ9SUIPWOUfEGE14zh/Iq5yziNN/4onDNoapB/FZ6MFN
EL6iG2GRbNORuDs1ibWn4d69iEvCHUZjzYQwvx37xJx88kN8jfbnCdfQwKtJzNlu
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
PcQwTd92ZJjxJw+SWT79lzMcQdqlMfWLpgSFY6ygiiNYHzrYBGhB2zPeaUFMzca1
Yu+8v/ijYE0LO0CxLZbDuRFfJESc+PYqfbIfH4zcxNybWDjqQv4fAoJg0cihjS+2
v7SxajQ4cpm7Ku2EIzg92oVO1jn+XpiOh1TVC0iP7HvqeKu11/+WEzZ1fkTEDFrW
GZmtzD+uAl/+NCWHtx2D56NS/Z1pLlYsi2vgMN8ixeGj1g6KagX/CVeFOkXbqlZk
URNzL3z+AFAAXW5VmdfHLKMJ3ZIkcrhx+Xp0y0aKLfaUaz5Cs3eX++YcK9jS7EJ+
GcYlTZ0yoyAY+PtRuHssjA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5392 )
`pragma protect data_block
rPs7M5HmdYEIBVgt4+gUHua4XWJoTQCyDQ/lMbckXHxjUBXYjvIiNJXUoZzwcd6a
sKKTh/p2F2UtyWIz4HwFS7RHBxIevYf5TbTJ1nObO59TXljx+lF6q2Q9pLVw9gFj
ksIxoV5I2Fqv04mFt4unl3vH7G1Id10i/GLhilvut9BxC84IIdHpVm6xUMuH/pjA
5oV4I57pK0+tejmKU74sC5I5kcZzbxCSUKFCEn7XxfMN0kFMmbIOlCVzZ2vNYzA3
t2Rr1S29JFlRK6DRQTEZv3Dntc/DcejW6UrzIdBAJjVAG9MOu2PZJL5+qpU2GOY2
WZ05o2JjTBZdUlqVPUqsZCL2RSvbpc7mQJ85Ac2mvZjRcK3m4rllIrXsONRSWHrG
/1nFUo0XVukgSmHXWpOqgtahICKOpjugbECSbsbMybYLZXYCfy9UojSrVqmbcmNw
e1jLEI/WHoWRee7IE+vxP6Pqm9Gd+ehwLY2Lq3mdt9+U5pUeDVRt0fadh+TA++7r
y1oY4QXLqwssXKPYDevLZRv/kBe6fUneYKQSfV7iQSx/co8LrM2u/LiAcIOgDkby
UXwbuncTv3Ccaa6ECMqbTfJu4TFfhZazqZxMarWICuV4eS11DyclmmV+Cjc862ts
JbsIF7Bfpr/ColMKMH9qNbUNsqowc7UhWwcvS38GJQjZun3Bs0xPSuO6tjKFBJF0
6nxMZMReYhmZQrkQFDBM41oInx4CwSiXC/lVEEQxaucNPPuMFGOfhSqmmsNCUl+N
6e00d712OZsLdY37umzJmcFCbI/nP6aWEBbCbyBVvfaPKAL7Rce4eC0PII6JFp/F
oRlF2L5LzAhALwgGlDoMClU4kIok8cEgx+MJbuKds4ADihmzHIXnXDmNgSm+mlFi
+/SxKKZKmoWKWnLDVH2klP4hmgrLaASW6lib4L2DdCzgzK83EsxLenA3eSaESc3j
ZUHD+LEOT7TXDSRzuLmFMzsZt8+lA3+EB7euFeZN+6BVggqBaWTcNw36khER/dnp
Ow559K05+7VnMESopA9ZlXBcHU7+euvEklTX+q+WSqLc3zB4ij2tfKdwUPjTwOXM
2wooARi4uJrsffDvh/vChTVclT5LketRmoGeQ0wvvy4mw9jKcI/EvDV4tFF1cO1K
e/SyisfFMv3eFuI7+kX9LCH4S/zPXDGdRDst7BAsxBPVAckrgOsEDgEkLvUV3zp+
A1SNNGKwmPNfj4t96vX3xGtAmXb156LR5zSos+K8/FCXJpEQyWvZDPlwY+SrYgS3
0udEog8Hdex+ZzrXceCwM0jYkCH9bR7TkTbsFz6CEqFwzg4sttJgnpAP2hAcD1mN
E7gsgje+w/BRjCkGqCLotQzuo4O9sYtkuFpHQFaPOcxQsidxq6umpiYEF9eI3bx9
dIaGPwVuVYyvLg+EB34fvNx7IMifE4hfxVDh8Diir/hB949juZQ6CHamUu+ZM/QW
WsdvdNEJS4lq1HPj4jzDxsvC/pfyHghkTSvl1iW+FG49MZY9cvcauYFUAS0H4zSZ
gy8l44FpnJpH8DLRyHO4I1OwM7pEOozaxHb9YiIgcwUk9/W8Cd7BZxZERQPxE1r4
op2r0xGW8rLMPV+m20spqltv31R2XtTSy7LN+/SgeWr9J+bjzMwP7oJd+oPtdyL0
kGVPpXnOYgB8qXX0BhjnNdbv9MrB/lf1nKtB/GcvHfUihM0OWqdYaMF+6QjmXeyU
QDGI6VJn/w7qpTezoS5ze0D7t2Dd5bP93Sf6JQhW4lYHNzDJinB10j9QXojWo8k/
LF2l6LBsMZxGDFLmoaGqd0TVSP77cxB+PQF+QKmdur2R5JA2Q70YRjXsa9ScAO1e
rCPVS+m5Fy1K+f2JyRobif9YTvAWSvmokRpBgNLZzO5G9t0/K7ZMhiP0V1EYZA/J
NXfNQ44bpmVaUqbaBRRXuVuJgsiPNgzGF57ZKFYpVI+Apc0VEPWuyJnVMjbgdL5a
gBKsing8gBufdGxCA/9WcrKXI0kjqpOKO8G9dKHKrf88mURWX3HfX+7XyPLkUau3
/KpPTcAK6WowkTOm5kg9Nx7IXsiyIxY2gTqVpcK6l0HbUYoFuGdteMa3WOVtvZFF
lxO5+KyLUepFT8WTI8nLxSSNq/kbvjOlcpUoq2Ih7fpKFRSBQ30fx7hidxIL2nQq
l92AGl63uLDSRA6hGUl9oWZ/U0QAcqIgayRNaggZRwc39YVXCqWwDiAJeQ9AOs71
XdWo/2WE8t1ZBZQDRO3OQyQqoo8zE4vEstmCMbJ/8HTkE4uLEfihNmhL6ku+Xtv7
YmHR9LDsbEArO9n5gsSV9F2hfVT6PzWegx3ORWofZjirJ+1LblerwEMsilmzRGIt
Tq8aJccTqJhGbZ1sPvRmgFpCWFrJUCLSJAcibBQFdV6zSuKbya6Xqr/QxLsYwmGu
8u/M89mBy1tDK66pXXduxkkILk2wywcs1wX5Mb6hr0JR0bq61qRf4kidYf4Ig9AY
nHXYSykzEwV+EHpP2aFgwUC4VlmVISPTie7CtvntSfyxTHH8XM7zsW5pNSLdJbuR
eKpQYSDrhX3XbILThod2hs/MBfPSMWTGEARTUFGPtXoFXsrirY7F57EBcOwMaMdL
le+3Cf1DUVSikk2X86WaHzfysIh0ihbgSeVp8B+hiz2P6w8jBhmC5t4hPZUl8W/V
CgOB0ncSs12I7Ux8ieraMKg8ACSuo4g2W0NgztxVSffyZf51IT8t61P4sfK6MjrF
fWTfNH3i86Fc5AjoG6/Vee1fGfyVGPnE9TCJOiyE9F02U3hN8HY3Mcte0sWixSMX
BIeY5qexzytAqpEQjRDTp67s1j1jHDAyMMwAleBO666PkbZQSwmgV1vtpWWVEYgr
0hrmKwvhJeCBeP4+3Kl23oZLXiwLPfJQ07cRg21PUFvnntcWOI+V8J4Ot6y9GaH3
0RxV8fouWPO7SJq889y0EAKEQuv/Ck63sIV3dBrqOIvzrZhsSfAwiJkVrbPGv3Eq
q8lFCvJGvig89sesRa5/iE5HutUSMUmpvngXHf5ubMi3PMMVFxfnKPr91nZWKvUF
VbNN34VEcBHwhNt5+0IjeLubmpKDIxCnzpBekBkYkFSCU9mLF5YUsrBJtkQNUC9i
zKUIThdaKWCpdCmC0l3/w6YdwHlllxzJQVkbF67t9x4LD+qxnQIzAKsTedM4lYP0
WtUN89a43TCoPf9JOG7mtcZ/YnJx82gArojluyJ33pTKsdVPAjaPX5ao6X1JDxDf
/2cMisUgfdQRIsxBMbWxzHmzDztEiQg7Izj1nwTvjDY0E6UU/GtS+uIK4xFm0tj/
XWiWdnNIwl7CTl99VemKIYLSQczhEP7XT1brkG6pLFOmrnr19dkBKq3mp0W97fqm
Ir1DkE9qFTlK2wM4txQtcC4msKAoDFBsz6Ogk2cqXo6SbEcpRO2vVTWLYLNUq4fn
4lOMUuAQsvfOjj7Zi49kA7P4zrT9J7tpSShf260MFoXr6IZ3dbskyQasydWDw2yn
/z4fepEpvUm/PZ0Lut/goV/TRV4X6bU/1iC8oEI1waWlyUDieR9Gjlw5hugmmkWE
bb0vXczvQXphikSHOMWls2oL7nDvI4dr5LPWJaEsI3CMmL8oCE9LyOFeIqn+M/rK
pS1PXBoFu/DxaDPS7BOBhDF7y9RjCrmWWF5vqnShJRXRH6q1J+Qnat/F3enyivZt
zL7fkuM9RD3yB6LkXmX4wTEB3egOGgeEpxQNwbcMLF/NbFVwrlYCXxMTjpvRkMsc
w3D1O6mn4ZzBvpdVlXOnbM3MorM2ta6z0aYNCidZfqiGUNsb3qw5jVGeO2fXsuHR
L2+OE2hc23RrykerOJ1RfM4A3QuJlfi4M3I8Sa8A07ROeicLOSVJ5ES7IQFLdck/
aF2sqQiNUfonFK7B4M2ChR5ZKEgUbOogR6kM1IE5eU3XTo0tMlQr9qeSh0QyrPn4
20tHfwN9Ig1K83LJO4UdKLvL7goMfdHIYZNZaf6rjH21bPi864JtFYpsMDebEIH0
vp6mwRrLpCXewBC4ZDfQi1M6Y7nSQ+taXAGa6+rf3OQNhD3s7jVMDkw4FBr7UtXd
zvLs7MsKMVo8DpMoy8p1Ru2VB/OysCq/MK/kOIhzRoN7M1zFNl57+PiRWwNJkcuq
eFL+cdnYhNoN+0Fckhq8x1o2ywI8XhJjZkUrD58Os/RVQEqUgu/Uv86fk7IQBEm4
W0ugnmsqzHVXEi4PiuXBl2TWU3HbOZUev6rdMORr/c7v3teSic5rbM7litXaYTO7
d/zMO9xZfULAiIs75ETK+47av6JEi1pdTz1fIfwtjbl9Uk41a2kYQsO5+FdBfGMn
nqV4mycNt85g+3tPvr1YfAMoKzIZwD/bknKtIF7ROuRjyy58+uesoaS6QbNAtreE
d7WirzeUMv+XaZreTZEx7X4RUCx9XDbDdh/Yca6iAwscSJHbjm1EBhM2Xbcq8Z/6
lTmCfLIyyhk6MkT3FSL195ffSiODXO7emCg9LrDqFRlrRn0x7PEKjAce0fjUueSp
VUnyrNBUpjTHxsxFMcbJW0chiwtX77asRcIhWi/VGn32SA2CMFR86qqbk4MgB/mW
7UqFzX7W+1GHt01bsKFslN0LbSAAnGZk2OHVg9xfr3ZTziSEXQDyWFxKQkCO6pKL
CgU3y9b1pRsV+bHn+PlUM50Av6Ih//Kn71VgVlKQNm3W24/ZgwDHQH+orfswNpEI
y8OfSWMDKPABfm/xeTCHOXnpHI6mD/QdrHN7r8+UBWw79ar+JV0REAKU7quFvWvJ
DJNNlSJ4QBVqH//QXpA2/Y3FGPCTxf+vfoAkxvHL/yzxx/9uqtUzno5Si/odH9b5
P5ZXEtov+rws355lRf0XwT0EdLay/Lz4td0tV9G1IIX9FsGPPRqZPUr1+h2NsnB6
H57kGi6vxPfXQnCYiGsw2LI85ZDMIb19LL6tQx0MZcFYGv9LC/wgJOXeWCQFyxE3
xpsEhVYVGEOljSWXfvvOXSsLYyRpuZbuKSCpCYKLjit95JL0AnBk7Vk1cdeqXgG+
GTALYcVAgX561ioM1/LJmy4Jcmr6vtW6JJYYaHbFAQ0gduLizkAURmCxdG61KA6r
kvkGYyR9JXpm6Cti6mDQ/J33nTLZlfPuW7xwY6J2PRNd69cCcPB13AHB9id0wChb
oWYcxb05zHOnd4xXbb03pmXA6Uc9Cbd7Fv6YFp8P2aOcysiTDiUjDQqXDm2w+rH1
jSV0oL9Z+WLK5yEcT3cYmUEmHitVlDQo37lsr80HTyks6KOLmgdQ7WpB2JAC9Hfu
Dts09fG7QnPsn3KA42kBd1uLw4n0X+mMo1I9MBWmAvRKUWimO3SXddu7BxpSzLhA
jkoVnKEQpIlXLRgk0RWlGAklIfeCGaTZ6du3PP7aeyauZWVBb8W+jFGwlbYjiZO+
+PKZ8jaGI+CzZ41BgskJWxqJhrQkz0cMgV/boava9x97PQiTKhxonSi8x+o1cW+0
JTI94wpjilJyXT5ZztM1UtNwtc7iZFEiMDerKC0ygjQmu2B4JbbStQPdqRTqvN0A
ZFvKCskpMjjrnhghV7Nupg12tXvBdRPFZRB0EayqcCwpd7hyskzHdpU5UEz4Uq8p
J07p5ISJaI88V8K+djYd5AJUNmfBY9E6AR9ZXpvSGimTUKkqYfHexbKpfondsqkx
mJaw59G2waC64tlc5XALEaCQNehpv2F/qKe+lFFM4mJnhBs7AevcCUPl5Vhpzz35
CTzHu8sJYXEAZhBSojs9GFc4NWEfIhYYHWd6oLyJRW/560B2Wqr8DWM1K6wrrELH
F+mTu7BnV/wQ0WPpRm2+0DCEZhMKAg0x1pSnhDrA+FH2qxBxvj0nthLXt1tnDWMG
8hmUPvQKsXh/NLm+GRem1Ld2qCVLo++Ow3ZVgcIdpovVQBINH2NncxvfidogL3sc
RmrNqguvxg7F8CFOkNSJu3w5MHtQZeWEFiVpirBoj7WVEaBuvxui6FBsC06oMt/w
2R4MMVv/+gpeGwqaMtyHLLwOmCKLbK2FjKv5JyR7j2H9dUhx0hLtzWztetl8vauI
IWSdv7MuskoJEHRmOM1tbXtYrDqYqZA9MS7I17BysWyM2meyEx3OA2s4/Uum7XNr
uJEvxczodYYySCSXrxoS6KpyKi0CmG5sIprfy3ihL5ZmDvIeyh0FsCTXbM6NKKvu
G4aWE2o6N/CWQHijqLE2uKTq8Ibp54mm56Rny6XZZDghEGSyJl2b8Bc2/u8TY0lx
pAOh5ROVFM05h2t/McjA+ujiTw/Q+/XDUMYCmHfZMFfV8s1pqQkwIW3jZie+YQtJ
d6fPeWYCdhIaKZIwjgw7jDMvMjv9TAtbve73iCtQdX5V0LqJa6+3KXVCdyYlUDjL
uW7/3XnbjpGbIedqqTTvsqw9t4XFTnJh45/N4O5FUxj2tDgNZUg8GM7eYMEBc6dn
alflP6Jxji+fwr0S0fG3V+mT+sOTjw26jLfMTsNDgMwmm9ZTwqRgEJ8LPPwq1alE
Yl/J4P/kANeRpLmb91eEe9QbEQOF9Xi83gRsf6SFA7z/C/PCutQqk1cn6CvCNj7b
RyyVcNK1ItknN+o59od3oBstzoi4+0DCWbI3PHgnXtNIDv4aJS/uSAce1chUT/Ua
lG8oL+2SPzTJ5hggH/Bl/3wBn0oUQAq0tQzgK68LeI4E2cuB78mkkdVsxJSHpD40
RP3Pr7TV8nfb735zlzSHqF3ZEDXA5KBHvnC8gFYJY71ccpRr7ZXM58vnTNXoGR15
WyUPPNgP6mHHX5kooACSXvf+63pRgTGJNZaW0ZevTekl1tLghz2vfJKqD5GwVgaS
SBgE3DLMb/ySsjPQkCXUk8EFn0u2eIg81Ti7tVGOZOHTcUi7cRK6P6ivaF9fhx4o
CO3mGcxAvtXDZdjDkZLtIYC9ifmpqzNrlXFgqxjTxFgSNKMsyZkIKIBMHI9+kB71
Ni6P0le3qq5V8dl/K2FTaJ8VuVQmGieeH66C/BHb7X7NDouz/1z3sZScIIFPzB3x
D8OaZFgvqNexvDMyqbsfjSSxmTEfeL3q/2LG0cwZR1sDoqPJcwUsea2KjCQ5TgFt
5oiPbwD73oH74Vy1u50H+5p8YIiIraiGRtiNOy+P7hATKRiY1g91RBiGFMee1KC+
u/pfMHFybZO4/cE/Iu3/cw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
aYqiCLGvKU3i1dF2vlUHbCyD6E5aPpwpoFS/32cb/Bq5T+LTs67fuxYuZgq/z4p7
Lpnk4g09gVeS4+KFl82QM2Qcp9UOsIMb+yE9+p40AERta2UopOLBhnNJE/7AitZZ
P+Q6hClM9j4mVEj+rVNlZvwHaoDTsE7S8xv3omkJT2egpAmVKcBNhOTbTOmAYVm4
30g7vqU7DKCzr4oZTM2txBnoECkeamYCaNkujL7cC0Wol831dYYr+yZbaofhGK2h
25vMmWvtlV2aD0dioAi7FzWAEWzPlu3QuWzTsJZCtLtXBll27KngpSQQdvzcZH+W
6uZhVYmowfZQhDc4k9Nxjw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8864 )
`pragma protect data_block
hhrJbcSk1CCQ3OJBYT3m3TOxXW8qBf8Ilmx68oGEcpkGNtN0eCKXoZP/sDYkKvDs
GyH2k66qrWNk5TCKrVQrDe1rG6Fa2Y6ZGoR9k84lxY8Z26XC/u3MS9IrsO3Pts49
8Zzf074jLmuH1KaqBdMZfBB485Oqc6XB9IPbPS4WKaFolURZaDTBI0vZaZFb4dDs
gBHv8fzuJU4XE8AgAmr5IESy4a+csnVYY6dXeTSpcv4bHd451/0AkkvtwuHBkwUW
JtneavQJAmat91d849J/ElWqovLt7j+XWj8Xk1MMOmNmrd3NubpsEbPeQ+ds9h3p
FXsbJumzuSq+h7+0J04IUQIx0C7LCrwD9kfFpznObnm8oOv3zVbRpUcKNw3tuc6v
9t4mDq9t1jFmeFy8xkA+S0BQuF1EAm0kw6eeIrs5ne87mJ/SoAXUUlNWSKJ5fzus
5HpmUftVmPdh8zvExn/plM56+Q78f339GJYvtViRxZFiLGXvSGPOObRmD7zlK952
NXWnMvUAx+m3Pl1MgAUeL9Rrf8ajr8Y+Q4/1TE2zbjok0X4OcNBg1i9VsDF7rVf4
mFebsI11iJMTWKDm+lNmhGrutc45itlKpjX9/bqx+LK/XXNxCr0odkq+GcgS2cBe
r+kmozmk3eUH0C/uPpZQN2p8WNWlHtIEccTHRyUE2bdw9oGoZ+kMudELTyU9yzVO
7Ii0e+6ULFvW+QErU7mTA3Qh3FzgpYknLQTB3ni3Hmi0uJHQIzDWNNknAYnv3nDg
lJ/qiPV61s/tdl4+28kNlaUmo5wdxbdlPQb1PoiFPKamUxX+01PsNvDpWlERm3Jn
IjzLDi3LVK/BVVufTDrLLLe5a/7EtS/6VvWct7XuqA6XlUfPYoDHxQkBBKIeTukR
azAOPhffbqtCkxUSGBhupU8cJWAnAhjQlwBI0bT5+C+cD1YbP8Nqu72pn72wcp7Y
gkmkVn00KaBVtuXezs3fEeKy6HJc17S9Na0fvHUpl1bHFyFEbLJy6VBL3YGeMB0U
KkVwXbxlSoc8gbi2011PyTnJtMtl/HegcFwVx0/BOfWD+mFRTxnkmiGrF8mQKxnt
QT0VEUbq9vRZRGkZ4oxBsZp7WBpRbouvPQJtHnjVanLzNhYr+qI+yrLXBqO8rUHE
xN9GJ5eGTOgqQIcz5Zp6FkPIwc+L41Ut2+LhqrW632khZC08fQtJGluwiBfKqrbM
a8HnDIMetgHdShjQMnLb6zItG2a7JP6VlwvU+1OeDmF4G6pdvou1OYl72GctU2NO
o1PF76k20z8zF61vtIWf8emNYXM0Om0aH7Br164hqwZ0bgOYiEkf3Ltk5OMHm9NW
MtslIQtILvLcHqUbWL4gUmUAkUI0NEaCRIBWUd5rWMGnPINh8pM1EWypCHcFUWNM
t01wjT2DZj6caRU2KFQ//jCR8gpv5zfwa0kt3+/CqjQsBG3UGs8lyTp/OYdnRZae
jhBJQ8hWhEAgrEF44HN2OMf6xD7ZGB2FnsGXnkDoW4A8TR8lLuCoKkei/NWzsgO4
H9GWNZ2hzwKyZL38FXgXfvelqVVR+78EPSYXVWYLs3t0Nve85j20vWHa0HgY3m7F
CdXEePUEdkfqtLB+8bEBBTMf6x/S4HRvdS0qcIeYYksVOHX0I46+LVHWS1H/l/YG
wwT/ccXJrcfGUWCaEcS6Db12Nn1PwHywfauySEouDRusr2phDfvKIen4hUuch/nr
uSIUhqnFoVxm/zMu2YNEREzXLwNTAXHWZST4q7AjzxOwL7nWjB7C5BXIR9ZdBGtv
nIFFIpQdyN3kgZkLKmWHiIJXzEF+eCX3q6EZ/4t6UVCXqUB9XYWHGKx8LV2w278w
cv3OrjXamcEqfx6JUsLxRUaI5noD8zl2lwf8km1IUo7TbqLrHou7kod7Hfz0G0/2
p1pEgM5XA5mIYLnAaR1+HhbARoAlb7IfAAK8tbaLwtxHgQohtBQaJluWCMlkFo3w
s2CdDYxXalRipfqdjptTx+m9p9v6kUSaHlQdcDIWWj+rRJXABtVSezthLOL+8+Fl
pHpU/DdgmLupwDx4huRdB/xC3sTjplvtwOwh6PfEDZuw2gerIWXUxZz7UUmwLcI/
+ckDb808vURJf32JgJnn+afawwXGiJlLhczTs7hRhpE+RHniEFRKQoRSKzPkCrrF
NobqPX9/T/iV1OUMFX/qxCrwkKqdswXrssn2WLEAb15C62M6s7wXEBq0pDVA8Nc+
zmOFPARDsGkFlS9Dkac5eNh80dwq+3w2Ae4dRqXNJZnAwNLpWHpiKNsTKSzt5RsW
l8OYBCP5wq9c69yqUkYAToMRN/cfAhZGsS0ttDAVFhHYeiQs7TAYnnGBDXuJ/OfZ
YYKzpHPtB9ECn0ihTxVrhc1YVxQrukz5c0DvLRTLYIqZ58dYGD94tE0wvDpSndqe
t9jfXc5EGor7ySaJ9qnLcaEIlpOdM8SI5YGeji1PBRrkLx97RKviF800ohZPRKRR
hjsDy6jRRWzp8x3efS4xH+NiZiz8HdHQIHvY9+aN8cOuXp8HaJZ4VCK90lrLrDqz
m+Mp36rWXGa7bodfHpcmCx7cfeMszvDcjuvH4Q+mx6IUziPTJpL9MY0Rhxk+0KGh
uBeqIeYKmZ0tOXmbp2ZU4Uw5r6Iix+WaPr+rPvNzo5WxlJeh5mXFQomstIWVTDYz
zBIL3mP/mb9gcTwTbvcTnbt37MVc8cIGadE4/eMNYbhPwcMXoH+yen0B2p5XV7w0
+s3Gny4AF6YfLSBAyBPmMMr6emU92Q1CJWMKXCsP59UQWGEhFPaHzjgE4a68hgSI
+eMZyfyUWK85dm7oCAyPRzHg+kKWsRYEcRNgZojaLo39BKwsAwo8NHafzvYUh3Aa
jqBpIQdy4Zqgz2s6TaPmQNCK0Kn4Ueg1hoO8PySBoj5x49FwTeWSic98lMU//2UH
QdamYe6hoEB/ZoYROnNH0/SZ6pDu7e5kknQFNWyqRSaf2MyCN9byLzETK3nJdaPI
SVISHPa6WD+yXHP+snDG3FG3q7kFcM4SmVeq3qMVsuYU1WBsxBHEHwhs+QSowKZw
HSsKK8BblXSGtYJ3+4DeKY8cDaWT6zJFuyBjeAylg7A1ae59rjhWQQj4o/qsysmK
VQZUB1m3Ua4MBAccGP4bWZfYxB3PHvHjMcORxYRL9S+hbYnlPZ/LrdtFADugSczX
DVfDqxbvQtPNIOxXW4BHIY+Bb/EOXyvPareJlY+5eXLMnTMJbQKTDMURzywKrRVb
XSRPTyFlH/THI2VGajTenNHVXipe2ZSLw0akMMUtnutFn2m6kOS88khm6GdG+bkC
Tz7YSHf2N/erik63mZLP1jau4qUSdlNI++TnlV85H+gr9SG7xqe0T42MjZ+ijnl/
yRbPpmle8+My3gV1rV0lhRSGYrMkK/bGSHGJbZadjOa/BGvR2AzvQ1FDR5MTfZ5h
Fr8ZCVxt9XOpmEhWi1xIp3I5w43OcLaAB2xviyrXqGfGEw4M2bfXXDnx1WN2GTJL
bsWCoerHi0koFSWzm5DJo+y02hvvR9Dd3rGbMjJXtNBNOr+own/zKmrbN+gl199V
k0UzqhPOZJYEUl7SI4yxon3s57gfdkoYkUVanPniripTicEmmFMeYgKwegT0rjmS
k/ck8ITPJY7jZROFZW70266H052FuZ+IHNoXTwtZF3YIu0TPrGyzwK4+8bSy0ok9
zgcTnjsYi3QY/szPvZVIxftcq7iijJkxKM2+4nfNstJQ7RE17TX7pLj9MBuL78Dw
7lgTuGu55c7p+ulFAcR1ST2lKKzYJ6oj2D0BND9auQaoYwevriImLtDYXOD3nUwU
/IwYibwLDJOVucQQfhvv/PIz2pwV3QyZieXJb6NHF4GpTxCPdNIGBlwxB3fzPpzP
yWu/NBSjy2EU5NDUO7jvij4NKXfN++Er/VZXw0JjpR9V1bHtwFxsg0siid0wM1bm
l9lx0Vn4J+HFTBmH7GH4ppp5VOiBiRg9FT0wszTrfdrsibZUSSgZOwDB+3v2Xjrb
k3WHdg6qusJrC90A3PZ/1t3VPV2OjOiE924pddyAQBemWhpJTnVYDmmUFF9b04NY
i3udlwUTdmu4RVy3W2oVPoffAv1LZC2vfweJsujcKslNh2tcOeeKeQ8Bv1FLn24t
Kz5mEH73fsY7kKF/5wRsf4AOb8IfKySrf5wiPXwXVsM/m3Y3BGbkls2t8MBE/A6z
m/ngs9jDgb/a51riiIUYJ+Z/8l9bjS2lVZOCKA+SrtqySfXEsBbN4+XrfUMEZVUJ
9hc+71SEJGhnisH04Sru664gkXWK8iOz7FwzcYuJxLbaDIKA9YrV+TSjEzIt9v54
rU1+e/yOn2j1oNdp/TqsNv3JYyVMqARzv8gnVCE20rkJ/tLdNGqml2JJhjub/LQb
Wehejc1yVRbIqDW5StMW9hSx75l3GiJUZkSDyP2fwg5G3gGRtR7dxvLAhjw/1b0K
7NSQDw03B69y433sZsKE+ROs1epOnEgIi6MJhevSMxfiheManXn6pGNuskN9b/gc
SatnD7d72oCd/vFnvZi+gj2MT7HivEdj72DBWD11nb0Us7UERK3KUv6MkYPOO7Qt
VlkdHARb/bzHSTSAwyUmQt8b+q1TSX1f1Bw9wFyQtpGftr2S4yYHE2WfgWEIuabw
llpra9PQ57/EXUDdayJ/t9Ums4glVmWLeKDIhSCwxgRysfqXJjqSK7eQUQnefr9j
HtvJRaquV3lxYcQZlRlFIUuS04bwT5Z3bK8qNR90aUQkx/RnFGyJmSMHSk7vuxdS
FoNd6Tjgg96hDgUjzJLKcFJqLeRB0g0/+hbWK8DPDuz2YfEpgJiCZKA9zEYyuIHA
KQZz3AcJ3r9K8C+gltJP3Dt6RZDg5f9VVYyGeAOY2/ItvaBbf+dP4QTj1q88G6oq
GZ7wYXkQ9xi7AOKBB8znzwaTOSC51WaY1wQns4bKoUtp83UaPOZWUc5r5eUXvY65
4fEGXemY5pFBLdgHN5Gtq7pXlS59ho66T6IE6uGifhaIpE5pSy703Gx/y8Mzs6zb
4KtZtabUGVe/MbvgIY5TWeWEnHv6QtO05vdVJDHvTskETC/uqFDuUSy7VlDN323Q
d/3SFhbOfX24utdbtWgGGbm71oCZJTm7AChwS/wg7W1COBSh1BXfAZQLtfUv4Gat
jJwnv6a2A59VY8k5zuUXZF1HgUldUnGBliiNHSa0w1BF7S87J/6Ytkiv2n+oSUwH
4rqbH1UdYizOo4cJQs6ohsKlBJIQHYfprMcDF82BdEBoTv2knzPPcXKwcsCRltwI
iexeSe5e67TXYTjCHNoXOGhX2zGPufcx8E7wrCPHP+lSf1dj+SpnApd/duk00opz
DFz+o7ynehiEQap3JnjniomRJoAtOP5gVs+Tcd+mhw9FjY3c6PcgG7ygPObaKFrW
G/Oukkp5TK7MFZR6LhIU4wKZHTgEHFOk47k1A8PFDhpVlDouMkoCDfQttPPCKQr/
/TIs/BZCT5Ll7cnOzRnOfU2q7Dq9+liHx7A4lsgIpaK6CMQ+pq2a6HMkmMhutGZB
E9I8B2Hs1TXxXwO3PSBoOxMa+oshulbHqrtgVtaeiySWkb/UAmPNNrR5wi7vcHN8
XSX9+G2FIa7mauPyP/iVgVbGSR5b/k1q0sJbA6Y52l28AY+tfiNPADdjB1BOQbQR
ohxI82rPwVG8NLtCx3awl4LxYjwaymtrX+a5f7rNA96lY0/BvK3virksrgr/Qyyn
vAk+7FSjzF7c51PX6GPDFubE65/2pWh8THO2uyIGQBMeGsjq1SHHJ90l9uYuzx8W
Zk12Bc2Yw9izz1VyH+BgqFawRZ4a4gNB6K11etuXnCg5/tyD/OVvSzKBTZXz/Qq+
jgU5EcAztOvs8xFFnYg5NpxUfSWWAf2C699DtHHkADYmt/944HJGF1s8NrT1nfdZ
p0RY45O2GpOFfLWMH0bf6z5aWLCaRtKX8oKWVnlbr9sp2LgVTE6DFt275J62FBDz
CqEfL8n8RP9JwIyNWzwpOvNdyaizwYz7h7hh+6XY8ktCvBcp3lVvQVahL+kQhr0D
PH8ImABE9c5kbExiFgxlCL1FlEl14ZWqGjne/sBK+TfoY7KsvA7IbC+31+gat46s
nVTf+cbBEODCsQeMigkzBzmGJJWWoxkbhNI+ucicDide+NxPNZKmIGJG0Tb4D1Vy
7BjjyFl9ZeXWtenswLV4SdAsSMJNrlYJto+VpxIAkXKizwBJpAaTOtdTjSlkcJnT
3uzc8jc1FOgiIG8x/uBxEuPhK0dpy9vckolnbb5VmOccJvuUujjMVnRqaHjkI14E
TZb1KaO8hFGF7REkcWibnHrC9k9EaKJQJ5ZzqHV9AqzAHE13/4htfQuBGtZ3/QGy
MJma5OkRZCGeehSCMiamywe2qf/AFrY6kPb5UT5BEp4WiozHgGFCHVkYufdGozQG
6Y2B79ymlWxGM60aduZ+gVtXEKLr6yiGFxslTReL6wNOb/2r+oq8LvOMsfl2YpVu
fPl9l0dZ1oTNg9RzuzpIWjBhAUp46JaC5fGjou4V7HIf5s5UzrOj+oHPShLkOKuu
MPLrD+6hfxy4KMZ2ttJMi0U4+QtiyLAcjio7V3xHRpEL2n/fuw9xlrHaDK6oAj1q
m1bunsePMKjxdVDCnQmjjGNCgyf9ufGbd6QiCEN5bVqyEp5f9xPWYtCfLtf3FPHl
s6XkyvO9Bzzk9AwdKsURsCPowy0KPQN2m1IfnnlkGsRSQeEmUhxbvvXsSfhd04kW
J2zLAzFpIsTzOaeOglvKXokXrTHFuAQcaT/ZWyfxN6boCbfWdF1zNWfFVXPO0ma5
3ebrnvhzl/jyKgbDRQvFq8w04GGHalhI0fMM8Ohkm2hiAOd9VoNQreQ9hooV7R1B
2H2PqjLQqJz5X90KoloDbdpYoTRg+o4JK6aHELgSuBRtlF7pYUr0SS41Qw/i3dGL
Q7+jgN6LKHhapd7RxA2GJqGaM7CeE75LnrLhhisL7sqqvOXH2Go35oHgF7txFtsT
ae2P/1rlHAb1TVzS80Rf0FBHwyd644bF7Ja8TfsSBRpvoSPcnALJS2scR15Cu4b5
fRyuZ+Yx4Xmh96aEteyIVEnpgKgDYCTahKLgqnxvHkekG0trJ1NwLhFS8B984gNm
8tA5IXAT1uoU41/xk0jbrQs473RdlZY3zJ+Ra+ueTpe9A/6Vu7q5MvuX7R2eKyXg
s3VQWvYZjbb/hi1/HYQELlHz3u3fo+m3+b+R8WOh9zrdtG1dNNucSDNMZ5F5GYl6
LWvw3AD4eQA5/KhI8N0VHvQu7HAafuYfcW8xwaOhm+aXS8o8pyvCLca7vXknxxiI
cPihhlZovZ3b4qB/U5FWad9bT/CIGQEWPE1M5oT0d7dgVSbLxs35Pol2zUUpcimn
I2HAgHHURTymS/UFJjWyHcnv02DUBwziZ6LplcARUPtbHjjF0vR9GN/HDs05juap
s2PkRrwe/p6XQtcdA63TlH1Z7Nqg98EbLTxV6m9/+Hko7duQVhKAofsMF83FWexk
QI+JKxjrCU/ZcZy0M2h+6klIhWZHURekrtxHrbNB7X8fNorY5NrdxboKRhmkNGVw
1YYiPxxJwGSNk769mbOnkWSRGVLTGBHUzzgjDW2krK1qC0Fiv/5oRs2IosQB0bEW
m+xhk0L+dB2FZcaYRfkMCHxgyKcF/RFxjmOHvyYCZD2IWy2juvmi3hXnihxmPMPG
2rD9a8TrXdUFeqfAzJINufIWCdP5qCo63QsyQhNmjpMi2LJD/FP4La8TZovNzceV
dL8LeXbdoxFZ729DrCsdW229jzlZuELj/ISHdT/kipnk9ac6pZRZc3WYyWlxO+wX
WQu3othpneoYH+Fb4PXQrB5MFoFAtOvF5YdXtQ+KqCRKhIrdIO0N4skuYO6V2o9+
P1oq7lMsSvoJb/vrHFQnT3r+/TYJ0onGJ+mPuWiPbL165tAbQd16F+yqL6b9qTCo
LlBClZMovRmUhdlslW/mbdiWY1WfsPItEf7geGwPLGAn/6DvFAENBjGtOdq7LwN9
BS6BKxljSXcE/eyhS/lBN3GlFtE4zA53N8WUd5UiWKbiMrfiPjS3IbnnVo0FO7/d
l9Zb/B2uR4nK61M6eSqnooqYw1tRyrH3HoSLqUg/vfVCznQQhE/e1CQk6gWleBRV
f4xQl6nf/DTrE5tTklkmw0eAfltPKuDit8IjOEQlD8JNJaro5WsabqAUlGrx/dUw
zBKFbS6MPfygepQC1P/mvac2k7IF8WGPjDOc24WYii/9mNNmq2H88ltVc99NRZ5y
VjGPYvPGJ4umXnLODOUAytYvrovEjrPtfKz21DRVMcCQOtJtLUnLWil6hNr7jYu0
6xkTBlddyjTkljTbvte5VXadGworait5+G8qVcLFVLrcVK/ZtKXwJgJL9spst2LU
9ZNPmnzPH2a3CEHSDw4zL7/3MkB+EowDLMx58SWHwT0LKSo5BvD9IBgjg1uIA9lt
VuLuN2ZhKqr7g5YKZqeC0eQYX+OTBQ1EIeBFTL2YveK91IskmYJtEDKrCCdgqUH2
5O3HhSy/mE0glfMGpXtKTlTpYa7gXaPf2jTH/1pbwF0OuP4gCv+LnC8iEBdIrV3G
bhQerOWKT6VsfgqdVrk8aGknE/yreH7InooW1OJ872C5AdDHhKlljsS1ocCaxzBf
PrlViUOt0EzNSbNpBpRRFf4KqpKu5mqTsu0qOagdIqObsL6LitZVson3m7Av4uQA
mep3S1l7kIAbcF2+k5UUyzBWjVHnqK09HG9IT7xA+CLbCIZhh4U9j6i7a5nbAcYz
4f5MzngrGJkh77Fe6EkrZJbSgjGmKV4ajsFatkmNwh9BmJG1tkQYz5tYDlviSVgP
OVMhERSiufyxLLBxxLKdKS76m4BZTziBmkPNImE/HKF32HAFp/y3g5zDHEJXZRwk
4rI8wH4TnbxELNDIk1EOeziY7X/Q6Lznc52hkaZeVKtVlE5E4lf/KjpCuq5tpFcK
qs3jp3a0Ymiqu7kFxFDUCprwwkzJX4SwJ0CHOmBGD5P1AaZ27KVynWnbDs1xf6wJ
99X5Y25PkecBFQ8yax6XHK7xz/LbfCM6NxZbeaPvA4zUBk0tcRpXgoOLMG4Yn2pY
Nq7eJIMi2f5lBuNTMBizl9juhpkxCQp7wAg9Z9l7F6OCrbenZ+8IUlXFNs8G/ECW
2o/8E+ok8xWWr7Tv3FK6Iy7xBiifcigZYC/rL/v4P5RsVGZFbp4cXxpKhWm3bWMF
Qjj4qy2WPUqQS3bdz1IEHMEWLVr2gDvinFJh9ydr/7PEtxhP1w6iQyu4TT08waa+
UGwW2ach3cgr+FPO+ze6GJqtP/QLHx6y/p0IUh8BUzoqLF4IfSCiIOGk8Cy0Ilxy
bfSuFec/3T9gI4TGY6WQImgXQkXsXFeXnKf+OdHB7PihZT+yuGpqVt6nHs8kWLlU
FH0Z2ZXxOIzzbSBVVU92Oi7BjcEDzlk9VgYfdhb7AoeIJ1TW/o8nDhhuS53QsMmY
mxsXeC5ewyCuBUB8vS8msfK7NmKRZcMxvisdGg4BkKQtsvlxDIlPEIJDwJ/LcBKn
lfXFqY1RlpuyKGqQC5oZrPKegQkQawLdIdpvZWIfbFSWHDiEUH6V7JIFCZZqABBY
qZwO58UdspnXM3i4N4cFwYQMKojCt3o23B+NjC9Rggs1ykE/4M/tRs7Ae+J307er
JHnhIa9ifxljlf1tWWwwTNoP1LpVzABYpsr12HpfXHtIPedgFnFtwt5zILRFzIuX
D3qUYG/YscfUmaBNi7djTFvgwNXaHIK/1Ri3LbAqLDoPEcFHIS7dxHYApXWjyAbW
7QNHe8UtEIPwb2qHbKUTChWXDDram65ZwF78loziHEt2LwHTovc+MuRKRiDJQk01
uAU7Aq3hIzKq1cJkxt8pdT2WV+x15IeUTBCnCiPmUePPBdUBknvCxE0YEdTiWII2
gcmh2OAdTlJP4zrj9kapoxsfnUmsaMRtTx7VAUwwbtQ17iW5HgX+EkGa3hCcOZds
l3tZVnI7KxQ4axHZFtMxUr1EZ7mxCXORmkhBD4sRmXBMBOGDCsc9oJkMX/lQP+Vb
8j1tMWjyLiR73jiIK4lI6lEuL1qyDYGBgjnMU2vKjnG8VQspMWxV/7t2BzewKuLm
dJsBJTi+e99W6hpt7VtL3sSquoawG1lc7USAKRz9sBMDIv6bUx5ppnuBPIj/gUfO
mVx7ih8Pfabv7sN1psMEI2Ik7IwaHhTaCAsv/SiDhEhKcmqmCVe4yDeAxz+8vw5M
noHltJwRifgjsYO1Iuo+WtgFFpnYmRR1v4OwSZW4EXbHfVceHQv2eg5x/BPrAvUB
RgTBNPsFoli9nq8h8E6Y5OzXJyQRiNwrIANHWCZbFenSl0MrAjBozBWHi6Le+c+U
2fZ9MeCX3sC3NrPt1wN8Gpa4C4KBbcloCCfwzzr06F7kmUrAsIbaqLnGgu1c8ONi
sZN1GphV71r6m5MWjpGO0BIncTdoUIiQgWH5I/w9qhXajEkGk2XrE4RivH9dQT2+
dwJEhQub9sBCZ+yv53fPRlCotzvkLtPjoGb2mBAyTxC8fgs5w5J/blOIIpdA6i7w
qEF2MLkyeyUgjAxxmhb2b4ecSpQmlWbWLs+Ms5WPI/bERksbeaDwXFxFOOAMeLwq
wwyb7s7kPrZJ5LVM4+6Mp6XNNLQapuFodtvfZHZQgARiMn3ae6cp/suJHcAakwNf
KkVFrpcI/f71SBRM/u1eAzEHxoGUUurlSwAb8MoPfFtXM27qftp5ghFy1JFcsnfa
srKox0B72FIuRAvymbK7JtnzuRwL+KpoOlhdkNnttKoZM2ENeXPrs3WZ5RuLcr4n
/jVTHSgluAnKsuedknNyrbHfelo3lPFB4y1sB9rJC+RZ5Z3r3ETOqc+1RtOmJFk3
BPPvL3d2Q+8MvToL12fF9+YH/UR/uf/5t6X0s04aXgDpUfnrqkD2WkVvYUPglqlT
xsDiQp5n7hVsD8DCVMAIBGBfsjqXSjmX2tymuvA3pD95qqcbyfTfXA1x+kdoIABp
a7gAGNkZ7RCNEUFBPtmKOQIpiDo8rz4x5qCqo0PZZDK5LI69tvtJBP/nwBL17OyI
fGg3CCsTYKcqakmSF8NBVMT1BB1kYtwTAUhLWZ1yUqTix0OEGbNjQBHSAHVrNSN2
XMNb06TdOB915fPSUlUn+on/PpF/NxyqkC1m0kkXSLN1/a8dnTteOjrHarx8bUJW
kChWu2dqPyeJUBCQxN1GBqzVs1kpEWT0hg1Ih0c4/UfgwHUICzOnECnwbduOZeJY
x8yBokVASWeZ32iuJ9JaIMVNwhxOT1ExaoBnx66gaId3Fa6i36PYyChY4uOYen4A
tZkT36KhEIp4uliufcDXp2N5H0dS5tYQ3lUqf6n38bvtnDTaUNVej7DQLC/M+MFw
7GIwb6lbGLkDZCc0WCHW6wCvp7MUmXPgS9OKHSIk5ewCN+AFzWSXT+xF6nCeriTp
C9hiTgmjFDPGDHCGKaho2hc0mNMphAfUOGae3tjpL0sIfGRkXQTOBfgJD5jIdXGa
vPL87a84mkWDa1KpxGPIIpj9I5A/o0W3JGGL5xSVNOWhF24ER6epllN5aX16vz+L
h/HaPYwPrBri2jnQsxA0kJiOn3CQmmtRRB+HYFgkFIp4B03P8eof6lCMx5PRn6EY
msePS63YdosHzgEkvbAEm00D7EomOBGAllgf0/JI5yCc6d2d+4S6Cq8sDroqbjcL
ZhmZ6+Abe9/6ZFdccMxjIlQ4SrQf4RMqLEcISfMogmk=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
T2dLOv3nEiQNpN3Y88w3qsTynlPKqV1nAUYrgep9ubSvFLnazJmG4Hzw9Xfk8c3y
e9nDjsp7IZA2OsSIx7R9qkhtnk8eTZIFtAFBF1ojyGM9oOZRMKWPXQ2bVqU8WOfM
BxfXIB9AcT5YH1mALNHvJv/AXe6NHalBDOpoDv4HdlEAER6Zx0gIvWQbp2qG2HCh
81Mckn9rPVa3hhqBCagKMlpedQQA9JSgRIsqd3Hfw286b6xVlmulUEaus1pDHs3n
0y2Y10Wda0buKBRDTfoP6mN8GNOYgbbvNMWh5kRnr84iw127xZH0syBgGLnQR0oD
ZVclub0RvIGNRqWDOSap0Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6272 )
`pragma protect data_block
ZZ+qsieP3vb61SIVtElvo03Xj2gwquWT4zoNcmuod+De3YbogaPVCKNazwbn9ghp
W4IB4KRw29rib12JmpPDQJKAmSOwe3TsIzixkVJEJ45mNwWCM/h106f9EMue3llP
mqA/KO+1MSIhC47wENq2B8ttMmylzgjztECkJvoiqQCFhkSzhFeeUpdiaRm43QBj
Z0SW1Mww7IEOae6mwcgwWPJSiJ5O8LUc8vvaOa1lF3QfVV5E4GeusEPUNYzzZahR
LqJAMlZOgTADL539hAoRLNaze0/QlDNSOJiZsADVDFVMhG7LJijPu2j2yXItTz8s
o8ltcK6TQeOfGhBHxzTDHfo63JzGiY6cGjkd/qqv61s5ToOXhLBAr9IhuEmzgTQW
OBYbz5kSN9jnW9X7+Xt36DYmOIP6RPlbEh4ZzNjptkVxw1v9r5/i+LMxjlRCSKH3
TuThbUFsfzdPC9hBzTFeLFWpnWxuHMZvr5WI5T+y0MJ76+t1cySCz0H9Y+rjO9iF
9sOpiMVBoCpV3k/4TqfXNXV71ksM6lhHGgqvfBBJrYXsanXZ3FMgKUTYqgTsK0L0
f5X0hcbQcsvpee2pTyfDrhuS2mU3NkhxGnvIsQXbVaSbVKhkGydBLh2nzLlnCNGg
cuDh/StMXwxupsZzt2Hj3+YJKE6X8eOsAeZPaVMN6MtVklb/y3Y3LznlP69LATqP
6clYHYv5cRpPmvVG6dm9v22lZgFT3Rpf5jQIzYby5LGNnjkCnEQBsEBl8dri2Qcp
3N0218i9wxmVxGx3mqLzfb0Z/AKDN/SvS9U6CV6xJnpPimn9T67EL3AdJopO2hXw
6QJHLaG6Gwe9XKMqJrC/eEU5ZGse8Qwm5Chq4jqjAzCfP+Uso/vtsDe1FkFmpz0m
Vphm3FzDMkU2LW5PNxI8qcdm3yFjv4/LwlZdTANIhWDUXS5vHAXqa3Niz1uyzrU2
76ss+tCCRvl1YY1X28RZyakhrzd4+Gc7MXcQpV3RcDynMhych33IZieWrDeIaw4u
GCFTf88tpbNWFmJ9XPkLstPDvyGdTu68JGlW4nQdrrJVCwb+pPpS05J62AF7rl5Q
TFCw+YCvblsYBNPeiw9oCDRZTSfe3Tsgp7O4UOq1LknShIs/u4bLdIllPbNfD0Kj
m+VCow8/Ln4rzlR9JeYBedAT+0GLETjOO3saf51zJlTrROBep8LCa/yxC5yv3/9a
NKTCwEtEPJzpH+hM7aAH4kQSVWgI/TG+rotDd018PZ4HrhFNmbEP3ewKWqSixMjT
PzgHmGWkNH6TKxd6+MR9HixYQAJL0BksaSCyQ6CvMr1cVN2wAdTE/3RHObjRs0U8
mdbix3rGCYMu3EyjWeVcF19oQeOjWKbtJGNBROVP43NL1Po/Szl5tm/DVkFYbshN
NrvU+fauA7DWrS3JHQGDOWd18moqWAtmK2lgSAwDjlbyh/ccDYm0Jo/1RcJEoi+L
GsanqieYn5UptXmPg27id6Rz1Z/SHQJ0hRP+c4ocQBuqwbYPl98S8lyPS5ih63WB
sqsTVdCiqaEwc31wvytZyzOy7gEwypuv8Re23w1oqVdMh5UKzWM6F6n2ZeYRiehJ
fV7ilRGSTQIOFB0MluWXS1aGhXfTlMiUdcGkvhjq3ZSimbot5HM2FPXzwvzdqtwO
RMcgSNcUVnriVnYs96bzWSrvYNHLlbm9KW4Ty1YmWOtduZJrhjPnCJOI5kX7Qw03
vxv26Ct7YLoX1cRbvxTGpXCLFY370Cnfgd4NrCFC33Pye9LTaZqwoztQqBsM7U3n
SHW+puactKPKApS5kc7RXlQKrbvj1r9+Avqny3naNrljU+SuOxNqc9J7672mbEFi
XLaTm33SBoyNvXY6exYQH2UFGa05alqH4u1LhvspvwAGCni3BOx0sDZ6TTMurp/L
i4/lauBRKLFE71PUedATDCQ6LOZzaqkGQp2zX/xjc/YeKMIpw74pqXDB4KxlQYQV
Uui5Jt3gqTpflxO42wXlA36pZ+ayKXsEF3zB4YiXkQxYFF1gecKMRW4adzmDj1Ip
TFnBLW4mIY4eis9aQnROUqZySd0hnSIQ1fomk47476r6usUQ2y9jVE3PKs4GocM4
G2nITWyAgHRhcl5Cz/ozFGJVYHZ0y6p/F4dy7v/m6is5CQcbKdZfxb5Nl21oQz79
3A6HGzIOE2qpL3hvxkvo5pn8whR5x4e0b4Udy0gX36kMdmYnoqHCtPkNI7VngEom
qRV2+FwBZKimLy6oQQfG+/WBugR4r6faiULre3rDBI7TQ54yCudrmakwJp06a/0p
HbPN7gnkR0Ktge8+mJaxd9OFuWJgx/Y456HGMKAtQ3FEzMUJmBGIVRWbN55Jhc1B
zXOkRf6nnjrF1tMFkWQ/Dk0o+wIGT/GNcK0UfX6TC4okMe69uYZ9eiyWwy2Y7uiq
2nPO10nXEdhIRyJcQThuOg49ke3/Zq3vteZHgDk+Nyf0MV3+N65zuB80GASACIps
QbsYpnu7NV4RSM+k48fUs3q95K5NU3sIgibNogAWGdHKR89UtVFBeDiEzat+lBaj
AYZyzmeb5dmiQbcnu84DHlqpfMx0lmcMoqggVMYeFOmQUDXjvQdtXfi3e2tn+1X8
C3XlSMp+CTl1MxOSZjToLIcbwcZ4bIRIK+U9lLSg3l97T0T7N2NAReeLLSpdIIO1
IlVhTHXoqS0MXbKL1tv4WJKc9ijFb8HiJoz4Rtg+uUqxjniJsj4X7XukGLONT2/y
ifRdY9L0srFsicTh78jnYeCKisth8TuFrif8km9eP2Mnn9fbe7NOvqXy9YO0vQiv
jlNvuYMGuQxKzMiPi2kjbRTD3eE+xLYl9KL09L1dNMEBXE3yUVG5YtKHLm/up6Cw
TCJRa3SlZNO+ogCR98liQPTOEXa7ZqnDhpLRHcj0M6UBGnapbxBsp67LPUeqcdkt
9LwrO3i9p8DiWtfw0wCioSbnWLew0+aLT1GPuemtbSR0Jn43vFloYtljgo0rWeSj
2na+Jd9TixlieiAk/MD7UQgYPIRsAGPNogqMFr3huqYRUtLjUsLQT75aJxDtJ3cL
cdOzzunYNwWeIhGvqAJJO9qX8TGBWFM3ddn4r0PuD7iYc5WKpebASBZ8as9KyrU6
le32PCzEN6VYGhCW455zSiGlNmiJMzt1qfnz8sRzPXc1B0tfmMAnMvkvvfGtJY0y
tvdmYBnC8yvHCkkJt/6rk7XuaZinUkNMYCaRsfyrmr0eWikL7lYYXrNwEiSRKlWs
llrCVHpbiRJADmyOic9HVUGsAisdik/hHmTle8MBsL4fqwp8dSRqKbnOzpaL5v6s
F2U5h7ZNqGtRSyEBg1FG/GJ03Tl74m6Xx2RdV6l3dY+o0u1f/H6KBZDq4Hp+FTTf
LSPkzC+52nL5mt2eJ/4blSpQOySg7AS/2065Bh9uG+WbXmNKw+zCAH9P02pNfaPr
CVwlQzfB0SFCCdA98k/Jur3s2J9Qn+a7lTvM+ZLXZz5GTVxPuHITGdurhInFfXJJ
BfxcGP9ZiMAGsw9yLkaOF4w68DD/cy8zHN+Zifu4/lHqqZf5p5Iv6cKBKqwxfXaE
zOPdlNhv4c+kNEGemzT0BFn84wRdbUNz8/ELr6v6sE6dI62vjJnRBdKwSZYP15GW
iGEkrIqw6pQOSglAzh7mguyFFWAKdImI9MayqqOJAr1yQKvSl3pK2xOTW4nUWJV6
wJUfTAM/lE1Xad0YylSrcwFm7e+vqbdFyT1kr5hNQtM4bG5kCX6lQ3WeF+MN04lj
EtsLZu1eHooVAnQpCU261m74YH8gT9tdXWdKwBRhyKQSs7d2+F+o1j/vgWOA75Oo
sXcdIzJmzdnA9HLYgNwA+Yqo6/Q35jjeNoKOk5Zmiq8hGIBIhI9kaV04whiRnIhS
u4isy+VciPQsLPHWoN56ZVdCDa6eJG3KSsRlliNTcgGv4JTKFC2RIqoCIylA31p5
JuD3P9wLAwVftxni1fCGEY4v9cLJaYTb+YORPp6A5kkEVbGXu8C8Krs+8RvH0g/l
EWb9aoWS8IOPEBr0hLI90/r3SZMfRzT7SN9jgQyR3vdTfcxARVioOQK3mDL0ff/X
Pb2rq9yrrnwprNxDZZ6s41wYiDdE3Ivu2rptZx8aYK4gvcewoF+s1nQT7i7bZZKj
HDDfUzRMV3U6qgjmDwNN0fwWEs4W3CB2yVaf+aZEtPnV5tW+IqrwoUG5erpEOhGl
do+o8SjxFE0MqHQzYskFS67Ko21CLIGVpzZmnXezn/LAeXzmKSunZ4x7fHrUGrG7
tZFgbr9CyADvge/9ZDnB0Feho+ZRmBEGcjryX2TxhGkgf9qMqJngjLJgkw+KqmUP
yymjm8bLKYRuSwbCa2jIzuNvCs7+ONc+FRjUiqY7W2UYe91RgiWuNHhxYkc5jsna
iFLVURrfbf1Wb9eq2PKx9Gt2rsM3sPfBjxyXRipguJnY7CPmCzm5fuph5gZcxQEI
63HLfMpZhRCHFEhNdvYSrKCU6K+znp9inGpKUzfivxLR0FI3LHjSkk7LfzTpeYD9
q/PMHm2S7dELOEFP+CKhFep6IBCbL0GszrOHRlavNZW09tI2UEI9Fa26HPiAR/jA
/LPe5P0vnHWqEJ927yAr1H+MrUc+jo3WbJbd0qwGQeCqbzdLMGat6t7TGCACjNO8
ZvUBLqwJVxM3vJum5BwfxHg5DqIlXUbKRuu8qZA+wzC6Zdcvv1KHEbyGMnr0R1jF
RvO6SpAKIWtXu6hGV6dmsn86LXR4iQqKgsn/thto5jPM9PbERNJ2A9jwPQFRpc64
DT4eldslYabk+2JmRdj3Q1fHwvZkpJILvq2xuQQDPLwlY4CmFmvZ5SDRnrmO5q+N
YVn62fMQDJF/a2f4MiU18EgTprbO4hZ/8Vbo9Z5EoVxX8Ix0u8u9UlTQCJfcsbIw
aR7NFdE2nU2iDtMPKio8ItlhuX8ATN/2ixKXbjqbE7p3qhly2/skse+UDkl7LP5x
hhU6gzBwbG6m2N3MhjWInm7ehniqhe3jbGuNLdxom33o3xJ8P6phuaq6DmKMfoiT
yoAzR0e3/VljRlthe90L7gXAoOq3EoRwT0bdshiTUcFWKk4dLZb372CiRFOlzRiX
bNV3c5AUbni1iJ+u4A+Vh2SBVAUl7ESRy329rKqNAqXbw6oTADS9bvnCaAdCmCDE
7gm43txQMUJzvtPCuuntEDbmeY9WaN2TrY1BHXHvgaO38zgoWgMffz95agDMTj2q
Rn/CUHXfYuXAZ23lrWEC0WaZLobG3dRNleFCR7DQtRuPd6CUf4KhywQLbpynvpXN
Ao4j6ZoXJJopsmMWRo0o4tpnr8771+NAGljVJAellQ39L8zboXiJud7+0/pySLyI
3WNbiCvtYLsj4gEn2J2xBJlMkIjN/k9DACrnkTeRTy4DQ8A/V2EjICtRgDL1rZQ2
96+Nxdy5LrWky+b2cVsJ+VRrSvqj2gLHx9KIYlXUOUBegdBp15GM8tnJ6gPmtmC0
FzVWJpCvpZ5rCJvZvp3xC+gI2D96w6sTwAnFd7krFYX2EZlsRhZP3H+oEjTFOroo
3tPb4FRf+uT4ya49XiDoTs1ayiLQUQ8iS+ujWozmnbsuHqmHTzgHgm1FriLNu7hS
KNPZdvTF/4nvOMIqate8LjNSBznEU3kpyB0C4w55ym81SDvf4XfEP9D7DBMb+lqD
WlzafITa6SOuOTjfr9NcpZIFL4Dhojvzh/8hTmBS5QzwFcAvF2a9+GjDGUW1YgHM
C7ZXcZSDK7Cs0nAOD8udxxk9sfS2D8PIe6dIRtJyIPWx7RUHwQgcjQWViW1zMP3/
ZcgeFaT/FpRN5Vsmo0O71+P9FBV8Xqu/cjQoD/9hdd26Wm17yzw4azo8pVXbWhdA
bQ+gey4qW7msfgVZJO8YWJQZw9GiLvRlOBGQZhpu+apuDws+cEH/DNaugOKjPeyk
/zPfyrbsFBvTedfLfKonrCZZGnXl2br9JvJYk2EaRiFg+3Id+t70+EwDUR7gTud5
xvaE8zKaIVgmATs6kdG8LZK0lJAAb2VfSHvG70TGJ2J1HbRyZaRYqrzd2Vh6x0IZ
v3AnXdScvlXL2tSjw14XSWQh8/xzFyb9JSSoUWb2EX2RUcH0MsKXtwAzEBB+K0eo
UwRW2K94YfDT8K162JINRPbVEWibXn72qVePcVm07JO/44R+i7Wh2VZRoj2jkP2B
uOAuqCr70Q6tPFv2AMVKDHDoMY+vJxSfRdyAWg8EHV2fP5TuCDHKhmh88Pw4/oHA
t8LZm5+U1C/SK6E0E8S0wbYh9NkKqkNoBIdEhGR61HkkmU3lx1pqb0xX9puWvEJe
3rtXpjECcxt+f2F3YJ0xvb+REVImd5iw2IZZxY5IkyUdEisBPFs6E2FxyGnw86mb
hJpvATq7vcf8saIqgjUCQm0AjfDkxPvxTCN+5MJVlrq5VWSlWU2V8G+IYEIJl7aP
Rh06Xgv9YphkhLCKRANsq/emTHHMshKLaIPWoe5VVSz7bDBzeN8B8fT8cfL9ICFw
pwDPGMwdy4zST1j1eYPWR6oOBLT7jzdYxHapT2/mhbd5Rtom8ZOxiurrYl/cU24J
23xoG97OAIVHOdeOuNUUMB7HEcAIAn7bvZfeiwNMStZchCxK8akWAASqwWNM/uol
+nAmJKTOcjKg+ZZDFam53CUP/NlMR5LN5O0UO4MNGJiqxw+BwsMMDTJyOxOsbK+l
3qt5ilmrb47/2AmYZvWJzmh0wxLlDBYZB5FNmFm/qzjS2cPb4/DqgyewYyQyt41d
I/7NIxDhfWn0iuevmgWtTCtp5oHgRavPf6fdH/XMEYsGp7rYVP2hG3slIW15iJ+l
jO3f99QGSFE0j0anDtC0XyvD49tfMs+r0MlDk8jHiuQJZE6xv0szPYydtmchbTtI
ESkS5KvQsR88z1bOpb0AipqmFCkCYBSS23JKgmmF3AO2jLYieCbYCHjx/Kb5u8Lk
2jZ3gViNHfEprViqydCt3yVpizf7umcVNbY8Qmz2l7yhvZ5h/R15ETyd3W8oZJyt
MMmtO1zz6cXjGJwt4Mc54lWRFEXTY4o/WAU9Zlr/LwEMpze99mAP5NyQ+hp0iiEK
YIf28QgL900oxHyQ8xGdkxhqxlh1VONDp/MfoszL/LerbeSdZm3c+Fxj2P+X/f3I
AqComCk+w75WSpENg8/5vZNLyPoQm4BdqeaHGJKG/MMukFdDEw2PdQswgaoya/wi
aD/8LPiZ6UgPF0dxyCrcypp8gQhEQPsJKq6AduPpoFuEK7PymD2Y21SgPqdBw4Zv
6wSZ4nT1qFx+cKNkl3XeIRjKwqjegRk6V1fBCFV0zgbsqr8kl7jI+21lXBqPUiA7
wT+Na15ysOOhLTmSm7FJYtiqkHuohC6Mn5od3Kdy8cYr96QkTZiUFTHapkpK74In
m9bf+XLe7NO+OJ1yf1pAU6aKB4zfyrKfW/5XmvmfDxJqV6QR0t59nsefjugXASHj
+eThOvONXwgGZsNHSw8rxEghMKYTxUYHJNiHF26M2totIoOckfhhIxO+kmfu9Nyv
+ytua7oVFJhMj/UoLlpgfN0gLk6KwB3RpLEC22DaCFU5mRmQLQRRFf8UrTJatUEO
3+S2uj1ASLfM3GtslSHVEEn5UCyqpTLFDXHdQadFqtRfrMWV9Tj0gJsqVmVIYg1o
A5SEpWGzls0Vlw3qhoApmE9Trpl3MTQbWwUpXD/KAdk63EfDFMU+1n/ZwHEXvpd2
0ZrfCGcAqXVZlcoIY9bnPAD6k1pW1Axf4LzhqdE4n3yXvu3K4U5tvJuxRoTNQtyD
XdR4UFlBxf9M61BXnFbQ7izfSFvetywxF1MNV/0R/sFbKn67eOhIm9zJxBPqZtlW
0KlJfUCiX7LYxrg3Nu2a8VAiLKLFSjuOmClg8ruTg4bzBw6gV9ci/sy4gdGB3EGJ
R9M9LJ85VUEOCN0AoOAFuc6HNdmrCyekZPOW/8Vd95/gGT1FNqL7o4Znodg7B/HB
WC/wVACIrwSiy4/V7JrUPoeLObxQ1RFM8Co33KGRA8Oyvw8e0VErZWRthSeDH13D
o208wSbxZSe2FHrOisxt6cSshBb8rUb5SHd4FxaKELyJwBvlw6+wxRT5eG60sK74
+1ELKIEQsfLuaykAgaOKiVVqWFTZ5i7Oipryjz2ldJ2XyXZA4mJNndLO+6GvEwLP
TePt5QTWomSFk++IMiv31S0vXJ4VNbdW8MYJO8qgs6ycZLjYHapq/FGBz2SgoGMp
Mc/OgkcWP0r789VfijN4Wm8bUTSydxqYJE9o5Cr3LsKlyTvr6YK1O6NThQjIIbti
WtxSWNuJdEZgx1ucnXNZWTIw840WlX4Y9klDavXxzgM=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
fG/Mqh0SErqG4ix2/q1Du+JuvpD0IFfmV3sXMuO87NhyoNiwl3hV8S9DAonVVWtS
uHHCOc3hDM0Q7AQlafzqQFA0AMcVlLCFJi6/eRnDn+nJcMyDxYRiiqCjqLjWjv/f
6VMGpZmSmll2F5yBpAXQUWOhkt4RehDgT+VTpm8JUUsB3yeXf9BbXYIWDgwG/YjR
8ntkFclm+3k+GcyhRVG1QrXC9gXBaDMu2hVzZAFtGNMm+0Mss6d9wWSzQtK/sC0a
cf5UDxRSdMG469spABww+6GSAFaRas4zQDEJq4mcFVN07KipH3stp0VppKGRu0/t
l4B+VPQ/GK/+IUd7tk7msQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5424 )
`pragma protect data_block
hB12R5PpjyS71FC7U9DWmLXMSlM7BgbE1EeFUYxTVBD4AU/r3z6CLGu77EN2Z0E2
pNny4qoHdr0q+c+80JkefHk+r/HtgI/jAYQ2T2c/jL4A2IPKiMJXPS1rbTgjYTQ4
5OUDXJld7W+hGFJLZOaSSXVaKx2TG6itZA870Z3LKO0uisFJ3G8g4lWDLO5ZyYWk
Ku7D4Z5B1IV8DetbX0up6N+aFY1QK+tEC4y8zqbcVvAtATX3QSABNPNfZffeDtMw
RIHyALLe4W2zd0FUDzx9ACaS8nUhR3bRegxmVuI4PxA5nLlAjAZRBLgKb+x2y9ib
UKVFT29xTdw7l9fLXT+ISfkmbqay4x3lg4k7bhJ3QuvLhy8itLyk0ly+ow5Sjl96
yWtQcqb4XaR9gTKWSP11snvvdxaoxlB6ahTlhwmoC5bMTx13BUGg1+O07u5MNFsi
GZhh2/WpynaJlbvNMf154Yq5jcc3PZuNPv1QW2BSXxCntYeaKG1Px5SixPIKhVPP
X6MnGVf1VP+3GV/s++1WlhbQsee9Pqlb6YKKfKZ4HzyoCDWmAk41dStcK3DtjrLF
PgBUc6gpc4D0LKk/nniNQDOka45bt2gr/Ha/i1Mk7QPBtGbSX1WpcyR7ZOIB50D7
oH3DYAOCOXMJBSxzpFwHtWx8dIkgFOxz2goCBNyD5xG/PLVDyw8agqbec5nCmYY2
/tXZGKbUK7tF+dhY25RyQYM3pjGVV0qAJZm6Xr5QYhWjPt7djN9X2q4jiHnR5yh0
9XePfLY+FOVeU64vbpDub9o8nese83l3FICd6x+kLJ08ukSuvcWhHMLoMY4H+x2p
1Czs0GY3PxWM5W7CVtB70L+U26l5FPwCHNpMxnSYoUuJOiEuYzlfQytpAuR8UlqB
0o32A15uGfW/iwxeSCq0Gw2FXaumXDjrLGzneejqC7P5GgVUx+023f9fh5gdwEbh
F8qO5JCvTO5N+a018lrI75EJ5DfW0yRLuArNOVBvy2p8djjdj/4l0Wy/0qrvCW6/
2My4OvWn6zOBSRAENKgFqcTp4f0H+cGqNc1AkpA1O+XuebjwMmH6ju2EK3DtrqJX
bt4hP+JRtp3366/KhfggKgY0+Hs2OjMRkpUsE/SunXGuUA7quUIIlP4PBQNnXqhK
XLLhGQ9+Vjp2t1GnH2BFEG5BMyakwukp77bi5b0XGAOc57sFtdIL81CRs9A3gy2Y
/bvMvKW7KiU6B9ARtVjIRDYPMO/aXozyeZvtgaFSaeWE49h81z5thDRR/LYy8Ykw
IF0SnrSvZosZ9Hp2Tpccdm8CB8EQsPsJyTXXFriKZw0R6q57cElM/jOpxdlvhHSp
9/+gEgNH/TL21sIzPl9IHiqgqqaxkACwtnkNZ3IoXngp8s7qVjzflbCIO2kY+PhL
zun4Gp52zPOM/b9fsXzFPyZHkWvnYPdyfahZPlp2KlEkJTHwohMoFDo3zN8ty4n/
KXAxAcarIm4aw2l96ncoy/yGKGCcckskX1h7o2x46iUSQ7ebqJyBb/8W1B9Xicm1
WuV6XqqUSSqJTGCNGnXuBe2DxBSHr+aF0cqj9HxAn1SNgJXMuBo6HmWwG7AArGpJ
ixVY60mn4hZPDSpfvdrGBbm/SWleoT+OplOGuqOAkCf5ZMza6Kj1vgssonxytp3O
jAGCOk0RAzgvRUvp38k2NpCsoDVuO2XIiUFqMFWq5DeGyZt27IznsnXFfk7zRv7E
XP9d1ojH74J6IcNVWFS/uT/vrCKCuWHTa0NDl87j/ocg4hg50BT5aZhJLcphKQ9j
Pbuni85/Fy7GAAWb9QH8d1FdTbMwOXiJY1Hs64AXhYMnsQru4AGyGl+6MauUQ90D
vhgPFihHHd5S8duxQ9xbhKTJES2L8vZkfn5Msp9bNLqnMI6rsmO/v8PaHLuEhZhR
iyiSi1gKDrco3jYKcj8wehbbAd4BQFDIFyiNlQjNPJIllo6gd3PqUoKQ5XeWVlYw
KRohBu/aUndEI9KnFqLQRYEyRivanmvRfYXsTaGRsHy3NtATE5c48VGkxKroURiL
pmhZZDkssh/INKt13xgRQxfL1ZABEazoVGu5+y/CtnpdHwCXr2RALGsz98SXeztT
31IS8ZB8nHg9Vu8nogAlVSW6STO829QgIydoMfeYAav9yjrAJVEX/d+RlSNcLqV8
eYoYowVBo6RCByg2V2Q3pIUXzWYNrs6CwuL5S5UN1TT3chhAOZOU45e29rEqIdIf
kMrKNrL/Uq4MWl1TYwd1iIlppbK47S1LuwohZuTshBmAsKxq6pcYBB99+LnGaFLq
2zHqIfZZmIWWGRd1kDAnNXhGYXvqPE3rUdsVWnboLpm4ZFRGl86PTkUNIZcmbDqa
Ed/EAcnEafHQdyporHe7pUI+o8DBFAQzXvDLUHq8N/XzwWhwrlSokTfkcp5D6pw3
BHVDTnrxku/Qw9AjvKyFTRkrNY+p5b28bQ/5xobnp8t60NVSI7PVBv9Ku80JLv9Z
OlCFaEfZMEYyO6tjz1NrmWPznVDDwp3uSRKclQWT/Q4TyY13x0CrdAtWr2qTfga8
z/ZcBk6YI799HBhbouKQMHwacgSed9OHwCFNSyqbIlpEaV1WpyjGZx8qArtsydNE
4gUeWin8BnjKbd00yU13JSqhehdb5k4lkWcOplE0DysJtUitw/c1DPcRvIHCh3i5
oq+8X29RoQNqOyR5PTEL/5rPTVdpnRrxcvrskcPI7wxrsSKLHng0Lt5I44LL4ksU
H9NDttrtvvQcMulEO82Ikv4GqvHYrGBMUr/9f7Htqd40DaCVDi0flNGX988FYnV/
D4PFhOSMhjnmvWDAhoLzfkUdAFs422TB6Y11eG8ouet3Z2CCJdeB9LlhzFhPgFUR
gFYRna/33sOH9KLhJPrx1tfMWQcC7BB7/6sbbsZtDmCuNZ+2lyINpnmRtfWfyuIo
nE9j9LxY0NAFSYzYMKWV6gUUsV0cpu5sVyp9yYJtHnG35E46e174NJq+DQddDKf7
yccey2cZumj3d/tN99DQOQiqkC2PfWKbWXfB7mnNlaJ8+v0Df4SBIghlUwpAb7Ob
q9BiXyfqctQJNKWFcKFlGRYv0mN4K9j+R6vE7FpANm/bVkSM+RAixR5py29R7bD8
MxRdvXr0G1xh1a17a98oudHnKsvA1HLdCVS/zd5XE1HDrSTbTKLEsjy2Ecz6wVcX
KXQW4Gas96EcNED5IIoL/REMFGeSlcjTxI5xo+7hsMMjZRQaz/gKnAEhTj9cPuGJ
jO+35sdhIQw0tC9U0z57iQJ8d7n0F7zJlkoF5BqcIOnCz+k411FhoNH8Mxh6V+2i
f9kLvilq87suygvT5EPLQXhsIIEJZZ4FLLiDqnvQGqeeS6PxYhJdHYx4He5zHBnf
INdLaUPrjG/oX1OGJsNhkcDlXEQO7G6mt3LziDi6N5eoOThgHCMO8BLJLOmMwQKn
nYKVoALcYEVREXUobXahnMp1IrN23iQBeyr8/Pc1cO4kgkT4gmmp6LgT9FIDuiTN
YXVTJ6+PtPY25EgQgPQQT25wOKPlSwYF/oTdHMQ5fdbOtxRM0ymEfBT3FVQdcD0a
WF03bDuBHqWnnUArpn5CVElsq2+zkoiVmh+F7RyutAjgDNEGd2gWWToroDse9z5H
FShoMVsoogVC3Hq4F1fR99T4TsP/Zi0CpcJ14p4MvbXN7yev6SAMaqoXbHXdfagQ
hJh7ypPuuizfJkzhWH3xQSftXlIwhrNDY1OVe2xk0Vf/RfDjf4Y2pZchF5687g5D
85jv2eWRCJgLtKXNkwNTqyQ3fIbgwNgdIxEpKz7avQrUARtMVpYEhhM8aImurtEH
ovXytXVxDnasNRpiqqco9nxkwDSgPd3T9BpXMAewpHfI2o8tkmE5g8gY4cCYfDaJ
NfDbgGgwiQAnXP5kG+1Q8FUOozkZ3oYzswgLb5uhCDYiVvq1TN0WzZG/TnungJE7
CtLkRESb3qYB5soEzm/+B11Zu7sBIzI24jTcoboHO7EpqWaD1R/m0E+EfCVAcTLC
St5GdAYqkzieZe+5krOoe8Gu8vCtl9D48KyMx7Lhpk1iQJSN8kmYbL4Wv7mkrXJ0
VCDBoPR0xl74MyFUDaZ5Fvh0n3I4bYLccD6eFsFca1TrhwvonAg+xBhpRhAYQiEI
kXHXUSs+WWwgy1nivx73TWy6iz2vdXU9tBW3ZYCSo7XNzh2TCEFEqSV1JhZCBo3n
cvR51WQzRbOEcNcpJ5fti7cnXa/XxuYRMQCHilRx58wBK298Cbgshu+QOOfAPByF
jVKsk5YMXRKtJv2Hrk3/CBTb+kw5vbU8u3UGBGMi4h5WFDbjC1CuA+kfhKMQES0Y
FXccg+KN/gBo4l1IIUbPzu9PuVtFtLQRdh2udBaBY/phZVg56zSBOfeFimYBDlPg
bBQVird8Byxxrgiqk/e08jOZP/53pEP8QzTPJLm8XA5Wz2cVaMrHmC/zQK/qV+X2
zGPYtqgRg/SSKGH7H2bd3KE5UxrT5BEuGQZbyjTu/S5WzVeJ3X2fALL9EUO6r/Or
gc2fneb2KVCFvcKjgNPkqNk5v+q0t7xlHRZfz+XOniKKvhXWRmLWqhv6hWPx8B4f
ERkkPI2Kt5TkPI2vy6Y3ttnxIAzYha/BUkR08bKjkTbilT/sQx9YPc/2bIz9cvnl
0MdhSS6XC9z2+kEwLWgIGhIWHt/3bfQ7UeGWVEadRJBMWDEBq4CYD2/8EbmC1rqy
fPcDhMFjkegwULdZPfu+YO3f10rHE5OtSGWwJtkek2eeavAyRC+25LkWRz+t+VS7
rrlMZQae4k0ro8da3KEOSsg0HLjt6HhbEIVtFbAzcDC0XBxgPEUbCZ4KnX74Qqbr
8SzyPnAVJ7AV1N80xeBbyes/zRL2phQ3sgp2UM6jfnGtPXLl8LEe/Juga4ge45Jy
+RllmT1xh9eEasUAOxZol9CG0g+C2YmnHkjX6Ego+H/V4kVRWrFUK+WJAAf3bVu+
2k2vF12su6daEuSHLguUEeLQLlnCFkKrQ2sWqkQ4GooaaM0SsxNSJSDfkoX5Krgk
jq5b+SR1nVXCvLXiAziD3sSHrg15VWqdBuzIHONowzYKw6NX8JnFcq1KH1Tvu/sw
IrdNrXmJv9sIl8xiQcBORLW1tNhzxyVZdpiRkAj+HDb0wne1EiKU+jAFxW4GhMTS
ZQ0qSZH6zFwa2n374uM/4l7w6vV5QRmHblBBpP1q8oaq7Pcy8LKTjRI55PRyTs6T
Y2dspLKGFjXZHqY4JIbwIVvYShcH8Pxo33XYV3aC9ztEEjtf15R1ZQX2eBRc+Mx6
yZ/xAX4vcaoEfS7TDogp+XXawb7IWhRvxx6gLTgtt5TzJf+xtI7QssDrZ2Dak2iH
f8gTVacbceLt36Byqjz/rz8ckWqimTN10ooGvLTxVPddeLmsNojRYUDFzDNolAt5
/jwRexkDkYT7O7F++qTqaBPOfBK4vNpI2CBdPA+Zfo3f259SR0sMG9DD/+hlWNY/
HUF+LilPEN5sWJovJf6wSdR15yVJ4MVdBPf9m0YJbJyj3EkJS6SXTbGLhdDgKVQC
9D0XsILeWEUk3u1q41RoIXA/5lSsGjYFjJQvpfs8mOyIkdgnAGpstHShHUw36iDH
0aldzCYanEt3BLCtR1ZPTmi+DOtopFpX6slp2XMcZWFc0DSl24wSIizSp8LykkRN
jMqSsm406L7djA2uI4PgOpNn89VXqsmMsMpW5GhLjOUAbf6RY34ZYnArhQX5GoxB
1CfFCirXRCMRaxKGoX6lOwMyuLpsHHOVkbtNEJ2+hVDAcTl42+70RSS2dJSZaYTw
7gNKBnTcybK4WLIzr/DZbEWw7w1ysc6TnqNHDY6fPvPWYbUtYSiksrQpsKt5PAwm
GVgyUz7SxNzLl6F/4fXvszqx2TpTQ9yGu2YoFIi/07v8WO49bJLV223eeARQ5IyA
2o5E0pi4Haihe6iwfZyTRz5xTIq9KDeiXbGbPnPpjLzNOWsbIj4vs4efTtAaBmNJ
E9w2fF07Q8KCWCMxxybmCcSWARf43+hgGEorY/ArybdZJtC6HxeRbR2QwKCpcWyA
2/TSMgnRD4vTSSYXgRkWvqmmfh9WzMXuRruzPW/b9d+F/yxfN29QpSgGIupRNjyg
wYjCGDgtcRCnSU8bfCwaQtpCoqo/b3B9Z/nnWX5DwvlP5JOepWNLT2vF5Uvj+cs1
wLR92P2Gh84/CWFnV05YJFDy9OCOt49t89bd3iy8Tx90YlXPa+7WgK+ZYIwBtOi2
/pj1nnR+bkcXFCpzo/q/KVI9Fc6itxC0r1CUCnOhoQVeUWgC/2J1jJMqhAwFFxxz
+rtGbQ01ArjtbIrzBXs82qKU/QP6EzzeZsOSLgpWSuNkDQ/6J7tmEucZszxHPacL
oPnwQ96U44XlnEQiCVgP3LX/qENCr/k3+B3N1N3GdYnezdS1CQSEK0Rtoh7s8Oyk
rCke0OeuJfZgguvp+4NxVv4zybv3WdFg8mFtX88ZIA02Kr/qU4lL9G3Pfa/QjPIf
5ty6JyfC/XLKI1Mq7GLdUN0mvhSeoiVLuaMPBcenhwwPQKqpHlydY9oH1G1Ia2qc
FFn5uYYWwoPbhRl7pGQ311i3cFk2NRe/iRJznCklVqvZdLaEIGbzRYymHvMWTI0Z
E5YIJS0jD+LzRxtYPvNuT6LW0dkxT16X26ci+SuEMdtREKA2VCytt0yCouhMy2Al
G1a4wYwMmoYO3lvyeFJrbJ0XTDAufAJ3qW/EytJlKOs16JL53RnNeZ1ImaVTeDtr
k8EXYIyHMvDL+dTpgQWC9k4ZZ2SrIDz/kIU6WZYfzbq3JAqm2gHOHPWQNMWCJr3R
vDzxC8X+u8cjqdxnEpHGmvfnr6s3dFu2OjzYXkaprDU9R6yNF2YfKLRfE034CEec
BSy+DgtjoJjqMvKR35ij/RubwlG7LMf/foGRxUdu2J1W4qF3AO6Bytc6orYuf/lO
lN0bS9+Ev7f/Z4MfCEHYLASRCzjdsbCxUWeljmrPyUwNDj0R5CtiWr1cJ5iRlCaf
8kAzI4iGNyUSJ1FRCfX+YD1fIIoSqUcFWGRxzXA/fatFdLKpmMK9ENYzaGK7X+Ty
f0l/H+N+Jw+QFY0/WrLgYj9cFWYQovN/GkcIMVw1xLAIecZolMwBXmrXmbxGHVZM
EEPB0C34FOSEW3AB8U31DPGbpiE8uy7S6e/3htVBOYKB1YutnbcHueIVx4o8aO9Z
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bQRQi0yWnkP8pHk18Q/8IUWPQ5I7sqCwbwyqNtESNltOVyWNzjRr0ZYPu5a5sJ3r
80oM1Vi2Sg8BnTVa7mqyS2lghqavHbW+V8LyzdgWtEb67nmOlEiLAz9TIq6oJiAr
5I91Qmyf3biL5Kt0OmXEXcD39SXaAYv1vQHYP5RLbhXoGOMbonevFp8HeC18EN03
e9M8CLX2eVpIWai0mSd3Z6JyS1mcAtC8qnmAg5TSBEcI7QxHmsfKDFghafms/8Ui
ZaorSnKGLsTunfPDeSXoCuCmzkCNP7a7pn42oLXiFL6YtEb7NHdNrW/S8PGz+ZTU
absrQB++sBsLdxZkfPKsGA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5664 )
`pragma protect data_block
cLcZ2lirDfpYap7b2pmtfCmc3iskMWu8dlJu86CuYTcsvl0AuAZlniI+lu4nLbvu
5SIcw5446zaJ8fPEJwfeBEtpRKdfd3wtkbNcI7CtO82foqlCz61p73d7/YIo9wi/
UZv34sHomQfdEWg+mo5PTzzKhX8utoR3f5Vb7UDQmyQIz623EIjiaC8dWIcqT+9W
NF4NEQy2i6ZUzGoi3RRngdGO6NnwQWRm2lf0Rn2cU505dg7sAOamGjok26zrLNBG
GQ6vVB4iKDedUSW16z2gYC7O8ON7qDHCpUubiQujXvEr3jpnM5QXtppdw8S83DJr
+T4w0s4yZAXoLPz4L6MZkDUj7q3AVDKeGW+VxmO4CXbFTZYkPgjWK5jSQCQoRDk7
oDEKcqj4Ej19hA+vZ1G3DuQUKPWmbRNVsVI53XCmPq/Gv46V7Wdkx410cJdOd2xH
48sFBNo/VfEDfOQFH3GrR5ZXY/8VbYUkmfONuIPVRJCK+sl4nPraSNRa2Iuya6n8
PKa5AD5pq1My46lKsMlwGV6DGOBkB1n4KfD5TX0MOMIzANSHoNh2qm/GjTIz677M
vm5daC+3DXW4okUWKiEwJ61Cv64vYPyhgL/vLB3ufs5mn9+ZujK9iDo6d14EPqQ/
t4NeZnHjAzYKPhnwS3nGkOQkRqYfTwUx++Kq22XO7jeWN2lKbBOn/eGhPw4Zjdiz
asrBLas23FFXd6DZ7xPJzmBGRxR5JnCV1Jp2mx2gi0fm8lr6B9Yr+thPvKph0OC9
Cb7Opj2zd210cZJxpyrQkvyY0zFQby+95GrUznehHfIm8j2VBVknyL9Oy/0wLSth
vW4fNqg2QmIjy3L6VkfnqRRvXZxZN7Dc2gOeX3MJf4DM2GfsU3s93F1b7t8uTHVD
/0z1atpCOltd8jNp+EZqZ+hcLBR5LydPjVXJeeK5dq5rIZQb2MuanJIH9gfmEPKf
OIrSsbytLrvKfhOv9WvTbt1APn+alfCzeFnm2GR1e8ZhgN1rYB5dVGPcyhFfc4VZ
1B41qtxOjG0bdsvhDZUVGLetGWY8nx0eQbU009N/F4H8xxcMi+1QAYd/H3prSRe4
nmrzUiosLiLz7USpJJsOFFrjE+CGN2zMsq77qiUpoMKgnS4nMl6PasKO0/KN82ZQ
tzYJjElbs2T1UZsfZZUaUnQl5iU/3xm2JvpcoFzW4maPcKr8NXyWFZTL4BY2hz1R
nj9CEmEB98CmbxX2Q24Gg8ERwYn/CnGqh7emh+dsyERnebQ/auib5Jn0h0Hy22Rd
+aoe4ENy3EMUvHbrwm9+gXJZOJ8rJmmICZtXyNmyTDITOeUwP8FMBk/N4CS/gpx4
emkacqxAV5IQskA98miRwT+zC8cU5aa5SYUD+Adc7pCgnqy9yBYkrJDPTJJqESxM
bcaVLEOmj5VSeGQS/IVPyf5G/vGJ6diyKwhyxNxyttgNJn96vB7vlpg2gOJo36w0
PGEXKl81WJBs/D6ATr09MYORZs9JLSIyLEZHxPYGEMmhCqAPcBTuNar1ffJD6u4K
8CRWREoSREL1fQM7n7PHnPgECsO5jfnXbNzNsn+Rh8wWFVoIR9WR+InkkNQlgKFu
6HDdoWkXY5JFvtkzhKqfy1dPaZjd1opaUL1qy5ftvHe2KEttJPFFUR6zxKvg4ugi
1k6i6r/S4hzG1xpz6HqWYvjP5Jkn2k9PUWXEHO4OMUErkH56CWUNfVFG6OOWzzFQ
ZPXM42N/J1/tYW/xSMNmz9hwNnAy1u6sLVfNGwi2Z0b2vFOGTpNmhVzgSnpZTvF3
DnCIAlW0jt/ITD92HfeY0qXXgPE6IVSJPAwDwdj1Z6vWY1PXWaAuEv0G7oo2x/tm
rzueMEBo3t652l1pN89uZOplOwntUvOu4G5T6k8azNZ27IDNB6rK3lXaibumfyY2
qaUmWEJP9N9q9ru8nL6kjBNYCtY45e+uQMQDqA+KVva8z+m+UwwOu9Z4iTQlgSR2
tjUasMERUh4pf5brCrw7SS5fzraCBZuRacUGPX+1Ce4DTnfk6VxDKvJ+Fg29n+6B
+cnHt4cfJOTdqAdaCETeM0zXWCdMSO3XFeqOZVMcCjN0NBtCJdsCSucA/Wd2sDeF
FYVo4ZcX/1QBCyaJGTK0anT20YbyIhj3Dy/1BfBiVYNg3aGXLbXx8eRoVHwtEsSF
g+bhW6TO0XSlfEwbsFlja5XAuLsyEmM9WofvJn31NFef0oO/qp8ICZxcjtZrDA0B
QOZNpop9Boj4gfDTOsi5dCNlbuZ4s6TjnZJH7CmxX6syIcHwUTTC54WgjvMQCoZp
hFZg5Oz+mNOMXG/DXtHXgumqZ0HaZqydXQNCfUp7A8nUecBfDEQPB/pzwv5s96aQ
qhIBzaE03xM6EZfqfv0GSmT4zytGfeZgxBuPRBRp3+0zRxxkivz2/6Btmr4mMvVw
p3u8Z2rqkJ9ffdtOaopGOHSo9+cvINuCja+pI+59w15LuTcekR7WTeioSwUOl2Pk
HC/n6vg1xpG/2wj4OG9Ji/ugsgMGyyz++Y+9r+0SXyY+wgA26Bs20wT2pDQVL32b
CgT5WNeWpwRHiG1M1Ag0KgbgiMGLV+jpzZMz4nOzkmeE/Q8NNw4PHvkNaNDc4DXL
2U0tQrbfqGKBgCwocroG9EviDRvHp4ZrJdHUSR9HoD3cHPnVWS1BF5I/59RpRw8l
4UpzNzpchE5xYzN8tvh5SV0/xL3QIovY/Uq/+oQFxdv+OxcfFEi2MOdYQHhCJr5n
PKyjCXuURR9TRFf3VpvTKGjZKCP2+hn89yjt0Oz0NURwjjBjf6sLYJaOK9ys26cq
0i6jWpJNlGHQFyP1mbYRZNWyjEs3zuLz9EvffhRo++FdSUfmgOfAJ83icrIXpdfm
EqpdmY6qxhZz7zYgGEdUqUjvLnieWH85En3kurMAtxIMAA82/lw7db77sN/DrOHq
QMuU6rRs6l3bPV3mAbf2uLe4rBfIebnOChonieUhwKzbJZkjQjZOlG4E+H/4YG6S
/pK3fUzoHZuvDYDr+Qn29t+TnrqdkFMPmWO9h7wqpXCbt1LYJvIlyVFEPBxuAH5M
mLenL671LKi1a2mu3ZgOQPtyoAnTdUVbgoy8077w7goUSx/zhZyyv07GMe4OQcO+
Iq9BaBg6E9szoCaOE+pW68c969CXp+q9gBNhjvNLuGcJNYsJm8rG+Jk+BtJEYmSq
QPEENa+y1UiDIUILwEjNtE5Sx4x5Sc6UQV8AHO5dGaxe9RyL5MkBwjjiPbNtOJee
BrJZdvnKjrp7t2/jMayptG9glyVNyVdHZp/hG7O1WT1kkOT4+A28wy6dQqFTKYav
2t+7YhqlbXiqJKiwLFDxsCeRHMtqMKjuNcNvc+D3KXSYPnK/05ymttMi4IkBA2ly
gWZlmJWn8OD0mkpW202hNNoznjXthjyq3jlRtDalkBPZw5uoyhE6iNRpW6lJYNAz
C80KKdPzi01agdlFu45GIbx0bphU9qj8LRtLZAXxk2HvNuOdEjrNNxl5X1w22Dol
zmjDbuEKx/XDItcIkK/lBVrLiwxaeHVeiUamPQ1xFu/gynLbO/Uek2pxs8mAQF5r
V54ZiEc49z0tJyx9YzInI4raks6wgQPu7N4dwoBwPcB7mOFpLHREkremeluWllTV
zQBoYbULrLhoiHqGAYxWtnY7alt7XSeeUcPgi8mW3qvuFgWmUfcrNVCXGemleKMh
Gy+3Rai1APcW7s13OASPpz/irHPKhNsZPsFAtW6fsYaq2QuT+uYq/QyjJKMFVi7A
srr7rovH9SdLpKQ48RmdSW+WPfol5evTD9ZyL4tE/L6OQyNJB1pG0WL0P9Vy/JeQ
giDi1VVfB1lxKMGk6AMTRCt8edwi/s6i0um356ZTSJSQ5kELbS90TmHGYiQy+UGf
JfnaTnvuhvCr7v1LN5V4Na82lr4bC/M5gjMJ339c3c517RfkKp52va4zKJcswaE1
ZfVoHEf2isE6HuKpJivDLm6Ghg9ItVg4jN45v56zn2PQbWXgp81UTwoHq8SEbC8m
VyQLV6PiMg9CG7ervL4jVbAmMhXM+8T/kB/29XmhSX38iq0AVRDur/qsmtVPANKJ
1YFlvSuaIbjv3vhqKzTFxE03mg4B/D9KnsyidEDdt2zdzjjTADNUKUDgdcYZsfpk
7ry3V9UTb7KiRDpDYvvANA+WpRprMNd/GsaOuv06sPCV+j1IG+1itwEfsKEut90P
jjcENZCd4Mkf8HYTlLKXxTkoW+Nm4JX01u0hLAmWnmAdEKzkeYylpntGP9VYNQ8p
MFXXkVIo/IiKoYWCiJS4ROhhyjg17LEUZAavte5EFw3LRVRa/oL011kJrSWTrxE3
EsSjMES4ol6/Y2goEKWTfc5KSp42YuNrZUb9FE9dLBkjUHzbuwL+yFJQNEZXzmWk
5Z9LJ9FyLgvYcelDdlalpntQfJa/nvx+FxZE4qXilWjc0mwnNjmNDMTGgHmzSeJl
b6Qc0AeAapIkfYa/vIcofYP+stz93P0LoT/sUPtCnqtsV9OjqQsN/z0Wh3Rfs7w7
tablKMqRaGDRs3VkBfb6RrMFTikcVCE2L4R9+QEO2rYon3zmARBPWAs58YKBot4A
APBd0F25l331Ep0ZYVK+3Bsxcp/8h39MPIw0vbtIVhcwU0P3rPDUQg6OLCe3bila
rXwQIqROdBc+7fUQwGwvJBmxe5lPUH6Vt2MdOVH9CISWldIybTouujex8Yi6qvC7
SsUnPQGGuDLVdn+Kj2QfQg5neIB2pBWubEWitqRzRXaHugmdeQ/iq1WoWXFCDRrY
srLcGvaqBtM4BfILZHL/OZ39h63pLy3sPUYHs7Fd9wLJbrV8xhakC9vzl1huG0CU
GUJBMh6Vp7vanP+iRsuGgPRc/7FnZb1m2tLmBcdOcxgeIUEN8AaXAPv14pQ+YKsa
4XZelBuDu82ufktDAqIrdB8uhmemEQ23oyJF/3YxqExxVPoZk9dnc7teLWGf+X5h
lnvbxwm3tiamtvX2g76bSoaMfGn1m/O1s0tzRYAeNjbSRGKf/DSVBJsAFtxPgUdr
9IvaGfdBjioTZktqcSSn8VKWxw1fV8v/6n5LpMGJ3mmJpliQ0jMa6aJRhEj0e+ai
zKsR+VrhFMbukalNosVnFSijS3AnCGUlEcom97pwCj8F9h7U0AJqtLjl+ROoMcCr
0xyTc6IR8tySdQ4fIIKbwpxqAzAEtvr2QJCkCyWLEdbYtW7JcCBsXiBhqAXmFW0y
t/cQ7ZJcbQlQEDGpTU0Lr75vRBMQIWLVKCzO4ad2J/1jNjtI7h395VnBMMdEa5sJ
6V+6XudTA3Zg3DUzU/EzB5R2lSIDmC4y1qZK2EkimTOXV5yLdHBg5DKKHQv+8xQX
vs7bYgjSTws62HfGLBSYJC3F/SwWzDKPBxBZxYYl8xhn6QtWOmh6LCTvWf7hI+lf
Bkf8MZMVv6rZIgVIoxosJUgVs+3K102WED6LyMHlpLyH7JvkTlgnc4QwYtmJnkRW
/hNNoTjpQrV0pvualgTNRK90lEXRPL6qN2kkW4z/8Xg5504pJmBm1FxrBGsXeCDl
wZvO+XmhskT5i9ka3LRf5DFEVEjHRpVwcEhjUBY5ulJIBLnn/s0ZoMQaZnvKarmV
tthye1SR7F3gP5H6pMCCRimA8joiLC9bGm6B9nBW8XYsYl4Ldz4Z9G7N7mI7TvcB
DLKbYcq3biXeWvna03a+NHBRFdkDK4VXQ98se5uRL8Iw8rltrpMC7sooEce7EaCE
gcCgsNCRbSAnlyzU5L3tUcvYgB6D81mMK1FgprAnWFv0RVUn/V3trmJxwq9RD2uW
f9pl5d/tiIFmcuUsRQTUSR76rO7lxlpYZ0MUR2jM3Od3B3/AKeeP5b1xKJcFcFyu
8u6eKESJSgu3DzKj34H5kcr/MIkV1yFj/tVYaYhKE5Uw/EI/y4VRyJnY88ewKkCO
5fK8SjxL5w29x64E0HCoUol77jI8ZWzTmIoHKm2lsoLukbMP7qHOW/scJOWNpHDd
s/U5EmOgwddw4NIsh0lW9iWezzjQd2nF8rBXDfoudffLdWs5sAiefVueElBbSCeO
OJviEB0KpPC1/eSbQHWukCqGEcKXEvjdD+SMJhjrGxfU+IiESSfrw3ahBTmPI37x
oLFiUP1LzelYEfCtC01K0JSFzwdAdM6pIE4AOrmnMFb7pnJCj1myo7WbN3fPwmZ+
Y2ltbUIX6cqOvOIgeUtBS0U1ZDA5srUsvDpF6rERVzlSJ3ysEuvp5xruVSEuG9ax
agptCogl6IdzyYZpRTbnOh84XY7HZAyp0/thlVnFQlFg2IQVp/VDmSMzh4zdrjH3
nBHq3Tpzv2HobcbQEeSUCy3nghWcNLICbeRI3woSO3sw9nn8EonpSR6l5K+xQ0Lo
Z3zjeY3jCICj+dFbos/yysGpKW22QJXAy0TffkZlYqoIk/QKuY1VAjKq4lzPjCO+
ZgDLgExdbyiF2Gn0kkokQYPj3VNPRnV6O2ftgX6TNQRqhuzjWmMk2y61qKKFFJN9
inapqYSZwv1FSU1sgF1T9owDCpR+sD4UHkJNmPDDWmrHTd4pzvudg3YN2fJlvVrH
rQbu2cxSfFL1NjDqjS6oOA9x2Bp1nLy5G7fqCGasmF7iD4IpBkZQto2mEd6yeli0
xz58hYaaz+dk3npuGEagYZdfI5r0u55PKum5oTxC/6PJDRm73q0DOqVVJl6u4Hem
Y615jbSHV1KGluCfByiuwMg2cDIFR8RQbANjIQLkgg8hobbXyGkbsx+vzqw6V/ff
xAT+C0fwc+7xcXX7mJG27bdNXUBEHXJ2NXopnJCdlJ4TQPdvk2eSqWX6fkUURrwj
Rlf/bopYc0maJbQnNo4CkTztaSTvGWBPzP37MsTdRlnQ2e74BlF+jFFokdPbWbss
8XJ7q2oIqainp0Rusyx+gNy6H6bfYGmCJ1nLHDhdoPU75sHqqhR8G36zxsShxixZ
WQW6U1PLA1ym61clRjswgS+aVbq+WAywWkUaGUB642u+ZT7PtdRvS3AHyndnS0tR
jM9z/dljvhrnwOYJlcqyEevR0/ft3BZlbBblXLw3tJLqhCTlBHbidoVgJr5NdWR8
R4P26zwXYtPJGt1j2gCWQEx0ZeEhSDo4OIVczhhHVAW9gdyNM8wbdl+iji0FQ9z5
nkYF3pS7CXaan+Kv2NZCg/avkW4iTpdUX6bxXSivEHOBQk3CEeIElcN6nLQ0gFa1
5QDImWhj8M/whszAFRVuG0i+veR0ahSaFfahbt/jNakkMjbvZQ/AkvSG6Jyxzmps
WWuFszcvokoywDoK/wmaUFpJtWWOEk8g/yfn9eGlnFyZcummkjCalhdFS4wcNvz2
ulLI51jdBONKwvKPjxhJtgBpw9T+UnKihXQFMj9zUPm8er/F0OvoGhlTLr12JGSS
C66i3SMfaxol+j+YPlhdx+1pOZQq+QymYery02ounm0Xy5N1YBGtDu8GjfahoIs3
oRtH6bSi/eLFvH4l8dD022enzcne0JbmKfMJ3is/SHr/ipkcyxrHTDtOsInuNLag
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TNLCvWenMvGmyRaRjsUfx9zKvYpYg6HeikveCSGtJkxC4/zh1gZm06d/9339AW5y
IFnV4vuDoBadepkmaRG31xtxVxo7tIikS4fFcomjAcDw/NjGFvS1Y4cpnmP2bsiI
2us88a87KLUKrg26dpoPlEb+5tLMeAS4n7DKz8UJ9VKbtFNMYfxZmmiY2SvwReo9
FjBs9cziSW7ocCTCoUjCwSSedoNDbBVzcQxtbK4YYgfOCrqrOSiiRCod8HH6jOTQ
WOrSXBYCD5qJOHyeTSD4caGpFIn120Xp/xLO52RUMTjIg3i798kEzYjVLrQTGqI+
ZoF8Cw4ui9hOrdSTqr5RrA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4720 )
`pragma protect data_block
LC5ly+2a72KC2ZuW8NCIt5jWw4BNE+YrxiDwQdWbq9rO79kU1wC8SATrpCDk95dQ
cFQMdN6TR6hB7jHxZo8a9klCaRmY94X13gpZsTJ5e20bziDgaMEOUPiP6Q2dEiu4
WLkZJsFLGdILlKVrq7ghy1TOZ7Fal76ylmRZot3pCIGS7KeyArJttFEsaqIvC6e2
5JXWjilD36/MNKimlQZ0yrSK04QRVyN+NEsE9FS69Y0bkBDZdHFh+Ad4h367tA0Z
NRoQ+OEfy9ho4MAU+XzSM6t58YCuZ4jVdOeFtkXtfQv+G0n9OQTzBsx2Y6JRCRne
OVdIEPpObhiaYZt+Vh9ZCD7ajYnUPMJpVXs9lHnQ/XumGCSPiGgATMkopBtd3nfa
8PjwqkR1qyRp3smDqkB0C7w6J1lz1toiY/w+V58af0I2gyGHS67g56hApQP6XBqo
VOHXxJK2s2y3w0ax+HKrST+/k3uDMqanORq+T5AV8daY7/fP+j74qma7QmK8PEHx
1JNTxeigrSMYvh3TIVw2/g5aV5nplTn8kARnDhXbmMRBuZQ6pwF30nN+0DK9MyE/
TU9Op5M5iZ0vzW8IMmGLt10kqqcbHfTsPdki9XAhTHnKkLDoLJsHb3qTaLtTiZib
NtR/n5vWzrBsxf3Uk1nfJCtObtgToNLGp0ZWKY82Z1BMVdaA+6lpxImBl8Jbsm2n
uzoNOudPALVyw1GAktkqQ00zXVT+upyFOuFVhis2undueJ9r3D/XSY0IpL+YNO5g
raq4mzS0Y8Q1RjZRK+KIa8KEHP19aSsT26n8b75azxFCrU5mapxpunVvWj1YgQHW
8cxwtBHu4f+Ajf7/nVtuV2nnOaN/NC9psfjAQkV+xicJyo0tdwQRb7NWWeYNslf+
jHCj59Ilcf1RzkSe2xqZOcl3xvIQYCkV8Z8kNBTTP9mu0lSdayhcUUi4Gu88f2H7
FEtYnlxG9ZOlqMcO/NpxwkqrnFUgMMbzRM5eBL/I6dfK7nvJoscDb7dLT/4314mA
p+8ys7CII1Z+ZVPteQrrbnNvZwj+ZsFxTt7+Jo84V95sKc+CNmLyLxYTbOZZ0CrS
yHjaH5791tejOKxNzG1CWcGHeFEA8JdS1zOjPgn1kskbwRp/QTZbTaA3UdJojZ8j
dGp7EuJpCQtT6xjNyQTbbs3Kn0gAH4yynL5od4CKptQeqBh7UHkjAmDBi3Y4LQ0U
uFTu6naaTylFpJH6ovsMIc3rP+OJer2HBxE6DOYVba+thgnpAUDTq+Vs4MFaiafK
17fRtwOx8aaYweTFsmhgJfUohF60VpwXtH+dRBcxuqNfR04WiNRuRYAbzlQNEiuO
AaFf3ywl0mXddUw8rX0rgOM4fLX6yHMcMjsbXifrDkBH2xyBCuMSRP07ovGcCwVt
V4wOpLd0vvpr0wQF3Ayv3S1iNuuZwsM/fJM2gPUZ0EUqwiyCUZbiSm4i6rStST3i
rUQeZAejIxykKf5VA/Rv8kBUYu9JuBNuvO9wVoXgg3UgGG0envi7QGGE70gXVqu2
/RkDpVxWg95LJU+/VVQX7lomVmUUobOwhuT+MEkfT+yXZXU/SMv+9V+yD4EqmNSZ
9XR/pTyvsHp2dxES95dmO9gS30By79B00C+3HBH1GFSHS+nE3thQJIBPY1sGm99e
y+kbtKsJuoz8g8WZiM2hQUigh0tkjV1ezNzRyaIomE2oRAcgwhMQ8r5Vm1xOslsv
mzaA5Y9vduBgpkW/4MpFmJ3U2Oo38oNDnHZrJ4g/k7mpS1Gd6OygRGgk8Umj8obW
pib1ok5kmoI7njJCyvwxOaPWBoeVO6ypnUO9mMLBvHwPXAMCxbpzjHeiUbx7Ypdd
OUXXMT2efOnd6Ediv/x+/GnKu5GWtObhaW1GjK8j4CUe4J6G1fLsuRJ+dmce+RWM
yc9tGhoJXMES8a7H/C5GQKNBLdgBEmet5QboI1Jg32WZN4LRVzV+450NLxiEleCd
7DzHsVRU+yVmQYSLhLc9oy8eTdx0TV+3wW7WHoHicgArUbJtjlEOqAZGa1Ra1PaH
TEKM++0yxj3Cxq5ytfp4KsE/nyva3UuWBcdYLOWLQpiln9t+p64hOng6l6F64mbQ
Q3fx5ZEnpket5ejWQOOYgPIpQiSWeU1DdMhJixp62Y3sHjKIh/KrKCrW3EuctpL8
pSHUgKANNIqUgR9uUTy/bdtjCszDpKcJqtmYRTNZnDkRUzCkygogoFw+0QgcW1Vx
P/1o7yOcBbXlxwJqpBISJB8xhA0EBJcfnAcOsFHhVVI4V7CKG/7eki6dLL8N5tzg
j8lHjW/wPRdyMAp0XLdL3sQ+/2+gUDF+dg9jGUQZkTFeAh+G4Z9VI9ZXVaEq5lo5
UocetKxHAiPkQPYzEq0Mt2kZpAJ5VdYQYKTwuSWSd+pupXvYy7w6CKyHfZBZdVst
eOEXtfJTDEzJzz2BZ35kee6d0/gfulo5IpucdxqFKTMAYqBtauvUeuOVMYtEl2eR
hPzh3Z+uqTu0z4FCFF/6p0K8TYlJOOshlQqxNa+OOKyuQkp47Q5gvfKmGU2qTBpH
80CIAayXfUdadXQfE+pQVIHQlQDzfNbzzH7B7eBPDO6jqDhezjgwwG2YEZKBe7d9
0oQJROHwXvytPX+/YRvCOv48XpMQrmazE8aM/b2X/zE6o/7sC2uzVwzthdBlVD8o
kdgct1DPbRFK02s0hPV1lu1SiKaTzs97dFgEGaPXfs6jUWni4+CiH9X47HRPcaUK
zCUmvANfHX7uJdPV8J4mCsycnhNSCBevYH+mwZP8Q8E1Sjzc5M77b+mQSFm1WpGN
mGelTSAx+x5KFcyu/B4oTdV5Hbxwz8ep3Vu/XhB1GhReDj91l6BKtKYdxUIpsVZ7
h0D6JWoNpkDqO2c/TVFDWRfr9odbNBu4d5nfn7EbUUjETb6/TdOK6Vte9hNQyJ1J
+Rq8dPD2HfW2JPO+b/ZEB8VYDCvf21gyjbIABc5U+bPIiFRv+TlI+ybz2dOCgcRy
QCdcCNJ8bR9U2MR2o1KelwBqaYduJHLERcxmxBgQnzK9ARCwx3IHDtU/N9dla1Xh
te72c2lNJ5BivPda7IRwKejktLarUKcZol0zUAcgp+JqXpilzFsGJUojfXMSO63v
89z5HBmz0ICFg3TlV+EjaLHpPtAcYoBALQZ8iTkz5yoxWF115rULidOuS8GDg3zV
Bpdmix03ks1bfOQ77q+YavORjpk5OeVI6WWzEX9Q8+52D9Zz3rJ2tYhoBmrTGgrl
zvoi0pGxyVxLnETliJ9ZJfcI/bzLi5UX1kWqjxv5olpLe7g3P1U+UyKjF6zF/5hR
54AXhsVB2yBX0iksb8YvSQs7wz15YFiEt/yGVmrpFQ+Mfx/ffVwhvvaL5oddMOfp
mvew/LYhtrRQqRzmSE8nB6IbYp89eU0tnEaoD2L6wy18NNcXXPbwibQ8GiU4V95D
ZNv7wDXLI8D+AGk4gMZABhcLIEsQNmutzGaeBOPL51/6JvvITYPjD5Z3oUZW7RX0
ROPPDgKjjiC1W14ICghYzt5wayf157UwrAJY4ckIiU6EDaDSKeZR4hynHPitd7cF
4cK+sBZecbypdte13WDi4KaJrSzHIxBaaCY7vFDtqn2/guApa08PuRg0Bl1e73eA
Qd90bwTk0l5JqK9d8q+FM0obl4OV1fyGdtXyB0qHxldJVtPwaCM3WKb+kXJPfxfr
4544kUw4mlri9MGTbSwoFvorCQ1RROCfUXFMXamqaXHDEdz4tiHG0PMsfkqtXFAy
fhQcUsXRtnBpX/XE1yOnTTS++iZYIdcMq1jPNhRfF5indouvTNpq1rrXMDRQ4Evi
wPWwGnUgmCNUB2Ymac/5M3ZqJBsLmtrTHJf2TCFIQ1Ynugt5iTU/sFSo/Vz1oW72
ftMzO8RG1LGPPSOF5ALEH42t7dJF2jTB/FXa3roeBlR4UqC+NBrkVOBk1Xh48BCv
yNvDNeMzcUQt53tX6FR5hn/bkiGjO2rKLrbR57rJ83GghMiSZuI3Ew1p740CEAEE
B/Yi3a25mfGnyyTLOdCzwx4FS41truxXAqaQ/Cha0QHrvcbxhMaUnTGXi2Edzldi
THFyESUwRE8W7subzvXzSh4Q6LtTC+hhCtUVYct17zgbGDG4fUJutOUAF1wywgUu
5LXsnKhgpcB8nRUQXWyKiNF0m1mhGKLk5wy0d8QJR3JYe8sVpR6xqQvT/TRtZagQ
GWIDfUON+z7noCD2nFpJ1tBCWDEbu+QS+MvK4+KbXc8Dz/wNh9P/YiXRbK550iZW
QYrrcwggZsPdvbmhlFCFNLH/zsJKy9YIRImhRRurMKtHcbSjIfWI7Fn2i4dDwZAy
Q3rZqlIffVwwySxRVTRh+8GYtWbHhqRiffSx8xn4yAz/QKhoN1kp00xfn9DLr5Ai
SuVpYgckOetEXQkJ6xp9zG1NjvCKtcRHZbPdGrSEQTHXvpAmPUcfma2GEaB3Vzit
KHOHHQvZAyjx5Dac6VqevQLJdmBPt4GccScgjBF39CfKNji5KB9mHRwOitAV+mGh
N+hMgaT0N9MChBNME7/H5hCr7y2gV9Ww4pdCIjmq0YLwMKEw/nVn4EjFAxm0uMEg
bQwxoUJSii6e900tXVr6acsPMHYC+i23FVhDUncLsSVOJX7lsNVNtJVhsHH1tTqc
Rd6WLnms3SmAxAWVYuq9e11GHz2wKX+w6tZmahGDMT4xoHu9mp4y5yoGybWdaHiZ
b+wZuT+RmOnkRab9ft+pidT6il1n3AS2Kxy5UiFkq6dWH2ptdjMV9o0VLXe7+Xcg
+tn8ATZz60zdIbcl88eYmWOV4kKsr/xGHRKqv5n1cvWc3755WfdvOimXNBoQRWXR
/ugj58W9OoV8fPWI/bsCAATZ9kwzgNcNRScfeC/IDvYkWCyPaUTqiZV9Zejmb79z
14bVAB1DNFbZ1U25EmsI/pPDtg8sSKuEvAFZFjACRIcIF2omSB6KjtZk6ZkMtg51
Pqhi0M2hP8JfW4U1IEQk7nROGVUDX8djvYR6p5WR3JQS6Iql4yiHvq/OD0/64537
W5XTLpuDhz7upl4VTG6DKK2Iz0hmZiwiiLTL7RVileCS/Cn9KZUZGUEK9765mzUp
SB2fF1GuqCTYMi2vUe9CjvRWpWSoR0anLnallMbesNI1/K5GdlQUNpULMNXfKiMR
aBCQQYJ3QHMb9IY1uS7l7q0jw9np5fGJKOZb85+0Nic+2935l6vda6UKPc49+Ds2
kFuLMXGLBdZd3i+67MZbVplQtZOnf9Rs4HToFoC3vgdi27FAMI62C3L+jbC+8mHz
w0Zk4NerPo32mq8HvKu+KDRjqLeEPoR+XEsEj6EfvptPytL6zz78HZDLCtc84x//
wfL2MT+Fi3lOhVQc5xyVa5hDlZbJAHJYW7nNHK7E8I/6IUxIEbnTrwFw9+Sh0LG1
l7R0wYb8N2ZJW/dnm5Rhpi+ulOqEct/y2rHzLRjMOVVgx68H4KOxff1CGOrj+SJ0
oS5WwlYyIVkUABWjkuyO4xGKCa/tT4nTAlf3/+RwjRuf7FxmmPk3TvoHj3ZEArlL
qArPXYBS7ytso0NAK0yOG0zhgfRFInuS5B6n9k2jwdvWHAVVVRSHAmIBNEIhuNT1
SVbuho93ib9v+h4pXdEGUNwRlFBooTNNuZ8a2++v8Ms398XJHWxUYQatqJOt2wkt
+4YetlXV+m0qI5vW6/GRiCXqLHHaosH+EsqP84OeVA2UsUToQUwIpEohFGthyvzp
nS5gWjDjENfJk8JursNz8F3CIuYYfqb+XL3nyanF6iQEsEejy4SoIkTY3VRtTXAB
lJFnJg/Z93ynTQfSIpsvPC7BDBBwrRqeubPW07B2rM1nMBwnzBeMODcHgrupdIUr
IVtNUqhBCJpzmRlmNY8HOeKsE13IxjWIVDAq9qyYWkqPBA0ODeYEz8+UFaIITc59
R1i35yetbMfYOoO0oRM78ZQZiKjgIcEbioeSOO8b3p4UkI7P7TsfSETecIMuf/JO
a4yEn2m+s54DIMXg7ebRBp0KD/EzqIXDjYqJI2ALPFNKkjIbfpVMQkapvlcKmMoG
MrDC+TrFcra431TwVkF3RQG85b0q1tMjIUDUaogeq9TZZb9jgJXTKRepGPklF3Gc
q+4Ftxulm4BU8te70XqmQxDtSpnM08IBDV3Zsv1q+RQ/Afc99P/kk1ZvmqxBF+Qp
XBm19qb6Ku8Vz/lKx7JNQRRglsB+UfZr3oejbeEJpPW0boMXavbkOpIZnhDuhALe
KrPn6nTbzX0Juqj3Y4mZSw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dy+IR7e2abKwx+gEg+zf5lF3jZuL3mETkhOl0vAt3WJ5q/E8i2NEyKPMjVhdIvyR
66SOsLJqUO+41m8gkBWS3ZggbS9WZi/jTwAb8PA1oX5QQ/6ylzyYMVMHNrfc66TI
VYSh7DqTLc4dXsfB+Si28Bot88BEurUaBtw4xehk//7wCQ4TlO5DQPtF9s5p+68d
fvylcfMXWNbgTMYEE3ihiFfDwnSW1Dgl65fxc9Bxzv6lpePty01YdjmN8z/JXdQ1
lC3mRpNe2xxQAq80SsDvtK/pzVLZ7arPa1n7zO4GdzvSgdt1AKpnJRnxoHr81YtE
RCLmaIbyLf2r6WzcdcO+BA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4288 )
`pragma protect data_block
UUYeKrH4fzGdv4P7AxCNVMTJ3xT2BglHy/CRS8rSH1C6orA7U9sx542TmQhn+U9R
lSYvshHimUWipMpZH4PKICSj9Kq1r4LJIFt2B2+h1W6yJdfL/CDBE8B5foUpYeto
jNLr+zPOyEbOtD+xHC3ObGXnklJ4EoDZDYcBp0BZis+v+pTNUMGlvE8mVCIXmm48
gFF5xTxm1R1EBgEQYfFVzRZvGl6THNMUzVysbWleKH1Ecv9B6mje6Tg6bF5TKzLf
UmSV/aNQnhuVKNqWJTT+iD2D+C9WunlBrwLCNsLmTfJFdjMchjtRotwKTPrbZHaA
l0IkeLXWvVirFwSiTA+Eow9Hllb6Elmo5jyvz3XpVjaRgkM3B1i8Xl/tQCDcvhyb
6ihCYIqRCRzz2GouYFXZDlhGmZJIzpJXn4g8WMQS061vg3QsViF0KuHtCndtMpsV
y+f/ZmUM4HNGumex3JaIVF4pS1fyZ4UZ1hlv0bR7dDqQ0rF89RwWf3ZxMau6u2lo
i76rl6ZqWX9GKB6WBSg+mgTmPXXRBcyHVS58HKz9dwrRX3S/8M5Vbzxwgkb3EhqN
Za/q9KIL8FxIRU5A2fosu1h2mtIkg/QaXlrRRudqpcMivfHBzsRIlsR0/v/JDXtv
nqXcZREmPltmulUPFEOPcyH6gcYQJYbOBsRAt2k7sQCmA0ov6UC4AE4sT5lcMfYy
LucvWI4PVyVfWT/k3NXPh0zpplWCESPKJ7NjDJOJeLK9y9/SVFky1oaD5kA4WK/F
lw/6Rjj4YxNm73AoBaN2+R2kP+Oa+/esDfz7X/vbo60PcTSIqa/EfAd/kY99Z2+J
frTqsasEQgejXDMmpFu85H6hNstXiusNultPdKNlqnVroKAmsx5Vg3oD5atWOynB
jjHFFdrHNRZuJpRY2bP8qK9LyXV5uChvV9nCgv6RodsqOcXtpmh6cS20HwWmEXoN
R+BFPWlky3fEmsnTtItx02ARWYI3NZ59gX30GzGaxhLUeu+Tz+NQIKBdAHCcDHsn
giwcMP2Y/c1/1qkDdMoxrVtfcpNh+dSr/aACPzopePazOCG7UPrSRgwmX5TxtN1g
aIR9D5H9ezKpxBW46UV/haRkXU7WACvIdCAYouy0U7dBXPQoB2DHLJp9pKNt5NmQ
S7+o9MbVKjy9lIAmXQe+1miWv1DhfKCVzjMEVaMpbwGUgiALLNN7bhaya3wzew5E
zY5miXtgmGaubE7Ek5VOvDUKLqIhgJVxVDbbMuKxhydabCYbiXJii8x+Idg5TPzu
QZG48Srj0SrNs1xTAsidN2jZ5dsNsRczcvzhE+vqw2hmykCpA0KlzJygJ6w5Sy1y
i5u9mC7m1wrY6tED6jsc0aYkh+W/ZqyXAsoz8hEwU3uevH8gz/S1iPv7CZ0vGjwV
8rUNjg/z85gSvAXI8Y47PmRj+sOiuf2u+17rSTO/g/DCEuAOYtoPFJzDUb+N0yUq
W583Zd3CSyD68E/k8TWAjiiHhsqD5l05Q6gPkuMp//Qv20ynrFyqqbaBcKYykS/9
cnlabLJqTn6OzQ92andNa5mywyd00sMO/QufifxqMvCovrPVuYu0WXernrDszlFn
RKPK8LC1HQHwLdZ6Mk4+F3+kLbA7yCINfRmcpGNx46pjV/ayFWlHLR39917gi3r5
3Il81ehTSNrMmungsFmYSdogxIcfP5dtZv/32+jq/g+h5YvYuWdv1WYbJiGNfvg6
ET6msoVRZ7McRMphCeTeCZMGwn5cSPeb1P1dyWs3uUXSdig6vhUKFNrju1/ift9R
0idoa1FHrWwszqARisDssZUOMTKCFzaxtjuZiDgRN88RyPqJZ9PQMDinaH6DfQhf
lYmJ56+heNEh/J/bA9dkCAHVpHOHcnaDMSPqn/oUR/DvDFCXLNnEATAQ2DjPrikv
NaKrtvlp3crrgjhDJcJxg1fAM3UW2bEdZomVuCXDdRQynlMA28+KP8yVKfde3ejx
bnUTTXRr5oxobtv66iBrJVUWmFHh9TGAeZGAv2zHpALvVUOwj6iniaSiu5rMMu9g
rMy73S0u58vVe4nfeVKVK/vJ+sOzEqYpUN/M6eo/enTk8ASr4LyVPJmjdxgP/A79
dBtKUakD8SKTd2fDHzDJ8ue+1BgtGx97fAIvgtDrOrDPTLQeIgZHAnpC4rG93jWI
tvMykLdeygLr49+9S557KVu7f/aSVltdjqE0USSm2+DOMImWVDUMlrJO5qjhGE3C
O9GpD1/SsMEobS78E8Oy879VKSs4PiJPQJCR1UoHF8+o2T7+IgJBTxVP/KpzxZ9l
BIEqsfl6IoLtfYmR7LKySBhQcWgyZxZzQeopoG4e+33o06FV2z2OEdncbaaap4ap
ANPF08ob6c4ib08pvh3kkIAvhmbV6f1qPCipfA7+AGkIJBQ6NkMv7jEYtR+iibky
abloQgLjt3k/RhlNUC5FA2xsZq3VnSUc306a54LNvoK0g2RH9j0tFPUDe3HeIwIG
CjDIIyNmIMb34BQ1wnbBZRpX6XyRULeJggZi/57nmWPwNQ1oweVX8feTKLJ20yeH
SXDBEj309butWNYGqa9lz9a62eLLw0Uza1926IF/JitUszx20eJxnfpSACDVjcHt
+i2ZUVUJrG6Wt3QI2G/lVBYWCkda289b0dFOrDd/sslaJBtfnaYf4MDXyprltdsB
6qWuv8TYVeXFlQSt2gfT7b7m7BiAT6abtBIND9Q+fCT5ziCIybtQUsKGxihrz0qj
NjN2M3WVzkPvyiadXKvRMb5uBBowFzwslZe91CwE0visk/aW2xZzCAs5S8l5kiKY
v32R3cH46ZWbJN5wspWgRgB1TOasN73QLax8rXa84RcjGN0WKODjB9Y9jPLf7cPx
G88snPsbCuIosxhRo4nwAkfeDPlwpjD/7RpcKwYhawexl8ZR6Wilf4oWEWlgsqP5
g4VJTK29oSqKPRx+K5VBYGVjgIStE6hzFlxGDeOh6qDIhRWJIf7l10WROpQUdvAk
OZ5+4r9n4IbwcT98FueCi3fBR1o5HhRx+5JDkwP//t1kI8E8dPUEKlLv1TAFn40A
RC5r430OtNZNzoTDXFbtVGVtZeqIEd1i3xsAJiop1S1ap2TEzelUWP0oQtX0W/r7
r+a6XVQM1iUmZ4toTFbvxCoH2CqZtm+gt72lHGJAC5z9qqskzuth47JMi/T8eC6I
0pF0wLDOICPx0Ha1duLmUwBw54QhkKoF+pvCXirjIbc3zXmrKYYOKgMLbuvDoXv7
72mlwlN3SIsMqANSCZzMfZ/Bd1/WH/VUCzA6GYZ5FCZDlRsNJ/sFiR+Jnnj8UPP6
4zhhUoTcHBuSXMdZKvwMv/4v0ZRHsrKdwpKQTluQkAjhVCcuxmaLlApTXk+NEpT4
f0RLQHG65U6+SLCjE+yXshH+Hd3IRQ7cfBFxQL2PfDbO+VbUhhFgZyXvQodSNnCP
hrnqhC1OsA2iXE4syWmlf3U/xx08lOuvS0/qvqHDeRxSmwmXe44kIqODxTlNAh/G
lBBgtIEGFOWheQNCN0KTE6KIHPk2bP4kh8IyiI9fD31wJBUJYEhovpWy5cLMZEg8
QHSVt5MQ5NNSbPLa8kSIuN5UJHJkyWFDtES11fLilGUCjElng2KVI+P8aELHxv25
I37O+MUv6PplYpDj80gNVUZ3FavhEtiRZHY+rK8Adboo7ASgFpb6SizE9NKoP8pr
hKZcTaVhlRCUkBUFftnr9gZAatZ8bRN5BUAqaqeZC+dcCIsn+Jk8ElqqU6h1Kgh+
EdjhsmUSMDzZDdsZPveELCN0YsvJmLhxXcaf9Zi64Tb67n7qbwzPbKVjBB6Fj0Vc
bmvfhTvjJumKkWWhG7hnPiSmysoqdT4y063Bzvqm+Rf8f9XUfVpecCpzLD2hgfae
svYCq6dGxvyiBHmv/YzUXQm+xVmoi7q+cCb+FpMbs+eyhQpqLUZogVBxTIhjsfII
i5Z3d0rJwvshKUsutEQ3zIqRYmHqGRsOP8GWqIK8cg71veezfVN7tQ7BCERNpqK9
gOcIlxyyH4mSI8lvi/tsmG6vQvOe16E6YKjkR7lFYFCjNQnB8OJe9iRo8sAf4tWH
Y4ePHFUjpvqozKNx+UiqGLDAQQmncO1FPTL/FmwJYS6rAax44276XGNWyRmyCjK3
zVrkJnQPvoyk5zVbdcHCOlZ7NYB6ItRA9KAm6d1uW0SWeXppjdvIE2G+0nhwwAJd
Tj0d3kOp85BFjxCIBEpjR5/SN/O9ErGv5F0+PuAv8EHiwapM0dd083wEetGOQnkM
6L1d/6se1PVpwucVGDJzBN5xjUTKloeArsMk/1Th4VaQecwne6g4PlNeo+6kkTM9
vqFdnAH6MqVWGQvZzDXHWv00zAzHjmaCrvDI7IHxeuo/fwNLQctg/0I7tmVLgodP
7TbASuFtDdTiZRQqvCeb7LyV4j88JaxwDex3nrcW8D/zVn16tIihtzmQCtmuMs68
DZS3vrcWchM/iYqfgJBRPD20GarAuu8j9Ff/IkkWRydGI7mKMxUiYiKkVMkpO5Mc
9vQNfwhnRJGo26y+vhkZpi19QVZT0zlKtpULXl7DsVwqewXsoAXY4Nxs4M/dpbcD
W8W7XXL4yjG7MDie6Ryq+4q+1TJu5/p/m7xaw6JcGWmb9+xtS/1w+YrkmpHN4PW/
oEv5EoXxohAcesZCCrs47uGOr+UzYIuuBY7bJoKtu3jvE4u+ji3qxsN01InjHNEN
PXlXK81GgvVlLZsv1mDdohGvUc1aUXRCsqX1LELEsG6Aj5mxRyhAOdrKMRbBfz33
xtx6mrGHqq3J0f88BxT7j8nQrRRg+XR5LDLTJISggzDuavxItcBqDkeBlqDWlV7s
KXN5LrD4ApQQIChsI7CALlr16JPH9WYdiWFePjHGC7vW4q77NHSh02tAQOLi6DNE
tVgPipiD0GzWDemaTz+lhxioSJ6DOZIvhHJ2PQIDHydDz/yGZQbfqiN+TY7vTatd
0yPC6WrTFAHkWV0PmIn4k8YYmQjQmkxv9VVm7J0ixBua+EhyF/AhEBcIrrvukk5m
gLEQ/n/itaTbOCi6ZCQH9H7QqPa7KYKhPpfEvcGAPU/pwGU3lw2DIMbqzZgQKYB5
1If+EKv5fok8RI74QZ28DIclGBjjk766odg4igyIg+YyHxivsVXoXLJQFbVQvlzt
dNUc53uALPGOU+IIU2ZMKtRsygJMooD1vc/+nHjlzUaAhUWSWe1wF9Yy6QgQKhfE
3Vce+tYm0aZMIKOb7kgyUd+lJDE+67dSdnB8xpAQ2A9/ovd8yF0gZ23fJD0GOq3U
ThOpkYi45c0hRr1A/KYEXOPthp/DmjyWvRV8ZYGUvvtAhCh30fuFdF/H2kggfoRf
k8TGV14UkZURSO1E0vyNM6OedVkjHLW7QpVTZZGkjg4n4cKsOgwkoGHp7xOw1lun
9ZDcBDffTn7HSOUwmjbmbbsTfp0Yf9u29J8kDZih7/FkFcASHAuKdKJ8flAkire0
MqqFS8QQwlLgkchv+pqXMZnyHm5Vd/l3SFCE/3oat1tktViuHpnJQjHzoYVJUlp0
KylrQMK6n+8knTul5NuK1AwINWEufI5RHCkWLOkBNCqU2iHSw66dm+6NFybwAfGX
1jvXleu1nAq/ANqnU6JaY5gVjhuqkLzdPNfeYNnprmL6TQZzyu3Vc/pM9V/XQxNt
SZ0Gjdvn0KejlCaCxdTZKA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RuMYPc7nU2WU28gUogce3tVP5wSCOsDa6g/9goETRzFmg3EiJ13lzyFvUGQrxHb9
NgUmf28TTQP/mxRChsO++uYgsV2BvU2BzVEe6KsvRAVY+g3RoqZwDwpGx35v9GM2
dZ/EUkWYWQ2d/5Ak61lCbcH/cmrr17mv/W7J9qR38lmQ5+1xyOOVG1ng7eFxQuoW
vk/x+eKAnR//WZRI6a3DfkPsHtkdbnMQHG4kNGS+QVNisse1N95sLVoPxYTuK/Xj
HnLfisVlC6PyguGedDHZexUmjdONBhYrIrhlyfMMacIsuZDWkQ3ySC2rK7iNc4Bz
RnO+0aXgU0qIOe/ZhCadoQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
In6TBz+EkQegU6BgVKD4fcoAhKYoQOVHG7UJ8AoKhtjAYUZm8eEHGFF/yKMT1JJ/
pJVxYDggCIfK+r3eUtjtu39d+KGyd0WtGAyMYMcWAVZUV7sQ/+Bs22lNHyC8j+Fr
I/6jkRPPE3MN0pbmIqk2gEkUuXgbey8wfqXMVbAWvieSRYI8j2jCb7pgkaD09Ryk
wj1su7WmlQEMGpLel0nB6w+pkP2FCqFYh8sDLhebgIiYVEKT7a8sWIYE3N131Z6y
KohfhJumJmmhRHYxm7q9Z7qJ1SgUh72u1T1vCplVyjzqHGMgu6MLXLgQ+ibwx6yg
U+Tj/hRIJjWhg8RDDYUtmIDQSqqJ7ke51UrSSWNJ3Tw1Q9NpcxOZEVf4icxddpez
7XmHHesYvnLhG6e6DxR1nbsudWlbVdWxK2qTo8qm3r8ysYmAN1+nRfQoZGKb0Ld3
YPYi/W4rZucIgaSS8i/3tqdg1U1EHo3GEJ5PyVqF0BcKnba4Cc2YJ49T+JVZqdcL
bgkN/CD6whoKWiACBn2/IHahDjA10d54iZjU18lPM/ac6ZL/ENIaPLD2JhlDh5bF
lyNrGSx5NFWRKXOfIRGsIaR/p/PP6ES+333s3buWLyn1J666+Z+R67yvp2rlCXyw
yEwCS/2U5xDA/j1TGj5iWvg+iEcqviq23OipRc+7g+iw6HrtjfkJTYZxBcmxCkZQ
wcGQGci9kkoiM/xBQZIPdqeIzniJ3+Y6THZT3vI5B0NsIiy6Ip6AKFBoLFKB6AA1
K/lwRCKogdyJrOLBMDvLKbQndYqhcWvqa8No5naZkpqZn5gbizKSF/YZ5Dzja08J
JgjTno1Q3db6Xtp6QJy3v+S6FlMqH1+X7bM7gcZCQeuzGxdj/jkZTt9ziHTGT0h+
CXW5xIRRJSHh90eTljzFGJ7WyTWoiJnRvJQLuzimxiDXRWultGynn2JTcELcUHD9
+rmNr2ujhfOBHxF6EdnURzUcvbl/y3ojW2nWlpRAgm/n8gaFeCBBn7JpvE6Vmthu
rEdIEbf1m4E6TSTM5tSpwiwYWPGE+LzxCnOJHgJfC2/LVAl6R0lPGpgitliSbeXK
/r9H6W9+rfhz1xdErXzCMh3r4ThY6aQr26Ojq+tvyGgXjytaPDdz0taqXdo62aR8
np8UYaI+0JJ/2ElEdkMWioGw2woEi+qMPDjNWsrg6bOB7WgMh3XiuMQr/ikV4VuN
hR2IeALlGA4TJUp08Zh0iMTCVHPS2OM7djL2DG9/aPsye7LgMl6Jbcfk2qCqK3/l
SbDrArZOOeHnRlwLkMufE1eqJ8+J9SDONsSJ2OMy5uWdLALWXVMb9PNhFrI08Ax9
iABtaLNDR7JtiHIYdnnW8cw1w453zOkkgJWdkoIidKcjPAN+2RENlD/7mK2nFb4A
Lxx8ov33ULgXlmX7vs7875+Th5m1m6YzJM4StglqCQ4cAf102oz0OeWnWEJSHDD8
rfI1afRoIYNfexAV78rzqe2FnmfhlitnoIqThIBBPpal9cGDmK7erXPQWawVkcL/
WxqP2a1Ve/RauLR6KgOIL94AUUH4r1Vcn96RRsxGkeQXWINEll0bMXsuPcECccZ1
KKp1EpqynwcAMKopRX+sSzSW2ulnerK2dn9maKzL4Gal3LCTxa2XoU1N0en+HzyM
Fo/rfigkEq17ZzzmjOHmG12RaHt/xr41pj/1ATBmHa6Di+f+l8VJ4+lPWKi2+U6X
X8uqJZkm6QZmNSeFlGxl/KGr5uR65rfdMDOPzWOo68yINPJw6qz+9a7jj2hBRabo
ldWtl8wOtAlFweoJwgJ02t3zEWmjaMrOQ/b80sJNghozh1vJpZf29+e87R+Lbn8S
jSiF9fncIllfad9r2k3WRa0hTgFsRkNe1ejXtNxpdQl5Z/QVfO6gt5F05cex90m+
2NkeoMhzPQyjCl77Ejp4P825rJTDTKMcpTTeiahew0OJyTwEEgJqv3BGLeIOGUPh
0DISdqvW7TA1YjAmjyJ2opPZW7f0ICdnBrkW2jBl42fRWOA4gxAjqTlkeiq5FDYa
4jQxX2iN+hjW40pXLRskRfE1WGCR7HI5jN08YDnqD3P4D3Ast+hiAep4Fnes+Zt7
2q0Ymw5BRwt1JCVr1vbkTgJJs0dG0mmZmOQhp7KwosaRUPs4XUPKzPfmT2oSy0L0
DcvbxttU4CpNPctYfRwqcdrwJ6nIUVzyvtl++zTiLHogXCJMho7ObQCBtCusB2fa
jGiIBcNh0X1UxipJeELy6nVATnYnQ3zXbIgS3shsNJ+PqvA81Aw5OrN2IGXlyVOQ
bhIBPTk16g5do/5yAm37QMUiORB7Yisuh/Gyb1o+hMh8E0BTiV1h73qyMMM/G0Ue
hmwAhWsJat6YGpuFOTDzKBwExieA8cjSGJ2hvySN5v9GDzI2YFq8ruVJPyc49pkX
kCOzNOcFhv1CGtYLtJp4FOKNjfv7Iwfs3NtoPUtorCc6ATbusIR1QmzFxNFk0UD4
O+iHcgsOUfz9Nlp3b4yJ0AOQ0zps409g/QpkbKUS3CAo1u+MntTHKTCTCqbnJOEW
VsXm4dnVlzSwLMaUgAy+c084NKv8em5AX/7Lig6zddvakIoZyMMW4/4GBSGkaPEM
72drlOfq/OWg2gRPQ47gflf6I8sEOUyCzFsIDTNH7Ll1e/cWKOiWQ/ywr7Hc+AxZ
LmvfxRk9Bx0xWPdKkjEn0BjXZXYyDjxQICOPPeRaLlLZImgVYaEH70qHRA7bNRhJ
eeQOb4PJSsgFqBvFQ0EAYRcHWS1rf0b7SHKnfWVVyYPgCEgqBfCGXv2TTiXgx1x6
f1BMurGhcBnfHZI1y02DTU2wSoMviUZrGfbCxqEtwjEzIOr632ksmMTP0Y08WWGQ
4UnFAW+6cu7inrYB2veXv1qBwcvSn2md//w8/6/BlHUYXAXrlrZDvWI83IW1f3N2
HvcYUFV9c3pw2asNhBCavyCCbxMXNbUhu8947gTStsU6G96KKbXd9f0TkTAbfoMk
mF1+QTbFnG5yJXYA7v8+pPlcMSoYGKb6wZaMNpMOeitoyJ6IdOjO0H8h1ICm5rs5
mfHygeblOV7vlOU2v9KTQbZKPM0Y50b+C1cTmQoraH28n1sUNAwimsSwwsjSqL9h
a+gnFcdxGlgS60YMl/II3wR3ofzW4Nz5S0eAjJU7r8ogZcVLEVkC6s288zLmevT+
YTd+jtodBUaNwp4LdNdEPzM3XE7nnynIVk8iKA2K5q4XwHmluMMqC7TOWvVoiAyM
FDBEtRhw5K4SHeiFZA1KdEeBD1vFK6TyE0f0D6O9gaM2/7+nH8MmNrncvO8qnSBx
nofsU/ZCCD2rgFFFghDm7LQtVUl4lMekqJ41O/GUxmb5N697aM/YYgj0OeOmaG0M
QLYHL8/jvJ6PuiNrO5eBLmXEgujikJWCu1NHbEeQOZ3kaYcyXT0S+39TGBFh1zVq
CnYsm4OkyUQXwIekvBhucY7QZdBOi0qdFmWRb587MYx7M4eSO1i6ORGVw7LkyVF1
RxyEJmW7n+kNQjtVsvAC0F/4IfTB5kitlrmJjCX4bQ5GLbxn/X1i4bJ1+2PU3d7r
Xo4wtPd2drzeQpOqeycDJ9Zs5WPrO2FlzzCTvqPlXTT1OTBFk74hJDTIG2uzAyU3
6Fa/O6nU8D22ssZTbokO4eMaWmuvHEO6m7phyZ3EVo+Jp1ubpgg9ouasZdla5q3H
1YQnwQsS3nRHl3GYgIjGTWnkybO2IhMP+fas8DAmqWCIM1jjtxXf17of34+/9jJf
xPYkRGA8RQj/eT6T1PQeZqJuI/Iar4loYSP+qObp92s8YQ+9YaT9h8fwiyt7DgaA
MJEqUlS4IU9RQ2gws4B8VGDlrPSy2x/JE4Ckz42ltjj2LWdTX1T+Yk9YyKEdH2ID
R9wWMPMKAzDM/Hjd+iaWmKkfw6rJasV/E3n7naDmrm0X5HOl9VULRaFyOas/rOgz
m+Eyuln1/VBHAsnWosfEEgKL87HhxXcsNe8y0oyFrSxvdSAwf/gkWAArZtUqxdnu
QMe0TZr2zlhj0GeXbj/rnfUITL0aSNxAfKdROxL2A6jVS27LGn8Xbx5A4V5FP9TK
PbxAyenWxmseyWiXY7D87R9/TKhGyJQxMAcE5yLRiZtqMZzsZsqGKPTT53ytJYIS
XgS+frtclbSCZvTZa8Ua+Ah5Q2jwhzCUTStKx30sRbThL5BA4HBEo9UrIkuGB7nU
zRNPulAZMoxR8EbJDGPyav/WuXWynPLSDNcGNjXZ0xbkosr61zgRAgPNX7iYXr5A
WG8G9w9YXb4w01cYmGBMkIiPmoxHt/MKKKLXUsouDsCWjctgJA5TbUw5UnTQYHlL
kEqcez8yRzPogh1GDVi8ykadJO2TGnaLqyvaLxgyxMte60oNR3ctJx9jvIdZFzf/
f/6wNLmqvaJNRVNCDO1y3ZuKJDBA2Mjg5szh7dV76cnFtrl902keeVPZXRAzwp26
0217TJ+tJT9tfQqJGRLtNX/CxMWaWkS0u+/GsJvvTznoru3wz1YjqOTPrHpuMHe6
nSz22VvAyr1J2qnm+78ZizTLRByJD+jdYhc2iPl4JVKM82vyxikPmbH3fo8uyB2O
ZKOHhxlhhXsn30xwFcI4YKOUlOBruMumU+d/XTzTseEmLbui10324tWinVKppjcW
kK8jI9+ccZ1NM0/XTBW7R7lBRN706NLYEyB+N8Xzl6Ktrw2qXoxuHPRntl71DDKF
jDliiapUuhER5lyTyBRp3LNz8MvezPNDOk6b7UtZ6BIIW5FoGNxws+KEORMD/yym
JVIVDPZK0f1WRJIXrbHUmbCCmns/2hWDHTAra4mCqjzoHA0H/zuSXsAa/AtKnQ7q
IkgMyKBFGas+9ZEkoUTSnF59q+pR6eTH6yBCh4MbD3iDS4xGWufHpYowreNdvHW/
k8hxqT6T5pDPO8yT0vfS6h0zf/LgAVd9UCrE6Juwtkrr3NTD8qEtJA0e8NVPe8s+
QpgK59zBbHi0AJGcd/H7TxnRGbhnzdXD8RrxI7WUcMdT9l/zIYt9sV9CHUmVhr5Y
LB5AZjbRkAkWXEYD8jdPugyFrpPQcymGhnVTLDBn6AtMONHmECF5NLMnn6fUXBQb
Qlp40NxkzFzUqMMWDDT0hdn96zfb1u59u0Q3V7lfllE=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cgGITSPo6EuxoilQm1mJOWsLCeEPZv6mkzf8eEiraJlDW5iTp32u1rACWHYrLv2d
9CEWzJOlBCvFmSWutW3n36yrq89NMNgQwogZtsf6KsZFc/nFOIP/s4muwi8vPXL8
FEdMxIK9D5tJLX2FDnxyFWEy79CAAx/+h8TRvlwJMzKKS++FrtD8DciA0vvDY40w
XYrJQCUoaTSfWQ4hA2drgl1WnpskkoZdEcYqDIhmg5B9j9HeyyhHQbO7wP3sElEn
U0LkPEbBb48R8uW/yO+D/VPty+uwMPtDL2mqyciNDftEyjhjL0RxO2zzkgIY4nT2
a+j9iXaXUUnEQ9/mnfZtFA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6880 )
`pragma protect data_block
loPSwkGMUh1UAyMrKp+/v1q+T7hsix/pW3+m7tCM+Du2VElvDgcjrjHLy0pvR1Kp
B3Ol/f7wUDX+xSiQfAInTv4Bym0C5EkiEPFXO+u1Kq/7hPEQLEBKMIsDpx1cH2vn
F3qOM6wr/QayULtKqw51FljUVNUGvGHTE1gvCrQd4B3tW7M6i0zpUBSbrgrWoaOq
3FAFbLe2UU49iCnovocddZkOj5lHzfQRyFhBPVRGJucO9w/d8E4wFtdTZuFb0EGP
9s6jmUf8Yly3cqWNPpHif2i1O/m1G8CDS+I+GN4IuJfALJcvqH2JWxlEzdDkPpm5
pUC3JaBasM4hW8l7fFg9+hbjF1RW1daqCCtvRhPRMQDe/9fPdreVtqoBK9fSL79u
SalXwDDutmJiusT1DiJsd/tHNlznEQiwWoJQFPfge+zrQuFgoeAkOyotw6q1XO4J
HjJhW0ixchKtyvCX5eMoHHBSVxVr5D56SZj/iyLGtGil9iJH1Txtke2NfYtiSKBe
aIDw4VaSpa/518ebdPcGYwCwFJXFmtgJa0pZ4JbJIaZEmB7soxhaDi0syhIMZC5r
uQEwj4H5drnUHqk8jrxuBGp8Tp6BHx5YDyyVSs/YTbUhcnJ3vQLbwOxIVgv+2qiy
YBoVKjo/xyH9CmPDg7LFTldOMNLvlC9vEY0MnA0I0pa+fthpo15mNVy94tKYLNzJ
l/nRLl2lQMeH8pQfiDzx3PMnOnn62JJStVfvBgX6JtimBZdXGlYOVObMISMvAK8c
kHz3QSxPQWatSZxTPS+3Kwz6qH0QaZl6b4DXBwv8VGcPirp1S92Fa1Pwb1AjaTox
3CJct0bzRF/0bCqksYAGrdoi+1/vgU2MXJrYtbNAzBeGwdcCalt4cexBHmb+wXh7
LOoFxD16kbdmyWdOtuO7nzhnAZBBWKgVrTOJjAUW80uZZOznVrE+IbIRLUJMU9NC
EINfg/lmwB3jb57bqq1cOZBQVSbteaLKTvHZJ9D1X7eAQeiD0wtJ22rtl35cMIfM
rpW27jNgg8luPnCdG1+QWwk1NLF1G4t1D+ZHmzkow/h+YlsT88np7WT8ycVCzBSi
Iws1vmtl7QEKFewBNbA78C7Km4l8B85Os/ZqQQamYwfrGhO4G/7Q8S+orQLfkSaG
yXNf/Y0V4wqqg0zIFPYM1iMnTI7SmxaeF8Kk7Rvj+6rv5sS72MdHBNg/hHjOxq+L
ntnJO9Cxq1yDDWhmGF2GfopTF0jqCdkrwtdogQ4PZYQqxTx+Ilt98DqCT/IaPd9n
yZrP42lCQBn0Vz8eHI+tEDrw+TIeJ7tIUHn+uQAPfyJiGcEDT1f2qebPKRnPcgpV
hau2UmhCYtxAkv+bap/ivNYzHKJAdqL9KaEXRsJPU70g1KVppY1h/quYGZ7Iwgn0
LpwzLhF80T/c4A6pNwqSR++oeyQbpFiiG4wM1wWyKoTrCw2+ziSQos3VliBpubs2
em3UP7OdG4MV8HGwHjzGlc3oV4Ahwz0x9+M/LD7qZDEhJKLIT/e1jNrWghNeI0We
EU+ZmVJVgZqujIO21m2Ay7LF7Rco1ytEPg8riTO8LJQ3xwaQzDs7O+OnjSAIT++V
DrZttdQpaw0+j7LqRCPdTuTtM9N1poqZX5yKGkrz5tj3nc/oAUqCKBzM61xf1X/f
lkFzrDCUx5mUMUqM1Mwhe+OjNUnJv97qTrZyhf0hM/2b0g0hIji2w7l/GEmPUe0m
wb87I/F9OxnOBojQCenhLgujrsIhTO7tJDY3EpMduqvB4R/fzSvaZMxcI/LBrkyX
rJP78M5aS3/o5BU34tDm/GmjxhoJQkCOamCFiIpxGt7lgIxEE5QkZ63TAQRzZbXa
Xj7exiISlMS7JFHq0Kh9YDiTv8AkmW2UgWIOwKS4YccorNkdwpQ1uKUee5AcwYcy
O4IZV8tAi/nNYWB/7rjPFALipZhVzd0kCaJbt+9SWvN5MH3WFa1ZCTXI5n2ZKfjc
3Zxxb4laar2DBG+J3eDMpgDwN8RVTD4sHjSIEgMo0xifRdZUYfyX7D26Qkad82YT
BZIBjcWBJYQGzcahXoQcQyZVYnhiBUch/OOlCLxvfCNDSEs8u1EYfjZkFeCMkGxV
5fTn/kRvcQ+7I7poyMHGk02aP8X/48iLxsYbFYNyN4/VP2yTjXrUHd6qYRqHoSJq
vcz/YHYVV0Se3udVGOYEY9GhTiBZJnWQkbhnXi/abKJCNgkrY2yg8yGE+lAOGm4J
ToKXQtwfFLdlgXrSw3erKSeFqXu7njEx6nByVsjMQG9f9yBj3oBwdrLO5skY2m4y
s3xkZwL8Q/w038VlntN/aJAffPCp3nW/hBUFkdk7FAEL+2xfskEWgOwjAjcj6lGP
X09xoHrC4qHbgS+Ws3fNiZh29H7a/b/CXTuDiLaiEEj/9bvezQPZxSDj9EtjgF4H
m0Dbe0rHsp6v4RkQyIJzkxqFd8zu4FPeB3wXIaPQIpG/6GMR3OY4IluQvhF1mNqv
1gTg5waDXj1r1BhDHog9BUK6t2vq1vy2dAC7Wxzho40t4GLShxIzed0/z8bHTJCF
9NNSwCqqHWYGoU3GEHQfdPCCWvACj2m24VxUor1lfc7HBIOfEd2kZwXO28ScP3gU
8zoYB7vTJhNbPTtuumzrxVST+pNcwqC9Q7yeTvU1jlG3qzhBEvqGWBDfrtAV2oZK
8q1OYZ67W7skgQbjQm/bcNozbYLiYd1mtYEiv0uOEY+Bnb0Y5eX5L5qz5sC3/YBh
Di/4BILUOX33K/sWRFSlTYJ1jlxE6SSWGA9h66Xld2Jwb+myZO/nFOIaeD21bmx6
Vg53aItgt2tS7d4EiZEcI+nE7aoNnoP+MZbRzM4gvFYW1flkOKy7UXVwf6GME2BT
TpqnuZwf4hIMhmsZgp42FGsKve9B8eC+A2I+TPG/IyRP7UXS9wVn3xYMN1MaB0UL
4cDvm7bMf42ALa2SPqpeFlDu6igDa+p3JnHjpFHeLpwhCEbZocn3cdUID0Ko3Kjd
Uo4p7ueobYOKo8BFlwMcdPV4PQRZoe/8LvHVhYqq6MPLdlzUa8twZyppVtV4DhXO
K9XTEpsUW5DwEBLZ/FjDv9svYuiifeLmZ3gHhZHyAtuM8cuwtseeu+Y2TI4xOsXK
SvXkXj237oF6qaUMsNhrI86w6YBwn9yizlYSFYznRNR+0Sf+prJ35Dc+Yf8GsLnQ
XjJ4GMp9F+a6+72B3ZyJtIF/DWwhe7h9cfGKP0whNaoXFQmJKBoXIj/KMiGGwA4o
1YeB9hfx5p4YG6DOPbmZM4YmEyfyNETHupSNX7Q9dG4FaSHDq2fmVKhQsIDqvT/8
ysVh6kBZQMqZLHuC0SOGtO/ryuE649r49va881fjkuVl4oBXpfcx60SK4GyfoQtK
is8gV4eiouU8OBxg9Y9pEwtFRGcYHhtDD6c9VF9bdgMB6BJ/aVQZFAk4MRkgUN5P
heb6PpvP95m6WJ2FLH69fkUQyv9jFPXnEgr1RubofztiE8L4fyhqSMbx15BWqgI+
OuJFY1hw72RIwTtCWqHw7HZawRAIObhixRtdA3P+6k2lenNgcgx/L3BIwTyh9MfL
xSKyWhfwSv8UgBJa59sducLeYae6sXQwvOaSuXeR8HgLJhIh3ZqBmru1u5MZm4zo
1YJUGPd1UncfPQipIcMY5lPYKRHOVNFRsyYm6sCC27rbaO0nf9BXsa6ZPXBxznVd
E0EJnmQkoKiNr+SMk1uAi5SB+jFpGd/fVnF2askVoJEcagm1Upjs9+vCsZ6scxw7
2JF9WCEFmpQGp9BTx18D9p5iN8E88m4Y9w0Z4Zm+xn1+WhTotTVWBIHSJt9bh9yk
jBnGC2Yr5rrE2kB5zRHozq6v1rEdPT73z5AI14tZnUcIhB4KAtmC+xLdbiJ8AAoA
46yJGFgRbSew6J2EfSXaaLMKK5p3ycWKhuI+67JKFZRfD/flKhUpaiyydYnkxagH
GXBgUpooOdESgE8kL32TE6LM2/RxK6eZ2jrdP5PoVIJk0Edcsvy9M6P9UM4Cfixx
Jbq+kDhd+L36NWdWr24akYG+27XmkDQ99nc5CHaUvAWpUqv7SFJKtTyI23bc8py2
cyQN/9yF1TmsfWXK9yyNyZT8stikSdkcOnPMyMR+5F95jHTSYOMxU+3AhQmeNZr4
3BSJGBaf4pmf4uQtANAuUZ2LBGfCkAHrkiOf8yCGlakNbQ+V/fd1EFWJgYYK2+ar
B4kNqkvXNzhQatDcbVR1kKfILfqsEGyELZv4j19qRFFSQIUdkmMQm2xTW6bn5/t5
vbSehfXPVD94N8zYGYotLhhySDGe+G+OJMKGX5yq5jUarTt4AhHJpS10GVumhm/R
CL1WH0Ar2U50G45/xfHPI98ZBFsrvXWA8pAs7WrV50ZIQzgaorfuwNFjdXfXb8eL
WvvFSZSXmfkW5qffQFzEAb8BeFcQd5+wSt5g6bl/AniHAGU+ccMtDdhKXajNPoEh
jyJ5Arr6W1R+SYEh7F/+YKzGt4AguB/rUrNkpTZVXUHO6p6sjhFo2h6j9mGmTRA4
ukVcmzUW8Pn2mDba/3VWEDjm+Hcsw5LiO3ptNq7oZXRGHqpOpdkQYEwTR9uXUfwJ
1tPufbVbd+zbJGWqd/0TN0yA9WWE4QwD+u0pHdr4TNraBjLGpYQQ5Dja19T/2ije
ToSBywBjih7zrqzb+FzQYkpdUNcv3nPxNWHvikAVjWV21FtXWbu9Tss51g1RUCfS
zHVJTzvxR74WLpcT231czsZ5PrDisFJu+VPtcovL/LKw6zB5rhHuYtWn068cWEZi
8MjNsGRg5z9aaGRuAbHm0cFOlsjUtLkEyZhF7OR12KQ/IxZq/c4UIeLdp1qf1P0u
mk5lIZxpwryNrcr9dxSpi5J6ww/Np2V1r4eU0s2pRlIu1CqvqolzKbJdQLVdIKa8
Ia55AqW04bPOPE+PpSqsFFzD3Zq6kYmLJ5ACWRIZPDIQm+YT2QLOYtwbvBki/Hts
4lMEzJneuvmmKVn6ecSLqdKVX2PN7J5zIonMYZPGPS4WgR9vQmDwB2J460fs/dt2
rmQGs7r2uNUdrXS5POcGy6ayYKi3I28Nlv1piursPjybTk5FO3Bdvch3rtM7//YD
WX9FStlosWCBmwxWRtlwRn4J8JSN23ffMV8jDUHRgpsWq1nCwGrjXspkizrhg6VK
2XY2eHyD4Z1OJhidedO/2E2yvMg16b7mrHHRb+0zx0fUH4T8VPbiER7xnEJFzcVm
xeCj7WmDTsqwnMwCO/aCVDfvi5OsKkOVSRrYmfh2FZo7GuY1uObxojuC8wjui40o
RbupEaUu9imwGIO7Ts9FLCXcbI/Ms8e/WvnYNIIhxNVYpu7zmY/pEWBz5aA1UN0Y
9am/Q3XGNRB/I7IV0fkoSDtUYMzg5itukEWJ6XBaLn6RZRnCRSfl43bZqad+G6t2
kyO6smYZztEbRwN2bh88dAlrh9LVTL5C+E8pyVzk1BjP2Ji6lRuZXXTmNbxpz/Ib
Rc3/7W2mjLcA5S5wIdDxk+YtjCWE5r1EfDRsb7FybgEt64X3hnZAPfY4i+REEa29
OW3zFzLq0jWAN4PbPoaqWlfNjpVMpLTmKcV3YnUYmNTLNUL+SXe2CIPAPImUFqZ/
peS9kff75f/L6m5f5AUuxwYKZ5xnIO/GeOh4+9FulYZ74GHdNTGGxGLPNLmxQb8E
c29crIkudQsSWSuexEzjDSMjZTqVUYZTzzYn/qdyX1jddtJ1yH2SrpLacYf7jTll
cHrIBMpXy08uxXikfrZbAqGIb8/PWLAFJ+DWt6DHiC7MLgeRBLrZAYqPYmgIoiUs
Jq5xDXk0T0M0UPs+/VvPK1DKUWfomcVvoGS0KlEZbtjGrf4JH2vBPyfkva6o3Be+
NDIm4qAnGBeteFdxw9b8+oNUbEew19wC7o23guZu+dfdqTXsHqzxi518wbq4eEZy
NQ/qqb8gChnRm5Yz3EHaUKoKsSG27eSn34TKnyMzFFqnvoOMRzTUijo3ADV5VgmU
aUcYK/IIm58jc1DPxgqKwSxUEtmGpvN++yH3lbKgKZ8BOPAkWHlCCw5wqK0eISHH
tJF/75FGTJ/slJcubY+GwXe1IldnLnysUla0XR+T5PzfUpDcRIVhstqthGniDIx3
Q2Zp6AYeeQY8tetd6if7TMUXXK0MlIL9kf7YODhncg+ovQi2+3znuk6P4zVLQXRZ
9uyIWiT76tXQ5Zl5ZHvvGCgo/yyqxmGDmnRfeZzknZ9keSm3cMS9mxv6o2ivUBVh
nfuPM5EUuT0/c8C7fq/tYJ5yxkMbRbT71kSn86oITlEg7DlOSIqRBEb6kW08d3xh
2ryX9Y4gES+5UlMBhOrcYPOw8FC73dZlk4OwJv1Avi2vr0cnfysArqOET4xiyWJ3
k+U9JtOb0Y7j3VK749BRbFNelCpwoBVaoEzKEgj9Y7s3M0JIW+7illI/8dOdOUAt
AscjIQYyXzfeYY9hCPC2LlHSk4Pt+ptRKSviMgiPfWp7kXMEWQMMYYc6Pmb1raPM
auGt8oTVZHt3klQIRyzHQzEeFZG8T/ebAgM7dBlsfsbCTIqjBeGNirBJN9CJ9tll
GbmLs/vSIUUGEYAJ3D86pSgCL8dRBNxJrTQZel8896C3Yu8kgMngfnMRjUslRPrd
IY4NKa2nrOCoSNO8ATXyj5bpVqkPvfvaNVJiJDxit1qucEMC5z8lmFlyan7ZwXsE
PKHlr30CFYhZUBMnnN7yv7infmRQNRxEk4Ha+MczUIq3cGlEOAIforjKUHzOMpfz
VC4oAGdOPDr0kWFHY9WBDvU3NbgSzZHLm3LbVeRSATXS5/slfcEjjIIpK2OULs3o
GLWJqiRF2EtqepP0J9JKBKX/c+bZv7b/cZMoV84NaF2J0WSfvSZcU84AYBScYwun
nOWmeA/hgqmnQTyGIsJMJgwITrZ9vderBfra0NAQox6OuzIVcu+00ZlZGkQP62BB
fu/QcwVKgbiK8pSTul95qbHLQjETswa11iIABs3udzP1faMjsSz+xQqJ7t7eWsR0
F4P5r3OdDiExQLJeKrGB1wgdYY7t/Yq0dz1f0mKcf95Pb75RMMXw8CJAeM+jdzeV
4qMBT3Pp75oa2BL70N7u4O8bmSX9Mh9IYPQyn0U/cg8MCzFEi1v2am8GoGzJ/N+b
f6FtFeuBSelEJnKla6SSxxNdfdVs5Dcfk5PhCM8ZqlmWztm5nGJQxUrJDAGEjmah
3up1udOWnT2chYTEypjIBvwwcFJAQJlcWq9ZKQb947nATi+VP/tN0FcJYS6AmOBy
zb8FpC9E/9lAa8rTC9wAzin/nA4h2H/2B7cqxyipDT3X5RMet9xHTNjXpn1UEwj8
tJHOm3ltF1KGI9ueK1tFVsLrHUWz/iYZ2ZDM3M5Fz3LZdW6kzvTKbjNAXD0ZMwIX
lKDK/dqB71E74RskBG233ZKKFD6sAWyvIp0dwErqUPoFaO9EjI4WIk48QHkVe1lU
JmdfHxvTj5g/8WzyNPPUVj7mMC81uMcVXSWBGrP1mog3bccZItuKiOAzTVyx2Xsb
VrGSa8mrH3cTm/iTyUzwdKTF0r7XBNJnH9CwDHPomSM6HvVCgcaLbrU63dt/TfTu
4tB8cbE/hAxCPtRda5EAWqjkBvjo7XBOIwwEyNroRGfTer9klDeZWtPpwexMOopV
M+vN9ACQkhoDY5i4Lh0RTCW7umiw/qH0mLdltW7TPsKov4rLejoz+s5H7cAQE6bG
le/wEX7fh6s4EhYxwo3+Of28iJe6wlEWHO+SNO18hlRo881MqB8VLMpFIYFHodaY
vryn7I5VGck22kXS2HmwOYV7CYPV+jnsDyztppS/rIOP9HaYOHUGWQV3Pkz86sFp
jV8M3hlQ0BLEpBoppvTzDaUsk8iKNyjGHOkrI62Z+1AcwoXiiQh//sarS8NEXB98
Xqd1CZiRGrNUFW/CfXAzhPWudiL7uWqHaOt3PNhps7/vlOi2TYo67X/aFP4FrSe+
DCqWDkNzRrTjru3JkUQx81x9qr9XHtrCnELYqypv7jCpNDvXlWYwPi9pXJC11HPE
7HPfXLFr+EVxFmdTsqspg8ozkVf4/Sf0vfVfb2hr2wV7yJy7h4iqEYoxO8FDqoAm
f9tvWU90UCD7rf0yr5kelVPMOEDHO5ApWgRCYGdYNt/NfbLE6np8rpDoOvnxKSrQ
vUVb3OzQSubQ++zmHLlPRbKEebsI1JWE0t3iRmoC1p4tHKVkPHIBQM7WyvZ+6AD3
hI9a3ngb0QQOtgxAKahkE7tW4rOX7MGZKOYvjUqYk/tLOed1qgUgo7DxfddyL9Ii
IJrtCovmSakc7Yk2xUsCYkyn7Bn+CIOvdpZ2xrINVj54gl8+uDXuigk5E6qRUekC
4oq3dwNX1CKp+WDVFULxLkrq2n3qKmy0rw4hcoZyVhrIHHgXO1reVmDTcq9FvbDh
fIeNJ2mpIf37G4X9cAyRv7yernrFMK7o144wJ/DBVwBlgAGtoHxhWIbu7lVpNR56
xXBTJm7brxgkGoCeW/KQkE1F1O/1g2LGzIQcxifnKsmx1B/zKonEEQOnVR8wbylX
gf0qgfKUem99Sxu6VKK9I4X1D7blRmfTORjnwby3KiDiGuTuplAuk/TVrZhZ9GkO
+W0JFW9kD6DTN5H34C9oNI13bMEANkxKZIbVWK+MQFuVm/C+dfFalNtahWz8eptB
pOcZ+yrPp5/zpXegnjfr767lHKTgQSlNCQqquEbV6f7RKjZQn2O8xLHqKqgyRG9d
GmtZtArhNKIttwpFmvQG7tbySXYAuH4x7Gq2ksBWb6PnojhIecd53D0KyPn2ieE8
l4bisLU8zGJ7MJNuB+IkzU9tSqnxVn6IwNhsSZGV9N3tgRcv8wsjUT6DmFaFtRBd
gEO3rxZtAksbepHWV6Pwb1yP081iFjO4CKKwdY5C8vpm77/VnvvwIgO/SxIijLr6
U4IZS9/zDbzOLKYF/5gGax8zPMzUFZftgZpCpci1/lRGfPNn6clgevaYhrNEMZkT
Eiw3wIcxldePyI5pNLmkssDZGAS8hn+GUftunyrddWBetglUyQE7L9gqcmwMJgGH
JjzvqYYqWwg3t7qkGFj8D6g02M2pswFqUeyi3vtjFlQAiHypT5y8OJ+MrZhRCJ70
0koKAUynfikrEUOzLoyNZg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TOCxd27O9Fsow1TFu/Qrsv8SY6EDJMI35Hzh/ZjfsDhxiZhUp2y0v7SX/qwyMxLs
YRsqR3X2cl8SCl3YpwcqIpDUD/LfQcje+YKoG2bD4FCaQrBn5O5Lmu5XRjdOBpGd
2y1lSFcK+Oehin910VKuL3uoURWfwnRFz20uVSOYQC4dmwRrWHZdfCKCvXhpCh83
3epBqHsG3kBBnCrcjCf9E9zwHgYII+G5tcfTZst8Ci8Bq8r2RprBamqaDPHYcjOn
I70tv3IjmhldNUiRDExzbUPW+hzpplsld/DjiLzsMj/MJR+8MahhzDb4qNgvDvtG
XdqPVkGbmdJJtkFCtEUidg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4880 )
`pragma protect data_block
hOF8Zx1uzK37cQDaC+UblTvJm2iP6IHsQnM0gt/8wECvBBktVQ7pETwx0LeVKCb+
wZWY4odTM5zFHXyFaeEf2qN217VIG3rSPqmJ6RjNNGsfbJB+9kHZTUcCBkbkS660
+I3d85EZfclwpyzkof7D6Q9Kbnd5/IorTch8ew/AoiMaowAJ3i/syfLc0E0seqlG
b7oU8tyz9fEDQ3SqmjRSIiD6kVl4chsKCrX58gxMWEs7FR3s8NcmsoDc2v4F224B
OJw+AmyhdGbUw1tzuk9nvkjCBEYs5znBIRFMxnbXOpqI7Ht2friTHkDu7fP173ui
TnnjQd6tadl8rr0/4AtI7OBelu0TQ9RphsgH9j6bVviHx9zGGkUvYz9H+Ef733Kt
v+wAVlr7T1Dyb0AQzKJkRPQ7tBE/JxSAFtxIX2B/0LFT2Idq4MKW7JlC7cBhzcPf
GZ59Q5W4umzzQWA3cRTzSURF6vh+5XAJro6pN+0xOGXa8mKo+NY4yAH70of70efr
MxSl5UKG8qgVJfc+wCAhczIxFYcPaRyeuApLSyjpbSiZW230g93MMKkAtZwjRTBk
O1lrmQZ2dtGseXMaibCPskCpg25ThXmbGJQxXdE+pJQdIUYtFuxcQCtNrz7sxQWL
bziMP+WDUs+lyTZ5EJzS58s1BP9E+BVIQpFV4bXwaLxP2gH2czYnBMnJebdSYmXn
Jj5+Lrl3lztryZYp8E/XsPSHALgJfobw/dFtHH8glK1GRFbeBVrQYTF1Hn5TEUv3
DFD6U2W6am085SiCezLFNMayr1/VgdpT/8p3lFryA3JeCQJRpM58LxEQRasxAv6B
Aysan5DSeZb7BZ2Jn4qO6GtJ0IpkOuTMvgY/WBv7sELoMzrnm32GjDHm5qOZePqb
Px/SoBqRTMNFfC1yjP/yFi++uMnoEmTHfx2lc39Bw/fFAVU+i8bPulyDhgu69KNB
tlVi+h8YeMWo7YXjG5WYzm0thmPLGDVs6NUndfCOQYrIbJBnzL8TKyxQXSovRfog
pfsajUoGhstbIkUTJH2BF3Yh1JOJsrk71ZH8y8oycldPQ+ayrk3xym0pbUHgN+xh
v2tClYY4NyjK3y0l1e2rFK4V2sMfMkY1unBstL+kIigEJL0LCf2IWypCeFt8wiku
yyreghR4H3zIsCv6hJKVLrbqch58+/q0yauEaeuq7xancLKzgJxN7+AE2mmkvaXP
zUwF26fS6ZpH+tm/z+duWm0zhyPzTB5hTextKAOnA0awLOXqeWgxs1PBGroasVx7
8TILaemJt5CIRUG8wW9+eNQuOXtMd/jl0zJUUqJF151do9TDNM8a+tDTlX9UVKaA
LtawF/RWuVVi1m5X4LMnzOhVz0nl6jQ5ZhO5SBdTzQLMK25AkLWY5nVfmaUIpCe3
4tKLVOEkp1dzcrgRK35Xby2j+seNydjnqQUIX0o/VIs7wBKvCXEXkyeDackAtgtM
i7KMk0KKmZAsxnxXAdkkX7M7JnMnXiGdk2SvWVCQLMm2U3LLf3NC65VYdq38Kqha
IyK0kQywZIhUq6lhGBYvBYIO9Emp88NvI3H9PrDZsnNAZLxxFq68r9+QSdYm3oCo
wCBFx6Vg/M6/nS4ZhHIu29vtejytZcTTBJgwHeab+u9WPPViJ4tM/8OlMpar3vZW
AQDEDH4xMVeul8wQIzFXJX8S7H0fD7E1kX/LOjK/saGSnQxW1F95OCI7PuzfFsJa
vpTNVPkPucWI448sYGSjN88Spc7D9m1wFRmszlL3yk8DfJI5h+1TP0wix9qqngRk
nSwphmnjoaRMm1BSQ3xmTOxsR4T/luoB78V3qlDECfdlqsvCtOctDn+Zv3lhDVbF
8Rga3JcrHSH2xi2FtHRmZJ6Qe5cxfVBrE1Dojn6XmvdH+3NKB6LvHsHqMKq27r/R
P3xWAxOusvBVaoO1bJeKT3fDikCIM2XHZeyJsBubssKeKlgZacHDGdS0i7IlE/uJ
OGRUJqBDMoGy4Z/5EuDnnVxjXW3ic4y82vOMWpI4kC9O/9rjLMDkwspNTvZ4rrQk
WYRwv85kQ9Ave6eqrvpq/Awj8WFcHMPEbRrLb+PAQ/Fq2Rl7rbVpgmtg0yTkPf3X
dDX5dFDPk5PR+PwO28YS7RnPcPVcu06HP+A1A3JbVPcEBggJpU2f9ckvl0jJwgoI
mUSSQbXKIvJhbMxMjVOYQ6ZH5LQH+zpQQODDdxlFPcp1/EWg8P/8TutErhqQllmk
0ssxujb5MKtVSUSmxNjIqMQApslGlxSqqHYeXvAhRGJYH4RAgru0AHBG/9oDLRmf
aM5vrzuknFQy3LxQCAZNUqdxkXNXvDo5PKHt+7TYKfMCFuf6MuVJIBpLft0EO6Jt
85Lis66HnB4uIpOVOkC8H1FcHo3vDnl16op/REY5LOoQArjjz+/E1o9SFmKZVerd
sCwO0vyKAdeheingRR2e/9BcXKCWbA/4l1WE+vpw7NbadPWyVJHTBbw1LlgSE8I+
E773vdoY3we/WwFeXo7alOynFV6o2t4qM7ehfy8vNd6az46PvhRuCL+VZTsSe1dR
XiMLNq4b89Y6xyZvC7GNIZELqIBEX0FzkMpTPB9pndaSN14HyBgVTANAZ1Gszilf
gQf+1jZbYdDbN4ErycYbcpbYF1j8c5HFjzOUBb6IRNcjd8RVTAeMztlS4P7lZMLu
O2OItJFu/x1hf7gZTqgD0i5XCJu3DrnbP7rmL9Wohx53jYO2M3Q8f1VAkuekZVmJ
taoLtPnq9kNCFagDy0Cz+pySZ1zaIuGO0mRmKpx4SXim4fHh59nYiZhvOVyKbGgG
YEAJa53Rk8hd8KM/ZqK8nLLrrxhlL7kG4a3gIBYDmbKl0K/Z/QHhBVpQ0aifF1wd
1UZSEk9tRRaI9NCaErPgLu/bnw5JCo//jA8keHl7BqivBkx2NoQriDNrHKaCNY4O
o+xZ6Pc0ri566QjCH6FoWA2WwV6/P+SdXiZDjE/5xuiobTpA6swCSbiOatNJZQj1
s1rHk9tjuTme5q8JpKHufXtcFXZmdfssBisU2ekxLXbhPKfWTDCSnTV51GljbYjm
k6wJi7lA3fokot4kFE+SE8lInDf4laYRnvvP/QvPY41XQBQRbhtmIyaFwuozKihZ
668YtValmTecXCH3orYmaZa221VtvU+czr7TdmZqpC0ebIXlqN3UsGoMbpjh74bB
vZ50oQTdjdNcVwvAvr4SSqe0LcBNKekaOSVVFMeJH8OxE6DSiWzTvnNYE80uK4f+
g03rhRRKwrqTzyt0IbyyCaw0NPWHvDCskhPfqqu2Qx7uDkyOoeH0ppI/Srt9e5Jt
4sNAJKFQDk+el2L0yINJEd5miZg8RCD9xtbi1HRZtIyuUZUuu2KACn+5JFwpHmVO
AM/E5Sl3FkC3kfiMeXd7gUAtO7HLK35csnNe6d2zS2Z5/qIKG3AhO+SkkPDbU6rm
MmuMAx1HhqUjSqloC3LjPBBVMun1AO/NAGaUOPIv5Q0xhYOFct2tMzotbZmFihFZ
xzxt8vghAJqdbqRknb6jzHYotRAeFYa2e1sZe/cZQh+ecgzQ1OtZSrwxHo73gMb9
79qP4ZGB3wcCcHacFNLcKDu7IcgNhLH20c0FwQ/A+kIdy9aHFtMAExMv9ljeap8y
mUNaJe8sWajZ7JZboo67l6mGsFUgH0+fjXxH0IyG+SWAUPdIZeRfwExKMUTjlzxZ
iTPwlrETFnxFQmaWh7tlmWlpZLhA+OJawkxnus7Khih4dGc3PwylVfsdSFfe+wve
woxojElCSL/nw4Jc+g2mAYIATvlgvsU5rCeLIVXv5kkOwFNMWWcq36MD5+iPHPK1
QwM2y2ExhvieHfyu4c9kEqIz1VYBX2HXFRs1in2uRJA6jOQ9l8+gCUxWMcSLUXd8
NMnmqTW5j92hjbx/gHdNDGAw58zeq8GQrjgud6mmd8HZ4LMA6aRx5xk9TjNleL05
4WaLawPS3Pc1tCBO+SIlbMqsEBTmlFB/cU6UihX/tGxzMZBiD/m5BCbYDtyMGA9Z
3GOEAgstMbbaBznMVqi/Qa0Lnc9Jifvft1IIa2fll3byEYxGK1pTrLhuPNoMoVsN
v+hfIOS7F6lxa1cjm5aLPeBNW23PhHHNuL6igdqLVkCZDrQEM2d3Oo9ARz4Ej9lh
jJzJrDVIXCSdUib2lmk1DIarTPD864SSvlEplrNrFr+AKGjon9cWDAgP2JxPrsqU
qAyNJQ5UYJGLPqBp/z+FogwB3ReKaPG0TuMBHt0SQlJERmIsNBIxGiDXW5It0Vvv
cHa5pxYlaEn6Wz+iCpRXnwR32WPto1LktIikIw8N/qQjFrFNpUYwhk40XMMAAF1+
Rspw2c72MDsD7tR41qXe5wtAumP9LPiuXvpKwZWeSZ66ZqQevTmbyqcfwdg0kX3D
Un4zOlKHgjLUNxj8q40R0itMVXkVOU0sstflN3vpDeA1TZtk2zX4q2oefJsHnO/0
dBaCCvsoRo6trV29lzz3x5QnuS6Rm6Ugkro/meFPSON3cOQMxGlpQbvBYvQ8JigY
wf1us97BtDC134PDIEra31jt5fztQBlCB+bEs+6qQKj9xooHDIHVprXRZj61mP7K
c+RYIUSs/7tGni/x6X+b2PGpkQWLk93PlK5ePKlsuL/XX3RIUunW24WPJ+/eXqT8
LECQeGD1XjDoH/5oiA3qa+/6YPdpSwHQs+ggeMRSnYWguBTZHqajm5njQ03m4F4y
GuRTJsGhiRwzKnKgK0CgzgfILpW1yZCOCKmu4N39v0w5dn31qOxQHybv9zClL/wD
P1+G9R82TUadBWtzZ3g5gvk2vwRm3m89cOe4DEPUWSj7E9GrcMDbvnEG3G2Bppgl
d2x/WwyWokqCUh159GN2anyAXiM/gC/AFuprpdBnK8+MV3p17aVj9C7hWO9srAqf
fMSfQfujPygghgc4+Vc2YZ76xbi4Asox4ACA8BvVJ9FyXDoc7Z6PlbZJWeXwrfpF
AnYmDosuKzhaZqRqGqFOg63HTW5V3NxIWqd+GrX5FnaBXUmC3d5ztzJ2NdEa9Ey0
GSR/A4B+YqY9NrYtDlwdlkt6PvTqIA1XMmzb9CwgB91az4XoJDAyRb656aUaLDQw
vHIIcdYNBkkVgSnFCtMBszD39iNu3mtX7OZ0+3ytRZeP6gdYOoBj/vXsM2uD/Fw5
6Xw5FDHPyxXmW/toBJeGWO2Txx+vkBPnoQpG9g6IzVk6euO3332nfgyhWVCw/ZVS
jLtemlwVEUE08U8Juk1taU1dLtPHp3OKfR0xp62v0HVqWDDRYyHrb+wuyxnE8vrM
VvscWcV40dudZM8si7tRo+x9l5fA0xNy03JOSAkZzDKCBNwnUUFfZJaciUCNsQ44
m0oVuwHO0WmevbLV9vb6eNLUOj009Ws3OCeqcNxH/RJe+iLeqzD1Kt5/f+pi3GV2
AkjOVrdjacIRoREXlWZNzAqR4+krNPndA++zkHSDyXJEKvI0nz3t/qq/3yaV8LIr
Guwj89B8rRhu+ELnaT8eQ4qCVR/okmoKQPw2VMxU4/lldrJj8Gm4EcOqxfkBs6OF
1VWLXyPCG04nqTYfOVW988Nob4s20obL+D46OArWZdKF1qsYBaI2yfbqob8UmRQP
T7E4EOOmNR819zlPYEJLs6g2oZqdSFPPCT7LJQLyFATKis8d9zCCDPUxw0tgglxH
JSL93LulbVRYV3J+fe5SB5oaLkj+KIbagkfpBFnXZXhsfyAGpgkIyODGhH7zKv56
7ZIfzJ9I/BxRCd//annVLJDXciDcRHdfOtvtC4sN7gHyCxcXXwSOnIRMmSXgKHxm
/ZnOtpyfRyHLWqBgMdmHSl3tYNv1JQDTCqahutnW4vco9ITlIoAkph14M8/6fgWp
T0MtK8nvvswR6SiOY1SqlxEBCr4fdS/L7RsxCuBpWJGj6fNayopjRvSMgZOteawV
55OZXmK0FtcpC1cnprU2yqFSNPtuYtnWx1AEZTwO7YEQR/hukc6ibbTdtaLXpIn2
ErSozZwpCqes2gj7VhYfOPu91jleaphCtue6zDGRPJG9kDg1deL246dynT9H2IDz
reVoSKtMNVhXoCFwyov3++SorCCepGpuAoiPKe1XUQGcUwoWJdGwZ0/TYoO99kid
7Qzvy5tPYAhx+wZwH60DmPFC5kl0Q5xqtV0wZFw4j9dDb6CArMi3FJJiNOisUpwE
tpvGeJtLWNON5JDpN4uwYuMBj1MZnAtXouQg4Lli1oM7T+khx/7R18sPOSXlQJ5v
0gnE0EkeGm/583Du5VznYK/0RgpQ16qcuwhDxG0ZlTscMtff84wEgOqdgRAq17Ck
34mDhU+IDun5MquhV81+nNNsqRdv3LVj+OonjHBUHv01Bq2p9dAfZnDeUoSQVxg7
V0YfrZvNcT00JtROkMtSp34isYVKwI2F8N7ojXx4bVnb+MtT7U7QFsloY+DjgibQ
pPr7Qk/UEgwGyuFRjmIZHz4a/pTc6hbNbKhsNcLqhrc=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Dw4b/4JV88/miqhkwU79lrjVXUcR4cFTNadfcT0LAPb+jg1YxP1v1335/rBiTNFP
WcoHILXR9DJwM5E5sT9AVKvIYH96K773JTZhAR+h7ON0kqrkAaPzyiLtq5mW6Okw
ZbLo913aLbwBgadQkvceCVzTBZN4TQ6yIt5+zvmiwG3YsI8iCYI1MAsoM5nEi8mw
rviXTlyy6+QwTceYHrjRI4Jyu1eD69Dhs5pS3MXhO6+AIMnJQ7c5WxDCAjlgsKHX
8inPRLFktZObNeEVtSK+JTyA5OuWYmzoF+mRHFWc16m8jXscz61jjpED9H46O/Gy
Px2Z/cX0eEuY7U73tv6eCA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8992 )
`pragma protect data_block
3fVzupC9LnYFG1EKM2Q5nOLHBg3hnWn2l7SrMf9+Mnp/Ic1eaWvwAFR3fbqE4jdw
Z8eoP/dV8gcypVoPa9Avp7FT0zLtZlzOXr0C7Niclmg3QSU+Qkqp/0dAJBGKrZjK
jFm1SjieQdLSuxwGcTuW8MjV+4bFEQH8xW2AuzQ0JDMrC3U73WodFG8KpS09Izsy
glbclDn9EI6EWvbBK92L8MJIqlHGrCuzGMoJUsO9uksRQq/4nxxr1wHU4Tyf8DAI
OYTiCZ7S1wczvxtP6yfN/M8Nu9A9sM+IYAiwVTX5aS5C6XSBDNoENff7ke4ot+b4
rD7qZHXI/c8rbq+QPBUVGaXl9PipQVoEs/Is2oi7Hs4kFdzV8M4vNRxzZoGrrhA7
ALENdlPT9JVxTG8uXxRVFh/fbButPh35pwkgEdgivlBVZNqAyCyHHnEDsI912qJV
wEgIzvVX5iuWkpSjpgS/nbIipIW0jC0PDdq0GKO9QcLT00Sq0cdPiI32Uygc9ac8
lembJ0kUSNQtqw6gmVZwyqGTJ/zPwPq3dSnyLkWXkcm7cHIInPbxXXGxmfak/GSS
mCQyjmGDtA5df0lpiqchcmPULTWkLYf9AuuWAJajATWl80qMsG8g11y+DRLuHZVn
x3mpF4v3PPf3sgbQjFHvSoGxYSZaKwZl4Jw1DlSCwOMoPq24pli50Sev8zmlV3Ba
KSwtoeBfUpPloh4Ip3PUr9O1m0ElNDUC/VUmCpLGEi8bsC/7o4FzNUfCAbkFIEgo
c2YjgEHaDUICuSCKPQ2k/yNdqNYAcYg0AU6zw2uA9Kk1jS9jD1MsscH/y0eHphv1
F8lGY0pkx8UzV6RYdLmTCjtrsZm/KUu5sdNqnw9KOu3qFHNxgKVZHBZUKtGF4YZx
OByJiLUWJK7RIWGhhdUcyaDSfLjRE5rTXYeFQD0NIexifTYRk9YiJ/x8dcBH49uj
cAOAJ62vubTxy2e35oKDoVOH6LFI+V5fiosUzoT5XHrodiRwUAc0t+r4bLxiTJFS
xdm5k9pygLSPmSLy/qzDSM60mGjR+1zwZ5OdX3fieRY56iNAvi8eCMhjroUQe6ZD
fiD/efeAbfybXe9Nwam2UQ/eDN2qFABmIPGnbZGfSDCvrOVPvklfp7G5LOj3nHEX
QJMTyTPQV10OJpQnP/cMK5q3XkNTrb/H4g+oGuGbWuDERanAvWOQZeu5kkUxSpuN
X60M26QP1jKHaFP/P0b3jnSA1WmYm+j4tmK4l0tawbup1PZTcHb37CTdqxqdN09C
+wm/PyGFqkoM8svHjDCLyed7eE2hScMhza9l23/QsN1JwHypERZPhq6sSomB2g1t
A0iKvBe2fFLBZTSP3UKmauh3Pxtq8FuQNS2t0LCLk2mvi4tAR16xVMYWNBZ1mYxE
qt+nRUMVIftTazE6hfooRRtTNU/v3hIuss9nQ3b8NHhdmHMHJpFUJMV4fgNJUUW3
2Z8NQHOHmdhvh0tpjBORSUjBs9rbvx+Gu2QW4ubqJ1VlE0JqBa/iSBFYGioGNsP5
gxRmEH1Ibosc2PIiZzUwG7d0ju9fUlHFfGWhbLwzq8iYgniSCWtE3MV6rsFhBjbM
j6ExTVgnWkVz0So19VCpMk8Me6KwcGo42lFqLE+hxgBB7Qo80AI/+xDj9VQgi/KE
17dUrUWqeJuwcn8OT1+QlK59dmmD14Ln+HliCr7V8J0qbaPUdexiPf7mOVsyUFbG
QhnoGRH53XsrHJnzxfGvjiAL0fGa6qrgX35a+HWnkRNUGQ61t5RbuChUnV1aSomq
sEFObHJLKwxiiqMIcv9wRZ0g1Gn++0Bg0BGLZ7UZypzSV1+BHo3IrQ/DC7nyokbG
d1RG93NCpnqfoh9qE6N3DRkSZkTOkBwl8S+qxRtdqxMmWoZY5Li0dF1F+1UjzWie
vtVxd054ZHpezMFnJkHCsGsT4BGjwcT0c+6VwdiZDGqvMEcbdrbSUnoBNHFl/HtA
WBx62n8Am8D6/ezi+huEeVKNMEYcT0Dmepcxw7vf04Bu3UhXf3gcKnvkKjWbe9JA
pqORXPi56RqjAdhUx3i4Vx3fK/mOSlSOhoqV63h19S7wmAm+kuTQqtfNDaxPf9bF
/95GvmYpXElvzbAq6NcA1ynne4XRkQJVz1byqRE3kkwRpg3EAKingLrNAp7oOApe
7CdFVFatNmhYBbGzTBZjOFItkk2hSS7ypve+f3vX5+A74ui3zYVlj3wBwhZrDtBk
jFubYffP79MFjr128xIOdn502Aevb7CGUm0Jw4fvc9Lw8q9KHL1dgibB9Y09pSMU
7mr0IXFgJPTi90OJ6yd0K6Dy5aQAI69gHkErRAqffDNbb4nIa63JXChH4rj1JQwg
7kPolfz7+QN/vkB6KemPKEHG8aI0TqnCqJ7yXhDgNRE8fL64wygKuiv/d3BehvEO
j+FlXfuImg9gg1uOwnDZ4sIZt+5NfkmMiO96lgtjSQGD4tHVNf7++U8b2OQR7oPp
1ED6JPFlsMfrVq5C8tZIYpOjJJ4GmaeNr1X/0Gp1PutJOaDxVonxxosXwYl9ZOCE
9leW1mr7X3uC4iAKjDdgXJk3bcamaVJQWWXMChHjgbCXCOkPve0lA7meCuFEd425
TEEB/4/2MOoGko7IF6Hsyib2cCjBCafhPUq0CD5nL9hDv33p1w1Mt4UruJesKSVw
+TxUoiTOhI+S0Q0IjWRnsYCn1Y7EZYO4I8QMECDy5GuhT+pzjS7ttc4K/RuzIDh3
zh60meMVniHRmwE6byRFBwZ4dhI4IjCBx63JdqdmfnLQ8BvxsTUhdtFhkQpVl1Qe
C3D7fAfAuAVXNyXrBnHivOodjjKHVPOQF69TEQ0aSuLFm2OK5rUmWHLr5dGe8bhd
DCqDCvfA7OIaZbl2hx2Ye7Lw1x3gi8shQAPkt7OLlpirsD4rDUI4qXjqtMHrc2zi
EjoDPmZU6qRnPDDcU6n8yOZNuPv1b6IKCkp3w5ExeaiXzz7rqL/UQqlGpPAtB8nG
qhxp4SsiatTL0mdf9Lqfh7nH1oE15PA4BbuSChoe/cPKEPL+5dZ+x32+oJNoQhzq
Q+5i5Ps1GHo+gQZFcjkRmXpqzU4bU7wWiw9gVlk4Y/tI9bhfUfJieD7Og0J1TMJi
YiyruePpgJE4fgSnFsQAyZYP2q7IjuHBwt2FZGPNw8k0Zj2NeVbWcvGBHfCie6OZ
b7cK4jDdeVOUP+yzu1heYWYkL6HPZ7R7Yl/TXT0DurtgD6GrFhO3vwtcjzZPbzNC
kmjAnUcsCtY0YF8n/RSzjpyiu3SKIiDWKFrgEubwGB2FSzBT33O8Ni+meqXQ/bFj
sobBC2iQCoDyLj6fb4BNi3Gtc6/f0sNTob16MAv0WguTecmesDN8rc4JQxYSRFgd
O7eO4tTPPqiUDrNtVQyFa0VDMzUnFV+tB6w133hPEzdbaF83M39xi3eb0/C2OEVG
A2+cVSh/CnmCgc/bHEvOGvwYzKGIfi+CWOpjAwxIomdPAlbbfzEH4urJiZvImdCn
yq1r8frEKh4eTKOnyeDVnpk4Pl4Pb1kdDGoBCAq39VokjboR37mXc9abeI9at61Q
09PZAt/vEnI9gN/GE7MVHLmrEVWO+DRHT86SN7xoxRVWjYCR7OKH6ipHldzUR+6r
ldyETzruIQw+qpkPNCHjCeR4YuucqHhHhzDbdy6+33GXdbA+QV3cNK4zfUTfTP/T
QA1P3BQqLkPOvQTc483Bg+kjP6PCJwoXywWtLlL94RC7MRJmboinbBXq3WuTbxxP
jZAmbJW9/AgRXDPOqrDeKYGvefMMecLewaIh4poAZJqBxdo4TQiPdgZ1Nb1mkGp1
x1K3Ppg297VVX6cFsZH/fR9p3Q9pb38zEGoLF5gf7kAqb+JVgjREUweyG9TVb0MJ
txWIBZDJCOmqdvdePSRtARLnJxRVlNmCJ5iL1Kvk5H+YnxMQaof+8DpcyweaoW06
mwfjkaEMD1I9pc66kWbygr94yE0+U1PITUSG2uR84IDdTvMVY0WCiVuJiRD8HUiT
WT39+6ngW+zVxPtIseGEgbLP0XvGaVBVMUhI3Ls5ig1x6XaFhl27Pbz48PleDCf1
ORksZkK5wtWLG32RkLLOZiSZnOfvHiGZBQ2NPkpVFQE36AgKUgVyIBboBnTbJHtk
4iIAIgu0kszZuVqQgkeovR0eHK37QsWZYBUIyxzxwfbk7hodV6LMhZViskvJe/Fw
g9UMdVW7FX16oxtzvfT7Zq3WhOFFS5J5hVB+Bx3KgVnz+fuTdASie25hF4q79mQU
bJm4QvXJRalsvyw0AKJJdkc2phzdJ71aCA/5rWUIRPjQyDhJTneg9gBz6LR69KgX
Dvs/+dOOwdxxNrS0NZqr/Wt1YepS60sBeedogWZKise+d3LX+9e5LqQXeZ6qyMrt
mG7IhxFF3zyXTJBACvFTk23ukpI7xjV3bcYb5v5gXaZYcmTYyQ3uko7mhrY4Jh9Z
ukgJGK/eDj977qbCo7hmLGQiMNF71hObA11Z0PSn9TQBoKDkHt4OEtgNVG9oaSkN
ERtWu644lmoa5I1FHWRxP/TWiGaTucQG77h9uDK78gf1l15PKqIBAEQrltRp8eZu
NNwqzO9TWoT11hIlbVwPLrmXx/oHaxMyjwol/04OZ6S9HM1Vlgk/hdG5xAo3aJgW
lFrlFDw/tg1gdG5naLG6tuaDIB5FEBEkGPCgutq/lSj0Xv8OHnwXqygqWHzc6Yq/
aHExqMeT1OvzLwRU4iBjerDb4TMpiIZ0zoxMznf4uU7c8SsM451eaqbJIlVdHLMU
iwmrUeRdlw4YOWZJDR2ixWoKPcmOf/m8et0Z04q1HTXrqR6VgncDA6wmi8fW8jwz
nnsA5Hv8CldoTcKXgIUNiPHpidIcrmo8Lghup5XyqDslPcZS/bJvFD+7WmzhBHhg
FiTrDPzN1gxMB1c5BmovCN0LNySrmhTGgjUEZs7p5w5qlJQxH1kPVBNxpn4tfb24
aAtXAp0Pu+jyv2zYG7nCDZh3mxu2ZR49cuMuBWAgdWMCPP41uZmSiLCy6Y/qT78t
FSipxRw61I8RKZzbaALhVJcJvvRiBN6U+VR+EkzD//DLrhdrKWpBkPYwZLrFxrHi
O1sFMpPcFHxTRP57WQ/pYoFol+J4YaDb13Cyr47YsPSCkMJrhPw1vFwOxOJc/fYM
EOMi3cp1ZuoaRGUpT1/xCUwRRwKQuoRqhyU3VD9zjBT5LniumtGrQe3S/fY/abB0
+FCE3PeOJx5f8NZJyqPcfLGhLrNMS1aXc7JJCHAmiNe0vc5H4XgthTgqx2VekPa3
v+H7LbbNhuT+gEWmjJrmQoC3+3FilgkZiuWvnY3CH85WvXAP9jWrA6I08WL+cg1P
g74Z+pd3sVM2hTTh2pmvaT4ltGuJrozNp967Q4urBW4LxpRqLNUj5W42xQGgCvPp
oz0JYzkdXUrcDxmYeZdSLmLxKzBGP/ZViiRPES/1PklsDVKdJ24YF+EYO9G3WtoY
a4y9z2ukm7PFoW4tBaVxcAVtgVq6zrh6Z1WmpjBNlw7pmky60F/kN/DDG1q0jsUk
TSLMMZgSoKExiQq/jaFp8Ddrr2SwDLp0MHQIdyqupXrquNAWuFyO3jfjUc3G5qN4
xG7PTAP4Os5rKm5j+fENwyp6DdAexAxLRjQZHSBFgVHfI3MkgOGYkUWey3iF7VEq
8/owuB1CsubaNfQb5tTA+tSVbimmKFP4yXYv6NoOSKyv/54Gp0lN+xs7ocLN3WND
yhs0zQ1OfZlsQUm4awVeoHjHjGo019F+HCesZqdWOwhmT4ILbHUYfrLuV112QiUo
XpjRxBijUeZjQ22MAuZOtwwBW8w7BqCsvmQM6gCdsxW3g3otfv+EQx2/oBUxxX07
cIe3IPP8Z5YeSpo5C3p2/ErwEAXr8lNAD/3zHT9F0AWLbt9uvvZgpyoL+Ai0MlzV
qoJzS2ijuYGoGNU9CykBVEyKtlWcLtdY0RwoXMrTgdnIdOKVCfOLiVVOTKsbiwe5
V1f8aPIEZzy52PKY/v2tcRIWLjSIgrljbWof8sbdnsnPjyoMctL0v+z6Wn6MvvkO
fNq1E7kLxkHmhIRfM37zOtL9c5/4Kx+eHfEqJcehwDmlvNr8fLAMqd42ROa4/X8B
6BtWVAN0uIQATw6BD4Yd3PckKCggaMoXnETFM4q87GVxO3qMY1dZCe34JfT0uYOj
wlqhH/ufpZWM6nnyKxYPCgvZcZvQyjfumNnsdTyz+UUjBEseER08bzL25UtJQdhH
+EizOwNivUMDg6zctCGBEvQoF7lFSaofJ50a1viP8y8SBs934M88HXW46R8tC4aM
dPeCG+rm0kxSOGG9SnnWitDLRPCUAYtIolWH/u/3EOyw0dS+uKRycdPb75FXyLwE
4LbHmJdYxiFF4VPKbN7xDXanLsJWHH1KD+odNqRFV21PnCSC53jnb6SnXE2jwu1w
GccMpE4rj7g5xPcwcFJu5pCgNN6CjXI6UGfFPKKMJqPz30JeN1N6x27PGPUkLFaI
vghs4NFsRBR61bdU/+BV6l+0dhYGxaqA+qVtHclcls7lhovCTzzbaMMe75jmoah1
VEu+ICZgWcUsNrLH/REAJeXGkDLlUEV3mVhCRWFdrSW50s4Bo/gJ1S32j2swWlWr
i16NmN32lmjX+vTFAKw2XxCsspD/S/TRIoWUtjoPyaq/3B7jUrzzehD2cr+BTmoV
/svxrETA5oEVnbkvYzcaPSqVk7Em8Ezx77vJOiY/pomJZW2kHL3ioDw2Nn2Y7qhp
jCjyTvwQbcPs6NuHcjqgdNs29PQEutlJcrE2nMyoruwHPfHgI7gFO6YZZyhLRZev
LFcs0Q4bB7zvoN/+5q8Q/hzpm6bEogS9YymDUFSFVGD1cPA7U7PNCCABGnLNe4+N
7Etp5M9enPoXS60l9K4EOSGtS7TI3yWMFKi1DH7NkxS1dcrK2PKGSCGJOspR6Gbz
f9R4q03Tgx0XJsRM9WR1MwxIBSFWFHdNfMCGDpggLMRn/SepASDK37fnnpLlyz77
4luaZXCjlsLlJ6B5q49BHqpF8w4dxepLyfXAxmtNiT93e2LWUxG1f6Rrb8vxh/ZE
h3qXLef15bnN2V1eBllfkM3zren8mFvFVyOZaDgLEkKOrbyQxA27wmQlGffb8wl8
cYFBki3WT4UTiphMyo/qiomXXtrBUy/A6uR5tAHL/l1Yx7BqlwNZtJHyXS5wRwS3
NI+9/ntcLVD6kggb2PNcc9WmFRU0dGjEagggO+kTRDHO/bdc9fhob0zmSNGe55dL
UFhx54GLf5zPXMQcHLIJ3u5dw3q8ZK7FN7JW6ZWrKUbH+vZZyOMIvnZhu/97/3DJ
WgGhrJW4etr/zFV5n+WRYzZyPP7GiJpvgkS+o4ecKbucM2wNFzct5o9A0+bUa93B
mU4utlzV9IZwODlg0MgXn0M/u4cmiA9gda2PXaC3KFmTKeVtwCg0bzwesveHfXfL
SMlCAkfPJIDKi3/K8kj3G/2RTVSadK1c1GbwCZ816t011JGN8kW4p6Jcdkta/Yw1
J/kwzlrroGEwI0wH0TFQw2naXfkZQ7TrHGgkQQ8pryCh0uzkFXj7tKN+pQfzkQDq
8CdTYenKXFne6nm1qKRNwKh95Dvvz/geJlFVzVODNU6xMpj8y4pkRVE+DnOPejJM
i9jiTH3aAqHlWtqYMV2/4eyUQRRcV0oafWeqORdYTkyYnPt5R6+KuGYgP4Dwr8/A
5StY3Ca71dj/FHj2/bTuP/7H3/YKV7ueyGujc1e3U+67ZhHFN6Fwu94pOwXdHepZ
JqjgpTKEYAzkTHLLm/FutVGBCPm2MaYtRRUbnPu0+TGB2g5crt8o2l7n/+wiD9xu
SGyH529I6b59y5CuwUh3/Nk3m9EBfeZ5wF+xjPeNTAMB58MhyXtMAaexnl+CZuF+
Syr/2kJGMm6tQGb9r5ZSeA0HvwHnIBuvZCa79AAxnelRMvuSudnkt6EYTXAOctR7
zqXcUFagJ9xn84LjSx9YXs70O8gPRSB2CcKRT9IWbK/W91WHb2en8e8qi88BJzpz
brcGhhc/yvT58ZyEZ3J5RRaXgbqYZKDOh0U5UtSllOnosDB+fZ281JH582hyaT2w
PkyJ8XhEzxxeM96npX11G/3a4tZZmODmZiZFMvscAM2SfJ9bm0yf2q58MRuEVVvO
/eC5riBe5J7dYOXQq5QxMJYG9yEeJMAJxzfaKyKwzI3uexwMGQLX3Fsut4TmOoOl
TZFUFxYW/GkF2Jx6SccBZnKfGc1TUCGKGCVwOMvD2pSoHSCIPx2Wkx3SJggv0wnW
3LHbD6KFPW8y3p7fPhHgksbzSm1RfvPHkdSGgwQs7KhceZjOrc+lbFvoFbpmjhtL
b5oG/eRLNy6jpDERtGDmvqzxd3Iui9zgyrBk0qXQPxjkGSHPe1uoPrCbMp2Tb8l6
ZeMg/CnLWwnPW5aZKRhv/sLXR+KVlg4jbujY8dj4FIosLznPklJeTHlTObBkAmLr
DokZo1tDB3gcrRkDaTRm8flNu83HywrfpN3gVVu+8bTou0b0Ke2VrOCeU+QQHH+z
iGE/AOUBTu0Oul4B4H2t148Kg8cRywuFpeGv4hmq/hzplpnJmFBsb56aBhRkglUg
/38iyZe+7YsAPE6P1EXkxOg5LZJGyzt7TyP1d/VxBLrJ+dwnGl8W/I471XagnCob
lUlzWQ1HIvE5eL0AHY8JV33M3VeHtNA1LNTEtMxAIlW+TMLfw/XHlAMTvESafE2J
ouRzdtIpaCn4dTt9hn2D7iZijowFTH7lfXWoSwc8ehVcJIRCJXMePEMbb+t7wtEE
qJkW9+8w7Yqh7M9FbKrQzDVkoQ8H/rhkzQ9DYR/Fq6YUwKCVLhURYFGPOp4ivTr2
zLkNo9hWDYh0NDxrxOi+el2HnT/ERZVvYZJZGPwUkR/90X1yFtRXrAH8TK73HdOE
PNYbAG9vt9vJLFwFGKF3dThPG8AAErhQ8ZnATTiTgkea5BpVfAxG/abp6zVz+COP
GXedgPfFdXky1R8u4AdypbE14rdUGUcV8NywHD96sP6l+sCQhIcztKIjZ+Jug2et
gHoJFznYODJZeR881wJ1NQt3kkYrKn41ElGFofR9yoCrirpzzlEmq4JFZUP2NxX6
kVNSzPY5FCQTE45Fm/dW+43aElIvjSjLIGzqcC5ljdwoCs12FMSotcn5pjVOZCzi
gSy5lFRGkwFBw0kzHw8NB8UgXZZbS0+kp4tNZN4WB7BB6ZKZ0wBvuxqaueMiR3Yd
0VdORQ3hjWS5eDwcNY8ue+J5LQShjha5nZ6rmMAhYZLHMUNX2lEf+5isPXssdh+0
TuDPTS8sGo8o/hFSeL+fwtVQzGgA756M+jjyaoq0w3yYQ8vwXMpFWBolg7cHkupX
3nWALMqYKCaR457nJzGtoxB/sti791WC3xtOc2N0oujEpsI12kXSyRfrxkNXA7Nh
50Si+OaTtYg34avANHJgZz4wapiiMgdsr2NJXO8s3lSY1OYLfubokc5Aco69z1f7
Ob4xV1r1If4rcbXVmVskrVF2oyAD0qGjB34xkbpfI5RXqKQkTSbDkU9QdlDgMvCC
9Fe9muPVWNU6/9bvKcyyaG0ZwYcQYts731q6UF3s0m5wo4s7Prj6IpVOtmXgbv1c
GAEfTlxWrNT3yfi6r+8BHK3t3OLlXs6MVoJX1STx/ME2yDmwlebi5nPkmrwTPXXS
jJ4X2cQrVRb2I4RAiJMh93SLRsUZPqzR/9XGBE9pYTemQt4Q6LHE+EDFneBXD48Q
Cda8O+slxpMrTL4Pcff7fNKdDbn9fw3enHB5rA0ZbOOlhPM6GCfgahSF5WNufHtH
Vj1fdfiKIiY1iH05NpL3Fxdb2ltgYAr2GuQKemh76MUIPcVS7q5R/io0v33Ns1HY
e1BpAjeycQSHSDGpPm0gJQAej9KteRsvi75qVbcKUVPRMwpdvSOesuCJlfg+MQUw
Wus5TfHa8Dfw7h70Vyd90WuS5hIVZRlDwXt71/DuHq+6BZdR77WC84qMp61dqegQ
OYBGoBQiwdvPLnlAl3RwGwuABf+UqfSWvtxGXPpZt5VhcJQNYtqXHem7sHBbmM52
6iuTGErBbE55AbR0lpBKKw5/mswy3mKPWU17EOSoDr2PQbGhOBIzpFlOaNDIh/wy
QLeRzxCTJU2MYDX8uQod+LTgvZA1ulA73LHY1BXTNHDf74l3sdWHd/2xcsUGYFkT
/vDlMH3TSH67c9c8dL0KtFbhxBwv6ne2l0Zuf1F35tJvzTBhwGiFLlp6i2Hdzbwh
8MNkBbOME39chKVI89RlwzXDoLwQUjHQZscHyn+VLVmlwFP6yu8uSF1mGznBNDCA
w5ZQuEBeYUzKQwZV+r5NptxnRf56HOfUp6UOf1FPlR+JQtjcySLm/uyHUJz8iFwU
fWIXsWttgMrBUigwjZlucRTWVBaj56+95vZgMLxR1ard1ms1oFDtxH0vz4eVHugu
uEuCGRuUfm1spO6WlltTN8NKBLvloiElZE1k7JD7/Jy/E3oo2CuxY6Ee+qypzyVj
hQ1Unyj/4JSd2v2xFi90czpZsDFmrkf2ZpZXAGek6bcHynwr985O/Ye8EzgO5A5b
36ry6ss2jz4EnnRRQ8ky1CqozSiohTbkKikc7GeWVYWeJ5+Pvm4qYFhAJDP+G2KF
2vHXkvwbFZUKImnw/W1sPCQ8EcYfjHMDbyyWw86owKnyG3XMzB6ZGcs8pV4MjHXX
OpZti6lfyiIbC0bKsIxvDBgoLc07Pt/nF/k/fEemj3PkzyJ4pWGool8CR/+yqthG
zG0ksxeRBVLzS1sc5WKmUNaAFgphm+BAfgUfqi2wMHB+vLlh4LizGn+X7YggwAUB
Z/EvCblM6KHgLkzSn3rNf6XRP9PZgk/isitDUSDeFDN2WytAqcmrhPU1UcJ7Tys6
tzfRqe6ImkXic7F+dkOVIdsMTCFkSMfwQH4vcfJ8CCiOEwaRSy4WWtM/PDqx7+V2
4c+ntg/VYNrKK2RJUr4mUKFgoHUZS6qQ5YEROrin/H4X2yP218hLmxZTmHDvruPh
Sc9AxRuh6lT5NR4E5j+wHWVC64DCO+f6MGHwzFzxDCR8nBj3yxClC+NrhrHwp5Jw
l1W+B3Kv+r+LlzSNpKmqzNYHBzwGza2aBmLPtaZQWhfzEAQw+wI99vAPxPhVUcvG
EoemdDlppB2EFYdSF4Ot6NKQuSVNoX6ANI/HI0dyFNnmp3Mc8aEwg3ZsG+8Hj4pd
Tx4f28iX20dOIkUFBdTc+RPEaNmaIOn7T845aJtuX1ZxV7vcbI8G4IVTQiA38r9o
hqo18xSTEtWhV7GyJnltjpXllvyiZe2EU7bMFuQePezs5VTxnTh8NbrhKPKc6Uuc
Q8ioY8KS4kCgMbZUjbULjO5Aer030cJ8PRQBDO5zC5djX90V09EfjhP3aeB9JiGY
/BKG01BUYL8y9rno6ONLZtSQh5N8oKPvXZgjqlmVgxgvG/57qOVjQG3ViSOTB/u8
zjYKuOBnLj7n7UdtJ9Bhusd0URzFYAc2uGNdgs3TA6sv73Chn2FZcYxt26VIgn1l
Z69k/Yr47ru84riDYN7ExQIbLrTF8Y9uqCOjm4XYZcpkjuVcgVZRvhc6qCS0ub5j
iYcx9gKEp7bj7JGUj7+0EprQsSCDna3vtTHWfdecjDeBc13aYTfILA6xR7FaF2Fy
rXzaKgAWMXmc2g7G+seWw85hcWdrCXpUcnvlpAwPoi2fBbE7MSUQBbr5YhOzl5fy
Qgcr8OJ7iQc0pvQuo5byf1MIs8plJOom/Ga8dY7NWvGqdQ37vC8M72OTHGBqIybD
pJGVMa5Jun9NVhqkITu1s5r6wrzyAIUsF+vc1TAj7KZsIEfI7s03C9vFr9H/ln4P
02wF5xR2EPYlzr2nNJBFqQ+9OedFjibkDoqxKUSVUlUNRbPyua8gBlhppUpVyimt
x31kbRsHmBudls7E4ZcZBw==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BKzndpwsnuhNnfxZ434TQ5xaU8tdrdIBYUXJu8rnjEpuxjuRy1lyCl6Y0FzGMMqa
shCGrbgFHBNrEPqXFUujc/g66oQsSbk+SImOoP+H2aYv05nnR4Kzx2wQeiOcjhm4
IjcsqPWsYtt2lKUSxjbg4GXXr4GxWyF7+M7mjIbDhHWyLL1ELzkhh0zOyOMC7Ems
5s1mfMgpGay/Kh0nD9zYkk1M3y1EIBHzaoqHdOAEJ3XEPj8Q1p+o99Z3cIuDq7Cz
lqzHjAOjVqTO0Lx1DvpBjYiJwmcaUmDVaUlcigjE/qpdoXYTp6PLV5zY/ogtkRkI
lQvi39o1IR2VM+dzh7gBRQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
Lmvf/S+hfh6Vjb/bkVs63697/H2gGdfcNew2xXUDubM1rYjIZ7gYRKUsbbbw/4QU
0XA2lkXTmn1M/zQJp9gnU9ZFQ/wMsy6e4DSbAvXiXksOuyhqNow9aGwPxN6xguaQ
1/Gn95mX3yIe0IkgXhmqFZt3QwpnU2i2rAvHgESzcT2sDbc5Kmoobgy3PNXAl1Gf
XtYZqrULh4Wc+67b2AWX+nYL/aLUzTWYhj2oB3tU8lqh0nbgO1uekZxAc31gn3hR
j6tIX27F9jPSA0G1J8S2A2h8uPge0zl4tWA4fPzJi/crHng1mqIBrGWSx/GqQBZM
eE4oGzI3IljRXXmFK0Nbd/jGppiEvm7M36jYre3RQfrNiu3jWY+GSLTe02LCPzuw
D860cwfpaUxkQc1cbWGxUeNYAAaOIRjwmjNuwObEZ/Mb6E81HgEGhM2jFm5dzYE9
CjIDu8h3cdSzdW0uH1/Mpc1GNMFfgg60G+2qUQg/f2usQnmrs+08xhwMuYzr2hT+
GtyhD96w0IjIAaHnLP2UKIjFlJIFyY8NrNzCqQp2mMvWEH/IBAbB5MFDFVao/rSm
WaHdFYbdkPLFEphlC2Ynlg4ocdlGa+m4hppSBnnLzuh5FSBCoFQlV79/PdqxFxpz
FdO7fvGJBshMZhI3pfUOBKJ/GN1hnjlIiYvHCPKJikKsMWfJ4ENxdMXmVcBjKuUd
dGKtZibUtWma2SMtpDxI5BGn2H7Q195zeeUp2YSN3wETuHLo0NoJCyMsbmm6VUZS
6haTna1HbqZyjeev/s4rVUmHmBZdzTUrXXCWGxSZoBw8ip2GR4rMjPMI5uuvbdju
4mrFbQsNpcqyTJ/VSWVWVSjjZpvf02kcpSqQ37pUcgdy7imHhk1KWPJDVDamRNfe
Ee8bNruJX33Ynn5meVEJxwzh8tZpOUU8phlhpC43nvvxs6gc+QRwtLBh2t5ax4D7
Wre6rHYWgYtAyIVlqo8/n+3O/Nv76F4aON92H2sIBzaDI9MfD4CtMlgo2RczsYPN
wcwa0ftZDIc8pOJev3MyNEXoN4FlYAu6yy1rY0C8gqZeVa1zfiUhnTcHR8Ty/JRR
IMxElwo6h05X6xzaDUqeu95+md3J+pAB16JpWeD2D862mS3mQ3IitQrkGcD39Fpg
eXYZlTg0UhxLui43Ie4uyhFv9VOcakxOvJ2GL6Ono+W3CzoNFLsjhd8CasJq1pUM
nJuFhDe453feAM+7mMpZKzUocyifWskBX1/rqMIGdLGhnadXpDJ5WAWZitlrDzVG
1oWbqNHKeYgOxtI3t8RMskRJIaGIc8eToMlEtbPs75bIaEvyitI9RuwL7709vbQa
RcR0MROMPCDu/WgPWT3y7m9rjGnoqv0YxIuYMU6NUOCrg5MHDtUsMkqT5sgjxgGD
KTWxBEL+YD58tjXfrqXWHM92dsu7D1mBFFvg60NBxzXBe23BPOtqXAPc63VgIRMo
xVtl9W32MFwvNMN4/a33i7jF+2kpB2L/YdLUuTyE+Tt8M0PlTw2aA0XXFStNDv7v
wIlkUkdG26zHZwVv9W0vW0NjUMnIMHw9xO5v7+qHP5/VsCm8CVqdM/8CIkszb5e5
BH7ywt+87If1AVZZCCc+tFySffAmWXOYOVvwQAdtxshnrfkYAzWs3805jPtIApos
nvsLkw1EChFE3McbiDk7mL+9E+9qtltOh66fjD6xjZfLDFQT/2CGQjS7lofc7Ltu
7z+g9rqu2B16F0oeoTF7rhR4fM3DQ9trSyzi1emTX/aav3C1+DmRyPA+hkSZwv8n
g9Vafw5Hb/4tbjftDC1NwuOHxh7/hpZu/qg3TIQGbhHZW1UmTmqj9C6BZSnlVyss
GfgJ/WdqK9UYRj4WMtL89em0tFzRibSi6j0XUceEJKilyffPXxKUzrQCZ57oRO4u
/GNrjmdOG1hdB41MI1L0Zl5Uj0Ta3Yhm+NfRJHqrQ6qzi5SARSL1VVocpBHujVna
zwXYMLZIqf45O/I+NvNlgFKZF85Y5T4kd4ZNiKVHLOzBmv0+GrRvVo8ECk2mljU6
WVtPti+Z52upOoX7OebOd53ukhER6PCUCJlspygYvQUasBA8/b4T7hT12rMe4o9h
wf4wbOdCahzTi8zquzPQ7ENrU7TeghnHXn/3LufDVvyH62ijIAcksK8WmYwHc4gE
ahwFY6TezpKfpfX5aAbDwJSkOS+aQIzigDb9G/K6RV7YOlyji2yON9rCIf5Fr1uX
/Q3EGHHENPYi2kMlFwlj0bX3A2UUEoa/JdFyt0cvbREg8yX9Uq5AjGCIFqfwBDRQ
+UGWAc5nlVp4Rq8A+NTsqWc0mk6e3VOSo5Vgv4KT4vzg7Vv/xvIXcPqVHH7Ft+YI
DQBOXmI+vZtyvDMqUKQba2jD+kKSptXV7sV0+kAj1RZoa7NYseDOW42oF4Az8dU7
+B0Mac7qrguEgyYq3oglDaYQ2YX1urP398lZ26EqLntOL/O3WCSCGx3SDpY5WlDk
DGKxjfzzEMnEb+2IGZeNUzIFS/z8w73T9iXR/I/63Ncinne+UUn0L7GHo/2QRYxk
bNoDbADxDu61A03k5A/Q0WN1DEvgnUP01JClB+lMIgLiCPsiOJ2C4GGfexjbUUeX
yT5itgFSyI1jNbQotdYEMoYQJ3KtKftuUiDQ2Ms9KeDdcr6mgcxxYWYCQIM4fm1W
HYq+f5E/8Vu9YvV2nhdu1xycyHnwliB1GrcP4uIfogFrUo6GW6eaIGCjDF2JgY9r
XYSDzTi6LXuMdeZjtIMwCNsh+hQiLq+znsVFsd3fWQ91RBPiwFQlb8+4gW7H+OB9
O9t08lPiygh2Xoyhu1jKBY2sawYxC/hVYsUqmToQgySyJjgTL9nacSFZNTmNYai2
k02ElFKo97pq2Itad/H1X9B/BvA+C9kHI3fyCT+mlzHhQRq7Htwi5BB5V9zhM+nu
SSbTJKSWzLbXQRCEVwTbElFUGXoiGTZCdXuXlAbwg9bqUmzbBcP1fyZq1OAUXRWy
Z1o5nG9Z6f765oDUmofKptjxjszgTKK7b8l5sFyxgBYoNQiH323V+DAEhZaVweZw
Lbdp9CGghwDCn7rfRtz2UfalNdq3AGnPSSzyIuKYaCZKGRY67fpV08Prp+jUCE0a
HNEIMRCBO0npewR3RalvRdi+/HX6ZFJUIZ9Pt0uv8DQuTvJUIz5IbHjymbzhvYoi
HL5HB0l7yuTJIzcXt1FTkzraWie8GYWGny5w+MvFO38FcwqeKC2Jmuy4bYdfqTgI
pqwvBk1LZS6jBP2uWXKWPLGPfVBIFLUgzg0ymrOwcaP4uPmP/K6/a00OeIv8VJ7e
2X0GvZeSMgicN6GXQryLfa/tPuLJhd4U1V7o5aEF9MF08WayA4ckcRXuz8nKGzjN
sme3k0e6zBfgLDtHudQyxHbNMHRqCRE/bEIahFkKTsxtibAA58NXvhgTKzpx9hP4
VZyJ12imUrbRizGWRyK6fCNqOVNjNi4pIO9k9vpWr5wfE4PXr3DUiNDRJRGdPXhy
BdO67kHg+olVC8GBbgDzuCBbdL+noQqWUddnLNoqfjlSlS2THqMLxH2kHUJF6I+A
qxal0mWVXv/FO0htP/E/mzpf/iJfBXzN+3h9Dd33ZtEFn2o10VP/nuTa0RARry5x
NQPQpcc46ReBnKtvbSmEDdGnb4c219p5STeADhHEG7VbLrPEg/Mpk6d+atWULjQr
4L55bXxxuzicJEygfxDaISiftxyjByVGLkSHuzNGorBNBAMSh5Cc4+qXnD/dYW+m
mx1gcyamjw/4eirF8KLlM6Jnu+5RY9pnrrTQDPAV/ANrRLpluPvOS+4w+FrhXxbQ
x9nO3kEyjbxBbcMuIGEyXPSkqR01XxgWXSz5FAr7oQ4Re9qS9+9OdXJy7TxNnV6J
DlhlOsdrOIGm4bSZgZy/3wIDvWv/czTK+Tqka6lWg4FPQlFeWRWDUSDHHYdWoAnc
9eHxCUyENutSX7tJBGJQuTSSjyx3DAslETMzKKYH9chfowUHvCbzST5u7Y1KCW/i
STykH0+7NoTkFidJCzp/UrKy0e7tC5Tric7Kd0ypviHNcshgYfORhL1aXu4Y5+oH
M9SiPkesG1UlxebC9725/05KXVadGLNSKutqiYcTqcPjIyrAzVtZu/FoTshJ4Ogf
wWLgn2eG1K4LKh4vPloOrrvVJ18iXKjoaBXVaDHpZlVMlcccdRs230Uc/0LD1xKG
2O8+TxR7OCeL+vMnKBlB/M88Tq1iPULxn2DLoD0jdL7ye6FrzTHSripJ+ZsQ59dm
9QG3SvBfHPstEtzZ4annwDBdWO0agrZLi18YePa9sjhxFEEsyGhrvvTrb1PHSLZ8
MxEvPxa+slLx8PtzYj0YO8hgsKMDxFUq8QyYa2gydfjYhxUIUnpIqME+wZOSJjad
9++z5IAYXX245LkiO5WcmCfCBaIDJcMX8BzDnlQgP2OeZXzPz73m/jrmDdmTl7zQ
nUj1+OPJlz4t6K7gtfbid0gCCAU9/sAFiDwfAXvJGP5lVkcCLjmuDnhoQbGTfHRf
RAuADDKK2KLsEpPuQdMFT4bKAeXYdr5rLOzLmkvH9PLkzGX/TuTNPwZS6sqX3E4x
tcijp+/gv8ymg9AT81xBVNQONOlrq/vxZsF5cnyxUGzWJjLrbRX1HlS66ZMqEqsU
uIrnGwsiwokXrHHCPmsusT6wSKHbd00TI7YErviV5zPdIXXTMWfSZujEupE9LJtn
wISLMRUAlakE1fLu2cgKjRjGMvJzGVTMT5ktzEvXtgxNg8vldtNZw9kunnVZL4Av
f5ZI3TL/WwgMEKaDMB92p7WuDOS10rFgwUfnH46syomddCU40NEIHVVfjuFVnwel
xMeTbYjfTmqbFg8EIQOaY6tQrqKX2S7rnubHkBfq8lD3Gg7tO5jKb97F9oVMcMTZ
IpHLNRrn2+zpUw2Q3fKP/64hi7pVs7Bpk6IUKX136NPpz+EAv7rqknQ9z/1G3oiP
jcBawSavf6K+Y5/1qDBH2Bgo9qiejxPtg0vY29FnPojlPmAg9iPoUWEIIOay62NV
y9u6lUE2Hg4s/WacgoH28UMDxKjb9FfJKVcTBoQeITsLmDsJEBJixW3mGWsli9D5
TOjmaVZ5mCrxC92Nd4YBiAhPEGz9TAHEcViRb4WXP78=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Az8XnaxiQE5yh8kN7qKe2ctE2NnGJneayVw2H1ec4Fg8Htl+sRCU01vIMvEKj3gA
B8ljBgdWZLhLMuJXeaOduclYiMnh25RgRXzCIKWDkzGV6RcsqPZmTEL0MX0skksS
fA36KEQs756aBafjv3hxVntPT1+zZQNAxG+CXdB9wJxNWkzx5tgNGC0NJD6YHz4u
ez3HgP3fi9G/QLfgBRyBH7yZgpprv7wcWAKepCZ396vMLA06JQ8G0Y7RODV6WVDK
wmSIRBfeJHO5//8QtL5YcNOi0I1aD23vsmJi0N7ZtrQ5ultKuSMLxv+TVxHwvWiR
A69gVMB1Ko5TX3554+qNNw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
ExI4JvY3+0E1S01FyhVlU92P/n4cYNEzknekiRp3sCHXFgHHKEDHRricTifv81lg
BDNRzczyWrNPMaEYhW+v/mgN5h2c98BLUW0nBhv2qxer9pN0FDpIzC1/hyAttZFx
Wt1ItBwZSB4k1ExRQ2nmXu8uud5pbwvC7iDAGIyguJjzimMFPgjH6ITHRwye2RIH
vIzRTAUNW3IMJ7+ZncVy1/w+gfOkDqK3PZF4KPQFa4GajG7+bjlnmfirSNmLAwCw
y45bQai1mIhiip3Ca7CNK5tCmI2zj7kbs+asVTk0ehgLCa95eR0BoFVYXSCjz16X
efZOrVSYrb/Fmzo1ZlVXDUs/OqER7exVUu/tLwleT8X1WOHsrxmDlXcDfsdsVWJY
xp5O9RwipdBPdS0qT2T7tYCkuwZ11cC1g0Lps6XcU5ciIBfEE6ru3U7qzgE0SiH8
xcc7KjibPkvWYgIgQrOSn9zwWhvhX8V0ogj55gO/vpS7bXNmsisTWadg+q2MU+n2
DEXB2YOiVZPm4qaK1Sflt4fTizDIi/QT4YYiZJXBdxwiFUMIcMS/E2ABbaEy+96V
7el5sQQJe/P6pac8WV+qO85ILnYukby1cO5lpeL8RvFQf5IuQpEPkC+fPzih/17q
Yawu82oh0l55swOdFbSF2GYE8x6ctsQ+hOQ4i76xxYG331nX3U2Qz69ddyuZLZE6
OWTr+0u+REaRc9MBpGUvZENgVE4nFjHnsn2N8LoUs6WXJI7ynt4jUH66Ku9COupw
tzHCI6ze2qGmmU1ZvSdgI+4fDiLHEGOsrDMrbeDNqbT9A85oXFd0sbu4Zo66Ly0l
a3wEGM0C5VwpgwvDtAO0aMyVYxhanBYHD/1lrkOLvLN+X+GtMiIIdome/XOzPsYP
dzZJQBKIKNifbebD+Jdft99QOu8HCCdoqZMIEQX0UiRObFjTJLeIr8FWwtYa8+Rv
QmjiGkUJ10ggVz/W+R1gyHkQkswizNE85RJM7RRkS4ZwM2Hi6vEyzIvb8P8eiIJ5
gNZcPJ2XzjHHuhVmiEVmrlkSYRUWgHGRx0Y9zPXHxA/U3wWIUtrgOcaweDJ7e3wA
10Fy8BWnCsNI+RHa9cTfz53vKwi0NHUohZNiHqxvoUd1e2MAUMAvdzjA4DW07JLb
WLWuYDAPLmHnrgXlMY+7TJr77091WbinKbq7dMaiPdF0BA2R5aOcu00AghyqyLSA
Pzc0/LUC+dObaC7KNhNoYySPqP2bufMrqjX9Oo/xsL1Y1ip/2ASv5/N32Td/JfBC
RinFmepsHP68Mr/DLkdmuY2j5jjaSaHeLipOANgr3BKfyQTd1GA7+GzINEz60lGh
LlkQiI0LwkOcTxPeT+RWcHDEtIfXEWrOQGhQdXm7UiKwSmksFKDRCxyyjf84UG2e
62zXnUkn2QS6ftCulbwmte8u0tUjuUb40z5nsCe8nYu/MaFkocGX84jFztWIjsIY
2NHpOQD/P4qzCfvuRKm4rn1qiBH8MnMiLddxUBY03aHLPGxEsJIIoReBS5ftNzs4
CaLWBea0iMRrdeeup5Np5MnQVGTRYfRgBAWYYmVp8xP2xUbKzCZzgMJ6P8Oqp8vp
7ccZjoE9Hd4TJPxLgixg1WXncI8BhPTL7cxzLtjlSAY4p1bOI7jCwLASRHWHas6h
oknv4mkNKv2LLT8ZIzY0uHdhvMxrMJYojYKtyt2EezYh5HnBgoPQk59DFvSISFA9
gEFBXfyDONZj6b520koz0IArrlYHNxMEOm4c6YWTROdpaZJy5XWJRkbXbs4uMKhQ
BIETzTfb+W1XRisED8UEQd+CWTJ5edO4PG4/j6xUhBhQz7tNh/ACk/qLgksCANct
Yp551ygnKdAdnboE21GojpB3qiYgezKNDyXlv2GqAKxnzZ/UU1hKF4lKFnV3W7OR
bT8KBAm0jbUQQDekuLpj8IjQ8NJhEzfzr44hwp0kBhcbopH9UhQMdaCh2Md7KV+O
iRRVkpQm8wGKV+7l8XEdcAq4j7Vxkz7ojzgwIGD0yToUnJABZDGU7U/qL68aBhp0
VVsTSIGNPUYNZM7BmQCsKP+/sJrWICUD/3yJGPycjA8OCKIbq331q5Ua+FM+T3Pi
AkioR5Qakuxva7pB3ysDZrXFom+sY3Taf6CPkEQKOMd1K1iVhxYbvKWtlk2SGi1g
8se+bzQzMkrve9Ci868qD/XQ6eKV2vlv+Ddd7gtMCpWRkVzWWA18KmnU36qOPNcH
k2vB1znjBkolKrIMEauop6J0OY6+6JKAk91toO0LCxsMKlLHF6uCvb+198K1VVn9
RpCvRdW8HF7ajeXQ/LZsJwyAyfpv7YFDfZ+P1el23OI3fZYKqNr4GRqordddHoMf
hw0VdMAFgGveS9H/vyGt/B7MYcky8dHsGXpEBl3IcPGKJZXHsvdEloHx6FZW2Lnq
uqLS0AJNgTnlayZXvv9J4JzyN8yzAA9bk3RcgCqP+b997sB2fmiirnaAwktD5qbd
EnMi7sqRXh+JPLZqhnyBtAAnpcox3o2KQtjE3qJ5ORQVrOF7fytAGMbnWar7vSdX
xqiLE1IOcD1BaWZ1IrNEmvAJ15vA9O2d3CwGD1RmWBg3OOTHAUyORtqlxrAS7rel
hfCL6uz5fHNmk9NgOfmJlD5W2qDeW/Cbyh195CsWD6djqccjEcZMFW17KZwUxwdt
ebgRG1z3hI7MGj1KnNUkhcdDiPFUGoxAyG6SAraMeyu8geqd8SVhyMWNJp7ECDVW
U5nyZanwIwoQu5yUacTLKgV1qjmiOtFTXURjdRW4X6HftqvEOoadmQjXLHFlh9ea
KuQYW4W4LrGdEby8HdYMl0JZmLHEsVO8AjFZn7WNbBbpUYpJ4NGr3ID9BxFfEQv1
n2HrLBRSccdvTgz0um6EA6ccleEc487MHLMpSLALXvgKeP6wx0u9PhAsiRbT0WeO
6QVrKGDILIK7E7iXnuc7LDrRBr0HKN5bYdULX6uhwVAzaTWtk+eTYbmCVtgjhg+L
TaPLic5twQ/yrpsp8Z6b7lzPImSoAGLJBtKswhkWNe/R+qfgoruwROHUIgpA3m4z
roKb/ls/Etm8Wh5Mz+DwLVSDwaByw0/sbEiG52glsTogEnDOrgNNXsOPkEDV8AAv
fAAxWdq2C0nygd0uDXpJiKYIqpYJvJ9Yf/Zx7P9w1u/eBzKOBaiR4VE+XvI6v6YF
CAbcjASIeYbpbi/CfX98sNod8+tqFSg5gkNwtb/g3E3nFi+ZxIziJd+CQGR0kL00
Fwu4Wne9Esq/JT11H3PjM1AcZCGMHCzBT26eFA7MdYFacglBOkj9+tjMTrtilZH8
TotedW2Jm/AxRpp+F/JP3pCvzo39wyqpfO2rsJsy1MmQMcmkXM0qWQB+lWDxCN9L
bkNq9AKS6ESRbW9/ECEvCJYWM2FSYlsKbXPEG1Pp6Na7Sj0hZ+p2LBajd8pRjIu9
WHTYlXeCWGznbOXNmijQmBVvKwmGDGdf4Dt+FWAmP3R+s2pDy+Gfcui53ct4vObX
ktVuL4mlrz4j0qLv/Ft+atiAawlTkP1lTFImTUWXoaRJwAZ5h64MRkSz1JyF/7Jj
9cPF2H1HFLB0md8hpaR7WADI4KEfiWTE4kK/ZfWReAy/QEA7iGP8ZKoCFK8GzS1h
ILgUl2fl3cOyRMn8QPDBk/TlzyzA7z06UfIpmotSpIdDBAOoWMjtoI7pfcw+lMh7
pe9L6N1Eu1BFSDs8Db1sMvJL/Kspv6aAL57jv8jfqrWDOoEJ0VaECx31sQH7ZpgU
oHn2iX6cyu5Ggyd/UC8Kq16zyAKIRPLZTU4RJk/r+w6np6ibto506Lx6YAoZFD0g
WfeLq7Btx8+TTaxsScPHSqpV0DhCP/9qdYzt25t4lLP0a6jwo54zYSFidF4lSGra
0peEUaCrSTzPmKjiydrN4UcXsT03R8d+OwnnoOEcuba5EtxTLZTlX97IfsZQDA2L
9AsiIK02BhAfkiNzTESf0TO+nRJFlq7dKPiLhUdJH1tatzEUfj8P1rgzeRkDA138
dWKfwyXL18L7ecakDIRU2ol/N4nkXopV9dfMqaZV1gScvHqIQmHYwxrdfxUyYK0S
AdX9BNDtNH8jtxt6bTBYomyQeBltJJQcJsoqAtJfoVo2WADJpo9qWV5+yfviyWho
PJ6YlSfd7CE2Bh/5tXFplPB/PdSK5QTvy1bcM+j0TzaOcH9rTR3pJhmAkmrHHNyh
RnpyE6cPBmkM8C05VtBTuilrUtlyVs5Ve3vrUXLp5SnyXmZehtX7F83IJXFafuXV
QpeP1qLJnNvKmYs4c5ecLPkyeX3tUf1cil9p+ldoqH49Lv0k1TpnNU/pQS3l/Iy3
JJ9VKWuKhSXLDsO+d3kWIi6EdMSshU+T4Fw300EK4fWjG/SRij/OrEm+owguOlS+
MxCkN6V5ztIM1+asBUgdgWJZZzeeEoEp8zR4CciMP+6g4poyCLhx2UAQxqxRMUpy
xn9LNk+Vi1c4AYm3DaUTDcfn/ZjdfXL7F90RJgSnG7hQO6mQfaQ1jjt5VQVykJz6
zqxpSrz1s2TdCX/yR9N7KN8FBEdtxQvrxuKk+H3sKl3DxADJwtxCbPKhwgwYX1Eg
zR3wh5pkcnd3nWl2jmv3HlnkBrjhS6yZeXVHXOAabblbZ/5DZxX0KKT0evb15+sf
hzIK1wqe+IGhE0s1L22j7dMGlDYg0TGfsC0a8ZZMhWNvrg2jP/oQsB/0iP9qmSvH
osqmYUnmguCTQRqGtXjpL09ASWkAJVMWeOLZcwWs6JAnp0fIKDpkwlk2HG2SiDDa
FRwoORMEXjlSyA2DZ8rPPDtaL5xJ/GvBYYveb1II76F1iqQanESAwVdXZIJKJL25
6Ym3TcA1X/+xhlaxA2H0ecHfbJBzUi+WIiGomMELf7/z1sWTBWqkq2eeqF0y+GOU
DogxRswB4uD2WpoVkTJ2TVXEhebYbZLrJcLBD5YjNXg4MlA0yOBPuBvOcwNL7FjX
rKHsZvPmVb1ozA8OPCNyglFcVdT1/nLScsksUmu6AonqAOqveavDBY2PgMxghzrT
qhVP1BNhXpeC4MO8u/Aj/0gUGuKDEsd+zHrPc61HYXodsOFD4AXEiIS8P7A4tYSj
+0fp2NHqwzIP+jkT7qXMJThf/Afv6mnZgarTYcoqyBQIwFjndqiS6yzNk0+PIrcZ
QIDFP3Kn3+w2YWoRm4llIh1gZMOz0PRhRwgKYWM7tHoFaZpeuwkY+hPJzRGho8xa
U10B6CdkOHMwuL8Ha5Lpe7i19GYLjpnddhTe4pKomf02NMNnlbfPUXd4x7SqrYK3
ZraDRmuanu6rpxuzMMpl61vDGBP69DYEnlAsY/vnzMzfCpWZ0WjW59ioQxb4VPs8
7Aiew59Dd/DZtSwoa8hvEil7qMcgWU6Ep1RuM+VcLbO07CzDoURnpeTVzHslAgGK
Stb7gEP3rDcWS4ZszzMlDwL8/P+4OdmLQwfkSmBeLYg/YxGPxQ0u5Fh07giAFwBX
3mmB/etjgT93SXHfseGeFQpNSi1NVpCM9cnZd8wuMIsnf9MZ7XpExzST703l4q6K
bZymCXWbibT/hEu2E3I2I0Q1X+LI89oA01E3XAhmIfXXEdHd/xuK7mMAGcFn1Arv
dbSl7z1+YePtICaUcFXGuZjGyoaWs7j023p8G1MNwOtlV6dHx2dBIZRCZmyaV2Kq
tw3k8+jJ3XMQ0uFDGx86NO/RCCxnz5sMYfDRwIZg+9of0GPIoDVWRz9hSRSv0M42
qb91M+K/m3VF4GmyPpC5jGGQ34joEc1H+B9UaDulQw8l4fivRKOuYsbqwLW/sWcg
5IL9KVt72NfSywMCyp+uV1D99p7J32Xqc4F0lK5ixcS3n7Xs8guEU2jpqODgf/n5
G+fvSEC62xbrhUbxCAIY+V8ac0Bn2bRibwcVFO6IPpTjz/9zjN51zyBOnjg2D2FN
AgpfslertSehKziJQogxdU/1r68QCRaZXu37FnyJXtBqvzvA5iDKvCXpPkBMSZOk
4NDS+iKO8mOQ9P+qXZL0fYzT+6+byxdHNYDffsmHbAw7QzadGye9YbndvuO4ZoMK
LX5Fgguvx0g6dKXJjddNKcpjl0Z+IUrZ9fMmfVu3R5MQnJbQEI4DT00kyCFS+ys1
QT+a6aHa5gtEXS64mxqYtqwTirZt+mkHtl8GqEqOMiO7fOm9j4+abOEjXPgYanKX
zAlypDx6y/xQtBj02B2agRV/ltiIk0KEfd6WC+tF0trY3SpnNDg3+0yMuQ51f6hk
pmw/y/zM5b3Y4dPxYw/OuVupu1on4KBwSMKZ4+Q96+USPDadR4GNz+4hxnCuCdL2
I8MzLna8m0GfsIAVAArhVYbtXJ+08hmd90AhhC44v3S+/84p9TdMh7YJQVnn0ozb
ursNUZX1ML3QHi2+cqEZkHIgyS55DCE1qdVAW14qA5wdGaykD6l6tLC3rzHtPqqc
n/uIW1KOmREzkYPzxNKkXGVlDtOgQyVsfoDiTWZoUrEMi33p5ZYlyuMOO6pfTUF2
CuWRy5YRUAiAWsNzRlS47lsYG0lWE23zxW6Mx72+qhZA4SiBn076yr2jWecFImje
jI8r4JZSC4oZCSgA7YqN8p9VywiuZX9k/MZlB3c7jIm37gDdr/mp2Y9OTPCFFNNm
OX2kck3GK2MnUItbdXWrZ2HYQZnzYnvuAIhr4zJ7rGI25zQv/hgQY+CXoOAuy+S2
WhPbxv3bdAdRIuw57mveMHjw7kIriEow9f0/9hbLQOC8/rovIUY6SSv0zmXNLX1e
ltkbaNICL15T5npWz+WrkdUCf1oBL/tEEWVEKKx49/0hTuVtHBkZYPycKZoK5Gyf
tukT/hHpMBLsjzki9a0fhbiaCQwA+RhWP73FMlggXMWAQNZzIqo9oxBPTRoGqc30
0sAqE6rbs4ffg5Pzid60fXCAowCg6EShB9eTj7MgKv6ESKxgeP29vxGfR35ism98
scrA96VbA/327RZROaQdPwerQamPgvvBtW+eAgCXndjpInz0J1hLSrGwJDgF8LSZ
lemdWrz7Pt3xMgqvhUJ2aUMRDVVhqZ39lfxBFo3VVvLN2pmpOyr0YkmD0EHRTncf
buZXSzmffivRAD93n+fFUhWgJpI5JxL4ndaO1LOS6+Cv31XNWL142SzilmjweCGr
yFfSOHQ1U1VCaZ+UJkHXCwR49c84yKyp0yc9gp4HaTPIn7qpqOoEhuG21XJQLAB+
EKXwoLMbOOJPlihdOqD2x7u4NK4h1pDCID7cpdQJsR9zjLrmeHU/7VS8KPKVQAjM
HPdVuML8Qc0B7KykvsOID+JexfzoUSJXcRTnp+1oae9oGlWpMLYPLGSne9oEduYy
K4v50O58D2gtdbL+hbqxa8YFq3IxOoPUftFxVeBFobtL7ubL2KEJw8mLpSn6ct/k
6hD8Q4P6zB3BIVhteiEqgOz/PYWtlEazNyQYucWZzvMckRjnZxiCmJuLRG34bMvo
u2b3mXCRzjO0gCdbxArI01nEnAMjU1hS2qXozSI71Nk6LrKVfBAX0IE8BMKADcTZ
atEk1lrw2C4HJYulbRwvvwFJDCcNhyxgPkya3pYROuj60t1+/Lw5TnTiwDkanUGb
juyHZANuqHFPPLF6Cr2R89S8q6iSaY5kGouUqa7Q+H8v6ZuuiiqOcXKcEVRKEGsK
ULdTak7Yw5uZggx2YJRljefJlsfxSZtZwiwIEFgAQJojFcc90uLbMqwoyYg8OCzq
VZxfda2YsQz7pIAChRjNp/p5zNbZpXXqUb9kaPyHBU8EZ4SCdXp4Vx6ItoeHBp10
FnpF6KGe+GtauE1jOeSLbDa7hE/IcO8tJ+SMyOtRdjhVVde3TVOlJCQ84a81ei9d
6hj4NvJ7J/1lchuFYbhE28+kNmZm98ZceHz24AW5hutkK8YeJb0gmNn6KrFdLKx2
9afQqNaxubp1VbGs28SqJSSJYpuNjt3kLF6MX6eKDce8isz6QASKIKEpfSHdvXcK
DKr9IjklifqYJn++getEnKFPjwJJFLYFRW5hv7yzPLN+p8JRD4chlBog7pL+DXoX
tBTy5Lbr9xkJ17pDdjEVWe5JfS7LK0j7bOu1wsAhSnUr7/diEZcS8CqXUjLJX6Up
R4RuWeH7qp8hip+2dIKHw3Fxk+7MpPkHfW/6OquJeyTgAxKP73E2bi9Orre2m5fY
B2w9ohWaQI/CMUW5RnNOMLe/yjpdXBBtDgQNUoanJ0nRApUXa3xTcymlY6A84nmj
Zf9RwBBNAjSorT1UUZmhGC1v+ri0n7MiKqP1dFbzOHUpSdW97ptjNLqJmMYK9O3p
OhF/nhAppYhGJhs/V+neFt2ue+/GzTjHTHSBvsz2rdcm0QJ4fX/zFmBes/SCgqz6
5vwsEeQTaYJGMLxZ8X2OcVfDx+23zk8xTaFs01gxFcnig3Ixr3qWZSrt6yl5FO9V
p2dkLX5BvWm7b3XhWOlcJV8y2FfzaMB2aOOPrI15uyPzatFn12OFT7WKcaYbAQp0
hEdgNLcKsNo/2S03qhTvpPpDIS8Qkr74DIiw9Qt7izHd28vHNu36EXCzpTmQHTak
ehtJH6B6xLGVUk77kc2LuGF3PJX/RqvoRCYKjj94VLKb5PKP4OGUnbrUnkDT6pTm
pBARYORVUhKuOJQvuMYsQjogNsS+mvWri2aaW2QafZ8ZG9DlqujY6jNaH5oNEXhI
zmtpFxI1jHohUZ8acoTmc1SdqrtR60SWiWsVtjYHAdBiGfc9EbFPfEmTk1c19gQM
YQ6tKfAHUFEDzzUUE+I+xDmbbcAaUb1+oAAMo2lX+bsYjeLLo+X41sIUqs8kIYxS
OpCm10IwyaRm7DtTwT3Bf5LjD5yskq5B81oYNEDX1ZBB4Oti5piHm2NBQFt2enwt
IT3SrgaBgM609nVKy00onOLojLjzm56GwoB/uI0FZfW6Wdxc+Ad25KJUEScPwREM
EYt7frN2H6e6Dh3USlM5DqsVPqGWPE+B02aH7ErCf1lbYJ3GzkEa/lU3nEw/ohmq
NiC/sPTllrHdNBg9vbLTkC+19S5NmDdBlgYfnhfPBRhcegSHv7C74coYb4dMNM61
E0zg6nljW0N2QIuSVuzjiykCx8D9ub+88vRzjlxCqT+ZstXnnkrvSu4YPzNvdTsF
06YWCNV56KwpO/hmFv9d2MoiDmKe1ZAoI6e0Kf574DUMop2Np+lFBzcimAcPCMWR
HikxWsRnT67aBUwQ1EfQOBaLw68WlXrjSw1mUun5BVBwhnPQxJa3d8B8yY52eb/L
1NDovi+KPmn29Vm6+395wlKYtv217CO65FOA26uOAeuyqxw5LHf0yuYT5bl2EWiF
d4poyt6apEAYU81hGBbEiBAoSAHxmV/uuTfzTmscNsYbJmqp1jwpF960lh6SQ9xw
K4dUJ4d/YvfCDSxRnN1u1J5P/6andgEhNpUMzZmpTvFSdnDEp+8iJbzJBYwk62dO
RYyKWyq5S/YTy91pIv+uihRMzO8X73HRM+Hlni9EDSYFHaZGbjLKl62WPCtnLty2
1SIgBqKe2XXDGwI15Z5EHPUwnTsQpPI99dw9dw2vQImrbm7PerEj9YCDlg8yw83V
Yy38K69R+/lNPAeHaDBV2AMScKaLttayXvCNlK2eCWqUU/4phH7Um4tWzu+gxtLV
n8HQQm1SL3CaMR7MMvy18F9E2xHCQ6X63gSXRAsi0Flxslhck1HAckqnghMkoQ+y
imQsbmx+A0UFJ09wFdxzQ4JuTC5cQBCIGVOn6t4DWArDn/Dq+/KtlOUTv8MlEMZj
bhWj02ScRxlKPOEsF7rgd56E1FW8SKEhS4s518NLcYIb02ukTtGLtMf+XQ+MHLmc
3Q037Dp9RvrvNxBIRqWXRGcYF8iW/5Owq1xGVL74JFiZubizspEID+UnX257bpPq
y95izn4ONdngD50Idw7IKyETwvjWHo7ZAYkXg6hoJjDG090FuYUrmrQ2T1RXp4JQ
BOxJNtl4SqZxfr1lvTBK2ShrkYXFWkgEnyOetyuWvZKyPXyAJJgZBy8iXyud1NZK
mylVp9+EzDUykdBiSRxGWaH2EuaAb5E+DtQhZojaOwcnOTO//ZcNbh32D/S8F9y0
CoCLtqOePR0nqV0YAwS21seMwJlW3OyERUu93f5TXddt3gOUJs8f5a/3fxpWH3Xh
LIg1BiS+uiAoEd5GRxexDpEsWqf0pT6GDqHA4z+WRlWL1rO6EkGZcJOOE2ecNBWP
65h5k0MAcWYpl6dP6r98ojVlLXZZsMS9JxSDBhj3dfx7dpLEjQTKSJRIA3er7Zku
GlfFcsO3f25WQWDba+GDiDOXGNwYvURSaag2M8+A3WJ/TvTOhWiN2WLSl09TJd1b
v3Av2bKnaan4avkDBPV64x/EQ3+Tqp3ERkC44lli4OA7BQIg6NAGCy7b0mh9TIxP
/nXNUxAgL08eJY34wQunkYcrmeOKW6AhXKbBd46azUcJVN8kq7bQt42VZT898KJY
5CNFj811jUuZeM883ermxsRVVR2m0QIIz4sIZmdCfcxQ6dd1XXNGBY4pv8s81cE0
OPkB3BaA6F9XlB/66jzBz4RAKE8k8/29j0TrzdGTNX+KwYgnZvgioFNDhurq0VWy
cHWf7SEg2NWH4z9SFq3ML9xM42r8ic0NSpnIFt+tdSjdA+EjvPi0Nfn7eay0LbVG
AhZYCly8sKu/lTVdFC6c56AGxszVJqVoXqTcqTlAys9fM8RuYPK/vuZyBoD0VcDB
CKpIJmyAZDwhmCos2VxRceFipcb7vbO9BgsaYkFgXkoRxY55FhyxmZv4RVrKhKf3
ZF4lclcWJjwVzNBwEUkjqdOpEGoPBu+SZ9yZiVwu02kMjIp8RI9Q+YyxfAAwdcpw
zW0RGWZjWgupXNbvEeV0YuFH+KH2po1VjOFnrr0Vj/glhSxg0ZZ757UFW5UUK8g1
HOaVYqTLYm1OKkEx1JCMR3ODkq0ozpJhoU7cuVtzQ9keWtNVFgd2MkzxenZP1imF
Hy0i8DpD5qf2/E6Goir1K9md0I+ni67/N7eWvJwW8mv6IWwdYnB6n2lOdGWL8kkl
f1FW/89plj/ZHhQLexyXUNa+nzdVuxUz2eZF4wJDx19S5cEIclSFLuPXJfA/Hsrh
S53wiX8j6m9fieV1q3to9w==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BkX9/rGvwmK/U7dB4koSVz+Uv4r/xq8MITADjzJVL15+RqQSOoYSY4OFJlq/SrZM
3dxXJKExs0miYe+lQ9fWifrlePiN4ClX5Bq+m214Wb9RIfW51h/WlX/zFrG+9VR/
gJwO4MwtpsjOWMLm5Dt6svzSDaC6g6swLzimiSbxaN28gKSUO8v1iskv57Y/oSr2
w8msm15Ae8naq/rBfwkvZJJ5FFOKSpr/KLxDV/zCYJqEvD4yvowCjKj0j6JJ3mcN
YQc4JvUaN1G5VGxasTwXQZoyvXiypP3+ODlm2cpT5RWFMLettCzKh4oXqIfcSaha
6Pahoux7J+61xIEoK8StHQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10640 )
`pragma protect data_block
C7kvCawL7ASuzxsHC9dfED57jr1+j9lVs14TtbJDVKJAJemmFs8XPEIJxNdDHBI7
XrbfX8UccYgSTWpNlK5iY0/Pauc/3QvsYW0iQ38oiw0cHHzOvJsRsNuv58KcKDWP
ewbOQCvvBYeyreKhyRak8N5VxPAKLLjmGkzXB30C6VKJpUXMO6GmrK0ciKmPA54G
V+/CoD73qGnohdSqURXMurG1DY8E/ltcN/u1WNQP2W8VoMxLbF9hykcC7n9P5ezU
nMEFoK7Krua65O8YivqMbMyRp74+rX/obxuX3t8DDyNXYhIu8yjKb//64wPo8qxD
eH435F23mxGAY9+H6JtzzjPBp1J1ylza3ehoQBePdXNWnQ/odCk7znKZ3FU1G49u
IvcFweb6vJ2MVn88useAtvr5Kqso+FehpaRVGi1TQjdkzI9p5b5FO9oCFm1iTqof
MIIrQOSnRy1tbgJ63FFcPfE4ayWDFxHoJyCNXKv6HqAfVFazOmwS6RL2ap41qEOg
IcPH/sgOE1Prm2Etmj8zTfJdLq0rx4KdW6FdVGUrVAN0LsS1GC5FkhR3nBSzv4aY
FpTw5Waf9me8hRiwRMrwDsXicXGcrkwQ49psLMqVVK5bKf5lUke0uUTXb5IZ+edb
7tqd8Oda71yE/Ur3pS9I/FgIyCwZMmdcvDYm1SeVbv/reOlmE9d1ZpTt6VjpQvri
95mFWAQiz3x/j7R9MBLY2wZlKp3pdIIU7eJ5zA61A5JavlxIYlVGOZl9qdiZ0ByO
63GmHK0K/m2d9pQB1xabSipXoTLpbW7BQ3yNJU8T4qqvI0ny0P+wi+JW9bNHDxKQ
5xGxqclFpBP35k0LlmjbTgESiCEDf8lP7keefuv8BdNoGoWckd8ugbFn3XJETBHi
tovnJUBdzAuj41R2OfN9ij3rVvVWtxV98iMMnBzCsfHK5yNsDoVH0fCVl/bW03+/
peATnboYHKIOO2KTJUM0Spfzqw+uJ0VwIJ0z1K5zQWioXoskl4per4Ylovc935DU
sZjGaNjHZX9vLoAxrjaq690UZk296779s5/ZMElxsDHTfvkYuvrGByN8ZYlnjMFu
c+uS8oJ0J/F9poXoLkF2nHNUUJJuPzi8zCaajaHfa3ZfhTSO5+GqlYX9xgOKYbv6
RgfUyx1Vdge5mZ/6MVzMnnnxKt0DDn1ppxJRGqNSAq5Li8zyWiFhuIF/RK4xcOVB
5zUadfQUCBrJ1NnYjCqPfe9qk533ZqUcuh7XpUrH1pDEo5hz4E9or6siow9iMdNP
xBCZ6L8ftcd324dE8oBeOB5x+qZ8aAowb0bRZ5jrAFDPyVSa0j33nDNAEZAflB7j
DEm4oWxhykjSx5odjAqa/5lxlpjVKoCk8jao6xtQYnndFXOeCxNGYTnwHA/Zo6oz
Ftttl+P51P0uO8MTjwaJhCBd7X7uBM6HXry9zScDrnXe4kNPT3SG5kZwCHQC90/X
46woJ1doOkvn8suD6YH7iCN8fwMSHSDMv903YRXFlZh2uulO0+TBQk2WcMSTfnuv
kNHxrkhgbLYbTY+9tTrlLdxtATCR7tR7OQfkUI6tfOSUZk0mJR9tq/BXf2OoW8Y4
e5wRGJQ6B0FC0CNPeQKv0zt56Re+QVkgeALiCPtkCxy89jyggnxy0J7CJ0/E+88G
C259xgrQA9I9Vc+nj2a/6c7WuNVM8BJx4TDGEWWBxYtNPAWzTIB3nj62D+xx4lr7
ydqW//D9X1YOdVVZdxMZry7qJwUVetQDLKEG7MDBAWV2i17id2HNELbE3Jsh6Ukt
uV6pZ91tqYPGy3vbUWqmKcfWS/M6v197kJBdmnapJLaN9pErn+xefSHVuKRPy7zE
5hH/TiyauoJkUaObETFSC/71VjsUJ3Ba00AUNbvZwZj1nFNJgl+6tl558TIuZv8Z
ijzaTHj+7vbIlLC+PTEBI278oJIn2r0dpMY/hLMkz6ZaradzsL6esZGwaya+lk12
utY/briWeYDsGheR0QmaGerVBliw/yrZLR4vF/E/fDKi4VyG23uDJcqBJfZvOKtI
FqpistHvyBzHvSLSRRQP7glHuK9SzbPY153Sfdm1+9JvNJrcONMYOFstGrOskof7
/vRrPi+x7JcCyiDBSWUoqdObVnlmMxpBn3DNKKwlQDxRS2U4lmA+Bh4QwBP5Jrnt
Uu0dSYDgPqycQwD3XajdpB7k5DNlIz4cE7Z70WNCgUVSH7Txj+fN51LIoToEAdBU
gmy9Yc1C2iLVk7NkE1Zqd/knuPcJsPK7eAiGK6KAVTdh2N6DODJBRPknBlb0vd3+
PzTdVsRCguxOxjGZcbhfIaO1UwO3s4HGLTCP+/rs6H24kCdU9N4qVIYrjuArJiV/
TfSXsXDNpSI2fX2g12TqJjDTrr/pwZu2APmPK4wq3BrDHtXdeFASskDaHbE8t9qR
oTtdl1PVjlL/SiuL94tydA5+ahFppOHRrw2f8gDpSfAoqix6aQ8fHGMTtot5GJyg
V+rEq8v5zvllgHIptWy0mWr5pis+9KOfYTBxg2PiVnZ8cSjz/1gHpA89F8A7Uako
WINPNz92lkjsjh+j/9+ZeEzZkaL2m5/cnTHlWHatvn/wVknppCicoNNrzL/lX4dC
df30J1U5GYru2nj7SD1ERNuGvteNXVCsouW4vzkg+7VmbOoG13WElj8T4nb96VWO
j+dV/YtBJduegSukbotFPxv0h+wmJVhBR3jzLD2FOIqNSytPf3R/GIfeBJLvla+h
ka4Joj7vMQgnU0ls8W7w2GTMIFXra0fC3UOjEhEcwL+y6LDEVEvCmDxX9siBnGIV
cfezYvPE7GM1gVcVbTQP7yjkIsu+PwgcafAKrVI/eZ0tsCY2d1zlFoFWo79gOePc
z2LSh3sz7y5pXyXPCOAwRvXgELqEeK3pDQKSmW8x/XrOC3fDmeY1h2M4CKz3rZl6
zoM/SeN+S64tk9DbeI4AZPJGeVLRlAJ1W9Ozc2/fG0W5fgJVWKkrl33AGB5Ap+vt
H1WvJzj/IGFlctBOW0dLN6tgKnFUZ+Dx+6NOmiB6/DXb94WW1JALxF2LJVrr3nJ5
g5IvLGlU3wt7PizzsejwrWwgTZgYIVWrDMnUjYJc2IMau/WvY5167v1Wez4PbTdx
M95N7Irki/S3oYd2XzZagGZZ+krtjwQHB9tUVqNMNaByasUEmIL7+hb13ZV3eGai
7Q9pk9C/tIVSrK4cvckTlm1L5aprYmY49S9PSTP+21ul4YZVMGUu67k+j77C3ZP5
vuOcHZ4VLvu3bF5rQzbwT05fc7U7PtGH15aXY5TOL8PsTN0HCP2hXHv/r29ptmVu
NvcOfZwidtSpS3X2hb/oTDxL6Bj8Nf7hipeO6SIFxEm5vgCLfOuXm7QqW7Tc1VPg
rVgH1+Z6EdZLJegP6TFvrMTJY0zwLkrWkXVqbP895LPvv4mhinNGbb8Qwd1eBYpZ
vKYQu1g8/LLr10WQGwkntsJVhunFL6TOcwHNl0Tr3Pj+Fb578erX7NF5fxhtkkJG
xj8lD77/Wwv/rqpAHSQxEZ+47xHaw2QeTI8DQT2x23wDI+X0N/g2GwiK7ip+E1TO
w6mwHmPHkIdSsKlIaBl6w5flc/AdqE14TLIlIThRt+C6mib55sHuvPqXAfTU1QqO
9MHRPlL0M8GOhctcntEk2mcxIFdTnmYS/vvOlvCBwQb+uanhtoTeUkmXyRoizzXD
6ZuKaMjDXAxzzEvQZl1Up2tMyaafW5m76tQRCPWTORiFki5dGm9MNz+cGRScMdhl
zv82lz8G7eWT1bWIznvg/rBq7naJaajzlHDvdLcVxU7knboD2dCJlPbuj6S6QAps
Vayma/QrUNcJ6Y1ZB2wrjHpngYJqKWh9Ev0XuMj+c6/bNM6+exdZJpH5WNaLutgg
mfKfTLbLbW3TanJpzO0/4ILmpP68i0XRq3fvEP0e1zvBJpbH+P2pX82h5HQNDeyO
kIWoZk+ioBXNYWgHfvi3c5OTsZhiIlfRwxADBsXuA2b4LWsu5vPVV/cpYulrttrh
6SBp34i2gKoPm7eX9i+pMRtNpYSF9SWDjTI/WDKxh/9cqmTS440YRECG2Gf/hdhp
2Za3voxRQA259N/ZLxUBAcrkos0iuJ9nkhuq9gHgsqSzf3YmUm9mlMld+4oXwhIF
KEyj02M7fhm4/q3kHFU8kmL0bveaeMSVyEfQOBdEZ7A1C0UThLQbzEns/e6qyAoH
Z1plRS1RjrFSBaqogMtWTicOItnKmXRU6nskK0zH45dHfc2/W5ZiN1zfuo9te3Te
8/7xNkIudMStBFDlDWGgPk/L5saEzTig0slM3Ui7y6/l496InOFjB36veyTl940X
4u8sKyCtTe3hwV7C29X90wg9CGcZxxVNOSM0shnBR+qXhccJqM5DvcyogX0G2lZU
/jsbk/fy0+AU7Iuqd2B9HRcFOQ0FFbaywEAneE3DoKgx1RcidZ8wDOIES+CMZwfY
ITllkqO96W3tdjwibm8hjuHRFCeqaHxpeabg4YHeZDmKB35CpfEDjxpQ8p/eBKwo
6WULCRjxX+QV9MAxB3zVs1ldM4Uswn1flPzoFlWiEvIIeO49fmcjc112f4/HcReS
yaf1ckSwosTTi5ykJEvUc+g0LE/B0sTkM3tvTPQ1giyeMXl2a4/Sf0N+8xd8y0/s
4kjWWPg0erxYHw32vfjz5tfXgLfPiIJF4KZgXV8BTlZUHNzDpAy3o80A6m2Vwwm/
GwnYYWK0XeOlUNIgReUV+t5nSeJdUHq0oK0At8+6DZynAAT4dM0Rll4UC0qHaML5
AcxVbvX6TSLzjkWMvekj55Nr0OA8VFQwMXMObncTyS1aVUmpIhqeRmYYM5HhqCOY
k8jaBaQEKCczhbf/FZcIrPaH/6YdG38ZtTX+5lZSqLYiSmHmZJoUIV0xNpY8o/8E
xHYQE9IkuIJgcO1jg24k3uUB8UDNEPhnX9OaPwHDrU18O9YCqoQ4YWRR5BgKPo5p
FYvALILkhic9TeruVGr0WoVr2ccwyksVLXNiJTXU2zx9TNFCkiGPz9RD/mVzMvnN
F7bV7LXaryekF5r3iqCP5/aeNi7uc8lPSlZHuDnqZ/WQBjSvXDH+KIyeRZAY0nnt
0p2qtxsVFY3pLiLkx+6jZl9Nim7yPXSpZlxBwxtwwyjZvhfitIMkQLemc06SGX0Z
FLivVQHpeQL7hdlfzAhYW6VesSqono2A4+/XFagPyAjk0JHXkbGjbgDd9HBvHYQ8
h7+66tnslq11R7+DqZlGNm1ppzKC/M8W585dWBgdfOchJCGC915sTTa3niGXdH0g
NG9WU2cp1wGbnP43QzVDtlME7NU6KtTfR683OJ15Gt6T9ZAubfy9N0V32acA/gLH
+Ij7HdZPuWKQiu3xgWDOHAxofKAfrtibZceJRQ+pFu2kBweHFBpkqLIddkThpi/v
E2pfhK7fREWW5yA1MvOvX1LNpcdtll7Tv18sXs6KhejotOrrk2Wm2vOjY0Zx7T5u
3v88lSPiEO96ZkUiqkDhDiFsCyNiTCqEADfVLqYZEuCVb+1zg7nqD86U1v+kdXx1
37kP5A9bMDjpMRoEE/UELlu1UOeYf2ESJvF4Qg28PUSsVP98pVIERBfdGSCWWE/Q
TZ7JSZfMPHbXWFiygT4I4PNoQcReQDimZZoc653r159OPo/b7KMDG47I9jsJ9eRG
nE/EX4psX3qlbi4FkFfduH/IejvmORB6slQa/TkucvNHSnvVTSDooX05fZylKUVN
3UoSidTqmWzeo7L1XvbESSMSZEFksArOkYAtCHz6+R2J8Oto7nDaN8zxAndqV27P
DQYN02aRGSj6yHBb0v8oS6q41B/9VYCTYZLph8kZmUm8/vDMuIQQPtV9MmwB0yV2
lKYatwbmUmwNA3+AO/mKONZVsHZfF8GsgKGPF1rUw83kaGWJ7p++imp3maLB5M2I
XrtGDscP9ZljLSwNZZGQMh/a9Ky6XtF9g1u3AQFfU+9E37nbHJYmhQ+/O8YPJUlZ
TvSf7EEjW81GZe+/vf5YptnLQIueeX1/Y+O8yD4d5vpiVlrROc9Db73aZHJjCH70
uDh1s/TqYiErZp69h1nvD7yq2Y8tuE4vCehsNMhRNnvR4bZisrBsEsox/UppcGMn
4uxIqeEWCL6hVTFZyqhEh0xo7KwrWeqrnPPbINUt5ePBCr3KqXpNUTj02/qyixho
jqiC5yRaOzMTDRv1xCvB2OPyHkSyzeAD6rsaWlNYuB1FK4e8FLu5RBcytYBJJLHE
qYSCNwtGzRIuh+byuBOds66ZRd4uNTLHIcuRHXAi1Srhi9oPIwyHLh3EzkeOudHl
tXMOQdRaDdJADfj0FSpiLnGlYS7ObD6oz9RVBXGhLoAAgXdYKm9xT9f9bUt9dOUe
XU6BoDwxMS38fKVqZf45XMZuNvQerdIZEEnjeYsQzerH8FeJr7ANQJmIXJ5B7vqp
xYt76rbeOorZ6ThyiUbm25840a+3H04kbg9EaqUvBBkso3lp8Sd+L7eua9sBc7MQ
ahsdFQcpz74hkPHWKhPzfteucbNA5or8EoBQwSDXjKOS3SBHEQG+btg1Rbbm2wTi
RCVrRu6TgM8pq4vzqG2sLbZaFgJhb6QbXifmqNglRaIuSwVmaxZC/pORarqVnSi7
RxExcCUTFaBrRLpsFUWT4vlrHQW5Co4FAy1BR3wtDyTPLyoKi8xnuks8Po0sC5gv
MU8FMpKpLR+71OTaMnK+5krcMX2FILpJ0vNDBenIWZhNpD5rp4TJr/n2Ik8p4PZ1
H0VtqhNLoKem8mYlAzy2dSykFIO/M42wkOAArETYaZvIX0OT1qZQNuhvfCypFLOF
5H9sVzcNyOHkKuGuOcu8Jip0U96fKgidxNr761npowqp6F3makz8nJ5C3bks4+Zw
KDY9QwrEWFI/MfT6VjxbPLh+BLifxdk7CFXgkbwm0wuGusHpN3196BIJjtRU/tnW
PQ1KeiNTRhBkFkEh1GeBMh19cNC7j2nRF9jvOYLiMj6yD4+MxjvFQIuzbtbNerGd
G9mUqfjV48LY/sQcqeVX73hggRYFbm4gIDLnY5UoOiaqKVrwogzAzyn98tlJfhpU
E60NalXrYQZcQFH2Z/gp9LIsqf/9azA7d+x3fPISK3Vu73TxNMSOtLm8BFeHFyqd
nME8R5+PLm9J5vfjsCeoVEPQDt9gLrC96/6dN0tnm3d6gm+1njyoL3ch2VoUPekl
l1Oc/HkHspR/3pJQVInnAUfQce/HKmjJ8qCwQTqRnQwpNAL840KGAsh6NiugnSE6
lmvMir6xsNlIyk3T1DfFE0J9GBn086QwKno995fM3rODfeTZ4dxKKIhEmpCD33iS
+CCbQuQS5U1sR1rEzB8dnYqq6eqDx+xQCy0QP42lLvFyBxWvZMBOZpCUeKw6rDv5
L+6dgl99AnztD9UK4oYSwAemQGP+75hQPR8+4JWGeLyds0asV5QPSdP4qksX2TwW
UqKpRxAWyIqy2OkbANlNAEWUK1Ic6lXJms7CJKZ51qeywWL/2lW6wAQcGxId7WIm
wFXRYWg2bckbS9iWiHQc0QaqHxY4/IotIHuDRmsbjpeLYrdnonuNZNm/+wipeQQb
c/JQPlHJshH/HCrOMklV3B4N3kbQwCD9KsxcvBikxOm6WnbNk9V5v9XhBgyUjFcP
8G+HsNT2WI/V3diyeBxeYV0foA3e56EIjboO/Oma3jV0oVu+xlJXQXNR9n0hid27
bwUI/DXucNsXEC78celsc4xprzZ6515daqgaBss+gE+LOmzfwjv7l6FS4Fk8zP9i
EiSD3k5TDCApUd5VqwgnvqgQ0qbuzAbwt7UDc+pfe+BePLfK8vnpwO/T0BS/DbST
qEOMVzxf3puccuMHbmlMlZOIildcpQIudGgydGU0qeXZKmnmcXzdCClrHkEJSz4U
sb9Ltjdjz260/HBS7Q9hbXf8FEvBCB9sEbV2U6PUiS4aWLgjN4naCWvf7f00WMJp
PbpaGvA4hZoTnClw7YlMKy7b2OKNsTW6v1ZqsvmdfLsjGu2KH34sykee3YCSdDj8
et/5vmBIqve8FFGiWOVcgcNef7UtuiOZfMd7Ko9k3tFk024yJ+kru40UrEcYyyce
luZBdGNqpQxzdDQpVYrsUs0/OaqYv+N4C8onkQjR2RxxwXolpxyAWBN0qXdPciWO
StSWQn3XCP3uOppff2T2sn6bbd7Xwft1aobQsMTamdn5USeJ7hUVS20n5xGZWIqj
vXO233mNlLZpzncPlgR17MNxCNgFTn1gUSO2wU2JvUxTSzFl+Pv5759NczF35ND5
VY/ML8JKzYry5PEACmXsz3faDMa1CCNDR60TAShlYLE5oyIFaU82vaq3UW5+JRgs
Gb6nbhrLliKfkFQ6jLBAuu8b6Br08cL6KNzvySm3FAnmBFHnKWDtasQT6AEPxhc+
m4f9UvDFDWPXvIbqezjaz/3yXqGvB5WzdIz1Wseo8gdiP0h2HCJ+GgXUAoFrzrDa
5/elTfIc9M3dkce7tXOknSFaVJ0kK4V56c+F3HWO7ClDQDengTDY/fsfKYEeXhK7
mLlDtvVi0A025hBe7BZnYd2GWp5dT5couFEOGvoym07RcS3iAA4AM/zi9Kj4bBD1
ADUUO7YfCyaRuuBubp8feRQAzi108mcv0WdcZPKjXOnax1pQ0p0ztOliOo5wy2Io
3pqSCnaokkJHt+/CmmDskcS9ti10LhhIvT0OtXqIqq6QHCtpiKVd8DtFytCqL8Xl
PRqvLzojBHVg5v+nqkE/72fMd1Ic1D6pVdGWBVMoLvPy7+FtMGTeNF3NNWFIulxQ
3/OGv5zAGjZTRr7MwJZ6vJo2PqhJoc3zLc4RkgUnNoNiMy6cifcOPbI26KQ4nR4x
qFaOfO5kdq9uha7a14se0iusMTmp6/jalzuHrn2whQ+yGyLLqCQwwpG/y2zTtrJY
Q1bDDtA37ON6A+O4Eu+y7KB/5rDtaIgpY2rMB0LLb6tKiYQhvtO6eBjjutkAdKem
OnKg81uynMM3yvl3N8CQOWWTtw0c2ml+FWW337Rk7iShdEf7yayb3DTt/6XU36L4
Tk0barGTKR5ezQBJ3qPaMSbyNLbWJfVqp5+cFGLtKrKVSrTUDxeQdoW0F6TayoUP
DF0ecL6a45pnVxNUqQS+jBTjJ1NbvorLSupKyd8qTSq84vDjiEDEnKparmm5qE8q
fFtTTVTlFKFteiF+umiXnM3CiqnmIRCjlc7lG7NfiZcqIEZGFMgCxD06p+7GewN5
ZrRjLGs6yyfQpeGCRfG5RI+rDaOOaF/R+2mVLZWbzOBuABpnS3yu0vv7+k4ZVsqe
8jZfUl3/FEHaLZPEFbXU7b5sxwqeO8g/pECbCTSSZr/ObIFaA2iHRfWQ77em4oiv
7xx+RHGJtfuORtyMJNse7eatROBF9WveST2q4XQML7etLwgn5yDsGa2wYHT+kV6J
pUKIA4IYrfuhi5ux6BWO14qOig1Y/shRfmp8TfZ8wIOtKWi+QWflQRt804lOfvRW
VIHUvWqXjl0sYpGdhb+4yvftY1A+pyAA6lj7VbLHjEXb4BMs4xbtEXZtfEhp8Z2W
axypRGvNyOJOZWsfAFXMYXemtOoY6q5qAHcFRACRC4GwZMvYwTgmFpG5RfdIrhNh
uQTADztFcdxcE4+tPxj8VJxTGXfjWmHrz7sn/VZHl5WhF96KU63Z0eGQiZ4d6lMC
ex4LQ7gpZRjkrHO+p8ZCfBgEqlgt/4u3yhXeFhKknYNpbszB6tmrqlxQ9XwUoIe5
Q39ZaWb5oQJ5ebT7axKrZ/3wpccCu5NOE9RKZiMzKH117Gl4fuAIw56gZmqRc7zX
o7oF5eXmxjFDna4iAqoKZhLWlrEPyZKjmLBmw1t+ufsKuENbeoM7c+u6c8MoYAbW
tuYlek5api6xERpozr1XeEI9SVPLYYRtYv/YjohUtNqwo+fiRAxEZ5SDJOIn6m5G
gGtS7u8JgU6UKTxVT/eGGirg+cCAWaXCb951ZwVLUcnOXdojqyqeidAxOeH48RRm
oJSWekH7d2N0jfHN5JZoEDGyKHkIWNB7kFJ8BCj43gdJR+yQnaTAcNqGtMiOz6CV
EBzXGIQR69coBzfKfV869Ly4zIxK0SecwpyEvFzrqYoIRx750Ggw/VuSt3NnMTeV
Bg2b5T3NGafTD7a2epyoD1kODPdjHeV9lIMhXcmrI/PDveuFn64wLnTle44rfasz
uvda8K2fw7WeULGSgy0F7NqXWAlPFw9jbRDm/PvoTgTSJhPGfID2Sa/K4iaqbW2j
6XPP5fNpSDi8+B0xkcX8eSAMpV1d/ZmbWuDnq21+LlrksMGeiDZrzd8+ruhCFItN
MB63d46A9sERgDnSLkh21gwZDpTuKJKRTWOU7OMRKnCtEk5UOOjvnRd6gvc98At6
9hg/yRivAXrtZxkDG+REuwXxV7BB5C9sFOFqLZsFGTwv0FZSc//Zbm7YJgJioNk4
ZKO7hGOZ6Fq4/CGbjxwzwyZp8bzn6eRfvtSY/VxH+iYHtUvU2yltJTnjhlkOtSFi
uKJQ8aLP+keUpdhrBor3kTqFf/XoRkU8wVeW7wGoN3WTOlZC0b0PImTCJGTs4L5/
+wu1dFvrppcxY9/lMEqvjPZirWgB2n53dFccKLxLF7XASguLufiSyjC3f6aRVOv7
W075vW/KdaKINo6L+MH3QtkQ3ySzloZnyRRK3bFFT5DW0YJKNQl5tM0d8koUadaP
5UEnJWdRiBe50OByGofDpExYfsk6OeSks6EpsTsgdCE40+jyZd3I93UhmkwY9LBA
PsuKvY6BoSk9HCcjv2mRnawOLBQtzvSWEGU2I90wrKCCC6llmqCs8AEvQSyb+fEx
tKywPyCnv5mMiX2gvMB9I9R/DLdj27ejhJQZL6jB2uQ8nCwu1jyKK/H99YgiwAcq
jcZsF3Pp2HoYafdzguXwU/zmTSro8dFwNF/214BVqwub9SWrgLsuM29BbA7AJv1i
IXiuV3yJO2Gl6rm8RiRIWfsUzkEZE5ssij+zgelfRWAtaPadWgllPKaAcxJPAmsA
mfAb2BPOzONJmkYwyO/DGbMWbvBdesJC1+AtfjsGQ3SyYoPU8mAZFJOLMDBjt2mv
URjCQhXGpIqJmx62y7i27FHo/UVV2djjQLm/NVhroo6fYnnL73PTgzQJ5AlhTA7R
il+EYge4XBy8rend67YBh6nWttlfjK34GuwXp+P+uX+AvvWENV6MWRn8gHJU+s0+
htJv7uXBiuMlK4BuyLTyIhC4wfNTrYWUrUDAyVgsjo2pWGgP42Aygxq9uPCTfpBb
IB0vcSMb1/eE9wB2pnrLdgXCr1GVeBHGHE+EhI/8WC/u98WO0EhGWvcDdzHZaO/2
WGM+y7g1qEj8Xhb77t58D6iTw4X1CV5hEigrzwhtqSjqVKMtk55QgwrIt00M7M4+
jytWB/SrGCNaC06spNSFqAQyK9jf4Am8opkedEvXxDCv+5pjInS+RwkqyhP+yE25
45Fdr9WYZMN0AuB0jYFSArkurhJvYzkH8KqsQHvisyqtZjtyGJvy0h/1h1Xdu/ly
dJRQix6+EFHWkffIrDVjNzLHnx6eHxmW5NkZ0Sbmo6643D1PDFlAfBrXc+54gLxU
Ch4d48k+FP4CpquOK5jenQlg4SggOIodyt2a30DTjswocy7bjyyukKl2+IDdYyQH
S+YRmDOdVTJQ669kXlm01gAfUXcU4DoGdby9X4QXqP59V+9DLJNsR25OzOaoQQJq
6MZbgiS4blgXqJK6Q28Ekh/wPJ9eB6yZIRF/a6W02ku1SZcpOziMesfNgmG+jQ93
P3RSa2j7JmHBW5JwGxM4AGXtuR/7YO+76p23XYSA+6Bzvtcbb+Kc6gflOsNTZCZ4
EIQDb1XLOtuT7nqCmCY/7P4/wHLCmFxrQiaypxH+//YgcT1JqZ+PbFDKf8l4z2cd
yR6W89Fi5xRVQ/PvVgb6VfCCHxVcO1m0daJznFnczKulwuqMw/OBYunkHtR15/Wx
uaP+TGLtFBkLmWp+tE0QDJRWoz8VhFHIxbo4peZGbMQRMyXCO+BgL74u8LAkYCFK
TmsVWetOdZJmjYZysxcBci1q886zG5/MM+7d/TxBxI4Eb6K2VsWnBV37UTtmqHDo
1OoXwX7hdEqIC8CGRwNIA3UsRnXJq1d8I3icdpABnGmTrUDdSSbIH8ULrt7pa78V
axT/DNlxQXzduefatPjU0knmjsSMSn+4LtGs9S7Ip9zzGGgZ01+W3GYNyfYr6ujn
VIEH6j4tr6/L4SayRjhdBhyB+SjRmPXVjlcE8IlgcybfP8RPZQ/xg1uxwl2AE1tB
xlnEckin+OM36RhcK0RXZzI00kWBITcTtdZKYllmOZg5SYHIQ7STVrt3KbkiyQRd
I+WYsqe12dp62bu7lP/jaKZvDKYMdcQuzE3++Pqqs6LTQY8hJlPocQIyTYSS5lRd
/af7eOYAUqa9onLlAq8bxAp3JNpHXTpISkLMd5oaoON6RjXweF3/I7hYYKsPHYKT
KgLJpZ7eiiqOHg0UTHIHMRCZMJIb38+xkYz92fZg/m2nIE3EkLDf0kKo1OmMeGVi
+0S/Po2ykKQKxVo9h9tw5rvzPPqhDfFe6JNZHJOp8+ucgII3jYv+RwLArgQB3Rpq
+G3gIbk0o0VBgdzYrG11lzS6CLswVzUcn0oTZbL3KFiUazp0OjKep73JNSZYSB/Q
HHL16sYbWAkfwx25Uiht/6/9GpQFC0ghDgkX1+s4uKejLF9ClxhBh02dG4SUVS2U
6mmWs3TPc/8Or5mp7Ed/gM2x0sYVXRJYoQKfrPzugT3ep38wXJhRuW2RrYzVHcxY
8OW+QaFNDwL/8xqDq7TsubxYHjn0NsOilIWHgSx3c95OeKH9vT3LdrVUhPKRbkbh
kaLBB9gUQJQRnZtWlwlFoh/omBV/AF8Jj0tjHa8Jh2gFxHxV/ChIWPuW37k4gO6W
ZU7IQU//zI0k7GUN8EGSbhswZaLdRbszttLV8lrSd/f5qrCAJiG9E59YNdLSR7kb
ulUq0Ptg024xvqenzyTpJl9MRm1B6OnZ84xoGjEEAmHKEaq1kIDQP/XCo9D1riDP
30k8C2g7dwGpmnXrcjw23713QzgAwxnPoYy37SRogaPIHjnCdf/e7GmWvLGOpeK7
JwysH7rM9GftlpPF6JmnwPfMrgbSfYsVI0hhObJQg2wu3FjidC7E+U5LyXPG8i9V
rhyzLnl90XDkVaEOcCAaTgXeekbzUXSPVfUCLQcX4hi0Mk2HNZo98FmRCpS3cUz1
AhUznOjI3qy4wpoVXnIL3rPxcpD5iQFNCH6WSwtiKdZAsBtENcPo99BfiPLwQvhf
qwTjrG4NnSMiMmfO7l9cSrCnSFar6DZZBBFePYVZtZfYe0qy9+0qMWm5YKIGUb+o
a/SoLEY7lJjncNp/J1EEuyalOG2M6KKZtwNM44VJiqZAwM7FbHdoli5KneB9ZDW6
YHaY0LFaWfxmEiKgQQeOovz9n7jnoubE2b+W44G5z6lv+vM6pV7nYPPLGIMOM2p5
k8FxCyPTTHOg8DB7AFqwPP0U2nfoumePnQoa4g90RlwlgHSHOzmxZdWGPyHTxMjC
01PlQgaSX512/bFIN6q38Q1JvzyKVVs8E0H5+yV1m8AW6gm8w4dnXmhzdPJasKBZ
W82kO+Z2Rc+2jFcS+nbyHyHNcIvpAQqoYVAcfCYMIGaE+WB0lOgmfrQhFuWIxN6Y
VOHe/+Bo/ggeGVtZztRLiiEn26kSHoQBmEeY+amxnwkFaQ0b/qakfxCkbkEh+QMZ
tkWqLfsdk6MHJji7e7AvMFJVniTACPSfFjT23bIcEKz0+lJ8QVBnRIqkwcxOU22g
5+e7wHlG3BEv7kPtrWk/H1o/jSfzSpPCSc92xyKgdi4dGAEs0dwszLTOZsBNQrYd
ziseqZB6YWky64mspk/qOMARVf2EipggY1ks+rGoYbpHv7ev6p4RaozCp/dZ4gyR
MbvrB7z4VK6MNBmHfv6mL6Fd7Hytk0Dp903FFOn2wgSS7NQvuNJZZzM3WhQoydVA
p/7NCQkA2qlvIoJSuLzg1Ou78XizRHBxzDZPKulQAXcdX7UtZ6wye5Jf0R00F63q
O+ouHMJVS7mNJFoZP6f+V/cAiF8Jy3X4jN61RQeXC18=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jC0L71j3qHC3P1JuMdI9in7aq6I+zRcysvN6ql24AC27+G0OhyNViqJqJOtAN4gB
bO2vl7WHj2qwHyfetJN32xkt7qfyJEL0nGo6yUwbWDF7XlJ51V19ouW5Jqr3nOal
TnpBYYaepcVqytGRatOOyEvT5/1b6l7C5L7FerpLuV8RCg2eTbSbi2RoPJA+x8kO
L2pF3oG6r1dp7PpV8zsk8D334dbBfnKnoygHPnYWjmEfjc5VA1k0DMoZ8FgpEpcR
hVuwh1nrV+Qf1AT4PUgwPogz3Qs0VD6zbUIr5VaIgnFxZGt44AAJH/fUiOsUCvej
bP7O2RcSivH73JGFrOU/eQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2704 )
`pragma protect data_block
OVBCqRpU0AwqW98UgW5wNgJSOH4cmEAg4Ko3EnYT9jZu5zxW4p4PMDiDhh5q2ShL
3phwH4JJHuvW/FV1plg0xQj9I425a7k5zWR2E6gY6um8bTooLJCLmCbvxwF0DBYb
FIR1tE4FsCgmAiEJCC0X2Ey6Ggxo1zSYOLO6Dl81egKA9p89ri7qpXfR4zJmoXx6
BXPy2wpy5g6eA6RPLuD4GFZU1Yaaa+7z0JPamH8A6xrwAJiatge/Vc6u4ETCAoyr
NzPOLZ4O/FGReeEZp0ckhLgWfR3FQx3iQ497xXSFDbZHeyjZaJ16dDcxQyIzN/MU
RJlX9ujjqrJow1pzeezYUMw3p5QXTJY5Os1VREexXzw9T82CqvI6WjdAwjAcA6RP
LcvQL2NsA0CDzxpkkhBmRrlr5bCzQQ71AuEPlC3uVIn9pf051xniFWgH3LAl9PQ2
Uaz64O4XcaL4mCtf4Saaf5psoq+gKn1Z71xZJ3j5ZkPpT1n4PUSlhPiq7Iu0m6eI
KT67lA9utcle+yqtCIQQ2AcBmxRA01Fg1k4XYKHSkovCooosQmJWzm8isN6ECU9z
638Q3/jEqVojIDbtzXgXMKIuvcX9ChLrr5Dnylkmf4i3045hrTwCDdtm/VLk/7rp
OeAa+PSyq/rN8mycdWqdoUMd1g7vEgnby6UtC84GEa7BC7YL/7vjy8FEc9rKuq8M
WlmxaswBfIC5D3DJaJ2Iwwio6xPWIuUSdfvjAJNIYbEpm3oTyrGgL9SFoDE9gADZ
gAISQpNnd998feAyDVNAWi1il9bxm4ghrGaG5JfMoxO7Hpu+cxLT8q+TfzKlHHH1
FlTBOvuDCsdN4LcES6TbSoBnQf/A8QLcXj8vbpS/5ZzaO58TbKA39w6+4BeJuZ9y
r+znTDSh1WHTUfqQi3MywO5lXEILO6fufbXmJtTtiEqp4exFb5yaMvHNh82yZzSi
grELfkRMx/mSsAzKUMph7Qy9EEbHXe0dazTr8Tbj20Tx+AyqE4oTKJGUF5/LkPih
yQBEZ80ncGVlh9gTqMBTA0CEOFn+9pkhZxcnzvze84lkShvEUKnpUdWgEL92PIff
XzcCzJgb1qCxEOuqzEk5rWyoyZSbMoLjGqkTdKWAENmnB6eW/FAfz3TreFaNVh2/
OTmOVlvfMAn4D8/dbPfUutB1xyoXBB5GoQhjHgzutbqXjkCCQcWBI3eVjG9dkYQj
B2t/dl2XaaMatuUUuzR0U7iaeTS+x0HCEQjUF882eH/6hQbxpXjK0AFIIabaaHOq
ee79USpVY8AILigOlf+OCz0Os3xG+Mgvsy6t48YDD4xBIruZStwIaogyB//o5uKU
kMCUPKvu+0dtI+Js397J4BGIweXvda0AFv4UYvQ+2LPNCm7/XSBEXcCjuAOLlqRp
1pWkmEQKHit4qhPADDrXiPDYj6+mlnaG+ydYHUHW/9lFs2HjuQBBZli3KmUgg10k
NYXBEUEB1nSUCp593A24UwbsoIrkVpLvdA5o3c2ekCgU6HIhkIzVaBGbzQ9LRh3F
BnYFghY0vCMZqFPr8Vo5+GA9IylM2p3S7bRKizSA/ghaw0dgvOt7x3UQzuTtWqCz
B8vFDbfZ8JnIRhEezll6W4p5l+d970wBSP4r9pOs5bNmok5ArW8wsGmwkR06kNgj
DS7NijaHN+dEu+2/V5TsnGjHlgEYb3m1zxF9RGCheD6rdN3+OxjVkf8z6+z7aQWw
URLBFmap28tSw8xtk2QhASKMXx7oa6/0ai5qKtJpwy3FgsmhoYbYcRIETzJ9IKrL
JZcZLLwtL4ieF+5op1+ahdIK7f5kfpDSHmPYVSN+wuWnTPEZspQ4+OPQqXivvMjG
R6JeCcZfoX/txUcZzF9OTsjyF+fb2H+VhlQS/R9klHh4Fpcv8h6fYYgLeC9N/t96
Se/FgmwJIwQVjDHpT2tU2Ou2KVwiOORh3OVj+lDGzNP3UiK8fYy7UNlJDjJUtECS
0Zu17HzFxgZBjUGZOiug3ciAknEHgurQFsDhf8tsDkVX+zc+cY8Bv7FWqj2xGVWr
fvMpvdcyg82/VCGYfDeWSbAYnJszI2OiuLGDmL+Yp1NBnNcwuezEXUikIK8hXsHo
NNSTSJiKphvKgSO3NQbKRyo/jjklPfBq+3GohRtrkJ1mOtAc5D5JF241IqLL/vCm
0SSJcWUV5ar7FKqFCBavGzFIaRd97sKVYnVRoO29VEWcG6LtlgFiPnNPxc8xgvnO
92vXOJ9u+9yVrWJiWhdKP2mHccmGMh+XtrC8sPUhPcriM55PJk1TphB+eVN+FcuU
7FSPd5kbzSyK/wbwFhJexH65sqfWCfHyRROXZ2LYIVl2CnRVStGXcydei46pAd54
aHI1PwHLYhHo7ibXqKCieAAZMHuTJjhD/7k9ROZyoIKCkXZrrJgOlVrj8V0DO429
mLU5TsQ/B13G6G7ZhbjjJozd8T7+8V1qyUpAYLtoZbbL4valUMRG5bn7YEW+Fp+w
lxJOFq7K9nF7ta0hKpdTNG2Z0rPeCGMdtdwD9ZJoWBmcvqyFAL1ZUKtWfhcz8J9+
Q8yKxrCtuIZYD1WnZq92hyFedOwxUbQtRdW06UmtFmFsehf1DIqQuvdclsOPXAti
2GU3Hi3Tru67l9VrFzuUoIe9Dnx8iuqmudzPDdRY2qvrEpBhP3xx+Gk6BkjiU8pm
qYFa2CuMb+9nTPJpCJNiz+G/KWIRTtqlK7r2kWYMKYh89vM/VBt+QvPNk6klhg3r
u5sKdWSap+Nfj/fPWdxStjURORKKR3tRzz2qpsnngUiIq5rOfUJFL20TF9mkO0y1
aERAY7TS/1+tOOC5cdoiP6uSYTr/0TR4bCnPTAU6JsEpj2GXuhxdkXroBcO+1Tn1
5eUB9GFo0NqGGVJ0f00ITX9yp46peN1NS5yqeyr2sgWqdw1tZTW3ssShg4PYtn0K
MVpN2URzrE9bmW0XZxZ7LEKVeIpkAhPJ77PEyuVn7jIgbHPV+gL/tspTTjyRKML6
DEoz4mbmzrVVXOTOV8S3/RxUKBZDHdmw+0O9IuAnS9l7gSaTZ30XdRblC3T7gdw0
XDnTncBt2WA+1y6Oe2kI4hwDMjlPAUJdW1IgKayV999yndN76p5IAkQEHs2nYSGF
g6AItzPRkN62QLJt0EMJ532GM38QPXrFIv05akZUt8NnDTKaO+po3/jjZUqFlUWl
/p3qqtT/eGXSbHQO86GFNzZduZleCEjECr+8R8KrTdhZHO8gkRy5h1coYEOSwOyI
9EHnnraXrS50miHeeyBN67QYOjTX/IA7WHoOVvkHC+F3XwUwq4HUC5GeBvj1KqK3
hQkKLvkhXHoUfE1ZZbzJDy8brTMP+WinG5odKJq5nbWDX9lEMZB7UfqBak6wrwR1
F8uLdisYNwsmWIno6PMljKCR4HFu/FfURArWeyn/w41f3Z8xwTuDcIj28O+nXK+/
BXmTa91EG9mX7CSihAebVZCkSFOWAfNfIAebe4lMxsDeu751lrAVYJ6fuTniRfM+
j8RC7NRRRTzI1J+74o9ilcis9mQZ7PLuq7fv/b+q+PN9TZIFvtMFtrRJp36K494O
lJQ4GN4eYb25zwteadBY1w==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jYpzIJ0PP0sZrG+Dxt3WdE/1OiKsbs4G6hQyAwMdYRsEA9i5U7zQn0a6KlkU6VPd
k3RmetDtIm2rybKts06/ZaRWOAidMamb9aW3ziGgwDwmWQ98kewPTA/a8B9mpMg1
5VpbO9iHc+WZj4A/BmwpfZ2d7cFTaRseNMbw0ZvahkKwhxvFrikbcLxvEEUhw2TQ
ytJ+bUt83Tii5aeMVPKmThowMALLBkmHbfts4/p33qyk2nWR4C7EbpwvLa4kNtqM
w1rOppovU2UXHHMrHIrbHdQ55KqmqUIfIbT+eon44/fHwg6Bl+io9fxAr2/CaX7E
cOZYydg2d50FyDXXMgY3PA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8048 )
`pragma protect data_block
tjhJyP6EvtwlUFMq7fA2OTM7m0U6a3zoq/S8GCzE40aKYhCeb782hWkxIG9eINAW
rTH9gYL214QOkQ7wkziVMv2YR0ozsVaNMUJhqrj6wtJbHLW146NSL37dq880INO/
cb+zg6r4EV3xQtlYraK8/Zarp642fZqisiFU4+xLC36EsVlwyfftADGW/oAkiWGU
swrbgcawpyQRyiFdve3mtZu289c2qKYdWSr7RNjiFIgQABEjVZr5wZP3GeyZ3jql
jNEhE25EwwEIJxwApyrwrt8HEbDoXPbCDWRbSrSBPhu2L6IM9TT7LbHS/r2pjo/J
nhWz7HIjqA8NB5Ewx2nLrJUViBClw10n/dSpURm1u4BBBBjRVfW8fi8sap86OMb0
v2Ntnrjb+B3LyHQmuB0hvVmKQCXYwg/aSsElAGASwQAvkpOBfQ537cW67j6zsEm4
0VX3nAccKOv6X4y+2wVy1uobJ3GIg2nmEEifLFhTi/KeJ+YvToHp6jxaknIKqkG2
jz1EJ1KraZkAcOgWqOybkoEfWUlK6b3YDuab5WOlKL2umqF+LpVh4Utu8ZJ7u4pJ
uKJX3xhxuEjMdZFQ+M2+Exj74vDVzaBj0hIPBJqp5bYLwvawESN0xA5G3T1oJpuW
SODH5auGMl3GxhNdDKYMKGyjD2NhPiNUUMt8GDAFQtzc0C0K0HND6UKQ+Mb1xKwP
bf33hDJRMJ1Iotn3OJucmd8Lij9NnqIyB3iO19gqCN1u771MbdtxMlalQuSwtCqt
i818T6eXvFjkFbo9Xkt/Z2OsBwfNN01zNoPGbZ6Xg5lkNgxIdIIGg9YVRLb4HM0g
LXt9+REBKL8xyMpaoWPcIh3uR6rHpyKshFJPGjMhROWfkg4Z8S3tHVqt0FQ0ah1E
oRhqUg9SfSdwarzJ2zUdT151EA1Ib42jC9u0vtFSEnlpWYFpOsm7ZYC8vdvuGyBc
9ZUeHlFZHjymVwrOZKtr4qiqPzZ9w0qyVCZOR8QmIE5WFplZXIqDLqRP8ign7zkc
60HVZi8ynmtHpZ+VfoCJoD5NkszoXPwydVoXEx+5gaoEAWyZoBvqVLy63XGI5M4H
tNZEXj1xIUYVD15drZRtxBnPaC3XIiqYdaj+31RH/oHDJJXHNfeE5Ar8jKCZr3HF
HFPVQqYRvzXvomjmcbd/fLQtPzNq9+7aYufZ4Oy3TbcdR5cLrt5SmbK5mh1alrQl
zKTZ1D+Q1VkTYWyzHiR9K6bjVWhouAixRlIOm+jJ4f+bnG91ppIDZ6MHq22bdgNy
scFxvgnmy0PjTe4pMvxzzJ4sMKDin9EdrFH8wHZLDVv8SkMyAryo73EUWs4oSmZj
1fJ9CqsseAvVYh8SoLWrTVVn5TlABgzNy6/0IRprADAl8meovGT/vlboK18UgpiH
TtC29yD0epQpuL9TZVUhMwUwpa2wbEfEfrKyMwlftDxXZZSmKHSbPw06gKyHeMJw
t3tAb7a1RpPm2j8Rd8Syhx013Cl7vvewPv3mlwEzcuJTK8OzWnyLoi7Q5LrM8pTu
HxlVxr7yDBORjTSWPDHtzozgxhcuVMtiqm2o2MMcFAgS2TdCY1EU7qdKV2APAPAU
CMsH/qzMykfKw1L94pLDJ+c2D8QBK0q1Zc4zQp1IVUo704LMi76zfo184VE5Omb2
Oek2LGbQawMkt5sSRHoCCkI7bdHC3Iv8D7UzfG50aQi60rfyZX31tQvXCI06dbnJ
8AQAUf8ZAx3G/Q4fvyFO1Cpn24Gaz6y1BKZE6D7uo33VGsdt/UQpo01nzFX1ggz+
Z9L7Mz5CpkVLkQigqYlmpvq0NkYubkW/vKuir6gmKw1HWA6tSM3Yj1xXMGSL+7Gf
G3SdJO6Fv7hYD4KhLdgp+OLZaAsxRZQ/n0JeKdS4S+xGaz7Pz5vm4spSnYuOklPU
KH7hJv+GpZrMJj+P2BeDlLnFzO5eGRs4SLQVhGLzmFERRIN3qzST/JLsv4O/H6ZH
sqlM4zMaiN/0uSL/O8xiFDt8D/4OwQYRy8ieU91XWW8Rm2Rv+xz21hhA4Bm9dvvC
swspy2v6oe+2+uPnoN0G0OstbnIE6HcErTg9h+NnD+C1Z+2U3WMC8Jy22zkHV3R/
cy3u462+WVUpV5Iq0WnVKEtcLWy43GfMI6di3AEL/ASfRUOWt6fXvvfMDqkYh957
tGSkp9W9hcMl1YWaxUapm/sCqddtJ7eRa8f0zfDVMsJXyTSqHNRQb7NEyWF7gpYk
+7P11j+gIRaBmNisuumJ6AF2fyZG6U4hzKcXpJsE+1POJVS8PoDZUN47XmwOm9nu
YcUrt8DKIfjZWXl81ERxmyMxR69ZR30H6+7SowGMm3xoxt+j09umK8/hR1gKQUn5
H0Rr95p92RE5fibjcPHyDfOESKyEC8SfuzAOSJ2axLnL+ZJm/uw6tsqHUDKuGOBq
CH6wOc/UtfCAD73P5CGSlQ0r8r/Xl9GdFoKiF7RrhIfZI0dasuOAaqxYepxFbAkz
JRvPxm2UiF38k82ckbJwsJ2dyb7stDoXLsHx+wMbf9JrFIu6l4UOtEKVaNTHnEDS
qstecqqe9+MXvZ7kuiMruQnXAe9YktKJsNgFfSIR43iHKT7VuVE+ZJQ48SHJ2cFt
u8uDu/cc8vod1JoB1ujbp+fZ4SIN85mMEiuEr7pMAp2XqQ+tOmu3yba0BL9cNZwZ
xW7PXlDuOAh4khp29V5RyD9kGpmvBLj4PHIFf/4/dTdMBD+WumcsblJrKWeQ48Lv
eZnyZ7SAFB2UzeAOPn6tXGWV7GGb1yswlXFZqTjUeajYniRaelOnxIlZ43wdDiDT
SkvAGF9s7u/j+v7TRtengIbd/3d2pL1fA+5W1q3V/Hct8vljgBIAaHhUXKAy6Fnn
WK3ie26CbCn2YotKJgslsQPnUPPr+AfMbFHBTG0SoWPLOdhRqEoqdFGuAh9IVHRX
YtNakZAKMOP3DQCTyAlD5JQklqdOq4jMsuny3oNHI9g3O32v7zzr3cmvZtGqnsB2
ilzccT6ezZtdPiEurZiAwjhgiIyA/dolACYhDZhxtoGw3D03Qx+cCaavI5iO0lSQ
gwyzkyJ4Xs2K0lD4ggcE1UYFX8silLfhuvgopP/RrAb6o9lRWuNPdJlGPnlaqiOF
aiElv2az5KJ+jk3PSqEgN5nCwhJ2o3tKTvfUTejTMEEFpAPyFcU2sGke5XfhvdfH
KJ4xLY3Am/lGy8Fa3Jxx1lXraws+F9CVZepjFq1JeHWDPpCmdmYwFGD8KhBesz9q
m8lEnqSl8duDhU0PGg/BrIgBwulOrE7KHqrqSAig+SwiVE/UGkOxePl13NxnwnpO
9Ev1Z1g0MNEcluwjmmWCTfKbySYEMNP3Mo0M1NqZFOpCQvb+mebqQoSc6iWWjG5W
Y0MGS3uGhhAqH9QZ7giR4IRqkNVVMrSsVHHgMwW0HFGB4Bz+JU9Pz/qmO13FqJFC
zb/WVfM/sUof0fPRF9Mq96zxStR9Tu0aKZuyb9Ro36vMYFPsGV0hukqGX+eXcOUM
mdikQ67taXLDOHX6FOEFI8vAJneOS7Q8y2oLRGnPIlcjhLi+EEqem86bKqqhL8uk
EU4x+JZGG/wEI2c2q9m1mOuGuRPebOAqyaa80Aop9Gm7563XhsgKg+2eCkhbt+oP
QqfScvaykzLVOuzS5YmamZHQVn+zYjEba5NCGX89H3esducrmVo1ihXZUOG7QX8a
SVIPZ00TbbPWuDFXjeN5hnGYDznbb3jx2SMqLNfSQ/XJx6Z9zeFI9eOvzJBaTPXg
NpucCZqrXpjK562OHkTsmVVFiyxqqDOa1Ao0CGHIFvnrRhKt5zashInt9pLQGmOl
my1Ltij/O9q96/zVblyR4bsfsnaDD54W5anXgGDA7IyIGbvAsqlTUiWhHE1XLg1V
G/+96mjnU8WeXGPeTFBp9JH4N7tKXiwfvw/vSfgMZCLdQP7nwdeQYXxt9cx3Ly7W
zANE7B6bOV8+JozFO5894j7K3PGAq6W9BBtQTD4GdPzdxFSK66cGL71JxT5iEUUp
HUqWocHzAGv4N8VPo89rB7aA41bCIAo6JCH/dDs0kdwZ1WVo8Qnyp7+I0OCbQRA1
8NXbbEZVxiD1kUz0AsxxRtSi61VX5M9NMn26C8NcaYw239aIq/jZwSiQtcqoWPHx
N51nkt5byljxsc9ww3OZ+zrdrIERIxKylncc7gvka7DXM3FhqpuCumnpV0//886G
m1KiAf/ERfnSa23ZVUc9VLQol+n/859oFbA7rsJsaN1eDu/UP1KuzHglFU/o7kxB
3Mnmg2Lv3QFBAeJtCuJv6rhwqbnlpCnorf368T36eO+O7+BXT9pitzzW32dcC/fw
EMwB398sFl9kHLt6gVniETujJFQ+rLALLT4AR+0Cgp8+lJLzbDrWhC828DH8l5RB
3W4bzyydPYOvvg1R8/owU7iNsgdyAYbxIO0U9EI796AfcvtCAHDp4wwF2uyzPNxG
4HmbcF84PAhItTOwqmhg/sAPxHChZH+idoZRusj6gdpJWFrOgGeHiGB6Cjj/xkZO
ey4OkdRhuEDx8L2x59JAq2SRRjINbx6Nh69JNTol/VZXzsXtY9al1KQNnWD/xUF7
KN2sNZjuiKEDOOOxP0JV+gYhcqTgH4XUDkgm+Pvdezivjc2iE8jH0b0QKmFd+5IF
w68pgaww6GIuVj95xXmmvqdMqz0agad+06zxTDqm710Zqhu+J44fwbWhtWustu2i
T6rgYpnSFTTfHhWDy3HAyKKfERjZnl+ATq1cvdnuaV1lpG/sgbWLhN5Fn0ov62de
JAjp7kvHgyfqKUrj2kHyVYob8xIobkoONY7y4J+zyTP+OFd/r1r0JiOvyHbEIYhw
/tT271IpkfbsJQFfJjvdBNyLRQl6bM2b3h3eFbi7quP92uwM7XFaasjQDF7nbGF7
Q/jZycIgPyCSeXI+Ys0rn1fA0xr2ykbmsD4QXwKwIVcjwd7gy4zNlKl/ukSnzrOl
MAVAen+yFMKf/JVOLdlPHtPl+VKZ4nW2u7Ar0gDyckGZl1td13+CaBGFOPQTLif3
qx/z3QmCwIwNcIyDUvqphOQIDI+n3xlN0nz8wwoH2ePSp3uqntcyvWlLtDt2VWFd
a2Gf67zOscKGCONBO4nSpVpiLkwGRURscWhNw1LdKiV6vJ7FbGozHHyi2tYoKf7a
5bmwZuROaUcumpcbh+grA8P5qecENB+wXgMVlt9m5rTVT/AX2JKEn/gUu+V0RJRi
paR673W2WLIXdgz27Lmt2gg4Tqpww/CB5cwY7kwd23mK/XezY0/P+LEEVOVdSKrc
llhLF/YC2Eo22sS3/aLJLkzoZuz4+BV2ikNNn0HjRKk17NCII9krFz4qAIUsWmMW
LQx/Wkgvnc6oVocWJWzJPMyFMgPrR3xaUrJ5CBLXrWnXxzzGH2FhvNYF3qOOYSor
JOccY/Zb9w3ljczReO6XVrZvzErYfeJxwWZLE+u0Tw4VP/npINoLIuxPQwnaKGLe
BVmk+au3+gNMEPVeaScvWw5pe6PIP61fDIHuLDB9X7BKJWmWaEbU6IsuSMxycytT
t/b/n7u+qOTkYfPKAonmHP+nWXDW73ej5oHgJjWpHGuiq6HGsN0G+MZPoAbWEtJ3
QANX8DU78LP3jTyhgN9supTWAqgcbzFNjRYlVy6D6e/05NWtaeGfRs9HqN1YavH2
g7Hdj+tvxvPI6CgcEtzzc5sxLzA8v8bZrax7cQWdApdB3IwL/ioXg7m87Bfd4ErK
dn08cKk0zAitTioRfqqDhXa2NJOitgn+FwdGlHm8OiCJ10W3Me2i3m1KbHxfXP11
dgulwS3ygXrqaqw4EN4OeS/LDyOWnsQ3Kz7miu3d5C9xmDI+UJf8OEQQPuHsbAk4
iHDOgLoDyqL1d+mtOoZ0b1WVqvUr8Ptpc+TSDhhhGOYdCSG3dY8bxpF+QHP9yIxO
vER2lDnym4GOSRUthxy6DPoIlXyj7/bEwmiVC+6YcMU7EjbC6+V78E6/0jESPMdr
C3pN1dJ8iU6lQnbfLP4VA8si3060pZSUqRbCqPSYTOgldkdyUd2xsTjtX1NmWVgB
/gw5FcL/81WDJMYoCVCVRio5P3VmIiohCZ/m1OmoMvSiQZEy66hZlQNikv79p0lL
oT8hb+UWvrK0PzDs9Mf1nhyo3biiw5WEBUK4tegXjtYeTdq+/Vdk2ItGzEl8IbIg
50shzBUmZzM9bMr6z+GmAnHMBaqImFfniiddC1zNXLvKycHn32rjhlW/tRVWnR7F
3NAbVut8RhHOosG+4OF3oIC+TZ9Xb0A9jvP80rlGctAn6tH13ajmeYsqCpDpCVqj
PCKb7Ot5MGQRgYzFI/HYcPg4MS1oJfhR/xO34wnzwsEYRlxuPC9G+IFtn3Xo12hm
DqTxCeugYzL9PQfFwIw6ytq1zfoLgrJNSowUqYYA4z74n55XXHzWHZIaXsoow/n2
6OcCa8h8blZpQopFPFGD/eD+GSE0dtDCx5VMRho0QBRpycgt+MBu1EQ3e2QpH0ej
fQh5CQf7atTd/datGrKm+j3tcH3k0crWj5nvRWYUgRQ1VsAyEUMajBxWVxcoSUGW
g5+QNBanKKk1pmQcmLL/ey12ykNczEqK/mYXLED+UKzdokUyqHzojN9dvRdVuqUf
iSaHugvQwZ4xJ9NkzWrvY0mswkcbdQY82hSLThB5f+Sso3/44gFUzHfEOtnSS0Od
D/NWJiO5KdLBhVEDiuPbFevfndwRiW1EN0q3qT0t0Vodd5u1Dqsc0I8kbPA87ZRV
OwRAtYHFuZUgQg3zbzCKajRU/DbYgi0XeMfiUcyN3J8mrQWqx3ZLveN+alzECfvl
v33cLVIq2u7bfSskOfnRiWsTGFkF8sgdI2VHO1yj5fwcWgesVg0IbUKNIX+2kgaS
GsgIaaKMxAKiNZ2fPgfI0gMXV1YxmtEYFp4pytfBJfwE93f9RpIharMKul48MKKP
KJWB/Tp3SavwvbSlRnTO1wswLdrz7Czvm9FeKMhLVLg2LxEMCSr9ufL8023d38iA
QLq72dQzjjdUvWKRhmXYnOaOnQ4DIV+HxjIcCbFZGZ7nkhW7k2TzLkfb8uukOp8v
USnmvEP5Ni0JBIMXcY4wor94jgdghupE0MbHY03IoWPj5N96VxpuKCbjwmGoAAB2
OjcQ12WOdXSB6uxT2VNcCLVXbANYhuAVG6SbQbX2Bux5Ma4iOxCbgoDqeaIrWk8i
ueBpps8hUP80+g+DQAEfmEQCCT9JrrRevsBBnmP+HlojowUnQP6CJ4y8g1PBdKO/
IexyGDNcfnx4gsrLrfjmCQS33fYYoHU62X+sDntke0aWV3/VKaqC5ak/aU5FNueT
YObwaV5FiKQv27X1bu40Ho91O/HgeRKU3oZfv+8DshuIufBOxI6YLUi1zR98SWRw
VokwCUU7zdKrXKds6c66lS7l6d6aO/0HMWWw+hnt1nuWHTcJ794jnsob+2GLU9qE
Bd6ZbkmICgEGVwG1tr5GrwJDRNEyzbEYegK/y+OxukzNnAZzwsXbec5cZfQpVoDd
5+Kgd2GQEC6skw+GOE6Xa4AvtvN3dQaxRSw84e0QP6Cek+2LPxZZZq/v1TKZsAQ6
NjuZvl1l+oxdE1hI5EU/rihICgo3WIByIJzf2JJbKfgWlws+aEQa+Fb1yQvkifd5
cyF9DECD2Hd+nVxq1ZK/zrv+zGp8qu88lU2R9fOfYVzCavyq6q/4A7B0n64+LuFd
5SOCEOds15U4JqgoCE+Xron2mB6CXEFwyf+a8WNFczN7FSJjxGFoAIZQGtG0JUb+
wwYMdk+8dWRN2goTsGfp/ibjyRI0dawP6LiAIO9yx3tdvjvOE1dTE/Kiym2VaNBG
C2ho3VLoV+UeZvOZg4sFZw+wMZDXu5lgIwKhShpHh3nhuZb5dRHUTIIPDo9F8wIg
DdtBrsVMmvU/JKX4rvUnrSkyqWFSALmBAEIEfhmdsHQOo47RiUGiOizdm1/z0pZ0
xluUxLzFk1waX/V45kVv0OprPs+UgMX87Fu2R6W2yQywNmQkw8yBVZc66xFCEn+d
vkQKDSkR48yYLPgC8v/JwX7VotKwhjurmTX4axzDFRwSDi7Ah/IgxBlK3Y2lsb2o
OdVm5ho3h/k9dt1YFfWy2R8z77pg29V18l/63XrZEMGxjffMs4prjdXO9VKZI9OP
LXr4zjjWAGTEtBsFT1rIjtRum8pUsIWa0kekX2Wnh+R1i2TbwPh7KnCLZPe19KVw
//6jE7Ej0DJitDdLewL9NLABKgp1sVGX9RfkW5szn/VZcUQQtnZXeszN5SgGZcEz
5wBMyd3yBr+D/5jp3prBnV7/1iiwPPSzJvRwuF6Vvmb+/SP39HWanKWhgDeOeGYE
OrZ6wO9CwpYeOi/LqUty+sYPF+b/lq34+u82Hz1PvOo/pMBq1HYwMYyivh4kp0Rc
kVyYRrTbzJ7o4b+9jbQ4ucwdpkEPp7GRhESrr976SQ9PtGaEjuW62hW8okMAtUZ8
aZh25SsnyYHQE+1lZTcHVAkSGg7rdnA3IT56r96jlB6X6sAJBdXjTHaEMuBL7p1h
PUyqhgN490QSw+fp06Q12voSvoBsfoJ58dbL5ApKNxwPr0qICVxhjOe2uengZ88T
j5X21LEIukClknRkwjhSZ7pEWfkmuQb8sIhH8qj5ZWlLa6RihO31HOHGkW5Q5fQU
XgLaZEZbmJxjRz2nvP6f83lexGaibAX4zk+RH3gsGfIodWZbFKUsT4YHX/9LGMMT
N3A65bARSSrp8O1LTVqodzLAyRYQINz7Vqwxir/lyf1MQR2oHvSTuZQe/5XIY2nn
g7pI7HfI4Lbb23KSUH1dm+9VC7e85557nuGai4MXB15gpXDK1s5q8oZgk8zTXCIq
LOyrv26vvqx5QeaPRWOxnE3JuZGwQFLd4caWYTCpf4Czp4pLLoBRnSdFGk1NCFyA
0HCKUr8NR/nv4eoLtDmx+SYLxRUdXjw/WVsIrqMB7hm0N+y5AS9S0t2nIqARJD4j
5dFPJtxVs04RBFPiDC9HcvFWGLViqIfJD6aovdB+1XnVY/aO+8SMNRzQqIC/qkZ4
jj/JY+eiOcjoCR3RLg1EC1PRQY/jCLWmkWKYe8NzbhpxiKGeAAg6W6v4qQ5COFWG
W1REB1o//bHyMedclE2WGycBJI5s3TW4+3gkz9sCJsQkK89TvmS+A+X61UrnebFJ
xVyc+M8qaPf7veUiWnIUXyQrkhrm6s0/ikNbb+zQt4/PWx0zfx7EkZKhlQoE3B3J
W5WxSd5qrWi6j0Y7zm16dsjknn2fz59PGdhZ5lEuxcuuL2GvndNr6y4RBBbkwJKv
HCIZnEtOsCpKcm4j/D5GhlEsHF3k9D+FLvxRNDmsp7U7nXUu3PrJwNLXjQZdD93Y
CgrzbZJNVVTcUD175cHfcXbJlxMePpbZafD/LKxMyzYV9jZI/SDqbDVydHq3I/CQ
EoNsjFVkZ7p3DqSqrhfzphWkK8Z7Mjba7iktRsnEe5GG4vJ1eUoYzAMXZe3XEDou
hIk5746vCC5yGPGj2sQe8oC2mgCkpGHyffao3ig88QoEj/IlCT2x+3F2SNtPdSaM
f2+68/BEkCMu7lmrk6PG2xQTcVbcgeoUCQVnkTAJ4f2WiLXLUUq1V0mq/VLxJ10D
0LKFcZOihayMqrBn7GQK6rmLiVALJ6FoT5JNFEdXiahWtLK1XCmwEtrHdKrh1u0n
gTDzVtCANjT+/akzYrrE1P1r8USjPFjPAc9vZ8SN6lOSgmWWYzHmz8XCJgdEDDsi
8kVwb3GQ+pAa0EbspDRo8wPC7u2QCf+Rqz5oYrlPCayvp/dtLBm5t/MvxU3AIIRB
POJth6n7OBI11SsJpWtdz3+3Y8XJB+h984zCM5MW3uWRDov24eXnYJxL6VXdXjpy
tXhWdhgS6bPnx6VKWSHJRXNAPinPS3WqfAcvmmL+5jCe7OAbs1TAShqnvpbfPDFG
JUdsvqdZdO6Zr0p65ax1yhbphBMc7FZFL0TjobJ5uDyGCNX7f//EmzfBfpCUJukh
5owYrgANUffl0ne+JJm9fY0dECKmZ7YiuedSBLGUGS+ENGGqWVCr5WM1UopMEKH6
OL51vlpIl7Nv+t65hPpm2Jdgn9nZvMKhcYJY5w1C0hT+tm6mSiqarMD138bgw2UU
L9cCKwnyn6F2XhlYCWzdXF4CEzpJ6WoB30wuXSq/8/zB3PkqTm3L+T8bNo14eNt2
iVU/ApkjuxwusIxmNyiBuyMwGBxBceOc8jYl6VAehw3ryGkZQU1CqcQvWj1EvwLT
zReTFnzzZ0K06xMifgPm7wy2WDsDLHQwqY4r8vIWSspLkIxitd4n/xN8QcdsuEw0
WSqdE0lT5G/R7IGKjHK/gSQhWID3a+ME7+uem5QULCWvx9PASRfH9U4qqYIwx+cs
6vOsi1zEbtnF5LKqIbUxIcGrbhzclUhVkfhWfg2vR08Qe4ba7oSHDKgSfsf6HnpF
4Y5E3JH/rwPYvfWiWa3Z0o7ZAHYKSABvph/FhZvqydC+VKupB2a0hYRkEpjAAQsU
79pTCU7G5CrC3KTEabc2JblKzMGFoqgJDjtX5FhICpSA/xrPee8FcCK72pQNAiUz
qYQY98yuOT1ezpR5Gvd3IKBfoWcstscNfoC6r8t8DNJJEX3oxtOEW/Dzpvge+K2K
MfU91ApszXOUDk9TuVUnJFuHGTAWY1FePXi4VI0xsTE=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jauF3ebLgD1sOXuXiwYuXpR3qVxQ/Pc+zw8Ms0LGHQtaqvicZA/+vjXsoEZ05Yal
xBJzf9gJ6abyUE66LIQuIQiWVS3jhoCkF9NFOnZ96qQKKQ7RnvHPJAxaOkjujpGG
5wem3CMv3GIqVU4sYxR/bi/kNlVjmg4YWlnuVd13wLTaIVvr4G0qcQz6HlOT0KPo
OZFDWzdmmOJPuP7AD5uxlBSiiOEIYogaUL6Iuo9F07KNQEOGzn3w8QVLll4sVG39
MdcxUqOs1/ZJVQw1+N3d7j9NauU0JnbheafvO9t9xX3F0OdzxSYay4OpfFEqu6Od
9Y4+yWBkChpOINSrRFFGjg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5360 )
`pragma protect data_block
B2Z5+P5DtTb6Pm+2Ei9uQ15Xld2RXyvF69vIsdXuVwQl69h3kFiuyHDKcb4jqP4d
CNXoxgdCZ0fNTPpMm9hR0EsFaUrAWWjH2zZYQng56uJn/fcixURaLLOPW/NyHXQr
8a/cylNk1YO8YjnkpBiOJnKtYZgPaPhGOtCIJ3AQkGzsPBSfubtcbRlJJEIFMtJK
xjAMeKBFNTGY78Q+dFPzh7+3GiCJ0rP/ybBS/8UJBIlSo2dOgbuu70xnIGOE9yGp
LoO9cZWnvgudsOhn5hxvId+UROuH3B94xQ5nqhQ/kQp1dJybqGRTNk3hsUjDQ2C3
rVxCqCZNVRI9idQOo25Crt0CMMNUSqdyudCRbGXMlHtaQm3DMKwSMuBZ+CrDwHND
/9H2o1ENC5Kw5J0pIilz9WtZAo6SAMcSuv8p+DI1gJv1FeJdyaLon+MvdX802Jpy
sfp4H6zXKaXqa7rHkggiD79l8/58+5Bz3wOqrZ0l0NeRvwGZyK/gqNQUL8sHqLbu
ZRdgO7XGzSYseQsvS/+DKyah8VWFIQEOAu+g1+eUkPjjdCbtTAn91UDVjT/hpn1r
0Sky5tWY9MwnUSoR/51m+EEKOlk1oqkfVbMJwfsvO2Wsh7M1AetnrLgeNvAQ9vVE
aKhiUBWJanlJfAsSYcTROMKRK1kG2q1sjfHk4nt+P4klZwsJMMIdv7KEGfvmVsft
d6jXXSlDRY3Fojv/C9xAislIpLlsE7uhLiDTZVx9FTf+Qm6Fie906W+zdDfKwjiZ
coCmvzFfkheCsNQJ/Jcr/r4/MwJUCY5lwO6Z8nSceSAgx+gKJGK78I/TdMqZiKe1
R/GNABKQ5/HKJrIEnor1As55uqeCTPhiL8600aHSuAHdl/PToT5la6tdAYK9NRPQ
aB/IzSCM5Rohgj7y1R+CYGQ4dGw2EzckinWOJATKW/QwsehASvugXFdxoQC0Wr2D
//EJPNNiqzyvfKZR0DFy+1Djgwgo2E3tkAo3at3bTCMHrQvaa26MvDjYdlLxfuk7
2P5+MWTEWkuir+r9VCckhH6ec2b38Ah2VZwJSfj/8x2wGX61KcAbR+WXfhxuDaKG
l3sQVq4AZhT82HkAjLkwFOteDOh4FxajGtlpdFcYuz2Od12GjO/FuT7v2KTzZGnz
ZURgLoFAXkfUrwKi+2IHc+2AUuTX2BH+OCi61ZsLYA8azqAW4Qd9UmIYTKXd1vAH
uMuvF3qutf2Kx5YTpew1vNthGs2rOlYPctkornmXUO9uMv+XZUIdU+T9TujeRf6R
2iSLHgWUeq/1sT595sO0FbsVhQOsYxvK2l6t5oevL/90un5ikW0IBnN1oeM3Zs84
FYcCmwf+0AcoQRHUFHnmwGOT9Y8pthSbCQGh9r3yqP15r6qcLyjtkp3oBnbYZWiI
AbnTRBl0qS52S6JvhQnG1RfyW9+qKlBBOZRme9mNQenuLvIZNp7x/M1HqiBZrFix
K2SX8B6pKsh8xlxcvz2dB0c5Zx/IZCdyZJnHtwAdN7HmolfBa9/PL9Wbpu6kZ5ku
ZRfdz8uFv87ajtSfOsHZTZ6Kf++RWe212Gqbc+wlOnPUwx7UVvgCFeNrNwI66tzR
5kg0u6K7+VXH5fLjpvWEe11U1ZJf/efr7I8O5dgkWjRpPaUXPvxzrdLwhwNCTnCB
rLcq031kXtCQXhB6aWf8ElYsUP2j/IMbqvlM7WY7L8pAPvBGo70WFK3PK3R1mnBG
YVQ4OVL+PUanTKORJ10Ut//7AhMNMMKNHuxQPUB3kcOLaKk9sS6kLMHJjokS7L0Y
TnN7KKa8HkZ1LLQJvVW5CZp15Bud3XBUo7qt1a3OiYUxOAFpOJ3H3HVNQuJdyIfI
MOZ79srJJYd8vvXrhQzEW8R1GksUnTbeWmbcJYTABnzFSz9EEJHenfyLdxaGMyR3
SjkwakwlX7ShAM6s8X/aZVygv+yApvWYyhfHaDnFE6GfBdFuNTMV1Y91CgTqz94Y
X4YE1tsak/6slle3GFETiaXIwXo+iyPBo6/UFlQxePE4F24Wjf1rRyrXxXbsCdIk
ytEVn1qPjZLzLCq/6gRoi3LDOw01byt8Jji2/0K8isTM9BGAxqiQmmAIwPNh2aLo
OzdUZtjEj0c49/TeIvn9AoF5k/Q2uUE0XmySmP9bUYioYIHNxEYZSk3ixvHpQFI/
9bPVGc2F++ELlh9vrtVMUyyJl62mAwOeR9b702nvbCdZPoAcHltrHg4zI+PuoK2m
GbFBhn26pjH7IToRkxsj8iO2rEik/Z6ZawL2ee/MBQzDGyU2G6A3b7Re8J6+lhiR
+wV3WuuhnkXuP635EtJBksXPkuN40yemucgdRqjkbxlAihVQOtj8/vYFxbi0wGk0
q3vjHsipXwSl+7SN5UXTrUh6mLm5C3yjCy3682qU5H6+wvcjy2rW0bMwAbi3egXK
++RcuWP1i33RD9/NgFQeFxN5VP4LMRBJ0cdPV/XSxLpCIIkGGspxoexzx5bSqYSY
puYDSmYpojyYxcRzLjUHznXkAmGVc5Te8m+OacvsJOA3ec4B7dH5cD1/KYGx1WoY
n038GrvEzN/RfyK3FwRoNCHxuzMySQ55B98ZATKdnf0Mu7QRzNC2FLQcu4DAcpAr
HdJQ1kEwEBZkPONV/qNq4kI4bTPYxY22Yn8eKKUuKBwQjlRN/HhPGDfzUdUeMxjO
tJzMRukQqMSTetTo2QX07kwmnvqFa7ym5cfIGLfntLkYZ5OmHHpJS2jUTDNMKQal
933gdlZk50/nXBuPODBgUPDhpD6QHR3fnagV7tbDsPtmpHJjIScDtnMF1vJtTE5P
OHTTnN3rtmZIGCsTjd72O+XOM914HwXM/Tzbz6PQGmT+MMaSv1NxZBqe78gc8P2v
AXmM1nZAuDkQ2Lk7OoXKD4DWBXnfSrDS2vL7H95EtjaX/6+gn3UF4etncD0VbGF6
A0zETA/pm4mF21jLaxGbMOgBnJ4yY8Afj9z4ObDPf82r3THhDvhVtocqipBEtciy
MdsuSk8GZAvqWWfEVFL3X+Tt+igB3idJFijdYcxoDTJDXX50qUHRoSxZqvfHlBFN
iEsc2rcAtWSpmETMwpYAddBeEaN17rAScDNsKpeUeLSPIAN3q8dmzwazlFQbdeL6
yUDitqHgaJ2EtffNh7qXzJ+NJB09TwBDdEsm7Dl8Vz/GJ4Vr75ofI4KawZqgwTtY
yOPhO/eSJyDB6e6TWOPClZA+U3HYtH+A84gFc/eZNs0EMuW0bFigJdmYiy4dBwSC
DJ3nWOh3aYXaiTh13Nb0lgrQZ02hVRQamYCvop2VpFs/pM98ONEuKb8vy+DGQI7Q
sY+35x2sbRash0ZtfZKmcTDNjx/p3QeNzWv3Wf+UoDIGa30BhiKTslRB5K68SbrT
WSBzab2G/m9g/yDdEDvB4lC7uaC6xzRjgf8WjEZsTzmZVi2gZ0pIto6Vve05LGB0
GVuWMLs6GQI1Ut2K6KDvqBpXFjf59o5S/VhMgQJNlS+HGAYmFPuiL6FrppiX4Z+g
3LOQAkhB52bYd+YmruJPtyUwd88k9gBtGMZxdF1bb0+BGIl9dtryHAOSgWvNYqja
WfMnRAJqc97UgwpveLOgEJXsN6vuXuj+hkeuX7+wt8X/F2lmZjQkHi1z4y3GG6Kp
hIpwHS3sHH80vUzwSDENsSdxR0WB1dOhVKtbHlEJzKzyZzJAiVJhdyk6VwP3KU5+
XiWmkC+CT0WXSgKIgrCRJsW+oOKW5JygViZp9X1rH8i7Xs3sKy214nmmweSnyd8g
RRNfAxv7LmV9wVxBMgeEosoHpJgBE/ui9ZolgLNvtc6Ry3BcuQqS90s9+LzFDNEJ
mTNO1bEoTM7BROHV08m05N0HhFzhTFVVVlWUw36fjUsj7u/j5zDEi0LCGMOUjEFQ
hO3zpMi7XvBRp1r3c1RJ+qL0jUKQ5xhpAkMjlXtL82paod8EBb/4iVahlg5ly+Dc
bxVPv24VB2CnsaYYLUxGAvFkKubbf1ZokVbyRf1wgRVxn1AuT+msIVSc9fpXL/bo
qrr1OLA76v+Z3D/0qMgmZBtJ/q4he7zqJTTZ02VsT/W9CETwge/liU3bbUIIKobZ
JLVdGxr9QYrc6JpPjkXMyTwmql4QW/G83oLCLaJepjV4LoDgUQI78KyLQdiyLbV7
un0AmBBR2eGpxjg0vziSnZmiNe5OX5Ap8hFjByq0mAHBC/xA2xC6mMJgMcDI9uAs
vymCh33i4DGGwVc4D2T5IB2MGths17DYizOdZWPLB/hC3tbT8/vpZEYeFvPxXL+W
o4WSOJqzL/9mY11JUGVxqZBDn/kfRVXazgbt4FyszW4vNUvbp+yh197c1gO0SGfT
XHGlLSm1XbH06nlexO/wZ6P6SiRtunv70EzRibjKBycUjuKEdFin54hsm7TefRRS
eRcLxZQBKiseyGnvjkzqtjx1gpLmWUZkyHyxamrIbqDulJJrUdXZPVTZAd4Dw1A1
0io8+wMSPL+GnDg2ZYLj5Egw2dwBxGbiITVirvz8ScPneqG8t+9+LpJQzHolwUkr
7xflBQc4XYFamAd7FHX8fxKuIOaWmebu9tGeIWa85j3TQgrsc65rZi2zbSq2nSQm
hnFlqJrpGUnwcV6mbminNutfMd01pIu5OJygxffY+1VPLVdaL/MeSv1pRQojlvsy
preWrXtXopSfghGvn8o9dFMwd+zbwikVlJSyjvlMWJJp0aO1H6j5Ddtm4pcMUSAg
ONZuLiYT7IHQpkhBQ6Oxs+3hTmwgpgWk6Pc/v+Zi6hY06cKXt82grxOUL0G6kwSO
rqqXVX/WzCUagB8SJ8fEW4GkC1s/PSe+hrrbQxSiwqgwKsuaV6u3rNu4tRKUqxUo
EbmRR3nZAfi1zD/3+K16OZD93E9ArCzUPXGEVGtpiELqkZSKsIbo39kCb9UU1Kr/
owqFNmoroYSUCOO+FNwZiMa63riQlzSoWprx7cuBzSoAOMkMzzcgKyK15fwrY6jo
O9uCRYGZS2TbT1I65SRmmiD4pDggangACGxhIcdbi0jWZaTXhrfZM053apd6unPi
LTMBRXqt2KMH9TqWD2lfRCD2cdQ1HDVLn4fk7C/dykWr+dXiovs7z+IdliK1tnib
mRm5OBXMCxV/GJ1MluED+sI/sRmsUbdM7Cn+K5oQJbwzF5+m/InQ3ojNJKEM6/IO
QjQjI7apkuXokzqezBf1ZftdukB4S1l8buauw0jfQZ53QgehFa7gmaNzLvy/5gYp
koKCkwrhYDnnNN51E5KnaLzojWI7rjfFwuk5scAB5nUlTwMQlCCaj8u5Xo7mbKbV
5ckgGx5ZYDtTj9HJSJoFPDnR3wFDU5wfFlKeDgA24t9rAuA1TezpYTjCkXM5cqzo
ITOW/bwG7PdSEAdDiCsLCRug6gIx0+JPsnoon8i9Mos6AMdn1jtASWnDNOnxHZWz
+Ep9ZNlmnXlG57U4+YQQ/B2O3RLtMwExayxS6qCoveTgPWU7FDJqwqboq3m7HF+T
6OiVg3/zGrE/cM4AjN7wZB0IiLtmsKz2zulm2VmUEfpM+XJiBuhwKg1zxVn/mLMf
dDJL1sNBE/f8aOkuACrDo45tYUpwvqGdWb3iFPyw+cbjUwyYVqD21i2rRwoKiCXh
4SyveTDOr5aeCpwnCKLy1A2nON9UV/xlaqsvblq5DKnrkOp/sb9qQVCzIx1+E/Xa
aHn8oqq07IyPdnxxI9M8OsO1nB8jo17AEsL4kDdytO0KPdmK8vIe5SfiDzFsApC2
Ht3YpOqmCiT4+wqiKRFPdQXB0EHhXlRHQGTgWoEeHH/QzfpSZBVnjqg+Cfvkhgj1
kqavPrtMKQjE8t5XvK2NaI3UFIHMGwlJ6bUQUw7J2e3sLgpHMMQjwRzKcmbmzZ4z
j9ZkOHXZko2VER2GVS2AchoVX/dxayLxd27YqtmGhwQdEJtp5ORIPqa5geKLRZEd
2ur/HV0rzGBpbouWf7tj/l3yZfz0ow5l1XvgyY8ORpzuBdM+511lrt5yZHAM2p7o
jxHYczg/9tSv3qeyDD+yDKJKNlyrRyWFr1KQbJTM+EvmmE38v6JPi03o+mDdD4mq
68wrTqxUk0ZWIadEKFuYNtntvZHh4v+yS+FOW3iKV/PsFQWoR742XEBN+CJIhgkN
/YD4XgGqqQZ0DGL81GrKSSvryEvoWhJW5C6tyvUr/y2voD6bUwRLtTEfnalMWEUf
toMdAf5MIBa/+SndAKsoHHo1TjGbSOuabkKYD5+AZTkicVWWiWjQq9LSg3O37fGe
ykaiNZHHTi6hlE1GQryXz8+mqQvLLuy0Pcj63ci0fgYnA6W/MbovSMTLIF/go8h6
mXJqMHtTxQIrimz9blzchp1a14DhUq6hbrRw0gstcQtEcS28T/j1XW8Y6kB7RTPM
XqZ4BYV9jd8uhttNxLqpBwwixH8jb6eILKQz+HWhrHz3SqpaOS39i3OxkLbn7eBm
D2kYeANGXgK0x60tau4SEfBmJzsSD3XVNXBdnq4czjYQ/cwCFF9fYA8soHjoiwbh
k3xOsVzomTZW10WG7RXsx1vX934+ck5f01Kl7zom6lyvfJdarPikR5KgPAtkcdtr
hToWCbbSJhCcHeHdgUmEiK2N5dWL8hm5DLChq10RrhPLaQKe/38dadyZHat81IRd
y9vE/Z52/Raobz0P0Q4HbClboYC9i8+pJjXZ6E0846GMHaMb9ZLB/Udl/avNV2T7
qB0bDlaqt/kslYm26KJ7HRtRDhE362qeFw8ZiDRiKDRa9kOHttioNrst7HNHzRvG
cdQutw4oxXdhI799y957hebpXYzFs1Hqbeo7Eju4P+lubM7JAL2rrfwnGrtL6oi6
qm8iT+6CvEROA+ZfSe+TS9kKjYedM4G0ynbUIPm3do64tmFO9idUMQTvzaWNNozK
JxN8/oE101i/AdVGayluoAu3qY6eUfZ1h4JyF0NMD9WWw6SEN3yNmLE90ahavCce
OUEYGJLLXQVBw+k6Mq/axfnM7SnqLAybbE/qSEvQo8YqXTcp3rIUYorAMyv61Jm5
pjE0tjxSpWhgSmhgr/48KQBH85q3O3tacv3XPXVmD2El/Z1M7wQwmJ6EsgFRWBl5
fNH2yHZJO6tqM+Ezichwl9zxl6mPlSPSfhKmdxKzZ/I=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jywlE1LY0m9ChxSIEsxIf8HnXnNfg75hZMSPMaGfl4v7A41SU2qL5ItFl2Vsfuwb
//53MwjAmlXwiSLU2zAwOBBvr/Wl0jw182lOHkWqBA8bFlUpyOEG51JIbpRsYS/y
kILF0+BllSUmQg0NcRPScwtjeEdpMlzK6gS9k7NgP8ITq0Z2NL7bYyv0fqA2intV
97JTcAMvcmSOkrz3LI5EnB6Z3k4d+5J7AEXsG4EcqoqcLwMpjvaSXu9fzzW8+oWc
TnpgLcIlUsw3iekugrSTJkJGMzTSId2Fu7EjL5Rl2ly5llZEkSkDbxw1vXHt/7Bq
BLyg+jMO5SD4GLigpC6U6A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5904 )
`pragma protect data_block
PlV8TzJaCEpsoxMPlsVaniPzdcKznFKnjhvpT5Ew5TOlkSFuxsV7daR60CPOFfz8
HsJDvadZXm314F5B5LH3o/vYM+iZXy1tCOxlfdxlbhjiMQt7iqKi4eISutT30D8K
K87upDIz87thl7gy2EbRumW/VRD1B47mU6P54T3Q0CDu2u2y1Fbn28UzX5L6EKOH
3LnhVKzGvowJHfBwhRjdyU2MZk3Gw1B87CSeYPAotE5kfm2FIIQ+cb0knGs5P8i3
8t4TxUfSY+F0bAyavZr90bmZl4ynvIgvfs+hl/47qtHWCIId9K+vKZOjL8dGg0sr
08brgi3tYh2tvGYlzwuxfu5o0qhpMZ2t0h9fY7UF1fpywcw4MhE9C4/GvEoVtbww
7Xt+dGvsqLFdYZByTaGpCUWHf0xPzI99mXisRqjR+3Dn5E+0Rb7/FzPseFob0ck7
PLEEhncYz+3ZcZ99HhfXjqLfOF2MlHXbolkJs7zJZ+rvstq45ITMlr8ueOPsH1pk
rp+/DDXlwUeqULzdl3vwTqeezb4LQKL5m628OQq6qu/BcCJ/gtAulw4KSdvxZSuk
czGOXqbAgLc2fABFSE5zuGOGnDRN72ibQHLteCNLVVIiPVjTzVn8wXQl6FonQGu8
IINBPImXv4P+wnQdhaYNMegxSFis2knvQrQqt4/iCxH82s9s2cXQN86gJBpg/9C5
47DcTU/nVWoJke2sP6DtHWbRlGkMMkER9jbqNkFI6CYI4O6DwgGCm3OEsGtGsidj
Fbxox/3PztiKcGkAqX0q2g4VgcZPDEd2YDCyl9BRAmFMdeLwbDrCFLnzv04boNx4
coayUCh3PhK/UNA8O079TuDUXIneyTTKOHq3Z9CHP45R7HxqwkZihK2c4jRmAfAN
6jPi/pTRYQuwyHCnKBD4PB10hr4l/qI17jI7H0vvrjQU2DhjF/93OJvfsblf53qx
XHrcH4q7G9RH7BgmFSSdQYTGEJOFiQe+/a5Wfdks0226/ZIzo2l/yt5rl7IIAQSU
PvR4tTX/gUnDQYlE3ORJQP9Ogd7fyA9LXQKHAbhkQPT80Ku+WhJ+T4Ux3GIFFvml
455oeg9eApGIx7y3DE477K/R0FwQRFBovR7KCfJb/rDx5VYTOT/WATz6puDmPkiI
7xf8R6RY2hO+018N29eaniYANJi3iVZQePSY5HWObZLfcXPWJ0rOPLtkh/lRBs1Q
HvZrvGhrlHs0TjPgP4yxMw5a+YBTIezAPzCDKJWGgoDktsFMuJKLuGIZTX1eFpEy
o9kqKmXgGgLuve4jp1cca134QAlI2vEAKycjgwWYVMDFyXnWep8i8UmqX/WjFipV
9p+dnwCyd5VPbkqtLRj/S8gL4Vgmbb8YDr3zkRErVniVURHwx+VbaxIiS2KgPkOS
g58POfXJFV7cujA0MufaCuoFr8Wwkbd1izheRCl2oC0xbR8H4MEsm1NY0PB1ai3q
t5oXJn7ngVNlhJznhMRKWjnqHcjg8w5Co6tFMnZe5F1mBhfYE5EvmnVvlbyTIdNd
PAlIWBRRJxSrOQJAHiYAcI01QzFpaXiJ+rsZtugRaNkjAiaQgqbU3lWrgmym3SBk
EOky4DNz12CWU8w6+pgZem1aDtpvyTugJM/3T505cO+DjBIuwGKDm1M2mMCtZUGh
la9jqKemwbZkco9YjLtO/x5mDwHIfaZitqHMJk5icrNyjkHDqXtcsZoLAVba1uil
qGtJmoVcH8TR7v3s4i+MWzjDD00ARhN1XlYz1vTnqdQVqCf9G8UUhKSrG0sQhQsT
aNkKqEwh6iwjSZYoft1rJQbloT1LMW5QRflKuBu1Nsq+jcjmoBIlumFPD/b1Cc6p
7exY7XpqPYwS4PnDZVAW/IFxwb5I92tHFYBQSgOqroYugv0/X0O/KT9c6dSf7BUh
S3xeKPGSaqh0rUsSqt+ZcqzVx+SxUV0CfxypZsh+QunKRW/+BekPvUiRKwEV9lhC
Fs9J3k1M6S/LOuNyjFEn5deL5lUvfDo6++qMLuZILC47R6yxYpmNpQklNcviS/0V
jJUuieROVz3egPBjFZb7kfjPgB/PCqHd6DWQIfBMlnl5QRvyph+In3KAlcfIj111
/FjsjDt+2QkPJIMZPUy0hHm1oifXIes5PqWnV476F/Fjogc9MmyPfy4IXyMckbrR
zk6IGOETUlHWvvCbo7284fpuDwnpZhmZgQukiRcNLVnL3BBYTbylVRACnRwNMIus
TdXgASu2xG4dK6Ix/RYeMlpIHvN4X2jzGFitX8iVgTy1j/KoMJuR8I2pdnUUiCjc
HqrOpf+4ccI/I+zb14pPfbjGpfqk3/eh9WV8tUxrB1PJjG9vQIHWmmxxBViec6Oh
Y+29hM2T58MpVHq8Smnq4+KL6EyRI2kmEZ2f50pC9vjAY+3KvPpPlyOXpHXdzBnS
Rk5FSZlt+akbDWh5zijdy1spuXzoU9/zcHwWCqT2iX/nE1/S45akoXIe4qrH0LN7
Sg5aGDI85VUgEAZQalhQUGfNN3sj7zGfZpBJCST4d+XnMKgOh6zte6zDrKng+bFv
oWd8pQ4sg94y5naEWK3xYBh03w/CYw6dPo5DdAbewKbkBVMSAekvdVsV1aG7cxQj
fE5bOEz5cFu4xV+JFGkLLAt9AeiHTMTXn5Bm6fZ+DibxcB1TiP3y2c0yiIGyl+mN
E2akHmyXlgUcfWRuiSY8lLrDOyISzueyfI6ERbX2jChH1LtwkqV4/JU9IJz60S4a
swzLRfDGDWUJkiFD+o8iDEtZjRbX82qfGDkHDW9/6bQqwPhY8Vq/9mPgRLls2uwj
wJ/7EbeQ6D61lRFV0j7uPTe+6AA7I1vzNLguPTNeTOFawapzhXJuUoBAlS+Agk/j
J+sD8k4t6QqWSdEupCiOifL75rolMCvDIxy2b3jxGFG22Y/eRHES+TjjZovkmHMt
ldTPEY+QKDsCVBetl5gB56eLk0Mp36xLSSfczluVl2LhCgJl8SJjDZfwJF2W0Hbb
5ipyA00162dZKt9xuJ1wWJGqfEih2WoXWne7qnc+frBi4J4JvamkNJeJAP5kizi2
11utd1/I20bnnrCjNU62DisCBonh1q0f0JScNbP9iVbzDj3eD/vlhvCyTuOUxa4e
FMRWSuFuEh863Fiscpt8nsWfuYDREMRhliPzHk4C+MA+uw2H2fLHaHCaJ+bhF2fI
ux/mcESfAzlL7drutUiv2bTV+jH9/AzCNxUgPCCHczusWBPNEoNLn/iIJ0OAFUVz
iVzZUwBJYneEAESVgX9wfYOZIRc5mlza35UIDD6IcE5mlI5eUiaw1Dl6p49Jtl08
yyQV5J+3qyxTL2+XJsgSd5eLE4MKPoNUIttMTL6djYm6Vfczh2gXFYoXjLvmj/7m
zHTV+t6kyIlmhyCOFADTaRXo36vK/l9PISKvmtaHula+NAGm9pBTwFrWdndB0yZI
8+vgzNEZCAFtIZYFaeQ/Om2R37KjGL/lKCXtx3o1Q6f8/pfsd6VHDJDB075eQVuN
LIOtOmTWI5H5OBLJ/MuaJNO8IdbJtXwK/z8Q0+vzfoTKnNNz4zgbRr4iB5vGzHyF
NmdvUmuaqoNHWECdpp+RhPPYbYjzQR3sa88H/I3McJISWMuU6OEZmhG/Mov0Dm1c
iwIVMzuTMW9zsfKZ7euKaAe0evCzysmBF6AxZqkM+GnPHMqI5y2pb6SCTk1DBJjR
rK0sGEpBM0jzpm9ic5kM6SSM0XIaGQRXywDZ7HZ2KUUSYaDfOfXOlsMQf4zpAGek
frIpBTj6bYV38Wcvr2OMIjQaJD2Ttv2yhH7npTBMbFVc/tdR920rwuHLyZ+zZaBa
OBnZasfdsfFBkP4jpR/dLSv2v2o7TF5HNeYcecdhBOJ6yBsIVrjtNciLoI2sCHqu
nQpvTzHUzkGiOCYpYtvJxEDuqAs+9io7xqRZPMgxfws8tTp5U8fhKeDmJMY9o16r
uzJa+ImqN2UTvGbaoP5x4X03SLVznNGP7GU9sDpuJsNeFBhKX8Y50j4ghUECKKr9
jChp+8LUcdyNLKc9hsI0OPvuq3VPTdc/Pv/XMmrPlSoZsJ5SqIURJW500FkdMRqx
9UlHThmbUl+d8WZ+hnh2RY4WxV4proPp0kbsp3Tv8ysrDAkR/tx5SSZRbl54e0dF
7mmwVi4JtyP4RAwS8wS6nLT5hapo3R8BwRkIJb22PAsCu/2VrLQySBxOwZa9nLNO
x4d9HCt7GOls//qGQp3SJPdt7riW6Dpn8iFh9/AcKudBByJpnp6Jsy61ZFzBerKe
KAKnnqTmrFjSvAPgXVpnXCbMSbKOq0UGVOrdrfc2gHXyLgsd57ka4UFd9ZfsnOQb
w/4BdI19lZoucLARWBYiZltXqkG0Xn/DwgZbD3wJucUEoVp37oej0G/5GMVOJYIt
CMFHZc+o7mCE0CruoeAPcojuOFQZ6bKdsif+yUxCkC1UQzeWUKSttoxP3cP8jvZw
yUQ5ON9T/L7J0WeSPUGVkkRTQTO9Mh0SyP3dH0REDBZ/T34AL7xpi3giYm/RnvcS
IBvzdYLdmSCf5isrGSXPqynL9sorlyIBiOz9bH2u3FIMhExI2rJLRWd8VQlMlNnA
R9FgBJdDlvX6SsFivJuB0y2atwbtLwJ5vtv33RqzDfXWHWjEWx0Ody6IVE25Txas
VHIs792hUA53jMt93xbpEwbFyY42PzNomraQbP+1zEvPbOKxOptHRC68tcNl3ZdO
qYgsnEpnECYAb9urzF2XsGNyKfJ8SyJC3QP/++ZY8PId7QK4agTNtT61DXqBaUnB
trmpzJGhhToFDYzo0zFpLUn8hJ0T23VFCApkxq2g/qMvKaxyXFg7hv2mOr+BR46o
jGIL5ax+MyrS+ES2ccsQGT7ITeLUuwFoYz6LuVZqLfGI5dDTmJwCeyb2X0N5XvmY
ttCfz/WqxYmCrwWDQflrfxhUUSL53ObMEzqjm2zw3y6V/sf2iT0dgnsUux1ECyoV
wd1onHfWSFn1uuZnmf4qx6rV2WuI5AhDhY7poYZRKVsKBPI93Ug8x0rbX0NN2mop
etTtOZqbw822f5kwD2D3cxdR8hLNun53NxnlkQoWapzceDjfdxXf/YnKul60kqLz
xroqtR5SVGYc5hfIMSzZa/fzFXQSjxot9JoLyh5NgNCDusteZnFAtCMJ9hwdLGqO
oFJdYTz7AWDirGsWpau9dlIW6STkb5KKhyyTr7sdYtY8CVjZJnWUuiKhyk3YWS4c
F6UfgQGavu82m32cezwHp8aZyF/8+iV1RlTEwGJez/FwRHTTni6pJ8v0cF5n4UyZ
8cNy/BfOj3ZH1dZySRmQsH5NfCWA7rRu1QH4NGl7NIseNvo/BX5soG8zZc17O7Ci
8ctQgHNlfwWZ70JrF2ap7Xkhffh8btYRQ3luQTf1p3D21ihPEUGO2e5Wxo9enS81
acYV4tgoLHrQuFHnL3p9CpNoeeDkyW1NwuaOxOFD6Rnl2uyKtWooFZlexgp2e24F
P/YC+hSlDxtSSRNKYcU/xwedVmS9rWgkeY4Ry2woAzhwGaGezsPR0Db/VCYb2vKq
+p/Jmu8n5i3xwybUeCZag1rdCG7HQMd6pvZ/+O2kCTb7N9tbHfp/Mi9ZPsrC2S2p
hZn96ZfRczQI8BNNc8vvSMLVb8iII0xFEonlIOiggDDF0rTEztclSbHrjTK/zMJO
qZGOFbgWaQSpOYvQs0T+ZkUcc4EK5YdUjZcqXo5AA1xteW1nic3ojXD7TbStF67+
MZ/VBGYxyOWisFT71wpIJ9U7R/jSTcF2yvWMWwDlzO0Ii9Gw80ehGa/pee5ENVf8
PtjiN+Bv7Dr/Nd16+umSc/85HEV222XAM1fwj6Qb97peIkI4+hjgMmbPjEdI5NRF
mD6BAxoK+fKc2/BwSu8pL3/pyqKauNCaj7gYdwwz2Rk+SZDvjTRwZydXGpggMw4o
lNu9SBLG6q0zU7Q6D28ChbgD20VA740nGFMQ7JsYUoJbF7i6ctXa92i222WFk2oG
2d7Nh3nXF1+mYwyLBlhAqizkIBghLZFlSN/cSgLAXor8XsB3D7oyaXZ5nDHBjE0c
hoZuLghMKYSWpsuKQ56ghU8MZgvzw5Hn52ST866LRgfwInpNBWyBsZJOhbuLK9Oq
gYXqtWCgEMecztK3Gpvy/vmqhYc+QCLoxd11IXxR4B0Wh3v2yPAWFVWntTwDISAg
H7J8KEodmNlr/Kww622Ec+30JeFotI/CiAnxtieAJORaOC38cVZpVqI12fmqTUtf
fPrzzmLrLtlcssjxhpRk94chY+YfyaOOd+QHJTQlzu8eZOki/4bURI/4qygWWdlS
vpQ4vvFtQMU4vuNrFL97caPax3BEyz1//zY7debZFWvpW1yd8X5cNg3+7IWX+oa4
SN0OkdLw4EAKJtswMwQTiNDZQmjy4Ar2OkMzULxr9GBEXDAYCoESO5wKGpbdN7R3
LqKCAhjaenaDdhcDENq8lfmI8V7i4C8Eltn08C2v4MC7QCdRClrmdbS3UJDJ1hLh
hrvpAoHevEVYA06EgX5l9KWf/z9nvVZQnItO6qAQ33MyHH4aTUch3eLsY0ptelr8
tBR0VbzpeIVxCsUig/IdiYQZQVYg8m0Ap20NrFkhWWyLNiAuORitoeaURnV8qNWO
yJTKv9Uke1vu9dw74lQGx6y/s61U8KXrOlxI597W2+7xS6XhqjYE03VTp2Crqu7A
bJ4V1zqzDzJsS/Fbx/p9V6++VPxALeo1FGL/hERk3oA+icydHRchGWuhy1mTZYmT
uhnKcFKv7SvJ2wa5GPXX5qXb/+meIe7XGrM7KbAURkklXA0BkvAobdyzo4VZ1QFy
vSbWI8gQznmuOe6CvyDMBDltscFvsSwcg5P8fh+J97+yKUf9d5dKt6Ajv59KGXeV
L30JYvzVk3004nO8OMQxKWEi3cvGexwBGamzjEt4lpQAdYhzMw4cAa5/tkYNOKn4
LpHuvvXk1Hrl3OihZKjKmL82DVnbJsYKBukuJpFoiGBmeAQgXBmYhjxBywAFtAIr
PaJJF9lynxadziJiWU+g1AdDkJrUrlh8HEO4ZI+J+uOqtMtKWsKjlAYnNWzrAKnv
ub9sW8OhK9yehDMrzMKUolNVO0czjobUCfST4e42uQXWJZbtMfCRu+uE1e1Sqd16
UHEnWx8/5JMddUx8J0gKJYqJfZj74EweBSxDNclEn4DXyfYJB8gdwN5M9rKMaw8P
ZXzHsLZ5M3AgSwI6EAShadO6xPEUicB74GjXRB0nddKh5MxIXF9Ahiip0ZWf90P2
7StUJgMRurnmKfGm4h/GoHYLzg/OSPWh5R170TpyOyQaAOM+GJ8WPzv1H9TGdWBS
Wyu1CE3uonmDl3sP4TxxwwEpom6iA0eSX5StXUxxF5Wku4OgOT3Z0mt2w9jLZcE6
JsrPDEkgKGAC/1ipGA5NFJi1RxDNkLUmj2JetS9/YrNd0n4NnvZT39yWJiqdVp5P
3bcCd71TsCsMJnubPBf96l2C4dxEHBj8fe2ZAQMyuPLPwHDc+TfUrwASPWCR1ELu
6cjZ1Dlc0xn/AWhjGVhZYU/llGctJXxU1F4WQme2wDK+WhIQpKEn6oaGjmhLUkq+
1e9Vtw6YPNReglfRlk1r0+QLwJ5UWGxHGrVGEi8hLIf/ffxIP+MWJAy5NAIRTB6g
/nSImEmwuwY6rPi0wiowF5B1g8OlaBJCV6KGzWyCVrjMOg5v2PTfe03xWep4Q1HJ
nfjBunwoIrpj3cDFZLq04YbmHyPRms175zunvPAshoYQ0xwMXbtpJTm4CNIp3MTB
Wmsl4/wuP7i/m53Fx4pfSMB0i+Cwh/bKMWrk1m6Usaa+OPjkp/u5Mw02HYEk6cjQ
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Zk6lCXi8elIliv0moIc64CCWoTfYCCkPo3DA2O1Yr6XSp3C4rZKW398opGMa5J6P
Qb7Qye5wZfsw35AlxqUYy8/flul0HBsuO+NVx3vOl9jF5GW6/QSEbc9eHn0wItNE
GSbfye7xqzeIhewMLsd6eyIIQlLKmCkqysV+AMyGFUlZBuRey9GxAX3tJZGghI3n
m9/j+yVUQ/UUDSFJTY6U1J6o9+C9O9+Lu/i+YOLJGp7fZlACOfoG7Th4lcFiEMWr
nb0MwhH48RnDt7jV1APZ7QjaciRaBBO4N5x6DWVTEsg/ZecOjGMcKqxMA6piNMCM
4P5yATcMN/whkb7MDmihyg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7648 )
`pragma protect data_block
GycBb64HepBesJi9XjOqkcH96j8hchBIznMZl+aygFR3tsOXobq+JoUbccAadvDp
sm+ElnmSj26vgJF/bXvziCAgaORi99pr6/rJbsMH27+ElxHy5FtSj10ZGS+RgtBE
NxDO6NT2QOMdeEFIBL6DLE5s9lwoY7kN8Gyo83Z8ZjO+Gt03YB0CcSKdlc+g27lm
RWFMkAEOOQwXC4HArmPGXl8khYlsfehtpeM4LNiMK7Ui8Fpv9YR0ejMzmI50FTDU
mD6323vovRCru5pPeTyYcxai5BMMAqQiylFQekBx3Ha0MbD8lYUdCOMHlMImREQF
Cb9uUg4Zy+Rk8sNTy9ZDCdwkIk+IFSaRh5PQUMDLGy1tHDSkcR8ex2cGxNZmyf8U
acNFsVA7Z7kMElyA9wpJ0co1VgYIeOseMhJWeXlIxgUoZGJx1dAsRC59IBSi0iH4
TR1g5jy+FQ8MGvuSDxWMcQFn5kBNWgV0ZkKG9BAqsKcEfr44k8dftlrmQofBWb5U
7duW7UY/LlvmUDxDOntuIOU3qCdZGXHqFiNQMZpzoPp5vc7rfHzLrljFtgesF/4k
FGOdM5lBrUipAXELKVE6Kd0l9W9SEHtFbnyiMnQtp2zpXJvmZwf0HLy8LJ35FbWs
DrHY5OWqRo9XmrOX96B6dQjlwtrwJUdWFZaD8zLpeRd2oB9jkjUOADD1JGlKcOaC
4xZoNPLmRoYABZzqCEKvzSCY5vpeYlcozD4FbcdTT+B8YIzwcwa8lLXe89V6rRsQ
rmS/MvlYTFYN+esw0rcB9YyC3+yUIVhb8k8zRnn8jXLEuCDo9OhAtPL2Mc1HMxE8
o8r40KIisaGG1JS8ABTmEEPFgAEDjeSilj/7Y+l0Ojot1bVwPjNuQ5K75N3Yyu3a
SRxH+6OrGeoF2frRn1B4XtXRuxM/rmHs3K57fB9QuUHkitLDYSYPAZHU+xOpUde1
u+DnSBRPC9t120whoumwdDZJ5yISGDx8OmLjllCPtjZSEs9bxWMx0cWvwawZbdy9
tCgPg6qS3ugEd8S7ecPNJVSxgIN4bP/yBV7fJgONKbwxacDATXYVv+Om2G58wfS0
rB29e4kn7+7ryk8s/DH8ycLJjrdetSJ/Truoh/HENr4D9w0qzFCGen+yvIH4Ux82
AL1qlIGYJRNimwjys8RUfZlofGNgFFhP2z+aeYXrWByp4Xvuvf/tp4NS62wt421H
0Mj2fH1uu4S8lhYyYqOFfZMRMICfRg+JK0ImpBI8XcdYv+BC1VF+9SRuNAZZSeg7
lfoVQkdZu/Xs7vViXPXS6KL+Hk957eURhjCL+DSWMl3rlF6PabSndD7MfjY7f29f
yMWRHjrPqPxf2Y/R5b8dABeViJQsCo7/UEPT8TFkTGaEuqgemdzDrmKBfcsy2PEH
X1rWUK/fulpLaAjTzXbdSLImCoJtwQ59O8HzTw5NVXz6scWNBOYgwT7SQwo97Mc9
yY54NCRlZ1/TUhFhEYiRmC2O5MfnpV2W5FTW+L0clZ//R8LQjAcne/NIpXr7Cdzl
CBR6DekfGUeKX4mKlyputJIymMbt17AsXor9Pr9qz+18GglXCA5BuNOdu0MHrXc0
ugHF/vjXLkU9hQ1PHTAyxnLQqH7Cg5yTnr9OvNmlZrtbkFwPSDUo6smGwwIya0Am
1ORCYpC4/1tzAOr45RkweR/lad9l0fG0VVpU1tGy40iiS9z0UluDBtAFaEAdaUiO
Ocj+w3HYxQgmyIypipx/BFYHJ7hVfPK55u3V2z8RarOUYJ84V0W+R7jpbaQbMwHt
1Cp+UwrcO9i9EAVA8b+VsbvDs9ZeJIthOVnbJwwEupZVMJSPZwOIrqOlpg/R2sbI
8OId0fnlbGfEMPA0fv+Y9QJmn77N9nUnd6kdbcLWWCSr7UkOe4o3osrRoMcIqd0I
GqWkkPvIOEzuV++wepSXtJxGTpjbeK5waZ4NUgG88mLVbMttY7/ZM7jwFIeENYS7
W8j9sUsH4nl0PU83SE2ruuv75lvazg4sD3bWCmfdcF/UbOtK1yWPLqN4BsV39MXx
0bp5OKgr9NRQga/NiFqB3TrJAM46QiOs4vehh7drsyL8Nsa001yKRxteV42hsTgH
fH8nW2cbZsQTodeGu6EbDR33VFbulrp1d36+cxrEUUDtV4ep7WNZJQbpZ3kP2roR
KKe4+5Lg8oCh6vuuF2YwdKBdu06hwsclnfHxLbaWVhGjRJu8eD3nZWaG8eLRMFFi
HDfG4wG0Oxi/aZIQ574W/A46H3vobYgXKKu6VJEsDRaKY0EuNwy1m7yJIvJBe5e4
WtO+oUnBJ+fz62Q5sJix453kkfrehjBxanzMH9jZhGSwoT7U5p2MaA9NwKhnsmT+
UYNRApj8xaFUbAys49V0NhXgqpbcI8bDZKkg1oSmlJJQD+uRHCJIL3PAYly0jG3P
zTucCvZfm19sZSd3ntbGqVujLW1N9LW2agIG/DUT9L9XA42rwxbY/3i6hW+2Ct97
+boeVsVpLDr5lIg7D5l3gA3Dzdaj3ah7uDIMtYjNiIJGmeDNwTIO5JpLBJu9JpZZ
mMiM4NZRNlh6BIg3nM7HgQC3kZZYohDDIG1/2Hgp4NrYh+p/fYiGui8CazJn0G7U
XNIjMYiuZVhj1JWUbJjBUsatqqN68pHyJLwxUYGuSlF9WzC3RAA8uCRhsro8z9TQ
jW++6NPhhOkwp9QQpVVL8FU+02PTxRRNDQP/oArlCoKMaVaZCsahGnUOvPFfkJJ4
UjH2AQIaDxOUhB8YYkNf+r1zl7l7FwrgwIS0g5eSgVTZH3M/pCJTN1IuJyaicT9j
sG5u1EKwlKTfBELa47EYd44jYq1oTYERFlLIqWbhhaX9qWqm96MCSGFk3prDsbK6
xx3JLVh/fqVSfxI4tCp3rAu3Hs8jTllw6oAbjqUUcpH2MaxbrGaY+wrTtT6XLVTO
IwRg5Cfs1HJEW6ubjHYB6a4fiNR+71WqBAnaSCscN3K0qgbd3NRezuUIBvty2Nwx
ZrNL3xWkJ2ZSOCX4Vp/gdeSCeah5TNPmIR55SkUGjilLWp6Z536CL/1lHzsT+jbL
G0V2/jSoXhIubys6rMIPRIh0EpAkj/P0Qn/wVQ6puCBKXHBEQoeglb+j/JhEK5Kp
so2zecx0hdD0+O3wRcSM+UDJiVaHNEyikH7iRj4xqIAQF5FnLu0n8+W0rRzJkVZ/
lAQKHgdV16M6sdhEAnbyVIch8Yw/Po/J0zfCFfGCFQGCF8f5oRNlSZVNr5NtAZUp
sxbpgaM8cCUmUecYqSsKk3Uzur6Lg1k+Wuw/kpmiSaCCZcXENvV9OngrJ+jGfkbf
G/lQ9ieyX91pgk9yrjrNStYRLL1cPgahiCZD8yhSDrC+jTwO+fbSiEdxYWiMa1YE
2vyqajPwtthQ4qNMvAhtoXsRrMVxGGhwmW6/oBR4Yaby8xkLqgi8RUsphNO91Yun
JT6qfEOnjRZopjqrHPrxZHAOAAtBs2vsKWXidis8CfsPlcTR8rnyCIlTxBbO8zYw
9mcEBvqF4mpCeTn3idyMcwx+ChU1oa9/wUpd8QVsU2Wo02UaVHLOpmH2KR39XdA9
W4ImlcFm67Xcb2sRX3sOR7LlQcNsmkPyjglaki0GXmXGn1Q70g7nRAEZH09jKrc8
G9basSqTi0I16OiK43lItFL2AR+R5yTffVYl9hUTbqKNJvhbG1k54t2NI9+QGfnr
HJUsJmDofSjgks2KeHKVrtYHgqbNeu1CHC5D33m/mHxROSodIeq0RjFtwJairubC
dZqqkClPPkKjFJQD+GEbOn6JtejraMQ6cEB+HzAe5ecTBWBT+WE65xR2JlyLu0V0
ILgbKmqK22RJLRHzAKn8xlv3iqg8j5A/5mVmoIzZJ95gbxww+kr5G48vtv5Cjrt5
58kqYLLbMP1fTizXgtjw5YIL+LNvGLD3pdbkjZlXew9yCxQpfMQ3ckH7CONxZs3W
/Vyw0wlgGoUeFB4G6UgmZnM5ENAT85XtsabDdoINP9XYMd7ExRNcLtYCzZBeiUtK
rrr22qHmFCHM7mk8Phry9b+9erL1UkCoILW0HzI4fftSyz8zCAL3+6ExsmBb/B4z
WY/KfKN6YoqoETt2NCaEfTuX608j/WCzdqg26+HqxyfmpLQm3BbnaCIRuG8XUZit
5GPN8+Ea7wKzylPqixJjwdipWXDZio91zo/yzVcVMs3mxuvI8k8CEMRGmh1WWDwN
N5y+v2CbHrgDiMJEkoyg8iB64YmhMtnovarDxUZOfIN2tQg3NKGrqtLhZ+xxcIqW
TcsHtZZLfOxga80YYHv96O+wjTl69Yp0axZlwoeT6lA9QRZyaf9UknswvpUsJmNo
tqyaDHGU4UtRXIAn4oQvIDMwZO/2wOHxgW9j4w+NlL/MkaZt9J7inIzdQ94VCbVe
6296n/0KeVONwkXEi7KLIBcPDZrr1MoX/gbrzY6RL/Z1zLhaEyx15YcnUHh0/13p
ReWAmoh9rlOtF1oG9ZCfIgYGSUc6BeJ7oXmjWNj13VQOTnHJAvNnDZRTV7vmbJNp
LCiITefan5gQx2oNHUd6kqoc+M+W8EKWXanAgtt2s7ZwKMzd6hUwIqh4AyQpkTcf
jANWccUUv+0Toihazo3X7cLKg5D4N+HLWpaxk0dskqEVZluGZmcWdkmJBy42HveH
NFb6RS1iFi4tzhB/PNCrU1JIrdCeS77Scnw7WwIYtPya0B4lUWssivwfqIhAkPp5
t0CC+4tKG4nm865low6YD4O7FoQUC+H9mm8fGCqgfGmBQCkWChNYMeLZUd5sirTz
mS/WZdZ46oJ0sWudLPzbqb87VrNOZnFIpveDm32h+1BCI0bPuP/y8bbj2lUIcR/l
NgfihFHHNr4YlTMhLq4axw9noqXyoWURo5ezKsrd/Ch1tWASUyxZOfu72mdCQOqh
N0aO41nUamp0LfTBjCJUcDz+/muQ9VsQVAV/qI9QknFEd97MfPh99EZsyjONOaKZ
Gk9Xi9w53P6Q8T9j1NYUBa9+WLEV/o7wxPl0lIRXx2/Y03P0TrH9avpb5tmVYS7e
99FYWz/IhFZT05Tw7i3RTf9ymZuyAFJ+MCX/8H/PxYKvzAGY5Bdt2GPMDooTWW2a
uRIBelnzW1k3nU5DkTwvB+x6C/Z/Jwg8m17/ah9flrRAzcvPhrq8Z5dtEbwCguAg
+NopB7/9qnMsp/0xW4PeGlpik89e19eBEbqfUlB6f9DOeAUWxneU9dKSQ27XyiAM
xTIgKxsqJ6Tb99G7lXBCIBxS9KRf3eExsUDZp0sLiQ73Sq6/QpzEVGKQVMVz8ghI
XzobLflGJYbR7h3Mxhh9Q8o/CDVco9d09KYI0BxEgjQKHBSdMcOTx3C5tH1Blq9z
w8da1GqoK+K4HOEPSB1bQ8Oqykh9F48Mz5yf923jpbLJnQZxMy9NYsToSb0+D3tx
n64Yyh5N0c1Jq3nGmvrTkMnFYC5P2sNe6KJARkcEwPgnLY+4AuXEtvBSO0BFjZ3B
P6Rs3QZhYsotUDPRZ43xpT4feg0dsUkP0jaJuItvlFMe3AzTL2L8eQuP/a6xWy4v
kJgNZUW+VvuXDw2fjaPSk2+5p92hBe9MPMRR9/uqOBzzsAFoSORMKzr2WaGNqUt1
/U2CZnUrkvWYQFF/wXuP5yzhS+FlQLrdZZ4svfapfKCKhGHsnUFjHO/9RwzQq+qp
Fl6mO1MtXOHlEIXgX0Pekl/X/5ncdCjcA6CQIUMqG2GMGqwBuaExRKM0AGaeNlDi
xU8MpXpzRkRbNQ4DYg8r+ifuXgl+m9aiF8qY7mlUQ+OM19BOb51c1rBP+LdPa2hV
OcELfzftyVQA2kuN2YfDWNoiRLGXaBOoi7WWUbV1JgRvBSeOZR8MAaOpMVLY8DV4
9+TzTDXrNO7iovjqidjG2Rs2LnE2JT7g6zrXS6jc4TlMaXfrWkhSZlpB3YdAXmzd
TVke7ewYXYK1P//NshDFqGACj2d5eL0jqQOyvbQa16fRaIGgtaq+eF2aq5MvF8fj
a84CFcOyFAycHWsakxGYOJXiyncLb9mbjsRdw6ESaOL/m5gfXAW0GSXkTVweYiDI
8naUI5kUXOCexlRj54Mjk67ATFcYwO+RPNJ1CBQzQCudY2BRe/oiXZFo2B76H7kJ
JIZzTH/HQU0aXIG1eAqRM/vVYjOZf/rSGsRHzooEhDTFMJ9+wKuP3dkS5MvbDi/t
rbU9Fh57PaiMzDfmvLklVxI+bN2d9bCtcc1me2tqhLWelu2f9gRqbTL2JUqEgWFl
/f3oux0XwLpwH4VKUt87WeAKooHIVhjyH9x0/Cc8GyS+UBZCNRSxE1ED6GqZ7cia
C1UdwvNy+6Umbt4PXfW/74AImP6LEEM95KXBWsRhQGUju4RZRfKHRtN4O62XZUxq
Oa2r0K6qrHTxvKyWsBxWtdYksEZjzQbwt8kFD76aslJSj0SrWFQxzJqpiYwMdFol
qMivDeEF4SYEn5iGe6NzukSHh8dhcywYs20L2F9VtvdRvuLGslSQkk2V9fTVggA8
2TSwLTphmWzC0oX3OCntw1FxGqEHBrc1/o5KbVORuZ6dDKFCma1slvd4Eny09slT
A4cVyAuaEcbLo9RvkHW7lZ5WKB7HFkDE84Z+hoadsh3jWwBLwcvrS7b3yzhSwP7B
kvenLNewMRPj8/Rv7ZCpjNqiObr4bLvKZIQwqEZKyFW5UEKLedj1PeZhuCQCtCEg
U8Fy5dNO9cEv0sfOmBLrccKA5RYGLPmPIp0dCXlgn87C9YUdKGfKVUrvfNNrvUa9
blmcoJkOl2Dxo9N2gOi0DWrrWvKHaDA3PYQXoR+C7GT2cMEiR2fsE5TiZBM43B0J
MBjKwI+JzToCJ8K00Q4UYt9yu0jsmvSzWHxrVLgI6jbmro9UEqmr9kimfwgAAS47
BJXLsco21gG0L4Cq9vzlMjFmRMJ0+ITssNErAgAOXNlCaBy/4h9xNER3SHhf7U67
6KyP5RLWsnaKDnheRIIoD384VppI1RGNN1WQgaxhgZykVLzKkzbxXOsrA/FvMtgP
9Q+tMhvud94FDrlcIMl+JWrZJHocij1nP8OCyAqp+3COIXdJGRpHBYHzUh/+ZTPU
/I+tSbj5a3mi0CEIChV3w7adF9bQjgt5O6J0keQ5HOb5CPocJn/coY3qQ0OD9zg4
Hb3Sf14ZpaPmNUEjje/4090ziyCq2ga6EOe7t5TzvCjqZvayxRfngpLSX57hRmRF
ZMcJyqcOnX71Cxc+yULtXtfsmZh1szXNcuhNvP30jDgSyVCV2TGGhTOxzPdmGncz
WezqBh+PVIrFv1Rn/9qwRyNIoTDpGTgkOWLh2YdpNTv0kjw8Zcci3dAZwglu0XAO
I3k4bzw1+beopNaStvtcqdYjnsu1yta5zVzaw1y9bi6b8wpoaorfv6j/Xa+RlS5S
3qzLVtVhSzQ6fADaPAP/aJxAdlQ8eIHEP+ice6XPy/mvAuUhSl1c2tFaSz/w07nc
8Vzxr9DhbeDlpun2gX0LA77F+llNCUHf0xOR9ApQ9tHpCG2J3NXsIxmoJOgkzwZf
RG48evw+21zF/G89bQwgOxxCksffObrm68FOZKm1D31lRBpIc5vamx8sbUBJVYcH
3vXX4TEEOM7XFoucMBgxhTB3RO+ATTzVEXyzm06l1UlM6hjOTZNC2ynKoN4jKY4P
jbv+ez7ITbHPxIu8GJ/2mD2iPDU8K3hr6La2CWyhEjizh+HMZH7MTPFJuk31E5/D
sUK2/4wSXa42Ew3PsPIz6NMjFJYBxVyyjfGYwCNnwh2bd49b5GCl8CsosVRR7mrB
ktBgI+Ugub89ZU07XOItUgGb/dqbOZD1wCbI84qFK8XCmLKQ10QKDhL/f+qnJ9Is
NZ7bNL/1VC4ZUf4g+gHEIik2cTfIUGhoGhYpgKxL0SfWEGc41fsZ09YlXbNMm759
qDLyzhm4CganDw0h3O2ziUY+r2754EdQG5JJo78CJUiefWjBw/aLgygej4BqyQBX
GVm/KfBzeY9KFJ5GE90Zceot/+S5qimL2ltbhTQL1RH7vwv9RhTJycxqg5swmkLU
iDXNhyiSeIiprOjSD8nZzpNE8kojilf2lC3HVLLkv7wSlRVaVX0gdfbEcRfoR+KA
a47+Wgy3xsR83HGhgi43wSG8+jabJpyjRjN2pNk/p/S/vdNSV47jVvf9TiKFPlVx
NCI8maXg439LENzv4cfTJK36zplNBoPEUcSxAaFxi3jQZLBUl4p84hC5ItfJH1Yy
0zB8mevFkBAD998V7ilp96GYBSzm/QJONPpg6/s7WjChguMKU18pjNKdBXUqv9qK
YEpO7ielsFzyKDbRFSGga5LUVSghdQrk+rBvIxfDNqAwCe0xW3ubyuX4bNyEVJUz
kIJRt+5bK3/g/Ki8rpvo+50N4/8mDtNTcW3oJf9tBNvyW36HjFniNb2CcBQn7r75
bdRQLkJSmtKL0PcvgNhES5MZ/1ubW8gT8VpV5Ut8zVd+MIfj9oRioPztcjxI+RHt
kCHnO3gZU6K0jgez9TvloWtWrwWDLD2TN9LIeJDwIlzXHnK+PS2re2MKjDq0gBwS
t5a+JzP1BV83Pl1g0BC7z1261dSg2SdC7aCAM0KQPRMrIqkexzHUc0XJ//YIm1Xc
tTnrLbPZsupMtpjEp03TS7ebAuU/ToB5BclJGQlSaQMaD0ZrkK9OZ3wz27OExpEy
PMmKQ1HQpx0Tic9TWogP/I53KZT3CcleCi26Sg/59iSbUB6Y8Xtk/MXBqN54LOpm
kjszWwvR4Q/i17rPfUGvpaf9xOd+7Dsr7nJgciYAevHXYeOaFlYdG9E0orvabLIP
b4Tt5g+K7jGYn2dE2XBdADjpYL3AnzWdkcasRoRHlJ4oBvGeZagxfqWa8zvYBiJ8
Ud0qE00Zei2R3CGYogBT7h6IT4OIo/4pvHiRLbWIajftLiVrFWAYFsEPkM5OmURK
MI6roNCs1fEhl4cKhFBvwdLJvMSAyb9FS5rog8NriEAyO8BldvulDwjFUANCvkrZ
jP8CccT9J4M+nKtitavCNkSCQrqu1lDwrSxz720YqKPZDySp3q7ebkWxCRO8tJqT
JjjHUBP9s1vwKjT63f6FzEPyCZbfusMByUl1AaDX7HA3DEEJ8z1ANl0jqAVr7Oij
NvnQul0IZceHvju+sPXc6Nsqkog7msaNGtnk4F8cfOoPeljYcHZ1xqk+fb+G0xdE
srrb/DNE/rcb2OiTQQr0mdKgm+2Npjtb7i9piJT4XbL12InnxYb7SY0+FtasFpXu
cnHyrf7cVPAMg9oaTqBCwfn4+fcj4fzh8jzrPa8UjquOTPns4xcNNjMyemhXKQko
z67Hs7mLVwMVN6H/DDOfaZ4fRtmnX6eOZVUp2UOmbSay2wuBlm/Dtyrcn2CqcnCS
Zgumqc5bDITC+bOUYDq3mMYj/2twqEMdPNeAYpD2Gy80uh19SM41mm34hSc+x/bM
varMATip9xY7osl6Wj7KNn6JQOqp1iqDfWpjvPA1I82Hv2NQd1Rr+oecX8tW4hJy
XTWaMc3GwPDwRW14SJd286l5AOIE9QDFXNT0Lefa4c543uGHCpfau7CfsWfLU7wj
TgK2oBnqJ8RsM7HffDN/DGS3EDUKNLHiNylTFp730pccvFQ4TaZQHTNE7t1KunXV
QOteJGOih87XIhHzXJswBb5gMhK4WGpP7yFK67R6Pcic8RVBJoS05k0V/o/T2j62
PeYTGps/RfEdFp1i75ORfViPR9Zgm5ZPUF0dlnjOMlcTVg5AznukbM4rHg7KFzQZ
sXJ3PndXY2lu/2fm8CbblJF/y+bJg5+ChwSS3wU0WJNyEpCtG07i14hfynQZH8Za
VcEYckJihNGR56CU8L/3i2L1aBsuCB1DuukTxriKpa+MCyFTVAUKXMbLCH7cs7Ei
uJJ7bSPxd3eWYSNjdsZcBKM8auhHUTV5IlS2L4rduquF7UL5LCW06S12cd3uypEr
P7L+y2x2IX8S5VpYmuBeZ86qalkiibwdlsEIMW5JoWhCdK9IDvNv9I/9NQn1wFLh
X5ooTWMBLcnr4juUTzdteoSdZoldXdiYOzhLWlme/J+hpVG+quddYgLGKMIZcRak
RvqI+mkfmz1NLIOxQeuqrwOk2ppHk9+waKTAX4lofpv4qKD+NvE2IQk8ebA0fPlM
u7URz3J1Iz68DZOBoOMidw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cCvD7GzOG2pPE5p1RoZYTAMUgUv59xJlcFbeni4GYZjTvEzbYdceZvcXwWmKkoEZ
g/U/MQoyH6vH+QEP6yDR+OgDPvieg44aIRasQwZ/roD3DLAMUF76t2EPamWltxLK
FykCYD5KksJhUexlaZgOtgllq6+Fm7Cdjvx3Yj9vSjWtQIURqr09vVIuu84lzDPO
vIfPlTsJU7SfVZZdqsgeKSLUFOwCh6wHSho8Q7HwFcRekNB7Z1OWPWmIcgZN+pZS
DojI9AK7zbyXujMb74z+eJ5cs5JmGTeTpZO5xJyTjTU7ldaU9v/H5AOpmsgvzycr
ra9evtE0mMPA0jylBLxDYQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5632 )
`pragma protect data_block
vKAd3glSfBBDU4WRd04RyF7ZY08SqrE9qOnGGUpV87QwuV+a/6QxnTLfqCifx2fI
imtKaUKK0HSDLwyU8nqGCuC8KWpnAg8Hgj15jd6FF42qvp26WZ6vNSNcbPmWrKDt
XIhgsvNkGWuBnUxl5K/3Ymw9bq0MFOaoZtgUqOPjdltCJIu35K/FmIzk37IWcbNR
uHYO1fHvqg6j8Ew6b0l1KaIbcA8KedIg0YwwKsRfRBBunoEfzyeelmFCTek3WiKz
WOoTIE+qwJnqH7FuxxkZfG4zbBJGeCYmtfxmT6lKulBat6Loag6ZYhPhMCLHgOGF
znBke2yQIFi27kxRd2440GCX6/5RmHJpkVlP7pdfEEC1DZeWeyK8nofXnpMd68dx
Nl2fEcm/v+MdkDIR1HzZF0YnJtVeRYS29EFCzK/Yf7HHfB9LK5Q1pPKFNJXV82bs
jz3R8BqKp6QTPDzunSW5XjmR3K9n7Lz/BWgQYF4yLKWyzDNa3jTedugOS0JoxDF9
unIQPak/TtYOAJ0QHc3Yoo2dD4cbaTUjpymlwnrjnET5WlaqmJDnU6HX1rdFLjvB
DBFSXo+oDc3/swTZHo+6gVM3ZfDRJYPa3DVzpLKThCi3jz9bT10hGs7R6eChogsL
NLP0WjThRlXuYOkDWgGu726KJswYAJ+6+MvvVEqrDvKbWz51Ns7yL8dQ7X1HQUr9
PilADt5ZUaps4cMr+SfBwzx4VfqC22yRn6SnvI+H1ErnmcGaeOap2ZJAEyucMTPu
hpB5vsIsBQI+rKw2kn+ziL/iTMmeO3bfTI8D9JLVlWIk9E0GXkqfGepfoLqP1Dla
9BWGetJ4BNYG846AY+PjrY4B9GJZ6eGK4auK3KZrhoFv8oxj6CuWu/rdAmbFzK/5
w7nDpS5c8frG809fp6D7ic2Bn4AkFgBRKBjsJHQib0UpmEJHAwf7EtJcKJwp05q/
7bqQDvjSND0iWzI5KPpsfT2Imu+Kjvs0POth+hYEAbieGiL06993ofxmskVXNNSp
4cPCk80pbguRrbnzWYW/pD9MmJ+fuU3xxu4QaZmERswSdlt5wC5SKFbqTpbLYtXt
UEzi5SUPqxfBUo1e73jM6tUMSIO4bDOpMw6Sx58R6DV1GJnieUi9SFvJQYzhZG43
ldVcX+fmr5KAk8wsyyeaX/kOPfJ9N2seQnSI1cXgLvSX8bimQHAPwfuM3juxG8Iw
jeZIuK87HyW88TxdwePMDGTVJZ6AgmF5stMBFVwStJBp1ZPsWaOMMB4swx155OYk
zLveDbJj/2GrPsfScLCKm+cYj2dxs0egadETMNuLJutRuPIF1LdY4dQHev1SbEjV
wu1kUpcgNPfQnATsGJ69pBRw3lvV/C7EB59B3dMkHhs2Q/yS8pujIkb7mSG1XZVY
nqrXApAyeKuR9x/aI9SJF0bI/An37xmH2efDXNDgnOSxA1RVqy/JcrK+UiQ7t3eL
1ROSHIFrN1oDyCvBe2bMqWrJ6gSDZcxB1fsi8SeLCT1GSTv+OdFfdnYc6Rgpie/6
gBCVNsPEDYHs/kemu536ZKkuwcja3+pr8FIEJ1Z4poD0Up3+rP2a1jvMN1motsSo
TscMYncwlrK4x5vOxpPinTCGKHBUmL4z8baxEBH37aBmEldeKnH0QSaFr5Z5x3yE
Yiu6GJ1q3/8ZlZF+kwqTt9F0swOysJOyzq1eGEcZfQANmvumaqJkexE+wYZKIHEx
XLNNIXJwZkcMO3gSWl76znV3zZ9LaLBZOgf23Yh6KPnXu28JG12LShQAXIAhviqe
lmfG/6xxwaxBAl6KtDilAksdTEdzDNWFWjTXrj7MzCGY7TjhLmcatn4EE3+hCgU4
h06Hsdj4+t1oRCVnts2NDU5TADgalnn5y+L1O/1i6y9AFCNnwIm65dJndgtgx7Nk
yKWRRZBGcdItIARLQ2yxdGEQOoLLu2Z8PqEnuhDdTl/2I8+urCr1lEnp+RWlkfQs
Hy0y5KF9wmFiGZZhCTSQRHzXgshm+NaH9gsFCVHtBECKHIXtO0+j0uBQgjI3V/zH
GmS2hgt0JFGdD9j1Kq2DfDDYgfxp08sKwDMXJ489/O8se8DJe5Acb15oiGtQGr1x
xq7u9g1Dih/vRXf6E2OvEKWESEy3UEbEJV9YZUFOsHHZVk+1RH64npaBevmELJKU
A8yWIn1jakuWJ+vfh8s44zYizOnVnAyHVU6EdclejeZTTgrLK5196FIS3V2zGEua
+LCbWlkdiXq4wtI/m0Zqu96J85WtxFQiCWNpepqXt9/8Jz7aGl4gSqJRbGt5S0sV
WZKqvjtMjsfjJ8HRHu2p20Yljq0kUI7S8EfXsC6s4RcQW3NXYqksxe3KDzUKUqNm
3vhJ63bbBC964BgNWdFZkiiDoDws4d+AxTht5z8m6dfkLHzAukX9T3LevB/zkmn2
GOAkTebrC+Wp+CXr+yuCOy/Cjt5zfyf/Vj5CixFy/oREsfGYGder2EUlgdgWTN4i
KdYptdRc4TVYXP1qvJYV/DC/gYmGqPAqqlSjs4HCP4nXBEyMAlyM7OyavLV99phc
wn7EaAbMihkx/2jQXcvuKD2C7dCWg9MWQTKkYnB8Pm7md1K4rIA1W+MMLNRUiBrl
UHhJejdLYk6u/7nwWrvdsDKkTJV3zqZLbXqRMQv/0xhpkScKSD2lk1HgdEJ0k/Yi
1JL8XaDd38MON8VdNeC8txev5P/xgaLY4fgdgEA+HnHlGsGnF6sEQzUdRtajxcMr
7qwUH9uCOJOTvIcAmDBwMvXf95jh0NoLG8Bn34bdmQtnSflq3p2Io9DlAlr3Wc+7
rQy8jmr40pj/FLaftza6Ej4yWXY8YQTtio3c/+ZpAQDF9XIoAqI9Nj5iY05WjaUX
xQvwhIVenyF6mhWbKYSETA/cs4HUwKvxRC5aTP73gUb1frYw/LnoS5Q0IKRrOS0f
iPFgGZSDqfqd5WGmFVhRzfEahAHm1LRbVY+GPdYFOpB7gQYe29psotBvCvwNGzpG
8pOInz3CYpHblA+D9JPGKgK2l4MW8DOV2ag3ug5bWAzSdiRDv8fJlZ76PEQy1bnG
u5fMrQSCWwpqUAzFsPnfIMt884E105bntIr9B92KgnPRWDGq1ttfLtZrvOHl0ouz
kFz1/XugvW1HXO4y2j6M6EgNvVXVsYgZTK2wdJ5fN/ZOtfXq1SN9A5dJJmRccuI/
BkxqzYnLJEI/EqmwAO0INQVHK7Nk55GTI9eOvyCWo9qiRdKNPNBcSNPTLuvSERQH
aAWxUvvYZoNG4ozhAU7s6T38wxpPsnd76qlV8acpTdrh6qoe/x2xkdyGlBxwSA5f
v4Z8YGcTTgSef5xvqtgFXNuO4jm+TnRtdBH5SzhFqJaUP8JW2FChnNBlqDRal3Bx
BoRwI7uUvXXMSSZbw3vlAWP7XqBQFfDZobn21ZFi00PBqXtd72LLeaTpDUZW4sa/
v/uUONLnaZh8kZwfeFmO1nezQ6EuAlUe5O41PnOiF15PuCqqFMmRHRAf6nMZ1f0B
NrOugqcnqqazznWQlVa6MMvZ0G+6TNAkdpAqOT1LNbigrU5FEWOmsPEscVTVEL//
AlgLSrikinFLyfod9jQE26BZSXq5ttFExFzwvJlI7CPdnXZqLkeIY/vD4cS5prux
LbKinTnWBTgv3dLVPQ59jLi2s8AIEZ19Q7BdH6K1oNfEnGK5We3VvppYyFjCGH6J
6QnVKLv386SEuKPM7M6QAA516/BsUdYq59todL1OYjELyN3zKwwm3URj1KsnPxRr
s+wcYo7uwnNp0fnUDq7PqEzGulhXE1/El+Br0RyM5pamWdHWWs17WtvhmDDa6i3L
4QQz/vS/ObdL5XqYi9dv2mhu0+h9hUxPg1mefwarblzUT+QzGPILd1PkqdLWH6Fu
TsWJFzurqv4R3noB+XeJ5787xKGY90gT3D2w/YE8AXGOpfHEkViv47LhlnlnLwRH
Nzg51NSlgNMchULfVw6XU8fJAxr1F3fXA1Bw8Y8c6eOCR8MnGqdvP6HD7zJbMpss
JJ14T5dwriiRqls4E2+tjlex4z8Oytet6/BbNYpnRxWTv5gPCZ0MLQmUQTpKZ2R/
2VxWz+hkLSWxv55sC4gjPRt/TJo87fzX5QqF3OvRmGZWQK/3f2kNrPkjX45njcT6
Cm7dTkvopiA2AECHq+tHaBaeHS/Qbc5ts5ePh5Zf/6W5KEkFx48a5XNo8iN2Vcqo
9U+uwfcL5usY78pvgpln6Im54H97IMGlgVO53v1DH3B7OYi/1g+lxCe0CvWtA5VB
EVmYrPEXfzok11I3FzUY389SR0GmDB4F2gL6QOXwuP+DDkFa8MjFsnJFfEKz7zjD
f82PmocfeJC4/elIYZ00U0LMmV+pHG5kcwGBSqiChEYV7vEpDz5DxuQ5GpA5oCl0
cDlJudQbShzZ+UbDZc2AotpFIyTaI4UJk7ppSCm0LYxdiOicuU55jNRJRVOrzhgA
s7S8NJa3U1lBxFpsJIHjJfgfz7qWXOsMRI44N9jt0vqiFFYwBoNJsFRm03eAqlou
WD07yCOZcNfKrRBUKUzAdBsXs5NqT5867kgaf0Led1jGDgTQStIPSApy5nyo43zr
FNZUoKvT4EU3QNkJdCtPqNtGSYgDmEo1XJj4mig7QDcgaISZkBGP8FeuSCOG6rEE
8SR0jFmQKK1KyRC0z4pzGAjP0XUws/YGE/DOlj6RiNnZNOkRsFZ+3rwRV00TXYmT
7YRWcBMv3nQe4VhW/Rjiws9aBuZbJ0jpFdx0dfNwpkYM8PgWIYKh52pJhTwR3OXM
fBpmNtBfDkPgP68qejnza4cvXxfOGArLgV8hrJEsqRWGqK/ztGwe7Um6YgFrOGlG
OHeNNtXEzmqUYn+WBBbGGt++2fEYZU3wPj965XtJ0kkSsmAenJvgwvhIUmAGiW4Z
gQilpV5gvoya1ml0DhU7K8noQXvmfKfjD1cHtQLaqanOma4dW705+6bFE//CxLLn
ofSLoIi426hR3S+X8F19+236OLr4xS9hy56APyr3VjSw9xgqQuDLyxUDuPBJ4MXX
/L3IIvmhT3CixuKGspDVol4SA2ODo1oaZxcFctzfqnZcTNIbkkLSX1pcwacprznP
Nj0SFPLjUj/CSRZXkLaAnwUE/Klv6C7oFd/sPflUcy0UjV57Vl2VOHLNGc+inA1h
wngoIZT+Mt9IXwWTEE4XDsHVS2ntSesb97vCn+vKPrbElE0DVvW3tcJ/r3PxEHXp
QtALZ+/kUnaUv3iaqsOUZXF391OEODd1CtmScLzL4HrfFduowYI1TtF9iuhS6T0l
/CEAqoaRw96ROufhw8qTrjEKuOtWw8kOnqyzNe3PdPuBQCVOjoOe7JYATOtoK4Yb
93sBUL38jbsdThs2wqWPz+YjMssRcEcLsXXuKhBZh0FTBbqmpFlTcU4uA+T3Sjif
F76P33O2vWXBHOMXg+X5E18jzjyCWG+2h5Y8mevyXsMwNTrZmXKFfQD0K46aCv6c
q0L5Df1QG8ni7UebQzT7eugPjJuCrqUIFChhKjlTYgk64Z7T7gVQa9211JpMF2ak
nCOq5vjxKDDGWOEgS00T04btTwAJ6EIsqhzaMH2P6CbDo8FtcPMVn7cx+PuECvK2
iR+z0fOm5a3v0unFEJBoqMT83y/QlIHlkql8OMADoVU/piioNdHz1Vt6/8KIhcpK
EQ6LJHTG0sP2YUDHZecefVb8W3V0fo4WBt1cb9n4MC2stxmPumKnyUocOVXhdGBM
eiLC01SDmYZGtewjnWiIE1UdLSTL8+nT7YoUkkbWDAMVpcakMTsD5NfQj97LCK2t
21RpB6iqRyGlWmF+b0aHcbWnMW1C+ov1trNXfrG8OAJRs3CEPYHk/EpZWPZFb7yv
pYICn7Vw7XWY9cbNpIbPRYDdutdKfYjapy/E0VinQlVYo1GvJLcu5QbpDoTxOsns
9Fe/D7WwIQyEkvpDs9AChrOIbCab4nzKJuRV4eCq5xfYIDr8Hpk2P1ihJxBUyxVc
ijg30Wb98rILWiAKi5EHFR97ETGiZtSytbN/q8/aWjjf7piiVWW82mnOm7d0NtQA
IYEsrx+f50KqCBJpDCXQsorhuHoQNBtV1ExFkpJH/FQV9ufWos9uE0IjbYxw1FAg
qVyVFj6v9eTvpo1cgCsuSCkmTEbmKg5WfBuT8SUSMb5Wxw9uS8plHfBuIAEdUu40
u8JGP/fFJIBnsxl/QlRVqC9gfR3VtVhTgn+Rs7M9hrB9hprc/tgw51D2onA8UR7r
U5vdyJdktwkQ0idr82aG1c7VhbWS2vUWEqMx/BUWnftfemip1c1Eg5Qb1d7MZzIz
PauiDSNFcigRu6jzF6s+GEfBg3aTjO0LAQ+099R9Ct7jpAzWM9uevgaLvhzrJQcO
pHIQ4ytIHR1tD9FsZQ2Asdtin/LR/a6q2lDXpPg2Skzd4fMa2DZz5brbZiDwmeUi
LU3wrNvTHno1o2TjqDwb2L/3kHZumxIoEU+bkysGxEWkaqRA2NOO92ZyEnGP4STr
5eaxqeZV6Ycgnidvf1rBf3CbfFvat7wA5y1wJnaYB3Vj5HLCHq0/U0RkyFOOCCJM
HmvKzSOD+ALjFx7Cgp8IOAx1jJetVmzTXZ08IeV/snfL4dylusRj3RR5cnIGVFTm
LCD67rHYt16RIndU64md6hFj1pIcSGVCUTMVThfZkVmJlpgCvbQ2f1IPBSbm7zvm
+LRGc7YIr9cUWphkbNkvCukcc62ab/3jYNLse/9psbpO+ST+jlSqkhyScY8pAlOi
CClf5aEDKZ5cxwvH/9vNznnN/PNayu3o8DW+BOK/vfwTy0LAk0fn0DN0NEaWOdnd
1hjGahz4NhN7VBpcPRVGTWMc2I5Xq1VpBOqdpimbjPqBl/88PJPsNbw0lteaZrme
4VwzNjTts+nEJbjlIf5r+1mXfgJB7lmUIilSsYfZN4AuXVfYGLvj9iaXYvIr4K+Y
mtq4m4Olm9aalJF7HBLHdha6iwD1PpkliONcSHpdpM8IRhh3HSqECgxC4FB+LGq/
TpkczYWZLAmAJBfyWyshQvIwAAI85FLT07gE2TTmZELqzVZ7qtHhmmsoZNKUo9GV
m5XiXIU4urUIAAGLDtO50LnqskuKahovhQm1UEVbQOL2jhsS0DS1hXT02glSvvHr
3Jyw5cESfLmlYq42yuxRSddmX3v/cxeuH8qsPwCeQIQnGWEPmUYUmGYiQ5KZFfKe
5btK+qO4Wo5p5Irxwn9pxhSmJY0dvZaaG8Z6ytimLxmxUNGGQgf3ESxqxxSk0AH0
LsS3pRV2J7GOUYULWznW4LtkBTS2u0cNhQT/JBldZrBzXgMn52BDjPiZ+Kzl/b8C
5Vgqe4Y7ihNfFlnIWKF69komXWjReZYdHFeSgGgOnBJjkMzWeakEjXQnBKZGUEUF
K13WlG9cg8dbfXJxPWeo9Wd1XaA6NyMskW5zpPnlxYm/+TdYjbpX9+GPQid0MU7e
LfRPIMMf13AmNUuh6A1cDA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bUTbupVBUqennX0WMfjEvQyDIUGQ2N+8MR9Nyf/jpLj9dWZ+NDhvrAd+WlsczWjd
hCs/guZMsZfGF//ho8RZ4YEqVpCJ8SZq4pxz4bydvE1ikYtIRT3QvCcj/GoGqHgd
I8Tt3CiIlR5Aa4SfZ179a3uHnz+MpOzXQjqEM+Zw+ktzg4rVMCoxwhf4ECPIepRx
AgH3Vh2FvIRQI5AfmZxU86PoYXK9lnpNXrJOJul5Lhg0XoH/6Jo44wDt0nmPFl8B
HhdgsfaIvFFXj7bPwOnYcjKbzWuGhQhMx2yGYldIeodkqDEeHXzQICf9aSR7TnhQ
OqYL81C4RCF26W1o9pxCZQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4928 )
`pragma protect data_block
CUSLJ32aq4+doFDpy2cGxl7s+Nnmx1u8pdlmuTHp9FPoem07o1EM4b/nAxFuxoBY
6ojsyAr/iIyLANR6FJ27pXKNbBDanauNTZzmraSpNV8qe0lbfeOfdiGwBUle66jX
93c0+dVJtRAniz7rV3u3KhOywmL6F3FQiU8OtcLeuc/MowvM95Kjw3SgmqgRBPYc
gEtD0Up/+R8lrrGef2HhmBkl4IiV6hYomfq/ydlqAtpX4XdLGjvdn6vUCAnMih8w
ehUeFCBFvwea+WHXHMfHwtI5j+51aH3lvkjLU5ERz7Yfuhldj+JiIJHe7SqJakSQ
FtGAjN9PWTWww5T33IxFAhb8xO4dHUDL9wTdH77ofu5QP+hzotMzw2QBjLxiUg8P
n2OEzwfbpXuyHtMNM7XqfDhcguvxirkvWw1KECWknJ110ZHtOnOs0qggBDHZMaZk
XJMJxYAQf2oLvKVbbVkb7INYQcaDyUGwbsGWq5G8ZzLH1US5j1mb9nwaDe4EmTQx
Y6rEtG4hWhR+YLaFVWMPW9PqLJPqnuBOUGt+oE1sAf2M8VDTozFO5HXoWRYDmvKS
Ouz9ZU/Xeu1L06bKsT0hD0eHwoFPgjMyhThsj+1eTH/aqhgGieq5luyTQqmCzZ/S
9VJA9RrNUT6vq5Eo86re2WACb30yBogiCYjDW0Zck/335YUATtlFsd906dE+1yt4
DMS30iKs33FZSNjKLGZl0/f8I5PXlKAcYt7hCxk3d5eSr1zxHGUrGMCmNfCoyREb
ds7I7nrHcxNmzacgmHugjdcp6m4dM0K+BY21pVAW12oyOb7gm3WNQ7T85fhMUtuK
/vxNM3wwqtrEGJdN9MvO2paLqAdYdZ3SGKzyn9XFnVoEjb8n1JXYJCp/cj/tULR/
4uVVqpznVuV9yWAPsJrI6f5yt2e8giTWTHRzk7wt1/F9tVKbCbRi3qae7Q4L8opd
f73o3Lpn+ILGk9c7LCt3uGwg/jdhgyattgQPOflQlDPEbHveb8QqBaVaZIh8cBy1
EUjYMXD9YX23psc1oC/cBmY1aJ5Dq1eXQAmTH3IsjISHqPG+YCkf/xu1Vr1lwIcl
0YOQwmUrYbfBD62NaFCcd6fdIi9tOBK6AOEtcXftYrGzW+s191AXaGv7KWLafEu2
OhkK9hovKFm3vRAJi8zSfV3Ktufkk8mUyBLDsvCw5T/JEP1f+VGH4NlRlaiQydSq
aMgoccl8Vvw1ftn2ztBDyCxV1e1d6OZL47mnanicOHtvncmtmlgAfTcHh0j0xSWJ
4STV4vnsLPs9uiKMcSX/R8xGE7toU9QWkckl2+gTzKz6ulyrRNA6C63UFJ4deRF+
0GEG3ZWvidN4u7mkvyoz5q6uH5fRtF0mMnbT6DjkA0+WzopkZGhRiO5pRae7NPEc
z2QrYmyphnbq83/J6l8OFGUa+s1TLkypsV2SvhM9LXuU7TVuQLVGpJ5Qe71z0DXN
WsHRBdGeh1nuyMdfyEHaDmZX/0iV4b/k0AEjWnvz3qouJulYY2xI1F469L1D2Jyc
ZOP+s9edAHIV/2TIMdDLyGBbU+kn2S3oHRA9WteAlnm60Nrku21K3CMIaY6MnHg7
mMp3JFk3ZeQ2sMG5flVwLc6ZX31YvDSmluHyabyCjLxe/+hz/S6Zm3VB7nFDRjXN
tw0JKR4/oyFj7D/KPwRlIEemma2RrGHpM5B5LC679m6GICVODLLBCmI8ZWpKfaBu
I6NWnHuhp3F/3bUUyoSWxe1n3HVQDVSs20EzJ5oxsqJgkHVL9A+Ab0yIuzoGmzlv
ag/tOKIoCN+wDD/zVUlMnhuVqz/7QB2bR7jxg7W31oZ4cAncrmduiywD1doDBpov
o/ZjOJJiduvpLq5MgdvYCh+bera2uAYQNu2GDmdKgNXt31tpOq6aeC21ETktm8e3
yQMH4jGJ2vsyn8/AB+Bl97s+yR0rT/S9U4QLbigVpWFvlNb36MZdydtg/ZGQc2M9
eyHniuxXutS7odVLl4NoIrjnnB2oTtX0+/OjysPGJ+rs7dQVA5CLk+1NPzPmzYjN
nCWYQopmlpZm1mCmJDnWJKXJwNhgb9/Zt9eZGCnwn8MBFHDc8Oucd73HYmmM9J4k
MzSbD6PfoXMKEaK2kIhH+VFdIwj754/rlh6yszMU84M0DkS00wmafGklEsEz8ghc
25FPCEekVWJ4Lm5czKrWMAkTpPcpplSzXOU1vAb1pvhrO+XF+kKg75IBLHCEf5hv
bTfOp8OZo/lioEBRr5j/MVbhfAMMrrnYF3g+z2+bXKzIJ5mYPYzteMxCUw10bOby
wbcVN3Jj+juX643adkR4xlwQSLu/+OOL8Ghkklie270wXw6kIc4qvfhSZgOHAWVX
5lZTwZBrVOSvRUkfBBWe8M2Yx33d2uKSf93Hd1Nogjoqpp541E9aDT1NphT2wJUq
BD2GQJnVlpb44QZtiI3R/yhxJjo49oGsrLEdcvuXaEz5SurYCzTss8loI0GIbllJ
RsSqltzQ+UKgYjshFlgBhlv6dvfgWZj/v6Hp5DDTOdGhXBNEf5BIWFFg+rnvHlSF
8LkYVsRXxozC1Bx7udMqTzCzf1zT5ujOwYYsuQnvEFY1aTsannKSXE8wDkTYOk5i
iS2I+Fo7G8lUvjcvJuJHYPv/OIG5YqSS8XqZrWXqDqlHTzEwLUJcsc6zl+zJCDAt
MC6rOKJn9bwRJqL9kGdmpKsvSjWbdIOqD7AUBdDaSeohrVI/xOl6R1mC+PaGqlnx
wIaLUdNSu1BsttXaxWRai+qqG3bIQ4OFL7+LNw6NkgYWtSjVxO2BQutuodKGfRJ6
ozZW7dECbWcg5mjdWhkjfrbywbwzDbxLLj8LsqZAPgTwKn4lyGEm96IMWcSIqMWC
ushOh2rJ3NyIXf3KyJ49U/vtlYwFV2otTeu0u1P4LWWioUU8H6xjPFD1Pfgt4V+Y
MhgSIOGJ/O5B/N1CStBqUOi2t9K+eDGd47oQd4kxYdvC119LQ64ZGFbtX+30a+8Z
S+MTPnc1S/fBBBkoW+BVRn4u4GmGqnLwuKtYtauu9+q6poRw0xYZJLfLGDEa7Qkp
1/YUCoBWQ3urpfyMYKw+X2Q8iGyEwMxPwxOJkhzIDqys1Ht++vEHrK1h+7Fdgg5E
MziuopTilg7IG1THVdwOld2SvR6k+EyNmVRs8nDhxKkXIw7JHGVQBUReXtbthI+3
RVApux3R+dlIL9C1QImN9FABchB6iWQQVtHpIMQRmjHYhYzuLH9w3PNOq56aXnrf
SV4S/6B70FreUV7qdAjteHSsreNTd67PsDQMw5pWwuofAteDAN/jCluOO/m1CLVK
IVdX9DEW2/UKP7+bk2mbZ0qkGRl7+IPxNB9RCwTBOAtflbDbGUu9cksVLDQIBzoO
eJyB0BkTqBZFii9FNSQkVIeWFktEq8w5WVoSLM8mePs3gTJY4qWJGAuspSUILhVt
IgHd3fRr2J1wea062AwbgU1ywbsKM9ZHD5deLO8VuykXf7l2OjNj+/qSU3kxmokV
wra16o6y3gWmFE569MAVTNZbYckx8kSY8Xvq16Bw83gkh8gUpmnecOY4SmZiTE0r
19JpfI5md+A8Z75GvHKreAsJ821BnoHwo9RKX+s0ijrw6kJopxggyrAAg1v6ExAN
oodfRLFYk3I9Gore+/yY+c+7I3BnnH3y/H6+4oe0puzyjwA7T6vRQmgCCZTAUUMf
mYWZf+aH8dYiwBaaukhnXhvJOT+Lp2yUWhA5dFBin5Sav6VX5GAEa6O2kP2xuQge
fq6jz5/FZfcq9N+tP6+8I777HFGxE3Z6/j1MGIAAY9Qc8wBCi0wLJ7T0KsBH5OOt
+gn62Dtf1+mFRWcq/ITVvk09BHHz1EpfBMbEBB5Y8B2sgS2rCRCW4JVKhJ00j8Yd
52fA3jbAB5bvEEQYjEC/h0NhqlEqaITIaC0rXmu3wOVqpOreQgykbz5jxXg4fwEO
JQDGxZedsBU9legW1m/jrMhOJcUxbu7caZO97BJym57qv0J/ZP/6hdG9PKLbc8r7
KBFcWlRTgaT/Ujjl3FHhLXcWX7Zp1oEj4xhJ3MDPUuOH3dxCo6n15ZROon7bqmc7
X7fn61y2dJ5iQZEPw1+5O5e8JCjEinRZ6JdYVKVBDRyGdHry+NO/luuLLoM3aQTK
hndqd+/b5DK+I72W6zDvRzRDUKJ/cM1krlkAV1HQ9NBcM96qT45QavRxCWmiQ4cD
ah8N8mATxLBCfseJ08RRCYcGkJy0dX3fvuvfyQxYThnwJHCpvZTM3FijOHVsQ29y
UuiXiQQrGJE+Q5URoGh6MyDqv7Oj4i+VFQjc5g3Mt4S0yXi8kE+3SPCHb7Q9QCT9
fbR8mzuTJ4UtIppzFwymqJbDN1qXdYYPhoh0Qy/aMY3zlHZTTQDm45yZJlLE/Vzf
lprjR4tmNIqV+hqdHSvlCWKqWCn98vTWVPEwnrGgWKaJTBGbwQb8zKEVuPFDvRKa
E5J7oYxuWAORzGvV+/IVk4f4eOWupuCyrQi9yeWzZGur9EA3JaH1GdIBl88+0d15
libC6uc+R9+DkixXczNLC01rAjORbAgbMDkSlUMmknQ6IMlZ9rOmwNQV2qzJefRO
c0M89CRl2TEOOu6LqOvzlzCLkCAx9+VluNcwHCiJP3DqhvvEzVzqrlZmOmq85K/f
cPIxzQgJNQGxwx0u15bBe9OZjjxNWO07APhCCavVWzCUD6QDqqNC+qqdUuNdBqPO
q6n9BoPU8T6bVABoLtJwtK0AUelJ0QgzGZ+jn8+V+Gq5fHmMc+ym0t3tK+pXUZJF
KLhyV+NIschTJW4/XxlbPspJq9fS1a01+e7ZPJEl+2Iy8zRKIRtXjU0umPOPESOo
M0PmaUO0HYJqIgNsqY7AVw4A3Tq+tAud8bVg/e7BTX/kmBcJef6iuhsLiHSYnl87
IB830ng1iV/fZtE8MNGdr9Y4Er21l85ucG763sjWxnNwkrXL2fLOXcbV7MbLl2A0
xKKHghZ15lDqX9+udCarficJShPySf9FdFCH4MgbUZJonDZ2kySjflCUyc+n2mHY
8WiYSs75aZ6ozq4Q4yymV01BAjlOjxZTMY/i9Pd/Xlf2blqyX51EZYzrv3sdXcL7
HDF9Pd3+Md68yMZ/eyFXxzksLTkh6tNaxPk6LUOZYOWLg/Sg7yEzlMKp/55MlQ6c
x16JbMnky6Ef89p9BmQI0g466Z5KC+52uC83ARzJw0ygKPJ6qXcFq2ZcaiQaFx4j
SjbOMXbNGPBE/r5t4wP9jBKdywu/oDUhHgSrbUINtUWIWDCbqo6qC1nVsIDRnVn2
8IuiItjWayhdBwbl9qSEcsO7PgqlgKVIWzo2TsUjAu+9PHzJKqyRBIYPxUbYmY4g
GGac/7bulSPwwbvwRSL/unb+iL/nMGxh49mSzJXIC8vjRZfUgdmoyHWfpjYsnc5H
mvrB8/XVulcXU+zA61bZwVdkH9jQfP/OFV+WuoDEi5oWf0uLZKYInIqeN7Dk/8cF
Oi8Vadl3PlE3c9uIdr0WATYNU9T6AXoDILaoZzAhs/saEZ4bdeieddme/MwdtmeN
EeAYZxkgeFr4IQOEBK4w7c0rzwcwJdfZApTuGFX2h6kM0gfF3ujhOZpxvpSWuuZN
A4760NUkwID0uE1A9WvQHfXg/KYV4ila/q7wKmrO60l/TIHMLPZM0K4lJeFzbKIs
MioDslmF1huKb7ALMyKbF4lfbxFcgeBAhBHKKWOvyoSfIPUOJwrhZDTi7224a1G6
J7d9v6JrAP8Lzb1UZD64ExbXB4Pmnlvwv0lWf3CeuOTuwxtNskGf4lx9b1ortkEZ
xfrERN9G5ltk3Quni3Ed+BcnWucmevLtfyjR1MbbI3jI7cs/3C9W2KL/yAbdqLJx
ytpRGfgwDfZxhtv47xErBS97IKdSFXM477Izf1Su8sv9mNM18V2QUgtpgsXXaZTP
L+k2OYeNOLuznUElqxBhG8Fpt7B1XLl1daxHoIQCRTjVFMCQ4RR7z845+oVO6HMg
Mrk3/cpW30KgQ7sZi6MbMdSNe3CVEs60meVGvJw5Uha63+2LGRZBKjdjsInKkTO4
uo8VvPPnlm8CVvkwU9B8QkacVhkKDJPYPzHrDO/+DS8ahuMLfjJE5vQdrvhpNioW
M71DxsluX49ufVqODdrpsyseOwEAA6flW9v10TuQAe5KVTrOlNuEjd8eXsUUfwjC
UICeHrlVlCmsSl63+/+4bKwOPqD5L3Ksm7DlguC++aQFrkUC70oGWcmUzlFjLcb8
7FmtTYvNQ/z2gDBRooQEh3+2wmv2307OKzLnHkIH+BLOY6WG+cqm8RWDfGwjHESD
cBU5eKi9OfRAVf9J4vM5hRKC/dD/w1pAY3ixMZY/PMpqfMRKWjgNjFYHXu5MOYHL
WePf6w3HnQf9qKoG2pWT83u098R9jJ2D6MHgvDJum6D0zhcqBvhcI5GEnTW/GU2Q
mwb+qWWTD8gufoZeis+wP9kDiDEY2B940FuouWwXBm9cfv2DRW0eiTK/Me4SRWk1
y9FDJnZQOcZrosGimu5c9B0VTpEdpEV8/1VL07e7oOE=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BqI4khWhqKTqjfFge3oTDtvj2dLAfYoQz3WtrmwOmD8DmT6FdttilHj3trxCFcRx
HPxLCZRqSGQbXXAD4DjAqnxrPTpRNV7XQ+kLtUanrLdMmiulU598sCAcojXWm0Le
CuxQCWeogwF+UUxfv/EjkZGG8T1jTF37tGy0VfiOMTeFTc6vHGdD+jnss7s1lV9H
+XEi14LF/AQ2t2Ka+Xu84XIV+spDR57SUPeTjOI9gRiaGz7bTAj1+SSozosdzVyl
8WooEHcNv8hLfn8p3PZ5Eh5JWjCVuhoBVp0jufNcF89kCKPbaAb0iFKXGwInG4BY
o3WW0mD9RZiFKWLwiTnLWA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9792 )
`pragma protect data_block
AbmCSmQYziWiI9ENCq8W32SgCKFLfjPKkBfSl4dMVnBtrYojxoZepmrE0+leMns0
Hsa+n415krg14V7EpEaxQjyrvKy4J6JUp24VYywy9UTodvxU/b319finpK7FQlve
PYYGHepc4khqWEQz5SFDr5/qM2mgNfi94aJuxy61ZutdZfBvJN5qQkpBl0b4DEhe
WPSzZZhXVMlhfGus/a/oJ//5a5sRCXGwQrvajcwd1SpypmI6ak9DddToNOiP5Wih
oHvdMjsi12D0ZbcDVPPi5Tu8sjLm9xSdTfZopWP+p8zKa4aqYmBYyS+DVd4Vre18
TEdxxEh1sNdhTj4D5QV+4pt40Ibsya6mal8imADIQCaEUVVOuZv3ZxDFVLDSrnVw
FSmbyKBXHXCnftmDBgboldm/3tb+fttoNaCQg+Iwj3nEq8Je5NDQ2hALC2Cce4Jo
XhdjQuisBFkRHavdiI/rCmNW84XCYSXP7wr/58JpRhrGgRt8PfjD2X/M68r3o8Dd
t00fChVRHXNZEbl/Vls7TedkfCASNxLJdYRkYwS5O+b4wA7dfu8EYjYAQWlgW1/j
TG9UwSKFLMgSFhP9Ww/2siQRvtb+iwPywGhKa4MyyVxs59AtMw0UoevjiHpu4DVo
VT121I9EQ8nSWJDxaXUUuz8OkoCNH2xSLpPXPU6CuMW6q+bJ5xfVbB69sShaR99e
ag+5FcAMyusdRNOoHuWCEmnisN9JHukvWeBm/O7bXLFsGCeR6rBmUsHPZVR9WQBs
BqDye6dCIBmIpIDouN2LKkI6TiIb/9fESl2JsmUJ7qTeQ68BKB9fLKsqC2wcTTa5
WfwT5bFacb0o7YtBmtOD5ST8hbHxlO5jsKZc0UmiI9XlvaGeSX90ib5R0XRfaCT5
zflKFHxCT/7OZYaZhZIYA9eS7Nsjvh0kNhH/rieOviGhfiOGWsvvNuHIkZe7bTtO
QfJ0HU0HaWrHactRWsFhN22EcVWaq/swHOVwcNhvrm1eezcqFCS/R0qyHLRRBzH5
5ALWIQUwPEsY5lMD7z6O5HeiRRX62tRFCBJcNDQ8i4JtCruqKOlfqwnciAVaIoks
URV6acKenSCoG50kJacYkxKhhNuV3Bv9cvW18b9nu+OatYO3uCJYMBBUMpaayKqz
JegVYU96ZgTWezWCG13IBxinLCBOIxJn37/SNHGNDBj89IELWtgB+svjs0H+WUrE
snh1DE3tLhQttI7y2dK5hjAbJ5m4nwQgUTJPuQVhhPYOR39+beeNC1O31tj4Pfpz
0K2fyzwwY9UEspP6iNfZQKw9VnbzteoIkJ2DtHIU1nndtjVhWdwqjPjfYa1FOUuc
ABrDOJLDFztvkwo2TJYQ81rILMtrVa+IVmJKyQ9CtKvDONbrcrnrgiIBTNQOxXjH
FJ1NGStwLGpkK2Tn9yFywPSKByfjt1CZJ5IM0UGizL7ajKFrOEoyFh6PSLqldRh+
kp6orez1NPVlu/6uk5l1h0d/m4GEOTIEOWlmgL4vB47/UIklkFYNdAmGsf4T5syF
uEGi+V6lrE/PDkey7wIMrTQ2esRqYxphjq5eGd3HyYl6asABvo6Y0BLOXybB82jR
l0B9JyJGiYg4leeUyOTllhwlDa2QYPyUx53klYpFfNMwTT2w5v/V5PjD6013igIg
RoKDNzPmiaMBNWjZEDOjfjzzC0VDQrZTAGcxsKpv7zvR5O7uI1G9IbG4LoCJ7uMn
KM7i1cuq8Htz1TxG09RGnNCv/DWAo2kEzeYLFz7oQMiZWZEMhY7lkTtn1uuDSZ+A
mEZsyK1nFdzSN7O3crYXSwK+nj6BxRfDIxC0uowxOGRQ0/W0gyS9+u/ijQ/tSClq
bIxvhaCIFxtWbITlUIjngPKDvfTl2nvhQqaLyLOCrcBI1eDUvfU49LkM7JdgUaoJ
dg2FbAfHkdBBe6B19jt6L6EkKQ2F8FyZCrRFbINyG2cPRDL6L/2TuBiOORAsRP2Y
mpQaa4gVjBHQOuwdS4rlx0B0Pow+8oJh2NitoKmyFgVUFGabw9WeizrlBrS4ZfF5
yC2FkQwkXgMYpqIbP6C3kPICYwITX5J288Dl6B6BZHeO3C09uo1394Mi71upaEzi
aPa8GZirLbu+5SZg+O2s+0YvMKReFAKckX/ucsnLe+GomOfAWglQsFIzUOgrdxrS
Tj5sETQSjswIeMD/wWip64kolYVV/8l4qqfExY/4gYlKiZxn3KooSAwlltWR1ZBP
6sh3op/MWPrDuhmHeKD3/wFJlnhhldPAHHP3jVcLTs1Qdmhm/rucQiFsWPrzNqDT
EktZ9eb5l5RQZ4wR+p0cmP9Fb9yevB23238MvUXKjx1PvsC6ILuhKnwIVrU4WBgf
j/qyFleXNRdv4D5JaYmHv4iDRfXmk9telBT0AaHENL8YpvRbHKGn9ff2GQHstZMs
dbZO7q01nxe0YTZ0Orfyfs4oap0I8ZuKIdAV7ZjnZ3xjdoP3ONLtL+u5U3mB6U4Y
urR/VLQCL1/vq6qMfE0DrfvQeDQoypPulJz2LWdOsd1s3NWaeBDoYW19WJm6IWGN
vOlgYQAnPURkQYfwPf9hgQFDn07azBRbEcG6unMJ00gHC8H9bzS5eXdBsu/yFWbn
TB8giwv2WekRExnXSRjPpEl92PaCh3eqD+gGhtGBwQr//JepM/csxU9jkbWa3dqM
65BFCJFUnXQ6BKJOSeYHjz1hSW5j+2SmArtWjcdxV0kRUYT0io/FFlVpR1Gy/kZg
M5tBPUKybPHkdT3Qyy+TB+O1uxRLIWlqotV42rmxT/PdtNR80QiiQYnyP2Ok5PNA
UXa91IKMkvtQ/mI8A93cvAV1dTLhPCLKHy7sPHO100hJZgFKsBd+1Q5UwDC6iehD
5BeXUAfa/+2f2wKUXKzKrOZvuKogILpwzKhqbjDhjQfZpzisAyo0J/z5aJOSveXe
H76UAK0VsIjHF7evIKOd82PMARirO7jtdfZMnafwfonwOamRA+zM27HMOPO3lT1g
UJWivUC6TsAlpZIm5v9FNHC1lT8jfDLNfe7NuSFmNQDTOkvVfSy73jeSDBjfS6JO
xaNvFcAkL5wzvgowl+2ImjrZ4B4gz0yUS4TDVA+GDnMGzuzAv3rQg24qS0LDYWF4
38MOjsg/e7pxcCJcduPQ/Sb5nGdNhgk8Umzb/co2D9eAWj2VKEgEx1HvK+Hp3Ao+
KKXoSbGmtbO38qiaVIE+a4gXBH5HAL/IhBR8K/sZLkazyGIc6CKdLQalzut9Qt8W
BorrjCh9dfelX2VVElcb3zr0GexnQ/PAA9cW199Q4fS8+/46zzVR2/YridSPvuq5
CPqM4wdLahMW+y/KmT24cYrCOkUsZalH8zYWYNnpvnxJ+hkhSvqrrrxJR43g83b7
Td8wkcBwY4mhj8ZgpCk/TplBxpldeB47x5/xLFQTM5RroqCUskq7bKBvvX3kawhF
voW9EtY9OCddzOVtghsdNEAmwpmhMZclyOT435QHbVge/V7PjJ9lV8D1G8uQeF+W
dnOC7NL0kGf+SIAwVYp4EaEnhHgVfSVgRJ6QoYOKyPNUjT0mavn2hGD5D7VUVV6r
8CkOrLI8MYoa4mnuDONXADPs2w7CdWaHhVl7P5FS91oSP1KKdk0eWGsoYRWGJgiF
9qWlYajTzNXP12L5Kk652vCXNJyy6ZzGEBBUkxRWoXrAlWT+m79WmHJ9fO44d+fY
gLatl8TlqtY+2I2Lj4Ppz2jIvq5w5ERqm+p4+7GFzCDwb3OoPXqp8t8X76S4GQvH
hU8cXQuES74fSIV/lpGg7cmxZw2SXje46G7hlsGLVfMDf+PgZwxqUR1k/808a7Vy
IGkEpBNFKmhidq8lL9w/kzI9SFyzwZ/HRTmySTVk2w7LBySLnNBIrbhcKDiKanhj
/yBgyANRX/y3fhbH6O+0FmZOQb7VLnAfwHamjYKixvgFPleAYt5YorWLU26lpxTL
iqkEEiH3OXM/9F9dVKTv9/Lk88LPSy6v2ATYkPTnz4GRDld7C01dqKez7ZpnwNKE
Yrz1IoG+4gSL7cI+PU5qBeTmv3F/h2F1dqiedY1QTDHqhNjwUMSb90UO5N0tDqam
IWG5FcpBQrts3+BY95Gb9QCzg+Kb4NhFg0aAihV7tB3F3iwb1m4skU1eruGaRPEp
QusTqQyakAYaMpZ4I/YMMRGvb2tTca/CQJHlSHrXGCkjOXyAxledRSg1iBMFhE28
jMrIwkBiugz86bdV6/bC8Cxf8cIPbUDMxMWyBnRyPTA4P8SuoD4lHtDz21wzr34t
cEXBdYVczRPlJj20TVzOPKZp3vGbNzBZ3vA/WVXB57x46h6hib5sMT7FrNtH+3f0
57G4Zy3on3CEI7jRBz2g2d2ArwssC4aNg4uVQpTeGKbBNq4iD9RjyKxWEE2rUgAV
WscTDDlspN8lGiphFucnSKV3wtdkLu83lqR9WxP6ZbLUF09h+FeLG+HplqGOR3La
Smqb8shaBfnNVGoqvA/HGCINL5CAM1myKRZgtPbrhsaoWO8b3G2moOAxBrjCQBLV
MEsAGlytuKBm95oV3fLhrFEfqTORwfxFWVk5U/dqoK6rxo3s0oEiMQPt9gZ2pDsq
jNLsrVK5xKotI7FVBXa3BzkpSVVmDlnvDXEtKQkCbTLQXJ16EzXuXsvQJlU8zvv8
DEAckZNelTz1k7hh7R5cafhKqr6Os7X4zxFwR1wLYJ0RdrQZUApdxSP74YlOja9T
V0xSej3CGeddNoRwm4/SxT36lGmIkFMBZHQP3nBEZUhLw5EqYRpQeYIqkBcX7Hs3
KAzj8PgJa7cqhGxfqxFaye98Vxkc1SDvRVmZ5rli/UGtXqzw1FrnGRoyEkuhC6iv
5iQmb7VcIHn2eaWIvw/Sp0XYW29u0LbfenXSIUcD9cSU8hxbfPB1CAn+lOEZae4z
pSzOojKnHyPalSyq5FOZtrOZRdzKvC0WfJ0XnF35AcKxeMdegG2CTFTs0kg1pcoH
htLTyupSUIH6ofujY6uZ13RRsrRfpJCAUIhY6ZjzFIv8yid5v2CcmU9N0SovgBj/
PsJd4/sXqcwhwDH6c7ApOARWf2Sz2f49hWMpei1nRx2va1bHPPTf3Zk3SqKmKnJT
jnoPopKu8AZnwX7ugqy32J/3i/QLHO8da4oiDjdWoP8eTjld80uUGUUB/d5O8Fsk
wy3LsEhwFp6krIb+jVvNN3iov6umOei9bNCNmN4agLPWfzJ6pEo5saHJBnYNvenY
7CPgoRs57G4/Ba4Du7Qre4szTPZ8ttF187fU6COF5/Xzd8N700uzBEQUbOGg1Vzv
dGAMlMzzDVj16vtTNQW+aLTCw7CU63g43mfyvLDNUk3LLpWBVR4R3ZACGkziaqIT
0W/8dwRDTPCSjAMUCuNlRW48LV7j3+1RBha1CUcJG52Mzv6oIH/SFaz26RoVACyR
8FBZ3yvU9IAhwPJZ/GlsA7o09Ulw1detANlSEuoETW7rPrt6UBOJ8Lmx+/J8kdkY
AY3yyRAtuWv+eEQ+uj5uNlsrw8FdDK1Ryx5luB45cACXI5qQgbdIlycE+tsTqgUR
B6FCt3Chey6Givf3UxyXE/W4dXujM/xJyHvPRPA+uSVMZ0HMZ8P64bg1COqSNTEH
+Rvh1YSppxKpU2gOAdOTHkd4RvbV5IBWTzEnn6P7GrhXWRpmSlTaNIgMjhHxBkF7
Pv9mYzrnmTHMtVWWMIdtEW3JDr8LnhlMxEE7MJkmTiD19mYXnvcLMfNO5dXeD5zT
MdQ754xjrVL7eS8EqYXTVSRkPMpfEZkKmBrsXzpOg8BLIgWXA9WvlI9Iqkhclvbv
nUkeC8hAvau/8X6ocLYu3PVt2e1p+jzFWDiCfeiwa3+4nUGXmBZIyB6X/8nU9jOe
Lr9ZC2Qr0iBuPZ8ylVw5h8/R/gXNaxuqhGxNyBJsQqiEl4f/nhwsHWNJYEIkW/9A
9rM2l+K8jcm77SE08vMSP+m2jLdY7EENFSffUlFdLBYl+NSJkK4sjcAyf9cnwY6q
4jY90R/k0mbtZBBlb+7Z8qWL9S0BJ/3tEg0R2qeLJ0vP9/k0xLnibCZdwz0FZ5W6
iedVjHX2ylOBDdj26mWupFerjg8qPwX8OCGxgadT9Q5o9TqFkyX/2FIm9wQEAYiv
R/6xtN9yCGVQu7LOGTt3fEqS/E+ICAuha21xAGefjn0n9Y4DWVj02qycHpb+rMni
Jg407BsOh2/Q4yKzG2cajeh6EK4vEqK7b90QrDY93ev4wHoCNgPOSs9EqGjTQNUW
0t9b8Cx4v8O9woHQ8eifidwb8X5PnONTyGby18WSd9Y1gUxnLvqrNWVMMrbZJIvt
riGIm1uuY+UsbdSVGVtELQ3GSXf8phxCLmkxpPkCXSVZlxxZ9AUN8EdiVfIpqiNQ
zjH/gZQOe9mvT1OgEwqdCbuJO5AGA+m/xuv44ecd9H/b6XHpn1AEXkO6BRLP8M5C
AgwBKT+0moqJi0FM6qE01N5qfqZImAwtiZjuQ6Jhbc3ExeaqaN78X1u/FVEt4kD0
Hvl26lI6780Y4sAJTSsaUqL8OTm0gQbzIqUXebxkohUfR2+wxRy99niMGvWw8zt3
GS4XZvyNz99ibt/4aN06sAEkeEDWeHYawnRHDFrLWFcXHYkSYfSFgAbsbr2n3g0m
mKZYBHTkMTwcRHFyoxLsepI4keOypPKwapt6ap2YGoORSsvpnkLaTSMZYtw4WwWb
AwEFMZNJo0jUaJJcdIHn4zKGq8Ykm6QQRbcLyIsHsn9T72vnbpLN7tAqWkKNtZ7k
5vbKbctp/Pr7WmBWCYNFkQA35PHFjiYrb7MHd4hcB9bzRf0/IsjsnAe4Ce9M2zBn
aVrQkbi0LhHBq5cgip45BR42pxPNk2LSqfAWmxGlOoT48du8PzukC0RC4Ccq9uQF
1+vUZKZVR9Inu3VB3X1pSdoVRBz22N0FBasUFLkc5Og8Kri8hT0fFDioebyt43xq
Ad/0VSG5akCJl6La+0AnJq1H0G+iHs533A41t4lt0BHiFcXVoM0WcCheUyk2MZHM
31USWB0YrZZ6zVEXt7uKhgIl2dxkpyTr5/EcIBQLMBhAop5Fe3qzT66uQNPumyej
Llg2da92C0+xJkv0N+ZTimJjVtv68cmpSasTUA/kFwOmxvNqAd2j3OGOcBRo+gaT
9TZJZuCJl7cH6JwRmTsiZ69ClI7BF7CfrOxn6qjtHh3RprpSiB3e05lAfiAYpanI
/X5lRgxgF06q4SBAWontnU5o7e681gXctENP6gnBip08xRAdw7QGN5bgsxbkKeWr
mrXBho5SG5wnlkMU9d6xgKDI3Kh4eLEuQM1xJkopOxCzdpKQRXfGt35xz7UiklCU
TzoylYhGDgduvQcb7n7ZS8cv/o7lGAGLGf8Zhw0Exoaz2t+Ykusspf2zwVRQsqn2
DPxPQ3qa9zM/oMwbHNAzWumx6dTH1TxTrJgJO90ReRCN0cFAwVSsBpPEo3PtnJZL
YRE+W21umGb5OxfHC/1eQE7Q7kqpW2cjHIgL2onZrHooeuR0DyaJ/wHmrl13XOZZ
hS1ogFkoyeVmkviON2NNOIa3ttTB5QbI/JYydEk3QaLpLlHBG5g0L9BJbWuS7YpE
nKKsTMarUlgleUYsTytGYMfFoAiuITtazBEg+Hg1m2a4X8BMdxABbgfnxitA9VmE
velfrtlCcKzcpmiiW7POsjvvqxONH0CdpFqpqKX2vlz1GlzYu+nL61BFGW6JgDpb
Cmh9CNrvHEe501dM6SCAeBBLSj4bmWvQjYq700jIF+ME4k7H/dxnSkjQH47VJVDY
TUFYzIrFPSei2bJDt0P507k7FYBoElKH2zjE9jNH9EHIZeoFhAxluoWNIOf7MuGy
FEGrIwdmRMPbw4C2MbmsPSjNvWMOIq8FKm1D1Vj9a52raIByGMUXjtDlTbuQvvQ6
Xsk0MqdqDNIaBhtu414uObDmLRqR04pFaHYQt3enY0Oh9J8fXtq2sp58Xm/8s1Rf
LrQ+ge89JmcvXgxAoFoc6WgJlaH7UK+reC3RqjYdQRmAxkssc/1JnLa8JojwoWom
/P0LrLlX4tdM9ElcrbBo8LO3jBnH2YMA6ktw505Dbs0sQXes2eDCG3Soh9J4WYh/
RMfXc1SQ7Mz5Oxdjro6YtvIlnp8Zh/VLl6dLz0K+VMGc2zYSlciKMCzBkvn4e18o
PIeTr2Pu0e88M4yRkbrNZBoGoYlIEImKjcKR/ov7AL9kjkbsvPKrA7HYMdaPseeg
lpntX5oocmMj7lGEfDQ+fv5uhh99Daj4fr/o0vKo6MFN6t2X03LlUW5GzzfKJKqG
nxBSvhqUoMP2t0OURtTwcy1t/B8hTBhh5oxWG9mn4wxnFs1rQ2qOLq9I3eZ4THlm
WFav/Tjq4IKgtv3ac03qkjz7XQSnyMc640tdCk1n3d7838RQfLecraaIbjM16sDe
TnV2YQPSz1zUGqXyA+6v8NoUG4DQPD2odxwT9Xg3foYcUSY+crJBm12qnF6T04gD
CaHUDholfm71mc5MCH1R4B3HfbdxtxSn/816haC+mfCcpub9bKZPd8QUOniB4fcm
GdhhH/cG/N8oS3Q2We9LEulCjD1f08jGbwNEqzzxd5Po40aVPKw4re43d/x/qyzc
FfpzpYtnpnJ2vuy62eNUAxXMqk/EdT7fcnvoSMCLD6PUJIbZ5vRPB9H45PraNBWq
1Wy8v2X3/sBE20O3dJFfURPqWCT4FVQAN6zJrVkCfPAjsH1j6oRUe7r0vHyXcgpr
axn0wiZJN8rMk2A9jH6KdVDM2ciHp7QlUiUndTSCdzB9i5OOFDAstq9jpgqfsTOl
Gmf7Pfi/NCbZMaingakdPfnf7kDdnT/UFso0tzP9iiclT0cBSUKcUxamNPRc57ft
ox1peGt8dQUKZRPHX7TGlgN+BLnGmZh9OImS7/wU51m8qSm6sMfk5Zzl2Yps5C90
o74US2izzm93+S39MY75w4xEpPAi5YOCskIkqtTq3Co9fXjbENsSHwBDhBrtbimO
UPO0zgDQBo/qfkyCeejFDGJ8r5P3tGMLtQprCdXSo4VXCZpKDvZkX58eaYiQPJYa
IQ77yd3LlTg7YbvKEAPD70Cd90MLJIEsbrIBoa6sN2blBuCG5RrNC7RqSPHpkwFD
nLTO5dujWe0ly83y9NGfQ0ni8lrd54xQhBspM1ch+IQBBgV3ROyEux46zGrkve5z
Yn7lSrveEhSP2k3QMvZ4rkaoWJX0ffX2axzGdcQ6rAyzQBSQ1dTyK/XppB04mSEZ
2bT1EK1nqFBcjsv8/ZGR8RlHlNjWW9XUoLQIzDhsSvxw66A7G8p78cXa74Bkgqbn
KNVUCMjzBhMLJGtU2CTXxCNUebhVHM8cnnvOnLgcf4zaPaA56Q4Ik5i+JclgQt0S
h/Jdr5QS1sMrmVUy9PqhzWQlM1fM+Qd6Nkqil1RQ5ErRNAqIy3R4UII+L3NE517r
k5/HEl/0olIdEeLC2rqono/UDdj4st6zO95lpd1VBGOR73/HkaCVCVCHACNOwJIh
xQjfD6ddCp9makU4nfhlLZZN4vcckGS9LvR19JosCEr4XoRGj2h7mPRC3mCrOyJk
zYWNNpv7X+6lxEFJiZlNaX6ODvU3neu4iDZnG4whTnLkkJ8LaWuJU1PaVysjy2/+
WbgtHYcSJjHigkWanjz5v4eRuy5VT17RpWUvDnt8zTMF3FLAmoM0Lhiqbmd7r3VN
6HTpgYAkNuvQuelaD4bRSXE58g9YcD4qpuEvKvVoJJm66ugbxmSEs+EHc/zpDI9l
AWS8D3k0DplSip/uuvReMlkZ1zwT0XCZLdy0Mte338qkXDTdZRImGIbpR8BZgM5Z
/i+Y+N/IwrReyzoMNjceMYAcEEX+tg4q3EQWqTW1vrDLmFTDD2tpSz5XnBov91Wm
wgoKk1bkNU72gKsRFpGlKbOQmYVQLMmpZICB5wx0KWfyWuCkBDUUxZWZmcQIEWBf
ZkN+H+P3bDlwDhtS63jDvh4ATKuOCtLDOylYi4DjtsVY7pi4VJ52lv2KXWu9EfP+
Aoyr8dQIIt4B39RNj3GGbMHd2G2qpSn0ICuSjnACLEEMug42/xsPctwYyG6P+Rnt
Z6ob71f1rtA9F7gq650AyOer8cRkzih6oWdRUZLfVREoS34Ru015V3o/s2+O9bmo
Zz38a6bygefNIKmULhL7rnKdpf9UUXoj3YZQ+Oup7VONUMyBH+77yLfrsvsi/uXs
UTs1K2ptgT6XOEEsmqsM3D4CGbFgIV8NI56jZcC/b7ByUKFdVeUb1DWKDMeOGihN
O5xDOAN6EPn7jopAatmZzivD7HoRq6z8h15LOJLtCgxHCqxsmfW8rG0jBglZakeH
3V/ZxsGw2EHAJgW5UqZO+PNt50wS3qZDZvflVGMZcIzjJjg76RWaYgSmKxPbkIMH
63zLSiTunp5pJNuUfCrB4Bzh7TPwiMWC60Vs2UXdr8YQJyacVAgd39uJydb0mgXq
aVytV0pt18cytYnkqu7BzCJUtaJkwNtfbAMO2zlH+IJOSCl4DBYe3S9XRkzGJ6eX
k1Km5SqCaPdpVPJ6SLg1QksR9os5zhxLI7RQIDYffp5qlqRr5K3NC7nVZOKP2CE6
EUyAFayjM42odY68oEjCXIq1Ix5ZFkDdDhn4pEFpOEIZ3E7cumpYbXZvXl2ZP7KC
Dxz8dZyW8xnYf4EmBdTBldYy/WCbKLGi6Gk5L7k779HWoVa6azI+txKs+oIFXQj1
eZCa3Xtnl/VFaeFsTjDaEvM2MG6FmrM94+DEWUYgjytPS+dZ3h2nN0/RzqxHdFJW
j7kAHoYuieVg7FQHs0zCPIYuKbgtzIRTdsctrIj11r+JwEzkZPMAfIIJVxJO5wa/
I5HhSRLoQD8ldzR2PdsWg80GvYh1Gj/tnSebb6/7TvG6eSWaGDBx7SYumJ2s/eRR
7HHKo8RJM1DpvUlgAeb6ZRXDLYNWZg/wnUSstDETEfkhcChxUEr2gJz+jPGJqPox
Qp2vh+xhf+9aajn71RR6DmN+5wXtCDCpJ2eGrDHbmcpZ/dtZ7ENyz/WrkeN2fxnV
Ezr/j1/nEYMxXfJoP5PYUvUTGwN9CqJEpsq7uSqR146+IuRJk0njnEcT6RaOkDIn
ZR95ZK22VH+5R/CtjK6YSNZZNCTZw/DXMDWSKlmFQLnChRTTstgkTv9fVCWDfu5t
c8g3dmMdhKu48d+h4IlBWdQZcYiucDfEKDmfbYONFieojyeuIOeGU9d6fzlKBYhM
nxCzbU4DXnCJneqJqLZ9t1ZPEDxt8d0Q7nVUylu09LVT7zqcMEWIxmwh9Y+C7aEC
OBoIa2SjHSwFRdSx2eNqNBrxN1tncGKLVEJ4d5jcfbSHCWJcslHrTwvhwkLLURgu
nkfJtUM794wxGyMf1vTaGgH02YFGEq+bQ2edS78SjwIZmjTB/6Bcaz8WkbpVIdu1
HM+Ba2Onzx1//fL7WTwTa2ceB8iAevXqPCF7bEopmuGSGYrsOd013xP9PPAPtnih
c94byOsVkJlUTcxO1KhMp+pCvoYQBY2wM+ldMsKdp3H5J5d+7qGZvUHiK5tzwqzy
m291V23bBi+XFTR57/EXRyf1TyN6bFB5xyaZ00OcD1N7+vjpUmoqwcZVSbYdjxU9
NnpaDDxVgmToOHiwvBuD/XRwlbYd/fcj4Z7KY90hTkfCPSRGPg0AraIqdC7WaL9V
PenHwZez46BMPP463AGqeQgXW5zzksFKIfat4hm5cchxqbcLY77cnU/gSCIMvRbz
ngTlUqlior/n3g7osOCCXWuZOoZBVtw24xpDXOMk8eOPafhhHdqMixa3ArhLmWbL
Hn8LcJDihnqf4shtvL7lnjLr3wEVwpgjkEOa67H6fsK9QEVUHeGtO5cQexsJ9NGh
ktqDnGEjtpXMdjQdpCEC9Wr/vpx/C0xCHRyv+kzVifANo9tXd51E52Vz7C48u103
tjPMYtvGFT+iP21TmpWsA5t+HcULFpkD5FKxxLIXwVIlm+5knllSPYY7v+Cr3nRv
LW/p3laX4htA6ym951FMTlwRvGltwruSjhiM8MAzqoAFlpKCLxBMzRA0FXXw0TIk
Efc87mKD4Zbcf8EoNc2dsFHDf8jkRkhQ1hAdsRvrS4/yZ+xEL419UN9iFiRURZBU
dKaK3jKDkTMOoXX1fppL06U7yx+fwQTkc1bRWk8qqyZqIIX6veVhsBdHnp/+mAwB
6K1AJUf1drQQMnWZ3MZYBtAmnCf5v1BdzaSnrAotHe08Qkhcw4bs7EW+pK2c3903
yISBisp//0zIg2OQGG040s/WeL7EYRAyvIVjQmExLMixP2r6Uj3MqKYFQhogWzs2
9dNR2hLUOaMiEKpGC3VsLvqVISgJbQTlsLCZX8KKxp/+5lKQrixjr4ePyscu3TRZ
OhhdQgw+7FcbH6Cj6TbyJ/tKGobtCzZNRjwoGOmyOrhZu+t5WZbzs3PPZbb2J0CB
VEi1BCE71cjKZkvqmjSjj03fg6l6wQnbE2Gy5F1gtQpJ4sz/FeD0DfhLjw17BZyk
tnzbzRAyjn0/v5y9RV6e/MoLlqNMvoop7V1Z2xCS+3ktBAMdz2cFpd1mjn3GscLY
/xNKzuynvTvRmfEOE8DJgNUSN3ahr0MZ0HN5N0g36NYG9+4ce04P+9dGoR6wIbN+
sdmE2pvoar+UAUhUKrj5QqiCbrIUVfXeMmtr40gH/vFOsFOaEjGBWJa+elSjXo5U
Hq0WZznQw0dWbY2jiOvtrsKFarDwz8pfv2haMUCwkNhxd43Fj7dKs/b9ex+PCKNc
NsQodQKPasEbe1ZO7da58+XFfnL52TzN+NFxI/kuIUzxaAygHOUN9lgb71MhhHF0
InpeNUh4ObaCM378YnO2b/kWKl+Llf9l4+t0MLRa8zJZ35AhDKwgN9AaVPOv6XoS
kMePQADzC0dKGGJJE+xQS9bqM1s6SX8DdQJ52AzIu0pjUN6OmKcoXUpUzN4Z5DeI
QIWvoai7lR4/fhqqncjihfEnEFw/2wIIFXrFcJ0bH/EpeZNmFwW7oRtsZT5C+etp
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bdJg0vPGj41/PmXEhP+sfjRJWH0kYYt9Lm10Naf1jHlXX7p+YfZi5t4OD+cSfPkK
ojGPupteD6ZEwQ4ZjIHiVF9Ywnq2qg9EIGHO6IJXl07BgBR6BTS4/WAEkxhB48R2
lwWqoi8z0AR+AMP4g/kpdKXt0lFePUu5YCAGBZywAite0hrvgisFYBeNiodtUxdB
EsutLUYn6v/JaWSdhOPg3+QvDrxhlMWx07Dy0nkkqFzXyNu/vGkX9x3ObMGb+XU1
JBYfqcmQYoAFiPBtTrL8X6FoFLxsMs9MnQNWo9CIXXvW8AzEBylaBiqJLzAH5mfI
KIxCuJnDC+MstV612GEs2A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6256 )
`pragma protect data_block
f/8MgKj1mfH2kFrGqr+wnmL0Cbneu8avGBbz8yL0yqUe6ooVXI4Nu3PzbwcOyk0l
fxXMAGvFo96AxTMzW6BOHsRjhoTZE422+EAqKTvAqpIhfvSVbGB3FDZFxWA0xLst
EMC48a06tTVnWNu033Yw9lQJdunVQdMTYnZVvTqItPYnxAbGfIfFXG0DxE7IusIl
JsLAIrbJNAz945de8w1IxK/96rT2Oym0NPkVyA1RIgQ78G67G4txeXDffv7/yN8v
thRoOer1WlUxHlb7jqMT9xdex9d6byGv+RRBorR63Gj2Gb0RtYmfmO7uMcGNo+FB
/tzf0l0P07fuiGVfAX7q8sgMLXWCklg//62FtRwFgj3uvPde2qjIO8gy9/iotV5P
8A7jkDmQEUtevCdwoY+4CuDzrw+KKbNoqwdhHI52J+ezbWSHAROwukG7zl/pzfWO
g1ig/OmA5Wp9Gw5UdfkaTeNZwU54MFLutYw46eQu6/Cb6s3eKPqol7UjG0qu/zmb
G5hZNnt3iOAkacDkGveNCyH8654PZxp259wK2Z+iiOQKhGxRNHghAKmQKR+RV0Wc
ac0VfKfW8HU+IekeScAJYG3z7whYbXzbP5AeRrafVHgRIfKuDYIntRVYs6nJ7p1n
f+s68eTLEBJ0AmJtPoCoTndyholDL3GQqLk4veYY/AkDjMylgbqB7mtCmC+lII7E
n/fWnvykHSEb+srdZDodsS+Mogh1a+mmKKqRILn9tngmHwMOX3pohDsSjEQX+zR5
SPYNE2Dx0cHXcM2OiAPHDYBfEaJxTYPe2hFGfRSzC+yqTy9JG/oWEJ9xKQdtKFJ2
HpuXlSm4Hmdr/YDIcCRqlx+rMXdVt4035csZbvB+UxzySfKEfYWohz4pMZ/KZaEL
GTvBSPldcXpEfwiw1CsYoSh2z0d6gOUGQKNHVRHntbYyyMY5R/d3qGFuw0916Vk5
2bkyhJGPtsxp5jzeW3xmxZ1hB9cr3oYaaiQF1IWBgFK8lidqYPxAkI0tJHxGQI0P
d/BWIZIhZqIBFB0DuxMD1akOsdv5a8I45JJt3U2LcGYIDK6v1iJi/jqb1JfHbFQ5
wJrPS1hperb09zuQctokzv4pNnvGv23iKx8uQXmCpulF+LZbu9n5+fKmaJPBgw9a
M7o6wkWTBJJst8zUjy2uWZRvpaECUyRxOkMk3seFQbr21ZlO5Bgf69zfXvgYcxFr
G+mHOnByVm1C/tSiHW+xzFc7m1JyjBJUCmsS7BmcWIntibAIkelQjtc4NnehWIJf
k6EIIWNofrEfVtl7Z9ceaaq3m18DD/h1qR5l3oRsHyesVRR6QO2d+dssneOwhgw5
92xpEkUILhEGAhxNjQ+fwD2zlsHsNc5kpqJ1UlB7U98JCCgIt5leZGuIY2Nn3LJ8
tBk3c8FVzHNEYUDpGH8yaB/u4UiZWoTLAdUb0sdWHaZdXE2OiqPIeIZUk0YC50X+
Ls5JNqT3c9UOXrHWQNhgxeUKkJhJHneh8sE6y9QuMnGyOYz4S8I1l1NuyAKWIKbu
Ip7Lsx/sEFBYLAZ652Cj4GUtqY2osfPpuniwmiuEK0Gp2Qyu757jQoGKyRGdzKym
OqHfqKnlitOeCzHQ0M8pS7dp7L9XsgKWFCVdFbQeB/QgklAqT6CDlPjLNr6BY58z
N45v9xbYAjT2/v1tt0skqweEJxs3SGJOHH9pu/kczN+rGvNH0/GgJI5jNyRv1DlO
roWeo1XJuH90WZqa1HqNftWxZIRkLvzmQPO2lefIHLj1BdGkkuYkvkrJZDK92VRH
nEIDTk53vXAPADqB/80LCK9VC4liJz2g3UtLxxhyHh1z5DFYcIJ29P8IgEkZdfu1
vQrwfhLlo6IsCDnuGxbeFhnGp9bufpojTqiriEfOjktT6eHSDJvYTRpX5fuOd1Vs
rfVjccMftGmLAvyUcdk6H+SFj8cJd3N+TMy9dscgq4CB3IlJIfzLrkaWIvRdTeQc
X29YPKmUFlPZqGOWWVZD+sE/WvEtjqKeYFJQDfB1i3fzpiaUO6Ka/YgZvT6ZZbq/
bOcjO5o38SAY5XqL7u6JjixF/9+leoBTYrO+2GQiFjNvT1vbbissBNkG6BKXwc4b
4U83Qeu7p4H1sQiBZ9L/p7w4lGIcQOVok5zjxLZtdaHPUk1yb3zdf7k3Cqkbx3ot
VnpDW6Ne46ieFm8062yMuJxghjG5jVIefCsUxgE4oEVVA5DcWekRGnVoU97U1ZR9
5JS32J07ljbOlhVfS4UeP+1GXcdUBJhVIYU5kI6OZVcfl2Lpi9KtQF4BuPHWbDTl
JhxlsgiLWeTEZE0zp+5Gk7V/is4GpWM0Ul6xWV8CKHwH38AlkOKSJsvFvuMxpW6v
na4Z0tVekgeOrdzq2CuOZyr4icknygR1HtlVs2/pCiyW4uk68DIWFZJ2RohUC2ZZ
TK6DDHppA6d7tNz7VpgqQEgmmo5Ku8NrAMxRvTqHz8PtHTSYxBigKTSwrAy/D/ed
fwrnFIanT57hSG086dv9RRKsotkFxkwnJ4PSId8jqVM3ic74yUYPcKzYRgDCfpFA
NhKRNVAJS4o7iv/Aq1E09PcDI4oHkmfbVrkUmOJR9V+2EvwEhIASUuwDvJ0BIZ3t
Nt1GDLN5dd9jsvS7tM/mumIkZcdOETZ5I06/HeAR28MULZbHVtkgo+RvpfeONt1q
y27XqRcp5bE6dHrdvho3P9Z0JzoHpYvG5ATexNNyWszpwopacuHe24xsNUBFjjgT
EVwfug8WMGWTe6eP2k2gJPnNWhNj0MiDKDm4Oj6rdhQQHg3E9LbTIEIh/4HeI1uk
XS2Xcb8MY+btcJpiDKfR+IjkU52knaw3EE4q4XSN3jROdBb77II8XKCUpmSaDKrW
BaM6mob9YDviRTVfaWjX3UNPT2pX/q0y8s68aNxZsSd2LMJty3AGiYe/rgqPDEYm
Cq7lz/XIG9DICrNMOEDWrVkv3vKH1LXvBVJ3eu+CXG/FkLjA92SgoY/h0LGhQ1/9
QwvScgEGnJvbDQGIos3e2s2e56yTHRRXeYP4zKNotjJh2VjqXBwQvczv1iddFuvS
azJ4mXhLRMRU9kb7aff6VgsKRjzYzUaPpXxtaBdPXlTTsVxKfkUwcaeo1/gdiBNt
sTIAFwqy0gXERyp2ZXDhkylOL/qfrfFRp8HpRLlspSZanRwVqlkjfZ1+vZowxwXd
EaEdYiwjzQ/BXz5/slWj2MPAPbfxOoSyrc29ByUAtdp7WuPrBEOm1OZ+4sKQgAA1
NsDSgRjsjWxnWS7rfErqO91Im9nJT7SXBHldP9jgRtcIUz8pkyYvspvHM02DlZMw
icogthAkz0i5rJXK1qOsy6KOswHCUt+Fwq04V2pxtjlLD3KAJEqTIXQABeuNTuO5
t1wrettDmKk1laK99TnMvu+/4b3NsSmzl2Dn++aTIW0ixzYEfidumTria+ND9CCS
juDlKLtJzoF20LBp19vdSwi9Ge8xAGwU7apQ/FluN7iqECIUyz4E3vlknNWf9f3i
jywOt2ixWhhQyjz59g/ggs+yrvW4qg4K+swi2bqA1e4a176DRFzDpkzrV0EfF/n0
tpt4qYp0WVpg267vzsW0Z5KknHDOEV7Yr+SOlEJbQo9tF7tE+LRLgH0uywoRHYXC
AluIput0uRYc8ae6hf7oQpEkobrP0ophgWFF5s0bfwFccKzxpZDiDkHN/b71qmS9
LJukAPqY7PY2D7SE3rFjSdMDU6YM5uRjDXAG8cFo+lKidyK1OnUbEzKMi+84KvTS
ubqbKqqjq9udZ0XBk1YnrSt831FLQLai907Gmtc9tJwnC8Nt29GtvgHd6Crt3Bqv
xY5GzsrsDyFpXXv65mwu5bVCrU04iuN1n9dstarYqRXlMnQBPCCJNP84UyYuRxEk
hZZgRFM8zm+qmBk0bLowC5fXwE8MN19goWp6ighuGq6uxcoqeC+AumhdDP5gX+Xz
72hEWFHrtJQVENgK6yJTgrEr2YXMZZryMaI3xjrf/yxvZVpFsjbcopHvL/Aj221Y
yfz8LL23e3mx/VXO8S+q0bxh5vQPqFL7EtF37K+mXQDDlXZwdpe5qs7ssSY/rUnO
Xi0KgPst1rJbQV6Cm8UH0ZFsSNjqh7jmrAR8eFSWdtD1idK1Ga2AXiVkWXbgOb+5
qSbrNf2FNmXX0afYlUwYIjK6rr7ZcnBd9er9LRCJBNXATMBJhhnHnMnp+aWGWaIz
in7uK+BXWX1AAUhqgc9R8bSrbpL+n3PwIVCFTcdPsUhIV+l/ZBS99g9GTR6+lFe+
maKtJHk3MxCNoYvi/kAaDIsOJl1K62rrUx8EXmaYwAQpwH1kYkycYN4zTzmI5IKe
kEtp/cjlroLfquTQ/PLDfbz2h5OSx7fgFbsGHAtWceYDyakldnAPyzgwm+EN++uK
oHm87TuiBvo2RyO3Q4fynVroIditJz1hpdIbgioZfgi7SY5AaD5btZitzaR0lgbq
d+IgVC63wPA7wGVbhVqXL3kK/1U6zfVa+TtHAoaY0Si55k3ZJIQ8b91rvB5nZe2t
5hC7rlkMKQVAZpLABski5VQFcYNaalARBxaZow+7sLo6v00T4fbGqdoxCGw/90ir
6/RMrkDTip/WIrHu3Rdmw8oJBWYkPMkzfatsPXClNpeC2yUFGM+SppU8CCPhvS/S
7SehXsrFZ4TjBmN/YWIWTBjlYg8qCsUJHBjWxtsowgRZgi989S51rAgec6qZ/ijn
23/5eEm81DASk32xULjuGQmSoZ+tukpT4iEPqi2gimqbz0YjR9NB01zJs8G2/3ep
A3c2y8h9tPUbOjqvy1pwOn6WhApnc8sm140P2pCtjZhsV2ElV9U2W4+JSoFvepIb
sTQ7iSxW8kiXQiIIfaqwn2PIF84FWZ1IQd1HTOLVO5E5Tkmcv74NLG3JDWlAQE/b
LT0MelFBCJUPOM5LzdVwJwxYKGHoNP+btGXrvjciSjk1VQ5zbfpgbRr489OfNB/q
zUb3npzidlvNmEPwixre0Ws335R8SM37KzT8SVN5Y7XyJsRSqb/SD7h+xjhvJPFA
UTbnuUn+VeVAuSYYoR1fPMCXvG8yVNJ/6Ze2wW8qcnwDrsIkLrkmb+M8FrcAfsEy
8c2SlU0kcvIX31GMjKtKLzsdtSuzuj0nFAYfpV/VZWsx+FchX1YUdG9nUsn0iy+g
18zyp8eHhBQG4yQopghYUOcmvqER1mLt9g0pt6Vix6isA7Lb7+RNAgGJ66oWcaB0
iNclXLcxRq+QIXOWQmXs4S4kpFnrSW7WJq2lGU32DogD6tRglYEinDTqBpFLp9qN
iaj/zeNFOSpY/vEF09U/BAInlr9bmIZsXyRL6JPlPiKAjg4dv9k+NYYTUcHVxVJI
UtHmpD9u4PLOrVpVv+ATs0gnXOV3qelXSQD7JHQhv/XRD5ddtIF/h+cKuuimiK0J
FM7NarBJywOTaOZ4UEvS0YMehu9k4wAJpiEZhggAvmEafod2zH0js1wP07/rsTFk
hNmvYHXv/OV496E9ZnXBYtv+kqNenow4jctpZhsvVdmZ+83UAq/M2qZOTHBmzlas
xtVZkLVctsOs3jND5zmklLT3pUjzUw2k9ye1Z1tRs+/VVpacBtQZ3knj+hJbo/rY
5188dLNiaNpvirek49r0wf1yJH3earCf5vstwCKl2DJtwbX+nHL0T1IylVGPDHOn
oFb3YOyWh7YXpK2/SoZVcWK03MNFRKfe6oYVo8DoX2IHoHj7PS3OUW380n54UYBi
sGUC4DmP6tKWA3QV3Qk8TcQq7v794XQPfdcEvu27I/aXTLhhSOiOiu12Dx94YnbP
ZnL2f2ivFouZ2TY8c9UlQV3KyF9oCWHW2a0U7VTmstZTdSWTD7v5QIxEvxw5Zk8v
o0BqI9GBphldAjpMpP5nSIuUNrDSvSy4OWPui0l/vuZvkF4vv2AP6CaMr8XFIJmn
w+lKeC1SaHSH/woVcJLIe4krTkRTbs2qBUdBWKvUkhqXvMfXlD4gtFDz5VH4aA/t
JaqFTHbT8n1j1B26zyVtSFs+WHx8NkWQ73F4j85GcdOL6Hw5k/kSQce2Q970RuA8
UGz9OKrMYN4/c4O1ZLjzCyAm6JTBbwTqbbRk5U2v3p+ewPfOE+NXdoPZz16GIG3+
+YMEbH/rqCraJsFUdBg6aYjH0veMmdSSR0Q/hIspB9I1DrhfhemzuOadzxQUke/s
EGlaLNWUaG+MaNfzX28XMyCPBSOwz2G7A10tyPAtY5OHWa/HykEq2cdsywUwPsNa
2CECvERGcsg6GP+UqUNzddl89ZhWzR3CNNhKH4Hg0tmgPuz0NRx2QmmhxY5Dk9qQ
TtnShIXj+ZzJBQcORChjhG/omg5b3C10+K7PuPbwJ8pu4w3/46ZRk1WVxgDnsytB
64Mj1vdYORgYjetOfScgDSrt6NOb5fkiUHi8hZDl+0jpn163bN35Dhn84wXKXcDK
sQzorDaFbyqMQsjCL4INXLCNED3m/dSVmG1WQqLSwp+grfQ4nKbj6IVezl2irPSS
K2Ef1qmHsFKVrRlRJ1AftktNpj7uDt0YvGm7MsTdlwxUWMwYWVWIITgx/LHmNzKX
s3jiY9iqmX0e75WIZJu325CGDV8aH0ZHkgi9EJ/F69UbIp96sbJUO4BhiIkrUL7U
E7yq+vU+1FJZX9vemcQci0llriLPGTijy+qqtD+eELnW0WVG3DE1imm1m5I2/SPo
PRh7oleubo+1Vtnnpfy4Kq6jREZGmlLReYx53nHbosc8PWekHpZ1nMYRIvth6l0t
2iAdGK4XuAKUJgA3xhG4g9dgNXHEd2PheHrmTQNQeaMCi/6C5G1MJDHTb8/9BSXU
hTmc4qnKY9nYBT83gUxvvbF3ATlr7kOKJPQsvhHlA+NXCr0WKS97/HavcO4iN+eM
vqvhuHg3i1nWAJQk9QKcWdlPxjqqyEQc+Cxmnj4QMv4G7k024iMIBliqMFrcTfRL
1NvDlMQjePP+JNai0ktwxLXP/crgP9VJFY3opylt5XV67GtP6b1fp4oyxORMwdT0
RQLkDQ2VdBGxkvLDKYGZO12uvq3Ei5D+h5W6kLc8OFWwCdPKcmLB+3qudNLJiqgk
s9XFTUhCuHMZUGSAN99HsMX2Q6LBN2uUvWOs00LW8RwTb7aNlSsWt4Hsk7PEuUag
q17cuQ87srLp+K5KeYrs6CDhYk96SKmMwLzxGOiqqHmoOnJRp6Nc31E9O57GGbXj
t3IDxFAaHm4aNs/BZX6tc0U3bOuU2BAu454Qh5Vqvpw7RgXJITRTfRvhN9oqcSph
R+iKfoKn+S9CQec6n5RzCh91OTiZBIxIs+wGfRsTHrWybPnXokbFcCna33RDHkqM
o+gotbzOfoY6Wr6d26hmVSSqMaGmgUJ4I9F6Xsocxmmb6CUSdOhHvsOJrVdIgcN4
UQHzqJJK1cy3PcAVxWgYayBUV6362QQeicIY0V7bqwz2TA/fBuh8Mox6bEF20mVp
Gj7RVWtXj/POrFFnPcnCagYemjlNXPPJ/wpSdlzitbGlf0C7vrrplnfLPasn0fu8
fUIxgrTUzWExaJDswEiGilKOefHnrly9NJT1B3TsOSl1/cMGDJB5bp7teqOHdyCF
dPl2Kmb8Lo5/Jq0FxQNhQyLUtxidGi+tRgg0KceLyIm39vPPBEmgihycj5IzFo/O
i4d0e65qRJFH4Ye3gr0IZ40rTZjPwbEsWISrPChPAPYJKWw35Y3dDrjT4vWaRLL9
Y37qjDnfb3NzQ1k/ey1ehdhC4nlxbp899csDEKX2yshMkD0eNxAUZZjv7HRXYiHz
zsqnCAylzTH46jZa6959gXBkYLVrQOEEoBavXD3LrUkELpLeHUvOwapEKry9QEVE
McnKSqEXWnru0N8szApTyZHHVHT900F4dLYx4R9AwAubqTrcdp2D/UaD4AzbHmCa
p4KCc2215pwJ4XdEylhxN3ifIf6JWDNxG366z6TJBWxyPQR7+vUui6pB7pgBmAIv
bUfJx/FAV2xcqreriimBJgWkZ82NEPwSvNHvACiThiIsNe0c71bmmxfsSdxLkxwh
6FJC+7Vn9+RF0xPWjZxivNsU1kbABkdqZzwQqzWr1S79rmYWG8BoIVwBnqTnNrFg
t+q8Jf5KPL69VPyWhZ8KcbN2G1UkUipQRq6RVmPvp7HyLTuzLN521ZI5JxdUlH22
SCD5DGFx/ZBwXjHbnCAvy9Yn+BXcSu8zCUahyQqj+rm3A1a8MHUw3gtp4nCWTPn1
1DG6TFHzQw9T26/VRArPF6x+zeq2UUEjFPYHM2eRxKbBOJrlfO3cr37LMhGMr4f6
LgFhy0F+p6N/43RZ22i0lg==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
h5YRt2br33UAh57vh7lhtUnA2FIKpVRWfZUZE56g1dvbpj8dwYy00kISC17nyVjk
c94zTgt1IaFkZCLyPx9oPDovH86qbAkNedP56Vn5Si6T6mB+yvg0P8/ll8EUlUCi
fmHzQgkvSlxJsAqmEqdr/e03IdYLdpAKJqJeFl93cRYU6IvgZIBTLmf9DK4p7/1g
ERzUYapuGd/0qSxRUtyt99eUklQkP9TLIYhGFl5STxZfaSRVQaq8bpfttEHy5HBM
h7f+kdKa8lU94EGZM9sPagLxr3Cb94xTuKMo5Dwi4wfRUQR9ZFfboobgQtQMEtPQ
gse+xmqWVdweyHsSTsKF8Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9456 )
`pragma protect data_block
osjvbav/2TkgphBCTpErOV425iq/qSzrMP6ZU/C1uXAke/driN50+jSMyKBJilV/
3RcleyBskACSr2SbqRWvTy/aiyurinaRrPi9SZlBslpRk+z3aEEK8bqcr5TMd6pA
hBCvogY+ZMKiIEsK7MNwCpoBCxa7lf6RY6XiY3N1+s5neS4J7v4zjfIDs16WZFW0
eFplnkZjSLAa3NAKQ3pPm35SsCwYnX59EQlxnJIluulcNB9f3JwL6RZO57ZgkxuR
KF4KYbf4rzguUoOsoIbmxQ2hyfnD3IQnqg0Blb/U4MAFkxFOoIPiYRpzghadgYp+
uIaZWWrkrYyrbcLkJ8Gi/cIBI9Q5EhIZz1rtKIKCaAJdxkgRuqD3Nvw9iym6eMHv
McJMKn/xrdxyr7tois2eodZ7o9aWxYpz92zWMkhX9cDEAC4dNNngEaaVtXvxlIox
lXkZ8WiuZewQb6UUeG2dYdk9iXzv26gpHUDncI6NQLohJMx1x+8TTVyPOoILipCx
fUuXan1rAWYDrxIAKOmLCqodiKRlW5LkIOEYqrVOhC2UXW3z0cNC7F/gPiJYAQYs
lyW2FG52jon2q5u9bZc91iL44DzuzoevenO206WfnRMZ8SDR2zbgaZ5E6ZbnFVrt
ar2ep6NMfyBQjPfgdcawGcFkDrjT4Wa4/UNpgk6WhA4AIaC1iBKBzMcFdzWufTcX
pZ8yYN0ab2PV7ltYpmJjByhbSm0OmNrhYgpCnLeM1UHUUTx/fpIrtek23VrnaENq
asWgnEofKS84ek8LPQ9UrUHmoHEVS+R+Ott6xUcEBoky6nhfA8t9I9b3YmtyHI6M
5x+2WGDJpOsG/bqAVrSQqBgj5+hduaX1l49TbXdk5K624kG0e76/xZ746nGKmCcG
wgZCA0b6VTklBygrpYp56KfRC+z7jPreG469HBnjk1BN6xSebZ1/jiVYI9I4EBJs
pDPWa3Enq+W0brpn2F+Ps658tiSZpl4leNhT8hHMkNfBQtPFj9H3+9ONldLuw9bq
WJWU3rkWniy3JR5qTF77KkW0K0jLPMIK5RZH4NRZe8bWHXTGQMSraRlXGL4D3plZ
JkrUmUEhfe2hfjltZUMwjGkR5TwB9L2LM4X0kqzFhSUpmaLL4ZIV/E0Qiv8lTSZI
LJXuu9e1u2+BzdOYB8lBrr0hpjielyjoF7ANNapQAzYl/2VQAQrwCZTp5EpsT1u+
pR5iDTKO/JiDLusvIKIXrrOmGxuEZsbBMFVpOdHhauBqSaqsCBMwEujMio1SoVq+
06xwxDpacnyH4yNz+ma3NmpmejovDsXRl6zCVmg1MPpJtD8CNjok+t9t+gCWkM0p
N/ViAogTannjnhg6wYwQM6Ajv4RLM2hak2n18gVRVTnIJaOd14lmhTUzRLcB2/BN
W52gfT8kpDDcpm1y/BhFHgZIITsQQGM7XbWlWciDitJTERlpk/goOYJNjKs22miw
cY2VWFliySCCWwMXCKfowrF2gOZv5JQNfGYB3h+TF+qQFQ4am9Hot5bAQ8o/frW/
sEh+8yBnIzD8OPDfoOQjbs7U785kJ5KLoaa/FwIlxQEZuIexhxi4XPAqlpOTUA9v
7A29X2Pq92PBcdW5h2D6Ms/ydJa8qxwM+MRdI//zm1wPKLBmNg5b8uW4j+nvAG0r
z4gYAxLdteXQE3b4MkbHLa0LL48BKF9YVf4N4IC8AvvfhaJT0/Zycf+2p0a6i5p/
BllIH2suS469G0BaX0C4WTs5SipWYdXWp7aar9hF8nK+rOKdwfutb1yW5FDxOE96
WaeZc/4vb1wR3ZTuYlWkQe6zxGYP4wUgRq4+zZ/r8+7htgMK8aKjko+ddAz9kmYr
r/auU3O8FpWLY8VHxS4eRsG+Bt90/hU7603aJkbgKyjQlhPbxsC8ASttx8HLdnVq
2CWmrYhdgDrCjrHzrHOUc1tKqnXxqy9lTf3Qcb+Z+kyomjJkdYvUnyqysMo2lnS4
iiaAod01lJlLZXrioFUblywJr1uvBcJ7rNUC8WFskOMmcdRExstOUSjnusk4mWIp
cKH1qe8mGHEz7LfBf7V/kkxoQ3OdAXmmPeL/1IEnM6hyxY/PKhaBQ56aeFpXO/ex
uSkpH7ONE2mFEqCFRgbe5rkB1T42jZ4CDO3Wd4xSTj399UDeSA4ZjYdeIYYfU+E5
VgnD3PmfVywGV19KBEqovLOfri7BtnBaVKg/gJL+e71iA1/8V4L++EDvcSttHLvm
CH0LD2Hayo1lGXcoKYiWVrrf/SloxDDtqJ9Z5NXf5MEfiyCycOuPyfsPsEZOThok
6NdTEYZOWBOJyY1xqtIM1GNTKjwebirSZa3ro4JWWDpaeczrCguxr2LCDQQewtLc
bK2c9hplj9pSnbEQYjQExWVdj0G/p0dNhSdLV3JsOHpyF3ZXNlS7A2dl4N/IdeBX
nlwcx8fDiTXR/LZqi/h5/rhBvAr2zkbHv0r12pJPfP3QE/do2YK4dS/1lhWYu/8y
eSFGBDb5SM0KvqDZrUX1BJFtYNF6BcqHygqnFiYF2BXwr4sBZhlAQZH8bHA9HP54
uM1dz+QJZi4canTRglxOXgQYbL0r487i+SCvKF5Ix4xuKWKXqubZJtjXo6AoO7rn
55oXoNbToZDhv1n44CBtylEL48CFcRx1dxZdCPaV9DtWxjIBX3XD4qtujWl91xlK
EBTqsyd/QVpEeSG/YZ+A0VZdF/wuj1x3VkgGmdKf8wsLjnLmpqIpQaXc3dLE4ycC
VKQE5PwkjapFo0kUPihjWn4/qfpqhwWD3YRFHCj5zn20miFVEPjYQ6MBSzNizVJp
9DkUYHC867GcunzAPdZhfTwXKt02pUPU9Z7WaqS54RnbROwl2lWj0AD7hKp6ibrB
CSH1M8sNsqrV6pxGCRgsireAfyy/NE9uwWIAYIZYuQUzkLIVE+nEc0k3Ab7UsQmC
Vbjm8owq85kbV2EbeyQWPM4dnoduNHirGEo8Ord+CVTJ0mDCREWB55Lcz3dfy+U1
XKm98opYqt8pxUi0ta+gjPUpvYxx6eT8T5exz6cbdwupqxWSx/pVJK5X5t7uW6G4
9/1ThsSL0fcdneWOTKtnCFlds26D98vDVrMoXyCEVtHiN0W+HgSluEQ8BU1LSmo6
wAlnY/cDISgplMqZXqphoEDQYh0PPuhgNmCLZjDx5PtF8MU2M6r6MvcGXyB0r4mn
6hEzLagQj6L6XGV27r/KG0MPE0lQr6aaJ1DvUDWvx+73Xd9xW1L/bCFUF3UvHm7m
InR/UlJ/wfIhL1JN1AHpCtEoxyn/QtLCK27RqzNL1hXmlkz0MZOvgBAiYTY10Wxk
wtH2pWcuIOasBVhHkaRbYs2Znn3N3earGac5U8URkrVi0lTbLKAQDCe+KwTR3QVa
owow1E7SAzczL/EMBHa8tEZBoU+9acw54nKh7t6l76ErxuutqQHiYRmTFV7vjbnJ
Ms12iHgZT6onxnEpOIuGflY8HYvj7pwi1qHVR3icpLFK2CVbjjrkiOzJ7BLgGkGe
PWFADeWQMZGGIfQzWw0b/LtJ2NKXA/nWQxhiNM/SQRVBS7175b9llxldwpFNsihR
Rj5ilKML1NEV4V+GVZtH/w10ZgiwQ/9W3jHJzF9CAzbNS2ZLHfgrl5S9Q0Fbc66S
QZR5Tzn8h4uDWcHFeDcSKlqP9CsYYxweK3+YaaYOd4PC8z6bYG2yrc+eyCcJGsOC
/mtCKCWMx/YczVfh9chq21jjcthWKLueVW5iM3qD1VMp7oXuL4UXT6qPmcn+EfsA
fXDXsygW1Tepkn6IkrC/eDIUhwvMIfUUxPRhbnf0muSo1Aq8oSYgk/urps26gtQw
SDxSU8AqYok33whgV5q7jFq29wNsXmg/UdnNEBeCFLPr578qa9vDQCf8+/CrtU4H
uTdppQVmjn+n4kEpROtZsWGFjjs4gZ0E1BTBbWyNZeCpNh4tAaYKEHctSSijdVWT
zvas2t6WUFW/g+k4wBpnq3+6sfCMxUF0NY7H2wSezq7SNmUMyBwk/1OducUXMz2l
CBa7ANFvVvNwm4+fwyMjPBT+owGKitHeKxyhYTw43zHfaHGxpuScOOcMzbxjrpfs
uhOsb8P4VcL+CghtEWLWD/wILYaAQGu4ewgSGDidNbMuvBmbTwcRstaWXsbDwmOy
Nc66QZlSqIYvin+V/toMYUmdowEGe4flA3RlQmwXQ9HHICD4rARuBHOJK4aKGbKf
OpXnDVqICEci4JAfS791SqBWZGshVe8IDrdgNslTRwyMJwQgrlWTFuYxWPT8E1Jv
bejnljr5x+NpdQQwOeQJUnR65bIzmbXdFpl4v9DRPMciTB7CJpNlle1byokgUTOr
b7kC4s6E16tHgNJSHDS//QwvZDTcwupjW7O/dAJ9mOGSumfn+jAkUqVxvbfVZI43
CMEB8CK0fC94O0PJWWkxOsxyQjsT78sy9CjXu1Ip88kedC4aMm70geVuWQyImeLQ
QAwieBXcOhiKIChkd86HcbgvcfdfpH9mTQLeXoglJ56MUqdNOIwIs1U5hc5QV3Mx
pkQP4dpabhzLkr+rhDmy7Cgr/lcFbz5HyvH5IzTU1kLQhGyJozZxo5GxnxsMxmhD
NR5zu2cUQEQKQU/5hL9phYrRNHI+pAYJVnXTD6u3xyexdCQBkAPaHZgb0NeRPZ1g
lB0GBxvRa+oDkTkzTRJU5IvG18C95BCtHzFN9aTypenrecqAJBH192Ylcn750UuS
MR16s6T5+65Gtn8akM9oZ2Ob6CQeD7DmqdyPoqZSRG5Z4ixBundnm6VbEKUtuXk7
PEEaDxkib6taC/9zNPkAn8CX/CKAJ/g+d4XoWbarsB9GmhaIKykPcU1lpJc0hgyR
FA4n6NEDcivrpwbsyzAPzKaygq6D7dYPZSdexBhkfaXBlYV+bjuJQKCndLPMmAk1
JY0y7ytudoXT6CnNTT3nURIff7L27U6NRT6BQSiFtI76xtMPdGB3nY6hLZRBWQh8
f8RcrM1CAehVg55r+8u8Vg2BPF3zG4zI0Tr9EbzKYgSArSK/Mu7ZGmzlQDR0xpqq
v2Tf7/1bPg6WTQkOB37vjWbMHeWNRBra+5TnQm3bm6RaPpGuKe+Ib+04AXBk6qzD
5uyYpphaGPoIyL79c0cccPItxOZyImxaxvFl+82KTpJ0tEZAHCkhZ9tzV1gg7wy9
pNKI40xiPbh+dOtjaXcxYyUOnW6C7m2Yd7TSnaoT/ugIrsi+KmtiwTxG17nFFyVM
mz+n7ds9HgoQLUb3bO+R8CvmjXL1FIGqFBN58pRs0WuVcob2xsKbsL0n3gozi7+U
NDy7FWyQ17w4ey13H0OqoBG8JSvCApv6d+e6G00LvSTN+wBX58dqsNHukwxo2ImP
OFYMlgubjw8BMI0pP+VFVdAP3CZxYx0wnWfjuhQhCKwTC2efFqUmA1SLbWm29KCE
EQ47+Ldf8yX+Qy7jHNTaK6X0A1BPwPpqiMU/VUSBJDBJGQ6vyrPkD3+lAHKdbxhD
Pov4SrPOS1h69TbpelXFSn95l2OwWARuHVlv//X439YnDoGhKSmbiryaHhiNW2BO
csW2ot6NTFUO8tSk1zqTcS2jDifvvJnnZGw/QnnYkcQMd8W1+9Qt8ISbio3JwxL6
V60WV8BLxFAC32bHXp938376eBoQHGKcfjGNifoAQUFzYp+vuyT9PlVv+WUAFTMr
GG3LU6rwP2gA/CIHPRWxawDNh10t8SHUE3InoBsGCpthDWzgiTmUJUFR2NjsRyar
iNCU9uWAr/0hCrkHNRUC/bKFW6g90Z8LwIaPdglkrJCSBb9+YzKo9hCr0NJLhSNI
Gy3+AmMiX79Ro0S2ZDjz8SNVhN39ZhordZZ8TOVpDGf/CvxCrfOGa9pWR7KaQvqA
B+nt9ilfDwLgeoLKsU/ctkGcr4K5uPy0dLSmWEgSxoPF3uyu9/QUjMDOEvf5Lcbf
x0sB6mEenTGDna9hzm6bJmT07s2ElAtbhg/RJxsNrBzHqIWL3CguSCRxkYpxv4pf
Laclm6k57kzsvs0uWTWG5BcbZdJjHptY6TcfhfNn/JCu14dD7XN+MyYnYCa/vrdm
tjy1BAUk2ZbTpbm0wym8QYqFB7BT3PlXqADG6v0PpAAFpb4/gxaLIpV4sfb7uWZ0
YqYt4uM+jD15omlRKEgOw/q+6llO2m/vKLtuCJgSgsybrpDf5STL/ekaST1V0QAG
Fa+ABJICcxPVIdXZow8R2UqUG7WgZe4HzezBQmrWfC+U4b7JhHpXbqcuZrn8Vw6k
moKvq3xzmMaygImet3Huo7OCS2l0zivMs0JV/ZVugW6pIz8urdE7NWBBE4s0lXoA
Y8C2/xkTWeN6MoSptPR4SjlMxqeRnHfW7yUiH/lI4ZoXyvO8WNw8E7J7OIuS68Ff
JYcYa69OgHhfB+5BEV5SHQbDWybQvr5LBw+8cLTyQ1JmdDx/s1J3vwVHY+pbPryz
033kUoHFtU7d1Dvj8ORNTOd5D3ztb8LhNRm1wNUp7y5oqgr2L1voX6UhlrzZySWB
cm0cf2TVapHwq1un8zOZPbBPV8MC8qFIVD46u84Tdmo5acVEeEhNiVIoBUHvTjwY
cogyUblVUfHUX4VSpdTHgqK2+HpIzKdr3gSo0fttiNoO9hJFewgZcUjYNdVW7j8j
t3L557DCYnF5S6H/uDz494S5F7tX8TSinbprRlufEAUtExevl+yzLES0M2lnyZDz
4+4SDB3yDCwVB/UFsnYFylW0GIJPNh/NoYaOIGvEHkQp8NOBd1a78aL9Trd8bSfN
8jCBKa7/2Xku5Essg+8DMAL7NkNhfRf07mkHlyaj5DL7JwqaN5vaPiqkyguNAE2V
OijKFpo4Zp/8aYxFI1NGTQhRHrJwJsJ+UoLI08byFIub8buqyD5EywjviJimp+z/
E37fsfvXrcuNP55jv4xmvwmFT626u6pPlTGBkGoTkkYwPN+i/pJzdU1o2hRVXlQW
2LVzY4D6hXJMFfeRPRL5La7QTwo2xCRe6VHjUqvAt5z/5AwY/IxcCY1bSjAOi25C
JofPAxwGsK97asNRrvu95SMbE8lNPFbqeJCnyLEhBc8iSHugJHV7p+Zrh+5SsWRy
fbxoJXX6fO9YlyihYGv5f5jvvc+reJt+z9fsEX1Dq4RhDF2SN3gzGLMuMXX+3gDY
OTbDZTShrLQmr83q7ebY4kmIxlCte11kR7N47QOehsNojCqKe6YCXRsacSO9kFsZ
If03IlhWUanJ59zisKnXyM4R1J9eOMBvroQWf99T6TaDNGPOhZ1Mr6zd+1F1Qfwh
IfgPWQY9NRgCrJwf5N4pBvmsg4htqfThLobmtCYmPnAinRLvJq1JpTNc11+yUpJh
b4D2mYwR/3ISNKSSujR7B92+WDIjwxSZwYN9lC8VSShB3iUb7cIvEV1CrkGc+mwb
4aCZByVKRHMPw/CpJH7B1oIbxZdoJ3s+b0zHaxpIG6xmaEWqRQW2PPD80rqyTnCT
u94GXkFhrNSduGduHmQtCtqLN1CBNrP9bICV9+Sx2PzoO6k5OJImo5bOX6yAHhv/
WtT3ld0uYnAdfAOBPdVRE9QU+csfw5zyOGVi1MFmEaS7lEhZ6S+ij6i2NmEWSUZm
ybnGqpTPKRFKBC9z1iDgPJuA40W/zWlysMQ6wKk150rDQqCuGQNZXnGpPzSwAugS
q58t8vVn3ferP4sW6O1Cdb/B6FVZcYqzV9u14Rv526LheFYUjEU5X8Kg+4cfZY3L
/b2vKKh/WfmULnjNfxPFVng+My0atgpDX8tQO04W+LxX1G8AGhVGX6a6fpAa2wnq
4xB2Ye5vZHUws836zDLqT9635kHlMZZJu/BRGxnyJLy+QAT6Co0ch/etKeJrUPT2
FnwOKZka7HMR8EsEzZt0J/4tcH6f1jjOFOqjPRd4kgVECcTx3/hYqGZpTzoyakTJ
UlS/l9nSkR6SlxD76DsO+Yzj+7ZDsWFcWscg+g72mlx5Lmq7pEENGr0X8PkXNhqj
Iq0ZMEDvz1fPzYiRNHv3s6COvj1BFTDO2Cpt5fIAC3XWXkNWsPR3kVFyYObwGzLA
ukfKEPVmPxrF9wt/34SIERVykOewLeagAamZmwLcNSD1zd89uPUfZtpZdM4MzKPT
lN2Pdqv2Rrgr0jtWg9lDaJvixI4k6AJJTXyLXORIociTd7vdhx+5htjPwZcAG+tY
Luew4Ucj1zbFaw+dIYaxXnGsfQgnL73tyuvQkGL1lWmUGua+HW+piTfl6N8PMuWs
3sfP1CFb6bu8F/JHGZQuylAZhgyfPJfAV+rVRPHVFd4FIovDR0AOJ3bBv/nKu7vb
WQPSFHJGuVNdvy6Jw6Kv6qDWoGtfmuLvEeOqmwNAe3XGXkO1j5S/+nvYpGKylqts
aG0Je/TIdvmbFq1T7xZcHJHbHEiMLCoD311v9oDYOhAluV/WX2lnPCWPLDL2Kcr9
sTT4+NBSbJL4Btpd1OvXDp50fQSd/azMxzAD6P7/LP7B4yIWkx7jvANb2uoWckaR
wJBgFnXNtZ1xcP5yhmclo9m6oOsd4zf3U8A82w7u8B9fu8nxf9slY0ijm0kaEqO0
mOBKDu+BYUVaV54geK43QF6/xVH3+eZDaSHh1qE/S9M4EfyrNTnmRsGIv66C7tqM
ifI8E3wv3ij9chBwmBdH56vWZpYg46q0iBeRdMedrPfpBJIzXXbMIwdbJD67cevc
M7LIdZYoPjzme8LgrXRLbtUxbpV52tye2qhSY+U04AmgMJXuShLphZqulr241Hkr
hKj/3aC96iXnNmd167qtxggnYm2EVZR2ZWzvvSD+tdMw41AATvLNSMZvr0fkpHjJ
+irhnpckXNqCrwfxQIZM54xTfv7ivlscpOH5MSWX+2tdRPzKtyXTyUMn2/Gqtr89
rOilbBQzEZAjuJn3Xz8GF370lVpmqtsYHO7w0DoSDdtDWM8WgQWg/6xMrs5JUp3x
WvBh86E5Uw4f/vTOBM80XRPZsXDsjMZJo4nE0H9UtuC74AWU5RLJ66OBihD3gtSe
9SgXsdwXQ9q95Vw/OXCpwxy6Asil89SQoephYdz9j0jQNXHCvJzeYzZU5LieNugN
XEd9YXJ166mxwxjrP1exVUB+tuWliaJtfhnB/WQJIrlZy/F8bIqJVbK2AQ4wvz/D
PRYh4FkahmJ7+YOFvVCmDSalEw35dRo0oorYBGRl5HMmRPYesYE0Xixai6y7N8jZ
4ieMpzRFpYO4FhPdFY1Jh+o5QqjHj6JUcev7SdEGwlA4iz4S7GJtWTlCFqQK/fES
9r0Sk9HKYfH7w7zLeBc13NRj7ONhABxoQBOE2XgNwVMhX3kGfDwOW+EkMAH0SeV6
TGlxIOE9rPjpuVS5wsxUs2KmigrEfiSjrZAAXpo0Irt5lE0ZZREeB2KyT5nAEv/z
4bgokdHYGGrKrnj0cVsptxKpgVTSmFIrvu4LDZyJ+HfAVrdzV0ddC/9/UmyZcIVb
IF+YDYRzMTZ4P7dSpYMnCqdMq+/vcRhW7SpqYP0qK3IuJLKLkMiEubkwGR6AsGtd
Fu9EF7CjMP6yZGFRPXtczN++DyVXpjMW6RreVGsIYB7x+J59VEk90hdTsitMqIr/
aGKyGDP2fVCq3if3K83AwVvXAkeP97t3PK4HmtDctLiM3fOHl8KylrUwiBNm/rBn
uz8fAri986gL08GEK8x7X49nK009ClEdYxXyQU2b3i5esZ2dH8UqHxB8E5225zvg
IO2gtEBC6WrzoMUq8hNupoAFDLHqzfr/NnZMkiph/vaPy6Rg27rWhdBOn+J7vts3
TEjhsmEASFMSL89tBvd1C6fL0MvnX6G12RRaXvCvWd55j+xwVpPmNyD7V4M5uLNW
IC2yGuw1B2fJBNhrINJ84h0hozvr4xO0s0n8xO8V5fbNjoX8rgywhzOxh/3K2P8w
suB6NOtNT66gELHAElEKNxJ0NDsvRLbGrNg10eL2+0QSTLj8p2h4pCC7z7HTXMNp
8ATpjgCS9J7ohze8yEQ+p+WZAaa2f3PwKc4R57bOdk5KfOUDQozra06Qrmg8bZY2
CO3sqPG6Kn16vEUnIl96QNBi6BoRxj+J9AmDL5zXek9FcJ4Z5nIKSVLFI3rOPUes
6H/ZhG8PKo4U56BfwcwrS9VeCgWC91sU7sBV+PcL7D9woiEZDqyscJejy5FoMU6+
mhXNlKrWtCytljel2Ad4nyHTji3Z/WZTSG+2aBLneIezgeckMKUBtDKvGYUVgebh
noUk0A7aalvaGVMFd4poZXUfZIIMxjH5w9EFFOrZcyK2bDhRD10n9hxY9utUntIM
BaaYBB0oMAYHGOk7avoO7m79B6jtgwUuUJ7dNiABIgEpzzTW3v20LTeZnhm+393n
T/jlFR1wO/R/qqaQM1paz/GbddG5NIh0EGk6ARntV0J2gT4pETCm/w3Z7Dh+yF2E
HMmVVGi64HWWXn+YuEuvUDm71qoa0xqUT1XFhv5xmggQ2u46l2tG8XtE9KLuIVZk
nfOQgZkjwBbKbPckz/La90rTc8h9b32Lwr1f8NCxAJ33em2ugmSwTyegZQm23I9i
QVQcM3PU+22k55HnRSohq8DGImjBV+GefyafMvOThaqasv3fxtJmhQ4bIfRZn23o
sBeOq8COnn7+Wbr+AXDOjVYoD13pHDmulRDW/5ZkGrtcChsU6gMna9xfxkvVTSn8
qTdB3MvFY8L+v1WFOrzjH2IUZ4+vYdOfXN3UWOVuajpqre59FQjJjSHlsmwLMe/u
77QJkTC8klHucZzKl8rhgGq+m33uNXoFTbnH4/bECuhSTibGENeBTIDwCYCM4+5F
obqWFJXIAxewzFRp54EJnCUSvh6BeL2ZobfHyyoHTuz6OMyeUHIF3hUug3CSgG+0
f4mF4Lbm/pII8KzEtf1CY8qzVCzAsaxS6gpvOgdVbz61BV+yyutPUpDdZq5sNo8p
v8gzggHEQjPqZbmHgY3VJ2BwRpe7QI/VePPhvTeJkYTRzOM0O8tYr8xcOWii/Y52
BE2YQaOnhe7TLGNQFfdvninvce73grMVLWqByr1hDQOtXeTRBII7HJ8hQqPIWmTy
EnByu6sMN/jITPMiHZDtuwFdFWVDdqujlWaIRzrS7F/uncQTtBh+d1ObmopwFy/c
xSr7WYECzk5XZlGE9GEZgiAU3hmnU7VPcsT0yrlI3yKamrciyFPaIa0ZRq5fv80/
sunwBLfo9jVjQKEPGPtmPCym1rAq7RjG/PscIdJaj9p6CS7pqF3qhG6pjtjHtEYy
2rObdHuLQvjv5rFcOczTYxei7PKSVY1yVVZQBCRgh78HJlNUUw/j4eMgk71RTRSj
PMSIzi+H5wAfzvKZ7T6rx/rFy5P3a9B94dvccyzyGqm5V8flbPh99Q5DTN/cHzo1
ALPAJV4BghL/H/0SKtnrz9PzvdQKFPAaehoxJsxQ5wJsA8Nmf52m/3Eh5RjWzPx/
O4+XUBI+Zv/NoPxc/14IO6FNn+sDfdP0172nkMxNY2TCJLT+90SbYGohh1SsUHg3
2DDNh7O5IuGTLiQwGmcsX5R+Pjo0jdRQaCVFcDbB/ytk1sjU/FbqNskOKfYwyS4e
dhpA9aiwiJRy3c9r/xeBhIEsg+gHWAqgJs2udKZjG+DkC2A+WityQG1DaaL4/fo1
WfF4YMv9MoqHfX7lfKCAxeQLMcpcQFFsh56qWensrlV3uEWMeERKL3BPV9PKaMQd
FX3O0x9JqycElhvsXk7hdihsa6JCP5/1y86W08xk5bTNMJmwReAVWW9YSgPpLdkd
fSb8OTGBrgZL0feGsqhBkKLKo8QTvym/vWiHg00vLml3eIoJyc943o0fBT/MjmMF
HFjBzCoaMkFc8X7e6fvcdj5XgtYjuaShwkImHfTpF6Y4I4XJuQVc4fPHca4tgEcT
k9AETJdpV30Ai7fSX2IDupTU/gONlrVYs2/mvXuVwsSGnu7iv41i5pbJyBMne09X
aVx5b5UeVbdBFyGfapHQoGaEstL60hzJoFHg/eB0J3hfEbCOMRb52r1i5TPRtgVO
8GkICJeX4hQaoYDcnwkGV0OSbi8bdXyQ2l5Ch9V4I1RJnUE+hOvgqo7LYTCWY0yb
/5nIjJAJWyGZQg6VpD/+34VKiLtZLB8TL1nTb0XTcd9R19iSCarzoBx8/VL/O4RP
KEY3K5OCdvLJO56fu6DN9a9uM8F9Of8SSUJ8dquoNIcmd5wGMLp4V1eTEU380yok
xhHIGWoOyvl/R3eCvxu9A0+KvAU7e3NILdchnZTWTeRfjXJe2whTi3jBbFxtBWRt
mIw/sr7siwXWwF/32m6vZgxZYn/R4uqFNc4u3/YhrrYgFAaiCa5VXCiZsVfnDNFB
6JpKDYGJ5Lb369vKVqUOUkOz34TfVFhzNaKQ9SRrPoGjgbOv+ryArC+kCMkbLYy/
hf+CyBBWsA2zuzRPfIpqgSS3jTpjDMkBATu0BrjaCFvHK7/yga6NBlQw+ZhbP8S8
p6NyuUyxTbAxhqy+818AuBBHnKSVRczPbdb5b/U3arhtogT11fL5or0LlGwKlEfc
uJg8EZ8M+/vs6WHa0YlAgsAvzpWE4/9wVMwuzBo8l0Me47cjF+9n5VLDFiPQwrdK
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
F0pmnADoOCLIqA7f9grxLBEr3LxDikKCKDmtgZDHh/dp7DNpSpkxShnyEQbzDGJn
TyxhY0TzTmcxp/yd8k/vykyig4wJk8b4K+OXzuA+MdTf9aYt7cNkdrTFH3QJlh4T
papZkxefDw+91auwqKCvzOw8W6NM94B/CQHkpl64OqqYHyRk0bfJHDqsJceYOd9c
fG6dDllFTUD71Boi7M/4tcm7rA+vOsMVNDZtF0vIZPv9IjcEOf6gfxjV8KVK03D1
07Ern+/0gv1bDRMIdO0EPNDWNYZV0QH/QbZyjllV/NBX1PAU0k8R/RTZu6wnTyUi
pOOxVR2loig8PAzVhNmlYg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2672 )
`pragma protect data_block
5B20PeKkJ4+a1S0/RWLAXxLOq7lLWuQwFhMhYEJ7xGdsntvP8CCayXumcLWMjP9d
7HXAsDw1QExN0+eKZvx8l/L86p1QfQ0BJsX8HEQ16GPY4YzLwkdcMQS2qvxRcGv4
r5FhqN56MPJgX1fZkNtDJoThfjh/iqMS7at9fjOqeBltijSAgD9YhPLYJxfZlgTc
qSxjEqyj4Be859SRFF/UgaIWzU0xjif0ptOYM8/XMER6ZkmgnYYjTLUZpJgGzGkw
PuIPA5lQGJINSradZWxHguIEJMuooSDIDHiYocZh6n5uWMw8KG7HjIUgH42Wbt5v
j89+lpD3z+iuoxGl2ybN4pDVvL7KbZ7xeaApD0Bq7e7RUYOATiZBoOxj/HvzDbVk
y/stCpWVRr4ShtTuoEu7oqUzO9ah85O/28nQj8OpaGdAT5Df0hEoNdlJWeXQ18za
18l8Vqx+z+jZ8kSimuxYFNqSrxuPuW1ZfRvf60GNW8WVZ7iwYWHt0ZCS63/qBeL2
9YCTNwIOFN5Ep3Iv8S5CxzIv+dzigQ8ptcbJy/zYOy78c5DKbSopwwJdhl+FCnJX
Z2fV8o7T6BdmAH4o75W3TCIIJ7SfqpreUoXOOXHsQVqsKajA6cMeMkr1vpGfoERc
SUGUB/wvC3YhmA1XuBfCpssorToF3A5UNAiGhM4ekXUmPAl3C50RnyF1Fchv7aJY
8HkPCDk7RrHG8PJaXJoQgAc2RAoyOqonanI2O74Qrx0VlUJcDD/Rkje8AopFaUPL
elW2CK5xCFG0A/pEOiZrJ+qAjbCPG8BFvnLeagSfGDgFllCDMK9EiFgLlZqokGR5
LNHGYNw83aebCX8hmfnkJCuThX4fF29UtsN5uYQlyGI/9CD7VY7mkBasooVXzG+k
NQ6FgaBrxaMCPFSV3gesH2az8v32m+cXz0+JGdoVRyZUmlxMhQwX7YPD2+ECntlx
+BoKspqmQ/topXhCUESLxwoVuQC66qxoqQbvNIE8Bsfz/dEOoCJ8B0oGBB7YIceW
ZPDxijAUraV5pkbhF7l8U/EvL4MNdRjKlMqYM1/8tVQfYKnZ4X0pqBfbjCZV9B+N
esmqQDPreFiOTMLjRmnhhyjnqcupTiMdKCN3zI0I3DG4q+HqdWO0Kp14S8OC+LsF
j/fVr3G8QZqPjIEuAXKvC8/cuMMKr2i45PHEAq+wo8N/luqm1VGqsVBdnt4+3jd0
PAIBeYWJ9o1qIMBSOPiC5RmAFBdMwW4lVJpKl9wnRKWPCHJq6xPMFVkAoR9KluoA
v7RNQi3cZhLekCZFCd2tzt3TlnDhk1QEwIB614EV7o0nvZeHdfEh0dhxLOv+sZyB
zcB3S5605pdtxlwWYtlI+5CKR6DBZN4RLKZ5+olWe82xvx2/SdbtM6vUO1RXAosq
QqAM+p1J8pzeANGoKpn26Eg7iYh0P8ohWjj0yDTuPx/95RFVCIGV0fP0S+Cxdyl3
rn9BkaPNKxmWeWp4UzDvCWNtfLhHu2yIOfl313EPiKg84N7MdJiwIuOMQQfycdvc
RsNYdH78w3Hs2QgnGsZjIohbgsfUEdllpijfXFM1yYj+MFGz+NiydhX0/wAaAl2C
xwRpzdHoX23Yu+enwHvgd8PDdCA8g+k+7wIQIlUzItcoBYhRYkBYmgI8woekIkSD
B983uhQro21KfAgwbJpgVvJE4PmuZLJCcJ7I8Xzh6Wu4lEP9tGnhX9wdNbHQyjrP
+DZ3+jQE7MWEs9wX3EM8bIn7ggROctCddiHehtWhPcoBCW2zWgbKLqhp3swP1G0M
BCj5FQ9VB1lf2UcN+j499PYTCC7H1ynNGZgNxS98j+ggVRSJT0J2WT7sDUQO8SLI
xWI8b5fUHcUq5EkpabF1kdOtOLVmFxE8VqBl8ejud45S+Y8uah20DexZfp65fYOL
Z79xaPJxfuQn0SjwqO5Mw+CjC/HyP02UBSb1X3i5PKb46DI4JMWpZOlrSBOhzMt7
/AS+bYgMabp23UcN4wu1cU1tit9QfQnNLgWguH/AKJ8lrFq3c1rZ5FMF9Feqxvh+
FH9uSe3rKSvpefZquDX6Hy+N7lvCILnG3ApEUnXtKR2ZMX69nVlcHYgDTRUzNFmc
bYtFJ7qn9nN1csCgRuT28Yd6tb1pIKdNvXeLxjqgOj+nYhvGw8DV7OPZiBgvpDso
F3qMZY2EnQiCdRY+Nb7wRGiTKzHBqAiPg9jfHsHTwVyeg3GsP/FGW19fHsPJwY3T
X4LpO3mQF/d3W5V03QQ7f831WAO5MRkI4YZa8a7VtU3f+jd12Cn1vynozTIeFYZe
cNCruImY3/gHGS8F7BrIHM5S31PAbP71jM+t+RufA55axX9lWSsFS7ZGIfFH5mNn
VAisE60y0j35LZM019AHZwAui8Qmcbhj8OxkGnFibPyg0xJDHbRJbjoeWiBiZR15
QlbKQvzic6V1JJT7aP9cfCkHzxHAqAEN3EZburIW2iAau54krXqzliHm65R5GcEQ
WZT7VF71uty9Zg6JyISp52vP17aIx+SawtyAn2aaPOvcWMJ/aBxxiitBEFoo7FvM
WqPEeWV/pjFsBlD73oy6JhJXI+Ng0WlI+6jSj5wQPtWFSP5KA6nNiF7RFIekp2La
idSy/I/jAss4lp1pVZYnym8GjN8POumHSquftCrEC65Hd0+unSOaMwJStArFcx2j
zsmcMBYeo17F8vuPj/OhRE2duTnkhgqBPPzwPdCrUST+RwKAzgZ3zQ+18ltId3NO
hA1W/QH/IBmubj3VlLSFzCO82TovqBW0wyGHpu/a0lTe6cs/obk7nfgGPW5j4krL
YmyWGqDD+hy8vIFitMqh3g2zYFJfgkExifByfI+dO/MNpUYkvIdgMEvA4eBnL9OW
K+zwF3Yi6O/JOuOphLU8Eq70N3aaQKVUCtH0lFah8U3oUJLvXyQkR0ElxiJlocCF
XHPlcTyhO2Tp3GXQb8qZExVBwyS4XYXC6jhCXow+5wEutethuFPwZ8rwKr5N1mJQ
mq5Czw6rrugQ1NCs6Pv6PP9jAjyWmb6Q5WdZIAc3icsqdGT3HjFJsuXIoCN7lTeA
oOf/6wj1K1554gCJt4ndwdOOKyKe1P8lDifK5v1c3hylz7sXh6s+yeDRlq42ophp
BoCd9avxqiKizowN8MxWaf3r2AB4LTwTtzP8LCVuRbszTmx79ewDfySSMybEfm+M
u2QRH4fMnOHAP0k7vz6Sc4kJmJLwIgfz+5hJTKQG/bTEWtS32cVOJFNAZVP9uysV
sLYUmt9rpIIZ7n2/MuwyDBJYSc6SAOw4crWPwM+np6uaaEX958ZHro+erZ8gTB/G
ASjNAZoc3yWv70hPOwJBZiBrved+gqJQO15PFQf7BS1SDlatn5PuteS7F5kXK7Po
UiS5GpGZseqLmvWKA8hk1bTr7y7vpyqUvGOiHz4No+dJgnp1SDu5rW6gVykETgYq
L+Z3z2p1Liv98mrRyVd27jJoOdCCgcapDtjqLHg6L+/AzK1SZTD/6FYBY965CnBL
uJjtrRlamwF/8+lwn/pvvRur5g7iV26Hf3csglleZaM=
`pragma protect end_protected

//pragma protect end
