//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2023 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = tinyml_accelerator
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Fri Jul 21 09:19:24 2023
// ***************************************************************************************

`define IP_UUID _4ebc5de730f9a250446a9920a5a21a9e03a697ff
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)

`include "defines.v"

module tinyml_accelerator #(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 5,
    parameter                       ADD_MODE                        = `ADD_MODE,
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,
    parameter                       MUL_MODE                        = `MUL_MODE,
    parameter                       FC_MODE                         = `FC_MODE,
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    //Convolution & Depthwise Convolution OP Parameter          
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,        
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,        
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,        
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    //FC OP Parameter         
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,  
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE      
)
(
//Global Signals
input                           clk,
input                           rstn,
//Custom Instruction
//--Command Interface
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
//--Response Interface
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
//DMA Master AXI4 Bus Interface
input                           m_axi_clk,
input                           m_axi_rstn,
//DMA Master AXI4 Write Bus Interface
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
//DMA Master AXI4 Read Bus Interface
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);

`IP_MODULE_NAME(tinyml_accelerator_int) #(
    .AXI_DW                          (AXI_DW),
    .OP_CNT                          (OP_CNT),
    .ADD_MODE                        (ADD_MODE),
    .MIN_MAX_MODE                    (MIN_MAX_MODE),
    .MUL_MODE                        (MUL_MODE),
    .FC_MODE                         (FC_MODE),
    .TINYML_CACHE                    (TINYML_CACHE),
    .CACHE_DEPTH                     (CACHE_DEPTH),
    .CONV_DEPTHW_MODE                (CONV_DEPTHW_MODE),
    .CONV_DEPTHW_LITE_PARALLEL       (CONV_DEPTHW_LITE_PARALLEL),
    .CONV_DEPTHW_LITE_AW             (CONV_DEPTHW_LITE_AW),
    .CONV_DEPTHW_STD_IN_PARALLEL     (CONV_DEPTHW_STD_IN_PARALLEL),
    .CONV_DEPTHW_STD_OUT_PARALLEL    (CONV_DEPTHW_STD_OUT_PARALLEL),
    .CONV_DEPTHW_STD_OUT_CH_FIFO_A   (CONV_DEPTHW_STD_OUT_CH_FIFO_A),
    .CONV_DEPTHW_STD_FILTER_FIFO_A   (CONV_DEPTHW_STD_FILTER_FIFO_A),
    .CONV_DEPTHW_STD_CNT_DTH         (CONV_DEPTHW_STD_CNT_DTH),
    .FC_MAX_IN_NODE                  (FC_MAX_IN_NODE),
    .FC_MAX_OUT_NODE                 (FC_MAX_OUT_NODE)
) u_tinyml_accelerator_int (
    .clk(clk),
    .rstn(rstn),
    .cmd_valid(cmd_valid),
    .cmd_function_id(cmd_function_id),
    .cmd_inputs_0(cmd_inputs_0),
    .cmd_inputs_1(cmd_inputs_1),
    .cmd_ready(cmd_ready),
    .cmd_int(cmd_int),
    .rsp_valid(rsp_valid),
    .rsp_outputs_0(rsp_outputs_0),
    .rsp_ready(rsp_ready),
    .m_axi_clk(m_axi_clk),
    .m_axi_rstn(m_axi_rstn),
    .m_axi_awvalid(m_axi_awvalid),
    .m_axi_awaddr(m_axi_awaddr),
    .m_axi_awlen(m_axi_awlen),
    .m_axi_awsize(m_axi_awsize),
    .m_axi_awburst(m_axi_awburst),
    .m_axi_awprot(m_axi_awprot),
    .m_axi_awlock(m_axi_awlock),
    .m_axi_awcache(m_axi_awcache),
    .m_axi_awready(m_axi_awready),
    .m_axi_wdata(m_axi_wdata),
    .m_axi_wstrb(m_axi_wstrb),
    .m_axi_wlast(m_axi_wlast),
    .m_axi_wvalid(m_axi_wvalid),
    .m_axi_wready(m_axi_wready),
    .m_axi_bresp(m_axi_bresp),
    .m_axi_bvalid(m_axi_bvalid),
    .m_axi_bready(m_axi_bready),
    .m_axi_arvalid(m_axi_arvalid),
    .m_axi_araddr(m_axi_araddr),
    .m_axi_arlen(m_axi_arlen),
    .m_axi_arsize(m_axi_arsize),
    .m_axi_arburst(m_axi_arburst),
    .m_axi_arprot(m_axi_arprot),
    .m_axi_arlock(m_axi_arlock),
    .m_axi_arcache(m_axi_arcache),
    .m_axi_arready(m_axi_arready),
    .m_axi_rvalid(m_axi_rvalid),
    .m_axi_rdata(m_axi_rdata),
    .m_axi_rlast(m_axi_rlast),
    .m_axi_rresp(m_axi_rresp),
    .m_axi_rready(m_axi_rready)
);

endmodule

`include "defines.v"
`timescale 1 ns / 1 ns
module `IP_MODULE_NAME(tinyml_accelerator_int) #(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 5,
    parameter                       ADD_MODE                        = `ADD_MODE,          
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,      
    parameter                       MUL_MODE                        = `MUL_MODE,         
    parameter                       FC_MODE                         = `FC_MODE,           
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE
)
(
input                           clk,
input                           rstn,
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
input                           m_axi_clk,
input                           m_axi_rstn,
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
C1DX8N1L/vJpqR3CcLUatSVnXeiSLPcEtObUDbLuEEJZboeVknqf54uc5YjESr08
JxwqDLuun4bh+HC7HKjher7s48+d9vqJr0aZc29VEV3RJBL/WYDDtXe7IMa/hM7R
Czw/UztZqq23vUlfULvMmxTcEhOoq8ay4pFgEIlds4Td3gF2nqY6i9ss1mjzsC/9
CsLKqo07YDi/osiIjZgrlPA/Yhm9Q3Ci+XCoW2hU5Sz8IlCv89Nwkqrj7BMupiHe
A4QP8LjgfEa/Vc5jHm1jJArAb420MAc/D3BSJ4/bckVRWTRMsBuGEgmLUEVlat0O
pCehwZzYs+lfE905iSd0/Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 51376 )
`pragma protect data_block
bzil+fgug+gKEGLd8KwwTXne4sINgzp7oM6Uj6TKQFx7YZTH9sJP73lCk7RcJ4i+
dro/D09O5ay57LSFRPmL0d8eUjbMatj3NgZ5Hvmvwv5mHsyPuLcFhTDkCFnqNSD3
Fkt8b0NhX+VI9im/6143Pgld+lGYbzl7/50/g8x+wDvx0WNBqfZHUzec498sbBfZ
r6rSqdW2Lim1/9fqzDDlb48xCr+XnOndRPC1DpOY5jrkfz4MYTmUCfqdUowj97vb
kMj4K1URNT1lE9caw8+pfWA6AIojN7/cOQoX45sSv1Iq5HPkG658t7/KzODU2fMr
FW8zyEvlaRbJ096pOhP9bRAQ6WO+sCREOecG8zboQkftJsNDqZBhG7n2E3rVETpz
Qbf7znfZdkWftb5/+rby6sXD0BGbPsLTwMgMeVopYUiy6rhgTtD18Os6ZDq3V1d5
yoDlDcRQcoo7bUjWw69s0G/XYaouBq1zbDeUi1J/YC5RDGBrTasa07BVAtbDgUg+
NdFuboy62Y2mo2tjqD8Ronqxa83+nWqc4KydR25qvYzfiEPLWvHcKn1B7syB+nLe
t1kFy9OCCoOuCzKp0Przww4ObQYE9zChfMSt9P0Npn87WvcDJp4zHIzoq7UE2oMN
4DH9yLtImDMSWI4AQAOiMeDxOzQMJJpNVgaVMAMcfsCV1GMnJM3rwwlIJ9KX22pO
MAqlVrqEGWeTP4U2hjYW8rujuq4rliV5K0cOcVPZqUXx5/4ac7cc18kVzWP3CMJl
JfczadM4xkLNlxqtFDBihcjuy1E5j28nE5H83+iiU4wBiy/bU3YP/+IrskDB0xVM
GyqWRAzStIdFeGZaiH4V2tuj0sC+9VwIGEiHOwvvlC2m6hK/Hkd+qTjJNxksuhC/
Zo06xGCFt/5BM8rRov3xw+kRVlbdA8Ma4pWvzjdMdVpU4s6bbsIDc1xRI+zoAjYY
o1YHYjaL4r6tNrBeLLgWG4KhFvuBP90XJL3zoaqNsHLbxMz/t41ymgTUESHww5vJ
xaGtz2wcNd8dumCLd0GKao7Wl21sgHGpKuSnsRw2kJAYfKB+ACEPs+F7GBJRjXd+
kcbuZmOuiGusU4IpZJFjwUlS0izCFlohKUKJXpfD69I9Ywyl7zZDfrEKy4zwMCKo
DcPo3KelXlqD2fD5SVjHniKT6V0YawOKY2SZgx9hLx4pYI7HsxFv29GueLF1Flmz
Huu/jsp/HBHyHqo/+8oZhMT6z3nPuJ95w72wr5QPo4AZ16W8DhoKLX9zUrUvhO8e
LFjODu3EFsl4OCEwd1TurXHTBYgduw/xHxS7HyLY1zuj8oiKsYVW16YZAr1ntphp
/uKBV6L+NY2ersHSQvz+EpRP8KMDcKDOFFwm7Je1m66u5ub7CkQt0zgs1NpNlASW
Kzg9xX6z6BTkG0bznuZgglNm57JHwe4tt1MN8Fkzkx19faohZue8CV1nRHtB3CXB
+NuycuFdK1Gz0aogpLL9ssHvEjR409KDAR9HF9Y7Bjjp+yEvKhcxlk61uWI4U4PM
wlSTspCSD3DTLsDkxvS/85i09PZeJzv5zc54Y8uaf72LtB989oz5PERRXGd03lrW
JbPPRf2dJ3QKe+zEBo+CLQcx8nBCESQtL0vjVHjhbZXj2NSa76u/IlLrT8+eVyr5
4t3fPuwxdm4/dbIbzw1YjKO1BJ4eb+2ZMs7t0rmDlpjhAFDc8D4tbBx+aofWjoc5
WfyJ58wbPZgkxLmOMFf8Q/DvglPNgKtPMGyribNnejrYKonFTTfvka9IpriOjmYO
8qTN49I/AjZm490FnR/wXr0p/znU7GmfufSx7whPfMSoajnNqMWkQuQphOH7QC5I
JcFUnplnAWy6EgrKrxTUbXxTxdKMnAsW1yN2WRY1jAfkRe2oYtHr+BodSwGO6GOA
t8ZuqGi6T2M75tv037VlGCSttK/ZotLXtxLDRW3x+ALJMnKW8FdUuQUPz+4FUDe2
+crxu/izR7oKz2arWf4PmqoTtfr5SkkMyaVMPcGjMwVLe5LHuQznTXfbx/tJlZyg
SVVWbwqyqnsfpIhAB1bt6YxkSsJ0FNKK5+AzcxWvWaeb7Z6D/x8Usn1d6kp4QJxh
cU878OaHCNQZ14QGVnfvKfq1CTMisL8cAfP7Gj0g7ufZ93ybUw6+N3KPXRicuNEU
gziAn54zyZUM4ngu+50O4w6xwjJbjcspNMtQfFPbMm3Krykq0lwwgXwMgHLf70Xt
yd574qrDoHF96IUbH+3e7+6aBr1VZ9xvzvsSrl1jxwOL32aOsgYRfqk7GBDFw5de
w4/497NYQ4essleDNE1tWPabgYR6qYrbJ1ujaYrCI2x9VG67YmI1tpgTHwNLUr/i
kUd4z8eBw57enMBr0K2yp7hUefWeKrpFsH1NqbDY10xay53Gio5LhEYKQqoW826q
gqTN2YF95yUy4U+9k7WRRF92KwqsLObGl0fgmhD2ZJyFuaDd4e/M42fUpsEDYaTd
5bC0pgEisHi5RuI+IO4PRqvlQ4heAvnZo10DUBKUkOFR23erHErT6GUvxKl8fzQG
vD2TnNckxxSWfIoU48vqaifJCXh54nDjIN+ezGMfP3Obu61C981X8pi52Q200oTa
C/yriD6mwwd4M10BKKDt5obuW6kfMuqMhYLX8LgT7fk8St1ZkY6l0vR0oYATmali
uSYgxO8qMDJmNqvWmzE6N8ibV5+70F1tCkGCbCn0TaKVjBZ2I0zzKdtPYOoVmBMt
vnKLgm956EHBc6RmjXhHAfouAD+rqvMnZM3FpzRWLeVB+0+Fu4W5LtIj69TDwoZu
eOjt0bOBpQP/2/gAkCL6DiCNmutqOQ/4mI9CjjAtri4jLYHAnZYw7vxYlHmuopbI
eo9bNPYNnXdAw8OkyXpvLOPeqC57wxXauqRwd6YXVXevBfYK5AH7/PZbz0tVizBf
Yg5ReMWM6UQ5Sqb/oxLqkko+BpMW2XOw/vuY37oSvtmwOPt2d+4C9TNPQ6FVIcey
LRyHoyg9R4HNM99i5uWfe7IEQ6ufJuhqcMIOdhczNUB8Yek0hBmz4TXxz4JizfYo
93RRcSCNL9QhtWwrvRBM6z86y8x3v7UMoEOeztOkIQSBCerHMNXva7TR03qqaXY/
XiIPu8uez/MNwE4zATqLB2QvIqvdJWih3NSiR/QgAvRnzvc/qcZsEXqkGDl9xy5h
jPVStzdE6WIfnz6HiV37UKWyHKtgIXl9GFvXQjkfvOWThh5wsv62SeUAorGntsJu
6HoMsE5RQaGMJE7PXRAcXNV9Ryu0FIVsyWsVUeCPDCduATKV/ogaAfRXjrQjkyMv
DoL5JswbDF/NS7VoXnJ+rTezz0usDOK3Xb7shf+le2CZplPkd1muZcEiUU9xyoE0
Rb9OacK6SJjukkXCBCkEnyVwk1i89KCRzcuoJ+EE8MugcubRrQr6cJCEuSSAyM48
YVavP7Nc4TZh2+Z3PouNYiSWEMM6vrb1ALv03iYHQjd/4x7DxhwjMbdgRhZG4kHe
0KXVlYdv99O3kSgJnxsQ8i9uxQwjAJw19IJPFVTXIzAo1RMsgco4TLQm/zhJlnPG
khQ1UqjMJBBGyC0mctOrH1n4JgDX6T0r7l3X9dv98x5VtBZlrXaX2uNyjBC/+q0F
TzWY9rjKNkdbrAwXVtipRz3TTVv1YlNYtqMiS4WjyvBnHmH4VT/qn6+GqU2tnWZE
K+zQybDllGxltKLt1IQYrNoWY3t8H9lTJRtT3N+iJa452XfC3Uzwsb2jK3X0cMmm
0VSs37BRt3HN7sQlciRvDShga7vqRmGANRw3Sf8V6DEh/7T4OGDmxqssscuaisOt
mx8uFjITI5rcmot63ZumzHFjg+ixt5EYjP6Z2eF3BiqV9uTx5A8a72xyPZU6grDy
be3J4Hh3bSEl2d4a4SxPRMvATZB4IIfhv9AHIeNqjQTKNGCmwOR8jKdrqvi9syvC
f1FDe09/5LRddYaJgNW5YkzUfAYFKpy6xD6/5CQzV5U0yj+OV5OVto9t+31kTSUS
SrWfY2q/2PojMQQyZy2p9xvOXq3Xh1lLfbKPU9V3ydf7KRKR7tSqISRtJXBaxFRZ
JB1b7ht5uhW0pIt0Tm0F7CJP81piCLYNllvbOoMGa/mmAowV/J4xcSg1PxD77ioE
Ftj8qtUi6EDznm2ylMxpTsS2kb71aFp8lgxbHoVFHjATchhQBQH5Jp/QRVmKwTFb
bN441u/ApGEDufn+138GBNA0y8VrPXJJINxZZtptvMFBNEJKDasDpqHifFMgvFQO
lTcQFO2nOeBU2Xc7/0gmur9rhV53tugzAqPksf1ZCPh3bLxMjWsaT5LA25EqtXnE
tZT9T8/HJ83pxTJ5BaEz0L92OUUYPiqyGLclYDYD12db7gQMkTHD9kBR6Z9YM3En
0GHIro3hcjKBq12LOT0S11a2SqfwZGnt5Qzi59Y+0evUR3Dntzap5VItXPGFQQrW
s6XWfVxIZXpG/nXXvEeNzYccKJlnT09BgoeuXTofYsdrhu6S45+aAboeS/OWe76K
zA+5F4axq0/Di3O3VgySRQ5Lmx/thv+lDZRs4fJV3Jj8YVq2L057AquSGGUOO16T
8yAAmtyTCvlBODJkWWSzJqMYla6F4h0ITSs8Ouaztov7n0LnD4q10ev8pYh5gPWv
NI93bZcEAHTsh2jM3OtydQTUZN3MqFzmtZpggvChw8dBS9mlWYg+ZeeI42+jwfXf
xbalYpl8BWS1ABT2SEr/KCVQl2ahaRdHNnVJSwJq3eZovF85FZyB3vyXPbueViAg
9Db5+GV82rMBnw8qM1c3vBl5qrqaWgaJ5bT+9FXeFesr8zjdsjRK1VpCzBYY9cKJ
fCPC8+9rP+lwVoBFGdBvIJs54cvKvW3zmBBADLinZ9HK5hYFWzg13y4gFk10SnDu
FBLqewkjIMduey1Ei4ZrFtd4IvU22AFvyvwEjMlxbwk4IuYza862Xff8ZiPaEEXf
V9cMDtGKh/eXFzeRROa+9+Ny7qLefYjCocRWBMiVafQSZMwsE6tN+BssJpuNLpVM
cTIJSAt3NYgSIFeoEnHWnmpSGls9Fv2RYW4NBWY9k4Ql50moqF1ZORhoecuxXvNr
RVIhONSQRn/5ipNaR1Z2tItIntPDGi2zZGWK/zgxGFsDLb6WDWT9TK75ab+CxLZe
Nj5Uf5rbtWErdFQB2vesQNM00sAgFmYtHqQqnh7v8tqNdRZ76ftdE7vSvH1o9Lwi
JqUnEgq01BE/MnYGCMPrGpobWl+hR4FeI2JzX5LB4NlEoBmiHfcclFfaeyCFxUZv
AYDcPA274lfqaB8aZ5P9SVZJD0INlgRwKOo5nuAR8JWFq+j8t5Li6iymL0sNW/1D
es2vYbOIMAwboNarHgbLk8zAV+IdWSZDEA7mO5tt6bWPfarFTWPFCyt8EL9Dvc9i
0OTEezmidpGAfcIzowZ3aFI4YJ/KA9tJ1IyagNM4GsywlSiLk9EM3imTayTAQoex
rkQibl1x5vfj47s70vqWT1FbfXN/WiAKnUKWRcR5wCkNJ1G8/vXMTSYF2ucMZWd+
RXg1Y0yuTjh7ysVu6dzzXCYKIJCgZ5AN4UNmAc6coRLkMPbf2JBxlaRNmk4EbEet
AW6dAsk18Zstkrg2WomkV3oTpARTqONtaZeEmKuA0plENzXAyj7O5Sjl/Dqt4oPi
EbBoe9zs5So1RCxMg+rb9G2U33B6d0WEJnrVR5UxeUqHzQ8kQ2Zq3Om89DXskzD8
nheXNy6/g5UMF6urk0f6zSPs9JMOCugptxQz9J6OyFI7IBUsymeaRpz6L3+mAv6E
Z8A1k4/C5rtPlGHIDhg5huQikd8LzeiIe5nXpZw9hVbsbn/kW5zG1gQMyDmYGMUN
no0ZHiaAhjIJqasZaq7GieY2XYk4gVhsJ54pcl0kL6BBR43I51NakYK1oiWV643J
YSkdneeeELVBzDcQeV0icUm3kBrrnUWErKvdH53u+2ijypc03nYmJUL9KEsmUjHn
zrW8P2QW68JY2on3OL82+mWjAlzD6W9IquXqLZ7hbdfYc/hVVLTf7kZKq5DFt7BJ
O+qoU8CLFwHklutClkjWRVaOJwrJijkEB5dH14ShcAWIpCfAZgDi3OI3hhLFPsbm
jMs4UpM4KbTJk4fkoPK1DZaOyoqe5HxY/J2AYCuUvwCgK9vvEu1EINU2cuyAD6d2
NIi5RkGaf2l2PfJk9ccs+Q7yKGJ6mbiSX8qyZTnQH/aofht2cQzgMXl3e5Lo8N1h
JY5L//wrt35IaCtY30WVS/DlluV5rFXzMlfddyOezWJ4HMC0RVYIp0BYB9g8lgLE
x7jNmwOWP/SuzRMaYi3gxLQJiffh03JnSUvZktqK+HvpVEd2Lb08z4W6e7V9Og7G
bQEh6J784vjSkb/UiKbFeo9dQvJhJNa5fpoTucirbgMtvd7I9yXhlTtUyZ3HBhqL
l8jtArPSvw3XlYjhs5KxqQLyi5b2H05AxqH6HgYxVpceJVQ0NNYpNZllQLnu/NFs
2JM2XrBdURy2lFjm4IX6KTMgIuxY8Z63OeC8MGBsEezSPvsYACOM0qc+VicmmEbT
TOskKZXKKbp5ZObL5BI/1ksGlPsooe9/OVkmW9bATnrV6pmyWK9dGXDpma4Cdhkx
XC2UH4BhRGL+G6+wrBG6hI+L0hAn+b3sfSj0S4lfAVYNZ+br+GHLDtyXPvLHVGQy
a6ZrWPFPPFhWa20erc8yXWu4Mv8NiDE0/wZmlmw/MfVSLaHl8ha6wkFKuf3TCA8r
9PDGIVjD27Pai8s59HHUAKk+8epKyqyGVe8E+IfqM054eOeRnkrfCKx2hbhSnnPt
1l9gvPJs8c51cZn1P+6WC0AvdBhNHzcLBK5Igv2NQGsopWpBBuHPQEtD8y/XRyuA
ewpYeX3ytggksNKwxVdwCDJWU9O0qIa4+CQnUlLGkcYK42FEQ39w5wUicQQrlNlt
5Wh8IWjwJAi9wfC/70e/p68BZjRBaxHkZb38VS4xJGL4fbgBGNmox/fdCAYVMY1C
mIFh4LEceblUJaMkEZrGhoGFBELVIYUN6iZFRz65li0L6SeNo5Bh3ORJ4keZAHyD
mEeCl5u5CbEaOjS8M7hU6uSohEWqjxsUz+zygmMB5eU942FOUhLWZX3TzALTgUYd
60xy/HUM2IrQGC+JXdnVQMVwbvVO5z6JCzymiFkNy+PKlNTJW+4fG40E7i/9+KtI
ZyO4V64PPCAywFl9k35GfhVlBB+NMKhRuq/mf5rTYqMkozZ0jFpPYdjVZSTMbkfK
fXN8MBjdANWzgm1lk8F7HPsSN18PFSoaU/UpI2VpkKrO+JJ3i0GZi6ejecBgpMd0
zpUPf1N73SefwmOj9mPC83xuqgDGKmutOjE+olN8C6NVMnNhrmVGEkoq0y6Kt8Kx
wsDZnkksKPhTp8hw9KA1PGkgMEWcqHUchcP7O+qv4OpkkPWoMEpWKH7ZVrtRnUHX
RAHlY4+2/tGkFXyDShJrclYlPpmZQ9Al784bG3+Yl6DuooLQLdBi3gzh0VzTv/xX
nyMWzOne6WXhKbE7Sk8MYHDzIjuxQGkpjXQDmwlPzAElJDv29yc6rWW3fxhX1DX6
AOwjFTj/jpY8lwXukO8lCaKwhT4VF4YCn+90Fsw71XqXZ3sdUdMaSnn91GheLW8X
MPL6WN4aBZgG1G8itho5fDEPoHCh4sc3LG5L+I5vXk+pnm4a1XPYaswdAkC6nuOQ
P93hHKhiDMeqPpaTXjBhLiCsfNFUdiqYNGyGf+9L6yt+exSA/RdSNtGYHB6qq/xw
57wJi8koeQeN2mP5xpLvas7MJa5Og9TtiVC1TdBE7iLFpAXE3yEImzRQa8O3v0BF
lI8i7squcQRmadm5Ejyojo2HizbX7gposSB/ASCdYKT8ggrnysj4z6QyuYY9S8c3
tuqEhLNymOUKEueebWjLZAFECtBo+FWY+10S2NgcH7VVBlhxECyKhsLK5/kVSgfD
k7n16uQtSE7O13fS1dHmpDhklo/F5xBED0rGT8/t6c5X3Uq5oE8BTEx39oCXJF9X
OrH+JDMgLHSC49F8M4ad3r7CPIdE2qXdep7HQbmPL5BfdFqhwRNz+E7k++NwRpZm
vAw9XC28pnZlqsAwzUedCGJ95jqvvY8c3MQnmgwQi7swo+n+jkr8TKPhDE1TrjPK
dYexjf/vhGH0HsMdl7GNiftCJmLC+EvJvSCyiZd2IdBasGGwRHqf6t3riVyNqaHc
i4TE0PShOwIX9PIGM5kffxZKRauAoXZbBOerA9nhimGu6aGBEyjVUPIBLk3SefG2
xbhCLA3oUejHfxy9y8GmgirPz3oQo18mwilXy9Y8RH/q65bUKs2gEc2i/jG2L6If
QZp5K1FRsmVXZESpPwpovMErQlQ4Sb2vwdSOBLizhA3xgdM3MLIv2CgknTCRYl2+
BlBoDjzm0IO/n5csifa60AD/pyH0ToZWcYiZ/uCUvJNIrRWnQ3IDpSMDkTWt44Ex
u1+qsJjVtz+7PZfL2sFwIKz0ii+JKUtdDvrPrsGzhAxDfDpvdYBrgYkhX5ukNyyv
XiJtYuD9j3n2yy4BuQM/GFdws9kGAt/UcTCltVMy4wI5ktHOMoEjeq+UvM2vy4jC
2JeqCo7aCUV4Ne+Ozy8vtnRE3lr8PA1gioFNUzoOnzXKZKw1kZpFVomUAJqOgjQE
QTwf6PUB3xFFbLYkDrXwqASQ5KgOoSoL2DbBpAzGP/IXkThtmQwDetWvc4oYOa/D
NSElJceBY/blVhIo6LaeWytb24vp6pOnSA1/02q2w+3+9W0ontgxwcJuLnBrAC1E
XHR0szUZPwyEMC9gzouzIZUYGUwbY3q9NZ8njp0vOsAYyk6EvNRJgJ34AFq4UNtA
2RtCPh9ThgroJcN+5esqU+Vw90VJDP5pVLGAL2MZQJ/lNdtu01b3aOBXSw+VqAvA
roujH4xBZ5y8nXwNgAVnJazC0wM0OEOpsQpKhoAk8mHDntQwD0L7/mjcDuTV8lin
jkjDhWwtkR/uRqF0cyxfY4N/beLCat/dJZMwnLlW2kdZHP0q83ZPxrGW4L1Bt/23
gUL5fs42x4hayXwKudLbZzYx6q2BIO/G79Kktzd5nsb3KFF6YiByLLVhl1X0f/nE
GZi3hPXuREtDrMArwalxSdLKafcixwxIp4NnrbnaEqrQMuCZTL6KVIhq4h5fjUSe
+b2l8WLgd0VXdJTxCqtdQi2ejUEKT6pt+gsKNY3MapAnqA9tK2kdeSEAMoGR+NrK
6E9ORJ6AlhZ4XGdpYWJHoxpSBdRMW163vekIgcdKaBxP4JrIHCI+2JkAhokYDGQT
HYg/dFnTRQGwzoccAOLgDLBPUWAURo76BSgHabcM6gzwc0M0+hpnC0STIkiHFPy3
j9CIvXoWNvXWyRrJdC5SFt9Rksvzs+bh3wpWEGm+Do2wCuxzFXZa0zEMq2E4eSPx
Py8o/j61Hn4uyOVmqHR9GjYM1IowihNtrj6ZMbI5hJsrie7tN3lHfFZmuvN4V5fs
x3+WslNA7NQ6nuFChKfGmrk/aaV94Qk9AQR6YL5ON7Ztzay2r3sBUr8R/YHEmoc7
x4lzXlabX6jxC30iEr7T07mL1cUMxFfvAig7UlC/k2o0kvIih/gw9LRGC9IS7GPA
ccNGpllEMzMUzo9c/qzpLvn3J/CPT4GtlDb4f1a8wQbXEGLu05m7IQE/GSEmO+vg
hYN/FVzknK+oJwX9H8TFQ9vcSQlALMwP3Hv4q3zvD1gt9ioVoaN6fwrfV55iKXrg
fgB24foKHUFCLV0mzDcrcqmygBBwjqbwLtD36vBpkqwOBtVwEA37xbIb2s5Zor+G
kvK/Hxp+YaBinnAKcrnSF8x+iwTn2ngruPu8h/WusenApU83+kH62Q9iA6XJluZq
53SQa24JUacscFKu5JI96WPOQkivI2R7EKtcyhln1p5YIMSjxc5C2qDJ2pIlUYA/
xDFJ0ftRacLy8+/FXkuinwwvadmBTvvvnlUM/xo9yMkvZDCiuV0hR3FbDjIyM8QK
FrMVOUHQpQkqNX8nM2cngVV95xcbF9p287NCGlEjJ6Gbvpw2cDWnFO6I2QUruBfY
Zz3fhVXQ8yyGmtb/9u51DNsNOfy0s6j7fvV97sOUWXQWAvpuH/hS2NIZXD0+Gwo4
zbhk66Lxa2juyVfRqyhQsy4mKRW6QlajisUDRhY9jaq6sUj3axCesgXM4E3i+/nO
L9953YFg/wMYes5J1kuV/5SkmMa2L1Gfw7zxuotzKwi/2IcUaD3R1ObhuGJdBtgP
CKGKpd40PdCWRAxBaYHfXYcghvhBs931E2kC1Ir1THvVU7wk4IMjewSjnoxodQRP
DrNhacXhxb46XZuwA3XGXe54Hg5QZyVDvJ/dUEL1KpTZeMSpypKr3Pyrx/EncSqi
hDhlS5IzAtZUQfoweDI9R/buOJtOnzFj3+7rJduZe0ZuPDLpVXIpX8VmJRvSuNgp
GKDAqTKDon21leF0XSLEwF/AgNR6quYQpgdJGyaX37wZgmLWix7q/FLQhOxUcVXP
+wOer4H9wHs7YSjh1AoqyhOuSAiFKHOxouR4wLzJ3kefRFkcvq6ayuqOtDRfraof
esvYrplpvXlkIR61ejwFMCGs1/Dm3cySWVY6UhUGZHyXsW2mhmsCgHWMv4PQxTzp
RPu4UGMc9V/aVgRKIEJuKOZIxHlpJbFe5RMAa9/paNpTUoMLQRmBOpVeQrv0Guud
3KiY9wN3NI5OQHwgM6Gf9ELb0YhOpCv9+i0HFc3s9t0Fj89ci0pWVhu89Pv6txUf
kXsSZYey7hR+5Ol9q7BX8FInZgywKnR/ddr0wIfLVAYOyu41pTSJk7I0GX9GWMl7
kJYyHGwmEpIm1hpmaSq6+ikSusyDAZxtLoKuI4lhTtwftXAHK4JGCaaL2vYrH3q+
3w8F949iE1OK1b3qkr/U/MOwRzyoaaJQ5UIEbFAUvyFHPQpq4TcXH/BefdfEM+LN
X7QM5ZGsfbcxP5Oryke8Fw62RY/6xnz+052IzYpjWN3TGLWquaqPw0Mox1BglT7F
ssQP26NONzZ4Ucu2wpT7K7ltZDYbFAVwUs0Gp7OjEuQipRBbJQVYgOnckXqGeD2j
KGGgSmDyN6Zlo2KtxRL3HoK/ZRgeBL64QhH4kD0N7VBZ6TcKXeYRD5RP8wEQlPKa
M/VXOYqdNklxc8l266UhJx//K7Vy0EscbwBUdoV/w5CcpPXAUji7SHtJq3pqvASi
c5LIdX4UW8AvMcLyGCMkfdqVsIGtfp8DjNDYOQ13OCuPmFvpFqeErwzLXckk45uR
ZIr2IVtNDC+fhtdsXnswW318gX0AheBZCEgBDxAmB3rxBZVqv0qzlbX+KabrxnD4
kNPTfBDwWak4X2fxTlOJgegGn3r+pyKaatJRd35CQRCKZVg0v9wSMtGvNZVWPiut
c1EJ7IDKL2HMFVmNv79AcuUo7aXLUsxO6rcZPH9qgm+JpL4Xy0dLY7vhjL4hLzP8
ctgtEth02HY1JWgrtkY92vsrXBRm0S2mYd+p+8NKjHN604GzDb4/l6KV9glX7jG8
VO+TjK37X56LcI/pIarsQKk8KbxwlDjbwdFSOmsH/EXTkVyAkalW7Q8bjTp9M/Ir
+sgDXqPhoVHFdfygF7CC83zZjO1gCqWjh3iTp+wfiJ+0MiFWRAcBNlPT3b1VSfmM
hoWXj0VViDPBcgjrO717EOUZPG25JYjiwAbAmT7dZ1n78MoEy1scghH5VTBCiiQh
sF9FqwUqCOeDIsjVX6M4GY+T71aMybqqEkB9QCRn+QB5Co0UM1QiFZcsyB+L4kFD
ophP1Dje8NASOEnTn59Jv6ESc3nirGcqvBJNN6vXqTv4cMSqP69Ac2yQx6yqT8YT
6JzyjijXEdw3nPj3SO3ybnluFmV+kJHg8kyYXGXEENBjG59jM2JVTo3zvycdY3ym
DG5r66Cy6mL1qbeYm2lB87FL/HhokhUFEOmEvsvO14kUs+PPqq7Vw8UJNOqqkJgk
rgEEA03OUXijmkO7dTSdgZupK820Ycp1Uoe6yCFwNwI7cEtk+ClUIqyoG8Ba/eM/
CQMoXuWBfDf45lh5hdkIPbD92A1J7HRcMi+VWrZX6ydIF20J90afOof6M6Sblv/7
6x4HiGSGNYTZI3lzxdatZZPdkGsEz8mOQ/XrsN+jz6bU0C+dQwsHL6Fvrtv8SVx+
chl6Wlgwa+pqbA6nvNvPsAS5YAKtfIFkS7gEcyggm/XDVbI4y15lUd9mwr0IXJ95
FT6NXl4qwqvTxptabS7pkSvGxLv58G2N25uCrw/68i/5QxZMGVhs4T0g6g31/HFB
rxMFXalSze6OkvXbE9rjrFltG0Eot2lonnoN9h6wOgYtmfope8xPYgdTw2ORmdQc
/SF+BbOm6ZebWRaDhFhrscuTMt6b14rkkJHRlyKtmHiTiTIsHoveIv2x9bhk1nxp
DvUAQLzcMIMaPPo/PPwfo2E3GsULqh30j3VLTVCLAz0DOSR/lmvdVjR/d48sr5WL
eoYql4L/YmaAvYRjTl4/4jpXNMrgPglNbR2sHcqpCBZkTt/NJ0WX0pEsvw/I5UsS
WI21ckC5SGOmrLQmqCiRdnECHe+iQJcd1konifQzER0XC3HZ3A2SeDxs3tn/hMR7
3QxJ50OKZjGGlCc6Eck0NjkodELdxSmyLW2ciLhfsKPSK+P0dxKItheN7gp+XEF4
U9pK+PBEE8Dw8mJ0p1nye5GUC+XGQ3/vMWNzV3uw+WSwuilJdasR0GKfya6sr9pn
f2PDmt9xoq/nvLHWqH6a8QjTRhwQLtIpYfvPbqFH0N9saAUwZi0/R7skVMyN1vr0
LKBvFbV1NIceKy9PmwqjAJps3OxUckbDWa/+ijj28tuFksEr7C5hOnm4wheXhgm5
fVKS+OquxgB3515/zUY8ncskBb+PS6qi/NTUFxbLh1o1mAVOeMibknLI90KQpJTD
A2LL8wFbLGc7Rgl0QeVjrT6rINdah/bK9dYuGMoWs1EYIdcnFySyGSzJcNFVnqS5
S32relnqQ2JKwvI61HBdIi5Wwdj288YahEDjkRxMSEHGD3AgfJjwg0cTks9lOsk8
8+K/zPbN4+WoDxrr7oJLnO35Bh39HfwlFkbkIZ66P1bhdl+ljN+kNufuyvsxM7ff
hk6S6RLbpOIsn8dR0fsVuTVfzACdSR5uzqo1MLWh0YBPmi6r0u23nkvA9malULGS
/UgxCLTzy//PqqIdT4/Twoi3UZPEcQgs833+92W/0KqHLSznqFEOppkf+g1VEknF
hfqsqh4OkgKMYlNCOEtms4OYjoLDxjXcOAOXCTV8HhElVPwIqonEoYqHCqfbePxs
LWc6qksPILU+e4twPHYUDR3kzITOCyyTz2FOJpvFgP0gdfVElVqvKu8xVrwwdTQD
WPkoVfWWcS3XdJUnd9+9rpN1pchtRPC39mZIUa0eBOUroOfVdPTwN8+kbd6bo6lc
iUeae2LIZEf3yLUPdW4yc4CxxGDV1P2KSfOTsds1dwKhLebKKEnw0V0gUrSlzM3V
xJznDOAo1rJPf8vwYI1eNBBsmlBOYXnxXb4db1gGoladzEQMOkt0kItdxZ/AvNWU
D03b/0Lb8SPU0zzSsH523Wjz6A1uoUOTgRyBU8jln09YvLScH3cSzYI0Gx0jApc0
p4vInVOd1YReMz7G12zfOWHkDEFKEa1J0uLMLzsYmmuTigRDHRwM8Ynm+riYdB4p
iRIOr8aHa7aBsTobhMYQ5aaER48aTO0+7pOjZMNkbzLU693s3lG5R2IM6MJgM1El
FT9sGbDv/gycdsekTwAUq2CU75EOZNWd9yQvtdWsrRft1GPjryG1zmdZRMDg/qGd
EM9h988RolHyQC/3fzL+M4gp/wloXKVCnz4tN6oAzifL5up2kw8bq0aQcA3roQtS
Jn+sHOYz4gOmEePD9+b3wJh3D2D9YNW0gc7vI3IYCPN8OeIJXsurulPZXjb7JsXq
QjyICSO4yx0C482QPSKQJySI7/xuDxChWeTrKY31uJCpBa48KxNOJ4PCvVdUhs+J
Cdj/isOPIf8C748R4svBZQrtJ6BzdrIDC5hapUea2isWJuv0IDokWQUgjCXqD5Mp
OxmE1EG+WOHjspWkatcWWD5k5QArN0dFHaakkffz10w3UV0xzolvd+frMiOqLyyE
7At2oh2NtfgmD8FiwVAqMqwgKo3Ix7bs+VXWIt71/wTXOIRk2LV+4UktYCeU6KHY
Ohk4a5/w/e8MHPX/8GUwcOKQ/2w9o1aEUQeWs7xbsFZwuZUToa/Jlh0uMVwHa1kP
G9AGPvbtWyV95oiEg7IkNcMVOXW1p1+y/vTBRem7il43a2dbvKAX9KR/7FZF3P+/
/ZyXXlffSzcx6QvfR5yOm96pEnR8fexZvkBxeUJ0S/CLZMFJQcSa8AOtYa+1SdHV
IF3o4V79zDYXOLpNNVH4yzZGP29fZLJdSVxYEib4c4ERGOzEOpnJB7Ya1ZRw3xCe
5v6cTrCfP2mdDnUjAM8FyVJkV8KHFy3bloyF35aHtG09JZFspSBkhgGcjncDgsXo
o/B9qrp4Tpg59Tsp0YmF2rgqbUv8ru8nm3rqGvUK53PGhU+9qXKTfW531sQloKhL
pOe93HZRWnkTG/nA/6SqlcyoAQC/9sU9wx5nbA3rGvGpPF7XcMZM2mHL67HPnMfe
SX0yEqaM9ZSvZJOHP6gAB1NDIglz+nN1xPCFgegKMUVAik+KOzn9JCo9+9T39fdy
NDTj9pUv12cuKmznHdj8ejEv6LTjT5w3UsWW8/8w5sm3Hxt788Y9k4DbzabDd5ge
qoIV35Mshb6h+ZZBdworF7UnrVtBq5ZH7C8Y6SdOfkH4uQCDp1uS9m8YCiBn0Qzx
B/Ya2r8hBBHPzh1clnXQK6XmfDqpz4cmLYAWHRPQ4D1++B2mBbCP9+rKE2ZKBQNu
820FJrOrZbngv3ie18p5wZYIzNHoUuDJE34ocJ7RNAoV39VZ+nglBa5QH+GPo5SQ
yfAI6+VmKcTP204l9T0fJrocfbNKPf1MGKz3oZ6CqrdFZZnPz9NHuxTx+dG1+KGC
hxOyea1wRwSU54jHmA9JPUuBNBZDniUS2vta5YwVKgYkW3TJMy+kaPKA29LXKvX9
Wzpmmo7irippUUswosbuEbnU1VP/seJZQj/YRZ4EP7XsPLgmztkGvlv4FOQY3sKU
8kajhUQPSG2Gmtau4Vq+mmmIfBnkkGzusVY8mZBhCmx5jTwW7ioQTdsI/XToTLtj
pPm5dIMnkfDeChUMF9szFnN9Mq+9TfQcJViYAliA/UcURzrUAs3ufq/V+xdwTPYf
+YK4w26w/IXUslFc0KYymGbj0qHREoITP0bSni5/SnDB6xHFb/zTf0LNzurbYil5
3wzy1C6usDrjLK24PgLgDr3TiNarXyNvwnc+Uu9gVxxcvPzn3d3PtM76cWVlMoqJ
XSgOjLuQ8k4UWCbQ8pOcM9JsFExD0OAi/eC00zdUUhqBI3ERNU2fNFWaEKZp2HAp
scrdepaBks5/7Jfsr5/dEX/o2GTfNVFz8IEe3M767lrruwidzIAMQ1824r0uWV/2
v7pHqVorNGwq5Q/LJZNJKYMMXwgl/mcBpCfJpB64tq0w103dnO+uSOjiAq5ei+dj
NKMVln3N2SXv1l5P4XlvPCLsVaGI5yIcOLugrnp65gpzksKg/w0oLGprBhWw6UH/
MVIDfsJ/MI78/JGav38FtcCpVSH8T2VJKwiAZ0ofyFvof0nYkXs0rzPpuM/SLD9K
uJd6Or2gd4YDnjMpShhsEYJuue7jEH7kkEM+ZiRjOSXitYYqOtfpOgZtRY4BaV1+
KKOnGQxmx31/8eZflzyV8obcHt4zhGZSBwa4FXc9iTYITD/HPr63bmzHAYIipXnO
haJI+smjJG2yB2LqcvD47hBexqohJ4oSyGG2tFGqEPGsVg2SUSpVT5jOrkmp1YKN
Ix4HcZb3JbvyjDT3kbl9bj8eQvBdWxQIUkhPkTcepk5ZCQVbuW1D8Au3sisKqsy+
henmV9Ct6SGWMCZpqFIpDFcEzOwn5Ptv7Ul2btI87N8/PSeigKQR3SJvK+U4Xk0s
dZ5lDIPzwsY4GOsbAlOstcccfdihtYt8rkXQjgT1bwZuYKAbT6knPoHPphoNDfDG
6kC7S8aO3f3+za7T8gP1QJKbYBnOEQRxWJ6UO/LH+aKLYx4z/M3n68U2gZl8IQZN
MJgRJT0HSr+I65n6vpeXC6m33fXBncR8sibnqQMW6EtkiqmMZbwF0E2VAISi2sBj
N5oDBwyPg9tRpihjYj4KLV/jJ4UIQiZHZmJx388AhXCKEyrMy+7KQOd0VlQtG7ur
zbkn4JgdDBP8LcPi/+OmaYxmU7hmrDDpBNXsjdKb2RjQpH2IgSjfTqfAES/83p8k
S3OjLDnXT9yOrfuhf0UqzUUNVJ8tNE6gWjYy/8aZ0fAsR+0ikCig2Iyiaegd6Jrx
q2GtSbpeKlXT+s9ltBmBk8yOWt/RpWQK2RTe+fyMTq0OL34/AGW6lEpMJdXXZA+8
ZPAROjfVcXC4y2Z6rxqB23MXh0dTEZnSlyMSm1rXPDVqm9E2RJV6G/Pp+9obPbnF
M4RFGXS9zbktGR+fw+Fhyi/f3ijhK9UjD98V//QJt6ESuKdR06nRRB7PebglhrAu
RZUTydASVwbS3Lr8GXyjTGfm3UhmYVGj+WXkdmClppY+AYKctx6iHIDzhLmyYjin
rYmftqkBZv/gWVQidT5GzxwhIZ01tuKqFW0BxGrPrZtRAO3fWdXMGRcUDCiK9yLY
oZhBGAimqddpOs79ltTntc64JcuOSUP1wt8krj6DcYR15F/+nyVQPXNEj+OZFogC
jB1n4knsqnVD64nI8QvvWasRH1+QLspfV00gCsExQEBqRrDbMnZN9sf8qamkfvNl
g5rsWGhpyqqZ0o1Quw6SuCgMpCVkpZlUWQsrQAXTcVH1Ee4RrRfIz/IjQN/SPuNz
svjiQgpU+4hfOK+hmEyRkWSYr/w9iLmDCtFjpe8Ui0c/6AfudtswYHNVCsgLk0Pb
a0ix5n7rxP6oDxv+xeUboDwtUmvC6u6TVjyhK3ImpJTOL6DIAWTy/EfjceKSqngh
qICjqmnAPSuwtPKgslmnr8WqVKBcB3WZZFmQxRI6zy8BRYP1UQ/YMY8YxcYPwqpy
Ox8TVT5TBrOmr9I2iAr5r2SXmBsSVGI05MYmMyQ4TwvRN8mz+sLn4FZsX5PTWpYa
nPEeDyszSFq7xDq0RBHT2qYyEDQoicJGUxKpmfq1kjBrVEJOIT0/5Bj3cwT4vARQ
OThgSXeUfaXNVeDLwFhV8+DAuHa+UHapGGV3n4uW1F5o3K+xeheSQPWc0oHowy0G
utGtkJ1xGQgOd6KLACGPp1nEvER1o+RvnftZnP2XW7XnN7x+opvUKSz1TTM+6a55
6TOGlzutKgNUpTGNEZmo9tAtshODKxSjbRK7BINI7vNfms2NoD26SxTuMJRfMWsK
7/N/XBB5bnIE59kKbmFpWWYbRXMUaJZFMxHMEU8WonzPz/daETwISIkXkzutyysg
KK+lIEmax78yvZvaCz2Iu3FInw7Ufde91wuihGw2PACpwtKEDsanbOE7d5bdAG4x
DYv5LYlPyZ3PKKHXntBVmXTlFnNvu19kWRYzlnU2V5GJfNVGH7k30FNB5mEZATzz
YU2y+eQ9yeJTjnoB7BIMbU0xbBtOmJ/vi15cC0gqJRkFr/5+DFbTw1tH5f2FDlUx
LBgHwmwYrF2aq3aJH2AhFKVMiCTppVmnFM8dB6dy9oEJ8oRSkAZnguDIx9kWiNg0
Mj9CsekNS6qbF0krLjRO8TuLHJMaYg6T8sOfLZlIQoruVyqyZycJYSRGanBys/7i
1h+5JvPE5VNyWqYvzj6ZetAPFbE/sm1f9OcIMMChI1Jaj0458JGBfqmBuZD8+x5i
Sz/bTBq1M4U1p0lLkyADBpkxo561lJS6pFAvcrxDX2jm9YIGM2WcIgbKBsNn1ykA
gZ8YYahPpv0uU2zrjpFwe97N92Eh9Ymp18a8/UbI23oJO6G0xn7E/8+olb6H0hEq
NDzttoj1vAh4dHunieAc1K7edXMmTkCgF6BDh4SlB0JME4pt8S8TsF9rIlklfpZz
AgwqaoebCerr6cz3ZLy0vPDQtoFeOMzrspUKKWuQ36lFeG5f6zbfIfOtaS/CsjG8
gExWlE1luyZr7OW9kVfK/PiH2NOWdJbvzdUJ4NSCwCcmjR7Mcqe9lEKUxTqCL3LZ
UJO7PUZkypIuCF+wgxQYhKsJI2WUBIjTwQUhBlbJ9YzuRgN2aLcefLMaWd1qDt0B
LIhEgWxU8j5qcKmVQAhinDScVqOQca8FWI6ayvqtFx4xTiV5hTWfvQhX0Gn+bwgf
RmU7IPFBQy0Z4T8sQ3C9n18Gk3kM07tKXn+PEbOsJdCUYcQopEEnQGzAvBQDLVOd
fHHUipl0fyxr3WCZ6LU7CX7HJPQ293E92MCbBKUNR8PTzt7FSWfWAmRX5bXT4xJd
VOTsbDeFIjuPuWfW7X76vWFdSV6Uted+u72V4UGH+UnP+HWWnSlUoJ9aHrOb8z64
I8Ozxe1WD8Is60DsRqPmIMDrSjZJBBwyTk6kDV1ic4nlIF00qcaThB/SclIX6kuW
vdpIGZjkSiyMTiFGP2I3Qwb6XrdcdohdQxY9OvgDwrTWI2Mr7qOjqg7xvhxiiP2F
KDnaNz2VTDWyvNUA89oa2plcboGtCVdTv6DVdJag74ynJh26OvZBPEKTI+fGBEfx
CczEmQ2Vs3Ri/khJW0rONKG5uGkIBhs4qQxFTtLZRvFL6IYgaho0KHaDinyTPjQZ
P+R8V3EjPxaPWhQO1hokBw1Qa6rMSvt6wZvuGWo5fPzkvVa+emZmLP8xvBkS/Yml
RNJ01552nMmZu3izE//tKMIlLBEp3pDYJ7vNeHD0HPkqhnHVY+Cu3E9YElHqzMCM
x74dfZcvaPoLN5+lGbU3d6lKQp/3F3HiASdbpIfkzzGFA9VNU4PlW6rWSwYc/Xch
Kkz5fgpOmqh6HjhIOYNbrAOpMTM6V6sYWyp6Qby085ft3C6O80Z9eBEAD/PuoAMJ
Yr90oW6x+Lzd9O43bY1ikl9jldX9pZWpcym2q7Mw5bFbr0M6UklLE7gzEDlPA9KL
Th6NgmOQEr90BgwPmRTiRuwXRlGVk8Vl/qRyW3aBiXf4rbk5WyZbVVkP9nOwhFRq
Btmo14o33txj0S9n6rbwuZmKg3Apq73xDBRn1ntcA+87zfsD8b7K92dxDdVCjvpP
uiD2J+UaVEirJ/qPub05r3r3rEiSC/jG8wNrslXutirEr7UDx0GUa5eXJdwLWin2
vnfAMYVLc1ghYpJ/0I+Kn8i/0YKBJn27U1+k0HakecriabRaGtt9XBeUjo/2yGJf
3ASTjb3Evd0S06BgYElcj4e8CKo1hCrk70AX/tJC04GETlgC/1SGtOhn/X/nMS+t
5mjwgzPJaJZzbfE1NCorcU58Bh5epuQ4H/SMFJ06vDmUC9yUoCsxhRUUGLMe00xV
Fz12QTNietew45AC9J21cb0QfgtOaHFUEW1leUnwQlG2qHiFZSSb2r3kj4MD1xms
JEunagGrtWR036lryEQkv9Itz8OpPA4LiAnxQvJzpXkNA5ulVFEj5+ixraPSvCiU
6OS71fRtQ1jKmie5G+uDmIImNmNlXTBxVqz0uTisOGsESlLyaiC6bbQMyp+iuoa2
xQ0YP/Z6hHrh3ByKCQ73Vs6DWXb4GFrSaLHrL4eF9TcHG7yRaAsphu/OT67I+qzK
HZOUtCy2zaDK9K+KgjyhEiowt7EsoC6JlDJm6BxzbYq4rSGE/quhBBwx0I/mS8vz
sdfmr7Ps6rwZdInKmzVUZKsR5qIkscDHueAeCTTuN7HtsWKDcEogv2PLes7YCv3f
4vzVfXWioaTqZW7H4r8dR5Ulao3/B1wa+SlJVwSq1ctn7J4UNUAsGDOjbKCChrsI
ofGUN9/pv+P7bJ3aqkbLiRMr7FccbwhaST+CeE4NSdt6pAcGD1twougTJW1urD60
wzgE0+BXE/FTDswnNMdcel2HCMIcBX/fXqqoOFOpY3PbXWqV+xsmijhkLykpE9RY
qCls34MSBdhW708YGvGf0xeHNzq17DRu5FrGgY3alxjgVANCCbr06aOc2d9EvPqb
oJ9Mx02JvGgDpm+spwONzUcue3a2iyBjbYzwrFO8avc0H/hfLlJXGYicup43ceOY
izBkJLT1wDoxqJbOodkJtg6QofgMPU0xfzpiYOXnCubAb3rZURHKmxk+UpAyaS5S
c7fb/vZeNhKDC471Vm4ocCRHWJgRdq57ujqGzZZe89hBe5pOl8hx7UmowTE0r3Hr
NBi9qp4Ea9xO8cT8mK8biSaip+RndyzZ93bdHxDhGiCVdvS4MWhIwvjZsTcpOaz4
gtxOwjIogtzXGyE2eChbdPjLYMSLLUv4ZFk7n/EJQRxGFTOP/dOR+o9kJ2xf849R
nyemlbs12Yf4c1HtpsScMyqlSCF2qDkRLOS6qTZYPEVxmJET8f9H79KZDXBqJs+9
ZyXywRdhOtb9AsjJ0dRynimo/aIPRGf8FdbQyGFE25/mm21oOhrvfB9AmplEk7Oo
v6xnbcgjNaCeIH9paeljMLCZO/vnihtqju4Z1fjcivwMclMZbcCV1BjbufhFic6U
MASBdJfhjGZ4YCN+fqsQnB9A+1pJxVVZiNZvyzdSu0idHfnHq1h77+ZWG5RLXCTc
uwL48s6Vz7j3IN+8RMkmUFtpm71WV1ly0epr7xV/DUJfZfwsuCzttYh1w5TcG1WD
9bBHoYXDYxgR959dTxK0IZO9s4qfeaSY0NBZV5KQy1MxbAHeVtP/DQPu17iOKMkk
vx1MyQG+4BNZZ84Ni23PNQxHBCioQoGBlzPMN6dMiKErH5ElzDbEPeY/eiKQXuC5
7uNuED0bslIG02biqsbllyuGmPcAI9jx/QgRBFDbdOWNFAdyNwMOG+jufMYrQytW
whVgEeUw4N7RC8nskxIt0RNBn1k2b4Os9RX/luyQkmY8PsGAeFVGQLfPLV1OLtnq
OXNdevgtcIhHHU4e0bPNKxD6Qr2weX67Gvlv32Bx8oCAlcn+sTrzpI9DsAF/cqQW
iNh41NboclAqiTup+1htnzgVqfq66PFluufvwJEv8E5dEn+deu8cNJRursh/nytw
78BtOcsMfBlYry2wiPg1sd1/tkQ+SsKMmZTqQzsN0M6/aYgAvuNQTPP5Rh/zB9xb
TNiVZFom9zKsT6Rtyt3hd+GUtqAt6xTBzzxXTUFSJtRg+SfnUky1JiE15GDrEAoP
jchJIuF5zTNYgZmJtpsfoYJdlOmA59o7m3b6xCpfwrOlXH8dMkwY0WAwhCC9rp/u
O9ew7d9a6s7/eTnGOSrgXpj/8Lh8bqC3jpeoOQrn3iyL1NwUw68fZnLC9BlIfTNN
0iIVqHm130e7LVr2L+4JAij/6P0B5xJv3nv4l2GXUhWHUHhIbn0ZWP4jAIXjQUNg
fOciw4NP6rIoVGndxiGQ2usSfyyI7gNRO12xF5llgeGXJc0631mNg7EAa5Vk2ulw
8efUJ5YMAUtMDhgEFBGVwnzeYxZj9pUW7y61m9Vfs2YDvLt1ruY0PIwheicZO0V0
sWfVrUHff7Yw5D5fD+ZiUHTXKaq3LWIH9SMdKaPJt6QZnULwi7rCRKoFP3UZqQk0
qeJHdLoW4UJwEIvIKh9nb5MhWsTpQWH4xsGLAhAhaYGq72nZ0arlR/XDWyUU//ma
KuAUn8J+Ru0G4tzsbJ6PQ0OdG62/qqJ+59MUc0D0kbP/PkKaDy9v34dxmxuGP5AV
VYsEnJvPZy2ULNFGtSJveQpzTxld8JPdZ56POVxQIkR8skxNsgnnUBDFNN+0I+yA
I4KEO3Ndhb6mHh6iz0HQw2d7OWkuBtKri06Mr/lQMaMzMo9Jmhvk1Uc9idVb7Bix
5XCU1WrXopicKqGq8I6i8okFcM0kZXSTrsyCUCUJaVmU/vAuuY9vgDLTrjedUqlO
h75+9Gjjd7yLqc5TpPeu7600GOXChJi8pXr6LAq6tCalJh0YgQUVXgRuOuVIUce4
GFFE0IQM8Va5c5kgFeQxI+3lW6Rad4QD9kEcYvusA/q0QcR85FBli58+7yvpZ3NW
J9oKj+lbQn61h6/chQ7hWNzucc9YCLLi3ohzS47NbmufZv8A3hLuOoy1yGJjrP0g
jBiGB3VEikhXpJRTf8ouZ9M+C3nIfGv9cxHNXI60JhA5f9ReLEWxO2mpcv1m8eaI
RG97bn+g21bIt0vX1GRFI6xE/HMiSCbl5yKgulKYo3Qn8m/geO63/D6ywj86QQIB
hs+Z3lAVnynesPHA5Q3r5mj6pTs3zS4g2RYr5wJaki3h0H+OHJFzwdaXLXCJPv88
imUFtaMbwqdxTKjQOjus5aUXyF4hnOGyh718h7LfOrJnNTEvW2YcFgUSAY/AcWia
uBdn9o7R9CBOrGxm2+MIfcaB148SNgztiCcKfqyxzOp/+IH3av3YWTu584sxfXIB
0QLyslbogAdYn+ld0pcNWbRhEyhKDGOSc7I0B1SiUnurIrYbGL6B6VOj0R5yIBDa
rdTQDGVh5Zz+lVnRi44YBXLGBcx3SGg/HW67CurwtHqUaqE6sseIwZ6cjvhQCZBp
/JdUYDHfnEJhbQ+WRsGH4SCXKqvPescTg6Gvwqb42C+Lpau4WzeOLS0jtO8YETOR
OfY01OoYBXEP5WFlGZJy9a6TtwMsWZnp/kGmAidjHiCK+H1IF+zkY9oOLTxQVqWE
CAdyTLqXvf0prIPTU5TxfCTgOwIQiCbSbbLDflAocJZVEjT9390bINezae2du4wc
KkqOd5x4AAUW2EhYySrp0FSD+ZZxYcIKZ6iJooTLw1Y3xwuKbgIQ+qpdgu4B+e9b
N3fceO2faULuaAoqEEqDed7gmoDitFcdWnpXJtX4hhEkFvieN+EMd7/jW1rqIlT7
cp3XR6kuxnN6MFd5UFagNjKp6AFCCYTAnbCbIMhll9xtd+a7/+ZjO+yoGuYpaKx+
8VWYxME6L1qczim9+2c0g6IefgGBuK8fazoVFC8dSBv66mcsut9n4AiIFkzuSrVL
kgfFHZwJMsk7AFRZ+Cyea8cjAzmk9CoCrVUYUTbsC1USaGOxT67ClIgF52Rm5Oa+
zsevy2Mo9vc/gtzlcBGsPiUnzbafjwSGKBRdcqBgggINao174Etr4SrcPk/fQac0
gmTPpz7qgv69qejm0/C9QMZtwf/s0ymftde5Wr3jKbRqObIEVsR9ThLKT0ETJT7T
RB0J6XqNXznnFaGmEApMGot3k4GJUAO3+Jqo2W57LSlzAaD0MSdYWw7g9H2QK5Nb
VhYc+HnXYtz1tHphXK4eg54htTd/x98ifL2YHBGIy/Hmz3lOVCJCQ64+kwSqHp6t
t/yHD+ibFT6NtIbzlxvWozf0vUsDgN4C7Jw6+cPvO9r8JgcKYHxBLpsp8Bi5v4iD
KgAArNjBZmu/YxqGb/nkuxU/+3wGlDH5tus9/UV74YxPfN/GJJXnaYNJqPQZ25Dl
/IAXx4eFC0yO3sSYevMjzTif+IVfF3AVZI1N2IwPgLF8oaaQpn8tFhvsfxaP25iS
ZB4wcMZvboDjCnL/Ucei0QAX+rk6xd52e4eEcGVKj8hZmtpSEn/fgw2mhN2VZDOY
LNY5T+hH9oEuXa1SHJDxJC7IN4fpSGqiip+f0T61m8InJgXJUaqs2H0lndoDgARd
OvouFMwZ/a8I1G3Baetw6jilF3drMonCquNCx+F/zGmm4xl5FdxE++AmCVYRCY3f
4sBDVDRUZ/tNN80qGw//q7oRWyTMBfhModJRpThF1pkfOVUgjyc5v+mJ6trMrRnB
ngGImZdf8y9901/VsoXMJyshhEracZhqh1OyEHataXz2gRPLtd6MdXNuVsQSaBpp
gJjgsGtsH47oOQE/ZgIKdbaHpnVATlyZYvRzLEuJhE90GSXlmEtEMgRPPcmtSCxh
hqxb0nBP7mnQIUJCg8PNcK5i6/MVrjxtM2q1sGPs1RXcNguAC1J22WWVo+3puzbT
irsalSbJI9wrrj4DQ9Bh7AXy089jXg+mcJVtcW0h2MV6G1OE/nGa9fpDwyMGZElj
jNmnYy524OAPTIWym9iWqFMwSjMbQvjCu4g3BLo+AZ0pHNhaRLLAqWCQ73epG9IX
UMcGqOENwXzDS0MFvX3FrmuV1YYWpyy2HrKV3icaXHJS+RG2HPb0DUhcHOXDOlLa
Y3e6f7yTbCK+oYh3Yi+cdS6hiuJmq6m2u+DT9jyQiz0C6+5UHh+dXq+S3w/YgdSG
Q7mqkbB1WGaxLmSXqNDYpgsgFt8TPuQUZ3MObsdUTC98ISDhwU9tZ/1n8nYE2Klk
P+PUOQKja7XPnR0iATM0U9BQAu6OJVT+u9VtGpzpRCsE6Rakm0o3ZtdZdsvBTjxu
10HOtAVeSxriDoeqaHhFBLfCsN5lOUQeJwHsV4AO3Wjkyn+lxXJXERQ4s2Me4rEB
oqei7WiLUhJX6+NlRUv781fup37SHStOPWeJRVWv0J1hRutFAtJaFtUIFBrTUFO2
jPJmDbST3/uQPvKqthoVnGu3kkXB1Bv54q/httNe9dYNgzT/FaDnvJ9yv1IroI48
bU4/bT/4fzf5qMOpEBd/umDJWmdtmxA5yAEqEQVWELoRjKxw2H55KNxaoMH5CpVY
mzOeOWgMLvT2Apkhi2+z+o7uvJ4TVHGy//fOkms/7oDzPqDE9hlNOi+ov4LVtVT2
5qng8JPj/kleWOopD7ug87GOpMMncMpjF1Sn37eC1tc4WRJlAxjsvP4LxcsyE9Mb
zbbp8LiyINTyMfKHD10SRuF92UVqTKgsX+AfPXZ227AURP9ku86RrSteWdYKDGdh
ssr7rmb410NDmvSIif4/EGp9NBBiID9wCPkDYjN3lcZ1z3fGARQpaU0tta8j4Ng4
BufCIWRdMO+bD7+xijLvirJgivR1KzsK9mPmySK0zwgNdF5+1+9IR8787r/mj2tv
QgUzJUgnAu+2HKhvwXkCcvQpbKyNdIWF8iK+qDKP+aaJHVWMx+odCxRTRlf/FW5H
p7DBDZW1+oYh22Nv9UmV/Be1PPr/4OqX5HhNWPMVCKUa8raNOgpG2hucELiV6UQu
Mz80JQ7dvCQ3gnOHFU8WkVUOtKN/AZ3kn6IRRi8oJvgpWfmT1Fccu9cR+9pFaAUH
S9TqzHPD5Curqm9PqGxsKgPPlGgUzqaKnfFL1u/n3mJ5NRUWJ2BUeDpXwaJnmgn6
8ifqVbNqrTKEAvholRhQKcPJSZHoRFF0MLcT7/hvm/CxXnAJ6pHTxmqSqTLNzAWt
SmXMhK5CYfpoOqfjd+vDUP8wK4Zf9dMKlOBFvieNH4K9HqSqXUm4U5IGH7SMJ8r5
ZqfYpAOAkwOXbFFh97Hqs/UK371LCT5WOdIz1YAygFyGp85OGFRDC474fpwhH0Jy
yj1oOa9D1Uw5+wTkCP87KtEHBWw77BjPgGTfc9lIznAMp3v/jXHfn6YxYjKmIOlQ
rVW8A76kcsYZpbeiZ62PFjuRKWCKE703M3uCDcisa+wj792O3IFP3Dq/b5fM0Aos
wImg81f1nLxrVYVAoF7gubTNi81Xv3hRlC3h1SB7wL+xODzum0yuWIzBtwGiYOFa
x1JTEZ/5F/eXkFm7Z5AM5qMYinF4UfvdHVCek6i9oOri0JAJ8Ts2yKQiZKwuxI0O
Tr74e4mAeC18VNsw/au1sb2c3AGe8Oqq/YgzM1W/FHcT3kIkVbpZ5vCUY1nL1Y5G
FcCM43FeqcZK1ff0nz47CwK9xpE7hB8DXHlxTM/1rZMs5RfHM/rrFAGCgqYQjZ4X
re/RugJohgxsNa3BOeUK9EITRCGfhz/23MLzO1GcjHeOTBVwLYNqW/Ji8ggJsAac
4LrY2ofe0iuY9XUZd2gUQ3WRm4ifFXuhEZf5WDx1mkHYMUlIDrDVLXR93+pEgVSC
v6BhSOzeGEWrn7Jgn70T8vS3TwEwDZbueOUd2VykOlN/Ly8ClNBzFWXwUzGqEMBO
wvzWnoOIV2m7r+q0I9m7IpV+qjvgyxLayoxkt6AqCM/lVjhjrngWXLNE81IiqBmc
+5SIO9sqqA4ZZjgRi1uxtzjOjC34UBUPfiOKPu8Tlk37qXTJq4oO4UCPdHNnJHAf
M71U26Ubz3glJEZ75+ibfZ9CpJ4GVSRqwY4ZfuKVOeXIuyYGcEOF3wyE2kNa9T4V
7/9Qywb12/Um3hq1Cng+0KFlUVVde/F2IuR1Lyg6yLEHAZwSGzAY66JUqD/rhVAW
AUPIYreZ9WvgTZG2x/isIKNSj+lKQsNe37NRRrnNMzLgavJaWXC9AyRqQ1n0yeIl
TMSvew3RkS0wMNsK8DJeKXBR1jMXQ+dqEmKixBggkgd9rrfMqhsGD/lLp//294xa
bFeMrbjiakxHVLvrPRjIAHXARfsjy/QZxmBym8KKgn+KgXOx20T6fStbZYlxIOY6
B9pmkSLXvE2KvSEikD/eZbQO0kt3vHw6TmWSP0DKoVoV2l0yjQloN5WHcEDfUt7v
7/80ov9ZTsuT3WD8koxlKvA3uBmWhB6+DOB89lih/YMPGr9UZB3xkfN7V2F0mUB0
PoSIconyCiTeIpzdGtqQf/lDcB9xBprTn7OTgt3cEqNZYSO036zEKRzIJ1XT7NOI
Mj+fzJAUuQUpWDsh13C4TmimU9nuzItxP8rKZRjZcnxe3i27ZKz+Et2/B1/bkunT
VStzS3NOnE/Y4Ml0J6W2hoXnsEhiU70tPUV9ZHfJa+hCPqIumb7wMUOI81lK5xq3
yyMzqwg5n4YrGHzX/BkR/3VFLQPYq1bEYaVHV1lG6xIDEjqCirwcXDxYgq0XpZPK
1MP7153ILm+dpHRXHU7AJTzkeeTh5OgRO44oo1QvGHuczUz6k/QHDDN6Z5jD7iau
zFuXdcQjHyJPM9yBYbLsAkIfofjK0Z5ZC5S70Lxitpe0uOL8JNiKVueVGEbUX/kv
0FJDCNd4RLYpLG7xhYJqGv5Fy/B7rMSX6ZWwcqHU/Lk17HpG4TO6XEP/lPAYU26G
RUQHBFhRN7YAJrTNUuUQHgrqobf4L4mva2jt+Rp1NOcPwtkfzJLOR+gGvkY9qq21
+x311uJx/hi5gQrVfMzX3nSuT2RtKOHdrRnlukJLcsPb6BwipGShJj/sVyqMFxrG
mgOaCVztgp1KA1OUCZFnw9X2DlFpXi+ul5jEGNfz+ClN6uYq7OTxmL+oyKVX1eqG
ZKoXik2sYyXGEVMYwz5gImA2x9faKS/ZHvINLZV16w45PPF7BpuW7Tt4Q2TETUfT
H7he2nnobeXFpiy1SDn3TqtEYz1m2Tt5k89GRw6J0Ak6vPMmHkDs1m2BB/IHPaWV
vRWBvAgqkGFy4j6TF44urVg9Kc86vnausSM7V8hi/pVXp7pKo442VsRb8etfxoR/
D89Y90aOM/SOXNADgKarWFadzof8Wb7jX0R2jdKcKLQo3FM+h0G6qMNiKvh94e4I
mq07BgJVtW4Ig3m0AUXPmeAOMTwTxcme3fyFH9SyIGwHtfLJl2AI/G9/XnrvOgZK
giY4qNok0GHQhOh0DycV1uD3q4yWYw0bRBVUsLFxzKCIFFOmE0YTRrlnG5lSN96m
MWrRMtK6acbhqTnhVEuZti4oUKOz/SP85qifsG0cKi3fCKNKaOHacvi0gC45zQPm
3NhyDk8c5daMk2O40j9TCWXmBaZzDupH0WDwf+lWt8TzSfuL1wp5WYc4nkigJf6m
dqYPccpYfSk38CMkig5YF8N0N34PtyqEj3l4qQmawWGK4nWja7gtTOWzRydP0V1e
/6X/I3BbRE+SUzPXdoOm1toHjuq52PdWy1CN8VuU5qAovl1M/RIbX3J7eLRg2nOn
GvCc5FjrFqCyUaMKVOavsF7Par6BV2T0ElFoGLXsiHrTuaHd/e5rL8AMrYUTekEj
+keY9pywVDXeghYiQrqH2MTO6uegjLd2YCaed8YvT8g0eD4rFlLA7qB3RWiAweFV
HQgkv20aDiL4x68B7H+4BVDs1JDeJK8EqYRqBKCCv91dgxWNUm2C2LMe2Yp5LMhp
F6bcYsI5T4MOk0hq7CoDE1D07u0sFqx8n0jq1xNoDh29aTRrrxcp3vt6IznCWnyu
cw3jfAFlq4FQxJjE80I+njnoBUcQ1IQB2Fs1E4KQEOSlTFzEGhZJMvaHFu+DRJes
9koAcQftnt6Qpu0TrgTZ8bTjIlkygZcNLZabdjwz8ogoLpzsBGidzUUzCPXL6SyO
mp1xk6j7jZbjYnzXOJUWgtdStXlHw1NQPfpGCNrtRT+lyUTV3G0mJSQaAu4qQgFK
TBXrbMLHkCD0RWveHuwRbAmEccyhIHU2LsyVfbBBmP08VXl3YXv9h8PzsVSxyC4x
KEXal0ltwOG0hx4bycCjMICPIRFidesNwuerVhnWGtrZlpw2aOq61juP9xhydol4
MbHQiOCFzXcVTmpVOcmnBEE6EJ94zxw+qrA+Uuwz9BSqKd7SEW6rcTje9jnqQ6ht
LY8iXAUlDPYrU1UgpLFNGYE023cfjtlYR00GraT7qFP3xHDZjNTPw7Dtc/4bWo55
mVYyNJU1ceq/zVOcTPVroC72MiFCcnTcLT4KvnoZ/Mitj26pzjodjSIO7VpnVpnR
EJHOr28PKvCPWf6SlRxPptQjRe51L2F5RA9XI2r97hPQOVl0I5vFjtYzQPKZdNm/
SENTJCrbVfG2mhxyEH742fXo9obhx1eocaViu+eoLA1fDjzL4VGi8/KlT2E8u9GI
uTvt3ippGR9ESHSheYrXP02dkXnyZHnw33eYhcfONpoOYZ/wTiS3EMAZ/3JvpH51
Km0lkPYmZG+zrihME9TR3FFVsncbIVAS73hYOts1btTMtJdXtMeVfzjPIQfW4x/a
S4wqXnHSlglvmUeEL4KVELIBqiZJkc9BIK2MCFaIY5oqJqvnuAQYcZsIb7DUpaGd
TRoO1kNRuereBwziNMszBv/TloEXivEbKXe16hAZyjkm4HRVY+1QVO4OPgb3ZR4S
Kx1ysmRArDBpN5gPCPEYAucJTo/KoAQQ6j0hxa4MGafsot6nkhM53gtQ8g09TFlf
iVDwnYz2ameiKK7LtixG9Ap7p42jf74hdNYa/mz6YGB2f3JwIiWJHQb3Pb6Gvg+s
hej4myRqF1e2Wc3PzUqgMqGI9PQVj+iDToDMz6zAgHr+j91/ilQ5E1o3H8kJFTrT
n8sYKA+xti0n0alnjk9j9e0K8UzZvIkASP4GABbI/zMg25wKqelzurf2838i27zY
U9Su4vMYTJhBz80wIf594vwRSjgMIKr47591CnVTlq7St09CUs7qE7G0R1e8TFop
aYWUgHS8SOqk8YoibgU03pVREziIdtMT2MvueOr6xovR6LRVfZW+TzbEiDkvKw+s
XWk/jbvu8jnrEcvzqi0jFKTyV3DQPi4Y7j4QP7ZG/8gIYuCrzDC0YN5GwN/acMee
VG/aAePS1eEX36CYexEcBDT34+TBEFxNNBWSrollwIc+/U7wFhaBPrcj1chla704
7REGKY40HSH9vkvxw6X25A+c5W++7146rDUKZxLN6SgVoLwfssb6p5VwmeQNRfev
P5OajWrfsta0CW8y/Ax0EWmZErk61olnXLNpd1OGispK0KbbT4YzLShJHIGH20iL
C1tRpLc1+JgPfmXNUy2ZE2f+95TSEfBPtaLg1Tr2VV6B8iDE70w0heSdww4Jh4b0
f5Uw6rWZn9SE+cbiuBNaiuHKan2RacMLg60QNgmjoNLQoJw45Xwh/TjUurwb/vhu
vNtSVUtsarNgPUxKHtklZrnUYZpMnpQ52KSgzh7o1Wgkxjn5jvwSr+XXyYjui3Zx
VSLbJmCNBY2Khp33o5WwMmUPywKUGPws5Mc6V2fBtT0O/DHTba4N/T57XpSK1c2T
8XXHT68qCvwz8IPHXcXvuk5F15ByIUz9lAxjBUJe46VIHM7TYidpsxr4BJUcE5i/
wDkf9VJbO/FomP31JJlJlwr26u6+qcvuKDf1ZILOs3nni/3CtvV1oFfSAid3Z+VV
ifb4CBAxAQXMUdIArff/BlcH1rpP9SOcjhob6GPVE8WJ8AJBjkptcGroz0C++UXs
52u+f5K1nGiqGabqJFunXScby0Hraau6FbKyMIe8Osm6UmOmh16ugcujs8pseJOn
sDeoy69Nf3gAtC00flGsGGInEiRnOj00qyQq3SUWLfEYvPRhCpnSacY6Qs0oAYLH
WaFwTBpYWt/N/GPTt7OCtwTljX1iH7/FnJ2AbDyEJSKhZjk/pX9hL6CyDf2LBcK7
PebqNFtXgoyID+a0oEFKaHHS+6Dyl8pp9E6OE60zjrCztiRQCbk17gL7KENJz+oF
4cnKg76R832mB81aSRv1f7rFY6ghqW32mK1CXuCXjNiCL5IPfmp/H8IJfRZpt0Rs
rT3NfAatN9GNpMbWiVwEBzDILxTSVGWo9PzaPrXmZW5hOUuA0osBzAQ68GnDvsMX
4iAuEPmxxIxiNTrhCHoNmdMNtxSJdz7Xn5VoxRbszGnR6bkrjOiz7UJdG1HWM+oy
BB4jf+4X71H6pYXp121Nr7tg40EgicM2yFR8hM+Yegdq2LulKlsO0OKKkeL2o3Gb
8kF5eg9NMiWaIIHeWT9n/cFd9pddixTDqQQoYfeaitiN1U/bfunXEyzYLHUl4A+U
5oClrfutas+IFpOeomLDvwCpHqQ8GVVJU1oU9LgKUa2Yl++8vuektK/PbWh2XhCv
zSUF3utNUHs5S0hOYeMgTiG7gk4BpvNyFdCksbd8hDKD2KszZzlfeWDGQF3uPs2k
qfXHb0P+9mU2iP7MsKkUl7fR6xJhSMWBSYi/f6qAMY6M1rz9ZhAfOcBSrMDNtWZu
edoyatwDXlTejlsrstb6w+uduR/J0G5Z7EuINIU/zvzKx4dH0X9/a74NMny1afdW
62kKiHYwDeHB9h9UK2I39yzys7mBVSn/pe0cV/lVmOUCP0mF/QnV3MNon0eJjaj3
nSDFowZMtZZFsytyFVU6BF8l/cfGMd+ZYhs/jHYzlIaMlc/2CKQ9O4WbYrjNU9vf
lGTePVOX9wGYq8e+oBdsdz+Z/XhpyKIkzzp1s2phnRMS8BG5LEiWaSP5EqQzKCpK
I/5/y6VW2PtZCnxMcGdl/sVCtXHuJuayy/rnStFfZ4SOkZOx7pREgdlNmyL7xAxI
X8PZXfg9F0arzhsy2BvxP0c/zvuOYxkl538AZ8+juOLYVcDcTC8MgO/dB6zzAsPM
rM0DPTSe5UhsfWJWyMWH1McQrIUp49ESkA2XKsByHUC1TkhdSrwBVxmmKRymH6jZ
Bd0DpJv7vMnDIIWPH7j72UMf7NNCqdeq9qF6rV9J2MoYGMClyDaSbMqeS52BcZnX
tSNMSO5PdBLycV5bh2pG6LFoF1raP5eyE2+d7Vif+hXqT2cNDMby79nkKSIijrXK
zTM88rHzcUEEbW3ju18QidkXuuli0EH+UMOT+7N/yKuWC1jefrS7sYkjf/NmZ1Zf
giJYJ7xDe264S+YwGr/AsauWeZ6rCiEUR4B2l+PkAvwW0iVGF567mqGuF4sD4wLq
uSr/rplQ/NDWlje0wNbsFy3YV2KNEcDQ/56nIDr0cmLxN0xza36UE5iLbo0sb8vv
w811o7mqnhIEC98FCU0AGagXTEF0ogRmzbEiOh5PaHIVveeWECaji2IenUAHc/gh
/ZIwDH9jINyALbuZGD6JQvn9sRqgHeBDVZk7VABh8i73O1O5Fgp3m9I9bkWRyJ6Q
bQDJMYM4m+atyh1vYTo6l7EaZrJUWu2E7IaPcvKvEuQySYTWhdvN5lc8Xd1a24KY
aaAvTTQipedJxHjWMg58zPqCn/lfj3lKBJqMIOekuCOx1gLbWaFIX6SzYoaY2GnB
8QWkNnTmwvNen6s7JGBxqIdyIb+c99B3MjQXF5W4sgclPkUiuFY7YbeRaiihkobb
eU7DI9S/cTlY9YmZgEXqDtL1Ftr/Yx5F7Rn5mJaoAeJZI9SFGwKq4PBTILpXMzEb
YkpUdC31rSSijxz8ZCVTajhZKiGltLtSH7n6wOuYZsoWP/vk7SAOvfhTv8TriSYG
JHGwj894ogSgvTOWzCDCM71RdzcZjHCEl55O9sn1kOPx6IiiXbSIXIx908pWu688
JqSIp5HMpYgM8x4ebkoxoj0wTvepSxcickgS1PMGfCX7Am381D0rlHBUCEAESEUX
M3SJa87kkMSUIO2GBwkwTT351aUSJGP1Cl722gvcR4TAF2xb7EdTbUnTurcBCJVP
8H2dVn8OYkBnh2PCaXupbTFMQJfTMPxswkY4ws+GauiVr/ZJvrCTxsSkGhvEZ/Vf
jRuRZEGUcpSIV4B0rnSFaXX6bZ52y/2Gbn8jY+7wrzC/YqzpVwv27BFKvRIAlnVe
kDJrM2bjWHdOYeHmVM+CRDJznxerPrUzY01oqDlSssbIe+kuHvODUYk7PIvAnlzs
Q2BGjGYxH19hllkG3i/V7AZTejG1naDyDD8y3/vfdAKXrx4B4pW40EDk+DLIgg9n
K58838Mdo9r9qbYVESBzGZbA0sAREQwuKMvLG0DMixjMVEy4IsKiw0GzMqzQ8wE5
oBqgjzTxyakiac0InCctmTvTaWX9NnZD5Ty0aseQxyS30eDt/nemv81IbIEZQGi1
PwTiawkLdSl7p6o8wBtWHidHyFNFKOhPDvimT4fmeDxg26YpUfgJHU7VBESIGW3C
RzUhnb8NprrJefhh05TvTu1w9HnbKsmlvt3xe1T2TjWWQXMtx3P/G8rU2ZWpp5dT
8+eD8k3CD9lYVq6z9wostG2Uqx2MortXMdJ0PH7PT4k6yI7WEKrujLYUGfbT/WNB
qlBWUcFyw+fP6jm6Cv8CW7iWv82pE4i9NguZd2eV7b03my8d3QdziR23AJC3DjIs
0lg7YxeNdpRyNAento1uqjQbtMOgM93SndCtRq8wPUGHJgUnmEbZhSej7/BZfC1E
etPXIQiQOueEL/lZ+p/fOjMtXUKO/bGwI+bCWkrhfxvIxLnVz8mLPilj7zEcUITH
7xPX/fzSNS24yUgNL1Dn0f8iBsaXieGaBb15l46biARzU3KOV0lWQXvHWurb92Gg
vLI/GVizVoYuVDobgHIjmkN+fcZw8ytDY9nRtAMASleqmR+xmm1PwmpMDUFznjZG
gcgMXyTCKHfD7wY+SRlGPmqQQb134aVN3++qIvTEeXuut142Oe7KI+y5A9bcsFLj
raFDtNeXyQv7DPN1ceWMWwJuvaCtSSqU1A3F+mkHpLZEi9FSUEPcdXuRNELK1rhy
ueYiNvrgM1PVD350EKdipADgwl6i9DwgiyV2MtDgPSpBATM6GlHxKUCW+unllcRn
y9N9u6uni3RwUT+rHLe5U+ytmyON638fIAxT0ZpD8wq7LrdFIZUd60v3ldrwBTgc
q5VSGK+yDeCsZXNHZbmIeCtMcgd0k/7yfm3OfSZA6uKQut37ubvBiwParFbAYUb+
JLs0md5VQoUp3zkp2Q1XJLd9M7an0T2jWw1ArikOa+Chjo2rvveQLbpnR1jXBwdv
VnVuTWoej+7nSwmuWWJH3zg8lQPyehBG0Yp1vjFTyrdfHGEa9LlLjzhGhAZ+tgPj
wOXyAJxi+kejK4S+l4s3Q/kYvaiAJ+YYWdbGDzsK08tl9fhJ2RCdQLYlefNxloS2
kn931qZ+Z9O4V2D54tmnHIpRTy2Y6vXsUKGpk5DdPUycecja7QhHEFZwY05CdOUu
ikF09jhNtW8Yqm9XXsclZqCh8W8XuTv+g6jzAsmwnkEkpYa20fzj6s7wli451mCB
f8xOEg/uXNAJKEwwuMuEpxcLCY7CKYz4kOQde7BfOBYNbz3alFbu7Pbit5v+dZUE
eniIeTuWtDZg0geAPgRly1Mjmpdxivhs9q7uaKI5ENCr1lizhW6F5lfX5R9yV2FG
XUsfZVsLv5Ss1+DJgQet/YgP5nJs02jlDYkAAKPzoqLQA+3jUvRoBI59P0TMrnXS
+C/2uUSvuDVtv7XidfP4jjvUADiNmmOkQYn8fBfgYWcbfQb4oa97kkpR7aaql9Nu
xcHFPe51U0/PC8LqHuYuA0gRuKxPVGWbZ0JN6VU5+m3ggsvTa1y8TrQivjkUv6m2
4ggNADIGyuUvcM3l2ugZXAKXljbpj4ngi9gcHMAcWF/xqQ219IPaJomUhxADHH1l
5aQ8ZQuerE6F2Ruu9O1bhuZGjqz8Y5sxy7/vR+2qBf/oM7Nb/+ih9iZ2+rJPC38e
EIwkVi9MR8EXYSsZay/Z1IjKqx1wekEidr/NzvR63PZ/vT7sjDORzFQXbQxwRjdv
tnCeGtIIX4wSSGxmkC/SRfC6xJeNxb2y9sjTnBTcgymM4Pjafgv2JRL23f6uoMU6
5mJImm5MMsePBvDAnIJWuChH64xG5rmn2MSFzG1Oobvi4PcHp3ZgrABKlNZrabDU
u6952oLY8DgFWWTwXh7EEvQ2ssAGjKY4u3/0A/KYzyfju5KYmg7fwVctQVjeyR8m
yJ1jmRPM6jVs8AIi01KfP3dapCK6Fzj1McwgzxTiS72OUiUs28N6fuBhXMRe3/08
qu2GSiLhLv49XZMI51EptecAcuiqcAZVHhhe+nTjUAFdBIBGUpVHuREnmILxseGT
c9xZLhgdkjXtGjWeYBsoU5cKZ95K9j5kIK9CLorXgENuE0UxysiiNocPQvw/6KTq
Ip1BKdYA3VnNyHG8ZXbz+hI8caonqDocbLFGjHNwxbFbESMpcjh1ESPAb6c8oPYY
qLSud9jnNKP9yx7wHgQeNoKRh+mJ02YUvRjYIcwpqs6xKkPRt82cevPIYMOlmiuv
BQrRjQP3dUXMwuaibOnTpjW6mrVChDea7SgcHTdZzdzjNBhi38ksibzmsznvZO7r
Rj5tamzvHti1GszYx887LrUa/gGzJ7XpL4a5qkm1oA0czBA1s4zb4lw8QMhTsNKE
03WhFx1mfTWmwV3NunSnnAhbs/Dllm04VrZIndRnbmRPwMCG5P5wxhr334UCpzRI
CRa7vQGD9/Cpm117RVgQY5/DJfblCel709BzNC+y1G4sSmA3yvzDm7JDlYh4t+hG
8V4WZU4jfKGOAh189cxrIl86T1/w5k6r/e+K4Rzp6px1W+2VCo/NIz6vy2LsN0Rg
2FPJk8+5O0FNVIXZ1wLjgARBA2g9HrWNpF67bIn9PmYdmMpUcpJTJ6CZI2NJgKbH
I1bnkpK/xppfzvua5pGF50CgaE+O0J1OLal32xJlWXrs3FlJhVpG8ilTy1lXzDwm
q4ebWO/Bi5YtPJ8dOGhtO1iule+NYs92OiUMB8+RlqKsx1UMOR8MERxkYbzA8ZwL
Sy6VmjiTdh1OgCnxIm5yoptZ8xTHUV5fOS8MLRYGwxC/zCCyE/ZOHMNjD6KAzRrE
c1rx2ciBECaWFUtdao0XNmVpFdmihXz7TKCk0FpzSuOV5lSBMvH0RxqS+hrgzKcN
0DcIelf1luUe78NDxC2qmrBChELfcfPnJX5ESQeEaOqZNHBqFJMrqxyQcQ3MnNXF
zDmRMuTqOyX/YwCapJ3VIhXYceNxLXdwAFxdLKZy50w+F8PU6waR/eMPb7Lmomt4
tI7gug/f8ZLI1rTk7RmVJA0zAlPpHIw9nf3HTUSbvUdjbGWRzxRAb+6p/1zYTGa5
wXRmIBGqVnJy/T2TKrt/jCizag8IwgtceAEYNNOtqdyI82MAt10KqrPfHARv1GRv
1zLfedxkbvC1Y1L9BZPwslKkTP/N1xuKdXmcEuJsraq9MfsTArLrzqz9WNDZ2KYC
8d9nnTuWVOBR1MZPOoTJg6vqGGJ3jxBLaBrJufAr3SHLebMD6/8SJEXcxfDDXFFH
tj+l/WGvCWh8kOfhTXvezE2DEmJ9Rrl6RukbuESPiMvUaKDwb/wnhPvGqHNYjFg1
ZnzQYjmZKaMmpmpiAbcF3eTrxsYL229qQyBM8vJY1Dp0GTFsqiATH11pJIOO5WoW
EFPxbTBj6CKC+nW/Ut6SWWDAAysjXuCmw4/1W2E/LakYwNf85DnLYRsAOtrXIPTm
Zl7QBHieiKiXqY/6SN+GxrwthNhLcl5+U2RuwCaA8s0YlV7jWgO5p2cJchUojTqp
h1mPsvZ+c4B50aKhu9RCNLQIBxx+d8eafDHVnTlXCF5WDm4RFYcJMkueFZ1cPkuh
M5oVJ8IEOvYWWZNATWTyZdQI4SfQQuQEB0JAlyAm5DXG+hzc8ahw4tLPrP8bDS6x
oPJ+OzamiOqgVPF3SrkgYIYeFZaEqySSVe4gIF80Te4iaLxpCh0Bim6GovRjZ8Co
tgJ2W0LGmi2gRQnFVq2GLk/3dvo3HmTjXQ78qRe/kzS5ZN6SrbcrLC8oPrntXqHc
/pAyUJzNoADPK4MrsyC1w7mm5Im093IhvoXAPi7qTnepdgWf2EYeLK7jNcuzjl9i
YSF4f/U8pZZIFRLiCwn/hKBzCrf4xz/NPz6GqJSo9SSOdpdMyFHg5oQX65mvAImS
8mK+lfiKTXJCTD2ojesd1fR3CaTLSGgCeHMzis0AF/p2o0SRzeKog7WbJBv/kod5
6usBINgzkO0uSKHj/zPRpNSIQo5IZf7hdUqDpkRkEphNvBai7kCIwqR+xTD7xeak
Hb6hCPfJaO0vYBGWlFdCu2hBtlZ+ozJFANYZxwW3RYkosO/zoLMfbuDXuJJ+euMP
t8yFlwejgm4I7EKC9JAflEf4VyI5Q5NWKZc9vV+YUlNtX84eI7rh7YaWv4fA8cwm
rpvMAQ2keaLXkpP2BHdMCdtodw5flyKsC6SRo0mJQqYPJ95NUHNTtXFL01s78Xby
XyJtew5XaWFE4a0TXvXT1Br79Su5ojb+Efz9/hX7xemXbC9OcgU4qIHaUpwESqyg
+fM3o8uVboN6Azj1VVN6e4Bya5R9vTo5E1z48VnsZ9XGFI1RY7S9t/mvQYI9C+YB
JHg52hmoXI9DduXs6r8Pv2socPal6QEQwUbh/FvCmPtSpsDEEPW/hkUgUcQoT6Xa
nxDqqoSsWoTwbVcNpgy7+uW33apli+M2z5rVdg42FLxstIsbzv/PhwsqtEVsXdnh
G9FoKBAeRdZwxlch19VYDHDAxZaLTXqsicriS4Haes4nO67A7PDS5pEZQZuWbElX
eQhVj8DUneX2xovQjY6Mg4uyoWyFgIhrJtlt+hBNthUAqNni1kcN3kr1teCTP89f
s/trf8c1gzciMdndFO+/Eays9vnINHMiR8DKEKUG/UwHMRGPQrrJqjxGjYEgXamp
hTesPv/nRONv9OnjCCUp+MrgIGG1PZZVP+6SiLSCQMxaDytOVD7u/KzvaqPeTs+X
hbbCm4Zy30ueNPO4bp/HToMywvJJ+qSevKhUnVzBXRhoSziHZnZYWv+SNjqY6ugB
yKMGIWys0Ixm4w64oDcTx93n7MqiGxGfRQrDIzdcbmvTW9SD4eeqed6sTxD+ErBA
222LUDSem+xemtrdh4EME3Et3CW1BwXB8ZtNXaUsUDBFzln8ICa1DK9VRKX75Ebt
MEi97jVi+3WQb6gRDUOlZzt/xpswUEJCey0p8K1YHWUhS4bdY2SkaAHnpLwouUdD
EiPcUoHciv+DhqP65nxV8MOad7ET+/TFZVuDFQJmRU8BTQXYaUq400jvReghsyun
Gpl0oq6c+PG1KZQPjbTLvXJrVq82dgTVBVIQLHYSWQwIWnMTvwDrY6jwz/cblqsY
oAU2AoNOgXiU0R+SakrY7JRic17NRqlp2EQet2p3gdioffMOaRdWY0K0xNqhbHuZ
/GsYpSipx4Eyxyz1P88meUFYn8RWmjeRN+f9DdPzui+J+OM0Yr36BnXkQgl8S1zO
3819dhD11wis2FkaoLn2k9ME+pvqaY5LawIRQ9s9jlzfdWrUw84E7iatgC9UAHUH
A1ewXqnV2W+OFlGXQtFmySEkLN8T2d3JVdP+Inx2Gud72jkc0YLpgqduvJnWFOvV
gZDJUTcvNAWa2bEANWHdmVaWyWjrLYPEMmZydRvRP60vdXWmzOgZyF0b+t33xP5T
/0W51LW2W8yDiGZS3MTiIz/MVKg6Gk8PNKV4+4baNHLcv7W3iR5DWdZl5LVF58qH
KoUnpHOEIWfhmfeaOxO5h9CowIAC2KZLHcFk9KArVazYKQwAvAW6tUh3I1EdxRDH
Eoiylo4dP0vKfObJx5gCl24N4Of+cWWkwSy9UhbwVSCgcXbeKbaEzK0KZPjQM22F
YaqRnVbM4YvHmnw0MX27uAb1MWd+QZqdvQIcNxukRQEz5FfTfBuy1U6xCvutqO+6
jbbmC7cN+cR6CpQau9aIKOLwXkRJYl9KkATXTkgi7fIBL/iAtsmpX1J/Dcy7J8CA
HgUEUKMshMic2gE0AO3iQcAJL7gH+UfP61olDt/6RI3deORG+lFX0YK2P+WPCquh
PLmYFn9p0i82Lu1jw667lJ08Z5cZ8nd66uRfyhkiy//SJsDBYs5ps2zPWDug4C8/
8bSzWQpsuNUL6sL8/3mAPST1nmGtQbsHrWw/F8eXoXlr4VDNs+pKrxTrufdgdLUU
0d+MXr8uA+jeubi7wHIjMIvvMqLx50Hwz9SWxO+YG1dH7xsFNNSJ/pEpMd2v7Chp
4uSltkzhZL63jBOMJToRKKgalZ4bVZPFLrwn2tIdHph+f4m5QnmJtMpY7ig/JCj5
lQwMxlFyDdqBASf6UVZu/PtqS6Pp1Yu/R4jRDrUvLEg4+ekCJRgi46Eus0L7YjLo
V7zt+qcH6fDEhb63lNBCIQmDQjZCNX9CVK7XKLLTUwUJFAGqFG3Eq6Py8GX5s2sN
no2Vng1h7l+UaOtZ3JVNK2Yb4vsEFP/xihRnetlkbcauCi6h2DB3nDGk5zEzBdim
6HDghZndMXB2TaNMiIIO44hw2rcm0n2CruqoNvFf+409Mwdr2PRN3myqnPJpqlPe
I728vtsgpNu97MjZUmDn7u9Mt33vizqe/KIKXTwpqBPl7x0UPY49Nmy9aOS6bULQ
VETM7Vyf7g6/sj8Zn5cBus4caV5TTDffnRFNC5H83r5uQwadwIkRwn+2sSJjCXJ9
LB75ugBSsLaD503STK54JNiLPo2a1nJEP1RyrmX2Otl6HKnKYjfAMCcq6gmx83M+
A+Z4nK+Tjc28yOsi0XtxV7zCaJGTFr/zixO2smyTuoskwcljmo9SYmW+X1FsFzTe
raeqlWIRHRaMU2EJWD4QIprS8Lhxf2kUFrKgWuA1I62yQMn6sWtbk8oGUEzTFI0I
2hvigyBnm3ls/nYsO4yWuqkHyjImWK9X+WV0/XOg64IehU0lLi4vTpaSeT3jQuLu
QycElCtH77pW970LrlRXpnQZXI4gIKUizKRhQQ1bKfs+Oqd91YDZcJZrE8KndWA2
BPxOMSQn/V6B5H2PVCDm6I0BLPycNT+4/mB8Cr9td0RKmXmdGm64Mg9nswZ1Vb8B
FbFbcSK5/fDqj8uim5sExT1inPT6GNkKnsYpVwXL/TK3jtLiW5aaYz4Jks+qEOj3
YqQAJjRji6/0CYHLDTwYxvB4690DOLobu+qg26qM/pxIRHS0aa1Tr+iTuTHrQTNp
RvhjCcUqLkl2eT/9M4CSkhyxdcot/a6rZvN9mIwxCWn/tYXqQpwVtVW9YPK/c6D4
1bEzThYeZXZb0/sx8fzUpTv75AgKgAhB/+H2TlHaqbQtttlCOkt1DVjk4pV7t79Y
63drXyl5EXHNiMdV5RaiZgOi4lMQlU820O1UMboV7xma7JUmxex1zfWqTjffy5NB
zwHMJr0DakBIYcn9tf+8Jg+X+ygnYCN0oDWN0a7MrIt2F4k/XwGE8rIRlS6taP5x
5yenb0K1qTLx84gHSWV1U3I5hYnO0KhwMx1jRR5RM8heRVhZMqHePQPDTIcjYztW
5wuzdUjcx0V7YeZau8FRarYjPSxdsEZHTUkkwAHVSXjujSrPQaKTENPWJ8jwFAzT
IGxrzElXAHWAy08ig9pkSf+5NwQzHYtrDF+NImEoE23rnR3mbIuBKFvkoxKVCDjT
Xbs0k9FDxoD9A3zX9cLaZGExyvy6povLOZdv5XELYWwBsAvHRSidc8bcZKgitNaP
a6T4P+f0bQ5syuxJoT4dkduS/E785+74c9PzphM+O/CPAHWErJTttSmvLuUnlx2c
yV5O4wHpySNYo9QbHW/+O+xkxriJXdd4BAT+zaaB/9wm56aEgFnCC/YCEKiE4ANO
KfhevalNmXRr7weJEoijhoyTbWuT/0Cx0KRA2rwLz4DByi2JCuKBTaf8NE7vpfBM
Lwv7o0NBHUPCEKHdWRIEMSyiV5o7ZIVcWB7HXGmExyNitk34VwZZYHaqxN2h4AGU
VbIZ+h+hFikQD1OW800G0rC6s3haxs+n0Txrc+m1BW94l8unLDUpBBqeyAQbptu0
BUYWnonWffZpJGBzc0BSUm+tNeKc9ZgqZAKUNA/+HUguj8zHQyBKWCvp14J4KTf1
ekHrqJph++F1rlW7svKIy9c9h5XbrevQce6UZ0DhxVV3dEWciE/ACkisBsVyFY16
/Or/eh8RYcRNdHmZvzQsh+QhfAMLcB0JVpn20iO8BjlVQpWk1oYVFclPXKVAq+i3
miTgGloHYb+ogn3XIpySQ4jXq2w/HRR7GE2EyHubWHS17mI1+0Lp9W4kHsHU/nox
SaZXTgmq14mmjMyHk7veux/ikXRoaMXdZCpF4K4wVq5C2LNlFIpbTsweGeGHbrcz
q9/kxddeMWh/dLOOINPqR7fSmPzKROFzwsDEXCUOOQTJmjlNYZrOIoM/k1nptlTq
DSajeyXQ31FBTlHEkIRhl6qq4kLYTp+LXGRJcwxRXbe8sZfNsTe6mUCzJ5fI9Uoa
MKUegYQ+JWt4o9+PJWUiIlI9BY67eGJtlr1KK7qvXOeBJDstHDP2LNBQ5HL8ykkz
ddg/MVQdlfQ9HTwqocPi3idusLEDPDKyclt6yjnbyROPPycJ7I9HELsRq0ofcA4F
4HbCxV6deZUwxHHV6iAaQKkHY9HAb90/JZqy8tNjg2G6P/sJM4ZYxVuj+JHTsau9
cu71T0SEGXdib3cwcMwswit6q9rvB5oS+Hf+r461JZeRZZr2DuZH7XMqBmcqLpFj
cCe1ZZ04BZLO6iXGYLd/zyfmA05Cc5iTiLoidvRhftQNZSNrDZK8ewHwtIpaRWTn
wBIK6J5oyMU43pifCIbTZBEd/UcWulIvsviWDoaw6jURCQf93cS+ZcFWhpYZ47fA
P1BXWaCwtGl+sN6eL9X+FfXjoKq6HpnNkCviso2HHy5ILRXCY37ILIOdUeTaxOqG
EyoAasUV5zEqCFttXRo7BuFLsbAI0bCXXQRg6FLXGxSMFlJyl8MXybTT72eUCSll
DPE/JHpz2iWxtrk0pARzmFuKZv7WtjF6wSkORJOQ77oYXTE36x81sALSADC9+uRN
AYsiiXAG7gHfnv++LxmAhz3eZQajZWY7Qjso8FyIesFnd/XtE6l09nZF/fr8To+R
pm5VCGcWhceKGdwbOAD4/5bPshZ3I7y1x1MhANuGWWibhf5PGVltEE+O/kvDjmxP
kfl1TpEI/fKxQLKghG60vbTqIqsDS21BFRyZXXPq3I5I81fDl2eqDgigxXnmNYDw
w2gXp0u2odRrlidM2xVzkOt3tTTdXqrq7e+RRFufk2ZmaCQ48gSjWf0dZ7OSJCz3
Z27iwjwTwpQmdAgTGTODnvABY9rc90TA94NjRYA6IRMeDxQuR2YnO2GwBaqZMcnt
h+kjbfEum3BM2egauAYWq4fayUpwjhLK0FDdr1NfomGbgacCMy5TpYe1tYHa0yHJ
Fk4msOoQ4jQmcLe8MMoMEtBlJu1tYdrESvfzUvpGWG7mmK3yvr7sGHK/K+6KuxwN
TmN7BVsZzwOx32j9GGmB782riyrQZ3uY54CkDs/faw4gViQU4uEyu35A2ghcob93
MWHr+dJblFL/CVR7FGGknm6CKf/EXtliIZ1UN46w+IUJ2Dj2J1rRSwUOBb842IAI
xNuTF0c3sd44W7xeKMgLlH4T/PglSiStmxUBDbKviMe0z32FezqrYBJUEr6zhG2U
YcPL/NUXAd676rGsXR8bcQ5WQDwqqU3pOPbye2bX4QCtnFEroTW9lph8rtvM2G+r
YC+1q+guwY4DBR/QLGq2vGg5SgEDIbWAq/VDHmlHz5ytbYbPDpjR6AtmaMQeaJ/2
7fKHf5YMcgEM3HfjGOfRFqlTLfCDm4F3zPFNlIvzNHIXgOGNT09ApvzpbMRnk74g
nglhNaliqi5g/3EZPNZC/Dk/3xj920q9vcRLgqHmltl3SuJhIO9rc9a8bKak5auO
HnBtpPno4/tUYwush7UDGNi3Xn1m7nN1o1DnmNOAF1wrEs19HDTx6JJZjrIpVeql
BLKqAPclDzn505fQqjKdczjX+7e2XL2++UkR5p9soMrhnQUt1hsrAJK5AqUUOSwl
sadmeQ7dC1NkPSCzXyqkPuSygQuYV+s6JTkwVI/BeCJPQsxx84Clw19VGefW9phD
gkW6IC4Nz0yNHDqQMxua8nsrqp4xEZOZU8mZkx5TIET219GTWha2DBRvTFnoieDL
X0CCr7EG8iULSGm4wHEBK27PXzuIHs/w+WcONQMTDz2rGPIHIUpat2cMUMNO9kUc
kSTMKe9zHj10IcLpdsx4xXzWpflA+MAPKQ/zLp9uvgrGOjyk3PYnYuS6CD/+sxbt
3LpFJpnGF2Ndn2JwkrYXDGCZOQtYx7OAjjognrnuGNy+Ri9McPCXD5A84/kTEw7g
tCaIg9MgledYFutEJv9fE7+pH45YqBAlgaFZXw5Khdei1FCZXiUEBxOKUBYzPtmB
hsQ8vcQ8kyISwDmQhidE1HuHBWqpn3gtwyUcmEsf1Ww4hn0Rx6PSsG+D7+u4hLRB
SCWqqEm4xyVPndE1UBEnchSeB6CY29Wzb28UGVPCNOW0wmBubsCqYYWwqB89RI9q
bTdRZxaswlSa1DyA6yWavQugx3jBBcKc9ohqTamnLW8eosa5aYwnUk0MtPdURrNo
+tHPpkRcwWnEsqyCpUZ7UsKIFdvgj3Mw7EYS0lDHDGiHrOD2+1Lw+TtgNj3pRsXA
oAI2pxpQ4TMea2L9K24ond4ojWKl4lQwTmYsPooUQL744RnwC6A2jNb7QAtRzkmV
qpbTb9BkvOCytYwmWwiUqVl3I15liHXTpVIZi1hlwYyjPc1DB4sJ0gudfGtDYQkP
qXlYoyYaoSpXa1o/ZP0gTzBxWCsV6v/QdmHDwhyPMRXSNPv2GAzl4ykAX/L52SSZ
s6FDqEuQrInkuYI26qmgeKwh3kDNDrWm1xnMVrJ6VztVx4kUCiXLjNznwOjvMEnV
9USw5iuaG2BK/RxI7BmRdhKUaVg/bnwcaqwXWe4fzjAvkS25PnqvJqTqITak4/os
dvdPCyD20djlPDPGDaKwH0PmfCirIDNTv2BrZdcJm1Bfzk8Az4m7oyiK1QbhUXQe
iymRuU1zyacwXDN8ilpeYbs8YB1O+EA5kyXGV9ZwL81sVVFPFnhaQz1gckwRlF4I
07Ruj4E7F16tmbo0io8NoNEh9HDF6wauaovFTzpsOQgvgcMSK6F48AV9wppdheCa
ToK0v4nVcBddeavzNcS0em9jVg5qMfS8LyAWm+8Cu6mHRSmIfJSSp9BJ4jj/7xjS
EjzsswDi10L0OLHy9i7/BsKbiz8bXcrS30zrGpiZVu67v428NSKeBCu3f4xy4Yp/
3CNuk6dhn1PkJ/R3xRuuFYQ1xlhTFKb83u01ywEq8gUGPoNeDYCBUQ8q2FZJ3gi1
HtFF45vcyikCptt/nuM6jb55qxJ4rF6Ogeu/87CviOw76KPpWtqet1DWJWppSIHa
tb8TEdUYZA67RF8O7voXclEowqNS4D5imhpXMAwwuqYKaiVOzslaFq4O1L2gxStq
V0nzcHNtod5FzR+YwLxqFQ8uiRUoBxAjbkXkgbgjiD8P+yBEHg4a/CQT1TRQMWg/
Op7KeEVufGzIM0ac3MQqt0ZV3KRafh9wHXq4tH2Ys+LctY1g8JZi0WdJ/Q9ckmNe
Ia9U5mGxEl4/yyQHdao31wvXVn5U1QnZkPWPlbNsR2sPamJh0DwUuhFiAdQNKziT
CMOCuLIwBmv1ynG3SyNuzPNdBLX5TFzwrcCSSptAqidnpFWB1hsWD5SvX8D/xNSc
HzjGkEhVsAX9ki6FmD2TnjTwIzA0xUgDe2eVcafgF6CBEBMnLpVP7B5Jdw0tNkKL
o1bOpEUaQbjAD9b+eDU7UDunkUilo1N5TLNU6IlucWh1RkRG2RcvL/aOmXxe8Oe1
WcK9/bDspJlVFWR0H5/e5OhoE9gSOoMTi86KuwV5H/KestRjuf5MF5EBZ2GAdsBy
xFczBsctfVTA1z0P34grqQpkrpTW5UrGTWMGgGGC8gLJUWFhAd4IUkHx/8FO6/iq
nUQBh5cSApFnxVx5cPUIWuIj+NPKA5dRmNbShTkRZYelebEkoNAd1yE0gjxmkYDt
LVc8PSTczaVbAQCpuBaf7Z2DauF1sv+dk4RMDo8wCoqNvpfuv0J6ZX5Ntsrj9ru1
iPkoVALnwu4PIqfPFCSf8e4UOEk5ahmFVhr5HU//qkyEmlWzrSrQ68NiBwmE3695
mHuntJeKsRPC+d00D8RKQL/okt2hir4rLOuE6cIdYkes4cIyHEoCjSVhbnLa3yak
BhDdLDR0HErb+SHlHBGWyk5IiRimrNrSlxh6Pt7TE8DEeRtA+p8TPxBwQQ5B0PVB
jtiUAzfuxM/mRuW/8UuwMecuAX9cnKeOTFR3rDnCZHp37VX3jzrmXeyM/5upl3w9
D4PBMydOO/dwx+t4TmWkbPQznTdKpI+BWjib6/o6+zaDyR6JYzPJvdrNrwpXe0iP
0S0G6NQ2c4uRBKJTdh79q8WQ8Gv1CPM3HQk8/PM2q4xuNp6deSRDPh1oCh0zGHMV
sTmAIMR2mrbKMQwT0RyM7jFK+1dXlKavh3qx8cH6PA4L46EeUIGagSZXI0Lpj5TR
vRpeQDP+fKnUDH0fT0OfJzDx2wMANitePFnw5iK0bTrz5qrLjv3SYiIAI6kffCcH
dfww1kKUt/tUbyPXNiXilxwzl1y1NyTXI/XxBTcBS6y5ZMlT3ML+EIs/hLihwzQc
xUCFtol8hhdi6m9ahfhJMQBhbFhUZFXUkxL5KDtKLFfZMfAQSpvAU7NJQFSma/PY
9n0iQuOJWDw/rpwshxqvsJvuE+KPdSsXCBb8tWhhjHGAobWRNLs7TiKSckXxFBLR
IY4DKMvHEF72aQuid4oBD2U48Nywj746/DKZFDSd8zdH5WXOesvfjCDuWRbXBx0Q
Tgt8FUEtUvcQUqxIdUt+Jc1ORJeROKKFEwucth8abcbr9JzGkdfTI71iUVPGwMY+
MNEoK7kH6bz7yJXvNhHOQTMcs18hEHd+nRjOXYipyGOjDK3J4uBbAVKDRJ9YrOnz
ouYoV8ULqHd3B2twDPRyGvuytyqS3nF4HavTEtgFQpo0kPMikHRZcz0Xs+0Hb+c8
OIEOiA7pSp1dKcFfLdbSOG0EEyCCzIJtAGqux+MUxOAxlsvZKj5XCndd7O5P7vHu
T8IMiLipkduYK6bNgbyNWczwnc/pB2a0odKk4dRHTmjOlVoZQMeJJVO2zQffmabg
s7D2HpIQeG4m3iyqNH102PEHzv9EfHCJ0DU8bv7oXEkoOeTvhKFNlbu6SHKVc+qk
LQZVsFD+MniyeU/ABWGpdJIGGHBuSuUnTgqgzBPHKBViIrl1a+QCCiMFrn3R+4be
fHTID8xYDN2Ma70/XA4iSHABicAZSY5Jaqw+XgN8DO415uvymAIZVOBu4o2o1ryR
hejHrFajNs36wvZ+2LzY+Z17iR4pc8MdtEtJ8zGwjVa/x9Q8HCa1slXmCf3Fa9J0
umbTh+QDVeZ8fLWLuEBTB/IfJGQG8DbdkLS/4cG2Kc8VcrqGu12f/OhGs5AtPhKy
kn+VK2cHOUoVvgDz75iH7MWervhd4gsEF/6mXxOzt11bulXZ8aAFNPt8tGNnd77a
jqPUs4muiq/XVccSrJu5q3cAtMM2alf92pQigqxSn8jShXpJu1gIk+0jQqHtVWti
umDLoky0aWAOouUwwAjvnfxq4vF6YiqcM1qMKHjiU+cJdWQWPGkVUn312X5XEVkF
mc45BA6u39Ga54Yc1gQJWmBJHaKlsn+vnu74eFuBXVOw0uLbLo/f4QvaH5cHbX5y
6i8USQOSA0bUNVBmdclUoQ2FDnTFSfgIaxELaCDmKPRTlgqVoTKoH5NYd/6K00dJ
lX/CpKWKFPW5xLZPbYoPZUiw6fbRCei0ZL3tNeLCjEKXH2tOn+gHeDRC3poBJmAY
O3sE8vP1K1ReRG+NJFdaa/tAw+1C/MeJKjluUxASIYMbmnZtIhdJs99tnegrFywa
QlJhzVLBzhCIu7KUoqpuYo9s817hwINn8FU9R/4c28tBAocf7J/dFg1GyDPtbvcO
Wob3jMnRFwsIBUJJRXNsX9TY8WJQuzPR+kqt8lqd5fLODNkdPuO74Xl9tNqxopka
PDRSPUcmM7eur8dhQwFtDj7JOt2YRRfleGYZau9NqaXNtUDzWOazNC99MWMKLMTt
jwwv0B8J/zkVyNWyL/k9duUKLgL/PbSbJB1DOvHsBsmGx1Az5+P2gfBV4c4gGzlz
QF0eF+dC5ijD2lDubc8kylMANdz3EuioJxiGjldWgMjHI3RHBCyOnFbpCwfpWVRK
v4g+cPyIdbMOHEl0qnU5maen9HdxLxHmEp0bABYEsWcnXAYOXngY7wg0VPm4/MSg
BdS4rk2zC0MCIKS3JlLX+IikeIBqBEilidPNqTdt1wM8wGOqVymz6CsUX/AsDpy0
sPKMYSuPe+TTy0bAgNeu8Ww4ndoBuhECy2AZUby7BfqoZrj7K7V43kFgiPogTv+F
ibn0luxt3oqzlmmMIM0rjdTL/H1P0daD1KJYt2zl7y0NI2eslRAe5HwTMlmiuwjs
K0zwMgYJAc/HhFy6IW61Ym/Yw7+lmwNZvDyeULCNTVlG8+ssxlE3JqyyCfD4xxJV
NJl03AWd0+qFmGgzhYwPpPuOxJW2Kz3A6UBRNj3HivvmxVDkpu4UArb8gXEwTtvQ
Ienk/afk162wGePsIfVptAEbtqntBubfsgc8nZsDJXQFEPhFgOPPGKnCP8JlaITC
YEZQHnCzub/8hAFeWeqtBq6JvUVV6ZVahum832+xZIJMkcqjZKy0Vdme0m8qeUgl
cNgbHBLL8yDb27yBKvHQbpXpx2+/luc87wn4kedmJTWfx/LEGYIkwBWPOTIcbF/e
2lIpJIS0MIpORy4wbMqCILfDeO66XoeBX/G11DyAl7iYNrlyqUJSSBW7rlTuHF+j
BN/H8oQSt1QnWTHWtv/WxvL9Jjg4QnVYMEkFHB3o6Ap6focEFqR9oLFiOFYEr5o5
Frzzsg+OWaCKd5DuwEsb2HGYFS26VpLQa2TSd03UeYu22GC7lGShMK5euSuMeUiw
d2vehekcKHNXjN1LDK+mEKnF4Nc00SWEy2ZcayUdQd2L/Gf9MXzzLDgHD7zjwROB
kvgOSy4rMinFtehcQtQWbpbSNbMaY0igur9mxFROv1ZV6mgcVNbHMc6//Bqjw5+K
lgUe/ytzJc+FjxVd/7cQ2+gQ6+ltrMVJza/EiMmKWTmKoWdqFiOs/4NAu+0qW6DW
H1WSlALK911INyLh//V5L+oWqtrfPxhiuC/IzF68X9MLdDdrv9oADJ7yeQQHXfNg
D0vUtrCeByxd8RnHXgQIS0jReeKCCQYu7pQwFP9636lCuj89t/qKOhntabXwYqra
N5sAVAtsr8j57rS5usNtE9ct+FvnSxcSQgBpAX1M1lpAKqDSxHMTcrDUHXpS2brB
VkWRxCFIw9AshZFzkLjY6dqNt0gPIsXUidNwEzWzjDqv1448ssA+aus9JWO9uvCP
m4bkHY5njDiAKBZD9JrQf4z2KB3gs8Ie0dX+7fiHjYS1eX53GDMfHksT4AI6lIw5
ZvkIraJ7avZeK4bakTSr8McT7K2MkmVPuSZAyErGy2XaCjISmxyJaAJaz0aoNXJr
yLFGiqKeEqqqBAtN7bj/v7jjgsluIRkSko7qeD3CIbXtP5zrFSb82GmZQB2MJd39
AhvcEIhVPgdLPQ7+34+MN2sHdzsSLFmKSj+RIUVRn7N2ih37qS3Cup1L3fO76a2U
ZHRUIvEJUFsD/+v7orPTjKt8EdLp/ctwmcYRecoAhRd3WfFelClF1WcNvuTZl8Mz
kvRZc3z0CsBM6LSO7XACwpE9yzmBUN7NJipG4beNkrlxXOFiWFJawqhfOcFe41R1
xLl1Clg6V2kOtHPjFkwonekPyRMP/hZAPPKgjrvZC4Aee6sTzG4kqIgfmOUzJNtE
4e6G5pdpP6Yx4cJjjpxUFptAh7G0UxO9PSIPVzJ+/sR9Z0axPId6XE5CLzR4UG2K
pTW8Bc3FcCQzsuaQsjlm1o3O6ZyKBfA649FmCqzWemfCv7E6fUlcB2qM6mePpyvS
ffW/DDJxR8ge9kbhxBA4+rfiB+5k0VAU9h4oXdfKCbSxtWR/N1sF8tdctFPuz9bE
GJRhgjdYQKMiSlNS0cR0x7CoHISIOBsvUnHleZ11FSLIQPOjURDY2Ve+HXrsRr8O
TxnGp68PLuzE82KES2MHjRSesWE70GoqqEB/QiOYjw4nKVTZ3lL8fM4y6AELr3xT
UKqPPtVwbHgxRca+w4w7xEWw6oG+qyA/jFOWtLJl1IT6LyLLps3YjWdz1IFIxZgW
01QS9bIeLxVXgpSmjIlHoVVAilWg0M/cVcP+QoApIMMNbMhFyZFy4z3Vd4aNRgcP
Chcc2c+s1DWaO2bnBwb4T1fxSvDba5Q0ytYHJlrWssMz9S5ECJ3dKwEs6r/MMCoq
L5ih8qhZgdtpoFdvLIcXhaZl6QPZcLZvpr0URLSlw1txAjBF9sBHO/Qwb60i1iRg
fTeQhLZhyvOv1WHR4080APSBoctNqY77hLp8N/jA/9HOBpybIXARcjb6hg6oOBz5
qRBOesf7dxvGV+OqDwf1C2HnDsRKOk+eGuZvATCyF8ZrfF4wTcsa0c2LD6kfQWSs
q/cv8ufQVWBYxl8iwHFndacvrTpSdqOxftcZUk6/lIIVUsdA73YqPSwsWzDGumYb
1s0WXsy73pYC6rNQe24ClQl7xOyk7tzzn6+zcEo/pnk+ynFL/HUuaimgJWLqrxFk
SrVt1R8KUSpsZt98mF+d3V2UMIHLvZeTKaHOiMxxCg2/7w0dM9I+9Oiz6fJZGOKj
wlfP0LIlKyqJ756HDY9rMeYBbletXczFmckQuVXhQg58esN2nq6kP+mTYhZVIF+y
+jMO0S7MrdirBa7iZRIp2tKu8z8hcKlp/7glABdkvDsEQocRJzvqcz8R5Tk9HN24
4XB+G2MK723Czo3sY/gvhPf1nQbS15DCcq3kRjm4B+xRVQdJaZ03MVa5vLPTPY9p
aWarNt7BvExc4EsbyyhYX3OeZBJQ1ppxJQOk3qtEXg3/Byfgmo9SzYaZfbdkcLxk
eTxDfm2Va3R2hapZ9WCzcTGd327IORkyFLL8Ocy2HF4AlOh0VyzNuY0xO7WZUF36
6YXwItjDygBKjd4PCjLYT5htp6r5d2dYG1DYL69+YCIFM20aZozSs+QN88rvYoA3
q49RLCH2p5QdOMhwEJdOy2K716Ta0UwSvJuHYj3/l1f6nJ6GzUKEYKgP3/roTjab
5YJHHKj7SkeGUA+9neaRdQHHSvPVcnT5lEDlUN0jJQu6IGVi7HEJ2fg1T2HMn9nS
73UvRxwmiL3AoaYqwKdMtRsWlAJNcd+9IkROUYljb9xL52HsXGT4IYtvi1R6+2wK
eFzqX6wM/fhB0oHJWVwSTsn4vX0TXUioNkrVW+L5BPhKwvrmlzs9Rkv3BASscIsf
HXQmJg/52PXN/lDXZUFcOsFj3EWYpc3tLfDcZh1egbdoygJq+8hWlrVPSiNat7C1
fn2Vxjc8cRd3pppKbEqk8WBlBwBJ4yTy06SMtds2/1pxXZxrd3em3/Cv+TqgKR3w
QyOJ32dGanWB54UPi7OpS7Z0smpPhsiJ+j+yYdu+qmrT0qvdAyMRnh4ECqZKh6cJ
HEy85uOCJgV2KjC8fI33DXbvZ83kc3akH/TkKJ4o+5KxVAuA1MDGlfG3YRePutQQ
iqNep6MhIS4hst36BmGTHM7IxQ8HgCQNsTsl4kV96qcuQpzoxZT0NILMQ9W7Wv+f
lEas8W2H9ScWf53Az4jW3sRND4SrOW42On/0OtKHiUUxluDHBjJNPSt7Yl0KeqLw
I/VoyEpsWHXj4dqGHXYuI1iD5B5DYWP42gHtJtit8CtpkbO02VBo3lq1zEUQn3I6
b21Z3dZ292DO08Vd1VKLifpqLKIIp3m5YXoPA5Zadp776XGTM94c8Gzko6lWYRyr
4X/8I76BPYN56nzqRIK/epkSHmQ9ug9DS8v9o9kPf1ZlgzVXHBVaCDQK7j5BVLCY
xsef+0WMM36V6t/2UbF4vg3BQOn3rz6NfGv2Bgm/TW7caBG55puUWwOEmmNQ5aUn
dWGJO7zqQB01lQat9A04awdxV+zEm3aAq0BIwQkAshaiu4QDDl50wM9VnNiqCt6b
fow6gWBftQlkyTwSUFQx20FywsOkTsYFnhbTI1hQBjMv1XkmS74L02qgmmfZc5s9
GN4K5TgJ/9PiNQ0/fhZ3T8eoZoAOjqJWD1Jbh61iOU/fc6QmLZfyzD6aRNtPYWdl
NonQHAwXu2ZpDan6Idpca0R6MBi/P93nnXU0SGHtVMphoNtz3ihe4Cn+3LqPFP40
7tGhJMbRTFM3Lzz8jCBeC452idKgU2ELVDQP3wFIf+iZ8jMZOtO76JS9Ki5M3eT4
Ry3Hrn9j10HrP/w5k+m1udw7b04205AHwG5pqD5ilV6TfjlgOrH2m3YSWYMKR5dz
IMkmRM9oFJImY6EtSgC5b+4z5kb9MiEPnYiPzIHBb3GKQHLkIgE+s65AXMseG6cF
7yJI1KmZqAUN1ImsnQ2ZC8vpPrFhmy/dmoNXBUmhMHWivyFP7tQBte2a3+iacIeC
6a4Tf/GFh/pNDZmxZ8h2qipvmkM3M0KmPagBPiCzDuLrQtjtL51I4S6eBUrDzqsP
8XEzEnpBodgx347WNfGXkLrE/FGHz/T+/s85GhUU9kWcIBO8wJcgHNt5mhRz67Np
BAnq9MXoSputmewfuYnrrvzYc/70pNxr9SqIcwjdPvtmMLsyGFjmMHkBJATvZaaj
6IasuJACj9OQekTiXZaqYx0gIv7kCyib/0IwPyHCf4qczQFQLEKnShidZq6jLxfP
kirMkI51l5TPYOjv7L2VhVu1gzvGH2GAbkbmBA35rFas2tv/jDeRBx0KhqYF+fV4
8mW5S+F0EPEpwvZSDi8elAmovZWEJYKp2wQx5EEiGaPAMlvC/xD4x19vhM83f2Dq
ab4uLHJn5i0in64P7cFcNGF4qcm6CmuozLmWUw3EtS8MIPx+/wgMtQPwcnQ4Nygp
SfB430UL9eXNkX1Yvw/HEjIQuTcxorQ6h6faADSU8uyatLqwSJESDUUQ6wlo7cPW
XqEManr1LZTLHlIVsnN3UA6Ut9xrh6w7Vxgld3nCkn1I6WHRCwljLnB9C9MiFeqw
YR9y76siEqukiEofn5giQ77s9m6KBcn0DjrTSUKnmlsPq/UDTYUnV539chAvMHfP
1cOsytyx3AmSPgY0Gy3q6tUIUO03+PuR+9CvQWKPf9g7/ALt0W8smc/xG3p/WMfh
ihD9G+nm9tV0ezvJCcN7u57Fdb3BY44vK2pqpJ5BbmbDR06zuvQr4eNbFFYgguMI
beUn8sm/kdma2rMRRQW2lRwlJ81z1yjAGbHMwPEUbu0Nymw6mKsWMjO0fFGM2S/L
jmeN0X90LCjQMdhy7DqBRUU448EOfzWzWZ8/4BkkRr5uws5zE0OobaNCmps7tz4m
YPVzw7Yn3h8auLIStMaGkVjFQRQjFW21mN08aEekCh9d3rBQdGftfGp6mjDEP4Ks
Umclufhdgl+r5msTnzu93C/dyz39T3Ka6+3r6LmBv/gIrQO5cpdL7HCNIJXGCnhE
27H9BxeD9LDagGET/tg8zJwhY1TeRt+PvfJD+SM42eMfaBb0hm6e2344hQBA5EMB
SERC5UznXrJj8642y19TQtG64XBb0F0NfNk7mFGWaaIB2/iR8Js03VyjoMHtfTf1
dLy3dbsVIH6lNNk6guyVtp6bx9+wHDHiEhicsyXiMO6uiuzPVY75RV8eWIWtndJH
SZsazd99fFG7G+ZQjur22ojdnpKgaazrrJht6d1KRaxfoPoGxQiKmelYq3HCT0BD
SEzJmSFElsbm+dtxi++mKFpsvpZuNFu7zo2sxYxkbvVZyXGo1bVtQuOT0DAnNTkS
V5yjF5NOoTe48/RkgnUM3di/u3GVReOm4Hz1dXmKW86sIm5JKVoGXPzdEa/ls6kT
nPfVuoFiIr0g9E6POcch/EgpUtzw/UyxqCJR8XTGwuwZgR1x5Eqqe7mrl1R90sDz
kufyq3ssZGLK9whlL5LwUHHxgGWF8EsgvJi+v4tFkNa6//dqJOnserqPqOhzUSwI
ecv1/gDHIIz4icwT6yo6KXwk0+393UhVe2CZ1HANIxQb+ZzrRQYkBUQC60gZALn0
OtBWH7DmiQzFfHaAXG2qEOjsQEBjK1dVm2Aibou6xJj840xivCYRD9KKbgLBeP6u
VzHo52BsHG4Ls/EZTU21BRWP39lb0pnCObFKFufhrP+nWlcCfAG72GKo6W2UhS8Z
+rsxzR9ymSDVMq9/vaQU79LcCWYDyxXh8L4T0gHACVJBULONEf1Jrl6Q15FdcOB8
vCnN9qKKWNFY+bS2lQtA7Cx/E3yMOxz/KcOAg/jXjLnXP5YfyiC85U5heVo0FITy
/WUX9WxEIEvxL+mUbAn+smSnY5TIT0qJ3CO2q7tRf3A24r1/slgti88p2ugnHoaG
3cpUvXrwAJDdL7S6F0belFKVc9vZKC7AfB/4nW66hNDYg1Pc0IO5P3ZT3kA1X1ug
5Arp6gsTZc/Z/hzGfJi+omg6skqKuFLgO53LYkDKHtyx+nLLeZhpGStiOcZQUSQH
lwq0rcLtVrAN4u/u3c/GtkDupOyKcC05ZD0LjhT6sW7l0VEMf4VAG+/Lb9C6QUfG
J7IUPYyMNPgcDfYy5tk6/iBKTwt8JmWNqHVKoiBhq+1oT0XlO5TqEaCletjHo/uj
7GfVlOy3t6wIrcZYlubdD9jqA68f8fbtpdkr3wL836TlQc9YeGYIznnxJsMSKrf1
ZJUTO+5+w0LznLJEYJen46MzMEDzP8yvRyAz7CeXyL5GnrxIUZ74Ujytz1WpXA7q
E3JH0sI43BybAWTlRqsIIa+ikldIyv4vGA7nhtzbl2yKy3yUn8D1y9TiPQ2JbzSk
ZJTfBB5I8kmZ55uhQydcPA1ftNbCRbrjC6+Xh25c7YnDHJBIFNZPQ+WTYQlVCri4
WHB/vVOo4Jww6EAoqsooG4qLN1fn18y4/6QvcDb2+W6REd32vb8cwccOPwQgDuJM
HR/H8FEPbgzz5lE2maMxRN5Fy9iG+WAiwd7aEQVvP5yuMkqEauAAqxXwvAwKJXuM
98SiUmpJXN6msBCLG6M+RM2S7WrwvF1mrWHiT+IrF0g2Yq8V5JucPn7YOf+cpeEQ
a7TbZ3WMD6vJ2V95rnsgCeMi8226k9oR9lame9lL+7nrNi3e9C1lUvwLin+JxXrK
FNRK6c7iWcDXBBFebQpl9kvKmbG11ZyRpQ0A/+p2N/R6DZsvZpjrEC5erhL2jfc4
HHY3+iN/t8yRa9RRAfc5+Gk4EIuPF48mYxsY4xgdOkI8uJipAeWRXZBrtifvi/Sr
bVo5nNEKhCOCgpVl2vQhA8pB/m8XFQCfMrEDolndfMi5uimH6nXJrZbWi23lw4sZ
WgO0BGYyBOZSWd1Lk9plYEkC5zdIDfmWzjKtJj3xf5XjPvNnUvSDirueUvYa6byy
bxCdtSQsF3d+fdpzOW8xeuM8suHXqZKpB0iBgG8x2RZgZhF3L6Ixi7qlaMFj+jY4
BnYeHh6zhdSjdAyqxTpuZhEVCJ0KsevPsX2pNAKgoD9E6cJZsUm9n0QZw9bKW+fB
nRjwBJIxUTtcSzfkUQWL73wmuuUc1eui2gKwfJTZvvL/fGIWRo8d8abcIUIdG2L7
oX5whH2QZy6pDyO/ebzhmCVssOpTK0y4hCcax05UkRvxEYmKOy8VGAKAGlnpLLFu
3SS9oDwUEZZbv5G557IpS4/LLgM4kJc3pkATdU9VRYS8ubDxHUREExSZFNlII4XY
i9Fhar7zGqY9cep0KQR5nuYsRMI+AK28D4KmQpMxen7v8kvT2cf+eAksoUf7pgjE
JxNfrgO156mOiZGt7IannIgx9ymA5hiTRKwFuLVlhrX6qn+Mq22IO/rSrJRy6sZP
XassSPXrr2GILq0Cmus3oqVK5gbkHgJXgm/0jTFc1c72Eas7MOdqvD8J0fD0Yp4D
gdQK3QXEf9PgLN0VPglrW0HW98aP2AqoluwMYL7of901HcwZlk1/px5Fqz8qY+9k
lo+fR2/ZMZ3I9DEjxAMYX3fTzEzlkQkmz0BO14SqWpiTQ1Zzts9yjSdlpk3etrMS
2i+vidunpFd3EM9RoKtsV3sp9WxsRJ1a5xjZjz44qRPu4CtiztF1eOquNQ4itqlm
nno1HZKIDTzhNidXY8cv8mJNFPpB+KbZdlPVSJfZKPbfOIPnFGb9tAXDVQy08Spa
cT4doFdpvH1vT3mPk3bsKZhCan7eBoc8lENKnL7hdWLDmhLuOKAGsFe4Cut7fDNq
mZLPMl/or9zQajBHgG6cDPgp+TR6jL1d9QeSkv/LO8SUCWOkwL786P0SEflcxIDu
m5Guwtz4B1zWWHKV5GTXgRcSJJIhhnMVbiHjTsnGKTwlDgRUeCuAUT1n02+LQLQ6
M0bSA900NTaiBdYrGmn0LKhsYlUhdVMcbZSYoxLEf/tMhECXFTZfiwO052DQJdhW
tWCXgaMhUMRS0PeGwT+VPwZzXzYb0VKWjgL9uheotNQRLkd//Te5DN5BDiVSvgJv
df8V8WBK3eaIe8ebLqy/As1n6GT6bgZxgyUuWJpONzZUTtW3957N6e7fv66WmOl+
LmZMx2PPsTh36MQFRKomHa2z11NR1/Sef6SGZBa+znhaPxqRX6VyuRnkVeJ+qfdK
C+xuVQq6/Lf2J8PPhFX9CLfZfDfayyHEUMObqfKPP0wR5OT5tNYDAGXQ3D9Kalc7
JaPpVWSlXFCm1IIu0pW2B1QEWtlMDp/Bc1IiaXV9zNUcjaILxocTDWIm58U1v61d
FNs33vy4ZT+EMwmbit2mKc+6chkqKsUTM/1jLIL/zIcSJES69DarZxup4q7VRvgU
DvhC2xoYW96P8dud4mWPMRYuXF8Gi9vJbR35dusPx8y9pQpRZWM31IZUJHKL7mfM
09UlKAlLwdHT08OJs8wCHTIKglHwXZRYGGyZaDZ2L9m+t4U2iTkmuzoIFFvqai0E
rbJHBuutMNqpHFxvmS8qpWeOmk3NXNy6L/e8Yt2S7S3adVZDabfdQLtQnAxQyHpm
EbatjgpycsMGvmqDpk9EtyVxXw4f+TYZYN2ahLLk+OLUWq/z+Ik3iib1azGsoik0
Q7XpAWGvCyjzjJVjiK3cKAAkGeM0ujG1XcUZfBPGky/71WLGMSs1McXjc8NFktDR
7A6NksxmofzESDOWCTPiBv2jmQsnw308mI6rnnXIfx7N+Y4X3nxvX8GzE4rf8VRv
BSzdqJewKN2J9lzJAUWmgxw12RPENsEeGkCwu1TXKeO7GaI06t49iQEdgaveHLky
oZEfLLtRRD7xc66rdsMQLJ03Fp+PvF1jdEdbgIkHNz7/JmCHxj66AVORkbbv9tPL
WCrzuNp/w/tOyPfo57prrkQM4e7PupSmZm0ADmiHKEKEcTcuajSkBksna1L/s/DA
zn/vUHX77EUHI3021IEJjn1wM4AJQ5gvlPNp9InKH8Hh1dsN+JX4277ggcunuS8F
C8AUOZfF2k+dseB7R5EfB4sc/AbVhhB9K98iePFeaq1tolMwcChiROI8tFDVWb4m
tsLTpYLtLUuY5yV2y/K+IpIl5R6by1Wv/HyRlHRe/b4O0Ow/aYo+5P1zZvcz85G/
jCyZpUYhwMLjDRXIE0iknbe3fIWaRE2Jzt+q8zwlQILarbajgeNJ3vZbUnxZQQch
fUUhVv2y+RdBKBeZaKrPKHRGuo1NpDKNNaatJnusxuNKShgykQ5As3LdUKEvh/aM
4f0AtXvmKcprUgfHOC8A2kaQQM64qXph9AUxSYfSQPrq3VU/JsdYOerX8gpcKym8
giXm7nm/GAdEZV8WzZD8vuiZRJ3f8D6V+vd/RXKktEliuMyD9fP3p/jYSkvRkdmE
+pIiDW/5DWqkVYAm7y5dB2QBSiZwLjp+GBfjEhOTjUOfNWKjKIXFL/jniwxpYVVo
mG8ZaFDxjHSO5FcxA1pgSvzhsX7MqNlM2GAIHn5bnsvlV4kY6uIGEErXq5BzL75X
Rp+yNUQlrJ7Y+CkJJbXc+dfYddN35Sg6d8ViErdMbhPmZaZoJToIf+sp8qHeletC
84hnAXn2h7CDt7Qu0YGie0AI6OLc42oHPyMmKHkeeHpTpbAUaI3W8w8yE5Ga9Y4X
bFJ2XVtoHPXmZa2yJyU0RiWLQl6MzkVpIv17q6Loloq9lzgmN9cqQ69n1IrlOPyn
qMoeH7vWrshyhhb33leEX50zQA7cGQav8NyffS+T+1X4cU5Zn69xV5UfUpdgaoUo
vil5lUbd/u6Psi1yKSqcZMxpTItqYzW53iCQ0hWhvkvVzf2Y9sBBzEf6Zrnqs66V
IVscnjPgqyO2PegYYq/J9/D3lBKeQCuLQlVR6QX3rmM1KPmcq/irB6m7f0aSp3hH
W07+o3FUL5XL/kszc5asqHVXcZhgPuHZ1rq37NC6ekHuPHmPKhgxeIPI0/1CNdyB
8kpfWHCN5IyxdQdvEeQJ3hw6Z2+XojgAOq9EEblVArvJ8nNvktBIjXMJDawne1ie
QrQuIHIqDNPRLsLzSNMJB38ilrN8f3kLrZWiGj9NxxOCVmoWnlM5iIfD8t7H4D8t
vP9fOKX5/sDlmNkpCxjaa/iOXQwQct9ve9M3hv8rMauWtQ7xHikgO/lAqVbhM2WN
IU0JGWb5IdWCm3y7pGUqWHfO2vscYjh9zDaiCH2Y75Ly/e+KGAKuvTO5fxTGBu6X
LMrJ5HvqtvP4aMsaDFinyfT77d/4iBecRHPM0X53blfO027tyysdOFLt6MiywhET
6FhKbnJ4yxDPAm1pE6i7fb8N8AIY40km4jgLeDwcxFdk5LrdgYcKjxNkJIJlxN/O
WEP5JcHSanvPhfwUtI5RUwGDWvxeA6Nma1QvkGPtiAXnQKbCBUfQCKVJhdpmx1yf
yyCvIS8EEDqU/H9W2NGhB/9PcQwvuqeO0HRhyuOQ41CWvCKK97O8cttYJxLlThzE
Xl+rPaCBqv2oMq2y08/C/cJvssvVSd9jNxroO1tzud2QCJuHWIvWH/sW758PuC6x
/h7JXrJrEIwk4dkvnRz8Jt+6PO5grN0M0B7KxQbrIOrIXCoHm4ghKbUpvaT/Y/J6
7l2XfyMbAk/lb3ZxLysKb3awNsNMls+wZkplWK4wbbZpDn9jI4DxYJ+lZg2bTNbI
DW6+NdeBNfiYcRJoNbHW1FOYmWFQzyhHK/AtfsxzB9ia2C8fSgMljOahKyZ6wNlJ
EgXhGqJfG0L2cK+r2a4ryheTvdI3s09k2E4Eb8jAQ12CICHR1eIFpBjWCCmtjQdN
ZKjP94E6kN5MqwQAY/9pCEiDPYMG1wUL2d42O1M24Qe1WG1MaIDAZqnEDMLZFFlz
1S8AQ82+hDuRK5PKi5pfJ9uxc9TAsYKNTcUwt8qLxes12NFugZuMUqksOsdjWO0o
BdqLvypCHP366UtL278CkVLLEpK31n7HJApgx28oeo7xnaP6MMH0ALOjoklJBLrl
2S3W9Q+7rWfXxX4FjY5JDQaCB9ZXu1PmfYaIdneIzJgOBbXW2MXuK2HQr29omuVv
uRTxCU7cjoyGeB+y/iUEtggKKBlTPZ4EH0zWwdT4FZ7oSAmQbNLz2d664IDa23Kj
Zcq8S0Ko6o8wJN4BSdyBkmCJeDbIcEsiItsUPuB4zjTTjY+IaZXEQkz87flRJYHz
ARi6ITUoPFcZBGnrEWr58Jazq/gFhW4HS4iT4gRnZ3l3ptaPRqesbb2TEljih0tE
kmKRaZaVf208G+1uXg7GL2HZKu8kczAr2l0xY5xo4zbny/zbeaYiu5pn3ZqDZnw2
9P7mjCSi7LJY4wgOgJ6HPtYqv/5fgA071qREybnuhkWQHXzEDiZjGIrdjdXGULNv
69PFpvkny+HN3dNIXB75uyrwkAMOXNUqlyuQj3NR4rrHmIUpsb8p88Hq/egg0kku
uBBDwJhhdFKmMKiVpLpT62ApZLzRxQbLojCk9Zssp75TA7CGrtOaGUOi6nSi+34S
W0q4xxz6nE2nNc5KSYGRIZ9f8exrQoB3nVBKmFFYRZuN0e2QslvpOoVxLiCi4WPM
QYRIHuyhNOVM6HOwXrOqepFXF/dujSrUo7LP95AOEZM+8gwiKeid5lBiQuq4DPGn
l9CWfu2CtJDKZh1ggbRQVPEmSrMsY+n8npUCBpy4JWx9+ujMcPK6epqGqM0h4GVi
c/6tEb1SHdZnpxTc84WTHq/CCNTAyVulVurAmFS4RTL9Yanx1UYgCYY6rqn48V1q
6i3IIMdlonUg8uFwPo6VWhDbG80HqK1dJUMyf0Z0nX03Fijodx0FS/UIuzGnwlcV
5mu8XNwOe49BzsXVsaBY0JeIvQ2iPePTOH3tGUArQuQZc1r2UwCbFqdV2mlt1QMK
B2tOTkYRRsC24EIzSghkGtUx0VNtFiPM1qNtyqBojq3dsuGdmH6YhF8qZtoURMeQ
1GvHx2HInGoaP/qYdDaePZCgtpTWgoO5NkODiRSSvo9kYcThglN/TUS7UMkkmq6N
URoYLDi6+O495xcHXaRfBDWfNVbxqxIMBac0RxPT9fd8nnaRQ0JkGKvi4uSRdxZl
n+M7FJkjhGfdR0KwiIRyihGrnquxS6S7IaS1uu2fl6qLsqCc65Y2aES7KgigCvTr
wjQZ+ef6LNN1BtSlLNdmhlf+8FS+SoGxMPj7SlZ7E0t2i76gp+VCPw8EpR4iQW3N
zJdP1J+4pArfAYmoJ+Iz3kesjxFawiZ4ut3vMtLPrBszSCX60GNEKBm4QUAlcxVT
IC2wI+CQHvUMED2YhrBdsivcuUGu/GAe9B7Ou4NYkk3qCjk0ZqnNFCWOER9I/oKE
p9IdvnNlRp7Z5EMivn/1xQ5VEKm9Sz8s0Pjc/yR2V7rYF2ohMHYnMz50RGefUXz0
4oFOHsh7RfgRAY0HvPdMiEYYnDJKkcXpjvVpzIeQfZRFADMVH0La3o4AS12H+d9H
I6gEp/PUO/DRfk/lk72YUDV+/qTWh0Nr31Z7v4YDNoJcc6mnA5txD+M8oNRNV275
6tfejlWWnrOpF3b0KmQg2knkwp6FPG/j5z1iJ+n5zYgU+iqOJffHZP4xeK9W+mWL
nzIlLFIxw6ddor5kvnHW0bqYoB012xKRhxG5UWAyG+iWweUCeuH76bVhznaRNlLt
IhEakHuMf0oubMQUmk+mxDKjd7HLj5fMSAiQyAkiSzhcH8foVysDdyD7qgSSTbpA
5aQIdCz2rlwX1aqw7ZdZwjybxZE8c1WEishB6rXwcNk3GzEiNWHwIBorQaP9Akcc
Mnw4UGAv7CCLB7a04QtXP2FQIV9t1OIrbSLtq0skE+hKwjnxXsXwiq17klr/vrqn
QWpdLBtgPmH8RqWs9onG55VD/gojEw5TVh4VXYY9gTg33San+PG1384mZlZAUCE2
t8HjlbgpnjjQg5kvtbpjWuNTh4Bh1EnLItxfD7bWEAoTQJFwUYDNelfBOgXqhuWF
R6V8CaW5sC2YTBRNSRRMucTD/M/+JkrmhD1WzJJdqxaFalESw/YIRZBqU6vb6VE4
Bl4uFnPbt/UPeah0SzbxZe6z8b2rPPVamiHSqKfmS7kYAIjQ8ryp+rJO863UaXOp
jOHpydIw68ObIDHncVkkaQCAIOSRdjVqjI7bM9Wsk6981aWo2ZSd/UPLQMnCUuUd
WGbAEsgcrzQZCR9kK5B8RsdYQh2WukLQDSq6xwI0/aCp1DEC3Fik5hQlfdsj7pGu
vAbDfHW95lVaFGj2fmMCavrYwxIE0lJa6BRG+OGo6TOQq+ZFsBKAGbqtocaBnJZ5
/0QImj5MQ7e31Lh2RKf43ZOuwqgu7r6f7VbX1HV7PSEQMl39gqrwEG7SV9QBQ95d
K8aXpY9xpPaZ+NX0+CXOrQ0PcwiyzE+C8FD6jV3XNzWEcTnVJABuxuq8UobCb3K5
cp+ouaYEulDcBCxWmFp4nrRHYdNFrT8C5CWVYCWIU0tQhs5X7Q/eqzsrMicpB90L
wcOx6jU/rGIH6ZhfF9y+PpttgAcMgJefJx1ZU0ZsUnP+yryE3aa17s52doUWJHVx
FTBafR2HOM0WZlN6YQhsRy/tLMpQulmq5xoga1zkpnb7I91VQlB2JHYE0NklxNRC
evGRLKhreCvpxTJYzHX+PVd1BSAxJBQD4QeZJt1+5NxHijDraz9yADquWbZdYyyW
Ia8+p3kiLCyM2UI88jojEFSanXTMZ0v3Qrh+Akq9HxYZegBQi7ZkgqsLwR7gT3Pl
2Sv4GdLHwYrDPtSgSyVke2wCPC2qe8wAnKOtH/5KSc9Ql9MiUjG/sesnl5li2e8X
qhUrZenhUbawjwNOHf1icgXqmBEkat6Qrpfub/gEY3RJVzUe2qTrx1syPG0/cUEH
TBYz0sIo+rL1BGyb/YmUKgHxP2CiLemaWGunUekotGkVjNslB63ltjoGp66bTq8y
YPWz51jwIWhTv+3CbX7rny9HPbjorAV3PUDueHxqMlbqgzV77d3BCNKXs9Q6xshJ
W2/FC+eUwW5sLJ0z4QOMcYtNExXQ762ihF+RAl+B2xTFOvThoEpa21bxEeaflRrL
LKtilMPeEPlldmcX+s3EorpU4mNWIiHHDt0avTMNmenm7aTSUgu3s+gNRX6lhn7c
wcZ0qGSWO45nlzrYZAEVQWpqTFRtMd05pVZtPf6p//xTweVaNa0RwSyfJEV8NrgW
zCWvpgvX8bLVowspsFXx6l5zAv8v25jf6a/0+m/1giAGpWXk4DybTMkJxe3Uqbbs
MuawRhpzts/Hw2cx29aBor1elSvklJI9cxGUD1XTl1bxwRMMklW2MUbibOXnUptt
Np9wp4Nwr4AHPd7RyYXrWmUGKDSS83vNttcfcxD0pbPb5YE8iC42HoL2tVcOjIEY
XgLCap+WtCu01C5QAAdeIB/0YcZCIiYh4Sc5hhPy6XVDVza2i12+Ltm0ZPGxd4DJ
OugJKitfw7V5+Vqwm/gh3OGUwrVjvBnMASUjrO//zdM0De0aj2kiRa2e752LZc8u
He19C2GeuiBBk5jucPjummoZG5O95pNsvHYa0GxoPBqtymSMQgcyt0zvFhoIcoyY
npaxN7BEI9SMZDOgeTCT9+odOlrXHfoQGNTsw8rguBb009Zx2IR1qZmL9hkZrqMk
qe8MZ7N+Bm9ces/BBC55nsL91Kpz1uqizNcG8tQabcZuhxW1RWLgX5lz2uM6a8eB
65vOlXRnPA0NiZJRqnUl6p83Om242jn18OIrY+T8gTDuuzRyuzonEfQxiesQ31iF
9v6kifGfyL9xM3EDb/EWmWWbduzYYNAU03OC/2Q572sfJDKCz/BetG5/DYbneM2U
zVhNNNCBCwNX2BEjTHGfD6JhbNID++nfOT5EqDa2+27XDbBwxfKx/YpBtkv+2qbw
Uk74yRwuRlONDpwGwgP0dMLzwGNg1US7S+4vr3ovkqWjV1JUGt5yM/0I9CPj9ByJ
gOZpcEX+9qhQSlW4TC8yzUaYHoQScpYMyrE/ngD7owYQWShajgpQcZI/OXqD/3v/
dtVSwWQ22zlHdCCHDllz2n7MH42B365VxNBrrPFl6yA2jX3Tt08PF1Hzy3fYjc+3
Z6vOV4Fns+M6y163YZv9OPdBbucxb8d9ZQEwCf7wmayO7CjgGwGhaOzdW7hETMqD
EN6MiFAEm0JYlpt6b5ArsjWy9rvzLTAeasqwvvO1zK4I7SQAwTD2AdGFzdZdlOIg
dV8kyzHuvDeOox8+2P9//X1qMtFnrsu+KJQJ1LGExwt0jW4VoXT311Cj/tG/XcEW
0yY7iQrbulQdzdGERBf3O3bJ+ZlyQOpiHfsy5nGN30Ymp045W0d0jF27+mGHMF9t
vL783hUxfQcRzM41Tew+eoeiagctDVMWN4zesuRIxL0hVOd6wc7SJ5TkcvoEslnE
5HmlEMF4AH0ZWkQjCh+h+vMWetq54uexaR9frKtObuEXfzYH3InuJnOdEyLE+vqV
8Si2bTKGyTbyo7j+B5ddvhM/H7Q5KaiHI8Ec+1+mI4OMSlFTKpC6RMX0ohrcCiBN
l8PgXSLbS17spvdtXlCuEFuSn5brBPCoHYZkaiBQXvcLYEEk/BWu6WButBNK0stX
VMCADe9gVlMBeYBxGqWe4FAkT0Ce+60CeiMSy1TwRIEEUmcIHfszSKo6Re5A6sGP
9wcTEBgYTubZRWns7n00cRNlxuxUsabJzaJ6Us4QGqC2jDFbzSkyAXMZ8nP9oK8V
WdBk3tDyiOys/jnuL+x433I/ceVpn4hFy34K46WsHmIYv9wAukD+nrQDeqfdhJNf
K/wGxvLtugOLoHQUov8ewboSfgjBivOn3yCvTJ8l5P/PZaI6UdPR6GSyQFObEPO3
9xi2ZQnj6TVsaBgJed7CgYm/2qqJJy7oGQbpONERz8dupNKZuTc2RTU8iJvqaz87
aQJXNPyLJuFAA6PvCCl3knOVkcBu2X46rIajQzwBUffUqkJM1VfFoZPNdtqbJ9eU
+V6NEWyZ2nbGp4jTEMekzwIpzNGO4Q4EWY59K0gcuOtOkbCg0FD3VRQh5crIWy3D
HJQXo6PlRL2b9VfvhIofsiniBtvBEerOz4Fg9siMucQ5uk9uaVtor5k7XrGsVYFX
yKR8TuUiZYm9q1W15KqbQBXNAdgXtMO3Qa9qlKAjsbdBXJO4HvMMsZvK6X4U0kf/
rz4NccIn4jHG0yGz27USRBl2vn0e1JzGsfXUspmbDJGoy5KQNRTy05bZYggFpnX0
3CzPoP/oiQaaZOIiTZXDLRJrLjfpgW3LmUylMSwns51nuHD6hmFd23KFDqDiN498
iyNdA+Wq84xv0ZtrrO9900bjej4MZPxq+yrq5WXDwPNhglkzKgA6R2llgOr0H8n2
7cSpjMsyTgi7/VdaQh2Ov808WMZyje8PKN4m1t7pAEIvtLZu7fbg7j9zSC7i3HCo
7ijKk72IWh3yE6haP8juJ/JlteLtHbpVvYoZ76Cqjrc9jmhJVpJVRr7Shznyi8H0
mQDTJd3te6Otw9bA5k/uv41pXKl13+mcAHaNRhbKiQyOVeKd6huGtVzt+5Hyc6jR
YJwcf/XqxFA37D26VD/NjsaZelFhIJbfhSWFqsVT7HSMvMbVVVn8S5SlTIwz+dU2
b4eZLqL5aaAJkJK10Zu+rM4/j6DRopjbSphWc5V2VpkvSnBWPe7Ie6tKmzIUgGGe
l1yso1P7dilhS7iX853WOAWNeHxAh4CKjp7jBr1R2fdUY/AwJV9FH3nOQ6rlhixG
xH7JTNOj+FbvW2KTiEAbN5GXUkksPOizgOdD1KYSMoNNbmEIBapMnBYTBV5KvFSX
1xrEkHI4dIUB+8mUTFqFncm2b/XUe2XrjHOQs5SMCqatkLj0h+Zks/ftQFMkRygw
ApVAhK+B/6SoKgsqb4mJG34Yr/Xq1QRVxeIs6q92s+vNjqSpcwqEjEC/qCp0tXZJ
KjPH8/XPkaBaiem0RPE77exxqKnPzSCOMW7FFeP7RP/UVhfUQ7FpSge1Gz5G/gtj
NBQv+FB/wcU71ksjyvqq8X1IPssSc84CgjqjXNRepnxS/VTc/uLQgPJgwDmXtgbv
1rSa0YdmZhzbM6eDekNp+vnXPurRHnSLAsd6lmOawKuhOjJN1lTnNArqguiFmg5o
SZaf6ZbC4dzMc6yuiR685AcvW1iHjqSn3kKUZ+4OC6jEvpUMx3hTUkiLGhx/s11T
Qh6nQ2IDg7vpY4ljoqQVtvGXL+excnu+TtBOe6RJDJUHPMxJA3wkZ6R8ouVNPfNG
AyRs8avgKGDoD5kVbp+9Wi3fnpKG4JJjmv+iuSeIEmNmuCbXI/bYIxHs24kFkpAW
VawIsYvI5uYC63XJJqx0P3+YhWxz7a7sjNOtR5Pfikq9ijU9HG6Tcpw8qjq/Myq0
pjnjB+BmfMOD8pKQ78t3d+8uDNb0JDayyI0gE5UehzvsU1R7vxsnMqykFuNgdoC7
uZvLZzqJja/hxJ6Cp4tucUVCPZ36TbynIfit8GWCXC+h87aUoX+Tl1wd7mCvvl0l
pXA7E++ERO1kSNSnKHtKYV+yibRY+7XiHq7dFRJCtnJgvOyziS33UqPvX9CPeb9h
65ZVlwNHFRcYaktbCe4dDBaSdkUpLFiEA4oq7wvbV8ZCCRFZCA+F85Ya59YLlUgF
YCbAv0X0fTMP4VMB7J/H4WzL9Crc3oKsQp94JoMR/nKHp3tZANYsLKWNZDFvue4b
ssCi1kt6kOUBopWEDTCvgDOHONkACZ9u79a41eGggc6FpHAnHABID4xXp86zlRiL
KTE47AYGFbE5wT0YsugqLTwwqUmbZ70KPqarlhxJdAu35Y+YJtkHCLObMOMiwAfB
beC3PSJ+9Kgugh81dzqpGSi+mSMhCalSSvmyGLROZh5RG2aIjXzTvLjb47IKyvDW
cvsv3yMNaGI9lcByvHHqyZIHgLtQFH8z2CwKMXEsp/dznMC+YsCFwOQNFFBLoHdb
gUMJ8lZtr64lnMpdHsetZCUYWzeEsUhR3Vnb+LQOGPuNGXIr9FY14aVjyCmBgUqL
mTq0qOuGOgk8S52rY7rOO+YCo4kUqaVTCK4JD2AlikpZdH1KexO9xlPngb5BEXtt
/qkIlMzHiy9e7j0APNhrmNog0e0DKvnJTedb6qb39Qfsjp3UxL8Ef7Slww3gaE9T
23ejdxzZZORmM+c3eToif6uvnjbMI44UOKAqeYaD5+07UpR4ZucVV9C1bZfSdwQo
OdU2iexIcl1qO1hqLs/NrLJUt8rNVzuh4CahIPmE4pN3K4zCV0TBbntGw27l3A/T
VxHJDw02593FDL4OdDJ0eIHHFVzawrMAC2eok5WLKZJfw31jJ9+EVqF7ONa7MUU6
9p1VpXDAIW7avsJKF/U4orV1NBWsFVFjad2z1v9vn3kkXn/pkj48SurNC9axf6fr
Dwm0mjp5QUd8g06AAkJo+Chx916xYFvaNr5CHRdc4yFitrzYCqsGd0z1J05unkkd
A6BQWvTZcAHfyznLtACDEQIFcxs+LnWjH59dgVOLvoR0ylH4/3BVPEpOiPSH85o/
EAS2yWgmz26j2m27HzRJV78p3LW1J49awD5+/Lj8OqsQtsGJ5oxZJPBKJANjEWF0
5cf8u482jc6/Jx9QyYu9tgpwCgRPTBdLJGMya4jEOH8VQwPIu2YvpoOCMUf/yi/p
ihgSq+VCrTemVVuYc1s4Z4Y+20N3LkTVmdaeZMjGITSloi/DPRRh5K6gok6dnnKH
xRwjLHuj43uf9+sOgJ6VKonPnjqwo2w9vo/2v3Mi36yygLW9gzmcqbaqYjSx21HG
8D0IDx6mdtX+3N/GmUGcGQggJo5XvGBQCxHY1w6eBpt35duYNNMYhezcFYPCCyIO
pqZ5Y5aizDCttYMRpFZyV1MjzW1rJxy+n4Rpbwtzat8FvYV8tB1u9oIM4rDAPYcu
Vm13jQjv37jLLHpf1L3xxi0l1fM5SAgYMx15QQiFCuL79r9q9U7FBJurnTz1/SpA
XvM7x8vI4wneg+55xaCTJJQ90sKgnGkkrTyaVVxwi1YzM9C1kwG/5N13b4d5Pmol
V5u7rcVehXSBPARK3LHDxuuGry9ea6Lu5LBlyBw6U8Qs3FtI5EbuJBmudAOxQSBz
/TpY7CPtOUFSvBI9fcIL2UXnihSK5Jnv5MJNPI//1E5196pVroJDWx4FmBmZKFTN
OnXeqJfYA4LTA66bKXwuBp7w3yuZqaey8SmvvhkyrjKY5wM3eXh6Ph88a/eVFPQT
Yp2JP5M90E/xNvMhl5sFXivTJkaIw7judLX6tXfISTzi+E9Bxs4piK46uotMrQV7
n2qeqt0hOm4TjjzDEUWIdAOrNCEAhq2oLmaPHBsC7DNS9Kthej4NowmRJ5RsyTMW
+t7kqNNHS5/NdlMlhswBZIuMxr7LSYdF1Ww1IhOJ+Wuu2n4xhkXfOgKSFxB1GSWu
U5kSZjLZFd4LhhnrfrB+mv/nRXidD1cBEqKF1F8/geziYT6wFum0T/n55WfjDNDs
xyKP4BB0pTR1ITTbnDieuuDn9JeUzMETOv9DGWQFIfKMv6r54LssGgAFMrcVWhUp
0srnLuPMsr1sAnmlbmclCepwXVK+74+/1kiZAzzDqOvQdzyyiYlR8yNCKf77GweG
ushakH1Alwe4khFgLGAli4wpzKQj7mggTgkpTF53l8XZxnxuwIjlCSglRva8PrSO
lYMSEVaSD03UsFN4I5UsTzW0GQUiZZm7T2wnZv4uYcZoeWpIVDhB2Nv+fZ98CqXl
PJ/DD7sg2f/slaRIvjyU+/of8E2rsfvaR8/S/eqo5PrQjHkoHpAp43FYHhm+qMOw
Ia3kWN9XHOSdV73EIbULaYihiVQlO3EMvqaKS8vda4uDibZQsjyjWGV4KBJxd2H5
G3VjtcqExFXn/WwonblqJlFynGzrMH4qphtfgnrNuCkAq4hAU3QyV4RAJrwmfsZO
Ez5pBjJc/QvkKnMUCtcieN4D9vhI/5ba0PouiedDyv6vOOCyqVt5/DzM2kY1vdVz
wRLoWTEh+NK1e6dG9VXnGsUpQdk8orFKD93q7ODTDHXheTnuFr8Kz2BkfXxxZqap
cleYS/YUH74LkHsKflttDZ6l3UmbHwaZjiP2p4cR1muxZhMdXEQUVy/Pkc7OdbgL
yPDvcmzrnArrWqtO2BsAG2IyGzic9sNdRFv2tgg+fOM4sfkbFY5KVtZRA725mvA/
CHJ7w1OJDvAoMZqaS9SJS5VjsjcidyQ0aYr5BnVr7RmKW33MgLJcD3kPdbUK7SXz
51CMdf8pIX4bFu+t8vUspuVz84sPB/bFzFR1iWUlCjM2/AhV5YjPhsTbGKbkdAVm
bf0H2acnyin41NnXWHFuPGCCIHkWZpVJxoYjE/iEM0v9qtW4jmZacuLUJquePILE
Otzh9mp2WKpdKBFGG6i6VBviCvWyKjmstg4zAp0n25+GameGDN+vjesA2LmMRle7
uvU9bMxfIVsQoclp3SLGwncOGnniP827Sz4rGSrX/KeQc/vSKSU/inQygN43Uyy5
YeJVszQKg2bU4Gz0qFLhhzdIv3l+mb3H7kFvvjqLHFZEzuWsZShMEFHHgDpHC2US
kJr1bpae/ZPPouYromwlzOpdR++X3fV4gtDwHEvU67tsg+NowQ5039XhSfzDoEEa
mgBBMaef+O2UrxO7Tlg6eAJsaH6LBybeUGrvn9Yfg3GhATZ6KiC2IYLm470QaTLZ
vxE1Sp0ZElp2DEsUugvGzpX/iV6ZN1o8a6rfh3RnTlhqhTgmFhb92weZE5bSPUon
tuDzHCyowlV6BZ/P/xuBveGf2mE6kGa8Fa2GonGuGREEFNmfcsZVmCMo3JnmSzdP
nGSvfJ+cyPjvvfjVi2QNfrHrmkJTuyNiMJT+JJlX1yb67Wk/F5T/TBjNxv7wk4rb
NYsg9m/CxhMGTYDeXYkClK/Br78Hkfo7CQW+2pGeNjz8T52LSUKUjoZJwSsyPKtZ
JTQrBlTKjsfc6kW63Q5gR7guNO0FvAEnhZ5ahf/OsnaIPk82xHNXrbSiOiVW0+xJ
MSXX0FlLCieWD94uRCbZq0oPPmxMDuiLRYuum3wwelkPjFdIHdWD3JUn+fj3c7hv
6EvkPNDLjdJhwRopYzlwwcm8IAXrYQT+eT1SJaRj3vd2QrJKPmEZBLhW1zgYqFVT
Aw4LZ8reZs3y4G7d518i5p1uBorgdXOhMVzY2JqDFGjtrWIeYHn+Tfeyvr+Q8Utj
y0hCCqE/Vsy+fp4YUW8LyMuqHglhztyVSTdHJL5QVInoNeXeGYp9zgrv+VLjEdvs
3qcGGDDAfPFiL4pqNRuWcw==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
l/NRhmV6gxkV9w293qcV4P71DOUR7Uh2mLaUW40cV1aK44p9wcBQB2WqEYsTSw/U
7dckncL8TWnzfaI4zDIxkhR0snE71b5DmMbaIPoeCx+CxX2tWEBs/w5bol3l5nV5
9Y9MJBeguehwpDHqAslqwqkHyOD60AoKbF1BoQbl+t0uPJUoJoPgyd+I0C+CIis9
eJQdwuM5QIRIVB/y4qGJ3ZYnI9SLnSWBqy63aI+kcCr5/kd2SCmORMQieSSFphMG
7c3dDwr/NSC1/9fO0vN+0VFKASeSK3brMOpvCNGjuCe2Ab6VG7XyL0qyCldnvZw/
CmJEXRgAhzrPCbNfQf9T9g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1200 )
`pragma protect data_block
axO/a46jB3+NCtUf2KK+2dVdI8LWmoVjjq45FgfEeqNevz40O7d41LyRjdbVhuZc
beaoAUxLf7Iu36QxSDNgUmqmHYd6U3Dkg51B0evlz10XYhi1WDQzcxpNKbXozuRO
mmhFUWCQdiW63/cTAwRWW2nd2pIhri66EHWHajmNd7m8HhFQ70KjN5VWJpOPUeX+
0nW8ilZT8L4dCdX6yTHbwCP9l2idVgWmY2ZAqC4j3ENaaC1NFmKaEAeCx2MhBjjL
NXKKlxNXYX+arnUGweiC+HS9bCJSZJVGYB00k+oSNRrChZVF5Zl0RcfNyxiatbqK
UudjJGyKrFk5TJEwtt26mRaT6FxlzREDv+mvAuqfWu7YMHaArFsES37y8YMf4NMU
4xRuGuCATrlW+Se0uziBHMs99WQoCb4NZN44NYBwGikN/kyCuoP2TXUvixUIJVNr
yihj8Dz/uD5YC4UoGt7pIET1OeyMaklDwOPap/pYUrSkfK4J2A2HP2L7cqxnx9U7
o/JpkxMg2KoCxytawBls60HrsdAxWe3NaPsbTYyxxD8+E97Wp+dNASs9qKITv4bR
FPwstOrhQlZORwokxXUPzgO4Vz50+ZjND2gccaiSeUSQD4kolDTZ3DDJR0cgHxcV
+M+5H4ssm/ymVJGFb3/H/8f0W8yuBrUJDTBdW1GrVcywdLU+1ttfcNLnkWynVHE3
MP04m4TFBfzGfv0c8TdEV/UC/zH76Sa/LI8ezZHZu9H4UWuo1NVuEnpJTbcX/Wro
aIa2HE5dj5MXKjrBSO/0++CuRJv/ONMjtygkuKd/s/1/z0BKhfUgcs+TsZ4vYJ+q
7kLGyDkl42WLgbb4GUcsC7agLFOgAdpaR+1QTW0s09gHqZXEA4McP9XqDPbCQg/J
xnBeoIu0lZiZ3DJWcr3K32t/vYuHJeP6VeMn3IjOZeh+wkgrAZpBY29hAZho774N
umiXUXaulXUB1eGEn8Sobhp+qxAT2w/aHdlFKtnVtf9VZQqxPeF+VcWKXDRoa4Qo
cU8aIlr2WN2WP9F3AeHEq5NqoEkZGm/RnonokWDlwDzKvwC1aENZcdkRO52pTIRN
WbA/11Ul8y8Mb2pw4PLzTg20KtqN20ecAXYFWREnzMMjWm0yllWxKNSC7DAAEYA9
b0xZ+5HYE1oEp5ruXCBHZK7ZQ9JFataDqKvAWN5li/lL+2ovlGfEG1j1nP+gsM9m
BbSaXXjuvStt58Xb672dKrrK3XFB7edMG8jRscmSl1ZDIU26OzE240JmT+vpXplI
B6sAsGItZOkOWRU0P1nAT1ZMyY20pcpLoaV4bUtjxBAWhrQq6sRmB/E1aDNhe3Py
GQk6A/3+h/HUgqqgP6nCBbM2w2lBRcvl+lnlW3ocgF4s6HIWbh/2PJRD3DnKrSDS
VbbpCyT7khKAxdHm4FA3VATpPDvKjRTxVtLcysEAPNQpB/fJ2o9rZPJxLYhm4iNP
fhQf9Tp33jJALFWShi+nlLEKi2LDYsUInfJxZnnsIUYV31Ivn65N/fW+YFf2nA0O
zjfV44DyjdrHQZ1vbGUW0SyUi8nRsdG1wO3hiyRsyiiPcl9sFQnkHqraumGzTbhg
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SbadBYVlO52/xS5ye3Z9UHUPFfp0Z35scEcQkEzwpCOGIL7o3Djn9Jmtzrr0fpsn
+MEz+/ShbERcGi1kbfGxUjKM6L7FSuX3+3/NM8WSsViFLx7yUeVf+sCe0g6fWYdT
hjcjiRXCq7EdpPlWdWNlch0DDBLjjH57uNvZffJh0dXNa5d8izc+mNWrZhfWKgfU
HeLM0qW9NntQwuOX+9btBdms87Sdm02Fm0tUdvZc+fQ4VJ3i4TCTPgRLdKBitLhO
imxE9fMNcZA9c7pso0eGokHbkyjFlaHBzlAaCyDHOXXdVV69O5sOhR2ILJNGLO2j
rmRh3r2/e/ekkCZZbUfQtA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4672 )
`pragma protect data_block
9cNJ+4GohWArbmcZgn0fag8hES+/LJlY16PHpPZpwcMojK/97HHK9HuIfBwR0+xR
JuD9nOf7NEpgoZXW1TwCZtd715dQsVTmifX86twBjEb0tx7+V+hQtVuIfXAbHnoX
YbgaW8GmECqCj5Z4ftg41HQ+t7N/2Srv8H6nmH61DLAwbhUVjTKuBPudhxRg1OqB
MkOE7dnYAYBMhKBvV0W7mNm8m9+qj8n3fziXSCyufJx2XwnFOH6cljXG3aQ3o91r
h7p1FyOC+pnXmJaeKeRKDezjp7L7RfDy6B3C7Fy4ev7ztp40yTOT400ZY9firHcZ
3N6QEeEdFlCImIpCdazg7CxNMRbNVvf8q9nKP6f3MIIPUx0blSi2b4LZZgjQgZJe
D/rzJHgAMA9CxEa93jR5JXMQtkmtgYIbZKdUTHd9486s9m0cQMtDiCFuxl9eNaY9
0Qov3ryo7bBBLWmZiEMRp7X6oO/I63gV5jac2/V/SKq2Jxwt7FLIsG7FFy4+bsyV
bQHgkxd1TEL0BIfDvng5yN5df6+VgVMD5zkVZgzcVlbhr7ZcVLkhhuboZuE+qygU
LEk1nQN58ZbpSbf4DJsAYwztK3vU/iuG2h79pF9h9dWI0Xl5HQ/AWIu815eGLPRT
t6+722i2uYM+E08PmWJoLAfZD6BzWMRPNgX1fdoh+HjZRuzgKWtyEO3ZrNyK2nLo
f0L6Qw6ZfEUKn/yNI1Akp6xt7f7MYLp5ADlA67DEeRYVaV0yQ6mW6W6TRiMOZTkZ
bj4WsAti/baLUYr7x5sRVzNvd2hw2qQnaJxd5iYCjgjlWvl5rCPbaiFC7M6aWrqs
NtxDRqqbjTV23Aihs5qciazvvTs7GK+g6o3ecE0ML/SiSJu58lZ92lRTl0mfCiS8
/L+XegTOtxIOLUCarKzeHDki5X8fBJsQvtLEY+UgmGxK/HYIU/9/seplKRZ1AXEJ
eY0vCbgMtV6OKMiamU+N1BsUXD1PO0IG/26qIg/3ExKSvX0KQsi6h6sbRSHYLMv1
K/O/0uS718MDX56G/Y5/3dQNZnIUIYEj6gmUYi/HEcZhQ+R6U5hsk80jgMwEs2sF
Fn7bRmYy7aPGQbcP6XuSeZ+9RmhxefeNaYvRqTKOVcTDHTZ1MTV5THQNQlFOQ0Mg
ytaT5OrgHJI+98qhV+MC+f8+P7IXTLUR9MtwzuYFXLA2zRTO/3wOhPoyLlfLepAS
MuQ/kd5lk2WcHWysBqshEi0g2WR63DKKrqdU4oWU842zijUB93OH9lpAWdSA082q
HHHnxuLHE8xqab7yEo5+vWyLYj8qJ3mk1FeId0MeACsC2k/mT3Z83cQU2rA6CL7X
PQ1aEhmHxME2V0VClMKOODhnqTSLQDiyocZ0Cu/bcz0q0CwA0kGCyLqSM4Ar6Oik
TZhsFnHma3faFVKwJq39ZHZkPYZ34pL2nr/G3O9RrnZNFPUsn2UvOTyqrm5lq2cM
f5uqj0dacARzI+sYBVwgumOnIiN70+0h4hi2Utzi+zAYAUW0ZE/bAIwXwmIqVpLi
250RSnLNBBYvDVdjc5tC4o3Vxy0S4hcnDXd0gfSUJ3Y4AtFtjGZTqC4mq0DGx55+
3pAkIeuTZDYLmJqQJglugCZ1vQZ475fdu4NVQvWTK3ApyrpPgtqJlTmSwBJ4SKOV
ZWwnKajrP7Lxy4me39EeyfzAmGG5Ut9Qf/tQ7l0H8SbwIz7aWCzAvHWVmVTFN9m8
DMldgBIqe/Raqw+mReTyF2w4jD0H9YzUSGf2wy39Nep9tdGPIb4FXxD5jO7SlCw2
teMgGSaTeJLRuCfYZj6TgVtlDJWOlYAd8sHf8MWtIa43e34MUIdEJ6SkqotPGVJl
z6pzQIp/4tODRlmX0w/5ae2pIhjEJj54b4N/EPSxZM9EjBq1XFrEvtEDZf0yjBsx
iI9p7WBWLsteCA38MuFOYCxJKHRELLcJUkNKsAe6pukFlKcsW32/b3RWiGSZB6Cj
7ED/rwiRO/cQAH9+lVqfbD1dvEhQO/c/5mIRh39qqL7wkfpWofv+aUE1m2bp9tgD
M0Y50ABdWyyUJgnthKobDw2nP4SZDpVQonF/SeewjZduKqBlgwita2BS5e2KtcUi
mr67Pc4pkc8u7i0It8zecJh51+VZ/uEwjjkh8Px8Rx3KVV2WE5HSj2zELJGt3l6q
W/MFcq3MVrs8YHY6NrP00lQ1bp+/QsE3S4yGjwIUAJLv9fBPT/faePIiz8LIpPCK
50v+R0D1Mjhb8U3mX3xRMtZ7K0FOGDOsXoQdIi9NTLViIm7nwl784lO7E/PtJfP3
3lnJbhr+wi62FgCwYQ7HgoSMjQxyORVNi88hI31PW5qpRBhX0tb2zG5AAwzpSUYM
g+2FdnED0kHpK3AwzqBhRrdenCPCIVtipUFv116XgdcHCMx98X24b5f0DtOU0nyC
wm94kj5sMQIankzDImW0CxQzZltbXCEnTb5yC+7snLWNPKMHLOVf0xoiKljjpPwb
9KTSw5Qa7m8GbjHcwglc5OQjQ58rnq3Rgzp4EBBXWsybTrmVuS/7mwzsK52PF/cq
cq41ClDZVaUom+6AJ1ny1gp2OGaoNvqFqIdhAIPnOp/zMaU9hxvI0/nKbdbeV8o1
0cBwiS4s+Fi3FZjtJghUnX6iB38lKNYIlCyCQY2meLwIxC7MmGOtooxW8PSeklX5
M+VHEtFefA1CRZkyEcY22O0W3tcwWsoXqZ28luDixkQTLf4fxkuAoNh8YnTH6MlE
0MHE2C/v0zT3i1dh0diD2AfTogJ71Ecyyu/i0aZOenw8qDWHKnsh6vebfe0DZlr6
8qnxWtcCQLrbu/b1j3sj4VzAgtBOXH55NvVvOwe3HwTRD1mehGQSKjlj3tIyAy0+
mtljF2Ej3sKzKff1/fePJLCZudLoG/uipIMBtimjduQFR2SUzwCJ8KAC2qZIn6iM
Uh48GpzrAsgrg+Lp8F/gL7qHKnnwfdX4MYtkRH6FWJ01m70QaXCYPLzUGLMIkN+O
+ABazuNazGqCwxqwEh+xIPZPn8X4CUbP3R8xdzPu71dwGyOrFdY/xUca5tdC0LB3
4xvG85aWHHoOtsI2IsVga2AKWXxe8vxqitOhGVxfyjgFxFdzmhsSLlsSbRBPzLus
yDjMINbXg1tiFA6nsfkeCX3ZrBkUTUoWAefSOf1ZGCEjGwxMFAMVJkb5RZ2gxyg3
sUISyfAx45vPjIhiu42wN3z3U0+3Mvsf5GdnFNgaVbfkScTpkaTsr68nHYgP4oxB
7MITFcU37ohPL0f0krLcg12m0/d4aq3QVzPvexN2jQo9zmLWt10TLx40qxN3flQ/
PTQG0zm/pzP48lO7Ra1Xp2nANN3GReV9EkuhdnEDasFhBar5De6vwzyu5KF8heFS
SDivoHUFwU8Joa/mNZ9Tr5dV1IjvjopxExr45nkzsLMlGukSa+V+mQKlYdEIHkn4
+Pf7TenrPGkDbDHFvFnhlv8xBbWeSNFw73rVcj937A4klu3fwTU2MbJuqRFXlvHH
xsEZDwglPMqpyyfSShcQC/nSzx+xELsEuPC6MXs/CnI2o9GNPyvB2YvltBPgkR7Y
6/IySmj+YfjS2bqRML7eLed1ioJOBWASt1ULg4cWIBdx1MQrEhHpPWhNEPQ7vN/7
CEmW9RyeDe61rrTd7qpeptwFz8tvquQqYYOmE9mZFJ32XzBjDBIDg3wB9fVl7kFf
wV43e3RyWqEtbb2QaZH5nGZH/r6C1GF/SFCbEpZMPlCHTj9ZZHaZh2GZRM8hprIP
j2fhzeV2Edf5IJcUxfvYvObGwZuKFawoyzs7SnKxxCfe75Sfw2svaHppflTzogSr
VJJ/GWoowS60+WlV9lhtvF2l+RIbYOKxRUCI1m+d4Hpv6oOHjgcNn1Qz2LCGgB/7
kIQ1i6o+4+2WZ3NrBxD3rNFeBJk21y+25o5rl+QVEn63ow3HffZZQmAIiUkWou5K
FtOkj9hSaHEIWOSZBmYoGGnx50Ve6rwb6NMH72Bx5BZ62p7VBqMoiWLqtCnHZUO9
EqTG5J9M0Qx8vaZQmX2DP7GTPIPfnc1JtflpTcRKnJDw1aBcA/+SSxLFVwGWjoQc
WZblJeEdDgUoACzmrscfM9JxzC1RN12amDKDo2YJFmaCPmm6IpIvGgi7grTCj7KY
P4aJT4WdWlKVsLZDtCWJb40NCh4nm6er5TsIBF9OBkni3dxHgTXjdEwGt1bEjGy7
v6K535ykneSetdMUgtycWZXe99JFdGq82sv8UaBrL/gYtny3UxpZB+YzrA8Fe8SX
4wZCRa3KNPaeIi90IHK1akAw0O26B5oZLz+oGZxoj/hlVhWAqjZFagG2cGlHoo7Q
4W1fmxAPoZpEVtDP0vEWgdnxpJwCK2Cb7x6M/eEBNsPUkWrNhuebBcOk9kKl7jb/
RRGU4yiuGyygQu6jOnIFec0Ho5LZA157RTWsIli8aTRiyBu3wQw2ULmEU66vYRS7
jnFvSlaCBReyCZCgtPyO5quKWJncoiiae+wIX5aZ67GmX+fG3TCAR+cvFnwYiMd5
zxsmlPYRiD7Ryk2x2jw+qDZHjGZ79CMFOzqr0LprrEQ/iAF+DVGb/qlr6mohVvLj
gWxAGbx4Lr73a9XtrzSO39MJlTIvYTTCyO16N6scWE5DmDd8XcPJHUX9uBBAEMIJ
EhrNa996Gr+nJDDpByTI/NGMuRv8wuLLJYRe7vgEw/n/3i5kU4mngp9PRerkMY4j
kARSi3lGmBk67ZxZ78w9Rw8uNwherk8occThtghw+xOC8/hRZ1sP0EzzdZN2o02w
iqUMJnYCuQNFY2M4OoDLwFROMBrBotraIdXBGfZ0flCio+JB0IStzMVTT8k6KT2+
dVVELPbRLf/wVQAq30EHHZwk2BrQ3uDLAsNrFfLZlBjHuVsIy4jtzCl7y77lBWsn
+6NA3lNxUlxcIsn8gW/4bhOhU7tEjP90jVhOdXIyorEtY/yPFP12hLpNNdTv53RK
wgmddosAa5N0kFQpiK27a9HVvquH6p/uPnbTdA0GzCxT0nxEWvxhmcDGrnRLsenK
yzMvkXCLYedkAtIJJtXiRIUZwYwxBlyl8pYLhUMVdIybWVBRt+xiVAtnyZ//udQ/
y55futY+AQqpysghbe5gx+mRa+4dBb+jM4+0qxQOnBn7msy20F78OiAS+Tg44l7d
mJFoM8MgLfd4C6AmDwjNb4VeeosCR+xRcYhsPJEAcXxOqrGYnRVSUJwN4nXa8yrQ
TKMPzrARzV/MDmg1azpi4hE6dB87bShBWdni5n9rFQd3tEhebys1X9iJZX8hQdlm
BwqbBrNlYinuuN5Jt+WbdB8Tf1TUElfVN/dWMvDy+mLNcB1MO+5uApiLMFn+X67x
yLRxkv4spFEojth2GJnQ+KjopbyuhBFyihwEynpfb94pMOG+AAIS97BkDxES95eV
SDGIKzt4I+tApAanrg1TkmmOaUrvtSS7yslSfZfd56Jltdx4/V3ys4A/HlZIFU2z
/DdwLLHf9j/3LQmmwwg6ahEDgPSMWPy6i/cH9I2pqfbNdWBOMh9E9vlbtfOemx4G
gIqCNQ6lfgZkfZrRlidyKEmpWls8yg/A1liNnzy0WtxTYuOdYoQCbKLLscQ3NXmL
S/0Cf5YqxnlseFAP/2QJXgnaabe67vz0BD2oBjOKZQ3Xcv0Rkv1z/EJYMqEW123p
PW7za+e8wduyTHMqJueFulrvBsViv1mNy0bqwVJ+EGGd7CUGPKRt6laTTePhunkA
m2c0tZw4YaO76NTmnF3FcMVC3XVg6OPSbO6wH1WXNk7o+vYf5TlUKftIYyC2vCRV
ulECifxab1lq4mrctk+Gf06UbNZPloujITK2MwBMjj+y2ofB+m6AXq4+A5gMxVoN
K+WAoywnytgPGr5ODnIEDqwMtW93S2L07W1z/qLDqLwzn62RVrjnAM9PtBIbsWrT
3Gf95cm4SFyihqIzPY3fXRcvMIbWdK6LlP+cZym4XbyzeAjgYnuyV+hLIHOKqmfq
9yUj+BnHsqCOhmDmlYIniJiJ6/6oXu+X/lCGkLarKOAsPwIDdHcmU0Q4mtaEdTiv
p9K2czh4PvNLTqPcVC31UCcO216UYILVjfetTSqiO/Kg0IEWTT4+jRgZd0tGo2na
19NmkkvnA1Q2HXlzc9yPhyDIjMBhfWRbxiMURJgxgqAVdrY9fDGAcf0I7ZXHXvv6
N2wnYRxtRfTjtMP1jMwSPA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
N7TqNZWF5Z0F3H3q42vMyUL8ft7sIZQvS6IzpCoun0JacDtljOL/ZL/8M7TqnBiW
qI2syXr3mvzoa5z8XDA8MScs2gDjmXLyYFxV082+pWG5E8QesANdF1xYwcN872Mz
2RnWjYIYErs+uD6TpP06MeIm+RQXHQcMe4pZEDkmsQzqMk3gz27XMLmRv1kkseD1
RUF8B/BQiasB32T2vdr3x3iEhhqmDc6o2CKIX53s2GtyiPtHpeH2AegJYYGKPptl
7cAaa9mudErHCWgFgRBG5Bdcjr2jnHBppcVv4WdvJUG2m3I4wsYmqOw3nQLn6RZJ
WWT5Xva2ZkDua8YP7LKcjA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9344 )
`pragma protect data_block
2Hr5G1dQe75EiXjEBG2nh7VS/jiO46gxqbbGDcXlnCwqGp+XC1jvddFrT/CsbKKw
oY/JWpTWVG1yt6M2agyMeOIBEIPqJJWqBnUg8TL+jFJWtggP7JNQD2rZHFhDkfEU
CsFVKktaWTqhZKvoD3ICvDJQWj0JR3e/ODf/2vlreOiTikrPRmP+FluGrsEQOFhv
EkQBpNbxUUu/tyfZC3JOjCKqnSuxpaqkE69zRBfUhseB5tpcrh7dwyvjU18bP+1v
cKWHrx/qu/hEMboBevvKZglYH3SuVVl2D6By+incSM8+EdXl1LbmzkAROjHSsmKO
Sc+VjrfoPaADhHzzpxlqcMhmFJBnlznmijwu+Ed3DZnJ6hWan38KMtrJxvuvQ5pv
P4MyU8BI4PVQSnpBUmUSsp5hWNSpSDhTbsbaiaaxt0/tw6TfL/heYtUxf1On0wlB
1bAFxQHBJxAivIY7SaO0xF/W3GeSzweZXGBrab9knm5qnD047qntF0e+yYFBZYbE
BEUgpUPGi0+VI8XblcBRbQ1h09R2Sjd8O3ZPY+fJBJl2pt1WngFbtu9Js4lyu5jW
pWU5YTuqL9saBJklgqvmmHTXwGzceymnfaJm8BEIP/2HvwZgX+2FVYc9sOY9RDRI
dsWLgZsjGijer4NOYQM3T0NpIhOwtJpXPeOAM2HR6gg4WIgZOkv+o/gPPNH59xMP
wg1CT1rAzowd+Zxeu7fph5S9wE2Sqt9YSY/KGEiUvIj40gk2xQqf95XSI1iyHclC
//FlS7kYj2NGN34kZdohkkw84uhynJCzp7bH7fv4xPx5KyyDg2uagbYjkxn4VADd
kI8zlsOqrJK6erHXZUdMC/TbA3ex4C9aRwDkGUMkosRyZ8OQH63qok0RlBaV/sCk
yJpNAEzUVUQRu1LJ9kz6MTNbii9qRUiOx4nQPl+/CD+NI0fDqsCrdqgfmJESOtJU
Xpb8xSfwlFxNB6cU0APYl3O2hqTNh45BLJTs79EVjwM7dFWpSov4z/ah2dj2rjjx
nUnZ6J88uIvt4jtLmL72z3VVvnkiyicGStj2ZPs5aoCWPGh69/X+29G4sHuOIO25
btObMDMsWLgsCZuAJ04xHLT0RgvfTeMdXoZ+nlscShnlKvhodtvL+rozsjAoX7ZL
1G9oiKd0dzMGFlybPfkdugehvu5SbGHJ7OgRQd+UGvGURkEEgl/d87/MyAg5e2RW
0nso4EnyEkl5GvRjYfmDv+ckdxTTQEA46UEzxUFWphS0v1OPH76JY7ogUki+H/B/
EfL4dQdicUeIXxo1FuxsRcXZXsq9lZ83uAphsg3wh83TDIRCR3a4Vp+9WF0Ko+z2
VxBD69hbm6Wt1EZSo5CcCS6FGzReJTM4mU2dV98Tgtq8GBwvHFn3Yj7SUPJ9iFH6
4c/bqJRArfPTnYWYrzdS+IyHttU5E2WPgUhp7r3PGAvH79xuEoqaFo/aeK4yLyfv
lo25suH1aQ7fCV4CIM8edj7iL6CRtaGc65II8ox/+dcBTq0XUeZCV/NNlJIsNHbw
5UiCTGQJsni5wvxHLacIWc7tvpBYk4oCF+/bmiLtUPszlZv9v07VZIKHCHKUapTU
2/SR+ErUFcvKMf8RXhuy7x+84T/QVrXnMxaSocN5cr1k2y0xSoLVEz2wMpmKsV/5
vIEP3W+Lq/E28d1So0K00E/q8chjxaMt3tSQNZpE6MjnDIVs94dpsJdRzxVlB/R6
JCVErhY0O4cRZmxwgsrE9r17AeYo4AlpcENiZhKH25QflnW7O6yV4gzf2UElw1bW
7KwAs/9DuQVKtYoWBcDzIJ74ZLlLTSEJzNnfUyQSen4hJS/UhXMvxse2BFq5FbWZ
hz3K2MT21fHy6QRXlfwMZdx4onT0p40tgLKD6SOomRen/tGTSi2xSp1SWmkOl6If
yDy+kaI03RVX8TWSTXYgumNmO2dqCFGKYFYBQp+b+Uai55IFA/b3GZeml/l1mEKF
m/4rwdagWt7qZ5QMtaYx9U+vh/WJi+LdPYL1yOIqT7EbpDglkuS6DYicAmBsVoDR
GKIH4hdDwHEKuqQnJf+jTM6LZDEpea3zYaNIoIiqnAh1Ls4BDFIF1xOo+9MMUOkC
6FtKxY99Uh8uxUH/WIpdzAHP7ZRRXzkKPHxmN+PUlDbbfl/Hly1fj6qn/XreP/AC
XXfwCillCS+HvlwcBjMdKojD9LMand+uKi1wfeBikaj49RcmKalTnJUpDCk9yMPP
MmrPhFf908ZGmmJ10/yF589CsudqEQASPrFr5TFmYUeJZci6TWb/K4uFkE4mg0sf
PDIpS/eJiI8u3JxwYDL8/VcDQZN7DVJDhagI31ZtYrb6hZe6lXfT5jB0hYiNblsf
J0YfCOgyLSjyUlRjMsdTYQ2vrn8sthYp30RHUp1jduG8E942lF6VJOPM6BW6qiaP
mLRY+WDQ9h4dTS6h8GCxOvoLguAXkh/mACWeuwFdc2F49iV0FlcSMgF+DjRzR06k
IcqES2h25kCumnoTqj/PxGmQNoGvYbVFYRfQzqc0UkMr23rXPI+J+sVEWY77coAs
UWR9V9BRSWfWcP5VDGSNvYnLtLjTZE0JtRD5NONG3lMU0BDotmXaSguo+pwfxpYY
f79EXYQG6KEneLICL5gvq8z40F7GWMh4q+6wRJj0pMvH9PmbEWsxwBbCgL966Ts2
ZVq2sQi609WI5NzBHoFEX20o15//jq3SkLaeJRe/c64lozLdc5BaJtQd8/UInP64
gkWIs/voju78XJtiZnegA9icH7xk+wIlRHFWWVjqBOkv7EDk7BQEmCbDK/r4dT45
mhBxM3H3Qqm9Z+sz1+F+B0/iTEu/OjFbe4HmtxtJhO5u/njczkOYTHw4wsTP8KyQ
6vRzKsRzS2aRB0LPnmnDIiHXnIfFQa5ImSS5tvHReVSkCGla6kIMNnepd1JZTnv3
fMn0g8zjTjm13k9bLXJy89kIS33aBu41qNlkhT1Iun8m6RsE3Z/NvCxmgXxGMv21
s4joX3Jeptbt3loOGGPp/t0+zqrFI7ofR5/J2B8nd400Zk/d8rR8F/GPVbvyCe4p
VadCBpxJI3U/NWPrsJcxwaG9cnJ1GKJ8Dx/jISnaF5EIun+U8ikYlNXIS29zvp0D
D0rIFUz2rsr8SEIOcF2afmL2La2bG7CFsodovcQPAVY6dyIH9EWsti6HymhXW5xQ
0jV/bb7fN8XysbrZLUgjV1nxEJpRdnga5W6i62jdS8DU+GjPV0YIi7v0IFxHe7Bf
Rp5gMfDkiR5Q2+RMfGSSrkkS+2a42Blt/+reElETvdWwAS8SDNNVaVObqBhB3MA4
bzUPveuR6fheqGc0sJDmgrPrfYuTmnL3ExWZobWhaNduhfLxRUebjB+Pxy8Gn5e4
0FjDg6aLr0DyYHgOx9Eesg8sKIYOGtwvpRCX+GgJg7HW5h3VFuSxdf4msuwfBJaj
n02FxatSC1PkVpRwp+Wkr0lwf5VLypVkErFYZz+hFZIsFknBTlwUXIAhKzfFwDS5
WPmrHH/fYqr6rukLnBVEtddtmtX9c2uS9e6CUP+2y88sCZTx+Neq73HhRFAXW8mv
Qgw8ENDLCSNCb9b5lafrrn9oLjqAzJKgIA5EoZeFBhlzmE4/+q5psYlbnXsj1ZyY
LQQpJTUd3DrY6Cf8HJXPT+o0XZCiwsNmpRf9zvaKKY1dWajr3aiQ6RWxYGnWeQMY
tVTdwCdR9wzn86B3FfhRhqQFi5AQlxHMANZ6CHpkUTLb9VTgZ+xQ5M97hNd397xf
KsOpa3KGgrXgyaUeR/NLwu7TLuBffHzjN6awbb1XAn6qD6XEC7fALKCd8qzHmiWO
hpqvNrVWwzcTnJEUXoVJ4ZIjQxFS2JtSg3yPkIYpa9BJ9HJ20ocZNdQ2fApsAhpR
OhrrhsRLbUmAph5lviTVpkeTenWgVl0lQBkihDks/+j3Ko3fsWphOHnYgXC1i5EC
lAC2aGNTQ7DgVWnbA2nXfoV6cKqjqmm5CUqkH0AbOxqZ6I0K7ZAB2r1F8FVNHn5y
3W9DYUNG2Ypgg4Pdxl7dlj7AQ8HCo7qWMU833Hs5LgIK80TTyZmhv6JIKaYr8dF4
fRDm/y1rj/1ZrZb81EoF3YLk6XYUCbqfttmTRZ8Ttqx58nQaHbb12IenRVdnoKxn
nWcGeUc0EoNxQO+Bh7bYPvB6thv2TWRPPr7DxFovIG9aHg+z4AnSZL3iNp4EYfNK
kNj3vzSAAXyBJ8iTiHenVqB+KkZZdi6gKaAbAreC0F3VXAndk/lMZYDllNpz5/go
V22ZdIFTo9uM7KmTSS2CEub0qkgY2VDjM5OIMk1/raFaQDMCG0LUx6XeuGezU5D8
VL+z1AmEsQiZ/RgSxxRU6jcJid3DU/aqueuI0xh1xnh+yvzFuQ76p3mc82qp/vFa
8/9xLqqkXDj+mv1qw+g+G5jXR7GHfVCT1xpE+7htQ6npYe0P75plysiq/DrM/v0h
JaYwC/VJgSJga11IeJNxYsQdIK0oIKOdYjFiNf4Gh5EhBYwpvQ9wZTmVI/34MrkM
T641sdjE4ozyKgt6r1b8LGIp7Uei5VO6sDEG3UuzBhN8jXk+TLyyY7lUqXua+6tI
QrWNDt0CSxpiALecMLC5p9TpjYOyUfAzbB+Z80enccgjbUpqHJuyXHwmvWZlH3pX
qLnZIrYItTCI3pbrwVPS35+rKEZ2ze84B9YIChbAuoiDtakwZhlDWoMhMTImhQKT
WHzYnTJFPrH/2PZUIt5qzP6bBXebh5lmAQLTegkeuKf9roa6qCYIGIQl3LMyspLm
Mw6D7AeRVrZMNWKCWku/hyKuz6dbxhqYaqrlKRZkewOHhTLtVzLGceU8UfxaswD5
Avk9764ZNAObam4rCHcTRSBEf+M7Ovwxuzhpt9nRhVZyUiBlhAWBrAkknhA4D/t2
inTnKK3vo48f2aKYOv/0yiP2Sj1evqAPWYgPT2FBw0y7F3NA1MeKa7/Vn3rjB/nL
xPaK+gEEF3YEQG73ARt0cCYk+URLRVuDVcbwe+TH3GK3Lmu97YpdON6GGbiBfDBV
rcUM/wDdaT/PzvVPutmFtHOqSyQtN3YzoltL1DYCu7mabiojyJrcQG2luC3Pva4r
psOv2s6LcvRt/R2PI9qSD2gErPYS21LICjpSn8uKJOB56PdTxuqaFvIQnW59LqJp
KyrmAPEbCldlw/WAP4/rdcyPHkcPRfnoLeV+QCr13Q1/KOjpdGy0hH4Ef+wgASlH
tNkrdQp6mpYBQByVbgccRSrQnwPEtCSuyJnSrtbO+L3aS6APKVLidtUU23m3xhMa
tGCCAADKhE4wpIg1oECvS8WbmRs41gpsfATeugreZydUD2XuomkT6io8HNugcQJD
Re8VV5HUHAbwZ5oOeVLVFWpgjEOT1iZD4aV49JB5x2ZmOG78mo6DsPxhe7wahNYy
x1nA/NJVWbREDL/Bl+8E0Cac9MXHDVStiqNbIETB0aajTLKNce9qpGbOojVwYas6
Iz/Wx78wsSPY8FvLJcDAuSOuz9mFtTQwnuQ3R6/kegZl3UBj430nvPRm5x5GRiBU
LNcg/2rlgVolVJJ5sZO05HLTes9j+2O0eQOFLuiigDMQCTk3UggbWV023neMuAB1
yf2FhGHPauXalZcv1u5p6Ht10RWDJB55QULt+JDzv6F2ZhyFqwrNW6F5xGqjN2GL
Il2DW/79zC/6oc2ZEImMAy+M23ALEdXq3gURjZlKYDu62c642Zp6o/lJPNhts330
l2KIUJl22Cg5fuOAkM/g46Ts7qrF/LKTzv7QeRfKIu5LH/SGknHLOdIyChUvQj4P
tLSZprcXMEtUOxWTs9DBsssxkl9p4V+CgoHw0oKETksHy1MPreP7R+KM0mFiSjKP
I87D4guufx3qokOIhRjw5LcIM+TXtQ+LVeZzxpGryWPtBRVW+Y3jtkmENTpEPng/
zvGDpLbZ2QW6xOb+5D0rYOyKgcyGMOegmfag2/jAXrfhK5XyKcqQ+97vbFp2/pVx
qwINhLWIg8NERsjtkYkHzKwCrHshxSmU9TRnm3Uykz+lKDMCPW63wZ+5Ws4OykQf
PaLcHeA3+bMxnHXXjq8vjRuisfXXm2Da86YpTHkie2VmF6NWdMhPRS/+NpcoTMRl
Vs+9wECt9b7z8TiMz1IARKhrClAyKC5lrTK5mrolkCHcr1cmtxWMjb5ueR6272Ps
uVkN+E0CPVBVdu4rWsi47EGC/eTUJwKdcG1UmuwqOxhPaydfvZJ+Kk/YNA+xWPPf
SFZFlsuGA1r7LGjSgPDatyd2aS6NRkZ9Dm/0yS2mV/xs3TBGS6krJw/S2a1taWIY
S8VEh2utSIXLU4zPonGbovdASv5GcWhbl0x0fQW+WQImHDY8AXi2sFpqQMNquPWh
btaJWw74/oNuBNShHZda3UgRM00XVanZgkS3LbsPw8Hs1mex95zBfOkrdDRB7Aau
JwMw5qEi2ZQrThRvpVViIjwua3CDtB9YkE2/tHoHpG4HiQRYM12MP2nuKJp53/U9
BQoeC2tUEsA5nfHRpBm9gBmYolEIbfQ1tyt0ZesDaRpIPsCe983+WvBlHE2/cj2t
cqK5pbMpWkliYQr4lABOjDZEW2mxW3GgoiSHMhNscC8d9/sI7t3P1Nl8iLkmo6hB
54dPLegLUv76E375wcSy/hYvlLIZNc9AGCB/ymkgCV5Q2nawzqoAwUQq+SlF90ah
6wD9DRNjq2SN8uJvu8jqIKkpqkZCU5Ffg06favP9rNSvl6hCzvnPKRzAQw/dTww9
Ur9geQJ7MQtNQBCSaWyK17FwKu3HxPfjydz7ozOCQsHZJa8hmXHQF0/lC/GEOPWc
Z9fvFZ4Pe52An0eN/M0xlNWNZmfMnDSLxZfMW2F74jNIX6EQMP8fp9NSkL1EG3Aa
odHxfoKxLQ3sh36mNekNRlR54T6m1f4v8BXjj1hKfg4Jmu0ejThfgGWZEwch8CL6
hoYihwab48NTYDDr0vf/6GvJKikVHj5R0ossnXbt0oU0Isa4fFMxHyTo335eh4tH
V8++BjsqLDlKtZ7ehF+yZabC8I9F1mvmd/gYTSMJOOglRCs/ZsOCxpTCjAA8bzIp
mmBNt3QWVdegAUt2gZf90AGcemssT5HdZ+uqMnWzmMg5fAKvt7wcH6LMITT/K7F4
4tSLyEBP4TEffnRUNx+Fz522MDaHD/4de1yQ+5wigTIinD5zA66qP0mpPlum4BkF
bBRKrloyiwhj5meEgQfCFJGLH8WcWnwLNai1WyrOwpPa9SwAyCjtuhqVddsl9exM
UP1FpNq9d6sx33j3ibYPodtmg0UjfGtTk50sh6erVKlPlY7pPmdXPB3J104AXHXD
viscfLdOTa0yQAySscrscO8blBQUql9kffUUZ11oUghjR1ovuJUj0h38Zd99dbim
k4TPNlWqvfFIQ6ltId4HFXkEzjM59H2g2TLMwENRk0r1g5j1GlSNckNA9uJJ4wjO
uUUapnN4ApDXKcQ0rZRV8MLwp2qkvLmZ2wM4QR+0Ctid1liiRpJ19Vhcnat1bsdi
rfLQ4WwIodGpbEa/ZtD+Gr2w13mg+jfvjinsmTmftdUSYsSuQRMb1wws01qkSAul
z7v8Hh8AthZskpDBdoyPwOQ2R+F3sb15wlQdqrqT4qULS58MEP0IZOWHM+hUGKyz
t1mkc4inttx5HsVMTmocBUYNAx7RvhvmL4mN+ceKzWqdIO1G/tMfwLuuVxCjfc/J
GHKNnhSSluOuPqcn7fjH17qRa1WOgwn3MlzuFp7Sv6netVfMLMMmWECZJMoUOk5I
y24Rpqsl25azFJLZqRaoVEb8WiZ152xipkPK+rbOj4bJ/Lt+xbmpoBnYwGrlDIJz
LPr05w4QX1xB8aRrqlfw4qIumU70oficomHijBSPioh8wagDvfU4u5PRXzuFxAQk
9D0617OCsfY4PUaUgtNSZzumlgcZLuzz3emi0pviNvAVif8MEHJIvaRUcEt8DUe/
DXGrLA8P2jTYmegf/Fr6TvqX70N/hRjyEXzVOvSF/ldmQIVvtaCTcqKpns9v88yY
37Ptx99YOW15FQMDGpoCxo4mjuS/QORKWu+FzVTQ+2++ZjaSIxGW0bjB3TdjUgT+
ZIDvx9I3DVEAWaZwPyyobsATCJcnupCM7I2V0ZgGDvX0JTRSwORRyBibPgX/vY8/
5JtqvNVHTqSWEK4UqMFCD9pEODkHuf8tPUuER9u+3w6VV/Mg7OyOvb1+h/68FK7y
x+CskG6sU0X3C/gEggLFcZDdsR2VOjVc8XYECIMTbevoQr76rRApp43y5WS87wCm
FjIe+noGOZ8ZhUlWCCbXmNG/hvtvbllLu5Et366ceiCC09+N/UvUP6jEKnqNxYyE
y/w225DTtPk0NHpd2fL2+KrUcQwyIFmllieGdh8bLri7RiFaHLyKRKupb0gh9V6c
KWgAg9RZtSYDpld3OTmj9G8ASpS8/qhCV8pSKrW0cWeBMf7qcn2DaKvvMGz2oyVb
jhyNSqrgZTz9YE7j6GrzUH37pUrp9QO0oO9syrw66psaySU1tj4R16xeB9kzWLFJ
EVRd0aeze/QUzlIHhkbC1rrAQZI4PDL9Tx/wK0XjPIiIb8ulgMwBMyIUZDVVxSXh
qrBRU2fRrHW4GC/V1V5M6OiKvQM5TnHrmnZ5/O36l/SX5wHe5OIVtB1Gkydjc9OJ
3+jM5U/gGZi65AD9uKTFnH9TdcWrc39C/kzuneQEBNlGJ6plxk4Phm2c9KiExHcq
nE7VZqSlI/5RkBneAFFeUWZNz8uMzYwaWktQ+rMz815o2CAeCq/2xghP7GglrEOz
chj2Uat0kwYNFswUc80/V2OaBB4fPKf4RZ2HNjQR2+8DpZWSfUNCgF+DddcXYu0/
62r9aZjkf6tQhSIZGcLJDDeX5wDoJJZE0Squ8ZU4qTplJHlp4OM9KQJFcCvd44og
iPwXJg3xIN8qlC3lWXAK9vW2uHjNhJGHzyg2QZ1Gzt/S2eTZ6TbACgIauXTgQulo
9lIt2TtqTW2fdbfGe1u5mIdXvLVoykb5w1dWSW5xLsGJ68GVZyKXBLCYB7WVqfmP
3yC/XSq0z/G2XkLZh5s2TrGmg1u7XiZi5fyZDQpwL0QA2WP28JY5KCcOELUGoP04
8TOJ/wN+B0JGzLe80b/zueHmr4PJfyb7bBacSrsCfbzBMpI9kaG+up6RQmhIIYBb
IUXQc6sVICYPi7wsTQN9KOQgIRP+nhjiUW++WZReCP+DskBpJqvxOndGFc1/b1of
rC8A5KdxZphFwxjn5F9vlCg58yfWKAwH6EGvGZ1LdoZOrdlj5UxaFQIaNK56Rnhy
4/m161w7H9sSHFyQVg9F5eSCNtGy/oABZbVsZJeoIrVZ7KEWywTu5UE4/duDVKu2
lDjaWlXu2njqirhfnqioaEYQhfhzD8BAOpkNZbFMkFJR8UjXMObXdhmZd6p4x+Ob
NN/pqJruGfEw2fj/BPUzsSG32/NnlthHwgJRECNz2bjV7Wdhm0wifX0Se5wMSkDd
Z8HqjqedW0a3MLnxZHFIl03M7yneqQ93CNhAH8ObWk5FrdifKML+tDNzpK7eRrxl
XSnvb6YJi99bJh3uIQvs55dLuhu52YMacWLlCR7bOtqZhaT4W/gf4HunMijd/JCp
QT5P7lh1LdA4I2eiuCOPgtIWGrqEgbS4QZp0yGyz3JWaxuXC8AQe3G0ouV/nKWXr
9663JhD04qE7z16EZr7gjgKXKAybCsDKZtYgX0+7RLelwkeg3EtgQrYofTGgl4vj
00k1katnjz2SM6wwClwvKMaRgwzalt4LA/W5feHb6TPX2pBpF4rqRGypzb5Y8ftp
q/U1N/bq9j/I+hGHLYsj0ibg+HeIG3i72omex8uSLEgR8s5Sl+3mim+woamH4vYy
qkxjhu7RgnKnH1OTZqctNguEeMppHpmMIDTt+LLB8QuMH02dwm5iCD4LkMPVoc56
whQixNGk3A2yjfCU4HxGmZiFM+HqTx6kov4pBQIFhiRu9Vq8KCTqChmOh/1NXk2K
IynjVsBQn+xsDl6qdWha+1dCpgiG7HN4niA6gbj/NSxyNGRDfkXA5ADjTRlFhr3/
rzgQINZqtcO5UQr3XEGrob8tAIQGOBY7iM3pBTCuRFlDIrCjChvAQ1P7w2iZ7bUk
9Dx+as9bDd7s/qqstIUse2BtzbdzPZe41w98oY0cDmVwTuo4BT+o1xXGVuhqKgAk
TafqOw/5OpvSEsvkFGgLh1LlmOFHc/0+7CewVady2bj+GGgTUXhHAo4rlD28HGVy
F1PC5vZyvTCh2/C2bcAcpaNsoWqub+bZTYbc/zCT/+yrFGdJUArI/kx94t9OW8dH
eTE57TAH1IyT7NzPs/X83A6vGcdV+9PTfZykhyvw2+p6kGyrpXLIA8QrXcV/mVmE
egizBKUF5tFeZ9gRLMk1gU9np+HgtIcD8pLJXstJimjzhIUc34lVuYjMjIIEPOFz
FfNJo1GmveMafgAyQ7C0VMgtqLUSDVIWH1ODKNQJsxOA6m4ioQX98XMGRBmBS1b9
qL9VvQ8j3TNy3gWEN7BidL6tJAplV0EPVOWojMmKPo4MX+jzauJvjxYG6YJbHZAN
j7yMETd9a2QwPP5ZBBHQCsa90gc5SpZW4BCyrGCNZ1J5767l/Yj2hQpb2dJ/PUtA
Lgdpz3p6nr0rr0GLF2dxv7CrjZBYhbh9UA2TbFemAY5euAPPoBqtx33tdDY2YAjd
RjWJtdYvmrlPwdHMo0QTb+NRYbPsez9DegsgwkvfwIISU6zI9TookxtxT/CZSK7Z
4bohfMsoP4Nha1Su1tSy7dQmqhcc/lnq7i6awVebF0aS2FLJ3cKR4V/2yd82f7ox
T0IRcxliX2Cf55H+SYuO9bH3CoehMNbdsQPf6SqU4pUoBN9es363AzxwMz4kacPp
4R27ftSls5COaq4QxNchdH2tZAaMdAuufvhnl7blTTk+N9hq5NY+AOTR4ECjR5Yo
cdJzI+r//Uo9wXADjGiVncBh/zFxn7e5SNADJBexJQrdN+0IJY0Bk+fiB5l1KU4v
DZWqZIgwPvfvH2eliVDJV3NDHh9VUzDG3o7+TRe+4MdWe125/m4fsn40hcK66tFs
MyZw0E3fRMEdt25ipAofbbpFEZf4NOWMrDalhV+aIbVq3OEqPAybAY3bd6V1rw+6
S8M5Ii0ZCkjPRqBw70fsRPL2yVUsoO+DI4+5DB+9wDrgBStOvzDndV/9gw3Y2lqK
V3HZeo2UDolTQ6qNIgkGYSmdUoag8zBLaPxNnfbUDAy35SkasioThmGsSdH6VWEG
aWrSYVNroDPEmNRThqz6MvzsVITKR0lPMrj8FxIF6ffNNkGWmqYW1Z1HgjEc4Xvj
YHZP2/vFWNHg5plaGlpeGDUg1MMAm1YpeKOVWImfF7XBgqSxrZD8/+tOxpOS46Rq
wSun0TNf1Z02pe1J84TTdV9HHV/xSm2U53wjq3RtDLpB4PJ0/D/tbLwGCuqj3h5B
2Sc/TzOpv/FqD4G4vumz3VC73+jG12AytJUMMnb5ouZZdrHacm3m/rUcn2fe59v5
IM0ivWMDWeVIQ3ArWZfyh6kn/uo3aDAWhmnQx4tAJbULbVbQQKPile1LszYzLiLI
PSuQu+GiWw3tudzeNG73rKbdr/MJXTaojsTTikJGuLjZHpHsAmNDyo3dVmS7/Rix
Up3akepbZVT7d/Fcx3EC3eXXnDX31yYKbKjtGJvavo+7rGDm2WluiS5P6uDK7YOC
tascJ8MgZfUnI3QqNso/X6GRtMg5+B7TUKSGZ2m/tZlExIxJoYKqlBCY69aa7u6Q
qY+zkMl7XgHlyFiPeCS56BXF+9dz+sXzNFVYWQlKqyrrmd70N7wyAZd0oVyKtHBe
g31ug37jQxDOMVKbhgqws0Qc/eolGtI2AI+P494iwzhKf1dvj5PxsEbdvmIBniNd
RLN6AN7t0ZN2neW2SL/RozgbI9IZRIDSFnPqQM9kjiOCCxAuAbxlkpBq+mQkuubZ
MdZVwBl83D9NfXoUi/uddK1l+6rJWTwlQIRfuAjW0dsHoJCHASHpKxr4i9RV+cC1
gWxBkxl8trj3TEo7PPmZL3liGx5PimCkIdgxwuZJZn9JadLHft5pkOwIXl+ykoCX
qmVxVn+DbSHLkcSeUOOzDJDO7atpPY7ZgLv1O1G2lXvQhZyl4sLj5ASlvjGnKgf6
sgDvWqSM8LQHBspfuO4WT3SNKEa7PBWgswZtpknGtBRFWsO/e98Q2ZtMTaMWv3qQ
XwXXae8xgIieten3kX6OCyXCLg67ETYqWIA5ltjjWMLSNTAM1s30zZW85wiRh0la
zCCO7nOEzpBVMWjpA2xrwVU5SQckMeI/YSHDv+qWMKXMgIZM7OksF2DdxuIksRhd
Xdw0iOsoQs8KO1JdF1zbCZwNhufSfbq84MualPoSSZA=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nORgtpVyo18u0Oh10DB5pjZfRU1fiZutl1KufWR7txBoLqoXC7JMHV1Qahxfhmrc
w30whXNoNe9aJM07T1WPfiWDK/t6sUYhza+6y7dLSRo6wfoiWWUAHr5jRhZBrWlU
n0HjbYikURc3aE7wd1Z0YQAFJOZFbFTRahP9cA4D8xMGeY+/sv+hI4hWq66crvRE
lOb3RBCFSsfapv20U7qtEJyMAXicLe2+Yu7zZewpmT9g6tg/fg17SofFh18znO+W
tHKqVUT7oI+MirTLH/8fGWnoRJ67vsvn+jxwbyy4dbB3snKgWplg8de5PykyYblo
d9ey1zWdIAx4+ipj/Uqxrw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
HRZivxlwAxl7sFLSjVQrXajp0Lzkn9qJDbBz6prU8ZKozFRl/d8SGtbmCU3fM3W1
ZUQDX5PuNAXwzsPBR2zqxVldDUxfmXDI/EkgeM14vh7bSDgstXvhChBfAOVu/sK0
mRFLqOBaR4k3sYjedEC4y7WyvvxxtXs78mdXoe/5rcxmPL1zUzruRT+n6IIJjEYP
XX2kpLAhylZctAqLF70iG2fC4wj1UyK9v6FPg5raWiVDCHR8UKpi7B/BSKSl211g
mXtg8ebLW8G6gRbVxVQa4o4DFU/y9qm/yvv88aK+5OQM262zi57H7WhVpRaXnkEz
gUhIR1yeXE0yTmJsxu9YMWOAyvPdhlV1r2J+PetELqU9vgoccqVGKJdBJoNgKWMR
ylRYcbyetgSroF3ByWIVY/0lYhQ6kV4j5/UJ3tPINxHJkxUnnwTS3ym1qZhsiE31
siEM8rqthQ83GRU91/nF42MMp3bv+hO8hX0AHJKAQcptyDJUqnJp0r2D5jb9Hf/d
aZfhTbxmlgRM125lH8qKBGszmlbWftI4DvHXAFwPuILzbJ8pBNj3X3wvUe3rAIXe
W57d7PB0uLIGTmJRDrGwS2lzSWWV13FVil3Mf6+C6ye4BmyepjdhewM1yAtHuZ8O
tXZa7wVDFfEXm71Gezpd0EG2KvW6UN4zsJDahFi9eR6V+UjTZEaygjfpP7PTMkpZ
AHiVlrHDUDxbq5TDlwEe6yp8cYSRENa8ncTeDH4hOz4BfvsKUEEDu4wGXG2HX+GN
BeKtwVDCy/ygvhdD8mRcXv3OZgyvRWs1KhfjKw3umLelVeB0gK1qEEHYqJM3xDg4
wKEOs0QZsy4XINL8hUe6PhuUtrWMt6qsYl0UmitgPS5s4rSiLNdHWfaF9UTzAojx
pBSdPH30kxQnSKPzbOH6D8Lt3jc7vb2eVHy9zeohiq1e9+WljBVC3syG5M4NIpt8
Q9Zit6K4nP1hdH3k4u1pM6rJPf6g8ompQTvLv8ZoL169W5ZxWSYjuYe/N7FcVSB2
uFTXl1inQTOJNcfwSGqBCtsNx7TT/xlAiHwLFo8GNsJRFsx1X7LYY99NLH7Fmfa1
uiZn0g2GAa3hzncCbcS0fkEFZ/KCpALkBadrWnsg3Bo9HUvEjZNdAzh1mqNhYW5Y
Kr59Z29QrUo3pnoBpnhMmG4I3meFZO1+bZ6sH/7haPltIinlg1vNaxUc7pxuYtPm
lezmxWuAk0yPHdyDNFmwymeG9YjhbHTXb/FP4aBwYRTTUahtV1bz/ULdfvNPowkK
C0grSn15flhmd/RgdoZItWd3AnFr4h3KS5syuhT1BkLXSwPhrV8+zBwBvrHIBTzL
fkxRBhO6JyIeltUtttL3oslzgXavyeh/Adui2ci7nmWaobCl7E7uI8M4ZnOk3KGa
kCbk8ZKxFStYTQyD//5gZHqvWzPY3lqZofzZs+dDgrzO2ZAdJFuzMpYdqdLF1XNM
xnMAP1Zx1i9bg3/tM2lSB+Gt5k0fmHefR33M9QNWZqgW82bAZtvYQL94jdSHaEOS
gvE03oUW3F00nKLVYFq/QeqhN/BJqp7LapXRtNLDCvWo74aziZgHu7LwTklUL8Rz
2FnoHksCTFxLxpB+ZVD0IXOZ4r7Bd3IWGWQ6NQsP0c1Ld2BRSzKHebMFmqjJG0O7
+vHOUifxnz949TOs93KGRBlGm+KSEJLERIW0JSJIVzFJX/d3y7eUrHoFKg6Vd488
6+b2qiLBo0qHeZ5s/8FAYHkRJAx9pEVQCuXNvxAt2Qf3kTwd7Eq5ApotKBuAIntN
+/KJtM6McYk7GvrqIOC7BqIDNanteC/Jn49ksRJM35xwGsLiSkccZ9hSwer2KbLz
PaZ1PNYeyZLhvGycmnhx5b2JsTOimgG7m7Pt304wsVKuj1rDQQPuN1T2I8vidUc8
C2xA9Ux+yB082QK1gq+aeZ79+ci7n69r7GSmpGpXlvW/WlE8Fj4APs0PcnMWhLZT
vA7AtR1Zpw18z7y8EryIPN3mhMPeondmGx4pzZuKKhqK+sGwqmx5OJdbm38mVj0Q
+ZE6XohSSLmtNR/duWu5VtKAK3n1jr+lhYxkd7O3S8hEqvfJqknOj5PAIVHtfk9o
XpcccP4AL00Qcm1Al/JlxCdCKTwj3JoJe2O4VIxYLwcY5RG82PzE0ya7U2DaATe0
pNwOmrFokTPzuMnFaicyywd00EL0VinODY8tNVhXmNPA+ZGxNoretOjrqxqpaJ44
1s5voA68w64hr7GBn42X0wCQuXfygI4CRHGxrV80D8BfOxw1J4bl2BC8WNBnpjUI
7R2ci05Z/VdoPGev0a1HS/E6xVQzcH2t34UbQPJdU9ierr3xCxOnkeyr4GkqBsFn
+UjoaDNkQZdHpY15blBRpisgU5dX+/4ZEkTA42EjrLREv60lga5zuXcD7zaeQEO0
6WPQzqaEREr7YIyDZKZnYJ0pmSP0seuvRYxmet0ifK0AdAoiuMhywAdFj4nRcjI6
Ybx3Il1t3E+sFDS1qqMOacu7AnLpThcad4QbWGFrudR1XaerrEQ7+Ce6oCyDl6YM
3w3ACYwaa+RGBavQXAiicnBZkeadLAW3Ql3HjYd+WT4KNexhqEFyXKFQa+ovLp94
dZGsU1hn6NpaPcUFeW/+FCzNmkEL74WbnlfaFtEsxGGppxOV2uKK7uKmSSTjUE3m
nryRg0/jRKiql0h41lsLZBHTZl3TPLm5QMhxmoUd7AATJZKqXDSV+lE577Wd9I2n
S/i+pjOCo4A8twocIsw7gCRBymi+hBtM5OwU0gFEq4SouG3Bl2CgEROHsR88YQoe
CIEGlmYONNexo3e84Ena9rXYSqEASYXFUVV3rdpHPibLsyctmJ767uqoj+w+fYyo
qnVTG01vxObhNjNiUDvPc4OyGimWNJjjpsXzy0Ulzop3v/WHK59nuCZddqfs5ZJP
RDksou7bKbxPQogOLbfTIU81dzpu3jI7RdEvAUG1qHM3B/pTqf/6AwX0sVL94pu0
ZdArNcYzLXGX+IGsu7X7MEW/ydAPE4mtqFJnXSvrqUKjAa1yo9sI9YNxBULG3Br3
PJ/GgiXfWFcgWNRTvSkB/IdZ2Ki+DU6+5bBOaYavyl71YMGMMMrHGfDM2YeT6Nnj
MehSEYoLeOH7l/T4ZGiIwI8afi8HoiBXpWnh5M0k88jjHkOYKYc6pijQzL4s/Tto
WN1quqgWAgBVe2odfdiY/0VJv7QiSz2b3xZPIi5VkF2lrkO1Qw9M6aQkTUpRBj7q
/Aq7azcAOIrZcwkwWDwPyzZp1VOblRps89Df94x8yhg0d/hfD86TeC5mmy0PL91i
tN3oHvwkg33y1BvLIk8kxVd7pFi72wiwr4U8VsSbvJUubBfY6w4Xu7/5CfPKqf8z
NiRm9Zx07WJuu87/nAYCvvlVYhksCPvDfuWkrZULQhNNEvcNh/LsMDq0OwML5N1q
u3s2tOWS0sCo5+NR5bupfKibzvM8LD9j/EORI4Q/ZypfrWqiuOsjsrQ7kpyCn8wT
RtTQdp8bD4pgB4IiKaYZefffPiz1/WCxQdag2/Jeptc4kYPU63bifp/gnTyaUkjZ
9kR/w/oFPJ8YGyvqte3soXtpyo2peJwJMtrjFNgFwqYY+hyp5jslrwv4e80vIJbM
KShy9gI+XXyEqmSpKUVSrRil+1NJ0KqKzM+9xrplHMaHv16tROYb+2oSWI4qq8S0
9DO6c3f5YToXFmA154Owv6B63CfSqgtqsS36zDrFfSBWm4iB+8RpswT0sIEgewnS
5FF9jnCCx5ENm2w8uOnFWlcQ1RNE22NCu3sudDldJyjDkbLCd3FzrCPmrJFTUdIY
XfhCuqFhm+ZHkwlpiU6rcjdBHNNm5jl0VdjfUKXHOFHCbkqQPN0b4IcWpPoPx/9y
tCBdGIbchPwT+gP+vEOOTQCDOIhJ/VynjsM4CVLxOn7a/mlUrUDTAggxORUbgfqD
gIm61MMKoUc3gsPxIAAi956rNxS219U8kN+K7pGcGodKLXbosfVZUPl5up7Kbwnx
HDlMGqVHDBRbLyfemQWB55UFrPUEahGKseQUaxt3HqB3AWmHCygH8puCna6LFQFE
Rt9J2SWbHuA3bTYILaFUVJcj6siNoWQjr/dD5gKqF/cTc7kbQNba8TOhI2ZIzbDM
epC07cwGOG1I8lU1RMg9SFm3sDMZkjrU8DOhksBoIgmOmhMgKs1TM0d86dY8cxvA
CTwcOlf0O8Gz0Ymvn/xUZkBkp9ExICyTurbk+IZTQoXdEoJ9dI4vJnZzi+GzcnTu
0QR25wGc7mQ6xDbGTtUuMLTJVKzs7Dhqs7VL6mGxYTDaO4NxQu556VIG5c/rY4Zg
NqHDIC6fJ90XnF6b3VCprihrKap/oa/KEk2LKTHMX1aOXiVAna4upZfQvZSP2ErM
CPGmjz+lbYqAXbF24k7xfOlrlAyAV/cTlo7/2ygAAUJxgky2aiX5xqrRuh+L6g44
GJlMgvKrXDn8gFyK3895OWYRcCDq078M7waWu0kwG+kNaOSVuNBTQ6z100Km4Nh8
sfB5SF70leRILkQXaVyvuPvGhaC5/mqKpTio1FlLOQBxd/I5YCk9aWaOhDQJrAPO
FPPsxvjL2n7Qxrk1OHfXXFQXWGIprhA3Ee8rayfymioCWt5MP7D/rtnvmf5isRsI
AX0N38SegIhcU/ZiSm34r6G1J3rNW6thBahq5reWTVwxKVu0blWz9fm9NSihfKOt
Oezv9Y2OLsWPBGjvNZdb2MC96JTnorJjRc7Ig/DUyjPSwgri/mjON/g2bEv002BY
/C4aClxBKM5PIKZ5Njd2cLvwWNiNyvAF9mzeytOXSCJr8WXqFiCd7Qu47tCrRGqm
eEpgc6KChhBn6FRk9yGm+qZy49ZTndCa8W71mK8f225ZUMm/x6xKycCbHFxI7UQG
pSIlMAJHVWxYqnWqK4o0iBISvkpZanbPxk9pKci30KVvpZeQgsFzHSNOuuL3/8i7
gA/363vX7KDPIznW+u+R+jQEKdXz37ksp35bA+zN063nEB1LVBdK4uLcbGdU0Eum
hb8cXfjw0iMAI3+IlSOgN0PHy5SpAWHKdOvVf4/6pA6aiAgdzwcKPomRukLkvwYb
HL94bDDSimm6/wLb3/2GhzYwGoFj9zuNJMuIIAMfXhfkCgBFYlgAmD2bf5ptxtI+
aP+u9MGFMn0wbyJ3hz0//4ItJgalXirh7T89FLmGhxqOxxTp4+LrXHYArfX6yQMU
QcTS7CXrWzrqs5pLbzuoDETW0BOGT9qcJ2QIm1Zl0N4w098JOHuyVOHKTc2pk7Nl
jUk5rtQ1vv3v0xZy0DFXLor8fIafGtGRN/8LXGUZOvmKmXjWQeqkGdw8gRvVay2o
xV2ng7QVRBStYVBhZjdSfWbAtjiHj35lWDcidWcl7ziguzGwW9XT4FgSk7xyj+W0
VgGyaqhh/NAdR+8nmezrlSkyrKtsRv3ARnyNdv3QnumxTMf3fyWx7rXvSuXrx4vS
pi4qaa8sw0VJjLKHmKoXFKeU+N3GOO+jsmhm5KUg/isiLnx10TRo1yhJw3y4QMRc
WCw7gCWyngGf0sV+wzliU8dTHovBIEK10ikYo1gTxYKdtwdCE2bkaZ0jfhbOXmHL
5AjO4h/tp7zsTSghQLqx9nsF0s63e8vsOnIx+LixsXlIR1hSEzI6YILa7jtLNAYf
Q5KpoeHjNRTT4ex6A8CmQ8PwSMm+gjR+JcFweO74Xs/7ZoNNPXI4Cfp8cfE+Dfjf
Lq9ZzLm0kPbzlVUu7nDwLhVGtsGwse57kCu8DltIJHNHrKV4EMo5Cf+gI5kD77h0
Ud+x/2dS6SH9OAh5Ae8frLHIHJ+6As0pU159LIkWxkdLHKUo4ZIJ8RZCu6yU/oO5
cZ26anooIPBzGzVBMlhMXhshw6yU1EaxVIu/Hiin1+97HtpbHUt8QkeSjSFjXbA5
HMJx3h4PcUf+C3FOX2OmJeKdyjlgF3rRtEMAn8ofzEZ2EQYDl6JOzFieN1eEUtRw
YD35R5BK0Vl1/RZ2DW0NgG8zdqgS9csb2mu/pXneWgRBk4w1i57i4bcS5QEJ7oAZ
EAuTR1+x0GFpL1jC53M/ocrsZPg7qXn7qBn8kwQR7ycpLN++mpkuFF2SY58cC1UX
smYR2Vmqr0RSaYlRR6/A2yEv5Eky6xx+wzpqOt+TyblYqGS6D0UkQ4MUwJXPRvFN
kjz4vaX/Mi+KAjEZqb8B0Tun2NikoSlvbOtdSoGgTv10njFcSha3zYsXQ9EIEKC2
N3Aki5A6dKwL3voHA5VN9tP0Em09s4w9dKNJQBS1X7BAwAO5klUiWByOeDV7T8F5
IRKl3XT+mPHpPZwmE7SsdAkDZyBmjFDDnp5dnTpbJbUgIETBibNyd6A+spCc1d+n
5VwvgcRjM/TXXnRLMtzZAjT7PrdeD567DK0WVvyQWiB35tu9slBNKwYobULu2eRP
Bq7UMRphtJprWq8ma3CdELI47UtW+987m7B4Ox7Y17lMDlS6/+NLfmC4yq+5SnM0
bfZgwt579QyHo1zBM5rUhkm7YXuNhSxsiUQTMNilpP6fEFBMaQYRpp6Njbjo4VIp
xh/Y8ex45mZqr7sQWqf5jzUd4bYMA2J6gzCKjuTDsHbRcyqXeSJnnmpliDdWibqL
/PQS3rPKEiaUBK39BbVw2K9lqDgn4n6NcN+C9WJmIhr6vLJUyBZ6H0+E60x/Khsu
OAJZYs0hTOxcx5ZU9/lV1Yo4u5DDQuqZI63QJip8V45UJ8g2kw3TXsQvVs85hzjc
4kk7ZA1Zi+It3KkqJXX5JC+kdGK/9Fnx2NqQzU+Z98mBUyw+AMX/enmBCQgex8/w
jFPJe+6VUvzpZ7hCDkBCj81mH0A/z+IH9UEtwhJdfsdDWpTP5xlI65KxH5ZgAs58
5KqAD8lFSYLs0FiUuEIkhbBHCYDTZAHDiPmb3ZgCv77jWMqlFLbWc9v06374Ysan
jvigrTLc+ZIhqiNP+FVsZSt2HbP/ueYc3i8SgrMC3fGmS8r0ygS8IzyMSIrSXSub
DCrCAti4LIvK4CS0Ov2S3Rhv2OeqgULD+XJK8ruEwTqhq821CKAEZdbsfbmqfOwb
A8tlfr9VLzMDS12QfO8WS/0c5s+EBNo4FGeCr5j6XUqExV3RYL3IyufQUo75aRM/
37trlbijbO7T53NQw1j6nZCVCDpZV8RGGv5QgeN17gdpPpSOhF/T1Rccxr1GDf2M
4uCaY06HVfBnYqSVDkQKrjuEyiTghHt1PcTnW2qjiefatCL4yWxDIa+bR6eRVvqp
cC3jRmWgGBKk5wQZmFJKZ947KgrWcUhL43gQGKzuO3TOSpT9A8annoRKp68oBO5g
UDr58FEWM1Hw8BI1yZ/6ljTOMIbB/oZGBgQR6/j7EWP9/ECpaLLpWiVU9fPsSyco
X13kn6Q6CJ0+pUdRUOuwiIGeh+B8+xKUFTsZaxRZfRw7wacsq4/0gh2FaDcwNdzs
L+53lzf0ibQRGvsM0iJ0W7Jzx1wsri6KG/8wn/kLMgUZm1j79MiIabEzmJterYjP
YZPfPxaY8pM5E7s95Jafj3M9aymnaMubKVsPKnFEZ4GN6bjUCL8BuNLxIku80Qjm
kemupsELYLR6nNXAhlWEDPoRo4bGSSqhfEHr6JdrSzp7H4dolSkLCfIRU4DdU9IX
Z6V8Cc3qwoj2ASM7yn9ADQeEbr8M29LuunrsvPeAGrA1CvdGQNNlLZdmUAVBG36D
RCToMM4lw7WyYzyTIvu8/G20S5d8vxpy+EAEjCImjSrs9WySEok5jy0fCosqUIoA
gSR8MF8OE06leL4vLHBBrs86YJ6XGD1EIdfIvN2mzlogcdhBz6BMQmkofKVvTQMm
NqOgi3AJWcQSuzLpO13cd0T8t7Uppoa+uf+UoC9fDwBeXCvSqQW7+12p7Ub/ECcR
YIa9A1gkyvav3AlPRZI/6nrDakuPa/7D04DyDe/tTCPGcdiqZLwLo8bmX9srqtTZ
APB64xRwYkcqs2S+OhG7O/Ph/N+Z0or76Ky6+6goymCAOxcKoo7LIREuDwfZiEUr
WqOivFRNBs5baINZLuPTk3spTeyI/KvTasGt12QOKQvn6C0IspRttalIV4AhTigB
4VkCdx+sfcpjutQsZrhZQ+pugcux375FZg+B4KyHJ0me2CFi2zjDiO6ZOOGnh7oB
izbKbfVsFg9dksUHIPolgvYFVRlz6QV/5s0IaXmwMBGjB4sdCMsqFejuNYTesX+G
pyZ1KBXaNrqNPZDjCe3oEeqoVZDbiSb2R2fz0+/Zg0w5HZe+Rd40dpHt7N5YAnN/
FTu8EP/Mir0Wvs+s/0a1atu8CtceC0ba3CFIpu54hl/ZFNh99DGVMW8oId41dyKX
xyqT6l18QLeUSnfRz9SNyzElqcrL0b58io/Hx+2rS6AsCxW3X8vSHMsJfjWuEzSg
lzCmouKbGecC5nD1bvAxSYSVxlrl/+CGClcJ2SLn5u55n5FbfzpseOnTFerfj2RQ
MHC7zyYDjjxvZ9MPKD8FR+bA9rvsW7QjtjpKreflKf+OHchAEhhFJEPvmjMpZH+s
qnBdg8HEzBCvTp/WfJm2SfmVeTZTJMR8+4G2t0MPqxzhVYAxnrhBNS+ezKBpvq71
4enDhpKGEBTuWF65PoxmfpHjg4xBNgdXMZaMsiCdDvBZALN1xFQLHOnlhSVv3CD3
6DzEWlkE6iOEd1zauglR3SKsJOWcZ20STpv1Wa70any79xWE05IS9zY3sxVrE0kZ
+vE8En8KTAqbE8xpWRHc9I2bngYS+13fHcfLd+WNJW/5OnDaqMuxWvIro/0e4Dn0
eoKklqTgF6P2YN0mRd/D6UFkhuh0/zM1kTZboF5ykit6tRgpVwwKw7yUULHJuooz
ZrLr8tNLxGS7wiHxzlHoOvV6Glx5ChDmhRsBpPR7641gisMAqA+DPl0XTcVUm6e4
ZB4BzSlfMJ/uJ2L/Ru43krBwm7zvfRIA4yAm7wxkzxUl8FjK65zvdJVd5HykzMCW
+qT1U3C/BwHms+lTx7g7rqzu/i5hWl6+sJ9Mdfzs/yJcBj2pKapfa31aUZw39E6f
B+XyO7FiCUiQH2aw8Ot8XP6zIfpanzjq6BSzt+ZmTMtlbMjZ24xDuJKxGPMvYRr1
H1m1ueQ1uhh9ghqctDdBgHmhJQAF9XSV+1VMMiBUxS5SvRkLRYwBkpYwTJsSR6uF
CJVhHcbywBhYF5/8pAjROfQ1Wr3Rxz2Cy/ErhlTrKRK1Rg5FiuGFKiIG/ltp0kWE
HrtRDTtKKdqUQ1pHW6Wt+N/y8CK24fXG2z3wGaWgFxbSS8/sXmb8UtvToyeUbsk4
V0BItOt+K6Z1sZdvS5eBnhsi4akzseTVixpERlyP1DflD1tbpQjeei3wcwFmqh1e
g1IAvySaticcIEm/BkR0URTXAuxgc6UeU/W5Xi+Uh+jO0p/hANiObAH9vgJNSdMU
qQ46KgcD2YhpwjAFHQszfvh5MeTyJBly5yne0kDDGQt9dOOaD++P+qTC7wpxXYFF
NxD/b9KzfqYbtMfEOxenbSD/AaEBbS1Gifup/Z4lybsrJh2/fdtmAy+OBJquEP6S
uEc5hYuhhoUKnaE/lzLq4Z2jk3Sa6JITM4vQSaPtXJz9WRX9xzPwTsdxs33PsP02
KHUhiJ7qJoWlppRPvtWSMc+l6i36aw6O3eig23ixfZoTodTWX0p/wikX1KwFzBf2
006oL3aD2WmpCDks/+BZ2VjYxRc/Ocmu59KFqyTPQtFyojhbHxXFGOFZEQ2LZIJ6
ZxB0jo49L3g8mQ+vL15wfy3uSj4B77Asj4TOHh/oMiRPK5/fAk+JHvD7qX7CzwJ8
HRvLKkn6KfZsLb+tKyE0JFXjqUybJpS1znh9W/BpIuiEFekoOlc6TumhPWavt88F
eHAKWqfCbYfx5+Un0OBV2cz8Q8OGVu/ePl0Kxsf3aP2qZKq2ZKkO5qaKB1Zt35FQ
hdqmXTQOtRm4Mw6CVOv/UHpbSDMfr1WbqmO4IPkfZ5AUhBfuzw8IGBFBT7cEu95c
+3pIUtt00ba5pSLJZPSqtSkpuQdjYOsOxqWvcZhtubR67p4A/QMz5PQ3GbRHejVf
flwwg5cWT78jxnvtpXIU8mHJTnxOeCDZpySrdH/ZKrjJ7gB4CyaWaPcVyhVB/a0P
lWWyf/Rm7P4SfL/FvxEKNKAuQX0W6OHvs8EgkIG6MNVWC/s/mIHU5JcctIo4Uo6y
viq95Oo6YijlWz/9J40hlNsfP05wBzqAzz+TceuaqjVfdSlBvQddqdok4+i23a1U
dFAFBsA5RYsmuRLLSHZpCpiJZFva++qYwS70Fp+SpUm0ntseVr15n6c+eKTDYO/z
1lnM2Piy77w3UOmj7F9NJrH34ShuoSnITu7q0Bd/4iJZ64hcJhEqS9sXlo8HKoW2
GJV8ZYB2d6kRhMPd3/gVarFn0PbE8I7dUQkHm9UwpTg/B6rdWgjIlLENpiZRJo1Q
5srOEy6d0h/jgu5T++QCNMBwKun95o6Ha5Zs/cwJmydHWdlS6mSJryiUzEqULISU
VV6n+UrDI3jv+NzPMDsCP/xYi5JQrbdwq3gST1LILz345CvoB6QB/U8X/bz1eXm8
r1PPsggEYdyZETpoNmoUfyvwmOSus/azJ05ep65xZ6RWTfjeCtfhcwvnmM2qwRv/
UeiHckDe537VquUfGhUpGToErMk95Mwnj/1qCR5WuHivVDg3xjYsLBYqlzfQqQmr
ESppMC+haYwx/GjBHA0JrKtfxkU1Xo/lrh5Gf/OYwgHXXwB+a7ERHT7+a3Syek4N
ddZ/3kaMFAjIErS0x4G+bkoS0bWPEiE6SvzIARePbMsOa/OeILjMjEydfdw0Z4r2
jKdYIc5oypmUbcCiuX9WNvNIPMq69x2CIOEGBg0HENQ8pDwd56MMr1hdgoXYfGlz
IJOsAS49Vz43bIapWigxRSDCTVpFyCy3sTuXdgWp3yCMbYG646BF9//Idm+V5O1d
jnjXTjkwG0LPM1+iYyb8Ty57TUyRSrokgay8in+yaMkG8SO23AvnoZ88+2IdQeds
TjuSXVVjJbuusDIpjZLqDXxkpLyWPDKfEMF0AYBXPDwK6Mu4TFwsiA8yl+qTpG2G
OvPahqquNBm/NlqeoJUk/g==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
a/gPHnDWHZ6+CY6ORzQGmrYEZZWaz0rYzBUB5oIHXnbAGH/KYmUAGe/Qh5GGn7R/
bLk0ylzTfBSpDV61RUwaIpqnwW2sPmGEu9PPfpURnTaTrUlTerzhuXn4BEDQYXe3
eQ9XB2lx9oIk3wGfDSWKTVG//eY/kimo1uL+3Q59BowUk8kUd5XWjymWsxzDhvZ2
zrh3Yaa7LuyCfd5TCgLX5TkX2ojR/YphsG4owHwmB+SU4rrpw91WJofMDeMl/kQK
blkFWQiZKtbgS2IjSMQuOLs75V4LK0o2DdrYTvoVa6Kk7LJ0rzcnnKSiHwMpd3nh
9HrZWVi0lw5Pt01qacOYpA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11952 )
`pragma protect data_block
taNAQu3bu37KjQR+H7zrWI+8+PXtGpHLUjZBmhGJE+P9CAZpAbwqM0sMhEEdjGmc
TA5XlNAiByiR0MTXZpJUVDKN982fQ/ipRKok6AIZuDNNrvQ1zhxfqIACuFHnPWu8
5JAN7FaenjilTKatT2OxWvM5viddeZ8zTfZfVOQX9D/8Zx7a1bvd2jUpDNEf661m
IQxLpzKWebpOLBnX2QRquejf3KX7DqqrbBI/ibi6yEVjQAmIcUnubQk9KGZXxlAN
WOhw88dRgTaaiYrYSu9Q+dbnNPjsTPQRTTw4gXL1lxDVUF5qlkj6ArJ06UrWRVDe
yUiudoLLLStkbx0aaBdRa2y5mhvGMPppxrA92Rq242akQ6BhpEEYYaZm1F/TiYT2
Wo3imAnrgKjZN9NG5t/Ja82s1Os8r0lc2XdixpPb5/qLI0dfH4mBEjOksx1Xemop
0qUOMWZcwONoeU34WUnnjIUAlPeTZ3YBYoib2PhKOBNHdOhOsqkMfjAKb4JPj4KZ
6ElJJdRRZbgH0+dS4xYSTExv2xZMMYwnu12pN9zDCTI9F02+Nml/Svp2bKIfRr8L
5tewcbLwY063IIA6zZzk28gfsFCP+8kGnOn/jkrBlvGgUhHrSnIweSuZWqqx6aVa
jyBHJV4kRXQfxSRTnJTCP2/QiKyJ9hpQ4/S2qEYdNnvCIv9T6FAdLLubkf7jG15h
AWdh6rnT5RpXh1/X44TItO4GY/hD1/wkD/xEfI9DzP67eSmVQJvemQsblPAO8PvW
0mAb8nvO+1wtRLhi+WwOH0n8V3bG5wMbC3jR+yZqud03XxsdFPGsCS0ROkvoxIx0
FrsPauTjhmlwrnVLMw5Heddrr2W6baZ3GMOqdpmQlRQE67ab/cfbcFcaOjc9ysWd
mG9KyQozIf5l5EhUinBI4cuQXZnGbrmLMF1j2z0qjlM25sVLk3Olh+UzUHC9w36r
Ql1bahg44SzeGSMqH9gQ8SQglJ71LRfeoxLigQM/4oLwgE9DSQvw3UJPN1KK2OE4
0wzbWBrWanKsv7WgrtTqRYavp73AkGB4QFreaNG3IRXqtQEUCBnCAqHSuLPqeVOR
6SuqIlmX+SwENxhwux0BePlHPXKIqNAZd5/2IljA/aPYURCJgRlJkM5ng6JpG97o
4HjJ1/aYIhHX1bKEkmUjH5gyxbm1Tn/GfkAWc2ZkZZ58hVYHzxaWwiM84vcbQPGT
BSMC7Xqn8pB2o0Q1VPFNogotyAgHoWFD7eLN6owlb5ls/H1pxVYWXslLd07OXCW3
FOPrB56+PEDlzcqOJFYiFiLnxMDNN7Im5BYGpn8OGfZiIyvGbMyyEgax6u7VtOHk
FNbSIc7O9Vz9tjjfZGkrjAffUPj06txCQzkngfW4zqsq3XCbvybaNKEeuDoiRP+5
KoWsES9xTGCxurCELr6k31X1AvXSsCnQNBODx/iovNUlMn1vof6cxsDM8tG5N3R1
hIPyEMEg2rgroLF/wnl/5NTuT8RLsRB5z3CLEH7xhhLtAmIJhRBNXtKQARmm8oaj
mMcp/yOMnrt73w9ND+2e2BiNvmUKqpdWXgVyaEDez9CDPJLwfBZJUM/oScSdMtK5
C1u6Kpt8laMgbD7d0R1LSTLC990wtnHuMviKr9sW9/4kOdy67WVZYFp9AmtEoDrZ
pwr/xXvBhL1eJqU179nyVDUL8qvrSxt01rycyu4SFTgzIjhrYrZZaN00JGePAmXe
azuec2fc3KQPJbEytz20w5USCOqh4ULAKEmba5F0sBsioQbePloZrQ6ufAMRvjuh
iXTM3VS2xuz2ruDy01L8E8o3f/vMj83Z8rQVeF1iprDt1nW1u2zfx1zqckN39FVf
cN2Abx+e9kp6ntNmp2xcr8vI9DhGqYnwL7RAvIPkf319zUnI3Z9YbWBSzvl1/BBf
3/bvFSaAyJcnrr+QsphUd682s/0VpBgr4iSaHm+UBK4X3I5iL59qkLWzzltRkWLh
1QSkGXXKrSgPmlp7FHems3y7j4BN2pWqKm2egSS8hVX56OTl1draBPb0YBao0dOi
az/XB5qZ0tqlhyTKsjqnd63ipGVRwYzGdNTl1jfGqWrTBqLsoAGWcutsCqam+hrP
f4SdSuuzrE8wKXyyHu/pc8Oc45isHuoyLggRsjPAq/M/paVsXwMctcSVBIgAxtqG
YU/8t9Vp+7qH9WMFJBLrmKlIt/XAss/U3cSgYtsYnQT8fUMoXSvff/E0aU4Wfyio
VcPSZ1pQdqOF6ffXZhSqZKAqrHmWT1NdTN0+8z3FVzpWL54LO4wrgFeqN5Lvb4f3
D0Ih4NwDWyCS1WLUq20Bs9z0ah+L9w6igm2Qz8jLv8SPIc6ylUVhTGs/fybc9wI/
C6/ToIHqCRPSo8xkeL8s8s0W5RttdSkintrfeO8tXWeJMfGR4KsoG47WXC99TejK
tZYRUnbPXbk43S1YT9uHzzTyooqHJ2Rxyn7odbdSGjl77YY0CCc1xXGvxz2Jn4Ou
/mX6zEY8oDJJSborpaE6Cc/itrGzhcFKw7av42rrBr4W388M5iBO+QStInTv8c/F
Bgt4EFSSrxyCDzWD6KPb/nxuK+QWnHE8bH6mO9xJoMxeAI+NsIDsBADZM5D7MN+U
jwfl0jmxmRjnSXWRHSTe+Rjx5eE92y3bUcbv4yf33Qa8XGkz4TIcLPNSBQhU35nb
SY/TPp9xnx0gM+7V7A8fkpp66miyDG7TQVRMNvNlWrKjD/SshEXm2OqFouKZDRRi
eYkwIl/Z4bnSbDCVOnhlaWe8GPxPsbtZmffC3GS7LJ+KVLIfiOcjBgSiwGyjX3Wu
Yqqnsq87XCSn4El/HAjBU5273+MuJiRTP3i4h5LNMsHqxjx+01cARPz/XeiQS0ne
y6YC2zD4weHH2H491MN49u4ch6rC6/snoDYsy7SOzSUZhegCLbewioaDVowA/PKX
46E52tUC2R7wg4WFDcfZGd68qCpKJwvdDtUMW9VZ6j7dWX8hpeYTvMWl7o++cwbq
AD+9s6H0X3N0iaITPGYjfUS6wd7/x5PFGaQRdaF+D23G2H3GtIhaZ5faRzyNMQCm
rQtSu/73MEL9UBXltv+LH5JM5ZhW4Gq7uSF8f+iY5qPQkbDjG8wHfNEnX1Zl279L
nGQ9Iz/OyjtAGIN7usNaEkvQ/E0IgEzLf+h/x3RzAPZok1Y+32femFt0Cls494bP
MKBrd+0JMRxi87WCMkSQO8BiWOLwp18kEOKxq7PCD3a1cUNQZTyrerRUIYdkjKvY
C6jWja2yvEP2NkycYTILWVkA1QDd/Atp3BhNV0xDGx/ZhmABuuuSgraYeRZlyMO8
1UkGKondra8nSMMrCZAu1cxNXnHEXFvXIcNn054TDqhHzmzdAjbZusJAZWwszEO1
sosvfUGjX1mWmIgb2L1YVz5KYvAqmtH1SiMvPd12Lw2eKGvACS87h1P2k+O36mQP
m61xhsQ2A2lu0kK+kJRSbAFdSo4htSEOTzyKbIWSda7MJsVUp4kGR9SAFhgVsGlC
zehCfWaz9YxKbwktsQiLDTnOpLv8mCelnRFnRNDl8A4LL+NW3S8ukxe9WR43eBph
fBIvCn2SS4MIFzsXoFuyfFVO9tp3agj4O5dcDf/8nBpqD5kElSy/2gJlwhWp1nzD
612jVZtWmq580qyyO0t9aR+Gy4f6szv07JuQRIVqhD10YebV5SnoiJUNAeaOOtov
aPk58tuvhYk6cDfFvGs5hH4zqAIOT2NwFZuDVMkdX5CJUVBtjsjcQ933QC0uvNXT
qQUONLGUOgq26KQtOqPjlugLH4+7hToDXyXs0Y1YEqv/ldDYUQIdq6YrC8RU9WVn
q79CzQaC0oKCol+5Uo5dZQp7Ynj4N/Yn3m1Pba7Nis/1X5YOfONORE1JCE+6RcDl
FOb/Hudn51Vp+bplQ56o2ouOQ+zkjbM4Ttp2opFAMZWj0+y0aYT5AhwruU2SIdDi
LTfGSqgg+Q1uZTeFVQKr8N5WBIGSb+9vuyND9IWfSVrsFQ4vFb+gl1MJJrqXTUgF
sQbohGXUYmzHrTbhPT3GeZFjKBdegswAHe+7gCE9H2rxPEtxf37dNJcCMxVEiOsR
TJKcmYyv3gdtErISMX2B8fYqydWtnCBNZx3GQrrEVv7moUZnmqHxkX3mfZRsgCa+
oCHJerEt5LNz4sQtmbRIUrY7Tfy91BLyzW5sayQ3fErbRuYr0IgsHnK20+/dXeMr
cllq8pAnx2nSh96L0VY3wf7ZK34znvZVOxf5K6pt7CeRrmkzHmHJUi/LZQRoq9sT
LIAeHmrtBmpW630jBhOeC/SeF4B/nZt5HgstD0Kb0C+s0jM/8kRl2M8kwr5Bswfi
kNZ/HZPd3z/o6VdFlHOm9jXzMocNXGkAHdN+0Gf1uG50PfQLXIi25d1+HHWNaE1z
Ln8TTAYTANpaI6oPwCR9hAC2tEgYj5dHRA7imjKAjjCDlYSUcguI0ZtLohjSqe1G
G7IHVefgUFnxl5lZIrXPwweffBA72/Tn7YCVW+cezkOHmefkHLXxzgiMB2MI9M5J
DFAM/qgIGOGZVFBbvfPa4Mf0Fs7p4UKxSFLo2ZwSZw10laZDOGtbpmtdn0mAgo2J
iEtwXECwdI4OWU2RZeszhLVeGREckXU82+HeLVbFELjbtd5jBzIgqvpPp2p1WX6H
lIericQG1YvjMBxxEBiEqrVYUqw4cMBKV4y5OT9NH4TttyExH9vmkWFTooeRTJf2
q+lzIL6GMRYpoKJhJTbclowoBUFmcheoc1pXs03GQYoJybymvRQWzDLjUD5T1yv2
fYalfrNHUvyxCHouKdqDe6R0XNoPB1k5leGgm9HI8oVRc5oghEBFGVHmkpC0XVmM
mlxaU01Fq816Clg9JAdMKEbvqLPdukeV2r4yDMk3frxJO8DOJv0fGHi5rI6Btv9a
4HcDpodp5eC7pOjjfP6993BJUeujn25bKoJLWWsUYQpSS4/IJZK/mROq+ppT2clS
RtWoe9qWGU7GrF0F7xL8hGRDZGQ0P9xH3IH5dPCworf5q+CqifmD9Nii5lqd1SVd
jpbFwrruPu+Mwf7/H3KxVsYROAJtWMXWI+RUHK0IwU04tMt23NJEVXM1MSRc926w
6G2rwTJcS6tlTDRtcgng1Q/tRr003ktZnurYZknrGVU75wW9wM2johnyvqedRxqH
h1OrtDlSv1R/zPcZRmlmXTfYDojTElh3nGjhiIwD7hiCOOpLA1BsxLB2lJmZvLj+
O6/gqMZ8TxPwWbQPdYUlTsYzd41z8xrbks+Fsv0suea2IZZy/Bu/a7CezvqotUtx
n4W/i5nkWMrYYwM38X1fiUDTFMEipFvrgtASqiFGqLC+cNQPJSB/zk3YvX0013o1
l/XS7TKYWp3Mvme8Bd6498qnUHE9nIwDQ1nzfOLp/LCgJfZ4IamUfGsPg+RtJ7vi
dAfQiWsf3MMlSw7v2cZIyzjZs8Cg3pt8Z1kwLYmTjoS5p90bSb1nBOxbf2/yqFPv
ri+ykglrBlShq7Y33VE+cnkbx/8ZJO6N6GVmlTHOywsGCC7GYFcpy6SX6BVLMQ6G
a0X4I78WhBT6PjuSJrbhfX4Z8Qdxt1OxdRmbzYtHQxN9GKrBD4P31oq/oxS3qBKO
JoTTXfGVpHp+5WQ+PvcejMdsJyPw8b8Z8t9CFabKjPcfw1BUddQ7IfQDcLS0bVKz
gI2z+x5IOWUBoOPk7oYtITbWidzu17EaTbD0X3syGAMWlU+AMSwV70wpo11mZzMV
OI4IGPgtzUaIXFPOzZeNLnG1ZdUMj1nkndRQ3Sdp9NHsJm1p4FPZU1eLUG4SgUNn
z7GbSYEL2zRooXPuSoZq4GE6GeG/5D5tGWOsCrU7FGkMt8knSAGa+F6h22E6rlu2
cauyWertF4vxnBTM0nuak0U7sCg3bJImSf9/lyUpcBbbQf9WGU25HdmMhRIsqsFi
o0GFucRy84Fhje+a3pni1w8b8TAPT9CbgIIgcJhVM3AJ0Bjve+e8WfhXFA+nuoHv
oSYk7W2C11Iog0lo09A67LRe1XhF9jDjLHodvR/CSHS9lDknJ9+vFScRUMdFUcXG
Uvlf+GljKHWKXPr3OHBRZbTpUK6KRx5v7GUpUeTmzMQJeAchLQy3HfchcULsjdY1
CcfZiYdtE13chPZPaD3fEoYtxvYQBGA0rT73cR/gi4p64vmBsLLKvOeq1xvxh85W
QKBtPg7hGkV8SGSOWB1tFqxRjXxDfmbfBGMUzjWAzSJ8p5UgNwMunqgwwe7ayDVl
lzP0P37B6X4AN1POIuSz1+xPMAPWxq2q9+E+THtsfMmzBPWqECTYLNhBcOmmuKZV
PsEBHKQF8KVOLgH8NAymK/ZduloXr9fb4mWEfC6oVnU4UUif24a6eXNgzrq8k8jI
89wSsTkooPUZR0qimNzbOYqiqX/3CKvkOfV89R2EqcNLcyCRXmYEPPSiDMunaJxH
FrlgwW7Nj0ozuVU9kcO3VINKBtH+lJ5Asu9QVzKk37ulhUG54vdhVDN3lPw00++A
4diHWX5q8KskeWZOhef3CVsHVNepBzfvBTkZz/mgjSSwfOHAXzYG3AivtVYRdoxT
4YyfvFH/xQWjbPqyn+GmDoQJOV5HBWwUT39Rp21gFMS6YoQT921ZX+NrffExnR8d
C7ANBc4Nn7L4k+K/OUSEBEAmy/lAnu6aXsPZmfBPvIPYnMEstc5+SPCbjY14kNtp
yBiM/oMtDT5FNGRVpmeWLsKzGN/F5Il4p48PfjZfqh0EG5KqTegJ6zK84EkMxUY8
x+muA0EzTQ7cEM3ZhkgUdCUSw+F4IaFT2PIlV9gPSRSIAHcbNY9b5bk+9gW+hMau
l5bCHcO5AhbOl9hcSSo1b3VlHY34Ir30IuXBy9tpwsNo9rI02gPvKDF1NY2ENxfF
zFvHea88lRMHQXO33OhsWZoAnvmOl5/ttoTLsYCtg2Ok3f6MXR5elHW1QCaVmpRA
2LVvDFAS41NkwxSo0X4eQ2NbpjBbnTpGd3wcQQJ7gL9Ybxwl6FwkT0J7vL1OJYNJ
eSVoZcegXlRbfaXXYtt9dgJTJcYbtJe5jMCN7+wNGJzuRSAsnOi+RH6fPTTUhzlX
eudLXkOmYQ/AiInPXQLDgc2qRGTX2yBAKzOm/RYsRfr495j4jCsYF7bJT6TAMi0I
/qClkF7CXAgY4cwqPomT001lJHFrRqkLBB/DlTO5kMCjTiPk5mh5z18SCwvOHROz
kdiO3J1xhGS2Ke1VYCwqp+iJ9IMddpwtg2Qw3pZRdnaBg0X20N/E7liuiHt9bxbQ
yGd+z9KM/BkL4gOmPlhvfyOBfySVERnpxHxCTeE1OAKEwEfZDvQacKx/sss22rVi
NbfCBKlN5pspoWxMRt9iA1JndPnUQI5P+mEx7wv3NHWFIew5h74shItiX+3UvffO
GSPPfRzDC0U0bSQ8QCSaQTWOwmIimZ5dj2fzmmft+98ok1rhhfMDV+nXqU9eOLaT
IQtodW1kieDJYb8UBzRt8wQxRfCifStnXwYpoHBHJrLTgknSf+ca1qTvSbUVSvxK
zqzdHx/W+IcM9yQdgo/jgtkShPkrag1jw/KSgHVFxa0aTW8lOjb8swTO7f119RNX
ePWceZih8XnFxjNo/efbHFd6Q7vsoYg3VBUJfaLgICtwslTdiZxSYQcTjawVHXsV
ylXk02BDs6MRZwpu7di7OBHO5cFUMGQfF9tMsY+qLk7FLSnwL0hCqm13ihzISHyE
tK/eiVcv/YjNctbSUew5Mu6JjOjyxTbPHCM3Rd38E/wsNqIVMYQNeNUo8Kx5QQlD
9YJucNVIs3IJwLcZZFTIiOv/bp1C9JRRzBVLHdEp1BGnB31aQmoAVj5o9REv2nNy
GX1HcdnF4vUsE4gcmtInd+5At51tD5hYZighhk1tx9XHCh7DZUBTxc4teCgMuAHN
TXspPARR+WOMA6oHdy6Pn+e1b8OIM5bizA2Mr1sNA1Eol/T1knCVQLuvTFUPRkhC
pPyUy6AXIzrgux6ZNIPY34/IN5wiMyCIIAoEO9HJo6zrcC34w3IFLuwOweUzfELn
8LgBHSnXn+79qsH0zkHh64WB22mf+shJ0KrIVD4CNEixx71Mdy54xn8XD0llTQxE
1koss+rzC9/5VtJKNECSryzpoBCO8H9ogTHNUP27ZT92weWki48dNjVFZHrnHk/Y
nJW/nJEWYEcU5+d/kOHn1x0+T+qh9na9S8MzmlXrYQMjSw7Wdbhzm+wFJPb5ym7G
d3sLEZ9RsJ1djnvwjYwN+XT9bEHDoITAx4/Q1bbyUHaQMv0SI8GXIBteMAgVdyLW
NqX91vQtfxnuaMWHxb9CcOY0HfEBzx2Ta0iO0yjC6ObYFqIDn2+ZecwbButaeOnb
fczxSw7jG/iT0saFUg1iw8Q12P3C/Uwm2PkGvc/3LDOeJf8PFGfKpf2Vp/Cg3pTW
O+mR9Q5Xa5qupyulL3GRGQYVyFRrX47gritfHawHJqYivD8WWZZvzJJrqtlV6FrF
P0iNCHmciSOXiW0xMs08eIHaNCbmWKMvFmFVzS3XOB343l0U67JUdVdB0Oz1foY9
OUSDago8lQuRFI8ypgkf8VbZ4wc9f4f/7t/EHLE8tQkmhqlaxInjhWatF7bKom+N
OIaz21rqVZCesfjYzmjLaeN03bjEJWJDfWX8q4xMHEEXzzYD8RxvzdgniwZZYKjR
OGglgOo83k4QAjh10M3/2DyqARbMy4soWN09ZSZS0TO3/fILV91MiiK5v5bdA073
KhUd1nin6JTTBuivpN1Rv7236eUMLBNjFRaPJEFBxDzo8P5Dov3eSlIDFDG4Ezxs
wY6GnC0r3XiU4+78GFOfvfhTihMkCtb1OBK8SuXRXMpgZvZLj7/TYrcVAoTqFAKZ
8tj2PYaP9yjSLLccUU+p+iLH6uT/XspXMeD/AtRfqSpXOWxs+QL6NCGKjENEj1HC
jDmFqxRnxJ5729+NSyY/s8wdPQBOBZRYz316xbgLijBNpPz0Vk6+rT6S8PDNLQiI
RqsS6kLgxpO7bY/LYxNFdwdca+J0gVZhOuJ7+F6t5zgpVxZAH3PYwAMHw5ClAk4w
pp8+QYkklRC0O7/xXgQygJLg0/EHJpyRNpmVz7x7RbfSogoR5aWrZTT30ke2Hm2P
R5OlqduF3rU9uROoxsm7uhoiPP4PVAvnm8+ku/4RGp1w9YwiLUnSkukx6XYWa4Bl
0pcihLXSe8rbeez/EdCRwQDQ97ZgILvGzHcXvXP4P6GHgEFjvihr/2P598/Qw/8U
rlzCBwuk7pCHEqabACF+dx6gUM0qKgShonwYbtbRFWP9kJFHF4v4W0NJmnUowSKA
1nJ/ld0uBb1SEBYPmoUjW9ppS4BEFh0PZajf4yuxnk3A7Ensibcf2tOV6L/xWScR
Fu8Ll9eIQXtSxuZlwLEa5WHAJJ2xjBTiOc2vG+WJ7v2q5UhFXKc/o0oKrWPu5PI5
lhi9FNMgohpW8JwZRpArpUJsg6EXxXzgBrMUq3rIgyJkiN5X4+i6jLiFbpYXwJk1
cAs/BYyYtmN0itam75Wrisx8Bs20hvjzndBBFNc0ULun8r+ifzL15i7FbBr3Vh8T
wGc8NqL7x4TltBcA2POtXBosTdcaHqKUR0ySjNCc+fcd9HS5DIt6RDuFUsuNqT32
v+DlZxsI4Pc9YkZYnOcohB/DOq0iHzUg1hvp6RB3x6lMLPdFFrs7V8rusIafuIlM
ipitXuTZy4o6Oc1WzIiW47pDCBD9Ei0vLPyDdOjNv+0G44mhmWUpyf3x/LEdCjDR
ZvkNXE900TCYrdapzlNnjYXgy0E/I9cJX6CM42aRDDdhGJhAezg0esvaWMra3KWU
KV2xA2uwA1QfHmHbfKQEotLsWdmfCtAd1XOxIEwCcA/Ag7ptyXG2tTCxyFAkkXqI
pMIuhC6SpkfgxoKKF/mYLXuOeaHYGtoFJQsImjYJgsPeCQVmsl0VNp4MQgMU5+/A
zL7Xp0huLltA86bGl2I9u2SiNAu1V5Vt25VOyW3xtldflPHzwnS5S7uhm2/+o3ZF
/E7JammkKmTgjBCznPk7uup73/QO7VlnLYhNZcwAhD3PC1kmnnTZOtbFjGpG+Eh5
63/wucCpA85AWNU5qNYCUeWRr/3LVAbMQrrC1FiehsKfE3dtCe8+6jReJfENXLVx
zKoTIKjAXSGg8SlIWkez45Lyqh58JSVSYYAS7zKX5nowDbtbU5j62jg5DhkR2CTh
5xXKAetB9R/nPL8xOQggCQHFci478UGwAAPMnukK8D9lN4zwQoHCcOfEMtmdtswB
fbQh9kiUmau45zEWoN9tP6VcyMs9UnQi2PWX3O017tH33nfy7SZ9vwfvBXt+G96I
N5VaP8OvpjBAPZrD/fgVi/2dz9XlvEMQ3Cc75uhwpEwZFZljlxWiAo85jojFWmhu
49x/DRTwjfG2oalT2pHe7NmN3/P6/uKoN7c9vmM1pTiBKEGSwmyO/Th/iSHkYwsp
lvFzsumzMO1eMbCr5WknKnnxgAYi4otFMLJiM9i+0wxk6apYiak8RTJveSCatqx1
quDh8a5V9qOTj/cZP8Ymn1xmS91De/tkAlQcyZa01fnmo9muOFd5aWhNWflXl+Kg
OW5XvTcGsuk2Aiv/MS62s/TfrBBCBlRmOv8JMMn+4k2wEz9dCz0VSvVXyJkANxt/
rs5zPVB3RV3Z8pTTP2UbFqZLezlKEXks86r0924GQgwg7lAkFapz0L/24A9+ZrBE
I4DJGZX0pAI6v17FVRkhUXNA4omkD1WcpQF/5kQ5bK8BbTB+BZJ+MQzZVdvUqAE7
A/ISvSGS0LILoIj+D/ZtYE6CFaf96uiFdmUifjS/lPJRdhUPGuf/YET48m74Ns5N
wEfvJCLzNG6ZEzko8KMt9ERW0CjRGaICUwPSXQoJL9mRfWmoaBIQ9BmMWfyI6c+G
hfQnLY4dDaSTHfKzxsbwFxUDeax+1SQZIv+cY0/ndUxpCRYQ/CYSAcEuTi/VB/a2
xXLxQ32uXoL4EMgzWEbluqHY3CpRPhUkmc48TNsyKOPKEyQIXR2nth2g1mZsbStE
193lLWp2ha/lmiMeGEmHf0juEnuqmYhmN41nwMeEimbGso8RGD65KF+DsFYDPw6t
Y37oWYLLXLFXyfjsGtY+c/ilHdh+fnJn9Sslna9cgLnwEsn5c86RpLtn3sd30ccU
8bjhCA/s0xTiSTTGt+0AHGOqP/67kjTgY2wpJP62voUwAgFqa1JopDQkoKpODB0q
daG/YdoHdcAXkMmyIH4u8Ha6A7nBJPKsp7fA1SCIt6Ksk+wqHrGOf51x/8XqeNYq
QzdaMmSWEBWQegSJLgYP94c3tmqYauQZQdaaCQn6PmW6YjvUY+6ROVZbbW57tZhO
l3YYfQlSwkttMX4tanGjF0vqYDsNh0pOx96oMDM64dfeSE2nAFCCT1PRFKraAEZM
NUh0U/UVuCBwxkVXokKKEcNqlKuG96X+Y5ePy7/4IsNFm33Yu+pwqvKh+Hbsxm23
NUFFeZY/nEZsmReR8NRfhEBr08I0qqqh4wJKmdlfcvf/qChRAUcDXfPcPbC1EkHk
HpRDIA6fAwhGIqiT35TWHIwV6lw2s5RiQh/TI5aFd1zOEOMHEJR99Lf4byjdfOXW
SGg4162OXAqFjoFN9K3lBerVYx529eyJUZ1mVcYXFtlDYedditIt0DD74+lCpPfV
7/WZ61TScb9E8zeiL+wKkTqbYIEbUb7MnJF58zkXFiUzF185KCcD9v1AA3s+KSgD
LdwJyi0oicK/VNbXU4X9Cxc/ehFhSwioZNWBmbyPZVptKhxrIV47TBR2ycRf23Ca
DB48bu27HlyvuxuxVNaJzv+jFNjSwE5JOzq0BRBqwY34861imfDa9SSVU1+jSR68
AL4nZvskVTxkJnFFLIOb3lc1ZsLZPgNDiJCeYutstR5JFPYmgikcdZ84dWS6GJxk
21rFmkAPQ2pCdi2mSozq5H+R2NYFTeVv6p+Gk/vQtooqF4gMhgXHE2UEKJHt6fgV
v5O64qKZJt6UuitdQbs9r3IsTEx29oOWc678+I1LIi3d3HcCb/IfOXtzNdZjV59j
PLi+9HWx78MFz5uJEddoXH6tCy9PEU7SEDi74iodDrLAeeTtMgKS2j4jut7Plrlu
t4tDWlZDvGYZo+LrP0NfpKVgWJavbb4VVCIkv/P4dFu7iGeVW+QYd+n2DX+McdWa
eCZZ/Zg1CHaFNT4aBdBic6wnAdm8vAX4nhCI4JCpMNaYSKqWVTyPr1oyuWMLJHRi
o34hcqkP0VKbHfWMnAfpyJm1cb4DqwrVly7Yj3825am5+AlnCGFAY/07yz7Jd9NR
X4IGhaM+yU5jDBlMaZdLl0SaQIGxK9qzxX/7vYZbiDsuFhs2fEd4BllhYj7QwjEO
MIoZI6tLo9o4RUydPuCYMR6lD5d2F1tM9YMZ/LBZIiE0ONIWyIkfNZ4gj0vUp2El
Q+t/6/SR8buHggQu6YRDUng8RsIwfZyVXfvmSRmPS2Sx/N4ojvfn33cDjAZuhy3L
TaFUW/waUlZ1wiDtGXJ+9JLV09miSMl5ol+vbh1b5QZdj34FIzro3iaACCDWdJY/
zFnW8nHEu/A3l+Vg0SegpR6PNrEgDqohAbAz0ZUfTZJONEIkwu6NIgWRH6ViucxZ
ARMY3GOMu2V7Kt2BzvGv4oO+/2XZxhY4QWaZFyLAdDz/DKy+kQHOXzHjOhGKbkaa
CXVyOiuvq2FRnOaMsE5dNChNNZZ/4PETmbvir+p3EeTTpy+oDFZQ/YwUDKUegY8/
wSe6cibibuCyz3Bjn8X/C3QcJ4USeKaHeW8hTxbS7jad2T/Ss/x9VOB8FwxyWdX5
246kVOIHkm1Tp4+vWTDW9rDvzMMXcCuTmyTszT4Y5Ft/OOLRUjv6dUf/+foNgaQG
K8n6Mpa8PKVMin66Mhs/oLS7NdWPPyKKQllfab0ZcJ+09XTRRRGqXQL8+t30oZNJ
fmqn80rm1jLFHdOvYJ+AuZ47raSgU/k5NO0GoewfSYxw/hZwp4KO+ij/2JfjQAsR
c+Yf0y99ic8rT05JnOpJaLi2s7pS+At5wgD0+ZEoK8kyPNsqrDPBzv1KoZeLskeO
GB5T8MpWx573TdydVjzgo+Ua3P8RKGgCG5VtMykn2+bc1x+EmmOVj1OpAq4yyJNs
4r9Reyp/ehRhj7wylgiP3Gw1tudqxXFsU5us1OstZl+zETKj8OAKEuGzrdovrXe8
i9sumeP8vIE+Z0gQiYYgNTn6Wjd1EllOj9F38/hrFSQI5L8arm5a0UXNd6YBhRn8
9lDJWx97R2icEATtRzL2TJlNSzNANT08dDE+6zprkCkRl5BdFHn8tDKqwdfU92cT
Xpwlgkr+WEL0gx61hZI9EHP3UHv15ESEDndopH126PhRTRhZYk6D83ztTyaAdo3Y
P3dXoXEHlnuNjXMhvGnzHjhhn3n7o7O0mJcq/ZeFWYLsTKYrDS7K6hUujbkMcchG
ANaa2WoKw9b4HO4yH0pcIxm8xNlBpcbKooCDx5Kf8Od9U7FoEfFKCkDq715QWkI+
G75OAHxIUjV/MFGnV5RjSvlcLkxyIDqaaUHlvHTVbtUiThbglyzTLfaKOrqgXiYV
1LoajgKUSIvJVRTiOc5j1Hjpcj2+V6do6NxJDnh/9QD5h+8O+kxTdLmeNZk0p4Ni
aRmxevbD8pNmo8BkhXKFfAIWApnRL5iJIW85hHJQFfDJZ8BV5HQgEvBQSNvhqOQw
Dbj+VgH43NqJyx3HRScRqqtlihWtswhm5VAtMhuwLoNI22dUASl26lk7RZtCo3kp
fQ62EiiQH2IDEWx3Jic5qKJAHglQc+zqNpAqEFHq8jZsxBwG9As0NK6GIioGDAcK
OxPi4QL+KQTC0ZV3AIeAPSoP2U13mFEI4ew2Nb090ZMmpsgg0r43jSMsgDLp29nS
PwKzHhH1u6napFDddEiwEJdPwVPaLAmJEPsU1pAN/iycgiMG7bGLZeUgKobKlsi8
edHqJIjWnL4uBUUErdJ/VXgktMMMzAhoDAD47aMtvbWA8ydDs4oyC0imImQfeKxV
BVojFpu31m8t8RgUreoFYKtz6M2TzIz4Ogw0eeK1dQ4E/haWKLnT3HYnp+4QcKYj
lP+vKVVP9V3Z9J13+6+lZk26dDTDLv8Et7j7cXQiZpw6Tq9qylPDLe8SD9GAaWpy
eeBOSAiTC94DBEPXmQ6GSPqhnMNXsD5lQKajIIzGY/u9x1QjIZHBeyKcpkJqw/IP
7RwNGBEr52he45xu+v9idbet8c+1ENe4fuo0YkN3gSKnIxlmuHr/gw68WJ+qSql1
4pEn0Cz6yEhUb7f5tLXlnaiv4BbtLi6lLhSAMdUAySrK4USReSQKEdjs5pWEAX86
OqK5X9k+wORH+FFzvXRgUSFIUKYaLNo9sMy1YaCTYuL52D9LKskxwcDCf71VqqDd
7LdAuHyXZRHYK4cTpGdYVreGYv92uafMMqpJxdB121TLr92i3yHi+GuXmuOhmao/
A3Y8pMsfI+13BrZu95SthSxkjoEKtJNgBYNDqQe6ZtfJpjdxCLgufP9kaleeAewu
oAgJiBMC5AhDMcSbG3LxT1imgsKCyZhbzhg5bqQEdi54vPQW8EXF0eY5qZZuKDsU
XkkA2xsqavakdrG0u0e0TLH7NsyN+SqlFT2ukVYo8LPVQjnFii3Jtd/AMzupB9mp
wjbTwSwhXreFuFnbpoN7HzVCOWZn/hgcew6Ei+6lxKgayBX5+Lu62yxG4iDCfZsR
2YmqR0pXRMyppge4zN6bqiYn/GmZTVB6fp2qdRIOtIk6KlJ/LJ+eirMtquvusOOF
sNCrpDWXjbTCd9BHo6gXeD/mL63Pz0DrQv9qrtHTqqkM4bTc/wo4H1ekycbAWBrc
fu68xuImOp+MNXhEoEut4Yqdzul3qo8eeOR+Get0MGXw0Gyb1/EEG48sGDZ6PGAA
YDYkdu/3DWzeMh2VTES7kcB9MyKtLsz2Y+mugPeYMQ11BMZWc8x2M3oIu/Bb/E1O
nY8BlXJ+WWuGJHtsqb2cn6Wc529tONcBB1TG0ru8FQWe/Ys6BPpDg1xk/POVsRQF
F/4atXWZIZ+C5kxvDRsriEyNAJQ/Gt5PoQj7Gptor/ZLFUVVEKbWTnAWC5RHhNcO
Zu4fY9hfZBYBTVUgIH2vOephDyqS2ClhhLkrR/HCLZhNByHKoqbDhrvo+NEP8cbe
1Ocr5od6Bj4OScnHRNxXI/YLy66AmQTXT4A1TRUK6eZWY4qDuyWvVPsuLT2MsdKc
3lC0jsZg0YVyjhOzMtuH+QTrEcCZFQikENiSc3JAXCjY1rZpoG3OBbJ1DIfKSidb
9/xqXHaf0DsT/Wwjc1cODkC1ytNfs4Y/1Stc3MzYqpTD68ljrZTA+BRYiS0BKCwC
6yjPeeswURAEdYXNI3uwcBYOU08l0y1T0UTCAcKuuCFuR7LxdP6USKSVim3//ewU
EY6+yc3jYwpNXx9gjCa6K697yO/N+mPgybERINf23d3q4e7YoDVP3//BpEnfAUis
ylovJj/eeqLhOs7L4T2uiP/EA7GVcz6ADKjvkFqSopmhQasZAzjR7BpI2JMEWVhD
ziY/wGsZFwshJxq9WZHFKe1K4AC7QL6xt6OBeHmwScirhD0SbtX+6QBZR0xL2+co
M51NIyQJwyhxMnNvCIx6n7wjoFWnlBWadAACuhNexbHp+pswHzswj/UPS1uWKrDz
Np/t+//OlVjUUN6ImF8LpL2sDxDMj9BczMQyB59Is9oUxlxtqsdxJnoEwH304c1A
qU+uF/fBFQv2NzHZl7zRO0wUOCYD+iducr6srlOZ2x5Qcv3/T71wFkuzyTQR6Ab+
mVAPe3H4tZGLDQ0ZgNYH2u/EzxrrhGRmmpxgiQwFp2i0fq46fgfq8662tqZWhQbc
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
MAP7F0d7XSbBqYSvUdqb1XoN9CGnYDaiRucVBNf66wJNhiWJ+CPq1AjND66/lMXX
7F8tc0Gdv7zJsXsgE6LDL9jRdweNbhOK2KGzssWgJuQ/q9gzVecmklU+SVMX9AGs
TvfBiU95DF57q/Kd/yaclnsW7NxQAOKztUGA61RAgE4fMueMQ5sNn4DLxenyyimz
S3zLOzXLrSOCUJHI2GGGPOLGAx3cTQUfcKkNjePAs9lONzQy06DAz7lQ2/nRJBrg
53nlpAWJx4PT90MKL5lVaEvdr5lVHJF0bLsfAaT/cIlc90wDYCk5FOo4oat3c2Z8
tqxhTlrfRRE63zHJzqyH2Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17376 )
`pragma protect data_block
ZWD4g5AtLy3ktasCerbZ5wNTcoxbw632hnOHQ+915FfZg71sOcs5K3/YTFKtM8pv
MZFUc5ozuKT+GRgccak2s4krd0Z5IIg5MycZ3bCOa5kEjZjgdch46GchFB+Efnb8
dpFav7zjNVraKaxtNWUQn5KcGqRcjWdWmTIqH+pQeH5ztxjuoM9iUq+Niy3Y8DS1
MjQa1Ct8h8s/r/LLzL0MKLShY+OXbeCfC2eWeMS/wX3xcLmU/2UPm5cuAqL4dDnp
GE/W/9Yr/YEIipvctVt8c7wWEnQ1y98/xvDHLVy5EcMySrxkZU5ydY6I0JS+r9JJ
EE41Bq9APfB6MA/2Gje66O04+l8051KfV4jMRPht7n2Wyih0ELAvmmEdqKx4CCyU
CgoCh5Vk4NHwl5HWOcA5mAmQg7n+/46VNfzxIHJfDuP8rlmM5pHX8bnlpaMpNdTT
h54QkDF5pxOm2xWtrDfNaYgKo5qcxt4FKzfrxUuBN60EjAEANgKlWlb1+cvSkdZ8
8YqsddeZtbUFGI7YjiLpA/gfmwzNSWa5010TNzCSt3e+23kvMGE1CDClJge+Ippz
7Cyq2WFEr+fFw8EcvOoS1YAEmE82unuAt2e53lrirjT+N8zG5mh0QUlYV21M23rh
ufyG6Gzto3ARqUz7x2smoGjlr/fHn8QViI2G4tKeHPZv1U0g3O/2KaPNKo3VYHJg
buhEK+32gIVcG2/Eli6AIOedVQ4yw14L673vJJaGC5yRLf9gWlhSH2wJ1HrzfiL5
gfB2kvln7v+TNnYzaYbnk6EMoox743WXPwsfiF0gAnRk7SnYt9f+GcEKEUAh0WiN
9d59/alAOrntLMWYicpEahxHYS0I1sPnd5ybwmmxISi1Aa36GevZyDr2jdx35HmX
0Wr3qAJzvTVlrMovrOvyoUTZLhw3o9wFWCKb0wiNGV1UNr3JG52MSGLjt68eWOFc
EO9oiurDiyWBXwtg/bG7O/7pAYHZ8r3sVp1AG/Hnzk3nBVpCetobBe/C5PRkhrJk
9S+X6LQztUS6H0ARDhe6wIzoJthEYz1agk8MiyqYkZAr2AOpLTOZPQiurIrr0+jH
tx/aqygezS/buHXif4u2KgbvpZ6J1fBKjBD55xUJq4R1/abij/HfF+dMln4fUfq2
2gLCw6tgdcjAT6GWHmtLd5DuUYjU3k14tqokQ059SLu3K9qMXlIsXMOBtR+83vl8
0gy0+f0NrK3bisvQn9/oqX45/sPMWPSH8BP9NJzsFpgDs4QlFTJlWi2UMuCxtDNp
xvWgJk/r5ZWWItGIA/navhbP3CiLPAahtQSO9TnkN+CBD8Cd4An5ASbn6pgfJDrU
d3xEBMcm8SnyLTP93JTPMRGeSbsVZQiZVoCfoGJrHsg6r8F+FJ6OJCYJbmceQNkD
lS5ZSE1GH3Z0DPYSyhonHewAQjgyflfZp/x9i76UbYqiOAYHaiYlPoP+UXHXvLXM
dEJ8a2wVZtT4bTBVlZUZ1jk3CPW1xKjwjJrxT2qGakaAnjBqiI3M+cwoc8iXv4bO
ga9XZoyVwC8iZLzaUyc3R6WyAzJD0wyHz3pwvb7YkC0GNAwdcwtbF27MQTD8m4rz
YGu2JagWU0ShfpzPxu3+g9zWNxWsqyO0le87UWi9rapzNOcwI7RWlOI5vl+cvAfL
C264zqDTra1z371xejIgmEECB1DmU9NqL75BnUPWkF64XfbK2Sw28aTsKTJu30LD
3fbN6/ojw/pfuu1I/+XNtLTBhWslIaF3KHe8uqEnPaePX5lrVYln9Ly3gbqOXI3I
zuivxnYD5AQ6jZDDxvdTSZkh1ZgE3VvcI7lihnH8UaBTzWJ2PaXRZcW6xgbq/0yY
hnSaYBRkLviKi5U7prmIeNtj+HWnoMYVy4UiSJ0P2tuqYT4/678FPlZP1nKI6upO
9Ew/sCWZj+QZizKeOSd4/oQPHLFjfignu16KWytHu650Xid2ztFe31m6R8UDT1bC
N38+XFfO/6BO4Pn9Uth4TmX48fja3tlENtVoKfrRPp0No1eznQ/70/7BbQ1M8rvw
4BfHRu+08ARikzUx9knMEPg2U1SiaKukcHo4nAmiVhWm4zsgPIE1QlgqNyEpevLA
npwwjDhI1+Vj/AO9VOVkVWTi5IFv+7cNP+vKNVt4Vid3VN3Mb8g4aTp7aoytvGbY
QM8z4mdP+3qHf7R1LGbvdZU4wKMcGSNgXIqZQCqbCqvd5Whowd8SeCCGgI1PG3ie
G8ibMV0xYeENTPRs5yYSk7jH91YzQH53wBUBteVN90Id79JOJRq9pxdYTfugn/2f
o8ElWhoweiqKK+MsALRrrQ+/rGsLWKJsZ4O2fvlxFp4N9Z29nOjX+qZpLRvWHVu+
ft8apLzo7H3kd/NfKyCPdE9B8WuewyxuJTr9yjRMQ+GYtJhiLy7/9YftR1fibMw9
75vzwmpIVTQpI5vD8GyIn9KgpHaRUgBm8Qb2JUjEmJYeN9lvPz+8wfi3x8rOMHno
6dkmXy0egzmoYpENNVsXO9l4YtNmqJDUlTfDlGtFZ4jtzS6NsgBRG7etivHzeaSO
sUJJ0x2xp979aQE/pS+TSVa4QsYVQauvUNKXKJtKtRNIzDk7u7hCOfmPmLJx1lLA
xd7hMEYSBIjWLDAl5O37oYa8kaN7oX5yOhFEbUlk6+KGbjfw45O6ANF1lL1PtVd9
B/TNGqYhLfmvl9mCKGr6QqYi88054mCF+IXBbLAQdkBcOafNdDecLW/uRC0o6Oik
IDenp3C6NitZ1m4kqx0tvirB7CDf/Q84+arvGaQNVaTaGjB39ByrbEzB7NlAnYBy
COfJp1LzWt6S1yx6mCwWqcD5JNvMvLhXSPlzUvVqfO64+zmf8J2jAK7tqM+9Hbvj
rpcEzVAyU3qVyADCiYqEquXFj/Qt29Kgxf9YC0gDf4B2hrG1zGC53goGlGV92ZWu
w61d16Hv7PqbBz4Z8PRPG6uMycRW6MQiMWOTYz8JsX+Dyb8S59vBbj7158WF0JNM
VjLHK4kFCVvIaVjCLP1U+Hl+4iw9cuyz+NeeQbda5ukj8FUmM0cHC39UhR5mEro/
C0+6fo/S7lkdQAAqDSKbJfCCvIkpoIrHaD7PJuIGlHXeFPuOMuFsynHzXxL+FMJ9
mv7Nib64+iWp9yuVXfZIYkC1djFxKFAq+me4TL6xG0br1Ue2w1gt9VtSWzOCKY4+
o3nxzaH3evuzq4SxLVzjXULHC2hzWely7dVxV0mPZM4diN+t9q+uo7xm5lE7imqm
KP1qdqgqO1bYHIJEfsbHv6iufqY5rS9Y2JtfbLqccm4naOMRMNwhhcOsFsC+1Ddh
j+STcWWNKkYBmlZPMZbq0AAQnm8KNl4wctdeTvdiZOBsBYEWebTSTNPZAHO1rif6
vUvNQiPEmz16J79TnYUcd4KPw4DTno48mV6WumsKytGQWhKETjztRzxeRMGaRY9A
oGx0tBwkAi6N5S5/nCcQ7fVebpXi+ZS517W6iO8ZJn3Y83SImNtkwEv43aXhmNGQ
02dDB/X3nk3nRABRgLhE7TuzKh+7VxU5eClJx6pRBwl+UbIXiJ4wBss2XAv99fT5
XjhYMd4/IYSHh0J8KLwCBiEbatBsoBvS4yr6srld5U/1kyuGkvcirdVgC3uROgui
JLu6tKbc1NSGEI+QJQmet5RDy7psoCLDWtqdTgFd3TSrjqpZ+IkwTtiWDNmQOzVz
gXnDxlnuOTeZ680T2YLFLcOlVEuvaaZQxFs+7lr89HCnYU5CTE9tVdzLJWZxU0T/
z44fb/B7aMFX67/WOaFH+N4GTSr6jGt3HQR7ds/kyVfV17823cKva9DgdSew7Urn
qhxDnHKqxdC375ENgHM3sfCHxLWI6HC1RQdfh56LDw5bmwbB71bqBfbvYzTOTnZD
XdMWXLjzqq3kJKxGk1KvQui/qmbmgtysnljugPuBWHWQhMBFlyZ9O8m4hHOr2gsw
BDrpGssgztmmYET5JWJTRA0rIaw9nkIsF3cOtZ5IRVt+0OErvsV5CsKahuptMdEs
IxO6leJtKqec/WxI2g68/Vlwi9uglAql/G5GRM476OzOb447OXZ0FF6P0HwiTdtd
6LZf3vQdVDLm4y8YwlKag2kFGg2ZrcjRDV4/TNtTHuUaOKn8a60h2fbqLoJq9O/3
1qTWykDYS5Aey30wWEn5s4a/YHBFklAKULdjrMeOV3dKC34fBJby0rZUwSKFBCJe
K3H/21L9igbSm4Wb0pqcjbohD4T2Ho0LjuzZBIwf6lyNkbkH/8TRVO2t+f6yQ2Of
Q7DYMPxT3hr5XllzBU+FAk5mnojIvXj7SU5UB8C6q78HamrGUSP/a7c5g1lSC20r
jkD/uokhmOZ6M65ksYpXdm49jr3azYSe6WyLfC+BiTmv6kv+RtlTW9B5uK3Dy3ut
McFKvHpEmuRVYXMj3PptXD1n+PpS04oBQJ2d/uLAd6mq3rg5w3wXi+C8hq39pXKE
Jcgzm0Hykp3Sr7xeX8EH9wjyXRybtFL5y+Ql5hBlTLXhAD0GZjGtABQ/XuYafcd0
nKHrPg4vgZUWBh7Ohyr1/qgy8Q6QImoYt9y8L1bATEJSTqoGrveaoAz+RMo7A+qE
RoE6OOhbQvnmykIGbAGn7CHdQMejAGp+bPs8nBl59SgdCnE5Di0Aj3ycjQUtz9M0
H8yzbStLonc3LX3gjc9St4yGdhjSD3XyjlzWJtJsCGENKOOPtJi07M0sHkyaN+Rk
sYbYGE6bMObY/0MMD+0R0vk3ex4M0HzdyTil3XlvdE/t1wO/bUU5OuxfPRMwHXWg
W1ZaMq0o3QKHlnZLFncoLTA5gBSQ8weTGBGf8sWEXpIJULaL4HmynXfUCbfoEiRU
aKgPeyEOkzUOd9dreCVGuVW0qcj67lYo8Z81QXjHIjrytEGoRcZLPRRx5xHIrh+g
4NJScKlBhn6BduH8+RzrzcDMSc2Q3MFBSMNQYFESD/3ojyskGtdTopRNmJq2/X/j
Sa3cPhc3YaSHC/LKmV/35cJHSF4LRFIvoA5bGNlhr5BCzMpmDXDTdWIl1+Nt58Ms
/CaSM2wjLyxPkAIO8Ipqh60sb3JFTke0iWmHIGVv/dFAf/VjXsV+dGQCfQy+7wti
ajstmLKwDcw3MMkWeiTJjPylPFCUL23DFj5ZKWgseffx/6ibQWFcGJF+8V4wc8mi
VhVD9humHXOXJ1jKJK6VCX0c11F6NsbbyskyXzGnETaZTAhQmBpjNaz7tubaJqNV
0zVH7bA+GigLgKXaLssJRGkJa/QXq8j8bo6aDE/LHkuoLX5xnUtNafQEds4gG2tH
oQc40hSc0TNd8w0zQ01RNyY0CMAo1fvuaiOEwW/h3C+khmVBsd96IAmmQEDImhLJ
r0C7y9iTEaVIxNvz+dFCyUy+3BGGfCZVGeBVBD9B8/Vl91d1MC1Y++B9W/6WkocX
90v2PyHpvcSSEzinLZnONSWgLATtWpGSXjnHmWXouD85CDfOhw46y8HfyrWgnOjY
aH5ZGp24ls8Ndj4bJ9JP35vJaZQqWOIIxiVPeEMvUKi123EL/7ao9Quu68+g1yys
5+gEhYyZ45SBAwz0visxlQ0UghCvVGa6e16JWMEs2FeBGjEFHAC9hbEGESHqWOlX
C8XYbTVeuIt6BzzWFqHHHTYU6E0QybFg8TYvesecTQB5YyRK1t/cTi/x/+QTdVrh
81Z+80/6gX+W9LSVv+xK4O+lGdB8cQbWQehws14u9z20eFZHRYyTZGa2J643vUqc
BI/kVi7aZ8r0GgyhyEFUF2Ycly8B6s5Xvl8j1mek9gihep2MDFtqoMv9o7/kswvK
eHPYCY0nS/g++eJeZCCDe9v7gxIGy/Dtz5azlq2glIEF3lnR8ByPJNMI4Nlw5J62
kXZyPGYHSMbQ2P3UlvIKE8UHvdo0XyfaVj17SMjwAzf7Uo09agRGNpXy8PmDil99
gBiI7zlj2Jq7iRykpHxYAauz5yW6Qs0ka61rfZnC2k9WWYlN3Rb66ydslLSoujg6
DflhvxblhXMgsVfuY+QqttnTv3BKGtkAbVY8nYwi6bzmY/KEYk5SuXhZ4csyhHXY
WkCnixPxB/exqH4BHe/EGDU791CvWqgJfgQBJsPUpkS/lT4rtvIhEmTMHTGL3ddd
4DvFxBLBXDTipUTktGHyTb2MHt9D9dM4Tzyq8/lhHNZGS/6AiDt4da9pbSsZfKXF
U6w/YJGjt/UaNmExpq2J7Rh6Bu3QCOpEhR27omqbeG9iOwgzQqhWVV9CX13IT0ML
p2NfRaP09hgVtYyOSZTsK5eBKBE1TtKmxxlZTmSkrsrIqVR7QswspyX77Gogsa0g
gCjTXh5+8lLeA4+ZpyE8TMNJrYUSkyD29H4mpgylGk4tLYR9gdqk1iacZl2VZl/8
Q8U+fR3EjQmusTY8HHzrn8JJJpIjAEEw00PQs/zpUuaRiyXB4S6a0yS34bpFh5uj
QAudSq8RF4IGYq/Un3r7T0PII+AKlNBSd2oWtflbs9hNLgPlFJ3dZxDCPYKKmd3A
OKLSCBXidF4VdWtDMkfhC0+869OnYJd/v50zfYwBHsDt0FiXzkNDtebBOV4RT2fH
KC3DSxRaXVVseUl+ktTgumYjsmPysXfqWAyOTJfWHjCch4m05DeKIjGMJIKjQI5l
G7fB+JDjj3DNm0p3+Fn3ZV/piekWz8lHLh/zunj/OOfaLu+YVnIg5h9OfFCRR347
kCefkxSQ2nlKFMxz6BXZVNcmK/cXdO+vjI1XBmEOY2u9wHX+5nvr59QoZPpj1463
YGBuYQDz/iGaWkzYcu4oIp500xDA//0lLhYfkcwrtIfaf5sVkykUCe/HReYWS9Ep
u0zlYFPVAqVTXJPvTN/9+fjefxAbQn5LlLadGirLDKaq1gTCyNVM6MHXfTi/WeSo
HETrq7r7bCNfQuzjRMo3TWEXrXmxcaMdFcKOnLagx2yRAvN7db+saKYLcg5N1/HR
HQ7nJQF/h7Tp7tGO9/ZaYB7HnZZ1NwiZkiMBhGWIOEk3rQpfKZYYocJaQiAF4b7U
o/EXcNnPKMwgFKNpIOpdhGk5gigqUD0iMrM0ZWaxaBeXVVYE2Y61qXgoP6Op2Zta
5Quxi9BRKnASG/ogNncDODmW7A56eRM+H6QidUy7vrNDOmO6ObgLezb0C2hfDm5d
U/vToeORgct1ZFY05VTC8r3/xWPCp67JMTSg1/WxdsFfqneYAZqsUa2R++slU0+L
0EWBTf9kCw6F/ozPAiowAf7/EqWQbpt7PHXVhy1VQICmAI+OzkA7o/XRwvqyHPgM
z5D89hpyyZQYcYUEG7BUXvYplV+r8ktIDH5HT5iqRmcDyhykyWleQwup/XVTyvpk
IA9B67hZZR6MDStBHT40yB4oa3ok9FbOaZQYXv87ZeVe1+bNIVHYnahzOcjqUYRz
16Qg2G2AMIiw+vYxAkaxyC0k9V7pY6q2alAoLogtHc0oxjPnIjUqVO/ahnbAs0kp
XCocRbheE+vYX+2CsKN2qno0HXFLvH5j14ZBIrLlWVUI/xn9furBlQ9HEJXNlmFt
72vSHCHRpe3Go87+dfmCiYhQEnsIsBB0qMBZkNIVaa3R6oLEvVZT6DD3vzrjKEw4
ZFHy6NC9rv9l3JE8SN6CiM8kPTF/O0P3iBf+FFdlolLPUoj3jkzl3qOC7ZZWY8kM
0Pgz6PsAD2VA9UmVAkvoHK9P1ZoHdA+RO8NWpbDAU6iWfp5T8uKMnZLM0jf5JAP5
gE91J7sA7y4tiElI7qdgFW6mZw2OSF9/yxkiu+8LgA9o2Krx4Q4D4ND0mOvRkYcx
669uLSTHvwL1Sg4q55ToiyDxvFNmPTqk5GSJwgrfdzYYKay4jvLNjseRmw/qHqzs
jsPb3OiP9+FgSNwOh8GY3r7LLrzljuGSpOvR0ipBXYN6JczhaTidZGxrBHmbafhL
PthExkTPPxTFAQlfRThNkZgD/GFoLjYxQi0lRrB2o5B1tM26iA6pI/d2lW/AQ+eD
vTq+jG/JW7a5S8lroKeqHeGGB69HZIz+NV1maYqKqQq0l5nmRrHTxUvWeNA3s8I+
hTYZSMlVlWS0SKZdSW8Nbi8OlMffF9Sk+hGIBj1Kx8uJBC9l1houZf2KyqoJhivy
p70evYGSMvw6v58mgkSHEjcsiSLYd6X8aFkMdbcOv+QQXx4q9JZ5NsaTTTsFSTMt
YatOAaLMaNYx9HOX2PmWgErz0vd6kS+bcep4x1ZPcE9Ux/iWXk8GmC5DOQt30PVm
t6wnlxdeMEPsdYRGkDDMyj9J0aLqibLbWmTrwLZFD+VjSRDSOnDvlFf+MRxNRPOn
DiI6AuE69QVsA2lvPGnxj+xG+Cf8fdMmG3CYXIYFe8TxzCZGHFMhA2TerriynYsa
j8Anb7GhbHvp9KNXrwI9hyNMXuvNiEVRBz+0TuYZIVIQ24pOpjEv1gq3hRFe84zu
5I2IEP9XgsTg7hgqyUEUlMuMYC2GfHEd+7eHSq8q+YiDTdTniBMp6lVq6CL7nlXM
8Vh4p6S1DWft5rl+ae4sXyw4Po6KAYkuzBPcy7NwTm84yP6I4rW/53lmiTBs1aA0
rJgw4WgCA/XJeD5Gv4w+e+wWnVYWS9tGfUPdeSOjOSB4e2znNV+VuGic9NQ/BNDV
bHivylJWOZDHQt+t51Ntnv5JHur7cc4NWUJRBlUjqO8XHCyaIvVmOOck11gwV7MN
6P6xRV4lfB8W2hVew30SqouFmxmYpmTltzbY4BhgOdaCdCXs4x5dune4UBKWfvMn
9u0UdYowBGQ5gEvs3fXk9trUI1XcxQDJhP9b3Bnf0CT1YGli1zcUujsagyNUA3mM
RXqOX3njtErgcNczcie1/2BTY49UYexJ9C49yyCvOT4rNJrvBXkidHBKmrhuYBEX
WzEgWLXkKwioth1JGLiv/iMHSmzsbCG0MBEhdIXkO0+AT5b02xTUTdpmiUSt+qur
gmQL88gZRELngL7IvbqzGePS+DG9SHGTlXcaPIpGlnSuZ8NDpFY2hza3/DdxG3xI
fBi5r2Jrhbbnri7CMqf2rqSkB147FJuYFnZ+gaYhXg9GjoBu0dcFulK8jKflY6J8
RVfsk5uxXwS5ZYBpeZu25wDTJUyg2FzKbfAFkFbUleybM8ql+kjdtX2Q+MU1oFSQ
07ss4hGcy5IdI0htswpalnVzSKoTRaH26o/dNWLtJS5RpFSwoP8BVBGQ4LkiKxn9
0Qa3Ku3Ug2Q96ubQN4MjmZk5Gje2/w4CTW9NK5MWC0ltmOiV+mEpK77ZtPnpKCTN
D3TMqfqelTKJfyghdiIKsP7zd+CGroULAtkofIFioa9bZ6pdiiz2u3bgHDZMUy24
QP0xg8TFxjpHhPGY8Mew5MZljS2yq43b8hZ7AolNMMovGhk95GhMwdgQd3Z2PBNu
MvcUQ2nTcQcsQuTjrcOPgcili4LyuMrmXMsTpw0IUNniS8jq6TaNgckRykd79ENr
PiRV5MdzeI84LQIufPzpsfOhCyYOBPiZg5sg6ztl5As9eOLISF++9kejRRYJUEF/
ZNgrlsjI0SMPtn4SZfP/hPQUM+4Adg5z2NvPoTCGEh3W5R6J7nRoKugiC59CAhzm
lT1FOHZAJTrd16XQRO8yHXqwOLkqIhKRQ00YOtB0rrKhevq9TUQhHuOSXK6qbhV7
HPayRTbPNv/fvt6BweSRMGGdneoQzM+RoKszCHht7o+M2QKszkAU8W4pafMM4I85
PH709ZbT8fddqESBGOu1XQJryn+9Pa1x/vjGMVPPNwvJUZBYrk3dsDaGWLffliRV
NiQ2DRrzRmemgCGJrAvBxwPxZ9o4LPrZGGormRDJmjpLc0XrvHfnFDkrM19gHoa3
9LgSYGjjzyTRpULrKzTBxmkKt+NXDNDZqIBCnjcNoGwUZXXG1it5JK4MKG+cHHNR
z6iZm9Oz0DiRletWJG4rACLlfschklPNZP7h/7KFkHOCU9udCmrvhg0OgkXpQFO7
jjPtwJqxvyESY6rco5L4p3kSQQvBBlgAlBLmGgPe++8jqBc8uyLZpggEcwgILvNH
vfAufPPsQcweFE8XPyM7lHrjsK929MzzvdKG8hKWclCyfwKsqlym+/CHq2xo4PQ8
6FYl4hmPSL8Rm3z2a32MoMuoF4+UGxdYB/jJu4XseNEUHXofIufJoxSIi9Zkpugg
0p2t1EK9XepLS4jn7GPv3WmUKLkyNLsZJpl8UVVPmRFzAy1lxBgoh7/axYkpfPG6
eV+VVhBS1QyPjwWlEyO3G197kAuIAL3K82EkwLvluPG/AsaiL2nnnas8ab3jWCJB
APCEciuW6FgwVj6riOgXpbFauRy5Iu06003tJaAMaXhpAVfeQ+fqITorU1XsHhDv
J8pNeBXzwj5sBytK/ep+yonKfml5rLZz8n/EgTowCmL+hM2MPOzjQjrhw4H0R+r6
GbL4zNgH3q74BITZot8Q9txtRcVnWgYr8e45ZE+9NEs/MJiL3yNgdGfT/gVWlMyu
sZcYwowhG7miDg01TZZ1u6IcY7MwIQhZPMDs+brA1G2uCKHdKroNs+t7ao5lUHqq
zI/P8IX5aiVTJTgdur//3TNPdg8X5xiS31jneB2VNMCHqG+t9qhbSNi3tLFPqob8
WIh9M9z4ipolvUrpy85vMUMVdwAeK9tkIINNY0UFc7HOqkGF/4M1tpZ2fktx+oL/
U0jzwaRYK+/cVleTTb9z9jCP1z3u2jBoM6fFQo44XFDk+HLGS6lxPnAPUquyyI1l
gAKv3aAdBwRJ4FP4kHnhyMsQszzU+n8h+gxJjAVwz8hRjJtL3NE3d9FCYezobjV2
OuVC2y269mo/NoGdLbng2S7+k8eJajgt7Q0TPxm489c6ci5+W3QaB5htaBRHArdd
mWHt6R9kBIxmxwaI0PQmmAWZzkRZo0AuBJoWq68WIR7gO9poq4PF4zFLzE/ZDuHH
KCcsUHzwzzl9OeU4IbEhIf6o9Hozg6iX0R1uKZ8aSASCfQolk9KtRHh1ajlYxGM6
Zd2dXbGh7gSl1h68A1Lm2Y7r/g01CRP78RNolnbbL2Mj6lnYMqlVhLnt5Q8YsqUm
sfCtu19HKj6o2qRb10AJ1V8V1iFF5xyohF9iQ6ukMdNRtUFQ+LR1ayKqHFgsp8p9
r9WVPWL9YOmGT++IJ/nTBwX/j5GJHxgnGu+KCY/pBG2uFFxdKBIfrpxrTCFBmTC2
d23eT01oqaZ+3aptSxj98rfgYiU41TmSl7ruFzwQFnVvf3y7sHdNU3x1v6bfR5MS
c4hgkV06Y6Xb/7vdi5v4snZ8DNDeOW3EJckVKVoRdoFrqQL9+AAzU27T8AERdU0T
TaMQLkAX0H5ywjLIJGlx6Mcqh7fwuPSRRYsakTTDel01lELmukEvdBZ6CCVn9JTL
f7vtyjiT4nGv0HWnXmGsF62D6FZ0IGcsJkhDNY4wldEnSJUfmSznOGjP2+eV+74N
yyaXwRC6AAlcV0Ryq6XzBqsy2IRI6iGCJqNjpxXJyanbqA3Mz/WNp+aCotyusPQD
TKmmTXecw9v8O8onu3UsJJLx0NOAmhH0celW0GnPBt8XXbf+sWkfqi9P3+/4FtK7
7E/h9hoK3KT3kLn54r8a3VuiXs7tM7a0CTJ3mWZPFw8nrWNnla5QEupl0zq4xS2u
y7oOnttHQ8NXnZREsRulWhvzn57SGKtmOx4pQCJooLZDdvsB1AFyr5A3jLEqH4un
aMyvWowSjwVlvLAeAmWjF69iybuqxUm0YJUpj+7Y4kk6B99y0JWEEriAmAFrcp/u
XXslP2Zbemtq3RCciTIBTAoou8e5x+XI/TeYe2pwXep5MjE+9IFFaRF6aTAYd45g
NzmR3rAqajEPsBPWxmRhArwb9VyHVWPLBN5sVKoBYojeQwUcKNKXUdMY2e7MLvVl
4xaLLbGeVaiqBGRT1XdV2M9dZGp/HGhwlEBmVkuVABHCjxpc9u69/qpVS2dl2ffX
/cCD4Rr107kvSvcZzCAH8THLGA1WAluoaGQEkmBYHn52kdGkY927MGaDk6Y7fzpp
W+GBSsWaViivqEipxa4cAP7ZvizQrKtSlmqIqTWJy/o7hjH8Jougpve5WfrIYdla
H4WSzdGihtiKrWg4gcFSsITBo0vlk4SD3DNax2/BjPXztI13eUpdEVsBobntsI2X
W4Q2MZNl7dRap0aIsvnUcIGO5osXi3qch6QpMbGWSuH4s09Q8YV2sTTx60I32TZ1
5LFSKeoY31VagUsFE+eE4Fq3cuWueKh279LnL07PREkaCi1RZ0y6TRQLCy+2yeJI
kfKtxlkT8YfYuQIAI3E6cmzFEtScnga2A0k3iSX2JbDxzrlSH4ssd7jiq5naOugy
NCzZaE5hzc1vvCtv2aE5DEqVOPHyrqjQMviWcKfFZwukz2qu1H7oi4s8V1sxQadn
0/OnHdUoJBlK5GyPEy3bG5EqG/RjLqO17XH5KgTzeJIHlAN4FYUAcIf70Gn5Yu8V
XWo4AbGesznGgnaYI3QRh2P85dyvDM0xQoOgrvTviNDuhFctSBAbmTkkfHDN3Gig
dbhg1xVQsD1Aicr3yA2lnOFkL2Sbm3Fsw4670eolCzIvmax0nnezjLwqpcJkSYVu
WY6S/M8nLXiIGNlFhg6gOhnu9i8HS693cRqdM3mfa2CO9K3URlNsqyesnraOSGNx
snIsu4/LViwVB65OMUDogHQsZIe2qE9I0/Uxbt5ab5lVI/Mz1ZqGbkAL038wugXc
MeMT5wJ81N0iVRNFzuNaY6ly3HPer7RT5asYZ8w4U2U76oYlgrmj88Xt5kBkU99X
047VXTIjCI8691/werjfUZSNac6rNKbUGveAbDmfaZx24FQmzEAyQjvcMUOBcFvQ
6MtdUeaItkulCfm7nGRmAWek51GAKo581oyjwj3YfJs+q2oJbja6ooZ3x0A00DBt
PYuQhm/5vfrN5bFXmi6fmonLagVZCeFN6LJGa0MaCo/TiLF2tJEdygSJill6IZG/
XPNkmJatQIUlv/0E3+bWmWEjpJ+c4xbEdKRA7bKj/RHktxA1VEGkZ/Cvef6X9YWJ
RHqKa6Q2kgNTfjZLPiW8x1qKjRR6PvoXHVzc4VOgoLmQD1gajOk4IMUAuZEIj3hm
e3r7GKtTJaf1GyI7n2z/+ixldqOOcyUg86hKs1sFWfuE7hWlBkC6oH9SH6S14hMe
1QvqK3LCW5rtkyV2hwAor6qx8GbpKBHHakabQGoHsxLEs2fIJxYdr+sJHYicPv0L
Julmmyg/VWGtquDvyvRZynhmD1UygAtXzkEgyC6oakDp/f9QXYzUR3wYjV0nYoSN
JrlL718offJwyedQIwMf6azFVg4bcj75gA8c+Oi6fpb9xUwKsnI+CkdRIF68pgjo
v2/tVJpeozYFxC8CpedUgpISWwnDlQfiIaL+932USqVFvzRK0p8T4UI6VwO8ZU23
GHvSTBhOtCkdjU9ZqIuYuueOa4+tg1fXd2CmNzS+Xx5YzoW9dCUAG2HMDusvyN7P
CauHtJ3auZuF10p5uwD79zVMvWST+oYRp+5sjXJaTua6VJMyB31Kp9yYisBQxht6
4eiQdEN00Tpbhps+ZfWUVx0cuiGZzPMICxQZBA0VXi0jOJBpNyJ3/OE/WFp5pS9R
FNQEQMpS4Hux+xcCIBpzJdMKx+mE7oATH9sL4rkO/LNFsD/wxXnBbmrp2dV5q5Wq
LsRoFO3BfL29dKVcd5CeCLLg3w1VHanFTju0Wa9RCsf8ZdaMthDxHQgS77PmUt9l
2TRaES2y2yRmxri2dQoSM/muZ9hzKig4js10NO4Ce8v3JRfO8E1LAMj9dYrq1Hu2
Jc73dRIcNBN2gdwdzperpC6ytgWv2Bhbuml+VpJU9x8PxxGPaCHqtECWuJdvhb34
TmjIATMkHd36j8aVgPPgFx1+V819b6CRAFAlwrv3Ol1jTN6XVkynBuq3diZO8c/s
838Gpy3IBM+GX4JdVf5DLIbXGjaztT/uL+fABJovBsahro6pvG88jnfsahU2huBh
7lgX1+gLmrCWqrOciBeCPc/uZ9YB5VbxklJVTtLnwDqSimuSYrBvWTwxmpmWwkHE
fxk60a0lIszGvMyI/J3v+cvJRinD0Ujxj9ULAY2jTR6OrdAAs8Ojg6VqW253ti6t
xWhtNsYtntJsUH6OGWemba1cNOH4pZd+bZa1XfhW71msc7nWdINADe/xHyfvY3Qb
fw4YgkUzdJ2xLJ61y04aZzuGCUYEO18rzse26gC9mcQIeqMWwoqqgLrzK3MpxyNt
+68a8GDhLzFuRgpJ5VQAXu1ZK669UrjieKpjAIZVe974DUXOdDxMd4K/cRjivlgu
R3H/FqAK6+zRgp22ASX/1qVScJKciVOkLHriliPZT5Idq/Hg2qZbOq3rMmDC8mSu
BiBR6CnktjO1vqOKfM0+5ZCj/GV5WMkM7/W92EYoHO0Z6j6lwGZe7LThDy4VlqUM
aAlcR7zr2lIbNVjc0Rt5PL9L2+If3L7iSPt+n8ifq5q/tRlNWJPJdQ/zZzjg+GZh
zuyJqnXB350s0qhgZgdGabmvDbtAcikPgQq6leUyAHFVzGqPzL3U4DWskj9h7mm+
kOt0pJLyNH4eFwR0nYquBgIM+s0Dp96nmkjLmcXmO5boefsgD49j8U0Y7mUCnE23
BJ+6zOcuBZQw7WlOz3JAEWXVUFVpFXTPSmGHleD8XcVHMBI+TZSMjG6GQumauovj
lRf8U4dpJeUe9Cf+i4dBDSiqUfp7z1bnn/hMj50s8RXaCkoXUzsNmXqztwdhvJca
yUQB6wlPGHuN3AyXgkqMaIncLrEdqStgFCn7B8mKIqPxQGt+pQBloJtYgaFJX2Qd
ijJ/KYErZHpDCf21ZpCxFencnOnaGRKhL4ov3lq1S5xWueaKcFzEqTJyahm2nU8+
tLunejrA/z8UYCTPf7+9ruuzZWxucG+yFIOvICriYPfrHD7zYTxaQo0pnDRCJXFO
jNAKqCYIRqPDlR0MzJwSIDsdS/OnGUP5lQMF98yiwprpqaCXBE1a7zHMB/OQfmS7
rARf1+LPLoWkPw/BK/FgyB0V+ra+2wU8d5C/pYxvO2LDFLhQB/bUnW+pjNjJpmKx
YBX3Y4cejwDMEtr6IlUhwHt2FHSHSBzvmupBiDyu0uI2EDgmwI16jiJjHLl0x2gf
6/ImUoZJG93MWt8nxeYjE/F6f4EVaNC1IfelwBuDp0/mO/7/L9ezaaR0wfjUpP9L
d1gSklM5hHK+H2MT7nQWjmebp7EKxxEpIL3rIJ3y/gV7rZ3OgFygHIZ3uvzdJoQb
/WyROC+1rK/g4plIXvL6tmIdml+/HuJCjtaegWnPEMrnR3N3fFh/zeY9pb94rbjY
taHd844EY0NyMzWxgS084yVvCTPDrSDHKeGDZ/aAsKKwHTpL1jHSB8vzVgDbbzCF
/bIMS9/OaR+OxqjYgi30asMV2JAzFqBWaHmaa60HgoBOm204Q+ZYXoOSu2QjRZ6j
61xshsxqSFfGt5rzpI3Hn77ZebIe6gvBDCDQf5Q6cemomnGDuJstKjWzVSmaV73P
5I6xwHW7iwasnLQoYT+ZIfFpaVto4VJUDAvET4CIcMZpXwR9shHcEsH/4MBfjPnH
iaPB8MnSSsR3VIHGUZznSBAUwWaMmhtWpfo0eRYKEiZTTcolHGD2I8Z/NaFuAeZS
RFKhkE7gskArsx7zWkozszSnca6DJAnSM+yOEn1tohMsDdx/D4ob+pL9yJkxY1ix
u6kr90TdtM5FJAVjIl2FTol+s1RinOXZQIglE77vSSUPxItLT3DDlFOFfaHgiZ8N
uKdf//3lX3RDyRcaoWeRTPDuKIv/k4xmkbDzQXWiVKCyYCrqLRdp0G7q0EjuUVAs
GsVhi6XYQcgMmBTyIy3N42LXgWx6n816PIwakpZ0wl14artU3RHxSKVEhZ6kQHGw
lvy6/+Pt7zHnS0uLgkIo+jxRJiU9lCclav3uTvfoe2GvGlMbEcEX5ab33lJx1yJt
7cPFfncxlcIs70UXjhHLHWglxbyfpkaegPqTa6eciQrajWvO0VSFHICjwh3iN41L
xsoaabhIajxbU5Fjq0XpROtv9t0bg4ltMpyt7vD/Op1MQwyjpdIZRqW80fWAlvEG
vrVOLFsbUOqisJNsnJ7orPiHDBOBm63PHnac6k4eM3F7tvJaMbVB6EfkJZ48aVQe
oRDPlOz9rrWmpl7bBGn66lFdyQ0itR+GUdHjS+lknCi1A8Icm724OIVHraVKFQRf
FsaizkvnCTfoqpo2X7NE0iYI7UobrcGqraaLM03/AdLolSMekLIPwt8lYic6/KSR
HRoEgftbrJUfS+b4LICkGIXI3NqUWWaYCxgm0PP5+CdxwP5PXA2ekoKQW/Cjh0wM
YhHSwy4c/M/oST8iN5U23rprTLqZ3Qe0H7Zp8otGD07XMyMFFSJiMjUOWfx9sqKH
vKn3YCM2FFjIuqy6qUGOvC7qrUNPuaChbJZMzq/4/trBzmbS3ZPPkHiLfZnTWvcm
iEJIwS718gyJovdO3n5ZQHuvfjY/GpPRt91z3wcm0OeKWHbZF3IJM8Gs1J+6AXAp
dIq32Uc7meXD9jjTgR/nYfgpU4MId3pSoK6g9ZwSQBakYRWxYYjy5ESUrF0/P4RN
kbPSbZMp/CHsD6073ivFA9BZXvhGnkg3mn/kKgspLvJBbxXn3+IJxBOh3nYYh/Mr
gH4JAob0STT+w/YNCwxmxs4Vokqr6ghfaA24vkVR3lUAcjuHjmypcP1mYA0y3r/w
Fp4Ini757WCn9kGJ/ZyMaMDayNnV1gGhgjkbdxBSLpq0kQ7aFuPDFz+yaxtcownR
sSft+4udp0+RGrs0JILd7xisXbbiRlDRGjsPQnQOi6/zPvYTxNewC5lrtYIKJ6s2
gNPsiliWeflOmrJ89N9v8Mhg+u3ciwxL2uHf6YKJwKLHm13ZrAAJoT9zA0M5xta7
xcBxRH5UUrw0S6uojutaRahHSgoH47lDvLL5DeORfCozfRN1x0F1hcuIv80cp2vk
pV2frU7nnVvzB/L/VpjvKazjYLqSnH4+BDnk/I0U0J2m32y+tDeE9ODvTO8PoviV
euJ+2tHbW8KOMmaFY4E7klk62Tgub2fXqDlCVJhdcC4gNv5FYL4eTzq5AVTj99JE
Do8WeWVhLVlNj+baldSOAMaJhYkuBYCbtWrKbarwUaNDMj6AB+HYB8OMBIa2Qwr6
C0j9InqgTc+RQ3vLdgb7k+2ze9B9jM5AE6epErKodvQSFvnxLegerhyvWBrVi63x
vW5hkiUE523VN+IK7On0gDo9EBK0zemZeVn0fQkSt3eYlIjSbMQVMruj5XQZ+ioX
GnUcDwsPsi2Qxqbgr8ESHWyoZqKz3iTx/NLVoGQc8J+wEKN/TySYZWL5FBEYuSW+
5Ofj5NQlGp5TO/kdZU6xFVtvuA1yvDvga7xKTb4FySh+qmWDBShZiTgP3+wxGno0
wRGQCEZ0WKQEMfGoFJQ/srUu3IVCMmxzfBExVnqGllCjz4K7njh8AsAaZRR7SrKh
7cEfarIa9x4iyQRFu9MWk48RzvYHN8DV9b3oG5vYkBSyTi3qFxdyPDo8r6SIodAi
S7W8SBZpvGcRaoQ2luzY9iP1UmH+vXGRow0NRMYi15kxonaOfNCi0HFjt3zp9Ud3
m2LTHRPq3ElJ2S4985psVcwtOyzPWAjjnOHtdO62ByYEvMNGwl2zL6sPF3mTAkTu
5NqtYlf3Mz9FONtNHugIqffsSh1uEmXeOL1PuhMDO1ux3xD1UWwbwkzkD7aDKJoc
OuW9VZRNKhk8hZ++U01H1pB9UUNTmB02/+rkV15tsCrATBqikcOocweBcxYk12dw
BQG1pkyRixDJlx3FnWipNzDjSWqaJmoRjlKXw87IZ1iwJfo3VOAyOlxKSGypXeI7
2W3d0qBAZYRlCR5QGPRhGETDDNOG3fkyQR85z008eOEscXqdrwP+5GieMstLqSvI
6zb8zA4EehCrRvAKZY1V/maNMAr8z2uAgxpKZI01mpIqVwsXFYCN0mnNld0Sydcn
JShnl3z9qjy6Ct6oHOnoVsEeDOSBvQq5bmqFnLKbwkGfOY27cm8i+v0Ym9b/pXcK
VxtL1Eh7/p8Ze7Ivdn8UEu71ND56KnQclbSbT7G9SWj+yeoUqOLJxaM+u1Z9HWmV
OvnD4W2NCfhZPRsMbAs5Xml9Zefqch2NXgQLgNKwuYFzNaW/XUWsstUw1mbX7+Q+
L57KEwPkWlVBAjsg1wgqU9GTU+Zc9q4a26Jm0mhBew2tHeKFriiKkf9RkzF0i7DB
ryTS7Xh+29+N9MMT7DoaRTzasuqB3rUOvJvMNExeI2HIH2j6S3rfnLRQLd1yBi1p
UkQ6oXO6Ar9K15zSKMdWTKwu8EF1pGwTYfX1a9X/G5p3IY4/iEYjkGtdV5f3K7JL
Sphuk60gTrQuyK6JpRh1xvlHpIJNHQQP1zQFPdt4KX757eTRic9u3oT5tmhRA0EP
BolRU29XjGCpA2xRbJVqGOtgpLaTvfZvZTVysGIaKomFBrIWV8bMpl+9xvbCjI8K
Xlb6cBHD9ahMYbf7FypYvuaIonhTeAh7tuhappRW31RSfqnOS3KpmpHD2GS+jlm6
DhWZlHmEJUl+LTFL4Qw54JitZDZ8u3xn2SJjk9li0AbafmRiZzZYCUyiMjrJ5AUq
1V5ObEE3LgXAMqgyDEB7pw2MIjmailI/88lONrLB2+o8yfceFp9SPAZyjj+YnolL
xPxL2vAqdrJANWTQZLlba6Lxkjf5uqOkQPKp9hA74EcTUdFYc4KncNHIkUrTCGM9
EMxTrJSOWdQunJm27FwXSBoAPPsG6nmayBIJo7hdSkmlGBJx80W9kTF1hPq0+Ltb
+PjcBfSBgKp/EzUmzcUu3PHAbnOdSb2FhQ3lIb1O1MJviP8Q/IiKuGKT1cLTXeLF
Ptk6zaCnomihjVJQyjA6/bJvIlLvOxexNCftfEUn+Ev/icqmDOS92yqcC85Y4jpG
aFwa/pS7/hbroaqD4pGAEPwgI2b8HzbAEH2gzofD1DrTTA8kxHBNLGmksdo5pgwu
ezzkuKVGIs8zBkiu6l7kXN8BSFqGbg+LzmKkdFel6d3Kk+I7rQTR5+mSm//d1p2k
TcE+NQAbh14cQVhyZZuK2raLuM4NQSVEWf8JehJww9f3eeLpCGhSDdGt34Ta9WaA
S5ug56oetA+iSs8+6NxJ+eOIZjo+bgld1jUgEOIeQX/B77ackzZjHkMCyR5rKqF/
kRhx5Tah9EZlc7ebAhE6yyBykgQrhaxVYbn8sViY9VUs1WmApOR/vVnuu3rgJtz+
5sf25yictmmFb1Vg6PxTHRvxn2ZHWb5vZvoApIoNBxga0jYY2w2EYDfmFDUuGnY9
blvMjWZsql9N8pXlTy43YLRXtmXCbEyEHDwqkH0mgicJ6hQXUF2tvpLjkmfD8lQG
oResWckpz9/Hpzg7PbsAZujoaiQoxtO8CBermTwqQ3QpuFi+hz66xgoGsLuDEOCG
MDOfKsf44Gb7Wht30zk4no9pBqjKOWKb98OaB5GTddbshKHgYJ+F14f1M/yKNuMe
QSOp+MX0zzNwHUoKyXxW0E7cVH+ZIFJ1yrGsTVgczAMr9yxyGD45JXkt0/xrXMd4
QzdNzFdF0sA6Ln5WBdc7FA78rrYqr/iLzulXpgh5tgcX3HBsyaJNM2xq/PLM4ZpI
VyW6WFwTAGap2tk0ITqUbrC/glGMUhEy4wSEG/MFD1SG7vdM7f0Eox2np6BNE9GY
Sgkeww7fwha/PfmFfon8dIM+c4GjSgN2EOkWFXLDzymcIUPp+at25NlSmqW/Whmp
Yw2vwXTpRDlC+p/TPzs2Bs19HKddrZwjKGndtU0I2GfMdAlDUnqO9vlTufDU0EB+
QdbMIAdSiFHEnlqHUH42i0oqmVniG4NmktmG0XrYLg7+T46nk1o8CXKfhyp0O1d3
7FDodkAcbkCvCngNk9YlDfC7b2VYGpA5/t1ccLsuX6BkyIJM1aSsSVAV7NVB2qjG
v3bbhhX18Ie80S935FA1WQFxXQmqYO9g6rM3yektVus+EWByglwd4Y0OLwJtNhI3
U6u8RG5lx9bcTF80DXkpDVEJUXVq1/qBFGmgAFEiAwLfSme7KkKxMmyDOx3JQspn
iunNLq1HEUlRgIikXwX1DXuCq8exGcel7fPwzzsu7MJnHeczK/qp6+nIgaGpW9LF
a5RgFHxq5j6FJrjLFlGGND5/J7ujHFuqB5+h0UnoOXEEnGZKfH3rFlM1po9cZxms
gLQgSotN90p7KeZb0tQjpTweYfi00+2jCEwZbZQBKsCwSqmPQ570/K6ncIQw7cKD
eAJjztcOwSWhrRzdMkTXpD0w9Js10DvxzKNvv1ZZzu3lGsg+lLyDZ4A4PHPaFqFJ
dmuoD4N47XBcgfjtYgSGSTBgOc3NlpyCdAMSdhJViehbOApBp5fdpqeA1DlKFTvv
FjfnbpmmSBC+aMz9VowvG+Xv3nen7DlHc4vL/eMqPrNQFyOEBSMUM39i+3CItJop
albLDjgJU6YNkiHcLMhICN3pv7+F//ZTPrKicP55eI/joumbjulnDYmPxHNwOWdv
Y7b0wvkDc7X7DUAc1NAyjn6IAKOHio2ZA1J/pRXxmb9nCoVAJ21tQON1O2r0CzX1
ic5PnPQdkuK6/EI68dGvjY8oGJni8DtY3TxMGZQedYnLh7i43R31M5Wo7rk6bDL3
9VMGPoKGnfr/n3Qpklk9JnGDW7OOU/F8WMj0vgFVMgAFwlKOs9TX8u5b+qXslNrk
opeiloGiwqjOG4e4uqfV50fgACfhn2duaVyB+5MqgGex1cwCgOB4dicagEMbDi+Y
D8+nK+1HAVX4Sljwhk3VmzJKs4Qf9GlaBzT1JmkRKrxvm3qHmK12MdoonTvfSztk
Hn3mzKlbPmHOfq9BqmgjMyEZbHfUHhve9kl2G88IYmGtg8a4nLQZjbdS5mh/RIG2
7xhIGNv89jwrVFtqUido9yluId83hofjhVDWKnUvkizZgjaCEe8TWI3oaFWXhSZT
ucfE2sSw9dXVgeBRrEnexH4PpjIIEBoIzhxUGANtK2Ok2RjHybZ1ijhkhyo1aiOv
yXnPdED5h1FQBV2xcN61oZc41K8wyh5F1Ilx0fmhSK72VIZD6iiPSaDKI1rg7Kmj
IHvHoQ208Ex4o7SNdibDmvAayyJ+m3yWKaCJUyK79kvdXVulpgKU/EgD2o6hKXlR
tuwzyawBnWcN4aJZfqtxntzdUTEaMAZm7hvvCRWvjGjCZLsFmTbj9RwRD4hGDz2S
G5VC5vwLRhyHYe8vClqImOaS+ZGGSWEeSO/JRTBt48L5DwL/xSwoZvL5VaGOYoJL
OmeDv0GHGOXnbIptQqYFrPAmy1UP971Ee3MQnpP07ceO1sZffa1S92F1byQIl4Yk
pAIzvE5QebFUzmUH20aO8lxwQfJoNAnce4OEraAKaDgVTLucgQ0X+eCTv4OuutQt
Kca18X6ZxamdmcHKv1yHw1pfZRaNvjD6JGmlgKL10VfXVc/P0JgCaAw0fDRndTYw
NmdYT9XS5zR496mUkZ0wB9Ang6zdukDKKvmKc3Zzb8URmfPk5bR7PgUdDDjCZIH/
Gqbu9DG+45KTtNs/YviqHWPDOaPQtGkPvTMwhrAPN7yuAiZ5MPEWKK2klXJWO9ju
lnplBj/+Radd9q+DlarhVcln0CECzp4WppDoR4bfrSVKuIUprXjwfmaHZiW3K2jK
6FiFY3frAn84mzkUHiRNIhll1bnMErcoOBkOi2aV45LdVKfheaZ7SMmYy6EMrwHE
b2QmxNB8qxmJPxrQB+jKml+2KFbQEDyloF4X+rNC7olxlC9NkNVhUse/0WU/LNYc
JrN1EJVm7qc0+MBzF1yCnC7XLLThj5gK0l6aLmtC58VLrOHafkZ2gnd/MEb6vKhp
1kHn0tAKwWaqQw9RWgmBaHo6u232cfbmW7YXJ6hrCOwyrM1vQHDP3qHkbaVfcjg4
CrEJRhHDPIUWA+DJnrAilU0oGslCDcmc0Otj0QGuzDKMlud9mVj0oNfMsVzHxO1f
uXSnzy9pZZtO3agcMLsgdn3D2zAh06Acc2E5r1A9PbBbBbW3Fd2aDPYM4/Diw4Sz
5Iof/noNW+wT/A2opT3iqsPTwA36+Paw5jbUOuqei6TOo+GMLYCOuo2cWhHc9QAy
nDON/2rnO2AmmMHEw8h1PsTjw0dgl9QrSiJxlBNzsLHwyXoLHAYKUJiZu/OH8nlV
k4B/50l46kLfKzz/bWTONZVnkQNeGFA5z7LyNUDzOxOZ1q62wfVfqFCXlpAk68+k
bkl+UJBsJ2Y2XM7uIrXR704EZ5iQBIaHpqe9C50MpfgN55yDY3qLhXO9Yq90izHt
YKKtedeflaED2S6rMuOWGhe5bf2hnnszXM3e5sHMTiwtfFQJn+HPAZbwZVt7xtEM
HZ5rwo40SAkIvTQhh0CEdbooJCP0dNkAWI1wcBrigQM3dhlb5HQ3lJL80ru58YI3
2jdPBYfS4CQOIhCVMazKLhp+SS1UDb37EUAZvJW4NlDEgVsd4OfnQwQaH5MAFS7P
wkASlsTBxfvEnYSStsbQYJSDW9SASHtsBHkrURgNU//xu2HlplKrNfAcIF57DXhz
bne7v0n6GXZ8qzgwAx7a9yaw1YURfbRS7c76cdXPvpqGs03kVcvQ0dXTHYVMCWE5
axf3HnvMCcmjEJyVHpoBR5zZcq/icccOxNKxNNFeOOgLL4wnSL3Q/PkJD1yh8x8A
6SIAfUG+ACEM+AUwdyvgv8EjHoMfqqrslELWEdCa90WCrcadZATFEPkoLCjCcmdW
Qrfe0Qv+iytS8bO+gPHVWZw5a02WKI+CvObLXf17GgMmahegHZzRc+s9oKvjJsF4
5uCE+VYiJDDMDCMu7DKTwdf2eJckc8wIct90DW7osBS/8rb+Hj2/12CfiPoebAKB
4DImZnrrYqhcV5A9vCnH8Qb8r63eGQDbfhsOmEE7/h+S7ML2CpR9qQd30lUzmWvK
3WiuE1svMzOcBNNH8ESoagDOVeUb0mkenxXIWbyqDzbgp90+vToyL9IOr6MglQbx
I8XyChedn7DgzQXES+kz4PEJMORp3f4BzpVohYKSQpA9PCTw8LQ1bT5FqxfyZyZ0
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RLd6rM8Kkb1rKUNYB3V+1/dNHXScGmYFDpRnHyP3vxfeSy9Ab+8+a8UaReW8wPB3
TzMbAYRRptdDJ3+1H5DOJP4SHHVKGgU+y2g/m8FctDvzTnfWTIi5mKBaacB2tPWS
uZpFwNY4I/rceX+kna+Sl4frTXmY7NUxdqAdo+/HRtcU57QdoGq918gUxBcQrkJT
c418clIKCcN8I02+Jy8EqAbf2kW+mf426nuCCqUnAxsEz4OXh8LTqaRiQdGj4G+U
X9EJARamgZENhNA3w/W2sT2epQDyQXOagZQrFw0/ohaw6sPFUWuM//w5iZIGKSUk
LPg2w5taYfoHtdFjZKFPFg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1232 )
`pragma protect data_block
KTD6+Vx62Z8in3sQVCyKsvRcPjF1l3N82dgZg73s8ZxJUCGsZY//Vigqr/+wQcva
ekACAAtqkqt6zzYtbzpbusdfu293YCnmzqoTE643xaXzQ85Q6oLECZVuNQ4BbKGW
rAKl2ph9I32hWbnzz7k5YE8sh8Q/7SkAprGjW/in/WdYF+GzxEY8si6if1t5qCX0
nV2coBd2tx9NVgdatteWUXaImvYKkCACFMWE2ZTFJXNlxjpsJ5waQlk3OM3cjHan
74Yi5xfm57HbCuVGMJwtr0x1P5UTU8vksqPCFVY53P7jWCKdtMby82wA8B3ewZEW
gUuwAXHSdMhKYP1Vqa4uNWUf5sjCQmsz7xhsm+0Jlf46RKmmadFPJt/UnNT7st3l
oNmRXorm4S96sKnbfRpTK7OqvkcG8Vl7jXMuD/SoHWutIfg80kaRyM3PjI+L++ri
RvtEbhhotSjN2DP5x6PFpACC0QUOpmry42Ce4ZyZcJ4A/pdR0FRO/h0Kz8/w1Bqw
jFo8Zo9+NTH/Iz+UNBco1dUEx/Q7kAKo7cTuXD8enPQG2M+Yf3/SeNlqyvYCLY1o
xOI/7agr4ZVWwRKncEPcWUlrjnU3DudGngNbB5TyNsM0sn/GIPPfBRgMv5yetGxM
VgghcRgkw8DhKx/agrWMjCasBYgawtB9ngPgeUl56qbXkRV5sHePOMXOUzbTW6Au
b6yxFQ9gqCwQ3aMDcBXNbmHzyjSePPGe2xDNAgnxqRH1KwZPfp6G2Bohp/3npaqj
+9cB48XKe8CCv6m4Rak8DMtmdDhIDPEt2sNHdABj51dr2dBj5B8cqmUMJRrfPfNL
C6RWJwZ3gEYIJxHeOA30HUapsHb1ZQq1MTyKjatNmNC61FXUzYAcf61WT0Pkqr03
QBvblSx7SSvtYYvXjmiWgSU6MncNo3WELXGbIuoKRcLkVhs52mzdE25+D//D9DYK
duL3IQ9un9YFdNuup1pEqEDXdeZkm1cRzgJLLaHGQ79nN63KU572hEkPOmelK++S
RWikh4TDKYGB+XmuxjK8CYyjtXXWXIU8t8KH+OU2TBedrPGnDcfXjyMhsholqLTg
2017wtuGTYjvoaaQfwKVO9ZW6BjXgU9OfvPCe6X33kYzPwGXUOvDvV1bcBE9Jwg7
PZzngQ7x35mJjajtuTOFS1hWAgC/2vE9mq76rgfsfIIXeZ6zPcFlQt1ZC5c/q5n8
b+8cUGSmKNtq1nYILfqzSeGa0oF78sY5FtzE+mYx5it/TCZ6otqcHuCoxO/W+4BA
mj18OCpL5A0s7L4RCZeovr6dRQC65mJkesfTHN3tQCSO8TWJs7gel+rcYEFfLTGo
UGkf/k0P1+9BzzjzYZGMDr3pGq8AcDTHKeURNxXBtJIlpGdSewpBw5xRwngt/xWS
J11x3mzIxxhGnfsFRYAbzGVslHQvkB9lqA5L4NLiquKmGaur8CLvm2Xb1bRrK/4z
FvSJtzb6CRHiTVnqSJQmte8JBrqoO+E5M5PVPJMR3gtJHg7IwtYzseZv2huSVXnB
E6wgtZ5zPFEqv5rwIEQR6wbWtUD89gtbdLien+y5q8jha00qb2b3ZeNic/ufdLKc
3l8GpWJ3hQMpx9k4KvWxaginYysyLdY5TOiHsD0VcGY=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
QumKnJGGWzIONFin3wXznrueeNe0gdGx2tM0ncJs8eN/jBO+V518ffg6bNIEa5HY
ekIu44MyvBYxUXSK6N9kcB8J+b/67LHkO+rgunL8vPV5PZAW2oiJvzq6eKoWZJ3S
/fdVmXRbaglU4jPBvno7ukxlMgQJCwg5vegzqHErjykXu3Onx0rD0DqN4h9cym2v
DcSEZ+67Oy5sTg6f0cG1yuQcvWI2NrdkJXtQuZpK6amkbgdCMVxwG70UD1WqJF5v
cBP050cCCrUjXv6M/qe9QXVMaMHVOd4qcs4/EdJO0zBUkAjYlpp4RpjjTbkIi+xg
mCrd46as1z77i2SLqKF5tQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 12144 )
`pragma protect data_block
m8gVLBvJdVDy+HFponqiz2uQXzLp8CigexTVNPSHJguwlE+0b3+q2uaNF7SrMHCv
+lgtUvQkjYFZd/yELsAed25q/1H9DyMa1pTboLDV39XjAQJ07sk1ERzoz34ZExn9
ed3JhZVEeTrJ+S0Chi67VJAdYlx8PiFQJoYy5a7+4QHz895/CinYugp4755Mleyj
NepKYe6gEsRWNpZsOyJfcDHDAMDYfG1V0kTM1dh7GDl2kIkHZCEqKemOAOJKjABy
fjIUDpqoabqdizI8ZPrrZckQeTq1jQOsxgDkgZduWZxdE9eUaTnTYl9NkqHS+pit
uHtiPTa/g7AS2jOAUpo6Yrwz6+pCe+sVHBpEvxIixpkXV1KwQBVSNCNylnCn+mPC
tNjvDwSAOrFYVQ3y84gMOPyUB8uubCWnEAcbAXcz+5A1qvhoge+3MNSg2EkmYpIt
/+h9k8jlh6C5eGEhvvYxjbP5K1g6jLfbw3GQRq0n/Sb5M6LnvvajbjBzSyUGEKQu
pyQZ09bmJQD6ip8saxyrGnUjF2Wm4ULLfNq5u84SgncGz4ASgGliL6mKBr5FE07S
VIfw6vQCZODmIJkzKSemWiXM5+epSYtIgTb9uRr5LrjDRC+56n1D86sPKDUy3AC8
MmWNosGbGQSGpsZVhO4M95g9dTPHaMx5+BiaeieqQl2iJUfKYqOqYCDadqPR55g2
QZ0O+0rNmKqqujKxZp4wKkxfdcHxnlYT6Scdopyy1CBiHBNWl3ZBWLqekd/MzxhM
EI6M4UsY9E/dnSed4KLBQnOX6FMLlPVk0Mmby9g1neoXt0RTJTt2b/W0PHGyOdxN
08Yvkv1s9riB5MhKuYgK1P2c+lT9v4UMeqPqGMlVbFd1jIrGbQoN34Tsr71Ard7T
KfF7Y0XpFzo1PIZ+8DfGYn5iMyLvhAZrT/oCZzQftxGU5G56lv578MEqbuW8UiCK
labUO26DLLDT0dDhO480UC/mdASlcmulVWTX/bYmzRT23TA4BbksvzSG+lMfjHpJ
E2rc+Jh8zPe7X/AnuJ2HqOwp32JYX+1s3T/CnmztQEJ6e6v2iyRNDubNlSBE2qac
vC8R3Y1rdQ1MI+zN159Hpg8V2iLDCxTEWPchHbAQerOFFGwEcJqv51MrXwnIAtsh
BOhoPy/afVxchgs/CDQIhvfxQFyXNto3JoTXncdH5Rhx6PI3P0muPA4Xsw472Wgk
aP0VKDBmABICcrr9dpRtFT1UZEJNxqNqmf1yfRFEFazRGPsoGxB+15vqV87LeEcT
wB1oJUOPDVY0/N5rUASqrrilfmlRGk2/aIpEnqAwl7IU8jefg9BWk247c42r82sR
WAJi/cngRIWWHRwnV+Ch57+49zsUc2tyB7yLJ1J6PFHcEDzMWvyUEtZuuRJUlGf2
xG/z05BJtW3G/VF91sF41xV64hmlvHqXSOkkINw2Ds6h8CgieA9ScfXwjge6EZfD
FjamQcMqU+oXs608dyzEhgX2a/9X0m+ILfHK0hoLgO6S0XGRjDfiLsgGiCPg0fxo
7z3C94yCDxBHL3loGRx9DSux+JocqwYs5aiWiTurZiZ+e9OU4LgxUnjTt4ThZ0LL
p9/t2P/yWn0LNQ2TMMPni2uw7tJRlitqB5ETgInwDO0SqB8sVVJgk2wf6PMSaq6u
4aQrUcLlzAweYIgG66nSeNy8N6s5rpS1JLQ5aCVVVFO+I+VgMuy3D8mV+6Sb2FQ/
1R3c8ik9z3WYXsB8cBu7LG754AVA40+vTK4wmJYupq/n9G58RybQW9ifkdBvnKOF
MvBUTmk4d4Qvj43KmG9U/bzm2tteZSzaYnQAt1Mw9TVDCcmlLu3JlnDhOJbrdHj4
6kI+QFxfwzyxwyP7Oj0subud03iypERXRzqb4zBV+iQVJc2s03H+XTEfDysc53Ro
Q9ycF6FiOFIvINqcCfNehfgiPEpR55hq4SU25jFLurdntYXroPnl/Lt6p1CCdxNR
fRXKoJUo9vWXfk44WEC25IByR1aJHHEWmbAAKNHe/ITW5St15d79i9GO4230OR04
yRDPvURYxyu9UIjahTyVWa8U1P/+dPMmje+hgB4AZkkEeqcjPStgANQMkl4kPcZD
LV+7LKRNZCjdZBcuG2rCN/f8PRt1Ve8h5nhP2pbyFhciVsigQsR1307DeqBesq0V
xkswHAZYNLnZ6HPblhj9AOogFEK2mxBT5Ed17Ogknfjbv+YpCrGDpjuxjjF9ZllJ
UWDjEzcIZH/shzLj+yhBgFIMFoXDs7hgZ5FIulysfvbfhJu/boO3Adi5DNcjlnAl
SaO26BM527x7CIwlRfWCJ9IUZs7EWnAsskicHwYQo/V4ydr/za9CDgjhBDiPiz3s
EbDwjTvALRTjzPagq+IZxUOsmmdglQoAWuwwO0AN/7J0pUNKaaMY9f0klM1O9TVe
WChsWYzstK8h8HNbhEi8EsHH4RB5cia8m10SDKLPSib3SleSxsJX2Scjr81ZNQha
o/3PbA3O+4JZNYcFOtgHVb7AnZlomv1msw6hn5aOGc8afv42dXNv5fWw2ZN7A+5P
XZZ/f7laIXITzB1qIqRSLZNFagIGXmqB3Q6t6ClYO+wMlBSUZ2qylzt4MFF/xmQA
ksRIOwBPG+7lXtUZ/Sk8oJwXuSP/ohXwZbTJgp0WBW7KoAiNOqnOw+aNqQ1X3/w2
i/W20eLivBEUN+KEchnVfuLEB+F1V1/oz6D4UWnsoAtjBoCstF0LxQfZ/5yNsWhT
HXzIXePknJmYI7yVpKhtWnLx+wbtbJf1y+p9EkteCCM6JuMYqO+I+H3EU0fqZo8B
zjBXOv3CHCUPAr0c3N6AAHyU1XKs8vLABSu+Ops+3ZJSx5W4dNl4BWuDWDrcK+nX
4+nJaMYfW1HqaAeyynOiarE3k4PHz8raJCk4B9j8URX6eR4zgI74LPNEiyBS8W/O
WHidP4719aDSycPlMcJaPqkFAx2VrJEJWi4pm8CwwiB4WEWwdisjeq9xLM4DevG8
o+njCe0JOIWgqCp6AaNpN6hClOtQg1aNyoYCWSLISxwGN4tFM6Q0N4lWhhqTE99g
PAboXkli9QBwIKQdj52F2IwbuYmnwFmfOj00LT6QJ+YnYtt6kZ88PngQ1t2Uko50
YS5VVU9w8YudJtMzFYnjKwexwFYpZgK0AGhqKVHBHB0KK2zv5YwoWzGND98IIS7f
RVFsuPxm+1ZZ186Z/YzVpDgmVW+D+liofdkcDjY0W4e+JmEirRS+mDVMtIpefKoP
VWha0pjDco271kYgjfzh9dTEjZW3OUqZUeceeNOuV91wojbzMHWM/BnijJutWAty
utv1JIiUBh/gZGNwoA9uAifDVKTiTYHvYNKcIOUjCZCxcPuJwS/CGSpTIM4Cnuht
Z9idH+iYOiTQgNBbjYGYKKJA9m5OkwyALYn4DMutSdsOPYSyq3xDPuogqYfBtVCH
60GNoYNmAbVaA8LshEUzNx1pDn4u/sfS0xfDmWBx0pSSS5uJnZflcqFhaoVD6dW/
f1Q/Vgbc522OEw1vPVz762JT7yf+z10UyHaPE6o+JHzWF/MCVUxnLxuwNXGHkKJg
LidmI30dhBtK9gjpz5G2HBfOZ5wkKfQPFVU/Hl/FQ90PMa0BUuw+jw/z1UE+7TG2
9IVC4WCxCn+XLsmz51cxVlNyVduiIcQPS1xmi77abbGkdyy45CFYpXI9UDFDnQtY
c6W2UXe0DW7owZ45FlU99S8yy+e2qdcwmg9xNMMd3K8aHWlMMnx/tSgHe3k6QtA1
iHVHAhVWw4Yhm3adcvUZYQdM19d4JBkkZ9Wnf/NTVddW/hzmIdZOw/7f0DrRKQze
zeQQDkbrsD1+/mjcatMGdm4ldn17KjQ44tkK0ylCDZgrXA6ZHj4fqvsN7/khVPUD
rT1Vzjzr/jeDSyOv1i6LFfBdXkeF6hcwuX3tf+87/DB/QhNIVF97MpPg9b8gzEm7
sWOL1a1/ck5cuskHiq3oDiJlvKcOtLgzN7vC5jG5wbPQZAkvR/ZFaARv1lmY+3oL
VJuZfYWUrtvA1u8qlQ9WSPpaZ5SmD6kFXAq8nBwm0YdST/iGFYfWIGLD4FyahFyD
IDJSx+s7zlHzl51Bzpisv4bsVocop9POzYV0qEj/w+WIBQ0p/cnrEhLhqd4DlvGa
SveKxYOxYuyQ/SYGO5SzYVTb3YbC2v/WUd1CBmoHt/ytfKw+psDKaD/E9ER+E1Ln
JtrqINtmPuA9lKIWCzT3f07OgIgBhLrm5pK/wmMnDfeDCMUwstwnjszlZePbIFt4
tyP5/tKlabD3ZyOHukaEaHDC9lfi8KIStrh1phJeLORbrtqyiYnUuN01AXM1weDg
iJlrNrNGVWwxFBI/EqyY0gr/YS8euCT2KXqJsKfurv8xHvvE4IBh3eXRERNPSxZb
gVgddygwI7b74SQdZqBpXUMlfyiTnt+jUxGch5RkrPACkGR4pfSLkJGhew9zHZpb
hX4kJ+xcvlclmpglu7Dq6KLlF2wtuJcOtiA2jwPOsxnnDESTZrPSE1cAsFQNbSp1
mEEnPNozfrq98JDFMGHVwcy3PNEPcgWYLZQYQrmOrDw4LXjL5eAf8jr/QeACHsqF
QYWE84DR35tjPOKC5/KZM2BohKgNwC0l4kxCi8Mk0s3EYsTGFpnIWN0rX/il1wgS
0dHp1eLW8+KIvfqGjHTRwz3I3JenG4knnMCmfJWTubq+5q32QYdOJXiKEyZshaFD
fLvFjDbsumBK8bS/S8FvnJxcTNbCwEywhxC7O+Drnl9iZe0dto+QBkqaEaSZAc6B
yqGDiy4bwuk7pfSopXiH8BE86E/+3DIxOKrUuA1+FdqTi+sXCLdr1UmGXgCXrNZq
b/FOYg1NAIGJxhTnTONLAjZP9jerWJXbxJjWAFrMkyAJxgVXcurhFjp7sa7OjJW7
fiSZtRgsO0X1xLEONrL5CpVrchv2ohU1pN3BkaZJffRGzS+glQOQ92TQdoTklrSX
oGygsBKldVbnjjDrA/EclZ9N4qFFQTt/+vWz2iPfs4lVKzevKRH13KVzURlN+gP0
A6SvycoybEGnEDN57TZoXb5S7blDaxl5pRUYYogxr2VAKEtkqINRJL1XqDncr3eM
NBOkNj4wfeZvyaLyl6g8j3EuOZdXVCy/eWYlmctRbmuGW+qVF7piIkiG+z8PDH9H
/J5mMCN2K2ZaUiZrHhUe8nHrvhw2NdYzoNlTyG3LcZX3CcucdI6llyUovqtFK6DB
qJXX0Ma0FogOZClT7Kqh4/eYgNRwZ/WDJKhkLU11+nsHsQKCxWUFtvHYCEY4vG8y
L2ya7WWhwFOuQb1UWHLeLRZVzi6kUQfnY1xDjax2a0Ko1oLGHWFB6d2UFzdEVxek
giCFu5fRtcv0ZKvsKm8zfJJ+2j27GlbEBy+wKRnpwW7wcuNuK+zdENo523ZnNhKr
vypVUcP2pVIvxMehpCub9pYTgL2x4JJBf3DI16qL01XiqR2UhPvCOaJSlSrDVe9t
Hzw/YwyDo3nbHsA8EGnvs6OAVi2KRw9Ia9qltPPGbA/2OZYsgAtPJlB8DSrnPZ7m
Mb4CMAICNwN5D1MyX2+R+0evdqHvU2X+z1fllo/fSNAjINJM2JKbaYaDsHVYJZMM
wq/0/WpA8KJC1qT6srRfvjnxCx7fCln+UuvdaeafA2SGdEsbrBDLPwT2rbFp3+JB
VZVzhexxPJDHRi31rAwN9yv52AIJ2QeL4eZN2b0LR7YAxzHfXsjlkJLXDiLwQEf2
vTAnmYU+4EogCHzowIXX9o90UG2mpVveCBHxPJ9aVjAItIa+W16QV0Lm0qaHe2kE
tlF4guw76H8p9/9s5rkWC4gOSOsgLEeFxemtk0fy0471GbbWcYt5Z/8kMjAB7D2J
cJtPaU8nfSvdiSdfS/q/SOdSZ0HgVSxRQvlfJyUXxqyb9XLFavfBy/DTeapCg5MY
+xNzZNLXgdw+K2K+L9UYXHZcDV6/367CbWYCia2bGsWUJy9Rs/93DGqc6jufOUQg
BpeZEl4uyx7jUKnoFwIjIfxSkE+2WmC8iKovuTdkeJumN4VQsSMlWnwnVOpRm1CZ
ntIXf1fVWr0rtJ4nPLc7OlJj8juMUCNb+IeRHIXnPHL0nmUPOLU6SJbq3LlgfSEc
ONWN+lC8HMos755MVxNJqSblTn2wpaH3vi7trhyZ2IEfRr70NRwlNnpjZffC6v6v
xvZyYYOhGfLcO3M2f8MpQqwBYC4ILA9RwILi2UNkoA+T8Vi2UwpCxDQhLk3WsW9/
/DkDjn5dx+n3B/DgIQ/ZSpxeLVKxfOg5V58+smBil1Ufq2id8Mbx64ClxxiVSmRg
patS8q3EEnzYMzwskB8Otr5qX3qy9iKjmaIFV/O7jd9jSP1PVh/rC4kfjydGxZXt
1J1CGCfzeuQu+cJ7qbh6sZcf4+RA0frwoKhCTSJ64W2HuPnUfBEOH+cyzmWZ3frA
eFw/yBsxefYvtxAzxCDp4Gwe2Qti3JXIGhVzAo33z456GMWvY/qnzMzCSMlM8GeF
d/+KP7inNAFC0dbJy+jNAj8ASMVWBTeCyhtI3zwRV/qqRLJ2/e1sJmWK+SQLO+yZ
fl/8+BQBF4Kxdm5SdVkZIOhEA02+sCYiUdu/axLpGAYRQhhEeoDxjuA78DJBIm+T
UEw+4PWTFjWK3iG+fihfXqT9ehTky6ebTnwRwtQzImyeZWeen+Hqcf1/gtwgR4be
vIIDVtg7RtrHv286LRYEP0k+YFHHFOlNQWssTZ8XCmywJ0NLAcedtFNvOry5VVKB
Fft7ibKaDNnaCsA2yYILBdLOV7zq78rLIqP2BCOkuhy3nfFZKaXKZAB2aAKwXMTX
qmo/OWza1b9HCKo42L3ySEQSr2HogylMGwLMra6H4nR050YM09omAtHfCOp7eoVJ
t7rlmIb837aXWldA/rLsKL5cP+MPZVnCKiEa7lz38RLQBD/W+KD2i+j925I+LdNG
B24mjNzgd4Jh4v915xBcyGqJsmeVjWIc8stxL0Y3Bbh0HW+jae/DkdmrZQScs0vh
6EA8FjaRLjMRzzYqNWXRwsnouQs7oDP+iqixeUx0Xpi7YMTm1ve2cTjnygpgCetD
XyLEMJjAqncMBSF8HJ/0W9ByOX4pqJiDPgZwKgWoFcIf1MkHaFV7bisg7o6TPPCJ
arsEhwa6hL0vaAd2A0t3FJWTK9VGCuXxQza9x7CYYzajbiswhaGPKtUCnGdVLdyb
W2O5I38kghrwxGSik+xebpO+i+WY3/PJH38yOhehzphNtDry1V1QM0gaNg02mfy9
ZeWs1yT/l7UQx9bjlGhpfu+Z3ldLPIkOBYGYFQCkvoXfkXh+zL0dOnttXa95kckR
IBOvF/0Okhql9VVRoAt9B3pi6CU6bdjw6JFo8m/kgHNL+JOtBNiKR45rO7xYekzw
a+rtLXUQd2K++/A1PZxgfxePJGKx90O5nTBlRCrcwSdZ/oE/rOj8nZ4yoUTi1AR3
h7iX9THq+FPBAX+qn8NZaaHXecoSizszDckHbOSRyzb19k6HFE7akkT4TRa2ZA1X
sd1EGt+KFjIbxP5HFYUo9Vmj7NY2tK6uBykAZphgzpvx3lyFueptZHUx1NUv9HIZ
pTso5PnUylTwj7DrJrUrn/DN2xRjIOdNEF7PiljpBGBdP/5MZZcyJoCyKt/JyUVJ
vyctcGhzz55emd5UMrKUfpPHqgpHpMCvNkH58jRXvHQEGiF9raXkX+XEuTgOObU5
qdX+6jzH6YJBTRL47DG3tFdccgb4fy+vuuxSBUV/kh4EkYpQkhfqUwpFeJtx1ZJL
eNqJ9QMo6vJ7Eqs6L+84mLEo39AkqwxAtK/ftSDzEESARTJYfe+Fyn10aTl4WTuG
aRhJ+UBk2L2x/EubttbwSANpIMuiKpkhnXpNuSEo2v2YByFYRnZdJ0ZIQuOK7kcW
cBoeifxqpnoGXpEj4ItoXeo1gU0Ay5jaIEnXv9aAQhP75+GBjKohLqFTCuAyQgwU
6ia3TTANRF14zD4JBkJ26wAUAZ6d+68UV/6JDq6HJS5Xf/zle3ZO87f1rNN6lWiX
KYwvwKRt352oed6a8Y1nEi2N+cXMI35zhLsN/aLks+4Qy8w25NZHlo5vagbW3ivX
FNGICd2Fq8/CaNINRzNq56rRqMkJevdNum8AIVONBYR1ujc9F2vVeaTepqmTUEpL
dEWxgR1hO8nc/cwQcFibzIVj9IetHBBYMYDG5RKiw8/oHuMrgrX4TT1d17CgPFpk
kEoTQCOWhvH9cSmG7doIZYE+XqeYmrtNv6QczQbZdkHuYJj4X7CREnJ+OpEMqtef
pM1vhntjTyRaQ/S+xxftr0DY1zQK0C4hgR/QWumHhPGM1hgOHsMuHNVluyZod01+
drAd7Tdzv0h++NMu6lNeB4vr4rGZ4wYXbYN2zJr3bV4lCy3HR2cOnT3SPElTh9tu
Ym+Dwa5suAGYMxZGwJyJwCcIi+HsUg3b9R2ZAvs4NS0wE95WGJjcCxpBDobtaeXK
vMhzRme9PR4fkI0QhUoXMoMi3B7LtSBYnhj1nWzSOHWyVazkKa/LSaEZxidHrGnT
OETvljmxbBFmrguRmrLCLhdg8cwqmOC9/WjJyeqZdaxlGaA8tdU8dZZjPgfajnjU
L50H/QeCjy+INUfiZdbCb0KrmcAqbnkjtk8wEZQpiKUjNiuAxJrfTRFpp+YPClhs
h8bIbLeGhxave2rnIhA99m26vnUG+vVlaZ76yGy0SRS1NzKIPW6phTNMJ8lJWNJ5
0YEpn0KGFPceKk/LgQjkNQKOQHs1TbXLi9AMZ7C/aS7p2ez3dO8XUbfPEIJ3Fx1N
1hSedRf2/aPD7/ahG5viClfKkYmYy2oC/gJg0ivj04BYi9RgXhmvvihDAtEpQ347
6y4o4yHM7d4mIZixXbTE2RbyaSoYRmREyxlZu5pNoFw0xmNTpEu5XqbIyl4piyYm
BiaafuF0EhSdYoDFeB4zbJt3gHu+XEuYREY0oJENHPQRUO8cSkaKPvrufr5//bZa
58leEoY7JSI+XwnwjEN+L8vd0AtP1eN8ziwv5XX+M3t+rpPs6ZuyWkhr5DuMDKU/
n7A6dmbdqkD/cICGzyOv72txQFT6fEyC9aqjrj0R3h9xbzSJIP/0qHvJ416zDULc
hAwXmmP4fIogzD1YZq03v3nNrx5/rjMusOMfiM4u/l4XsFD+wKpDg2m/BQUPozud
k1Io9lcX3Do4bMLRQFS7D0fe3XRXUylYPNYrv+uXKw2u/Z73rtuYwARHTeaOGYqs
QRLzyV+NSRQgQrQSu0fIJQv7NzIKHFrUq8Y2PRV8Hc0wzLue7xh0d89mKt6Rife6
4hnKWQ0YqZBxTrf0UnRhEeLOnep32SJpUxxbvZGKPiUEtVOj/aBhc9W/LmUliotS
D2QMvc6/mooOYCtSXKiRr84DBoNMiJS6smkqB5M6+Yq1aHUQtBikRilrh+vcmF+x
46icF+hq6CSGdd9IlC5dd/lEw4dEj1EN/vhg+p11K+azU92DuoOh/o1ZDsyD/4FK
jhj6LAQD/ajLaQaZMxWpCWh7lViNQB2EOt3L/66tUMwKsAKHTbRcUJIIrlSUWZnf
+rptcOx5H/79j5MTdwZsueeu6qq49o7EwUklBf7agHHr+T5n9iit/26zd9e7gGb9
kfU0mp1INjTMq7oQCs8C+1yuv0AklUflJYDrqX3Q/8DH2NWAG9LkNEmCFM1Va7D0
h7jaNfjvmsZD6lKwCK0J4WC7rFzJP/zt1uj+o7rMYanQZhiLEpoc+t7Y6xUAR3pC
74canHsPOx7ffGyuRqaf4qjAFCXXy9mNy6rwNoteMDqVri4F3EcJ94lQ0hbccMio
jea8fWHoPuibtgrKGb+T4SuZGxCOigqnBNkLQZlLDwgIR6jO2ERJ/PtX7fMo3jRV
jbzNp6iFOGPg8aBxnS2dVt2mOtu8Aa3UMSYxzscBgY63ukOiOyG0jmTyK1vS+/UN
oyk6f1kBuegqDT6mWfp/FeoyXNTHziEqG02kyCfgxjft8Y0WBKZ2AyhAO+Pwz98s
7JYLsDSyf5Ee8yAHxVSu+HkaElqBlljRY0O2tqaFtxTMnP4o6vrNKKWqBd86UJ3K
/8Pf5ALONH1qIJI+134a20RugLCOiS1c0fr31hZACgePOoZd76WHAilx02MNBGVm
8VW+E1nS1hxr9MiX8mAMaKeUF9X4VxhbF5BM4ufJQmJIN8BaFLXZAKosipkegIv1
dHfdXv6iJZExEjL2Fov8w+wNRqsnFR7i7cAH1+AII5PzqYWW/f+ab+C89xpTqvbI
jvRWyEgBICB7vuNtye2G8Smr6PgP4UUWj8MsRFZU3FlSSs4Up1RXmj212sYXGknZ
3ocqLGk/1J3a6VIIde+yeR0p+E2qTfj4QXKP+lbmfN5wmKnK0pKRkxeW60NemUe0
HCrdUK6z+wbqyKBy3tI5wNcIPwmFofWMXDelitKSRbxvjMxYxmyRXxHNVJmD9E0p
SKIhHrEof93fcE0kiXodkfvUzQvgQmzt2ESfC1u+QsnY6BRd83pGloGmt/UcmAOe
NulAev6cHvr4undPUXSVF7uRy5glfcO9oKRZ7LcMr4Y1LvQ8iPKPeFAJfKvhPcuT
x41hso/cm4NaNb0CuZDi/chXxYwolbTK8Bjka40VBp49ykhCFnNrzmxv4cgJUjn1
MFTSLgi8BsKX2KHTxfHQ/O3iAqkWKLXh/Ko+EqHZ/3ln54KbaSiQBbZdy5WXKrIv
qMsI/JbBthat1DPHieEnA/Me6t2fBCsEZs7nNuowFH9s+qtNqkebF9tL5at0RqGV
IIjQqNsdhO4xDiBtRn7pq5QMvuudmU3AThn3PfeEZ6or/7WciuqkCb7Ln03hwVDy
/bwiOaJCGeLzdkmVcuz8yE3ORTdWEFNgMCAT4fZ/FjhrYrBa+ApgMKInslQk1vk/
j7SrPfiZa6JO9zhR3P3nFpJri4efYYbAqrmKCluns+j3lWfKIW3H26QVE8UgLn6o
vSQDiroeV9RWTYmJziLJesfAKuET3+iJGZJ3vh+Fn+Fsp3mM7FmKNYjdTJdlAeEf
pp0Xq/dqFTUZ54WptIWCLyCdGG4L/4ZpOci0RPBGUa4mNM3A3x7CZ1jp51ozh3gB
IPWlWNvQcfLmru+UKsCRWsysBk9VKj6eFTgjEHpLNMb+yNxuFVd7cX345thm9AhU
vR7Pv9bDF4f6+bWf/gmOOLSHXFIHh8md6PLsRqAf149tWCR2Cd1uJKfU4q+7IS4d
C2Ss8n9BNCGvKJCe50n5/ZDZ2RhNOHqV4pZ3qS7oERgqN9xpzRUviOD7Km7bOjmA
pQQB9voGHdXNwx8w1zOq09JX1+hQ0lxOMP/A2FU1LOU/9pY+QmG2MOZPAVfZuWTX
0aXj8WWKwWnI2l+eakd1Kmm9H3vrK8kUWNYAk7X42TnF/E3oGfrQpAm79y7lNCp6
lfHSLHYXWxI7RIhPCcOXmuD6j3xyJCceTf/rsfiOb/R+tZbf7ExBSosUivwe6jdi
5CbBPWUCtRscCE8x5TCsovKX972JxDpZH7zc86lqXOuopuihPHKlx0HuM6FS38wQ
gG4O6SMkeyMmVb62PR7xr2yeyeyDkLTv13WPWWZBupSrPv7/UQEOiom6nUMTeMx6
3rZVLsRuwnzCGTJS+Ugfp+MHU1XEvusb5J/VPiD4DFJU89SMn3KQI1n2YImXVsdO
X+5E+nz9aycs3P4tQBgY41uPONleFvRQNyvEYv06Rq/sA+mI7mva+zBYRpHdbsUY
cjrJcxQe5nrqO4vnNReIHAxIXC41ljEKvm1M1ZLILOtfxfTgtZSsIybhR8xkgNSV
RO+S5cAFyPNl+ZI28Iu/yDNDihBrjKhqI23vBaWApLCBHswpXV1urYtXwUho9VAQ
uOZZ4Bm8yIh+SUKdn0iYWCdLukibbUGaKmguPKpcx2l7c5qTJCc6gwNSjJ2ANY6I
kE8v3jwfDrdTAoOgcH81+utb+mubWTnjRByN4rrirMIAM1dZfeIxRL127Olt5riF
/pEzAElGPAuhzDzXX6WKpMpcbKS2SglKEs09126GMLJtfaFbgi0J9IqLuKsvz6CU
egBWBkiMtP+2JWy0KEfrVYPZdqJ4ebt3MZn7DZA4lAvVN40pG6n1mbDgZj4k0YYI
f27+RqumbzP857/N3vql8KrPugInS/8uMdXUp4Gg2ICzXZvOxX+vqYkNxLZNmJn1
4R5WK6FHn9Au03WdAOGzlWer130TiLKvPovC/W978+BLNm3RIazJQsA1U8nke+rk
WJuXGHyjVACbwBTmROaFhWT6qWE4a4F83fXj6oYSQfU0wx7RBebZqTnK58Q4896E
C3PCPlUd4I+iNanBgR2wcQcg7YKjS3pV4ITlQI78DAnYAvVQjHyCkskKpdx04MRu
IcTppzUFWOze3bO1MZSlf5PB0ftYrRfK3pgjgHrhWPeN7klUoBZC5cPWda0a9xNK
RH8pNYD3YwbjzaeFiT+X22bC1MDaW2gwLuMyDSZRqzja6Yts6CkaQzZPzJUCc1EF
I8OfzlUubdPZ4kdzKOwp1nSeTmdLNbHeGX8te7jCBfeJiqqtiOmVgAroEA74ta+L
NGodtTlim4k3+dgMCCXnzfuxfXK2fcVZ/4rplmlzOsKTv4e+GMYpSMlNZdGI7oq3
Qb+mpHNUdvyglzyjWkt3U/upJ/duhDXEdp4LiD+3KnJbi9gfVdpwUbs4BVluxy5o
9i7aDxWK9cPXBCALkDX/RGIox7IGtWvm6mmTXkS1bieKkmWTGuaPBpVGyn7SP876
LooDIxS2mJfrYcypYlx9L8tV+3Mr7A7LS5a0gS99ohzfTv+ThbwiX9BvZxszjPxJ
g87NzFn+1ZcqQUkZ5a87bd8q2O2MF/OVu5Xim7oRyc6Ej605NVfXEV21chebqJUD
XaCqoanR6zlZZBrnwjxhmJIF/zbTRZImBl1NTQgkp7GptRZlfsopzGxKZ0+hmtqK
mQN98O3O+hseioNCjsokPujga9pFgK2d27OmI2XP7ht5my6O3UNF5Z7vQhh+GGub
S8dckv1LcNBW2F72fOLN2h6pF3rn5TNyArmScPC3HkHWkhUOzMkd8IoH+jihMWdO
R3p44BGMd3izjKbrHjJjtNeSgLpNRSVRcbYWykpsbBddvICOSoLkjDOpqjf+Al4u
8O9b+cTkOHtTFgxq/3AURW/hVW+Jt6ihnqz+xpmTTTBgmTT5X+qlKrXOEy63bu3F
te5sq/koc1horAxfu1ErTKy/39tBdpLm3gWrhaB+0iapAifSQZWDUVrWUvTj42Ik
3gSNGqpZJO55h3WkK7fiJaUR1Yy9ZO1B9cPIguRznxKY04fdkIiLgiguQsJioNGq
aV2EkUKaqkQkeLealPoPytyNRcL6wlWmS2M4Zag2EdpSD4wLLghvVwvSm9XlcXgQ
wEJraeWuxrOr/YOeHNGPnm8r8G2Ta/nNWTz7KaNTsowFfNlouSMGLhtop39eEGx3
WIH52Y4O+PgtROGxAsfzZ7dmykWPXxO9NLS6HhJpmS+aLeQsT/+qhaQeHNvLRaId
AfDZthiFboy93T969edWAER/JhRoXtpIo439oMS8wVRSC5QSz/HiyrP5APecOYuC
JrtqIlDjMJmbwF3D/OrFOLOWPP4+LRopeIcIgI2tCgMLP9WjonbfwVJxSTuwo33k
Fk8XS2mvKcKvbUeCNgFgMpP32senBtmNj3CT2DBJ724jVD3i5A4kDZ2vFElac3L8
Lx1v2Rwpb/Zo5L0q3L42mp+MCrPTCiiQqUOF6SqKyksCPTx8X5ohRC6W8pQ89as6
d+m8K1NEvEZ2NT0kpxe7YSjuVTDzTOjEEV2m315pih6t/0DuH0NwUj/WBx06pHxw
1DbpgiOQ4bQ0tl9qa3seBKCA/yja3c39aDvetaURwbkxFAzPuR0MuF/8LnnrlQfM
6lSTfDR84Nx9nNOHHzC5RKmTM6FJB0/XBs4aipDQnbopCiTsl6cB28Fdup62L5aS
AnjKjjSwktwgPRbN7VDrdFoXbl2H3pMfhAGU9xRHVljgMY2lN8AA2NVizgylNjBW
kMyTWtyY6dYfc+mBWXLlCeQUP8140SVtUl2VvNtamK+arNP+ZEQvQt2bM0qG3WNE
kwbAn2I5C2w5vHzQ8zo1lH5Cx0LNDRn0O0MKEspMcBpBeAmilLKrnQcqyQGRIpWb
pxEOxxOLe9SC+LdRAOKk4XAvIz5zYT0fhAGffkItcWQJANFhTSH/TjLRw9NPGnZw
PkKlXjKgqUlcvPoqrOJeat6VOaTanUx8YOjvIq8WOj7m8DpT/k3FHnMt7A5Qr2eY
VzTwdtiNfqmkKANLB87JrYu5N82R/IPfddADeNbd1BwaVnXZdYm3szKsK0JSYQJk
Gio09iWAQWPDXMjutl74SPx57ng5kEFOBUVrJ+hQSNWa3Deqq79Fu+bPMWw08L/V
jNjlFTSOEUFmc+9zBki7zbsR204QmuSDxbJppD8XJnl/K3encuWmOXH8p7aJC7yP
ZgQkcyIMAYYDrFpQFvgI3L5c0YGsluOzJ6V6BCjuCkcLgiee7O+/lSz9ayOTAlll
q6AxfzJvZ/0gWkdf8LeMG05/08HvK9uSLsMTR2TAmRi40HW7fCR6++cNyVz6sZIv
vAyAlTYNov1UtRBITx0dX/Htbj50cQEkaXc0XGwf63Int4dNeHt0MrX2ZRmuFS/Q
gD1ZYEeskjMZOrtG0HafzIydExC55akzPG+DWGr8h1a8AMnPZCktwFbYCGtPMNJE
wJW5tBi17HJdyu8yUQRNiLPYAos7KYyGMxv8D6wnok6pIiqA5+Vo5qAzqnyomu4M
oUhhFPlZSRAaeKfEHMlxXoPTcTOigKtwgZgVIga/AQTz+YRsz0gnJyBY6AfGgSax
OlX4+Fdg5/8DGBdnOwV7eS+HOz64G0cvbKhDxA+c0VUzjDxuxzGlHIaiu/BSEkgR
pv84wnP2fN2yp5j3MbTR8czBJOaw+4GABNWL/U64xMzAgiX3BQIpIm14nV1A8t/0
cCxUzQxq9xxGtvRqso3th6iXVqtgVShEVdU5/yLOIMu7IDvjZLCzj2B4T9vIm7Pv
MCwCIXRB+ecrE9Aev46TJZ2WqFJyMRoybqjSGE5HvTVuYjYOmOoqBwgGcqje4sae
pluc7rObF/2LBA/WirdekmdCf1a5+Cp8MQ6Q3UOd5PYGnLCXP5Lf0LWmCPUZUvVg
9xy8LzOVhRjfIClTzRQTeKOfzLflPq34DYobTSneVWJOTFdfOIHsUaJQ+YN2MEtx
7+nB3p8urRvgoN90JE0C3gljwh/AUqgZ8SMmeVGJV+pIyMUBurffzacKMWKTUC+O
NkmjBHTc7B6C6gw3ogDTTW4F0ndiSUBV8AhJz0xJeS6Suao6VMc2nQdjBrRltAOU
3ktWsC4eVAOM3iurOeb2aCT5dRBSSPRuY0qhGc6W1astLLznqJI29eCbHUN49bR+
Gi4oO2cunpVjaXpR8HN3+W2HqbC56gL6fh+OkMuNkiQNPl+jeuZzIVU9pxMVJ+er
ZAzo4l+LnSlAqABc70KlMwv8LGHob6uEHFr9qiO8aRIQ7dkfvIuwJOXh10HKLqmu
w8q2z3Yfz6dThtJ5M0jwPQcz6g8u3d6EzZzpkVk1TExpYkZ2ca/qHRG2ia9CBMbu
HfAUDkVMdSLklYgLGYEfSQzq7rzWvJsr/GR30ic308Uz3ennkVhfpBrNSxeqtHsW
fm4v/gAeTcwYG/g3tQ8eQaDbhEShQf7UJSQzgoRwmd+WtLe7hAAXqtQmlA1pVLWz
H6XIT3xHQuR38o3PN20ye9UN+bwFxZstc7KMTQZ+ljtP/xIEdwKSZnd0l+IEVDnL
VXH2/IHVqP4dVnf/2R0rp/InQLGiMk9JEjEeQEZwolqZ8qhNd5ElsLP3iaO/qtad
+bBdkJuRz8qfN38/uMTnrXFKWqcFqgGJ6wqK8kE0clFPr9PHaD5ElY6XNjdVT92U
F3AIezXD+oBXs0IQzKS9A3mcBy9xHrLHRfStUXi7Zv8+ucTzXyzDdqKvRkBDXgP/
/W0Z5g/5bQsqX9VouzgrIFHy6fM9pOl4UZGC3g9emkkZui0njXZu2OpFcFKauJQ4
xgi9PBseDfNUd+Wk4SCxLlHfEJYVNvLhQjTHEFhLxz5IdWTufV4BJs2V1Fkj3T0m
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lu5FKzEKosRcva3dBLDPg4kXkS0lG3oUOp9GWIYJCqaxTX6uapIc3eQHC30iggSW
/it+Tlm6MLhFVA/wdAFn7FfCmYQ3KpWG3qUjS24ec3IGifPqrkpKt2jKPaU1M9q0
lH2JnEMWuXtDoWZVGoqVbJ/nrzP1cYc/c2/zxy/8VbXLHiM56+vuksL48WPLU2eb
km6lrfykYlKHvbh/ZaAvBjjscwMeZTUvwviClH4OXDz/AVRBiZO9YEx0Np7hKzfk
RyMZ+Vtppf6kDPU0w6wwETBsKSE82DYG3hUE77sq3SaCWTgYKLG85SvhBWg15kj1
lKH0W6WPhn0WKBVqP5kKMQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4528 )
`pragma protect data_block
L3drkStwCm3yXyU4CsHUBcoBwzC5N/pgZnpOV3xYMZKZMhI2mYIZ4PpicbI1bauK
ETcIu4KvpMgj+nfCNF3CtWVy5EWkJY2ZuXvlEfUxUKgAwxgGw1m3r3NYnjmYBdr1
Rs9QUIwKC+dFkdXYc2nTfxQKuDSEIQRzosT/EQHVhIyMUO+CPuKpOMnZE1MnA2Y4
QyoaUJQToi1H7rR1R3gZsUMSH9ANJMnfsJBxKYYAbjs2d79ZqqZq9zYlT8u9FMK/
pGD/62DBxiaNz0Jf+XmgZ4PSJuS8amYA4zuPo1iqHwa9IRzj2fN5mbGwD+K2AUfP
KdBokQkzE+/UDNRrgJLRi8cXPPkmK6z/TPbSvq+jbHh5Najn3etGBG2N9oR7SZeb
koKtkGIPR0waJ5ZybnbHJ0mmVrEFU/9G8RK5U9lCxfRpZNdSKrFClX+VTfp/oszn
J8AE4suU7/O/p86eDQH1fGom5OswZTi9GOR2IETrho+JBkIn+sV9OlJtBHcTuFn1
7Wi4Gpif5OJPuGPtbF0CNiBAA70V3ABD65wBAGe8Pg3BU47WzPtJ4omVAAPyXcZw
H3rh60BjQRVpURxUIXK9iEg10BDDHPYlS9gA200efJ1y2K8AJXJ0NIsFj55oM7XT
mk604N9JgwyG3Z1drqRNiyPnAYd3oaNhmuMUuP1zbbB3mdjXRHyGjaUV+EQl1j/x
kq9XPvVEYOuJBvFln0CmCU0aKgJgxxmxFsG0FRirxfYpnfEelkc2bUcxpHK3cLse
LMCQOoEQBRCiwPi3ykYPQ7kRWx9pvBfYVxCjcOjpqHQ/1eq4INHPH8BkayXYbh9o
0rEiKVcxdXHxYuUk/VdJKvOtjMTjPXk0P5PEOM/Eq2X+LH6bjQYDMlpyBr1gaE+g
YzqSH3DfxWDreoBI0COBbkGVzB/kcUOuwFGfTcJJF8PnI7buL3l7KJvdTNZwmmnF
rSb8SvLqGN4shXBOdBaQENw/nAyBhDIxlI6namOigId4D6zHQGPpNc9ty5CR6Ec0
E1NyLZ63jLGFwvkcsd09E0AEY/4ECYWWO38fAnHCbDwWu5m8J61+vA+Z3aYktT2+
0/Q6eHTRUMZlJEx86jFyPUJMRujGrOur/uumaeOnh6AO15atOM+ZwHMy/+dkOxJa
7O4qV40Ht8rBVhz3vTDm2zt/94O/Fsnj/4kdWszdb8hwMiVFCAds7kiqVKz2jO6y
XAnqbVZUiA4noaDJRSV8Hn+0VMn4w3Va+2ScE5bwaRw9Tj74wKo1mBJrCQfeUIES
E2+pFcS05zCEgmA4TFPVXvqvWh8QqmwC2WVjk0avVJUc7yuXQ3g2EbsT5fgGyt3M
qYOBq3sUroXQDO6bEz1pF9vSWK7dxcokZ36wMzsQcWkGvIof1IpEIa2lKlUD87dw
5TxZ4cdnwMo0fAqkIu3zrwOavbdhlr8YJPqw34MQSNZxPNYPf/OLQFKYyExfgJE1
OWeB+VMAQdSristbkNzeHGLg97LbFKoe6KjT9z1YP8Ipa8ek01aICTOdf6WIrAtx
44Kn4c7xqrllLZe2PIkKzNK6vrPoI070BP7pR5CfX9ZCYrykaIHEaoBE3LZeafxr
bhyRrqwNaIiEb96NxafHb3duCBmMLW+PuZmuyfaeWPZCzSfWmjPuKkW+yKZ9qUOo
BDP6R31IXYO0JVAwyZZUaLQL9YK2KFmiCvuShD2ClsiYHI9cmSPg7gu7OD/JtM6D
301hWNfVOlWa/uER2/f9XMk2fscKC8H/Sx1Q3EqeQx4E7YJIqQmkgEgV9qAeTn0l
AGqcykqo3lq1/89Gz4Oo0KRKMcCL+jqSpXXwjxbIvJjYtLVaKl+bvZJUD6nyCttX
BNu/TjwC1WB9LxV2CsT6xa0Qvz4y7FkfANP4QbntjuLVJig3qaHLgvIE9Tm81SEw
DOHRLWFRG84Yen5bqszNQfhthspGYOm9H24iippiBgkYTpL7iE+Is9SeMKPfkdnu
Cby/BHIUtFDPe5r9s4SE8x0lT6LlZGVNTtTCabllGARclSdCTr/qLvWZdGM1haOQ
JLn7WI5Lo6jVc2tJGx6U5TAtnJvsHQ5jdfqGtnxakkxae0S2cPKF9unDkGgGfJHN
FKYaucve2PYyWhSmLg2iqGfeU9nEkm4dCWJt9H0p1rh6+1Cxbuwvoydv9LPMbpy5
OB6eIDMOSRcxcAg6Jeibin1eWoRDdjEGoMHadcHFQT+8+MBsQqUL4vYR8BhbGJBB
Izs+VkLnhDesgxZ0gdehPg+DrtBzXhYFONJKsgG4G7jaM1kLV/UpiXnv6cNlhyGn
22XRC/6IVNxbzm46QJrUkk81bmYztjDtaSJ8XHQc9Ruv+9XTimYXmbOu6oMS9vM4
9HjQXspaXzt1pah7l7WXgA5WRcFhSUw5Bv1u1BA8dfrY6IAMm8NP/AzW7l5y/MT2
g2BSHFXVEGVJCjca4qHeeZt5ghOjN6af8KsbaUFjdnYZ9c2eUDb/cWof1o96tCid
uCsjnrZIRuKRUE1zajqUtxOK5hc5XVHtUCgcahKvasXhtpIQOhYr+DDbCURsrRwh
JB2tMs1SVltatLN5IV9Fkzbtk3JPaR8og0EP/RDVhtiQrGAHRmTPvZHc4HVC+9NG
tpXAD/be176K7YQsQeUqABORCoi1SMEWIL/FIsTK0TnfkqqPZ5G1Lzfi8OQD54FU
DsKXwPSEKO23iv+o338jM32DoqBEgILcACvmFBm955JiEssdeygAweRWsgxYdUHd
Q/W5CCmXIOnX5/GZNgw7faFRU4nysj679o9i4lJwVaYy4RnIyfojt8PmnqsSSgol
deiUkgHFClMSmo1M7osgnFaOhuDwz/PK1oVUpO3hXYqJrfKCqzPOV2FiodZi4WF6
aRMXtB/r9lBk2DDODhKGfNk6vgRn6X5sa8NvUB2UZSfqNaa6y6QmMJ+270Xg1yxC
chAC5pq7Ni/w21lGIHk2pjlp7hI7kbw+XLBEhx/az9qM7V2ga/YZgmKqQ8GETN0Q
ogugaOVFrkWXysia5S2R0A74jX8ayHF87FO4aCu73wsra6jGVXZzTpEH1LOLO5zz
l3zUbGqGTlueYEZAyh+TLffGfZ7RQ8viCytXba03XJq8eW6pD6CrxFBb55T5tO3k
7q2Q29cz/SdEywMFi8LYUr4Z4aq+HMBbwhMVHQXLsKFJnwZoqYntvhQ/zUox68l6
fKfoL+ixYBMlMzKkSodUXd4QOonmtipBrpBrNPJVb9g2YJfY1mpJ1dGyb09wo3SK
nFV7uYIrgayGhGBEz1Im9UKo9l6y6wmWqt3mkfFUOksIgWchUJ3aeF9Lyez86ZCa
Y4Ibl6hgkfTc+VjhN1uHHm67vKlNyX2MIFxg7agguTF6GWLxy0Gad9g8u7P3dpsi
cD8eI6cP2Q8rB/LLL9ui5ZERUAnAcYVivsb2gKzbIUfdyqwWo0XBk1BQCIDEdkTz
xKEHjo6W/dpKAXZSNx47wEtOQ8SHTKAKU7x0HiEK9eVowypxpX4tENXxcaggG6C5
UmSFSUih1Ms+pAavhqY7RP3JznPKDEeFCKTXztlr95GKHkkMyZ0TbWhwazBbAqHt
buSCy1ciaxw+PgyTYE1h5nSbsR48lIHNkLgNTjUyJjcGxPWVP7eywU1MHTGGWoj/
3KJPmLX2jh1R58Uynhw8AHxzETc3RKv2j09Cpzl0cacrUdS/89zky3P9uRW05w5H
MsaySJPTja9IcU2khavz0tcVbUetrQ34mdqG89Zu4doaUAMq08vdOKeNsB5Hg3rc
U9nBJL2SFclhO7oyP0uGzrTP4D0q1yydLxLbBk7vj6Ok8TsZLHmMb6KKHiODnkOu
fWevYR5DTdxJjV/AkSSM1npO1C1GrmBovhRETpdGoQnuBiS9YJU2KgVXAgDePyW2
nnX92ulzoKCE80lK3ff+yLj7bUN/9yErvbPV1m7u5i4DwxUotOQt+SKywUwG1zSE
xiQRpHzkg0B8isFPK0jK/vTEeOmAQFYRiIwkCWvWdK7fbYtU+ZV2PebR4QqL1l6D
nhx2jxWr7+ElxFcKHVNxLeaZEqXuKSHlvYaxw5N4WPr1rIpGAEQpefajKyU/rjwH
VSTQt10XMvXvxNah78gNm/xR0qDpO88G7iN3SGHDn/VLE9xAnyFOoMvAIiUy3L+T
TMAiP09GJu59o8L0SsoQT1CRTQVxCX3HkNgm+lLiRq1DWRA85lKbwCLfssp8TWOa
s4P1m7PX3XDYvZEnE9X9ydIcHaAqH5sNFgkI44P0q/LK46m7HXnvMKLv1HPTen4B
eqsZSkflQNAn07fbPqaPC41GcCI4OJJDL/wqRquCbJKZJEFuQxelKqwjpjFhaPgP
1lyxfmAC4sNwQ7nxMHNFf38EcJt2hhmQjtYY93JN49vlN87r/o7n1vszJO2jj1aO
dEbLXiKW0EPUO9L3NSMWCJ2eMQlJUzrkKdWfIY716mTiWUA5qLeomw28Hi3jf+3o
zBUY2qLLzl/VLbb6gK54Af3jS7etB96AvbJu2ch+oSWKlx1FYeIaYJxQUnc5uGGA
pNEU+9rMl2Pq1t+wFHj5dBUAaPzKVG/Z/zeqUQPCPObWu/A6hhXTOnpMFgckf65d
XPzLuGcXljJAvIcHM++58tf+DmrFWkrLj0QQ3DJyLQ7LYs7b6GCrKssEELToLF/f
kNYNqR/PaX4J385O4r3IHXp0EuajAjcRY9nh8M0j62KL5J7yuEUEjfvJ5E1wqVen
Odnfl6S5gjRfuyiFK4BEbiLD9+jDDvvVvky5QnAN8u/GWwo63NkNSVtXfMrRTjIH
ZfKNzGhJrzhrEW6EbGQDv+9DebfWdywiYCJ+ucToNg70msG/pYx9WkFVWuo7GLSl
VB+7DizCVSwa1L0ZWKh64UKMP2CERP7jJ8uqmBo0/CEw0tT97ZgRt4jBXTdEBf73
dtpF8nR5Fbev/tsUzCTN05NYBsZ02fXS1LUOxKFirEAZ6Vt80dd/MnfylCNJsk1A
+6lsD5wUq8KzsQBJUHzF77KAiW45VHrJNj1RQ7Z71fsaXk9BsTMqQMeoNjNzWT2M
TiOPvtFa6WNtA/cL+GPSlyHuZjUt8PNN/S5q/A9Q04xLMTwkxUIaQWJRvBCUAtm9
+hqrYzi6EoSZ7sBcW/ktSsi4+3Cp7lzEds50RWgvLiqW3c+TlQeqxKOAgC3dbG36
mf5He1SMBsl7Az8l6CW1fub458mDIsGYpe+wvqMMOFTVqKVJPQBEMOgAaazX3omX
TpybIc5TWyqcOojTqQcnUTFhuKAXcI4ml9fW+FWlybBHvvfBevsPERG7KnAlzEa/
T4PWsDJ0fwLlDt0oD1Jw0f9xUmogJtWOpe0UmR3lC4rpxjmFQ3/2PqZijUnxlcCL
wWE5fgqhjsWLAJHmUwWYMqmKroTKvk6a7FB+9unV0eFkxvQLM7ZGFuYQSVKF9hHN
Y6362FzFUXcRhpod2tDDKj05nL9RbT+LUyEwuB8/gDiBhRnXZOnR1TctlN5Xqw/G
YMOTM6ZvfsYxO41gKuv2AfSist2aJMbL10cK80YEf1y7S5ADSt1OHXE9aumU2Ap3
e6wHSGBUz1bTIhpMW8Ca3J6i7UX2O9Vt3g92qhEd6H0ybFGwfkxzlrNwT9TrNkTY
Jn6PZ240V67z/LnXXZJeTzD5o8Zp/cjCMvuw/C1MMIdh0y4oZciJf90SEJLdS8wi
qGaylBzXEpXRameEtAAB3YrwePc6Jlq5ULJbN26vV1FVIWTzbCkvvLZJ62qG6sL5
Q/ldYCVmXh5l7Rf8kOmHFlU18oAHU7V9TZBW0HmsdRBlAOdi0yVVKCMcMBzDrFg0
aHtuJILDb52X2sbPl+PWYW/QUeMG50+ONZedFgdZUyMQ+UGYu4UwdAkWc2y0KQ/Z
Gezghx6yYeEtWkVZ8p7z3b+IZyN7kdBgpyQ1CzQtuUX8vVFnZDA0xR9RiD9l/FxM
ErM1OlQe74g8JqeZMG6pNVprP3PzigZKg+k0vaF9W7DnBfI6z0AiDyw0UOAd89+A
i13TmsPHewBMIkHfrGODDg==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dJ8/L31pty0csr0zoobhSKvMKUxTZrJxRbB9l+8+EGpvVOXTQYuGOAbMg9APVjJH
ZSTWxwHL8bFXqIvqWefXYlg+IAxc2589XVPqm7E0KuPOVqirjzjWK0FLeYlcK2J5
t9WJoUfTJUsf8W5d1g7ZJatWyA6jVfghoowcg1vOCZnNc7XMeeZk5jKJidxs5zbj
lZAzBVrjUsgjONi2m75n5Yq1aKdG2hqEv5qGMdsjVA4YVlKrNmT9WalJYAwxd3cC
kaFdQQNZCV827Hu0jEt9ohqq+CUHn2BCvi0BDPkUFk6VzSDBBLox+DQToZuLXgoK
fvzB9yKl+rbIZZsKaHUl1A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9584 )
`pragma protect data_block
8jOy7ZRfxFZ2/lg/lFTaZSGYBEyzKE0ont/2rhaeYd7JMC8ws3H8JK2cj73F8RTR
JTdnBPvi4mcziN+OZcPruEegSE62HIu4fLjl92hWbrcaib1Uw0ZR25fJL4bC5cLc
9m5vrLQNFGQailwAgmavMCqPBDZ4ssaEnItATFUXy/hagnUXb6phXGTy8mMbXzMG
JXEV0DTAtukpfGPPUBwvb4clRR51XqfOoIa6FBGJz5pUPjcjvy7hs3UkdhxCml1p
IEcoQNti1TTM7QrG8TI30rYGw63IdNV15KRMc0mQ8SxridVigNb/GTS2MRJfe9p5
Qtkdbzvfg6dcjeu1QsheQLARADmsmwKLbickgrkEC+V9FB1IBZv/oheiNEXWipgM
AmWLqZjhosusNwWIRpz6n6KkXpiEOOPlX9HU2JQMNlxLNPYwr7q7Qb/nLboJH1DY
TSNGROcjKAltr8BuarsNvkHIzqW2ovUM/XGKLhohNzK6RsIDrXCePJ7JZKqz6MZq
5S+hDRSIdei277TThEdBxw1flQnJ6VVriSyyxhIv9NF782Kh4IvDoXzOMYTUNZyA
f0TtlCx+yY6a22iJccecPR1W8iptHi0aOAg/lhniCyUhUM98ijMSa4Ns7gRzjNFj
d5PxAtYzmj6Dl4feZW44LLqb7vHar1ugnDIQE2NTIHThN+7LkngX0sRPAoVgVIr5
dRL5kzGiRoIpWjryXcgvEFxzw2dXg3sCtHnwVJoCdlOTm0l8yJ6glALZ8dtPMnDg
tCZlpr0iZiSqdsbbzIkLvaCmTeJmo4MMhc9Y+HJvQVpwU5xylgYNqwS4JrEtW9fi
lwkFcIsLrhRgDdkJkGHg8tbC+7pEVtU0pT8B+EvVsAzEWmWYbmO90WHzUbpTzx4+
tBzTjjDa9O/+ACIwkbKlB0QnorTAIBAjzG13o34nALPqCU8L9F6lqR01i3CbvBCG
VUezr/VjvekGFUrx89Z/hIN9deQjOdY19zxRIyiItYrz5vUu4zTq8LF1XveG3SmO
UOc6QQ3SMed+q0Evek2a66Gb7Sno3vfMmr+NfyvoQ+SSIDdoP85PlK73a2oNdgkF
JchGUmofxATL3ELERT5E/fCkCPzs1YMDABBYBPKWAGmdrdv0tO4Zrczh8lGwa5mL
qe4RSrUGdjzzxA6+QZeohSfSSQn73HBbKyhsRbWDhchJsdgI/Hm3bl01np71rG0g
L8kHdZbV9/79mj+qcwd1pVV60N8uy/z9F5O08y4iB2I+I9bX8iXQ5RNnmjKIxmKk
KgMc+iUR9/3ADR/b1aXTuCB+6UTUjIt1EBulKmrs0HO0Qq5fCEuiUePetskIxXxt
Y2cLLisOINvbSUZivCQYNyIrpaYgyi5k9BP02q0IsExhqn9mNjH1TUveg1bHZiD4
u9Vr2e6f77kiZHxoTuDAM2eEZuFBPc93GT7GQPoOs2bIZl8ZIzGvF7m6Y0Z5lzJK
aROA48+bUMTfJ9JiaNGJ4VflPuk7sW2c4AlyrpkxCR7RzGh+lZcWnGDWeDaHkRGW
jVN7nDyMgRsAzuXa5Ifp7WRgJqBMy8GhyeqqJrvRWpDowKetaPrAev7DIzN2JKJP
bj1iqCy3vl+Ky3rV3ACx88ImuhTwUvPxe9SxRlsrE4pMURdnchOR7RSfUCck7fyg
59rt6NRaspDDe4YwOy1gvih26JDvx9pukWCIcLAU+ypO8IMHBj0kSyxif7ZKIDlE
K27QVXsLIvwulcabOUMSeUTWSKiUm3RDLEkm02xp6kK+c13E+R/OrzcwFs0x7Nr9
KC7bZrZ/5Cz776htYbP1beE84yz/rC2PV1aRN2LJiKpd/6E3bAMzY+BO4+NLdVmh
CcswXQBwFvHuMn1OsPLQ5+cRGHTrSUZRcjw+T0lW/P/r4G0N28MGGSFLWYiy2LM7
6EA98OwD0Mg4uHc68bMeG29AECmBFr/8bRMldMNIRleE8vjopCLfDvPQfzV+uTFh
tpJGIjHJvNU30cwEDS1yJZ9tSYKwShtL+A1sAe8G87HRatBBgvXhon36hTKWCwRx
HLjSHHf+0cEU7tdLnbGyaaizWQZ3YZlHBakehJ37O+Vwxd6vC6lmb31VawAfNQ3E
/guSyibt2GAwp/cEp/wFA1O9ZkVr8ifnMMj6u2VFJI9XV7e/NAuCkq7WMHzZi3VU
0rY//NSYG8XrASg2EBdLBnzzkAykPg8N6eA7yRd7yZ3aVnhrZNvGOVvdf+kxffu9
3q//mU6Yzg/3NIy2qLbtnlNTV/5rpzhRJvNNKNmEBkz26AW5CkGwdZtLXZ618xOR
5ZfeNei2rORnliB8m97IGyNlTIEIAmDyIRdzeIBw7NMjjVW6UWBZKSAIPm5mwyIZ
/5/slKkEEhYrYoqRAkgGiHZa6sERCTYnqpzpFrx/DwoAb6dbnA6Uz3Dl2f0t540+
5v5UDQsEUQBilfQR9p44RpRW99DldXOgJ3pO81Kfx0tfwPZYSYIficomw9O1oBlw
F/jldJjPKWIiCAV80wsnqlPQ37pbaxKHAcXyFI7eiXe+hesLY7dv8ZA2WL1Ymp8C
EwM4pQANsRfHXeF+vSn9GhOsLcYG5pb34V7FijM1JIzrTRw7S5d94NCNACDPpuse
3s1WilgH5I/XTxuZbMf/t5lyAzk5OMFwyaEk23rtI7Ki5Mx0HctTShhkhn2h9jih
iBeeWuTg360//cuihmq81++j54dKLz6BywK1t8AftX/ZhAVIaEuTmHR1uVwjP2tx
R35j3pYMZRFKHRrNf+xbRIzDm2pGJL3PTQeMIM5i0AJlIROPIwMPi4k0oj166CTw
DxrRAExch3DycJk6J8/PVO40VObDwQ658T/gi1u5B7ZWu/nB9yej1kCls0BWfv/+
ah//yVA5zAbc7bP9lblMgHcc4rA/SCjErm5mCB3Y+lRzvfLsTJk11NEqydikIpxm
/JGhKAf/G61vhKmXaApESl/GHXTlMIQWBTaLEAhc4g1tyj78f1rN6kuqGvTXwRf9
DlGCGSv0B4JdO7Z+50K/cwEfr+vVGJVM2z5KLihw5SD1t01ef0Did5wAW8eryMmS
NraLab3/LLI+/6BDFshJqHIKV2ono7l4l7GukJCe0U+So8ekQcakyov26zxzt8YW
o8mAHgI3tgg5bLlt1Vlo402T5a1HSQ7hBcwa5rCjYrkWsRTxhDO+W0vGb23el0vF
yD8/WKugzuXomF5kszkxn65aWbCpt3Oq8/Mo0ycotnbBKcjYBcPy9mZEoqFeoVEf
alciH+kcPWObRAYeNes1bkhBb1erq4aAf74FoUyKb48bb9zfJDrSloTCRWcgr6vJ
onviajbl/5zOzrIv4X0xk+eyvyrnT8UNHNhDpP5KE1YXP8g2AoohGK/mkXiND7cM
ZfMpLzr8xCHbAgsopIVAfFc+cB3cB4TncwediHLTx3JpC0ys8UdX39mZ4HTTbBdO
qO4Y2z2qnltRq5YoR9SZCmhNPisj84Ewxu1lK/b+BMDHjs/RobUWFUWZXQrrRq0k
wGizdqiCLX168GGT7vl36940bYKmIahW7GHTUhsjHzknEswvwQ6S4SOnOeF16HlV
JhtKG5YNqbiHTsOdUoIgqyZ67xt1P0GH8iXNvkdvuAtgwiYk1ZwrYg2rw5DPl67y
9UrkZJuNMOE5M4LnwUWBlAr0QtiKU57eRX6ReY91v2ifsUHNpoyyJyI5VmzGa8U9
l4wXblCdZdAiQaTfQkRLYPsWfjSGSkSAO7FDzs6xpXlyzVoSWMr63dsY8WmrAe5M
C+upyBrfy7J55SV7dkG2zcSq/Jfcryaf2u+PJFYHWtZZC4brDMNzEy1RiKoNsn4S
eHarpxtScu3Mrd2X0Q2ucryZqve1U19SIFvHHyx3ESWedCiFazllXaPDpd1DGQlm
tH+9AhEgvC32Wi+KvQ12GEIfWVQ3dAaZ7aubT2nHJLFuMGEyx/W3LOZHEChsbCqi
XCTNt3wl8cklfzGze1+9p3wxf94M1HF/KUVZq5SzE8YYC+Sb4CpUEBBQL882HIZX
KeuoLGMooKG+CT9eKMPGdDg3Fngs1pU7eu9BjBkO57+BdX6XZmtA9781EOYvbzgD
MNVFiEg/+Gfwy17WSvsEqIdPTXVc3u2V0wkEMiriun8hDyHI3zoMFYgZBkBGKRdn
OvcGa6TYgMsKs60Nz8nfZN/sFktM+YaVR2do+iUHjDY+QvZB8aXeS84r7tPZobFo
TCcVWPH3szQz7Y7/CvD5aM3QF4z6Ur4ImnNaAyZLw6wKg30ThGZXt+4T1noPhwMP
TMfW8VwgilTAV5+HlTDjnaKjEwuF4rNGnckuPpDi/qwOPsUyCBq14MmRqeIONVDR
Bx82aB81r9gw/AOjGOnLrevJyIVjjoboNoYVc48vTG1pH4RvNKV42KsjEBtrHcVb
8YF5s4Rnd8v8F8gPhuuT3uz8cmaanCkr8MGN/A94AWVSvkAUG5WDaiqfyecD+JQ/
DMuk+sKksfrJx4AZtCYSs9FQONnAyY8u9ezhqxIbYDcQZokwS0+X5WHvCgDS+996
ot1L5hVTGFJ8AI6CaoSB19ec86a1jlxt+mi4hLdW1fGuAi9KNsSibdLoj2h8+Vg8
CQ2YXawPIi/dG6p3XtxNe62EJuUjRWNkW9DFD4VF5fxxBS5iNINSj6ksiiUvgWsi
Jat/xCW18A85MUP8J6vjWoKd42l4Hy+sz78bdcByBjRs81hEzsVRPJroIc2MAMZQ
VX0xU1ftv/pbgbKlayuxyJ8U1EdfyVxO/OG1gArKxxckS8+Uw9SaHA+H6pC9A4wu
EfhsZnAW+fL3C/e00CjhvEmsHkYRqoN5jscBRxPKhObsv6XlvAVW9FfpK92FV5vP
P6fxV3iYhIbfLW2kcIsSuZSXtfOIBsedoR+5w1ZaeLuH/I4BaRQb2z5dlZDEP63n
yD7OPbWBNz9d94qqMCOOA7/QctLip+ONdBZNaTUlZqUj2eqv8mrM/9pR0AdBprSi
zWAhPJXiqWiTs2HZQQr8nTnHJRCmgtxMoRcvffy97dUnwioQgcpJclSH53Bwq4WO
G29pjtCP2r+EUnaf1E/e3Sb3h0qn7vCxEailZbMAXr6XNOGeSyMiQrLS1uCy0fAk
zJ+laFMmIn3d4vFj0cewvRwu0XeidL6XDfxaW9Np1wSK1hpDhbJLxNSZ1qTMXCyp
MHEV8QiFatD09Nu1uehMYxM1+UpmYbChRd0/w3D1f2l8bbN057q50uLJtNgnGp1L
gq3OvqNqhiyd/gCnTfFswI9FhMEkHZoa5HEykEfCi3PtNzWQ6hdEQ7kmkmVhf1s2
f0MHlBRpRwtAYZPrBc9hdDbahWYMylFo48FhlIW4CpEDC0nop384OXar7jkBeSbK
aoS5o2znVfOtMFIFtevC4Dkgx1Ld7QrVuyg6cje40KYOuAGNdp+wnUd4Uu+C3zUD
PY/NU8Mfao2KKbYTRVovds7DahkJvPhVPckpI8AlGpS4ZLJwvfmx1Nuwz7czDVn5
cGuDNpy25kX8RhU2EfXmI40pzu/mBwS+20sI+fG0kdLEvRCPr3JmpxpWh5BdUU86
sP03xKms8yKglnunuN+qyYy11ESAvdstIIbz49cp9kub6Nu1enRj/6ec5u0I27Qj
aZmd6b5EiL1nlAf/jvNWAaWIuLtcOxVfhmOlS9ro5V7yHBoNf7XxenQoudJULLJX
eK9Yn+3HWhn+CnRXJIZ8HyZshhgQTN4ztxZRfCrjctUabYXOGl1H+5Zr5yGi7R0d
KYxH7mezIhj4l8mzsU4dUcetuLWrbh8I9k35KkZQuNIaf0OPfHvNqUxQ8gzjCZoy
0E+mxOCYhrlxCs9AMZDoCFSOK8Rnhp/3vPk5IRvLH9wv/B3TdTIbirzj++02yMTs
WvyQIEBqwCoe0mwMpSnafhlTN1goXIQsYFHWPzI5N3gL1jMwCrKBcAPSWACsMEgr
wdLcqk7aTyVQX2GU+/t3agm71PCAP390ohi+H/h9pAJMkBQ5QfV2f46GqDrymueZ
YkYeNzj0yoX71NE/pD3JZtc3g09kDNARJme4fNvHdtP6TmsjY+yl4nUCu7oywyIR
k+L3l31yFWZWxZgtaADp42+4DBjl5C7Md6UIbBiCi+QWxqBPl0IcP7OV4/oJ8CI+
xV4nZ9hMnzaYIivR5l8KtOIw8Rp/+lI0fgGluKY5aAlbvdsP1N367tmMogD+CB77
2SkZDY+LvKnH0vcU+z50FJ2sjEjPtb+2fTQgq132/ymzjOWuwlIaKEznghYsHrYy
/3fgngmH2yvIWjKLmYusJnYqKhA3xQGcRbG6AMrSUbCCYmzSeyJMbwVGZixD3qUL
9isFYp+VUGcAIm6JY2XECurWjPha5k0i+ZbCP3cWtSAbsqnJblGyRDHg6wpY/jBG
80FbK41vDvdVrkdH+aGkGswEY9jy2qvxVvTdllyBAs23CjjRNjOeZqxbM7UMU0sZ
tXqi/SwBrxUdyegMHd8VUnRUjla8nL+8YICRySeBpYU+picjy2whUihWw2DzH85m
9aZuj93qnmHyJOQsuY6ok0Mc6Z1jjL9aisR9tTwIGrC2KG1bFQUuPSZOx5DQd12v
FInCAwfw25/ChIkuXcfGbsjEwoOkbTYMrDNdQVq2XM0cHLubOKepLnPgjOP67/73
rMwLIGjBA0J0cJzGgqAjXbptF4khYkiHfebJWCj8jEEJa7nDy7G/pnEAOSP5ds66
bSgPxLrmIyN8YqY0vhZXBRE+A+o43s6l6iB/VpCc16AUd/9Xf+XleDLuoiLW/WoH
y3lcbWZECEAaYwq3t1+2mhj1XlOKicii+/QTPoGrzhaVtsd5LW2UvNIy1szMvUkZ
9HAzEvTSxJ0ms40jg2SBqo+oottocMRs5+4TmnHgXblJqqFMgZ7oThfTEiH/1V9Q
6m9clYcHQL5sZgs8i6AnXC9dlBxjfMtP4sREtwJM07E7ee8ge0sC2yczihIqvfGt
ZTaaZeyZlDljh6rvtrUgv3bT6CQUu/i+i6YPf0eLFo5PqP4EA46sqyrBbwGTuG/M
RXYwkClSlQwBRZ1UIehITLsTzwJW9wA0ELYhstJub0dBWyS4J4MD5URFAglr51IQ
hR3Qmr22lIfy6fAD1v3poi0KWGDGQchImy+u7YwAr0IgMRPY3lD9Sq5dD5+7wlTE
6gfHBiSbUsd9dfM46y6hWO+m9nUnt9p7n1j9KVy/PP0XOUvvuhXJv7KFE49UAkLk
z3uh5cFw8rxIh9dyh/eBgbHtEkehi8wiem+jPK+NQoPfZZXdC/aI+dVjnu3u92RH
Od3vwQH68lFq0ZtE8uo+k9J3oevnnWvBUAJocHErkJM27d1i7ll43R/NoHku4MM8
7J5j4T3N2pL9Wp6uX2S5Tke7/173myh2xDUXCSuIuWpcXqU/qKsSOmG8gQfJoqFf
q4hB+qbK2nyTt91omnHknIQfhvlUTHfmPbON9Mxt7K4P5uTWtlYtxXMOSDvKpRd3
atAQjwOdSVXG+4bs7esrx6b5DAGGC/xcup2YL6K1epN4n7n0+ghZZK/fg3skde6l
pehR7Zp/4c+d0/AOhEf7ZzPuwK1rium+EmuMlORgVa38GH3ze/l9ubqoJ/86YOIO
UFfnHusZfh8Q8mcf6sHTzEh/RzjBqzUTU3S91BmK8bHR0WKzcjSkmTpBllmFYfAG
H9yRlvVhMC8QFJagplZ/Bef2ClKw4U/cxyArPCXGRCzl9YtcbuWQum5X4jSeo49s
S/4KyJFbT2f+4940ZfLNeg1vftGmOqzHrV27oZUJyMsWxEUk/B9qrZpUMRlefr12
NulIla9F0FnQgq9pVQQZFq09K9OkmKc2u+mn8vqPKNyg1Y2tAvNlBy+JPjxhoABq
bGnD/j0mPSfRiHDcxcMGZ7q98CK4lOQhL3HvfVc7ZpRQEPxZoM4s/cVs26ltLrmN
IpSE4M9yBWTG+J6lPWHC/6DWfTEc4H3bKvaGoUcmzbhb1n4KrJ6gc6NXbZAUvGZq
/DSJWndNgMrEItapWsMpwyQ1Zd3NXyJXyw8UoRG70V8W4Eivk8ZAnxxpjVIldiha
D9/ovFgRsV8pqpW1+cXCx2tipRA1BN5viVB5kRc8mA+1v9nMNANWotrFnXoWOuj8
2OlsemlWRyyl7EcqPPzY1oBTEjXgLu4HjQZAld08OkWeuGqUDMHh9AAZiwpxYXnM
HG83jxoemZVGwCVMmglECRqugA/30qZZs2JBPZPLQR8LHU2q53lhOdhnkMrv8KmJ
lBW9f0XrD5EwHg6PaG+jTSbhtuD/kKH7MxI1/jOXVfZlFmcS2iTrICQ1L8vr4pZI
3HjPz9WQAQYHjfA4JFRI0mgJlnmOLtZ/LaaZ1TvXi2RoVWwFNfgDK7sQuQQIfGaJ
KMbBGdx4L8jf7e1VAKgxXnY9wMQlUnebGmzrhVj4nyHZO708OasaoXh0IWLKsDBr
vZjrm71uFvr4vjoyLx6EgCAnJtV32uiiTeeGR9J5WgSz1wP1NIMH5UkHlyIOtveL
egM0vZJva9lpARWubYs9SkNCKD6WH89xp/DIK2YPgoMTnkzh9WBs/QVpoUuHs6IK
vwNphNHOnr9MTavjlP82MVSZ+emJWwj+WAQ2/Nue2v1kIif7M9uI8bZ1JX0/lznT
GQG+Qa1FrfIzhbOQQbd/XwxE89GrgVOs/Yex+KVy5QZtExkOWr8B+4MWh9Y85uS5
Y8bIJaGadxdsd50+GRX7RI3NJf26ZSEICckdstk+FuE49+l8IAvi8iefgMeCFZQG
bj/6szEYC6r/gwGxCY/HUojb5OwhQERTh4pq/jNsbDCq+D51YRdJ2IxnBA3w8Dxl
oSGEOH+uMQZSfT/gT0oWlqAVb9c3cUI4/9o5BBel4fGjC3DYsF9lXmcTj9Zgcx9g
yy9357n43VKRSA5Viuf9EWNmcR6UQ97iLp0g2jgvER09mTR//hsZRqr2eU4iC0So
HicET73G53p86BlKu1EZhcJQRdahmILXZIvx6wp15K3RVHqC56AUt2qMb5VVvovP
4uWbUJ9VKGjey0IKb+YP+WjbvbOYEVwnhF2tockjH9rUWZBnqUxEr32JObIgyB7N
O2I8PCoSe8eyXaNPBLZlmWb3+IjvKRU66mHKSHpr13ceYPaRTwJUnrOVX/2OWXJA
+M6SYMLSUoAvhuHN/FFJ/aqIIi3XNBfbEK3vu6oXPHaLptrHRocP+Zl0RCPfhkrZ
CiRfzZRakpTSPxHs5bdC+MUrpgtN7oz0dzhZGK0mbA4u3cfKGRJwRXKWdtAHOR0P
16j1wM519rNtt6CxFM/KizrYpPnSEIH0e/9yhOMfutT5luUCy6E6x59wQ4hoY2Cp
B0jz8gCLCNjkCoXaJGKdXy9aWWj82wOfxbBWZa3GSFzBxPQPpKeM5LZQaK+PeeTn
UWfDC+bB55i6ttYjjI9PjwzL62VudXXp09pwQ0DHIBbXkXnW8NroVzaAF9OXHpD4
X0FZT17KvYFBVsPODSgI/jpzstkzoFH+atlCMcE53C/yc86FF1y/hD/SLLGK+XZm
LAbPDEaq0odXnD1zqpeIktJd7kxssPuHf6/qpoQIiEc6RxLp4MBRnMY4ozRwMg5r
jeFVRowxU71AJLk3qHdRV3UDBDePsJWQpcOAMGY+YqwR3BXFFjdT6IDD9qSaQRaz
8irupa9mmrsSQ8xh4TjBcaYB/Rgh7ocgU75xAU0O3pYwETk+20QOSUNaek/eJqfc
xUTHu8fwhB6Rphjc3iZKCiJlRZX8szPajpmq1GNIxGJqcDitPvAVFcwYIiivxqNN
joXgzGlURaR0e6Ove1MSJI416bqdL0EqmNyFY4qsrUc4928ma/AVhgO5FfK0ddSu
qkvEUnlvu7LN7j1p7b+Jt3TKECnldumcyL06XghyfqyS4pI3o1n4RbKfFm7SNUno
02iiE/p+aYT2MKJVu9azJ5Ue2Lh3wilk+PC4+4bdfv1Bva1VKUOqrw6aQuu1xHs2
u23q5IzgAcOsQhPEpz55uSAhk6OmB+X2SzavyUaxj8KBaL6o/Gn3syTB1UAsKS6h
uOYsn/HCs/OalBRg7LadKoNrfPLygChZeGi4ayYYFF0b1p2l8BXQreGFCGrYdZ/r
4TkEobWnFoZmqtSE1geNtBCvWVPuah/NYmVa4YW9fVI/WdB0zOsE5gyDq25Xcu5o
MHq0zZJ8zX7p1zj5rSOTgn9zQ+S+U3aO0EKsVaod0YD7Wm7bAQTmPrYsSJMRRnLp
3ZaRPb4zApixsB0ztJlvtn8ChdgenbVRy54nXa7oIzz0vLrS8884Er4c6ETadFgo
o3z/HBaPXJLArbIZwvxt6tt4c+HPNWKayh63ENYY85ylXqHU9ZODQi7RQW6E1xMY
w6Jwt+781rKhbkzpvNSXPFDUMSY3qhB+mxTembHM2KzDNT6NZDFNqvNNbZuxk/g1
Rh3iNiRVHJpJgAVcJBLEs+YbjcIwiJp34uMRIGipKnTi7UIz3a/+z6nTStPypWNo
LeQXMnGDljh41EO7VwcpQ1RERqcF0T8KIC7H7hxyIdFYyP+V2EayiJ3NwpmdLdzZ
DaLCaRq/B41cgujguXNWavQ4Y42YPcIMVb/djjcBqZZ3h+kkCqqmAg3N0cdQXsvt
8Ebymr7GpfG/0rosiPXb1jAE0YBmxdetf0xpOQ49wr0AffFRFNTsvapFdQU8x5nH
pYvplT9jlwkljbnkqqoIjX6/i1blAD0L6DOfba+1FD9VxiiZl63LUxKp5bKYHAZD
dY9qyyHQo5bMtFFpzgGkJqvWCKSJLOgCgxmbzwrhVryaOi9kOtui8DFm8A/WJ9dP
xgIBteTPJQZZEgb+Vda+9eF+N08yckwRMoD1H6HGSYZS0TTUvu7stzgwD0Fwe2/o
IjLTjjMKd0vOKoBqlhywsJ4pu0VXvVAPrvIXvYSYwDtW/Az4OGKDpMDgxWjM8b63
WuIXRuvhwebTiuc/BdY61RSVHxUw4qzTV/aI4diydPxSWx4Y4iKbU7vtw1lTwxya
oXYHoyJ2LLJCS0Ywzg60+nfS1cfRTRuqc/kARAL4oBjdq5te+rSX0+YLYvjZxk+W
nwS/3HaX62O7h8gJjlYPXgNS4lkMvU0qLZmAw0IXfOi/byMxdNJik1txyQtTz7j5
+tpmDysO6koY6KrEYa1euULZUvSAqg24jm9gWyqpk8s5LV8fSapGyFh6jhsfjlhX
8heaRXhGNpTC1/nUY0uyf8hjDZuCtfGaS/60jf+ysQ0xDG5ReDq+lXZdADF0E7TK
JDDV+2hAz3hJizhrUZurba8Oq6BWxWT73S4aBQhFt03c8SvMHwGGKJFiW4TaMUHm
7awVyKhde8vXdBMoW1LzmKXHTjT/g6I6/p4nwo27padh0YK10h/jnQV/xax/e3Rh
mSn+Bk6GX4YfgdSEnBCACLEf26AyI5Oiu7Ud49v/TgHCbDmce2yooZY/NHOo+ts+
6nrzqoia+KVuB44tJioCpgphok1ow4s3FRtHFi3XHlauVlOJW/8qBjrTyYnZGzen
qjrmatUuKsZn7VaEEDSUC1h59BMKIR7a8yMDSMPnnwiMjCsNg/9v1KLKs8ZDYzYZ
zXuB9q1YU2i7ywk06MO4safZIe9Csv+8kZcfJpHVAjzlwX3TZyclYZ2M+oIh0ifc
iNq87gKdaqNBiw0bGyqSalrwDxjBU1de6MWuma9bD9b2dHaEGZlM7IkPBjJSFt62
jHlYlQTUt6w3MDYuyx6OhsBE5ny6zLpaYd3r7ULZ/7M+EyLjO+UDO9brmB6YCQ+4
DpgWtR/uk7mYeLegE8PjIpUsV5JzivGzI5qHWpPCw4ccskeRcHvT/kHVfD0kN+kJ
GeF3+aGSgdf9YHj9Ez2Uf+mA9v8gV41Gr+SgPmaQOlybrBfI5PFcHO35fo03aIqu
eOgXzS9JYTr5ouLd51PXvxCIMmdok4M4IPZa76UH6XLYELffTuE1d2gJ2SCDkYCu
CAeUmW5TgZc6TDGkB/SpvHj5kJMsFnlyPE6TqHvGMC9WOtZmRgVQBLTbVnXTKSOm
srH+Fp3ffyTYAAQH1goq3nM0CDouS5aJn9EUKIlxSVGQ/o78jTZTQ5Tz3UtefTLp
ahr6OSNgaV9etCtaMqriNyA5n6tSoEU0o13M4967TRtgZ4jpSPSkYxKGkx09To4G
mSmZwKjdW3Ld/jTBXPYkXdouXpbpqa9emCp0uBrRlgjO5N/vBV1maedSvZywrpyB
pI+eFNFjqdbDupC4k8Kmih0z9uxExMbdE/vq00/5rTrk/Gqqa84X0YnN0ILu2vpx
0BkCIduvUhCpoBuHivR4bxH4F0JvQ7xfLRwEqRrRrkZvN/ZG9xTnZes9nPUpNaL6
yOV5tEHEpcVqfXO4o0lBJusD9gCWQQ/Y9hwzxhctNkNDIgdrL/595/Z6zMKxdQvn
Z9cq47rYZrRAHVbZeQGJbL65cPH/3FUCwRdpd0M6e/sOtQdhEo9G1yfBkG4tzWyM
bS00hFHPo4nEESWeskNUDc10OYsZXLhmn1OUHtRRlgsYpnY1hJPQTKCMLvP/SVsK
AKjCbXV/oFOX198GYiA+4fcAmQpZDFJ590UP56idUsMlTyn/o6Uh13Ni4lPGNuQd
WK/NA2bZoV0ivCR+FqXW6qmftxHImHTKx22cQIr+82HPrhOdnx0zm+0hu/WqKjIb
bKo+gyHY9MtZ5D+ZynZqVkxGb8qaNMs565RSYJP/mldObE41f4mOSLhboft1YUWo
Xhz89ZnNbczGFms3ulmCluLQ8qB55qBQvADoyaxk5Ac=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Vz212d0As/DLca41+chMLVDWlyvFEi1bHZZl/ySc3zvxBCDf+eWW4v1r6BTUm+QC
lUyr6AkBNO7o6Zv1oj7nxliYkKDOyY4hQtbFzIl/di5/4t7tTZJjHJuhUtkj00TG
zT6rjlLJ6g1zQLuKtA0ZNu0JzoIfIv5jhZgX56tdS5kCtP1Jn5kfncjE3uWkfCke
+/g+bpj5vUdenpP0QpB8L2CVnV9DvBcorGvAo56WrfyUtd7npwCzwvb/9HBmHRZh
Kiwn87ZVSDK5I2ClPr+PRaC0wCTrXLfayLOMhP29rEsxGcCXCkk+rU8TCy9Rj5b6
DpraeqmpIX6ycCHel5WMtg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8096 )
`pragma protect data_block
sytjidCTDDVPhhBolYtmigefkjwAIL0mK6oSM0gToykQChPCPGq3KAcFZ5UceXNn
X6hD9WIwN2Qv+OGKERniXSsBN8+gAR7bTWEuRiUUkZZeOalcPUtlXAxK/NlMGlhC
Gnaao/5nP8+kEuvz/00oCmGhF4rUJ50XUJWUH3hKHmYUcTkq2O9AGFW89mMqORx1
byU6p7zOyJwpeBISuHbzPoJcgZHHXhh5m6g4KdqJz8Kgf5/fqMS54OTZl61oGhSo
06zIUlpc9t2zmI9cIiAE4NRIB2yILhF5NxpJG0HfyvsYXVSLZ3P40H6DGf6364pG
PK6jS2+LlRJrJk18wTslmLgThKWWoMz/iVY4091aHPfG/HxkTEUlof1vQGVvy23q
82VbLGmxtxKqL84b3RiIoGmS0sLegcEG1Q59MOwo0v9mWZG+LfSiGxn/R6FFkDm/
KWuoVuK4nfG3nFAc3riI8gOMvHFV9oXGktXYFUX+wk6b18ZeFYNs1hBjIeY0kbAM
5V48hkO5tF+hFHRiZCscYXV3WfSlKP51WwllCASLrBrBI7w3JElYdViIWzIlgab1
aZJY58VkmrS97UUe2xVQ8J/QQVjZUxmM38luIoGHcUNRUGlR2br3GDic0uiAySWn
vhIj7zNr6olaokMO5IiYdka+o9LxkcyziFzDEH1Ad4s5ewITFAfMYkdClfbm1Yk7
Jf3LNKTN3S2ieQ+EFrEBbNaZ6t4dMwIb2g5E3Z9CH7jv4JS1ZO/DqDAXoW103at4
QQH+trR2+v+zQdKp/d8vvzyoVV+L5nnYoh3CXE81VfQJdAx5BNIZCtlqx7Z0aHoW
jLg5SpHfijB5t/mvdfhDQwDfqq9yPEH9hix2SFaCb3XhLW7ZgKh15TvxQ1N1cjUU
8Fx9qiIFNpdrxeqASinb0wMHGiPZyMMcobXQp/z5woqETnxMJs/g2LVzMjVRvwBV
WtGk3f3FX203u2CrN1psuJAeiWVrdfsgHmwNy94puBvF7Opr9RbEYadFDMcdhSiq
I1atXwOeoA4qxLYs8if/MLhzlvj2Gt9QwrfQKkA2TofNSAJZP/oskgvw7pYpfO26
pukd7kGrQjG6uZdLnw7UoQFY/ViG8ZO3jxWTayNp8uSowGn4r5sUE7BZkXeo4Byb
JtUlN0oV2ROGBebFdsrHawoKKzKBV3b3G75r4W/aeZyCtHJTn2XqW6oiZ+8neRak
GPMcuAcLlMSkeLan3wRUjWUMHY53HIMmmMe8eSlDrzxCc6RY9QnD4lk7fwMMjwpA
aLniO/JDvUbrHFzvNmzHktxhIlZL9Kb21ceR3f9VQivnLwFNOP+EeawBgRaHhHT3
xn/w+e6wEZo8Ng6qXgCxgMfBXw7o/pMrmMuwB8MpMAHeKjHMdy7Kk2yEp+WvUfpu
qjzIuLPPGsQc7+baS4L5IYmUvhOvGADlQ4W9gDCczZoZ3DU7ahAdLKCLr4cmcLaF
2arWQLxNbK+l9y8OaZyZKS2HWAfzzqqyYv7VinoZZol9+IwuS2l9/dIMSxmZ8RlP
wgxFKNpfW/oVy25+1RTorbNbfOU66tW3dSI2YxSEpGURXLcF5+eLFoQPxPOisysi
xWmPWFCW4gWKVwP1JeRTStKDInwz7w+ESCtctzYBz9CRbI0bpU4Psb9uvxmkooyY
ATSd+MognjIZkpSxzpRbUgAWjFFo7f5H49lnQRuVNyg/QBa7jJ/hIIVbwv0zQC90
a8QYGbA4e7qS7uHp2NgXzr9LqWHFk90eBO3fo9Dtd5+G4GfQdVKLMHiWhFZh9rKu
+ZOEbHWKNSZOUh/RdZ4ebKSAlzwY/tYeYm7Jt1rJNxmI78FoOGnJFcQ2QXN+zqBc
K2bO72FGm6uZK0Jbd1TfIuhYLwsK8+yg6wIELGlsFboSOe4r5a55Yek7a5MaIh1T
LexxqbSducYihVLohK74zXGfZS0iuSDTeEutxDfSveR0BOYzLYZ8qypRYg7ErOgv
FguVZPtSs471ZGZArq7Obdyljq8aYOCpfY7uGXj/G5yX8FYtF0mPREqvWFr63yEw
JS0sF6N4acnB34QCGZcp11VQRVtDPW8mpx2Z5JNP07S6jLzm+cWI+xKVHylgSSGH
8q7fgYsGxIwWsZtBVKp5h8PolmaRjhZYk+MxzExVCsP2PY72S+F7WqIhZSJj8Bmb
sXCsfyoeb5Vk9h66NG09Py1QDnhOQiW6jakEwHXGts7EAE0owJOToIeEayoS6VLL
2nVv9Xs2V6KDXq704CQp/A0pLSFwrHZQWp+H/RSX+lfH99gJaQmECf8+908Z6RW0
BS6aPXmhNTDvWb6QCNGwWDvNFMLExg2QqCi6LQalGWQRJPNM60hYBRovUwx32wQv
bEYvB2Lpl/LDmgmoG7Ymq33ofvZFKqvwHjJGcx3vFGEtOZ1YPlaR3mZtWMbpDy9p
zvhsfeNXOOhWdlG1s8RdW0Fp8H7UApIqUBcMDtRpLblWWBFnF5BP2Uw94EaWh6EW
xIKtOKyPubH6AXw6ZLoQ3BsBsyMu6CO8AmAzROTnunRGLKBLlLdPmFIY+VoyIZO5
55OSE/RcFAJdTDg1buLw4nEd36YIga8aZOf5wUaR0jyV7j6ymCwta/+HNuMu46Db
LKzweMZPrGquC95cbL95qy6p9uVoIzFhySyYa5spUctyQMSYkzT4vSvXMQjMLIgs
CFq5VDROorb2GdbD7dEXKOxAm8Ecr4JwR2q8GVALTDGr+zbQjjlBAf7MTMyCLwO7
cFbH8i/oGpDaUrXiJPGO8WnMW7RoGwsHgwseir/+VL+20M+75SG7I6mr6G3kLgAo
kFaitZaswN0MWnl97B4yzIOEPp0NhPl8EFsgPfKKdCnl3bM5FTGAaXPOjnqDLcVF
wYEsDufqsG1UNM9aI/w+vYzUc6ryeMApTMLZBJKWHvh+iSUGl92p0RHP/8y8Y1Iw
pVcbKEO+o0c/q7qxZg+GA45glpgGahxr0n4qPLg2/JkIMJznp32efjkHzyPVUU52
xbhP7avizngqOBWKzzvuQ7/97ipy8Rw3trfMGso5yASCpIAOBn39YZEAn14tu+qN
V5B8EgfosWnBbs6GOYh5jEvKMNFCYKXwcWMhLUc6UDZHBvDM1Y4ABXd4ILO5PIuq
Z25n1O37YwEp+M6x8pi9mHT74mUYoKQptdA4pP5wFW34e5dZ9U37NHEd/Ziqzhck
oXhEFf1YIHzuX+63aa3AuVpwVl55dfG4YT9A87nxj7duxu9k+eCXwBOwMRhh4Yqn
WOinDEuoksWedWKuNnacoxYHnqi4f/NZndvcaMSYChxjfx+xcLkXAbdE8YFA7O9o
aPNu9PE+sXwIR36sIcz74h0qqR/ZpyrpmCSjMmRTnAKVpYDYt+khTGVyc6Ink952
5Rf4/1Jt06w2XwH2rJh/cn5VQ97azbg47VxmESmLjn/exNy+v9qQYMM3hwbv88Gf
ercf99VoOA484KCCyIlNbx9Q9PdXfuFArOluCeoujIOD2o3qr5yne+anOXRGk9DG
0MEtiVaWGyhrpInNPUKCD+7o6pq3tintgLvsrY5gnLepB5MDwVzFZWXbw4JkykA+
5+zK2TlVKLZu545ET+5Z3El6O7KIvYuv0XhJbAVyWeOLfYr3NpZ//U1CD+bKSjhO
r6EIds1U+nsH+KCxp3S8RV0epy0XoeIdMAzFkUmKQVoJzDNA3QIgwaDDbeEZDqxt
GgR1If6RcMsrhnbV+cU8VtzBxMb5oRd4ioJgxAkIEkWbIl54aJsDYekvzl/0bmle
sFk28tNTyrRxcJXQJHbWGfiaJkRHXhZvXGAYdnL7DtYZveYd8GWYWsdw93/6ZKMn
EvknoO2MFdHb23clZDXwRQ2S87Pmpui7fm6IB+6Sxt6mYmx8+8xhkP4w6LlGnHRA
pBNhqEKkx6ew8/jyRGHIt1hTJBr3ueRM3pLZjjDdJQl0UzlIQkB7JoqqHJxPx8nP
mGBND+DC38COIc00MZunz9IRtf8ZfYq81MN5kFSIW1K7c4uOpQ2l9enVliEJgMFi
oN8vRyEZek6SZoCiYsK72YwlnCEUm3ETFaAh51P2sLihKVGuoCDLD+deAGrh+Jz3
TedihHsxDdr8R/mpBx6LNWy9UIiJtuMc66X5f1keV6MLFQi17RNLlVQwlqEY35nK
fAja00BtM0354f/lI/2rdYhC7Bpa4VqD2aknSDrFc1+zUBhDRnpqoHVHAOVLe4cQ
QwVJvriPGCk1yUrmjuyl5zrSTBPkXRBMUKpKqwosTGDHneyUWTQQHMHFECLBxCzR
EmlgS96IaTGJgD8b+dTAeH0G71HSKQcleFB5aVs+qQKarrIMr2IqEUh2XZyqlQ+C
JaM3+vJ1x/CZpcjPRj5pOG8St4S37qMLz+eAujLIi7ENPXPchyXiJ39jdNHXOQx0
v6n0UG4bmXzw1WHd45zncAjcDVz3G1D0hjElbScAMKZT7ENPIrrnBUmmeMFNPr1f
3dCYfvyvjhFnqWPQI+XrGRXHtD7036HfIEH1nwtHIxVgKG/b6WNy6yUvYmCXF8oh
HUN47iY1rpbVIZT8e6jtTZW7xqctRUxtByCGnukH6Mstpw+keC/1Fv79haIK0Po5
1hsJilcId236wr9wOLkytQgrfwKevJREPHeJZcreVRq8rO+dD8lmN2oooXd7pk9q
DSKEdHEuOXq77LVj0Vkc16CsIHPHDsnfaTE1sEW4edNAGKPIgNwIxjeZiHyWUGZo
fJGXD3MVdBmIzOCivelG8mhVf8pGdhyq68/VTwFyHD4sH2THiXMNLLRht2BRDRHv
xVGmt/byuaq+hQj3ieAWWnmrASDBHR2OoAhI7mUWFmN4ae3S0Rg8P1R8dWrDKK1x
gqDWC0sgYKuLmlJxZUvsjHe/9ALWoL1mCEcGP1uZ+paxbecMw6zHwfVPPIFfm9Yp
xPXD48KDK0rKdC9Cs4lUIvJ2OsqGdvgZ1GxJZRD48wFfsEuwEvmNFALuYSsM1/3M
vCdLd5tJgpRNZMj2tYprSo5Y/Mt6JIzqIllOj2CWPp21jdW5jVXxazTbjl0Gvdoe
5pv6WIj9itzv/+UaQdyrcJJhM5+Gcg20xZ6FKhXSdG0u+I/PD1MAPQ19P+ZKLLjU
r8SpOdUEV727ZAQMriUYcFEr33cArPYXRJbbsZcssMnvTPQTxWQeQyVul8x80K6u
K6RTk0bYWjI5WWiXiBlJNk2yFZPX+B7gGD4SffYfLqMYwBS4jfxAx4nQQaWiReUS
+htL2HNd+wjjyXfrNl40DdYdHZLZxU3mCXBfq8TBRzuktitbDp0tT3Z32mukhiDk
OwrBF2PRxB9+Vg5tXScSq00UbhxrhnWs9F1Gcsg4meJ/tQLhjfnyZ/dnw9esZBYt
qYj2oiW/zXDNwa0ZLsCUhjomfpePIamo4MPWw4CcCpNYVVt7Gx3u3WbcQ4mwg+dB
zrBsixaLGjmLAs3ZqC6JO8llOzZ3DNkKFpNB+mj31gtEuG50PK9inObu3Jp7EKWY
q3Kra5Ea8E4zRjPpIkyT+6wdNUc7fGZn7GMbKkX2ofTFnKiwPSazXzmZSqLICrXE
eARVOy6Pxj9BebK5bHr/WVqENwLNr+TS3UcyGZti1+9jRLGoSaeYCjOQG8G7h5dg
yXZ7UCNESi59SMgww5xtGsnRT0zmE5it30P7EkafS3i516R1X/IpXVke1wLkVrnQ
E8mz8qHG6Ch27DfUkqWBZDGW/WG1UBn4OL5Ju2jz3TW5uGer0umklwnurxJzOnbZ
TXKfihgyIgUcuYqa9cWb+xw698+voygqrKcEv7B2NWyrI/vlMidSJOzlnzITp/02
mWoKGLKhXO2tml32UH9jcdMlSdkyehFs2sxU4iHInivg6yPEnGhUANrqbZPYvdhJ
ThXNZVVjwnsderfOvlNnMOXTX+bSsf8tIQFpyYcEBhM89Hb00PJAaaT+us+dRmj9
oH64ZuyeR2Y/GqyZPJ7ksR7U5dD4FpQXIjRx58aazOYwNXFcr/k9bSZRLDbdSk4h
kg4jQgYCr5F96g2nY98iZoT6c5fU4goGKH4BydlyY+4Ne+ZCbKqv5GkLBCbHat//
apaQsDtEkD9HoK5s2DGPxg40mk28+e6BkIOGh2LunqCbEmCqO9PUoo9JQsjRUcII
k9Jo3yQS06Dv/Dyi9NijJZ2i8d36DGBRDVCDn4V/BX7gRpjroEKdOB4ru7OQiYon
AIDyIIN3iwUlAaABeatCAC189FN5LgblQXoNZo4eeaotjgZOZulg1z06fX/JGDyh
pO8ThqOaUr8xJUTnv94GKvNf4AobGr4uMoapk1A4rIB76rHvnoAEwmb5+/NKhdsK
Owe99N5OczWR0EcIBSdDKtU0T7/Vfw18ZuaVpqX+vpRiwlDujOh3QOvZrY8CnRp5
AKyZe7nTECh6wQseLgKx8mSkjMAYQC9rKIr0Os4mu2tzYW1Pz2UD1YxzlqZGI53h
ofaEY1fy66P3wt6EpFgoyDjA/HIsKr18M+gjfLt8t976/UNuCMeveMPchFOVACI0
h9f07XmDTfE162VprSWRHDPv/WRz6EfDeKnDWsWkw8ybONMXJTXTf0xDpN+JPm27
PzlSGLtt+ik93VSUmipjqW7JsZ1kwhVjAmpK6K6ZBjzezB0KF1mw6MsNnOoNWAsA
x9UEhD0u9+LJRH/YaKAWAD3OWVDJU5A+XLFVmOo2kEuuBSbJaWyL28mJJAAwFqvu
5hw98QnbgqwXeFIz9YT3Y1SgT8jyaTpLvb+6TFn2jWmSzNwT2VNYc2NAZSjVbeYV
i6GxwMziExCzS3s+N2W2er8dax04m5/uHJGTSeZ7A6YfOY/bZrV7njuI9R+zEidG
uod7cHt7jekEOKO3pwFcXRPWqG2aB3/I4SpNKJGhKfrkiIoLIQPzwHsM9V62jr6a
TxyTKqVM+XuqbAs3FwKcqVeaMGbT6SbPL+3gO0K/VlaUMpyWEdur9oogu8XcRSVB
HZUJ9np9r6iBS6Zux5cB/tya+CXDck1tfnU5NfGLkyAk1Gw6T62vs5idD5cFDd2a
DVoMZd+7bQqUyUiIX5FCHsTDYsBf/MobLkW7ZiHZEodLC3aIfg9QZ/NZx31ESKN5
UY+tKUSeWJAZm42MijvcJeivQ6q+Om6P23gMDFkYK2gvnhsN7kXeDEcC2ToI0JrM
h2wjcSrVh1T36l/F/Lg2QMlDDG7eEfuihkRYiHjJrBUzYrmPD2ORF1HzF1239qSC
ca1ZHcJMIBwZIj5p15gSlM50feOUdDwUFWhXgg3gcSc43ef2urtRucMW3vCBb3kk
GzH4ugHEpBmYlCyyV4vqEzRoM8I6IWovpRy1x+L1Em/xQdsnFbKvl1C4Q1FPbyLp
goPQOqT+3rYJ0gSukckPZsQEZ8OG96EjV3lbOxILbkHc8xZJI2CoOI1MWsb4IQlg
6FKQdhN6zT9xHdyvIotaxEgHx+NAD+jxnHMJ3APcwVW1Q+9/8Vk2bkVSomTAgJx7
qI1oeIKUw+qpSqvylo3Ck5AE6RUmhf5y5Ur4R7txlndnLS2j13elXaprGU2f5E8A
jdrPICkEKMpxZ1xuqxQfG0q7ePpdxMKDsypAb3dHbixp5y/4a9BOEzzi3X+umMUC
BszU+7/ALjEFKKG3FnlGq4rox8ZW0soMMkvW0U2JmM0212UUrkh3VCX94+4/d4uP
luXN6oQm4/JAAoBx3rSicYBuPFFhs4u4Kw/EGhF6Ba/yGNXbspMTouV/CEaHlwlJ
r5b6jTd4EGrH4cqkgomr79t2mcXwpQMHmM4Ge7DvWhP8VGdo1f0tsQMbfJlg2/Jo
9Vw0dXlklLwDLViIVQb18tdFCP4oAVJ+lczZee4Rb2V0rv6FjRhiEpq9zT/4ZBm2
YesvqKzkHKq3o2QKLk0vWYjFTHtmRbYuYKoP3DI5nHzejobSd2oLz23sJ32Nxz6z
H93zj3o2RL/pzoU5PJ1i3XeOVyJ+Ev7NkpCMW00pKdlpZV2fLRYcUwNGIFLJrsTn
mf2oZA1cMzURYtgXU40zAgTvT1tyjeznVtu7HTM73Qp5jmelgEjdADTBg2AxLVwJ
H3wb/RsprL5OQ9HpyAylVJvQ7S43O0K2RaAVmb/eU1NAjCsiOx69LO5V25mhioTb
SbMZueaVGzOO3tj7kytf2sV984FPrGWRYuCQgKuYqf5bGQ5NNzQzxqWL8m5fTP9e
dUTifNW04q7yGHMRuDR5oR4jpOhG6rQe60RgiTYzMuaVXw4G2nzgM63FRK/E5XwN
xULs3nCf80Gjvxl+YUcdJf6/K74jcrb0wjO44SIWHmzWAP6eyU1BQ2uVEdZFtzIl
pSnEfu0tIhqcB/22NMALFKjY6GyQDqt8XuKOSqFafahspmcnps6qeUtm1Isbvgv0
hReSMfL+FEUHRXb0vgWh0uXLgRqtgtrv8UY6zFLcqJTNdj1S9ehvGAWfMKs3GDu0
L6JhuiA4NZqNqugvOqH8a2muB7rntDY0DuybenzS0zvlfHxjmMnL4q1qAjFrGT0p
Gw4yLjZxwdI57n3HroU8qfPShAAodNka4CwkMgv/qDxk7mCTjjYqDTz8C55I9vEk
XIKW1EINVgRBMedlqBXYBBZIDc2nzC0gJmu6cr9Att0/n3a83T8QJcK5I78eccNf
wRBYedtvWDFruKZoXe07B77MjO+0nP6Z9lUfW10IoFBmbQ1qSYCYguISULdYmX4L
fek9rCMCekpLgSZXhbFDSXsUC/FiZxES0p2HjlM+cFUSrE6jNtNe+ZD0J0OTfNEe
1VtxeCV1o5jEJzKL+AFAxmSdhxJDDd5Y4lP5223V9/F8hm+PeK3ERNx98PXmXl4E
LQRm9kP1CjdT3NuzTHX6D4M421aOpClGawU+/0zCkhzoTDfYOoQXRkyKuJzcbdh8
co1lzi2Iw9qkcxnThwAGYK9ZjySZl3XYpqBsMj1KZiYc6ZkEc+9wyNjd7DWF+JdS
axIseyNy1RnxNNYc6ZBKzhh+Klk5tzJM/d2RPHsXoMqy6ZJTGHSzneh5/Dhr2kv5
WZkNU+jrCHoRxulJM7VtAUtN/68PrzioYiZNw/HtY3sCDKOg5gIt3eX7xtamfgaD
9R7ErURgCBBZC3oIkn1qivvYA5VDzd/bCChc8hNike+6Q5iM8KY4SMK6GCdBGnkZ
BtewHhFNkgPoeSMKfXgDl5YXckwKmiAk8n46rBjuRAqZOKLA0DiaOZL+pQmYOp9M
aMAzd6IMekpZptW42DkD03Dt1rTiLdx6Et4yFNFw1HsfvbRm5lFNpujO7Krel5qm
K6fVbhpxZmD8QNxVsFZKUNIgD5fdNc8tE1+iTu2hxZNCFh7GeSYOjgyJWRaS6Br4
flsEkPxyJbDa7tQiZbGU3Craegpd8aIC5gP4bz/rkk8t3SMdpVPyX40D0rP/YhRS
o+Oe/xtvuyHNFXGCHvhNQFPbt3U8BQnRmDXwrauuXe7ENNkDd8ZFyK5fjyh77+Xj
gw5f10sWnBLiTBNx4tVi/Ap7+1oRC9DQwHll17sPYxq8x6sANbGh05XzjWu5m+zH
xSy24VdSMrlUsfP92h/IeaBeI6dUm/+uKKO8+Ycz8Uh8vAoldnPLGOBEavQ9DRhI
tXVFiIwdgcU9qwJ05Ibwt+2D8yokCoOCJ1EwiWAzUStj31T55s/ZaWqWyPnJUJ3y
WW2XKhgTVtZtFtjNSs7CkA42GWT+9AObtuBuXP8DHKuYQQL8rq1CdKqlICgYxpGE
65ooz722YdvauDEO601L1KWeO+ZYd8toSDHszCrfG4kDBXKUXsXbfQtIFvGL5zM9
LNlccZ4CcR0trlUOGMZdVpir+9zo6w18QTXzW6Y8Zs/Pqr6bMIV6tpp443e4xZ4S
flZAFdTjJrKJ0lzvPjLCiHmGnj22efXCz2iC5aCfRsXqRZP4UpLTKJ8R5z0VVZOs
W292xN8pErfEJ9cxp28eLQE1IzGr1baMlnYNt7sfazMRNpUUfXFuirBSwadzfZKk
P8Um3gXMHqN5lrtdUX/oUhEMMo42qj8Q+h24WOzI/WMQkGbuIV7Z519gKu3acjU6
Tt515XzEYYI2mmrEqTqceZrFmmFTWgRpF1hl06spjvWBPodM23SDHVLnVFdqTZv3
QM1GXIOfDjNV8XMYUrSJotpi+RTpiqBBZVozT9wcKBotngdQKbISxB4NxPnzk2iP
hZLQ79CP10o9PGol47hPckprioRwbMkPpBY3tcFW8WRcstC3mBNehPUFHOrhekXm
h8gRVFQGmqXybbdR8NktMFiFhtyMRxhQA9JsoSkjkDovUDZx4q2HWwfHRheFt/9Z
VpMxsjmFQAKio/oBi6U8YKftNBFoSjXNPzykwevyuAiOUOZMKW1t8iSLzryHjEkm
3CW2ErsoNvGI99gnkP4XrZRUlzxozrqO037pYuOmrutPjkGHl2/L+CXqkzywE6Mo
fE0fTt2b8PqCxlZ8mYDzHbYhpZElpqDbdfsXP+814S4fcYWSnkkKhpuFQ3RDYWdp
rb2jgeY6xKc58T8rlM/Gp5mhOxX+Be/VokLrnudswlPRmUcdP7Qw19dWNLSpreo6
Nl2qFGP5IWIPB72r7+PbxX+CnXIQqY27ZwbkGIJGgFHmjRq8YbJD4W8kD3/OG7PB
wbDBpcnjwzpHEWzxqc70MJdMTOVuJj/P43oOy7op7mJte1xqsR5WJkHdOnsOT3C7
RA4mkomFiVkksABnGh5h44hJ/Lb1S2ssHOO2AN4C4Gkmdi7AhO8UteZbQkf+9nd4
2aVGv0UmYcKcvsvhhyW199Is6LI5BTxY3r1r3ICrE3s=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hRJxyjE8Tw66DzbnEWy2ZgI1aUwwRAQC7x+M6MIunWviSh2dm2XFq1qqU4XuOcPp
kRokPcJsFsTWMnBxMHvdDXsNpTgE9Z1hrlv88fB3wLLcd2lBM36ahpIdM4S27IDO
UWHV9ch+kWXA7Ur7GG9eKA4iL2rMVroPlLoDAYe7ytXZMANh8zA64jmgoTm+NiSR
3BWv92TE+M5ySio5tqG/rotga/uNEcci1n/KJv4k2bCpYhR0F4RFSSJwbo9eif3b
1/wU6OarftcE8jHvW81h6kX9B1q8ZYWQ7XXAqu+8f5yxIAzGlwEXUMuav+pyVs1E
RykylQMcc6I7ePalihHv5g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 20288 )
`pragma protect data_block
22HpWQpkFvPmkrfnb2UqocSkX8ZWYvVtL8IUe36ktsx+y5PWyOPavkmgHOAJjBq7
ebMSZRNcsM5tS9QPBmmpJN9RXMXTw3Al0sxrmGJI1qvNAJgqcDT9jjvBGTtuvk8c
zt/KA44of40QY2RNybdSU7sgsHmQV+utMAh8U15SWnyAf0z37LGF2FAEq2mQh/xG
ofLZSDMSee40XQhvaX1+5pS/ofX8jf/CN8hy8/3QTdmvmLqbHLP2Rg4ZQ7sQ7rJ2
9oQMKa92Mo4OhimkhnYsy6bon0m+BAdBAy1UDrf4hYh/Of8unmzM8pcuxMbJZP/y
OuIdg4fNeEMeVzPVgvB6R1m+/sgROZgYvS/T7TSCU0bwPw/l6Fc/tYf8JHPfnglX
5znEUS9kOCJ43DQFslVbP8Mz2luWRP0eCnVB8Vs0KOytqHKfLZ3pdD1aG2nEoAD9
L+sUsSS50Oc+X9pm4oSxhnJVDPQoHVUI51Q+vdwvwl9Y8/Y6nM08q6yV1ckLNT8N
+UTHjztQ8htpNT+fmjx7GE9nPsbtQXE8R/EEeGVCQFG9J6sNvAjsXkBByO7XnHI/
19/wvxN0+ESNhhMsB/99lhJRzaRK3Hc2/zm8yHVy+nNXHd9ctuByXE+yFn8zeKIA
Pz+Et3joUTPquO0TB/jP6sH5cvSQOmdkctdktPxnrYC0VgkHTahgEQw+d0gwgANM
3TZj8e0lkDYzlxp4AwTO1MYXM/3vR6mlLYeaImwd4kHq26xdGUmCTQJeJpxlfSct
CI2//eOWxIVWJG6tE//GDdvQdSi2/bAN/+Ut6ea+Axjo1muBg4iOGuzgCZq+Rmlb
DJuZNqt6ZMrOyZit1WA0DZcWgEc7pnZHNkaTyPklb/5wZmlIafPRknjq1kZMa9Cx
o5SPDm7YFxByNj+6s1SV4B2g6qOH5Xdh0pYVb6sXNTojT+Y31SgvYhz9pJQGRXZe
di2cT39rjFEeBsPtiKB0G6V+RjnsMpNM2Rf49cZHaHV0VX76aPYvUpjblk44WHYz
ee0TQE1yrvmkshdSCcPX7mY+LZiVf8KXaF4jQDNTn7IUR6KL+sotBfZgR6N5snHw
EQgTCMB7OPKVg8fEIStRa9+AFRn7wKYrJ4YHP3h7G+GzAPUY/ANPL4f+PgSL8QD8
dG5l81H+XFX7iV0XlRKH6zDkXRJq/mjLYAZcxF1c9HARWKHq32U9Ni9ZY1EYt02N
0eNPHi7gUFg5/Gm220WMAsUeuZEvNScO9T/nU1MKoy5sbdZck3E9egJd5KvAZpG+
KB+5pErnnmP/FRr+3+ZY14hpF0NTEIScRZ3fA8C5RyKBawHwIKPbBtCWc8ZDo6lH
GAyequTiPobOeZGi/qKqzFjTZ4LgU1/gHHahjJtnTWzpwRCFLD+XoYBvz7wHf45/
wMoe7IJGfMPzG2+fKJPP7JxS3DyXrti/tb44S58gDFpZnueWg2NGFef6s0U954XY
614Ntg8T1wNOib8YMCFovN3aGqotjXZuz9zvxZJwa0SQKCH9OH7UsBcDtT69UACd
lZh7On9qvN76KLjNFeV4TyMvF3XwFxYJfUB4T7vZaIyzFmVjDHdoeQqMK/7n1y1P
QIgXjDdtPY6XwrpzQVT7kyHAPD/hyBTyGsLlyEjUpHgjwe92QtYuzw51ohOMy8EG
M8WrtggH0WIOQhrFEv4uO72c8A42jKgx49SNRjb9YWgIY9MFpKXm4G4h47y32g+o
Bp/He2NnrGWLseoeGEDXLrWEX36S3g7GWMrrTzarkIU0daGcx515YUgzxf6h5J5Q
iiWUsqCeNtuaeYDVTixNtegbDouc8cjwR6aQ7f1DhR+qMh0h/aCSGM1OhFs8RFqd
YCwZe2PSnGm3vWzNlAkeov4+fQkWe24V3GtzjKVmtNggEZZ+qab0VzEildCypeP3
SdAYp9hdPCmCaFPqiwAq6/Qjz9VPYjxwwDokjvLV8eU8c/+m/7MceI2gGMSs9Kfl
gSMDdsHRlbQr4ERrbXXZCLQCmUb3oIlRdtMtJrU8RHNVr9/ooZ730w788dE1Tgzq
GWwrF2bFPzlTQMbxxeGzL/5Dq+PeV3d4mMPOI2rMC7hdOHyOE3cS6GxaMAznyxbx
eAKh0SxWa2Y3tM3TZpLw2X4ePusruj5Byz7j6C3nw6TR7tgU77uENt9LbWfgKUcG
4H43TTCjZdQRnmGsmUlIpDHb+CyJPBQQYSvtJETm8ypBuXLq10LkIZhS5idhIccQ
lXkH0ZzZDgDAUoROAA8gqhk09JaEYVPMu+sHAhHRDWP4tjJWfK8l7UK7vtHb7g82
pv7ZMK+oXY+dVxD2sLFxNyBYz12F1Os74t2E0DN/gQ399kHzKWzkz9ekcbZojnzK
g2xmg6JqGYQ12phq9riY0NrxJcswq/G/msB0OqCG8xnmtSRjdYwBiMUSHKxkTluZ
bUtW92RBvZVIJsGUSz6sUrZ8zL0eaFus1719ASg0QPWy9FwgmgOGnmEBHqMWAImT
2NQzKTV5Hc7mSp/6EmBaO4HghaA65m8Vy7brhvnSK51rZKJU81jdtX1jreKiPKsx
nult0uSyU+YUyXHrStDnVS0xzieepUBSH+83Ft5LsxnkahmxOXYBYcYAweSu6c/k
XcMZui5gb+YUhiO4Lvv8byu+ZyI+0j3vTccK5u8cp9tWf9yuTH1M93gZUMW+nK0V
md1pkC3LnED2E+ZHjMVA2guAcZW2vLOXySgi6qH6W7wrlWS2+3mSVQxU2EOW/RVv
WzKrPvTiPH9O56aWgZEUl/Cf8Rq6puLEakmA1zqhMZL7D4dRGVFsewOVtesKtDyl
/KIx1Sf1oI/tO28GMGj6k07SrLuKMSMpl7wK5/47MAEjHSNjRChqjm3FSvzoDQzr
/3g+lvncOQt5nWR4wt9PrPCA0i02I9ASRkbRJ5yaKi0pLyDDKpJ/4mCmrgWsLvhy
xNCZ42e2pZUcBwM+gGccUNj1iU94agZnESOxzX7p+S9cuEMWHoiXqV/ZAmkcYnDM
PbZXYyIADlCAIs6mQg2EVdKX1/kckCBGQ5MtGQ5QQZFOU41lGmgrzaHWKZz/k+rR
H/P9S7+rjbRFR3wo8jeeoWo0xwuA+K4YIfTotjZ1xocEDE+sxJKUZu0g4jPpChhl
TtAiShRBp4JyDHEmP1QxHnTW5QPAwZpgx01ErB13VOCff50K9R1vd8mlfG06e78Q
JUNJ8zpcaPDE3Zun38/tnpJKdtXHvXxXBSoQXc6wq2PY4wyuq+G0XaiQni2HHlid
jfcNAwhPYZVc8IYu08EWODGMr3lwxEIYMiIxTHC7omNRccMe/GWGranWw9yCJ8hb
ZvcwOgCBOYPCZrnqmb4jG3JKh01fnRXpTdrBUY8g6W7bVo5vgXMi4qGxmKyehYxl
tpmI1xmgENLjQq8hmszNLrZksMkV5wLo/JEJJpa+k4GuOc1XfAq1i2gBCPPSLdyg
hCQAbFWMuaKdZescUcbJbXrn+n1TMMz4N1qaEJUeVE8YN5q/QZpAgmnoj0Rg1G7a
N7b7ts1TA8zM2goFGMrxI+fPmLhmVvvMG/jQDy227GorfGcz+vqOlz1i/kVsQG3Q
eR2vyRMNWWT5Yksw9pWgWT4B0Ny9l9R7c3lRDg7ytwuE+zsscB9Thk+wViy4Ue1O
CKJQEwk+rxATWrXcfOTeXeMlWgGaeUy5SDbtJzh/VNcNeUM1J8Q0cOaDxcPlsP4Q
ht2oXTuyZ5wd9qQKGW54OsqKujhWZCq7o1VFwvGSzYrwDoK3lLJe/LRyOiZl9oWg
HAn1V35wc0TQUgN31pGbPHFhNnFQ1tYuyUdO8FON/+PVCnJnQRp7ZPugWdEPqGu/
aXoPLU/t01whZERsurNL15LF/O4XaaeITLiyonFfZ2u0bq9EESfSVJxcyLyZxuny
SjuNHuN8hMvcd4NVlnqYoGlH41tpVo8dBnJpk4J6gP/oEBGuFlgT5BPBkX0VXnR8
BBauP2Ur4NXsS7C/Wh2dyS0kIumGtEsCLN9G53jEyuWcB/+cwKdgRWyQdaHrfQUp
YIvxqJhzNP24QWrXyMOvt/ozYPa1WAi/FrAR+/EBiv68eWDgxnG9qrYkVl2dg1tO
iaX5eKXKdmgB7VArSDGOns9HW6b2xl8fzxqbG/Qw4vxcjmutXVW2Gc4dWoG4oGwp
s8eZLLIOf/QfxGIQGYrm+uUoSMPyQ/uV5LsUn2JzphcxOiLHyWUhxJqLhy6MiHIY
4TJk9zzWFOCpSsslxClmAZyDVl2gWTRUR3c+HNnuJz5lPgg7G9nj+UJNGVUC2KjI
DvewHoK/HH09Mj9wLvEsW4MNnDRyp2FVyAt1t66jlGF7pWBS/w7BmryKkPwn68Jk
XH4XJV1iYfOVgTvt8Hx19h9mGHdWumwryiHgpIDNso/jD6T3l8vmRiDDeR6Wtz7E
gzRL6rBdmTG3DHeEAryjCmLaR47VBp7MZXEiuWKD+CtRfcoc/+KUPb9YuQnO+XIr
VT5pl6nO2R+KnXJzWp4xZEPU2J0WfzeTLpnfJIr92YBKanemWZxDB2nMzgRa8ELN
OxGUumh/9TLt/xB/+583YgpKSRVilT8oPWoyMGyGgW3zirk8HVebPXoixqGgy1bR
ZbhRB/kxgELbdmUgez93958Zp/G7DsCgLU8xVI0hnUwsiuPT19YWJZwctJm/vbtk
xzR+wOVn5y1GPEnjvuMUdc1odNkB//luCq74J5vWqguXSEo9lC21a8RD1eZQ+Zf5
j7Ip5CM1+aexUGCZ+8Nm8gCMoZoqXsYfR4oQJYLyFD73wpBiwiJvtVcV46p25DQw
3+rlPfJLn1rMICbbXrk5JeV5X+mjrg3XsdViTXJcaVLp9b4fpA70vSGgWWvFBtZo
lDe1SkdIk66154ySxsQpWW4CV+NhJely+xftcv1qFFrKJAz18o32O0tmH/6iaPGr
XHdJVHBmROO6vXYnYgM+5j2OC2chHYsxuTL2oOZT6FYxX+ilCUmQOoOTwKczdkOo
bG8rwZ3gisJpJLsblkCrAdmNW3n6JsKcMhP6s0/L+hfObUctPbnVcegwV3sidH98
w4a8tQbWL3dr4LnhhL6JbzEHFPgJpnSTvdZtRBzRt5tAizfGaATDXjWVeqs+pmt7
TP40qT+l8TmeyvwgjrjSbU7v2YfQ3qEZOQM9yPJ9qIB4Zdm9icA3kIAD4EJnNqDh
4EyAHtA7ufZMO5ZG2wQo8jEUZfVvNP2tuKoXAbJYrV568zAUsDIVACs1fl7n7wAc
8eE2fefgIm57zkAGAsj4DQeO+EacqFadWDH8p/h+OtBWZMGaZvJlCu4p+1GU/JB1
ac6nfnIHulqxQVawnmNVD/M0F2KHixCJwjf1PSd8doUMGLAlbxLLn8i/E1SPnd1d
9sA1Q8D2s8uDZ7U2RF3VxHvK5hkeaA9yiWNHeGX5QBdDup5g0f4TNYojNcgO0iPk
hpI+DRDHoja1TvwmhVHJ2P+8ykokA/p/LcgdXHVC9hViMhe5a7ZYTJ0XDcyQxHxT
APr6U7J+IDN/SdNaVsq3lS25sDS8L9xKVYXTxjzGN8n51ROd91LQf6Ajimsc5oHt
dj/1XYzUYHdIGE/NlRi6faVn0e41YMBq8symSIV559YvUOtF8tGBg90I6JEyTopL
0CIukU7WM0JYkPs8ayk7+wZiO5F3594x/fG9rhuGLBR+p6dQpIuiNzOjJU06R6t/
otimo8epUvvtg/dXihS4EsvwT+Go3mLNErnnIdiKQRFq5c5PDHlX+5qyCBbJusSK
/996cPZz+4bwK1b9zAvhJCT5sMbYJFE1bQsr2tkSn9/ohb7EVNZAtMV/n81eXoiE
HPxJzpzocb5n7/BDvaV7b6luAMq4DmisuwSk/zxTQhdtWq19CLVnmfefrpc2hT4D
NhgdoUr8aMs+xMV7dob7TqLhuol0xWmMFOdz4Gi/uRqSy9KwQAqg7YbhRbRoPT5/
UjdLVr5Ed8OqTymlBY5kDzbQplPWDbqE4BrUJ+29+wrfjMNedrWVe/o2Xti9kLDJ
jG07eqXM+P9zHJR/3H2HeQf+WsUns5VpC7t3mHxzhPLoqkFgohXyMrv78ej6btBV
uOyyiTJdPCXllIxxmIhUtFZCYTViia0Y4htYDlpf4rkh0LgJj0dB5oM/f465Sw+c
xRYUqK86tO0bWMPFyB33HVBd013hRjPRo1qGtkEzlRTxBjjfwAhZuqB1UIeXbf/R
yabELJ8rXdNRQDM7ZtnXCavfddviRK9su9oCKGal8NZeyjbR62ubbV2diwYZ2/u4
NmwwRp1aJSkuAfa8gqfqh4FSyd+ZcdgVrnQ/ffTetT+92KwhR/HcaSfT2kw7+gHJ
CCEddMn3fG8Jv2bryx2jOGJpbeO0Vw59PZhIXgDwRnEPsb5r39+lGCLNloMjNOwo
iPnIhAcTzlieLJ5aKKjBbKGR2WNRTAl6iHuTY9k5Pgmr631yzAOnC+tdNOrO+s1Z
rhgK3gUEW3EvqIGjNtPua98R/t5Lnm86HBf0M3mjZBbho5+4qQlyJ3JsdjUyWvun
RCIQcax8ZbKR4PNUgFVzGChH5/L1YDmblhjN6riG1H3hAJUQuVWh+pCEle7djfvw
24VqwCyBvtIX2ldeYBN/vIRBXZVqkOChiWztH+Y8SiTQyoZE5ZaK+08CFRPWzKCt
BJwBGOWwAd+V1eKrk5UnMepBFuIp6XpDgmfblamnBCBipguDsCLefPeNwGfTnWiI
VEOMDcouUPmdmhyEgiIgT5LD7oUCFH6OIhTT4MPeNvT1Bsn5iL9FN3hiZvtCoxs/
K+yYd4lELbrZh9hPLqUdbzZ3OGqdI05VmUnFfhPOS+LwUqD5RDTwNbdaMhuSy8Qf
GQaGOSmPWjIEMjH7sHxYEFwdpjyScZIUKGHEm55Z2tg6D3QmGmmfLPp/xJcdahvM
WBpjmwS0T5lrT82RpTW0WYfvIaxuYoxSVLqqYWqc3Qn5dTX8IbSa2Afr8EOzgYOx
6LAjE1K7JUXQt/3rGrlJM52D80vPOB742OAarFmpu+YsziTwg8hs9i75AQTCbzXz
0fHu/71XIjcWIr1nNYDhpw7wMsqBE74jqbBsWIyPbs3BHQwP2lGd5cnqHp2mK2Ub
DBx+4tpl+8CPAWjuynUC4/mvbtkjmTEEiszKPwBxYNo850qbZuC+H2q9+e8hrPGp
QCSU2OiWtrDAejS2E9y3zBOTSojEK6hPtSsq1RTzS8773GGXusjZmCsCWmYa74X+
8wYGYmtzUxAnSLQDKMe0Hmh6L7v/K0EX5orGmBJxsCg7LmDJQ+6308dd3OHzdr0D
fGoi6ExFSNpNQ9MYYDEcFREZNM0pE44olrR+6wmklm+06O9OeMn3civo1yyntRVA
QlYYL3Wlhy85Ghm6bzK60btQU9/XwXJUKLW/r8gp/OmAIJJgRTqx7xMIRluesqAs
WITGmOcHSIkvGmFBcGk1N61Qw46UF7N9mbbHmeKnVifR6+WcRFlwiwJAfEDAsQbF
TUzS3DqGjh+muhUusW2aDKcrqbIOqbooKVT+kwe5LCqJQYwI+6CMqyoQLN5c9wt2
xYjg+Mck8RbtZEePWjBsoJqsiNPLkyCdaRc8zcrUh+Zj0aWWqqzZhl1Vr0lLTdAI
4CaxUEojZJBKl/xCjGnhgU9TiIxNqHJBe5yf15nbW0Ouutzb7tmhZK+pGTgqI3jW
09L5iHqn1T4671w8sjKlPlgSWOdu71TszkHbqLHkSp0AyqVWUu4gCHkYybfC9FD2
RqLrQQQHldGRfZ3DrjpwCcm5PPpbNLD06nU0mMHixKTliYm46unrNrT/AoQi1NB6
jcgA8keOmqDojHSeavu8oNfy/2ieXCFQatcGm1b8YooAqpFQBEDS/3QM4ugRNv7T
VnHo4Eeh2c3xm59f+RRhtZTGsmYODFDw8t1QaGvhqdYf5XD6januzOQi9bPKYxuy
y1jWRmr3MMG5dl7avB5AaYFQ/QRDSOLDsG4YLFVnUvSxgI7Avuo7mRfABZcHNz2Z
Ouq+U3mI4QvPUE1MiKiwQroliyN3DBl+/N8Sst12662lr/50L9HAJLAYuAX2n215
6WLGovb7ZOBHWlaAjsY3Z0tdAQPkRbV+IyjvTeVqvKqPpu6FpIgd2sda3xDG6RrN
xm3SH6K5eP4/O3p0HiSiwXjJIgrMTSkjbxUUW7rNojRRseH0sbJ8fhj5WAjYX5Dj
UDMQ9hF2XWbpzwGkMD3t+Ie6i9kYZJTXaSyOr6XJBN+BfrXzICDwAx4FZYXFx1kH
+4lI62nwrcMk3CXXhx59tAuBh6rJjDtKJ91EgQ7kuu98X1emNhF2fcGdaIl48WdT
4biET89NLk/oudXDdFTGGvpqmAkUiE5EyehYlB9xrGLJRGYYa4jZXlOTc6kTm0Bv
Xl825XVgQz8I8SbV0p26iXgMnW4aGaD9EWVhjBR98/L3UMFXjH/7+pQWcrCmd7x1
oE5NNmq0v4sLWp/Jy+ZrNOdtHsmXdephDT048eeFZT1W4ZVnHi5JU82A3xsNKhAj
pnnOrGpn87vG3gFcTJlIQWbNX90PK4wxxZmk13RxP+IXo7bGos33GOSBDfVnNpJP
98WFVx0/m0nhT6XvnLzQkCOaVQjHjZpUj89bf1Kc1nl/Osvwv34D85EmLiKEBROg
XGvzEBEM7yiQqOskd85EtyvJtfntlDXxSDR2Tzy4Yb7i4nbawdpGcueCBYcYHek/
+8wut8OAEkh7NnApSOWJjsES5OQ/6Yyh5mxhPOLK4EOjLInIBs1v/C97RHLce+sR
3XjQV/5kbdRXivQzV2S/uAhPw3FQbFNbLbjF2lke+5UY0LkAhBilXnJkG3IR9Kof
qWpLgNBDey0EhJihPR/bUeW2qtZcVxieeM1GEa9LGxqCYJ4T94CodrDJUifnuLtH
uCjL9qEaPpb5E2MtOoKF/dve6IXY9hp2n+HfieOPA+w1o4nwCyceWLFYjtIGNiWG
626Ryhe7bH10vxtsYjj1mTNIKV5bfDVVa3G4g9LEk5HVAwBWG1rFvdmqNlZoU4/4
9ZsrCbFD3duJzg9Cf84Jydz2IWv3aWaCmavhalokGtae9E+yEFUSg6pJ+xRxt2JQ
7RxSzPf3FkcP1TpkBM0Nl4KxN+q4F4gQSZIcNevXFBRBlyXvtuDsB847b4eb0iPK
N+s8pQ62AZmaT9ASwyDmt+Fr+a6ll/pILx3gwpkE/5z7SV2rM4r3vCWhX/kYFkAg
3j4Kmin3TncEL1lgg14lnObl2xQcJZxRwBSMh9YMR69Eiq4Q6ydqIBMYN8skOU0l
aKx7pi8hQRppTGwD2RIGnlj3rNaZSEpZX+3Im5H1g401EOQ28nnKL4SuDlrLWybp
JMcMoH56u7DluEoZ0SsWnhWK+cv+yOlaEHRVbUWTVpD72A7vImTZmsEjnXC5LGfG
zRxwgsm3/lC3kt6e+06LhnwH4pZiZ/UrdV9AFr7aKGzVyZ1jYyDDkkh06EfAm2d7
TK1GuR7pvO4UCb+ou8oH/2WnbXPc6xdPREydHjEBUe7Hnslywl4IZhX1LHvyFa7p
LbaUT5N0fXlS6tgx7NXBNTz8druD1zg7K2JGczDNqTvIhC+Qs+dV5K+AySfEZR5P
Qn1GFb5kDf36jEe7ThlmL2RbFFKw99PedBrDRRy543K9u1vI0JeEWsEWxrfjsFk2
vr/xKp0mJA6MrPpfbD7XGMGy9BwICPrTZy7kKzgZ7yU2U1n83EyZkd7yV3tyDac/
+WUwg0mvgxr9AYet058pfJOmxx3qSilwC8NrNs3V8pAgOHv71Sy6sxSTipxg77Rw
V50mF7itSwkzuB2W6tEwteyxgmv3HQxGb0e5YmUl/4yscw2VzZx+sSIvl25/Sduj
lZLlTro6g1amM7Ki8OUX4f3kinQ1orEil0asQjuPVWn+uh0m1wQYtjttfl4uWiCo
FgAExopEIoo/ipUcRZacmxeaIAmMKHsXKN38JqF92wvsrJl5Z4CzgAgUPOTLnKhn
j+mt+d7Go4PtzCYUl5xVRXfQ8cbC+P7QIt26/jn4UdNE+9exSEtopx9lenaRXxLG
NcvK8vz9T8JBuF58w7Ay9fmzsk4dv8mO1D31ZAEvLhMg6bLQIw6/O+NwQzogoCYc
RL8MG1y9YRNYVCm9aRIHzcAtfnhdtcMFM+26SIv5MoIND98W7tGb2Fd8PznqHLIS
gPhZ/cud0XkJ6ybnR0EriRdtKwy3NfUxaTZcIybnhIId67H3sUI/64WoLCmccfY+
HeJ+v92X8THb1lq0mvq7gXWd6NhYYBHOo+PDnGQzjAlb5TQWuZ7pXDo4xzbB3ndC
fRzY/ZCnFf0osd5pqkUosNEVXepmqQYD/0o70BnA5sbkWTui25VEFunNgvJrlA7t
PhaExXcYOc+mFy8keRjl7whnEmoch00CE1Ar3UrkKTdObG5YAu/i2Ub1UUsr0yQX
8efUa0+u98d4mfNsWOZz6jIX+pCro3OzcmxJND4pTEz1CK+C6yPBMG8eWeo8qEiR
9m8HUjDwXN5V18Dq3bEoYuOhLHLN7grDbSexoG0deVji9UYd1xxOjxZcU/j9y5t5
0b6If6GttQMfI3WzVcHveMvr40/lQzhPZV44K9REta09Z7TP0gRVZw3t7OevnGyE
fx7/lZCaecihHebCF7Iqs/N2XQMada1USLaMWDflzcsZBGV4mTgn1LiXO9gfda8p
21DN01GqNCHL/A32zK2lLMRy6udeAN7VLekEt2skLT6Lh1Rz+FkboVypHkCWvc1N
8CMfhvgpL3u+NZxmdPlv9Rgzdfbovxun4mnfNYIQ9FP6qGjS5cRGuXMY+SP7oyvx
8C5fyvYTD5yGB16OVMw2bXbTpCOFi6JnDVTVUz8KxK/7cooCLBYEdr3h0B51pRj8
2YrLers3Sr59OCypqq+0YAWoRmVlg2Om5vhw7k009m8DTTEInRrM2eYKOKVgSsw+
/V98zWYS7V0u7ZEY15Q8KOqyMgJ6AnIFsqWnwQwMsY4rOY+8GAyzL9AJzg9eLxyB
hG6ljRPjBsx3SbzxIdE9jlXtIL6PTI4pEVMrs2YZktY6csIo3pW8Atba/mtGwFix
msE9DgLfwGZoL6+QaPiP8NUAjw1O64/Z4M2exuZp16ufx0BlMEWRvVAK2GA5zEiY
jQhB102SwBVDC1vkevapkXbuph757MNxhFRhJ3BQBupFieCS4eSOMthqAPNe4P/u
U3oNDkjqvTeIXJ4az6ZJJRtirklpRDX6o/ZZ6R52I3KjuTjrIsJbNiFrhz5P1kao
DyozstV44tQHnCcx6xeg64vS2Ns5hR5mrfOBo0OYuBFMjxxDK86JLXvSQQHY7uKp
2MYKm2v2UI5NZ5JKFFHJuKE8ZQx6+PBeNQ8hCoJnmMAwUXp+bR7NNeRH21ZMpkte
NrEgzfvkVXDqn0pTW7z+rEwcsBWp5Ko9OFSBz+cXr72LFRaFmQibtUlhTd/8beWu
SRgaRJ2FJcqcFt12W4GJ8THMTOa+VJhZNiZ9KHQeaew3QPw4+1EPcmPAjmlO+9Vo
IzYxB0tqVXWWAZmnIVEvU1w1LRrGdwmUvsgvbQUeYQXqGwTNaoRk2HzXW4iWLnCZ
wROwdb6WkP2FP/s3lVPGkZ7FNFcG0+iWkrtVRTDf9UNj5+qBBcRQmKVys8HsAhBb
FVg31PzMgPyuFwCGsVTNk/X1xHfLrdr4Mw3VtmHNRklS6Ub2fnzvC3pgJUNNCdRN
7hrCqA+3gM8x/EpkVAntkltQi9axY4gleDnbfeFrd+DKA8wZ/gwEcdQhKj6g2IIp
E7QuGRYDni+j+9C9A7t7nkPW6K5H5yvU2LeLUNn4tmjqafzWsmox9p3qMSwJyB85
BWOK6hYautRxZH6WuedfWBGcMkxqRouv4U7WdW/qzWaGEwiPNeDa2JLnoKoAKNtN
nfleFdf2eJht+/4Zy8TJdJKeJIqjpIZdW+kckyaphqDVaSJqGjZJcOqPVz0901Zv
69qp1+mKaCWGd+tQBW+vdKkNN970aGXq1Fy2w0XTteVd+0fXLXjAcnPJQkkuP6vt
WbIENdISaDBsgeFdywl1V8ldWjb28sgxFiAQqD8It6Ev/wMh7MY8Ei/qF6yZZg3m
hnhF/yW+wBSP0VDNA2GnSXE0LhBn3HS7hAa9JHMsIhtGAb3sKx0aVgMU10S/vw1O
54rRXA68n4kMbCnklmtZconKMqlpg5Q0VGVnCczQIavAKTHevUHF5WrSkbEdbPv0
KBINxRtuGkh5tF03PC++JQk3WJNWYjH6UpzQynvz1BAvwIbae7ykIf5GiraSrZGj
KDF4x8cxZkV1Rmg0ssXpH/cx2qgXlk0gaaAhKp8nFnChY6HDGvg80UlbDCdxM7Qd
xDWzFM/hki4RSg4RdJEq2leuKaWNp9XRB8XQAX9HOWwjAcCgcO01KXhDgw9j6KHj
OozP2YHZXEIsMLh3H0fnDbxfhmo0i5pNutmdOrZYjZ7MdUoS7i0HFqgaf5kxFU8y
oyGCHDEqqx7FdWowvrGVJ1jTH3KyoS2EjpcPQbSfF0OP38kRf/RGXQShdzl0atYk
z1gyeBJ+zdCyL/tNPcw5W87j1h5yH9uwKYALBS+tWzIeEl7PhRc5mCeR6yG3dX9r
+ALjAVbquXpunM7tM8Lcrjks8Ay7wHh2BTW2jIs6qFh/S/fwtplAGjGhC80tpXHY
j9tgm2/ThrwAx2AY7UquObd+fbtCNHK1H9+DuJ7X6N2JGg29mMb9prfVtN+GygT+
yT3C9WV5IFAFadahQ1TSpq9OplKMr4htygcMYC7kcp9v3WsiSsm39aKdLAv7KQqX
l9eBzFeEhLj6m6/WfTlDThq73fXrjnm5m3uJTQmnKwUni0JtKLRbCB+kpbWgWUWK
mjSIxqLcdFI4dIzy/1UoRKxeQ4CO1PBWqsMl5QpjcTzk8Bkd3c1KTUcuhBxvbcbN
YfvM9f+sJxa50wEHJ4Tcy9eQW9l0oFsMRk15QiZJn6fp6NdgqeG+BAgbHRWMOAFl
2ARLbj4VgILAjrsClRsXJbD+RPFgB7FJUQWO81L/8D4Sim6pfH4i8UjrcSoM3slY
D2vGmmghcedvzLQ2rtLMdvOauWGjpxGoby0UZ3sx9+KLP+wB8NmGH08Gykvy4WSu
ah1OKlpUu/RdpibWSqd6PzTQK9ycqvUa/d1+d8kTUtg6iO5xmjrDdBgAMgSQEc1M
TBIEqwyKmUpN5BpjRAJ2F7rBiZ3BnFyb8+3OwMinqkE8CO4zgfAYTSuoemR2zeHg
oH4qggUvtJr7X5BATzmA1WVU4xXAK3hCKf+6qSR0ODhFjLzUdl67pQpb9DdxCqrJ
mhOcEggcbmn/BxGDhZ+9zpf+LSPxvYmzZcb9uQGPbk4kJaW1QHMBxvuzPKxhgLbJ
f1HEAgkdB4fNbwssbYZa3IGC78XpowRK8InjmBSFypjatkjBzO2xbv/3qxzLA4It
tRoJAMkP9STOUtmph3nfeC+Hv8diwb48NbWH/zfsQuXOWyMb8Ux3otYp4DqzLaPg
/qx+zxqBywesd2lWWg0i0QYS7QQo44Y8dksQE83BHoDrqTi7C25Akoydy9TDWEqn
K4ZUmhrXolt3B6uVo6fikkhwDF1vV2S4wpq10h+TxZwWKBjsP6/SwDpiuZ1oK0Mz
UtuYywr5NAr5lvL8vwNG5f1Je81ZqI4aFrOmvF4t/7oxy9FUUSmrGO8Ma5xk5abL
HiqoUMOBkUDU53cBVrma2Uy4VIkDhwC7UqPDK11orsbiV9wtVqpOKpaMfNjb6o4B
8gCrE8lVHFKwtsqDr7IL4mqbwQ4TRTy8xVakkmrzLIQAxdT8ObwUXHrhOaUq6A4H
KVPfi7TBfXdcDr6ScwIu2VERUQaDnKr3bD7GCJHeQf+OBj5ZaPiJ2pmi7GQfpx0y
1bIqt2/+ivkBfvovRpUEwi8h4JbeYWMqG3O4FbVwH+UzpqxY+J0cr0WsNsYNgmHO
0yZBaftHxxy9gpid5FIGtJT1q26V+dP+KqoTaQwTjw/wK4wF1yCvBW8ReY3unQ+T
TiJwwS+C0j2z1POi/nquYCHO2gTbWA0DhpaXjGBQu64Yi1D6xhNCziAfx+XhwsmC
UbJboq7yFqYJzUAkW9lVn0qhQaC7L0eXArrQEhDNe9lgl0/IQegevZ1ZBJX6l4kp
svWGexwIvEvMkteFJWdHGMwKmZDU6GnvTwRpYZDVWpDJX3nnPZIKYuSw4tt3+/is
U58+T193j6dJSF54GxpfO7NpW41o/FagakFZ1JoCQI08r/fVhDWet16+NEutOuvC
YX5gggAf7zdh9PoHkD+Vzb1qrbWqETzQ/ObOQ5MilyxUsAajcC5UWGDAs4oWkfde
KzCDY19h2na0JZHRq/eoD5s/UQPvlFO2v7DxzgqoP7AS7wMiqizNxaHHLUeS3WXi
oAYI8JS7uwHL75ssRIZMoOJ6OOykALdCj/70LEuIZJ1CODznpUhB4+s+d1YcXNoC
8QxKCtFwBs0nuEmJukezSgLSS+TDEff+FVBXUfDQnX9AhvJkBjlhj5dSWeS09cSv
Pji4rWKcK1Eo6UHUtVsXxVf6P759NHv77xCKz0UNChdx4sXFAlCPLKXgc8gxaupS
14YOE3ulCBoBbif7NCAOY3eT+/1qgfGPaidpTit0SLHOBEtDjoaykoFq0XpcEt6i
RxXN5LlQEwHWCvt9i3wV24NkWCcUt/hgNAITJsQa5dxGobvLRxhiqErVbPJJw8qL
V/yOkMkd8FamlJxseULRhRwV2fJIwgYKcS9j+gWfF8tMjMox35fRoUrOwEcYPuyH
2g5+t3iskQS4dMjEXwHi5T0XTQnFLs6FmUVMEmgABcGylYf44BQ1ha886anrNYSx
BU/sbPZ8Sr4nJAmJJ74OGravRaw8YMQwZqA/wDqmLf159JGmD1KXu3C7vTVVIMQG
Xx6Qa4dMdls5s9Cb5D+lF6LTt3uO5comfY9ZgDUV9T5iCrupVH8gP2saIcet52FK
bC5bE8QwNvojxPkKJkgc30dc9ZRhkoLRKcqGhQaq+bAWE0vzlvs2MUUAhfSn41mT
nFGnAsRRUy7NYEmp4K5oZPmOIDTaum2/maluWhJLLy+ny8E7DMJwUZNn+1ocjX2w
L0ZQtOJFOCUE9VDOCk1U1O6mK6ZNQBRlmSWjOeZ9Frm4wrZ0SNX/55SnNZncYSID
jBJrJii4DUzMDP9DWEMURVsIWQwuaisfgprUxEPSG+a0rMv2sOCIxhUXlQ47zbn5
x4pCr4YaDJoXfXleDXcEkUWomxTDJwNHFEm3uL4PyT4zURm0enrMYyfn19XI8oCp
i1wmp/Oe245eQk6N4ZBfg4t9zXqSuwhXBW3XkbHuRrQjDYK7OQNX14PAl2NWyVv0
9XV9OWPyinKx7SASxnz7J0SkX/M/DWCRoy0GQ7mWakHvV2PImHxXIqROojFYpot2
0bpQ1LQfiNLYCp4hAsavj/7cHiJNqrzQGhqf7Tr8syivJp6yXjmzc1m2jyPgqBVX
X0ApV8FatBGWHqWHZnZx+Nkc91VUz83X7L8mf6LdR9Y3/x3nJ3hBMEZZzYlu6RoG
ugcOJYYL6y/u9cGgQONYKbkdiWDN+MvcnHPmVDdQ3EkLz0UpmQtGBBvL5dTOkVbi
O6LeNX0Ug8N09zPCMxJeLkqKvKv0nfu/Jka0A9dKMtgUD5nLgXtCc4DAFAKUtEvz
+C1XaCi+HJhe4PVSiXRkwgFEujPBLPEl3XvPYAv4da14Y3wjAJUn5GoKjp3yp8mr
1UQrSIq0JRl67e2paYtBL4XlA8kQdLZZyA48nvZJmZgpN/QQjjYJvW7UcflahIeH
d6rCAFRLevXdm8r2WQnI6QdEIuLVjFmsieOnQ+imI/WSuBSQpdRqNP2nBzdaBMgJ
eAQyyrdCqVNsrUvuo6i8Al3NhHTjK8rMjnXsxfKb3Ic8hTEJj2m6HdBOjwAIlLc4
8sSuNiSRvaT9jih/m+3/wX0NyTC73Wek2ojqXad92DMA9MwyF2SVVK8B0iVZ/6Dz
CXH3tKx7A8St/5TNVKzvBzjenaSuXq+aN73UYJF4pM5mNewtDnpOg9HDxuraIpB4
IFenuOGaTnIqzcKgthrwGBQXhebeHh0atmP1Ug0RTSjvTPbhufsZaBqwp4ZPzAGh
C7uw1TSC+uKM5gEpz/4cFfa6Q3LFZgQwGkYMsjxvLKDX9f/OfkGvfYzTU5wOYvHY
93sccaTVt4RFS+IFqoNEZKgd9HGDxZ2pnazDQi1Q0MPch5OHDOBWUrw58rlwBjwx
5hQcGFPmmdvVGrzOOyXch+ftJQxXFiVRHamGfEaQ2XPJkB4Z4mYQPt9ciZPkOH4n
J1m4B0IZwkG+/evim05hOwgqxjJlmMfOlgy1hUh1gTAnnD3kkI+NXwzUwVK0uC6H
GutZu+KPtfQqUL9CfuW8Sd7VH9yxWFHtFtryJO0Z6cEtVr9dcHZlWgK7Qbhjb22v
SpBHtR9q+WeH7Ap5BAtwUvdCzIUUsm55EvwU1vPbac9cShFvoThhnF2SQhOHR15n
5vo6qp41rrCWisUmXoN7cSzxU8NXwNEWtv/BKY3J7Y3cM5lgrgvGpP7SL1aU4GrC
nUsjxvuWnNh1oSiEMXrH3m+PsD0EXJ3wM6YKNba0od8e0vEsQWgyyJlCGgjrPNsx
ICbzyF2H7RVkib5nX9hEIz/AasHzyzxIxlMT3ccjM+Y3EaqrSOmgvE7HcaZyEZrK
JkC/E9+lYNKpp3LrGAcji627YwfSOmqoNiXndhoUV92GaJgmbxB9yK/DD9y53jzg
ubUz+4DnlhNdtd827O/dFePDRtWZ2J8m6kG2dribzQYvxggCC/2LcBjYUOBCOGqf
fwKYw8PBiOkCkXdm73TrjUd0rdNZfMIMx/cBVbTeMQ2KHM6GGrNGnm50/Md/B1Fp
Q5tTZvf4qcfo3NBq0uamwWsb6HQ4rYVyj9I2mIF5Du2zMvnmtTpWDPHna+Trmvdc
JpLlfkI2LylQcDfRSLmsbqwAK7+pl2ZwPLUP8tIUEX9yXZrLS5D9byQ0sZMMeiyM
zIQoUhqbKJiVXG5WFj4K5fZgsHEh8EU8ShVL4xPW8WWGeBRf1tkP+R/kP2ANCt/H
3itmZQkAwXq1qfA9u00DMeJ8yMukAQLeuR2V878og9yHln/2JuFYwHValn6VC6Ox
V+ZHw3SM6IwFjjH4fYOA5I3m4hEnFf6DWoMp5cULD7abrzkvhqju/qWuyYY2NbXa
P8nNrUXyyoh8JLkpyFfNHeYMJ0WFTtjmQV2gpFoJ/dECq+67Oart6PR1xJQZn7yI
Cg7Zp0FtkDNrU5s98GT478PaNHpYj6ywcDNo45NONU2IGP215NH/rZ7XGWWaCyD6
/vtfzo4a8+iMhx1l52rD3JjbHPRxDg70FbZ4LQTIg/V5pTXWlzKCDHL2/EbZz0Th
6E6ZdkfKNKOIE7yCDfK7bVQ1AJichyXhwOfIV8qgLKcZA8nSfeW6NJ+gMTLEELD4
XyCgGE87sZfTb7xLsr33AwwBMYxLz4qRmnaZdGjDpF/1xIt3RwvIYINh1SrMDrHF
Nk85S6ju7PY5CFsHByveWfwZKexDPk9VERu62RhCdWh1KeL1UDMudD5t7NAp4KCy
6mbnmuoqR5fpR3VjTj5+TIUWt4fiXVuUOA8HsjRsZPryjkVfILXNp+8jN9Gk04o+
lE5x+DkxvD1VAfMmwSpCrVNusPd+8HFAl6HPKUzJK/ykT0X+zxE9jpN074eefGSp
YK93psxLcIvFli6Jitm3Cs3KghY1UiWbNML4x2YvYID4I5g8fEKC3+8LoGrxoYF2
K0LxGGxeTo60FZ7byPFuXiWmiinDSTSm8FB0BZYQPb6El/dr5UZQv7n41wi1hp7n
WbfaeV0sjIySQJ1RZUdmG3YoUi7V9Lx7KT5DtdgTRGAukj9b8tNJSDoYppHofFtJ
FuzFl8sViENQHeoBaIp55s89NfIHcspjVUA2em5SkKcybGCtSUu/Spt7dgh8D6kb
XIGc1LzLrhEzss8uUYRS5NuyDBldDnzpKiOzfCH79Yhwa9zXeQYZt0W5CiWHiOwi
KcQQMCR8IDae3HItUy0bF/FSPGFD0vKA5uV9v1+xTT3Lo2NqyRJxCAfrIRWMSY4p
3+QkIiTQ4U/WL1iB4iSKso8mDN0W7AfqUrZ3UVquWxDc8lzAjOO8gYg25gJKPfgd
7t7AUsWIDnszA0cSCnjOUwsBkRueydix81Ccsjomj4epMpSF1ILjpUaprxQ0Kyu7
ekjF51DAC2NhZKEYEbEZwtPBcNdRBep3V+aGNFYiFBuJWd6xMbxWtmWrA6j70HuH
euahLcq3XgZER5VCAH39t/RQ4juFmXWNv81q95DrksYF8XAluvoyAa9tI02s6Qkb
F9zoJy3bVpkaskVJyoeBDxPRHjuoSfv0ME9zBFDubPqJGffP70FGy6XJDQ1sBAUq
BT983SY1uxmeJdInUh3jQI9Mq+ROcaZtibR9PcwYIC70QoJtkalKt80g/fZ6mZEX
cWTY51ugeoYZw+7/olj7K/smZrNZy7uctmeEDrFm6zwmb7Qw2mvo3Qqf10sdSKiS
BWIv5u1jCcnSzNx1vCNdT1CbCLVRz4dnBhxMUxxf6I0FWTUM1nBKBSeYs6lhD+Lh
1OrdmLeEr7jf/+jxyKEdBBC3yFtlGhrEnN9w4WL1RnbVrg3WK4E0sQuohZlWKqHw
rg+Q5etsk+QJsKkUHhpJeeqdGWFJyWvNQKB7aAfk0nUDhlM/+7BJm4h/3XqlZ/pW
1YTH+HjipruUM/B0byMD0yt3JSiRQGAvilEg2q6px/jxZokqxYOVBagRbrauvSF4
1w/7TTh7WuXGKwLQbcrpdopG+jt0u3MKIL3FwzfRTvIajkGKxm5FJWiaK9ic/BBr
o+hTt674XuU/5MOybAt7RsY3qtDIcOE7izVhCuxIJsj5Dny1e+fmuWRui7nUTv8Q
FFb+YK1Gkg9r9s9o5Voy5hmsW4mbRisxnLyeowNU8Ao4gTMygpWUmVCwq8I4n7+d
hU8Lcjfn3CeRL7dRAH+vKKZIBVMFYcCU1b7JtAW5hl0iChDhOpGLCU//pgpymqA1
/x2BnV89dcevwY7Irb5BHo3EKj1z+qz17VGYYz13pfoAHEtegUx6hN8nzCZev5hY
bdBmAV61YeB9KIIpOid+/rDabBh3WhuaAh3hd8mgW6vFLh+KLen/iVhJCoNDeY1X
iBDwVhkuywC4uThRrI/gpXSG9UFi7PLB/71MY+4kToqZuV4zwy+kYtpDUn3zPyJB
ucp0bSgEEQFjzQQpCaQZuvyTB7gpjZLa62uvFo+AoqRcgJO0FZ6z6lv9kAvFPkQm
7idye24W4/9K90+1vG6zr5vjZ4/X8Q57wKkU5Cqi7q7Vu31xXLGlx2VJQG3hrULP
ph/LmI8jxIEhucRWP8iEoyEumMjk7PxAIYjcW0rCUJAZdsowjKumXYt2u5fbS2P6
XmHkY3POqMWJjX66OqsEx1EaRCIXK6cKSA7fvfehmbqqYAxVp2ZuF5S6RvUNpVPl
kqqn7FTePEUNd9KvqPomB2m/32c0j0h8sGkkdwh1CQeDsOkwAt3hhQKGXQsMbOAD
+mv5WD5Oe5E6u0+/UY+KmfTqmNDP/4ouksgx8YZNAGU5YQZ1J+ZJuJKFzSLvXedX
onTNHeTTDGqIS6lmKIe6KmKXF4lrz8GHUlmQjb7qGXVZttdWCVCn92VZBwe7TaA7
YCRrIT5CmBfIa3baWYX7KJBbjHhXt0SzizUtSderZoaFNAXfKyU7itF6iulx0wWJ
0lvBF8nz8PyH31uo41lS24vz88HaiphCzKSXnF0S9h6+5OEuk95PFckN6VbB9FKu
JJxxL1W1Zb7kzZGZFgGmtRiC5n83Bve+ycN47ZASYGLCj176hUOeH9Kc5hxxydGj
dbsmiayLs6TCsNwuIXfl1ivbqrm6/CqcBtr8XpVe5G/MJpesZheHc+0wAnCrBO1i
8XWu1YKeW7UybHp3BMMVkiN+xk4bnMuoLfHD7G1eGrCR3ZjjekLjZl3IXIY61fT6
JbeCKrt0kOeMOgy2xfqJolPX20COI3GFqYsSgb+w69gQ2LQd+s7HHBXeODS6ur/x
UK20TlZzdpwCPH8rv5x51g+9Jq3YiEBcFO3DCB8KCLuezg5gOLHzvapRKVvs8siv
KRBlzFw+x6OORbYfoWFTnAP6Sl+LPVbbHIYHF2TqclNjrUxsm2c3nShj0DdbPOC1
yI++Um2lnfsYXaVvigCbxu6rRWzIEykrqWKY/URiyN2hYmgZvNE8k6ge+6t3e3m1
rOKjOuoolhzV0/WYFx8uwHTW3vtzgZ05ma6dQbEs0P4vZfwxCnKyWDgdNwlh355s
uEwOAirk1Z1A2+3nuVrh04GmrGEcfIaDSDY04QjVsF/q+tlvlsH1pYqtrh2o9FhG
iX2WcBUhefsaUbrRYmczaXYbPMdolAbB0OCFmhrpA4gBBCeab2TU7wgGcOnQxB0d
IqPkgxE3GyiY1SpZ89IBiXxc4u7KLxxtYNua0lk/+yLkVC8GrsBCCo1cwj3VwbN4
UF5m6+dTNeOwCZJinA7I6kOvgsl+FQ2w78Op7BdADNUa61lY98bWhu+3TfPDsO5v
5DUY0rfJ5Vw3q9VyS1e9eHx/QgHsG9FN0BSBaGwqtnLLFqbzHTjS0aopeCaDjsfz
vyGdQ5F+bzpXjA/1Mvfw8n7WMkwMgiFktsKpYoFVPhMnKmRhtqG/UrrRPg+Nou4L
qiYTypVn867fopEp2FABs1ZHEP3NF/kn762Ezy4jXARsY1a6135vryKLtwtL+VFy
qkwukr15appDkIfslngixvy2CxdWSLhb5BgJQPl0rj5BeULNdBmJFJEzra9CNzH+
JYI2gis0CzdnwfcES7s0ZFT4SWPW9+kV1M+O68snl98ZOff5fC3G3P58PCO0r5GL
sqlDK6+XoHLBlf9zuG+Ym7UlGXAj/xRr0ycN6RhBtF/3qByRPvQSSMLykuh6fC0k
mqMkKRGjyWWF2ggB/i+hWcHTfneYTHtXH4y4LvbU4f2HtjUTVdH8CDYlnEx8jBnx
/u4xzSsIPNZw3obL5lz7gVVjiGUb+UBUqdEF1zjzfdf2EKz+uAD8A7U1XP1kXA1F
c2IB9uG6M2BDWhIV9Qcq2O7rb0peOEa6iLJqFH5PrBijw1V7kS8qzePtUqbBoxKF
p/m1EB0cC3h0cICgHyJYb+91D4zCSIgCQEstr5k5dT1+GhXQgszKJDutsGC3zLoB
+IBSkjpA0f+XPHzqwHViJVEbfOh6b/Nkd7IhS7oGeg6ZAeGhWlVL9U9EK1e1xfa7
A1e/61T28S5M2oIIw9KN2qEKPDCNA+svXZ+vt/hImlQnWdmU1jZEnjK7ROxSmPDR
oX0xYMkjv91xJDtaeClkJMr5dwm2GWYGDQwmFRMvPKvzWi52XR2QSh9e20285VNh
y3FyDewEgTF2UxuhbKHC3Ea47Hz5L0hMykTlFSIS31bhhceL+yA9WtZlGPRv3b5f
/+sp8F1lmK4Dnxl+so1hGaubOYLY/Jy3g84rulENo8Ww39SREsO968m1T8qdwBJJ
qN/bsvG8NGS3fZglcI949uv1eImZ6p7sGUbytHW4MAhMjUosxLhWTicQl7WZ8tFY
9GTH/kQeg3aLXisf3U7hECSjNB+/IyFoMpFCwMSUJ8Yo6t80ed9t64fydNH2GHgh
om1JNOMnLj0Wtcotn0TGiIcGbhWwEwgkisEjabIYCDqYK/7x7Eq3TiMOm2fEzmlp
eotVBcsVZkS7EUng3y1KdSWaTXPsPHxR01sasjUhS0AQRBu4x3PAjD9J79YWk/A3
CupCyLMe1Na3n6KI3LH5/IAVQRgGT59a6j4yScHYhVyWn+2BMf2xSgQ3nJ4Lxg/M
9INCt0CposwKGL8q0C2DQs7178GDkB0UZ1xtBZH8LUYK5w0lafMwic397sMjZy07
CTvuT3VnZSS/aKKcuZHPh/mAYVNbi3UAvOFCJfO1FitHfI4vT6oVmhoKZkpXsI2x
9joIHIBJnCaH177Hz5uP7d/7nNatSW+A5sBTOZa3ZvR18cQoLSI9K7b0Fxo7rKoo
RJwKon0vlmpE7EN3wrW+ssq4Lu3LhxpQSqqy4iV4snHxc7saqVdrgKNCQOiRVQIH
xcJQp/jhY60mmVOBjJfh2vruxC6eBV9vjTYo0YckDNyfIQo97IaKONOEpIkfUv8G
FZKORDnk5AGji9P35Vr73OTaPSFtlQA93bpsasPCp2jmOTXDocYUa/UyBYvexK+Z
JlWRoU+ekfpVAjowRT6MGgxWsz2xxsJf7KdX9pmoQ8NpqT71sM6PBaF87AW2OiyA
SIuxoS2w0TMrd1Q5JuJtssMehADN3EutEZGfpkABdSeNLKpi4moZeER/qe2dNa3M
tNRRWPSQl+tmV/S/jF4t55weWBva6LT/yV3q/3nf/GrEWgJkDDpV/9RWbScjGYXq
eVyKzisNItgaNjV0eZueNzbt5w5MlZTMeNWcNJsAtXyJWGxNwEpzzEg5Z9jKbZjl
XIUXIa+gtAb9GH6rop+W5koOwRbc37NkqOZhNJ9/zCUomW21QDf8Vxd0bw7TZESv
vusThSggyBt+ZTlMY8jWGAwxBsJ3ju8acM1QpRDg3ie1vbqSvmCw/68kMDUmOrrH
SSqU5rOOxuaEkE6/Xm3NNvz/9pHqCs4W4FJa2SNLbtfMtMc1rE6xnUcnTBMups/Q
l+Au76C4IdX+eSu8aO+TG7fl+NCPD4bFHEi68bwvluPX7j9QTLp28VdKKOk82KXM
hu/lJygV/bsCBZ8XUtay5IClb4kqYJZUjr43ut9dqnKcpb87ecoo5lGti98lUv1G
4Iogvf39olUKx5MaD+1GekA0bJeHauFqkuFA/Gr0TlKQqn1TTDqvkc+juHeQRLPA
o4XCW6XOKWVlfqRYZy72sLHZPIYkeYQvTlcMk8FXGu6mvm/RL4YKSHxxgJZTXaKP
H3YKd8xFVczIZclWSZ9HGWvIS45Ty951Es3Q9aS7M+5SbY2HArQT2KRy4qR5B2T8
6LT74hxioMgB4JsfngVQFTufUhINMEsm0Mq5jhAsl1jb4Sr4cC9ILFs05nsL/SkH
bgvlr2h+crd4dQXrD32U+Ve0VL0jpff3QHTJGpE8ThD/Jr3T1wTcfRvzB6u9MySf
6AwZjflk2RQ17GgLRCkO3Jssajhpwcb5W6s1px4MDFGq6PrE+1dCN0SmZpm45se+
JJtDPNMMzFYW49Kza6ZW97wLFbNLUnKVQFNUYIHYU69mZ34IfuFhclWEtM+e7M25
c9RChNlaH+GPTmKv1fXA5gk0bO42jjj9XrFhTN1lYp1Ji7hBfx+naPrXiXXu6K12
xsTo4DkeIXre9yrIheLMFPwYCrmqtPAcWCn9mlfkvYt0FVkxf2Zx23hlf7eGz+eO
PMfxUPFBzY6rBw34/XoEjNL4CAuMrMd8NwYwi1GFXeTTw5OyV0VnoMJST4vKVV85
2miXvAqogb0lYSQj/LgjoTB3ppsapubjnGuxlIrIevK6mQivkD9Ms8ZfQMZ35/82
y8CvXAQiy19V9rJBHyTlXWTUIEjDlc/7ChOWS5wrg9fEAEb7nX0ON35w5AIOQDUe
JR02UZ2lDl9wnUHTxc19SkhRmPLtZzF06zZionjfzjcBTY6OX2eyZvq144coT8Gn
FgxBZEdghukoH87T+GZFqENj0DjJhvpf6SLtoNks/iLFIQy1a/dREUWidMVA1zYS
+E0aKsl42kVuYltk5CgKgvNlBTu9S291GPzxKy7gCcFzHP1enuxv/c46I7gijOlJ
wIo/nZpcqB/dqGfTOveFvJl3SJxKFuwKhvOFZIT9aoBRMxJElf3UK88ZnnuM0WNE
BVQi19Xjjlk+17R9s6LJfGywZrizNZ4fEBokg2iPSTKW5btY3mSDVG5CxnCACBFh
V7i2ztvzVUXUSgvC3iT9z8CsuugNM2rIgXue606HFX/qHx/s3e6ayA7FTGxGge8h
0/K+5UIjPfpc9w+osnWnwcBFNafpg1DT4fsbOq8ceM/ABn567pjBl8Bo9C2HNjuK
xOL3slILqf50MIGHsT37/zB4DA1m3Kw52to8naF9PoUOZTtR6dWYSI86J7MqOPRe
NM9vI3GnihiWYomE+WTDdXhYVNWmHSM2mW/JH1pYSUizy1Gj5QmwVLgWPvFwjtP6
W5BtvtjQY2U+hveqqhvOGDL5imYyQAPwY1F2EisY6f7kOZgdcT1bbP8ofYyRQPya
749Iz7T0jGZYwnlssGsQdi5R9aUI2fZSrrpDQach+EKMf0oo4vsbwbMod41/TJI2
uc7ph1cm4+NCVqw5b8kFZ7x5OhU6gkAR/aRUE25bfRcKhUVjMWqbI+55lGZmx4S3
6Sg2Mvx++hARePDHuWpD4cckI/jAObtNSJ7AslHyyqGruQgmcUNKyvu4NpLHu1WS
4CK1RmMD/nu6KAoOOjenaSet4Rvko8uoodtPkz5mEEfjgSFdeiBnWKjHwzUAt+V5
Oe1qVeM4noxwI3LpvnOlLQ6ag0Gl/H0UFzaXjCt3hA/2vuZge0qqN7xmOkxwudP9
Tmt1FuEB2TCnpK5tKYvffFdnWpNzbdMRW276z9tiQtNe08X2/ZGgO0FjxcgTCc/E
3q3YLP1yio+cLPYnjt6t+1BTzksIaH3jNwUDNzq7bfnRUXcAUWEzg1esCkT2ET0b
VgU4Ea9ijvGizjqxHFjMiGw3UKFfAeZOn86kcyRPr6SyqjLhtvFusrZN5u2RHfug
561Metk2+/j56GUsx33/8YF7kj7GZmDafKFsWezKk20FrC/X6VjWzCYisZKr6j63
M5fC5dZeA8+B3zTB6WWexTAJCs6y0osqGN8zwv69dwV6JyuPA6Y4aWW0m7Awt/fE
PHi0c9EG78vj7qmCt+zzqW0Bv8aBZZ6JPAr7loW2GqUaDG30pi//kbmY7LEV+kW3
FGFe89+sspjrnwVXK9GcBG39czKeyGUzVj3ZyssRUOPl8mFlKuDz1M7a3WUS6Sp/
wN4PnvTdnlfWw58e79+HpiL0mD771CDnXUb3nZyzXB1EgvkX5/vNZkjroTr2UDmM
Z1VhmqnQGc5NrRNAwgN06yX7zRgESc8rJWRoJp3MQ0pLumMEs1oNp+ANCUvhAXje
/HF8y8s5HlF3k4SnUuAtbuNJUQVzvcjbkLl/+gP/isaTfF1hh2Voaj/QYR7YcQp8
YnG6IbOnQxEdCaGu/apqP5T+JsUAh5E9U+2NjDK5+vRAHRN5E5uKr2xjQtj4TED8
nvwfFlqdUKem87gxAFWtMAnPb7FgmMcEmXlZwKhW1Vsvx8YMXvylfA0UJ0h3V9zo
ZMD13Xz20y113Yy6yiMiAKaFWRqwUz6WKrvwoz4dxPbNI8i7Y9ePZ9rI4ANW0V8B
TX0mqZry79UK+zhJteMNv/eZ0NFrwNhLt9Ros+K+ZWcAokyDiyZ7I9WtprZdyk8h
Pi3GcLYposB1ou8aEL8btRIhaJuhXMbWZNjEgkj0nU3K/vCDhf0Tiad7sn8OzfOd
SPsGCRcOHVg0jBr9vG7wWD2+HDOlxQzBQXnjfR+3me5P7OkcGYwwjSA54zjrMUQx
RYBnt2AcIhRCqXKo94XR0HLnKtOPzMYmFTUV5sgEuT/zPoE++PtRHvbxrl4GfWpu
CJ6PcWzzi5TU2BQXgA1Q91U/rvhsBKERMea5PmBs5hlB0lXbzj/vLwKWKnd5yO1s
MpSz1BVx/PqkmIrvre45FODnA+7GLQgtINZUKDxx/MIVbi8BDcH6t2jDqry+17it
bH0L3ZTM5tlsX+/2rcrVSGwQxcJIyOZHEO/rhlwsfw7Mm9ZEY4G8nR0uWFrQe91E
7mzz/NLCfOQ1t3Y77HECEoahk2wBMZYHT0KM3lxkw+pPHiFbv42LqKVB4r5qOiOO
jWaCrpDO2vUXtAw1OWrltfsy0Sclr+Up9/UBwGlgXu8Y9Q6V5m3iucJej7lNlv+R
M37WFlfVW96Xedx11cOgPWiCKZAar9qU2cLRtr9oDDUlehTO1rRDddjMaVnNN7AK
Omg9v+FUDl/HtcOv3kL6WA9P20lyQhOYxZ4r6id6VQirVoxR7oWdcIWDNG/MPdxd
ufI25bkibhwH0XbXiLlQiT72hmaLmbtEZWFFw05SvWubN0GHF/ayVcrLPPhX2cdx
X3QzOH1ZdUtXUsxDbHvG2efYOyRIsMJQrSi4GoRnKoBQWweGNLRyZtZ1XAjcBls+
dVK8vateNqKhSa5hGKEiwXJPM0HC+fAfKpqF/a52+6mbu/Go5hYj1jN20lUO22Ek
NcGCzmNasvVM/Z//Y4EFR7c9t9SUwxpx6tLOYgDBrZ2MZIIuwqZ7gJwIr7YpF7SA
eFwc6QzdzjZPsEIaN/RGawu4P4u3Zg9ZVcLpGw8ZDlDb74i8h9FJFBdUYxjsgkRX
sO6aJh+K6/3HIG4sYtYvotqPMPSoaWYbUkt0OubifrJaHIKUiG7rGOvPch6JPs9V
iae2ZxWDRAZFM+IZIo49uOerzN2F/Vx/AJANjp4gPArs6hMvOI/imbgmx4DabrjH
dSlHu0PwSuP7t6FXA/iredpKwqq9cGvoAvFPAAgt3oOlABTyphqO/GDTAcWqj1Fn
uZ7qcWUHdRNpVlEGv1XGnr4PcWVRxeOaU5Itn/fyBxD8nUz4hqHxMMyY9xS0Ct1N
SZKhJKrTZ3vVQojcABFai3k9HoDujaGr80sO0ntbOFi8YtdATYuES268N5gdzKPJ
JM1rEm8MMQDB8oIvY4NOMBRVvnUk9wdk9CXmUB/KrqIupwupH5WTmLD635USfApv
VcwYjKkxQPyhgGSMtPQEQZVSmXjTnKMxns34IpoNsqos0YF6HXbu+7wv5FKZLW4k
P0UskIrnjRJjS5F8CrelLqLxIrSI11e895frDJQ8VwnszKYXSvI1F0I1Bdt4ZPFI
g+eBCXCoPUsddoLniQ/Ihvi0lbFMu70l1CuOwvJWnKXedfwUSpjfg8QFPs90vYrY
A70NMZVnLgVbsav3oV15swDkupoO0EjkQqI3FvcEa0I=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
O7UV3y9mpBsbYf5zrH8Q/YpT+vnCbd1ZNpFDfjV1cyQLiNGFoK1kKrpnrEL9sdfa
RofLe4t4RZQpyQvzriRa++gXVja4hpGxIaAUVKTWi/o0EQ0npgyaTA5gnSijt//Q
Yo0RSmNAds8XvB3mJAlGRyVG9un/1X6uVX2PkptyeOxtSWlvt2NwS+Ui/gb74r92
FI1Nw+ao7VH0Iyfu4QR+Rd7HwU/96eiRfuURn9yh67zAwh69U9KCYK1K1hM8PXYj
9TRtvtxOZHznY1HIJbqk4YdXCHtCf8Ibx0Gx5bKPnxc9rQ9P8eGcdjzfbgUcYsNl
tXob0Qq96PGUbF0geLV8fQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 20368 )
`pragma protect data_block
fJHRZx9USb8te0RfmlmtS9CCpKUx4bUYMGQFWQx9RGLSCAsKIYUdGp6Y/NTC9ch2
FG8TTy39uXoC7r7q9Xh/X9hzzwUoHLlM0Ce2v1AqCIbfPkiD1b1onKw2+d6s+TLH
GriGrej5b6aw21ZRRQfwiJd5bIAS88Dq7uyX8QTl+m7lb4s/D2apSUiBmfL6J2TV
cw/LDii1VybizaNYu1sSdEPedeBHUUyddp7GX+61qgi0PqRyBNUcNQAYZWltEzZj
AGbMIvzcgL0GmJcKaXAuWsmmlZkDnI0a0ufbdFKJCUSkdcSRihwNd8KhBuDTz24t
L/Ee/t/iNsmPQHw5PvLnXuGJh1KBkQ/N5xjdOzl8FaIz9tPFTGKBku/zgAXgoWhy
IKkQi1Jqm05k8VdFI71r6f4OnPi3mFK0Rr2rvEqtvDhRpMq8lHxzZg27knZHsrl6
yK/S6w7JxZ01+0mGXS4BXjSyKVfBO9yI/CIOBDoAVZcK/zZVdsDIOo1Cu70HHFNd
5P6iOngGKW98m5z8+8RYuNFEMzvivJ7NFX8wamcKeg0ZQnMgN8kvQWOKLET1PEXr
4NGD/VzL0FuxB4JjTsbsPE8V+Rmrdyk9wHxt/Bco48FYu+iNEqD5OY3QK+uL6a1K
oZ4FCqIND2hLD/VKS3XtWoQXBez/3O5SPLQBFJljBQMX3Afb2EI46epyk1+qLSqo
CgeddBZBegfI5JiJf6JWjS697e9qWtFW4ef89pzUF+9nB+YZfbFYNecuvthYG44F
cWUrZeHnEWHBTv5LdrcXEBa0es0zij1cOUDakyVO7HgP1kJwLkw0KKbp/ElFApVi
FD2BuUbEt7NKWV+w8+QItecFpQRFgYTscUreGyMAKgli+XdhY4xD/Z/0jVNRGFms
TcVtCr3hfkFbhC8o791WNH8UKKGGGY/OTg62ZyjDZ3Mdx4ITybeECZcgmeo0TdEo
XthRNFSN4OhdxCk2CZ+8X/MpMXccrK6ahsvXLWPiip+CxW9Yv1JkI4WF8CIJGyL5
ZKyFBOWxaAO1UqFkNSMUgw9uHYyZHvkDa93FVWvgDKph1ohKNSJ+XXdhEl1pxBNb
/mTR9suIGkwRgHfNAuLauAXZyL2t+vcJu+g1xq9n0pGnV6X+P2AQ5EqFJg9XV4+h
MtXayJlvV7eCJU1eg3/8tdxkRUfc2H/GgmRR1Ra4nlKnHZJvi7gQYBE4KxdQRuUa
kMPpbxza5Yl2HndbMxExaI4ekGa2wFKoJiUjOE/SCc0mj+M7entcLXhmLn5jQggm
EtzE60d3aGVunLFzmPyivFj7PwmYcbKtg4Q31J+qf4Mda4FtW+ZjAtDAaVi3E5Vm
PveNjfbe0j3XhSQNuU1BoTapuORMNU29Cq7VnIUh2F1Dq8uJyVQtoJWivEjq6TqQ
blOFeSnQdsbya9QIngpHjp6+kxyZEMzLxkEqIelIV/M9sdXNLg9rvK9NvxkCUWuH
nzL9Om1/mzMeaL/ZoWFlUQqVN7YWPFpJ7SA/cIaijvyQ5Wcn7uPm04VJ7oarXj9t
ZTbUp9zbVjIJnxhC+VzZl//fQwonqp1bz06pvRIK30TI2RWffozMK4HkyWETY2Uh
5cOLvdR6vaPBVwZP+FHUGY1sFNVfKWjSRwQVq7kGs4C5YYf1PobVbYRprlPuEWSS
+5FCaLrvSNyjDSpMA4oaWtYPA4jnXSilAbyZP6OBdIVmxwFHj/PFq66BFSajUCHX
sFn0wYoZfzKdi2nPAw5HJAjGUmm3tViF5qsy+5AhFcef9LeWtrCijpEH5WzyQBLY
/yZ8ibQnQKxd1jyCSC745+MySzfgZNuG8P11QQzZEglyCr32RHyvk2sgRGT4IrPn
AqmLROuL7atcjnm5I4v/4MAvb3HTyno5aDukl64/5bMmpGI3Aw7E760fpUSd4Ju4
dG+gpJiUl272u/w5ItNvYc5OiAt47wFYAxSAE5lkUqeQMvUEIka5KFcsGgiOVAok
eulQIyGxG94mwBT86RTrO42+xTU90FmUskRehRj/ZwHutBWoCstLimchtyiV59vw
jTV4oXVkBHP0vy2XsAcJ5ttjG5UtYu23Lubt0MZFlDgfoyJ+EvNKUumLPxA50RFd
R1Fco4Re4dgPWK/qPpOJuxOKQXFd9tCkgK9m1xRiwPat4CtPJepmSXuNX3auLZwH
soGdDP9Ku70Sr1Y2tD0b24I9pvGXRhzs/cPqxdqhQ95BezMIGdsrILbarZl2s+k3
Y8ijUZRIC1mKJV5EwFSPn3ITgqyfLvQtElWX5agZ9JmVUpHBiJYhJl+ZjQ/zr1xP
rji/3uFADa5Y2V3+na6ne07HvaRhGv5mW4p6tLBhnkz+wmv6RgFSz2WAABWEaTVv
9sKSBbvk/YKfPOlAaERSaZQ9v+/NJ2x4kmFsMz3JOrFH6yYzlFdRib7CcD6o1JFo
oVH3LWSI7Aym2cZiwYqmfFS+BthPQgu1nyRQWmP5I/VhwiRR19dyJc4PHWN5Z2RD
mqW4ZnQqXW34u+nOYOKn320xs//A2F2vxIaFpqCM/D106ORlTrunnl01yDEfdn+v
RrOEXfrTIITnJgoJZEtXYah08Fb268YOmrFFgsP7UtOYHaiVdcE8B3t7Xa2mUJGo
2j35YQUqdctu+uokNtk/rRaJ2EXNjb7NpvpAU2+mZEnY1n1xPkV6ddaBNrysRt4a
UMJSaa8cDaryI65ErvalSoYpe2TkGsp4jAliowPtfGj9seVHclgHfQPoe9Fd5CRJ
zeIEXGyPrtA/E0rgryVcpRnZlj6HtMJ6595jZ+KXDzNOOANLgIM7gIf2RpABmJk9
AzvzDK9JD1/dpA3JDQ7IgB8n8ESdwmTHa5695xlafuP+uar+EEyNpvlyGa8Ojg/Q
n+JpGrFpRisF1PXfKKYe2VhJPN99/CoiuixINERGaqy4993RkUL3JTyBf01NQf9P
n0wYGjn4bMFrxpDIs7kEG6VFGZDwgqjdt5jJZN6Lv9UM9ZJXlDqIC2kTqi/GvFka
tfdxuwzkneFSkEtewemijxnHphSMbEojkh8OkEXVHcxz92uSnzVKuyrSzrAmxcHM
T8Q16/Ho+atQn6QjXRd2dmcsYwOPgxDIBQ++dqyPa4D7evAkoT32JS7WTsZgk/pK
kOfGd3MS9OYJjElTx6ot3WGF0AQOZsVreYAeBhdzHsNUMWTvvO7kXlVGZTXqpG8h
3P0tK4/ALnmBA9XIhaj+644lita5f888ldwVuyPsDlsvTwYMH2nHhzbPI6u5DsWo
6w6EOokwLbq8mDxAEeNjEtx128QBLO79h8K2RIpCbo8cBUA6fvNP5zZu9nf0wJmd
l4lpTy0VEi0dzg919Z1LqtaORGIDfy9+B0+3gwd45zWRUoc0krLU26V140FwzqS6
qo9CsCSqsTpr97GmaHhfZlBVgFQV0PdBfjS1P3Z/yWMjTSxBRHkNeSfR2LyjiThH
6qg3QmiuqH1bvW+ggkOFgdx+DMs49Rl2I7n8H07s9tjiGu7ECLw1FtENgATXYwOQ
uxZTDqEuryjl/e2jNKoDByXUsnsK1ZPjmIODsoSGELnW1wBKXbo8qFSQ2C6wAeNN
LfLTRB0C7MhPa7TW8pDNzNIxFhrnUfC96DjqJIeEzDUNsN+dxCZRWV6iVP7LS12U
4GlpRdTkx+0rNA7z+Rt40Ue6QgHGhsPr77WwU/AwexuTOJKgLIsldVwom931XKfy
7gB3KL9YMqyMHZ2YN4UsBlphnWgCCmg95mxHhV3VjOSYO/eJWYXNYH9h8ll8iZCp
//SLF98W8X9svsowOiLc3m33tHOYaVwjgQZfcly4K1xXdHX5xb157sfZOSKMm9Bd
zAGK7vTkPpNlu4VaJOzUFFHL5tnp4w5uKbytgHEmb/Cr9kTYLmaWU5EVNHvJvMo8
8MLym3AVH6g1PrCxaLaS1hhUZEW/Uw4QKiqFrgcw8mQb1meZEdZVeOVCKW8XQVkX
OyZEVksl9qloka+W2inSgESja6cepMKyC31KTE1MXfbyA2Xa4ATIy11vL0vIZsNN
/9hxpkW5t/MpEVunw43cdUN+wQdg/897MGwFziSehgnpS5SOJN4YbTDBqcF5M9ry
2+BnltgXEgc6RBynQs0e4HQ3nUzOGUFFFVZIIO4s/cQBs9rz+PUOo4By07pe37OH
xXsvaQH3EqYqSNXEvYRSDQFHYfBAmA958Ohw1+mLki9VbdpHi+hz5CkNdViJzBHP
R63vB/SXhBbPa+Yw2CyIV7IE+fJelF+V0uEobAKuL8/ex01s0C1Qrb+lhClefX5A
AeudeoSrUyQb9DWqqmtlkKliPE5+C5BQfl9DgdNXtc7H5e+ex2XCkIxfXzmKBoWA
Zf7O6lqaXzcgMu3Rgk6fQsARVYUiliaE/FjmMv3ZYcuBoVOsDo8/0AF1Vhm4Eyt7
cucgwtfYvERzDjXDo+VijiOcKu2Xu9aH/m55EGajiI5MJLye64NI5F4VKtw/qvh6
xm3c0YSFC0OAt6LUeY6GMMD0RkCSG+ICMu2a+2gbg4VM83xG3do9GfGOpE3YNxyR
P7nXptYSd1a5Z8sEhylnB5sFErDTW9EIWrbYT37LH1ZWYmU1OoPHWUPodnXOfNL9
bU3B1sgm8+cU5Ijrrk2/svcZwOFUHSl7toeSIcWfcKKD3YUG3S3haGRKRfBRwVdJ
Blt3AA+SblD2kezuEBrFJ5yjHUu2LJPorvf7UlEMDXTBz9Bya1i5VNrWZ5e8eE4X
hcHkjTy9hgZ4EKi90e+GjN3oT7A5FGH/nQj8O5TvmmKNS+9S4fyCvjyzHCkvFfHK
HMktPNIn/Uy0BBGlV4b+isAVBB+y+OvYVdEoX4dbjPfTCC7pPMr3ysQPrRaJkUbx
L5ptH9lTJ7EDQeVpCmqgKHQDl8YHJ1+vdPtL/9+o5+SJRCgwQkv3FjvLp4nim75Y
NbstBvFyD1MyVxO8oZiyar8JMQNOJlQLyS640h/A5v0HgJu5UC5LX76E/eupw7Mp
4b5GUotbENPNVlIY5MSWNQ7CWXIaV/xczYJk6dn+RtpMkeD5je+QWa5bZ42Mp52p
DOOsRL+/aLWF9v7sfQmw4Rmp8fHxYH/DIm5zW4z70t74iex0jHmS2Y9CCHVDw5H6
ZqzUhKOynjMyNHkUdv5A7I80RBVALZjNuZyc/mr2TGnUW8HqQ6AXpriCWwzQ9quP
oSkk0gik++uPS4dvp6JZLP4EHNgR3Qn9fgLRuVIuEEzVCTWa772fJQMYysHdKAPO
XoI0ttULK7l/Kn5DbOTPAPC4eYCr0ZerdnnnhlpnYkx6oQ5Qk+5PpEwOZmWe5nDf
s/4lUkr1f4m55BkKUudOxWOuAc+zj7Oz3Shpvj1HhGgJA8WhNp/RrsjDtMbCM76q
Jt9WybrdhL58vDD4ZvEPtXQbe/CrRvSX7fK1BoryY65b3eLSHEyjEWkwTVOlslbx
jT3QxEsUaNwz/4qaWUzRUI0w/jGdXQbUIF1QjOtCSrpQsLopLCBC2owwhz1lAnxR
1xqUa98aWKSuIZnB3IiTsCYfqYbvKC09flr10FbCRM3eFw4QIRc243KVdTa33N9T
/QALKowru/9pNC2J9XLbGpuUtPCXLkB8FlwvVyZtEQFZ+CAUSXiY+lVvZHw0Hn7k
uTl86bgFFU2VflXOTCSaQMOc8u9keY/LT/lrbO3UqlMLGQ+wrXUC9RcLbjEuC0pp
ORsAuVoo8UuXuNzhArlPazXeNaviu8Jh8VlrI2AwKvMd2wWWTZsqekL70klSm//0
TdEI1/8NTbTJqApxHulLPiRzAz6R/36G8ahjKH8yEOj937JjGDcrNkLNPIWdGTnT
EbFD9AL1kZ1Hqf3y9qXTmSaSnbbW4IlnQ3SfVaxCerRIm2AKdpVcK6dV5RkNbsmd
PcLOiLTMyPGuzrCjvlLD7xtXA7A2Svh207NVXYc1JidaAqfE/lZh25LuuHwyHdXN
n8kq1SsuiYIPquzGWQkYMJh8IHzwnSRr4jwgPseGOW9HbeJZCy9wWvlGMGCZnUgP
OXLWvDiOPw4J/I4thl11GPjT45jO7W4RejqaTtDAG/Fga7pvgpuQlarc/gGapKsN
MLR6cT0abhj8o5NofRfdwAECUmC3StXilw/LZhZ9JtWS6RnyIziQdXqfCsWspYrk
DrneTEKgPPJNCiDRsJQ3bnzlN+y+yhV162197KeyJjUMv/4/PuX+6JCyOzpjiax/
Q4b9WWs7qADxGaCeOWB/z2+VPJKfn9JM3JwwMWrB8l76JXPPPk/iGhY3gz1hSOpk
7G+H9v6h0Pbuz4oXCb8EceG9cX5n/ZWQnmWweHkt9yOwOHExHV5mx5BztbT6fZvX
XxPfPwYULl/BtScTmRp1fo4LROcuRjxiTwdCRGLrqUVu0JQD3qLbH97qQy5D9H8x
zYoB/lmTWT3o0aa82D4W+hocL3nEuAxw0DV9I+g28KEY/V7ATJboNZZj1cPiB+dU
nAudG+6Eg8BLr41XUT5hFB/8EMqB9f9am4o4ozu6xGBl0ivh/20h7Ng+V4BmMiD0
VNCf/yew3TgEu5MeICe5st7XLY5MENjFKSgzfJ2FUY+LLmRT6EV/L9ZrvM8kT2wQ
HInbWkFLepXsVkKfbZAYbfaze79fJgTexddqYMNZDEjtfzfOSg7fGJFhYVSccq3N
lld/alVfbH2DB2nPZLl6eqBim/PRVaOkkxV06hBly7ysmOSizbA6TyrMom1cDog8
f/++XC8718ARaA591dk2wgBBwommwja7OaBzB57AiPiqFrr12v28CG90kXpOMPGa
aJ43GU5TUmCcCy5aYheZOicelJniVPGIzkfjncpl4YwVur9/tDapuBZDj7BZhXnu
yMvO02Z+Z/Nkpk4R4whDvHZqhu9QbNALGQvnYqOSJ0gn2N/7yqZXh9AxcKgZKdic
lNvMBRuGWpsCZQoNb+uvWPqEr7Tu28P5gpkyIoHFNzmexBaaQZcHEywPMneO/wVI
mFPRicwZv3359rkZlwCXKJlU8T9v0XkxwHhhYCwuReHLoPYoFFqSsD+V/u5L3CsL
eEmre8miPSaC7EmPjcfO2OWMrF4/FhGTF0gkic9PLaUT53ysZ/cxxZGoIqx9QEbI
r+7oMcXAZuQuQX43lTbWwNwbNp6Lf+b0O/MYWhyBtoXf7y7+rQEN3a5eofZhaO1K
/a+pVVJx3EU1S83khD24wf7vDzJp5SCF05wnClJPKW2m7KWpqiRaFwszdNkeiQ38
m0l8ewIOzFe3aYNZ1ZGztZASJFK29jQpDhyQ8yYlXD5+Vx+oZHbeQ2pyI2wiio/j
P5VE2/5XFZT/5+2XPJlWZ9aZ0VcdsefXqqgEm+/oHaXgoOAvsv3SCJ7pOEWIFDNT
vIhH9pUI3G0Nt9uOi/i7IWnAWmMTIsNm8vG5009yvhQKevRIEcFEgf5p+YdgjuGB
s+Mv04mByyOdv52KeeaPPfQ/WwbojpKRLojzj/JLOH/HV8awpzwgUzNHAbw9bnmg
FOXDwLmdT96oaT52SGL8ZFVUy9uC5T4agWGZAQ501/Ua6lx6ohGhcKtIYkF+9teU
xg4bps2fj0JVn1HYtvyoF69YjvcTGxYg9jKcpNyt6PCgspUt4Wzyt7hi3VUhcNZS
57Bnx3W0fp0DANAY+Jux/D1ynczwUaU361cY1B8MAijthIbuHeiVYctfszmxcPww
ggZXZAmWXraJdQh2R6cejyHxqPkduRMdWUgUoEIXO6jwJVo3BP3sbOrD4xIIvU94
ctJ4C7HDpoySM2zDBlR7p233rR3PD9bNEHYUsmSRjboQA+zbtygsOkRriD+KxDpL
Qtjj9TfEcXYCMCfySxrUvbIXbQutAiuGGdyIZCFYC14Pa90CXP5u7R+3L+CX/gEU
XOiAUuQQzhTG6r4MlletYkAN+2Ng9C4OZvrARJHaeNrMnoWEIeMMUQo1j37UFvUF
Ks/JPqbknNt5lKX7xYQzfYacDZVPl/tKMD6ay2e7+0V1r+Me8Iknf7C2RMuoo3ol
GFCR+XvYRCawUtsUArzYPyPWOCKBhRZGI039uIOfuvutg32v/WifQ5ZU+aIf01FK
07rvmSzy7U3+u6iy+EWD54XhTjGp0KommjWodf4x9I2DgsvzfdtZCtvIE72n6DC5
sLS6fPICCFzRpVVyzXIvgJgtea0Z/OLVXmf1DD9YPG5K0EAjplsOdITEvr2FLolt
EXC6aOf47gVYJL6FmVQJ3Jg/DIVTHxDRqqsTCr01+9P6PCjhGcD8GTRYFW1PABrP
Qi+s1Izwkholowq53NKYMjYMx4wpYT0JQ7z5Z9SKALV4J7xmoYUjeyz+5vEkIk//
lrwobMCDWmTcwIzDNYgkG8eoqV5kXMjQoTr5SbJbZiU1Zh76EyXP316LN0prrWAv
PYpU0zBXIqeg/ZGYlzrSarszbS4sq/pOeYlvM1YqJUU0bkWY0xJCvJ5ojukTJ3YT
Y21BDLADjPRFgIB+tJYrM+FvkJ43FtZdrdYrWxHUBfTdOqzBE7h8SEFNfgSjY+5Z
31hJwhIAS2jyosI7251EsOA9GvnZ5kF30V0PF3eXjG4JuaKWTUc6ogEyI9yyLFEI
VMBlKgZcrSr8WMx1856Np/lEzhYSQ6hy3xTR4FLKYwYqslcls5XWqfos0ORLcHOs
fJ3dFXW+F0ekqH4j3Nzu6qpi2OQ+CrM6ozbHnWn/Ap1MW6EQrWo7BYhTGm3dmRD/
ZnVpRAbWUIJB0mNn9kf9PsYKzWMlz02buwCHgHSNO86GlNKHWpUNxu3o/JaK5YMa
23VdQhIdIgIgCmKp2FlwNVmM2OF2k3Odt7Dk7ymAQJYDHem7gZ6PWtVtSSdtMzFs
GXy8MNhFTRk65EqpS+jwx4bgTA8ltlc7gjTWO3Q+HJqTNN8DGLdMu5QySDlkmas6
NwsHzb/FUXSpbF1kHqjDDLHWNxplKW2I4GtkFYiDJV7xX/+/RgsyMu5ZzGWqBT8z
Debu8cMBcJrAiMvH56lbexdoH7m6MaAwzEAn535g/v8YLcssmlc+EBCtL1eyUiZB
YmJA+E5XBf2IT5spB/dO57JQrNBrrSj/pdOVfhia4bzh7cisThiHyJVaWB4rkIjJ
xnwWTWLPWwva6MUy/oHT1sprp8H19okmKJbTjCUhVcbJDLKwTJNPfZvcwRIrqNCn
UISM7qGe3Mznfr0OTouWbpOJTZrqLwbECgSMFRMTYL0c/MkftBpkHH4qIW1T1p16
VeRy+VK5ke1FPF1QukwwDOmGTQkE4imFVMM1qXUbkNzJ/+n/gFhYXncfI0etDgFR
4BT4cUhCli988fFNoDBIJdOZ9E8pqJFKjzQWsXHzXg5iuIHamTEGu0xxOGu3KvAv
zWS5mVyJn2gEgwlVb7/LsRBZS0ghtsHwolMfe8eRLsWjY3Rspolls/TISaDEBlBG
uDC0YgiEUubWBn7tjfNifHgqGe5vKw1NL1dkYxyI73+qcHN2b8YNoHeKaeFrGZMt
dMR9MsTBwkiF/5KauVqzfYk6Ygi7JquGnN/+kVwfTNb8PHa7nA8bFn+fFt90LCOn
Zj8WE5UNbnrFwwVGOXeHVu+MJuaYKMVblr3CRxPi/I/XbQyMhdH+RWMzhx6/arxR
jmekdC6eGIP9MQJF0cwFsjsiwq8DHi2Gt22lz5C9rbywkZDJZQ2ZEeqnZy2YLIQ9
0qXasxIRVlNzkbPY9Q7ghwUKHfYtcezpdrkXL17sC5a17VVNCyGAPzIFQEOkRO7I
9fbA3H+FgkVWcuEnYfIebkje/PNn3z0Km4/qbV9zOrc+qL+BaKrvFrvYhC1aAmTy
silBJVApeOabOuzW/Z0Yl/ch7KW4KB0zqWs+ED/h/aimXXyNzz2f4KurvH9GUhdE
fkErxhIsj2H3zEnMyQL9PCwAQltWy0q2uqnh62zYAcfTq9OFlSiE5rBja78QNPRI
U4BuZX+6ckA+jtJa63DpYwHn4We2F0o6qgVjQmf2YdV2ywyKQY67ed8KSSCnFOqA
uAM0sob0b7ojj+UW2DXaJPbze8AhXpgWGnURko9gzSEZmdjwP16yPEyz5vAnvvf4
6Pom5+t+rFSsMkdkODV5aKaO3F2gA2JPbw/4dvN/o67I/rZIUzok/0S4/FKixXUN
Zmze9mbCyyr4/rdSGadi/LXm3WBhhSLO9Eu15lShFF2O49yU2R5X6Lz5tNral889
u18EQVmJpWu9wNpJsdU47TNHAViYtzen/z5SJlgCcfTL2/tuPfNy5ert961BaEQM
SPzU10yvPhCfxNzUzUqZ04xm2lW9Lmtxrxv6QI2BAZK45K0OZi90qgGeiL9bZajg
8+12Uf8aqAR2BPuXQ1s1FH00/b2R1D+fYx4W15wjB9yY5bYC2wDXFeXwaVvzGHVe
OzF6Hr91fJHl4+8C0PfcrmNZUHwqh3+a7VlZPb7q6miQi+oCqQcaySgq271y9I2R
cB17ZImuFnVHOhZ1XL7UZ8FPfzF7KQRGbS0OLcTIuEWoeKn+jBqVbkHjZMw3GO+I
VrmczN1nj5G2iewhGsfJuZxLnIBHzGXaEtr2vUYmBlOyvtcjw37LBGOzHGZYMuWf
MWOcSnoXtUQ/4Cpv/AcAVvQULm+gx5Zm7vFzwF4KMKIaFQVjlvQ+cZFXlx9cIsZJ
PnL8GeYtnXods10ioJFeEvPdzI5GfUZIqN5rm8Fm07FvT+mtDuBiUAHO5WrkEI33
svCM0hXZ9I7H8Yws4OXJ+yYWZiC7+DNjL6f1NT98JsHE/NghFcIcTdn6U+my8Pyd
vZ6f+kWT2BAleptCIQKp4SgodPw2xQGEUC9byf34QvVPhBQufmxps3Oo65NZ3i00
LeGAAuNIuX4KnAb2W5U2pXcfcvM3XaHoZFsYOMqy9M67CrE19STi0Pg+zQt59EEQ
nUEq1gVaVT8raZ7hK8kVlekZHFZ1JzJkZsDVa9pBNt22R7W4xCjJTb0lHw062m4R
S9LWYHgiVGicAl8yg1zDl0JFJ2Xpb9vUl9ex9MrQhtfoxrYddg9AIcqs3YtDPswJ
7CoQkXnlNULHLyRHWv5FZHjYv/+urKAJSrgyeaPhxb33OI1WIrB4VLty+GP1D2DX
Edi8twgPCX+46xNilHn0vlmKSn6webRp17dR6HkXIWyhw1lA+fmgeKW0KBI3+FuH
z0loo+UARhSfXovx/PHRXeGvharptaT4PtH/xV7yh4thuu0ZBBBzh/aQY0xLwUTA
/x/sMPHEk1Y4/4i1UpIiZVpDP9ot8fJwpKRwHGMpRkaOuKSt2wF99Wvry2zRimmC
odlCnKt9SE+CHYYpfjjrVmKiAWOdHhyu06jee0EYnwofqyY9WtV5fmZztAB3MKz6
EAtNS93IeGf70SJcqbiX4JNu9vm6dC6zfIWlYi33JcLeONpHfJjtuHoDrOD38dwN
EH0IN2zu6bJHS06qZVoAhukiaTK3JfDherryjtSicguOx8vsaET0UhXcPYx3GRoH
IqNNsYYILJsaRowQfVy5670XSB8HgSSeNnAsXmzifGlf3wLfP+tgw+6sI0o6hTmP
DUqGZtoc8B4Yz9e49NajpZ8t/XcGFD7uPs5mtMh/jnd3IBA2W/C2YBC3Z4FZl6Lo
02F1SlhRTdTEIVCk0lnpENF6OR5/EZ+5SGhiN4yXJ01SnDDntuPt7J1s0WwJ/hOA
CRfiQ5C1D7gfhgjMSshCTu7jCwQKGNBRYvJwhjNfT1IqgovqkX8vLFcghH6+9e3A
XRJcyQXqPLJYmOYFQyw0K71SQ1Azmpe7y4KwzjT8xBFcxjMeo46GSDUL64167biO
oDI8Mzja+3A3Ev2KUG2BpqETUnKxAikqsBU0Vw54aJ6U+u63ugK4g1h/RObX6QJq
37JE8oBzs5HUBuE9j4W60nFigIQ0SEM6c0mNPTCmwgi2vIx9o5vHwD5XCy1O1kh5
dC2ETBOnwoSx3x6c4r/YNclanIdCUk5MZPAm+X+KDbRMxvdnbDVZ98pUDTqJfIYA
RvpoMvvVXT5R3AVteHtXzfhred4F7NE+DfnVcFScr23oAPE9CV4GIyrDGgwia+WR
/6GjcAQgZPUhi7hN8InVlLTRwK/pe7GkPJDMS4F15vj1IGileIYW8fR0UWV9yvf6
iolnSUQdmkHIHV1GLpXf+AFSXWDsQfk5bs1EwMSZ6UjlRhcZUnB3PRBu0ay6iwa0
QYUfuf97hU1WbCOX/XJAg2RME9bYZfSYTNTWfYmdrGK+Kr9uNgi5rztzEbAd1frz
cfoK8GHyHZqQwWfYVvswW/DaeK7A4Iv3vD0U51my/urKjPXUzNFzVCbbh2BmJaff
d2RKrdqAi6bQfGSu6evfgGh44t0adkVU7KsOJU+jqmDQ0HoyX4LI7CeF0VdQPi54
a74qM+Gyj68M6LXXj6rCc1bgt2qBKRyrpc6fZvB19OEva5rAd+SLzKv8YoRwdhr3
GEtBiyQmaaTLrgHzGcyN635ml9ff9IST6vMqmnXPIMPpWgIqVtnmeZYaTodxoXpM
vv0gWmzs5FFuUYQeDpDIXk2IrX0DeKO25qu+eG76ykzCyMuaQlXvKsiLEeFlJv/i
01M0ic2qqM+bvN+zS94UGK8xqmrEHvvgUj65iE6X9+oHAn1YRURvlsXsGTcE9BBW
Dkl8l/DoDlsmoKstj44te942wD/T3oNu7yhVPGU3fhm8WeCPpyaIBbeh0O+Ge2vP
GE6jqsjz716yzg8wYHjyHbN2rtO6voSd6fgxeuuOpWEmqyUo5HhnkL6zrlTzvY9n
zCE9aJ1ckc6rDGBdGzUmO0nZeCvWrh6Eu8cApxZ0RY+7BAzrc13udcKzYo78zY/k
TRH6VbcvNgZHGFtzrvcvXM/jMvxua3aNS5Jbzj/8Ymh0T1kaHOBBDhF3z7nByvyc
thas30DXXhI4nD3IdFdYasvaUdpR8gzmFvgz15utXrvIFT5iQpE9jZCXK5goZ+Az
JaweTxVU9EYDGE8RO4BpXS00dJAx2zKgpGZZL5T6IkK+Ltf51Ds+oLXLPyq2190+
2lEb2vpmc/ZNswvuptXjUikqdX2VDZPtJd2wF/I/8jv5Kh9uCpul5Af4PRNYhYeV
CgKwmf5zWSOhGqbDmVhK9aBmsuVZWbq4XttlFfj61C+3+FBKpJpxnO9+dnMtASFW
BlV20ihFbBrilTfs5MCvQrwvP1Tz+heYYPnlEFElhtKsmgqZUG2qPyDPxchRFkCb
mu9j1yHfUeleX5bCQLKLnyNQ45CMNvY0QkKVwSTsTQXAIcth3Wt5BvFNaytHJUMK
oZXTDsuVOrvxJUQ92RV8BOp/BOiuyfJ8PGd0n4h1GMu54S+hr5DIn1MJnkUsYaD8
trYZJxoKN+tyab996C+bs4yPML8tL+ZgPJpHcXG/9HUUBGtTwQzp8EBZ0Sc2zFWO
zG/0CsU6lLfQ1VmDB7cfKRAxE7C/sNx3aDQashQMbatGzFOutrjnwiMp5DjbOA0j
+oM+GUXsZx390I0BY79NpNfodw6iZAM3Su8hFFsIwFT2TLivPKcm4xTYaWtukvR9
KQ5kMkzgPshH7ievWIKMKofhjV2ku/jqWCbwUtqWqft1bUV9wE6jPh/53s2JPyXB
gwvIjIELuLRWBJ67X92o4jUYaeowut6gLhzUfLhCpjbK4lWaZ/K+4IWwKt+3HgEX
bQy+P61WvHdo2Y1QhhSiqytaY566AaTCUo4CzJkIpwXA+B1lyDxFl4d+JTv0PB/Z
tyN7xE1oyNlEniqguDcptSOWRCysea9Za/bPydRoFkOgKJ9P6MbeJHKIuBlrxGvS
kUOqxfA2XU4urW292NyUXvEtDiBkVbZr3PbWHXp8V+mUjU2HBRz6VdT1EPTnitY/
7jj9Eax2R3VCXCVH7vA9ppcTz68WBXhl+iR9Vu3JiXBeDdoPNODdWAYEM4UcVG02
gmXUDPVjozG/dSe7qNlryf0+ctSD5liF+rEXOJHpOPUhDtYF60QBWaQzS5RmVk81
kIbr6l1g0qDCOXPZEk0OZUUvOdll7a5RqIjsySrZ9bVqA39ePOvsiJYSpBVtlL0r
KpM7hbKNQ1LL4lPbNVV0/ojK+ehBGjK6MH4s95AJ/wTw1t/MOFAdCYy0wBo1A/SK
idGZ/ylW9S0g08ssojDBqabKJV7JDLEwR1qkLnZHknV1wpRS1sOMQTsznkkCXnVt
RfvFswglywrIbiO1wh4oPsWzmBtI3Ei84T9k4BDKlxcbiPfaB1xJ6Q/C1l0QN8Uo
WRgIO2bWObqJRzhQwomSDG5+qqV9a9A+Y152N0R6ac5SOgYLhucUGKnZkjatQueu
L55lKvQEBiO5lKuGOezzQ0bHUeJXFgWJeHY8mWVGIUkAeltxS6eSXxMHuOO51KJt
mrrfzfhBjt7ip5QM1/3NDd0YlKxwgu7Q4KBqx4xT6CmLQawrvbxiwy7Li1R5KE5I
lXtQTncSPPZze2ZLQHRd8gKyfc8YjdFbR1dhOKXNONoN6zFU5I87TbhmNP2CeOS9
Rak39YXfMz9NASmT4fLFWjb4wZo56Pd8C6mG9DKZmiMqxz+rs4fI2ez5lgqdbANB
+ojGdKXUC/u/iYZi4092uY0ZKlPDjt7bvOjl7O0Hsj9seGHX/GOoGJo3codl0HhM
QddxbnlGrq8yAcW9H/Y6oRpgYlsO6ealYaHFcllp8cQh5oSXcI7XOVrRLzlKOQhm
nmKFaa5rnOv+6id/wzoVYPZMqoAi/PpcFJ9HXwR0zz59AVElOkOWxHejHiF/PpfQ
6ig3MghdVaE+aLg+tOfENBRr4GuCw95LqNrkDnmUNbtAq4BbE9tb+sdb1QOfSmia
uiS3E2anaDcdTU/AP8hsvFH1o2o2xqm5BwEJbR4IAJJHLl3UCOWpMy73Rp3lTdyK
HFE0BUPUYD1UBKQINrkg+rfoCk76tJwMvYAgLcsQ5C77G1hKVXr6kMLjjEcArU8W
CDDkFwQx0tjZFSncwZSsdi+6MayjIoHYBs1hPrFLinjr+zMZTbZ0NV81apLD0kNX
7MCgAu4QGpP5VZBmnD3bZLAmstaQsY3SMIOOOLAoMyeNVtoDnH+NZqxMRIXI5f9U
Y+M1TbL3wzogmBtHnGBJRElVJM7wJBXosVDsknbyfZM3xHw+OuygLoP/lQYyNTY/
sXyUdFkvydTohLDHyxzSX0l7Mmxs1o35QJecmpb+Vu19Cv0/w+CFn3DFOgAaxGAJ
uEe1uWEBfE8WEiCtxhEDi/Eyg+TDmtYzFvV3ry4XQp/x/2liZnu3z5lF4uAYa5md
BiHyv31VrNbOAR2bZnBdh+3bGNpYY4o6JGpDhTFx71f/I0p5Xutg071qTOQmLH4m
y4RndGckh4pj3GPcPxmy1osdbF/iiNvpB7bT5h2SW/1+Dkz5LuMY0tztV4pT5T+q
VDl2PpGNRu0YTUU45lD73thkpjWtiwbPp1H9voWeJ6td6g7aMlFizpCV92dK2To6
FTyLhyymdjXwXjKkP59GlMfLYPOwmuCHmndsR362051o4oKKNNuWC7X1B6H+vCYP
XHgSrzr1qRoWD/8jNvXvMpq5veCxAtTVs3LuU0nCfgRJ5jDJjrgiJZE0ZQ2+RoiU
HY94eRS1OAhyOn72nxA0z7O8nnujDNhrarCegY98V/j2ibNc21rtv+shXZmXAIah
lfqYta2jzTP8pWDzjOeaQhxwJFB7VjvjCyofg+R1sviNwmeJN2qaH+Qwr9rpzWr6
DdhmT16O9//FjpznxGD75nAavDEQ0KjA1v2mckDAESPPVQ7pynEX8m7Txx5RmqXL
s4cTEcXBZ7/JsfxNsV7D29KfDu313qvWC6DkZlNFT9OBgPQ2Q1o8A1sDxVSU65yE
CEdjgJJqo7PxZDo1+EY6/llPQujK/BO6BrWyvbhWmrK9LFIIFXIx4pjuBKE9euPt
yoNA19vpLIOSVvdQ7gLnUcFA4N5VzdS0ltBGOVfWvJ+ukehp+kmHz+WvWYlZSt7x
1PNkfAJd/vxLmoJw2B5Ztjf6pHpiRlplDzmRtVqahcBg9/P6uNgsVw3Qd0gVOb1x
BEgFf5MDyJRcYnN2BpF93/hkkxt6rkahv4YJCWlfoMNUh1A93cvtcAmfVF4N16Yk
138q+W3bS4SZxWv+E5XMoAiX2V01WDNkvvw6dq+Zt9g+0ghWxSwE88GoJ06aIFD4
D75UimiTUurgQJH5AytmMgNQWsdirZqdvWwiGeaIhwmkbVsUZ2T3ffm5JjpsLL6P
LwfaIEyVu2Q2CdM0NfgTdgotnIX3wEBSKgOqjIjtoAWjePplIHdFCdUKycmCGCom
SpLTukrUlojS+az/lSnmk+sOnI7C5D/Ki3g/J78BVVqB68ZK56uHv9TrlzCPr3nx
i+KaEkAkC1w0ZQxcenHckhcto9GA0pEzy3bTYYXYi9bQ6g/hicA3ZklWmc1F8L3g
T3Z9bgmsTX38qKVCpEUi41mH2mOSoGrScKytNow4PM4wdrJkPGX9x12nVEkfPJdq
5o7bUj2PtMr2YfzGCZ8R5EOu+YkadReF9H47raq76Q/wJhq3WfpbmEFaa5R+f21P
Gmqplqgb107Zj2a6gvHKAJ/GD2qOHOcmsWgkRD8K7eDHqYsgQVOonvBgWFDOVZYH
KYxFKD7TC5DDmClwKQcO16ttTi2iyZFILqDZLe3A04Q2h6AN4djvKrub7s8da5t0
rcK/uRIeNWGrZVkFnA3biPiQIwkKsYbJiamCVbnr28vPJg/JHtu1vfs2rD8bosth
LT0Vhylj2+XMcQ68it25K+FMImeD8mj2R3aVSrgpw2WMhPvwHjp6ZcmWQZWogdcP
Gn7grfOX1VlYmLlm+qItX95rZE/2NyiowfHtkMf79cPHVGoOqUOOiV4XUQh+4Lhq
Syf+3XRjbXq83t/8fW5sGdMt9oYTVq3i82ndGv5ezj2cQmCI8ajjvcRpRzcqTE2C
t4WBJgLlz8+CtHAYtA7khoSJdgSQKu4w4VHQJO1eGozsWsr5sXmy7xuR7/0dejJN
hsflGzwj5jh4h1z8Q9svMDUBXs32WYB3VScUZOZ0ZiAlJp0WtAsKVM8fRLvQWvXa
nsImznL9CXCmV4ZdWeXR1ffKKCNTcArfDtzPVB1l3Vtpb2I2vcRHR1rMI1kLDjUz
MzT1wrwZmWe5VQ8wW6sRhWJRwBpdqhTuEqSBZOBfIEnDYnQFTnEl+0+/YLI2rn76
hsr2l3Q/jB0mdal1ddph7xqpFU8m2+vb2t7+uV/dPV5tNY/uU32qj/EnVrdHFdDE
LkUHwRBBWURNEOI2oR+cWp+E2p7+M5YDd4ZVDQdc30eit6PMXKm018FzWb0o+XYe
3YUMEHQ1ChagnVj86z6C4JB4nQelXylS1X7nlZc94yreDaEDs75iCvnNaJi5TZRs
2fQRxpKD2WCePHqUvgiYLatHObj7EWcHiPI6lK9IIzUDh9gs3OVnoG3RVW7119/h
QpMMbqkIpj86ATgSsHwvqvKeWoa428g4vOVUxl6b88GUG088Cj/9me4mpPcEJucY
vJhhyS7chILP+0iu3Kp+NA7JIxkgN4k6mE4hUmYiBNwnYR1wfMvVuLOyAXedd9xN
PQqmWzixLLOG4AxQy/W7VOfhrJUbxwaO6fRYS1esWiYblbfWXqe8A7q83SxLdjTh
LsIxmtF9czEmPYXHFBI5w/MSHZiqrUDRk5Jg5IskRxItLeels+Y3PIrc9doJs4Ua
F7I0pWtKzAhdVCxc1yEVvBsTU0SFCdCBan7MGPkjWGthLkAAUDZJtE5UPtrF+cDt
CQHlaCqPixkVjnA0pjNm0pf+FsNNbKqnxMfTCoD97trLdta/4qGATHh8MZ2E7xKn
OZQV8bTC9uguIsFDrexnM2l2Dg+O5ElnBk057lwiLTRM05U2JEw1P8z5kylqMTHv
4xM9HoKg1oeTsGaKVD4T6ARKbQQTI3Z7Ox2SVnpj3QFzvsAp4IprD+A9T7AH8vtF
dTdiuFYfTaHnv7YNz1JOvxNogtVu5t3l7YZJoVmuJ/GVEH82D1Ql3ne4MtsnHFxq
qOM3m3IYfOo+YTgjuhs3mEIcgSd8Yf5S62Qgrk3qnVnSu2kb0XaIiY/NZ/moTmWy
HPWkf94jwZiFF4z8nDAqnFs0MgQWIHE7vaEifJ/b3unyb1NwPa1rhEsHbl1KvBa0
uY/yiMnh6dMxamLxoj9HYhThUP/nAZcCIM5ZzGmg/2o6xxnWTp2BQfSETmHlvv0M
1QQY6DDGi2z3GK8tjiyqCuOy92xHvsqTbpJmOUs8bxQLKA9AKEwkQPYqbtlqHlAj
EnlBcEUZDAOO8c52yVf8RiubWXV08TZ/nQLDqMnx204+ueHF4GI344Ayghmz/tCW
klEU+O9CdF8UveS8NG+TCKQkmvU4IlHJwfrwQzt0dYWzpnegz1/f9POcd3OAc+N1
ffBBKoC4nRgVYuDxFttznN3gKsEqA5uvx+YwPjrZf3uFw/jApBKkQCI3o3Zc1rZ0
5nwuFbnuikBi2JdH/4rwrKhjdDlp3azmRwhhnzNOXEcegKhR8HCKbcVqrYnBNcew
gqI3qgyERYUUQLBJUTNCijIFMTGrmPE3yPhhCzryRhtl/PA+8Z56CUkEopTCPlQJ
Lg0ApMI5MLeF4jNDZyn9H3dxqQr6KLriCNCJ22iDIJFB/6Vonn6y9xUvDiQwxV0K
Ypa2GW1MWNsUa/7a1gmu0H0ssfTxOG0ShmCITuuRS/nyPixyKHtl5Dq5rbc4k2jp
cyErth/Cn/azBwxy6qPOmHNhv6KWmUaQlRSxhteeaRrSKwwDCxo4vHabXl5D+eOq
gHeldPQ6a0QnHwfDVoKS4dtnCzWzKL4/bw91VVEJ8gCzJO+4ocdnLkgYigDe9PM9
w2X75ankP8qk82dOHZTD2ApyGJ379C1xD4sOaOdWnWDmXUyOUtd5fFfdqxFPKvl5
qfXxpV6Jhrkemg4L51arpWMw/HUIUI5K+gkpmj2fcwcGcbIlK7NPlc8Z0JDO/53A
vkrEZPMaYUdzuvOxFSFBjgukPVDfSilXEVVHXPaZEwgEZgQjKCrP/Cjxuqyt3Vxo
3cZBGi5yvgpPHBlHVqxBkihlAIEH6C2U5mDrf7lh7OR1/bwo7l2Oj88L3SIWJW9Q
wLw2ugVxu5tB2rE4XxwzBLVI2YWXQpNL1dDy9g1c2wVee/B8Ws1C7jLsEcGavrPg
CEFIC0VPACvUCaK/5IFmCAoxTpHjBI4nbHwPlQYGEKL6U/f1MuQxzd75QvNmonn5
tOum9zaGOoKC32hGwuCw0t0v3T3D0hXSl3ah1oadSbvvs6YzP93FEnAlPFcW3jC8
UjoFkBZQySL1BkV0a0WcmKq2oPEmjVaJAs19gm3Rsy6Be1URAWy4BklLwyuXAmd7
fV+982C9nREElhxFUZggZdXYItIyd3bWGmP52KGmJFtjsO9dqjNUbuQSh1861Tpx
J6n/1yzVgaipf4Cxki8O3O3ZVN6/Rv54/eTn6QqABL8rDEIco5axqbcN3v2sbrK0
L+8jZViJA7gM3J8qO4L85+AjbHE5r7lB3TyLGHh7FosuT9ydIZoPeU00+XkAqdgu
ozgOC7DFNl/bFfKOgQQnVi8urNR1mf/u6On2SydDbqQnWwgpoTUM4oy35Okzp8hh
6is+d5d/g6Pdme2QvsWH0/u14jBD+GHuybl18nABSEA9kwwPt9W6yFCcQh3mrF3F
9A2F4mfkLUKLbqnrc54gh8NlSU4H7T5JbkiTlXPJV7CEihjnEBySI16t7AHsDZQs
zM0V9gU+VcFOLzuZJr5UurGtRvI4+6kgvVSbDs1xbOnpaI36D/OjJ8kgK1X5Ez5/
PtzTs+pjMe7Ra1TDlaNz3o/faFILVOZDM0xkA0+/u9IGMX6xtDdZNa9zyRNyWUz6
8G6LZ8abrG+L+mm0goZGFYlEcRf+Acj+RRpcg+CyRL/c2VJL2NZziCnGbnk5Wc5x
roLN0tNF5N0GkCGk7TYvce2ulUEXYdiQ0XrvEqNmK5BqmRkkjGEjj7F768/UJKQu
T4LUNxPhFjTxW0+7Ae7XHhJU/wUW85IabhJoPlWD1UEJ2LIwoqziSY6UxX6R2wEW
b4mIJdpxAHEkIXIwfLMwG2QpcjBOiWgglBDaIqHswgCrsmKuJarNbF/WwtWKYFhx
ptlT8Si2pxam8H+Rvf8cDRzFmamb4bBOv44wr3U/u5Nzyi1nFHDdx6YrfjcIpaYv
Ms/414y4Ts4BezVA+WA0jSa+08vbFkTjPxL1r2MdBYYqBk5ZPL7eWvfqqhgTEXxm
EyJCH4QUi5piHCNd/feiybQUqdziOaXDwAlfnFKE50XYlo6Fe3KmrVUB7s4FmSkA
6ZDHlf1tEjFU7ae/sC4h/wiodOANyk2nxOiMldjd4q03ZyaLaANuClAN2CaFVBKn
xRZ3F5IASue1U3BrHLB+yqXLOE8LPbhSsUl28AwTYVQVuCpg4E9kYSFPtti2GZX2
NLLT79jLnX4RQ94a89hIUEETs308bxuGZWyZyLR8nAAhsKdgVXXOm8YavGQwBaL5
3I0WawNKs9o2+IXdVGHSlyRPi13Q6GWpRcpUiiyYuq7QF/0J5H67EYmEmmTwOkvY
Fjc0Qf37UJdrMDrJRQmrhmT85JXXPx7qycTL0ORyJksue0hEckMl1XvcOnfWy4gT
G+P5DbgnPg/0w+zFpiFYu0w/ND5QJx6Z6soS2oL++D0mxZ9LB4meaCAJuBPY6wlm
V+z5VR3iBA8QB/ASQx4QAP/sAxaKX/vRBpJdGow51zmVpIA56TQizfouaR0erCN2
CJ6g5vxFazMEAGTRZogcdfAhTCrEi3nFy9TdVT/zQ0EWqNGek3KUdeCzbKikkfXg
XQY3rxbvcuqt6t1SRJ8CSt0Pia57Y7pDSAshjogbGyH+2yrR1mcix8E3Rki+zpz6
01c1SaTfOQxLDmSn1Uqn5nSTnt25ITDKVJnJTOAwx0w6UOABRcazXwTc+qZRUL1U
qRqheDbBs2F/Ap9cG0VwUw0FvjSj2nrVytPCMzXHbQkhrxoRmljqG//Yd33aHu3z
vc+jnjY2CoicfXWWOftTf3ufU9tKuaml0CAuenBMvHoFzbqZPZ1+g8QQWQvRJnD5
FjyPwymcz2zBRx5Mb/r5BaQUSV6MwY+MyVobtHUkDUoBp174ACJejKMUEgXl0Gbj
qj08WOpQeLNw5vbLNicLO9HL726xhnmKd87iYHHyQdsvbzyqwfEgNOE0O158rQRB
X1WLTzLdeuaFlgLDAc2YIRMUA1mSoo0qeyTQkzTyArJL90O2+iNwUMCs3x7zIcyo
iHEj6H3HxuDxFsbkROzbnow82ktSXOCuQv01N8Tm+svoqR5KFIBaBkI4eiIcR76M
oxYz+8zB4+xXpPyafO42ENDhHOMw+2pM4F9ZyI0UnwbpcE6nzD2AVA11X3vFngrP
vpYMvvrrPIC7yzqcmdBVr+fXcJ6KLIwEsWcPmLuAEWze0xLCNO05ig89Ux9J3oGz
WWax842T+GUPjKACKCDM17KvVlKlRZhL1G0z7EyYZ7eljAylQO9ZCWfuR1g+pdiy
IsAPxlDJRukLnSM4ZklBaZ2oEIBsVwDBiuzhf7XC08pbt6cTtPzB++AbLgQs2KhC
XiLJWvMOsZD9kbktibq0M8ol/qei3yfG5hOAZgYNT6rEskuP+EA8hjGcm7ciPVIM
WrSXVyQjTO2Xzg2ndsQOuz39ShzQ/Otff8OeA47SLDi4soUDHiujtMCsxBxQBXnP
msbFBbxoTJlZTl6Jjeak6KIbxeHDspuelwCxNayLAbhQrIBj03/VUFN5zcrMkkp5
nlUH2jDAZm+I92ViyjvyENjj8Y9jD3s1ligipY/D/J+87w3maUW1idxxZ7HiaUkG
o9hEoU40AucoPr3QwOU7mk4XA9YlbV5iHrs6FBq4bNaCwSPfZbRXKrqiOkZLOxgb
5Hkp8iHVtN9sXGe+FOg4/xxL6UCAg4ND4Lsq+PVsMLh6c8J0HYuvdDh3S6auCqp8
qNHbslXs8FFmlcwo6TXhY0h5V3hzzF545s7+U+vWya3y27yA0+qLuuTR+Fn4QXu7
AFqog8TSwbXtvEx4WfEmvk9kydGfLxA8/VGM4Csb0P1ZO/VE19PLJSZWots/ucGm
9T5BRN2f4pToj9QHhD29zXon39p1ZiaUVkf5sUntbBRKVV1JHs40gtZJVw/dV8wL
DJ35ctBtRcN7FMXvcZX6Pvp/vaWdXmASNwVKW8BruNaxOzi7JT3vr5oovtVNlwdR
NjQRXBBR45/MD3LHerkd5WqWFo/lBWa3wTjBCiKhHqA+QOXVzA1UxRRo5Row4Uvw
fanr8J7utnhVjDLPlpON9lfBSrOPKjrnvcnCkM9+X407kgz1ac3f3WiRHKOe/lMb
KZSXVXO4Ay2/TQC3aMHrQiXoAepQNTtn/A8z1MrMGtLLBvrFx5PuybyZTM0vE64A
+0jdxFfYn+emclApml2i/+7aiwUuqY62WEZ3tVBy4hMM2d5RR0X46RsNk1/HKN/7
/aZEBNUfIMHvYc+7xkUE3K0HOHBwlkuJYLy6MuxyJxIH4iulZLaEnVhR2IQVTFN1
0l8YtvisbTiwA04r7lerBW3CqiOFbXy986xFE+RSYmx71SxF8eZa8QWK1MKZUPbR
nx699QjHU0rWqO92XVD8KY/kXGcTV4+8Wfx37k6yQ7AwPbG/ZLF3/RhdSs032wMR
UtnuB0pvon5wnOdIojkdO3hBdKMdUejsxSLSUp1/YW2ELJzSDRSGDpKTlH4ghRt+
jl+Tqe2k+69CK/XIKWdif9IikG5f0Sc+c0Zk+PtjdhlMXd65jTrjHhAr7l4Tb9Rd
j2dFa++pV1dT19CGqdMsHoon66NgiYF2NM5OULSzRTUfztRz5TaL0tXqpQywByVe
pzPKI3E8vUBOkBA7SIYP2MqI8UvRsYngoFT8I4OpHQZphlb56qNvU6fjBcp/UmSe
sag6YjIPkaMyD5NseSvPrK+6YpX76/pvqOp3YGXlCzuezT7DrY1mRON+CNbwKSlF
kJdA+NwJKgJRM/7/0L4Sx+zba/5LJKBHvBhUiIzVIDagLWFcqK3a2ktC8o44kohG
QN+o3qlw8McF19iRmzN6O43jjzTb9jsAyPIuTEVLY9aBZJJurtZzgI7qQ06JaXKQ
uBoM0YO6kJKnT9N+bNOjMyCOdjJch2LNWKy6cLgEwSeFwNPZN6WgA9aGfhhgAlwK
LftfnKOq4GOmSvqkdEFKlloBb9Nuwuls9uYwHrmgRpO6kKoq2kAI1cCda934zy0h
p8mCO2ab4JWwR6CXRXePnsXPgwi7DtPeagZMSMOSMi+U/AQU8Ita90ZjBj/rnm4U
BlAHs0euAT0KuyuEocTOGLZ7TnImLt8z7FhVNnwpxErWRrBna5cqs47Bks9uzrHX
mstxlxham0ImnnFHiHFHcGdZeLmbYovdaMsE6UQ0vFfNTuLkhWqj+NOCTDLN68bk
Hndh15hJ+tnSdMmW4Vslje3QMF8L88KGU0/aborYoCJw8QWiwvHAW1WOTfPM8T1e
UkwWBwsIU+hZN+AHqWl5gNGmwhzCRbPe765MrXqAkRHSOXUv1SQzyM+LCdXMzWpR
vyTOy7a+m62ZeCDPrc+xNQXjwV4rTwL6nG/yN5m6AoqtJz6H/NB0E+Cuks5R12wY
pSupLXvGIycBfe855m9q8yP+wsmLkDuZsvcEOKKgXeW0SSVcuhUyf5y6NQG7z2tL
kzF3q+suJ3cMvkk3J23wN8iQIrA8KdrTA7zpI1QVeVGpChfwASTXmj0cLoJiagT1
E7daVx3AZKz84nu4feM6usPlpSao+ubHj4IgHyCo6h6yn1IMIGvAXnrjYNPi3LAS
xTv4bVhApMvMwctLSHlpV6KioiL/GE1on/9Z7y+l3LgE0Wbc4nOOV4EX5/BYOwJN
DBWIqW+RmszXc8u9iPOFFYqNRSnTG/zvt7EtAfPOcPR0E0vPKj7ZZcq49nqdZmn/
mzIy7dAGDVTy1bQUUr9gH0Pe6xnkCCIY5dkUOidFWkYKA7fTPgGFzdtPQCvfyjlN
+OkpsZI+2/HxTZwLX3rJdQCJnHZOYLfcVlTF71IH0Gc+6YYPADP3Fgy5heI8Gkkb
BV6TMxKpahy1OGy5Ui/PZjwvHfiUVWA0mP5sSTA912qm/+7ezFl2VLzpc1IdUsEC
y1b7YG+xOwjRHxIfXmORdo5uzrPPxTEj9WIt/BDJih4vrxxu7KBlp4Ivgzyi8P7u
NEveKnMQtm9nk9dHjxmWVJfMDeXjYKs32T7gaRGkcap0YMYHk/p73QRYjxfZeoHA
Li2RzDx5wfIaAtb2SfC4jb0bgncB8rAkUEDRFWsM1pg/1wkCQd4XrdH68TUl68Ic
82+p2hUDWzCgKCiKiRgx41Yt5cEeZ8pxnN7/bQqeRTMAjGXCeKbETij4nCexxstu
JcryifJ3NUmhkM9oNFtn+QYg6LgNwYZOcawCUz+IkhoiVlptNL6Mbs9fpGHu559x
c9Ag5ZQDM7PRYkIAPuhxSFdI9TxMIUVWkpYiUMlZin+jaeuR2rZvq/KvITyHwxb3
2ToD8/dPgP4CQI8Z3H0pG3wv1sNeQaAP2YltOj7xmXXldi7GgkZ6boOj0qKe2w3v
Ijk2JSCHARQ86ZJ4Gyx4+87gRGCW+1fqh47TQ+kJg1VuDFLLXHZCuGToxRHiyEb7
KjosYdAlVhDdblpJt1bxKDfHFeTcsfFCgHP26J0ZcQahSmPDmedGPffyrPKjFmev
RTwUOmYa3m7Mg2ryomnO35EfVaPQf74OabmCMct74dhMndspJxyWYlmfg/U9/0Vj
zON27oYD+y0l/siLWZONpVI71cPErCLiJ//w1R7lWXffxv15LAUuCvDA2nzxUqKl
6CyESuDruaEESnnLaW3tnKPMMaVxNXNfI05885rBhq9tMW/a5qMJdGxVgkD/CTI0
MmvMb+rLGvQg5w6E7cGRvmSLz47uKkpWxwEBT7FO2CeS2VKGGH7FD/hrpUFbDhSO
8/Be99SvOu3MfALlNfXjv/YmCq//tS7c0gm+D2JU6Zj109/7OpEbghTfF3iwG+b8
81xnrVpniZT/JlMqbhDLTUmFbtZbkf8T9UK4wmlDrk9CqgXEatgRlPwllNCmisR9
GPDz/ei0UXt+j4Lw7m8hnQ2np3Qq6WlKsMQ+ecJ5J0x2x6OJHQ+cwtdiABQfZih+
+93npm5yIvUZBNS5kjGloo549bLzJ+BFpJ0PMiGpqAKVBUx3ZcAKBtS6e7V3tQx5
HEubWp6gSGLKOdQYnf6uTsrwpSUFWqL5SF+4sG8zNtCOgdzlyMx4wz5p6BJg+Zak
6evI0kpKFbRcZa5TZWugiR8L2hae5vm4xxBTQno+cut2ggH5WIC/GUeY3gDPDv3+
Nc1j/VNvZJDsVr4CRA1jBXoe/rMuYHSsC8w7OFL8XE48bvpOnoKQM2ghpkKG3srG
ubYmQyczaJCu6keD2fBP71VkpVZmf+3AVjB2mfvFtMVrUxn5luWS2pP48I5P0afl
13h60QcthcBZEi6XVV3CFzTs1r1R6nSf/O8/jNc91ctvUQNWFZrj80qkvNGml/BI
P5uBC1CQIIix9BxWntiw6WPIFoO4duFnPWIN03zAjQKmFKpqSvQK1w4L8JalO8IN
EE/sLH5uL6Ocu/i0+MfSqlejIeFcOa56Ot/7ed1mfoVwNb/USRWFpZSmptUcH7SG
TbAaZjXhicA6KKDBJU8N7SSghpglL6zQHznjTlnhJCTrZjrrj48jkyM5mzf7X1qn
PalVAdFWV+Od58n0MJCGq39rr0hpSLL0tpq2mIjgQ6uNXTxjupcO+V1vDEnIi15u
+AJ9LtQftd4AcTGAfBtqDFRGw8OBGrKci1GTFYsFz/2Pq0jvd/utkHP7ljsDBbKc
yA8SSpL/0zWARKf5LL8YPjRb0Jps5lfcPwE1cswVxSdnltgEQr0YOMjvZdK/8fY/
9PIi0NDhNI9bS9oN8ktDC0KmE3NQSruXXXTmUeROZIOxeHf34uXX4Luexiu7Soqd
iK7x11b43p2oRoCA1LBAk3zQnJii1mNh+2/u1/HvOfgOCj2M4XnqaXj7vX66XBXB
+qniRpwDvVIcWPbGqTDbIiT+GRY5mSV7uiSNCTz/C7HrmvV69ymN6/+6uQETmu41
H/g/D0ujDawYS6eeuDsPEeTCB0Hw7MkPY6R5I/sI2+Ub4PzVSbDSKYX0G85G4Xm8
5kDOixI21KdxFPr9+XScf+VSccPxuAbQ5A4xpTL6M7uuVafwrV8EDixFUCgQasn8
3jQQWszh5cTUDDBPmPra9CyPQweiBvw29QGoOZ6sK8uZOhzt54OvqcTFnswwfdCP
KtRwAYPNtpoNbrYzzzFPK61k3JtWpVwKmmgmhAc35jJXavUQGdFLg03k3bIiAUXk
nEAJa9gqqqdFkUpBSbFrIjHrBVKl+lZGNasbcQbElD9Z1twunfWO0oNnoosOgT+1
2s6ucpnRkJ1Bbae0luboUSoBKRxMjqCWb3caGhL0x7QBzobk3sBRFxfPR/9YOOdK
j6oGwmXZtKnWnX0kCiJZB5qLWEg/uRsuOMch14CYbJNmIvJY9BUms1lHuXbraGU0
bViCJgGlqKU1hX/CIg+sy9ojKIaZmm5757v5vpqYRS2aoLRt0VxDaWgCSDpvHe91
j1GCIn+/M8ofcY6Hgfd9F5oFQ8aYEbX69HmBthZid7LNHC+dfVj0rtjdKwJNJ9i1
Aig5asuHyZXv2nkWhy2wU+P9FtI0eIUAbAnE4txkbzz6m6zMxW0BZytzqVCpXr7X
r+y+nOYogNBGgijKFjvTsqRkQuQtD1vrbifK1VZEfiFhe+p0xedSMavKkx1oQ5gM
PaOTaj2cscYGIWBwbkbWWInSmD3lCDPID+ycdKDHHY6W2Br9/Nqb/123UtdPNlVI
tgM0rSw55WarEnYlSdT3KuRswvivuUchAZzn51YGj/GWZP+LPgs8HfXjuCtaum3F
Q4euzMbIcwGxcnjIqtnyDImJo/d4tCrBcb2F3bMeSDNwKjTRsf6QHmDpNxhY/aHN
s4QHc56tNV9bMEHf/+xs7igxbuNHgl8owDOQII2FZvnmfFZlEsgc83v6019RBX4p
2I5NzyQHAU7vGbKkA4P4DzKi5l1POcCxK88zPeswuzkbH4s9gCFYAT/1tSon4vFi
02zLF6LEFhXSc4aI0tFCjA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
d0Wy4FkWvikX1Wk+aSfxhm8QOMV97HxEG8nHMCh2XHG9hMM78yuMq5ot4ZHb2S1y
4YLsolXcn1LIHMDywF7HMUG+4OKhwJheVK7rVzpwSFfIjXTIhWjFaPRMoqdriJEw
g8QcUsvp8zOgkAXwkqJO2qBzDwxztaLLGUiXfymn7Qx1/toe9sfYan/RiOkeRovC
FNQHc/Oo519Gpy2xa5A0y5hIcWbFB8vvQkI4EHQxBHXxS/yVAGwf6+duDgc9XFAi
y/SLkbygTpt75HzxfACzbnpxmAOAIlpdtPo6lqD5BpY238NQUbJ0FjvTL75eQXom
qI0vi1/qlTBuPYdnbPENmA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2016 )
`pragma protect data_block
ltRHfUDeBzPmVJh6Swb3CAuUuykppFOTv8peO6EoBHog7b9+YmdNDRVpovV2IJQh
nqv9pv/BejO1/aLWoHiaAjDVgWyEL56JRus+9tdb8H1RhpswWbJE4HmRoLcWm9OX
f+H77lXCK7xxx5Ka1xbwwNYKqDOGa7/5vgY6YnGtVIeZU5G+7w0N2NTFaufbm35C
zapHpeqHGvvIOGQKv57hFJ4HH/KIzan0aMFQunAVBuJa8ckrnRCuL4/ySjt1801x
IkHTeW2HS/YFcO4Az4waIjmWBwqUCD25E9u//nKQVRLll7GuA4ImMmQmYo9lZ5bI
MMVPGQtva9IGqt/NhTdrOEk3d/w9EOodcKM4LDiPKcUzbLtldh4qgLE1vMqC3O61
rvYWiY8yNvr2SNub/3/CSUxj25Ged2wDPkKbWRu+4vUVwoO2gGVn/Khd0F5frkxH
Pz6FS1yYDxby+ecGhFXyqMlFYeWxBucFr72545n3PYO+KMJbw18TuHCgtZfXNx+e
/ek1T9l4WTks+ITqJo+C9d0rX8SccjKD78Mx18qI56/FJF2AW2SNDHg18bRFh3pP
GMfuyY5Quumqi32EWY5n46w31+l/86OEmsbrTvhZZwfFS4GQASFd6HUxNWiFB8BF
9DJfE50mZPCTRa9ovPKOJ9eRS8fhQpiLtpnyxphYjriFLNqmrIFPYz/VnP4JIyyL
Vbht17rrIo5B4xeiK+pHL8APz3KpznzpBEiQVc79L+rUmWAdi/Qq0NX/YfbOExol
W8l/PBcCXyjdNVXy0Vxs0Fg0FXik449TIlqg7APXdApvPBHO6HoNCtDt4xebHlY3
8j3KWWL5ffiMuwzF1n75U8yhBWHdsUryfpY/Qk+Rg6RNCPKQK5N+H+KJBgvAE6SX
HWlcZqSuk4al+ZED36jhph2bNu8Ar4YRTdU8Uku5lezF8zIxsz7V7uzvUQNcF0FE
Du28e/QlfzMtMSTqW5WOd74nd9MpsAufqlajS5Zly3N7o2UkQvYrCkiBnGLTWWwU
oJcZmWyuBqOZS40WK/SFlG4H8548TYHTFKqdWQ6Czr2ioKvcAk/VdjbPf/JBenfR
wDaVJKU9B/Xs45lfwrVpSf1La1/Ci/IfcOe92yI+9RJR2S7M4myJ9QJBD6lCYv5C
y0oqCTzNaJ+PyBhySNESYIbJIPJyr1QX8SaXo+C8hFp0JZ3fpbD4K/di3u5iqK2Q
9f93DyWWX6edN1OXXdbDo5E7jIGPSTGzGTfPd2DFYOhbhVxPVYoDo0xR+EU0DGt5
oA260LMaPVX5TrmzxFBlClOjZyyoiqMqbNL8MkSsMXOUzk6o19fVBlFs739kBtIU
RG8ryoFM0WVDN951d5tvzUudlpEtgndN19h+JZxXmXZBKTkLFGaXe1rPa9tdKVHe
np8F5N5jvspQ8kdF4ltSWV9YAKDmV6n+QmjDKKOiny63K8JqjZAgF9t63SSsVrV9
RHPvS7nznqLIJeH2n+mGAogVpdXMKX8k1iqH8NKC/Iof96UjR1sAXpJJ9g6MhO4D
hQZb2Mnyhx2R7yWOfi1xlQCLTpf0LFAvxvaJEdOB0vKgEH2fdOG+vWm8pmbMPzLe
FZiAekLx7E33epyVJsmdGgOfOklfecVFtD/9UjkGrLQ7PZn4dXXMYYVydJTKWGge
55ezzKq9p4+b9hO6syKjCoLYqUg6ldieXZALgLz2k1t1dwVx+8rxS8sTqwL3hwn3
yLRGCtpjSpZy7kzq60uq78jOXKhTgC1OH2G05sSNbEJLiyd04Dz844ldEpVkPFKW
RVpPg2EZDuZ71W7FHLDMLfPxfKzcZOrREHmthA4DVijuHL0djLEliIwDb1/s6n8J
QJEK7KCGohNu5JNBHYuW6Xx7LeqPHrF5kBiMm1+0BCWwC6EJxJ32AGq2WqHmSJue
3w6iS3mxjq7LgbwgWSM/AdA07iI7aL7isMrET2MgkB5Eo3DrNqQAaCS2VJAexPHa
epQWk/nG6jsUWGYS4e4OtGJKpn9OwJAE8G+WKQj1rw840oXUjC8O4MwI9/CSZHRi
A4EfeUUHK022Y66WnLBAOoM3CdCT72P/7kf/d8K7nC9hJZiLYSGTeAWCPz4Xqiez
vvul2cB3Kg0ITQkHG4rySTnX0HyYlY8EBq81J74QN9ovoPGFyi8jt18hR8OzsBn8
E/ovcB/72VEoDDG3QRmJQ7Bq+QzUH4Lk6IZI8jpEPKIyPWHkwcEP8Pki8azgMe07
gEVfLHCysemIESfCBa77Fpgnfu8LlMSCpBcQzsvXYlJ2bluwvNimn5yROkLZ0RGu
tussugGqPOYMSFU8/AKz8yvb+rASj8DqFquXsghbbFbA20CoGUUAoUlmbNiOcUX0
Lal+vB4WeC7F0YOgABnZSJ5LUdF0Exh8RqeM47H1Y8w032LmP/LXGTX3qxY3I/6Y
jnrzZv7gU4SaA2V0GuBO2mnwtU6cpzj6mY8HjeKRBwb1XPKndC8lNUF37Y1sjhdO
10Nu7trX3CGTZYd55/Lb3Mk1NEDcairjv0y8g8fZoxsRM7oZIlpNnOl6KgihdAR2
aWLAvkkF+/sK+hZcyPOqBad5Y1De9FLFXAgj/GmzF6k/97LzgINbz7Wsdah31C1V
BtoL3N8si4nFz0tEbIeWXJrgb/bDROeCmmhFeXFtgosIBIkfrAWC4b3oBFwttVq4
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JxUNmqJ1OoK7X8qilg1daBujmD1sRvYq0XB0DaKShH+3po5imsiAXfX/FytLFfvY
ckXVH+63+aNGUF8n8ExN1I3umwmi/PXgvBAY8fNELiW5nJLRQWOACuD1780+WWiD
Zwqp5S4o24he8KU5ml3X2/wSwA1p1oWtjrHe53Cl9JBVKn+ZOVTiqT3EugWjmJlO
3ZA/TteK+3km0HCvMOuApuefakyb5I7kjAT82mp4htEUeUngU36dfSxEVo1XEZT0
3ugs3b3Eq2hmsKJUUYBuiwkMyvW2IvhnzXDQgS72/S/qIuPivJh8PaReo68MP0NY
XOvBpQSwWxb/Ny3/rwz8Vw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10976 )
`pragma protect data_block
xf7tEQ2nLENBKIdAAVQaVswO7JbmdLAK64syA8G8Zc6NVl7R+oFn9V6W2YDXP0ys
nuBUnA6ef511wbbRyj2tQeExZM4QvL08ux6CpSyTK9svl3scXTt7E8Wowt7JL/5M
EKm2Lu2mAZTv1M2ZwENri0X6YMnL3hEEO3CX2Cnu3q7VmNN3w3ikeuC7Sd9EdJvn
ATUzpeONnmvnN/YRpCL5QJi8O6DOouImbCFGNMdIBvUis+Zt/XYbhEezD1z4Jju+
o9/599K2qZU8gczH33S76gQMSVyXhbxqvN6hirVzApNxbjmwE72+C1/NcmMn3pxv
G59Gkqcw4hGrqO1dKWKwUdqzHH1KfwEiTHWVGq42TknmV1qi33O0+SxaJQdOD0BV
AYTdYekocdprdMCDeZieB7d/qySrmlyKr+/g2bD2SUfBZwNmC01QwMZR9Yf0cNsW
0YlybeCKjkL4BlXAaO8ed09ZLOmFpq3vgoKUMuddYxQYfsu+ic2cYmZTvh0D3Gma
ByCDPC6sbHvZEr3A1p5L49AzSL5JHncnt1rrMVLEjoYeP7s6tL6a8lCoSQe+OJYJ
OsEmfj3JJnI3Id8FknacYcVYiyQYdBPO9cEUcSlih795VPq9gM4z94L9spJtjk8N
zB3RUUIPHmID6BKDGkQNG142Fj6dwvvxHE61fCJ/I71QheCA1tzAfWz8ZbIFAK/d
kxnVaSaQUUmxj98thsBtESID6py39TM8tVYuD8Gh1uOE47e3RObn7F00st3vpso2
f1GJGMGVRyvX1jXQ8hyouIdgGvkJ9d8OZ51Pj5EmsMs18y1/w6wRb6ZYJzYvUF2B
KrstzCdfvysTHaXmUEy1iIigM5SL4Zz6GyOMYp8FYlGFA4DQFzkBY7r1z0xXStNS
UspJ3BWUt0uh40AD0oBtDGhnr75OnEZnO/Zhjh1WqfDzCN9m7CGStejJDFSjDq/M
s5OwcW3bV4+YLWzmpWR4YF2B6l/aYLXgCkcwQiHeTn3/JOOmYcvbJpqD6OHpXTSn
S7yDQ1+Ma2EIZ+2cFUmUkHlZl4Af0+mKDIJLugxjpmIgMQngKHZ441RR1Rc1RpwJ
JwEb3kiRl77QuyccrBAy1Ro2VPFXqqIbDwOm6jJ3h5ZryWnSpW0i8/IC4jZRO/+F
c6lKGTIrwp3C2Hg4AZTr6QaZbKA3JO7EK0lXaQeijzAOYe0JXGoeCl//admOl105
f23WvzEqq+pQ3GxI5QjbEuHIFcSKrkQ1eoI3Mfy/YRtB6ZugKyll3p5IGN1CQHTG
zIiPUSgirz975ykiVUEpS+03pq9ULaloeejK6MqvZO7kInYU/TOjeCenC0g7iFi4
cThoiAww7puutk58wF3VsFf3iKNkxsAvC5oH/kmA+yHkmr8ZYArJznKZ81m9hUh1
z1e2BQ0pzqhj3MdL4pQeJhfdZNExNDQpl4UTkyduejhjbuUGeXx0qGI15qVL2eKH
NCOD9IeV/MFYzhhBI3/ZboX/MH9wwucAPRAKnwjhf6zx8tvYV39jH5z4DvarX+QF
Cj5OEHMY8uclXOeu4GiF8pGH0tkmsVuU0Jnoh6oOZtA9GwM9IOl6dkaa6+IeWNyo
ISDFIdTCwI8TVfkmbSXEoDiwimKOAQRUyibUso1oj0BnA5DYUeP5RQirEqhctatV
xl5Jx9pvhms514kUaSQi+/VwAGBXNTei7fGnhKRBT3cL6L4rK3XJEHozhGOH36S8
UZemxjOpKGpEgigoIf0/pk6MRxd4pvOWjIJS65cuI/0QmOKpYh/pgjSD4lejsXX6
el/PLLaJu1XikZgL0sQmxO1A7Bm2Dd017+1RCgxDVW6z+x+JOHdXL/qrcmQd02Td
jnZLIOH3JWaZAKenQr4XdSZXH1ad1auxWkxX8YIu7X992J2eXgBKReovPChraTrP
nUvwG2HfkulFBuyoJfNw3eSpY2JkdKYN3y7N2vITy4nO4cvPbhN8fDjgQ2gyjL6E
Oxv9icwdxvIcG3OD5gSQX3Jp/SU0Cj7IY/kOoerUnGwmwtnSb0z/2qDtBcUqKpVw
WSGot4UvH7FvxquhpmNSQUMPvlWK7bUwAt2yfJ1IWOCQpcfvGlTMnW8vdrXAvdkT
QnyGmT8GMnvKZoWraTdrONwXijef+jrGF1Ph0Z+xvwF2LBtkk6elXKjKZhYu9Hpc
jfs09Rh9BD4Zrb44xi4TAjELMuExBY7La2rGGG1BhwwJZzns64udZlFwccxbOhaO
5yrW8f6TrRX/fIs0WnTQ4dQSC+rAL6TSICYpH6d1h0k2QukfILG6FJDIrAyZX12O
pyY0YnbCfuKFwg3dL4geBL5HfM30Ao7e+H1CIz3M3a3ynOKaLRCmfIHQWnILa+Rh
00DcHhRLOdfS95GuCdkTEDOgseVe42+SwEXz6qw2U7H73ICtF9QjSH4lImdnyn2U
I3UUzgs9IRANffX1ZX4f+YFm7viUrdyMsf2oIgueZ4dXGICjoXr5xujmIgBECl1D
10Xo/p6fs0Z8N6nL3YsuUaB7MSrJo3G2KBQ64ioAnJZqsd/9JZ7n2e7VXkgeR5VG
sF4JYSev0HhCFrQ0LO/mq6pM2kgpewDtSH+w7/3DSwMDKZHopUGBiI2JXr83Prpp
3/pGSYJYeN0TTCuQZ4ueGurihHy+exKevA0hFASrrEnx1cecCz2PAKNzCL366DOk
1Toy4dycSWG9iLf/6keuHoqqdn/gg9QxJn+JVojVX7lHbkMhqTG2QTObZr+EMDTb
QBNZ/nR+adw9ujqB8hbfzkUbJ8mbzcEhZvSyObh4TRr3ZY7Mi1VWnBTSLg1c8kNL
Mqvbk5XiVcmuiuU5m6/Pa1mjgvR2r5jA3R2OuWFkkihDwGRoUjR2hzmC9nhdlCrT
wL/QVZdiaHjm/L/U/bjh3012IeO1ZR75ccJEajTwNVfUeBpc3/fYDQjaSKUmWaoK
97ArxZ/9uLVHryPkDNVv/i4Bg5WiYmhXU3Z9b2u0tca8WgWHSGOhhOOiOUmT3wBU
esfJ885OLBdtdsQdBsuVFvwuSNG/ur6y5U7rolA8qpxA/88St4ysXMTPjV6uCMHI
NvpayMg/9FtKidQu3zE5hbDHJqp6l1RdGF4FRmKt+5AhOA/nw6x51v2gYRxt7aEL
hYW9sIwMFNKkVD/0+wxFkM8xk2nQzbvPubaa6F0AaQJ/9uXwxozkLcMYSq2tfMlH
KvKP1o+3X80/cP/0XuS4ySvVPPaCBdHntFpK/9EPCN4hD3uaJGKtpdEsbccV3Mik
PanM5IgDj5GEAOou1HaECZMBsYdbkhJmYzJJC4RejhRZ+b6jJP75U76uPe6x0tjO
NoXaEjs1xgvH2FInWK5Ur+SsbWzorOB/m66xbilaQDliNmFNMvOTK380VVkQ+lKe
J8YmowUkIfrnraRm5xS7r2nF0GzI60A3vJykHiwHzyeTlQZAJO1J6Of26rQ+EGEw
Nrtn39jcCsdSAy7+8w3aj42brwQrG7DsyFlfCx/EGGf/wWwVNtOojaO37gKiRJlI
qIOgYa6LhOieySpcj38nZKTIuiDER6FmsZ7op3eRrx/m+8+pPIfZgcwDpqgy7B2t
q3W0DKtGm1e+6h9Y1rTNRVQ6b7VxqM/j1rK4Z60fOHPiVJwwwabuEO2bxy7uyxz9
iFiDHi+oGIG14NHEBfxFjhDmfE5MxxBGyVP4fP+Rtox3UM/JT/DWA8qn8064+pPp
wvvq0e2pdH/0SRxwuA50QOirQhmc4PCVihxuvGSDb+siUMqWlauzVlxZ3AvzPhRy
Q+CJ1jF4yP6oZCsgxBlWxVnsu4ROGYf6ru00Ww28DrEEc6Zsu+ZrJx9SRDRZKlTT
ROL8PQUTpu+Wx1rkC7VkWx4HVOnCNNdpV0wZ1qVJ+2gVEIgk/ajFtAuGR8KcUWeY
9fcfnTngJfmxGHsSm9eoQOu2HrCW0n05elnmqPJRLYyn5ePSke1FJVXMnmZbqpSr
uzg7B+Ry4mYcmAKlsGNc72/ljbHfUNtY6+nY0lOCHL6NZDc46as81IA1DQZGZeAZ
lHd4TnUhE8wccjxGdumkKUy/5Jy3IpvECIh0CRwhQ67IFDiDHgBmpD8WTSNIAKdn
13RTWVW6pQGP0yifDue2fIjS+h5aDZPfh+x7DCPjoi+kvXSBW2EODbbVQtS6Gw2h
07TTed2IHhp3r0FXoRkVtoRqjPZEFNNeIekLozXfdvvjqNdnp89Sr9vLRtFPC/46
7QwRBFp5PFf3C2k3mdcJVSra24kXh1Yxc5miHbFfT1BilfO871TybKJS2gyCQOrT
Fg+vkfdpju43oQjXerw3ehRNBOGOay4qGoN+egj/AdVqVZMuElZY2kv/taE1YnC0
+pI7b20iISFAZiUrt1oXilQpVw14Hc5s80Nb++fPJdDv/CHfsqVggNts5aU1lQur
5NXhc5vXZlrbBCppjsZCGjCk9V4e5TushOTNGR+NxNcxyV+7DnBdRbbLfMlYDFom
vzoX9lR2Us6TQgzcrOABMjchXLo/OGsAB+F3Zjt8Bzgjg5Qrfa3wu/SxMN5CRAxz
hna2uatZS2Oa1N2UYNyVZ6UaNUTE/LM4dxCoMdtpRBWYk+sMPcDt3NVJDBDP5ukF
Zt4YWYUuA+oA4mnnbBXok4rzPkHDx6CBhrqXGd0yZXPiKoKzRf92cP+OATmkCjBG
3mZ6VLRGTchBYtYz+GSawZ0NDqL5SjmfDD982hcqkTFu/00bwevK2Wh1wA3TOjCJ
UMLAOu9+ZCIOBRjN0eGsb5C7bEmyiek4w3WVtCG0gtxwWcpOpWc/BQWapa2ZvIqA
bT0dPCpfzGiJ0/+eYkB2N3S6r4eHmrezcuJJOh1uZfUv61qabtRf6LtJ6a8fis8K
gVUvXQGOz2wkIBS6jNnoPEEqqbjLIObja12GvwGJxP7Eyr2l7NaT+LFsMWlv2Luv
Z9RNRy25uSzZmWKL9FO7wzgBapRbae2oGaILRG8XzFs82ulqJ34NJnsm0odLSm/O
bGt4FZEtmk/GiTqWtEL2cMC1K+P0X2Jbr6Dsqc1i3vo8Z6XJmlLJy2+Ju7NU9FCn
CpG1L1Fs3o9wxCwq4n1Ia+us4TXnWysUXA6BK5Nu1xeFHV65OgNIuvVaFdxpMQg1
B6O3yTepxuSNhp/M3hQBU1+Lwk6WRztZhitJHzDbYecpMMwoC6L/cxSWgrqRuaNN
Yi2jwOzBF9uyGJapi8xPGErQhtz+GDRmE5zV4OFReMt1yPZiKA3k1m9Qp1doIfQo
6QlQszZWNE+516hXgSi6Smp2d4T7q4jfhnoW6jMOF6kbAXktCfjEVYjqC4w3QTlS
8M7GVFFAesTpHlui70kRS0QYSMzwbqIo9r2UI+DIBbF/6p8ZwqvIPaA6IxLVLXSZ
2oSFrgB28ZWPuMGzbjczaDmmjQNskmS8DRGzCvA1aZ+pBbw53lzPzIWcD89arbLf
MhXkRjk0BmQGWX+TByoY6ojThTI0FM4VRBTQ424NTEt3donqnOzMJhBGpqxTr8jZ
osHlarGxSEOhwyK8rN0OBciyRNGAovbER9DPhGguoHwH93xXfRMPuBl+bS0EXsV9
RWOwKIgZCd+eagqOIpdO97BZX/5Eelo4Mp8sfwysYlM6OtUfZfoXB4Gs//1sQury
xGA4Ri0mJ2QWm2ks1TVL/fhIZj89v+9gJ74NL52svtA/gOxbTCs3BdXI/JmFkCAO
f45irBTPIBACJW99vMwW6Itq/+/5PbE6loEo0kgI7FmB6Qfn3YuTCPGNhzMuXu6Y
CjvcEZs6iA8dkSpy+HkIB3nz31jBXrZ0dFl+ev66obSWcHZV7nMIa4oTjK6ou5Uw
fojwAYG6Fj8XyNRsRGx6ZFNGTaliv62kq839imUM5LCOAjd2hxwP2fzLCDvUdO6x
BZO/X2ZVJj1VPgg81s+LOMP6Ae03iqT5NiXtjcmisgV4+u3uHXAM0NV9bZUWNimH
Azepa3smat1ulA1DEYvlGKLBkQoZjhyLele+yqDrSDA1ODZZhMsLyTp6DCsiHEsl
+AA3+LgLp1wJ28YIsakM1u39DMbFnlSGsM9FDPjnV3dQ69BLn0kaGZQPmWjBN2J5
/cBVR6VwtUz7UHN4+xaOWKlVbl6FJjn6AQpTykxzt9ErhhBI2VOs6DP48iwOdTiW
kKFKyhHt4xNx00XbL+uCL3ifs0awWpYw3JwSXeqKe2wS7v9qxTywJiOmb6mzc2ZF
cO4R1uhm4QuEZ0j08+Sc815FNz9tgS3juf5/P2NNUwvS/E0PoDmJ077kkpF34pP1
twiZHtQ4oeL9FqsmEKF/9GDXzPgyOrRbrvpP+sHjYVXez9WMyV1QgwYPahq4kZKT
fFm58rPwgagtElueQ7chx1MhOk5NvPEjRFHtbS6viFDIcy3J8i3n24myooyyWeom
a+C+BdWbsXKY4nGCiDsmq7FbBcO+Ao9M1X+K8AAp2cc8P/2VcEclOaU2k5lyhUFR
eZD2OCdRvLMjuJ3cyPEs8QXaNPek+NFBP+rPUjCbYXLDVAIjqqymB3Fj0uxuiRvl
mSQz49t8AbErU3bCnm24tZhVJYQN4Adq3H6Ieby8vNWXDjlMDChIg1L9vC4FAnME
MQlQ1TiKfSwz5PsM0VJNf2Q+tO/NFsjer0S5XUqKy1l11QIOxcWOmM2slyuCiz71
49J4gjzf6io3id4FNNHPqULL1FFRaOsefabXW3dPL02vJVvA2/qD8P1XFx42v9ui
3QYnBbLLirgHcZTEcll9U9upcPO3PKNrVIM7zSJhpunf24LyB1A2AEaCqf4Jr2Ph
q+4J+Lmc9PGtSOEm4pKxq582OdW+R7EyYMjFi6yrtkGMSlEQNjM6qAQFvdnwiUuB
VdQnv6N9G4uXOHOYw+G+DBNvYRAw7Ag2lru8Xt4BR0yeANm8tEhEI5LElOrbN4S6
dT3f2foRo2XBCs1n8lLlqtGDaNczkpHiKjTm1S5GVJba5pKtUQ7ufa2i5LvXum5z
UTo3ASi0G0cJ5ub10lrQJZrk03NaIjV8cbnU5HLFtcmfLj6ikUWWRco/l8jV9OXN
G04xPf8aqLqH1GItHBC9pCfzCmc9nUkkgRzZxT45a1HcwIi90nK2fe08GqnIV3YW
P/kkcIlZvgoeuTzQ/7uWgCaI6ozl51qbV8HGHSTOpXvY5W95tazILD8jd+jKaua3
S75nDqbRaOOVCMto9fBSpSQoDkNnYgiU0+8evXIRQiAaJLR3Jjz65Iu7LUAVethw
FsJvz+WxHPhrXmJ02O72BE5bvZTlxWLjbdo3w3jJfJB1ggjCN6N6OttrZTN0pcJ/
LNO+4/Yfxz2H9Ir6NGdgtOBRt74KreU2fh45gWFe8Rvs8UjcTTi5l/iDS3R7psXj
oy/Hl7S8jJsjyxMDc4JZdsfbxMCe+WZ1y9EfxTWb8VY3ZyPQ9jAtaV7VwY/0+UIF
7Pw4I6vAtI7MQluFP5YFLUTO9/k+sl8w1naN79x2q3LY7t+cH3dXHtfN6VOqCWLu
W3x7Wpc5dWpQsMkmp1VO99zq7lk8XpWgdIjtRDfYTtVkzT7en/dH5+BAufKNv07l
j986y0ykRGo0tqYqsRo3/sqmHd/LnMyB38qCy4Nh9Ckflf8QOKwzo/FKEi4sDljv
yTOwiptOCbJAgVRcbWhMo/wrS+E03EvnlaZC/YmteUvUY6eJ+0j8v49s2NIheVOM
xC7xM0ofpuA9VaEONh3i6ORAC+iP4ftsjsH1ttRp1/QV4wHwL6SM4db71p/YyAqK
J0yY2JS61NRmfnwnkrSeq3ZF0aYgMNBbRZkIXCvRzmFkbhekGshRFtviz6++grsZ
3FtdP5LYEyW1V4nHD3PTIq7k7q08AI1Z2faOVU63C35Y2ripA91//YSzGShzF1Yp
dCAPjMegMDAtzCaTy9IT1xNUode7rYhiORz5PCl7Vr6EWI10uSqmFQVssZNYJEKe
M2UJffT8QsAB2SJBnLSGdhbj8MPa+tsIHtXhYZQ9tiEqZnYRlna8bWkk3Xcp9x/f
BIDwXgnQE8e0uOUXCkmH1kYNeWKhT+qum8Bgd6SEXU9UroK2TaWP32wDtEZEEf66
TzOEZAHz1PlnnqGqw4ouax/Tp1c+UhkpTlIzcCjNT+BEJ+byFjOIfzFTKOuxVpUa
LjlPg2FwX9Fj2x4tsPxZ87M5554sOsJuaFeXo08iTvsvI7Z3iaDnXWfUbTwIqE+8
zpAFFtRrMowIxxfgbraJ6yq48mGM/bcv3w6h+itM+Pg993CxBDup83z3SUDETKa2
M9DM7Pe0NY5oUodQ7BT5vFUZHu5I+ofORk41FXRFM81Pff7Szq3FrQt2l6e4QObO
Qbzvzb5feGJro/YH2LWGRMhGVyWbRA2uuwOo1piMHQD6fVG8ZU+IyUoXSuv0PfD9
CXdsl22Sbvr/P96mNBK7dDhCYAqaAWzX2vSEAxfA4rJV5PPi4piPdjAs8H7kM0Wt
G5mOhA7Ke6G5ZIlX6QdhpjsjgGpjTYy9aJLCVKehofdoPhnNr/B4vJLWDY1o9ZyD
ekd4X8HqGTsHqBokI9g/WwPy6uxsPBxhygrT/RcNj9dgqigEF8zGrk9fh37mLIkp
4jH6X/0yLum4ELGsNvHpWEPu2SEJQzEVGXUpSWo++TflyknO8kwH/fjK0y7kdET4
kWKaSUy9Kq9Xxpb54tialGTdAJLNIpBDQz3RypAqkgk2hgyMzp2vEqpTyfGugacF
uCsj9qd5u+M0hZpVW7byEY/sYHUM17jg0C8voddBA5Ux0rJPFk6zCboVGVzDcCFo
phUJwr7DEPHmCLCNZps1ksK6t3d4g9jSv4cAxrkBt3mYTp1IFHiCEzObCMmj3MVF
ae0/Sqs7LSCRVSPJ/PJJKQKLYoFMxguFGp9dl2Inmf4aBoyBYKCOwBOzkTOOjlw4
DkmoTIrUljPat9xfBEdV8prbF9z/K+50p7Hl1Cy49ehlZbWQRLPEf5DNSS3Kyd8h
ikEUvBx4yBs0FxykCSVtwexKlGFa9vnyoLguQkiubdHv+PzDuMc2hFKZUI6Pc2lU
Fz62SBuSd6xs71x74JrJ68Xbw8pjAkhxZJFbOUeoBaH9oPsEZnCavBHEUtPL+4ei
kb2coyIeryw3WLwyKCX4R9wRRv6+rfx5fay3QKzR1MSIhLcAaR7AJbtoVWWS5/kr
a4+PAJna05FKhiEE8dI2O/fh1oF4zLn3MMl80rjZwnoPPyn4nlutZW0JEhbbJajy
1MeXdSEpiG1ICDR1V1nbgoAJYfr4i+QdpiTaTTp50DxXyGSye40auz/Ydp82vU4p
mj4+0i7gHuBLz5YmF9j6MgQYmQr0d82oz/qGyi4ohgCM63Qz7mQSLltM5BdjEgGF
qKeX31D3kDCntVpbajnolGoaZ23iLJcYOP5o3My0VMV0eq5UWlUU4ThyeXffOfmx
sEH64Frbwk2xgOGT7TqQRK08IQrnR8M+W3rl5rURjJInZTtOLL4qSk+vNySNjbDt
jbXiwlqtZh3oPw49asng1x0qitZWMC72zXyq33X/VWXakuyml2LcrZTvLc7LgjXZ
1pVrPTpTD4JfFCfx2yVqiAW3HNEvJCuMyUl8XUjkPCRh6Lpx6Y/bgiZLMnOoKXNT
MhiG7Z3OA748h0IeImD2qrMFEEn04vgH0A1VsCOSLxtCbeyocD92oxFa2NrfEB2L
gvimFH3JF3tv0RgwKA2/UJWxesEC2d7HWakOMASKN+c663gR3Q6LM+11hRxzYR6u
Yi2Ly6gNlstQEvFQYzuSKHxhteCu3RDsvwmnVVi4Qo+XilyM80ktvagZR5VJANxK
fXk2MxmEDSoG642Sj0zaVPX2yCaWE0rxpzNtGxSP0zsE+SgJ1mgYJqqDzyKTpvN8
0qK0XzjeuUdkSA2eP/j/CnwvxlIKMA3gy720xB+RFpirr20V8raz5XHqjxunEjlS
6jZiPpekN5Xu5jzlwbFA0GFdWqeSpT7+fhMHqc61GIq0aZ9Zb/cJAg56IhQGehQy
RBRfl/UygC1iPNQ/86Dfe2B5scIGPR5jZgpbcCaephsVIYh4h/kJKbp8se0e7XgS
oWbnBlNgAzIrYezB+3M+f49wK9OwKuE7aG5c+ZVAW7IlzRZC+45t4bPZkf8qkU+q
AgmRMnZdEpTTz83GhlPR5E1fG9EMFepkyQ2auXzTVeKEm//oQvhs3G5gnTEfp8Uy
jERhj1JNfjyeLfJB42Onuf7b/HgLtkBm1acReWu1+xJd57NsEz+bvgTm8tCy4KyR
Dr0getZvpJh+Ia0B9fWoDHEPoTCyjDHrkWBTENvlkCJMDpt8+BXVNvw+7U+KP6z1
Zx88qE6i5gSItk53MDRJNuik3aq0CLqmZnpdkPKYeUsLieRt3202MLrRsm3J731m
DkjI8PPJZYjpqfFDGaTo7enZNm2oUK6OqaD9gpGeuz5yOfKTiZzstNGSSG0Kh7nJ
3NOAd30EpQxuDQG6cGeDWG3+Z42UrU9A5v2pSQlmLjNDwGz6dtbWCqL/YbtAPeZC
3EEW4rXMvcVDWkknmu9P1RmY3wwgPKKAFlNzBTpVeU6+j4RGRco0UEv6FSJniGak
vLQqZsHP0VZZOPifL5ix+ZqI3ncZ8jWHfYpqlkl2dvGKMQJYScd51qch7fh0hBzV
zwbF6a1FKw9ZhZuQkw6S+9PegCPNE1WpCxqg2q6PQXBCmoggIhEOySrhlNzkRrFr
tXkAGEWgaGhpYIDKOrFTvCvQC0dRj0IO10E5/4jQfxhscmn2oZs0FOhOkn5ZJrhz
B29xtfs6H3RgOg/H1CUr4xkoTXhsOgrCgX4OS6H89Dq4G/XSRTVdO9RculjkFVZF
lhQitNPz6oooxC0WjL4AmAadp85bj7srGoA/7umJM1S+sRi19PNAF9FtyGZypKB9
78BVFMDM3WeFUtKWdcjZEbf/ZFjy1+MHE0tQQ9Umybf1WOLYZgPZh2pDjtEo+k+j
W4SJBeOHIrrf1wrpcF3fLMQb4YHCd6AR3cJSFUd3A90ejOYxg0s7ybP/Hz/2UuKG
hDyGqBUn4FKPDWqZJlAymUqgtBlpfqj1R6nEFySlKBF8RP/flzcxcVV6eFXH5yOU
wILhUk36t31Copps/rDpUigVLGBRRfrdUsn472QaD5vH3XT7ixXd3sFWG9Ej/6Fu
VJgxN9sOB6n2den5SUvuMoN3mQvzaB+/G1avatCd72KtArbRS2CT/ztCvjKsAK9/
5r4/O/ROUkPrPFMWutEnTu/aaWB0A4YOncQwpuseRHnhVdKZRKhXJolAeslTG6M4
119vufrEKfOHjKPJkdZUcpZgmr9E8kMPYbWEdY4LMJhShcMMealJWXSvAVm0Sifk
jflzlGxO0FdDnO43VPvlZxTlsmIObZh7dvm+Ei0Fz9v3fCj+9f31K4i1+DfC3bk6
YDCvnswVadCNnZEGBJ9UmtAjQrNROJO5dSoymsmS4mqYfXe8b49FDBh+jmftz8i3
wBJQC3DN6P+7ZysN2bbAUJyKeVm0mfhJDFq/IayFm9TJG83vfPjto/Svti/uC9Re
85VrglxX8jBbTSch/tdHRAhLRJbxFe6Y+v+H3lwfjEa4SEwKL1m88iRT+1xRQ5Ju
zxclBsVdmktMuySKBpjfYYhziRGdSvcMe2/ClEoPLb9oaYZEkBj816EQandRjn9w
kDgZCtpK+G9egSFg6tmmjgdWpn/kRxWvJkFqcvfAQzAtwJVHDNKprRh6tGZ8+9Xx
4mypdxnnSbUnfkap8eA9HAU4n0gVPOFl3MRU3BcSMtdHW2PAP/treOmMDoD3yhQT
YeB3koSIeZNYY7UciUbFzRKx82hTpAWsEBg1kJmNO3o/hQBOw1heX8zwXULS8U3z
rT4Bwn4a35Hvk4EPBllCxvi/QOpNNKPP1aDtnxImA2STaWwQPhDRt721F/uHabEI
w5ALJdFG0gDlmlwPp8KtS+rafnP0edbscxPmuN41ORkm+x4HNztB4GEPHVEN+rvs
FI1tTZEMlwnu5ab5gq1tOi8SOzkbMUaQZgv2N0eZyzlbPZjcM52gPg7TyNU2Yy5m
2IdNbcVCGJkbD7rrVTKv3U9MGFh1c4al1U8xg53VKSTr45FAkZDiPp2oUmDJUDRs
h/0/Rzy4sfNrIbu5wXkUjfGd1Q91TPTGlngrMo8MDinipq8fEyRLwdj0l84tdXqN
a6+f2BR3boZrePGvZajaIQg3UV1D7xbuMaJW3fUp8ZpxLNQ9WZg18BrF7BGRxPdB
jU8tD0p3dkxQZ//YEYqhHDxj7Gr1du9+RPO3LKwHbmkb0720PZ2g6lzYtHLcjP0U
PkodfGflMzI25E/QkwJCKZddjnSa7nTM1B1Ie2pFkinTIMybVBGTMLPhnG5pD2as
P/z90NVpi9lpWzC3nfF3aw+R/bl4tDPIMhztu6afZCpU5vs+wmK8rzIuTX+d1+e9
1T1TvnVQJZLjQ7SKAIO1kgVYw1GV0Psu4GQWTxei/j8VYSnBwBrAxw1NfyjNfJEM
+Tf8ArQBRk12H7kvKksczWrPhaG0Eo9xLcDxOEQPRgvXo6gIHOz43VFgCtH86s63
n8RCrqR+Ad4rdeUDOqCmKZQ3soSG3zeXTKz6N6bQSNh5iyEJseuKsTfQoHUprH5T
uBPtdf98MKDQmZ/8pZs5EfFQDEAsubpjgmtPDQ3S6PWXz69B3cXMgYm7ByAPJFXN
h3vn5pD4QdDBBj+tgTt3MM+Y9x0hW+j9QreiwtV7OqvDMBW6rrVS5UVpOxZiEbUN
DQdkw0OvF714Lv1Sg8rUpP/m6FQS0wQjXanCVqXsIeH1W6UsB5J3il4FofrEPni0
vpdnDrrBwC54EAvPdnPt7u01uOoNgcm7jJXJB0tBfYfeojW0MagIJ/YTkXPdn88H
IyOJSPt5UH522EKrbHalPM5v5cui5YfXha2Vo/5AwCPpRPgtJOei8KmMDbQ9SA4h
gSg4Lxe5emhjVlZFJMTc7PQR5wtvzd/4tnLMRJce+UCDmUX/4Dopzf9ArrVcly5m
y236NgyyNcKBP1IcEjwKT7Twz4q081b6G+G5q725M06DOqTbT4k6o+IPUZVPAagX
QUjcc/cOUg4i/44kykA4h3YI+Hk0iWkS8lPbG8Wtq9rEmcJCWlXDkNrq72s1xxPf
zlx7Vbi4NICKFdTikBN+S69mdKn9WGlmZus7YlzSG2kQTWGEG0HyO+woftBAPfMh
Vab3Ph0VLs8ACf9bvKDvxZVhwKZ7KKAwEU1Y2rFx+nhShvhSSfNtSpt712a+Axwq
q7u2yCOZENjnr64hsYVbmLst/ZLC+5t69bh9WGwZJ3gLlnKKUpFjkuBhQdNr+MyU
zs62vOEx4qOJxrWBTnOzkCuOY+PDN11p3V0SJMcO/tg4cNyIqimhxlP2CvQmfvtm
iDqd0mactypcBPTdB62AmvWUjJbX61v3JEsV89RCLOMY/owWX1GOxBb7M8+xPkKj
6YmRCMHLDwRNBHi/QFl550vc6tMiJkGa4qH16zvT9RgJtt1FheY4aXxTfpiY8vru
VZpZCCSGCee9gmBysNdUEPHEZkZLZn2PLBaPedj++JtUzyR4cevQ39/0XzATpwDY
KiPCEZP5bemK81tsLNffFgBvT10wY/VbrSA3xxUQXe9ifL4P6NZuoVGrB0zf7yEz
Bj35icJRuPg1Ofs+YpS1OBN3tYx8PhU/jHG0SR3BsAx5UBuuQIZox0Jvt+anq+pm
pnkInZRUf5oCrpZN8Tp7mC7g/vNHW8nXq2aADSJw6XHsEpivf9pjpuRbTc3yiJhS
UMbjUFqHubk2YKcoKWIwDOabtbKLcVxGtCopUl21rmJIMpM1iLYbrjWGw0T8GNY4
arEypXn9pWokMwSTecBlG0EXzvGnNq4D4Lh/5WNRUtp5vBpRR/a/CP5OyGnSrc/H
Mjr2F1aHFsBIKEuuZilrpiRpSJOjK3O5EBE8Og3maCWEjwvyMhaxLgGdEEkZIVpR
TYWAJONZLPYdfuWe2FSGHDfLh4JihAze30z7hFBPaHs84H1UPlu1xsx6X3rqcvrY
fRd/aI0uB1ChHyYgd4zvqYswItoKnAKQqG18tSnz2VE5F5tlzZ3aqSIf/weIVsBO
QVGEPFU9vY0Oho3p9jWtNl9yUhNM2PKmhN1YOC3FEpZ0NYF3E9d9OrSR1w0/1qzN
EL3F6O6yTG/iQrtTbC1HRi6qmXy3blVk9WVSoOTWIQ+iNj+Te0S8djTen6YJlyVT
HbpgzY6SHNEyejWVTN7WK02CsAUFypI9N/yDURTFQoHu6B5h/HD9M/v+g5qdEoxH
enBP7CAkVD42KNztuiBsyi35Mu/BQzrQkh0OSpH73YN7Z2L1r8B1ePztHyc7coLY
o8FGhg/5ZMUlQxzR0oQTXztM44fss4f5nz+ALiHUh9356C4xKOopTC/payud+P33
jTmt7EsDDjjrRujQ/lWCmWEJ/KUZUNsqJPMJ51Y4xc8lFBzyWiOi9mH9WgphMr8R
Xi+c54ErXyDO+FDbRLejNocWrySIEHsOzv+28KN+2cAqTPmoPa1Kimu7KHvIG6RC
bebFVEa5VkfRdQx0SGnQWhGLUfo1LZ33JQVmpKIVI3Ce/rbIJ56PnAWniI3541su
BOsqOo8cZBt+wtTk1YhjWl4Ikl/urjE83r1MNaXLdB0=
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nE1ucIAEyzT6YyvyLRDYjIDin+/mLqK3ZgQ8stDhB3ouCKWMtPo7guUfEPf6LPD6
OPCtbLVYBakquaW5izCYMoKuWn84qXdCzRB+Pp08TP/vOV5uhWE4IgWyxrg4KU7g
Efosz9gu70A+brUBkJjooR5NLOAOZf208uPWq77HWott8ktFnH3yvuKTN7igO0XY
LTma6xQSoUJw+F3oV4OGg3Fqq7eFx0snYlsWN6lCdq8mLlNbksXSB6lxcVIVeVFo
L/gampJ8OI9fT6O8NbpdGslFkvG2PEjnvpCR76r6Y20E50JlBjqMhCSzBnFmx4lQ
rAXSd8BnpUYvfrqhwo10hw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5040 )
`pragma protect data_block
WiTV8h/1MxPhdP6dJnoJGlMXFA1JExEOPQNcj1S9Ib1WfwJ/LmfX/v693vKKdGiw
Q6Hj4d2yeIKml/f3TOAFMxDRLJV+XfQdGOc9ihMPW3muuscnLPcIJ+Fuzoq417wu
LTovbVDd7odSqmDVXUQuF6QRstHs/XoN2E3Lz85+9LKbx1IcZbs7f/7VXEechfne
e7mfqDudnN+7Y92IbiKFbTxR17otTeWmZffo68AfNF1wEAdDUQFYEsrP5aJqqyH0
Lecl6IukLM7aBjrm2panIe7I54+Vz14TCSV9VQws3VfxMcKwTeqI512ywAl3X/SL
0Fjr/Tqd6ekLtv+ISw0emaStLdX5Xl+sQmRWnuxXOiNujZkXRHqch7Tlnev/m1jn
wxphaGb4zq2nHIXFhuCCDLDBsRxrOOrRaredehSyIvPXVHRj9IxR30oBkS8tOENd
TVpu78V+NSTMKOLuzJRYOJFc8iPpESZWX4Tlgrj1SdcuUCEjX/rSqlWV5p9YQ94M
+Yr5YGxg6ZaXW9IL65Dn1reknQ7VtdbG9nAdohCfW9X8OPKqzQMBnGjdS1yHPrcf
hMKF2g/zd6IJcUF857/CHM/iRuxUnnN84eObW2O6buEA0kP/yNXG/Z8gxyGzopeA
ao3e2+y36cBs0gcdoV5qCH20GJ/IBhQDWO/dNSHH9a9tkuoixYeRPiO81DNIXrpx
cmiR2ktUBdSzJasuoo7VPWwz3PPA/FwmDus0BlkEF7fnHPngBytM0HFalt3SAcJD
lrhkJYRfnrDKymn4DUKcxCEU1KvvpXTInmq9FB1A+joccSqNqUa/u3DeUOZf2iax
kebhzG6+KMmWSVOu3jHB9MtOwkmay82jRmvPY/6cSmJqVTJJCzAJYIHl9u21zDSu
vKELsPfBaSPV0KRI8vC/8A9zfcIeeB31WEGWPb7ZWXoIEQ6ZehVn7V8Elb2Bq6un
G8l/gQf3Hi5L+2nNqWSBUjaSuM8ffBBRcuuMcxp9Qj8o4gwJYuj6iPk41Jw40Ric
OkasswtjKkorYlWKt8O4wKoR0P7JSfgJI+x4/cYbZGZm6Hb45Cvo6xhXRzxtXfOE
FR4sV/sFxJHKu6rOcqDBtFZPmlnsjsCP2T0QEQtp+TI1f7ygPllfAh4WJRw4AdTm
26L8WbPA4NLy728xWqj0cQQiONHzEX32y3W5Z+Pfty0zbGC+xtWZUrj71dXw/82X
hlJnxvNh6vQtp6Nh8ZzzIQ4jxbppdQjZ9uSJKwxxiXMWE7kQkds09Yym/7kRibqa
mLbhekiTwqRQok0x1N+Ehz8RcrOoc1qkPQNlKwToZ7fMp7zqu73mSnn7jzvQnxJa
YUHZs30f5Qw28hKQFB8no4aV+rZykVekPGu+RcZsHJ3g5sJ7Ny88mzeaX+qCqoNW
SiYrDBoUnVH3Zkcv1BY6qdp3o6lI8E70Ihva47IDmiBaB8+T9Z0wyFA4yKlly+FS
98taeooLwi/8ScuGBelAZxi94wXj/PbKcoOT4jSFCQD06SMPi+uh1yBW2x3tqVwj
czIZ2L541YX/bBZyIB/mmxu4fCQV5Xe5tPaB4JcnnVLnhqndtuP9N4VC29iefZfX
v/ZPiECwtbdMswKm1/b7aJP60FPq0TH6Rvsyyvu1yD4LJOz6aKuRqZAElzzPNKG6
GxaFTHwFCeHlhp4rdP1hITKCdTFLdJ1iWUD7sh/HNqb4u4aBeJMxFMcMOGeQ0LdJ
+TgtXjjN2WHSaWKV1yPUA6YetwTLH6u0c9JKDsF8X3YMDWT/KvRFdVZxLQrzyVX9
9RKOwk8tYfmaGaLtyIPezkS19neiT7KjXanU50ldDWzBwzmxEkchOjdhchErq5IJ
YLeIA2gQZnIwdv7wvJwVJbOTbfGhlGirUc+r6JX3oq3GCwuaEWHxBMoRgf5F+bYl
TkSBYZDQgeF1L8tdodDJTQZX6oyErR7E3nkWvvI7Q64kqoZflPJksJxZZrsIHPrn
K8uRtWZuXrlU346jy4ghvUL9qNvxk/UIa6FvJ38DKVwqwT1JiQ4BHuLwXFz+Bq5d
rPzplS8GvAdsJUuVWLxpHoyA4wCLKZC8u22qE3tg7eSoAFbJcBKgWPK8SuUlDH04
mOXxAz7hi3dzbUOaHzwYUK9UHqjxcjRx5S6p9cLi21maUc+Ns1SwA+fLA9hgOnWM
KNBFNx6G5ezaYdN9PhfDFbgjAaMEI0T68ow0GaMPwJjkiZ5JSPhWPbflyc+D06oM
3UftKdbiUNHvJrMEUtKd6CHmSNE9sYxeOu+M7E1Fos0QzbiEWPIThk6jz/LsSujQ
jGlfmDfUTOy0dNUxZ6diZY7M62FK1bHWSHZ49TcXUp5M22HjL89ANhg06EZML7Bx
E8lHdUyqJJ7c2/kPqCq1y5GccoAbRCN0lHO9sRK+CgndCA8irkln8Lj8D9bECucR
TggFh0AXjyq4bovdpSbLu0EhCtBJ8tnWcadkrSDyBaR+kw0acIQuYHvyqk0+VytQ
i2tS8K5DPL6HV7zU3+Q5nTbv1GBO/5bfN2XHgokX83iNSoStQTUpkGBKHDXvSABn
FqEy2/8jKipasomVn4yqgf9mnRti+Iyp1sfYIB2KpD7yC5VO4muWsah6clKHENBM
w7sgNN1/9/V/dI3MQHiN9/59A/74bcoFFARaCwap6Y4brRWl0fQScFBO5aMSML4v
zIR67MIhgx+DI5lqG7ky9YuIVtgHjRa1v2toKdoglmgxRbd00+vw/tYm7GmDz6g/
no3e+R8zd4RDwqDqS/YKHiwcerQaiVysrSpugkTlM4zKpFiiLd7/XyN5dexCAb48
7Ka3ke35vaisWVOO8DIBPFuSNbr009XERMnKz+YQN4jU4F49rzD23tTYG14ukySc
o77RzNmqmdQA3TBblXQApahP2T6WV6AsGWv16SFut+hCLHZFLG6/76JANxKVNBD1
zZVqx9PyHcnExMYdb3TsPQpJF4FhJp0MlLoZ9ZKx1z0xXpKxu20FlnKlMLG15NNw
2rzTcMjFEhIS0kbN8UgaWgV0OxdxyrMkDYRlSzANHiA9GdEL84/88xi2qRk4D2SR
/FGVWsuhlyKK8hVIm6X/Qx2d9RxPM4KORaC48yj9mb2+aP5Lc08ubUtkJxC83BFQ
gSViruGdPx3Jzcz8CFMdJxIKp/BBNd/DTAEI1kZtkVHwU5XhFVkwRs0JL9jz2T6U
FEyP0GPpVf77hb44uZRCOGl6tZT3KDotIgutMHf+OoBB6y9fi1eqz04NTkRrW/Rf
AOkfAl0t+t2kWeovkThF0xshn/viJtVfiQV1Ap62dMOyw1tymbIQoGl8bAYHFkPP
odDBRYqOrBLpaJeKpfPiHSCel+ztrtPBH2qFDFpOVU6rQ5HN8T8GHqqf58WMl1bU
KSZKhJz6wCuZTs2UXxHwgnojvtXxHJYApkIcpn/ttI6e5Q/Ed0QZOsBnrQi8pYk8
yRV94Apt8u9ijgzGNr6INFt9jKI9IZ3OSW7MUQXlSMup3WW6+FXWRy/ja8uS063L
rKHxfD5Xm13xbPujfzz+2fsUuzBBVDA4IAsNM1j8jhcNlEpKj2b9E072y/9LshSA
gxIJ0I7FjO4v47w4ygtMkOPcYdthIkH7e21oXWFBWnKAmh83XIzoZLSKBfR6F0qL
E4pheTRmEn4R4pDl2YDdG8fHV+FwNM8Yv94ihFMsFNjMn7HDfGiv3k/6sSQcmw9Q
phyBDOKvOS2vxAWQmJA111mmWCUFm/dKCNCQtH7CkdwiPm6I8NwX7ayFu5sPEI6/
qZlJ9iVJzTeiVhsIsHi4mVNs2I/xEqTN8rxJCgCUCo6jSpvReXakX6CRG/jJgTic
IN8+x4YvLpLMvjw5RkhMtOnWPgC5AREyC2sWemUgTMuCItb5XaSpj4O0sZ8CbY+E
dfLTvaOvrVdkjmTYY1MeUuFYiMZrJ0MDGEjBoPCfWRzCaraL3ZnxWaSkxtzWWupV
w8hXEf96ci3akoAzT5QqIVxrQOnvEE5USey3C/TQXbNHaRZ4WDL06XlBQ6N9D8GI
etIIaZS3zB9iUBDZ7btju3JUAR87e22wiwEhPHN6l5Y0U4pzh909xl3SbA/ESLo7
RNN8BFZ4A7M5RNCOj1CJA4qXqsV4Tr897HnlzHGejaRWNo90IrAVx1ZYxPiDqeWc
DaL1XstJEVDOsqFcDAgCYlIi5ZmE5QRH/iun1woK/O3WjtFddkhwrsoIsT/3DxK8
5bWpjybqglmV3JY71zeqnAADtekKluxXKH1HEEWGtSEnolyZy7ySrNhRD1SO8n7g
9CpXuOoN/29GtFOFbnlsjSEYEZbGB+fr6VJktiSCS5FB3duwsJ20ENkbBeUQ2f50
4t+1poqJ2qxEgGE0cWV3o9tZrrNDyoAmrUnSP4l3NtQmm+a1zgi7mgH006YpJh0Q
RsTRnHW/mFcznzqfpApUFVwjoIZyUs+4KIeBGJCMSTC0ADwhTQcwSiWIMkpF750d
rwS5FOFYC2opzzs+WHAHpVW6uDHUUyThqS4x0GX+mrQQDdaymrSSH38pXot+e1Ex
UnJLn5xi0PssqJS/OQHxuCnYrhq2SlqhBdWimYtXm7XU/oxzk/E1/fZlF6WvvD62
Lt4saz0yTuxkm4BjjTU7n12eeC6yt9KVH7VVQzVXms6ZRwp8Jkri1cAl0H8uzMJg
Lq/dg5MF44DxXkDCBF2EI+TKLSi86U+WGd6s5RdsVTq5uQ+lIGFNiGH94TwtkZ3I
6+p3UncuRvb5XpQdAeBmDU0biq62HSrxi0o8acXe2pxmaz6/T4WlcgxxFA+I5uBf
4Xvmrlw8hqiXCdbWyUQHdd77fVSNqc45ffh0r/n4HgUZQRhaoJCc5Ni8CfErb7ct
RxzMQASpkXtiu8qCfbPdb/yfQPAmPS5DwYyDAin0e9Qnzw1D5igV04w641BideFY
SzVcZv8kpDjkq9VKCKjgiRaDeQKGOeeU4r13785XMI0UmmjfX3wVDQpcg2pDm9xf
nudfBWRWOjMlh4OMi5u1EbOSOd0bOzDW2BFCW4ubrJJs6NGEjWZiqVZc4NHiELD5
Vv5DsBZxdCvubdIRxmidwf29KtQ6LU+x9riQma7XpRP2qGr0bjiaVdooiZTSDsLq
7KilNlP2xfRIM3Xcr8b1bNlcQ2wLnvcSyjY1wMt53vjuBbpJtJdU90CNGBgAp3VW
8Qlq3Vmh2HZAoxgAo2ZjyCjtQvXFGcGBYDwHMcBIZKmFpYqYIihTADsjMPMZjqTB
W/6mnH9oOoC8z8+z5BSTy27yGuVK9DBmWilRS8wwF7iDSLxEQpZU01sEijqSoeRa
7sMDyduvRgGSpNO6WfKGTkMQSunDJLwOZv7m6Um83Ege/+AItPF+Y7seY+JFsbXD
sBqiW/pGqRzVxNf2jarty88kGV/cBYgx2gejTKXAzgvu1LNY5jAyjX13JeS2Pi+8
Cto/1GnC4azraCE4p1Ufu7WUke7hElMBhaA90ogt6/lc7UMRfsmPzODpnszbb+Km
AAUqWOUCr3Ow2aJgnziPhZ5Yh/a5wada1putca0oVO6N83EuaoHkHhEL/Dxc9fgG
cOutVFsjSl8/+H837Vxvb88gm/vmgNN/L0ZjKizasBczLYcvCD1tKVbgOqLo0A3P
30lEkhJNl3x675KmDEZpg9+uT9MRxtRcG/2xRvwnhqQhpfvNIyG0O0zh+wVEFHz6
Tew666GnMYUUGXW/ZcGh76uAoguhrJ9WuF4/AymUKWH7kOsSqztDRUFqSRilbR5a
+IlvMgqHK4OkRzEtw/3a25Qn0GWpiNOxldidiiszADsR7+vPQ3+CYZt1/RjGU96Z
IwjP6ni4H2/Y1bqyIry96s88ymhyIpWlBPhUjG58Zgko35iIxmt08SuSKYMVEvPK
2kScdv1K9N59xKS1oU79QwrbljUK9GzDakUIMEt1m9zzfqJStqUP4w0g7H2XqbfS
fi57+s+V1InYUfKR2pskL2darBWVos2oMrURQvZa5Xk+b2sg0JlffEtQ3okWXdFT
tMI2TBcEmd9/0dY853qTzYjycVT3HmsO0nMf9iIZTtPh9CW81C8N8PVRGBa9DX0d
RF+RRcnM/oLp71AS+TKls6Pa8LRaz3oKQsNWCu9N1Ywv5+wBexH6bvXz/ctzXbgx
J8bzvv62vuEm14C25jNsXz0CC9k9eeMQtBo7GowO5uxQI8kP6TPqD07LbMckd5ZC
MycTZr3gHqiU0PtLSY6BcUTqPEnc+RJu8QP2kFZI+2jbJnhQX/8t38zflU71Jces
lRg82Wtk1V+zTWnXhxWYqS0lGUpfdL22MqqP12y91pYHowmTkdvXBI2BVGGbyjOy
gyOX+EQW1jsMxIPs/sao3/LtlKk0bEpWjf8nH3NPx2ZXYY/JfQhNz7U6qX2ojWnU
oVCV9srFmrYDnKcZYbkaoigHDAahmSwCuqofGaatWKC0F9CeEKTeoKpTdHrXvbQ7
oTj1WOpv3Uy1FZeZCXAglJicd7lZxn4XIBb3gpR9Ocj1BM67wa+j88n6buWaH/6P
pxHyOaG3Q0o8ebCKN/Svx7FTP0O37H7AhzGe/kuG4ZiuJpE+CLr5w1XIqHERZq5j
+g94aOh5WTkFmjR5QYdRVsjRg/pVSgy5hZQbJR5WnUveadoLP2bltV2K+Lbp+e3+
2qaKpevSvnALkEtUfxANlSt0beuop8FUT3j7gXIwFszETh30jTEH5zQ0Qxk18J2y
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HuYC68k7pnzC9gHMc4RGwS9MM5lKT0Mx8b9+wIUCdWX0QI0oPa1LBV9w2dr5Ozrf
JNJFr4WGymwlVDzNkbgn3JAK7GzwMUstYfrGaqT76fQoYRJwzEA4SAdW3wByWumc
piCDQPvHlmYXmRVrCgH6Q3vE/LC09L1ksTSyi8HDebY7uw5M4Oa4CcmnZIreYM/O
+zfyE0nIgKRMLO4o2ieJcaqa1Xlcg9ZzPeTgwLYb1eHOMMoD2LIap1dl0BS/O11W
gmHY7QLIBs9Zi0n4brMUTAD/OUa4d9GwDrDz0SBfC7F5lM6Nd1AzGx57D6n1EGcx
8mr8fky/1CSyFtOlbW3wBA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
5CUctd3CBm+/X561C4PoQ3TnJzMaZU3rJ0hT43fYUaQ8V9/NlrWIME/vWtVslJUZ
esHcirQsdPRzko8eyFmROZHBULyxLtvG6GOBIzfZ4TSLMAaHACv1VrkYI1YSqjuq
wUZoX/V1U1Owtw9qn6KGzsWcCoH6EdCCiDUQg+qEqXqTvh9nRaJ8sEcd0cz80JKB
PIEZalYrds1ul0W4RO+TSsy66NJ9lfz4NfEYUudK5/LqRQTFreJBiWr3qTdKQdBd
n0KFNYx8xOCeeqeT8lpg7qpzV1nIm0LiE67xwIHQJEc/xcL+5fQNrTjsQ7mMWXku
icDRsIRRQFoxH17RQZj1nJXEW2DDL1cKtneyV6vs+AB67x+II3G5gjIl/RFNzSKU
9DFF2aIKZkYMW6b2IaZlyBxKTpSj+1TnbAoa9MW2vRvaCBvfaCJQVyPTaOZ2J6N1
5QEFPYQPiHwokRRVsq9SzcEYLB5T0bvC4X/wLZratL5KvzMYAyB2mNKIrrF6wxhl
BQNYKreKy+GYRndK8v/PNQyavShidlqegb1rJMOmVQKeja7F4lHZQPK5A589p7u5
NattFyxpQqOtADzz/Bgkh4vM0f6wWL14Fcw53xM6Cc8XcEWhN8w22rK5k/dA7ED7
h1vjcjDEx7arb1xa0cK8+4KhUucw2M09Lf5ZMp2l8P1oQSt1P9Yilfar/qGMhVpY
ldX1yfKITpRjniq58OA8O0f86HuytjLhBmMjisvXwH4Zs9uvMqgwyzop1f2NVtcO
vogPgsry2Nj+h2sMUMfl9zSQ3JQTxeXCBvlUCLm+5mNsU2rhtNLyDkB7MwQqo3+x
hrim0n9oPDRuWIx6u1rwzeAoo0Ls4d97FCilq1+mI5c860V+cOsSn4Yl0MCAUt2u
piYz28dEhYnfth8NInaYcQJfdllIBRkYESxzgKYQ93w=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
fxlwe/uScLJBjdDmihzdo0Lkj6fiHZto6bdIs5mbiI+6mU8eL0UE1uclw67/fsI2
ML/a1T7+L7bX4OCilqJKTw0tkKdHr4YnjVspiSPGu3nF2i2D5vzKG5wtjrOrLRv5
jpphie29sh3LFg4V4zeifS4PUyYldM/CIGn+BKoHCTj6uYqBGJVqU0OrdgUz6Fhi
Hl3RrGYv6GyQ+vnB2/D4Mc6yc/Y+MBFJ8fTlxXdbUcbualhRvwhxYwnOWqOU0JuE
Mug3CuQZmOffSrdbTp8Wu2sX96nxLZfJBfmiwDXX69GKlc9e4Ii9BeL+Afj0q/8I
8R7IZOHpQjLiRrsDhHflZA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1792 )
`pragma protect data_block
TpJ3tadkFMmE+Plsu5jY1sfWGhXMRkD/8FM/D8UVZJGzxs0EwxcEriVE+uQvauBW
/XcCTM1g6T6Dn+dwd3G5enO3nR0UJDBsQrtOQ3MYE80kYlA8aaxCRhmKGkgMUOa8
7kSuYgg1Cs22XkusgITVA1Q/cexH/TMXTyEZteuM+P1rvsUQEmExfalcrJNKLnpB
c7BEhwI0AFeiiiArFIPSoy+uuUEjvnZg+pwKIrHZluR9V0esY00xwIrJOpeHU6D/
I/ZZvQBGmmQUVSvJc/KRxIgZdf8tijPpg8suyRWQuwq9Z4BbQwMZ3XM5pfxfoM6A
yhCU2clzu86x7OReJcNBM21X8xtlulHeIZnwtNRTNzJYoEIEzHgfiCyWY3DSKvt6
LkDEiL/w5OdvKzjQpa+wsyn4BfXJHxjpeFUb+B9Ml0bEHv2J+Cz9lcHbugDc7fJa
Aa3A3qC+df8jZaVEU/nYwNSw2xVlHvD7ULUoBXPAtLFL2MJbr/5CoQHkZx0O42+0
I3R7AS2ziaJVdxr5Nofpuk3xineHMbH0IpX08tsKW/s0vQC9bbtQLBKZhKBW5m0D
N/XFbBMTy959w5GSh8DoMvGXEKI4PSx/tzLezdNf31nGi5lpIIxSt4K32blp75ay
X0KtaFC+BR3u1p+CdTsz0GQ1t1R1jdPLkdEbnCJ4lZTq72gqhab2bQB+SS2Ucnu7
Zar5btoAgRxqzUg0Ts4bV7gcPygDpb0Z9GQx0bV3yd+CGr0z1D73cjKx7A9hcJH0
GWjuOnOOt26LuqzB15s5gzVthWv38H0U3tG0dirUxJ0XLwpGbC8dabQgs6MdaFHC
iRdJT+hz4v9277VPdCS9uXZV1uOZlpz1u0yfAx5tQcei5xTE/otqXwMJL9hfN3dE
f/heTEnuW8bR+sHNSa0EDNQpGdyEAWheN1zgjndZ+7O/blMCyPVz4lSwl+qJTcKv
DOmDC/d9Rt2Y01HxOAkrfS+Up3dNdedTMfsRYXZikZ1ulztXc44phfSvmeZ26FB/
6/LvAxM9Lc7/pxAAYN/w8OIZ+DnV212PCHCorU6Q4OXQ6QrhbWEFRKagMkPc285l
RH/prKuEicQx6mpaKLPWVl2M4dwEDLB8hCFzoMWmycXomFe5rCRu+sCJAOCGXrxj
kX4//t0QBfqiVCWZ6MTzaxAWgdKFJfkeV4Pgq2kpjzFe4d0UWFNGpA4+jTPzUhHe
KslSzhXlsJcD8oyVJuHWlrseHC65ZJbE7EtU3IX/cDdAJ4PqDNFoL+xBLJQeAPHz
2C+0/Tz6n3w+HouTLXsUOvTrX9gdhrA2PA7rxDnMsQH+7vhZmnqGYlkyufdLyXni
C45YrYHU5KCupODPjyp+4AYMP+dKoJJQN//3gCXZJxhqya5w6WA8ZgSdVdCRGlyo
HfMNuXsYginsG0kBbexvV4m7+aFlg7AYcQuQ85TKJumissZLTCv0C7uKeTpeq69G
wlnv5Zfmyaf9kN87zn8FC9buvkpybrX4DOWfZR3Pml6eZY+6WZue+QNmefzD8+t/
/Q7Fb4B9oW3QbUd4MgFVpkCysCOFHZEF84Ovy2LVn1F1dkot1HdDx0NLtndsJqft
NRQ3S3u1IqP3053rrrxHx48FpVRL5gwSjzGlnD7v5O2iSy4nsYDJ+NHZGPdpDpER
KCsiVsZ7ZAQBIPmE6nBKIc9YGKT6ShTBXT0k23WpOIJW1obcN+BC9PPe0OpySEZH
DMfUVz6eH5C9dNtyMPMuZDCEqEQwYfRVLmFkHL8rar04+0AkAhCGa/pCfG3ANiIg
Bq/fdCao9BbAY6gUQvrqPva+iikwJz8wjYO/5gtFPQ+UsHFtX3PkPRWp0vhu3MpA
G1vTo1b6zGf+dR0H/gcyKzEiwI+liL6oJO9qwQ7mAkxd0VK4EvTltlQDHYi4szFb
/2yzaOWlSg93WgmCjzEyQnhYi/H7DSSAVv0vdcqWgGtnHEh5PZ0MSTAVOMKzand5
LJfKAkJVpqV4pFPOlsmbCMkLa4MHT3aaosfkTpB9rlZaUCbvfcl5ol4HXcWzmlI+
pgNQRQLEy5lNHT3aIkWXlaCRnbIiNpSNXVoek3G2OWhX2O24+uW5GxMpkhUdkbmc
x+LoaFbUpS3nOxr8aml8Eq42QoogVJRyGkG0QiuW5M98ujm08kzIEnrb77kQxT94
5LBitbeomNGgpPqFeIjlH4BJASIsOT66yVGXG8Y3sle7zl6VKukDwExb+mDNPZQc
ou6iDLXdZHDirTl4V7PrIUkj1ty+i61QZVbjFkJa1RfITCAuVLM/3u42eNt82UZE
wJOGtee33aqYQWlD3/oqjZvRmfVcucdchzoB1uM1Gc430PLai/uqI3ZGBr/Lgifi
a5OAad2S8GOhcq2HAqYjQg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
C04DrsI17ymmj08t4V0QF96Yq8u6d/z8UjL1I5RLyiHsjg1UdOOZ0foZJZ2oG88D
RMd2jJKriTiKBRGhkei4r7ArrzgXAWocVlBRlDkb/uNgwUaAPEXzExNFwlTePc8y
91DULU85hWXAscQwDUlaGWDhra7mccmTfvlHzWgdXFeDjMCn2t7xw3S/9fYo5oTb
+9woxNjwqBYZ35QUT6ZzsT/4sDGy6IEk4FaI1EjKKxQGPKd0xE01lkzhmeD7p8KC
H2apQsydbuvVxvrV6AMm7EAJ89bDyo34GeJwXqfdvPa9vcraFnbyeTm/jyls05v3
N2y3Uxepux0n7vMvIBR3xw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 30960 )
`pragma protect data_block
Qc/fCHAQ0B+y9zeo7anv3ACa4vceS+VP4ARk8xAC58CExkm5ELLM0xtJftv798J0
6lJD74cGMN10qNmp97w73Kl0lotmKsfNSNKjdBgmS27hw76pmuxuWzA7veWdEdYi
yFY9jPUTa447apxDDcbvHUD98QOrHhfGr9ONpXaJZymWqY5mtWKw6S7fWuMKpXri
bKQdIR938cn1C+bLOgnT5vYvZEyC3hJxGCt711OOEm8FvtTWSoO2QawsOZSLsGrh
cCX6gF4cC+DnlsO6/Zi/4+H2HGtLU/jfJJ+4WNPJY4YY30vYrMz8G516CjprObY0
fZlk0KnrC0BtRx+bzgkIN/EEkv7FOK2q223UB4WwcIzry+05NI60GHiNgob1F6Tr
b0kKfkb83E+fXviFKLmZGUN/Jp+FjESjMWqBAQwuYXPx7+gRxkPBW/uVagcE2fnm
A+QrLdGC2sYXqENIkZrSLuhtbXmezPS3I4RSYDqnPMTuxcfFvOPFlYPF6zlM2alA
RsRFG+I98u7ZYnWB8qZEZu8UZoP+uUcqxrEEweYNN2QL2OoMIndcx44F16maW1ol
jzFSOfMSnNB3ltIDrUX5KCuN6Sp8FxEGs3Dy9QurJYZQ/t2dTtcxv/wJXChjykfk
CWTNXXCb0N+iv6PGSJMxsSRu09SlRSB7JyvBjMtFJRKi8+/+lajwCxtTh5FZOK52
IlrBcdiY19mBdJEzSHElypE0QIQ4PK7JsqdhM/gzj2Z/EAznCabKse4zt5acX9CA
WspdWZGL8Fum7ES/or/P19KxHZNU2K64XP+nt5N/SJTYzM356Dprrm+gin52OBu2
5CPsey+JTIymJLMLfFW2NOwO9gvYaSpB4mF836ivYUu1U1BskXs/O38DynPzuZvX
4pFutE1o43+zKjracmCKCr73i/mBEM33wr+8iezjXU5CdtKgFufOZiY8e2MGquW2
s2x4C495kHXvReugqRaS6TVrnzVYi+v5rvV7R3THWsEPBmCU7Hu8x9EjlS2I7JNg
wHCxig/CQGpnH0Yqpg1cG8t/Qm+R8v3G1F99vMZ4Jg2CpmgoGtNc1833XN4OcywV
u9F/bLzcKfMvbTSdF2qpnAUYbzQvWUgVywxWTCUxIE9bt1pbk/T3xfQT9hRP6lq+
rQKBEs6/5NiEDoIlGrnVjQmrUwh77lCSAUmopt+z7QZhtXuOacAa419eO8aq3KDr
zB18PNW4Fsf2ySmsu5lBQ969QGfETZp3Amps/mZPxc6aAdiVCzxs1qH1XhBuX1iR
z7xkgOYQdXv6LAnRW4ZlWTIuNqyy1EiDAUlglfS69afKq3RnOzQ8EbQRJ0GrHjkn
Od3K6a1zPAcVk7stu8S3/OKwnqvQGEzecJJBoDDzJQBPss3AK7smOSXFFWnESZiz
n6IUeWwUhFtcaeFOADlo83zfpyabdY4pRkjeU8QifTAy38aCMUtF9uNjmYreS6XJ
2pswxpKtAcvg2tsrIDoO4+pJ/mZW9TwBWEYe/QqFnUOlXCg/+1p6cZoETRYN59+B
edjKMVo5aEZZP7T1zjpXfjMvgc2bD3nq7VUERzaKT4UrO4SlFmYwri3Mih6GPmOD
jwXYs/V2YV14Hr74JL5saxXMulVv8OtlpZUwtgC6L/76lVz41HUCvZgxK6qR83HM
o9cYPzVpECa+4o6hSUVraSgIxGvF/bqCMUPfqXh3/+ANCeswsmrgYXqvMbySRhlE
XHo8Dw9znIQOeCEbVirJGOPZE/A2GREtSyl8wkLgssn3awBvRJlVMHVfwgCf6N7v
EfQ0q3aZnC3lQQ1m49rEL0U78wHwn9kPQt4xWhh+4wo5fF9wFztqP5x1fhyPl0pk
fYsVwL7pKu/4EF9BjsHLyy0Mgm3l0wE9D/FE9+2DzZiRB01LXx+7st+HZbBl+ym2
pnwiEkzvoXg5IzEDwIYVfFe5+2gPEiTd1XNLsk8CTviJEKsqmWM2Zon+VjHYdcRu
JnBi3j/AWCSXLMIBvjqcv5SQulbXCt1f5SgxRMhL2fNQntYtCBUk2vggpft0i8n1
ut6VxVTBreG5nS4YfZrGZabY5nLfkYEx4lqcwPD8PyOezJxM/1qlri/napqaGC/n
yWBN0HNazVcP6ucDU5AjDKQencq4sDfBdP+BCD4IIygyo3E9uJ+NKRtyRhHsXRRw
eC0lbwHlKgfgwyy3ruUc5qCPiTnLgmvVqR978lnBi9+9fcGIWeT+IjddS2DToOHZ
Xs9HsQBi9LPnG6GU47IamMUtqEdCDBKsezFLqtta3vXiiMNX8UabTz6S+CrZuQ9p
bnEjnhzy90XK8dBvPnclQmDk+cvn6hJfVmHFt5vDxQVKAzr509LYZI7KtIyto3pZ
5nqAo8mnYC7TobU1/130Yzo5caO4ys0bDJ2HBSjV34KQYLbDokK2Aablm5BMBJU1
qZLBO1KU4s2ej5qMkPsxmu/ucbkrhnIqR5NZnO4YFo6S8vYC1RERChZYlua2BE5z
bOpcMj58uVv811liwLV1gwtIEvfgz+MoCddIHDeQ5KYt7hzRYud/xUe9D1T3PiOu
c69aEcY1xa0+acLcfgaUGbdkzN9+PSKAfpggS2bmgbrshzGV8cxhMK7YePDw9Mwp
A7Ct6z/a52B31NjfFFC20QUmiNo2+dF67acWKmIvYvotWid45VeYvmloreE8a4p6
i3C2bSPWkyb6oVUyML5vJLOuqN5wlT2PgDCy2Z5ZasDdAQGsd7MaW9+i0m+4vPWy
Y3tPEyRcCJfKcKQw5kJPjIaZeDE+JyvcGJfgQ/4Ua6/wh3pZKMV0Jxi+4OrXlAq9
B7/r6XS843TDmFn2dgx3INpavqYkJuU//PqZd6jZ3OJdwrHbN+qIb9dFR1wo5lj6
4ixpeZMf+cDpdbYtC1FdQqBEOJ4/lauCveI96MgXHI3L2QxbL4yM9CtVkqJvtDOE
AiYTSbKsQG9fU16NvwArveTXKKitbRQQ2MOJFd+TZmwmw7G/XvMJ6bnOwbgXXiyx
cnfYA0g5BxEWp+gjdhPfgBt8oDprXkIbl3UB7SwpP6CtxMSshRLLVUcOLp259VhF
C7sk7MZBKrmb5WA+h0qh/QBJqel9gDS5I3canaPbNt/8LHGHG27O8jVdNR19CJT0
oBTuJ8eyEsFRKwAiZcCva6JPjvi4DhDO2WAOjTiyB+IYGXUHJLLdpJ1PFMbJbwyo
h1LAiuzueG1ybS9boPZig94V7Yu860HLaimlQich3h7soMIs0ZbokcxVtx8QcPMD
OmNYhLv8Zt8ymwsJN17cD8FHq1w3FAD8P1vOfZUG1WVbJjI2gdsR4AFRjoc5Ob14
qY1cyOo+HA57iEeT8lPWLdkpmZPqp+ismQur/pddxLrl0c6mDO9/NPHh0MKJYMF3
EVXQEeIEL82V9kiabqaRuGfu5sSpVqpuoeQr0RHxh2xuOqVjFyAfZEKjugrg3U6U
0QO8QtRVuaS9LPxH3Yb3Yy3N7kmxANN/rfZbYA2I4nBKFtpm52DhfSWMCb4Jzyyy
UyruMdimHr72A5QmKmGuMe9oVg6UAQcWTPNbyMqCwytq/3a+wXc33fx7jA9Hzt91
dbAF/BhywYp13AvfE3XtGXmVxwT7NbyPiB87wUNzqPNsaCyPi86cZ/v5f6WbIDMD
XQekioDBs8hNX47egqD1GDUcCgsqrSNdM9kh8LmyihLXkFn7UWyXhZCXUIk+/mAe
1sacMYv6jhVkuwK5/I/3akOsBbBbj4AnicG16QlFSa9FD/dg03iwXCaYwoMjEpkv
y9uDZd26NuDLk8RaF0a6UfEw+P/QK7FwMCu/TqrFzl/AkuIRpmGGvFMu+MuY6qQZ
+xk8xYr+YRfu0U5fH4pI+3Lp5D2PLLXAXuNMkLX6p3mshqZQr6FIN7l/F76BJw7u
itg55hnsyPtyZctKJ/btDSINr2xD8wiFpVuWqGZI8BjjGI505xrcybUSLcF2uVLW
QIHO722p7670oUfrTbOVIqBMPtzyL3FWdD7CIc7RnQVHLTiIZNkI0H4qK+G4YRle
xocWKzLOd5p7mfCtLk98aEM5cim2JdAFi+hWO76vAyV8SnASagmSPLO+dm97YVk3
AAEVciLyuTM529LjaLL0fhpxQUhVER7W9CD7VybDmts0RdjmeZeu1UTEulALr1B2
cL5uONNIxC6MicZezNl8/PBlJgk2RpSuvIB+MvXHuEvf2No0wV4gyFKaGzcMNjmK
4yehtCbcru5TV/Z2WA7vtmGjMQFOaSZ+9AbCXvKMMdPDpBYtyrMBjGWP9r4Ns+UR
Va5SvwRKFTAfRluksH/87miAN6tTuCJuI9dmxzUc/3kUypw37CY0kG5j6aVheqpN
obolaJ34ZhKOA1FpK2N/X7f+9G6SQdMtj/sAa25HVeg5ifE5pEK46vOfsahg7U39
JeB5WPvB0dMHsiBEBgsN6C8fyZC8dJR8Y5A1kMI+zRTM1EbFjLk3slr0qeXlDD++
stKrvT8thEzxaDsA1wtJ19yBsTW/tuVH4au9JhyakV7X8aXyOd1KmRXeS+0GHtQa
rUa3Y1e6JcrUF+Y+o6Y0cM8f3QLN38pH4vf4lExriLyIiW4dMPXYTSPAB8GdeS1c
gjrXr7KvLmnqngCFfXS3X29cSheFerXF8cZdxbKPoLh9bdETgGmHM7jfeLBsbWuU
/QHRHn97iKCNfOcsxpwKb8AlEATN1vlTQlvkT2qMnO1CAaGDIXEQlZ4447VcQlQe
A1RdYE+eSC9f5mjoPUYeLlFuO9rv277bNUpqreyjdEgldI4MesF84MSBesfBkik2
8rEags1Hlgx+rfWeusvVgvTycScioAUoHQUXj3jZdg7GM8b2gC/lqEI69D44UM3v
leBgAqo0W2nzvXge1+hoI9UT58c0+5eSU2jDLdQjpN9KT8HkOFeEi5O8DkQXwk8F
UwslC6XRI3Nopu2difyC/+0KcF0t+YEO1Ar85Sn8y/F+BUwFiap/nHuUeO1LoqKR
gq641r7ag/RIG63DFlD8/MZVZC9BDXH/F9AGo8SRNlJ8DSepIJCSVW55XdST/Him
g/8590WmhreT7Mr4IWp1DMjpgXie8Et+9RWCRfczXMSAeUvQree5pxj+PWCOyZ38
Jrb4dm0o0tDkzx39FgUupIEmlv0RioBtN26SyQkOwZ5mPPU6t1Fgo9gIgTrsdMrJ
+AfTNY1EGI3GOx1Re5/qCiqK1+F0UjYdC9ort/VuuvoxUnfK/Uv3rPxrNntPFUYl
LRi6nmsseQ69MjhNrQHCaJQc+QchUFm3BzdlYDoizwievRSdz+0b5KwvSk9bTLmE
mHD7wjPjKmM23YQEq61dv8iJu7C95pD0MC/4WHGuujF96qjcWKTzlkYBEJCcByhc
0m4KRwYlKxnJZUvGGawEtkHg2nBokT4c9bWzWUqc3OvpuiBgjwYbwJB7AEHwFrka
dN1o6hNnhRi1FpgSNe5VMTgzGr2iffnFl0OF8GxECLylYrVJcslFsZgqHxDsnry4
qDMV5sBve5o/dt2DOIj20384pSjehK/fTMqKbWG+OhgnxrobrVCZmpiR3INUHDEW
hi73NV1ouy6yXr+eMKK3a0wEtduJZahkEEGzZ7X5yPun1JGobhUYuIapM5GlLK8K
yslpENMKCL+SEMG/76PAnVRzYvGmSBWMwC9T0knpkjE+DYt7kgD7+q8mQLspjggz
0oNry+JzECamePlhMDm3tDVOUajD701iH+l4K5qgdVthDNBzKY7pLQBMwaFiCgDH
H+Nmm856E6ou54SXbGvtj9wIiZzdljjZIdXoHC0JL0xtDWvM0TiO3zPgI/ce55DB
nmvPFXtKICh7B5Rvy4uM93GwShT+lBj0qPrtEzD59CyBzJLgKkH8tg9lwqrm8MkU
2ICjKlJvy7Epzcef6FfjXIrceIBuvcP2alz8C7kV49WAcTlxUv+SoppgrNA/kBMm
vKM1/bfnfkvGor0DIi8OxQOAKgSOj2qc6qpGj+x6GOs3xCXHmVRJ9Bh8Mgoi05gB
X1yl+CUBPr3PzdwMAsic8ZsSp+liSMJXbYrikiOmSSjhPzoucUAuIo3hErDhv/rC
QJtKo1GN3MZNXa/KTCn022vSUk08CW7I8x4eOq6qatrOZJCpSS26vQQIS4zaTEgp
NwFPar/YroKcZOi7y70ZqxvSo/mQ2J1+VdAJg4LtOOFII6YeNjg1UX6LpdDFy1d0
dhovuXbhoGyR12TEetdSoBqtdog+VmgdpbtkBBeKiZTMEkcvp3VALYbsfCAibgvm
lGJzkqx6wosUr8Mk0QB1UxHO3pWrloWo8aLEhlkiEG3Mi2rq0LtunTqW6rf1n0RK
EuhuopjqeWiSOGnJXxO6EQgXXPuFtnlQnH7S8dnZLUBh2Qqlbb7pbpKPqFBKqSZB
KebKw8Zx6Fn3kzRpbFiLqSui4Z3eVNwdyqgPN1BDPdo6H9E+fMWEYZT/5X/6+e3b
U3jltQkHX7MdPco9jDZnSuPqN8RstuljTuPTICS8Wlhy05Jb4TJp8iykVppFQnDS
gbJ74m7TUCVw7s1rYBR0+8aVezXt/RaJFfBGFv17/hFWrRGTtBkwv4Zrb/tLXPLv
lLsy0Z5nreMZH9OnUdVCNyjssAsuu0g48nPH8PKIbDrYIN3LZ4FA9dCWz7oilEcO
GLIWtM58k/FvQzZhhbb8WL2pMNIOdCJEzFqTHLAReEzQ8Xl1etXntLWH4oTY/icV
yr3txn17UMGbbp6U4ww1+CjlgHVb8TD6DKFJZ7vd3GHOLC0uVuayi25gyriowwOB
NyTIhbk9JfvxjFd+JgNIRMmNX9YjX8IEfQBLYvA0HUTYdPebMK/oL5LnM2VeK0w2
gzJsGCUrA63xD8lJ6NRZzR2hRvmnnsDualyU+QRs4cSDgcFa+vKhSq2UkkOQG9F1
GCYEaLCUQHnJQhqTKn4p7TmxQqGHYsYx7eE9pIpsamDfyfhB4ltYRVo86SL8zCbZ
iKHkER196fOqVLRu7zYEFHt/t81+ujmw0C9IT7P3qDP+9/UAVl6bT5/fh+9ucJJe
4cDosd3LYGLkXe6KdimNycWNbYpIyx70EiLda4/ST2s0mwao5UAH0rKPy7g4Pfcu
Hxez2pYlKrkiIO+mFnnOUpf2K2tPy9pX3prWVhDwxy14LCKEiR20WP1AXddEcwMz
JZNE2kFRpdQy6EnGq2+6LS0geaMmWusfYIZ6zkq2yM8qlxbYjhgmAIGf+w1f9iaQ
W2n4TzQcekfId4+ffXcVfSzK2hjg8MYVVgrDWMa4VaGb4KJPPdlVJd01AScfRlBC
RxgzJHHWDE9cDT3/1pEoGWpSQd4fFeN5iOmS2bjIe71rUP0T7REQ9mctjkBCa25c
huMqNRLoor2tMPr0de5WmhkLO4XKMRgJbhDp3dXPsa1jnkImH5zqws+87A6LoQtt
I4DCzj1PwhmOuz+o5bmfhJXTfxpOIAmynbURJwRcpRHNq4PKNFm5togUsi35j1a8
MGSTb8+D3299F6BTDzuzDo6ZUHXaI3g+AuwAuYUOO8PR9xKqcACRT9JMYvzg6Gh1
wIUl+GJNckefTBQ7KBf4TIFLryWJNd29g6sYQwZujGU52MeCI+soiqW392UqJZRI
o9dwIEMCs6EH+qrIE/HpMi9BEN8mipOn8yCNXAhQb1g+6uWuyLD9Z4/AUjHbI/Td
Sk8Ph6/yT6DEtdEYOxZyew4lKTJ5X/Kfaw/WnvI3Gyiq0glgGIAa79VeJRUS20VT
o5HL0gM9H0f0mOTTJ3n721bPLqE9hqivKbXAgMf4hyIwWmHo5fEVh+DohzaPHcu7
vB3kqi8N1ELHYVhabtYPryMxA4nLRJwgaSc0T4LY/YoBRqXmD8qlDku+W501GTst
M1qV4DU6QoejQgSxy3OhM/PdYB3pkPyua/UwFkHY/a+si2+fpMIB68ySTLuRojEj
art5xDu9hTixUonjNOsBPbdKwoIB7/xizBV4WkIVXNSPEBBNl5/PNjxinYUsBvcQ
OCnM7Wmx/x12DxcOJfm2xo02cUhDFvfFwqKRG/9OtQHk0Nw0eA7n+zx/U5CbARfG
iyv+DE7EcSmHID2Uhh/ZfE7kYoItywCCywCG00fJCRbrV1pXuARPo4ZLdu4Lunce
ltMfNo2q4LMlLV0zEA/to1rmnZsNTX4WKV/TcWPF/KmlALI2iUyLxhtooZV36RAL
c7q9YNcF24+LyLgR4Ec6Cn/nr9T0En05rlHw66vfQRoA4v2NtNO4IkpURtTIvW6+
n9NUGeSuo3SxW930rDwbAHuDN6czz8kKxHjfysogqYAm9vxtbbSJcMUvTdDVlTbB
+h25MmLrOcV7PcmFfPePgc+/77xRZEqv49wmMWI3lM2e0/vRiPvoYkrFstKP/NxV
TxEisVxvojT5Tb+DwI3FtkaZJ92cZx+gEOGNSN7iqr/f4gs8s1DObVxcKmF3rN18
95R0I2flNnX1G/7Xzdjv6h13ewFEy0WyUkQBpTHwTILMKww6FyNS+f47ygVXm24T
i6WKTORIxdAdD+K5bHP5dXIwOYfwChhwc7nEUtjA35UEBwWkiv3/TWb6oYFj7E3W
M8hQIozS2Ubb+eacntR8XUPOFbFpAAU9AjR5UXEIdrQu2Qcyy02aWelYEibjoeXV
iLknHK5naIjXk+8iwEnilRcxEeIX2WyeWouT8c8ckUhKTjXxchiE4yjZSfhZE7wm
NRueK3Pad9WJ8wziSWNF1LgC2Gp5SvajSKFWwRtbQTCL2PJA9jKfhGV9OLACsX9b
cKXXjHEbDGh5aHC8GDqq6YtO2cZOInT6nENairwgSKvmPevHhuh6aOERIi1Q/Vo8
aNDY1Tl8WKlS3zSEPTW7/GumMVaZRu1HIQwLBcbAknF6RtESnzZQ1VL+6y9Qutzf
vQgCV+UseSFND6JdiQQEuko04I2ahOZN9815XHWo3WhybkiQ9fxoZ0firHNnkhHx
VtAipu0UE5J6tt101Jk8zO+L3wxD1eTmlxnQFs8dxZP+snxuFDdXLQn3/AClcIbG
2+N/dqeFY2/zOF7g4ZlXEWXuFFjg0ZchzHLdvhAXzb+hvPC6L2kJ4qj5M0XQ8MF3
/C2M2OxDmP7GkUbxtn47gXqRINCN+Jc87MjPq6F4Msl9f9pOSzQY2X2Q1xxG+qET
7JQg5TwrOi6Uop6VFESZ+Yopus4yKuQi5//NFItrT3r+80qJw20V4FG99SC1sO4h
C1u+JSOLNC2thMMBhzUaCm2pxWW33s52NWv777NjQ49C0PMESk4vipfRjUNBfrZ0
eO6bi/4PI1GUbbSHcy6KUln1x4sjIkYfgkonZLLIEzeGuQTn8EYmtCojuU5V2ANt
bIbcg4oMLDxIAHhPXEQ8CZuvIYccgCWvbOi6WjQvv7csrbNOGtAGRPTQ52nL/Dgg
0mRpDh1EA/jA2TsxigEdhANWTPvU73w+ev0kQWpL58fbbgFrQ9+3/oNRTNfZCQDN
W1ZN/UeBGa4O7V1t8xA4NSbKq/wSZGpVIDmtRUPU4Thm3sCK3gOmOYJjYqgVjkhu
IM2OhUpGGSCIJtTVSKXX8RMDD64PoaJQGYTnjuHOM5ZzepXt0jM58FRs00gd1+xi
PMgo7Pfc+SYkNJiGziMzpKVva1LHSYfFe/Y5gPTwYFLo4mfcarMJgC0nZ3DJoYDy
IKodW1KQKroCp1zxmWsIWmJKNoXB12NcfHVxl8ZTlx1putdIeQXQxO7sXfr3UYEk
EtpsI6xAPPl8MbDcslB+Gm1U649lLxFAX1K79GJahfaOxPQGB7+yEgwH4eBMs4fC
SXK1wql6pVavYfzMflG5kWZ42o4WG/ujx9PRCVECmimjQPthTlb6/vwQKAUDgIg7
TglhssEMKDItpbCNhBz1+B0LVJauW0hIHcqG7CA7n+FnxCkHUB43tZYf4ruGRUgI
BU0OXvX83R2Z6lvcqolLKE+OAmMBI1RPQK1xc2I7D0SNTK8qeh3SXdSsoV8HRIoT
eTbxi1grR0IyMmvhXHdEcTBYtAyzom2GAlEwQtubOBswJ6K5ycCJqWUltwYOgwsE
YazsWjihZeQTi6piF05rWDSJy5FL58qEKNLMGMaNKspkrG4dFBl/aUMOgfl6FpUp
p4jqpV0KnN8MJpoPEgUUdqnSRjvZ63fR7mwblU8kU4n0q+qO/YeJY/bKcuNUl/eh
A9yDmY368T8RJeMC5Ack+warkllDE2ttX42fanwXWwOEwbE+xTKRLiSPxMXpqu28
NVBW2+HhlpiFnZlgGZF2Bq/PUVt5VUhg5wvmXVsYGzvjGw7Opn4dFykWQyLqTBl9
N5GA1+tulh6ip4+MJ8hMj4XUrICpKd4ttZe8cmbJwB1i0k5yr6HcBNuRlGv34GCA
ygRZY3YdyzfTH9szJQwtGgWFKQtWfVirrwEkF+iwRqFOUKD3aNYfJbjEgiYDP4Fd
qkaczQDT/DrDHUrt2utS31yUvuY+KOsZeNgLoMFsV1XOeG6PXLFPdnr5Zju2Nq9p
68FsmhqJCop+iFs/Lqe0EabBMHxJIIdhD73dh3MIGXR5gLjW00bOi78KKFOInXHO
WEMUI0JNmLXrnJ0JI6xgDSCcnkgYFCr5BkVvHscNcgWHUzCEH1fbKJt9tCWgPy/o
DmdWje+0Pdo/+7g0V8oU4AIV+tBTDaS6UQKWTk65HacngBJ10RAN6LcuZsGXPMe1
FU7B8fUVXARuoSXU05TmRf2juid+Df0M3Roz/BOi0Zn1ZrMIAy4u6K6eiy7tVX/0
mKYzDbkY6SuJAUV+FEDqL+gXN9LI6r20grXWGfZJo9LUohfnPsKabNn6g7IjcBzP
aNvuHVULdEMCOWM5CRm/NwLR3A2Gg/Sgnr+KRZPgS0XVYmGHHuQ460IfHWJmd8hD
CZLvC7N0+SEs/pVY96ief3a5QrmyjZBxfAFsLXi7XIfz69totQVk8EEZdeiJBRgi
Uj46lAHQXI5qyZliZBYrov3BZCOv+0Hr4DbngMfelrMf2h4zi7YlFii2gDHChWTi
Jk9CMFpWAG66UQqvmpT+MQknIr1T37Ov4WpFwlpJheyzPXl/SJ+XV+KWFbKduFIq
TcIdLLO1W28pXYCKoqMIfL/vjkuAaS0p/ZiHtttNOpb3ILW70dF7Jcz12pPb2PeD
SyZv6bA5QACxy0KsaMumDc66iZu66jgOkYuERmT+noOC128+0MOpBMRoLKzLy33c
NerDz1Yi2o3mJ4MGaxK0nCpBPZFTi30PBrhzcXhf84w4RvAC3+Tx3ncL1cjphZ8n
Li4SRTAk40vdotSHMGnEgc+ryh8UuB8ar2ieQtjO9S0NBSLCu8hPr4kKqk/MIBBJ
1Zv5OkKu5CH2p1216JwHJNLwRwwjpI5NiLRGVfoUE50lXjOVZV3DuMakbvAQT+pv
fGz9QKrV8ccJ5uUnCQV2K7pxDXpUIhd1T/DUysB1LGBc/jCDGp/OzfshchydG1HR
v/6/3jMwmaDv/ewFPCUQ/ycA7ghLV41BzMQDKToenLkyImHUMrISByD7YuAjoUjQ
055PyMwq8uqsCnlPNIkSoY5fQYV1n1ERFQLJxiuWns6A8nknvPPjJyp9OePA14w9
5oNO9PKC67SEGENpYPcBehd7AqOJXAm6AqLF8fmXjr2zQ0oKNyw7Y4IgcD2vUcu+
Er8Zk1uOByG4XkS1YMPyyuU9DbC4xnXuk1q6NCPPBAo7XoQgdfeuucOTnYLQoL0d
JJXnAqyv8VhQOXhVO19IO0VAUoFZTw9Ia5uMAr8Cttsz2+zhfP8L2Y97QySTaenI
q/3nEHdh0Yk/vPt1QzyN1HSTDEPmhPyVOoCwRO+oFOo//0XekDmDrKinVuRr3Dpd
kOpznMu427Azi6IhnBXx50sHJp0ILgJpkFh36KMyyulqcKxdibWqzqvirMPt55R1
5cf3fQyD2pSbrwPvVsKznH76vssUiVXsapZAiCVmSrW4byaEKerCkV05MfCnb1tk
yiFvpWrkUp6/r3frYdsdXAOwuAx3dOuxxxNrYA0npDwj55YBrFy+w4R3GwIVwDQI
kBOG+wuDC4BGr+mv3cbMPrPxhO44Ey4cYCElS4rmtmkM81Y3KSUgx8W5uUSXyRca
M3c+m9HdmbDQjK6MoJoubkE7c1PW27SGUp+DHp4GbmArZVNz8ujpkBdbUtn9SpqE
QXN4DnX/9qLvZQbDewTFfC+zQmwqV3Syrup+gvtamF2XVRjYTu/xG+w5UUuH5Nma
crtjqP7G1qq2gYVoUeHo3pfn8i9Xf9s+euMYDNkknuKLCSVbIQ6NGWdSzNfRGLhJ
UiRSsRR3QAb6xYk/MA4rcNSmPYQywll4uvzBjlu19sBEQDdHkdTe7ok5B8ZolSvS
VfmbPMXrELVheavaw/MBcSnAOxaHrEqGCnvUPxLbbQKXhAs/tXQGWQYTxYefuqsa
X8xRx3p+4iX+F4bncXdUVew1J5jGHlTN2YVqbP1KxgufnCrHUepIBUmYVPPI64ic
Qtcb1PkSJ7zBbjdk9tU+gWckRWFL5XZ9MimGRn8c1XaCaoet0JDkB/P7fEKY9pl8
Vsrse3zPBfoeb/GAKlCpRhDgA0RUpJEm5ioNNZRZ8tj2OuUU9/Y/1nWDKhseonE1
iYinz5ZazxvCgZ2Y872PuN1TN5in0RaqavwsRhrZRYeeV+9CvFO0sqerA0bQPosE
WfzpcIj6ALpskm6AW5Am9lpj0xw4X3NZPUnAynk2Eat1fCBlXI6/16++10vS/aU4
61isNgvdZSpJ5jNpF7kDqyETya9WQdGODnOR5QLYsb+O3aNsJUnF1GIShjlLV5L1
tEscE6iYav30U8eqssYVAHRrwEHdKwa7o6EKa86KDvzxQKnSQmnyjF1vWbLVX6jH
qFJbRjTwoGMBoV6znDxEFad3n3hjebQCUAlOuKdWZ1cvV6LiawN71lgppJPGPbqF
VjkRY7bLonhuJEI06BspXAbXELoiA1OFb3gvcKkWWmZyVSYY4Pnod42MAgf37ps/
nAmtmh7H7anR2mMSi5lL7gKSA3R1ou0v2H9a7z3pory5OdPGrd5U+xPJ2asUa8N+
QFgHomrzyGYnkDFPEsHULKpuWpN8zQXqCcG9qyxGlpP2aULCzckuFUQ+ZlQlffQh
NMGEtiovnOzwljVURjRe/Gk1bcQaJvQgLOSwwiYRG+UwaD4ZuGHIC6FF7h0S9rFp
bnsXQE74ciXnFNbwS5z9giWJrUPcIOGjkM7WpIJ85K6NHLYBCCrsw2t3mfNwQeDC
9XKdZAjDMDC4bnVRzTQKod8iBuxFYJ306i+bgtQZOBdlXIw5I/ZsJdkRZww/j6+J
8QsrYs0pSI6aI/mS/nhD7OMbflcymM75nda9MEiekxibXJHOxRUfZuz0Wn88Esh4
CmweKUKiQjJxLS/RmYsuXYbetwFb6cIPgMOBDDhIgprox57oOyhWJgEPCqZGTUyC
Ktq8AEb9nygg/tIeEWqU3Ms0RFYRcA4T6FbF6Ik0bwqDcn7Hpz1fg4SnnDHjXAEn
Y+/mB1DIOMdZmvfD1wtiZjKbMdRxpLUninN/dT3OF29J85HK/oStroU8Arm2p9aI
6ujjf5AhUaOwvLkNX3ZEzhjVC3xuYDf14bTQ3qYyFbWoH4AqL97eTFFMhB0EgWyQ
Y1EFkY/Atsgqtnw+fdFQMKmmain1v/ivsuPX6sd4fkKGASa++fkWognqLkp59xg+
K9W8vfqk3Qdvb6C2dbpefIXrkGerxexWeLxb4+KkX5dwZYoBh361NZpXkzDTsnaN
9LbEy67B2MYw4JwHPd+cLaACR3MZth6Qp7HBeuqJUbcHnnmx++BiqCUjeYj8NTYM
LVxiztk5ZmY14NjDc4rDXNCOw7hXooYaPg8HOvLQerktWMslqp0VHTweot0SdLCN
eJdGGg5/ofOjtc664+PTkTJtMVgQd18X4fGQCAQFyNk2bi7bPRKxTbbwK9hay/eP
1qsmDTsLSIkggmh/3RcNSmt+BmkbuJGut4zxEziMmeP5b3pWCpigH6vnMMETD6/s
gqH8adEvowl4+104wXc35t5+y9X9h75WdJd8uSclCv6T2nAbXAzn1nH0YyLARcaC
hFfDpLLdyOq5S5Q+YngH4rP8EX5sV8FndG+L2VePIblsV0CFcxBh81pqTctNNDBp
6/vgyq0ME2ILVVE0civt61ymkTRPl96zpq+RiAhinxMy2m9zt/0GT3M8bRAFx2V7
MHI0AiULOqYMe30+MUzHn1S0ucPxxHkQEHiBq/S0cUIiHoZO5tQ/IYiwSFkSbM79
WpGYnogQ2iWyI8gy0kz7EDifscsuOk/nWsO2SWZGLGTNsuM5Nz3wQAsDeJDaE8rG
GQx97XGbpp79TY4eNNqIONWrpidqSfD/rEJEIL1pPzQ061PKC4oatlfMy++RG3DP
vnRkKW1xPEex5GKF1HAT/yQuDORHYMs31jvrHqWa3CzkjYL7IVdec8oC54zwJRW0
5yuQ41kT00gdjmENYnm3L7Yhtlelk1v3yKIkFJuedlNytQtR8tITliBOw3TaAIvT
Ivd2nIU+01EkbMvKPYdsBcpI7e70aumvKnPi3OISkI9z8jYyEiHIpIUoS9zwaepq
jBL9VFJNNqjDjuEW/3QFEsLlXNGpZrN2Cp6Q8qeLwLu47Mb5AU5Zbes6ct+sCPZu
U8kl+UyVXhMM2C3+TWIkpAExuuKRwJ3zod61C1OHclUoumcGDgLTHrEFA2OAd+iR
QJcmE62Kz7CD7CAv7qWNbkg21QT3vxwYX6/VHOnwg3wVLAeUuj1xgXz5LYig2QmV
Zm/bPkxpfdPpWjNroSWzYRNmsmaYOUYCj+AutsXcnASBQGAKfksOW7s5Qcl8J6i5
F7DuZA6/GZqxtLP6xfYrW1PP/3LxzN3iX3Q2bm/1rId/l04K4A0mAnuWS6DD8zSb
6gQQA1CobC1r/QhUcuuqHAsWRlGYyXuj5IxdPKnA6BY6zMzs4RumyBLOqlB8Yhvj
G8WaPZkvhb6l4KlNdb50yRg56PoLzYdcIQQxEm31thQ57eOHSFzyNfVvn7ivfeyH
2xMTW/HHiUSLLI8fdpHpbEvvhAmkQ4cWKu334c/1b2wc9XrgHQ3J2g3zXMi0qAna
aykEupKr786qdd7DpnJsUmKNQ9ZB8sZKphdkL+oH8fzpGQBWGCTlp7di6fI6Aw7G
lCJOUZ/TbKPsFLP+wL9hgl/XyfPcUrSNxZuyZvDqGqSQd6wuHrapHEtiTc9B2arD
N8hUYQwQ2iwR+zCgcBDbHBucENw1gm1rdc8hQCboYvztHEGisqF0yZDjNTmmbAMu
8LVGD5smYCd5IgyfcxOXmkCZH6cHMLZs/mE9MGPeTG7jwkq5dC1F16FhozlYoFfM
RitAC6l9GOezyv3ZqvPcGPc87F4qyjzjM6iqjhSX0z3VwAqkNGaLEVsLaTQrTg4c
sPHrnyWN0M28M2P49XCvmmtfImGUCdgvQKh8hUX7XXfRW9ISR6QjIAvdtlPYKRYm
1BUZ1qkzBH0qiAYWPSUwAdLtvT8ZSVjHbpbdwQLkrdQ+S5pdEAXdcuUYzNqVwRv/
hUL+vRc22AS4GavSnnWEQiRyFtDnLtat9zpVQx1XDJw+3sx7xIKMAaHryE45y7Gj
6GxGGqSr2MVzrimA8uu9ebT1Z0ryQ3F5Awsh8AZxeITma2eIhFlkrLCMpLgJ9Qyj
S6RRZrBTrIVgS/TDapdqR3VJbw0tYJhzCFjJ6z/RpUKsGInHIHOp+93wfto77iDh
lZTtPF1XP3aPZiH/lkfcIBKeaOOVMiJdoDa5bL6DiWBqyGAixJi3icJghbYeDQMO
ZYWZrufwUEgTMWDfpa9D8s0OHf/dTQ3xkhq7nOHdQPqnxPNpDtdeM3hnZ8BaOHL9
L3PV5MHlZEALREdG4/Us5GpIi5HwdN1GernsxjBdLXa48GVoy+QQS4S8pFn/t8hw
JYB1Jjp0D1VDZvsxk+Gbb5Ic1R5qtGxLPJ4149HeBdOxUK0q39X/tj6ea6BPCyIA
IeoTyuH0yVsHgz1I0yf3GExza2T3wRn5Gqk+GaTWvZnj8i//ydI/Yxy6FTjzCBMF
/lER3MUPyVJZK4tS2s8FWnrRJIZFLLu0cPy5urB2bvqnZJJaJDo6/9hzA3TW9ouf
A+PyfoyO0IPgAHFSFucD/k//MosVQ+q45uRYZjp+Jv9IYKBC3T/f5buTYk2H1v1g
aaglvjou+P8FRJ8p4bcaKFXAZWlaJ6pfA+FfT8KLgoxnNy5FuaQX7Ax6eboLIKg1
+yhEW3XEkWJE1iRkK1gulNrByCelVZ2WKLbZx4x2QPvzLtt2ak1p4C2WW5EU9d0V
TBOzTBXPvpwMUDHyxlHTRgoDeZ/GGOBmk+ZLsQflK5VHOqbNTRfOUxCI+BQiJICz
tSMVlCEoa14KvbbE3PAtHgR1f0UVN0+EsVT0KnpyVkJ3uLd5YoaUDckB4OF7wnya
rs99gtAI8kFYD2yakT1pOUb9vFO5vSL1w1x0fRdCBQptKLvvpPnaaVaqpI9gFj3r
caJjL0z2pcsM0r59ZQjBeSoy29uyWYYFeL1scWFQYZCT1GtfcHNHnStU2XaPaKp7
jX0ZjGj2co8MlyAaQZWmjgUbvj1Wk1qFTjjOB2oYD9hic6h2qn1F/iRhwfibDivN
0KMf/jfRbbBjpQuVRQu8PPKeARz+IOKnrDWTcB4zXiLwHayirGKAmMUkwyXwsygh
2DdM5s6d5ALNnQDyZcDPCXTfTjtc/JtKFvVbEvEZAe7Lt32YYojNvAmMm22USf7z
ua/MeNdzomd5+y+6U5LWvC0K75red3AVeV8CnrOoDum/7RtOcOQ+721agbvp2CxJ
W979U9xbWYcc09QhguBL8HvkMjVopiR98/dODLMiKb3XMxPnvY8iopGPSkapIULq
tJIZXAWg7oOhAPdk/Oo+MeXjTJPZhk61KuQL3T87qslaQPMnR2ZfM3jK737hgXa/
cpOdQXWy3ZHLwokkx6qBs2GM8soQw2XisNH6JzOGeHjs2Mm5xRmsplE5ydZvcjFg
h7dE/N3dWuQTptNYJsBo7qTri1w0XFVv8wpCh4BRt8UwzmIYD+hXQC58NylwJry4
mgEpxv5i3/SOBZAynbYQkEXXdRjYzRXKJvXzH5ygbm2sM9NRdttYa4AYL9wNVcgl
ynnTVsRTu4YnG6Onfji3EwsMsU4zAEwgWjWtjz/ZeHB/s131j+xsVi4gCVX/8bx9
JKL/K5OaogLHck3PXtyKvKlrin46V5Tz9zDL9NTwu/kEafC6kp8nwf9z+WKkDpnm
mUXOtjFEvwy/CK64/6xfM8vid9WDKUMjk8GtcTxCOix95oUBPDNaLVCKN4rTKnM+
SgCTV5y+tFS5rpGmGg5kIix89i8jcJzia46d+j0Z4PJ9zIsodqTJo4VPt0SvgJgN
aqlW5ipo5CVMnijMHKxI6PDuzeepy9FoD5cLTDDogSgPfLI7ThsH9sluxCzr3nIu
WISoJk0kJtjBRY6jBnzJjLfEAcEutJfVZvLSPAsskiN6XMC2J2YsE62jvYL5e+5z
p9DmgmHgwLfRBQKFvk+tXQAFM10ZRzEZRod2/8zQoA0dmpwDUqsHn/9K2vUfcfnR
kPvYnSTuZrlIUpK6KqMAOP9D5xHG1QihCRtI1DHbaJxgtzUvH1VFlJKsb4pblR/H
lIxjby4E2JsXiHZChpcdJ/nce+1JaZ69niGMo6pxcMBdEmQe8xf2osRFVftOQw3U
T/7OZaczVv7GYdKk/8TbWfcTsUv79Ove0VUtQG9B4pBq+RH/O+m0uj8swe2c0tOd
CV5yjMCx3ICpYFe4pra3kBnWAtTmR9ygQNWZLtO0nDUl0fthlxX/4Ah8RMK04A64
1tgS543bcqkTuGojJWATYpINXsoBioZ9+hjfKpaZkSky3QEq78P9dlH820+UUcVR
g/yitAt8FZzrfWC+WoTJnLRErQt1Lj8yCBM9oJyRhOjEWyyWXnn07NtwHdAMkNt8
l9h29qm5yhVbFhiKfAa0EgS2lD7OJl/Crg+0BUJOmT1Qv1JOgthBjDp5esbhhmOW
6YacqyAvnVhJLnRq0PBOo52riypW/z5gh2ponhxQ6Rje3OgpzcHKEC0Dp6I34mXm
b/SPes3e/cKy7TA212oYzEDRVCqniNvAB2XoeOhdFWY9/EeO0mWivZQf3d5bWUqn
IUhtqlW2sCDO1kvVbNxsC+pv0juwHOWQlgdvI4DoxLopk7vUtcQ2OdbOWcw1MEik
LXk+ea6ATm0B3VAuRHttA8ysIMEPSWO7G702o/SsOFc2IrF9BUAC9wvi4Rs//ERE
SqfldWQVGdj5udS8Fbl7tGF1g2qK4jCVCzfwn1BO3p0Ykzid1UwLF46NRI9YPC3E
6m8J8grUJ6OaG3R4klKdqU/JzetLbO2mikpgyOWOLGCH5L2Xmq0/4hxDeO/ZP192
9aLimmgjzxmyo2oPBhEmJXSIaCL/kaxAXdv/LzMrpIdua92nTqLTcacfk6VPWr2n
+D7lgxj2LtkpYmk0/f5O2XvKQDa9Y6Kl3VDBTFmi8puMdy6OeuQdD7HzOQdOnhnv
g4MwfJ71/I4wA4OvGNMcl1sFidMffyFUn1lyyP4tK7D8spvjK+zn8l39qpplS81P
usjV4QLpBaoL9Xz7FHwwAGhTMqR7DzWmu9ZhB/vqx1dmQKn+6o+fm5lTdDxJnYNN
vGezeUUmCIrpv47J+WhkHYZk0ZD0H6vkLeh9pytjMD+W2ITOHQT8Z2eWf3sjz7TD
HL/lezK7ePJ7Mj2XZbA/4zz9a2kG7OH0KHLo/Wkv7Hj5TpeexilXH8rDWo45yorF
yD2M72FzKSoIf/o5w7BpUvOf9ABXeFxEmZnLD9fhMlbHIhUA1qbelC9ORw1pFAXx
e21GGyvYvZJMyUKscVHwjUD2DWY9/cNYzN1lusiSTbnU/nCYiytDf1lXDmeEK5+x
fi/x9fMBSVlkO9773lPAadVX39QlZur1JYd3lrS0OS8p0UXKoifQRv6til97Kr/x
LA+r0JaRLaVjlm5/MHq+0MQ80OaH+EKfrq0MxjJ9YZkNwUxcnyZr3A/g20XWrnu2
z3aKCaHlpoVXdlq/XvVcWHPNZz1wx7sW5I8Zr/OQDAEe7dFtU/xNupst9JjLL1nF
KkFrDCVeprItbee3yl14mnTuiqLHkdPCwi7KkLqtgdscZHkITz6ZTgz8hDZQKz+5
aJ0D9AUXKTzscTwWIkfEeELut57XjlA9aifpS+evo6ARIqNZaIkI7HjlGy7bwpNW
oB2t8h37E5J6sz3U1acj0ylT2ShRLNdxDTe6JN/9D+SNlZ4OUSYfksEJNMN2/4nU
gRx2DMZmg11JbpBVsdwrX8G8iIPBdyponZN6g5A9qpd6Pe30zOciyVlPTO7h6Yeu
IjrYVmk1cIP8q3PBpA6AvCieoah7HAzruEZMG6mUyevuu9SUn6vT01j2nqDubESD
lcaPtavq6LkQsiVUFSauMvojAe+9EL2jEkFwwvmjM6FP+YSHLhVy4NXsrleCruUa
E5ZKIxki6x/Hdl61Z/ACfOAog17DOZTlbIN+N8ZRnHm0u4fxOxSTWp0+nkANv9oi
bJEADrh+Ohf4HOH0A54bHMnokibYU/vPFKPmKxYQO1PN+ze+9ouJG3fgxr/CKXyI
ngKRXuWNcT7zJtQ+I30ibeLuP2lEG5wYWjlVa4RIHU0sCFq73cFw4t4koyvcp2gs
Kh/8ZM1hv1GTDsGTLn6eDv1PjIpIpDecxaIvVc3A91+u4tbEN15FG6rio33uVW6K
GpVIo3KR6aKyh9s1srVVlvKvwEY0gysuuSA9fwsrMHWszhG1MDtr4GGBilObLXpV
tMmn3jIGefaeFsog4RnoOw7ndLZcY1smIqN0Rt2xdKoQYYy1uTSXUMbCrhqcemap
+gp1MZkAHoUdnPOljLiCAyrjB/iGRL/R5YsW2SHK8g+Zpg5B4Fo5XS1x8N+fREgO
2mftLcXeV8NOtXp5MCdaZIhFNdLpLlsPkCHB3QVrnP/nP94Ewz5YFygYwN1bXSKK
s9i1gXWFYCKHUkRpRKmqZYNspl9OG43Tw8Bn4Ymfm/hov317Xl63QS0UIA2u3Rmr
lD61iI46rhpV5oLa6/J/QnS5ikjUhhlfMemn0IZMCDiRLpGHMObeFUmDBUKG4pG/
+SV5h93MOglT0140bVOvndvcAxrVSlF483MlON5f4fMvQoQIozP2wuf1XNc67pk6
M4lwRNdeSd72znPO6NyEkDqZlNgA5YzG2VnAG6IX/xcdjBWmCXg6vQz3iag0gw8E
BxagZkN2COXsJ27UA0fCo5hyazmaYPxb4u4lJYp7YVXtFUFTzkFcuoHp26CmkFmw
jsFy4iJLtQUxu9YK+aTadWBYT715P4zqKkbPB01EH88KcVuOdG9AiFKkDoCFpAWa
dOZffH7C6KTiANkhk9N3J0+poOIGkQaCFa290c8Nx6UwOYrNS1kE/JBQNps26zPo
uY31NuW3NajqgkK9mBlMHS/U8gtrLZKOu8+yMYo+P61hMppAhQkH8scwzVBnkHo/
S2XAKxzLDarTKLJDCn1aKroQleXoL8WXeyNjmkTVn6lZ4pugFEIS6IW1vWAIYVNB
4Nv1pmDJYF24gRVZVxKpjLmoFQZZ2YIKIlAWDwRRsUFgFEDIJ/Q2qXTxg7buV2ER
2aqidibtmYlGWY64hYzkwB3y89UB9wNXE6RBWqUIKWr0czGjwkTHXN8IqUjH/XYK
WKXtf/YWVSZexMpAjdkn4WFFT2E9BjyBE9YCWeer+MbZiXipoOn+Jq8ODzGzT72w
XpAYYBaw/Ixxe/dbZuvOP7e+QeoKTlLuFrHssjQtNRGpgLKY+Ma/ONM9xZLVEAJd
PsTsMylNS7nnwtt5JsDMHh33Xad4feZXIkaB0Lq5m8uKIsDf0L0y2OGpHwkgKF2n
wG89dtCnzEWJeaPButmYtmAaN5rgzAkLwqdlDdlP8AeU7A9GO5BSVHNXHMbF33nN
Xl8Txz6EYmuQ/EoiZUr+IvQ49w5fyh2GdGuGh9HOy/hX1XTcrlqO167mFW+uYrqM
Vf+zsOKOCREPO/GvttHZtJ/x6jUWra8wl0FM67v9F5+iX2Lkmg7q3Is6Vqqzsxj0
mML66adEAI1rhQH0XfMGBAmXmc7PhWFyRvvipMA3GrIRJhSdlau4N4Dk5ea4WrPU
GKU2Kt3CAkpQb3iSU9M/duIGlmmfVUzVLZBVaYchu7Lc6JnZXZDYIZDrzgrGKO/6
gfO/v8Hu7D1IhptBbHmHogZHNTqP4a6IsdeCviWiTHy8Rzae94g841v0+MjZ4sCd
NzFgLJP+lKQ03Fi95cSINmVZM6QSzg+OJfGp9kf4CswVmOI2ZD6+fyRW/fLTe+pO
vQV5UNhDpHQ8kpygb6fEpOlwpeH9G+v4B62AGbpHS5uFjAt6UkHoiawtkODGX3h+
rLOnWAYgvGzukvffRT3BCqIEXwIXGvQVP9KQOmmrg6mRVZrZaTkeV/JyVSVdMZLW
Q4gG6ahvqGguFiu/ExwRQSO/dBzHioVEhzeJLrwrwwve6rJ0aS2pOBTw2y7GAjlf
as/c8gapyPFLoqvuq/1PmDrv3rBxApGj3EaJfusLCmNys3REtsrHOoW22RLB6gvR
jgHX/L/2NqlYUM1zpDzlaydWE/bdB/BtEp4Ax0LWA1/AubqA1FOO0eIGEphS0ldk
gKfXE/2pc+8LD5hJ9uL9nAKC6Bh8nhJoZLC5qaTYs8YFQ1Us0MAqPMxbzcG1CmJc
XPfL1LnjF+OiqbrJGAb15Ss40RryAqq+T16fOP0p/p8uhutm3UONtGRVZO9t8Fiw
Aa0i2o+5Pppr7LwbF2miRM+RgLMZWk0chpp/rd+ev02V1LJRGNjicZGSeO40264f
kLEpVmjhGLIIA8OWULdpa32jbFBKCSFSX2Yw1rTXXHx37Dhadwj9Qs76z+KU5RNo
j4MJ49AltaJKdPDVmIv3JGKujG8TG54oWosElEC80oQPmtzcna/pKfY3PqpojCdv
ge0vNUzSf3T7rRH+Q883w5lB8+HOZd74kbzz5EJbFp8/w1Ppox4neJiTyP5XUy3K
x2ylnOVyWy3r+4hYfaSA3zanjBYpW8dtuX6J6s1FC9f1BjYHdT8+PzD92PF+1/sz
a9BcxJVOjbcs3MGN1ZiMQWnAYTRGzPyGGrP1MLXIOnImkm71iztw0kzDzrQtggty
v9Z0JNAbzZMk6pkBmZRIu/edk6y+Mo9qRuslkWCApGgjPNkZFcgjLg4VKHgReX4v
kQi1a2i5T/voxU3g4X1tHhbCvWvqG9Pv18BTBVmrDWRx6ueKR5pYYIw08To+jtXi
yKJ7vIR6I5p3rkS+0GoqyOiAWgwcrACJG4GjqRKN+dMvT/Oz8Rw6OCd12AvP4ir7
GocvUWZLdED683fvQUR9nVs3X06z1QCv0cxSn2guIbOboDYteiDByDzd8y0hthVt
vxgh1ZrCTGvpB6hEO4ud0N1FAi7m+1Sd2KDl/c7iwMc/wCR4K12Cked+pyowPZ0I
sHnAri89H9R90rd6PR19Caxtm/9wjPl9KsTnPriW4O6fqIvCXGpHTXihtqziknu5
vCyE2rCnHioPhWI8jlvGqefsoHipDGOt8/ic1bKUt2JkI3nMKVFXp5iewgY63Eh9
FecQq8NHgzO+LrPEwXJlcrTEH1PmNqZRNPnJgPXY1j3ZFd3cuJNeNJiy/kKsZcAW
ICjIncAmoyK5DzlH0yGBpgb4uM8b1KXKCE5NW22yV/GsQzXvX1AqAVMhmETmyjEh
NjBx5gYXusVHiccuN70Dk2Cr3ctDrXXu2Ulc4pmPNzCxXakADBreEjxjoxOpKTPk
S0CWkmvwdlFy8410GASwaB9I1kuiD1SXNNPCCctkn2Pk/kv9EUgMFI26BWitty9f
2LnqZoZZ3/6EXTomg7N4KJ1jxwr737MrFgWKuW79dYqj3OGDu4zwqV40a3li12pQ
Jw5/JllX0CtuysB16oBHYvNphEewEwjXGDfckzY3ro2s7G0zA6wuUvXKWjNfNp+D
AXPq71wwdWtGz7xzMz+4yR+aLiqo8jVJphMbksSgOR0ZVQaOl6LdqP1Z+scO0QaH
SWkfcoyoyaZhRWVu90bWPkcuLK+h4ippPX/aIK+QG7QhRBoM1h1mEBDOVAdmWPWU
56tn5Jt1l6mMDEKnnfk7QdNkf17X2IX81xeZAwsr5hdLLAgCxPZnACE4pYPOBS28
O0727b5I1KfWDTEKcHKe7dKIvxDKTm+YQKUyPlg6waZ5EM9OXwW/L41S5He+atlU
psknZ8xcRm+cEvLcvrSpRY6ni2WaEVK4NpKz2TIdfWIhyrt15D+g+nO6Onl5hn7E
fzMkttki2mEvb8lXvVNa6yAD+oAsHjQ54T5kxalHU18RGU4PBtb2Ng5o25rSAC17
nCbMmbJDXy252xuhSbJKP3K4JfPSyA/x7X5sJFdCs3xaoyILzu50m9T1H3mKrwQm
5EJ2hLS+4z3H0ZLDU4QPryudZHNF07b2UTdJTPffyX/BLm311rpAJU5UNuKKrf5c
qvzvslD8JmxkWA37N5EnPwY0HrRDf2ThFp9j8cO4cHAIdJY58wPgBm3sps4lE3j0
cq8uG+AwhxD9PRxopbfZ/8Lj6UUFflXRr5n0wyTrswYTFBzT24CUQxM8rc2Clt36
d/4WAr73ULNrlOtOTt330IgssQAXAxf6/RUDhJmsdHpD5y7ZAA/aYEa7FSinSC3o
Obi2Fi9kO5vvSGUUkTOjdnwfAnaaDM//qYROEtc12lKAQG11jkBZBoQt8rRMrk7w
JctDN7rfe4huGIxhB6i5oCp6D0e9Y+undbiRVA25PDj0yS+Z95s5IbHzGt/SaTSI
3kPJQCSq/4L+q19g6gtysp6YjDgDUgAKy2QgFnzqFBxhKq2hvFUe0s7FKKGR6aIw
rZ+RWUFmrZJ1W3dgv1fOBpoPG8mqTGAYCFnFaNyn3/iiW4dhO32WhfZoRdrJDMLa
h4bqzOWa2qu/eVBGlGRDujEg45bwHg1r3CYzrF2RGg0wv3wsBbxG0ZdVPkSpEfk0
u6mZ6EZMdoJ3EFV8QmyHwET4mJE/eTS5t/jNaWnkDIEeUbssbm1lzKLs+3mSAt2V
IhcyqRe7eYGt1gMAR3lhoFCA2xWti1T3cSxDudvhid7QsAS4QWqbc5nlVLBqcyM9
Vw8zGuWdX+cIo/H0+fq2V3DrFnRhWJGR8vKSEZJK2PDvU7iTwotYs/a5l+G+a0lj
9uIFKM83b0pQq5RrjSq/jQEDzy5lx+rJ2DXqAvwIxR4NIhNM8JNi7eP3oOTjtbpl
hJs5/MECQk911CEcrd4VxbF2ORi4CPfV21DrH0xQsMbb7xwJQ8YnJAucJ48Wnrrn
wOqEjqY1L3avECMDR/nRqsZjQBXIXRlGEGMqtgerItYm1dRE32AQ9DAwAeH6YK5N
rZ43Rtx8kbAhSHR01ZI0gy9GMUCaW16OCiivAJ0Zw6ilVWhMUspzvmPYnCF49NuH
JW2EmZiU3EZCPvpdpZMifAICzJAuq6X2/bdHiqTuTqnuKQDQjCqH7VjOno4SZm1A
xEDVscz1vFkkJ9eAlpIFHlpiTI5OZ4aIpXLn2mdalsz1YfSpfOHO8Kzow+m3WUym
V9OyaD74RPH5xrjLzcy+X7hRDl9m8TLp/H0Ei7z4JV2+nXdNpqctz7PvxNIy3K0W
naG7RiccH0rjs1CCs+l/lKq/1gyMQoPZg49g6PVqwapLZUP6hAClORA/pZ0g2J0m
+VpqalVjZ9XebsRKtpzePtWSZlmpvh55FwvGiah95x2KHxbLdPxqjYNjzpA+gOZ5
O+u4+ezzOwK6b+Y4fmfxZcuKwAhdbhV5Ny0Mf4xx4XjK/qQMEAmHnSh8rYs6Oy8i
vxPXBE82Ab5odQ2GXZZyQhKFAvY2RRasm9s9dT7vcuYakofeH2aOBJBwuCQEGF80
s931hg8Ndo4EfAJTUu1J2ghYXutO+IUpo1fg0mbA6kQXoPwLOLkOBuO13ncBMJ3L
xKpjeIykpuwh4b3tnVGd/gnlyYPeqYL28XA5fSlIFJz94Y14Y46yOU+lteMvKYwq
lrgpO9Nplzz1cAXoaDyQ04DZIrSVHSotHllSlxuLuLKvpExzJVXz8o+CD5fHBbsm
S027Z0/V0XnVY77lBMgzAXJV/OQWE8j+W2xYHfRogm8Cxza+u1RcxN4h9iqtegx6
BY/ZmqcBR2cdQpxn9A5bIkBBP95Q+BEPrYeZ//Xpbekws34OUvBGeoWe+hVvPnwM
Kw0uXi3yVb7ZbsmD+hU1pWmkrXiRNQJJoemkRDcEucg7EQZ+2h/nT8fyb0Nya4iy
15T41lMoNLaQ3mmbbyG7Rt9fGvJqW8YjhHu2QprJ4lZtIvdUajf9fiL9+iOhmqLq
R8kNEjOP3vio5KfTuaCO+hakZulM2iqIyWekTfEFoBgg097cGYhl10p1zFEIbbyq
+SL/8018LmCEs+fReOeUBY3GgDAFTYeFVc8Ll8mHM5pZ+JHiXKTnXkeiiVgVScJp
vm9fA6vybMBagSwWGGoZkEVZEeN1qLmI7OBTEj4iW6l+axFThjChGx1hsmPt7uec
KEUigR2G5uhzrc3zgCfJlqLW1iSm8Y3RxJkdagMX8gshyvF41h5soAiDClm7uxED
DA4r1DqimhP6k+rtYvr8BhLyz9xxaFwPI9VGHoVOQvI+MWwSWJpywe4TDI9Wkkst
78SR1CacDByea1l+gABKTYU4adD6QYuoKMeYahsCJU96pDYnoLKaZbMbH9kd5Zip
4GqzD7U8aleinxMAPAvNNP0mt2+ZtzNQZM/tdHalnZkdDtlvIpViQnbsfDsgEgP4
F+mJVOeh2CaQ6f7nt6+K0DY3BkdjM3mZ2xuVmwBRF6Yu7FKj7hbKkFjyY77cQQtB
VowokT1dNEGkfy2OIG9xuoET3HUDV4Nmmj/dnAy2WnvIy00KpH+t7fU0xwzMvdpX
dyIkkbAWHB7v1sEIkTq27dZoc4LsW8uPpakDq4MukmyXCkBJ6vdS6xVGJRJcq46I
fBUImHzmCSWUzIeB5LUhi9B7MYr1Pxxw/+0t85oHh/4IKRHww7FZhBT25IAEASXd
7fV41ajHRxCyNroB1YfnQ66gudaB2VWt4kpk9fQi6EqWaqjyGrUbQM0qCQia9gUY
MRAxe9/8d/wKJ6JTNoY/6XqlkqbHyrGgkqdORrBkrDCdj2gDqMrNrGGNWiTuvU1s
Cy7YtamaVKHdMDB+vjmOXJBxJXr9sfgRdqlnfZo7fkMwzpIU5RUPOMoko36xYIy3
1j1bejM6SBubWeovYPpOPDfyDLFyVHajuIdMmokIJv7lPI7U1CElT9DWpOOcy/Dy
lAz4xlhleK1JExG7i8gchn2oWAgpVfLQEskWxYWYVWQ4qEm92TCPRGsUAmrh2FZJ
VY2D8e/sHgYdXGJSZFXXP2g5Fdsi0LXAqMkdBBATq1hI16dO/8jZtV9sYJBXAcTN
asSGeAat2se7bwfQjaidy3tX879CxWvPLm/yYNMfk0wKPeHkt8YSkqGSv8aPIfwd
U1tWI5VmmE5kS2nxpHRwy1f8nLld1ghjTS8O9qvtDYxoQlpYhLy6Jhk2Lp0twIs/
JtFTXNkr6xEGRuHP4TUcIbhbbA5ko4h0VWhSHakVa1VSeHhAqN16nucU+PUbMdVi
N2BwLuLhpkurWjJxNj0r11b8gxVnv7R4b+cPro0oxYiLDASq5//zZ1MOBfY8bGzf
EGjHgCjkDTYC4A48d4MT4IJI4mj14Eaa8c++vmQ2xMwWO5LvxRQLKJte95quM0LX
lV6HzYQnR6sdn8PeYkFVQAZfpPjDh3jZKxJthzoEZ7ev5w+FbVzM+dFoRAYSLFaH
XKqwDSy9UaGyTPZ+dtM3E3/uA8lCHPzS3npANm5hDyRFzVDlBcKDY92wRWsNw+eG
vOUzGoyp0CqYjZadiWwbxZaD196wIoE7PnOBH9x/RpSgqhmAbmcYe9IcWylLoQPl
VwCXiE7Vs+aPueaxqYIx72qCfp7XY23SqovjWT8qheRbwtntyGLeIEmr6uwg+qGO
1R6RU5EHbQhfy1oVnzeZkj9YcwlV3SrIXJ2FcJdMnJrzeGN0xuQ+cUbSsvUqLn/7
rvMDF1V7wd6A4OGm/tcrMJLl1b7pYFqutUg8ltrv5Vc+U/MWkZ4RzNDWcHbPTpRC
B//Im9phbMpYqEM8F8EbUENWZZ8GaF4rTooglGN2Jkbi8HqzbfwuTYnpD+SLqizS
5rU96f+pDMrjgFfJNgkwR/YKvBh8Lya3eAa5Qd+Ap/QbsaATDnSvOXsrC0+VGPl7
R/2hP1v+Tcobq/1BlI0HWXke+NiVjZo9zFL5LLKKn25GPL3muruW63v8orZgPa6U
pto2v4AW0Zz+0SkYg7+laPpzdU/d0OV/NBxmVOve6LZAM5rR0/cy6YmlZj0UNck2
U/k4mIdecM7QYpWl/GWTWfyeRS3Qi5rLorEWN01vgCXFsUckQUE2zPoCIyDh7M5y
BNV/HTerhRRHEKIguMbob+YX/wRFdz/peH9mwOE8JN65qQ7XBclAy030DTc5ZccX
C6RxymECkLlMTWVyMGYhsOgANRMC1cZIsSugnNBv+ChuSxODmY4AqM7lQDcpDuwf
4BoG8J8uaYffHbv3b8uSjvtQjksAK8RdFvA5J8V0gx07K7uY+bKmnyNDGHMWkZJd
xM4T9lxsv5Vdc5zX3KPHqixyvJIpMBc5nNMJnjEwwGDcdIFFcuQ0VzX66A6M+fCo
ssBuiKo6gGkdJuOsAh2nfyjL5ZnXK6TAcbJFN3+5cDV4rhxcGU6NzO7C5RqyZMIf
KdaXb2VSjLLJRKaZcsuOSth+VBzRpD5VOKtIIvQ2ykE9/4dQ7Ems4QVJEz1X7OTx
MOUEj05r+ILcTWZHtuI4l7xj7xqJ6TzFqpc6JP6+U0dM01T/k3iXEaxeo/+E3zIj
aCYBI+QwYjuEWfp+dzIaLUF+UqFpVdAaM9EyqbtMONi4h8GfHUwEKQApqmRBdqk3
PVMkJSDY2lQpCZq9ya3R9bUOLw8VgJWV1rCSowj5lJJ7nInsmkgPJ5GZ3v7dAMXW
6F/vQI3FclsiJmqkjwwOtKGPZq7qWJ8m9apR+taznsXvlMRd2k2Nvmqn2ddSBrbX
Dnsr2ckkKNy4X4Z2Xr9byM2hZSCvDzRTAd2qHEL/MPz+IkcLpqMWhvwWs4w7rB6E
xk0FZ8y1VV9FXv4HTTIWFcDZqNElGeqWZoUB/SyclzCFM/x6BDGiOiyKZeD1n+oP
xnZzGsRxnDF5W4xH0go9+LoN4NMqgF5mlUZcTj+0sfdkgcjHE4YJP32Ehqwgn8VB
36hwJCLoMzpGS7tLLgxs8brQrEZMPiBGhxXvtbpMHZfRZlL+2gqL4k+q7fqdI5+z
c7J/YAbsvL0MnLulMdVLJPuIjH2Na6/TNovYGwIcShVgJJBEwGG570mF4c/Zy/oZ
yBb3S2TfeGMhOG5Je3emU0rekURRXxl8YzrrMjMmLoa4kupIFKTM/0r2fT4wDaTB
K16O/Uqfh9wSE7qZNfjsXRhPlJfl8LvoXdFEhwd5w8OU5dgc3YAXj8wxY5rWmS8S
ipMVo1kFWJzS9GrUNYZ/0t/4cvAdeCYzLEr4Ffchz1mkDtouJ7ivXbIUExpOBv8X
Kt+H68iGx+XXwzGhX4VqlcZfcl43KHeYVTx5RfpaDMh088EYdiMVGxFLinImDk+s
kY7ZANIF7c8qqOHbtEfbERPIfxeOERqmDX27yXC2P1Azje5H56W0yxXDtTYsx3iQ
jKUXqj4I59ihI7tN7ZTB8s6878/sGWYaABHUCySTsFj58hjMDA0aaAWA/587Ul8w
WDf/Z7ayARjWV/FJNylXBWpDrGnDoW9H15tXcvzRMJtt7+SP9q8uiGYS6iS8qHbX
4mpFU2Q+qi8bFzdVsm71eHPUSwJdOQ+tMVTcy7Xoz3gvnzPaUzjf4mPxmwoBAk7K
QH2T30JC1Cl/QbFgbOo0grhRsvLUjKZWVfz2o+CINCCdT+Fw+4CgH17IDqeLk8sm
+8gZ2BoHkvkAa8cNkVbdKdlvIucl+GSkakTKTqQISpPhYzUFR86YJK5Kd0nOQGLH
HzBL7BtokOo3XCyvmLlpQVys2zjeq1h8bt4LkFdMXrunRWVqEZXCdBWdl4b5V+t4
W+64dIzZRoTB3OPjq/UKYoAiBqS90hfuY+XWa5ITrbau7lWtsCMPoQlNUWYZF3zh
V4/CbFZTAZzvEltOQnmpYd6NWsCEqdXC8vGcTXRlfh8B3HWvdtiASWFkv1dI6dre
cMfjLUlOtc5UP88f3Sha816XnmkHX5+xc85FuxLfyPS+8i5pnMg7PwENmR2sa0oA
8hiuurnuLX7KqDJ9MP3TIuaFG1eYkrviq7U8n9gvC9OKK0ZgjgngYCx5Bt50HErx
dDV1mykrS306ZUttCTQLLiJohZO8ClnbB4Jh13by2r93G0W02ddK7fiItIfk6cf3
d12VdfaMGgRyDJ4fJ236VG2VDgrQCFhZTOZDYPZf9hj8OQ0ZFiGxo2te9vGAIkOV
2fV08bBqGA8OFuI02RxsVPQfmVak2Axi/pxEinqvKNtc3yuARr+DVi6Umidu3Yp5
fQK/nwddQxqRKLwjNHc10TxtPFgES+GbnorL1lF6gB0GpBv8WuZctkkUecPzc5HH
DFHKc+zXX+G4ZuUL/p6sUBpQ+3be5iyXB2Do62rzqVqyg98HW3lhwQkzklXieogq
x+gS9qOSx1HOWLc60XbaWKLFaGntjEFxGP62DD/h0B9vCAy26MWOoFpV+/7IhFEO
I5vZHRMcSTx23Ks6hy0aaqBrDVJSeTOXNA86fs67sXjTBSHp2Q9nWQdFCgbIj57+
29Gwu98VkwQVHIC7GvM3KtCgYndtURYJNMZXKTcIroS1lIgqEzghqDG8edahXStI
+Z4s6KNjNurDribCLkqtHx6WQ2YgZp47hxojVuRyLi/+mSnDZgGqmJu3SRpn7dgM
oEbL+1VjQlzyyQOfug7RxrpmF98mg5oP54RL6dQdUd1pa+6G/Uxccdcf7tD5siYN
QMqdjXk8fhfOI2CuWnAsc1hzgodBzRTzAynaIzX6YTZxs80BjzuRWDmyCDOPr3/H
gYhlG5wUYHz/28HP0nW0OhHXkS82bn+wsNnC7VvR22u8HGKxdsBFdQnuYVbeLWKd
sv2OOBwMoCgo7LeYg1zJFseudcbHwLiDSRbQ2Da47s/xuC5pLCl8VjaAv/o/UcEX
czy9Vf1rXhiC2B8J2KticuurRpVnpthnY243gD1NnjUULT3KUUe+PZPWzcJcHJk6
ItgEMXEXnVBzR+TzQfiAE6FSJH0WlfD68fskoP7jo43noyaL1r7HUGnEFC6LOTTW
G8l9nOI72xP7e2Nt61uQdNEfP4shjHHPtI6CfSpwfYiEU9Rzc+p40r7DOdrADuiP
izkrcNSLE4p17MsFZPrUxLCeuh1LSgE7cDUgBh4ArqCAA7c662+dvNkbyA8vNh8w
Et2lE+BxTV7wOiNN39hNwtPv+ViqvSpVKPnLRonltou7anQX9nEsZHu4J2Go/0lH
4bdXvDe5/wlRcjxjj5TnZ5IuOC00KhSlqO+UN/7VX4wdQ2+PjQEnjdTsta/e8bmH
TMX4GURqeioyTXMpmYAymDG7hMZCbM21xx30/vFipf2AOeR5mkLNV4IbHQ6bXrRB
xmxo4G2An2mmh4DhHBaDA4SBIi2KvNgTJ/oKsVSrc2+Iy3tY/sB2ciXDTrgUUNXo
03Cxhvs6ua0F4JIavd7cyxTVaVv2W0ivso24CVezTFC9+38JTm5CiM9LjcOqphVD
mz30Uq3xEwKvlB8hc9IrvFHNOlVaO3S/gripW3jPgYN2smWBYR+dl1LKsWfBSQjh
tk2zvRt3gnlHdDR0DAWm9GPEkYEBk+cheKNfFZ7yrRqK4mSRJNnJ3LaiTBaVifHP
ltDWyZab9sBH9w+4UtAYWMQ6q8WxtN/mk/2FcXK+/TbdEHbPnEc17OPiDHM0zLh4
MIdn1tw7bH/AwnPjIpVySfkIqXv0C1vk/eNVujLRixYpuXn2jrSzsf3BtEDqACAA
w2F5tZW1Q28JmqqFc2kgIO+n+WrRacdkyRzOlfw3IrDFQ+yczk3/udFs9j76ci2w
opM+LQMNfinipjJHYJKlCU5iEXon2y7+AR4VU3rmTQWQ5jnVW6eHG1QkKsk4sUVN
ha1OC36RyMmQsQ0NhC6xbRtHLVw5jNqOvt3BQ9T+7/FGlilLWGlvcFyyrgsU+tCm
Lfz11UNtMlRYk4rCsbbx3dDn8/aYHlZwvipnyHgNnsqgj5P3JgFQ7SSzG3mu+z/e
qvZwcnZsO6qXRvjszH1ygfGLZ6T3Xoi6+X2mkX8inn18EWm6+tvjyuV3Q23yVV3l
0f7ExqaeDyFSaOhHaroZdZZAEFyeXqd2N5Ql5+7rDIncyNYGPNFXrUoU5PSK4Jo2
1Iibmy4cd2mxYCQsuilc5NvxqZW0MhNhYQ6FeoPDLvfvYVCBpbznZiEOdlyF1cUq
EjeUqYZ+9PSetesVnr+b+4vkCt2iAlSFWSXtkLlLciywZ4HHTDD5j4apoFTnuACk
lwYg6bna0krkHo4MK1Dbo9qJoPTYeENV1aNgtlJpUaZ4mROSqm7BVSqzqAKE2dv0
pkBsb2J7YUipSas1ohNxPPFyqz+0EuIOweUgHHblBNt7yxd44wsrYpnU8cSHBkl1
cJDy+RlzJCgjhA41zGmNkxHX6M8bVqzTwyKaA531cg1DUSbMrITobrTtDu7wwSxW
1xtWJrqEni6AkQuVRDNyHKhhdRIs5g09if4PvhxtZRao5ZEHfYNF0NIDobMSA69O
fybZiY/ZQfC9cus629+YgDgDlyWnY05OZoT9ZGg/B12z1d6P7KyOT21n5OSmBESI
1Rw9Oegl/tE2Ut2l2APlQWWw9BGk7Bo+RBTepknM2DqhNWvgA5JN8jD0TSYepRyf
TPpROCl950TxPmIbASCxYDhhKNp0LSwM3mGswO32wT6HYuxfbbdDIZgvk9nnPdNo
sB1wqSSfiAb9wV+l7Cadvq6SRS4+VEMlV+wSCH1LgPKadffr7Jh9SMyKdOGxD1el
6OYQtLyuRxTaFVgiTP+jyqUW/l02qAjEHc53jiWryBzIcI30FgtGJaplD9PtAG2m
1YftfdfGpIAO1GzvVNgfbGlrOOH3rjUyuLqLP3JQdrbpMdekaV0Zpd0YjtFDXTqQ
wYVgJFipRVbjJsxPajbo8eKXHqLuksifNi9ficH5/5oKQ3yKMlcuwQcgPtorq8/n
nwdrgfmC6QX1Ukt2Gja3kufuUj1Pkqi6SVcHbCsYOozHcfA+wqSYbWZnffksQdvJ
IfRTGgfscGVf8Cv08y8ICReGfgoOnllwmZe8+ib0dVTGqrrCoOX/fplBOum5rrEu
0AB4a9ZqseBycFySe8njr+MMG5yCzJsDQp1OcS3EdCwc3r6m1wX+TBLrUhKef+b6
sE2+if6RtGK2UhTuuQbDWhWVW3NBpgAuh9gQGrxXMOnkjni4IMh2BpnwtbP9f1ie
OlXLruNgRKSUMPWVOxTUbMcq+hVMXu7cAdfa/+MU/x9GuvnQsuwUdhlBVSKwyOKb
gLqGSZa54oixzb8dLtfzSfa9i3XsTr6Hz3TspoRc/RipyUWub5d4F2ZYDOHste9P
23yasgtmphN/EuKGidHeIDYMEnW07V2pUMAmez9HzgCpTTtkWuyB/5hwLiyVM/wW
7zFb2dAZN0fkSMLkH57GcFQxevOCVQJ48NNu7TFfVSpprcgqFt7uv/Qt1rK5hOvh
tGGQL3Lbsc1nzGb2Id9Q+BvCTY5tYsmheIn3haze7WGtf480/RdvlKSN1tuLLmc9
zOZOhxNUsK2zJgJvcCFkmmaxxQFFPxd3le2RuZR2A/Twgtuv1Sx21He++MgfdnJ/
AacBzc6XQFOuOtN5UjhL8ZVSVw8Wza03bsCq3P4w28Tw6HnRO4cO7nGqWhy3Fba+
XszyTENv9Y1dH0kOlLlFITmJuRwnM3+wrXxvgAqdb5yafb3a6ClYpkk6npTdqx/n
ppKOCYAWsBqGfdm/kBBd9VanZCtMI5KUHFYnOfIg6AlqNVeePlqcJwH/8UO5Aks2
ijzQtLmtn0By7/QX7cw1S3XP0cq3xm9mKQOuki6qH7X9oSWuqiTwIffcZH9cXOfC
wpPlOJ7DA12gnvgGcI/rA41jN2QN8sWimHvN/bk+PU8q0F1atBjRIdQmyR0+6umQ
t4ySeG/9VUIsITtEa/WqvTTv1w39VFP7+soLwT6nK5LXtRzBc2fEUAZKR7EmgAiJ
0JrX6CvGMXETFm00p0QQfO88XMwzCJrc9FSdmyJok9K/pLIP6mX0HCsRY3szeHv5
+yDqWJuAH1wuXsRzvZBcY9DxRmwhITVAeJHFV3fRaGZM00bV6kEwk62ce72/FbIb
DT2UXBf5ioekLBbBrd9n2WUKDk52UgtSfCwpg8XUrce5Jdold9iEH5Xk4JeA6WbA
1CymvhJ9+VIm3c8FGJwJjdc0lvXrzyQpMYK1XvpSzbIkrpB6e5PWNREYl/fa+RBl
0g/unX4T16KWd8ZNHNtjSMf9C/UB7BRhx1GdVfoLmoTfr1On5QteC18S2RrFAv9l
5XDvmiCyP7j9Q3QnfMD1cvWzrK1UEANny2CP6X7R33ttcZ3QFEG0o47PribZkton
ipAaZ2HtrdKh8rjsLr3LO8NVhcNmqijwF1mv02QTd4g6tMmqFsLXF6yWgz7UI1eP
mxiffphk1kq5W8F6osjD3ZGn7bnmW+Ln6YYCsRlPWSl1Dwy4QnGPu2ViNMurk+ox
GYtjx+TemnsSvJpOF7JwOvPNSl2uGjFXAqvq4bMT649I+KhR85e+iXbb5mHZ5My9
b9NHIMt2zkwywLhBr2E4eFwvKqnDaoQVr+Mu47mSoRjdzSBbuyHDkUz1pJqhPzZs
rxjT/qsAfX7SkasSOk41BhEmsXByOu/uy80ExRf5zaMbF5jlFJttdpO/PTb0S8YJ
4ajdOJq0ErmyYqaii3iqFyHI6RT/KtUK0HeU1PC6J02zCvZ4ETeRb9pK3hWKTUDJ
WQ6UpbQEP4tUK60JSr9ryfYSxpzbMsp/0DkzTPoZ1ltRSlF6CJbD0Gl/iCGLbQPk
3EhRkdaSAyGUVyDUqK0L93B/3vXtLNjkuFpDaEbU95i4Zqj3e4tBvv+ywE7ui9vb
GVBBAVAYYqd/z0eebvh3wF0s+7rgXt2HuM6Yb6UAcvpcA1XfrpGq8qdU6EYX5nJd
f2yoGu8G0r3Yr/IDdYxLvY9AOieXhui5aryMo4ubAWCeuEU9K/As5kRgZaBYY1QP
fJlUl8VQRGXQ4R2NsadkwImAVkYoqiIQZZ+nKBQt2ET72Vw0sYguNZBWBzYbLgaX
Hi81VpUuzLhd6YIoqUWzFsVuewKrLmECeSlC9k2e+XBW+EbwDTDBSqtXgLxJ6H/W
srXLM1UMJ0to+hUaFsev3BpSTwRAdOXeD0LU3jxL8Uj0YO7fRfOOiv4xTCnSUvA4
dn89KSMgwDHz0CksuxunFNhM6T46aWiSHn3xnDpZ/1IzVJJwT5VDo98C8MUk+Lqc
qst/v4d8KgH/u0LDVwC/pQxqcuK66Vrm2Uzz+SnMcnd1DvtloYAQ68TBUmUBsSrR
/JijmeQHrIkUPXu9KPkqhEHOPD7Rvu4dkPmP5M7XQDS6UaMr6iJCexOIoNdtdMTs
KmE8G0pGqmGNVckZz5h9GmciVaGT69TCACTwZAm57DuDqZRqrRNoRJ2BWOn1Pf+K
DEq8b9zHSrJdiL+7Hr3dzxFySRclsTPpOOtf4+j58uHANaUXXWINdnR10LmrbXz0
Pf1+b9kKd9Zfsj1ApXTD+T59Y961mNI/hf9A9+CJHI0TVeLMVqMeRogNLHuH6NBY
QW1nPJAcSHfOXOM3c7QUZWeyH7Ndw6FIwSZ5wiWm2oCQygeAdXLDBMQcAYJIJytd
CvZCeYAJOpllHwMFH5yOoSk7dZd5PEmI8BHYV5fDMw2PQ4Te8B4680DIYXc87XeH
gKDSIOZb+7QbmL2e1LKrtCDqgrnd0mZ7FZ3t4fdfeN1Xn3JCIroYKjzlR1phC5IF
UzeWjJpHQai1VG1V3kTZaHjzkefQaqlrisKaTnbLceSxhoKv+F6hvZ5KKoEo4Zfe
XlWOO1REuW/RsghPlaeM8wAK/7FvIX5xLevLpPU0d/PEu3WQ1PfF88JD7fbW/cnE
p86jWppR5UQKoaEvUluQS46diWB1SpsDs2gidbUvMYQUGMUGbYBRhoEUKhScCmzE
rB1oM/iQM3YpB4CPm0f0QO05Lb1CTHit/m9rvWxBH4N7jXzgD5RNTZwxxGoEpqxP
jMGN96aqWE8AsO1bEWZAjxsO4mlr3Vw5TzLNEDLcmurlEtZ8Jf6fcKXLEKZOyqpP
ILID/5qurSOIVaF6lfAttJxv7O4eDRUNLUZ9/u2tFBmsd4sdPFEPlpA+7K2QBbY5
q+om3GLyZVLZPfovDp/+UlTdA1jelWK3uLrknfqH33SCHf0K9zLQY6Bnn8zpCIuL
MprsTNaONY5eo1u7XpHCrG/ZLvUukqmKehK5tyPQDmcFQ0vxbxvC5q+aQP+SAxFa
NSB94hhoAaNUnCTQ8MelZx8x0k5osX2iJqp/0IfCKWZjSDgg++jGx+1t5QHnSAhR
RLjuVXYZicG/o++p7PbDI4mZ6AAPR+q5Lkz0bFJEX/DWVXbhFwwHnecc1so1hH4g
4PpcndQYudLi5vOsbD4yOswGBd6iLe93Jhi0LnhPtpyd+T6uopwsAlZk/X1K5DZ9
v38yheEax1CLq5XD/tCD0WFfsuWgYxMJ19e9RkjHNDHvqJnYHNZnpObW4+LbFnRB
XAPpvy/o5+RcOZSWK31xTokDXbWV/U14xCE+/KHe1fsVXJkM0to5SFEcEY6Hqrr5
PuosLtfHOymrPrcXRCJ7kE4QCIPxAqE9FkHpuw2G6KOc/9+18iOP/42K+dr2yGe6
8q2xiPU8cUAiBjGTgSRB8TalT+xIM/4+10Z5qnmG+cr+qqXmDHlJAcXiARwOEADA
sijM6B4nC1Gvlolvu3fPpRiiL4lBkHb6fd8vLmAFMRMVJ1xVuZ/LXst+Jo6kJ2xg
Qyj351h4hKH5FZIx3nsRDKCWXOrrmzU+qodiWzeqHTg/pdBXhrrLFfMilF/eI2lY
b7NqX6ou2PnxP6zfsZpg40v3DJODjwR64vD+NLT3c3lNwxqEKXndGQ3W9PCPgDN4
EQVEapDoMOtwU/r5HWi3UD8D6mYvvfsnhGOzDiB4jcOFsYp0VL4+4l0E25RMQeDL
zmcjxeaiA6X9kEZrD50yajXLgrAeLk+fMA5bzcGpK2QWB6My/qVIFdS+N2SUmeCm
g5shJw1Q5/VYTimbKG/d6jygTR1JPcuH25GHTVn5MwmPAnpCt+M3c3FLjMapNvQh
YNEjs66GdTtmM5SCMB06rEmkAH4e8FHv6Vp25mZc0xAIi3VA+NzHJQUvjV8QQ8gH
Lw9C99Evi/u52JgIasU5Fsc7gFiBIPd/iXG38QtobXsyZ4EodiH9yqJWp+lKcgk/
RKzxZEGMNG0ayiX473tIsL37ksEaUVG3rcZFARGeGALNVtg0yt7XjhRtpeC8lBXJ
bdNw9DERUaOjQSIt3gov4Lavo9biUMczsRY+oErcdV/vDui2wJdRsO1fsD7u7cIT
acAVB1e5N2pOqY1bBsdBVwFAA63Xi3TUq3WXce1AXCDlDOIvN1XhXru9O02QWMv+
KtkM3iox0eiwIcnHIxPRjSx+jXTBvDyFAfzBWSpn/3uAjbrdfDNS4JBdlY/t6K8+
ieOZmCkEPYMQSRih22AwDR8RUDmQ9DCHU6T1sdjELzdAdXf5DDh7J3hzKkKVFHwy
9qU+NZqw6MkZoL8ZoIHKoePQUVc1RFcPe9HcqKOk7KV918Vw/r5O02OrMy5ipe4G
q1n//8EwacjZA4LUAwwR3yk/0WtcZIzkd7/V3141QXSBVoZPFqSONJqF4eW7hLFI
S/kU7/G1t34S9zfKFfbiJ3JyjKBFoxkKz8V/OyN9GDIeCGB7GpZmAM3etfBERlMl
EVVGcmhpm8JLI+DUHzeg9E4dgfMZurUYWaOtJyJc9meYcJJz27aRuBUmzCv3bGaj
knCx6UopytVqo/0/Bf29txZVTAEnQW0W8oFSwnuAUppE/e49C6B9OoqGyXs6S5oP
z4L8jtBbPMTFAtC6h49ZnBjd2XCgDlEN1gtMEXaOmg/ESxO/pTtfB8ezLbenI+Ds
tvB6ivxR1Yt5TI7X6uYUIfjfSUmgPPxpRnJf1pHyu097jNC1DoOJuuKDi9Plu4XL
nKjtAM+Dauk7V+c2D37+MIP7CLh88F8V2mlwS6+m3t8y0otY3x088M/HBrkXDFMg
UX9B2XFAKcBsVl0DdGmRC1LzBumrNn3NADIOdAIeAugmugCO4XAvY6TbrBPpJjp1
IgAXATIvKUnOpGwRvd+Yxgp8xgwNldb5aW6xhNUbcKwvGiVijjfhHwJAXYkoHe5H
WQoH46/DbAtPDqWMz/NuRxaduozZiZwsCd8v/QX69vu7zLJErd39MjQl0xGXGjlq
cRGT2etnqhTl5ARmoZ6MMoPUesr4hn4rHBfcsYrAxfQDAwn08ylpPGewGIUCs/fz
Rq1i9O+9nSx2RAnvxPKNiEWJQs/JPrQP/0ucOgxZcpL+GzQluxhRSHuDlnm48pnt
Pgq2chEtbyIOLEn/Fecs9AONMvjkdN0+T5EmJ9gzLxoxpiHB5BsQNC3UVjgQmLCy
GalfeUL0+6BIiVipC3H5tRgam/Fb+iYexD/3RiGl0q/JYiT0AmlXcJ5OgXW/1r+T
mtG0OpkOIWXTAgDTmsbK1ccRSUeSituufFUuZQktDz5cwKLpQyvt3tLD7x8bXGKr
qq58ogYQFq20Lirw8D1D7tTGszwmgbgHdKl+QA/bqkMQlQXKitYd3n2ISKbqNfw/
cAwhQB8K7ztaW1QTuUqFAbvpiK2UgwLsqIgikwDJWyr18jp70oHhxcZQfcq9QVSt
qARnlxFEAA21L7aTgJVIhKMunYd03JnsllF/MecPOFe5Hl2Xm55NbtkXnz4TGM72
eqDEWZaPmLNP9p+Y+LtqRUmyANxFp/Bw2aYAPb3146l4uJvY/5SVsf9vJpDD9+vj
eQO9BGaNsKHGaBoOJHwYmuphdh34F6SVoX+E+eZJpEhx/ZfgVWVftmuwzFrOzIC3
Rp5maNIRDXEzfxgxJYc8C+NK8pDiQ4iNhbCCuMHNIyV2Ei7Us7AEQWe6GOCkZBI3
SqWKOxJRFX+IZcWKQypexW+pBJNsQuwi1nH1/HwFHJCyTQEWrs3MozrIJSoe2JwD
sE92Np63+48B37K7nlzW7pw3vOkMWy5lyGvbA3ujKwN3lC1hXHMdh/9sdhH+d6jV
ZNqf2umI7mu7L6T05mwrtHHtxLPsP2iszRQzKGqoC1v9Dqg2xXU3bE39EdbaPVA7
62bE4HmQspnY9kZeirj4AFatocClvi9aZRSAlZFLSwoN1XmysIaiXEFhVhR1L0Qd
YkihdOJhUQ6JMGSSz81sQrFUsw19T3Ivr1qJSOliIL0DbcrkkJLbNyhugS8gchJ/
5pb2FSZxYkybkNx73EXi35ZSQZxlbKn5H55ls3HlYJSjlygNEFJnYkqQTBWfYLP8
Z49HZje1bZBw0NlDhQK6bw2wkVzFMRtvvNIEWgFE/HHfRx5KZ9uDUYzc6TOSFPgC
6yzJoI1U88iOyHIPeCkShhHyk48XI4BoucjeQk23fjoM3tjR4hiSX+yNddUigle4
eGsUhepKMun0jZytOyWGAj8Px2ynUAfCScc3/Ld3ZjlNuhvqbSoQEOPdHgj+ftnp
hW6uJA3zXkARacHqLHs7zXadHK4VX/2R3VsWh680EKcvRxZ7LiUDfpwRES5Ewgms
lJv3Fz0+L7cvJOyf8rRY64eHroZc5VIBoICOj0QxgczcjDBsbx9J3Hp6yu5ILu4Q
ZCG86ia4xWI1KqKQQXVNxxF9FOd72FONVZmWrKcwS7yJ3yrVBp/eeOCM6wntEv1P
AnL8ZYyfYT5VckYH+E4SpxW/jiWa/5CY0TycP0moI/7r3YdcidskaQERUgX6gE8Q
JASU93PazO83pg5xGGrYmhT1O7pu2/4Os8DBo3dov9CLKQagCISx4NzKKRC4ixUi
Oaa8q3avjGRS64E9UTGCx4TzVDwnDb4vfFYc7nJsvD//pGh6xBaPNx2swEPCxNua
R+3d1eUanTMACsoW/MuE17erCHvjm2sQFfwiDMPZBiYrqIPAKyt6jkkwFjITgRit
QeJdQe1PcaGawWYNnF6s+Yf6ladltfSSpYQaYuzjYpSdBvyxuepABEMCU7cEriJj
91fePbvqpbOEqTjG6lryIWABQx0g8Ir0+nuJpyzqtDDKsQzsJ52mP+5UkgWgnAv0
gUI3b23oHCAGZRvqcQzUTzU2A8zDu0fECq5LtoS12TqMMDBrx/7h82o8d9lP0fll
M66y/gdt+dBkhPh4/36eZ3eVazTe0uGwO2VMATqYE+SFLnu5CJhnwPtONp4apJgZ
cLLzbDLBLZmKwDirb7q8PXuUAXSaf6bZKt7RY0I6lp5L4K+n9Y/GpnQmzk8yrVcT
nH6i6nrF6+MLhwIpyI1wXFoLojonL0Wk3IG1I3WVFwTtGXPis3k00kj2EjMMvrTq
AdYbtEP2BepyCgWzHYjov7O7diuFx6tLdoHNj/EAfl+HHsu4JS/Kj3HN7WNm58ZF
ZcZ7CTf5lg9SnvrUUGOG4HhnL9SQ9P7bmWfqwpRXNxeyFurNEBoDmNqafOOYEUI2
FIjR36nRyEH2HPidyBRbLLWAzoqlSj41nit1qDM4P11m/9Yack8D0u77OvA4jKN6
rgZsdQ/2aC/Toi+rbPpZdsoOkrEBA1st2kpoV92IvZbIdgo/Md4RgYJz5fZZKA+S
PoO1zeF9K0y+5PVkFiMenIdlUROZO5Ll7BGXG0YnSDfmo62YSd9A8HKzobwMp5mr
bLGOl2JCNT3hPd9ro6ihqN177eQ/Iwm5BVt3qkUKZU/NZcw8Hlm0HeUzncpJjjp4
4C5CgvUv97SG1XOWh9lKoadrxBgNRmhCGnw/y3sxakFVhW8kqER87QP97UUXIYkR
tpEJaMzfEKOlHN+TePl7DTeBQuqV3SbC/kuP8P8Ktma5EEL51tedrPduDvlaKMkJ
3s4NoLvRrrR1IsBp/FFR+hyZAxvSv6NkSSayT39rb+QxCyT6VOk023DygV/yZ7r5
oeCj9Lo9WW49u3EBYrfGpC1en6IRwlgieWhI0e1GghPmqfaqkudrVFkpDoBljr86
fC4QzMo08uMlRV5RKjSUS3MiyxUolJcbY+Wv9KN1zcc5k1ioufBUaAmuNVYcaNhO
39dxkgciWtU8HdKC/swTfPA0Wl5+CHvZ8JVjAeKOYnmEqThWvoNJzZtRI55mauae
+O07H3hkEg8uL/btY2rolMhg/WYMxkt0Wnh2ja2S/59Gaq++IaZIyPHcgPQuRfQO
3c7MSPDg7DNtvlAUgOiL0Ju5hdRpBF1id/3oaDMro34gBSLwytRB3WuSFtm9Czbj
H6rL8YDjHWV4CJt5eaggDERh5uJWmF00CyTKItXfeVDIMS8Si3Ap19p2NqeI+Sgb
p2IFANA3jEPiglrBJ+2W8XXBc63FvhS5SauXx0QuMAfnSisD8Ecq6nN38li+ohA3
f8cvlcUNymKPVlklA6aQgrju/vC/p81NA1rthDxbWHyJdQulJ+0SRCwQiuJYXGD5
2r6W9Wq4bfZpo9LaXB+JhPxptJXiW18cKDkcL8htvRjd1MDIoiDdknOpkQXaKbM9
RAwyWIgtbhwag8T0OCD0NWS98taeY1Lkk57qO3yhTvQ6UIwHOWeexOKvetzWsnXx
xzPSQizAvd0uJ6dus5U7vI8fAfkwMtH1TEm+B7ZB6RClvcdJn5XSh/owWXl/vYhx
jTRvk+bXXGtMP8+ltWOtLhCACVgHMxBNZDohhbDYE4nJzPpZa+9JA9v+1LQ7vpGF
edbgddqVG0gpKUQPMfInu2o0prC9zoIv42iesppahbWDIl5up3F9WYmItmAR4BY5
YJdgtdYMlWQUO8bZLT7HaJvzI5uiS9X0ZzNjpBYFB823zKxqe01BELgwhTB3FdEx
w4iFPayUndwB5vaMuXhM+CZeYzhix97J6fUjFzQvEcAMNWYGAk64k5AAk42QthcH
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Cc/M7uSQyfEoGl+Ltnc8FRWwTGYjOtaf22ei06mJOtTjCXSZ08L44nG60fOh4E/5
IMqaDAuvdDVzxh7PuYH83E7VHcJ63efhohGTfncj+COSxakTdIbYtgrAIo6BGqOV
/lD43rNxfj7++tQ59zy/slRQwe21nZtpZ9+CI4OnaBhX0tfOoMx2vqainfnpd9nu
tE8KAQXANLckhhLyc1Yzrm5i6WJeO0CmOSknT7uew6en0iFw04McoURIWyR5eelr
YvB+osGjfUpJ/YJ+wQ+udS0vaoktwNjyhDG+Soucf2Ew2HQLO8Snl7ulkQbgDXhS
TOTcTS2oRh8K70ZlpjUJ/A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2864 )
`pragma protect data_block
+bBVIY6xuuv49JIO6WjZVJf/KTGD700mNGoI0SQlL8Tr9O9mKh6tgxurOL0uMnz/
COX9o8WaAM++Nsf6OATcLe6JzJe9aKRU2leqs1827e6TsK/wXgKyTviI9Uc02nDS
Ol/9AE6k0egYjdtJeDQAZS18MiT45pxyHSDIg7DzEikenTIzzK+NP1Us/GzeaAEJ
6RjnZHmlv1KJ7Q2gchKIJLWM7/8pBL/bnGPKC27sEDrXqkckbjsGSJlBemZ1kDDQ
gOH8AmrJCDbH+fpzwuWslo9snqLo3TCYX4ny9Irm/e2nCZzkyEWzFEsxgL3w1/Np
xCoUjUOr06psLDvisRjd3HJuEnO9AN0OcLLe27B+Y5yKr8s0YqYEpl3SHPyfeGF0
KI8+FH0KLGlev+TuiaADx5iIebPNEPpF774ZWwmw1c46ZXuamXkl1jS+QtMnXfcD
PpGd45uHW1OVyYSAy+f6cTYuoRFgL89/mJOx92K1FZysozv7n7BbhE2tWIKNPwHQ
v819W/HLQbNLgYstflnYiZlxFrgoPU6j3yMkaDEd1eeLTGLvxLwUaoe/7kSejrSH
j0tlhoPp1X1oA/yE4C0C5MZovf1yM7WoOR162qTAjY/KQ8ilIxRvLq5b870EvOgt
AXy/g73XJIfc7RSt+RDK5HT2px62TTzonnm9+lmb5S6TDkm4X4ItiR2T3M0/yWsT
JeHtCg+lrZCHgz16GJu3w4pjciH6MgveSYPQS+LaoLLU2o1jfgNz6BGbNWQimVCJ
PJ3bicRpqfjTiGKvziZRkEPBrgqOEOsOliFZCLt7xGVm1mBp2tj+KyiBOmKWfAKt
ptR0uIi3S3lEa3yKbtykZXI1vHGaXvq5AvYEwe+ee/R5j2j6rC4MtdYAVXvrP6XL
YxAGe2eP6BxjUTr9XZZ578fr97qH4dv70QAOl7B1be052VFkUV0Whj390jydNGn/
DMl1/3CoRoTKQ6vca33SuAh72CJwbdLgIwyBeM6ZcEgjknO/pbs/KtdG8/f9DLTW
7z4hBZEaBaYyGPGTkJ6CkFTrcpLPRen7+jklfWgRyQl4K1lx+rpZOYcBhGdJoPE2
6FZSN2DE0L/3+fqd6QHQNpTijvhqZ9i5gHdjy3MaYDkEdLG4OjFusbqAiwWu/k5w
LKzR0Fue3Pr5jGBP4j+YMo6qE6YCcwDv+rf/NiRSMjVrek5MzlqO6Oft8Zt5/XHD
/xi8h0f/rBOxXpXUf0dKJFKeutQBfM7Tohj1msvJyUB7NZoiJxQjkslqyIRmMndA
0Js2F0nJwPh5yitqpJpl8bbGO4bhbDfgm0Y3TNA4JTbPbbkvslQUGo4ipPNBVKCn
POUq5c2QwpAgoB8WgwO/fVFwnBGwgL/ieiZ/c99LmZH3WzFzKg2gCY9M4XKYchv2
181500ZxZ3Go3iXAh1IYq88hMx4jHxHNA7zvYKaXqHCcu1JXbof/4z9MN/IqcyZ6
/Sip3TNuSOJecJ2Ux1S1D1xnLVhqBX4RBTH+gBl1GXp4EyH0ffbYzl281uRti+qi
bj1PiUXVByobJdO5GHjSAqsLUCtBvyt1NgFtKn1Fp7SW4/77/BbmhOGrmozpY1So
NGrFU2UOWGPId6VbQWd56Zo+605i1bRlZvclj8HbyCLo9lDjRwPi4BN1ygaJ3vld
Sd6STb5vp2Jc5hCCYUJUBAENktfBr/RAaW1riSH28ny6migL8bG2pmSOnv5ApfQP
vxt6yLTdseraAubRKaEqRdJ20HgcVwZHf4jWaQ5Upg5pa5WxVr7xmebd8uF6Z6M1
8FaGza6W03PDC8O7mjZ98cxvjleQKjHA38tOnSQphOUcBpJHuY4Cr4OAuil0U7DX
Qt2/WIGjtpRTR25JXPl3D2Dzgvy/hA3yjxfmTBTy/9nIyY7VxqihkSHPAWDfVz7Z
Lr9XT4WtFIaWHwqthS//gqukP+w5quLjgtA4ss9DnIrbHvkTbQI+Fl7VkNt2TU+K
gszxKxrZJIAN+isEZpnksa/ylFd0k/2RooJ4rn9rwP70PnHY0G/9ECf+Qgs94AgQ
ptY285QTnkAmyIjNY1FNMASCqPNCDUkjr3csVcD6LIs2hYuhmLCszgdZ33Zdod6C
8wuNYCJT6ApcIUHRYypOntJvSsz7amNPoCHuuT92Ga28gX64XbmfZ+J7i5vkAZH6
LaBu00iDl8PqtUZ2sHbBGy2fzyTlYwXnZO1u/txZelyVy4Awd/EJcC/PCqqlXsQ6
FZV4WDhrMBu8ffPxB5DgM6mJRWMcmO73vy5GhE/AG8SxMRu1BFngS08kM9VrAn89
lw3HkgEy5fwcF0q1EF7IOLsyUvX/6IFZt9XsK4mvaBWVvuh7CXyR9nGVa+K+ZAHs
sF6MJJH++SKTZtba7stX3d/stwKRxproM9vh9XCHHA1Jy9BwZuy+riowjakasnY+
iojdehErOAMl7C+clQu6NXZlUjUMsgCB9hAS+5hJp3FwabER00bus180zBV0z7Ki
wG+4UgmTVgxpEcfMZNzq2HuDqIjmmn+s2TWqQVBb5BB0h6i85KWFryutUhhZtxgh
OUnXofZ5YWufob8rmzX1OhUVqyNrNA6xtalWNA8xaaeB3EWvsijbvAismoslSlbT
qKngYdzqv+IQftCFUNqYSKYuM+BjlY0/Yvw1VU1V/+3Y+ENaDUzByHRmhGcCC+Sz
xF77SRfU0cfzp1cyxbrxeXQAdCBg1qelv3rSMU8wOqQGLklv0K8dCEaBaIPunFsS
n7U7dyFZeXKp5h1PiZ3e1nxh2X1Lz6E4LKzz2v8/sdjtzcN/9/ZsUwyHevP+GJt2
aMr0Vi37v8x1M7Ci1Gl641DDWXXqS0Z/MqhERw3sP8TYXNOjA94pD8arFEY8u/2z
kqq5vxPxj6sSmhLa7iCQSZh9BNsKCvd1Zo9xK5r3uk2ByWkrMQ5hT12VJgV+ssnx
RjdGHpkgZtWC0zJIi07mQBVZs/0+daJqO74TEbwdK0ARBmDcgr2jDFg/WPsQM463
xkmtHvaHzmVMv3PSLvGC+yG76p8S1DVL3y7Zkwrs9Um912htzoyjVVsUR+pgm3c+
DBANEELrxRuWbFycd07mvTZD0OJAZj4Y8+EpoSEOC0ZeCDmENK5oWKOaqONF+/Jv
QrwISWgo09s/n9lPYf0G+5PzQLEi0eR1QcdypIXC2GW08w7P8YjnsBVjvXLetXih
XZMAGM+GryqNdAgxbMRq7yZI5erM4i26U1lkdehc8UyarJd9+GV85Dv9OZ0WyUTN
2n39qZInng+39aDCDck3Tu2T2uOUtG9xuISpcjy9egVuJ9/x8jajA7NVidIWqIKL
oYuK/Afs0vZ5ExiYeKqX+9UiPzpLMBNc9g1FPN5elb/4x40j5vTrtUuAixeTRVki
s1bBQKTDOYCWHQORoH/RV1ZJHf3DD4E7M1I+hK9LrD+vpYHHIoKyyZVqgjR8CbSo
wkxYPyy3WdR6e3jK6AY2ysD09BZfZFzdkGAaFa/+qsXKNb3gqildHeK+/fDxPisT
hGOY6JzYI+T12/HRLLxFRGT0pzSr/0rMNeWs19YkHj8IR6GR6mntvCnFI60brp4F
q9VhsyCbFsRtVui3AXvyUh8rNErn7c+5IfD+mWbyu4WWx8HOBlEfzyWS0ipE21fr
I3mdiq6HdCJF5CdqIWc6n3lH0tuD8fWXvFQSRE6J3dRD2OgRletf+z8PNUTaGTRz
PWeZ9YpPXk1PAlVEOAEGRfOsnZQASm7BCNLxBAxhZh31rtyn0Oo/B/sjMw4hLUt8
a9kH9HCOyUyqKStOQ8lPwwOq8CkrFgRMeXxyltM/LOU=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
fbvE1uOjk3I3JAbSz1GmuoeaWsX8nmLeNSTFQdjt9E0mwzjh53ifZTYH5kTsY726
WoHsG1nzGJhxVZDOTe3noDlw2d6L3yrnbgmPxxnTPQuTz49i/x+BJN8fs+FLTUgc
U0Y6aFr0o5cgG2jLVGtkl4qDCTu4Ly+caE2mY9KW83WobThxkKmtG2xm62JiJQO7
boXyr/aRhbKklyiAiguqF8u6gEHmm+GxiEn/0M2iu6KBSyQC7/rDpfNKptQrKlP7
NpDbV3KgbDRChBVcB2+Lu+LnyPmRZ9nD5c5pGVdRSUEN0sT3VYt310VGLpo9mXGb
vaDbW18wL8PHtAN7LcBE9Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8704 )
`pragma protect data_block
puVSFfo1Agh5YG23aJffc35KELHwe27I6B4oPbhsVO8kDXzfHk773vOCs745M1LE
Lm9wMnAfMopPP5VIQdP9nq0np0PjTMLZt+U6MapmLLQwbuemkTf56qJFEybYeAuD
YP0rXEX8dhXtcpgNx+lXFIojy8W7T6zHPn/2blRqOketVQr+C3hat7Gkx5d1QX+9
N/i7iEPKk+j8yYmX0pRrltMwA69VD6afpUJAT+OJwOJ3FaaM7iBEdWsQNI2XZCal
o1MfTZMg0O49f4wo79Ynw0aLN2zwvEbN8tnnSMTTLygWxT6V2jED7JcBw3zn90N2
c1Xvh83/Gnc+5nE4vKciY/lSnVvPLY9cpJ/YZXjzAGX35FkHMl+mJuh3g8/Tuz/U
zoZVYM8wrpocF2AcG+fnESo/SyCrqn0ISa0dprUrDiZaTVGrMxL1ya/SOQkp2f05
uimCH4kR7X3yMgP+6bUcAVrR6cRjfWjuONSf+jskWExpioYUK0mE/KVUJTyo1pIQ
HI0m0h6iadkGbKmqJmAhWpyuf5ck0YPf0zzc9DBGJ8o0PZ1g8weX7bYSMol8UH32
t4yrADVGgqNn3USgU1+huiVJDtEvSim1ofwu4G+7DQQ4QuKvZlEcNWGkdRjXdgW5
vE34DP4SsKJm982vDXINFu6e147rujFSDng/3yf5yLXOj0SXDxXwQDA0VLhhEBnP
MUA5FkjxJEAH7oNwLHeGjx4fiWFTizXsnT+LlbJahBtIYLFn+/nnp/5Sdo/x8jb4
sh0pCdqcD2KsJNLCf4e3PFIeRI+XwbJJYgLd5W8aCaGm7+AXbqZPClVQFkeQ0I4+
OMDd71NLOyuooDx/3s4OqqUXfmCUjLvimCnS/F5sqrCMUDSeSL+4t9vMZt4XbNeO
GiZQ/Sbft2aCC+0hIE+15O3ACUd0pHpaqw3D9LXig6CcPDfsuwykbXfJlX4amGV2
R+U+mTkTAPuSHB7cR49SlH39wEDMXDl+4vvEzEMD1XSdR13XZZiRsYGyV7oMCPwB
iMNHCDALfXm7k1eb/gIrmoAL0LNHM48sRszoWtGTWd22ZCfZgsi9P5cDNnCOv9DT
ZPZ6I+slCYtORoqq4Xu8MZYrjBNDVFOWnoEi5Y5ZcIW8TysDp9wat+Y1yYzX6OL9
um72yLXqrM+zi9kRmKbo2xySnlP8SS3BppupSns58oAl2y1Zr+JoFBMenKSZS5fs
fl9pnPV0KaSxDZERCtAqakwyo00fCu5hRmu8nGGzyaXEmPdXNUeLQHUhKOh4Siv7
fAynn81SAOsBbqrRLLFxj6rB8UmB8XaB+Hbc+woaybo6rRYkNY8gvKBffmseIOBt
BPd0GJAoCUy5clPD6ryxQuxbyOJQNse6gAw+d0apKtQMEqRjUcv1oSEvSjSQIuLN
BlT5ZMxMoQRpDaDGmYUCxEHUjecvqCQcSuYEYZiv95P3PIA+7jcHE5Fp0YeWjtmg
P1irL0ZS7sb8lunGNJRb1T0c7EHmRRsjsLIlDmeTYzo1lyewILzDG4Cw/u8O6lSk
AjaNbF6MNwtc0NO5VFjCLtoPo4rmpHjjYwOkcGjnWsbI67WBqd43mUgdicKYcv3w
Er3oWNePdUYkWpiJG5lA9crbXVe5f87dADxfFZ4yb/E+kFUds7+8WjOFDbeM5x8S
w/B/38U4e0qNkHtTDIqp8LuFDldlpRGI5uzPeLfNRWoD2w56NYmsfz0587sQEYDQ
g1NZkn1W0/E5snJjCpvbuzqs+sihC0FY8tjA+9Mtd54w1SrPJz13WrxYEA6PugFQ
kjk5AhvL9tz/QPXl+p+sVo9ae6B0/spfeFJwt29rmo0XuRj5Eswapw6LYHTrwwZD
RuX3wDZ1UESpBYmbfUQgPCx9r/G8y+AT6uB9z0kTP2/jMMjxmYNSqieCis82HzTE
xAkvHAZF2pnhuv1gf+aK+f+n9YLi8/pQZ6ji1CRBuRNlQALg1mgjdcY2S4KNqJ9m
tAdCEVFulfggC1uzHGVGRnFP+wE1D9pyxecHLCbkx2efkTej2tj4O58Q+F3/pHZB
9K4/giyrCsvdYEPDBI8G6h2JFuTp8FlVoqnWXQXKiQ1lJEwgnPGLujIB0PPDBAnc
lDidTa0sO1UTpcDsN8kJyIhp/HXsqPxFufRYT/D81FH8Yc7flHxh9joPc1CydWP/
JwhDuRL0HPlQbo8p56Zplj8WqMu5l03X6JAoez1+JLz30Al0qAPTIW4gW9VxARtZ
y3k6bBrYAXb5EH5/ESgbu05zDIGAZb8Ca1JCsPFUAEhokIEaEkaBLn8oh5yC6hF3
puvcfH5KpY/zs4AhjKRNeK5Hl03mKX7sdSAZkf74F1AZZq8i99RSHtu0Nb25E4mL
0SJlONPPFIQC5Yc4/ULY4gpeNd843ooNN7OjJz7KdpqWtcwZrGiJVgl5cbW54ygd
5c8PqE48W4EeeQpLAVqOchmp5fCQ0elreq1k6yFbxRhddArCs5CMPXz9NgPRDfLq
/1gzPHW2uiz0PwdXKd5TQQ5p7Rq/KSwusGVremLcIoNXuG/6Fsg4IVsCmyZV2ZBt
MVaY6rajTRtfGjgJMi0r6A/4TDwEq+y98eslKi3tt7JyB3TDbTQMQpJhtksKymn7
dyBq4QnJJkCD4+Qs8umIwq39fjfh0hHiFlCICU8MiSo+orSipnYvINlW+W7jYDcY
BlSvgkLILA3yzxhHN787G0BkpX+FjnYMmgYhu//ZqAbemlyywN9Fa21nbfXg49bV
IOxS3v/iN8yllbUbsNpzK6AkudOTeIqFji3E7rXjELFmsir418yRjkC2bIQ2uk9g
CL1kRGPhrmlekpXwWYF7z9OQQxO6kLSvSpRIRx36aO/aC3NJiRTCkpwPol+JxiwU
pMXehhXyJ6UHVrwZne/5/q0O7/ptASawybrocjMjmnZWdDQInnWb10X2GRoe8fQ2
cpPPG2DV9Vr3vcM1c7UOsCjXRmyHfbhu9CLKnng1QPFAjZabeoFQVrICRg2ZQgAH
rLf4n+rVukJukDw4ue0Yg9NKjTSeyLIH1cXDi02yXl9Rt5vAI9tqVuUUKgEcpSE0
MaFsLawx6Ewj9+L2CID8VoQVpnPURAW3j94e0Psdwv26in3ZWV/xkxBtNsrbv7OB
KK04xzGrLOIfHYLpCCklFDG0ARjS5ozC9LxhqX2CWBc5jAfAl1TDnVq1eD8PaSy0
XXXuBRNx4by+sUMw/7l5Bg1uNRy0tOg/mKskNB0mVrymtZBPAVbYUPZQxvqt3BB4
jNa90qNIYRt1+u1xSkpegoC4MrPdGS2nYYTDbUGTsj/EvsM+LYyKsqfl0mSinhqi
lqbEQHHwYCir0umflYIV99nxm/OZfKGcNvjT/GsG2tTIwpl+NKiIa7Z+jrcNn85F
MQdfj2+iuT21ZyM/LHNq3RvmuBqAgZSS6FzM1rgX+I2yuzVcfsSxBB/GFiB9y2+p
R8zlRl8cLgOW7Z6gW6RKNFotv5UDA4sKBbV2FVmCpredczs0CfsbGCZA/O4thmop
YFSTRSyfem+cdLP+AB5kC9m1sYYEmmxKGPchDeNUTSngA7SSd2uqu3odoX7fnhMn
0gvIkwe6DY1bFHY8SifieXF+mVLhY1doI85GfDHOtkrB1MGbfQDl1TlcT0Y4LXUK
X/Xtv7viNLYwhXTseGPc6+Zbq7n8IIA1JApaoZIQSNF8iFItEOM3eJyQWKPYggU4
3AtDbTDksqqHVeksrBMdxZZMl1q0LRDBUdlD5HF5NK85YPlLEJzmVWgVVDTfp2y2
qPbsczF3rsr58DgAJNN1qDk16XkYjdvEtHEiIwvyy5mBwB0V60Ej7doy1TN+PcTa
/6/O/8CXeSMOOLeBRi8y1/Bs9E4rhG+u1tcNYLqxYn6smmt2rJZ1iIVwUIJgP/AG
lWEYGxq3BiWNYU8doA04KLIoChO+Hs7LCMasNxQpbdZPx/8LP/Wrvunrq18wCgkW
RhCBU+Dy6K7tsiuzBcnyi4e7C3Bpicl216htvBlS0NKv4RNeO4xAzq49ARO0hr12
xt7WDontWQf/2zGk7z8qELvsRhzX7svjbzLJQ3YLxYvhRpXiVxRyrsu/37iCbdXJ
6AbKeKkomaLYEAUJIXCezqZtzUdzffFk8r/yYSQidMv5vMYBavtNpdauyxVF96Kj
4h0+n16In0Ekiqiva1uoYSw0GIpGLw2kT2Y76zojQl04yFKiXOeWDzr1vyi5AC6P
h9rCBUSnEqCLmRWFRjS1NbWNrItsZwyccwE5ywPqugCATFumj4iium5QtcasarYM
LUfY+xlPP3xSthooaTgwrdZWyaTqxEvoFLy9QghHx2rkTVkaa2Dx/u1odQBqDEIB
B36tOFDa2NiPkNyRjigDfi74w1ZpTMaITFfEgSMzt88vGedSxqHRBXV8flu1JqxA
abiTCNjvHRr3IGAYWiRWu7Qh4P0h0xMrxdftkN+AGrZhXUKjisLwCjvufLrORVwX
G4ZYGgNIREe69r/V7OEJLkXNdn003L48r5skDILjaermXDGHWB+aEnmg5Uizu5Fa
DtHF/NgpLCdU++WEIqKM+X2Cr5iUhJIy99SwnLHd1I3b677KMSuA/yw+QcbCi6Lv
318Zf3jTmJJiJOTj0xWxkluo7TP4FKhKGadwjnB7y81J+848L2t9XXZ28GKHjnWw
EXxSzgrHVQMiVvszPZuawOADkBRjIbEynjCH7VmOUxwn70m1Ehf7+/LBuGK1GzBx
+mNgSM1lyxvbQbY04BH0e2r2Oq2nfUzsmOq0Vx//9DOU7dXAFOMTLLRybZSvzcyA
LA4L5AbaeIT0Up0L9iw0vugDxy9ftw2cqE9t0aOcWbnmEqMwupXPT3uLS/CHc9aw
mQgs3fzcDj/7mD4JMkDKjhPRgMinYWQyMkaHo6+NvBub4Kuveyxo/eHquSZETepp
sPTFB2g5HiW9r3K9LQjca2bZrhiFb/FNXhKvr6+ogYUUoo425MtD3ljZK6IBiecf
8jcMW9XLUQICiLePuYTbVH92wX89WkORW0o32FD2aReP7mulznAJdJ2PX/YGx0yH
l3qVqG8jcHXeAcby5kZaQGd8h56vNt7qMfUu32QYU01YnCBjY9dE2zkVTPOROFWK
fyTesmg3/s/i7UVuA6erIgjYipCuGj1TA7BjuI3lIK/k20rBxn0sENxNd8Lme0x4
PpiigL40cdd3APpZ2ZxXf6TtJKllBtWv0d+PYHLOy1qiTc867s/NmFIydUgZ8y0v
2kWfZdLuPH6Dfv1xNP2VOX/G3qZK2EQ5X2lacVb8NhLPjDks+YBX2mU0A8l5LKz4
l2qDoYpuqpVPN2W1Q9Rtuu2RcdRn6QB1WNgLwOUZHY+P+vmJPA9PqRwr/olqy2Yi
1gpJNPPZDLshB39MbqCdaaWuNvvZ1FEOe+/b2WjwaILgRzs/vWogfi5854JjysSQ
UyS1cJ8x5BTQfHJFB8sllGCbnQ2W3HmypGdVmG413bQ4GVCo1NCMq0y/4DVacAi5
+qE9RK1NirpnX3E3Uinq4FnStbWVzx6GEM+gSD0VVUz0PVzO1JpLNzdXa2ENumRm
KT4+t/HeGdogtqttOlibpmRp14UKc8EqqGvHWyzNU7k0TeTAN7JYnADypM2H4PCF
kYB6uADBtgV0Y79xDkL7MoGi6Ecv97VJylbnz0PJncc9lC2RbUytv+xliXMBjAdD
2maT2I0JJvTiUEdCReCVBli0FPKeNq00u+hxFYscLm4wdEQJoO6lhQNdSwfEYr6h
xIM0SeP33Zb4rbS55BtK76fCi3jK27fXjzMittXJYcqgMkioIGcXrwCqMX6ceRxf
5H45SkCLHqZCtZP/pObfU38ftYapk4nKN1GTDJ4tzR/U1pMJ1g470KRtt19alSgi
NgjQ56mfhY1XxN8LeJasy85+t8qchlEK+/QOUzenwd/qF0GhL/NcVBnXn/cKcxJx
oZ3iOQur2ea46Dc66PNqqZ6B6lQbtOuZGG+mt6A2cYuZIdyWlBF8Tvgnv787co4T
RJ9HJVhPmlw4yNHPh0xeG7nSPs5bNbZXJxD3+T0NZh4gEqIZhtjZz4AEIn3tbjM/
BsfB+4QNuQH5MvM5mhb3VldywrIekQZmINtS1SokkCwtG1QRO4uPFt8jwVkU9mN7
yWNOO5l+qTZs48DWYGnRQQIXb2jZxCVS/xPaZPUUiw8MBA83f6hUKLGmI3wQLG+h
ikBFtbL2iFCsTtwBj5z+ZmkFi04oZ4ZeI5ucTjmGaXBQInIVggfoNuY1r2QaAYeg
5r/1wutdxqd/0qMxYD+xd7fzAZPs0ATKe5R+cAQXqEgmTOxOSFIOuvhyt9vARYZ8
wAo/ZuKIkXNUsKaVR0StJChEwAC+e3MuKMkj+ruHPhKEMLucLQIBW6TuQw8aA4RJ
qpG6dwAHNu9Pxgbh/fqBdcef/n/zJ66gh8H4Xl6z+M4mh8GbUNrE1+fZ2sk1g7rR
nytNIs0/4FrjOWFpELvedzDj3sfvSrO4Lx9R/UhqdybtBRsQ2p19uuBO8rDUXxbs
rvKwYzyT0bBsLHDyNncCC5BCT5NS4PRx8DCw9Sld+1nPhH8XBZHhz1sTZs/qFlxJ
15UigxQ1Ys8aWvLutwckwDQphZYHxWeygNYsnrXgRvvB1ObeF7McjGrpwwMRwfkw
cfyFiEgi1+1cddhB/9M88qIM+G1FkOVje0UcRImgZnT4qbxbEcb8qnCWXXckZtGD
xl9Q0Txf72a40PorpYPW0wcHVxjbVyZg1eliBdiLFddDlw9QneeeyF8MZCKLupdL
3IJQzUAeWkLSNoeSfPnjuHb49VXSmz6JDWTLlJHyJ3L0pmMk+Fnp7zKnzu19aTWV
7i7xvWBzmtmxxfMYdRJqMhpJrGd14XCXYYfAjYTucSyexW/GsIom1nKRjChA8Uw4
+KDLGrd+vRdMbgn130yuo4XKNF9u+odGiIh6sC5ZzFMiXkKJ5UnFbeMskaHFKUR4
deI/hGjChoId7kVy2E+iEM0Uj/FfttjzRR9eYQF5dOaEJC16O9BRQV36d3ygwZNN
CJmMt5o4TxqbVPcOTMLA1TqLSJScm7K1kjSUNh+7KS+ecxOJmsEcKPxNHXGbGwlN
NS2mPu57ZDdtkhlTCBhxrGNXJaFNznrjUlMBpwPpsPJaXt/1ApwrNoieFeo8Tek7
T1woPLAaBb7THQcGTT6K3khJzsAjSrXQ3hyoFSPMx8VKt0Vwx/P3Ruo5NpZQ07Kz
zDeKdKSKxEpbubjU3vsYDRblfw+Yk95ok1HXtZ4v0ha2B2Lg8kChoryGtQyz4iML
Ii50BDRU1hJRSAfKgLlVkp8AU4/N6+1HXAwPiLAVXUr4Nn9C9aOH3UXShnqvoG5m
BwuPwAIOZztFgIR6KsoMs8C6Cpt8DtyUSkG1t8HUujfPI2EaCD66nx4h8Ktu93yd
0m/oJrj9Yl43saOWVFRlPej2MFaFE+ifQUSJADNE1jZ4tFkoC5Dhsctc7gi58njr
uqM/7SiKOtdORYGdigZNeS78XpBIIbeTrC3kqBm+C0RYf41cCIUYsmpqyDB+QKv4
otHzf33XkILRWEjLdktWdLNOby8SF96WGhusRRZ0R8EzB80Dj/w1bSwoFb/yZ/gl
4Sv/WRanb+JS+nXSndQ+h7C275AgEamRoocZ1wIOZ+zDfP3RQOgkvJTQ8dNlatbP
KETl82drNfxP4XhgSyeMPIIMgDZADNuLmrrprhNn1UlQUcPSvtDRDzgLWMG/hQ4a
yLapE2v/xDMDqEFu0i3LwVfSw7rUEcI6JM5PM+Pz4Jbl+F3+G7goPyWxgHTrMhyR
MFkIB0sBiy3n+cBLIoNGQ70spUBZCFKAZR8uqPSpshvrPCxNwLiWwylk3VHK6xa9
tdsRiC0J3X6COrZrDsAy6vsDCvzt3fV46QmAnjZsMclCvxiySyTDlpjnAP4blnyB
R1oyGrGjAwl8gqlgQ+UMujuL/MTRDvWlSNfm9Sq1IvTKQU7tXhZtpS2P+kvVilqd
CWEuaBgS0y5qmZ52z5a9Na09rpQ1Q6SFDliXAcfnBUDSgVOgs2MSccduNIH8U4jO
rKkKDaSNNwJQcSHv1ZCL+BIrkvL0fcUpNRhzQgoPYkJWCxgWlngKjsM5ptSXsgSn
JecSzi1h3JgB3f/4uueDJp8c7eUKKHPJktg+w8FGolBTgDXVyNmi5JtT2ksZMRGW
fBodyYpWvcrx2QC0qa8Oq8k6K3pwUE37EDNn3UEzoPGpzdPn0kS1yZdAivXHcL6W
U/l2QbgtBPrIgVLJGtO5/r07kMaaNeprjG288d/Ipuqr1eAxNOsrgmSeJ0dhgxQl
+sG0FsznzcEypDHP5+MAoOpiHS2HCazU6mp5UNxU0w6w3EcVGlsrn1EZtY5AwRYN
0TqToXFHdtR4Axfey6w2tfeegsQTFlYFYAeWtbii6IfTCwCWvGMKFwYCiui7+lUZ
dfl0bZPNGQ5xpZ3l0WXCNJarBaMu/6WRgzzFhjWxlj2fmgtWA0tdwvIaeJt6rRdr
Mo9H1uzXAyom2toDiSkBqXJOHle8ZoZaVVseJl3FApUhIO/jWR/sooNW43RHym2R
TEhyj/QfqtTFUc1BcEaYu2DRWIU2/tA3aOg46e34oDcIyQQP7Mx7tu2mo5dAtjIr
ZNukuYGFi7aBEJRQynPHwDz2MCLhCnIb+O4FZVAdfW00XWCLhINw6fZPQ6FNYMR5
bjWYIk4RxCq884fIfvGnuzM1Ilb7BnH7tuFCjIldIvgy9R0O6k7aYM6b6Bq5xlNK
06LGaueBk+3LSB1nGpscLmokNTeGY8D6KB4Sd7Fb7Fy9MU8Q1zt6rif0OMGNud2J
ArqnmbE25sIvW6/bSZ7QYdjLfSFqZydTfIUPfQ8n3VNtxNv6Rllt8b0HgqMC+HO2
SpM7hOg5lAfgzQ27PWZCCl33FSuRcDdCp5n5eRUdHNk9Wo+1yfkcZ15MbCw3bu7x
RpdKWtBq/BFXjZiznNzDWeKnZ76DUY3QQr6cW7Nnu/zb85qWCJQaGIjar0VRkNX3
Iq6NYXQoCggrvPMs4NcoTOl5hrCEDdx6lB0yfmfcopVg79xMhLEXjOuFaXZ4pHC1
25qW0n/FMwHOJ4R3Yuv++tjJ7bQkNPzEZygO7SLz3h/vgiE+6lai8PaTsjZizIU0
Y/8qqKBeZUthKWyjVlMDQpy8mxE6ZtILpPIXYvRxk7S6BPkgb1DLwzRbEkd/YAfv
uwnn17JeT6iIQQyv8mUZh3mvm3DqOMY2NKfYcwechA872u8ZxmkTboNtlQTKPvth
ThBFhX+lvaL9iop2z7r98WCc3yxnMscEhZmsA2cBCqkbf2SKis8gGX2eIN5Jwo73
27fwO0qBIQDI5o8gkTdVjODL+8x50Vc3FecGD4vA/YdCUV0qyNoh+haErcbUNKrX
TQeoC3/HTf8anyixP2r+g0x3Mx/5RT2f1kkDera5WHYbyx/J76w2MouFe8rY76Oz
MlnTvRRjF1oWHIKB3KkU0i3n88UYQ3M4JlZJcOOexlD0Ue4z5eWJrEPEp3ctEKBS
QYDDh8MKwGNwN4lNlPEl7v+SCKJ54Pr5UOBFSdBrV095n2Sk47tWOx4i3zAZwaAV
ZHHTRttp+FABdDCnJwVLtq+rTTLRCcCdC5y7nxri6ibB3l8Ea48MLRgsQX2P6FAd
YuINkxPspKgBUgotXyEBx3V8bbOFStjgVNkyeFBSb7/QSQN0tLtZXqK5qjCveOcU
Kx8Ip7mvDfoK6cked7b44hjdYi/xFy9w+TrRxWKLzAKHKS3WqSLYYlb+j7ocv5Wb
P2NH9TJ9brqqRZ9utFKyh1wJMZFv0ImJMv+PV3c2BTILn7dPq8lCt17SvRj5f//o
zQSFMtBy7Dt6b9AWH8i4PFZY8irYrsQgvHczwJVOyipSii3wcGRK+Snb3zlpLOmW
L0rlc+mgnZJtSeyEJWalBhSxcCB0u8X9wI6T3u1afxnSYBgKMbbawbiVmL4zrrv+
tDcLR1fN6pkAoATa4t+2DMmrXbS7v62FxhJPIAN4fZfi4LaodaNu2/UAyy/lxdcA
orRVbGQR4QQJtaG8Wg458MdShdiPE3HnJxFo9XdPVCVU6FEfFM2uWeCg2/7nfF6e
uU7C+qxBfLAGwJyDrJ8kDgSMtoqE8ttlfllk/8EsUIavEcH35J9vAEjboLwzoMpl
+DejINGVoXQQVHhOyVQqVu1DOJaNh3CE73slRgle51SaAZx52qb+rxABigsITJvr
9i6QS5ahGK4lJZ5fqxPbPjXXVP4ty20SdAPqQis87re2dFrAp9MXJDQDqXeWEPW0
Urnn1nWW+Q+5o7bVv99U+dq4g8HJAMzqOfzFprNik1MItPKb1xZAhM0mF4nabgBg
QTnqOsBMaM2S9NDlqiRHqOy73rpUO/MxcDZbOmMEZTVBHhQXbzwZohS6cNOGXHDe
2AHL8DliFJOvG43f3ddpiIhklIhpmHa0v1u/kiaa1rHUO1mHKFGMP2zZAnYsqAlP
J/ZFWWfrsP1LDQA0F5hmbUrHG5HI29pmQPhprKYJlpi9Zzkg+Ili3Y7svmHOIxY7
+1aRK6KmpXPf9/WgDJWRMAsOobED56XoNF4sqXpJ7NmbPH0wSnjkHOFveenEk33Z
JbzIJRtimIkPHxnSnt2tFp31a9HycbilB18nNrAwYQau9Nk9cbI4TboIqLXRv4Uk
595qH/ulO/t5bq10pNGOkBKwGcKaoISeNYc7TR8JI1jWES7gzV5WMcQ9T1B3WS8U
KU8Ct7NLIKvu9xhOljU6V4wA9ixn+GTVH7bwvv1UF/NvayT59VckLvZOsGMYPfIX
tdj4drOQX/WJBaoaRonOvQKjpIB5PmEvs4t19NTwgFtyAwkvVOLKnEXmDxH6Qsgm
DhNUZnzLTcIfRF8KrmN7th3EzWsNvLLAhrtIvbsBQ8lblzuRcHcZ0UoblJkah59k
cOj5twHuYIIOoOi4YNhcLB0+rq63KWw06yhIlSYxnMisaNakhcm9HvvjXwgOaQSZ
x8GFozxQ9SDyK5vCEA0E8r0WAls7lLFPCFL1Ix6D8kd3vljB23wUXVsJtS7wAmPa
IVIr+kpPXpEBYlGE9+j9m1ncAZRr+WAdjbQY+nW3SW/HeQTjp2PYRmTVtO2G3U+S
UjSSXb6WePEgXWjd99/IZeWe2ANAWoTV83XMl8wrx1lvjE3JmTyQzzpLRSCB0hrv
uwaCQNwj4ghDEGhxEmXHJSCDyD/Olcgr3haZkiNNmBWujyupXKZRJqli1nsgsSd6
jso2i73jv6NGbM9ICnS4Ist07j+RWQLSPHaV52Q3rEbf/etYYkDcP9LxbvZNUqL0
J2vYr/tWY4oXVLl4pLeBg9LASly6JMGLFplsr8vPy2i0IdUVs/vL2Cbvdzvb6Zb1
BmUo8JKIW3A/3KwxuFvoUwUFfvSfNPdW8bFaJx4QdQj5YVeEGi5WMgPNw67eEoRz
08vMVyy22UXSB6EeC7prc2h5+0utdPSEaNVhVa6L+ixNaoK4zHJG/QGtHekR+pQI
TfPW+rHJ1V/ggrT8OeUcLwC5FuDlax3QPQh2xfKfmW/oILuKCcx333LqWCAUFhEp
XWrUbPGUpetkT/W2PCeVug==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
QUyYEn3EQu6K9XqEtQRO0CSQBVC+TBQy/eH8V9AOtyuWZVT4xaiRfxSc9xf/S/T2
2H+SxZo6K/zXBpu5SvPCHZAtKKBVZ68loE8xkpeoI2Ntojyq1dowKb9dk81rtwly
n/GKxakIUkWWZXvKjF4PswU96Xh5KIFBNO2lG4HLiKL5JSMhKTEX9Df7Pg6lqigG
0zSTc+4KTEtW/fycXpnyKERN1oOSVg2j7zIAm3SCym41x1rogUtPp5RWrVMun10l
/xE7j/6hpT4wbxDxKaGzOJFsOMNuXDSAlhTwOk7x2f6Z6GqVfzDBHV0XW+6uPB+Q
mfQv7rHGV7jBRsqKtW0XDA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8400 )
`pragma protect data_block
JrXtr5RLd3Lz2s8lxcNqUQVlAje7xfmWjFR2swsnnu/yOgDKmjiahW5of/7VWa30
oN1Wsv8+azfvzgjjvBf1h3TQ+xH7372maNTxCcEgr6G0MGjqiJFh5CsQ6U8PWZm2
LkAerDqoF+IrjzGjzeSG6IJ/mU1Ua5qIZm68yd+aOw5hrOjjOdVeADmOnbTu+pqH
Sp71WGjwi/FEjsgRqfNh9j0kjNTPqDqWyFDPU7WTYHi/a9C0xEfNEjHfxvX80DGF
lj8vuHtyzejvqCKbSjQI2mJ/Uo2tDf5etk0BFhLj5sOQnreHav46zGvWELCQtRgj
aP/tTHqxjKNH6iYE4gFaFEwLtJN2ilYEuVmBEVfWNv62im1khE9151heLVkfYxUn
ESpkwcgBiwX/I57biYY87F3kEQ3q0t4Y2754DNxiJ1HhZIybbDYKVj+9WIbdAZXM
JY51gm7mIaDy5FuMOyCmDctgdhNMux+FlFqaIryN6V9vlsIFfFvn1RbIBT0OOJdJ
IYMKPG3lpxzbwKdAP/rB5hQybWQZTNyFkcOGEuDhyJ8O2ov2SYYsmGIVJFLKzGyI
Ttwm6To3jr9MU8113AsUIZS7WQO9FUgUl3QLEL07XV/LO3rWnJbGlBdMZ4ZwxBlY
bOuCvHiXCnxFc7oUTqnuEFjoszUdephC/uyUb7CB+AL6L1LQIWBJI6qVFV83tyHp
BQ7VHgvvroYpzSHEB0kOgi7nsBfPUQSxAH8hMo4r/Mq8z/Em/VoGtVHk6ESn3/I2
OdMS42TPhpwwNJS3may5wvnaPrnKzjDlPOgf3LnevYDDq+2R2GLJ1RRfpbg8+3q5
zhcCrfoWCMNaU5Bly8sVEqcxfilWkeFr2a84Y4HyUPdW6954FpHKDydW2BtZZ307
4p9QUV5EWsFb0rb48fi9FT59Iq1PicYLrVzQ7CGIrvmqzj1Sec55qObudWinQq3b
9D56QuPHFzwdo+754qqaz3ac9rLzLoWQsnmbXatkbhHzR35hXDRtV7+XM5n2ZqNN
dm2LTIZWu1FSgxjbwfb4cixK5bjVNBkpiemowKLWkk9yjTR43JwUVV/VnCctoXHR
EqYrg/plpOujDKvs5+u44bq4yHTaNZ9VCt9Sysq9TSa/GK+MGIglobmt30k5q38M
60LnZjszS7GWHd1tb2xebnPtMaOxaf38Q8H+fDBAmmFNrbMBI0FJ3UdK9WdAgIWW
ij3A71hqnMHifIRJzVlq161uwXZ1w58fOszyI7luA77RIAANIroCRvE1VJHlGWWb
wX1dlWzc/x+lWJy2Kiemk834Ee6tV/fCqRKcEFEjtgMRqC79yP/AbAUhyN9HPT13
LcHKuLJBY1JcZt0lEZE6EwK6qe4XGJFkUcpxOKk6npKOAsl3n/K1bVawR1dPUMZu
o5iNYFoW4mI03mRmsh/sTcuCDUvqn7oKEjDDLhpayUHEniFKQuLD68byrxVcE0LJ
Y5FTXo99Fp6hwRGq2NC/7EPD9GEA2431KXk4lcICfItdCxijaz033P6XBctFIUQW
XYSFtBGLybeM1S2JFDMleVBIVj6S8IAS8Mz4+MdSjf2h6129hzb5vT9knrs0toC7
OPO2uxx/12ulqii0f5FTsgRNO8iPjrczv/FyvG/OmGOAlQAal7ypOCgOjo/SRROZ
MGPUl3GkenrzDo0GGBvNB3hWYQzjTVB3DogHo5i8ej457gyP8/nCliI46Jjt6CfQ
5EcKJl0VDbDox8kYH/i6aFvfO14P9kYTUR3nkLf3G2fLn3oLnuJRympOh2VSejiw
q4Hww5/RYbzcguCRWaaEIzFTJMf8IEyL6+1DZwfVPcvhhd9vx7fGlMc2Iysp8f9o
KrXexu8jcuNf3BLX7+diWRcWBM3p1oE64/0tZFkTSzb7I13WTm6nqytGUGFUMcAu
FYlcBbgy2MpFFx2I3ZbJVP58YcVNqclfNnSvvxQDsh+rqlUUZIRVIhq2RIVIu81C
w5bAvPwFB4/q6smBhehrtSuOfMUZXegzusVhWiYqM9DUtsUGiZ69jC3Njp3O38sj
O+3Oo2E1cfQabVTB2Pk/aR99ht398T1J4jD3lmdNKh0lPATNjscoHpzCNmwsjpEJ
MPIZSuwLrDngxFXMN0UUC+UEH95wiA5BK5cL+P0fS7U9MrBdhbnWpvFQ342ROO3d
PzSnh5HMlt6FsNLzvRS4DpVdPSedgGyAQ6xjUnKH/J/cdHw0aguwv/AEnyjwb7Bw
2tH589BOnUU4fzANEgYaijsnbXtOKIAwqY1SOxF4dLF6csQJFm1e5O63p23OToFT
hEC96PzcJr4/tJL0xQ6iVIneb8ZPh4OePeuQIbCZ4E9Ynatdjr6kfstntztu+IjV
Vpft4BJHOfnnQBuHXpmhqQVvgcg0ym+Nfx3goIT/zg5b/YusziVFt4YcE/z0kZN2
xYB3iFiUOxZyieN5aERsxlX2wWhTT3ehL5tFFwi8LqK2zMPs2SM+V+zWtzNZkJXt
dP+Md+e7ZkwD9EuOl5vjqNC8X06RwQA/ZESJ7Iv79Pi5ARv5MCsy8umWjjRbc3Ge
kelzjDWByPBh6FhEWuH/lhLBXAELAhsrJEpwMPMn3VeGaOytY3E30BUWg5cE0sqZ
NevlW4rTcr+3DzeOav4KK5SlZpxsX3rc7EAVM3QWyDg3F2WBc+kRlYM5TUrBE+sj
Qys5Te+Hzz/H0LJmBScMZh3kV2Ok9XI+vFnJtv8JBdmohY3GltZ/Htt9Jv9rMCr2
EDOGCG6Bs4lMsACrdQB0rxPXzNmv//dQPeOx8x64zayZIep7H57i7cdEkJcvjNBN
edVVBBXoCpcf1oyJlV8s9OparsCEv/+4bRoCwukuOaOdwPNJIjEUkyNKxFE8j7O4
NZyxeBNisu728MN/w5auoJlZriWBEK6AmJHMiGMltJ6RZZARlgdBfUj9RT4dU8Go
lKqtaP8fMC6bhBkucFdsYZaP8M07ygIqg29uE7a6Bm+TZKl5VnuphYtKSMCvXEma
kjsQJrqIPdjYE41Y/T8TZ3AM/Cav+iAKFQyGarDV8aKzwgtpEVKddmE0md3mjjNB
mXq5kDqLDxOYNl7YoyaTff8fe2lsTW0q3o/dxQIxJkOiOgixbkNyqWmjZQ54UfxO
uUfRy/wjUZCEKiH9qxlG2YAkAwiw7dPoqt4ZUQQjcmpptAj55GI5BEGYKPlDTd7w
2nVUZq76IOq/2aiKsd6wcJaUcKFeaMmztU/9mLcl/dt906PJPdLUY1b08yPs5YG5
KLZ4Ddv5DNkEsdSOuQf/nW4pPYBMXSg6uocVnPsAfvr2yaM+DgFCnH0nce0dZcPe
PrJebWYYVGuOkURvGNi5ZK8feKod+rOE/IhmuZ2vfCrlJWCNME7PR7ROFU3vrIJK
MJXhV76MRIP9S58CM7VgutvMDEHC1UpVH18g8UvaPVN+5Bdxnl3skwz08rbWtjbR
ZuXtYK90wfvDSZY86BX67oHWkpkMkN33MnZ1jeHbhpSDFWOngvSVjT+UV9nsT3Ye
b2R++gXPM2ten5YG4k6ZVCCbqpPe8Z2KpKf1lX1inBUwQWYWGZxJjqfsddaqMjWP
dvJkxAZmAi1fLLYXElpQBWIOk6EiuZEyFZhKwrvYg10cjh2qxvpAzXJfA4/vfLV6
B07DLZb3wMSVrTrDJEIV9Vp8J4O78S0G6f+TKckhYHWXMwh8wHdymFjVq0pHZW9O
NVxYf/EjEMA/C1xdmZHm6zRo3Q/cDnoG+6MVblyEN3uraJf08pCrKW94aKGK9wHv
W3f7eU1D+wn+1zmzeb4swh3dqOrA9zHyyW4p3PJiWUVCq1shipCtsh6FjgfJub0G
8JbGYu4JrBafeyQbhPrfmt6JA1UvunfS5uya/MAL+yaqsvrHsT7BKIN0GP9TVv9F
p5k3Q3k9QzCMoAUvnddmplUYpDjQVe8xqp2JTlCgo0uDiGp1zfmcA4hnvxT4xaQo
oR6EjTjtoopI5eCEmCA6MYmuJOy4A7bLmFIf0CgZhoSlmRPPGeIWJiLlXdbt6MHv
EEgxaCu/KNMGmiluiMAI0HIvn5aVT3jK4FQKie5Uhypug1MeeP0jWfHpJ/kV9RDU
aPZ1uX9q2fBRDKUAz3dp73qIqHj/DX16kKdZf4ImPvtQ3BX6yI5QcVXHuYM2HQM5
7UOpnT2kiGVsWfs8eGuDaZ3cOslgrzvdjzUpGRSLcn0vWCqfrIWGyB+iBp7egPV8
eBWAzj9e4/LXyTqrL9OZrf26YUrEzsFT3AKoAaWLnn1B6TRoon/Li3qhdjGF64HL
MzS1r0ysC08OQTRTc/v50zsgk4TVSG0BEQ0hiS0MAA53Y1Yqxr08udpScrbsK/Ei
+4zajP8xgvr4QzpYsmprF8pOs7SGF++++1SWAp21xSbIYC3eFqXYdLvVbOJBtZ20
8E9vaZQ0ZaxJtlwMoMEROSB3W15Ror2trLWyBPvyRZu3ig9pXcU87sphlT6eeCTd
0AISbaGs7WNTEOBloP+RAJasBirfXEDnQ9oEllpkxMqywyUxqgq7+A7l83RRkPcD
31YEcJGsw8d6Z3vlPrLIPJ/nYCDzlzfRJVjSLWxm0J4mBd+6BkWfEk0/QyUH49zb
rJ2KK/ywU72isvKOOzx2qaY+zO+Wp98rCSnNe0sQQongp5m6aVDos+gJ0+BJbloG
0Cp0b0wA48XPl0cMWsx+XLMQ1s/xLKshlG1fBoBA1Nw/bF2DWxtY8F9Uct3l9xTw
vb569AimhZPvx0o2Ps7YKKM9tBWbKsXOgEc+6Ezo3flDdM64LasS/IDtoKORNS8x
SSVrvK6b/OlJ7AM10MlDEEHoV6sno+8sr1+nDYnhLsXX+jTZByrIGhwkxpBgGGZU
mq0uzMwe4mOXIWyxjQzjsl2YK54qzzFJFOS2xxx5/AwuSndTJ5eadnl/xyoWQnUG
nqUX4M02HH6DlccQ72MaGEQPDdn2+xbtVpaHQilEuoexv/ukD7jPcrDLqBGnt/A2
H0NbYZ/JCusetViG7AJpriHNf4ZKNfoR/FUw2S+MKR51Mi9iIWsPxpZ6yuNzqEAg
VwKb8ctbSwtrJzT8+ELQEp9H7IHoKD8frNdcZcREd72ffoGWQnANcssy6C6tZUvp
tt7/VwTFylbBUmHpd3gdtvKD2U16fK1MPLspBxwglbVjkoGXdv622oFVPvv9NZ0i
tcktE4Q/Dnpmf5aTAd4b7Fil+CW/YEb5NGOB10g3ZmrguFY/1P3uWHtnwhTrLfQR
wcf42yf/C9YcszfZ6ti7V317GJ0jU8eWUcBAMuq0bXeBUkYkfm51+x1P2ZRDHUIc
QLZJfUkorbWndGBO4zXtbi/7R/RH1dwdqtdFcYabcxsnMR6nb66cj41Tua6P3phT
TYMZxzBgm6I65PrRASXjk5cWEFDm5HflpsHkF7l1atbKynHqJIe27vMl76JX35GC
U+Xj0o+1DtNDo4B9vFMeb2tUlaYdFm4BdXv6KS7BIa0yZli0tIY8uluBwqVmooBF
CywQRgxhl3YT7PsXr97HrfHZ3YkBuECXxsCkZlk4k2nsnQtWXqMqU+Ub9skbL02L
qwokUrogbncNCg8zlthFRLkUy0Y0MdwUk8it/TwGlP6BBQ63zLw+X5Fj1EPMXUqW
bc8tbmn2FcYG5fxHW9ySRxcPeiOlp/ZIu0G9yHHRC8sSD1FP42jWa/MKXVsGeeZQ
idjGIH7BNwjsK+bRJfIor8FjDKRtvoFSlNXWOEQTPnNby/tu3xm+NxhM35tDCH2B
fk3hozSrVEGQ6DWUYUqxdMcGtuDPbHdn4yr1ilQxZr41NG4CzHb+kxKBwhMSJIPS
fqrbcSdzAZnRGBHGRPgpkpEyaKRla/epaYIOqg/Art6nQ6UMkdZ+/nujJPDefTuy
XDk3qsyonWwZsb6F8KzdBxW5tn91r3/IL8WC/EWKQmTrUKTI15xzncf8nitW44P3
/O8SozUhu+hTsAtvX7TgirnEtpYpAQFKvng8nN12BiwhrJkiG4CUifV0dcVc1CWf
4zizC4bdR9eZJfKhXAP8+rhVE1G6OIFOUuHODtusXu37gIZBZc5LLmm32zDTmIgR
QPj6aKRJbhKlz4zsPc8Qk9FhuD9JwPvJIe/Z6TuEppMKh7jx6ich4OsnHihyigKo
yI9K9egOWor81MN/7aiKHqrjM23MWbuy+TOVbmH5T1gUnZCHmxzXxrk+VUrg+TeX
X8bkHvgNCi/za0rCokqLpt0WnqJgkUeUhU1mKzk62B0QzuthyLMFXRxjcdtDxm7X
N7QzJgMA9mSYEKp1borOVrTDJKIfEcvWwsp82CpCdvsbkuy7gyCTWx6op1ApcsWm
JOEwMuyp563IFwSMQCMv83vqJOxAV9S66mRGSxyBB3gwVDCZxdTEtZUBmVY/flF8
u5mnQN3A1xy9O3zzguPvdIjODuzFYoLKt4DuJ9jXdOq6dygtiKMz1O2PcCKH/VEX
YuZAZPeo4LzNSCCr+QHq+rkPgYU48V9YeJgQfX7ju36dMrr5nZYvjYWQH1VyB3a1
Rf5tQe0CuY+PMcFNNVSMdFocclGrgRMYtkxgs+RttZtnf+s0I4PfqtsdaroVYcbm
6wrZfgXvy1QtyhLchKM7ENtHa4XoN3kSJAmto3g6vmVroVT3PBW1P9ySlkD8EfPG
Tz2CzTuJJpDYW+NEPCbTy49qsmL0C2uy8C5V2vigAcKN4Qu/woDnT/8KUsAWJU8T
uxSK7vNVEwDL8oH2HOGGOdpKmPcjMHvwgSFErzGn2gYCBbRV+jUFllAjb4z4cAao
qjTaav5twQZ0gQk0PufvOqT47UrkWYDQKye0rhHPtoAptGCiPBeCDKT051BpkIEg
E+vu5fhW+4ztDv6fgfl0UekWAH6LGtyMQ4fq1QCrJtm5KcixQ6K08iXkCBbbCuyX
hb5t0KXBFkt4jdXugNpbl3eC7/K1WgaQpW9HQklgmHBobeID7/tKOyqYdvj0omm1
RpI5QL/6nPPWsYDCGTQFC4rpZVA5ZOU70V/lMMujh1uz9jRjbonZnNiA0B901uqb
rd1TSLq/DFmsDmYJI8CojP5dTxp+c8/mh4NRyUtBjgI778IWJWyxZP/v3HtdsRUl
6CXzP4WnNpYCKhbL7OoROojdqba9vr/baHIWFHRzZnB8+AbGasleOFQwAFAtWgLK
30JfXHgHA79FNwQQkHQUpRjejtJxwpQdd6WYRFKBbBrL98nb70XUngDRc3XF80aM
4Xps+zMwLKXg9e1FoUjuQdiEqUazdWA4C+UaMNFfdOkigtFdn30j6oyAIkWTP1n/
FEKriJs6smyspZfVwLTMlBf9bnPFFbkaPI8KcGMeWBTiOHQOuSBsyjez5Wdx4vHd
1lmXsite4y8g7ul7IzOfjJLhgKpDkgZ0zD725luqdm4IMLH8NAZ7gwjRaYRssudF
MG+uLYRmyp5QwsAjHIcRppPi/erkruw+eB+3IcStCgDlqWg/POveVsZBkLcUjllz
cp3kfHKGe0oX570pLF0cQGcw09D/LYwzPM23c0DcNKUkVrM6qTFAGcqPC5iDNkld
vR4ddAxih1sCvbypfIisYfrKRLc4qjhIlVYPYOElEctIo67q3MHxlF3o1a0Ccpww
nbojTu7J3zUU1gZVGDdjTJXrwuwurm8si5BgcjA42oLSqTYQocCxEzuT5x28SkZ2
CjbPJwlDvgNmOuJ4gPPrLGHXFwkGFFnh6aIvngZB8CjcpzZu1MJmUdm2JdGAbCY0
RKFQcPtunw0Bq1IbHkffduXX6nMfy3SBuJ2CN2HN5YDeldYuWSQg2QPDDpoy3VGJ
f65Ls+3kF05ehvCov65U0LnBFKGDjKDL69EWq4os9EBAthJ4b71ZGymKDZMStR2z
7Css+QIx7N2PAh8BUJrHTXSYtTgxFeRAJMMAE4sKX/Tb8xViFulkfQkW/kfvDGe8
WuVnflvBKAK//cEMh4u+I8ieuWkUuPrDPDRHj9dLj1tqBREVhERb7Vdb07UQSZZF
+LzFmyPX/howgfRgHlVie8QJpbObNQJA3JJcCNTqPlnWgVwmBUMQlDg8BvzTbYzo
HR4c47NyP1K4GrQgDHrFOCxDzuh9xUacyBis7lKquPMyJeOJaYG6c8wi3NON7hI+
Ro9WFcAKGC/GfpvaP/8BpXX3W9CHfw6TLufei7zciSAQ44EWFyUyVbtjaFcvURgA
R3fA59UbWvRNNoCA1AK3qXbcTM3ESsD9DzvivwsMkGZOatqA2/+hMY06wiFd9M/Y
l2Xi5h1YNy6JpnZwF/ye0RcqsrC7b/BRtgLXBLgE7sF2QhbKD2OJrloelEAU6DsN
FcRDsN+HS0CETKaK5QURIl2lLX0IIQOtTQbc3/zopQF1Ug6f+3Gc5bIMNHmOckX+
BuWxDYqoy4kr5lwAsLW+xTZxPSTolojm04eadVuzc5wAD7kkkYtXinPOdKu1MNG4
k+PZlrMpnOchDmm+zTACGys/NqbGwJWTjjTjj9+fCc2bIftz9k4DXv85wuQFCZzr
zTK92uk14Y9cc5FI2xqP3j0YzwdkaygNE+Sd/png+5/aMbMJgYcRs2GCEYFhGGe3
HQ5KUZQQmQesqyzFqpqqd0Mjs7Z1hQM0p5dEXs8RFV95ixIhLMl94xnZrWbfxCzX
rIjZChQaokQ6nFJI0KoJXDrJvvo7HTEA3pZ83Yx8f1ZU7fiegyBkdIDWPKeqEDn+
+YKQj0WUw94s9+n0ICHUxDtkpSYSPXze9Vnf0gfsXLDgZy9zPkARSt4fmuKQCEhi
3YESi4lfAhjuWLhDqQKWx00KUvwXhyFe21X3S4Wh3gIYvGWgixrTp4kVFTT4IQ3d
A26+j4WVwH95F6neIkjgNCtjTzsH0DRsd/GCth8AiRHT96EBGI6cO+28JwwiII7R
n5fqH1SROtilK0AKhPw0ZjabFtBNzrDQKgmkRA8zvSgWs34Mi2Cn+8BULXNu40Vo
virK8haC60T8TWQb51fAlfzsyowlWU6HuNZ0/yj7koTdI3m5EWIpHOCCU/6HN5jb
eimWFEkKFRDMxXxzznSqYAinyjZoiDTT7spv0c7R0vieGCoh6ypCVif6ZYhvxZVA
OZrqvxGVpzD7rP30avmGXXLKVw3taQ9jupRKy+40P6ZAQ0FR/LFHWB5IHEzLpXpr
URweVoFI3eWww4nC576PS+JbD203IFikK1u0GLLcgtO4QWHG+K6cwtLtDmcbVO7u
Wm43KLRzGk8bz8as1cnCP9V+5MdhhnOBv5TSck3+I8EN7b7O0YMu8bkENqN+A5fs
4vNufBYoZ8Cvyg8dpVXA0rxXddh5UpvV5zZyfjYIo7DJ8pPvmCoNG/EG5JsCSEXT
NFJvlikcTnwSQsnjBKJnifxCBsp+qj+CdtlJNBZtg4k3swYJZ5CRjjNJNMDP1BAQ
29k5DoCTgAueEUz1FLewBb6TbNxcemvFMyHD6GU6FzT6xQh3ykS9W40eNuIiJTQP
ImaB73zW9+bTPqJ+4N0fct/CCakHcd9o6CvDhviPqmqbwG6802ErLavh1+jXjoxK
foqF1Kis8vSS40idXP0M56ZPzYRI8YNaOkJe1v3MslofL5kTH4dda0WXucQdMckC
Vf0w11MZ7aDXhbhcOjGT31LLAUg0tJVwrGda+mlqElB2YtaIBdO918d5MT5H8iOF
xtVY3znTiPzEvcOe+ol6FjYzGT6oFTA+NonXIvC8PKxyDzBiM4xrl5RJBniCOB6D
a8z6hyqBrXU0aYENXLjlPbs7ZmhRMVPykCyMxOaZtw4uOto21i+Hi6MNrSwKJJ/E
ZXc1ni79LUGx67dnfxu9epfk+bgfIVfYsyZIMk30BKwk9iF6WEirSSTV/ygap640
4yNJ5wv56ffAfqjCYipX1w5gyILPpq2qPJTLLQRI7eZbI8wAHmUPJDOtcY96fCWE
zcCVmGcf1p9FkNNLzgle9YU9DNMiOY/JfYbyYVSnUh6tobiz+2nJVF/3NwevyQZu
AuUfNTdGbuT+rxsCLP8g9lcuGWmurKEj5axnQVqhg47sz+IgCpxdiK0SfHoqVdg0
dEfd3qRUougeKlOZCEB/Y3bEsM0MFXwTLyC22JVga2wFEsnJtF7N7LWtdJNJuICV
0+D+ilPMwy0VJalZeFsgmkhsrcXZUSVj34A9mo55E1RcCKQg0c2fOIR80dxPl+eZ
N7SaefmKh0+GeKTC9fpXvG3706DH9Twe93G3OIIlFxJ541r4WHVBuc0YiohwP+XF
qt4NlXEz3tZDb2D9h8sR2mb5PUotqjBFI1klD1N+QPYs2oaJzBbSgfh3IJ6axQ3b
m+3A2PYtW4C0/oO/QmDNgDz/z90x6pELmNd+4LIW7Pu2eXlrLsaATHSjdEUMUZO8
rTsdGzblEIpbN351asAny3JZxXzXhSWrm7Kj4lWMqShbmRA7zm8ASn8fQvWOO+iB
8DYI/BKHhOdT3wa9UVc7Hxv9JXc0s9JgukrV+IYCbR0w4rE9StB4I1b7cdZJUoht
0/1VFhbB9g2PTs5pWvGWnLbfCj9HMZHalK/3Ga5RL3n6DPeqcbQWbNeO7s4ozRN+
9JrToV8jBqd9+RmMfqFf0hJCHeJ2VkxQP/oCU2N8a5A2ysA5SOdIbU0+xhvNb7Hk
T0ucGbyep2hR+M9TmEZ+6NdKrDzCaTwPZ2J8fv1g4d8mgpaHzRpNlx/xvG8ZqLIS
HryQYr5ozNaaISuWf2uvWq1wkj3yXoZH6q34O/VwSv+lC9s6cxryVZltxdyIJxsE
hTyNtWIY59r+Kzz3/b4+FYHoKJuKtfV2yuno1d4ChpYdNpqMqZLa3B8/k/e0k+l0
B50I3TJcTzszF3+cvJ8B1kNfJlsouZxO6PvdkWGg1TE75OsoDd6OaLSj0rwePwRv
JwyOSTAHyCfdgKZdNSCQyDjs14clAsURU5KSKvhPGO/H3lYNGxqnyA+iN7BuY+sE
ywFZczaYesFG0kQ7+1Hbh1jEZDJB5fymV3pn/QcJGr4Gct7NpBSiPcBPeb/T+sPL
Zvlw64s4cLNe8CBNtBd2CwDocALNYtHzizjVFrAzKBDG2W6aTZDpiWPTNH9IqzjJ
bn1ZpD7AOkUe5zc5jFQCcpeE9PvQO0Yxdv7xPsgIexIBTqn+qurwzgl56EZXznhq
geO7VNWuhRzSXzfiIlZtrQDelrlc8tZJRxyqAsrdBAwSKOs4CmHLCbL6J+uIhRe1
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
IWq+LyDJ7F553qzRqx+wS71P7vMFgmDzB1IEgpsARX2SZHKmgbSIevCyJtW1KWI3
BioOZB4zSVgq/IPrBM98AeL+pdXADVD9qndmSszESzbOcjZT+fpxVQ0KwYPtJHsP
6Z9Kn6U/FPOjbglOc4xSik/XWFs3Er2G9qKALc6EjPs2k2w5Zp2S8G+feqFsphrE
BP5HbUlWAHjH3XkQ5vo5x+0qPBWBwA51yl5bczIqx6LNlPkcbUW1HdP7JAcYNBJA
P+qRS5pQv1f+AX0YOfRG1LjiQ8+Jm+61fGzpvjS5eLDqOem3UeHTx3S7d7vyZWI4
3trHyYJtHApfcLmz29iRdw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9280 )
`pragma protect data_block
JSepR+XAQBhwdyR9Y06IPggWnS76AAy7/sryoGcIukn7wvgdZK9As/05Q1rJJdmE
h613r3LkSqlllPk/vFVA6KPNGMMLPuZQoIRvJfC1+ftZZD11g0YVCQIXTBMqjMpU
jGy2+MDasGvcHtz4o3iKorq6GT/rgEyVurR7sgblOFOCkBjV4//Zgx2adk1Yxc1f
rfiyJrugVTc+VByNqvnQ/1DDA6O5HqEBmXb5Kr+eayCVnWTr+s0QevEOkGOH8b8H
DCRyy/uN5qtsAA/7PfP9Gz8kUtZB4NWZeetTtvGi70Yf0BaJONJ5Kv9fIEVTovnJ
ZOv3DeqERH8m5c7f+OzCfA/GNq05MlQaIF8BkOEnIbY1N2YOSMjSaBOTKt7G10eW
tajczOv6+kNEexHhzRd3/21eWcv8ikdT5MozxGboEY+XjU9A4RJVeLehdYMFLA1B
7/EIJ3gm29yrqHBYCgJuHVvVo16NKI3NXSje7WWgv0LhNXU2STHXTWWdbIJdNnqP
P8AaVl/bOOIN97YoYYjBgQw5MQ+4BVgC5Nk9q4hqLT+cCYewGrLqRtJEsy99YSsa
qlVLCa7A8p8uBQh1A4ghNaNc8O8XDJ8E4m3cNTsUn2SQMLslxlvTRwARILSPbu6G
CznV+45ETFLUMR7+qCu6GI43Xlell+v5mrGYsMNZn6/ilNzqudu4DA/5DJ7EJjEI
lggIleH19RpmCpx1C356ePYtA0T9AbjfMWFYD7CiGUh+AQv4uL5/3wku/HFOIPev
yeeMzvU+tC6gwyhONx3eYcA5zJySdm2JdPamldLeoH+3IYI6ia2vBj88CzFCy1Lm
791Z0OJBsoPahFxJ/hkTWk0aE6hYfHaLpIAM2AdQtotRDJJo7tDQGUezErmR/1t5
s4k1aOqtfYEWGiRLY7UOJkYWl+HaTpLuEgNWjL4yr9rUGaWaGd2jNf7lNraPkPfu
Y5QObVBTyzvdTeBg5gI9LlvX3vUPLAYq58guoJYfvnyYsUU4f/ocLckN5ap4cG/i
oApRzmYM4qNRjxa6BpEolel4y4VsLX7N7t1pl604hlTXAR4bzZ7WCxnagoQjQIIa
+L8PcXm5SRaqc5tc4ze/rTOy2EPnUY6xAF/s/8OYfaRuIpJ0R3ZITga/1/gwncuO
8hAzlVpulymNvtvWdh9KH28ydv5CJTQW6UUqCQpDuemgiqeoREsYbJeIHUwp/gg9
2WC64g2PgpPCetwKlVzcA4yDNLnoBAqeYgkdDll2rcg8+1fGyqN7Gw64ugOkJFjE
0HhicXrwoAxAcKVnpArd8RgViyqP58nCgkUpoMevzq9NXCj1PGEtcjzmdAJPca2L
ljqFknMXhFr3WBeDpK3LkSi4dr4k54u0NfA4+4RxGItGPYHMeTdQ7xy/T0/TpcXh
alkBmZDsXBgBMp/vYoZjRm4/gsKfvtdFXsxst2yiHomuW/nkRA8hkyEIa1hcbbIB
BNER6a75mWwIbogM9OasTEelVXPttYDcvhDV/0HOIoZapOnu/wqSkO/7zuelmE5G
+xYVD56iRHPmfR83ogJxLTU4u76dV0iqQhPA3Ra/ap92Gim6CUJhnLwCDOT4o4SA
rq8go4/lqi7mMHYjPlhzN32JA4AwxLYv+MfgmNfDjTKBD1ypHA+fLhrWMiLMQLcA
93Pv00L4KnmKLu4NOQq34aPSMiwdXbP8PNIFdy76IJSG4jooZTyUpZHscv3ms97Y
Sh3DABftuuG/HdZd7VLKh1OfMSqzY1XHosAbyOvjMmCoXcMpV/sBoeyW7iY3cSVt
FjEKuFTdSflgSNlU4VmA1mWgrq7KmaNbs2yqOUJWs8rdao8xkr0dasp7zGSw1hF+
eaVkGXJ10GcyaAGK3Pw2BMAjgcdQUBwgEEVFI1z9qsrb6ZFuxwHUgoBV9OBE0t+6
V1jw00eLrcUaf4gF4zYVpmgDw2RNAiq7o2Adcn3UkYZkKuyVFQKL0veh0BKWbI+d
zX9eoIxuWleMPcCad8y86hJOtTss3kdx9cB4oOvTtPn8qZSV9t1rLYXdJxZCeuyx
QuPMf3PrlcGNouY1zkoXCJ2S5ITXlAGLzIyasXKom5bdks5PUrTVcLpxPeWB/6VO
ZQFEtBDkzH03uQl4e7makPVZZlzhCLQ9YyCLEHc6q75U1qZSkOX+zUaVj1uNVDIQ
loScrFptPHQUIyLQCsOKjchEEQm7huySVIw4ccAlIDA0PJgx9eNIJAmGHJo0ru/8
LoffgxEacT3Z/D5Z+HhuvFjASVfbE80NezcRpmyq4RkCSmt/lD6PpXDOXRNDGbzk
R5EOK7f3HwmYjFRH5lJj1//voXHjUxZcvYDdvjmJ8TcssKq49bUrcg+ItYxvACy7
R9/acy5Gep8gIUohGTA5iOLX4xv7+Gz90JmMKNgO1XPeE8UKuEyJrHHQnirey5/t
XrrdZTSATPlyqf8C7ipv+UV5CN+S+DJKmrFXGyV50yMg8ltTnDVp6cl68Bi/IJQd
r8NMikmzAYFAfSvajfUXaXAsn4fmHS6WAbftBdQOStc7y5rYMvBc9Q+yTtU+tc4q
bt3FFt5gfyGkHCAPYxernvN6MV+gzEThGLtp7Q1WESsBO1HT2/+yY0u0i4Vu3Y98
fb9XU+ts8/iyolOhdz+0ywxh2Mty5p8e3ZFJVYdhYz6HYESttFEsaoaRiz1kachm
5hV6B2nZFqiSupCoh2GJe+ZKVTDsuGDtkX0WnV1W3abl5W6RMxUjve1E7GPEQJHd
WyxCiDMjUTIytL/BG5DoqdcOLIdSB1UvLhA61Jd0V6NvKGu+RK6OXGGUqLx+ZrX3
0Im3bopBHNbiwQsGujKyZ8DRZ5aL1NFDRbB1fK3d6vbddkZHdSbgAiz8+rIuJbtt
Jg125bgNU5QazaKfairJu6IXBoXK1mAGKeOc8sGJNKtP86LVGftImaTkowbTS3zj
apEaaoLr78GjyVu3CWOZIm8cxTFfi5+w3G1/dfVMurQyhKEIiQy7BFiNQ+vUjAUw
85hCaGYVTMJc8i8edFVluJSZ6HJC3umJ+z4FvB59c5vUG5TxQ0MCr+oZexUiBZrq
KpqVh3nvO+UVMlptT00/QHyF0dPEsltxfvc3pp+snknxzHINsaQk84PK4KMQSJUA
/ppICryIGCB/RrR7fHiBOGXgdL4CPGqBrj2FtwWpfQ8B3LImLUSi1GlccaZqDGuU
XzA5JBgVW9UbiW7vGi1N1yVduXVJBwL5edsQmsUKx7yzimKIedyk0jBmBZc1g2ul
IBrNH0LNitHm65vB1V2RqkBnmkPzSDY7A365pbyYreV5IYjJfANSYVtUU5Xu4YSm
j+lpLodpg69fdnIgeymeb19aTfBuE7+LWGTlo14oafl7rgUWan+VB1eJ6uHNjU74
eePljDAGBgnzNFyU5i5fYivfgBloAXpUaCYCghfAGLDT4LKRl6lh/6PaxeKtkCWT
3pzWaIMUQ+Yd/VVVBlVQPBDjk+U/qVgllxahkV8yMU2OE45s/doomzC528/ZF4JN
TX/pwMNBYxz2m72At5VLkgvl7xH9EG4ALPu2uLd5eGPWU6woLLprw5klhI+3u+wS
jjZRmfmyGZIF6LxvxYl+LB7p5bQKmdzlWsn1PaXXWFXzNMGaSaBmgWSFcccikKQR
xziZgoKBAWblYu1LQqRXHh/Dkcmia0+0gz2EWhNhBBNOf1GJVNqkmqNRUqlDtNN8
YOlJFUmcdc1VFCfapdE6yQ7ll8YCEIFi02jLG+r9Hwd6bhch/gWz+TInevhf0EBU
lzx+DwbS+f7wNyJ1AZKfnWVCBCeMHQoRtNtY7w1rVGi7DLjuRf12xdpVhU7GIsO9
IfY6/KLD0e+wKvVg7AYe7XtMVH9YgSrHr3J+15yiBsA8Rb0nYaUzhppLFdKWpRVz
GKZjwyLydxxJZ1GeVeVkZAosJkDSicbV5P8/RuOk6i9R49KD9nCY+XHmNb5llYeF
Xy8ChSz/2KOlsDK3L9tdFHKBnb0g2kTa7mU90hq2y96Inbv44USBfpEl2iZnPTtX
24PyeyVkxbewdBjbUJXhsAVo9ZxM85eifthXcCATVWNIrHr50Pn6IeX0DoaYQy+M
eimfWpTXBnPY/X0qJfMVOWFaq1lmr9hIsod7brdqNHbSRrJ53mieq3/yawWwxIH8
Wqm8MFyW13eljKzBseHU3vJAyPoaHL42OH/VCPeGeZmTMgFq5IKGDLZw6Jg11sIo
xRgWXFYAPUo2Js3p47g7ShfOYrQyka0c73u9Zp51oeVRmyvN3o3XPis8e5kKw9He
VZWr7OUCP1Qq/82zRIrSS9+aQTjt0s+IUPIfiveYhNL3brZT8OyEB0G8gMHwuHu4
omU+db2ZMqG+no9iOKhE+AbhBVwjkiPHwhxjTMQaCsYDRLMdlV3rZUsYY8M/UyBE
Fa9JadZxYDnJSGbl12vxa9bWGEBSmMCP3E/9Evh0GURFYWv7tkKYS7TTaaomlRno
thBhU7BNwnU+2zQD+NtW5UaVFY0HUOKSpO6BhyxDCyFAyF4o9ZcFzIEGmndEfUNu
GR3/7cwWXMWxhwIeQn24xJTANbV14ig+Q1VKuITfVTZgqXnMAAAQyBYwRXJDkRka
H/7HMTNjAYNwhGFJecjtSK/OKqHd5JSfUy3DRMvOw56oIE4HFUPxjFVuMFK3YLuC
cnogXWTPkBrY4UVQHcGHOYa0EkM+rrKWKC6kNCTYBwMeP36PaNRkmEJdSufWL/ct
F1d5v3E/hW4du5orkp0vGVVpIHIsJadOnwTpfrojsTrPWhdQn3v4i9XNmgMQ3qVb
0wIBpNI0KXRrEI+Hed0Pxu7BDM2Y5LX5jQeeJQ+Zm91P1ioCfLbdaJiCtwEeedvD
SELrqBa4YJC8k96wkZnEVIfbEKEKMUxmtaVvt5LzN6hUEPQN9Np04HMQu6rLmNlo
89J2AVTM8VFIbHa33ouqHkFh9CHaI38uzO9X7VX2WpM9aO5o4xYMQAMddKt3c05M
UsBs14n1ZAAzt8Xcl7u3GpXaHhRy+LXTZ1XvtQb0WeD99EkPYvCR2cyI0tI4u1XY
pf8H6fmlPEXVhkbZHr2Oc1tOJID1+01reX8i670+f7AnJ8GFj7/grd6idLhx0br0
dI++XXoeaOM4/77esD7fQZYDtduMLK/XvTJU5g/kXunTZwz3UNcH6hwPhn+HpBN3
qVofVEA76m678zmCfI7+72rt08l6OJ3fBh5fCko76VpewZKf/gmAcD0RqdumhDnu
+YclMnkN0sPqWDrt4qQHie25vSEBEHhUNMZ0OmansaRRJXB22Wt7qovMuB6dzu9Z
Z6wIe6VmQ9hpn1ASoyIM7wTXaa8aK9qnpci3lgWkUCgyGBJVVFguPIIee+4E9ntl
DvorRYOxs7PiJqUKD55ivze1Tqh061T172hPZQ2eaRWizpdVgyrn1JJm+bRraXBg
UdDjt9lwdf8dYrn1hImVgKEW2mU6FniEDROJVol3xg7rpBtN9A97fRU+I6dZSgoN
ftHXKD5mOE4M+ZE5Y66d4OBSLyF7xlpTR/WgjHCqhvCsfFFZleIWelG+/YviNFJ2
fFdX/E4f5DQd/+X/K1/ZO4/4bZfWX0B75+Z+6LWIEQL6eK+KMIJbUgkwyioO3uzr
+W+y739gumO+GJ+slwFbxlbHdZmjrYTD9uGSc+YHL9dG3Syorwrg9qDivU/TSuAV
cQ+Q1jo3lnYTiUXKi6dKTaYxElMAmI49lb2JGEM72iwxFaCemMZ6IDouXKJ7zQca
t4PVXllSLeGTWUonWAD+DpMsWrJ7cPLPmmB76wDf5ZOgeDjAnK4qzklNu++SeAM4
cepZYM99PzjB39hvqcpWEq9fsdm1v6H8QZN/YsDMjB5a46QGVbwvK4ZJ9xSSYKAZ
ZDYffWX+Vt5+SEh5OKE7I6EszaYMTZKtZ1SIaXXSmUmdZ0MWi2v1WDh45StkeSgT
WLBL8meRU+QqKLH7Fnywzgf9i5p012IVtkF2zDX/aqU2y/crjQbbjSHOgIkYGeMC
9kwu3LvOLI2UjCuLFOiYrcfSkG2y/WsauAtNG8Ek0F0o+g7l98VuQL6Exs7ML8ml
AHUQcjHvZKd/ZSunJsvmcUQwMhwGXEJFfZmGlpYnxDlcoDCAPH6HnRaeDwF0pSgd
nSSSTgPq0sjGzUW/Uv6VA/hPcy5WwR3Qt57XpqaBOGU2LPAYT8AoxrQyqNSZnF/5
FYQVclk9vAe6a4ZmJRI98iv91jwuIIf3X02EMI7e4JSjnTwTHlLi5ffyH8ol72hy
YDfbbLFAl3MsR7o1c4DX0afgmdxtlQixHyZFYMYgsNyaaJZv0bBD9XS0jeRLMc6e
D37Xo3YPKex2qVsVtHzGkkVtEJc+R4TJBYQx8dy1Wlok0dR3uOCYO4kPNeDU8lag
Mgq2md1FD+cs/7Qt7Fsx/TkKl1fDdrh7/JiTxdtFnQc/3kkIkuqzO4LqjgOMh4Jd
BM0dtRPBnQ+ueQB8030CUd0edKOF8hz5UoPb59QaOmBRVuuu+utaHXq75D9RITA8
JdkupOkAkVNUffekEx8+V94WVwRwUZoZIruh17HZqSKHWSxc0otozyFCIHWRiJDR
X9ATi4zpMjDNIPSZ0pIGBzJtZ0xz3PYjqrcEOotvBZz5YeIaxLJ83NlJN/f6XP8T
8mPXjwaQHFNxuMvyczEZHHtC82fVJix+jTddLgA2LI/qf/bpSTUrPiK12E9v2ClK
YasBIoPs+knjieycTX0psNF83gfvUwKaOYQlHYHg5uqkpGCy1Lv600WbOVU7P9gf
j8VP2+v3ha7J/a9KAX4JBqOsp2TKUDqh6P/2ZwxRwum4f38ilpWF5VDqMUKEO9Xn
TWuJYmvNqLDky/P/Dg+Uvf1RN4G8Z9se+bix57IbbsmpcRLGKIMR5wEmEEsBBYUi
WklPADgpDb8eu+49xlBxSq4o9eT8Qt0I2vreK4mcDVpB/Ghe7yFgKg4tDEnxjFko
7VbwqSGQhwgzLWK3SizE3kcsjSohGH5VqSYlmdOXJHMyBexz2i4gisTECXEhGY2E
S9Euzf0GFZ/VGJUwZdo8NI2vASBqd91I8Bt3y50+sCPRdgwS/Kt5TIoj8XOCPFIH
fuXDeFASPnxa/cUHxoJAGO9Qv9Bx8KbBFvRGt3NJXpeeHWijkN0NTmGxXAvLLojF
a4mkR43E55J7QzWbvB5F3Pwc1syJGZ+S4Yuv7ID63Bh+JWTa7AqHMW0YSEzJpNnH
MybIyTrAJsjqSD9GDOZT+J+Hr7QG0xehEBAeBBqkzCi7VjlX00H0jf9hEfT4HhMZ
NWMd30MnNbRIhWmoIJ5wLPEjP8W9PcIcF8NvTgmPg7Hc0msLWdk+x8zwiyS7KsBJ
fuK/Q8BBMEkYjLwDSisU8pycwa9Ul/6142/679ftDJWV1XL749RurtOYCDDfbYm2
gyEVKyLd/RUzGG5WrPdPxa1jiK+qHcH9cOHeVo4gMBfoWMbT6q3MlC6WMDMNpKLe
h53C2ICgp4NWsjhTtYDSdjnRvzgFzIznq90EWw8F1AqduJh1mSB+SmQ+hHL50RgL
uk0e3pyR2ow9Zm4AjqKiXRmIwbnoFakO7b+B4FBvYKYIHS2/PXHhvhS5UjM+iTBB
t3O9SoVwVg0Du4m2UObyLPFLZJ8sKjiTeUeFmxA/8asrcypKp0sKD7ucb+pfTAu7
m0LvjpKB6kXpEjPuB2h4sRwKZeKAVxP7wXUM4U/cGMFaTYKb8AHEUtpNnoMkVabX
WRcFXL2PIfB4VAS4DWQwtnujuM9978g+5t78P3k0ffpReQk8dZDgU2CZxCxLR6NN
Tp5IwULLdpl1zypUCH+sL1XUMKXoWV6/XBQs8GHuMSKVAnwWYuKqUnujE1bddq7P
IyLuLFt8jU7YcFOUyA9imsnBoGINEqvAWghCZZTsgqK3X/CURMu/NIGQGbf2gMig
9yAwUMnzr9oSuo1xrIbJGcS+/s2b9cWSnw4dc+vXzTUAURdnGOifv1fMcCf5ol3h
6lOX4/nzHwJEzTL7fTbedVHuVOVcel6jNRGAiTl91UaNB/N1EwsehOEsG5rSCimL
0WUwupLQRyKgo8HI5J48hI5PeuHcbutX7WoZwcGWLgicwIVX3sIj0xCH9rXAJCM4
L+MdzqeEbwWGxYhlxhhnLC3+zDLboSwO0pGKNgiimd7Rr53KHOS9xuGDWfnQtwmM
zigLyZ4GUgidkzNLkgM73tQhaNddELfuzBlQ8h4S/GwsgzUzFX9fmeWQ5tlYghPX
XHVtOMA76Sbbvwm7sk440pvdqHG1ZW6S/n6Uy2vf6eAfKnss422i53/Pv0wuCv3a
t4mZr88bB00sU2f1VuOwz4UfxMA/EXAsnKXseU6STuKLBYF7eEBTuuVSv7M251os
HJ/cyWt2bcoGerHkUNU+/Vz3IROTPNAvYiAaq1a+OiHW5pjm3996RZ99jIHYTPhX
Bx8JV/sShOPk6DZw/uhadcqZKHxc4R2lY0KmtZWw+PN77w5jj1L5sXBci6c4LLtn
1Hb9ze1DChatVuWKC8I7DiHu4R6VEr5LgeJ6jaybyQgIHxLuRy734b1i3RFzP4K8
8Vojx0+91hSzb1wleTPU26r0dhSNsAevYDd+Cq1MJH/KcWfkRJjDjItfIFXmBDC8
0oms323N787tCRZdvGUkak6giRBftzNX8TKB2ZSlJnMWqRWWnm3eO5gT1LkTN/Ut
UHMTz0mVp2KFJxuW3JuQSniG1Nc3+CrwWa8uXwLy2gTbGbyVJqONsW+Kt88s4zIM
W+LYvSDuwjeptnmacIIoBhNz3T3Gt8kwyvzgMQKB7jZTYtWOuKlIHGRzMBcmm/oJ
Mkl69mfx6k7CS0iraV90vJqpD8jklqd2yzxklqOj4ViPuS88DQyI72/uOuACBvHS
cdRLA+GiHdS1mgmq+ZbeeICCdCMN9v84wPISbUvhCHMhcWFZcXhYBHbCjfLZw/sw
4GbKgBsMqXbEWWhsFjLWQmXDxCtqGLKZ03aTAGBx6gvy/1KlsxTTHrm7IWq8zlcf
FVOXAFju8qENwPokTkh/E1/lSV17XqFiPuL0VZVmnYrTmxCBzyM6eoIMV5yiQFfb
9oXw50YWPRTdYY0d5/aFTNWvv9CHHqcdx4WnZB0wfrJ44MGyeYCSjaC+7w1Yn3E+
StnKfcvnnIXYZFQ4QqiM9c5SGrkeFNtgrpW0eIxJnrlQM8HQO2n8bcQ/uixaUXSC
o8JPeQ/YZgNEzxex/3tOMpnu/PxFZnupywrtR2ORTSxX/SomVPeYzMjXMmKkdPwW
cqpUvMMUErUXleWgOISpcXvsSMfOGyJPkA7OkSAHdymXw1uuOz5pNzFUceH0sT8M
itxpfBCyHhH/lgFNa9bLvOyGIgSKNQc084tB5qhF/JIXQX6mfMZWGOsA9VCKjYJ4
YGCXKnZyKE/7ZmDpV9eF99oK6n5gHmlnRCwYiy6OpmBXMmsKUEtanKqrtr+/JQX4
VLMFaqDGcdXv9nxPFOSduSAJZ5K9oGMYQbiVWrlm06nKDNXW+/GVYf0L34ujvOcf
NPKrzA7qFOv/GPqlaT7IQ6S6HrT6yRDQS0lvwLLLOmanFrhj2bChUaKlg0X4rAB6
fNfsAHxGCL0pZSVG3Np3zepQwKBawHDMAZkxu2/D+2LRTe1B3tBlKo016DpZ6qEx
H0zESQjLjL4pqk7EjoW3Qqrz+ybSU9ee0EnNwdn9+JtnuUyZSIVDGpp6EjIag4Ck
7/NMWXtszcgKf2HVsienOVSvXRGfGT8nAXDvp/eZWQGoN1lZCd+lg4O4q5kROBX+
FJeepSycQ6clxoMfUSzoLKxT6tXG0G3JKXXVK7cI38tVh3p4VGtlzCw8KW8fNdCM
/sIwsbxNBzEAD07guHiqip3PNQPaHwXJxt8uAcR5WlB5Nz0ArkOKQvZt/YwJ2WZh
NJfNigUvK2rPFU/0f5cPR0dpmGodlNjqsZqrcdk9LkXNDZCNpwARd0j008jPfzzu
1yT1zXrOAoiP4mW0WSfvA09BEK+ksSPkClfnUIUFir3NYDnmrebYMeHuHVKP2Tsy
+g9Js5sFqUSJ4nuKKchOes1lKfwt87LPvUcQ0hj3ufY7o2dpiMp4bKaTJHhxrBZx
yT0rfCqwShKLUEozE9YwkpWotqS+SUmUfW7MoNOEjUohVImBxLIpMGrVcwIJ+Q0o
XGK5wWI+KBvFiEquVssINL775zOjyc/VTHUNLL5IU04+VUqVVjp6OmqtQT0828Lv
aJtuQ8ZyHjkiEYqCSrURguXA0TKcwk9xlw8Ic1PFEdeeQwOUuWzacyKKtfgfDu7X
bSACOkzQr8H9siZZUiTEiuzf1CxzF9t/KmS3e21Y0QPmVkewGuMPeYEGvyxkTiBI
UnjeavM+bwmdmfv7TY3ObG48cxpVuFS92uOO6kJZufjmwfR5a5aq2eOjcbS8Dava
HGkyH9G32e9O1Mg+r/O8Sm9/NKJSIcKlJbtNOKxtmEdpfEMAWFRc1tCIRysoSPf6
XkRcBPs/4nne4w0JgfRlYnRWB+URmFQdU9MdQf7uGg2ow/xfyn1J2pTKFag338EC
6vJLdHlZ50gjfgaREz4DIMiaj0MKOK2N0sBmpJ/dksVkNjpBxJX50QUcoawcop2C
6JshuJGNdxWm01XeU3bzu7zUEcPTyMFgV6kwVNe5zEgqPI+DHDKNkkhNRiSglNXW
HLG4DjVbeDa+ouTTvny4VDVJFdZCIuXyEMlG1qzkGHu/C7McNc/v6FZnvwM/MyrG
jAQhE8aL2qWwwYITMFhqyly7l7lAT9oyxlISCFhWdcAj1McaRJ2HMTCR/hZupiAE
+OvgSPfwuOdrXdPwfwkA5ZVHm9SJiQanfV5Z/05OCrJKZiApPLiyX+kDvAQ/cvLb
a0Wp3X3CE9wKPAjlcX5drHQD3vf6S3PPcRlN3NGir8zXGy7nckfF7iHVknZg3vDP
VbdQBSzG+UC8Mv8vu+WGxTA9Q5y7s0qkmVh6dYjRlG1s5zTAp3o/hK+gDo6vNes7
+19snFVUb9D3KLACPh9KfB5TNPZzwwvczWQJAPRVg0h8XwX3xCSDwh1H/XjLyper
/zU7SMsR7C7y+S9wqIL4ka1pNwF2kRSUbgpln0dktJkDls4KUwSFMKr6H1yA/nRF
BkGx+D3yGodJzF7NuIqNKgaD0fQ7y43splyXLu3+QbAn9wny7XrHYR8WBsLwERIH
G4aChs8myN149hazv8ZmVepug6TqAymqFoJPm8yy6J0mFHalJ8GWbaF6iU4RdkSQ
okGpxyDtsw8ZdxEGstZzB551dZPRGlfsLlYEqcL9FooZT1ZPy+9mvE9opnY/EhlM
RM6R0ITj22iyHWwkVZeLcg1AapVG8eycalmEbYqN1TT7dq9OwAjCZQD3cdNM31kN
Y0KcWFWYU79lyQ5JcjEShpUtDa+eLBVHsvoXGGr8gr7MDSvRoJkv5IEn06orSBZp
2Wtw/gKM9i7XgpUHQaaqSZd8WjwtG3U238PRME1DvkU77sMwiDOwp42v5DzQ/TCv
nlMzgzK/4V/mRs7duKCo4B2J0Xg8wgkr/tJzOktx/cb+oZG1oKjHRfYIhxxlxLfi
c4XVaLb45mB1fMcnMeszkVvmFiYsTUP/ilQLC8d25saDb/wkv7R2Pbic4clEBhJ5
FFoOQsDdPFO5gcbfcf9Eb/ce9DGYLuLio/tdpoEPheKTjKU/3nqXu6+jVi+VKFcI
K8qzPuhCrMzkeOPqnjrDNL8SBK27Lnn5uQu0XswndljFDdhIDRr5JSoO+UldjCRO
Ucaeud2JSZcoIB8a1UtwLrXmQfFp1rk5R3ZPA/O1HlzJom02drDnQZB6QTJh8ULP
n79WGngbZRkTGcnAi3rlJLdB6svqjcn08bpBBw4IQMROfFf1wKrkWuHSONbuLK6M
ouUg0IGBfQWCwwiKMCAn3IMR6v6BX+CKih06TnxFZkNxX+HxqxJEOs9CTT+JTpKD
D22mgFnbiMqcEEvkus+TGPYjuObIOb2V46EAM3Xx5uer/GqfGTHBRyHJL7dyjwp3
RKQkIj+in0aDrpTtjWYHBMdu/W21SyaVpHwZ8OC5eNUhjJ8oGj1mXISpkhY1+Nru
spanTF7k4zc1iCHtP08HjWfDvH9h9SnCXxUJ3Dtq55pbW72L6hgerMGSxD4bgy7F
cR0T1oum/RKhzKrWKWUPJe8/zCPiefRnvT0OZhw2ZXYQiAWbUxhBRiaDognZjf8f
XCqVwcXMdkDuG4qKp0ep8x3igEThFqTIUqvZCv1W5GbzLgoVJMQDbxZYePM99aRA
fkuIHg3IUNskVuFbT/U2pxgFlVFGHsFzgSwH3a/3twSPwuy+Y9oMHx1EbBuiEqF4
JQTW1YGkNk3JlsaQZvSRTg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lGqzS6ZvEeKXVwwU9HbtHJXO2qqdybtyGwRQCMuPBZ/aqd91+dIFa3m3tSeumwCB
xPNd5PQtprmePS/cenyV8/4wX3DUmARSYbDFzH60iF7kYgBfhS5dKhcxiSPoLLgH
8K+GKp/QlaKdQXyPZE36tRoWo8AGJL3rydjN+Wzm9Ab5oaSXRwUdQt1tSSgjJq9q
+e70kze1juWBStcO+C+qvHwbL+4FIGgO8BnJwE8lCVC4AA2+pCc6GxMSnw07N20z
5q0j92D+4PLxwiw2bDxzQlS535SI0/X/PhSizXj+VOrFFsyH4QyC9uHqr52izW3e
Gs6Ex13EA0etxa9YCvOiEw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
oqIPyJ1SO1AzzWazr/zcTGeXv/XLZLtqsgHk6zDoxtd/7zwbDPU6cPXMOvb9No1S
jeGBnVdUaKG6s3aTFzq9/XoqlttjlnvZcrszB+Z06nUypU8bw6hdzgXLY9M5gG+p
vKwo/fD+oHNYvCqnIyOa4gW/HBJGQiDdRMaf7dftgXEH0bR/1LV6hXIZLUZlJekX
PlqChfTxPGDT88VbRtprPaTj3tFJe69LsuBD3RoQYvCBwfdtVW2E5XbrnvNqYDBS
MO4d3zMje3DA7G/s97m72JQmplnIFUTJ6Q8m6sgy5/0yeQgqaTI7WnVja69MMLrJ
Zm6H9n8LqFTevqUQEpDacsmkhbw58LITdJAN/UeHj5rbaT0eLNaRYvAt45jHlaU5
aFW+7npI/scPG2NqOAQGmm++t8QszKctYEjsidO8Md9ZSRNBzmeS4PT3mBiJEAGF
8WuhYdn3AyjFntMtmZ8ndPkD1zpyr8SqjwCklpA379Sdv68DXIgfQsF9L4HA9u4V
/aVU5PdDsrfVwf9Cz9pEUotYxXkEVXMTyrk5pzLkmIm8EzEYsuzq71awtm/SN8zE
3RhJTlZNN37i6vPC9S9Pu3KaGY7QBLrjqCe+26BUCStR4gUxDUUbaeGNJWWrQ5Se
glE5xVESeOJEdfGLHEwrMskBM7UeIviKO39C/BFhT2LaAPJzdOQhsRga45E+SBNA
Gp+L/J+zwzrKcGCfU+crWAkQ7H0zEIWXfzDwoIq92tNBROzTFFe3tEGqVcrsZNsV
q4jnyyX87xMAkCSaiuV7zluwU/QutFBKIGLvYmnfIle5GralX7/rjk086/vKOF1V
vB0k+tF5Tv7WNbIhOg01wIB4STFioZAd+nA0FIID/4gxt5mj4wLZlsuu4f+LtR9Z
HLeZisGOkoKtgD0Ynj3swqIC0w70VTcgaE9vdw5ojHGx9CYeHVeDm2J77Nrcw0uT
31jAJnqCacX8ezFFoA8SKLTi9V0SCqSfxBbMfyXUDcr52BP62oTrTpOoXtBemrKl
vORBITAkB6VRYzCp+0U/KRVHzgbWbFWxGTP+l/kObpHSHxeEGNN6FOpkIM4c+Bfj
+SJHQmXFAxopBpolJuAsxdLFPy8TdQz3gBEUpkDklseBJ9hJ5vUR3/Rh7ENXVsHX
GzUhL366VuqbAVk5TapjjJd0j6gtkcsoZXInJUcXvqqweJUIpd3tYQTtljWG6I8Q
oAR9IGKYdKXRojZ3zrTAiJdJd95JwjeUCZb9OUdoxpTKvth6v0W9vVSLgw7e86qY
87ASCO5oc7a6Du5vSMZ+vLOj4/5pXM+oYPIjjCBUj6olpxlWZFQ10KPZ/If2RfJ3
90dBEHgsAqqQMsKf7m33a1bAO/6bke8N7/oJ8QWMfal6XQVYWn7nT8NRMqg28gz+
7ARZ+7FLMYELA7psVbsPi3/DfNvnQHR/tKasn88VLbSVQpIsbeX8fUiToxCwHP9b
1PkGffT6bfjdGfSZbYr91YBahjBLtq30+ZK2C7P/5i8wi4l1dHkm8jxkVDWdGVXV
r2fOBn36HHZqnjV6lj66QMhSViVY2Zo8rcHTanQ9goG9Om2X9el0C+OuschaIXTq
RjRYO+0IuTANTplpvzZEPP5SgI3/6JXBkS/21fY9xZc+uwpmVwa2dC4FQKdMfwx5
OC6Vi+Bslc//RWrvYZvHPPmy38ddrZENohmr4h3DoUSBXAoawuyk0ZKd4WjF8sFH
cvpA7fb8woUS3B59uGlQq2ij0w3anIRzXPbYIBtrXtOhvlYwdkjGXpCcFe1s7khQ
5KM+RYnL2JHuWEh+ic38yBdwnoOh60LGOTZb6f1/JHPS8jF11LK0YsS2DpmSo6gc
HwSexBMSmFZEWBCx2aR7Esfbpuf/mLgpZUgiXaWAaxOeOAhH8gJqtFMkzM0x1OpX
Y1Wwugi4zwRPw7DkrfxvulKddSt8XbDUjvfPX4Umi5C+PSSqwJiAADfdS14u+VDc
pQeNIfGNmavDHGh16CxILKHSoe5LLPdARidQDg2Z74JgduXjM8HlK0FEZj2WewIH
PxKD95sMm48MFANoH6QrBFZeP/hMDo6FhK/rTmKGz8LuqMD3Wp27c3QBw8z9wQ2Q
m3Mf0F7vr5eJRrd03S+KCdl5efkeiHr+JxAe2hkeT/X6P5bInUVeH9vsZHWgTDQf
a/PMevR9Bolqka6k+gQxY8UZJfJUQcYeMVXC+lu10yPOxQ4+1VGeASoyZAlZ4nLp
m0s+1Vlca+nh2TwCRVqF0u7emosl22mkbMA7P98EdONe9lATjeS9dTMNJMfJz4xy
MuRrtZY1xZGvaxw+LP+evJrk/VpcRz97PFf5E6bKw4tLt7AMm/f/4Xh+jN+S+hfB
/SBccCh/qafJMcH4fi09X3rLXcfXlsrtdoZuRZZIIeQeLrUisJSrGV3bUTfy85i+
EoMYCorhqn75HUm9b0IO1lN7aShBcHCD4CO6k1GIR97CNBdYKIjJ1bbLd2FQx3ql
afzfxNiiUPR5teNZ4bJW2Idq8fwr9Ijt/Xdz/2hxJbaVHYoDGVLkpMkXjQkqXQIs
H6m4Nb+IrKcuPVSlDi4wmiXc2iePM4CLrcuekZ0LHBIxJdm9vqQjNTEyQ2iAgHwI
q5QjM7Sbv5lgC2vPNaLdxe/qxwid7PMZ04t5DlxOyKUzw8ku/sOa5bkSIHXGlkP2
X/QxVs/Wtv8vvBEOIJDquxK7M5vs0YZcziOBmT4eczmTwvCtkMHAlufrCxTcqE40
YS0l5sqn/sF0HUi2EhfDYmzw3x1S9ewNd8Ad2UzavOySYpjW11gXu5vcJ4DNeRQS
SAmEY5plEsDy8opBDD2m3mjcMlgr3lWHK9nVkxmEoejg5TMyDN97R3D24HpEoctG
NYCEs7pzEpvCJpnK6/fWtMovVHGaRFdtE4Nf5z79pJp8jeLUK8ZwKOVaDJ9cmgIt
8LuLr0PMUgJJ2YVa3zvChY7uRiGrOx8ofiCOZCc6aDp/qgJTZzV32/pDmpf97KoR
xGUETrqGt690WDWn4GsvsXJu05nbEOF1opo12s7yli1YCk7LC/A3pAdMdcHKJ7pE
uKRnXCVS2YKZzdJk+fdsomK40p6Xf1pBF4Qle8Jj3pP3B4rWq1NwHab8XU8aEbLn
JY9IWAPMNlY7/g+zvO3eNz4v8bLtLwfwt4ysL7EydRKOSybny/hbTSoEZ60cLREW
/jBWtwkCgTnc77NT0fI3a2WmmJZERrO+LuKOzxSzynnj8bY4ngGyslKzGqgnp+Da
hUC8fhIa4044Lr58lXxvC00AFC9L/wjxlILaeVkOShj5OREvupsLrsHYg5YDD6TV
3UOgky9AlnY0VLuCcVotJR/qQyZZen4pOFCzkok7NbNZK9N8KoER5m0mkOvlsbf1
8wGUJieCO5TYtCw2wB7BxGxfRWd27AAsYhl3jZVhUiRPWJFyde7yJPd/GuWWYo72
eI4Y/rgq9CjPCUSjQELm6qoW4AkKae53QgzbSxOTMO804sC6bGTvsrEonWmVaNhg
xutF+38UUtPK57jgWNqCO2PG1SGoVlU9thjiEJXRb4g3c0tNHBioMwCXjgxa4oa6
nSt8hYa17LwjBPPErj8B6dsYsQ9pYxDmYYGM8NrbXaTqpTAHoYKZFqF6ULp8Nc5T
jr5GzaWmqRpcDAnCd7YMT8yFgaY70cV3TEX3T05pIrqJLYuI552RIHS2JJ1i3/mk
m7FClWfW8Le9EglY8bwFWYFhdEsKCRZk5O8q1j0VMomLKxmE05A17ic5Mkzj/eKA
KgnWt7U6k9rMkFca3v+aA47VVpFSISuc1c8bOcHaKG6b/lqaCDAnQHBtJahL119R
ppYAKeO/2AgBjjRbVmFC9B4BkFD0+GjHpRxxykIOeHclN+UOyGQCEeRzkpgAWi5U
WL93FUrryfpK0B/9j064cUJXaC49G1vByKA4BSN1iakAl+50dJSxNDZkJP7E8gMm
JUU+ArNVvcBxhJriNpG5+T/G2w95Jm099q0UoO/jM3sp79spIZrCpbgjiixFoPA2
+c7Sgy15MK8aEbwKdPvKVYwh63D1Ih0ezKx3LBFMh0eDZD1GIC+Rjj6PBtDxLZeu
eHAqKBnvR7+i4ikY+L1/5MV4IDmZZyMR5KtsjW+KPAhlZ9fQ2Q0bLmIMDNwVV1aR
2RzLdszGpCNBI6lXpUT4m/eREdW4BBSdhCMURtEgvCibkDEjO9zvW3lrzcEA+Oq5
ScKFZZa3OzUog/OEi3mVDA4ka5Flfhr6mxo88wNaD+t3AilJ9yGmsv/XhA7pNspk
irz2xhGd/EKB39PFkeK4xS2VMbIMLikELRYP/JQFxuirP4tVta+9c4JtRHXr8xRl
efNB5u+onyqZQRoGmFdYTTjwbTIN+6ZnHwopz+X+HVHMLEGH4pG/Ww63iCHu/pNU
5w6mtyPD5NjKwD2w19/Fg6i+/TQxcWG1eTkB1g9iSBJVZQTvQBMnyuoCiua4t1E6
MdERNl+t2VFXPECWx6I+vVmcPPGQ79te1D+Jx5ADnd3jOlzbDUdkPYfnRHDzjRGB
jiotFB3yJYjX/f2Rht2lV3RiGeMuZaNGGYICX0SWjjE3J/32daPZQTuxKrM0mgGj
WbiOvM18mLuNP/qsrlz7KHqQzU544dxuktmGxcenaXC63jek041+M2uCkspv3P5q
NQ4nyxrdMoCOUYHXs9Bwgb8DD1rUfb6S/wfSEw3QdW9sUT/TIpc7oiAnLX393lU9
RsvjEzdM/W+CydoB93xDIFKO/VPlRV4y/RL34GLLR98VamU6cwfqvTUzikQnAfru
0DnH48TUB606+2F7+GjELDvbuk+ZqtSrC9ppJy7khnk0SYJTLXpB8zPoASGMlW/v
odEyPtkDkySaxYeriM0on6KG3zCegKj8W4ODyhx6DFoNCLdnyKvuJi95vozHRV0W
Ms8Intfv92Q70bZB0MbW/Fn68maqeRyEqDzsoRBfPNDKOIR0PvjVYj0ljN69MFK/
2+ESCaFdWC42SRql9dF9y6DKsSWSxYv5I0JimkCpGA+5ll4R1PFprB95tyIqCQ2C
ucOPxpuSNPZEe1hY9PJRPQ8LfRlcQ4Y2+U3q9MII4zZn84QgC/6Rqrrg31vXOadz
J/sZm+3xeY4OmqJJdcTR/6ChO5deXHhV8FabxvH4aV4OgMtUbR7lc/S5YKK/zc0a
mfKMjXBdt6NcRx9boI0zIpgjlKzzDwS8hqrXw1+8lZA9/CyWOB7jYlSHMnw/DyzI
pmaOUuCkJvxbTEYhcUhDx7Hbm4TazKrFQLpRRtnCpvhm0e1tzf00OQxPxjMRk+fs
tMo+KhFi8VyUPJnzXAVSi9v6RLOB6djEf+f0RTi7vBY8v4fxal/4ovwMd79kOwv2
yh1WgI5al1sQQjQQzL5czvqj1scyvTR6Vl6uijZVDHSFmrIXQhRmc0MGKLSBZO4s
0fr5h7GaNpR5N48GD/QGiasiknqsAsbGurm3tq2kGiTPb9T75RksmYztGjvRqtc0
244FNywW+VWUv/up6YhgpFPQ8BxqLCqU7sjdE3Ja2OPnPFSrO0NjBB/cEpIwzOFD
WsZxzCIZi8CxF+ypusaBF62u5nL1VIfycmX2Pi2NZ80hI5I+3eSh0Qg8dAz+MlZb
rB2jPzIzDe2Yb5WOvGkFvf9zFVgzPLLy9ahKBVxrMQCcdV7A1OsEW7jkoLgOjZXq
PFwlnkGrMW6MkKM7KSrcj9Qql92RX08kuvAUfG3q1PEiiPXgyzDeBAEGvWuZsTpB
uG2W5pgg2iXTCkyXfoxYWbGMKKZM/GK5olVj0xUIoj6Ix2dUUJ5as4c+lKYOUMV5
K9AVn5JVF8wemYV5hLCWVmOc9C/33yjgJugPztTAbpDesrgAXUIANKOggRQTxe+X
2OG6seVIOH2YnGVFJSh5Avb8zYDQDesoH0IwWLUsSi2QVLmgrU90GB2DcHd39js1
sWLZcL5zQ1gNZJSBUzRG+gR5+XxyxugWD3ZSt4zGVo/oaI2yKFP+y6K/nW2G05tP
8lOu73yN1vdb1SD9Zyc2k36v1PaUY0mpdWCYMUY+KUTz9s26uK14t3pkljUpTeo+
AYoqm3NGMB8yRQTXEUGAaF09PoMOJxekQYfsmEEeMssOMR4tXHHDnz7bHPp8+6Ps
4FLV2oW6fSL1U8iYDzJOnFvBZyfqcOm6ZEojU4/AcgzqaOxKmDGWLgqYOV1j7IPj
ri5c0MG0pq9O+ZdfhXPrLYSRQusN//ESeZzrZaDVKvKy/hwneH9zqHIKxI4sNS1+
/+sH4PVvElKA4D+6nV8IqeNfjjKKYVsSoiv+1PwTFXDYizPT8n8/t3EIuVSuIrdq
DgU4Tb/waI+Ysi4H1L45oVkDPCXl9/4A+tUTwy8ZzO5TWOd3mtYR6PK6da/DJeKe
domif6XaFghq61G0sZesm6mg7oNFuK29ihZcOaPmWykhthd9Ea9efmv8CTjYi0a7
EXcVU+x6FFA+KPhuKfDcairtyjUYDsXhLKVmYKuW7ENtNuNpUskOwWB0p+Kwi2LE
LSAgcp916EyfU3r8GH8CrbqrbAebXDiBh8ex0ZPj3EaklJC0dUbr7W96lx/nFx0Q
WQID8bKhXN/LX+F2ka8aCMqP1v95fcQu7dfR9qIcERrTSViNKGHAiTRy0iGE20Zv
696LdfdzVRJNvPUjO985s46CXvzGZ4aWGum8S5imdMnJZyGGoNwZdxBMtKcuqhpN
883+1zi0JbtJmde85D/7XJWS+I/6OXBBtiDrXCO6SYW/A/gil3EBq3hwV/zdJyM3
OdaKJIlZ46NphuZVgc4NIYh7B4X0cGU7Kosikjeh/zv2dusU8DYKsh6AgcnFUuXl
1itpw95URCyxV8VUQs0TwFo+IHth48m6F9WcjNdO6ZToHDQs0ehvEUdVFA0QsL5L
HH7r+aep3psmPeBui9zL9/lrxeGDqjaJ52gKLntuhRFt1AFMbA5Zcp/OyS5Nhi35
1yJ/0USBwEhiqhS/Fy5KRtgHExd2nhI1AjcubzuFo+503hQZhJgsWzKSnpSc7BvD
gjdOhc//XzfD//vZ6mEMBg0OqEbCgDFuOBKh+aOqMsPUNazcmFl1JktUxKBYyp8l
Gi6FUyXK/kLVGjf80KLS6gS+a8lEp0y9kYgGa8CwBR3urXu5AuSPGQmFUkVl+A5y
PrSH2A0X+5SrJa8nF3voWqJKMJQprTBokpursB1a5NV39wNEZoKRVwI/FpRT2/GP
QS26/TESZMW82zP13w/cCAL9ca2pYVWz2xGE2lnU2mNRE6hCqSlxrrQxTkbicauX
7KtbZ+aOx5GTvxV7D1n9tanxfp/yTgxcgpZCT7MEl2ELwjoBk34Bm7opSSPOik6g
ONkjebsUy3nWqRBrJO55tlMq60PppVhdi+CsM46p7oOKNoORNoYZtX0Y6Et/TyxI
boGoln1VthDm8qMxeZV4DwA/Ss5pgMKsm9tNx5uQwxYe7HLhdvUGsqt14EiS9jHl
ERgVZFRPb0gTv02d9//eVmHjtHurW8+p27bbz3cW3Q28mgtSKpgs75qla5kjiRuc
xJFYG19LpKN9YxNSuDhrEvJHxcxgAZRWtDt/twexgJhsmWApMRX9E2ANL8x+Lomf
mFTrX74IUfwHguQFdqSo6cb8LWCG8V5V5hoOf9yTtGOUtrmr6095F9kQTewVVOk1
b7WxtttOwIY9p/0FSXRk6TyMMpNikBr/R8dizhEwYGjswT/2ABsC6dhIb4Y8QU3w
SjRvfeIvhL8m1cv6QkrqL+Z6aYJ8y/zJ3JyfowlTiTGByAJVBXDfqQZRpC9Lk+y+
p6oPmjahi0Nnksfyh7ozje/5HdTiUeHTWVwoWb+680IhNey4MNFfxCQLE4igegdc
Y4xjlUI2GRdv4v22GFop/Hpl8mJU83sF6ZPUwhutg8Ogmdrl45amK4BGJGeYITsF
ZFtU3xVNezVxRUXM1ACr+4W4WZsqjFqPc9DAxqn44ja0FmwOOQbYw/x6/ymjpRV8
kGSvA+hlnW9Qv95nPU7w/7OpCdUvmLb3nuTaBc8111ECTvffEAiYwJhtO3ZLda2H
wjYReiMuPbYx4zlje3MDx6TibaFRuElOkrs/Ljx1VP9Q/3I77w5LrtEmgeOLGkq7
KbLmoplo/FAgRhv5QEh7DcaTiLna0rZfizW3nm00xK2GeI9s4Sq1EA3PMteKeKSn
MsYiRQ3GZkxnLQlusjUJwH+eRmvXHZCdjdRQfkz34kr7ZWTUWw9lwRWWvat99MOd
mpRgq0q9CAFHPrJeORCE9dl7zQ+g8+7m7BCFGVtGkqkUy5N9VHd3ddwgo1CT4/B3
tgbCsdpfitSX+F1uDd7zQQ5PEbira3uWkOmtnLRLpgZEvrFUZwCbMm9nQlwLcl/O
zlBznXCnY462tLJFf98HGNb4GFm0bzFsJkvT0mSRrAq5tRqAX6xVgVGifarkYWtQ
H1DPhFHNe7iHzOftudYV8CFrUlaHuCfgotiUnrABFe++MH8CwsZxvkaYZtpzuUzW
6w8uUe3ai75G7/6E8Rvj8ZJHBxoqJIcg7HGHqWfgHj5BOTNoM2yTg9Fpc7wKGA9J
k8mRnZHKRwk5Pzy0PJ0BRCWDi3aAJtwaIpbUPTcGjZyUGxdGHEFVbq0t1CZgHnP9
YxpgvjSmrFh4gefdu7b/vIoPvp+9FtipOKYXoKgeT7qybjucQE3T/lJtOWWwd3zy
cu1EleWDE4eD7ylWIL6o3qcvYoDnRlrKHbCGKkWK3WmS323o/z95Y4qvHbJtf7RW
vubq3VYRpXw2nE1oeojLZzoqEozpY2GFYCoDB3bSBPL8r2J8bBY/EfE3ihQ6u5jm
xmYEeLjaMvuGhHN19NM3UPp6XVnzOmlg/PTRUBBhBtBjykPlY0NkyPNJtK3vg71a
s9KYYytbZBYUy/HtNXVhbkKnXuMNcg89HM0gJMNahIHsu7gCvoPFwzpK1yLN/lU+
nsrSo9JTttt+MScUDkd5H6wyAJD1gLfX6bHox6nW5o9XK/KyoCdg/fCzY756JYLr
r0Xqb6IJTCI/XAWrrExAKhTj6YU9vzFFRSqHCR45Ywdh9sZVtJuTlDjPx94djgOM
kKiLAuvWJXt6WQXKkNCC2SyjLN7bEu1XP6kIZvG4HVpFlIAI3lMMwUG7I4ZO7j67
zA+o1yWcRdFnWW/KeeYTx4pBvzKv8YlT3W5fMQQfzEHfZvKOHOVaI3UnN0TkNnZi
2j7Jr1fphFzV6WWv95asLwlkDWtV0hwJ3zWtNr+sp6+XvxyehRUZT6TKhM4PkALM
KU3TzQH6zSrgP1Me9OOkvI/Kmi+D3R23hO8DUUeIh5FvEu9qQbepdug3VPgg2Tbw
TdFnbNL4DBSCboCVusK2O3DBcdBBhg5S10yM42pCN2Zx4ZMWbInV2nGwbbt5h3tZ
twWeibUJwKmD/h0KSbztQILV2T46t0S1V16lGG7xYlSGCXNm6slLtyPd91ZWNCcA
Pfy6b8POyYzd6hdCW3EXp8aXSrUpL/L5SbdvJEbCi8Fgqc1f4S5zaC4reflaozEw
gFXFFDhJynX19TjVzazJi+tnvIE6XtiZeF00JuFbeGXTWOBZztVeRcdYOyoOxhVl
QVW+5n9T8Gvybc+QlYu0NB+8CZlPwSP5+lIHbtPO6IebyALuDU2smP6JgT4B8Zgu
H/176vQGSYW684VyrwnjlgutWTzA1xTHneKaHPmYdrU1p7G6wJgwKaqUyGiop9o6
BBR7evE/lTyLh9UHtqbrvwAZJ92tK6aSSFsec1gr2mS3x5pSBfT9/SHcRSNPID0I
q3PoxbXQPgGvcDZ1ua/pQSdRJzUbg6im67ARELQ5eWQbF4matWm3tA6uq/f+4L3V
R6d1x/Jl/QOjbe+SW1DFKGpO3D5ISsqVFJ6NNWa6NdGg0C2v2rZIdU8y6KVulF2D
TkBrRVw5vfMOlNAtyGeAyh84ds6eGVrLy6fxnAFq/R1N98lk96t4Wvq7C5HvIYM9
U24voDpuaQBE9ByH7f1k/Je/9jJb/V8Kapo0gmPtvUKSUbcdJqEyuAj4pHjy6Gl1
q+K76hkthIbyCNxsA9rlDDg+GSeJlxgRocL4auubTuuEkIO/6OYi1n/wwojJzQ+D
g0uq9F8/6VTu6rCeNV3ntTiTHzDWojCnx/BflL3ZMioiCz9JgdipTfL0FjH1dGMr
vvhFpJinBpVJEmfD4LBsO9XNuyW4ZwDKXQ2a1tx5qiz5TS4yVyZMS/G/6aYcMDOd
09Ped/4klMmmL9q3i3GY+PJQ6jhvkthQoYW1kjklTxyci4ZvLfR0tCkRHKdgws23
h0fL6di1N7ySIjIMP1dGb0JrzmQiTy1Ppnxe84Gxg7dy+/vYvtYO+SwJHPd9e4TG
rwrUlNo1iHWGF2d5CtLcdsfygCSjehT/gFuoIw2EPu4POglyJuP9wfBnswi8Hshb
95b6+OX+BAXbOeZsZaoOft+uIuH/ycUzUIKkZ+UIyKM0lJlPsdeQL7LzZtVvkphf
8BS7OpJWZHmIwUITbdAmn41xR0hyUH2LpI7t146vXMuqOA9RXeRxA4hD3fFt73as
7vKYlJ4085RmQpDD/ZELVncYXLn3fwmsidLTPriaJtwft58JaAPLdm3RJe3P58WV
vMht5Qh5q+sXIOzymMYye28HDlI8+RCeoeerJPpy7iQ0pfmfHHKgQJuajhVtoiOt
7hZJ3A793+DrfSz8Esx+5kqdnGifYXCwu4uYhNmN3dvOs9FMnNjj3HvVpNKqTFmV
Kwleo3Nb4LH+XCc98AozHG0MnoWYmVoF0AS5+Ap3BEzY/PyD08wWeYR99hBlZXJl
EkiYsqIsGsvPeX44+kNLENkusWR6eigBDuOlVcHYcwh1u/94nu34q1uyme6azJB9
kgkEcsJon375oFhpyp3gp+QOLCSGd6ihUH6EZp9CozDsCkckX+DVU3guhUIbTqzF
a+USsnLUrPYQM+yOrs7fctvGnRCNumsroN+IUPOW7ngCz9LY5DWI9LtadCPcKn0s
7JJCQ4QRTHCOevOoXk49kQCuOkjzZBgSX3h7pCIyRFW2Jw+F6TdWuuCTECrfztKc
m6lliD9fAsBtQ2siyhfP36IAS6u9c86uWB0jl5KZ708x5vJPlJIXFfURic9z99i1
GKqt0vqragc1gjMdBDTG3zrC8SfXcFlqX4/bZD0C6nq1qVhQx8hXFRFM+EJ3z/pb
79ZS+QeMjhs1z0u+n4gX+A==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FIG2CExSgi20ER1EiVud7cbtpdfpqrtcGSSIyp2tg7kodOJG0OcQZ1uLLUbXGaIg
2DesTQ7DEu4YO98wbUVCFcCxBpIi0F7Rs4tF1fCML0nED0qo+eu3g655Za+QUJ34
M+D5dpx5D6aYXMLWDWaIo8tD6XuDeX7ZIMNdrRhLhuhrX6OS6RSm91VJYTTfnqP+
RfFSsqfPpzLqDX1omRQ1+3/6chD3v4gtLz3UbXivbjBJpqkz07vwn1iOBlvgpLDU
qqFNAUSzGSuLUxL10/GLAVFGdee+iYXY+zCt1IoHaBd/3BDfgeo5rcYKoDiUS0Iu
ICEt+nICtnLRVjwP+dg6nA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 27200 )
`pragma protect data_block
6szt1kZp5/ZN1olqfXz8+19cPgcWoLKNsq8MV0HrAdnLSRC6NHIiRt7uI4GqVJjQ
L97JzfM+azjXvkt9PBo0cqtm7D1S7nm8/RkJNQBSgSgt0Lq0RnalQ349HUJh2GJB
nQgSbJPOtvD+sB+Sckp3fLHli9BDBzEXnemiZKbr8md0hR4EuJ4I5eYzaXyZnHUq
bs3LSbEFBabzQvHpjagavOvQ/vlB11fLHXtCe4izS8QoXmhdA808RcIVB1BtVuMn
h9xaCyuuszKTGKkkxURSMiycAuTNfGLXvY0wylWgPxq/0qIKZ3HlvL0ANqiHUT1P
RSCSBPoF/GjFlVvl2Fg9yN6wVNo75p7bZMkEP0IIdMD1OIkOPoJovzOJMlA/yIFR
59u7ZJDDpVMWZWJQEEhso72PyuTBrWv9tmoP6MHJ19tjsxF6u8TKMArOq1BEnfVJ
yvSINrtIi2hfrwOGfMkHXOqn7UVTFWujahmxVBB4I9PtskpRNFUzN8gZ72tcdRmZ
S6rezc42BThUXPIGF/6eLUDMhxAylG1zZpzDlwqBjPvKt8abvTf74rr0XgiMbq7Z
nz+EgBU66qBtj7H6a6OCkThSHPqHejRO+TlLo29Jh75n5XhV0a2WuRaeflZMFsgV
Fodjeh4ouEHvB1h4eFZH5GvaB1OACDqiSuhv4tu5/pUUCD3F1fh7vyjfa9FBjOua
OKKEwbRLcMS7aIh0gN4hMzLGH56FP6Ipy0XYWcpDZzRvopf7vTwA52sh4NvgIeKy
itJ2FnXIXqzfkdONFMQH4EC4hNKN8n7fVvj8WTGfnV5Mo+vTWif3ye5nXLV36qhc
9Xe2vzE1EnHwaZBZrGVfhVqMSbvGxstA8EX9nvnMn+URhbXuYDPGMPrLL/ewSTKH
AlRqwO0CvCueQLjw3WWk9HE2KukFYlx4J3FeYCWsAtObZ6InNj+4A/x9JLWOqthp
iZ1eeDeg84Nh5VNR077DA0lZSFSyvDpDP8MoMK2MwfUD4+ZxlUitISgWdP+SgJ0H
4VkwE6kjJxJgMkBSY9pUoRDsv6Xnj9e+eURjQ/upM3QXrHkqKruEIGCaPIz7WnQ8
BOd5RPTCpP4mGl2pVk3CwNxg/Fof4g60qnupI0+FuAerSWBIPVJqNbE2APMmCoa7
Z3BqIc17AFXDzJokADvDMygfqw0ve69HmbEWF0KGsIhgtVwy51lFRSm2Ag6WYIsV
MfVRzj5jERPebQs4cqdm/gJr3Jn92dYeQ5X5oSRtXl8/yAWhBxcyTYw/tIPcuJE0
jt/uEm3FUKpIS0TJzsWZMeB9nZ7OmvHvazSp5jEjatsq4i5aOFZnF0YuCmJ+kJU9
mHqoZ0LlkvW5OVjZBs413yOAzeRKKWlqze7Nsho50gok86D5b60d3u26Gfbbti/z
8SGuM8DWA/XDP1cIGGrILca+2FW7Uv98+cvY5ojuWWF3qnpHDFdEzUxD8NrFSkfh
Vc/yB7/uyS5ZjDPie5J/EFBjCpNSQn8jAKhOBNWq6cNjxONMJrYru14GxrUNyCzG
bWQA7B9o9WWhOyJu+iN2lLpDH2nHo3CubcomT4cyd8aUkCz3genFsqErpzU07V7L
FsWuHurjiY4gSMwi/2bV2Tc8gQpDK5rXsuZ0RD2mCf3Z22BiSPOcoLtzpvCQ0Tpb
4+NhIC3a78E606llI1FzUTEpzWiXW+idDCHOEryQowBf35qKvReVQ2VVe7FHdRve
ix40mDDsEqOMDAjOSkw7cUdsxtYgUTqZ7n79q155Wyd/bOYGA9xv8cwVgSdysrlT
kuTHgHWz4sP5JCbeaMjlCK5csk1kJtlGduTjfJiLqGcwAtdXrbyWHc3zW40cBC2U
Y86e4oBjT/TIe2AhW4sYF9BZI8j59y1GrEwsIzyaT+JUKwA2NZ5LH3nssSRqAsBw
rgYdXsu9MpPXnbbuqqwbrWENxmyRr5Onb2W+Pq/hPflQa0YVJ7H3VzBCJWeM1z2b
Ww/nHw7AF585HOux+43hJBBZ9EZPpraDOT1+2qebY4/aHGt8fiZbmXREOAEQHBEE
4frnveyjHfp8eGrThJwQwRB7ohjNCVPROLccPK9hgF88rm+2aRrGBcydq8kgGNsc
ewK7cOI0l+DMVTT0AtRgByMQ8CKO2vcwAT67Dlw/26w66bMs42ujRQnzf06wH8We
6oCBE45IVZsHz48gawn0HMb5fXrBFbGWvrgKaDIVQGDqTmy+imkz4zExknDPJwHw
GLg3K1OCXCoTo3NIWlL8U/c0GKI2pJEt82glWscCYfrA4zkrx+INWk6bGtJIPyzG
iyd3jyH3XgZF2D74xceUrU/MfBO2Dw2P3UE8ZQhHvpnokCPbkxcX+ZRHYMZcIbI+
iRGnVYXNrSukG2nM4EIgc2HZR8F6iOmLJ/LinVZ6cDcZu7HUPgzmh+4E/6NUs5ar
5ndshSC5hZsBq0vY3dl+h1esr4luW/0LwTNRczyqjm/NhUzqKCoQ4bXgrwXgrLRS
tLAyCgNpz8LyY2hqkcDkRM+QsJoE5T2c8rEAkunpt59XLzADr4/aP9HMvvz+7Z6Q
v+S02F39eQ6yx+btbQ5w8KoWqaGn5jkyQbvMLc7I2+eW8qtzBNZzPpwdHtrMIUQi
yb27XEzYOcxZyLTyYRYCOmvWKSZ+qOCn9jkhpzUjrL3WJpLpLHNH1u0pW3ieRPYN
wgeuZC/TlJ8nqRDKiJZW4+ElXXGx2wDdwKEI1Rl6ya+x1gQyuy+FhSYdaTArqPxc
hX6qcEiCNC+MHevDmFIc3rmuJgvtLlUYPLjQMhUrcYAwD8jDZbZOYEXYKa7/0DIc
ldwx8bvu7UyfTl1KTiyXabyAtuTm2U+qE1DeLqWNt9lUOWLMpnMUJYLt6iMCXOyA
bDP3nlete63306Kiq8E80NVDpz8nLFTlz5Vjofe6D2s1E9GSl7fdWOPl0iB7f8fT
jCcFfpBCulOf1P3EzzyTNnNotLXG5/uDT5fLXQvFaAfmfMDq6pUl9DB3X63fmHYn
ab67uNWGBEX+OTqnYjQo3SZ9Ty7dQDGzdswjWLNpDh0fbZEtdDQjY/issunoM2ld
zxq+OBl7QjoTfb1a4UKl1diBhMoTMf1oLfBh6h9XTjM5YAFxRZY/U1Jm74pT8AnM
Oi8f8NIXwKy1Vkuv0JC1Vk3XEfmDLgD5maZ6OmVcgab+a9QY9eRBeYO0X/VK8vGx
peTckuuqiogE/+lCJIZTcqoD8fhMiXkxNvK6yAMpCVoyVzAR9ABf866OUU1lb6RV
Jh+dqBd8fDwb0LZIDOpoIEM58rLdo7/g0ovz0NRxUT62IKSJbnPHHnQursk1hZKl
qpZCON71C/hhw6I/qzWQYndKpyKIQFPVQCSOqEVc08GU220JMWBSPmMU+hf2vdJm
nRg6uOYQ15JDC4Ag+TEnOwU65sDgvsz6d5fyvc+Jg/2HeI6fQjXemAaHmAm6jq7S
61EbPNfirzdHIDGPmnG9NcTDIZ50GVHDWfeoBuRiCrkN2lHvNDM2w8KI5Tkms27V
Q4IjFLvCLo9O7QztkMXPr8gPfw9j8f6QMJiC2itpxaQtdbnVUDyeEoPHkBefGEhb
uWdZzkFGOMEQbLPLRq/wGeIFpr7CDopvrjAQu4I/r2LyN/HqIid20lpOH6t/Yf5L
Xk7vgkYiDVT3wVEjc7SCAZm/U3n46rUwBXQZRqY5LPQO7sTQl0dnw3S8st36+PZJ
v6sEJ39IspDtOr2jxOUEjNz+E26WBuaCrx+6aKPn3fHG3bUN90Ev8j4H/jCcpaTe
WDVKB4syo8pNSXV6PQaweO+YG4WMrg9GmrBVuizMNoJrASPhjEijPDZCHZRFfOIw
yu6JR7uMLvpAvLuH5SV8MHmJW8KLatCewc1y2lgatNRisQW4Q1DSIvaAh3dGZPg8
CilKFlr37zOW7jtQKaPnLtWH9NlVl3JEPF7IPGeQ3RpyKQKJCw3Iv6fjjCpgM/UX
/8xJ5v3TtIvsaIRPqrazBBBfpS8rtU4m3pvPXBXd9vaZxjCDjjsNGIPaFMRJbOCe
e4xjWxN902h0fI5BuIAttAlCfHLlcXcQnE6f4Z1fokwEXhqiKVl91sV7y0QvOabO
LSD+XLLuopsOlMcgcIcrPQ7R1OrXL0q893Jja1ROCUwdzYaal5qWnvZniOHYzBvQ
pstIprb1UTK0vSfmU+jqls+cUZq8K1sQF1O3c1saIClhoB6WyUrNdAJAz9eFKvgq
x68+jv92mjMdTwEPU0EOpfYGQU03gT/8BQ2SHnYFL3+mRSqF7S3/h2RvWxuRePaG
iEbllaDA+q4DnEvTRLOjK5Te7JySXuTPQnUWNCWXnawM270tATap7p8DdYNcjjvh
eoj7n+XSLp8tpY07+NelCiTrjpROGzBB7s3yIaUGJEy/X3KvFG5IzbzY8wfNl1vH
yYrYOrRAS7cz6byvVeac0XorTCeMzXc4Iag2/+ys/In4P5N/IjfhfWq+lDW3+hLH
VuDweu+5elWmtKyUavsCG+/ab1jEMJGDXwFvJKgmlUTh3iVtcgnek8OZAbXFCnPh
lRIUWRUtxGkPmzjoEgl7nORbHHdX952CVoVn7qlHUV8XpAJYj9BTFcahTUy+lBQW
ftYHCEafeYLezmVPt/FjAs5tJD8vOsXCTgEv+N8oGAVvMAGBQ7SM2v/vjMuBu80C
RlsfUbkFf6hzd93bfSMBbnoRhOWjX3TiVba4iBAGB/s30ihbsrJK18RrNUzwm35f
2uJKEIr+Ns18D1FGG9RngPVOOgf2LTSsFIxycNnUKs+7AO7J0S68ZxpitGjJ/hQ7
mFeXibjAnu8y/691JoVgenBfaw/uIpr7JN3udA1KBSm01H+GKv2yY4D+tWBxQMIM
ZJ7s+QTvxelSgUi2O22+eUVfNZ9PG5r5+WZrywMb8zpqNOQ7fvSWP4ntpHE30roc
Q2W8UHSWxwQFSyo04ssar6izoS40k1tKnwmxzvYhP4XLQdlSkrFVDjS0Ykw9wC/F
hzqcelCR8seBdddXWo1gm4KZszMUh0tQOntwZjMM6qi7c9Cq8oTscNV62A01FvZL
qMtC+yxpSrpaMwnSfN0m0OO6+RawR53s0bR/z6fd6wwQlDg2XvCQ+MfzrqRKOdzg
53zJb39stVtBJuUenx/IohXEbvPeK/MBQvdDCls/5BP/6i7tJFJYW1T6zI/gDn9a
NOjKl9ydGGMyH1q/n+A6gnXe4W2C5wupWpiMjA9zAJh4BSpNpawIzGPiMjubuIJ5
lr/YV3jWbiHaKX6ODFw12M8H8FvsygwcaK/yNNA1rSAQNwEUfOX4DbtSvIfT96Cj
45gLzPDxBdvGU4Ksp7SpjKtUx5uDzkxdk+msHmvpgUz3Hbl0jgzxF8XJtBdM3w9X
Gx6k67jB6xhSF4vj56m70LpKXz60+4397ZavBIqd60+vHj0NB58cRR3ywfKhIJXa
Z93iwytGPhZ7QHwoZ3tB+suGENJruNHiAqMJJaiEiNRKFaS3Y3wIOS/shD1mFcEO
Qq0c4TckTRIrkjd2Ox8JjfvaO7h7/wSIbYVMALArlM07Du9M6m5sVPNrz8pnjdsw
7sdIFmQ4NJVHjjsPcmfZ6wryl+plTjgq3k5O1H9hRNIbAq1E9834453ns8n2aZIw
zho2QwfYzftpM5WD3qJrKol540xr8MZIWCPHNe9YG+rb9wr3CUEyolhTEiVYxN/e
vpMuoYsZAzRXif5/FETpONEkRgm0zxDlfW8TR603m9B26NZMMB+uxGduq9pA2I0a
5DK9G/WbYHjL+uidOrzpBR7pVn5MIPCIf9YwUYWyrnMJXgGQJSVPUec3qNdHqOUs
1+dw2FT5BhACLJjUQqR5w29lA+qp2M87s/4flCuVoaSy8TiohUqOF1n+PjT2FmQ7
JYooE0gjLfJk89ReyAs0StCtGD2rYRNMOqq9LljFnFO8lfRPVIZKwBhdxSusmy2y
flFgwjggPhTXKCqHRNlqsmN/TxrR6gZDkCqDBLZp4aTaB3Nb5PmyKcXHI0XtK2hJ
vzmArDRxsykzVx8s1kDuZhnRTNLhGVh8kmJ0AtHDAZJEYl8KF/ZRDa+JvQOZazKs
xROLhy+hfRWL+iWAz1PZWwwOucEeyCAR56pL3Zh0IQ/xzYQpHBUFzXX7p8A/DHa/
1INe2YdB+DX3vpKcXMjpsUun+9W+qR3N6bJvWK+f7D1sD2z+99wqPTwF4kFlfhbU
/myz5qLKDgmWJ35QlvQW0Wt8M12CoiIpbGxbRqn+6WeaCGbylpgmxdR+XYVXTbln
aEAUiiwL7qrCqryaxclKCj51Tq2vZL0IAeWtKXQmxjHTCurX+FXSB8Bc2+kYSzcs
/Z9zfb5tD0okhz6bmKJMzaHkPzig2V/SUjIEAlZuoC2uC+TJ31ArMLKEQGvmqfoe
lgopqN7eXBphjJ3AJfk4kMgBH3grljk9byLM1yC4YkO00kcHVy6uGjG/q3kUdfgD
JE5zKM2gbX4HOPWqoy1v1pM5zO1LjyCLZxyLTTsnvDJr2OCA43mT7C99rNSNNCTy
V2dII0YzZwYmDrA+1NiWRI6ztt0cIR175COr24RvfW/upWu4l06xg8kdD9M57eOA
7oeaw3AZ9XvE81Ic3pt/fHpITx3BKKSEpAxw3Y3phCWfslTclNXx0su2f77vxapS
J4TGNW4Kadur2bB2EFdszCdhVIGQLjyLkYiB0UhZH2ctMC2D35hFimMzVlEXKblF
2SfpPTrSyBo8yIl+vLYbyWWiyYB4dPYstpzuErFVIb9b/4uLjI1WmBh06KIhfJhV
L/d3T0HENEdVEHBQ668N1jpiZAXmVBIA6PR6HtKpG73ksrZgvvLCAGl+dDjltI5S
3ACvtk/57F14A++fRhVQ11enJIAWUA5yXNrNbNdazqpX6RYQ4KeREK1f1w9tXl2Q
yBkypni7CF8LagsdOgfM1KQ6hTjDlEVF/taUrKkayMD4mxEnOQj3tHNF1HXuo/ag
DImgCK8KArJd3e0Wtee7TLimQ0Tnlx7dLjfbyLWE2Qi+RiTRHghXZJW8EUbGcIvQ
ERbBO4Vnk2WjxS29TMlCZZ90qDPRkhYg5qUwwPEyw8/ZqSR3v0wLjxssLlq7Pu9M
G/EvX/NBCKeg0s4lUgv1RPyXxdyrqMCwgrTMrPBm4tqlkVmIIkihNCGkCU55C7xO
n3SZPTOGSsnbz08KMCoIn//cdKQiHNutip91IwY2+i/jNtQwspiFh5VE/Gs+b3fZ
t/TntmqpvVsMzT1zGbs5+dX5BdXCCGsR2pU0O4pVNSF78vPBluAZg21maCdg7DYH
5Vy8gDd4aKbYH7b0aXfIuoVnsXvvy9yX7a7YY2WqMhmKNNV5mV1fw+AxZBhRz+/L
XntNUEawdO2FlP9XPIZlO5+Y0hQY+a+1zYLHzAzC2O5rrvKO2kKv3Vqe280ig84Y
4NrbyHuNptR3vyHhUguFJ9vSOH2CZN3RkiP23HA4wQ5jpZxR5lF/+54VbcZ1ABxN
Q7iLKM2lX6eHhjnCOZEOOCx7OfmO7cSSsSvQa1oIj7N4uXwCXTtabxGELzA1cexM
fHEEoZiLp8aW4TMvOwT30c2vps4cPSI0cdRHl4EhdZHiYk7J0M2MzX/JwUewNyu9
fSSxl47DiliIzCnb3x718wSqgalLXr+pLFoLdCaMMV7U8o00AGCXqxFGytxq7IHL
o3E6KfmAf/a1Yk9VZBO4fx2EO3AUgQJCGJs+IHt1Kwb5DucdRp3k17L//EIt8L3o
LM6Z9KzeGeu1UOaZ+dzVAw9ed0rulJX5hx2cmGvscyKNqbKglLYYL32eIGiocHyN
M+u1oPnaxeh6D3fC7sOJeBh4Bqkmt3Vicp+MCQGXn/dogP/L5i2W21nldTr69Ckv
Ktrbq35zX0Sh9WdeCMGkd8yDEu7fZZZUeyER8U5cdn3QgDUpnTIgvqfXaccBPFdZ
RulLw/csdSswJcgJh7gMYJmNngGnUFhfWgHpEZt8FFOQcfTMg8+Dqj/QP0vXeghW
srTn+D1ceGx6NJ9JnlWymzjsj0MF4TDK2KLsPAHgAiksZjOnpxGeg2nFD01ieOhL
hRn3X+QeL/N6R2Cm+WT34jWr7SHb7pzv4ZZYUnvClHCKLa+ZFQCY6dWsRvDJCe1S
9z+Wyex4e6uQ6Aq1c6o3+x39/moq/O445awxwYSqFLWsjTMkb1ga87Ho6RsnhI/H
i2YU6c1/sGWTnIFPs6f2pRpwz4lMWCQGnPI4gAt12/tsm6PzsXLwwHKlvt1PWklX
6iraZWFQ1q+Vlt132EPRFIWKr+Bpv6ojtGYv1UStgliCWjhkxrA9wjtad33ww6ml
E+0zuENPd+7IQR0Inz4xftUpCYUVudimv4KDgleKU2F7Dnla83oI6sOIZJjwcjQV
QJRMgjdhp8aB7qP1qzLWmfnS1FXRM7p5eteN6MH6vO1Sjx97XuF8Dj1b5V6tSG/J
lmPg5wnpwKK9KX/k4dTJVpMPMVHXXJOxn0803QpHjlzMWHIlGcVLaJb65S7IzsgS
bGzpJFP6VglW/o+ysIRwJya97XtTCryxZUqPXsqgh2o/ZmKqrFNn3cutaRsCL5Im
ei1KIRpCDZX/Y4K5TrEpkbIG78ruj97uWqHR7RAod0uYGTK2K74yaLvQEx+y4Ool
4rQyOO8RF81ne/tzi3EyLHgCo9D9ibh9v91ATwwvjbeS/MWTEGs8pfXFStthdiKF
Qrxngm/vTlfsoVDAcPyP83pI5WvIgOLdg/iwtik3aDdUicjbTgeUaUdKnWJG/A/S
cfAXaYP+SnB9JR0AmHrx/FlhSA6P0+c0CVJf8EEgxiZPZ2ta6/fEM5TGJ/NfR7mD
0Tq5Hv4MC6hIQhHO545FIXthnlLAlgO0TQFgpL6CD+ea9a4CZ1uyDAo5yXxQIyZv
rgocRerA7giM2OoDOSNy9US/Wa+paG1ne9Mpss+d0wdBJb3uHo6I6GuLWXiRdUMK
8D495/73EuLaOTY6q8GCBEdfWV69igIp1GrRO7mdMoMcIAS/gjpoamDXqd65n1O9
5tL5ThixvZi/nawyre7g8QS8J69xPcU1W6LFZs6317vvFOxMdLvhOquU02hHWERs
8KA6K8BJ6lL48ifK5VludGPjcMKPnqgY5AH7Uko++KfoYmcdrwCh7GA7RPfA09XQ
+GEZc3rTGKeXHTTNkYWJkbEmOSdjBEJHcDXhCl3RV7AL9HpNwyL3f/IlNQD8Uavs
hePDxGatKXz2O6JSsOqaQwXheSFIm0wQHipc113e6W6SXzFpqRbtMYBxTyTqXiKN
zuheBeG9gvENUXo6aA4ns9FOE4Q/SHKWa3ndfTimIyCoRNep+pYKVN8JsfLHehUQ
ONrap09FKKgFi4eOaU7vk1Jp2OxyPIW/WDfQGmH8uCV3zFqX66DonqtrRgQwL7ab
T2g+5tae/1IIUUnAEu1l+olbWiOib6ej0HZV0Jfrmd7/4HwFOmloHMHJn0HwH0jU
i0BclBTiwaUpGreIp/CtuocCl6oh05VVlYLMSu0WdvcPczDH+8BHMK0ajvpNQxKt
3SH0FDfa6mpReis8nsJ5+eSL1hK6UUtGOwS5zbw+dkOZrhgZ4/og3ZBbM8/Zt3j1
0CjWbELgIwNyvfoRxhxbCIIh8Q9syXlcJUeiMhy+bAzGZvEVQWVkzQ+4elFINQ6N
Y7KOzPnDr31VXTKCkD7TTdcO2O3rqDsm7lEKRgzgzSCeUA1bqCfb/WqH2Ody3OzC
B4RepZ/qElQhKAwvrU+DPDmJwAAVLhYjiYhSoNuo7DGDyXLZ5YoTq88YWf746eUm
RXNE+SZW1npyc+INDCBETfKzygbK+Q0nfSm+/2Yvle+/6jMy8a3WC7YWtXx3YTeT
m3ta7KMPvXWkJ5CqaSnY7g+FydhJqYFtAYytXOmifpBeZ7mjESK8VCIKXhiT0v88
Om1m/9goSV0QQZ+jqIZg8XU0OYIABB0hs5FSXkUy+KrdgGGcb8hKkscmnkDhOCOB
U+w+zh7bt3/0Ftddbd5J9iimr6J3XBj6tAmW99FRwiaPc48GrQeCCEyphLT/rgDR
ChOReV2AfrjAWEp/o37c8SoTDnSyh+MA7l7pc3luH/6ciwnyHjr/UeKQPxHZGHwW
nd1yVaxixveZTAYTUmpi4UcaNnZhpV5XembdUSjvAB/ufA4mg9F1H091V+qpw85e
H+F7hpUV5mE9Y7Z5eewGL47WNDQc2smQO3WlnL749vVglzK+Es6y9YRK2XGuSNw/
OhGj5fT+0Mj7DbwSJbsgNk9+0AI3i46dr8tqCoqlkshC89B21GP7KODzt429pyxa
2JcXdSItf6651kFa86Mtra5b3jCQuQngJHawurWO7qd1lOIyDdf9Lk8nmH8hL/gS
Q3mvP7cROHnJkL2DjrDVFkImmOKAnK6QdyGd1QZuWaH/owVdof8jSkrnrmYCjaDz
0IWW1gzHqOmn7STlUQp629eb8cURJmjoUDbNGhGz/BRtF3ZSWcyHCTOEFqcz/t3i
ffXJcY1I6VRJ4OiRJNWxdeKt54HcqJJDc3fdlQLVNJUUppGeOS51SgY5+WwUkudV
x8iyRfuEmzqgHBb+th5ALib5n9ZcxjvOwk1RDycRh9r3YAYYVqEDxaUvwK5+zvVL
GuvJy8Bdjkaji7/JvqAe4RKiJgKF9kGF8HZqeBUsPY7hgFlFshevG7F4cSIG3zYL
997d/7YHKTSab1gsWbUu/k2Km2fzpeY+9CXkv4l/jjwbtO60TUY1r6Q4mNU4Dqnu
pAL49eVcyMdTKEZVMjTzu4nwge6nJPyL31ireKWrQXdQWJ8qdukEJMyv/3w5XIgu
jLCMzSx/K4ohys8raQyjv95KCKVLboIugMslB0c5cz0eFTBR4Fut11FpERyIHgp/
olzv1wYIThHzRyR7LL0FOwNDibzB76yWZDdHTZ4qG3RNdSb15hqaegvcnGdxOwM+
jqQ3D0020BA6VUgb2nFpn+jrBp+WsAZoJH86FQd3jZ7rz9wTCYsU4Mt8ARhTddOI
EiAiQS3aiFpDmrbvkmXCuk3Ys061PBvj4VjqhfqjF8cJn7BBVxQNDrFBc6HvHwnQ
+5FWzxtSuJt9lmuFTCBjV4sKdyITEBRljpGiqe5gdP/PGlVyUwpuCFTcYiY4wSN4
P2g4+vkdNfcDy5OZNyQpKXSi9sShAjYz6pFI98lgUusYNyJrns+yXFXWrwawzDTO
Z0ndFAhW7F+r2fXpt9bC8ZI/roXBSdw/+3OrEvh5jLbyAnASj07B6l9EnKvSljQs
Ryw+rRLaIpF+Amf165sGbseRldVn+svNNUiCvNhnZF56uA4ltR48GO8BxX5wgckS
p7DnARg3DJh+lWeySPnLH/rTAzrUQsPs4aO+OWdx5dLBwjiafTOWUY0m8GTKeEbo
bGz2nC9DhQAo8NZfTDI+bigEGeurde8nC9m9NbAUufIQWJUO4kzCFDqrL5glwJp0
oxo/44JPN67aOCq53h4El8rB/owEerofEXxyP1eB7D5LxW8MH0JKnNls7e6X62GE
kgdOWt1ZxV8waBVq82kDtW2cWGgJL+mvMRcSpbXraJaXJ/pWYbAVH2XOvxqtoTkl
4oN7GmsRpwk38P7umuZsx8JjA5m+SBuF1z8xZxHXv0uBT22D9CQIYu3Y7XiHnznn
o3U6WAjUsSXdIGp4KeeVkSIX76GdXtGHnBZd7THAFWt4WNZ38I5/7tlytr/RUqFA
f0H1AbwD5nF3pqJNnUXBjHyoMNQFrGr0mFMnSPAAKIY0KlvBdp/IHFLWHnGCZy6m
7eTLk03eDG2lvEDnZ9uSP5S+nWwtlY53GeTwRC9eGgQy+ejvNtdJmhZS2KD5j4UB
yd4qw7obxj6Kk46j5huJh7lZLB3fQMjfA8roIhQgsXc3dJIxrvNaDVd/NTgrw8LI
8rX+8GoO8swOC/wf+OmVvbdGPzyOWLBI4uMfHA38EGBuKykXEONxUu/DIVyB6WEf
jUfAUrqVjX01FbCPwSGTVeS/95bVaeOyIcczkDOKWqpXf5KqsDxI5z03HvGdoemG
KTb2t+Nxn3J77TT/BqyEYCzN8s74bsaJRppDLs42kjS+gB31PLgIfJpRYpsJrD2S
t1hyb0JYx8Kuflm7mVlnMXnoEpfwkoPyHUVKNjSse+AG7BdahRwKVqHVOhPAIOO1
2L37CixAlsHBjWmWAVIS1tsYrwqvrVpRSub7X7UeEfEnp24eA7QlMroq1qAXMGQf
+7jjHDcnWgcobAEJkFXbm2QTPKOHnJSHJgJHfXFZocVRg7skIG+ot8jJ1roXeibl
juiaaW3ourUT+qrtTUydNsuCf8DRfE0Sxq6j6ZSMLKvsxczn4SQ62esYpWlg5Sm9
cXOd5vC8lv2uv5Mf3p3TU1y7Ql1ESnDhIHSfba43tllqF5xCD6BTpf6NQDKtmdec
cDjQlOa444Z9P50xSMjjByqbSE3ae3D7vLoDmSipYqyk+HLn7xF+e2+ChZ/o8IQR
XHHojyvLdDlFdLXhT7DHn7aZWpWaZrupT2PRSSMDZun2oyjuwrp7bGIejubRtLGh
G04us/8tNxX2fml/52kxSBEvnsKj5rR6+mpinsBCDn8ufy7uoJeGVpb+aU0crmsJ
EpnbFKYJgSAtdRhBBEyogLGJ5WZGpvqTVHaADlwKqJH96R04EpUPqLq6Fo6r6I4o
N/ZmxkfSYcEg3hueW9xIi46KyU0VO/QNvhaeS7/NovdT/eUlKOZ438tOnj0LP9pu
ukdiN6mJYyM5YxaUkb+OKvyzGfHN1FKc6Ok8SLu+uKlLBA9r/cCC29ONagv2QBH0
S6MdmPRHnYvMu5GjZNEkDdmdj1TUUxk2xw5TSDkWbUUMHSF6FqaaIJEPZcip9zMm
bZYPLs79CY0jguePFo4qVxUVDAZojjWSJty+bODxkVzbZwpaAf3UvYwvydq4LSfe
dderX5RtzbzJXM0ApFGJCG5HYYEOD7plIKLNqgRt09dN53t5o2+NYWOyyR5jULfs
2Cw6E7Yrsb4xcVm3S2M4uwUmn0ikhmkwiqRi1QWS27aOJH3xOs9Yhf6bD30PQsuM
hnGpJkEtrRM/zwh1Niz9SKVXMrtFPkc6rAGQTOxyOUn6THOVa+nsHg+GFNR3ZBSH
AzJ1v1flAeseZrTgBO6bJLqKxqzSDQzuE2IBgDCnNu4sVtIdeQ26qv1z9AdFTnWQ
CpynoTd7oi3MfsXuhTwTzSZGg4pN2Gj7g3kC2zEx6kqsEnQhWTFMT2cD6smCsBdH
4w9K/m/jnn0KzMSm2F6gjQ+FphPZXzQ0/sRNrdkezN14FcGtbCq0BsebjQvCDuug
s5h2HY5a3ttvE4wwSJ3OJs4IGBgOrBNmFUDPepvq1dD2M79B5qboluu5hjMh1SVb
2PF34ePPgJF5uYOpEn4ppyL7WtnSWA9SENjsSogmosfQNvgty5x4h2sP1YzkELUW
kccFMHZtcYwpfa0wq8lWmUM7POqmQ0iq/buTwerIdmLneYsTf2jybmras8Ukdn9z
/Xh5wuKqLZHHNnu3VeMTzLz/J2VgMKRWLbFJof2T36/azxY1qqE0EVxbYNNIqJJq
dTuNPKpF/bcLuhFA2ATAE6YqPn9c386LXUarOqGKYnahvYEI8QauTQtxO5+bhlcM
hyB8J6Q1b9ujaknGUnVAw/L5kPO2dfbZosRT0OQyOUxXSmX2g1spXcocSn7I1W5S
zgzrUZQaiZWXsZAKdCt+5nRXXU/3naLxeMoPbw/zWHovfluR1ABhTlt9Us+mWyf7
W1gOrh08QK1dIhlreo6bpvG35B4gHqQdswVOjg8e6tXOgTlKsQRyTwq9YUCT47Kz
sYdW68Ub1aWCoQxRArTVclZytyuDhwOP0yHTrFt3d7QF87NsBnI9pMAbvRGyyYpY
DY+1n/KVuQRFfpgnVH79Ak/CpU2ay3+PJiGtK8dBJgVvD3laIoFiXPiab9w+LKxl
vHyvFKQMveca0cN5oVJ2uTC94TVqAMCAjSw4NGUdFcZmFTBwq+Jndv3RkGPtB4Kw
9q6N+BYkk1X1mDxHy8bLvqxjk1I7RCi4YLRE9YUM4IwLIm8nNgw57VsBeJcHm5lc
AJ1G7/GpdCBh1Tdf4MpmsJ00pdbZRICK4l5Y2Wyn4MKQcBBA4WyulRsAv9YmTkWu
C8q6oYzNN+0FsnzJiUXmgd9D+RBT9/9og3bJbPpDkzcTKH0OKpyOkhEcUglwNl5F
9kVok9TESESo6fNrNfFjsWl/+9CgWBolQkokhh4+gKEVU1YKtt1NdagcTfLAZvnT
fMmjW4+BXMk0UUkFdOKmP2cKKPJ0YTcd+Lk9eTEpFiQNne2ljGWJLpR3gZCZp6LQ
wKgS6gZNiNrVsCIGKhJIQ/aAVavAe3Wm2HU6Wcr+9ECU5rc0RmR1Uye3D01sjcXu
COjpu/EQgCynhOT6F/ZhuRtCuRQDQKuy0Pi97EysBSctecWKQ2ksXwje2xhQFizf
O/LkGaqV/gQowgHn6sMSe4UAubhTTWc9zS6xfLcC9/FpacWWukduV2lT6Gp/YaN9
+BQg+JNRVdbbnRBNCjrQEJHd5S5czKXlZDEpuJURP0a2oc/7Jn+bQ0nrUBwtWWlo
An8ANNr4TiDErP0wsMxnW5PSp25b1kcrttDKC+kTmL5hTEcmA810JUoyrivYDBWY
2n8JZL5uswBVQ+RSkXl489yUaeEMs+dtLZMIU8UKHJeupPATwsn5YN/MskdMP4Qs
UgmuhQMq/D1wpWGvskzB+OG1rhYIoysaaRqgQ3HypwHANh8o0yt6f+DJ9dP/Fj8c
oH8ADm4jSZCKKbPMnH3+STKRnRUUCR2sx8tKQLfnYz+AX4uPDlMqPr6LmRf88BwF
faRlZUSpix7i19P95lVXOb4bnorKL2YBZwMO3boUqcnCHQ/4gsQadS2BdVz9cpBM
0gUiNX7FVrRrsUYniqkOi58rQBMwCfxUaCNEvK3VVBsyu0htWTF2IVBmOYE3LfqT
Y3/GyO3RNt16F66PF78P90NlYWvQr0NIOc39981V3VEuVtkp4b0o/g+IDQwO5B7Z
+TiR+UC61DFZR5J7XTVLmFESqtxo97DJ/tdDCVK1UgeXI+OBhsa8aCzyxm4kkU1H
+YbvFihpIOefm1VCSjvSZaGbfSqSWL+5kM4L2N+KjtGSPwPrh9MqCXI1ej3wfAOP
qIw1u65qLwFSpJ2BwmO8ZrwZnKe8rt31oOK77pZClu38OikGdG4qIQD82tisFx2r
UnurLW0DLYr7ew4ZUazi/0fKTqBedsX/gGRUNjDbIonwILrzhCku8HpGH/2bfIkw
uJlJ6vEqtn7v6XAfq0AWa7ygPeIEMHqMp9iaXyahiP4JB01ijt2UBqORJOEYhNVW
I8yPoL8E3Ew4w/4fR2fVPBnO1B9I0IM0nNDO7TnA8BcK2R9fzVjUyg0dMXda+uQl
4Ckk7uJN8ZagKgDwsV9wMQWFUUjTggG4f5o+2anZepGPOWaQBmSMfnK5xYEDvX1R
0T3LGGydM1dU3+kj7Kv0S3MLL9K3vNoJr6Xc4stplQ2a+AD7gbmVGpKS2IJ2DK9W
8ptp5UggNRuAxL0cM2Tsgsa9T884EdjBoIXYIW1swXa59n+s9UPQ/t+hI0ODrEJt
YvnehzZzHfgqKjbu63wd4rGncm5T3gB0/zMBJb1/76T7dCNtI0tGNRJJk89J+Qgt
Q2Lzs/kIrJYhkoEFS29/TFVkQ7p90sIW+eF0OE7w5dT8USMbO8xnyrfBfS9yGRFS
CPBg5ne7k49PK+UvLFKkMwNCwDIryHL6fPX6Rawp9Ielrpmq8rbIa9q0hAe/+Uy7
a/K31xSMN5JPtlN1NiMB1xT5Fk3iLV6pSfsrA5JcPhEPliasr9kkfijlx/6mq3AR
EjiiXr93FB0FjlSeCzd5VzJGVDt48O0Np5d6CmwdnrbU4DDO9KIB4wPmkulkntPK
9SdziTmA0i9HHVOktZsAUxbTtdSug1ZpqZUvvBzFwB/pWuuN5KfHCUBxTDAcl4UU
I4D9y1UImBlkxy62hiTQR9Kz97cRzeqA0cFebZdh4R8pGmN1+v3yW4it+K8N1IT/
0TaGg5UT7sBDmF8QvVSF715nS/yK+gdmrSENQEBzWeCnCUrCy6SJeVkDXYdc6iCx
Fhh7SvDBD01kTPzJQEBszA1AjS7UK2n6tJAHvdcTnRZ2CGHQd1eXJPhXZk3S08Fn
4NplxCGhq8D/UnoCf++mLw1Tf15232okgkO3807qB1I5U+PhuA5/4YlJ2kH+gvFV
tUqsUQD+bC/urEetrUndnbzbga++RdpdDOwoaHSOZa84I4ZthFJIdFJYgIkAhB4w
U8Cy/Gx5TZ3YdSFiiriZ1ewvuf+IZSiUuLQpN63reqFsifCdxPtrqc0VDl6l0CcK
e5q8vd91b6aewfQsoIYX5KnwVUEoKVrfahtXlYwSMkjMijt+999isKS1iGu2anSe
dQ/w0RkIHt9lilZz0VJKtbjr1j0CYohxyRpdplRLzg8lcQ4zSc5XZoS782skYrt7
y0Rp18kw7EZFwYjzmGvSUylWTvi3hZkthIZP9FmbUQ2ZGaSZFiZd7Q+Ia2R12ED6
B4vGiG/TPOycvR9J4KPMDg/KLLg1KjnKnlxTTVEbm1j0Cy0MwF2G8Uof5BZhprl3
BdoWUQ/bFQe+/nrp4FJ3yBkVUmRXZrTommryH8H9DI4EVCSNVaSLzSZ4Mw707EUP
glN4mUyNnnN7nryeU79jOmRraGTlJ0HC9RQYw6jn6yDnkbUVWWf2hxj3KLcaiRFe
rOvLXlHOpB7lEQXzoj6lQ2yUKaSLPfGGSlWQYxNez5EOFKU209yLEjjqi5FYpU/J
Ut6R8gUuNm5qnjDbvRA+zEamYly3ucnqSgjBcaHMWZUDZ7qLMwwtMQrXNA2kYOAq
xxQD2VaBEEeZrYRORAkvcNi8w/znLbFRiQ5BYcHcrMQBthfVPPwvD+gxlclXSRlz
p4tcgDT/Xn6E+oI1mpfYREronSaaenQ6J78vuqkd1GAocVp8rrGtHn6gSrVMSJha
9umWacxNonI5paX0oQh9D6NyjudN+TGfhWfYF6XHYgva7xLQgRD/saNvWULgxQLw
NjDFRIEeLLmHS1qzB5v7LpoOJAdk/7DUy0HGhGAdsrNKl+XtH2BaLYz95HXVMG/d
hoo1nBH+3ZQ09Ae6pIIOlFhM/TPdA/ZYN0WjRT+fZZyajyW9sA8xmjb63oufdIia
evhuuwlnTulau4ElzUTfT2Qdwz9zvUeIEW1urxFU5l08jarh06FzX0WUtMAM1l79
1QOUVSKESwWXzL4kz1NM98qiCONOwKtmwDHf733ZWHTKY9cL0F2jaVy1MX9g/KoU
3X1+7L0EjsJ0lSuSN6BRX1nLCmBjF9CqpG8AHYKxyplY1fJlIUMnp9WArVWGbnGY
Bjv30tR9Vk4e/gnPcXy5al8Mt+77imB5VwsEu/G4ZcaV8rYgPqK8pEIC9cbGa8Qt
NzOdCVVQR214MkHNuOnrx3YiZvHxzlqsiHgLlXp4gE+wQuw7gJZ0fOJRTv5kv8rl
puV21xAlHixXdNUaAgJRC/Cje0DA29X2OcgSyDpV5eevGPTPKsflIxov6q7OvkGy
QHFTcVBAEaWsWCGbbpG1Y2+SVgglqsNuqCZaV36gjXtNzD5fD5usvf1IYwcxyltV
v8SIOk+OGXmGhlkEg7ATotKi/B3t+3+q/Mgx3xYrtCHVn1en3YXFGPEmjpK8/cV5
iFfWtw5ZnWuwGgphk+AUXLIwJqRrXVv221ED4XBnZe2C9tjdkgEWQ8DWQl5MURlA
iAGYodDjNVwQHrKl4AR3Jg5nWiOJAsf3mBQRLEuZWeMnRj5i64/0oEDR7iu9ICsK
U/76X5hM0mvXkL46CvauCY33d/txb/bhJ2zjnyp06biCDYBGugOq9SdVg8o4Q3sM
TI30ggAXV/2vEq5jTEfvMXwmFVZL/fcBf8m4b9jf+83vmJTw9nLOv33f7Efx6L+X
jG7uw4cASAJXwrFQGVwJIVIdCRSgQIzzvXIwRDfGfyAwL/WkUKKVRkudb0IhNn43
dpl5FkzF23bnJUKtfIxq8+zgrPlVr7POXG3134hsOynATWpolGZZOohsEb9ELSQG
tXMg5H+1DpvpG4HO4/TUDCZGit651p2wYVpN/QpR18moQyjZHZ77DvLOHFDqul+9
FdnpdEfl1JkTgTMWw/zcguFgS8E0xQvtPeClwq5Apq1C1Ifddpx50HNANf1SwiST
Jlc8GWejtYqCiIkjE4R1jQdI5omAockmhdmj9f6al0LFCvZcFvjnC5ajOOxA/7qP
1kLySrM/sP1VEy9BTvVFLz3VvPqLUlFlgcPRns9OyTLqixHoVewWcOGZNbdOoXvG
qVU8RbXFkxzOmitWZ3g9PeXEiwB1NZneacKM9toS5BKxE53czWZ+Ln36CPbrONQQ
aEYhmmr+5BeZporJBGFdyb95vDV5GTvMZuVW0BNdns5R0eypALpKFZeQ0nOKeUQZ
Tt2j57y9vedH+mGhIgSFremPFP2OyVcKMukwME3hMwUo4+uDdWToZe2tz+7Wtfcc
zXVtZbVTdCTzYrhHmTWFqlEnUalYAsa3QjaQaURVevCoJb65pBEjJ1RAzkm/KLmj
z2EAA9n0l5JWcwDVtHKpJNXqf12xoXXjkrq02FmNyvOSyx20KvWqLdwPOe6sj8lZ
YY/Oel3pl07JCdbBrTbMnfYD+/p0phW/1WrnpglVZ6a7Il9ETfgMQaa/ETyXFxOF
Nzp1a1gAnHS1h/GgPCyQs6JaSh2116BHDPy9DwepYP6C71jqGa7mLeFcpKQjI9bQ
iA9JX3zjVssT+AHvhVMxoWnQFB/tLp3RZbPl6t9FX49cMW+RRuKs1js4tLdtpSkJ
9MgrmNa+9aB2xbmq9WePJrwVhnncA9BMc7Pw39rWgkADvHmCId/HHck7i4s53UaR
2eagBS7AzMrqc66LvtU8dMho3JbubNysoS6KK9iWWhTdZN9Yjxm2O2TI68Y6YTGE
6Mr+trQM8kYlhh/zPBxP303rYdmLkh51w68309IwqWdOak8mc7I54WkfD9jMl59C
TlhxC9Oxrwc3tqaiAuXiQMqwVBnaI7Rt0wKJ4xVDhPfHlbRg70R0ednTBA2EQh5a
2pz4IBUgZgpKqvEeWCKM66sC7sHx3gNz1w7j94uhtQWMtSMP/vFo4tYz+8X5VnVD
vY7LrMwcb5xhYnyiMza0N2y8ekBOFFWv4hRWwnDUYzyMCiBZGMHz7whD/TGlnhrf
iAdr35+2CNm+hQn6FLfgvpk9QBfgMJfVrdumUdYuebcfRBgGaHpXharCkBxBIyL/
wc3oFWSH5LeVVjcTybzYSVAwa8FOe8huFIPlIDhY3PXdv46adWE6an8TB4pZoPyi
0KkcuD+b31uhGV8KPyHmQjDkLH7ponFui+vfa/JuMcSHlb+o2XPbgEGiKB9HrIcm
3SJEEfDAtHIX7LMs6BwQL9thcx1iIGVVInhmU/VvX/oHjoD5cPpygbgVJ0DNyLCZ
dj7IfUCBF93KksmWbwWhFvRM3RAZ9rqE340JF2Wi1+bAnwp/aycaFRO7JAb1D/pA
IY6DhbrZ7jivMTnkCO+hjwV96xukreMo7rRadNbtaX7MMdjnvB0AotnqS3puz3hL
AWPDvNyvXlDIw2LDEYU5ynk/AAoDf6HYgv4yDWME/IkcJkLW3WHcWq2ULWCZoch9
6jzKwszQrp1F+ooTFEZDP+s0mgoHokuCK1Kq+AqXMe1E10iWYzvSktOUnJGMrdRt
aBrhoW5/S2vhlbf3ijhd7H7+eXzuBb7MOzHtgKXjuGwWainaYhMDslzQlaOB5EMt
eGnQ0ac6+OR0UOLw3mNrzuQSQuoZFajBERo1St7Op2fZ9EnGgkpeucDE/DwWyQR3
jKSKFc/07racxREYfCc6ydAKYHhOTPUOsA7+W0B28A211K3XsIdGwYhl8dGIEUbP
9TkU31fk1iljF0eK9iikujibMGxuCjPFB4cGnR30ah1TBeqkIkxSxPR17fMr6YUs
s35/d409EIrsAb0a+6UHf/kTCWET3Q+X3OLRit4hE+LQLRmVAQG75waR9VLT2OTo
9rSu9KU+vfNDSdr1uIH2bmsGYx4KhWqovjjpcVGQ0R9kPri685Ex3pxAuw0QL3Ui
qifEWDAT0/1oPkKhvlPssQURsZfxFXGGazcUfD4NqjpSsTpwkkf7CzBkt62SATsZ
QXFhXYd/2iAhpKqttIHq2HTWnO1Rq78BSUZcBOpjOG+far9w1tkST33GG3Dctw4J
+Z5jQb2gw0Zcez3X7KYAL+hKBnW+FLXEnb7mOYBGUyb8sQdKX+ayx1+1PrpSessY
z4a57FrADJTr785G2VKG3AyIqIUWEBbS6BRFBP3RP6fows32ls3PGQKEOJCH2C16
v98QkYuD//fytN6+SU3OqqVWMP0bES1HqGz/vOQfHHVh9AE2y/5a0F0llIhfaQrv
FFFa6yVTkJ9cF864ttqxjLP7lMjmWu7ucPYpvRjoQvjJOtbCCtwcSPKLYdwWcLUU
cNwysCcIt85TehURtIiz71J7NaqO/UybutZYfY4m9J1FhC5tDmuveH5sqjvoHYH4
tikJjtO3DjJguTcYI9iJxHiEm9QBiqJNVy8nlpfGSQyDCDcoW8l25Pubj5LG3Fwi
0OKSmA5lSloqhp8NtaK/JE1dNnSfQhzELzZ42RZEMbq3vH2XGvIzfQCS+z1LpvBe
AHhbHEV7tSuDHUKMgIdD3kPROLdh4jHODNQvp5R5j+Z5zV5ZQwVjdpU2eBf5L2ZM
dIMrHIjVTJHQgKHSCCXnMS4WhO4i0DI2p64BmHKzWrawoP19tENpucjwSKAApzcy
15LlSMElzOIFlG6ruZYjoLEEVAbKn8IkmOl499AcW76VWKTBEM3AdEBN/wDNINa+
Wq4aEyhvX1ftvHQsEtLbS6H3rOtsGOkfEwVWoVYPS83vOpIhRppIVOWMRFsZeoda
HoPVw+/C3yOQ8fEGnpZK6dKd78SAXwKbZwsy2wcQWEzWHU4CzCbfqes4EVie9bwW
27m+OfWi6/mdPQFGz3uVdaiwOazImKsRUsIAnjw6I2ovnSc+SWd/UQOwRV5Jdgb/
QAerlQJhcbqRqhKx9McyitUd+7ez35c93JAxysHX6Vrf5+U6/Pw8Kd17LK4M2DQY
ib99YI6jAHcuAasVizDG3eGtuRQgs/n0Tn9uwB3/O/Y6C7QvvCZlUEQiAt79r6IL
/btnFBN84BALooz45qzn+sCoFAL/sJaiNQugbK9MSX6/frWYHUcPXNRlVangjacX
bnB0+0/6shbhjOKpjOSFew4kgaWPf190i9Z0K9dK8b2Zy9c2auDnapQAUHlaa6mE
2SegDqFKohj+5YlmLK7fZkXnKzNBL/5pJIJeYIsGY0AlCf+68z0TsaRNinCq+wwv
ScfS2swVLKscgSRLEo370rIPQAtQR+VYD6AjRhqQudAoKCVYSvwQY7bWg24C9kJt
6PHMFNpKaxEjI4PDhkbfpWYSoM9LbXumPXr9tX0PR/m7Jg6P0eRtjE0iTQ1yZcL+
1mcs9wJ2SzVRyjAat/9L0hCsocBp6rQgWZ3IRNsMSDW8G89MaKulk999qPW1O4pi
IcHohnUzf2Z7rL7F18BRYJBtSeDfYHp0C6fmXZPdNpcz0WqJAHmYQtKEbj9rTHmO
qqWvlvUQaDrkm4+hWSv/hGJY3PDU3R6IpZmKPb+V3uFlSHhUp5k8Am5s6unIu1EP
5udp7mlojfLyEVjqQxKHNBRHYRxdaagO4jzrV7GfNa/7A6DJt3ZK8azJJaygnoFJ
GtUkp4VvZGJNbc6vjRervb3xg0fNFOqrvTEqDqZQz5613NeCK/RmFs4/rNzTeJGf
y/Vb0l222Eg9ahXC7rWaCC+RSOkmziEXhElKK8uU4mFN3holdDIJFtoBxkMzNUm+
U+dwS3izgayThC65cgn1pU5kQmr7kSmEbYQsLEdn5ZFLk/gbSmRBNL24mWnCjGcH
ucH2zHTI3QcqsR1GgpIS9dskitqksQpAFGZdeiwclISxD2cbou/7oZ4XFo0VZfiF
kzButATHQ7+QIRcq1rp8haKOyQ8kZTDq4YznFBn6aTXINY2ejsEXZVijFS9OL7MZ
oQgDD7JRK7n/AmdqeO4W3CRuCgF3AtQOInjRdE6Ypm46lt5mJpSdLabsP/4sb3S7
f1TmVxixF3r2/zZjVoEvR9yIyNe1acYXBoWoCsUanIhew1GnPQGDrhskfswCbahG
b6MzZz31wZYIGG59fbYlSkbtI5YXh3C5LDIvD/3V/deex2mhSOyBycCYm2HSHU//
f2XkGYUNv/+joIxucrgtMGHhMNp0DPGWyFOIlhTZeVigN7fhQaXMY+myRNkZJZcl
LoiFQaieJKoVFf3QAdC3EhXw3q37LFiPqEUOfwwnJrKqmEaKpVhfeL7qyZnajRI0
j29Vmi+hRG/4TIZfArXLEGuPH585LLCHX5IXVih5f0TMQBQl1Iw/Fv+gUL//pYgw
L9ZPtD5IiadNhSOkVqnbXyeUzn3y8OngXx57bbcEhs8yPxpliZki/ZBgBIHIPKwr
qu8usWgTBK57Ff7zqKE8PHMDrXbDINcgFJGkO6h+siMPB9c9Ysrh4cnD/D7EDFD7
aZ280sipXYwcOettvMGVaVP8D6Z8EL7PkGePWtHGpTMXaNBn2WpYnTMIhc5U5/yg
2DHcYndNchxON0igp4e37KumdzcjUlz+1jLMvdKrsKq6/LshWXcfHP3GQ/u/l1Zf
XnOsyEM0i7jnRoVzbAeVcQcWX3v7I5Ym/UbUdJOGePA1VqBIgpW8/SljRdKRhPN4
YnBR58H9nik6d8727Nia+yI8tUaEdHHHE6paUR5sKPqfN0vu4AnlagbjaI01TQCL
+mkIoWjXc4dS74vLhIg0LDtQLD3KuJjHOiohpLLVaQFohxHZMfDv3OyVwZ/f7i11
i6xac5UaB6KIDIJ3HdSK/FqW+vYB1106/r/yhqvXONGqJ44dxuhEk97Q3Ae07UN+
Yp7QQqnH1o09qqhM8ldbLHxr9Uh1GgDvwcekOJkHVsG5XCpsUeOOlKsO1UFyzcc7
YSUWnLIgRw5PaFOCynkBvig9hEBS4GxvGh3IlB7zHSoUTxkc1j7EcE8jmZkua01w
uGDVxG2MWSCyaXpLPbnrqBCgwNPZT9lpegZ8A/sTp3u2eB4EbnxgUskXHNMEvDXs
uLQUUNa8P4V6A+vA/ZdyI/a4e54xTDl34BNwa22XdLHUodNfUcIW97zqkxIPHiuP
GGBZH/uxMroLPHm8yMSlzers9nIrm2X9rbexUnnJx2pQ5YIlPSGaacIxzz/rCYWI
3WlQiLea1Z6G42PWYXDGxq8oAAUBQYy+kQ8qXmZ4B1m4zEVe6+ALzVTpDcr4MEKu
3nLSjHzMqT9GXHfRKveyEL2Rw/DILXUFFY5o60C/NmkbvA67s72yR5jPvLkShzCv
qWoxjc14EbMPnCrpTVkSXscsZ91Gzi9nUI8yFSCtgfoOlO31+MEqss8jJmuTdGP2
sNWWDzxVs3bv+eOcIHCC49wxdC7TKGsCa0FPguF5n6nyZJeaABg2o+iS71OTkw/N
Xb28TK1o+jMr9rZqFMYTKhaX2kKJqkiVyUiluhS8AGIxCuBXLwYtoTPYKhFALmIe
+vAy+v4GYv6dvSnaacYUa4KZB3VSoOAZBYcddfEkvoyOM/X4l/k/0jT5EljBTRHy
m72fNh32mulypPupAAGW2FZRGNcQ/YNhYBj2p4iX6z5cgJY73ZSQLfF3l5nRGBIw
6q3oiJebF7+7VtYrMO+lUoay830s9l3K4h14DFXG3de54ez46dkSSy/y/spJr7/X
GW85kpJSfUPvpOuV0OVEbtSOpeQP5RHwmMcW8Dmff+WDqDEPOp6BieH1V6FC6ajD
makqxm+M6hVk/84K6Fdnbq171xjQXMl0ETEhL/FwVVUCuXHbcTAnxsOJxp1x7TW1
Y7qEewuUxhAVW0JikMfqq3SeMPWfEPwIvr1UYqcq2KccLHp4ICgVPh642dxhuacc
nM5/TZty9cptviDdL9NCSwU49PMawR5iXasVdrU8WKNrQiAJX9TcKw2/XuqUZflG
G3dV9TTKSmTVD1d13qu3v/2yZv4PmZ3xe9Eiwi0KaBq2cBPm5gFS6+qMvPCZ2p8j
PcmzIjNfXMrm2zsHV0pd+2BmzV5C9ufUTgiQDKpKtbAofWnj12S/3FiD6jQ7na9H
/N6D+krG1pLJruRhyHYmp3k4ZMyCApM1IFUy3Jd8Y0Sfi+3dx0sRX0LWmL8ZwVie
HUO/7jgTyct7DdP4vXV2dQY1uYgeacZlsvFq2OPy1eNTSa7Ty+BJx+FAG4KmIKdA
RV0uCA7/S4mNepMb7WPSu4QIFkBZnJgTOYLWxYC1a1uOo7k+vOe5aWlxQNV3nJri
XkA4JPhyl6ZhdDqJTYmUo+x+6J06t+oFQZerE/gIvApYhq7XQuK4soVUqvGqgIbz
LRBF4C/9+XicCZ2dq9u/VclFRcSNPPJfSFOtzuxE1tliFojQldiHb++PFLdtf+36
BH6EYiYGaobTyhYdXt/bfn2is322T5JMdCUqp086Zk7IFmGgnPmNxLqReqL9j0vh
H5/9ShH0ri2fbWMEPTj4+UJQhovdOE8kLhkg16DmAcgwasbTMXCJBUBrxKoYHqnF
SKNOOkrxAdk0Trv8hf9Z6836LoPUQ/5agj0hht3h/ze9CcDepvqPFXsz+ongu56j
V/2vyujLxCj82YidYdhgxjK+ebjIUTZ5ZqDokQJ02DsRFpDyT2K+us45+j5Ed1KQ
nQesw/4d8o/pWz3NREt23zDA8EQEN+mOiKFFNsRqmvY/0oe1RGzwyFb1lQ1NvxNl
uib8poPruAOcSzA1DI6l+WBjE3d2evh3//UIe1DsnRG3YyfBKiPLuDMLY5YsCLu9
cbeEGy2gTafxOvBFnoDstfPQwsKCcKEiMzt1trfBCLf77QxthhcMIbRBwpr15xrc
Nyrf8bvP12IIWtcrbHvOz7LORbEFlMKhxWX8sO7+jHhPKYpeqH8IbRganibbCpdf
RN9oU+ZXZZ2NEJGoVklr5ssDGFKV286bBpRulJGn8O8bckhRirQeb7GXIUoxWl/w
yewTn6zIlk3eslqkFeq6gaRqimsbyAEL2mR0qkT5bmJytREMZqHL66XbKBTm00Ts
V7pgQtGYaTTjZK8bpUBzbafn8sx4B/7u4wI2ecc9yn07mqiY2cPuCzGNbqhPaV9p
Kd1MoHaFLQ8sAqs7Uov2NWuL6LlTfKnhUS125+YyG8pyOm9QMnt6GQfa2dVX1UiO
95BL4ZCvulL3Z0HX/edKHbirSgdPLPZ24fxrpXmPCewRnaK7T9t8Ia4V2OEApIVC
8noXvxoyROsQaFfOSYTlp9ex2DfxdvrhN3v0lfhxSRA5+vN3uwzaFxHLPRsghkx6
B8lVQzZC+Rc0hurUzvhKBogk1R/DZ81PN/EBFcEz6X6FkVtXkVTzmA2b8aDJf3EK
vV9Ux23cW3JwtegY0DUL3dabaAw3qgzSOeb/dz29aR218YpLgLtDzvixLypB7fst
8ip/tNIfIfDq6JWZoQgonHIardROdRdW09Ghh+gbflXpkf67I24bS8nt9uJkMsfp
cnoAJHcRfk3A3/4+DRVCOG6EDCsDfp5iFRPguywWqgA/cDItVygWZkfY8pDTwQVH
izOcZ051KIZpCD2hyRITw1nhhUc2KFQJFJ3vhT7ocybeXSFjzvX4ZFac6sgvovlq
gTQPXQoW3fi110ysk9nLo6dvujln1gtrgj7XCJQVyFtjxCzAdtB4DCxU9ARIcyKq
7qXlyKa3cV2IsKYRQv1zh7zOhoE5jysxmy9TgtE3DO50EczrLolH6ABjbk/ugv/b
v0Z/OdskvE4gAeFUJWuORwxyjJQKdsYfvXD4tL0z7jZAULV13pl+Fdj2UTSm4+pR
F+8P7MZOX7Dp+J2y5dWAllz+R7/Ek8pIAIWEFEJ46fgmSr1RfsgZJBtU5BEBtqUU
qWn925kp8zRe4CbfddpWIOQkSfki2jxhV1L/NekQD0ZzmpuMcIWq3mO1YEudY+CH
1l3b6daRCLCBvRT9m1i4/jp4HTA1/3AiArI09CsSC8SzW7Lo/xwGhm3LAc2r+GTo
9w49WB6CL+Kq+oyBeTbIeahbwB2iUamn6TjriIpDqLn5DboURzdmBA3xvgYhNF3h
V1yzNA155HeAmbRaNujLat4G9bJJPrNK1dXaRflRxP+qs3dnHx0bIIEfUOvd0Is+
5Atg/z4NNRd37u+H6fxxAqm8ziLiWchLNtn4wrLXXTTSTpr1KRUc5NNJ5N7khO3y
zbeMh17ZDEt+KALuOB5V7L7MMfAj1e6pYGwhObWX5G4KtZmTNWYyP7IyrGUS6RcZ
v03ZlWCUL5jNyL/pWxFDvZqgiddR6g/pcmX18wZhIFo2FP+pfIjtZqE/SvpvPOe3
wdUio/y5iuaA1/O5VLI5b3OLVIHuqmHZdwKkNK3uxfsoyzO3erBfaI5XZF32TA2Z
hERYwI+QxkDJpPcmFKlzIAMovAxNEbhnPj6wYe51XnXXYDcjRfXUUzr8Hch0phJI
iSIbLCzjMeCPOpIbkIcp6w0u/4LfRurY3I4WT7NkLNrwIQ5iMt96k+Oqs7lA4PF9
InfdxCQZtN+8KTXPWS/b3SX1lhUQ/x5gfDI0Lb4wd1WGJAPoifEQgCyfNpRkgUJT
3KoizB/GBhvwIQfMMihO4dT9bQI8WPtVrXPEEK+2tVOw2/bgoqlP+DotEKBUOpT9
UunDM3I0s7HHBxrO2zIVTclvt35HkkYGVOwl6bbv0egJH38fLrnXiOj1eDdsCWjP
pCASPuUs+1WT+7ymPwdngfdgIb9FiwBk+8RDqnbkLW9PVfpEaVdp2KzCiUhYoL/W
dzKlMmezqMS+gkz1tOge18RgCYUEoW7g/zV4pKkE1Sv6gvjBJUGHQ9VFgs+VijM4
UKVftFDIp7fQd4iluxGAMz9mfX1Cq4RkGtLshTBZawiy0cqB21EcxnJQDhcNqbIZ
yS8j46O2bv5khn3E35UccpNOjc2QHwOIe6yTvnnwJgzatAagyDytJXGx4gNTFYj/
vNvTcCFFQSnM5FnkMsb0peYtsggpOabyT459fP0Xh2MBE0ceDEGaMCpU0E1Ic6+R
TU/KA4R/tmGugESHaiIVnLsxL8S+kYH6beZDtwSuwcTDe3rQsvc/MR8fgOB3lshL
b4TqI5i4FfpofnZv1y3cA1NzVTFXBTclsaAWAzPj0upf/oAUczrvgx/qqmQVWhNe
48WM8kC4sv74qzA/jvXLUhNzMZOsQdDFIiMova2YE494j2yDss/2zBbNcOFAEy/T
CFGioM3IhOd2N59cAhWddllMcsn/HcaaTvZ5MvOocis2W8hK1IRSgrpwBb2begXE
xXkT87DqCDAK5SEBs3ZjQTgThtqnqIDikit6QsK4yAa03AncLrqId8iEzcr6an1x
cO398VRQI+tOlBUHw44SNgznAw62/n8lBQ6oLcoo6+PqVb/EVR+CRHHYOm2cgGY9
eFS8hmboTsE7uyHRfhOMQnDQt67TzNOylWCbwDxnYn3Qc6so/H452T7kfYKd0gPb
1bbVsNOLItauMUP4hwekirNTO7Yqjzx62qtHP7kMZoxnhkiQ3BSXxLc/ci+k7e46
qASFPcqWr2oFvPPZxp3mZPDcTKdxXrDypensUZgMIq4rXV24aTdELitv0cXTAWz6
AntGmJsSEJOijhSwOEBIw24W1fvlwdwnwDBPBtkR3rHHAGiKUjPECrzKKHfY/shL
cYa2Ljdncj9pH6aVF5U/sEYkFec9fuoZ4CRSQn2trXsGiZvaDRMNvBn+z+QioOcW
f2w+FM9fgMulxLXOCQPbYV+TYmlcSDKC+i3FRax9Nunn7crBjuuzf7iTasB4cePY
5JIhhEvWH3A0jgZNe4Zb63FTtjdtpY88KEjmJVkYKqSCtR4ybJD0AwlLIp50Ywtr
TwuUMhntZj1BcubE9TJTZiDo7mWfjEeAPhXm9mJa75zKMdTIOAj3lGVShker9a1f
hPfB9M60X549Z0ZBgFFIp3yLPSQVNoXhKUpazZyQcvGr061aLnX+awdmIpxYwM83
zaU2Ii3rf1FKO60kmPNSpuNy1a0T5wimpsqouMKlk5VpcabPgWRE5ufLJozwDrnC
JifWitjWMni6xhfLsIAso/SlIK7qhVzvF1xJ9zcxRQe7PYIAkh8UFe6b14t6xRpK
80uBpd9lxd4U5qfJr/HN0xX2LX8vnDwmF1qyVE5Rxzh8lW7jiVe0dTpclCVmavzl
+pdvza9QcYoUjEfFIPZQeIYWQBOezIaVnt7ENa0HlaA6fWTBWMOPKCIH+CR2Inwc
4uPO2Sv63cA4KLOc21joFsrMaN5Pkqs/Qqan0sxAMdM/8vx4x6zSK3qKiDgpf81I
HsORC+vAdnmHZ2+H8aaypP9Abb5lqVCuWtHlxQy+Ab7xtGmwXvx6xZmmwdgp7Wfh
5LwOO20nYa5GxVHSwXmOP4XqASzr4cDeF+T+uhl1HLI2L9CrhrwXRw4rzlVAWue2
QIc5hkDnXmckfyNsIEsWpPr5IhbolWgwZGaqSdC2WKw/7YGVRLQkcq7moThaU6nN
P0w/r2/A+nZ2hjIwfmljDNb6Xt5TIAZI8/U3c68TvLk8mqk3dlJJXXDCL4jzyloc
GVpufyWwuf6JYRyqcw9/lIrIsK8GUuHPbsDsnhUTpNFbyIz5iAKKGra/t9/JwRzL
0Lt9KxzAGqegywq+pCGUwDNb6lqKgcRgO85kkN9FQNLuWSkoYmS31bTHRRbu9P8M
UvWedLuWcnTKY9ElkylficiM5F98ISjFw+U6v7BbgVU6CxJE0VunpqkxDX9yFlqK
NpTklAJKUCmfN/Sc9Yra3hOcpZAhoNwWafRNReTBDOCAqCJ1fn0gDT1cXb05lrba
MeXAj1fVTTNnKhfDWPHmYudNu+ac2Q/5KErC1rVFDoHIij85a0yPCup9vS2wNlWe
7FFAGZoAtIVBl/d6SYQuUkcHOOaueIRe3ozjBzjW8kaZkiaXrLPtv/CwE0CU+Ged
PGRZGptw3FvrWhMppkAuNyfyfK+8ziSwCaj3OmTi2yc+hB4N5oPcLUKU8A/Tnzwg
PJt3J8Wq8IauBKNrWTUdW3lqN7t2FFC6l+O5eC4tL2xszhDTO1tDyyIyncBdWEr4
73bl5+4Jj+mXBf8PkL1JFOrDo+ukzW8SV/CwrIE+2lllmFKOkU4YEgAKOEi5fqRJ
meOHZKNsMdp+J3xs84y39c8gRYlymuL6jZJ8F1/+jDvav6dAW6hSq37BdgaqpGbs
u1NBVO6B3+WogcWfquDVBABbOtvQWDjLVBU9WOJYg5CPvHVDkhQ0dk/F2h2WUweb
g2q4WKhG5ScQX9cVn1ARcM9aW/DEVi/psfPGQdsiD75zEbV07QSOMfCbT/AitdI4
/K3eXOL/iOBtkqogqw8hX04mXGJhn+F2PRpzzXqno5ZCt1MsaJaOteQZwrKlbwjn
Yln9S2QEeNDeD0k1aWIdCHpZf0DiZ4ZmNqxE8TqtHRwM3HCwejbqEwxQpJJFzNbC
Vxd7ixtpwjXHeUo4ELBBVzPuuQtBt1cYT5rHuSoNBi/LSQu3uaT3RIJF1a0X2tL/
U8O/IIBSj2btjFRlX4iadI2bIC7iNJHjh87n4z9sdGC6yq/zXNeUJfI0HLfcLmOS
MAnhcvLxEEfxSD77CfUIEofDRkHMf9qa++OwtJWXq+GcjIdV/6nZouOhawI6PQyy
hu5WUMbZ2QmoG/4xUT0wiW+Xj5RGq7VVeC3dPZVADADKMtsjltUhKU8bs+p0QVPL
FYvg4OcNf0QPSQBIop+VT3y9e1FlcegB/HePLe0mMp6MG8NBRtTUKevcpHsmiCyf
KTDWYtiBdvQ4uk+CZX83Ec+JWkh966xQGJ6LWUvUy0Cci317xjVK3wpCuzVJ7PgB
0ZzmFbvbFlH0p4O++ahQFZbpbXNXfgqjVcqUYgdqwpjQOp5bU7QOBM3ANQcntzv+
S06dmHqyfK9uH+QOPhispFYlseQJzEucUfFe5d2lFYL7cuFQNaE+5gpevmQHi99T
zUgNCbOCHeEpq2UqiV47yOL/KLMdkbJkiL371JXoGfpEjCvYVXij+FTyP/FmOdMd
CP/SXNSLs2Wq5EpYUvCBur7GQB9KbnjfKRa8FAF2ACPdHz7s4OmOuCwZfn598AV3
dJbQMNw9ODpDm3MkMDDhFcoTQuXOVy3nRa8KfuqpODrAZQpK3jjJ3KsmJaxzb1x2
8XuDAtA7mWsQi0+PPRMsV3Y+91SYLVZsGuCcuWd7coNAKIiqXsj8N634awWxaZhB
jNWhk/tOaEDHpzEG7lx6LlBcvckvCSmhjjDETrGRUh+rl6aWP1iar3ZX5hNGEUKS
BSP90jibcYxQp9OR6jnlQ0W1n29FrQsTrlzReoWXVBn5bt5NhyJciklI61mU5UQN
ZuO0nDyAqszELiX0iz4574osu96FMxHt81/v+qZZEqI/7dJR+Dighcz3g65iE0g9
YDkJYnqXJG1dlzS8YJi4bzPiDKBc5bMd1dDHpdtY0Hk9GhA98d8aovWv5p8DAuzf
pnPklIvdUKW8L24OlYqCM8m2TJPqn7S41MqPWtLRvQm0sCyc27tIL2uO2LyQjm+D
fB/2NkgwxV2mWC1F4a+I/sqBpA5qPnRWzbGD6AV624Ynm+PQDvX86YQF41NlXdRq
2HaE0j1EZWB4F8laiuAjVnrPLza18j27BwW7OSfrvSYrTCVlkTsqjrkruuPNN5Kd
XmvaIPsbZVVAszEtyAdM/ch2ZIeZCiHvYmfQDxOuzJ0D3qe/KiD6I5b8pNjr7CMm
f4c4vtGwYTlUyBDMwsv5pq3aNdhfRNohV3nZEVObjZb//ZVQwhUfbTOdGSTJqkUg
iWVV0rDy0KZUdeHI1HTHsb3PYuYVI2hcJlYWHz7SOiEwYDvxW8R41tRVV9BbJ++j
0lk3QjsPTZY14XW2Nsdf9hUeaG7HwetuiqpAC0Z97n0Eyijafyn1q024nAtRWZB5
pi5A0KV2OrGYvcqrRodJw8sCXZhHOWeEi6tUx28PZzV924U7v4T9N+4JlByFUakf
9wLG6d39be4o3lSXUb4ji94mTO4D078xKHEYBgeObkZ/52tOHxTbIdkSfzqa++lv
iqN+F+0Hqt7WhDCPHW9FDJGqVaz4IkyVKQdUOp3YYvDTvQYHD1Pur0dxFLSiyDiL
JWyqey2571qmVWmAw/5TGEoEiTHUjkmomGf23jSYOehGMaJJc0hTQzdimQL90z4P
q3ounYVLsEjhXbOrUfNIV061gOdJni2uSQqyTiYdhdj7gqHmHiK5miNeII0anseh
FeFM4ZtBRxKLN81H3ThPNF+yrOTBLh6P9kp1wJcrVHT6Y8KAJurff+bXuLFhSPY5
AInMCqvcX3Evj92T1SjBky+LS7LbM1qyVAQdQDbIGub2DzWMR7Br2oiAl1XoWQBY
h+k4AMA1qUnWbK/biXCul6Rij27a7h90C6OwstcHNjYzYzAV35ekPtZ3LuT1GL+r
4VKEmsVNzvfFEfYepigqMlxq6C2Q25IoYQZi0Pq+z7stvbFE5P+dcqg4jpPuMb5V
KtLOCLlCnIx38NvAbrUJgyRFrDkwircpcdizNHnwp+uJHuCqEviCDSystdkb+5mm
0r3UMN+oZkseNPLB1Pcs3zJl34BHjQmuwhuFGlBwsfzGuyEppRKM4JRX1x+mXIvh
b200EYoU6dMzatDcMCYjyfW+6ln8r3ygPI5DWx7hJY0iGJY7HLMxDzLwex9QkrE+
VLphURP6GkELbf0H/cZ3jeSU8hcjlILbKSpz4CG0j2l9MO2EENHoTD4Dn+F7N0JS
RWpu6j9wqeSZc9QzI/rqBCenZh3vFMpxy5NQIvjZDPjAKBMNW0P+eO6WKtx+22mh
cHePO8qo2Ai/8ysNMaucn7xI9U+iKY5Ho+S71oqxvHWfzJ74ny4bERPgtBaa0vgW
ucoOBWO5m7xVj+9zoHOwnOsYV5TqtlSHaCI80O8YL480OZ69qcNBIxodFk/6uMJE
b6AmxOf58aPDGJUROT4k5FdzejkOdyxlAn1rTDSWjlN9tHDgP6UV+mZ6BZj1rkfK
v4vcoKOObBo8sgQ9WRTNov5UV/Cpnjm115233MWwpkFrcKN71Z/WZhBaJBKcHNNj
GOFSm3YOGwTU2lJ15CbMf1/nJHHk1ovUY/la4G+nxAR2EPi2bVWjiF+65ld1PED4
dWp6ndPKNT9f9b/VwEhfPy4X87OVUjbVEDnUGYHG1oba2aMk7vrDDvY3du/zhyt9
WiXk7nY0af/On//gy/fp8Ghfa0F4oL17A7RpExYsvigIxJYR0Y1D4juzlNzNzEMn
PG4QheuysNeTYTNbcgYfbZeQJZ4544I75p4DWYKQxZDXqmFq0hOQL7pCLwKeUtMP
TIFJXID07mrgSEQWbXP5zXXxiYuJ44t2XqeBVgLYGJEYaiDi9UnhGNxGcy1oB1UW
cRirKL0uN9mNRyi5yJFdqmGTUFtH0/Csjqd3TV17xMmOmtsqKQsO23SKr2KufR7G
g+0qr2pdhLW9Ve6keoTLSlhN/VdFYBr031T3Z3ngJ7Kbc1sMOmQ44vXA7kPDTu3j
qB5YpcHHkesIJPRI4wBipP5OMaxAZKg5SltMvcIqltAFl48nbxQ43M+UvMNPxWlG
r/utNLUqbq3gOVnnxV2Nub9Vj2F4pW3jQMEZnHjA0jULmArFqSVt2kZ6x55r9Fbk
vyKdtsqa4GIOSzDNKVcqM1T4tMQu+SMGjwySItnjv2zE2N7YGAZuCoQThMfaW/2f
RCRGCg3jI5dnVKqA/Wbg85ZVBbTIjNXyzpaoU9K+Jer11vOI05sExei/UGIFehNT
SZu0h23V9D2pMofz89CGNltevmccKG0MSSsaZh6/HD7S5qOBxrGPM2opOL/fvAb5
NjsIRrCEKm6P63w9jlSMoeusb8w9kxirJlCFgPTqvRncu/ACmVFP4aAlAoWNfHtT
RIbo97Fi0rJMOeZoF+oXFKHhtzma8JG07X/3/eo+XHdjCYJsM5DDeaU31YsKZMBs
SzvCn1yBtxqoMfEXXVCFqBZq/DcGf5ydEO45lQyBfhlJAnvj4mGb3fWbk6KGdUIF
DMX5fhdGHDS/VgWo0hAGqHfHnF0MkcNPvrtg/13Y1PvbU05Tg+Auo53e7VjYeH0j
/RaGvwN1XaUgXVe1A9yZbaUAadIoOmxAx1XuFcbpn37Bcb84nY3XgZMxg6vZho88
Jmy9k9d8v3nP7OoRvIATt9bH+lBiH6k/lkadbn4ZR7SMVHNzEmk4PCdCqSD+8J/o
sQz9KLYMp7Nh0pGYiTUky9ZQ5O9xAXSnvLDuU7IsHYwKLR0aTpnOiveQHSWbYQa+
8iA0W36BhHxhZw1QxzFpOR+wsVunTux77MUXWBWDzY+etX+xq7KbfBiZ9yBRzbdC
12pPCUsoM1I1tZCYX4cPqJDjsYpH8wbiihFG4tN1ihE0Gr6qvpCLEsGFxv5ME6zI
3E3T+v1W7Sg+IFgIOoCV6v/aNpld8XvgZVaI6+XgmA9e4jcql1PAm3eBXx1URncL
u0u5nCGB/+vpOaZOYuKPRugFGIbgyXTR4W55BpvFD1l4ZCeYx0IsdzTaAkfQOsmY
5k7DI3Kwi0NzZ7EWmcXmbDp9mieWrh/zxDGfSDxadOVWatZ+S0bAZ09SiAtjbVJr
A20Al9QIlSQZEf8HYn5ra1zhIrFGc+xnRzNywVeqnW2jvQu0Q/Ynuh+5olmfcJkd
/84e6BqZdYOWTgs6azp90rS2fF81kz1lB3EuXj5pGzrhs06wArqCh2Zhwpvn7oQg
9fAfCYYGVykTSBfc1uifKR+eTsIthFqS/cpMBmaf3o8yvdi0bCvvcnCV2BZ/+aJ2
EA6jtY//8BXuocU2n+Nm6rFp5rneOXLjg9KDCzKISHkIckhjEC5GwElP2VlkUoX4
GvS+8B8bPkoDJ7tEFE5Xj/I1J/uUt4RdLv9Gc1B7zkqedWUbDzhHqxHePcvvv5Cx
lIcMR5VcSk3zLf5o5XJ413xni04mRTxgK9vRE/zByXQ1kxXBkvQz60N8+Wl2LOPX
MdOCbluUQBGD7O3UBE9cc8+CGKO8JHgKkW4wu1WZufu24cXRBurVgVjoaOT4CzHs
i3OwZu4nQeUvf38DxTfQftErHWSR8TpgN6WYdJkq+S9Yvav88XdDoutlOGrkBznQ
54ZDjiJzQ64OEbG9KHk/BskhiZ1hznKFTq55PwQh5wAl4RHIgtTxV0guaMyXgJWV
WgMu2lTWLF9XaCBV+YlkrnCgo5oAuUWmpXgk2wMA/+cwU08Iw7OkdHC3X8aLJJGD
jmr5zWvTy94qMj9GknB1l92yPkZo799EojeWcQ88Sac/Piaei9nefPhjDrBKwmOe
6jqZoTnbs67atWQmUyoTSwO5uT9/o7dk9FCDVG4EYSHthIwzxuMHYm4CBXe01eQJ
IpslYWl9ifo0QVuR61bNdgfiWusXDPtwG+EqIT9zdn6dCQltjnQ6AQ2WOjD/mUz9
R/GAbORWmo0l4FK7pFaaxT63rSKim1NByFFM498il+yM5aLs02mG9M4c/r2aBgao
o0l+mZvNpV8ZEHqfs8LivkH10YqGIsKiU9j2610JGYgvopSDf1FaQXkHhCcQaY31
g2SVkBV0zAMpXZdGx+nn+HbDVw1UMWqqlLaUkCyYPVdHYqLcnzRUArQAQFqL+sUg
POKhD3IFkzAns8IQUhzrbhsOg2k17hq6RcLyH0sp9o8rBgHDgFteRQwzhq5jcx3m
/hHACINP9BIeDDpI89s7/gwz7pKzIr9u5nNt/FB1aLtHhVgWw79ljNKR3vEsMqkL
fS1SEh0cqTOIUcrJNt0tBCezRmR55OFfNCP27V9+umLNhciXWRAYJbDFSqvwYKWw
BDYbc2uPv8c6id6AvPc4QQQm0ywkVpDh/HVnNFotyxCJ79Ocdm4dFraliHjoABI1
LxPy/yUBLV5HDqDSqduM2b1rwltFY1hmEmpZJO0x/JUiAoKXOaPK0/DkVgRZlB9E
OfUcKfcsvnDzbLG9oJ/aW9tmLuIlGXTPrXE4sMT9MEWekxnsgu2gILD4jYn3dvtx
mSFi5fQQuB9qTMbbo3QH4NXgpnRq49JeLhWSf+PshE0c2vbRGYHlh0c6BBqSGd0C
ML8bIVHcLbsudxIdqIumGpIcoMM99Sf8678/OafLN3JyxBSLw3AG2V1ky0fIDwS5
k8M9uaPU9nYgHW80gGGgU4Oa9yaX3vLDEpPRvrljVSIrlmtIqezqm5o79mf6iS9f
37LRbDD0iwXtHJnhpwguMttFJhCw+FADVdkczyKd7xxUw0fE5uPfW6LyyEPMZUzh
382n1k8AyWuJxZYjskunYzOMlO7vr8oQCHE2QRm/3I9DcanXCJ3ouVxYVNlXjUCI
C4pgcP4ltTfghEvNI/HbhUnD+QutyrMRlO2Mg4om+caOVj0qiLe9VtnEFezof0vY
cgOJt1hlqmvUhOryClFNTU7MVV6x+A9831iSfXRzvrX3cvJJBdwvfJruGp61dXDW
wIEgLFeF3ocq5BK/Kxp0h5m7j2SJ7dgYdfWBQmlOpvbTT1B1fXKeaqXROzM2uGcA
a7SYggAU4LukE0iTWw982PAogNkbFoh+5WGK0Xpj0ts3ynBQTVTi55szTihTGSKk
hPeO+cO6Iju+z5nR6tTyZ9jmhEJABEcQn+FaJjiq+yzDBEVmBpBFfj+rMOUYolt3
kIEg9nFFOYppErq9r7yHImqDjjw6tRDL98Ult4DJo053HO44VfxSSnSo0unRiKYj
Wh7HL7eHre3gGIoTYE9drxaX3KkYTcP7vkJ7PHe8h+VY3NcfVtb3wNOTlE7avVPh
wEgje9kSjU8rDGI23UUFRnqi8bKO0xqB0KeSDXYac1xgpwde9KXqdtYmBPc7PGoA
mZXdgpnEl+QFG+ESb399V2dgJvIZAufspfeJ97WU+8qvFNX2o/Tw08yVI51WaRxv
+jST0ZEmKO2hkzJ6dRXVxPqw86kfK7cqsE/YzlouloFCzyU8Gu93m2I5xPC40CAv
bN7Sv8OhzyWLtGArv4JprP3Br8SKtRZnulojJeRcogaOe6SzLXWl3tG2intocsvy
Ugms3nYpFMqz7PpWPBWg/EJ6wqya9I1bYdOIwjfl5qM=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
aYx4MsCUWFE9Cjq88zj3CSHEGf+JHd4wGw/fto6m1Rd4doegSBYQ4iFDS1InM0Ic
VGxLH8CLCN1BPygdIUNbzGURbTN1fZCo/FfDP35tlN6RS01HlhBFdzGlD4Dl+kFz
If+2cAEvQS3XFZtog9C+h6VxUHTkcIPE/ABNw4+rr4AzYZyFve9PJSn+hOO+Lr0l
VlcQh+kq3Q1x3lSLX8pweOm6AJ93AfZyKdOpDMb3xaTNL53l7cEhNvxQUHmnXl+T
BaVWM3nJrtQxQ9JJ0ho+OF4s6et35dvGYYS1j9bV1dZf0Q+2H5ZW8dOspuX5TX6C
WKLuRMNHse7xUF/5lRG/Lg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9232 )
`pragma protect data_block
8FDV6sq3fTorKSVONnaWIITz+6QLFtWZI+cgWt/KPf/0YLS2raLJUjESZ4HF3c7s
VXPXE3doFYsbYhZGt6hSexJzhQe7O/d5i59u38ojnMqnnWnsAjB3aorzEkXusR+v
o/i4RsRRb+ZNbG4Dxnw7ZV6+ULa4DI5MEUAsyDHIAn9nFf6jrraJCZ/RdRcaGwTv
NJF1B+QkHJBAAXz41uBGytapUk9Nb2/gh5GffB1DLRGjwgED43gxpuWdpJRCzf1I
FwMU6I9zLAfbLN7Gxen6i4wRdaGLFbjPBnN4k7Os+3CVHAHLioV4o5NvqxNerp0J
UO/Efl358lcQ5OVJJ2UKLe5k4l2L8lVaVHdn6R+nuO370qgmnrmsXre/KolDvxkt
EygXs+v83pvGBLreuDdQ6WT899qol3ex47zzsJRpaeXmdWsFs/khhEO/PBpt6kIB
5fG6wVF9XI5QwwjM7y/Brm80qNnZf4hKQ2pJicfrQqBAHS29BwEmwodq0bYCWGog
2ly2Z3nPx0aEPjekInyLEJ1Qv0y6oZSlAwinzyITCMSz/VvDlZyxYYymSD+aCdW+
80Gj6Jzeu8F/czFcuNcm+16g9wyH1afTLM08xzh9MkywgHzOhLBKvay+Ieua7y20
suBbEwj1WF/bxOHnmIR+gtjhqao6Sq7Ds1HllWkvzUxM3j4J9mQlG0KV01i9ySu7
475e7AfEJ6igogf9XnLQzVZ1rLNoExVpq7EWZq7X8OZKAHoL0TtGxcKm/VxdJWaq
2IvdXmH1nSi+s4j4/b5XwG4rEgfJc74ScuhkbflyiqPaSc4tHI5v9cbKgt7N1aVI
o9+zll7pR6BIrdJUvxoCfRfQ/4jsWfYuUIXBtTFBDk06LAElPApiTWrLZOt02uGI
ot/CX9P3lBz3ASnSDJIWus9g1jn1LIEhwNDyFKVdNGVDsD4rzQ67nsOM4dqoE+cc
6YXfR/+kcGTV2AE/WRq0rOIJeVl4D1U8GoIhOURKRiRiBKxJ8MZDQZeUP6AnOBY/
dQzSUSnexYynsvagan9W9ZNtl+9GNBbUJi3aEJ1ajeFRHXu/ubFhMnV8vV6c/g1p
TgigaSvBhsk66jWhY1ooH3HofFcq4dwUxzjMmDL6Biof4OIEMxlzEue2Nlmm4/VU
/TulceFq2KO28+WK+mND09fDh8/2hFtGkHsU8jUdEcHyQc5d5Ys6Y0fsM5rWPk9Q
iL3OgouclzKRQG6vVbjvK1Nqlu6vU2KmMDtLHe4MTvagPLosdy6LSVCLGZQt33WC
jv81Oei/BLc0d+6s8CMtfSXt2o1iMW1OtR5/x+aYRIxygqMIsaeMpKeW8v6ZwX3m
tHyKqZfCSGSqn1V2SIN547papNtzZEoMNZI1hfmdk41RA7Wb99+LRL6QWPbU7xwP
HBQMJ/K4ZR/pORbjWmXN6kS55+YH9e2U5x5tGMT0VWrg6yojLfp4HBP3iDWXKGJO
cZgIpvrq9KX0gb+Vw586u5jABXbSM32Qr2GolUI/OxG8LP+BG8r85YY697ybnkl9
fR/HTTtZPtRGaYjmOdZ+zwD25eOgChk2dz4YOlzzVcwqRZln/5IiopBjUcL1b2WC
01i5zVLuhjvJL9bHHTSufrsvkdRCvZfONTseko7/NPNL8SQZhqd8ZNFpV3pd59GE
DxVC5DJTT4DvJie6hu4VW9Ty8MiyD52rrKNxxPq3msOUTUZQc4hQCjUWp4GqRWx+
Mtivo5G7UXWQEf93lQUM0mHsDG+73IOdiYmIG8WHqeHHGJnU3jSuDficX7BlAg5E
yCqSJTGc/olAb3cahUMOuMDumHVB4W4HyYz7hJMUKUCa9R4abSQ6wfsGqiMnz7xt
KV/qv1NxeKhc/SYy6y4pine8iDHOgnP3Kv39HoSxKTx1poPwJnzslmKWZ2jpjZSn
Mrz2T8JX0EPEytx0nenLdrfS5XV5MSQSMd7ovXB+XLQ8C6u4XzZgVs/75gF+7RN7
688w8QzUHntV0DPP2P1ItXF+ITkvYooLI3veqiHqWkDkxDUGSUoOjfwmWIUIOuGR
KCblbs+//E+j51SzXXqo3lDt2dp7MpvpkDorAsCebiAqOIzc3ri1oSW2ekfcRxN+
4hnAFupzjECykLf0kTfuZgjZ+h0fAu6BctCuIOeIXtTDQEQ+8DpO6ZfugIaep4SU
ElE39UIg9WnmWaAcTdQfODdSDea29VDt+YGNXZ8XyhibVijGirT0Ah6f1wjOiE5e
IkvD/Tytm+Fh99D7R8ORn0qc7NFfYJqux6MiYouLhWL8sjjUPJAUoviExPDiX6HW
pawP1ISkaQJ7lXYq+iULKjFKsZB10oHFgIDwdqBOxLXwRaUgHOc3lwyLLEO/ETwG
7yK6ujM51CQNHqapBNuY1WYaSVhcdQz+FtO1+rb2hLjALkm7Cw3M/1Nl9CnQ8Ctq
NQmeHsQbTnP6xyvdrx9KSR/NRJb2QIU/yTmAk1P/oKPvDy1LgAWNzox2zGoJO+1r
2oi1yKJjJ3rO3WkjPsVYskeqrobMs0QVUVbWWc0VJqH9LQK5K6Zq6wkQJ1bDM5BP
RL+USZCaS8HPlNhS4ovx5uz0m/9De7wpP2Mb6OF5Q95aKuBNXxYS1hzyP5A7D5S/
8c0YRI6yucW8zv+b8yNVGkFfiYJynszL/EQbr01qKFEusLsYBm/Ilzi8/c/5I9l8
3WphjNdvHL5WYbxtGb+gm0IxdoTQj19+OrcicjB28x4nGIo0ifl58e/wfJ1ICoVx
n2mYA9mmmt0Cw39B6DmhYM8r1dlxPmNqCHS11q40s6bg9yfbowxfy6sRl5jcdrg3
9ktPagu3I3GuIuCrx80ONi5pmDMq1vKILjerYP2t8cy3R175Hzcc60d3hNkCRUvS
aGXL1aWeBcDDusvif+9Q86+KHtFBYQrPS3e/LCUhSqvDVRlMeWH//XAd+8gzwxpr
2iNaJncROV2Ok8bRaejD7wEUJDfU5DvtYmXANwMXedmCE58lfgNEY3nNXk3VbrxT
vMTAIykhNg77yeNLLUoYCmV5vSUvJSMdm1Kk5S3o3tH0aUe2ASRFpdcqaWSGhhw6
QzgTDS/D3XNCis+uL79fv99FPyrM2z2v5Ji7n7E+/LLxcNAzQeAKHfs2icBiVlTS
RTgjSVNuKBLkn332oyCXxw/NHcBOdNpGK7Za0CmR4ya6uKoFidT7FHk0h/+qlZhe
Tutua5BKuPObsTiNLr09+D88X0aYIu/dhEtyvPaf1tsqzWZj34ZBt+zvSfqHcbMV
DaEwGfxfhzm+JcLiS5ivDu+6OSdDN3F0zeZeg+mu80MaZ2JLlkBcoXEcl1PrJZBA
rvMNdBPSFJ+WCBoNSZ8CRNbl3uiItRDzthOpsgp2EyS1oSVnKuqWmLPmIMhp9nil
tIYT3mPr3za0ZCh8WXR36V9bv6BRVskPsAVW3H5iXkrl61gardIEbEtfX2rETBFP
j1SkWgCxq8NqV2AAQOGrlIGINJQAV2qhEOB0txUu579NtOAY/qlsTGtCjmY7ody/
t2e7oJzWhY6QQWgItvns5MspjdPDzaUIMO7lpZxL1ZqDE2GUg1V6m9TqeJUNAmRT
7GSGdOm7uPNCVxHS8FJ3z+Il3l4gUgc4Ke2URYvp43cPJX4a4Z96i0U6IKxARfyx
T/GXhCXnqEPHBuZ4cVzSAfa6ReAZrCZVmFqcBcuJGnLaJ/D8wIUCSvhFPO95d/ku
song/DlLKSZla8CMmsWpnYA4+Pq6ajj4cPz9aOOsoqlV4nrGnP/0xduOgPvlmdDW
/apF7nHr8Pv+2yBMCT9/WORWyY43R5EfGgt3jBE7gzmJdDU9IHkBIVopA/mAZUvy
8YcjeECnRMmH9WlFT0RncIBXUPrjtkdgN+WXdjWlIs7gyxGNU9tHZwwH12zZxQwK
ZHI2N63uxVW4O6ZY3wGub/UtuEYmlZFwL3GWdf8auCL8h7Q/FdGRvT8gs+Zung4q
Dv4Vw7+hxw9XlCp57qukqK3npO06cJWe0zRR1lX0MzknyVRmu3xGZlCmI7m6ZlQu
tqIHFeGaP/rTFSUbeBycehRThP+BL+ypDxaXyg16hwf+pxMAfyTpEm9dNMczdBpF
eXQuIfE+IZogY33SAS8NSFZNrRoDbl1KjVF27LrFAEGiIe5SRHXW4+2FwKrOoNq6
4auJotPy5S8rq9AQ7L6WZsis1RbbxkK31S7l0pv16BlYs3WBFxbk+Cu0VZBcxaK6
7MQlCb07tLfLkTeCR7OL7av8R9cudy0/BXKhaxeCeKTE2xhGMeniPmaSWp/20GCp
mYHNONxnvRZ2/1GCuhauYwPNK15DJoUsR9Zzp8BdK/9gbwr6B1H5YU+Zo2BCpLCM
NuNhJgMSOzE/S5yMkcAG+CXCca4cac+wJpWNJPeXsm4ArAzlnbP4Cji34EOGkrvK
EniIq2FUEOhIzzEYzTakBSLA7rfoafhgGx59Ct3QnZQRYIKOVTkcXI540A/+wJXt
LKCuy55PvL18yeVdzPOczRQutMTILohRjZ2ijTFjA7o28KPlfMvCJgRRUsgZZ2Du
y/WocylJ7PVDSfZbAbdzEzdNUmwjTxUgoP530xlCBF1rKXsRra8zezTUwoLmwzLy
1+w2IqyvFE/Bf4eXsreG5InwIEkChznaITvyA2EE8kps3pnVvd47ppRxL83JmL1k
/Qso4G7Nu0sxhEEM/Gr8xc1Yff6ix7louwvRenYb8qVW5WAcUjbEXthiqjGYjR/9
KblcY0BXJG1nbmd/y7gbg3ZoLzVOLRgEk+1VMNLsKbNFoU5HRiixRJTZk06qI7Og
MvSaaJcypKOsuo+5M3JDdJet+fQX/giGpdeoWFe9R13KIoZ4ThQRjEExZupXvmY/
ab++rfx1VyZZdZhcO+Ws371ZhEu5ci9UVaFW1grD4pdDNK7XMT7yjIe4o9Vtqi+r
mtY6gGJCD2AOH9oEkO+SxZ+t5RAgRNvJx4SmS1CvjBY2yfn7cx3ixiZ3aeeZkRWn
xOesvBW1QGoo2S2Vn9B75a/KemH1Y62SF/EiZnNOx2uWGPbxoO5z5wG7nhY0/2v3
QGwcAnGXTHKdN+lWDi7erErD72ZbGJNFvaMmdoM0LAnUoe17MpRvgWXx3MUVO6U2
Cy67a/LjLp9AfjXjgYXI/sHsLqtE915DEnmzC6FlrWC0h4M0KwLKY+31OQpQIOsB
t5owFB5nRgYFrWpNBBa0BWLxyLs/FSgFj2f9eW9zlClRSexONEX8iKmvNh/FjAFM
1QabHDVuTzTOrjDryYM6cNxFJq7eaFZYtme7Q4jJLfuLHPVCdT0UmPriYUsoWU+/
yNQhtuHhQO0KOonOAS5iXMQoD8x3vKmSMuqrwqYROKXOdBN9DAHG2eVxDK5UYiKy
H2QpMz2tmj9pQ3yZZyE8lsBeL8dFjClagFUq92DGqfb9Jkcb1RwKV6cU+jmlo2zH
grzZq+tzEB8HfCe+6q3bSd+M39hZrMCzxyC2RtGUqeTps75uz3qRezTk5JD/Eeo4
QQpPjFvDRBLpiHz00BXl5wGQQYd98czzlkHqn67QkT2os3e+s4mAFHR3K3GRycoj
TaSfO4fpDjd7/Mcl/6k2Wa/z92X6UTlWiuskR7hAlFxUS3i0XvIYpkj4v1rRyecM
louwNatb5EVkUzalpqmZcUmNnST1Bg4gsCJTtJRo+BmVrxYMeWDnfE/laduqctsr
VgcagLGFU8890qMzEnDX9N4B9j1lk9XL7kH/cMS+utUTLQhZBnkqqyxsFF4/AtpN
ZfkNLaT+C4d+nBz4vrO1qMh2RuMdZcmrjbsLh9gV21/SiEinpC1hJVuui50gfaMI
oovI34/qyxxclmtqgz5jahv3sgPI1HDDGR4bPIXMcH/Wg8f380/95TyAWVStOqUy
j3+E051P/kMoLFEpJ98+Suu+JCGyaLFUJuZr2zAQCm9ptRzsf931upswZMWDBDWM
Dpao61iHK3u9RGX3U89yOMRO1KWZGsJ3ALHDs3hCNL5LDRdxDFfZm3n1bzVg1GGk
8/kQQb2KfmZjIcT1tjMCI2rOIVm3X/WxfCbq2Uodl+Fqc86qR7BzNlguk0oliUuu
1rm3pSMW6LHLVc0zaZ/Emx3jhLImI3IVL40EytDnBOMZmkYJk+msetWvSHH9WGAz
gcibhLU0HBrilXOgdNrJ0bfLXRCOoz93LL4cUfT6km5ZUeLKF++H+LFaVI+tJf6y
uNSeaioLHNXNl4avb6IIKGxAuWbuPy2BY08GI5zulHfw+aMyb6iLRI+zSTZc9ZN8
ndF32SoInjEtyh9oeOIgEcXouuD4W7+aolmav2I8p6GRlDqeb77+MFgg0ZzcUlsO
bSn1Px5+0EtwyO4C3w9taV9WMnZzZ435LB8GP5DoJR34ZDH0e/EHOZVA1ajb3s+l
PtxVYp9CQ7KwWcMncgZQgEARSv8Aa2sCx0t2rO/PW3su3OvDn/60BP2rrWq4j7cs
aHSCLMRorDroSPyGZm2miLpvPtqCcX2njwXi18oOVKGshmLXkhy2+a0LlVUP5441
MXKFen5go7SKsUT9Mk9WwjL6DS5eiN03rlG0FeRoUT1u+4PLc7+OyKPq4XVsoYS2
QaCn7wDQXhv+2pbKSgwZ8+qBbCXGVCpSAaQvFLGddlb+ZcjhtETURFy3Vpg0yhBw
HNeBrg18dprVuVzxM6OktlyTExVRjpw8o+1BWldKlldwEdOUXO3V4wKMPLWBHRhX
SykduovhxzU3BxdzbC+cRu/cRM8VBeB96cNeqVaJ+9sYX6j5a8MbDzTsrMaA5+PG
m2+mh/d8dVkivqYFry79nsTc6N8/W7+cKknWEII+Sm11fnk4LC+zbHgQp2nH5t4J
dg4zdU2KtT6rHmdvbxolt2yD5tqn/hQPCaBVRVHw1OZEksM88ESrs8avHvjOo6Mw
d4lJww7lbCGZQV+EVNJqu6AUU9pI/LDeI/yBI3PDfxpPXPR64YL0lcnF7QxloVXG
RFRFlD+kiTtXr4ri2AWh09cPOJD8eyDPHYSZM3am986qzKQ2Q6E+sQn4QOnIfrQT
P65qbhIAI+BiuTUDc/Hw8vT0ZlE5cird/T4SiongU5tAWNUxa7B0vSTM8y9iOlG7
gio8s3NBnypvR5TjLtvxpZV9kkgch6+1La7kbCZq1rDS3Tl5ZxUkhPCW7zRPN124
UjkPfIjcyH1sCnzlXafngVXkvIv6B84X3rFfNRyXQGftloH+6ABAhrFKFv8jSsRV
anHmtCiZpym7FI8E7J9WHCuTZSdyNHn2x09KXpQIrY0IuGcHSt8PRX3c/VxuSYrR
CMZqYTFYENBhsQnnJ0EWTjeknwyrtBeWqMf47kj+NjjoXf9ykFRTEzdkXOAniZXb
2z8hS+fNCieCviHSyxsVcbvQilteqNvh78gtdQxgsfdyNfLJNlh6+aIsl2oFSBL2
H3GZFp80GkR+W4ToextFRGOX3QLXWEdT/msQ6FQ1HTPfcJiPrumxG5YpnyVv9JFN
6CYwNkXDep78Eq+1V2zIE5OR1vhipSU3nmng5BW5ZDFH63xwKHBiojeLRc0Molid
HN2KH4C/FfEoEk0MPU4sq01QtyHYbCy4zlM1ogCaFuNKoyIVoY+I3J8uie7iBFd4
T3710aDBPP+J9YqGGX7qzHsa/7eM3fwYzaDr/NTpCgnUhfudiE2wsg0D+45vCzjh
/G9z/A7ewikw6NdIs6HSyYXMrQwHfFYwPIfRRIOKNtd4Ojd51dxK77d2/UybeEGX
l9IiBDhmJUZmabo06bWUAStDhmTw2z+nJxqHR1krR5eA+1wWXy0c+G3bq6cCFGXJ
kKILlfjX6M4X+X/AVmylhFGfDK1pYjp67sennG+TDZGymKSix/518Np1OyajiAQf
untya9f6SBf43Q/LSbtORcJRAxUor2afImcvq3L6OlO0y+cjw88Iww/GXI7BAw/g
FhdFisU9iVy+bXFqshHUnWdfV8XV/PyDM/6a518XznvTKByfVkbymEV03QbeWyJu
8/OVXp50vr++enD/z18XamZdYWw+b+f/jzkjy/opB65qbCfXg7RmrIAE/AJCk2tP
KpPe7mrvg1g9AHlW8FJNG7b4fusrcwPTVWhpCY59Jl6U8xBAuokqfXv6KAM2toOD
mmMPBimywVaj5zRqIQIm7S7wKQgAoAb1UZ0dFMRgpFuVU8p5m2bN3QfCKO7Cjgj0
pbwO/5Kdf1i0LV4gFnl6anVmCh8xSmj+6796T0ZSAwHDaOFkYUvgkJNeeLxggcLg
a+CgBwp1TG9qDyhGXphN5bxy6vSO5H4QPGxyY16vyNLhdVRC1oVGWzPQ+S424T+n
L675f8OBMXnYDm5F1aHBwFpvLWjpp6UIWFZlAwRTXbRd8EVK0e8/GKwcnnVEe0ZW
AcQcCoDLm5wyj3mjYXp3em/0aFeYKA+QZrOW4z7ibdB+iCNNtsC2H6hdNgDN4XwO
ORL+sgoxWlBH/KyMVop97+rDCZR0sOcDLDlbbLqr3MOt6RXmVq0C8agNQxN4PDrv
y+URFxABaGhOwzWOhvf9wIjZtxIG/Eib4x4nVKDAJhmgWFqaRJVxtudbk9vXX8kv
W2QtFSxWW0VWGCrWII3mHXDwIlp0UAbRf2FTs+a6pau2wByQPi2GwYoBbEZYKddr
TrLMDHJqUPjv9i/BZJBjWSegI6Nj/np/SQN46kwIOE/4tP1AuNxN4MSGeF7j51O0
8T3a7knWREv6etlmI9Y45fg56jQbx/wqS/H0XZxXAT7cEeqybR9Xm+YbxK4FLjT7
c7TmEabh81mwpaR9036sOLidVz4yc1/zlFvp6yDRgoWhfqyH8CfYQHseV3pLSHSZ
+gtgobNW2Qa3NyK0aIt/ZO74F8gFKsw9YvHNQDdufZvGNGhrLIua+Kw5qfebp+So
Y+Ty4d+Q3ZvxCYhp7lsTNfhveWDW3auAd8Fyo6/w4irjNyW8uVz1UqOTnnlgJfSy
FkqyMaFXxcPL1RAgwRaTWuJTywJ1pkwM+HeLktw9GWILhXzZvGLNFefvdgtUlPFW
LYT9WIz/5WA4OnmeBN2eKLWgY9pTbIchxn0rCpHfCWxpENWvmwYm2NpBdXFKiogZ
PNjA8fJ1RLUoEsynh1oVwLOMHYDVBkHhReNp+XSd4vHhSVnwMhiOWZfgBcWX4HUD
8l4n6HzV1wkSBsFt4dBkfj5aWXrp5HoYA2fUYIvme37GuosBwyIZKe99ohJhg5Kn
1VTqUAx5PQnJpHBRK3ZmGH2fc5GVZ1oBBQDkf3oHtLlCgqyIJnb6uws6qqKtG+jk
df85m9b7hznqrZFBJHYL7r68UrOiqKIlBzr797bRjCi7WlSugb78t1PhmJSBHPYH
oAcLOWJSwvDF22XYQXN+QFnQBmhh9mI+QOZxPJ6AZ03Ds4UYFLXBa1thIknWScsB
iFY10EABwEmAqjzwaZ42BmZKnNRzMvvoVJlTS60pnpXyGXrPJq89Ea8FwGGqC4Ml
de2DNjNpPOGQn81PwBpWHBwb7oe5ZUQQKvGrvKu9tHPJaF7xUQDlWP5PIX1uDu4j
hY3QXSLZYKzXENgO2cpsMjriWAkREqKwFPknfso6JgOYL8axxTxNVL5GwoZZeTHK
QmZw1l+vp7etLwbAWZEiebtSl3Zt4jIjJ3s/j29cShaPclSqcBTd+MMTpAAEaFlt
nvF40z8v+PVUDPZx/SA8ismf61NcG+kFp+KtzmxNG09u9F3tgtCkTqmYbaXeSPz8
YMgzIpNqkHh/bE/IqhzLlHuSOC22kJoqyALBqpLI5BYZ3s8dg5ze3eNACW0HyuAn
V5bcVOhd1BV9bXykWnIJAipqxVoGSbW7HC5Wv2ByUgzJ+G/HemuV7/G+6YF994MB
35NP2UjxlIuVcX7Yz5OwLYhiKC9r8+War4GBuizLBinVRuTWi6kBqUWg8KQbTYCE
eE6iyViNdT/r8vy3vRb0da5ZnIaGPCXnSNphSd8b8WXhn/7zcNVZK2lyR5QPST0i
5xoqBr/1GMpJZGjaBSLZgQlcxs2k0qFCbJDcXySEH6macnjsYX+/i/pXfN/ir+An
s4QspUOA78dEo++EeFwLRgKr7Rrv4sV79yi1wQtffwuKRqXXWgxvLtuwN5+ekLnD
Q+zmhLMRD+2HGN20jEjxK2NXOJAlsPZo0hC31aHBWEwZVuOe/O9GhjPNZIFJigqg
Wj4INqvDKM1PY0SXTictyp6QrMnOa+IZJPLJJeSd7adklG49pmuaeT1RrudTiSo5
5rgLF2Hf14ipjn+Zz5olE7OUXVzIKuMgNdydoYzaNhgmWacI0p8UurmuFpmtVqdP
zLOILylPL2uX1+a0WX6b5zzSo1yTxBWON8MLnrixOmPWxahjtmnQTb3rr+q+GwO0
zGocznmxmyJ024DO8L00XDn1d/oXywbGMIjLEKu+SC0j4YdgkLyIIRtwuoNRrmzf
I/PxeAW7pjt9y7NhoLC/VtlNLZsvxpBc+KqJw7zcRVBEuAFpa+6YRXNbKAuuPL29
M3s74Nkag95F9FE81HsdP5wX6FtcJqaILqrQrIkYE4DtV4fKfQgcGh/usnVS3u7h
QKIKq5KAHJEOyPo+DGVdrBqc95/6e5feXu/A1CuJTmgn632jCgERt47EeAD6J7XW
k+AdSTIcSi0cpEPDsGDlg7RNbmPLZ7+Un+WvR+e3PWucMCTHBLiO/N1gZYMW+hxB
EAPaPRbrz1Tibs+iI/KjAqn2RlxtgAOknKI9Jl9laXwtLu87j1K+crMCSUH4UHYq
SDFA0G02aydrN8PjxlowXXBSMly11JVVDdpV7ki6VLJ+BpmlkFxXhu/Is0JgCUFI
5pxJKpAZBn5WSwfRxSBWKH98eTZnCgzKa/0YtcAYjxbNmO1xobm2cpSfgrt4qSYp
yK9eKUsTKArSWutWdyzS6vVrFR81lDGnOXagdjV9kV/UmNeZAwed8Dncp5dvb1Ro
1gbF75211iIh/shFneWcOjcV/pJH6URKfna7c3Gy4YIhAjxTPRCp0emEIn+svjL4
2Wnrw3PTz9OS7NGpmV/KjqpUom+2kQVM3LgQ8lGcdujdKGCr5NPwawq7XrxwxhCb
kkQ4Xw86DobeZfQku15oWlwSLY6gGnNokUzcfw6nvSpAizByyR0uMHayEApnh19E
ke/S2CGIHbodeNhCvnhBy61stlS8WMt6VbOk2XnrCw2kvL11raw0UHmegRsO/MCE
tHmYl1Bh205wK93pkDQH+UhZGBXtlIjCHiTYImZOhGykrzJpdQ9lmgH/MXOk7o3N
NHcCv5TeMex7aEqOf/TruyV7bKbQ2gIL0VvccHh9zslmTTcWNpy9/nLIXZS4dlIz
rVJb1AcLs/unmNioLPJ1HNHmekdc+BLRvlLGm9ml2/kWF2A5PDV/1oMb+733zUbr
MR53ITf/iThZbZwJ8I8BFLnKwylbHoBn5cjya2RM6IHuBoWHGuT82PV69zOWgO/7
JLRfmvv6sYZP8aZuUK3LoYwoI6zMB8+pS8FqW9NL4ssjTD0cOqnaJaj65xICElSB
pWk7yu4gQdmuZpv1GHr0te9Q8MkDzErsg+lJomFLSUUSH2fzxQlBpaROdQqPFlOd
miKh+FmyWY384Bn/HYFpHgVW6dTg8yLDmcY6fs5ezG7ZGJj1csmmzjX7RwDdOZg1
USiEtyS4/yF5RJji8tOQmpoH5d/dKsbu+8QYoWrTTnAWd1fRjBmm13Kl+qKjhn0i
PZO7dCyeUMRHNYJuxyGZ/QqMN0hbhFnWe2soeHJ2OM0GK8gmPcSPQcpkR6JMHHo8
Y9MLIZL6hyWUzgII2XBHiG9d43QCRowP6EP5n84QidSOWNrJVUL9iGo+ke8WjQQw
o5KYOqVC7ZD7wMAKsKrqUdLvzT/kqOB3wGEj0zeIXX+mnP2jN3DNYdm/14nWZ/n5
tfXnbk0OWtRChj6JvwgMRZm7xcjxkuKIlsomvDw+qhf910ztYC8Z5YY/mpz81H6Y
2pki7CxHjtqhjeTqtUC1AJDrHSnWTut6QtXCueR5Y80fdAx7GPpQO/fgkR0J/Az3
SDFYFliAmtYQBvRnjVqksfyCDP4FIjJRPfdThPu1DOrZkWTd8nCHM5/GpaakiSRk
7o7x+H0pLliuWAeWvDMFgJUP+NtP6XO2JXHdZblWw/aWhXqTVfd8nyrncOOlL8By
iEv1NDp+t84+IPfBPL6KsQS+tOPgocFS8uZTifNMydWZHhuhTLeHJoCkSq8j4UcE
GnD/rSEeRvs0gw4RqRsOut23NWd79zlbz/ulfe2QtI8Hc4lbJZrwb33JmAhJGTD+
O7wh+NRJvw6V54LNM3DElQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
iwClglTMTX9ykJpsES30VMAhe3uL45aufPdCAVoAKPFXMJWGz8BrmIYUdM0y8EMR
uYiwyhNNVO6RyeXbxbRs9FE+kftzTcBDNNYN8pu0NH97VPLgedsG8YiiscvRo5Z6
xdxCghQrUW03CcmTx54A3XxPS7KkhaolTqgJcEr1L+b3ltZQfU2Afk0M67EuRI8Q
xCNgc9OoDOrTlD+SJ6ZJ0SJgeQuccnk1AIuOcYofY82D1Te6Z04Vvqkm5GAXNtFP
JX9IzbrD/qbPcxTXFuA7AbTG7LT4l22iihjot9ntIVQxIuA5HqoMAVsxRwqPuAW1
nZFTlJNF4MJJ7aoXRqsfbg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14640 )
`pragma protect data_block
T/D/a007bz6JUAGBf/LZ3XyyC/vp/vDMYyDOJ80NEE9WqoEHXpbih9FJAiHtXOBp
uGwp5SC8dpAw7TPj/mCXXNGzz+OCn8aOJs2p8iI/5Ega33N+xUv+zUHN8LtuwKV5
5T2NreTdx5X+huPSI6umxJgUE7sXCO8XhTF+PxQjeMNC9HW5Qe2aQ0PxO50KyOPz
sRsHDV0UDsV4PHKUHrGwngztMd2WSErLwzdev/8gszCqmUg8SA/ho5+JEeW2AcqP
/MNHGF5RRjoIaHhv10dHwrLclO8EVjwhiH0+jcfH8yvz+DxjIicVIp7jxG9QyGPT
WB8VI0aVR6P9qcZtQWiK7HFm9EQeH3VJbTFPa8I6iYpbeR9a/a9g4jaxDQykXlTH
s25RI3uNH5moa8GeQVMZoAllYyKqyZ3iIiE/1iMympXmjVForiVWO4FN4tl14BIa
tolM13saZOp6mhEryoGKFs8ACCyul/sBpCKs0gvbAN93Xrsx1A/VgiM9Om4gfTiW
TIpgWycC/Kc/OHS75Kf5CWgiVMFNBe2ndM5kRr46Es0YesOxri77lzqSreb3Y9Be
0HOM0cUcEmAifIyfRxPKwO8NqzyjrMoNAioAW9x6NNAZ4Z2iw1RuRoi+r8SHJrpm
VDWk4KN++2jaSLYi/8cH9GVuq6BqeeF2pyidiECJEP1BTb5IuUrXPHy52jNrUUrd
2n1GL+5qtY5NXwJ9LKmJS0O88wZ5QjAsFgJxATGW54LcUGEsoRJwHDb6UU6nnKOI
4Xtt9vkym9rCEBDaHzzBag5NC/8YSQL1yEQnNZdSOr0GW5hyN1GQeQzeyopmAca1
lW1mCA6zq7VzSaZFYielOMUCtVs2NzKpRWz5q1hq7UVbCEL7gW9/m49AThXlK1+I
XQ327iB0kvob9yjj1zTDLuRPmBr9IgNg3ujzyMOk6nKwsmZGBPkxYZozQWNIuUYZ
fGB1aun/gXV519XvUJfKE4wKtnxl7SGlZUQ+8CWxOuerEJPe/wN0zne64G5+SAUg
1EV7j6LvowpyZwA1hi99CL7KZMlxzto1/qJosNldzlBhV6rPzSeNizBCFTQVhXVx
WNkqZHlWkKAtZbvK8UPzDa3SUxP5JHuNH1QF2MKwOzf4pzKal7x7iNkyEotyK0zq
k9zDuFjERfX1teTu2uE4fn6lpnE378vAs+qQV3BePPzcgvB05eoycLUQgu0G5WDL
TzV/RrEyMbViyZds9akB/0bTOl4obn58qB6HA/+quwZH+PlaxUsADy7GcEPLMevK
wKo8MfL/6zTCzGQYXYc77cp7rZZWIqwxejB76XCeQd8xKnFw+HpTNwidxxXlxvfq
Hp66+ittwHw3Al4QqO/OITRiRF8tG7HAjTjX3SsHPMv52FNiCPHzbX+Wy4d/3hkY
PYNs0zYUtYECRRUa+oVqS7/KGIzNPNEsFcmaCCdVbimqhpgTHncJ5jlpzNatTgdt
kay6wr6sDRZiPcKFnU8pwIxl1+RuWHfO4GMJ60QQOk+GKGY4/vojBj3FPYKYkIE6
0DfW8dMzdvMTFCFhwyVvJFulPxyShGlFZqPoaoOY8tI1JonF3lqJuQ3So4iQoy5d
wYQtJW8Ophfo19z3pHuvw12yvWiMtMBU9vbl9Egj6S8+Xee25VCq+jBdS4qhoxDq
3QpIbNAmSnbJfErdUWWWft8xKj5H0tLWJ6/ktH2DMqmRfJkBLZCRtwYZ+T/G7L37
5w8QHCnt5qK7KRrwlITyPHLD+ebv30+y4GVjtGfzohDkqLP/ASkj5DHjlJLo6dx1
EgqbA/c5b9NZqbzR0hk9n+P+lsguLK/9vaFULqC/jQfFRr4ojo4HQTqrSDnXtqUH
3YHek6x6eDTZubRRh8QNBKHgmklJnqVVU0Hk0gayiBOAlMIHAquNhtstZMYolNUL
6OmRjMTDMgpSi0AwldV6ieFVKZoKfsPw7AwkKnFuJTbGUsmI6Nq3lckuvactNLnx
hFTAMvRKA9/yXNtxUObD9V0EK4Fk35/XHrnZIX5SJsKX3zvY+5tbYVQl9qcYr3vK
eHu+t8gg1YekuS88/rsN+GQZDsD3G4wGN7VRMECeugHbADcU0xAa94dGK3R4FQ3R
dxD8GsTfbcIs+Brv518t4zXhgEMQkDuaL9wFNVa5/V3kVO5eqPoC4NaUH6EGKqTQ
TDcUdRWYhQN0FiODCManuixKfWGZiJ+Atv5ZDPKmZu2XnZkfJzXcm19uSpPdc40x
zXzCac4Zp3mKR+hJN6tOhnhQayxhxx4cfUNNHCwvqWY05QCsBRbUeiG4y+RCTCie
SBHUtx7nE8R2geLnH0IaxHEHiNzLr8KyAaUnHu2aecsBcrsUvQJdHGytn3jy9u0i
XpgI5l5KcJG1+XfCy30c8IxbLMejqbhXhUT0M2OFiL8yBz7v64ctuxcFD6wNrQm3
a/uB30M6IXo8bMuC/O8TP2lSc5qvoLSJOkqQXs1ARb0R62Aa7C9MorTsgQv10HHo
+prFwmmCy/OugnfiPNfqYygaOdmOFw44kcc1W7h58msPYUSmKyf4n2EM+PfoRktA
UC6s2haq+Exyi9Kv5Yj1foB7LmHw5M8izZedt0dn5+4WEqKHkxkaFrDi41UYTRmn
eBwYBwNby065mshU+SCkBmIy64HD5CfhGkXNZc6e4TXgWWRpWt5q82a7OALXTJtN
42evjZd7eR/j7OiMBNieeDTB2nhcAk9ueohJ7XsrUye98ZnNxG00DQgz4wMoBdmO
0wK/sQwSjvyBleA60l7SnOroFz3tPUl05awLlVOxU//Q+zkz+PZZOkAFGwUzxOSt
rZM0iWB1m5tR+wWKg2zgruWb/TTWRZsin2l7m+r2roLJMSqXHAd2IteFAZMQC2Am
D+1XVdSIYIqHg8bC5qoIoyB+iBckbnMfGZ8NnTLnleBAzFpNAet49HUojyteABFL
99s/0W6KLC5IY3ZcdmsP46mwf4LvfCtx14esZFWO8nyvn5GgkeX9yvH7+q71c9uG
vL09kfJgxNSsu3ICmceAnrzOxD8uUplQTdzdjkJ0AoFpHasVm9EpOkpPei9Df0/m
4QSekRsDXZuDbxSW1juUOlv/LHD/wNTmevmmlwx7ndlfzREzH35qUJw4iwSn18t0
l19zZ009Dpc8+BBLh3J9oWDA/hgzrsU9etHqdyFMUoEcJBRoJwmTXJRGBnLo8i5A
mFxvUKIz4SrLVI3mzymdM8iyUhMrZ32AWDEr98s81C6xJrIRekLy4i8ucTKyA0MJ
L52RHF+W4qlFSoXMrDQT6h2+TWKk5v5eKBZpTB4y5ZqAQ3h2xDMwLMK+lVzUgihy
3+PS743R9w9nYK1nysKJ9wEVoGDoX0ID0UFAyiolAwUTiDlIZi6y1oLc0ms+IcM3
UO7UifbvYZ/ksD0mnCKp7tBCHKDRekqjoFFUdAJffTy2Udk2myQ8omDoQFfyyeiG
5A3FcIGDDQ/DpZv2ABTxMmNFJH6gjvz7f381Nd2eNnak3O7jKO5yiBCEwRQtQoJ1
D71dnYmx2mN38lko/U/lppDsF8Zh4ovJW31WC61jJUR7OLxApcATUhG0BHzfHLfl
6E4pP6wzX0+3KYOnvcw6vqCQo81Ol83o39StrPe7in5VeiIKNmn2bDRnUWgygQgW
oLaYS2Hw5n7Jvg5nzIOxLv+4x2WpqT973m0TkP8iLThnhCYJ32QkIJbuVMZtsT+q
qGwue8+Jd7rSV6z5cKLAScCgCPo3wolsQ2CQX7VzbaJ399nWoYcHAsbIVBjz4lXT
uCsv7XOymeh5QguYOXqcHwHsjFu+mT5HkqT+SC1IchfGvW78zhMPVj4RyA07VLd3
gJ1+Up9W9GWzuY+hQlCKMuhuJcoPwu91LBMIelPDz1k9A5XzAjZKo5E2511q7qFI
bmjj9g1Bqoj72cdVKlU3O7WvOQNMk2ZvusD+SkynfGwo+3NSC4iLPGraVa/72fbv
T8D7ZmcE0W84YChkoWq+MJ3SOOY3IT6fjEWXl8Q854k+27mzvKMGl4eSQo+66xKT
h5Lq4aEyuCufISL0la/e6UuC3tHfXTPSFnvzEKM7PCDQNWdjm3u5yy/dMIb8vWHj
yN6m3QdvwNOBFvE3Va1pn4JhlbENzmGTp955KX7DnB2/lT8ZtOvPqHs1TxcedaQi
8haCFvK3TYAuP6nYxNQtxVUnuIB/0lTkJSYj3BcsTYdoTv3zdYyoKCognZOyzENO
9OpYz4R8ad/Irx3qHeYAdL2TUAiuYE3JPIwjq5YV8Fsi7O3ppKbg74IHCPCfK0C1
2kBXvBExVXbQLxD4pJfYkknz4Ff6Bq7A8p1P1rvVO8/gllpZ/izK93Ef06ekQL3L
z5Ff15OHqVxZAQo+bd6x+lHbE0Grkeo0sPYcAB4oeDsl2hkiFUZfFh3woeCqpO3C
jHEGK+E3dAR2MoCdsdfGltRzgTbFNKtUD3H3Gpa3QX6iQBpTamR++OtAvMLtRPxl
t+t8JidoEuVWJwS+HDZryWoxiqyanFtfavWqCnSb5zAXzDdIdsNHm6u1kSxGD6LK
wIaqgkrSLJ0IwaBeKSZwGQ5qtRt+QxqnE2+6BpBRBUmrVSszBEa+8kgC8Khet8Yv
pOJ4Qr6wrvVCZz60/TgSqEcBlvV4Fk5VpNtF4F/96oWYdNEUoF0s0V8fWIqD2Tmu
x5wmBA87K/nwWmPidoqzaWNirSf9hXWE6LNe0c7Jk3fxPSGDQ2FNZY9pNCcSsc+T
B3TWq87LyNd5IOx0BC2BmxDIm3b8aLIFe7a8dRTtPXog7FlHGOr/O0yr27+nWOrQ
wfRSnYXsXrKePvoUFDjb8/W36kFu/uEgNXe2weXFFbSszZJyQdljGksAu9/+2M3m
Zghu1nRbgh1CKveU/I21MzjGcCMfUoV0HOSUknKvUxnSZht1bw/fYKjKfpDjJb5N
6pOLJyFTZJRMXwMzX6u8xDoBIwcdwbFmHjwKLFv03B24h/48Ja9JfpN/a1dCzrD+
5QgWps/kolKbgmTVABYChwd4FT5YqFRQSGz5kcSMYl4gKhN+AosyQ+EMiwKScODu
xdBsdfgFCIC1zFV7DnwcXwmTsIwVLxi2HXH8PWFUAXH9NKjIhiXq+7k3Tvc4PmLD
v6x4/5TLbLORiqERNtJWEPwQeVnRHvp6rG1QVqftM6tFkojnWU2dMZVy1jZh/mE5
kYiw9n4MBPO6PyVi9SQ1iA65H4vkO1cTUDbJ5xxtRLMNDwkquz0PNr0ZzS1/FrKs
XfPeYrXfv6a4jdwvnjOUKvfjBliiUyWjE0Ea+Xo1Dv0V4l4vYjFfIDg7v+E7D2pd
j08oCpv3wIHRTfazQuA6g0esHrO8nxAqSOy2KPFGUgamfgSWZ7+HMw10Ppgsje54
EeRSQkvsEenBUvODGc15b4ACi1PSz4ljGABRv2hhlRDvB4dYrhFjqokHsH0Y2d7V
8lx8XXHH99lK0mrF3/PDbSrwNSppOpmh2LQjrszFDjj/UzxWnLlLxSPLyW2kIfud
FjpO8KhRyW+/YeVydXmVxqgILkvP7oFZ5KlvDGKG2nDf6+fYnXMaWmQNCI6ZwXQH
bgv32sKxsIV7G5EBEHI9+gr89uIBlwSdDKyPDXhyJP8LLtkovvj+6vBrV7eesYtt
B7s2aS8LJFUFJ21ZzZp02KjUDAGm/WQ0K0bi9gqgSDQKsd3LeJ/XbsZZax0dwUK7
9OBuBK3/8Fv+K6n0zjy+Cu46zcfCXaVcjwGq/H/jg+NHttfA5Gd/NFaxtgc4TYYh
M9AjeyBWKX+9YxLH9t3VVvTefOBULYkfAW2ZeRPSTWFNRatYrjv9FCkXaV6YOd3j
rbBAZ4Ge5gUxCOLObd5/rlmP5+pnYybwhfaq48xOqdJ7LLocd3qkcFdD8Vweqx2R
Z9Pni39KPEGnlMI+xjMSFH0lzOsNaDGSFAXvSnAVIOQ5f8dxFWvqTDS4vXDwqOSi
upI4cAkNDG+fjiTLqeOCgmwYEQvc72PC8l6wD48k6SX+rAbwYtjl4xocbbX6kIlR
ebuj9hW0WMe80OGAKRpkXQTEseEkKLxzd5sm4Y/2cMWhRDa2jl/WUR1BmXhBzQBy
Zm1N8MY9PHY+p+My7LiqPtQbtvxXciBSWAy066R7AzREQLTawWOhcMBOM4WefvNT
ktjrEBefQUS5MmWPDNS2MFp+5HbV1ZC+lLzeMJAAC6OelCdf6WCZfjJQj+qCxyB3
gSK4erqF8tBefi0ApsV+P98yWQ6LpuEc3Y1pNqqXfLHc0GubZhx0tYqa6Xf90Tmx
pCVNIqQX0DGU0PlH4bk/XdwVuo9PPXgsTaWUrmLMyOeJzm3+SChhME/YNFU4LtS/
j12MxudvVxITGIpmndg+UHYfDYVJ3+QoBhJDNhz5K5k2RmPhKvudh6qYD6HeGPGq
cSP/1kczYK4SUaQ5u/PxiH7U+fwndPXSqQsE82TDUG6USo39VJNovQyImzM2pmeH
PETw6jCBQafi713OtQytbduNlSh1zn/mbF5JFUnABbkRVzC+IAHHpxNAh5Oap1k2
bXJLwNEFlxps1UlsZyzdkSYAZiz+zCRyny/uSQb/fcBkLSZNhy5xHHKEzqIibW18
wAQ5ImpS7Q3JeHwKQ4ZWylq+MVlA28L9fOT2BGboJTiM6GXa0XsjJy3jDHp9dEgg
CpANe57+/IRCvvnoYSPCes4AgUNYUq6IxDjW8EGqPJdTEli6RtTFmDSI9OEOau1L
j7zMrAt/BTLD4FYJKeFfqkYMH3luM5Ob1X7c5apb4QVRdgymzymEUKLWpoasPW1h
REXJ85vGA+5mDpY3znvpABO2LtE2kQKlrLhukTq0NcPm0DpOXEO+wJWHXhK6Pxkg
gS5LSNtDeTxm0DXuUWIb+qZKrR1V0uaCjOD7mRryv7nc+76HnH30HY0kR7Vn6e0x
oAY8uNTrtOYbEwCm1E6Lx0WsqhknZqcSU0LdqUbZq/qpu7uaLcaDyp6Jr7K147y/
4+ht70ouciuT/hndiredW2DS9y+YFjHz/FCDRvJJGsTEg+kPuE/lietnjKU/HPDZ
bz8bVI/IkCUBt3/bKkIwEat+joBFV4OuUIW8S3DnHNrBR6Inn7Anpe/3NlDtZTeh
z8ZLt+Xy1C8fuChV7nlkveM1QNAal2Wwv2NF4H57NwBYWZ8Licuz96VnFCniw4s/
PsBKqpnB2AzCTzbJKeEXi5ppVo9f8PnAPliXl807dgBtLxZK8YgzjLUgwxsx0hOX
v52uK2PKtf1Fms87xmHYcTRcqrDlZE9IPKZY/VtmukYoD0MQQ25pdTpJILH/lv58
ktQEbDU/YzSc8eSTyRhb2Uym0wEDI3Axpu2l41Bie2USxWwCwpewF3vn6hbpLa97
gWJL9yxuobdRIkL72rS53VvsDe3UKgRkrpCMdrvgxrHa5YjX121cZ5uwj0qZXKL9
1+G/o0cdY7e9WJB68y/OI+VVsmRRnLS5NzeJOHOfjLFET2sbsDgDw3x/gQ2TUgSG
Pb4uqU8jh09ZnmFAUWeb6E3UsFCDAI/yC2LWxLs2GRHLSZYZxxd0k8lHoGzkswe4
g11NuK+q4Fh1FEmj4w/YCf/E7MaBr5U8JjyS7Gko7VpIWRInhJYIgb2SL1jNnhE5
Pq+mZ4ckPKmnjEUnHauLudRmTK+GnGmFsci/+y2pX+wVthcd5IdFRE2NxRWZLC/+
w9ODYcaiFPE129dDuKYn7CEKThO33I0pPkfDp98e+V6UsbTMTY3m8euyv7aedOqQ
zCJSzNK1OhayGNTcb7MG1lMWHnsobcO2SN2wYFffeXq2puGaCQbvCEFJUYw7x+v/
b9sdGXDUlwATK7NcLP0V3qqPEPE+MLtwCoY1l8cNGYx1v8bdjNDzgNc1wG4ZpUb1
hqODCIrYbr7pUDbGb9AzBBC9vB+z08V4zO0N/dcwsU3L/H0YZygebVpPV7YkrKXc
+oZFwy42s4MuxmDSPpsWAZy3L6KUjXzulgsKLJsYqi8wV43gH90NDXXc2dYobjGJ
Ho9d2RgV7J3ZuYgo4wpm7pcE75Q/0f5v12/auWcmLRc4CIKh+Pyer6yY5rRg2qBR
fhGig9KDmjxFmBAPbaBhpUxEtE16F8hdKxIU4wRfCKVexwTnGcF/n9NGYDhZu0BE
9D6QWMIkI1n2jkA+5ZIFxJyUpqB9IKsIYInEGaRlWxG3lBl/iH3hjJiqP6t8SEiJ
7pVUbDnGfFalr8PQeX9h8EJ3yn2iXrFWAuf/TPkd2l0V/s3JxY4wJGA6ndkvzFjZ
NNbxZqqMybX3RiNjOKlEbK49rc7zylbrGp9ScVZU1d15TykszPVupglrqm2ockVD
Pjce3MLSo1d5f9Yk0rxBGctM42YIfXe4dTR/y36IFYZSgb40THt98H1/sw6sEkCN
klUvgZrj0Cd1IILEdJ+bK/zGKI3n0NCEJwQu8Cv9qCXjdFVoJO+MqEpJwdMcHkD3
F1rbcICFQ6XJCYnb5+kbW+FYU49ITYsUaax91REBNN+PFSHDOYlv5PlZ7AOdPr6Z
xvQBtyJUmK185qQTg9NA4RmPyJNBarBbH1pISV27yITEe7fN1ZG9mnyfIGxPvRiu
WRejmdwjtFe5g+Sle9SSQrsfHPOYirMatXySv3uzosh55Eg/zHZEFUzRzzJXu7Ql
ww3keaCi/7zjlY5sf4t2WB8Z2hlYLULgED6Y/VVmRxXfyMS5L3ZHEC9zxIsJVOlF
zQXl4Qd9BDU1AvVIUhLLc5SUDfaxtYbrzCcl7C+V3Fc9etWtPTamIZ/nrf4SINlu
yTRAr/Z35NMMUuaLZ/UIejL74/p3BgLY9bFsBW1MyC4Sce/TKOSU2Gv5n4Ob5oZu
hVCNLi0i8JQrAx2zVOAA1X5NmcNATGBqLk3cmW3dulmlQ2aUBuvsWWbIpkzyLFMk
tZInYS3FSIiK6RTOm46UGhIbpwUSfEA0f8wMvskT0t++PH8X9ZPXcyT742ChG7vN
PCi+TR14c1QZhi9+9y9y24aBD3yKAJmE4pfVfiSCS+egUjmKqvNgT/VHy4dF8qjn
DO1/QIAIYfglCbrXdgZaoieuaTXNdSj+QuQVu2A2G8y9YaEvFGpUCo76owJAPxRC
LUq9Bk9tmw5ZWq25PjMOaN89GpN7zWBBtheugvW9nZup7rjKi0kMfwQC+lnwcV1b
AF9RNXUxpR7RXRX5D8ea1YMEtS6pKSqNgd0vCq79s1gdRLjpQGqBR0sIkC3WOyfC
iuPMEhss1Zf34rEgU6DPrlvGjrIUMfobIOf2GeowPqz8KjR5sDLvoNfbC2eD56bF
lclDsdeePAJ9WYxht9TI7Zl/MGEatsnjkQWPN4bigxIn04zPdaqbJD5+nM4Ogqy/
/GgVswgneQ3HlT+6GZO/J+tqXT6QHhb7WSsX6Y3b4wZYckcuod56R2lnIsIJn8cO
E/VZcpEspb/sm8ZJ7FKwOZ0y2cTJXiOQGAkxMvmRVSP4IBMYaSt+YzJisjcLhLjo
tLeU8RK0okFIBFd52Mjyv2uWVYNGElLCW9hYPyPpZGuvEG6e1gnqcanOUEdC7iOc
oMU3hNCzIc7J+l69jZTUaf2WJxBEyjhKiPaHA5neEYQU6mS6OqZHJooBuFZSinTN
FCTGkFABk91VfzjaUadw8Gbu2davq+9QFLeBqJl6yYAtY28TTRJ2tprb3s+ecHBe
8JZRtOMSmrDgP6sOoZKgEcwo06ll8P8Ye8G1p4pTElCs60UNt2vJrs0GInxSCntc
vGaQToyE2eMg228EvIQqURwgN3fKxUjzaR7ztxV3UomT4qCqw+O+1uXhEPBnXUYl
Q3M85F9hBocrgLOsaedOd7niT/5zHLrnQeTAIdL+LmKVfnJTbXvCKjQ59q+7enLO
MCfM5xQB9v5hjQx7wdQOETbHurDHhcRW1CK3Z5vhqPU073PpIvf0nbbxz4HoIZGs
j47NFPgP5o8qY1pzqJ7c8x9k4EHIqxg4h1fJ2NHFhkiuECpWAN10wNtKtPuRVl/D
lje7ckWP+CO1YUY87Hf7jHj/0kAxhsXSijS3jgFhyD0ZR1Rx6Bv0a7ZOfvKp3rfH
HS4KV9HUwiE7DT8Q4nUmBNfRYvaNW9eUttvzBYsxpM40kV0WAFmuc9f4KPoWINfg
oDqx3IsALS8xsAnKZmNFhb++CWD0ZqpR5qAGMy5MGRSpXLFdEMpJkhvGQ8cFiwEt
qSaAZal/1Lp33h+LwBHwftUG/itHWJrkfH95waaGkmTsB4UjJDmrdrW3koaeTlnw
c/PWc5xFr1XUYEEp92XCB65+tcvhJaQAU3b87qVm00tb/Q8lMMIOhjytcQezbSNi
ikLO/9peZX7r2ELq8h/IwF+lcI78tQHVOuB+iT/jNKL0QCujjOEBk6apZgKKWDjr
ga+uDOW0h0INYVYLvOXoyOCtOUNmNF4NhSBaBA+ll/6im493tZ7Pg91zNJKrxmUD
I9GbQkIvqJZK2JtRXgI2HjxghChx+FNYX41Qcvet63ZpcPWKU4U6MGyMQ5BjUm4t
W8uDfzuoaePkAWWKwnJvY6TY1nuy347OVMIRHXYyWN45ZBqucpvxDYlRlK0WJYBd
1vgTWE9QHvNse7xP32IjcdKXINeZwAWzn4DavgTS6qsMjnS4Y4r6LG0C0H09qq3x
oy0HWxY1ksSpjgN1uGJKNLMyiWAuzm0EDIXPGI5eriYp30iQCX7WGotpNsnACgG0
22dAELLX+a7kl7wfHuyjBFWeqoC2LCQKclniJiNn9azTnXVsmqxRgsYgo0pWz3So
5kQ4d151h0hDTOJfSO4iwfT6xd2Nh8gEFxZjpw1h7y/72T/6PVjU6YxmBKfGfhHi
z5/eRUhvgkacZddyEE3irDykcnRCi3t6HOh1pqUzaBszYDeqYNIzeknI6tvLZdFP
xzyieqFhvdlIyXSlK6i+2AzQrhuIAl6vIGGTYNJZ03vBh9x9ppUtW7z9XioFq2+U
8fYgc+mQnxPDA9Jklkpg4eN87t3diK70+CWm2vzBzQT6Jw5kRKL4aa53iVaRgSDl
HwM0M4oEgWzv/uDHw2Tm4rc+emChn3XvvtWSrcU/4UPrdANG6DFwkFJe0ezQn6nw
DTlAVp65uN6IvnmdG9S/AHIr8trYQM3y71P7jL+FpbSMGt4GdQ8/XkEuPrFbRAMU
WkxYpMR8fBN1YQTQ7WTidLNBsZ1v8ouCAtKw4Tzlp7Efvb9EsY6z6lhzqxtSSzuB
GhYOIjEKUifv699PX7eLDcfILgLxrr5zl3HsX83mZIT5x+jTluNQKxSJE7ckNMyl
cr/gemN6wLMtsANWveqAVL0t04HduSZtxEssYkFZF65djj+5dy+SDawqhNj4+clQ
xkr8lsbFNNYxnvfMaHgFHdBuqxsI7iUbULMVw8KUhvh7mUYX1k852jZdupcEnRHC
HP5wz5h6JT4abPv5+DGV537cxiewGJsakeeo1VkEmct4XlBIMptP6TROMtf08vqn
QmVenSp+oeeGmuX28NyGbhFcw0f0IJ2FP0l5/CDuXvsCP1NzbhPmZhweYGkbyq7e
YfYHWEFPooh/icPbN9EqrKuxXoNCmZHp6ElWGLF6TDnkN3MmuppHE/K4h8PZUP4W
i4apYms5E+9H3EZaP4oGRWmkotkklVrK76cmNU44b5EPrMXCkvXaJY9e9jVa+kRD
hjHcG7PRBZFlN4Zz+QFnryKdnsI2IhGyzwTOHOO2DK9LxVgzqncxY0bSzVFhglVT
PJCC59XAIh1k+O3OWzd60sqDZVjV0Hlen6Iwk8ZrpXcT/PTyp1SRTD537IM7+mJH
YD9O9bvbc0qQgUnm8mbPCqqfpi27cHuNPblF//03bkGt0XPBcJMszx/ToaaOAJJc
wtXgYb/tj+23nuTx/4tr0cQ9P5QARKyrniBx8lCx7tQEz7kcF1j0RoUIu9HDEkNn
4ZRQLYbXU2v5LCavTJ4cEuGOQthmYqFMsAnzGkQVE9YFxGwB8b/NY8BTs2VxGxw8
yFyaOPI/i/3SJjL1v1D8OBMXUkEpZTPIXkqKtqYQBjn0OjWkp65ZTrCnpibqkxpK
9ipp/DrZdLNE9kkbC08Vm9a1e3PvdsrxF9W7oX0qpyFVka/sBv+fIV3AnFXPMuQS
5OE++oxQR9y99WQt37GRkuoUJSKj38Z/+sNZsG7Ho/H4REN1c/L5g2cMTfh+3m51
YuJOGiGHH9+p0cgkmaJOS/39OkeqnaSHu38kcvl+iiyeylQGf7KB2zAJTnU7hrlT
lBWIOld1ZyX+LB7e/dO0deOQBNqM/kjOmgPh5TmejWNXeZ2vfMyChi1SZ7xPXggC
H129CF0NG29J9+AsGSqL0M4Hf9IgiwrnCx9C2YI0PA1Fa9GNudhSuUZYv/sgFwE1
HEYjbALp7eL6Vpkl6jBVAt+ZrLbMg70kbVyzpCd57WqISO48nH4Mt0Ydohglri2T
CgXGHhQFZVfwhU4Otlk/zjqf2tWP/Hvfvj2kLsl+AE6o3dLK1xK+ofgCU+2HPmgi
jpTqpSK7rhsZTsMRV5Ya15Uzn+pxNS24hPMRsfNpencrLne51gezEcjJRv6eXqUJ
WFfHCmGv2otBeydoXca1jDGm6dxdpSKQebj+l4w713tnnwk0AO0X8ATxcVNUOUpm
juvumVfHkVbYi/NpDa7pajjO/XXS+96gjS69On5Bnz9G0XUZo5b2TOTVnzVCUcdN
pfYO/KvlxZal1Le/qM4erjiyX7NDV48MqmcXzbci0rPKv6i4cSQRNaxSswZnn0c1
L5HfbDfnKpaOPPjpYccOm3cNlME5mlEIVNgghdQobkvs5T1Zzsu7/AEANTF2NDyH
A7bWsUiNLxj5tUCa+DfeDnezcchLmdl0GcL9lYLwSnXtFphytoTY/75xnPA3eDTX
v3F26l+/tbF7C0k+CXbaZcaMVhlUigmYt5+GjcnTdsLK0WAGWTEbm9Cu2J/TujRL
lhsFp9Y5bFjUWYcRIu5JXRjUBp/emGty/Yrdl2g0bikHN75K0JbY4vqxzyLAcfs2
fZn8g6WesWYgqrmaK/CI4GOvWmcAzM7xiG/03LGM2tXX1Eb7N00m7OzERkcDqe/t
BOv31LywI/ig1HDIANnYCiKyfUnq3f/lLQNQWUYUJcv5CSC5ulp1TQ6EI2+KDFm5
mMVc32Ld1p5VLY0RZ8sN1+XigY+Nh+dQVMx1liBgYmMs1aCOhRekK2jFWA+Fz/pk
eEHOE79VSeUGNjK0wPHYKHKnwvtMIWhQhoRahvcKlgq109vQyH2fvRC6sT4C5/iT
6R6fZUAPp77KgFhv4oVg7QtiG0/TW6k1pwpeYyuZ3jnOmbp52iu/NBTavOhAUjqN
D6sHoLPo0ByssedRpldSe/CZC28CYVHnS7da5T0hjOFqn7ut11U9KV9s8oLotqcp
it9WCsYdjOIus97/nwOrXGPnsVgFoCYiBG8z9gFxcxXi5OaXK+giLib7yfExM2/Z
U54vVO8R3N5GmLfXDasS4WiEPfB5ohmJGbQdwpjZWre9nQUKKZNOH0crzz+NOnG4
asawYT44zkmGMb1H4J7c5IBoWarRz4eepRxlJg+ba0Fe1NLGkxIphlybr+dGUKuu
/q+oIbvjTI99qMAv8WuuZ8m/dYSs1YkLOMRKVQ3vKS7o/T4qQpZE7lwRi/2zURFV
skWEUo+wZozwzvRfLKAqR0uo8rtX94r0LfF9KLiI3SqgZ457f/mPSiaKxWxyFZN5
kej358F+jnAVaHgNhACMXKb92If+RD6ULf7g/9wzW0CLH+sU2YDHA08dHG+xF750
OWFlFmwriS0OeKjkEGLc2q3AhjP4AHF3X/NwlHYIl1IfFpgv/yPnFMxNQU34PT3A
hGYXokPF+YTGZy0zfZPEq8VFOaoRtkdcR+i1vk7zvZzAZ2FoLo8eTmdV2fWxWTBV
i6IGKSXj68YX2eS6P/m52VBifw0xhD81oPaRR3URev41RmoNeKMDJnDIdDyZetK1
gEWqixsFbdfUbE+bsTHtPzzESOPRpneXyHEoJ1BLc0lsncepVzv94NP3YOxIv/Jf
d6aVi6MAOG31ZRtfyvC8Up/BhkVdH7DibyrDFUA4LHibLg/AZReum383dPJd2o9R
A7FBFShKSFsV8dAlNhQ/s+bl4tXaqPxHpodkMlmX26291c0YQgLWgOPLVV5kcPJA
SQ6fkfXkKSg9+q5mLcRZn0+eyBCeq2BRPp2RNrmvU1dih+FydTxTfLnRbkCscWIq
v4J5au4YIDOl8cm6JEkOEilej37iyZAo0oVe2pSrSXYneaxe4eoMBy3xGiSyXqkL
rrtHLbYEtSlI1Un9ROrD8WwbayhMA5mFqw5FNYyNOMQ2Ik3gRK2R4ykjNadj5+CP
gkhL4qkfqnLxb/pI4gGhUEwScE7jsEi5JsEySYDCHXcWlcRtQM66stxT92AKTfrZ
9F244skDTGwU1DGGzNRjK88tqkwZVqn/FyAZxz1C7gAaSczivbNXevM8PADNsfDy
orJYkGPDK4RWalaG+ytu1lgvrq/gBnVT4ke88o5cF66ZPRJPAV9zzwUbGO6NZWLT
hOBmkA08wJt/KhGTLPfQzCHGPu/E92Am7VMxqchPsNP17hVz2GLMfNYJdsxyu7gO
ZLVYEiX0B0Zd228I1fjrmOi/QUjLVOF7cJMDnb7NBN8OYABPHBkyZlTqlhDxFrLk
RFdKk5WLaNBN62bw9pTL7gbg1KBrudkUMHuA1/ZCg1rU09GZYPffRV8d5GVR5p34
Td1GFrkAzfA53IdmOkSC/eNblbTMDy1JeV0sZ5bGFxeY+2953qRJD7RuSrh34XSn
oZFRuoNswSHDfSgNj9SAi1V7PRgR4qk8edzHKct/35ERdW6cE9D9CbzCxJZtg4Bk
FMHH9lA7Lhh2uqLAirp/D33gl7z2sHUZn7hi00gv7AdrzGJ9DJlN3vVgFSTeIqQr
uVDILNtBz6CvShJBerx/fa6IER+Vp4sED/uOrJKvkwdjb3Dmv7JWuwKS11THW4JT
fkxLjoP78YN0/gYozpnX1qeeCB1g09AxwImREnS4IA4ugghAfmr4R/Ish/oYYsUG
8eKfsdjCUfGWzF0HKNlhVYGj7mBt5+wfT6Va3jj79v1S63qcLnIp3yAKW5lHiqpX
6B2clmRlVeByXz5eX2hleYeWfCq04bLxBycpE9EXMB/GeaRwumNYt5m5zN8d8BMR
uHefmvKdx7+kz4EhMVmTaUYk7v+2WNhlYE2SzdP0vPcGuMRB5AHJcK5Nu21dsDP2
M2C6pyDhaPtod/yJbC1fwAKiD7aLCckDvlliKIjf/YaxvG3j7K8eaFbw5vp6yKOI
fo588Z4pLMDEf8OK7aPujDdTugwrNv/XE2cgq3tGp0XKsyjFHgssL2XjJ4Vr/1LP
NIgpjt4/s9uNQLGFAZHhd7PykmlBb7LfKo6njWmWqV9XIkAU36hJBuGcMHk+cuv5
kzd/ciQiGfwMncX86q8/1mGd0qub9v7tf84rNbHLd8WT9/xDwxlTdHRP/cxl5rCn
3MJ8MGMBHnx/VyeO1JNB4np00nTGn8h2sf2JumWEk+ZfIAHgX63vvvAKCpiok+8S
PjzoBKO7uVUPRx9sH0S64dAk22QFFT8ErEAnn4pQEd9RFgSwquVgfXinm3y6vzc8
iLMQQZ1tR7AX0Jj5Ajgf03SpwBvoLp789ijJfwWyNEtAerK0yiUPlFDwVSuvpQyk
5/ZZr1RfHz9TxPyOy72Lkvap4IEhDKwGMpr9NO5xXcneIagcnDs18m0YWUg99Ssm
yajm/JbWvbxYJdErSrTuF8YkAVInTqU2BKpZr59dWoASHCpoDa4OUm5aKnwUKsHO
KXa2kdZCnS02iNKhK8Paj1gT9xp4VX6mtAHZwHINSEqSoi93DL9kdCL5QqUCjnCy
2hY3ZrqQjt6Ntq6TnNSqDAsG0XstDr3yTyLwssKa53lThXd1OypmXxdL/LNhWUaY
PFfo2bZgKKOGo086FQTnhTBQEeQhV6uSp5jf0jvbEyjMZIhjLWD1xj/XUjKEj8D9
EohDxF0sViHThFbVFkwZQLTdo1AS59/Z9YHhvbv51O1g9aGE3czaSnFMZf0K9bn2
/edq0xZ3fP4aS2okJ7ASJIByX26vTjZPqy/yEEFyrBkXGH+9l9z0DMFlB5Ro05iv
AutvNWRPUMIckGS1oKwLvO9pArfIFGlEZhuapw8wTzNoN5IUtQMenawR3cVD/T3/
y8oCz5Z3I7kWzYZUmWOcEMry0+eJiVfkTXDrru19GLZ1/yjP7HI6I6t+CvEbmdTu
L5BJxE+5QC6FCAlXSgYHU4tL3POLhfTNPFxoAM+qhruvDJ4J1kytjjqxFUfX1Bwz
HFfvuCo7YJEmK5QmaaF0nxa69FLpJLYIUUVcut4JEeBPAmK2w+mb/6s+hTu1Jdxp
+iVYagPzZIRE1Vbssc9nafWU80CWFPrrlF9fMAbIwPuHBfM+XsPXNBZDeReqVZXW
pbVQpKf+3Ng55SkijcYR9pLnvNnM/zLL1RnMGcEK4CObp/0hFNTKuJ6fB5Va1U0z
uQaVYKiwp2yvX6H7bykrezp++2QkxHyKbPyUIMSp8UnQnizI8Beo1mRZdbPsI1c8
cKL5b0oW+dRzfsYLgHDRXdj6xkJHQG1lWzFUOu5dM4sfiUPFEQRB6kAfqDTxP+0C
cIkYt/oN4Y57LKBDzKxiR9GadpU8NhZaPpznYXesky8zjB3NMYitfttH1Jn7lmWB
ybFOYnRiThIf+Y4ceNsf6RLOdDRolx7mBpRi4nB4xqvXOccKWTRP0fBSei6IyBka
KXXcpXzoRxvpa4/mRHbgOhQTdrLiOrFJYwQr/c5uRpCM1323YkZRecJGa38cNFfc
Ii9elheW4BoD5mO3GkvdCFPN08fWF2+MpgKw6+Li2xx7olgEGhSgUQM7zzzG1jST
O687DmrT5IYK1vRiZRr4BYRS3htFf7x/4Cn1uHL7+jWaeHB7hCOMnEVBy2VhJKrm
aJcbUZ6Mc9nCs+GGwiMcLRN+3ChP/SkxFAtz2y6+MlD8Ln8zdzE3vaKJK6fivw8O
kCd5p61RZhTjqlpht/q7Mwuu4OTO7TVmqhECk2PoTrLiwe8Fh4KN4Xul072AJTr/
+EerSDtLbyzNpGDLmC1Jwmkg+IC4hCRcOFwDYxQdiicJNA9zrckKaZ3UfPfFg+o/
UiFZuL4gGnZ30Y34h/4n0vsSagX2xpQP619kLnDgEsIwK37ZFxjKTPdB/5mrtNdB
ShMooCij1tFOZrmM2F4zjwZmCWM6Z/DdpPLfoq4rVqPJCuOE1a0reqY+RdituL5Q
KA2LP1CllpiZIwKz3eNWlHUbnjr3rtQx0Q0p15KynMsQxFe0AdCW8/TRgvSUyGDJ
OMfNZttljng9C+aphjU2c1W5tZSWjY7QzepAqgK45UoZpCX1K003aaokQl2pOiQs
eIp3ylhzuvBO8NODIyIQaZmWUeK2ZMNrjyhc/MEnxQwd2uGMdIF5haEwKrvyNWEC
Pk53HnwdeXSHMTErVDtYhr4M2gmdHTkHYsjXXde7dxa+ICHoIPCtSrnqWSjOrTU3
qT+T0AN48segNNU3OtZBe9JsZgw1hT40aMKWvgvC/0XxewkwGANocLrcxMBFk4NI
rQoYkvSzyob+s4VQ+5p7P43LX833vFlLK2R2MU0M/CP9MYX5M6T/Bpj4a5Nrrq8c
xbQ4ymYcz/Pmij9EJ4pEmjcLOll49kzQLfOeQ7458u+4fvXy0WwalzgeH3UNUgZx
DRrrC/ar+3SGurv21tB6jGmcJgcG8K6A5g/kndSvZce2rVxdkP+3UytrI2+vEbqU
Svk3E8efJV2jckayiCm4fZK+cqd+wWKVCKM4LTvtSFMTGDKWOHEB097FMO1DJkIM
KwVri9N6uJA7UNZvMHlyz6+ykZyl8/MFo0Xac4MKyHpKcMtmji3ePbHUDl03Ft08
zahbY6JXyeUxm70wGlGm0cdICoqnn47UlCNppVQRIyvMeyS3Gs53c4CzD6hrzjET
UDm26lI2UW4JhywJUY3bZOMKVuX928CxHd4Q7en1z76XBEQ2k27UTc8Eap//IYmO
++g487nL7smOla7R2rETNUCMz+xqQ4SmKhNJTm+A+OjZCmWfkTQtj3/w4vPUONil
I/5BRFxq4SgLaItR+3bC65Op9loNK3ct12LMBEfZqzk+klRm2T48ytMiLMBdjROk
+s5qWNOrqkglSZr/wFRbt8q96+w2q3psbOk6sFFKj5xgKHA68xf9ZaSkAuib4Dvq
KPL7YcSSB7FpyYL4Q5QYgkZpiERwycV2PuKbUu0mjeRmp1NNNdXElD1fmGtocq+A
XC+bWcmZ0vHy6uhBQNsrv4ispF0fzqUTCdzWGUhgcEDFO6gxOI+j33nVt2BBdR8j
dIXpfx9GSgBMffDo+1Z+vQ3Wn0l8chG7y1R3NahmcFsuRE2w5fFxpDeLMVEBp4ZR
TV3k0dzjc8Q78nB4NywXfso9Z4hBkVResFD78F6ab6Mv29DAjuHCBDMob7lVQeEk
1oOnXsFm8OwSeUgNGn37T5bw2UdG2EQJrbD993wyDzM9xiXv0+lBYlBKo/1WsnnF
IAClbkO6GSnC4Sx72g0ibo1ozScWvfJQ7WIyeAH6Kc/iY8zA9cNzjDLPHAxYViTZ
wuUkMUq69yid/ho7ztqhxcsPgB1x5j+Duu3IqtJMp8D+B4RurG6ygYTnEYYCKfM5
11PIrGW1C9/KB2aTZ7z2LEo0ERQ8Br8NPP2FdvV+KTGDtk8ynPxHP+VtUZ1ahyJg
OqLqZQA+j50EqquMZITBfLjvn54nxzsKDmsXJ98APBJC4dXrS1NRvFb3lxpDa3iT
08wLVUKmrieH5xRvHtao7QU+xiFjHxGGl4cRqghIelazpK0MuScrZu/4h04oDKbL
ZhkMyXjusdZTduEfs8AMRcEhxpZzKGU1AHkwRXp4ZVevCueKSNnPLxxeAPUoQoFY
TLLtWiudVS2RQfm0K80INs+jQQJPVI73/qMPwohE1Kn/6eaOAI2cqx8cThNDBRbk
XLzcts/1H49uQW7dKxmV5CzAxGTplUrGV1tJ4oDVhNMWdxhl/ne8RLX3Yv6rW8N2
EGk9+r/qHu9KOBQ9Zh6lYozCnj2tyuc+Z9Lbf5dX+yPV0jRhMFHX5c/ZPtFWTscP
pkRnKYGIZCKx0Wq210bmCyabgEMqZF/SybT4AHSVg1xzP8u2sgkI694u3dOxVeU0
VLuWUV7NfeB9+TpFg9wt/xECk7QvP2hsNaFcfy8ehu4GXkNXm7g7L9jv4HVQTVxq
t1auLdtr8exuE0/N3315rp47JDO4iKustPeq/6MgB8Fbrzd9PKJmTFycHb3OmTA7
jWynEacMf/x1fcyY9TREroqg+/Y3x2ni2Oxdsg0VX3lpFKh5Fsie3ItkrCatBvyl
xvkbER8P+9xvsSNNpx2i8I5aNVhswDJ5gMAOAfVWTcmnDAUWA8DlJ+f6kxBgdBbE
XQ2kJ40TQGJIsCC43wyx6ZWzxPgTGmF+cKJIRCIEAOzlgO3U7Hc4rgSOYVudvbmz
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Hh/fg3FA6CaAIoltz/9rLsSu6IR9GWvuVaz26Z6axQ0k6VsOARyLwIP7yBa86W7z
7AXRWtK9QtFe0yseSoIyn/VO7QWwQZZB2kFaVataVvGzQ/FCBbSnKqCGtofnE3Yu
mufsTf3wsbe3xsBnK9WPpYM/2KCMUwZJon1yGhPXscYWfJfBJXhuUUkMEp2TRHsC
T6cHWvz3puhdHtuCgMpcwkwj8oNZKohjKMATpAFPpzxmMpNIKZJvCjaSOU1TcyUw
8LTBOK40whXLC1PI7UjZSMHSAWSMJBCIZrYmcnLxSqi57lA6PGCvYKm231gUTcOc
TsSFPAzTNIoVaIcMCun3Xg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 21648 )
`pragma protect data_block
rZflI5lcYG4D7DsPxEedVZ6mXwHhnn/ukGSGlL+ZtLn/5qH+FKMbXKIk3S+IH7Rd
sho+DKkaue2RLHqNvyIhiwT/otZ//kR6cDWgOKcLojOFruUT6MvZGHqjjS2oUTha
Xoe2/y6uVJyWewkZNu1H8ZtL1DalSmHSsigy0NGTCMglujAFVMso6L7I73XTonWG
b5xaBdMgjJatX9idmY6O9ukxGHONObqHuvkbx57g6S8YGTt/W2tiCi46Y0Q/nI4F
PbJxEOQhdweBhoCxALmjvbxmzIkiMkclIiqqxQsBnhw9YahXdPX32NFNA1h/QGcu
nGCbcn8vND3mvv3YfcaVTHQjgRDo+ImYd7Pe0ARHKHqHLjnpQgy/Z0FX3iXXluht
uXmajkcxNA0omD7we2NNQpim7z3vmBaa61+TxFwOvLSspU/qNG/MJ/jiy5EIMAIP
UMJ+jXEd36ruJKZ7H3BT7istjlM2KPeKbld4xPeqDX55yFKBmJ+NJW+RysNAw8LA
6k0OoszWF2veKiv+zDkvoZYRl0T6mhugT1BoefaXK25EsKM6edQ2bKhAxJFpvu1o
Rrz/zZvlJQ7LQiUMTG6234Pw0Dt9eA0x5JU8TJDZFcKUCJauSxXDu7IABr6NrNA4
e1VZjM2IgMljBRgioIArwStCyDu+Zzz2E8rClCOjR3tTbmVooBHiG4+MO90r3EIl
yVjAXb+0e5OCRUIOZcXOX5K6hsgghaNjp8/NgqwDJHW5XHT6SpGKB/OQZdqkj6Vd
07jiVZ+E5aTb2e8/aCkt83Ga1Mh9I3fNj7FcIUQa6HpWc5n3/1Sp+woNS0hekcqj
F6F/hcE3gCXawF8+sH3Qouz7aqPxqVT8hA/51plAEeBbz5XcQlEyB9Nu6xPHdSbh
n34wJGLEmOfIdm+oomCgl9jT137TZDyuevtSuSaCep0Ghw1QPSGO5t/HBVYZOAn3
RgCBugoG/+WEC4MdNli3NexoxE28L9fMxxb9HBqXbTxO+UmGBjqq1fMQLHXKSCyn
73TBgH+Je+QtYLVliCJ55jeV0TRiHsj94JuCb3P+joHC+Qm7mcPemftesk/21JRT
Qu8pKeDBBkadXwko4RNd6hIwzKIoiHCB1hZ68J94Qyl6GUMk9XhHyZ4Ezpb9UVum
jmRTeCueBanaektNDsiIJIbbW/SFKFvmb0aGdoZMDLIxYdsuBAKiZtWsQ8eUoz3Z
MuQNIBL7CFOHkK2jbSb0J8wZ1KU7TPTIVwkZX1mWnyEmGukY6ZlyvWXr68SIf8mN
6GkVLlF0KRONyOlyUZsyH31PVv7jS3aI0LpMuhh5RQnR9iPs/wEICyTcl/kcAQuN
0aAPbefbzvSRW7HgoSDibY0hgvXxkCJhrHqsy4e0b3GVwBrlnOEiwQaCwHk98CKA
ONsFeqNfig4UeshGxh67h5SUjD3CvA3w6NT2EY98M4+LZID9gWUwqwrppgJAZBa0
9bdrVGMCUDeL8WZn3rA5n4CUIWcc3ntBQGf0OrZcOoJ4jZT2GYrHlLTr8CcWp1pL
e05lqanhPku2q5VcKZnbBlm8SZvaKLhgCYhv+gPSQYr4WOClb6CH3zzM9WlV3ve1
hGSLIoZtWsOw/dzn1r6pPR5aki9ikUU/GglYFIBOx7bkCqiTbLlhXfPyFa10mgLW
YCykDL+FktaGyuiwKizy4I3OnivplSl/nIq2fAz+gxd5rFaERzdjPCkMYd5A7+/1
UaBEHlaCTEdyr9TSRXYRIoJt2G6spsJmjqzUjIf0Fm5gW0B81WSOOtD8Y6Tliycq
iWVJv337ZNReRgbPJy/nhWLN3X4PHECbG+PGmrx2vKVV65WR1HVOiJg5qoGHdio+
e1Kyuik9FThnFyrO8LHc51cYefi+XaLJXTV94XHOyJvvjygop4Xqme1VyFF7nPFz
TGo2lSumSn+IJhTh+s5Mjx6qtK0wGgo94J6eHViRjUni8NwX/V4ZlFoIE2/dh4GY
rHBGbM++2vOz1X8OnPqscxtpfxW0fim7MbC2wVZ5RNKx9iD+qwyE+HY7rRZg2sNl
twe+FouMQoT2LGw64yWJIFYUTZnTJl7laRuM+V9kaA/l6CUtKGlTqserh89tjxLl
QOhkLtxE+4hJGS7GQu0i5tSm1UvJl2dETNU4q1Z01e1YqJEZdLcqJIerMYi0liV9
NrPxoAH4jKEu8As+FaMkNzYarvrn4qe3FTWehAnFMtgUwAYdtZeJ0MKKZhF9CpyY
VcBtWyt7Vg57IXrR8Nn1hf26auulmlkvs0U2hhB9OW3nrRgw+CO5aWHFVOqzQEFE
3RmQCmXIJHLafp6iEy7rDjQhDDU5ugkd68B/M2VXIQSyuRQvHJb3FTvfTgcFUYqX
kn2uyOxSLOQVtzfgk8AzCnop93sRFmacwiUfcVxeGSbEyKwp9mUapshWxtjEzf7d
57WAO3+bkOgX7fbLo9SLT/xSQFMHpUYrkxZREmNa65NQDaCcAB58alfMhAwryUSW
BrE8YL0raqnA3mSqyFMZipJcJ73Q1qkt5+uOSH9yoHmNJCKEMZB3pdR3XHHwGpVz
aucHRB7ANDwFG3bYpO2WN++DTYeyt4JgIUIE9hvfWlUBA5Nuh1jPiaeiieJIv4O4
2upbHiwwf/SMNfNRQ6/H01ZsX4SdPesZxgaIo+M9sR2mWWWe7AEj5DwHY9g5BGev
fyN9J1oiE5K/uybfzDC0fx2pK8c/lelBQ0qeFbGhRzboYgPrsLOjs1sbm5KwHwFx
+Zg7QrcFbCHpR1EgZEZ0dtmk0vzS+E5W+QJyUtOYMHSKwOvI6121DnqhksUbf3qN
EY7ph4M+wLkHqu7Rm+8wLBLII8DbMghjKWRdVDAB1hkJVYhjN53hG9sNLckCfion
410UKWdE82v+uqj7+OjjMKxCwzcTChqugR47UtV2V/+IlfBB5BpMk27k2o+kI4gg
w464k0wb2tAhs/E44prTBB/tg9JgRY7xfgcVsSzKe6UGcnoFglKmL/4YMdnyxlxU
41Ra2uCeXZMze65RzZVR5xf84w8m0dCMDUraI4QQx+Tg0XWF9Amw0T/DRDTUHnjA
zfizVHLqAGWmoUarvYLdXcaCLMqinYvgNviPYKgxZQfj8qVX6q/FPysN61Dm2xWS
XAcGDYa/kWDho1cHbeOMxWKSu2oYQJxU1gN5+iM8VPGq93okv1yeojWGu22Jz0XM
T+n4vKhg20DFmn+fZu7utWA+KA8IYCsKL5+HYLz+oeVJwwxhBrwu5Ph02IfQCNCr
q9ND5ieiJRqJgrj0JbB1gXVJELHb9aYuq0qUPy7snZFi1BHPrCApnT1LKqHkGiK0
tIgdFvIYitUSY3TIraZSwg3MWW4TNLVx1UK2sJXwukSeFCS/lNU36JNc/FOJWH0O
ZToXeoFht9PVEUtKtgu0EDjmKTGIsJI+zem2irW9SOff7Vsb81u9RZyGyAzP5FzK
w2Ex+jsrkIFRx2AhJcvWc+0G1EAY/jC33XHjjfueTbuR4c5Tfgn8cdLV9K5ILU2a
KcCBenGXMV1Vk/OYUrh1tzlZ33sQWw5Q6H61boIASivKtb66jDSVgYRO7m2I90H7
fc4Rc6vSPvC8mkUpcT76k9noTocmBUXsYahZjn0t/ycorvWlsgUwzwLyhx31fp1U
j3yFSQupzv2m93qjIn7N1lGtgKxoEU1NTAOHxxVkcpWyPX9hMtzXyipLMF2tZ2wa
2ChnPLcDtzBCeGKwE+e57x9gHODQBxaRsarlCmAo5Pkaw/cA60L+sRgflht1NL0D
AaoHxAfGjtHOjlkJ/nrK6s8LmK9pzdseXXzKOIfyPr8nTxpK5fvdCt/VAKZvsWXO
q54yA9xTxGMxKgYXxKsTV1VK57uPs3Jd7FvKwycLb+A/4C55aFRthVdYGLhmeWi/
mPpA9WNh6W8ISlJ9v/NoDFWHmGirUOT1APCzEgKx3MwUS+Zwk5EZOF0dZat3JPoL
T5B94W6ABApHrBe5YKTGG515Xy3M9yn9KRnbdkWtO583nLtoldTMrNgRIoKXqmUF
dvTs2G1SuUXZXhr8Db539c4wo+b0fwQ92Ndh8k2l/6B/hUhr9jAbWfQHVmtOghkc
eojkFTYQTym0Zze/WoI72p5GlIJZOjO8FzV10JQrTI3cLfhGGMHFAuSzk6sANmDE
s0XoBf9b9B5TlnKUPF44PDIArqrhg+PWuHHiT9FMGxm4Zzks/SIbnoxNoC2uE9PZ
9woE95TBENs1s2WPIwSF2IlmcXgESSm6R/3YJjA4tdXqWqkQSw86hO5Fog+JV/T8
R8iM63MUeZaoeoplJG9JGU6yUlyPgakHHBxfxhRtMQUdlW/B4CEPWLKIHS1sFwOW
+rPXzick/1LBuS0VQPsZd148twCnjfnJKPgdZ2IX/o1I7NWF3uBRqTopF6WFiGoZ
3BgViR2EikWYOJhIuMtwtS7uZb351mKDsET7X2IuuW/n1HADBi1hqPDQ0RWeVDFz
fh5Bks9YiuzomqGG/8AMKwtg/lAvmQpQg/Wnkq3tm52Mtm+U4X7xKmF2oS3nhPjV
5GzEPjxpAODlh/N7c0kf1gQQk5HpwFpv9R1xjDa1FqcWdKdUaunq5/b0M+062pnI
S0RUkSIHfUbybbQJoF9iF9dXhf6UVxbsVKtPjq0NZeCk5qpYNwaa+NAKUyhx+SVQ
SCM2Hugp7LWfOOm+gGjnacCvhE/qi/juEniOFwsEplkEPKUxHiQV4WFSTlXoxd+v
XVx1uubbvvIUEyhQDhE96Ozv0k8stWR2hEywx6Wb3acQs4oUudsz/dYtfuSZ6r0p
6ptW9BwytpzrbI4bzi3qnqbFbXnlzLxVKWcDaZt7jjV94Im7vp5uNQ9qo2+vUx2S
YkuylBf4MInLjXOCvOcdiN1rdUeYz1LvfoTRi/sX+QAFjpMoRbw7kXMKhU1OJasl
3gtPRzpAEcv963jHPyBmYgEvPDDVbO/48XjgFipgf4YadWKsfLlnaZHag0iVQAIR
wjRL3756N4SooIsxEHZ4jWDTKgeSPa6jVDnYf6/0G61+LZVhGBKg6dMO9BcvujsD
I6R0pKu+ek0OEf4JBc9nGxlg9JKsENBtDQNGRRBU1v60iG40lkJil6jSemVjbYIv
JfO7HEL7IlW7UeGGK/3MclSlFyhyzRzKKPnOIT7Pnei+iEeM4CnGYVSSO3QXuU7S
UGXHP1rMVcSA42NNo6vhV/lc67m9Pho5Zx8R2bm2c0zgkNnDrhG9rShA1/VlTIjj
wV2VmC710OYxCnVZgVZRQOAciKevIRzBFOKQIsZa9wL47FrsDNFAclZbRxSXQns0
pc6A62g8xfdhUbdmzpH2pX6C7B10Q4BExzxBDfxq/nYM7ySj/t7BEwQ8cg7Lpu2S
+HkHfgB5BcUPOBAeNVQyRjJuCbM5b4D9hhjWx8bi4cOfrUGBtDz8iC1MlLa9FjlP
NAH74MgaOr0qsJ10QQNXtAQcUlCmw/LqJv06O2yu64UaKwrWOR1BUUhJamzGcCHy
RhvRj9ghuyE01jxmaXr5HKA2s6Yaur7tyfNwEduOsWBJE+N2YkJDpSbvoG8UJiLh
zBKBS3tQMl8k36i8LeUONv9/x1JxqDCuPr9/iizzf+Q1WwA/FgXGjMDLAqapds/x
ah5K5KmBBSZgObwJRtdFfA0DXWNlFFI1h3j6xdVabudoqOnz9XmRCwDNqAsMHPsn
P9BBrEOPmJHIwm/JjtFtuaRKc/Y+TYqr8pAR1dz8Dc6Wg7SgzgWdfaG2L5B0/ALo
W1MKXU8lOFK4yKLAlws3PzAZnT+WY+1xthkqNohk2ObFMLOK7z5KAzGb42RN5KqB
qoeuR2RclW9c27Sngn66FKSuyzSTS0+56C91kxziHTQNYwPOcuxTg+4Ll9RDI9zr
vPJioHA7mctQ3+wg2QSLhSHI63+xF8FmkquibgFtzsJG0ZuKZiR6nRtJ7crjrPDu
qujQJpXAxJtHO9WcUdevYhx5Z8Ge8Ad/BqnYZAoJvaznGTc4X/PDKtEhHKqbJw4V
NxKS23BW1P+UomgEH+GrOkdKxSV4GkUsXaypqPfMfhhTtvnNs50rD2S9it4n++tM
ftrG0AC/rAceGxgyqZvGCVQCRxIwJhrRC7qVAq/+t4JBVyvVBtOFgUIrb8JKSine
yFfmzu17V/hSg6WJITO80TTTGxk7J29zyikU5myOp/WKvsDjb7gU2ufW2mkSi+VH
1pQeZ7MbdGPYhJSJYMkt+0Ws2MvcZl6m1mqKIzU2jhMnc6nYIBBrezsE2ko98693
Xb/x5P97WU/C2Yi6TUvsY+tHeTCQawALVacgcli7/6TuNiUB32lMzdzvLaTHYAS5
tXPfa8sGPRrwb41IsOjNEpuhqg+d8jTlGb0DUCDVktYB9//qzm2CdA34g2c6JJ7G
25MbxRgry7zylgc5/raaQXwQyTrEVnpFpwwAHxsDGkgy+7DsPq5SNB389nBI1WLl
lsRFs0bdmnXLwet4DyiyFHTWtpkmLvVMyCqDqm40aE9rZuRX5o3TeExJ9DL6sjeN
71eqdJRo/BKwcOVPYzg0aqETxq08v323cSOaFgYSiWbkiq9ACySJ+zoTfScXBcsm
nlW5P23+qE+h9UTQ/jPb8/yFIIdekFWrFSMb3emKgFMyppFMzDbj6dGwAMUkbjBv
aZ62dhGgM4+UFTNZN+h3JSX+m0Oa2gbPSJmAJukzkVXhZ35Xy1IShLkA+0BvcAvH
wYoOemCfQjaK632DllWVkJk4MpuwDQUMvyzQeBk+5xYJEfg/TJ4wXTcaoRIxguZI
BY9qqeQyFKVx4o7JsZWYUJSDnpj+7gBQORgAW31mGKFk9VRjEHEE3Hm2uguzWW/v
FCcldBq/FdmfoQGcWXYag4F127w1mphgqW4riR9je/udiVycfeKZTfrK2X5AUARn
Le1Pq+15ca8Xz/D8ZYuGe0QpcD7qsP5j6b/zaJMrm7B/1JlhgN5ctJi5L81xB/SN
Ou2I/zdGBmKgh+eqTRPqV6qeGPwoxO62XZxJa4X6/W0fjvyIqq7Nsttp7BJpQA4Q
LGpsi8bOFf8ViquQWGe2hW9w7bjkvkO8zQyCvJ74bvZsMuaMSFVvVCkVZv1Kb/4s
xTHtTGAAd1DPSIaposJ5Lj59XTgG0iTU5hOcX+NtI7I/y/VzDtA0ygh+EK/Hq70I
g2nC805NMWMnCRMZXTWhdc4Yli9K2endQc9aoBvS4K/elfPdzvXKHgS/IgOriuvw
3uS/88vRcKmYv2NMXRgmhPJRMLGY1wq+jcYtq8Iv+GiXO+FUX10boROiQbIARKYS
5jhvGAU0vK1yxochlBQdaD0/+uwZkJ+/+3bcmx3Hlz3sqNPMijFFhhQqBA2NzYIW
3QXTiv4PwGc8OIl5YeS7OC0ALlMrCZXp/Z8CT5E/0hSVR4Jsa5PyA/S7EJBtC6wF
OfZbMMXgx8fL00AZKVBgaOSdBEFr5NdX30KxAKvmWHe5J1ieXU82VjLv/GF0TURY
j3RdF+71VMJIi/h3IT0tyqEuSHHkwmX5ofDNtcWilAZDJV+pJy/h7xRfG2pFk066
ph8QxqrMlAs/x6QmpS7AfEDRs6E+oosB7ZmFOQ9V5mCSy7g98Ijnl53CLNqdJmie
YrQQr860Sl9AMYnxKDs9GaOsSgZ/bU0YEdWWG77wPeTa3109Y89NAtUoNYhWmjkY
WsOIaSKuObrqyC8fDSIQxEuG8yVU3VMMp+/pOQos+zhJGF1XMsu3QL3l+0hqaJAq
4EhyNT4Ax6Db9b62n3ylh4fXmVHytcZMeI+mCz+zAUKQIW+HkxtNS4wrJ6VQIUUw
huD8BCnICHHIyU4fpg/M0tI1r1kmby2uSsf4sRhU69t6nonUOydP1qk6goMMe70S
hfSeou3JgjQfG4yMzFTbZ7hgbjcNFQC/LJDWm0O9Nq5DJ1YNs+FS32AlRUK8GoBv
/c4Fn4/ThPhPd/wDe9u4XgiLqEuxGVfjXJXF9QvpBLpP11W3I2A1ueUEkY5z+yYw
jh4Wn4XM7LtpV0qkZyr1E0+9KDy5Bi26WEqQlgsHOV2SdhaqEvI6jkQutLLbLNl7
GgqGiuR2oqm3F1nMVmkxVz1dkYQtWA4zlIPWBrFHFJHKi3XitHwziJUCPy+J9LPO
dd5SxOg9/p0HpDoEHA02bGUiZlFyyNvvClca7pe38YBlWs3ZOPkMmHksoDpIo3HZ
RfQ2luSouqm1V0gubysl5DFRRx1GHQX6TwVBV34am8MUF04APQkLQS+8JBDtZ0NZ
ERCuxO9PRmGTqZWmYDdkqVa8WDWk2Cjp2Enu7ao2fEnlLQqOEbe/CKvr9a8Za/iU
GzyiqNyk5QXcxrJakyxzARDO4cRQ/okjUHKiAKuk3gZPrgPTqRApooJGa+KTzNnV
qWFDW2+v7mOAvgXV+/rumzq0FHivQD98023PIQRRuLBYdPieQQfJK5C7jWSYpT7i
NKOkx63uaazAGIH8+cMBHDxQcMRufexnHYz3ia8BQj+OLu1YcujHO4qCRIupsheP
zQbrIICrghP2nPa6XJ6XzfEqXNvJxPQMFemZHpbEQ/STlA4Up5/z6GVTaLaRn72w
IWxAnQuu3kJkmbBmCjg6I1UeTcA0+49EHzGeCyRo3aRNZTB2k3ISbP7d6uyiH+vE
W0iuttuP5CIbb9A++OTNLX3KK0mEHDNe7DDAr1H6rX/y+CFXGtpm5TCLc22pXvA6
pds/ooicNgaL9UYCx8+crEuMB5x9Q1esQ6Gqkbgg+XN6ZcoHEjOt31BT1GLVIrlT
GXfO4RS39mK8h+ubQ4+YKA/6y3TMZ3s9TEgnADUeGq0+nt9ONchaZku3yJb9MbpH
W6D0Z5uF0ypYDMcArMIa6vl083R8lzHuVGd8i163PTaWRc8kAIqXQQB7TyCaBBd2
XvzvsKCqzRfmU61qrs2CRi86oGcRBGRZKdrawAY2Fp0GFbEi/HvpFQvS9OVOz3+o
08UW5MU1VGY+hxZhad4x1tyHpkYOfBZGnpsjJbzEekQxqEQ4M5tRBfjRatekWI5m
tjMX1ph07CsziSSCKOHmjngZAC7jdAZbOLTiU1T17xzS8YM0VRiGz4NONXtOCUrX
Do4cggkJEL4pqwBP2Z34Ph92NyzB4p+jFAmPW124qvWyj78N0LHwB6rf988Pr11w
wiARMahle9Z/POyNiM7sEgZqTXQzza6ZutJ4+UJw0xSx3nbKPbhGBNEInbs4o4UJ
DiV8fTSPSXPnuh5w/mcbNfjzvY3Bh+6I3KYFaE+UYgLF3YuQcjLF9vlzFlGz6CJb
3zWw3sX4Nd+qkCcJz76H5QoM8k0+X2o+XeLWWT/QgaKLzhCP4ZQY8rRp5UHi7gam
PNITfoQgxG6xWC5FLiMz8P14PWug8N1K4DUK8ikOeUDY0sx7uX7uLz9oUH62Qq+f
kb6mEP04QrF/3u3I+g47gcXyXChP8VPbMtc1UZS/j6XiMFnpw6NbJlfSB356Fvyu
Z4luyaTK+xI9UIlL/LWF2EnqB+WE6ximPf2OZD9Ke2k8vKARybOINdpMdGJlRJ78
A5/eEPhBsghTccUv7hiWbbtr7x/38hIfNjM47Cm7D4JPK+Qtm8qIcKkdqWmT5R3x
LvfDmeqH6jJKJrVKyhWE68lZPpiRKUotGj6ooliU9fhKIxufiv59mLT1XP89jESP
wjMBssM3sZ9Xz5N46FCbdXYb/QHGG285whnFIyIed685gNB9RKvpAyFy2Oby0jYX
DBwJp72F7tB0/K5aqIW8qmrV3z/dH9ZJeqFbczKGd6Dz5xTZZirDTCLK7sWOs2Tg
oCn09rz8MfXfkQSlZ5BsWiVjYfPjklE2r3TB5tjHdBCQ1bUm0X9f8vRX99GtX9Qf
sTv/5YzqH4RS+RigRKVGkqBff+PT3WUolFtC1H5n0GIOhIXt62AiFZNGvWpMKRBL
NqRKiu4v6BIRNfSWHiibkrn23i1j1nXnfxkJbAbzx0e55pwsKrP2Iz92uMQ4a0A3
Z68vwb7yS3pzUctlpaixwtMipadP4VIfkLU2pw2ezIIg7oVbgWCkOYOFG2dmcAnC
DBeSQzjiv9tNyqY3+YxQnqdXWswPMq+E17QxaMthOMf5I7AcgDzFcV9ny7aOdAay
B4/xPnB3GXiWddm/+LcGiRcAgbo0qorxCDTUMiex9DMH3Hrgz38bqzyTU04jd61E
fDZ/USugjAWOlWsCrz8Zrw1f4QddW/pTvtITZ7P2tEaQ6IqgYdckmNDFYljoH6Yg
LaMz+0oDA/AVndO9Im6aHorpw2+QzLgVq+ysmfyJrdaUW7mJf94bUnyikBNmcbP2
5mn2rKaeHHsZ59+pD7DggmwF2NYhle81aROG23NpbLhRKC1RHhJqzD2sd0ov0Ywr
y019THWxfVW835HuSXptjGLxBMIeRE0W4ZHQ/94hR/83mZveGoQinqtWagRvn8wl
8sW5fZga6nvDsMp9zVG8E8qGuIJAl3hkVhsWOE932ZUQY7y6NJGLmtgH4sZ4gdM9
k++wDRPeyYpqP5AViqUng4rdzcTI5hlmk/y0M6HTjpWnWhJK5JIwdcYoVrTVeZFZ
+LNIsRrIswviAOM0o1yvNmqmRP9AT9buxKgvv7AnQvUGQtM6izuwpuII8FWyqVoq
0AHdGHyczVSdat8Jo+zJ53KkXtn13+0Lcqg1yn5k3GDcst8YE/aParVww8f+x+aC
8gmyG6joVnrfw957vWUJS/ezuVw/bKdaB8ursWPwO2i2jqoVg6WrisHAETQzK5pa
6fJJyx5yMWYj7RS1u01aF/OMGt3sKIlGglZPrIKSs4JcAxmEhhwtDKnp1QIYhe1L
hwDNpKuCGyl9jRcf1c9xqNHg9nMKT22fJd1qPBnkTkVPRppCjJkYwPDuOCutK2aN
gcjRiokqoB7FCBIMrzFeC1jca9QaeSSKHSOMTYuK2h/WeOO++d4J+km6GztRAL4K
AjHG6FTADjp74t6L32JaTRAZCannoz05lQDbUWF0CREmNDtLVNTUu1Qm0k9t8ffo
N7TBB4nlkmRMerxNMbCqoAmP8sGkUkjyTcNRLTKQrhRDu4AJbMJRr/73/1xE8+lO
zR/TFMV00aM/9+CRvExx2ZUPjD+dN4dUs3/c6p+6MKwUUdISj8ApGgeC5McUPEeC
fnECqVcohsU7v8NIxIhmcNOsxHU7pTKxCGLxmilQ+WWvLHD+IGtT2Zgfh4M3+Im8
8CpHwhCPDI7rEebCiJ3rsf+QwS2sYQYAja6SCfoYl44wTqFumcfIQ1HI24PMO1Bq
p4oZ+b5Uh/GLfnIH6bU7FnT45wQOPYrZ+cXMYcuQjFfYGdkVd4QteFU/AHWK5x6U
g+7VGnWSYlaS/TRtswp6ylq02yBtpbFN8OgM2iYEwWXKB1mgv/Up6FdaEiJEfr0X
qKy29E23L23WqcXwgZE/x60eIeJjcgRT/dXTtaf9/1DpydzqKqUK6iUkpglQOZdg
1AbSY+rLVNYZgPZubf/GevmLcA6XBw76IjOlQL7WKFOVK1J1oFJYS1qPnK2qp2/Q
J4JZE+9M6j5ByBaD+dhMdthT7SKiSJfwGCpvP0tHFkn3PPUGrH3hOfjinj9aa3VO
a1HFoQRhGm54zb5h6wBgdzjEs/rJX/HVnYBDFDuuUpG+ycuzI+93Lyc0llGRjwjx
SiMXvGZrCrEz91CtSnu3/n9T92h1voxwXs5CsmKY8oNHxSe4Jas/qsPXYsoSO4Gy
kvF25L9ATWumrl9Qac80+peUuRXSUB0iY8PRsI3Q9Ybq49tvpTg54ykWuAuoSWew
X5LXtO802JLe31bNtn+QQnpJul1AEqDqX8SMxOX3+zGWuigbKdwcB1BL0ocPykkJ
l8U85BSR/v/saaeJ3eLBCWNRHVyL+lzm29TuueI6K0/KK96DVIRIq/yuu5RM5JYh
ZLz83r4KIezUJyRf3+L0qHm4zPVx4yTb741Z4acOVjlCcWMyFLYEKQ5+JOrG7ayd
q3eQVfkVi8FCJXgD1WMP5Q7ztuTeqvJfryXaQRzwC4Mpqi2C1EoBtjojcVYOJx0b
P7AMwovVoNrUnUbtzVHWG5XBD9nB86yRWuVMSIEPKaqWVQ4drHepnKY/D1y6CZY6
SBTJIGXP93pBmMyOC+erVUYOM5UxrSIEiPz+h7Bv7rskiQb0e5zMuGPgcHMtY+fb
FlVCDS1VdSK6/8fStn99sSnGz9jrTtJHRD8LST3mRdZV/R8PKL8IezQ8ZITPp5Xh
6Vd87DSNRElPsQu2sY5z0v8fRsjykcghscqFFnqAWztFVP9yRh0scVCvofEIHDGs
x9jwBNnlBRhCbAnwGlyTjC5hBFflH3R2lz5j/AFiVbBSzdpXognLXF2Rm8bFMOVz
vZZTonilNYklRzO8hHhZYvAKmuri9xoCEZHq/JbmBr5VtE5c6FDGHcWdaDs9P9Wi
Xumy6dEkIUXhi22zHAQT+OPCG6B1GQCeX/TzVG5zhzH+USI7bvmPYnAQI3aeyETj
64EuqzD4emtWadUb0qrqKYUTHAi695rxVnc76smZA6nJyqRBYh7GMXL45pTvAT6S
gk76EppcFoppuyvAjTTpqHfcO0q0WzdnK2UEkmkqEqHEPr5UyPbLHA9cmt86R6K3
uWAnL8+rh/DdFmm49F2RLRT/3RVA4iIlmN1Jn7L85MIsYWNKc/iUSnN722Epspkx
ykr5gSkCf+u3vWnchn+8gVLvitOvQXHfMLyssLU2QZCbAymIrkgKmtJ9GJFcQKQz
/zg8sRJ58zZFPm9zXlJVyw0wNZmVFqON7NSXkPaCuGtTPDyi7vE5DZ8j5hXuF9dW
4SEjvGS6s+7Vft+9ppP8HcR9ZosDu1M4FnSmx/ybaT8iMiIcYpcp2zhBN681+VvZ
nfq6xAwfA/7cbYcgcVsfItfj8lb/HqbNjAZNwvoO+b7psR8VfOR6ztq+0p62RqAa
K+oMz2S/1Utq0vpBnO6C722tqI5dwfH+1xCmuq57hl7gI2b7lU37NcvyRouBxiCJ
ntHY2K5pwFJ4FfDlTMu/LgEL7UXYAUU7eaiJfX8MowghJz5R3xn0Lpb9SPVxVH5U
v9OocKnyvPqmYjhxp/oBQNLIrEh3mMC7huAom9ZL95rh2KNAvFM7o0+67nA+Dcjz
qof2WKWAc34Uoz3x2tjOYkIYfy6lSYzSPHYcjN1qWYzoHeVFHHPRK8Z7JG/6aloz
3TAx3yl1mhdn2svgtHZKrzy7YNxb3eofw1oE3sxPQZElNXc6DGL0ilC2akl7O550
OryGoDaDpz6B0NJ7PYm3wJyGUPnBKqHl66miNroTh4TAq0o/PG/vaTtxsiOzLpK1
FSblARX4iugEugMRvZJMZyYJ5TVN3b4gFoiVp82sHwUm5aiX0/xNKaVNVVuqkfP4
FS5J3rOh5wrZ2mSF243Cc5LsUYLZGpQzmgO6UHjhGY23YNeDg9TPBuNqhdcLpcnH
tdxqEJPP3jAvPRwormMcCHCb8FXCzUxyBAVeyy8qXnv/jRBiUiMB5R+RMykV/qo4
fbdifRs9GYhtdaveEEmqirJRQelB2dp1KjfGoIJ1OcDvRtM70pTDcC+aADotuZdA
mjURBO78j6w261HdeeqtwvcfI+Dc37NG2NQNJhJY0G4eo3zicv2GwRlV/XaWq+ki
ITWhLR2rfI1lI8IN8PSCbAJQHLGVnIP8TKdZxNFfVCJ5e2OtUMqCLdTCazdcRu4D
bujFAoWv68ruFzgzLtNxEh4bSIcu4cFVvgAuNurfFqikcFe6p6OB7Qw+UA191r/u
laMX2rayMuJtKO+VCJIsUC9RqRRWdDvz/QhuYI1/W7DFhi+BQA3EQeaMThoRZ7Is
snrNqNHfb0KmdhD73PIwe9Vn9eAyq0b/zdHweJXcX8TiJcLbEwkc2uUUd5FJIP9Y
fCi6iF3AJEJZlZCWMGVUBNPlHEX0SZlgI1vvn8rLgl2ql3RYFsWSkStit15eZGP+
a/fSydfdvFiJdJmAOy/6gZ6vs+CFU3U7tj5W+31FLbB1WzJx3cNWoVVTKEuuwml9
gl/nbHjUXUJ97G7k6yEgAUZyNmK1MEDClMue7Ib3reYY1tDRCY1tcT/rlTKMmSI5
R7HI7c10noFFmAbhJQthZjeJd04Pa0ugtEvvq0frU0G2+7C2lCHCSB9Z1l/u6lhp
6miexMC9yC11YRBluKOqgc7cIqKBRFeQarcMxPmTK5L4vHLlj8zkZAJJ1fu+vS6Z
B7AKoblq4r/wcUPX5GqegeEd/Tsu1IyYfletE/DmqRheL7idB0+PsAN0GXrBOwW7
fgsmXeAIcNHPizAAncK46ublKUbd1fqyvdVTlCzKrX5ukU52lVVJJUvF3v7Il+Ng
D7mVT/bdaXrSKWVPNgcdrk89ymOQfQrkwZySwZSpvd1MDOX6K+0fwk9l0LnZWifc
kDoKXNkdEzsMpJVLc+5RbhBZUDn0u1tJnasSrE3wTZo8mzGFYVlIK2o6dOLfCyT2
YNbBB0W1VkiQs1rbFshuIE9Hs6BDF4exHjm5jMdzGCNhB0ySuX8UPcimKHQpUC4s
EIpJSBNsEOP7U6KaLJSHCqpPT86+OWWn7JsTTMUzkT1QI2uS8EBzRXRt152BHAKq
zOMc51zUy3RXe0GMbAtQndE7ZCev37cuE0jqA22wlzwtzgUZ5x5T+R+EELOmjF3j
c6j4o8NyscPJL3UuZX8JKCqYuxE8kwNBRHhbCyEqccupCSQ6XVGHH+UaM6wbOSeO
d+5O9nogIdL+0dTCV7YlWQPzS2f75t0SRoi0VJr9YyduVJDQItUMJtHWRO76aCsG
QERkx3SKEkpFumdc0AfOSz61vTDh5lPa3g5CJElFjqXNYcZUyE5aunov9golp8WF
bqtGv3hzBcOw1jtqNclQEdszmWc8ox/tfIqWu01hhGjOIgscXecQW+Fo6DRpQAyj
J4tihclaN1o6BlvlretDir1bBPFmQdyb3/uP0NPDsbOpBHJO+eLJK+cSmilqxfsM
A77BKKneFskYwy/HW3a68xUKEgKwgfAqJxU+teTClI7O06/Q/YBHpXQE3QgPwEiB
NPLwpU2nCcrg5Y0snFtFIUaXafkDORqPXEJaXIjBeMfkZv+VD4896wDtu9aRd/gS
M6P9O3vhA9BHPwyWN5FWgvyTERzdWxOPi4mDp5MLkk015GTA+g2e+XT//00MaQgJ
CzkMfKjpw7l6i28r/7uIGn1n7MFFPt1X6sClivYlfAYNMVookqjUYm4x5h3AGgor
5UO3c4Kbi2i8BKYBbDO15WQVzVlTGGpEC2imPt0HtwokvSOB+7e5AFxzGJFhln2M
91Gx1whFZzZWYdjxae92Kac0qmDaL4hbiooksM0GhMocdZvL/NCQdv3yP7f+OGlu
lQzGBCyNVaBv/5upt/0pIOinAlBOrjvl0G6O65PYmrS0MYJdCI7YlCU1shpexD8B
MLt17aVbzxSN7R0LDbDXca4Oth/6FUoIou+rVaeeJOYYeMFlKjXCw6DsHu5KRitm
WiC0bCL9OFhnxClvNKCQahOhOf9gPF9UZ3NoLTFNw6FzKiUGVOp2h45xLgxNV51c
rOjK/LPKcZYDfgbw+tCZNnGLhLQM0yhPOLo73BCR+7sb78vLlg8Ujxwq2NghG8TL
bfoRsdxUIiY23I8yC+zboc952sJymocsVNuHrxgkGQ6SxoGH3DbmxcyBLwABOv/R
1MwmjdoJ0zOjrxtpC6Pr/ygEXTvjt9I1Oq6Gaz1HQbjOF+ZUXlEd0aF+0i1+shIU
kCis51TTd1d8m3TNBFkDQHtBC6Y6biaymcBuTl2+1otXYJBZPe9rswItKD3uVdrB
rZJyd3SHnqN6lF5A1zKaseZB+AsD5xyQLICUq2ThYByWXWBgeU81/SZmhk7XtOri
AvqiLZeBUnHssLQ6DXc3OilZWmaU/q2rlTrOm3b2inW1EgL+XL5SUdn6vB96dj9v
6Q0oTkjoS0BjxjqTSV22qAoyy9tMJ+Kq4v/LueFFBrv+0gB6nWJOCsfTyjln8J+C
0i0/1pFl1FvB1ud8NU+qaKayjG+j72iqljjHc8LLSKEH/L+uMYXj9HGg5rdnC6S1
FcRC+bmqwif1aYFydfoZnX8R2O8VUFOgyZwyEj7LePwV0wl+5tbep6ltBxSX+HmZ
o3E2sUAJ86RVTg7DWEOgHXYOidkOGoXbDsP/lOAGxLyiYK/XE25FWbrVjARATxwk
GCoWeVk79GaJgzFp4keyR0qvZ6ud3cXu3IcDeGPRH1M0WawTbbCV3vm3j6sFGuig
8vL+ErCX78q+lS+Sd55F0nh2+wB7NlsBgyDSCW4J904xsKYomywqO9r+axFrnaBX
TfeZP0nX0Ln6RrrSQJWIbpw1PujUm87GcHT/b6SeHfFV0XWuZkqjf8FpTtiIkk0p
tIP6aflbnYFqIhbuyDagfL7AYa41zk5tq6dW+LNPncU+iOaDNJ1nq5WP59jnRTaD
XnQwzlSKwCkeLKLuuVbnSfF0/HIiIU1EdoFBj67S+GONMqLq+f9dFaNWa1BS+x/D
dmOcXYC9BttAjvIkfFJ8Ssq1BV8BWM+UMYzmJInCP+wa/JpqSvzb8/Wh3gGOYdKI
h+KxGljuNero+k532y7eQOc/rLpM64dh3C3q46B7F24j+9OlHKRuQN6ynnkLGHnU
HfufFWnhrBprE/2clnXAbNQqHdysOFaYJ9vMNxSVghtqhK0qxHa10lmnchBD+giI
dzqkFZpgGlWJmVV0Xc0KuIUC/PqvImvjNXH1RhUwDqlPoUfCZNQNhSHszQVvQp9N
kmxvdgtQLZInF2w04JB2XZ4ZyzatGLOTIYZo9bkmVAV54iiTBwG2qMSp5y/A+ms4
1YKFbWUZn6ZKtadZWyhhaKypGWy7nd9n+G8vjN3PxyhbcGELsFJ1aaNuzr1hkNb+
ipBcWE2rZAUUPAdS2pnmXf96vHLaR3diFE9FWNQn6njEhKm/kxJIYT7T4qEp2W0e
ceAxUtAYKj3FgZcCtULNMSINf4l15+yFJiyYCPywSnO6VfEDz72kwqrLYSPedBVk
V0m/vvPQxW2+HAq+8PuS0MhqewrDHnuRZYfrPFk6SkPLSn+QDgTh1krPFJgV9nn1
6bzhkwTmyiUE+7MQJ/lb++Aq9pXAcydtjGK+svmaY39/Yqq26SaZd5wwkzmArnj1
Cu/PkOqf++bkFXAD83CX2pEpsv4g8I2Iy05nK75RoFDm1Km9RJGnATMb53R6rBj9
l0YzmrvjfDmQ1jBnXV2iGkftmZ4fUJmGI4NiwMvERvroMF3L9VW5KrtCtEgTkxZ+
qrCj4qvSz7qiFskAVQhyXg+ICDkkAPkrYt25VkK8Ig6UTzJ0ZOwe3n8ecBVceB5x
a9mCjjdQwbdG9ViLU9AVDstqIYIfFMDqTfj6aC6z4PCYv3m2XOU7O1BzVY0VnxGr
IDwC7A5Tiwn0wdq13yCLIBU5/fZZx+/E3IeGZvgaf2kd2ggrpfMxbc7TMz7TpGcq
VxCc7BBZZu+6XP3BK3SAn+t8bAalOUx6m6KnAgZJD3CZ9VaaH1F8/SlY3VnU7cF9
VRJdU/8WByHnepbU3FQBOVqgFan9amrZL3gPYU8LyTXQA6/QHV2W2N7A2nPG7HOF
KtQNn2Ym5YCkIk+DhFy5vjwRTSgccDiBV6MlfMBHNRokzV5TPFzyeViIh1aXa+j6
HU3fPCj3R5hVGwG9AaJbWSSWiXotSGi4gD6iBKYFZ+pqKeQKZYMxRxFHSSlBjPWX
MaWKDyoCV2S0scYcO27FzGdXBRBwQlS/DWwkPmG3yVbYWtFWOUMTHI5mKmcFh0HW
vKWXlghDDj1KiF7i22TU59+gLFPpCy1XIfwsFewmjEgRK416RVMIs1sI4Ks1ChPG
WViQxUmIHddwLrHyhmDkZPT8du3TOGl26ii3BLPGfrEuhH/YIHLhbByyuW/pl3xl
4gJNnN4q3yFwX91PyrJqZEtuHbGtEzew3nILgxSkp/I80sBfxIqZ6mckkW6KIVSz
/kTnYUSjcbZyAWSHW1BUkr8v1xqygS/Bs4OORMxxm2rQBS5RzLKFY7YcgHCRYJpI
m56AOCHzZUKo8yON9+BiSmkAE8BjNMKBhjw1UKWNp4fXdCZU0RHgkLtqCihBIzrm
fqEhT1FDWUcCPBvUyY6I+oDy2XzLcyif7BJncUTuXAUJ2Yurw6rVXBZN1MK7NpeE
aX93VZ0zfnn7FpU/Biuv30+kTLtOsadCgN2rX+eUxdYyiXL2Jl6JexqqpHODWmqd
NytwnKX2HLaOhb0Aos5rn2GpwcAgnhf0YFsiqAegDUrjnwOEwn2XeCHNbw7rp+eu
7pQgqHPDmEYFuzPqNKCp/Sf4wq9tBkmueU3sFREe3SfSsyeGangGw4rB79hoCjFq
pcU0x+5IsnYZLzaePUKGJRimP+cSPkTp4nBqjWi7F3jmO9hhTAEexo61cIAdJd2A
Au8B4lBQZlLrJLFOpCYw+ucrwCwNfPLdpvOOBl9CaCr5pg1Drv/Z3xaWAaISRcuY
Nl+vktAyTfjmMeQ/8WnryrLHU6/p8OjFxzm/aDgaaOMs4DItho50W9TPE+4pd0vi
2MUtH72gqhsa72A8vRMA95pHi3aqKxayibL9GPQxPvf/WHnteXkK4dpLUNZkvXsq
ibDQ3bIaGBU3in425QLqREb5lMb6P72sh9q9EO2uBkX4mPlhPYelhB1npNuHTEGd
mULIfpd628nyo10QI/VXGOhXm+kxdsDBIuqOYcAb/Mr7KUmUpNHYTChITIqyNtY9
s8C6T/CF4CD2T/H8goXBwHWR6xwAkokFF/u4aJ3eN2/Nh2qj02RbvwVP/ZhWB9z7
112Fj85ZKfITKAZirvwI/yTgppz8YwfeRZn/xvSlCwZERLhpvnm+VDW6x4aCA47u
MSX72bjtPizFsw1ncOw78ZWY9iDfhWA8aqnrC9rercw7+RRkjn+cwg/miW7XdclE
+xWUT9SEpIZKX3OAR0OhlP3uBrolgu6C2YltLscueFY/cthNdKpzU2GfzQZv12b5
zUfbnqgW7FpgkG4A9KAw/sU6kQULIfHcRzm/6pOe/3iGNX08m926FRb3TMe5E/6F
uT+/QRU7bYSHgsg2WLAaWneJdtRLaqnBQhFIP2MNGBOgBtm1vEhy2NeHWfM7xE6e
N80tkxAy8mEQ4d0WhgOg5smxp29SovsxPdpe5Uyf8co4LylP79BUlBpUAs0dUTu2
zWoCZfXak1DHC6KtasxbpjEwb2nKJfpRBUcse4p3Er/5Bl7nv83qgJk7ig4kmiDy
oWYopTN95NCHFr0mWTY6N+R3W4/lAg16RdPeFVeeLKEOSAWn9vkOm96HA5ws6mxK
Ib5XC81+YCCmnv6sBsatn5hT4K3852dUNnSvVq3nE241+Z0jYYZ/vDcJjcFwdDoL
jmKv3M4G00Rhc1Qv1097W7vQvsx4ARFBYNy9mrya3mFncMBtVK1mjAPHJWofF5D0
kf5NcwZtOKM/eG2mGawpQuHN08QsyvFefi6BbY7KDNe2hZHKtHHLJeqKXhKDkWrw
stKyFBRnXP2UZl1O3B65j4bwquDoOUj5XbXOFeqAEggEs4edCVDfgCIZcJaMCSrm
I5/pqeCHr7Lcjq4r39IGj+kQkPmVLFL5OjSVKkbRfiGH2OvCbyuRuS+H55krgvYy
k+ML66HBAH/N/WUDS9cKIQwvD5WULEGCVSzQHYoj4lozY/V9zlzvX4pC3XW/bkjr
D2DydcI4oBZMsfyg1B/MZKsyjGdi2AmrGi80YdE0W0NxRWR9CnXmHU9Is6pLNhWo
KQPQKtu5daO4TkvDdoByKiQV8XjsiGu7qVGzs+8eQ9E7izdxjcWRa/aRcaE/tzJf
ljuj5BYSp24yf/tuJ0NX1UhS/nR+jMRmOYN6zE9F7/P20SOgNTyMlYgDDSdkkXKq
hfJeIn4VdYaBswI1LrGdbsxDb2/cG5DHqBz4vWp8l7E5Bx9K8BCtL3GnkJ0m9BQs
L42jlG6FtgzKcWFFKSe0z6FRja4ry0ajOFzPh86+IbFlhoqJIulyP98i5Gpbi1UP
YTb/bUa3/OVudx5xOFW76wilSEwGaAJoLfft7U5hl+oof9ofxmLPKgsYyHD31+PT
0Ete+Gj11yABrLu41dfnxrvboxYiABvks/XC3MoF9r6XKHF+o3TU6tAhxS4tBBZh
Hriz9rv972c7Y7jr+qiA2PBnH7cC7ZstW8QddYLvqXvkxQn6DQvmVxG5hLHQQmNq
GZdDK57uWP+3iYNp0+gFDPMoFk1l2R61fu+1c2w9cGt8bNvX3aQbEibiVU7S/UmL
oZ3ApGlkXpkBA2tA468yHPZzoIFWTfXAzkxRgp3muKmq7vPNC9j5cfmrrjA1L9e+
bEWJIWyfqQ9O+mJNCJdRANesDnEeFs/6WHcN8yDFeODybZ45gCuussJ8cRpt8g74
Z415/3vmZiwG5R2bir5SUu7EMjl1yPsRlK3LoseIL7Mt51u197TlH9HtWk9p3ETh
wTSiVtlNflIWRpNezxIDPtt1iOpWMzZIZAeU2Xt+u4r4pjxUhzwYpTsH6xk6loMS
BuGAEOjIzOYTnKCJOt0DNVEKuZBFRNx5txB5beQuYTlGxtAUdLaK3xCDEPPgJS94
+MOfblbMEsHu7rNoC3cPxAisaZoU7k05vSlVYmnV1LvvzVi+Cf81y0ZOXit+M49G
Ve3Agv7ky5ZjG2GTQCw/lYYBLrfdWLQa7HBs7i2vxgPapsm7TkODR3NuUZCHQzS5
HWZe4CXCh0cUFN75MyQzhWC0u7X1hmIQY7cbf9IaI97KAfZLOKE9J2INniZUrSKb
4eFxwAZJKXakT4+/s2XLfPcR9LctYqJOyheEsMVQ1NKBa9IZcPPyxei/STnDtIdv
bZmDsEF/QvzmDp8j0J3aHj8rjKBU+D8tmKmUq4nnn58ZDLjOxTJMJdSDOipvE6L6
e6ijfy5/hH9vxXc2hK+KU2KlK/Kz7CbW96YFbHOgL8fJvm8SrRTNV5Uqi6fvqVNp
LLLU180D6VDuka8h0Rt/J+ZZFSqBhZ2RKpnJeT77T24F0NNUP7Mye4ejAeuRWKZy
T0AeuratLx3cgh/J4gGF07oSqYIB8C98Bp0oi6vAe9G4jWaZ+wfDFqdByS8sya//
I5ckFGbcMZcVrEeyzKR7Q+3iAh6dkzEwbPie6F75WzawGBGBLO9HDXoh1W++Cs+A
d1JOsoRSJDksTcS3XTDCZeumPYV8PylfBp5tRKDqjwQGJdNMRwgbJLBtQ/VP1bjD
skbRWohAZikVADHzLTqpbNIO6H/C7oBC7E/DBiIBtJT7wAKyIi9B28pCZZs6nw6+
K16tpz6CKrjhNuViGM9IginuOQ8dDIKp21t3cvF9PP8NFW8GCC009lw6jNCGwY8C
gI+a5DKpZ3bfPCeCDGH2SgF8nX0RlvRx9Af8Gk/fsS9uKhs3JM/yedKwpLJfW7vS
eCeNHNRsrwQZXOt4P2JlzIb6BWZofrMTvvFKxSRl+ZAcpMAPxrvb790uqOoipGFx
4pNx09RU8V5qQfVywnOIgk3YOKiV7d8fuNH/rluRji4jit2Ji6Dl4k/CtbF6uU4s
/Aua11ZXq48T4GqxWXtcMwLuh6vtPRG1FsPjYfbHWldVEI1y95NbW9TYm7lMs6dA
4iJDKimuojRCUQz6PBfCaex+TW3RhLoOd6+nFFjk27hGkFfzQwpIFkrhzI52OFwR
jXqoq8F/2+q2i+2lm/PsnVAnamhr/OeJb8bArYfL2EXm3UvgHX2WmRlHB8K8mUl5
nZ+DF6X9WoEV5sMd6WkqjY2Ysp5CRZzRbCgPPG7nuxFGoiJFigztUF3h3/FKhMPK
wNa7vyL+Qyn3OYnJ6auz15fL6T16qPWI5goj/uAMPi/Sf4VzNK7e43JkaUR48aT1
xnwdVaApDyugNaVoksO+wE0EP7KbcyQjJOGEcXkhI9mgMSGwwxf06caB0VZJ7Fqi
9k+a5HLWZ1+oyL3SRXneH4MveEDcovoQFYyx1YPMTTZcw5K2k5bKyOVs/8L3Mtjw
aHT4aSXRkpBzzfdBay/xlUBeV8eF1mVFwn4DFj7/Ditw5g8DF8vIdHGqfdo/YuWV
91VtjraUfsGbp1ONFUPXGy8/0D6X1BDCzz4jusGFCGV/F9HYp86oqFMrnUTexy72
sWW9ShQIM0j+MP6c9nGQqsUG8vNDtJ8vwMZhlRIxx2SziH//9O48xurqv2juRN83
4iZTa88JqhqOsvh4gQdI/L6yw4DyAtw2IF5xpgUG6723pS1dvyS3pDVhQljEOyeS
lfm79yUdQgr/5Htuvz5JVLcG+2ndNyowxsgN22PNwEE8wCDFwqOUP4LsC59BFyz7
TZuchgVanYuegYcbFxxcn1cXEkw/qLYRhi2ZKOLAs7zrAnhPA5gu3400souf9jZL
EMth0QuPbjTcFhQfRjFLEWRu7FUUj6pemQ4rinOJdfAGf4g4vf5506v1Yi1n1HCW
91GIVqueUranKiXvH8LTM6Ugtd+sVMqPqDcxDbj940BO9MWGF8ptTFPcWPhO0hq8
6Q0TnxNUBjejjxDyLx38yxpqnkwIVYIGBDV3To9G6UBzxMpLGMZQ9DYzEzQsYL8Q
gSN2zAhpqR20LNj95B82aRgue/attdLT8peSWbzCjTaQI3wqUeT1pie6iYOEhbl6
zPCxVuEx8RQwItsBcJ1DE3jbr3O+J+6+LwUF5Uvr1aapnXz+i7D49Jg0VOre3wCK
kGqydNfMnBiY4jVlSlNrDC2v1Un66ADCZfi/kIIvBLgHQ0IrRitsj7ZBK3l11o0x
8wXyqx6p6F4uBSCeLLEGNpGDJdZGIv/knMpDloDf/nau+rGVX2D3ughueEgS/M+7
SCNBSDuaE50ZQ0Mg1WyJjrRkjwQFGsM2tPpUwIrkITqxjuYVn6H9MVN6FyeNTfx7
qVMD/zFf9tG2JQGX0wz8uDn/8lhZFinBqLdJ38njeLonds6WoatuAJ/bCo85w9b5
y+SrwwQlmk6PLs/qpOGQwzjo/ZSenGotjeg3Me5D8Uv4aiPeMTquXr0qebpxvNHk
hhUL+oY19cX7MlItjZt5E3r5xHZf3C4dcvqbvnyKqdAU5xtScwsL5IzOfu0Hadmi
5UaDQ8ROPgvIxB6SPo8XQ5Fp16cWf6IDdI6M7WGuJ2MW3wO7cwtpZtsXkW8Y4C42
u6qM1lLz+rYjQ1obp5gMDzXDkA/8c7QbSd7IJtiaHOeIlSGkuWZEmThdjd1Wz1UG
3xFZ3EdrRBVkN9EKZxJZGjkH8CsU3GNzjiLkG0IHQPMtRpsGFgEvDznR3k47HS14
VLpZcsrs/ZwY50WuaoMOCXWMY2ipBhKaKM7LFsEOZb7FRO/GdIVeZWzhXWs1ofwx
YmvJ9uWu9QwjFhDVQ6R8TPeDmZp1OgFpdK3V1VRxn9SjHdO9p+77vD4j8xx6S8Qm
kUlpC4qiWYXYbyywLRiSpaCRzWVwVxITlzcfT+0pdxKPkvUl06QYxKU5rDwzfSM5
+eTPVgfg/NxeNNANpPEHOmpbs6XzZfY5BLZLBXz4qhIbvv4SpuRO88sIy1APq41s
Oan4aGK7OHFTI6LUrdk1rf8iZfWB03AgpFk81DXfi3W8NFgs6wtHrxBC/jZiKW+4
df16/4GYI8BiWWaQffdzEifnKySTP8tYsLUyqxPDm7BkFO8w/QyZu9GK5ThZ4Evv
G19xLOufryqoYNazbRQJ6eXXfJ2Ctc4LPsqVDFsAEvARhPCnqfAxT/OjSYmWp6UL
qvxYo6ryJx3b7dcJdEnXjZwHk53V+sy1rNvUMG4XI4YjhWs2XnNUyi8fXwrb/Czg
N71QMvJ5SaHGlGpFm979y9SGqFZMJ1KWyh5jU6q6PXSe4Y+0lCvZ9awESONozBMR
eqUVgc+5kiE8EKENUHT1xFlS6Ptb/EMIjixv+xbDhXAy0CryPHKZzElCWQND1K5O
ZM3KYZt7b7U+93a4X2Nu3HtUhVD2bKnv1DsY+i/0bPMzW9gGNfglWDyXVvkEbecK
Qp6AK+3/bTqEvOY+FWwzV2PMbyaX0dLKTcTRAprqSwIYO/j72arOKHmoJxVCE3Qo
sEA0QgG+8w6vgl7gE1jd2y9uSTZ9ao0iAFbYZgQFVPhTgX6NW9SIiYrTYRsOdCE7
DN7tXsnymmwIh1Xzf7LyGPRjvYAcE8MH/I2bEB5cMbxJbuiVBwdxO4Kuv6KJWit4
8QXF9JSDGKMFCcud6z9IbVFPg4HURVQEGFjERTQJlB8LuG3ApyCbL8DCu7lG7Kkx
C6yIHdWyTJ9fCAcYE2dK3ft+KQ/hC/K2TY+hSEUoa/Vimy0ieNsy0bVzU9X26Pxm
D56hliPXWBqdkZHbZwPOxGvR6V2rVcYXwuV/rl4QS5ivaAUQilnGbNCzR2Trz1v2
RmAttzmLGoaPkMZPtncqzRY2a0ecz7aNXuc+d8bKJuXqBNR1qIoDc80Dp5SAVjsA
xwXwSF0bt+KaF/mWexJawYx4DtTwznVfPHD9WWcFVjAJ7NCyI+oooT0Be/oZdzXQ
s572qTf8UnrnMP+ECN0RxobZuj6PS2dS2mpornRSldO0O3xZdSJ4mcv/LMiNp+tI
KFhvFP9VX6eKoTabDXv88py7P4GuIJeQlvcREG30i36BfotnunJu6U0wf/+tWlmQ
q1wYGKWmca95WFFk+EuqX23Y5nNpAd08mRBaM+IKjswKBZLtRI+w3eaJh3K1ASMw
RafV1yKBHh3Ii6867lVHPCo6iPveLNNtyZMuiUSaXH3b9jTCoK23IbhXiI5PB3o+
Ldij38sSBxBeOBAwnMWD9Rwh9wRQVq+UrWUh25AXZNEp5FK3yHNncjwOn4NxNEWR
DH3uy4lnJWIs0jzR1Po1jFlX0pwT098VW7jzX5YqB+dk1fhIN0g5uxf10nGbexbx
7txJj+G8dhf4IuVft0Bgl7zu1FFQdKqkg7E7DctGBKdTi7K6YVfJRfSiMcD0QsKh
a67Ae1BGJTCi0aaeIfkScPexOw9FscEoJAItC5n7L40Xh2X68SQPT1QpyRZY8Mew
fkrLC5pFC8Zx71FJ/9fGXUfSS85A6RHhnS/8AhEUOqVEQ17DRCBKyaJ+j9t5odtG
uPz9SxPc0hfVmn49QJME/fc6l5+scCUQT8EJ0nCvk7lPwlitKg3m2Wp0i7NkyW+o
S2ymJdI81beqZSx8J1alFI4zYY2AHZvDYVFD0cQBydjT/Jaci4AtsqAPIBHgX/kY
oeE/DPBnsA9FcRIZsKWfQWD9glHHEN/rUeyT5eF0vi1E8CIS91UqdHysnzX6DSN1
o3SNRCwKZHcdzgxU/i5s51YRbXHoZWqKSCFczb0ApxLICQ5HP/NfYcwB+JQI90Ec
ul3Xywc1KvvahNhTHjJ+Hghswu/pQagyV9Oowl4f3ZijOrD8UWQlTBa73C+mN4yQ
aiEVMGrU1tfQP10MYwdOM/V+G01gCvGriDnGA2WmH7lidT6dFQrnZJPdW3a1mJeJ
EUt2W+Q2KzNDgAaVB+i2cBjaGQ4N8oY3/v9zMFxVg1ZVbraHzI+EBYIReiCV9Ivq
cXIIRZ1L84+AG7Lmnrf1niLVdtXcCt2OSghGevcDaQxaWlsr/LnCOG2BT/i0ZDeD
fYAndDoHhf93zsgucCSAP/UHozg/VBbnrVpIgrT9WLHzztns0QCitSrspZfvQtUF
Ak58PTn4c5TBuv+f0crND3DZhVSZDqTwxApwc8a62PqtQs0ousD0EQKctrkNWGCv
ytSeer4B4+aCvpD/Yfd64acZTOqFGhdT9z+fvyCGZacdxlkkl92eYNJJJkhHzmz8
i77HYyEoN6DfFZaWjw6TbAHQzyyu+90Pa6aAJEsrJwWZRJ2GcDc9ddSXM3N1WU8a
SMlpXDVRol7Ot2z7cIrRs+KfEco8EdwIrU+9WOZQOdV8Lx5ZaV9uNXJPoh2DsbhP
tHMjWcOMyxPHesnTNgmoHsoanmGcSw8tjv745VU2pGK58UWJnrYq9A4Davw1VVvM
ITZFtHlyWXpn9PgQvu3N2FJY2+E+WtO9pW+z9get1ZqF8HA7DYp/55Z90CwPxohl
CFjBmgtpYL/zOEXprFCM1s+hkia1S4D3bBL9oSpWM5/mJEHgtnTM8SaxCHt8CwnM
r1L3vYLxRtvRwnIG2hLzfaR/kASchyxytcZGMngbX6BPH/tedQ7H2E/RV8j2tDix
y/m3nWYvKoOSmqHsL1hhbRN99+LjgvXHlPzCnu+Uz6Z3bGBNMdzKej0L2Xh7NNk0
jm2RKKwLqqLwm1sWo94zQZNd8Tyu2QLZkBX0WrIp3yf4TwtooMWMxrdDYR005btg
jP9C3fYzOCR5Aewe3LdADKxKeJjan9PUMFjEwMMHDUqTk0SLDVVAYHfS2Qavvm+Q
5fr7zbc3g1vcHbk+etdNslP3YS/1sx2BaiQYQQN+y5jDlt332V1AyeiCXLQTK31g
aPKY6UAXG+gOSZrzAcQqew5L5qC7/f3FH82bw0V7v3MAR3GbwHis+r793n+YU2YJ
ckbqC6oGIsaLfpPlcRTFWDleNZDTuRDPdOyi/7mnIjLRIS3u4kqtAPC6mtQuL8A5
GM4l6TzNMYzHo/lnXLGprn17tguH3kOmxYKcAc3bdmORLWiWplenFCNalcBKNRvE
XBYXamRMT7Vxl1ZS/DsFxhiXORnbuXtsdwRgbWZOSW9cA/GFti2BUs6v8cqllEcI
t6w63fWFTDUIPBD5kC2rHZUj9PG2MznxXyTziIHdJpF7KUINKWqqQL+xFtsWZD1w
FM7D/thheZRnxLBNQNkt5nzzydiMygqs5oArUID6JuY6FAqUCmqBb2RA5IYetDgW
Vb3GJIt+hyRjYlgni/UQktbbmOdek8Sptg/zaGniQP+ANI/X0KyXEEGrVHpNmg05
LxuUWGrBj2/uD+5DHuGtHDksm0usKeA4HJQSV1aPCGfmx2dzbYPxmknYkyi+4Wis
gmWgU9gkn7YgcSytG0ZlOeMIqsi6YeRG91Q2oMgwO/uftvPlUUvSusnakGFMnt45
KEvzBvobzpu4jJirS+QlMaShiG2HPDk6mQE1HncZShn0XHfGlG+WDKhcv/SbjZJa
k27DyjHVS9kN/ky1Zkh/av5pdpakp31GUdRVSGFqiHpgR2aQciGzVUlICMM+9Bxb
XwwUTA42/F0ksffsmrl847bEj2K893JPXPTyuRT5TkdwTHWDrG1Khwd6ouMhI9Pf
9F1hNm519XMJRuzqD6ayiQM6/Tz0dz6320dkDsAPwydagf9oOzZF6GBuAXns4Ops
cWkX1/tNInxf7yKmjQFuQnoXuCf5LP2S17RObcI+DONc9ZyzBytsVMkBuB5bvXbP
79zPvroJYsZzqz7WySNJZRjq48+VPtogOU5GxPB0F9cbELFOhzZeZVqNvWVClJpY
HJsoYD4dP7Yct7q18hJ2qigf0pmMX4S58k7GMXOSiO09X57cHMBmSeMNGFo7VApp
IQxuZohO/wNxR6e/o09VUjej0oywxkHsz1EXlzmeeGOtVHfdy4wQnY27B1SQ1ehX
SDDNTQZ/fqKbx0GoAvPatRbN7cIHYKO+UivRJoHj0bzs42Pd09JJCu8el3pPU4th
hVI5WMhELfnkz0W7mm+RvVV0oWCKs4iazQLlAI7ZCbHBBPxJwF1/Yvf4W6yIZdce
kQpWZDwirZBCmIGbkMMui1aiXjf1fcT+nAWR9eBMTJQYKvtb1pGbzp6BedfZPjix
EIPUyNbEZ8GsRlwVY29usMpTkvNuirM7tFFChsVu4V6E30LFFPAenxron3Gr2rF8
fh4MdOSrKBKePHoPr39p1LxeNf9nC8izyNayJU5cqbL+9YXUkunn+N8FMzVh8cUV
aJgjlTUf69m83ppWO7LBlfYcmbxV2D/GfN3tKDptkH5lpsljXqooG8zhYPrmLKOr
BO0T0kfBygyrpafYA6DGK+RLtruuLSA4EZPr4mLm3PcQRs6WtmD5FM+2iWPmFAwP
BwLegzdILJvAHTw77Up6PG+wtC+WRFti4vDEgAk/IAYQqQBrNFNbV0fuKhGUSm5B
KMFjAR9iO8AaxLmlNdNtFf2UXSO75ofivzJWIY8+fvfEa2nr5/rol0eVQFd78jJN
QuWDb9iNRDzDWxgEi43YqErb8t2cILDNHmo/oNsIZo8Yon6HMO5foLpzcUFsHnqR
HDvp/2byClp/Ph/i4ZkLHmqrq//nFSi+Poq9FRK8H6+cIjjTLnRCUYeKUVa3+wz+
FDMz6Mzmhi7MahAdythazfiExZd25LBXZoOQwjlzoTe/X05VBtQGfm9j2lbOiBjS
3mKBTURnNP9DyQwuyWO6k43308D5XO3ecqwzqbT+pR0xIcc18qOAtb+gJZkPYZ/H
dirlMKdrah98thqii1MRCDeLOOm2a+SzdGsPPtlIKr7172DtQg8klgjjbY5uvRYo
zRjk4Fg9VYtcGTpoSCHfoh4ekW01RMPrs9lKOsZ1rUWKj0UY6jch7y+AYrxzk6r2
KgCGGgoFalajcDN71n/SuvSVi9+zFM1MdZfTBjQNnga6mKahm75h1hPM4FjgGYlf
BIXSaV8kcu6xZiJ7pbZjcxeuXDNIlpLJ1dbWkP1I7NUFoLp3QBGNikt7z+qbJscQ
U6JT4O4xKlD1PpRbknhyX/M2RrbDFAOw9GLN7x4cDURDfTsiNzo/YK5Nrx6Y0uer
6uUUYCjBI6b4iOv90V2nlCW8Rftig3ClY5+gBDYqaXgNnVljo1jOzCncEsmL9thy
tu6lgL64e4eryhlfw2nicKYhn8vb6ISGYh/HZKTCFFsG4oXELjVVycK2ZBoAtjSe
pSGgf0zOyQjiz3jspzC5FyY827sJDP3NneV5Rl7pX56OsPbkIU/6Xczs7ShBmNhU
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Uc69fnMkmPTtSoLllFU+5V4LtMjY+/ZG6C2W5yNQhdFZGhNu3QuXrJP8Zz4F2PLz
kxDvWLlHnWWtbFa3qnSCmei+QUWRPhTqwfhaK5H3/mGq+DST6cSM25SwEUydne52
HzdC57cmk3GUtbfDQ7gxipuVhv12CWLmtGQtK77EUIx4vSFieJjsaTWNfbQ5bVYk
oo7PS9WKpg00c81NAakrukBTLj8x3crTthJ2gR+OhPJEXu0l/zjtptAvIOTM9MTS
qQWSTfPuRzraRt+U40YzbU/q1bvzYWD7wavq0cXXhmZ0nC/ncX5rLy2Aj1IfmfNu
GlqtNor7+vaj7ObkeYFoCg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6496 )
`pragma protect data_block
8Z4KoLXGKwVe0wCBKj40Q0z4eeY2ryFH094euFy6j7SQj1eeL/zJ7DnEWtEtdXKR
fpa4ZLkYuDJvGUG5p2lv4ABalVdo7Uy1mrssbs8lMfdm7wW6wXjsBxsrEXXuDuHX
IPu7ryNyOXw/ELg4DQbIoWgxM2urIv6IdopceVQbpQGnTG2ha/hwAq8/atHliwTc
jdM1O48GGTzaXK3Jd/6NOgJfEytjC80LGIvQdITPDxtDGbuNBZI91NSkVVxBibH1
INHm7Yw6b7OwzZTJoFOwBrDKdf+0Jk4WLdtbKPa1KCpRcRjntqgjNsT74d0wtQbV
HIipmu8quECiCUIg62wx1XUqIQ7AErYq9O+dL2tgsnfsWzX7+UJ1zMOJx/L9/J6U
roX+TY5xSuGEh0R/nGaabt65pqoEYGAVGUySJoYC8VsHAW+Yds9cSdjgFm1fWwo8
WzhCszDZHhKrDXshmxeP9CC8LS4B6MNbfbZWCv+4+DgCigknzBee4Mb8IaR1LgCO
zIZLAKKGl6XlUThttkjgHGo/40HRyASfV34uZPGHbEJE8imcjwbowWOrizH5XY5Y
IH8xTIMVfCu9g/bjavX894KbWNsLs3DcflKcziJkD3vpGj8L+Jsx/w80gWbSy5PU
HpmDD5xS0PltBk42sz0dIhUi2UgIhUWUQ444mdcycKOXkQYg/V3L3HMV/oz7gaCC
V71b+MuXMoH8rt6EiiaE+XmTIJEsz4BGov3pVUcyo99VMiRlHPt9Kd0rT0wdQ4pD
9b0OHqmudIwUk5YVDWG7zw+WBIKjyrXvDVaxheycLRy1EoKRs0wfAoosjvcjZXEh
FAeplVOSTXOx4RNmQvFs+bVJByF+xfnLeLUDj5GWLXrvCnGxipu6LtlFBXQhW0lc
/g5PA1MZiwMgHbkNuT6b/bLHQMBrJo0ntx1NlWUQci+TUj/GisHSXxWFVy5XqUeL
Nnsd4HFTmTheRO7gE1uCXh7/JO1ZEB8CPUmQ1dOD/BKvQBRHdMcOVQDkzP4+E4FK
pd/NSbClyp2Knf7BnUJNa9+lddwwEe1fRHmygMT9q+8Xp6BvkFPmLX0n1v2zXo4D
pbHbpqGK5fZdTQMZOwDKPGG93clYZZh/rxKE5J73KNkf/at9DoDWD5aKoRtHKLIq
eRajY4PO+wMxOY8Vq0fQ7vpCr6MNBsml6Oq4Mk4yiOERAU0lqYqx6MLBqd6oasDP
MICTfa8f941UtM29JjJyvE29nMSw4i88xNlF9wctHvgSlB1gYBNvLsrPuz3ppGH4
xniIwOIRtUx2tbAGNu3ovGnOxQxgKiP9c25sW346oU9AsFO4qnRO4tGRuUWAt090
fsGfQetxCXrqonaEgJG8wKA1aJZB9UOIDMhkK0epK1zUb5AWvcGIE7AK040C+6fD
A8ovDzLpl3ldFzeaGAFt8xTR/orAXNuybsvamm5KQBgpvsaZHCAapdDQGlE60TbA
MKONFbLh9zA3vwJ/qJ05L4oc3eCarJfpYAwT+fc2THn7e1iczdUppb1I2394HvvC
uvUgQCLZONif5/QvRGj6tkB1i4UHnwzeu9w4uW1cxeA9Q3D3Sxdrt7m9C7zsKMSt
SbEBJQUWMtiSg3e0GIqXqM1neEpvnuEGpeVBow7fvGPkP4+8kG4HMR1KIQIdUVhX
kPCXJTsoDbk6tVyONkjYlAi5m4xVhscLLerdRiKV/lNCEzBZ2nTSRM1n8K7HtUIf
RBdU+UHGV0epyHHFqZfhv+A5MGUf8OUsV6vnB8maSaRkaghya2SLmK9IfKeS+X9g
DIid3JvujqivHF/icAglFDzdba0JaCesCpyPzOODSVM8YDFcJOn0q8Txw5bLlDFd
ixtqNuTr2yicEIkX2bfNGOF+TZTNU+gg9HxWkWgcxIb1/4ED+3hmSO01YdaU0TqM
VbzkYnXuvC9yzrCLJgVHwRPJAAhZD/lxP3Jnz2L3LEPPT5QMYZsp3ZOzmlsEvdms
i3kMK+qSnPg8cBCN3p37NuPPYzyBng4nxgPShUzsjPmRUOOPdY6WuEljfoP0BsfV
IODkmhXWK5vf7LlWW5MwcHQm5P323WG/Ha1SLGCHQzOMsWLe/HwhgDVhdL4uu5nb
FS9fJTGhCx9pq7QiMs/6liKXtI4pCnEDmuIm6bQPVSXacQzx136OzXImoHNoLTwS
LKNcBv2M87ygaGljS5VU2Jc1q3G3Mo7rM5NMYniY7Dp8sekhxuwG1udNNIik6I/R
4B76F5/mdUuiz3TIcnTknE5xgn5FfDZZx5bJ4icMm0tDGjb4984jNLKpYNywESUz
/Y06iepxWLInux8Fs1gb9+hsa/IWYMkgcynMkZRPqd8R9NRfu+Sb9cOd1m9olewH
K/4gta9FhO2/DVvXZ8KNvCg99N/Iluf37sXtFaDOYRqes3ejJtoMjWZuDmcJyzTq
MuaUhSmlbMCxMsY+zCxvwH21nDBmmLR9OqSiwipGj7KvH3WgKRkqKRiLj/4YsO2b
/0JB6y+4MMDrCzJTHKuYiEPS2TIucJrBVMagt4Oz9o+Jx/uV/mAdiZQ3zpx2tQl7
u6+g3PGj+0GuaWnEQEa0a/6kNr3i3qYU9FRFcg57HYfzCrh2mfnWyI0+/s6EDZ25
jDLHfPzc6AbQRSF1TEi5A2DnqN9DRnj+X9+PXL4VBMZ1HHKGCI2/M/PTzoN+JRxR
3q0aAtt00QYzMIoqD6J49L1cAhnjrwEqamG1fx604naZ5OgW/YsqcD87zzI6lC9d
7Badzd7+y9eLtA9QwN4BScf4i5u48AtwmpZBOg7pmf0Ut+phHEOJ7kzv5ZLbPSEE
P2/HGJkxHr8+yh3q4tzRZib7mNwJSrLYB8rjdgPNqHiRsKjPAs6NnU2V+5YLpL+f
y+h3rq3duRJ2Yc2EnIwqVczviC003Kj7sfpQrAtDdacWkwpYPs3zaIxpW/ZhWSVb
OUSzaeyfxdtoGBNWx9MwuHYNttSwo9liFhEph8xpaHKHvXnxaoiaX6Gy2ToVVK+z
3Gt+IceFBsC9oFoDuTt+qtmFFFMdCWoiKV0oVT3QwkyKv/m4TqJzp0FyV0yBedje
sqrwZMIaV8bR3ElkvIzn9/DC6Ay21M7KgGq4Yq8G2dvL/mS6hVJaF0oHJ2Py2t57
SC6FMptNs71uKAe0yEmzJJf6NEYZY0RgYvTmHG/b755hIQ3YJzh0KWT0UldkLdVS
yGrBFzpjRL51wNnNbLYLvMbOHQMosIVX1+EABrwKhOeQj7UGkefoZNUP7k8lBrwV
xEXCjnYlIPcNOtO3wC8NWKsHvCOO2Xwh2zYbCFPc7Ysfk6xStTOGc8zDiJazluxr
93ieim+p7951B9VgOf7X3xyEAFBPM/F/UHLvUznU8PM4JvmOibtGzPy2B9JCIdvh
b2KfEmOYKQNYgTUoLiaB5+NO/xyI1b/NXSBMHYRS+xtYU7443m3gqmlANShzR4io
ejqDwpJPADuQkViDo9PSQNVrY1avNyqT73Rz6dduUdD5nNRcZDeE2HG9K2lbD6t0
BDicL+QxYS7D0jNk+p7HAQnudZwB4ODbh5a5XWppgNItP5yc/mgdDMgt3HfzMNtk
VeV0i57TDUm6PkO5BRjU/KFHdAnPm5KWsy7ATsWjSRkYgx7xGlAaTTtHeKvt9SXp
Q1py+bYnl4ea0wFSQozWdcR4CcI/j6mhGiiT/V/1/MfoGzEwNJahZWUU7xbdAEEd
IYl9NIZyWO3eHzQ9k7eQRgamaKjddmYlDgGzqoQQ4TK1gIECgNYErFtZsawRPgRS
RiAgA+Odik2NPaKpotmctcPXWSBHgK2GGArFwSorYjlcD8v6/qW/LXs2gjBtkI75
kLNuDZPuVbE1HGKVis4lPSG8bTuimGr/va1p870kQltO1ErI9n9tJswpAtDvscSP
DpeYKOl+ylqJTfrNSEYQp/U5UGed5Jgd0sE5Xt921UMNOfmQcq0F9aP6snd7Nji9
umUHKLZh3S/qqalX5Lar0yQlJ3vhR/08i+QC9C+xDIJ+KOY2+WYstbZ2HZwpVI4u
RyyUVXDCLbDdKzNd7NOng8QWftfjaNeOmwVubf6kGMrnmB+dBb7IvU/wHjxs0CoN
OnFxC13Cu45TmlG62iaYJI4FiGyXVvhb8RStPYaaKGNz+5ON7Mkkr4RZ26ps6h1v
UGn7rgsi4emyi2sI5isiZuL1VInvB38B/WWJsevd/wuyNF2y8bpZA766BywJH10R
YMLNOP5j5cUioJG/HZ348BrNeFkYNLYZuaGhpbHYWWJlrTY2Y6W4ns6kWQAgR3RN
k3lJSOcHUeYdWytCLOpxkdwC8jUqJhJG/gNxG5mDS3EXtOqdtTMdrmCsFZngE9rt
vOlaHlNQqhLaK/YvUVxXHY8w5TR3+xqGMw4bx3RxEJJPlFIe2lEtonQwwvKcim5Z
nhh89W0Wvw5d6BTyoUu9paW8bGMGnKC/X9tMfZKIgcUIt+OgZt9KpxPZCWXOqTOB
LwlgAYXJSSZXoLYs5vM/kx+cujpXO+My9qHeznCEBCJkrihsspXm7V6qPdI1PCLI
lX+HuwLj/nE0SwuGcdhD7O++4YCKKFFyaEpHwA4sz42OkR1GM+RhxdvdGxDnr+08
QhPBDWoe11lTanV5c4hy7Pz15k02uSccS5sratr/sTrEQYKvLmJGhV1aRMRD8vWd
4CdkRwh783H28tQRdz1OjreqF+pv2NLyS/cfg2tp6gwntzehxRTxdYAXHZq3pQbM
p+D68zDbKjdIBHdPMUdZoYZP7ooRNHFZzj4PRcX+YPlR8rs/GXIvbb0amzG+PcuJ
J/QZQgzw+w4AWwlMOvk/xd3T5u5OUTkyC+6v3P9mS71jcY9zF4aMlfQ3TERBkf4x
JXXoK1/74ZpMWGkA4wMRZWSF30n7qXG4a+evgP8ImUE6pkfXM8TIMbxHmaprjJm6
lnRhHFO9O3D4ePylWZp+gI2HTTrEGz5UI9AQh+cuVIkFwAewE3TkQCKwf7LbusmW
apR1ICjePyP+frIKkY20pfBqpDvnwYGAs6JWtiOZ9WzYlP6CuG1dJO/faCxdAzIw
fhezb156v6IwCHdXEVKWo1Cgh31FYNHO5IbpNh2l5/DOFOWw+tDK0nhbhnb+17Eg
GwJBTlLvQvN7KDO09R291HTRnXsVGcJW0xTt44Lg98fpdpVbFQu6wg8JfogybOS7
80Le6NuIpNfBgt8fMhfQ2485ndgUAplcH8sgvtFkC0CBT2l+kYsfJk2JA1w9gfeO
Jtm2augGTbBMZOG7PRMioca8GJyRPAZ5T29N/8BECpGxdYu0z2Uj5xzYpAPHfGI4
YGEeexKvzdtMtFDrwPuMbnMdY1jXO+Y1/oAi/jYDqbGOJ/5omYlf3bJuMoyvLk79
zTCL5Yx8wHh+6kbZ02edETfSJOfISFLqu5UIA/gm0eIAIxM/yOcgzJF3GWhPQyAf
CwrWCc6sHDZitJ47xRwhzKPb8q8X0mrpAUO+p6XiXCK3/NiPMS2uUv5aGGuH39D0
xfSbXEJT6nWqzwsjTjEXy/Se/9bhNz4prltDPLsMZYMXKs1LmUnCjEfdvODBTSR3
46VUexrd5HOh4lKlW6x8OBEVKRVpD8rn9cyAMr5eBWMD4aWH5HXeNQojWdVFNfCn
VrVXxxlyONtcCDXDPza1kedVgWD1PlPgGdunaOXko3TR2Pyat/Maa+oz8h/g7bNr
w8W8e2GToKZawbz+ustMVvYvRBP4aWyIG0vMNESSj+t4U3S/9drorjcSUGErhNls
xLnaxsw92lcnRYAEDjQ/Kx9v+gvwKRd8mmRMiFZkr3o+i0XlPAEcK0khXm0kBx6r
fUtY38+B57g1NCyLXaJ5M6cVTiMXssjNkhKpfu1Tqi1Rh179EvX8rDo9MUPnGw9C
M+N3DBLgzv8aKe2Glq8qFaARcHiMLV7kOBfTll9jvFIRT9gi1OtNH03woRD1DPoA
eIQJTR0WL8yOVZg0d+pal8uPJXV/6xPCUsPtk2pFZ2PBJfz6MwOpz24uIJqYzubn
08RqLFgAFeg96MRmuUfU4hWa6wK2Yertqm3c9xoLfok6nR1krImzlgm49KGZdw7L
u4vXfC26L138JcrtMpSG6a3dZs9Ol/qaaibxVSJf9nXawweeijXC85DkANU0mseZ
nWo7bTPfqsryxoQREf2xJtxrTFJ2fcT/+w7LRkAExi8JCeOuDvnFitqW+1In4i2/
IDkg63xR5buVzk4/F2FUeus3D0dRc7iuqrBwTm4bUjoeigVrTFSQVl5c1jYyc6ol
8ONuyJaalrLgD/9a6P0ZkDL+QkWxqBBrxAXBbFqZKzlI7qOdj0874pFv5J+DAzeY
9FhKFn9SdJrFBC5//STKKXmAUBa2+Sm8uxU5/Z1dLHlKbqNypqRCWPUXHUqqIQlx
1z7eUNWiQjYPpxv1Iw7NWtkNkeY/r6oMi+74bfAvT3UgqpLpuafURKayRVFQ5s36
IwUGrMyjCcWYBVKTrGEhCkpHHTZi2TDzPeyTwaXhiB/p3x/q8QxGyDa1UQVJHoqu
TW22c6llNpI8P8/IqH9uAWKHBGhhSyWEf8vwm8Ke7Qm9rFTgDgEGNYP37VDUTje8
mJLAYa7e1EnQtWRHMB1RyDhIm8WDVIfkhffuMxhqar4DWFntmOyPhl3fyLKGDs9U
C/3RRYG+w2/Zl+SApr5T0wV3cLRnTLA8o/1+R9HsBqUVhZikiCDmAlw+MJVtYohb
AiqbYDQmwu3JQCyxzUvQzSKwgLgoE+96jeneW4Vtma2uoxem1pAetm/1MlFSyqfq
pkAjqEQP0ii/JYXCNS2n7Oz+rP0qWH+omJ+XiKv0ImlK0D9FCy9Z9cebUHScqH/d
Yoj+YyBolxa1/AKtRTsKBsMULzv5+FTxlqQZGul08QmXTflCGsguxQLA14wgTJ65
HVWpg7lx2jh6C0+a067LNEkvpEqO3uMgAMlYXQlh/OTWRCgDexAx3rsVMJv2Y5Sh
PTTSPG5T08dIb47zVp52kTHpLibWk9HmUrVqYaMUDpmwMN8NduTHTxWcvshtJggB
c1echVWhGDgT6lUUbrYTP0zXhShRUFZSHMQVq9mpWB7MoN0Of187dCUC8YUeCFsx
4pynyw/qejOCQAdPt2Lc3THGV6PuFDdPKXjwlXbKeScphsESix0UUyck2M6EEoCT
voE9bNrSOeffZml2BBOyz3rO5YvRX0h6Pig/Wo+zrmPrf7pNanDsIoEinHiaotSh
lqkZeUCdCmChjTHIQl16nsCaBS/58FBSrGfhwggEhWlYE1pvqD/wngiKI3lIczIM
VzJAXHlqrbGzzNOT3lyuO6V/rd3ngVjtxu7eYBM0+r8ae26hJcq8gmJLmMoVs+4M
OgPuw+mtwZz8z6HLy0eUJ2wakL3TPHvS/JyVQj1YzKRIdN025IBoXk3mPuvVZawV
0v3VQGMNtnDyOKSpJnx00CqXIBCf9D9Si8KDuvx2p6uS77vKnLp2NEQHi2j4o7zh
OVlLUoCVTt9gocVWyNtm7BvITz71tWQ+4tHNU6WGWOWIe3VYViaVDfr/kJvL1B5M
98z5coNYNXKWJuq4RKHH9Siy9C5ajWXbqM5/4nKJw4KsD396YoZdtxsMHb+B6TLB
Aj8y+ayjMZuY3EwFXiesBiBVZquuLhgTTMXpFT28bV4oaHCPkTlY5bpAWHxcLXDR
bo5/yOJCa8lcC/Fcly2cgados5Uy7yLu0kqC03s3VLlstBq1Mua4YjLCz4zVK4LV
g1iM6lGGEeakXHtBXRhU0lz83G11srzwKE7Y40th+FoGy0GegBM+ual36N0pt3K7
65li4qM769heZRNJ8SAYf9/mCUJEhwfXx2FBhcwgTNxgFspyoS0gCmuwZYv693W1
EjFfaN3fapij/xuegs6LoRKACTt2HNJ/dnAkY0Wz+sgnF5ZV23MlZ72fKWB4/+/t
egtqBzFxeCpl6AXbbomqxX+Ie48wbXM5Oaf7ZFVYQRYxrglb5fVJHf9oVsLTuXOF
nZwBAVGFvF8b1z2XnkMGs7GdV8X38JGB/yKQ+OUoPmRs9e91rQUA8dw+x/54g+IA
9gBnYHIpXAg5/EjBu3O6rpKAdSgDMKM7A7wn1+jn3DAdPMLMzLeQvl1VV0N7FbBJ
kSmRPN8ijegTuCkJIYztCXnuIG0/Tw/h74iXeZa7WuJzAIAEXBLDQx4DyOV8c5mT
0gSQFt25DmOgI4bGhE9oUZYXobDUGPEAcHpy5mlUV3u8sHUFC9SaipasOccpAOcm
o/nTN6MxzQ2ZDf3og+xIJf6sOObh+H2JSHQQDMwX7GCSgXg64R4nPLgtIXtc7mBR
4AEEgkZym6MQBlI2G4y1wJiHkBfcomEvSWplc4coBcFjLdVwrcxKtjTTBWYPOkkC
2h5YwyQlK9KUHjUMntllQEl/eoWSr0Ewsm3YW+h9X4sw3dgyk2qxiO07OWw+Msdx
vFDjC/ylt/h3yDlH/1sVztItdHZEca9an4bnSqvult4LGxcghIbqYBCOJ8PFp1Si
NQxtbaH6Ho3Uc4jg0VSR4UvDQhrCvTyJb3rnFTMRLWwpt/2nIavuoEj4wxZDu3hv
m23Pw4v9ywBSWHrtEka4lKh1Gy8K2UY2ioTVA3rAs9XiR8ivwf3BQ70EcRHVJtjO
82VtARtMUCp4IzsdoR1flA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
m01bOq0WfT0aP8xyfCUdSL6bxxoJ5FuOR900bzVEuTizO4/l0VJJT2Em0ymJF4Ez
XJ17RqPjwDMkDBlXfZ7NaQ/UjlFYo1mplzvGhFTFQ7umPpUAtZZ94Cv+YDdbmROj
pkEdkmbp8DoEl78LShuMfBZV2d1ZpkGV5m4UssMgasiY8CvcSOi/+4vrLGDZOF+k
SQsex2YGm7lDGkC7D2Xjd6OX0KbYsUJ4z+lBJMGiiKz2QysPwnGteSsJezNs3kM5
/3hzfEn8QhfYXZo6DOpEimK3tW+uneoC/tg8LqQKWv0KjJ0RHCvoV7IpnVNvwFFR
qHS6/gaP2bCp8wnEwsoe8g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 23728 )
`pragma protect data_block
Sitk0VJE2hhp/tlwDa1GG/oTRR9By9AJALkrwoVMjyGXOWdZB48E+UH0G+y/TVSG
5XfaGRnkUAM8MhJOYOj8rJN6KbGrj4cbbaNwheUPmiVVeh08SDBIehjcwd5JyQFQ
cSAXhMX7WQwzhoLXJz3FoO6tuxPMtyQNxAEioq7eO8qhX/kjfW4Lss45K0Tu5CPw
iXB+yfIN7yggQfM5S1Xuzpk1NALcNec+/SfG+phLDGYmflPwr6SDtIUO/b4SDekV
WzNRKAUwtREwqyx+ogvJFrIzdlo4Ay6ip2xgroBUL9wHJABwP8SFnPC2JVgKzauR
3FW0B5CK2qKDf8tmpkdNIedf2SmyF5nZVHRc6q9EUYBElUFO95zZwFEck+s7D0YS
k8VmbUuvP/tE6+FGL0nlwz2hAUg9lYp8oPDoyozrmHhx4a9050jBH6a7WShfiX5s
+7YhVRlrFdyJV1P8LG4Loe0ngdBHtTk1JnIVa9w6F+Vl6EspyXSbUcJ7iy7OHsyo
QTcV1MfJaPWKth7QFVdkoTriSvYfnHg4/U0d++4aNq6vbBPBrpvAUypkqmZW2mEG
+b1Ym1Mk/ePR2iF9OiBnKLiApmqbL0RKb5buNL4rsVx21WkTdXjEd2SX5wPzL5CN
IXbRimUpk8y8sWFykxUuetrGA5X8M1f1t9kumFLw8xFqNK9Ju2IAzfRBJYYCFDgB
DgD/7VpEH4MMm4ydEdOpyiuKmslCPZy/edi5i/ypvA2v1lNz7VkAaQzZVSkVZ3Ew
ew3b4x+qfIiDvF7y7FPIfZrZtyzKWiJ2OCl0MnjGTJRH/ahd1lRrNfThLCCCptEk
5KtdC111VPgu9+0xf+cbAUEGJndskS2oyEv8gh68uyuS2FgSVoAh8mgtOr05CqOS
mQbLsCsYpXz3RJSPpaAdZJu1kDBVcCLfVsH1dfZkScG67pGi5Xn8g0mFKjt9/I98
5GvglL1i9zOJzUIyh1pvUCihhClz2X5fR+q60Q1zpo0yZbFgSsu4RkHSueeX2K+7
w+pdjYMHEKNt3m7key3XLtwn3NdadvtqVBrDmaj31oGoOGbxwQZlpseie1hcT9Cx
8f34fa43UCv2J1CwGjbkkf+kHVUyCmIhPULxuFCBlorkKqQbtHCr8VPToirMuZHt
H5zc717FRCrJKohAYQpI63bryfpU+x8gc6JrchREE/lnI9D2EQKmaNq8HPxUEHez
SEV1TM0EGa5UCNRcO8pSbD5tXuxRAnuZ2bi81QCUJRXEU7kDExB2Bhfhq0z9xhA9
X6YPgrWFc4mZp3/A8N3MOnKCBEJma7aW6TS2DZHSJCetWwLEnmIdvJGH8ty9rCXI
J9lr8QdP8TqWXJ72EY9cUtQ4AJz34LY4Nj2MDjJEbqHiR6Cp2XjS0L8qaPAWmpPe
gaG9dluidYghUt6wzke8T6k8mdYheIM7soHy+L5m0x19i+ms9REvrUByBO+dLAGd
ZGZWwQ+ZlAxT0sg8UKF9mWkt/LnIIeaHAyya9AyFuay3ZbSOoInHeYsnPKPMNLzE
kpHZgCPNfta4Dfhu+A5YbbpBsAAVbeXu3awkuJ9pzIQW4ilnAmeproKLxCxfONJ8
SQSEChUimXjFcx73NQTrf1B6YU/u1xIjG8nCCMMjmYlVggKJAtaac8+hduax/I4Z
6WH8Jk99kHXW6IIy6DCHeloTxPVnBXqSGCq9Jxgm4dW1knI7/ZigSHBNtXihOBPK
AGQM830XlqJaZ5PSmhqNiSbyMkTFPqt/W3eCHVfr4YzBFrUF8mZ7kcL06V2ChXjt
tkyf1K8xXgY4hkcWec7CQFoXkV/wT7nF3wrFjif9gmh+098uPoszkVFTBzaVZD09
uWF9SZRTZ//kJw2MTpL3foK9Xfn5ujmJbSRzLVOBccUutBdpbFmoJAFYgrWzwZ8Y
SLXlkC5gjZEsF6k0zYTgiXjcn8ZwkKrpKxfjFXCLSm3J6MfoGPHUg/5egJb9ZVds
i/CmcvFix2AtVA5irDk+wjVDL0HMAsDUImI9Yv5mLEn7PEWPxh52mLjdet5qyfeg
XJv9/c9XqkGWwsnh0CPcNLMBeZ97OSkHATIO1k4I48XuFvt97SFqG39Y+gp4qewO
PnwZZgHZc16P7F/cK+DIHxQZpdffYN7Xx68jBRN7+6HsHVMfFpfEeur3QDLB0F/U
TnMC1ZmofSPP54rOQkrzeZDBVCl34QJfpuoPBkZpCuiqtcgODV5xYslofSVnsobQ
R5NqmNpeIHLzCgoTYqQKxVNZ1gmTpBmI5VqMarLvudzBQ9qYD/MhlTLy3adwKIrh
xXNJg20q2rT0tFdr8ivqansb0Ovo4h5mJYvKZPy3hJGii++yzJrFQMiWaE4iuQ6y
WNiT1y3q/2Rv4CUAoFGOGEkg7N+WnZBsygadI6be2ib/bxZi/hMJ10J/TTT4TXPW
0+dElSPs+BCfKItoyunPFOXoM6CvFcWuxKRQ14gVp2lFa9XQVujw0N1CJNPmb1cK
9fiUFXA8iJ52EJU7O0lO63h0hTOnfdLO9d98JoLGfkT1iSnEHzbzSVxfW+XcLq0n
O8DAqXtg6+4jYkftR5CzA8/vpSncbc81ljIZzBPku0Sp4eQKKhD1UEMrWffdJeKO
NGlWDbVdO8fStgzf5rz83/KvxcwK+Wvu0kfyX9xKS+MZsQZ21N07qx9RcF59jUbV
fM9inUtS6gAsBYHWLVO/KZphoPR6ySZ/TlqM3DTf91eqST5nW2HWSV6XijCRuMdv
sSZYisEftEMD1eOhsO9rcXqTr/00MbKH14xTFpgRzJk3QGOIbGYK3mJQQqlm0Ccb
+uzXIFCLt20ILM+kbnncrh5zGwgjjcjRu14YFHrrWRPrT/p8LNJNIGuw/ZdUgNgj
f/3oY93YeJpB7i0dTTYxwCG+hzN95Q/VLlgtvu9KLAGA5RgPX7wBg5siEuuSgni8
RKssjqw95BGK3nHTTsZFqC1K+PVsPjEpXwhrns+yALbonmCSXLRyGhuZ4z0GXmN/
WqI1T4gda+rTDy4AcHQ3oeVGoNgQKBHD5Gc9kT3qrmc8eGsH1EENEHVeHeQxJs6T
/wVSO3sOSNIisdTOsNeFZ0TIy8Utvaf8nk/eQZFhKn6POgvLdxvk8J71FkpZHR+N
7zAm3tkrRzBuPDPmyD7jm0CWKRU1T7bGasbJE+fXRzi3uMDNgFVIHdxskonjvrlx
20UxBSBh2jMPjXEPh0dA3zf2jp0RgB5y29lCZaQWVKfW/8ZT+BW6uvhsH98D15up
hyAMpL6vFSrnLZ+lTWBCpBQD4Wls3mD4PS+NlB1lPtJlYk1Er+iCYRG6cJSMcKDA
pajEPaj6KJbjLt12xEzNKc/fKyWOJfP6euRuvkjaFizE4gQneC9UIVcF0006e9kW
EkrdAJgfWdkhrccFUVZeunyAEsrygxdIVV4AtsPhLIWonHgWvDC8I4nS5mrlJ387
g/7nOnajJYjjlvLRLbEApQ3x1HH55LjcUmlEj3aqK3HDhj2V3AzBeH9NgLIpAV0A
aDSVNaWDgHkzVId57QtmhrzL38I71hShLmHPQm+5dmSwIbOQuhk8h5EBk+9Pni92
dtgPJB4kKDRcb4BsNrnWIDTW6nIvr8iZUufpwAx9rIl40mfC4130kmIwVfXlGANV
vGxVZoffEwdQWNf4KArJrDnEFEDf3tUeX+F+lnjvewTlLpDYtjLoZrZxfOoWwnJ9
jDiWGy+QMhR6+etFF9wo7xedmZ2hKwsI35FVuNLshWsa2y+jn/5UyrL22Bn5YHv1
WjxaUVzmzynoLwBFYQ90vb5R4/UrjO/WvlgvkAn8fp8q5uxiWxSHXxcNSWbZjYiZ
Vv9eKDFmiBArHFGWcuiRwyVp9t2dwQEvGpAEL4UbdHaLKby8dwHabMXVtq/CkgNv
J7URhnTHEW5Le3goPpOb7aRByUPVW3OK9U3aJ3jesc+Hox074zT/nTJzvAmtJPYR
2ouKypnU19yW28LT/S9RnTO5ef5IPDBv3p/rY4Pzk9b3EKm59X+wlwdcRrqZhe0x
/HM4eR7VIYx+Y9N143IdFMDsZeioPNW3udrRQDP1D3Cwc+b1hvraZrmXpORrbzmF
3Z4D0mdFJ4jfCelk9XrgPbdbozCd75zYrKMADk5ybI3c/i6Kqj43srJ2QHzhL9eu
SQS8QyRPFoWPQf+kBKiQlE/SFvhUSwry4qSE9Im2d8QmJdSNHLcnSRVpNW2DehzO
p15rLiPmkkvCimzdkdg3/ibFV2JRxkfOILbHJ+AQyW8spiBIfj4gT7eLzos+tbE1
Eo4w2X80FZxRVEtCqeww4O2nb/skipiyPcZYzx/O8qvK5SXGC/IeC1Rc/gCQiDNk
ni1wNEH2/AtTgYNUJQXc6OeXg8/wMg2UM2LaK45ZV/WVsQD3X6Qbaj0JkEkXAH5D
VBVVGuaAPlpFm1EFKWagx8+K5CX4SeZDctDB5AmS2RX/VjMIBAU+Hpv3hUKMWPdS
i5eA9GnB4D8GnPmfFWxwB9hGNSRWvkmPbRcmJ05MRdiO1qDdkD+1BtF90vAvuJWA
BhFvqqCMahjdAcfdiwNuhYfF5HmB+phnKrxvzAdCtl8YBhB1MdraIA6N9pH2eMzj
2r0pAzlYyc9slg7BdD3K9aoKBBSs4pCct0dtSQRz4IDPfP3x/SgERltyDF6SHcKT
19UqGYWAZBArZo2iB+JO2dLhR/ycNmy7NkZC1rKGIL8kcsBl5NT1Rpqo1dEE7+cW
9J5QSgSWkLFjj8mfA28jwDEgR0fsgAq1QfbCplTX+ufawCMZUx5UJPBtqO/M6sY0
/3xyaOwO/RAPkAcNQ8zmadMTRgAAZmNsOFZSuKxl+NE4N8VJNnA8lwDvOAQfiePP
erLItNsqS521hUZRQjvQ8CXEAg9PSOx2n6MwAY2ons1XU8hdVOJ7G6wqKfUlnyJf
arFQyeeOvsswh1LN5XTQi5VHs6+pfknzbAzzj6nPccHX6POcR/dYd8TWL51YqVCS
yNX0B1xvMXLl9NUzCfMu0bNx7e/QQ1gctoiyu+p+guetV/HPbOKgIM2Y023pB9ku
M6JSsIoALcIzR6AEF6urQ5pld5SYa/aMg4GLdh3JdbBO2YCbsQH0BTbrT+n7z/eH
og7kRi7irSZq3g+Bcb5aBy1IpWlrsTvDeaHNBwR17mcgbSB+jGkCI44wdX1wEn/q
djdqni3NYH4aVQk4hdhOz9fhrC7NRQPE5wHaiJf1eEj86w0d/rc+ItRdMFw0sNEo
sJHQJLj/BV3UoeE99IBAIUAoCs/5FVA2Sa+SAL9YATlnS7opZIGuQ789Ept5RWlM
fH45/LDVzGA2mPnqRRMT3xhiAjTTrr2IxE7UCzHjV1T0QKiP8CZ7yfnYGoi1prDf
RNnS/UULsXIYaIL292bjqrluhPoA4pTN+EGO9Za1k5nBDl694wwfFLQHXxfvEm3m
oI6NQBp5bmtB0rdWLTYfrt1RycGlwbRBmKMjkqZ9pYOT64XnOod91Vw5+ne3k7NN
ILpgnV6fRancJEbrPwad6raNFdEs+toATcH7f33ZlAu14bJAz/oL5dR2DP9kOZKe
WSZRGzq4EF3AZLtluMft9q+5zaABZTBPT8A1q82Uu9vadtnaupNFE55CvsnCNYW9
Ykb8jA1R0uYjaCANqBM1anvOEoi+Psp/orUkw4NNyCd5Mznvwxsz3bcZpF/EPT0q
UoOQ+YjSWyilfRodwAcMjMhW0aB1QnuqZDGBz9+2giHN6aPBbZrujckTkJTesp/W
clvJOBxfptLYZqHt3s7/rR3zC3L+TCo4P7ZiyOZeoyOV3E4D8ZaoBm6bK2mThn1d
jMOo6UApoA3ZZ5XcnTZ4wAt5Bzh7OdTI0sz+sAhxFM0yT/jXsbq6gAyXgbmCsqp0
4dgGJtxPKGPzNPFoOuAfvTZWFpM2fJhL78Uel+YrRm8hacj72t5Rbgr3eBVq0G+u
3K+FVA7pWQ2UbmN0fyobCl0vJG/uHA5PCwdGybLBawbrdtS9E15QKF2h8TU08B8p
AojgmaNMUgkrFkRSIrJpc434v3UI5rvaT2va+4ELIQKrsFNax9MUTboPXcWd5Q7C
tGJluAnUckw0bTtWKbryXT2dKmA+Slk/H6+NcUTvH+fpTdEQ8/xor3XOip+zbdul
jhbWolvsJT5KXD/IYr2ZBG53VL1KAkfAD5NfihkfOlZ+e/2hsecXM2jERJrkT0Fr
NKHUKXhKJRUEia58ylBclpBXlCXEsNSWULn64x3KaY2bcacYLX6q1eyXemiJgfRf
ShiEOnyr1QMi3W5C7ZbYaHWR1htWWVHFoXp3OsP26M5BJeWT72rXKCLEU5QyZN0w
PkAZlnQmpusmUqdHrLfHbT/GK1cUKWiha1SwuTlpDfQcrazrd/9kj+5WsT4ruIOo
d7GjQ04sdRm/ia34laY3P1a8L82eGsem1qqmYDd2eZFN7iD6hsU0YvMZLXRrbPU9
oGw1W0lyVuxtmYtRu2gzwtC2JX3vlVWL/22U+GNDiGmVyJXNnr2FTXrVZViUEcVP
jERlhUu3V7y/aFut91gFi+umojRUcSB41gk+NZgO0dDT3uWULD+Ln1NBRfiRvm5v
cOhyDQYZFGvqnqlmdFwZyDzadmqT47The2l6mp7M3IDeZNdsmkZhgQ3MglYs+DSf
yKBbhuazV4O0sHBhq9SStClJp3k1ONLVHlNgeJjdkCPcCsmkH1koef0WtWBLpoOk
YWysSWgjmmhu/7FMKVL+MPUuvBGK9m/ZSd/HNoLo1PH/qqdKH7JKWEGZ4nffEb5D
gcoxqUzq3rHlnIgLt1sZYbqg/9TG6vXDquD5rT7sgDaJxst1IXMF8BA0Pr919jO0
/O1lOnGNr3uA1q6x026/+CStTuMuzrzYcHhFRjxySOqrVguWaNWxu0JiQg4NYF1W
Huxzz9X910fEljWEyUo+jG4bX4hhb9n8ridQmgK8cBY0N+lQILMoH8SB8ln8c4R5
+0NeBLRbbHedjqbbxnL60CJCN+0/PUNV8E/KKOq+IWtxwhJsI2Iqs5R9yXMlMUGp
kPn2XLMhX6Hc9B+aW07m0/uy+I4CKvh41EKSCldqD1VhWqsRAyN09iPfqhbx8yPJ
lucBKmQGNNIW4tlq4DyfbNMJMdnNCVSoM/G/gXJQGZHc9iZC1GvbMbohDkOdHGEG
UwT4OWewZjCjNevFNBMxvjRIG/Kn4aqb+SqfgM3HgSO/bhNdM9e6sCmeLkMlChS5
iBVrozWeD2GmjLPE6dsqqq2Y2w3Dwq5eW3uqfIrR2lZKIlK4SriclF1Dh7xR86+N
PJXCdDdsdd8WjwxMnhT7Of3/JTRNQVYo6fs8VuEmMn447Mtnr8Hxn1sWxfmbdaDy
ItdOXPlCPwSBwehl5oiP7kVSEKOuJiI6idxi+Zp1E15GGcTyIdoXja+BFLNhpx+8
6q2z+Fw++aNMdsUv1Z+IgIrDVQ0UaTgy5sGf/sMaHj/KggHDu7LjVQw25oi+sFTk
+TOEhmcX7fic2lHWVSq2qS9gzXjn486GF0wtvUerbvTPrhj45za+NXVXpJIawS0p
f2fw7RK2Q1UFwqlwHbDquzdcBhqb313ZO+Xi3+O4rKHuo4ohJaepSgY7W6Z4Se7O
51YNFbJLntsuf6hIJGNWIzFHplbu6d6dJlAeYn//QN30acQjdqqmmsNaZIEZRxNe
VsDzzksPw0qNDZkA9qEQojgpjvNvHLX0DTFkgBvdoVevFmSmwljx/LmQGdd8tYYx
EcdBJUyXRFF3uXVu4VLe67QxnyvNTgoa3Uat0lGLMGDDofEZSJeKwWOLJVt++uiO
sRAqnsnakx1xvzYg3LfF9UPYh5XOtpYzrexk5TObxLpKpAT85Gmyd9lEGz4U9sDH
DGRhbIMLosGQLQ4kdWHXIGW5t5J/0voXmSdRXWlkIfECg530x64cT1oYOY3g0gPJ
bMCHlwsiqfaI5OVWLmJIeW++uTpu7y547ea6kSLu7cmXtazTaVfkDWHQF7PAOWmu
n+TXqkZPXackEdxDlaoEoCG1De3yHGtOJl97a97Qrj57Hu+WEJlUxkWhALnCo0Tz
fTxQeDxnyKp1kJszRjRnCg2x1oOULDKal5bJpMY8iMwnMFG1/EBw0SH00RmS64Oq
bSITyDBnq6X+Q697Mco3HXuJ5ybUqEr8MWOEFK0v/U+0078f3jiley34XH6qJH0+
8ubxMVWu7TKPdZrPd/YUjvS5AAJIRcxXmTgIA+OlRsUJxcMdDiWYPVhWPLFLW5Tq
Gk5RNrojlxJkGMfxdsKIkxwCedpg2t1/38itdBfQk2fLNOvts32aUCLmPubVhscU
53q4Ru2MHxV/a9Z1YfkxJrhZ7mU22r52ReYiatSEd5SZCRQiVUrL0GPUZmyCvTl4
8WV5yZLXOMjf9Y/DhEN0PYWVmfpbeiyzBF1RrNrYJqcReJc/9DT5Zt+AOWHyxZJJ
1zOqGc4NY0p0NYnHNAzriDqm45rvESwCg15wgptk3iyM/lLSVVJZPwF11L8g3FPC
8oY6ez2nS0yIRmrPIU+9DRc/hzOIxKjdW4SiRo2c7SoLXeDU7VXjmKVmQpOvB9oa
Rxv+lkN1Rve/SXbWLkAnPYBx5QUC6aRJtlZ3kop8TwIJGQMA+URr84w0VgLRSCxN
BNBCCUD/nUQ7OtEav1j7tS88RO6prqJCnxqg+93fzJQV1eS6CksOSEAmbCRQ1J4M
FdJgsZs2f/Ngn9TqA1sAlS3Dw1FCi4gK1jt5kOUPzGyicWdoCypBOolIg9zamB8l
9B2FNU8INFFlnsXVJ2ynZiokOXd7gA9t1V5K6wasgqkMRgquCr57ZREg/p/bSXSU
jfzv2BIr47KGMe20S+BMQHf4j2gm8uqFeF4drY06Ibw2eTCUi3drp9KQjdSrUNAU
LFLcn4YrwEanUuvBk6+cwM+WOWDOTWICFfFp6uTQPZhPTsZ/FMuNeJ93P0rFfjgW
357dS6GevE9uq3Fv0Wn6AzFLM14ZKvUrzBnlSG/vzeErYSKgACo2RxX+eCVAM5u1
KKsVeZoB1enOpqdbL77KEB9E/ujK8RhZHy/JcHatLIofVXhyZRwMFa3f+T2LuKch
CbMngeoOGH21M9oviQrfwl6/HUiyar90zNGrqPepPkgyV2VQQfSc664WFPeWSAxe
Aw2ipXXC79cAnU5XnHmtGulDurkGOX1BjZ7NdW4Cs4b8PUihnq1A7EuxGIDASrsH
xco52FweqE++E9DgpJ50NfxZtsCzjzLs83DbsFrI2AZiCOi0K12OI39mvAYX5ql2
9LV/YKICkmPcPk/sKrjdywEPX3ETG2n3mUfy+/1Blhdpf5F1qyozWf4J9d+S7qZR
8dPVWfZ4euigZNjKyKKtjs1/kIIW4iz8mWn0bh5CI7jk6K+bwcOiaqwZlEyvxDmh
18eUPEdpnLBtqu8zg1p7tBmLRgiN7kJkfee+MRL8jfpkJRQSYNMVD8V5iAIrC05s
CRgwOxsw4PWpQkkK0qD/l02Fho/6EGzk911U63UbI+f8mu57j5fOj7aXwX1NOysc
tsaFkPc9BFwOTRf/6/RBDlDqV5zCoHT5UoOGkLqwgxk3JazbLKEWIJwFOBrkrA0X
y0WMqi2rYBomg7nHru3Bo6qNIqkF1+pxyxhVRg0gC8yGbdQl39SOK65U0XbSWQz/
HVlT76kab5Fo5htrBXUsXFxIF/ew+Lk/Xrmu4je3XKehfHMOPt40vrl0eLiKtLvf
qO96+7KJ1X7bLx0ak88cobhDMrxNWU9OpjRdUd6nDp992lueCIiqvDe453UaOi/F
2ThEMtSn6iEEfgprBCMQo1+8HPoQ5QNO0SQLHj5dSyQhig9a7ReOECj6AD1G9yAX
lKhUEGDp8Mj+vifXXoubuyUNlE2IWi0B9Gig+9mmKtqxMANfVQhFDntVQvlR1wni
dctdpZMc+dcRwxceFbXVumLjZO2sUnsIRREMvQ32Hm8tqP9vca9KDMZuKRNhUmvG
vq1bbXMgQIIHalwYgYbNHS2cJYqwd2HrVetpbvTTcFyNfMdxc/JAjt7G1spPovnr
2ZPJv9G/3eh172n88R+23r5R99U74BwwDLfFe1Qqfv6UwIC/JVBkwDq2Sxg9H9wM
MLeSj8G4BIhIFdL4FbdPqz72D/spgyeBGWpGWzNI2g+bGCobWJ1fHnyr/BuWaDyt
uITCEdq0CRagy2xAt1Lh2CTSqeRbEYvrvDGkskIE1D952YMZi6izdxXPcnXpo/Yf
pdTj25hFUazr9Jvh80plaRBc5ngxtVywi0cre9ZtaCvhQJ+7E108YlTwX8ZVwxFG
jVF/7fK+tZIDlyf1AvlrhU9zzLs+6lIxoqGMO+DUXPwBR2KEejzqqOuRi32nnIlE
vqsrzIPLPPQk/3vYrefvqdR35qVgxbuyj0ryMJ0hnWbhRPMdy9YRgvGKs8YvzKhv
+cWYnmAJW01g/ATOQldkZCfZexbGMdzh2ylLQ3uuPMQapuNrRPAHkbJgWErOdMyj
5vrqGzXl/QIlsFeTBrcrOCYb1XaS1rYww2CI1umE4ZVJAtR7O5GczbXCvWnYUH+p
Y6B5W1woI1NaR0aEDqrw860VaeyXxNbuO90dsoZOLcmBnz3RCpbZweIbqRzOUS3o
c+JarqKEqLaJI8QXnEyR9LckwqMDY1/idVHo6+KC6Nx6NqgtSrkASEFKqqrk7fx/
Jcb+oBYXUSHxg+tKSM/k5apUuoO3DEkf3Z6d2eaRusvmk2794DJh7mS91aB/TQOD
mjHQjDMaULacjWbg50lJpDgvZvN5aMFShsmZN+OI624F2kJP84ezdPwBeCEjo5k+
scZjChxBT0BjorB4mSyUSqMurIJKgABRqJ2EiiS6GQX+4rz4gCar8ZBCLzlIpN/f
2cLzSmntU4JTyoYS2XxX5n44B++UjDlz0XcqcsUshGIQ3440d6C/l0I2QmD4h037
SN2nrEBnqRySGh5M5Y/fo0vDoejsKADv1PehAaPXBCx0u44IERtOqypvlxGvUM8W
tT7ym6O7KuSx5awjpFgVpXDgE5QOm4Wautvs4KLw2frtO4e/G09kXX8zuF+22LCC
z8PO1KScc5nO1aHJ0GncXl2EfNdvqCJoPosHXnC5Kh1i/dvcsJtVBByWGN6AjmEl
W3oyMDj7n6J2Ak/Gtf10H8wXKkwWVLKTVUwQOBZaKmK1gqFil940Fq+4H6kydqi0
w5NZ57dRcyXrvI46CpLArJ/Iw7HBumUYSJM8P9xZzG7CWmFwtE/p5Kgbcj174bzi
ONKNRz/4P+NjihxscvDlhMz/xPuuXEGyfaqzmzIuztuFeBXQw/EdKEAFbkH8THD+
fcwvQbH0eDCdmeHff7HE31XKSRh673lhJovyT4YnQ1vhDpADg+GiMgefsmO35ULz
8Uf3ti4ZO04pcqEtsvXZCvalhiZyLYM6B3d9w0t+8T6YBnpE2gkS0z9tLUyn1i6p
EtjwBtxhCTGmiAKaYGHnEV5BNXeCpcOLGVwoKjV9E9dKSrXIESr/jvb8P2Qgx+8a
BerRWK2pvOjVQ3YcViko/yx/LNCAF5wbVKxf6JU5BRW4ei+vKDRd+0rdGZWlGE0U
X+3RCQYyuwRHI05HTeyNKREXIGnTceRZdv7M3op02INrwvJyJ4xttxTw+Op88CMW
pdCIROBVYe6P2BV7EthQgvglwyA3gNnI9NLSh6Egpbw+YeCp/MnX6mFXod0YuW/m
S674FFtczHoaFWpKvbeGZaw8nuC1dqyjUBmZK+IjqqJDVjm9eM/t+QS5ybqXOHL8
3Eq8XrqPG9yldKgYS1ipM93roqAt33xfyiyndVHB4hL1nlhTRIvfr0bTKNTYpB7e
jLM7/r0WpNWhrPnTKrvg91bBALXI87KKCPQY8/U+EoT3Cmf5aSxb3UwW6GnQJGHX
XFYNQBA7pX7KimTUqEUa88EgwzFcu2afpEVeG3aS10r/3hhwG5J5EDFasTHn6N2j
+k7jmqCt9m8AP8S6qDcrYaEkA41amJoJWsCZPqItIIGEGDG3bZnApPfPjUlkqviG
Fx+Z4qT4Rna1yCHt3djlNoZB4/1+6/hlTilMN0phKeq8hOehuXy98X5MkyV7BgMK
AqJGBosayOl+OqqQlmmVPiGZ8UbwGlZ6d6J7JVmWWSDQcElp6kJ+IRzlGpTygUWJ
UAL2hSNcCuY3pq3G11Vg/R1kGetqOao0e+HlBzvD7JNdmrLP4b6ysI7p/ljh80lh
dAOavujymttt7emCaikwERsP1eM3lmcX1EzpFkrnYuiYd8owpEct9PpbJdNv24ub
iBUsaA1eYxYE0Qj9fD6bD6KaLWgTPkFywpYhHfUUnRxmG/wJO1NW3bEDJgQ+LKgR
CSxHZgu1HBfaFpnRcsxhuxrAWcn8eSYWkb3LrlOuFGgtLnEMFwmTddh8fgdthaua
Sf/dZ4DI7Hyi3vGicpKGplRKF3l4ZyET8cViMfI+zZqd1q6hsxAWr/rX1yThovoN
sZcrGDSvAGq/KV6pU6fN9IrWTwNETqdp5z57YQiYwkeWStgoPw11IMZ6+pJei7Sj
Pyy5ivk5DIp20SV48vjI9z89RaMIegR4E0/57/ee7rmoCK2xMME6X7TH0SesCFIF
lhCCGB5HgoSONUXLnYSC8cswY+wJzb8cwpK/DTkA1MgaAqsyH9NRYNJ1Z5rd879E
DpUgIKCOOg1h3t7hDnaFc1Z5NHMwhA0T75o+ggyraeLOwpG4v9akRr58+queEHj7
SzUCBRIR351vl+B9cIq5Rosj+q/784Njt6nB2zsmkuIb3VOWoBWMSCmqvzSvumsd
9jGLdxQR6rQuHTjamAgXrlbLthccf60BW5kNSuZkdmbHPRj1DtpSi17It0xpzhuJ
WvOPH7IOJMAv5Yleqp8l6WVqkortcvZEs82BDKgAsO9fDYayx7fH0hnohoLns2WS
32wW9TcmSTP5h8l1pqxe8tCc4FKiszEp88q95ybI1Oq8gGwwLgqGmthoG8sRc5mv
Bx1raSR/mDmT96zjkryBuj5ksvYKXBhgtjGR3UXf8tLGaY0V794XnQ/pcTleaMO2
zlejgcyktE7boEfeCmTrZsqKd9Jfa2xGTSvvQlzJZf2gOz76T2mLdCPq42ymBzh1
KaNqvbMHRoDRbptZbVz97teZjOhQMcUqF/41l0FCLDZhSSWZ+CNRZNsPEHvUape9
gjsOo7bepPWQ5dNqSB8NDvQ78CpU6Vehqn3lcXaxCOm+s02RP8X8g793hZJ6ILsm
Aojwam5+OBxvt9pjwQXKMGTjZ0ZXCU6bTDIMidGW3h3B5LzF59bhlMLtY6TIcvBo
EKM2eGLKLxQHsZpV2oEecMZJsgwsEn8BPf0cXq778duySJZWyQKcuxEkg06jWdqL
CC8oxUaF6zMnDb1QeWl3geBKZ3snkCZTxs+Zs23QKFoR89oZ6zNhIsIgbT+9PMvB
qNZ58o2orhdrICWuaUB7HQqGlvArnU2Ofb20IQki+D+79Sx6GWHnAljkXxwtk4Rh
joOUluPdPZoAwFL3L8iUNMWdCgOYOKK0Mae1J0uKwMa4jKVKyBdGBDqm4kXE57dR
tm/dZwgRxOR8/2vSHduFb+JDqVoBNX/6Su4DjSTcdxuwWEwONu5QtF4OUgT+XMNP
AwyyGjiailtRXIo9eM5dIoLRtL6nEuDbwkkUDf5EIK5TGziTS8KwuA6jOGQ96tvf
kUDU13tfRYRfxIMa4CoArZe0pspAsHxZRR/zjEexrwC508WAiLKN5qim7EQ20LNw
WIopXyraELlUMBa2+qtA3NbOkYHpHm5sa/HOVFWfO9PHf49MYgL+3m59Nu4v0boe
tZuA6gp47dhXCgIyYpdGX75qCzqCusa8pPf7Pd2vIrplpOZf9o8Gsg+Y01UB4wr2
1Sty7oAiYhZ6WdDBPYutPIaNq9FOD5O7vhSaTZ0jcI4lKBJKXmX72rNx2Ch0o5OJ
lUGm679idgAWAl/kWzqf7N79cStKSrIypzli6zpoowFOSbR48JzNrg9o36pGpvSY
wUM+GYsuZtpP4tyjJpPogWzmifYZmMkmwLPqN39TGt9/madm64rm/VBwFSxwZnMk
f2vrFIFl69ISXVGVJ4zudu9l+E29NbgsbwK4SRDuYbXlja6ZZGMI4gLPMNtpQFqL
r2DLOKp/CrilWhS8wE6H5hONLdNodHOgrZiayWPO/x1lWnEi+HH8iLgGJ3f/OQZr
qeXYPLAyxAj8RVpSHdWbQ7duTNwpZdu5BNSFyzt63hluAtIJ+viydPvoMHWQbtyF
vJjxyN1Bv9OvvfZa98Z3hUTMk83YrjagYtWll3kexMFYHBxmz1Bp0cQJKixkKoPa
XZz0j5Lo2YZOH7HucP/HfKhEJ/B/242+wR9nyoN0bJeOL1l07BOMf7r46FGBzaXm
suTHZB7qCKIHjlVNLN+z5pTfr+IWkKcN4VThnefyAHPjg8+2AD05E+WjNYZoS1qn
xkSjvKBM7fI3lsBnjNG0WrVEieMkPfZsNpPl/eUaP5EHHgruf5bAI7GaM/oRhW/s
JmX3ZxZizaKljRkZuNDgAun7JEzlWWqpLwuq7vbdFZKWRyfwo9tD9/395UimF69n
hCghH5MfwvreEA1AnkZUW5sTnW4avl9p5G/KjLs/OIVl7HVFJgcUXYI2DYTXJ4G9
mu6ISmTtYClj3xfExMqBHJaa5Sp3/Y6ShI8udACbtsM8qVpdUZE2C/sIsEcRTuSo
z7QNepiYc25drwuc/sQEoSiNryHr6Obln8k9Rlm+M/tUSOM1bmumWaInbn5Y3Gqk
qbqoJdYycu3azYnycKtgxab7qjsomF5auWnwRTHxYX65rYcUQ5k5fXmBdOg4I20I
mTJB1oSoXLrkWeg5cUU/31DSajYJ15qslpg4FAJRQmYUl2KlWIvrFagP/meNL3gR
nTtsA55AtsT7MrH/ZM9X32TqQO4jkDC3xdWrFX1MRDotjpjp2E2kCqn0cHRoymXj
+pGveLPcvr9DXSsLo+8/to3d16AYzuEWJdKJ6AKYiu4ENoIu/8EXSJq+H9zvCxIq
X2JJrpN6dmfHwZdJEfF30nJg4FpzjGaY44+5CfCIXexeROUOJZl4GWi7h+nhXHB8
nISFyqzWYRD3/yw8LrOXsspnD/NCrC4RMyyXMl8CuDuoA2a5hYcHLWeqp0Wai0kG
8KcQ/uqBTzyE9JdEXVmKKs8KsS+POdkMWQnGEa7OvwUj8qybprRahmc8FVvKS5y3
FQMCqfKrO3PFsPqqrRk4ZjrbR81QKX4gcs7YKIXtfYc0tEoHnyxV2SuEM9J7MKdo
ns/R65Ad9QMRT4jxZlIs+0DF1Wqb47jFWI6J5UB8kIKnXV5436WE1BDwNe0HCdLv
psCO57pqiXiYN059qHBuCS5WBgl/Jp9lZENTU8m4DiDcY8k7q7W7eN0KAVi3rvu1
FJ5T0Zb56kf+PlUVeHgnMqrJERi8PczvhjDIDHqZJNEe/vhEYdw7SecLNCs0PP1T
vTUs01vB6LdBLlRDwDhxKcB1ZeRSOHeSwUS37TO99gUtfci89+vaKVm46bAYXTVp
Fpy0nP9SCJBVrAl40NE/NJo5Jl4KMG6YTPO/GyLSHiZuPjfKxRj+4juTnPQ/6am4
QhG9vZHMYdnY5gFmPm+Ow3dBAWqT5mfD0sN0+AqihOOEsdBH8JNCgW3lZnhP5vbt
M74/i1SA7UmkzPWLttoKRx4Sc2HQ07jt6/Qwv7YbmGJ7RvwXJZBmLSWAZUQsO3Aw
Ty3DlFyIpebdjxnOR2VpIcM0CbvHGd98JMl3KTxzTm1Rmdg0Vl+csRtS8ySHfJz8
H1E+yiIQiEY2O/tuXp5BpFMvIOxXD97nULIeudBdFGAT+cN1VBj1/ftp8eGRZ15W
aX1mBFDJ/R3PowMhnL3dIqHWkUvQZqy+SEkLRGPQUCenpwlJixhRAU7tgupaOygy
fpoXnaotxxCm93Nf1Uf8TLGSxXt+t780khHHM4/YlmzLtIn+z5pDVPaTkUwnKkAc
w1ylA4oSUpJamzj7TyKRI2wo7yfdYDF1260Ix1/48GYfV8a5NO0GwjpWZpDxsjFN
MAODaZxR98MlNR3Hef3tr1WWq5IJGxZwOnyXRDW0wCqzxDmM8iwvTayrHSV1p9ca
WIxedGh3CfVnJbFdowscIvDtUZXz7fgxF+41iZEe51ZndSDtqVW9BbBDZGHO+sUl
BRLMmjGHnOaK4AleiiB4zTjpYv4zwkrAPKhrXODddn3zNSrG1YaPsjSp5rmipkf+
GYQBYJHkY7uIyiIa/fDD17vA9zdhxglAFpFWCRko9PP7xGFzcQHQHdw6SAssqDmz
oAHYOLsejgcZ0TZtzEZ7ojkwlArBzkl9lyYVOa9SZKMg5bQdlSea+FeoNNsf2bph
Jx9zGimCyJYhHIcrIeQv4RYLyUjlG2MZlTQfZb1HxcF1KqssUDtLJdYiaCO/SIVC
ruhhkcJIN+XOXrf9UT+Afs3XF0z6u3PAAjieQTDuEnU7vcSkVQk6LvwfsNOPbi3O
anpRdLsA8or51+QGKZPUheOBEkAE8BEJlE9xa/UzZ1ow1GeeSeswMjgblOhibCLQ
H+wih3rcdggu4a79iTLlARiAQkVAo1bY58uJClrJXqTR0qnge9L3Z9M4VUYtGWKs
P4yFcDtVNUpvW/bJ7jafXltdY/ukCeeh+WxQ1w4bkARs4x9AjjRULUHrdKT0TGCh
/1GLTZHXZNbRKEKDbmUABD8YICcsVJGpp16IlBmyWxUkC3d7+3Ps7KrT2BGmEuAA
rtFoKDSq8Exr0JXpJHqz79PWonwk4bR6fVoYzokV7ytInQcwxswrkCKhomu5wXjC
Hlx5KJtU+fkr/E1cDGDMUsC+Lk/YWQO6+WbdVY31rTmLzqbxyyrzaqJc0+MuTU1+
jodcnXxdaBc50YqxJrV7wLPLd22ZYCwGQZedvYsdJt82YcB4rTcX3PzdmLs3aCr8
hDeAW5p5ELGP1LkpGNzQkvCqYUIMaWTe2lbBJW7Q3DLSC5+LDrJgwuHHWLUGHdL7
mPS766cFod+qsUJhwhYSTp9rVAXYtg9BZpCs78m5GCPJK+/rVALJrbyVnCw9SzEI
MvnEaK5TWJjDActfIUSq2UE7slVkB2sxjYpRRO0Cv+prSBut5U0yXJ+z0jD/TL/y
cxAjqblKj0xqYareDGlrAdOR3t3VB59K8cR3M7gbX+QCZz3fq9fNZyEBH9/Tm/Z3
970+8EojloSrHEo3PUbqMwgCnCqGPgT6Glde+j8bRbRkKT1IneaLE0XtP/TWR/gh
fuY8ynjl6+SmUecxtXC7HNyRQ1KoUeDdAn34GpUF12ZhJhO9MMmUMFCvhhaOS7ie
r5N4+1pfKliHq9/FNHyyPV08g3ucUVA7uNHQcol9htoBsSacRm3qNckzBJE9Hbcf
2lShCsvDFjoYZ2KTmDQM/RpIGpaZlxVuQsqZTDq7WO4ZQBhQeMQGlJuS9oT4KLkA
AzCVIkdRHOkNo8QcWwRqbwiqwx6Gn0MO9Lt4joHVseTs9YiQ8z32tOwMs6ajCnFN
2ZCpT71n6wFPCsvi9zLevhxb9ar5eJPddzc2YSTWdsWxPIGwUlVKBqOFr4Z/02sT
dnnhrXB7RaWazro6dgvTU7FjPAhPFIffzJh3wZekaEQ/LVuet+vPj6mlnTt1n2bY
zRbTr0JNOpj4qbgqyYx/Xj35Q2LAChdgR7MH0xVdqzhedQNJJ2LmnG5QsOjcJT0q
LPKHiPs3zZxb4cyGdLEgCCfUWruhpcB0oBVdHmDLem7il78hA7JFmm55yNJJ+yRx
KdRdmcqAILqTnh+zyPmOeHVWtEa4NBABCQMOHe2q4kTojAoOb7Hygte9WqGnJYt/
eRr7Qz6+Hrzu2BPIs43dBEcQGgIuL8HN6CYWJh8dYq9bld43iJ4eHSTl40o91Eke
pwAL8L3Y0Od+4I6mwxZQax7b9pmqEmX22txP2xv/N8Bc1JFe8cFpULXRgm12uvWZ
6tjhzEy/p1Y/azEqv/O49JXGP/o3hR6UNsb0i/OxKx7QuRCXPJGkV4jmYonpcfUR
Gb7PpIOgSWRAvl3jZTeRm2hKQWOejwgLA5tQmhYMNNLUcqkQzQGWHfv6yHArgYax
FNnhgSqWLcY1DG165ptZhET8eoP4EjTUi4sULriapQ4ujEAaAPue16FRamo9ovhA
Q8R4wZUmD28bc85wm/R29t+tErlMJ4l6f/C0lotE/Tf8RwaDWtlpCWAP/+vm6Kta
DegssSmNL0W2954hhwL1e2TEP0yeOXa1+gEJtjZ/KXoSYbwHxVhcXpDVH4Fcx3Yo
lASrYbkccdpTNsSinnveBLwdOW3pXJDfCiPgsnljuXNLj3ZaGolOrRqgy6oJw/mT
a9ojYmbTSReb+gG1tqKJ03gaQRQqlJ4BnMhyK1YNyXCWCEcTJhAvSyn/UVJL5Y5S
332Khvx1LpP1rQZRGPAcOwRuPEYkGtiij0GtBImZ/i/liAhhMBHYnitLxHM1V9+a
u92uxhVYRdEonEcUkJ61cZ1IGU9LMDEtjX7R7QkjC/z5OWFVkIkv8A9CCsOrTEui
byQGIcYps73WMPmJKLL9MJVGjQnwKeEbFTdzYsVwvxdUhgreWHoJQD7/3Giic6DI
TY5+0pcvxij7Lr68LVTT7utw8IddmBCDxgixL8pKKDmXrOi5m4zboiuej19ZOWeJ
jK9XkSZtbbaDUSixaV94gw4QiKwGL4J1HQJq602HKyhXBnvb+SRhoYaR3P8q8Bsc
ezZTcn1rA7HkjcOAL6iSByHJZXiyCEqNVXBfqO1OkWIEvrEfIrPHWbv0MKEazf39
4Ap8Km3HT+GhHAIpZLL0LpIApUb5YpRM6q6e1gV/Gk6ARVaRzFsdMuiFAOazCHTT
9pybivTgxcElSh/Hf4lhlDu+x+WRUo0vZwwxL3rnDJAhBmumwBUKRX/ivyXaGDE/
WpwMqH8Xg0lCNDPcbk76iWr0o8O1AmK5D7vmw/SRbjgcW2Tcrj1xW0d/3naRmeMN
NyOPxgCEFCbNrO6Km0pgw7dIf1orF/2Bb8vgsswRYcRVAj5eHuuEDbu5elhLJo8w
iSZ8FE2/yruj4gn4myKqm8cPfOHABcclXUIrXGi98XIhqUgkQ7Uip/+ehVSsSa5r
syqxO73CbCjaeLQjMCWHB75cqMD4XTDXVIfNCqBZ7A7lB1my7d8dMikz7xcYGsc1
BujvbSEwOV2bbTAES4TMJWTIpv69dfYFAp+CkI3j25EsZ9q/jPbCGVuHWwhIA2pZ
jClumT981wxN/06rvbl9HM6wyuxG1XJ9QMj5NJUfmddkO19uQcEXqpcP6921b1cn
xkWhCkUIElQ4ppz5GsHhW2B9IYwZRHxPx+xThXXHia7zZlhdfkGSck3HfWU0XBlp
W3oTYkdr1P1u4chdyaE3LAMYtuyX+V0e19XWBo3rotg5ArR3c5mXgxh28WaNxxQD
TlYAduUtnve5/nKZ378N82vsEe8QtR6nof24LVF9t3/0K9uCuNjhNx/I3NqVH4Vm
eyYvf+Qrgq8ZeI5KCuzSDFih4wTd1tXB1PU3iFdJz3qrnjJ+uSnGzuka/EBbhfZd
kPUWeFrizQhXaI+AlfU6k97aWvH2zYOIN47YbTBgJEckxOwbudgz/fggbN2vvPK4
LJlSB9lrBasQV/GglPw5I1hOAEtmRLiSLgQCXKkap1UjShB5rivEw7UO21RwN6Qh
GAYpezzQTIqD06FsQ79K5v7MG8GAr/Ju90D+ffYcWxOxLzRWHkW0HbMVALgg22dD
E8ia5V1URkFNFni8zX0lJgdf53eBZd2JVhi513rWbYYtvqSxzpV04yUFc3MrCrLz
nUAAHop/xes/KZh8CF9FZw1QPkXsF8rxHdNagP69/BZA4VdlMkn9Zl58qs6Qa0LH
4/TZ6H0xvHyWeacnPJKhjAQaFwW1zv4+iCoTH7p4AxYciOP2SnfAJGYdQ8TLp5eI
pSfDmhxDCBiLZBNBVcyubFF8G4VXBy4JfDOWqwlgAr4nioECeN4n1LSA/geEL8Et
GaTts2ymvxnkbOJCO8IFG/WnWf3z1MEYRguctJNEwkK2LdHLQJRsvLf+c74wvO5e
qXnd/IHzpELSUC/SzPuHHe8AFPMPGdwD/haYMFiNyocE8cWdTySTHDweznFploc4
gEId/Q4TFeEODP2PGr6K7uw27gg3GVlhWL+zdQ6TrFH90nGYTvz19XsVtWoYth9l
S/FFrDiW1Lfco8o0RLjQbd4Szr2+aKZwmZ812G97AQvTP2a6UrKgMGaKJ29VzZZK
u4dbQw1SoHr/9tjYcgWegHnNmJ9x8Ch3anSvHsGPh5niAN0xMDxdujhef4L/eERy
xuGTYTuMUhDhFTjidCYqH8Cv7M38Q5Jgg9Z+aF+GlWSZyxdSDc8HxRf0WovwKxdi
4lD9omI6zA1veeY9vx6phtVv/6JdHYYtbWmp2ooUOsSioPsaODsgEIVoe9GmA7nu
RB3lpbe6JWGFfvFbpYo1ZPIeV8ORHaO1RSqazp7ksHCdhRwdgYIEAcf26A0VtfLD
voUSetmiOv87fMRcOX0MLX6MaRCD5nE+1TWHI8ELCHQndpuEzWiCf0LhEuAcARhF
qnZqqK+ygBwbUDFagGNvq6Ya4bIu1mwDIIB59TFGTxTkFEdmd9RuQGIt8ABHyomW
xJkD1gCmysP+ODMJKM1rn41Ur98p+0KekijwN5+pibQbPu2zAYVZWqt+uGZZ7dLw
PvA+lvdpDbtfPXLJyV014TBYJTqtZ109JnvZw+gtdfrGlFZ+aD80aSW9ox4fTTIj
GpIfaTyLTy9/79Zk1W+H3v+/BtEYCtyJJwXuFirnHuTYjy/LfJ9qLs2HRcNXJfH/
TDB84a1OXtX7qoCqBeoNMVWY85+2Z+qYQOdJGo3thLXO+C8Ro56TwLmYuhftIgy2
CJOb8wFpqa2kWuN5NzjVw5ZJbEsYUVUIv+tdWTkJz7dvpxGfoTYOHJwimfxExiQG
QSzaP/jMs28Pm/dRmW2HOi4qL3NDaLiHgkwMAvx8Qs8TH3H50W5q25GO+WC9ZP3Y
5yaRn6GzYJwakFxGmvtd5U8hD6BSnjj4dGBbuLDtsRtEfj65brcSyElTvlcPDn6/
jLUd2rcIZDlK3yoBwYYWmtMp94CHRkatkCJC47EHlGh5148fKW9VOtxvKjIMRKr8
9MeXv6hZ1jSZ7VkIRo22Z60kZxcwcNB/h7/pgOgZdpPe7+v0UNge2CL2nHK76+hu
7z4Eh0uMmrrDWVcraonN/MyKkYv6twblIJgAmQWMEjrXWcK1JU7/5FK2/Jn83gVO
l4OoZAno64rkPE4hewxImKzXsXjOCP+IHa5KR3bb66JhyKOsIeUh9FN92w2sOPql
3EVELWKpbK0KY00791PT4zU5v/W/bE688wH/LvZ88V/QRO8kN7UpCrdeArSj2EL+
teOLnyy6BPjYgT+H0i46z1Y6XK9MrAORf24MQ4kragPkLGW9n65h/0aRm3R7tfKI
MVLawngme/KvRIcUHpk3i+yhDNVbaMS9F19xG/I2eMYp/Dce2MDCKDSNEIQSKqlK
/H+d154BbYe5vg35W24yqrs9M8nttnAR7ZyHvLwA6twRnUhyGnFd0ccXAYZFEEXC
EIkS/g3Y51pB/4aNeF91YYM3IF6i9L6q1AEH1LzakYBiW+IqGkRREwXIh6/bqPQo
h0zh+CnhPHhdpVjrNhS7irX2pCUps+vZK8AT1yHh7DnXxE7pOAC5txq6tnw0NP79
IOIZRJQ07YS0USXDQMFnJWmP2dmUSUIXsc828lsB+epFi+TKeXOOdWAlrYCAv87/
j8Hq4FgnSOKvy2qDQ1j9PWYFS6E3a7LfiuabajwDKhUK7zkbLMs24pJ9O8sgs42C
QjB2VEYdAktCfEPP2k8AZ0MpJ9inrsgwdmLJ49VkFYxp5gkUFx6ivwsyhhQ8Pyrt
tChj1D3tZ5aURJDipIl0gmDrWKELfJmaSecky4qNlN0fY3stjbwueYJ7JjzaEj+E
todlkCl69c21wWkKWC6syMNqD15KzXu0hiHcmOzrN94dXsgswUiGzZSw/L2hlCB8
/1NbcblcLmV89vs/l4yTqi6KHzft/o6pbk1/+YWekR7MAND5Wx2YK4MiEjOb6Mq7
hauneWCuOtjV+eU4dmCF4XCulk4XjL/tlykTd51x69rwwP7Tv30+mTlmGvqoEEz0
SUgZxVvM0BbfqQjRmPoTZKEPp6CmgGLciOCnnEp/4THx5uChKvVfjO1Zb0r5Oq8M
ev2uiPPWIv4JN0naF/3pw1NEcPHw0NkZBPU+nizhH9knHnfNRPo/ULLa90mj+jxE
hP0Bjgg7/v+/g/E79V0WrB7Gxz3nOj9n2ZlM+S44yKRkNncsbyKfwGkgftHHDjBI
+j0+94FLRdKcsPSXBl71gj0uuSFrjrfK6oSepBkrH63H/ZeeCP2xb7AiAi6q+IIT
5FEqeqUb9WdgZ/97DcyGkSwCP6GZMi2lws9l4rXGNH+3bWZ5v/enGhmBU1AobRwV
w1yeXo0INUN9OWBYnX7/r/vZBh7oRjOG49GGJ/yOOlJn7wU1mcYGFAXxX2hmbdmV
AJBa8frGwNFCw2Wu1G8gaZPqXW2U7vmZzrmjyD7zApaYKvq5tgfXFvZvSnhTOw9w
mRLTw906H95GBh/NQ5vzc0vFlXdlGk5WTvOvyBkz7Y4M9iLo485DJ8iE+yw8xkB0
BJ1YNoXjPI+aX3bo4isy33F9mVz1rn+4++02bFA416RpZSkWZWoofH2u9uWq4BUo
62vhuwPOLHOiPyh7GafqoUnaMZ5rN2/fXx32ZZFRD9sS8Onpld6UouQNOgIDqlmZ
SSv1on4lKK0JNYrEdYV9Jy+WPHsQGxjTBKG8qtqXtnjBhAbS+7e4xbgW0IgbKM95
AZSAjWkWMHQprbetMER0GlE+KIyJk4etQAqHoiwx/9VoKlIstEJs2ZvTaAYVLl3H
VZcQvCnizNlpRiCpIh+FedPEETLsewRKRUBsOj1vyAzvSZvr3TMGma2UCTAg/CQv
NNCm9NC51Cj82+0wBuuoDNZXPyPCUAhOHhTUoKbj1Z2V2wyE9QM6xnacaMYgMEM/
8h/Nab3u3/GQdXjbWtAowBcruvMzCcPYOW/ZYsauPbId4JD2I1IgbKhBiSTyyxg/
3RWw78oQMGk6VhT7aciXLM0M4DFRZPO+mBK5C5Ws+Ai1fNsvjyeWQD+plrJjdUnm
k5XRQQLd/27jbvrHxu/dLzGH9M5Co3G9x49R5gRVQEuLYLsMEmIeuV10FXf1ExTE
Xoxjc7hOmiKVIucC06DQuDpnHSijHFnQsSMZEIlpvlOr/iVcyy5Pj+MiA+G1D3bY
7cQpvXI2+1WVsMIrpkebVQvuMZM7LLa6DJ56qpth4wo3vLpoYZFO8+61duXWRxwE
tCKj11c/JjsSlWS1e64bNn/AnhdXfJwMzvY0lRtKudh7O6lYB95A/G2yPKXIW+K4
5+PN+KEP6qVxdLCMeL3aPRvN/DZs3wkyTceWmZcNrCz+T7FSyayyL9Z1Kv5V6MJE
DhvsrvGPPRfobrho20ZPNRGbVJrR8XJZhfcaBrKmX8CjjT6DDE8j2M+d0TDNaMPk
r8NjBm3xuFzmZsXk5FA6QdoH7aL57Cbmcg9DkWkro9Tdx19t7k091FQf2gQMjBd5
op6mFQeANEeToY9Tpk8MZh3hWuB6bVc08N3RdzAge+o7tJG3+HBjKGTvvLkfUjXx
hP2tiSpqeVr81r3WkRltcoo/OwwDWaktLRHubRK35lfsszR1ITJFNrJ1K2B+r59J
UzsBrt5xAJfVr0p/2Yb5ec+Q7kCEu+JKcCKNI5lXYbsF//ZIO2ZlUOGu2NGlZvM5
nc1SrnQ7EIvEkf7ZhfGIwSwbht9hpGid3rMqWOFmt1u3LuM4+BiWD1zujBBulbFR
8vvdqrAxrrnEKLG6ELekzJiMjdvd1GzIs6ORg7QldACdlMiwPanxSug8BQllFHgW
ceSqcXXFTUC4i9izUQK7oZpIR/gZ9GrSVhrtQLOU3ihFw1RLmyOxwVYULe6Q1QaF
Jay+c62HDld5mCN0/tL65nxRRQ9U+W9yCEoDITMWRvNq2vJGIYD8GViLyiAzj2Xi
y91PkLNZaGV7HwRp1TDQrjynhJ7se5qcahUY76DmG2pVvD9b1KbGsRidlQn08cxb
ZYoag3zxbAAnMc9R3Jiv/OIgT8yyhU+WL6pIy1GyemAIlIQJHDdY3e0fo3NqSuL9
TaL4IhCFBbh+vhGuJU3+r2jRZBvsviyHLTkn3wCqG70XyQrObuhA8MviUV7mvNEd
UUJfgjkmI1oX2HhTXlIfH+ZuWKnFLvdWhgDsooqtyGqYzF5CZGMKVkHwKXcngHIB
VAB+ag15tJB1JGKFCGYFQWZ7JDhYa5uXk1FA9eb6NpG4IL4UDGtJpX1PJaiI+10Y
+a+wOa4LDo04q/9xa7UVLqF1G/GDBHISTjB08LQsEQmdAV8Aag9GxWvQlO4ZC7yl
Ggr+eD/ncKI/Ejr3yky17y/M2DcDf1sRwjsRC63ZuGX0sr2kfwUtlWIG7pl4N3Yk
uOJVqH/PDW6s4nf138qts3gQ900s17f8gFAqB3HaB8y7S9XVahUTTQxfrtdbz/DU
zN8TSFbCRTRK1R0TxkgeLgqZ5RWtIqgDgGiMrdO9xUL5PAO6zx2RSZL0D3rW0Opf
VxxIoTz4VIhsHpK+NBF8n/+6RKKqupQ5iN+463iviIyvQGjNiv5Ti7PuFUY1MaEl
9odc6mHbWuJU8p5/9KFn+I76R4y4Dgl6FQAVRmjToMGoOX0RymJy8Bufxl8Wa2fu
hVVemFRcSGtknoGZscNwUz5USbuQU9/EYSRI9JPfs7NLeUPdYYvY/BxlrWe0FCMk
jEvHHAgoKii+6EHfFfdLt61RTx5kR+3Il1elgj3ct2oUxYwt4TzJRTpG0IMl5j3m
b+HbOJ9tcnUSvZTRyFjHMQ9nmip2KXfpdeKVqoVEIDWfmQ62uigeJvgbw3Z/KjTf
xgDfzMZzuyW5uVlvIJPMSskdBPmLQodRtU+a7oIXLldgH0SrT7YmAZT6cQ1Mm3vZ
Jyb1KLHXUwjzi1NfnQOiCz883jAX1KtQGx6RFB5HmZ5gZ/A7DUY/kCy2CDSJrb+Q
j+8Yx4rXPDM8xwrCtdA4n+vtJ5qBbsVmJYZIemb5cghlxmcw1nlalI5rXQ8wys+J
vQZDepPSMIdTk8guzuOYEp77y1DkBq7rWZ4XBzPTt4EDkIZZsRomdkogaKSRIYyF
VdEvQsLSYlfVpDL0ygxSzCsohnjbP75YUzrrd3CdHwVQNKCR0a6QgE1Oc1mSxtSy
ouPBYeLy36DybDOjmo1vpJamubBhT3QhgNOFw6zJoZxfTpE1mYa4U+El/mpJs5kT
SWAsP7syT+5+l7BK6jVmFJz1MQbYeLUbkrMXTDaq4xITe191bDyt3JPg4U6lXI8A
FctV59FdJbX46rqlZv8lJKEg0uH+seNbf0fLadP1yD4CkMXaWCwL7CH+Qmky3LmB
ZFGsR7cU36+cgYesQeWOZobNSZHltyrrrQe60WGYWxiCaKuM7Hal8vuVjbV5hRjY
66eANRhksujO2eBh/ho3VVY20yAfeFpxuxakDHxwx94AHlUldFQKQHKKz0dTDjP2
HjqD0Qad1ensC+XlUU7pWFGHQ9EoleGiPhb7Odf8djwVDWxyF2reUzfQlwaDYKVt
RpleJJudsiTEvk7f5TSZEy7oLBP8930FoGLVpSZWI4qjpw/0d3Nnc9Yru3Bevrg8
bBbQ+312a6clCnvCuhQol4kU9tc6XyRjO6AP/aJMwq3lPBeEzEJSopPKt7g9JeLu
YloEORVRkXqMMsCzRjfZyACuJtMaPU6Erhx24wew3W6P8Wma32bEZeSVne4FjRbd
TUHla96Je37bbsZtcD4k8uLSsP8NEl8cEktFkeGIkui2jC1UNBnYh3XJJmA4FdLW
V9W4iZFgn58LKkf4QxJCsG2xtMx5mlujTg3mb1i5jml2fnRVpnkHLkcJJHF8Taqb
0iOngT39iM75hdinDIRlaFvHtUASu6ZGbattxWpb+zm9clyKqGcqwHqj+XIQ8eV/
Dg+EAH1EFnfGs/xh3XvZ/Q32rnID1PgS6ygMUlrRwAEXxeBM3WIa55Si/nD+VEeG
Tnm4D7Z6kJAid7VUTZMbiaAeMtDZ2eR2FfvrisEcrPsP+/6Mb6HV0qdSmr4PGSlH
iLYA0XRfgoSaNn7iNINty4gEMvLbHECAht1Lf/ibU9xa1j+sAclUxOTSL/4TtCNg
7gnOPuU2HrHFvWb3I7rFg4lA9mxeXw0DUE7h6lihOXvtnsDQkMoxiXsAFNJHODdi
Wad64rrm88QuWcZuboHPCNJ1vVtaYG0SGGdtTW7kBj7XjKhsH7OJGLnBBm1t+/Dw
JeuRpjX78BcaYub/tPKiEfLPzYcnCpkS3t7H4QFsJeHN0od4Yd7O3e14L+yFMbkN
0ZpLIUpIEGP0C9A0/Z3XwiKD4J6QlRngVLFkrl/YEDy/Y6E3glyTJ8/Q8LDfMDx4
pYI8mcjNBCTTFFi1uBFm+kZ31joJ58/REVzG4jebUMYLTzpDMDYh/b8mxt/LqA3y
ZFBN9iIlfQOhv3Mwj2bx1ApG7f3Bozs+NjMR1/54lXnzWLc51V9wK5j5nSYKqw2A
Brbu5vsv5FHknZo84F9QXRzqWSvwWXT1swPnO1wt3JqnC0qiOJODvLm/Qe6bZguG
6317eMAqRNiuqPi/HxiRmYNiiy/uxFFEAs18iT4WGXyO1noUeuMK1bndnalryLPc
smmkoSeqZ+XXlklkcJ68PwALTonvRQdZeBfsUr8pjQNgLGXnxuXqWkg3c14XI9Ab
Uf5eHJavNol4dehm0xPijCZubGv/jkJmLvsmo2h3Aw42eMmZa1b1Z8a48kOagY2U
7jI85PUWuJnXsOonZ4D+/c/vr2zOoE0ZhDSSqQuIOf8wXOTxyvbBHjubMnT+NAxo
DZ36PiF4GG1mVr90B1aUmVpRFAYo91v/8jXYGp2eFR+IdYYqyOFmlZM+h+u79KQQ
RKplK7ELCBd7GDhCe+EklsK+PwrkWgtY3hRErY2fqNVLf4H1jaNGf5lgAbI+pjTk
js60eHr9/jizfbs5DppDX0X5IuV4wDahPCMBnLIfKPueXq1XuYkact7g4Rwr6YjM
n7mBFf05O152vYfeUUmDeaGYm3bfHi0KILhOrJxlauiZhVp04X0mj8CWlTCFwp8O
XvaWVw3+wyMlKyGbfg+0PowEKnP95ruqtPA+E+nc36c4FdA1/TxAIFgY5/TL4vVZ
RGQHeH7ecqjArR714tDolJ6Ddq4qo9C/jf9XajYS54LwV6sg2G56BLsBNXydERD9
ximIKPs1DQlPcts3udEnf00wjOyAqmokkyypQxy3BzItcAcoHf6LdIsOdiDJR88v
SDTcP4Ze+hr/HV82vqT7BKioPtwEOlDNF8QqJmHt2jwrefvCRFRxJytSEPOXldFX
/DmQn+vxxwaXWR0ijtK+osW0rUwAhxsrUW0+Y3tO1AfLOyN9o1R3IWDChovLF0Uv
OPDwD5W/qbtVHuu+505ztiQb39NtHnpcXCL7KBjiEtHAVV+k6ruCQJ9AyX+m65jA
oUrHIjy7kB4cRGv7OkT5rJUzfomULcqiUNB3JEclBUBdv614hAsQcCRY+Ne3NSDX
10nfuQcxvqv43i1pCgRwYDMSC1Wmqb6TUVDaM9ay0IG/4P0GOthLppEWYR1jChUg
OElel4yMyywjrTp0JQAn7d03Hi0CSrEoQ7fOLbzXZzgAzba/uuFm0kqfiV0prwbQ
Fc/bN8dC0A61IzKu8ITQnFCe6qI8VLt0B5boc+CkH7N9ErJcH0/zRp25xX2s7CeT
tLz7SLoT85qa0kbdw6F5y9dnsw7lvE+zlL2s5V37GQAgvsd6tELUgRn+t0EZCjp8
jphM/AaOx9EuWhvbH/NfrdjdUJ2hFvR6A2ckAFtZ0rh+4gv3JxIA47IZMkI1Slwh
ETBOKN6hLphwYBKceJe5FG0DguPEBZjAB+loFd+BfOe6w3U7vOFWC7V3rgYACHma
3YCLhvZESzUFopQzHFGoZeX8k51q6LAV7mH+iDxuaTsNECaAFPBgZgAPn7h5E6fV
rNOPslyjpwYUTYelY8z/ofGol6iB00KZ1hTzy796Gdf7GEK1+SHqtpfD+Bc4ov1f
zJAwy8U661+OC51gjYyDOFVnlBqiL7WwSIkBRWP2/paW7CzONtr+Wyi//23HpQUA
b0UeVnH01gC+v8D3JA2sutDT6oCk6XhaROg+e46KTSMPST0t9HW1jzGv8SThJ3ql
lLd3ZV7AU7pBfTb2YKzKWJaM5yKbPj1NxCKPZ+rywxanakudQ/CmfeAvuscXmLCI
2mdMz9wNLIeGzHyr+UWYxYFw36DgIN63DZBETFAq/jyuD/MT9dN352Kc+B3mNBHN
V+O45hmTtkov+F8Tb5HKaubw5p3e3cIj67yvu3gOS3XIQLV2Gd/X8tw9c3LcdjZt
HW8tmgpdH0PjOkij+y7BINVMFuU6SUTwD+ZmItXW+FIImRbSpCJHGsNjG1m7Qhzp
Q9O5o+MaUnVxCDlqyfA/C0uuMqYQ+tSH5p2+Tx+VSCcH6mDVFkc6TxA2hGo8Vm8x
F1xdg7rx6BPrg2YcCN+IHGvhEW7B3nMbaQ3d0Xo9e034VFJxcoWR2nT6i42RvKn8
xP34yhRTrTvvXu57L3s/uQgM3X7Ga8411vqQv7SJFwnVPN0jQ3hhPAR5o/lLT1fF
dCfxEzIThHVwC2u+fq96MJbZ9nfLAGsI5zy2uTqaIbwFeSMUanRPGLqOqxzAM1Ec
SC2NfMYhghZwsm3Jd0Gbjy3OT0FdIpRUXLxdHyGBih4k9hpkF4tyWREmedU1MFKj
b9EmoWCZcFJS2ilrz4sEEnvNGwi0C6tsQkQuF4CalJI1A/9XHeeDXlS/c3vystva
WDVj36PbeJA/gZNaxK0pWcjeX/D7s0myzXbOCl5MHymwyIQ0X+qP2K0VuurjpgQw
TwK1YFLrwR6H6vYB/tL9fYclO7GJUxiEiCptisazeC9aB5rtFn3qOArTGyc7Ju+B
hS0PX5FzXE6E9eFwM0IvFciPSMxmPs2TihItIfLUVB5r9GIlnNkZU+930FNk+6el
eQJCejRtfYEXGdvaOJ4POuua7EbdeH6ARCB8uqVbWUdXwqIvd3XYMTMtlKMY+087
F1zdOe4Jzi5BTKNcmg03AWTpjxaHcKahBS0dzdtGC89oXSRKV++PGmb/0i7EWV87
TlYcJ8EAmdjcMDY8mYXVAVA6R5POWze/0MiI0Ea3A6awR02pozJc2kjnGlzJUC6I
OQB4j+lZ/TqIl585rPTiRHDAMg9csWEk4+ABjDEzVWlEEU2phkQd9phQozDrpDJA
gU8RY/iakH1t+l4K2yKZ3G6bB0dv/Sveb6Qqx0uUDFEQQ0T0gaxQYX7x57a6WyRT
l1HcGBvRvPh+0nxcs/dZTI4P0JdKTpcKeALsUVwHfw4KqCTTibGIAIZvFKKPM5DH
D/XlD6NjdGx6QEzp8dso4mNObnmwFFamn1yA7BV5VuQdH99n3NerYeXzb0r/0j7D
jIaLPx9PNdKKGlZVUsXMEpySRLPt4k5jAsSotYkLj0udNK1G573t7Fpu86zDNCYI
lbAdExuLkqjOjJpchwgt/TwxnjZ0J4vjtV0bfUEjDYDItYS6BTX3EKCXUKnl1f98
fyy6uyem9CmudimY3iKQqIQcgO5QHdwdkIo3cWhKssxvmEPvXCxg6gFCYIx5ymfC
9QS4O1SFqX3Jl1PfZKP76oQ5spNgGn0XFxIWNFTBPixNMf4MHRsZos9BLZ9TeKAf
4mgEEuSVzu/2A2w/1zlVz/LeC1InaQDMFVjs7etUMwckqSDUNJH0EqlBga4ObmvJ
bZFLQbkg8o++kTyYVK7WK99ijSHFsyxPz60nJM1zKPVv0hMukM1m0csvmE1N69aF
RniQt2qblcaNSCCsIc0gaGDB9xAYNeblDAHMNmwwh2jMj4y8zMCDXsWVxU1N5q/j
D36TYlHw0OwF/i1boWEcF/5QjMHc9i5RIJ9YXVJZ3AqIhamNhiKqyt2LWN2CKRrS
/lpQt35jyDMcn46zOr0BkflW+PCDcPzUVEoyB05j8/XtdbctGz0meXYDpfgna6DG
CzxM/0csYYUdl5fivtP2fhY7FhkCbpbTsmAer5lQ+GVAI6bxpqv5HJaxxHgX1GM8
RDv/Pn1S1gZ8e4Sccsth0kYWs4+5XV4OD+EHLOfuYhT000pcdp+rOw1nGmRijo0B
bqrwl/6ZpeRdW+4LieEnZ2WqNIWA6Ch8bInRyYGD8uR4+qYSEilD+zT6z2Qo+awC
+SdgedvEyBG13DTcE8DLEPd8rxj2AzuIhuP1p+XcDiW3d4VYDlwGubtKeere35P+
hmFlZMp3ErhvnF2rJBtMPw0uQEEIkZ62/mqHSk4OD3ntcWpEWLehZCOFAYUO7wcr
LTdmsnc7cu8k1bLUjo/LFJXCN3K7Uw1xneaXVS/XMTckXDxFulIt+Adka3ARXA6f
scTNfB2cUy1MQG4/hmGbLxt+5k5N1jPr6hOf/AYQNWxaApl2MG/zsjKpmqZXk0ZC
FWGXMPTCNQRV9wI/twL8qNrP5qn82FWXn1JhtlShepjUlt93ohfVu25YIvRSmIad
nTpEEYHFGy0iD4TCFNJCozs16kioVWPXyotUWCuE0R3a8j+9onedN3i0+dgjU0Ee
1x2MlUXlPyOhkrfL5A0h0lgmSak/k8fF3TAztBqpCgIV0Yy7XAwcVNpPo/V/ZnXS
MAc+Jn5lPoMWwXy4IqYI+aXg2v5mNPmbeR2mHRnVCsje4CoEJIBmNNWRQ41NqE+A
qva59obaplpYUpY5aZRY0vLXjLpAWUNXpIuHPRXMCNbFgpSTxwjKLgkYryk2a1+j
oIe5c+H0wxkBvxcI3YvBES/nsch6fFoYRd1ny5oabqppn4MQHQNrNizoSbIj4wnF
avWf9rXpw2j6XPY5Li63BP7LAGIyfTtE8B/BICPwR5+Zg4eKNZL3ETFiQGaRO/qy
j9gDdkHnhiMEbNJmAQrdmBzVvOly4gw2Bmk5Ly+zzKUv9lSKBaxTVoERAzoy/YD9
m/b4GdzwHB9wkYaSi5xOxsThqznJEG+jyzFaCR67mEJPEu1rFY48+A/31WvIzzd+
CWvc2RAUOw2cLwscRveiNm7/iubKweuy7q+R6sAcmwHEwuuJHrBbEBywJxHaz60/
NK5+S5BHoOMg1wZXJEMchYDRBUnDqJYtcULR8x49vzKzFbJAhnpVEaTJXSd+nhGr
QjKJD/C1JpPQCv9KEvTB54HzwCu+Tv6kyFcHFyBDvdHtmGvU3rVyWzW3oiOOVnC1
1sGLpXFbipgjoB4qqVxQyy5FTYF4Ix45H+CYXDEQwESIsSrwoEwlPmBgJ7Xwov3m
knKWin/fFWkKFYiKj15a94KZBQ8SA0ho7PvqUXjE6zQw1pWRi76LcdcIY0eysfLx
wlAZ4JZ/8/SgYN2BXFm+cGXpi/XQadjQqF7uMnXzWItxrfWm166DSy5/3lOQjgOw
h1uaZ79lFkljtSz1EmI35w==
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UGqwjIJ92wlxEVSqMs50zhFBbtInRjWPsaVa2/HYVF7Gx6wilbxAd58JV65mPmHf
fg3kCQ2RqM1V8ZXkc0JGra/Aku4oa9sYd/ZON/Exm6THZtULqIge7tDZnblz4f2k
KxGHQ5zoJMxQ/6PxZ4gN2tNKGKJCMhXEUUFVYlVNmKbvTYt3Wrz0zfOu/lADmqud
MPsRTTKvhKGmG4Pu2JTMS9ssv4PQDpQ9CH/cmPF3Nk2PjTdoBFmvYTbGzUSxngUl
sGelfJpU3/7vU26weUSekX3X9Yp86hbY8RySx57z23chf78iI09QoLlJ75ZtAYVH
0zOZAgoyOSy3k97t+UHpNg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5104 )
`pragma protect data_block
KfmPqrOqmyYf2mBHklB0gXguPqJ9cULiMillC667AB0/nMBQRWWXGNyeaSObkp3U
OY+XW4tOzFn+DZqbQHWhBtX4Ot1MfYp6t869y+YqZS6t3aeqHNDrim6Ej/gqnbIU
eS7QYLcZoStaUkI0Q9o9v0gov3GjXG7wGWjQ6/NNlMZhsrVlZF75T/O66c0VoQU2
0VWyh6nrJMTbyEvc0qcU7P6u31v6sHxzl7cVpeW2JS2dDZ2oOM2tcAjuxIg783Pk
wGbhBAaATPwbs/25Fl++xRZVj8su9hKRE+rcy/Z8bsR9V9t8S5ewsx4Ga///OoP8
c4wirGGSYbfABB68108pbLs/bD+CDzEJ7v6ky5viSKZtRkF99IVYKQ2yRU2AxTRc
WJm7HrkNUFhFzi1KAWxCSCAD0WSC7nKp0a0+guyEPvrZkklR61zMSPTOFqF5oWjN
pis7TsYADvHWImlJfvCsk6R/yWOqm0s+QKmoRiAvA/fTGP8TKp91DLPmKgWfiu9v
5e7Zy5Ct5vuZbD7NKYsWVdPGy2A8HSnIoZrgQOxMvOiuWfFGwjmFOlEDXnkk8FjP
toSjEpcBKvK66JGRBGqVtDDhm0HVS1TpLb8UJ1gPms5Sa7owYEAHCsmSP1i3xsNA
7IUCP0ow1gevtgv2fUvm1OtgYphvYx7qu6/JUo4Sv9FcUfH6O6mZ1gsWtXg8UBMa
BGlChhsIS97TYUzjFdCkRgInFrXS82XGfhlc+8GM0enigKztqMOlKOqpbnEBDX+r
+igmvDttJdBISuhN6rjBSawwDL6vDOcVj49Qd5sbDekVNNCDHWXCL3l2ukmNiYq7
9LHS7Dha+BbzHz3Jj5VHyKz3PVfUbzveZ8Le1RWk1PXhdaOvcJUCYzIf9teqdgIU
AXJM9usT02rLxKKaDS82WmWerz6PHYjv/Ttm775pReNPaJLV8ghRRRjiVVLKtsP8
HkBkwVAWwXIH1g3gs72G+AkBmNpwuBq+20w0a879x+BrN85KH4ZonI1watjCDZer
mtPoOIWgOcsklMCRN683L8ND66ncrkev6PQmYCD1Z4sSGbdLqIQtIQ2zRWN/Qal9
BZV5EVXmlLKd5MSD1KXDusbncyGTcJ9FBTjQ0vJUP1JS/TuSHymthW0L++3VWtYK
K8Yp4QEUreL4TydqAB8mRC9uVvJzb/f2OKfpVg4q21De59ZqUB/z+Q38Kh8mGoBu
MXnT2eRNt/etFaDnzB68LisAxSaCwAzisTZLExoR8c0+fLB4kgdImgfI+Dq76y90
V3wQ5KHi7S7K19mQNawkkIcHMCtyQzweBsyqK7POJnqiLAu6wYcmodXC7eTZtjzy
dAX0GhCnu4+mBO6TNqd1HPk3qeKljMvbRvaOQf9NkkDg9Hl/RGFkPQMiyXVwv3VV
H6i1i2Anysd0O+fHee/zsN6WNczhZBW/Ve9JBswiY5XVb6SPPCemk/tLS4WFP0TO
D+mYN+xRg3xzT7znCFOyAOnlppQIRBPQwYAH1wOTZf0XioDzBM9jnaBnCZ6mhDUw
med2eaTfVAUXY5wmr+Bb2elFQbH+FjVaHEwuW8Ku1Kr8zCL/Z1J4Yy9T9zfQUqvj
8Z+9U5mYPQLZgEIygbrkilG6VSUqBQY9KfE5xS+k5VEp2YQitHgblOu+oXXL2lm6
AVev23Z1IW0X0i9+ZQfzGhrYB0FxZSt3IzVuZFyaADqYsC+xyPRFJ5AYs+HwbtHr
3vfu+2eDDeDlXuXNrfKQDOGDHhT4xsLh1Zl0dNEvWBvr+WpNxNACe6/CbmcS/3uy
ZZGslUrB+b8VAgZbjJzJu20iV3k0vw9Q7sGgMdmuDPkMzC6sT+Je2zQ3akUpaC5G
6ccjugUVUeOD8obHdjbwDiqXmaX+VF6gFetyxVLxczBrg30ItIVGr8MBwvlFHP7Y
XLUwg266tuBSOJFWN/vrU8AoOzbNp/Icl1d3aERYNUbCKdRv3fn9AL4ujqyMheil
LHSOhdH90tMBsdJbudqIB0CjZrZXMSj+rLn/z//Y8NAlKISOdMQFMvXtgoG+iXDw
IMZHpxmjjAGv2jZ9/FG70x5WkpHYuutIlJFt5u852uyt9Qpyla1vQCkLwUnmUcF1
9oX7DpWU7lVxSD8FSN7dP/s66oUvQJ2vTfe8/IZizllaEItfUhh3J1+xmPJ/KerX
qiC13UY+gqR/ZgdkOlIS47tqqxzN1+yaqkR5hKsWQxdUZL1XB2dHZq+lhjbrYoNn
n/3S3CLUl5tWyS1R42alL3unTBUhhSHdS9NSMOHvzXgQnI5ydb4dbCxWSViqHgTN
c+DceWv977EBSiQHDpFUOeDqbfHSr2EGQZTeF2+uKlJrKWlCYymdonfCbDP0FwoO
f3NbkjGHydQqW8VNHjmBsGV7Nj6V7EyDfnBY7dQwqIZHMdNhJ0w9rQI7p1WaCrm5
0W8W2nMcg/qrC/cS0PGbkHgXgGjf8o2qrfKBOesXuUlohQaLXKeIaNa9kgYj1yv5
0WjPltSziCScq4GLuYMcYRb2BwW+4picsFXUY66GLaL2ZM8xjR9lYSw8hw3G1rnA
ypxWQs0+GqKwYYz8GwBBMv2799jOtk/k5iWvYdXsjjpp7yTfntNrIcc3zf3fyPS/
qyZP2cA4het5SmSi03oZjC/iZ/x65IEjCBrUL/j33shBCnc3cdElGkfax80Rquox
GTDYIt+NYfrVTjLMC4YB3SszahhhzZb/XXcNNVWPzxtUDFymVcQ37P9s/olvkKZP
jVqjrBl/4bS0UPGuWH+M+FQQn9QrquRKglHtMx30E912IDnJvEhZEgr4/AQoZQm0
1mePd20UwI6aLz7WJRhPtC3fLFkECwYb/ho9pAKT6vazEz7oeCwACFGaoSRUmzME
pBhzE/0j3CEz10FhqD06EhSOroKeOrdpICVbXFFfbCK7S0YWmoK36orzM6iYcPmK
pgb3ns8kjWfdBkwN50p/yTSZ6iDaxeDWuyhGXEOCsQKUS2bu0SL3DGBkrvtW/8Jk
3Rhmb+SemRsulwAhmrpeIN6XPvD0mfyAuf+Ib+zDXDW7QAyPwokKq3VLiBF48kB3
dXy2g2kkwRk+OV76nnspxEVmlOI7O7VLAISKnlhMFTa0vDdah8WTtP3HKh21u/LN
xX3F0K5suuV+kFx+Pgr//hSIhgZvARCZEnZVjBhx3//Qj9nXF3cwKUZQJ1jyqIRS
MYm84eJGBiDPT/eri0e6lUOZOeflc1V4idV4bE4shBKZfyTwzNaCKSYP8WXJPdn4
OGgvHc1K79VLBYKd50v0F1LYg4GX1QWwfWiL/mTPaHfy3R8xZO29/RYlGtGjbKeA
flYu4TsXJnsUxSpx83RFzk3kR/3hhy+plC4MZWW69ZRAGZ7WR3+ffMmAs1qLzJY8
yKIDaBqr2TA1wqJcAuOjeJmTIzSgLPQC/jr3XzsAM+UAGjp8e2R6vzon4eajFjJz
0VrMZJVQVFwVubYEXKlYgAYO916l7v0AOCuYXN5neTwDWuWkgmPArFtWvjFIm0yO
XXv8nxNToxnKRamX5PFnCE6SE3gz/3E4mGjBJrLCu+jiIwRaiZjbyc9yFiZzRnSW
UxHoCEnPLbVEfz8l0Zw8uyFWMnJS31iq8XQR3POnWzBawLOPJ3psNqnksKNcUyiC
bVtNZn7xHEbd1d/HCcb/DsasXXf8wV5aHOFRpMvbyE2a59MOyYSPPgtabYKgAY6n
Sol+8/+mFWU7AYOef6lMup/2d9bE15PzHEWrURr2GHG8Zaqdk8nrWr8dHcT7mGT1
X88qYdaNNS+K30Y2J3iRG5NR5tVEEpOH06O0FnG1HZGoIRF0rmdI+AyZ4EbKKUpX
sNaP0jG3PDRpc6v6imYLzOfdp9PTbIp4n2WtzXuP4FMFPl/F0oVfyHENqg+/zewZ
/gLuv/xNGV7h3xMLFPU4IrRxVVCK3YZHWsTtTAv+Yas74MCN90yCpj6mUUYWzu0n
OFhwOwk7rFoEVfzCTDKpxqEtVkLIV7+M+upHISWHIfUU5DarjNWHUDpO1kLqoYKL
eUGWO/iRowOv8ssfZsapHf8pcbkVTVqElbuT7RVM3LB95zWWqjvlr5Skh8G5grln
AI/ybjWmLE8hYf2UDJRAmst8oKY6Bo5eukTXOkUhSzu/flIlBlYfccmuBbyikf1s
pCgUK7DR0MdSUe3xLHJ88cKSPnwy5Mn25FBJU+k8fDlOZVFoiivuyHe6GGrk3Y7+
bvJF/JBTrzhnPRZyATHukqH8s0t2NTaNz2TUJHEs5ItSpnnMYkTHUY3TDOrOuQjO
g4VTP31vJ+UpB2o9ygL5dhZbcl5JXR5ZrVA2ZAYTL4hv4CWktsAuO0x3N/SlTIb0
Hvd68FuJ/cSS+8TWYQe3zd3sGjj00Zeb80umHsDtzSZzooe76be+wnagIYqYpKYH
0Y4e926dRDk+wgf9uozGI9hAczfLYfnjnWcW8ExksFuWLTq1Vqp24VP/Y3D4xbs7
ZEycdg/nWQgLkFVRwmeHN7q3hxpx7+N0YrEeK6+gK4PElWkKPDtp9nKgfcCE37DE
hMnOvS1W4lX4kzIcSEcEF9LwuYd6AyV3XvHSv0omPWaayzFCOR+NS2u6piFabP0a
7il9fhCV7sIFSyP0DcZF10ZmZuWOaFm6CheAIx+S5nZ+Y51lpXy7tO6l0bZpfNRp
uEOT3Cy6d3sHnPqWW55hMpbonxfo+4KPBx5GYMMIZBYs+wOnGDAj8JHhZtbPWcib
Va2+yQeUWd54ujMUxRw5SZ1B651xNdCKFWWK8w3d6tkdyjY6Mt80eOn6kwOQwHQJ
0kKbbmlbLDTzOQV/J5EaYsoLtwE2Bjg5pUeC9kN5UQq70+SOUmQ8mlOMzjpY0CR0
0lilt76uIo+MnQENGThjHmPTthW1PgVgVKZnW9/ynprAfaxLT3IHvq7TDDYf4c9X
9qKYoF6ox3jmTb/R5bnr7OsjIhLXwkjnOsKitRV6aFHgpQ7PpYEI2CO/50b5SokS
JDWwBUNOfAgls64ckOBW2Jta4N15PVwdGJS3nYn+AFz8uwynHL8oz5Kmq+LIillE
badM86gFU+TBPfm7zJtMWZg1tvh5Fy+8lEP1ONL0UtJBatlGq/hquioUpIUEaqX9
W3rMXoYrpFu3RR4du5bI3iZmPz866Q3CSd6lFmWm/dh9DAFikG1NNmyD11+jvTec
o7zp3mOck2ORPxhnNRCAR6++ttHnVzBnYxZ0h6ViialVXIRNls/oN2TVslzUr5iQ
7teQ0c9Q+13pVHSfXtGaOECTTo7E3PgqqCIq1jd/4wwUvP27/aDXA8/pmrBY7hDf
8xuUzMBPQSVyKN3dwd+ypjfN60CMlt6w3j89I+/kKyqPqcV4v6mcrVxvil+gCruM
8GCnH0W/iX2onLz4Jz56/wCOVcG/EC2XvjBwCEUjMsABOCxfiPVlph2FX0XWucVH
UV3QALdwgFDdVEdXRY00NE3ElbuRJarjXjwP/OyIK7Pi81Qz+CiJUUbX71drxE0X
K2DXcY+zYsA6BMMNXVXS3ZYzd3rHd6fjHQ2bpSgNauHZr8bp1ylxTkliD6srcKhV
Pccq1GN0PnNLlGXYJ+MyrhLlp6LJXfEsEaasEe43xFuC80ehJwwtaZP+HVadPJqL
Dif3TBdbSXcnOSnEWZKl4ibDJdPeCEZVxO1DIboHTTj0yEQqIILkE6mgDfYfDvKl
N4Dphuj4TyobFSewGYHGnSkwCePOpRe3eJ2+B9Zxhhv6y3N/rGUVMrodGtTnRSAC
dWjuzlnIHUpZh4+hGAKKmGu8Y/apk7wMdVuhKO0cWh5aRywKq5vFU1d35HTzg8XG
O/DP6RXZF03VBzghC9NpxXmHIHdLF2ACWXmw3zSsoNYsSEQcjeTx2lE3TDaQOKfx
wE9bHPNYaOxFFe6S/32TCgA0lF/EnhdCUb8bKtAY82nr1TMwp6pupHVAxPnwqcAc
rRwPY6x1N+H1kgE6DLDOm0U+giSz00mxSM8o8JCckwKNTNJdLE3mk++9nxB5eyhR
MJ/gHiXdjy4tyKuzfvDhceOENzpNU6RgfuPEuvdIU6ejsP1MFAs0ObOc/4863jVR
toqvlSNgp0SB16m0C+PRezY9LOpWqyVRXAJz99daq2sT9LgQ3/CjcpWjVwxQZjfh
EuSFFyfGa2dRyui43EZtdl5TcGNUPMwgTXSPTtzsoQgWmbuXibnYEn7DXpwvKfXT
kzoL+1kAEL7yqF7sFpdsmifhOle9oDvS64V/bfsC3lCe0IaJplNmagktL4UUKV/7
PQeLvIP9jTuKClSt1j9VnZf/0i3dNU/ibEd2aD0282VOb3frrubA9QgpAeqdQbab
+4I/OaJt5/DyLk2zAwk5E7y4bcZpplOgt70/zy8M1gALj62C7NbMcRlfEcCrnewP
/6SANOEn/2dsQf6PWsQhY6M0IJQVgOfE99OMpEM/EZPLsnXjsCbdv9WNdp15Z/Bo
S/nSv/u+vkK5sDfSsTC2c5sSNN43fsxiaPlAhMkOwiJhQMj8vnYD2LXQJq5qyr/P
KGcLx5/rypVFazZTCh8mDoTki0jJatT1gm+6OBzOXHOfOxesv07IR+rj00fNEcfz
/GcNukh251xRXlK+DIpkCOkoAPv2LauHbRxC1T/DjFlwT+eQpQljuy+uIF5ioDgr
Rbr72NFDJE6y5XhJqtK7Fs2rRUCA+AjPGoJs6a6K9KaN+WVAR/crnOXXy5pOc6jR
+NCtdeFbw9us+N2wCrj4KsWuJn+Xzm4cAUQeVVxMUW+3fYQe6gG+M5mwG9z+Cn8h
zHmWAqBghRTMp8QsvtEhZA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SRWX3SDJI8w7yYiMvozOzuilhYc+tdiKqq+3qQEsLLu4egUEKFjwmX52WunWz89j
YVvEC1WHRx/sYcqnnNMVUKej+Cu0KK+y+M0qDzoh1MbXP3cCdHa3qu0dKseZWEZ2
yXJDrrZMclMj93tKeyr8cVkK7ZmJAy25Ifng1P89G2AnRS2bOrx22AYgnOn/z01L
KwBkY2CyY6s09Wxhi7iWlEOpnXSJYtP9t7Mdg107JmxJTWJURvi9dwF8G36PNx09
MNbU53t/wnFaHxS4mB53QoCISfE7uvUiEV1LWLDu/gLOOO+52fa2LzHs1JSP3g49
XiNDuN6NUaLlWQH5tJf9cg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2624 )
`pragma protect data_block
G9NbiShMdEqG+up+yFYlUfDRPSNfWdrjg0wzjCQ5JIa0urqJwdhqt69ftUT1iBUe
UNsaP0j2pY7G0CjWpXWfcUrAulRjTYCUe952eyn/JpC+Nb4XMc9PxibC9fb2spQ+
b9g31TY9eO8dz78pENxq761Mqf7IUlxtwCCShvXFQsyYaORm9jrtVpWzm7kXKLhB
acACuE66iDJ46zGzD2O1OyS4PQEKbFFSvVnQcGpu+Ryx3I1Wjuv3HvWJi/H2oMIJ
zrQCPvvoc84p1milZtoSaAZ4lED5xKaG1rGNHLE7brxKZ1ksjhd67AiQge0Ix3Qn
qbOUoSV0XmWgWaCtB1+yo5jrP43Ktu5fWdwSjfjXJ6wmo01pTNjOTL2YGkrQr6IW
qxNUTSualB6c2Zptci9nonC3ZoFA6FPVeKKVLEawxfJ8ec3p55QQ2Wrp2NDpdSfS
YLCGUnaSMKoC2Xw7JDhfAxghi0/v19An5QyNoOZ8FpyrBWeTtlDOtjFRyl1SbCGk
3fttRP8dO5HsXBwt94b2g1kSmWF2PJVGENdE5TsuxTo3zdcGuCA6OXvVSteUwqqm
pO7SUFU5NuO6PpOkLSHA04UydwiIZYjSk60NC5lKNksxb34FDiksBSipDLJjeUvn
RrRUOcrTTOOa4NXw1WV61CiJgM5aSkDkQ2i+hR/nVh2yql/t7vw1B0X1XTjbfPjA
n/pU3RfJSh42VmJu9eM/dbUTaoNi6cU8u6wZw/f6hZjm4ioIVPKwPFKq4RkquZHD
h6bogC9bGd2JlLVmY0sviv73puCrQm9NuTWu+rxpj/WhKY75tUCqHGuIMr/3U8L3
fGJw5S6e+7MeJh8t90lnigKlXtJKddKDKCJkOXmXp75UW+H/h/G869+wuP/eMh3y
Nag085VQsDze1/Z+yBlmloLaqcownr4zNAQN6T9pvnnB9xfQy8vKsbhbrMhP4oLn
DYMUh/idfg4W9r3tZfyQebUTy+ukG0wNoq8dr0Y2Ml/PPfQiUl/Lh5kFkBDWw8LZ
q/AWOmhV2DPxK+W7uIRYgG/C8oKyUd1Tnuz2wVYmw8OJM1enuz3SUs/zSh2omACZ
xVtXNjuH+1F+RqiAWw2pY19aSeSYt7q60ZYIydSCAjDjrV59aPj2qXs6mzbIDmha
YgIH+rTp0Xeqmi+eb8/P5+PrPrYhzcEY7lRb+dBIdj0ntkjheclnNJAFKsSpJVPm
wq3hTG0yVfjsI6VmhaxJ55X4/vdUjUzX+9G/8Cwdq5C1tQmh4ZEJqU3u+emhhC64
cLvEbrsCb1vlc/sDysbril4Ip92PB/JQLmslCsk24nmQ3vwFjoKbdc8gguFKlhOm
1YpforQm3rYGX+ZA6986unl3Aec6cCV2bdcAAWP/qew8jnWCy7W6RmbdkBZRn/Yc
SKE1Nyqzs/frdGVI5jFOHKcpW3rBI4OCbSHsTDu9M1dptYN3t1kCHqUpgXiOLXwv
2u3vQsWU7rhU7AOyM9AjfjLnhCSPxYK30lPq31HyQ839LTFYXW/itXDOoV8947Jj
Ol9nqfoCmH3nPbe0v5aXuw72GnyUb1E+DpbBwpxJch58dTXf2xB3+qGu5PfV9UfT
eC+6flMlzr0IWfDkLF8ooNzbURusxaGbv79lTs8GwycCG2zWPAEiv0/FjIfMUUIE
qA5uCRi+qeJXJjxvGJFdM8e3m98NybKPqtOLXGr7dT8+dnokHtqIVDb2tYZ2+HFE
MgEmvA65UbFY2L9mEugKrxxNYngV+00oCsQqenhpyomnQPrNM60cHzykLjcHT31d
wlzIMbNIPK3c9lnaFShePNLfRDCIcJFiZMG64VIhgEsUWkMZJhvyeRIdZz8p22mD
CTNNoZIEj0yDfJ/VhxR/T7qvViyjcGCbD00/6zfTAbl9GTp1nP7WKATyLZx6ITV3
VFxnioUaVjc+b7wRev4dfU7FGF6Eb5L9ykUSvmqeQK3/G+Ic4o2O47BXpw4E/sns
WzxTcpMC2qm67h3Ue8JZn1xk+Byi0ADjqex+bcla8Fswx2sQfivXnRCr+/E5VBQL
CB4QNHyBE2klAfyaO1niPX2NwBUMK6S7AlpEUweoNs2lGwMFymj+QwM5O/T/icfv
cKQGrNzD+EXLv76uNNTtwlxKgFy6sPHHoYMv9ZH6MYRvXZL2qW1pwPI44WGPxsu9
mm/4joDVQt2TimoY7IU3glRhn6avhwXRYqtSjQB6XzVXjxhLFzGRSofLXCGUQPdr
JyX1Ghlx9Ab6lsDFZ0UY/bvyv40GnA6AtFxzDuprJLnHpY6dX5QpFr8cHEwj3gBs
e1vBSqNMwGPUsWI2mqvXKfMaqT5fTDaipBZ107l+rpHsiYWbHnwl4gfDwVCiGe+C
2PVCjzMriUbqcUZ5CBs3Woih68OHtHh0Lhkz6JypMxKqZrM+YM+a/pzyIFsjoGbB
jaFh4dydO+SFKmTGEY0I00AEmDIfH3XpG5j3L+5brzwkGkOWXaXfopbKssCi9b/y
4LaUXGQexqIF+w9+ajzUvT6Mccu3C0px55xgOvQ/gr+og7GAZ2ttxs074rpAcUhW
D1Q5zGQm8E9AVL6bCStOhU4rORYm60wgA8D4NzLf7tvjg0UQCKxEz5KRr3orwQVn
Bx8GEIpccWqDowebcFWblBbcrvE5qHU4xwHdiOSEYv5u1M9NExKvPW5tszi67ge2
p2aKAOf1KqxysduspKKC7ZOEcuJx/tnTRY/3li13Lyk9/pjKndG2hIxpFGjVhF6j
sk7E4UAnPBmUGUpiq5AcN0M8023eonfQahoV0yBsz+1gtsuyXwwBALhjh6N1+Dd/
LZUMy+9gkidJENlxL5ZdjPfvhuR1FpOFNpn+6AfkUWOapRGkbyRht2BbH+55An7D
wUcokrMN611ehKoTvvwrgcksMbRc/Y/Ui63CfFgJ5ljHoaztWirTO9IGYrisbSES
3w5iz+J1jtflP2MljG2Mad+YAikaQVy9oxpcH1hpmzQFtnpuCvwbwICAfavYR2GZ
yfEY01erP9A9kZUxeTvN+iO8twONyjrLqKb08Nmlhn/rGOKcrK0GJ96juIHy5snx
yNR2tQyhbSC4FcmLZJoWKVGwU2m/oRRyAbZ0g73S8IZj0NJKN9MEgxvBeOUiMUUP
qrj/S6fYsvT1I9P6xYNlgNRc+1OyARZ7eRQp3Lgkix3JUiYfpG0FgjHVW3dipX78
zPojUrBAFGXDSfvnxMOQns94/wX/WfZL/OYKlH3MF8CdUwiaINeig+YeEwU81ASi
FycgXbBXXroU7UQsO//MQXPPQ8CjzM+nVIA5pETYct+VB/QTbhZkRKa4A+g3Agvk
FVpepKy7ZnDZjAJUvQJCA46Bc+/GBCHDbDsz3wzp761r/N4qE/d2iK+xcVK2i006
WbB5/vK3LR/6PrjuNdj3DvaF3ZWdlHQ3VMqy1BojL5/HIzK9+gHjjlsfflSxbTVu
Td/0isQn6YfHTEWBB0rbW+IG56ucO3+akLfD6yTQlYE=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ndahK3qRILVNEkdCG9VkvdxTLGP+QkPnJz64IrOVGHLgSDzyVTloY+CwFWhLYnCw
Z/PWozCeB3/fWtYXCQscQZZiC0VnOq0Ih6pb7se7puMVYPw08T/ZkcQnCIEroKkQ
PIQdTWT8B8f6u85+P1ungkbu76IengGl6gRq/NTnAMotOfdgnGej5KDXVSvLLbsx
Yw0ObIE732kfXY2ymjJUg5YpwrvFgA7frw8b3n/hOinBaIEUqOKgkLXDtVhX9U48
iTpALp/FlJoCpbh5rYf2BgW1ml6PLnWeENxVgWL3XBTxiryC1XvQ4b4afbMxiToF
oMs/AkrMYg5+a/HPXVpRfw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17824 )
`pragma protect data_block
wA3y54enEqydZgQPNfvPu0LssskEMHAJLU2LbvKYVwZTJTRSEZ6h17VfkopXKcjZ
JGpRS8C7eAtnRg9WAiVWgfFUseJUhUNR2ASLLvbYS9yMa1R9Wu5+BJk/wY7iGK6/
Oq2b2el9q2ZDREO40ueYfKYjRUkbrHNaMLfaDGngAquLmf7Kkj7fbFKg4XCZoKbC
Jpi0MhOVto/yW4MdK+U+qct1LcKAA6y215qN6a0NKqvhZICqMPW/Y1/ZVQK7+d8i
4gunsIW2l+I4dHLEXEW/bOxL/YBEYkFRNjYwzy3B3fUL2/gpoLWqUMESkK2EgTyj
4btjcqTL9E99MKzJqVFqKCL80n4bBwlGPTNR53ZSbhImkN4yGMdFf4Sh8Cr9Dni7
xuXXDAlCB/2VZljhFePoxAOaipTMRKz7KtEDSo3igd2wnm3VuPCqDPSxxE9AUWa9
zVv+Zjk1CmkrfF7JA93H0TLgO1sORrjJFLDJaQHfEl4e9YK1YnAfwlEqtE0Z23ve
QGnQgSrUkOOo5itm7nhXqgqgNfDZj7sptiRtm6L12BTtbWmvrJbGXv0XK9fpuH0i
RdwNY8yw/i/v19K6w1x007eWAboACK54vJDX+XNaBIju+1iScgvY+XEOzDf0BLbx
yT1AWiUg7J38M1TnVuJLQFBlp0bCTg56Kim5n56ZKfgZk733oBzQQBzJMPtht58c
pgNLyMLHFD3dhx92X89ZXymW4GurR+UuFph9Wju08rNixE66Z3yDBm0OfCkXMgdM
vvjSPMvtioH0U7EdPKgzwf7bIi0mV9FXA9Sz/+2voTUuxbX0aidIAeczs4LcXrfP
bBewTSjBrlKZp6E7t84h3LW3imjfzU/GFPXd7POFtloQGMr23k11AtSWxwIVjxP+
ouowOC7HlzQ9OqkcLH9qYgvPi1x4R3UnW2/f8uwO4LsEAfU1NBd45e94ufBMBX7V
cDOpxILg74mNHLvPp6El0RNATZ1ww5sOis3QkKrRLRv+t0CvSHNZkkujx/ztrglh
G+DnhNeGvHAa2x/wGggCiXpI6D66dgVlFOkkE3ybGEumYiXAu30iLDEX4iT7nH9f
DdFaYgU5+pHbaJttMbF5FI3Hv5GpNcgzWE8XFp76+d5A9IW5Cl+3xzUh/F495v8h
EEXwRDGlCleA7TobkoyIRwFfxPWRElJxNwSTBfWzsy38fGb5cxzyJ1/+mTHe/Or+
FaB2pLM3UD2R8aWkWBcgORQ6qGIAxsDHzCLP0Cu/jovAb3DYiwbjL5d7hhXLOA4n
vEpUk6yVZV2VFuDf5S6pKA+sRdLNU4Cly0MkI6hBKVVtG0jvtYrUJjWeTfIiZLop
2bR9TLUISHot9magVLzDk6lboLz6X5huuQq/l3a2U8Xc04dQl/8lFisnTBI2PqWL
Hch2EzNqlXYNcdbhtVe2HyiOy2iAzxPsIjBEKQ59sifWGndDT9rmwosZgNl8K7NF
FEPmE+Bw3wlvxW1inMZLLLMesc/DPtOq/FjJ13W+v1MFa6RR8vYm4LNJJGQOkoWj
HGSSjH2m7j0nNGIx2wK4kFCBWUdErR4ASnu2WdsDr3zuJZOZb8w/DdxFDCVzYDYu
cVfLihkATQSyzFf3icWz1jeW90JOLqNvBQ/Nf2CaQ40AISvZWBHrspVs2NQHOJct
7drcsmVgiJ0Q5nh4HR1K3wYh07wjqBRobgygBbeRHKeL/5KY4oe3xBoA5OU0Ktvt
dgWNzwKVZb3x1v8x7srj+2C7zmXhLTWKDfS+u5vjGVkWHgyM1lLHq2aTZf4a2iSv
0XwOWwv+O6u0kNXAa6qwu0pVPmYNNRAD1UVyz2HiPYYw6r3ZZOMl1qdUR9KA8Tl4
Boa0er4sx/JZSP6hoUFXsbrEMVGCytjxbig+VP0IXCSNY9J78V+FfeDm9WNE5F7t
t9VHiiLX7wso7YyMNPT+6j/zDwmN2oAsykwgSfHCAtnvjYpQ2IWW4I/X0mHbSvty
pysQx1rtSId5oMFvcnWcoIW38GCM1RNP35383ed4FgEtcs3OYSDV07B0qdH8R4e0
t7p8Qqanbx66aEceAGMBSV+biE1DafaWuVtKccJSs8x8+el5bhmRF3WTU8AOug0c
7ubLPpiHlQU4dgHR79slnjkIzNek2eaZ3dWRY0D7x5Me611DHWCiV5Ypv8MrSoBj
QsLp2SwBOjHPjsWeHL1GDAVzcJBTKojeZ61io+rnP4K5C2LVWb2Jyxk/LHbwq2Dr
Q8AxvlrqrkQvfLrBZkTuSy1+YLBQdZJV6/qcv/r02Of7jYT53FzCjT6PVG8WGBdW
vU8n1TirWhVoECofa9LAuVcXVVHMdPn1Bc9mMJtmms05CJ89I4sTIJoCHR5GzTIR
uLWH/9H3XFijAdzGEOCaRPQN6IfpF/2VG+WBCrC6iediOVzdInBj4t+yH774Wn7d
3NI+BDHyq0TO5nxJZ95Z3DkN7Sty9cbKk/6Rd6F9PX36J0MA0UlsQAkVoms747AA
mgPyh0Z8AtMYw4KkhbyriTCZSHpfJy/8CiI1vqPkfUbgXL5HLi940Y7k0yr644EX
G3wRD6YfvVgS4sd0XdhqF5+b7oUR0xrhUy7sW241zCgaaUIKrod7b3iTHV0g5sfK
0Of6rw0PqFdjHa33rsykWNXA4Ek12BhvmU6fmsINLYrIjgcTAJZIdK/FJn/YZmD4
U2CzojIQZiDzecuWXHj9KpKZ10B6QCbZtrvCZKlH58gC95vfBXo2rvpZZZEMOvOX
NsvjjsN09Oi8ykEJH4ykoWVazmb2XM4TG9+Tk0YQCZtPctIWm2bMHLBh90tmr6V2
MYrSTxUNkO74EW5WS+X5e5vR/iueUOMf0SdLTv3Xv9BeFQZY7wTm9VvcOSPm/hIr
IRWC2eTaN/etihn9ubKamyyTcKUr0SwuH1RwsH3RzLrSoXYkCPZ3vDGZ25EIB+GJ
n8lsKbwnDlS7Y6BG4IzGKrMrN1arupN0e0tR/uFWZug6ISh24iQLMXxa55Puv3t7
QYbawSoAjwIrztPI5ktjn3SwsIuMJCfP98pRf1p2d9+ZbMCKh6JRo31HUwYSCGgt
sFnbDX+HE1wy3GFAJc1xGDpzry2ZhQRDID4D1IJdXadq4ouFL8w50Kq6CfhmpYk+
Lvx43udsHmJeGFnZe/FZyrdnz2ZMA2lIf8/e94y5GD/wRaPbA5YTALkBb0pAh/Lm
waKtBYqnQ2yPlAwynCSZPcHSyOU/DcEfnqHC8XsVfGpHSQtB2O1NEF9fO2U5j54A
JrXY3qqy1W5+yB7xwgr+Bn1OvOOAgup0Sy2Pv6CFG5xIHQyn70NejPLzMBwRYj8V
9wp6iItFJ9Tz+vLgIGh3Wl5v2EXXfI6TvLNiZWvOfnawX9JGPk9twzDU7mCXxngh
PRcVXIBR0aw1SPTWV17iB2X0WEJYCsvw6yPrMBbJ29/EL6bzbBYMU39NZXy5BMcA
dpSilaG/a2jubhWX+qBU62U5WJqO/yytdsD4LUj8Xu7QcumuApMi/fNC17oc71bg
jWW3hGrF6ukEPBi1xuwA0KvaH4GFqWVA6aJAAjnNRD4duR7MDMo9+nHHStF9KG57
SZTWL8y8+evn26fgQqWSucoq135tDUVoP6QFG2D2FHXBOzFz4dmR+FINoaS3MOEu
lySBywGegBIom3P0PX7aDI8sYTrMpUmduIAQiCTBOTe8Q4m90DhmimTx9rRuMsZ5
os7/+5UgxyAcyZfbgWueE0eHxIrpY00zwMk5zM1uuLdUvcqVYQuuPdjf8NyPmjLC
rSfdok5BI/sMoRIz+Hu7aL6bepkcyQLAro/PrJ3/QEA1jGQpFbXfUYc6asca3Dsm
+HqbMNwJTy86I7Xl5Xxbc3bioqJDNduvb3idpiQceQiC620XfLE/neObNB/ySIHn
+/x1oNcLQVTTMHuipgwnC6USaalIk51RablLtbsh+Tld9wVNOCLPqdvhM8FME3Yn
b/lN4z7+kpwrrWsG4qCZxtxfOlBdsFWuk7y1jrSuwlpCPlo9zFXzAWsrPzE5Mtwy
boY9wdr6KQThidvVrGOM8vTF3MeC2dzS2+u0z6zX1u/6r9w/VzKXbdp/IryWIOZC
gHreKvaow0abvNJV39OGxq0uPj2ubeXyuuKP/i+Ix5b6gtPwgeKINWZonewtQJ7O
T2FP1aetJ0EJel7KQVLGp7b0Gn4wK0LA+1gP/EOio8k5z+XDSZjCm+GhmwT8TjsP
c92Sgc+O+a5oFcN/nCXWA8rdYEPhSvfIn/RR+ODjAEh5LIYb0c+t5ht/X1gSLZ2c
6gKSYw0WVIqx75oNElYD3DePW8zXlgH58GX6H4dFnQ+aOfSJAgU9ybvok0ooSK1X
IBXCE7RaYWx3pRRohTg1Gn7NGXo/XL4YCMibKjlrPNjtEiR0v54qG8zMvVcB5gx/
Uc4+8INQaGlYE29lN9l+9lbmLmZnZK7b4zvMI6ydSOgglXTdXSdn/1/s1aEYBsQz
povaMieQI+XUneefivJEXK30sq65PPbpwcHZ+8UrCJ6vKFdU84cypDKnlM4/ysQc
XSYghiIIeCKgLQk6QR0yWfXsh3OwOABkE7sE1+Xp8pMo2MnnSpbE4KRvcrj9dseb
ZLoAzKq/1RlUf49nZBBkaAn0dzhe4Lg/zH11kPeEaZWiL7DhIPkDvknfwzWov+kt
oOY00nyZEx105l53z92UZg7hw/HEO+7u1HDD/egfbmYPLitdzrlvzgyqzgDDuH/R
DAQCdFF5+Qzi8yFNsQO3xe9Ts9IvsTEL0WyvDk3sXsAYhSaadks2BQIH2MG0FUoD
vsVHWSJRhnfzNYtE/iD9NHgBN+I2zHl5WcuNTv3BcR0VhlV+AOiSqyDJcEsLRf7j
/7SapAZcgmSyj4DsadFUw1sPDdkqwRsgcRG9QXXM2ViUwPJ9NhWTvCQI7mE7ruqa
Yma84QG2OPOIlLt6Rm/UdSLmkmEeL3BIJ/ylzLLUsC6cJ5pVjO0oCftms5yPhgis
QNW7d3ij2IsHVewapycseXzvTPwukBpi9N7H8Yyy4HOMVX4s9C1hwkCP/u8oynhq
7pGtRf6u9+jLrLrLbnwHm5bB97Wvo58vGzrzZ0kFd0De2sbs+02eg6lF6N+9kYB9
2c9sJUFXQxAGH5a8ErH7RlG78UxEmfYNFAcVnpjlOunPKFlkYje6R3h2ryf0ZtTM
7qSF987zkcxcTZd8SPfAObc0g1Xuk3i4SnHDn6RbQLSVj46f7u++MMZxQiGE1sc0
2i6wsaGcDZXXDpzA76XJ//6Jm40zFoYi/VkUWG7fxWiCcs5Yqs8063YjNkZGFDek
L++MU4HOIWN+Gn+6JwlHKpHxliGZRuYgnZw8urK44OBzAk2ZJhIi8Yxf/MpDPZ0A
VLXfIdwkrgUi9ywc3BuTZ4AC+AsZNrm/WWPtoUSTQy02Qgn6bM0B+SD1pTaWkES4
fUDf1fJzwBBzg2ubqVamtIWub6TtclzRzTXiwDt2myADqiuOYCPiF8czduxSgXiv
7ucToOYcUMdkf6aVzXhBGMpLkdALn9pW2j0sLm1OtTt1AMogVjyqDo4S++sAyaY9
D5bbtIDzplzejKuUjqYKRa/B8U6RSLhz5bFEwF+GwP9iHVjJMGNbSxxPfgByub5B
obNM+Ti8IYSFgWi9rAKr6vse8GJkYFO9yaw9G6quT/mc4ANTBXSucTz+FfHYAwKD
c2YEo/8tFyTNW0Qp2B/tHlO5QXXuVNNHrzvYjFUkMBWmXlNpbjD1iRmVy8BfASuF
jt1LYlaiLGEb6fLpU+FaN92Sf09k1u9x/UpJMAYCTpAL2W5wUgx4KyqpECFltL8G
B2X+ZZXvknv2pvmJR6NxHpNayaddSxbaf/jQztSiX2dcR9AWd+eNY45MEtG7AW4s
eyzkEe4pCKTJSne4XSuH8volPhMnXGQvPsZAi4TEkEKzezf3+eeA3PdZaGK9oJWO
k+3P2mDPEnhH2o3u5iiz94SGq3OBYfZDeaTOC2lbsQu9u8QyssJz+rtZipc2PKfz
eWWWYPLxbY0z4xDmfSJ2lP4/InrHwBQvhJuziSvAc+hTJN5xrlj/7DFYP8BSVhya
kG/x7KZFifWQJ7THBNpm3rvxTA/4pNB+eYtoyF0h/IjhouDtt1nS2UUb1d+p6FKV
06zRkuD2ke13Na8WKLqGQ2HuJhes7hhAoJdz6U3AvnWtJHjQuiujb3+aGwVLAZLt
Aw4XH2y+vtdQIO78eNsTXuJJjB4O34sIVA3qIn5WJWJBu4zRHhrnrRnCMWjyyfi8
cRGoTL5/3HiGS3a8Pta2MPLAae8VNyGCm1ECCij7RQf9D6V8gq6rrXcIXukIW8lQ
5aj2KieKrAzkRBVDbdjHCvmTRMnUMiYDXqL598RAXcMXP2XadrIUXzCGu2DGfw54
qZ1Ze5wSGmfg9G9sJQ4kpfo2n6FiCrewcvA9bCVhchg+MVYD6pyprjc67y7w/P9N
oY21bh8Xc79FUwJJg696nM1lxFAyVSX7OSDFafjycJdzgXsgPgyXzGQ8ODmklntG
+5AEjnutWOGVE+YFAlA5Ro6rOF3zUMuhulSSE5lP7QzrCWG4k/O/0aBX8sqov74Z
xKv310hA/p3P/HGPa9RtE6v8+cYDrCh2PF8P762/OoGDUnioqNJd7YuUFiesWGLY
qkqz287rP6/y28Cwgw8RAJA+ZGEwmHPDoQJqFIzeU0MW8FTz2AKDG9gicAWqb+iA
0pQqTqh8utLvUyH1YENonlOBRIJ0aYuUhdxAey9vY2LHH9QCN59nLWD/alH8seLA
Cyl1E4sAsajMuFQJ3725SEpEt6JeHtZBHfV+H4/AY0K3n4b3rvvsKKhzuLxXI2w8
+mlXj8hvBhmyXp2plop4uLiJ+B0NYGQy5o8JZ9I+vXrxEBkK9PI3qNqJufdcuyNU
NNKzaPtrkDuPvBEn0coPLYXUPzGSLcVmHPABjJgKdjMRrfaSIj4Dfhfm94IICkr1
w4FKWNbVTpE5qKnarQxzBOpWlUTn1If4K2ZfX1WW2mYqrqGQP1wKy+61hdRH/Vcv
JU99GOh0ZxeJf8PcLpl6QwqyhFcUz4cLqwQrSd8E7GX2OB3qnt9IeCU7Heys1pNi
pRTFKJ2cHb4xdUtAXJTKturle2Gp4naC/J/hi2W64pdYIURsdGvrnhP285Hw3T04
ydzuEK+WBBvSinxZme1BxlMk21EaB8S77an/uKDn4DNMbDV5d5W6dJSjC5BxpSGk
C63rkDt4zePEVAHY+Ujj6sU8ySZYw8qeU/CJL0dwqPlxi8bz7a5fJ+Df6GT7sDYb
+z/IufgUaLms0xZqjq2BzKr2RkuNKy9nJCCdgKh4Xf9aIZebS+kvHshQD/danhES
gi99Nn/wcrsweZfXZloj349qQyzoTkpSd23z+wYEUzPw6Y7AhmJCKSPtWP610993
YNnIgusFrB6cr8zYwEYlCIV978d99c5n/Eiexj7o5WjlsalbxirgfLvoqYrtoCA8
pv4rdOSdGq6ZvxSF6jQAnUe2FPtL4qtp3A2ZwNaV7ib5jFNEgLzWXbJEC2nVZqMU
btJygeyD161qJ+3tGOMw54FqPoI/VzSiTzEdTltFY4ppwdNWVWbTv50GANwlTlAF
W3vXJUHNTtGm8UEiLdnqlcRJeYB/nweb6xvHEEHFpvzfE7qoLAKMc4IaRBuFsnM6
ZVEL3QmuniOyO1kcZdj4GHsfeOU+cADcWXKkJ/yXpD5+mQ23TrLMIhNuWWV1sgTi
wVFiqHMTVKnRz+y+04I0jhM+oOhP5LiN+Im+hgJJomnUAdAGvJW4G4EXjsF6/qtb
jc7hHhEh0EBffTeHFY8YsJkm0zQGjJBqZgSvngUUN6XSIi7Nn/63isQLGsqbD2E/
D2yZfb/YuRb8i9jFTbKbLPMsaoLdOExCBWeir06fi1VLBpvaoaa/AX2+t3sK+Tcg
udyhj73HvEdWnFlzodAgCWsDmP2GpDqrZlqWtCXZev/g0j4ErwkQzgTU6yJvNFl1
Ox5dsvAqTypIPfQ0f4H0Lf2tRLDYsJOh3s3incMO/3wuzjCFMt7Byql+lePC/i0U
teHxHn9IEKeTWw0JpRiZPyP0pZqP2hy6z9t0ZY44pMm4pkKPukzH96EdzgCsjTYw
61Re1/hTrSMRlLExj8m5yIUEKoqY+ELZUg92gW/M9g+GJZQ1OWIUlZBXf87lO6M/
kMN1dSgYrJvtx4JCQWWzjAwhUj7+RT7+LAeeJG9uQKnkHP/BRMaJ7mHnuAWn5PRZ
DYFHGbVIXy76JVuXJnUzNZuJxLlecyEEKqkfa+4UskJjXUv8xp/IWlYQGnyv8Z2y
M5Z8haWU6qLMZL5R/6AXoUzJwYzB5CMvN2uFT3YZLlR38b2vl1M6z6YL2KQKE6Qx
77tYAniKoi+9FKOlHA3O7J7ZeYek7R5I9Sus8h0U4AHmjAq1WfDcqKBnb/KUKmVq
imMP9C4BnDdQcYJbFRwUwqMaJ4pQUAaqO+5VRw0UlLr/Aa7iFdJzGpSdsF/WUZIl
ClzY/xVUMxUAcnhCx13yhXP0aVGR4ALkDysN2ZZ/ZTUHHwNUv/m5/L4PrOpCWtAd
5a1h2JPHczeo5/C049i0Dkg6nOdrEXZsnk+cJJ7lFted+P0wqicaLX1Ou0u/VnMT
DaEMeSgUW7iWi+hPiwm72M8yX3eck338eP0/HfJ0U3rcGK0x/Zo6Xf5tbhkFqoba
EnL6ZKmP+qas8Cbhp6m0CGELfOfSgmO6f3n6aqgTlSORnia1JQtC7c2bZYnvIe55
IRmIzAGOE9djgbbTUDnqOSFgnjFF2pE4LBrWWtJL4cKlgUW5Pn7Eeafkw5rngQyS
w+Z7QMLNFct0L31rL/ydWNR7o1QoFqOOhRhdUrhJfnrkm7DLjMGo/Gmj6bb2lIFw
ra6X/dVtVqnaVucM4ZxBgC/ChTpbw+WxizPkUlrTfsacuhsbyXTDtNgPU7K/mDkf
QeF90gGs9CoUUOYZg5IwA7JH4fbH7lTuJZwEgZuGeIHG5g1SO9+N40tL5KCyGkYc
O4dzGE3TEiVcbdpa9RUcgDYO7CvBZ90JrkchKLgobqL9lhbhpNRNQuhTT1pKTYFk
7BgMJjbc4g0+ZBVMAx2JUQFuum9vrgaizv+1YxXjsSREJhr8iCNZVlYpLsfxqBe+
RvpK7zkh3KwLMSlBGn7wI0bUC02GFmMiTp3HY7TulicCDhW7Sg20dEwEbdB5WDWl
EEPreeDqrcMEomDwXiJDsTz5LKKuF4WOZGAC7Q9dZVa9XexaHe9tFhobiBrnRLrf
mVrwIkBSl5yUyy3sOq8Gd19NBUnnywXCgY1cY/NLUCCgMLFs+kYhgnZ4OoPI1Cau
3s5+loLhYUtOc5uPi46BIatZFmBIuoZJKzkqueZI3pN3QHUtI2WQ5nq/Qqa8uPJi
bG7lahrLGCtwWizdQj1Z2XgstcVjGOdE0YOxTgDaSb0g5v/NcwtoDOvuZsybCT+k
5l4/Dq8z+2aGPtE9zrlsCZQFeUn+9hBoFoDIqH/TtNoCDwuvosw67Ia9wgurglmv
jSJI+RwKq4i9mWb/tMVYw/UzMPZ1BWKIrSHTBV7Visai6LdnAqp8fwBB5CQFeSCI
mgnSE9d1fBwRbgBF8QAMBMTjwBHyK21qwq29Ay7xHw7r2NxBZBTx4BLM6FcAp9V4
8+yGJkyEQmCI4VH+FHMQQ8SkDqB5lw1TLryiutJBwPnCWzDuQTbSQtXI80x6J4cv
j9tmg/BwnWW+XRGUucGL2L8bkDzXfpsjJji8pRUaMZPrNB+TzWtG9Yps2FfssYMS
ZqjOILecPxaW3TxkT+oUo/GI4L/rLXzVIUcKLHcuuLCYz8xpf0kFv1X1S7GHUp9z
1G6mJ3qHMHvXDfVEVmyrzdASIy+Ju9F+O+klX32VbrEo+XAnkls+CXQ1/enXckP4
oSiuqZgf5v2fyZOQe3xvBmI4pfa25TMtmFSAgGYJBoUO5M2ePFfhSyajmUWAH8RG
c4rVbnEceiVL+c6QSZaus5PvcecptR3spo23WWyiFokXetdqTRrkZkSf+ABMWyDQ
a+jSLDUKOT4uSYP3oNGrJx3lC5mL31Q3zwvVsCg+5LeP0TO4fDTgvHqGFcwyli4s
jdtJjYxrlyIJv0K0a/+n+lfPqzBHwcZY8IHAQQpHnn5SglqrmaBAtbJ/Efp/2feK
J8WR9PFbgjHnpQVH4ZjXtzecaIecWRWxAiopKc63myf3PmfqG3XIloGlbeQvk12L
xl+1V7M48YdETJEQgp8aQ/etnyJd+38SjTPxkIwxIY7/hUqWcBYQVcLXnNJqtI8h
QKbsEINPS9Mhvvol78CySPiUNtxh+asOZMrTWq4s3bi8C6pXY8gWa1rzTHch/x/L
3ggyZPVXtP1jAEszYFwICKCHRQRvbd4AQLim8Amui5VE6/Ja7Th0eYT/6KdPYQyB
fqSFbWiBgQntzT5zfEIZB1+1FU0aVCKerP5orIdNLqzUvUhL1wpIxvpXnlPkdBCO
tK/AbXuTRnODVIR0bbSPKvo//JqE4nELaSLjJUtl8dyf0IkViniSc0PX5vzOUf0o
1ULdJX6Q8j31ucXWrt7vifYaxPISGN3TL//I6NMG6B304DRPrXeaRWuG1uQXTcoV
OjzFsWI6Hp2wpDTJwAeJM9qHv6GFpoKNZNHxpROcg9kQFplaC6nVQ/ZLBipgMW6i
3xYX7q30wGJjc/uxNA2mQq5quDB7gV1Dj/S68Dtf3UfVAHNbuhhz90mjGbISd8Gg
DTS7QNKxJFduc1eGwc021aiaRUXzSHY2g0Cncy68DWQyMS6OOdD9YOTe0S6kI2tq
CCYQqA2Gynae4hnNXnGTf71QIdrTzglx0QuvVfZeU8O5en3xQLS2xIiuVXWf+Yfv
3yAuJKWjnuFVE4dgJIQ782mmvJnMj6cGdOf50AtOGIrEqNvEIuoGWUEdPNlIVA+P
tSJ5fo/JRrKnRwpKZ2kw3wR0w0zsR1247KtQ5hayXbmj+mRmxv+pfmZBZKASxlbx
Gyyi1HBtBQd/mXuxO3kA732tkws1+Z1cxNOp2G3TXBE+veqtxzXapPw/5rPW2asP
sB+C4VqeYekGQx06MHTENt9fG1X4EAfdYQg8KOkXhgFv0uMtvawGZGSxbra39ah+
Q5G2STgBtn4h+HW1XAnJHfmHKT5Oxwb1daPH5kuZSSmi6X4WrasYMLLh+PTILJoZ
Y7YcRxCAbsUxljKLK1PMDHrKxpZ7FWaL9Lj3YRWo3pCGlQ5+l3cN67Ppd75hxu0P
lG4z1YVlC9tSYLQBxPaRwKJ+lCR5/O5XpIPLl/YZ2PQ1Y6b9N7FG58p0ClDBcK5h
4+rHEftXQO0989LBYVQpNSrObMdCpzPd9XGS+dzC/rkpqXxCLCLPUlFy1KpzsAgw
LZnbe+yWGQPXRwQWs0b/VlN4ZBB2g2hlKQVp0zHgXDAzmxEjoGqKREedi60CtwJ9
ztAtmS6Z7Bu1lt6ywd2XG3Ob8DLD4Tqys2l3BnUAIcBZygjy0nbmrFiM0iAuIlO6
x4CElY2YiFe2xVVFwUqCXd7QCsY/31DTChWFddLh1NmDcpr6odgAiajE48mg52ia
B6XAgOWXhIniNBa4H4KFcmtYkz4Bmmx/y4RNU0zLCwhlQltmtq0D8wg0taYj0Yzx
Vluyz7BseGN4dj+3gpZWfrKM7GGm1lEh/i2lM2Ma0t0obWCqzZPir864dU3U7Mkq
W/hzHL1pPv0uBdPQUZAF7fOuJ+qZhnEo2HY/QYnTi76Wq+ruR5UXHDOSJmtV9ivb
kgEG08L7XtUfJK4k9dYPbffUt/2HjxhSsOoa+zcDixttqtEc5PFxR9S+j/d8MGs1
yeR4Xtkih+ubhOp7QCt3YoYY15D6kT40woVLLaXsIdmcm89D8krO09nLtXSnXiJp
bypUfyxRyZm5AyuWdxLimFfutArMUkfQD8Xkwwl1W0OY8CADwlxvYaYrlvHXLPJP
hIvRi5KAJ1b/jHZ4hOZiYqY8QpPJ6jRKHU7WHUBnAAPnQnSMlkiwK99rCt7scJOL
jQvjwPtFZ12N7iO7wlMz797Br5NvpFMmYl38GqSvmzvYknEqPoHx7zdQvPcP8yOG
nPDSYwuaOCeq6q5W0Ts+YPovOjgmrdPsxqUMbv43EAqK2Q4mHyLwR3Hy5BA7eJb/
V8GXfmbA3LBCkIeNoNeWaVAJ3w5dwerBxTt8pakpdro4rJMojLEqCnzLcUxKB/Yu
lY6gBdxFtkLUkg/oqbUQt6WhYfTCh9+nqRhyFLLrXEEwPtNfKHLJHWC8y9qGHaNF
3hmj/ioj+rX8g9t7HMSpnPLpSfBzvr964AWVx318UZNZT2jyyEFNISInf4sFBHOG
Z3++g0AKsQYSbtRns3chfIyOqapF5wJI4fKZTV9uRRMvlMzqpBQHo2BwO6AldyzU
URbn/9kDSFNj4G80mkHMyR+UeLC7jnfYuEZuXfae+XM68v+M0QzVhJhcPX7C3Azr
RE5iCvOaDM0kIPwY8Rd3m8+nhoCDCw76EUXkdRQYDYk8u4Ezh+cbXnsDGtRlS9De
F0NukwMEIakN++H7MUIkuezM4IzR19vW4NhxJB4ICLKkwSDi1XkGGu4pwO9ewVdA
h0eZVxUAnq4YBVgFa3PPc0uw3fISjLFrB6Cn1MjMVGwh6QAiPjIXEQGvEKCNR69k
fHkqkMkJwkAqyeO4DcYvhHW9vwBTvbASeYyW7KU7mKTzZ/33jSJq5Ie31O+d7Xu6
UVwAoSpgS7zA3iNVI+rGR4TTnvcO8AX6iWdyIoZsNRzpH6Hs8NPfBmIxdmhWpSbB
DFqwF5MFI11mNZkGgzyRaHHl/xSId+QjPAr47Fjk9Wwpo/WI9azImLjdg5GYeDI+
zwaZ25JkUj5X+HZ2isfccbb2pn/JsT52aJBhUkLaacI1paKwdIk5RZLXngun5+y6
1/Adrsf7v4M3lz58vOfIuKmvfR/3nlxgXfgw57pPDSnzYi6K0lav9SipjoIKlTPv
01h2QTtUYj9h8AxQpH3g1sBK1k5IQPmo+POaIYa05EYIHcdoV9fQ4yk+D+802RQm
3Z24fxgn5FAPAp6AcO5xcFj2tx43wL22UfDjV2A9lmkzw9cSH6H47Hcs8v5rgqs6
dSp3zNIZQ+ef2krFEe767AvpCzfQXN2X5jZxQjVJvJOvnTG+b5BQ4CLYfKNiiQco
IySxBSRDF8SyCXLpXwfBlEfSq46nV+NVBxZ7oUfKy2C5MzhbSGZTLzDv6LudeC/R
2p1pcbwV1roaYk+TuUEx+3XKOMhUay9/WqNnb2NutLpDQHMwnP7YT4YDX9Mqc+T0
CeuZeYKcY/2SF+M42pXpUf5INPLaZXZZYjULLANRtSIyiMTfv/kH5RnQ+WcjfVO8
v86XgoAW+L1QdCdzQTE4jCbWsISQK4olhlImrqs4SAHqGPJ8JhPLe3XltzN80Iao
KMRG+PhubuAFbUfJVMuaaqf5C/5Ai7oyz/sM1w+2aZlEqb1CZQZEwbED7y7B/hDB
d2eTFAA86LjQNphrgf7Rq/P/WFIN8wC+05teS9WQ2ptiJPESB6nGKy9b+Nmp9OQr
6mV3mAhzknmvt1A+kInnYPJrl/4G+dY4p0DKZIz4f4IDG4ujrZYb2NwDYg3+q2wN
JBgU3BvnnQJVO91x0Vcwqj/PuCuf6VBAcw0Vaad1/rK/0PbDdn4WCfbwFpusOqZT
aoW6AzK20suM15XsHV8vI1+x3lJOh+oWqBpfjygfCZHk8qk9CAEG4XFJizrS/Jqy
md6gAvfuVyAZ1IKcIZKKSj0ukeInfhcGGuSSV9nY/B4zLG/khTlMRSvdcVhgMiJh
Lc0M87uEJdzePod9wYlVi2KWHNRn7HtIovCOWOzRw8uwJfFvfvPaZNEnr3sgmBpR
VEu2uftK3TqZa9nUjZipEo4Qt3jIfXDjlI57gnZrD9tFxvZ9TGZBrlBSWw5jl46z
uCoXry2TMW8jrTmAE7KqjuZQbNuWxT0kgYnEvZ0EeeTQw8XDGjvMV92mVt6oW6ZH
QqrjsJmStCFNmqzS8h7+XLcumtIUxrI3ND2qOg3xZ2g7rnohTQhLcfhFi0fSZmMh
GmuagCmbCSYyoR/Dl+uJRxYlS2NiWLRtzxbCwx//hNsT78bFI/C0Llcw+hBVYkzQ
Il0icHR1sGFOD9FYh3V2lWzPoCmsIUrjZJ8RsJa2zlNEsFQOhFdaoncaFflJ5tKK
4EIEt3i3YMO2YaA5g9HIsLq2OlOMmxJADBsirCYtl191k9s89gp7f7yKUrZuETbn
VKsXwE8wTwvDcGOFxwzqp21OLe32S2SnKfVVGWo6TGoI/Ago1fwQ4c0Kd+bS8MIF
oO8f1D0lxtomJxGDX8jeIVBPYn2eNnTtHG5OLrhWdss0dSAx+nMTaYrFOZyeulPs
sMlHbGRqd+u2AsCoSiJ5smvIe4pppzY6fkQcpsUFmoGwLIxG1k/UrBudJSIPiGB/
lPuYHKKFulPp4puVsmHZdoiqQzYmN9CSwQeeLlYWMD1D7C3CwTbNEzsWdGZCMr3x
l24YC85+LnXfNpuSQS/7vSP95yPDFtE+nEJjv+Wl70f+mBow/duo/ERivxJtvZM/
yD3lSUqvdyrFp0r3hJy7Ni7mNR/AksoKbi2tUCWcXDXfjeOOfNxcmJdH1IlO9ol1
GeR+DZ/vLBhhzOuoTLME+gYka1ZQpuElQomIIGUV3ugCA2dccjWb/gJtZGiklqdz
4oPEYms7ER/QvefgyjvbMM31yh2JevKuVUPJZR5+KpLNIoDGLj6SC7EPESFzXNSz
IoAgPUcfg+1EvHd8o3Sc/QQdwvlhgKNWmt9HoIWrG7EwOzd0FLCFu2gG8nwNrDNM
+TrmcyEFviU9JBx7gw9THe8FWlmDQs2wv7Az06oTDjLPO5OrA2zfMYBYNTnTUMez
LX+6l04OaoeaAUykOIas4Gy8ZYmX2ry95l0xW+DjKk+H1Af7EWFmMxka2u2yZ7/q
yGKWVEgAWgHe9Gjf9tGw73B0a/luBhCZqDsrZ0GP/+lYnKW8TT1El0Yv2qMv1IyW
ReXIy5sOzIZ7zq7qTkrK/mCMZ4X5tAAIjdhC1NdEhK+lJzLzAa2/gk6/N1pBysEh
H37EBZnBiaEJPOcETABnHdH3aflKfQ69FXe5zsA2ta+e7BID4T6RRGJHVhBHKpWQ
Iau87qX20lc3y44+LS7MnyIHdcZFs1aMIDdlZUxJxobc48KOYmdIOK2X9jU/QpSp
OltBfpLwH8R56e6SlwBGqwm8DsBia6DhTMgd6iUCzvQlnDUWH7HVZstIiJqktIaz
P5cZBiORqaE9QxGD+tnTkUL1FpxFjqIPeZxuGKpAE3EeKyxqT8xLZjax5yWIFj2Q
3Q24xjLsZPJfkIcbxnRk2fwzdFAMkrjadOU8RC9SPH8+K4pwEo/hXHGXcdvfodTG
O7YU+Q0kB/s2hskMDybC9pMVz2eVfYK0jxWUGuwpFndpBiWnnrd2nQJg34jTSm9M
C90EtPzu76SSLjk50/kjjtpeCkU2jtCaHQUsa2mqN1jy1knjNT70hHlcDsjG7Eum
lzxf56nfAvh4DogAt2V3Mw6fJKvboAU86qsrWEqjZ0GmLorSMoXF9MIA/6c4rkn/
pl+yXRAHpTCOnCMYh8Vtadtvf6VWso0ZapGq2NbhNVTHZo+L5OGGzj5ScvcM3KYI
08uPQTXCwctUudr4C9eKQh8YRaeUoh7BP9H/QOca3JvmwKUAI78pGz1POqcmfGQd
ArmIHL04/swazz3JmjXmOrimJd+lUzXu3fvvU71L+3HfboCPP5aBThSLeRhLG6uG
maHwQoxjPC66EyFN/0nKF4hOh6zqWaKNT7nTR/T1JSXRD3jdN4z/IS0fUUi8bmu4
aLLWlUcPMZ3dzQVuIfZnpatu6Zmu5pcjo/608Epg0DUpNIpN9VxPFhgNhnFqebAs
NpZr3i+VleyCTtJV7mX3nJkXeILpKHxAKosIiRVo0HucpegV6e653JRDyrHnkF07
c+g6Ue8iEFca7IFYLgh58dmI/Uqj9H16+hgh3F9bbT/41jA6qcECMuF76amHl6s2
T9xnvk0RgZoUhpAyW4pCp0b5gfDcxjaJPPwANKMgrE1advM45M5E7rGMzoS/011L
SZi7cRegwdbzlLbkD4IdXuj5YIMKYTNQ31xHUJFZtfG8X2KgQlju0JQZy89j5Oy6
bTQw/8D5c06wrFM4ACoKKbFaeUk9ISP4ee87EhAIO1FPcHSpKPmthGzihbHI9J+8
Vq1L2kgtJZQFu92wlDH0vWvi59KD7B+sB0LnJZ68CBQ9t5zyDeQ5wjWyKoDP8laX
CupirSLbfQozsiLFTWrWubE0+DpNd31jvAQGkibkMN19vDuctIYXvwEXo8pwvIrw
mGy3zwklN+CqI4ZDXY5VZOyw80jKiw7mRU9dfMOSqXOqM6R/RIZjsbd/gYXneKkT
QX2gV4gVLtzXcPRYhC2Iw/KwRewGgemreAINsOCUeamiH9Tk8LwxK5ZgdcH2/P57
+iv0jMNe4CgJLYyEPgrWymh50yDRaxz3LcrviOD+sHC1/Fa82oxuuLhEj2QMIHIe
izmAOQq9AW/6gQ3p+srrhEAv/vCy4QHpdzn59zguuphuI6S9IbjtqXxyFazAtRPv
32azpbfPSwgZFpZRjR2BUmpb3NA43UV57o0UfHtWxQt+OvzcTXpIewJHbwjWjeCy
vaVR23odqDwnodZXm18X9fBtZw5RVO3M1s9B8sHXSBGPoBc6YlBHMw3/wb54V7r6
Xu18dvFW5YGz8l4xdD+MxHVFjMN5llrttLR8S0vbnmlH7wQPkE3ix5q87PLI6YVD
C4Jb7fsWfShDJ+CnFC0h+dW+Keqfj7rbBQIqricKFqGf8Lg7Ky1hWxIvLav3du2x
tLBlujkkPek9I+Gs55yyrqR+qXPz/f8SDk5mEZvd2wmLsGWVeqGukbysAmLGt+Y3
TpjB+RCPd04cTGqJaXlQpg4u2Qj8sfVI/nneyyZDMs+NTeDUPNycblTeznjbQZcK
SHBrDe6I+q9N3BovRw1l1rtQd9Qp9j11/+hhfZx2QRgHyZvTPoOp4o9YTPowvn9H
Ngvss2TG/2hb6iwheBHE3nvRmhygIP9rBGOI99pI0RgGGZBaKkiKVhC9f1kLqikd
Ym4YlTn29/znBW/zSy1vv9Q/Fno5QpZtyz7BR/7FLXwxVzilyKO5+pIvmglP9zRU
Et9DcCjlFsgNTZUZMa/c0OIngXXFZN6UlE/BSrBivgd6UYGARR5VWle+7tHsSrvf
CtU0iBd86vwfFvJdQ4g6c6v3wTiwATY2mxb8W+kAHZRjM/W+dEDMD2a6Y0eS2XDR
UbwO+jvXMo/ARH/VMDi5PGo9MChV5AHBV8+dyPdgW+SAhZqCNyyfga+bFv2Kgunn
ObvVMPfHyU51D+VjrcYyFLoMBFAo7jnnKhWZG92f5aWNXmadQ8pV/1ihNyloKrIo
BI/yl15aFKURhwn3+SLRSAS4SdKcBReLoPtike43P4VNt5iuTf26MFBGmzoP8G6D
mA12X/uSb15H2a6xyGazc9I1NEyrcnc19lW04gd30rLDi6ffLWCiM0JEWqC4avkW
6jRSiiN4+08C6qN7uEIJeBrqk82jxx8ZNuNoGS98aAGInv4vFYRCbz1BU6nOaqw7
Hpe+nFc/DH7ejuHQCFH8naJq7M3IIN9l3KrCiEe0qujz4o65Pyr5TGTxB4FHtKmR
HeDHEyrYC5MlI5QOkfqVE+D3piayYc6KoALJnF/5Fcx4MnkXKfn3ptHDOW1PV7z5
raPp78aE5Rq9ZkCBgByc8Vpj9jq3gLEaGHH8WS2zaioVhphk3a/eVD7pUSLaCbWH
37kNrZo+HTEQx54JHGwUrbtVDEpsHbxksb5+PP/ccK6K1I4O76P/Tisr6/St4U3K
Af3SClHdkv36V0TPSNAmz/EqnodaiXZtpmiyB15VBE3sfvM2lhnPjMPS+Hhn+Rjp
13uugamfFjXUSeCOCDxNHw/QNFFxN8NXl8QDCUcteb2y6reSOJsW5z19ggcI2G6b
IFaqHYILVCpfF2Cyj3CLmb5ctcA7dFPbO/JZc2p/IER7KWa+XoyxNLohTQdNuVzs
Hnd3PngTval+MigwiFVGHQFNcf9DD83KXHaaDZgkB27HMT7FL3Fga/rbPU/q+Uus
6TQVbEMp2hwG/bcuqknutgPKhfaoed8kG/cfigiw6OT2x2ElmWOTD0MegXyN0is3
AAsRsx9PRSSiH1sxdtb72bsG4yYxvcJiGihonAZp/M5EsRbXWG3FfZRNRwQtEgYt
oBikGKUb2VvCWvzjqMpSBl5mM2oGKJOCTKjVlodwAeaTF/v+ozFRPx2ZqepvltBS
eUWs4CNXzSb6B2TG+xGdZHs3h+oKLD13KNHf484q+WwJw/T/zJoiUKW1wlhSSnvR
0t8Ars80v/Dh1DG4U2Fwo2vzlxO0p99kcK2ZDVa5yv6vFKDex/g0HU/faBur2EoV
6AiaQIWl6TzZSM7tT5bwBhR++hj7+krc9TiUiAfjziKljnlnicYI6owQGS2elBtk
RmjJdMEph1/U2YM482An+H3YsZfdbsLcEgxpltey5pgPwuAs5XGMp3FNiN+/3EFT
WbcE3xVqT05nZdZu27ONl99vJ79nw3R/r3bL3JN5oco2OFEmQFcc31Ufsa4TGs+U
iXlIDkqa1ZWvxyO0Pw7RbOK4DDHnVbKgnCXEgrRs8H5v80t6daA9es/Tfx00siqf
9TQ6S2iZNuzPI76ausYkB2GrO8S89X3D3UJjF2NHe6h067Pw+5vVI1WPIz5hFNY/
Rt8BSpDcp4vPtfsv+i3zvWN047xfSR9ysIXDahcZFZ2OYidXNgSBf6gaO5XUSKE6
OGocWtObjVcTvdEV9PXTELlMyJtIBF3vgEeFYCsUOeGtck7sk/59Y7EIWVbxusRM
0V9cbDoq+5bHTHTO9NsS28FJMlPGr6SydvdbuKNrL909RQjEExfcqVoCbBxInqwO
c590UoEnfmat443XSDzHRBkuR0s7RRNpLRLiDsVE+wBJyvoBbYx6UfYvODWUTaIS
H1+YhfCZFSKSiZ2cIB8JYoHK5VEt7ryAggPTkMPQG21G90eOKI/cDsXjvl75gkP6
9rheLfWjo5rO43o3788tquiU1wv82/1hKSPvqVobQVO/vLRmaNyfhQpNUjwPbTfc
Irhc7WBYTkEbb1au7WCg0fUTDVkkzgnlwUcb5FlRrunkI4bh7eVQt5zrqHbl4VLR
vnj/w9spkapz+Sp0cvf1B/jpAyJAuFB37iIZFawZSyjeK8yHecMGoNIdp4nXk7Re
ZFLp1xPaQee6dgPojiCStA/riHS02OcMCrhSl//zed8f8w1Y4WLEaBSdmpO9AsGm
en9hMLy62bKIasPICCURoFImjl2i+SuMSQPIzWnMYmXuqNWDTYA1vHw0ofwTlF8o
2dLpgJ4+bujHjpIFXtiuaKcLkn6A/fRx527goEq6nLg5QnZ0PMIpj+lwv0ouJAhe
19iELWqoKeDxF+xpna89G9tl3DYXFI/1zcb2DREOYcYDpTi0dfit2O7o5ljINhI3
LWeo8K5bPB2l6Wqmmo+eKi/I6RqzytM5BEeoW8XyIxjmvLZ5mDd1gCVDwoWv5KP5
C9HfdRNS/s9x86VgykNhaaKANpQf9BU2sHfg6bSiDGepc5SK7OrCNrneDAouJhdd
0YVRQa4Js1G2JUe7yH8SOr8bekfZoND0qH/6GGX8X2HxSF+WTX3pN7NWhNDKBWVF
JppmB3L3cZZ2Q54h4iGUoYeN0CPcDIDTSY0z8iDNFtX47oEKLe6Q/8hBcXhJ/UNe
n0ieWMhJF30GmTnq2LpuoD8dZVvkqw2dYtOlwfmwvHNrYK4pyt+4ZFNDFqy6I8de
MGESg3sauFhAACofLhKbLO6cFBK2Ay1kg/SR+WtyTcI8S600SaFvQCq8WxhgobLm
HCHYgc9RfcXqsfYMCZPahW+RqS9HniB5sG0uHqdhR8Wv5s3SARyvHXpSQxzD6C5H
ZtuoTyr8bUO5KdZBdRUhkSQThSushlvdAeURUn/pw5BGVqhp7W1spS2oqXOJJTMu
e4+BCVT1MsdQvvLQCmOyhy+7c1pDp39jZI7ea9mmOBRlhmAmEd2oHTg8ru9nKZkN
vxzld3RHyGM2Ftj52fq60HG64dmljVWBVRq4KwNQl+j3bryB63ddO8953COVmF8J
NcYysvQ/MmUFjMHv+2Drmh/lZ43JccsVMyMb0fMVnS8+paFySP1yiZay91CwTK5A
BtWMrfvSTdLSxoEf1yXhSatWiaL6uFBszoFlQsFJ9SNRMlZWIhzIjDUUppdScVwI
mgp3O2Xnqje/NH2XcfAHZUgrY8cZP6h+AezJOClMorypizHuAfM4VNHcouV8FCCt
IpTDh2RgH0VwW9J1qGmF/fKuOxbwhqSw6Vxf7HdHmlzyVc/m02Ao0sdXfyFjz8Ug
kDRy+OfnISQf9W6VIg5VPUh6x26GH6wNR286m0b9gDENyHpUHsPAFizjfhHqfpFW
D4uNusxuv8fuVLWBw1iKM7ZgKc5KkuhOUGKQT9wNURCySTDm72i2uSfXHn5IUIk2
wqZqar8QIhXC4FQDw8PZx1ecWph/Rrz9gM9dl9cKFjNhQPsCCGRH3XYc+T3R9PA+
PiAUT9JvZDttRSup4m1CeX3PI23kGwKPvp5MYHDrqS5u26+BmeMbAJ6s95mzBfPm
J48d+5uIkEqPjsq6zNU2iq8XACVXtpw7aeCuDsuS3ZJx54iR+XKM8lsFH3tfHSHl
Wovgtg5KlLlabaEzGNdsTrKawr/S/z5h8p3EpYEI1jDIsJCwhAZ7TacXhWgtRALr
pVKlLqkNKftzFs6gMIqzucKPNtvY9IBPEpvIU3L4ADpSQ3UbvwlDEGv+xp8H1voz
FObydsrYbB/QoikJYmx0xxL0vPyCHsKLX6XBjbcTOCpu8NULLxXid8T11Y2fCjaY
HMy2xzdfpQgNreke+ZETIrHDLXjYQ5jQ9Ka6iXBgdexBT3tgke9nIiL4tLHKBDPx
kF+6SUvw1PsU0jGMsvTuXmSfEhd7w9QuYuU7F9L7uUSoUX8e0WpTb8gE/raXlkCS
jX+KXb/KxjcdAk9JBoP7+LMHHYyAJDRISe7diCW3ezFeh4js3J488vQ38u+BLzKd
nC8fCGTKVkfd+MeFG7Zxe3WMF2SUaH7gU21YC3rVp6+h9W5l9a6wmQgHCVg2BuTc
2ETzmxT884/aK4I3aSkPSs5pL93jUO6CRUJtjLOgkEFFUXTHQj6glq1Y4UipKC9N
nuadMnv4HGHiwaAdZJ2HgFZ+HOTMcJup/SblSOHum8pe7DcMxEg15N8BFmpECKuB
h8qtnRX8Dq+26jzEhFH3RQz8Y1NcgqcbdFUjD2Ecra6QsCUNUsxc+Qqw0y+/kJJH
vL9d8wNRX3rH1zOZn8qsE1agTmAyrznYSRlx1+BdOLSwQQ/OR4mgb+9FA4IuX5K6
rwQ13ui3E8O0U3qZyZYVkOFQu41behOp/8ogZnqkEAikyIpaXoRTTz6CBs07qdE8
2AifSxY1fyvIO17L1v7K1vGSzvv6U01yN3HxMnuafRFODICWYHbbpjRu6V5BcQzg
6FGlSnbMbGq7mSBbG7lo3amlH2nFl54Xe3V08W4TMVIbyvhc6Hz+eqfM3J5nA9Yc
olBJnvbPYrCCmytWJqxwXNM5VdexYmNYVg9jX5Uxh6pJCIWN/zh+20jfp1EdUTuV
9F46o2zk09MLlmoo8tIw/54O9h8qtVXNKy67SMu09BsvyjQpCPqt8bgldjf3efNy
HrooY632LVaUc97iewz9dN94vbktj9c/I0MQePNQ4YNDfeqKNfT7kAVHhuzxbHq+
lIa6WX5K2eTfcnODaVvJnyvXByeM6J0g3IeiggjCQyic9RNYhNYX6OXFuollpWBR
xqXrWo8Lcj0zJ9BhjCxpxaCofW83sOeQS7U0fuayVIoLBQZaXYpQDa9yvNvKrBrW
3NFD2ixoASRr2JeKuuXiqehqyJlcc3DmLrqZZNap+p13XFPhThr+O7h/isi7/iHp
exqP+LGKYEmtj4q9awoz/I4gqhtqeqrmXT2D6PncqCPunxmy+Pwbm7/p/hwqgMZo
2zUVCdq/vPBVqAsg9aklAqOM4fny3huiI8ValQBf2qCcS/0oQqSl075p6OUcovoG
Cixwr19ShynqX+RereM8uxDNJ2xMB0mtatB3m0GTPb2Pl2bZmU/orlOK52LEaBDi
qk2g4AtoBGMH28LkbqJG/NkKUyPkYK1sX96nciRE5qp14moburneXGAaT4sfwhFf
7EzXlnE7VY8c+8JXpbJ4XH/xKYpGs+fEo5Xv33EMPXONtJtzctNrsc088gFQI05m
9AZuuDO85KH8Y7Ss9TudF9KO8swrI2xCcyeiJkaMvNSQgDEbJUiJn8XbxchUEtxd
B1qkzlr1l2td/FQiWf6DzE5GKc8iz+jDNSNYXwVaakIYYFZu3joJC+ZGeR2HT83u
s+wtNO8Y9v3JElMWDj/spD3k13XXGOEn0/qMmkEnPHe5+XAOeODBmSWSM2Md+vQW
Uin/OSGZWJyt+oZmHamk5XrdMOSgsy95IX0yx3rEKyKmxH88nWTawb8dU6eVrUJd
CNdlVddT7u92C7DZzfQP5mcp9HfXWL8g4dGbwD2KtJ4wNjxrnmwmDEALk6ZA0X4n
kJXd4qjSdDU60jxlfHuXpvjHZaL9RsRWQiFIOFC0YIb/lmB5pcJtfuqnouQWARvR
2Rfr8NDI+Nau6G/C5AMvHxrDf1BnN6botge4DnKt6nJkhAUzMjsKVsi/LsHEf59D
SRObvFUvCO7UQrhZ6rhYxRKmNxna6YmhYuqZAv692gghgZMtBm6uYDTi6W+PxCiH
0Q+/20RIAJLyGgtwyBwF+CEl6rgM5ZRDBgkvCWwmv4Z4X4oVGpbKUAxgTrQbePO0
lMXVufKFjhiz6NZY3yVsWUSEHzOyr1OQRLiDQSubh7vVi5Kb1htsLqjsBffgQx0g
6WgI8zxRAZgls6fWkNC9TPJMO3P1anRBoxxlLI5UPTs4hk0FyF5NiGXDWv6/oYxE
1JtUXGaCgHkPA8cYzUmJ97Zc8JmaQXyQrmDE8mX267FQYF+eEQ7UmzKQIp+OkdH2
CJ6XxlDemI4/REibYnaTRgyxST01smtIal2m6vMuHlEqyphcXPBDVfuvxtGzGJFq
H5CHyKEjKYiKc4NVksXqXKScXhoX4wa9DjZJIyPLH8lJj810WjRMjD10S/lPYSeB
TeH+/xSiW7YxSR8+B78WVqQIrrXLvTP+cw6hHApG0H0ufBm75Zgoepi3eFzFZ36g
F8lwvamFr99vCp8TQ7ZHfP1Bt4DtnDHHa0K8Iqy20WR3iPCAXwqvwjb+7MXCHDFI
HJ6OFIFx72i2ZLeW8VsCl0wk+9lA00uaJDfcddRlHFcvXNGSjuZIBS61IvBpwIcF
UUC8mOVIWcyzU4/Y8M53LP7nm891YuthP+DBn9/n3GSh4V84QnxDjzzu17DeJXkc
xeDU2Pr8qxvk31DdcMAMJ7pXQAH+OVC1V5S3H4MwmD67VRn+5TkISb+lHVjEY1fa
947+fYtTBjMMMxBJIvPU5h9NS9VRuDL/4USzd9MB9lzgttp4gKx42c0eTMthaU/z
eQjqo2usd0t5ydwZbkD9b5mTc+EdYpdpelsQlZDOIoghqyp9FXC01o22155p3dNO
b/MnuBJ0d3z3UK5zGZqT/w==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FqTHAbMXhMXx5sQ5hB0ChD++eB861mnPIYG+eqsla7/7p16lCDmgd+sz9v0VwUnE
z6DHAzLVM6FsBJhZbZYfUMArNsbesuqlnFK2rKWMF3a0V5AFmsczoWeEyr0F+sLy
ODcOgwhXl7ov1PuRfprYKXXk2xGc9+ARB3cJi3aU5viHAaLpC02GKCO5qkfeYCaL
2QMOC55ZXt6+PR97ZYQJjI0qw9S7flaFsvBC11SrfjqLCtLQddVOC7gLE6ync9fA
inS0AYTLocBiri1QOrdfqA2aY1X8Fd+uiUEok68NzZDpWpgAJgkPHdWbTCXJfGOd
nzkd8fWCIffw4BUVQCKCMg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10416 )
`pragma protect data_block
F/xLVaIxn2SUuI/YxxXfbql9TnBIYZVRZaRuT7TKXAtX4DFldPmCAbD7wKFQBKo5
9bSb+g0mzrAHFZaIx3jhRAR161Di3eTSZzpNnwSi7swQWvyERKLuQKgtQqgHO0p8
Ar8ccrVAVXx0jEQG9z/jxbRZJUCXZS3ziC4HqwNP2Y1q4M5earqSNeTyNVTXiebW
qJRh6soo6TBtFD0AMEJtr8PIi3qVgBfn7AICniGx+JNmtB4Cz0B8aJK7tbsPPp54
wCMUDPO1wFHXjIgbARmDGg6r6KoosaDTVLLIWHCT+gUXZN9Vtuuyqn/8NFCqMoPy
DJYkMHUkf2sVEHdz+4y+hVXGd17UIpXAyQUqBIQ93W0jAoqVFw87ZTK9S5fGGOuz
w6z4bMai0FN6H3oSN2CGh+YyMxJFvgpgkUp9I2OFY+BnlGABoVEral9xLYz0aF6p
APfJccr6mNNimF78BEsqfqy0dGlQ7D7E4M7cgA/6ApMkKBNGkES7LzWfSS+jkvt5
OMfnk5hHgP+VO04sL9YNJ9XxSlPNUzbG5YMzAFv1vXmVmKxgAJkbqMFqhdm/FIFm
60H1giv2wtYkxsJ5P1Mp4J6T25aTuUZ4Ydqdfv596itwg7uCSbk2tsKw23JTk0AZ
owDXShJQAUVSodhJ1KLy23aViunIK0gVS/9E61+mJM6OaiOhBGCY/9AcaF7dRq1a
929Nq6RzGxn+6FdBYSoP0k5HKdWGS/QJLB2kaBJfXsZuqAd4qSF67iElhzxEvhUr
UoRHkVOC5hqUei1YbNBimmXePDaFBBGHcE9BScG5KvUmYJTcOsKeMNUKhNXbwgP2
uyPEYCzmKt1Hh+FnYOFw/9zyJkdfXqtoQCJUG/884kPttIxCpXkb75w2QPM8C+q6
WTFwchi/239ToQOp8sBaS9JOJ/md4lYgjXWOgr7Cqov69znJdoF8X4oNQGik5fXT
K/OESXSZKqcFsqkduCywwA5i+rMVoVb3tgzZn88jfvvBKUir1/eG28dgp/yNyepA
MgE+qBixAaMfYt3tGguX3eFCIpdOzLAlan5jvErnKQDlk5Sn0mz2NjH3XLpVm8mg
Sra5p+/8i7EjRTKdGWlGhPXYZ51l+cntnqI2n3vQkLEIzkFk9WJAv3Vm8+p04PXM
xCrJtiANs5zXVEIYAxYA1jL75sIiFq7Mz5+qpyA/NyLAQ9KIXcP1twlGdaOH9c6O
eVS0zYusTJ+D+zUeC46J9gOCix43wb/wMVuEwQtXGRvNWWIavX2RcfkkxQVwqnGV
qPp62JC75GuRt0cDOZcaHVTDnd2/t16R7KBhVCmDm8dqXaxUj8GlqYcS2H4vbNom
/vIfGgAeozDaqKb1RFtQFYKa65z415PWFtTCun/eijQsEaIkuEqa0oggn+Uk/+6M
HGpTq9khh/nkJ4yPdbaHKPyk9na6eF6YbGAR/e2r8NDyXqIKMjKWYXEuSRqgOLdP
MGhNRZfTp6nTRskzkYQ/SJ+nwA3cd2a1SeFOiquhSuRHpNQ0lVGJZJTtgWw51bMs
ZYVGP7XX+CDWlkElZpBIO8pII/LYwJ7U+wCjgM2Fmb1zzLd6kT6oSBCzjfEnfv/w
wbEV+mEJRqH9AFs9KK/dK6dhuzOsbdw4j18sjqu4vXwH1G1NzQohjTMI3Vt7M1C9
6gaCOaTrAck7uCOChZM3Vnu6zt5QcScUQYIez/UK3bnHdTmifWLhfaE6Hek5DvKG
CtB6e1jaluYIOVDzxgt3rAx3wMYxQvc3O1ESOZuhF7cYGoDU4ua0MoF5wNW0uAyU
IBYAz2IIhBlGAx3oecGRP+6CU+67BKdsrYi90+vtVh4FkS5hcf+Ndo4ejoTkeL2s
Z/Glku4UqKptTibm7wmxbDHFsyanNXlT3h/3DCsPg581L+zIEnVIteAbGJ89tbHR
YesLyCNPnhD6w/UPWXJeCOmKCc19OhceEYvGLxWS6wCdmEq/HriPUJxOowVajVhp
yctNf+P4a0zQ9PCb29TAFPpFk89ukFYdcDsNabMftMOF63atPEvsmLxLhOU6SXNQ
DgkVxyX93P2LCwAnJUOmXza/iYGILSoIJzjDmsjR+3twLUhJAzPDOBNfeJyhhZwx
hXXa4iPt2AjN6hWjnsx80I3KyuR2k/VfdF3YC55sFgRMguZONBJkRxmt4KRj17AN
k7sUWOfptZfS8cgxHDKuhjaN52/WaGui5Q0Zod1L4JNvgJX2JZOpKzHk4wRTYx3G
m5xEzYLd90wM7AGwNvQChXC74BHGY3qlRDx2MbVXyex2Krnk6f89apc7u59HYvMk
AnhosvfDXZQIcT+n3quGmBlUjq4qSQBmR/n5wpSMkIPcMpyHKMf0xxmhG1SSmQiS
t3BIBbDRG/8mzIB1f3BSacqFUT/AcrM3hl8Ees/NRg2J8n49/w0zHOvPNS2JSO+3
XJfZzzLu49ElC2Q+9XDSV3sNxkm4FDeQGguv/hTswBC+pKZV8zUDZJlKDIFavzYQ
5GdF8NYRhlaJcJ5Fw9d6Z7ohQ8crakGhP2ASf6s2KFEYvcLNwsfZCZn2nKOcui1j
a5sykRwBWyuAOx3aSxjRfhI0fhIOtgRZOaiRpkG5uz9boacYsVQiDtntiXpXk/3c
sJUxw4ZNe2fUISM8U4iFg+LA5Bn40sQVnkCD2tRMcTV4a+7AdOakb46hmCoImShx
PO59dfmVkR6kpMSIVIS59/L7e5rqtJux06AGxRlIK4jkpyYWe0fjRvN7qYwHwr6E
icv0K9i7XoHzN7OUQR7JayRrNHQP+H+GJ/eZeG6UFdLTOpI9/of3Zoas1IxhZLle
UMWt/oTjk9gQNZ5EVB5YdjyVr2g/WAv0LIrCmb6JwmDcTb/9Vzm9KVxIcEhzoz1k
6nTamHQfQEbdmLtxW/w9KWb89MRtz0IgyrS39TN4yowuCz8oqY13cuwKj29nvkjS
kLp+Pbwr2NzWg8KiBvzryiJKnLodYr4VJHMe0OwHIy4o0EqP4bQDN2MlgccOBFfM
AYeGR9TNnmmHn/RIbdF3ufTwo47gQMXoITgvacROYjro5eEZUU+2fZXsaLXhjHlv
kUvkNckIvX0/qGzIt9h6ztXGNKRmNmFb8qYWgODoMlndEfLCmHSU/zb9nNQLU0Vy
W/ls/iyb90tgakxl76UdA0gpiGlTbETH77fXdkrT7sLYpr+VcKtDS5Sj5IgPe//i
NkVnpsOzP8e6WJHsbpkIxkF2blhwGJ7CM7wkINGIHDfX0oPM7TOE+GwRMYsE9VNp
xy23+QNaOkmV7Tyv8M/Z5ow0mkPYIOORH+6Wtb06BRc2l5swT/EDH+fU5DEC6an6
SGqkN7do0/Pl26hOPbbP0wCm1jFCkkw9Iyw6N1hZCdaMTHXOqXoplyDT0T7bX9JT
ruJ7xdFsttj0R4oLsLJPbWxFvnFhJOUOeELf71shtAMMHe3k0TZjkRHEW03IGljn
sBfNmYvbvFzxeAGP0cZDtcnG7BFwSnlwEmBpHzfKtr5j70IKSIxXsXq2BvBpD7Dp
FQyRnebitUAeg9SWl+vMn23v9nX4MlRFcJ1rncBL8ACwm2oGzkZu2VB0Dr/s+my6
WLDjKPHh/rZBaqF0sKE4XwS+F40uAFe3Kh0yAOTL4coSu/o5UiXQNtmEmCSoE0K8
wNjrClj5aQpum37VAn492Cc709TFbsSiV5XR2H8HZ05MQmRQ68UHwJ3T6FR1GX0h
dfFqrNaL2tNjt5kq59f74orqKmI9gwDmL1P+Lr4euNQ6Xx6qTmUeAFZMUKLq4cIW
zhami0YzN+dfTgnMqdeWVT7wBgY6Uak+cUQUdrHf6wNOG6NtqZ62vFC9QYYQlNzL
cmU6WSuGK4Ux35KkQYt1j4/eoW5DhMK/J2rteyQrNUcaBi0Yxy6c7bFDrEmLkAdW
E3UwzQuf0uDJQ9nxFKdSvz75rSffZ+kH0WxNlDTmeiV3gpx7EuKL42otHCqu/m5d
QAXE+rgL0zxCm/z4/I3i+fWZJPF9Ua2v/+bAlbiIPni6SWIX49+BV/oSVuxm9ddi
4bYNBvwSJ9w0uCW67GUoaZj/EysKJCuG+J0kRlZQLhD+4tT41m1Wu/NVz3uatB/h
2st7zQlJ0J5vgGnFNIyte2ZXtkLXLR7pIRwofditPl1fgu/DIiKLGPbT47RuwM2W
h54B3N+87HL0Ng/OQ1fO6E4rw7x1BDkSS7iaDwC+FQusyoJ+0NU+AwWwJ/zWMx5J
11eF+XEMlmHLsDASm4E62fciVYf1tTCfaim71uJdFGnz3dBgb8EN5PQaD/Bs4wfe
QQrKL/MTXGBwKXO6AKO2/ic5qsQ3aHbuom48BIME16tyJ3jyZhzKEfFeDbarZndv
xd6th1bktT/MRX1MFt8UIJfP49OFjtf+XB36+gdcVv/gP4ffgaVwZgiBHuAZcR8P
FH8Adm8MjbZyiketKnXN9ZRaxyTuwMehvs3yuoo4xqyK/ogteXEsd6ncB2gSzA3f
E8itL6tXf0GMW9QBvO0McsxjIEZTreJiJ4lidq8s9/WSnz/Xw5+3lvIctZaLVTkw
E0toXnPB607+pMMJMBUxEVle/24vJ8iL6IsSGTFAaSwkmC5l8wbk2RGKTsM1h9hm
+8qg4B1MadQQOsPQC/RaKJ0Mip7pWkrzCa1vjj9MTcD5cBSYKEBhP8cwbpf+MVjm
OrmOBqdmfNvEThN+liQzLt2w8/auqSa84ZTAwshbZ/aYpr1Av6bg71bV0UD6rHm0
E3Y9wfgtnnSMPLT2jX6qDWhR+AtwXc1qSSyNoiPkuCuGIaltP0YxcaOVDitzNTVM
z21jKLM95FiQ7OIRGVQX2Ed6E6og9tkNAFcyoFWXS7IJltlS6yPY5xGgsItXUNUy
YMgzWo5ui8YPfpQFtzNURqtPyXuL9wEea+0D95bz2qBxT6wd0NjkbDT6ZFVo+i1E
CxKL3wanL/SsJDKi88TeCPImUuTddHPGcrMnCyvXYQDzVaMvBdIggad4g6O2/aCQ
WBd7b8M/CB0MqOINEE9fgiuXsLO/+bTG2pQpSGRWNeZiNkSZrX6BjcnuXRwc2f01
JCixG+nG1WtB5kCeS4s2xEZ5xP34BFEDw9wZes/VsoLFhZEsuDb6sShUckj3e1k6
6HPAzp1/65ZNf3DgNnFiV92cFLXu4Np8EhELU4fr106QgqwHME+mhZvKwJZ+dA1c
ERzPGRgLYcqo0YREYe6cL7esGkZRPkSTYv7N5Ns2X3o4zyFmRDf88CnFURx2Meg9
SQ3KvlJWDn9HZkRaVFMQ60JkpxR/itdwRxklr7k9F8VZNekSgRf0OlYgZEmemMOj
Xeq5AFKsO1rjWctuEvGZPDWxwSiMipAkzo0gayU9sdp5b4fjuLoUaPeANJ4ZIG9k
AZqHEVuz5QGcVXdac/sTu/rWR/E5m0J77axcHs1VyU7RBRLuitNbGgjklPi04B4B
FFcHtv2ySxFHKP00Ky41z6nR/5MPDTRTsfXKmIIlhHuSb7Dbtu0okiXzHeBID7T3
9ipsGda0I5qn/8MDKCQUk9Iyr+AiWMIBKZ0azpbF93wQTHP5JrjEOSpUaBtAAVwU
HakvgM1GE4mvylRNb62t+M1n1DQfNvdvg9EB1o3UjwZCOrAIe0EOgO7Qa3M+V+Lp
QFzVB30SxL1vqwUI+ZSbe3JKUU9Jn5L2wSrxqC+UdH2+GTW1ejIFXgkkhA4t4GVb
1OWNWqT2GgH/+cPVGNWOxH4+SFPfl6Cn9d0V+6J6zKMbXR9l2gwdhqNad6r2wYEr
NTV1xnTOHoE7516/YHPdm7U7YzZVghRYl/ecwvVpc9G54lnPr5xsz1JrSbCGyKoz
LFwU4NmGKQjh2oj9qBefMNByUVUCSJy/NZsQA9DvM8HqXjU48/x5yqFDrEmigua2
iUcyz/0afMdlKaaHtvxMbBPTf8qu1IAkOZGasae22HlBT8gPKt5weofWpTF6zPWd
GtAp7PUCSNsYpVWKcvUs6yDhIN/gyNarMvrmjBM8UhpM1tinOJT8ssyeytlZIeS8
8714Tz+2rckS+QTlkFZ9XswMZBcIqBm2f2APBk3rPB7Yl+G8DZuVtibypnCS7gKj
E+hETHuTc9Uj5q2n98Ngo//LVdjYJYAxJKuxG6khua6NRIyndI/1xhx+XrLE76eb
otGjVb7wMhTEkfqPBq6HRKgn1sYWxOkYin7o0r/7VexAnlT2vbNJ72ZmS8aR0Lki
I86SfuulFtJI6lRONCaXjdDTGqDVgYdK5ycx7x4o7ipOJTO5k/Q9q5antiTRlgCE
VtLCZaXs0q32ocUUcT9s7BMOIeSMtRStEFpEMu4xlHh7h43IORPVJG49OQriRnHa
+/rOw0B+qh6wWGvWWBPMqBfY530aWKBpyO+x6bRqlJKLYclDMnRhd2dbW2CjBbyn
l3iNggLGxCfnEeVTUlg2uCyJUjL+giu+mxaS9z/LgKnyA+qg4Yn1NqhADDKUgH/h
Vu2DTdJv5zLYUjCMzuZ9VYNTquzifjEZYK5NVQlBoYg1J7T1mrwWYAZoYhUIpeIc
J11ParRquegIUgCHOWVb/KDoYg739/VQciyCVRfKhqlwuEsf6GLhmcEhmA54RVNT
QGFbUIjD3MDuEopkwx48Rx247aIOOmx84YlcSQ2M5OnMkzpU2LfFqau7055fWQum
aPc+yrhPPwWZGUslGNMDpkJ2U5iAJNb7pIZwqMKOOLhagmjXZNf1coPeO87z8v4U
QMgGPPk4NLaTHNZMIVuiloR7DlkaOma8SvhsbgOOPeniTzHpQC1tkfiql7MZv44F
rkVNy62s16ihO8dtYqOZDyCEXZcekj/HKYXkqbbPPg7XiE3ly/V9pAGu0g2qKBt9
AIHp2RyOJKXKuk0iJnI1RPfShHTh8BvP5sWENL5hWceNkgPL2vfFEen1HOUe+ZWG
h4tlFsW3x5zYaSLtZmqGWETkEseMBj03hEFYZG1AICJ/1eOnZT45d3fz5w8lq3Zy
w8RT+Nc/xX4cdzN2HcXn699mhh8cvaVx/QzmkprimBzM14xHRzO9wCSo/qFFhfDJ
3Nx+DtgzUzczpPBnrDe7LGm1DjST9Ya4NBkhHEeEs6nb63sEE3nHAohWfeFs+/xT
vRO12mRnHVybv6mRHuYBM75OdZrncr+U4zUFskIRTxVIVqN/uyxSzMj9cK1RIaH2
htAK+Rtsm+Hm/lanjrXpgZUu+zYhnov5MUncSfQ3SaYtuPM1zL2ziRjD3fecX3Ai
EdE3EdC9ZVmsgu6NAJ9Cxiovv0slGm0y2o3CjLDC3Yu8REUVm0bLhKx/eD12xDiO
BpCg9dh/F16pss4xB+3lLQa5wjbY5Km9Y+bHqA2RBh+RMkedkfzipVYjeGX5leL3
F+C5MDYO6X4SgdIHV6FdqFy7d/F4H1YFItBgIB0SaM63yuYv2AtDASkRTqWLbgkz
yfFba8T4y0Bv0uOSXyj0bML0mF3gRG8f1SBkoL9imp6qZ3qZftrdUGqQG+h+8wWV
2v12MmaAfjXbA2PjHqHlMHOZiCimG3wRvYvb4bIYWPbP+7dnj1/hyzRqnyWn3iPl
rGC9iJHCNkSnE7d9+jAOV8MvYbkT5Pc0kbjV1twk3x+Xnp92AvzJ9nLBqhcn3ZY4
40USgnFMLcd1ixEFlAlQaV8uDjvQn4O6B370aksNe9FZG8Ay/oWhk9JezKu2PvTd
yOnRNqRjhg//peRejpFK43uq4Rj6PiFEtNv14NpKQgBLk9BQhMZgTnn4H2111ZyX
DbqUiVU7e6pQWshFiduJhH1MBTlmOut2s51zjZVTVKG+uFcgKP/UFL0YQyG0w0Df
rGEdJqRyqRLmTdv9gNBihLsc1lcg/J/s82eU+Y4oW9yk26GFwNWv/CRTsjUDRIFN
ZCB8zQq2oCsPIvdQ/97cOISXAio5yjfVQuS10aBQPGdlIFvgLcbln++f9S1y+B5W
PovtyI/ID/oJEFGD1pbjZS7BTxKVREhATLlIUwnS/QZIUCVzOm/TFXrgz7att0iR
65klIehSXX9K9tPFlkL7WKqmHAznqlvzE4ejv8Nt7dJTQUbs9OEluOjbUZDdgRY6
ZyhuOsoCzmtAz125QTS2toTKqJ3xKgukgBSiHxHvm6Qd2XUhCkHF4vMkpzxVUkx6
PIFrxSuUBYzuuZuerpvMQmX2ShWZdoqnuamfagQqZBVHCLZ2u49lKutOsTWVcE3t
5b8qNcfCsWc9MLRweuqEhmUqmYwRVdRoi/W3AwHadJlOLhscT/qIoqUWB9OazCR+
/Xeb3B1FoosAd0LCXTf9fK9Dc076cJKt7rwUn5zR/ZS4KBDUf9B6FyPl989s9EQ9
pqGAQJ828qBP4qDPSMuNNCsF2LbdywxB7IKOp3sfEdMOxzxMAnRd5YgUPBQbKw+n
kKRSvMZ9REMdjpOaYCjUw2p3CXo77VSznU1YUpny3+tmVWKisB1PTN/qJJEFWN1k
jfFbWX3QlheXRu5obrR3kZfMJ7IZm117OiDhQjpka/Yr0AL3hlOBzyxaT7AHYZvT
fB1Zt22pQrbgVRlXBEQnNSFnxZUU2pOUeMhsQvcmzgJi6G5YbQxv5AqcK9nU8Bj9
2O9Xq0WujCrZybXhU2jG9PU7aeu6I6oLnG/8mcPM0hCgygXByqwh1Fk7cIwkoidP
HDTnaYKbfiZ7XKm/b6Put0vRUyhQhinVIR/qB2zbNLhZwRwOUsDIHPXEEUeeCV3H
KjpGRYlEUA6T8ewG/EFNo+CLmUZA8vRAhbP6OT1GXhijS6GDRmNTaNq7LlFeOUfx
vyK0IVCinAujyuk7mRYMMF0K3AdYfmdLm9IPi3YX9r3SxBIsMAbGn3od/9wSzHOB
IdU6fSwfqmIWNACG7oQ6jeGdmDn3dNBacxtQrW3/6/IayWputF83qLoOqIfooK2s
1Hok8Fkiz3QwddmCdrXCTVxq/Foq6NiNnyKTd5qMeQj1kvbrmTYMkqWu+XO8a40E
htDKxpN1qoKSfAVljElRzOFOb9PB0Y90CZ8jjC2fcyh1XdipZF5ypPIgOVdopBaU
7o3n+hyyr/LGE46Ojx62s8iFzH8O7f6nzAsjHP5PYIiUCe6ywET6buv6qLcYnIYq
8fIuf6EqrZfqoHQ+emYxZAlKAxTy5Xa8VAQ/vGkXfr8L6of1IBl6nEZtUTac7LPS
QWFgf0Ozwd0DKWh8YmqH3lgyQ2xiK+ikRae9hacGRJwZuRiwE0JLxKJPPeRCsXJT
ltNh7V7W5A0rEZEzqe4UHrlo3ioeCq6dOyLuU3Z6U/THE13G1utsARSQ8XkCYOYq
8x46OG1jwRiVm7WMkSuROmvSnPlnfj8egoJBBeXf2pjLK5QCYbaHF1ouLkPEPu+v
dAh+BkPHp72giwoKQhSKterq2pz4HhpkmHgBl0nKLn74WvKitgOim9XEUoFphSrj
V8yl2m7gV84T6MenUf9nqxVEEFT1JW0BotrSTsBwJ+g4QmsHO2fQiNMBuDRqrXkN
qQ6/ScOSkpGmLwiR+2Te21tirUBUngWB/4pmVInsF1Q3Plr/X1r+3cr93PId3cGC
3HZC/uyUM/aUmXs1eBq0TAcarJoou3MD0cSVERv9DviEL00P+hxo2+bFDUbC8QOK
rE4P1Hw64IuL0GGfGuhe3pUnHNMcUvDkaeUQJkyLGS5JNf7ShEygG7RMAv8TY7lu
6t6jFdHCHEqwk+duzdKkDytUXXPd0m292jINn+QXlohZJhi5ChlikK1ohFV7+2Q4
3i5DSRbJiySVFhoYHWEl6V/7bMn31/q7W5WIzTNPsvYUEFaNIFCd5og6x+ywRdVf
5cFBvh/ZWNID+tTrO0UWpeOXaoxZpc+AbRMGmjNqedI7VxXe/wFOmL9ize5u/UnY
Bje1pC+xaVLWJlHb1ZTT4fHE7jOZK7au7Rp4odO7zow0p17Ww0EbKPdonxQtcNWX
dSGrUvXh6ZWN6sZZNolKk2p2JiE576QNOLX58FOxMDxgkuBBvruEq//R+IlK88pv
U16URx6xP0Os7MTQxlMwnTkVQIiWKUxZowtH66AhheAPOkCXwVKugi5QpAEt92a8
n0Rl5YjFiAxZ3uEIlB/NBisUdDCuGr5nDQJwtRRxAf1/CAX+JsZB5cVliNJgX5U7
9Rnr2bJBq00Qy9CGJngKkQA8xugSMrWsBmoYML+IGBbnZRZgdYXOO/MnplvQUj7j
CVZ+8qRsuf24QDcBvHP23tKBoRYw3iyYVeexJWziAPzI8VOSOL0lIu0Dw5eQZ3b5
/2Wp3WooxLuo8kWCLBFX1F4cj12nAe7UGIftbjE0j7vns6OuinPoOZxmERX9iIXh
Ceyf9HcEoEVD2b8fHQ9FHLAcI21MhTOd3kVgWdpLpUok9NEpENbC+3nVIxmTkyPK
XztH80kBvsBJM9ocp2pdgH3DpDvbzYVqx8a/+JuG7QPZAcHml12RgJYvg9ddZEFV
tIR3RbPeIWWYkDR52KW8W+JjWjbcp3r5gyRkGUbCGfeQvLoF9WpxsfN3I+gSpTMl
CxxrRmMvG2/XT3XXW0y3xvNKQZXhrZgo9NerTaBhrGpCaS+llLXSS4N2dTA8dKDJ
YWFSisr7yvmJ4B20Xy2RWrw2WDPI8HKcZbNi1t3iZJwiAzDQZ7GZOh0Y2I2t9MVN
K9N27yZm5JkFCJI9LKCINjwbaO3AhUif8NXDGcRcTqhqQG4JY99SMIgWH2tESUbm
C6jGs7YVCpfw06+1L0s9esDdIIdiSqdSifhvk3yUO84aJvlYvLq/8ma9FSUlKSN+
V22MizaZ7oPzM6rw/ChYPuYtkPafCuMUHDCo0jTzeLHEy7kb9rV5Pe9EQIVI220a
HufKSz1Q6/7ASKP8x6G2Q7hCVllIsn13RpqcE+00opxWFRaAoB1W5L3MSlGyvyAJ
TjQEv2lPAWBCA/JDARST5ecLmoYkQNr0hkMkfPdKIYJNpJ+IDdbm1Bi5gQncPKSX
hvyCqC4cRB0Rcpovcngm+DRGfqnzuOS7SHDaTg7WdShvJ5AtVkU9xk5SCJIBVb0b
VzPULnBe4eZccalcfoFWm3vdlENugIyRZC0mRWUeJ+laBLD7oIBXF9IeTLr8Xhsj
jV6cxsxLgCRR5lpcDaWuC3OO0i2Tox/4UnjJmf/1EL7BjNidNZOE98UhTNMOHDzp
WKgRmaqru8fLvuXwF9ZaT9lho87VumyP3JshFHx3goNArkkf9eG83+Dfyg6Vgj1X
Z6Vx5ULi23cdbswv5UD8TpJ7RGBLydXoQ0GR4fy0riCR/N2t6RRdvh5wqEFav3nW
jwIV1y61HmYhz1yW7HZscEjklEMHbzSsbYcT/ugn7bJdsbE0WIIZgP2LTIXTTaUS
uAAkEsn9Vv8SmCYtntHj2v1/dhYnRP7xlYqAX+L8HSKucjwaZbn0g+Ncx2Kv/4zV
KJqMHQN9UgCcqSKXzSat1OZAyaH8KEPP6HgevGvAL0gBTZMgJ5ixl9hEIQAbQ3g8
kH5YRYwk9W7GI/lKOFJ9zDzpQPlPhlctI5i9KUYDtDkLsm5GFFnsIw/Is5YFR0a/
U1oYe/ZWHEMrMJprLEfY/nJ0OeyoXQvlEGX7ZDs7SRwo7mzPap/oREvFlo/NkEoj
8KFHO55KRmTg1+75W+bjT33F8zxazy4LjzPTt+1QRFf31qys3x1gx4RmVK7achV7
uM8imdgWqSiSyoX3AhbtiLdWGe0xEnmB7FLm0IwPt6OOcYKo/7oTj56NVb2adXtw
0yRhJCcWeuc/Ga5TRE0EJlurd2TYbDUn8OeppSXuQ2d8FL922UVUkhKwo19yuN+E
KkE7h+XGzk2QN1XsRyqzp5RPKb9UNHrOhkz16EqeOAbC2XJFtD59zCH8sTWIKkib
Gq65wDJRZxHxJwyATKauXGXIM9aq6CSB0090kloscj7xnAqZMKiaa0WR2bJITw6j
WAdsUlxuINO2hCH+aTANWaK3DGOQIVVZ27hML8YowyskVJ4OdgvGnIfCbDzYL5MN
+LsTf2eHjGrdaqhreWrAutxIOaPzqB7cJfQDratSxQi153A/Q4XoEa5g2LdRGhUh
WfD/9Dt5wggqsV23f02etUikgrSqgGK/1gMd41PcylzetuW4JvGffTL9LIcni0yy
gCAv4L/Oyuk9LQIx+86NqVif+MduS+fMMJHDpMSyh15tbndvzcQWVK+TEymxMaSg
kwYSYb3BynAOoV2wS58sz2RZNkZbl/ZVk4nn2BpPNVhJ+Hu9UYa43kQBbsMWlaG4
PlbTOk1b7fBJRnA4UL2ExWePnEdvX3KaD20sBCIM9AUrLtUvibQHsDilJLFq9s9P
0Wi+KW91jHUpdcgR8/5WmROV8M23LRAyalHpcpmsKVm3LXD8dlzVwE3+jBcqIMhT
Ltk12YFbHyU1czwK8LRWoWdv0Aj1Upi3zXZb3m+Ke+E7VLkwDiMQTusEbe7FBgKx
8TcYhs2kgMY+DT0ZK9AqSkY8U8Sb4nheiQONA7K9LrqxIz4K8BX+Eccy+4XSw6Xr
mLnXls4+wjbHVZNtQrSlRFTI3K2AECH9T8MrM2GmQnEzHk8Iqylvpp1t0vgWzSlU
YtTsws/WiWAQLNAZ6Ryqi1wIqdF7jorziCcuOtrVds+FT83cAVRMqRKtM/RC+xc/
r0TnWXeUwPzr6Kx6cjVJ2aWLADKujBzIJ5L4QQjYPIin/QsOLzH2NcIwLHcPNgeH
ZWkgTS0WQuMcxwjSAxDkI9Kffy8CZjWd4g2Z7QQqwVSSgtsyeNuIzr33CR4pqexB
uYMrRZWWiHLQfhs9JvUUNNq+3g2GYaDZY8034S6Z1dQigxZtk9wZE5YU1LKkEz1n
KuXMCiO5NGJrMk11bx7yI7b/Kv0B2Q6HzDvMjqSIRygMaJRHqvkx/ne0eqemyail
VvWifHucidEFQ3koTqCDnJU2twhVK+GyyHwlkrNxL06C8/f2EkUA+ufApcrjgl+t
enh3UBgBoUajdEh/dhZdsZsgL7x9HIgtFkfYQ3G7ewn0D4Ak+FJPhdHt9TKA22Fh
nR8/5Umn0Iz5rezdvIKCBo8oFm40GgdZDXnOPVb2VAeZFE2h5VYs6n97fXgJKFB5
Ze1csmXshtKpnSa2ntdZYQ/7vs1LPOykDIcVesqm0ABQPW2VkWRtDXUiy3NRwX+2
66dQO/tyWnMQ/2bZRypRUA0fiIER0vad24oTC1PCrjuByeEa9HJMQtCgtBNRalxj
rBcAJHHz3yLhoCKu5IVgmK4pmjizMJF6UDGga0tQj+YQEmtnuAV7MXuYjzllFew3
j/XggqoAvXbpzsJgShySWWbqe0xZdaVOTyMMoiplmhSJ+DwET5jl0u1GgEF8fCbx
TeH8GnE0/lbbrfEAmzvUXEgLog9P5xnY+YkOxc9PfGyR/MQQ9os8SFQWH6sguUKv
pwSP19nMkZgNXAX6Zz8cUzKizVavf9+P2H1Csi9RUlgBPzisFbNDJXDevnBq6yC8
BF/+EsvUT1P7dkxgQsrZUIxvCjZ0eNjanps/E1Jt9X/SIrxccbu0JNrxdSCD4dBu
u17aQHoY7gi+cYmLLO2+6iRMpB9NXAJsvW3dVyN2mmaEsLOhWgunbtQheyTN+C+y
z49/fn+8qNaACadMYUVN6sf2RaNLi2S1SzdjXE0riTV42RW+piNGDo/wbVUlsDvi
/XKmzfC4R+wz0Mhhg/weLFHE/MVQ7tXJec85eGZGVw2JAu2knfL41lP7PdDtw7YA
9NVvrW0vmVpVo8y3AN3xfso4PJyN5qOV/mmzPgBpiYjvD28J/rxkHUNGBmsFkB6v
z0/LmV4fazcsgpwSc5xDO29GBLQVZcJmYbNML6bN5EYgsdT0TIAjHVK761aioFdr
HeSGqGkoYGMG58JCTVDAFWrToLZnmbOhniUP/5lbai45YDtVeRaN7HLyCsvx/U4F
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VtIHWytHn4mDHv8dok5dnmAn2Re3pl5d3F2lfP4ZimcjqVNyPPjYUca341hRwtDm
7ifFns7d7ld1+nVB7nMcucF/394r4LXAW+qthgMnC94g7vECaB1VUAwijgqzpM++
C0sZV3H+ZaFAx6FI/zkevJ9TqpMvfn7ubWwSMcA6yGTv8Mgr3azcJn+m0cNOK+i5
+Ner5yvILaSogFJQAIJeJYvf2wDkfcqRIoOwO3btcQjFDbLjavhAruaa05SZ3L9/
5NqXKVQ40iJ2vqI33aXeqRMA9SsRXYrWorNmtnqqXrarvLKhSVNTL4T9Pg+dToGf
pAwZN4tttLz2OFcyUpPGYA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
rBVitAtVQ629BoJ3dWLQFt8Xy1zKNAlx18I8BmJrcCNk8J4JRzz0FH5mSSGM4ugI
ovxnLPyx8O/XafdRdbGY1G4XvT+uTvxE+vU8ZEoquJZEZqAYFFnO6/ks70/Ky7uW
2AEQF5MRaRcEVj5hGTlKyyX6izCil16S4a3PpcaTktAXzJvvZwGaNJWItNB/tYgI
cj1rx6Gx+QgiuoL5lo200hX+hC+p1fTri3BqgjwePGOJ3ria2b2yWa2qqzdO5M7J
jOmyNAWFGHd60ecth2y07io2z8vczY8q+/sXv2VI/Sw84is1e1rg8VW3Djzr+yX5
0acKU6SjShziK1qVRuZbIoLeVZoGvtAZpw5BWG28FK6j78RGpUZ2KF/jUfA/8htU
nlTdJjrvYpNvYheLPgco0+AJtvwKq12/PzADfbNVhAyRrWPAVrq+poFSVI75h5Ab
9ihPr2hPpNVVV55jtgIVKQ45UfEuMcLTZhkTzF05eCT+iqTOySRRCwcixdOKld6C
KjN1XSvi9bKdNfCMp8Zpxk+YEs6+h7M/qxb1ZQbT7H6pRj7JggWTVUYzodizJf2e
DcJMSdLvwNyPCuFAfLlvnxHXGwMtfr2BhSoixIGHPCTVH5+WCE3lkxI1Oigh66b9
JdCyiO+Jfj6+k5AARwq5izWB7SrY7jffYuQvrJtAraHQLYhm09rRtpjtsb6UVBN8
RDKRpsDi9EgyslVm6Vnu/hERw99eGDTnjMJenDavARD+VQ5TNHjjHhqtjqw6YgFQ
M+5qWk6674rlZ+u9X9aChVAShpYWxVw9oieDM1K2RGRkvMMHOOBBdWM1MCqqmKu/
RVzzHOSE7ivjXLsOnUu3FMqK8iwkOlCMUGqs3Si/A57SaXUO3W1JE/qdBACuXgqU
DIMWsUKDrrz5ej7XURksxn2ZOlY208syUODX8RMyKjmv+r3fMEAdOUUCxEOMLaOq
qxHqXSgVQwmeSv5g9MTYm9p9fO91OEwT1fAGQfhmNBOEPWl04azJ8XmXr67JvVha
2UQdHQX6rcTXKnAX41hT7osj2IBmvXTofV+PQwGbRhjm0gdgYicc9PJhm40RBeWU
heeEeKdP6pAEe/qGA7umzIe0iaCeNbc239LppKhJh/03i2wjjBCGvE6BA/u4F46D
GcSVFzptuQBwe41EFh+bd61JF0MAH20gD9jx4JkfhLABpOqT9MalS7P/gq3C6p4X
ehd9JBNtSQRdW3vtXynaZq0eOTZdM09VgRBnof8TMqNoudYlpkuhIgn0j3yMNxow
3ulwqceCVEv6xmjjRm8JF9qUZqOiJB8MHpCDlvP3W+ZahDkA13BBhgkGbB6b3L81
HY7giWy7NQyI9dAKpcGG7N2jj4eVh26iYWgV66gAUmpzhPXOfnfCZpuNfB5MCrmi
aC2GJ0rmOY54h9V1owKk6XCQZox8rbyVsth0MSc+MhHscZUyqBIJCcKglva0S+SC
oVhi7MAGMXHQg1chi72NjqskTao8KS3l8bZXgABWkiEvrHKs1HMu5kFKk1oZKocc
WM7cjvm/Kem//PPqv9f2FapgEl1zhiJDT3G0SK6xmXjdKQwGA8Ai1oTOeR3mwIGC
ONOhLhTVLkX7NNavNcH2g4T1oMoJ61VNq5nBZ4kjo6A59d3McwRj7cgBoo+ZAw7o
MSAFH75PMXEGD/z0N0QwKBaH4TiU2sINKbPL8/wlsDUDgOmlVZ6biUduAQ+4DIer
jP0dbMQPew30PZ0oixT9/mY/zot/2T+rS0wX0FOHHyzoAquENPhrAb32R178IcmZ
4daRCod9maMl7gDZv97bWOnVMJb7ZRefN0WdKRpTC6tgywbu/ytG3TlJ1Z4XbBdA
09gTrR3lTD55549SHrhOMJG0jBPZCQa2Itg0aWi8VGOqAiCLOVjFGaUiF8/foYkX
8cAkm7cWyVAnZtur85Jpza0pjcLUf20EYcIw1Hp1cfWLItdRDNdiImZHzwO8AK0Y
182elZk50u3KSciJJXJMdsKqXUh74RIEikoFk/r9ggWGLLu+CngJgGiCtSr2a1Bd
Q5/zLPSHPFW4OdqqhtaAGmBeHg6YGtl74vQl++kMY0gWThLPEj7pv3MLKBXjHiGy
pJsgfQtRIO+iZAMCDpiAB3ss+skgmjMHwnH4aQDwB9Fe22Hr8+c5PiYS5BS1lpJy
+EKMMHo7DEE5NXCzfSj+ciBCWAYN9OmhdhU1R54ZlNQgHcif7Z0Wj02+ZTYbR0oZ
Ur6Bg30dlGlkrWuSCH5N9bE9oQoOOSUGrwY9ghiyAdK5jVVCPJZ2QOsmjKd9cnO8
Wg+joJEV9BjNaHS2XCD1uDrEThYK3ZwhqPRsGWbmM25g1zHq65ov3SNXaJIajqsc
bBW8IpwBLAhUqwM+IAaXS5xwwaeqUtP4lRHEalJ5g9qtmpmHmTnbXCG0Gk/VJSoG
OOHCngAimi205ksnvG0VrP1DCjfcI6rXGK/jd/koO/RVlOQqDMzYC3vPuobZ9ZyK
zB6/Zqq9zgJFsN0ce1VXpdlAzKhFM89xmP3eaD0S7ubWjLTz4Wdu0LilDIG5uDS+
6uiQyzPsEsy/nhzOSr9uWcLdosvMRWZQasBHXr4W7PUiMrxp93qpBrWi2rpWtwDW
qcU+gT25FGPbf22zc+Uxgo1Y5r0jY9xoIViXPkWsNti6b/Trp2KA+UNR/OEO/yrs
834OhPy0SEhKtsn3IaYAwU2UjpJmMdd353tgyxK0c7DY1DrYT51H9YvtwE+CH8qr
iOBBRziVPQ2rX7kQKF4IuDAGgPxLEd7RoEo9Oj+3yhcctbV60EcQF1OupLIiFAn2
+aZYrm/Ny+KA92uS50rrX9kAO5b6FTb5Y20UErm5Naip9GCR73casE95n1FdntsH
9Cc42JvNVQMyLZ4P78SDf1g2bQfBGFw46iZnrh/vqJR3TMoVn1oOfloePuyqCOlQ
Zz8aYxCZwaM65CWM4sX1gIrrkRS1tURnotNqi2gixWI14qYCjPlX+P/lHbEmG135
XRlDWRVsNZadjrVt9B7/SE1YNVkI/8enBmEVNUIWrMiwyQfyxdVYhn/6FIMWMpzX
TDNFoBpt93+sZVRkMZjF1k1fbuZ7ReEOyNpPjDu9H3JnJHZHRIP48aFUzXwQ1BOu
9rDSpgTfBvFw/uI1019HOnD4jHfhqEgCBfKJlVyupVuLFqwY6lVUCljBbDmzYNdN
qcob5LT/UaxfqKlb7PSSG5YozJJqLiFbqWsQEOKG26zWGMjHOA+Dav4x2BHSN744
+wfQbQzLFYFiTu7OdtbOIeZXa1lgrjrzkjelqRXTLNzwubwbq4TwRy9uZllyDiCA
ETV4asgVwuJrJ6+3ORTFitZnuEEcR25tkM9Q6qUyP7UQls767HXD0laSELukMzT3
m77Ps7wOSUDwAF2b3iBhWkFGiL8r61Nqur2NMcegCM74kWv5ugKQGD7Od2iLHX0i
u5SKuQIde+TFcLcLNT/ZSol4gCaVwcV93ZdULd9imsllN/8f0VqWTwM66Ydyyega
28dlUJvp5zn7ZcqXUuT2gZGNZa4t3zg3hAFgVzwOIVBM2otggUth+PLGO+6m9ExD
1I6/lz3hV1nOfvbJj4MKZ2JuLPY32cflPtnXL7ehU3Owd9jVrPRKN9m+3kEtimX4
rg7RxHW0LCLCj0WxPSE4lKoHGDAGWGqe8E4nvVL5s9Ydid8oGEkr9UYVHDP+J+SF
FjT2R26yPu0MWhBnE/Gd7YqT/HGYP0z7vjkdZsNKfL/kZ/XXPJ4lZlhtSHwYFNJZ
lN2KeeLctfmdp/3VcA10rpS9dvIFx2ThlAiU2U+s7y40Nmz6EGeT+lffr5pLCSeA
wh2p4R4r6f0I3Yx2zw4gre/yCQiPt8AH60L5K99L7XTMFZesba4X09UUNXEXtkoT
WuX7bj8A1QbPGsybF3ddrFZa3s+WQC2eVEiAeoOBYVvMQKDoMA1yWkD/Uth9+p4F
1aBI1MTb9WHHKtbRKP91SUhLOhva06XzkSrSNzPqnGgjPHxdeBYg+5Webm++Pvw8
ss37sSGrgJqH/VIQ6Gm6OBJVdFFgPuQPE/+6QU3w0kiKchsReisYNMvNv+FTdGe7
040mW3XlC2zbtCeN4bZCHpV94xtN+TvoCO6bFNFMK/DXyPz8yy6SYMVMzmty30U/
Sjx+gk53nRBUT1Ki67FxUec4fAl+sqRje1gqUZ89huyd3GrsM4LBVpXNj/MLQ3tS
enaPU722lBvrLQAT7zTXKiuTMhLD09hYL7ciLQXLLDYw5OC1nwHfckwhPEqLlN+a
OPf5WKr23LzlUNvFUlx4w6qLQua+6A0aGoXLz8xcGnKPxpgexXst0weP2ANGv5Tn
Nrwcx9Wd21q1PF4usDIRQSyPXOHPlE9LKk/g4sQa5Gy1e0pBpmzV/W2PbMdAEKvy
awn0/Am7nelXEoyNl6Uo8LEx7+o/XWPSayfVo2FD1miPdLK0fcDOFlDNQtUMEm5j
Okn16Wk/NDQHgDlrkFe3hYLMVp/UP4+mRkR9dw7ibB9Avki7bDIdqU8GvuFIOuyp
BYhbdJzVatto6ZToZ3e46L22SuAkzZ55eEwCSiMdI9bv+HifvIuvKBcwl/Y2d+LB
YuLVT++HNIW/aWaXoFiCtgNx8PabyJ+YkxTh9s7PHNH0aXxCHif8xuf/3fnV7Ia9
w4/dTgt9rpeA7JCznrQba3Oq9JEirZ/tEfCL8jruar/a/DDPSDQd2nzVgxIZR1yg
/def/R0VGIs9IIJccQHPFZqusklA3IRjQLRp8VbHixRKki4YRMVxskFY8tfUFL1Y
rW/VIdiP3BBwpZvTVbE/RPawNtb0omALqu/w4dKSU0OHBouZraAfTMsi2+n8PLvY
KJTFNtF2KcaWbHA861fJabPIlXAPuSanH39aQeMwZQ+F8ZiSFnXQAUN6sNINexsZ
1Qg8xsUJJzdSfGXmaQQE5mPgMLi2rat0WpvwUxiGzWDCin6vJ/DTRxGjeyFSKNfr
9F2frUt0RBXXnKy/IYsHrKy6d2ZrK1Y0BbUZG3tFIvGGJScdz7rsfdBgr5ua5KJc
pQRJUVMXftpIkDDKDorcAdFoN/P1uwiVZkWYaC9AZKSvhJXIytsSv5y9sHogG51+
rAT/IcuIHRWrLdI2sDr98ZJ4OgnaKfUqVIIOX6HGkYTg0XHfy8hTd0bI2uEf04+b
RwnFa8vOYI4VrDmmbA355Y9WVJ9cIpG3YAypD5Oh5hC83UQbvhfqC3m6+/h60nZC
STYC/qN9BiE2a79BZ567093gQO6GdtaLP1SKyXJQd45GQ7wG5vlovSXv2+NIHAoB
yAWskqfUAWwTq5AM+kaeZdTsAntJNxW4ARXzuP+YGWcWefd0gVoDwO2BS55uvu3K
OhMkuqKDgHGBTGOHrMDkGPYXgKoTvcPkRyY2JchQManns7AfKqYN7W1a16dhDJaV
ck5Zdgw8F3X19GhQrAUfZjLGRkMmFWUMIu2sk6VSSB/M1vqY1pAoGItg1m3jcL9u
bQJcGm/HrsI6FCR9XkG5xXYIpxUEFGyClKvbUQdyLopchecG31m4zlhV7NKynrvB
kyviKuINXINaHwm8QBK0vyMYpSq6dM7gJX/0Evd/Iy/8+B9H8ZWzMjf2yQEENHhs
1YxSsGPrkWv+H22NOZ7W/GzmC53/nw1eI1XxzdbT1ipsIduC3pNZ7MdiXGv4Sqa9
i4j4weKRgzhThliat1IiAHwfPA33tGkzzxSe8HjfWy0/qbbLZmqw3SPp6BBj8Zoa
qcUHTt6k3RfC/xk9ludvm/5Rsu7UfaZgJJaDhhMTXSe57DOaA4lKA0+1iTunpppt
zZbRr5Rmf+ShMJ0zGL6tuY7PPCA360uknB02ElORzXeu2pMeBMNlEOJE9TuSuNuM
I/xJN2u/XaASMnoV6uAAl39NDXJgj/nHdg47qhRLsup/JsR7TrHT12MYSEDDC3E3
05sMoKzyvuzNDOdVDJcZKlzwtox+nnO9pWKA/FEf8jft68OhcdlN1Qaf1sEMxdpp
rRsdVd1YHETatpJBH9+fso56JVOOD+d8hzFhz2mV8VKWMHSTx/JhbDV5mGZI7bBL
uKNJaIfQ9F4skdUynbHTxbroGinn84MqPRw9VmdtDPovDcxsTIISZtdu6IA84reC
hsqn3JFePQUxaVvA7w/HdjGkzWVj25U8i+Q6LWX4P5aNFQVBshpVZMT7cmRnnCr0
RPZpD8ETrG/FTnca/t/XWYwzKZ+KgnVbbAnjfYRbRxjHKxyyo+9kV8hlfqZx8CYa
gpNjLGFyqt2g4/y7kfsjtVOVqgnJpB87ZiIV9iSbbMlXb6Rda9+wPY3jcewgJC5+
kdEmjCUExMtgyNCHzZ/210OX/SyujKDAwDzqcmyN7qjbAzyOPLC0u8S972iaZVw0
i7xD6deEt/pcpMoSio54tTbY/cLWRIFDIZtYbHHiVJQFC5BBUNXBw6cWIPwFehxM
82msT7WhTS6N+DwQJ4uwOtDcZdI3rwzW0nHvNztx0NRKDi7TD/nYy2CsHw5Va+Th
I3gxAMluqyn2/k9sloHu1Ke23GaIGJ5GbhbSvnhgTrf/GLPNWxYQVhlPCH6lFjYP
KHlMXdhX7/GfDdJISX6ThutrxIumb8/X2DAWLa1dYa3QcmTZckEvW9+Bqmjaxkk/
jqqR2pvo0M1VRRd6T4x+9fBd1jDuS+M5Tac7GIfmMGD0Pk5PhaZAijeCvyu48zck
j2hBZpMtBIRdXDc1HdFl4fWgw1K4mmCvfrfkAVz+mq2CyXdfKVoIWeqdIfq8N7xk
7IR4rwwl6CLEWLfHlom58RZlEdlSRflV8ke8OdBO3hCxnsWFC7+mNbf/Qdeya7r7
oZWT+/ZUIIYzMWjxNobBqtygDqFzW72A4lXDU2tz8CE4OQE5BE8xlaC6hdSCAKTI
1hJLclQc61PtTasLnaAWvSThKBQmkAOj63acG9NIU5ovNA119yai7FjkdiH5uFSL
P2Ec0I8DAOS9Xv71EA5W+j6yZUOaYEFrEoXkwnYjIUxsnm8Vs8EAGeK+B96U7QOa
QmHaGGR3FL17rzU3Kh+kk0yJsQjr+ph2ugBZH99LhRWfl6BuIIz1D99XO927cZXt
PIlt5Qt491JEizmpIbjg3VcNqxmHoQKi+XzB4N1NjRYb+YNsoDsdFaxtzDJAUbmd
By7h4cMXqsahpPL3L4RKUCd0xwROQiA0khTsPJcOVeABcKnvgwDtXmlOT/QD9fGH
ttf0bNx6EmxfmEosorRdoT0wGAWgAeSsl7x2j17EFtq/JGuCw8YNocheecVoMx5O
l9bxkc0xBylRRtRD5kdqLRyvfRfMpiuPNcfaIz2Z0LGrOaJtPEC74OVnGvKcBTIZ
STYGXTfZnRUf/xiFC4aNLF21vN60ZAF+A4BjPXWc1E5v0Hm8DpAjy43b4/bKeE9s
2x1JwXIIebd8QUyqNNbyIktl+SYBPGrGpXTP+8R8i0NVMBw1z0pKk922Nti/j/Bl
RHuyGmBGYGBAFCDFUy9NNE6sOGBdTYZbvjLRgqCUUHcRnODQy/boN5aC5sc37x7v
kVb2yLnp31BzuoGF7eALjXGmRldf7LK6ILJkAOnTPQsTiXUZjHuzgULSA2Dl+ICU
RTFoqh9crsoQv9GNC8djUJ0x5LdECEx/Pk4S1ouPa0VhDV0hyyofZyCZqO+wU5Ek
mC11ysXMmGeDy+Gw7OvtjC0nn7kXd89SqiappevauRJdn+RKuUVKx6JvrYwnVra6
BuVWqzDVfkWjKC4ZisjCKqFiBQBEwFOmFNWM9HmjgIoGw7m2j0iSoXS000e265Da
c3h7ouj42XfsDKGQj3R2v1GpfOwL2uIpT2CrU4MLJAiiDlOO07LL9gFw7eJd2SjM
qF/oVkExfo9L2MWGWDEWOXW2yEQTftpRFdFIFxDNZ2dsQAbPuz8Kx6qdzrEa3m3W
cuKAFAudlKD79QLg14DRD3jdOV/NT9WqBX++YinvIudcex/KBbyLPcjmH0Q2sr5J
AMstvrDQDMGGQBb7w6zKCQ==
`pragma protect end_protected

//pragma protect end
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Cw1xoX6r+/SiLjEZuRQ92okfDd7E9wbqwLxnpAyu3A+oEGc7q86FGBo4g+dba66N
qhJ6yIcMCv4A1SgrfaVAC2ZMeqr9YkKhO73jlXtfY+6yunNPrkYfp7V0w830ZrjX
ceUSKgJV0FI3ffoe3ZWr9wXyyVG4oiOdciEnC4q6DGnHeX9LvAzT0d/Oz0rflmt9
UPHg9lHLSAHGGZb0QBhm+5CTlAELD2viOjYdBPtYp+p0yBJv0ZEYCQwRXhGyupkk
o5J3cQMD5EqdqmV4M7VFc9G65TEtrJRM/c0zTZapUu6EwP4Q49C39JgmVxHqd4t7
TYXs/LypLhTxgf3kEJB9Tg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14480 )
`pragma protect data_block
ngF5UoG5fGkeWU633BnzXZt9IXmuxgZy3r4dIANllIuujMZQfi4uSWGs67rzHX0J
s/UY9H0n3pEo6w0sbjg/t9QXgHBsUFPkfUKfTtBycTjlpKxBtKPvuaP4RFSKbrVm
PXmStnoYs+bj9pZJ6j3J/+vQ7q4nj0MXT8x4KWJD/90NVHzvot+tW2KGLA9e0P/e
LMWjjc9MEvTOtKZOUK9O6R/u5W/vhofBi6rRCbJ5O1runK/19uUSc3y1J215YhTV
fAgxy6XiU/e1m5hWpuJ6O9HfniOaY4TaP0BWQASaUwwPvX9bbXDg102H7oRUfjwj
AZPHjvQ8UfU4V0e+LvvRrqPYigobtsCx9olmbFh3XvB2ceRO15UupWKFIVZBKmmS
Ba0izRK0CWMInb1zQeG2lKyIFE/rWFm3jnXZYz341nUE29VKi+ZWxSFpzQz8N4uB
sbQYgMztj6rX1rCN5KRNHRnEVVl86uffJSpwrlJWRUftkVoM7SdGVy3KzAZdiNlX
0VuTj6Udw65JyqgalCDx8ytzkjJJTs6RbWTBAcO31KDMhe6KysbJnUJ95qSf4lnG
RfSc39ILQMqh0NdD1xC6jxc6ijVdgAaRvB9TpR6UY7kRzlIgCiptDmNyqOfQkVUP
pAPtybALS1O83fCXjk1EJj66JAjy9JSbG0gKiVY0EnbVujVFjeRrJBak/2vD4Z03
hyKWl5ZmpBMd/Kd3bYmp8m9G8hgQV/6RcRr3Tou0OHYh34mS7W1j7cktqxREn2Jd
z2iKeV5fTaltN5F84gcfROGBOew4tQyJG3HvLGiYcYZVXEvhhLf0fscvMjinRCvQ
nIKMOm72ksTVog6GXbLLq5AEGiA319aoc+Mj7hlX/L9iRDraERYVaXt9FDyNsUoB
KFsWUeb+rcaGSkE7jhwi/AJtrZwZRlR/1C7APFx1hUHMZ74x/FdUC8DVV2jCk4Mu
IOzJZTTKIHdBSc7FTTKWp734LfLV+Cx13rvZvl/gRWCJNnC7tOIVOLnn6aVvhIhJ
W5sv0HrqlzJHU1LbBG8vsb+zIfn/eIfOGB3V9JRgH6d48aDl7It2sSPbW3pYjvWV
aclgwQk/F/j+IHKiwbYwWqyrbtg4YjBEpQibqqJ2MnU9be5G8usPhr6QnSi9LTsQ
yHIhKuKDmbVzuzRmh7OCeMwKc/kwuV+i6zCFmZdbXuD6Sgt+wC91Gh2U56CetJbv
8hpLGk6wI2Vh9PodUS+WSz4dC/6NNDtNUVyp+GxVCDrI773TNFEkRc5FIlwlHPow
YcDkNQtO/VfWHtrK5CIjqbgRZ6KH1hCwXnXVkJkGsFLvxOJkoFWdGkR6vZRYuFZg
GzdXtarW7HM18vBfc/R11etMTEI2twzCYz09fAbxf/SUZ/Ib0i4OWS29L970ceFE
wyX+WZUrlTXL+hxjIkioN4l76GGsjEm8y28BIJqrcdZQCd8otd54Zilcdc+XOCHB
yB4E8rFftFNFxk8e7kq6AVN6v+F+FgCVl2D8Y0K17hCjQiQuI4VX7WV/YDkQg7Sy
1U9sGoBkFJoNbSry+nav0iLfsG1QQK/T+/84AwlFnqUmxt7xt7qjgW+kcjGXpAqY
TLo67Ado841KRhKCP54C+h/8soS+KC88JJwlUWvjhcupqi514cAYveqbDlPpbjI4
MubA4D56sfvnrMZHspAMGnhgB3chvf702VCH80DsdMBqQ3aHpqLl9VjIbQQGUQpL
uKAzzs5jq2MRvyhBcv1dgdR9seFyIiejoJHhx2OyA6Esm+9gDbiVuCJ1O7WR4wOg
15l7YnVMEByO4Hg9Zv++wC5hHrEZp1s3Y4zUe5XTuN2iT3xvUvgwnPU7gRKeQRJu
5SYYJOsFIQJDA2VmicyxMTtMMuzqNKgO8ty6t8zAkHqgzsIfmnuPUyvOPhuVgs0S
W2Td0JS0m8hHy50gVWldKANjqnrFQuYIUQ56kO/wgMX4QjuHnODHJJFGVNScJG6w
RkLAEUP2f46MRE+JUgT2HzhRBDosjjTc10ZsGmud1TnRCHEKkE+a5/xRZFieYTtY
n1qsyKzU/GCxFYpSD6giAauZHfxfmUkXmipeTWWWziZxUDckP8rdonFTk/EFwe64
HHjvcfReW6VOFVmU/7V9ZBZGCfyZeRFyeAc08QpycLaVt9vvLf4PE5dTrn65C/B2
9OFc94mRRf3VufduAgSQ5NPD+UgObqo0erAYyTYn/AX4O3fFBfEgKX7KiHIuQ84e
uiUTqQi6PWyCt4pxFmRUty9Qjmf42RowwxxI4Ab3OA5Qjh4qluwiIujkK8zuoj20
/p+5DGFnKs0glDNHGdDu1d9jkHRQ3ZpOJTcGGF7iCHjqjcexGVQ0FaLdhGBYU6VW
k/5eW896jnkXvV/SuDfv+c7dVgVNouUiDeya6xRrMJvUfSdIkcBrq6S+W3knGzDE
XPC6DkvcAXDEDmttM624f2ib0FOybhJUB6pY83+ddBzw1OII5lQKh1R7GYtLo7OX
8BsWGddk3Wb0+U7GyH49r32EPoF7bqHXsErwrtS/xjEH5ttaRW4VHRa4yrnaeF+z
cfvrHON0R6x68D4dehvn9N7IlKYumPDtEQbfMh/eH8/DyAOrQhDZj37c7N0ATLqJ
AV7eQudmxBDREMNyXq01xkoU3uRegbhdg0GIgu7SK90TO6dse3lh4s52TsoHBWuG
RprQQ606aiC16c4uy9oOVK9YGy87iG84pQ1Bg1Z9zFO/CU0iIN5RJ7V1Jjji1DfV
YiidmOVkFFi1aRkbSxjQPWyM0RyGpe5BG9Dkf8dgJAcI8Ftv53hSqcyLK7ob9hVc
WiiSLmED+verVUbcvZqvdknfP4dHlIa9GMXNVBQupeqq/u+ceGTZCf9YxwoDpc+c
omBgm+/ENJG1ITuZ56fpKklckrUfACPz6TXQH+bS0r3is7GnLecIbjB8/x+TY+en
FkqgxzWaICKOj6c3ZKzVvkNSkdr+LEwvvvsxfvxkEkoT/0sJLAB8xxZwHwMAK3AU
xMvMLVVrsjVEl3r9QycGpLeuLvUR+WtcOFZhm+l2aSw5JZ8/EJi0LvGIG0m+6Cjv
NVEcZVHd7JSFrAM7UtiKSSSy+9IpuLZidEeCikJj9eSAtd8p5rBFE3x3TSz6a1lO
OK/BDs5BYKBdaCdhVBdeIQUSHv4TyLO3Ea2xaAzeXQ1qzBFxQQWu+54r8DkfPv9F
wSbKyg0NL62WqUMAyZfU3NK/urSc7t7g1UpgxCBzIWCGPQ1QhtnWMSvGUi+rflFj
rw29LptRyIh5alKk2HmqVJYsoiqZjKaIqbBU9qj1RkE5D+Int2utkFwPMAq9Hx8f
Tngt//RaRXuasP0hkbVxb7O25cruMdg81TLqHSd8adoEEaApVJ6eX5TgbB3zzP0f
dwb+SKiFTxCwZrt8jAIxexbjLu4A5BYNM9hn2/K63wdhBOHY9WVUBo8zdgVE+Ptm
kbjjm8sRtPBYNj0vZlT+gFWcyEEHfpmTQ3cnhJwNJZFPCvtkOBsMqutlj5w0Mqwa
fvVW+iilGryNnILZ+3f0MkSwVuJZdAhrQK3HBDdb+0CT5FM2AjieXHInGeQXMxve
unvSTZkOy7jiaT5WUDD8cLRLdVbTPreelA2b3o9JMjzEqhmWWIISlSa0sUquz/sn
H6aokYvxfuJlWWibyNyqsEoGq+RlSmpPfRvEaGi/i5nrLHSTS90rZffiSV0bq+W2
ZUZDIuBWGZrWKgqZhdCnfmFt9lZtrrpb5PB5SsQIhLy+8peczvapAyOV3q8FiFRD
T0qoUQyjrW/sdv8XnIyhkFdfEBDbgIvKN2Fv1R3C0gDHkDQIXs2X/a7HGlIeHO4Z
tfxSR+hY8eoGkoFSlhewHtsJ4Qqh0fn88///h0xGmqC9Kolwp4u8TkXEiUZ4Op0S
gUWzMmTTm18WzBP5kubhS5LD9vD6mqArQDPaWSEe5X9u3xH9Ip7FkmkdvLnUnvgw
+0xigMIHIf9d6d74I3Z3uOB/HlbJdKaCuDp8mScOZ34r8OsGbAFL6oj/Swu0x0FC
fcev19iZXTsf6QJ9mHqYLcQaiAvbj8s9xGogY4GvAbjoFnTPr+9L4/CvpIQMh+mK
2gEAfzzbRqn/Tcv7GqkS28fb6LQR99HLQNQ7FKOLCmq2+r/3k7cgnOW2vPfTtCBP
nfcFy11hixg6eHe2CpcMyDgSj42ZnlVuMQvBlm/oFRmayok7vFHWF+cQH2QcNu5Z
UCYV0269Mag2mUgqrc9kvpv+s65byFitRnOLKE/iRsTn7OqCjyOScsnSTk7Y1Lzx
sR43YMlYxqpIg9Ik1sIQF2GG+AQ0bbL5qqQtZT/JRtUk/o1M/eiMQR4VYXZ64SI4
8ZHX7AbU/PgCp48fm39l+DZkU0UGTM8cFM/v2cqBflxtk4pPoIj8lhQkoMotkpN3
THH32CPCgTR/DAwUe/nD5FCM+llkxALwq+OR0U7v2zfwURCnkNXv+8BTCir6bI5X
n3xfwH+ytisG8s2dSynfrGdbCXh+xTQIQ89ENatIEQTp7JrY12mh56hWpMql6kG5
lEz/f9vkx8xNrolAOdfeigFRmO6LHJwOv/FSx4/dl/LOAjxYZgmTjfc8DX1yPMli
0KsQayG1LNvcKiv11FjnEF5befavIYCOzHiLPHXM6R61yhpkAWUe4CGTNbmuqlak
S1cBInYPMjFCqb8sln3a358YlR1JZEOJIxn5/V6LzsKLGXnxdD0INYHUE5Uo2RC2
+0aGEsFbmbEF4v/58su/5kegfJuyvz6Wa9rA0Q0p+F3tbt7kj8ypXgOpIarXmdNQ
sHds9hd5MB3dtuyyihTraaQwMyIiM+8OqCJai3L8gadznlqlhKobncMQ2SahPgml
Z8Hs/bdmSwOK6Jr4DZb0l7Fnx2geu17v0HuAf6B1JwHRzYf1xNhDcTr68pGDcNBD
O4LVfpHhuN09votpIVc7aWbYUsOgUK9Janj2OOlDBKn7nOSrc1Mg3bSe0yNmynPE
c3DYGPSavuSUyLs50EgpINfwfka5Uze0CYiQ0jg2cvVLaYX+1nrd/0piHNQxAn46
uDQDDO0M087CcTb1GBlxpORorON/PTsMp7Hd3ADXc9SerSCdli924WIrbIrZqMiQ
sYQkcBiWYME+XeiY8lnpoxnlrFNbeRwXxCIvCuCQhw/52OKQ2/asesoDEtEfvQuN
C7LTdT1OZWsnTeWV+tMN+55frmSHp6zHva0aSptmf7duFlQLWxord5kz4+DLHOkX
TjdslTjW+uakyADE3PT6ACNm51TNTX0l5wvbj1lmZlsnkbj5M4yc7JRj0G7bJJ2o
36O5H0G3e9GuzQG8MwTCHT44tys6cRsxFjysvoD5V0uJEmFQ/NK0I3AEOmod2j1a
P3PV93hXbe61muhFcu22IELRBri9bGNen2GV8TBmWdeyADibRkT9ov/2Jvu9p5t/
2/bQe+1HvfcYx/JI2uQ8RaB3Z5u5pZDpJAEpZB51mcUPLyYnsV3XJYu/ag5SdkMh
BRDe/bu1Vn+HEbKEaLElV4eMxcR10sI1wm54LTeN9Kt/Pt2MlRNRJ9tym2p5e0Yl
r4pr7SJYjh+cN+ywQmaKlHgMhWGW9FTLv8BCKtZVKi+DopX3Y9Gjg4VRFJ6EI7mj
KEJLWGIXryzZF5F5IA5TkXj9vMwbJR8MKJ9n1NA5DXt2+nWnaSs5Fd4QwkTUmmbU
dXwAenhoI5CuaOxncP5pwjiEotACklcjB1d/QHAsQjpQFF7hPJqjx4ddoxilgcYr
OJW7yqixtCqtvSJZ8z9t5zeEIHs5zUiki+h07NsAn+7P/4ZW7Yh1PeHLRJjYN1a0
swSoW6+fKxTFMiUMvgnvGgaZJzcmcLPJ05INNv5hiar3rLEheQLdiYHCLTohzaO2
/XW6AKQGoNT0biprtm36vnKgeiHH7ltpWSpGaNS2UvdsaGgWpAjoApMZiSY+MD20
6loCeXFgAsE2liExUNMZ/Ens+XMgArKBjaQMQECbQHQoJIUhF3IGeZRDNCRbUlA2
7cYNCI5k0KTqNiXOE94O2z1VBsUyvXV7qsdn7dkuXmYFtLaX18KgD5gxccpjcdyg
wnePt8z+0nNcicSu/BLghNNn1f4zacOCqDpeS2t7fTvMrsdJ2h9Nr71dCZ4aLxMs
8KwypeGKSKTAyNuJRyNqAXUi6CScLLci382Um4hEI7uMPVchnsA4Ok9brfOlnZtE
4IhsTofo50H/84bIcCYY+39EzuM2NN8jFXER1mHoR8xfe5VYx6NydEt1l6eUzQ84
3dRn4B+cceIShW1rpOg5ANrY4B/ymDankzQg/0Jgd/EZyJem4/AlDCjRX4q8AM1g
H46ENhdDvENwRnB/5wbGuBg5/NAoMLNZ8oPe058/UJodgys24lTF/Q7hytrjHKFw
ednMX4jJbyyr3c5xeNJqekHDRxJaFY+tE33qCg0HSRXhJKR69K+T1qokMddZqQTz
v6l/A7PX0bcbNs9iddbCOtKHUoXEzNWPi3Rt/9V1MqZ2dpBM3ZrbtbxOMeIMURrV
X2VDQ4nyHwvce0dufZqywqEQStYk30OFzzTSP17VPO6k36uXrDkOnUXJtbYWvp6M
q5+5y+i+TGRork55K9pr5nQa9+GJufrqDDyxBI1407o0vVYYe2+DnbcP8agYTCMj
GKZ8Rb47//212kN20gdvy8irgCQ+IHbyk12q/ZCYUOfNXm9aJaO1hIAnxQOPXMhT
SeyFZ2VK/iuOaDRse/Wy9BzrXNs7VY1pI3ssd5zwaJuQSVKTQzI2GZAyP6tKGJ5O
o/9fECko/sMCXkoP6ouTE68ZB5wPWJXeI2LTUIBGkmcuD81UgKhpAJTHlqMHZJfY
GBdNFL8HQidQj06V9fO5QCooXlVHu/BXikb2Xfw6uuRIGeOg+hTMURtlN20KNKGs
EXlJehNc/TZNn0tz6rRPbSkU7TPUzG1ICHcK6IXf9fr9RDT4inBerI1oj6wRAuyn
DM72RDFPQxMMTlOWITtclMvyX5egNCWkzjKOjaF4c+SdJhaFP366uCAL/f3pXsSq
JTUjayzr8fk83VQ24NKUDo4JYfvPvtuKGa2gb3Rj42MgDwGkkhQPIqUWrHsqiYSq
L8D8PDJsVVfIDaPiEe23HmQtS/MfcA1WoJXea5Qc+IUBnvlT5M4duT2B12RTL98h
BabOAuMD334BbkKnJtSuGl4IIOV2rtrTt7NjjraBWZc5Yp7Ws9CTaKXq/Lnr1i9B
i8/A/USENrfDGmHlUrplc82joxll9Lks6Z7rBm5O12oCHV776cDQtUdRtioebm2P
HSi4vBL+140a471MZOzkm+VBfs0vHA5m8n1kHBiR01zDHcHAB/nEslISB1rVQ8RO
PJRJJkDnGKbNr9h3voZZKaitPO6h6Koa+nlYOERn5ZsCBwB50rhMzyAHQwfZgBG8
rJ6rycyO6sD7zSfFkew0RaS25QjOwjn+cn7m6SIxxkBvt1c4SUQmm1W8DRhqc6t9
rBwHi9+0ep94tqFmGpDeLrIwRweE5HPG603E+q0GInB3vf/9l8N8e6bmKJ4SbBz4
4JcJEV/BaGAnNaDbCsWdYVkE8E1Nbli1E5vtbWNC7D3eZWB3UCf2rqTKpQfBXSnE
x0tRrSQAzJZVQ79mbZSICI63oaL3AU1fGy5qDWHQOE1P4VSHdcrgnu1UVykK3SNc
ju4vdHu59PI60YrvhwdLNsbKbTChdB778CciKHrwRBz+/w1lWM8ECaSsbWtNe59t
tVG2GLDxHleIdkYemyWBaOkJ8DlsGFabuH6C5DQ6Wz71rXYnINLYGevcztWjA5Mo
/UFq7aG38Ub1CbOXW4akSeagUVEr6niyZQzkiytWrdCM6x9D4/JfuLy+0A9ZuGKv
/ofvMmLzUGa8H+ZqdR5eZTt+YQtiL7SbaX3oN8ujXfUr1sKVybC3Vqd+37CdD3TN
9HbvxtPH/4krUh2qttZTR/QEC95BGXqXrxj4F3O2AQUqXXSolxBH6Q+SHqAgqIAL
C012lSj+E3w89pijSJZ8fDO107vq9cJeUCnC0zTYu3S80yhb65MR4SBZkQ+x12Im
BQcPwUMgqLQV+MWijU9pEfo1JpOC6C6Kg5uxd6+3Dhql3gucZRDTIKZ1kIxKupYn
lJdIuHIuu1H8YIzNqerlKb6KvWCqvWkGfihVBUgdUujSUFJC5RC8cZas/Fhnbuhw
BqmtbPC9FPpuJGzcw7c4oow/fP/Q10MItBSQlQ4E6+J8MpzEIHdAonbuaSKbhiXu
IPja8smiITe4k9HRHQEQ4D3d+SKAxHQ9h2NMPHdwVYEhibdbT3akDLfVGfEMIxn4
2KACO042WxaXDTKxHPyX5KND7trCIpTPC6s997FtHpe1yWIbw3J5OEFuBpZEcf9z
xhwM6GyQ2iStoqCJ2By6VsSL3cc0/XX+Y9o8XF/CTxd/oiMKOUJETEs3ngBXIdPC
VRvIFtjCKsfyWtcg+1f2+s/+xBuz7vgJwq3s7pbMHAiL8ft/C+QQ+Fzue16lvG+2
TtDl0XyhhgDiV/Z33haxtCXIQZWznjkMFrk+qa8QSg6Ltdg2eZSb7n0BxU1ir+UE
nBYtdsDwkKgUhE0d84M44dOCok70PmfYxHsSlpn3Wohg374RDjMIeJ86rZb7vy8u
8mbIem127/QYxyLhCObjVhL58qz25RoAc25SzHDqYKSqL/+K11O4tauqoBTpXNkb
giOx8WWRl9eD7NEgE6jWcyj3gX9r9966NT5O3QcEqIW8ysiKcSrZP089l6dCFyVu
Ei4rZqd5183i+pseM+/hedSpd1059ariwDpoOTpDI2cagrjy5pH52+zvfXWRXzP2
UHBBe9FSB2c7tfbbX9HrTCbzJNNcBXcaqEJDAIzeGm5cHGnLeIAJh+Ps7+/DqgFl
W0pMvlvJvlQe50BxaFdtrB/vj5ldcD8jRGqP/iKv9qGyxFxvCwaT7zhnBGqv1YHg
86e/D5K/6ohGD+yLfWuymsW0JOaZtBOdC0s0dPWWRzJWC6FAmUhSWU/Re0ndRZ3W
tSuEHXKxO9r31eemBNuhB3ArOvbYG+ZBUXcFzt3qlRMLY4JkbVgLXDCVfvER0rPZ
+Bn7tGoTz/Oiq+7KG1elWzURcnZ2vms6ob+udBPyOprNOQnyhkjjaXzPCmLJnA1C
RMg8WOeSU0xfOlMqnzKVLmCvh3+ypw6R5aHYInW8BzVFd/iFAqaTPFNadrC0eGvD
TXM7xDGCiZyas0gpGKTvKqRk6z5BzbgL6oyDPuxiJw/SUOUzyZlZ7/Yk6GCmAE+1
5/Nw8NVGgtKnYTBOkxkohPtOBtIeH+iVL7rzQ75CKMYNegpXsiE3q+cyDIEuXzzN
AKTD6ipArYMb4MOUTbzi6aijKLWEDzp/E9J8Z8QFl0M4TUvwrli2xVm7Yjwbu8SB
4d8co+QJFosk4ZRy42IzRT8ZBpbycRZb22aeL/zKLg42uuq0PwRfp45S+z+jSjyW
cEp3U05zj3Ez3V0HM3uUJ5l07Yboa8CQIC1Mn92rKHUs00rX6DwKkl4r6w4FW1QC
JaSMQ2hDL49sesl1LDLTnfvL3UQe07c9EFvd3Tb1UrO0GT+01e6p63ADhsCGpIjQ
Zk04IsMumB6ls4u2uWd+sNaLhklcX0srNjxLSoiCrdrAYEp4RwH8q6FkvWOsmJtQ
AnLnzuul+Io0CYimjDSDRFF0y+Y02uZQcntOjjRaTkU1yyAOkb+c5uNemwTs9SV1
zIyDfgqKhaIXbd2hf53gBkEv1aNTVYWv0dHLkbmfPv4+OtkYkO0mmDqLUmMnxrga
9ElYov5FARg+CdNvlBJWkGYhLRlyeli1ugQQKfUqTl+BUZNouFNtQehnjTxG5NLg
ch+r4rFLWB6F8lfSBEsJypkJRfH38zvR8cTV2ruTZP+yimjG/4BKwb3uWvroIEfX
tC7jmLaa0cZv7z1DXtJKniey//lMWdDctCSfqe8JrIQ/Ssofstb7S+8zqn6O0gLQ
LuxQ0VbI6qURmTr4sBhMuxyDWjJjnuwQ3BS7zNE6krAsw5kTeGeyzA3yXSH5ln+W
FW7f8jSX3OTVsRY9ai/9r+qXQtvIS86Mha2YlxGdjRbZMWqwuyV7K61ZXEZHzWig
Un3t67KymAbBTVypKG7RO0SduLlbP6z7gqy2juUB6K2QCzyYDaYfxg4i7GeQK/TZ
ZpySut/rjOJetlcMBAPU4j8NfY7npoNk2Gy95s8Kdn/sv/Uafaaw8OP7J7Y/ldxw
VZtwp8OmVjJx3+cQQtd9eOGyyPNZLaetc/lQp27WyYLmusPc8+4MHPZUaD4wllyO
y+vTKBdDcMelw44QV/AP1Y2jfvqbINZMom+Ohjw6vRz/PkYMxdB38rRCUSLMa4cc
9Ru58h5GCVd81apTpzfl2ZEuo6JvmQOErcl9o+RXkyiWWmV53hHSKrqVy+hFpjUz
bXfsqQn852SU4JtOl64tnAKdtVAHXqHZxG+2QyYoEM2ZBht2sS/yXj9cEuRCaPv9
EUpOTvbAJO+j4ctJJKHxVshC/dnYtfbE/EzmYgHwjySnym8dm3RpNNUyKwlUq921
C5Bre3wwyWzZJ1IKodMrxgwCDqAmXSQqiJSTuJNGfQRopDUulUvQ8faXehzetJ5b
dZfAREyjOVnWGODUkvv3EdW4aLxA3TWnzbfLacLrPyIeV8xu1tpn000OugOrJllp
m5exGoCTUV5jAcewCL6OiPztahJKWkiGcXqEOXTOVsZLD6eNcQLJimWL1eWnBKBZ
ARXid5SJccaGb6ibJ+FpFnpVK8WSdy8gMSXJqCunjxdZDi5NGIz5ssuok6vc/5tv
Pb+UWCXZrQKnTHBZGD95wgPmqjVG5XF+HTy4Dc4z6SdfrESVeJEzm5c5oRVMfKaJ
6YSQex5DiMzBzPgOAww2ET1ufrYJ8kktttOiF1YaBoYXVUo5QFBLm74xExirXa3b
Er0mMPmbVXQtjaAJmxiJ8Xg1OXIUzQkeDuIY61TZjsswEbMQUIIRD9qeCSuhE/FM
u/lHf0W7jkW9WmtN7pWC3NjA9DSm2iT+UJ3PmJJJQqubM3aw5/jjvZRZo3FWcjHm
RpXM1Jz8zbWZchZTZqVbmxSd9Q+/VZwnHJaSFS4boxhe4l2d+yu7i5mQ0PmuejNZ
YkaVEY86qd8aTEiR/imn558pJuTBJrm5MHUkKrmwq31SWTTzSpLOdeSukQyRhQU0
U0PvGyPx3I4RCQgL2QuWhj8hb0jb9eCtDYDASixx+kUTLucb2pTI/oophWz5vqhh
tevFKTFZ+76VLuah5SQ1PlsdH2wlhWoEC6B3PGVf4Wx8DX546Nymfywu9j39O0Ec
4Xh8Px/N++//40mVrB0VYt2/4fRvvIuTDhoi8StyVS2CutWjgFPTjoW/pvsPGXbK
2oCluTyR+30p0+cvgPTPku6hG6oV9+dAPuid08O/WNJghnphyC9h0EDtdwpwi6sU
lKBrS+g+6AhDxhPxIvn9yRaQVEcoycgUr0ul6qic3TMJn7EcRwc2KUN1/eJi70In
GAg0qiSR/hmyAXAay77vOxivx9A6in6Tr1ogVJHZks6Y724oYasFKXhMrgAW/L1P
zMSebZ2s9Qpp4o5Cg2zKx1YfSinubv+Avc46QekyvX6UBvYcgNlCtShwuvcqH9JO
9NLnXehrQ6PcPATJcLtab8sZ+iueqbp+tYwCn0FXKlSkMXK3IDkBLO8GPpn12gIW
WBcjtT+PZWshK8dNDJ0BpZA9K46/LBIKDGVzEXUbJx40jqXZa947vxozxXL+Bh6a
v8bEuj4MqPZo3xqEbsDxhLfEdxl86vg3EbSykPzNn0BgmU7qqupGFHX2CSHEe3oc
d/WWWB989IVgecEz7b6MKiWCOaA7Kt2jWwcDFA+vBTuKGgvLtKp9edEVJHQaZdPu
AOzbt3XwXmk+g1uEKI3y4jnxdWsYLEMISW3wYj9AXeu+yXxeYPvBh0g+RWHqdw1n
QljuyxIvYMqYJvcSwhsO2Chs+0CTlBJRj4d0qniJKHRySi7exlZ/4ZXvSV6PqMMh
Edi9LllfWWWJ/PVYPZvw7srvHNdY36pUOWHyeycQrQilrpqXy/Bs874qwIctJV6v
7Oqhl6CLMBlCNZU0KF/3ucElj4jXbYvUk8UPhA7QUhIayoKkVLcGT0SkWTP8erFQ
RiYrbQi1iDYY+Z3zZccwHJ2/H3xOAXdwFdVnLnMsV/nieNLCOWqsP/VlHwgUQTb6
0Si/c8ooM82gFctdenHmkXgaEBaO7TJrRnPw/oF0LXL4+tvo3PuozdkiivN0XkCs
3zSvkzpzgCT9C6bl7bRPHDUyos/zOA2Uz893ONwkfY0ydbp4Qds+Zl1n5Aht+8P/
/M7wSKeysvxhsebRfPRVTpf1ERZfG2FE69ePYR+VdCdhgygiWaCGygljV/gD+EJI
gzFjjtPG3j4GWGySyd3+OoXycsPjCYoX3a4zwGT4t+OQP8BA+494gr3YkkJHujmM
MCC7XxHLcCrxX+VW1ICsQLE3z5EP1NCs9MREV+sM8LszEofV7rJBrbKXkQZjVL4b
eVAcjQfYSH0On1jEDWOcr05O5dRJcvGqi6IMTcCMykKGvm1tREY4TIYmAZSrCgcA
6ttPm1V2u7WnUxjUoZtxfMzEMKIQDz7q5I5Ippax00EMuNbRgg6BR/anonun37HR
0EXsqm5n7y5XiCO48TLwVb91P9S72xskWOOnwFDffUPs8JbdghLqfe89LC9Ofb/j
+zoWnTrixrDAYS2PhYkD+8+cQyGgj/kztBlxa0envZ74lWEgIdXAbRBnjvEkliba
VU4/e5MYwODkfM8zuXQ0E2MpAL2FYjA/MfXNEKsma2Dbw/pNSNBDNe28jMW3mEKM
wdT63+8/v+cLaJz7NUhVTmoEeaVu4gR/AeWEsCcxNfzJ9k2oZ0wuFotbdpBfD5vD
IBK2YlyCCzgnC0LUEzUqDt/TO+/ySEzxMG6YIT8WLOb8q2R3NEALiz2xjLmZgXw4
2Hlx0YhUJfbAq2a0r9gtFstXPqY5CUdDOThxg6LTEUdmKLxwwMKXvvLg4vXBvkcS
K+gUj6m15ILGno5G06wjhbmTtqYlra7v9WZhMgof46spTf5QRV7HNczOfuKPi9fX
q3VGwYQSBRlGBTvnpjkM9WUXJ5IDHSOC55aG4GUyw062LdeBgPw53K5m3EhrGZEk
HeF2AqeT2JI5Cd/KBAGyktbyYhDH0XzLSPJRqUHzkHm3CP7weDc4kZ7LECiWpoDV
uq2RObNu7CGECr4RwJs8hm0KGhV4SqNEHO84SdioxdIKmsm+Fw8sfozUUoAeuUlS
XPhxr7gB7iB+JrsVRskuoEFHwYGGw8w7syA1pUVJprF2880sPtd3Q0TwsF+WrLeF
snl3RNZ4uHct1MJmkAnMnsD4lrYJl81FftgeCmrPSjRoLUCk6tqM2HWIkznZ0yU4
JyocdrNsgbEYs3i96jLJaRR/+rIb6YsEH4J8n27b2+LVakWMyiY18S+2e+ytsypZ
ORb1ztw0yz5clKI1jwj1g5aszUY0q/4hdsGLD36qA83nIpnYF+mgsugCZ+ipEEfT
IKNSZsTNiWg5AG43Y3JoGzLcWi8tLIdEFnIqPglamHaMUHLL9O/UMoktaWTrz1U1
9OWhgQphFjq4Osf+dDu0NEVD0Yg/J8CswI4PVlcBKw9LQC7xblNMbgkE3CP8csoz
XfFMBLJcnOIz5KR5+lQ7AxfcGrVn4bIDaezxIngoMxgjvKT9+X7TD3C1IjRVdEWV
XJ1mKY3XwYQOzWjFoF60a4BRbE0XklK6iXUoaJdp3D4NhUJVh/rJvzJvJi0v0/2u
XUI1E8iIFZdkXdUw0CykECk1S2sYCbOkZ8n/NcocF1mFy/YSwuQsl2KJLQQH+7lw
BIm4e7umognqonkGWwHIC51qKZUP4+yR+xn1YjM97bYXU5o9eDpsSFjx1gA8zH7L
Xpp6sky3wz/DgVfrlGzv06knq4NZeWDvMsvHeuSCetCWGgXsUhilkCAb7lqJrs5z
YrSuZv9XRCS/MrPV6FvjsE7ovccBVqIaBcJf4tMavnBEOJVnHkYBrl/f5fvqHErN
ea709J+QWgHKsY3TOaWDq6SgkD0Fb9LPOVfmilvfQHjYxuncKRhmknjwonHFMVRt
lYTg9gowCKgXDnOm9sMDMMOLasDNVMFNbD0kyiZzHfKrbI0zKzdCLcvqip4+LUL+
ktRdV2BaUyObP5RWuA9FV93OVOziDiv2YTAEZ/LBiWOmeDHeHFJtsEQ2ISSvzX+V
9quxM1o9HBNymqFRkLe3gCqwgCrLJFUux33fuQ+EZfvW8PHgSEBebNqq4O+ISb8t
aOIhEDuOxeorbbxdguMdCTpNoIHKVRfLaiaJrw22b2u7xtT7wSdMRoofq1yNvbxW
Jb7gnC++Lef5ywp3fylh1KduaxqQDUIrMPfzzKQjkxVGdsdosGzCy5Ba+bjB1EvD
Ha6X8EtNG25SBXov7z66B4OynNo+OUMowGyMfWBqGiY/pOcN7N6MFGveYSBh2cEq
lRZgXOI8hPH9ai7HE0h5PF3jX51XaS+XQ3Q8WUvhhF1i2JKrcp0af0JFjcDP8F+z
+UXlpwE2/pxGN4olBPfjp9ip++dSiKehpxZhlxoHUHiVRiovbwqrIRGUu/5sYh2O
zQsC0baB6+vkLfpRZXvBtf7Q/ifOaleQS2hHdCbcU4lXowk7s2B6qNIPHxGOI60N
65WPxhm1aMY+MU2BmTVY9KBWDkZCE3A3Kd9BQKASY/p4UQzDiEO9uiAcnkolYCQ8
/93O5KSXMhzirbWeLltpGOGT24n2Uztr3dPFtsN3Z3VtrduY6YabFeGC4E+tVCew
jLvgdKIzIOl72S0jNiBknBmatXopShsxjA3wvgiiQlluZO/LaZt4xjCpWVRKrm5L
DLFscNtL28vEXZn5muhSJupWT3QzmF0HW9fArxhwxCrqFH0AF+ARQjGx2LKOldaq
Nx9x17j10CZv4hr6jZsGYmqKH9urYrWsoGhWVBfgBGXB276762yhSErgjLwjgbwE
MtrA0RDmGMEtWXq/SrXHjzXQ4NbcGJIKO6N8ZL+QnGvSG4W794U7XsmGaRJlqA54
gte0S+rQpZOAi3S2P7vn/cZzApX1+iaY81RGiYUeIiy8kGbdGoeu6Q1FX3RFsEO+
5CMcBpMlWpvSLJ4847+kHWk0s+kzxPKQpEHKS3jVdHNd4BlLra+IMyZ60vT1W7Qi
A22PNeZ3aYikVb3eegPuLawXJgbNaN7Rhvp+iOFh9Xz3PiYUfJIeeKQonJHEI0/h
AMcUikkUPwZQ51P862dvnjskRxfAhRrWhMNhC6wEz8ANGxT4+D90FI0RVqyKNY6e
Vp1SnrheOgjgRl39dZ4INOSxyCveT29VR8BjR5Fz9KaXrIrdZ2Bog+caGl4M7AEE
X4269krBsyRZiFt0RJUHbBi48Hny5K2MnePotYOS+j5g2aFRRUrtZ+ikoyTMLuxs
AJADzk8DZxPYt6wggZij8RcyyILFoNdYFS7/d5FfRgDQruMj1gqMTGljpf277ZfI
rW2iUqky+6E0ylgiujeDyMruFDKYStTPCZLZcCF8JE80wTs8qtXt5u1xAkuw8EVi
aDQSvFht2ArSCBC2pYxTWoxMR5paUvkt28wyRXuzaU+tNUFXLejy4diYc0ifaMTL
kTWFkUqfMTsL7bOysoMN6sMtwUFSIQs/Sp8ZK/9xGzEN4vvGhouLcKb+rT9ajF5C
0SvoB6Vo8R/esnvRWrqYPXakpLAmv2r+aOjnYW8+NXNn2k1hJMmsAG2Uz1KqULRI
NHcmJxEnme3TdaLb7ppR3KOR2ufO5Tr9MYo3k7BFIjR6KlPoafaRsTv5OYdSlZu4
J9HMggN1Pgj7i/CrAZcOzty7uG8Qi4LoRnIVBVL1E0Xg6NZEriQUHEu32DXefm1l
JsE8XXL8s1RjZeRqURrhVkaCOazoSbtuHqZNNoloonAg5hjYZ7GkBLIGq3MpczYV
QvTAeGfdV/x+Whz56LlqfbEsKmG8Jnfa9dwn8Pxhg5i3R8FFVmfaffOdHTdI3S2u
SW57zGs6RQfm/F5Q5D5hmDIOBIGUDRB9A6ErxNhGGn+XFrEFsqOvGrTzHA10blDw
XTGrNVhEchRyumRVJXzvo6/3/kko3kPkBLH138eRWTgUaURY+9Ht6LWnp37ht+cu
oxviCtBpqvoZSflUCCP6pV1BzF+nGeilOQOwfbkanicAogsilKYVuupNGmtmbnZm
FaVLLNvwM5lW2E9Dfc85qPKP1oQkGfLJ7g64eYdGeSQvj2u9DdguWvSUbr6wJXJY
rw+caNgEUVOP1yNc8DPbvWEn0Oie7huU7b1zce0IwI1Cr1JwpiXl8hYOvf/V90eq
1n4TyAnamkdTJSZZZOx+ysiRkN7DZJ6bR46x1cQVF7yhhMLkJXp5t2xKiqvtME5X
Yyg08UvgUU9HIowuscQXRNfvz3xudozvimVyTZh6tdDX6vOzAKxk+ZlPHkWsmvhN
lbWHPe/L1ntBBOzv46NSfSnUlwMzYrHqet0RA2YAyGTklNZjzNKkm+fTAhl/6f3l
bnEEK5hgPqZT+L8P0UWMYEovYlP/J+nUWBJc3M0giDgXqYm0oh0RcAYkA2aXgzhU
INm1YFTA2s9WTXTDSDRyel3xnfDcXROrxNX70+8zB7x+VLjCvNxFjav8ICRmUtWN
xqBm+wf6QpF/IYtcyLTv1z8QGcO40wqchccfkua1CUitZ/dR+uYDLfHQJluh5oKC
P2s0ek8oHFdSSgBTroSlnrVHtK5C0A8tw3LEgewQ2IbTlNp2pOQi73kPqsYGpTBD
VL7vxSJDAvPTn2wIGaRVfVyo8M6ofO6QrzDqH9IQVxWGEVnBtzNvonHhR7KWY/8i
ZkRS3X99H4cn/NHJKtYMxCgwDCYqhsghB2EPo4W6K9WVwt4oGZSi4faf+SLDucIF
0tkwGbr0LhAeJlC7TdQkhzklC9SZLDxZzyOcOeJdkNbm/M5ulkG5GtWEb/Vcn/kZ
F4JJATe+7kgKxMeqxbrxn+3RRRxJaE+JNGohU94aS3t2PQlCkue3tKCt4fNNssTd
h4fbNNfda7B4RrVPjKDd3qkL3rZobz5SVtjdf/Dy3wnXET6qqv7uQjscsM7brO2x
LdzD2MqY2bhOAhdvBkffp8+Q8U8I06HBU59kqSViUqdsbz1yC2iAiC7jwL9uK6RK
FHt7xi9/AQ5UUGqvLb248ezbAQOe373iQLL5G/R4khokBZ+Malh9SuRc8drCbdU4
MQkOkLx/9t0+jeaMMUxI7dIc3/8Lr4QN3oxICSs8kJHhVLwlHdahoVBN/RotB8Us
5K52KY2CbW39b1TqdZWFuNCJx5M0cv76lWGlkVd4nw9LCnjmsOzwoPkIWeSHOKKG
76pmEU3QOFyCI5WhVJWr+SSy/i75LA8VwPR3StjWs2i5cduAdsooeRlGwRWSMohh
bANipVwQIemgRRUtZaICLxhWu7dOzwaKKrD01IalS7ldaskxz47ogf9u307sY4pW
HHCT/hlr+S+n99YlDIRPOjYYhObBEDXR8Ou6PWvFQD52uVDFLL2KbYK07/Skcpr4
B0y9jGRseQV8aCw4G9mCN+60GKxXWP0wEKcaGKWVp9AcM38dh1WBu6a7c2VwJVmH
3qokfHRpZlgueJk2HRIsaYI0OtymMDQPV0nC3IGSA0MetxBgHb6ETGJUPvsM4Zfo
EnfU1xenzVypmCOqPHJRhRXOZtfsaz9XX9YGfeILOooOz6i5HPDSIQV+g+lwtiIH
IbBA1n2erWjQ67W9/IF2qgdye19BEj/nPDosgzTV4fTt3n7JIBN0IbFsCp6rSp4p
YtRiEmPO1GkxaLl1ePi4VplAEmhw1DEyNPgCInWRuna5HNuxMdW4FEA9haqR1NFy
b2K/0zXnk6ewmVgdYlxwEiOAomyhV+wbHmk7Iy3u1spqbZx0j6zfzbqcB1rWlmlX
ubiimyInfR3SDfTDbl76UxZXovU8uqPM2Ly7Gv+XkMN2jhCiOdOrOZr/2i1YtkX0
CznVOmw4ff0uDdDM4V1mzPD4cruYOO9U/LfjXjrGuUdH8NdRNHfge+17RpVoQ9p9
EKBYzMnjRj6CaMLk97L1gz+jHVjidoe+Hl8rhwtmVTaDuQqUzClCxed8QQK9akeZ
BkIWgUScL3V9lRUYHBtf1jzI6eGlZNEAsK/1eXAzwOVerybEavoe32J98B9B4FMI
ldlTER2KjsITKJNRx2otvCfZcoPy83O6jZVDKytVcqEGifUCbQR7nIXofB8VkW77
koWMzxgri+W6SfOb0OYDmgOLvtYxqhRkO6kCf/ERkuBTAMhi/2zCR+n3ohWyiqDA
G123tNt+95naX5gmU8z5DxboCuMr2ySkKX3eMS011rA9UMNMEsKPb0anAB27vnqE
whVLN9hr80EsLbCud8BqDrxZ5pEg1u3CLdRti+F/fpzjrnq9fwJ1dbyCvgLVrwpX
zNTls+Dfn+1EV+dddo0/WTuHtjBpBlNMabVEre16Z4V8qd1JXNaruAkCWw367VCJ
9VE4AZwrrguBGNVwB9fWHZabK74r1/rQwQCxwa9NJZy6AVSdh79ZNU6vIe0OVWOZ
c7NXx9D8DZF5cFVG/h322j071RijgM3phaFvGvigibc2efRTaTgyc3IqI0m5wzGZ
1DdZ5NJeaxzW6qsl1i1+DOahaTEPckQyizSCnUPY4CMKdCimhPywvQlKef3wIcgW
BIrpvRcPUtVmwhBrWtM17/CgH/h5zbpj8vJjD5J+cP/Y+HfmOUF3ieNX3sgBXKxj
FOIL3fHwarzY4jvt8cWVCjhSFgd1Gnfa9nHqFr5aiqOBRqsd6hWNh0Qq5xUKibcj
MPez72GxaxFc2kmwZFr6oJa7grqcduTUaLeCpg6hBE55tu9lRER8BlgfUjwxdVYy
ue7UKcHO6N54yW1aFyfkbOjA9ghRTuEDL743F9Nq5LmgHARJLYEnBnBCzpMsFf/U
mVP0ticRrG4pSaZDUie+ZrOfqsU7SBBTZqOekIl92fcQvqlR+ngyrtsUvSaTVq2Z
jA1mVYYrEW0t41NlV+E+MJjVsDfF+Nh1v89dBXA0xZtX7dLkaXOhYpcpRQ8vMHtH
cdH6S7OutaQ+RltEhqfuaSTllr9RdmxeeSzZ9Yurz/XyPX6PjNn7rxbSPZplbE47
A/4FKxWu7jBWAM1l6ciTFA7h8CjFo8rZXPhzysqOGFdPIrh06DupBsyMdQh3q3/2
gmi3uJyBqy6B9xyOFWpiaspYVUdjcqt9NjLtQ/19TDc=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
XjZBMfaJgrK0Tc1Ubesgb4ZTrs0UiEyujx5WS0Pt9TlAYOuvNzeoGjikt3xoDNfE
wMT6SqSn5JHQDiE4wUBFPFQRBQ7OZQP0lyq1sVE1HgMEb/8G7rKEtcyfSekalY76
a+3uA8N1/DlZytlf36zQNaxSTJpnaJNXnxxKARXz0vR3VZhPLltIPkNFVQt5uz3I
J5zgC7KJO9QeInkvErzmcVIorcb/vI/RVzQrI4LKQzS2j4n7Wygv5SG8Yq75sMFq
VaCw1J8NLbCqXx2ZKWUAomSizx3BSFpp3k0kAXbq2W9k0l3egFIYX3BO0RYfkcAg
Iot8JW6LG7dIy+rnlryFRg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7632 )
`pragma protect data_block
djVGWR0F8yfHcKIRgGlJnm/X3swCM2pFvlcXDXzQ3tD+HpiEF7nTcSC5Ug0MkYH2
JYGlGjWfLYa0AE3Xl38j4c0yfTHDFjtwgmkOGjV/fJElKyhmL417N/fpNwB06iVk
PqWIspO3qvBAsnHEW/taXPwEh2rYV0L+sl3SN7+DemYVQ3VqLJQEuL6oEsrTW9tz
1qX7EG1AEZ0A9T8pyu/C8mopwgwEsbRY4cUkQzzp0InsaIXa0StQGbfM2tr3s0UY
fWKWfrnk16w9Fw7XyiCTN7nBC1GKBEEyri0x4FEd38XnzhdalURPUvJc2cWrFI5K
8ANyzTUNfU0GHsFu9T/EnZGz3y8ogq2sQsv+a59FET8AupJlpFaGo9eBQzgrJLwK
JPL1dgi9E9PoeMIm63CEkXligwJDZJgh/1NiNz1I6WcW70znQoyCGvSO4Cwa2H3l
586Rqt+aWED7F8Jn4gKctHNAnyVWuxXhYqibEw2UL1HXgQPzxJB0VPfBtSToAb4d
2s4PIuulb/OHtvHFR90jEdJheXHvmtzsZWHLjM7/rAWaUMO1LjFeuAnqI+tzyJzC
Nig0jtIBUJTNdOPM3jErrR/AtDZRDq19qZUO5CH1uSHv/Kg05uPSU712tS/QUHJi
mmXxkY7yMJA5zLBLiofcs4NqgnfaKT3sJ9lFg7so65uNCfRAYxyNlaQY+0+xNCHW
eP+4Upd5Bl8At1/etBkpcUDQc1b9xrrxBvftSH+UrqP5+QDt5uRKjFT1vEYU6rhK
vnMmbGIkivdpYiKZmfbfqJJVFpHsCG8YpK8zc3LRLPCK+3+hXMkhkCH+hL8LePor
ZBVNqycizbLb1unTRQpZho3AhAAky91CnTjj8XKzj9BTf+wd68/Igw6R9/ysCufO
xZant53QLAYfS6gMNw2znjpKfMEy3rz/+kwAECa4WOPnCMxzNmG9GJYptnHhGD7M
CmER0H68I/wq8/O8XPZBKQBOvnKkM36tq/pVJ1+36dBwF5vwxibHQZG6EQ9pd19R
UMpSxgQuTabwkQ9XQ5HmBWz47GoscfSac/8IYcWKqKx2fMxdmgKkELVuUVILm6b0
gkO7vVJOJwAhc5vIaMv/sl4sPCUDw8ROYRdKzr2kAy2ss6L0M4UwWLaid+fuYdit
oEePDksgbzQp9wBUDjTwdUBP8JCCyX91qsG6MowaeLxKL2M4f2H+aGWe2cdULyh+
OKqItEf90rjy3xtpr/9LXJ/JaqwfUKmh+fs9AaVxCXxQXZ3bXeXQuNV+2DCHfjIM
9QqWYlo0nFLGVix8bfDlOf2Os4HgG0Eei+eF+8kEIL8SWSR22IZc4UQcmAn0hLnR
7Ipy1xAObisP/eO8PlrOvjhD3CoRc+WUdFR4HyPp5H5mNOBu6BoS6DUVkVxdEFWk
bZ7lMeE1YuV1HNVcgtN63y0vF5yFlBH3aI+thKuuQWv6W1PRHz/MNSDkKMcrBdTV
YNVSJoKYVqWEpssA8CujnIsYP+EdJBM1jMfjmgQ/v4s0vvKIZle2NH/71+R17lHO
r/fwabjpybV4Gw0B7NJ4lMkpHLDU++WF+frk3rKGwkTRTwVaFREJqzumF3waIPjs
uyNvWTKvT+hilseLjae60EHJcWAND5wyBZIjmbSqgw6tVf1FB1bvq5jk92P0ywHB
yjGdu/O27tKlFsotVOPOJW2wIhBrWekdJoZ5+bpkR/qYwY7euSF0eQQbom9/qgeZ
jKVQ0IubtnyugVwoW9jMnPdjBoGB5i1TURFOSoSup2rB4bmNH3kZBkeGD0/y8I6y
JvhOrsUAs94jdUuR58DM5GSBWIXZOA6bN/GXV+jw5giIHA5aaot0eTVrMKGxvO/p
Nq53GLoiZ+KFXUVShEzzAR+2FjWyc4epEqQUT9tj6SiE3KUw663QUdqsHrQiQa5O
zEfEsGEBgtztbTc7+TaxRE9BQY6YRFF2cyoWiXrGkRZXadUV9ko2Hq8ocB5963xX
nPoidwdw/JakBTfQxqDAVj3pV5bye0/ds1MgX+GjldkKa/BT+5IOgZE18X6fiJw4
LltHe+mSmxX6LhNy7ViTBqcfOBzz8xhAt9tsQ+bWqPIObjtYuucy66lyHzXPlkRB
yjsaNX4Fgxb4aXlJjFu/Gj1zQrCUELYev8gPUD25W0XahORt26mhcF/6xpYmbFOe
/I2VpmEHk4v3af11DfP+2yzvb0SI6XuOBS50IiDj2t7Tyn0mOhCOV9e6p95Rx/AY
xL8kkXXgbuibGjddI0b64a3BddF+Q45/9zPZugcpB/6lEt5J7AG4vY3C1aBhErqR
WZ4t/oIAdHUn/liYqG7xInlNCvIukz+LiKi8XakPjFWcWY/4XhO9ECi2OfftwJPp
tyvXp4mw8y2rtuFW3pAMmtheeKaIwkUAa+7iuhZ9zvtN0VE2ep7aYfWVBISApupM
Q1LFneS9nTtVisPBoiDHo4qT/coTnpJLy4g+Wpsg+IhXKuPOU0i3RzmcfAlOUFZ0
wZ6Hf98zLoTKjtiW6ei4ePXeMAxdEq7AGLinx9nRFC3JWy1yFxD6mvYy09dIXf8N
Ivf7coDnRu6tk0aXB61YqR1wUwKAEqOLDK4MtLuaorrFsP+sOhpjOeXoRX9pH879
0UuWZHL+tqSyzJ+YP3J1/QgmZ3gg03/AMsge+bOZB1KXKGJHpN0PzxE+VgILnzEj
DCJ06T+Vq0oHZLeECleRcIKbx+c9RDqc9dLfcrwLvdjkY/74kMfomzcQhgnkJsTN
iN1xgJlE60Lv/Q+raVT1GzGRJnwoTnQ6Cr2oEk53GSMfdDj63Yx+8D5u9C9AA9jX
0G5gSolK7N0m6W0GSqeWOWCAmA6T0+gLlFKrl6b3SmpYROoY69UZhYYn4wPn9OP8
UvYPCo/1qzpM4RQX8n+mZ6Ug2ucqivgE1JrpZRhykRrbnWZ5vgCrY5V3XDvoGQ2A
Ye1SEX9Ilmcn0IAmMYqBWztoIo4oS+VgUK+gtsswXRxlg1ISiGyrzeB/0He7paHn
5IlGA/jDaiROTx+AQUOmXQf1gfUC34FCbWyOaFriuxCFJy7dAv4Bb6+pHHPEpCTR
D+a1U9mbu8PSklNOg/n1UufKVWZ2KC9BQNtvqgIX3hn1O14leg3+mSfgPZuwGct3
uW61jcO4tdS7Zh6mqxs0BYiqo4E+GqAINjKBB5B7+gekJr+pvFhAjpRF7yA2bxnG
Kexy+aIOywLXxQr5DkwiUuS6WpMy9ZSwsCxWMSAwYLn5v2gPPnXU3n3LFTQtUg+R
5Ib8GwcQHPjQsyu0q210+TBQxEdhKzsl1YbzUAcofME5HMsboGDO26nLReMjYwc3
zfyuMqaWXajDLeadDQ+A3EVzRXl63lSBA+kPRMle0x+iYOuo4r3qEwQ2iWCNPrgY
BydcBNUJ62lFyGtHc2Rd7itdxjMVnSB3OA/NSbTza9qwIiUKrrkpz02i0m66dLYs
KE/Lw5IUxUZwoNxQTuawr8i5QHVuICOdQ0oMcZsGc5UAfaVnPNkHiPiRMoojVbKm
3nyPQyxbyo6vP07/RqMLNi9frsmwsvAmUIxb9EAx/EfYjwY2nTn7HlBCytrSAX7v
Nvu9Q1lrrYWM5M3w8xRIdT1PQPk13CSZoSXFK8lsYUc6t1xIKfW6nNiikj34XI/v
VpLn4c0qcq/4cZEJTzj8IwYY3qh+EWf5zbJ4T3NWCf5yXw84hH0yOsIUrJZUxwI+
xjYsQfgkovLzIV+3vm4K6Kd7/YdjPde4ANb6IaVewc5SORmmgcj0nStuUcrnz4yd
giungCadM3dkjGgWqv+JU0aDS76gE2ceCMDwDCCa3CE9bLdmLjxSRjRHkGxpWzSd
STAzGQDj3CS0Vy13B/q+oeodD21PeL+dWmjcMrGRSaokHIn5CIfbyxabEYUF0nqZ
nzknEhzA7OJu3/yPBpk8yiQhoV6ZMrYZZ9YvzgsB996ung1xjs/reX+EI/HNs6fH
e4OCtRh4uvbSs0ooR9ugnLyCmlM2I/icPrNhfFE4RYIFrt1nVIm6+wEw2vuQY/p7
1ZJf1cQoCrePfkkyrjkL8psgLwt2VY2ypjJa2GZAj5m+L79J/njHqy/ZJBftcrD9
+smf3/EGEn9fcbCuJEIr6Op1kKFEM3HQguHoMIFJUh4k5zg6qzAUa0gnKsNf/qCS
VGcQEMnSVE8a/QLjpbKyM0jZcIDhTdISMrOZEbUTCI4dOmUeHcJd2p3W4iIFFzSD
H+uUDUsZCQK5D6xHLQJ4TRqH2JBG3bI1nO2+h4PjmYPADfixyfq2Xn/6rLkmCJTE
waJIoCWj+4dy96ti9EHKV82eVLYkoDs0pC+iRii8UHlKGUOyrXpd5tA0jZ74b852
UCrJsV/oDarCoHoRSCBmx6H5Tm4jwR/GbYGbYR7ghYP6N9KfWJ+hYtvVE/I5ai9T
W3yFvsuTSaxlGC3MnzpCmaib1MGVMXYDtvsN59VJLpjD/pmxCtYcDSi684ep+OkG
l4ki61TrV3wMSjli/HLiSpNdARLK9VaqZdnTCrgsPq9MTjN7hrR4EGOTHOvGPgCg
GOL7VNJYgWFhEYN2AfnTUGLkuPBCNP8KfraJLoAFpQdI+o932MVXcSkZgvUQKT1u
PQjNzFsKxNcMG8aPkrIqy2qCfN1WqqginLx9tdbmcmFaQ/Bj+n6/j7MfmLZECylG
1kpqiSIhcobWrylnipLXpG4iOaY29jKQ4FcdFbABIqVm/XPpN3kbZ9DU7AsRn4ql
ApxwJPbcgVSm4G95QroILBKztrOr61sVoGjJ+YYwXUCaQDt9MNdx4ramosDCuZWb
fmrNxeuQ9BsgChgMaKpRy5jVQc15bbfX79pNddCpXsrOmXvRbr0UAYnMa4CJcq4I
snPPXvUAFBMnFFqMUkHlsU6+cl8jWXoRkygU/+GYJcDniyl/V8TKOlmJdErCHnj9
KkHfGotV05+8ejcxI8MoO3wPeQ0niB40Wb4jXzWGBvNCS1cUXS2yrEQcUcHQQczy
qELNUTKCUpBzDnvvRx4BojefQkAKKv4lYEydAx2yGiJ6Ole39XHG2lzOYeFfjKSB
UDLt7K+HsZjBSaKTDSvcHYvqJIaWKxB3EjIbN9ly1qIImz3CVihj5HNKG/k4y/kN
pzhFNsU6g4BnmdZKWHPMo+WS92vETEMm81jD66jkPYpAMAfHvczW59nNSWe9JCvi
tsG03IZ4evx0hz2Y7thtMeyDlVT7awricKUlFYZbE8dGeaHKs6KVLa7IxqJ8gp7d
ir563Jkd3wMymLRYPMV6cCHPVTCov/erUAm4byS83lH3vzZVJMFHcPV+TM3AcR4o
5jhU967fKIF6Vbs+F9Bj3Rk6nELsm720ITaqSyaXaTBYuzX0AsUCD4CNlnpFKTyH
PMrnsoHRDQ00ye/8uMiARo6uZM2zorT5dDE1M/0nQvUrB4y/6vmgqpe/g4rUTX25
CGn/txNlddGokuuuVD50daYEg0wQjm3XMQP6SSOE8UCsG8SLVEr0Ia2XVScfrEcz
gKRYWXdBm9bHW6NN7jvIZEAOUz0aboMPD8vSrWzLilkNMPhkdxEhzNgjVoEhoAsx
4jntTykVw5eltWS3c98svxliBjoMbQWegJY9Dc9BJ949piiVAZOLQGcoBklwQxrh
tE1EUd74AdAEvfUR14on9gwdquR/2FT5GnDVPRAOFi5ckejvYHYBL+jaaOajwPHj
PaDocxnOwsegDyvBK8iRf4/xRUZ7lKSdYClNr01rSTCCsSj3G6kcHiM80VRpgPWj
WN+rC2BGYI9tzFBo3BdmUxtVhsgX79xyDGskMIvgLqGp8eEiraGsiO1Ff7UNbIQ3
dbvPWAtS/j+RZf8vlj9tnbSXmBJRM9HTmEVe8k9IGITZDHuYMa/YWnVl0hN94WM5
x4jz0T9dqjItxeziRQiZjnGI5sbuLv1TR2P4RmuYrq6J2gQy41dCHM12FV6PlOKd
UbWhHXZhnm1nGNGl7csH2cSkIz/WYQVZ6bmJp3tl08wtfaRMsPi3k1mihJ+ETkNM
qWeo8V28JkGrzMLVXnbR+RUyH2zdjPw2kPkvMuRG6ChyTYyOVN/1ZRQf3ASFzoaC
u9/nAu7b9Z+bCftGTPyLZ2UApTUvAywjexD4ygJA7YKsfK4AqWOPuuJr7lhWX2TU
d1uvoNSr868aiyvaChwiHAJWAe6Lp2uPSzcvt5xz4pC7RQdD8xyno7v+VisNql1K
lgy+all82eW7SdUfvcNBVxnlAsYxMyPT9PB0xVOxI4Izq5S1wxvcZdQPPbehHs3h
HKo3gnMHSk2sfOHptNWXRrownvZRbyokUbZL1YTwMyqSXUjunoF7oYdlcPDdVh59
Kvq6T0MHqsHq6VuRQuqniE92RPHK52cKc7QY8Qfa7IevZ66J+ynNS3rPUDHsuZrl
Yk8vNMgqyVVx0fx+B2LDD/xRPHt0soGEfdcjNUAN0r9L8vvlMwul7Te4FX00Z1BX
ABXz0b07iET2koti8uGJ8I9TlHKuZRvF/DNfU1+p5kfVw5NL1xPm+2rhoeMJp/zn
cqpCKnHtzSDljrG/TzpXQPocQpF/vHiE3OOsbExhWJX4dn4QU57oLmjls8/k3TBx
NLn34QRe9xYj40rzU/LQVDqiqv07Q0+ZDnP+pQt3VPSQ2sqj0suun2bK/1Vv61Sv
SS8y5MEO3z4R7W1YfDtf7tmFermK5p5e6aVEwu4UfsXbPgVme5bGkKMV+O9Kg+J/
uGXoPLbgZ7Zr0401STX2ieu6QOCvrhmFAtbhU6v5/QM7UTxFB99xhDxr/SRnvDzl
lhjCFxJAQ6wmNDvrDMcqJmVLhQj3uaDHVUZjzlHKRq6KDNdmg3T802UHYvLYz1yQ
1E8O4ufqfR/tmocsw+4CFBNqQYcTsOos3cKGRGXw1vbD6zWHsnNovEmKIGtu8yEV
FxrBrPIDSD5tRYO/o/2SjfPtObsgHs4IRRNNTdgFX7Y/yiBOuSVwzlrFnjIIgkuQ
/BfELHGLSeM+l3izGeZ4lOv6bWDJ3imQPCkkadsE+2rQL98q+9yaVlpza19xIDbb
w3oS3wO+7jqW3ssqGngoHdTH0GIZsqlnrr8a+xn5qXx463f2T7cgx1wlICIYtGXV
f+TE7GBH/VIZa9d/YD0TQgbSLo0jvA8bckrco8Iz2t+gDujw8KUf9Enaiun48wDq
+/5TFDt+W/KGrM3ocB2rSVIh0oxB6/7fLpBwCV51pHjJlEMVHQH6KS6DRYESpuBF
aVnCuP9MCYcHC72/0czZQY9gsn5cnVG9k7SDPWbsHmZ3O/FnENeOyvXZvodxOUqu
zvdi1ra1OE+Hllt4vYLL0IuRJnGA+dfywJGZtwfaq7ssnf/oH2EC+lWhkRKcrGhk
g0BP8zBTXFDiIOrXbBHL/3KhsA4QGFMVhRkFRZiEo8wYgDNj238+vsa3RM2y5Gq4
kSM0TCmoThPSin1LSJ3WD6hYMqIhUVBUz0ZxONX8mGFf9Eg2lfUPNlbwrJ5mCvDi
2Zz6ri6kbnTpvNlR+8K8gsfMya5VleYG58Xgasl8g6Tg0dniRI61oK51Dprs7epm
B7NrGSsgDuOBie4Tjf3YiRM/hQWql4gn7KwKodGaUEJNds7nFOEsYqNTLti+iu5E
gBpBjFMDkpOdKg4zvOWpfKRX3sCLRm2VkzPDYNrSpWlHunS9bGnklhW1J8EaDhhx
zhr13hVjvmEqYpjcotKVwH5fiDNFYifBQd4Ak1c7ufWzKNzMr6z/TjfjLYbgU16l
HZvgPgKbugHEjSkcnBYNRaOvLls8B3Uj3Q+Rlmnhlgj5gDF3lkQ0knCf8pOIA61a
wEM6nSAM3wj+M99PV3T/pNzeBWHYpG5a+GpOJfe3A6XKE9Cf+ZO1EmwB/sXn5aPm
eLmqShClqoUPfHXXUb3/y2JhOc90h6to5uoFTsAEAzYu0TzcSMVOxZkBLl7RP1w3
mz9/IXMRCi7ZFqBuHVL89E4tAf6084IjzybG50oA+X7KE68F235lBf3dCCGgmLSs
oHkxUbZ6fWsYtZFyS9gTQGYa3RRy/+QUwNN2abzd8dttWUU9c8mwvZSaQ+9WEWZM
2NrVJKc/GcuN1vdNpMievZVvAXR+WxwAsN3/6qvQ8WF061V1pdd2KKExZ18pK1qj
kY/QephJXE2wDt0XXS16tauxUcrq+1F2VihNKqxt3RtiVJUJQCrp8mL8xtHJ0jjz
dA3NYBJp44l0cjAp+p6dZ/15aZ31pENRJozgCvzUdH18aLaU46AiP3NSqgKD124V
22p7PDPVLS8UpYmoZk1JKWW7vyRYDAUVxlI8GQV+MQme2lbdueq645WaCfSBMbBq
ciITyLz5yCs91umvzmdZm23PMFUKvZJEEpCL5GyhMKhc7RumTn2ByQ7yIUL2n+iY
0w4GOUKeNOjDQhnBZeFFLUEIjXnrtX3eNzsAI29gtpIMG90UgU1rJ7wgYfMF9C2a
jGZeVEYU9W7usQxAsVjIryEBUqfj20XjH6agfmcNBubS+RjoeK6mVOLhMW+ng758
m05AXOEOmZfp6YYCt7nU4OHV9de8B5v7sS8qAjgVfR1tTHpWJeMeapDrBR0vYaMW
PSEvyVoDrgDJdOIEH4tE1kpKMylQSgLNSYMfJGb1ujBQXdeFLeLoP569z1IoxAIe
ldXX9xqngPPwqc6SPSKRphkqDBJsGXFBCynasPgj+WVbR6sEalrpoDTov99WWT3U
KmeOuw6J/kx+HcaOyg3KgUWSEa++dwyJWZlXF24/YCcWMbr5MQjPJDfyrOpw0gNh
MKEYpdhdmy1OSmHK0+eKRg3KyjDdbStczihj8ZBnGlTjekNzGOlQZ06pZSTJNqWe
Uegyxo4rH7esl3F7WG0INsSkzg/Kun6O6dnRJDFd6o2qnK3QDvdWS1trZcpDi8pw
FtQY9jk0TQCQkJ32oTL9waejHbRUmHxM1jogZMXhtykdERDEymElrRvb8Ap2Qa4p
iK2WDYHwGav2NmhCLQ64weMrYnf6E6JT91sPo6/tVV3s4HhfTqz1vWQh4ZvebzGv
o9zSsbuV8nflikxw016Ra9TcixsqdRSkqT9Nmzox9IFvEWwKLVhw8peJRs1f1dEr
zFmE1pqr+w4lnqN3flSk/odoMjJOcYnKmw4SyUuoPpvj/fFl5JzjLnLfOLF8Bnud
zFxKtwiETVTH1smd+dtxKzzlK3RE6zsMPFMrNCekA89xQgNW5GRinn2YREgsVKRn
ixfeA+Uy/dzrymMn/FDV6LTwHRMGa1ZwOUdw65wxaOdNuYyRk3TC4/KGf22Ld4vb
89QQtOdgnN/xTYRCg3h2FFUcocPDyaWrTZ3DGIaLpU4Apg327nOrieYymm8mnRWg
Pzmr2PCYlpPvvfYVIJnM94XRRsFXn6IE4poD6blqNL2D1wQLdNjahr1aZ5HxGwVq
oxd5LH8mkmQBUBi/U/5NJI/gQ3Z1l/IRo0WpQellGAQOpAZpwwf2GUZJGKTvAUEK
Gmnn+e9JWa44OmnaVmF+aILLgojg2dIxAU5CjD4Tgj0j1N+u86RU/lpTOB8TtgjL
eYrd57tVndGBD0+yuUoGl3C19gl7dCHPV3/fNehXBVNGYQXGBdYHoSnOxDlWpkDa
5tHiVtfzrk9y23nuob8jAyjYH9RK9FuthKJOlQMeMbfGk5SMMJ+ADVxYQFR74TUn
wMwOAVlw1PKS5TK2eiNCvXAGR7LpfoGDT8CtdcGV/AcQ6Dl35J/F92iihmCx6Dnh
ltax9hwLlMDC8ffCqVREFaVvr38KfW41O37PvsL/bTd5tmuYhffvKds4pAKwaAO5
lrZ+8A3g7wB1r4nUckwJPTuKMn4cC75ucHZSqoJ0Ug4akPz9fbNzrXkd0TdNZNR2
woG4JQoYRg20g8pVHVPDi6rrN0fH+rUW/bQmMnIFZ1i6GkxT5TROCuaurosXYWd8
ekWkIfVgnku1nLCa+5HzyQYBopB7XzTX3Z2BkLweDhJaLmIjWg09JC0RlN4xe91Y
abCXGiNJAgJoijZRDs9dYsMqASt6kkAnr/eah5SZoxm4cnnnKrh57wbDpAAxGrz0
MGqJZcCGAYq3xtA9p74oGbdVEz3JyA7eN5HhMLPrnQggHB+PZhKDcJ9lqDv9U1XL
ONPcFNizriTLVF2RXyPXQq06Pf2vDIKZ385bv8BOaNK6Z29uPZ5/s5DXtWH/KiP0
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
YFvfn0h7mcY3XRTlhEdCo9u829gGwUnmPsSFQ3s8TTNcn7xOIsiSVr+6do8UfWSL
9jH6RvN/qt4j54MBOgPR5fO/UEGIRONtrJ5TTioON8n/BcYJ99vrFhJarfg7RlSl
4UZEbFm8R+mDkFPXvlor5/+m/UnYfMO6blmYRiRzP1E/E+aLDf47H7nRBp2SepuC
tJtFszrnQNPNisvktIkasKJhgm8uUlxY+zAUBDVj3ge1sQUiDdVd22kRo3TiKkiM
VmKzRZQA/XCAGgqIjk64s3hQhes7PEmnmw0vdemliNINE0Y5CkQQ4noHFG0G1/Ch
53oDUHj29CNGw8vaeLUxKw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4768 )
`pragma protect data_block
U0bzNn0rRJ9pcILrw5XGujmRzWxcAhGbR8/sEwoQxRQ4yOA/ODBpaLcNnPCLxHFi
TqNic5apf7CZCX5B97qQCj7NAdriIh2l7QOwDGRBs2yS2RmDUd2SZsR3HtFmdngE
NBgU/0svtx2s1Jfvsl2ItP57N16Jv/r8GjVssWo7+nmNuvI7nQeoLThsTXiqGi1J
JbXg+q81AlvPKgBb3tON2SQUdOa1AN2/k3qxlbFxRCDhp/3K3lodMH6NFiQfT3Vj
O8oxjGMaXsGRUjB4KqqXqORM8uvgurqvS2Snh1iI59zdxv+FAvQSh85kmudMrbxx
QwlOrTAN5+0f1BzP8elasGERxU0wPHk+2mlrNEd0GaWc7zZCTQ0aethSjkLU2wUh
+UDRzIsfDEO8oz5O4XEkGxXxqm18AGJmC5DpBcB9O3hvDm9UddTOv0hIYYGXObym
JcQ213hT11mX9I17mMJBCkBhTXxy7ZFgCl4JK0nKKwHE4UwiXrVvBElWdNcORf5X
aSU8KTGOkN/ODRkWw87OaRkWFmwYrFzV4/1Zz18gvmMOVN/Xl4xhwjSEv4zcVJvo
JaWY6KOrf7HooZhKxOUkPXW879tESWHbkMTnqEMEKRcXcGfrZMkk04eCUAm7idf7
fgbugbQAd+OOb0GDE5XBwQuJ4xEzsyBPD3UbRTmzcEquZTzk8teEZNTH98yqXh3Y
OF3nMU4CNtXH2F9hhEox9lWx3Wo/mpj0YA6/GIG+9qisyYPSma58kwWCopcxxl30
7IPGvbEKEqR9tDW5O1EialA/sA8aeltBZ2MqWw8XUlC5rKb0EE4lWr1yqIxzCglL
zBVdF7GyP6FNqpKSHYzsg2p3IAUtvTdypujh8npiSOQ7e/MOI80/t3/AZ5ncmQ6A
4CuA5afVMnNZl87F6UFZeCE8FD2iwwNP9/iZ+3KcXB8StjrQJqIOYGvwSg9n4Ym0
6fPoqmmpCNZCz9cOF4tyLVVryZZ49VcU5AXXe6ppXaDwm+HnQukB94cprWaxAwGh
TF+G5amRTR5RW8McK/yeRSpQ4Uv2h7V9GzCTniFTKg3BMzKFroEMR6N6VJ6hMYdL
MI3+/WCmG1bmjVdbz9eckSAktpWxCpQFeSAtOlj76x5rM5JDc6qhzoQ9IN5mwoG+
ubwmS1p4uhBCS/GZgoyms50iXMkPctPTlEGSjr06uBnydFuCaFzVU8kGqNpa4hxU
wx484hEkaAjQDZoybtzaHTqsFjdSubqhAh17jnZOk1V4rXQ0ewlVKE0ojUT+Ko5P
mz7iIQwsjJ8i5lZ+KyXTZ3VycJAktbxR0fZ+8tzWtOKy7Xb06ntnyQnK59vDWNu4
GllsutslAobyUPLbpDxDfNkQi8t7jZ2/NR+3/TiNpkpij7ENufr3zXEE2UIdU8l7
tAwiHJ206Ho3Y0nWyPlx1cbY5U06ZteJRGbVRA2C7s8Mcvp9OiG5i9QMBKeeQmWB
bRkFVtGet/j9gLu5fDM/O8JkxKHE2j2XyjhJonrdnTbWJFbk7sUXb+0im1GXXBT/
eQ0H5M7sI4ih9VMkEGdeNJDzK3iIG02eDEHZAY7tosHbLlHctQyhFF/EawGql0aU
UQQ+HNEdyNYUDa4ta+Ud1Q9NxX7wzezWIhOahrcprwSa2k4Aq+heAKTNoen1hj8b
TqYcVFNQeUKGzcNIgkVM6XpBXD8nt1bl9WnoJnyxfwtr4y5UoNOzLk+AX74WeMKe
Wrk4aU7QU58mF0wsw6dWfOnhc5361ebEN0t3m1C1x1FZJ1wMOMpwBBxxutLuCEJR
IMYJZ1BV+ScuTsP6O06QPhcVwHpmux1oqwFlpLviZVEie6aO4DDqzNYq1al6RnIZ
v6AlDV7NdYy5fZ3U1f2TngYeJC6lLKt0wd0SC/0/qfkc1+mUwDQzUMmuL4dqNKRP
kA+lgvVWkSlvCiG48Ps30AVI5AgRTOftPui30iFHCmMdXFC80xq9W0t2oAZLMM/1
XGBNkQetJSt9qvs/BQj0OBM9C6mbThSp01ASloo2ZFX8YGtcSYdcVNa+pY0CRyvz
WpZfhVYBovHha+c0ULxapW4oumNmvEnEdf1kjTn2/nnVeFqLHNvUQnQvwfpbo0Yg
D4Pp/PQOrbAB31JA5NNuChTm4BQNDdXng1/mmf8lqhsg3k7HckU/NYVmwte/x4pR
z9lH5/p4790JdA9dT6EVOWJT3HhqCrFyM3E9eOV/G0Uk0EUk4QMcEO1HiVAhtjIB
UwNJflQ6lzoqwpwlaVAh+QBv641UINH9TLo6uDq5JSCVkkNEly7mdy0OsCf06hSI
xmIsZbYHXYUObQC53LwKprCIz6WgXoo6CUn8uGqAsT9GqS42hbqMzyy3H/XK8w34
O8Pn56IbBVCeWm/hwfCA4umcJqMl7hn5M2tXCTj+sXylyAUiA+XbRCKGT2fo5lLw
7H7oU81P4hi/pd43J8pzUc9H65374uRdSWNuS5GJD7sYrhZD32e4/V/5ExvAwPDR
tvJGpEwaQF8lVlImm6oUT6IrEF18G4S0pM3fb/Xj4dg/oFf9jsRpx/QvsBooihmX
9+HPvODKaDOes5B9EcyLGubrhjIdrc1cYo5rMQhWovs0tqNes48R7ps7oNdb0JcJ
ycY6ERpnBvOBFgHlsVf5pyRWbolP6EE1ajBA6Jw+p0VR37bL0H5PPDxgp1HnMPVp
/YrOnYVowmuTu0RWOJDKZSVRenZ9ORkVIGzWGTKB1TeStsJW/MKAwloPfP+EZfGc
dPBi3RnwrSActzfLZOUkuIWUEwHdTIXQRpJDMH93s165UCtMV3Cmqb2cxz4g1yr5
gDm8hDtrESnaIlKnjcC1hBsdu1TcM0Q3pSQWQZh0ZFyRKPhP2wHq55DshEb6kS1n
ENdG26ZhUoEH+f4eoB/dOM0p46EU6vwvPo20ws6Cn9DCO/GTyuRwvoN2O+ODYRhf
6Na5rzJSfdjVVq4gdgI9lR7XcdUrB1ayXBIKAnEw/uaY0TU8z9Appuz0RIzsGKvE
+16IxaghTw9IEyxnU/R1Y7j9jNZ/8qqVZpgTYe6RO0tADbSYjTFdpQfhnuod2eMI
KLi7VLIKYGunO6zrUDiBydYXv3s7mpWHQhPSY4+jDxGDh+KobM2lsF8uOz6zPTWH
PlRRxkpTuOZz3p45t2ZfdQN9sN/6StEVmbj7rt9nHN1n14cwrIrOPV7meKrCyjuF
JeYWG/FIl4I41dY3GakZ929dfFfozviFZ2gsDr7uVRBWAXEBTxDmgosbCtsIG7wF
UrF/ceOsGDT6k1mycHM5mKLzaSvC18tQ25w/i4B3sNgTm0QsBVIenABstc6fctjW
m5/1Grw6xS25ZR/vkOcqkmkOLOwhiq3x9CvrC2TeJgjsuQWgcTieWStVKDXnTRnD
L6r6VXZBZS2FCEULLjDABOm6X5SVg5aAIQETtqh3tLV3+BFuCbp27UhVZ7IEJiS2
/zEGN2bwJVAMTygDwls+gEDeBCjSC72uhwWoJSeTzodMQbJ9VItolP2NLgTL1avI
UJD+CQXJY3K76ykz7n3KpdXphvVEP1EDDz2E0bIGWzEyvCAkUE3cFpOAXqoNPR9x
x+2/kOpouy1etnL33ZkFM89kzzNsPyuQKfLshVVxl8Hw0CQ0gBL/PVIfEOYPiwgR
xpliJiTxKPbGiGTt8WWDulTGoQxsZwPyLogB3OHvHcUOBIo9448/eUORePLjt2ZX
wiDwtOlNG/I9ECvYQVRqPSOv5L4hJk6XII2jCp5brd6NriyDSRuYt7HseizZQSSn
tZpv/dWF0QgCivfbqq4jCcAI/DzSB4LfdQJeatAG4xMYB23aT2o+qSAd68DSBtEM
yE4XyIYyjBsvEr+olt2FQi/70Q/CRg71Mm9IXoUPQml0K4GQE7tJsDEjdNws6vQa
lP+YuEww5U2/dmBH52sg7XhQ0TS2lzAint8/BuFQ4gdwk2HQTQFj+yEPfW6r+5Gr
QM9+Pc+xbQsaMlEvMy51jUh5AXcQ1CwuulH6/55YQI3KeBTqpt7z9MayTTDYbPn+
0IrFkVNW4F1vEVhiHRRxCUCQ9bPFutNV91nC86Mr1p5aOX5PU6Nujg4ROTX2TGzC
T8b/3SlNZSywttnBPtBtgAONkeH5Ho6LkZ8hJzI/QOpgGbZIiYyekM6xeX8I1Wn5
WYEYrUOAPqiU/6+CzHlSegqbDURLBPv82NwSYFqGrg/K4KjE7WK705w0wSDT2ULC
rkcauqp57H21qhbWjuvlXn1eGZKVHA1IJZf+AszyiPNr1ghMI2WYPS7az/RHDtaK
AnrFMukkD6TEW3MdHOdsOrTFpf1sjGCSLVAmDE4W8dhSjnKwZZTL201i5gexcNu3
6MS2y+U6gnTFyPBFXnHteNNeoGzpO/AX/DOQOUQXPopnahIyyv2Do6kWGRAu/bar
dcGvj3C9cPQFKVJQSW9XXB7KEF6gbT7x++srqmCui8eWUn07DrRLfRkmiMlFJ93H
wmpQKxLQBP4oRAsChZchvNkxVO3hOpi9CtEk2IIkInpsr3wvenoRFU9CwTzZALDW
Y3ii8TifM3YKIRU5Q0rc1Fgg+l4ToFmrevon6+9Tth9YYH9gn6l8i7tXbzzP7K/n
oBnl7b5GionU6hYa3GuX+Fc1JfFBLTX6KZmnuDfigHg+pBdAAYea05c5HeMAls00
MJSkimILZz/EwcaQ6KSR9i0G0O4JLtslTKd/leJbFTMrzuLdyDvF9ZXlSN4w6XL7
3DeJb4uzELXD1FRkwwSIRvNkojuB5P0vb0uXYWFoWqXyZdSdstQs1x6iP5IV7N6j
eZusn3TAppZvOpJ2NDl2gO28tmTuO65dvc17fPjVcLeczVRKLkCaVCNcZZ7Dk7Ve
oJjXiZeMcz2jdd4tbf/ZKIl33ObF8pZY80z1usRTkH6Jz3dG7ooanQAM6Gwl7z4v
8waIHbUUp8wffY4BLEmkWPOvyNEAN2pJwWaUTK+peWEo1meifuJuOs1rrz3smh3V
m2KRaekUYKcC5RWNtvYxLeihay49z2Epk+DT5TMFc6+y/HEJkhSyNgiCV1pPigtm
lTNCfe+6NF4h1tYn4N8hyaoAA/1UDUMQaHt5Ab1aNxdo3ALQKKg5ttsI4GSwuun6
t3MlmHVp+3qYxxa26MJsRubk+gz9HZyXE2yJDj/B5pGACW6gmWCSyw+shUyH3Od3
T6qIiz+Z1E1JdE4adDPNQad7lf3DpapGXDl5aA1S3oqSHcZLkPFEaJHBtN0D8iBY
u7xnkMaq0m8xdmdwNV1nReNWEeGSxypQEjUr7JEGfU8sqG8fBD6LQ9WtGYmqibqt
EFteJj1QU+Ck50Gskq9nKVXstRpUU1GvQ1wuWcfB2RQBaCs43yFUMeWrRA93313s
u78G6S5DLRQ88LVbXVoGXfcAS5ICgKmY4yWuW3zzqzClbBTj1DaGoEh9gpCx3XZe
7pn7QN8cXH8jMRaydjY0sYrYAJ8jWt2I80SN+yzAtLP+91N4AtAHO+YMNOAufzlk
P1fnbt7RAvGRIXPShR2tGpPMHbc/xGR7sBPemSnMcbFOOIh0yowLgNUVHp14Ylim
mNhZT4HLFY3De3FJ0T1PL/3QdolXvl4KETK064cC6JwlGm7VSjGZyn2wPFYRVsED
YQqQITTjkItNWRR6d4pf4H3D5T+4oRd0ONXys2CBTJ06Eq6hnpifjr4xpo+bQDB/
Qb/3XI9Rs4F5l3bsy1FeTqF5Dy/URN9LIeoYF2l/MCFtgy/g3t+6HKHdrbq7CcnH
tICo0b6aOkiUUJBXcTb5mX1DjY2zB9YcWafpC5C/2rvM+wwrIwGqI9j0rHNlzrij
NrjYHG0/c1ZdH7sJUpcrIulR+KeotbvLWAf8lbxBGwSj06QyEz8CKV03PAKKgNUy
DVv0GUnYZWxz5vaEHONhgeFff9FUhAYLYDRr5up8nX7mhU9iiJQziqfCIAfnUO3W
9TrIqNFobmey/apT+t3qn/IwXtrqD/yx/hM4ig3cWnX+kaLLE6geHCaz52e7H0Z3
LEEshUrswJo1MToPDguU4zvUdGra7tAkcVkgmJ0uaopS8BtsC3jVMP+l0uumM2lJ
46t2+Goif8TGduiG/lDR2vQz/U5t7M5mELEYSJYd39f1qEl/LE6QEAjbn7VCkAUA
QLzYGun17csUfBf22Iur7+RvitmMIwFceyzJy2WskPIglJy3u74xvz1bnCntFTvg
zB5Re9WrfFCtF5SBMVcSb3nLoCuwiS25u0cR+OmApiFm3QWIGZBCfFUuvrqj7llF
yznbbtQ2ujXogvArDU/bA3Rxn/inAeIcATq/nPXAZnniSJ26viQOdczPewToJfza
M6WpQw7vtxka4OQ1iCIbtg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ETA5vUdCwsChX9QWvMAu0Ty5BFD4Wwr76slUMwRiPRR01Zt3/RWYVNqaA0oumrq7
AlMzfSiQTGGlR5tbjYSgfGIXpbL2NxYjngSvaSx/M8DrhiUdBsNIW13Zan1iassv
q453MojxoR3vpMKyi1UKuiAIovgEslMtLeNBDpDQTbfZIYXo9raP71YG4frQrQUb
oAmhQugLDCSFaEVvjtQjOfrvUHMXGXVGuJZD5cZLknwjBZHDsn+5Fi8JuJey83VU
oei61RyqRcFv4aWuoj/oSgXvidCKZgTnm2Pfx9w2FKRJvbAr3YIHr40tdbRqMdCe
0x8/VxytWgrRe70M906L4A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8720 )
`pragma protect data_block
kEBd/qM/T9qt3eh68vldOWigKOwrBRVxZh9x0d5+hOi0C1dctCDF8gF30YlWjeMu
HJrRxmaIjqTTXkF9tOys0K9WGLgQeVhADVJ95Xr1EW7VGLJlXvRiH2uKqIioceuk
1gMfVIvDkTJcsSY4yvJx+WV7Db7kFF60OTg6JMESlGUAgKhOkwwXj+As+xJAUIWd
CAQtnNVxvG/42YYAEjmvb9EDAfcZezNXVncUZ9yL4kcUn300Y8Q9dJIj09M457HC
SsV8oaIQa5c+qcFzpTeEndh39y5vtdOnm626FRB9WgUImNL0MLVwB6eHgeSaR6u2
0qGHMTwdKnauiloRfyPNQ0+wAEm6tpgKxA4YJu2hHIJfuu6l/Q1tlDFfm50RmUxs
r+VcuXv1UgjUtZk2T7s243+V1ItVmcgLb+PseqzZHU9swqrgFBv5L3IHSLK+E7Dm
Z8lXGHBLq5QdWA8lWLAw9MYFWz8HEKeW4sRPZlnasVnMTInbrF5uYKgJSybpq8en
rEMPK/gnTC9tUjaytAZdqn8bE1Y30cSqU4PrqPJtJmRkt76ZbNnyNqnnh5zUbnvb
2y7u0Dh2cid7TiHrdJsNRaQv2HLAt+xZqdaTOZml9DM+PPuKKr4p02I7jhrYymXv
X/UKHsI8Cn+fBIFhCTC+nCGvwHVIVv4MRqVSj6ru8F9qA2I1HmSsBb+n1SnGzX3a
pomt6z0AGKQqbFdU+CcSoSNw1fZp69hplsaDCKgD+1cOy+Wc//s4bDRMMgXIYESq
B1xKNnmAWgbrHK65ZoOpfcwEnSjowzgYW9KUIKPZR4dMU//K8FITExJO725IdF/x
WGKvXflERJ8rFkgB8QYJw7Wkliv+eDBeft9/8DxeUHPYHpTcGwWnolkdoH0IT8KU
JBLLOJnCHi//Q/FDw8rNMfHBqeuYElBJEjaArjw2Ti2gf8jM8j5yMMBqYwytXy19
CAwr5c7q4UnzCD8p1LMAVrx8pALTd3w9vkbUsCIFBdv38xdhg+TiFyVs4PriVw+f
B5/M4xSZqc+Jutl+VHc2ZmtF5ebdNmaDKGY90KFmllwfkqgpcjs6EoAuO/y1Ef6P
rf5Iqu12S3BssfFes7mVoAqysw1CA9iWpp26QpHPQ8vidgOfDCMe1XBBWxLWtjrD
b8shDFGR4BIV0fBo1I1lznnHXmxna3xpKYLAAx+8VobKo8n24vyVMqedBFzmduOQ
nwFuo6U1Hb6MPWEFReFvVrkDdsc1gHSyt6/0IM9H4jAqkKyb+ECwhYedIm3qEF2Y
jPt/rjsDzGN4uG1+hyiHvq0BgBUJAd8Kcdr8TVvGGU+NxDQYauKTfB3K6TRgAyOs
Q+hRE9MTqNmJfUAjOEb9PBOa60H/XjC2ONZPznWAguclJOOIrI9J+U322yu5933R
O8DV1riNx5P9VGSLfkrYFcPOxd3rOb+DJKfTiT6VCa/uWpia/Ip3u75LsT4ddyUi
SzKiPQRaew1bFPwyHUw5s6NJLDEuZWXzq3WpdqMNbA2JEAA2g0+B1wDNgmiRAZyg
YlhrUCvs2fVZeTel7hgpcH+VPNnRkvSwRvJkJ1MOIfPwYhkeo/kPsqPun0sfmSP6
MkShmSMeCvUnPa1yIPoo52PVlltQ92C5F7FOcsmqZaQGGDj90WKixE1DPQ/i9RiI
hcTTaAsgfRXQ0trKaLZcLMZwL1s2lQ1PRbovcxDh9FAS66NEfaNQuSbWL5aGMV36
uiGES5+g42xep15OjYtc+u5YhKv1970VVB0VzbK/HDsoub2D5MGDMRxWSRkPJXsy
H3NFu8NVHqB8EH061FiSFvvr/jcCag5JHXWZpbuXZv+g8LS5FG1VFjCskUfaHJCR
7LFTT1HD6Wu7flvHULiD9G1zOYViwpkMx0oWc5+a2/Omxpy3ZxESR3eg+2UOz5hV
CPWalZzvQdc3yarw6U+tOISgJB/fmWc75ZKBw2yJWg5k8x1vc+RXt+Al/ldFIUIa
HOHxlvQoIpNPzkieT082p3ukb2JrSGBRIkVlt3JbCVI10JD0TDy4GzsPylP88ibH
lJ8eK1PzBl/84Ur/AShuvZqmUz8BOjIL8PLIIyvcVOD8VUqaxUUcqngFbJojPf+I
vHDLS9z38V8oF03FhxtwlEmrNfRiWOp2HRrhyT4OEhFrpCb9VEIzbVVKAYKRxFdz
3CqEYv8oTTFRIXP6Ag1jVtg0TB7xWRbwdCfFZJIJ1DqSlyd76LB8NJmDK0AFtfV6
4kJM2xpoXzjUH2c5tZjCEnk33lNPF9Q30y9GLOfWzWHV6s3ZJLASx3VXH+nnbw7B
rcDnD8Fo+vw955p2sepFSfJs6ND2AfcanIBZCepXhw0+H7We7dmn9iMLGrJP8JMb
sZqSioSyRIoF/bqGRmPsnlnkh35CmWseOjld2faSJZuWXEZGqx2o9Y2e4Jy2vH34
kKtPA8PYm3rMGKD/8faXBnoR+mAkNh38zgukDEg6ah8smVvo7yuphTlkrLxtrpV8
ccHkj4GFiEzi+x0DZ1ks2VhZpmow34g4MwxfFGeNWnraInNbWbHNQCV6QAfbSAvf
Ho4DTP3pYK3seL7zJucLpImpXkgo/r7BtEXbWsOxyDE5gDZTkKfMryu8ExAVtKF1
cxrfN84eUS3Pxu3j6wkreVEZIKspIEbXzyNA4YgYjqecYtTK0sF263HljFYFTpJl
PaXSTl4fi1oAq6S8tyFnzS7v6fkURYSV9LK8xGLV97GMY15u482yLM39g9C/9B7R
esL4wo9obf7EegIEmB6oygQe5EmrhnIqG8/ZfuZ8/xq1c4wQEiMdouTrc7883wZK
NUCvXUd8Wqe6UofsfdpFXHscCtNGi/w8YNd26sJqYzR3iE2gtarSFRsJZ86ZedP7
8t5yBJitGinTioFV+aPBVtgLR885zY9cp1SK9w3GpUlYAvB2LGrmgtFZ9jnpPnwq
4AHnKfZIdloo9jvl8NiGS5rxR6UYZrYXiBwSZDz+/0V1pafE+KyrRpcJxdqxhMNZ
SntRFNOe8sWd8BaUNFjcsn60e1MpO3KqQ9WQCN3QP04hvuiipyKux7yDOt2HBz4Q
DvkHuuysaqWtAsiV0REneeQtsWs+MhWScEVp8O6iwq1KaBs/ij8+VKIcqzwZPZSm
TiHyNWtUpOq344KDgv8gAyo7wiEu/J0g/P/GNPcIf98HbYc6MlDLb894t+tqnpdn
Zc51sKXGSlPGN2tDfD9VARIfBZnCYJWi4yMOyhT4iBF9AUtHXjDdhxNKzVbDRCmE
HfLPekC522zJl0cOaO/JB2rnr3uvOJrcj1UohhnGbak6h3mfiqz0CpI2d6Eh3ES4
lOtxwSU8RhnO+QvFvFafml0ytoyhX+TWGQHMAxK8r04kGvhtCwCOj+ou2VTPaphv
0njMbYsn4672kFSYvUBLtTdfl/Faelv9lesvBQLiUkUGncbTX0CQhy+D/VMFtlf5
jhCTpsR8nE/YBdUJPf4OV1MDuVYnoQ0c/9Ihc9Y/44Xi+ImLBOnhdbCqhsqrVoO0
7vBnbA+uzUU1EzY/Qqx0C+nehh2taiDPTv6UKZGaLnTG6FupgHDjpx2kNh7ocxLq
99Jf9OrwiwmFDd2ufXEdtmRBLjZw6ZHdJLznMFLhx8FAcbh98Ufk8VbBapLdCx58
3XgixIDTYnrd/hVnX/yG7d8651f1WNu6KF+/GhFKMFF4e4e6byemNHg/m2mLNjgO
CZLt/izvNNaY6ZuJZ/Q1vULg+hengvUmtnubMrxfP7XtiyJ9TpdR/edt16PZG7I5
4NX+QkI21DaWsQZ1U4aSw2/8z+O9PpDaTbIWPmJPbue6AthW6uAQB1D4ehj/G2cK
ttV3pt0oulz+BLJ5tlRZnhJPpKmXW8NTfdvqHgkAv5cuK9LC/YmRUCtQ/ZD01Sjj
pu+pgmstz5BoyaNrq3urOEO7UBgxPxh9OZ1BxZi8YYp8/UY/SmFCiGIQHQADRfLe
s5a2WWt6aopLdMrh0ssjGKKjuonj3rgy/LkgUgBRpW8543wVfGCAXpf4p+hFj98z
JmqaU3dOpj88MXDba0FcQjZsBf9+8VCXOpLOuFpAVd4fVMLrOiKjJ2L6G61b36n5
GzmHAf6LQGGToJQUfYHG8EX80XcQZJlAWFBtMDz3NyK9i3ULROZE4lxYGZET2Gua
WYPudAHwneZucybn2S3F0J9scXbYzrhM5UdEggkMTaX5mIxEz1LRxhTHjpfXMgVq
Wcu9CUUoXoWfyAFSqS/11zRHX7zfYpkesROtgSLnizUgq8mcC1cPD0idkASDLPyy
NLguPRje0v9ASG99aBZ3HrzszgApKwd4WO0AyeUGzQAsPE8C7+JCPn7vwHbuWBMX
8u2tym7CbajyLWz7oQxwGbf3CCV0G7u0rjFkwe+FsAb19bCNfbbaxZpMKCNWHHRP
UKblxi4+tKUdVOPNg31BQ8dAD9OCEZutU2JrK0EmXI9h+PmwPgXhZtKaMNzveKoB
VCxuiovgqenYHiyIPAqBJDmVzATTnroTGbbPuI813KOZrsYYl7Rk4E9GZCiL9tBj
AmOCJHdesGeGV4gyJTwAEsI2Ma8quW8sLiYRFGltY8glP3TJg4+BRgiDJ0YW8o9g
wNW8Ti7xXC98orORHSalnOPiNIiBmMsu29aDeeDc4rlItLjkS8OBTWeROvb1efLZ
xUqWD6LiX7+lxlwOeRNbuQI27Mf51iJZ2sW/pVPWIg1RzuHB/N3hdtPmW5Ki22RT
uKSx3qngxG7WpQU67Dk7hCEuxvAsV24hxpZUMlpLYY8saMlW3vcTEzPbFv4SwExf
ICyO0+kHazh2EAWBvCzoObcCyPbTvhGsgriq+JvNdgLk0dxbrguglxJDAmUrDR8C
F0DfV6NS888O1OO6+GM+LxHQjF5ik0Bn2XEM/YK3/qinuRzP96/nQpku9yAUmd4q
gix/9hD2qFU3ptio5wF/MCvxbhI0+G5z4xw4+8oHJbLa8rohGCSrK1OhJ1UutM5V
ztMqK/hDYEGRXZLiu4nnzETkJqWIKC8whFmVVYo/stn9XpyhMAzml2cVrhxP2Pv3
onw5/b3DS6W7IFgR13JJkk306CAdXx92oHrPAbuGtiTmP0LVDkjfyo7mXDjlv463
HnvH7q31rUlbQD9VktAq5W54azzyiG9eK+GDtEUJAIlZ+in2GgT+0XaAeg0xyo3q
UAI1fNwwr87PIx9uZ/qJ8x8qnqtZPWGH0wmEx+gAJe7GrpTXm/j1wBWD4UUxUkEb
iOIgDGGwoWy1ZfT7/W8lZAHs1FYh52LDUBcYIUifaoGqHnI/5+XZppUBt/SY9yYf
kR3uJcEIKIhVFoWBqzwRLdX/x1a4SAdTbK5Lc2+qumPqBb0QcJYQwFgLijlTi2w3
PZT3RP/6883dRtEcCRb6J+Tl5pkt/kw8RjA6YB4TmCja2zdNP+CoVPiS2PzlY2aq
E0nAL+TV11Xf5ABeKFlQ0i0sUnmeWoCvtKSrv910lYBes7lvNNui8gUtvGHDwuAE
kwWfQVRoE5DbZV7KbjJpGPEmwmHhXQMUR/YLNV830y0AWWNRkKUCV69CNJsrxxFd
CzfW7UcrlUYpzDqNF32f4VR8/S9Oqw8Xxdf1ZR90VoCaSplDw1TbWaUcb4rdeoC1
kXsGEMjUvuqTAbYReZt6oVL07x+lRRCyC9o/vjQpaLJsc7xf3S7GA3H1a+m1lNco
4yOk44hNZ3jpje+4bQupktckSFlwGjcAB60zETTUvgwnKEdUhZ8oHmko8no5mvzI
cV3MVIdn21nxsog9jUoIU3Q4wHr8dyFSOsJd4jxYbRqvKX0NvRlX7z6FzpBYRN90
0VbgR9fOxlztpVIIgPZHnN3y2HQegrtf+ebeRz0giKvPa+SS67abPYJcFHwIXKyE
eZgqoD6jTCVDz/hT/KwCQGX+6Erez50bbJbCwketlyRVjuHCcT1gf1IX8seulS/3
mAb2cwiahLKXEsrbeIKkjLuZCeOITcSXlMXBNeBYD08bDl4pkAp1B77UxHyxtuJj
SH17UGUhMRztFVpzpy6I2GXuO1EXOqAzHt0uBKnRKdtsvmbJqXSn6XsrasGI5FBN
8AZ5MItJGuitbYvlBjohAK0jHSUojXFqL5ohcUNsEheiIA8XdZghW+oK+jQq4QI2
vb+ieNsHxzpoB5MgnAjnDCsvADgQ4X/Cel7/WDGW3d12fUrSDErYqWget6NBBDmm
S8DkLD6qRmBDXZjYBL7GyyNhiCq0hxzIuLF8rFiLI7DkGb6KbjgCALebEuViWRT6
H05timx2bndDWaUup0cgZIYAVabKAseu7ADSBu+69JVwKzgDkeTAifIJHbqFiFVK
ylQqjO4OZlUmU+34h0Jt3MeAeyJu3dmalEjuCPU+ae6iqRWFR42B2w/S+ZeSxU3r
N5jfISVmKj4j61bsxc+VFw5VavVrI45gXwcZ/2MuMWW7yRqAsG3Cnpu8R3k9oXSX
tdOJ97AlkcuTrehVCQpRrXqGd5QTLxFobg0oCu6++eD+oxDoG3lfH+dixPVJTcqx
Ao1XMIt1PFH1ykml4QxA4yMwfETW2kAwnw1iPPJvdFSDElb7Eu9tbOABWsc7Sqcn
jwXQBqbG9jGiA3l7cOT/JPb8oHbqSaRacDTfYkbhC4SMMDxBNuhdoUd39yYLgvkD
DHTYh0bTAONlVXTFer10a0BgLuDaP9loSUMQWApLWbLv1syWGlmIuurAtjfmq4oF
NEtj1q94GPkDbLcb3/ziJAypjksMarnqFBzbthZjoV6vB79xxGneRHe+/y9feQkv
Gm5U8XkLVDBBHFMFWdHzycMLpVv/99WSzMDpHUdgaXHOj+aci0q5QQJFv3ZGTDn4
m07ENMaRVXR1S7/mgLENLieSUHsqVMamEFKcAO7fTtifaDygBYXNR7KOEByKasxj
sA7R1dxKndXtkN//8B0HCF74ETl1luRR7jF9KfTW+SMPa1az7n8dSIjqB3lU6n9R
I53qJZnwExKu5xH6oZmy8qqyBB8hnK7Nce4r5V64H/g9mmESTY69HBJC57hfOPXK
8IObbyFwAkSydu3el04JwnHbYAYIwtXNQeMC1WAWEeaQiNDPCh20fevKiFHnGpGP
KaxJdkpXJ/Nd9vCzOlqmbt0Qo7gGisrCkyNfALstljEcSpOx8uQ477scfZu7OHKJ
/J9AT7aJqftcUUR6BvisyxhK0TiqEiphlwhD7qp/vdGGcC8aqAdiGm7xyPbtvbCF
nj2HHWxpi2GkOonRwM7p18C97hDv01SM90yM/9+wtVbsncSZkqySc/HKXtxAvjYU
nbMYRRnCNoEBdXH0P6I0t98EzKu0aTsi0JSH/AYiTMbXNJZQ9MB7F5ip0re4R47Y
QaqjW9wCrXo6CTnwNIdt1BbJ53wr2Q7iuqSIh3t43qa1nesC5xNhsEb6RfDHbvo/
6OHHoNsIpu4ktNgnM6EpaFhP+ZweKgnNzEdjIBeU5Ym7Uki56SP8krj7KN+Vw6qV
3t4yp8hvzriN1hToMQcG5c8DO4qrfh+4lkuSf15BvBysaBv+HRoyzqwDiPPNWGh0
ngqMt08+bbNjU+08TdKYIqs9KD+dbV7re8Y9MGSnfm5E/Un6Dt/SZx4eaaE0KKl4
dSmYNAsui5i6rWCNYTIU048/xKyVKNKFOckh1Sej6/DWOZPBNdkiBRoJrVF4GKyt
zdr1XL9K7d9hZQET7DEcPzY8RP+CJ4me2AhdfAsA65x3YdT/c/Y0Dk9E76e9kbZR
kyh6Qod4UbTfFNuz98upwi9FbaN7SGL825k6VTK4kM7/7kWev3GssLUwCF+Pq6U8
s1S/PUr9CuD7K2cimtTRtsfju666SJSD7M5st2Jct9jgMYGxUU4g64iE1DozJSVw
4fdu2eu9XHDwpG+oIIm2n+qMCZv4/CqE8UBVrh2nuJd/ZfsFvmJ0Uz81w3RQpNzF
xT/LWUcvNruF08OX1HptZDnBO67G2wIVAAj9K1CJYUHEfi8B/7qSCbki7eTy7Kqc
7dI9ywDn0ijSvTJzVhEzHORNJSYgIpvGc6AinidpYVU1jy2BqBttHcNu896x7RNA
kLKzXuTnmdYh6/IStNQZbrL6A3CIvfZHL5nQ4nk+RX3px/nyTvOtNiwR//naVIQ4
XlE+p4lMhwitavS7vafovsj1AGkMK0GNN2ZHUyoBIeSGF943vjFLJoHKTuRKoh5T
SosEghx3tdauxA2q6ZYMym9KCyGu2Ooy3pejy5MkeiUaD0tIqQQmL5h/6wzIbaJG
97pZla5Gfj00/lNDtA0aq7i+Vz89Pe6PaOvvuRE8zBZPQ76Z/Ej2xvmkJBTvjmdh
SUF/jOIgamiWPDIYAJjMUqdTDfVKlqe1xXqBOD0gUd92uJqhZm4abvWM32tIhHlY
Gni8do3ZmxfV+Byzjpc8wSvkVMWicebzERVDLJuIuKaSZftMoU53keR/A1ALzsck
ymSUE5FrQ9GkT9+UvrKcsI323A21EKyk5sbWG29FBGrKNCXFL9LCf/4D2Im2u8uI
OnK1iSQDpXa6cRPNZ2EEBjRWti8k7z1G/3NUnCnCj5U1A4zvnlspfGDL3dSeSARr
mqQWBTqK+ENDgU9NaiIc06XeRiFZBNk3xTDCQ91wJd1dX6cwxluM23FbI0JN1uIq
clglH0Wk5LSetP5OsDHws+aEKGnTklhAlq2jXL7MA9AbpUCywUa6Uc5sdkxh9ZQx
MW1AHKeDEx2TNiqidcsgCHlIeaKhhMgsuA8J96o98XVvvThcu0knzHV+eIaLxTTU
/L3corwvczvgX78dTYKol9iKCQxQSuCO0UcXOGdihSYoC+g7Utimfpe91XzRHW6P
Tn8et+PRv+Vt2gbhON8Ddq6yV4VEyU4moUtST2GRRErEXhlJ8eR+JlW8BwZAllR9
9FKe/h0HkvEHGJVAs6a5IHq3h6PIcIzKshhas+wxQz4zPhdMSv34us2virfRpLwf
ezZzR4totnkOzNDj7nXRQwx7HUz1rwPzmUz+3kezOMOUKpC42P9u+fyLQLDEJHre
3efuDnbkchOEvs2YWzH0TaW8ZlR3Qqnl4YCnf5pGe3Fsv1vwRPO1QZgWx6zg5FFq
oQoU9bjeIqYO6Xra4NuYM6ZCAf6341MRyk4QwvKLYdHyKdyFdseRzhfAguXDUoVh
giApa8zMGcYmUqyG3jfJ9wi3X23sPMcHM5gxFSrXF8xhAec0Dfc5uamIMJfd792M
NBV35eJ/Eby02XGTeWiA2OpZ6tfzDp/8056kS+vz1BRv2O1Is8TRh2y+zFVjKBeu
TpX0n+c6BNPAapF5xQ89Yb+gi0IDoWNQCDES8DQPHlMEhO8rVlqNgZhEnbQt3++B
3rLA64Xc58cQZH6L7IUNotL+VWl9zPwmqcEemAfC31G/TxLMlD+qeeN7xC6c9DP4
xSgdgmSS5TYq4XPq5EXqFXtBdRvhPd8+hYmNK5Ea3XFTO64cC8BgDMEDjJvzjazt
wbnPZixvdlr+nyv+mvdhKwaVd3kMYX72nH2rtMxtMQYSNKKQQ/vNOVcnwvb2WmEk
fIu3ew31np64AONXXP8H/y3AZiw9bVBYKLNtkftdGrG7N37xIoOOLR1gs+ka4tFv
U37RB3xsnuK2vGQSIX4DTvAuOT75kaAPx7UwgJEY02mPpprZd7jW7FYZgmcgjKHJ
uGmfVYCSKsZcyXWQxJMzRsn9uGqukDJlGwX1r8E4O6OvLBN2FiDSbePAngDfqVXN
DXBSWB99amzEzvqTWmN3gwLjueQLktJb3a1UK04xAL9tYLV8dts8blbJSS7OyttA
0QagqJkD7idW99Yfwo5tcQvyDVqMfdquFl8hI0oULrWPYg55X26pICVtik4/djg9
/Ub+QL42Q8xLatpwjOUeDNkGn4u2haxfBAvwRWbMVsXLxngsSP1w4k5aEC6WLs2d
HNTpcEHoREoEk8rcdqFPUAGe+ulqego6k0Gy56bKYT30CT1SuKjwnCq4JRtzNzgO
TkEk7PCQ5PR2tGUnWxhxNQI6mOT8bejteIiX/PI/w1McGkzqI1xm9BdmyKdJz+oz
DjlEPvHv+OJ+wgJiD/WQ4n53/D+uSJbur6tATgCzaq3tKT4M2THTvOCHZ69UWzDE
iL8TO8CWe04eDDFrCHjf4e9ZPeA5LomGQxo5V4FHzKnEi460PKXkjrOSYaLSwJDE
D1vRQ5zyPY3oroyzcBKEgKsEjcak4adnJU+9pduv9DhFj5dYQHg8KRBfuFUVCG8l
kDIiMLRoqmY8cTQVoxNNBvU9C4+3c9Zb2MIEC5KjV8MHl2/MENMkrLljW9JQJR1z
VmCQM2YsgfH1SEZt+MuBHK9Wu0UgafGOdboJiDTBlNSTB+SRKuTauYt9k8aaw9iL
D7Y4bB6XExTK/+WWsyHSCyjVFJVYhXnGe2D0OLMsrLJQm0mPQp2eJC32VOiwFoeq
RylJE6IE6QUoULT8FuzPOKstAOn9eeSIgDRc9HWbK2rT3+1OHmQoc/J+oh4LAFGH
u7U9mcPFDh0Lkx/o8mNaQ2r962N/uoqT2T3AXp/lNX+EntyvVcLDw/AT5c1eAkoG
3TfVSU2Af7p4mOlgQGWivIdg2NWMuXOMABTC9i2oZS9sAhocHBpFU4FpvSec1C8m
Cev8COYOk1iA+BCRjza4WUq/5umsdVev0A9Kj2QWG3w211ENSZlzgiICd/hbj9kH
odkhlE3mWcZfgekcJMK2jFHpEmSn3sjgnFGZ1sJJuywbsMFyet6KG4ed1qvlWYtX
48W8ar0IV02KFhRYpkLOuosNG0y77Ma5kipTtKtLyApWFcUvxbaJiXMpOwemOKNE
BWN16oWZ/LepoVWJdma4UwEEjeSyHPYPg7Qrhv1GOtzGPsVprds28Z82YWLqVtGF
xjEAtL9Odeqzh0hGZT5fDPh0zRZQ/NemzcBCZp8Q8X/iDKRVSx82BWSYuZODEdIF
5kP8NuqILUW9HnbVAeApv+nrUK53idgKdfa1+A8FF7iNzlua98d66wsBQvfue/dA
3Nw4cC8DXVRoH39Tw4m1XwHxr9V1cvSpfe2wGyFvl3QBRXiEkFGIqX9y3wrjaF2W
x8VmARKtZoSCvI9Wod+ye+3kwUlY2GhMAJh64hraEP2i775En2ENPZTXYziaja9U
kSbQwTd3aGSmHiwFJdWhpyChtLW8TQFK/VcPTug18HkmAAyYDjSm6YqQMjsPWm3y
dricGJ9njrVqq5vbnngivb5R+WY7lJEtBOP8tVVqAvX0p817f8WdudpBi3+fE75z
XthtV+rilVjZfGzpdCOeyO4peL8wycaj2v/lkU6UCXdSBm5w03LUiYoSRHxirZK+
JaSjGe7KrlZLM59lqiXAG6jz7F+lgAnNeZKZNkuSoKsFy4T/rAgTeeiqI82mDPL5
A/Fw3+YXypy816vi+FcjGwAEXkO1Fg5YOIp9AFzJ6fnPS9nngwG6GXvMoNzLykxf
Dsk0WXcjl7uVoK2sMN2an6xdYdoCf1c8yc66P59n9dbCCObD5/YsfSopKZGuBcq7
4j+06RyqOK6IuKTcPsD8QC+36CJY0e4rrvQ8mxG9HyuKq/uf4yNf1xO6j77Kv8zU
d4KZ13OIsannUsbO9qeUaMjw1L3LQ/eGDFDYtMHpIcg=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UD15lsZ7V++MLm2WwrmIYhdz1uZc1sBBMfTavi8NV2RFgxb1jmWIk+FNwhW8ON4N
1YMBEcze7YuXoNPMgD9eqYARhmWexBDd8WGU8LfuaBPks8MEfM0m38rcmv2GS2D6
BKCeI8rDv7+0T94VkYgavRii5yVxtXxiCSPxF54qvPomsGRd4tcXHtqQGe2y1GhS
hKnmNpAtnDu88LmhQG1GjnODT1CRF3EFGDac+zN1GB2rWNhTqrUC5kvJbj9iV4Zt
Y3NGSClVHemtui/xhLx2q+CD4snYkHuaqxxes0UP4aB23E5Yol7bupoJ5nq/Eqlg
m7JugdXKPlBKKrHo5nGwLA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4336 )
`pragma protect data_block
cC8A4d0+5+nmuKPRwUkR7dYmjMO62nRJScdAKWx7OpIJOs4d8DWQB/uVg8r/El93
Qm5G7L8H5owIcNPmuxEqO8b31oVdWeIL2XbTpleZIq8MRvwJGCHiCnvOXDpOdpMK
shQXtsS67snZVpXM8zsmwern5lw5bE2UyCJvJkKNVB+/29sCp5VjrFE7A3n0zSmR
mzaXYhKsfrhpFTW8gcttBG50MDHXg4OKollCEZasmt93NVGdJSN0cjJ18SnBoCn1
qecTmJy2ERfB6rE4qUNcWn7qjdsO56ig9da5ZMylEZ7Ge2wR9cOUjiMX8F+qU/Ms
BvDyDLdFRS2uHv8rl8kmgss3wn9wbAm9Ml7ok/AE+pw0SJxQapBcZN7HvAiVYTVL
tDIbxOlSN5+IBru8wtNBzQYrBEgZuOMLjaf0Hf7wNqSQ7TjmBu2s8majXcWRQpj0
pt3HIwzLMiAS3moU8rJ/QJaK6SlqBml6b+T4IKo9mvGfoxDmTMjxxZ13JOmKdOed
Xeia1pTZcdX/cVKFQGGz52TJVlrF+RPYMGDIuokrT1ezzc2Ke9rLo0qzFBJEEm7f
rlzx/nWPWBbCikLPRGy2yqqTU3x0n+SxfHmHFP92ifTgkyjq4gCNgKJGkrwXC1xU
cVvhgZ5rXk98em5cLi8a1/UJcc8buoFkS5szJ95cVP80Q+iZAv4Jnb6cKys6SPF9
XVl5+yN60TI5U2599B1w2vhc5ltzd0IBh9C4+baOicdxs5RZxEkLumKoM7aCa7vX
gM8yiltFT2OT3eh2PIzYgwcpkg1xV9sa5TIaVBUZ/wLasvz4yq95F++j9UemkbcF
cDdzkTn8WeRLm7xWNBiUQi9/CvNjvrKCNnWcS/+p391Zcc6OVRI8BwPF+qdg1LcY
6M48d5O+4JRuKmTjnihS+H3Wh31D92LWQL4Gfm/9o4uSAbBErHDLcja3P2oJB1G/
IiZ0LNxJUnuRT1ShjC6E0i1OvlJ7q86VM2wNXyw5ygDw1PZCEqwMBuj362uUvzD4
hxDizKcGJDQNLpS9Vef8cx4HrpnFU7UwYZPY5eVpwcqiGRTOtTtGhA/xMMx5GE+l
GjlNFXsJGn/DHSIq2yiJZcpmnhKv7kAbyA5O+IqKOdGhkmoTuMVk+a/Rp42RdPN7
16pgmwIOeORX3v70FP1pfr079beR+cXz+iq/p7+zaXLKCm07tyTxXVV2gudWLT45
70HETqy/WpzoB6jvKd9GKam4ecAkDUsaQ69NzHNBDLwf8KbMydG1RkvcIROn6TgK
eFR95ZO3g8gx9Nv+Y7s8p3KiC1zQeyIj0/N0f6iktmhUbg8WPCCGRJztK32pvdgV
fIfO9AfZOdfOvcmnP2xjKsGnQt7p+bnOx+sJcKFayP0ZyROzID8juJyEvtWJQyfG
xIVbNBRR7C88aOogvs0SuiiT9ZbMXm4dqHA9ym2Q+Q/9fg7BOJ4Z+IXWxZJngIDH
4k3Qy05bdGmr8TcqHaOzeCN1KiE0uAzazJGL9k8fc3ZP9Romein+Wr/8WkQ175L5
4bOfPpn7zaDoRYyTpUiB75P+E32PuAQjtdIXWFd0QCdIRcIZaPxDUrqsX/ptq9MZ
+yiAXYGKKRVG09rfTmbYddD94GFh7JrDJWPMKaITI320R3rSkVVamZqZ1AtJ4MOl
RMvv2WI/uMSb+O4X8zftScUvJqDOyMiVwbPX1sN6RcXsQgwo5Iie1l+pALxNpb1q
6T0wqNrTz7MbGWvCLpApPBHOJxAfmuVWoW/XISgYBIickvugiC9FsnafcO+rkDWG
Fep9yyjRRDNt9aF3GrVRgEIwXSbvZu/g4KeDqCEGk9V3eHVuAj7f5l5zP6LIETk/
Nsa7ApzzNJGViv2jLffAUJxUPp8lhpC2aO/7aXVF47pJWyJg1TUKuJ76fYwRIV+z
WJq1I4tSJ16NE6p0qf+SulmgOFLPbq1s0uXpJ4v3CS1lVOX3vGN6OqHNxgmGKhdY
2GbPbyX08EfLvGGbVfTIMcCOhJHfqkU/UgEG3kN5CW8USBWSEGx4KJcYhX5PGUJC
re2zqGavkiw82zWXd50mfLN7v6ZH+h1p0buT61GPUxwmmkeJ3ApQe9ueNDF8yOoU
QrzvprM4UAsjzwGYuCOYhorsAOuNJrkv1TZyYTZDAWGsy8Rphww1iGfCm5Fb7yjf
IWQrVoRljbSRjvafVFEkFygeQaGqDSLmICtl//o9jT+Old3dUmq5tzzT4i4Retdm
rUSah/nqEoCewP7rT14qk+YGR5WI7Q6s40248owEdUYenkZZfsJLYx8cCPZ9dq0R
bPckq1JlXV7uyI82Pt5OJzoftU9Q0rXaIDhG46dx+8d5BXBJcWR9uX1rH9wmKodL
Vg+wpVtojrQVL87W74Tqag3m3Jzs1qOhFbzx9D7uvGGvjZbPBqRSY3ZiutTOqkTz
9pZ+tD7fA3fpC5qBHCpPDGwdh63rocZPWpsEP5Q7nrg9uLO8fetXMrIsBiN0HeIl
qJC6l5EKnUxiSWOxHgnzwPXnKeVB9kpwbHGCuS6WB3jDqpjTp+Lh1lXA7HHxe4vN
CyfuoNBkgMVAvWLLFoOAkOojDq3Xq9FUh4UFa6h/HaxW2M4PM7rxY2oC7WUWlPcj
WnUXcOxvaMUurvt6I5hDwPBIIXO7m0E9XmxXfJW9BG+/hRCyOtfuJikCgvrsUZa5
AJdBDRORH4PhiwlXyPzdrn7YcwWnf3K8hwHw6pUoWqkBRlwfK0tAsA2lIdjAvKZT
JhEbxd5yfWl2OgQS8aLKTUawjH4pXBAiOvVp2Lfp1z0kEHbtmeNdusTo0sGrhtOD
o5r/FQnahKWwKGPzhunwzQxK9OUOtu0A+x4nfaAYlOx970uSjINca0kMvxOk3czw
d/kSkLY5TGQJj4KEnt00ec2cPJV+qKQdDyqYamU0KxYLBchVu7+bgJNsPX6SPomh
tdDHcUBRQGDQ9kZW3fVLXb5ZVpVn3j46HG0n5MJpuHLMx139Fw6Ny6p5kx/h6Cpy
xUu9nbNX1y3uosZWoSNkjT560/H/rtw88uUaOmj9HOtxIyuNQNhgGPCGfMdKUIa7
Y0PHgU7qzH2Y4lMrLFhDA5DpESpBB4nl5W79y7acktGldwLlHz2vOjVdDaQmUeFp
HVozAjOKDQ10ykuSpLIUHngK/Egv2/pYEGc574MSm7pOe6/ULM7EVslWaW2NyKLX
+yAcgGn7P0gGxS+pkpkhNBiFG5NZWTgTcy6lseaeM6FXXQydUCEdSKDezLBWxjgD
j93jLTD5Q8SbK4IOd1W/0t+sF1sjwZ6CMTGnICwKpChh4pZcLoBQbyxjBfTbwDjk
8JdVEeIvWDSlulK97dI5Q+Q7ruKKL4Zp1O7ajC03bZuaunkHOspbktnZOdVviU+r
DA/m14sj8XKN9IhoelAPwTO66uUa2OA5NCbEWLYmv3yX/ThJ3gvySPr41gPMOn4v
sKxfddkpLyiEcoSe1qo9/YGbp7GWQjQd46N3/nrMgJpC4Zr91ErApetq1nUvRVZq
1oInMBF6T8L1elI2DM1znM8UsCG6IxcikRVxI6k9hXVxpYJ1QrUdIidVspq8OhUG
U2C2NR018V9i6YS1VSAR5QFO7fSjbVcg1FhYxaCy3Ze2JmCw2/wyOuB6MczAkjXo
GYXs6Unhw4HHZ/W8sWLYiqcUdmQmuGNPOYM0xbZOPwPhx/OY8pE4UAhK7xAHhJo7
jpW/z+qGZtuR+yZMh8LM/zkNyEC0iOBnwJQaGYok/ocIU+YIhBu/w9Gb8SYszud0
YWXyNGNvDUav10WseBZy2Zm40VeoyPu/leousfUFIdYunuJokCqo41rPnmJ7gUWc
5IdFt8jxLrHxqK0nsG10X0BSFEBB5nD4PIPZlVcpX5gZfe0CXHNvSgrWENXa1j0m
MMEusqzDx1h6vfWXLCuVyMEFyX7bz6Tc2yoWX6y6PtqwEVNTAjxkNNfxHwxdXE/r
vaAB7/V2R4pafx3eiXptKp9B8qxUXUd59FDeZrU9Jpt/Rs2ige43oD5CfRtbydMR
HQTif8lOU7rC33cC3eA/ekKwzN0Ocfauqbp3Fd2EGe0nHFnKE7cYkNhK8V2aFCzr
QWbRDPDH5gDXfgwklQR3lgktIjp+sYyZzyPAI4bpkOI/NGu+HcBMHh2P/mATUlq3
dEBzhhXRF0J8Jf/V19lu7u4/puzhhILUzZFCb/tyiZ3Z2SVYF0jrXFfZlRwToMRw
2Q+zr3Xk6s1HOHuKazlHGR+k1PZvAe3jyKKJt+ZOXTAoBVBHqFv1f0YttUkhigTr
sLOSXydpAD58rI6zK0zYq8QS6jX1Zyp+72v0sN/LsOBGiKb3CAlcSg48ZEALBDcT
xDzfrRuDDjgZr8UH68CpyJBHO4oDt0E+el2s+6WV0+nfZnokMevzVAGQsWQRiM0m
oBDSn7AM2eQyQyeDMI35Xt9qNAvifW/8aXjeuA8TXOHwlSIZ3Sp38WOf/4rTpPbM
FSeO2WxirShy7/ZREACbVhApwPwaO/0+Lm/us3qttM+O1Kv3MLETejUg4ttTyB5l
XkoNcZyl0hpYVK9QZoAzUrJCztMC2QijerfT3VsZH456A8lzvNWmqxTtLc0i5Gkn
7HiIZqr6Qy3VyJcdMdSnd0dJv98duYAkQzW7h0Mp+q73/h4vcV/yECvms0qUOq/0
1lbEMg9uBWCOhrgqMSi7HJVZNPTPuVtcFuID5GS3p6bJIutOLRApncTM/7IM9ato
scj/DcSOkQIfZkptomNNPd4oZtY+SqrI9INpIebKsiQz0OyVQB5nfid1xSW8Hk1b
VEPEX3qrnACR5XoPhZUiw2DWaIi2Q+z2ihTtWLIuAL5E3OcbDnTYFM+S+0wGAQDO
EK9Efk722p3+7YukVoz1h0FxdGONxLKrXphuWi8ZHkpOnuZyl1mtYpVHoEo7aaui
6cXOCorl7GpQLnvHJQ3zdL3URbTNC7lBkt/G3Ssg9NDvW0rPiWETizvT+q2lK77a
WQwoVfrHqljIQNubw9ewmqawA48Nr1gFqgbU/g4+UIBGCUyOB0UZT2wZo7iPYOr6
pytB7TZMCXJiErvLLgkGN/vxCfcJ2cY7hteaVl/P07ysHgnDvsXvLgkV0iXh1ZaR
/oT64pMkegZj4XQExJJxajT/y6d5/epfDrDPqaM6o9sepU3ocVkVrzo0hQ2sw6N+
xh9SejW59L3A1FRB9PEGnr/JxZiu+A7Cjx3RmvfhgLpHaLhrN+oYb0R8GKX+uJOZ
eHcZ0YhRJ9KJcuVaS6LwDtu5s+6mjNw2MZ+0BRlV74ps9uBkK3JLca+kM+lgZj+2
G6EIUwKsxC8/Z1XrRCQUgQSvXuZ7MBagkBl+J4aSdbgV7CUayr0W7u6DdmsD4FPl
bskyALfEJEitD39/jSKpWuDGofgj7dsKQabe9aFX10KERJdzd9zhWK2b8lPx//VQ
3AXI4uvAY/FfywiT4J3ytSqPQUNtuudon1nAhtlBNeh6KHkBYmcE56vrziOR8CtF
z9BotbS/EkbvKIL85vpEO9nNOT2Q/JfZ7Jh9XsnRQN4f07UXfJKa8uenrJ39LEsL
Zzpt2Wl2u77kNu1K/QEq6dfUgn9tzOFSGGuJacTPu8YX8bE5DnIPaUVA5EEu7qsh
qbjeRMqHOR8LrzXYWydeQBHwTNUH5VY9/EvN07Xf+bX36rffqWlH/f42JTJ4HO6M
T6qp2oWJMyQ6TtuVYZXi5IR29W83+aoHElE4EiFC+XE+l+TZX9I2sEoMc7wn1Rg1
9877cA6a+S35JaDYA8hrMA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ILDEe79eVaTIRFp/0ixw7J2brBPtU/jaDIeRfodZPWx6d3dWeNuIvQLjGRKVTtFt
o7oPTK4JyTQQWpmRSgsctlINemLtldp3yQqNmluCMEsU/juhB+TZCB3g+clceias
Jwl2JS2a7/Yp9VPAnk931NqC/8NEWRId7kBSfXGPDQCJTUOcncBHpmh6onFvB+N5
cYkPRhUQsIazOvdnl46fCc3TYPCTGzlRrIjlrRiBAIIVDFZwISATadVS5lCrSmt2
z7YfgyRdqc9DRP6oKKL1TxWq0r8TyeXCP8l3uX5AHgY8NSKVjh2ETwyTXM+U8NFS
O3rNQpHKTAcHWNwGxNRcIw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6560 )
`pragma protect data_block
m+rQ5ICBvzsdUDSAwtSnnQbGdI43fhGUj3VQpD/OkRYy5Ez5QvrZ/R3ZTf8FVAKX
1vl4ZYMAyH1iNOvSc7TC7Vvel48l0XEuIf4/WB+vmb2CewGp0K8Tw4m54qhH75HL
Xzg5GGiHSMeOTKgKGtJjL2y2cRmdeB7VAWKNh1AG4fuyiXN4Vrr4MKtfUnGw+Rp2
uQ7BlTjYQdTKaIII5c/Ge1Eu021Ht6GqSuvpkxFLDiB1wLggrCcBQf58FMTdJMRd
PCn75cUlaAHqOd6x+jiObxwi6crwSHfCjBFqRmy2grLSH5vQFyqSyBYuSmYtkqKU
SCpPhRJcLU0lkAM2bAR8Sf4tiBAX+3vWnZviwEUL/MwU9a3T4FbPPd4OUvX164j4
CAZ/ojWHD15ycApIr1jFmR9of8MOGAxniEA3OTe6nPpK1pEodatLEktNkoXKFoLZ
wfHvr/AUdD8W2eOIUsZMWI1ySGzqCF+QW9RHdr+5TbgXNUbTQlOZcMMFEH5EN2gC
cHq1PG/I9CDvLFJAym7fwqMn32arFzWi06j5HLUHn1aCvvanKtxiXu2SH+Uy2teU
wcl9Ggh+Ae5+j/YzPcX4oM/0uRJyOFBOHVtbdTpGCDbxcLnNfIw2Sxu6fJlais0F
BKByGEh9maBlMADWVOVyA0vP+LLwF5GIma5qI/w3qtdkUzDTIBjANJNr8LmhPYkr
uJGWgodXltIIXCnscxOmt1EyPDtkKpH/8CqKae1xHlf4esHgqspJ8X17m7XBU8Is
wJSfYfli09WX1ptxiB/EhXJV9eOMSE4a4874j+qQLplFh1VEBNIsWqnkWXPAeChL
wI+Ar/4CZQiWggNsbzCvPxdl5tzZ9N+a1AHIVNWo33gPpvJMu2RYSJ3joHlhuBib
GWZXNzPgsMCKJZOlDl4aQlAJlaASyWv05QWdSVfbNIuXHB7mzrN1u2ogGy806/Hd
ru/J9fQxhLTHlpcakdZIFJ3klw8wB3OSckdzz36pIuUnfYkq/Hd0bn/8HciGk9m9
5tJCnDdnTRIa50eHmE1y4a9bkUnyOPoZ/FD/OOShdJmuhXV/ODC7cimV4NZgZgra
d0msQnw4iRktA17GsqqFMezZ6dx51hLJTeljE2+l5htsr+CPYbhmIZpVjiCAc/yB
iF+fh2C7wS21E7ysyvc63k0qe49JqnHXnwOut9h7ZgeqfWpw6XMRT3BmHr8LZo2m
ofuPHkUFQWyb7ezlM5D/Su32YAh7a96yej60bC53TcFayZIc80FPBdH73WpTtVnu
/hChuRHvxLNL5VaWZYtn6kLWTOGh2mHCi19FJ7KRFJA8ksWnooQgIlXfBd+m7C1Q
aL7RzJS3xZYU0hb4IcXC+5g10wzpADp4mzkDyC7q+wmTdTK3NSnviaE7OjDhqTzb
nl63oBdTMB3Rz/uqCPGNa4G2H1Pfh3c9bP71Wg/m2f8XbXwZNaHJtnqaZWFT9iBy
02vBAX208YnpRy98y7g4DE7I/jhVYlUOmPGQhkwJQubfxUaokXEcRKvWrQzt2QlU
Nlzs1Qj9020Bqa20w0xxgeOHpSC1Sg/c7AgH564CLqSiVSJGrDFvFvuQhby2jH9J
QuBRpBV9aVepsh14wkNzSU1p3YxCJ3/M1FX0j5QCfq1hFdkxOF5XbtitsBcQyrHm
O4D9IdpBG7S1t6FSXzjuGKfhjDuN/YWLU1slOdQmvcuf3cjVGlcAfqSyJp40lGGk
ospqinz9o/n+l/pW63P6jezGFVenuz3PQ3yG67FF5cio1p7VDdzgr6R8BlvC6Du8
Js1SKXaPxxaM4oXI4pglBsf3pPsxBUwGntGlqLDgy3h1aghTJp2bt3w282VLjwr/
rkR8cTaWMNwu9/eJ9lKLMFDycqt1LmN4a8tvJ93S2EJbaXrZXUxr0HEmojwaL+vE
BD998DMsoNJ/ReA2KceWNR8KBJpf9UjsxxGSKa3b1ToJCAVC5VY67u63ZHtsIFnP
W6ElNtHxEP/Ll57QoJklB5GZc5xNTMD0kigJ7O1cqZZdOTEFbtzIrh72Daur03Be
9SfVyC/GiTogehK5q5NNOo3tm8F20pHz9pEMY4IPTn0gAROtARlOFt6vmVX06TML
ulDhrJQsrxfvRR4SdiUQCd9Q5hn4UGXy3N0UQ83484roGFi3FFfjBv0nmOeEkdLX
9epbdaAATY/KI96vNveBAEHV40GIdUKH8Iwo4Xbj04ePgxMv/7H/ugszRNoKua56
Fi+z3usjqA+Mx5TXaLNvZ4DRq+1UOFqxyGMDiGtqJEL6G1Tx3H/kgqxrZzhsFPHW
C7oEBu9mhUnpmmz6IsbaCR/cK9W1a0caHyrmHwvY4s9AH95Jj4RwEZNPd5ekBDXQ
cFs5QcYLVWIrlcl2re4+lBs696IorVByhD92HfOloKkobVPpPS/O085YRgtiQGtY
Cqto5fM6rqVHSbsXMuSGez4MxlfOOkRCnayFm4qrIZisRCSl/xUnCOmQcFlkMIb3
ga6DJum0IVSTN47wMOLH63EXqIpFjjU2LAbmonuGGzCO6+PwmfZiHhIaTdEXQUA6
ISnCgJjM3Umi7WnaBrjKr1pdJ61boOwHl4T1/SqJj1TXxoGl1E0OuA3tHcJY3W8i
GkLvNh3qnWEBaUmWdnMVyKARsaWq/mY8JWkX+Nw0OpO3txJ0ImVLUMYl/IaZPuFX
bUu7ZexX+KQv8EjZopIacCW/EuH0/Z1Lrha8xms+bh2vcwFrshP72DGPeydmwnc4
5Md/mA9tDzqp76m5df+4mMQz8fBZ3k/o9L6q3DsP7iXutvTFzSYtqBAwt7GIFtAA
8cQa8fFzvK3QH1RLaDhwUhbs7hxEoH4V2p2299XboQgmFLUqVnJYu90my+qB6uUK
ph8kDDfAVcsqu2hwowKodt5APeqnyb1jyWH+h28Y0zs4/ZTj0iVhQxlM9Jwq21+u
u5edFjy0UoIcgsdxH4tnkZ7PCh1bqH9nYZ+Rop6Yd+3y1asnSmUW2jg+a3xO87Xh
QLJ7HJvCN11bodrMBSDCKnad2JBPfDks4dhMSZAqruuzRQaLSX2OMki8XVFR9+us
Nh4qhdjLfRCG3V7Bdk4NGnJOcqxrwFKtgRWxuUdx65AgbF8fgNcGrCbQ1SIqzY2g
NHlJPzK3xGBjx9g82/4yRv9LjFwpp2vCXyG5O4M/gKHk7KVguUzamfEqx2NQagL7
RZE1FwWKiojtBV6kAn4MjUFV0N5VJjBZbWvOyXHe63xH4wyLWQXnWIJGV07sJ9m9
FSyAPgiBXSx0ik9PF4lP+pFaatp+ttqxCUFFh4JnHixmCwNoxpLB3+Jn99ZXCw3c
bMLn+AaJZ7u4IiJAp/XoqiLL7aUoSZTS6LUHVMyI2Qf4sggEVYvZFVt0Y9l+YD6H
qm2dq8WQxoXef4dIc+1mz1+FEBVHlfbzG7lLC0KdKB5zyOrmPxEu9tnDJkMLFqmV
A1ymkJ+jWqCvI9RgNSqBX1UrfhhDodyz91HaHnQJwpjZdLxOer7ATnlqpBJAEso4
RgCTh9xFxc8dDihRp+fetc+44XeZ8N2l6BJhfl9O8Mt8J7/jVBztOWfH8Y1s/Q82
iZV2JDqVtTqbTIhc6RmAW2rLeA6xbELzQ1dhve2ZgXFXzMG1m7glYUdSM6a1r88D
ZhNH+bxILFXO9he+uruxX7eq7wTplV51hoDU83vAqsvoDsTKyymDvAzITC2RlH+o
DdkCjp/GDmtMiKBbEtMHMXbyfH5C3tgbmwfSIGphKm3H5wbqVcJM1/cuaoGQHOPX
Xzv9VPRRsLOmQUBZ1/kAuUNGg3W24/RZU/6cFUJa4QaVJgYIXBoZ41pDbT7lGFAa
BYYvo5jPQvIUYeZS0l4M0oAgTXXO6T5/wE+F5+/nVVaMbMajuJDZf7kkgVBOjoaK
u1h7rE2XeE4DtSG8Me/4hyN1suLLs7QhHSswYCD9km/HyCsns8AACQ5VnR131zzN
U7hF2ltbMkMmIImtxJyKTisxWEEa7o6b8Bs/40RcL4BgYftnjKMk+0O/FLG1n0jy
a18J82d1BANfB0568578ChQc7VaFgLamuxb2mpq/nwvKaTWNsqTIVlx2hg4fKphG
vvTwwggBCM/hjJ1Hf6P7vxa1fhRnA4QSnJaEaobx/sqpK2XmlYoV96C5HeqHcgqr
e9nGpuLsXwejMZ7rrjZTUN4mnooHLu1JVSoDhqOV7l7YZL0Pyx5w6ECAPiBgusCw
cj2XfyDZ46U8XHRqnwULsk8HZaSH6GRv8E7R6w+P4evUG06wdcdgXRzE8QuLH9Ui
DsSoWf6uGw1x2XTXFbD0xHew9926sY7MEKzaU0nDOTBg3Y6mecYLJqeSxZaSlKM6
/YLWcUEHH23IM5rH7C4nz4Xx7FgdzPdUZx4CxQIUY1TpFeZiFtwXQu4K1WVYtgKd
3BmwBvkxCdna8FdW8lNR9U0jpSVVHyeeQ3uoLhtfFMs3lkgnq/cgfY1QNUE9ZISk
/Ihdfb4Qx9837mXlz5JcLS0l0kZGHrGEGpFgJCP9o4bxOWGH26vXZB1bJZPKrteB
C6nRbidmYWcXpH4QmDPvOkJ8zopi2sTP7bENvbueWrvsyM3sEdmWjYJQiiwqTYrR
XD5VFHtjPOceIEChv/ZkzUuNyFLQk3cerdgbKUVBtM8+dAaR4vJs/o8Cp1fW4Sr9
3PxdNNNEpgpjlPRc2T0togC5JR8jgbEXi6IfpYsiqboUXzpoxGqiTrBmMP7dX8BP
k5Zbd5rVX3RaMD9RLEzJ5wzSUUaP56HBqmDTkwHM7RjRSGY73MYmDLBUjRAejM+N
CuFbe/2renvqeAniTaDrq9diRi1NmN4iBkGeuWL25e38M6rJgDvF/xX3H+7fSe9A
RjXaQ8Zz8eyJFgPhu7rcF16c3QkmR7OISGghWlsvUd9/cUX/MkCzkrC/0f0oXwPX
TMDx5uYQlOK5oWZ8UCUFsfvTAvOZqc2Uwu5GEMgHRQkXeXb7PaL6mW8nNhtI4tiA
xNsMWUiQKjT6xHGo36ad8NuZaKYhTrNGBiht1cevTsnb40/tA4mNCIL9RcyqESsm
CLMFOAfXPvtNCZLs9ITDqPN8mUOJdPWL0MoSLPs2OtxeHxojIrhfR7fx/mdyHBrd
SDvg2rNZkYuNMHdTd8CxXFtcP7bpNEljMmiH9WsuDdt7pqnIcPczyx3kmxnpy6jX
vNJLzp/yI58orFoC0NKzipqRwjoo4gQa2yxfXF0j621yDLCMdNqW4fwMZk3UAd5Q
81iskz5qiQCzMIMX7jDDzsB4NXAnvWBflazRImMX9LG0S9+hhDlaRxPJLdvP7gJe
okcfSPvvpfwEZQ7XZxUlFlpsXuE70ZHYE2w/aolyRvNABmWj3pD3ZK2/JG0b3Nqf
aXi/K0O+XVJDJ7vvUsmrrudFbqW3eJ7c1yr5H9q2/L5tAm69zvlbMHh4L4J+wk8W
m12h+ynVoxAWxCBzgx8RmFHcCQN1h0mBDj2NjtDuIdIgJZCczNrV7SpcuEIa4cjh
7ByJcwGqpkIC7l7T+7ujlecpp4mof6dU9D2g9QRQHXUOOOUGHEJv3CL+mnqdo7Xw
linwCLWbTGWNxiEsDhYMjY1f5I1E7jP0BBlxgUrWygb18v+kzk8YLJJtvMfCQ6ja
qHF0U6lI/ryIXSpTG9Evil1WAFnZi/1M2+gqm/wMWa/7gFBmnyPdTbQn1ZJULntw
YOWpQzBmrp16s/auTqE4F8WhV+eXOuObZ2KfZHnjhnld+qVYJnW8QmLCJg9GDGQU
5YI6vDuoc3woFXtO3/trPHapdf++jQeXmFKXzo7S1oBLMBhacLR41Vj73NjwrFV4
piKnpw+XHWAclJIJ7qO53VaDXN7o+pxVZPKgx+X9NxZVm0BrproaKT0mabXNMy0j
bXGZsI85jjO9ymVrR9nd63tx692Bx7Bje6kB6bAUKhXa9XZCqpFl7TacuGbAdcha
kgbEIG+dwcYVp4nSjo4B7PC/Qyvf4rIveVvGC6nl258/jEzJv1giefb2gQplc17V
xU4Uu7KxtMD8kyeNU2qisrc7kjuS9gkuqh6PpcotpyM3nYlG7CPy8sf74MEfelxz
LwvN4HebfZjsl1jeHjVpZv9XB2DxDtj5osQm/eMlQe1MKYAyMM3Rqyxe+UKBRtNw
gR0K6bu0X2BPcn3QQH7okVObhhJtLEN3ogaWxPTcX97m7cd+HVOwvxxZkUNmV9CE
4PaWCtTZpMTKYAKPiFUOohLhVTyqn3YWLlT1JuhIb/rF2u6XUKqYHV+r3NJGQxYj
99lgNbFfAS4mVXPsLeKcLGhT/F1flyyrpUCkeTEGQ0CSdcfyakxv+O5R4ksKcgnf
f4336EsfCZUnba0GP28qZttzh7kQ7vC4N6xC/XUzw/6QmLiMk9z+5avYg4PW+QDu
iLZqwY1OceJdfDWfRSF0XizXt2K3pa0SWwXEKCcx4DujgCU5kQKz2C2mOzBxzfdG
RGOBverfkkpWvB06PtbdZKTqcM2FzO3rt9PwhRXajy4N+NsfhNx28LxDDj5lD0wd
jv4tTQIVDW2279iZ9aGyp67nCYoYJT6vXZJICbWIGtdPxx1JSFRhn+2eurjSDxGt
R4+S+nIDs+0xxHYHCwBLj9EN8Oy3LtdmRtM5umwKVU7Cax7lG+SiiDLFYrQzcFBX
wO7QeJRNNTU+Xh7wea6rxxosyQfFbJmMayG2hLcGJlpfDm3FxojLXp/KwGA953Xb
Luj4isiqY7h6GK4iE0cGGRpmH012i5n5K66GsnikXWk2ADaTN4sqJ6RpQ7KcQLJ/
8Ia8ikpgHT3e+NDt7u8AYrjIHqmUCuq8wAtyjfInkvm2PilVsCkqKNQ+olrho/E4
kniX+xCufnJOW1HTRLuv+EMfygdrRPFhsdsV4KH5Iav7K6wau1p/qmPgV3IdQFLD
GNwXmJJXJOXB1xFQ4lSQK0bTIATXXpGv0O7Vh3c8mO2pMUswuwbEQzCxXVfxiN72
tNNtdfp5QY9RgcB1Wiq21xUY5aZfyM5hahkgICVjbSi6TvcB9IF5n9sCnMrCgxhY
OfBatL5g02G1BtopLQT0QMjwubuMAhEoy+Hc9LbgDxKS+uNCJOnfZeUZlNDRYOrW
vG6jWMTfzoGN+pChqnUWZPAYNe7zJTgJld8A6phP6s1XjzNpHCKdBz8x8l+IuYoj
PSF/rUOWpq0wFqq2Rf31DCkGf/KToRF4ztghurkMqwmNrY7lPlb/c3sy1+cIZwkJ
0/D7BsBLzdtfb9LGCBJ9K5vHCRnqadqFuP2yB72h87SI7IpboUu8JAuiXj5JAT0K
g+5uQ5QbZ+eIqEUGdGzXpTwVXgPAqHUqn3FelfHswCWur5KO96SNfmDV3/n3BaLg
h9bOGWMxI6+fRAP8Utr+gF3z3Lnrv1tQt9Jqo/6yAROTJSDBak46hasKv0qzFwOZ
1LGOl0NDTXFC7tRbeunWf1F+7lo3w6gWV6efg7E+IGHQ68wl/XypkQsbUeRFYIRZ
Z+wvi0AYM8Upf7oUeBvq4T9/sUaF7WtswqiLreL+u1yJzqgPxww0IA645J+2fSzC
+6GmQSrfHFeITyMwnQKVhplND2WXyJVbEQXBILer1AW6HEbjhQmYCPFHatat3FBv
TpkmTVFQaoNhQ19qgsOD03GakIPrBy+MwNHqD7KP6YYxQIVehmgAeAgZzLdEnuub
HSPrwP2RJ8CecgVe4AylYkqu73lxOX0vZrp76fg/rQTFOPhWDaxpNSzGfMzCF4st
KIN3mDPPJMMhEnNg6UlmuV03GijlyCWvEVo2xLPCBeQepZtvF37Xt++ZopocavVa
qt63LvBQb1N+hWY6OR/Hq1J0cscJ0XhLIT6wN0eCEPDyXBbBcJrSSKQE67PAHkZ5
v7I5IDMdpktxrD37/k/D/NSI29GrNf+YLOh1mRdee9NBAiGsvjxvmF3pkGpe5uXL
yqJ9Xv3QpGclCzF91h3/vpxQuYr7R9rfLcd+kIxxDTFLhTxcm22SeocG3UaGY1zm
mLdJT1SCY2SfJSqulFEJdkycHuguvs7N64W7s4KalaFMZDlEyrB46X+gymJEt01n
YVLE6prPASoGT3Xm6cfbwtoxw/CZlLvHtvjAuZhMdE0LIf4020mTzUQkQ7GXe1km
48gsWcc/4cDW/Ds8bSOxNP5H81i3sMiGzqQy3NcoB6fWmT30Bbdd0afqZG+IikLZ
A7m2vG+uAq1nTuMqi4B/9W1hDKuJU70Zv5+J1CTJEaqX1d1hH/KovYC1gCGJ9p6r
MV4IajldUV2QbztzSyr534834ZbvwOStFDivMK6oFw30BN8UOcK6cdaWIjsUNzyK
SfDXTG5SpHFCUF6ZTzlJOHt4z6S6l0F/4cXHI6IApfLhXSqQ6r7AvAdCw5GwL0sT
PUxHaUnJikEPO0uhuG7ucJ/1UqUwaNHjoq6J+iiUgKqhie7UeEwP03+SZp26hfbN
urqROOu1p3b4wCKu57zFkj7GwO6j3OOGDPtsagop+HsKNknJvVvzk5R5r64myd3n
MLOGq94fFZtVlRK49u8hcXO/7hqtDeYoB6g11CC9xrNfUVl+nXvsoNylC0Eqw5oh
lQqYtg0TbdWVfMkZ65ULx6zwTMDuibKgqOkfNQJYoL3m26DkAO/xw/A67hNyX8JM
rSw71ePLIoncWKOHDe0cqwOnET/WOxZyQqLcuqvPnKS80v5Dat/6/9j7CFr4d51d
6dYQQ1vcas2DV0MGNCFpAVInuJfF116NyYhRwO7xJgM=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
XcR4ZZmoT8iT4Nx/WZnp28HFuF39qMBHwfVyGZSfEQLE7p/guYAGD0ufCYI99Lta
quddR8feV0nV0PMGlOYLU/h1OqKRM50FByscPKWZHmvUFC+Rh1RWLJ+qO3yg5dBu
XO6bBk8oHDX37SNcJmOjryZeF/YSCdIkxzTTjrKNYF2ASiO7xsDp6RhN4CN/Nebg
1k0Xl7TpKhFSGlF+b+JnxUt0pSM9YLlqNLugzLcwWIKsfCC7osx5o90Iik97pMfA
U8G+T9+V2EAXY7UZRD/qxNvTvvfxL0ACc9XlPuQ4Kww9qBWvOB7vT5oY+iJVIGwM
X2NbGp+sg5InHvnrv2WbTA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8928 )
`pragma protect data_block
uXlPPI5ZHtoz8QwVVGW5sZyLZ4Pp5Vi40bHx4YLhmxHVjK0RJrqhGAbIbV9Ot/wy
rDe7yvuEi5FHtgaxZT4xm+DGDI86HKbQEDfdRsv1YOj42CpWnJWlpqplRkARWsyk
IbbMYhbYG6faunw2LsQC9fFliBgQ7XYDDELdcPJlK5OWdNGNxEJEuXoLRxuZaGgQ
ENZPZs09NFYEgJD4m3g9oEhyersRCRnQ0uAHDumyIEmTUPVmw0tN6FkGpiHv1mvJ
aMmX5HZ4i228v4z9HZLM/qChCVNRcTtuwZeijCQnjl/CiDPXPRotruGK8dibYhok
7QDSk+W5BZVdUDs+y3VTPGb/8SsWBgYjPI4HeQ4UzuSSWJ6KDv1IEIZO32Q430h4
sIwx0UXkrkIsf9dbB8PpMtcPd1uWnSup5PFoD2YYlpLwCOThbOFqiPOqHt0O0Uq1
tg61/HZxxrXWeH1EjLuIeUd3ShiCx9hENsgB5rFhpeH+fy1SZgUKOjMcbJL9NeE3
GqbmG1rSGW40yopKp8Q0QGxcCDYuVzK5AEU9XiHIka/+SYjxQaJeOZpvY+AFC2w8
3qhKfiDa3fAX16wCdkNW3m4zSRMgXTyn7OroAU1Yxlm/UTcS+1CtzPmYFhgOjiqD
VM9a60dOrfN4i8rUAwtz+Wiu95UGBwH861FoFiVLYDF1T+sQcMhUYvIQTSTVXfCp
ydr/1Zmet2ZUOhHj4ZJAzLC9hwttGp3pUBHkPU2nA29aWVqpIctbT/44Jtevwo8U
rwsjwfP0Vp57uwVY+tbahQc2NlkopLG81MF00Gfp5tpKjfoERr34s8WbTinPsTNX
DyFypZ/aHlT8IDpZYW92jvLPlXikHxrUn/j+XvSsagyGR1OIIYN0QwLVmYJOqh7A
7qKafATJ9ok7+4jz2VH8AZ61QpjND1Xn0Vd85NNTzKqHQPmQ+1i5fe1txf9RsIVJ
esmTO/oTUtSQCsqcdVSRXvCzVAeJBwIAyi1G45ulQwDyZvoDKnkBUTpCpOMlDhcD
TeySkwBgsJ+O8SZReeuhwaj5QUjTuAEl07h32CQyXci91xVl2Q1WkVtm8GARVROs
StxDSguE7p1T78o4zIMO3cy7+IsmF9LMatO/IWeVZWUYrZIdZbB8g0jTZOPNLJZ2
vsHJt7zT99mHUnvtdmdwDC4gRFOIrz6rZ21B4Q4VwJdkPg+oFizIo1vlnqhtmtJc
+NwxhRAEvzI5K/ecLe2axXgUs2PBUyq8B9GawZjWNW9yfJe67q3Q7dcGQwulo/Z1
tZSnYowyGb0gE6JL+x5jPxQKNhyE9X0+CcjRgU1+/HyGZo/EUUrB4fmjhTA9EAi7
FCOn0+BLFHLxOljXCQb1bjX1qBLxy6Y+zVBDncRROsKpfRnScNqSPNHBmpqahGSV
aIld8iupeOKW0Z2Dp84HVu6bEc+3NdW9UDBZV0WRfFtDuFTL/vBZuWsFUVb++MFG
nzlkAsBn7x7DFJpyeMoc34WdHoOGbLWPUeSfIXeLoznAL9A+a5V3egLlZ+Z5SMrE
0jzwQK6BIYZkHc5qlsqz5wnRTki4Ar2kkokdRBRQTv23ZJAylnb6br8BvoPomTQP
yu0/2/Dys7UJV6UUyzCS5IdyqaoPVdYUfWT1bW7DUYRzlUBdSgqmTULMtgBCbpCe
hsFYjG6AphetQ6fFEwur+p42chgEPbdXUWVixv/NOotRw2bhsesLr8cjgpWiQaCZ
nOWAu40NWZCaT1e4hVsMqMN9dZh3E+xQKnMLd8qC5t53XWRPTxZd8uKZh45GLdik
atSsA3fXazONX2pQ20Xz670kDLbV05tqNMc8IAkpFmSR3kDNFKkrRzqN7S/VPAiw
p1lMZXo9WgfppF3RQq7g6buJMnysOiYlWHshYygq6c86GjDLFI057rYteSoGpKH8
22Rq6j1H707diUaDFAwHxd42ozO/ug7LTZ7d0NKSEdt9ox7mJkmIJ0zEJGuDGBgB
W1qNj3ovz5a4OlqKH0B4FUpdu7kbtxjObW+2tRAUTzdQUWTYBieXTrajSk9t6fWx
Z2vVac9zstkKplWSVhc88FWz4Nmbwhajz/FyVO7q3nF+M7orUYT+i/GUox3L31ak
WtnSeh7NOy6IMBSAr2EWBgOuZehFXAHF8OyXUnXz/JPdgvBxttzKK7hin22Bz0KH
84dXyu75g8vX3Vx+E03gyOdHJ31EO8q2k3u0Ap7y73eRhyyrFhXpASwBpQwORgsh
I+jkXoWMwLy4z7PdWMgegUibRZoaHG20CVS/wN+SXqj8V8ifK2EbrHJL8DJ2YbvV
oShVqJNWnlUuJe2R4sFs3IfMMMyWTXjL1IkmR37T0icHFWkiOtL5ACL43q+5KylI
BxM6LeuIgQg1FA8fNMGInacGecKo2TqJFDzBdoaaFb0/doPGS7Z2LMuFrATkwxRH
nWoGJu9aKk7JbE08tt6Zse5Iwz08BWz4j9bPZXpMBmJSWfL2Tngg1068Lrew8AzH
3aYHx45tBluSGS08wTfZRwdmSExNqe9rq2ylyiHK9+01KTtQ2apCLuTFawUUvIkm
fKX6XVhsYcwYtLo7K8U4B9RWB0pvZSmVSvwk4eg0oSJwemOmqBJs8shpnoR6CrfH
WMhDyDLDKQ+MVFQ9+zNVMq4tokM8n4YLanPG5lmxNwBHA7N9xRUieIjOTbvEtZst
3AhJU6/KvPw9Ya/8X69DEBY96O8MngsTUTY4UO6sp5NVWVL25lQcHN97cVU9Ql8r
b0OK/hSp2eLa+LxyIs3IaFqPWasMCSesvrD3m+OKnpBfaRJSfzh91OFl14AGnGnc
j4mgZSlTXRvr6DHPQ3EhM4Njnem0VIMIcJzcF+XuwbdjSMA1HDAW2mdqKUCkUPuZ
a14a0EuxLoO6q9SyPloEU6Eg5snF8JnQ6mpOFurTxKi2POThMzsPl5YZGBBcsC89
nAs0E5WN27nCzozJYaWPsW7CzRddiXVikLvbidPqvIcgJY6bmSncsBU3g59OWK3M
sPHBtXqyN62oqZZQJoJmQHF7z854ESdqZHmdII++oGQo7NkmE444tpWKK0mS2n9S
+fWcXgjVvExJuUQwWfKi7JlatCLwo73Mw8RtbB2KQSj1Zjgxmlq00xKjje4x/GoT
UGWfLYToJzB/yqJ1oUyJNT9D5cObgln+P6tEXBSxCHKlpOBAkHEuPyqBJvGEWi1k
snjmkkGX49Q+gtsvuvCxU2ptWfpU4GBZ5gRWUzJFb6DQQpjZTrjdUCCUeAc2hiAM
mYXMD9vaTWmje8GDZHHz6G15QMB824nL1llrbttdJpubc7oKcs/zBoxFk0F+EFND
mpRCvsIGcAbd/IQ+Wj6ZcCTFEsf2E3SV6D6v17UW9YmAp/RVEec60eOLMXYuljk9
U/JTn5D2ZkYYIRxjpnxUNfDdzXSJXYGRC+4gIc9OpKg/n+AVoAp3d7QGDYjos8Up
HlG5qUnuaTT0l5AqhnHdX2R/Z/hjB0b3J5gjip6xSOFkhcs8n+4saUtngfqEuDmr
o8YuWwcYRnBnW2gp+mJrTaiE9mtQhEewbRKu+1KBG9lfEKLD8ZqXDBUh2Lr4jkrQ
0KsNJ99bRHGxhV5tj5RJCc+kD0tjgy4sCJyjpq91eAK5iU6OxRHQg6Sv49olSxJN
1KI78Kn0cV/WQXti0hJng3HUUd7DzSd4RiQt2U/dMlVgVascGji4DL5jfW4M3bSn
DmGY2tTTbxvPsLv87Pou6QilHPPlWzBKSZdix7W0XO8+dn4F0Yj+oMmSRVhLxaSJ
uHSmdBNKkC8Pm0cGYdKa4ALu6x58c33KDp9yV36qzkdTrl8iTkV7j67rWDbxX4ma
leFOExWBR3mloRKHXXGZjYXdM89q/AqOsu8+jYL0m8+E2KpGCM4Q+ACrUpZUAFyk
jeRto0q3L4609vg70z2ly8RkJUq014SMBu8Y7MoiY7FdMnRvRuaZCGWgTS/ge+kQ
+QE4wNpc/US8qFbRJrQbQ6oj9Bsac9aDPX1DdqFlFw1bY3bW4YYpt3W2/NRtzIPB
S4xBjGPZHPqMIwc0d/Ln+dKEaJBpoS9u+5z0wMcKvyOvr8Pz8KdaIN1XBvyh1NP7
r7KdbI5QHyDMVFBvIuMeRmOwXT3Vwn4G/YHo1tGFF3EpCJCSx/ONQaKBzh1HI3e4
2zGAY+NQhsvbNQmy/4eH9Mu6jbEDL2J9zJnETRNmiyDC62Tf1e8OE9HvKkHUoqmO
g33OzYwI8pnOQSVSpKbXsmaniYNappMQzrjapTj++QIU2dNpdHmrGJW83eoCCP30
BiMGfBfimuAl5HNPy75ErO6nGTn2eWsOsNlxBSXKOXmCEecDxFnjQFW+HixDXlH4
dJOcDM3MjnCePPazFq4Dqpk10uGjcjXEm8hRGDr+4N3eBh5tsJQOQVW6gyZqldzE
UZjNtPn5lqydPmsDEbk/r/8g9NrIXFkYyVOPIQXaY31nrtIIhV6JqAk2UqiVkngn
DxmBqJN2cIMkZd8P9e95diQC7q62zsi3eI01li7lbuyfoLzgeDxawU8wi7pjOmYs
9+kL97ymfjNaXHhl56sbkscP1tPtw2ztyckIhURZpPXyh0BH8bBOVZRvRY2H/63t
TQ7KZaqrqoq4Cy7Jly9WnS7kRPR0Suh6Ge7D0s9Xh5NY9kVim1lbuFJwRRuu7xRz
oK5tHyY4BC/SJoV815wlgHsWT8S63h8ENRvMlnH2kuphrnkPQxaw7KF6Niv049SH
CyB48sWROKOws2VvWxs8Z8Jchewz9qEs/oZTLLgA3YNs0a0qy1iSguZNfSTjszXX
8iyqyvnfuQmaI9tGBWtOlvQIbhZGrGmXHwNRJ6x3N0K4Lg2llnP6ACnxb2B81VZN
9F7BhIwtsTXAS1xYSLN4kFkz0uDUVVgPxHaKCDK3S0Gx4xSSM0uvwSJOBRwyfU1r
8AF8ZHCYzdXwfW0Od8J9ByUcMZoUXE4n0v+GsFOfp0QuE5ll6Z/5biGqKIy4JCXk
u/yLeBvpjp1oBRe/Yi3lr/ZtG/OP36TykxzkGvHCoHkCzGd/0tBy9hTTNhUUKMvj
DJmfED/J8bJ3peAjUsYHcFt+5ecqP2rWNnbc8t9IKo8XQEQQy6DU8NTefAjDLh1X
+0DNaTrqyMd2NKhWfJHAGv6EKMejwrqsnti5vWz62Jcc2MqGfAvQMBxeBkYxBm4l
DxropIK1DLYiMLq6A29QsOlD5viRR+prFcMk07mM7mO9u9jLNxW9CmUgGwptdzyu
ShwaGK1gL/4S9NEvJlPex2ZmTZf2YzktiQPtFJTq8a+lfNQfQlIsKzs9A6WomvwO
TjhKcbttSglTkqIlYHlYXoR2p5+4a5jnF+6tCNknGGklNXyy1Cv9QkrjpeCkG32A
e5ooMK9fPdoixquCONn7lh7RvuH+It1sqK2g3t54eOMG2qvKaB4c6Wfj4+X4Wa3b
bQKJOo8lBFyxebOO8/8v0bljImTUP4qE34PA2M8SVFTj0XZnj4myhrioV5InidFy
AVaIEWr8ZzF1YHigj5UPPdOPRw3BDTr5XvchI/L4g3Pa9Y6+gSZfw4sMEM2ab8mj
tf/wvaM9KjbZVyrHyG507770DbZeYQHnOAd6+VzQue6wQCQqe+PdQB0114Mx8qMS
v/I7Ty+yG7YIU2Bx/4kwpSo3sb1KxWCAw2UO9TDEPAabcyqNx3ruyWG/ZwWBJz7/
UOwpj093iSORxboRDWnlDzj9Ref2vzsqd/1I6TwjFbM+i1jeoOF2O7+Cl6iCrbks
TclDSFWakkfyoy94d3V+7SnVplDUMl45nGWAVTBof6OdUmXUd612dxX0Wgbd2zcO
XJgng31we8X2e/sYeqkCpspv3KFUXPcGliJTCbwdEIaMp8U/Sc3MzT626YapCEAw
1c5eoGtrV+J+93cAjx2QFtJeFsupwHaeK0dmZFLUaRMhEEFn6sg44Z3pivn0FzQI
HnT5UTOhNCUbqYZbdF06JgNNYwl/mXsrxnaz/lRNS2vdMvdDpWuxROtRYmfeJPNj
zskGC4VOveNf2pqw68MiV2noJKf9Qfe65aHk4CU8EIGCIU4gNsVPdiyVORLd5hNA
xS0cIoe4ehEJdfcfxHpD4VL7wpArhqqQcfZzHw/qlIq9axITA8ClgTRO+cfxfSQk
NC5P9HFKMzvCiD1WC2gUzuQ4rqwv9+gglypmHSMElFa98gXq2eRMwS68OSX0K+vy
yo5G4ICvMMWiM/kHaabOf6kMbbVHTwa3Vrry7x36O53Jzj40B+G0w1VwimqB/rd4
Nt4hSSMlCeItZEusfu4ttwRmIhiLbKIcDYr5MZzZtMfH81BJOxjD7/Tri9aJbh7z
AB36a42ppHaDVWbYrjpxEM/U3ZdfIyEdMU8OsDZ8bXVtEbhcZ+Q/ppqNMNBTixlB
OXXBNo6/ecJxGdAXmhdMBXR/WGJiKeZFX/QmCuVzLuifXmEcuSDGCTAX6HTQPwOs
VJ5Z7h9eKpn8Uxqklspyi4EnIAyNsdAMKqsJ8VKQGu9qKjx0t3rI2gwyvdl143Br
RHfYX8QMvUeDBEg0NNUvUdMjX/tP/fqwsyAD1JeroGho8I2bp1e+3kEGcNyDVaG1
JvBX1WMLAzzUp11bxgcgCiUMF+dSBe2eeSqK3HxRAHuSF05VsBoXA36pTI0mn/CQ
nfKDdAEEPph+HP96Hv4of5oaivRm4OYODmUZ9ulEQUF7ZSc0z1L8TVHwNjc96pB6
UkXCianb213EdPNyGKaT6Tq3/+SVCsxnBSW3bw27xKnsxyIcqDUywaSbYO4i7Vq3
/b4VEm+2qbqJBHjrjLfLDCRydHSEDwI8Hc+Z4KyQzpjcNVy1ZQCUAtT4F/NaID91
l4axxwxLJrJ4GsbmgnXCicBXwHTCtQz78U9zURCOfUCpuAq2znt291DS3CtAyY7x
wRQUx7t+nWN2DQADQw5gAvV0ezFLMomA4WN3pl2ZH4eUmYXq6vHrvXkE/bnukKpH
zNxO2Nk3NzJLi9m4kaN1ozLja/0gdXfw26jglZ7t93ztcFwAfiOjd/hHuYOQJ2iZ
PHLKcqMILIysCLz2lCoRWjpH8AcCfLGcUsVpc/Ndgt629OdXZpJOv7QEDhEXSBa+
llbrn45l0fTR3jpP45lTX+llDPlpBktKE4b3t4yKKurJ3/6XDUbA4uBMsjhPxs2P
RPpF7F8UWAzsCCIB+9gLwU7HdLiYQL9LgAVR6coURgcJuepAqY8TQGpxVlq4xBER
Ya6pRDFgOADbpKvKD+vIQEQf2RsVcHZRaILiwAEAThwWt6oILcj9J2v9c6bSX2ri
okyP/SDOj5Ot15iKp9XFBGuYtG+6bmhyIeofNRsodS/ZWG6sogtjZjetwA81LDnw
x0cKfECu9oLn4NlbwQQcNmb/18LuTcPNgYijH2WxCGOkxCWnYlbhWXlnUphFYCKf
H2o6Ar2eOlKyogcWL1JkkOTN51//nRlUxGj/GuY5BDcEEsHRe0clXu85iNyXmt/q
pLbElnRadytZmam+CWaPibn3/pX7z/q/1+PVpAZ5JNAd4mcgewHto4PN4WnJ7ykn
0q/1xyg89xhDl94MSem+37T8exWsFkZBrR3dEciroWegTA+YrzVgdi9plle3o1vC
YXw5gqvr64yhMjAnzMcAmy2Mk25vKCIaPsxPr97ap/ymb1mIzFWAv8g+wyhx7JzR
3lzDIGfuDDIwMwcjuDjXPdgcyNwuGEHxbt/7viTmzZnQHX8IX239Vo65sOU0fo4s
Kk83JQIGq8CKLtPxqPNnrD2ZlUd8PI5S22QlXMxy0G01gO2WDCHcawqhwdRRiiBh
7iutgEKuQcADILzAlsoowawEYOJctjmiQeg1HQaCFdOpLxcBYUIr1VzsC/DF23+F
Nwu2TgsW2MW0/0wVyeNHMiXWFs+1GwVbOxcZ+AeIYW3ILH82FI0XM7lgyxbI4mfO
TxuEe66JEgYpMEMB8yGd60CISpRvzKG3iTR6GJtMRlyY2BDB+gzJzAVj3cGCIgHD
DO3mYQqre7v1c7Y2MtzfpYdx3Ep+DVo/z8J1dOkCPLu8KJn2ZPQSPAjmQ4IjTG6p
3rQJjc94U1zninrBVCWbO2KMOGLXE8zqoynBKSlW7qIeczOYeMmN04Vkj8H64U1s
+o698Uzd/Rp1ye4XWZTOrHp5XHG6sODjr2/8e2z3f0lmngW24k2la3o3OHaeTM7/
VWK6aHuw0JaMvjJayuCnK4/EP2FYFJvPGPMHuOIYmFJEVp3YvXo3n+Eo6g3k6hkn
4z+7f2lC8/wjDQodKt5+9JaLFfvgRSPByQrdrDLW96QG6nuhOsse/woeLFNlonR1
XKWvLiz5QonRMqtdm1nVILAzPJw371k/6eDRAWiluHpBGiMKt4WDgqrNlHTtpCAw
9fLkor6eQdKol3ReM/BViQydoOt0Fo1BmZNsYWmSScJq1UdqI3+sBz0x6Z7sd0oT
n5ybZsnR4C6WI1Y+juFO1Iboh+KaN1OPe8vx1nqotwctHc5Z+b0geSP3/EV+gbG+
Ulhl7yxdJsWqxoH+xMtt7jU4LHMVVcs/otpwJXS+jZfEAl86x3QVU/S+Wa3P9jxp
5BBYY2bJKlenP83rWxtj6aXNg+ZLVcCY/uJiQsGNzGcMpNX3C7J+fMBQ5S5EU0tn
AD5Diq0kznvNCChtA0o7HG/UALwVEWeLLJhbgR03QKRaJMgjLtAXhNVJopQX1hkM
flJkCMQZuZ4UPy4iEIcKAh5KPbKpQssoFzjbyCyDB7W0Qo8ktj4N6GvLDdsaybnG
zekYhaNqU91qHysziBGh65Rs8csmu6WFZjJMOGC346+TnTFAQHkSYQl2YhdfdAeR
3XOURQquSiTQfU1kBsiRbGO9lNp7d3+J5j1r+7dBaZzeB+I5KYfX3tEkkH3N19Lh
Id+JxKbnwGjxT8xXQpEzo8LSUJ7ex9Nv4mPOIIbU8YoDdA0wdi58Qi/FAj4Y9wDS
/8pkFhzcye0nTvg1qX32rTjb25OG994+sNe41babETE7WEhZyH3yl3BK3HY3LGNX
DvxCwC6XB3TBZfH7kG/4wSihEPHeyv+NNfa9pf7JQaG7Qm8di+jk3+OzWrWBV1+Y
f3MBlfzjLrJ5hnMWnskjGK3IIjoVSvssTq5XvPlBlXZ3siILwKFW6elkqzL6eWdj
pbKnRUePlFcp7+ZcFhrlM+av0KhVYpJEg6Fm2MY2SjYXyjTIeABAZPd/WnTPy5Ke
KV4CYxlPHSSvOyHdKF9PnPk683BVOlfCeTpyzYyfssLnmTln1exIUdoZHgukWTkI
38qMEt2OQwcNxz7VzXJ3ocYLq+lQe0tyq+TewIlYJwJaQWtTKd7Pk+xcWoVvIC82
xmqMEodPcXUfu6VFJSoQpRtJ4aLSaFv4a26W6KMNxo2p1xII0nsPEZwNgE/SwtY3
Y1wJOz9zJnJx9dKrlqv2BJ0H0SC6eyusRmYuBnojn/yWNFST8eXcXvNvtO4IfZG+
Q1Eswx6Ts0s82N/RpOisCX6+KHTsrxZzHv+GWSKIX6jXqKvZ/cJi+YetIYGGwpLy
YkOD73e0adLurlNbyXL0osZBek9qhPkq4cJO8SuuexGVmnSW6JGO/RSAv/ZrcRu3
M+DNmLf9GxlhDacHwN8I15M8ERXGawqjDT/qcLc5IlIB9YKrtESkrbGQnhj6cP4i
glyrxk8Ot3qhW5MIq3yE1Aurq4tPpv0Am+IT2xYe/28l4nSgUOFrp6lMsS3kTE2x
Jj6ZxG5pNd5ZFLuzC0LOcI706ywWy7tmkcC/KMqSV/MTKs7nmAWT9ckCjM07H83j
3g/RePa3vA7ui51xNWxuux0b6KF5IsYlXoCcyB9EohgEDh8KEE9tmBYmmNao55Qp
q6/fup00TpG8bdsda5OGt3M2YVViyqwStCZmkEjPIb4W86eaXM5qtMKrOHZJVQSV
6nETQLlOhEjeblSUc9PpWGPjZxpg/fhx4u8rfm2lJsz4ArqDy5TODUjPmXFgdmUA
P2bx4sODxFXUuhUYBnL9FbU3NhJAfI3QVfMAnIie1+3xJUYK9PAUz3t5F8KSOBoA
2AwDsQtYqiMTvCYcoXZqyxqVrxA6LlOPEToOo9AdYWnW85hjdXQgo5Z2hxtmyjRd
7CY0gA58g882MnloRM5Y34z4+hMg/0N6S2ysUPWGJiD9NJkIJ+V1m+jRsSSJIyFl
zoPbQZlkHMz/S5/nLDFJwJKNNwBNx8xdPSjg6UXGJUWKRWBUI9WJXdtyJWO+P2j1
Lzd9gOhhRgWpQ+Rg+294tcalwexbRCCn4C19VNwSlOLtkb07J/9o+qDkCIWrBR7O
WuYUJ9F09U/1LWH6WqCaABrE0ZqeBuqSPYpyjDMmacs3EjyndH7+A77Tpc/kNb7J
ytJpg7D519RwgctlfoQilLqBRYyO3pvyZmQtqp+OKBd56a2DPfM7XkTHV3Ce+qK+
g/EdaATdZw3YoU/Hkd7bOvndiXzJAaETY5LVf5iNAG7eKEqT89R8iS2jptyp9ogT
CqDP3CAlL8XQVhrrgViBkK7aUrFCLhzYk78oq0jSNliCK7o2bDhtH8HyV8nUUTC/
NLlNm9j2Afike3HpC11aatLdpbtYtf4ScmcQYzCBZblN5pTBuokigDkxx8QrBGK+
9vaig8g/TR3loeJfr1FrssHr0qKYpPy9YIurpGC/pJ0Y4RQFuYrp3IpBIubwS5zU
btJ/tnsWzD2bmmrf23w2hnvEF2bZlOpOxVb3e6VDiIFOOUIMh7R5vfNEPbWLYVXo
S2txTMF3FbgpEDuvC5eGZbC/VkHJbGhXp4tOQqMia8VpJnZx4L9SR6GCU2Eo9QUG
B6ZC2iNwYa1RPBLJ16tZJ9sGIVF33J0z95tqxlu3Ix9DOn/PCR63Rz+VSlvLXSBR
XjXMTpW7rCN/7S7fXMX5whoKX2AWSVVwNqcXxLqJ7xGs7wPEe+ImJF4Ag3MBlwaE
sdMLzIaHThj/kpMjjMoVD5Y/QFYc9BaaF2s7i1vrOozSexvnUtXfXv4jw9FZMEOJ
NkVohLMYi+QAEEIAMJg0IgSLlrwvuqagYgegQgr50XNdHEVkT6IuYiLngoNOhFfo
8fxCF2VUG0+CHSQ4X8umw+89jncSOCFdzHeAYHSFWDDZiv2ala7fcTeGh6QHGf7K
eG2yHkFbQSYIYBnmTFuLlnqeWQ4IdEuyKiW9i1h7ubHSmPDbkgGcORvwAb434YLR
EdfRIyy9UPaNG8h0lEGcs1OxT9jnjPqiVSekY2ntFqN1+r7LytdzhYsZUGXyhqm8
cXctiD39cg4/K0Qf1OTm0NxMyZugrwwiqZSIkFkpBD9ohiS1BZfjsW4eK6ZxT/Il
zwsF4sgxSR2zA43o9zXIIHcJIIfFEz+oigbdpVLlcvrbriY7eIO97KE44p98/y/9
lulpDyQihJhI1lhVEoethNIAS17tpTWlddJ+hpDuKxu6wSdDatqT7ESyFYM8JpE/
PCkX98Pm5/OSwdU3L5Y07NCylow8/ICnvoTej3sOeQTWnZy2DntbMzRHgpgpcsey
0e4COd7/mLUww+/3kD55p9N3cduoROf689nYf2e1AwfbUIkffQ+htRKMexiAc6JX
RyrBa9xKakevC8OWJQsHOxEFirByKweuAJyXl9ta8wEcyapWh1Qsy/IFDV5cnyvk
SzKMbPqRzYpzS3D13Pk+j3A+usSEQ1bguhgnC05JAfFu+T3eGlwwl4YxfpKX5XBK
1pVzDxQBbhUnfW/w3YNyWgetFVgUpHGdTn3d8CNR/WxwR5rb/EwArm0QpSq7fyUa
6Gv0qua/I0y295isVMdrAJXwmq6bVmkLg8uWPVJC2uLY+7EXS64X4E+tvB4P2Sh0
q6lXPz6Y2NkuV/Ofv1z+in+fswWtFd/dBJnPHd+NoI4fpl0/++m23rR7V86BzgLB
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Qco+rCRy4XuDd/vT8UQTsefMfc6+2TNuRCS9KGbprTE2mYsSNSw4Kbozb4nSa5oS
TmgC5CEfCLR00RRf9vKaIPoM/AOnZ9yj7SU1Q58VHAJg/AV93aX9tnZymw/nVytZ
6Wg57ghDGL1QBFq3IhxNbMjztdL+b+tkU/puNJPtwYoYkVsx5cj3MCbxQ9SYtwHo
CRV7goyS2kwPKJfxygDe4A4rd48xsh9R/XM+r62HhNMTXtAi2nseRH31zqlZHKTF
SnJjnS1B6AHPzlmD1QYAS3FuzsuU5btFiCebDMvFb50UG7fZiddrL10IsVZQvY+A
Qi1cfpVF3VPYkGAulSU+cw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2912 )
`pragma protect data_block
kfRDCtNU+u4j4MONvkVS/bM3vCIOzNTD+UeQFY4RoJwAxV7lM9bK7nRtj4EtSGR1
XQagZkwDGPVf4GT7EnZ5PH3Z5g2x1ciNUX7em2YxgImRrxTSTUblMN96oF4aJM1J
yvzqVUyzFZPhkb0YQ9mE0NgUqdSZK1fzZcMjaVqsN0q2FBQyBAYLV3qBSYJptRam
KUpqRzDmebQGUj9oGAlzGS0VXSF8jdZdrhCk2bRs1o1oGb8eY4ZDuvrETZJ4S8v+
+Gp3o80Xgh6ub4n/6pWfx0lpACbHW17sPydfFUZclw1Amg5zErPDQ9Fio2kEz9yU
/ZpmZiDTKbQMjKcCA7f49L/QF+LhMOr7bQqg2zOlQjF3Et3g5nkKW4YbGuiKjEgL
633XsHJS7MqbdKIaLuBkwxwFN+3KVZvG9+S5Oj5c6dq/o7EkhdqzoUv4qBwkTpEB
AJOIO+Nh6l9BXqKflJvoa/YjRiOuM2euBjSwevFIY6pK96ECV1e6Ms1UNpBecBAI
2D/FCn+XrNyz/Qm0QRKqHLsp6Cg9IQS8fZmK4xQmXcOEk1P72U16GpL08HZ4hNXQ
hZFatJxMvYLebRqDMi2R9n2/qo/3S3v42ZSaU1wpbYBH+LodQmnOSll0PlIL04kt
Hb30/JFjqZqw0WtlzFw/LOBza94yuxgry8fWMm4n4nCfTGbixEGPvZlrLo6+IsQT
9ckwDc4qMwg//k8aUZC4w7zDOTESpIIBXUAnNJ1aWMrXoKO1VNQMQ6/vO51+jPKt
LycBsDTuJZnmYA7llARWxuW4159bfRXLfZy9A0gCq736KrP1xOojYKPfTiayAP9B
qikeC4i3g0ZQVtN6/Qpak9ik8sRoERL3Fjw9LbWz32y4RcXtAp+61MOiVoFH8/IQ
sNFSCvlo7Q/veY1WRxpxKnYijvV7JTXqnzWsJEIdxOHc6Cgp11i7HU8LNH737de0
iJutFkVSpKxkYv4Q0VkkToIuAQisGw3m1RDneqRMNPX/mP0OI+NvJna7t6iMmteQ
eoSLrzrIQu9dUaiRC4hVbDR2fIV9TIqR/fL8DrBo8gCYsbXRkjMBnVov788huug8
NWYJZvMywqDvKNyPS6FGOntAF8PKd2APzGk7MlA7idwSzfKBZ0yyza3Y9dflM0Ua
L3QvetWUZO/92zelB3xqPwwfNuAl7bXaB8HuLkLq0079zV4X/uKBfCN9tUR3Qdzq
V02+a7RbFkE9IfcboPn/jUCK6y0d8yvqISat2zGUilLz3TeYqovXKS7s6kWFUk+8
EDO0KPJ8Au/bbErixXRBaxKQaer0TW2EFccDK/OFnolzvAnV5Zq3HMkdjXDRMqXz
8TUuZSZG5T8CfMJmfzV0VAU6Vs5KtCv7hDpJ8NWLGY3l59LsI2u9n2LFfJ5KEU1y
nT94NCAL0wxDYZt5JxMpOxoMXIFln7G6uwnN5DGx/suNOjk1ZI6dgW1IzL7qpvuu
x3h5xfKaVO0qCWugVpmAqlHxujXTXVWXbxYhKQo6QzwslvaBmdOcHTHuLHHLpPAA
z0Qarkv7JZXTEJb0TFp93lMddu3j7LDBGz+zMOiiTxrEjfya8VFDE+fJxdbCDM6a
RHe/C/uQxxL/OkaFYMK2tMIRhLp1ncU4VpXpyQDfnq03GBISJR2cuZ70OZQeLM17
vmh8PAMN5b1C4i1gjt97yEiG9P7tpQCHWoDkm3W+sOzC4YSUr0F5CqhdhQ5FhnSa
CtccYjUuUM8o4g7EWvbKHgSE95RyGJlFO2LwKQj8Q1vK4faR6JXOKXvQUEb3TgrI
r1pNu14S59stZv5Qetjk5iP+f7aPS1QWDTrAbBBHPqA1Iko1KFWfSkx4FUrdwY+7
sKjP0KwtfvfCvdm8Noa7qVJFkJP2bAyUNBHe0UJZj/NA476n5UkGFzHcxxxRiR0o
haMV9YHSgOr7KVdd+9QjHmoHymvPuMaq3khNTy4o7TWtss/bJDYUP6Fxu6GMSEH0
m/k/ZeNhOvIQHKpaRfhML5jqoNrteY93qA3U8WBvjDGgE5+e3Qn32PZP7jYLx2t3
G9oAv5OKFMIdwYNRQw98SaUpwiQvX0S/c0nFZN4yxEnvHYK3nZYjEgKGB08Q5U3w
uFMd5MYHvgiRDs78hwY6ngkT3aWLoQk8eGIqrMmFMDFMHUryP4+QXj3nxOajm8I1
Lt5BrCf2SIO4OgLnIMSUcbYQZSXOoqbbNBNoD8BYXwJ6c+r7WgKklnaDzwVCp2Ax
8LhFrK1676yTBn/QuDgTIurgkh9JHA5araFRugPly1Rg58RHZO2Xf5JxpOxGv3so
PdihBXrhz9vS9+qbTCR6f34pm3lD2YUGMMD5bw/ANlLCJrQD4b2L2R+B+gUDbtgM
IweYySr8DKfZt6tdabMnCUuefSAu0OQLatAkMEgFcZaQqCtGh4J4J5CxEOXHueDw
KGFrB327IkfD2mU8bCj5KevZBTOEIV0l2yuDU+s1T3IYXsQvDIFWXsVRiJP5rovc
ZHn1qpWBTqCnwQ0rF7kAXgX/VdiX4Z36m9wxAKIThcWsJX/dvsAmus12SQUU3xEm
9IAmT6mwaMtdFDATWtYTNrT65C4mo78fb0ti57SO2a1lhPEeok1KII2AHGpLIyGk
IhWGRaX+7CxMBD6g9NhT8qvskFdGgVFQ92peBEfqiMwO6gHZsEsgoWbdKKSFyfTm
QM+DG/AuoPM78hSf08blT3NK25CaARxq2PaV3M1jogmC/Fbfjv3jKi4eqhG6GnJV
BUVmp9Pj2dxrmBTU20lJ8hGTj0FshOrb/VPOTm/aK9hgvEkGo5A3zPjbysfrruGx
HUt7uVx/4Nmc4TnrXcTJ/0B7J1QN/ZinrS7+jYYeYdaxxWjh+gStkxtam6MZRMNi
P7OsD+zMOtqHHJ96jlkgxsqrSn0/QOc6J+5SdP1UpcmOzvLg5Mn47xYoyCSrMNUD
hCQiv5kq2ylF7JDcLmIqUBbrH5dGm9RPqUoX0GcEqovgehyXrValXJ6LzU8ppCjI
hoSZuS7f49yAsJjSVLO1Cphg83ZuPBJmcGNcEZhqPLVVne96uQEufp9Ycn1oiMV6
0kpQ9t8pyKSQLpa3pYtk7WKCQ4TkPtBVgd1oWCRHS4/QHjDMpNJuMMyXX1z8/oD/
CrsGFSOXPt7AbT/ziULs24m7VUQGYCTN9CbKYz653fHogDoeVzkPGNj4A5eRN8fI
kFLS+v01rwSqmmLXZUVv0ri+py8KcKy9uuD0IrZtpRNAnvmgc4ZJbp9dsfOsfK1K
4glRHZKlc0pXppbA/1n56RQ8kz1DzToqTlWX/5G/wljpdOEDgz75rBCsxsX+6nju
ByhoV9N/L2pUHQGmXkx9Ey7Vk5YKkzNIBfszbib5FwFNlwhadLnmFUm/KpzNARmd
aud7B8TUnSsfjuRqM3HnS5QHSwpVMbXnsj9P9BdB/JGTKzgI/tkQjFJ/i8SNahyu
TPBXR/58Fm8D51Pv88xQjm+SCuJ3aTwnHrjZFeMuhLJTuIKbem68e5pSKEEhKMdz
+MeWKHwtVhesqr7eh6aIlXbVcGIm1bvOxY1qSka4OCBra0XpMwNjaMFQrn2LRvI9
aCRj1PIti2K4aIuvHnLTLjH/l0PJN1n+pG6lJ0AixqCqnRlWlyHcKCPt9dA3hwRJ
agSeI+wHowTgMCvfFR9QqXRBPi/7KNz05D9FcyVLWbVAoojlkElX/hDbjkPFVdC1
7kdxSWRaOLTOqtxG6U2zluUL2ItEgGNZs6LQpuVU3NdKsilBLhOIOTyh6sPtKvEt
Di0nK25E5h1TqHM54dzMyNOT2ELHvdTF+dmGDtTph0GeKGPMjfZHvMKwqtbNKyH6
DfG/EICLH9MDHQbcQYyHZ/dYZyu/TLTJM9gKdRvkV7I=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
KM8sZLzbvb3AZ40XCy8glvkoVRqx/FCdKA08cPcbEMHTksWNqtZm6FU3cEiiU9rH
ttxCDSnTQB/D2WvW/apI8DlBMaR8o6JUO2jQKCki4p+U6zYdY5mwYoaF25rRQbP4
ujUPrrMyek+QqwE6BDzKmQ6nWWVRZip306i3zM1SHD7dqlaYB6M6bnLCgOncPcU4
SUm0moLQgXwzVAxSJOCtO6RCKLH0SCfK73asFrfwt+FI4BVrcVAkLnFzmsTMwYr4
YqoKQ7Jslf49mYqg6fRn2G3Ov1uWawdeYsVUUCgnsa3GnClf5lGGJqgvoTcKbBRh
rf6ZjSxrKWmbV6CZpownrA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8016 )
`pragma protect data_block
eBacXWmKQZVe2GcWI+Tkdi4emHWzE7dReuLuxbwZHiiTQ07QCM/XY8elsoNkAMm3
WAsdnl7VvE47cEOezMaR7WGhaF3RSKfda7QH9N24yZ/i2ILbzCW8EClewCNs3pMA
tB5z/r9hH8wYb/c3rtcCKhZ3T1zt0qJXmAe7rk7fxoupYPgqsICHQpYifJuS/6VZ
KW3DvE/4qmSkAzcHNdQqn8GCIKvJHs7vnnPcv7wrSkgNJyHvimsh0RNRQQlPqFP+
bnDVo/TkrsdNPuRzL4lkYo9uCr/StEea1+X3XPGf6Kez9heNCZ2nTijRBy0TOiqI
X73q/qpaTXuBrpjQzRC0OY/AYg2S8F1PveyV9IKw4m/Ram/1mtfs0pM5fft1HC6/
oc606TmxbKaaNKA1QIv2r881yyk1gdqNR7I2pnP+GMUamX0Iixcrz3PzWM+WKlLe
0OTSnSGGcOCRZW3KNJgVZC7QDkOZbMXSNYtNjSr4ON/PH4MW00ZJa5XvrbYocGJA
/D1sl2rEyY/e/MzFShkYJQg6DaLdxkYLmrshmrHewt7oejC2NOkjEjIkDG8tR4qP
hCYE2I/Bqw8SIA7GJniKurhN+QvJtov4gXKZvUIInKjUM1Cdd46CAdByqeoq/iOz
gNVzex0ccfcTUnb9hBU2RkOyGTpUbSthrG2HX694bqONAtqt9TKytbuuDFIEK7SV
YIwqtIB8LBTmqjj82SbgiAUz8pifjYD/MmKXLQN0qmh+7gGUVGfR0Fg78oSIJLgl
EBpObjuX5Bedsqt1FZ75bozcBfNeeXG+mWHjlNl+LfEthur03fvpmjIojZyeqU92
WygP1nXJtIv2kkLabfAHMTWJrq4thPwrrJG4pHdb3X4zTZH6zYiuzf2RpZI57fOU
50mIKa0pkiBaP2LcJsKG9gNqGXKn42F4niqbAZPUMaUWbcUWb7KqrBRO5waeiy2h
FQLiUe1rz4RFct1qtlLx0ydKHlDjQg8rZmFYWEz9BCIeA8MeeLMbpd1hkfXR+dv+
qHlmug2HiOQSkgZYOwvAqYpq3RESvOAYaaOkj+sGuQIckd6BD6ON2/jO8cWP/AVk
KZiLdUN3nrXS/VoNI421JNoEmrdk4JZ4wW4pg8KJapuusXwKDL32IKTsgeu7smYi
PIdpwfAX9ntgdB1NFJ21jF3qn1uMZ/WD1nKlQvnk8V/zLpzAPMgF8UAcVXos1i3K
zOIHU0I3VPv5dxOHMILletyrxjxAIGqH9xyoZzKGJa3/9YvenFVXKO5REWKt4+QR
QI2Xsma/BKNrjSwD9C0+GOxvPudCWJExCKWR+iSFoEqsShXTAXfh1+kf4Dg38Vtk
T3YVU35kKu+NXZbBcvXk2zSb6QuyLkVrmMuNtxauoFwXdkBOlgq0KUOzLFBpsOWB
TCt6BWz0kDZ0NdyTnj/TR6MsJTr0ed3utEdLZkKdubg9X21zEYUi2mY6WcjkVW4P
wHMTgJ2czJhix9yF6VgSOQnrPO/qQBg/9ua6PBWSVh9vopL62PT4QHgdscZGeLDL
3dyQD0/Et6hdcYg+7hoYAMwpFEArgM4m91BUeqxay4xQGr5tVgtW/QVMAbbb2IAq
pPdOzi9u4TyXP0wlDu8+o3qsEGJyBVdnFhZ6eY+rRStwEXVJrMeHnKBaa/VAGKwS
l+dmMRni+7nWoSU6PZVOLtaGvfHBbRrYSDEBlJmh65J1llROjzcCA+1uciztr7c+
jzDP+/ubXxVh4HCM5lw4j2n0ydfx2VqcvU1c3ntI/ZICyx8hWF7+LePJHK//EJHd
w1J0Xj1nAhsQlb178cyo13e4V9BOluVvFjxNNli/+D6hBhpGm5GdRzAUbQrPyZD8
7ZiYOlbdlYYVXGI35hmN+jpeCrcS1JLwk0mpdiJQZ0HU0T84TP/18Z5nRwi/WI6F
RfT9Mv+UeGFSOKLcXabirPBuJxG0GYGzSK+ex897ZyDFTxH9MJQhNLxWhk9Uwiqz
anXwrm5tfs20f13QY0fYQQ8kUBoL7Y92UU2pLRRTqN878WHXOh/75pFIbXi01ERW
aTY7aPcMwEz52OzQMbz3tKCd3AXV2/wIG6ncw70uLiYYv/VVhtqAXWytEQsRfquv
Rw5fjy6usX1RvhQO2G+u0h49eVZOF3yWni5HkBZGjJRFPEjevbBkSY420y4+1Nvs
SWSLbTkJ/AOgv83ARuWwK8fbKdJAS8wcxHvlKIVODqypNtZ8ufIJY1LUKjzc0CbD
MgxXI7lmxhlX75qGELEyk6cEd6DjSZrzzpwOlrRc9ZspKUpCskS3Cwj2i1QdAI2p
nMnWCayTQ9vD/RNfO6tzbGQ+wQDW1mEGDI1DSYoFNv+X9excLD7gYoeAluBEj/Sv
vdx1hZD7jxWVCSZ3+fzN25nqifqX5DkgCAFKgbNNiSOHz6RGZR7MgORShzElwz9P
RJ4zPBjzK9hEizvVaI6hAV7uLDcjLMebBd5BCDXFfcgwNNC/gCDDlpLFjGCWVYtI
bQRsOqzq817uyR15smcmLHcrSK/Lokj1mUWgXFuR1KDZh3rDWkBKlqdDKCFnUUzd
ZIlzT2Ryya2Z4Jt3/rDGVMR1kbMMAUGSV6aIqpv2Vx8df0XhuoaCzR+MosE8MR8x
oK17PYCkEiQvSOJIBDOiCTgr4PsIXZPx3ZNNh39CJh19fYp/G+rkIPoot7vibAo3
0Qw1gBRlutNy5axcDLnwELMUcPCVerSZFzflberu/MjaJSOyn/qyXdYt36yQIwq5
3sOOgEVgcsT/yxD7+/h6KMhopntLXe8x80AGW1XBdIcpFMnVc3eQTqQHpsH3AUyO
k5/TJEsmmjSolsOMWPVwTH3WDrMcaWZH4seWuUCuQg0hdWO0ueYZMC9eisNgc+17
80gjJ4EUwr7fGaPwyWBiRd1ZoP+QFW5Nj9c5yr4Ti2tMUmpcSDwvcA9DKWKe1vAy
fhegpKue5zr+o2DiiDTvxDFQC+lGeEjRUHFLaenrDCTKJ+RKkUc/w5cdn4ZXpOIa
Z6kfjtMh+gfPYxi4LBEYGw0CImmlF/0a03ZxyI1DfkVFrcgnq99+E6bK0VWhrnZu
7E1bz06HsaWhUFi8OnreYFc937lIFGmn1EIbhL79gc3xcs84bYX3aI4FxLTXt71j
9fo3JvnFIqrvKTd0L4DzZcJc9sBwC3ldbLesJ1omUbKOwueZo2bUWs6GVYInryg9
kg3TeQiO6OfwJRTT8xEu9eCPIsTb/vZE9WhmoTDe299INWVhUfOuyYKYfRSX2KX/
+iURbuj2c9YZm9lRVFcwRFoFH1CCpQr3f1wHgwhMT3YrV8aOlUlsHcUXquxdSQ4W
kN3eJHBGbfF2WU+mqb4YpHmQ1hMzvDAJfjQbhzi1lFaUeXiBWGrnu2ZJg/h7naFt
V5AMNzH0xePR2U2oTLc9X5kLJOPsa9KaIk8f6TGsWYA6uWZL/A3ZJ7GOFwVrkvpB
+LLvLgWW7EUvCzjlDE7O7b+DLAQBoq0358bJn6kgv008RMre9MKggUF5ZklfvV8P
peomaJUBgcwWrURMfHLq01657ADf27fw1AM9gB0U73r5uWEvjGiBQ1wdlGFJMM6I
b/rBAfixgKylW1bgIAwP9QDukNHFqgxTdVLkT4eTvSl7vN3gsXQBTPCHRt9a6wpI
q/pPC8MgESk8M19fvVesPBFhLHPd1BOPBdJtzSfmU3qT1yNwGoToYuNFRkgMgBwL
D3bfV1RK4G07PXgRll6NQX9bSKlC0ZTMesZodeuC5/4Z6rVh66XGzfjDa263tw3/
JVYwnUlg7OI1gaU8gyjouRhd9zmDOiwgbSO/y9Dcpt0ahLogkybj8p6OzHSTTezR
rUlYhepObBNvidpc+DmGlGcz1B3vMrpl5A9Ttw9C/KuMGx2ZOQhA64zM/QhtNijC
iaFPPxqOKHCBE8q4getQGdFWT5C72jTHQidTmwokZwzMSuU+taGu5qYzOFXF+0Tb
V54F4mitCW+xDm0KMSs5S7cDsZwc+hSftw9RSsj/KiHqgXGr9aqO5qbMUwe47WoQ
8xHNuHWZYbfXErnj/wHSu3d6z2isGSHOrRHu34c5rxJEjKu0WfqPxQz5bPWVO+H6
jp4KjbqhXMSTiZ6Q8sbsjGzOgNyw/DYMglUZDmWhFSllgGF/dtQOL5xSeymVeH8/
qYF8gSz/wBQatT15Y0rVfGd1pA2G6IxCpzqZbNi2DfcyWJBB1sm/ga/2DplITA0T
N+CmH0xLnNu2isPARsorLtjIKetr+Wd9KQN9S1YzGFBEWdKQwbTd+J8Bpwt102NX
tb6AfWhOM9WvUMYT4drKGDI0L5bqmdKHyclMCdvlF7vOdpYOf8hBn9nAfEZ1r+XR
DGywp34lqiKQBlBkWe9Mo57FS+on85E/5eOXcPvp5kkMV6SkEZgt2sho8yMbpb15
dpqqrA9aAsX9puS/OCpx/h0ACs5VR4xaL4Yp9Jv6RCp5io9aicAsLVLpWqYYPYqs
VbfLW0QBRVOiLVP8YJFeVi9WnhtMjzPMFTqVCug3uVG926MX4cQxzPxiaR+mpaqV
R9qnX/TnSF21AmeRpdI4WSnLlmt7chKv9HiIx9O8g04OPDaXwqvjl0J/HtIMuDr8
CNrW9ECLKozEvOQwvI+gXIBY6KthuUQF+P/4P0EF9prijVM1krleJhCKxrERaR0z
cDGb6QU5gaWu3jzXCKOhMAlTxV1U8rOtZUNe41DFl2loc7Pc5KUAehs5xrwpSCqL
dtl2VPTkf/q5sNg4LJZI7yrzBD3I28nKufBwRMaplApoF5cMqbxF1N6jOvoz4nUA
zADTYuaiuIFe2bh4ogW3g3NGb4AfCvFs9y9P6OmWOPgSjlwxkdKtj/xPFMbBhHGg
h1FEk8QfSYShB3nj15gxhqikoPBIsdUqBSWdoTKeF6XhkVfmgCEqbgSDZ9lz+34d
mEQm8EhyDkVI95zBUTqdW5KFW2TQQ5wRQggICtKfYx4WnS5S/zf6rX7OG8zJJSlQ
VZ9MMfkwW6bxa8dhqjl3P1YifNb6RsiLJQZRMZ64R2bxAIWYkra4DvCHHUb6yOwZ
rcF4SqB3U/yTVNR8TubTf2j0EUITyVrN+eJ/SWQIquM/2VuBY/6XbCjJ9ozxoG0n
WK1rM2RWo7SmVHvQ7UfhmDKzsmh9b83piFA1GovwvKuOeLOWPLMq5tTho3cGDAyK
3gfot8qHDPHHhOEbFpDlbAzJ2pkZAwnxRkvUzhIihE29UmxgnGm7mvy+OcuBPZ2d
o+nge5lkNHuxCtJzjCXfTCpTZQG4BlCUh6OcFRuvIQKeIdmGAVMlwhzDi4DLfBJJ
4Rwrf903NzcAacuHZm9pPVbXyPp85RElnVsoEjTU8RpuP1jM+XKDeoB/2c5MJgwV
zlTzC/t3nVKLukuZpMyhZdCBNGZzc1ASIhk2F/A9po5c37e7eMsrhstJWY1zMEIm
2zfyoAK3yvM65SMKqbcJuRTVGge4ihtbyy0GLOjDCx8FtISVM03y8ZLFG+anjtvS
neClaw1Ck0pUwffLGGUowTbmyX7kuHV3Qpr3gT+2OjHYGT2ci6pCxFFxGicp/WyC
4uwoFPe4/ryXrtfzHyKqFcqNBOB+1yR7YhX+Uzmk1hlKrNjbSq0ZvIhUWFNdCa/H
7rTCrGQuGWuGSaWTZZsFtF/zQJ491AlHvUcgQHBh+JsBcRaOmp/Ct739mh/rnKgT
GVK1aTpH+m2xfrTmQot6bMB73Rq/ay9WKWDq7K9RkwfBzXRs8VMOrqKEDDQ8ozK4
4VNRlu3TVHUdR7odEaGuJjl4yAmq4fv0aOoDee24a7PYJFfEm4Z7YzDfA6J1FWGm
i9q1jyRFmaCXN4q1V6Lk1vOP6hy10/NqoRaGJJB1bFc/WQZ1B5rbTApT99N5z09B
88ZtIe82Is9J6F/CyiYjUkF30g1rnF7ViuRRZ6lPQo65gINBfTcta/9zoA3/RtaT
ppyZA+DSxX3mUBLIbPl84VHReoSgaWJaht9+UEb8CITAi4KfC6LV66J3FDHDn+ze
RBerkVBMc1ymvNH0nPNGuCojsq5ksuPrQIrXLikTWsmRsAsnTlP4ik7Uu6Fccn4y
fkMpS5k9kRl8gWLvvyv/6RIgA3K21P4MaG6ww+TKFhNKHmgapIrn7EU0apcCNToZ
0mE1Je4Qk5cIqlhniaaiQ5+uuGX3deoB3tafgOfFkYvCstTM/wdGwjhHxKE0VpJd
AcA2YQx0rO4cQaOXs21DH1G5R9o0gOOhwrTkqnkXfLFjMZiBjZ/wQZVngNuIYKab
uEgeu0wRdGBSaZ1UEfMhGVdm2uzEGoFOGwwlh5QbgTmgBxCMXHaQTEFH4cxpw4FR
AkwPZ7xxyYKgoD1oXf8J4J+J38cxrxSzicE2nAnmk9/+vcSZA9CADfQWORXwwj84
a8pETIsJtQp9OW+lQc+mYDhutCEhTeJkFdyBPY7fq4iMlODstb1eO0vTiG+Au8gk
q+aUom+hFn7X39t7CumptQpv+jEiaC9QYqaXUvUtZAeY52llRDXx+aLj6ojeYhhO
CDZmoRw39HZob+v/Ja71+9c2jcsypg+4hZQc4NNpPMcRUs/UfKpVfnc5bh2Ae5H3
Pc/zgxa5H47NzQGjc+NS/uwmIvTlT+qXaD91HB7QdooPCNd+nXE/FQUkR8oevWqX
dbifUKZ+lOWFE1Jaj7yexnYVgTQeJieUymYzYVFCQQeCZ+qdc7PUK9AHy95ukaA8
2kUwTeeN/TYrzXhBD3fWJ3QLqOIJDcmBQ5L4LtF0OcMGInoVu9CmU3HVshfWizsH
7gaGbE+iVmHKTDPzY51xpC/YHIj9fozQ+Wy4KCg5v6u8gUydWmInok+GxdE9Z1Ly
vOH+GmT7Xj4N8o0+IIzcmvTaWUN1Ky5tZkpGKVRHyvmjp6zzzQy826N9tEmjX7MU
G8/WvoYgCY+aU4+VBa3rWoXPjqPF6m4WnTM1sYS0YsuBtpkSwsuhSVWVjzCJAAfG
YsmWBIRVjhCAXo1fzRjbW8TLOY/NSUMZu4kq99PMXl/+XsPjdFwDLAQr0RqNm0w6
Jbg088ipN2gEfgISLfeH1eIoQKClMi2DM4DnQLx8mk7IT03qEmKVoEsavTdbCV/0
EPwOtW3mPBwodKIixGp11dzvu4hL1bgyQjqZOYmopUFKGZ/QRSpgDU9rFK70vwHf
3JzMm94HX4tBwRtuDuHhPp0tTIhM9bnDEy4cQFK1i2LOKlP9CesqDMJiKX/8W/2Y
dNiZifpHQSwsrfNecGKL/xYrKlL3SlVlVAHdBK53AOb0TgMPKAUMXqbdFTmjlaVK
u/kF2iqA4Bk/2KDLPAkmtBS3Q9I7pSUGai2OZcbVRZ1dAE6MMQJSpaP7WyJmxrbI
mWqaJ9280oeEmeA4jbHGXhQqz0HVjmEQnE8sYmHhf88I0124VS/4Vlm66NHBFkHi
KkZin1swvPqZfLxEo1nz9ntfvQ0qbEaFbGrgDeERBttwgSnXXC3FM1ECh0WM0yL7
yqOx3Ww0jrKFBx4vvG7WJcFZu5LBjxmqtDGjih55xXYxBKThrmKodAqymIBRDdoa
BWvv/tjRvAv/YU9dz8cyV8gUZ7D0R2U82cyaLCzC+M6984V1wW4yhaGWo2H0AF6c
/9G+bzSsVKigWlAq8HeXiDR1nC+ugyavcIU2p6hE34GdNUCl3ZJJPy7eD9WP4N7l
khzQpX1YGqJRdOxvdWQOpyiHM8GdswCLtx8bdwA3QPbHwtfHYLm8q5dfmkv9rJkT
0CrSJHOWSrJjhMYGMJBDVquf6EJ2mgVFrSpdQFxJuwz8yIqSeWv7Pw3FV1h9IAR5
oDYiytqb8LfjE41y1fH+iMWpnjil8t1PsWqY4uyQA0osSolv2QwoLcTBAtvcPhvw
zi2lJ524IoaYccGRPrUK4ZyQo59Zib2ypzjbTmZVvwO6krqUvEuEUu7k9c7LfsPm
i9g/UbFS6ppqs3ejIdKc8FAcp39hDNIwCPHLjap8olMai+I8w+zNdQyzEO3gZWh2
GidkWuyA1RQu39Ldt9WEuC/9007wMDKQRAaaMSsEUCAY9GrWAK0rVedpjeNS4Mhk
XBK+1w5R3Zv97IYOPS8FjcpD6A+a6AUVHR4FxWs9X2+9jd+RSRHBBJZ+joZ/sukb
ZEcYBZQbkratjk0ldXXrkX9Kv5oeDDuGIQo0JeOEJJfMvvevQXBUWPiz0Yp04RQx
YMlKw1EL0aoGWXqNsZwSLfY6clFvndWgSY0PvCJGw8cm1i6WyKtA+HkSgkU6uCSm
ltakZKnj3XLNfSF/fwewgW1Px0ZUuDX1oLBpdtPGZVFNcaKOXfpHqmlVkS6oOK1r
6t93xqsho34O177dSMvXEcAveD23qkwAycJW3wQW2PtcH3C+K8Fz16aUk4BBAomh
rzv+XDuYRyKMX/P6jnRBBWLJhVTVyHZtTdQBoHKwj+H2KzEWNHkYhu7LrKzUQrg4
VAhFtwvMiVRHpRqvEHmPgBxbzOz7YA9dzbSfY8/R78pddDhGNj2OQd9kfNRWrXhF
hq4Z5Vn7TuGU3v1E27Z/QiizcwRuu3iCZZsiOkdxsYpa0fUwU0/YEq9FTa/WghVj
u0HNagtRDtW3KoLnnaKQIJGLyoPyiNOwy0pndbGbY3AmKC18CpN8lk9GVB03ueJ+
2LQG/abLYS+cxz9zB56ANXRl1Bxd1HZN70YN/7rWn3IhVVrUNz/Rt3bZUpowum/z
VYJxXwUMfN1P7q2oQOu0f1/ayNKCjKzg1ruDq2Y0tfOj1iMtIUXpkvRPuZD+BgDL
oXFjwN3vYV7ugYmktj2flRqFpVYKaiF8L6Ml6Sh1rL0AqOHeRcfTMdq3Vbl/3/Jx
otzmqk3aG2hX18xgupem/cPlwFCGgmrPF94o3ZRO1AAkMctmDX7Atzmhj8x7mrtX
SuvzBtXCU1nIS1AUaJ8K4MU+YwIZb/ttKjL3pgATvLzJYWHQEEVUVg+43AgWBiv0
kKeNTU8ET8n09cahhAZ14snRW0wyc954hwtmf/caV8at9VAudijSdXiljjIbc4Su
AsgPc39x5bsTkPRn9qvCaw+T+tbui1/7bNaaHhyP4qK/0d5fZuj/M16/af/qSuYs
t1CesWMaQJmv/C2bge7P/a4DRWUrzcetnciPIOoFWMK5fXvPe8fcZwMTVb8UPIYh
iaQcKXMc9h9SyMeFtlGCwYLzloxsCvu+5br+CEtMrVeAeZO7M4Jo8S8QX8DWLoUC
OygmD9oM1E12LGGBQ5oQ8MuBHhT2XB2SskgVUVLi8vkGjyxgCJWBbOLZAGm7irK0
LsxHF1ZtMPMhhRN4x6OHIS7vzkswnahYx7vX5/8sr/HJictU5s9jQBzIOt21SbQy
R40w6wZjVUelJrOZc13o0KFC00+helZ4V+uaRuYkb1/bMteWMDlTV/fT8QnNPrXO
Nr5e4e+gGmOdOuPoCNtveyL+VWo4ncH1isSNLxpgBgzdfhVl5WKKkduIzEIRHF9H
ijLm1PVCaQzWxdiw6PpIPOSwjmuC+T5I49nU6NsrhB9aS480BDK+L19HUmedhhBz
T3XPcd0X5dKddT0CI0tRrwYmN8DDJgYeLs2GpRRdS2pnOUc61j1MIwsh+8bnSIX/
VKZmazecB2Lh46ZMjsMWidOwhESp7yYabtoCfrvNbPGHj4TRBrbIsUSyB8GyC17V
5GMfWaiecRd8iBm1e1JJ4Cc7J0MUNY/sQrRcNaQgCUOehj9HkWQindc7DyfieS2w
7uRSxp/Tg0YT0Ok4Em2kFsqlx7jR9g69YPujYshu3HjB3x+x6kM1qrVJs/cw5k1e
+yRPsZSqF2whwF+rF+5/2oCkhzG/Ia2D6UwveVkPj2UafOzuf7f1MKI8rrFvxhsJ
iMUVERfJp2nZOBdkw77jG9bka3VPdQqEAhkx1Dljb2wzMzYqcIj41aEu8RPNRRl+
cLCrzLcvdrqbFq+VJMg/lmz4FkW5XaeCE6rlqIZXfnUOel5tMDPjcqFkrJv195dW
GhKUJoFRLUupzc4tZJm+cw3jaoNnb2SfunJ/Qd/qGEVe1KeFrzBdCkU6lGO1Y39E
GyeZLdnICZjTAirhUKMzGjSBjlVKFIM1NN4+X5zK0ylmZYiDcxNFnMJj4Q1SCZfH
9jSLDEFJpa91As8iX/M0eA2i/2A0TynlR9w4gxGp5IhI2k1X04Lq7mnJR5rb/9Ug
QFo3GXEwp1ZmPzNN44N0jT8zAlh+4d6z1BkHIp/BvzlJCXLjLfuXFhSLmil+Yo86
NHeeOfDVPT3XYRAsu0Pgv68O6s+d0Pp93ezIij/DwZ1oIJQC2AcGyvWunEmaRAM9
MkGT9+n+VWgS00q5AV9MXl2gA4K8tFuq7Wvoe/WCX+pNOvbDDzheO0l7yDG6oFDF
EHog4nUyegPcDMOXf4vyT9CPrYAS/Rf+gdkGW40cjhFsD0K/cOdBzr3dGXMN+W/S
UPyLAZGE2DuQuOULA+eG+5txZYI7smdvDlR6UKDZc/S3oOogpZdmGOV0R7kMhTIa
18byHO6kQgO+Wozdz2sIlBnGTLFFgQmeU8tD1/G7mur4gD0x7t7KbmWsraj/DzY5
AK3Jj5B1K27hwGENTnhwXbVQiY2MzSfPBiXjr+2/FsXgNEE2zntSjgqLOfCDaYLP
OeV60at50xQTk5jgxwuE2C+O7ZX5F8Q628ETxZhgSucHAhQfz7I0kaY+1lfO0MYy
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ZDd4Mr0WyVPH2b4uY8CZfYefzAmVv5iJFALZiVOCVhUZqK5q6ZJrfVi+zftR5xgx
PHW1BeZtOE0V1dgyUYLaYosQIApcHzebq782gHPF07HLH+OHIDTJLhlTdmcVhtyN
0Ey5d9TDVUcKRnK6Uh8p396L4hP+oLZ7jdGR1Cn7a5GK0qiKltc+hXQnqq13lmuh
8oeZ0dTU4wuufEUelZsXF3NoTwtvKonqX6HclfT7E9p+p0SYwpGygkaOVgW2TNGp
tKvpooxwb3YYcTSp98Jq43qBrR8EL7hvB8o5yec2klothdenKiQZPxX9GytK00d3
O2bSNQXZ103GHmKA7kZgUg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5392 )
`pragma protect data_block
K0EnuVXd70vzcmWXamaZWOThr1s7EG9OJL4zIdKqAmv7LB6QNKE4/NuXpIPAr2kM
4hNa1M+bT7UjHGDGAZCXz8bak8btuR1B/NyfZGkHv9yrmI4re/tRDDoX6Qn8gYlN
mp/51wa5ssdrLXtn30cbBfCadH2FuUQUOgkyiO8I+BkbiOzISH09EOkqIT2KpSJk
SNPRlHzSazryBbOzLZmTabwC3bKRVW8/TkRR9Ch3RGU15RMOAbS7Ynq4NEgRq9KX
jYgF67UC/AH4elaZ6joz8RtV5Mk5SuMoOojQMEWaH4aQleOpep30ftH/EXP14Z74
dQt5WorzEe37XkhYgQfFvhiI+FE3duy0MMHFv6mNqVcyfRr51hQ45Xq6jujVJssd
Agn4V81a7HRdhJaMzydqAYJVWol9Kln9lDm405JmDIJTniHPGL/FMJ23jLp6eEw8
BP/ebHS1Cp+6ZcL6w2SmwvTdTgsuFtapZjS8pIvUhaDzpQulpkj7M3ZyP1jNKxpC
0eJ/7YNy2fStGC+0nA+L9n/q2Si6J/rtCL4D78dqWuvd7hcB5NqycMuWBFgZaonW
/34koxhfGhhv1HXwIIsJIeXdHv9ZZ4KOSR3G++jGHKVoIfhYms+skIljcTjSSyhP
TzAEDtcVUYVGuegVZkPKexgvTJJb83+wm4hP2ZJONuUPH9YrOToMJhu9T4l7Xuso
UJNlcrem3HW5paz85yWzDs5PF2obvh5C3iO3ErFM4YCdX23qBGMYqEqliLpUwizg
zgmQ2LNveRPpmAT4YA73oWNBz4P2rCYWTA6hCbFFCeRraHR4a+zNMLwmX/pJ30Jm
UhcpKZ2dHJ5M0RUeqXwCvuHMMgjxXLqxep/4yEHfKCbcmspsLhQPoe9XfXCMgAyN
h8G//QIO/gIY85dHlmnOrJRsS2ZOwaMHpICGC4lF3AU6MlYxq1NeD7CjTnhiJsvX
HSJwm+IQWjwA7k42KDjaE/O24McrCU+Q8k7QtE1ZlLdTdq2fXKVPSC3eq8dmpmt7
tvradFQnE7wgGpyp7yARyx6n5dmQhXilwiAzlb0uw22htxFZHA/JEiyY+kKuBgUN
0MtDzgr+boBXF5Fjj1YmExfALkK+yFlACYRFj2p3Y8611a1q/Gpb4Wp4AkNMjmm6
wig9FrJRTmavx3Tg8n2npFH2eqYE3ju+5orqVcHbzhG+6r1UKSpYOaah2ncX5o/a
C+/9gPJyV7gPtNPPw4wimhdwPDGMMDj/kf+gIezuCT5DROCo62hUtLgI41yp7G5Y
r1+eoh6q3zjK3W7vYZcKrAxquM67zc0bCb06MEpWev1WB2mq4OKe2Z3YsJsrb3VW
VPXr+o+luFRloWOAMr1brhzCUM9poVZuIRA4Mi8U4XWj8gv+0XajtkNwrmmLP6dX
jCz9kPUkp7E+NjABG2DcDupDibf/B4cAacO6Fm+QzZzNn69AiKS7zurDucRJnxnB
52duME2K7cJi5KcXSvsRXMd7Mzwwy0ojBf/tH3SA31eiQU8zBT5gWjiW7IpA8+tO
HEMxfk8UxhjKFSGI+u4OUhOBDWGkhBEstetznm3Ov38vQnBoQdkiQMKZ8GIDgD/d
PdiPmkF2GQXGPlclvcmQ5/3zjP/PYUzSC+e3m2Vbipe/FDl9ZMn7hoI8OFw4c0iV
S68RwN6jlpCsS4TrHbqb7wHQcN00kZAooSuoeRt6XofPtjeuVCvvq2eacvDC/WUS
iCmXBtI+JcFuTc+fYPMIjWIobMvT0shIcFBbAjLMlySKrekSeho1yQqOlwO87mnO
5l2z05iOircgCq6xbm8zvccqLc63fS9abYLhSb4VTi2KyzkQ7XWx8/b/ZNx3lmRv
YrfUvXOOTvLqFOvQif88KVbd/GqxDXPuqRKoz6SQEAuUAfNRDbd1pNnrVjsjYGCu
1X32y3oPrLBQJhyeYDe7hA0R2dJh0LfHe+IX6EJ5FWJx8xf6NBWuCkBJ2xTk+f2s
PrM8z6KHZgLPoGdh3y2p2rqT8YGBGS1rMsq1XTBNrLH21/tKkHoZkGBtGoCtD24C
O3aXZYR5qwNw6Wa6xtNR1iygB5cXFQRTxrF4maPZWHGIA7CtKZxmcysTg7zxEdv6
lT64XycmlX1eRyc30UkFozyr0sKRUDxyDdyTlVLVhVKC7TFRmWfcbZ5EjYOQR3LZ
etD0xN2pfECrnoCX0AnhUFLI0zDnamnQ79HI6sLOwjGNNDuZAYh6pCBEzIBgo32M
URBAF3euIlZDdJznYgpowoL/sXAobKeylrryulLVB6rlu3VQ5D3iGMrOYJsRDqN0
7fH7cmR0qRouKc8aVqjAmzDU6xV0dYDXUnlwtQm9zUxIGR9b7a6kDwPaeGINnd7c
VlpbbiiyyZD50He/Iur+eMwgn1T+FqLktUiJt9+ejtVs9uWDvb2hna1OUPhnFvO3
I+QA9UADx3WanafgzD9Fnto5/qRCW50DVStWdZLu99f3PfQ7ccR03vRgvhgwQqLB
DOywdNKDfHl+dDnBAcSdjxtnGGdz8OBeJ9Yddeuq81Zi0JOrbbOtjdrdod0DqjPs
BfyJkDpsmAksX3/LKj4FBNeay8J82QQQSiPxZLDHrYx40VJPIIiXbdpd4hVR5Rf6
KAFKka9Wmg+GHBX1IaVKh2FeOn5SFAAQg9jt+JTfHlmRhlhZoeiUrnsHpAX+gAzH
jng9OirB7DVzj83ZZqhodPuKTxbqHi5hDXk9yoctkG88515/ZLNWRYjsa56Cw13i
rcxh15NEMLf9l/YgvD/RTf22q+69pgtjvfABeYovRSkFB8+xWYcqTvA9+PVJy7q1
iaZphR/eVl3pH6IbI3fTRAwfyc78AduVSVBjA1xb59vSViZE6gETNGB0lqBd/UdV
FPK5c+ezP4+7B7FGhYTc9C+ooqnMlXWNg762tQLU2cnd9zyvGtVBXuwC4swFYzdB
BOQzkGw5xI/UlKjScTJMTysDmMj/lNWPZuunUoEL8tqIWLeN6HvkCt4l2c2RtMqa
r4kD2Syo5fSofFqCkRwYYr5LoWiTrgWBPG4Bhpx3U+fU/+lY/p76B8VH1Jfkadue
lezaxG0s+0YVSYssctCCUYHN7r0byi12RQy35to9UePRUGohn1qcPUmfzV3vdNad
TJlTfWkaFUF3TibBbZR+JDgq0N/wCO2ryKGZfIMzku7eadflaY99sCROvSy4UsKp
wTuWEsDOWnOcgo3dVd1+GY6zBjKth7rVd3whgGxriswYRRXi0JbYw6JhwzJEUFyg
SgDLcOqPkC4Vd/HoffD+IUCZhMNw0tpoYnW0o5+1p2O1US9XMGAiYo3DoIN+YoVe
2thgck0Ozaa5B1mLmPAauzNQyO1ZTtxnrKIKP6FOB5CVLXe9URmZPB5dWqLqELOu
U6xYWE86nb8fi/g7sYeINbJldE+JeVgy5meM8dRS0o/XuGJ0/2rZL4GNXln342vo
qqB7m6grJW6G1TbbZdj5YfPRL2oFzB5whxbRF5TzHMC7IWHx3duKP+LIVYAJ7o0i
FUnXsJH7iRHy2QV7av8vdMmCSHdTWyoAQv3PBT2168OtzTOU0qywBDmkCFQMtG1H
aLAOHdG673xNLpsR5/Tei6Y933aADV1ofaHl+6WRQhFIdfdzzfiDWNK1voTLaz7d
04Qb6sPM4VzlCl28StQ4CYVnH7R1n1iFFNxPvR/eWjiZTQgrOhz46QKDGiXoI3jJ
nXG7qsZErqOhgEtu/ZN9QELMeoeRCMpaRP+ffEfWLWZ7BXjcvIVggCqpviY8PbK+
0sqr9gaEhsABKX3PwSSFb+D2WxNRhQbAiRV4Off+7SWoHYXxHfMMaxzbn0N8ZJEz
AUPFOQeQsCuhDHwM2lkjNynoYbb74MpmdRhWGqHhgnqqBZvsWkUxw3Od2FVX9bNH
v2QZgv5d5nC9dxphEi1N2g6mWBUz00lQE6KU0uAG87x1CmyG88iA2ypcrKj2+WM4
0eU7y0YwSOozl1GryxQq2uuQKibRrjx0DX/G6ZTZCXW/lCW7KJRhPygvmi6/y2bL
wLX7vEE16H41AcN722rJVED44qHi92EwWx09npvnaynEqhI5soJ/ie6pb/xOgMu0
Y7izHfnebWU4dQpqvtpYHKVsypeHkpYSlF4Rm4Ye78hUJPP/G2veyOoAU5S6hdw8
s8TIbYAIIGdxR6WZiU3rsjgskHGjmTB+eRZtA54AiW5oIt1k2oGSNHgktWZdY8Yj
5dOsphuStARXDXf0mDmhefJ/HfGO/sBzNl+sGZFcUKx6gAshqIKAlpD5XNM+Nb58
yfD5gHCowI1tmLqibXhTkFAClC8Ljs4gbL5/z0RKiq2bJ3j6GFwlBSV3KPR5B/RV
LlRh8kkS3gXNSBoGj2jAPOuWCP5xWlL/BN2lg+57JkeUTz+GTcqPD2ZbwrZo+Tcf
qebYqaD1PALsN02SIr+Ct4tllMPnsyVim4TpZ9IZMaI8KcOrjhpjKYRxQjadK/qT
sNR5NJpJ6TMa4R8KZejgWYS5PrFOGOj5LEmrMkDcMO9ewN9aRMZ+un6U2MhPJNO1
qfRarfedDQ+dD691545pI6e2wB0NQTq9BaFenQYiXwY/1f2GcE1ZU8Hj+2cLbAGY
6tDg1Fnl5t9Wp64kB3tgEGlYnYh4S29hHoJj9DWTg9Eaz2N2qP3cKvyfAP3tG8me
lBfXz2DNc9ifv9BTccu98JEAEPGN2J9opUoqWqN3jpZCF844fSA569mZW/e4Ir2l
rBL2+pFCkZ0H+Kd2KKmFl76buSx8jep/pyn84XjnEHrqDlaJ53+AROdRYx+/14Ed
BI2zymZ4JkwN1RRQd2bqW8L3HlA/VEuEl944dB2OgOLtqraYEVRCwH822jj2mJrI
W8VwNqV9C3bAyCUggVG+fR6kQNKoxIgOxjwEe6KCKoD9GoqEo2GU3y6X386RH1+K
dVLA3yu1CSuUpqacICES1ijEtjkyO4zxpVNVAqMVYye2MnyoS24qYrxxHI26Oexc
l41eXMMBwoHJS3CWfNWPUnk+Aj4Nuq/hBbyWkc4FH9g/sW6olBPR4BaQYKCu4yhh
/xIZ1OrCq2qiK0VwgljWB7kgZzhJ0Xdx36j8BUvUziujWVx9+ydtk66xP7hl0kCm
3HpN2g3t/BwJA5wh/wgWpTYW0tPuqROufhGx56eTh5FCx641lCfwY/6q2+84GWv0
r4neQo9HTHnXadbtjn/ZzBuBX0+PuTw1bR1Ql8W9gOQYDPJ/WeSK6oVrl9BPbeuC
ufAArA0ZDlgpb3s0UULQepmxifutLXAuMa9v694b78S3y8wGvYgCzAJVKQK2nZBg
IKMF/7TbQPa7ZmlinCVV+thSzQ4CIObDgMRxYnJHL6TnLSTIscFSWlNS4YbVUzwd
CEHlIHhn+ULoVqv84TwaSWscPYYFuSWv/u8TT6vqu9zcPM1pdBHsosSDD3fefNFt
mAzPic0v6Ok7patr9J439R6zmQ9PlY9VwfgDKtC2kI5R7Ryg7xpS85o1ARqWxNZb
OEA38ms3Yl0EjxbQnRd5SAljfk/iKdw00OV/fFPt5v5UFZalZZ8Ldg3eTAJUBLG7
jDlUMXiasX1lTHJww7x5ZTplAaBkA6YwikdomJDAjnoth7Z2lxzcA/sc+qles/Q7
MKtsZSbC7bxTfBO48cumcO3qwIiKlmRuD/RMMTJ/vua1CPVeBolwEFENHAiyG2wI
zGcuxohJhVte4YTZaYT+hddU0khkG2jA85OpDYCtbLZcGkpIL2mvWIShXnlcAC0Y
wPnWgTRnugdndSztOJmkOUIKQkxsnmwrSxajh1NHOAjLgNuYADqNwY7REeV9sB9y
ogoG4wxVTqEWVU7w1yAoUPkhELL2OUQ7mvFe3+W73T6u8c9LOM15CQlGKn+/9VeR
Sb4zJL52K4JBmye9cdKf3BGnwq8LBmw1g6xX3442tKpd49Bxog6BXixKK69BB26X
q557p6fjN2m0Ylhk8FAODR9uOTZauEEFs/Z4M/b0WXi3ZlOmYd4AV5CQi+WjX6xm
cyEypihJNZII8PYSAqN6O2pvwgtwnR46XvY9zREGBXdPYCmPHqBFHAsZvHjCS2zi
6bAZv5l3SqMEZHPBcQVaJ1X1UaIsGO0wtFAWw4N2tQ4LgYZer6nijvBzOYFKyyOu
9KmtDe9RObjN/Fdg/lJiyvmpxK0BJUhjmlCyhkzi6IpAISaB1wbGKCxrnzCtZY5O
D+iqsBMY6h0RqHvce6xJCvCKJ4mTTJ5NmPyAiWubcMgrjO4w0x+QCfQDyM+wVESi
UbM8W/hGOgxgI+ALsxKJGT+JBOqD9/N2Otw8UGrXjgzac3MOKT9lThlG1ePmeoT/
gKn6uAY1g5hAsJaadYtpBp8+vfLoHefv4JV1/1dwiKwMYRI+f8OZguTBa9pIjjJ9
j4Mn66wVnqrsMuHCXaXPOO1w5hkByJxIdOdOQl93KIEYqRoxuAVX/uriKjnJdS91
CLQvqPEv3Pdh94JMfwFXX3tSftqYkntXJ6loa8aK8arCaERktI7LjtvrILAO2Igj
b4Jd8T6HZyEV5BPQsAfSrrMz2lr43Glh4Qxb9B7DRxPLfiWPAm/JRQhDXMUzsxnK
fTDeOKI8bvFL54+C7PHIi4eVzCtSnZllUOf0+x6Ry3K5VVSvfV3XVZt1I1dIHfqF
cA4kwtxv88VKE3/Qdd9R6j0y9qhyXJLvJkg8XUS9QWnZs9JruyGk8ZyFRTx58jO+
CdX7BQDVRzjD6cE0oG23PkIEcoGPVIMYJEERUyNpmeOMLglvtx3ViAqqnATg2cVd
f15YQW8B3szMLtnVN32QKYnVPzldaXajNjlWeamhXJ/1NUwKOGEnIQo0q3k1vhe1
CYrDNFfb3s8t/4LPPuoDfvlVhFAa2PncayTBrIxKH27xWvTYDaJ6sQ5LO/lKiu+o
8rQLofEYGdfXCCCxGcvQorRQVCKyU/OyKeeFkCdungMHIP0ma0v43ZWVjBVrhSwc
Gp/6FR5uAXGSfI2OQGyGX3KS7oyfPJQ/sMObUykXLZSlVbLnP7g0qA6dkN/jZNrn
BYrlwBSnHpf7Ud3c0jZiA5tfBlaksX41GtOrWsrKv5ztKzdnsRmKj58PUCkCS7XZ
7pkezfIP4E2Y5AqO5q6wT2dnPManJP+xXrcAMN/QmvdfKd4xQsFpLflCmiSG+bUq
RELEkiHmKleMwdq3KVDe0w==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TJMwgdyCpusZjyDgDaoErEoOTAeR5XKcc4VdbEikA5KUABT9mmDcUHHqPFEGoXdY
WP1zHC9EjRxjT9B+Kbw22bOP3GUXmgLYHksZL7DLj0XfZ3Sb6+ZEGWHntc2IH7/I
nBiBl7HMI8Q+abXoYGmrkEqISxRHr+PtuEyaJ/R3XkPuryak9kSBXvC2JNHVrSx2
MKwPqWynCTd5E6ubeaYXCjt2ShSxb0TsyA2c27YrK54hEDhI8qDZIRMRa3zT7e2q
qhZLcM2mJpF5RTwPwpOlZXTQ/B4ZvoWfcxyO37UHW9d/ogDkSuRepOjR99DBdYj1
zlFhvpcUEmmipM1u14r3MQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8864 )
`pragma protect data_block
Rn049Rk/cOkwLZLLe0TFi54qkDitfXfo4hzkLs9i9mdCvSJ//2C5zO+9VThCSW2Q
pR5OdAvDMuzi1N+HTv5KGfR+mGvn7jgTvhLdj+bDTo4CJpy5nw/sE2TpNZ1qic7S
90ebTVxV+qN2UyVgiIi1DtG3ORqWLvQzGfZ5w4b6kBcTN1UDB1jgpQ5AVDZksuqR
cSqGEHxxkpK4osELWduJ5/1ukW7HBvmpS1BrrS9VPYkPIGNElbFLQq6U7VVKT0fx
15ZQWYG4T3agHslUn45LfiO3SJevON/wGPYZrz0btsxG/QGH+gkGSFM9Zb3WyvA1
lhEVsnykgPrMB9fwY8KVfPX9BMb/XKNj5PVE5OwTzFF5PcNZJcx92uBvJ6JI/i0E
9PyuheCc4Pgznd3vevwZwLw8Pjm/ww8yDDKmyerS5AAtA+FZZszlgx5GrXDg8zYC
qQGOPslklMY9KYtrkpwGirfBOpkjX+/3bGXVAlfk24hMpOFsH5CbT8R2qT3NiPsT
ecKg2Gk9/5840g+2XhP90kHp7UOvMfffkZg9MWonYF51criL7F4eBGOGXJ2xmNyh
3d72KXgh11tOVPeKCgTFtz6ubSg0rwtp6Zy4Qe4d7Cha6bbcIGn9HCpjfx+8O/uy
HW3PujpHXOdj+mI3A7s1tadqv5uy8zvR6D240IHLOhDXNxPo2vWRXP6irW1ROv5E
Tm9YPa1c0NP32+HUkG+dOz5FSZ+40xBME5B7EKA1AptFFSQ7f/ArZKi13PezUSda
QTbkJqBKMnhYbmUecNaL3M4IFHG8AdtuqZuqcuzDSrq/+USan7pkImADD7jurNUR
UoQSjZwjUsQTKfau0QKq1onukS8UjyfF4C+87t4cDQm5HLSCe11LSMQd9UgJ4RIT
je3/s3V1ArN+n5kKetS53ZFub1w7teQT9+pFag4sd+yXiujUwuweoUKue6KyWl9j
e0L15u2IF0wxEXQ/govH0565vx7lXZuShfWBSStHsRw3pPlYsNVVgEVhPNs1w+tz
eihqBSTngEd1e6+YxVSCedI3h4b03qzW2ezppi7YTOh7zZazARDcDSl8cmwI/qtf
GODNGubuIYjV26Pu3GCnm/Scl9wHJea5kSOTVB3yjzrcj+b3gMZu/3ol7rtl2H0b
RvYqbcvhzg3M8TiNisoqelkw6fCOR0X1oGsANAwYGn6a5evuH2gDB4uf0SHPLCZP
H76u4J+eh+KMHagXYw5oloXlYZVVIgN0DlDs50GCgJjaeK7jr+CKKAPO6oYYetq3
ITle5xMAJCxsu+KopzH3EXC/6wcoitTEyZhdB/KkbGKN3qrBOL0RMgTk3ov6hsCK
1Hhh4raT6wCYr0BrHCuX+XgDxZoFHRKjE9X+eceMnSnFJMlJvTvgXP31GaX4wvKO
kGIIFi8QakDSdfpYkVTbkAWrv/ljQBryXipbrOVzKmtCI+3UU+5JdKefp9goG98B
p52gG6/PHhYEgtHnw6JWmP7bRrrEke8W/l7p2Quf6baHPj55QYZH6yEdoNTyrTu5
utcQfhFo6FvqNBw4DE9SSX0jy4elKxf7iI8zXBmqCWWcQDj9Zt0BaTOoRNCok6CY
KKYXfJenEJK15HeXHgJp/7DjEPS37rZ7qEu2JjsI/aM2BlIEcr4m5WYJ1FLyQ1AX
m20kS/le+p5dXEcxucYl/DY/ZdkUFDAnr5JL097+4jBPayD76NGN1E6dmY7+Uax4
tVgMFChTMhYoZTwdhIyUVKJqayV9eI80/c7+i0KxDPUZCU8MwFJfHkhVLnajy3UM
hXZp2sS3qw8Y9Sm8PxWIurbsnI9oum2u+h9auhlfOkUBwLoVevwYvQT2LiwydJd7
x0p5Sug1ZxwL26qi/Tw/whimz3wdjyDKWQ+KQ9n3we8HURhsgSiWetPBdgJbvdT5
1/iv8IeywH5Bb3I0PRHcY8XrfV9v3wBMrB3OedelZIb9zCATrh3U2DPNIUA3+nlm
wAYHhh5g/l5xPihtQM+FWnZnHEeLkPzWBSZHuty8OKiQz4CBEMhbGvzebvPqssGH
Svr47jbtISHEBPVs/HFTB+Ds3kyljj1JwSg8UrY7Y/UsBP4+2MDY5NT99PMH1nlS
MR/XY5EVPlpejdP2ONhh0unCCjpD03ohjREn1eg2xV8fw+Jo2PNjQQx6TsQnAdlt
SvixfRq5VnB6vD4Pa+60KlzNRt454bUmtOBJbT5cQMEhGZ98UtzdnZQO3QjWEJwv
SCLNJExb86maR+AvxkVVBjw1rQxEVaNySRyVIKOUMng/l92RaF7FDwfijhPkQd81
sZnsDaZ87RqwMIHlbfriqjMkVPsiNN7hNY+tiHMRhVPSN7zlZdL30Y7d4D6oDgXC
gg34a028p2H6050kq4OungLg8QmfbnIv148CAHO8Wd3LzBO9teRTMvSg1Q9JwSsH
GjFjPcTcAj6xEH5x5aK3qg9p5ea5RanJq5TwqMeHq7qHoObHJ5m10EeCAWeXhSb6
iMMnWqCjZpwuqmWLcVpW/zGMpgLlQs69TPTtI8HKpslbVhmEJwIFwPnS8RWAkpWs
H26A4JyX+fN1Oz+03X07maud6dXghG4z4vVGQX6Q3hrHlLB8AfH92d19R4bI1oAe
FAVRHy597mhgb3d3e0sKnY0/7FASmbXYHr/tM5EDYDO25xElVYVKD7NBKNA1D9vf
fVcQZtbNf0aQnEDFZono6m5a0Ep3Sx80YH6ZmAzsZSkUfvibNlp8XVA5YIvrJQ1W
TlV0JRHmnf7awvK0UqZwClHF7S3ykzzfrAXhkgOl5j/7U/nAX8HBUMJWx+9slxTh
U0T+EOkFWwkQXvQ7LVawz5maNDzngADo3z2DuaOI3UhMI0MRi741UlmeZUD45z1R
9Fiplo3IcVRRxFLiwkp0egHGmRL+wAvPVi8Y+Of5sKUV00lbxwuAwVc4+uHrFA1E
BjTPvk5j/cgAkC8hC5elmHJvVNVbfrEggAkxbQUfAPLIfLeWfGLS4jk/0USL9yY9
4IC5C41OVvjmQhd5I2dscE9tjWrf60+CIVYlE+LqUxH2AVOlLJvHJGK3HY7Zyi9o
7morFx2b6lmgfS2Dodf8CmXvei971t5PYbARdQx3PO+Z/jrZHRNW5zzIkCO7qyQ3
D0Zdr0Goa/xVbzqqnwJgAz8V9O+nMY/EGpJxmqQj4hM+TLnS+A1axOY6VLJgE/tT
3IV6WljDGVlX6ZwdFMFwq5a5BXNGrxxoOniIwIf/x+5YWSVC9B9SIO0gr7X+H9XP
9pMBgDs3cXLIjYzlAQSM8ogfFH/U7f3D+9OYgZkGWjlL3lNFJuSGWHMx7LVWy+pt
oLkjXna5NF7s4NeHKS9F0ScjLAA7ce0ZgGxdm63qIV7WWER1CQXsR/At59K7XMEO
wUgvR4UtRzcGCjJdGTetO3aSm4K/XIX2pB5G1m3vgLArF2b+zUp/WRdlKr/WcIBP
Yw2v/j5qHzzICy4bEVrxlWDDHapHVIAUITk7W6zZEWnZzypB+9f5CJdFnA1qGdfe
TvazINw32ut5srMMXFgqa3r0aCfYhX5fHLl9MEma6ofT7U11J0CZIwx6h5vK1QV6
H7RW6dsMFdOZ4UXxZL7niJdTE9CuN9H5AAX7N13vRMhmxK7gT6do37ySfNYpqai0
wrrPRqJK4EJuXdLeA7/KvpGBwT0NMtRRyZyRpygE1d3JjyfW7I+1opdNMT8rSPS1
VsWb6kUeSqzUNHbsZspPtTZFz4HnghbQXNehYPoVcEZZPt8elAMyQOgBmodkSkDW
2bgn5/GLkbHp499hIVb46Go1BEwTFWFU+Re8JwJ9nqFXeV9W8R77X5Byb0BCZMum
teDqUEi1D9ZxfSP3grZEQZz0TLp8MintDni14/KZKDRn0TjeQ/ONlDBj8nNCHpwC
TGVW33q+VafNVHCygqQMyuwjI5bP7O0LYoc/ItvoTfuWKnrFCaklNtk4OHAEfgQx
mXnp0JaI4JKo29W3lFuiSxY+FL0pZKCcplNvBNf0izDMykf5s9eiULT3PKwobYTF
uKfz/2rElJDZc9ed2Hjyp4nodJmIa00HY886pV3FOu8TQZ0x/Y6BwmT4yTJ7a1j9
J883URZxSZ6Al6wyj+XYEFmDu+I52pJ9L8o4ZQu2rCHBVj2FgabY3E7d1nFlVDjj
g8Qbqv8B5EoBf6qR5u2iIWSt5KO1E0iETrzQy7QpIphZley8pADayUEMydyZoeoo
Y8mjIKdgMsC9S+A1waaE7X/kDOJb/7LowJk2MHRngWo2Ivr/A9d+FfnKoGItJucg
C8fnngJAW3GXIsCASD6Od5lRTsJ+1ooZvH97TUYpAI1xe3zxDpT86Hzt8azQvqxD
uZoLViwjhuZc+6QHPK8OD7BrLSqb0t/qxiJNlRzCXHnfLjlv/4huj0PY8ZPkK38R
ZI0hnyCkP1et9u7SH8szmxqupkIPCIEeaHezc7MV0eylrmJcqZ/5dlT38yLP3Twd
5jsvwKJJ1Si50+p2L2qYPTBIJT+Hm1zVHY9RlY5/fe0dFeeYxP9c5MWNPg5iDR85
0Ui4oHIMiPWmDTBLPUkwJvEnBjqw027kMyqvDTGsHAn/XLLpw0T/ZtvD1csdxs2n
OgxT4B05XNyUcdTUxsv6pTOLGqEPvf+fJ9Z9zvqsaHTzk9rQWr7asW5WUor57yhL
m2hB6IntLaO57iJfDExvBdhZttLtKd5gYUFhqEfzM9wERTGtA9irKuNz2okNd+pl
3Y9I5meG2Zevu8YBj7NitgJB4IGRoonDLg5VkhxQvLbYJ6SpvWIkMsm6SQZz6xTo
KJcimXpg6ZQI/5tcq27zoh31vBSSC1qYX+ykMlWBip2Lxpter7aiLGnyUGsjnW40
x021kjizAss+/J/o/KNXCR2++MqC9/991qFiP5EJHDIFHxGav9oGAWUpBt1G55H2
sPfqR3f5CCt5JpGUlVWYyTWza7RqORf16s8WemBy85A06kUti2/YL5w9oJvFX+Da
Mwg1xt0+FrL4SO0yj9dEw0IHhgHAXu8kCrT4BQB0JYpthkS9tSvKJdnUlwf8xX59
htVDzA7750c3wW3OT6NVlICss5ak28zW85NGqtWraxVPqVjLfmLiuS2rYgdI3fHM
np7UjdYkztNFJ4TNH3mpduYfgrgWi9/u2zALXdJDTheW+g63KqV7bQbYR6+0KN/V
moAQ69paFIr59dmxm5kBYe7xj6cF6JSCJfeT8f1wc3h3MkuYlsN9WR2YMmQBEj/V
Jd4tY0W4Rt/H6BHRGd9ljiYXzX55CHOYHjlOZJTLhaYBd47ThFapsK1FDv9AI0MW
ykCA0Az0gWH1+S1jSGgXk6lSRn+qekXpIJzJh7fG+3TcZRCzFqt4fsEUrPbDFRck
6dXvPn+DJWI3e3WRQYrIU6dxxPglfSSrdYF5QJGjYxzidoblbKSjYipEDHhH6gxC
T4PVAePgpbSQQh76JO5g7dl8Ap0kideRRPmBJnzg3zR0h+x+4tZ+ViU6gFOYzMEB
y1CyV4sLF1lCgLmR/yM1k0asoYZ4UObZOvGfJsAKZN2XTRh0BXM/HgCqtQWp80J7
ea4G8pLnD4DFUH4C7qMUvTO3yxnZoczf4DAXgNOo0LDBzuIHzRlK556ieEZOGEcw
s7J3SP+zmA5hwKXMNGLcQrAcu8BRzxkxQRrTQJo2iZT3xGI+dX0JFw9yhAF9xJn3
qs3Q5Gy2SLjQs/FNVhmAVimCKaOspSRSvjWDOQuUY6L1ZJBNibHhsubf2OB4EoyJ
qk5U3c3z0w4MPEcI09qjhIlnuHXMwr0d//yFWj4Fz39+b8aNqLLYigzN6DGOn+qK
XGzfxrLblyU8ykrQZnNDO1+/nISA/VNOQ5Dd9fGOcbVEBKrh5e29lwGqRiNXq0ls
0pSJo8izRvzfqd46whm1kBFk/ax7VenHYbigoNTOuF/pJoy0rpOy6XA4BenMhTi2
oNckvDJHi2XheT/6S0xIhZYO8EeNQf/6t1iRDrwuPy1PCcgziL5fViA3SsA1qBCj
MlX5AdR/ODYWB7pnN/4h2VJllcusDwRqZ8yjCzTIGDbRYQHpcX5IIZSEnX/enm/2
wbS60FuozJiGfqF5zKmaM6DKojQ4rV0yk9P2BnwarW2BrDT3ooTZy4dwHePejuiP
3ZQbedJQseyLITs0KqW3HhKaLYlXFAMt7hkm4yLfRjIPIDd8zBaKEzQ5vXKdaJnZ
ap52swLqPH4diAS+R+NnayHwKjj4UqTbzJwFXwB/PUtnvfvVmFiUn+DiPENFmdX7
N4fpaaSapd05KMr9CM735rolFp8lANwovJak+hl8bpwThq7jhkOAMczAlTgflYKo
mKbf03QtV0yZTLpFWTl65dBuOBY0MSdmPfQqwCwnybrSvon1aN0nT6nvnJ+Q9W6J
8pDkVtUgOtUVnmdm6UQBFC6uWbsLvOQPSy7xipAaBT7q5ydG9yGG5VTB2F7srixC
NHQhCpFbXMchSJOHAh67jkA5KY5vMoR91qc66QeGMzJZqProWyxKB98SroicEGX4
J13Tb6qxlNcm9fuyqfc8x+Q8rQO8re8n55gIMUzOn5mPT933hwA8Uk6PYcd/t65t
BY+Y5n0agxzLp3TI/2g3XKdfjufH57ru+U9bzhQAL8oLumIsOgbC/i2Iva0Z69nB
4NYZFBO+krbZ2Aa0441QXVMgfNMZReMyB7V+MED1xI19C13jmxJ1WFAt30SW0pob
J5FV6biX/002qM5EI+ds7MjHY+5GAJymHl5zI95JCwTD03APD8f6FR+VImzthjis
HuwTBEkQufHCkfpsbn+fzrD8tZaWnoNtxTA7gXI6bKe7Xy66U96LGR3iCraZV8mo
m7qVMmhyvYyhrgmYSZJs2V8c3IoMsskCVMUI//zOOOTPfiPEEOJLDBCux3aaSaIQ
ydQaIZPlohE8rnb6g64hiZ1uzmqen40NIJoaZBEVMWLp11Cv8zuCXw7oOoc4gT96
65yityJIl5hKwpiTSGOx4y6QdA9Qa0+Upkwod5dghFmPSgwbx1u/rL/3WfY87NGJ
gI4Gvi3WywFZfyUJ8XgvOUfMkbFXIaMRxEFbltWjfNsGgw9u/qq4slIt62WaWoEh
rf3TM3qPW5WQJ3v0xUfFLSt/r/gSkJR8lLrn19YaQW7/FBWfZqivWddZqtqK84qY
kbH/1ESXtCGOzYDf2jt8b6qRM1Ku6wIzne6rqBP0wN8EYKMFfIWhF463ItnBXnjt
wutF/2tNPxddLkmMbo/NjhtewOxjdDVpiUGtFAloi6HXOrNRGBCMJK1AGoENRzvP
dTeEABGmtm/J/AKwrvkVSRdMvfKCYpb0kvYYaaZqFR7xNl0gHqy4L8If2uPGB4aZ
+OYXj7Vrhjwambsmp3QJcaqnQLRYBfrKeleMeZ/SOnywE1zX44jbzeIFzFN7f2hT
LsWFYzgCDkGpRChiZqy8/Zj5EOi5XP4w1xn4+bfF6JerhfEZUZG5FIGn7wLkjwLf
T21BxflwVLd7ZApt80XC2g5muipp7zJpDqOpR3v4ISiJCxfoqnBbogQna7v7RDoT
1pBV1olaBPJciWAFuFqgfKWoC0urgfxgsDz+uI6pdFOBujLCFtHX8OtNg2WHQhcV
/+GNRSt1vbkH8JzyY5EmPesjnCD/4CoZBhxcEUfSDZlH6+1z/k+PBCtBJYU7v/yZ
Jo0EAy8QWEbAZ3WoHcxq4cpUsFv8dqyzB6HHOIo7j+fSlDG0hcakV1b9VAHuD2iZ
hTviJNlkNWB2Hwg6O1gHpA2s1aq3fYbunkLKAu9/n5iwhYTm9CZ91z2QUc4+U8hQ
GiYs/+khGsoUiHKwmtShAzZnDHC0p6fVhwwOlatIaCfkOvSKg0d1DVmqJFWSO78b
GHvSWF2ybC+STvRKJ2affqx/iuXvcDSpuVoSwd3LZMj7/D0LDNMEBWZFI2TZOTa4
3z9YM4wKCsVzuOnKKlglfoD/otqKc8wDF4K+xAjysVkqEBiJXqjAEfwMlDJGXWvL
84jmXTbRgDnGv5YaR5nkgzoV05Eh+oOykj0ktZUxr+O+/w/M71j7MHSH8Uj3X6cX
G2S+geBZgPmhjf4k/Rt5MEcQM3K5NvyRUQ2kr7AFKgpRlLvqymsZww60QlSCkvcG
YLNXW9jstqG87hOXcUxEgUvipGX/XiKvtAV8+9SWt4UxBtOzcC19VzcbYUIgXFX0
G3ZAz8A+RECYMygd6N4vyNhkebFGbptz+qBoE959Y/6QxZZu7pPmXyVrCOYkBBZ2
cEci+FathPd+fD9qHuHeuwxFtHzicqcT/s9Eblesk4q2B6c866IlFp9MRzi+Q2yi
c7UsXkRt3O2unimV2EWVE7TEIJtN19W8ZoX3gvDrW+AnClcyadiNYR8IC63MwirW
jeAxBY5lHu0dUB8laMDESmDfvNUGRm7KDZ/tluL3syW65vGgWBEJGUUYVokU/p5A
y6ty/Yb2cAZ/bjUlIcw++umNVH3S8WX7/QYw2RbooEe85QaUi1PSPTIum9gDMwOf
lsN6N1sJTc2szCZ8QiX5XI0c6F9l2mSdJ0djXS4loi8+qzccKyxqjpO925n1CtMM
ySANoLjNyigCmOixUPWRS/7bKWnFyM493f4nXJbMDT/7vNSs7dkUKv5nZWouNCw9
7iR6lEw2jB2FOJ4JnRhERzwNj53DMh3bBoOcp3g0dYAGZgPlTeEunFePlkkfV1no
WD/jxl60f7u2QPrsarmn74d8pQixbaB9QKpezrcO2OlUvaqBmC9qp0d/xaAFzo5y
QTwgz2AcCeWiRHtBgDAb4TXpIvGf6d1Ht3kFR7YJ1rL7wMw5ykfcQLrfQPoU7TEZ
IMlCGSMkJTSywIY3w/HxkZuu9GTa2VpzhIMP9zhJQrx3cYQcdvwEoR06XxG0V5jg
6WSHjk4ma0l7KSiH6CPt2uv040OuG/RV/EqDnzdXC7E6Uoo/ZhP98JLYjLxmiF16
5JJ0ZgOZz90IKFE8s5PeY1wNfqNwGjwnyVzI6KRUePL+FZFrUYxHzDUx08/UHaMS
4O4B0nXmCteCfv+0Wb4HujIm3v6x/kCs+GG7jcrvgjYTP4nixL7ZTOHi4LY9srDe
oaqBN5AXmHl4kKf2P0oD+n2Byl+OOpH4aHJJjvmk/RkNfXFeNTlWNVeiRiyy6h+T
eWaGnQPr1zigyEN8sNi3ZfZW5YWAFpoPZaa3PfrcTuOf/SPfIBnFhzop0hdOUJl/
NMVu941rFnOGqtL0fN2ZYVKjXe1QidHZJZiW/ROrGGHLrN3HKs648Asc3ACqExuw
YrVVa5gFflwpnMV/SNBvKxnpHKmrO37HImndMzq61ef5GotqJ05xpwsopW/Im4gK
glCyccV6x2HtAiQt3gwbFlwziCFdi7UuzU8D6wf17NTFwthqueFYo0A2pLoWe1Qq
T6Rb3vu3k0x7cZmJqlzQFvIk8UjoxFt8UATBUyTt9ja1waD6xMbwY7w8p1SMkVdB
nDBkesKYGsaBAfn+oFr3kPlkm9j8zTIOd84vm/bhDiKZGCNhmpfcBOJYkwXt3Vwb
3eAJeydo0S3I6QSfwzQD8yum/r5yCtGuyBiSCQ4KgrDITYbGQf+VBi5Q2ztRtQWq
DNGGqJe/YRZTQq53/43y/1HYJh9qrDNOezdWwDZouKAreopWhKm7jMkM6/uekWTj
nSJINwYkKw0zMWY6EkeWz0Pu3lIzdrnq+zRY5Tnt6LS7RKFBHjR9ghPlIpSVXtmN
LnxZpx3mMvVSHyZWK53fpIJCju+m4WgEcv9T+FfqwlJu7aBdv+LafAzE1EDIewLl
rpxLi6/LgwbwXVxGr7lKdx5sGzp1z/O1PcBN0hNqDeVhprnXsHX/48+wCdt9GaX4
Q4OmI73kdD5rForNlkbZs00KbhFK16ztk7i83p7b2+bDw2nAL5PQPTdrpbwO9PF9
Dj2+hs3QhYBwf8sTS7lldKpdwh0cf8FjjxK1c+NDYmt//flP/JhJPRo8Fwzw3Hyp
KRkTANItnbjsN9hsIgsJ6lVqPYObWOeyzM3aCpGowjjZgdrFvk3bMTbzKrxrNwfQ
LKaBhxK9l7VuMNhfZAOvZtfrCw29t9pGrmFst3vgtqxWq1ze8kd0Ab/pdn6qNNmI
YheT4fvxVvfxMzEdRIQjq4y/AB2KVwdBk5UR4peCw+w2f+cMIbmJmLtk1BcrE+pb
4ZIrC7pMU1MvypkBsuvnwme79sfk9GmXZ57QkWrpdUg6B0KH9tCBZXvEf6mg/wE8
XauxAKT5cNQkike94IlxBASjDMVDunY+KBLZEqm3IhDWArTSPe2N+eMlHm58f3CG
36Rdeu4CL+Hhxrag/fHL1hfgQoafm3KYqLlDV5m/r+pdNWsffNcwqoZOjlGfvvtn
O2KCGL4W88VxyPAhNFWP3l+dipF150K5pq7zuNRTY3/p7ppfE/1EERbL+r7t1bvV
4P41qTqA7TQH1iTfGJgrYTG4wCLwrv6wCu34lNcpQXyF9pvKTJMxQEpMNEVQ7DV5
m9gp/qqeoeQh5yjR97YSMVMUX/RTwTAyZ4ToU/b8Sn2jRMcdDJkgCg89g5texArE
5ycCjr8ieD28iAAPJ7Q7GLQpyDvMLUIJYZzuxV0d5EaAkctKKHuVHV3yMQWbNov4
hwlYiYS75j43MgYn18HVLP47omPFIBcmfbU3uXdJ6nNZVWX9+5DvAVr16peY+Hnr
w1ZR0qhIulX77iSoL52UxaEJEfOsl1U1trRGcavJdaRWkePYq8fb/nqiOvHOKwy/
Mks4QLhgIlCLyPKXKxPUYdFWog+rjVFijLl/qDLIq11ir7fKCKj9rZKNQ6lL5Z2k
Z++URTgzpzxKUTD0wrq6ZMSKV98RkXy3EM7/Gq7re12FL3mccoD+x+m2XNjFqysH
EBjFuz+HKnSwnUQrmQz0Sixc9oK5HFxW4BjPyufcwyy/1MyykXRdDwPFPHNcjAzX
y+EwCzEc860fZ9nG6NpK+gowlxkrRD3PcmKGZHu7nhK+PrCulnYKG4XYklSS9vlc
0bJBV3swF2KzFYgFYBZvx/SNwP/Q5gOBHH4w87xXfb5oBpIcXrg9YhUkZvPnhPDv
DtYMuWx929HNOMUC/lmqanbjpfstqcOQOVZw8ljUb+O0rQxPnm6KE36zpQg7ICdv
xUOnuhgPhY95QVqCrSusrQQq0WVS4E2/+O77OPHaIG45QGSROYVfRgh5WRttcQGr
3PzdMeRUrtwqyfDbo2YAFQzygbZNYNz08OUYH3VYfycekbuyTgtQ3dwGTrMtO/oQ
yagL1mYt8NbATTdFXww3ztMcmE6oEjKtCP1DLStDEbifG58mC3kRwDReCjExesL1
m7YKNBMnWS+2CWc7jfqjaxyZuRa2Fjek2I5D2rz+EhfBttVY/BowdBmC0ZA6mFGS
lNmt1E4+2PLlF36/JeJx4kKr7EvURoeMUhm+4dWJbapOswa/LBQXvvekGZIlr5H7
7RsUMnSBK2UrjEEYOFPavoPD+lEamR7z3bPP14DwBR8VZ2/iK0w+KPEqtfdKN3jy
l5P854Lbn17c2bwHfTkXZJK+DA4o+XnRAyKhQO7PG+ouac6vRpTCY5ib1o4PSc+f
DJXepSeDPGTlKjRXAMRUsFZ3IpyHFmkShNcW3IF/JiQZPniXMvP0ljfiPvjEpr6S
k0acuLbyjjFbX2rh8qq7s8ek0h4FPv7ABwurRPsRrTJLQ8rFIaHWzSn+g+WY/nZq
CJ6L2S6twpEpumn2lz46q7XUTGQJkSDP2Ujj7nTCSanYBVJ2Gygp9i7NDVodZ4qp
/Met1JPNmSI4JyHuVHAYSCEPDr15YCzeZBYXtiN4G4Q=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
G63ImOZMfsILHrlWsF87c1k5kB1AeYW1+GpfgGuP+7wbFNpCW2XQx+HvgxTi7u5L
TnMH/6YnS7bao1j9OMSWRjan7rHZ0TwrGJzDUwZCLM4NP/O3MGRdF4tV/8ZkmuW2
xuc1mBfO47KR10X1mktLTlG3aWRRWwv0evceh4xlN0FE6C56fQR9Kk+zLHYq97WD
Gu4m8TyWADpxQpVAKWBwV6pGQzeQ9svIn+qXEzFUpMxjBx1OICyPTicdpO1LpmNU
7KJpHg9s28Yby1VfTM9UC9HzCtj2A3WjQR0Ojo78cA2Oa1UpsJboUqhPZnS0Tq5+
9aOqhbuApNRmwugF2U4Tmg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
+moNvjYHFtEFmw6TEXYHKyRXeINBIdgyH3mLA0AUvP+vb4rzKJhZX5XoZ4X87Gib
FzFyejS6WOOfRBfyA9+PQEFVh8kQqgCLzwdjERBo+F9K4gzUAk5fccE3hqMUHn27
VpV/k5U7NuAQmn1zf/xpZ0Oj56g1Nwr/mJsa+q0qINxrDDa8X6yc+MTydeOVFvCi
QRNsBhry7wB1cRrU1M+Bwzj3HXVGKkmKgwWZ0BPPoeOOiVWiauMo1RTDxMyk6ffv
bVDi1v+4/6f9lgIQaWbnEQsfj45kQGA6xxQVLgdvTGJLyVxlo6HNV6FANuZCATDd
XrLoWAAkf168NV+QtZonux7Xj1zLwAFN971ZOeShQ539CrZnIJDm6WCt/N65KeTX
ZgSJI6bz+9myCzRJCeQjW3lsT70OV+peq3bMZ37PzcfThDRhnvY6hpLIN5cwJjTz
ISpVVAxExyAoDRDjZcBCad8wsRhJFbDdkfYh9kjiehNuBxQLPGheFzoIAF6D05mr
Sq+DpSCSu9M4+Wxgt4HnR3SkIwwRMK7PTz43VMNSHLGF/6n2hfKX117lPqS2+BLX
ImLHh2Tfwq6GXCUhISDlcZomnGuJAmC2LKLE8rN4/DxIbFs79OxcF2ReBW8T4ymb
xSSPpI1yyZGB4CYVQn6qvoPGoqK2LNOlBKfSgMAdH/ZkvH9WpTmd90pIERRkTaWs
ky1vfOIPXDC25Jm+QS1tnud4xpe9k4brxSTAmu7C4rHBWJQOdF7q56Y+rV7D5zQi
ZLYfmf2R8BHV5rGP19DyYHvvMCGqJu4hGOlxekaBmJE0gX5xSCt2rzu2cEd58Xqs
oy5hCmyPtmFqdeYGRnM2+L3J7pjdKdJ0C1Qx5E0XA22TMeMlqWsNGvsTcYknwge1
0mfgIU3jmKLUyCtC34vIGXOAHuxaN5S9GMzd0H/9NukGBnVVrqD88L/OBCUqVMay
3LkaSS0qRW7m/bq81FhhC89jdc/oXb/HhK2FTnbggnb/LvLbSDsDRtharz9m879p
3a8J6zKRvsdZgwe3rTZDXA4tELfNgLqUTaBdzOzl/AzeaCVqfkVZ2+bYGaAPnRpe
E5pCe7+Enw60H35WEdttuLwEnDuW/tkWU3opqy0WBJ8F9k4TapCmMDDpMUfs39gr
4KvXbqt0V5x9GBffhZoL4ZT6xtRRpRRunyHjSPjqPnQJUiCHjdaxhJqtt7K5Lesh
DR0eIFA+nQkGDwNHiSAi8/NfIs4Lle0EPwLZEgtnykLmHdOGxwsWE41jVRca51A4
KsJGuQDG9LvCDWnpxkTNCxyN2kiq1XtLB1hI0bqIg5rHxlCqN3vN333o8pgGeM9U
lNGsainVET1hseM9bBe9sMJH/ia12en4jmTZD8yBt5IlLu8GGHeNEazHL2iFNOdN
pBDmhvyKObMdo3wUWs/GNex0ZF0B3nbJpCOE2wRUt8FS7D8shftuFE4+VlIbIJyN
d6XexIF7pX/c3eaL72wpAIkVnvvYXX0Xhm4VEVnn73abCzs5IS23se1Qq0UDKhKC
z0ni57fCq9WM/Wm+WLYhCA+AcpXD2ggLO0uza3MBu3KodXVDrne/OKvowQqrF30T
9syugWRV5FXytE1ItzqEGpjOT4grTEgdjDVG3QwKTgcvvRa28DX8OtLTDB+nGT6n
7DKKND4Gm+3LDUIPG+LtQV4hsS2seV7i0pMS3iuHZ/d2bELHikcMVnuddJtxDL+R
314PIfmJhQVKgwal7X1fHEPBAjtP7MQmfYC2iIhcEeL5y3SsJdtawImbES6G+f9i
ERftBkjb8RngpoTEZety2DV9riBFoIh2DlBlBdCabc79Yo9aWGwNWWov4E4DNnGa
uk+0RxnmrUTBlUcmcsn78QDROJz232hc5U5kfGk4iWrDo4YKDX3nZAFajes9yCme
vJYjbtHoApadhIv2ksVpbK+tYeQ3uXWjpxVOPvisjGsaoiFjRYse50cHuJ2kzYae
EYmmQfLhIgugzuMk3dc+IZmPJuwPfxb1p/imP2IFXyExR7OcE294uhQaLYEva2Gm
O37UEGEQxQjV8lK8UxhVPb8326fDvXuM/kt/AXsgq3LPHenM8xSLpr7zukXoo8pb
DwL2sgjX8mfy+AsQwnd0F/UJwTUBX/JXPcG2+cQNsfJwUhylD30/WP3eBws3cVv1
0fpZjRyP3+0kY9usxCXi+ZpBXbg2K6k9DaswrcgP7yK1MdffEV1wVdwY6eZk9baX
WTlnX402MnY6U1WIOugUL1HmM425AlN0/BxWfR13VKUU+tF2B8c06GWsbaGBFOOU
2g+EF8D9ldRxYpQWBlcyHewpOLnslEXXFPqy1gnBl2Sv1U6N9n+PuAey7YSLyzA0
PWEbentld4E36hnK+GDsSDSKVya8G3qF5yz1q/1EA5F/YRRtWMq7skVwrkwBv1kB
CLuyIec+baayg43iVxLCfcOk+nM7ysdponP0U2+XvR3+WXhN7dYxEpNxTnuKwDjN
QUgERhK0/prPL5yQUpjv2vSR/VUv1A4dFBGAt1kE4qGnnr0BfsibhsBjGfe4eF3j
nAdYc/SCMGz8tKZi5Sue+qUy5jTE6yktiYC44qJYbNkX8VbexfwhNpa8W6z+ryaR
hAMM+1GcuPj8fcQGgfqkcUrm5q6q2RMpLrsY4S7vbIQDTo8GBZsK7GrrepUzjiRZ
DekG/o5UgNMbpoBZ2J4eOVhtLPqXYR595uaTO8kUPAvvYXV+GU+EO7SmtJq4fnF/
dlBGi3/vG6lSAWElV+JFaRKG/PWoRZIIAb2T5Z9jvMXvvYdvS7phRHN/HpD9OrxO
AhAyZMhHrwdxyio2nEhfVPP8YzSHoj7qrFJ+sbMOyQ1fABVkenSQWeUu1GV1yrQl
hoXFrosjtGYCV4tk3yUZ5gadClv7dBAgrNahemSZ7mKznsMGbPALtR+NZtgKpxlc
hLqaYC1Xl66p6IMhpbtJJJTET2GVi+8xhGaNs+733Qg3/+6foz+uGrXgLVqqKPAI
y5r81UY2shRhyTBmlrRUkeuKbC6/0Kn0PERyvKPgDRXSoh7gwiOcWzfq1scKffBk
Fy4cgQ5LDQM/8CWF9IVlUh5JQhDANe9u39gq+e3nIDOn57PFbSVsVlgCvsctnF+L
uGeGAvFhfY2/EBsmkqGAaxyAdNxXMynnzSHqaocGPKMvYhbkru9WBFQ0DJPgKsMN
ovInxGUvH+4V7SCfNFUgu6UFNB7vhgHZK07AyiXetSZZHwbBF924X3lYnb1mVbKr
x2RQwYdvw2BEddJAQIN7LsVsd+t47BXB9/2G6SBwxZJacltJtDZfZRZqC+culeMN
YMIyRkQO4l+SzPNYEL56DUK23BNTKzSbroa2yCzzmUc04+nURDhQuHr90Wtv/CA9
R3XsWvDD4dhtWzB4bVjzA+ou82STnHZJ0D2W68tEahAcn0upfQKsMULBPz71JNBM
Z85p33u/YxXeXVoIvF3QIVzT6NqQ5ijQThyNJuGC5KWoBRbdhlTZSht3/iYhpMve
LxFHmKg849X/uJgTwyrUP1mSATQjmarYWPZmryW1q3EJGp6XGsz4q6f4KpcVaEoI
BVk83Kd5pAzo+yQ4zsj6ylPaSwBS92GutxMco9nqwiR8u8rmzyQ43gAKkIMGfoKy
2YiNl5DCmlHRsIMl5EfqnoyXUuQVZ4ew58xVWDwdxADaj4anLGzSEoFqNC5fD5NC
mMv9LBnBFlgyC2WWHWszgS9bvgjFYt7gFpq7yW9+sH+FQvjTedUIY1UokEt+clYV
moLaRNrbYTps5eNLtWk9fJNMoYi/qXITr+MA4ZkfHqQUrCaNJEwuXvKAhXpb5p05
Uf9hOMEvlZ1+Tm2Cg2i5FlSxiajwM2pdl87WJ4IkS0+dtglhGveCVMXMYxzJ4Hvq
UYPfMnqjWZPW1VsB+ZFkINmw2JntIZOQyQd0q51myM3sy2bNX43P8ak9VfWF1vrt
POByiWCj0scaLUS6f6L2vl3/ho+WuvuDudxbSUJMvAb0aca0rKxbmhTPyR3Ti3rc
5GY1zKVtlaotP7KTbPwcPpmRrXVet4GKfE/4zPvIU1oyIrK8Ev3X0E0WlVQcR5mO
VNTmXW/62rLUal9GvBf0dPPwqHPKnI64JxEQU5/WmxhDaer2sFJXDx9tJx8aodD/
vcC2GEPocMdzY8LubP09dsheNV2kJQvlzR23ST5l4BG9Yfzi+Ej8v6Mpcp5ogHHS
CqWsn0gCnjUX+oPWcvujSP3DnMDEtrt4VbizmepupHoI3yBsbOSP00L1FqPOTfNb
PqQoA0LTLZKtsF7kOg0mD7H/ocBIoXJo5PmntFXXqZkBBlKU+Yg67cWeSgdSnxpr
el6ojwAB6aZUFifLRNZXB8wfQqIzkl/gNa93xW9ZQCjjM+h7/0EvRlhEbheGNndr
ZHmRNOUjAGQtC5CM1LSIT7pxIO3hk4JsbEAlw5g8T+vzZKNZN1Yi56Wh621yuEIV
cJTWQBJoia0pYmtTcuGSkeKPGvCtf2S2tswQ4qyOM/IxR4GCymi8JTjWyTRw/Sax
fnwHe7kunEAfkVvkRZ5aQ46gXTbQtdqSAj0qiq506T9bq8webM/KeMn1n7V63oI1
kBLDhG8iv9YFd1UZnsNaDZEFWQWa6/4gTJCyP/H3UyRcT9GYnzFn6SlYaDPQ9pq0
IebRinGHzGc6Jjp7DN5ta2Bdp/iRnRTx2DM0dCc0g2iVayb0IWVTWbBpHx2DnRsc
AO3ISJYX1TBfSkkIQnaBhBiciIad87HVQV1ByaP0O2hu+B7cvz/+UU4l2Mh1Y27H
hZ6q8orIx1QK0cFNhRhjjrf8CHb3PNXw/W47NKqmJD6fwq7vraCscDDSi4gPa39Y
7gBILpM8VE1oN8tj8msIBQFVBpFMZpP/7XCQXn8G09QnVBWVAkNuwT/eWR7XnZpL
rBcPjiRXnC3+Kpj+IEpAcijnmB9o1Ut9K6EWWOyNRGaGkZ2JiEoLcL3+eQlydp0z
Ymu5vZ3+wCdaFwsolD+NSD66MJgOWgPAYnrNy1tdCkj7+PMq+hQPvUkKB90bkGMH
W9sY89xvMvg4axueDksV/uUqSLzJHBrwg+Ki1cwZP/ZvAhOc9F8mJUomAz6s9t0r
yslx6XBnIBLzS0Q3AjzsAT1IoIGJhCkpw8dzZtoVMxs=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lXAxZLkFO/s1cN3zRVQejzzR31lqD2ET5zi5gmdXwBl/XUXEX/6WDY8MHthryPEE
+htWOfottRrLvHeUHuJmTBhwEsoNjV++14xcb9IBs+ZppNdXQoqUkKCdkTU/UWaz
bVHD4P18SqJLoUMx2m/i8pggTa9uUEEEFthtpCuh7f//CgjYSvOR0njNE/qOjlkT
Qk1KnXTATblqApUd2LyGsqRK/L2Wb8ygeZCdc0Ili6eszCKKLORgkMw1Uu2M8sUb
YnJ9KDEVOo7SyvmYNZCgCLDeJEsP5cb2CMEZFZSislS1kF5F3HxHbeDHwEu7uDLp
yawpEGWIssPTF2kLQv4ukA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
/mVnWyjCOfkvG7LPw6cKHxqLDN6DWI2Ye1bJ9ERUt8WeQ7GmPAY912LCxU9H8yCr
XwcwxLxQoQ1iGdvOxQewYM/neDQKSX8U+s/td7aLWDl38MQK7DNLdafNzqlH9Lrn
McJYguxKtbnbHTdjIbloKaifNkIGUbXF1AhRfP4+S3Rw779vvDW2ishIyELvidB4
sdtAe8+SOtFcAaXAj0DjafbFjJ9sPEoUsJ6JSlAiXwFS6Qd+W+y0yL0PCacLgT3X
QduEP0jp5bgtqQLOJIdH/bWmcXE4KsybTFxOQ7K1kz7qjrdJVN3HSOvdrwXTl923
HJJs/u6vV6B0J/VFgJ+15lYqyBWCH/BPTQ5bC2SiAKRcWbYqYdjejOas1tU2KSk9
NmHPhk3GTAOhlx6BxVp1tbCu7FbC0fAG+zZEHWGTUl51s68KpomYaueBIrGZb6Wr
OKSXFUn0gYfzJmi6i6e85L0Ot7G0pQmAYM798t8AyGs4uTp6pKaEMlylTmXpGnEl
HvxetaGQ/g7nrSt5kV/yXKAxMekre5GaMlle/UUGqeMMri3kFJm1or0PFMKd9Yyw
WjCMjAnwfKTEXUIJQs7m63TsMUfEZ0AswDqDVb40PiUSyYXtwPIrI6AazfQBtupJ
dLhg3USgrm7iF5Z56yjlCFj+7wljFIQNM7q2uZa7ANp+M0nGsC70STSI386NqWHU
lQgm2b4vl8ClM4jhwX67olnNM1b2YUHo56iTw6W/H+PUmmDBqZrx3+sqhufRZSjx
GPHOZT+uapZ4VQU3JrLWu0BBQQYsrkMRgFFZ286lmv+waO8udiZ6CSWFptV13gLk
1VSvDbT83J48r601sV35ZRovHn0UxnvwIG48w+jDCX+OIDDyvAYMuk/jYHwFw1Eb
Ii2Y0NiQszDFvd5iRSNTvDCOMoIk4E0w2/2ex96Q8BvVuB5us1PlkZ6eI+L/qYiR
9iRxymC90Ke3SmAnHqp8JaYj9iYdMTHZhHNJ2ISiqN3msHCvnlvL+B/DR/VLcJkO
YN5OitAWkp774KJBwYWYFJ/38n+O77BhukTAEG9/bvYizZGaYE+RaktpF4zKoLi+
zP1uOyH5OTfcVz2pprdVForfBvuq5UFDOz/97XhL/D52V7l3BXbjn65QmneSZsRI
XcGvsOljGHdMc0+ft93+KWb3VyTZakNqDiZflk0MxLdMQAljQey5Ral5HqwDYrj8
mBZdg1a/OXqigTEeXuR0D39+4dLDYHGjRTqda1y/DPiGzZ3Kb/5zumdFms5lSZ82
Kk+p5gNJT4FQHhWxa821xOVbm5L0BbannMYXN6DnMjU2B7LYrMr7QP4nHnh4DWdH
ForhxdwMkeqST5KM12AzD11vrg4dzDbb7tB38B/odcRgL2F3YuqHeon8DxrASdIn
SUFWODTtC9EjEWQzSl3sfGBlbksqqetP7A7lJ7eN67VKALgeM3gTz0o21kpHF0Oy
kV2vI+POZUpi7d22BTNXQdqb6Mp72K9pXEYjDdmCPtAHLavzHoMifBc0pJ0F/MvW
RhoyFZIo4HFxO64QxXTyUleYE5pLryCZcj+1oarpyyNRUns6n4sZJA9FrTLswUX1
iiHJcLaK41jKgxL3wtIcRDmkulMPIZ6QYt7gYOF246XoSDZxitFOryXaKPJFqktp
8hFrHFjmawcHMfSnGiDIvAGU4W0+NNrcc3U9PiL4SqwcvJugVIWTd70nKFXJO89+
4dXRdcPRs1arbtuOhz/FSST1zXY9B6ZAT2nsjgOFUpErEjiqyvcIFXmI8H+7rTwC
6NgjvJ/TuXnFe0iqvF/ZhS8/1+0QJLWyy6fLIbyXNu11PXSY3HOSioXovl+iDaoZ
KW2HYoRQ2q/HtHvbGQRUSLf5Rc5axIp7fZhbw3E2V3SEHDZVU2orwF+EddV/dqKv
SP1BAzxSdmAoMNVusTUfWAyg81pPgMNF3OjOST+buwY0xUhytvMq+xzHOyZrMvV+
Ph7+DwMfLVbaDojlCTvW0ZVJxskAQtOm5fYC4nvQ8/F1ipxVLrEumbFFW3Ybjz35
fwx58dx8hHu4QZvUjWF6Xgm7rS4RTGtOCNj55xKhJOroc+K6qhSpwlCq3Wp/YFBp
/s0WOar5UI552MZe8q6j5eWZwMdxAWSXqXFs5+UuFKxG9FB6tK1TEM6TiWFhNMjb
vuKzzQdidl9Jz3NKNNTYMrwL5YwRNsdSCdTqOK8gpsAPFqQo7EPsCjXgOxFd1KcK
bFZ1why9H510BAgK/gV3BtmmY3wXr3SKOZPUaWqyLiOJFvTjO9uFE9SWlbB33A9P
WhFEmOoIAIZTUbXfcwOQ2zuvTjEngjc9DnmmAkcblFm4WNkdOC5SRGI7P0zFrDwj
Vd2NEt3tUyON4yBt3ZhIUqmK1YTZNGPkj9U99R1711+xg2dCdOCau71uwDlnOpZa
XsSWvsboGBoYMiX/tVS2JClxmr+svURT1S84f8EXGl8Xs4BJXDaqnx4wzy6t3KoM
khNFWg9SmC8+ml6vD2HI1Jed6IQbEZ5rGast+zm0+5xWomjmXq0NG6wf4CuiNPqB
C9/SzVgvVqXYZdZuXOBJOCvg/KjG7OQSMSI885ftKtz6K3wZp0z2iB5FhE0oZdAX
6rVBfjIp+W+xFCwutbMBt7gsXUO0HJ8wNp67w1zOmM1wlWV1O8Ps3PH0Ee8QU42Q
0dJXKFW6/HvNvFKYBCikJhHnutJFIHWrA2OxP8x8mqsnRp3rGzBoB6Ydw5rgP2sd
oQSS6/R2Tph2bpH0IYvGcDLKXcOimz1lTM25qop8cYRINkvr2g5B4jvz5kJ7wHEm
58NRmFTxwnwO7ut2mbnzeDUCqNoyjhycWmy/Fsj8ziFyLLb8+hKRtF7zQBIA/ejd
Yw1YlyYh06RLWEerI1ACWBp8YO4bwQ7p/aAN8hKLh2M4mDbqMawGXyaAxTtJKG9V
izwh+EXmnN3ZrF3C+JB/7EEpxDKvOIJrNlSKJCYd29MMeH3DdQhuQ1CVAlAPofd5
34ComgEmGCkCe9QB3GvDuaTIMeC1DIKFoGFILgHn7TusqobBsV5lmYFre18prYb7
Uq7xZ6uHbh8Yp44DYmZiyZAN9Her2lIvAtgLQOkzb7rOjKBcT91GFMLeSMXhbqzR
rR7Vj0zQasjAtJATMdFWjdWr10Wp1HJV0Pw/M+PyfHtfJl9m/IDHaSbCIWNa5FHA
Byc95vR6kU/fQt9oH0w68g4eZqV0i607YhgJkNLDKQx3ki9nqcrphS1eFsq3EaKx
KsE5SGI5mJ5O1+s89HWKRRty3bVn1mVEqdmQ/LrLM3JeoGqHiMDePk8WtGSjI59h
r71QSaZAmCB8v03iDF9v46zGbRMm9GmLsgoCZleQ2KgNOxzLF37NLgZ4cmnj8qSp
uedpjZRbm1t3yUtAoprIETtMUMR5b88bs+6kuJ1Yuor2UsxUAM4u+IKKo+qXO4Vc
R16hFj7d9jMV9vhgUnbbZ43QJ9lEGGCczMO/j0KUdUWd8MChCHXlPMTwOqpno2rb
9kekVeDYqD5LwmO10CBYOjf5NszEg2Lcgn8xfHeUSEKCsi1yzz+SyePDptsdsc0f
/8S3xezpjS97qfQibWVTwufxK77xv/GdRyqJIr9DVnxE5KufyilvJDucCj3TYxFz
BBwg0rLzaTS34mCObWJmYK/0lv1NrdqOzpXGs4vURHdjfY90akZKjnvjDQYpnH47
IewZc9IKy0mu37baf8gF8+brDxHswyOsTODg+8aKDQ/3+qa9a9vhU3kIfJcxbyxH
ju3mAfUVRDPUKvDKdahgLel7iAE49BD4Nr7DO9Nm/bl6ZhmEZTlr4mXiuwgGmf5B
ZebA9Q3y1S1Ytj1lPmFijSGyejnta/iH50Akp78vIPIWAIAqINcfSBbMvPxIK1Hn
7TGoLcDtlDzP/kkH6bOCI/DdrBylzkLgen8jmvawiDopGIysPzqAAwMiyvxRnTVU
HaoX2s8QIoqRK71kSJZUrcWCVvvSCAJ+1J+rMySby+Tzu0iqwzDeCYvFc3ecXco7
wGtTApIlioVoJ3N9CXJ/GqLBkNl9GF2wNucmRIVgDJw5fqW1A8Q0EPv1dY9qooPG
br2gkLf2gKq4FfrUG9UjrddbuTpDYnCexecTgU4zObkPAO93XfE3eGmE0AnB72Dl
I+0Jxr+/m89T/CA92TBoIOKkzzYjrXY2AupCIPmfU7URnILUz2xxGAkgfO5J+VN/
YcZceyS4jnwd1ZwobxjDwiCrl7qwMj3gpjZP9C5xFk/Am1o8e1+WQfuvs636NV3T
rv7OFpnrAcFqsfVN2dI3XNKz0WsyZh1Yw9UoGssKMVmfodPJP4dJuHrdkD/rS1AD
zAyYXy6m55pLrsBuwMrMqID+wLtf9BMOi5yKNXzoH61zfQ5F4+UTDYqmss8RnOm+
rU+YblHuFNmRf4WM0j6AYIIdWqq4SKQx09ewaMqIWPQtLkP9A90N8Oe23FSdwlJW
JgxzNUDWHexP4K23DXRC/czW/2aWi6AgypJQ98CuSXtxVp4F/J2Gp/8UW9jyKIim
KLmJoIbhyjs2jKdPEk4TQOJxI3to3Pis8ddA5JKYu/Z7hR/f6IusMPjlTXiOVMg/
qZ2fnOXkpsDAT0vp5SX6HJavNk68pepfNmCW8om8w+jdPqi3tRfwGcrSLqh0q6SF
8XtXsT8qAg0IkJRIB0LBCu5N5eNWcCE8V+KHZoWKMIDiop4OYzoOi/yWJK3uInXr
54QLPsM/KuSefW7c/H9DvRYok/jc/d09mdovXSRpLyyyF0Q62mNXbZO8mduXsdP2
kYJdnd9MnrKkKbMejBTbdH6KNZYyy3EkuoCHZKdAtXeh+EZMq7JX/SSo+3pPdJ0c
iKocvHNBxwZk+6DMhOsOsIE3818B697SlQAhj7y/XWB0tf+3lfvyadqdAK7qdOW3
A0TAPCALp3yIGk3GMR8OU/mpXY7sg5KI+TuR+g2OUrTYp9fZhY7WduT+PM6jAX6E
ACzJgofWpC2gRoSUX3Ol1fI4nJf8SXCr7Os16fwBnFGlLVNj+PlaKxCK+yWW2zTP
y2rcPTLmb31pM/P9mT+0tbQqY7runzcLFbeNCRsrW2KJhHaDJ/c1HwaCy7UxZKJX
e6oKEqv5UyFtmplDoie6/hbH6jsUD8nuV34d9e3Sg6Lpmsz0pVXxiNj4eSG2OvXw
/wydPNrC0k95cm5nq2cBeMqQ9YgMoi0P3vNMxlO2Sa4LxDQ1JwAzAICNHzEDwtjP
PK45EDCH+LB5fC+t9Wmst61PXV0Lz+GrvoupCnEYjt8OEfCH8rW3OA47D3Uo2nQ2
oU7/L6/2U+AGQTIQFsdwHb/M2bVHtsrk7TJ9oC1krErl4XAoYLkqiqtSi7vIDurt
h16yXclyjvDDfW4tUPuZrUMeSFAnwyJIyirGEfGDiZVXNn8adQLEAUTTCdkZhkLZ
KbNwCry41ztz+F8IFfoDcs8Sjo7NMBrB5DnqKZf1BZMKYt0S6cluhn9uBDQX+NFh
Eg40yc5Riam4eppsZruWXfgHc5UD3+9yWTrBzbHTLyRJ0nNm6r06fc/tbcMlFRIU
Uzhw4T5RZuijacrHyIXEkQ0kC5AyzTlrBEMZIiMFmtbYmC9j6dT7BLsZefTFLUgd
SSD8nxoVSsN1nUvJKnS/ljgfcJz8X7uXwSRLh6YZ1fR2OmDSzZEBFK9abKWAZ/w+
Jy0GZzlahI1aipzPXplwXo/qgYjp8Fq2hZ/TNArLxN2dxuAgpZgYVfRgxSii3vK7
/ql7Y9UFXWZiyPLGf8wByUMvVXxeY62T6ZohkeMucqgFXCH5ee+ey54GNF+QurFj
ndTa6Qvf9ycwq3qLLOSd+UCRwZi0bkhMalS0OR9BERHCeoD3G59wus0Ia16Y+g35
j5WYRORJTYMNf6ko5fJ/5Axmyd5FjjlpQgdiIAYif0G6qAa5RTNyo27ZO1s2NpIw
F9isOjHh3cUmMoPMPcLHs133+oZfK/jZBt7XzuxE3CGV7FG381tQo9xVgfjeBLuu
OhQVIOYSZlS+GNPw1OW8jLx3kOALN6Btq1yPtlrnCVwAlF2RvSu0KHSoSYkgMvBc
3GyrHKMVGOzxNItEcpVOFAcmczpRkxxsxN4d0Z7IvjmilP92pB9m6iW6nVtGx2K8
5w2QEdpkpDzj9JduqKaxZR38/Fke8/iHLRxhrWB6CXk0RQ38ca8IdULZrV0hLBkc
PoJKumkO6Wuz1T6+I02HcMGkNzdRahk/YTrce26Z0JQ81quSDmGiomuw/1m2AOm/
dauQRWab/q/ja6xKDJJAlT4QFSrOCFMGYQBTHb3mSnvh+u32RkTzTqbE6CEuxu8C
0FyH3bUmpO0sxvR8jIOOimohq2EaEHjBe2z8tmpf6rrjoEhzvvW67xwvq2dcuhDJ
Tq+AOcS86pz4TeTD73HV7i0BKEjcZwuiOaYdDsoJ8e1Lxr0bPJEduY1RFDZo+gxT
UbLcB2XMI/L1XnGCqBaBYqG5ovc0F8ADWOOo6vClHZAWHka1CzGKHqOsywTq11Qw
ef26qpPLAbKLR/L0PfbeEm6NJHjOteibY4xHbSXMofFLSfrL1haF/9nUrYZgP4gS
wDjkPXEu16yAo7GUBKJUzQVeYhlS8lE71vreQ16rDIKD5bR9fUsN+PY8zG29gxpV
D2vxnFocgNPr3K6pjBVpqWAlW+PTh+Kkd+hQ3NYDxrAoMyUXxY21DVL+FOEXtFSh
xqlKsKIewrQa2aiMGObrQuLcPWvcN1ir84I4/pt102TCbUK1lIaE5PSjiqZZTrDt
/ZOMsv70UTlr1B6Vc7WLhIMrK3N6xRXU5MIURtMRoTd3GoSNVsbA8YQ/25IWExo4
OD/0O0duAHrCIdfQk19rNfRHHP/V5r+rpaqqyy7SQ2YdwhEyMtDnvJXrl/GzS5qr
VbNi5dZZMBJc0FhNjHH4ln8CDd+IFBKk5Ks7ORVQmhewa83k22O+jEnoeFOJQuu+
Q4qnpP+7pKZEuEb9ikl0w3GABkZYmtuNr49AVzZqM0Gl1p8IYcHt7wSpmrKLaRa2
UGoLw6lP5D0ZbUoHEQpBINXAwM8YYugPVBlffvqfZ7DB+VDLT7IqwcTS2rzqv87e
oh5r/l8xanvEH3E2jTvNEZt3dlgd3HYGN1xu3XJ1SKzQSSLPJoTU70AlTDAFcutL
V9MEJjlwasmcETSW8EXuJcX7RAN8VPDIYZezuYjFg5Clv1OSLoInPXcdunnBZqk6
6r8Jc+3fcuaKN9n2XTIsXyEykfgo6TcDy8UQvx8eHFZIpW5T59td3eSgruGHw7I8
p3UeY3lpM0SkVs4dL5EkMAtjJdtIMcCdNJ2k60jVDuBOrFE3wdKo19Q8X4v04CKi
ssGr2CXFQc7crbsyHiIfnm8ScL0GSCZYc3fYsWjUaEkPTtNUDBX345ZABHzWoFvO
ts52015l66ubDYycr1ljbR+UH0Q3nkOHlhCFbp3Khgs9sQQndcntxJj6O1Jbv8qw
XOSVOyGoab8O//c0YgsDXbnqzWNb1nuVNdZ3C6mMcWzn7YoccuKe+bIIULf4CnLm
hW0heJFVReJm8QwdiEVi7qyBSZAN+mGeO7bGr7mbYaAqaXAOSYCZbpPmp8AAV9qw
BRbi486MJQ+Bn8eCOueMFmoY1RRtURQyaW0PHRx7JF++w6jLZFPsTv1COCQ2IvOF
AHEYIoF0zFCLcr+nBqsQm5jOx20I7FKnA4GEcvzr6xgnfLvqj1tvMLFEkXhqkUwX
sURyo6CAerrfaYrXY7ftS7aJo8kRI3CCgOLiK1sZDs1sGYntFQSPftsgGCYQfgqv
oue+CzD6P/gweWrTWWLyB0pcu3ASZW6cE1STS4r+CCEJ0Yvi8Ftn/rbvJOJCCtYQ
BzJQM+JLgYbC5yOJlDkoyVqCutuk7yS/75rCLmKKS4993mEl9I5izeroFHUBSqQl
ueAApQUj4uOASofvuuXVJzNlbvnI3cc+3hFF8jg3RcLKLtIzEg2XJ9KmAnR9J/nl
+fu66y4JHCopKPfoAnoFXqMpFapD3Uzz2UPsWCNuhYxh4V+kSM9fDDi0Y8xT+QNu
Uki8BGxgQB05AvwX1NnWWWaxxrY26Pfw9Or3++nrcxRYByDolKuJN/DtOWJvjkH2
rAtjMUskMDWMnkeYLG156i69TPRWM3L8dSAspLdPB241ZoARnroNfOW3MRd2WXGP
ClL4uySfC3Zn88FVVSd3w3tM4GeLeFI4yEFVINk5eoyXU4J4nN7R7f/WSeuKeYdr
KMI90hg13RoMG6CZTGDTleTUXu49MI52yV6tuQeLm2Zr8nl8Hl5mAl20wWJsv7Pe
8mfRwPUR22WXo3ar7Y5nIyu/srNR3w8v5L+WBKDyGvpW7vy/hUk+GHLtoU8Z6HoI
lcE1tcW9DSietNlxHIfTCT42VddzcUb+uVd4f9dl/lq8uqN5W4QOUwML7OYNM0ti
mM41ylnJZvgOu2sA/KmtWUBjP/lOc7071dxI4ZHRss2jW7q9R9bysVKcj5RAGeZA
xpe5yQEOOf8fUaQI+wlskHgtEcR7zsEDuSAOcRlQ6Cydyn7zdNxeDbX4j9ALBhIx
vJzyuG+56SWrICQaPGVELDxIw78XEqPHCylFVWjPCYlXlY/97ssDy8qCzvpeU6LH
kGDyQ6TXK+zobYrxa93ijfLdqSBaIO71VZDc+udhmIs1ovEgqrawKwfXzZn6Kst+
OtLMfGYCxfGx8UoV01A5RmDnr55oawULVdj9O0WeU1NJg0Xdcsd7V+PeGL4AgF7Q
0sZQMxWAIFcKDWBBLvbQyWQ7VlW64W7Mm+NmZRGI4g1HkDrnMAj+3OrVIxy8Vm0k
UCHivIuw6gdMQUwPg+4X7h/XrIETSjZODZORxLqCXTXb8vFXKQ00vDHYHNehoUMR
bfXXs2zZhwf4iJ1XGRLzzEQIjC39yE3H+Scrajob8umHneYLJDkVkBOWegD3EhKX
mMNDipqOp6ppJiC9Z2lhotWVoFFvA+xF5zBkaSNki2j/tgWRO3g1pe+zOAWLYCmj
6WrTvxd6yrJq+hHsIHcYSpwrrf0+teyRSlp3FQx6KRXlMqQKbYL/BKXtwPrUB5VM
wRZhqOpLnqsou4l2R8Tn/9r+3/Mhr1UPyqtQhhxZcm75SRLb+5PcVXoTaO6kxlG0
84PxSgDFMOBFwr3jMKSzBy7daCaveXQ0gjZpXVnUzWwQHgJvUg3aBO+kxyBR0sE9
39bDQRU8Q2lGJGf3l+1gzv45RyfyGnfxLyqMMUjO9fllLRrPxSSVMLGc+4zzC8xa
L52EDAu41mz5v+5bB5fgk6TiaHUdnVnRTA0O0CyjXXjaWSwq+iKAfuhalOoYnUdn
nwvCKGwJM2ly+CR9J0Lj67pBlKxjoFyNLPmNrtoTuRycvKK46QcXDKp4oh0a1iBM
SQ2/Tl6q7EQLs50So020Yq4pdNLb2lOqHLquT4DqTi2rWl1pwedKB/Ge6xbfjGze
Dg+gcZDXDkHamI1qyK0PHk2vfKOmBhIv8RaH0kFIShg0Vq0ZxK76LV4MBpcLT8c7
sLZjsRxQb5Ngznw83lm9csE2JDcPRoOXpPR7RyvhCQpl3Faco5kj5PZeOqW+AeNc
CrSFbTgzMPry+FL1Kno0YUY74RxdbLsiE2yAY58W6PyNEZZroDtD9OanrxpMyqAW
zphBg13ZjpzQuOCh2V9OZfE6zstWJ2DJQSoXhAa9KdZVYhbUmejUWC028ARgv8Jx
Zn8psvWti9jcxqplaCIlGetZ74yDWZbShKl/co8JO2Xn7OGEMkiVIRptro1XC+3c
FwRwb+baWKshCWU/iMSfmMM2az/bMDabAztv9lV7dPjn+hP8uEHFVJGGb6MYLBeO
97fQuJ/FCN+fInhuwYjqLkjFi/jR2NQ205Tr0g94XLaHNf4ymszzIP/XbBQNgl7E
YGjZAGsBmv0Iy2fK7qcAp6KDmIUO6SOjjidwFu6b2veVYP/JblB++eTNIQ1PQL9Y
o07HpLMiyLsIaqIoZTuKG8Cmbg6Ld1yL3unlBLCuazRFmzm6T9+bt8KybFPupPp9
sWJK4OjN5dQ3FjFXZE9Qq46B7RCLb1Q1CvLB2X9HDbU3eAGoShfLkJOTd5nZRa9G
wiRNe3RyrQN0kvsYjuZKsL38faWn7PfeD4IoGJddAGW+JkSIMp1+tdvlZdBmSjsT
1oEmlFecG7NuNkyKb0pRvGRbjCtFtxzFR2rsKA3EedZ3CRp3YXssJkpj7vdCM6im
a1hRJtKs5EnLYv5ecgeq12Hiqs7lGFB5EOie3TX/as+oIVHVRKo+MwMGYoIR4PT7
n5ne6K38LP3ujwoL/P1x4G8SMw4y6UocdrMVdmi/Ng1p6SgwUVhXB3jqffnU+b2w
1KSKyElNkzYLRYKhvGGl/72E/6B+ilvC3cHuzd/2nueH7S27PqamvZZhYmzCXlnF
WwUV8LHqIWECw3oIgBLl5KIjAlCvCYKCDcQKwjk96fFboFOaofsnRRmLqatltG72
4G+NxH8wRV8vnch5WDED0NVEvSp+upa7R2jc3G6uKbC5dKZ1ydapzjm6GmXqBZuV
jYmphDhs+JXAnAK8GumTTbX330QsQqGsTVzzrrQxphTDuZ1vzKT0J6QNkz9AXEvh
UtDw5ShPI3jb7SH1KQLNWA1Xer62zUVxIz6FXXbkBYFKq0GiIkD6oucOfuwjR1rU
+2oz7rDf0tIbigLzXeY9QRe7GFN+zPbytQixigb0eN0MONx2m97mDE2uAi+fAGYP
aZjbHd3W2z1iU+rUrrrGYcMFEsF8NsVrT2O3337PrRtNRhbAM8KW9Bm9QCTanKS8
zgD42WDcyKZ1//AnPVXvRAldYNZsL1/+iQWOTYRb9Gd3THCIaZ5ZsapvHLYPSeC4
/VEMOTQeMw9EOGKGUSMU95A8cdqZhX/Ik20tMiJRE1AN2HP90CwPmJCFHRbS9ifn
bGBzZn95TFQsBevHX7JA14dBZpu/318v2CX6oia3dsd9KX0g5BcrRN9CMZyRxqf4
HMLibQMuL4xCHzp2UDikGnJnEf1IXQkHMHJHtXOhJ0h32SDf5qR5+ks38bY4r++6
arJNAV9ZaNmt20FQlpCD3P6QLsHi+uKNfTPJEozTbiIKqaym4LM3L6iLxPTeeeZZ
51/GooX+fDzQiOUAgWizVA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BimN85wacJx5PN12QzjxprqEaz+nA6mx09OVrjZxGGk4ZxwytoINbbVbSbEDw4qC
qkI0s3zxmAXnT4XaquknslT2sbN+GUNLke6UaLjEk+oPd94MwF3mkjhQtQeAhLSC
cFd7Vn27ROx7hG994QV+8NWmNVa0cp/RDkFLnKuQk2oZK+7PRbV9pCJs4yQA0NCu
ya9vPdcwJvkejaKELSXXu+5lwbpZzbTSm9T16KuKa1l9VsK0ZERvjM4GcmEN/j+n
9OuW0ksz9+H69Lllg8N5VlYwJN54c1vLiBsV+c/05osf0wZRtLY35pe8XJUVEKFF
Vqv3oRrpr0x1+JWu7NpAxw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10640 )
`pragma protect data_block
+pWhQ0XFrLCVCBc0irM4jEXAeAFqJ3me59oPzYsPWEtIhdDtMcJLDuRN0fCrT24K
xVtPrFqYwO/MshqYCH/kIRtsVg9JrmrN2ssd+cZe0EWMjD83M7bYxvkoDHAETFuK
mnSFkXkXmyPosg24QspAgOd0NhoIkgCFngjuvqypSTX3Tj910vfnBIK+8MP4OVcX
1nuW8I7168B8s48CT9flVdpmmwKPTUlieW2IDU4Uuz8ebHmHRlpTpz2v1laeQjtq
wS28xkR4LnL9u2zTL9FgewyPh480QCJB/B6M5Ot9Xlorhms/+atA8SgIg/Abetd0
LlrLk6eIQ9VIIMKgLI/ZteBFllMac/KEjB4PUw75vUIwBi0PakpRJejmIJqZx5x0
lPImeEkXYKrUiDgRKcjDnt5GLQamgEtw/IPaREYAhAH6O9PVwG63mNbKMrBgB0s8
b24GipLGKmNkGxbTi2ztSRWgyl5J4a9mE7JyV4sjV2fCuxAtVu1NmFN8cTVMy9cO
W5gNbRY6N++u0STHxyFmNjZpd+9RecphLGfdzVMa+Q9mADmHHBW7o0oaqbvQt/45
Cenw9YW9WlQc8at9x6sf+M9kQ+jyEGTXKJXSphge2xmXRqGqh1xsqUQn06K9mWQI
THWTkYv6eHWlWRg+ihv3I7bjy8aQkSI1w6k1K9mE7YcwX+utHZkz6VQAMnVwxiw/
6jKBW3cFmZEOKoqUwsz2X36z8TPETUmWBwrCWpFCo9Wm9VaByW3fNvN7l2H4Y5mG
8khJufjJLYGr3W90Cp9a+BPHyMGw3WQYgXxfjszi034O6vQzxn88UPBYj5bAIf/E
Z07ObjEzKm5GWJGfO+f4iIFJARktyk+KCeFPv4g0pQ2TQ9Hhsn8rQCWVSoHIZPqE
G1iOVh9mXnmCBUezGlnM63kF61yAukv2D8VrNSWotHpIRbkcMfZ8k1aXRfg6sDqp
ZQWJEkN/VpJZahQEEvyNQ0LeEjwqkA3I3llNttuSerOes+KnRbYQTfgncADx7ENd
7IJ0U9Yo3JWABdHFiRDiZihbMUJBnbUotfX1SIQxwPZshn2IISdiGQEVZfaWXGT+
H6w9tAnf+zQeMqYwHU5jog6nTME6xc0Lmh/LoghNKPhO/Q+P1OOaddIVIbCMZwKn
xiKm3489rEE2Ie0bz37fBnYS3PQ0DNzE/G/4MSReUXtpb9aWLWtRc+QzCPRQGOWA
5m9Og+XvXn41dEUkJE2YxNjW/S1fu7TB9nlbs4/+2Ip949tDMe7/h0koJ6DWr6pu
g3N7YA4vXuIxX7kWQSHCaHtDEnow1IsOfMOqhkeiy6mTEN48QgSyh2v/a5osJcFC
3eAEpEHcXDINcjhOHZlHyay12d0HlRPrnOS/x/Bwuxg481JGUKdYMvktzVkLFJnZ
vP2ud/zhz7LJP3E/ubUT9KJAuH/Juz+4KKnt3bMbCq91sE4VK8BI5pQZFaYWwVSL
ikNm0jCspsP9hv+GHYCKkSuoH2TYzGvn+t7JxfsOU/5mh//wXIs7EhsukRknec5O
iVpigLBoQxXakRs8Q3hV1Hpn+39uXtGw9oJb8SngnUyR830pbYcLe0EMJ4zJt8NM
cIOiBKulDOLyJ088v3igP2m2pzBaWmk4q+NNmMbUefXzoEZE61EbCpuX6GvbYaPi
HaeqCyG9B0sR23mPmcfGtiXg6eedvfqzMNsJpU7B050EuCYnqUWIBdNKwj7OC4/8
foxEaKLBI8mUVqTO0FWnevDkwj6CAyENn2LsA2AzY8O7qe5uugqiZBl3TgrZphHZ
6epv3myFfPS77pq/W/BkO+zX8NjmSRXeAaGg9i1vyR6urptMP0MIlNZB4mLRU9Ed
rv11lbP4gwXgzy+Js9haYlYdmBhW6J3ozSfNd2zb9NsB6E/w8b+/JjytS7euQ2IJ
uPpq7FM2ugISlyf+xmHgVQ7hm4MBuuSthMec7A3t+p7VzeS5NKcPYpYA7W4RtjX5
lQ/onCuH1QZLjy1usmDImWrwP1wzcYRnsukG/LXdcOnrnFMtFomewmekEkocWQ/E
t7mqPSQ9SQZIPytWhS803sMrlyP2V/zMwA3EMGODv/YENwPsNtzhyaYm7FVbNmEx
Hz2tNgbl4Mnnyutrw2tKZzGlK06FPA15uAsW5eJthtUQitfr5x1RlJ2wjJ2rQHu8
G3Go0MigPleftALR4d1t+NJx/Ii0OlxdvOcuiXB/AoW5E1lqLQr/xp/fZ4PhK4eC
DPQAbumbCHNwlbdjBJFs2ZAi3E2+aZggSNE2DOQ63gP91cL7Jbu3DJTVoZHfrUxH
GDmuyUwgAGDhZ+hA+mqPqxRiQ2xdxB3HGvnEF6dsS7UufwSqrrVRGUC/g4W9YxBY
1spa5+x8KJXo4eu5L8c+QCICd77IVZ+EF83rD7OfIHExqxCe+h7kAgPx2XFSOWTv
LCKTwmh6Jd1VAm/3d/JIuDbOIwsTfUtULvToZfUM7V1l4uXfJ4ghRsCa5eFkVftJ
di+2vXqVcSybx709Kfvs43dggtcD3pp3EDKPwH7JwOA3D1NwfAv5B1A88H6iIjYD
zw4sAZXF4poZMd/dyGM29IsQzsTIv1LEVQtTXjvnha4T3BoBpBave9y+GCl+qxt+
QraqzlbnLBZu0KP04xXaYKFUPk4BmGy+SthCNPMy+ieFEzjCxL38c2bvk746XKx+
+CtRYPsiXQumQH1Q8Tv1Nc+aiXZjlwx3lhIRPezQJdGdGJ+2NRmZfMMVsVMXa9+3
U4plaMKfVIbrq43FhoDsxBrHgnKQJaErh0swLqeDLd6q/wd2PK8Sv+Uc9X7BkIXg
aDTNU8xMMnhGRlBdqKI8YTeqhaiBfST/eiTynD0vxFvzApEEpd5lHFP5i1gJgbU4
i0DxiF9+eHgBNgZoTAPIrtjx7W86QLlPAzWLK1DZkdb+WkS+Jf196zze28eX10b/
BXE5AJBj3jrSJ72ZAzS6NNHlqWzkot/iTIEDAO6RIJXSN0a7V3bsf8EP+ynLGEqn
6V9bfTG43Zklo+5zJEJYmtQ1yEpBVkDVo5V3D2/93/mNoO91oV+F5CpK8/2Bq09I
URqgu+vB9pU3rZCg98YPYr1SoeGvOCh25DkeNB8etmYsui9YHzAY29JKYbbMc0b/
MOXWJmx9FYj/Pcm50r1hFDqlbSCXUPbSHpC3Vn+oePXArmGAPMfagSnWiwRGcuv0
DyHA8ctk2JZ+mprovxSnJlOTAyZccN1XmzAPXjbvL02YHK4VwYcalmFwXHwJP6dp
yKRehGEC+GsfsNEjzFOXdKnQSnMQTtFTvbC1pu/svFlBEG/Z9KEXy3ug3nXBg6wD
UrdlKM8BNdDt3lZ24MpKIx6qHHErl/20020KD71lU2j2KichIg96zeld93rRlU/6
nks0k4f7aIOPCHMlbl/zh/vT4+D4nDOUl3EVrZyKQWpMat4GzbUNqYCgPn/eZPXN
M0PEj2twDYI6PH6z2UFO0tp7aMBFJfOd7Qi87qPoOFjoQ47dgO+Z00bHBYcQwigq
1cmLopJeIN6O10Em5A21gVHps4ArQi0amO+/7BMSfVrhKQCoREm/hqNHAdovcjvv
Y0cOK0v5lcosWYTGzJidat7es6NjxXizeP/jrWJMeEFxfFvlVMbO8b7Dcz9C9Qyb
XDWOvX6UjmSZySnxjuca5lCTc3wC9pruWa0Qp2xM773jh9UDaPRSDOJpcOJUkI7z
DQHCPM+UAdZI5zHO6WgpRXaGtyxu+dU7nPfBZRI2zU849UlImfDDdl42MKEeqrVG
+sqrXxWqQqHIn/aIPG7dAL/hd2W1SV8lYsR5QPg00j9qyzNfCiZUh5OrPxcJx1HU
+x4lUutA2d6e24eKNyOyDeXj/9IxCgNazTRkcdQWtiY+MZER9JWfyghs7A5LgSn1
Dbivca9CS6guuYPFNfdwZKM2VdBReTy5LmoXBefZUC19V36ejkdTNCOouS63wXer
Fq0DbaPw1JOr7SDqVjzAph0hhd5Mk1cXa9b3h3V0Xbaniog48/dQoJpi/r1uq9Mg
hkSuJbR3Xt+PrF27ifmYa+pBHoOv1hFhhxZ4ilP34c2UBGFk0++SH98sho/nH4H1
OPcwNebUR9Kiv9ETKHn2TiwgGAL9cZaztJltvqLVuwM0yyxYZLzjkV6MqfyyB8sN
onJhs5xUmfxM9z8p0edd/qBvTzNF7oOz2Nwk5ffdmbm6FWG9dsRo37gt8C/FQbOi
NEzAD5W1m0AMJmsutVaCpTr0gFCKhIeLusGtn773+LJ4Nerizw7J1IPi0lYqpzOP
omRHFzPbNTX1BmdbU1yBrp58VH7g/QoWshZi0+MPC2+LGog5W7IutSsvrktgI5o9
uUJltlC9bRczlY0g9/HbJG36SvPdEytm5u0PBmyucQ1NnCdz5fmZeq3I/xrq+hhZ
pxFrkFkoFyTuhG9CfAyEFsTbu4Fghq9E8oZO2gcAGf/blI/wrv9gCLRS083NY7q4
VEPH81v11Y21byBBxdKC/p2MBXWbMay0q6rwVcH5MZqdIRCSyXiAlMVwagKRvUFy
tiGIPt9+Xr05o3uYvs6hcnIZF05r6JsTiBlkwszD2UTTGYjJhjQPidQSKZMbCn7F
9mWcSHrW8KTWdzcWx9DqXT/nhG9gMxnAnT6kx+UDHHBFfzurILNnTXTqW0iqWKT9
JQtq0yS99FxW7zAAAShb0FT17m3Uy6gpnkBhwgv1o3bh+UfzDk+Szc8+M1XiA3fW
ATDTKdtNpvORVpqXnm5ZPy4fGIxSxpDhIiMRuMIa1vyMEdZo9ANacZOIghUiO+Qk
QKZgYpuj1ByXiWDqpqLSVO06puwqGLqVWEdIh90zkdcFnpfOxHG2JLe2aOQ6M+V4
/nuBJh40e3Zz87811gTM0IOAb2WKgdI0sEazLDekkYAcljXl06DWOXLlqj0oRrvo
OiYhHXp3stnjgOKgRyg3t3/iUA0WGswu9cLVDokIPk0upp0cylazeCPT/kqpZK8J
qGJH83T5brSvkP9FgAiYs7vpnGk4xXFJEUDVaRO7hJBAPaZKVYi9r029ZL6/Tnmz
NEhAC9rXp4BW+XryLrGqSpT9ck4WuSrCYm2u+LrydOs2LTVbwvfLawJKlXOnjmxo
VDCtQp4iCLPlO2bvU1FEollWA1s2OT2P8AGXLmhg2wNU7ISxsPUjDDO/HKQwFqsz
CEtzwAHkHMzJwJh4ivUF7NeyiGGBvKcVLVn9H2YsJueoahPVO1OHMNLn3/GquCDo
DG1c1CnjBP+vkIgsROLnduw4mKuEUxXKzEzNf73LgtwHoC7tddF00ozzzn86G4nP
mY0QkB8iXb5cZYHXgUjVexKT3mo+vSC0bWlNZjRCq7iWk44GV9g1J8/8cTHkx171
ZT/hYBMNAeblK1E2tirYGgxbYraiQxB5q17Xgs7GDkanT4zRcHW7IDLPx/xYIYFs
7neZ5IrYQUHkF0C1WxJVt/XIcxB8KorqGMRcG0E33hTSnQsbUqYhkSrbUsrgNg3Q
X8KwB00nf3KsS8tRKvocOPVMJlWlsSSJX5qjJD4I/717HzU8AASHSabd/9iAExAw
MceO214PV13NXm90RFaBMViUqQ7Yjn8gJsuVNgcMlbEMYz9TQC7B33WoiZRcXVOS
ICmu7jYXvPfwI0K4YmjAtuyf3fyqNiRVNCKUZfbOR/4evtlbzRh9xEvut1ONKpP7
O1aSnfF4HlkKxL1HiCJqqs82iWAGbW0HWovqdeK9PuMoQpox2Q0yFTX87q7Gsar5
h2wOGRdEdXFl/a3G8avhrLp8J+2x6o3t3akjncw6YGxdub9PWWQOhpvWpuh3x7n1
c/6z0MVqbjR5fvQC4GcMDZBpYiMK6NdJbWE5og1KzL9SB8pwGI4w0SPIViZAuvww
HTlPkDpLwfmx+fvASJHw8/IuUW14Jg77voVWWCoUHVQgBH+4yeYO50K8NYjc9Hkz
+QfNxJ8Bjdk1Jg578NHtXWMmun0Zn79dbvnNa2TicrnMGtmwYQrwYaIYn3bpmSPp
OT3sk3/nbZhLPWPSTn2xnAsJcDRCyrzhfZ6Gl1AEdJmAaL16dGeNcDqGxZHDvh1w
nbp9vdshmbuZ2WPOHDcK2uEhq1eOMriGRkiNbi4RBYT34WLHO2vr0oGFAqMswlV1
65VuE1q6/wvyL2y9gJlau1iqf73dmTDzpEvmQI4nST3CE++hns8xXoLaDXPz5dRV
eiVBqMa82ygZ00W7Io2o6UGzlaKLDAQUQYHV3Ev11cq+lEq64Cd0eNrLR+8qlAc1
P4rmjark3z8pk9uEPUeFy0iNYK2q2A7vhyvpJyOnz7BugOlauXkCr8Xqrs4ZLt+7
8U2qU6VMsjoWBhMPk2PoN0VVRklpL4rqnraS9AHRR72nERMh1yEVQvgFiiroHYI7
RK1p3LNKDVfpChwOrlk0jFCw3s0gDFlMROK6CDfLDOtiTz9Dp6/GvX1r0KH8QgF8
o/bbOd+MU4i8Al/C64xva3ssJ4nPGB5tXuJSIhGLuBGn+1SNO1Bc3oDKzIHvkFiN
ld8qrhh29mJT+HkNVwa/9HneEZjDo5cyKY6Jqe3RF5Ecy5KHqfTwMxOMLydjRt1p
7fgGpH3uV5b4dzCcvYIgWBQgT7HqxjI4mBDJCi6KgweP9bsw2aqDwKUFoM9Im67N
Xo3abmd4W15vod5qv0UYAbVK14TZDIbvPMQxPp+GfGTlURLkPw8W9jspS4XGkxve
vxRe1Q/Z47t+NUY5eUE8GCpU2ts0UNQW7GW/beu8o8iB2bImKrFLtn53sdLlGWc9
g4LW5Ev2cjQRA0QBXvI2vS4j1fwhEd2jTz393pDrlrj0cQ6JhnUpr9FHIGMnZWIb
+6bOqOja41TNsGatet+nM5fqjGofKqOmOqqVs3hkQPmutKSrQ3CkS+ILi8uT/yAQ
n305t9k3Z0QcrGmFHRi3eBUe1O73YJurxrpOKf+An09elFzGve67yBQuqmc6cpCn
HfTclzDBEf5ujGNnzFyp/3MY7LoMFBwJaOOm3xgL0SP8u6TwdqJlqYfX0Uwzd4PX
9r6qJA+Qu4470khxBbBIpN2eBqFlOyH/VFzYSei7WWoXx2tNgJj+l8YjvTLCGx8u
ZPqnjUIDDs+1rA0RmWQhH7FAO2fEz+S1LroPymFYEuK3XD9Zb+HtppwO03LKcXTU
TUfbNnC2CgycpY7V/pWboEnXIqipZRP0YTEx8f/zZgsyaMY1EYraGHAon2WnfPzA
+m5uk2vggY0z6z/LI6aJRtOpcRTbyKkS9W5zoj0nW3iZn2Hi51iUtGm8g3o/tVkb
jsl48I8tFTgEU93+hmW5U2epm+XkwQmmkeaT9uIo5r3fAh2QWJpStsBoFQmoY7Rd
Mwm3B2GUC82hqD4GmYgQ8vtVZrCfzDy4Sm49xz7QJxQGgUzqTjhNjNnUaEEEFa1T
b10HtELq7WM0vzt+hzn3wsdEhC7KHjr+Soc/7W+PCiqjscrLZen/HUMHiB25RCcH
OHSMoM00BGlaKGO2/l4yzRXDCmfhE+6KFpjMuVN4pqjT4i8aYeVCfZ9IZt6jhZhy
qc9skev+zxN8XJB5PKk9wIEQ27r1z2f5dRSlJo2EPgdTVm/3HYgcUc1yaSXAY5aN
bDoqR+hmSCdZkT9+hFoXUcNxCeLoS/S8GW7uqJolUidYqLz+N6M69AffAFnr0bJb
BP5TsHvblxU4pydkF2fCgho4B0lx0RMKBGU5eapl2mqVQLPj9yUBO7KGC3V1Wl4w
AMTwE6jhQJ5tU8esAaKq0VJ/PZNKFidYLFLstRyf/n3fRbz3jVmqSNrejLwJIVuv
Q4rxneO1ywAGGAhGN1FWVgeaZ0W0NzBeiEteOSgESsg82KYhwwXDimTcIqhdpS8O
/PvJ0CYjz5s+iwvmhiC1E/ac15iwZPWBvWneFLHKb8Rir2hhwgZ+pV3eOJ/OTaP7
QeMscrAEwYLBgWZqETwBe2RdRgm8Uy6tF94qRF6pTVtlMGIjV7Lk2WGqN7BcqUI/
fcR+dE6IkSlu8wXKuUAVELi2BWe7qvcjXcErCclLJOSAaLhVK4OCjaxrBRdAEOvB
i+g9EVIj+/9iQ4H9HqvWO+dtaxiVKfEdK6JTVt7RHsRWXctyZKMFXdL/WkOmzHNX
vSeuszCALeBVBu0W4yoZ3KjovfPGrRWxvhRwbsKq6NsAmyOLqIyONIPZNvmqhlfH
/xM0NRHgFLeaVQ+ijZ1+JlVTvwYqEjhq7fHRJFc8UbZE58JFXY/HzeGrgF2EOLVx
8vzF4XCyAQpLFYTEnG6jDo7oMoaFk4gEBJ12LNzjk1UHWWXvWbMRj0Jw+7ek13Mm
RXN9XLHgayviFKVB80HNvqN5H5WJDzP/KQjG6XXNQQpXzfAXjOElrLRZ3F6GFfI0
oT16Itt4U8zJSeUNtG2CMxapca2L2viNHaoFL+CZTgGAzJutRmFKvMDqn/fKtU4Z
EsdnQrxhA3d/PmBtkgC8wKCEvPevAVq7pokF/WjZNAj+pUasSFeusWJKfZoC2obF
GDl3ZZ+t6GAFzmR0Kbp5WpT2aKkaoCOgxHGKBG1jlUPDJRYPWOt5GNznl3Oo0GP8
O3uvQfWxIBMRjq6x8PqpMli+O9AG3C88Ya2niQuZXM9lzalhKidwled9Vvf5VEAN
InSqXmLs+HJR8bug/uY45Endip0R0rhc8pmx7VwmnEhjvdQUIMQFOb+KlXsT6+ly
9aq1CZo8g6Djqja4V0BpiuLMyPWDfZlz3GNmIdQK3gX6GSJ7jQ6h83xisIezU5rb
NFZoQ0bRt1w/LnSvypecGEIV8SmisSoT9V/It4LRmlVGvwRT5llg+80+trlI47hq
lbX40MI1xVHZNyrzqE6Z0b5NCCU6AUCU4A2aAe7Q1oqZTYVFKeWK/VMfsTvUcizA
khQBPA29hnBKU4hu9sUdmbxYZmy9DhFnJefQmTG18yuRxol2SfJQPaczOqOT66hq
7xn9G/CXzUpMC1RlbzrerA3cVXSbnOc8haSqjv6oPr01xTcg/vO++JjRQ9XSQixg
rr2PfYt5lCuYvWzZIDf+NxhbiMo8vYaFWzqXchIaYhMEZMxOf+UnJptR/YPhIRL1
wC7vx+ahkKdusvUS3ViYEyd/sQsEEqAa9Sf1EUXKJixiG17t3OWySLXLCZAQgw9i
5w38A5BARuEtM9U0kI2NwX+Oyc3/W8H6n1e4EGWmeDB+SXDm6GiP1JtHmK1V3BgL
0ydtb8v3G01VCi+/rGI+plfwCDxgPClDqhKDLN/IVkBz3z7p59TVKTWFqAeignc/
/9Sz6r4kzV21wTGu5unKLRG4NzDrrwwaH3lAN+JOGRl/uZ5iZ9WqvhxDF4Xh5GLS
LpGWhDs9sCoUnNjdsHrR0PHUXuS1BU12RjJBruJ7D8BDByW2o/qY9pH33V/K+vy1
xEe0iWbPCA+cH7FEsWfgVDdR7zXVumgDfPhGatPDb4MB2jUKeuGMNqbCtlygNrt0
YtFXMKNTXas/uczxoTXRMl4j2JLvXg8XvudqZZ9wrozz6uIC4Y6GuSzD5oj6en9f
0PQqeUi+1V3jzPCyraXTbKqiHpSZPsLQD36znXD/bKuY6bqIcMTFWE6ewHi8IT0f
6tUvdWMqFcDtGqbBnF2huv8iJMODlxVGFsvWZifp/b5ut8KCy4bR1HUjwZK3L7lt
wDkPcdQosA5LZFca0UvDfcBAjciTHyzm/fwIynb3g/6Dx9mL2Klt52LhMncU7DbP
KPRuk/Bx7VDsk9kQZrDqiBkhVwNBVZs1I/0ESSILvgvuwGLtRve/B0zG5p7sP2Xv
bt8KY9hpFvPZijL4lfD1UDiI48W6v/MC1dsL4dfICokVkGFMjXr9x4lxLwt/kDlW
y36LVAEnWwk3YVtYCilv0o07K1PI10kbdsOifzyhSA/RR9vE490F+eYm3xYa2/9U
jv1FoO4f3MxRu18BAXeWWxxLjt65/VDOycUNua3CWP7t1CEuuED7Bi1Xgp86ZFi2
N8efudFvtlfssI0dJG55ZZ7qRKtxd0fsQdnN0NUESDNu7KTJqm2JGnfMa+f4tkUo
9gruei3DXNrVi/UVgVQx9NeOEM8FGKlWvNtvTKNzS0w3/4Ji9oPxgp1n4crOEm8K
etNGV5HxIwLXQQE/WGOzMRWWYwhT794bkFmBnJPZ2bQBqR0OmeUc2McZZX1DHogf
hiFazDAx0PRaha/Qq8vdTslXpJ6QBKdOrnCJwuy6laiLw3bnFMqubiGIGBkVGNjU
FCvfJsVbCwYXqOdKNzO3tLNOLR9bVRSOgi7D+q04V1GlLPr9FPNnjIAv9zyPeBsG
1nYUVd5WN/vWQQtU5mNc0HblEtLlP70+f3eiUjZGj1tCz/mEmcjMwoTPIdG14ZBB
kTGQ3+gNOpcW8HzjCPakv8Fmb48K3G0A4f6Ss4mPmd0/KZMv21g+XhOj9wcHCiPx
IZBx37Ix+6Hu+vMV7xwLeXgYa5c9OMQfDUmXPFNLzQfcs/XSlyGVG8cpU5RyWBLs
qp2NzH7t2GuftC7MuuWBvMGTv7l92k54uwQy4R6bPhUad/DCbOc7nT8JqqR0NkvD
Dx6yiNLodwr7fJJDEOodmWglo/DYiJlxODwlC50AcwuZdoX6NpauQxuysgNQg/0S
O1iDT/aophLUOPvLHIlNAmtJlSjh57tU50sxzv+TOKqpA18JiEhbSmputzY5bMip
DM6+GvAfqQed6ihKOtiK556qTONk8CPY8/ZuaA28Y9JF3aOOK82aTeSLlEBXJ4bL
nhDZbkHr4UAuWX/+mu45TTqsFHewKfkX5SNDnTAbhFa/uBz4SfWqn1tAeFrbVmYE
1Xk7X5zrOFzUOLq0mhrygz4UYsoxR2VgwZcreCLiL/I99Tw+XEVTdJPuhhtuNU54
djv/89NeBYL2sJZnsK/F4lmPj0GyR4J9h+HQctq2k3m5bJTR9qYjQ7w19xIC6YGI
QbaUyZjuVwUurm5ueguG6Y8zjmb9jQvFGQ9YAh2TPE1QZdXr7r0xaKP/Y9DrNxW/
zUFvqCInqt4jux8iEdbqZvT8tVmSEU+0YIsVEVxr96ulex/wT+gea6h2sSVP7q88
y6MUiaAlxSDRZoWEpnXN2RIy9Ltmob3oh+/aW6dgAUZlfWmXn+2GmS4aaUiNQyXb
Va4O6N4NBj5pxMliUXde6tr9L/d6tS7wOTgKdQflig/0OM+x6NW0j87gaq43lLJq
Gr8H9+hU6k5oDHTQKPC9wUuVWijWFsifRXvLyb8kpsJbW5yYfkw5GKXagTOuRYMl
dt5pzMvf47HA4NWEXwZ4nI5iaGKr9+UNDMFtSnV71zNb2nbd1VbmyeiRMlq6tX7J
QonkGD2a3RohgYJm6loQsde8tVVWE8frJ8GHhZIfOdcFe3pOEjSHRNq0g+IYaDNY
qKJHtMqcYiBoIe1Spri9gFZ4Y9z7+KL0bu9kpw39U50nvfY4lwYCVd2vPViiAH0v
mWnZ7CIC1x7yvlFUFVQhVAUCBC1aHS7MwP27m6+OtGGp0Bet+0EjT8EBiRmWYGNu
j8Ya8DpTJE4GumOnw1ojBU0sdhMb2CGjiTJvz/RnuZOhqN8qaKDCJC5RtPO1fCde
qds/LnD1bNsSwBvZTdtBfGCzm9KsK2sM7bpRtud/lI1c+zKvhOG4d1ASU5bK9oL7
flTUDtbJd0zddkiLMRZzNu40aHfMlpyiMf+r5mz/BHZvHLhzevk/Hhfb4oDJnRNt
OLaWGi/UizCJnz0d/XoQd73VAoD+Uq/Q9nBjdxG0pLme9r17uZqW2vqPJoh+t1rg
9hOrVUzeKT7gHByDj/5sOzcvg9NmWKbw8R8igfQxrangEkL/BQIiQDqh/WkhEkno
ysxkTSklBGLZyN0DhcgE8JvHBWlGFdmKHK3wGgPE+/iv1E3LSqACE0FcSYaoUZsu
dGKgzssZ3OV6TVrExV0QzpIkt/lt6KXX3oJzT05tH1S1iJVVJhjwM3/0zlm8o8gS
CxzeiH7mlGzCrZrxa7whtyThIePIH8diNye37H9BiJhMYEGi47DAQxhzWwMFYEVz
FcZn/o8fGlm4kjAf5XCupQTuhRHttvxJ5pEE2AVF2GBz0rA+4nqGoG4aDRa47Nzm
btxkOb7lDSsXt2ol2gpP6GdlQAtPtpovzdlenQtFPV47J128JxinZ2QPFLwoCQ5S
ncrDDiwjYrqoSo34uJrmpBqTFBhSNl5ErTL3V21WCD5IhISN0Nwg0GhpN5y4cPIx
DQTo/Wq6umgfx0vzEVbw6/tqr9vXjo+MMutKHf8z8pIpn/UqWodD7qHcTIMcZyTB
GKx7oTRlXT1X983PdeUQshINi6usyR4QGUIoZiTmVf/LPJbDGMqdpvAdIBGiwV88
q+5yPdN50OlyLwtOkjs+1SL0jXchTAWTpnosjw+/ex+XyqmJ0QHq+kQnDprgiZ5E
S2rOglpppdgmFFz6p3f844/n71wnYWlTp5nSuEc2kLB1aofUkSPNzQzozKW1TEZA
5JeisZhMOCIlm2rYGI+tXSLr1Zjdl/UD5pyqAajg/JzyvOptXt+nb23YFxOYaemc
9cmhzmJW0bVnh1+QP7FkC5k4RSBpriA14QNnu9B4WcelIau2a0DvsEuBx7JWaODr
zJBmFhsMhtKuQxwkZWaGb0etnjimcdImQYFH9/hU4MHTrqotvrpcMLpdzBZHtYMR
isc0yKOgF9yuFXPewt1wkbDk+D2hqykOMT2Tj7XEGCyPKiqthFVKnO+bDECErm1O
Nmr2YtFxV1hHUPvKwr+CfGx/w1sIf5jFd98zAgcf0pNNvvzwO2Sb3PKQ/3jNmEii
dLI2jkIENjAF1aQ66Hoz3GBVMPk7f9dGRP0XcneuWtH9HJImLHqcYliLTDyE6iuU
lmwDdqrz7PozjCkYcBNZyJsWW8A6ooDuQiax9fTBGrme/es4dy3j4s71VxjeFYXC
hQh9I8156hmqHchfnKG52vN6+bN0m1FCdmvIN9/fmQR3eW9uHqifD5hOlxcGS556
gy8I6OG1+rq7NBKoHpImQ5JMzVggjiyHEbXBBiuBvXe985rxiE7qTbs6dVJFW2sk
cteygZqkDpV/44cM1S4DO4I1pfiZX8PaRUfQv8AcQUJazyAaSLtvjWR4jw+zmF9S
VndsgM88jN3sTR/0y+nwlbthjAoZBFirim2Gq73f8FM1y1TgdTD3bx+LMMLD65/a
ZQb+YebSd2UV36EfnV3k+ptS8VX1gX8tXAQEQgN1V3iS7M6//5L/I84uEr3h2WWi
eihXgibnYMBgXApK6xFGTdDJ97BsNb1j16u+GeH3ocJj3cvOBunTlQ+ZZwfeMATY
mjpqXd9JqJHC6I0QEV8ajzpmZ80PjYrmWWtR3AqD/eY+i99bnKULGo76m2ZRxSg8
qeS30i0DkXOInWP3T3wyspwIplviD6EuYgpaNtsXFgd/XD1/LuJ6jDmj/dmWHsHf
15xx6zdEmF/2iOArhgrgLQp5RFiiA1nz7pUhcRrtiQXL/PMjGAUcxcHwbdsI90cM
vOJI+kVlI8BwLtsn74PCXYub+zMbYh3P3UKCNjYNXTTBjQ3xF8nN/fZUXoLXDcc4
0zcvCQJG6bAOKHfwPHLiah5HUMEbQ1yAKjEo5GXAXOhqWaDGme/4iCwCUimk7dqg
//10C5nR/dZ4h/feb9axKxyKsTkbhyUBJVEsM8j6Y0cqm3Wuzo5Gm6mabteu6OUv
zacKQVsJZBPbwWzWxiOQAnYNIPgQ0eTMPswR40G6OziuR9yJpYK9Ojc1xaBgHAmg
4VPyvupqHULJ/ptQ+uQnXPR5qhXUcl9H0iNnYaplf9UXd+xcnPm0sOPvOYib2r4S
Wovs9QI1o03xSoa76eAHOzO14AyYK5DdA06cnWXwTDxrVErNG4MsmhQIieVTCnfP
GWyH9liD/iX8eyzQbrKPHFDPgFOCchXmfqcL+Tib9ZBAgzYzBrjE3eoboJ+Lmh2d
7LOi9l4CnE3khl1HAZyKqbiUipyZDzm7DTanuVVwRWmXxKtJo490vj5LzstdjisL
8Al4W9odqTxlKL2FsxiL/uDfyC02jl7SVLg+0FcXM2QnKqrTCqbz81Y5kS6VUY5n
bOpl1CUvjp0S1dqwufSrUuUzzEUtMJ843cBvigvp7s+jP7ChFzY44nS1eyTYHXZe
eQJ5fRkTPA3izTge7jyGO8bVXf1qSvRxEeGWCV1Y3IU=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Lypz11MvOD+k5xpo8FGOPbvxuYh9m3H0TNwGkzgKggXgdjyIwhbKxOaD/MMIiDdt
8amijtBWN9sbUeKqS48TlWjJ8e/qFKy1EXfJt8yKcB78zE5wAIuEmQhPuk9QctUU
o6l7pLQUAmN6sGRV4tWYb5qKC5S0IqtOtkZiFIrxKMMm4pfV8VJhmI4IvCE2u8bD
u+XQl3IseFtnHpdIWV80u5jSIp9zs3gQnYeMk3MvnQTzbyZzOvx2FTd7GM684ChN
Lu4YvnnuyDnahu5JvtwswG/xlE53ZchAn/IrtJY4rlpC23YGmntXR5OxPxUaNFyk
Jh/PaGWtmPNeqEG+FZBMSw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2704 )
`pragma protect data_block
LwPfuXMgiSi+OcMaDlhim1JLR9+GkMJxDMYRJGChtNYEG6Wz40piqIXyAeG0O5Bn
HaK4Gv8kFgIyJHFt6zevp29xtJpfvTcxjJb/lFSY594labxolUWL2RYqWL09JD9t
okHacD5LzJp3AXsGhNZd0+dpRAV6gs2Ubw1yThcVWfbDtaMdU1WvGPpsILiU3Dfj
i7pPzEkmstsGY2hILBlz7dWNJLNjToD+uL+Kd5r7dFzsqT/xaHZR1T84LZ90/qqY
gaWgF+R7SF92TuPHcmH/ly4GERJE77Nt7zpaJ6UZvrohr2XPVVp9GUivbKOWpF41
HYEHzmwLX3f2dDAWtTQgm3SAipSyZnYjz9aEILVayCDvsr1PtuL3FTE8dvY8LkZ0
FqZydvwGSFGkr71xhAM9i+xBa51lc7Pw8FBDceDg5JHaQzvaoMWTXbEyKd6ykQO4
QrjbfFesdydBbVN+vW+WxGZjMFr0cQI/cYyqkqw39LkCmRafkdg6iAu/UJanH0lt
YNz6rz7iGT9qG0ye8ZFXnkCWWThF56VrASVLy3hol1t+sWsET8NgHxZ+kpJdyYbV
tID58haVok5AVVhMeWFZEYc1v2qfYuqG0JW1X8DJz3Ks92CK4pI59g0cF51HFS+T
daeUZkBGkmhhA/QP073sAdLY0i1JfReOYnshv8e4QnWXbjltt0V/6GRtoqQQDYrS
+QYp64WN80kk4jlY0YYBS7R7U1gouh1FXwSh+3EN+rSLEnMmYYc7nG2krS3umGdh
iJVsdCx1/qsfWyKTRzGHXnqHkR58uPiH/leh87D2W6V/GNNCxZRyGNKsZ9QGmxFg
IIG6g37mpZvyB8dqswOV/Q0xWUMntPBncPTvYC+pWFq786ZPsKATsyQ35KhYXPue
hg70vQWTBbJScCl41EL1YEvKd2S0q7SneKykKjnG5RvpVq+p8n4xrQRjtqICYFb8
muqwtbv/NPNe5izE/09bAOEwg5j2nw7U3aCFXG79Hmg7YyKZlAQji8ctJwJ++Nry
VqXjydB15ylNfXuKvG59TYfievF1b2VN69NOOVEWawo3Up3/FXTXY26/31w9a5KS
Aab627G+8mngkkJkMk6Vdtb0eghJEEH9dQHJ0RRu3W8zilSpZYSR5YwCje7bpOQU
NFdNsFEqcp2CDp3SJRr8Kp/thsqMo51neU0g6stsDZWB67lRxQjSKotuMJBM4ogy
bS+TjVZxRjtZP1dnZWJH0eEHGU2Tl7VKggFA1evTx1C5i9pxeLIdIGuJFk9ImmDo
SvYrLaJp/uvGuLWto7lBHadRJDL2tiBIEblaSOzOS6ehCwbolSVNgJVNzaVbVAft
qNoqCeDPnCYO0Fxe6TadHvuzx3lbracJci0CeKVlsg7NzUt84BP76cIRtyWaQCzI
UhkBXytiY9YDvhIzvPuA2orn/pnskaNL3Zksp+za1Ky261lId5hDrdvPQv4LwvFq
7nApIipUJGDrvBLTumRvsMdJkKV5hnA1nECVGaGu0VRNbaqizVxfSPDmKqSN+sGp
oPQLCXmDEGvcE0BfD6uAcjBwWwc8PoYNEzl1vdOJlTSdU8IJcRq/6oqgWExQPQKi
lov6IO77mVdf6G5Re8Mk415hAiCR9gf8V0+J+tHnlNSOWd779bx1w2/Vxfx5Ch40
8FBzpMe3pOn5R9BrmyLbt7I3a5OsdJp5db0ItXvaoFUMGTZqUXZYIBP6QvTx2k60
ZQaHc9xEA5iqyPOmdaw+EIjtzq+lAHzzi/+j6R68FnC9gpKjeKFtZzxP91cDptwJ
4nsYuCbvOqYeIXvE3afo0Slb+lz3JgqxuW0xwIsAo+strrGcqdRzXFHv1rsRFfR1
s10sAXzduYFyWDQLu8xolaByZQa9vQ1G48f7RrSqDDyHyY4c0PNYOtaJWT4yY16W
pl+HI+N03Ygie8dpmc4RksuxcHSsNPcpAuGNJMoUIB08BO3V2JFYncXxHOH+d60Z
US2bUjsNLBawTWsH/KpKiMn2ACaFuCDCa5Pxi/GKD6PDDczC8bh0w+SamEnjd+3b
bW6WoILbffaj6uzqkN6QAT5wZuwKvT12NTbvtIBmPiKDuoIKNMEKN2hL4PZUTqBE
iB1713msysvB+G59ZVExwdYJ1sLA5ouK2rjX4rXvPDku6zubltaZD2Hgrq6QDXI4
iChzrkpVnQUUkPkCIPsq7zhTXwfty0pD1hprZ37uY4TzGUxSQMEqZGHR55Dc2f3O
oMz19i+nAAEqlis5Bpm3R3EEJFcxUDf1EBSRH48mQgs0jvxTcIt77VDltXQTK1T/
aEKFFsCHAnyDC+Amj7MZavvrLgRVb8D3uv7hcRW09FtoQI97z4sdqjCI1Zz/DjTY
yqaClfRSF41XMFy0oszRb+3CJsHl6kTo7YlVSwczdluk6u33mS+FTfC7tExZq0nM
QYHwFNUTk2CHWfnoMkEBwIgmRNAQEiqjIvlG4S3hzR9d1EirX22iYIUSL1bi+TVR
Z9E7R2mWLLYxsmmEGDaZ/7UGd1152TOR+9uHPNHfc7IsDRhHxZRzUi2vwex/GTLH
5NJp/bCie8EQT9WZL2TQ53rcHAD0EGuXRWnRUg+TByq6iyYA9jJf3w26txrav2ss
3JMfAbBgSPt1UysYGsq3Y9mrcPduGTcyJNlSOwEh9L+BEVrietIZbqJMAZ+F0cLR
OBXytA6AVE6wqnh2a/hij0x36m4UQKd5Fk5KWPD9wMwf81D0WCiAMfJNsX7DEEt7
PRFrkQ5e/oRp9J116ATMGmR+H3ugd0pAch2YAHNth9GJ+lKOpw6Cc9Exyq999O5+
Gr+bF6Pf1XpNPMX/w+JrWJVYlDgF8p3YRJhozBPRs0CdKdSI1p84yassKfYXugj0
C9wK599Yg7nAUEWaUWK5ZjnyosN0nenx/2Cjisq988jtjvgkVhVcoEP7G4O/Fq2P
dcriBp4x3tBymJYUjw8yK8PlAf6Tz2vqnlcbzQZkebfZ+zUWQEvp46xPAcVjuErW
UoeBb3GQ0k0iXEkCMfAE8L4Hgq9oI/mWZawUi11NYBMLypbwMeSpYm1F4MHT0Idh
L4KS4K1j8ZtV/a3NOGcEDZOA3tA7Pr1MUZAjOfMHbII1m0UBtgDQxTUjtIwZAq4u
cFCta3m03Uoj0AEvPC8vjZxvcPaEnKz6CswwXBv8mHupMXDmniyNYk4GFdX+WgU5
7dkpMdfw8n6xnVvdeQVn9BBoxtDC60S8w+xNkAx6JQiM0OKVkZK64CzwBZCiEwHr
wIfepxfGfLeevkbgQL2ZTXi42Z1rG0HZoykhOcEaagpC5MYXVotG5TVIZA5aVESp
2LBwbn+E+Ix60JmhM8iz//ZL3Y++ILtMKi0O/68h8SbfdcqFtZ3aIgIk8NxaOYL4
ZatHytZmgs80yUXmL2/nVuQsKVuW3btdYgiz49k2iU9TO9iMaVPDzMjfntP3C/06
Gd2V9fmdX2UBcmkZxK8CAfJ7MWWkQBEU9Dqpzqg+HMj2FxeHn41dpuilsdhzP2bD
FDBxQJtsrZGwpCMR3tkHRc6y5B6TKRQMaVNMlIuZNxJKrP/24EVmRTUb/WYtbhcB
tQHLLe4RVeMu5Hq2ua0sRA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lgAdpRyDQEjzr+j880tCwJJ+biRYBkE3F7GgV1SOxdaLmr7e8phuupV7FMkGYYv6
40iu91mNAYU7SyvssPZ3XUt+YyraPNVjvQUXjOp90v67gr42oN6uE0bbKA2abivW
2NlkX3W9rA7KwkoLQQaw66+7O+ytXu4MZeKuReYwAp6gv93Vv88oykJ73n9v3wfP
sL+DcuwNOUI6j9csIB4buqM17o0jSgcAouDaokzLLOarKr9nu8QqpAUJuPpKmf7y
hAXe1SVpJfEl16Nom2y0oj9knbBoqW61KIeLcNhGt9ZHnshVyY5hAJlSj1JdYMrz
F+W2lxGu0Hs32EiNXErOag==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8048 )
`pragma protect data_block
rSGagcsR9f6G6RAPqhEVdstVraI8EKNuQDaGpIGMavqUlFcVOqNwrPDBC6KrKOtV
d0jS1LL0UZhHNQFBzWaERTQeZatfOcJ29mXWL/fKg6aaxI+Ad0sEYyBNEhd0oRfz
x3Ssd/B8YRE+Eo80cRVd+mQLFhT1ik8zA++1sBzCHTwMXAesnSEiqNWVssbriLJW
rnTDfyopRqSQ7Rd3YeAjIo4cl5jvgzsQeiY0tbikuKdo3awji1cPVBpbJrvlH0Lw
2nj/Exo9hdCndWwsz0UcYYexQ5uM3ujo3uuPy9Z8ANw1fyKalEe4UrlzKhVE7IVu
krHKRFYbUqmgCW9fc8nactoI4Rfh5QAoe1lJWzEPOktRPxe0eyqWHIED8J86uiJ7
mVLSSH+o9utame8+R+IIm/TYY2gWjaQiFRKMqAZuaFNiRn3/FXyKzQkEP3nP3rKO
yfcUf7SU4wW+TBugaMMpToecDegKaEEqnmqBXswUWtFFELdD3o4XYKKTBfj1NAZs
BvDoWb90R2xSAMw3ToyKIMgsmWC6WtRPAnTMbTBtqYriHUlDkilg8hrUt2MC/faK
oTpIUeo29nC4Ar76JfBt9Q/HGBh63Ocxm9qUIvio/gmmLRbLf8kBJp+0qg+cn7i6
oAdleWeshOaIZgnfftWx6C9GPYbEhwisac4ztIPrME8Ewf6Rs2TLtfejKLE8iej2
vshm85oJ3v9BI/+ncpfLJnG6m9BWBl/b+nSw9B9rnNZriSnkLSUB103bcXaFBJ8Q
icjlNq1koBWsMf1DjhuT0kLUaVk0CIq3lqFOjgeO7N1Dz56kboZ3QQ/6B84NbODF
j3UmrUBQlLjEc6yXSDEq6UTj3//ttaJdDiN3Ipy6W0DdP4LYYrXcWd+S5DXBo3JY
1iWc5KOooyB4PNtJCML8A2iNZW/K2xfMG6WLcFTVDkQwvZTa2V3KMqvMBAkVRFtg
9VfeDY9mVQNsPwOgMslPJdwvFjQTVyxOIDbYgzw3CJp9lL5oRGbkYF78Ra1ViQgh
GfOum/WVjjpMGE2pH0gMI2fhkFMMEa63gxxAYR7FcIH/xjThzlK2pTjqUHTziUnP
3ldmePcAgv+KE6oNtpnQaVW709Q569gxOwg8GMr3NYJRaTrzY2jbjsze/A/Srii2
u/tb1dZbSgEKthM3jmgy7aOKm4q313+RM4567v44X7cek454LXIDbOFtYWlLa7nS
dYozHEXMx6XOrMqxL1miFKLNMhCevtrHXPAlbMRUDxjpHnn127tvLEJCypB9HrGE
zCdtSddZWIXkaD5Z2Rg87xv1L1v7RoKXWbRXUYNYtdphb0G7/v1UWcYh7w11PRFS
u6eTIG2ToscgdecvOria6S+fI7WIL5Xosy6OoNFoWxEXQH5A2T+BJ7wvRKGw9afU
2jpMOqfxQ0kQLjffpZU+WrWHyzyDgTSraw9W/PY1r6ihZ9dZdxT9884TIiF4kJov
AfYgOcsJcK8wFgnaU95iv4aoA0pQ4/JPu9KDK80KNx8JN9mI/KflSryaOXzFQE7k
QiXVU+G6vOmhgcRwbDAfDNivaSh/QD6gj1DBmYR39O/Xtobh4zgLWyE3HrSvFpyO
/tnMRMVPFE8Q0ddq/qFE5Lg6j9uwvSjtrj5252RT7GcYc+5eyeTQzO9L/Iguvx3T
78r40Qwwe61dhT2X67tZEalbzbyXOvv6UwFhLtr8k7yfXPnBfbxh5GOICuSDcwJz
A08M7mtC2N4Dpcvf02ErPAuVuF/ccIHb8MB7dTFUcrbg7ssMK41FgoxfcbRUkfCJ
/iJZqzOQjiJ6+nwTiYoHlpxAF9MjwJgKFKaWxcOvD72rPc1abbpar8COdQuNJLAU
K2BvVwLF1naF5UsUky60GEVhcUXaxLsY9pmYDZtpPUlP38Z2MEcE+5OkHksuEisP
ufIRvBBRudvFHCwlpt9HxIudIjQa4onkUvZ2YLhkbVvpTN7Jwc6qj9nqkjgyUYRS
UZevEts28PBJ3+SxQJ9awuMJai4t4d4wrVhLNtPWQbKJTGVimicMrwp3ER6s5Nz4
6B1cLz+VCaAXdvJI/T6mj3uLaGJuovLYPN/nrGmxc1xuyZWCQ86ycl4u0oEA5T2a
uXP8LB+H/UecAY7QwQvzegM9V7TU7eP8gequDi5Wh7q1gsCQvCymhnaC6vPmh9CL
5YRDSn2M4NMXZFbIAy8QLkGmNgrMLl7k9Wo4TJvhLV0zciwsr/dADUKNwPscu1zo
1+mPbuN9N9vipj3ZOHRF/vxEK5JQQU0SXsHwbMMHRdDvjPnIG55dEzsV5KFUyxKI
IazElAscNOqwe7rYO88H+bGN+QvE1Zg8lTMVspStudmDhifKLHgNACZ5n0a5iJnS
f1Ndql4RlC31lHiLj/jhC/BPVEtSZkAHXHEU+aZftGrqv5lLDJOc0CbZyWXmrs2z
cD0XlLJi7JvFCdqeXGNKn0sDdwuYEmzNV17koKjlZjQwSVLwJlzjTDv9FzGQ31KP
WVbRjleczLubvv/5mncVkhPsL2n2OyDzMfH6RlPnUunNAbZVMyHf820h3ZCZKd7s
dqsfAP95AmaJiqsxzuiLtGdZGgSN86z0qurkDiN+cxFPms6y1zjypSkr/6UiOftm
Xue10/CD9oV7nsSN24ZVL12O5kwilIn1wSXUsakyLJsy3pLKxN4gRLLg5p1901+Q
L4CHGenKdg852wsQh49fxLjCkPoHEpQRWpuj3dSDnXqoEgtEC6MtqdkvJUkyen0w
DTZ0cfP1iJJlaK5uCd8T/XLiFOyzz4+56fEyjpnIjdErURRrg8+g2Dzkdm2j8d2s
0h6dNCk8ky7/gZLQcAQFzDgsB/aElrXL9XA+m60GcjMgoefe9CBvhQ/Tg6CR0ZVb
ESrdWBK8Qj+P3HAaWjqitocs7dW2VFAbRBhrOUaHsd8mk20jJNWpmGtx13/LXw4b
XjD9hXcj/NeDJiXyVZM651CLNomRWm+/T0Ytq6+/qRiCU1mGbY82AnWI9AyYM4hc
pAP20WTPt9MhNtG9wAtW3R1j86slod6UOtdRjQEmOzKDjx3wosZjAjtEqLu1AjAN
+MbVqV5J82ZcuaKZSC9VA4Am7gC3zzNt7JIJhMgI2J8PIgoq+xsLH2MxgkdQNAEJ
H7tju0XYIHG3YwbmFWpoD1Pn1s4/ZsG+o+hyObMdxdDt0/AvC80pQPH43RmbvTtc
BGB2EciXQ6DSxX0/MBruPegr7v5R82aRrd3VaHGclb85h8gCOy5wvqn6Bi15nwgu
jb12caWhjADQA/QjT621uStBm55JoTYq4CNqLJZeh/Xpvo3xDro3H/ajdVugGfn6
e3HGeEyIucnktpAbOTk+hatGb4Y57OC9OkMZshqXr/ULEW+MTdN5xpMsMLDR7BSG
ont5dpGkuujAtWdGvaNBu4AJVG9isyqrV9KvHV0rebkdvmIsj7rLzki63ATdLdzY
Kj5KhDr4Nc7YKXHcGaPsp5NH+RtGZgrLdmUO+VHV00k8W9r9+109N4G7U6X80sJ8
HYX2jdsVJimE/Y5hQqTmExvS92qn3o0nR+GBRlsC9Wbap4+SuMPNVNQEEP2nEU6k
OoKpkZrpCE0AaJxGS1sPduYYzN9rkNMHuKgCbhAS0BtaHoeyM+b57iHfMz590Bjm
+3BWoR7u8SHVNNZ1KFw2qAc1M4mVijTCeIQUT2WB04evos4wUtfmMCpE5EIhsSit
tVYU3t6og05pc3/5kVcoOdCcl5KzjjwF30axYK3Yh9aPNVcLpJIktdI6hHgKDJgS
1SDpZYRl4JE+7/YbTxHXVLVSaaiFCpzefX7e4CUIPh3JmSPTGRZDNcjy0Y3GWgrO
7N/3mpOW6tr1ze+OR2F30ALXcbfWkof2p8RJXATYr5XcJiBoaQTTYexS/HIJJTrf
dYnW25r3A8gSealKO4AUIcdKZQkG2aEDByMPfpASZsxqjGGnzZQ3zCrDYMqAoUeg
fJbcaWeSfJaJIom6iWnyZS1vtZTFASSjka08lSVxaOw8KVzHV+EnNouPMl6qL170
OLxi32JAauzvy9BIWRVfiOGVueXcp/vXcesRpCC4Arum6sUlwrf1KGCB7cAvcRR3
U44cFaMkb08kT8kBYE8+VMGCFNLAlzLPAqCUpxrlRSmWdWZ1DzZZw6/9Ctrp3gGQ
MtXC896VpqzpSuc8H/YaP7PlPC9qCEeJf8PIncdekWwU6ooZK97TM1JB1hNGx0DJ
n8VRqigN0w8Ap3OOCJrSQePfWtchQFcZilpaspnt2DBMNbyBI69tD/fFoM3mEdVF
tMPnwteH1UwISyqTTbwMLlVuGZkDLe1pJzd7Dy1rKQ23xxCNuuu8ZMCLjoh5ZKTz
ZEeNEP5knjV7+LluKDhoRNc3WIQOCnJjwZQcAe52Z+lqBK2rPnxyKUOZBLlURDe+
5PGY1FEer+lv4hNq5LUx5DppWl44AoEJ7Lojw04RHcTfwA1QQE/PCRlEqN0cn7fB
Bhi4MkHfrypV+3PyLBgYUdzrjt+r6ifwLy/FJpx/C7SEi8p518eVX6yHrE65JMXR
Cs3JWxwMVmwI5f4nE6Ucc05pihttBGcqnUV7twgYrNEYPtaoPGG/iJW9P1JHGxM9
XsvIt1LZ+e5xzJo3/LspUZqoDxAoTc4xsw5A9k3GWFO5i2aWsbxgy4C33JaF5vk2
KR2Jsh61t6okeJLeeXgWz0SxvaErN6BBlSQ28JnAl+Mz79LN88Geghq7fQi7jc+u
3QxpUqwZrOZIMdNdXuMK8gdfYOnYxFCinxxKlZHFPd4ndZlU2aHEyyZwRgZ52vWP
uCweAy+Qt7363hwgT7leIkoRe7AcL1IhsdeznaTT2DyKE8QoS3bNnIfHy6GV98Dw
5vOr4V8j/fSt3FgLZe47FRc9TN1uHvAUW1zdqZzk6ym/Vzd5Py8wHzw6d9DwFxYm
Mm/LKY8T/lMdzF3zn3Bh7cX08GHQXLuHg8Ph4tLvDi20QZJbWca8l6ZnswHeOkHY
R8iOHEFXVpycPMyAUBdtXTcJziae2Pw8Ie8rN18EkTKBNApvYBSYQMIfFL3DnyZy
9TSkSrIMl88oDejcHlmR0nlbvX0Tnc6kWG8YguaupYuRaZCZbg9P+mBinSdvUUCd
zV8BuLaNgDCEEXcwhglKX/SjMxWkYLh4Rn2Mq6r6QEDxjoaOH3xM59mgBHyCQ3/f
+FHyHBZ4mGT2tDSfHSAve+UsW6NSWvjGPHCTXJhggwvAEKZlJirV6QkgU7RUabHg
KW1xmyphblA/l5RFe2lnD4pHbOvbgNC7U0xDW0bIk8eFfOouFQVtapY1OJQWHDEm
RWk0J9tB9Rz8HfNvZYoc7c24ttXRv5GkmNPVw7I0EWHpoO9XqULculz1MAZ9qBR3
HoBJ66sm4OBCwOfC7VHPr2mQu/esVUJ5wsiHQ/Xo3dgXcUlmQKMWXjgHEHAbjxNz
dbZ1srk8ZklYyHdIsOGFadW2e4HHUIUXJDaTqXcW5t8qfvugFAPQ4JIe7oBTRHCf
BdnuQy6FG2lTqf54GeeiWUUFbVLdR7Ssy4XqybY2uIWHdSa2U5+jWPEiPR+6M41b
fQluGjxZetK/9XlaZfqWtItRtFSsTxToen9o9ArfW+taq/bx9AuJpMl6dUWYvJaN
UjB+CAyTg+kBwBvWhFXYhMuJDK3hqTLabKuP4UEr65CT6rv2wvF0FvJUl1M3ikWX
CK/b7Oxz4F/Wn7Dj91Lwk+FesMJZUJIIIgzvHFaXA0Op5QEXYlE0ZDdABNg1F+/Y
iP6eTUTznj9/oYdNnEVR3m1+Nlfti0TRD9PXApTzwg+SiU39Qmcy6DrEFCfYYz5M
9DNu4+BbEzBLX8Y1p0G3EE3nUNbSrNJW3A3ddepOgPxMAfJ6FMTsusliD7mWhPrh
tH32WcxiputAkWc6AFcgyVrmZjzsjThT8QxraaiUu61L4DUTYTflYVgC1ro1tsjQ
KrVu6pr2yZfEQNrmlIuKiDb66EfR9z0/eFpEj9ZesI+fu8FK6c6Gdhfjk6pcATqu
0zcuKa7W53nLZtg+mbViPSkqiwGYrhdvsAJFpTkFoQI7MXXw3D3xekOoFuuhAduG
gU/V26s2gDmFJtP0HrblR7SUm2oX3NJZ0FeyCCFEQHozZeC9hsUT9n28iVShfPuV
cTg13AXD7a3iQEizUz75XyJWh1SnlgYY/0gc9O3Zv9sIhZJpfdQFdbxLvDidN5Uf
I3VqShmvVUb4bLjY4ftBeXq6MvTvnRxj2q5H8gRRPRoaNeWDoHZOZjY1YapMlW6H
P4ey9w5WNPfN9LUjlEYD8uQqOOtgxdFuNWEXHfDMJ3Jd5esuk4KITqzECqOtwnkX
/k49GFEbdWVZ2mEHGmpDAn47UpRwLtogCtgCmIaYZaeRe4e7S5lNy4d2yOcnbv2Y
h1a9X1haRBL8pbWeYMYQKpRG9G+KRwHPLjGeW9DtQh05JeLTdMo5T6kQG458d9x+
+lxt6ijrzNQUIuJQsLNDKeeGu1LCWRnbOiE90Lj2wIb3sN3Vf75hGJD2WgXh65++
CmzCzm/MmHtf5uEkGnkQ6YLgfF1FuXjN2BBDNj4ByFgiAxc5BPqEmJyMcovNoK73
wZLisA4f4ccoSCtCuNn8+nhYAppFadC7t0LpRXHeBIJLWWhaTGpt/ktl31rWH3PN
747KfEL9qYWytl+EpJh2b7Ygm/sw7o45AyT0lTgXP5EztpFZrqROaku1cGgSBE9/
L6KuNJD8XyVRYvK/u5PE8JLL43zHD+3DRdOmyA5BJMti7ut/GZJ2XEbJvJvJGIwO
Ml579gcmuBE7BDpJoKm/9NU3XyJr/5lxnuDg4J1nLxA9Wsjm9HMLWTdbPVHKhtoI
TLvmtAzZB7dqA9w87rfYsqrCGPWf0lRPd8Pg6kgisN7GfdnjrDRI7NEe7xJMaqif
Bzn1ydxZ6gcQ70IQKByByyUh0dueJIbaYaKYiSDm2Wh4gQDRJH8hz6YS9rnD4Rtl
Q0Bd+tgWWI/4FuosRXkbzy1qqhqMlaGAl+IzL0fgW+Kpk3PS1dE57tHTgJwvEjDu
kR+v18qAxOKTEuNjL1BkDS6cKx4uIWf9YhykUJTfTb+Eyrmj24APGTQuS78baRR8
BZTeYkQwNR+5g78pFNYM2x3jt1XwwAlWdwoj6xvtIrH451oTRSS8kI9vuw7iiYnx
J3jNbkyv9nZ/IALbt0NJI+3Qr/OVgrvSxYV/zGzvZ9LKX5Xm+L9LXg1PYGa5Owzl
ex7ySZ/Lt+5IAbaHUIgwkOy5/0hiinBG9j6MYcR8YmmusbIbdE+UTonhWvxlzgg0
n8/HRNi7aRKDAJoqrZDNeJJIZIKfaHWME8RvsKYKpAVpvdCYsuvOgnerwzo+FNZn
/00NDtRJ2CjjTXGdBAd+8HD1jLL70tYhpD1tz9/ZK7EirvXa5vSvtXPsNahw0Wyl
RL8BBE8tBaAcrWEHo95wMrUNuJSVzVT8T/9/ZkMfJQGLPD1j5WeqrW07h9OvanJ3
Hcwpq3oaRea0SYiTUa4RIzrW0HMFRgDUeld/BmkDpecK2OVcz1PFh3gdjzrYcVns
PnBML/akMN2nkngUvkZ3m1GOq8bmIi+wi7foAgqpkewh5K/P2vcsg2UWYuOwctVT
pJxnu4YjycyAoXgx4LfFaYow1tZK36LDIaCyV/xkkRkOSFdxtcdfACYGSL00ZK+r
QgL4zHiRoo53KRkB6tv20zhCnyqpz3BDSj5gOXMxDnZVt8wg4wGeDA3tTkrySdtQ
eKLZgnGEqEigym9cUNE9gyo82Z+wTJ9YHDjrsT7ed9g8vH1gK8nQrr2FHQMWUaZB
n9IeDDFr4enosia5f0QWOv/84WK1dDpHN8l54EFwSOLZkPHnFBrbz/OTGTS6QIpA
7VjUV1pp23+Amvk1eMeBg6vQN1htarSiSw8PfqXYNuc7fN79psyNCORZr9hjPCFf
sQJGVLFU8XzplypA/6sLSRDhMGM10vGpBP9FqoWhj4cqWr0TTAgT6RB+488w+Aez
cFcPMv+4htV4j+BpTCbhT2BXhGwxFxFgJMY6VnuHh4/iwO6LQ7CXauSOk69ZmUSw
fKkCWhrnR7BMqG4RGHAi2uUzTP5U6MHoQm4ZWhpMPY5+lgFQDxGtmm/qW0QsQ5sv
66tnIXYf56Zc+SNv9wJ+505G3SS7GM1t5RG49ojzrd3in173Mv5d4BUXltK3n3lc
UoqaKTQYrgdvxYUNRCHgFSTWXSg8rsc5HCMBRx6o+ulXi8S8J5lwZQIfir/MAJ5T
e8QeDorKF+DGw5h0ajBQ2L8n34GwieQFQ+8NN8YHUTWVi4gHKiUTkEa+bRsBsAio
cg4KXBAsbY9r+2jZTFR2wn04YVhWY/quypgPopEADRbSHx+G2+Jiz6oGbYr3StWd
yJsjWB7iXTH0amjDwpWKXBxrGPkwC4ggCHdSG57Vxc22L3KsZnGi/Ec+Tt5Ex3JV
iHfyrqRqrqlNo0/Fx9OnWbAAiqMkIUMOUrzNtOfWQnh1sMc82OwnD8LHYEsaFIGA
Co+nCq1r5Vp7v8DB0KjsOqhiVQg2VvV3tTsN+Qvr3EUDRjo++u91zltuy7TJKTdT
Fg/roqtJTiWD37b0EdXFMbOMg+xuWiB39AZGKqINot7A5I8L1Krfq/hyFg3YjceD
VAPWCQ/VVyQiGYzJAopacAZrPbUOA+iMEVKL1bRNbTkOcHYHxeTrBSBh10QOwMfN
Coi2X0xif2PCU9IIlH34N42G6NvzPFp2LmUPALdjrYO8rForDq9DV8zA0qx9ZPq5
QexRcdbWlExyRYRYLqj21/E0ziNBUwWDuFQxnIKbDgm0MlEm0a6aBf65eFln3Y96
+FdrhhtLlGcxgjShsGrKgAedli//MotB4C6zNrg997q3YvM+weZutBZR4Hz/FJjQ
398HATPHbOwQkLM3tW5RcY9KXqRHqJHnWmo6mklKmGQdVF7/03oNCyt7jFauCyve
SzVgWWLIp9xykspqD9ntK7SrFZ3mKfJ8MGYKbiXUSPprWHdvzdoPJR+FwkprgMVU
OThGcUQZuZCw+4EDZabzuA3qN/GV7x+3+WCDI95UIqWFphlZZcwujVfBtsBjEyyt
6VQ7UISwgp7dnSpPCGtjX2iv/WSRI87OzqWyq+wQtakoCGMIep+0G/3eu7Ux2+qD
89OfjgKnI97RUO0hBj+bDvCYktVbmEne/RcrCf4j3VV1WHTcJaCm7tKqvGw2ffYH
kHDM3K03RoOTuepk5iISN3xPNe9eTvsvnSSRpbu5/24X1IEpeH7FpMGezBVwQo2w
SgYq1zpAqXFO/Z3vBVUWA62g732ah1tJAdm8Uczn/58CmN20K0kuAUHK5FSHh+vO
HjmcTbrsUbhnRzA89O0X2f3N3PvwnjLV1SyshygsUyKJiLtzjdcX1PtozGsURYoB
DcCm6hjHzbb2PHW4jp7PQpzD9litdonCGBkOxiv+iE0MVBJF3GkpkC3XAaO5A/qH
dK3f6bZZavTgVmnhI/T7rxEyphBPSt4RBnIn2E1H3lg8eqN0NbcEXLHbow/PePVR
XPDpuAAY34POISFLG0iOYC65GQu736XoTWZt2X3JlYtu8TOz2h8wyuXlxlvPnH0S
ZDqugn1vwLi0OWm/NGeZwoAQKFsb+vM07geYbYbhoiYmGvCaz37rjyT+fLTC1q25
PM+43+U04PA9p3M921/bImsUgS0iLxtUQQssaipZEtFnZFckJwyr5d9mtZQkNCFz
+ZLMxc6yD0Rbxhq3g8OCNvGqq5oVlPejg9T0t+2CTWNxrXM2+HnPkFKFSB8L5gzj
OJH4pHS8tMS9H7jcOoE5iZJDmhY1MFtcKnyxLHDYJKRUTozZ+W4uJSsx0nYc8/gu
KHNPMNvGOER58ak451lS9Wt9xfQJ8AnfBWwh7U/+EAU5+o3oUfnVKNq+9yP64WTx
+jvB3rmr0yW1LxLYVrv536Plwv6vPOxzz+YYw4YR15tGn+BxTOUc/0YsnAncqr6Y
dSFEYT8MVExi4llEOJeYczX2v8ksD9dypif2DKGMfiTGmqm25Xp1Wsvwh/7bOnpD
WUNnLtyXPamYeJQMMgl8HqxosLgSbGzDBGm5SWpH2ZbMCtr7zZtxQDn/zd74LvFh
rgc0M0G3X12QQegV4CFTOez9JhfEVreP71CJDG0rBWNFaX41auTtl1/0qxgRAFxl
L9SgfaIjqoPOikd0RLnAJjmZaseHZilJXq6f3SehxSqVwYpQeRr42ZFcCKfXK5BF
GJ6i4DgOimG8VSe43lkXEVUq66RMKgOncUaLKhJJ1hNRdWgc/l57103HU44+2s4R
4lCdQFrofSRTM5wyyy9zUb1kY1/D5wgEhCGODnOyuEAWWi8VKhShCS8SIVF19Olj
BSxrg2ZI8u61j1uEuyN5WJ6NeIZMh0vrc9/SSW+Jp5oDsBxNn634XkY43b2jMTms
mMOvRx4kkJGGP5M6BbOjNh8tY6jOwAvP1o2jOvYsvsgBKU7vnJ2ijQnxLn5hwJGN
/TBEQlLxQNc9+Dk86PFPs6E82oBeAh0AXvOmdr8FIkuosHuac1AVLxQ9Ix4QN792
GWScouLnTs0SrwKMe5J98BD8lM2eNHhqFUpmPua9vAPuvwtacrxgE1Iv5zjV0Nrz
jaIK+EEJ8I6Vs/lC1gCtnhXNgIlV+ifG531wM7DJc4W55YHLQplcJOJU1P0F3zOr
2ZHq7R21SC5/sK9FtfREmud9QpG+V8ymRUy7CXaIvrU=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Ev27hPnMUpQpq527Cn1aksxyaTUylln9fyBny7t61mcoFJyBD5hGY7OSj5LN1CuY
IQLFs5jrGIweByqEhvVeFRUoZ6EayjfJA0n7LxH95ez77oSlkwuT9gBjNYpnh4ql
oBTOjFdLqztktvBKSFPKocIT4GsaLJWymUshJPWFMeZZBiJZ1FK5FiEnsEgI19TZ
/dn+Gf4+fx4/ALufRIHylMMd6nr2AzFoK451hVngCHaL3Wan+Jcf51J5nSo6Zev9
WdhE6uXA7Q9otOw6Sfws0PaYpc3VCgWaq4h5NmI7C3fmXw3c5Ar2FgUt7xS8baPs
I6j+ejO8z7rbw8M3wEFnAQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5360 )
`pragma protect data_block
07qWr1tcqtkR9yxQbouwMOvY0yqFaBcSI9D0kpGWzQt4giZpm5hioLRSAXmVwXxl
en9r1Ceadu0SbLIc6m8+wECFipZ3JBROhSYT6Z4LPpqbdBrzF6Rv5CEJPpT4fjzG
jTRYp3wS4p4w+dNLQ/3mju1c1DgyUmjy5D8ViOVF8uFA8J1VFeahKPezOMunjT9U
SGJYDlmu3V5CVCbyvJXFbXUWgcVJ8YWsKaYjiTXJAGLXYVxANnPGdTI0MnF2jdF+
vNsqQnzkMx2IzZdr16YNWlvBk3lupP45RscsssKAWgZ1xiQ8KMdjjE6glFVU1mkN
dXPPqxwkC7zu/6xHPrwIw+pYNrRbqy2e7PtEqmDOM6a0MPokUth+NMVZrzEbZNXL
9ry/c/8f1lV5Xay4ZNNY76VXVMu9jHe2+B8z3O1g+sUj6Bpg60RfokZagfElXHer
KwOmtQegpXMe8S2pYsGgNqYlR/cDxErSPXB1ZukzkueA+/3NSuCv5kezJaYWsex7
dsCHx8tIojrEHRWvd5GOsmVGhRQJbMs8uz/WcuVuBTUsmq5gd83AHnZ0vwjYzSqn
pxEc4hT+cSvFC3QhujYrU4/2V5u1xAyJO4Z72AIJcYOspZZ5ekBnIB5N21QIXBGi
6zIkuOsApCI3oxqKzmSXYSdhKN24yCp+TaVgIHf0wZGox6xOI4CyMfQ4kamTdGF3
T4ZNbMTrdC+W0GXVzTvPKXUkVWEb25kbAuuCfA9/h1OKrTeGCDTnjQWFeE/LTQF9
VgAY7TipfeEH3ceNBvonS+dsgrm0rnBWDc2W7sPgIUT43XogXD+rSJFUtP9nNKu4
DtOuMf3AM2wRdkiyYpvE2RR1DPNhLlX7BO1Ntiu8pBilxOJ5LNjOEP00FbHvyr+U
dncc31h0QEs3qlMUgJxbvXKOmU9iUjuoRnqtNw2lvArilOthFDPGvAYFkKhJbtLJ
0NgksIAiP9QzokVzsydl3pOj0+UCuoikWi2MLGtASwIpHc/O2WFIw278pV3wShvg
NczrjyJ98S/QdweMrzy/6k6Fe2eqWF7V5GCEHlnlN0/SBqGuP8m5lF/AAmbTaAru
LTv5ZwmzVCT7fDW85NZdC9+aytvgWR/vaDt7J2nzdWT75Jb0wuGhIHcY5S2prk4h
NbHeZUTARlOzEuFae9oXYd7qCO1n9/ItzNd7yHIHDJhDtl0Gpe0WqitkEaIWxtP5
ayEbgbAR+z4sTROrIZY8mZERjKs7oxrnaQcAi0lpjVzJqywMgoInF5hdnz63y5VJ
TjfR54PDnXNE/BK2h+2paaExV9CkBBFSk3uE1dHwog+E4goE0JQlXfh+5DdHUMqn
YzbDbZR8GlW9WDd499UbNRxz96pIs1sB0IPPNFV1pg2n7UTCJqve+xdgT7tNRMTu
gENoragXq27NzAbIe+yJNVV6OioXqzciDLdLS0y4vajYG3ts+5bjtgkK5F7htTbN
9pmZ0rB6B1OyqsfcTY/WKjIo7cj5mgUBGVFtCH3PyoZlRfpqNPcGlw3AhQ8WikDk
hQuG/9ttATYXrwtKszKwFV9d70Gfb67SNsxBzYRrJ27aC7vBFwRXwi/Aferqhy6y
tN4QcOTBU0m+njUPLXHMqsgU5SdOCSyQV+aMT5BtbZn1coryAAAzruczxpF5X9jQ
P5H3TkSpzHwVdgfUXUJI4yYECkgcxxEDYxKtKxaS+BfK/Mhnfjjn6oVChX23n28i
CHz20f5KXUPdDjcsVeH4FQ+eV8+t3CTkzdAL7YnNNFu7zp6+SUwCTksNpM8BZhtQ
kUo8hoRbCT0cmvJQpCq8q2sXntCIug6apAZ1Ddcw1zkCDLcEKo/DhYsr9D+nthno
SZpjH1jQwEI6Z0iJ27zLtUE3J3XrQDEpMts4NbauTQqNnlRIe8ANzkjHQNKsDrzk
zlELh4bYMfuVzvznyxXiqWR2noToSdAFLFEIW6ew7a8KGiaYiKErXK5x753BOAb7
x1KPWrQRmkynnbjEdOmfHlxZdT4POuP8ACsrG3OUHReKF5o/au7lUnjYBxEtOMA0
2GzP4uMYy4MVHfX42/oKWBa1ObKE3J6fsN2QyoGrIEiTYkYtdE8bQi+T4L2kU0Oo
scQgkry5Rsub3EJWROAK94VzfjrU6paZyw7PmaShAUpa1ignXTHQYZ5d9+VybPZQ
rg0rg1/KMzRcEjp3ulqpVZgqy2h5kSHQjg/tiNo4fG/9UlRQ6lPQscY8Hz6EA8qP
Sngv6mEW1MQxJQf2ij+F/OyVESbWb2YX2csCr90//EuyZd0lwwNBrp9+ttop5AwW
axlbsz8sK5XR1YsS91WEA6vaXf6hI2Wi0c+fqpvHrcIWbUitwL2/IkpUl1z1fgRL
jLe2VhzAykNW+4ooTDctO2zoh4t6V1cEYglM90QLK9p8koSpmh/rXobT/t3SzEtr
HQJKQlXNv1D1lhqM1n+OOLan50Od/P0yzievCfxU/G8A2kGhRhSrw5PtSDbO+Tai
/EgIfGEHaAwNT02u12xql6w40Itmvg51lViTHl8iv1YyCY5Zu4f+DK6xljnDWiVo
ajzyRUBlFkoxqBuWpCSpT0S178T2aW/JjZ7qUao4BPhVOYM+ZMWDlmrwASOStQze
HKiT2apGnNQtJxiFA/0cTT/lKocEE4AATICOhLRsUiaO/+t/+BCruuPP1TgiJlBH
hcZfc35XaRmgydkbgLlLeOyUmrbgmndUeLhX+gzRxWoUkOeljYNdueFgi3J8hUU/
JJ2GiIjn8Q3jS+7Ei/Xro61i4tty5NKv6jIl7/axNVt8sPCBVkSTVEOsagT3QQEn
FySEjR2ifgqL+v1zptPIJKaLbCQGG7L8qB4Kp3e7kbBX7lCoCVrQvx2iMKMeup0P
ezAWnp66qLcCOMsYjqKTNJzGZJv0YUS8V9vBksoB5NMU0CEZPNKPd6ta1o8pSYPm
csWWKXuhnovQCoQ8xa3ZcEUVCLRl/1+ot77NGo0bnRcCdkS98PI7dAlOMKEacDJH
UM0OdZUar6HdJklaNFy/ua/UBXfoF2bej94Oa6OspDtAyG/oOWBptulqkLqa5qMW
FLxdW7MErTZBXaO05GopwaMsRNw4aVsP/+cuwLyMlIVFgZ7e8KmAjrBrfqyptoyu
cs7fl8vdChiX5rxsmtVSNZ+upkQnXaV0iWjpBpvp8tN6YAGjE7WB6R13y0dqcggO
WtoaqqEw7E82PSI+spS/mLUvIZzDH1ZtgUI5x55H2EYZuqiBUulgZDKAZJ2AWkpw
rIwAc6ouHt0w70L5FJIg8sIpGnK1yf4ebFAkYpafaIOhlSvXP3//MOI+PL9tu379
6oyiKVHXluXuEVUxsoCTYuDkQDCeoGSSVNGNDslwdtPaPlqyZMT7efCJ8IJ+OJtD
WSi2YyyUjlln/c5/FvpxOSsNJVNoUovSnoYDplRk2nntTMcnkwiw3ahlR8vAhx9v
neC9kgb+RoYmb/uCBQ5RnJQ2aFKKlOG9p1UAEZDr6N1Xmmqh3G0lwBxywmjWp9rf
4NZ+ZxC+S67rtB9/z/rRUxlsIpuT0UpF67vMqfTOD2OswWYtYOB2EDOcXNj6/h8H
yZK8qhmzufnbaTAmEbP5EJ0i5aGWLcrGIiA+rHhMwL8A+HW7AIugW4tJZDFt/3cl
Ie1mGsdkfoEImWp0BH2xR2Z7agftFrkJmkz8m83mqn0SUr705ULxc17Yyg9Lr8cL
AvlKhrmkCBCEFp8qOVGmqlP1wyNI0ijPME9T+4FsQ/vr5Axk9gGzEQ52ygmavs7G
+mA73SGHxgbgkXAhyms8IwKPXzV3A/8T82lqZpO/CXYqgOmO+cJLes9LWdGBVga7
MM4UpF8982HKJC3A5g3SNp3raPbdGtsGNyqbgyWm77Ha+GBn3P5TUaFQYvwsQGLS
R/zyshXMyUmFEHbyT0awWjgQHx3T8bXyq/AtnfwjA89Ub1FoI+Kpq0tjIkM+9rTo
1GK/zMSDGuKzF038Q8Vxdm2wFSHrqNzoDJcXJ7aPB2jD462ZTZgyWfUXjVon+q3D
QocC1BKdintxmBvR4iyEY6tso0aL07zpE5oaDCrpmCD/dCI99FmRTYGvTBLSCBk4
OJgaqaEarmjGf9oCYD+TZFX5WQcvRJ+D2kmfBubAArz2EDJHirkI+LIEWBDye8jm
TMxZI5oExsp/JuCvDpFYjbt0rlRhjUQiwdEE5Nbqf6Ln2ZxgZt9D4Px5rOfKS0x0
Nm1Tkis93WxD+U61UffDEY8nXaOCXhhJL4XBX/Qj1BW3P1rnSiAI7ENSV9g2sfzi
eD8AK+ygXdMwos83jMqbqOqzNnkHZpf606FPT16SRb2MCGZaYvj3x1MSzSHe2EVw
8oMyn9EDKYxrybuxxadXsd8TuMdsSRDWfXG4nQen88xZA8HLDnxwV4LYj2URNZfs
iQfUMmtVFcumbBiPbMdBQRqqTJfOZpRa7KXo97YaTLzl9AUv1K1aGnj0HprYtLYK
IwK9HKt8Qv5bKejN5eZXJSYeXpu3PKyhmAFEpXzF9vQx2CHfMy4W6RT6mWRx1dQa
puHDT61uL0/mcuFWbZaaRAQOKLE79JdLQtRCk6zeI10WEIoRTSs4yDEuCfstbhvK
kfn/fJUAa5avEo2QANiX3QjFQcNsDx6zMMXmIVr9Ry7niSy+TcmaBO/1Bwl2N26W
Wjx8HXlrrEqYvB0lAaeDBNrGxeYXYsxPHhfIqtEzM4nzJySTsGSWb6qXquGwVDwI
IjDVTHIHTKorpgl/BHGupjOBK3pQAAiO64qIkJHwscC/klPxAMARNyBl8cAMd+FO
IHR156Q0ag67Ll2Yw69CjMYZIGzxeuUmpMTNQmER3bxSOr+ro7eXvAn+AbQDM6kQ
+HOj9SzfyXnAQIaWkgXqMBGp2KscwNN1Rq6t0AJ2l3zCBb/Q2LBcCBbKGFYTQACE
ffTuIG0Mar3YSAKnGIvii18RJ/SSIIeuag8LnuSCdELbNaOnIHxMqwPU+xhIM8a+
29LD6WCmGaiOekemzyh7RCjAJRheA0vj2v89AS+grC9Ry/CBitDZD1ulgKwt+owI
AMundR3F3Q5nQjF4spG9wcGe8qQFTGGkEs4d1iO9wD4Vg4+/gY9o+DXgco8ZaphE
RKEDHdQhlfzwRZv1y/jscLsU7FddZA19qMeFP9w9ZcehkVgF8h7u+BC5UzNxzUww
P0gKrJDb7oYG88WVK1UVEXdrrs7+pVWcREwrezv1sM5Xrknhijme7grNPbGqZRma
r+FomtYN8mso3lk2wTSpe6icVDd9hpOKGObzEc67j9OaTZEBm9o2uy1WC0egR0gp
vVPnfRKEPuOe/Nse6JMmXaiAdaHbznMZVn9SbSX4E84QiUPbM6R9/mr6sT0JovqA
WmhI/M8WLUkcRJhAhzy4rBD21XFPlDrNdZySJ83P+3IFScisVOP8QD0Bb2C/B56C
GDdAq7hi9gSZSEptkTcnZjEslrGm/DAw8Ctj1/E2eTDV7/Il9tLFGDWymY6X3+2g
ymw/XqvW1p5jLUye82NHkzaet1gyQNiBZ6NmYa1fIzL3MSAfNGy8mMF4YMLS5Rdx
p+V64WALXy8aEtcilk/Qkj/WxtaLqhAOiE4J2cIRbbR8fHJLumOk6l6C9KKUG7K/
cWdBlTYgsW1L23E0RWr7CW6MLoolIPLHZKw1WaTPvNe9k5ceO1RK9hayBHzgDx7X
yDmSCEgCV+mdGy3Nn3dS/rGMvtKVhoyhO+DlIsDoLvPvFAM8JM1+HeyBDGOvQQAF
xYLYUUzwpH2iyHF7pAPVTx/ut2F3ghVk5+D3QCjk4NIom5T7ckD3gQpnZNPj9Lez
ArpoeTFONlNpZwMveTRpkgP3235zEGVjLm6gL6T3tvfJSVes4PhaJL0WaVz/xzdI
qM//oFjwsn7axRSRZuw1JGMDI5eyzUPy8GepVmTJxfRS85lyyHxNpLs1VKFCO2WD
XD74tM56Po2N82Eak7Z+vtQXx4sjuTbszrT+pLgtQGuupZh1hpXwy+BVpypRKz3Y
jwl3FWfnDKulldcbbJ0P0/pTYKIBSSX0+PIafhPpF0v+u5cQwWkBQTzJxvir4w3L
kjj7eGQla1voocxqc6IUhYS/jEyrYipWClnhDbEhhKOuPh4MNsGtAUUs9ndwn+vA
zvmjrIzTJnZFJTr5GREkhjng6NBIbsSNB6N5RKYAnB3+5XwKq5+rAlsZ5SRiNkbd
c/dfknpqNM6X2oN85qx/JvcYR9qHWFjrlB6IxKZJVpD9U5l0XnlKDxWt/MzvUkrY
1WGZoYB2InDKraT7O0lK7NSV5+cg7t8d69ugKojCCwwNjahc0oUBBvdaKGhu72+H
I2EtwJZgotT/gYSAJKv1aQg75/T+1t1ZwNxGmDloXIePtt+xbKkwOVpkoWuim5qn
tFc5xCe1Qg7KW/EepJwJeUfncAZBRuZ5JnRRKJsVXVSSk+c49EbgqYUn63h/wwR+
yDkLeegdDi+vD8hn8tH2vU/nc4ZyiUxi4XKCSpyYPliR3U9gxITQFehIvT8CmxUb
Z8DwE3+0cjcEW5m1hWy0zhRZKGxygh31dQzqn6+ok10uO3fBK6GHmVdl4RrwPFF5
MznYlKl8a3/Fau43fV3XAo4HTbUUOUGMh1uafwA6uqAhLva/r2ruODZkTsyN0u96
yowxo77ftBLuoufkPLlggq2flCl5bSqrjrWWGtfCTW5/IWKdgpLZ0nRsK5kII5UZ
vTK/iHpwWIi+ni7xyORXQfYRIWlw5MLkPConkgdzJCL1Qc2qhnOtgYUmI4vyp0Wd
2hd9ifyLpFEIAzfS80v1a82/DGC4+8v8TFAOy+DQR/g3eDCgM1+Cwn4WmLrknsyH
DJ8DcUqiS0dD2S0/8t78KPcBrhYdJABOOZSq9PDOhrP+vYdFIhI4DUhBqrc/47SD
mv34g/KgprG+SjPYhd0XyMcsh3iNnxpOnNsgNEtyF3esXjlb0Tqa9l5/cQjHxpy/
YZj6nUltG0uQMcODd9N+yCYjio2wvHRiBbMmIKtSGLg/zKn6Vr7eAmWKjIvCXQ+J
1hRmURGyQMt7cI0DB6PnIn65hhWGwNiBOXE0PIvhaiphSpoZdDCCcpzDL4zOAmi1
mvrxZqpWwfHUMDp07elzGRbgUj8dfhS+ipOZCu2Jd4M=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bL6vTctZ3HRit+0WvyauBhR4KduwWzMsFzFXX6hh9LfLOP4zomYSF4HkeCTRKdrj
lwvvfv/onz1nWwbaKuEzCbNcxWCi3NnaKRMCjC+yCrDOh93nYZmssGxLdDnM1SOc
kmnVFVnvVX6bPeiuMi9r0F4TSUd5BJc2KG25HfX+PJG4eOP0IhFjs+fce68KafTK
LQFlZ3njuo4rH8WqXrn/iS4GpprRSag0efRm1BmiqgE3hod3Wg5Am5B9lznmtgsg
g2KnGRY7W4+EJfYFnggIjdBvSQN90At1ZJYL523xBkZV5eP4K2wNkPS5lkT7aFC6
9EfN1R0jiqqzbJb2tEU4yw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5904 )
`pragma protect data_block
PcaIbXGhwwuFsAZghTorlj2X0NLlH5p2bdVYd+P+m8M5Eisrw8b4dN2QgJFhgKE6
5NGYHDigQQFsSQZKhsFK3Hl7/rI/5lRUb9utH23Vv6M2ICrPtnSGflTGopvKQRJO
yZKINCAubnkwdWqRnZX/BFJBwb6k8i86LMoVqnpjsL0lAkSVCrbNYz6pGuDzgUCn
jkdlabhiMs1GnqWXxxPYY7Tay4Tch3MPOf0xQJrxymdsuvxFQuSr6fov5QX/P61J
6wJKDFYwl9UxN3muypl/CpBeNg2oYkaPsAN93wsYy5g82h6l/OfpZGvih2q3b4QU
CC6PCI/lSbmUG/H+/7kSj1raUFzbtJxZsfpHwzaISODaHxGdhyNqW8And1eDrSr/
GMW6CR5S8l6jTPURY7IFsHrlCVTegAek7HW+ItfJLZcMu7pGpawJwitFNPNPgqHN
3mmx+R3sMIoKc75wqIP4OGUDoU37GP3lLXgPCA1oyw8jt0BvJLYoh5c1HRDplkdn
MFj3jB0MyUuwgykoxU+e1Mc5h9UliIVarliln2igk8/Mm1NwhA5v+L5uelypSrnS
Wk+gQJyfDL45Tj6C8X+Q1PMCqwjFmRYSAnve5Z9nKZ6yXlIl7tz5axHRS8pd2sxN
DMlJleyhUALr2BZX36D1RR6BJSdXUwI494QNxfiuJpGEG3mqvsJt6WMXwzx+ljHh
/zBdM39bP22VPncncwkk1TB6JbPMTdV25RWJM91twNyiBRnNgsIeIim1Nv/HOArc
EclKfMRsS4TQqWkUQ3ISLb+Ji127Wyo15mdBIreKLemUzL90xfpFWZhoZuSXA3e/
yqYOoKcpV6QckH5YqcFsEAOthHpO0emzcloTaTv0UDdB2mTw/I6D3dfJJBLROa0V
MS2qbbEe/oqFqY0vGCQxiDTqmivagq0pN/j09LUvWd54sDt99b/vpfaVSq+1WddD
ZiuZtbCcr19t89k2fe+raQUHBtuSAV1M7q2pw0Q+5aBazQTh2NHl9MHnvsVT6szm
zeBn8Ly5JuaquNp5r3mDciBFLYKCv/OFehr4SiLR4d5XM5HcrfKfjpvktyx0Xh/X
AYvM2VhCiLXV8OG6UUM0RPK2pwdLF0kGEI0J4ZiNkwLosT/N9qkhacN56/RvoUzS
mMotbbnJWwfbFg06jBxo/WuARfK+2YdF6hjDeE07Jc8MGhCAJ4hNz0Kwcdu2ObMo
qSG7JP2rk4kgzKu0suSnLLlXTdMhTerfknrKfF/0jccx0b3uDUeOcEJ42Ig2S9o0
j7KfaliJTLQF+GnDw4gUxyd3YNcASTbwgt8LP7RA/b6LiG3zA9o3DmKUJL/5KZ5s
OFB5NmhbT1IC2y5sPuRdQT6kDoxzewfGMyXgJMuWnRx7ATvEAgidwLOVkGsak+UC
BKyEYzfM4+kpHMb9LkuIFDYVapN990rR70rh7Lv2h4TBbnzSx2uqjehhRhwr25sR
twoHnAJ7mrSugcrkw54lE/Dk6CDMy/eCkxRLIjE9xO3maU/9uMcGTKiPwrJAdlii
2BBd9DaHf8GS9gtkS+tuDi7gtXioNwBKFRvN+2g0FeUpa4ZDYQ7Q4/MEIybsB+Cr
DzokNPJS8IDWQYHjBRKK+BYkXmOuOid05WVQqAHUti35BwX0iwZYSAr736nCGS/p
rePBGTNzNETPSdIwaPOjUNjkjT8CXo9xW2ADpoNRvW+eVNI2rsf7FS5gX7VaJ1Gi
xYHW41f48sPaoXuKrzgStOJ0rsedM9YRS1VE1NeLGanRR8azV1IZ6C7igJQ45Vrq
USPuIl4XliQDlspaSKbctfiL9VTJqPftbiSzk0cFzKm5vo3UHaWWbzjpFWCX48tl
Kd/m0E1omdr3A6I/Odg9lnkZxAPBtPE5LrIaj7PzGDB/t7SHIGvjwx8CqXjfL/uQ
ZEXSx37C4dXHFZHWCUa+c1pKvVScO3M8+ItTs2PosxWvCvBp+BaFDnHVHGbkIC7A
AmejqGYPBAGqhg8/gtimgJmqtzSoC8uliJU4QvmkMjSF+P9mnOuXC3P+CM+VIjLX
V4GIXhnWNN+Gt7B29a+qwB2/nU2Pwo22mcoVheHB5RGadQTqP6VTrfpKXVk4PLU7
lufr1NWKNCpmBOVOz+sk3hiXWLnzNg5X/D/mP2U0wk9Ebj41YJuiYZKQPcJTDYZs
83FIBnj9HU02Z+ijF2jGI0vcorqfSb4U/uW9X0w8IA48OT2h386hR+GHqZSnNceZ
cSC9sepfRMctfr8WQalrvZBvrNoqnK8JSpDJt8XHBrSqfezuZKVWr40LcSiMU1V0
oBtV4+6SNgzGAw63v22P8ynbjvqfLWKqE5CZgdsgRJ6h/Lt3wNN2DhOeqqNGpskE
m6qYHC9xmkRJiYeUfp5HrfVO/qtyuGLSXN9c9mJzsNTlT8vmqissw0EY2Hs9+PRN
/jttbU8cpPeVQKVQgi8A7dXBdrtw1zLwiLy1mmDcWMwqPSeh9Vxdfxv0/7Nd6fFc
h2btwxBwWYWSRofkIFOc1023YnhG9kZWySwP3ESfxWbgUzzANUaLurYgyfZ6ti/W
xE1z8h3kIrbQj0u9xoM3aLzLv4hoHrvuuulm6PYv0uIFz86a/bkX/5hCmhmzESEe
1CUW1DdS5sgG4MzQG4DH26+z/aEfHxDxUtw7o8u4sM0+Q+b8yMWGStV8E5j/4FfK
l17GdFwYB9vVJ2NTnhA9U2Q3cakKo9zSe/MFUeeJZ9yT33NSPr5mj6LLGX9iJyjQ
xXbNgxNFBIDBawqXB1xwUMlJuivM7R36i8AMLd/s59oXDMbmZCwdnc4VffczQmfg
8BKDty1v43M/B6OifmGI7wN68b4T60kxP4T+yf/UrkxH1ujPd0BLtjqFdqVWar/c
mZeUlXlE37ZCgwW03N7gZBbWNPgilKIfw2aNid+e1C6rc8TT5hP3/N1fx9fHern2
77j3/3Gz90JFCiueNzsELENqd3laiEZRi5B5PU3CMjDrehkZqJQL50FbQ9xqt7R5
5bD1LvHQWrFn6e2/by3hBdN5prvXku+CQDdcstuJMpIdEu20FJKuhtRswVmOUW4a
eUjFZgC8Q6GLeXfQJ4tbFt2/zUSxZHsWunzd7DUxjP68WtbIO/2jjt7Oeq/TWh3X
vaZjrJbCbLBnwoARZ7xcL2oDG6Xy6t7eNZsFX+RdH0vml/eLWoIKIFXyhCU/umx+
grUFZo1irxLLS0AkZ8bc97BX3ceyuuGLWVjUz2j1s4PNRoKmNmb0VLyyngfJwhhV
/ZZ8ogQi/81ThXKsf6Wb3mZ0SCGCg/FS6NWsq2oDN3RxkX0G84/9rNNJ/TJ4Puj0
aGXkhhs1DVg/unkCOLz/TUwS27OSzEgH5ISeYC6uu2wZbu6wjhxYYKSbuHnAUaWn
q7h1xZplPZbi5nadPQrj0ANNqnUY0SNoCV2dBlUts5qe9pf/3oPibZZvgviTgZjX
fzh3uqdi1qlRdKYPA9H9evhpeFGvYgsOnk5sgZC6gmnyFfKXGqOkkmCvgop9w957
rKYmyIOVzYJnSBt4x95POKS2olpnsUSZEi+SS5Am32vdMSxuNMeB8WhjAKTQI3Br
9nnWuv3zp65lvijaOGn+Ns9l1wo2e8d6ShaQn24A+MmqUtvTpgCriDfX0gLEnVan
1O/08UhizyCXyloLdFqX5gFakOXexrxPNcNY0PtcilpJO3b+8sifv5gVPsbTZ63S
6kAFoBjP7MXs9TeEedm8wi/M+6gWXlnvmjAj2JobiEybwSx9PH4TDEmWAkAiR/ng
n5P7x5WBoGVxXMWezWsQom8VgkJ1DsteeyHxRFwyMDsHehuU75/qk3qYXUxXclDx
lOG5Uk+FoURB6/Xsi7rOGFesylQT/O1nzo1g/C1vUZzqyHTXNK7jl7Wmt0Q45zkW
Krf5rXHfNQ20DkbfhqCGtl6WmJy6YMX8fbmaDAYkxjwj6T7wJhnQygPBT/8YfNHj
3jfvZ/Np1iIOw4DsYQ8XEzscbNl0FuFyJTGg5hMu4No9E4Pi/2xIeyCILq5gYhmn
Yp2vx82BumYsvd8NgkJIbaQdLYfpl5vxR3Gwvlll4f1ITuOLzTb7uv8hlSHHmPyB
ILupBrQgTHmz+ji3CD84N/9CmRofifxHdm2OoqJieYl8bE/Krxh0HTAC3tAGvHWq
YED6vS1VSdW8HTUYXFk4Aq7z+0ekpXUkhy0ZHPq5IFFPjUXEhzZ7pE7FQyyxee7B
sQSSjd1s8sGVvuyKvz4hQBw67X+zlRikdYGwj/qXJ/H59PLHFh4H4+Lhnau8CCAt
cYVxzn76hnKizzwK25qkyYFg8iy8O1NF6H1FFBSr35cp11VuZX4J0Eae/NIZCpzu
AOHO1lhqYkCj3I5YBdJZ14HXsRyNrGJ+kocoSTt25RPMnU7rOHcuaxlBNaohfG4Q
elAKGtj7bu3ewT9iAcFL0FHuU5sC7OB2Ki1UpFKdh3DB5XEEAx6qXglyEmB6zJlM
WTnYsSGf9JEqe5VQ+RDr7JlPuY/AsqogiVq/rwHTldTOvCpMpV1KyJ9cPHePJcTx
i7urMHM8awOHVcvpC2tpPwDUOK8BUzUFbGgbxc9qBA1wDLiG0gA1hV2wlYwLQEMi
0YgA9oGqb/A6cT1xbNn1rr4FcVNudckDrG+OcQ6ybK0UJRvCQTrhF1kJKpAxvdzb
jY5ex5OF06+LQi+r3yXPAomK58UgzbPcA29loBJ0v0/nQ9V+Q+XbxUyPVItpJnuK
KvngoUKW4yy4NukfBwoZDhbZ7jZiX540aPZF8DSRNQXytIjAgo6Cb7ji6bc3pNAa
Y6iaar4FVbI5iY6usZn30TgIqF7hmmkzunR2ZvPbbNjJu6/FcivCLpZi7YPION60
s6kqm8IUDMkTkuWhIIjLbCj3fEFpelIs7PcQPgKXwlFCTIWlLhnARje6Z2aYIiHE
hACNpMw+0mmha08lT+PHA8d5CRGJ1tpRYSHpuhIuB4SHWkdLDDuaESiTpGZT7lWa
n8GMO/xW71RKlTLgxlPkaIbv8SaQX3OeAaQhynTrcOea8CYKIcSQe4Q+rEdEqtMh
qQYcw0kXjeG3KgbNjuNvzfj8bfHYjZph6Uz/on5JX104sD2SN888VZhaQ/Lqzr3a
PvOqQFCdkFGj5y1NmflQ6Ei3L0x9sXO3Ia/MWyPtAj6p+DgGAE942j+p3KMWr1NC
KPR0/8E8boLkSbKoMUTg9qCNR9u3oV2PJ+Petac+EnIMFv5hxsBgqiz5HICG6cZY
c8sy+Y0lmRX/9JtNrW2SODM0V1E+78BwCusIFFA0FhNJ2DQ+0wMCR4J2dhh4ifUd
uGRCsvriGMqh1OalQbWtOp75fYi2qKfiAJigkhLRPCW3oKtDySXi1yjn6b9IVFcK
xSSDWQF55+C1Cx+KoCqaNZiqErn8H58vbNoBNQp39VzW5VDOBZsiDQmUIUFHJC44
57A55DGciKQfa7RRQI/5j+x5fD6IR+V7sbAqEaUhexIb6NWwzdLZwaWTlwFmxh+3
ccZBkfe8NQsTadVjCHAp6tA8EUHaVC/TVD9qDJr+lzsPRprWgwcVHINLpieeHNXb
nBxiflGeYVi2TByaXirKd5jyy4KuoFMp1AJzeKLHbrZ7jFPGDnNmSWAFOmBwozGY
F8Axqr0VX9CXhd22Li0crdM9SuZlGFnbu3r69CbpLfOtKTsBSpEeOOF7eGn4HZrf
6/EHOIFC4weMrEkE+tup4eGFyjzeg+1EwncC1GreSueL9io96Y04wepV2/d9Vcsm
yOTqIdSv8gWQPQm6Yaj24ntJ65/LT81whtlGY52a93uNxvLpStlfgmQwVYM2bUJu
SdEkkKu0z9BFpxpFTCfJ0+fytnLRScv++/bFlNG2OfNWKpnVSYqwcTzFzQOcS/Ob
sJPTE/KEVihIfCyqd1lORv7b8uFeuBVgMjCxoOPzQsNMheDR7mgDgYlybTQ8BWHu
G6j9BKQT1+kv4phES9vQyDQju8fjg2GeIphqUFAZRSAO5r4Ld76jFrAHLZwZ1tPM
9AJzbQRfNAkSDxtyIP7DiDa1z1G2JLKKV61Of7LlfaMjh1d4oi2enpqyN0zAqsji
bFrh1EN1l5d9YwV6xeaKIWeMZjfqK7CE9BDNopbEGJW0rkoIWvpcTzy6mWdptP7M
KANf79Mgp+leWotKXU1VVjcUedYlKUf702Di18IRuwmO2vDRc8WJwyB9W0o+aiqN
MFWO4758xAfZASWpGLZlkkanFH3tTfXU8T3xU1hSvAWHRSdI+Bo0rxWPHICAI4BP
4tantKT1uCzE0QDddn/7A7/E2HL9lM5Yh68xAxwguwFUEI88bKBbp49Ep7mAhHQ3
9Zmp0xxCgyfxfDiDtPv718xANGd4STsjbV/KVCzZN6uYbIDYwjlRSagC1vE4N3PN
2JZ7GJfRichDM+saD/t57N2L0BYmU5j8GxzZ3CdsGTpyJzbmtK8iqAmtnkpGPq+f
Om4ZCfvvL5Vy8ozR8OhKipakJ8gQBK7g+Re3TBRdh16lX2Liq2EspiLYuB33IYrv
OXUB8QnJ5yl9w28NoueUFLHNxnuW7FnsepAS+T8hwXKLqJ2Qv2kxN1z2wZ5z6Jbg
+utm8OpAy3JIwEAtHcFOGcWi2g5Pt+Xiw2oFTWBrIbHKljDQ6nETaGApy6UynDT2
Hs/AqBOC+YJYshHw017E+66y+I44EgrCDvxkravk5k/NuJSTthmeZ4CeQI0MNZzz
ZC9Ku4AbvIM06cDJu3yDtxkmX9JK4VvSAnV7tkkREO+xk5bYHVQcDqrHt07KPEyp
UwHI/lnLHwT1+4Io+8NC5MEVpiRy1BNQrCX41QdCnLnnxhwIVbenLjv5OKjQmcrL
QB6JFEigWUZ3Nc802MWvkspgRNmk+SDKijiKQ5DOQ/+kP4WRu2n+WdWq7QAIREAO
J/zV8GNdcYl9XJseDyXuRIzRqnYqD46QyQG5M7OTMaGBg/l7sC7+kOCVc5RVyJZ7
SU5BUhxCECKq/E6+ztZpq4zreST8iVqtr4Zde6+D4FknqF8Vm1anqNnb0QbwKNWl
s5uKDoIfRnLioJZzMF6Ptds7K7YMYaYVlFhlSIlBQq73k9qDe+7IJNVFtYagm8Su
ZvvOpDeSVpWz5V4sgI3IIoeuzdFPQrXqenmGCxCplT9KhQfN4nlxzX+zG5yquT+1
BqQQ9U+/4jFRZ/vwbYHLPj7zDAW2zSgpBsd4Vq6PRv5r2MnLG3ut5cx7pYrUTsy6
0tLXFoxCNHFcts8lBy3EltuH7JU6cvN1QDMEmRfz3TdmH1+m1X9WldSiUa65FAQL
uViYLHx5EpuG2TPgHq/qE+qvMvgi7OkEA9kUu19ei/5FmolHx6OX/KGxLIVEsAtF
3FAqbBA9mRwBl+JLByU8qXF2ozq2lMizjZCtBSYui/yLv4fihPRMkKYM5luTRaGr
DWCrltXLfqN3qBSdyyITY5LDQzPo4IZhPbRQYRNN3g/xfuAZ0+TQWR2KHYXb8/L8
ynL5Kqk9WzqrrDoxJEryhdfOLOAWysbd/C5tyG9zjdwnF2qsKMQz6fMxBZZqDXG1
FawrzczOf3BXRQ8k1jR/V9sl42+ikZhouQWnZP7S3yJk2mqRch3ppToAgpD8LIcm
Ie1HJwW5gBLF6X0nznCFZqpk1FV79DH3WwNRnxPEBld7Q23g4220VnemUwmBZfdq
vKC3nScdX6Sg7Tjnda4OtTej/Viw48RKruL1+LOfdVumedWLy1EfoUleM2my31z1
/MrjvzWTi/DZoW0qkCN3n2hWCw/mIbAuPr5yUoyaHrzo0AwXN4LbYmrDCHjvKF0d
mqVtU2Y/pBSjk7gAakyPI8f+WAyYtpiaBiF0YBWYa1iS26WzOjU1FLeQJY0CFCQk
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
c9r1fhnknvy9NHkVktk0NmkSTqv5CCo0eK8Tv5aeznky/Y7vyds3hr6WQaf44H1z
ubW6jPZaTgImXZG20ARWdRehGgLVZFj7TPvOBu3c01ZpHFXeSDTE2p4412xpbsEc
nE1mZQhjZX8t9bosGCDNF1ZYZ3/WwB8UAgaOZEbMML2Jma8/8XuolSUB1pPOe5Sj
vXH8uvmZzrTX/kxX+ToSAxGrO9PD08nN264Xv0sE+ElF7EVtDle4Mz3c5USI+2vM
7IfJYvk6Yub474LgeZNC/gUofABFfdQMNZtaXe9QZ3Ze0WEOIyy1wdSTEyMk7Ssw
L3CTyUUbWGpzvz91NBzZNQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7648 )
`pragma protect data_block
YPM1H7hEcD3Wt6YC+4dIxsW97EGBOClBJzebDiBAzUAgUqcx7iULll5aVkiAqHjP
ZWmrwSDYTTjc+0N0VyjCeyf9aQ/IBauuIEWK+kbQtmsJ7kcqOOm5K+JB9zJU8itU
iyo2VJQr2pHWVApt+ikUE5xC9+MzguQm5WTEannCYD3uKwX+8ivlohJiOT3KxpGq
yo1JNQFRDDTfAe7Sim2C6oo7SdBS2wO9gILthK7Aa6dcIiKizsBrjP57S6JlKWld
ObWKs+S7i+bzjHPJJw0YmCoR/14rPsmoA4vp0Z2Sb7gRyV1XKNkI+6+uWnKEkC2d
SVnfhWDH7Ya2rUr91sPRDXI8PR9azMnnwKO0aNUu5/iZORDVCI16UD6vv4IwXzcY
l/BvmijTvENHGPgK+3GCRsBFlEGiJrsKlFVncyv3XJ7xmSx0q1LvYqG3a5ujFnv8
htO7qiXA45DV0Bz+wClWIvBytPWmhIFblp8fYzx7EGpt/xCsCp/4PNbN8DXg/niU
g7as0r1oOgT2WSPu6nL6wJPIhb9qrJ3bCXHsCv5UC6B2/DWvBpawF+n5rcQagaEv
ZMrnDqxvp/Pq4A800e7MTX4ozf9V7OZCiFptxx0OkyC8NCIophnDKA98tJ+yu4L/
mSLXj6LXs+ulHBJkjeIJk79nQJ+EBu3B1yhvFKYBCYpUzr3ceLkXgn4AOLhrsNC0
WW8/YGazpkYRCytI/QwgPxxi5EbOnD/h4dRVx4/KSRQq6oBpJ7iFQ2hNJ6uxS7qd
EEGUIrE9wWt1wXqsooEnQgmBHe+iyPVslaUPxcrW8xZ9e0aKeE2XxMFJ0prPRHjg
Kdc/4xoMfuNeODMLCjvUytyJNMWXU5ITvWILADpJU/esBMIRKYp/weuj9fmll6zX
4x9GFSWwzC5dQSxRLbbnMZGor5ACXTzV2iBv+SuM0J8l2FYDu6ggvn7aYzVOFOgw
a50ZhoGYMQebuhasaWnzbFkrJjXphAR1eJnnYk+0LVKtJFpfVOQIhw7AYMO4d0ko
Xse0zby8g0rqtEuC8St8SAxCE3u9w8PiJ/vtNnXkzpmbDfe26ulX6JfvsnVggQME
8X03B4KlyC9TOwU0y/PINMd5HzKLXb8+EicIIyOf0Q3tmjbfneElmswvPqklqea0
e7eHw1z1hXi77HDoO2beBQj8vhADnmAmiNYSuuCQRfo4sWvfr8wFvDVDgxaJxyVd
xi4NzZJzXruNqhdDIfMyATlR6sYCwzd3nSznju0cwKDuPA3CYEehgXvjYhvliUYN
Vr1ftSYHAQwIWDQKcOMteff83jjrfSiorZDzxCWj+LTImHY/RU1pxC/o15AOgUnj
FGCxaj+cRXxy/RV95rwJcOPHD4v5SJXUs3kIgA8rOUnL/PbbcwpBXP3kZA/onalR
9pJtXDgLO8oU1RQLyk/j/o1YeqbO2akgPEcVdl8hES/8X4asq9/Y/HiTV09pZalQ
aSGPb4Zdzq7kfeespdphLlNJ5Uuvqpv6mF99OzYKdlCn6FsQX5dXTZP2JLKDTAto
tRuhgBp6L09JS2QBYjoh3qn95seuoFDVB1EmWLUzLkmBY4hsEFi3qBo/wDk/CcCT
WLFP+r3x4gdon120DlqduQrUbgzemS9VL4W8mbH0DjW02C3OHGn1MLwvMufFksdM
bsMjk7weucAP+pfus7ENZFPUqpGH6w5JNk7aRjRBWR5TLdNpiR8mJOk/OhdCZrQz
eDxfMZiVNHbmHlwQ8u8xoQnblLpZxkJWWQdXtNwolxfH1rBaLWCXYwICZ6KyA+Sh
T6XQguLQFmi6ymrbifE5pJw7Zzrz8JXx7EudqzhtsTdDlNy0P/VtN3OHqk0oGqKc
2vhb+NgKodAg2Z96zstycb93K/zYI6wPk84kb/czU6Z3qlP95xQjrID2m358N45A
Yjr9XXetPDcCEcprGKxFBs/6BBs09oCp9nmdwq23+VmLtGMummaskpTfd1CxEj1J
azq3tALH5QjYunXlDfrXqf8dNSC2vS0wg117+D7SOpuN3Y9K6PvU05Qo3HuZyauG
XzTWYVWkF6OrpjxA9NBMxg1qgbGFFIjycphb4LSAftmhiunPKz1/dFViP7APGnzz
qS4YglBBTZb+8F+FJhnRYv5NjpMoys5wXlMMBlYCr0lIGx/2TZ8hhl62I/1hs/Sp
cP5xOaZ7Xjvp+BBIDNG9F/g0dcKL2zwS5ZgtQUep79P4cgnQ2vo4Sjxk4xueiqL+
l0QVzB3fdXKf2ghSYnPG72mc29ri6BDK+4d0ZmFUMlLdKBuiiCT3XtF5GRO+16eJ
dk2ZcQLUCeo7PvMscs0e4yDIfvzY7hKBAHZkpWB/G4Jqe/Yc4iPwa7N4K/Gdo2rJ
qriAI6hR1gkCo6312H6Rtx0lqnUi7r+mhQExZYdrMkp5u7t6HZkGtW3SMD0CxdVx
gJ07ob9FfmvjDZIKmd7SgIb+1JGyCijw+prEGMYEfZAOBSyPrAMGhDwFHX6bNRv8
JwLEuUxo9ntPdTPR4zoQfQQHvAyE9bQ3p0R5BTKbaaFW+T9+RRA51xmXx+n+/Iu7
ka0WkcO9y9bjInr8DhBZEZRqZsG7JmRF5ar4WcOZXg4N1XHNxUz1MEKk1/xPSGsP
7Af2BZ72RozzMtIo6ZX10WcDTgjUsrj9q9oCUqHe7SdIHQK5i7zkniuCaAOrQrFC
o8PsnSBDxPfKEnUZs+m2KJszptXpttt88gJIgX9T+cu9oe1aoMCVM8byBjb3inIH
w/yZwU50SrITbvi3cRgePAxfBqRjwXzbfVDZQHwOEV01Pw9wBVezM2iMmKXMAJlv
QDZKEonlvX0iZcbqqsgIEn9DTYigxRlxZRpcDNbWaVwp33Y4kq8wG9pQ8HZOxm86
dJnX9l/g73lQBcpU7mjGaTPe87lKQghevGQcdG303kmysUtMd1Q+wnBcMShALySx
AUNzCiVqB5HziOpZkk0foKSTcPVny4fj2OIxdXYG3XZWkztzBOorW3yw9E5kO+3V
WpjldJw5lb1hHei7MQV7bG82QjnjrPaBQQ3/Bq+yqsYk5a2K9lCyymeptM6UP0M1
qJAmTVwuO5OY4dP70JNSatXIZNCmKHanICKzMCI/LuMaCkRSsZoqXZWY3wbLzCxw
6NHdBRe87o9WkiO/liNm9dY6MX8BwMjsrlGDHQsYT5tpze6YZ6yuVnzM4IPXb1Ma
eIdlnUYxfaRI2KNSHNUDT2rks6HOcf62yWT5vOQBkLNFqL2zi1ijSYQ3JyIFfihQ
l9Op7Hku3woeHKaI2zbDy7KG+ruSd2lb2ofZUPClhakhLWre/C7L7mjBEZiKWoEF
dnWBkVQQ/9NMIXFHDCdUbHwuYGLWjvA94Z1Lht9zV8r4ZnmZXPr7MIV5PTreNM2C
QjTCsPQECeyvPjU1ehwrqYZOqHjXNr24bDOXH1935ygSm77LNfkXIpmgHTGWEFvF
RyHFsKjM4ml7zQL10LbTD+YcCcY6Keyxgw88DsDHqioWLl5Jh8/5qaO7zy2eLuVu
x+5Mcwy0mDm+NrF5CCI9ih4wzTQYoqrXRk1bw5STak7aNiOUGGxefhATXH1I+t7g
3ePn9cCwlRef5qUAh7jTHA7F5btgi5cJhUvbLZyu+f2LLqeLjjKW5VKC0znJRdDV
RfSqC4oB/I61qJkuUFjCbj2pQVVlLIpEEBhn56SD96+Qepb4QeXA629u3LdSJkG7
mqgJkpRwMRrTwimdppNH+mXMmd6sPxFKuTCF1KOo4q7RzmFmFMKiPmZ26fUVFw3L
TJ3OHjUYUKSbVBCb+IYHD/6yfKjwZLPoPAnlw0DwmOJdlU6w5XVTL0iosnA3UC23
IJ1BoIYPKY3JHnRQ1hJGSerZO20whCVQEXR/y7+z9MrqMeHHOaHZEHERA+pOcoxK
651Yz60qQruTdZVOdjSLoB/56Rc8GkJbIfW2L4DECNq1OVyK03f95IqE0X/w5en4
Tzwh+vhkKGvTIRtLqJAX18lYNqwWKd/ER104yk2GcwZD6BoDArYlOu/mc5Ll7HnP
Jg+uAvYeU9BQUAKQqpDsaZaBIn8u+gSWSYoEftAzm/23najMKJM+N/Ed/TB0zKs1
nJBSzOtWmMG4Gdm1FtmsQdTW6Pgx2I20mXTJONRHCRLcMP6MQtGFdrakX14vwlpG
SWLZPmcdXG2tO+PccucXUgnLvoWK7SV4UHePkz9SnyVRDbIFR9mmFiGH+O3gzLnz
oCKE46bNrjRt7rx0Lc/4qCVWNQElrx+31fnZdbNihmA6Q5CCV8NJjDE7j/tHgWIR
V1UlFMGPpajHFbTWN6qhHITD3gT9g4I8AbRT6Aqm5Rc7wDum3OgOsakAtm+OO6ku
QxcfUNE96wOPv/GDh2QWCqxcvGHYvTqqvi+KIEEKUInoJeXVaOLnzBpg73u/xau5
U7Kx8KoPbHu+tOprCQzcYiN6SRzBA6siXgWEvBGIKN4rj4OUzTxXAjDhaPPd4iWn
BSbDkNk05xMXLqngmo7lVdoOLaIybiNsDn0RZWFSsz914BdLgoI1FBfqJH42yFBT
u++N1ivDT///rP19VOxjDOHL+YXnmyo76a31NPeT42aN/5QD+HZsKBTIyGdvEUI0
4OJ7PnZOjun8VIG6A/pzh/vhlIauj00ulwX8DVlHiRplC5yNZl0HR+j2abvhV0wx
9oSW/F0uFhDZ9O97LaN1e8UTOD6lOLInNyY0VOn7ZXKeOBBAvYn+rIHui/Qp5KoJ
IVfv16a03W1KS0Iiv5kLA7JqWY3gKNkAvEoLHQTYPwFMDnOPXta9aYGoMOlG0J+8
VuSU/+mfwUyekuLNUB9LX9hVlX/Gp8rYHgPna970DWweyx7gRGMrbBjPn7bHReHa
f4UW7cyswJ4T7PHd9BsaQhkCkHLMwVQV0oz1IuS/3s8m8exR7+uG2CEw5BdDwPP+
wEpK0DIvnN+vJrM3unLUwJW8vQdLhn6zGR3k959G15jphfnWTKvCvFnujQISW1jD
6H2oDGAsLho0iFv1BHGSYLps0qQpiliI8ZsB3kqdywiETFqTiHhplBmlzW/k2I+r
icok6rzvlnumnXf8FJRGVe5EMdGLVMYOQC7Zv5ZM/yqIsyXaqFPeJ5lvvm+liREx
Di2dSQQPM0Iz2FJqmtEN8SeL/N/0PC7yWMbZB4zc6MhA4BV2WwaXbzRWXk8ow4Dw
9n8WMIiHzwbOlipOlobEWg0C5X1OXGuvQ2FMg7W78+06C53kTkm/csnVa84nJJWD
jq+Ns2CRBrgCHN/MtuJ+hid37UZ4j+UY8im95bDHYdGJdRVu2Al6bjHSS92FYPc9
exjevUYk9PDmU2nqDTuijKsnkkMO8t+E2eID5mwdGbP1UQUKowfmHo6qO81YJ9/m
S+oChsbkXv6HAedwYzzDXyabgOEyZyaRXmNsVUL54QH+YURFkfHXBz3rQWXPZN7O
TitVzWVZaOiNNoX3uyKG5C7oJ4a/XDxEdCS7ahkfnVlmFtq2pqQb86zZt024dNVq
oNQTszrHtf2aigIE/uKTMYcE9MIhn4Rj/1YavgPaGuasd7AIwVcwdzgvBDscPfFL
g7E1D4SAor3FVtZ43pwaFFSi8cJuzziP5laTP2IoAWV59bILgwIelOTH4vzjx05c
wVyYgX8ki5dKrlECcFgGLL4RPndsYBbQ5ljdnPFh23pbOaxUvOgHxSCPSke2iMos
VhivRTqsgTP0lqtIbbBb1eTs/RNa7jFJeaBbLsIe2vJ7yx7kk4bdwNKLc5r13RWF
Y1KedtBrfnqtrnxRiUMY2Jk4XWRQ3uQYMjbJGmOL4EbG7D3EcocIpGSK9uy3XLC3
ZkOFyXZTJdbvE4nEH8Nc2zktFxhoAwBFTl/zXBpA3ddG0lUwYr1OF6/DiWe4sNgq
nf1iBhZc0+jH5Db+tBLyYyFvGmwkqkj6HJ6YlSGZ2sOK9MqdLSibdxswiNvbPtUf
ePg7OdQZJ1Amu1wmjD5TtqG5LfrajbAGTys/ZV57LZFB2L2HP9buABzKD72qYjGy
Vw5IFAFQExdrvhqu1qSaKb0WOW1sOenU6VCw/DmXljmxlNF7HossG6bQhDO4RuBY
FNpXjTQ7z3pCBbhkHebxaoLBUzXIoemRynCm/g/tV3hTBIjmmCMxRym06noVHuir
OVKoWSRhXFzVMusFQKfmSIYE2FNykSWKgw4iurJFGA4okMuBwJZLsKIVX0iwk8hd
3xPm99vCmyE3ixPG6ZOzkRt3tMssZ0f9cTAgjDRHXzKJd3MHyB5E/zk4KNALNmLy
8U8bcsBFP/j0GlJQhyhK69Jg9ujJ26CwyAlDtNsghg9TLrw0Wc0UTtNpGfA5Tfhq
FulsPNNquoRS5t+yYWqn2NBc1E21GjDwVCdGkzcHj0kqOT+LNr/Uc3xi1nhj8VLh
B3kmxjnUXVFztX90+NvdaZIdN9/c6KOGA8ki4d5/DoEpYU4ATBpdsusAPjo03sLf
hKyzmRWsOqewseuJ3s+od59CvZA4vPdqAHkGAs/e62+rgbFRN3cWTzcx2pOZOQ2v
9DI7Ybv10+XQG+XOgaqML7fhxJN6hzwpx9lRFURk+IORMycto7yj2RQpABzyO7Bv
HrDhAqOt40whltgKe3wxwfzO9+HhlRFTNzvaaW9U9pkHoPZ6G+5n5ZJMLS1tcpj6
dtxs1udsgtEOVJ47XxkbqC6Q0iBuZU2waSRypeNC248m4FvgPQ7dQrB2/iBnorMB
IHYm6u+mhb7VDC0YkO6DLvn6F0F5owwdfv66xkw54iIIPK8bGLx7MP8lwJ0BiSyz
uoCvzD5CPCEH9d3NBFmo6iMU+vhX/dQFt84uDAtEBrwEqjMMh/F52c9j1ND0rWcr
2Tjkf2v+/XGyHIs4ir9ofZiqbRovVze9/M+8xByoWZAOLR+SGIAUogqEn1dLeJYs
fvE1HH7MvpMYrnTQZQxdRj0QjDnAUjQ6CGZgRCSVkt0RWlL+FlaPE0JAwdLFo04t
kTyW8+RYH/EbkgH5mQFzG081HfiUKE+W5Srvef4O4rrykOp2Qx6szGNGMxKFIx6A
CN1l+xmJgQYiACjponAet6dfAWfPOC5C01j0RKafLiuAV4BjWYCQZD56GPzIv7mH
w6q+kh3zAxOl5FP+7YnXrAOBVHkvOwgXXfn5uIy7GS3eXyC84gPBVCbnDuw7U8Xj
8oLSMiWP8AlHTaHWYQzG+FsqZA1rEzWVCxibvyJYkMW2n1eOg3ngCec2KcQrq5PM
djtnxEt5ilYPdKk4I1C/bWR94JcNifYpj4Wg4TGHwEA6aOblqu0U6vTR5M7cO87v
MFuoYrw5SbzLeBfYyAVCyIOsVG2aaPvtpicQy8VK4GT11dF0+LwbVu5Fh72H2m5f
Q9XFNWEv/TBrXeswb8zR2j9qCpni5ThtIIbwilhQZwcgaTHWl1xor9YwRy/4Rpuy
rQ26nGU2tO2uAZ9aM4LTd/P80WD3l8toeNt5Ce8qAL/eqKwPyqQ62fii6Nv+6VT6
/fexzfiu5OMAuuUp1pW+3W6voJxVoAycJHvR9DpWum+u2/l8wcMkL3oDNgPgahLM
uDAjXY/L6zYMwoGK/ZrlRYLhIPx1eEFuRaYVJYWnLBq9zGC3vvt/dmkuKKX9c2I6
NIIbnpvDXTU+sOUq2nmIgtNaWj6IhA1rPBXoc/MyQ0sGNb7cdJ+bgTWmHFHU1zQ1
YZypC4iKKuSVDeSd5AWNtSFw/kW/EnycR7T1DFTktwbhD+yVAY/1SaOwH5I/htyx
PL6xozkdYKMKdGRoxHoP8FPZyFtLQID/KbHM3ZSGXFQ0MZpgfNFzTL+kPbMyDlod
uQophG6btEgQZyDGiSVabkjf/2aoGFH9woILxaY6j162sq5MgfNwhYEteajHMR6d
EXDBIfBxkfqjSzZxvhJ41gsmej8pTYKBUg7BM7LAEu++AScDp/aFLc5QzF7uybV/
0bGSeqzbP++UoWP7cahaeIxL2gHQKh6f0lT0/VvwcukEEQ69l94FCRVvkhmabHkS
HBx5HdM3OQpm7R1usjRfk0d0k9Wy9A/5FZ3le7gEBe8pSH+Tfi58j6HCKepEzCYx
mzE1cPyuHUi3pIkNbLby20VPq5J3aqYrbviV5AwevaKhm2jQVIgug7PzrpRRYahl
NUxfgGztISPIllb2PLwPNsLCwUIN30vXFwnll66LyAMiPA1m+C/HNlu30WuMUXHF
KnIfqmsNKYj3yScR3xR5Td2qu/4amRmoYvxQBkbtw2Sh0m+oewF0N9cP0nFw5hVj
/Fe9wx4hJBVWEVeCAQxnCR8vVY/XkWQSHv8rU4pFMZwlmwhyT2VskY0n6LDVW4oN
5IBJp+Q5bCLRvKG83gvW9YcddiZelcibjD1JaLnZ2dljK1zzcQxoc6xvC0GenSrr
Gn7Rjl+p7s8LDBQmsy28Qo27Q+RUWhXPWSIN5OWNsObznoVEdTy47QIFLrYmLOoM
puCNdB6D13mqZXYrmGXdt1uTHUvPG2gLtNPMJbkP4/9K1GN1f1k+/zPKaRhz3CYw
oVvDxudj4OH7K7Y8/sW8EqkE88oW3jDiGwGyRtp3DUyX2A+NZukBwjyNj4OxBYIR
FWTrC4uojA/fmE53U5TLcle8ernJ14SI86NP3682PWacvP48ijbN/umo7bPKv6Gg
bJUNA2EXLkP9Kc1qQbyyDIWV1eI91t1NfPjCDz7QEuw4CH7oajmzGVb29VS7YEa5
zZx/amdVsXvcTsRMquTKQHK+MZPXGGu/DGvUskUlOJZ4UD3OGHwD+G/mi5r17Jdu
/t8D2gi7qcqpz9a0a6ks3BEEbGKC0aGZQiC6thgVY8o6L3I6gWDu2H+OFsKnhJmi
EQAdwLujw4G6fEhrd73t+7OZD6EIWrAIlpX+xrsKF4CeZvrj47UphWUStVyQGWY/
YfHYL1untpVAb008RG79Zi84GToY8nZrP3HuAuuBUv9qoifpR9Mdx2/OypMzbauC
uDvsSG+Lv79tjPV8uBWSX9mHYBu7NOlSEtCj6c5ltReSDY8MihWJ+QsQttQjiSqj
7nyfrmrl9NqeDu1fpNcP6sBdoUWK6AmVPn367M1Z5YavmiUeC+Rp7qENlLErCDj2
JVS3acHOwANthlGJHP/yvTMikvdQSMDnUhctpF00yCAc3qeLybyYgMtJzDaXXxtP
8lVoI1dBXFVuJUCjhKbSxl9LuyKiG9LAJ1gtzZNH70jhzHAJVWb5eJ86XV7ro83Z
FLcQZ2MVUo52Z6lMlNfyMhnAH2dybqWcevdWt15i1ieNluVhOSteHCU0vNHYAFJY
jNcxJ4OB3aCZakACxv89Ra774q1paSW6XAGfsChMWqNjD8YUOgpa29WBVVrkdkXO
vqdxM4ZB3F1KzL/uFvqCIT7e2f5VTzCiM2r3aUiAAwaCv8urPYg0InHRSccdlOlh
fPR+Ra8CucSGYEHJX1V94+8w/LDinqhFBauJQs2jkwF0nIRhFwDkL+lnytLNkpdh
IA+ljTnU4ZoGEoTk2dOmb+E6uu7w5Q5Ky1N0dSZ2ahQdZAgcCDD2gjaP6xxRq/jD
LT8bTuK2t8IIqc8PTo1gIRwRhe9UtZh8cte8jLt0jwdTHdX9SRlSvHqaZ0qnFRFW
sVDjU3LdkMrjAvRoe6y39wT3dLpuI/WfUSHJaTW9lRjwVLDrAnCjdOjL0783VFIS
J8KniWqHJvzBXOvt2gUsXML/KDb555G4HLhPR58UB54PSDbY0OgePVegWfResute
bTQADhi0BNo/j7XTfG9Cz3k3me6BVkJ2BQ3Vwh6jIE84pmVVuum4QTAPaAn5TleI
SDQNR/0O6K09ym66GkHbYOx/HlzPuX9qmED9w4LElRi1JqZswvsI6c4l2nohw9/J
EswwfGOhLxoNXvCys0qbWb5oYiTIl+NTCQ4AQoxEzJ0++8LGnaTkoanW4UtbTRIc
kFZ6tBIUk2tpk/Sb9OoR4p8RIy8ExD75Od2LBBBIMiwOpoSyXnS9NdEKvPP6binM
gsaBlnE0HGIoj5QDXjnMk84ngMkiKoBBujBaqzsP1mv1XPlH8UrIjN4WrO9o9Uqc
/tjBve5Wzf78CLukjk/YikgeaFUrSqDrtHbgpPukkPtEEiowmMn81KY7CuKDdbqq
307VzRytiGxJHtSJ51SUyOluEEuz/riXa7hb+U8x1iJAcokSLmMQMn9grpCOetbQ
aEHbazcYNBrEgfAm/ZRI3w==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Kn2goq7OOhezBONGm+4ggGqo9583/VlaxlNhFwco0ZPRLkHqJFwnJ9neuM6RpsPX
L21K7rAdThQVq/QLaIrRcZ0Gv+dfMLx/KNCCjUOcqKsJXmpVqSjoZaBECnHzfmYL
VZeX8MFah1SQIDZdYRg/pQw7n2XlMcrmAKsWVTm3BNrufdFsOkgmqYfC97uyspkk
xZ4DJ5jWY/LxIArB/W3hJfbKcWmFPZgttRGqUVtxxTU2VsM1XNzujnCqHqci/VbP
cBKAnRiDCbZzBbojNYhuwNxD1YibS0C6E57URQFFBFdUNtUHZuKJvK2TIMPn9hP/
QN+e3L40PWlcjVA06+EICw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5632 )
`pragma protect data_block
fNGZNR1xXsjSfOWrt18gu0Ok8qQ/PCSVR3+PGss/WKuIvkMuRyhROeIUYdQbXTWk
EI4ZEdU556ULB5JZmPEQX2hkUOiv99yQ92CVH2hGg4jWirYEM8AiVJw+1I3OZMI1
4qHiQk6RoZ9wDZLGwEaqMmCzw8rRXSR4FId2OFm0XJGwQfRwSzjuNGYfn9VX/dMr
ZL1um5UIyW1e8tPGpObWp2W3NkFgEy6ZfjryqcWs9MfADN+K/+vutyIVpHdcSHot
Gg9qdyn1iE8fkpu04l8xaAUv9iNWoJgYK7C/xtkm7QVwUYi+Z5mDga/T1r84EpBx
uzX/VEygQcPmU/XOM0sQDcH+yUl9N+gwu5zHa/JZeF7or9a+V8Z1y1TI7ZWGuo+n
tl4NEXLYIFt+KbYaTnCnSNzROvk/vuLeJ9WtFjz+GuAeXXBbMHKeMPo3ZaXCQFGp
hxiHRL74JCmN4hJeDwghaRyPFqVfnmnesHOmRy4LlHN7Po4staCj5YPVvumQXjc2
T++hIdYmXwNAqN+SrAAeNle4jNLCoiV4YPCDVYLEea5NbMyC/SzV5E4qsB0pXxwJ
p4L9VmeY+i60Fe/rvtaRWjCXn4W5wUJuLCYi9MkMthk5RXIh6Vk9IuftEuTAMNz9
PGbQOEyNq6snJln45zeWLw3rfTb9QSHLi1V1QAeiLopOvACmRDHMwPTonC8dXsOB
SWLNeD8UVLO8ezH8He7xW3emW3ydXInDzzf1c7TnkQK1vJtHRPdfgyTwSEvximo8
fn7037jnQMp+E8gbZNQoo2BbeP3mDRxxWnyes1JcXTTE/rBgNf62Yzw4bHMHJzEW
8zG5mTt+/0hI4jOxX5vqlepgwBjnlJn5+ilitG5syUubhwHKAj7N3m0RVfXekaTc
VNn2BKYfd5TaQavbkryYteb3xtI3n5KFQaDlGC0uhuUUEB7bsnhR1AG273ytohb5
MiK24FlQMwaCtwAVfVC89phwPSCoBsrb8G/53DsNOls+pX+1fHGSPjJK8k4E4CwI
69rMyEdWSmLwO+us/XVtABGhjpaBMmxh7mgaCvpJzgABFYH55/TrJdqDhBqYzuZs
ahuCjuvE1C6d7RA4M/n3F0XRihF59jRMVfdw/lKErf/cFcyDJqT9STMT1WxPW7Lb
K7HPAAx7KXtYMe4aPrgyD3AG73zpwspuK3a87hLvhUf7Kr9UEirJJKD1WGBylbvj
IDEMb4kzb6U48x8aUtwevPpau7V/6cnsqH/M7uGHAaHQzuxW3zXf5ci4JFxG5sDi
akYFTE/X6h0HyZtuFEC0hcbCfTrjBopMAkVTTkGP+SxZV9zCh3pixUyZapluYol1
Ri3M3X0RAVj+s6hZnkkblik4Ya3+Ch8cQJ8MdnJN/EJcZso0DJbgLlSyIP7t43ER
RtNQg31WIR61c06ZY7EjyrIxhnUD0DGQfnT1VmRRaBCGrCb45eKBzaxv2pJuK+8M
DNisbWvqxnP+kZrtWWgUi/qCI0jo3rvIOkzqbWXAsROVOItgcoBjPlwwUwgIJj2F
wwArUbJkfF5VPjOtXx3EmPifa5dtfhm9+bFug/lnF7Shpgd3i3ARlVKP3CbUBnh2
kio0bony7Jf5VKfggXq5661K74x3iJomXj9Ouka86iLA3D2yU96rIicgNrDDGE+q
l6o/mHki6fGUxdOBXx7Xn7jZH1h9BE+IPPLryJM3PIkUqAfB++tsH8FTeKCoDNrb
oeYYDO+DcVkti5jVZU5oq+Uw3vvWGLSjjGMq51autoRi21e5R7Ubah6P02KlUi2n
fEXHDx36xsYJWFCXFM2EJcUdgRktEgiJfYqrpsr/yvfnK6JowGPwMbJbdt7HPwnQ
z3DMxxGJA8nfErBlHTbSvlRP9QUD9seKP16zXWcF3SvCcVMohDa0V3plyZ1w7Kvn
XzTS4M1vUPVM7GgveMXKWddkUT3yvoa/LeKIFYRSZQTLwEx7Trh61A6QgFeNYB8X
Vo67C70BiyssJw2W2KQ0Kai9p1ta/wFZ0wmXj3vBDYsdOOYKs0u7sokpw0g8wQJI
xXhLOd/rNAXMXz5MvPkPNIr5cmMkAMgmDablri8K2zxhcIG06bSy8TMzq8cGKtXO
VMF7CQADvz9TZjw1NnqP1MRiGLyiJ9/zGXOxizyFseW82LUK9bckWeCcxGjA4sRm
U9/SwzjF8XBkgjt7IAb2X7LflBqMA2u0w10niwgCbT0GFEYb4qnqlgoz0k3wtUZo
NdJDpFTtHZ2pSaiC09h2q5H54T4hiXQyGyTBfKGYvlDt/+/pnE4he9y/nK0zJbnT
tC+Cu9A6kQtLU8WP7Z5eaL71xyZSsfBjE7ylD1tFw7bIWbw+t5aLN3kWxzlscfXb
aXCKBboWNYg5strmq6s6TDK+dDCGB6j/N2YDhuxGaWwl/hVA6b+S6XsIoO4OurJz
UO3CYPXcEXAKo16nBqoTI49VNsINAuj2aVBVhAWBY0RbAUBMB1BLvTwevt9y9Xp7
8S+KSyf+o/WfEiPiSBrjyi5evvTSSW8lY640p5Opa8VQHlS43+PT1K2+Ki1YJ4XW
Dopt5x4+rspzLauQawOQj+jnrnr46sonViC2vlBCM9cjliDd5wby3g7dgHq+c5Lv
HE/6OmwPAyw+gLvNpks0az01dAyvUE7HUtwpAChRDX2iGGvgOM8aDx624CYjCJS9
qq2Qx5sXgxj+hFGKrtrqbvCETil35zPhOW4y4MLAZnpWrJiRTxYGoYhrlUs32mMo
lmkrfVervaViDELrMSa661MFCDQQT4z9eVwS6ZIUX/6U61wDxw9zU6OJ+xBqWWHC
4R6dZrNngb1yVWOhkoJZZpZMdJvDMAMvg+8D+keiTHkljGn9wNDEnnjz1L5Q4acQ
hUS2h4yYVsk0+jncNVNdmnFBrC67cU4bXzoMZec7WA2mWk5o+Wh+KqDxVGs/2bad
Bth6yZcQWYj96ruo63vb1/cJemqZSXnGnxCjNsRzKjrIxB1QPRGcfVYStuN74qj5
UlCFeIpLlsdm7JpJkI+Nb0lqZnJhBMKQFjel6E//+8OpyusjW8SicCj1VuYdjaYX
WYVfVcV40RgrpLFOiimJmuxD+W3B/MX4zN+w7hixhlClvT6ok7pSlf2zDh1atXe6
mjJkJvjcyML1C07w4eb6yJQekMWkjBXASy2wdLjgDsFKY4/3SI9iet9s8aYejwTD
KHA5akRQmlM3idRgijDccycEOxTzx5PRwnnsmhl6BmpzMmcDvLu1Crav4/na0MgO
GEMJLPciLyFp3Bb12bY6E2J3ts5s8wEVB6MrlTG6od75EeDOBD646if2WymOGfQz
ykw4aGySnCoiuDUsZVGCd+w4ghW8jvs05YxT2G9aX9atRtjSHG9+netG9bsNQ021
TCIosrgtE8goeMtNUxhwM5i5R33W/LGxeX8SDVrgrz0pq5KXt+bmfy6vx0rZKVE8
dBdnhkHDBEjw8ra2JxEeLqaZ4vCOCZyUd0ZUWd17hGXtBjN6yn8zzmF8oylcYTKT
5+7CclyZUsvg/aSiRbmZ3uHXsgqUR0e+05f6Wbbhx9QRZk/rMdjLcfsIUnBOnY/t
3MnA5MtYBG0uHB4bLP/OiaXtcSXgQpJUb2g4h6gmN/2eashDTJtX9ZZ+jbUTUH/H
Uf9EudjYQy1G1fBI5CQQBVpuO8W68JmTeAxzjvclpXsT7DBE6+y8Cvqg1Mlgi7mp
hR0QjucZuz7ZqPIRRJh7EhBBG1A676LN01Pi7omohtpxFAvVyP7f60god5Ayzyta
s45HRAkWP2UbiqLuhgHbqevZU6m9ntqHNWehrV1G4axzdSt3D29gNU6rWx9Oa3pe
ILxMysWUZNB8GgAjJebn6KTws+joZ3e6c5apYPdatfxlbBRuNaQrmJVaQiauYNRw
bGjW+oLLQeikdv8DGxSnfffLryVbryn0fIwHJHZgAADqLzZy/IyTHbYP2t4fj0rz
LJBqi+mA4rDtg/eaiBwbI00/Wf3R/2Dx/LFAIKBua+a2xvtS+OsFBNwx8rtJkYxh
rGRgRg2Kz+vooAsJUQYabg3KMy6iL02/PrHnjjC32HSWBehshtbs4yhba7bGKgHr
8sVDRPj6S2aJAQpD8DyUlvQDcuHavUyv8+7Sl3RQoslJt9iYwcro/XUrzOjzEHAR
L1QqELWU4K+JINi/4NZD71FfGzGc9JhtNGjNH/nH5eRqHs70GxRGq0CPaq9neyMM
8HF6mP7Xzek/5+HVDBsyvzjEf22kptts+zZs+gtA2oNN5hOmHW/TiKNmeesfTklt
gaDrU/gDNJt+VweWjs21yIYRwTAYvoXAw2IZLQa+DHEopAjDPjPhPigQaNBzZNdO
DBU44n888kPu5/pCqnmPI146rMWj1u+LUxO+qntXJZr7JnIwB3VPTE8qq1kyhTGd
K9MYYvTbCEMUTkW62cpj5TuswXqzhMpgHRzZH21yp9ck2mYmwW9kW697iyx1QCQ/
/uXQa68CvAfoZOsGcqDNd3JXH5kgQmQdNYwO72BhxbtJMUfREoPCAw7rOdwBtMMc
dwzDoOYxSadt2cdp8I+yRRdUyPehC0Rqna0fNWEuWQdfGzhq7KltXD0QNBcsTvId
PKNNSG3Vd/JnQiK8Jz0OZ5s3s57qpsAFL9IC9ZIaE6vVgiF7SMSQWqSXsUhACOpW
v72szrdUUmYmxqAnm+4dlMjtX3Znf4Ui9o4AEvFHSkro4rMHgrmk8aOQEGUfGCQL
ceNi8pX7j5OZdzI5KkDCIn4z/UCuqLZ895y0o+U10pl8VnOiwUTQvrrCSsKg3G54
gw88OfGGQ+THzF1lMgyJS8J8ZYfeoXtUu50YKE1vtmZVwFEuBJ1jtcv0QnOYFjae
7fMy5xusCB0xXa/oCLQpvuDX4/LbTc0m8iuGlWqkVBlnWYyX0LDctpyvPDVlC0up
rs1qxHKaIOTqiqjHJRa5j5HXhKdpKT8mqM+EbyLNHwsXroWD3areBHftPIk6+f2i
qThyij7Qwd0VvGTDCJCppiJ4MKhMCmVlwSpGbUniAbxVRT3eAYxQEzyOtJHWGGbs
m7hBcrE+LMPrJQWVL26eJQeNCe1oiKG2xPcLk02oVTsKVQ9E76Xt7AYbIyUNbloy
bGp2HcZ9eSPM6mQ5GW6i3HlDeONeXEbBpg/a2fq9XkD/1s9vyofhXyLdHHaDxr4w
c2x+zmzIUzpUEi8cIR8Uf0X7kTdjucuNmVSJvGnDgqK6cM2GjzpGKJWFlcV+BoyB
QFrj/wI4I4TOyNGnU2oYiWDxjLmOHjcddHc55v/U6lPnMLwiODTd9WUXgRrhmQcN
pqJHwAB1WTeXJAQF9MyUTnfBW8Q6dMx0VT3Li+Hq/ORXzuxgedbouVAkBH6pDZId
G727gKSPuwYlSx6GAsUcE/aDRE335KDthgV3oeCI5u+kveq3SteLDdv0xgVOfZJl
SFz52jmMG1N6iyFz/pT915awKJFIK/U92rBbWjuJAR4w3IiV2Eh3EoHPCrVkILmF
WGw4VSg3bP3YtqbwqyTDWWof2nZDjAkJ6lNWRWAd9+MPaFLq9mtRYEWq5s8ULsA1
+LHwt20YNoeg1aGpEPLuwPwSEAaC6cBqb7i8/2r/lsmNnOR2FZSH2lF1Fgn5JEsl
8eEDKrcpFu6WyoRgXuwVmoCc5KkTgdjDPBnEZV0BXemF2MKOBBqfMsjfjdzB4dB1
AvWznScrfVTEJyrg8ixyFHRYBgM2wLGJWT1cKJbakjpheksBgWi7ZaL7YIfmz0B6
CGbrgspeVg447+WhNundHcBgSZiTGxADKsixBbdzhazQQchPzrNDfg/ROtLVR8cn
b6vbH2h4+Lkxfy2TkcYv2XZFcIbBHGFvLbtYEiUfB2yayueeNGnRNyTIjmNELW+6
iFDNVkezG7GTCadb84dG1vJeW3YzVfomdBGBoUZHa8m3OljKWXIe/yYTC+y5r3gm
nVKxWozIHOwd10f1DWENVdBTEZSxwJ3Vmz+jBDo+7RtSsL+BpwtY1boFt/NxZr0u
F+FxQIQr9BqGRDWtwDDL8481Uqf66l/uT08TGOcIdiYLrdExH908LTjmOWJN6rd0
HCADI40WQReaCxhNBmCV7hWnej96RvG/nrtijccMzaML1FuUC3oVykfEuzWBC8tB
jDCopvEd/Al6nVfIE4WAhitfbDCpT/V2PQhORNTjzzpE2NaZqbpahK3+zTlGh/OD
Wfs4AjqVdwak6sf/CGSW2QBMTCuvSXSdGVkJ9pjXLZJouDx0eVg0RWota5tgly6O
rRC7sLPFWFdG4FLh7yjC1BU6ZwhGs7tWcCI4K2jF2bQoVQwwQZwBBCry4HsB/+hy
wD+rY6FoKFPAWb3V0+s2m0ia0a0kehIM05/7I2Kh8Lk0Y9l5YvvYv/q7hZoMyOAR
2RbWCzpa8DJwnqeHfGOG7hiRMiOKS/7VhaqmDhM6RhuRPFW1FeQGqDCtlIQdD8J6
e8+CJ0iGTvgn42Sv/h9hQgFr2aL4Pev/syKpPZZDplW3a0ikpgyR2vH8mxZCbedU
uQX0Drbn8dYDe84Wxf8QrPuI6DlODF7eMQLbkSYJlrhN62G5GIwXWZ9p3BH27S82
sTIXEPJhTLp16Lgi4/lleo0cwAhJesQ3WYM5XOCGT4k5PwEYelsUEpbighVDbquA
aAJ/NqtBPX1y8Wlmm2Mg5nC7b4hUJ5U4QqEjy3kZwv4KahKyiH7nOYMcGGAFq1kf
57VZPnU57GrQu4kOe1yv/9LEqedtUCmRl65BgOZqqhGLgKXPRwvNBT0buxzpllEa
16ORzqFzew/vDMXAVozRs+sET8olUesMIEBDvl4vUuC8AbQhfT7/FCcYw29EqFez
2kzo82cdx4YFGrg8hxdnx4hJUWkQ0IRWgs5BIrknKVsUr4EGRFyZGPzjO/5EgYim
d8XO57ssX3bXWd/N7q48A4tZxxUSKwPiwWY+0IB1iv6WrLnHeDyQjKLbPPrvbeC/
tmxE6gNdQtY16t5hWZ2Gr5ECt1FpTW3o24zwZF/QnTOTYmXgi+87daUqKxKxbizH
+16uydTQeVN0ZsBOsFKiCa3aZHVwgIOo9jZJ7g28ODoiwGHTOJiPsdUYAsfUPlUv
V/QEhC7WjXPQzTUiNrlvRPKxQky4ZKJy/4sXriePkRYm4fb518VRDTEgxSj5R5cm
G1yXfIMwfsHMbj4HbO9fltA/8pAV+1UkVNA3UVKFomuaf6Bv8iGoe2jR8WwlIBYr
I+LxOt9v65f03F+1jAb4SwVlB6dzzDmN/VpuPbzj8UBUJVQoHOFUgXWm9VEu+OFh
eWRSf1VubPL0R3S9SC4fvFXX6Wsl4pnOqxyv2ghN6Eut76FokMD9YHEnxV1IlrYE
wwV2qE6Yf73qLlJsugpZfaRRSpY34hvxIHeB1EUi9yoWdYV4e2WrFoiZIByBwr1C
oGs+ojAvlnM+gl3U5XIXp9nsaOmaMf8QJbCUM+o7KiGWuC3CS8wGmQEL0kJS39Jj
7NG93GaMhMVjACxVthSiwg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
MZmWpvuqeQcoHUVhaske8IwpwAb+eqCDKLIjcWmyRpiJy+tHY2L0efAPFcB5ocZb
glvtOBw6OJZylAqAI0wYcdwxmSYKaR6E4+nOIxGRPV23vSrMPrqpuiBD4EWA6xrR
ibI5Nl4tVVXSzgsh4F5LecExgAOCAcaoeBwfDbHmQlLifzBZm3YCcXZP2QOESyXz
8pxme9mFoEvHSJ5bCaAmad8B5tH3BPsT+HVw4K9IjnTRboeJ7HZFZChPKdpAu6t2
HKZsdd7YAtDzI9klODlSRG2lT90DyvweWTEpVkaOLtO/wLzY8WrBnDigxJJyc+LB
K0nuvaRPG7wn/c6av+trIA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4928 )
`pragma protect data_block
rNRn5DmlU8pMdBQJPeDi7pbX6vMHFifv4A4safAjciUOTpUXob2bIE3DFAO68wBD
6nmFVdtfPI/xHL7gcYxLaYDOi53cTXqnW5OcBe1W99cJbROn9E1NykOBuYGD15Q7
WAKkVOfBiHmG3TSgXA5ejqTSNY8gScdvnpOSvMKdjoiUQO22lTpppTJLl/yNxT0d
OnOibpXd3X8JITA5/fY/4f6CG6rW/6Qe17+SyEVRZtrRj1jQkukWL6loqfSJyz7g
2ozvn2Ugf8+hdUad9uA4bu2u5KwUpzDeYBYEWjIeL3AGg+/yy/AEeSPkxmbx/DAa
/fUJZa75xLslHrpGZ5bhSFHJfKLrrdqIPQsEZm4q8VoZABqdLAzIKdziXEzHMqbk
Ois/x8yjpNcAdIoKCykaqeQiSk5TiiGHBzOORV5tvcFPOMisia83P83n8u53CfTM
/PVb3IMBj5y8fmGJk62ObdXHpvs3bQXv4y8YC3Dv4o4D6sIaxSahe2oGjg5FsFO9
TTTFmelpq6lmu1VNikut+u674OGBHqCZsgYXpqXqXOnSXzcsaftPB9IuWwa3I5b9
F/WfyMw46MoUFqKYTRMabTpAArFSPASm5f773KGM2JzemNSjjfhlPbhDotCGiCyx
EhQAsYJ4kwKaH59KubYW8eL/SIDwFMEvXn29vqkmGkZOg6LfnBgWJLWoyL12FZSr
Am8Z2MNW5cRS5JQBq5HyZ/552P9IP+gP312t6e2F12GB96rvl6aSbS7W9L4QLVCo
vLfE8wUMl+9MhCIeLwrYaERiUrZq0ey3UrooobHmLXWVYEfQFXgiXSrOlm1uMJYz
S+9rt5I+WSPfDxM4wV578oM2ZVs+leN4Z7WCpM3xZJ2h9dLbS/kS2XfLWORmmaIY
MNRrd2rhqM2ul4ft7nTWJ008FUJHsLh+zlRlkOWeFO+xcw3ksI8/tSDWRm6kKEt0
Pvs7yVAg66r/3GFVOfQyv3zfeHf6Sy++Y4dRBmNOVKcayVLq3S50dZ6KoIlXdlIn
7fdHVa9mEqByHZdmc1Cs/lraTmFY3D4c3P0t8ZM/bTSNMHtbvvXFAh3M6GpfvH/1
mTM2vjn4D7E/2px7NYlt1SQXvljhEHX2Yo6yhBvlclo2wSO6YmXE6biECzAeyS0O
l4SNEFLQ8sgZynKQkcVHVHZmcCpH3X0sNa/LcY6/rQGAoLtVQyTx5ZmBQeltkglp
gOIahVzIN4Q0nplz3LZ7lsxjLyvYb5CbmLR1G+2mURFh6RhoQvn5nqnHuuCizD2N
dWNK4V0IvykABNtLbWMuhzW3d/5d2x3/qvzr+I3hBcg59okNcmo+lXnLlZ/rkgvW
q7fhVLrw7Oay8Tol6XR1mkoYRKvb+aC4fBAYrViC8HmKDhoWzwcCX9wU3y9hH2fk
tKD+HWGh7WsDrEq8k4XjD5v7vodPjjngS8VqPK5fAgA0c9F2KXij//RS61E8dh0h
mRbcKvVIbfn3ExAZbjBZbfEZ+4hqKTG7RA/mLSuETxwj2ht3AvygkDFTS3SfXKT4
CVXHCpEm0A5n66FwHEH/Ct6F0KCtdLwANnBd5FA6Sq7UQ7/R5V6CqUYgW9MV+OZi
mSZvPvPrM8G33xl21yVTolbncqoix50HnQxiHlo5DxTI7KEv6kkFj0np8B+9ccML
2X+noTXlHxA8zanr0nf3vVocZmz85E73Q0l0Xcp1j28m0T75RFUM+6bcsfziCKeA
8MrtOZxRdNYZ4bERg+S8FujNSafk+FZQG0X5LO+q0YtY1LJHy27MQgwcf7U+lG3+
NFk3OsFY0/ZqqPHFETLNR7KVqvyX50xfE80U+m3c5Arkx9K7ICoIbkFKV2quL8tT
IoFo12oJC7FF4BPw2MQi+IcqUYL4z1Alp/n2xtA0Rm5rg430m5D3PFE82IiTyOHl
vT8dlyKpl/Z+Ns7/h7X4IHVhT6lQpqSFqh6aAclhM1ycc8y1jrBYkzFm8CKfmksv
cq4FUfyzemsN5uXoq4cA3uCEaywEhp8rbFjsTINQXKoNSQuR3xBHFuQMxtz/cxGZ
M/iRIKzY3vnYPOMNhFzR3V64F9e8kFHXl6a5MeSD72EBkn6R3WKv4O9PjjfvRndf
Kxn6pIQJ9kR05dydKTMSVdoaf+5sXH5kr/Rw2gyAadk3fp5kWpPNV0Pt8wj5/eCJ
Qnh+2N/ZnV2GH69LvoPkKtkXvVf7nDxSot1LnYDlZ5Zkzy9Zue53ydOeOUTqk1ys
2yzwJKFhVl7gzJr9nvYYOKtvmnp3JB4SR2VFnxeHnfD7H1ZnrwiEcgdFU7IFNbbw
m1t4QjgytL5uQNoaJXdQeFAIAYzZv5U2EgfsCo1xZpEU7j1dntl8wGBule3xSC1J
NuEYEVKVLs5sjLlfsbCR89doFwEiFZ7Imm4RCO8vDUlkJSN9Apozu0v+hYHafZrO
X+p4Ilbt0IYiqG6Lfmy3eaj0+NULyahx2G+eu0ZYRdH88u9dDiYl3aGm9rXHHHGV
UVtizi5Fvk3GKtqLAdTMHH+9TMgqbZd+bXofZFWFxG0gnJ48MvtXgaMbMU/bXeoG
tVeH6BTeqaapo2rQTfi3wlNjKtaKcyOLqoNduQkhDscO33EmFR9h+v/edWbW5qwk
sZu0KbRG7/A/P04Rc2+njSnTOikUt0/JpH/862RO7SP0R2NxB2XIWATfo0ARg7st
ZpBpJZA1wf8ZMvxu9Q9LfPTqSPNkywNSqT5uhTLasPwS9ZBgmpYkzINPfuaScNvb
ZuskikOHclFtyn9pDTKsuZZtM4ri/xWf2inMxCmZf2T8W4I4xdRKtOu22/k/rs+R
SPBaez9ijCf84FskxMSvBZfuRYoAHg8INGuWP4gxHwOAs8aULLUac4tpdZjZRLQP
GFiNcMtctg5CvNqfZA63eXoLxgypIBS60Mxdu9SjsIWaPvbb9DKjjRuQddns6Q5Q
kqzdwnwU/N4B1jnpKM+j1m7tlrAS3Tlom1h+kCEFMLGjr7rr/077b2V38TsaNIbj
n8N+stRNbm7qH4OX8/Xx/8rRs2Lj+4sZ6eWwPT1jqjuvSp2AUrmuhDTkDmb9ZnPP
XbQoOLkfx0gpDu+ett79X+Lwx0KMqX9mku55Vbdxygvh9CdhwiIGHxihdXo9mBxj
nwWhC+kB3Lq4ONE5GTDP5WqVsHiA79h+FqnVdvBPhl4lfNvXsL82udUStCgo56dC
AG3BxXXTWEFBPTGKSzxv3AWlLJ8Ha62/WWkW57DNVV0/ygiYOjlZjYD1JtY02KuY
El7Mp+qv0RkMYg9UXQ8y0WN+Kwf7Fbx4CnPgDGOX6qpFpIT5mSRf6IR7untQVOwe
I0ZWoXuLT/ZZG2NYXf8s86/7Sz6qZlpWMMd9gN3IyEbZYdEySG1XuPAxguwjhqM0
7yLnVZzEEuc6LgPiiXcV9Z1Uz6t+SK6/BBjZlaIpOADpm77W3+q0eb+GGJKWF54F
Vxhu3cMuQNAWgHoKs1SVZuWwYLtBgGHHbtito+9DMqSth3bVTmShnEScpKpweZHF
Ibl3zOLwjWxJkuaJhUS5+zbSWXa+Hpog9fxz/bhl0yozRdLUy4zTbYR6UxjQnH+r
cmMM/A0UoOekr+VykQonoGJ+iylG79wdkMftnGyNEkemD0hWEeTMv6jT+nsDoAaI
NvIyKXWKd4NBLaW3xqLqpvTe8z29F5/u0E+fcxEGwVzJRbnQI6lt5eFdoWaLI+Rx
NKd+4wqlOxuLDfIE5ksYiav+2TgtO0tv5YWHH3EsynoS/t/8GxyPy0gCsTrq+u1I
pn3yWUY/Ff2TUxt6u/iPtIUXgJgEXMZQ4B71Iw7HpLMSjbtzw/qth9ipaLMGBMgG
fH0x2BdQaJD0UWy/YZLBJglO6Hb/TRBcZtfs0/RtdFQrlUaLCIJmcXMi0Yulh+Ro
xtGlFUXgmsigUUGtKT35phbysBSFpxi8y405CBBGGbKWHHE3OeVlpwdbABI60gIl
03zl3RbEXy0TdE1BZucKfAp7rv7cEwD/mw+JoG04BhoL2zYQSxeAxxbz5xjYXVo+
zug/crlZ+w9olpHDSnY/MaGPU4vFtokMaCf0qsXyFOWS2ti2XJgMcIOJMdOf9o63
YFWYmAeKiEXBtakXdM7GHzQwFDdcR8c2BcSPZi8Gu/Mnq6vjmseh6IjkhKBiLvSa
dN2F9zWqbNH4ebjmDdwC1y/vwCFpLqp1I0q0X32LVdLkAQ/ksxmFxP9cX5OY/J1O
tLvew33p9HE7Q2uTcYYIEtosSGhG16VIafVoPFbXE5n7ApP20RZ8DNz1yeOnDvcr
P323G9kp4JZNrVhsXZpwckd92rUkkAWdPYBq1rRePMPFvA5ihljNxP7Hl3G+GK0t
jVygDjeE69jbuajmL3Wx3WByM7HRKCTfmI10J9S134YgMpjhFVMAI7OKXYXZf49Z
iW9rrdED6MJNRmBVnOlBWyfzXjwtKADu3lICsIME5aLX1bMG+hgL78I+vxbmhfAO
BYO4pZdvGB4HeyJ6Yp223ra6jMsgjdkPiJWCReVeAQEyzwhavfffeeOdpXFn8Cd6
us8EpLkuGRyEPVkdFgPYMKWMsj9phjkRo0eUgw8vCvKPHXgb8+BuQs+hq6wyuapS
cDjMRGBZJx5KGlvkB080jBzGqFvVk/b3a6dOwF9of5x44mF3IkPDR2T73YnwMjJG
eOt04gtQ8L8xFXRFPwaN+H3KfxiGEDB5ndKAC4HlXS+btYdoejoEhJ6JqVu0YMbv
D92vwvBrxZ4zJPRcc88v5xsKLKmfgwhie89p9oY96MDYk37Iy+bvJLjoOOpchkzK
zipg/O6o/NfvF1g23kJX7VOFgWDRg/Xf2UiKRdMEFxSgY9yZnApIQtRfZTXfZhPO
9oCZMU9IZbacx1JkJ+5o7zEDqwTZEZI+NEJGlDJsc5Hv9AZUvQlxV1JA11DYcSEC
HpruJgirJlW10kQ3syicxGEwmTrdRXBPCRag4lAvnaonRjP81ZjQt9RcpxhpNRNv
6gcdig+OOsn81lsuqBRS7Xvlg+Dql7s+nh19M6R8j52VFcwV2Il2+4TxuQ/T9e1K
NIwZMxEVVOcXIWPQmsFJYeiXYksvaLjcDgX8Anpjow+R81wrM7aG8gZm8iVgYlad
I5U3diS22uvD3yA9YmYfBW0TLyKrHpBClttGgrDlTBu3f/i0215O8eq5FFeyqjvl
64ooVOYh+PdylAC6F9g/MpaWnXfueNduOIpK03udnJ9nvymYKqfqNOWafWFxMuyK
FwvDJa0pUTi2AX29GooGUvRbGnP+/Pknm0tmtFwxUNouFTstn+7bZgpfwnDPMVaC
sYX5NC4kWRdx+KcU5m1YgZv37oOHEdOGP2R44O1SN/eMrEB3gs5zNRy8k1jjaIOq
43UDe8oY7TOnYzLrclvzQBK2EYiVUfkpaepo00kYhs/fIvVf/s8OFi1HmDYdv9YG
WG3ovw0UjaTq00wca1nyozXVyl3qX6z1dU0/h3dIS4SpvhmBmMU5kwatMw62LU5u
lPwn0NaepwHH9epDysF6c4AmP7xgKcl6mPQuPjIxE0bOUOc1Adr/vzXM+AuyHqaG
prs93odF7q0AQ/9q0nphFSg7NDjO6fYpl7iutTVPmW1U2SWzFw84AI2c9vcq3mny
6HjC0epXIZGiddnu97SwjtYkEIakk22VmvMDC5sxwQczN3d5DE5niek6pbtFi7Ht
uxlBzVvOIO8ysrdnp77wl4Lw6Hsl42PEGuLxj7o3finHvNN2bbks/mt9eJWZEK0m
bg/VMR83ts70Ytm0W9wWdlPxRY68KU+4bUdcytbT1SKs5SglFp1tB20jOGSQaYm/
7LAsP6CGTfO8USe5FJtNP1ysPKzEyWhp9HT7fmPuKBr9V8dxBvzebDsrZoNowQp0
jYiBuXSa1aDLNVqgOJQREBLXEUml2VCRGgK0yVP1L/W/a1rxdwT7RRCUkJZx8PhD
cZsEnmEcG0Q5GfPcEj7Pd6QGgkO1ugvI2lJOjymoKhZ4rwqGuIWLHaFjp55Kv3e9
5zMcmGuWHN0UPLJE5d67wxijmiVmDj3ToC2DsDE8jtZ/ErRonEmmigeON+iFJy0+
snw3OkxCdOuaPaKzQKOmhV5rMMNoH6dOQzr/+uEBKgqK200pcw+PlRUU5puwawMn
sxEBa2B3VAYddTRYsARt60htUHIMBHJW19oxj/JywZYiHWAN6z6fxn+TCWqxODH3
jQAH+1q6U3jh2riQav+fwaPlPZp66woHJuYPkqEe9q70CHHOdjDAgT1L3quFyMs2
WBPI0EjxRq4mTqaFL+Dd0jcK+CduPI8mbKAhl/H9N27lbmGkUtj7OWVSlPYfgSgk
6vhb3wweo8ZhMwXRWoqhai8lP3Z7AOJzo4CHukyutEanYU15iqpiWnP/g0g6fC1l
OsqROFcWvi7r9ypbdeRDnKdCR1ZHXoJuhe4cEBteMh5Zyl5XRoq7lSY6uSYzivN1
oBhDXIdpZiZQuJukMsliVmK/Rj1UJfjsOmwULGJqNbaErwvQFQg3IazYtsSDiF9V
uP6gj8BL6dYXx+Eg48LzuVA2/W98572H79Cg3FigI7g=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
n6XN+sX4MVIOC81Ig0cd9lDaYnafuG5TS78c40kxOaEnt9jQjZck2oPD8MC9sWYY
M6zzXg34NKic0pASqIZ11Qaj+b6fQb4ftnLEMDytzzHZFEahyHTp66TCQLqfJjVd
lR5boecLjFhNQSY8nNJVgpDq0U8ekVExIiSwg+0bD7UmxnlV4uwfiqxGRMDYVG/4
YNw7Nbnand/zTbLMZGU4WjBYwM69SJppJt0AC+koG9762W26423tMh8DuGIEziM4
ly+Ojbm//1Qcm8pT8Dxa3j64595JVmcktxBUCsjlD6eni4duGMJ72C4D/7OnadtN
TxGmxMJ/+Oiq/ysFBpGjOw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9792 )
`pragma protect data_block
2dmrGm+BITtF1L+op7XMevBVcjL1XkcJLRKaX/HwKcr+JTD+TeMNNalsFTgzX7No
/iXLESDaJ9BKMjwPvzNB9aZbiI0YP2mVzHz4pCB1/guV1xCTryKa+i6a8nt9ej+K
o6eJOb4e39/Epsate6JJ48TGxkomsp6wSnozOjSpzetozUch8Otvcei71QlooKOV
ScLBpLoiSr7VajJP2RPmkzrB1Gawt7dhPCiKJHfjukCr9W92jvn5S5GzF+bLW3rC
m2o1U7rl7msNTxgd8USHk7Z8PnajOzhxXJGMXW+cwQ+R2KLyj+3k5fN70DKQ/d4C
MSK9DonZIE2eSqo297PYDlf+IdMLRcDKPRMc1ZIN22hK2T5nWzmfQgTtOybXI1Fy
AKIrsXKzrKMV40JR/Bkbo8W3RfyOn7lkeQ17cuUxYb+RivrPnFnL4Ejgft8DsYAM
dRDYcT+dxlghrQA4OM3Fash8DgoFYdS+Z1kwRb+c77s2qZlwp2qJzyGaw+596r7A
xY6igQLIZ2t68rWpLovB23kbl7INGQ7ZrK6SUHeAPGXfABYmD6h4BWkwKppE3TyI
0e434AEVyS82PvX3AppH4PmtKMjqFoAnqB+9W1BTBqIl0IIqEjXJu0BbVh3nAdaW
uki9dR1cw2GwE9s4tSoJPqy/Kr9cQvUD1yM85BcIbp0wHuTwFnswPVRXl2xA8gUo
3WO7+MyuD6YuHJ/eDsMkGzqNsmrexvKb2csY3Oma0dC0s8s26gGTblRqIEyw4tcg
GCtIdFYOhuG7Qw4J1Xj5fF/WoJVQKAUFDpxoDBgzeMJB2IN8FcuLELlnZ9wpaPkP
4BzHNM2Wpst60BC7hnQXUByl1baV0tX3olds4585mquvc7kFG5cKroyIWQay1Ono
r+fbQ4jwNTDLhczOX/RxC9byU1WTB/cQFEYDn0fzXDFfZmFyz93pWxxNXW2FVoJK
51qKeAwgk28KTZkSQp/V6IsGW8eCBI4d/LkmqvWo93y/wcvZ5Q292j/Rk/S1my7e
GKYkYoKmLkSnj6mN4JZ83q90LkdvOpHJhz4DzfnOb4bJjwE4Cp3l9FI60IO+hmrV
16A5BDhtlYyIm0HN0NQXnG5cCImHHE3r/UfWkuvtJmrJ8e8GghCivi82EP+7ZoBw
hrlYpN4gCR/jQ/oX28PS5DD6uFoWyejvnfVO8di+ANKq/Fp9H4Ek54Ocxh/FSYNe
9Vz3XTszqOrIUGm2TFVTARRJ+m/ubrumsx2dp/1+6l6tf2A3w/FsF3dE3UHPyMOc
Pld+TCwjeLDeBE+XFNyQ1/PMrLHOD+GNjZVO2ptPD90HuMo1rnGu2YY1RQ6MNLOe
5ago4Bq8NLzM/ewTGScDMIQOGMZmQ3E3/7/QCAHiguuhKVK/cFoT1r9Vcm5Rr9EE
uhe4h8SNaqeASHS6vQseUPpJds490COsSl9p1jaS4uBiQuUSUs1o6q4fGPHshKfj
dPJFys47W43As9HaWsl+V35pw4RWCKgFQ9B0V782e8dY/7S28yBrkI+AUbjBPpcP
emdyFYshteHpC90OJnVZjSkeSsE4BME0ASSmEJ2R+q0WWPvvYpvOvS5OfL74j2jI
v9PIkxfrhkp+0fjbFsiZJVJhdW+w04m9raOL2UOkqrSgP7jjhYXRkTvGHqmVYqy4
otDJz6gr1mXuoT7cGfYlCPik7LSPwrkippxPLQuRYVRjkYEzBnIAy5bY4l6mchv4
UT+BKiUEWALnBAEFNmmvMT/4jv5QBxjfQFKpXVwydBT9aio+1TuTDmpjC1JEm3UX
rI8968wSpUFuDeMgTruf5h91A/tb1BsusazJvPo7v6XaI++U8FBQLY7iEt0Js/Se
8RmlPNspwOMv12hhtx4AB8DGRDnzPiiwpPFsE9xiqX2ubO1lCxkAXcz6WpDWSt/r
paNgZ5hwaAYLfCf/5fsKp4Rby0Xo5vWxtKUPAEjmrNAQHKRsLsLaZkxOBDpai8Ft
0d9qTRswHU4Nhk7ZVKfAotUuoW5Z8QF+09RokKLmf12bznQgAeQZkzRrIQK1mWjm
ONs6Nk5Jfk4s7rMv/5WYF3SqqybNyU0020bOQ/nt+GJw7094QIsuIfye5y3RQIy4
Fk56HVIvJGW9eu9P3zlZCYfZ0wwiF72tdvXghnf3y/RBIZqu8Z8bqfEYMXlrCZyp
e3rq3xWlwdE7XXvC0TzQXgw3RW1KXVD7GNMUoZqO+ISWLu/nqsdH9VO/WrkcqM/e
esyX5hzPMOoNGP/4jRsI5yEQiIKw0hPf3JFfg6kxWTxrURMBVtcJvYTuenHNTjx1
tiKDak6a3eZ5DJMwox+MsyPgRSbbdTdKYKGMp0Xd8bwb2OCQ4CrncoAwmcxyUKZA
sHcC4+YhNcSCJVhbf9vrjVhNzomzshyrPqbXpQbPXtzwHDdZAiqSBYUfrSKM9ncx
paoraxDRxLYGr1MwE9UnhN+6iS6vTJfwJzaSbsfFUcdCQSkL2ZlzZVwfWu31RJtU
F3MpcXDhGylfysNgoEG8ZDOJzRyxTJpoXhkIEgqR/ylk1ccjHmIJJOIRTKtJgVyQ
zp075UkpeUoJTEIsD2ptRufmXGKqoBYzaX8zTTs0UD4gABhoWQDeghIGkYe1BrJy
D7b4rLrSWE7VFESNDs44xijkgzc9gM49OGQeXcFjvY7OqdRRw4G/7wSrI85Wj1S2
fcRZ98vOjNrh0Ol7EootMTbzBPLH2z6zzpWGSgaYDvF87aOYlWclPcxzXR5GGYKW
5fEPBrWF7mHGPJ7AClPqtjoi0CF9bmb+mVU4JPjk48Gj+7Fyouqc/hs6RhDV6gNa
v+CVpg85NlkWk39Iu8vPVAQc1UzQJctF0erbB6BiXL59CEZJ5mL48mL/QGxbeDAN
m2sBKNGxLCRE+8yV+tbsmP7HL3CZFFs3JzDy098k/Ls9k2KnZEsEDDzLF7XZEoJc
psDHWJcnaCJTtXeeLBjHdwaL+as6p02xIRdGaFbay6LZAGnKxbNepByb3Zh0fbsv
0bnEH3aPYOhDtFmaBrZl5L4thVy80TqNAnTrrEkMH93yog1UTYCIBQtEUB+EM1js
i4OO5+/lNMBSJTMkWN6io34Z099Ph+BQw9qcX7QO50csgc68KOHDoNLU9JjlAfcG
4maQo/Rh5IMzLt2Y6CG7Vd7fevg+HK0aDyCH1ZBosRXcrUNi8jqC2OURQvOVgYXu
QNtCpPzy2VADYIiD1MCsYuuDwCyWJ/JLdxwBMzJjKCpIoM1zdWMyb0hEU5Anu75M
n+wxt2NRBN/4qQHMTLBkS4YcuugZ6x9W/Cozcl/WuVhb+OLnW+bx4DBlc7V+VmXs
UskWm1/3iRjdZlEetJXdBFkResOCkn8SE/DWyuAbh8jo/U5Nv6/xbWSYcis0oA7V
beLJLUrLrtLjzLVro9rGQNTdUeoxycGqhpI3EdEo+6O7mFX4tN+JA2dpCh4IUo4b
OUc17dQevt2KwxS3yld/6BKAyQ1ozlCOtTlne6Y26aHWiD2ggRolU81auf8wXuCV
97ztEmHXxdJST2KO+JPQlWUGkzt0IMX9w+HFyUwQEACEG4WtfCiZCXW83T4cq98E
q24il+XXTzXFfAE+kKq5B9ye2EtJ/ypUQsKnCwMfqSfDR8py8Jg4nReamQAsF0yS
ODp9umTd6P02TkKYbYvjpmMRgfWazv+5wqX64/SSPXHPE9E83Ll2nA7BIR87NMh3
G9bU7eKSdXYv8H54wRL+YuDiW+sQZvdjXYT+GzLtnBtMw2doIsnD4XKZeK7uTWeJ
o4Y6fNWNEswe6Ggo+OEXyl1ocrdKLB8yL5xbEw4KHEz+Fe6W3OTAMfPfhaWRzXr2
nRFAA71isHMqhD5Sb2yygUB6KtpWIsf1z7jyPDupNFMxVUAiNwpiwqKRuA9+cOfW
dJYJ2vRiDLiGVu2DTX05+EQSqcmlMetsk8qOrRIs1xjMQrOB5GOjZUoLDmHr2Om3
25VyldwfUdtdIarv3ZorhGOAbzPchSK+fFVp1cbegd/nI5DJmOUddf3/BaUFqrB6
KUwMES6Jc30HNYHYUzLlNdp1UIj/uUX5w0NEmUwCF7bdhz+deqIqkH5BPtKrlQ9h
bQ+zXW66+oRHlQ466AFnys38t41ckK8itm/D5mRes/6BCuCXSJsB+VTk6Vn+fQ3g
/0Y7xL92EdfIIZM53Aa+2GGdEumE4v8pf91zpyDqEZsbRFVfRB9L9iutdD3XovqG
L3866UtgqsBSNhuSa9AhmUa0RxCHcG/CdPs7/47qXSnPZN0UexsGUYk/dINsZXU4
TujGIZBkf5nrn1jlPUm+xjL1yAHVKquZjksnHKFUb5CYzO3A1ziYd+xZ2wNtLOHv
+LlQtCilFOPZ9Hi5UBQNcvHbr50NYa9bUNsrI7NWIafO2RZoRsLAr9eJfFiv1G07
DR0lX7MIWVcQAdFeuyNmH6f7KiAdIKsgHb8k3g/EuAum2We19DVMLY/Uls98axip
DDWsjWvyrGXfUF/nbPbrnqgckIve1g6VmARoAqa0oXlMWmKb6a+SCjK+/d1yoe2E
iq7FmeIksomTNzgzE5zNcf3w9C5EPW/oKD3mOpI2i8CoE8jLxZZb/sny4PzA7lO/
Wj+RDJcyUZruuz7b9r/qp8i0SOofJuyyNcwYchOIONQa6i8aOU4DEnpmbOSI1Ksc
huNcPqsipT4u3Z640XYiiAUXAVlnzoW4FRq/IBjRuNBMR/uURaTsyBmXkBydVnTD
qeLFX1gA5cC1fsR7j0UXZr5qse2O8RpI528u8QzCvxq9D/GlygmLqfee7uTC04ls
yYDybEKfGgRFwgxohWrc9gAv7ILmgEVcMJcHAP+DIYw71GAyO437ZNRrfx7ZR7Fb
ODW7uWqn7/1p4N+rpI+c4hyI+WTtMa5nUtFYrlG4sk0QGoW/uUWxkSRewjIi2P+c
Vx/f2c+alyjPKLtUQ4N2BYSebBwh4sHsPQOoxkoTNFdBdfVhcrr6UMNTOfUYjla/
M4Fd9DXG/+ky08rs49we1zVm9ThtNDjGHKvh8ohDmv52d5xjPezlsPXkl9S5EVT6
kafw+LTDkWFOMGlo41CewoMyfEHDAVj+LjZUkc99f+MKe+qP2cyNQsIEK+IDv8XZ
Z04x+pTwTiDIWRd4xXiAoacCdraMl5PPcUnDEM0GqG2wluNo6Gjz7YhMQeu79GIS
iosMl3Lg/1XUfglGZW2Q60oZ6oR5ydUCNoo1u5k1aa0qiEaXl3oD2EThYMxerISC
kV6chNT99+ThweKPS//H9JjGi9lDvI0WTIKS01OxbQ0ZjiDO/56JKjQam5eLMc1w
LauELxowAdJmMJr+SCrUzebwMba8Q09r9AFRV5e2RCPZXJiztf1Ab8RZi6eXH+Oo
xFKp5OV95XN+trHv+mkVfnnjrQSBIdgULTtpTsd2MN1MJGE5KGSeza7sVC7UJemW
Tp5zj7kamWMP91pFQNKLN2WMp3z582Ju2W86I5gbZJG2UddghjBQHliHKl/rOI4N
zLpgoTnQTZdwgfP58cRzexCggL6ELVC1L2WfCux5NoY55qFT4DH7QVSp7DTzgfUM
UAMHoKFKyw56bjPVHlcDwbFBYDXRLxdxr+yI9QKszoDX4+oUUWTuq1Pyt+g29ANO
lvbzq7Tbqu2z5yFhEyGPP0OO8vCH6zEwpZcXS3TQjVo10OeQcGjH/HBBWtTQgCbw
L2vAAdunY9dFoU56QcDWKWoaIeo6RtdX0NJNoM/uFqJHonL0s1u2yN5ykiZbgbRU
mU/wq0MTSi3lQgwnfliSeeQ5IoKupaJ73TrwLaLFGgSKa8+TWonGjdMz1m3SejtO
FUmwFV7Zd+F6/Fdmkr8AFUbHB6Siq9XX2XdDOxgzfxKzM7ppRvgk7/dJGL/44hKc
OiNisEbt+M/qDxPPToUjWg2uE21ImKQIAi7nGRhN4Z7zoYZ57lp/B64AuVutBxYE
m29D7t7XbbTAaeRdIjNojNGr7WUyi2CJVCk9jaX4AVU8Dx+qDxWZ3VBYu+H/mKX8
hcSZ35hUz7mgfsSXtQ/gKPzowSgFfQ1tWKog+pXvOOtRVqS/ou1l3IgbpiBBeEFt
UvydyH5Kjbh/S8rYzj594rHZVjXx/UEhv+8HHm82TY1izQT8wqr9HBPou2WmGvKX
ONXFF0C4D/dIxDYEsaPN6HmZ91T6BwRhHHxEDjeUzLDRqhbGePhX64OJEpOw0kLd
z5x6WRyUVuFLvFz1Y1mQo/1nqswovtqx5atxZ3lKsCTS++H/vvVgKCjAsxH0sPkb
zbdbYD6FrmAoDUO8BQp4wmnsja0CXCjCLjb4c9r8wzNixdgmIYIbdUE+9a9iYMK0
DDsZdy5dObzJZupM08hPPtOIW3gUZjJFCCghr/WnQlKzf7wghfQD2Ueef+V94ehX
gq62UuJ6O0xSwXrHkb0PLhLKn7s83JT9CFvpG45vhzMSBYAutdSDfQ/UMI7C39HQ
103/KTRoJBm+ACCWSMq5Hsxh5wPF6ABxDFXJ5Yleax9rkFtzGytMyEW0o77kl02R
517+hcSS82shxEb90fWYyav/D6t9Pbs5+unxyweYeLte0JrJVZtk30kqE2FXguyM
feJzkaUwfyYq1iB7Zpm/s4vH9JG6EWhgP1lpDscz9qwYMXUBqbhTDk3xwuMvxWRY
j50jHw8f3l4rG0/37jxCJT+CLkpaZy/ZY0k6YbF23epKtaBpivqthXHDJgEN9MQn
RE97jZW4DqYowGlQprBROyarg40Qplm98nhQC49bcV528/VCCqE29xK9e8cc+I3/
dL5p4TH3ZtM0cM+BxQYORlOa9o909WPgbrnTnmA+e0DAu/NKEqp7aZhGRxaI6fRO
2mhTRzoIKjns7kUI8XDKF6/iXJ4rCS0idMVxHO445rtUT9fsF/XwC7bTLCawt0Ax
62BaK2GehDwdWg9hdq1P1iWU4Tsgie3WmIpx1vyUECP+IhW0CbE/CnkdszSaQqvM
khIRYPnPQwGBvBhoR52b24pRWcejxHN7dcTfua6gDImwnUNy0LKZnrpG0o42HiW5
Z+5NVPLkR4n+agH7LYk7yWNVcJ4QE+7jMIzZw+1tqSvaHJnqxR2nCnWpa6wk4g2x
XHkDcPvItYvBX0ONmX7i9El+uNU6ZnY60Na4HjqCUpcgHDNu3nC/H4sOOj4Aqu0z
vmpe9STXWqNS6FmVXvPL9nOAdTAgckN0NFOiJBbtRTzvw+JfAmH+dFDwKTSiBfA6
O0dsdQteiKd9NCMll7XpdkhV1kJEpDnkz8+1UEzaP1Y9OUJSP/KWVNxHPaTDtgzL
y002cIDBp70Lc0uZW8OWm5PweXi51WkIYVNlxZyUTby24YtedwGjbzVdBS5HO26A
odAgx24qQsunbV+pg9tCshiwvKEbz+RDTGPHD+RjgFkRjemC0+NWBHbwUIYKDMd2
ApHNbKySr9fkwaDulFrQl0qtuY4EmBRKwpKc+RcP3kBT7LenUQX6KhXICYzFpQGt
qw9OC6PfFkxmY2T18TR5KfltKfpqKm8hdwoECzqh7WRo9SALcWwMs/B9bS++8N/S
QNCO8aKjZ5uVlW75qpXm8SKGTtxt+uCusxlbWF7mp3XOg01+1F8GL71CcbHOhUEk
6yh7HjmcTp4Kik8xuGgP4DribH3Hniv8WjWo/ELNV/gv4R1iAw1Ujs/LvzzHhNTQ
pEgwODRJIg5x4t+jpEiQtQCR089PpsWH2eUB+U82TX4D9BZNnFdrWIk6tDeJkJ9n
hQNJVVgXxqtyZiOugcAQhwoeE0WlLF3DVnCsYzZSiiICoLXJhVKhY6CxkUFNTDql
q0k+puMmmej2uIRfwpt9pa5polWO+qpRMk229+izoE1vmx4VBvs2y7LTLdbX+gWV
WmIPI+3fMqne1mH0sZ5g2tFbg7/QleIpNU2voPV6PE1RcJsjw/XMs5DiwA1NGu4r
VE3bqTrivpKiLGun/yXgQgrUFM9ZuEOdXeX8AwtMMOSU1AossLYJdUc2xygarZzM
S4cxtSDp4Kr3EqEURisrDtsUB0WzMF3uW/RhP2rK9FSskLBG0ti1qZRaHYG0MFDc
rEGG2kIErfrUQ96awE4u/rHeYHNXS27WmPSFZ1yVc1/X6VeSpZ4/piy4anAeEtxz
xBhJEX6XuRwNrimCbKaYwYeyVhZbhk18FBEM6zUEsbceArccuJBXLHjNH5gSpzcn
7CTIPvm6vVzt3YmHgCin2fz43/JFdEeYYynMBIYdZn/G/1pTrGYPdqcUBgbju7v7
uxHpt6MpIJuGcRJLOfBRDAppkdsZ4lZ4z7QrcRohw6WUjEmgsSTDmOapw54aP6yF
Vp3NA9cdWbHUsV+vhL/bjRpx8uGao7XqHUtmnlsQehBHq8r1woOXZ+cxfF18ZWiv
I2xqpoxDpWi993+iJclfWVPmgVBHh4mFur2Hi7xsObN5pxQ2GcGuuwpxPGgRzkBK
TVK83J0ZM6xdc3+Y6dQVJGUji5MqjYs9Rdqb0qf10TB3R44oFWla2YUnrCssT2mj
ooeKj5jMNn9SARzDlX19Ik6uKgajSGodKNKnEmUmGNjVhu8PVVSe2Wi58pxnJMfg
7XYCctL5t6T9IOVx0Ynw74LvzLfH/uXvhw/WSsBLZY0EmPnSEjfMiAcEsVrcEZcu
4ISn8M+UrqBffq1FmGgmDarC1JJQwzpdfArtApN+VNvXqwdNQ6eZP9QCCmOMrQod
ARvkOSfl8bDSGIEWYn1BdBtdaWt1yiqXnEolT9ULhQEalj18oR/pKyOCrks3Ehqi
O9SRagYunmesEln3ww8nBr3vF1UJaSYsqfNj0FcNQKieY3YwTLtuk1PE2kOSEoMI
D2nv5a/AR8NxOVmZCE3DBuMPZCHFhZ6RB7Pc47Xo5VTMmz5V9DHUyO4fZPcMA0pg
Ikjkw5rGPbC1fhRSm8hittV22Bh/+F6PbEK88QY6RvFI0UERusZX3qWVrD1yGSit
sax+pEfGLyHh1gkKmFC980r59Izh0gtOatETM8RXCxIVdu2RdyRsfhaEip4JP3gK
h3gF4SAaYH9+3lircooxf6STek8kNJmvp0PYCy8zsS1luENB5HGD6wWbpwUY8z2/
GskgOm3y0kKeMFadSr4MvHVBuhywePll71m3dD7JZ2WCkHo8vLI/iczRxtc//nRp
499HfEwQIg/ocHtgDrmeyecAtsBrRQOweTYdx33qyXntgeJm1RmKwncS9bzLvebN
9NouxIBHjGasWfBsfIyeWoyE5T29+nptugXxbkpS7J+E1vjgWNjAdGg6V5xeDFEJ
eRxIG4bfs/nM/cIceraDHdspnYC4he1Fxm4oIolBYLB0hKoweesn9q9fouD9JMkX
XSK8vmRn8CbDaXDpnJ/N/tY+v+3Pi5PB0HSrXZS9i/tlezxeN84jHy8RuuFXjq2X
h2HbIms2v2t08PGX3xfo+XESl9N+NRdLpdegQtkRM/fjQW5dcLrWrGNMpDj2rUf8
H72DwHYTunKLghkRzsBgAw/Zwmr7tuRZ9bOcbMZJ+zMdx/j2hMn8AbyY2tidNwpy
0y9dLP76tE2k+iPlJVvYecf0O4L4Gh7INqVc+Pzwgfak53OrMldZHY509jVtObkc
/SViW7F2pYdKwAlS6NkRdqnml1YfBQGhKmyIx+VdaIvI+LTkHhq6SqyPAk9/w++6
fqcZvw1AVlpbSTObzFwfCfQSiZZr8y+bQg66UbNomKUH6AoqjT+jhLKPbaPnvUcR
OMK6Q/Eo6+y0MK5fMkwXZVGZYvi+No7nsdyv2OetwRNxXK9Kjhk4Z5U1GOHTuhuq
eNlP92Fe2ao5KCC9t9Q5gNuz6hybRIgcu2keVQbOrinx+N4QY1fcFJ7xxPy/R5Ju
jM/pR9yoULia9e12SlzLSI05vX29SzIqsqfAQnehK4Jik4RTtRy++BmaCy/BRUVw
LFKBcgUJTO5mK7TAnCENzOFpr3KVwTVZFVXVLhqAQsqq20B0xj/Ky9p6gbOBsbJu
YHaGE2dXolgWT0DPbJo9WdctLG0en83yftGLkJOd16QHzZldbl1W2qFm1XisMICU
4Us6VjOZPPVdWQIXVCo49f0qs+MilfSPmS/pMor4TsRGMeafvmcu2f7B0ibU1w7H
B5L5Ol7/on30OqY1/MlS9ga+wQ8C0cE5T1SkAwx/eWzefk4vwMYukEaZ347g1gq5
6m3fEhaMd2dzDFNNPWHwo0I/FuWF7AjSmmxugdSVsxaG1aLUdI2QiLxwltGeh/Sr
PyYvmfHodkD1s+lGEGfBchbkqTbzzgUsIMRvr47VwnURqueLsQMr5pBnNoIw7c+4
4+aB/CVLSiT4XShYxdRDKI+35jrkMhdd7ITyJHkBQM1NX2g0uPmwxCl1CYIOrZeJ
PCEZohD5+bn0sJMf4SJlvVQ2qRPnwP2eL584TU4SKPHJd99fa6p9MhlcT0C0pePh
xinSDM9CB9m0auq5Ww1KGtRF7kZ+0hELYisEA6j4Y1By8YIy6ansbfKkFcuD0DbC
PrW2WcPKe497ekI4iS7gW8DUd8ZcOpU6LjzCgHWVyTeT/qyy4KhBTob+D8flwZM3
XTDln13yUWZpXOIpegOA8upVTmDde5vQbGYky8H8qcGtR/7XHnYPGCDsSdNqbCC7
bwXtVkveLObpcgx6nxG86M8zBKMNdFYdumLlAiXLB4Kciqy1tAHO1JotD/t7D4T7
OYyROWzwfgDhjamzS7DX1EhSTKA/EtDvnyJwp1DKJgY+cPz8xpYUZNMiO5ij+avV
iloI6a3Ncv7dFBDOdXOXfgEglbzVmupkfINdZ2tRtR7gsUOs2Spy2GLVYhgX68tk
UHHXrT+bM4lpKqX78a8ttTsbN2JnCyR7/8lBzhb7y+ZKzo7wVjMsmKtj0exhcpvb
WREiNiRVKskeifPeDBcr69rM2YhvlCXKdi6oSoGWWY9X1z5jNHrm2HIBgvslnMuC
ZRwJV72UMaSlxvDpymn7/HOJbTvQtl1PzbUpP1Fg69hORxPnJKyFEItq+SkETYt0
e3fzue1xyQvim8wubJuCJSXZ0RCKBwCWBnHnGneGYQs66Rd5AWpI0Kt5hskK20sP
L8TNQPk5qW0rBcu/9ccKmG5cTt72J7bMdQ7MC7QXVlQ5MXWwzMY0tAOcQ+unE4oD
G6UD/92PiPo+IokvCO+XTMUqPEJZewK6JvcSEWYwAyU38GtBD7cSzBJBv5mh0rw5
qWmktHMqn+sDQRN4PJ3ALFg2eAFFbGL3pH5C2X0Va0dypOlL+8rgpb4yW3XM10VA
caI1cL+36jwGqWW4Y4Wghad/fA5VZsyCdUkaraIJT0XodJpQEJQUVFUFCTZunVVK
HyalnNHcLP2O69kQ46WSjXs++CniFMZdNgH2Qdt+sg85zqPwCkFmBMmV6h00zUgD
ePxrThSyioN7MkIXoOZKZK7HkvL8LaCn+1asrIIclM+Lm8MgIlbsjCOpZ3QKrczL
onU+0125UYISe5KDFYArsD4bXs3DCkwCfUl9Zr/87BsscHrnvIwIoyMgYecrak4p
HsJEe4pzMnQ/mZEY4m3sBVV6OtLHAquf7DBl8+TgUKiUAQ/mVdc7Np5TwVkP+KbV
VKaHiHSj9fdlmxQBHc7FlKqzp6kkTpNhrGmuvsxL+GAe9zzAWW0GWwYdipihOEcK
VFnSnMo3YX7YHdf2LAgAH4OHHipDRV8O4XGVRhxjwUo3Fqk/DKMq6AG1/pyzGvfF
EP84wguh+sLLUt7le5fz3Y3k72KxSGOgh3im7hNXnufU3vto6ZMOqQ5S67NAUuV4
0ixUugujkvJdZmgPjWJc+i4Nj7jwHx5z0aAJigBlfBBwfrlTrifD/HGLs8f5vmvQ
uT24iEmI7gvw1JQD6TklDzK+RXZPd3GR4Lz2SX0raFtFDaB6JUBRupaMpXC0pvtp
dqIjzQzPHD/kpoy6+Vo+UMNMkNt3kfaMbMUL3Pc6M8D+7C7slntVOHM8MwD1lUA3
x4aFRueV2VswjtrD/XDd8vcJ2c2qSwQ48Hzh43KHHl+RL+pWqTmfkXUjk9vtP/bq
uN3yzbbTnfBOHF2Kzlf4LpjXn083aGkGvj/pradSju6oeo63XUaEE/Xez7+ULYfb
nQ5NYFGgAKc0li3WueDX6Iet8f1uan4+vlU9w0Mcv5+CqmoiUPzUMeDZ8VBeaVs0
tpoNR7Yxy6YImBqDKrrhRAcFfWqCQN8T8nvkgtWBobdgBhaaTpa01cXDZDQuwI2f
7E4fA24UfLxoZQ6QkaRZY0Zabxisk4uUjf6hCjMFgH16qUxiycgmS1ES4o6c8kF+
14yNjrgjR8IEDa+B19rOb0oJUm6SRNxMPOJ0rMybwCRZFVpjH9ojfAR28IdAe1OM
urdnjvX+XN+keWX4q2FU2OuaV/MyIOHbtS+C8GEttXQkHUQOJ9z8QojZywvZiE/M
UpvLG0d0gxJNLdEeMfgV7tgVnQQI1s7SwztzMbKFfdSetJTwxD2n8jZ2WzAKkgD2
Fj/1WbD5jy3IhBuUragQbFTqmpNoKSTLocWaQoju5eept/YrDsNQn1yhAT53p+SZ
daJlkRbCnjd6WkNNL60stnk4CupgTA8Il37dmBbY95GtTfq/CounwBrJYcCh3Qzi
+Yne+0HpFbLJzE4D/mchz/8/8raWS3i3MlmdkMLZJDShsuNIFTdnfnRM62WK/HhM
pmwuUDi/7ob82149tsXtyo0O0OHzUvB4VxloVhyaBRsbKYIi+q5unzr7w5yCgejI
vV0e/UfYu+BFf8ecTR1lUDvPiPE5PrQGbxg9Re4H3WcnsAgw5JC/LKL9ewXkpUap
zcaqiKZLROTpwF6dGsl8X1TkAZo1Rs2r8++oYy2kEVMZDtCGbWz+LLU+66kCk1iZ
0e3iA0BLGAHFiD/3GbnHiGOfAt1tJ3ucD5Ky14kvHtHEYCjamp/PPRfkYbr5rIfM
hQ1SwlLO0He4k4cwJw/TPNN7Gw/O5/dCGfTxjzC9AbNoW0U4+mYH3LKaPnDyogXA
Yai5BFvOzAFTgjlp5+FmCXTXtC/x4fUhAO4YBZyfnQLjI/AivBf3fOQAY40zDs49
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ZZxamlDgJbjaIPBDhJphUGaphscX4K6OFc41bOt71jwUI9veRkhA9gKajYf/25WO
lwrBtBh9dnoE9FZw2IXNsVQ1QGCgniUKWuROSnegtTlDT1GuXRkpwxP4uH+d2w79
7GZv9O9LC83l7idywQUG5hQ68xjZI00AxtYAnGlsp+cEqzUAZ1Gjj1WH/zhwrkoh
gdlcqab0pX/IRpFQ3dpksItIJIv9mVkf0f5qFgXC/06mlJa+5GPinOF/lzWZBfP+
GNdFqHgcOAjAI9rBJQaFoCHRU/+ZWO1B4T4NiFeeQ/JboGT7rQphwTvRWrI/Auf9
fPMoS+0/H8EKXhNcNtRDlA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6256 )
`pragma protect data_block
jatTAN4+GHe9Sw8C2k5OzIfrVCjQz503fD1tFHLzIY1xUt/w83cBKNZGXdpQ0ZuC
oF7Kmc58uih/pIBnkIsJ6sY3MOZefdMt8eUjL5kLyOxqk5XILX40r2g3zpzMiqvX
6/MexS61DzOFbXHGvrUSlLLBw8xcfL65vw7ZJG8SH667XtlTLggR7GkwzW/JbAcU
weBHgF5AP2ElwrMJNVa9A2yq+KxrNZs+ulOjwzXncPnnl52WxbO1KErazb5Q2Ufn
rB2CF4uMOHs+mrNjVLbn5d3QHuT4rbxiMX7TLQnaGYpiuf5Gtlpw4VZeFAxq3nt3
FudY3YZsnFU/9Rr944NTLRBMNiSvI95gJV2CknrPsj9ZaD97ejR80Izm9VnAu9rz
/FeIX3SahZI+z3oR6ymZZLmGzc9CaOKpr/z/SHqPgkLZNBtu9nbaNChtlIw1vFl0
OkJ2uCwP7bMhUUpHWaYnpNSseRsxg5k90PKnRWuikjBgesFSPKtZrMGF7nQi17PL
t1tQuuI+kd4/vHxfgkU2jZCIEka1XjKCPDHnGvEu+rUq5s5VfRZA6SUB4KR1acgS
Z7TIZJ30zHEEZAWzaA3vE9chIbvpgTbaA9hKDAj0PyxCkDE0Oqm6qvEW87eDWqZE
qkfKJr41XX9wHD5agHzu+5F4NLJ6tPCdXn+6qEatot+jbAypPCU5tD6BM4MTHV5u
LlqRSwKus15xWBTfHXeXIIA4C6KwWUVKy6knu0AHI/rABbQBBM29/a915IXul0jd
+sSH3SYtXW62VX+g9LYFwFlutIOsSFp2HOyhuOEEXgaD4L604Tvsx6QQe+D7JEY3
SXk+HZ4tzDzlPFIxUxBXu3BZR/10JR9YUd8O2a6UbYRp1xKt7yoa/hbhrY8OyDpk
3kfTwdGc+XInkv7pniHl4csIjAXeHrUyvO7FMz2MCbCrXdc2+wSWKAYb/ONpDAdt
KPnaA+zK57wKyXRi6Bxdef3cxoTSAGOJaJs9E3lFKqHhpIDCH5PPGGCNZARDInVk
I/+aT4RIMWqWGNlMte/9fn+3shAHAFyIg1R67JpxDRXChJtp43f+JpgxVgOu+6Wm
wyjCWXUtbC1ZcmIxCVqJQ4PfpJJyblRUfE4qWWM5PLgJAoBwma7J8TWCRTpDX9XR
KmtBE5N0Hu9x0WJgdHlxhagAY/AtH0V2BPRoaZ7Pu54jBDtoCct7XcSSWaHnDfaE
4LzmhUlf7OKhvuuL4p4Yr8p9W1eH/cPcoX7gZjpk7VQJLqgC2Of8bsoKy1Rta/9n
6JnvHcgSxfI5wWylANdRq2Pg6ghmMSu0CKiNnfuA930xWPX1v5AVecXRMqm6MEaj
56HLefs8Lo3tYoKsGiBJMTcmlXMeR2Wd+25EOIctN4K339ujB8gW5WoYBFDkSEu4
LHOuldt/furt2dWo3DrgEAjC8Np7EV+I0X0ivmbg5ptTh4tmP03vnaI5awRRYKLQ
ol7oaGjENWP28ABPNx2GCridgiXU6+lBcpIC+RSEA0YZ9cTtiaCyiHEqTjRIlMg0
9cxNRIwMbOkil6Qp2kh3mqs/5c0OuNO/BX6BEj87QCF4z4/Jqs6ojjqIuFzHT4J1
Ego/1qW23tYYWbyd0YAO9WVQBKYSYoWljoudu048kEBLpSG8+zL/km6hy/z7u5QQ
plKLP8ZSWeHHNbr+bMHfaJPTDGdQ2mbf4j8FN2pNTN7v31GUqdsIzfuoLI+nVOBP
xtF8Cky+KdkQ7fL2M8Or0oh+/uiWzfGK7p8RM7W7nkMnb45JCJyHGzECDZzCgibh
9evGAVsmJE+7J1QsZZ0Wj5rHiZwDMZiMpSVXVPAZaQ4kgLuUDc7mHePydM/NKYO1
spNRL2OT6nx7fG15EIAzXi5je2JoIYOKxAXrhHDcC3Cw9WgnmuTxUkTh5z7hZkKN
izs02rBbTekrqupxjDmFSHUGXLBsxrCrSFsPiMa/l6+nmxHTjp9ydsl1aTWYgMji
CrnAWmr16Iq5NUiYkBus5GQz1t1+SPat7dXHWBe3Zz3KjADXvVvuylZr5IPUXJTh
leu7i0LYg1UtSo4SWzq6GSuehwy0lIjCW+Pw/YG2XdBxCruT8PFNhYnS4AsO5qSx
ZHLrKbk56RgJC7Rkib8Fw7ELhO1QhCIB0TOuk4xTehTroP/nzYki15sjBdcUE8bq
YU3+H9vyeHKa4gDqMGyrVPlwXFErUrZKV51Xj2NPvFoNaenRICwJXH+PYO/XbqjK
/oXHBaaUCX6ojAJIBVzgyDD7Y4GPitv1VfU7SwSjES9sNM5XLQsmPGTwlSvNv+Mz
qrKiwYOSpGjYOSvdcPFKxfbcFVrSvZ7+qhPwEOxNQ0DkMHDHOTVfFXl05ojmvm6P
dv5TvkZmXN0jrW7aMIwCanNYEsmeG29Sijr+AB+fwSXHZa5vu9I6ihS4N+6H8lHs
4JL8Es2jYybAVVaE7d1iK+J5mTjvptDLYIar33EZLdhT6nx6HxL0G7QBiy8szZLS
t2pAcO0s1ebsBYsthQzgv3DKnTUa9BzBKR4BvENCUSDQIBK6YGTXKSrC7QHd1qey
RNL5nIV9Jgvaw4LRoDwqq0oQrDBoEA+tpNc3aAuX8oTCUaMz5J4WY/k1VLuU9B5r
/iPYJD5nDhfNCBmxs29L9/ZnmzPvYRxKy2VXu3vhpeJGpAhY4mOhdKnmxIYHUiy9
InFFb0+iQ2UA4jcAmm4tZJWvDyGTrJ7ZqdUk6phrKK2E9hhKKkAJ/bhgp9tSy9+L
0rc75VgpHDzCGTUZxPSLaJQot1d4nPf5W/+Z4GtEdvzRv2jgUY/xzqeAEEApY0RH
nT+CBBQJ+pQezujYeQXF1K1iVINy2mPY4RjfXqWzfyE0TntdVl7ya44Nwcpmlb/g
sYutNXslKNLpojrVUqFt5KLE1NXw6IQICWqCWRZLN+09GANUdyv/s2DRc/CzKShP
tC8x0fOp+eqpUWwb4G1TFPWkXaI/O/0iYB2rFDZI6ZihEZ/dnf83palWhZozaXpP
EQ5SQr+dGS3vt6GCmYDYdIbiYypq1iNaS8fw4kEJpEogeZqt63jCdEOFf/ibNU0v
kMnpDXXf8brDJMD1kPVmUj9en29nx9nWzqZv+mxKWjTrhw4irA/V7fRh6f/GDhX8
DMlm0re39LskgP0BVr/C3KGXzlwxPkVl0MwXpSZc6dEZooMW+15ODI0cUCd9vEh1
RBnriXESovdpGhZcDXPlMk++L3vQGDxFiI5KWGWsXH3fAtxx2qdk/hJoQH5Ruvrb
ZHVOw7hIZ4LmAyFlB40+0UpbsLgmm++ssOovKVfmB3xlPcmuGHpSuOOtvnuGl4MW
3zBnnFeMZZsg4fWb6YLc8Kvv4sIOcbLR+xHlwivDvU01WHKn1lMYJ2Zn++i/ZZW4
p6EH3hdIIhBiVU+b7SSttSMNBJH1MangS1ehpY/gsCF9r3eyS/73Bt/xDl6QmoVi
GfJDQXGluFZm9NT6wyyohA5dnSUUTM8kQh8q5k05uh6PCrx5hiTiKg4FzFiM5dYf
D99xcZdRl4Ioigdg+mTRwSJCE7M5o/6E7aYF8QVXcE+Oy8FwVkhDSWWHU3NLP3Bu
QjgQpHCuRbTleM8krmsHPLS07vY6HE2oTUhMz7fsfZmI+pqOtNJs4d50JjjiwdnW
sdPWRxEiWmTT56zj2aMmH+fUvZU1RFFo6x5DA6CSP4MJ52SxSKFw+gnJTmHofE3E
sQwFKSFUMwGsX62cCd1OC/FIFp99pyMLZLRwfuwz4FJEA5OkOAX8FdDY9yimxhHq
ze+HlP0V3Huw5TUvWNUlbRqZZBMDPcXVfoSDrYsXUbKqEjUTu+jZPlxIBQ+OpQtW
pfPZkRmMvOPFtunzk4KBtFvFE7JTxn6fTwl5rWdGgglzBXWrpFEjLpz1rzIh/DHB
aIV/hwI4B8RAFSO9VHzNQl/RU1+XVoVFISDLWDFuhb0AF+1grPcjcuxS+HbuvoU3
+Mzo0h0Cl3ketcJPRDT/acOwBBhJ5FJJXm0ZoZ1yxm2m37kJSb5mkAsNp1k0g4WH
kuU7jyz1JfYiKYDTJGjCXDyM+cfVDrn/FoHBykVpU1KNFubFL2wQ5cYdMy6aatMa
wtFN1clSaa3U1FPezVwHRXj1P0aW4PlwoqXJT+V9OfIg8BR5Ryr1IGmGqSHzjHtX
mEw3YUkpwFyBJj9h+d55xxsw6WmJWWbWxbUjcySrEc9GYdEWXNNt2LDQlUfFDBXQ
a1aqH8SN45vg1qjtd4heVGQDVarp8vDrJ++Za2PcY9uXSvLs3acJ9mPfNWCVOGQX
OTvZYOs2z8FtiCMysLbMEV/lVqjnteFZ2YAe55OZbTg6zYexD7ktwEAPZ9HccFgr
BPBke9buvSxSbLnb6yefcqwt5ZT1Vf7NsCsXrmQRcKGvRbz5CEEqjtzyk2NF32DW
s1HT2x1J9eTA5TZASHLxivqsJ8EUqs+a4EJEVWpXpW7LbhBYTINBrZOIeeWZUaH/
quOdzzRt/1Zc5iljQc9ZGemASElDwFUkiK3eY5rN2edwufM0gHt2g50Xyvmabilb
MHrgYYFuemyF+nmRRRQB1aacEmUj33j8qJIYcGNuPOGt1QeAHwWZ56PArfYcwyz+
VwFkpESLDGPik+fVa/eb2cfN78nldOqwbUJN+Yo2rgspMtb3l3lTXBktvYuh5f37
AQukkCwE6uKbjoj6KVf/MSF4WrBpHGCLAWfzMoS/q3K5bWbqPZjkXaqcWdnkY23Z
Qk7ynUR1Cf9twrGL7i9E7bLcEjmdYGvDV5C661EzJqR7nOm+tEjlLTub1Oc0alwn
6cVqlYOuX1lKjrG824Vjb2m4lELLPJohSyYHqfdPqkJAf9yD3+Qd3RvX46wm3nDZ
xQ/loxijsBdVLyjpJimN/aqzVualzqpFQFuF36j55vWbAjmcnTScotxpi+Se70ma
MWiBKwdc328ZpI9EjPAS6zg3fcqAjzGPqriY5D3wnWtkxcHvCFTbMkMoE5T3mOKx
aIAJZq3d1zJiAZgYBMV5JDEh+W6lUES0BBYA0xOZrgyTByj79CH50isKIposMtA+
lDj9fIciYykb5neV+bCcggYSPDyFzA4MCyrgARrEtOv2SBSkfDpoA56dlhJ4TbM2
vZQVZdxAHWEfBH+LNPiOBJ2PcB92vnu1nQaEKauTDds0kakyrxj1S5EuteBDSqDz
XMMID+9IvnB32BclQKM+Q0KJMYeQLiZR7Im4ACyYlDS7pxsYFm8WePlVuf37PHRM
UmnqKYPz6Yf1nM6ivJSzBS3bjYITnyV2Ho2VL1zWBx7oZ23IMaLC96CZ+SPbh69w
aa394Bz2X9yHShnMZmcge9WxbeflXhT3Dup95cerhqAl6qZHRH9WEvqDII3mX8TL
NdNktabNeH/7pCDxkY9TeoX1RBJRlva8ZcIf/8XqqlIm3IilWFPdExJTFxbFHyPX
0N3UypdTV0n4mjXjCoTezPn8YURiUUvK+JhAcLfCTHYdMrnBOKr5UgcZUT2isgSf
wXCpfhCgkDS8/nD5MTuyg5eCTfaaTP10D9SRRa6DX/GBuh4q2eloDWHo/qW92FMc
o36gWhjDGFUf97YwzStUvW1auP/Vhui03or5grk8wQIMeaR/cs7TM8SAUJarT3iC
ihla5etc+bNKohkE6sZBW6hLQCJ1jzQOW627TSLZpHeroEKABYOIVrka+V0MybC7
OBCC37EreW3sKbTzsPsnmPuzdsFVsovlFeQ6LXnEPTacbxUxky9PGNTAeHMdk+1G
ck8Gajy4EbJWomL0b6yjCCfk+SfeAKwe480pZUOCyuJJtbh0NlorjrU6/jcYu2Sq
uhvQ/GmrQYYEIn9/NoQvnGvG8/L+Tv4nIa8PpnlMGFy6l6dPoVbHP58t33UcKbqw
bDFxSSYmDs94rxkuFWWWCh6zjp3h1xOSH4dPZrWApfVZr/2+tmQXnHcEOjWlkGq/
LUN165ZZ+mZ4XvrFw2XzFNcTY2LUusSCkGQKY0zCdCRLYL1sWdDPi161QlEaND/6
UZuZxi96l3XYYUzdSC1jKHN4QwPm9bRFb2KlKCNreb99f+f/kV20pMz5nRwRaEg+
G61mYwFhsdWFEkHXrij8yzJTnRnE90dqw0pIuQCyalx2RBysArINEev1nztPuybs
wirtjClxwKKh3tl2sWc8/icgve0gxuxSD6x1Pi5XiJfLb3Gk0dcf2Wu8zI4Ugddj
giZcHAvea0/Zp3cAbsadtGtn9ZQAzho7c0EQDPQIeDh5huqjrrrHmlcwyM5oxUZ/
NpzQKUU9VIoarTXwjFEaBrFZCaRYA5Fjq+NJXVul3ZfpfsEIFanQZ5hv5mXxnZh2
Pd2GDgybpvkxIghpeFJRmhmr7KUdwrsNUE7SnRPzHbLNFnjj0NgUDRQ9T7M9jAla
Naj8qWOgxbW9IjpyAlPCWHqEIdvJQzAoGg3Q5vMB79A4njJY8mp+4ZnGTUtqZ1lC
TTNjJIzw8Fz2XfKbOx4PpFOB+rpnamsrGBLXGtMscODgBozyRQ5bpbysxHFX9qVb
W5mf2gBaWK8/Kb0KpK7gVikrW2xNWnn0Rm3AoPKZXcMD5uigAr9pISWXPd+OPWaT
In31fajunI8MUBapJ3B795KbmP4RNVgYx/XhFisNsmJFgjV/NFAseWa3iT53YZsA
C4Jj6A5+g/WWUZKvXCM2RYC8RiE/bO38PHvS6z+BJ4yjeHR9uScexd7xVO595jiD
CrheMjS8nft9K8CUG5WDcXhY8bC2Uy9l/owFjTwAY7Z2PFR6wjpexPbxzURbys30
zXCPkl/VgkLIXHx4RGP5tp1gUNs7oN2zBC05KxAa6kp7oqJ2tgBjAfZjoBQsIFzR
oQ/aWqcTf+g9S7TaJ7d3JpBGwzOf5jN6xC9fBwtfTcwSji5JH/x76DJD0BCcqk81
Hc4NXIGiCbrOiuYr5pYFKQXWIYLyYNhqsa0MjsA2Mtxfbnx9M8qS4DQ2jNs5wMAH
IKemd18ZF57KaGRKDq6OkdYNIkBAXmKyKP0mEQoBbmQf3jfQbywXRGnaJU/TgVgb
vaPjpdDRc8OV/uImYZLRJRaA9YrkSNIqfPwdSGAfxSekJtpOu3ea69pIcpJD+9fe
eR0goWgOkjDPjAnK8J84zpSjye0LgR3ytYHtmhCJ3Mi/tyJN3WZIEhr6VCJZrOSi
xdMtE86L4XRGwntcbEowVA0xrF5MukeVgasNgOuGK0RHo2OYlSx0IJhS6xuZ/MlA
XnXxRwlDNPW+NlTrEMP54f5HH4dOMlNKgxbR3yE6V3GBrrQOjkeQYmZ4X/PbGFWU
A+G0dRamZ6PT+aGS0rKuQy/dG81SDIJDUETghblg0M0xCdj4dwvLM4aGmlkGzbTV
vNpTrZ8AS7OqST+WvxRivQycHU+uHLyIMt1wzAg46ssE/x/XXmc4Cf8IWHa9LKLF
Y4DJWM9Xfgc+/XfV1mLpTkxBaCKaGV27ALaaFCU5kjOPPwgNkLRhEqb5gyHgpgJ7
cDrPaJ+KeIPjyBIE913Huk1cK6vka4Cs/Uv89NPn5wsfyQhZs5lbopebBLmjVSKF
W751wOUL4ianBeZL240TDltRVh143lss/DC65j0+d10A1nUVgPtzR0bAhq2f3zQb
aA2yXhOadvz4woAxkxlsic8arcdpzE2SLs/jBppgZcAG6SFJbjucON/3iaQEz0Ix
C5slwTzc2GZbWPKYRZ0l6EyGkC3zg4uPfrOfRpRKScFMnS4dMMggiaz2Sr6lBOp9
5Sz/v98PjyTKHr/EJmtIN/+j+C1IEiYwFiX/drZ/Pr0CNQT+S9/S84uCuZywbFqB
yL6dvwW/ksIM2q8wjK8gWpd4BfaZJuch8nUJxLzsWeIbbGiltCU0HR3icyX+/e2p
LqQegylzbdTAnowjGil77nsz5Dtdkn9P2z4DT2ELuJP+XxVWxIl9eBL9OqqHQEnt
O5qMw1NP6jEGGbvR5ueE1Qci1iRxq+Yo4BHm/4pT2wGU64X7lxD7GL1mkiTCsYjv
9AkVrdcddBV1N9HdTJErdYcn32IRwrsSgAI480YUqV4RFGW1EjwHMJUAo+xfDshz
yvhve73Az6F98VvgKJhaOcYTkose/0v9tnvaEFxHX+TopB+MTYW25GAPt9XsK+zP
3Upu60+4K3wXtCf8l4fyIQWftCjZ/qqvfId4E1prUnDE5Q2cCXG/HVEAPStcFIM6
2o5noumR3tdgw6pAwi4+aNt5XEZldw6xdNVEoqQn1BVxakFGBaxZQn5yNpGwasBy
v7Df64tYlz6WRbD2SLqE3WHUKAQ2c3XITSc3+TcTxUhLnLf1gMShc9K4nmyZcqzA
nmijYa23FQwPqmP92BXw8Q==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UzKty/iEhkc6/VxXGZ9UuxTVGhWJ2BGtcxXAaB8GUTEoXY4H00nu5jPeM93j0vcS
EEDx3EQNt34RdDOIbLqjv3vzXE5snxfvef400YT4sMKEK9avDhiDrqOc8g85BZzs
0RuzKLZRuGxwC0/ezV3EIgipqrXOyZapSqjER+V4P+S8kei1n4+WZKST/ET4Z/l1
h3jYDS0Ca7peXOk6/FqnjZbyVNQcK98er3tTpkQyX123gQPQK1yDN5x7DW4tAX48
MnMBDh4solA2GX8r4DAs0qT0nSCKfmFBrc2QUGJK2GShylMJBF40PnKRKU8M934v
8kFZvajWm9VUjcuxIftQOw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9456 )
`pragma protect data_block
3JMuon1ylUFMwyUynoUgE+Jf9eK8iBMfSddSq0LOb1vK4cIgOYTBkeZ8E/AlTFO5
wM/VgB4octcrldaVSVpXauX4xfQ+iGojIEWokEScOMs6gVNSUGOChyNWg41up2IF
DnjUWdBeQKkyKFIf1suwy6gQxytyKIB2Y5w/LHFk80g0vm4qchzHsJY0JHPbDjdM
Aq7gyh0HKiNAL0mFY53AaDBzRmlNncDbiIo4n5XDROl22JhwJ0j+O0/6Nqrzdsu+
iQqpr57ap9W1npZWYO5oJnjhJLZrqZQC3n7nEb7TgKrMRgakxeApqLQ5XTWz/LWv
ZW9vHSbN0y4r/M1PH8+/8RH8eairyFTCOhbpY4Ou1lhn68J83JxqdO2c1eDSjmkc
AGjStcUpNSwg1z1HFSg+kDDSPC17xINpmXBHZIrZT1OWWclwddlbKc4ScSb5TXjl
hHP9ReyUnd0qM8WmgMKkRKEutYWgFULkbD0cXfkb6bX1GJ4ro+ILNkxpPtLPyvRd
6WkLGeNPDZASfYisPNwn1Lfte2wdo+eD/QA4yXppcyZQL/T9P7pYaIghb0K55rVR
Q41fmBLPeu3wXq4HlEHTa6nZQzSEYH6Y7WPD7IDMwDSfje+xU7/5OgYWD89Jnw0n
xNGs35x2NRTU53R62WiKzdAbUQo3WSc2EmuPmUYAeUrThxDPJ11P+z2BBZt3FOFa
dWEIfBVgR/wFRuXO1PZED0HQ998Zvns9cbg3Nv7QmUJjP7a+uTvwlVbtFGd8wTiL
bU/d94uh8QL2ZWW5XZYNQvWKdldlQN80bgAHywLJlmhq0kJXwj3cioTpPGEhZKNC
aTvUHu7XiMF/si0jgVsa8oUWgcRagO87wM68dUi46DNZCvmbIxhpwJk4UvdiqZcD
KLlV+8A8XrMVkchhBxi196XTizz0E6d2TzMjNC6jpR8NKNVz1iPL+flXMRdZCk0V
0U1f3kf+K3pAPMpZg/oHG9hKauu2JYV3HOO1VrsdtVKaubhl2fltu73dGG+hHKlQ
Y0WmBbJtuEF2lo44nZX50rhsQrhoQ1vOIKP5vgg9XA0bmti2UDDI6AIlMdCAKxwL
OnCvs98ni+l00cQ3HuPpbstBImutiGQquiQDlBPG2nyNntZdIws4pFFVku6N9QKD
d5QmPmA7WoU9QfKQmPzo6m80ZCZgkH9hPglv/QTH3mDo03OIxL5YocdR/3sY7ZXA
Y4yIzFiEPv6bLGM2OtyWAtqmu8kzem0ol/2wyRs1DuSKCmhAiHVSkgSa5hYmyZRJ
HLgyEgVf9V+KYC/95jev8VLFzU4vXS1qvZaKeBDw7hJ0f5ZJvRetNVColQNrz4Sl
6ySiLsiBrAyYUMfw7ngtrFUKANWN/73L9x2nzXNyaLM/4EcRVHuLVgNhmFokz7Yp
KSVC198m2qgZ/Tb0DbhME6SR7HnF+TzeIZAdhEJssgmOUZK8ApadEYck6riOTupi
Y52q21JcQp+0VgJWN/ykmeJupwumrE0hRmoaUoJExPNINDnU92vlqtiW9cGh1WhE
zcFKq1hUngfGdGH5PpeaURv7YnZYhrdL6Igbgvhw4m8mdz0mFrOW+yRvEnsfUDhx
gd/EtVr98GyE8iN/b/YkfA67PsGCt+3roTRb4dwcqoxIvusSOlLq3aQ7NsFRTLq2
WczcKJ/uGNwaWofsQ24GiiJQJfAUtADgZtJlQcvlaL3v8OVP3XaZq3g9+kO/mCdE
ZtcXSBZv2p9PQ5e/pDGxE8HZZ7+G3Bd4Kl3G8m1SscbYC8ZERwNHsM9pILWEZEY4
ygeXFO2MkJG+TNUjwyzsOrXt1aIeuG0hm6GT5ddPsTvqH9XUjqWOiNFXq/PSt+Aj
5eUWCcdsejSz67OvapJW33MP1/Dg4NNXlPPOJvFy9eZU1iJDI6Jee1Mag6PNM4m3
FhrX6jtCM929mkpruVS0AVIWc3atyD3Wz6mf/9nxgPJltmMgqDu3gzrR1OqFa8bc
Ct34wSm+ZsMKRygP7hV39JrwXVH0wDouvSLaAMdDbbpXRXbIQ/kbzXiFLAjqFMJN
7HwBypAlZf00LhqOpg3xKmGW9SLBoNi10NBd5mOm2t3tXEZUtSRpZx7yOP4XEp0N
ZDUr/1yP7QIFVZjL0BJQSkaccBu8Z4DxCYG5WzHvaz/NWdQhyEKylW+b2AAtxPoO
udyjpCFICLyFzygOJp5sOv/hGD+YDm4NIZ8af0sO73fCdjPh3QHZdG9hHERRc3sR
xjqaXlIn9Otkru48bKSd4OXStlQv/glcHo0JtWXwFjPiNC36B9/Dm07EcIUxj7+V
PQXFS8DTiGzT4tVnkkb12GzMEmOkEQIFmCR9p/OEiLn5XGrVna4fyLwgkyWFZivg
s9Tpbn3tGBjV/3SF8o46xFPjdRpFN9C+qNPtpmhHmsJt7nA7sI9OWKHIm/tesGKZ
2uEPloDuUfNNHi1qmIt1Opmsr3O0kIa9rWItICxtLKvHyzqp6T2mlWBD4CBMucfN
zG3GD52oEbi/OfZGfQIgQd135mJMpgNPiWVdcbkS975AtDMx9quCwVg1kP5ovmLM
g11sBrIyx/roIXliV/qH7Iquk8aqQTpvmR7XcFOLG4fdkw/nW4Qs/Gc5L4ng8oEp
fIU2PrpXYuZqTWxhMXbT9hYecL0qsnwF7rYB6425Fq3fT8D7jciEqgvpzFg636gS
nZoU6DOBeTfEtD1dd03YZvUDzgnUgukHfRWMgGktgMJicmIl0FPqgvaAUNLBPAkz
HP3z6AQAqatgzX0/LCJ5w+NjhnHCKt+5HGwv7GTaOoy9eMR9SMpza9zBE1426l14
1Ajd0/8wbeVRYuSKsBLa+8SYSYa+xPQABYZ0SuHSnqsMKzGg5ePEbfdyMxpJhMEq
duDwi1YIzwyK1oG/VEWZyieJEQ9NRP0IVqB7mweFJuiEBmt8/n3Gz/bfl3h9UW3C
ub2SqJkK6FANE2MnpQXB59gLmd4lIR8o91nElpSM9UwD5Nx5In5u9oQ3ZngYjPpK
WXGe1+QD/j0gTxe6GnXDLHKmBuumBbSwVKwRPV5/q82pa13h64ZBo1JkL8/90RST
nb+LPx8n+B2l8MI164fBgYn4vboRusl1ndC3caZ5Qe/5uSUyOrEvj9fDT/QV5ic0
qNc6La0eDt4nQf24IIPhFdHCmPEzbe0qgqbgyah8sh3GbtcRjQoLbBiy38r/2KgS
IBIRpW2al/GvzLPuE1sWZKZvVn5cmjajhv2Lso3HOSdu2NCRyrqusXhGYvXAeFDL
iOoFCzff+jm84acxMRPjLXH2D4O+OJ+hHuvwy5Y3HkayvtBU9Zd+sAVIVD7TW8iW
2RycNnXBPaDz2vgZKImhRDad0r8kPnupG31HRwGLAX5A/S9TP0e+bhZiBT5BlT8d
cv7rWlbK6wyezM0Ba7YHT3A7Ri4YISo8BzABjxd3DFtP/ziPU6OiqeKeZ3V5Pm5D
jLpGHoCOfwKrZOSab4WEy4rsfvi4pgxKU0aG3kX0u7uCatk5FtNZokcA7Gq3sABw
gKkjcM2JmmK9OGDI1shiRLOGE8pKTrYzgByCIE9L67KP49VA0lFP9hJ311KAbWvk
vMzbJXPfMPsDwGrQnXqNxKSYJCSmuFI4egWgiPC4bK9PnhLka7EMbUuvA6se+5Jl
93goRqssJSJ0F13Sn+fY2jL9qP+tJVYIsGR2d5n8GulIHT7MCuERZk5qxakeqCPt
NhZXpvV9I688ioxoRz1fkgVrjB8YFiVTBtlvWWIwanB5F8vCZV46qiTt7iDbDtED
oTQjkf5N4lGZ/0kGSPrNP9Ce2VB1GhZOQjn2sGrXvgCzWOiFOTr2pPR2pnYEvrvP
kQpmYeI1rPyuWQi5ZVpAb8wI9i6fIe5Y11V2JGrj1e9JKSbq8BjTkKzYjIvkb5ut
CDYJUdob4NSDr5vEjSjrCbf9xV5+nZT+8lcYIgFtG/cP4QpuvPxW1xLtDOfyD0qR
WDvggT6UEJPE2p42BEaT7wwL2uko6gFhzyAQkhoD19VM6gTi1oZuxXJlR6bJq4kq
/x7iJNC3jKfTcKgkXw5IQxxXTnWOkqpOJ58e1bw6TdO35qLJnj4w7Y5TEYj2bGUO
Wb+sX1uQhUyQRrCSCBYxi6Ej4vzI7woPWteukOSqI6CbDBFKLKBzIywBf7Lex+yW
0VO/zW2IU3IqBMx+vg7dsu+lhUWI21E7bRunf2UjVxE9b6i8HjQa6wznZOzy7E/r
C8YrsXvpxn4IF6hCRDR1ysPXlmP+S8FgbZCvlIV2LNIszP9HcETKF5c3b3PPPNiC
p8eYschkbkSJaWes/rs/3Z9s8ndSH+DoAtQt3jV3KbkMh/ti6ymEGIcqdYYCuWUS
PKxsgS6bvi5jL89LL06ujDDdvPEPEzBFd8UVR1BYfsJxV2hMrGe8frQRVqu5DF8o
+aEZaj3VM1IZtaMBWqowhJhs02yNfiV7XX5VnGRL7QfhFKbKvNtcHQ6O+NFBsji4
TH3P2q5nzuzrUj61A2RtDP17m4eI9tHKAuv3I01R4Bz4AGix2sZtrEtaLa6UqgMu
n3ulcaBIHjlVtlWRomxS7y8JHpUUweoF8b7Sd31huDn6cxjLayaoAiEtYALtFvZs
H0Xv345Ra2hg2VhI94XIZoUgfKDnVsTZDjRNHwpr4fA3Te5z7krKmlNujeB1YH0y
bjffnwZpnxcmCQ8gHVALk+qkKaPP4VDf0ufmBU+5eGXN4aEtroH1NaQn/5Zh/C7B
EYv5dIHoQm1nBTUr487jsE4kxyOVjk2IfZrn05mFRprCRZeeubJPnN0IEyD1WgkZ
i7IrXLs4wvgWxBysWIiE0AIKomrUy4B9guuJnRdGd6Uj1cgxMgBhWdQ9vYi3wq99
7wS+3C0eLpDWC13ZO7UeeDmp3jnCo01nOPXK6fit7a+cyOg610B1xn0HcIMDXa1i
LK+2NaClc5megEXWBFIO1bgj3vom3EVLdAa0QvMHdLGBeoZJmaMdqWQl7ERLNvRY
JI+YpD/aMPrgoWr4Gxw3LpYVqHrDG6+0t/YCcqCfi7RofkEl7c/X7AJ2bwpb+2YN
OV6+rcVXYoUlPSJlejrw7AWQZXPIx7V60C0ac+l+AiW959UiFVEw1RC5sSDDCQjj
hUk4f5NDIKY3jTcfnUvNb11muFFMa4aSTRwF6GjRzI9GomKtbgiZmoOQeR99GA/Z
q2x8JGzFENCg/Sj1cX7xwHvR1cqexwW9vAAXaZ+/vYM999IPoI3wWwDdly6AQd3n
HX+xd//uvm9KyFcEVgbECFcnvdACI7+Ycu459nEBzjDjIu9M7iMpj1JApICXDqTZ
pGaRkXgVV6drU1ZCE7Px/JWGKp55e6UxDhffDZCB42sFU/QATtcABvAwqdMGOTPx
MYg2po3UVi0JVotFHnipmZOXb2+MNWUHuoj+iQq2bEQAIhWnOVcN5rICiUvvt4nj
NRXKhBWBqmegzNZEVd85eOLGilBx4sDYoGAJ6a/eLBIGwU2aRMFoDvf+81xdVRdX
wz2ztvWL+E1hMfbARBPr6d66kAeNvme7Cr0/FnMIrSTKgfzBOQ63crdCo5tHPhd2
blNxwQcC9GYJ9gMO9Mhn+nzYyNB08DXvMKse/97s1YpjBhV1Sjs5y0+VhnOWdz0H
fIm9e7kWZKgZlrcOI7sv9ry+8Z8981E8h46knWK8sRtj9wZkxAPzxC1x557qHK30
HBYGRVu33o/ocMcLP3MqyNMcBAMRH00NMV7SWSISzKESG04G78I2+SegkllLezNG
CN47SUanZzxSPRfXopHEgL2+VOkbK5a+jErZNlE7nqWdCBpGa6peUYfDh8CHZts6
7e+z4HIDWrvbV030eYSuyG4ECosa9QxM9OJ2NxBE5ElmDCZys6KXdK8dMmPfkufP
pBprDDP40aW7znKg3s40EITEckYV9jrQps8OyRCUfCSUzj3n/l+4Vk9SxPWjGU3Q
HvmEFQfvRyNcImKG4ncEBXBnilCVVo4uIVYz5dnSUGaU7T6H2AVZVRL2Zl0ZQilV
nKe2yknAgaNeoOiMmjrFjmpWtxxbba57LBzsB2Hbu/x8UFWT7bj/2qzemQCxykKC
/AKPwl381mTsO061TYxGLHLMd1IP8FxFykQZrWK7VBqcB1CLL0qSPgNf3qx2YrU/
htknkLuy9EayDEXdB86QikhW/vOwu987KJKvpCJmTirYn1ZR+zblhjDoQnpwWD9B
oxXijSL4b0pI+eIULd6Vw3mcGQh/T5V6HZ/+HhsUvfi7WudKShcCc33I3K7z2TzV
22bfvSTxpHrO2vXN+1KmRv3hj6vqa50N8o44wn6Gk4JD65Wyf4PhkhPs1E+sWzZG
CkHcgtUF9+IlRshKgU6ryhqXFWv7igHnkdp3N3ioaaFxLdYLYSlD/qSbj00fPRJy
7byNscFtJ+CG3z+yOMk4q/Ao+fOVd1VwcujBJLeWi9Nt0Z9Qu0es+HDgU5VdlAmh
JmnDn+69LFkCIfrtBYIHbC1dca782u0TLgr9tmy73AkAimqIOHDQTrUCcW+WHEbp
dTKJZr4hXD7ZqOfJMVd2BiuxK57YOfEDDBHqmpjolN8cqfy62ClSbQHA5W/57ZX9
Sf99vtNTygj1DfVOgy2k5a9CggI6rqUE5ATWS7NMoj6cR8tw2+CJW3UfGga9I514
8zRhcCEktWfObBEReEsqo8Vkdo3bz6ZIZ36nxvqqPXlG4VuUEpQun7bgo9zMJdqJ
WfWmbxUduViGp4qaoGs07RUSiNRXFnG81C/CEGKllAFwaExvl65upWHXxS5RAyJT
R6/NSsUr+ZXokPSN4QsZd9SpfIyDcTnSWP3gdcRvQoSGvCik1g/IBerXNkyUNJI6
Wnund0paKsUMLY/KcU+sFkKIMC+4o2unHaWbW3PJz2+ce4u2eGTQPmudLlWABSXJ
gMXkGflkmDmaNcUhUkY1aB4BXfuOMpc2fePJEAp+t5S2uE9r+fU+Ge/ZVI4oyQHZ
nKllLXpmz87mXY/c8yb+l0aTy0924UMhEKlWiZ/zyJKrPxreUua8pAlcS4k4WPD0
bvkV34wJP8tXGTJiQSGfhecIjeGXW2D3CsDO7pghwOJxNiH5BFxqMsPrz7LJXX4t
XXx63tQJDBXbEzO5UDaYz+k7NBWKbwS0uWU0+vlz3bbd+/JGqXVN5cN9XWvuzN4F
xqZ1GV91dudjpU2L9oAHU0ylbAG8ZoWzDGi0ZUKL2KTFyH3YSHBxhQBZm0hMIqZL
PswZMdeooXTVwp4S2IlB358KDQzeZt9JN7MrcvqS7sfZMF7CjAyEX86K8Q9jzWc7
YVlpTX+Fy/scVWcIzOCafZ6nXtLGG8phK7tylPkgSHWHCslz7ZvyCyUtD51TL2Dt
MHLzZ8hSZAK1zk744ekv82E5DjQ+Pz9r4QNfwQANmBPCe2EEc9AvY21yA862LQXk
QSNSPe2SSHM3NUISHL932XLkJgdwBd7ouryEUfs5A1Hidrabwd3KrhNqbQmkGCcx
MP/sGjb6lgHbYKqxYfgBnF90DR61UlKDMvV0ts1ydIY73LJ7Fz1bppspNxbHmeAs
xPaVCG1gr7FuBMl145c4TflVBTTkJ/K/XtEZg0qpWQRwModSmVAjUffETeJQ4GqU
Y5ELMRbn6Me1/hMip8XV6WTwN9g3ANwiiTrB3v8G+SVWYUQ/1G2iMZ1yVkarfeOt
DBkuw3j4131gO6zxNDzhU2ZEzgZGj843ToDPXF1zfCFlCehmNwVXzrQD2fZVX0W8
DNCdz8fcTX8KqeVZpHhDFoTDySJx0k+HWS9m9beEFYg74ld26SoDBm5CTnKPa0Tz
EaYX+ZgRIQRnk+b6+AKktE4Usupj1AJVO+99cmxzwIo24Y8aN4wyQT+FVB24EaPs
IOmW+Gh6Teb+Ejyv0WNj1ObzEartekrOxAhBSdAbvFo0W0eSTeU+gFrbgPT5iB1k
SSDynD0Rxi5oIR77m5pQ/Uo5hYhlvrGwDc0USdFoZAKVu2UwKkOClFM+OEiXiMmY
5BsoxjLFMsMMIfaJCeFZBNZuJmlR3RzTPZ8XLsrNjLoYgyHhUdfJA8sBIXyRh8C/
cGJX+dQevzv4M1qQ5kxU6tWQ3takgpbM80h9Nf+GjcIO2SShb6SufpI89iV+F8Yu
f2UQIkHSZkn2CkBX7sxzadvhPLziSGX6UpH3zoR85WP0bAKFidTqIJD1SnXOmyrF
SP4YJh43WIL+/zp7qGdriSz5LRYJJ6jR+OlMfAz3OlOuRR2IiMp8JZ6lWxMJqhh6
+adFRn38BK6x4iHRIFUw2QH+nW10CH8S02IP6SxZOinRGqmuI1pMEm+SPEoiw7A2
TaZQoMsuvvgMP/y0iuGieWqxTYQIRqhqXBILvSlNBEbcTCIqoZar5o0iXhQi9GR3
L8E+nnw6p5ShkC8xLD1VsIindODuz7qN4hiQOLMEPXoPIUXjya2zobnAC1piraJd
nXakNOInJtYiIQ7IpcD4YTGeP5hV3BqybRKhhVJ2cpHz1OLIQmIyVt+coFNmgPqV
bJ0UZB9FLdgWD2yFMa0741RAtB2KGmPxZCzYy3uXzGc4fHrjRf+g+zo+9hU0waJh
gX0+3AU60DvurAseRIhYpYbS5IPd6HACt054I1hciI6yGBgG2SkPgkSOcNBbxHfI
8e9fa71XQ1B5GvZ3l2a1Q2zGCUyJN9UthNaaE0t8xQav7mP7dB/i6+1OLJ2itCQ9
DTmJx0g3NVcfq4SsuJFMSzxnldcDAbbccHZou+apV2CXcRhm+g2CXasoplMLPIbO
+KUHJMtzUnkODKzRYLSM05DhHjmXUV6OsNNDIzITX38vlNuaPTVy0yGHxYaSu4sV
N3Dp0eyrsoH4U60f/Qv241GS67Pb8sbF8rTOcq5oB3+va/oZTIwHj7GzwRnxZylq
iH/JR9dSAC3cZlwzWgw50QqaRULxbRSyVlUAlEe3YEmeH2hujpPtSU8t4ww2lPya
fSnWmKMQtT4qng5vGB5Su9sRN4JWfLEjqJy1ZlON9l2neR4Bp97c3FZU+/UnfHGU
/8W7Cygx4LuZ073XpYE2ah10w+pnKyTGEmL0CGI2LIOHjZEdBSDeKstHlq5NszjV
TjdmIXBNxYMuxqS1lchQ4l7y0b5s4udjaglMadW3xLd3PTPl3Matfm/RtDa+5lNb
XGMOVDDp0lITRvLLyAi77VfVlxUOPrB9zqgBMUThoMhAHAs0ti9Q1RFGXgwUQuY/
TCBWRzKy3eSzcXa0YXPFjqJLerrC3fiwDhBuJOOhUbPXjuAoJCbgctXr+SKUKEmX
h86ZUe0ThIINFHluRZusQCZOY+HB4T/jGzLfe6kSPVSX8I8V4GHAWkTiNCb6bJkB
ewwJlqSHykEQqgr3cHvpeaXFCwBe0KFxv3SwK1JAg85Rvhaq+EgnN+BlPa//zt3M
WqXd5JIvm5f1p6aagaSqg4CFwA96PwYxiVOirlMchK4AqHWrXMygyinE4rImy4uL
GXL1tyNkZTlcX1bS7SZa59rj8qKs+eMLjnSH0yj1ARVS4FiZBhuV5xvZ8z4moKIu
9etEFiGfx+DrEdO7hVqlP07LZGjDpm2LEqNiv5H0nb396XUxKxkONJnTgAjzJTUp
MWuA03SlI8G9bfIPzR4zwKVao3V8+tazUZJokcqlOBhJb68QtHDq3Uob5L55sxuC
JG1cQM6+71ZTFVQcjqfKI5/rMXRXHMYJekhjnZreKem1sAw4gXU8WPx0mN32bfuo
cCplLJF6qfmhqHm7WmWDTYsIg1bP41q1RZOgOyKDbADSXok+64MUcSwSRCRGLQqp
t4ylPnKMWhJtK2H0GdGpONgcK32bf6GAix0yrKsdOdFkibeXYn3eKa4FBbhsawRY
AFcaw43HONGXqfGAp8HoQdTudd+6MALDXxl4yehjUqV8UJwtTRhAjLljAsqypTym
3hnzF7psxqKYiHS2GMjkf1A2fP+KcyM5COMcH/a6ap5Y/mjVpka8USsO1lRFnoMj
EWXTcwy+DzFm/afGomqQtLl+N0Q5BTmiuVkOK7URD3vnsg3gNbAaJ7EA52QC8mCy
URAhmvBaVgEP2wV8LG/zIodiqX82lVYXUAnOR15aUEI/6I05IWzRsMg8PWubFrAM
gUTNQmw/9Sd743YgQqe7mPQADeoXnZB1sODbtOblPeg0LsKkwIqxI8st0tRvBF8t
rt18mRBpVOUE2B6YCkT+6Jzr6KJeS8MLj6Z2Ab+VExowBDD55rcCYuwVmWhhk+IR
VHcSil+CQVqkK9zhKjKomQSV0KXvQc+6Ec4lIP6GaYPreB4mP7JgPg7qFtZvAS2p
EKv26DamfrNBAVLAiF931lz9Gl1Xb7IpfnsDMXcJdi0/SR79lTVjFHp3wjxQtDKu
E2entoBZiYNVa/kZi522ekhvSOOqK09Kpa5+7Vo9GMnxEPW4aYqF3hh++GIvJ8j6
Lpfyj43/TiXidjm63Xqn9nL8o1tOiEsnPot+dheSFJGH1UiDF4aj62b1RDcVlOUp
lzqHhiledNNFFvMj3aeUBtOs+eBW24ecBW8hytiI2SJZsTKvm61+xuP1mehgXhSE
HVyKNJkFnfnQvLPFiDoGJcBY5KumQ/XXyGkPb9R6tngtSvRlKt1FIl/LpuxX78jL
siE90+/FKzdOjklPBL72aFQTKfzdkxeufOYKrHYTKDs9HSH3O5ijJp9B6OVlPuoZ
oemZDXhhuoAPUcxjEiYxRa29I95FzlPOAe2fsZcF8NWfBBzunqAyMfP5cvGDFrKV
cOsisFh0awo0T8gCPxGmPpYkiJBqbc9w8erjiz58hy+qC6eFPG6BAi2jq8E2xG1E
HXeThgA4tiiSW5MKjEz/PG8w60KFIDCUvsbfT/zHSCAYnOIW54bo+CzqWE1FtZt8
pmtUsz9Y9QrsdcbbST4eaJmgvF0g3RmLf/nfxEbopmF5oaFlWG0HqT4J2BtSPPkS
1KMXzilMGaBnTBWy5yr0UTN+WSjotQoySvkrqEpQ89zRKg0X3NUUitij7fUS25m1
CNpyHoo/j2lNd5FYPvii5VRZDQWAe29vcStYV8BXxcz1akpt0IbIy5AhPTfZWYYX
XQKRCcPs02OzYndwyZU9jZxOepF2hnlDmxUj6diXUOA4vB1dVNOe24SZatiVsIG6
NFDXA8DJyA9p7WbGDaUkgHV38oH/2Q43Z4KIj89n/s8SwA1lqarI4NMxEx61HZpd
Oc74hWdmjTwxJY2bVHTUkVe7XigCTAV/Xsn5fB5pj5ViZ7YQJXhqmal2t97L/TzN
tonQ4TdYD+v8T7dNfSfRny65nUB31EbDbSZ9/EEDmgzJCscRLQsaMWx8amu+XPwz
EvVXurgK+97iIrrlCpfsIsGGlffQoNTCrCQ/sMkNP4Hy/icX0nrpE9+74Yii1P6o
LJg2Q2zZiZxJn+61wf8sp5wLk0YZ+nvEjOP4PMIDINT38CohZaNOUp7EeQNAJtsg
a1GUAVQsbwRW8kxJsX5LkgJiC46uTrGk1E0tbwbYGdeP/1FElVA81yL212GrWgI6
gZ9vtuzdxOmlAszFXy7ECJHPlUVbLF8q66eVsPHsMPaVqc5e3c4PfiDvjua9sr2E
rcYBHaFpLF1wLF/ga4OmCHL+fyZBsjCnAZfT+zB5TBo/ng8Whb0K9dH+APDyAzkN
zCwwPbzIWRBVH/tY5faM1YEpIVtUM25YvBBxwDOKHUp79sIp47mpE6+K4n4fqv2L
Uzjs81xc4vGK/A2pCGdxoQC9/1twD/RXOcCZFzeIYd1Vyh2jpA1P5al+d1o2Llkf
Df8kbz7peiVJQ2z4vRhOIOeDvKTq/RLE1LWk/yAxojNvWwKc4KGF/Li6Mbx6v27F
GLJr71hjxmdVgvzJrXawddSa3thoeE6KHHCOjsl8v5gFadpHH9Hg/a1ndgDHa3NM
/vzRwFFeORqecmIULfSrPitss3auey7qSBL9LOX1tx7EEaP5Lt51GT+wq04m9VVa
aUDDhy1uBQF1qH2bPLXqmmhYVksst60vQFnvhCrGVhWlG1YIEsC6clSFGEINwV4k
15F3ynFmFQJtFP5r06Yb2yTx4yh6Ee2SAyww6HtMC8SQo4Wdz50HW3rkg5KhIKQ7
TQwE2mbJ3c5Xih9ngluHFiLBU4px5Ct/DQSKL3aG88cvZts+yihbo7Ik4T/y0X1U
mbENJMw9qee92kFr6kIvpZigQJH1qfevqPSPtyZNZ50yX0wsxTgoK9nG8JqM9IrU
uzZGW2mWEx3gXwLcZukObJEFrozXjuH1DxGVNixKRQvHIHowEB4IlTxpGYq9mcCO
zhvFdpxNI1Hh5z8riSKllFiAeJ/rh1f/fvGodOcX92KwxAKAmk3kzsQ1llKWWhRa
CNrUvqMk+kMhldlgIzSsRKws00zP4HJgtCLmMDlP69dEvijcJXxETAGfQrpfvUPp
smBsDHHn4DqQjiMQTzbweZNFdH6SeXoefZEVTsNwtR7dX/xcJtcl/jcEVL92hKaD
TvOejW9+/0UexQVtjJX02b0j2IYKzOO0xjcuR7OV9LBOlEZLIZw++XXV83CMQtEn
U5upu1qtzgDCJz9tGLCjFiJYhwBoOWeURhOcOCuQ/RapdwIqakMhg61rhz0NFqhl
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
fRaxoPgrF4fO+Kn/DjTIZ4YhaRqWh5A1TefdxEFwGK0KfAJlxSQgu8MfutoTIyQd
hAbwGjebLxN30f8UMhAXNexvTn4ypEXMv5ZAFaw4m+RYr7BiW+zcrQQyhcpxcoUo
K8UrB+zvcHPWPOfKs3hNOsVFfzas+z6YL1MMIh81S2xbTCLwUJKHAJ4dfHS/WIWE
6zgP90/pDXe1/Yqzr1hQ/n5jaRPxei7I3sl/2W0L3C3BM3wriPfS/r6sIEiLhd8l
183Nw/ugpyfT9Y9MeHzxk/3aK2JseTQdZGT7CPzhSaELB9Vvrla1LzgAzFj/fYFE
WH7UheR/q7oTMvMApxyNtA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2672 )
`pragma protect data_block
xlcKxggCwQ/sS0RVqdmE4U8hzZu9So99LdhH0g6zakvCslTqxIq1V2sdUJkP0kUk
MguO9rZDNWm+ih+5z4LiaJXWh/v2hDYPkFGaesdP6bSRJX4lkAEjMTW9EqxUQfBX
Ff9ZEag3Jz/TrmnFZjkHPS6RbfFE5MhZKe2yoDd65RyW28csE2kJMuvHT+cOd5jO
zBmM/MMb2EFKSRjRVHfeLKEwP0GLI/JzTi80+WScHmrJuV6562gpeUCYUAHMIbIl
mvgsu4r5DalvGkkmXXDUu3HLx7MliJ+2n0nKt/Fbi8LFzwPeuBa/4fd+dldQf1mS
dQJ+dBme2sOhGKQ0H3aiD2Pgt87oytgZ9WQzlaCQUnEqxUW5VHkd84jYBYJz7+Ue
wZxkiKL8ul6uFOeBh9HDFIMp28GJYmoBkSUergU5pONFrCnOrU0cP3IfIOl3TGEE
Qfc+gOMCwS0AdrqRmAO8RpX/ttswy/rFGEPQGogKvuOVAqiurchNcx3WqPwkKwxN
s5bO+I6bFAQxLK7YA2Ztn9loQiIlgk0iybCLCErC4mSM5VRj/3ZJd9JZx0fjFv1r
1fKV4JR/7Tw2NQqzNzVKTPvm3fKRtvR/4BjwU4nMBvDNHcmXV6Y4x/1g78d1LfDQ
4p/Iuxkhq3xcbx4k0xrqvKFewiAvv3oCLYNPnysKnDsz3PhXIJ5OReHyEg5YFqUx
kUyAfaS4UJ5WXbdJep2zrr40u0fqSTJS9f4+NXSUFAeyHkNe2F65FXhsPzcwsINI
4oN1dEyzqdvJ1eNqdf6skNe9WZWv6P6iulP1xJSQb6es2sXiG1ExN/drR2mBtkhm
Gt2LRoXnkr9qodwAdvSmhJt8C7mo8d3FcbceYHy4SJP2xCa8Dv2hGG0gLKI9lXKR
O8Yz1zms1qtE7bTd1vwv++ndC92GZCqeFM9LvJ1tZzH8PJ097vcP3NFP25Xu9jDm
pV+m9Xktm23K5dcUZIR6IFV5MyP/fJJOZM6mctAvU275hbXNfMuHJGiJoP4oxHhW
37z8X+XNEhHcKr1t9KzUJ8VciD+d3iYo1C2+Ac0eUMFNmM4kNYA/4s5VUERS7r7u
MRcMpwWiBvTmEo+sfrlOeuM2gPEmYq11H+gvlJ5mCNWr3LDFCZ7boo68HPf96ZjC
0vpMF+GBoxaxY5S1qax4cI5MBPOPK4OUwxvpq0Tpc0ejqYjgANuhLGho6RAvnhJb
AenO24pY84zV47kd8x3jEvZJtyLfyoubitDAcyNqSluFqggfyTu6SQ5MwD5Osnaf
+CWGkLfbU8b1cGmkaurpS9JtiHMcAZa+FCGfrFSRmkV//qX2PtffhXsh6LvEyhNO
q0uqcR1E40qvBJg7FjUxIDtlE7SSaWJyTJgRMYD8xReV8k20bSZAyd2QplWaksJV
33J/0x+1+IczKRot5MKd3kGCUpqGtTzJ2lwd1bEvHMwvKk/r1HW+u9n2LtmXzhDK
MS6qxSLpcfk1n+OACb8ZAvtTW3Wi+aH10BcfjfXd3YtP4CNJmax/JbQLzHu47D3+
KtDhA01poTlpsbqJOLMAvq4ENaDUg64kkVFZSR6owUiZH+2Llgd19vTGnCC1JvuL
IKRacq7EhSV23blGnUnE1issCF7JGtQtFGfFGcyGcfBkqJCjHvlC96Fd2APh3xqC
F795wfJwb5fiGZ0l/iBq0ZO8BwkUdwV6iNrr2gDFGEnaRx+9lM1vOd7kKJY4CvBz
hLwhTByJDPZlrvLLkQAMPaJlIZVayAwkgRSUCbNER6CU62EqnFADWDij0uhsQd0K
dDgL7ByXzT7o02GJ2BJYbWS7HhVCIL9hqkaLg54n+DziADsD/q+zlYEgBgXARH01
g4Zs6EHM4piuNv1aum9ja0K+RvmaQN1CNrEKGp2hVAs7hHDM5GN7jOruS4Iahg15
9jwJCIM8XYxvXE3FlRN8SsT7JZXFNAUYpxTnC5vi3EleCYWFpZ4y90v3fX6WoGwG
w80/4HNGgMOjkcuaEKDn1tdtTfuAM4rq4RYxuMZAaI+TgRch7Uh5+k/FL/BjjFrG
jc0oCXdn9LJ3HG8ZaGnmtIGrk7mjHatp+CVM05NvI3iwRsclwFwu/QeydCmyP8pY
bikES6aEnWl0b6qi08sra+9yDc29CP9AxSIFHVyG+Z7dylhN/4CUFsjgA50xWRRM
4iU3sFxv+ITuCPckn5u0H0XIeu9zR1ZMpjLtKz8JrPpDNi0evEjiExJervQg0aMk
PqWI7cFLYgFwp2o1+38qicY7qY6dSaSrGnbc/z8kUQc8KpGSCAX5V3IbHyBx+h9x
8Pj+rQVc9cvFxlpOLSe8qpSgHZON813YNXZ07HnfHgj0g4i2hmZ1u+Iuetau0HmE
qFr3qbfLxrxg2e0/hHmKWvelwN9A5t3qIZHvXoJQSP/qv3GZky1aZG6d6Ge42yZN
dekpeLNp53oS0VlYkk2doacyvXPO0WkSxbsUrf4PV8gv0o+kEK/Id+ITeXZ73mSj
Q7u4r3zBQiuvbxhmF0+IbmBOZLWVkh2NZ2dHHhgeH3QqtgLAYt/sAZFJPurIncq0
2AkUTRncyPUXpVDsMkRsgy6c1xReJaZ+pjYqPphICxaAjjOB18EP6VchHWnsfK+B
ucC341DhqklKqcIhXagiDXugs86TqhdA/0wK4+5e3+/MO9xmKOK6xSQPi4Pq0G7/
kxT+ivO2f3g8aBmVdnb8mCEDcf+tX+LGaWAoHNekbQ/nyH5bTNwBmEjnqw5uieKD
tJxELc/nMFYPY6YlOvz9FEXhNMjpHVjYqx8fvdI6J3431/hnGmDgMox3HKM6qsfr
4jcsW4P7UiC+GTUfgBKskqjhsJzfJiPSgb6IQqrKdxoE/cCEoh6UZ1C/QnNhhQFX
ziOnCJUJglnTy4y6zFyFkYJcDZ2qCDNg7ggUg8W6U0O7+JOX4mkrIWmJasWcAei1
PbhMatzpAIWq0sIALA7gOYH1MLZAC3iWpGXTNUcod4fqqa8e2t0mzDIAkGhlxHhx
/fKOdayTWp1IVIoI/umx2qiJfngxLxoPKxCTbXAvw4jl1dY8zoQioM9epE/VSmo3
8PovUa81n3G7CzVSywIkqPUVWBxwnB0muMP0QGzn+OTjsBgM8W0+WvpawanA/bkn
od/1EUQl7vDZH+ziJgpvj141wuAgKi+CviiUIkx1BQRwlvcFT99xlIYeAfuArk5N
4nfkDib6HCPUDP/KP24LF6uk5F4i+oN7A3WI7f9ngUL1UKlFT5v0it0xgtFmjU6V
G8YDG2cnA5QyBGlg+AERfZdDLBfa78bTMpogUVlDazhzTN+gvgTq+7v5hv/yt2T9
OgEEuJKrWRizfmy7LhxxGFgSZZoMCyI7jMrFQD2AcgeFBbO4iXGCyQZy9g1c4XU3
CPqo9vJxc+t5uQKvFexY4lvHS/+K9mBwpV1K8xt3HD10mXxzCs8Tidgtu8AvMrB9
uxm10rvCSYWOVWWhnB+zdoOg5OW0MtjkUGaBuubmamZaWV8ZWvfFHJyre43/r/qU
NONwxGWk2nb2T95bcAG10fBqza039IVDLmZzxoQVsGw=
`pragma protect end_protected

//pragma protect end
