//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2024 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = tinyml_accelerator
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Mon Jul 29 10:45:41 2024
// ***************************************************************************************

`define IP_UUID _0aa6c7c6224453eb5782dcbe16593dc9d52aa7c
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)

`include "defines.v"

module tinyml_accelerator #(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 6,
    parameter                       ADD_MODE                        = `ADD_MODE,
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,
    parameter                       MUL_MODE                        = `MUL_MODE,
    parameter                       FC_MODE                         = `FC_MODE,
    parameter                       LR_MODE                         = `LR_MODE,
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    //Convolution & Depthwise Convolution OP Parameter          
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,        
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,        
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,        
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    //FC OP Parameter         
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,  
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE      
)
(
//Global Signals
input                           clk,
input                           rstn,
//Custom Instruction
//--Command Interface
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
//--Response Interface
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
//DMA Master AXI4 Bus Interface
input                           m_axi_clk,
input                           m_axi_rstn,
//DMA Master AXI4 Write Bus Interface
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
//DMA Master AXI4 Read Bus Interface
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);

`IP_MODULE_NAME(tinyml_accelerator_int) #(
    .AXI_DW                          (AXI_DW),
    .OP_CNT                          (OP_CNT),
    .ADD_MODE                        (ADD_MODE),
    .MIN_MAX_MODE                    (MIN_MAX_MODE),
    .MUL_MODE                        (MUL_MODE),
    .FC_MODE                         (FC_MODE),
    .LR_MODE                         (LR_MODE),
    .TINYML_CACHE                    (TINYML_CACHE),
    .CACHE_DEPTH                     (CACHE_DEPTH),
    .CONV_DEPTHW_MODE                (CONV_DEPTHW_MODE),
    .CONV_DEPTHW_LITE_PARALLEL       (CONV_DEPTHW_LITE_PARALLEL),
    .CONV_DEPTHW_LITE_AW             (CONV_DEPTHW_LITE_AW),
    .CONV_DEPTHW_STD_IN_PARALLEL     (CONV_DEPTHW_STD_IN_PARALLEL),
    .CONV_DEPTHW_STD_OUT_PARALLEL    (CONV_DEPTHW_STD_OUT_PARALLEL),
    .CONV_DEPTHW_STD_OUT_CH_FIFO_A   (CONV_DEPTHW_STD_OUT_CH_FIFO_A),
    .CONV_DEPTHW_STD_FILTER_FIFO_A   (CONV_DEPTHW_STD_FILTER_FIFO_A),
    .CONV_DEPTHW_STD_CNT_DTH         (CONV_DEPTHW_STD_CNT_DTH),
    .FC_MAX_IN_NODE                  (FC_MAX_IN_NODE),
    .FC_MAX_OUT_NODE                 (FC_MAX_OUT_NODE)
) u_tinyml_accelerator_int (
    .clk(clk),
    .rstn(rstn),
    .cmd_valid(cmd_valid),
    .cmd_function_id(cmd_function_id),
    .cmd_inputs_0(cmd_inputs_0),
    .cmd_inputs_1(cmd_inputs_1),
    .cmd_ready(cmd_ready),
    .cmd_int(cmd_int),
    .rsp_valid(rsp_valid),
    .rsp_outputs_0(rsp_outputs_0),
    .rsp_ready(rsp_ready),
    .m_axi_clk(m_axi_clk),
    .m_axi_rstn(m_axi_rstn),
    .m_axi_awvalid(m_axi_awvalid),
    .m_axi_awaddr(m_axi_awaddr),
    .m_axi_awlen(m_axi_awlen),
    .m_axi_awsize(m_axi_awsize),
    .m_axi_awburst(m_axi_awburst),
    .m_axi_awprot(m_axi_awprot),
    .m_axi_awlock(m_axi_awlock),
    .m_axi_awcache(m_axi_awcache),
    .m_axi_awready(m_axi_awready),
    .m_axi_wdata(m_axi_wdata),
    .m_axi_wstrb(m_axi_wstrb),
    .m_axi_wlast(m_axi_wlast),
    .m_axi_wvalid(m_axi_wvalid),
    .m_axi_wready(m_axi_wready),
    .m_axi_bresp(m_axi_bresp),
    .m_axi_bvalid(m_axi_bvalid),
    .m_axi_bready(m_axi_bready),
    .m_axi_arvalid(m_axi_arvalid),
    .m_axi_araddr(m_axi_araddr),
    .m_axi_arlen(m_axi_arlen),
    .m_axi_arsize(m_axi_arsize),
    .m_axi_arburst(m_axi_arburst),
    .m_axi_arprot(m_axi_arprot),
    .m_axi_arlock(m_axi_arlock),
    .m_axi_arcache(m_axi_arcache),
    .m_axi_arready(m_axi_arready),
    .m_axi_rvalid(m_axi_rvalid),
    .m_axi_rdata(m_axi_rdata),
    .m_axi_rlast(m_axi_rlast),
    .m_axi_rresp(m_axi_rresp),
    .m_axi_rready(m_axi_rready)
);

endmodule

`include "defines.v"
`timescale 1 ns / 1 ns
module `IP_MODULE_NAME(tinyml_accelerator_int)#(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 6,
    parameter                       ADD_MODE                        = `ADD_MODE,          
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,      
    parameter                       MUL_MODE                        = `MUL_MODE,         
    parameter                       FC_MODE                         = `FC_MODE,           
    parameter                       LR_MODE                         = `LR_MODE,           
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE
)
(
input                           clk,
input                           rstn,
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
input                           m_axi_clk,
input                           m_axi_rstn,
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
j+jzIkMnpyMZd5dW+epx8rKjd0VmETa8SLFtf5s3aYqrQCXuFN4fPRfTaOv007mi
J11xdyLOxFHE+yrFHmbJRi+kSqEq4WRrdhey15Wzt9rX+iVzsYVsHnzynT2YwKoX
B4cc1wTE3cXiuKx4ST7ZejS6NZy/RnjgTn/9E1Wia3o9b2ZHiociAXipE1kUpVnq
YlBSFIMWbwpOXMJX2UCZdNBdotKAr9PV4cCF8ZD/bZRQ/mLxcIRDhvE6ReKY3giT
M/vrlOKIqGBSvKgFqDbW5O6PGQxQ4bId8xWPpCY48rPQ9VF2OE2nH10U4KRfCl1r
F0pIar0tYN8SQxAdTUpYuw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 59120 )
`pragma protect data_block
HucJdtI1toLQjHg6mqjnKEeiMLPdcRJP9+Pul/G4f9W/Jw+76icz1LxOsVgOvhdY
PNpSHXD2YrM4PA1k9GYvu1pLhO3vUH0dRYd4vLR343PnF3Kg5m0FCWxZsLWG3sDI
Bqb29VBQyXsBjOE7dpnTxCdiBzB4EQhlMXMBtzycXafAthRn8cKJkLzArgzQZf/7
8Y+ngM7VYpFnDCXJSO6q/fsgCbjKqnXTSZvpRenQS6h2r6JaerBAmQ/1Bcx2xj1V
zv6zR+/2T+Vm5KlnkUskNAXaqO3Q7SHiys8P23XOn/dk+sWKuaO1AaLTqIx2oIrq
f50y+bA42nuYIdURtbYrZy54GUX8xQ9LhYdEnnVeX3GoqvTjlBn0HXlMEHI/R0W4
+tkhzvr5t3F9FjlyV9AfCQYNvUZe6783Q8Tm/H3dYJyN3GSEgqQzSvXDocq6ZAwQ
18NGeMRTPD0Ricku9gpn9S55FhbOsqleYWLfFT4jHKlD3RiiDljJ7TX7Vhu3wk34
Q7q2xu2YMRfg74cTDN4DC9RMjCkcjSNEiHZ1lJss1E1Si6KOpMUI3x+4rfGqfenO
qv1EPpe4IrLBeHfVrk+zlH7qZiyKEK87/9SN4t5KTQPCDOSUFDYD7Sopkz92mz4C
mB0XxkrUlqiI1oYiUNq925ONVPXrC+EU8Q/LTYnsDbhs28QXa6FdEd+BmNH3Ch/M
O4WN1EueCugTH0Put5Pq7NyRY+0pfQKbimwrY4gbhFp3dSvrtLKbSIZm5HX005hZ
vf5OE8s01sb0qlw1vq2wn9ZJTLfoNQ3sWdNUIDSUZ/nLGaPv10r+75OVj1ktpjmJ
SeyREd8fK/tVmrg8wmjOLvUF+EWU2GWeN861HrXQrpgDQfK2DKqMKjSwlzCOWVKE
MEguc0RR/e7DT9BJYIIMZiv4I5XmUj2XXvsjTz/B3/ucMCp0UTWLmRKjBE+/EpGc
vLWloGQdaOtt65iIs0aZr54e7GAUdAqWJnlYpHo9O8LW2qj05E0uzbZxnBA7FVQ7
9QddUE4d0fz/v24dJD5vrWvlTpCIh0YTDCChaMKli0EWI7pzKWiuv/6z1vfiVK/e
5WJNPc/vveLS8A0JTiXU9YdiXzwYsEmiQaGbgtmv3lkHJikaTL60jHABlS4/7M0Y
FZ0+KPOrHOQiepPBImnNI4r24BHERNyUy4QARwI3bHuiAT1iPJT+b6VI2ATGFxI4
LTACWqEvqjne+xi/9amouO9ldg1sYOGPzy2plaCO1IBdnJmX9V8EszQCZeKgeWW1
fZOICDFj3RkEnONQYaQBowoJdTXCsP96snGLIyoaS0WshGjyjRJm86hiCtguZ0kN
QeLhX/6PZ/34edYrkwIWydBPZuurw8ppcAhHheXKyl76TYYS7bitjI5w53RrNv5U
bNVOJWGBDDha4g2VqJ8bUMK7DW17xOB8izTfQw6ytovn/YwEBH4qpPH8AUNkVyMa
jzP3jUlLmdgFoFYubV0sQ4xEvr8Ew+9YcOXQZU3jYXlbzpOq/iIYXQtkIlHGuo2j
6pQPF/3yJmRds9MiBMO+vL5pnUEX0P9IYTKG9lJsyj4XY4Iae3TlScJk9awPcLZk
JQPA2IoIQibZofM5vuxXXR0Zev6upaewNyu7ZJXMTl7aVcLnIPG2Uy0vVzjgsmmj
+tc7friQYCM9nMQkc5mRqUsl1vwr0qRkfculWT+IsaoyRwUi5KDwkuTVqwBZpoDF
q4zYj6654MBdo48t7Qi4dYV5FXKUYiuMemgCjlCWBTeBRtVCAI5utFoQWMcu/gGz
luVXurmqs89A4BtgO0TgEU8cJ3xve79z0LVfrlXqZt4G9pqezeNmI6BZQLAKqbAQ
XaD2v0GnIGG5ZXZcT/V8JMyn9RCvF5tZaUMM/P1N3OQsmzw9iyC/CipI/9qP6OEg
9Wob8A7CyZlEtvupWEVtPdGH0K4zHPNliYGM9CogDgZ1qArUotuxwpDtC9emfwma
+L6dzg3hqP7HcaB+Zrd+UAndByVQjKir7F4SJaT2JlVG5qbhJxzE3Z1FtHQbyG3s
GYN8TaStppqkNh7cq6c4kAj+mCJx/Hr0J7KCNwVSNXocA3QZwVOAwqgaqURPIGBb
MT86C3OkuX6Ek6LldV5tNykryp0NFccrZY7+cizI7viCpms58kB2Vwzbyp2vm/bz
deSo+jtR1LogpZ47EBsOMSBCykfun2f0MCunoE8dx9TKH7qEqkKFPWZ3esfKRkqS
pDby/ckj+ogA5gU798q0W1He/Gl6ybj8dMWEqpth4/rBUEMed7+8P0bLQUvmvVjB
db7PpCT64Dl7EnU+CJjIr95FW30DJaa28YdQvvmvREydlutln4encuYMyX8cD1fO
0ZsbjOiOQeeqCZdvAhoQUdYtW8pp0P0c85UK0coZ307pSrPz33fwoptAq0NBgl1i
r+k5CDz/6+MVsXdX5ZuV7LL3PajCa7Tq3J3M1TaFA7/mp2PDrjlFKcFApf6oSSVt
HCBGVApZsiEkJ1eooQg4ah17y/NAHJgZYNh3ZozpanJosnQl6mgfCzUgopt2t6Bi
+QOhcyZhbrVHoBFrCQxQiR1VAp1GmiFOKkvL7jgctprJFVvDIJJFXsZyJCFcafuS
V91EZY02aqgSfh3YitYil1wqevsb1pDZBsP90syjooOWtUM+WrOdrzDheMtf0Gwz
wcCf7G32cNSVYlbBeMLvLieO95pexx0t5W4yOBe6yWhU2yWCxWDeHSDEUo4i09l0
G2C1OM/21B+B8RL6dCzaX1nuzMBrHqbWGA6FFyVxxwEolvooVUFN/MR3Z3VNXch9
3bGr1N2Ek0kCsCN7ryOmicBh46DqNEmqP/uqZddGWmC7e4hCSD7VUrrCQ8NccvgE
eEPDGxakxuB4+n2rK/tw/z7c9zwDufhDsueIcjjjoYTso6z3XWwh9UddKt6ORWHL
TUufdOT1ypdoG+URgUIs1b3n+zQcdwmchadc/NIlwo/uOCGCvqnRxsy3vAmzrXkv
6yrCL0USu4J+wR31TFO2DCDUIJkGE+Mt97vieBS7o0pEUE13lhPG6PkPEPciTw3u
j6UctBOX8QDZ3uIATkmjR2H2uX1SUcI3fmOzTuUL4yeunbMh9EUT/jnPxJwQWtKD
oiozJaqDKFUuAQta40P9wUK2LcZEoPq/KYPopoIBSiANQuQ84aap4QPmmvCG6pPY
/nyAK1Q4uCn3iOIcwDjLoKjbK0+iLFto5Ie4hF8DSVI39kuD8dXoltlabZFu2ZgC
QxVzzVbtWxa8KXMifvtT4PacYUADcqN5wGLKKPK7YO2zPwQUR6SDs/onIJjcb+B4
O+8fAIRF7bmIwoTgY4oN7inBmB7Go/QoWZ1nlILjXkWqRL5iqMFpXQBrvd2DnWPI
3uy0+Uraaau/1lRQp/CGyrO2RrFBu6U5VxwbEREdXFZ6E8ct+TDauyvpsRZ1f65G
14v83GzVNg/DNqebs2Pdp9TIYpaGZidFH0/F8FPN0TdNYWK8njz3ye8mw6mx6F4B
Q9FJYOCEgwcoPgwpBDkGBagvaqz1zE2s/PSeKV1m6jucQuC41FM0Pz8rOKZWy1ZN
+fBuAyqZIu4XoO3NHq3l8GaRAMPZhPynvfYGQKHqC4gs2UMFS6+qw7qxNz2AiP7W
SIwWcqUoGXiIHJc5aTQ9sJBpehhAyqeSZKP4o8dDhfHimmN8TQ63ogfmnkD2YWIW
KsSGGWPDybtxxrJWKUPJWn8PHOSHBkOFN2xbG8Esr0f+CNIf9fRA2NeCTcrOMrIZ
VnoPNI35tBEWbkymHwEG93ZZtTmMPFhueWSj6XtaLuDm1Hn/qoKGalONftX0RDO+
KKAvXN5Whwev6L6jYEBvOAnuVRA0Zcaz4sgVbvwFF/21SJQIuqTcYDrdIldWp5tz
YBxAR2cmnvY4RbuXo3xbFk38iFpZ37STCiKHup0cLLpTL//rUd1krxHTLCxw7EyK
Ngl+Z4RFAgRG8bAGk7kr3TpOYeVIYAoq8B/KHvVkqzw+xme/uUyXVthhzjFBYeuU
72TmT2Z7j2PMx6J4ZGDM5gu89y3Jik8BJm/707HZBPOLFJMM66WVtY12wVSh/riB
Of2S6RqJROXO0lzl782479SNBvs3OFGujRgRAkcKajROYBBxkLF4tVSEPeTyyhLw
kst13TIf47G92GiUkE0pyUOkLgXQeOfiVi40nk4AfpW3ICWVyc7CQGmLc0FnCPzs
3IOhtrvP8VQLHHP/NxK57B7Wf7dfIe0CRGJOFz2Mv1WK4zn060q7idQfHNbmJGhD
Xanz4+MlOB76T1xst017rnf3LOnsytgx6W/TZ+yVmgq7WhEzSkKoM15rkplPYjqa
l6WjhS0anfcC5Ykpr9awRlSwEl/eu0G25Ck/vBSF1Hs0bC/XymOpqUr2+/M4YJKI
P456QubcTybJ70MI7gIp4mpiTmm3ofnnqM37T01vjKKRnBuIAbFId7BF/MtD7Mvv
pjwpA60s6hCzUHOpKi/XIHE16IHIQT1fkiFB3C3kdhN5hSL0hUZjoLvHrRbYANAv
B6Bugx4w6zFcBSrocPYr0hJVH9QQE3wuW0sqtzMKlLiLuXxK8gQFTMbNLEhXhaOu
/8fgQ5ZXDDzxzSPUhRYYl5BOz/LSXIn90Nnmk+5qwQ4GZlRO2uuQ8RCRQAzkEMah
rPPfeNbqYGloC8mxCB48+yYr6fQMC9c7F2UgBt8jXks/nOhaun7B2Yzqf48CzSMb
vqGp22mJb1mlAuFyfSNzZ72yjJ7gxMo9w4gdHA95JNjyHwjQzOVhB6OBVhFjphHa
zQMB0T5YDZinBtiqD/B73U3ZR+j2EY1RGRqc1qCjmYgXqkhHYUP9h3qE0cqjruQS
3C1z+4xkSpKtV8NMgc+Ko0zjEmqVQiEZr4tyA+o4bxyC6XkB9RsoRD6u/Iv1VfT3
MYgdOaFJcKU17FueDTGukufiKpU4pDeBTZliGS2zBZyiduYc9Mj0pwqOZsWGwql5
loIFBSzYiQ/Xlor0cZeHtaUHFTQg8+o13DDeV0Ce7XQ/zfRXWVY40z4TawmueMc3
NioYWTXvob02+ezI4Kh96miGyoJknA/5iDdget9+8dZe/If/nSMTcz5ex4AlINDE
M0XiOKdcnSsh66DycW4T/rhZLly8xfvBnTZQiPb1LuOLGdktJ7j007kdjWd4BkNK
ysRxwUPWF6+ERh/SI9lS85yGLnU6v/UwEdenRVLMGNRwMbfFlCXChBzEQb/UjfLL
k1vHngb3MtPqjHTEYBhmXfFR3aELE4mqQDSKup54Q15ldWAV/7JsJULkePO6eFf7
KHfAAaD5zn74XsXBK4+DAabMpZmJrmpiPVdxYIBiPD4WyvpxZAG4mUBV/XOI3+Wo
Vn4cprzSomSMGcaoV1RFIgMHgB9tkfXsk6wdN6h9N9II+lcNwtufDoS5WJrNXSnm
GnWP1bBUtZwqkdsuvazzHOo7hL2dGPW5sm0a6NKdfwARhFNVcYAuoMBUSWBDl93m
sni65uSXeLnTJU8jnqdxvYTsH6UkQKNOM3CV+ShsGxZEf5SquTXwY/5IBcGk//Or
7rO30RDgv2g9qTR6en3saf6dIOD2n82yf0LR1lRHs+e1DJWNSptjJShTaP0dFX+U
Vc1DeCS8h84BpcMSFKSyrfOmgoYEDkxhB9YbWxedFbDgITC+4/HM4bmuifcjsxUX
0GDDGQvD06+20FMoNlZMEoPU0HdR20tvn3LWc+Xv/xXvcpYM4G0uv/q9iJ61Mth/
yMPobN2eoENM122nb7HWod46GKfuvZm6N6keDV8Wo31fJSzcGWRZ4HRowj21nqCK
u3xCKd6OIDcielZl4Sp3VkPyLAx0Ydt5A/CxHuY/bGeOb5P5gGPY7tb4/xyxTAdd
3fOBw+8P19vLgqvxlWgM2VZiOFzm9tIPz/H557sKSWSgGCyUuqKykLUqe6zoTssT
WiQpsO77d3XaOKXqzkZaZnkKbZbMzkVVSCGq8VPDqoT6mjOihNcCNKAa+3ggV7dB
InwZrolD9+4waaC+0BiG938BT5qsUPa3WF9ge9Nux/z+y4kvtqWnJ84EZfjcp/WX
0bzl4NON1TuR7a9cMWDDd0RkWQmLLLdtZKDtnARQbtXBfMbQiff6w3rRBG6/GUOJ
QOFMkW0oplOnAUnH/blSyZvGYj/0MouN54a9w/DQE58B925R/XNzdZ18lsCwsTsN
IyMrWOkCOzvudAGMYm9lTO7c9cddv76CdLYT4uCzNVQExOnnV5ec58aOCQsYv1H5
v3+nAJx9FwMK0uuMFbW7EgMMxoJfvifX3o9w8twqVQtkZ5MomJfaZIADKkPMFd4e
YiPxdC27iwuSyvtBBqHRGPFEezlId/qLA0H4FpnsKmho6lb/fkTir6xYHhYgEzz4
8M1onYAXjnKeVKTaBFsLk2jkBeyKdXunzhtTY2JcEKOc1Jt0+283K9wXH6jEbu9y
JJio26ePESZiaeg5gG2WJGlq9gkvk1lohhcMF4HwA2qvDxH9OIQMyDcsFA/UIvbb
fp0gEWV0x7HX9BiAWtTrcKZYg23gYJh3zHv9zsLMIPwI8tkRh5qfw8mP/a5RHV7V
Vr5XmAE7OO8iggPTF13NDNWXNBaXemEtCa3FWKkotRYtcnPDVDMqXNBkdPI8pWwH
A1sts/4xjDsLoF+CoJWb11CkZ+WuG9NdbdCVuxJPmFHwpyoZapLB9AjKaynuxXKK
cIusrheo9sEnC4LoaDG9pYQUFefYykWCFt6/y06PeXtVdMt0M8AF44xoqEMf8Qei
9RR6qfOsnJzsda5KZg7iezEkPIPcNpLpBKRGTuOUt5oAab2m2Y62NHlZxiZEGLLK
5tK54+ZYz/WxwuUfy2VaOfGOQIfnLoRA/SZ1VXbJdQ+jPEx1jPopDIrle5UD3iU/
V1uiuG6Qdm+hikrIPpYFbhZwdQ+soQKC0FE2L8mpvtdtCSJNkKD3dvB7Z074yEou
W1AaiVyldhsyl+KMt6Cai6Mrj7FqIGyoPtjAziHASXVRyon7nwyGz1ovz0uQi8dd
YCW18auPI/VTfOQp9qEpihqrNo6+YomCAZ994Nh7zmW16qbTrCT3iUV/hfEj5Wjm
yhNs8v5npP5a/69sfzlyU0orrtMC/GZABRabI/B+8IUfm0fVyXQmKoEb/O/RiwPf
eaNSkzD5I9dDK7zRURzMFg3RYHfb56YRGJgv0cTZYeEmp7BSyFSOj9b+nID6P5vH
FDKOHNyDvnChwM9OtLnc8GGXFG9ffvdGdJ3m690D2OsU8AsbfJ/1jlEdtTBgoAXv
FjYpkkMNbadw/0hWTFZfGR5cTbYksQqs/npdZR5AzhC7Ui52u4E7E4S+FAhX3WEh
tbmnLzlz2mZvGMGvFia/G+g0bTRZq90mHHSO3HS9/9oShqAEyYufyq2JarPq8jZ/
CQEd6WQK95RqWbpMJaVb/dWNDgobGdsD+Jw0Ns6eYofV168ZZ6YUO42y4zLZ4a5y
RwzcwpV1zvWfPfATeHI44/21P19eq96vSQ91bap2tlqBLiwb0gC4tl1Q6TMTbbBK
Asey2CBiKXiR8dr42aSI2rl/kxOO4SUZUuEUbtccgT3cATDwkaHOO8aDvsWrZLnP
VJ5UZlSKd504LK9nDysyCgKuYUd15G+PmeHWAiNmkyvpnmexNtvzAwc5ROfhreCN
pozdlri/HfsfhCVvGKu69Q7phAwCVVj60jxw++cYMJdhjRjQW+mhjsIrgrMKYHfD
ssglB/FwNJiy469kXxxYWR99BR8yXZlpHAzDgo9iDDVyuClNKjdZ0vPFQjZiXMif
bZC/sEJn4WcCJZcg1PrikWqElTZYENLtNGg3DM7f76lRHfNaCSzltklzA8Vv/bTB
wzj1ZnbdS9sRCOD0NEGaBUMQnGBP2cjv4zH/oAry6Wlh3c+ICjT/9v2GSwwInxk2
WG4+wXAYWH6xGP0Hu5jtUl6GqD1frPsta5dVO4EX8jBIGe3Pam4SQjDf8atmejr8
/pQqgfv0Ep6d99UCWTrvqOhYSJixamvKVY8fCqx9t4zC/Gkh5ggKNMMJw2eTyx18
JQgh2NMlE7NO0D7aIGqJPk7FOW7wPYt0ISjANGWAFGQkHh7kTr1aSs6qi1ZGsjK2
xma+G+d4stNSzY67zPt39hOJ6Fx/rgrp4tYIPWUvcjcps/zaimd4Qoq4F084ele6
LG6y3hLEYMkU9phkjKIFpWAlMb2/dLP/u+zIXRqOXlAS0UFzceA6ylJb1OCbY+J4
qyfyUw0Jcmw1zKWZ/2jI+zKe7o6H2A0i8FNZ2Pnh98M+9lmNfqtTaioBsYHAo2tR
rAbq9QLRN/EvBGw9rLIdldOvlSIQZf+rmTinpwfQS7d1dQRqMPMTH9SFCTB22aMh
NCPuHBbqhzyv5qufIoFzWZZayQuz0pO8QJ3j2I8O9Neeuo1M9n1o1f4uDouAADk7
4Osv2osTuiVPGAPVvPnvN6uYYCi9awzZysVKQvT54mCGhZ40GTt6mOMTsf4BZOTy
cQtZUYNbqMFPgkO0PDyWpexqv6r0RJGVREDLhVNV5UDimPUE5bAU4INDYb2KF3Pb
qi1rM2+tiGf9MOKgbZZXdUnLzU4JLnE/uDLSxDmkXJx0KE+h81MzhabXCnCm+Iw+
MmaEy4J7sKxAFltPuAScnNtjiz/9Tc0ubzE3Mhu2H+FIG8IrspfszskmLbjXgBs1
HgiPnCRL3mDj0fsMjAwApHm+fwzal/YYuy3ttuAARldQFFShldsiC6NetE3ZKaK3
q8hVjE7CcJVYdCxk4BZ3HnKT5mxaubFcaJE2bsQGpDLQ/xaVKKxDJA15UIaKZ5T4
N8XZMqf801z6nnjPbJh1WraKEb9jz3bUdyMS0GIjQe6YhM5xocK+AZOTIo8c64IJ
D+Bp5zqsJj1RrUA/Bv+M4bfD8kKhYg20kU3lNcLJ9Ela+iOXTf7Y3ohuGkKo96Ca
yZPyD0erfJXQUVFGYQbqkiqU7CykO76KXO40vTQQOq/ZhlxuPYoTDKFObXpbYz1p
l0XcZGyPjXVgAiYYdDMBih2hDl/rMC1ZPreZ7EO7kcXnB+tkRiFLhn/kgT2py/uE
4O+I3A1uLlZ/uCVAVJLU7gKGhubucYbeddh66tmwsmpDZg3X0KopNimfhSytMcWv
3etalJQqHPRTRnaCXJ9DXiE1gL4+fs6bmdpJoJFOxw7Jp22GrDnZTtui1M0kr12U
ne4mk4ohSObK4gvlUn0X6DJnlzPKqWjl7QV1oNa4jJGz9tpG2yyAUEgeTKtDDrLY
y7VQZ/014BHBwLnzfMx8ijgcdTnTpWEZrdb9rR0tbk/oD+vSYr4Z4nmA6vibyfZs
6He0RQC0GQtTWAMMxjt9DFWV+lWymCk6ptl+lQMb8iT2Sy3HuBPWfmlI+xOslI9W
NNF8K4RX69lm9JRKW6G02DN00m+d0A2AmjcZ3G22/dHIXPRFnaJq19HZFq1MSq5a
9AYGl/TwPVLvQ6cUeSwHj3Ig+yM0LfFfzWE2Md9a6hr9fX1F3/KSL2vxFfaB0QKS
hRbG2UjeS2HRbtAFci9CpX+XNR8j3vGMaj3rNeRsI0aNLRSGgzHd0NXr+2y2Dmqe
11nZhJZxXnZz+RGKo8Xh2+c9Km6rILe5EiYDo5A3qkZSTTJU5Kf5ANUqXCSdwHm5
fIsfnVANc2DIMPHrwp+tBZqQu2XZ4GsINX8re5jhApnsk70r3w2zPOOvOjbiUdb9
rOn1OFq++epioWR6aP0KhV6W6FIROCA7QosGjjEdIoHjxUZBLDIcXBI4H7QAz9Vj
cwrEaVQ3Ax+SJszATtyzbq5ISGQeQVtp2sCkBXs33Ny+9reAunyhFgKvpAbsmxRG
bYxQQlKrdcglfDhGK+Ty5J75yvYsnNsxgkAasXepWqLwAlj5cbYf2vxrVi30g2eI
/B4n8Yg5dEqR9ZyTz5b/DmhZZrTcop1cENrYJ9hZFQrQtHWIJuZTTPDHyVQoyJVZ
1rKAuf530PBPfDnlv71EzvBz0ikw/7Y9VEr5zK0YK/ca0aIS9XswZpVvba+DPs+V
mFBcg8nxuyHchtTaayUxdmDW+d6QFW8iT+xzgyhLVP+VlenQ5Z9xcEkKDaRJee6U
mssws38QCus1WVWcB5F3GmEMdd8bMITArY2uB2dAf4n5/SgEBoPLXQRkW+3IhkdY
tWmTaeHWQMKKokeKZ0rDx/MEESPuXM1W9WtEC5q+UwlXnYWPzPxlB+2AyNfIwqyd
WhxPyoP/9EhJ2nXUBvbrgneua/j962LKE+0EQ2ZTr6MP8TV+o4NqpkaEEZI3NYDM
afDL5KV+9m/qoDz7lzkQT0A9uEZQYJWW2IrREeqNCjPqPL3QtXYxsn0z0nV0JddJ
BL1e8g2K/LAZQ0rc9IVglTMiq0dNiJhOeo+ft49+lXrtk1SjSwbNa+pDtoWmcVxE
KFdoziNy3LtNaAZLuLsx4igt/NP4MbrW7lBZ/PgpoBtWilhJ37Lxn0vJnkTky+qR
WvY8+K6w7qFS1U3wABgLc0BDv7uLm8lDcx0Hu/9xcoaNSxQ0OwYVN5mzfmMsQBN2
NtJ5OoUYLVFZGdveC1dVePJn4cUjLKiD9G+ebCtPGn101inBHlshTbaAtbmgT+Bj
Aqkj4SGUYJXvTOUTq1UbjUZdn4BfahJBxPFNvyvR1BUbslFraX4bCQLLZqPfGDtQ
EPF8D+UoDbBBWBGusph8DW3y4zsSREG8Jb/uMyg23cpRx+bfayKdAA6Q3MT4+a5E
/i70Let593z4Am8qn+Fyq/aVMoqbj8DpVbjKZgQnN+BDJIsRV8WMoNy063SxwUNJ
j/z41dNT0LZo6HREoT7cRnXY/TVf7POXSr0crx3xse3hLRcY/fK5q1YBOniApgkQ
qRik0789QZUigAQK7ws4xvVE0eOvhcAVDqx6/s3DQ12qhbvpFx9mFfLlaKx++gAR
i+BjWnC2PulVz4/IvejOv8mpbztaJnKSlvUbjbTBy+LymSPRSQGHSSpzIT7vJa4x
rawsF1+pUVBeLxfaYyL2EXm5G4mJEKx5y1djVjiogbvict/btNFdoRBVz6opKSq6
+R7wBqa0sRPy2Jr7iHXj95Olu6C8Yx7VK5SKZdXAF8I3emzzaFSu8HU+erLnGO5v
w97gPnvbXuloz/hxrSV0DXIpJmPHDQVlDYk16LBo9UcfO4R/ksUHUdI+MjhIa9sq
FN0vevX8Q/q4+23ekWji7qkut1o3zNDZbYvoyju93y0++6AnLI/xDYuLS7845cdf
hRhlswrIEGghcAM+ABu2tDivgnCXsfv71Hu8YWiMmnbuk2D2g2iXNKgSItXI3HYj
UPWgyCespx7Z3tD02ZGlrPUVG9avEhhUlAK1Q1sd9bCqQa9nuL/6qUbxp7WaggS0
lxLITfO+Sr1jdQMHS+u3dIw7iBzjGp/PmLA8ZYhAjDKhGFoLyyEcCNO0wkGj2jk1
eG0XuwCpNrRpGPTdbfNR6bragTmczkzBUYarrqWHOscIEErZcp3E7FtegsP6ZD1f
KMFGKj3JXz3c51DFQTosfYPBwU53alJLm1UGwo6M8zbL2QbxsFgL8A8um3wrr5vX
vM2YkobSApj+1pwaviSBeC5G1JPn+T/jipBlfybdGYJLtgFLaq32ijNzb9F51qOS
vcn+S2YIOkEu1yWsuWJVCnhZ6KOjYW9mIj7NHGKtK4tT+r+5+Bsuc5ul4oDSrCTw
UK7tJ4AV9IbF+0tbenUEGfSzdb6hGl3z+0TOXwoAMPYh+u+EAiaWariVf0elp4To
1B7ZzZzlZQWP0LbOGB50Hx0bchbgdbaHGdmZsBsrMaOQ+eOZrHFBNbKMaiqRNN1+
oY8Ibz/2wsKRh3pwePwWiN2R7MKkPnkcHMliRVqjIZGnxxiJ0C2lEGTH4QEOTchf
4oZIKL68TdXHansLnS+DNfLSIUFgAsgXls7XVd2IZIflMZUSTN/XUURzMg3Uqoxj
DejCVKNWZsjo5HKzw7qmGlhmC7Ro1ohUo6sPrrgW/OQwWAbraxDTYmE4/pFByZpx
/oHUNAC9ekF0+hO54SDgY5GJ6Sfv09IbJbRmG6LYamL0N/bZ9dN9V7m05wPW15Ud
CP3kIgxeqcrDGxNIqTaLJJ1KMzrTwS1kpB9GnI6MuRsGDGEiBDRhcz5DXVhWwoi8
Au9gnJnkJGcWQUOAxytdVfS/Qz1ev8GjmqMy2rXv5AJbV2RbIuG4OB6KtIWd4JLM
tMRDSwShmII/jf8PqsiK18ts24oC6IwPBzNETpgXwkbxMEqiDypWn/34sk2AA/ob
NpVa0IcQo4h0AF0EzpJeAWFEsbZZpUFvgj48Z8t3mwqvVZBUuPNQ4FCCg4+0rfHj
rmJLPCl01QdPnphToU1O1o9GiLGDiREgGL/rvGfR0uNbsKryk2/PIfh+IsELG63l
lqW4iZo4UUs3yu5Ga9TMO2kl1lc12wq/F+LQa7DGjacx3Re4yJMAVkQGlkO9liAq
e9UHBZkYD/jL0Y/lJqSQEGMPfLEWKpMd6kY77aYO1+Rs9DGJOTQBfiQ/aExl7Fn9
tgd/kUSp0+vARaUP5MBo6ruBtCb70Rc10n8fQQeYyzNFaFfTNs8pi65Eg0Y9Abe+
0ZXsjgQ+pZq/yyA/YD18kZyhsZ/ASCJAHmRbq9hdagKgFqy2PUoPYmXjcHgyIUFD
vuz5PvmGSklLt7rRgZAdrbFH96ZvqtOdGpyjCv+bprIaDJ9/mknk9a+gk++leztb
MOCogi/rIbqFwICuiTCFv9GdbOhW78NX7TYcgwdYANj+HmSrQ51xyoGUFjzhOdCR
00rATQbb7S032sJU79iTFLXptyZN3GU13eejWb5WsxWqlWf0pbTc0GgwSq7iCTcC
6HM6gsnn99MJnJz4+iUCB01nRYNkhmHhYicM99IaMPSeU33QtP39p+zgehcSHbHJ
KdgwxiUP1PIPa4PXyS6n1r0M3A96+HfjEFZLAfUSWrNTSufJAWQFpAdd21fJrTI+
YZ7a+1fQdXkTg2oZxIKWu/gAJuy3qIplAL6p8jDNTrAodt2/jbNxl0LRIaG/fC3U
gNSZvJ+DAo3n1MqMD+f5HDk4x0dau0TN12ilgwbMRQsP7FtzIT9rqziSqEQur5uD
4IK9mYR3592X8Pv3gKwLpfzx6QQByPtgHSzpH/1BE5wckLKG3cTDt4X2ecqFd50B
TMr5kEUW4ej6GQU/U5pcwyYweEwr7bv5lAqp8u3N8iR9cTfwdbhF32/SYIYYlY34
K09tz13IZRnto0/SfNdIaQAJSoBe7MtkgJ7vDJBjVQ5gGeLB+Wpk9UX4dXkLZ1RB
a6oiuMHUS/KkWA0zUZL/OnRJZWoG4EwRwxKwCvjhqJDqIOanCKfezCeKycvKuspG
bJta8jUVTJ+Gg7hLN7fzBmXjhqVKX4uBSW7O96BXAhsBEXF1sYHtRsGY/WkVhD8e
4EItXYS6Un3OX4fxKOqfYL9HkDf+uhgxQ5J6tovyM3uosvX6niKsW55dwIs73h/g
N6HmpSQHCGfKm7Etqf+U/6Avxmg4UQP+UwG8MfKaBUoSga8yqYt5IgETJWGZzKqm
hRYKtRoWTfdZorjpFEugi3b0EChxVhhPMtGtUTbiE1nZie2xLpNistRPdeI+ogvp
86zlTlyH0miaCmIuZorKKFmWpM8E6V0tlU0NrpA+edWIzNECPdy16Ng4iXeGKQGP
P3Y/bxwk1ki4SdVIXuqXJsZRzMHUlqfPy2ioeJsUgjEhQU/GBlJk0FafIjDU9RM9
j6lkr+8EMjq0Pv4qL5iZoj/9pbgzTu+uhbb0/LbDNblO+wDQ5Q9+Wo9xwAms6Y8a
OFBQtdZ/5Nz08DJ4WDaiWPKKfh0+aGG7k/8ux9m4AKzZpIfh5BBtzEOUj9M7zxBe
1tRwWWiO/C75V5RmVElLidz//XKfJJGX0ylJo4r8ZaDVZjzgs+xjR87GdpkY5Mka
8eiaaG+7ImlY0rmd0CB1siV+1PRn5qguf2HcUr2Qx50lDtfuw0rrpLVZtYF+RIkA
1u1/bZpXlYDXMxOm23YbXoFvOh+nELC/OxdF+42/HDFz0mitAqGreXWhR4ozswnG
4cwholsdMWtOjeXHtkZe77JCHnfOkCw7zbM0HYejrMg9h+0kLsaePuKl5qZ3Qlts
nMikLMzuT4PPpHfpSc5Ra4QWACuSSNvrnsGd2Hk4zIEYWqH5QZ3Uu1Z/MamLFaia
+l4wQaZTFN3gNPNAHBSmJI4UFCeMDtSUT1H8/ovLl59MRJsYJWVUlWDYx7NC1QbO
nvS2dSNS2Me4U9oJwfnhDmLHgjp+wYFvVMDbri7x3+/Ue3TxjZl6hQWA2RHwVKts
/s2gEEljllMSOdSzisYxNhIUSEBVakY/qrMahD4O58a2K5A0y3cB8mbSYoG21tXb
oAof8HCGGgFO5fzvDiin+29srTg39fshjbYZzpxOXVxlQq9wyuyGYkgT6eaFPMUW
jjw2dQlBOwPKjZIU1vzTJMzlZ6a1/TA6dH1Ic4DDMvbq+zGXYux+xbQe0Y9Gjigt
omHuikI/DR1RotFiUNLQGxQbuhLeGDWl0RuNBh9PnqmCFx07FeihBd3STqN4ddkf
AVItmvrcRIrQrhBrvXOH9VGzkzIajEo+Ag3CzL1PCiUjcewzp6VK9xEkDyG+mnN3
eusfjK34LLOROfUpqg8Sw/KnPPJt6eIkdU/kLCotFkYaMPMoo4nX8G+XTyBymsr6
Vw0o483aYxPLu82drEUnJa9EBSL8WkKSXjx+4pl56C53fhw5Ach9zMDaKcA7Rop+
ZsoZONqQbLOGyHzi/NCWXzPWViQEB6TK/+b2RqR3zZelru9VYMBIu+AmazeWnyUF
yiOHofYggMKYMpDDI573mFq4cN6kcY4fkiMUFRR2gt4zWDIDpfgCVTOr/lHX/t8i
zvn9lGQ4PFsJvvo1KgxJDm2t1J4pq63g2rSaSBJmYan1G7Y1771NzAJrVWYUjnk0
ZPw9mJdiT9SZiHAIU5SwVUTqeaZzX6Ya4l6gt0tuvijzIZksuBtgpqQchhKUYA0x
c1mJgkfMK/86+yIfzZwOGbxQUtWjOJd+Ph1oNHxfbEDwNw8ploxgPIgpLsHgNcNK
wQ18ii7d1fV3duFGtnFksoo4e+vLGD3/2/9WOODyLXb+etWBqUoVxdoPFtRC+f2k
a3l/k3RZ2ZHo939ZLmIJi5eXxVLKJkWOjb9fOj+xSpXNKGFmgtn5PmA3xciHVE7o
UrZ3rC7q/qw2TkLmEjH9m3qskwyeT35QVgo+TlHUUzFImFl3XTnQs009C4RQ56+i
Q32jQdmzia7SKu81paBPlsQYln73daR+v9OlZFkOiBXp+racuiYI0E36HZR5POIM
Xn9iagUsZFEQfrgZ2WjE4kEnb/lauBWUJe9eVgELyv/JDjHdDqgsk94GTHkhqqgd
p3jIBbWTxZDcgI1HmL2+5MQzRYCjatiYC5trE1vUL5tLrHcRC6tHYjz9oxj3Tam0
waq5+6BrWTTyHNPjmt7394ooGkpF6Mzg8YIkpgfADNkctFM2/mZKsU7hLOxSeO/t
4t+pZIFT8kjP5uv0Xj+3XVR+5pUgj2UXO1D8KgNclSHLXD29XgssZ3COiNf9J87e
ZtbZUAz6PL3aOeABwP5ZklMN2vDRUpiODcscGrKlQkZL5o0J5q2fqHwA63dToCGg
beeMIaS3lBiyn6zoqC4VChiP5uZxQOVlpHQ6fQ3oUtIe8EMGQwzCnXaxw/A6+mD4
E8bASBtL9KgslH7Lt3hsrihwGrB1Cyi2F2f7je+HqGISKzieRgAfE1e6DaEdhZ8d
TpIAgNxho7z49reCGlwuFb1gJCJEmSs6L8icKoOgw8rJ+NPKzJXMDwGUWIhTnfrz
i93q6yuFvH2aV/tP52wyA2WpQFeOZPe19lmYtSz0n4nVaw5GCS1/GZXmxa9Fxr9J
ur2TGBPUb1Jw4wqIoRHa4ZF6UICFA51bxLfzmoHWyjgSpme4m/GuMviVhCYdKwkS
RpRybgEud+/ZIGhDegysw0PNxJZm6KSrYFiJ64xz9FsmA4EcmKKUaGxsXmKVW12K
9rGL/YEeJIJELJFJY3a0EngLD9MSMhXkDBSSyXCXE0mJGbMmRGOpKxXkn3SipYOf
Ai23JCwEL6VF90rGkFH6CTIzYEVz/6htuc2ztGn+xY/37/t2UZJVQdHe0fZfaAwN
hYWQY/7daI2WGcvYGxS+5r96Cb8kfe+N8wTGiwHvJRx6IGYyw65fEkfudVhWvBAe
AZ2WlN5z/q7WkEnmeMjT9V0PKNo3QZEeEC40aiJ9JRC1UmZWGVe5NPt3AHOF5qNg
tlvqVIcwpoaoyizdWZKZMTcu7aJ63XhmTxzbdnZfQBt3jOFSGcJWokDBpLIxbmNB
YtdyJ+uti71xBQ0WuHyHCX8tSdInFX7/pXHTJdCEZmUlSPDmVNsOvGrpk2fPk4rX
H5Ey89dOuNY4Lh7vVB/iSh5DrIrpNOrTfq6SRyFgFluraYenqsx47tl4POHNR3Xu
Z4jEvPeebeOLvpXKFmO9QYTeUSYfqFq8dydTqpOGUcsnXL3grEh29rgRziPMSbGs
hcgSYZvsh4D3ER7U3QSNjux7BFWx1gdwcepHmHvjbTtcvMWehAdETxm0eZ+AvBH0
OLfZEGeoYi2sne88LqcZEu29BkL1f/awKtw4WmPPkDj/+tn7nYMh4m2RF8st+EwH
e2s70VtFyDPcBiQayWU68d7Eg/ED6Uy6SOcnl45IwwhAErLZuHqgWIg0iHBWi44W
uxG66RX8+phmjFVvzJW0BYb/aJXggJXeTLpjwpr+B9uiNMeDbSq6E9U2s/3SArIL
5GSswc3LPx77zgTDI4i1Vh1a6AahijxOQbHu8fRJi/adDXHEoJIr49BMu6fzESJ0
2DA46f0fkmNLo7u989X3asuuaNFYVVY1khOg4d2LfgzCvffRcdIBpb3lR2ZQI++w
nXRC22wIg4CJ4ZaPWzvufNLMmnRwaBgi/z3zIJ1G7Kzgy9o6PstyStJYQnikqBiR
cCj/iCBF5DF6x1TlqaAmRp2LzNe+LfaoiW1uNGsYlIWtjQWtmOxWqwoknGDPs+54
CY07RM65bKVixkoDCEFx97G1Z2eEXPd53PrrJ7vtzbmLwHL0ui6bKeXOF4Zz1uCr
+jOBhEDhuxso/XQP1ZhXXXcHJwxzbjZnFxIWKms2rs+gQ6ev4CiM6Sbbuyb0sRyO
6avj/ECRyeAp8c51RF3tb4H75cGoIa5NNcLE+cAFc0hYvPjfQycFK9T0dnqpZdlK
fAQ3H1UbSzsbOguagfkL9doJ9EAfBCgsuMNMdEgpAsCgcXXAo71BcpdAIg9mOinP
wpYcVNwd5ZxWLBiPh3lk29+q1J0hbzg0yePW+wxWDfFomAaXsK1vLZVD3au3d30S
LdF5hXazeJpVIcRDrRSuvWFNwxpkgcaZ/EIOOj/4lVNDgNDgi7Z7YNm21gHrC1ha
1Tokh7982/ooncuNjFUITiK1WDOf2owwChOSeGe8kPCneqqDLft1D6RA/dkhBfQ1
IAU7LKBllAhXjf7LncGZ5r2+ptQM/uzb/hhNaRMQl4WsTj86jbiYJiPpAWZrO2E1
okxYZDewUbmvqnwI00BVjvDTYJBuiP1O4eWMBNU1qKc1os0RfnjAOwts8Rst+G55
rL+AD3YMZNFX6ekHK8DLN5Fx6N31fsB3ebSs3DC60/maq8Dy9DjPi7YUxMaYOnFM
9lKAEw/sB++H/ZOFnJ0xNEclWeI50kMuJ2EQ3FIEOvmryOzbeF1hR1ogo2jW00ok
L6pSLF8EDXzp68h24opZs7PCw2Xrmtmz4O1s1LcXmaiEXfSrglNcE5J8bAbTfaZU
QXHUvavMiF0Tahn0qdfiHkK0tye+W8d0qLCRWeSBnxwmUFwK6MJB+3EfFrUbhbVe
tbxPt6+7AKlq3aTfo0j4iX8m/uH20oRnN6+rTWzgdd0uCOrWXgFSwrUbRw068BiL
1fhBVLnjh/jCl2q2FwlMNPn/gJjLHwfrOszYhDEfJ5ULo73rFuyDCeQj6oSKBK0t
uDIEeXEH1ql0tJybxTVfkgzMcx/hzEIuiyiSbBCe++Y2jk8zVzpxXOfnFhs1US8N
IteKQbeO2ShMAnbTtvjnosxTyKMjeJM0OagkcWXm3wLXzXX3/4PNkaQYcx0MM7jV
k1Cf5NGvc3XdM60FaL/kYc8iXgR4jqwuMPqiwpj/5SF+V1RhPG0w2cOsTMEQj69z
AUkztw8quKJtpnlRRSN6HZyi4Zd2asZeDFFeTsW0vfv+HZ//cttyx60C6yKPbLKX
GB1+0Ym+pLUA8ed040Jb3sSPjPK7/zbOd3g6xzEEs8UqhfKDe053cUpALnCvxIb4
iGQVlKA/vOb+9411yLeEz50nPMsvsuzkoPmbgr7LujtIVm8qVJY9Dg4/sDAysOzn
jUQLF3yF7oku/p8nQG4cFSNemqjBgcpN90tb4u3V5nbdANnkQGAB0TLcxxcejCqB
aou2cpPJbszIgtEidiZGBRXshAGJvp31vVDHotgjJgxzLZ6/BzI4eUt71ApaBbyu
PTk9tT4/mFm5ibLLepgwlhvo+4RYgyEPCdCyGKlCefFNOlrFOntbGmkMitJrVmfz
xoc7nqq9ya34jOuFkQFud+eP8p+ARBpiBDYu32JcYEyw5Wk39mXG7mpRh6jcw5gT
7sqp3eA9kQ4vIOUFXeGN1dj0bXy692jzcFCZIkolojXuqYG3IKwqKKy/0JADYQx4
wCoVkV2huuxOsUeKWkNDYlJoG6shzQjuK9SF21pDUa6hUTJBh/1mFYw5vUF5OXsD
aL2hn6oGpnUOQdk9HVfgwoBzhHEz9mugB7ds1tQ5+P5veiPZ5i6bkVTI+oLAA30b
lvnJzNglBRWsMfQHtYhJGBoJEuf3PVFyTJ2MFvSRJix2fog3nBLbJkwilZZK2wSZ
uwdiNzZlvIimHt13vpLaRVJ+tXo46xGZK0ugvGFc4yEPv3Zp7qA9ZVRrpqGbgL1J
KQL/xvG7oUiVSVWOXNRMzUjOhXufjvKoHhHeP89UaMFm6sRxPs8V6xyKJGR/oSiM
eeYjOVWq2kipUUPyPK6TpeAXztQcJlqMHw3/8pwTJtkssZVVaQX0DN8wqe1OwP3x
xPuMvuQItyMCSb0P0Q4zMWXLpXvstdy5P5mbdbANKT0iqgfcZfg4TPLqeoq3Wpr/
8Zk6zqO5EBwvQUZmdJiKELUlixsGAFlnNEt032YeXY0mqjmEAfLbFzOue5aUUOiV
q7AVis0n7OgQ76dfFe+4ti1A+ldvg0I8EadT1RWgvzghnDx5doXAYFnreyYtjxDK
pqct5jq2kbF3KhrUXMsUjZdf5OMDQVHZL+UYMDLcSsXsrkqvlaI+3rcnZJ7vslwE
cH5RF5ecrhL9tZ/eV5fss0ndbwwErCo6h4VMnCaNfYkGd4XTerIQkr5uQs5zo9NY
heuMkRfFK42AFL8SPgXW/edZ965NrsGYKhS5VyuwK4/8U6VTTqoatMW6d25NAJ46
4QpvlrF1CRya/ym/td77qlH2t44wMCMN7YQ9LeQqr+j2eWrISs6BZ+GBP/LVEn++
FZ67QybwJhkJjr6bdmWxO7QdiBkU6blGVq3EymgqjdKbkR5ccRfxRf/5pwvGzNs6
DdRoWdV4T6FxiNfvFexlbsWdewSvWm1GQ+5DIYsaFGcgp4T67YFjpphNtwnIUhHT
zlvow3Vn8szRblvhovEH7RNWnKihU0Lnm/DnxlSlsrtwYHc1qCtHPJz5bgNwFGU0
mBnHgWwpR7JXJ7KaB0TkTtXlYhnIKfrkYnzW9d5N9EWSqg7JcU3fGBjiDsQrtM2K
YtaXNtihcPLT1IMR9UkYK0/GfhsQOqIDWHeauCQhEelU4mZjkaCepil+WxfecQ+k
nPg16Q0OXvwlmMru7YXbWO+eKMrXmA5dNt9LQfj1WRWaNLyn9YegxkSYsjcOdfZp
vZdsqW3oyB9UGdpqitbVx3SSWXpgB3dPcP6d+tht88SxU/ymwEKKxZKO9yQPrlaQ
WLc+22sVUEyJ38xKXet/sLoH4vrJ4bXEUwhvQFe2e9H+p341yaGMcg7m6YhK2Si6
61XJ1vCTwpRmOBC6V6JMtZGXWg/IYqLNfCQX65LKqmMA5kVZ+TqkhujjfUF1VSCW
FzJ91rhX5eBIeRxrQNlCo13quuhcT6Atg1hN108k4q3V137IKuEBt1pOeflSfF3V
Ip8QJUFtmX0swcgyESTJZ2+Mk2nYMVJc1px1UYgfIuBbOHnV5+NfFyDdXEWslQgh
ODTFpb7IP1nCxK75aQkIdLKJ2L9oxhm/y0ThmaJSZxakEQSpHzqKkYwyYX66DRNc
nYqGAM0AI/Sagot/Ly2BvGXvOVjaP8gmuh+oIqUz4PZkw8IDg2uI92L+L/OTEbgX
QNCdRMsJkD6/GYUC7zqH0uxWpXwOvZValfsZO11t7kFNXrzbXoCbDsWNA1rgYPU6
6Ngjwnk+6ydvwTHkHGuRHpA6izIC9lKtECnZ294FARHLjH0pTfNqedeTtzT536T1
VWCW13SLpbYynea5wjDyTNvyAORJ1Jln2bF8eAxN+hTd6nga0RNd5H2U2ndVJx5y
sIWqRt9m9agYWT+s34sfcJd1uxqeLS2V+I3gGXcoIILQsx5nUL2GhIKzcOjc7V+M
h0qRXBgGRXgGM87XwnAgGD0ZwFtYVrMlag1yUbJP5h75Qk0zY8vgQMnWPoP97ypN
2dVskqSnL7gHAQOadwoijpxE0gPYZCBQ1z9e5BmlfU0IMft7ZwS5mAfsoyD1TB57
vqdN/gnIlIPhtJAKGHCM3ble5X9/bA8VMNw0rvd9yjfvESbbXFBIRrjky2ppSqkv
/sXnnLx3yhDqtU0y3fdAKKD9MU3LsSTrNucXDWf/34Xs9ce8CjZDt4kfgmdpLZWm
h+IQkEb8oiW1crrk912Ji266aCsioc0jwjJDVQ1p6PUtSV7HLnU//FJJs/E7rFeP
59pTjD55tOkcPK5bI1nHM56onunUHtlVF+qhAqC8b4xGnGv3kdOGKOFNLst2+rlI
jCUKe5K3d8CXnK7mEsiNAi7wj6dPoloJj+dXUdfaDY2YsF6DiGHhLitWVKmZdzhM
mMiEuB78N/QbOMaIAvmbyGwgIEgmUJlUgANqYu+TIlEwWJewicZeev13nrWcB4nv
t4YERzD5qvh2ubC2mxUpBWLr85HdYUQhReQbGTj2wKpc0VtmPdrp23ZaXCR8M+G0
Mj7LYZmdfcx8f2UL7SFR+AFtlgvtOgLGwyiidyTebdnDJ1lnEmZED9BN7ZhIEgGL
NsmVov8ys8i2kXROksTfLp8rIW19OBJ6DTwQXXMUtFZ4roEC6J98HYyazELa1D9Q
2F9+Di0i3V0RVPPRerfUTPC0uyB6DxtFSR2yoTNfjd6DpQZ8u3I0yYWzoqlVkHr+
mAZjZQ7eEF73Of18GuoOEIa914XdQaDSMdoHGDmdfVcTcLlp770fs9xdO5crPEyo
fAAi1LNEVrimj15QYT4ODK8U+VFw14ZCLGEQJrLge3dvQi2IiCpTz7Opxplk8jTZ
eb/03S20R7d1KUWE+Q33HdgpqzEkEe9kGbkEyySmP6tObkc5tun/GK2s5DWrc2zC
1K58O4GlMn/MVOpcjIHbvdJykoUnfPVIIPng2/3O9+sl64pr9IE+HyOMfjy4W7gr
DfjeBA2bp3Zcbjq3wRimplXo8uK95WKUp2XFvw9ykhna0zb4mdHtpxCXcHkv+4CD
PzmjsS3vMdCUP8acjxTRJrNlI49/sDFjvE/CpzGfgN8/PqaPDFfytfjdOanuPwXI
VeaLr+pGNRC0l0l+UYe3wK9Vgkq7ioxnQ95M0P7Ci8h2hRaE7EC4AIdza77ls3N1
1aRWO4qHhvxleAofTFYbvoPGBhM34XHx3p06MnzUODZioJi75e/8JaSKC+2ZLQbt
oplv7fyu5EoQG0cLCnyxI/YpD0B+va1p6SHLVfNT8QvtAy2RHyu2ixt8buYSuWQN
upszUA/kILo1rMTrU+q5xzYuqlSU2SgNvhaqfhWDJ1DOygAY/QfxObaNByFB/3Xg
KSxQW/+dPS4azDkn8WFd2wnX3Q5d12SH2VnCggQhbm0roe426bzekpinNDDJ4nac
Roi9F/Mof11InlfHTerMMXcACUYDz0fevVSt0acXgJhBKaz5GOf4WhmIDu11hXjQ
FfwHIEAfL0ssZYyAr9y/LonQFT87maNPJT+WzhSdh7io4xhIj3cjw9vVRIcyx8OH
Vkh1LWAloFzuV+/k9cluQE3rOcQO8u7g46cD/9Uf94MPTq4XyZkQjLnW7ftuOqbH
D1jkNgtduAXIjlaosIFt/MNLNhrO6yfuRNOjFdh6pT9QidmJ53AAG/SXjWEK+GVf
umbkbz6jRJH4kBNPFN5PRaxEc9CGCcdYow8+8hOfPv7tz4P9gmooWm5f0vUK454T
vTxjTwGd29BkweHBp3Z9BnK7VNHZxXUorsZKLmtjc6UwWaS+8p8pU3AGd8RCip5M
GUlBOR03N8h5IG1T3s+bnDSIaKGXG0sNLJsdmSXkxVyM3dnMRxt/5VcG3vPA/7DL
gNvXhHt2VUmj+TWLyVd9yp0IuyhfgmMpjxZKzpqA+pnRDhJeNb5Z0FHbLzt/7bjs
NjLJtxguttIrQZyee4OdMvJFuRTgO1amEuHMCg9cTUo5NqFsEsoTnHiTaZLzQ/Au
f2QE7BS/FbwgGVd63NtNrHzYH2XnTqMqWt6oMdy9ZJalHgZ24XaA1H7lOoQg58eJ
kvCKye561OhKiB94kqUShcuRZ6SZkUdutv1bxWLd3EkgzqLwcqDd8Cgqg5D0grMo
7MxhNfE/lNDoUlvK4w92h8J+7zySdgBaoo2mZoCQLlKyG/ZnN5pWuZWTO4ct+4DV
Nt3OQpR8ofBb8nLGSL0YJ8C/Q8B8mhJsljkcEP6/5By7Jqa2tg/VxuoPHGOABvXa
ar/3RGAHd4u/7QNxxGqjoU00HohMaXDgGpkW4uZ0HWGAbRGFwty012ns67pp63xx
Z0ZvgfK390vKgPCfgDVZUpz21CjyJSpErc4SWUTA/BW2j3ue4hEUIySSQl0mSxsg
oW13x5UHTORW/CnGkO1dqoyKSKC189BkMV7lTmSKJb+2TOAaRBVzTcC+7Cqlw4XI
oagOn6KStKp/EDp5bY7aLRH3TZWCjNbCo0jqBYGuZjc3GNtZI0cUt5BSU3O/rAuo
Qhw51rrSitwC7E/TrsLCGF6NRteotFjphAt5G6ydP5vWjY39+QiTnmoo/+0d4qp0
yTf5gx0FCjAOpw7OMOSScit5zO5oXLByHdyqYeLlEW3YAmyBwP4o/sprssnslqqU
GWDmDuBrjCnuKD/oeMjbQw4qYYMIrElV1U9xprjhV7xNm9WLBXtpsfvS7NHAjMiW
WcLQ2bbaR81xBD9XzxMgwPLjaKj+z9BysPMLkei4D/wPqKCoyJkkcCChozWCnrAN
DsX/5fzveWnWY6rUkx+MvQYVhC2bhp6vb/D1utGEQHJDKQNQsxvLXQ3TiNLKCX4A
NDWvbkVpldh4st7DCLH7kynWtc0FoGBMM2arIZmmV6bXmrlflBPuQJrP2jmjyeqj
8q6LLM00wDdf68WrpVF/kt2d0fp1rYbgOOVcw6M9rPlGQ957EazVloseYTmXbf+/
qUZXat46kjhOh+qQvjwRhLdOVHXMmNJdd/ByvPjofmHtmtQ96moQopRWeyt+l1i0
hiVGx0ae5OSjm6vHz64Udz1qt0BFf+LjgZnj7dqZnOZ2Okm262wP2nx0uJAqbT4M
H4XWBw3SBYcpseSv9jfcjUGZPUkzKIPF5T9p81yRbdydsTideTEfP6MqcDoce6bK
4i95nYrFA/0ZcYgvJnh84YQST7HIKCa7sgm4HS0pmDYCOY/gut7mudO5Dvs96Q/U
HFAEUG9jDqm4bxo7Q+JemaGXD/yBPH/TGXdANoUCLMtzKfKQIEobGZUdIEdzcCQV
Gixvm8sI0/3/f/4pmaUXQ2xqVSMQngHhXahAjmH2R+8q+dd2sr/aQcc/jHJwcM2F
OdSLXoslEeJpHY4V2N51i/RVZQ/4J6Ak2FI5rI59ehk1guPpbHsymDbBc0wlOwPK
1OoIWEvlxXckXHr45y/39JQvvwIXvntKc4H0FnCarwJoIkTY1DJditEty5y3nvm5
PxJ64Q/4nT7HyJBgmYgU41//wLcZpgx55daJTC6nZQcsh1x313ZM/1nkwmt7Aock
6yd0aQMnc2cJGDxCm/Yta414ZIav1WvP7rUEI0dT4lwPWTxmweVbNxppfjmICwrI
E1r7QOEGuTyGkNpzgMTcHw1YAKVYF0UGx4QrcKSEAiGILq71rmGMFkxh3pNRZNOT
iG+iQ4fZI/oSYWQqcwITji+c1BSjGonMqhs/mQZeRa0IS263qAgCSQVuesExDwcB
CPqO86uZrdjrCT3mR0HCdMv+pyh2qzevI78xyfbPW4rzrP+VQZ2sc/iue0b8955T
r9hNcBORixJs8KKySkVuJOAJcG67g+sJWeXRCA6EmPkm8XLk7LxuBDcHQ2uRJjmj
Wu80J4cG20hL45Jst5UZW60Sc2cfoDnxq45WKNnsLCg61QFagXxJBg+L7HlCa7+2
BDYPw55blxkqQ1/mB7osljt8HSp46lZyHv4787vqasN2IJct+OBaiHT5BAjHMhie
L+rtLqicnSaUaaCvnCT/gru+6hMebZj4efPjP4uXTzaHI7pwHEFziDEPPCa/6KJz
VnPJREfqSpUaLVac0GZblKPHpnh8jwU8V4FpwHkS15XnKT4WL4B7MLNvRy1h67Gt
oS78Dl4qfiwZ6yWqUbNTiqb/kvdOIxPyM1yPuq2KLNoZzCz5g3gykjDFi9fvfhFh
VbVj/fY401hDoR9L5ECh54bN4ZcaBD3PfucUXVzChQ0QsADBrkFZVFuEJF+EvMI0
7ECqR+EakktmMkxzXqsL75IW91pifhyFL9xqpUeg2/1w1NJ3rTOnStriYY7soq8w
OPh93uX+3U52ZecmZVRTBjLZuFllJJHNXxCAUalN2Q0/xJvyjFDNOvwyQyF8tse+
+my5FvQ4yRD5b30NJQx6Lsh5hsBMiFGd00Z9RxB4Dr7EEMfWqZFWMK2YDK209snI
zSamLb5WKNw+7vu989hE3FZzjWh0jEqbKRKgUE1ZaPOHxM5zXas0dadKaBv7WYYL
RmZhohp7WDt5koBLtZcOgp882a3v3T+oXS7zMqYK1yBowVGyxNJif/mBfIuD6oha
9jc910uu5D6lSMK2mhFWyBr2035c2uNz1FmqqD7enT7oIFrSQQIDej7SCAtDMZ1P
Wp/IKfJSjpLwY42IcTtSfFABm9YBSSX12d27OqAD5ZcDm4uYp236OQRy0JKHNd5p
H2n0MgekSF9KjMcXzvAdgCu/87MV2S6mqunU8RF5bs/OZD35ZVCXr6hnOPtZHeFC
kAwrMK4biTESJIw8OVd4XFb9gtfGrj3LR1SxsquVCgM8MFFq9YSym7cK+C9MV5Rf
nQiwjMGEj6iHMhNtFQwHxLWaJXqxiJCRQN9s/cbjpl56SfSceCmIYCRvRThx1dVS
oXtua7o06zW0XqsmgEEijgdoxCbVMj3lbg/sa0HAFERG8BGDunf+uevTxc+qVD6H
ZuKFQwcWt2XCFW3In9/FVjMqnOake5sYL/kjnwKMgF8m86I/zVIk22ALzco33O6E
5xER4mjo+qXy6Hf8f+Tyk59CPmZ+LG6UvI9bHK+oo5Oz0W53ovPJbzeuTYlPzRK5
9V2xxxxK4R8wP8cII5DQLBNogfoR+vBL/mpqFVTQyMdX0sgcTm2XxaqvoMx6hgK1
trA48rjaqll5vtdQUdOwAM0u2WJ0T1kxfAAP4WJjZ90jTQ9eLqrhQ+4ip9DyiLAn
0sQwaqO5/6/zaHnqbXzCETwL2usqzZ8tahtx/3dVoH0stfOV3QK9G94V7zvtKYFI
/vxHhtw5k5dvVR0UwJutTUOamnFO9eAiLsLrpwup5jADaQo6UyhGa5yBZyspzPzf
dK7O8PdOljBh1cxoXZA5XZMjz5IYKCIQ/mZglDIvdu5KCXjv3mSJHP14SJa9sZCZ
jcjAhH5D/99HvZzgcy7hyGQuOcsVERXBa70H5LYYf5D5aKDx8Wk8ZCSgFHYHwtRn
sp9VTjvc/IyjJnJUjj1Jgty4JlNPCGkcHVztFjtolxihUIcs/vqOQyqgVeJ5CzdY
TFC7KvEcE/HZ7L6a4RjBdwnWJYHoEReyIbwIPLPwePAMkCT9Xg6t/L3ytjIv/5nL
aHYcsyXBJm39zMPImwxLOfE5OsBN8xmzOQLVvZux44jfhsUzJtoicn6hf6rc5Wo0
hcLrjYAmfJFpSOvcuowployr3BneOBoio4nz+nXeoW4+VeOINcCsRtPFCJoFT63d
C5pLaRl+/mGNfJAoYO7l5oLP9cUnP3raj0pSH+7Br1XjslZpMOtekOuHQ9Th4mDM
Yr0YQw2cpjQM+6oltD8aDTSWl5Y4SYMcVVOOEn44qQzlNPRA6QsVedCwlmY3MrB8
LWOkbJf4BzC63bdhLgI7cTR/Dj+XrhZPXC4WPkZrQgvaqrWnRaKAQI5lRanem8Ww
Pimnj/4fn7FDMsCySy0GQD076ZeV2RI7TH86cZelM75cux34hJReYGDn7DDQCNeT
rP1oGlXfcHU9LBo0PjchE48HnVp2BNscws5zaZbQuAsqrVtM/ZNmHStTMe9a+ZB2
xwyx6IYt1MlZYnho25PwIlRDtmueDO/zVtqxDB24cd1GRDFS4PChd+zgNDdZDe/g
C9zTUrxXIG/RHyYpJ+a9SyLr3MeR3v88EqI7O5CrOlQvYXoLnRohOKK066yLjlIW
C6JlH3glQlbPrJiqp3cVhHI5Ulmy02dgfOrpLZ3iaIl3ZOp7oU1GbRkkjGUszoe9
rA194n+nSO7XvVT2qMVRVPOaPWp73vKCUr9U1ZRUUxj5AibpsrVV6Pg2W4pS3PwM
TT3eRXrdwVPusQsnlbmri5EySs7ZDgQkHibfzgG+qM/u8bC/q2Rajzfz4ZX6SX4r
WoNJf7yAbayToXTK1lsVA3/28LHcbSqJzXOxPkhZWnVJ9hU/tOG8DNf6mNVVHFmy
oCqsXNmmlGMiHI6+Vett9xiUnO1E7BZ2RFtF2aMe9UnbxJ6OTsq3RXjiNsE34PQ3
DTrDi0BZEzET03X/PzC/J2g41zHs6F8DKd0zbfYQiZ89YohF5TbPlVPPSYqdN9++
quqSvY+Va5R3Lloyt+95ML6Y6v4ts9aJclUzkeZGro2iAc3FNljeORmGREIk9FGG
L0iQcLDsI0jkywrQ9BJMrnwVxikVK50tvDRFjbv2Ida/rvX3DAsrwJJsog17WHPC
lpxnR1KMzIK+EAToBD+wLLxXFvKhjftmUh1HKZTrwLqKXNbwOUhPUfhP5a/hVFcV
6Le6Kt/8FO6KHT5aVci4SWF7xJvixEScYUQqe0rutSBBNiyEf3fG4/sSkjRRay8s
+IIzsxPKotXpkZ07nyj8Z6JZVtbbkp2PQ1L9A01kjFBMCkLCSkrJHsm+Vs1TOKgf
f7keHxeO59GtpZsanLYr6ylYNHokrYPYKbtQMjDotauvxTk1Z/KmuvFI+AEaHI0M
rxZkZahvWbq47YwKLx5qxfrwBpNUjIgBhB4pnKuGur4zzagKMpHQ6Uo0oF5xpDPE
dOnACkn9jSqe0TAsjlqxz/3CkZlA10HPDHPAo0gyJyzHPUaqa2u8MnCogoG5NBGn
7Vcvb6CE7IRYGajSW+Pgy5NRrrzEfBfFBu8q4OhW7e4UDcIvJkYfjAy4SeSEVF/A
7V2I81XFWAxuDVmS8AyfQz6v2dDn+A0PZtNyPliL+LVy0ci/5viNuHs1v+1dVw8y
lULQj7Qjd9HRz+Eier9kB3JZNUhYf8mnLhp7Bx49SYELe+7VItTSFkse4UKFSX4d
3GFPEEZWosWHfp72zFxEl7VjvHWSSS2f+61T9x7OK5fRI3+Uxrj+iG3GMIjgnt7r
44ULKSDNWn1csDZWNpmcfPXiUU+ArB0aiLVxswkRY3IeoQgqGFEfR3YcN9OBXScG
hXqOequYlPcSRKLpZQOA/qZ+NDq3WlGqCd/FgukTZfTGx56oHfpuofnYy+L2jKB0
OXc28hugrH7ii3n5dlUeCom9eRwIUxhUjoO/8pDOKKHZPMfevedgXcnu05FrqdYM
hY2Cwk9SYco42tpDLGuCA2SNW7nmlpUWMVest7fJ08LovGCEAfS95E1+RJvtfSTx
XGo/fNyIM8xq8E+Ix517CphLmQgVnhswviQdHpFx4Hzn/mm8Z+/75eUnceJqgFIW
BodBTdIkk9RObNEu95ozmoy2fnB6w8NLyL68eaQLO7Vk9SGUrTUPFHFEUQQ6gtgt
QrxE4owI/Hn5q1QUGAIHK6v1jY0HTwtJnqBus+9TwM4x0oeT2zk+UcFnkoCyXOTx
SAX/xO5eJENFbTDmx5b75ijEeO5SHlQdlmWPPt/F5gLdsOUD24lKuoMMpuakvpw/
8wad5FTXeZOk6ZKE7HZMhygTokzV5FspvN7YXsdnPfgWXVaImY/Kz5NN9iTGEaKn
BKeTc4sgVc2lX9OFKi6VwP+7VWl3Ob1ZHLWpKYi/YM3+afmV5ZuuuPR+/XTAKTID
KtI2IAtxPaEbKwWTvG/x0/dJTzdZXqoCwibzB2ogHOmhF4P82IIYrcRcGbqcZX29
tKFzR3ij018ABt3w5kXrrplmoSOnd6YHByQY4yuw0NWjBCWF9mL8ut/0Y1dE27fq
DK8PGeYeAh5U+SDjbqujQoV6POlGNiAWlp1Kmd4dzH2QELdcsTgryQkSLBkXVvq3
owj7VFCUoSuMMhedhbvelRALDyAZqNOGMKlKVYLMlnSac9zyJjBfoPx0ZJQXGHx4
7lsTiStTY4v7OfDkBbPX/2owJ6gR9hqRZhOe9Ut1B6pDAwL59IK4fVqYHkZtgjr/
/L8O50nd0qLYGKn2ZZpgWhBILkMHFGgGes5wgKbFl0xI5LpEcwqUdJmtfJjheydv
gHSO5H/fo3xeaWR0O3UvNtDjaiJNrHBlbDyDZfMm3OiHy/486zzVYFI+2FasBNnO
0NL4CQL0kx554QS5IuExqIlvufOp49pxjHO7pmRl1cYM0A/4hFejkCpFE0NsXIeq
6iXA/05O6w6tMZYTYQJKSJdh11z6Cq/8d3T/BgI3MXrph62QZ0Cex9dU+XyTOO1H
3AG9Pl6tdPvaI7qG0VU8NQDFcVwK6p7wNrFsJQT4jOdEKztTRAyRCUI0VFljiALB
svWu0p6Wy0rueQM9LE8Ahu8UDMZ7qq8PosnFHmf7yEbIwhhdTLmvzwxvCzmBv8Yg
2osIswadq/w16D+Xp15COyASrWFU7KsCtlN0Jb7O18zo0o19geYGBW3o7N2Cb+5L
gMg9nJONEMxw2EDXiBeegzVWZmr4rLdzai8tpGeSMnRn74Gq04KQEFP9TQYSGc3u
6fCkmLif/C45A2VzKLLZ6FXsOh/ZFoJ/Ei4Db6o9c46Hnwksma9Z0WAe3UudZ1A2
DAb4r/25tfay/9IUB+/VSPLaIIqGF+zh3z6rgbcWrDWMbmWs2bG7eOAg6QN1XzB9
Yfm1nboDaJf4mef5sPrAHaK/EmFR3gfT0RPxXZ9YvvrCI65Bjm3IwoWF97goOlQS
NYFSwldj7Zv9c6IuhPcDtETaJdB+kO79wf6zjijFuJVIcWEQZMuKIcDif6c4ojM+
i/W7mHv9uzLrDNAIZ2jtPXPViADBrIj9blQMMygXERV8DExRbhmK454oq/1xJTON
fr8GsnaxYH9S7iBjdanWVjAdlRkVNsGkhMWA+ZKK9g2x4nhNgZWTeaLbg7bMQmyG
thv1uL7cA3ta3n/e7OtNzQ7t6yCJtJ+RRI76DMjI32KHFUTzMRljKgqE4DEb9O/9
KX28TScrJEsOFDOqER+6A7Vy1slB/8m0ktXgVWQTFp1Sw+yo173+9OlBvfPRjJWw
CacL5sG+zjohs9qotTcl9I2sz5s/6kJeK4UTyWkFtcGYPs+zt1dg8A8JDXskbyEz
RtjjNDjXWw2+Pkc4SM4SrD3i+HlASzsUQfn53dTLRbqCk6OPyWJps7xXK+MpKKM/
nmWi1yIMSYorF/xJWLOU5UtZ6Q8DBF6Jk24A1IyGpy6Qq9liuO3GXMDkizRg6rIf
2pnA5lNEFw1aea5BzczHcKZpoQYM9juhmAuLBWXBr4Go5nF4Fgn7bkPd02gbUyMP
FrsnV6oCGzjkqGKNQ03b0f98KhCbuBZbNE2BA4wfUjgrNa03fKAE3QByIY4VZwuz
ujLo3O5nyjc9mhxlUir1R/K5AoZ6ixCmkxjdJukrdm1XDCOaUjLIphvnjEnGjjb1
JwsRnI5QpnJH4BWVWp80IdmDh8XPTcnbR0adAyU29i67XomFbpUKiajfVb0X7Fnj
jtybqkQmx2gU52/K8O/NI1SXfQug7396xo4v/Na47GNg83XAQdiQ3jRNbbxOG7dc
NdnImCuwxtXaneTxDGet9USlmddHZqYPE6sV9nCUhufFcPpgEIdi5YMbcAYWEZhj
vsKwVZ4QSgq/bq8Ip22t7dLnMAM/8OQomWd9TBktONLUYEvVSX1SOU36YCZboWaZ
80yjX7fYsFz7qYvJnSaiF08Bd7qk/lVdIEmAvz6NEmL62nzcvUwpyZp5mLbg0tHq
tCbGrlddd++NOaix9j4tSkURnSr+QoM4e3qj8cVx6+pxXGrj9BFQWx3VxmFikUbL
3WcLQ+uk/KXcVJiiOEPjco8znAfBpESJSfHFaGC8mSYz6AzNGonqm1VHz3f4bISk
oRy8HjpF7hye9gDAwUXoe9XKAGC+rdMLq2iciH6AXs5v+S8ps+tE6pMNy1wgFfmC
AttVbvORSt/LQLy++AsV1i6czL0YU+L0kZlek+bXgaykbT6Q7rSfNH5VAY9ZM3J6
5tTlmja/5vNRmkzEomztgT9B2x+QVEGZjKXPV305FqPW2WFvdM4bJN45zfwee+0s
4FLYAuenOhPqWRmd0U1sSA/qPtV9GiNbEH7orJ85yOSebRR6sc00/dNbhRMdEv9G
llJuFKg5OLIdvWxbDXhs8b/gZPB6j936UMvNUGp/rpRDp3jSS3vSoIMWZf3dBxFj
ZRF84AUbmd0/5QH0otJnSaEp+EpLTBo34pOJxwE2A8oKFfLER8JCg1hqbnEmYV50
04CrLJ3n17wP/G/1whxgMlZqES6EAkQtL6Xy0sz7GfdGPraw7+OLkmmrHttrD5kT
7r6h0pAWH834m9ZKeE/JgPlbQtefzWesy41YhDIHqWU/BoQIxV6DjyboNFEdS5bX
Ic8ohT0NJXmr73akaj3mWedJOJ9miDpWwZaKGkY9yZlGi4Wakf7WzAydVx8vphXV
Akn9tZ90GOC2MwHfkZ942JShK4Cc/DWODR7P6zwSOyB0ERn6QgNbHhZQDNure1wG
ASkGVdKVSo24ET2RkeRHC6bS2BmC3zqwMgn6dv1HlXT9Ius9vn6jvZxLWHdgtN7t
UpqNgUemPlzSV/4qzCSAz1MWKbXDBDC4FmlhGw6lnOsctiKDNvMCOaK66XYJAvA7
z4dqlfwXxcT89vaERE5weNGdMnj8ZHO70a9upXXPzn92SIXiMlHyJh7VBMq6kVMO
e5ytrqNsfhwPqsxSJjJiBnJq6UoQJKIfI+OWw6kP7O2y9kNSUWsIJb2tVoUqFSmE
bmHzEsJ+Y/nsYclsQvoEYK6oCedXuI+JMCjJEw09y622DBYetWzM0oKQz9iq59mK
nMwfjbW3jADmtx/8yYx39rsGo5NnAldlzqO1jBmpmgfJ0YKCHI5ze5ZQ9DnSZTca
LN6OPQ64sKJzUhXahL1TG+iUyO9Bz0vuX3LOKqOfbxkOEhis88X1wLnQ0g9+avT7
yU8GRN45zr/rC52CxSVG8LJbnTGit/BzOVa6TW6gwDIA+7WUhbT/8IF4MCUmmvDR
n3SB7XoJfukoD7PgEiOWZ39/pfAaZ9hYIJYpILm1+FhXxDY2k6DT7vOvsndvSXcW
vxiPSx8JfEMx6vuYpUhfZecQmcOyfAIvNnFoe1ZKfoRf/FAk3qi+YesOFSbH2Uu1
4vqt17dytEK1PeBDLt2Q7saq5rGshaSscGKC2y+NPR9rreT1heSMDmEoucZIHQOn
ILZA4M6HIEYrhqRsnBh+Tno7Tlo3iFFebK8H/PN5QzmddW8ugdXhsUOqbdlLo97R
iND33BSSNKftR9jkz4g5gTYfhdS+4J4e6IpeJ9RKZFZYS0HUODakO1AI8geho4Oh
ymhlvGkCiPaQ3WujgFbkyyOs+PqbYCDloq0jY/5z4jAZPm1h0D3Wg2CWfh/5YVQ5
BYqFF6chOlwpHXCrUrQxc35IvI73WZxwmmiS0E6t6X8qNdhkdFYo1qO7gU3jPSrX
7IIoxTsbKe0Cjl0Rl+2BD6HoNeGrz9XUzPEowKHdNwTsKu7TZaSL6fsIgrwWugg4
HgDJRNlvNZk1A4iAho7q9tF1RdRiDHiLLWr4re4WxIUWJxaqG3I5c2VqAkvrlIGD
fQJVGTSFx7wDe6xjacBdGAdJKe4X1aiIBs2UltzWkDi9hDHttHXXkETTcrq/WmNT
yu0KeAVj1WrM2sl8CFoJrKic55uHncXJ9aHODABjehHlXdiSBD7z12o63geQ9f9z
KUujdgSUiM6BbTfGSN0KD1bSgGCl0V0N1vt+TxaR8za1nmn2oqX0SZubD+GoG4Gj
QBgncqNcA7EUjtwiQCMU42UAn3Oo9dmW/vHFiUjhYEXgdvrofysQv/867Zj2iFg3
sAnjXUFnuCvGa+XktDH5l1fWI3ind0OLU2okCI58AHHeo/uFvbN15SvUZqwzKcN0
ErmMjW1eenajIb65xk0OisqrNDZoBxkkC5cp810iIjkP1xbobuYQY6etgaCcJq55
4DP+45dyHrfyhkaIYotcyBjuwVdPo2NHjzChw7IP1WCJ21bsT2Nl8o6uzESqYDkn
zKc7zFmvOmd1bXIoaFOyVDk7+kWs/AtzWamQPBukIAGB5zgdlEg3G5mJASYHYezz
Low3uRPkBq5B2laJbIbletqp9U3B8f/ZAw2/GDcgS8ILo7rmOAoAN1ewlq4nefe1
uTdLKmRw/GAbFplK3F7azigy0bDqjXt/kJP9qNOCm9TrnRPK2NI4Hbkq2zr9UH4S
E05U7bfk+17UgDRDYyz/1zWy80I+ze1WfsVygMMpKIJw98P5dLCwBC3dBfivh/aC
b2KjnU+i+2sn3I+ZKxJ+WNV7x39BrlmZHJaG4BzkSVnjV4XdNjNPSd9Pl9CbN9t6
aXD3jb3aHaQlS1S+UEm7VTwZ+O25yhbYXIB9h13bd3VJM8MC/B26M8qLZAIzaiNR
lRDlLARkOqILkZrmR3fgJTQ/410+5O3I9cWW3jLgd43fpUEI/NTjYfYevk2tW0C4
nPiCZ+OFsgyNxeyoj7+PTnGjanpUEijKN99W2n6KArHCANp31aAnLq0uOWWImioi
SgMoMvKjBic743Zx2djAC05scixOXybpe6KNpx8UX8/yDYIeeEleHTZOwBmoOQkU
+Af66Hlev00ObjpG+4iHuQLrdoVObqGrEM0KHJhVJxfAvtTHm+dWYAp+/wJcFnRA
lMBA+8GajDl9yhVXQwoZTMtoc34V4k6NUcyYsp8mJt07xJtJUWcZQmZwDhVHc8FA
sesmEho7hMJimXN0XlvVhHgo/9XKtSDa2dvjfWoJ5um9b3RpSDQN1Q2H38yGXERk
GLZaAHXCurNXefbsGmNxjTwaq50U7OIch8E3EoftSYrDTmreR4uTiFXfxX/xbkvH
YE0UiSsHXTVrKWfH9Nz+GMSe4WZ2peJPBChVCoK9i27bpBf4BMsOr6O6zsFFeaeP
geBpXDyIAkp1FE/kcT+ay3HLVWwGAlISHOityaNV8Adn21dBT5IR2tyVYO6W8FO2
1Q9NNq4gY2TClwG+x6uTfUM4zbY52XgQSj34QMu0lkhCoRaOIyZepbLpuBjrUMbk
n+zSr/ggbq9YUOpem2aET4jzMZlhccUQN9Poy9gMi3cNInJtbUGGMM6FuNYuK+FX
/jlYasQ4XV/xCguxrYOcKPktspJYq0joeXEFNWrSYBBucDEw9g9YKCQBA5WgANXG
j22HAJOMvLW1RJS8DM8tZuVDRiJep/TFjbR6FqZPd+aO6AD7lp2VxtLcQLYPdkd4
1fp1PYGK6QNY2HiyIP/p2HiXBB4ia7koWg9sP0QVl/b4nEwkB++Dix4r9+QklG8g
NiTaPcecpawruvlPQ5207ZxETyf4EgDye0RqKJXBUFqFtUgDuiCISCb4A5FjUyzW
jsnW9FrXl7c9Bar7llWd9tddGCBY+8/uEnD5OIbJpu04mWzmnkLEm0t1lS2zZyv7
sYdVs6nHUENA0LGZNj70SGo5FzP+8N6GQPdSK9BF5K2cJpYbUgdniKPcDanM7udt
V3xF14fvlBetVshml4pmVi68hBA+T0WuoNCgu9DUO6e+lZx+Ns5wZ8K+KKpM6kFC
1/+Kt2pxAS95PGm0/gHZ6WzC/ioqQm1zGw9QKKpv01AfiqLIemqGfj0eFxyqGmJO
a3iRj576WzPekBomw0jt22xLNibAkOtZxyz+2xmp1JzyzaUTr33tLFC5Pw2o57X2
nownGqvJGV2w489eeD/waeqvfTwxS7ZkLglcKkyffN4A3pQ6oxrCImh0s2LzLBf6
Qj31LWR4Dsa0N16iQYey1Td2U9NLXEJV2Hlsj6q9ByS5A0XqfjNjDseZp0Fs9FSr
A0OCV9QT45FLmwKrMG+VmPZiLyYWVA27sOgN7qIt/9FDX1kRJ7XOPUStXJ1GhmY/
ifhj6FKjzeVcctIUpXkA9txlQ/BeU7XWz2z1ZoHbjeHDUeMzOEwjBaCA+G4pRxi5
uknMEmNvdmsf4nfE4Lg8xmtOaMEItu+3BREE3DVnIBzP4IAqJGgjz0fIfXXlMuSN
6A0RiFO7g+SBXf/4xQQsYCEnZk72GlOB9eljxuurQHJG8vFpXQUJtJDKfSUV8qHn
qeSNQgzYp7Yn0xBFcK8sMMfEY9s/aalSx7yBq/Lwn+jlzPttvjl3Sjx6fG1o/Y7z
F0RBp0T5FQbZiC1WUCqf7ZdpXpeWGKPCLe9oj88xDUZYMr0IQbjYzc+IeITGni+F
sW+PrXdvhG7RrS2GstJPzdB2/M2iyf2F1QaVlz3KgHf2M+5+8Z2VJ/ZRKNVBnm4v
zpgIcom4dqd/8Zds25lN6nKJJnz8gSRPiw5AG9vS3sItSIq5J5fGMItlAlGtgrhS
O/0Q3p1zBRgfJ29Cw+fsdIBldj0f67W8Y0F12iVe/LsK+3wfCPYRKS4fEd5412bO
0Lea4x2jB49gpt7OBrKN7ogrneZ7IV3TutvwKjzz8A5YOkyulCixyde+UfmEzQsL
Z/PJ5kNPaUA6qeJ/JnfSwPSHMAnoeb2UmLp38i6LhbxzvcRB0NPjQpglF8opZL0J
x3lNdcOzF+/Vm4siaabZj0Mlq5gQHIkHh9nNg3Yf/X0SA3OIIohWiIiMnSOlfA3d
aiDcr6DAMO96nEvU4lC/dtvRdnWG8Gew5h7t4tny83nAwqSYYztPgr9cs1cqLGCV
Afp50vbrpaiK6HUuIRj5NmYi0TGRLAj01HZXInU9KSeFHO16pIOqXIkjVKzpKFpd
fBtIqnGTq/ERhA9PWpCLP8YIZ6A6h0gYdnU/NDjyDnZbS+K4JttgXaEABRffCxCf
nYEO4jTAUi4Ik6UbQsWA0bNdpmqj3AT5alwGAgeQ7vqaApISnnuz83mP4k0WqzNH
kUX8Da0AqpX27vK8QQF000ZRJHHmGGXScdPCTUIXKRtj/YNuTB2R1jfjgK4HFa60
kFQXHImNu32FhLh5baVCC2V2CygTfRoiCxbNm/cbo+h+yVF6QhC1M5XPm7HhfnY3
Rj93FgAHQA9JxUIgbMNSWbcABg9hSf9xyWh5bvh8J/lc6qAd7Pb2UbuLtFwK75VQ
den1KbEnEjykfhdXACV9tSrG3G2d6fx+SS/NNOnofnKSB88wRRJyGmQuY+ecDaMK
c3ZUjjwvlfdJ/pOWKFRckWxgTb565Z1rZyeuRMX17PpdvQhXbzQmJDCFjUatQHYo
jsP0HMkMgT3JYasbjv4WRGuc5Yp5QGoAbzKygALMFzZjYBY+Ekwp1vcr84c2Fjh0
X2ujDztJvKM6Sh3DKzZCQi8n3WOL2Qvz+9xt2X0X0wrigJ/0Ob0i2V08plJTWydM
eeohFOCHml5ws56Wv3FGPk400ijwkmMChqXvEItk4buAWlG+lO0uqyYyzLog/w+t
+AF3ZdvBiolcWbu8NE+/2KhVTdDo6v2OIe1XdKITVWrM4MNjJvBmIfXrBXF/al+C
pGyxmNHkUWa3/QS8G1qPpCJTgoDKRsfLtOO314Pn4KY9Oa62cWNVs7vap+kYE5qf
O6QZsG/DnTFyVxVHjm3a5NidVjtw0ht9aWtsdFiCmDWZImpnN8YHaXS6e1bfqYFL
PEqJFfDNy6qZc9ceqL1kSSGWPGrd1Gv8dMQJNOt4X0rQ9tNLTpqO+6po4uDTX3L9
onCMyjmA2Y735FH/dSEuK9gMV3rRe4Lk1OfRWS9IGPe35k7EFt3v6X/YDhyU4qZJ
9PhEwZk+NY4fxHpXpoB2dgVdLgmYCjAvxUDHjT/kDals3WwXj9OYFqQF/aIajCmr
bXQX3AQHbFT+ZaEuT2fiFCaIist2FeoEO+pSVgHGQYOJXPrl31ZoRnJKPpjc/OeD
Ipy+RQWX6kdZO+N6e6Nnpcl6L586djIIUPokjaP3f0ixgKgRbge/GJVS3a3oVnPy
KW2AFktKTfhqWcrJXLSDXY1z42V3CTMz7mMiVyJF1cFb7FipRSnd6MRK3qR4YVpf
7VZGRBCsQhkaQ8E8DuSdq5UW8Jfea08s2EkP8VxIBZyJd49mN6NjyL2lGpNVNfao
UgoNBNz1DZWTht9vZBYnnmO7Jf0qpDFxHhYGLgnzlUqdZj/6SuH8XyULSL3nwnY6
NFyf1VAa+YEnWuuyClf2rJV7OIzEbCRa1sQHzSZ7GS7QDTLZQQqzUC5jQxVyWC9Z
iHfqtK7WpTOg/bKFRIQGg5kLodRfX00yQUkApU9kwSD5njcW9Z1OT46zadJJDBeq
GPaQ6tSQx7JfOMQCEsZVhgXaDLz5g7UBZ259fXp9KEFAGg4OIf4NtoWtcTsq8PX4
feATJ8i+0y7HXz9iu2Gl6K872pTMfOyIng/MfwXmRq+lG6Z27gDmBt5AWtB5Aw2v
LFV9pewwUnxG+wGTZtrBXXiX/yKE+wmz2GFYv4vgYxMSwWZIHNtUBqWkRWM/O6Pn
NWmpeJ2UdWaypz47KeIwGvbEeZwPtgdz3v+tOv4Swe9waGeR+pMx9MPxdlX/IhrS
1tbC7kpsAkOf3znoNVMSSMQ3yR6m3t7SLL9ZlLPL2guYmbqCFHIhvqelO3F20g6k
iQjmstSYSXnfXuBbvFWnIK70WQMtTH/CEm+QwlQLzBpWlWJjlNp8+FMz89GOUPN1
w/DalHnYd97psIrHMwombzf+zhE/gE2XijKnxFXhpaGRYcHXWYZc3mtu1nynNYFl
ey54RzFkhAB5EApeB8wC9EX5as4ovw1ijI4bFvc8SZ8yRg3i/5QxEgY+/EG3RrO8
6lvwxuk2e0TnZUXonXYqHucdkyUxsoozhtp29MKTRbp7dcCTJK5WyoAqoMi0ScGm
dzarfcZX5uR4vQFWtlDncbBlVhnB11/yWOMHouhX6jEhbn+RvKfBqZ3bnoCyJ8Ff
+2E6WfT8U5cNi/KQwr8T9qyVDSUy1mH37zsI7LNfm5PPk5o+wdj+bUzAs4ayfruX
jMYM83rYuhZDP6RCqct+ReSKYSEOewDlqgBZtBHXvzeS1+tpJK7V8Ulk77OG5cLk
cWDgrQdEVWWrtjZ1F9zwhpQ1Yjhy5SnExS80OUlxwomNTEE9aR8V4xsuqd52goCs
uGVN8qrPm0+1eEGkAX5LSF2rd1Jau5qfeLMPu6DGJOcU7QHCjf/ymG43/r2CmIFn
ak781izWj9ff7Dp90LV7dRgCEx1CppKU6UQpAOjDTpSH7zywW8FzuHctvFjsISND
o5Vrc5qooHyX8ZyO1xHwWEi9pVCFsqrU9KPGTMM8H/jlDbmloOThc72phG+Ch/43
ESWd0magBHzorNdva+2ZgMafTlSIEknkhWtTvVADtz3QFjq6DipW6G5yrFSNBIAP
rqjZqCR+1w6FqBm5BtNWfiCk6nlF0uz7e1otsEW1YBUy1LUZIhJP5R+GnynNX9u1
4umTkW6Z77L/QTceFQZWPxZrpCE4bKlRc1YMf8eTQ30ofL0so6LWHf9oqLlE0ZJY
SN5T87QkuIpTLcgnlNVkpnNCDIkqGMuCzczce8rH39q4f3PZtb/jcH5jmAgFLM+3
bVCwZWETwz6yTlWh/9txOQnxASk2VEpPid0zU2sy7eVeiTL+IBerKDjLAY3JdkT/
bn8wOE3G/e22LDPE7PFVsWBIWSY9sR7ohE2F/CAwuguFFDUfnthtVTfSZqMLje2h
H2cphrmyfJ+W2VxeecIyqd+3bPlWrQTRbDX7pXQykNj+3Nx3d9x6ek6SyPwVD/Ok
pHh0uiBtd4WnTOEuDF+vecIlRowKLVUz11nV7Ho2q6sPIMQIO8OdDsBcDPcm7pYn
nLeolTTY2On7Tuh9Kr7Vyc39me5oJl5yb5SrBs5dwW3sWf6CZUa6GTivNGV4btjv
nWjPautYisOuxDuaBXsfcbyCsARga8Gebzvg2WXuYf/1jtOkCReeIaEVoxwZLYNJ
9797AzozVaBYd6FL9aK8G76MhgZdxMW8+nMgwmWfjSIGtZxybEco+c4uAv6nMTZ4
08ac/8+BLGi3BAJNlydUwa7FElQt2NJ6CVtXV7MzcKkgPO86/WBFL/b5Ch1TKwvs
SlnJuO97wTH0LkStAis/0wKbQEAFcXCyxVe3iJusnSvS8Kule1RYFZCr7ELDI0AW
Es1XkEh5YaolAUz3FnCv6jQNTVwfBzlFSijx9idAUhhtfPXFBWd1NxvqlyZEanyw
U8Nt31pIzZtEt8k9uIwEcth2QsKnZv9iwpuMnkCiRev2JAlTkujoppchTkV15BHD
fB5RQ1etSMlocmcWha2StD63zdiCuGAdo1M8i2y/QpNSQR+cMbVszO8IFL/ploTg
74gNroSotn+wJdiCPsKOur60LiD7KG1ZcwlYYhbvEApibhgJHlah2LFPl30g0LKd
kj8Ebn8jVGDIBTDF0CNnfVPgz17wXQdj4eMtx9ZKViauIJEF2V9tLJ5R65FOnVZA
u2I10/Bpg9UDCY4YnWiutmfncPuM8L69qg2b99hpooGKTLB8DyeafCq2cRtSi8W3
ASbL854Ns2yTXgiq+eHolhjSYme/v16q0MMFN7fzNuPeaVu8GuRl16MIKNgEsE0X
DGOYLKWrMQIk8uRGmuZPS8XIRPSQeDZJhPy3wEWMD8JK8cN79IsXTNhoHTwwgwyT
kA0W3VUR03Ro/TPmJJEuvXwxM4/bLqZZcBK92hz58zeYlnn2doWHAFZUUdr0WAmi
gEoDLgT3FC+VKpO5/uzA3cCRUayFCCDt0xt4gJ+gYCcKWqErwCJ7tHJHyChd9AXQ
6+ykCaIX9kQDlf5Cvz1jHtCPJK1+/PVCGS0SozDsnwFUNglhf/L0d4s2euWsWpCh
voiJrJKHSM3730EUETR9ELXbU4ZkFu+C56QT8wAWL+Euuv1oIRS9eWDx/KmxZxob
b1jAZayKTfkJeLK6KdqKo3XTr5wpw/T34XSCRZcGu4bWtg4QjJ6ViqkLkW+XfFRi
Beu2wmNjP3DYrt37aWa/hhyUED+E9o153GIWvexPGgj8k13LJo34q8m8mw9kb4ou
l0ihcCB//RqroTFgfg3Rpkack3W2zk0motlLrUtbys+PPSuVI9JdQnn38/2AhP/V
y13UTYgqco/JYF+LrZXSAQk91BmLLKJCTZd8SgqcX8sBd6tFq7Q/LUSXIsjFMNcm
+huwfcpZKnWfnpUBKyR7Vyqb2qTEg1l0g2Y0Sfm0tEvDNvkKFjo257O9g6kfmYvL
9+SsyiCX5cuH07hApt0le1xmfbTT6CKdbDoAjct5KHhXn3ObtBtc2gq54GJBXWzA
NVQ7y7Yh83RUINk7ytyGp8Rabv5f2MV1Me7nJVVRlEJdwyn1Xx/nzZbsLN35+IAe
Joi75QwaXNLk+KnV9pcv/XdEvR9zCbaHu+D7EQ1Zdgo0Q84AggKu/OmsycSMGNGB
Ji8CgKnFLyhL+cdsWS+okTMVV3OTnQo8EMoqnS1So3xL4QvNmUfBLlqmpCkMUkiT
u/VVg3HwUoz/IEwivIwgAUl75WSSAo3ZAzs8BinlnX4n8iVEHMhQIv3m3UXbanBb
86TokxByIlPz21VzYhys5GUKijg1J+ayQipAH6ZUOqwNhLDitnGou/qDJlpjRci3
raYtQ/6UcGSHKANzyH1PHSMbqTNGsY28sabNlWcaVqd/RfpJBnD/u0IKmnemzMio
Mv6pLXG1C/KveJ429kGQjfQykQPyDr7meTRrelbSZhyZAwm8J8wifY912DwUztXk
JMNdLF3owt8WFrNohJDldWFFpDZIy7P3N9BIBRjy6EhkBAR5csXjJzQAAcDwL7ly
Bbsqs59uIPN3MIieMAMaiLn/m30dkAw9ypxa9vcrGF6DDqjavWgU5geOuLSiA8/E
QAkGS9Y9vwf4QOcHEECKpLkLE1xwxL1Fjj0X0VKxgE3lSs5gS7yP3GAEh2fX8G+z
sKsl0qJK3k092UmYwn3hYARElA+LBIU1mO0BfKYfDwTMJK9xgt/CQaGAEQHEaKpj
OxYpxg2WwmtnhhRw0scfn4CRHYsAk6kQAI+dEVTy0DhJ/3guzYyuxmA9bChIijWi
slBfr0WtsAC18iU8T4nNWsOCleuw7mEhhjD8TbzzMviZO+zoM+cPIp6+B7B93yb3
pDIDJc+C0nlxs5NxMuH9ZKWGl6x9PFAVCZAUCo4RGzyl51HKY5j0qL1CQkSqaydC
O/xGUS0Xbk8h5QDYe+BfulLBBJl3dG4v2jLyCV1iJ9PxB035/VQBedPlRybUN5lw
SwAHXQLgwsV6S71ZTDjeJY4cUXBRrjv3K7WitCRUDsADEpSShqQT6q7sJi6ud1+d
dYe3VQtVOTFY8oqWv4jZ5dB3/kuaDk+1330F9Xo1+yhSfy0VRqE+VBy8t+fgVm8G
ubcEfhcpExp2gUros+iaiVGidtil351r3SKPB6nGqck3ARPEalQzZgG7fNEagPIj
Bpw4MKic46R484lSMetdlANr/dPxWoCczvdpCnZ88zjwP7fMGedT1228FBGRO7oU
iejC47WYx7e0Su5DiyUHMXMD3eppifgIn75Bt5VFGvOdDwL+MJsfAIRSPW+uGmIi
tzkF4pvamqtWpBW3YU6QDhqDIlKiEXFpFnoCEltZqaDQjL7cZkzFjDdiFa7ejuX3
ntFfJ1rZYuItWxE4ZQHgJpzlX9GTP+8GHyWz31G0TMyYyfRkghZ0z8CUl9D+PxwZ
VCPzCqrGLwW54yBg2rhosX3Ss42ixUVAPuvpIKCohjZXn8yvJhtsNNP26Q6Z8E50
tLRgPtlTTddLJI+PWxqhg8ygl6wVl3jT+vO7VLf/BYaNgxPDKD6OB2aAtrNiN9G7
URcV0q/sdfeHKfT5S0+T4CaVruIcxw7Mds6lTYf1UXDZJfhES1NvLG+atSy884OG
13B/iCbDg5Vbkwr93lYhXjQqaZZQnd0wyNf7vybz662Sn0ImhQw21ZWsgw/QpaFS
Nh1GShlPTBmHrMovWUcs6/rHeOU+Qp1cXtNKNaHc00f9uw9alz4swQTovhI7Z7Kf
YFDYt60MPqSSXpL2rnHKwU8cwqpRR+V1MQqOBDXu+oKgIzbzBgewPLwAr3inCOl/
kEe4YnEbwoWXenWxYcz0RjQsKEkrDdR9rHk3uJNPeOeoN3UTcYORouMR7cHOsiq9
1tTODtO+NayqMM/rTwOxDJGztOj0Mb80uoCZic4XLjAqVgp2qEx9oV/Ml0UBKi9h
mt+4RQ/9lkEHdFeQlFA1mlmBSUH+ZBlp8EB0SMRc2XT1/Pqj3hofgBg6xJx6MZRG
bSW7qSH1l98lC3TSC8niTGuMJuxzRE6n2md/ycCYh7DJ2ZpJnKl32yP8I9zQhmAi
IPrgUi1Kjz3W12yV2bRNVfUVzMrEn5kPOk9utbPu+6u+96kXCEtF18qv8YCnWyfs
LJ8D611sGP5+OnclH7gQaDubrh0joyJH9KvfJNAVFUtx0JFRM48q3ZlCP+rrjIGb
BWQamY0tlZYc1dpr32eqfb8usggIQt5/8wZX9jgxJDRMBDG6ohrQy/sGswBfxir3
YwoJgjwhip3K4e5zKpHLg7Ib+egWpOjpJHh+WMcDGS3wvnvI5xoeFDek0EtevjOw
JDn0Lv0HwsRFy7V39DXa5Q5CjGkrI3eFlVR1wDFGVSCGQURStZ05+bnfHx46ncWN
L9C3sI3Zn7ejwb201WALhL2pfHv/6qnoaeuR4TGgd0kGx58FfQtkZbkO8PwM1o3J
A3HaSfZZevfFC5hPoLpTp4TI2RyQnXzyU5NyFH8PatjPba21cVtqkst1qi9hYx2l
Hv28vwoJBpsgyCDUN14Oz6yGl9S9E3mBBIhvLsDZPhwKiPjLzYZW4qhUeIjYuK8D
mtEOOyrFzXDvG9uZvMeJTmSrZYg/f6XrFjJfYy73H3LOD7J34ryghvGQ4gcdc1Qq
V7Y6/AYJ4D6O9rhXDM4lzjydFvzIUrT3GJd529xrt+/w/m0OAgrQGpgJ05SJwpxc
DvQWjvReRB9eFGDXGB/msDVyDvdaX7gHb/hVp18pkAyf2nbHiGaPIIbnTUMdu7qH
VK2exPrDKBs9BQsP3GCWWS8pUn7vfHd0MIDFIv2KSxHDAjJyqLOM/d5SV9KaPjDH
0NpHB2hVTfJgyhWAYG6rnmN/dko7vZQ9v8y34OXIiT8lm0RT1Z39Vg05pgSGlnm2
NoONE/fp4r/or+GhQeZ0z2uec9ORZ004EJajcDA9k6G+EwrOq3aeUuH0l9p7MnG8
fvFSdl8cD2JISlviL616r/sTSRn4n9sJ5yjWwJgThisqPgjwdEs79SFhwTUFYaMg
K2rXyJOQh2zSnlpEZtZuI7II/1SjfrvdmL4T8QEXX3SKK8o81IoddM1RnTxXGsFT
NeebpS+gpXrni6MyA/ul2m+cP/kgMwWA7opfSfU3htZGOM9Fa/Y70FrXOOXWMFda
MRbVId/q8SBSzFhTUVPijQ8ryDpjKqng176MslArWa2vrfjT6q7S6ULdco09K5Uf
yU4ac5HWcW9X5hNIeltzx9vnZO0OJ0lEuYBpjc1//7wAR8TB01DtnexXfI9d/IlE
G4pgrrWaczUOqC+W/rNjed3gjpwqEW4y+kwZvzTNjLYh5ZtaKQ3HGjA5v4xOVX13
wJW2iCYiZXXMNFbu7pkIKj8rw+cqudMIQRkZfSYHGag30MFh1h1v/vjWWXXT5EBZ
9KCoZRkbLPioEUs9l0rrsr3KcNL+m2udT71zZzYF4sF2GKiWK5pwKcrMfYL4HEE1
qrDJvS2tzDDlIajBlCiTdT+i1jMF+ca+EGB8I851x7dPnOQ0LagmP7jbnICtoh3l
red/KRhA3QljCPlrwffyUTm+e7BSFB6+GHg+8tiBd+0CKizJ6OBNNe+635iT1+tV
LXfOY9NQ7u0xCw4D8GWhR6UQxerV4j1MXM6q5BHOXbYyIDZpP6RglM+9wUMqYz5X
8ylNT82RQg1lWUiXeVSP8hqdcsYcM0Oz1t9V+OZBe37iVAMMlKCtF/R1U9zzRauA
Q43JobC8nGdYkD9SO81Upf0iKk8vbY6vsO7vVbakym808BZOVnFCU1FXQsTcyCqI
+iyn+4X6QU2IJ8JzZsoAn4WbX2RC+L9cBjMdPTP98yX5EPvOla6DVlysmv5VvO5O
qCoOtc3rshVr8ClnkByE7gzEBhA3RrowtII4yKVDcQ8fqtAIJ65GJ5JHDLPWoLli
uvgz6z7zohZT/U2I7m1gI6TR/UylgqENgpo5cSJWOAHvLEAnqhpRcwV61X7nMt0T
tKkTjikJXHE+hWkweR9xp6KMBhX8hj3s6qTsITQKZwkFQ5tulQUmihEi6/WTOtlZ
/gotnBpqmp7/8AsXt7IO/4ri3CV2vNZ3+zmxlnLphgIzkVDh0HZck5fFHnUwctxP
38D7pVv6cbJKiUpGPUpkvmwGATWN25myZAilcyCrykwewxE9bJx8MsEKd6XEifDa
myKBNM/XnUsKFikt7fLEJEclW+8x9+qiDowTlGulDqwSLSO0V6ir7gViUAiM50Hc
bZ1IIkLi7CgpIS5l71MotVLzLDqV1Nmdzgk22FJmsWYFY3M9getvIwMuU4nyP9hs
ST3OT5Tpa/IOWlodILitkwojDGqRYLPkN8+2e/TfxfCDPdANgi2+/rhJmb5Katfy
J+mrfxnMfvOX8mraKHxwb14IiJgIKruO7twNEz3C7mk9k7SX/ldR079ZChDf2rtk
N2H5dN3OnQ2ULemKKPJMawyoN1Ufn+4bx/3uOH19MCfUy1/AEGOm5XjT20lG2bvo
apBRvcglRND3ng0/kYyUO3Jemi7VJSQaOZCre9wtBO7NfUS01WqkzHb6tnwzSxDq
KY+CR2qmLTimpE6QQuDAO68YnnALdcMh+agToVRQIM+Y4Jk9ZdawwaNTFjQtZdhY
DI4Vv+FcpBwJzRbmRpbWFon5H5ARG2JSeidiGjJ93MVIcJcVawN16KvXQxMvZni8
M3HJkNDsRVTr8CMzCrYMGiJ4aLO9ZrXZMotjvROVS0P7EpUFa3zVIU2qq1Lkj9Ms
HVjKWy66bElC7EVe+TQPpE/S1OiEaVnZQTZHDtai+MJB/M6bBEJykWEXtjYOroIp
KZ2+9eIKLmqawLyiWiACLsUsuEnqTRCATZ/Ap+dQkaIW7yQNVTy0igwA8owu17yj
mSYf9bgQ755n37KZC7b34ylan2NpvHMYtrNChsJzIWbmQNlCUXHvzzY+Q237AIEY
qHnxDn6fTPYQUjVhmtu5xNz0qrO4W8cEz36Pd/s+OWuHrrpQ9A/xSY323KsT/oZ5
Q547MWpxNMIIsHnCmeYYLoX9Izcg0sFB4vB+N14LlZUBVJfshC7nR3/UeXekZ4MY
nlzVzTyIbNTRBIHcjbxjzbkyTLbNC35PLMdTyqGQEOJfJQ5y7nHUIWOdj5mvmiiY
lOR+ko2HAwv/KYNZL1XL+or1JPbbxHeDEf8QkKQnINTkwuQSkaOujnsa2NpLrMGk
VFFfVimJ/lbodPsOcJ5g09xr2/oK85pGPyMyEpwHAHOvZ4VYPWVb9UIVyY+7ZBKU
a86mYu+aGSBnERD3i/7Q4Hgc/Evgk9ajdqpOFVYjkWGxy7togpqsNqFQxtKubKlZ
VuYiDHaBnkQ6YesfrpoD1d/ySEb4S+xX9QyQL38LGsaHA2G4ZFvp8vARGm6KK05I
Og6wz7k3IxW6usqr4pEQIW5pdT3OYEyvyZ+NBiBamxiL9F2GAddJeYX27cGBS60t
zwKq7I4ABXRx5h4h4N0zf37k48gtRdjQ8w+eBb2kwxFQdX5Jyshil1dP9n/RNNE0
XtMnSUY4g+ibGF4thnXK5hMn9fw+R0lHbuZXGUtSQLkRA2Sg24PSGMDnrNMLiGTO
3eoNgBuVlNi+JNurmAkibosNLtcou7c4kv+3XX3rBzXsfLUdlhjbEnxS8T5dcsbH
zKG8LDIllLPm3vIztq6hC4QPZ4x51FDKcfRxqbndw7nA2/mBBCaMmJ25MZBFxiMh
EHD3/wcQvnPktDtLpM0Z0uI95PQr39KxzJMnGP/55ooAJbtkYp5/GTRKqhliiGzn
Ba3ne3pqW1Mh8GVIz786lv8GLCSbzVGHhZYQr8mxj4sfkw93Hr78IFPA0EGBRqaZ
9K80n4aLTLNvRqMUuV1evTq8pAlqscIPvlVP0XlyiD1tGaFxKQdIBsuIQUMm/Tvf
+t7bLQ+zOdBJQo23hD9N7RppXRnM3rZ90OFc6Z9fv+KLRIKIEXoa9UbqHsNGYzdH
fZBSHpkOhSJN3QXHJ9umR8YPeR+7fFVkBYpQVXvXtEMX53ZftnDW3rvvboKcxfdL
cwFuJtI/J26YRCXZIdW5CsvWEzItIeMWDMXVuHF2cb0auSB+NF1tsNer7w9IubbL
Pe7VNSVUiqVYIrQMGv8TZMo17Js/dNV7liobONzssXk7CNAAQDF9UJvrIOZxBfXF
P37FMFq57R2KS+8kg2DOt4WTcrsxnoHanEHeIKeDBPSXYe9KbQL4nX3IAt/V2faP
cZNEH3f2PrOrSKC9KK+78fpUwUxGFKBuImyOnuy45RSRzjgpZ+1/YpkD4cCqwZrM
MoW81XAczHZ6hMcC31YK8JjQAfu66NG1BkeUfBF/Y0SP+U2irsxI9w0wMgn26sVr
hYObLGa7VtNjuQi9SsQUObGT1kGL9+r7gG7psVQuOm6m1wPvZQEbyiAKU819r2lG
Bdlec/RIN1Qtd95iOwzuqGJt0gTyuHZHEl2sSqAizCOEh1XbDRcqWXjBJcohuA2t
Cucrjifwn6tXnxxX2nbEl7SgfsyYHogIL3Xg4zM2wS+0VFhjDnBqUe56tVD8Ueye
iFmGFDxNkR15bpa4JaB+wQvqaJki1TiTyGd6IvSAAINYsD/qfU+Zs7xxNZLhd0y+
4PF+gDFwzpJX9wo2FtRjB+5EUAOv4L7GrLLdvufZTeITBuVrlB/EUSxJc69yyvtq
rsCH+55OwY75WMVrN+ssWoF0898WUd8th/1JelNfEx4hNOeawdXJV4MsSpjAYmUX
03GiUHofaWcg9A//G6KC2b1M2LvGr/E03vOn2Ga3ylaohWASF7vMOUW9Gx2CtgdN
h6UfDbpDTXo4bMedjj69Lb4umZSKA+1vY3SBbYOP879pLcWq9He2jTmP1HYX72zj
kzTIF6kdwnVqkncjDuHNb0ZjMaCmHw8lFVKyRsruZICvL+vEchULlCoy2GeQoI+S
ADx0De9r8fpnNzoUexE0+iIOjjNvW9ZhnKDIDAFSKhpCq0PWOQ7CwG/AZB3uw4Zw
2UPi5364/Faq6sfufyOjeqh/RXrUMhlv7Nfzig3JJZRJGu/6on+AEAbfym8SFRuP
PmGS8fkpeu6ianStydoSve6knlEa99H2hxsOaz9zmm/3ssfwSrOhwC7mHC8jVzx4
ZREWZsTMl0v2cTmJdKC66MXHEBWTQOsSZ1XLZ7C5GxLbyz3rPMDtuuisFqtSTBTh
EqqK15+L8kekQFux9u6ljz+LYjQqFiIeGRrYTURNgSilEBiUGrdMMpFFRZz9nNwK
qbwd4e3V0q1AIdK9ssFjOGG34xRGF03hGji7rI+7hm3ajxyO3r+kZiYz2An1OF0B
bqah9jINFNwsNheLm9gcDgJoAaxJ4MFqmagJERESCxfBo0oz16qqEs8wwTzV5Nfp
XjITlNbNA/dwDtANNwKY5hkfuPOaKGwMCgF/2ONf1SlJi/AzEuKzP1WO5gtWwP7j
UrNN/erJqq/R3xVsMjY/QCfCOZuTzF4VnjZJ+kcn8VvnrfKuc51xBbEYwI0EKkK/
BRNh88p9bRi+WCHDQYxHkgoHdZuO3HBu6Q1OPWJ/dgO64yqDnlkbHn0qjtBi7xrB
IlDFxFEh2rICY4hb4kRK3bPmidTyrIJVXpVowFI+S2MX2APtT8zzl1dgcabXyxiP
tOngR5jLAQaz9cnSUEh4J1VRBLhJEMt2FoyPZXRmWz4qtF+CzEUMCEQ78RQXpf98
lwalzd13MVxderKhvA/d2RvBmaLtkMUPUPKR1Uzx0F+xxdq6X3Ld3K/pWeK6alv7
ScfdTdHZ1JCp1+sjvkarYFIaU4gEWUcEw/PUVI5q881Gy4SbDW/yb3rL7aER5Mfc
aY2mbrStSgjRNsd8JYqSLSpZUxjtxXThnFJRg0GY/8WhKbn9Sv0ctC4ZUaFgb+W3
w2yV/ZSjmSUWfK5MUmG+Y5xqg0xAmVF9ecTfpIW9iClczzsmVAzbT1p89ge/KuBf
uJw01lfX5jjelDuIAHY89cyWdfoLt09r2PLqkZayNwyvwiMCXSigHaPTTNwolhuI
NDvQiKpyEr16FxE6yANhNIHSCFfBqzbaU1oP4Y31xAibXETKFf2TRMZKqteugPAj
QUDqRTevuGgTiCk1yPHr/hv8OPOzWN+zKhfqnoNoAjwMvGbDrrLFXK8F1jpBe7RA
HgsWYCj3b3MsNcilpDfCeuaymbvBghPxn/987Sjq12DFUCynXlpiSFcgl4UPxkvf
cxfIB2G5NACQewtxSMBGYQWnJEUiUswoVIkiD17+i9jjzj4ltNrubxenH0D9FIWC
SHu2TLweloxijNvUJ+t/Xkk9NM66YKXDyfRqHxd19FLH6J6eWX4wW0BhCm1CJIN+
Hz3wjmXtB2JAwUtHXDgfjle1msw20ersdZAloaWgUDKFksa08bi3bv0qfMfvoA6F
NChM4nHhcJCghUKAjA3XUouMtCHxql49ngQw0iJoi5qzrLxKkAyxHBK4PJl8JjWO
0jbkuH9Y9J6tttLx3Myl+XdsZrCRVhFPgFBCLEXp4RYtOq+NajjiICggVqjw2VjS
ZJucrfPJoO9YgC3lunEF9b8vIszmwJ5+g3PNL87yMpfEl2AMFsqjrvTvMGa1LrzX
5JB4p7mpcpx66vysQa1wgp8AHGImIoeguy3a2eR8y/oYyLzG0dM0uBV9AgZ23JJI
9DkKQYAaM+aOV6ajwRnafOs/ISWDdnIm8elf1Tnt7v3Z6SNpn6sCSvFEmZ+ti2To
bg5l8QKVkl9PmuU8pK2hH3j3wNwguIDcqpHagJlkb/CFuCU/urtKiUxHLDqvGBx6
Fke4PvME5tQ8bNMTQx2D6u5SqBcMF5cdIoloaEJxxaR+NdXXVNxhEcvDTzfNkAUs
CKC9wKc/CRycFFbEH4NKOc85/P42lZ0stpWx52TAvZYdks0fCqTLI4Lg4tRXAWIO
vZmtq5A0TsBQdJcP0R7Mxdz1sl0n6jYlZOxQi7QZKHRHA/ZTfoTAsFoZW4BZDwa3
g7iaFS9YPpto9og6HfKoIxjUWV3E0PD7WrrJMsyAST/mhTE6JbkL+6CpdF2/kkEq
ShzMojOuSxNW/2U1fDbJndTLahwvPWB3vjtc40o+xA6SFZcsB9MPIUofPJwD65Kb
CA/kjV2plX3CdL3RunA91dDjTbsL1OJHZTNsXEbD28gzoYfdWryrvGnqxxYpSbCz
zNdSl53jJoS/kdU918VCPrvti43BzUGUdVXh7xsqdPDf5MgT213mwMK5hkXb6b8K
zATJ4l/fdy0SgK6bu5EqKLwjNM31Exd8qkunZOhF7Vm6P58nQ1XEkig64SzJI5wK
D2tfiK/IcjRBG0U/XDXerO+igt8xyS03dtk9NT9mBlcu4DjeQrR7/iqziUKsytuj
fqeTbhZOPu4B/KRx8uGXwpFw1RkjStepNOvbY9VAfyLY4m47r7IN9D/Chz+gh7RX
Txv+POgz4Cdfea8Bcqna1JJaHhHSq83Q64xm66QCl2+GihmmySfuEAjU7gNb57el
tYmd02AWH3edj0Qn71kNo+WGSgZqsdjOe5iaOm6ti+YFY7cmwuLQSHImu4rHdrKz
KumNea120duWHQ1L9eKtgucq2xgHKmVnaoZFHlVb+FmAa32I2SMur9AwmC4G8cPA
LpiTtfhgnjiglGzgB42jRJpa3AHqtf2ELpVGUde7vAn659cLcdlG3b3VKD6MZXjD
UVImfQTl1XrNnE64m361s4AvcV0ySDAURQRjF+Ii1FLQZEy+NDEjHCJS8nb60+Kt
OOSR9mep72C5hgqv+RU+EikzfRgkoUZ6AN/7e18R92w7UP7SKw4ECfWJPRLE7fYr
PbKuGZ34OG+x64N+vARPyCBwmKDpSdiP+hhHI82x16YLAqWpm+eFic2LEzYXWwfN
RTjS3XP2FWD0gaWI06mn61WdVknmaa+lfyMVibroZDohbJOCmaGuemn/N7zY78YV
nf2K67DzjQV3cG5Kw2qDww8ceQPAI4Qa6633ouQJqhbsjLezrgAcWM/wH7Rx/gX2
EefBETBhlj89aT0x9mMLnSyPpezmngVS72i7CAmorzQtcgBhFx4W7cZfnitiJZM5
O9VPI5TQeUJNXxRX4jjL1anpbH4rRFgbZHE6kBep5IFKxdfiLzst6sFn9WYoNYol
cjVEJd7lWYvGpo8l3d4wSWoFiPwUlYt4RwCZLaMypzq9YFCuTkA3+T6/Gz+CH1Pe
8Ph2Okpws9vNKwmX+fyis9DsEwyAmvEZWxN3tvqHx4AfmzjmPNw/ddnP6hgwjVjQ
zra0WM0OROvPTM8DKwnxBjJ2HcKI/LBa+fu+ApzBVWdY5BN2FuLPRu6oMElqQfUr
wSDIybyFMoVu2nUI/DAyTNIT7HBmxqniYfW3Ek6gw79v063gjHoTLlPCn9pPD7B7
uziDsWMlvkpsu/Fb3L70/SY4FCs1wje4XLLrqencoiGtBDn9Pr9RjKSmf05rq1Oc
gHs3C8wX9DBgtzKBY1C72uAZtGhauGuwLxSBzbBpJRaYc1kT06BubNMeX1CLcXI1
oP3VyztQNW85DepYY/8YNig6XCRre8jfZwK2bYk8VdZIGibW1IIzscLPHUhiLxe8
Wh9VQUS2X+O/xfYecHVyh3w/B5TqXYGFIxQFZGeTh9h63+GS7b+RMez0QjHzmApO
oDQV3SllCk+tc0l46mkiNCBvdbg2LBNZhanFRcpXYtfOmvKApQSeiTsrUxNW62q8
BO+BKnNjk6jclBH4CanRSXxOfnZl+TQGzAIzbT4fgsgH2Uj1tZGiE/og+Oy5XN98
jBMUZoDl4cj6Ils026apou5CgpUXyJvXToRs7lgT6RDL9QBPg3AtDHe5q8tTFFzd
cIZ/M7WtEdrBJYtJ1Fbc7SJ/ehZeNVkp1r/utQkBCA5hGHZQ5CUVOri809idMfya
e1J9uExIqH/JECnhausTtIUsYYyT+opChTK+bif6CUToofU+IpMrCNDfq0v5lOuO
NfaGv3pbhv0UPV7cM2c6xo8ZYRmscwTWX9zj8F8AXOrytVTphbrIBzmtrLn/oaED
WGPDJYkee+Rbo0T5GLr/haW1k3ayWGg7GHHIW1or/2WH7SZsPkni1TEa8rsP/nvO
Kvtqmixu110ccONd4nTj+g5zvzaaeoSpdGi//cdDvfZTYQiE/FtUGQhZoHHPIkpS
cKeljfCp9Yp9pjlVQExe4UcuR8sGBJCe5YbAhVMMADZ3qR1Y/e7wiBVjI8yYZ/gy
n05rJoUf3CUSTZg3BUUfgHvcjRWK30S/C5Z71sg1NuSPsg3eKd/+vzwR2qhkx3BI
wI5qKuwDJe8KoBd4a5w0ENyKZiTThgl3j5qUdZixWfBqiaoZBFlo22vHKFImlpjg
Dq9R6KdN7X0Pv2QnoGQK8VEUNbtWZgeNQkATof4ysg3Qa4j+PPcb4meUFCdtk7Wd
7CyNBs4OHh7JCx0a/FLCwmsOw+dZMVIZVj4594hhys9e28Ei4y+dRfcjeg2qbwVM
q+nj3wpEbnwW7MAejpYEAYNzYugb4gN6NL7uKsf9wfLWe59wlEPxQFpeCpq1ctAo
NlMGQYzzc0RIIZ+yMbBA6RPP3tkbUuDulqu/M273L1cVZmIt886i60hvKDrkD2kC
bBi+PfHTgV35V2dhqdRaJrPqh446GJ5CzJFesZUQDLiY3aWu+mVWyxzvxX9l8mJx
2oZltK9dvzg7qaQqo2+mS1TGWPimjoVRHsRu9SYFBMgh3R81tS10yPuh3PEGrl1T
7/ViV4+K53E/WYWaqeOmAGNOBLDu4p7/qcloYuKQrVsG3OWyVH1RI3Q4eJMHXD2j
Zrd1X5eLVd7oQuyWXRrMVqZ1G8BhkM4fqxZ+cdYw3nJCcmP/e28rw/otlshQ4dUN
0KwHMgCODyjqG2oqWqqEaJ5lJztv95tw+gkaTEBu4yHpIQZSA1dbcdxQWbB0ZaQi
YZ2FZU50fed9eSlvkLuFDJzZKvCoZMH7UG+Mr9wlpZGR8mrifUIawBLbb/sSxlZR
EXwdWKv5pPgUAsnfi+ONGN5DTEF0Kmlje5EkvywwT/xNQTiCc9VCL/QLtIxbWFDW
0Q4DQd+J2fK2+WkJoThLu8LA8EshSrsydqbqg7B8d874HaZ9gr2rKbjUaUXHVvtn
EnX3FHR4ydMMQba3kXiAYeI2/sPjUg5BWI9HialMTNevO0WrQ7qBxdbuTJBfn2uR
w+ILlDKEgxrq622w+DOKvzmat+FvrzFGTjVP62vX/6f4U00EdNuCBEFvBwCx8aMM
r42R9RusfMVIGJOecwOlrs38c5Ii8vKX2ulHipEidFGF9pqlfHMsjozFIb0O+aSL
lwQg7PQ3buw0QuXIr49RIdnHD/JEqQA9dyCpS4zZcHltK2XI60nmcp7i8mhb3Hsi
132H8leg2SyEJ0KnZpg5xWGnQvTzKHapOyj6aEQ06oy4NARcyAyqJ7WGjVHGkD1s
L57kUtI0Nj7q42M8cXJra4r8ntIrD8DIHtVKFfpoU7ekQboNszWMU92Z0npHO8XT
T+K5KvRvZz1kIxQr5ZNHx3/TgJrSGTCYuo7hITAYJLi9KpHIf8MfXWRJQAFIGKT3
9hu+C7XVPEWozZ26yAE5dj5BXnA9c6kmSiSMT18e346nW+B970qU9moIHYHo0aWd
Xp035ZLqqV/jbHCY4xIMz89LjiNX2UlaV0g2pET51Cc1Q8EbVJR0l+mbLEyj6Kxc
VUD9qcoipgZr+4J+dxZ4aelQtOp7UYj4EdmubQmJ0C8ACEvwvzEZpQzoqzAAX5ZF
Xk4Jz/H8pQjqU8zd6IqPyQb9anzFB0foX2MEB0aE5eGeokuBdslGDYYPM8qfWsGZ
hnWybiqDABE7ar3i8RrhGGAr55z2+v8+OQJVtZvqF/OLduu5tnSqPh89CrlL/6aq
8bGqisDRRaO2iKnlK7PkSW+0BsgGmP9ReqgVrb4m7aQQL3mTLUB/HHlkYz02bFDe
te/yky/XioCz7qxF37Motfl9pVLPFnlsOe9XQYX60DK+4eoGGFwBsanxfBg7PE0r
yQjie4clEIojZFE/wntH53xH8psZQ3U9/vbj+KzXt3DE/0X2ZIhTMXgiHbax/bP/
sez9+TOzJZbpkK/zh1jFa8gMQMAZXDOYVdSO3YUb8V3vj2VI01WKUVvDNvWO7CxM
SYB/8cvX73u1Mj0xZeOXTStB/s3sWssD/ScieF/o5nSqoFRG5ny13DOcpqJBbofe
rVhooezv5J2gLd6tptOt/EfTqxtjMIdgnur5u3PErhxUs/8pUCeFVEFTdgIVkm7+
3rAfbpNdoN0ZjVkkmilvtu6vnPvk09RUVDup6fP8YkCDZsB+TySyfo2x0LU/kBpb
KZCyLf2Eo+xzwQYNc/spVRQ6ckQoOLbpGVpNiF/UzhesysQr54yc4fRcwtj75hHM
f2EimeKdO5VGqIU+VLBGlSa/8L14vAo0qNclZWKxcp8MxUiSX3W0csegsHRNyHxp
GhaK7GND1r150pLYTieaZQuaqLrxfS/LNW63Bh5ELAM5wCPNi56meLlON7DPQWhZ
43LLwWJ5RXbDOZeqz2VeagZZMIa1d9IXl6Q3i5aKSRDe1V8UziIrRSpeRhOZivmp
nDiBXteUIQqO6YfAmGe6avgK+ZixGgu7vQ6UTwhYJfoZZb3L/VzdDc76z1Jow6As
KHrT6dXoUj4owUXdT6pSzKl79zbD9yNjMFxrf9KgYo46Vnb9TQ4F4aNbgPhlq+Zk
IdBLy4ewGzsJMPhHc14wpYOiFcQyucBMl/ZWdFo+81HvDSA26C6qRHI7GanJ+Nad
AqlF0mMXtgivAIBk9/+d+bURbQkxIJQEGSEHydq8r97mP9RPE9/QeZRm3egdspHd
AXEiFgsdQLuVv/Djb8DaBphNIP/Sqb/4PA8myM3b0acQMe91MajAmm+oVXlgGai1
bcyvYqk3NW9TSmM3Mg4oj/BVYJn1V8NYBe56tilgfFFJc0YfHkX00iE/41vejiXU
psHcFW3Tj+HNHaPAYudWYowVgqV/RXjwzpRmC7S6MyLl3FU/yG+epkyFsTVE0lOh
AltTr+vIGYYwoMUSiaPaCvYCsvcVWBWnlHvwgSe+K0qtPXQ+ao7wCdX/F4PVjfAq
QP+gP0zXuMa0Re7WWHn9LYdyMuZFkuROJkEhty8JnHf44rMmmRmtHoyp2tNArZi5
53BL0mITYHSHPELys9zPzY8Ia/ovlcJdGN6sqIA2MTa4XAdUdhAaS9i6mEDPMT2S
url9j7nJ4bm3BSdZ2ukClkwLamA7h9x6oEwMsgytqfBTLOwMr+jLJFdzRCQJOK8S
KbUlGN7Hs4Adcn8hXFsgwKtVDaqXvNqiRNkAFeSCYe1VDf3QQ38vf2pjlF2b4hcF
3U9sjKnBZxqMje/l+Cck7WFsxFyVK6O1i2A1oGlz8nUHjdZH/KM9IWWHOPS6qeRc
I4Rt0wL4CknYD5HR3/BuZ65lnYlqIROK6uEi8y3o/FBKkmaVkTYYx41Izeks+Jko
g3H2tt1QYVx9gJ1oEaF6qcEcKvMKvX9g3NheFw4crbMFvje//u0TZ84qk8+tVnr2
M6diV27HY2Qacu9gys4aYUikRRamo0r+p0yvilXWmAvUrx2m7HlNfTjMKtwT6fi1
1z2Zun2mFzQ0KwWfdkk6iOIcKARIFCjeV0TReNx1nHaNKtnHeHZfOYfA1vg+FwSW
WK+W96OyAVnnyTnFI4ajLn9ZrjFp+JXHHzZo8jlmFbNcCSmsI57OZjRu0pCwscr7
UVQ3FXVjJTEM4yQ/RR2KSnNxqxyqIunuP9a1F49N2ph75FzOXIx6mWd1o17aDzfC
OEXA8uVzLdB4Z7EuufB7GF1dZLN55Yan0oV8a7WTdhPlxvHDrLI/DtXB6onrDL47
1rVEP0zkGee3TLVBOxe7D5+Rx5Z4zo9A8vF1rOLBmkpJbM/+wUUxVWgDGVKIzeEY
A/Aj7mGlI85e34xTiVGjP197PYrgtqOtRmCbR95oosTY8Oz/aM4wf7MWagP3oR7F
xE/lLZY6fqsGFmWTk+sNAy4AQaK7LpxkaFyyc272GP6EUePaN5hYrCklJWgxwEdO
CY5xI5ttAg6+Ui9v0EApRpXrWcAfVH42vDkTq3aKiBN54gducu2bT3mDV6zQl4+Y
33ltGQmK48tuqlcn8ck5W0MTn5h1bQqfmVcscVa1kv888dZLSKZ0IZS1I+efe9kq
xM4eH50Cbbe/rt2bPl9UQRupRrZbmhk+2izag+Zyffk7fWe7pIeCSQtM7YRZN4VK
AMqBBowOpVROkco+Gkjmg+OnOQFJ4bSuzbLNHKLwSZtQuUoaD2ewowXa13HK+bPc
Lfh/q4NxAiJkwOpBltSR2l42ze1rxMUKizyHsnxBtipj143n0YiW6CYENIhDTNwn
WSnlKx+E5ml1xTJHOk9ABSiFFQ+9SwVRFC0PSNMscpYCoyO4WVRslQWGPjFYWH+4
3HHqOyOZEacSnYTKJc4jOhkKPErQSMeDuq2l6IK1dqHgSp7ETfIy1spVaxQvIENU
+v54dPeQXKB/W4jc8btI0Ltx+hxMCbepooc0KfsGkSIUPrd0wmPmNkUXI1TLeZcX
QbjfXNCIPD575l2gehlE/kUoWUAwuCY+M/VFdsKTpDfIYegLAPOAqGfwhdANmAw0
JiN9OiJ5HjW5wN3UMw6KJfkHR68SfdTF0e8b5FyZpHeT4eiZLcfoILUPMUJseEN2
evgi9644w4HtJL6lnuYBzX5iyzzCsu4C/bqsZ7y8PiDQhR9EjAhsgUMbRtTAwxRz
qxCTAWfVJR1dwW9Aq2dagUr993QAcVAeKVqMvvAWmQo/w00uGTdzbEYVOo4J9IRn
t5U5xqKZkzGTNg9fh3fc6ertz9zW5eXniYFVVx0pios2rCVWS7Xf4LjyDi7b5zVo
3sxWn2Go2CjPj1dUg8R00fjLKXq5l+mam+Wh84qJodOxs5S+ATlmA9OHUFl3pYsU
35siQm6pF77rvPgCsWtSBqQtzNHjEC98P2CrKg27571G821hNaGYiLanpwhhuaft
QaZOLPF+GAioP+gQXW2vXzzZIU9VJHf+/P6Rwl2CKI5foO/oaemLHgjz4GCgxbVC
4n1/Zvm2LgntaCAYoX/f6yuicgFzctp5cy7MXRxYR313pjcyGBF/+WhMWdb/m/Nl
MHw5T5+da4HRogd87UgkxnBFFyCn7d/ZISVUZIuus50iM6SIrnPNUIM37IVwgkOM
MJQy/d5SGUPfjjTSqUXa+3rDcSmPc8kD2duk7AZ7Opn/djJGWyK0j5DJp0I1GdjE
b0CwFdMAwzQX/xjhSelUXT3rTQS4u9elZq1JAofhER5UixMngMIE/rFrWX9ggyP6
/xXojNdJDjxyzA6ZWwt0aFCtSHiJ/kE+6eB2MQUewvRP9u0eLQoKmeUm/LKQ6Ul2
ZzDwglJNNJfrZbZKKn6bIYfNrJie0t7xut/9sKGTG8dgn1gNH/oNGp5Wff39/xZP
lQCcR8ve/1asPr1FIcQTOVvrTuaFTxj3itPxk7W42kZAPo7+kdiy2F/5/XmAi2bp
DDcGnXoImHMNN7SjzeIEh4Ruqmmz4ipWJvwYoKl0iA1JwGB3TUTSdW5DI9M049hT
1VT4CcWeEK6XDaH0mPNh64zdaYeCxZUMkHox2MLNdacCaDC160x0w2hGC59iJeYi
D56uweJagOtT/e2faavO8H6LMh4AJGCRwSk4CIQ+0GK8j8XfcjmTPAgxDla6DVuj
WthneychIOFcrP4/sNugTCGk018kvmFTVZYmHNBEMCeynIEayJsa1AqMF914klM7
EzWSLWKgCSAs+NYcBHgzzgZlDLDoywYP6S21+9gwnr58lypdm4hIPdZSQlA4+AGK
Ei2MBBLfweGpgRZTOsT8UoQtLE1BFNr8Mt4jLYrjbS9Z1ReQ4uTKpz/Xt1BXpfec
OL2Cbj6pnS9TVKoLJp5z651yKZqSUtqGQhqeTr0pr3nlUIRvo9ldzDIjejDPRTi5
8l7seQ6TfH86ZcRIL9HUTHkKci8evlHJrXGyy1nAn+aL+sC0UznyDs9mwEG6HKSO
059OGOIARUBeqr4jvJK1A5WL1uAMGn6UJpoDoO/+1gHpKA4EqMC69uhIDG7GoAgm
MzD0/iooMK8AMoT9A0U1e0xsS5XX4FFWOHWzZViyvlV2/Zs5VQusynwcUncA74B9
TJC7wDo8VBeDRwMKmPX4Wqe31BdawGfcj36+hSSDMhVeS9UCLjb4yTDyHR8d2Q4E
yrt2IeWoTDthwlkoUI2oRa/fp8bmEAUxsxv11hx6+VUNbJB4m26Pka87n/qvAWfS
c7XreOFaBrRlbhul6a3MOIWqvKT4Bi4wBT9YrrICj6wTbQzMEKFeeEETdp617t/d
HuxKdDhp8XQWglAmJr6F4H9e8igbYMIlYvLHMojV/BL4hyhcrhUg4FBeVtmPVx8D
4R2abbI0BpwzO3mwPAKVjYFfn2SPELv3/BkGkdHkWjw+xqwtgr5OX2tk4jxpPbGQ
M2oXvDHwSkEckTf6ydE76+Ih+/Y4xSgfF34AYVwCm34XRafkPpO2mBbiZruATX2r
vokZc5ZQB3ByfNOReCeaB41xXESKAZm/BEweB53EOLMEZUJFZIlAHD964wUGKJ2K
Ig/RQ+X7aiE0PZZzmqbk2EmswPhOnj2c9wcFmqft44tFcSPO9ffkjdaSNz+MhEAI
MfQDxvX4ziFcNXDAaKL0pOQiE4Wijr6WE3mATCq2bvPSpGaNv9P6XCKJ+FuNowSI
N6krCeV4lfgZzSNRGqCPOnQlqYFdHxcgUq8jq3ntBX39cTm2IPXMTUXKej82C+6A
2hVRjJTKv8gyj3kx8JkBN33ndcBKWmJcUNu6ntk9nyEQw2w2vuGkbxYn5EOeK5SW
0naxLFwsKkhoLjOhFv8uD7H1JkE8BCsofsj5av7iFYth0vwpLKNbojtOsKdUrCDy
FeAMLkkXYU6YKijcwHS2TGZ2CWch3kZVkh6lHraW1cJ82PHaKzNuzYp8P9TJlAEF
34TdApCChI59porBBL/HdH+TYU7F9p/CsQ/pGdSsKTXwSC+fP6hSZ0I3lGLDIEdY
tgz1OFG04lNGW/b3Gynn4LVhjgr6dA8o68guNQKi+RCehncQiebt6iH/GkFaAeCM
Rz6bfg/Lv1/loENYqO98caNnmrazsDTis5baHKfOzBhhCVakjTWHrY6HIyqf1dYK
9vY+gaXrny2LJ+hGee+GKPD8FgCJxssXq86Bdf43OhTyrSMFvrnMhGk3Ycar/EfS
ju/x9/dOIbEpyCVwwxuYk5OeHTGxg2HUEZi3JdG2/ctt8nEgrt/a7JmAN5OAvGrB
xS+iZUosrN90/4e2gc5feiWVZXD4TgIW+/MKSsHWuHc2zpXaRpea8HEg88rWm84A
MG8x1DGi26i1cT1Cjo6W/VcHCatttna/SxCvIfWCbJUTRkx01GLeaRjDcKhSg1V4
fneq3Cw00cZEfpH2aHOrEXGqAPEFRpwsAdpG6WkNZVHpQlTcz3Dg6GS6CMaiz2ur
HfIa2zS9Tpt9rdjCHSQ0bogmZqf8TWM6kP2iRiH+B6V1zTtkeRGUC+TGYodldDKh
s2UCmr8cFa/9L9FB2KQ6RSdqJ2zB+KKW03RJZQqV6dDPwLkOCBfmlFS23UosZIG9
GEWkdZU4axVtGDYpK/GyzXiz68+qqCEZwjKz1QmbC4JFrfDIXhgpb3LBilIafI/Q
dkWPfprfMKmoFNhPvsAm7sLGQnZA6G7JmHl5YJF1hFWl0/NmRk/W6es2/Xvbs16/
pMoOm3Gw6G5FQ7/uS5gzsBLnWaDM29/HajHFbhOm2EpMruZlbaqysMNxt2mSF0IM
bBgYb6nE2/erQurPddGbjEtYsUXBOalTklQ475Wb+3Ghf/n+yw8WdXAX6P3eSgoO
W6i7t975Ypb5oo/bJkHXY33lWxpKQYKQqu7P+b/nzs5lhbmIQW0dPLCz5IXf8oXv
AfPK/nsp37GB5BZ6v9B5h03JrtLwSrR3RnHGrLbesAYfHzR/KSKs4jDhQvYEwyGS
w39kzcsLeZ/mAzxg/vNN6Z3fnGLX6PQTqQTbHwgXimnBA64bicNsHeAjIYv7joS+
lTiMaWccZh3rTIuThkgVZahJxbBZa9DMQ0AVVymOW93M2Wl8IxiGbx/70kfeb41x
CmmJUyQiGkH03x3YaNF9FmZv9dSY9nKIG5jI4mmM1tnD7hX3YoWeVvTSmLvqND7V
gmw2F1E5aXvke+6olOd40+XXZ2j5R6FrZhEE2TwohXa/A4igaKWn/+qBo2jB7Egc
gB4gH3wc2XO9XmHpQ1ra1xm/1e6gyFr/Zf881PM3kEYdylEpj6DVxG45LNKq1bDU
GGAWgxh3d9qMRGCU8Z2BuMiEUQ6Qgn9B0aXuKIrWLQlnNKWUE3CRHoVGW3CSRxGz
S8xUTrE0OhkrDLDPaSDA74crxJpGIVXvPZWxAR1WXuw1CtqKRmWQDOepH+BTUvqi
VHOMUXTJ/nuMYUN1cxZr4JLKDyW/IGtLEtx3HSzb6E5wLdGCuVeYo9jdE41sk2RL
QFnzNm8fos7Uw5wHyc5zBdpcLiTfYme6RLS7Zail8vME4UIQPPhz5sGBxfpQRpEo
uOCyqKjCzBvj02WbQ38xnWGVaAL2wscEOewA3ObU1hiFtSL6Oo2g/ImQNnFj1e+s
dQzjf65G/eD6QwFfA3bUZg4MXvLkTtpjBplQgS/2Wp4eS6cGudMMut8g8HrKUqjQ
DIZpUm/yuQOso2A6zaesMGOG8ArLQagpUP/CdJgG8JD1qrAwHNV2ntjskcuVUWEE
PFFUYFnU1rISzmTOoUr8N0Eya1ABw5Vi1VsrPa90EAoP4nPC3TZAFwhAAe+IBOIt
fAUOrvU1sFwobJJZGpoIg6vR+DcvgKL4PaLXtqcrDGRci6w099q4xWrO8s7m5RqH
laV47+T2iBqE4ovIs/aUw40hr3IXVNGR8hdHnXe6jA0E8dDajrSmeFyDVnn+bEMp
JzNRQCHnxoGI2m3NOufky9Wgg4PTRN7DItgZHrjS5bhGt572qsuuOJFisqSbLXcf
EQ9nNY+LLF/PCRK1nX/BT0nGca/A0R6MyZE8goWcPgmA4z8ItlXilxIUcENagN7Z
QixjQED2cFRUjqv9uTKlm5LH81p842MmNi0Ly47R/XbZX2ACr7p+C08FXbXzfvnx
uzNd7UFFbOQGBuJgOFYIv8h3SfpiQMyUx3l7pEpOjhtpB9U1YPr11wwQ1Tl2i3Sl
Pc9hED9Sd27UlzkqHGPdvA7g339mD7DJaWAbhwkfZQOVONzFWU9ZKuj6VdqBKdqG
5BrUQ7xfl6Bw+4UbBgMdoSfQJhBpQcrfZAdFc3cH7CqHqmPtFmswvUxaMFI8hYK3
Tz+25YtCuWaNRdAg/T7km0P0KAb+HC1xtpR/7tauEzT2MHL6n/xFfzC3omCc6DlV
DPbAIJVpQk5vZHQb5/6KIp7Osn4hhVRv3mkcysDS1dDerZCdjbJZXMVZpxXzqdPX
N4zIwZFcyEzD8dI0sTI9eb37cujpiWVMnEIwjFQxpkQHRso6n/sCpIkF5miiE4FY
zJ4cy80Qzt5OmcwzdohX8MhPuQLzAxxKFTNZjACom9kroqxJ+b8c5y6RtiZB/tx+
cIE8it8KR83acmnBb6rvaIPo0Kh43T1Fstq/zq6MCYggqkHvlPK6RoPHby8+AYVs
Ex84HR4GiI1xDkqzLojDlwHrSewI33XMPAzolDJzFac2F1+pWtiALu9YULpg4tws
lreE2WsUnhro9BBgGVzIuCoPypBmGxNQ68aOuSVJhAvQcQOMz9iT2AhoCC6B8oca
3c1xZrl4zumgKpFSsLNK5MUy9YGkbH+XIBlOYcIGDbxpQT2cgEvmXXBu/E+wOcKc
JJo+ZVtvYyP0cuTKQS6OkGCnJBniQQNs2jiDuw34G3VdWY3n0SuHt9fhxi6Mi98g
vPxPyLn3/KhGO/liClmp49XJDIsEuLsB1kcMH6SRIPWh2XeS0c7/st85XhRnuTEu
XiLhHrue9qpo+tkhFFIq0nHOBEofcs4bhtc6J1xOezPEimV+8gK6jJDWnTXeZnZg
GDKQAI/3wEgaU/3gsmkXRhDksux9cOectvGO+SS5onHdEF2hQM/USNgEuKzxaX/R
oykRB/6dSOJ3iL63jnnWR6YwT/ZMI7+pBZKBqWN6p3oWr7Nn29Rg5b3Om0yn2Cwx
UDOfKUIVavNUYrAsGcY0ImsTvuRAglOJcfqD+1EC0vsEtfTBTqsAHQyIsVlMcEz3
q1CvCN8m6/ORfHGqWxo7LTCq37CdPGMtJZr9z1tmXjRRO01tzYN4YG4NmFJkoVaW
dN2TiTuJQ1Xdww3IeC/iq+sfKlxsCv6TM0pCWWXldi1D0rWqVK+2ueiZZjaaWR7p
xvCS5kDOPGEOFXj7AhCzzSkfyjCpJRtC2VJ7x3lcAp67U4vYokF43pD5bMFUGuOx
6R32jOqHMZ21igEJRd/kfCSgOukqMcBRVFX/VWoUq8mXH3vZzZ2XaEss1Qbb4B7o
wJyOST3Y9Fo4vZruG1eEys8L/TEmWuCk/RzEVRCtsoXxfnAa+6djm4XeSTVvd41U
h3Fc4Va8k6+a2JbfMdhyI86xYXVrAahfE7aD5WK1zwypU5PgGpPWWTK0W6GBxmyP
3HcbeNsXoYhgtlP0zmJ874IL65QnSNsuAyuBeUYwV6HEekBeANhoTFaUUa2x1m9S
8Lt1GNfF2AcflW2QqE+REVQvTBqDeDF8lPqkXHzMIFqgBtLG2fyJiwqiZ0ENXFaT
k2QtB+9RJWqN5pyZrqAozi76OiUCk/B8IVtoC1SsmlGDn5b9ROkpBewTwcZAuMtY
XV7oHsXhBvZ6EWJSM+0bFRP22+1zqzO6YqBdMSWmpglYJLJUZem6Y3al8IYlW9S5
486atEKg2iM9rJRgQ5jAt8cPO4P1nTz2Ypb7jcw81poHth8xVmrbkhu7QokhvRpq
EHtJTjQc0crJyM9BmVPZy89VGKPMZ4fpeibvnOK38+7KNL5owSjPAK+d0xsV30iA
6zMnCaRDWhCu31WhfV/+6SUUvRiYslt1M2V7epiRBj041WN2mhDyT+HqQFWkFeSw
h53AgSH7hhyjVIA+3kqrOLS6n8IEGi2WeN1GL9HzeDZTOtjXjmjZKzUT3RslIJDI
Ta3jyhnOFbR1WR1epNMxZk7aiPQXZTKm/LgXEK06EJLC3lCAHwdU2sctByRaxHMT
/ud2rmuRXUb0s7b5Fr7eKOh8oLKos7C9BSSmISPatSnbCB3PMT0S2jWGFAivRozI
eLNFFb/bOYZaHb/9cGSJOfEz707mHhIINekRw3k7vdBiSdS+OgsVjDfDw9Cmnf3Y
CFSjBJyeQx0wEdaPEXM/TLUyioX6wH7b51sNTJt3AQFgYc/R1JUea+d4O73E05tT
DJbn7dhsYx6CF13uTo/7nWFj7/ctmMCZ5ZffB8CtGnwpTe0vzX2Wr55JJPQqSeMJ
WDYyzP+WwhAqssKbTvbPju1BXnoIeFCkCx3ZVPrRkIGV9SOYjM4AxCcqZffQKet5
Zt0A650MglMCdpjPEFR6EFwyCVLZiuqm/DlJf+oi8egdq+eXeYgkO0pxmA7VrVN0
T7yZyq5hxdmKuaghtB3YQmcusgroA5ViuMcrYRQqmOWo69V8aaL6cpO087bmD4yy
uUpvyTVXf4MtwbT4VgKRBZealX7wkPcXKtXdPWjTmqv38e/RxdY6MS8HAQmgy6zm
iO9teNCctwkpIElW3zmABErlRpqrZ/i72r9/WatBrA+vOMjEbwvIa6jmE4qEXlLS
Da1yl8wGOC6yfUa4o0B/GAHuJ9H8JXKfeqPARFCUuOuGfqKatWSFrZ7V/wQADDxp
BztX1mD8IBI7yiF8zy93WXoAl58UxvqdBXgoTmHTWn3WGZSxSyqIVCtRcHU4Km2E
AW81EymDay4DNDZlfehbylDDK1ziVkYwPt9RlKqb6M8MksfwpwySmT6GBOxeHt56
NSfwHsf6KdfJO7/YTvxhZ7jr9l+RUNbXuqsHxehSGpOW+2qnlzZPi5LMnrCpXx5/
rtVldK3G+qGniVZxKoXXFNhXKQNh7HchxZ4CvpO+fxeq5mdGTEuYupnSiksbTlFa
O/djcWvmiGcuL0suAH9i3o6YYwKagvVB4LsQuS6cNS/hexGiMNOmmHMoT7OVZTj7
+TA+GDfs3Nz83/MNIBaKmp3ppsy2r7zmuZqtswXeh3jkJnavThnu6v9e5+hJC/CV
0fLPVUDqftWUJcyDCPORgonsS6K7ansl9OoRPt4mtKdVB6mvKwbFQ6Cy+wAgAlqz
EuNXY2gCzYR5DdMDUIvKLJ+E2QOdNX5wnhkpcJScEU6ZQyT8CcqOSQAsBDidDzog
XbRK2WgXZ71O/SWDMG1lH3DW+f/ELuYPDASyfsaWpXiIDDmoW6m00AriIlbHNmO1
3AGq9E+DUMkIizv73sxQuE+u/K8Gn/IQvlouZto8qd/lK0GqC/kMgBv4iY06crKc
vZ1mBOvJowbcXmOrFRM4Pkqako/L210qewQll6vizVs5VwHDelXf9A6GXgzjFVhG
9ptQ8LXIowEwOSQGYo+hYWd0TWIvwMcVPXv2uqobVWqmDBKWjTZMpo2dWVqK4g/J
RxhURoVTExQqelO1aPgVUfKmMAJynOnixt1qldRDCBOq73AIx8CYUVBY+e54X6iI
vpWAdYLsn54UpkyQijfVKmnGdJ6R0PIDP9+r1Y9mvgDIKfmXt2Ara6eiL3iJQ6Q8
GLAJ/7F8AvbruQFR6u2uBdafVBvJ8QyvDixM2K0IqILF/JO1VKX95seYVeDKLYc3
YwqXS0ERyZgiKDS7bKiTKniHQjn1JU8wLQO6y8UsHmnttZSKDaxDVHpouX0CSgnZ
jPovzOTpSpWQBNm97pPaCV+IabT98j+Yn1uVOR7WN5ZtZ3s2TImMs9yO3uC2nMcY
17MpofsmNP1q52E8cHe23KeN2FQm3d+mgi6Bf2HjlSDlNQG3EvQQCSjuL05voe8H
LlKU+sA0BakHvJ1oVgHXJr96Flbbx26TWkDn6r10uB0gbCCUJwJ6IkfhwNGuNuPP
49FCp5tl2iW+rzwXaOwDJbcYzcEruRRWFlRyBSwVYrMw/YwnigyooXX9wB1NY+B1
WaMgPEf6BgTjChteqdO52ljxxiHnvXz5O3lyhlH5uTiAlfLN7mva0SGPy7Ddm5ND
uJPHEiCGbYbreS01gcHdQXqD81vITRwdH4ec+UNe2yv2t4lwRLDNO6juQRLICSzW
lnljDZebVIE8MypL7wgOg1rPRyrveUKD6JOlH0+aIrEEzbzxeWyAcDOmi2u8pUPE
w+Z5v1ihm6QSApUO1miR1z780Yw0QtQEZOaePphajl9lSmGOrRdjQ24P9cdVpohf
P0oDZX9Iq09z10EUxGsYNYQfLnFFZcC7S2aCY9B0D47zWaeRBioH96zPRTFWoFoK
y9ldocVHDdNeKzlbEQq1eLuxig5/kwJ9kViej78Y8RGHPRIWtTfqqWwzXCkFKok7
6+C20Q6oaiGdy3zMCQff/pVtC//zT+GqxLwOJDt28DA1SB0IgIKQ2qOj0rL5neoU
rZ6rFlBL5pY2KDl7vcnqEhKkkyBLdMZMcJhQMU316YlMnm9POmtFltEjsymFcHD7
nTbtkYkkJKPyTIs6gzS1QBfRt/Fb8aMAMbvZ4sYhvjl9gGKnBb20fnwY9z32nFe6
qiaIQyYGzoy4/AzRdKLtNMsN35S/2y2TI4YovQtGizQypkNKJ8Fsl8GhNtgUsmjj
YQ4hdWua523nrtS6jfJV1ncEFDkXsIQqwFVo2ghMYCTXKhtMstRgnwTPVWcngsn5
q078j3Cww3mkGpeDI7EXChf+RZWGFy3LoPOOUewWWtnexGT/Lu7PrJ1rBnitUHQt
9EUlaQTmPz+88sKqO+k0yZ0U/MFd6Eoe9M8WgkFCKLvVGMsf+vVki8uAkY42IUUr
Z/28lMZmOpEiGOP+16diWF8okXBbIn1d1iDn6kAw0XJqdt6t187xW5F88lmIJUVc
TtD8BgsZoIQPwQgRP9FHgXYuDBInsSjx9Fe6MPj6fwFfE1LqZ9PmGBLDyQ1CPWsL
nqMxo7VcsluJBcTyJUL5ykm9MHtqmzSEulQNNpMOZDkuCdJBlG0UJe5FcErAMQcr
G9kIgP50lE1VXa5HA/+nWN1kQfmnmZw2xHFIexggIrUX5ZJC2lw3zGx0DLMQpW3R
p4qydps7wt5Dl7Px3x/rT9sDYU6qIC0SCgKUKoN1QdYtIinzPv3RT7dKlnBuSff9
yAHOw50xF0tuUtRR4WBnOg9siDyHIPLu1aiamZi5RxIfMakxcBSfv3D5Th3Ikh7a
UlqE9/XdTpJeX6TSSJ0ztcZJcNg3mjXbmTCa0sKaLLJkaPosUQPVILV9BZIwlZcg
iEDjSoHrO7linY7OUWu5hzj41cGztteQDbNrzRtBbB/KI7Bx7TnJsV/N0DKIWZga
X3aftkHbG/vbkSkH1pUgPxRur/QAG4r9BhyXEaji1LgxrfFImWYRk4PNyCD3KN4b
CkDJ36uamHth6Aenr9+vqbCIYjUefYTL7aM94vCbP+qGjxPqEQ0e0ej53r8LUy9w
m4LdAf8Ph4WEmYGiXOLQGWzUVkkenzGxOjPHbbBB86yLFBX3NwJo9KpfA8GLFNEI
Od6i7EOohmqSuRUicPinIGKASAkufj8vjyTYJce/ZDopvPk4xdIt/KRrkOHf3IRy
gnF2isBM8otGng4FPlqMpOqq52coJSZWiZ5sjd43jEGoSExUVM4pVweTP27vPXMg
m/F57swOyXhB0HsvHJgKqIhgJ9ONr8MmMujM9FXDWPtEnS5qaC/bMxZ3XMjua1pZ
YR38ACTtl0NIeGBxRSGGl8aN9ON73HVzKvMSVX5FHlWD0LgP1xmsbZDzTdrJex8P
0IVx+kPmaG+Y6s9ioHi+R/Pg+8lzE8GwJqBesrbEu8jfSyDzlaENRCnXAQXmn2kY
m4txWkJIAiZFOnhsOjuG6td/zpIxKW3D2cS5tTuVd0rQKrwGQ/qSPb7ImgNVceDH
zhncJb04vheYnkLrP/8UXUbshnrw70QJjWYzhrP0a60VlyZ1ANA9LCikQsyBW1Ia
2LxbrkdrKNvV2PzXCH66VnPy/Caf0KiFir/Roc9M5WsvHIZa6Tkg9XoQCIy1HVjX
VLyl5QDXmHTviUn6tSgNRoQTMdniSR+aR5YZLZy30QaNbFuVOcBzFVxe0rUG91lD
WAg1LZr3qg5d6rE3iuaTtwkg/NuZzvI2TilS3mGhv4fAxRCf3823Nh0A76qACDRF
zBGsDILH7nEsdj2IndZB/GfS+nqYy1EEIvvNzPyejRRAQLJS4St1luZB6fScbuIE
/m7jENt0g6+Tsbx0n3LoADn9XlXGe5ntpt8WKNImDG3eb7brJlE9nzlQd6TbNhNm
ilEEIQni3ZNuz76I679yPadV6+LeSv+CRZy/vWJX0W5QJOQdPMe6a+z976tCRQgW
RiCladFNoTUqkUmDDfq/M16n8DACS+71s7WB0dfIbz8QUsrYBNH1/YccRnYe5KTZ
Y85FBe12ZtxNUUV6UR2udoIj12UMZ8ndRnjDtxODflxJqWLLyGmaDqk3ePptypTm
QG6gK/DvmDnqciuj+v7RCK5pc4E+ky0t3dafuS5MtyMcFobH9JoZeaqD8HB1fj0z
NiXuYZFduoL59XfKOxmLpZOJndFhiNnbdtP2tytEJT+jFJVJJ789uDcWbidun/Qf
2RLOtEBhx4q2E4oQsUQCUngGjkdcJVqx848SHOzDdTEdi7umslpnyeEhR8qJupjg
XEfnG8EKzeu2N2lImuMQ9QH9Ok39+xFvKUBeRM7KRq4uFp0Xgbw3Z8ip2Tk4uRBs
rxCoQrlMs8MHUfnPTCkgMlZWjRHW1kvdcAkzmiUYKbUmhuI16VKqDKs9BsMRNwSK
0R7v5vtITaA+qGwbi8rlD1+GG9FPDaAdOq2nZ1ErmJK3256PBiO9pzWcs9FdfIgG
h5cTOOOAc56FkOTCItUb9itLcw+EmRo5VtsAoSmBOHabWT/2LdVoX8GAHmnXwJot
olOu9xq7/WYDEVtSZJvMEq3veHOOrCiBXAQz6MizKsBgrwN8j3EZzFEoT250VEnN
jQUEGXY91MtDPPnnI5xSeBM7y357U+v4Q3NJxsX1hWvE1T3vvL+tOz03i8s2VBvm
XZQSfGMhWxLYPQiuLW6tVeHAtmD5BxddlB0ZHgibdYUak/SainOzGYZ3b0og3dFJ
g9Kcrg8Aq9lyMPRNVuhhHZhnnzCyk/cgFK+GT8I3C52vweoW8aYq4ilfpTP7RtWr
7PxnkRFmq5fTo5y4Y4mNeaOq2DjBWPc0m14Mit+fOBKUuwWp0ixZkNbu8ItMqq48
yVbsbFQUPE+42EIHBUWD9skcr+yxUdWCctJBEmezuOadcMPowSrI8+1eFLmSEKzN
IHX9rNC3DC/jXLItjimOtjjt2Ex7PSlRKADJvhd5Y4b2FEhCjvnIVQJ1JfcSd9ov
eeweJW+dzol5zaHgT8aMJs3sos+oPh8U/7xopHBB1S4GUg1q40jrgvNvcqaJi0nk
DXKOdJAyBBrrdxxB2wNmhyQasL/tEouGOoYzw2U48kbMqzkHW4C7qZts2r8vsda6
usbXseiBPrEdI/P/gQx/hJ13U0H6doFud7xGQLWTUVjG37yCVLxtYX8mkZ7+0zXI
fVEi5jY8bMp2KABvrc/hnwr7VRrFXgxiSoK9J6pIAVxlROnwTxQabFGIWZKU+g8P
5xaKUJ61nIlcXZSiuMh2l7HTpqJiohyAXEtkRxg7h4H20yCqeYrJs/R4QJtLssFw
EjrxAoT79BZDsVb7PbvDO3Th5YXZNw2nqF2lrQ/XY913OzNsmKu9oUBR23d6lpIp
s+C+e2LOQbL+0C6XaDx7z2pKEhrBC88rlx6kIhbeejFIERP/LnyfJZ4fY5KDbnON
NPhQnzJj9iVK7ZgyaljKjmitC83oAHrgfKQ3adjFF0Ye1kzVbKV8DGMcneSKwZ4H
zJMzgFTdKzR4Ddmq0szwVBS5ysBaYQpnyFSTAO4i6hiGh3RNGhog0mVUZBlKGn7I
WyAOjJZ/h2BqI530obGt0hjRlerNpXWJlwBz5UggD1AN7P4yD+QeX5Z6Lr6kvmrI
8Sgqyl7LYK6EzW4hJG5iWaGXMIMPlWMLEe/2YeN1fw5PaqEqIowGPjpQJ3AJF5q5
yJW3OGqzLyTNS6ZsAB2GdGmArrcRTKIhv6l7lldG4qnGUIUzmPCyZBSPGuqOsfkf
leoMITUGuOwtioj2l4ixTzpDZqZ+X7RsEyCh0nJdH4+i4uWtgFKXsPjieECRRz0g
ZHu28LViy9eRRWWSfsfribdK5BTwM+rWrRM1f1gMpZg/HTTZYlSsJtwIZuINUBIB
DfUNsgJtTbqmN6BgFcTgiXFKv26bt3AF9irdupUb+wXf1ZlcqOYMToTnW7fjXZ3a
TkShQzSTYiYhHInl/oh2ijLLzoHQf3kWRfc6tDXHeLBJ5CJothXf0BS7BSgBqq3W
2Msc1W6xjHENqk1ZkOW8g1JU2GC8Wmm5455fVD2u1ahIRK32yHPmE8slVFB2MFim
D/QkmR8gI4/9AW3m0ciZtu5zP7RJNT3nAPi3/VaKQhRZjhy61XXCqV+fzHKI16bM
Ih1EPX10/eYKnyA2re72KdCVMiBKnz0NzzRn7Yy35IYu/E8fHlmagYF1jx2nloH/
L4EPGtxFqE/A0GEKbyMyyvVTZFcg145oTKBtZn/X/ScPVV0zc1pb6vDaiMN1j4n8
8LhYZD5FTZaUTPWYSTNLUlDe0Wj3RdPOXScbaT2cSN6Gi404/LfYcg8OcJ1AIVAP
jtwU7oKtv6epSOoBP3Y2QBxOeaqsOBYMpYr5Mohwly6gp8+xtNADtaevLT3gay4f
awczF+HVykSsRPSOTwdHjNnXQT9kzqXhFuLqI66MXFqyit0KcpRwTSvAKogvWaOr
cxeotyA+L/guMYZzKoby7Lk9xeezHkcYCCWK1r/TR7lO5TjFVRjlOVE733nOmvzh
i7B4TOmnxyrQ+RrxJgwDaY8o7yeQk2d9pGqTxZT7U37cRoANWL9rU1/YVPVCpZyL
1esk58JLcl2V9gpBCNUZVhu9c3WFB8JWs3IWg5PGMR1pKhLOBKQBTNSbQEnmgukR
yf1/B0nlJPTEZsIo8rkayktKQTuvLMkAfB1TzWGdisONEEpnvf9Gdmf6vHTpS+kv
0LIiq2mgKwXdaHvBkEnd8KRu6AMw57XwI5ou8OIAHAOU95qSVm4UVg1Sgl+ohz0t
xotNwo1QFapu37wHEM4oAuGAoLOFDr6nUCwmZ3rT63emnJ4koyvIJTnHfAdXb3xZ
ZAd6fCl6BCAKMYTV4vd/UV7Maqb+He9ME5WHuJ3Ezyq7f2wxPwKpVU1rsbA4qoTs
3zBJRXXcBvjpLn2mvnF/IFfQdp6XNyURR+dT+JyweRzrSvhy+sFg9iRcQk1unMe7
SXUMfoZlicNcRuBAMqOt3aZfPIgG7kwfoRsXtggF+LOYF6hA4nOmzl3G6ot2BpQt
UbpShWCBgvS7nV9fMwyW8BnRz8eLW7Wvagu9X8Tghb7YbrOT2d/gZ/FLDH1IaDT0
z+sUiPuJFRx0M0recgisN9B1SRc/6iTnT2NJATl73FQVb4AYV9OHk2WkC2+8OjSz
dd4jus5DvNFe0VKb8TY0WPrvsTEa+t91dzH6fhQtAwlcnYPc5s2uFnG5C5i1E0WM
8OvFDXU4B3fm9I6swVXZwNc7nshqGcifh9uM3IryT6f55VaXIotftdVOUr20yQKI
EmCgw9Vk+EafFB8y/sHDXqbk+poeNg3XdoN/wmVT3MCQ8SoUxZiIYhn2PfrzkQgK
U90uNTekbFT5Whx9goHlxjNYq0mEN/88L/PJUz7XItD1+s/YhgtWYXRu6S2GuHGN
ND6QDJv38mTMvcVR91ODSJo72V+aeKLqfngGz1HFq3RGS+UjQ9N1vAziEBOunoPo
fWvwR0V8O8v1VHXTsnoY62szIxmYH75cXy+2LXmQ3vXmPZY7vpvj1cl5xU5UGlVh
bOzcWL3kIddIukvT8yx0CLIajNeClon0UWzeaYxfWqjI7YujrKUjwwod4pHzanw9
QjZhHdzQ1lZYbpgXJMQ0+N/G3wbsc5MvzZPkIj1QgICxBMRrfLpFYNpkwSWgZyH4
9snYwiwtzsUIIBe6HreCj/8YUbu6Cc0aZhRGREQOarTLlsT0Avo34q3Q16pBTr6f
lFta8uXydGls6Kn3MRemG5opziLbAow5fSaGsXZwEi9l/oLMEZDjDshY7mZk8dIU
OXqJ1B/tPkLIfGVTtOYuB/Y2xdr6vjSDtBvfboO8EyzQntybeiMlJx8IhVdOZdeK
gDxaZ8whGy98NPrif5gH27Tno+DwQqlbpsEolf2xC1eOgo/8ghonRuvy0vwE6ppq
F90fpWX8y5zDIwZcJK02BcoXU8s9lVYi1VsZPRjmBYQV0JdOpzZwx8FCCyBbMngo
gO7w0s48UX3ywUdanRxXEA5Jnucwc914FlZxRTE71G4qKj1dzNIrgm8Hl0Mt+50L
dBM1F2I7b5nEqP/UEKq1KdGQvsiuHQ6kdA4L/lP/vIVM/4NV7WX3dAn98aPiZKB4
pWqfuwHFUN7VMRnFghtQNEO9XcvkP2ynMM+CkXZ223H11IzanSSi7CEHvxKoJMPp
q73pu9u3AHoFoVQI1BlDeNAFXEsXxTi3TMmG+AtRXhunEqTuV4OMLlEmaMXNKf+M
kCyNbRvYSd+Lyb25JQ9ncxUH8QTJpzcG42jBUAagJFWxEG7K0xHiAokQ5HdKZaRa
aBDkwNsOzhK6DYsA0CjygdIao5UiuF4FnXAO1qxU0Vp3FEcUnchtnn8WtCVOYF07
DrXZI0Qq2kRhry+1DO63/GSyl1yzG70djf+AO5Z+YLVzQRFvkru+FCIFDyvMrGYU
lbMkTbATtpWTyUFhZ9im2cBzC/Pnvk4p7p7djmz2PtW9r9xUQ/xjNBM6Fbcvca9t
EuXzU8EBM/5ZbC7EargPF20oe9P4A4uuvgB+qfaJxgAAR9S/6ryuVB2HbyyLG+In
OfE1h3zDYSjo3uy1avGi6aOvG54kD8g7LNn1t0qgXIgsuL+blK8jQhoGY1qK9YLC
BYA8lL0JtikM6LCya2kZFljjR+cYxbwBDUWK6VrWOCC3RpAVyIC0PnVmr/4gHTLi
qIZb4Sp2p62idQMOEh37dJLQSavNqrqy2q1m6ht5T7Cm0NKUC1+khk2HTigJrmta
fwZDnzXbczajE9kYJnRi1QcL8n+iNb8hZF69YIg/y7MJT/2ksyCiu2bn3tWO7+3J
HYrUWITJIaT+XjxmXvEuOhUCPtiXRTr17iSqqSihbFpDeO0XW0tRqOdW4lFopsTv
PCDMTJybFqifgpfGHU2f9iJuPLCO9x34D9N9qHLFgeDcN3f5jIHpk4Fci9oFhMfi
xgGl6UX+xwpo9RjUugeCi9YzsDl5OK8kkKfn69vD3hKafhCkedh0RDz8MtLRL65r
zwbQXiQL04BbAz238pQhn9UOfrhWgMnmllkWcmnaClLLfPrIghvvuG+XfxRTOn3A
T+tHVhWNJvUOrCwTP9/ROSJWfwThCeEIw6Vq+GynR+mZRtacswHkDetBTlQzg5rI
vu30J2O3nJxUov4F1VhSVGT5y68ZmWJISOP/4ercKJ6P1VzPjutkVEK77Tlyk85F
85Ujh6B8vFKmh7t9G4YdLI5pt+NU6xDXoEXaMTT7YiIIY/4kPtayhVy0/PWf0i6q
vNWJUGZdW44E1MFkegzK82EWcjcTvauDKHwB75oY4mAJH3O1fr7Cijc8BU+aM5S1
lRL9+UHwvEm6q+P2Q8LclmIwtFxFe+V1zrqFY5uhY9ShSkBJaGXY9GXTttG09g8i
mgwGgl7OoOMNpR3LJ/sTgeUGA92XuaCnTBTflsSXzOC3GgOWA4InuGGK0I1XNCZo
Hfe3RI8BUxVGyX2KxPwXLOiKOGyHDUvLsOc/Gahlmlv7wLWPKvC1tTIi8ebrGSe7
5WatOmW3Tr3devJj7gmJT5SetLfyxOoTbf1/Ik3EjFNgN/N1hSgnBy6lXhOIaAtw
uAckD27aFcMRpSGCOa6BQSQ25M8t5ORt4i8N5HGOJJ2b+imuq4PItbXkyUXGCgal
xb32R/g3CazvRPHqwE52t1s3W3p1Kqc0+bWh/lXUVkqDMvYNQT5kKQDQfzBxkmsM
LfVbVxg/16AJ66Tp1dQQMOLWIRGiYsKjAl7QQtjq/wMGyd4YqBKJG8Prn4RAG4k8
33xv6B5wkWt/oGcU9llN8Ftmiz/deCYCy0bJkvbCxZ2PoZB+oow0Vl+JXHM4j4gb
4xZKAEUIxNg/HFw41kdTc+Vmg/lYTnQSoAr7/MYziGz1AxHuMeeoH3fk5xrkePYz
WlHNuvC0d/PwrPBkpTuyk2lxQFF8EMjst1PnGtSy8zosSlkzMAFTuEoxPosJNkk+
OSasKt8ULAVhGv7AIS1+Jgocp2A7T1HZG6w+d2KMblA3n1dCI3zFw4m2w3SfhHgC
Q17Nhd9RdBkh22jgIE5S108b98/8vRJz1D6dJTmFq6rlC7p+E0b/++29XMH+pVqI
jm5bxxoYk3uhhHulS2UrSZejqwDmDuhDidSpOoy94u/ncoMPelvk2ExA86dcsWW7
pQWU+nHECwFk8w0LgKd6tHFgg7CK0QrNLsz+MS0vvpH1X3gvcsCdaDzj1y8yqjy6
i0lKrt4v4fHJ6tqt8jCde6CPj06LEPXYgQWnw+Kl6gJvklJ7b0eVKiHOKM7qHPmn
KzR2nOxK/c42par1uwl0wtkUhvsF7Ymz+UEwyKcmx+lCU9GpUNNaQa4SAETKjpR1
RiU2Y1s+fBxv/sSg5GDCjuqrQUlPABELg3x7jM9xtG+ncI2E2zaNmwQ573ocMj0G
WEIP2hxJykKYYGDETSeY4SOSe2ADXJaOw8E2XYmNJCb+n0lYIcvRMidzXdoTK1oM
KVz872Nda0lFHdYZYPrnRbw3U6isbgmV5aPnVQA4lzS6Ves7GUEZXhCuMeyp1y3O
lMar9ir3KPvOPKKZz8ZUlOqt+IGAAZFJnshBmpiY8aZ08pwj/hA2Lp9Wnk3QhRoi
fBw63n2GIBnbK5hwd4onld+/QhJHHB2MMJBKshbRrMVnX4FHC58l3MWrTmCJvAkr
zyjUQ9IRmVi0f3Msv/vVCujLz0lpGEA5HZ09U9/qJ0tO+fVR3LXr/X9AO8eTiulF
r4NysarVdhcyxUmYrYE3TiitGyk1UaTshrKPPCnFT63KTj40eIUkI6sF+vxcPzJD
QUKKx3BgyoReZw/cppXNSW5084salaVYuKJMW9i3h7sk+hdfhak7zWFsxR0y+wT/
C+6SCQOB+HCCLncPHkfME7Mz6Q8GmBH4KJT+EytIIP5M2CdbWNR1DB/lc0iHrZOt
ifmC32Vlaeq3kgbti3YU6hIHJzhp0722QbFiDTDByZxWqOX4twNq+PhO8PW9lVjS
B+R3Pz2V3ubTjG5/KXI046N889dAKm/OY/KpA18DGmhHJBu9NI292E7fpg60T56l
X3tlEjH6K+IVc+F0YvGmtaVqF4S5znuuUIF1NNvKjaxS+WkYSDMMOJ7bck2jRjXl
Mwx8b/M8oYaCYbCz/IpFJFpTrY7O74ySg+7Agj3cdhli5fkW54dnLKMgMA8r06/B
BPZFOCeHijwUb26gfSbqAZcyRbudRzZJFj0Peu2JcH7RKAXqEwMFEqFLswxZ2yLy
T4CNt+6QV2XemiSCMdJDlQk7+ES3PuzvgfKqIFgVB+5Wm9+CPDZhLPU1YYvibvCB
G02TUGbJhXPS0BP9pW+u+Se7AsgHD8QPsLlJWtH2R4UVWLawHeib1+yMiuoWsM3j
dUiXZHE5kRVQ3354lj8txB0gcKIoC3A0w4UlDixEwQOnjehQ0gTg735daUt+HZee
LMWe1/fmuDnhqUJaIElRlkOwjcWwV7recvxFIZx3lF+OFJmwJ6sw396IrdXw7twh
BbSSxyJ2x4IrAH5/Yc1CQuJBhYO1aaLEUzYA4BllB/2S9bVgRjbk+/yHy7eD6yt6
UFZYifHbBhu9wWPyy0GuODaZ+6KEsjsdInr8XY4QPFpusjOCuomGbgI3r6BSq/A2
IJchD+FUai2h9MmPTvsGFQW0hI/fNs3KuntpaiPsT3kHkYLQe1+P9xDpamvfGiDW
dAncALgcChvJFBJPV18GWJUF9UbMs0NRL/+etoCvYxj/BfKA4K74BPzrAgVA/OKb
qm7mTrth08Jp+qbYZBVXr0b41VDKj2Di6omCWJq9Cg6lM0ExZeKfOTsALo+mMwrp
3YqOig7w32bM1MKaRcaOAjrbUAhk1O0lyrrQA7/6xHnFFnWrEJiubaAa6LQPUo6I
oGTZ3WhAfhOwbPYNMEKdNIFdPKeIWaTXFskvVokLqynRRzCO6lP78aRUwKLKmi9b
V/H1MYnyQdXtRaxktMNj1C3D8/qE+QXNIroiU63F8M9ms8emcCRSOIP62YEtfA8b
xnbP7F95ExGotVSlxvUY55ZlbF52C1VAo1qZ7d6m15PkbCC979CsaZ0k3LyUpA1H
zrtWDMEWv72f2U101nCv/nK+kOXNcPI/uV0P/5vWoPCwVnXUO8ZTn1WhHo7NjtZh
SqyxXGMJpI4l0OuQ2JaOVzM1nI1HpronaCxoMkmowvhXrmV6t91gDEj259JB3WmY
a+0NdpM5LJbEcxHKMmnFJ4AqX9P9dZnGNIxbRjuZikQYmKIoRBYv8p9JeasZp9Ub
R4VyvlNWhVbt3BriVXj3v/kH7NRff6xocNICbKnZk3zXaOhyw4iCE5Ivj1bj2i3z
DrVf2kzkwXpKqYBVJcLZbqAFfR8EwHllkhvdo/uQPGKROG0z8QQJVirQsnuynwYE
9KI026GZ17V5hn8R32LN7JqTTs6aFJF9nNZ0d/C+jV2UMHWTxJjsf98jJRavFE22
nvlqjTRr3H4O1FhBkUiWiBiAnuqZ8dym4paMFvNZSben65qsFQPUY9hEanBpc8cX
qN3E+3o9kZSZwxciDTXO/NNUYfvsHyu0bC7KbMTjfOfgdyuUlFrxsZivq+IIT5BL
PJNX7jl+0rhSxAUUe5TseIkH11W2AYQmZXVRko1NNwksQk0Tk1ny7XAQwGvOz7FE
FkMusUHvCt3JwMXPeNSSFwEb1GaEWSYG8+wNClGb15iWXYxGdYT4QRbk5CLD30Nl
rhtNaRFBE6Bkbx2daCa938N/WJn79qW62GmhCl4yf8+L0xYJSdIZfw/pRcnhLeKV
5Oqhya9WCJkiMD4qLzYYh2b/W5BeUPcBSXJV6ose9ncFmzS/5a+C+gok+xG7XOLT
W8Ux05VHxCf70An6LkCzdkStEaBkAOLahH2sZMU8HnOlcnyfugjKqj8uBDb2NtdP
xwdHD+H45/fKooOQDIOYXdTv+zp1WDjF/IZNc+KmZFTLiu5hZGGWEnhF1uUPaLTA
wOBkrjX3V35aQs+AobBmQ+GZYRoQJt51P2xl8PwzMBDjSEiKOmuujnHwojOHJxON
+7eL12wXbFiAcgwrA97I7lycBdAknaV5pFbxydnfBiW87cLtt+OIkZ7T8YfvP6Ow
nhPLlGF87/gyH/KCe85+Odpek5Obj/T0AN3vDr7uKWYnaHW6O4KvlYLofcOe/Aax
lUfjTovtNDw5LjYYpiUn32UDXvv+7pCw1LlH+mrVsrGEvQ2osGMRfhwqszy2FW4P
JHuBECAb9P6oHWAnACfwLX9YAy+TzI5h1tLghaTjzWgJJ0EMxRuEcAlBXXAWMWis
4T54N/KtizJ+GUtRKKPwwyNYISjHX+kVA03J56u+/8mByhr39PSsbvEAVouCHyfE
AC8VhDvCx2+GXuHc5gqEOPd6FN0+k4SuSjz9T7u/eNccvB5c78MjRh6OgxIEHKAU
DUu2ylHHe+regMrb8kZxTiWZkp7YNTutr3BWw4PiTxP36dYjC8HQAHhIanLPIvP8
mpSEnujXchAZzNrvChNYPxShC7Wv71l6cGigZsvj4q0YexPYY0rA4Y5zuC8YfAUL
6DntB1k/+x7Dyflw04Hv07KEr+GQbF++0olP4VAAp7AdJazy+9qgsKA9MBzMG2Cq
AmOh3LCLm8d3PugKld4BU54rXs+JwaxiTUkVTlccs8LbTfRNpOPZnGBpg8bcc1vA
+Hxv2g0BhxQmluUSY6OiG+R4N5+4V7TA6fkDet/L6n7Y/og/z1BA84uroHrhk5Kz
1qaHau86fAiJ1yO198owqXlKLwlCGiBghVDzehN+o4P/N/wjpAw4jpJuCGQKA4N0
5ACm6sR9GClVPlFnBmlyuMdwWevIMK6zqgmVhbnfJKVjmo0otY0lZQ+7g0Uq+MSZ
wgTmohBapgJN6NIMW2ugxXLK8RvmM7nIWO+fEJTxgtnI/X1ju4w4obSF5FL5sUEh
N+aQVEMQVJbageuskpgGgVntrwet8GuC97msNbW7N598ti7OZ1ez/f97fZyQBWp7
8LGA71kFS5SRplo84KGVzjTIomx5WlpsQWPndVhbkvKA90lECfKaOD034jNvsP7e
mOewLXH4T5S2nIwaxOCyDX6/5I92MUIqnR4GWvEFhnH7lmEIQts5k0UFgV3HKjXe
1l5aCEPp7zMA+tP/VxnxOY+ZnQLp8OyDDZQ2AwXYQxVAUs3klxLQSXQdjfhEviZx
JO48u1+68Uhx+6tkIRC4xqXXm9IZDLkHTu8P2Hp0py0KfDm9BBWS+6/y92MOfeti
82adLcOjfg/xT4UDkUikRm9aajFpE2qNHIUVupjbrMOZeXVpNXwi5DnZ+QKQL8Ed
4UzXsfzTZ+MvRGfUqx75ARemjOTgmghtDrAoeDRYZY8xbP3nJuPZ1QxlXWX6Ung2
gwwY3ibf2tmAliIh5LvPlM9XP3hdfcPi3Wq0/IybNx1I7DuBtW5/McBa2dU71DTt
g/jbQdJyhrA5jcJMUci5yOiNrm6xawemWyGoaxaazOvw8vnHMYxUUjCs38zQbY7H
yIoqix+6DyB7ol7/bwrul2o1lJH45F+Lvuip9AKN909g5euHfXKAtciF3duSwbeF
le219uQksk8/JlGeV1CiNog57Gj/Fr+C8xVduWLcUx4RYRtFiSlnEowz22en2OSS
D1xmRwKheHBabt9zjlMuCQhgyBACm6Inlh9oISoWslN6tYHQPaefV4MMJ0odGYtm
qlwmlRlQZPv+eCWsOujjFZw35dOTyPcF+cyBMwHbzLaZCc1OL8LTYeO2uyHECK3j
8X8o5VGjhA83Zawy7xBecVD/fp4HCQsWfe3bonBS8M6S/qpTF/jQb3q+VQQYi3NO
D1ApcDL4zyYaRM89HhfaozTsU0p0cpNQDczePN9AI1N4u4uxtO5v2z94rEN8/Xef
JJamt5tT12AEBnV/zIrdAwMfKf5JdPp7okb6sxFLkEOxYngbE25oAj7uUljPAGLq
EOH10rQ8/9dIfZhwTuvfO1XEY7UmyCHP2b/61gysb9Jgtz/qpR63ISCViNGj5Ybn
AjNhKGg18wS9c7zKbmAJmWgd87+L6GnBgL0Wc3Eu+anfiVK/lqp9p7S4C/mr+KNK
/apCh7ckiovgvLPylBlT1ypzOw5VZDYy7pVBIPZTdVwiCvZiX+9Nf68Fg36o1lzF
RpIzWa0Il6rdmP8aBA3oqdznlFzPkqNgNT3vbDmjzxIpnRGORfjUELmsvVRYpUIX
nD6xextCFRYIO8nwxFK+xzDdFA3xHQ+kBWxlYvszGZp8IjN1OvEHtd0euRgtHq5D
w4BZuQMGfHHbw5CJ8rlIEyKGZCDATRF8BTOhhu8Yu2BD53iNdttSxLgcU5K3BmnO
ORVDW9qGDZaUtoQtDpKO1fgjB/Xz2Ne1gDkWNNvBrmem118ADbpinQP19tUr57+r
lU7vyaxUYtTsga4NCIpZqQscFa68tNUQ/AQvZqB53IRjRyPeQM70XLawhggmXi7s
znzUl0iyPRx61KQ72ColMhDcVvEhgeZL7foTmHHI1+NJDS/qj1NfCqe5T3OxHsZb
qQGpzDg+TfER0wCJigLqu8dRHliF3v+3lJWEESPIPH7aq0U4xLsCwYLFC1pPVGuY
QJQ7bJVXCTmewPRu81e0yf5ph1BZfhwWPU0i14N8C/9Ll/rT3vrkXj+h2PYPMHwv
OqSR1NJTZB5vxnp7/FJPRaPgpB3u142YFA4zoIfRmJJsqq9TUFVmUNXX7ym7ZMkt
DwYZy0INZa/yEC4lFshAklHErdN+wcXXxDT9XTYPtF+D1UBR39vzmA8BAQXGtN/x
V20EDNDbhoNomnEbnytEpbs8XYAiTIrzJFh6+8lTvZUDPoGsefZMn4I5d/6JXPHY
HXaFps3Apck2uW1vN/hnkRyFukpW78mWCuLNAJlSQ1o1DYE+sDQ4Ohycu4tTUdv7
QdHkWWYQWuVuuA+m7akL12xklSVT457Xdvnt2bGQ76iL7lPM2dZ0MRAAkcsXsHVw
HNswGYbdSth+oaoI7P3lfxpdlG9SNEMw+aWUweHHvLBMVmcI6euknc/J4dvKeTB5
ihzTQEv+PVBDitm/baPhmbUWRkQmjLQLdjewlZaXWMk=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
WoF5qvsJ5RGK6HLmYUVaIl5nB5eknYZSihswei6IXYVGlibUidIok/WTsYUpjdAh
OJF2wnVuu4Q30j9cQK3WzmrMWlwgppF+wZf99kl+05nf53NF2iLkiHDk7qYOrhs5
RHKMKVbp2nKTs8ynAoXHMrJnCwAmOZ5wS8y1TgvuArQl+lBtf63Ycbb9rsVH8pVI
PovtvUcVyBnQIOMxe7Vu6ozRR3xcuSEtiMbjDH4OiCYDjXOJcC9LP4JGbtAK72tu
uL9xIV70pTxGPVRH7J4MtFTRpPOTUMgOyh6XaljCOUgiTzbyDWMznp+UXxhgWESH
05wJhTaiNJWxNDSeeYS1zg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1200 )
`pragma protect data_block
Diirio3PqOq7xo6OcttDf/eWvqXop0mqAOuYx9I2U6gH0rIZrLqUmjzAI8zkvI74
S3FzJuq0071Z+A6NZlqyfnZ3AUVbe1nFXhtjR81ZAIKNBSlkf8nTAVBdCFS2vveL
3Nm6oaI8H/kKVtqgzIq+JruNRuH2d3+ptBz2FPCCLrxUcHakoRWVYuPmot/tnuXB
g212ROE1+Um44iu0jGMUtd9eipMv48jDTz0suo2/O74l5a6DRx353nScmCxVkjhr
otPIyBNf6iESdyPPXux1/+Gbkc5Z5pP5px3NppdlJlQwvcVJv88g0R1O2MXf5Mnh
imAJTwGPfYDoObU9+yc9Uifa7TvKPzl4a+sEdeeeT48mybpqDOA/f9Zs5J4iybcx
z3tUNRCVvQE79tWfdTvnT1ysh+0Zg7kH6nSJlT11Bzs6QL1/PKWl5b8aOzWjs0Tc
x6mXD2f0xQefzzurBfOP1y9/KK5g/Ls5uR5PZvov4sbuC2s6OHLT4cBvhhsNOTvu
KRc64ttsK2stQQBZMBhR5CCSjp31uKZES1A39ClIdjhshiiUGV02Os5GBP0da6HV
Tzeuz4FEpjIUmR+nFgNgp+O9pgeow9F0mDV4Axv5eedw6nyIZyOUBRx5V94IYtiv
wklGflq77r6A/7L+8oGWyor2y/qpC64NEdwpx+dNhjHrlLofaTw8ybGZ0qOcj5/F
kLzNKXEKYvqDhj+ZgHtFxFmHhT2WcO2bibk/MJPhGDIV79jPLoyNSUNfZKnT8Me7
aNchmtNvXPzplQ5W0awLXHL20GUNT0saHz3ylKBA3qWcaxKPuZjuAN2FB2hpEeN0
nIBZMhYunpWOQnubG1yfoNPp4+q3gjYDPKO9FxIPIXRPwxy/NPXb5zVwNEgAArCR
gQ/mEQHd9qgr9vEAl2dyxDg0IhpT+DjVUDjV0VGCxTEIkTjdXokfyCbZOBsyUV4N
GQiWPLq6iMa1VMQoujtU7g45chqdb6RpDFPsj8rUK1AOQf2+ewgyWjNBnr1T1bzJ
h9cz6+XCyqL/dsQTk9oy9qUu81DnThvQkTjWMwXthjIUOlHo8jsi54AbM6hK3RaC
Wh3KRHiFCEVMY/RQ4j/JhlM06QIuE6j1wgvyof5WUi7QEj20f0H4kMMwrBSGuWfH
Ke1ecD3eX9fGfpVu+PDBtar7ZSnNs7UeM4cCtPqQeRWVhoYOdfTLfGLmp2bqCi8l
cbie/r43jRUkF8XsN+x4Zl2pWtB1p3q/Kb8Jcm6Noyg9QDdBClOupr5iWMzqYZZA
IbAonYl5dVCSarQvbRYd1p7XcvEZSSJ9JZVyX82iUn53i4VSKgSjbduRXC66SDpS
nSv1IWHwRDi60rPldpN0kQji46t9YXsg1C4bbMPFJKYa6ObkzLl4yvwP6itVPdvx
W+lQOu4z0qivj5iTLS6vP5wJDF7yJkdp9Cpr9sSxQ+kZAu1HtkRonB6FroCy8zyt
CxAYWKqwe7xO5ZQqNME3bDthwTNyNPcUeNNWbUn0yK0twmWoE7tOK6Bi7QpgufDa
y6r0tGLd/fFA6g+bM/UAIZdnkEMVQNMr3j/x5quiF9J9eRd6qHe5YnIW/U120WLY
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
d4OSsfel5UgFCpbq8soFdSeTfWAO0t5NK7kzyhRC0x4eYOdFI4358DKgixzpCAvZ
z9tD1t7Cws/dgybegBW6gs+IsaFI8Nc3aPrW0FEYIrvOtEr5lpvLZDr7Nnpw4z6G
eBIgziioTQdqNJZnOU6i/NqD/VsddzQk+4G+s53XOPFSCKj5j618QLVXKhiNjBnt
uJdfAaySg+KGtece988HvGGppQoo/tgRQxG28vaZCUCq0DXYbPukMPd70QlpW4M8
Q2R/ytGunesdAYgIF4YvMb3v5MiGlBT7OTyT+UxJVSrWHF7dJyys+enhBO8x28nv
HJIRymQMyCA2zAHwXNO5jQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4672 )
`pragma protect data_block
hBm0j6hDakRBZ2H/7PO3slc6ukdLVyKNpWzs7nniH86wkZz0fUsk+30vInIIMH8G
lAXBcv+EXZFt6DoQ94eL6Zkwyj6WztuzKOcmtkZmffZ/S8IoZVgQRn/WpefpK9VE
V5WA6nUwZAr0oqwbBH7brue9SLbDe9fElas1GEb+3swMC3Tx7HLrZIZnbjCKLP8J
7PS6igNajwGUWTVlZjZgUkJwVpbr1jjKEYlJp5mPAwA3CggcNOaRytc6ZvaTWILR
gIkSdFi7uhUj+l2nVJ1BkZRvqGzNBfzrrCddMGULk7y+by1fT44JV/WKP/sO+Uri
+B3dKQYauS3oUwspNXtk+/65+zz49WtFcVZLHe7X4G7HQ6k/P+bfgAsnM0pxQIgy
uKyOPE8D2CV32dgrqEYZRBDcO4DfEEik33ZtFpsA5sHoxJ2xyEPVN75heQ16scdD
h0BTUJTeTrH58Te1KFcAyCm8R2Jp3aAfgIfHQ5Vgxzh5xPOq/nRcKbT+mLkC/vaW
lGpuXlPUgBGwnWwBSrCZKwhgCTLaakpmeD3hmlexCcmiEAA/mp6IneUWfb0VAYLq
9Sp2LE4xYiFT9EofpW23HPtAokCXPoQEiR+bmEaAR3xUZ5fEesD4XOMU/sYd2Bbm
ugTwd7dnUCAOyvh5XsnvgFUnnXZLZWXvHj0ew+7h/8jTu+8ZdlYLvHZ0L/yFRaT5
/mekcXnMjvgkREamsVKnX8IhetGn8qg4CDxluEiDhVUen3cB0RUt1eRBLr0oMRo3
O6yTzVx1CQtQ/FOsiMBKA9SFi5NI3h72a84e8H7WjaYxCRnyXHwA4zuJKwJW/UUy
g6nr2rF0ua+RVTqIyzBCxwazXuGlYpM8In0WT2s8P2kHvb7vYt2eQCkekKcVY7+J
uoj+rrsakzTOqzXXcCfCv37+PemRGXrbADX+8lU77fWU+KW5nW/hioSU8ukHQYli
flIMKR5/KXi1gT4+gwTJqd7251C8FYfCgXP4fydPg9sTCcHBflo0/y5Ut/vcV9H2
gy7Zf5iU4aN6XWMsczBRvwceQgd5nHDsZs+aV5gXKFGNuf0yRAtiveJktdSAj0cm
eNTHWIMB9fm9izUef+L41hEGEqljMXQE84MYYI2AWgvwM0TYhgh1VPnJ+Z8SJ4v+
hWla5OWJWily+xOLe1aBluv9prFTKcKSgAjrDY9SpkQNIIIhgGl2stUmTOK1huTZ
Au3ymQ2dbt0D+XD11c+lboJ1dCava1q88e4etddmWqjrkeLF//PgycdFLPhleOcU
18TCcsVa8kFYZqzUIf4yhEvzIbF8dmUvkslzk57fJ2FISF04+dXUXSabgSgeveHE
q0srdobS5M5zlXaeve6kDOQOBIA6pEFDIUKHbCNYgHYA/Q9hBVBfqZquqrpkZn/r
6c/n6uuQHS40k7VHiEErenub8PyF2jz4HyZzBGjTn/hOzyxB9TbJdpq3n4AWEg+C
ACIgixu+aRwdg3XZbFV8ALfCa8lg/IbLQTSFk9VX0mmFFSZrJp/PG/JuiX2L1HkJ
f7Bmk0aj7Jgr+JcvoiG338E22sbcS4PtVVwhpUW/OrsYlsQVWCiTqW0uzmJ04rNN
bzwuwyCKiszA65SdwibUYSgQxdurlmIyyic0IwnlpFCjRXe+cVokGD4w4xYH3yzD
2yHgpQ2if8W8seRAbx/9BiX86phzec/T5quGn/db7PGLvuS3f4TOafaRmHwYWbYi
tdho3uEoWmd/Z4nJ+2p7iVrERUMsoFr0ig9P1NnCSSGI2j5jR0goyKM5I3GJzZec
VNtgzwDvbtUMOEapg6Tyr9/ZI30LWA3KInugArFNwE2fDBjg/jL1gV2Wat/u10Ez
qmksQxLkW2CIzdEbsacPz2zOWFqZRQz3fY1qp8S3RkjVo0pNQ77c4LY601wG4UT7
rqbI/PW5aZSd/LhybPF0+3OzVklccWwJjxGZZPXV7VQG5FJLcdIMvbpOh4BKAZKJ
x6tOoVxC6gxQKuCFyNsKpdbZKD+I+p69gfqMDZuFMyAujJ9p038qMRzHTGgJm3ei
XtsnclN6NNUYPIhraIorgKZelAOQBD3LDs3+t31R5Dq3zgxrMGtDf/UPkThtN4j5
yLKITSDhNzQ1xF6OpjpPgTLW0lJWRuyO+cjPdWXu/mfCyFLPtEYUHEOsj3KAmDWo
yDHrrjPldVRFV3y1vA2dj0hOTgGC4uj3yfKHD6lGCzfaZaFfBKFrbYEYaZnIJbJU
ymaQJ+fGh2HpQpKZiD5o8tqbjwB+/JUg23jMnC066Uf/qSke8VuZjkBK8f/t/qQZ
cq7PiF8GLrOAl9gcB0t5tya4zz1FoYdqowcmiCaEiJ+twkSBSK9z+EpV4tuj4Qz7
vk9wTHeDVUoMyWMzXPXUNzoSM+6Y08c/T/pqBk/IzgkILheHSTLLXFyOzML1UfBE
k+tHvX5NFhN1E54dM0/VlH2LtFon1Qhkluca/+/NPERzLG6zvxEzfkFI98rHlxge
IJsc10p8Utr9ypMOESTJ+WLNsCPHgmf07MBGdDa5gVJGBuGP3MT79AX1xCAwsi2C
gZE96tsYMonX4O7mMbl35BcGcEIzgs/7gYukJLVSjf8wXcje+2OKqzwlN5z+kVJb
ibobSvhYWqMNzEwSB/H37xhUTUlhDZkWS14eS7lEXta0sGV6JAmxqZHDFA0Au9Je
XzX9Q7dAygS851mL3lIL2PGR1RiiDyGf4+KxHRDqnx48pfqi89AzHrkkfdApIu07
tiVF8BzcGABLcPVQHncp4XjqcQYZm4x9Q+rEoP49HFwnml3NgzEFG2o5Wcvc0adg
TngjXKhPwmFZ0SUGbypTjv2LsuBnRiuzF6A6IfPwGivhgcsHYmprEBLyf9lHGbN2
7aI40qaX4MGN6FSHj/r8895Kcw7NPsNghjSmY/P2JBPzqolLEe/ehucFRUK1xMMt
RtJWvwQeTSuYCGwI0sfxVNydGawiuSYhc/aeqMlUU5EhrR7fH5Dgd7GolZQJeHJr
mOk+P0U86abO0QVxtA8WuTnDrstGlgkk/WO9Je/kDva1ZMRomisGvAa6FYmDTH4O
MGLJosamlutrJl/z8spaY45K/Zjj5HVJlg+320ThnMRBOulyL0WlgiHtPsBhygv5
Cq8dRK90PfIQxDjt6uqGm3ti1G0uRGqFuesTwdEy9zP/ba3a3mZuH8L2M6GzgFcM
ybpy0g6n8MBczbRzC7F5MJSU/4aDwopt533cOGH44cejG+IUeHWDbiFf1xsYJgtc
nh450hsXv7IPC5ruXPT4F/hTxHCpMpO6pUafdbwEOJSbKhylPrYI6EnG4LzoV1J1
RizuztUTRGpc3oBKZJD9e/8XuHDyjj7RrAw9e2kNFXx714nUNx9fdO+6j3Oxix+h
TkmB5tbxXDRLbrLau7O/PcsIg531HIgOYVtSMIWt5nAHo06Gr1UR2EPbEnJo88cf
+A1SXYvA4H3Y8pZ11+5sJ4alNt+YAl61cBFdKxJJUnFIsK1NxWKxW1Rbc0RkZv9i
TuxpfcC9Y9vbN3YGH81yEG+qWrBzFMthBJRvAswTC/3W8fZKtwlJ69P6OJlDLyVZ
E193tGX/kyeorULtq1Zq25tDVUMLbdnIIP5QFPPDdPpzjkvQDUUbWO3ci0sVSydb
MJ2s1N9slpg3tNMDv5awpXExww7FPLKGLH78Bq0k4Nu+RimHvSa9jNrOD0l5x4F5
Yj5RiVERcKGdKeUOX3uPN2Qt8p6DYUTzPnB777G333S2FoyTeuodJwO+tjV8hs3P
Lt2KRvBFteHld0HT3nkAezGVPyryqvmromFprwF0VfO/H4WO0gQLnnHsbYJ54yMr
0etuGYEsbszASctfJmuH6z3YpHO7Edw2Ch7hXt8MV9wLjqreIgs6wHZbK7KThO6B
xBPeHMFVjRRgMx9LcQ9IoGwFSrWucEhgEUOmK0qQD0fGGzFhg1fUAdgMP4217j5X
H6Jx5bPYM+fzt+4PmreK8DjCQeGAVRyuKgtM5iqAXM3ud/mUIJsYFYTVRN9yUQ34
7GCS0gO/79X2qHlXvue2KKi/D+tAC7gLD1eT07HxkKFlOX4yeZTdjLr6e5KuW7Zg
t3WskX+zwec+bL3SXdCkbGX7+eVU2c+H0rleMuMhav2UUOKLbkH6sgQwAlwDmjCF
GVrurkVyI+74PvygOTM/xvy77sFGT5m7j2iwYxYnjOXU53TNrzVfqxTXIPoGHZ5R
ZTC3U094lb1khlCD/2cQY69ITbooLfmRH/y2Z+CPD//pSPH9PaNrwo5g/db7Lu4a
UTMufQBbKhEndObYvhzmdmRdAn6K4eBjeQBu22jTVIk5Lzc6YlHAW3UjPt+ox3CI
x8vcRGwsCuxgH2xXXjRV5/Ga881AdBVzxc9kdycPJtwixroTlJ7Ybj/sa1IoBLzN
1ZR2Pyh4n+0WtOFJzZGvRcOaBcyFs65IAYQtpfkVJi3cL+CLFAxMjnAe4+FRelJM
V+61BAtD5FDjpDr0ia0lrG+BuS54o2tx53622mtnr3Wtc5HguSF9uG7bcGvC1Moj
jleYZde/du5/L4PHZWMXsMnDrogr7tmv3bByXJW0+PAkNyhFilL9mwEXM/qpI512
5ndzjqDvtEr7s1MdOnN32MWf+IgFKDtEy6A6W/80XFwTQ7JlZmC4fw9wivfJyNrO
5+1jGo0nrlReEZPTLcevNWGyad37RNXxW+OKVMGxhxF8gmzd17hkIea6XPI4TVdB
9oukZyShneOdN5Xc3JQPO5UehVggz2ZPU6EJgFrzxNyEtZdveTA5Cm/XIa+DnJrN
uPoEJScb0iHQDKTH1c6/bR0351oaG2j4y74/gjd8c/6BOgtU2xu/7S2T6QFJAsOT
2QVVrvjtS9pAZGLRiB2BFHFUpqlwmjzXROyxBZn7Hv9/jbq5ecz/C7ActGyZ6AyK
oUDaksBHF/Nq/SU6OGuV4TDn3SG71KSi8xwJMXZitQB0wluGs/33XOnzFKMCDZh9
MZaw8QN8FWog3pqT8br7VrBRToz60gMmRcbcdxNfy83W31U/QohqVcG7oWR6Ntol
HLnKZZaOc2CjXFRF8Y6tuHDwePC0u5fWqa9OorwUGc1XOipTdCZe3k2aT8TCHbPB
9jNQ+0yZQnDuqNXh4+vMa2qQu1OW48Uz1kM+NrylWkjkBayCcLLcLD+e+rFwWpMw
2iWzKFeOEWt0i3Ne8EQF0WWwfkgkBA3NgpIN7bNMdt5ZzCtSBffaVhYBmp9UFXdV
Xiy7+rq0JHsJE5RiPYI0GbdrGe8cyQ0z0xDG1G6YivruBdOE7xRTVL7wMT3m2EL0
Cd+O/GHUCQv1XiXnqKjcgp+PUhfvLBXJd6M0iQ8NKXcLKiiT3bwsJ1Bb2DG9K8v1
m0y6KnhPdXVqDtgRRjy5dmvOryXVgQ7XI2NfX27WfKMmlpLcN/70tshRCe2Q/UtN
1VlGoFIs1tGMiFFwIfJA2N/u/XtbPPj9cpUlXQnUDkIn/ztpdt/vO0plPolgG0V0
1pqV4ltkRGCC6v/OXyGPKf2OilUQNR6LY1vdIkAC31BmxdK+kbwHxoYOu82A8yPW
AFNkTskRvjB5q6arSMnHBVHc0UsmypYgDqdCYnu87VBcWMDSvH6qpo8iT4QWgXOm
zQ5Z4rbTe1Es6tjqNFWccMPVPqZxZcBRjW6JP1utFKJG9sGs1WrqYKbTFgNVYhqC
798k26gNAPcTogjTYjiZ4PTmkEOSDAfdiGvv9FSdZRpij4aq/0PjmWhhVp5Q+v+V
QUtN/QQH4uTeZ9tXKxeB9xchwifcxpBUohFRTzKNvSTc3b1S8BKUPvqyv0fyhUaI
iFZ4wdHNvIdWJXMoFwN34pfBo86oxMaQJTBMW2nr+osE3S3axjy8otnZKkF5PA5q
zJTNuzGVRUdvArbEz361tcfyqmpGPTTmeu/ch6Xe4E80PVad+avzMgcf/VfEo3gq
7dUqi6fsT/N8Boi8GpUDbfxIwOclXPIX2MWJUv/EHHMDoHoeaqqe7Xqd18RCc7Dw
ACQfpsDQ4fNBACwQKvmHHB7a8oV2gz9ASXuzwpMIGBd8JoiZ1bGHNDwCKPhDGwx9
yA3JnM7Ys+fDTokwgHdwg/eBnnl8YbONoYXOLyw3dFIcSukr4JEdZ+71p4FLcGrR
bJ2fDHwPBjymaNsM9w3/DOv+UxqsDlUYi872i6lNzEOmEEELki8iVAmZwIRA6Hft
tN/a83WahnolY2Tu208Pmg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FCuaJMjJwmJPaQY9GonuznsI8rUNrb29Ggq30pPCaHrA/+9cwmUo4egYJoJosjrB
Anb6niL0DGsf/JqkwOgpVhgIGSgY83TsDECNLNBL0KeVkkq4c2sucwccKaLxC3Cz
z1CQ6yWRNkAeZyrSTrTIDy5B0L9PpaeOBeRnJk//Dx7yQpw1FYV61WO3nitbVZEj
8/dALwQ3FQijmKzJM2eTG5MNl68MCc0PiG2HqHrgbSniYMC7Zcg+85k2mRaOx7xW
k40qG0ZA0WLT/xgvWDUXAxBFW7lkYxk8LY+j3JJ44nHqTvZA7scVeS/YRMq1p/3Q
cpVIIAoc2b3tZjmREbux/Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9344 )
`pragma protect data_block
oyttPiDkWlEeptTjGt7f9xfJeMF8iVQKCU9o+pyqw52mEpjYZTBquN/0ozzwNzu2
xILeZCc9eD/kd9x4wG5VLiPzOKPcGaA47GGzL79pPM54xTb8DW9Dy2ju5txy0suQ
ME26Zbz0WIIIqgHIabpP1XCeONGqH85xN742WILGc59XljPgDtQ61u7GXk80zFlV
F8YHA+6Y9Jcwf2ZNLTstdTXiB6onP6iKjhP3IhZzW105V6no/yoDo/BbKFDXKU6v
UjIj1ziz5iDb8UT7BgluJnWeEBWMTEAcXAcQZ91tqr4nC2kKopf8pOr4Fn6la1TR
N2QFi1166FlqGuCD2iUrPJIz5o27uvKKCJG81bhP0fZUeZCk+uCp1BVwgWWS3V8T
1TVouuaHGmF+53EX1YXVPExnRbYL7aoDObuGde2G4HSLm5xHQKko/Gi2iae5l6cu
mwBu7fPVzx+Rj+JiKyPPnzUm6gto6jWySiltQaao/0TGcgplBeA9qbPXF9Rlx0T3
w3tmG9lH1ib/a6Bt5ZNmgHTCGBx8JS266NWoA4ws5qQV8YSuFVbTZj8W9LzbAgnw
3HsoPJJXQVPXFrt94fAtDMkfWn0xyEieQHbG+9OFkqE4QSndlPClyWuVCTAAa62B
RpZTxNT5p5AUMcoYpqPeVJltO/H5tZXJ6DO5kZU5WYmxoKrLAi7U30jRvyuc+TbQ
hEoO/VTBo6uzNCS4C0ubfDX4hTe9dULEFz6EYgp8yAohGAwPWG9Kw00LHBdhBFfB
synkIkucUzg5MEIk5i629Wu+sJVD7pFc6oYgEE7ezASMZLQ3WU8iODCWUWquVJdl
9Sb/gVY4UnvGu9r8uSC7b9yXjkcRCx1hU8Zz3jc3JUlpkCtcYtGQIwWFTdKwzPTE
YU8BaFRpRF1HoFYnEHJnhehvv8n37+gXMj3BDVy/S9JakDa0wEktwLzl2PTnTRoj
faYzCmUesllQmuNHFb44BFT4e7LDcnBTQfbepdc/viHTt9wYLQf5/fD6lBrAt5Bv
5uIk3JeSwgt2zbi37Tdq3LPvycEeTVbEeUlKuvUl83Rv7tF/87wC7dphagfTW+T8
oOuqq16ZytNkLbBDawpKCyMK2WJtD0seELFfOKWhOymvePY8LuU/zSbmJZQCHLL0
X6dkHavIgZoNXDuz3BCt/dlO7Rd49BQPr6MSsx/uhTp94RleD5hf0bEALtYLznxR
qVfAbPt+AKyI+lvNARr5o4Yszc81FxUUluu9U/j5SXb8vkJ31Ha9LufMJuq5lGiQ
CwpYGpzlYY3gQyWywKdosXYMquh0lqL6VaSDVYE2OLqjfmW9BYO+Q7ue6B3/yn+x
vW8V6QIljHmx43TxgbWC9YHl0s+Re4XOCkvZytwfFf8Bmj4jcNI0+YEsscRdGc+N
m/jAsBF5Tal1ONjglVDa5jjGyySTI2M96Dey5a8uleCPo1ZhimN6pr0ixzM4X4VF
U9rBf1hbwypLD5bgGyT+yHqzwyFi362elRHOjmEfhnZj+OGTTVmVfYs32k+QwANR
yz2RQQIzBriaWFKsElkNxGU6OwskiCSpTyhABXQ8DrzDWH5RJehNUYHEindU+r5Y
87nc2IJ1D2fcpo1VKFAL5o5u/PhAgZa0GI2ummow4vOqOyS+/Ay/pj5juXeL7ZDS
Ki8ni5ienOL2eYq7Ek09L1dIpOzv1b6nmt9eFRe6YbZQdZwuMUJiJAVHEfnqooSX
EOr6kSzfFgN17T3KxpUgcj+XewLp03YO3hx2ljaJ2m9cv5YlMQGKBdLL0UferyFB
SiSxa4wDFH4M4qRw7eEhP4X4Hy5YN6u1nwuVbeIz7cDYjiW8aAVOVhYlKL+X4+cr
0i0WAl5Jn6S0SAcUcd+CY0YFPibT1DQuU8r1JGKL6HUDdfQi7X1g4hnZfRqocg0d
Vt+hLrSsxwwwyJYa9Sie5JO720hC5uTX4iZGNnCdN9T2abCvdZquQ7fBXozQIVZi
hZZ6LDqgUv47p1rM6l53I6uzTjqgbcWOiOKV6lvvEIXzfzLIinRaWmOytRXjyaal
2kngFAYcMcREOEboE9eEDSlIEVbdPzQHj09LbHWen4XcHwRbDatTK9/Rf35It2ce
29V8NMxba39I3+w5W5/VRoqphB50Wyzc7eSdFK/lxh5+HxveZ0ZoIs7wDrIjdLqf
m+rcBio6z1Lt4BLcarD1MOA9rWN9/Tmkp3UHbD/HeeAvnxzBJLspPe5n1nj0ZoKK
s2VBmhxvMyXzgCF9kRvU4iCgXFD4FE8nfqGDp4Z5NlS3LKdy2NBGr1GYDY6A7Pfa
/h81KrgADXb5O2tCTqWpwRfLK2yAmF20Om/SC84VJJywiP0NGNI56nYtP4PH1CgD
MBRoiWcHgbxKg4BlmsEhwFb5ue58Vj2Lxgg26JVuQAe2ce42KkDaIcXXPJRKnBlY
ytb2LWc+H2QhGl15jbUw7zI0yGs3NghDA/TP5wZjwQGJx0aV73S0hzuPCGGRkfvk
eGQUGdFr00MS8Z3iK9aA+9y0qMavLQ1BC3W0YCSUFoJTbe/VxH7R8WXBPcppBB5S
GZ8JUgg8HuQc1Kzk04sc6KnskBXYqMQNnudH5YooOFS8vLrvm9wGBTCvtqWsUuHK
FtKP7yla0MFahvCDDbd+IkXBZfpLgAeWfC2CksoWwJ/3fAJaMTpsQfial/BX5RBc
Q3MrmDPwLly7cgy0s0k1bSYOPJ9AQ9+iJLzoVp5Go3VqC7K0QTCCRy9/9T79WrXV
8LC1s+WMbUmbmNRp0mqBeUA+yYqNg86UgQlCickOXVK8O8Bv/wAV3n7yUBbtg41z
B69W7epJL1BPvp7WTW4grYo8PXlrtWeqoLXKH5p8f+gv0IGb1Hb2C7zsrCGbDycg
6qVTknA28iMFGv4uiLs2B+FfjFanBG7prvGKz0WYpnZ+wzND6zaa0pCddMldWby5
dR5TMWm+fXNFDxFAzA2nmrUQtqjSH1kAaO/mRZH3mDW0b8WVi1TK8q9QdjJGJIa6
vKF03zbqO4UG3RPvnKXLQMbzkK8ElZD07+XtQQ0+M6F04Fl29rGV3Qia7bA7a1Y4
KCXrNVxy8tfb2RA09WeRM+i52MKnhLwoUrnNqKPdzrEi5VxYODyJseTTiQILLrvv
W/IXk1hdcfkuG6NyoKNWskzs9BKJW4DDCjluZEL5GhvePPTxPZsaBza6XiZdb9l0
0AbAKdzznz/auQO/H/TN6zySvOCMyOio6xbkbDRJAlh66+kX95OLPq/ktIq+LEsO
ONOlHsoCCItWhaJLMMgiRG127DGfI1bpfM1Gg9hQti/H4imbB7SbmPncfKwRkkuo
2KXCZNGjyHKZ7vTtX2dNJenEJNZ56cJMAqCePJpP73K/Vt73gjK122Z6mCuNSx/M
9EBZAO1r7ZWMgUuRf5ii+N3Nnj7/31SeVmuqNkkYYLhDd9g/KwY5ycSWdy4g2izh
ACXDcaXSOOcfaMzygZYXKCYFs/fhMoMDPjZ8etsohk2f3iSRlJ79M+axUb9/AX0T
is1joE1qiecy9ULb9tn2igGv0OsTnUcW0gJpuXKP3N7zutOg8Ly+r0n9lWa0epYF
GxEyM2V0k2TramYrpA2p6SOWKtjKIWDFr85GTapFlibdvBdzdmH2YlVFVhCVUZVL
6qc2Zhiy94bBZbRzF78zJeQdtrwCiYiX5ToStY2I6dswVm2NlnYd14jrlapO0nEZ
UDyyP/tvLM+Wez/s5erd3GyOoJ7bXYNUYNe+pvPwiVj21b9AthJqjP+pslv3c3v2
OZRZTimS32P84+gQOpoiEjEjojvYeYq6fIYGHQ2OR+TBk9e0nuPPUFu4znp9yX1S
vEa6ZHDQAadeBVSb1OH3znDEMV/BkcSW7IUCEg/y8wiiZkOqCA/K3kF6Dkh3Cdqs
WpzbUCOeJ0n/BdiCY6ESWNYKWgV2k/dHFfObm9UCbDV3n54ZtG4vqh2H72fNqvag
ocxFNNBELO7prAWKE6mHLKeL0B7s4ZwzDs6U//3P4GHgq6R/gH0l5AR2K7w08Qh8
ejaPfWnlK/fubm//ccsf0+0Anb5R+xfv9S4gKntbbdnCz1pCNkSLEKDkiICFbtGX
6HHREs3vBot5GrcAZUhsrMTg30XHiWYDhFWo0YXq4GQdyDVk8gKkoTxbpzbJbQjW
MY7yNq1iKVFJyAEyxWFVVjZo8mdbSROciY/jdRg2MUZnQool+bh1nH2qcDd+ztPm
C5mCD5KtEqQaBSpDbQjTRu87BwIkBVW50Ix1ygL2oUTPsP06mLEGc1us04xIVYIT
zaWR3fNpjQ9wGwMN6uTUzhG+B4HwpIXN9q0MQHOaCp1bbpy1bw0mB0jtb96Voo/A
xjz2SnhI5R+44BxloV40cQQHTUWn0X4dp3+ndtUj/2Al4IDgJy8fxn+Gpim2Ad+q
FGJBUp8k5xKY9XiNms7XQVr/FwU6xhX2ry2zd+dq1b1I4E3v9I3bcgeTJA6u+/fZ
Svr2DPjVNf2M0yGJ1EW+rYLiEEdtt92+EaNUietVUqV0lMSxMPVIB2E4+WJTHy9G
yhGe0ZhCV+zQw68DhvTAriEwQwKHMlQMbOrV94kNanvkySPJRv5+2ML16akab0nO
dlBRz+kxx2oordUXr5kE26kIyGUzjyo4nTK0RuJ2uaUIlDgmH3RX/Vlle1len3O/
jzJLTsiSimh5fZrxObkRFRABuG50+YFENEkxAM5dP4szLpdPdMgLqSGNXpcwZC9X
TPMUli35w5o0Sgy0U0ZNU8DZ31/5190AOc61qy+UsOa5uXUreVZ5JsVyq8ihDb28
WwTHI+vYDdnVWImNRIkuJvWbOw6f4GMpdXj/PAcwH4v/OXftMM4PFAH9CFMOtcar
X8uNdSW9+0SI+NBC5Htzy1h6SIL1YuUVf6HnYtzd+QfNpJLoCLXxmtzks34+yyqg
OZer9/LbAG5zous4vCEPQq3MA+Mn7lpscWdyotttu24iBWo9q8otP+AdPKfTWG7B
IiVlhyoCaYgOnGsv010moWQ/m5aGJY4U7ZXEM6Deljb2fegT4mZt+jJXgUkMpoXQ
dbxtgJIIFQEoMJewVjS0A5L8FUwGNBBn+t8SfQLrg5LQLq6/aUPBie7+MyD+4Aao
+ZHcG/7/sx/og9Mg5MfIWOvZSEW8kj8BJvPwGLLDMWkBVBnJVMaVGu32LEosz1eg
TzcSUrW4K1IlmUL00mpDiEtZTHFVnlBPZaNUfGiIMIIrhKM9ItE/n2w6uoG0LpEc
4nSrMNHDMSC2MLn3NmOGF0vctumuMlMWlNLCFSjubITTlbpcxO0gobKy4i3C/YWW
jeD16xRbAsUxP/e7aUMbaPwBNxlJyw9VbhOHxvqMLtgcun8O4RmsksskTCUGF9pb
g+BzH/i5HPJe5/9WJNYO+KK56Pfb9cHxkKok/9GH90KOZD+jasnbtI4ZpxmDC2QQ
QaaLgh1d1GtnFhSsrrGGbJM58GvhOTwnM5wvebJDqOdcIRxGwLV9gss44q7OHrEI
NyFi5vkF0Qa4tEoeXb+cfvFddfEeWToxZiMCn3S8jR57wDjxxj8ZV1e4Lzh/L1k0
oSe0jFXoDkc9MuCaztAlYqHDOnyVAeI71hcyuWUL0mS30/auS30qdl6/a5d/G2+X
GQXKQLCcxjZ58BUeA/Mjc0rInG2zgDYmHafi85Fv2ByC4qiqpccZEI2PK9FZMUdb
D2QBj6TGzWV7dWNo7uVhsWaVsKrUmhjua/udqLIiiTVifSWB5oPGfUPhwOEcyagz
vB0vAHssws6Wzlw2HB8Cm301vObxV27ZQSztsL07bDpvw2sxApFYMMcFXbEWuDqM
dGWN5kvxDpPduGYjLzOJ8Roe/TaQvIdEXv8fqugc5CGvlkXwTok0+hsY9jiAGSZ7
TMEVuVszmMwLxY5Y0i+SB8aprzBcd7QMEf6qY3loVMgOGcqvifpFLoP+rxvexc91
0czi1MXnJQGiSWZFFE6IrC5nCd8a+bkYwUJ0MTgtojNRiG7hULFpW8oW1XaxKGTy
mwLTGBu00uWn0yrQADU8YRVGr1Ffpi/gHky4ZPLzG82nh3bVFw5eS0BtihNadsWV
7FKS8M2JV8H4S81AO7/wGvlOe15OvQ2KYvoVkfNu5EB3Zt2jg9NbmIFHCeGEb+4k
C/j+74jI1uLPSHrTM7XNOniOM2+HHA03jsWMvVOHQpKmepiA7E061+uM6dBlg5Hc
YPlcpStpaB5POuaclo8k7/YmYmaGCkIdVPyGSP0KYEcbM78+tnQg1f5Bao9U63Jv
2VGCImXuyJMkE1hHgy2U14RaCRsGTZP3ymfcTDHX9qtT2F0b+lmmg66wmjjc7H6L
hdw/pb7wa6KILy1n7kNpLZfBvy/AueOZo3LSITtCX+YH7zXaPC6UwJNrG1Szzn6t
QZ5laR8o4ICrGNXpNucdEaVWg2MSNqmqHwKXdxyKdxt3HIYUNJ7K7K/PcFfj24nd
x8xUtDm8z6x0ED0wI8TLsay1v+pVT9k7zl9OulQOn/XJrINprYIeTxfOdoxJ1Phb
pO82kUwSZZU9Vz2gpYN9MiFTLC43cmP08/Al1KY+ymFVR9W8hiXPeddkSB5MpUOK
enFbLtf4Jn7iGBChX7Ncmj0mv1i8lXXC0+KPcZ6Tv4roSnWOWV9EbM3kzjvA1D0s
6U5AEF8zJynqwyrIHELeXb5FsqxcjHeOl21c/wTxQvt+ZzPSj1mMEKdky3l5+Bp9
MtFocnDLrXo45IYUvFRYeK5nllKPou04yUavJtYw1RMop9KMRw05p/2nTt09M7/8
9aQueXem1pXVjbYORsxOWdRFQm14u21fbEVt+MqopOaV7R7vULQXxqWgd54VbPCa
86h/Ik3fdoi//0dEdAjwZIwL4X+p1odJRVRnRNaK0Ck+sudESsDbndGVBJyrASUc
I+eRWRIFP9cH3XNYtsUof5KA22bAgsclQQ7waVjU682gKftx3OdQFSW5eI/BnI01
7/r/+jEzyOPdJMhXObzfsV0y+3Y7gkgTmNcal21kJ8vPs+xeukrB/V3AGZet+MGW
gxz1pOSKCtKaSjEXodL8fZ/vPidWaH+vyTSI7i5ViMzMGUy1wbI6+oyvcLJksK1N
2OFU3xYtaA53ZvHydIWBcY3okWH3W0yf8t37cCKoxuLSB2iGn7vJDYrQZBKVgtaZ
SuK2mS2MHSAvtGhQYw22ST+I/oK0Sg0tepfa+5xEEuqhN3EZOEUsbWmkdrLxC8y2
LwlyNUM17wrpR+dK60NhUiW7ruTumynmMs3RKXoa9z1Ox44s4XRPmWp0yuwCrfVb
6oo9jd8ipXoK8Blqsji9U+cbcOjbw1oH6/Qfm9wDUcvSoe4jAvYh195BmqGWtcPH
x2V4HMQ5ON0NjppyHjHGPRwCEuZuxiPmSm7wg2FFB5oXV+a/BDkKtLX6wsyYcHdA
apqDlXpXfcmokzMepPSSj5B47WxDeDg+wQO2v015n4NYUAVnfsWGdIiJaRSlaCPs
qxpkOHQP34ZNl+Kk/bIB+gajM1ybajalxc/adiw3Js5Y8ZCD0vXO2aQT+MVUy7vv
HaLWL2sMMuHfWMEhi+990jR2BY/MsGe90WCkUB4cQ51f5cOKIT4w+17AXW8RR6ot
cr4Mb+EG0NdrCPHdn8j0EroI6j066w51AAWx8k++Z6Viwmnv3Scy6g/O6SIbBYRx
Pnz/wlDCa2KNDW0dPpRO60BfkzxTd4W+AdkpMPoqGucAGeqwCBb+lz+ZHRaEbZDL
EGtiBrZ2zEImhIZw8UMoTKx4tMfigiLwhBwdiv4NpbWO3UjV/85PMGvU+OmiyIFe
4WY1zmnsu8tEz1HjB4gW+iRYMYXVX1cYRAF3Tq+AAXLTmzHPa9Y/XJMfOVX4nPrx
zmZf+xq0KN4mYdR9zRr2/SwMVA48CQIRKxyjc3NjmVxIVBGh+camsHqS7CDQyojd
awjN6Ns6ocBET81tLmOGJpngutFcNbHJCalKNLZCev895JWK5jYj1pDJhRw8q+Nh
4SO0Hh2YOVERbtcPlx6LVq83LVIwPGbg+/j1Glccygdgyq2xLcfftIOaemqu7i7f
lshTYPtGl3YIW6cJhbJe6MPu6SjwgIHFdTosdsz+/7ny7oPZSN3Yk/fZkSjIZgF0
wkiP3hQkenyLki/nv01pNS9tIPe21dAZDNfWqvjuk0GtLJNaELMPzoMV0ZwhhqCO
0TtKi/MF65LPc3N42ZbgcJpFePS4HzAze6d85a2XQXPd/x/JaDeSLNybtOgoFtLw
O1inVkVnyycKIxQsss6kZe9BxSz8A5nuhd/LNlHMhVcL+YpYkj+ocPsn3S+RIpyJ
yARVfF3W5XrnrzoUaBcjpwKR397z6yuiOgFMHTmzA7XS1XYW3n1OPK9EZRMuuhcL
24X+x7G+XOGUyOBEw2qiOizsH9mFc7o6O3i7l0sruduRdWGgAaU8ulajRTJ7Gari
0K5IedcmzfP4uxjyX202msVpsgVusmtOAWxHn6dthB4POMoMbIhL75y5FwR/+zak
WJtIqg1Xhr4Pyydm53sfUnUXs21j5KTdRPqhSHd0Hr64nR8jgTaVGC7Yx2mZgw7x
5bsiDQSX70QQR7iM/1lQRihnB5KtkX/pNm+dn8DI5qR7IHxOb4EYEF/NJmt8LQxN
t3euaYZr7JSTISWYpMFOcnBGNN5QFOTciQHMKtSzIpKIJBOghILbg60womTBJBP1
n4A06yoDVtKRjoHcO4S5etTenoyTMFooJ4d0zHA4IXTuhF1NmlzrgImTUhjYQMJK
xSvOO85bCdDo84Czc5JVKr7URqwVlCEe6hPG+mH6vaa2i97hJ98Vp3eolV5fivKh
fv+Fr6l96XSlgEiTUjXzpxvSesprgb5BG7oT3m3JEgKLQfO+3XbZIEuX929uAteh
NRbrZAbrcoM3Vmd11aAsKKBBb57mek5E8+NXzvfBZREkhUPwpbIAHXA7psO0RW4S
KnoorAsyPY/wM898/GL/6rA5eycW/w24X2JU378Xst10lgoB9jOZ/Eh5MQMh+u8H
ToNsJF2i7YLWtfPCxlJcItN10j7Y0zDtLPCz+q2mL9eyK9NLKRUS7s0dsBDMp1y/
rNTQPtOObtoB3BYH8VUS7CcZ/ulVCJmwOv5aQXrifedy3DiqoTtKzT9PWJYQH3Sf
+gAbmlh2GfKuXzhdHg+9D334n6QWd4Qa+3P5nTChE2O7VcF9Kb/6DRQhR1xrlHtz
iOEreOrspasS2mwo1864XtQh+cGhchGivhiuFzPlk+mxMLtaJp/UFODJsNmCBv8m
bZBmvm3234U3pw3VOOgXVG4jrnIqmIY9Z2s05ePfXi0F1rV1eby7bFK+iw29OlM/
1gDlLESypeeuEOQ1HvrP5tcoenk3A5Z1ZR4c/75duzXsRNlhL5CBil/25cdUam4Y
pAnVvLH5jLYZf6g2e9xclxwS7YrfIwBOgNxm8en4YFzL9/LDwzL6cxD3HbOS3TyW
+axCcHqtjr5esie+BNC5L5VPXIOXBP/0vRyBl06bMcUNXoptYcPW4nTYGkq2Is3U
ireqlnWuu94HElLPwjNR7RRawy4UTnzFDtGNA1R1IMzOlu2LAu747CB4TrPGIfqG
tcFBMQ9cu9OIQoY8Ktu/AmNxiCoO1UByJR6HOUmDbcTtb0kUcnjeBWJQOYYq5etY
xUbyoumhvJPLh9iZjb6WDkxMkBGVotHrRHpH4fNj4P/OwiWUrQy5+N3Rkca4XfFj
PxJrHD9kqR7zcG1GR4EtElUNVtorL0mcwCqpIuXQItZLONLaCGunsVq6DmQUCQr9
8F3gqtkk280tBW0cB8dSaEcr3ivDihUHQdg/ErcRQY1A7sCVlt4InBDL1PquTizx
jlGx0uL2a/+/SGyQzPXZrfzdF0y3m345W9YcoomFvXNZOlz1T5cArGswY/JH7C/b
GhoQxFIOXBEntYXrfShkQkVNPNBDw7q1tHvYmXOiWJuRJUQh9Qy0Xuxnw2pu70hi
cWKSR8kQns5EM+abmuBFvZAEEWj9nHzyi4Y5CyRHg8i9KopEM/z2M9yEHiicLnkb
9RTglxAiNH2GdShC8Sx5ju9ZdUd6e2W2MPtWf8pkWUlzyHeA60IoIF+91fsOqTRB
Pl8UbtxzK1gnYIFRmeLUeId9ugkql1Gaz2rCAUayu/xO25SimJAJS4+k/mRe/5jE
55oA0aiJIJD1MbRQ74mzCdbjW+ACCUTZ42/s/C335kWhTT8ycKQFAwLxHKEFCEKu
16nHRb1jyty2cycoQ6j+VYMZ1XosE6xudXLUoG4BUeuwKXDZXCLYReS1QRinWOLk
5NnkX4SlmNIDgo5/rB8q4Z5kJgVbpka8/EHnDoLcIgPf8OVK1FSBG4yfZ/cueVo6
zq42TwT4yQFH/dfPXXl9w9oopbFHgeH1gpPaD7Rx+ssQaoXqlP1UaVJsSdaIl4Uw
EjdSjhLugOjL5X8BI1nCmcfZoOhDCERpQzfjIRYiGjMzmSJCkDZefz7soQB3FqYK
cVb/Mb4YctQ1JZ3OXwTd635fPa2keNltaX5TIJz2m02QbJ8WfeIhDECVRINnzg4p
rfSLSzfC5/W368QkeNKWhlS1/EndygunCveQI5eb9LBNOuDrD4SSGL/RkCxKqAzX
+pBlprAR7rLVWBoLeBgpAl9CJz6a99HgN1iFL6lxYDDnlcZuEyeDO4O/Wdtv+I95
rAX47QW55ovDf8rSykMB0KhGL7oP3XwynwpAserj2TqznWma+9wChExqL+A6FgpL
POwjNF8D9zWipRFaAG87n2idjVMOmmaDf+iV97gIOnfYoyRPOjnRIAR9cUoS0bAJ
ImciJCDCuoAHjHQTZgpIGFVLbRBPQNigB4/Ve8/LdRNfakNxCLHEmsE2P730nybm
s20eGLiGrMGAuvgpQcSgvCueu08FSTYuGMJkZGL6EJUoOtf3pIWDH5XPuxvfoOyz
T4zfO552923857L8ryN+l26pxzq69UsTZ2MSZXtlN6pdM/3YVslqM05KtNAlKDEG
vykvO1eCf56VENiCWL8gPs7f4xw1MnVYr+bKR+AMSFerAPdJnbBJZF/OxYp82PMx
5vFPm4uy3xXTUObiEAy4WTebb9qP6DOPqwq2V6eySA5p+XtiNu9YtzgEdeLPmw9r
KNdyN9UD1DwtZWavap2uS2pBavrmXk84SDTyt8Oq5ynchnWxIbaPAHZzt0VVmAkd
q+Af6F8ozCN73glXIHazOuOO88BBuS0X428/4/cybwDeGI6hQ/iDFSVLUnf8a88T
399VTAfS5YkWS97Zzb+pMfbdZg80Tx0lYc4kpMKFWBkXjjjDfawZRMgg1y3tm3Jo
557Sa4CtnLMUcZiWgnYeDhOJrzaMBXU3tCkhk2UgWtsdRw/27F6Vr3Xo1kuHLspD
SUogDTluJATTkZe2xi3yw7omcfxSNuzEgQ25oxxbO8U1vqkctqq+Er8jCPs6a/1d
vaqTD+rcEl6FpqDXyZ07D9mBLU0azOiHTMs8O3qGI3PnKg+ZiCuJy7pqHS70hsi8
vCZ7+g66gSJqYGFoCZrjahDRsQOuG76yHUtCLD9Di/s7vmxrZRQXkd2RTBgLqYya
AlFgdAB5FyMH3uH8Q87tcQ/e44S+ID9fGMbMm8Xs71K+4UHsqucGf8jx9O21uyq0
RyIiv2p4VVmE4p2EK4207M6nh+p0hwB9Xq7fnLpdjDkoyfr1q7Xrcqf6nwhP5/Na
okFXrC+3k7D0DRF1975+MHLBv6SqpJTaU/tr1vKQXbHBEl9FhC5LyQS+jDW8ifkN
NFqRAut35li9PAflAuBd1s7ufOP4UY4eUDum5dVw8gjWZdwdjfQB7hDIRmdi/pCH
Gt57XOzbWZdsLV85LoABFTKjiU/3TnDdNpew3CAo3cvfobJJ9CpNyfPMh/jKc5ru
hiTS38rb4ChWWu4Ch2HDcwhkR3lgQN1QTl02c9Xt34uAQZdaICXAJGXOU/OL465h
Nv8jrSA3+rZubF2Vq1pZhTDaAcKfeAY6ZAlignHWGTP992ipJPeBjNMV7u39KTWL
tmtCBtVxcdFLiX7EhjrtSGoHQzKxLQDA81ES46BT3U1aGR+VB50EmrnZxsCiqaJm
5k0gXTVGi3bMww23q+Dxf6OemcWvlRqYWCMRNILK7I9A68GEqaE2fJngA53HPIy7
h2BKH70y6qiMUcaras6TEaqobVD+XH+BCgTFGh/bDhTI2XTqYmVEumy3dWkhcHg5
kdrSuibjq/5c/qxKLjZ2m0M1vGyVbFs/0H+DNDt8xp/lNJ0udKE+6NjEZ8VfPV1h
G9GrLPD+yoo8tEcAuHkQiBpXIzU0awkclB/7P4F9+qpZtkN/WtsZ+lI3OQR+T9yB
GVQpPYEWKbQkWumqvK/FwqiBzWPHwyzvRCQd8JtWt/c8M6TopSlVz/TXnmP3qP8d
dj4I1N0ohie9N2bMXyOq3ZoVVlYCSKZmJ0ofWSVGSGY=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BORwTtseE1hUJ4Q1kFXAtoW+kFh20gw4kczxNi5fplD2zUZvf3cOfqzACthUiYgg
+Lm3A9hIc3s/41FX04GutmVqaTjrxaVJA2fkY4YRbJ2xe++9G7LY7qjXd5323Zoc
V2gfsVkpz29jqKzwUdy0Ma+YmF8wPl7Po0nw/74NMk8e6QYkaZv8UelLCiBHdEsL
7SvX6DbnZdK3uMqF5XgGtSzLMbSYGz4Ykr+d8fGRdWlpTR9VYovLhDjn/LmkHjF0
zpIdF+dNRLQQp0I7bTR552h8PMRfAg1N+sNGqKvgxlVw6KVbZ3UVlnzCz4M7MTKH
iaH/wsX7MLOAhfcYri0zLw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10304 )
`pragma protect data_block
yBW3/BDggl8Cv0KYGJKNjWb9Hw7gfCG9KLfI6IPHwhvCjHhy7zvU93v2Nru1bOzy
kr5TuFTC6UVxJFS+WVjZEflqsu+ASayMcFzynkBIBpcmEQKbvQehe3CWISclPcPj
gYgh3XsECXSbTX+alKj5VEeUh3nj7hMiLWIu43evyk6kOnXclqpADhstmsUdxsMy
IaB8uVGHrejeuohIkQ2gtVpR/U9QvJbCntVtP45/mbyAdODzcBYUUYraxldlml+B
nkR6FKMMgGh9cznd+DPJVFfIVONawJ7VZLOM5J9dxoYt0abrn2kZcXDA/je9BON3
86b5LkY/hhRQZ5aycI5vZxLNhdl7xmQ03hV/1ZVDYZiCRhT5WDesZM9uOf1jnwg0
XSbq5eZ+2vpMxZA9Yovd0mH5+esKIAqq+Ne3YOdTWsC1vcF84NX76nzsPJVmn2na
LrLPjifQqCCfIrArbTdGd/MSlwfFCOlo2JjlNLirt8tRiLpYNEnMRALVHgIIep/2
hyJ4gE88wwPALF6QkxewE9aAFFU4K+dH1maV5KO/24jlUGE9MXOYpSnFAzFf7EUk
lu5iFLAM7Fp80whFR0sQFKlfi1Eq+WcHJSqGB89HEcM4BqnXycYe+phzkKodUqQa
rIScDP4RQngDPR5Im7xpDjqUOIPeGLD76zT6HWh92qV5AR0uviXrKTM8BdV7Q9qQ
+Ud5wOW1IRITSFKeZ7Eg6MarR+IoniujSuE7JxYYgzvjsrG5qnG11SfuifWhwwLy
p70R4z/XAnrMhMaIlS2og0xzE59J1KxOIlFDd6EDpgsfFZ/CaaOT7h05Dh2Gj9K+
WGTFEefP9YIU4O3kO6gH7klEYyP/CWR9iehirLbXMfHXe0eualOWtlwb4nlfc3cF
uVlDpn3yuPavs43hDeMRJMAHKAFRt8Qi7p3UbWN+bcZMk/sErhMGK2nGuoNufthy
lcqz911PRA74vhWx5zFEL1A+P931uYwswrp+xFNQorTCp0gblJq4E322ZYHE+uE9
DvrufOWpmw4/uaSEakKyxqP2tmiG5aDrZBTMex7+MI5uM4yGyByvcK6sWs3mFP22
Vyx0rtqotTKE9NXX5D/wx6v2H3PpDT2KHIDD6MfwBdVE9WttdS6eG8s6g/A7kDvs
UTdPkLNyzxW2Sz3t9EJP+6WlA1diPfzSFDhYAJw2JyGNVRDJ4rtkBggsoy3MW2g8
pWKPVRX50cDrOLuG1Si29QSTM+hyCaFayqTk9NkKyMVP0XTbXgDO6Ta0mm3w0ljk
cW0pqiMGtYkXsvyKERp8Z0r49FfUgV4Zfd2M7fEfiIk/N58KtovYqJr3TbP86Sqn
lisRHi+AJOV3M5fUbESsXl9iXUo8M6hvP5DJT/F1iXTOo+J3F6JngqgsA7HUqlHm
u6fN581A8k/Y8sHzbYVB0PO3KbVS3aqspAmEY1I0MEn/X1Sg12GDoCrLMrfwp3nw
xGRV51exjnhd0DQZxIaWXw/b1Gk3DD6qxWjYeBSELiIeiAgOnq5oMVD/q5vG9PBV
/ZVo0BA9PAKsXIviscAUau2bD+C4WyeVFTk3w8h4rhu8L6blPXsysRHNPbEgnpiJ
UXFRwQ83jA0ZGYfVnfUIY1vIJYsR3xj2IyvENK7aofZMX0JFUR2WT78MCoIR//Bb
j64zuI0KL//8B2p44f/vkmBFkNXHiJQu3SsuaYK2RY95xDfC8OxL38ZEeSFRq867
GtbZUl/2l3TrS1Aj0Oz4Evm5YPbCK2VRnrPDwJFETKroMUHouFQG4DwjFWo5zeuI
FonKBYUs3Mb2bLhsTr2toUwsqtkkaMB9k1Hq+zj1uBOHROI5Q2uAxdVYQWdBlSqn
mW4ALLbMEYDXjtZQahmoIgWB3/93q4c2/XIIa0fXmi9Q98iTC+sU6L7jo1Y2Utbn
NhxgP42BWAVseW0mUxJsboHlP6kOQ5RU1HxT2gxdQV0R8YkYVhEblgNk3hQNFQO7
s+nDa97cCG2d00vLeXhW1bTZG88EpAYzwC/PiPBr8jM/cTOsLFckm0ptRAZCE4qn
hZrTO/Dq7J+NuXYxhdCqrm98O69ojB0X42iq5KX/AzQ91cUTiErDd7r8kgQGAryX
ZiaTcGxmDehIT/CyWdY6bttp/Hg5mtU55E5Fen7zoYl2AzJJRIqy5dkiinWtOdTy
SpYZCXEwg+y1caW0LcT8gZ/jdaIbpm9S+q6KXTMQu6yzvddtpVa03rbtvvimntX+
R5mAQ+e06lOUAvQ+CXnFj06bKvNfm7seC/MjYNsGhZywv1ShTNxFayURHUBEcV/b
ENbyy9VrvyxiIYz4lTOjoCPHq5xtMjqzi5Oi+R0McsdVqHfNbbplJZuz8Dp6MgpX
g0sMN54wGQYcqprtwrQdTk9IrKHeNKM8fDK+6tn841OTexf+wMDSnCy+oQWg03yy
X9J0EPWh3ZKOP2R1zgVRhYhvQPFF+qu6aEYOgdjKPRTz2FYqnHKw2C1C9eeCjG24
vVOawJ02gTDrnhAxslobxbpxjFLslBzBRdr5Uk9TySNe/OS3C91vyGtrPOLZDXfk
g3DTNCL1T9YMS+5vQ6QL/vLbBr1KqUgs2/sDlSQ4rKluqvgjoX7V8tjfnUQgGvbz
lwLCLHd+snLx4Vq/WE6uMPIvikqpl8CsAzhupRWO+VCRGrOyTkK29POhU0ZfYhra
AH1A3BlNTI5SX6HIFtcPGlKCeVbMPlOIeUqln/9M9naSJolHP/0XgzzZy4gYNTcc
Exwo2y73gmd4LX/hqR54Z9VR2lkHQwiDRTCyrquBXj+7T23WHwcAc4i36vwsdRX4
8vHtko+bZdSKZ3lBWhzbTYmZnrjSZ8OwX7+G2+/xcEbMcUNMjRMSUMq21B5OicmE
OTryXUFH3WXW3Gwg4DX0p7/RGUgUVws+lCOuR/A+GNiBt9eNPlwPUhh9nrjX5gxw
kt3GST9Yp2l6mu4p/4QeCcEkp+k4Io7Ov18xFbYZzwuubYRkDIFSVUqPNGbWX/Fp
I4URa97CaQzBRhd+T8O2nxhNRmbNTRiD1QlhE1CCsbRcMz0i8ojnSe2PJBxwqF/j
nr3RQ/Wx2FeLmYF1WUSWugXwYzd9EU28xTPDH5LYSYv7l7+mHJrds+U0kK2793D8
0U60hAFZdgKDgHH+ucLUn2ExXZofTru0gKebQkxQ6z6AT8c0powhrQsGI0Pi96Yt
U//DX3HgNfRvmaYWy/X0Gxhqd6UVmtwXaapfxYCzCx2ystT9zlKGFn29waVrKlyn
wADtAgP2hAArU4docggRXcCslBjhvsHr7FoFjDi8reDAW/M8IrwzEAQ18Ixcg+ux
gZoaZMvd7PdyDjgd0Ayuq5y6ZUccqa6xNUeC8r6Jth5yjkQeqJurPGWtV1qOrTp7
OuMmLsQCqA/YtD8D6tt/JzanJ0yEdjC2WoF7tty8RBxzZ63Rp37InnmWLo44HzHf
NUG65xHETLybIPycaxGJXJE3qzoCoBNJ8bvl/1CyUdOuOQL6dk2g4gMxb7+qQQ/s
Y/F24gmCbpqIGMRP3ltJydXyROiCEd3L9DRrpd58aZ2epLWaRUse0DUvBsKgJFKz
KPBwTvXIAyo3G8BTR1ZAGF1hCuvIWNR0yQwbbyZM9ChaSI4zYv3i1hj+O8ZpfI6p
8G54mCCxrIwRoh8wBQMK9nN4M2rLKFOgzs6jlXb+O79T889CzFYWUtd++2xV/gdN
uUGBqrD93aNaFGJSDdPbUQI9EJ6M/8kctMThYBXCSIkTszuOAr8c6KipJv+yZqpn
EtgNfnXub9sKh6z+hmg1QxQ8qzHG/E0FwMIyePa+TtjHxdElS41oIfQjtYStKNkS
sRWttOUtUCUnGLGVZW4JF1m/qc1cdIabSvPytjDQO8Xssuh9KAAlCsr44s5FE5ug
gwJsvbGErxH/Le5xn6Zk9pCCeBkgLcDNrvQ6f6AmRnPdpA4ruFiDDGuhtI5SWsXq
otMSUZ2KnJRJsXxO+Vgc43v5w0jlbFIYV3Iu1pLcOXFpZMox6opvdMBPFYOIg7vf
yFRwKZcn89dYk+jtZh6+A6P+/I5Cus12Ic6OVB+mAOq8OclAdhNdrg6Lk5wBuReP
IdWW02rUBrICDAuFaUDYJWTTG3QiGnBcFGIXcW9Y3ItfJgsa2s8JKgoMCOBJcCWa
kGRNpkLgET97lGz86rAhAgU+1TOCbuGdtsak8LU5h3k0MLh6/DtbdYCynsVzVwfc
3jLG0hY298N/4I3AUFM3mMM+8M9VPGJTNOTvZcUbHEe4IwAitwI3aUfzJLM2ucz0
bIyyjTw+4C87VHNm3iVxdN5iIp3GxuUp9VsOvmtUgeEi1zst59HLe4FAvVI++Ju8
u3B7vU1Fuh1QKcWqZcZrEd7K0gcifnr3tFT1julE/CJ3vSeMF1ntA5Yi8DoP5iBY
KaGX5UiVwKlOaAp5NuuiMjjN26jT8ACXpUOEDdUq1uPLygS7aEvCjqRsgTzp4cbv
7/GUlhOTWsp8i/WpqRle0dz7wjkwRgLdu7cPXEoxckLwXo+ldAZVJRLyDeacfAaJ
X/p4v3GzKGOQGgxYoT6arpGZvGWhwoTIdW1Ue9uAvdVRpANXyoEIO1KMLrVuylKS
Ig67vKunrX4hcM3ZAydCtPE8t/jmR6SvjHQFNZvYg12Ic5/LqACsML6rIc4vv9xZ
7VI7g2OVQD88EEOoxApvYdlnSup8KRUAQTA7S7JUhplK3icQxN9fBGceuvbHZJJH
ByLggJzuk9M89j88AzEGor6onUFRPalFpCWGWRDUOV9ZRNXvfJHj85RKC8WNGiNd
5FSCY+Iu4dhJNBHYbyZHjbKBOi0I7e+aE6sKVOMrkrtalM1WeHhwqIDX+hpfoBkQ
n7F7P66Ksw/P6ZuW5BnXuoJhZVqal+iz/umHcZSboTSiwOuwAtn2UXuiNYp42zbN
QXaS0WBBcsjIHYf8OZ8EXqGRjF3lYGgSs0eiDnGNDECkT+gRoUGO//bRhH7dqY4U
SO5lPI5drQgYn768fuSR5VJMNWQ2uhossKoT6iHvlEJDhKmr6H0YtN/O2uPVnGQ7
SNBlLJrpRVLlbKBy78W+S9oj/J4hIeYDZ0KxW9tmrDUZaFmGISSGRLGxIkk0aQR4
ELeqMQTbwgoFncHqfRqQE1zoB2Q07mCncKAJozR95pVn6YiMmOkPrkZDn64Fgfs0
jzbkxlpJ0cRqCbmpbQwI2K/iSZhnmOK4KWKVs3lZGrsS/g3KE6232rH4cgotNtSZ
hirg9NVKjywWdxMkLBf/qC0byiLktTcqpVnH5UW3ylMBR8Be5w4I7ZyA07RQzUXB
gMkjQgBWyD5fopC6SIaNTpnpTXdbIgWH5VgnjJ3jy9WoxEH966s11Pjc2q23VILr
YEXuXXK1WLFWvDnm+oo2PRD1YolTCnJu+nwqHXdRsd4R7fchi+/LQD7iCPt6uvnl
325wB0y9AtAjXXafQK6WTL/HqdfREo4Itun4d8WKAA3o8vwL5aTAfXA8A9iA/h7K
TJx3+PO3GzNJnHu2pf1494mTwWRa1APFhZk+1fXAbMbzl1VHHCf+HjM4C1ceogNa
IoFNl8ARcFEKh9jTT530rviP2mfKCDIiy53hluXg51SLLUc8LTcqPpKhBO2ub1Ob
xcILvxrAcwNOmAm9vQbP6xH7AJTdE20Ol7Bi0qR+splK04Sox6kxZvByQgQZ+swn
pwsocPc6F4/q9dHFLNO9dA+hatTC5quSqPsIbszcxzdO89QZFBU/zhhsPNdje6yT
mXehq1lMMzmg5gY7Jn82uzAhPGNMT1RemnaR2qXhrhq9fjC60Q4gm0gW16m1YGIf
SL9M8V7LWhQelwpej4ktJkAxuSWQvwDf98nA/Qau3qZimHl0jLn1tJY7PVVpXaFM
NV78r0T1C1cDGivSM53u6r6eLbqvsNipv/ofXMv2Qp5RkpyQGfVVh0h1TZhNI9ZA
61hDphCgFfza+J4HV6WoCE7OKkkkw7LgWcX4Itq2oueilIKJFXpwhfKGjLGB1D1t
eHHM/bcN+ZZBwFf6Tiq59/GkMR+llrV6MT9hqP+scBQdhNEbklFJUSglsMqYsKnQ
NpzxHvQsia0p5pfjOCCjGSFlOxTNEq2COOHbMjDakx8Q8dgJLkwq7Z+lugcAH3R/
tkQ0t7zJVYmLeq7p7MS57d9pCir5WXCa9RIWS4+TY4e7/I4U185/SYrCUyaejJX0
hdwFfU5z/SIosKEjFfVWN3EF6/BQFiKBBykulC4zSVNXtGCNJ5A4FQLlWmn28L2P
2IbUn/5WbZvSBo8UFUBZRb1PTrVhxa1bzXh+KT+4IGPfJqpLWKDSe/a/dT3Vsuy1
sUi1d2+OapZ15QxvV4+Aqj8HEXC8pt1XsJx3AYRLaB2Kdh/cibM/s9X8cX5LA7jI
7s2kT7M8kNuWL6MYBGxe2OrTsPkayClkJvOhvVdC4uDdeWlOBctMTL+eW+4fHevw
G4iA1vuiMRag7Or/1bimaNBnjSoHp/NwuP01npVjSjuSXUKuokhQZErkIwF8juS/
cWIFOaGvS4A/HMwUcGDOvBND79rCd8x4Uafl1gBHwdPwcXIg+yXfcPe4+mioTkk+
3WOhVzdICKfY4Yn1jhMXHdIK0MZ+Tnz/Jpgc0HCszq5OwbhthCaP19RUJQ200guL
qBWqyH2srIuuXM006ytf7cMjS0AfvvIVYaMM3qjeDuINVO4QRwZMuO9SoCIACovO
Ux6bo0t1VDmNa7EYb24GaB3osM5kQTgZe7dC440YZ5NTYy6Tvg6GCoTCzgnjQ0D2
YPc7uGYJlCQIWXvmBdngpjINB6uOOzck9M790V/XbdtD43bMYsbLJahG8AXslPJg
3dDFYO9gqcnpSNhT0SIFUcspFZbsZ9JDscQnL0ImxziczLcdTydk4K4NHU4Oiray
3bxdV6OtLEv8LsdVxnGvjJ2BjId3xb08FGPI36R/PXrJwH7IvSerdGKc5HLIoGHk
HsPv6hBriy1y6PYJwdQj+fi8EuiMYwwKHGabNIpwKuip7Fgwg16YTNrO3EuEiceK
OzILcrCL9TW9DVQPKAEy6xEvjBImG7uWWQN3s/o0NDIZjfJeDakz7QV4LIJzjDz6
GYC92reg/VGYSG+x77fpd7N670NrH2eGWyFwh1DruSL0ZDoqNVOtGSyd8p570T57
udjS+tujq9vMSJA4t6mTb2S5PwWl7B9T1535chMV32zD4z0gpXN1fvlvfohTgvUC
RQ4m6YRepONH3N4uLv8sczAozkNK4Vtkkq/GPo6B575ds/m5IAWwxJ0KbFM8H3f5
ctt4jnHkH2YyN8ZAxO7GIntKbKYSuMGojjusccguxIRlhYgTKwSP4k5G+ddz82wB
0DXbsTj/bopukeNpx1Cz/HjilyUXO+ycnJrTUE4fxKEcmkw7v2ort5TU8xJig3Bo
p0hMJ3J1Kyvi9+t4Uyeqc4ABcLxYFYAFEvoHkQv96Y9bmMxdSLhev0IU1QI+7JAk
J5PeGyq4Gs8wPbrFOr7ENSU2vHFkhsTvZ0fFhw9PMvU4uzEiZTKO4nBhBFIIalEp
+FXJ1NY5ChH24CHUaqoClK4KcCLTapcXpKsg+e5xP9otNSvc/9IxFuvQJToL4x3W
kXxY4H2J64DLT4wAuX/kj0Lz1H6Ma3VQtXc4EDPqhuvz1tGHFUfjlwD57+IxkdA5
e4cXNMbwgJ++Zr6bPMZgXnBlB3WBbZTZ8fnzZSudPRU+Lh2scZeUqqWqtNFubzM/
KEFr8ejUemME1MS9rIZU7uqVXd3HuycXF21t2y+mlVrOz7gtQykvdxyeR0PDR7mF
5Ks27XbJ8phOaG8DAoAB7rSZgE6ynbZix3olB0ytG8ht6IZMhXl2cN382zfbXUsF
8C0Ysc6YTQxK0EhRHxNFqRV036scjRuSiMOZQelTdtxhW6q5vpfklKQdJZ8OLkf+
rlundZL4quDN0YCWnt6QRgkCtDdtP8JQSUsvm/Z65C5F4mS+U7p1GmRaOIb6hEc2
QpmOcGT72WDW1rC/PgH1a6darPBEqG35JfcxSy2HLB+qEDrYReKAzBl1elpiYeqZ
689ZVDHgtKSwxQsV/UI7jL+rffM671+COzCqsl6GDJmrmgSFMUj1xzCDywcmHsNL
3gth04rk920gDrEO3ctHDr4COBKbBbjVT1vRGNAyddwNe3K0VqoeII45NwaYsX16
whux3Vkvd6EvWB9ZNgZQYsAWWOBySH9xTEHyHRAVWaTWUDo9zfFpAua4xJu7u1Z3
KPraOpn5AwtvBGLDKTVbZzOERsO/odh5920DjJsV4fI08DDx2BZtLv4UVSBusrLH
YvbVRGtKCYVLJ/HM7HPMrgGuaH1NLiBUw4TSFANFWm5QKiD/TAHfi961WQ2qGJ/6
xDVMI+XbRgkv8+25uzCDQoU1Vw9f/co3LKsqdr7ERR45YzdwWQpzWS3N7EmMLrQg
Oqtdyfg0ste5ztYU+3O1IY281oYjekmP6uy1mTVo2TBByXKOxiFfl2zy4CWbhrdc
B8UCj5uyxeJgNGxm20xhc2DB2MNR69h2VEHGJhlE7oq3yOLqU2kSzfqA38FFp3y4
xHlf+iOX8EzuqMMPr3jySZ1N9l/RkoAI4GGku0Fz7Cn2pYNHlo7vpTeDMhBmCZ0g
fBvyvMlspC7KQP2s47XDPS6y2ymY71yGUo9fuMxDvnI2NCPHLuV486VA6pC7nsPe
HuruRStdpcEHrhPQQyJLv8FuZMIQzUYZ7v6keSI1jIl7NAQfN3pqqDS1WH4vkRmn
rg42KeUfOGe87gFAdQb+YykMynkE3Cka2R4xEyXJpQbgJz9Jb+Nj+V7wy+CqF/0T
gbkL8zGWeK8Ew8KMdCl9E9gREzFAGt9pDORjazftb6iFUBsqUpaeEVfb85jGZb7n
m72moMFA5VvJhAt6BRMZTj9sf19LHdi1B/TCwYc0mUYBltLIlviHmu8VnJQE7vlH
NyBPJKNQ/RntrUJfAVdoRWYGyYF+QM1FgEt5y6PR03moTfga442g/acmw+Wb+++c
BcsAQ8jSHh/SL/XxHAKjEZHFQUHPodAU7TwV4Jij876MmBMY5GnOj8zccMow8BK/
fyw/rTDAZTdRmxvBNpSJZ/7VVs9IxPfvK9iNDqEk7mgR33QirtRqwwqFS04siFXO
PmVlwWcjXiQeGsXLl8jyyCqGHSHEUAe+cd+weqkdvYY+7oAXqyEHNPH3kphR5bSI
97UtD+e/W9aMeIoxuobGxgx7LlqC1FTblLLi8jgDetdKQ9YnULFpXmUJqNiJWlrj
281MYlCmgz4pdCKlQlKZtLYPYjGUkR+Fj2f3A14sZSO71t6IGx03H2kpX2Vh53vw
VFQ8f6fwC+WychK4JUaaGubCo7osV+dHuoxYTaH47oJ3qCW8nah7m/Xm+fIwT5Qa
Mvy3Z9Xs4YLlOb7hDUCEp7GF9wVOV0TY8h9c1Hm9wJMO2FPTOhw92NlovW7F6CTV
PeAXb8BGEy0qx+UYO1obZsBwpKjWvDt5TOXvOKSH/t5mPkCA9Z4annZw+XMH2LN/
1dPcLH6RQlh77D4afcHRVR/BUyv/gPP8jDRuiHlJnvxqmEgF3aWJ8fh4Nyia/lyI
LW0XW1BaL+jqHaMVgmNwdmDkfmUxRo7TPty2TrudKhj5cAaKZs6Jub9Yl5x3UGG7
s0uy/XnSHgisXTAr+AGlJKAvxCYbiYfyi0o0BMc1LwvkJgy9s+gX0A71ytWFNut7
7aWErkqKJvtzMnG3myWJ+H5cpkPbu4L4P5bMVbSYwN491CYETJYkgkMv3XqmERqj
iKgkjStKbUihw17qbn+rHrzh1BhHZKrKjjIjUeFAw0sfG3UOCVI6jIyntkX3CK4U
mz+u8du4ywX5R+3amUTh+asLbvHPLSnFHo9poLVQ3FhyMz3V3GLCmSrDw0XkSzW5
wNYVeqgu/G7ithef+p8lhpEfWzBxBl3O54i5o7JbnR+i+YI1XkhEi3RSUkvtainY
X9bNVtV+tu6Wi6Bru9CD+yZRrL//Xdes536NhIxDd2OxtHahRKWZETRz114qBzCu
Dg/lqvSoYJlH6tboUbJULc8vRIbLrJiiqUSZxUVj8mob2KgbTk4sKyFGvItQYf3e
d46b+VB7RB0fO47JWNsHhNEdrh4nS6f5xcQIYGBrGkKmgkTWXXyOGnvukyifetwb
esHNgXoox+i2ZO0ybxmPSY6XSGFC3EF8eF/hye+/JSM9fnir+LfRAAY2X44ACMvG
RgZWKAwSx0YfYEfsQu9K9CkEFulGyQfNGbZw7+1cjYW5l/XoKkEh8AGk+/iX8TIC
HbdBKr4RJP4C1ejAtB7vdJVfxQ1uQ+p4eENXAonWAUuPUCo9zhEpe/3vM27kGJC+
HGTIXawIe9S6J1Nqrs4waX0NdRsBcwM8uv58ei2ummbTUYkLY2YYzed2p64XulGv
tBNiLmdOqjrYMx63fMnCKj98kXyRgnhaTKokrEQkqRToOu60Fuvd36sm2lKgvxLu
AFCtB7/LdTFa/xGgCUks6bVM4QzkfHFuHB5hfTvbWoUah1xqY2ToXoQ+9ygqG8Dn
hbTd1MO3dxGCKBQSsyPgEegfZ23Cjng4c1v7+JbE1qQQMvRZq8IwcKRr5u2gWAJL
YRb0/RrseHYW/9l+UOyVoD+ih9xa2RPGK/0LdC6BrrWSGz06vHQOe3rKxl1fZok/
onHDm0/n0t+oxIwIcDnUHiuwd24W2sfsIY3i6fSbEZDDuGfHnEFKKgr1Tiq1usuM
ZlUAKb3D9OCEBPULGPstciCGr3S6XMCoDUL/ODPl5oVvNVFmZV61LXY4LZSH/Jb/
AFSeThBUUSKr6ek5fpJZAzxOvwSZByQC4xVIcH0le2IKOPWK0Yb1mxHeLtFnRXHN
q5BrRqrTFwLZcXNPSt8ZHK0BiPm/xAIqhaEMfHooczJrRkiMiL5Qr+qHYolPD/SM
Vql4+ca4NR9igMITbaE7whK71RFVpQ7//uH/ayqozqHBe75K0H5dIz1raKuw8PWr
P1pRycBhgbNV0ycgSdlCZRRpChh9ICNllykB98ZmBZ002iw8s/7EGTCAtw6QR1CT
uRd6NFN0D/Jsj2u0svk5xZ2LrNrq3NfhKtORSOXeaDz9srLUhgGYW9lsYAAg/a1t
yws5TfezQVGO+CxPbGkgtJBbbGw+i6/qyjv5cj8e1bGlGlE9F/oe6QWQ7DesXlyl
FGtpK3l4tmtM8YTg6xqL103HzbP+vASxJCF9n4/jg8af0r69yCULXqqBo7nk0Iam
WcIb8MsubKfSyJtWXbYwLcLzBAi10gvz2ZFfDlcXEDoeRL8zZ/jxDAZI9/YDMotp
YAT6APkYHmykN6CS62MYATHPgjmc58fRkjocnPwc1NCniki0AUvSj5ZYhfTInfCo
9BWhpUGqv9P+cZiw/Gq+FWmYHXRHGAzf3WTTlBs4L11LivDSPu/O9yf6FqiChIoX
zW0lmlx6T8GReEbKS6hhFMvpYqJxYMb6HGzpgRvysE7alRet3QqzKJlduA2Q8QiF
/Gav/uUdvTLJuJtTVxmn5f3JS2VFjbUcpqwr6YbNheEqmT0p+ZETE3zNi7y2VMvX
vV82pcv276bjBAN8iJrhoLRhN2BfO1e07JjglOaAl1D7uz95Gquoo8P6FQm+Hqme
t+Tw8e7oT6s1ePpaM9ASxgvg/Cpbs27aBx1Hc32FX26RiS3ESsDkHsqHTaSaV6xI
5FdOkr9OospEZYz5i+1PpAFnhRLODUiC5jy/2Q6u8wEvVAr13LKl735LG/10iECR
53ZrrQV5RY7h25p0VsKckD24fKj46d60jaWO3STV4OQWBp4d65aSL/5Hg76bQl5V
Vvoq0ptvsYoTKjSUN5R+u/D/a8j3nPNbt/5Q4fK2vLSM2Kp0ZCVHS89LxBgX7iXs
/xITQYNiOKA4ErANgYVrFYB8BaNO9kudhyXWvhPLygK9KVnCQSyrLAn/yvRvVqnA
CetbRojDL4Ns9PGdfSqPM+ZxSx0gY5niORkk5nF6q/FSSArx4E4xrSbCh5CA0vf3
GZ4Gfsm5mxt4kK7Tvl92uq3MJsBHs1SvWmnmzVJJzghvJE1WYW7cKTzsPWpOVp/J
dAwP02CbKKZApw+8dQQoiOAs7GVl9YntP8WHNyOUrZO60wYzeR6Qs6uh/TYpe63q
v5tgl3hdoKNRz7JDuyhxCoAiGqvQW/PoVfjdiW2BU+eeq4g0RatWnLr1MrYQPGvh
TPJsvELL1nMSw0R/r3g+oxP7iua53bOFvxYi0qwjRfvZxV+hspzNZabtFUG79E0K
YivQrcPfE7XK164pDEgE9HkhYa3HVJbGVE4hEsJl1MMx2qqA3/q6Ar6wA4mKOpHX
tRtkopnWYeY8Exj4Q9CDD3k6rD1LnN1Q5Dfsbiwlji62y9vvjjbiOHXU9k5dvzRg
Ag5VtWOodZo2pD/g3kB/Mrb3HUQqRmXeCEwQhA3fdnDN3OtMxnKBzym29q4FVE12
axowmXrfBQZts6OCsioe6bMqhNvN1zwH5SVfW21dE0VZu8pjBi1v9xWVMusUcopj
tTZHBcS3xWEQ8vhmPUDjEGpBq9FOQF2mw8b7IqjX9e7phsuqxaTBfIRLA9sIla6F
8k8m9c2w3IBIyHXA+EOeEfe0d5c4DRO6RvP01EHllKTIzz8aY/4MA8fLD+kWDWsV
zGLQxjhMSYL+AF2RNuf+4SffMlBaFbBO/D+8OjVDfD11CP21MY9swMWcZxypHhe2
5Qjdm0fd6ZL4OVaOrRGSxcDz9RNn8ldoeEnJQvC3ZdAKEyVZsPtzpilv/ycW+15l
oZu8uzYcMr+EVkRtqhLzfakrN4YQ2AAigXikLyT2iFTHactK5HoqM6If7n3kuX8c
JyEQ+/p+HYRvHc5Tltp7COC/VCw7MLx2dhir5J4AtZuLVrunLbsfBelREJIlh8Vi
5pQ6QlvU5pN3JK3DR8f4fTNjWKy+Uf1wSACUsvSa6Mr9w0TpibAsycClOc3/AK3r
tqy0YCZElFmsD6bGzygazuMMx9mJXQBSH64dauDprqqYtKWtn2F4QNhs9srYum/g
O78nDYTWXd8MVk2r7Hj7fpK1EWD8tFe6HTaU07XrwfFQLLeAiipAz1TD4wHezERJ
rRvxcmd6kb5kix20WikteKJKTPrGO9qtS0ne4N/2hKb+HRd/arD3qqtWrcdQ8MJm
xY+UXg52TeQGt/YTtn2Ajtso2TFZOiK3GYPSiyNy4NtyskqgukP/Djd1XhWLVQPd
fMoMM8Ekszx4xc/S/cFkZcK1qs6rRKFolh5J3OsPhHR9xWkWP/byigYdQcIupd/8
w4YrFJqAkFbeS9iQLD3Tll0H+BoG7Zh0QKmrVHUgQeMrWVsiAV7YSCLqYguNOcfU
N+rMQgK2L8po/egs3gx8s0wEHXZleij0gWUtXpvyZqpRw16UZB4qDbeObW9pTPAS
WS4QCJkayYk4U8v828rbPxpiO4FjJpkBHvLdHzzbqwgpy7Na8uqTrDM3K+0y1oSz
AXJPfoeuA4WL9IsKGrBJdpuNsvCj2se/uSmihnOLuDrDsmFABPuQKYXB/iAQgTFR
ABriJpTq+kep/1pUVF3th6MZwgF8mRVmDttoOT0ND2oL+hef6nPfXT0hhSfldKsa
mUBact+ZwX1Gnx8HCLEdMAj8vA/biqTy/H8WHi4Da/esXuFxXZpDDJCWmOyY/waq
RXLQwo4d8SfrDIO5tDRtqyLt2zQuHuOxLUnKR03y2wM=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
INqLwtgN3dQ/efKRc/3E/G3JW5DdiD823xjk1zThTSyC5H05570Qc8fI0KT/Yxn/
cIZFcDgWZrBDROV1iaXrCjP9QOBdQ69f6Oh0PL8pESX55D9AA8ixpwt8H6Cq228o
dkmtrmU6vQzKS19MQ2K8+sj5KvbqwF34FTLy9Pap76MKrT+HPJEMRQkl1WylrFqH
CPFLdDSngzusfz1Qf2BWv5JNLqpe795tMkXVmVTorYxquiJ/cXtRV9/YQP7bz/zf
Qdg+fDYezOKsGw12UNbw/rZHaMUtZUFEUq3zHRbILr3XzXF7RhoDfrHS2YQ30rMT
wyI2KftUT9qDo8kKpF5Y/g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3440 )
`pragma protect data_block
nH8vUhtQO+auw3/9tDItrX6UOlci5R84UhZlnULhESuJI9vvEf7wxOEAc61J0kff
5xW5UBW/DqiscRy2/ApUWxXfTV2N22E0aTs2+vG9Q+T5s/oA2Nj80OuiurT/GLQU
O0b7zHJrqS1C1CdF05RuDd4ufyQqR28qkYva3mEdVQgc3GMcJUriEgKxvdsuHpJ+
9J4tVp+POTuRN+QmtGNIqpQAayHaQoMacMunU0G48hDcN5hZDq7LgpDXS2dAcHFy
g9qvnGNj9lXgEU3Pf7JeZ5ewBx2tyFNftiMdBwq+RF9NwloD7WTRM0w/VJukMpuS
DPXTkyezUvS3QK2AYKg/H1dKk60Wtwt0cMupnv75qFpJnxkGeg6MlFoUqavUcVt8
ZRDBR5zrnH2y5DHjqMBlodZnD+g1gry6A+mRiY6+Senc8x9p/pB/FzlLd+px0wVz
m9Gtw/mecVp9R5m4+Ijc0iUCAqNCtyorP/L46SprsQc0U05K6bdoXGPX+G3EoGTw
PpzK1O+5TL8siMkF+//oCILhuZQ6Z6bUBEZp1sEoJHpmsXPGMKz5csTYHUu6TkvW
ZTR52hz6jZKy3bb6k128+3sFC12pB5fyOGRfmMQD3wvYJNfCvzyh5moktAm92Wdk
2AcCjCjgcIroqARpSulNzSSxXrLdGdHUH+nOfIztVhBY5nmbT7cyfWtNwVFmKrxf
MysxqgKoDIBkCnQ3wHC8x/8ndcrtnnw1xLoAINbUpLlQFRNHZ7xXk7Wh/URFaAXM
ipIMIJUXqPycEAIbUAA9sMEi44nLXEEjpJi5OfHVkPm+TS5aDLzw4cCoZIErg5Ii
pKVhm0yPOzjxPm4GW/AhqlOTYVTir5Nmanv+aLuCPniDgd5mXKHll4j61gNkWiRm
4gC8LcSzWMwbIcb6nRJtQtshsYhE6RFpYGnWhRO49OJlDTcgptEJ0bWBv/srjDCD
VccQWKjAVvMDHtDZT9QEKygS9kCt0+d1XRJC3sqPcF9c8p/2fjEjyD0O1XTi9/q9
JTr32uT/S13t1ZDQ5a2SVQV3VA3XAzSzoRzR3F1HOLosaETifdscUYupUKQYDvXB
jSPXsrQeQMaH9cnT9ryPzLzDMdvmVn2IDVxrBnnTIwkD71wmczT7h8otNxMVzPmU
j9wTsZKX8kgIvq4SERFGhsafxoSU0/NgCy73PTBZrpMRHk5F8MsbKhbfgHlcV92p
AlSV3ulfsRbg1Y/0DCGHFyaFM5MB3MIslA+wKdNtETP0w3lWX53YMI++3PbqIQft
6E85lNIxAuIApCcLiU89hOyLpti4HbMG2U+2ZZ4R+zfYeg1wBOTU8J4tvV5WcCKI
W8TNAh80FA6fErcubf7vZEyJFS93RKnwgxIaz5+Y/e5zY1ErjUo2YMNJuWuPETJt
TvhtmCWZT5/e/47f6hZcKsDFCW9opmc2/ZS62/tPjKzgMwLAjkgKPuZLRAI1myrM
nUDGA29FVfiaC1WTAuaMT6MkiqAedOFBCjRLdFTESioaYlcC2rXILAkxVA837J0i
1gXP2A6ZCyfmiWhvRu/svL+tw7BKGJvl3pbdpJUENsM6KA33rngGJGcu4mJXI8L4
6QBYSuYaUMS/TnFNlXiAT67P3R/DJwvC+BEy3F69r9ySA3Ph8c4nxyVVg/m0RpaZ
mX7PBpo54yz7il7e7SxiZDAqHzhyWzM9mBc8aJ/3CDg1raeCbNpGbBOQsekFzC+C
eqYAs0fOW0TnT6jkxpUteaM7le7h+iESUI2gIxKfPw6iG6Fi3qJQ3uiEru58iJ27
nj93nTMwvOuua6id9Ndig3X2R2oly91vgCh/dP0bzzI+YWjNv7I0Rmj5uXrsQgcw
hSxsmJWALjKt/duW0/5tNUt9luryq0sHHsEWat68blBJyPQvA3S1tmFwRZFi9sZq
D5qQio9PgjNcu90edLqKC5N05/3iW6fnj2aPvZB5n6/nNO2FJZBcbByZV3gAT6xr
D/kHhACaCR26OKHTcOKjbQGcNPgLNDR5UdANPPZIJxqK6SaIj16iNkFbU1KYMdVo
zj+rPBoSQm8FP2Kdc9fXYsECZ5gDAPlrAbQAxSwZV0UrZqJRJHavt2CmVbK4mej4
8EiQpRZ88z7baWtfLVL7vDNL+8bmcwMBzJs/maersFrcUkb4qCFsGR3UkKCK1tiS
/HfeqCjzPnfCl97DzfFG+ngZ17xsAKFt+iYoCIeNGvDdmSj6+OlbpFSDdHPhoJmu
rz7npkLuQ8iCWWa0EsDwPQbXyiSdbuyolnv0CNE7G+l2dk4wt8m/RsJHXooERxY0
6Vq/bdVa4SI2aSoQn4ul05r4hx6gn7iuQVpU7CQQP5Me1DCxNYW3D2Cnu8x7prEt
16IlzEkrFV9ZOa8Ds26YSKlZZHVSmY5hpLMXh4+zBEH/nJWigjGpqMQQZSdUv/fr
mUWpfa+KvdcMLrE61qmi667fDjJb+fX1Nv3lIg8yMuzJAhNtIIQiR3iyE/oiaux1
Kz/Murwx887WBJaTEH58+Ktdh4+gGUvMTQFOxprJsjW4gjhaf2gRFj7P1Q4xzpMA
zsOOQpLGvMrr6KkSphSvYsT2SRVgxERkaf1kz4vlI3K1V41RRl+lVwh3atbrAd0i
s1lVV5A8iRCGS796e5uEhTQOc9biCKh4gj4VaS+qFSoiR2HPLStfI9eLEGp9WCLW
rKlecEVXU1P9KhEGD3uB5aj4LfHhEhQi9D8X/Rc2RGzl6esG/nnmPAUGCKFxjPrz
iJWqG0vC6GIgN3MeJePNcE3TO5KMT+BTFAUvpSdV9qdMCUMNpb43HRzU5Dp1vLkE
jWkWq66mi5ZDH9MuZl3KjKIoZ+7FiBrlosrF04oWWQKtdOLkUjV21aGXtglHAMP1
tQxkGegDISpZ2nIuQw7KDU5Iw7DWi/X3qOvIMSNp/vEo0IC0Ir0zLa7L8h6O9l6Y
x/97rEANT/nMI2T7N6PQODO0LMA8VJGAS+uBfrEEwiYovMAwV+ohj6QXLMiRnv8J
j0ARq46vcCQolDGjQLq+y+E97OPaG2pQ0LSCELHsmJR+P7fT9tsHH0JMDIWBVNq9
DyVtqbdInEMFAmLUf3thYNEpioc4KcdgQ/zeDKYCsLMfhbwQ8A4d7sq/aCOwUWPQ
cD0ypErkPtLBWgvXi/oym5mNpMAnimSwLKUWjMPML+I2pSAmC4wDHGjziozw+Gj6
5Ab/yvCnCpqmTuJQN1LzBN7nV6RzS2XdHVrMEdkYEeHnEwZu4na1b3XQnuQLlkFs
omHBFn5d9RurZGY8TRaMtpeAHUErtDmvtmddPRMePOdnsXrJVit67/NJ9Em/xpvx
TEls8wTm0/ucRKeMdQgAM5N4P2kRyH5AiaQUzkwP3/I4U5SnzfNAQ04x0Zfl+QAU
4rSn1Gu7HrG29LUmnGSwos7Ux2bVAN3ikaxeeJJ7l40U2ekdqwK5qpeKNCzaaW4g
7INxylvG0VCabUoda2+Lt9noCobujJa21Eza5L7uHSOhG+OXhGUvXG0zujfm97EV
0VcxWdGzI6KD6rUsrzWGRkCqXLCRnZ7fvr+dOBEaJwNds2kF1RgOiCxmuiaGHmYQ
r6S6oVklgxfvqpGje/2Z9nWYbM0rX7w8aNaC++GRcBr99IiUs49kdUJVUUIPBkL7
Sxfxb9pfkk1q3AfTEmKOJi/0B5jfA4qedmvaWAXx9QFNdBrtSduww1TWrjFSVYVH
otplir73pthpiN+TLkAed4JdnE90Ae3ozmJr3IJ3AjbqJ85WzMhXFkZ7rHU3aCOK
NvhjuGra5tYozq/qGCxHoxaTBhUSO+5+xNYpb+dhgf5EAx00xekRhsA3B0tW363o
XZA41Q9ezyexOjfXQx8PHo2miEHNu/hJdPfGKowALV+zJpG8VU4y8hU/VLEh7MQR
njDISgN21XPFsM1zuGa6m4h5FwQjHnBSZAVCgMJFh7EPjal/Y+oDG73DNX1c4Zpj
7XOD2ehIKD729Eikyxk1tb3Ln5iA5Gndl0EbzLe0UTPCPscn4iYlm4cM37ltSwCR
vNvTz4n+M6UlsJP095FEqdWU/xVHB00HlaUDkWcTXhYMzxJAGpKQDZhyCBKV+Cxj
NIC5OoiYf/hysb31obxZvjoV0zQoTj6ufZr7aWweE2h4djnMlnPUahIcGd+/JIo5
ztfnLjn+PxuzzY95Y/TwSLny7d+SqyMjLg7XwnMUN6WHpLy3erVqBNT9pMSfYBYk
+31fUYa/TOTIM3o4uhRlIYzsU3hC3vjhtD9s0tbAu4xu+G3Heg1R+6nwF0OmybPz
no2Tn1j5pZbIBN7E5G6A6G5iMkYHMY3mElTLcrveW7Y76dkJ8M+sdtmhPCxzQE7v
3Alb1IY1B2hRAcXGlGe96p9+5sSOvKo9L4dqxYDKJVejk4pTvab55yEgxANlns8v
u4mDpmh2zEymJu0yb41YvpEXbSB3k1704l18kQu076b6ZNrtnUpMTfQKbdmG1GRq
13ALUxcCnmqRCWUsNXnMV+nkDmQTZRM1Tu0QfsP2UP9/ndu5CHUvhnKt+/7k0UiW
0rrYqhqPAuei7RbqWHydXP+uDiEjWA4S0VUKDZ3Hmk4=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ntANS+0ooG5MPxJ0lyx/S0AWXU2xSPb8aUS6tvxi3kt37jltOmLsEhb6jpnICg2i
gck6oIMp+Vlyd7+NxbmAh1vt5KZZPGxrIqUUA28uUIDyPjdgTDpnASQa2DG5+mTq
wypPwIjciWLLvFY8UyP09weRPWlMqMnsluYKcKygTP7Q4mXQxBRNyYNm600eeFRi
CJ/fguLuuiW7aYRn++TgKF3mtFWJFLYt5QVS9zmZ7NYZeiPOt2jJcpp8MZdVfbnS
/z+2Ou/+5soGLU9mWN7+zzsvuzS0KX/m6GtRBQdMAj9eRK6eDflRSgPpdcf0E8YT
lHKBGZPg4lI/kAfS+dGjkw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2176 )
`pragma protect data_block
BiuVJxQO7QW5ta1r0zLoHaF6ymvRkRxaFlbTnHWmGgbRp8lnBh1xPbHn+iWiBbFr
yJl7qPkeKb4/bmSqVUV4dpcXsxchNz74n5+83GewQxLDor1qE7zGHD9PjsO9nd/e
tAQWIZQ66VDvlOu/JZFrZO7aumHqivZ49G+SEbA49n6+cDX5Vd9pwE0149sX/rLc
Fz+HLO92wJGT4gDeqrl5YLfLb7W7+y8pNNYrd102a5L0OAoUPYmY9rjXJqxJvFaw
xRyqJ6XjmZ5xEAqKWmm9EefbmidhL1CepNhybvrPZHX4h9BpV1gBsPQN0AfSEd0d
Fj4LPtQ6R9STzhocXd1sxgsVOBvMqF5x7ZmeyFNyka7x6Ite3DwXRt0rgpAIZYci
i8opjH2VAe2gtHJB+Jb6bGU2FLsQPo+2ObRXkDF5yeHT8m7vIA8ueW0dBigT9P1T
DkoLL25fcg+VCp0tgayalCxb2o4cOuNIwMAsfbcxiAuS9lasG7ob8uQbNmh1CFdN
YEseCmfuhtHQE06EJLOONfnWR/CGOVkQ3Ca6Q162w+XInIAIdPvXs9ZVX0b8qvtg
Yr2APTI6HAj0gb/m0iK6ict9KxJmejA2PYXtWXMwrBeo8UyvtYYZwxa/elrRasoB
eX4VHLSjNoWbVcK/Y0OrMxl3XYlWL8b2TgGuxnnwc9DiVhFVuWSVIqkR+ZVsy6dS
2Lj/LnC7J2j1qsFGQlBg/vl89TGO+NyM3q4uo+FvgrGMtcFHRD8bk9VZnj1XX06O
vSD/UtA+KopKEYHR0/QLNJyFACsMZ9Llx9rrcFNppMDSZCX6WolzvV4mlwJYxXc/
gxROXNcJ26852uPvtBMErRXkGHQPzarCGO/+psITedePu38+7Cg9Xtb39Nz5H//Y
4r/h1ecFHoqBwPyEC3XLy2qMm8vsOowyIWzAv+BOJ/QloyYUYa6gMovShcnT0iKM
N4EkSxUe+MukKpPRW7VVJqiJTy7e2oyDp9XszyjO/Y5iBzf0kLXk1O3kL6wA7IwO
eLP//XT4U1sBwY6HPhTAhk05JF5u1rsS8iiBHTJCPJvT/rPVUeYGSchxmbjWLHK4
p+K8xJSQo3uQEBvyrf79dt786HIHFfthrTOMJFCuOHZ8+bstatIYl5pE/tJTFwOI
H0aZx7emIIV0NjZIb9Q8uayM/9JwwZrdTggL2+3Qi5EejW/JC3Uc3vDLvaqRpJxj
ykdF0yCXIhmoiDTZMyVeTSkarw32tgY2fSJgBYA29hgzJmAhCN+y6+QZ949sk+5e
ANEr1PYOQ5p9zHEqWsMjcFZIedpZTyvyIfp9GqguL8RqNmpNUNhSPcIMPLz9wSXJ
38wOQOfAJVAuuoJ8fFccKi3Be1j1RgcUbLi69CU1XB1mTq0rg0HWPKTOGTbbNZsR
VDPaO7SXKabjYpO2oU4auGfcvEtKYZ63YDao8lkP4X/Q01ySAm+K+heZS+ecCCTt
wFr6Y0iwFnPKIM1oKUY97j9pTjOrygA3jq+SfNrbHy4q+djJm2nWY7YyyIxwfv0F
RR5clG/QRll5gQ72jfMDRYjUpXmPUj5fFiAcVKu5t/VVXx9WJ3ELygqn4kyuNufi
os4uR/XYvjAaVPz8Q7iCHj2rA0joMYNpjSFPkL4CxqAnXedWyuNOnYI8JjGdJolU
YX8yvrWEQcRVPJrXL1xEvfyUk0crHC29Sf9ZgLkJHqnEAR8/z0li24RtlRJ3DGDL
2SXoKX0lovz1qCikSZ8F2zEbbrPN2FjxZ4AwF4U7rk6WHUzB6Pg2/z0QUK6wV4M1
PGxjHosqveZPqNP622j9HBpsDv1dZmGJfemd550qonjyzWpPAYWf3ol6ulqRDwf9
TgPfWK87Oe60j+yw4jeZr2lhn7N7K4UGZ2JO6Mp5MbynTO6G42GzQ58eMBULZHSW
GgQqLBwTWHylbAgLnOAfWpbITn5IAKtJsGHYNCa/krX/dew/b6VSR5qrIMOXLsCT
5pwhGBg0TKKZo4QZoBJedI9OVwUZoghmldSiAQvvLc5vVcwfoXHDZ3ZB8+BrHtA9
ulo6AZENv5F0pcSXixHlJjolyZSdL5/D+jiqqgx0wKV+FDpwx+NfRs3UT6Cb/29T
qAQWZHw/IMJjb2eg9QpIVFSAaFDlXPX9vwDObTJWvMDwcowlkDa42tZ48d3YlvIQ
9Woi7vIK7O75/YOJlphwWYyBOPV3OliqCtpfgXgSwkeuwWLzQjtj0puzVhqhWCMn
CheNLLQFV7Xl204ZfO9omB3VFhf9pNW+IZRJGRTmLlcrXXWDdNBEIN8kn0SUR30J
XigIpmDb2Gq7HaxquB1auXUW5ywkeSJnToJGDPiSSTfOshG3y30BaPlDOZbCjg6U
HdyPORqZraLrXfcPEOFD1k6LrxhraCgiV+RVfPvNeZ1usV2nCd4RvPAdfnN3zcUE
t5vtNvz8PBWpHA8pjLTroqaE9TTlinLpoaXIYOssS7xO/S1t98ISZFtAoyDeKIPb
X1jOZwLVwDZYujHQhRAIzoAW7NQgdk9nowBxntKz4mvv810rowJaopZnFDolKVAW
3IVfBta93742yFjkUmo6C1cmYJ6G3nfYgTYzedlI2mxYFA4KF+6S8XwXVn9A/qey
bzKn/C0DJcQuR7cO2OQvSUhAZPEEpKl5EGIUFio+XrgH6rbDdU3MlqrwFgckaPxc
gi0RzpLvXG63gu9PYjy4ax4XPlDEK7dMEAmspWmXfQD6/qd9h5CT1/bM8cSNecfL
UyTVyQ1cdJan+O25av3mPukCeorAS9gQlFcmrXlUivoVcZwrtKAYz51aBcnTXSLe
pTchI3rJjok62OWzk8OWUl3Zu2c79dsRnTQ9O+SeOWJUBNTG35bCurucZ+5R6gfH
Sfv4JWeBGF4XTKV1ed48AQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
h3fNPAPEhIDIVWfdlP0JR4QGGaKx0m3u7lQOIkIZ9N05vimWre8886W0Ibu2ZCRt
5/WWfVizdwCQhDcS1DpUQAzRv2fffqx6NW50bu1ARZbgyzF84fD3nt2fSPOyivwj
iWBp1KDWeRgtyTZ/v1tljCOSU+XlNuMt6+NL1Wz3w/Ag7vjVAIrAYExQy08aGHsl
KaVeFJzkRkrHOJzbxGqf+l6T5rQlMoGd3oSpA+UdqBUFdvDHURHlpOCCUQa2+7Dy
RFsZOyfojQwHanxhAzx4mBUBQ5lq7pjtt+3eJmZZ+BDz2KHmnpD+4m82x0mGmyGV
ZegkPvv2PfATtokV2Bb5Dw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7072 )
`pragma protect data_block
rhzXCd+oPSRRbAZR9ArQaNKdSzFvMnFT+NBIsAxamYfoZBr2KEdGWeXVxYaurrMr
Y5IS0PZ06I18/Rg+yE4hYbMpG/YHcynwMD5iikCWQesdbINAG+UJkD6Y+aChnO/Y
T0F+Sk7wlKFOWocpwr9hnZudq9Xl54cgrxle+dHZRLlo6u2iTYgH8Fu2A6EHg/IH
m6YdKSQUPPuodjtWKG30c4N78SGidaOnQSYYTsgGa+4m4iBpmTOF4g2YqLp40mDi
RWnJBXCymPEMCfyZniuKeLX0FgwjSxSM1/mAOavrftXFgXBZdJheBWElcLclT3yo
9MwyaUw7/XwodC0Qi1xMCW2ulSYLupPhWkKcRRgTcbqtev0tJEIhLKlp6Gug4wU3
54kaidulRgI335vgZtDOYW120KjqDyDSDS+xO/oUFsnX9S4/8jcWKJPvegkrjvU6
qk3AJK6rD4q/O3FEXIgbPvuGBnuNuD3j+LQP0dB1E55w47QspmmAAU70H/d4pR72
/v/tJy6qphEX+d1ImZbz6/6PKMkbN/qMg2nc1JH0E/gK1snl8eLeE6TrRHqxExAx
JbwiBHAXyzAI0hSag4fpsPWdW4wFp7yL3oi8a+RgV6YGlv5ASD0oQjnonlOzmNZb
2Oz1kv6hFqCOmsLFDY3WYZV+FQZEW4tZ71gEi5kKmKuj3kRNDCdHKu2eU67vKLJB
AUuNV2p6pG6uMtdHTLTIPIpK5mBL+pWnnUi4pCkQ6GzORULQIy4f5C3FSoMdGT04
ENuvcad4e7J4XE36z5k7OUazCsWJPa3xYRiYM2VBKbVPcneWA0XR17zROCNsK/OS
sGw/JOM+OGj2vi7bx3fmdwvbdee/bA4FWyhZx1vvIaZ9n5DAszGvCIK5uH3OGcLX
BWBgYINUUmUgbq/muSF6xZwrBY2oXAhCpQH3ENAjdEbiM9YDPHoGWut1zeh1WGkg
FtX+6sUOyClXKL8ujwdI6javGV8HrdYcxKYI9ehInHSMS7GKjvlL9sfV0znvixYJ
GttEvSVqaxOywncbgUo1MO0Enu1RW1JsNHqfp82C7KQ4mbxDcpolmQF5tnq0h/zD
bO4BmIrrRpm4VwaMrg+2ih/Tx5Ao5E+238h5Tu8aIjN0h4vSHDYu8SUkj0tJUjrK
k8u4N0g+4ln+gG5+KkfkjSEJ4mCUk2uxl/M3Cup/ZPeogeC0JC/rYBhnjA7NcjkP
uIN9/jCBP4W7eZ+u45Kegv6cmMlKmX5TaKoc2zjB6AvyCLeTf7aRgtT8DR7VxqdC
c6RYwIJuGMp3qtnOv7Wgysno1mtpESO+xo/YHDGq8htld+EsdGWZ8h59iw5rrpnk
ptObWKlIfCbCo3vBRYsQ1Jn6WZzf2CC4wQ9dpeYRmxWv1bKFOb20aaJilj/EPnqA
D5Jxdf21/dIYERFigtypddOc8E63qbiLCBBBhJGuxQkalv1Ou5y0lntq9Fe31nM6
bnB5x90qXMvUL4Nbt1jkiaJPyKUMQ4gtQGVTlj2I0mzwASMA4ccts/P827paqBtD
D77/AUFddCCkY4BJP7XlxTm4Yq91IKu/egUPKzcEF+8KZIz5miV5diEiXuOeIQyp
iDYe6OSojfGrwVPss7n85socGbdvJtE+5LtcEzs99gbBzUANX8czw3AOTF0hzRre
8+PqZDFydwRLcgBg96eM2JuhlolCx6DorBq7aurVaWoMFjJ8ObQZBQeIibf1vo2S
1bvt9F+7g7MWEpl2qr8mKtq+95yECXl8ZtKewWiS8D5Y/zu9b9nz/QcPqB9HK9Tg
mZSfN92RbEc/YvS9X6wz3QwCasKtHXq48l7oUDvsCfB1VQY8mY3br0zrpHksSz4Q
xqwtaATz++3ZCN1kiAJC3ysl3xzI+s2I4VObedujo+gJCvhcaukCz99tFjjrVBiy
bdoJdwRK66C7EtPws00gZKbhlyOsbDuub0gt6v3gsItzA1Azllbud3ecmtq0dhpb
jteFvhudktw0onFmYTFpX+LZdV3cmtTKCaCfB0XaySJXo1iVgPYgdiYr+o3PGECZ
TcrH0c4zwdC0p6/gWY+rCIH+YIN9t7fXYtgW9Z0+rvbSlDWq3axYDa8AfMj7tBx9
2YJuMhBIJbCEbjqcHsmCek3CcfeUobpGTk2suI9KliQ4tNb2k1onHncXmmqSVx1N
GpFTZtdqNIraiMj8QGMXjIQ/OY/p7msthNdoYgWFW0mxfdKZoyArUmGXUkpdVDoY
526ytSTYoNiASuW05nDkW6R2eTXBeLFMFULsC2MXrppKr3nWtKx0ICGb3galriDG
BS7p4zMtbI0prY37cTlm2321QyBSsKcYNtsI+x3K+0vgJcx8q/TpXPmNw3/nw04n
hSyAjDtaREtxrr9q6mFfMrKwYwGmBI9ZzEsc15FvpEFtG8KFXjMkFZgIiHh1VR9x
8QdintukxdRaHB664RD7yw8nFTQs3IjICuW42PeV09RMDONJQdz44royU4mlejP6
5gXG81M2ZtqBOXCmijhCeZPqqmH5TdIIAvfi1AJYhD0aybrXQxC8t+t/krfPt+AC
8u4cGLi+ri5dYOA1bkkhosTsulPYLEjYPXaj0ORccljGf4YkBuaqO5BlTmRLIr7q
4/x86UXDpZJCRwquIgJmdQqjJBpynSkl7N9Ex6ucgiG+jWHTr1Jsst4k3adAU6mj
L+YkBRtNvg+60VDSuahOiM11aGjwCbYD1jyCtxDPT+4E+xIF5JUdg1b1ipDJMIgL
JGErp2U8MuNDUUMTy485F82HkADHjwuvptPfCqFMNsUUEYJA/n2nHQ0OKVE82q7y
EfXMUCZ3RtV9JekI48lYLwJumXzxy5e3mAgmh+sMtaZafurnOgr1VlmWN/I6CVqT
h3DYBhUfvuQMr7aicZKHL/nEUrKobX9wkU3POyzkK7SfNPDwzAUIS1kAidr5r294
BadVu8nG9x9/9I2m4pWIH8Uq1mcjWLvOBUP9Ajky41cw90RqLK2YOtC5C+AJMHXb
KIUQtXhzM/gatSjgg3PIB4Mv3QXbjqnNq33DIkT69dyOfgGzmVzxMoq5Yn1IYqtK
wO5Zq9F6TI5bN5trxPCtM6de/0t3xGTrMCgPr7yPZ9RPgO6AoNmAa5B9PkOkaS6u
6qJhmzsKLRcswwT2p+af5+4ugh/2A113F8b1MkJuIAgiA2K5zmp5IRChtDlCH7OW
KTeGnODLXdIsY8ll5TG+Tllnm5aVgVgrnejn7Ug78f02IsY4nhtL6uLVs29+Z5qF
g3whp2q+vafwPUxYTyQK7VrKbCZ22Um5YGufcZU7MxmZUcK/vDPepFb4N0YCT0iv
xHhr2HKMOS676zqfpcCRHgF2JOPio8hVs5JYVhEOZEk1rbiAzbna6EK4cqCIf2TI
5ABkMQ1tLjCuA3p+Zfk7Hb6xE2Ph7u7ZeGNHU/GBQSAwZ2C4u4n1Co0/s4ckTpla
VncFe7cnnTVj7xVA7zf31uN0jwXV4ma20ldDK+CpUHokLp0pYM8X6DOvdsljo5Py
Efa+82tZbMZjFXS+DCsuH/1jHWtATvh/sAkbeQaHK1UjqvAjS8oL7vI/3I7rjeFR
wn4yb5z3rjVyUpAEbUp4vevbacqQKK9j3zbdgDFeOIkOItHzUjyKO2KSVK8ted+q
va3ehjeeu1+pxrL6NuOHVGeMxNAOoBKfYHA4ldtgZP5049R6JQGnL3FGCAQYGccF
ytZB+B/ClW4y6jyWGUX0GFl9C7FeucHkACVxWceZEXP5cSe1R5C8OAKqRuacTpz/
6ef1l7OWitWfMed6C8+2GN9g2mWGXa0RfpmOH1vn8KFprnn3rkRENhXC9bYaq07b
bYAMqr8B1sMAS7aHefz320QAVJqmYfXznuU7EJtPLfrtDl7E34388em3VtxqTnoZ
wPY4yZu8Sp1ed6I8reHh4onSk4bFYVkI2/9DeR19SEQ2cnYbWk1ZQ1fcaN3Y5YuO
1YXjuU46RxrGD0g2mYEIl1U5CyaFqdmLxQq/JTf1vSFPKWYvhoRQYEvJlgHQl4hZ
V+2Bm77JQbvNrnEUYSig6ywBkp9rbayqpr+NVVEc6yRu28GQVdNKYfGRXpyTsFQb
koH0iNlWI4VnO0rCQbuebIpp5IYVKkaK/lwk+GPYa7216WdyIL0/I6zV6WL697pi
oD9b8biS9ijRFgZxXICUwAsJ9ACeM7xAXPUTjLjDdAILDVdb6MyZP5QoASu2cuQ4
Cbo1nXtFIC5TIxzMJ1YfqlZp5M1sCvaIRRXGl+gI6bBZLp7RcMEP3a/wuhATRBLy
8dD2cWnWE8vu0oc855oiBwPModxFnPu3pWkFe7kl0Wb3V0+EPFnWu721wh8thbw0
/HzJbNeIzaXLzwh7WDwWXwURoyn0igTcC29sa85qtHgDWDW6tAcszWUFv9topnt0
Bldj9Uh93qyIuqYJHR3OtpqMMl8EOhweQdI1f7dI4xfcqX1nG0bhiu0PstPPvcXt
Ydi6Aw6pUfcu4tejGfKSZp2egUtLFyDHXc0fGWbRPrYpG+VkazxHF+u58dHDSt7t
H9lUAGetFsVlj2VLGa1IU2JCKz6xpWA10OicttB1gf2xGn+puygzL7IppOsKg7IR
qUoXRHqvEYh2sFdr3Z3Bud7nifnN222cXRPinnkMt6YbH2Xeic1BNf4K0cR7u40A
8MiyyKdr/K59TyTTY8hQlJLf3Hb2Pzv3CKbdVCVysWo39ccQbWm11XlipDaKoIKL
A3wzUg6Rg8QxreJcs/GIaAv/nQ61PTw/T8ykfwFP3mW1PCCd1m40AMiUbUrMpMyO
MmxtQg0G894NrJfR+QipB2a0iAFTc/LOWsCBUr0EiYt/uERNldUHfUhTAw3NlH9d
kABV47HTjwXjb1roA+OXMAMYWzHwgYsso4DiC0XsAHDVuMBraipJqCVRu4tykSzY
nrZ25voRfaOOFopxAD1YUHZE5ZsVLffy0D+V95ST1hGcNE+V41p8Gn+09+ik1ab+
RoDnqH4JUOqzBDHBhMLrJF7vjQZ0K1YvPJHI3hPbiHOybUNjTpsg3mMER2Y8gpjz
aNOZswXgHzKVI/7+GFv0/HQY1gILCms4/nMk0KDg1d/L9geeWmoV4JxWVe5LuPJ/
yhmsWZPDhKjfdg8N+ckJ/toeu7xuJ83NyFKItwc05WyD4Sw5b/d+6dfEmxW51Xml
U19W8qey9rMw5f5mDw7xtcjCu4+lrmenkYYqLUTX8hyMMQb8IJ2fbkBp8NCky4AE
aSB/MoQ+Jv1ls0bhWqqbDvt4jDC6SHP671jH5fghPi0He/lxdWuO+JKtWRlrrROl
brCM+S+q0h+QB7brwPJx63nH+AMxq/Vnqo1+lRQJ86n628Dh6ZShA+s/Aq49jNCg
8hkjnlZuphAvbdBx/RL1N/yUsxpo7amAUtWSuOuXMn40QA3rV3VBQWyFG+0+tpXJ
bYxsmVMmcd2KcOs66zexlDfMdJg0ImUscrAM1twXZpFt3o5xUO9Q35NJWsNPzIWu
lL70U9CgzukVGr7QIglY5en5Zin/tRcZUkmDzvyphIkeICGFgncQcABfUft7kqu+
uR14cp+qW9Yd31x8p0buEP4p3ElDEA5ywxBa6guTMbTOgya69TldfOpb2iWkdbRV
76s4pZwBiQ3JGHEEIVxjW0XRI/hc+jIcNNZocRfzO1m6xQMhs8S14Qxtw1OJcfcJ
zUphazDZxV/15/dWr+G2vJkCpidaENXBJsKwE+KWb4clorvtrIhe59pjyyewwwAi
3cI2u5AgIqFfkl/PdgkT5HFusDB3Z9A/ivV6kS0uUf6OtRa2ekD2T+Mxay1IAxxC
UemP5W1SiumOAur5JYV/mD6b1SN3PCA9xe0frT3yUob0iqrT5bMMw0+m7aJytOUR
yxJpRY/+DKuYxEruHUxuNQfxYUeKhmTNF0sSMJcuxtPBzUkOFz1EI+txi3PwqhvZ
8gTnSGB3tXMuKY7/76gWYtlVtrhcD4bXdsEx7jhkgTY221yJQNnRvRGz1agoe8Sf
B9iAgMl9Usvpccl9wqSFIy7eDDSzHZqZCkZELxOLUgkd1sSNaY1pGzOMwfbj1CuQ
ktLl43peevi4fjUuzYd8qd6ESImtEVzSgHyv/UraXtZaz4oEssmkZHeLBAO/9h10
h8Sw9U3vfHR7ti4aFkkBYOVcwkKqxWomGbKr3E50vLdSH+1bsdkZgEkp8k1DEMfm
1k/TqKOs2BeUyzMaXs3O+hEZc71TnSweOYXuz1MAGrHqkEfUa5Wj67wXfSYccq0f
aupY+1SXwOGV0wyCS9EgTC8nE++w+Bih5B088DnvXGw2sZHBbUHahrLDdRBk4Bz1
OgqW+/i9C5C8Ch6nPM/cZMOOTBZ6SkMExJbk5lcRO++r5YlJ45lv1xk9wV1KN9e4
E7NWOajHNeN2HZAUX7QSxMlyC8O9Omr+EFPgQH6Z+AcQO+rUh9L9W1+kgpz7fm0x
oG+u4nC+w6Z3huYlgzba7fohpptFfvtcDznYWxOS4qrevHR//8/Jm1y1d0+yplsE
JwDM7a1IgwCnSG4biJPRLhCqIA5rInDosnmpLpd3btl6vJSKvUQI6kodSnFmUHb3
BKFvDrLWJh2mBU8YRX2f7+0YPGCoS7FULCJlMx20Fm6unh5afCefCKMfihXAWvEC
3FtMOSURm5CDPZmfv/LMlBpZ+MsUGbuqq5JzxlwlAGq/Gbi8zTtBU7ULkprSq3pU
RjwelEkbCLoWxFHlBqsmCqxYpjlq5ydwe001ooNvvkFPf90t2I/y4v5HDirYestk
nOe2atwkdESPVMmA2DTZ5zp7BYyVcF4P3RUmMSd0b2rwHrfV3YLhWPnmRTmVRUm5
MO5QNZ+ZnbdvpDLSJ9WwwHNMMukcJwsNeYJTESnYXhLfeuvPum03gtKFHBHHvDBL
ILal+l7LHd7Md8U86Qtcgl+aynNIV8LEY9yXyX/z9sxvqNFdYeJ2qZ3gqWjaFoHd
tXMfBmyzFyVbgYfdq9m+QduldoCq7NdG7dnYGDSbrWcItKeZbVXrIT0r0U/nrsFY
PoE74zYc/VsjX5C5pHPfbu7QZLq29XUGbFgOA/UHNuww3XSUsz2d8wa23Gg1OHcL
hmCoZyw5G0mBcL4Ilv4e41aUMy2g0o8Mv4FEBS8BpSB5l0xW8aCTdzz9JoH8dCpm
g4xOknTBxwictiba0Pi7laciYbrBE97lWy99UowA+IKppewNbMF4d2qlMxtppzod
ShhQTt4JYPDJX2JSO7qZUw/JZNGjoC/koNBfKO3gIYGC5oiLi3TiPY/A76QV+lin
/Wmmb4q9aoTM5/km22tg23mRFr6eJ52n/lGS7QHmKMvIRvAzrsBtRrrBBq+sjLby
8WCywDqtjp741rvDh5n8vEmxJLr8O7oDuHREanmNlV6LdMTeWS+udXdzZnyAGqdX
D/NxYb97MR5+5sZrJ09/POJrwCnLulg72bVfp1SSkTAFOSP8meCb8ibWDi6+84Ya
ZMCu9RItaovOtJmAhd1P1D5y9pm4OYsAST+M3Pp8yHjE1Fy1wbA4jkgqVYFO328Z
eA5ECEmy1BIVOoZJQfprdgM220B5yuUWhAwcTE0hvM5cQvkTvqBZ8E27g2HaVtUj
XIA+c6KfkRfE5LCCBkVstvYgesu7LIaCfR8we9q1EnBECHKYfM6T4r/XATam0Rst
xl5A673Almb/+jO/SE2Xxqu+qiwtMPjqa9Ay45liPSo0BvvX/LcrT+2Lw2JTIPxJ
fcMLqW25kRHFtUOvKmLgkSDs4NEgdy7fF2DPLgGu5eK1MysWcH8ERi5qqup8vutX
Z4gJioGrzHFKebDvPOnNwpQ42o93hhNHsjrKIEPQUZiF2+5djaCpGa1g6wVrpCuP
cA4wdYhm6I7SFDLmpgOa2Mym1YQSSRSqIPR1gK8YIiQadqwyWkTWtPbTSIvcZVpm
jTFeyDyktbQf63+QGJ3LOVSSi6taL3FdFpO2icj7Lbb7NaL6qZugXBOw9uJmOpDn
ulQd1UhWDKnlpG3jAgpsorxKuou6G+RPi8sEvBPUk1ZOWRH6TFaGglEUPISJCSC9
k04WQEB1K19wkiUT2vGZKEvWLwc4HTaHz7TpH18UJoM/XQBEUNdGFT8dPNEBZO5J
YW7qw2bXMq3tYaO3IvFihm/ohDrGv8Ei219KLZLHrjpBkD0EWn0vbF8GICzYuu6O
b65cHjRwK0zdJPeMTHVMCi/iFIJW4mdZ3SBNveTZSEGSGkLWKC+hWiG/c4whCkga
3TgOjxOZG5G/7g2J3q9R8rWuEybN9G7ZK3fj7EQzz1UMXNVuCsNeifD6nT934W98
iI7WiYiVMAr+RaUqK+2zUzTUHvEOWmw4suztR+Q7p4orBeHAld83RriHoNHo82w/
Fxe4S2mtBXQps63XI24o6OkOxkz6vGTG1WKh4QnUs3gAjD4ETJIvVmOLaGJMA8Rw
USdfjGg4NFx79puSlvkRxiA2byUuUSOMo/JMbIfXKujysWLTohNfgJZaieIIT5VB
xCgi5ZlxU/nToe1GUtnYQMT8FHtfckDd5vOUmmgnGSBsrmynE+2i7/+kQxv2htI6
afRcIJRRpPZq2ptRDzSDdTzTfer1EMKE/MMcRaD86NbiPIOeaPUAMUhSVmVEATnw
0hKSwMolMXltI0EhnpgdpL5mjtb5md0SXzHWI2nXmY94CcZ+UfGdDPmRM1V/4/LP
Fdk9CaKxLid0nxudqPDQqVxmj1Kuojt2cTubO6w7mPsGvcgUjCI39IuK0/XsYspt
yGAzhDFFOmKVdBDhxV5V0o0ip8nSQYLuIaf7OG/kvKsW5tI9aC9ks4RLD3n8f0Ev
0Ucco0PKMpoyLoAHrbrJg3B9j9MR1gd3h7ZyniO8DxYsJvdkoVy4FSPSww/ih8gI
twsQKvnkD5rIbbUhw9Dgxrnr2gwn/r5/y8YVoczPe+zj4de23JRJSYeAphbdZXST
LUDBjWo6ma99EChwZe+/m8QOjW+lR9bef6Dq6cXBZAxBwfFFmJjmMoZSMlCEDpk+
ctYYJ4KAsxT5cKN7ux7/TjUUc8NuUYBB6PZRPy5fxl3t2UAXBv/936gY090SV9BM
H1lci9uNBoyBrJX461LvqrHuv8OU5oVs7taB66suwY1UuGn4AzI+ffRh2s/KxxOq
6tdZud0xNzZcwBqSj/1bSx4iiiBJQMfmkK/mZQEj2ecp+CgXpU5rdKy/m7/QTW7v
ddwT4kqR+LStGk0mDPBN2qPQspu/7XlehXSJXHqAh3EGlbZgYtD6iuQOhUuBkzbb
7YddCr5CIAT/XDXYSeUJJYu+0bjZ2HcxwzK1Fhv6WuzQH75aV/VRIMuUWBbml5K4
VqsE76RNpkOTrm2y9G1AGORKIlC/hJFa5SIOjODgUJalvtEHR5518ZMzBtE3p1D0
RJtQttz6j/St8m0TwU1Rzg==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
IuspShdI9etovQNPY8sDfwZbnendrVDGq4Ex7HozuLLAYvRAgY0c14ORQHoCXSTV
vcc9QjF74AjUrpI5WJO4rdPCb51QJz35lEElGXMvDeE6rdgQ+MSilz8BbhPyKJ+I
UCz/dYt5uNtjIAACjk2fr759p1jMfrRbQDMGSmw89AiOOi6NoQqRGpJnE/wbnXcO
rGv/xMqlNGdu+MlNJJYqYS2tkXCbA+bgA1k+zaFR7PK/HMe/Y63ZeH0Fu9JEW9mY
MJn0cTShRx9uthvaXinsDjiwlZvDT7ffuhwBdyiGcNp6TEjhRoh2VAb+isPQUipX
iSJVPBcAtqDRux6lAksAsA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5424 )
`pragma protect data_block
OGqDAOQhjC2rCsg4sNAdscfBspB4iVMEbV0YoxUk93k8vh1pKvJOQowwxjn8N8Po
4equI5NhEImuKuk1xrhU10UpCQxdXS6lA+90SJVGqCV4PBgNebIMkeWv8CFPYOy6
ZcD2EzkytX6TRlO+K4y+49yeU/L/JwkcU3kHqSlcSG5Kk896NQFXd672v1DExsyP
UZwkfOLmhktG6K8hD+UmPVuRSIgeHZD5vIni5HsutxUYuS62Dhwi00/7eR/9dv7r
nQwIfal6hPPwEGkBt2bmhJDu6IBhVAkAsLPPpumW+nkS5fWs/SQdvR+kqr7AtszP
qr4GTsM3E+wyQ3pxPK+CQDkdJ2oSopbroBUuYdxSh9DOmrLcJmF1udpezFTKTRHC
awQqg2sKuDU/Hn9bGqrPuSZ04vDTSm1vL/YAAWuZvn2Ej8KFE2o7GVNAqsMde8on
sM1hbkfv9H/FuVfDqy80qLo75PBGROPG085+hEvRoRPGlEw0ucue7csKPXXfmFl0
upDuxHw5TRMLq19hxSWAT0GyZvaz37F1+TfvTfTcom37RStZVbMo4Qk3LL7T7DLx
FhU70QRIh5FhwK3GdrCdBrAZWWeDVsVO5pjXpmis8a+7uJ7v6LeQDaXCqKJPZjYG
G8rNTn6JL5IzrsgMgJ9NR2C74phEN0pwoWrEIUOZDKFXja0AGsD2e+kmG0jttX82
Vg2Z6ATOKBZIPudL25O2NZUqmFuH689pnUSANq4WEIJwjggqg/4AjSRLEWQlJtIb
d9Rh81f6+bQoMpt4HpZZErzAhyyTJjGs7OpjZg1JlWLNXA4wiarbL1WIQj6Qfbdz
ZiZoh+sQj32jBEqqObpDSGCw//2RB20oUcFEQjRM0SBu21u5LkzQPCnXFlBV7fzD
5GVgCJ1fgl/J3VjnryfC8IyG3OxDc/mMf2BJucbNuhjdxIQgPiHBxNy7dj6RJlbn
TwpO/xpXwkuBC+N7EbLjHhDXEhSadFbt61VPSJd4Nb03TsM2n9JXeferYzxlsxAs
frccNBcaiw2zJbKSTwINjTHb8QmHJWxh3HVasHn3vWY357C7NhJHNhlrHAPs1X3t
4R6zdndtaYchvJ9LFyZan+4jrTt7Rvy064E9j73fkMZmX+8rq91v6Z3x5MBullzj
o/LIfkZmGiP51EHsRONCK1pMrU9b3KwV0haqlkNgA6TmBQEpSVQ1yxEARVoK8NPz
ZJdZl47BgC3AjAAcgOZSenudWxS7Gjt05wRpM6OCG9bhzSWWv5qdS9JR2+1bbwOk
tdpDAih8sWN9m3LhXCJd8OKZLhJhl+RIsdCSjR7+c0V/mRjwBTS1udhhr2ncFmBT
TmmJrV4ufZn3sbM1quYrHOQ5bjf23gWP3/d/NGCBiFhgucB58xq1aRozHf7+swQ0
nffY3fQldmdq1ndAMU076oPoDn5cxlLLIiWMsEouOPpQceWTek0uxDX748bxMqsy
m/uGulCFPecqGQ4zg1SvQCNh1iPxqEi0mUVM91eZAaAynrWi/slx9jTONRsFDeFd
Bl+vwiNaI0aZevbWWHpS01LnwBzTi9SIXHWk+Xm+49dot5Vh7jkDuHKmGtMcVlJo
r+ccHnv2+7CcCshH/y0+9OspLAkaxPYUknWo6ClGVswhD7Mo/rTu2bDO5I2ICfT7
M9BIGf0VvXQaC3TATC4Ek4XMQd65TJ3au7YGLEwNkKVXBXIHVIlPeMI7TxWWpSen
79NDTB0YFtOnLoU/Osm7P2B6cCPk1lja/KdU+lRepc+L3khS6iRohm9Zsb5u4bSm
ObXgG1SGOV5FB7AgaZKK5cxazdCFGIQKFwjA78hTscDRS7bRuivRCAiz0PXT5wjy
xKua4+tssGjBGahlqUXt0EzxQF3kUhQ9ia8sbVBTpYQiRYCqGXgloHP/gYvZ0dua
ES7dU5aQerwmwTxL2e4LSEp6e+UyrNOblOUxw3o05MaDRzVxhhWb/216doFJB6W3
QZKo9W2HYthuUGsYoMDeBss+1x/2ks3Nj9AjKgobtm7M9mV+iB92Cdus7uZ00KQA
ZC1Xk70q2Yav1ggrl5e6nHTSPUVH6144X7cdl3nZSUk21zU4WyQvltI1w/UKREGR
Id98TMl/V5dUlTnaK+MWvcK1c4nYT5ivz5AzqsR8MdhU6yOopaERZbNwNo+35rDB
xgco598RlF/sNscUlaY8ignHDeoY8RjKYnyXVtQ1JmbaDGpVJtwSlPJJJJvcnTfs
3gHlLmyG/wgG0ZSsPkfDfkXPlr045KLDowtZgBxZiMgXK1+rl/vgOaB7DH1qVKPj
5++bEOFs7LjcvNllCZa6tF6QxaQ9UBzeX/ojd09RiGaQGLmEQDta7KcWB6FR0tsr
Z/3aHTcVhhsMqLxUO3lc6hwUeW+Hwen6bS6lhwc9Vk5JS2C1SNEskf9JA/kjoua/
wApKp4aS+Zsf4UhXyuf/sC8sbaEP9V9Fn9NOz9EiE/5Y5Ta4q8DJ7IQZ4O243QCv
4pd5rHBhBstKrJ2wPuAAoBCkY9i4teXL8bd0fiErKrky6ZVmpYw+oh1+Yi2tCuyn
WptS6baydfHy4azE2TZjVGrbNm8UTkxIZUt60RqiOjRkcVkaVVe5DqSGc2Q1/fGP
TPEFQ5tmEo4izLYZjl3rMz9SnIZfbC5FANAx7NZoqtlyPc2YAHNJvc/lqv3Bfu+W
d+nhoTqnJp9DZazPoV3i33oBJF4aQgr04aPqh7q7J2NCwpJPqbx+31xTGNzU05xt
fR9MHUJm508gKp7aCqwQGpOxC9wQhCReKvku+C0VVrEwLg46C/sLFnfLGJBElfmy
loh9h0n/7KIqQLcWbJKP371stjqZwjtF//X4Hcl7bXJazZlTolWmD9qzbdiIWYMB
LimA7pNBC5EboZCBg235MmXThvy2wW5/9LOty8okTvpjQ7NhoE3pEqslYUP7xnhZ
+w9xZbpp6pCFZ3HgRIbWThwTxHRtq7FRNw1xv/aRegWjRSzuNVFMsgOZycfPk+rE
7kfoeSKdps2aaRTK/QxWvmKeAQMqEqAT7wCRSm1pu8AsqsKd2wnzGHJG0We6jjDB
JMrn/TdR9sa6sqH85jUl3AzRv9jcwsmsApcTzjCJpHp/Wi+I8842bjDB4bbojUYF
uZcusgXKHRVUMW9JMwnPZSseXxzsZaqDHvoVkzUEI8Hn1liQ8JtanHEA0ux+sbzk
91AyeRP10m+ZC3Jwe4JYtobJS+ZYUWKEdNl/E6ZPX4TMkTx3UwG+bPxElR035k/T
TjhY61McHM/kB5yI/MiV/AXSRF+MR4HcolrVhOlSx+excTZEBNzSe6rVLSM5yECG
CgKCgCuuA1DYcYTt0pa6xd+Q7BcQvqgtdNgqjqDG2zUHfjVlhu0ipm2Hr8NOOhES
6Pz82sRldaMLd4fbRwWlhoF0RZscJXdQ4SKedQUeYXaGZa7G6p3EyoEvIruQQb1I
83R4LdLHFW+fPC4arBFF85WFKu8dUw7hKu3nXIvEn/37oP641R5qb84Dl+Ps+5kz
NAmxByN0YtpYIbMSxh7vDocl0cW9lWlNQWMBv5TioK8iZj32G8zcOXIZ/NOyMXW7
/OVaOYoh/6kPLEXiB1whNFh3ZOpdm6/e6MfPoxdWXUs9DF/bIkzXPOXG7CiUYo04
O91P8Uc2ZxV58EDpHDv8pqzkcCevIQw566i3HqliGT5iJaotauwR6HrOacedQYY0
2B48BJCCZDWYlXBpUjaIvou8z2tAeB0qgx3X5L1bwSCcGqDPnVI1XpIySjr9tqBp
WZyn7kDT0EexBMN5efS1+tp0CeKPL8ujvQ9EBJahIrfKI1djH/T9TUc2z5iXRBOI
WL9w7MJHmK7Uayj5YzUToEzpCac0ZdAocLsokxnXkgnK1RUNTM7sLExh/nc1SA/u
3P6OzgiSjsr0G+T3d0uYwUAi3BMq51E5EKntM0yhHVq15CxwBnyrcQvwKdtdr6ny
0DWmmPwW2A2fsy2QYh8RRL/Y2CIuJXAzS4DOz/88Onit1/2thndfiE4OriOWBY6b
OtiopuseAxaQTdu37isAvEgVURCc7xnUsTHEkyQSrqvRLbj2n7lkIb9NBFF+WMe3
Jzqm2iFATc9NZvBZDnU/dxU7DDanV3rHW8duiBxOoRkPc7Bg3+G5tP+fv11CefyN
QvNXrpbJXHiPTlrYsaRwnczE5wTnNdeNY2tpKODyShm5XEY07FRiBOjpmNotb4JS
tdmeQWq0H2sZZ2YahwRtlylgYUdVPjA3MXRxeoAF3OoRVvNxVOVMyGTp6AXJAsUN
xRnPbYG3VcqGvySCY1fq5tLpN+YePjKiQfPx3CuVzIdKc5xk6Yej+2JYwb7Tvtu1
YPLyID39OntBoJNb7KPVMLvLrfXWA+Kq+Siv+sKZcc/L0d60PC7t2j8sb8wHOz3e
iC59kZCj4UeHv6VTxGZY2dMJopCm7uhSRRkAlb8KCfwyIbGLrHeW7X8cOGYzEIA3
fMAQ9w8dxsJSNa5tBiKl2BizvrLGES+mqMU+XLnTVRXZRy40Jgr4510/bh0coCIh
zMqQ2v01svh+qGOisMFvx+U9/x81BVYUPuPhWYvckzfgVXmS8DIIWoFqPgGX7ixQ
6GD2IS7GLZgIMgMyuKwKYreGJx7ORHYwbSTEqlf8zgo/e7Y86DapqX94TGm24MQs
XK2YTU4BupO7hc7SBurspYsEm6Q3ki8X67PkU76AxdaMKAWzo2Qp6atr80q2ptaq
aaJumQ5sFI4FykIi4zKQf79gct98HHBwEU22309siQ9dE+kqSwHjvFgdlH8gF5CH
Ibtl8Im3mLQwBeBs6gA4TcGc/geBLjj1qgKbs6jNDcs9tpHq08qZqIhZ4uSe4kzh
3C3xG7blncOGcHjejiNsr3tXcuS8iofvWnVQfgFvKQTdwM9XNh5hhYDFdKqA/IE9
0hDJTlcfr/ckP8H/V2VaSADAfFlwBLlRSHKnTRLXAN0/+c6fVIxKGosBjkyb5Ltr
Gc0Qepzg/qgcqh4pU7lhNCOu9VM6uZo6EbV6MMmyxD6jxh9epIZCCg9abEKwx+BW
dVqjj+SplhZlW01XvIqi9wmo78ko5AzW79qmVEFHAXIZc3AqVLRwzNeCp0qFr+JZ
ns6nkEhmHyYBiq9ppsbFeVTZpDXn0dmtxHIYR8MWTJlgwgASaUQ7lpvPcH1RWPyG
Y9S4RGPWxY1Ww+jq8ZBhl6yoZuRwah2p71n4b+He9xWbC6uEVd2AY7vUp64CdR78
9M9/9wsns6CNI+n+FEPM0oBxKCSTthj3WXOyIhT1cuKhZCxGw5sYJY1YxKZzIU4N
Z4u8hUDhVk7HXC4k2Md2ljznJeyzcHY7ZWGAz9TYRHvSOH02oT25U3AWODo4lX7J
nqq5nPCg4+xaxMuSnfcO/K24vTFh+Fo2rQXEysJ2t3nsbC3uguXFmi9IChO6ZkDf
mTjjDMVxdbfOGS8rFEY67nisVhGnYUx9MJqa6DdFZL44hQkKDgtFgNp8AtQOM0kE
4v0/zyczcgO1K/lTTtRZGSMwjXHAcvDLgnAjXMz3STsc6476OuDDe2uldATC1iZW
fYqSenSOd4jBuCMg7LEJe+BMl1SEvpnFCbN21hQRzO2gcNjDuNfiHpCEdP4YQMt/
ZDT3bQD+Qzebu05Ho4lQUKDV9ZhXAlGpe1yFgqUiWn1Dex1L0K+JE6idfE6RtQKS
BVmaBiHmwFuZ4QmK+2jnBlb/XewOA493ZqqPSGNIL0OKg+V/HJ5DmUoQ2/+B8vbs
f4XiAssT8dVfRx/LV05eakEI3Bai161m5lAzPRgCso/6LTn8L4vjopyFmhR1xlXp
vqHM2V2Jul0hVOCRTy32TStu7JtMZJvIeR0r+U6oOuLT3TlkM5qsS/KwrFdEaB4P
8d3LBweiDTJhJChmzJlEIrPPe7Ma8Xr3COJJy3eTz9Hi7mgQBdHHDywKzpIjXjxk
sHFEkp+pQS2btQn1a69JUZjjnMbGweK4+v8MJWrAxmhgMG+aWGsJn/fr6KsNc2PT
HywmUl3waZHrXnUWYpNYUE+XT/DsuKoJKDinRNyCTikpCg2EhrnIXnYThfDm81VS
1oxExmwYxc+WmmSgEw4Yr+BjE+I2Z3o5807lRU8eH5QHpWN3QNoiVkwUvkwJWGah
ZZ+wD2yRGBIsFTJh2TA4vp6r/icpEM15Ulb6ewZK8MzYTSnb94Q5NDnejOm5sFeG
00ZoojUQEWPRNLaKvELbrCit+CxIFiAeEln1Nga1lGO6dsiaSVLOm7C+UurvhAq5
oaegQ31ptqivtOMryItjY06wHOWdE65nPFi6FHdVCc7Ji85LlGl3Z+PVFK17IKJ7
WV4vJlavY7UjsRup5rZLYy/NwlXOe3SlSrmy5+phEHFyLWTkYWQSn/d4Xb+RCbZs
pYIWu1pXA3aaydYrZ5QnyOWCaJ+f+xb25aqjmWdwfTUlKLOqWHswqRhSd54E12sY
u6gAVLxFNQ9iNPITq/f7WfS7C/w/hTf9VYCKcnQcBWJFwBOTt1zMVlYPU67TWE5u
gcK5f9BLXpbLh9InURFp7VwyQYM7tLZfwkHK20YKkACWLApbT455KTERYYJ30n9Z
tP2elxYwIwApbd/z3hnda8oBnbG2FHNJ6PjRPR3Ub8AhVEISisvMuAiJ1gdsbM0Q
KivRGqxNWolMFM8en5w4j4kvha0fqOyJbeMaby+3S1EE5vBZwPUnQxebYIPfMwGf
TLbQOYLoio9WHXrKy/jM9KxMDzzf/R9s1tMwh0VvLE/y/5VjzTzCiUCM7cBHtmjI
SqQFvViTpQtzzXPNHHRAEflMTU2RkFzKWTD78zBerFYIg45SaTbvgNsO9PmRGpRE
S4vF+4hC6/FoQg+AmtB0sBo/mhmF8VwZEpYXWgu9rBxWVACveFmIQJHNoouVgPgn
F/VMh6aoGHqqCKdESWZqeCW2ZKRMrX/0A2q6kvwqgjR6zZQFB93hY/1jGYY6BYg1
ZGDpwzuuM3e7AzIhabbeM6u9o7vKcDvAI+FVHANhL5CUaWw6uxsVahbT+qKCKnGc
c7Pyoqg2QvPsfjzeCU853aC5HpGy1pckQPnbcT1Ga1uNpZOhJENoqLm45UqBK3Ep
J6SLeXi9XdQo1uFy617b1qYNo4MCTFdlINdixhIHLdwX3wPMq1viYTDu6Txlhx3P
mLa0ISwMysiEi4xogRxTvmXXhJl47NQxFDh899ptjVNXmp+zeDIdf0m0wwQFqByb
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dwg83wnHAkXtnDdRBh70kCyZu0IgZuw5bbUgR1TAYu22aAVvte8VVB71pbBsYlc1
Mz1A5J2xDxUF/P8hiMWvJHqA3ldss2xPwwU3irhbsABPrFxmPUmpDrf6lw/F2BV1
NGszqvtP2DYGro+vcGotmdQyFdS5HR7Nie1GUPjoOfgwOOw7bd0+JeHY7jwq/VYM
71y70KKQGaMKGTUhKyx0aYKBbELJ9aUfMpaoLu3oNiND5n2vb1umVYtN/iITjnHu
gI6F0R/iRkb50cnUvmMGyrDXCDlocmV+G2fEmUygLjzXw9Cy+jML6Wyug8v1rE5j
yh/1Ys1KW3XP7p/o4TvrUQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6656 )
`pragma protect data_block
TiKQ3Brx86R8WgBVQbR8Nd9RNIo+wCDlJ4q8283m1fkfWcvQqTUyXK+LppVXMpN/
b+egLXWxksgxbhNQpnm4cz5jec0DSOrH/B4eTZpqCfeLMQgK6KiTvcurjKqUqRWT
uFPuK6PC3c7dDiJc4RPnjnwRkC59DrYLHAQ+C8ez6aFmkyU33k8Vbk4xQ5VmRTRS
iP9jryY/V92Ej9MWYf2pE3mS3AXsKn7LkGWcgZVlpPu2cz5wBs+fbvhglOKMnNft
KdNAlD+ZVj0wOLBSsADQGfohcwBi5EgpijoXwBmbfdxfoofeekANeTqSJWfgryWM
EDLoa6lvvtwjDNMTEN7yRkLCMjNZz2QKEipEFxEpNZFxO0u0E+ZNA8diZ9NaQ9K9
07JvZCpABJEfm9UTzEHVXO4sJgmHaOMl0eSWAyMnDiAkuFPE/aXhE2BLbjY3JUze
GfkI3njxYFrijycqIM9Vb7wRABSxcpaYn3xqAl9ZeX25vs9aW8cPlrXdPe+Kylo4
rTOYjmTL4yfnO8xdW+VD9choJ+XsihPjwhnQXXwNfXKpuPJ7uEXZttDO4204Ukv9
jj/KdxTMHJE6y3POqfOnZLQdAwj7rtWuRr+9gxaXz9pvle0Z6Xa0fJiDbqqxUBaq
5ZV2SZdUjR4p93SQlkm34n/sBudpOHxY8puFKAh0hffUwgkvn0oSXfPyQvzI5Ccn
I9nqS4iHAD3oznBe/iZ1L7OaHr2dBL71kIb9isVLii+PZON120dzctCZmoFr6LAp
iZSQxyGanh1iTBzZvYXfRibfMOgoBZ1NM8n5srH1kqbOaehfTmaCioy6y5YmTQcq
fj5pwEcgOMjC3Dg+rRbqmo+oZ8ek7m8UHNEqPODZDGueKcAWQx9Ecqi1IhtvyBhR
YvySfA84ihYBQnpDzSKQ6iP+H/u1UHbXavVVcbcmb5el5oVg/1LnzAmDc0ht1m/R
sym0CsU5MgIyPsagODNntOoftrXBdajaOLP3gFy+3TRShUJ2MCLH1qkdBy83KjE6
oBDfTvuAdfHdFBhAgVdEsjbhmG7pcDg91Xx0a/QlbZaM+rNiMONOF01XvvlIPddU
2ZHc6Ngv1aaB8QMA55jXGK2cFSCNxyfiQZKZFNt3TFxgn5DcaKA9oOhOMZJRTnRH
KR2Ol4DsJ96PyFiNWWgAE/j6wXAXtMoawxyumGFqyikP96nq0lkUX+oVxlRDqrMg
gK1RueJvgeXNyWbwUq/2gefvqqiDtTrgertInaCKV6m+tu31LTKwGYtdI+H4KKWt
xT+i6O8rrU2z6+Q3XddWIEpQVvmLKUidRp4bEJe34ZohUDWjIOTeQViL4IAfmbTN
GpjUCoGElK9tA7u1lNzFJbXD+ThkIfA6teX10vIinyg6eQW1PTs6TEYoB1nwk8Oq
GwzhezaX2bcgM3HpRpGJAm2chq3GtysP/a0ewmYvBvSQDEc6UTUg+l/06hXffPPx
QVh57HWM6CNdrUI9yY8rQ2VRZ+JVAvUUmuslhd0F09rHmX1mMeYxMeIlw8sJB5Wn
1F4h0BZIhzO8ag99Hv3xHbmH+qTi5FZ4ENyrhRdRbn0VOBUj7vFDfn5OQS2pgEj7
DSIJcP/IeZ09mrCZWrb847Hp3YhJ+fYFEhC1laRqk6DzU92jYgyFc14GLTqCxAsB
+Ms8e3JY0OatbGDdhFdOeYfUBjt9IBeRdlkFT8Yt9HBl08b5I79rsvwvPQYv7vvk
/6twFGCrKdbcPFS8VOrde7ea5fyIWRhYEnGbyUJfv/MQzqNgLhPflCuCgN9gv8Hf
4RxxSgziwUw/N5gN0amJLMOlwX/cJjbl/hu+CIEfC4HZPNzE50FM5PHtwQyO94q3
dL8UpU92qBwIwy5yb4apDotdtU95CRiSv3swpmqnnkdnxuCM/rSM7Y5LGoHVZm9R
iTJ6t9SgiOC/27HjCD5Trx/tX9pVC3d4zL7rEUXVwr6KIXPm73iRBjgAh7o+mmht
YoSVtnRKMF+yY77kqv1w4/l7Mv/40C93UNnuTR+MaolpWhtTRCoIIlhMGeRh99+V
YmveJB38OaW+Csenem1uJmTngTgpLfK9bPWbY6SOJMYz5nEvNSHzd4fnS6bAULBd
7tmVl1sQPic+hgNe3KKUssjQ6GwFwEbaBkE+CsAOjw8toIssTaYFdvzTvbtj+rIm
yE+mWpzV/bAg6PesLTwXUkeByfkllrctCzETM1VsYdy+iIB4E/yhaRjyqcgtgEs0
fNDDwbHC+eRrj56p0v0zsFuWIvVuX+dkbraIJ3xItSUyvGzrF0y4eFYB2qyFXtVo
6+/L4VbH8Xho1RriId8GDPx3uLprJrvWEdTW3q28IbqQIL67wYkDoBH1wbGjJ7lC
hX1/hnjcObo1Tq/aCgByBeOGPby5NHKBonoYIs8nTX43nbiP1b/BBEP3LCn5KJYA
3HVV9M7OhHO9um1wAvVCpe72JJ+jhzx/LUVtJhw91fZIBDT+BcdY2mEKi6NqK12L
XvZr4aw0nIWIXI2uBn7pfYG3RoEDaqC6Vwmcfp2Iu+irB428+Hc4tbEk9Iz+E58z
DJh5Mp89yZ4xrj9sAEjPPUyT8Nui9E7ANCLf1PVvvlSlCPSwLRQmcT+ov8c5ed03
et9ouMUZN3drzz+Fgh4PPzqzpjXLkWLlwDUFc6ePZlZHaZcoF/oRCZ+88JP2QTFe
AA3rz2bwU1pNfMXN0teA6tmgSIjVxteuQiuHbCLvEbG73upS/abJPhNbH8c/ORF8
cnT+A+Fj4I4q8Vsq12osceovrLdKuIz8r5VHfHonTOZmPTAkzLtQHGQ/5wVb0GnC
lCnuglj0YLciCVgYLLluuMB439O3KcuxilO8T8NLsZZEk+VZij+6XyjPtdfaEtnc
vkp0G8CMWHSrTw+BB06q80f7BJjrK1jnfKh3+4ubjqu/w7yHU2TxcuXj0RdWx3BI
F9y67etPPnGoZFn8L6pQhM9bFx37UxmjxTYDb2tjn5kPmADBTzM/eWNg3faqRPNV
cu0dmKILQ9O+6Wiyd2cu1mpxZ5tKSia7px+nu8uYSfezK79sM5E+oTU4L7lOppP9
5l2wRDr1gwOxXfFVIpbuqfdEm5nLUJAn94uYutmQUVl5uQf1x640fgs7RqwdCeyZ
84D2vK/iLmXHWGuovB+CRhsfezouumGhFMyF69rF5XLSzAhGp3Ux5AiUCQw/1+tI
gaVOfKySJQnwWo+SmMwza+kVD0mdDnStQtgzxjO6bdfjR0RB9fwn4mHEPiDdEFIa
ZbzvASMhot0YnspMSBZy+VO6xHJErstIOkhhe6EvmMCqMv55yVWgIV85+YAXD/92
Bt8Vp809Ls3XeisCXXt37TO880iCzP+hWEmlzKDx7UHwQe/yccnGVPLHT87gbkUy
RhKBuG4/h52ki1A2LiPY1ZaTxXBd6e6ZQ57CBeztvcCxJTKykUB+IyUEmvVZ4zxs
IjfIAuO9dXcMSI7l0qgonSEt7J24xbA0tSWee4HSaJ/UK3M+rl0hHS5UVlA4xryc
30dbdpsf+uuy34y4SWTEH1vvcSzYioUtRT82EkPjqTcDutd9DejZUPBykIP96tn8
guGK7+l6iDMYb0RlbUUc/Ylv85o5Z4G8tUlJqDlQm7FDJqj5vLVtBy5TsZsVbwIA
UdDBJBviGoD3O4mHdcrkdDkpi5pqLuG3avUjw64rAF86plaIrSewyMfmCvz3jwiy
vYjPfllZ99BYi/BzDrsTgNs+TyHSgWUTlE0VWBmjGPgvvBrwgGKA8cTL2cY/ht92
fl+tsoiwPdde5OAW5SN4zwTqhdw6EV4EF4AyX03DbL2S5J7AOD1cSSmEXY1FnR4r
5upk9TbxJHkJUiAC5vkJFqdJ3ALMR84dSP8wx2AlgxAW98wX4CHYFJH7/QDhkF+2
EeXdS3QSD/gQ+aJlDd86yhxQZF2Hn8BzldR/ZoPNOYlRzv3K7dtd70CuT504zoA+
XA3kYlbuKlF5HHIo+/fF41tMZ4nnzYlKME8BdsDr1lbha//13LAqx8Wg4pFnT3yx
BuNyxuAWF7F82vZ03C/lCALnhYLulyTzvNBPVs84S+aMK6T5Irbc3nImt1l9yjca
EN9pFmpeHztcAEBA81i4QViq8AIrbf7XW3zCzSNor7+twa5/31cIOfbxE4P0X6Qd
WFjg/OihrIprHjUX5R1SeRP9E1wlFdYLA5JEnbWEnZvCiCpSdCZCqXfsCNwABlOH
MUpWZR1Uf6QY5InvZ1LovcT6nUMxLu3ZUUjh/6yiLQcPWUzI8pmI2NDI3KqPZd8n
RSclhWtorI33Qx59tJI1p4D7VMum6J5oTtk04H3AkbrCfhLwHWJBj6DjgUiyvyCr
d+am6737MO9BbHyICIRIQytJh3ppeH4KJxIaNvxvzXS95RVZyKLUM6EaUrTPauZK
R1OZXV0TMttgIHOU68kN69jaUM7lkGiBzTisJxOFoW1vdEMVUIm5YUNvN8wdPh8+
IU/R+Vop/v5s8qXaGPtoKXxjdtGsT9fq+e/4/caLq23B/AqKWZ+HxjjwtbSIOuKL
Ohi8WyqVDBQNuxO6/2k6r5xiMddzw9zWjwEDIc0sBbn9apjQFLkgrHoD9VlyNNYw
UbGMjOKsH/Q143JYEzA1p92y43vzQ97kaVZ4o2fqsdW7iM3P2muTb5iq0yFHwYhD
n/oEHUe7vp4tSsMWT8qr9OMrkzoJ6aF+ZooPd1Z0pR5wjD6bLAfueUNV04YJDOOM
+0J/YMaPk1EimDFrx2I3UrjFoqDrOMqT6b+QYF3QKzpD7q+ZAdlLXSU+CArdx8rc
xlkjhzkQDi1+WzBrCCVHQOj6SQP9OUFV6E4xGovMA02wwk7nyVeLYg6mhp8DZz42
mY89aYIiIdDRR5JPnHWLnW9xelt3DdigTXZ5bCs0OAijTpK02nLApa6vD3OyDW5d
n/bn/mJ+wsdZjtjBKHFWUohQYeikPoLFAsa6Gk89fNYhx9jBR8MzdhPW2wlf7I4F
47/mt3EaeinIQcP/VI5PZpNM6m0yNmHhIVOPlYbAD6SGa09tLriu/RRoznFQYRkT
55CzXWWYeDo+oX31ara0sX+aLzLFLoqU1wo/4yIxpvuJ+SyAGHvxGKW11TWaY9jX
oI8WMI+oCAoxDGpcjY0gkQXEVLQAgeqRd27N+l80BlJfzIKWx/kiMHKx5GFoo3z7
WjtRca7dWJwI1Spg4+RulTlXrV2E4Cx9qnJpPmHud49uV5rY70Z2Q8scnspS9A+6
BZS86t96EWn/EPUxUCy3BGjxf0lAVCowa+2l1GrLO/3K2yiweifn1fSi/DRjUhh4
/wENTntZ+DRWI1sUhGKWswsK4E55PQys0Y/UTttKmiw+/cBhag6znLxMa+xBDmVG
i91JGvjT3NPe0ECmNLqZBd7QrcbibgnsAMn8BeChleC2WhBtDFxxw0plEFnb+HVC
5tG+kVZQMH8jnBGLVI3qaiBqN2a3GuhyNLinZpqhZF15JDfVW4vGJiJlyrrOUpki
1pEyUCTOyKYgy57vpY0vV07fyq7GBQ+vm6xEC6GNZA0YpTdjQJ4vxIN3ZpVcOEnP
YR+RHzTrIMEZjBP6peUGstJeEQK9K+7KAib6C9GRrppl2bnBVlmCTE0Zpf2g7KVh
+5vqPrkWkVl6Rklun2aCJYf3yMeMrgl0GYkVi3Oep/v83fzMDkAg+KIAuxjqvlu6
/+5vHpXPgyzte2Iy0j5IlsKdcAtsXZ2Ill6MXsJ5JaL+p7xi5eAn+jkoIG+ZLCOy
D7D9nJVTe38k+GE9pY7D3tJJIlV4gp4hySwnGC/J6Ps1lBZ6Z5py1tPgnxyGyl4K
UDOVbW1ImVghqCtFDKXIqAQ4Sbv2lDIWDs1ZDLfL56dRNgdDfKNzK2GRvclL02XO
fqVH789pmHK0gKck6K13QFqpBjKMP7zFDMVLR2pMAomvQDwRvcMybJD9fjYQ2OYK
w7h7nVndOgz/F508hKYSqTxPQRFlYFt59d0MO9I96lzXbgxC6In7bAviFNZq/Kai
ccQxMruNYOFBrPrBzCvkrAyQ9/Vl2Xl19tt/RBeMdBnhlXwMpX4MBTf4O6QE4/jv
/7SSl4QWvzgnC5NRcFteWsw9kiBPVuWXsoVDWk7IHBJXtrLlsRFfwy1tq7iLF7Qd
Wnaak9SQHSbHOR9V75Fy2GYpVEJlbiXULD3aCcm6SP8jq173Qu97Jd0WuOmzj8Xq
ArzlCLickdYVdRntvEsGp2QKawCb/BNEdkPZZIlkN5/SQY+GqxxNWKfoql59ztL+
0oaJmnAdBPd1noIOdxqTx1tq6IRoGy2FEUCkGb/wpyz6O4TUk2M4yRkUCycBj2lU
YK1hevh5RF6EviSWoIW6ntdsKFQ+Z3wwR6ynKqyzCyawW64vDb8K0YrvsRK3cQ3R
Tk0LIcs94/UuuHlRVoQIsoVxqTQHpaXMtp7HfIrYmfZVWa4JJwFejIN4M8QV/4FS
IJuOtYUlYOs0WfrFfFsoDQUijdX94jzWosUSj3/gxpZyyAviqF1P5iw17M62bVE/
EX9m1151w1q5k78xMQ/kW1Wt1esA+XbkLvNCXApwP1zOYVI6soI18L1mB6OFKM3y
naRs5gT5RAE10j2+zzcUETIJAvKUFfxRbcgcsbrB68y8wRDuUbTwwK1JFwrp1NrE
6jqi2C6rgOEWLEmlyQsgKR2G6iHgxhLg8Kq+7rkyReZe2mmKH9UijdhHV8sD4ZCz
zXvbpIKNsg6iICmxO8NqCwXoJ4GIjHjtJeibcbMIlrk+AkhfPsTsjSEMVI5ZwNL5
tUzXJhUizb0EeVLPair9HAs8r47zx/AukqdA6x35xKtyU3mMV5+AxpiTNypx97xq
1XZOSSaiDzqDQIJC0xAhvKeT22p8WQUPiDcA+xizOzdahGvOdOXMjPcbfRXWGw60
4b/BEzqPtMIXYTK7csWa7u5MyCi4R3D5a+9MBJu9mjnzbqNPRsWqW78Iry28cGuX
DRhi5e1s4h/1KR2/9m40wFgfhEyy+RdOzHJG90gj3jt6r6VpuHjwyg3wJimuoQPK
ISPyqx3H1uXl296t6k9AkjTJvp8AjXjjFZdhEPPltYfbwUc2GztmsyW37W2scd45
92PDfgpWTti5cJhe+K8D9iplHkf7HeV2+tLLW3AvFjbFZ/XqbHXOmDHUMNIntIrw
7C4imszARcLdULDv0FBw3rtg/dcGnwpi6gG6cHpgY1Wb9KtVIuKMmEgIaQ3Ka/BO
UWSLHXIBWOS5GhESbXodDh4YURmLDndQB4aX60hvsO7EoJ8xxBqKJeWXQR2NLaGV
wYQV9eEcyX3p3iDbfQ51cpEwGSIDX5y9I6G8rFa9a2JZL7/vRJ2Q+wnEtdd1PjZt
ZbM2RiCha80WD13WvmIMHsRD98XaobHl5O/v/EAWqJ4mc/zKNRUdgP5WzMvKoHU0
ucFjRqTJYvFr7lE5gbVE/oKc68GMcoV2chf+es8LN8A6+b7OHiWlbd+shRZnRnGY
AxGc/k/pDV88h1MyiDGAU6w42ye+DZ9vmbyXKR7POdz4PpCCwtFcqCwXXNv92xRF
ZVzdt7LgC41VsGSCLslfOhot0BUpWyV6phqcOcV0O4ZHbn6OpAPaBA9qSrFZBrEx
PFjkQOZU8TAL9xrNj/I0BN2bP1GVwoSY/k1zaUsAF6k1IQMLrOcNZyRlmoUwjE6P
mpfYR5rY9/gKTTdztqDLGj9/f5qffoogI+E+mZn/y9keHJJgr3cdXaxdN33KW5mX
BB27HP4DRQpRIxzxbMHgd020yZE6XUcLSFCM7XDUC1uruaNC+0omBHJs4q3HxdAj
mNIvatwceg4HX7NWA8+AW5eQO4+Ycy5YOLXzGHxFj04nYHuR27g8JSKzLcArAI5A
lM1V169wZB1WE2rq+vV6mUYAIkXceyNQlnI8bAGW9uwwM49BQ+FwWTcqyelnYuC1
HqDW87EhAaX7w4XgbqOQ7vE4pvRDpf/cU7EvJDZEHwRFwpmU0J3wJvkPVMuDWy9R
tjaOEuciTnsYKGrtls+KGgbdwG565s1Rk8vgs0nTGKn/B+Y08wYY1zA6Z9m2qTRs
VhhhBHhGI8NhB1ZxUZgILJ8a9Nxn4jdxRlOYFsh+0J/tvsT35yxOAsz+ixiwDKVG
ZKpEnz4EXcPovExq7+QlXB+cy5SRqKiDH5D9In6ldJUsiNrCr1InqGkQq3PWczgT
P89nz+rV9TJFdBpMMdTfodmLMhotw8NufyqZSN0p+/0puwi4uVcAC7MYP5+7nIyd
KSgeh+d4LvV2NDHp9/LpBulT5dJSLEI1iTLmNGzx/ZDhZrlpZ+bP5yjAFByesCvW
ZLO/Efx2PxBK1OQprXuFKgZZiHsCrgSfTU82CZRNunP40F/rV2684qzzvMOnvHDX
nJ24uzYemd4hXjeOOeHrC87WOJME93iPTxsw7OSb4j0LGDc9gaG2iVzGKgL5ue3z
RzLrTvk657voBoY6fRUQxmn5oYwCXTeRxnrVEK0cVQ519CtcNeVqg1K69TQL+a5E
B56KcLl1We3ECxlDw0/CgKJBmATlao+J3ln5xAz47pBYMlcbpKX6NPldoJSKDf6y
O19e9FMogK/vWDTuRMTes6Sa+VRT/Nolij/mNvyzhKa2lliTq3WQfE5Q1cTiFxT3
3q8HR+bJ1bu0Z8R7JFqsKaRvHaMIEeemNEfNrqOPcu/+Y5SkhcpHBe9Qa4vufQnh
S74UYgt4cVCryzmds+e5V+o53TRdTm7nhvzlYEWHo+drKKvaxQQplyc/z1HCbXKd
ZlqH807OKEqg/o2DJ6CPnbw2tycDL0sHSXn/ZZyoAMRreT8b1712ItjHbMNqRuvP
tI9jjxjdUL2jrBjBnQz+TgydGlW0Fjy6YPDlW39tSOA=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Y2yQnAsTHF5/byk1Qpe/hSmqLfMIriS8c+tuMPX4xSxnr1+MDukPj50rm4prPcY/
zUHFrO8m7VRLXcBr9ij8xttKRUUJ7qvaCPk31zb/aM8pIBqRh+aHRFrt9OLrv3Cn
UaWEumUCwkbOTuZ+VAxsNCk721RXmhtN5vTJSjgvwixRhWhC+5rjy8vyqM/0kzB+
F/X1v6ZZPYdWpnPsoUEo0Jk5mVyc36TcnOQwWQbrmrqSUq5dKQn3QH5zLSoVDIRL
p9laampOaP0crUk+7WHemrJNJMjDFCgvkuBHJmTRVSpgYb4cZ7mwV/HJDhSH18KC
pt4GDJOa+XzJ/I/4GvZbBw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
hBLRZz31Yd8oo8ZXV98aRmlipgoIa2TgQCb/Eu2jEHU3PUcnURj+V88rO8bw0yKk
G3x3jsdhpNbdmd02Xeea/W8GPFa4EokCPz4DlM21DH8Ynv5uPUY5Z/32VWAMSbP/
vwEnfRyxaDnS/vbSicH6LI/fmrTyQAh7PbgvRW/aKaDtX+cr+mEoADVVYC7A2uFs
bOvG+rKC6swyWLN07uI3vQC0Gpj0XlnICyzzdWhEf8nHiYkxHVE6IrmK7cPlImj0
V/RHZlkYRRuP5NGjJ9Y0cafg8HTfBEUEk0xP4XIvLIamFIe9elrNUlpy3o8HyGc1
+EMg94DDTmusLCO7qd6kkL9eU+8LHG8+ZX4o3GxT56Xe1j7Ss5Ygw2B/AqkEQHf2
iqz63cg5yaV+qlJvscHna/sg5VAxpTmKC5/d7a0CqcDuZ4wlH1Flyuc8ke0jPxSr
mpCgzb39ShZz6/Rq2jfL5wCPM0PMSdFoHzWtVBlZ5Zu341Ijwyt5COluEcaeGzWr
8xJHI+2uvQER+FQLKEuUJJhKhnhVZoB//mhhbVzGBS94eoHwVnPDmmj18gd8UZ+J
yHTox4XwQexq21w68phusvwsGUQ6+V7r+dtJb9Tmo2hhMHBqDeJrl+ubMz5YxQ27
zmQwtwlJ0j4C4vmKxvOA9H7Yzw+mEZfFLFassfhCFytfZtjRBW1OmDG8c+Q+4Nbq
NZNmf6yED1WNtgxGoZnu4LA1mlPKkwXOrWJfarQgPFzOzxW/YXVsk3s7CsMVZI0p
RnLhE9fjmjAuH+yBYjnnbB8/c39y4psWR6pNqbVEuc807CWWWg758iZVTvHMuiQL
okcVN0+SqOpdbl1m31BAq0KMC5wARtZ+CteckbnaEQfLPF2uznx8Q0cDDFJ+QwS9
Z2ej+sixxJtrB5rfhbXD148vL64W0ZgiMdmOAMsr1ba/AmnMIrzsIdYuP+vA/lwK
WkkNZegiw8udZIVD8ELZiJStkrsv1ZhUfrJnlr3/W7iIAQCQYtv54AW+fI8THiH5
VFzzXps1g7xFr/py+Ip9YxM47VsslNkifpP923LtLXZ7XEMQ7KcXIqy8Ekcj+G1/
DsKOiplLcyUGtH5UPFcDsfF80PqMl37rv+nwjuApEPxn2YRlslSYbXwEMZHkipVy
xSMApt+7NW/JBO5CN+js/hYWVgRts2E9EGkS9VRZTu2VBm6Kuz2oO4jDtfSXuCql
zo4fHhNsmpqo93m+SMYjWTAHjcycOhqWO7C0hJlEgFDD5z1XpXbrdPvJtoG4sk+S
vY6V5EUZRaRmWQOFIRnJHkHAMJaVzy8sPqFpUnuXLbISAMTV4vPG9qlt/kmkWyg+
o1D+W6PnJnKbgTXE55CZgfq6UYNYNDAu+gU93jtgcNE1dudRrpmeVXk4i8UEx+xN
pExg1CKdwUIHOOwTIc3fWHfwga5/rIhH255QR2F+Zka/xgmqbU4qRgkySZjlpLIL
6kv90T5XPTFriEQb+dm7SMGgzd0SWOCj6zKucqsF8+hpqsjMCKOWhY8CRPOzZqe7
bZgWUQ2OX55cVIWlV2goZLhiSE3Ct0dGKRPDk+DMC22Ziqj/LPb7/iHynPqBoGh0
/ECw5XU25TPOaUGLJrkoGZX5rZYEjeZ1s0+OZLoI+IEOxxgAnl9kLhy/menRSTx/
UTzHHUQp79kmg+D7UHuvtuT0yzWyNxz+XhYemsxqgEEFnq5MwFt3Ru8o26aFMA/j
4Pj6zp7Y36I9qy2o0lVlx8/6tNcOJ0Svr+nkSWhO4AhOHJ4uMbNsRmHRWyTw2mJA
hm91IXosCX2txxebuPIhTWcFooYue80kNRqQwFqysKFGM6VxprGOH9wJ654QvDpj
SV4b1zVkpMWIk75SDgQ4JcilUatTXH7LjbPtSyhAFUVGL8v4m/EzaT1wJ8v/6tUF
c/wtuld9j3ln4jQnTD9BADDSicctOVhtCvX177JrUY/2Bah4lYwvEIr7j4IFC76s
AX/g5siYODd0xpaxaaQDCPbkcQHSPaQWp8+vMAMq+rFp69wY5lgp9NsbFwep7P0F
j9bd/AtBXRZODsufq+0HrAxzb4IPwCfB/Gul5XKoyRHuNj6n1X1Tg3w5qv8Iez8a
hNFAamTSbZfGG11riDAgBCTLBxf9F0jk3j6vbD8HHed28VaTjpTviOzfVkI6FPj7
88QjBZeNNszRmDTSdaXVU0mpOJKjTIHJbCT9TjvcVRbbJqqh2Vl6Fj3HsWpaJX+f
gaH9TUqqwEks8vQlv6KA227G8MZpzoEz/lVsAHscPnKrA6XeXAGn5t1cmVg4T4d8
8ubl5eHSKubnsnBEGBDPNGjwGnZ/WsDPVcTH3XP2aJS2EEjpwwxZuiVVA0Yr1fMv
qz26WBwb1iWMjyXK41Ofr++skvwND+gC7wPyQ4PDxotMQddbI8AjbAPsgICKIocM
4wPmHt2qFgHy+h0v7Uh1Ju8PmaPncQeKFG5IKINL6jJ2/zwMOqpBiF6ZLQqfM4Hz
o5GyWoZCcRZwf6NmWWRgMZi+Sxar/8bZMT7bFTrZDyKRLKzJVb/JmjZWg1hOXv+2
5UFTvKR7UqARfeEl57IaxpNZBBiFiGJ7Jj45lSQWR7zZNWb2oOLGLLUv5lgen5zC
3ERho1Fd7X0rcDP3slWi540G4gVwLh6h0gpsEtog8TdMEs2YQOqp1e/stGsGvSyI
FG/CP3ZtKK2UTd7RGpDTQVnkshNNZc24fGWwQFwBHcz9O8Yn0Qc00+PyJz1HI7ws
QJDHBMKoY3VHsZzNH8VoQCZaVyB9A9Eq9ldc8vSSNGFd75QcX2tjXhhS6wvaQKXI
L4g+jhsfEdxJ3S73BQShNa45Q++cgemhpzBGVyKMwcr1miAM94Ch5RgJEMT3eRa8
6NtpYyZXjPfPxw+tZyptOhIbnlZeS/mVuy1qr4rPNLL0rdsh260+56DNG78DHfqx
HQNiyM6Q5DK3yuk14u6RC7gLVmtFmWzIWeB2BvHdGbwnDBZ+NQaX0NuTF3kuqUTi
waw1AT9UOIPFmGNiRMDdb/vLk70f4WaWfRhlcNzONqZSDzmM9Z5QNevIG1ihHAt1
ZuyRCs/u4aBa56fbvYO+NK4/+cl1UgwsdT27V7+vdw8cHvERMdwRBPZEjFiDHjWQ
Xji19caZGEzlQGbJM6oSVGOFgamvCo0ATKGBvlATYWaMMZNVBHLYO3EIcHEHxLzk
sq5BEMhSL0YLCAPQ2EeAHnhrDFuOERdR4ESrr1v6DdKIfp07CYWJjcMCmmIL186W
Z1V1XaTcifI4a+t8nP0EUaMwF/uL59Obqpjd6DXrMeCXP0q1pOUUpZnSQGFReIAN
MdD2rPTaZOupDTIVbaSuduKGdtVXvlDc9HCYnDoQrPvAkk0ks+cwWuZk4p4ec4Mz
8hzPFmYPYCtFlUgDaVoEqJ/GFbPOSthr6qKMG3wHAATGixD6jLBCKSlTQchttpkk
rT/WQKIAq73ojViiqhLkAtdUwLFWPAyJzFQiwOUeI1AgmBT3Tgosg2eGG5lnARUi
5VurbmWEdcult2CI/ZRA7tLs2M6WrwqIzYh+vXKHGHyC84fKQirAwe6+XZfuSzmJ
j1GBoT/npxonJ/XzHJmZ8anWlzbtellcRKZeBlTR7FA8e8dHOXUefQXjgY6InCmA
4l1UjaLSAcTF3LWlOZzzhQKh0GzwZ2IIMyXBtrO4smjby8zHgrEQzIPo/5AHZesB
Mnm9iWLuZnE2wW11zr9CwcauU59H/9aLBXwsBn8duNMk0eBHaxWoAze6fGb8D1wj
3eB07o0zWcawmfCCGOpk+P7Z8cSFROH89SifrGT6FnhjNUHvM9sPV+Tw/SK/tin9
61dvtORqaRrc6oqE7YOUhPhfV+5f0fSho1CaS5xIzOYswKhqteZAcBDAmiI5gVQT
bA2Pf2tOC+tUVO8mfNQKwnFawwR3J/4E7/gtjmUIxkemvhETlP2TnRv6Aa2onOzx
KxC/AfxJFmtE7K0aFTbrkj2/KM2Or20QJMEn3WhAqeexDia8eZ2sFBjxmBGtsr1X
V8FAZXkr4qEgU6s7ePHGini0REdXyLl8txpLCNYd9AvI/d2WkDKn/TMSi+hWkQUm
PcLoVur7gt9XZn/88gJnHPvJUphke0oZRh3DXAVQBWNFBK0T3R6RjHCT77epPCT9
JYTJewGsetkIdRuNxSHZU6tgk7sjLLzoQcaou3nu0rKFKnMZ5BY5QaSehUs2qN9D
S/T+LqZf9QhtnU7AZ+oZ9xOwmo6fGm61zH80o6WMJUAswC6kSe62JqlqOq3UtiS7
/n8pcyT9LEmff7461zC2XF/8UfcAoLWV5wZT3VVKhXmhYHtUUKrJ+StejvooDe/9
2Kq4ZjhH06rOfjRcXovGLLD7WmQyySraD/brlzJUpoup/nFyZBZCSl5G+19X/fH/
CPIABAEtUXrNHWDQE9uc4jZwbDSQW+11qNZb6+tvDtKEAv9d+uXzl4n4zNC+u0aP
acaKOMok8vTwYTNwW3zzPMCOwHRuRufj402SKupx9b2IcgIeq7T+JPI6uSh0UDdX
QFR/e8afanZ+67lUH1A1in6fazD+f8fWUZ62Rt11DQj8F73h3BtIpNx7bNXXwPHD
15vzUoqc/XDBwLuQSTaG8sqsVIBDuitsoRJ7FeCE55OU6TMJXUb2aVxJSBFOFh3D
A20K8wINTn4c9rz1+Dxaa01F8VsRhZwvwcGE/J+QDzdgdOUVWMs/nV7r0ANyU8Tx
BuZ/DWZ+CRyEQC10gO3My7qoJyeJxGdyYXIT/of7mJRel9ytFrs0v4a8qPk1Hcu0
V1lynoMH9OdG0hzTmBQcbSh277Jd2zIqTWK2o/qbvuESX9fPG64pPlSv4qmIKSqm
ScgnlyNtJTIN+Hc3+nGYryM+FGRZdCqOFuZ//+DStvX2/g5+FPWwbasehGpopEcm
cKcizsFwTSn4ClIboKMcUFBLtq2ihEGGijlzPbYdlp7ktKobQzGU+e06ugr5DdeG
HAiyjz9m8ydEuVHHMQYFAm0oxs8e9Mw0zhwQjCzuGqVm7dPSJY1/BU+h6pDphcRD
fXJHjofxj1n2K2CSZiUQsq08gJajYOXni1mhrODzIhsZME3i2PLhBMstOjqqnKXJ
CHPLOZETRlKoy5JCK9/lJmVxKIbhJtxWN6hUfqDH0SL9WSYVfwZE5RxNmXvxETyv
JQZhU7TtpRax68vzz7jMuNmzSYxjJiWMLPQTTI/rkN3qbKVVwjZNiRrP4sDr+DhW
4hKc8h6KyuQ16kxuqJgJZv/P07/z31YTEIq3OY6kTpX5c3UH1YBnGEQJW9C8b6fZ
RDd0/peOugCzmQxoffMHkIbHvy6EsnOXT/HLH++jK66senAjSxxJtfAO1hpWKwhM
f6eaO14By+SJkmh6WgHna+b2E+NxCjmlMhGJWW14TGsKiQnWZw/e+Y3vmFliy+GN
3B6XhbLO6Wjk3eg2XPQn4sGrz5zYDtT7jVMt8mpqDGIpjnjqP1oLe4yqC0w9xisR
BfERufD/IKRXZLGi6PrJwPZWah0mEAMXGP1H1cIzZxvQDCO/r955iEb5dt0uOj1g
+2FFJEgOcARMpyUFArDwf0JQra6gWnfXcARbr1CzQUsFCY7qy0uTMIArN9QOb3Em
CKJxG6ML+x4SDDJ1LcyfNdyotRRi8cLfunesYIfiAs9KKEArpMslFTaPY1jb1sXi
hbHhsVOH27jwZt1KLvdhqPfxb3opGbgehGP4Ykz+3GSY7WUMa5TNUPonpd7Pkv/B
AD8IxD0tseIuaot5mZYwqyGhrDza4Q8dRpOBvRUKOsFG56E6F4eMdzMl5r7cu1tZ
8+J4T2o6ILmw68LLFIn/uqO5FCYMUToBIQoVrYIgnpJNhJmBnS+tBnPni46+ZvZw
MPnWNPYem3P7kjD3gWVA6AcsQ4q4Z1KU7Y8KU3CcZyCcJyuI4GcF97RAIW9oxyw6
tFDXZZTn6M4cX1jsgYY3rgsHWwlWroNchiR06RNI7IVsPqQJ+Cq3/sdLBqE07RbX
Qj6UqQkzBsUQX3ehew+ghRhjkh52JrgtQjdo6zZBQjbpKDSBTtMRppSEmzuxDEKd
nZydwGzgvRgLfKYyJZlCD0/xioSRD1BUjsFAUT/xIgnjxScEP6MNRxM/2uV2mUaw
knD4yyXARaxlVwj3QHr9n5P1yLHu2DST3b8Sd2aLaL8rKJT4paezQgjqnGN/zhyb
qPxnBwswwSqwBEbDrp+hKC6BGVWHOkaYJxMcGYRV3lOwLgPe4URfAi9nExwQ+dSb
GmtdRLMObU8/53qQVj1uvGVErf4f7+bcWjQVJNoR2490a9i1NyNna7UWln62+pEX
3h8zDp1PBIKb6LCrryzPvSNAwrP7R6HeBtWBNINWx/XB7ONhaul9fcztw6WUIfo+
xp5xRWkbSdNUZJvOwMFK5exuhyKm7ALb+8wGoIFaRoRPFyxlkN83qbAupnWiELGL
e7r+aMqP4c09ZQzmS6m81MjxxgnX3oQqFATAiY0sKHIIGB+W6Y92dcqVj6iNte14
PjzAFFLS7XxEK4wLpZ+CVWtIsbNJgqlOcqvsxo8DdncwyPnHLV1XaD9z7uniFMPB
PUCnsLBz6vxnuUVGY4Dxo3+MJ2RCefklVO/nrLDhEX3kJFltu8VbT/E3yljzobRg
LbAp4JEsmUbhXWDhDYYNvrHBPQWFJivVa1i4gOGjOWGrjXnnCJxchWL7OK5ouafJ
WH+MybxBS7wcjge99TFSprPY/Wx28tonuhjAmgi+5CjQlMlDKBuaCqkP3AjC1R20
NKIWGYkyGOv2yUY6IzHnFR3aYDMtuLn1nxRwPPxm3Nril1JffG3wy+EM0pvt2uUF
+s+e6mZOgQ0Pz7a1VZUFpDB8M1595phTNfvZ/2YslNLKwl30NRFEF2r2/3+AtdZF
qLqpaB+hDvd/jryUHQoubVXEY3kYvQju0nvCgjnltq3JDrNWQ1sraNAhQO44ghfu
KLNLxG9R6XmXK1fbeapwxsCVYcJu8pasbwE3UzocmDWLdw/T+A2JG4es78CfKGH6
gdzPMDhbaNeO1mxIReDbjnIsDgo3ovTqYdnfb0bcQ9ovgbXjW69BGa8OCkNsIV04
3wQpp5vHfoBxpaMN6TN+URB9VeKOC6FLu5UDlrLbbqkewzPw6enHdYbbL7klbvPH
uwLlev53Qb/uJEZE1ciMBvIsGxuELGu36olwn0jkgoBXijoO0fSxhGKUOw7ARcTU
zsAmN+Jc6Gj9T3wAqU1fQhV53crg/FFRB1pfHyq8c53xZQ1VYxhmPYsyOMwWP+iQ
7RdrLlcRgFyMd/yQ0/ex2pIt23PCbMwkSnX2Xy5Q5eNAUnziVfVAptzp59HMFQAN
NqvLUowjC/SAVPL5O+pucc3OUE02wTN/CQe5ko0cKZacGZ8ySDlkGwR4U1+8a7jl
wzSLn/Ej8+bCe+5poGOsDtCCNvOzav2Gzs8p3/z/AR9K+66sFmZih0098ymfOYgR
t3rVS2JxtSIEFRn5HJqMmD2dWpoG8iOV884/Uob6spWDTB7Anh+sy+Sgjsg+88JD
MLJSdFpb1PsNJTkNXa8jz9Ww9GnQ+cEtOToKw/kiyMEugubay1O/+0EgSaAuXDdI
AQT1LlY51gN8/GgpyalHV0WXwUhhUonpNfjk6SQV0F8yFuHX7Fm7jIvR/xeJoe2v
jEtE13ekIVOIjBmL41qdjMiJvA8QsaAVuLMnETHpDQv8lX82D6ItpD6B70FiPXOT
UFgtc+1rofDAHxT6BBSiC6PPb33SmljxEUPLJkOwuRxDa/0EjXg4Y2u520yALljm
hEPcYDiNGcLxbZrIKFfE91gPnzg6pP7aPc6hRuv7qfjcFCLN2Rb3OW1Jzx1tqCwN
271QwRMzpXq8YvxmzD8eWd+0KeF8yLwvDJWB6aYFt0dfTmWB+epWvAi+duedExKs
S0ZJ2Yl6oz+2rnsGyD9g+OT78LgoT8qW+4CsnYEPHO5oBgs/FQYKsm+x8amDGnq4
XEYR9ffxnDWrfcuK202LwA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
KUmNc5PH0DWOLwh161mJHDHyHt/QxvoUoMj34cvZ00aB3jeDogvySRSwiDiEhAKl
z+Dz6p2cHKSpPsqA6MMRpiikgz8/T7G++QzjyPztLGArnZ0Dnk1htFA2qivfmrls
KNAScrJn62HQx5N0sa+g7wmPTv8YG6v7YhDOy+nj/JjjkYiZiQIXBM/XA4e5KN1y
pmwruHXLd6rng8GO/PrD//WL6IPq1brMgGg61J0USInXlkOF/+W9EdxnibkhmAAF
huL1cR72ayB8vr+NT/MWWIQppjgoxC3vVZbVgv9Msgb5cn7vOn0w9qMF7ESBhOG+
iY1kmENqJlKWtBqdcWpMUw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2224 )
`pragma protect data_block
UWpcy3QmUovBXCfrK3wXzhiMxxeQ4PGT1KQiylSxtypoFO1G5+ChFmhcTWcDpnjJ
vrroPZ5OK2TMqGBAT5Wk4sSUJeJsjuLa44Pp0tdb74EO63hTr3ELbMqBMgNLsfzq
6G1FGuCudgWxHBAB/vsXkUjiVVXGC6xSNX6bbyFlGQsOffXZ1E04BLG8OUr7fmqL
XfyB8pvHvd/3OjWsMk4agN+FCXTUSkZlSWjDQYyrLjT90nx8xCqNdbnqfTNebsct
Iuh2RLK8LNdie2cmWCEj5Q5yMByZJ15Dw8aoIqNh5gEHI+Ik8RCpBrUG4e+a8H2I
RT5k8T53MA0jwgDqElp6dNt3tPf2Rc2EkkEpOjGz+rgymOJR8WnxB+jColKhSURx
7VNjruFNcyWzHUnwQ5VfOR6BWV2YkQorXa8yOShCDepbFnKZriyHaM/pDVHVyrxT
tlb9/fCFF5dWjXpfE4sPylnFK62xbkuOeR9FM09Hjlq6Yr89X0qJfDeTTQn5Ct5M
aQhShHyQh9P6fdM0S0mg95KVN6t8MXeBEaQKkixsO4HOrNLEDu4Ld2FaYfqTheO2
/JlLFX5yq3aGDHl8Eh5BO6hsk0qEa0I6pBISI2xyI04bx1JI7MHZ7fARpLDhdG34
cqBRGCNK0OYUhy56DpZ4VQ7tMMh9RtV3X2LXSzmnqE7OKctijv0/fEZYZU3Moxdm
N+IHyIeoMa//lq76m6jBvkb+nUW5jlbZn19R+o3Lg9+N5Sm13+6g5P0htnL4R57b
D/5O0OR3dSe3YSyL5H9hln2WxuXjejoHV7EHoOYK5Lt6iciYHAbLhKRx6LoKnMur
4lgi8LtoumD/GgR8e4cxASMwnXeDv0H7BCiplXr0ZACj88Rul9USDjKXMGmN1uCM
ENaoTGIgRgqw+3ZrTgVI4qO5RM0w10Xe3je4UdkEzjC7oCVnrqKFR7cMUQhtMoB1
t23aOeQmsiTfVpidDtTVq5pM8bu3TN1dKr59KekzHMidY+S3DamfNDXk94L/n9ux
foH0KVx4jVNhuPsE+j8hgrESgof6vPmKamea4h17yDv+UymTJ+kOCwC7CiXTL06J
/u1rVXEPASvuv4HSMJ2haxv9z3odF/vZrgVavAtSNOWbcfc4+U7WRzwGwtBOWU75
lcc5CGdAWOXuC7jCwpoZwIqurUrjuiIZq31bor/Sbvcl+Cf7NrajRmw7Vo0FcKG4
8j6AUJx5V5Exsa5yU/wGEVafPSwm6nKycwn3gNVyFQIIXgBwEBknz0UnOrVKlJ5s
HvjJ4fs7iRdx9RZ99ENc0taEA96wdWKzkPZfq6hFuGzTVvGoHsiFaw2O2s5VrmQj
n4gZSrDBAi1m2/ySf3uGLLVayKdtHZaLXBny+z29m2Q7/wejzxt0k9At9se2iIZA
fcpj/uQUDcemEBbL/+EqCr3u6PjVLUlGTm4fU/sKrjBSTI72fLENlT2JzYzmZX1B
LAKltzrMhzU1m0HZ0UTuaLiuzjC7qYXnI6C+dgDYwrQW7p9r1GUh5gpUEU/Nqlhj
YCrSX3Yxsce780PUvUC1ZtZfWfm6YC2EmZxk8V2ICLVkRYFpMIlgWXD4vn1C7Y1P
MUJIk+scCFxviM+6q3BWyZBBkgOZTdYQ2KHAXW7YqgxHEFXc1I/uavk/+DrGkdPV
mIejqmEIsUo8gFoX13xRqmewNMqnae5Kq15UoOkHbMDbf9Q5U8J8PWC619MT57ui
mLYjsLZbEBpZGMEPHH+cOoBjUPjKGl5g4ff/LxBu2jZmG7OGYcttxYVY3va+n0YT
BncgOyrOZzR/wI54f8NTQiDrOgM/47hUtU3u06shJipKXGjU/Ent4GXxHRzm2j+p
nEQXT6WwUyM8LYSbU+luNFRdT6wEo0Dp+fgmTgeXET+JoHd18JjHStYlqww0syzf
z78e9ecgV2o16wEzlsWVWzxXr+85+U52FcCx1MitOgm0z2WaJVEgWuD6POLon7tq
l1+o+2tbQSN5PIsHVi60HYeIoQPU6Fjwn2nIKMaB8qQV21wLSjlKd0KLSnMoHuqs
kqVh7AVBq/6tRy5zTTtyRB1dbB1Wit9AGZf4VRtveTngABJRs0eigKM5Zdk6Dw9M
7Aa9i4tWDd1udOHPPAIm9LXHvXRV9JJzMpUEnAbuuC1r8zP068yXTkKtDxQ4Bg3x
c/PbkjvoWmvxz0dPTGW3E2RZcRGQ0LxPt0qVTUj+iak4KvyifUdDPbr41UC+zuoF
H6YL+egX3lpT44y8dOrcj4VNCus3qM2aQ0jPmcpucNTFwuENVn9NLtbcI9YKITPX
7fQqkcAJxknF8XsbGDS4HHSoU2vuyjexOPyoeRhIk+bEXn5Er1wWcU4ScCfbaEP0
Nyg6jUEnoZgw4eRdzCEdiayg19EylOAqnKUhl2opumzFa67uVsZXu2+L019oPImQ
X0YKlg7e5AZ+uPps7bRuI2iAiHwM5KnpEIQw82FCs9lAcFFtph2kMqNj+L1mzrQZ
DGrDz43oJJ7lmaE+caedMF3qgNzey0uog3mE55p5cK7DGW7TJZE5+PUgeWLUTYWV
aPcpJO4K5ulQAPhqyS1Zxs0tUeNvGbDHLNG35aPSKGj0vRzOiVZb46EBbX9HTEkZ
LhsJ8yB68T64aYUDAAFX2JCUC/8Fz3VIkg5MSNO+5MP8CARMcfPxeKtVPIsIwg/q
e9IqPbKXuu1Ba58H3JGppZkNbDS8/eL995zn9oSDypDUxW0Xm6MfNgKp34EaD4VM
cCy/9BB31+ydL32FLd5kvKdjoMWXq8kwoKrJrupyExbK+0F1gZKcFy4/7xuWFWta
1F4J2ZwxvI8uImB/ARi7OV5TlC+b+SISSW4BQT9ot/AjJlsVImESfBrSf0fraSGl
uw0hCAFJxd/34OmVUuo4Tuj1Ija1TOqNjCXvPXKWPbL1428WbcEcjCYJYk5uhauD
r2LWtcK1s3E75Jy1tQLFYg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lH2StVFl6WSQk+dle7yrh1lHfXyV3+88FFru+2Hdu3sCk3zQgVLNMlturSFfgZUC
lW9NQoA6sfE7nyluj2MAZaNi+6/kaKIbV9KOpRkhBfVBcODvNfGCoduFXEQ9BGM6
Ad7g9lH0qXXMK59V/9rgtUCqfOn5oUOGFHirfL0F7jUbgiFR9Z5R6LSdn7PvbmTq
gZJVQmjfEHLBAKtivawgGz2yTbIVQxTcHA9AaJLVsKMTjpBcciCPm5o1a6aL2yPc
sPNwJBd8zYBX8ZfRY2IWg6WAyhAVSLEb+e7RDMJEzE1oAvR+khOPrDxqfs+siYtq
hKeS6HpEAHYSVq/WUtauEg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9328 )
`pragma protect data_block
4pDW3Z1QdQmfpJH96rrWv5MEuhZgQHw7l+0dTnUSNMlVhwLM0ewJ41zlgFC+AXOb
VK1gLKSvCyuahU/4oOlLmx4oLlZhXhk11ZaffDzxcbF7L3bibIJKJabKnZUwZmQz
MtflI5TAkWs0mY3Jj88ur28dYx7M1JBLUZli6q97Z2UYKVsUdz9UDgUgjepFluWt
gdRBVDOaUhJKqUvxXEXpFsMjnL4dXGul8pk4Hl0lI4e9eO5nhOf26rSaDW/dRkZx
cuGAG2UYWO/mDmjfaf28OZHCxkya8n+BCzBNvVCCU78TsEgeYP6+JeoElCHr7zOy
d4JdTm3Y2stgbpXDkisN5JACG0cb0yp81fBm8KmIXevS62kPhyzCb0euOO++Ygh7
Q9YVpPwdb3h180q7o/bw/gzAksmNpCWvM2xC8Lmn3IMdXP0LaECMhvE3PxujSae2
ssG48VoG7+NIAilFpOIlldK4rDoZ+MOTMxFvy1fzEk2EZaj2Mdv4kEEZU2voszMx
ZAdlvMoj6q4+4y9VvTT2sJu3sJ1Tz89x6ch2K+/i26Ka7+zxN+AgwlKtE6q/Nj+p
B5dxKTGLUIUKnMZJ3PfbJ9fw6Tt4jYGOy7z36qIFUcBhrLbO+d33InQBWikvet2d
2GkCCdmcu2B2pXmt82akUmuzQPetwqnSsPhgs+5hBGPHi6hitxQuGS+nhp1vbVDa
tKFVo0lRnssEJuPrRhsr3E3yaAxS5AFhNlL6cqiy0/WgKNtHh2pIKJgZ2rU+jFXz
3RKPGLs0Xc8HW3d817uZlbR1YbbhWO+YFDE4x4HWcjGnwsNezqEpytDam+8q1DYs
Co2Gx2hOc4LTeHroltsw/acpFdYpF0su+vvxfNQGY9ENjHimqX/nsoAZif+6VM6C
Epqp4RdQ65KNPxagVht42bmBrzaDoF5hTvmOsRB0UnKtvVdKZgENYVGbTioVuqeL
L+sc5Lw+Ri4uuz6JhpNvWDf5bWJRSHcR2yhk8ht8vw5G4JzS8UrpjOq2fr/3jtbV
I6iz0295mKsvini10u3AYo+ia3vYSg7617D2Uz/ZNHLNKRyPPLrzHW9pj2SovaTr
OyYtADI6n8xUmvwjGS20hJR1L8R2qrvAKDcCOQ+3Sact8a1T19/Bbwo/5+t6Da6f
CeeDtt+4jI56ttWJfGpTMpIn/M6wdsePqp+S7Rp0lVWtyKnijV4SqNZ00wJ19xxJ
UuQoDxgrsRz1OJaQOCC+il5q6ljQhV/+uJt21c23Jxz4+CbLTfCuT2BH8Y3T37Yu
J7xu78PJasYY6n+GiyVsC9oZI6chwyz9BC8msHga4DQSzA2gISdvN5o00I+fng9H
2xSzeEVm/CmHPNrN70l6a/ZxaNy3PqtdvxYlIUv97tXBe3d2ZGaeXpdDy4jffLpo
sSeDGSXH/EfDCTF/ejVZmPWySDGCzbVfMRCbjTw0spjCRvC3YJzZrrSzkgLCu0OC
wbf0hbNI+pUd0wQhO7z20Ngaton4Q3nb067c4EoAnjfPt+fM7jCijong9fCoEkST
BCvMOQfRynRs3y7oM65CK4mvaFcWvNRb1dxdwVbw0e0KCq++OzsEOugLZ4Sd75N5
Op2v7zC0gqpmAwcPn+Fg9j1XAuoH6Wj/oN4Pe+gO7A8uqRp0lQ6WGfBhPOiRY+0G
tbTNpcmKNx5GqWdnYnpOxWbGvSxB+KP9ZFZTYenEgNiLk1dJD78b6xug1GaEeo9m
6paj8pTmlUQMWqYZlW0GD6aYgf0IpWDaktmVSwz6uqJFCF8/WodKzyja6AJHiKm4
AlwlZMPAqMFBTtNHWanMnDTNjfX2Tg8Puba1I1YFv7dLrc4ag9wdHXy9cll1ivXc
kC+pOosGX/prS8zTU4Zsa9qfRBICZoaPmdrDCN4fxYv3h9/+Z4mbOXoJDx2PLOR7
tS5mTDmca89M5lDtrBevJg89RSfCHIMANGPpWQOSdMKzPyXso15EFiPN2vz4GGAt
B20BoFRn1VQfghjslVFK9eDBIqVslStDXYDEybh/sB8MmWlaMkxR/fX7hFLt/CKM
TauqnFWW7yHnwTkl4gQhD7xYtN/UD8iI575gSKn5NHAli27304vZWh3kkefs1ctk
NEYV0fXFmiw54dt2A/aKnp54r8PUchmIOiyVaTRxsqL5uhbxNHzmH9TQtxdCJogq
mAwDR0qzzTklo/JJb7x0IxmxJ1F73LmP7Qttlxqy0PO3fYh1LZtj9K25mloglMfp
5S6kXsZTdDPP6xv2dawlYke1FtHYcUcDGc1mkKstXaJtCHpJZpSs19MTTV/2bCYH
Shqs9YNS+fLolicTzmdBNJeyCqcH4tUarRO6viBjJoPntONAYVxQPEaXabvrMnhU
VIT4zDEsgYOfJsRYVduJsc4J3nbz7azTyA7ETfo32tw3xGvvQwMOMNYRQob1h02i
a7YjtFkMcZZGpZ42n2RQJd5U508XI8BPXbCPK1/gQmet0xCeFEOEEZwOexWYtbn6
HCiksNSjGygjl4i1l327Jt3fMFM4FcwmFVwsvTJgZmqxzILVowBAyrYjcNpol47h
DxdD6ilG7oewHGDq5lEg/qFHNzROeqGosz7GX4nt30K8QYIR/7DK+FrNsOdWsdlm
q7NhNvNEkMQ7+d896uh4Tq4kftdCcLrdzO7XC7+SoCPDcDuesZufAO4WUn8mVMoU
3cMBPPiRDHF1bquiupIUXU5wqOeR5+gCB3lwOOp7AD2xWbJTHDIyc1TidmsxJyQN
uxZTE1goWMhHca6PoXpghkSnxmj8//CKkrWPuv4Zl3o2s9pt3rLUa1fA8AiOkVYx
rJeVfJxZedkkxuIefYefpSwDn+zQvYVxyu6tVCOjr/aMXC4J1mUQ3dl/nHPlDh41
n7jdUm2NzmjX6rA67UH1DrtcCMuc6ZPTObrXhPopJnnigimxu+DS7uOkmDbvEmBl
VsXfnxySt6FgVdZWeDWY8fTYwjSKyJM8k3vPUTH2Ti7nWzuuiLMPWn9w8Ddvz0bc
4zmCxidUi6pS8bVtJtK/Pz9crYLy4E5xhGC9p2rpjd6t+ea1og2AFzt767cKhwKX
luqYhOLrziVeEDDIm/rwjIzOz47yPcSdOcWgoLievF1h+NWmSET9vtOepsZf8TBC
gTz/LB2MzsSJ/EUcShm/PH1NxBgPUtrPe8r23sHDxojkRDGUiH1T9j2tkmpn701y
k4misolMmuJVjF01kzsa5EvhKazfAFy6GSUvMpNesR1ODEuGpfKBOy75cd0vEJyS
3YcI/ZRMbBueTdo1HXLeTYDDMOQvVdGFqpcf15Rz46/+sMxc7hFFkYLl3YKs+XbV
H4b/PPXIMHRUN4K0pxKY8kewL5wjUA/mkuNL5N9KAI8I0N49qQp8HGWi7TJ3c65w
ekfxMyw1QhRn6qE7f5CBI1w5QRIzKUNwQuQirz46WWx7wYiflanz94qEX00+dAbb
tLhGgKQ3fJ1QI7v7U89YYPgMumrIvwM0zsaXOTzNY4urtkHSDd8qLHF75jZyHZGS
jeWDmqEgol5J4qFqTjJs96m9htpgWM6+yBNUPANvlHdS1NfIkKFAAuvpEpV4YTxQ
XvTygzR+ik+NDtxVhi5rEAoZ+vHeqsNtJF0rgA8cXWcBUaSryiOkYG5y2HW3g9RT
RNTkcg8c9FUzblFHhvBgZ8Ds53X55HRe2jeO9tuLmPeP83XoKW87BAigDu9Pcov9
gX0BW5TJ83oqCeKUmXXGTtLI69Hz/3Loo+LjE74e+dVEQ0UEnaKtYdGKETP/s6OZ
KAlWH+JRRiTPdY/dBnYOimBrXj+6YlveHOEuc3yciIAhEVOu7GtY8xoKGquM5C+O
s/2+fQPFZMCNHyrrA9FadOrWg+r4iqFmLJcmLbP5w1b76j7HT3RtHvbbc65Jew1k
75KbG9wH500QvRTM4s7vrGfPTL8R6V7SqbIYX+cnFqYNKOGvJrTRkhpueQwN5VIk
6w9/Nb8oGEtds33oll0g2mp9/T+fN3V+S0utz8UbDkhVYl3Rd0LihzjfrJE+4lFE
ZhqiQ3Fu3toX9mdg5E324YjWGTJRN/9xkdAKe/QS2XVY20DLsFUcAT0qNnlhC9KI
5SAoXT0xvBplgeX3Q1UksPMEvaW5S1jbfRvq5NCDEVsmtRhr2kHSkHRhqTpAyGxE
4a40akick176czc6dLX5+LLuoYHM9XCb55c9SxRT4v/Bz33TdfelLrJ4pWJQbNHo
2pAkHLOMXf6HYpjs7vfWER0UHdO+eY/ePRIw3SGpoT5edLfivFgoJ+5qQb5k8rGo
FN6P4xnrB94nIp/mdK+hsb8nAFVm0N3EcA7ZYuCdmHH61XxPTI4j6LEiqklXsFhp
VNl8v2rAncv/ukPB98QEcIhf+4oeG+X3VATwlxbw91FL5wGnCdxI/1WrsqhaOcFK
oIJQb5F5L5lwBbr1VGECThNS5HwKP6CrOZZ+LmKfNfARz+/Cpyoi4rdDoAmBGerF
x9cXSTNAGZyrgUab1g1Yjni4v91JgvOlZ817BSWPF10XAQkLnRds+pKF38XK3R6g
F5QW6nh8hDCLCzywUW23+eMvyjlYVLQ3hRbygWuNGL1IcSx9V9yRB47wm3zh86g1
E+8AjeSKt2brdBOuwEKhQfxFAfO1+zcW+6r+N9yAGcJFjcvRF8qFh/20ATXkLhar
D/A7GX164/6aJeqLJiAw0+NfhcOCdyEXoOdIKwbbf4MNaHWNhxwe98HnBZAtILjP
rBCRbvwxGtUZv514j6A6F7ZJ61vBmh6/NX0EFF/d+6A+aWqfgiTOR9ZYyULqrA2A
b/uGndpr8Et2ElKvfj0Xn3qwkCTqdvQXr5Ra23nX3+zdpVv9Sb3lRnyI2cwOiB3x
7DBQz1WbrzCVnrd4aX/EABIVDpIR0LqY4wHVHb1VO/6oYaTTiwuoQpd9W3nVmKIf
p5nvnsukfOtha6jDmkzZZ1eh+yer3Yf6EisuEnuQegZzKqHQiG1t54DoTHcpEBxO
5yhsJeNZadGhaPelaVn+8NP31U7X5EK2rhioTT/K3efw3kvbqwUMtgwbNh61w17C
adlay/cfiZvBf8q7KZ8iuNLbHidVfUR9krYNC6s0yGGEegGmPsu/nj8b66Z+le2g
sSjpvx3lg4yRB4LjqGN4hxxG3iSA4cxQXdZ1eOyVsuHz9Hp6zLTM3D76rtHE/+d1
AwUAoyMPgEosLFYYTIP1AN3g/9ivNbErZUW2jhfL1fEL4tYXBGk/JTtLsbtUieXN
23WxfInFe1zu2ImBBmUmGrOIO1aR+AtHuUir32BH1JlZyKfFSXmEHtZiDYsiXw5b
vw6h07ZCq/0/Ph0/BCgSZKkY5WoIiKYcHQDSZoFQKmkfk7ZwKbSKyVm2TzqAfBzN
XNgEUIxvLIcuPYTCRBIOdNlVoNVXhBdcIbLVXve6Fe+E/L74YHPWG/AnphVb2NbA
hIw8QdkCMpEt2K3Lf+xMoDZ9DgwGcSH+K3HfYDOCkOScgj4OQ3VprlA5WZSlCzUw
sSoSbAa8Evkf8RAOByCuFFpguhWSH0qK/sqLRm8uq5HDnadEtsHJncHFqKcVGAzv
N7A4CcnGK7/Y14OEM3dChzTcetst33YJFYnMv0RJ5kFw+vuTvHkHohFJfTc58phq
/lboVnA0fF4wTWwXKbEHIq9xVIT74UEFgeCS83PIHQ1EFqxA6pEF55dXO9wXZ4vA
ag6ZoN3hux+YCdbuZD5/0MEHqygQkhB4eqHFDwK9N87NXzLkGQ3kxzHMYOGmhmc1
f9hm5frn0iOsZf2kQUwZmdXFdjjIBXsYhHNJAw+foMNl+deI36OjulFxNYr6CzL7
r1qgsNfZpEQ7oYSyi6gy8+uhm7odCQktTKfNzUpGWO7Jy/9pQgQdVxYzuce65/rz
MxUUQXZvo6FlTyv+tqW7Z2btLRvjM25p6/rmkUu6Sw8It2wEXXI1aCfBnInXdPQ0
JuQP6KKHB7zvlzTGH701dgosp+U0XSjv9lSGuoRc/t+wR7eis3qXeXm59Jr4N/yU
cVdNXe141qKVOuQtTsfgRCZdG9q/QGMAzC3R/9aRQf7Cq3tpXTQDnS8+lAyK71bA
3zdC+lUBj0yxNjt2vKbYk/GjDFbotCHEdQKuXdebE+6+PGIXpJOkXjfQ3bQo8um2
ih1F/GsWVJ32slH3cZAQoZy46dgqf85dp2ZaOFoxbQ6fQ+LgvDBvHXXMYkFMIdgv
psbrdC65bXhjpW2oo+PQaKkD/EDsppC5KC0/1OsEfP5rqZJkWVwQJkXnocxxHFlm
q+S3YAWdDElJ801KM+yBNYjHRaaS726/IVK3YDNbLc9PV6zkpucpkzP07VQcBXUF
BtF4jtkTES7mNHooyfYGjXDkaaJtoBvCxu9T4snuke4Fxnk40yOs2Kb2KVHz7PAv
u+8pT2so3Tzq3zS3Ushbg32pUMYG8dq/SCQWeP8uUm1el9zehlh7JPtrvXALqPH8
aTysY01EGtqSt3761RC1Bf8Owjn/e9DrjWuO7TOwfxbr8Wvs53Sg7maIEO46dUc2
XX7BzdPZZoxTa42cQP0H4mVf2rJ07aTCWAb3fa9v5+CWkaZugNx2ld5+BZTrriWX
uyjx/aKQoeK+N9mPwaQPUzKWkdP665lnMShqTmIkSf8gdBaBoxOjEUaGKrPcVEFl
KABmRHYaevBuO0Nk15f28ONWGODp9w61nqFwb5zwIt7JJG2uM1au5GJo7N9Fz+Tb
Oh9iSvnNa3u9PURFBgUOvLJbM9/Lb1i0DPu7qrf+65cq9wee8Sl8EAsmIHTsnyRB
ioiBAB4gAAVqGaH0noYwsPMboNuLUYIZfZwxxc4uN8+eO4RuftB3dkHeFCcj40GW
oRJzRz+ILPDvGqR23ALLxlVV+I7S9IEFT/0FBvfzH2hYnbR8Ia1glI+9x8neTiUz
4JRiE5JRRcLSoPnBlIATgPCpwEKJ3aABo8Tci10Gzct/rLDZduDLurO9+P0ARHbU
mCNb8cMtV6AiRPnmXlwMBA/mJT+BlvnmbBKciUN0NRjxl8AQewFpiL0VBgfLTBqj
0iViLo2O6BaDh/+20BofSAfhk1RaTBACoXRt0lw84CZDajEEr130uodqtZFi2AOc
YdDl3JsBkLjbg89XMMHnm40MSTwGLOGVkjD4cfS27GWJdWzrhV88KtXnD5bJbXD/
oIWVN4KiN/V9dCxcakdnXx5m0M4SpAvUa6wHnwkfqWQ2lQRuGsutO5KpCyD4HqRm
PKxXB4nFhJsLKzX9eEbSTuGmMCYdfK5CMEt87cWjCJpML/mw/t1KHzI8cz+twboI
fceOyNKUReRB5rxLtsNs/s9SQ5wkVPkkp8sYNVFswWjHF3bOHAl+az5P9AmXdlsc
FYQR4TBsuOnk/Sq2bNQ7BMa85UflTmkpKtKUB3Cac0V3NnFLFk+yRxtcN8Dm41uL
FalAShrfM/C7yAKP0YEyo//+cAMmzi8u5FahMm+VuUJ45n1aW0s+aHOSwsylvrZf
Pzl2CgIyMhQSHQ2fi4GHgWZuKxxrWZ770gNQ47ildMpQbzt0dX7yfMv0ZuuUiDGb
KXCaPxQxX8UeCvmxynP9rUZwFywIZ6bDVSYOSYBB9taQg3D7hMCRXbWMfJ33B1SK
//MXL3B8Yf3v9HzV0dK0t6VyYXfp+bfgNcg2V9Np6h843+thCUYvV9/fXJa+mh0Z
SYhDXrsOh+GPghaEh6Zw7SDptjkVoeEIWGpMLir+cVvfBiO5oYuFJzr0SAP//Z8E
r+BKgxGw8BRHHGVhlWGwDMCkT8f6Vy2P0RkDrhZhLtRUijhxmibwqhZzQJzZFiGz
a9PLElr09Gt1v8KWCTjWJtr6gKBp6u3KHtmzlv4nPMKtP4mFLd+c2qqQHNKYVite
IfXgIkXcOL19T6arKPkhYjL4aEux0qUkwq7144xOo8mmIAgWCqEQlAB7fUhnCoeC
WVq3Z8RoumOrWvO3bp4Uftv/8GNzufxAj7C+sprOdy93wc/J23qlsBSPhbnaqzby
9Jp3GL/ZVsI7fFwHG6xswjAkZ+dO328CPFTavkqz/ZTV/arhXAN6r8jGqti0WRyz
tz8WUZsnxcFqG48qA02VmNl4oKyZW4CKx+hcPmlZ3p0YPBU4RcvlnQ0nCshDGj1M
bIArpZryadFeI1Y3yep2ocouZ6X0LrEJeBy7ZlZSpw9QBUnXLQXc/ucGcBQqavqv
vqDLgwim6/QSEzpfiEX4NV95+wO+qcd8AKW+ANN4aD/0ob8rU7A3xQ0Mc24+rg9c
C+NnXQ1+uh3GP9VErFds6oho0Fh7d7md/rwhEG6E7oD1iyVN7/6Bd7Fc1hPMOt6S
D2H5vJLsSknXYdn0C/Wu5vrhFvQ9Zow2k+dytfJ23vCyT5LNvZ4C1k3DzbqBIm1x
Lgo7AeJqfwbfrc1WYGVf/5FiN7mYnvKbjdcxHjQoBkIfuDlig1eGrHX3J0phD75U
fOnwUX/PjtW/rhwnfhhnOC12BNn7dsqPYhV9qUdeLGrcvq1iUUG1OR4jqtUZv7pV
4olFySsrpaRsiD64fKn51BMa5SmKWhuKGRJEM8DSsmBMxeI07hhI5M+mNNWHRO4t
XSWnx2OEWaAj7IcPesbDiAqw0qjDnvDvwi2zNPNJUApCRoj4SZZh6WxpOMpQaeOX
pfLnGqeIsjj5VCUa6WoAQXCOtm/It1LLdIBkSSdUZy6ANigoO1VRp0OAl+eGTJBm
iRinHOyYYnghGnu4udVFbTMGrBmuAxhEw6ccuZH0ZkymTXsYB8lQJmvGtMCb/D6d
KoL/u2f85RZHaaSJ0RB0tNyn2PRrLi6BR/aimp63UQHZaFHE4kG07RuYoJJRvYuc
PxumvwCXWPCUj3Y/BndZOp/yO1PhSlSM2i/OrenkDz0oz5thZItTWjwlq3JOZHLo
/hxpV9+A24Oo0fzTCRbKIHsva/EIyuzM75aLysmrA+KBkxZJ3Sm4d1fr9VAgBOpF
jf1lfb6HTTqQRBlkrAUCn+JeyzH/mYya42DDAMyW2OC7kIj6GwMrIK9lSxpie/he
ceHap2wClnUFHBwUatdOiRxqA+Stx+0S6k/0l4nLAYs6fn8lwKJIVAC3LkGRpVP5
hD8Xkvs/g6Q+LET0LWoGuVaxovgleOaDwSR8/ErRSTkk7553g72iiKoy0hNXIEDR
fSNtzw8iDAV0GU9bRHEG0CJIymXksCEuNLPTNWAk8/22sVUUxsqc2T5nmiXmgVsQ
pTt4JuovXj1NoudNNhoHexeRL0uG9oTjichrHPMEC0EIfTsxbpeICjuM7cQIK6lL
zcGPUIcWXDiCkjN8yZF+Dwp7LU0J6SarZA55xCjfaIsWjWfWq+WqDaKosR+3RUsv
1rjQZKgAigTvuuHdnC3UE0vToCd4X3CluhYF2hLrAIokNQmEwe7H6K9Sz7T4i5W+
6I3+BdDx/3EN8f4PDJdY1S2A6K0UNUCmFfTG7BpI2Z/mI7yVE1ltFagCt4mviZm2
xFdKsHGNI2OSJFoZB3eeH50Ak387ZqJUCUuUMdkWNu9c36z4ECtjO23Cw+/Gk9M8
fp6771j7v45ZKpwnchycizcQorepxSLnaoQJvj2i2ceEnxn8GGmvNsuVV9Oqry04
0sOXei6QVQc4Kkv2MI/vA2p/W2uyIfyJM8mntp3aMhbHitRSHH8FQ26lyTG7aarS
fiTvQCmPsKcmazz7OBjAtGBJakypQPmWF+GROUF/UEAP4pS9JhbY1V7qJTb+AIFj
Fb2XynbyqhSeD+mqWnbM6ilr8jHjdGWH8ZTcyya1c9DB2vSYaCd4w2yOsrGxoLrq
vS0iy5U/+3AIUrNpKGFmV1TqbMADa2ysWcEuQofYI48WtRtb0g6ItvCkCIaCP62h
4DXg5CYFSbednTKnK72UY9tf4kqxB/ghZLepbvHVgVJ4RkEMPiHRHc1Oma4MxTCY
btqYvtkTYTBEtlmeOAjv3DwzYuSebPaYJ67YM04mqoBsp9M3amm3JpoZZjAS8kdu
/tnUcY9D0UMrwxBBFX+OJ6mdYwm7JRT0q9Nk1YTrJtlpzA0wLf25yMOmVlGSAi2y
hCbPnjLfi8NOmKA/inJZ3jNK1HYPPu6GXzsF2XC/MkB5IxNL//ttYTyilSNrN37Y
+4h7bCJ0CaNiAEEj3rFxtOG7TKcAe4VNFncVpoMY1Fmu9ooLPyhBxqesqNzgYHoB
2Zp/YpmfDzxl65lEOU6fNIJMbLwEibBFXxSdWtpvQMZAeM6P3EP4k6Pd66evysIb
c5lN5t69wAsxVUwxZ9SX+pdlmBdYdTz/0zAYRx5/i4PiaV8xa2/daV6Pg8+bRt0u
LilWa4ihrIU1wsnWmuHASe3qmcH/wn3TottXE4rn8EWLsDuX7EWfRODabHSxu/xz
8yLzbz+f+LJIOQJQzMiWlzhTWgQBlppXO1dI4rIp0NfWeAWpl8cj9B0taFjjkJ2m
8OXzH57tB/hQWJpvV6tjuf1KCCOZociu5krbx4FddR3FcvpHEIVUCXIXf9UYg/W0
R9XLc/1AFy3kZVX/QUcrVzhW9w7eMWJUAbTht11mEI/XAdhd3bGTBp2Kvh5bh5Ml
+Cnka9IRmdv88HKwurBlwODk8th41G5ftwvYNd1UjRtMWC5Zf2SbxUYpPAbXXR62
n4OyWZ1Ul9sgH02tVkC2NscJlh1Lh+GB27kL8OKw/queEzjUwr9pGqqYJSil1Eg8
VEMf2m1ha3FlV2bNJz5kU76dOkN1BOgUzY8gg7/mtOjKLGVaGc5gJvH43NTGEAWY
n8V0qn/bFpfIwYde0fERijtNkbuIEwcZC4Lfl6ryoHAL7gKEcAKwFB6rZ3Cnq607
XQUW7lUpxUxvM2BXMf/D4ZIeSKWZYgtX1CW+tkRkS1045yk8lTnqXhSxPRQz/PUF
D00605RJXixOIWIpLMlU4IW6EuwDNXQ5rTJ6YX0MRNnWCkG+R0lCwh096GIXZeP3
zw8CzYoaN7XulAzQehMplbSnLVWH+gvhdycBEL2l46d+IlsPBr1cqF7kR8ETmolk
7mmD6GUjUtDH3iymiljZuixvIF44hipfS4yEGzVx2o5AczhwsRUlSD7IjL/wJ2M7
M9HEyOxluv5bBrZveTYZwC0/EWryJGA1S/HSsss95ivkieQwb6mdxGQ5lJKQp1Bf
yUffBHCwvjQeHzhaNpMsoQrYQ/XFvTpvKhp4+zfcwinAsNOfdR4JCrzKuwqwYLRi
/uMDZYoYRRi32YF+kJxHGcQXnlk5ty0stYzafgVQbIRzzrQoxfokC0mkVzYVdgMV
Kfrh07RCy3DVJs/pRsDvwiS9rRBhpqvVIZgK+NzmW8ErINCQcCWFk/jrqniBOb7T
90n6Dqh/tm0Dvuk/JUbOJiJGpfGf47mTGkDe4JGo9L7ngciMtX5rTjJBih41IGAQ
drHR/g6c1VIRPe/Uf46UQzja+zfICa0WTdrMxiS6qIS7BtsVb/ajE3At1gWg6Y28
bqfyxs0R/tyy2hpN/XFdAdZ0FaOToPr4x6ozbuwdU7k+ZU14K0d/UsPXl3H0NfJN
Tyym9qSXhAvBac/+1LeNr1qTd1vVl4v00nXPG1lCI0hStL913yTfMxrGB0CqArwy
hOF5EJrtlI+fWWmEvv7N5yCWWbgE1kAmiinwmJp2REPRHMavskbfatVBlhAz0upY
/uvKImVsZTzU4PmmR2kPKgahT0Qalck6s++Vb6TasQBqpDNDjWUBXUk5J0XoFL2K
TGAHOkNupbawEyPuop6jg4dsktn79WY4XJJPS/+5+IaNE+yKjQUQvfgpElU6NUGy
J0bJEFv8i0ZXNa//6YcSQBH61+qwCSWKRTz63QKYTs5fMm1f1H+78ZymMxYrp9ZH
qGDDAT9tbVxYUIzhFE4QOQv4Vc2MmlDMl4RdNJRLXCTty42Gxa4JB9B9fP0D31dT
3mJSagZk0n544VCjyXnqetaCheq7AbXZLwfZfoBFkxL9aN1TYRpsELbPkHT4fzc1
3e2g37d4+M5NA/1kpR1F3A83Sp9rH4anSXiYb8VVmEj6wD9NVr5vdSkhhvHi5lUD
QZZtgVMPN8zF41REovm23ejzxBmoIMOrg3sphUjPq5weI0d3+TkKeHtpK2Q6yIvP
0FGhMvqTD/qIe6oFevOZxFYXlRGgrKL6+b09I2xUzVZPvvpwPQ0J5KIFn1r1geXC
oJgqZOkvhrqeLb/ELPKVxxI+7ntdLShuFSWg56yzEWd2AU8xp0VOH0hHEuBt1qrB
UaXCPdykMRfI181U46nx56NPben9ZKCxH6AbHhTzYOMTqgrRNIDE2EU4R8A1ezdI
rLhGIpSJauoVK5SMmI+PVaLWPTnuZfll8A31pN9dx9kquIhssHxLFB2WGlof1NqR
tyiZxEuV8agLr7N8dNytabJNR7eCV4x7cmWxXfCEx39xiBeH55NtFDO/yBNYYz0J
ZpU9614bhcrhniQJjBo0fA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RKfrUMK+VUOPqI75rmB/pJuyFodhrLeLj3KqFIEzvGwe0iehYUd+eUvjnRnALl+0
MRb2Wb8jiBK80Dug59c+rdUHfJktSpL773VJ2ncKi/sRTW+85Po606l53PZdluHK
EET3f9II7uoHMViPYdckUczHcLo3ZV1g8/VrId3k6slmAorxScD/scSXtsUAfNKC
VafqulMEmIEYl5lHTCFWZPGjLflTikP/CBHzNYrBOJ92Q3u9ZifKgIYd0rBkt63m
YwTucYCfpjiavuFgNj7GWMHfiDeLxviQUoX8gB+MleMvhY+s2tu0oeynQem6ohSN
MAIbEnCBtwqGFd/YcVDHbg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6800 )
`pragma protect data_block
9/uGrlHRqBgw1UTH38tnvQS51L7QNTx16YUf7B9/fIeg+AogoohsAdC3Tt0F6aeh
qHF+vPfoc/cOc8o6B+UuaIMse5OPMpOPncvP1S60TOW1hHe+aIg+Q67q0pRckCRQ
ya1WWrw7y3TCL/PFIz2DRzUZIsG6dVy7/S+K/EE3u/3OTS6BsrtR6pH8jRQ2UyWa
wlDBegqtwW4cxJ9/+lZCTk+SS89TfXrXn0fmzYS/O46YlovFvYXmbvLJEOQ9tglW
TlsCrNgSviAlPDCwZ08vDJm4eV5ud7Hx4MkKtSfg9L6vSQ7lUhnZCBMhLhecA5jW
YjE8M42S8vgIsDSh82s6/5a+Ppn4BhyxNVpuZlcHQve3sKPD8I4++Ib+Sa4UexAG
XeHFwsj3m4g8jelpqQ1EghR3pp13KJGTH9olnIbI1w5Iye0ltxTip7wRW3mDuLyp
BAXQe8btmJQw80+vE1oyRWHDAHkzyIXaxlDxbDRrAGTC7cogVjtBIrJpMgrOztsF
6yr4G705+X+2vQH0zN5ATcVkHTDqhIUxVNXrqSjk/TRz+W6nlWpefXGbE+4Fp4MI
DjTWtBwnDAR1U66KWHRh+yUTCEYasP865Vd1nMXYTxhrzxh68gYc8SKUHuGOqHoM
TjWEsPbCyUug4k4H0x3l/TDUXMrMoPwPbIoZaRLWKEh8SAZH3jNBosNqhFZ4oGYA
h38vz2p6dvLowst7Ixj4zXAP0UDKdRc6185zPYmtJ9JleImr52x5ydwfIXRaUnzQ
pf8bc23UU9sRyH+I7nUTXaWwCXAbbnfaDqhXdlAHdPAhK7FdK8uehVvZYOtdA6RI
m8BVHdF+Y6d8fojQlyZDHvvxXYXzjWLJDHYu+aWs8K0Q/4xYgGHUZDhbOVBtte7M
mhMS7RffwEvF4FIkPtTQv+OT0NsiSzWmn1Aof69lPaKtb5TUQZV2i6IAvugZU2vL
uG95AH85ccGB87Yv5HHwwIWu6Q7r/i3pyKgtLwKaAKcIPcETp4xpy+1dYJIep3hP
43aOn6B0x/oiPGVheB743BxS0jWLr/WPuTiOHNp4c23aN1JMOc2eZc8v7MhlDktS
FUaxuMoCMd92L3A/EwIY6/pbfAZ1bvu95353/c06T7Uq0zm6Ci+uwYFFREyhAmsA
cFMADbXWlVlymtFsQJNVdAUQmmsoMb905cnp2pUETnpN+ZhfvBm9YKBNKKM9JkBM
nrjE/5reW2vg+lv2BButP1FV3ymsF/nmjV0L8G/a/tMAOutxGmx3osSL8dBqzK04
XwvoZlLZbwx0JyTQRkrPnYmB0/GUm6Us1ClZkI7J24VaaPOzoM45lm8nOdKqRMUu
LzZn3vNBwpoNGobUJgPFIOBAUY4PQKfn2+LdDrbTz4CJUpkREzWS4fStBKT8bY/D
vjaYyi4fZ69QgfdVNjmZLm/jLq/fSSfxAaVWPuqYbxPU/7xYshdGGa4vfjuNuwIJ
YwRue9e1oEsCJ3yy9YQimKFGBlRb0Rad3T4ROOWzRe27NDeu4oW80VypyEeUO8Nf
LJm+HIcaBf+kh6WZdJ0td1PerOG5nCOAl2i+bgUxCpvY0e4su1vi9hLZm6agHbuz
Iag3nRWTFAm+c6Nsd7OMyYTKpYqtWlvy2oJv5HASM05/ClgzwwRCaOxZrfTAyzw9
syL5PiqYldK81PIOPiF1faiEefQqNKHobCbj6XikvrVThacwYSS+vUECPhnBTszB
74HOALlwW5NPBKwl+9GpLU256Q+UKxyiM5cg5U7i+v0z7iQ3nEH5mx3yOBbmzAIC
/JrH+deBede0vCZHXTn0AN3m7vtqBBzQ4lLE+eO8SFcxkb8YcA6lisqgBneAUKH8
pQEEOymc5E5/XGENJGZWIISc1CskxUl2tbiIoEKM/qTg/VuxrbUQk/jBk6lEqXfk
ewWR+VVhg8nnBkxHaxRpVgBDLbR7A/3MXpylbiMroGsdodhm6cTPHT5NkwmZg2oW
UP8upiCGgRMaiDT/D3T6MBanQ5MRtE5cOUQCQIZbyLvivVwvW7c1TzsAMwTKB6AN
01xHY20kVwVIajNBRbAcbCjyltRK7KMoswJG3OJg/wvH/Ya674hKLGYTZWQMCaYY
hwvpgvMabJ9JFfwvmRrZcfkWJk1yWnomee3orZfc1QxUAWNlU6y3SzSgZK5Tpeg8
kGFKwIYAaNa2xUxUYZu/PiSdENZ/DcwPtFqDyHw2Azd1yz4rnOS3stASMz/uA6VS
IJ198mb5nULQ80y1TLbprmmoX1aTEUSMCM+pfzp7stjg4z7XxlEEhYLNePT67xPX
8uTYvzei2SuuDm7klLFoklZlbAUGC5B0qQnOw8/E5c2sJ6HWpVqLwVrCJvWrYCGZ
jRf+F7OAlKpsOfYdx1bebSY12JSB7yJxtg3D1Wl6Yo+A71zu2pcTB+KbJyUOUjXh
Ea2py9htCLdY6fSHSCfFdLnRQWZby7Hm3UvsZcNoV5tZbftF+1zZutWYtnb9XMNP
6wLxUCg8AILbCHIrrFB3YMUQHPij+wM6NdG8ENRrKUXtoY4j6mWXNEKcboTh36Oa
TkpcCRlGED7ggqtiZMQVEM1tir+W/dPCsaBcraJQPbZVjXOBdiseAnaAb3dZiCGw
mbCm+/8jWs+LknWDIBDTuZ3SICVsB1wZMnsJYIsPYDJGIamuoDg1oAl9kDvfcFf/
Gwiev2wt6bL9m5sPo8dyfSKB6JPw0R/vZxEQL6Sx4e5STyPAbGXqi68V6rC7UBTm
6gloohee7EprY7aNdRyHmZk5IfcGuOz9TytIly/c85TOG7wGD63ojQGpSCv4dH/m
DykMhoZPctMeJfnWubK5AjRw5dDMGI+Ke4/Bz+S676WWi3tiTObJK3L1ziBwOble
9sa1zn6YGGV/L5vitYsZTs/Vn82BIdxrOacpTwYtiIZXT9t2jZK5FwZ32FT6fZgf
EMbfhXzjXaruzkT67DdARQ0saF2dwCWus7S+PbkZLUzwuUuNwOp5EZVVnJ8SbN6S
Ek0twHn79MnrM8hRgzwoVJsOsYwvHprZfNTIS9g8gIB/LzABM+UciD2hPR+PU5/C
OCnu94Pv27q/jONI/PVTmS/h9j47JuOSMj+4nqmzdhxI6Ab7iuhP7b2e56LgbPkI
8nCSeApteWhGDHSlhGOgm834rOSY4vNSLcj0h5pkPLq1B6qHnqJ+QKprGJ0hipr9
JrnelqDoY757ABVGJCYXxA/5eDYpdmZee9McdfhaMPNv/kk0/Sjc6c+By8zClN5Q
A0JtL51/kYiRtlz+hTgx4aJKT9hR8uedXOx/n1tqvIc7S8N75o+jmZY9BAl/bR5j
IkawKthx04oqejvqaCuJqNFdgtU6Iw0lhNkfwceD/XeDuqu1AYWj58LOS4VFJ4+J
TQ7U5GQbhyti7JJTNhqSHR2L0XeVckDif8QTquG/aUpPW7G779m7EyNLXB+TXrjP
7R+VCtVp4T9EEoISdmfUzzafJwb7DM8dXBCCGnNcBz0YJcQr948PaxQrMlUIJLmt
wa4PBaWiJBqKnOYAdMIZm+Y5fjPV7nNOX89p2m9YuptjfVVyoV2kLC32kl0gcG6e
1M3M/cjzwDsvfuVuvN8ph0XxuIjYOYHi9pP49r3MjlZZ5/s+OQjAZArDRpN1Vk+C
KNt3gue+L5hUxrCaSRhVCg3dHhAsWup8shLqpWBfVHWrbxWLZN4D7gf3iC9SmPbn
QgFoKQEv3DYKIRGq61fgjDmDw4uvo0WFVSJ0GOf4ZY7QDEWs/8rvO69Xuyj9d3m8
r48POGwHX0fzhMJUTl1nUNbpnGEryonzcGI0YrGBIoFEhYYh3NJTAzJE3Fh1Oa4C
ufEgMIInZVPljaIjQ8DQBblHzFzYiW+dRjZMMs8wio3r7XvWn165IyyAFwgE8te6
YyS6a+4DlHticZnf4mn/ealf6IWgy7fVa6IxtXd5yOEVTr2GU6iBce5C47L3NeHZ
lNrZ7OP5s6Jlbhe0oxB4NeaWtgradcjzu8dcZ0hdKmHIo5INkByDC+1JnPJVNt0T
KiS6reAwLR/dRD9LATd3eI/0CSfexI9nDv1Ie/rkfZ3GlEWl23mYulZOyUdDSZ4d
qXbT9GbraPyO3I8lpo9rlDnlixY0AQCRMkNw6Kr7HEY2RoqpiXlDI4ySMa+Z5et+
oZQGgDY8/U+wmFdEAM+olNsxvMd6hwjaa9CYGiFCAhjLEr6ngQVZ4wFkH5jMfW7X
rQnsBgr3W4QkRWQ8EeW4ZrY/k1yOB9ylqZkxGp0hAQ5BtFz1ykajDTPFlc7nFHUu
lJ7g4W1JlCHCYcm3u8dfssFjDSYimTdJkBouBH5UMevYgUZUFNKOAWQSqXp7FQYR
bU0Olq0KuxDtKdzM4sAT0QszGrwHoCUb+4a3QLp7deVo0XaLY8oH44/6+7MM3VHs
szSCj2KimIFO0NI7jhXTL9EZUjrRBDY9PdEfVVJyIVbirvceYnTwETh7PKMG4vRp
NlT+3E2QwIBhXH/yY2xsJgBFkYrg5Nbvr1+m05/DbgYGCJv4rqjOZgPAKmlJRmAs
s2/hbZRJUY0oBSNgfFeu2682okmHo4q8wy+CGs1NvdhdKXCoCsBDVqUr0Kofg/dU
WKKLhL5Pk6PdVLp5kx1ZhFlA0MEbwBwu41S9/D7KvP/3ETXKv+z8e4drFnwH0aY8
+hLz+W3Ht+A5ODUvjP4tR4pFT/g9J7Ig9/+Gn/QwNKEFSMtxEXGhcwJweyvYDUj3
nRk2KA/AqPpr+SyegQ0Rw3Kos/5s5ceHmhLGM7CcTBcG6sxNWj0uNerQkt24hcWn
hJmruFRmDlBP+b69FtKs6RhDsOVjxinRHEzDI2dc2ke3FLY8E8DYNU+4yX2Pu10L
KbAdZX5ZULWXPAhJ3FjRtuRqDvoyei7lTPkcTT2MGBqinWZEDwPYC5VFlQ8VuJgH
gSINr0T33KipsMvRL5Pgc3HLGrKvNSFD4aZcX82drzxnp6C7iumv2yfqI8U7ymPb
Etiir68AiyRYbWWJ5ONdUASA5HHuoRi9u25Yi40DiIPgyurQlWftdlAxSjzZoX3f
mjfWO+A9n31CTS8KYi2Rc1kmNqX4yj8c6GV8Kp5YzL6g444GKaq206iDfzp99GSB
LDKCzwdUtsb8ZWY0CLsov9vazFJnnTegZ+gUcpQFeNy+d8yY94PE8rxMqP8RMSOi
gF3TRW07QFSLLT0nn4losBwiC2SiQmJl1UjOQ/A5kxRcWPXo3HpPyrs4Yo3bBNas
9f/g+OQnmZoKqyviBdXtDUwC4LwIBhr5lGlcP575mWM4DORvEw2kBrsz86TOvoD7
Jdo7n2zgVOw9BRFb4ilww7lnpOWp1DlYT4xe6LVl3gUUSwq0V/eKS60narbU1GPj
zNGVLZJ3vpuLvCETk/nRkndm3kSuCywGmBybCAx4nl981XGRSW7OW94qNNCT0IQK
h+AnQ1bsAzN9prxyBKQIOFIsF8AHu8xHPzCGBQefNJMh6gx/53nPkqAyPJoD1ISM
q7txFKyjHUXM0u/AKVOS6G8ARxglyAlTm389lsihEART4Y3kAH+J54WcctNl1nkp
X3qmOLCUEZA8xPVXSK65I2O5gvMwN0VNkHntbWDw5Oti28c1A8YaEHxz7FtdVzAf
OrHguPYZWgvUgqzjmCOIufH487lM/gL7vmIdIAApTbcsk+RN5sDnbbKoEE7Eo+VO
+iWXxxgSpyAxVHd71rbPXgISmDB2wxBt5CzQZ2jc+VuOBhHKz517bu4FsD90X6Mf
6MgxQ86OfmPrx5IxbaQMlexASbQIJ2vkT3QQUBC45UY/YZQndMsKFNxiSccsT1sM
NuV5OJ44Y3UsFzOAWRsGYeFbSnoFQdgJSaJZTpHvkl6OoSKXpZJkAYMRx7jazlv8
sitO+8qWlEkr5MdwR2ZZwk6UYHjTFAGa3i0RuH9ugjdxWia5kMDv6VKvZ7NcjUqh
iwpHrhyNpQsfTEbolKt/nL9dmZUllEETi8ZCLzYHhD2gDTo8LHqj1hTwg0J5eRvt
Nohcf1MGZrOoKVih53pKYHCdVNS0cpq2UmGAKCy3vO0EktwNRKd/BX5yVH/e7yv3
UxqL2cMweyR6PuIiu4JvvXqjkPnpSXpwGli+ogLdr+39JSv4ydnJEHkS4qHwJAqz
HSM24AGNHfzgxTtZ0838evt3D686/hvk9MZQfhvhTgCQREIrT515jCQxYP15I10h
Umpm5qXERTBmspSWIZ7Emet4oJvCfq98eXLC2/kc+JHnlbooUK7Uy2wga8jCJ1ZN
uF/UPPFmoOGN7j1fBBprWli6RRkx7tlQ2HV09qqjRYfvkxZahn7LLwX078Y40zep
Z1KeRyX9E3aJx37sGpKPuUK0jDN2X6yGQQSJ9PmPD1BO10Nkzw4pRHs81bsmipCa
Jh9Ps9+VzIfxMD/PhtUbbD7yXRPSFDxsdssDfl4jTGdZqfNd3qqJQONn3zPvQ4V4
HlBicrAUjh9w6o71C6+EaTrYuPRqY6CWOQdwF4fqyLtS0c77gE4NeYB5OB5swGV9
KSOiSgxYY1gUsjHK4wwXZRjeNVx814MUSgNCEs7iqo/7x0KM7UUjFPelA/r89DRz
C2G2CiIEtXSfHf1AN4/gEnFKitdkck9ccwQHuT/zkuEn6ZeJP9lDXKTUswenslwV
CtwsTME2vH7Qm5IvKuYX/ZDv0X4AoRI9kc1Gw+ZOCc9rOBNaG0xJeJkBxKM51EAx
aDt0dzFcCjID2DibjghezGWLkQT/eIAf6SrI65coiwc1Zj18Kj8XflwACKEUDw+u
gW/33Qe+hHYBnFneJez83fAyRBlEfacMcPZ4PW1/LRrtdleFkthTw2HupAfycMdL
jGZCIPqC7xwaDbVpXd+xFNiZMf0I6KukMPxTxFJUJA9OInfq0EJd8Lpw5h99qfWq
o9vgzye8Df4LoAnWgIcyWMbnhiCT61Q6IRgPwB4nzOnCRAqQyLv8KMz1eNL0JoCo
V8htnME9G2Zd/p3Wk3H0tIg1t9zHtJrTzQSISmiFtfepv8iGd8mH9H9ROOYAOVSj
b5J88icUh1aL87SXtXM/8ikzcHz4wiysMalL8XFtnYyDaPJgq2i20RWoN0y0aExe
HBfSy5mU7Oh4iTGyk+sK/dtJ7UB8zO8p75JFmwIyxNhbY8TdGbp9s6wKHvSEJu4R
CuZB3fBDDxd5J4VvBHjLVA9iK46kT5/vC/LLYIo0X4LtSlrjXAvuL2VEAGCjvQ8Y
3ERem8xBemXR0IYn5csGhjq+kL6O6PcQKv9H2jIbr+P9bhEcQD6uGjHFu1iO3ywO
LAY3+qorvARZ9/fJAUa/bQOmfXR3v9ub0IYCvSQDnWY/3OWDFDhc5ynzRQOEpoqi
TgS0Aqzz5XmTn97jtP+PPgzZ7ScUWddhz+05npb7dGQK3dh1auXpi12z+DBXu979
diCn7uDDp9kQSqFr/QVLoMQRvPPmh3Le0L3rbbaGMf+V9jerBST5pvR/rGFfIKNY
FvdUbgN4LsZCACLl5WZRCflIjZcT1KhXLPqkU7pZ/bK94r8oO6pBXplc14sNsLQ9
95dptJWGfRa/RjtzNTnEy0IlQNL6VA4i5GEFmInn9ldurt0Uz+2vYvsoZhxyu6lz
ZkJ+agDf8NCslbjl3BDPxgBJ1XP++w+X+QjHk0KjpP6qr78Ph5/WAydV7bn9/Wf/
NbprZpZOSG8Ha8C0O/I/RSLhXOb2DkLdu5E1wISUqHNSlYFXEFpA4APjfxq3OA/K
K/XbyaR5Q3b5u5Gw/8vAxayzx92wvwDYonaGTj9yab7NtvxP7nce3or0RszNLy8b
2oie+2OU+NsSf9V4peyk5eJXMkWBr99kGrLv2pqiJ6N1DffK4ue4sdz88uKX4rpN
ixZSO8KFKrABR4NKbHcqmABbl2ZAWBKkJhpu0TLBFIUz+GaEh1ly+Nk9IUlwxNlC
GNykdAubUZCJQfurJcl2pbuAir+fw/umKAI2Iu9a098wUNPeVE5DXFamMvdJ8ORo
9SIhjZ4mK8QzPZ1hu63kN05/58gck2XrqGkyV41BFFIe0HaFXFcNVtXd/g6tMhC1
lriO3LzvBlt5smIIEegh011fF12gG+taz/gExaPkZXEDwcWtirtfCLU75mQmJUyT
WGM0YY3hEjBJWzNtCXaauCUgwVv6AOoyMu8ee75Sb2Xmarumw+tqjrDD0e0sFmQb
01DllVTDw4eD/ta8ereAZiko4XGscyUWQxJnr7fmneFxaJs2zC0MqvTMG30gAoen
AmyqTo9cvloDJJhTT2d0DQw5PnWPi3/sjB4pCBAllaRck4jESu+Q02Kl2y+XByAD
nQjuNGZeMrUdn9sQTNq8tKBiklW3RhXizxOYJZsy/7YFWNoIGGHditeAddQPUSRC
gIaRq80xM1z/eX/46cUKbbgpR/ZBZbbnsHIfkhyjhXU/SsIJpQKFqKvghcE/T7zZ
CTH8E5TV3m2Oz2nev0xM0KjzNTVa85gP65owO8lRp8yk2hMPhzeREJzcIYQhQ888
zlBh9LT1zSQ0vsKIVw+9sQyygdbtiD3dG8l6MuVHAGlBdUZF+eO2YgA25Lw1xXwN
DpIx4m+ECHWJ0gtZKfN3vH4yirBdYMxH6mSo4i2THsA3gR5H87NPOYtCGvRP2Acw
VRw9nWMBXw+MqIUjG3Smc18YSVkGClI7jdMvIWUXLv/MNIUEfWwTEBA/wN4h6JOa
rin8I8GXwJLX9XmKzS06MdxRTbAINUiTKrcBpABTVU7J6POq9OdWSw/glVYNFNp5
pABjXQdV0xwIMB+npCBWa+WkywCQDg+7i9iHxeM1xmyDq3XtOgXvobMp1cSArrVT
6dQT/KtLIjgiAtT6rK5azvi9cghMRRYza3YzzLs9IF/yLIXl9Yk5m68thf7uF4Ud
eUeadojK/Rgj+RsC6Uihlh8qUm+JyoVWEMVwpHUoJbEWKQuwHwy18IKmOwNN8U6H
zJRyN+0PbVe72yaUCXEEIEEvsPaBgsEcNscJIGV2b8qXICLsxHN3bunymPgxmXbM
LDNp/T3p6CZYT5eB+FgFyHu47TwnHMK7ZOETGA5kIKU=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
kwTSVExX1hTcuFsYNbuSkv2vHJR1F+uX7rGzHJ32VKmHj1ImqS31UHnS/m4hCUiq
pOI8BrimbwmWppYr0b558S/tDxFbrcvcgBaORMDu8F17zUDzFCYF+P46hYlKLVus
F/9b3NFu1c0u2eB/6hODRetc287EkbuVmXTFdWcP/E7ipy+V3TdhvAWt8A+RoQU4
VCxD9E0wDCGteQQeBBNeddLD98E5GV8BXqQP/m+TOa7XsQ7KtMNGRBXZvbM4a1Yr
FlT3IXtZ3v9ZthYdm/1Iy/zx5JC/QiCgbTx1pnRzs3Kv/OtRu80quSg06KcNDJJA
wTHPfKOChO53KbjPgj0+gA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15408 )
`pragma protect data_block
empn5bpGZI84AeZPbsrqXRBlI2hFMlaTsL1IOMW+t93YsGf10NX/mret9ZXu20pM
caIMk95LTnfJ55M6+ASW3p/mtkwLkb9xklIpa+856HvTKlrXhFCs/OoE3AKdJcy9
x9IPfxWd0xVlbh3aOvKEqbzx8iCxwHLzo3KxaQHLQM+cJg5eip3Rgmn6ttY5l6Wt
Zib04Acj3q5PmX/EZOqmkiDbw3Vz8gi7jrHFsXVyFJzQcH28R2oNXMMFhKiJOztF
cIb9dq0DAIRdtJhZSj6Fbb3La9VxX/mTTn4SNU4IxlLnzQyXlXkS0k3wE5l5lkWF
w2VgXqO84c6OZXfRi0+ENC49n61USeygzlg8OqIPom9s587q9qwO+Q9pvGo+qndg
W7gH1dTQ3Sg22FqkvhT/y1XNU23kovdxBMOs3rRnxQtZGF2vV6F2Be5Zk/6zok7k
NfEGShYkl4SoPjBFx2aSGH6dhbP2BPChOa4JasvJylN5Z68LHKPVQYhUSDINFyFJ
S3pF8kb5vSLKHbnr7qSBe+xFlr+qK0kairS7qXJz8gE8QqkcliuixikN05z904Ut
i67qtq05wGyubJ45MbRd2/uM/nRN9FZwRuxagL3dHNTbQKlqtQRX2afdTb/FdsPr
lmUc5FJJGE05TGAKF5rD0vf25fTeXW8Tgs6qzf2kliKeHbjqg9kmQTVnIkQjAUxZ
MN+cw6+0nXwGHaMPkY80la2d87vwpM7LsJqFLaSgVPAbmzBZZi4yUMBOk/Ko1jXr
9X6ZPs2frNY5SldxR3QN6BPCsY/XGjXJcOyTQgbC+Tm+6cCayp9qtvlQfACpWKRS
BWMCywjj7RlLFNKZQWqrJUkVxplF77vLu0KcA/FJRbc55/6nmMQFM/Eo0H1qrB7B
Psx2WPxA0O82VXWrGV5Uijv06DhnSm44fgZD+1uu7M61NbP260FdxJ8rJy70hALa
lk9sTiMrjL2Rbj6S3SRUuq9Eo7kAn5RK9JELChtC/vr4RV4Iie3Jc5Ih1Tmg/qeP
kARwERxXltGP0KXisttN/i/bBrsIq+8s853J9aWSBDfFw/Wm5gSGC5JRnkEhknlf
a93Eq4lhYhuYpeHFSJECE8pi/T+6rW29VmbgDHhxx2bIs1+eO7vBp/16B8xTy1yu
33sGIFytJGl9h0rdMI/XJWYa39Q+PT2w6wSCnLt1E2+GM3KLeVxiQREsxrVPFRVr
lbE9fIuF6acyEtuuKGDyAkrajC8Rm+KX4CWldNpQ7LwEaaLY1e7tB/bSi8wOyG6E
6IiPttggLq9CmLo6hfye4gLdKOxXSEvKuvscYQEdG2yzqw7zlMM9tF+D9RZ/CctG
yNSM1gkLeN50nUi0JhSUWFmQ6k+9GzrQd3WdF2OeQUbfdgRJOpGoQ3mEtIoSrU9J
+WxInfBlBPjHbYiw2OLYQGM/bPAFhYUTtElgIVPaNAR53JHOgrtEJ4W+/ybfge6b
hQVYsPQnnZCpgdVlgWyLngHIueQgQ83BwjNrAeTyQAfiprguu78mYLIYZJ9XlMA4
IufpzIkt7Mh3inuAkTSwTAmuzCnEepITCU8hB28XmC8LaJPnDZ/bI/xrJwdwy+A2
luMRS6uUwInMm5zDfWVDWbIgGnSkLcX2Em8vdsvTuhPJ484aS9HnMX2xdgYAuz5P
YVOIxIOCGvq0/QnwtTro5chOwzC4k65fdoTUytpmiyTDEsrVPWTgalyqXmq8xn7L
9NcAf7Tmt/mAn4/1rjgnE2VRKCMwm/KsC3lkD/utOr/b1Sc/eqoj49ZLcRQnDPXC
0SCf8T//enM4VL6Xuu8rbwPOsRJJiOdqseULGfUG3nw9SWRsbngTe0KB42/FUc5W
25SgCJZd/QvSktBs8a4jVQpPGc7h9jkTot2NPKKsLVkE11ZJM75PIWkuo86H+nCN
1fXS5Ya0ANl8atM8p3daFCQTLrHBSkDY2l+7HC3ya8mDdu5RZSvmBCrf3kw+Y+/M
+f+R6xWcZRh+vXf7Q8LpVApqsGTNIBMCn8ZpEHRJJ1CeVH5FFAJH3jPOYddLhjLF
j2at3467U6jYLoYVmnMGwuIGI3cIhGj3eQUruiEl6/N2PhHHKgpuUR4Z0Y1jAYJO
VP3h26npISPa2OOcRdjkHtNVi8yLwnd4NDwG2NyPTDHOgxJ75uoP0N6RzyJ+tbRA
6J+eAngJUXBA/0ev9xyYOs+f0cSeqnDTi/uHph1lshJ9cAaV3yIHxxXfpT6dp/yH
60S4uYkY7IEOJKDOzHdV5Ap5zlSTyDt+1tjp9jOSnJOoLCd13CLIHUz1W31iwSwG
vA9RAEq5hAkxsVwb0vxIOEPNDYS5u1iTm2E3EBYHyLCQOlDSShbz/Wx5CCgcYPGc
FE6TS4s6BD/MIO89WsFMASgyL2CAfvKMCEuk+FLzSQ4QDACtCXT8KXwZh9oO9Ur6
eq6Xhyt6ErwImQ93A6y9e3fSSRlFDUGVinspZ/IBx1ty7Rp31ITuXUg75BaIDyXa
oFaSGXLbd4sivwpD8P8bLXjYKvJCQhD4OoCuOUEmloVTjoolBMLV6fLYTbkj187b
tl+hsSyMnZlIR1yMHceXGXLlmZhpSq5eP8NEUPpHHsWqOZv3y+M1WMMkxefNwjnw
BZj0j+auHiW8FpewJ7o2y5/kTpfl0OanjIws0jtEY8L8py83MPSsSEilghQUCw+z
TzHU7SKFDKJ6n/P4gFOk5s0SY2NMPft6vZStGrLsjWurc0Z0RM8H5VpGJVbtDVdY
m4tv+qGg6WjTFcPLjvwbDY+uvmo3Ujlcup5fFmB+8f0+WF4hlOumIWH56s6bFFDJ
8yb5gev8rL6M6T7kBDmom+HJGTKMHyeJSp5EPYmaqZkOqiyZHHDUFi+PErHofEv3
3UnEZNNhUQvTC90dJIAIqzq/8J3O6cWU1ADmLigmtkn6QIsQEROnWPpGnL/mGs+q
d27vDuW4E7A3/K2pv4Zb7BXqSK76KzHmlYDzURf4ELWcLt3eKdqt2eFAiBXgrUTk
1u0HcDDijvoMOEtJJ9H0U0JvR7J//enrx/luef0nKwqiDagx+0rE29wOKb1FABjI
zbxFwXsm8q7IUM7lX9ogV5QythhmoOhEv91BwKKNTPSOd4FJt07qNTygxOfkpwS1
148Mxjr1B3KwYQkWPqIgRm10wHYjeypENbVyxXFjsU4FiBTTBNghkEsQmxlmsDi9
aCKMoZz7e/BRDjuuZIBE78lvR3PMOzaHisKPHDhyvN/zckETQ8dvaMeV0rj1AXWH
CFFZ/EWfJCG9thlO24wyXbnG1/oY903tytb9JNNM+oVniNk+V2kTWVyt4icp5QkO
jBWubopVHaM2t/rvwkykY4U/dw/+ur9+Rn35HmS+pHJmZOyrWr3gdIKfeZpsseAt
t0YG3BwEvnMHrI64DXpCMIycYT8bgFwemZsLHvtE4qPLYpbogB1XSK0xRtZ9Blyh
MOkdK8c29nMkiadtZY0MFO2DrtOpMnMhFRvCO25yQNEOU0lzUZ/HD2oeLmSo6GVM
kNu1fuEzsN770BhEAktqSC/H5Lq8E/2T+FNCcKVtNzcJ5MTBY2a8Is1ebcoTGKfj
KEri5ZtJrahPlSlwQV6XNEkXicMbqqr8/KEtEqkGIY2qPffEhPSCblGYn1q9RLGI
q8/OEI0Fhmk/384hXUkmEzka5a1Y+K9/Ojs1qU/pUSoQVmejPfsgTiPFz4jVJVNr
wXiJPn9tslEIPY71bhWJXNkTHPlJoHK6SbxKlfezFWcmBBzXd+cwF5E6Efj9pf94
PR2nEhTBDlQIxVw4UwJRZh6ohOaUSxn76T+yMTB2BIF8gah/CuliSxzk7XriBEYm
WqzlbskJyjDtsp5DG8kiydBksy513XfPD5Kh7v8AUBVsZw8SQS3h50VS/RHskRdR
cPU0aJJBZTPyQkgpnac1quYI9qxGY/LIzU8bfYujjNd1b/iBfwlOCRjWQIKkgl69
QWIbjxFlGzgXWhI2AI41h2OiVjhLDrOhE3hghg7zB4UEBcDnHEoFMQVbdSNyRuje
zBpl6DP4FH05O5TnkDQiuDWK8zVmn8RBsRHxVdG2XvozQDw/1Pqlh7PYX1Sfuknz
aWzvD0aHfgNHNEYBxbwEqyBsmm/7+noX9fp+a/5KPDAWKUcWiUwtUblbucrrLzF/
3MicUcMNKR8dncIMKUhKKYXlmR7jYikQKjx03XQ+cdLKnwKaaIIo+1FXrNOZjgDM
Y29sRZlDfcPvAOUo+/iKqw07d+h3/u5IzkU0KsA3I3cbRN4BtBqED/TChpwcp36n
FV3PPg3b9BVRreb1XNwwoDZNyqPP5nVdUyLrvyHP1eJuEHLTUjmYme8sQw54i1H4
Ve2FVJKAG4vNHLuHyBX7ybHICYA9oCgzPsWrdRV/XnO8A17AV10E9RQqDSoPihkZ
sYh3APySWrcnb/4CaqtMaJ8iBWIuuCvIBfdMsxTGWpxjquCv3SwKE2a0Wadaf567
DPGHJfkfqg5IFolVe5iaRjins2LMaJ8OigIPPr14VI1bNi0+tWNMhJ0ssHV7Ku2d
BeZKisYUabh7h+vvYTtGSlqk3uQdJJ3otk0u+2Nz5018vg/XfcdJQVLeAX1rs5TN
KtVrbkUC70SH5VdRIq46IdTkdtc6bUOfgChC+Cg8rlJHiM6GdvB3T5QmCaW418ws
d3Z2/q83THwLrsI+E5wiEzIYk6OBDxo7KraZ3nufkz0lPmZ03E4Wsyn6rfpbPk8t
76+93lQ9w1vWegwJkI65ff4/Vrwb/Zo6WiAqsOI0dhIE7BqOiydTn+Z1lI4BQoCd
lYVEwtzsSxw5PEbmeYfhfmt7VyBMTzbQVTRpJ0O85TDkmxm7dtTfsqKiPz+CM3sM
PHK5Btuf6eBjgt5hAS/XRERQ5Xp6i82I54R6oNrOtnP+jtFQOMxvaP639jMoQorg
vXtI/P0R0J6vRu/blIBXHqJwFO3gHGQyt8NyucGetXyTUX0tLLf96aPYt3N4YD0o
MPOVeInLWOnm3HKIF8qVOW2dKsMUjngQEfsI1XFqxOJanfvOBr8e3HrDMvG72Wl9
TGoHCKa8Nqu+0kbWcgZm3m0oZsHi00S9LOs30LJgpCWmHJQ9KCPuuUD7bL/8QAzS
2Yu3oPAJ/Bx1sYS6r8QMmuq1fhpM9ivR4cT/dhhEFiJ6MRAjsPkY6aagj6JF0NY6
emFKEFmcI9LPUrSamEF12oqOgESbeod3jlzvIZA7F6X2BI0vo2IH1wrBzbSvEaWz
M8YNVOqTHd9oliGUPoIMDgXz2jkA9BKnEQvZTv7+Pa/r72AEcLBwz3xVqygob723
e+2qqZzsolkSTixuF0VKh+wwJVLZdxFrS9w7UsykSHh2tBMWQktM0oyZEU/n2xTz
HIvwC6t/q1b4IdgrQJo17iW6MsBschzAzIznXlXCC1DvWhtZ3tRbQXCl2sVZtZoV
2dt6gyCtujGpOsx8VVS6li4FnikgKWyElyrmr5jrxXMFz/+R1lvptWhwpF4nV1gt
JwWK1MAfBaNX33OqV+u5mf7SakkI5O9JsGMfGimRuERpwpGf+6E6BJmaluSUaxa+
GTchj7rzcNpLM2mu3BUmNF1Ksoffa9kNCJ0nqA5UCvxZ92+tn40+a2hH0Omcxj+L
xhe9ket6APGvDio2HVHswD0bxTzCXma9KyW4XDd4TW81r8S+9V1eKMFBIqVVKzmB
HQZ7oHvQjjQPC+M7hXBlWWq9gu6USTtbvvqxy/hut2/EIWNMckdZOb30OURy4iAA
e404pLnIvV45n+sXTnXHnoeMp2apz15mMkUooBi6/ujswlygaAWxeSQb1oqyhy/v
TMWJWfFMYMCaVG3AL3ce8fozrAxlyjEhC9jyY+L593FTfz7i3L67m6HU7cXvzdWq
9CNTHP5Cxk1esVVQPT1YenKwSPfeSOojxx+JeuQ0r+/DutWri3fo014enXtvwD3Y
2C+irGwZ2UuvajVvZAAl7w+HkKM8iHmFTmMJMhGORt0AacZf28e4ozVMfJ02lfc1
4aj1qDsJp4EhZTwu8NkCFjZi7yJM0dtJZWZ63sAbvU8Z17QLzOWqEYLInvvZXW2V
jFxGcPFiE1afT4aTujafdsPqWj6UVY+CxDGfvmyHed6fypw4k3Q0E16zkPu3hvoT
7y1FUjgUBHo4xVsAvPUn/yszkBD0D8IffkIhBsVBN1Cxe3s0753hBbf+YZwELNiz
kMEf0Gg9DpQg02ZQHRXm5LcJL1s7E/xp9WMH1XlDWTQy+N15dQyQYa/cLWGfgcZk
96VQy55htNRVkW2EL4WDTu6fHPhYUndgoC5Hc1xIzbxcdAgZ1dlKXHtYkaqYv70/
RZqB7ZPCM6tEsAt7u0dI1Q3QOw+zlmN7b9xdQHyIcsrrX2e/E1ny9mqKcicAKe6Z
tzXiMV+LPoCeDmMiEwQmlIEzqrJRUJJ8P9pcU3bo6WxQSA97waW+gELzB+zaUMSr
/MMyRfUhBPPtzPEGryN9TE/aq0oqpsIBINlXXx1Jnn9WlQFO4IivQe33AOLJsm0+
yCqsnyQ+XzlxvXEytnuIRgOanuDgX4u/QEGKkOKV4mop5D6bb/lyMN+7xZMKOVbV
LtyE3nB04vKQPQ/ctFk5KNsLZ1RJzebJF70LY2pjRNTctHDEsgBkanK6GttDKemA
VsuWM55cwhfttludGAm5tm/VfAH+ipoicsdq1mV8xOiVH6gXfr6hb/RDGzHfkS3s
qYOgTAXyTJwIfjvpHsVzbC1rGKT2MZwwJpjSrFyS2nSXU/fUYmNrhUoo7DWqsLa2
a9Xgy9wG99yqcbpmKTvnUu3Yw7jr8qOv5so0igUfnHTZNxI6VLf/nAwqO1JQs8II
OH/l+ASc5AKvmBhttKeM2RvuecUiMevPFrxhGyZhvMY/e+3SAXknc3pPNPcgvJSg
W8Z7SiIPKkbFhIDWmcSlPQMbqN9DEkK9NgfWRp+1PIeGuXfaiwNYm0ZZMO7QhKMF
aPa+o+23WlxjwDLYNGbT4L4OHCJv4096oEK5GC8SfzY4rTT9CHx7OE+qK9BdHR9O
HUHTKsj4C4Ktf+8MPLXkC0Z9YzE4PHrBeG3OTZMp3n7JXaygMSvo9AhmA7vKHR1t
WF18eboBbreFow2GW1PcyMr5pahToXDonRcts9L1AMVcSezC/Hp68XxgKWN4V+3T
p7BJejiAHBxhkLbfVmByJ3NRSzHxbwaW9g31UMMS5SlSGKFkjg4xNV0Lzl2pYVd5
IJKpoLrVncewp5FHtFAPaJy2f8+LqEJyhzyzIQEWFE3fee8CU24RBvrP+5b+AoPW
arcVEKw75ZYOzCWvrfNKgIW/YwrTk71vXOMsGFa/K+bGxEaHHgoVE5kWw+P0wCGS
BUjinD41Z1fevXDP6ZvF51Jmi8UUEcRvFfqnKXQsd++wwuMJqqUpjO7+mlBw6/1C
7A/k+z/tqsAn2fjWm5Qb0uyp3aAsKNA6BSr1SM20UGuV0SQXwWw6uu86CgEOlyeC
+pDyfFBiPsn5oq5gVlJkQOqPlWIsKhT2omsV4d8BZBWPoUglqRvKsuXfznbsMFAq
AhJUoqZCXyRuwOM86UFYZXyTkAHBGrxQpwJ/tAdZ3fVJhQI+ts9NbPbOE24EJzZO
+YyDd5Gk0Zb2M07pKFMJTRJwQa0hmEAYXIabltWNvyWr3zpMKEkOJffnmcH0EY6B
d+zan1cpHoUNmy9CaM5mtDHjEL/kMhDEgBDDhiZ52x370XHxB3WjBjbFVstawbc7
w6GfOBqIcSRf/dOKx1uFr0JEY7AC3doF0V2pFv+unPVs5lu4waeoB8el8Mzp5wkP
Yw5CujoWX1TBNRVDBYMI2rTojOduhqILiw9ZyErHrk3ckZGT9v8iTQuGrCmAPVn3
RBAa4lSITqxPYUKfR4PC7rTdwGM0SGp3AWu5Z+HKrNLnaMLO7tQ+gFWLBcj6FbqU
NjEBc1n+ODA59pVNq0E7i1IhTwEBGM5mNZ7pPyUQL0lKEKyR32EAH6FILOjNTbnu
3q+voqoJaEYKciemqBuL4Bzu5V30c8JjNjWJl1B15xCCR1UpzecbGZ1oJh3Rfozx
gMk92ETEpk9buxd+0IeBBhoopGNaMo2ohAsj/aA6dVJ9+pOLpyN1o0PdNmj0JRey
WoIpf0zgmdNJX5sA4LvfhdYLrNgDQhAu+0m5+lOx2zqcwbjdSL88DTjcFhD6qKYf
0rDMHRfpDZvVc4vTbQ9yLO642ZhmDd8u4or5fsW+q/4lSUbu/0fyRiRlGDgmbr3Q
JisBNPaOH5G1PToQruFotfDpU6BgZn5+AfwhdGbRVCmUEMtCcJDoRbxhtxYl/OLI
g9r/hzCpC/BIU6XM+cR2LJc1aLqIh946jApeyzWNXXNNwA6MJE76CpaUS/DatmTl
xm3k/Z2IvGZ7lU69e1qUhZ/5MzpWPoLJrZ3RVRuUYAQbZQbnzTo0rH/nnMCzNEUk
/SU4de4ZeBB2WFjCHnNj4oJ54j8+j0vPehWLKFVrXD87g0CohAN9lShxWDNQi/Bx
2b5NN+X8EXc8PBBvZv+3xAG0aJq+W3mN2wSSf0X7BUsSmdQcP8q1gCuVscjSNjmq
bPFWqmf95AXnif12LubgowKpbTISYeJ7XrEwOxeU2xPjm8fKMTWOcc4E9JQeKaQe
h013qfG78XwIGMW6I9/16S6taefZTciSooXySxqhPaK3jUgyDtn6LVRyu5tqSmn/
QxVEyXYeSk9T6gg7OFhEtQNdHuAyAcNCvWoUrb31YwKGKovOKRTiVW3mV0qOVyb+
22IKzulQBdfLiKUaNUHLZNR64OjGtXc8aifGNCavivsKdA2fUUgs3iwY58H9cBkY
P+dJokpROK/3Dlj5mgYJA5W/c3KW+JVNby8lcCyxGiZ8NIkP3A5SVytNi/EZe7ST
uqY7wrI3CI0Q+gcE1AEkvX6iQBA+A4/kkcg3302dpjnn6G/K2qKuA9kcN1MyCu2o
CjqAYoQchWlDFwWqXpjkM+D/VWmOL+VeNFngHzgnIH2EvLd8H7aefJF8QrPSU6aU
QvjjK6GcKYRMMvo6gheafzOuzrkroj51ClPo/td9S9cDTsDumtUEeobIPuyi8OKP
qBjGTBb2M6mWWF7TtBIKnwDhfkXKQfRqlCzohHP7WRlcprtpjeMqS6W7ngUYAleK
Z48z5oHG8B3rxjAICDQvDU2vnLABV0G3kC3RuheaaOXsrCiQ3Q43LrOiSb851IZT
snxS8fjc1eEo9ejmEXLx1zj+n87NJZgB9pQYXpeAwW3lsHluCg81eOuiI+5zj1CL
owbTnn6KcSU7m79CQ2SlMvefdFS6ex/cXcJjQEAunj7s2OUeiQdtGx/ziWvRC1ui
3b96SEi6zWZpLnKw1J1huavJyJj8V1BRBpraXENuRxOop1IYwO0KvejbiFjUYF7E
EbcHUynIiIMjpAYnYg7WK2CXn6L7ilQRKtw0Npc9B2bZLC7FcOFqK+HjLaOxy8KP
UaFyUaphYWeICpqCW0nCI91ZSuJdgk4Yf8CvvPaOACcpvlo+a6oknZHx36kRDY2A
eneyro1/L/zsg6nUrcKDjzSXiyyA7ONZHeyJFNP4PaAXCs2e6EaC5hkIScGj3rwl
EQgfAZwvst8yXz2R4PuS10Rhr6OQTmZEH7R68rIJ/ejlX/4ogDFAyphHCvN/1Rec
j6Ctir5ZmMX5vz8QhaDnfWeOQ+CtUpftYppjgR/NywIIAvihxRNCxoIs6dX+PrTd
IPYUkzX3y49ayG82qGye6AGPczMleNl79cus9H9Rv/xRMFvZwQYPkwurnsCf0vJI
vnDHui9e0zyH5teJl1OPt9OaT2nBgt0uHWNuz8GzTcfKbN489VkhTyoPa/tJcxg5
mr4PSas/pbdXQ0iT5WIV8j6Pwedvjtv5T0OPsW7qt4ir5Lsewnpgh/YZCjHryqb2
EBjygsdgkPBaSIKBxonVEuQk1qWD9/IZTJIzbEpSpv5PsfIKAaZTTcooGHMkdLK5
LQSSBuQT8tOgKaSffdR4tnomdmj1F+pQtmYKAR/G3rXxSnOJIS0LOtw4ofifsAQ2
/5qzc2N5FFJH1bM6PZdfBNm2m/HBSvjWT6Hc/gOze+fbJUisaMkBsoR7a96dkWgR
GEv4tSF6D2c20n31tNajCKZSP0DjGl7i/xIAihO+IzxKppgY0E5nWXB4/2QtlFtV
Usr4KLSmYt7Im93qw6ic+8hfnwdm3kFifQOi1ybHqPV/uU/on92QZFkTPV1+mLtN
qQKmZS1Q55G/xmVnwfs2IfsWMZpE37W1KixinoAaDcalQb6LkR7yb6M1dgW7mE41
wx1sRXtJc1gSK8HN02M6QF/23ss058pu2/n2gHuA+44FPlQlXk8S/Nu/znQvGTHO
uy3qH21VNjcnVJ59SJmCQEedje6km3jj34fFiiAzowobW+7GBcJ04dxkro1okGfj
jMFw+Y94oKsQVjqcq2VdN1KDr0iY1rQJERFOiTjurDCUpS5OnXGZxuJ/TsW1l0qj
LGR3ob/4bxiKVYP0M7FH2wzcmK363dKk82pugZiNLCpw84fx4mTQiN6YfMi+Rq0R
/0L3qNDY+0d9POqHmKpZoUxuiuI/Zy3STNZT7KCC2v9ULYLZStha6vjg7qumB+wc
Git6etHPGFCmy+Vy5oIQuePp9no4K5CwhbynCA2vUvQmNPBNGsPRxKPTjRi/NJS4
mg+2UIefUtnKTuVBEvX9ZuoyWWRxctBuKibsJnZ5t8MkIqdR/3Z0GPi7Wot5fj1G
Hv2A71jxurGIIxjcEo1On0d4ktFbCuz0AS3oHsQNVyR77wrom/X3ldTAyH0a01SP
5y6AuTgyEZoagMM/WMr2YXoRxvAb5qOqg3Cvkxjv3A8qWMXTM13511KaaqyH00Yz
isnvo8N/4RdjCyIcSrHthRvqU93JgV6upubdeJ4AXPzBHo27fSOob/tSKDK0GfUl
O211Rx8F1Ijg72KYq4VwCv1iIx2xCJdA3dGGazQYdpbBEwedulhQfpa/OqzFXaBG
hOMhBiuNqX+bumuqUxTjNsiEWWhHp//MmSdaDzFbPVf2C86em9sPgbiqSZH3tQrh
EAoMIw3PMamzHqz7M0ymTXTuJJgLL+aUjE+hC/ZZKz4xEgF1BtLvMhdbgv51N/iP
jqTlABAK1i+NM3Kv5PuPvhi7BDwsG0pGq1XyetkMZTbWFbxYSzRZj3Akidd6qiVA
nCycBgtOkyxbB7kiTXC4SqeRVroI+CgM8PdZXDWF/1d+eZzHPNhqoShWGTRpHJPC
DnOnC6elTdV6WOK1DtyDiaEWQXslJoTei/OB6yZBmN6VIkEFmOXSzLWODkMvuUuS
59nDRjvvQ+s6Z4CtEpU1dsWr5VxZPV+HgAqzi0l9B2NIPtaJDc9euBYb0tDh63ze
g3ayep24aOOoYdq3S1xOS8EXD6LobOUUoEzFsOxbDxH+epUrk9j7GRviC//ETF6B
HhBuRR6oC4N9yExbXAwtzU4+MIxpaXepBWcczhoLKV/GCqKENRfj/yFKCuwYD0y8
LQju56NoMQBor2X82bn7hcF4mN53ceEOQ4KRAoMsod78gVimU9wpNshXrRHavG7+
tepYcDiM8s3N+Ikv/C3k5EvzHfwnHtBjr9hutqb1wGOXS9oQIhj9X56N4qTBGs0P
AqOJ678UZOwfgdgYqWQu3DWi77iJSpE/NbFF4IoYvfIYy8D9DVX4JFSza9qiNzOP
vSZCqEj6xAutRmQM8Bk3Q33CWI7gtErkfTPon2ur+kgWSChW7RcqGJh1OQcVBF45
mjc3Ejer3QW04FObDHji/q4Yog/jvUx8D0tLmEWH+xICA5YunM6TP+HAGX7WC94C
pxYhbMfh4cUauw+yuuJXmdf1NyhWfjgVsnaP0i04SwpS3ajf8Cyfc7219XPc11Rd
xYmXoCT/Bx8z6TYjMrnFAfIei/wdJQBvEdz4Fba74jSxqa/TbetOWIGMcXZuyu8A
hNkm2ajy91xY37gxL3qiL2DgE6ilUzY0Y1XV5ttuk+Pc/74jgv/X3cS7+eFPWCuo
cXUP6AJ6+9AVesOFueKluF4EDS1jfRDCplLZ8wpYDdkxhNDeSGXEewjiFc0JvOWk
1VGZ9agcMF61iqh7Ew+VJrE98Bli+8n5QDOVq7AVi3TWgZuKs5lRuhN3u3DB5DrT
kLxDiBgJWAq1wKSyUieQb7M+v/i9lzxSbYO1MRL7jaz7iZqFYNoNxitEpb3EmXZH
GFYQVqi82pOeclRr4tUoQ795mEM2EMSjnhytH1nBnkONVzffBDQsi7gk/Vn27uM3
uWyTU288pi4j3jHYXI9/NyJQ8ct1SJaU3+CQFnb2/GFhIsA4ZpU9Js1RntwJktY3
LOIcqgIKrw6fqiEb4tw9nyHKDnmSdCvC31Es2QQx5PHh7yzhpB2qDZZG3fzzEeV+
qKy1yGk7PuId8geRtyvpQl1QfcPZgNvPYpwsDq/XD2BZxPg+CpiV4E2DPmbgD130
PDnL3A9GZITx87NtQCoVcin1kGX3CBsakJ8kMKTqDD+n0IGaScZVO/eu3/sp6r9l
cu30gQCgu/KsBZTzh9Of5r0BYsYJd3UtpiUkHCscN211B/vw8kQPqlnh8YMBvt1U
atGrUl3OFqJgr1+aQ7ahJ+qwrkyQYdPHT7DgL+p7J7ei6LOEufs1i71jFL94yCmw
4upyT0xNSub1LnUEwvP9AcGSa43CABkQh7Cye4rZNrb+nzCktjx304XuXhXLKP1C
ZLnVg1ncNi2AmWsYGyNVnoETF97LZT9LG6eeCbyXGCrM1/OqmK6RUO0naBkytOF6
lG9/2EJ7rz5LSr+u9wrHExspNKPScpeLuhK5meLUsy+5xYDbmnHCO800KxKiHAyf
QB2MSgvCqBubVNpZGalk+upkCodvQVbC4pQu17wz00a0O7LjfpSaVUashA1IsW6a
7A+o6QTaCh4Z4B5HYmN4BCOki6lCtpDh/C/Tuu2mj8AfapkVsZa9zaYbgnXvkGeZ
xqAiXsGD2y0HDy8Qqao/YWClaDOXwePlO+pg06HeFAAew5/cpkLQd6pK/+I6xoqu
w6MuEfjFfIGNzw5nUP1suwugn2ky/GAkDX4X4lJiuPzcWcTW+hgBukWB1Ju7ACTH
4CX675pacTKYc+HlOAspzGY9mm9qqZxGsozvz2Ovrrqs/IqfDzAW3n4HLmUUbtIi
FPBAfsBhMc6v4COLI/WyDWUOxlwxzNKtcTB+wSUtP0FC2ggeX68GJi9X32/Pa/5d
TlsE+J50CIn8ch7kkWvEjwc3stRAaO/JaIl9J7W+G646ZdnA6cVn6XnmcflB9eK7
D8LWV1W8Vv7ZqlCzXIanzfxcmwrLLKJ+hmmZH3Mgx4JGODP1OWacq9f8sSpw+eEb
obmnG45SptoLnpdMuMMAfxKUK8sVhURw28ZvS0gkNWUYNpoqx8REEjXAqXJaX33t
wESIZy+9Qe8/eRjd6PUUZGqSnEoNJWsjtUwt3/y5ZOitayay3RXpvKt13YARoYII
19ZfcFL5ixNekIgQDxqjECbcUCkuXddWORkPQqC6I60lNxJ6WjprP0Oc2K37Bsbl
aneMLUjap7WaAlSUxcfJ8ojAhxX84edaFANVLFtI//2+Re816UbJJ2Gh8NSMcE7e
hui1XINjB6nDpEZIYXoxDxs3vwy2NiNKA8fwBU2tUzQ6zPUIzdoY6iazxhqwm2S8
3GkO4mJ+0GDAcSi6PD32ML4yaA7iVKjiGvMhamcihGxlFsru7Jhv7upl+b2Dfqkv
r83Z3o1tipOVpniyErPeILuArmxmo7WvdO+sxVBel3DbeHF70cfeyAua1raMl8ft
0W8aVeBccd7ZO93aABjXhZbW/ZQrsa1NGFSWS16jfw8qvxpZHsHfNFlVQECU2gFQ
EkMBcmZ2pBOb3PNPtmjZcuuJqKgjs+Pwttrd8wh7Pcr35DgVOjzPTSY4b9/HRqjg
tX3vDHqyfUDS0IQ5r3ht6sKGOt+NzbD8aoiqjcPDLiI7hdqo82GjayMFDmU6Qrce
jU8e70/rA44ZhurfdwnmVQXkL3JGc2Sm8T02Ojot+2FossK3TizIB2RTzfOxA8Yr
ZFQFPYXbyAd5xhmpeyXP6kYsUAqmzvVM79Vq6r9r2pq7tPcLP3pYqmgOnGyoxlld
uyob+Pra4U/Hn6aQCt5ikbBLd9kD5z/TayOj36G2W2WRPTr7zKh3Qfs3tkDVBDSs
hii/nA91V01bfECU3aKKaH1bD8hAVejfw57A/gWWh2+69/LnnQ8oF6uY4B3deORA
mOMkdwd04m1w2ndj7X3nS61AqONIKPXzpIPpjzI71tNFkhILUuqLWBNpRzHdLL0C
YN1D8ZXfLbYK2XLyPVqjkhYuIFFbLZEPYdcNO7lZprhiHUMO47QqikxZ9CPOshco
5XcXGy4ywTuJ82IOSunqhKsjvfdKXW4GHRBleckVXi5wNHvTtUwEPDPe+LpRuEkG
issTldo0RXKqW4yLqNGqVeXHRd37+x87gjTyajCycysA3HZxMMy7Yfq0dD4jTZPC
agFQ6UeUZ+SLyzPB0eSNb8Z1lXir8sxggERJ9sslrHR5vNFTKDhNjZl38Wp90DEV
aWhGCuAZqkt0Woab6IHYw0JkNOuQTdlxC02TRlQOUiA2HPbK+KlyXdlPn0kNrxyL
3WA3tZFgKKCVlvJXCDO11AZbo4Hhh/BzFfAQTF7QIiyTROVZaBP2PgA2ElpFJWRa
TtmVSm26P58bR0HP0foyfl73DRwkajte1/sSNyoQa4DsKfg5GkFGRKBROJ8GPKku
rzk3L0Zw303mSUaqtoGLr4KS5KQ/zpMCLRQNP3EcwuUV+NDlvMErRzfjSMsCTSM7
sAvPcC0qVYKOdACJUQF4wdQOCHMJDkiJA1OnxiunEFBF0uEMyayDwSzkSej1jG1p
LbfTIV29Y3KXezKXh9q1pV3iC9LVL7SLIDtPrh824x3ei0MsvetXpeoTq9GUiS3h
zCnB819QZqTYSkLwJ8e3IJ2+2x5EzkXrCLbLL1Cc59oV2ZlYi/oNxiwR9DLd79aV
b5tNUB3oiwTGP+cgeKqXkDOKBUsAtwJj6kVFkSrMvpFfmm+kesqZDSA1gc5JWOuH
IfW4MWvBN2kFXq63wXU5E5QSFnoiUMVp3msynwiEzzpsmw9Xh9eZ621dn0cMgys2
4A3HvVsQolPf7gPDqGGj4IbRD88E/Sj8ne8cKNT96sEVsuH0uRvXvl9MJKE61FCx
D55SFuKI/zQ+5hXFcbRzFb5hyRbgWu1V3F6HjpI1ncP/CAUC9710laNQZ3hMKDoA
AwuPnIj2MpeP+SfTl0EeOZIbZ+oobQCLrfxS/do8VyqBJMd+UyPTjaeBwD8BX0CO
n4Xz8NDhAJ0LwqkuzxKBr0+2p0VVaMzsmEJClJEMOLjXZiaw6bZLsut4uJgSBdyC
P+KpF3QStxsTvcQOCpKnZyszzCEMOA+pGpnuchT3vzwNIhCGkNbtWgSz7MYBXAf/
rvtP9jcOLaTNCdsevh1SyuQkdzcs6til9GxPZnRCwvt4aohzRFSHYJ8FQiudSrJK
7xFSSmtTIvj2zLp1OAUmzeCc0M+dTD1HHCHrGMI9L0314Jsi6oF32ZoZ1Df07nE/
iru4vJ6BVtiKRkdXGnLkhIeeeFYvspnVHwpGRxNTupDE67mZVt0OXY2WZkcjhlcP
1a/J7e9fi+1jvgZvi3142NZyBekMfFk++SewikTFdJ6Na2Ru4BPDkQxwTnQsRn6H
fETFDDnT9qsk7t/CK1iqlm0mshRvB+2l57C1MHFVs8QpIJOlCK+hRg3C46NsswDp
m9QjPi9mhRoa6VGTLRWCE0Ri+U31Mv/H+2nbeN8AYYfM5N+9DqzmzDuK+mQay8mW
NT4ed4S4ABbae/NYLD991z3mDUXzkb4zhR9c1QNzVdHZ29lyv3Nx2DRwUMT1Aecn
1HDNcaY44HHFQaEaH8ax2OUp6jNTEYpAAV9AmSon5akL+CdY7v8tQnhLnxsqKcUt
tsad0rRPLnWjUiE2vdWkyNzk+QY6V84L5vIMrA2hzVl9kX+otYNymONlRYjXLBl2
wL7XMBcrt+ydG/V2duNVZe1HF0l3sir67CkJGcsA05XBn6eqgH0RoNTro3aaf9j4
c+kQWufYBiNWKDdqSHk2aN9ubZLZ0DN6Ahmafx0kGW6PuMUTrlavOzL9GZSGnIZt
tMNZTkfFE1Jg8HTeOpFHnYVIYvQ3r9phxmg6tSPKvNU/wjNvbDVLnK7VIhs51kRj
ENxreTaRZzV9S1DnRxvRyxoMTPil2hf0WxLcLjKG/6sPVwrZ93dOJA68IUpOKS6v
rHZP51K+ceEXa82EpivSnfjgfAaxSXUaYVLQmCY3RaEJvsv8Fc/pny9vkxwCI67T
ElrePrFxCknEe2bMR35S540OqsH9hy+fP+hboav1zQWQ7PuMlFiQueshcSqUmpXF
vd06ck3GJxhKLDtf1RQqTkzSXsm1YUhNNBm5XwHkQEpi6tcHDcibhsMn8bMHrfjL
r2iXHAfU/h+BQZDEeGPIBqLRwRMceNh9SrOJEYKAONKJ7w04+cf8pHPbKxMu8ePs
PgBds3w7NbRoxY7qMJ+ZXK39J8iEVLlGt3JK+28rk+KKXW9CFnrTQy7By8TzSbf2
a4YWyZCKbH59+4gnClXNmhhlyI+LaquyfStFRpBVuPtfqhddf7Pcy7DdhkRFnm3x
OFLwrtjlHQ3F5SJBUfhj4h2icz4kG3aR5SLUhOh19xca2ZRI57gnEHa2GgFchG1p
RA6WJlK5ypN2TCwqlm+tFqO21679MoZjlfMOTwuXu17JWyyAGNlgGnpug0kHB602
j7tcznSqWik2MVf1heA6kTSXghyw08mTSNn/YWSsxEslMISoPbwhSbpZVxbf3hmY
DeDmQQoqyMbNtmMdmPt2J8has2ed38CwtnSO2bDisiZ9E8CBkOn7Bmn4sI6/Htx6
dgJNBSEixDtm1zgf3J2R7MAll0XsJIuJPaV6yVrw/MjWV3ZuL8j0GKYryB2wcL4e
MF5fo0fZflE5LWnjOvzHVLeAP11xJRMRNffKeRDAApcixdgTEXQaG8SLSJmbsHom
OCzhkTBUJwO8p3iiQj/eBRjlV3ZjeL78kLW3kuHYhDmPeVcHaOC2/OwdFRguco3B
qxXEDQFtRon7GScYvUu+K6raGF/ausBMN+T7+OBQkrNHsIwojgmwLrQ5WA56UdL4
uCXX74+Rhmo4X3dI7ced/SNYiSPM+ajVX34i3QQglXFjCuAUMjv9aiQC+/kt4lmu
khNozoQ76gyop1GKFJOou4twrykrVq0WFUhrcw4XaVFb2qwV3frBjYKkFVJ1sqtK
MMvusCSDfP+Mf23UYzg5YV3eHpgfdikn8fGuqcbH7nTBx6Q8OJXrldrEbtddyMao
HXnHPk63vit7nIvp7L6IKVEHvCUE/XnESnMY+WCHafuDpYx5Oee/R+8eXwCQfJRR
+3M8gMognmeXw8fi88Sj4wkUQmIPVP7vcHcvjvBbvfCTVrKLZWpVIXnO4Zv1Ma5j
yW+SUmo2G3DcoAbqHNBYUqmYNF5IEg94LkMIyyD3P1Rl5lJBw6wSjjjgJjM4Cqbj
xoVX+7WCJdvdSvXi4WVuhDX3yeipvkvCmvsZeHrUDT4RQAuPSwY9TMLCYPNYvxsM
exnsokREOwQlQNOh02ypK+ik67OICja3ultBEFhoQyQWi8Na9FHkMbnL7qYx62A7
cRVJ/yLj2ybGPYsJ7W12/cdS5WjNzW+LJkcYO66Io3Gfg2O5cvoPfBv8CtuawDX/
T/zdOvyBrqVWIMle4G2HdNCiCaqUrgaJsmY1MJFb+QzlNAvCOOzf/1KRF2kohY6c
40gkUuIM0ElCyFx4xOBcNNh61tGxlXExz7WINM9NBfI4YbZ2Jbh4lOIqMnUundYM
mBFaVINW2SLo8FR5ByEdRRVf8uEJnIqz0nQO5tpbsyMpcgLlufD1aciMxnjnnE2/
paRGvz0B1O+uVN39QR3noOfNMnmzxLpMjFULIhjz35AQsLkWEaARwRHnbuhdagdU
KRpHXPfJnYH9KoAALFKQw40tb3HhS2eRz0p2yvA7ZGzAF8h5OEf4tPgVAzS6Less
jPCANlVFm1nJ0Ffyc1jqc1I1jLQG50a2TfVUPpyvdscnJ7COO63PqWBF9yDGe84t
LItzkIHPEejiF9h2ECRopx+1oIiHeQ/QkEEPaM+bsQDjaaFpoGus7pB4d2kMYLTa
PDX3Z2jcusAMciWmbvAPGQ0SZBzL5uu/O4udkg8rOdVVHFAXnT7BVE+A0PQGbCl0
CTtCMKztMWuIacENPGwP6Crqcn75bVPnaob0ts3g4SV/xTB6t9YDlgMNzNHh/K9l
Pp6Wez8bY6WdBMDVjCuoQWK/hSyar0CqxrgPR9YlOhqZhXSnIimFWjHvj2QF3mVQ
6uRKZksB1vNQnSMP7+CDn3YGCv9nXKyPO4E61UsnBZMwlkWJf9xfILG0F53034Vn
mW6jxTfvyGtguC9sug/ILhLbIgmB1QtrSKvf1YVHJ9Pwo9sR3dbr7ixGRrRwgt4p
CZV2cEU4VrowkAeffIbm+4ox552uwfNTA9bCpunj10AonKIdPTHvbqwp6lzdIjdq
7xdMfZlGNhkD58p4Xklp3deVDLRwVVFgSw6urKudhwlgI2BoM2aRkuKPEUDJF8TX
cP7ExPZCdo9jjWHbk7d+GgALm5VzRXfwJtK00o5ML24XWeROL1d/XEZIW3VRTosC
OuCFDqMUpmksOmFxe+XhMoPpxHwHxAU79+wnrQp0feQcf3CDzH1CX/r3BdmNj4tX
CorbttbL+hn6OECZJUa6vv+tVPQl1TT4pPwaQMBUqnuo+Kpfa0bLsA1yxZIg4SFm
T0E5P+I8JKMk0RcjdGtolKQ+t7QOqlIuVSp+7KnXZc6CIwaBcExAH9wXY3mEeveD
TCBZ0dKAmKg3ZkPXD2ox2rU8vNpyW7M6a4f8e+zGvll2uf2xkOVrpIaMyuDsGbvC
lcck/wuSJ/HjPkK6G8GGLJAxvNnOEhkct4d5PkizGnEupjjR2bUpVt7WTrKKEVSZ
yxIcolriSEzrFKtptfzOLLZVhatrpRrmVd0gx5UPo765QmjUvnRQQnVPvMvnbUNu
vjERysWXC4LHul3jG3nISpFvfGsLiI6MmLRoNB1jiGJhesOy5dEd5TAA+XgPhA27
SaeDkcAzsvW5yxYRtyO48Qy/iTysiR5U5zOWfA7ipH5hQUadlPhrgdhoeAOVU4sa
S+QrmthxEVFJrm8hCSYb+dD4EVZPBqSZtXYCum6uwbaD9nyjAMF3IAwB467PdTi+
DQuTCXPO2VaDmsT99IGNUpA54Zwkk/95aJ4nS4iO6D48Va9YNOg9FM5nFNzHP5Q5
bCFfl3HGdK4cg8VgPL6zCNtxciamfZmT4IWj9uJikaWRBVriKkfyqv+YGEKde9fm
Cyrs23NlhD2i+glGOMDQuUB7OXzcqbeZz2w5bg/6g0igE/6MZUvhA4O+jcb4Mqv0
8hjso8Onf5OdM7DBNMvmhsxT719xJKbol6s3AziDZtElIB51q2BramnWzbgg831o
dRc8tu8lkNatRVCY+LG2h00mW8YXewr+va0bPORvVKd2Twptu941hWhghKDvcNKe
zrhtH2SR90N54dtfvFEo1i0MZwKyrSTqo8mLKuCsm6Jneoe/3+DucZO2SHR+orhe
G354V3YtyKruNT1EDgAPy58UFmamqGTMH8/iOky1l6XjJDbT2PdAu+BOylJjx8xI
VBKSZtU01hPd4VZx6ea8Wn3KWoQ+DMBJr8QvH5j3NNZ9O0ZiT3JzZEgmE3aOi0NH
5SPFIrBFNbxCUwQYntAG2yYmUOgwtv1YvhdFK13rkX2SNMCsNE6eyMymhUjQNhwP
1umbUlmFWHoQhWD+59z2jSGKwJ0ZMBGUNNrOrfO5by0JNFagiPmDKbnEp6WsXIVO
3ZnyaGxIqSBpY7hwYVF3sHD6uF/cKhfbq7gSfPDcghy33XqGSxwBnegZzBtoSYRq
oWrXmky5uCtKJcQxBv8RwaziU3LpzFq08U1JQ12DRp38fzDJRsa3oatejbdluNtK
7jmRkaa7eqryqJoz/KWjX7cgaDrCcG14Mc4Hnxlk7iq4kUOwvkYiUXYktqfG4Dga
KTMc9Tbi6ZrEzovF7xR0hc7ywIryoF17ZUV3R0WyLVxcMMA63fGoloqQX0m1hxcJ
HSyyS3kWkz1LO4UJ5wAz5v8AXekCrbhjYMKbNzj7CZzE7QUap4V6t5NABtFFjI7+
4v25NRwLFRx169CgrxT829j/qHAAotq82+hU1VgTRHIM9JXtgE4gT+2sOnusmFUK
tc19Rd9a+MJQsYdtv8RfiYggRHrusn4+eSHNfsKx8lDw5Q5gwbuVhOhFzUP5KFMc
djE/A34ZnCBkwtuC8FMJdvOx6txH2ggqNHb5KHf8spc4ya9HiO0lWJkephvUEKIh
MjKdY/L6rjKgA7Y9pxz71YUsg+QsOmi0eeZNjQDCRfgDZ2d5W74sqBXC1DsFiZ8g
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bxghNHxokwKM500pyLDjMuDN36xaPoeyphYUK4VCXSzKz/qr1DpwBPDgu1f3Lc6B
xI9rDMnD1c94OKfzyNHUu0YsBrl/Q3+4+aerE7tnGG81mqZ5Bh/6dw53c8iZvitC
dZkfmPbmo5L44XXTdS6z5cKQHCjwnqM8p/SJm8UxXSunH9ICUM6rKlsQcGL+n0BG
7QWG5bdvfKHlYE76CxIGgE7plHSiPBxKwQMoEl+FohBEGFjFjzq76CP7YzyUGJC0
OH1jiAHFeTF+MWfTjD7uOFVHl26zSw+wXz4rrYVbQUnEKBOTEGIAqvhN2bOo4CXI
H11PZhFs2It44+ns4byTaQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11760 )
`pragma protect data_block
Onzk/eTJLHsjEiK01+OsleyzgcuquyP3s8XOEtpwGNsdOoCp/CLsJXAZSPPLcuIz
D8TShgZissXxAd+7Bp8ZWfk5iYPuJ+iuxrr7i2j7E7P7f8LiA9ZIlIL3bRxFDveM
QQ/q+71hiZdBX9x8DLsMxpfqVLyWjmfmTPHiKo+wb/8TNWLSFXYO2HJtD0IUID8W
Tr0DUMD4cmku070goC4D5XkFOoHfIF5W6kmbM9YZCbU9jnuPhJ3mnZjvb9JayAoC
N6OVhQFq46erqYmCMPm1aspIWgTvaqCqwaKJubsIY//ZY4T0yHOBR+xYDjnDMt+j
Z64i/l5NB4oiFqq/E15sWbwxbKsSPuf0P4FwFUmin11HPe2GzgH+1Np9rN/viJ5k
cm2XYC4+BKqi95nskYMIQJyPZ30oxetuMYuxHtFcIy3kPEuO+2sbt8OsZXUphFJG
z+n8ZeT9PVUqxXSjCZeYigWC3mS6t6I35mCmRG8G4gDgWOC+i0YOgZmvozwr8AGH
AuECQaHNBsztybTtt1IHVXsY+fLpSL4NvrSvqu3e0qSwbImnuxsdyLTGNH5ienQG
xJ3Tb6BblNs4uRukiYYxf4vOYKVeWFpvGAbEIl3+/YFmX6OLpJIvX8454Bgj55L9
vc1mLhAsFSH6sDtQTNkURS3wt030A8BfNfZGok1A0bG4Tt8EChyPjg+FILTSXOI/
0BEdh6pNW5Fr4cvoI+ux78GZ20v1vzYw4fr2pXznLrwLMDvvRJaSlR+DtCPuiTD4
TOJ6/ld/OWz7+/pS0pedmGJD7sOPALCdjgz5PLnIWydDH/w7WeqyFZtPa07iSwJU
Nh+DcjoNVVeNBzKsKu4RraHmqt+L23aq9j5KQ3Nn4Hs5O7P5XtjOlE0fVUDVj5wz
6+fqP9zy5YJgS9jjveMhCcI5prv9QDaTzWD6d+rK+PTlupNpo1Z/URQtYsTBcPAb
zrvm7NFJT5SzzqlZc7Y3NbO2tuvoyCsaGPbdraD2TvRllIA9Rf4lsBsg8MfZbKmt
QFcBsvlqhHqqBQ6X4UQzpiKXORdfcJUXm042Tm01M8E9tTudXuTNqMpzLbexnuEj
IHUJjd7fDqgEDSGnidIEgeeXsWvJ47yJQRxknbOwU74aTBJS0TAXuPThPqHFe4TR
a8Il1CYBnmewMhGH0ZcM58XPZTb+FWYTY+vk8rqY6z9CFKvgcgfFn50VVEwb/iKg
GDagI8BEbzzaCwhyx34LCwUeo1MG2EwvLB0Cy4eY8PlxKaw2+O+RGiT4i7pXBB58
1AplA19IkgRUfG+hN+H3OmJZckkRpViQwnBmD5EdghnwYg/R3cZoX7aMXd1kDLBP
SI07/V3IrhvYCceDCo/6zfe7EisJWyrtOok7QNyzuaK8mbER9wCK+VmMig8jcgZF
Ful/kFKLgQPhAod4urRS+CPVm7tHjbAW2ArpHbkUiURGVU0MvLvm+OT6WpAUD1qu
kgtCqj023CND+Bj/siYH7RyFdqTLRlKQ98OEEjSL+F2krEd9OWejYGO1kyqKpeG2
SynMdsCF6ueowfU43UZquwl6N+9D6M9lr35qp/D2Ywo4LqIQpSR91OTKVkRCXmgA
8lZ6a3VyaWMRMAT68OHQdz12vXR2w70sAil36yeOEb7MsTg3iJUd9uQcRw/+N1u1
wQQMhb1tMT4/BDca0txOZRLcRErzRlx7ZtyDFsGlMgVNi4oQK/15449RfXczuduL
FEVBv2dWvoydLQtNjjyOOoh7/og721S8lKHwwVkVlcl2lQq/SPNX11DAc2MXLRyl
TNcwo/bN9QJP3rNvxCwccE43lyKUcN7OKmClgn9v8m+pNIuEvmVQNcEnGOJlT4jD
ixIyrAOdfzVaZlq0bH+J6+4GufOrQ3WUIT1FHV9uhnzRg+6D8zCv83WBgMKdL9ZQ
gsR+2TiZjhbt02RKpi7hWnnY0mPNHYJAYRopO8LhlMf8/M7pJmEi1r7gOf6Qy6dT
j/UbSbQ2Ur8ToXUyGdrhzDhjaP5MwRvjDDycdESWjhPnHsOnjO+KKkswaaCERR/2
MKR3sqzF8wA58I8wX7xaFTCYrEF3RsZNhfvHg4648o2Qz0FswdKnrLm6v/qk6mvm
iAveQHkzsEgz9sqXVoZ2OQrzJZ4zsI02+NSrBbqK9v+iippu4VuKduh7HDgarOrB
w0yGMLdHG0XAk3XySGYt75wKaZmu3Jy0k7MLGaNb/kt6nA4EAp6raSmL0l+BTyBO
QSEYNPeMGVbDrWpBJVjQuCUL6zs+TU6UNo75a2m0Nq10knpVYpL/GV/Lxf70xjgN
aXnnIHec8srTf2Ag3aabUVT2C+l5SWDhWTSAPYeEoQW8SC0fx+SjNO9UyLRGMuTU
X6UdM6PCVZVioMyPabYPGN1aRB5u8W6xUtkM4scypGWSFGvxqUKT8VvUmv9qLtXg
gdn/mrMNXl2gBxjsGgF/v03PtBC3U7q28UwG6Zc+slI1LeTYvXER5tl/E1WsXK/B
SSdiuiJh8CrJGj1xORmEbTRq+PCNnV+6TXAasUrClRRFKCqxQQP8pmvWwl3qFxwM
F0oXzCes0Vc2m1pq1AELgm0Ybvkj2xdVBmrs+Z1Rs9CBikitbDTuDtWuWlwVXCqJ
9CAtBx4ekzLH/SuUtkhigKmkeZZP9Pq8UFSSt7l4s3jQSzVWZ0gCXfvhbjtBbB8r
kErrsdVW0BMLNCNLI3zHa/DOUCmycXlmIwG7v5lpBqHtuDMIuMRENP+ugN5iUG6w
vLPXRuvKv4aaxTWsobUWKFwcq/r8pSkan8LeMaIRxHp8iEaf3jnkqBWzTr5st0wp
wa+jXIlPuaxoyVZMFokYZ+FHZ1Me3pa2SANPLoi2xEtYAv0ZVPGsC7dGVXVs3waZ
unhncYslqm/e7RCMSIOag2xgBsQO4DMRm5wrKXPTaxO1Wom/zBX3TH49sXe/u1Oi
ixLgUsW08ENrSvMwwCe+/qGwdx56AI+0wZBT5RZ9dPt+Z+REogo8+yMC5n0YSXua
+aGF7DOrvv+vR9edksiA1PsdwIBZUPFswy5ijCsbkeFCBanIGPZ9Oe16jp+TePyG
3iXboH6POFXqLnSpvmAb1cSbiV2AHaHuSotNGBhewCfZZHwHjZkLHl312FNrrkxT
Zr577AQR2VMnf3TNvk5socdk68oEAdhD0qqE4CsbHJNcAzVNxU2BgNIhGjxywuHB
0UB/ns9Q7lbiFkDKIV+un6pHyHc+Bk5BknXTwhSPNfdwJ2Bm4igGtWRoUVLKDpUd
KrczXTQzczhyEBSLjbiw9Dr2mZrbxMIi77StNcORZg6Q6+eGxHX0ulgfY3dzok//
zcocOr5+8T3Y6gb7X2YCakTX4FdsRJv2nrAD7Bns4zedSsyGqf3wdhSQOOQF3Fda
O40/FDXHv7ipRR24xKNqa1hRD1efYLG1RgOJ3d4KYo6jgKg3Vi3gNtkzwOZMkNZc
Ie6/EkTCdJl6fm+kDFOGRP2w8NlniQr5KNgOr4xE6UNPg8Fta/b6AS6joe2Q1Pwy
CEFf539gigRCMpZfwmfCg/hLfi8LvGzu65HSKtUYvQHE06plT79zqIB+v5t2hCER
mZhA8DB8aCP/+XeEsrgKRZS+Q/dCog4IYyLF75XXLjw95D2z1n38B7JDKg3gpDSL
Usb6p0f++rhfQ06KluDKGYaItiigJHxaResqQqGDsHXrBYnxSaH+AX41Q0YEESLB
EOykt2YawdyqoQ8gUDtKzzvuniNxwQJBCPZyCWHazXLjwep94xT+Yh6f6o9Voumr
ZJ9nSqtN0H9WGMwMOxIdYO4HDt+LKP4/HmXzF/alYxoNLkWGT85Z6WkCGWYNCrVD
B9O3Znashe+gRf4xtXog6jXW6Ckd6B5Mv0+bZgXwA7j3kv0e7sQIM8genuSS1z4d
NDZNtGG9Jw/0/qT7huCbiDNHZhjhNanGdWNKL2ep+P+rdiq5vKoxLJliSge1cIfl
CUirC4thXMZxYE2D8IqveSQ2RCE6NvzGDsKf22i08pWeVoqsfWzPxHM2ScWjhNC+
71z3krVXNMyiOvsfOtaec2p9vLJFhzxZLKBFSx6VRIJScfdLgo4Lq6EfYeCHfzBz
y4gfIU3cIG0jQobKUDBPdN4JYQxwj2vtzF9ej5IXDbl3+R+9+kUmr1bHtxiUU9je
WxkxSw/qlpmUQgUGix6fRtK+Un2hpCqLfLF/3dLV4Dy7xHW7MbHDM7Ys+MV+As89
ILi6Xb1UTM1H5a3AlHeY8pENv7vJBJfp5kcff8R8kCSRinp+UjNTB1J9v+gxmh9O
DPCETyVChdfa7arwwAJAsMFtHwldGcNHifawTn9D3ACQ0QTF5GXHmPOHzO2G88+I
UsZ0eKlt3t++ZH6m4QR+2aUhylKHtCBGqve5U+s3W47idgAXcTtoO/j8upHKEFsw
9JkUdK0gb25wnfqSQAHXPDMGFfr2cQKNFJ3ZSw+/42hGJ54n+6+L8estt7zFqruf
0oCkxPOEejAGx+9HU7rLVKHCNYxH9OLKPeN8GNbaF4p3v5WXMo4SS0vNDVdoFHKK
wvM6MvTVgJfDZgFs4Pg94PGJHghicgN8IgYMsDYbzzkTf3+fbY3bms0LV8vLSLY7
QOZFh7mnm99jEax70rLMApYYjHvbs7Vo+g6+mHXVop/UfAEaGjgo8EwF0Mk26dty
/udes0gkhR4Cl3e4JGXmDDmguuYpn18TNHg7TxQWfBcYDCFVHz/gGu467bFkfnzj
+TzDbEcoDDA2J+kcTJPNAFS5kyfQjQVi1HlDrBc94O/1tBqfQFDGr+IzIfmKEmtm
mlTfXfAuOwbW2Fcif/p35FPiO2YiZsTcEtJ4WOPsFrgouOT7VCznzjs4EeVxKeHY
I1opll6YBRgmUd//fw+DiylGfW8adSPjxuAJGieY/TXpWtB0NbsWdyx7LUHqZ0Wv
gQIcIvwybNXm7eUh9Ryru9aNcKrhmv4JKM9ogVjosud41l6vgExsTWT/WqsoeGBV
pBZXrHqOcr+A2zuRqsN6ZZzAWDoy+CMG/pyIhxnR/nVb9YN0rkTfKCVnWMlbd6L7
Mxr1BfsGZZlkpExVgEFjmWa5WLaaI4DKdyqiEB/1m71RcxuBLADav/7gc3YlB3N4
WZ4EBmnKETy9oJ7JlBQuM2gmvdSe4CRClRShw33rRMH4SU2xl5nbNHrwol6Tq3u+
bntp5nAQgJ0SivP5pEYHXzx3YkxNLg4lyKEnoWzt+PNzBksMfdOFGyBDilK70qs1
UKJ534b+1iS+sc71lVTLnlDOa9lIZ2uas69OqeXnBCmjCUeBMyzq2akE2EEph0PP
jNSDpxJicWXxaAyca10Y8mzMjGQcmg1ybVzu47LeM5LbItxrpnNPAsgH0xpQ5y/a
YMe99W2HHNtjkq3+7QR4RZfiZNqpDm6G4f0WKjKS+0J8FZYNA+CSkZf81hk4KRel
BroqdmmQA+IA9Y9Rr34/F9O2DKiT6WGZh+L4gkF0hwvYjvY3woUs4QMlJRNjPuy/
WggVe77KL9pNlYIofypgqroLSy0sbWugx2RINt/B6qgbt1DUTE5Evq/aDFbSRyDQ
hcaEMDm3oPGftrAHEVoHNwLyPsZ1NS0+PKJYRiUyeTMgR9FxnX2Hu/22vvb0PNNN
eUMoxst/ilDuMvCIrzrVAedBoB+W79CMAHBu8MPMATBjIjNncOebAphC4rQUJSVM
0csYfJvf3FyJ9e1Lgfn9410d3SdQNVOmHHt6b5a7dRtM3p3eZMJ1W5/fxQGTEHFT
aJgH/DCeI1R5cHdOizJWVxUPiQRoEbxAHyGOKjPLgtbVCxvbeD7KNJXIG6FIGB0b
rVgQGYrRBYs7uMpniX8nTkugTZ+tiCsD55dqOQ4jKEOpHH/OqnQotE5HLPNtFFlG
WCt6aSaGjfl/ZUK7lHyF5QUYoDImtjXdiaiHkwrzgimAoZ56NrIDJlkrqJUaTzUW
QVizdwRvzeWlbbAFSNeuzM/gYnf8GXWWvKiw7n4Hh+rKVl4hAQSctbd/64qbCmai
8JJyz6myCaGaL2qQBYQcBsmbxdpH3u7gij8rrKk1KLEVN+uTTt8/EGRiNvp6f42+
S355gPUH7FJdqaclbP1zi5wf0OePhinXGZlS5TeBZrIh8mf+t5TBe2LbN7sUWKmL
Wmn8TGpQZPy1EMO5Q3cvqiLpBEPjj7YMNYCBpGjHs4f8CAOZQTW1Dob5WrrmZj4l
eFWNKzOrZAlqNkx431FS/ubsawHwnjjfneF2Y6jhMevmqC6Em+NCVQ9dgWinfEsa
sqkT2oI/he/qgBJrO3dIrp4bz9pqeVm7aNwVD274v084ZKhc3LZ1ao5yV/iBrmW5
GSijcWaKIVBUqYXUdb1N44vF6O69NRExPDeTUfoBQrO6KNNL1vxTjeK1XruQeluc
/+R6sXyGKpDej6Y6sDbgLui/zcK9wguaSWHUnzOo0ib74azzD+Fl61yL9fVOHzNL
Uk7qibf0Qs9utFrOYKh3+hD2ZmADSXP27o+EIVx8hxXkpSPaerQ2gYpv/sqRRmkZ
jN1bcuFXIJtInKvBrO0Lr/CQ/iPeH5AdCWnWvRcoMsggkuczE2KbDoMzghCpPLPY
rAwtyjmY/gIG703kwwDj7GoM4m9gHuRhgFSUGfKeEKSh4KMEOGg9r74OSe/HbMon
tZlrGxRNZkLDPWxovl2GYSHgRrrI6uZnZKrOkmhLG2GecD7LqWOTbjU23JQYUQCd
9jiNkyxVbygjH5L3SdtBWqzM98okXSkE/agQDqgEjNi5A2DSIZ2dpOR8VqoUblEK
JTS81WgWkzp7KXbloPl22GEnjDoGP83yd6M0v7l3zE3sjOlsvUvOBl6x6EjC2yf7
QnLti7IcAjMJdplo/BwdbgO1yMzUgyEjImYOVtaKgf+p5fW+7vyzRD9PwCTllE4z
FsvCW4Ly+iZLHc2CmvAgtyahXVWrvNlrHfB5kwQnX6SpxKAnX7R6HB+3FMSLPbUx
Y8CVFvaM1EDKvBhVYLT+1OlcNF5Z4hsDwXXueYoKxN7BBJ7IuA90PszhCcakkIdY
2ZoFi56MvgBuzqfjpQvZ1c6LM9ZubUPp/pgSq28mIK13rSpDhTkv2Vwwz3Bri8oB
nOtbFA+2dfO0a4t1aLDPLJ9razYaw7ZexdurYKhBX+TMWE49coCDkzxpMbUh3Z4l
lazJ94DjAqmnXg8p9LDIX9GtKvHpK3+W2tB28s0PiP7HeiWKfcI4WxQDOyuc523G
pErc0ZccgaWNY0VF9T5BzQ+yghAekDx6btwaK9bhvIiY+fRc7bT9dyVyOaIH208K
dbPSLKnZWp8Lt70HLHEwpqHL4pKmJLpWYHAQODRp+co6u96SEIjU+qf2+yyF2zMh
qlJpnGFtqabGgjL33qKkUFvMFR8bFrStNfCDZeN9Vm04XqI6KgphZjexl3xBj5+r
BvAx0oolKtap8I+6OvxycOT4J/imcgho5MOZq8gy7GNsIg9oKxJjL4SVzZJRSEue
tysV4CvJKi7PPdlSKcGmJwpQ9L9f21ydxLXSvsPMPBOXYhiJy8zHcTX606o7cdOH
6q2f+cPGgLUYEiuqROetpjSPj2UzS3XGo50j7ylstfKlfKP1VIvldzoCcxhNITSH
tDISAqep76uRtVXgdEqbI7c2voT3ruXXWbOTNGOXPaI/I6zKctuVSME4nLrOtYNV
5fX2gzYK9xs/s8SBk4Y6j7nPZ0Tzi+avqtWZK9Ra32pVZ/Wbn4wJdQZDWPyUHxw2
Esqu+z0DjEioDa6tMlRitrpR7xwdTiIUtFRtTRO1PZEYnL8Q1jmJxYgvMGTuHuZb
JsvNXTWau3WLkeUlqm648l2cfqe5rqD0X6XWoH0DwBnn2yVnYEX6eNQn1TqAhgA2
16ZIMxa/apyaLW2jXegniVyxaKlsrbbbwSCgLoKfIm2PGdYGjNcujagpjnGvzTUv
+ehT7oPxT9BlpOoJvSdmt2YdDam5RFUTK+04VSML0rCa/w9TtbMdAFLRcF9p+5ph
V39Ekt5Nko3fSv4pyPWZ/leLEp/b5Lq5I+k5xQ0d/IEYOVMBYdp4PC8Y6KM66U93
gARHsy6qNf1csaC7cP5ebxAm+tRDci+rHUnydvQTOahUhTwHSIz6F4uvKY8kEIww
mUisKj1QqCuYsRS12tUrDoCIZ3OhCixT4Iq6gUmS4upPBfqdvuMueyCIXG6YQIxM
5cXt0gcgTwEJGGbwxRwutnSUyG8Eqe63PL2VyiJ4L489p6+08jqSdmErXTITO17j
nbvrxwmipfKV4OHKnMGZZ5pD1HY8qj9E6hMHas/LG2yD3SReWj5ezUn1RePf7tg/
W1QGwh1h6qHJQFg6VPiKeqO6Xi+zlPSd8cKGD+YoB7zLSB/BirreNwrZFKXKV0kc
/mmLK1Rr95zMe8XAcNR8OzTn87Ji2G6OJ9s+p55dMdWSyYUBcSRcLBk1Hsn3a0gm
u/sWaAyZtdjC0dPvAz9zpx05rk8uTKLffghJ2ocHkXONfLhqp4juddsxyGKv1r/b
12EPPUo5WZRlOfz0rYD3ovXs9YOIsEpVitTy3D4s1QVxBDczTjYkDx7LEYjuCmmD
5k/uWwAnrHqk1EBCsuXGuSqHmRgOKL4nSFUy0/Nym250Nf0Qp3vElkxxMgI6qyjj
jMizwfYQ3Qfn5d8sFrGnqFnyanrxUWRmbSvBesQrXYqn73ZIMs9aXWp7Smb/RSrK
h9+aSheG/3apV41ZcuASPmF/Us9BxbmDLNO4MlX+dq7HJmyFQLN6rp4PsgzLLnEc
VfHQ6uu9PFKHYqQFw4nqKiyVYhxoZUpJpA6Y0yOKMCGuCslEbyr9SMK+u93NbXu9
vuU0jlJva2NtPL3nnzuXo7Dc9tP4SX7l+ZEeo6Z7if3LqH5KUWB9kJGVbuH6Pt7O
6fbcu1OElps95ZvAFsLpHul1H4+88r/3ga6Mw8abc+Crbr0+QOvNC1e5I3HOXmtb
GsyLIoRmvNDDmEXHeUVOMmgTNa5DXO28K7WIhXR1PQHgQZvmNE/aHtZ+ACJaLH96
9vPpAzTJNVUOa1fKvzBMGb4Xag7OQObOibta6oJhW+o501Q1XiAHP7gu28+XnpCt
5ap0VuVIYHGU3nh9zZ8ibJJClqko9lT+Rloei5RMXBYt1B99zUUZO+5iaoCXxcII
ohgRzePzVVrsQvIQbv/z4tRVxIAcDASm5035lAa/xcFwGUlvD18M8uXVQ5Tf0fnF
7KYu0EY+iBihAdYlYMqoTBixuRHvJTXKNqC3vIKh6eyyOz1x8E4R0Fy05qMYE+DE
ffWVjJ9KsgGy4kjFOuOHXhBpENisbVBBLCTCtp6WLW298Ems6+RxOO5y4o/eKFbz
2rXal+M22/WH1L1wnjWKLnvIiXSVE8pr4JBJWbSdqZVOBteq7sE0W6eFR8Y/KGaE
6FEQcRzeE94w9zu+AZxdgFD8HjcQVckFXPPcLnL88XruB2QwIQ/n+P1jK0rYnbgx
Y6brcgHpV8a1DsGQt26gzIFC5PGRjSigzZvC1vWtKmnKXart3K/YRWyEatLKWRbK
l7t67HEIkN2JOBlWYbWLQgqlXAsOXiYh/dGoxV08ZUo/oEFk/0+Dphy9FHgO9POB
2aSP+AvnkZRCcdi3BUAqKnwnXUmCE01QxQBSjMh8CdBVDKfcvDwFnrfdkI4pPIEt
op5QPdqcvyZ8Gb3e65lM3kdUwRgTmB37Krr/VWzCozSQkn3LnVh6+9OMcbITy98e
wAWgtIJ76rc7HAK9JCndW7eufc/RoD6mgWqvG7Ui9i9RUJqFRMY8ILzFVkEvGnEU
GSic/mP7w955rJaD8PYp94toWN7qXn6CsF6QCtv7wQQ2/cAMq8wfftFqGa/cpy0f
zjTIMXhY+Mf4b/OetKRjHP5J5xveG5gU8+QfEqwGHGeUx52S6/liy5Iy6IkKQR4k
nhpJ4TLP9Yq1/WilA0qPs/z5/WlWFz/eDHf1fWRx8vaSykDf76nGlSbOvzVrm7Sy
A6Vpderp9jekDrUbmG5xxXHl4RkwbUXXyJ0i5RH+fdKX4eKvm9100b7tjwT3vwSs
NIIZnou3BDj+NEkc3U9UvpmFxh767XYFZcei6vHC0W8IAWm/9DcAmf45sLvbVGBr
F1+BlxSuV/DCZv6/mDWp27tXSz9FrSVLmpFEbVP/O5Oh6jHa1YeDuaNL4KxaMLob
kbFBvtFS2Cys1KhAopCo1xb5wECLOvsYbgXvAha5exQxfjNTslvemyjLAxFGTdTV
whRhDrJcP4ipyvK5J48XSuhov09izoC2JgzxFQjh+2Q4n9sxVZg8skHaVtzLL6Nr
FWXyhkDoTtcbxwZfMrtIdO+n/6k+CX7EP1fDIaInF5QwtPbgyaxkE5rA2UEn88hJ
1WUS5UQcd3YHNVcLwqFJymTeveaPFrOnZN6Uz0oekd4vt94loBI+7fspxDq+fwX9
nykwBwLD2JgTw3ZP+STCw20Q1/ohmZcWeaFFD+H4Aw3kWtY0Jan2eaA/7w15k1Px
datTXvRkJrrSs6UjojqLA+Sa5jykaUK9yF2ygN8qtKApr5+gZv+wsex1aEUgK08T
IOfJcKhqpVBITqPAp5fJJay/eYO5Sg5inYyOhwQ3xQOb4gnPXiK7IO+8BJuEo5eg
ooRG9NjJrpRX9Onkn1d8lkR/L4gPohTjUEGUfeen7hUGJMkirq0yumhCY2/4EtlX
UeqfhnJxTL0RQ9YrQwNj7BcpM8sAXO1bxzJilM5FauDVBMBnVfnuH4d13gs81uo8
D+QSzlRRm7LBM9QsQ/F7HDJ9RQnvsKsz337r9/IyCrKEBu726GC4CZvOCFZxskix
8ZI1+1tUx+x6aEouJoVzeMTnGTV+/u6BHprAPvwKOofFtHwS4I4zluVN888IIOOZ
XvM669USz07vcH1z+cY61oKcAuI3G+HXmXVFlkhEzIZwXE3ky0Bi/XJXiI4cVpk+
ehLOADJygsv9ViWOTBqyIDr8CMO4RG0RFxpnNOvh1VcQQANPKxtu+3YrYNbNa7FU
aOFAZhbjxOiEJvru8edJrfKKrit8bbMrYh8f3/JDum2HasGm3QxadjG7FNEa5sq4
p0X1WVzaDS5NpmubvxB7/+zs/EsG1yWwqMmBuZywikB6IlwuRu3J+fnDo/KioS5b
83quHzBEIVmB7xXZUny0gHxzPuFV9w887NH3pXQAgvlGS5YZ3LZJXakmF3gZuo99
aI54tG9onJONUTNWVdvCCAxatTNI+HSJ9zTN1xaTIrBR06hHnkEKgJKdDT1I2rOz
nvZo2yaqpJmsuW0i/iK66XJzkweqia9X5hENCYZSjMksUjQGwhg6QE6D14cFwqi8
lveu19ihgY/Q2dvzaWDr2LnH4YoLgLHivar6G61P1vmzD31EPmN2HslQrLLhWdMR
KQg5WIrTUrqDZEJwAsV3Przd2miOiJ1dLh6qivm/iniuUzykP8ybRYYD4v56RreN
qxI8N2fGBdYj7KDAgOqtUAViGZdLC8SRzgkO5PpCOqb9aBI9Ke3mLxUnqmTDPR07
UrQc656Ovcso8GAWjwdhoZqkl75zhany2RI6tpiouge3gKVYOUq07V/JMzV8N9kQ
m/AUMgn6SiAA4xb1UqRVcg2Xx1Tu2vCGEFJ0D6uHvC+yIoeRzKUxsaTaivdvQArF
CVIc8ZOrIw2s6Pqx9CMeI1G+MCcGytBwy+4Lx8V76Nuav0ZA8ZhXpdYS7eaLHvt2
1+02Fyalt1ggDYnhSgBJYbUqsu4SDLxknp/H+d5qC+5R0PVNdlOWo9shhjkrXU92
qfZ8yatNyQgE6WnWFQCUOuDX1vv1dehT2yGkLiv/WwEfJuI4Wi72qz/yaVq/Ok1S
cPt+34M7QrkzLNVnQMa4tQH4Td7+OZyiFmGjDHx7nZ/Ext/dNGuyGrPSH9InEEwD
voObsKBzof9SCLjIPrmjNvn5bJwiX7oKd3PNnT2UCw2bbRjf2lHmkvP/METpPkse
JdoM26T8ycnQTEZNyeJWcjufT9aq9Y98cDq1jKBWaMTh11Up23dOXUTbgO5B27PA
kTDt1e5uTAgeInocY6UKL58EB5a+w0+IizDo8U84ti1/ATOwANdCqIeYh19R4ofK
Y1DMQmZ4Xj9StyJotwX79ZXJ+FSShqutRcrNgaaQr3KmanlWzyELROKK5hZDPDjp
rUffdMQ6Xf15qfhU3o5PVz/oPiCdZMXGrwpWUxP01cXfqs1GA3/JqwyjdtluPZZ3
4iGti4RHtXkAYtpqJU8cEPDxo0gPXX2JLWfrIyPJHajeAkj+LYW2QYbDGR1SwOsa
javPZKG0mUBssas2aNdWOTvZDdqvDYUDjJgegAlBP2Aya63NsLC98tk4HGB8irCh
B3YSaMWzvy3j7krBPGBWkb8xjrGK2/iJYjgJmisE4kcV/usnoOO3guNV/mynTKDl
T61i57+TKwcjj5LcY/WB3QcktZgycddfSlNNR8koccht9dW87QW+MSL856pgxUGp
vnisJhDgJbyESivbyEDRy11dA/0FG8wmb68lAYXN4arV6Qz1GH+u/3UPQZB3Adbe
JUCjt56h79TU7zvwWRvU8yXD5lvef+llnbzTk+WFa7S6giTzA5kdfuxxVOWsSLE0
w9Wao4nVOx4GRvFoPkI0XRQCDixkBa4t6jBX/OGy4OYXoWcCB/rjSCX7yw6EVObU
Evtu1qbdWLTqMKQJaETGFyj/s0k7AW+hyArkWz9MQzeh6Atg/Y7FenqSDczy6TWT
ksl1xMtLmLI96iLmmpwMuasw+goWr2+a7EPrCI+O1nhOYxe+U/Yku7k1MiM/z7cm
1R7hBI2PDTiwI8H+3CaUUNNG1tcXl48H7HOBo6rvnzCx1qUXc0sN0vSuJaaKfaWt
3nK9XR06k66FiSLQ+tf8lix+ekmcej8PqTCYc1hTXwL0016Y0HPR+TEkAkgvw4jp
R+d+9rdUIPLmlqoM+hvUw9iqYJ2q35MtiacGPHxUU641ORXaP4Br5z1TVQOnH7ru
t6Wl4krULVAe7H4M40Cqohzsc9s4QjwzLBovqjB/OvUqbkYRtAVVMraYT8ig2t5U
YOxGFrPcg4Ph5uNFIqtrzVLHLY+hKY0cfamaXusDWzSHW+TWAWHVt5Y17XmgvwCk
+MZun+DijoILKu8rDtk55udfM4FpQIQl8HlYSc7++hBaQusc+1CbxBCbsVZhQJjT
tKcUH2I3fBHI+vapjGfODKg38+a75QwYdKZ3GnKPDJe1QsZIAVNVY5PmeEbLt9Gk
cx9BAh4Cymac8C6swGj1rWF+VhZ2f87vSExliun/zs8PZOHlrw9TszDX47ge0vBh
cDweytU33SanWQ4+PaTRmnUTjJr+QiA8APeWCDOqfl6Ku+lvPaCvXuj3bQiOCRFG
0Z8NPHP4MaDqyYAB/BtxfaEK+hEYTROX3MthxlN8sy7ITw5VNd7yqAK4YcgoSxIJ
M7JzZDL8t2Vt2/O+AiI6xHc60W2GzMxE9L4AzuWtFC3wLoD9HlL02GUhkS8UoAoH
ZkIH2sfQW4VBYEbVU1RVo6HT+JhDPLTmLvlZ+HP2HC/V18aHhAiYOtsE1rA9mIf3
HRXMDBQVasakDyVFsUINVP+KKw0PVAmB+CWfhEb7GjvJBrrM3HMylPtSV5Gm8YnA
lBxH/PT47UVlTDI0XrmuIUBwkOe7+gS6VgBNK/feIR7Hn8K1YRzuj3a4DSb5xIc8
5MDIRtrOlOO6veh0AOH2bNrHmn2jqwzMWb6O8SODY/3gpD/oQSWtKFrDceq1Z+FG
tvzdLYywAZajxw9Hp7Gjj58A5KhT403OdmVqp4Pt4hWoW0abIik0VhznywHQ8ggf
J3Y+eeueUX4wV1UVH3x1asZCi7eztjmn6UU5AjZMs7giYr2N8p6odQHFehx16Urz
8KQ+JEzmPAJnzoaMct6X2UP/K7YcfZ9L1DLzZYvuGboQCtuS7J82H0sMIpD6VKsl
OhcYrdaoiu5uzqMpN16wceCWq8xLFMoe9izuO8Pu76tnIsrqmQSJ0eZJu9X28NIx
7nZm9pv94sMD2znxoB2fwLvBsxdr/823fIuA/jleMQg8YsFX17txy3ZhKqCYUC4t
pnS7uL7Odh15sJ3Ml47vJFxYOTQpOjNfFxAizDZa8oD/1VsZsnxEwvRZYwPZIsJd
MzX6gU2G6WY9WwZ5pRVKHqJuo1h2iBVZld50H6Z/psr5Ww3hSasmiv9ILWa0Br1Z
r6Qa/YFhFOnyIMfJy0QVkmJLXjmsmOQftE96y2gsEojq9i8Oys4/B6SkU/Fdm8M6
Ol63/nDw2EAT7t6pu2mVbFq1lVK80M7Czevj6kjlUVLjyU3K7NqT7x1zlzZ9+lH3
d5EK9XupI+4qFNIelHzQQA2zDdMSi5cbhCi43IUIj8q9isXLGGjStaZd0JD3YaRC
SDnbrmJfsLu6bw+kWJ1xgTuwdNm2PTKX8LfSI9VJ2cbSBjRKBcYD2RTeVXrmGaGG
zRKbXjzCdBoiz18hYz/YHGBhJmZodq5Ok8laOJ1+x5SDnUm4HiKC7gBttJmmnGmB
/Zuc1gP1iCK8asZZXhxHg4Rn3jB4rX4d9y87FppxWEHZQvHaIWCKlxUIERvrrAei
37gYVPJzC0Ps62c8gTugKlB2QAMYMABdB4RuzxFXakYTSBndSb2i7F+ga58Zq/NL
0em97GA/csbpqQBSnI54scpzoLC25mTqM6U0y3nS/A9pocSvJCjyr2KFlR5o6jwE
mK37rPR4zdLY45wNfIwPy69VmOU23As+udG/A5xXcMYIRsqP3VSr9amRQDDLm2LH
+6eCY/oMxShQKiPLwElpk5265ZgtA2hjggWx96TK0boPDlGBYqt+TV1Z7c1DpBTX
jN22v6dm0k+fR1cI53kWi395A0ognIXYnDkn866nAmbgSAEvJsSiXit38ynifd7T
V3Yx5hChqLWmEElIkdcYbq8CkCVZPJHjzpFnjp3cVOgXn2wnI/z7eGyesKkdBZ0G
fK2iNHlfImpUwFCJptHTNJ5rECA8V4Ek/y/XZwH3n3zE5+Y/rphdkY0P4DP4o7du
qBqDZCkgOLVxlpg6QYC7E5WQmlsb/BkNMI7Gd4ZSmrWoH9VHj3yyxYMK0+WrvNnN
BisReBnZRQgh/O6c1SUdmlHDsw7do821yg9c+OMzeMSBISehsCCk8mS+qXE718CO
fKvlQ+9/GJkKUe+cHyQ8w29mRUfWlRvOt7AtysdtPLVoQy6cUDole2M6AQ3L4yY7
P8LgEaFeCB4+RBlaY/4ot3NHgX+zWjGBlXv8fPRzZlCUm6eWnVnQX2/IGnSAzh+d
HTdYOYrMBcgDgCf0cvn7hPO+x7vlUUsWBchzT4Y4w1JtE2+uIvGnszykKEMJMx43
qd3OX/XDAZD7CY2R+CUQI1K2EdZbSMo3Hw2seIlQ4/Eh0UkmLnXV50Do292rQ8uR
ZdWsAYtcnJje0nOymww4wEHXf/nBitjQ2dyFv6ufGTcHun6aRVMsH8OU9d643rS0
SxiVtu3F8yev7XXdKqhuXX9558V8Isgo8P7HqUNGS9g8LlLTw9Vb2wlxF1RcJMIG
3qIe4Xlb/ZOZ08wX0VR+kMyHNJ70fxbjHf7QiUU6BO1/o6b9R675AXLcjqP1TkEA
e46Hh+D+NwlyjVdxlrWBomkCCh8sX3EEsWMaujE7aCMGye9rfjSTEUGvGvNW6azH
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SZrLBoceEAc8r7GLb6EUVgrbA3foGdueiYupPevIo7xqPSKDb0dU7HVUhn23Fovc
R1FIvxgZ+Wxo/A4OqQ89pzsFfIDdHoTiwaq6nB8thhofTNMO/LIx/bYRCEx5hH/v
thl7e0Iehjh9P+O+b759ENrxQIk4dVXjwBsDFx4ma8ZtNFirWfRnVJ42fvR1QK2K
hF0eZQ6Riv9hX1uOzZEQVgBc0OizWeaEFCGhp56fpT3hePUiedmdD6oNl/rOCcVw
x6gqVsCX/tjzQoExyV8LknHToMxPsD/fu+W3UBozUQB7y3LMFUSdEhhD7GAPKJED
shPyB/0F1RVlj+vV4pLWSw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7520 )
`pragma protect data_block
KK8Dc5C8xMr5DklRkHlMhi79ik4V1NF5iAUpL72E9ncG87kyV+BmWNDLg1dOL+4n
dEp7bHqZxAHNuXpGG/5pxfX6RZHziNwVRbJDhN2tqcWL3OFFhpY9geNPGRBjl5M5
5UlpDcod7XgISsHwukNDdDag/yW0I1JW1CZkRFg711Yb8Gw1Q7iEQlZtA2zatao6
HcW9gsnK1zHZ1MMyskZC8VUUDf5r/HjLviuow1vh5nJuav9f7wwUkURrhhof03ia
qMCurEZ+h5KsugIqg6owypISwyrCyJ0lpTXQPS8dd/FVunkRejYhyqJG3cDyetWj
rmgUnZWa+Tk49LevXjOf1R8PDlgyPsosNBhrtPjktvB+aqZ5V+6topT76uYZcQfK
9Us/cRWbVyUYWKFobSgvZ8/Vpsj+07yIGwT5bvZU+n9zABbSARGK2Zt00aSJvTSd
AU0b2iGU8HAxPeqGNMGELt2+T+fKWmXd5wpI4/OR4QDTqQdYfFmT+1WO5H/+NWhI
y3i/9ef4o9DyOmbub0n972XxIjZmZXRlKCXkzm/NeKH5y+UDckslm+pZBSTRwVR4
XpMKOrbFS+W9+oCYO28g7QAnxTurfgJ1gu4ln0ZCMC7zyo7z334uK66SU4xwN/Yw
SYN4rWImsFFeVY9cyFpN/emg30pdB181YBXCNh1XyK/26zyKMX62hWVFCmdbpXk+
ot5U+PlDFYxLf30CuUQ3NLmoCHDmFA+/FCYZ1pC4oAEh4fnPIkqZpIiMkWYKGs0G
9d9ywlQGSEyWC1DIzxKZyUILGg/R1Ghc9E01OSAyqzeUbdXgDlIpVMjXvUlO7Qms
Md9m3q/8rZTFVQrU1FYtamRN0fREJQlx8lxqTzMO+Izi2hG+4l9w76ttLK/2Myv/
doQIaYNQnAbohZZHPdqGPxRNpqFOwY5bRfUW+i8Z30hN6PrrDpCYJ7Wc1EHwIgUZ
gG6xCvHLFXwDvKoylsCFka8kYf5H+lWnLuL5wukNSrhPmKMPRmCJuSgLzB+5Svs/
ozvpAbAEWaYTjQZ1ariOeNPt57A/CYUgHZfvyaBpe2Lit66lGtnUSGlChileeFhC
FXF1Q74XwF3CBoOfa04vjkTzbaO8VSOb7JGJKTB7MnIn/kDrKof16deyaICGzqbW
W+rjTDq2eeApqDmVH4Q4gTVu/wojKU3OpxbJBruysENzMHA7A95y1F3kRCm/jEPn
I9aL+GvPMcNOcilFBoA2hCbYpOj4vqrVVKVx6n4TA7BTAhmLYUuEVXhAn2Gbx6pn
DLWziCDec97J34KybwRxpK8mT48m+35CeLd0QrIBwvgdOZC/akHwN3MBTxr3KwdQ
trmWPtaIQxuEI3lvhvuqIklJ+VAIzEHehv0rLHi5klZDFWyVDqFIxwA5IFVvhOLU
jQ1f20vQU+/HcG2sAK+UXoS0f1KIj7e9RzK4S3s1DskCNuhWdO6kr3jaHT1XuaVR
W2cJdEB7viswJASCRixsYvmhsFi0h9ihTY+r7iJIhhGyylqO1AoD6xxbkOOR9TtI
EViqkdX7BYN7wrRHnFmvhtXN5OYygIkAmLX8vPQSoZGZfdFXnXDcv8IujVyYj+e4
O+YVvI28T6wVhoXm70RIAKN3V5GO+VR/yYCDOeikmFpk0KOwPT/01nV43EbiZBcK
f9wBFC4DyPPyvb2AgapmjMsTV+JuGrAG45UmUH4FrsGgKWpmv/6lOvjJBOcsY6MH
mpF8sehkuJoeO+mednV+X9uS3O4tQA8EpooNe3sMhZF5AbpWIq+M9X2eEu2vs14s
iU5QF3K8ef2i1OxMLx7eRtvyUJe/X1wp0+eqOR6pLrCvUZx8dwcw0Ux9SFZHNQUQ
c3uwAE6ih5v/BK+97svA1nAOWw7TUB1opZ+qV+tcLws/JXEdlk3gs9GWhRkKwofp
5mbR7GrX7ddul7cfssD2nhHMdgQ2Nz20am0UvPfc7O3M4MHA08m/Lzx2cMz2Bgq+
o6eMh8dAamum01IBSOp0oHO5BVVVQqR9OZ11r6tySn7h7td96PoOzcZVu4aenrQy
0Q1mSXiDwNUeeaGyMq1fUcwNr6eU5s7WALO8HvJzKxVU6BjXdtdVVMpmh2u2UxGI
692GQqD/8HiokQoqHSfmpAgIT34CH9LHFEmzV3pcsepuBJupCLvmxwQ5TvK1ayKN
UaF3xNglHGzU6qMSyfpWJsM745z5oERcqw3z2xd5ccOKbm6ROiW8PO+VvUPE1OVR
7WlXB+QK3SFpMu/xqAGeOg45R491pXdP5bIBbmRENdeM0J9XK+hu+uBIHBmFhe5L
ZR8+D/eW8rlYrWc0CUESyXug4N/3cHdVnZkTfvN0yTalj8iNwjKOu/439vXCei9s
hdydhWBlFvSFHdHQOWmFmu9kt75de2E4zBxu9EVizWToryjxh/Dw75UVcW1H1rS6
XK9zimmfEUUFIIJ7SSTMd/t368R6uBNWE6OYVxCWLbb5mx4X7adF2WYJv/tlrLyq
zhAmw/gGY/lHApkZ3+p3ZyOwRvFLV1M5ZWKBf5NGxIWyUawJQ+gJG4ZF3aFyId2l
pGFFoQnCS7b8ro8ON9WbOzVdAVXJAOoLdlySykXzrNm1hgjbhyRHt1/RI7lwYqE5
s/790AiQ3eHJ+nAnzo2QnD0L2bj3AoqGR46LYjavKifGrIV/Hq8W64Ra3EF2r4qF
M0iVbJZr8r62zzUltGRxUxhPzSltuK3mX1+3j1/50behBZZ7mBntOiBvaFwOgrRu
y/u7bdPo5CrtwP3tohHjky4X9HmEak4rcruBuyBR3nHtDSJ6xL/IbsmO3ZlKwbNi
h6K1NGXJ3xf3JRWUqTKHxaQ/46jEr9u9YNcj8BwWKvCfPRYAapV/xCHicHfOs3UY
Xxj1XHCIMWZ3021S08h+KEePMOTvR0V6bnlKN4U4phV0hsSSdFJY6QHPhTevbMJ8
1OK9XOvKkPKGuJmyplz3/57aEsQtk/F5UUKWYMRMDiOjQZP7SYnnSL2QeCvjvAn8
u8SjXEab973LPoRIAhIJ6sHWwQFkcBcAujVssTOH9l5VewN1hQNoajnkfb+uUWU5
dkGP4oWfeWZVzxHSLwZmFTlNrmZ+HBUMRVnS6v6WqI+lfo718aCPiDXX8ziRyZqt
c7jK0lFVnKmiNovam4buqbON+pZTwZ1l6yv5m/p6ufWXdEwJoueZUqjK8pR7yv/+
PRX+Dd0+p8K4sDiCiLwGxhaID8T96hn84fP98xALutg9fgRmVk76x7yZ6zrX1FMu
oHveKmXjLIwj2yvgd4wRQTbJ8OLm/PMzZOSa05b16HZTcaSTUb0dsHQ96rofzeo4
SI10u04+hjKen1Vml45EreTVJ9R427Rd49OBrdIkgRw3MasjRCw433PcpjuNLZSs
qSaCEtT0+AufuRksM7/NHtjnurA/3Uxxy00Sjkut1pnujGkvsvCNCkjt174SHuZc
ms0gCv9jUc2/T0vofS0Y/Odqgm052wK/fd73Mxg7FAGaedHopWchu9o3OfJMX2u9
8a/mIX2CKT4NmlPgTdUGxWELfSIV0nBO1nKjVUnbLC7Yk17/DxYyEpEL1TA6rNl3
IqAgeY9aKinybPdga4mxRY79ehP/aePKS+u2eUM5pab7xasJ2TsNtJtQ+RPOFeDs
iSZ/Y27fe8A9RHmvpTk/VolHyxdTF059yc3kbYbqZsxTC9o9S91loVx/VS9OfNWM
/Iv9SXwRsezzpMeDHfpoZSHXWakZXaJtDHuKiQd5U2bXVbG9axocsFoWIK9VY93r
jlsfmbbfoMV5gf0I2FobO73bvnjq6JDrac/Jtjvip00V/WV0Z+4Km2qP4+4gkQOH
tUtkMRaGV45cqCTidN9tbdQAP+SFdlcUCnZaURKVsYeobi2WO//Q9dSrXuclLy8e
VaB9tDATwbcmPAzNj0b8Xpe58UaycjB/OLYb6t8QNpdmBkgKVD+8ULWAH/qN3Du3
d/j0aK13Z0K6fucyJgMlW2pAZEsvBvlIxKQv6on87IB+LrIWJraqHGGikqKyYYph
ehD/go6MdnXDKuT/azNXobeggrQvPZgKAPz4UwXwipaofS3illsaRu9ixer3GBv2
20zA5xLebKLgI3wx5/b66S6bnjWBKz89undVlz+c1JWgcxB9muAQscXN4Vf7Aaam
75ZCEr8qXSMWN+N3mwdx/BdYAdN2E8dIlCdyqGgdysmxcno6RiEBKX8qnETv7L4v
e3cl+MHk9FPHru5qgOjwYlER+ivdFmUl3weAZXxMVrrQ7hU1Pn6wcGKEKoiPXWGn
Fs2ENCk/DH2E8g4Qju1M6ZsdWCQmwa7rKG4yDRUomUpDlekc0/eKQRr1osG0xKfO
zRow2efszMyy7T9hIPtglcPC1QMYauNPVIUs0xHhxOyUAwS3LPjpeEjS7Ko/ztl9
FipCW14EsJfrGNmVzyLfCZmCt8KaA7UtUUVNebUP0rX0EdChvHW508lRH2d5SdvF
quBVrqLmeb2OsKaV7OTpXNpHKG6Oy4iZmrOWJa0c6+wqkIvugSuv6dmhtkp8db5c
JP9Mt3bS9kBj1l+eWBJLiYIVBKCXasaGYB97ZI0Cuss1NdkpJ95L7prmfbfszQTc
S0qqzEnbQ5SKKSKr81mo8hNTSAIfzs4Fmz7udSy1+h4wlA9zizHpqCd1sNjxNd/m
YClhDcj3yLazfqP20GEu9eG4MF2C4Eo3giactG87syKaLQL5qFBWvy1lqlTVXEiW
4q9otmsk3kf7ShVMHVqg4FhDRMhK8xTOYhe2msuN2jdPeIL7vRiporadWZhi2vXG
WcvjkIjRTxLGTvHh13QztR39IiXr34BNMHYcCdcXFiNPkAHcYWufhM5TMrGr8ys4
S6/pWHYkn1q4WYjgDZ+9CW1FWKrWRbFB0GHEdxoTFvHqZjst/c9lxAo5sf6xy6oo
V9kJofdnZdzK72b+w9OAtM3Somg5sp5O/UJysjbTxVhVnjqwTbrWsd5r0bOp7xst
0XGvoW3qEVIzYFobqbw2n7QHo/k+caSAEQCERxH5eLf1PXa6l7kNvr1206RS/s3u
N/WtxElNKCJRaWj1K3LWpHiiGUde1sXKDNOU3XhMTfkq4XNYuuxeUNP9QCSb+wBZ
9uNSf6h4ZD/tZzfOqPjEMAj3kCvMXxgEredjFnkorHG6lBz9LqQJaiOvqerE09+P
y2Kc7zPWP4G1FiefImbdMnF20JrkLeVQ0mvHe9NwgVZrcfXBI4EsnE8Ej2r8Rhst
FFdHq6XzxIFTZhboaklp4JQMrTnc8dfGoD52xSnWIKl23jluv0Rn8TlBk7kTCzdL
v2YmQzAopqurFo8rG3DE6fXTraa+8tBvnCypfCYn49AMYVDufRt4Jz2QFbQj7zX8
HabJKmcGvmJO09Bf6BtYeYbF4YkLt8cJBAt65VVAgs2cuwqilM2lCrC8f6UVkfyN
jxzdkTbxS6qvxMK7J4JHepgeuwCMt8RUzFUjEjvoOH45zZPDJGWbHXwYqqwA9861
9OVgvly9pFvsPrV/THx9Kk/5GdMbmKSXiJEUvSZA/rcGp7vuDoB9pQhnzjzoa5ej
/nbnDiv3OD4XYMCP3Fgm/JH3vKoTtDqtQgw+KVJtYeW2FIQ1poNfaltBusch4CnN
bvZ8/BO/bZjYz2l087oFIqFvaMfvPLqP1bg2pVg/HxPdiDtE73IWxmTLNykBx6Vn
9CMEAhLuOMQw4cGn6IsdZLegFgAPXPh+wDM10Ro/2ODLz457XUUjoExv6k9hvxJR
nkRk84IiwGlxmH/sqYcyUTbtnrjRItVSgAV5rLAmUaqRfBD/YfxNR97+USFVQVPw
t2ajQOeNebnmwpbllDDDSuFyqKgX12vfbjS0k1+aw8uZh8pp+EJWXzJf1fTWGOOb
QJNnr8/YM9r2NXMnDBARYu5vEFvR5NGOnyG9V2a7c2Sti9J6h/JZaMNVXken3ERP
xN6AIe17G1UPKrOeQHTD/vdcmz1d/P152lHWjscZ62SGUgmM95Ibp5+ehyjxgreI
p8VoNd/b2lzBPLzAjuQ1bRsFyfNxIFZRKEhBkf+GGVOcPlcMihHG1xyjfSA3v+C3
Eb4QOzxx8M2g0NJe4TWZNeRqvdcyQTYPNqZvAUYFhlAJ5i4Ie8316dx3eTCb7scv
H2XZqr9JFgC3zPWNNZ/NxHHxVpKqWV/7Ejs9Kgp5kakgiyRPuqyga1UAMbx4Vq6p
7u+7gDXbbWOCRylNgV0Qapk1smzn1LtqYtTqYZaYDBvKW0EbC8sP3U2eFDuL9DGL
ZY2/gp26ku/eblww8huyk4wy925+DwinUzwbSoQM1XC0OPCULLJWX9savZkkBIMw
d36ZIU2oAVjYTT51GwcdF8yL/YfCYvagL/KoVJvv6u5YOeuiEdGOSTD10YMNfD0k
PIQJMur5QZ4J9xwOeZiItfFERYlrYoEBHD3QhjQkHAq3MjcmLFAV8Xgumn5Q5N1C
fhVaKxajnQtG0F6Zj1aMSGVjetp+6lYvRYmgMfovIQT/DyMLUUOpSto2i7dUy/2g
f5ws1zfDS9Yu4pM1dxWiJOcL23JSlcCL9p3+nuFyi8wzhVaEuBNUau8vC3UoIfdT
HCPFS3WYYFZEtIythvvIOZzsGcSkDQDk9eYNVvtBk1Rt768sQ5090GPR5ZukmPIa
KM0kbOcsoW0ERbxMSq0R6wKKWJrLI1UqxcUZFANyIU8zygkikQNr3F67DqJosVFM
0kUtQMIb+KjAyVBOdLNsKncbyBllpdejy8YE+jBn6e9iHmW6w7dXizwe/tCsXd3y
h3xr8QjgWGZxd3HDlLiJkN8hFpAXWsgjQqHDtTC/MSI1TAkT7xworr6Nv9Lk/+dv
claVPtEDl9s7a6MLkR9WSqJkhgynHEAHPtQxPwpwNTmjOz5Z7pikCI2JPJVGrlHO
cm+DkaTQ9sh3C/xlxPvZ7THq9O2wUESQFHeulcap2d3sDMaG8p+o0FnJ8bloVTVa
szdpXNuqZgujGOUhpsZIreZGhjMCn1tmfAimCpTVgcU23/M3lv0B/U94raz6o/qB
JZb/wL+DlAMIk3RIMkPxDm5d4CcrYsl3hs3rN0nleRQNFyGDfQg6bVPRsq1yD5n1
AOi6TcVwHIGf1GjlhmGHjM8rb3oLFQPBvtyM1KNf22qZud3C8zpbDG8M2uTPUy9R
qqOEVeEm2qfhp4BgBFfIKSgvZTCemTU1osFYRaDjSYkTGfPiGUGCGecj+Kjblc6X
drd4kAJOgglojaLQTKZpt+5yCBTzX4/rn7mtn50pYHHhiUUe2AFpu6M1k7EugahS
rru+U7JdKjatL+OrgKDK8xbEMNmsiMl0zJajOQ5Bjr8ujQpTpGmujYAyduG6aZbR
zJsJdm9gWRsEyXbJA9zaNxzuugHagF9Uqmo8je/rlupwfr7A4ul/Dr9ulgD66cyP
ZqsP9yRtYW+CfsmcdgQva+RFlhJCzfizBw7Lcop5sZ1P2WTNnKPfL9C0N/MqEVL6
MqUncYuiYPjqjrdcP1toVuk6y8tCO72Rt98sXoSnJfTQzFgsv+ngiI14M+3wljfj
XBCfGAxXvyHUThbhollcOWeEDYTwLjAVbklyGhB49bSBRNUkb0hiPV5Ef56Ih9es
YryT1V1k6LFUCIxXzgnocMgVc7RGhXsUm21oE8AAPIMRfyFTorlRXccw8XMxTOPt
MHOmaB3/DtW0OfL6mrkqkxgpg5YXKWZ6oqiBOoYMGZaYlgYkso7BlA8vdNOJN1Xb
ij+Qg0Ay9txcFX5hDprR8egonEL5VrZUEuRBAGAi8xkyLu8rfaMlJ7yHqzBO/vmR
l5Y6oBpUqVveW3Em4vzglp75qsXoF264m2Ao7LWTjRjMNJyVyJPFMZbglhDlpDih
WML2VHBGS1d4/M8TUIvCUWh3Mz7IWHMlsZ7RwV7sj238B7By43vJyd/q77N1X14Q
/i9njamzu86UPmIK0kjNefrKzCWcQ4Bu6bEDhMYhcBEl9AO9n9tpLdxnGXqCiKaG
Eofyfc1DJ04Ft58RpdsoQP8jYkgF9Ejqfh3VnHf+MqLNhSAbTlJae7iq1FZxib0i
HQ4nKBhdww32Ipp8Z7HrCh5+6uiTgn8bPLOnq1hcb07T/gZsnU2+3Z3c1tC/FLNo
uo17FPMeyG9vrxqaeCQM2AHv+u0zV2YGKx4yn2XVeU5og8duWFNqA0mOslE8PGRt
xX4AKW3h3YjpEQnhKKEQ4uaUFupWOc9zkLCtYwTk9GxNtOG1cpmRxpCFH+xUC0H0
EHjjiVnJ+f9PXJvUTLi6Qd269HEv0iT21OGHqOQ09hQzWyafLf6Yxosg+GOm2ppr
K5v2HjDctRR53Q3y+LOtIpeFKVANl39WCo43+1CC35HLaAhVVpThHSQ+K+q109tk
46dz7vWFuC+BmNt8veimPSdK1Mx43NoJgRuryv/oCNaV4I5ilg+cFF3Tflc5opSt
ZnrJKUQdKTKIwwJkyVpkMNkjbXRyklSEd+UQzgE+fNHRNZagfcbQB9lYdpyb5pZT
WnpXs0RwSnCN9aDL0KsTACH5fqBPVuqact8YBInqc1dL4dkvlduVMcDYmCSQn/tZ
CZxFmXgcTSFZMN94IuFofdQIhGtjQ0zab65kPEaiXUOSb0uJi3AvaXZilanyiBce
I+RhkVHLnUBFWOrbBIJFf81JT/7+5bisWMd+RxbrqKXezZXQ5PqMhHjK2RtP9t3e
CD+HANW924CKzJKT/88k14gQbXkFCs3abmviOx1f+5z4o1zVrCCaOlbHdTmJGx31
893RkW5Y4IMxVUVfU7UIuE7PPu+nCI44wG/5gnjBtO4Ka2Spbi5AbWRO2HMHaUZB
uaz9TznJjOd+hqb5N/R5urgHi5wvMGBKN5yw3JAoX0uCV/lBlKr7CTiyPtU5v4Li
M0zC/0PS42YSJ738he8tagHIWchNuaVcfd+a09XKIY+3NO0uCRyyq+6u3lLFX297
yzITmzv5ee3UtL7zCSXYeF3HaFCUKCT/k0h0IsWBYadQmbMLoDo6c1WQL/+0dpIJ
aU8PA9zXO0r8FdeuYEu3HW53fujQ3dhetSBT4y4I3opkHrOrOuqs2M6NPogGt0Jr
cjV9hwmgJfrxRm9RvsUx6H+2iDFYg9N83dz6JSqNOHCPZt1giRPqdvnItV//x0Rd
a9RjAtTbJIhhcGSKwsNijjOoqj9nrlcmOm6UjqQOYUDLwwyy59QctvmtfxpZ2OLF
J0Fl4qJqqErxjjupYu40MkSoA/SYxpdhN5mA+7SuAj3QMxbd0L0zNhCIWMod4DxK
0WhiIxzu4K40It3P+Ir9HjvbiI38eeQHwDViTFHzElWsy35Xs3lFN6IW7UCMnuSP
l5BI6852mS3DaNcEv4G7QzDJPT2dnzqHB/Q9pQnhYx8sKCbqIW/kp7cUBEaj+uvC
AASbOtpb2ALhYhs8QHh2V4nN+1qTeTXaEWTt/FeAXC1b6WU3Gn/WcfS98ULIDLCf
B/GspefKzc8Wt8rFGzi0yUmhHgCpDMUAkuaU4saqWqfyGa44AxVQhLYlLh487ddl
fB7mma0kw0x0MMqruxPVLVf5xWk5vveqEnoD/gR1meQwwNc0zIgf4d0LZ8jgXtvn
g4kvAQF/E23v0cDeAPEVyFwQu6VhaOaImWWw9SKS8RvKBC97Kt/Nf1hHsnzUcdFk
LrNlBgtyN293LD9a21NUAcMvhSODOX54yYJeTNX8Nija0zgEb/mgFCw7xR7DsNi0
Y8RWHVfJ2NGig8m6DA9buNSj/E88pzbiIkh8vxm2kEScJ3+4hobk48YVkYqI6da1
3DKMHtpjxjw1G9/6uCB1HEnO/KKk8F7chkWByJlfnUm2jIwhMBWi5QDp7wTdpy6j
ZTbocDzTSPXgYee2n8ViSrXJO72XUKXlLkPIpJUAvRid5DS4d11MXuMDnn8wAlZb
Iezd8213diG9HFOPtLdI2JgwzSs/AJ0LBeewz7UWv+mPjmI8D4c/tAmgPi+DnLhW
0lRGci2fmo4aqsoqNKTEBBK48LBgHLTVE3gbwBrMyH4=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gQOIMscy6YAoDrfi4cZjfzFKLRVEoJ4h5iXOz6BPfJhcvZX2yNL8EcuSYPGXPnFc
iwqUepFZPa6Jm2R7Yj7o9Ymw6aNT+CXaoVd9iGk0yV47DCf8CGq799WvUduH/lbr
X/SZPKt0eQlZhAF/PG+suqzyRgZ5HPAgdJ2a1N8S52KUaItvprwy9aOvmJdlWh+B
YcMsjvzlcCZKuvYLcEo2TbuUJv3YK5TtZp7TZ/8aR16QhBciLhhHKTwGwNMECIu7
QjVdbC02UsuPKahvwCvvp8MU2W3V2hKGJvnRb6gf+iFrRIlIL/dRwj+q3HevRv9q
mQRVMcp6LFMO+FSnhLrnZw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4192 )
`pragma protect data_block
i40UtXg/Hja+dZnYbbS7MyOxxACYsDOu0i8qB2xtYOvRpD/OCa8Uw8oKKjsGoFIK
uLZ4s6ACU3QohUzgcQ1+M9sqc4Lg43Cz6/YgcQ9ifH0DCbh0haZhhYt3MAD6bVYx
3CmJXsU20wFemskz6wV3arDSuPQOezvq7WMvWpsWM42rVMRCqKmgpfyTTQwJWED9
66gAIP0XkcFyoCLF6p6Sy6oDakr8Zi/QsfnR9r97vcFoIOdmuuoQrovS5CaKq6k7
zN4hClPz6DXNWC1CP4YOXCIXFzufGZoEeazzApi3W+oyZljjf1rkikn5MnjdrdXQ
PUZcR3rG3KxeOysQf4gJbg2SvsJJhVtoPBAXV8Kttgijfnn6VJka2S3ibpg/ONNa
BeQNsA/pTbMM4phCdWHNwqodlJjpR/levbJ9oEX9+2pi04ikHmCNUtaQy6K+GA9Q
il7869t45hJnAOOz+lbUlxKxHoG2TCj6VtaXQOgGKNnHOJSLleUpWsL6vMIA97mM
cS2RbjnXDp2O0EJyZWPy8tuTRQb67ngFt590UJ2VBrZor0TmE/5kvY/L02gLSjR8
jyfyB0WH+yMee4/NuObNnqVT5fNuF9xL3wVCo91jv+lJDh/P2HF8/y2wsurLfj39
H8uSYMSmR2Eadsb6adVsR4GpOclex4GfIzKhIaDSBDrOuZDOEq1eIsl5hmptPnTV
sdJ8+RPgpLi+EWFr4B1T9lJowu2tmevmNXC4CHxHpkP0kq6CTLuAQWRP6H9Zqj8P
knH4MRFGSTZ8YJeO/15D9x+dpApTbVxV362GtMzbxur+vfw1gFhrmxMnxM2b8uXv
nKd7lPUAaGeRaBSrfSt8xgi54nNlELoyFq0au2l62gxq01ag8/FdmKWzXuh6mXoA
/lW+kBlAlI0X7KhzacFVzdvZ00b56WW3kkNUUEDGlk2972XGFS801Rz4exLjou+5
xrsu/rIEU1YfE30jXN/j573xAnyz5GMgF1PUIb/fiLbrZE1uRltMO/npgmf37Tvt
0ajWG1R3ezNPh1pBJAhm2srkpMlLDJbVXnyTad+Ylk+u9j3bH/DqczSug1ui/QIM
/ZdboNXT03kXuySvzVrWjZ2VBQgyjfsh59wX4eNPigm5NzBvlY3BNoDnaSTeIlei
tSfGGeS2JljFzTQ6dkemb8JF0CBcqMOIyIBIy26i4qIifZdaP9G1EiYQeeu9ASbT
uuJtRzHc/brVcu6ENuL/e5WH4wC/a07hnWaCbS3Mbd8W0+mShEj/HnDi463Eoduu
LK9Z0InYxCJ4Ib8NUCbM8WA2kg3+0ULpHY39f1sIJE03XxHslXQISijc6KdbIpy/
AnAVzd6S8szgu+kM7SSWwpKdnJeIyi59mkckx4VlCy9j3pznS6se0tzz0gdCCPw1
OYiYJSmunQQenzI2aUNel9pFnBgGIBOXlDWWKjSN9TlF0RY7Iyii06FrVw/mpBnB
2IBn7u/2CRVcdVS5l4J6G2AD4JZLQDBjxkvtj0zg5dkZwA43PcqzZ4v9m9XpXqs/
AJIgl8UngMhhIyGiqgG3GNd5ZG4xKQfLzuWh914B3R7UDa0TXPpF2vKl6SxMV2CM
YgEEUZcEXrQYk7S3VybV5zdHm8RDzJHOEcFcvmV81CPGmaeGFQvhU/UYCa6Lhhcm
2Osl0cnIgIlM99ulMTI5vgo8EMpK8sy3rSLOk5VDsEluXN0NW8DJNh9NonE2WPIN
RiH/Jj68/6yA9FeNt4uHL2KTRts/uqKiVGkuRthxwrTUlDgTwRzLZ6G09YRB4qUM
1oXih1MCc9jcAuA2tzyI+0tuxRvuqwpTj3vmdvfgNsyCWmCVduWW2d14RSFx/1dK
8rmGOujV0jsbOkOYhYlsQXYAFDAx2rIQoOZpL5pUKUxyjoz97NyUMasvCtqLSdPL
Lu6zHk1JMoU5VmtqyDOd3+HKEyiSokeXu4iavelmZmDo/WHUKLgQqc8nTCEAtzHN
wck+8YGAX4ZG0Ezkx6DvOq73wYwUFRgW0/QJbljgAyYb4hA1bxwy32jF3WMWv8p7
47ngz7fIJIozTjv27nxebJoSb+Vulic/vn4QiNULMlMJOEOIdixqDQcLkGoJGQq4
mNz18fwtANmwHkjQmu4mWLcmuw76OXH/KMok74IOM/8jAgKwSwlFx4zrX/PTembU
Ml9Qj7hMdD7SKzRwWt+VTBJgdJ+8XlL64DJANZbjohlMG8TnlGHfOsirzK8BW6ci
lNHphEmt5Sgv/o6QWuL2QvANdUcHZ7KiqfhFvRb7oQi8Xd0rI0bCO5ZF+L9x3QAo
pBKpFPSUDxtXSQVwquYzY3mvG3sxEPGTNj727xo6g+0273U/ZDQnXRKyzw5bl+Es
lem/h9IN8vbEP001CkorUm+y9Ouagrfx0XJkSY1nrMp+pQ8kpt69KOPyE/PhHctF
mePTQAyQ2A3P/EQh6z7qYbu8MLV+kc7EmaKb+D29LdfMXs5WiJPfyn2z9HWikP48
rsn0K3KVyUUUV63AqHNkQaq0rMsB02RjEdMzVLAgRynS8v4Q4Ju6Ui+MOrrYachS
o/aSk8ozgNTjsAM30QN0Qu8Mn/vp3E1I/+sdFM6I1RzJ9pLChPi/A/RKtr7FVP3F
QzoPq6q0gAmnfRJuIBJalqYzZQtOvS6k4+qcnM92lnDc57uoniZn7lMZgsIYQfKS
+MO9FnUUtwl/a6daPWt14Ako3GVF9oLkotbvCyV67sBGHkoJGuuwZAwmybnk1Pb+
35j6/GrBadlXpKG9kUG90e33qfPHIC8lt/SGiku0d96NS5ZV++XEKy2NYCQ8uxj9
hpFAhhdwhdBaVMs5cN5U5NKEH8N04yVV9K7n5BqNooxFXvyfTCTNeWwpmG7AnJNh
2hzHGgZa3XHsTXqXg8IdwVAlDi2i+AxD5nCPtGRGQxkvHcn3nReqGzxyPx3leGcC
za31fNy7eHt2W4LivrDvo3UkAel56DJQkvjjBaR/jTvoYdB/kolKifXirP30OJTg
lpP/2BSFZcn2Uv/3kp70JqLGtj81kp37NRnnP7C8JmArTTc4GoNu3rUwrbTbo1NE
ZQvpUSOmT2EIfnr+s/SIV4DBAyrtwGGNjdk2d9CE0yhMyx0L7LklEvt8s2btM6a2
8PpZz6LPZvcQ84csyFRSSlbFny5HJDRNQXv0/MV8Y0qAiF0dJZgAw3TdYc/P7z/A
TsSYhMPVV/S+kIF7i8IDo/WxwhrGTb6EEe4BO/+lQAegAWe4gvK0rPLI8EJgLoc0
c38aZP6Qvy7nssrMJHMuNOR3SnE4Xxgzu4hEFZMK0iwzeBNlmlihw5Sfy6Hpxaxn
4+NznHbSIgDV3jEn4K8pI8qEVAfSC+w4Cl5mRz4aGyHWGss3ayyB+h1b3WSBNx5D
FmQQbT7/Hel8t/SapaAudCDB5jhDMCj7QjTxxZN9L/05PFZLYY861eTM1+sMqfua
RE5jvXNZ5H3zvi2IzGK5pHlJ9EzelS1uNe2bIY/HtVirHpYc6ByHZGk2qk0at9Rf
rb8DjMYfNfOB169niIrDvmIDAxqcj0GxszSDH47D1uw9rp09UHfaIumf1606eLEf
gq79wSy6Kbv8j4tyhDoRMSakkLXPHU26298jNFsAV3HdJeZEETmC4zae6LMMTGnP
n0sct9rrVBXi7oGE6yRWOjtqliG1BunLSoXATpQbYBfz7ZMNXXPLoGoRZtRom0Zt
oB1scO2xlgta1UTEDNpLBjPhdeiZQhsHoYUXzV20NTReXqPrmgwxuIEqzAYUdKYu
iUN8RBuxqVeUuK/UP3A58S9PYOpseC2/E3Ew5P7VOPF9JxsjGixzqvKiiLNTqU7T
31Dafxlx3I0b4rkRNXPG5Kwb1+Xsg5NqZ8tCBh8rfyA7JfiVCEtdCvkqHiNR3msa
ao93I8HjQ/QjOrT7k3A82X6fUagRM/CRhkzsTiH/tv5s2zEzrw+H2PerflsFFuo7
aL77SMhX9wtsKfIkDAwW2WMfOOgZbjtDlTN0rn4+1d/QmeyZXG0360QuOG7vdM1k
2CEiYzzOuvRZ3e6WO3jrYBlesS6ezZopWzBBZd3Wwc5ktsEhOy5zkuNr1xUtd3QF
yzkYoi4RQtZdBPdbmvpETRa1X6Z97LPzNg5ctLV8j4cCGYX81J+vp0YDSKl+Fq/B
f+i7soJs2LgIx2c5kZGDrnjaB80nknMDXhqhYeOeIlzpCTfwWwLqvuTb8YRzNCLl
hdTB0EI4i5xXunByTaDycscS53Id1xrMPn7hOh4t+Hlr3TxqjjBD3mbFHcBXdfcD
G9ofj4CNYp6cjlDQhpHUxKJcGgV90ryQ8XFzJCkNx+JTh1Y7Z5rgp60PJZjImksC
jEz/chysKcown/3K7+UobCNJGUrcM2Aoa5g3c7Vwipw25JthfQrMfl3TsMkSyVS8
nFpZi2pwfgW6gPH8C12p8rjWzDdBTDfa0kLXUx0MSKvjswXftB9zBeEak8/k8bFW
D/MyP4jl548/7gSYh47+2CZ1bPQ3ptfRPWBAOS5SrHHS8yIpgrQs9XfzxyVH2uQI
hHcHgHSCgYeTa0EGZDUSClwB8ee4YNm9ySE8isM91HU4jcHSx5XLRKVDku/XIggk
ujtmCBpd/smxFXeMO1oSrZTJawWuq1S33fQplETrBOkUWFyBarVNNLfU16si6DpU
ifFuG8yV0bOfNdBV0Aua/v0589a0jh3a+sLwrFFwTAW+W2OGZBA9ezXNqNiR1dmO
z+a1yAU1s2BNNVxilH+VTRS+oMuPW8oBm5UmZ1H70mAed+gsSfFpvPVTSQ/hXo8d
BMxD0UditUGEAAUE/rO96oEb0fyoTCqRswFTlKeCNHh4VrcvWkdvimnOY6cunbrI
0NQeXIMJVVdQ1wi8eBnau4Uw59BuEXDsxgVOQLG/Xe6taJT4qi7ccf7lQ+5f2HX6
Gy5PVYvcgHrNHnrf8WCZ26VEquqQ71FQ+g/BFMh5q/rWZ13kCnlip5ci11oQe/jc
8ketnaVZx64ZGPGSb1folVMjcnvDFfdRb06X5+H5t7V/+Z1Qnf5phfFSswhkyIfA
qtmvl1tI3KO0zz2DgbRm8Fts6SPtC87c2AWFqFTFen0OJSISfhI8ZxMRwaP21s24
SSBLq5tm3LY1Bpy4dS1yvqYf30qdPpG3KKxG0thD3N6LTGCkvuKJGfabqQR1N4Tf
i3yOEOuEBUQi1/qskUC0+aTbVqhDWRUecUVNbp1xddr/42Yagn6NMXuvvi2yt++2
1bp0EXK0nsLPaB5DE538Q4xQoQqgOTdCI5xeDRdzLrWUamVBnmnRDJUVPVh64fdm
nzkppG2Fl7o7jl0K0XkpmULvhMSjoLn4KV6GGT7ELvGHKFlCSaTof+2Inx6k3XlH
eSH+ONJz2g1QW8HaF7zkLcNQJmozGflIDYchfWaxAJBSPLffiU3gmZHef0+nux+o
dHIVHjF6kYVAgkctPNslB0pcAWW9tulXma11yJb5uVwg5G69c19V2Mt4L+E2rGHr
hhPlx/qenRRrCuIyzDibqJn/GVbg6nLu3nv6SxbY3QhTim1NA2AbZgCU1ZwAhY3F
fZDkolzBqs5STCxXGjIr+g==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JxmOyl30ecuDGm0XR2P4xcu019FmKGoFugtjZq1hJykjYMrjACtQz/dfFGavVusa
kL/UKReufa8LiP6Zf8bHq0g5R/eysLMItx9IXxIVg3/d6sHfCO3RO83AyrTCCOAe
trqrfJXfi6WIxsSXH9jCfubWr8cTKJG2EB5VsIuxpQYWB0WAuj18Iwx43lzPD+MG
z6C2gmRCpQmonACukiojPGnFvOc79OrWTQgM57RdQnzYu5RSL52BjiOz0c8LkFUw
d2wCY3cU14tybPzr/W73jcbVRoxq0dE4sGwkXdewhsTWYIBYcoRoA+XGnEUvu1xl
rT5NvmO9lnMYIpddT6X7aQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
BLtgnsYaUzu+iA6+rdRwVPK9tUGfYTUBQbwdER5mlpjQe7I/L6gPugVLW2HSgOUg
TatTmol91T3SGRn+4yErLBVf8VqwpySFTNI9DCHFUl0KwjqzmnZUDq7qVJqa1ZJ7
MZXLUmpAKXqmXqxAEciLhYMjqrxylqih3ATIU2FO8mIAjVpGkFY5maEJ2ilo9c64
kw/YKJ8VaJNueOLOXq9T/NrzDoXspnliIKJLJDU73ZYXmdFAooGkkHs/B2mlIiqJ
Aa/VdZDw9sGouatcuMrF7iwdpB+ejdRa1cZXUEhcmjLzbEBgmcxvUqo/4j3bXhEF
BGOX9EeRJYLjV53jw7qW1dEsnsNZ/MmlcnCxy91uYk7LkRgYLuBoSfQc6zqJ+aej
pYZc79jm/hjG3FpMDFRX8Wo73EXAeFMxl/zYzoQ3XKPS80PxgluAsF7KGh4MrSVi
VkJNK8CfgX2CX5k57ncEAQUdPiuzzhg+5qOtz9lCszn+Q//QXHv+B8DN50pcyf/w
2Xs2WA/LT5fCfb2FAdleA/VpoRQKyhY9hdYB2G/mm5xHVwUJ4GXx0hQvcWAkkHFx
0K4c2Jwm5RKA6KBce/+7kiWwrl2V7n42sohsE6GKQOlgUA33k492+LeRyBZSlZXZ
74PjjiGD4tYYTfunrds+bIOHEdQSd36At/j6khg7eyZBG7eQ0m2zIjQdMzB5koxn
LSbeyiUok7G03q4douXifzR44TYbRbb95D4f2IND/puMJL4Xiz1zEUcxVTS8pqBX
FFGxsbHtHAOyPhtQdN6AR1Ts4ZBMZXjO0J7hY6HIBCGF56YsY3mEYVjzGn+y9VI7
peuRQdL7N+l4LG6UEdWPgvBbVg1vmIZbEbN8totPjE9wUsejeDN/bob+bm70zttw
K89G2bWv2CWYV9q+TevvoGCv6a8DALBXg+WDZM0TzRdIEQzg2VKpGNgi0g94o+uJ
MutZHfGo70r2aI5+ZtVpfjsNyVmi00DLSsxClwo0fYwd3E6xM86xPXcDv3XVs61C
7Ou/P9QzdyK/jTLXx0i6xhhOf2ioVFp5RY19DQfQHwj43BkI4jaNx9KKAncZ9lNp
IUWti8R/NAgAp/UfXJHdSbs00ttTZEjvYLhM5pG5/vt3gzhLP4nUNNQpnlOW37KN
/1vIuwtfkYOEdsqTcD02EL96xsmfHW4FIJyBKOw+XqzaB6tpCGfaQXaVwkiETw2p
kXG5rcX7MjE7RRYT+Pehdz39Zo+lkduf2/B4FcRJB/ysZsb1BZwGmuIKSyK4RXXb
3BSdXs930SBU58Zc8rTTVw848vM520RCUWGUpYhQ021RW/Mx2rWi7RhgHOFtEWBe
CnZqwO69x+XtSMErl0F3zI032EuLLuqXFUADuYcDQn9E/d8zlPLFbEdmufzwzBnx
yqLi2KLSgKw5xF7pT6rT2Q9f5lYzMLsCfFqIpDFLDhHzZ21Gt4vLqm5XzYdDEbD+
9Gkb97lnKjZHYceNqS0j4BkYbp5yl88kEU4fJbgJZVHwS8GoLsfk5gMd/KawHcg+
2VzaSHwCkvfAEosQqEvd+1Z1eYKbogxjZtjN0yFf+Nktd+W8COkdU4wKDDQClRqS
P1GqCtQVp7ebWYdI34QKpWf4IYeSVsXEE7QUTpaMDPuJ91yaex7g8O2VbMd7t7al
RXPhYPXpZ690Z0HyFaqz/LYBRH+KaCTbiWReIUeAgm0MmFdTbZbDBxDdt9V2bVQM
c0O2X02zVh+YHiIinQzYG0dVaiFPHWWO2p6nA0TafFsJaeCQ216QAQGJfgqVhyXf
lJ9GQnjO/gxhHqdyJir8Z5cwPCba8GWUQeTnil7nJZtcKRuukgAdzB3s0RssZ/xd
66QMKB0xgmum/TIw1kuy7FRMlH8G6LlJ2hk+4qNjVWD6i3i4ObEDUIjzPotoslVG
tbz186g1e5mEtXdPkn/UEEHFAbcI4agoi7oc0Lsn21INJWQt85hvOUfW6xhDUIbD
5qs8PjTQKmmLbLYPqoiYKIzB6hUiEnKlZJ7JEyypfG/gPBv1W7+tWXlaohXTKlAd
EvJEpNPSzg/9UynVASwMEg2hm01VHH8EhkGX+RUjFg6KlKKEoR6SJSG09RYDzOA1
FyDq6bqNKXajjO2JzVkUGCYuysS1VKLN05O1XwXQOuPGcmNTvknEqCvlFTyKtnch
CcQCUTdxlwQRWtgFx3L8uwiSNvFLt3Iwwx3qRSSmQV76iE0ewtov7umtUxmzFS88
YSs3gqXi28b2j7HfgvLHzL/hCHtsVNgCObLVuhBs16OQjb0VBgRb1fwxG2X1kfwC
qQ0x/BRYOD3mJxfbMON6BpFiNyYSbpADNU9rSrKHJaRisQy41ex0iTotKsytO4j1
G5K4CRh+gWHVW5/rRmtOGINP7fXe4b9CWBe0EEAp/w5UEYHVjnxnKQtY9myj0gbz
kBaeiMWfcEyDPzhZfKElKbzhJ7OH1iijd6AevFkDawgv80MJ+iUMnhq3U9hru7ZM
5F8oEGGXeXXIDCzgIrKUlhyOBn8PCpGRmTHOpzQeNmMVSN1Hl80O/+wxiUps+bl+
5s/OR8Hk7QuD+13CXrYxjeLieapeb0WTrhA4zE3f+BZeZ3HqQsnkkimoSwvTMls9
1WawzGFBogYcDv8RBV2wRVs5SjXMSo58fyqesSvEP9/bt/cDB/BpWR0iNfKBIlEY
Pons22COse4DJEHultTe3sM49J6t9QbKPaM8cIjbomutc9yDyfTZW6euibJIei5G
pP6a1bXmsOxK589KIWsbs/9gkS1ddNw9dEvGrgb44KlqpHHEuTA5dSRxOBi0pQ4A
njJxm3cgcorbvGMbPa0u+QCOv9czO+XBADLhx6BNeN3KQplvquriEH9p2lslHb/w
ptvVgXXB794r4JAOdZqAWR1GOD9D9w3LKeBYC/b0QeUcVOqkXjxTfPpqvLsJRU5/
iKd5yo8kUwWDfxL7O0ACUl8ElJ7ALC4ZZImvp6u9eIVcoHOYL5Gd73A6/sJA9bFV
dmkwAI+1A6kiRDmRRiMJTUEvXq+BGPstQEJ98icZypML9vjtSvgqqDvmI0y0piQv
STKjFUFCbyJNV5Z0sdHQFnuETrroC3BWfs19CbOMjC8ukvMu+cKsmS0NG5A2gDGL
7LSaznrnpRdoJep4ju9go4DCiE2E+2Iy2h+cl5gtswzvdVJAiV52zE7ZK7CJVAlx
nTqRCkogeDjhTikWlIYRS8dYk1SN9CJHe+0YgFLHW9c+eKivxVvMqGVjQeG2tnDM
1TBCLdlJIjoy1gmZmLI7++TJ/ZhOk3Af1KIyc0s7BcI2BcLyTZ2IY6GjvJYxAvSA
l4kyjUxDkTXXl4G2HHM7pB8+zZ+DdtmZaffytZ7Cxkr+j0RQG7EGXWx+ZIcGfHGe
g/DX8iK7ER3Fdw5rL0STOpy6ehM3BHBdu6oeUSKCmHgR5LAaeG+3trwvzbzE9c2a
4mjuVtElOCGRyqsWwLXcXvyRNViMuqH1ZAXdOqGl0Z55ais7Yywc/irWBoOGUj/c
obTuUIYtu1v+6X4H8Yq3dXdY3llmZWaT8irkJbNjq+JNey73ajuyhaJhPFgcUHJx
WXiD6IieYKlca0PuadX4ry7LDctZYK1rSGliGJV9EuuIHfs9aA5Np/WNiOuYJdjB
7QLUezPO0XWuHuT8s9MwyngeDOv/vYImuP6ckLWLp5B+GN/C/d1buIhzXSwF4Uqi
t75UOokm/9sTVDim5wxapwxnG0laTa5up+en8LVTZjASDuaEpuSCmLNtfw0SkKu5
LY8DTldjtuxW6SeSBIVNNDZeyn77DtsH/DQc+qVaspPCHWm7PSASktE8Zwt5tMue
QAHTSEPAHh3ms3Bngu5DAmyiLrql9868Pm2IUo6Sl9xDOjrKP7c/xZ9Z/WRWSwG+
hmNhVs/DCBJ+n1+uta15y7JeVGu4oy286s2GJxrrbCE6OW75NEh6q8CaLE1O6NIF
WpK6DC5+iCpZgCfkSX0f1nC2U/JLs8R99lvFFdUsBf7Q4Ycnfc1k4kkSJp1q1uMh
ngtIBMgSgEqp7K99FYN1xD28EZAyM5ysWPWE4+QUwK9onZZQiWm+UYDhjkW2o1Cu
1SbEKaLqYFaMmjT8H+qyCX/jfR2hxGsk7y5X3jtaytSdvWrUv1Smq8Ua6xLcoVLq
0yzveKMLccBbX/Hf2TqNoB0v2T0/oFXYWpc4dtFnv9SaGdIy5+SAJOFPsCDA78DV
w4udHuvLs2RBQBVrAj5BM3nSCjTDxNLnRcW5Z/gxT5R1NSugQOwRv5Tl1RkPijsq
g2gY+6T1Lq+qQ7/V7/EFSq7WZNlWuG/gpdSr3dczL9KOiwuGFBXHTzaxBZSXBEjw
WyC8nLBqgtijD42gFW3PxFkVfKKMDl4hP66M7K2il3PWQ+O35c7MJcD5obM3lu68
2aZLUT7ZETu3RT5SQaVzuqUs/tswr1MxCjBHFfnWI8ikb/Z4iuRuCz6145tw8nUA
rcRdNhdHVgcY3QohBSUKBmnwP6DehJw/CsYfNEMvT8zF2Lnn13kC+BFqi4YBxLyF
78bC3OeLAU87xAVm1WPIWZJoaQYTvu8d+IJn9M6O9Rn+2kMjjIRkMCtbtx3v+itb
oZCBonpJifFINshEmpOuCQKM8uQ+vnnZc3s8Rm3aqpSo5u9KGghw4dLv8T+2iGQI
SoCaF8GoC7dT7PQLsuLaFGETewPoDZMwSdxz7aLHS/hJYEhDinDQxEYWErq1x1Vm
6Ikjfybqrn6xs87mbSZgdhWddSr/WhCSMGfDzjjVJO+pfrOBsHB9ylq5SCGMDkOR
BclbDzihAh/7cJuYDeSV3xV6RmyIVWani/Vq95wCbRQD0UggMHD6wWJ1MdCaFnp+
/cbivn9975D5MjMj5nzUq62TnBjFITqxQaMA8FkcBMU2rCHSbFt6G6hejERMX+VF
WUwlzUy60lyRWR46wGLcuvr5k1eobOpSIdxT9ufwc1EJM15bbf7RQZ6CJkg0i0Qh
wqn6qI0xQfTOy6RKLK2SR1UgMQtz2inWufz7FPRzJJDChprPBFo+GfXp7R7/NGCx
QXeuoPUL1ZZSi+ImcfBf1uvOiSH3J+3cbBlPvJAtiE3I4VH+qqgB6cGVnMatKyR4
CyYyTAFU7rneZ+EnqMnURGlVfbS1oAfUIiR/yp7i5+qgN6w1ThrAWtjUa5TowhN+
aBSVO8SMr/Vet562B2TA51/NjlLizs0qM97LbE+O+OwrAgL//U6RpDav4Z7XaT9E
UOAQuzdeGyYF8gVGZMi3jo0CeAzCGTYRa/QGtxICMAFjWkLhctpkTNoMdqIfve68
BpwPtX0g/S2PJ+z1AXBZgm+sHVnLfGTzoXSME1bSUrLAhgEtpDl+WoF+DeGb7hOx
wLy7rW8IjVFNZCXWZFj4qEhSGVkQhMd6XXILubaobxIL55OIE8ffrlkr67YnjF22
ltH8Uk75iYErzX2EHnGA/QLUqE/ZXKVHO7Yp6JWkl454NzudP92xaSLhJN1uLkiW
h1sEHVXgxY5FLe12CQJZZZ46K513AsUaMAaGjExDC4F7g8GteyKuE4FeUzI5fR4D
j2OsWjbF7ouMtNaeSrFNurcvtvZ6h4KTxgVzfM6fn7qjPZWzMym4/8MtoadO70BE
T+fxIqkwJo3qNKivSZtvctlMD8g+otAhI9kHRHYADYTXqJ1L0f3fLlUy2rY7fokV
vcpLMPQ6FycfzXVSAvRLThtF7BvdhxpKZ0fsadQOvyXVMydprxwhHpH9gMES7gAk
lCmTj8YzzywegnJCIZKHbROmA/sAGeIXTG+Jl6MQyhV0JmcR5ho5yQvHZ8fS4uC0
tOD/Jrk/jCPgMaCuu/6/HXwEKiRYRbLl0IgU9DHKxTMxWjsgbdvVqbk2Kpuz9S/p
zQf37Hs6c4Ya51pWPKv2yenr4AEVXBMdbW03fj0FiyUxlqeuzsETA+/lG+YcYtXs
fwTTteCQYQCnrj4wABjzK6MJggGZ/QHjp7IzWYuyRHkDOdPppkoiAhCqZA7j6pk+
Fq5CPGSGmZwGQWB/k4eulu9a3k7/X0T+TzUo4XkzWGEZHGtVnud+aBWWAs089r2K
8/12gfH+x6ql5hZx/dy7QWQDlSDZ48L4xTgiEzFPqn/qLTKjuPsCGNyguY7/6dpc
JX03eo8iq1x7jzvQ/Jd7yqSe70MVMDq591BcD+VvHRmejMQ3ybUWvMLqAhTNY08F
U+xflK3N/Tz+BYuycrJWb0Ekw7aJ6bWKaSbekuAUg/iFITqYPt6HV0sAh5o5+Pbs
oJDAYlIYvafIaB79ckHCuWFhI2KO1AXp9Qhv6Fr13WQ3Bi/7P+whABTpbZbE5tuz
WKnAk/KSjUjO/jhNwbWQysR8iwaQJOSCE+cYJcWYBMOdZ1B4gtIY8/DjPeyt8YW0
/U/oEzyUV4mqecNPC9SvfsGBXfJhSSqmoq4mTfe98um+cXkECyfCNmjlogEIEmXG
uYdSgzqQ2hQnh8V7PLC5x//JzN5CzvnKJS35RSMe0EENhaIxqdS/zBTUf2cchW8T
COHrBoLv3kedMJsduvbQNrXUfQwtdKfinku68JailvOZjNHDwoHLzxrwgsPvcq1V
4CwJwFQvGAaZ5VHSt/BoMTk+VI76f1xWrBuoTRKgwBa5LMC57n7OipYA4XEFFKFZ
PkkNUk8eJO+HTCgX1hwT/8Yieo/pB6+YwwwmphsXJiLQU8j5fAC8sdkSW++6jmyC
0s2JzkcrqgTBbuXwoXp2f5RhkHtAAPrjLG522o62xlz3HVyysoWFTPUsO5aIx819
8HSNWktmv3qayqYAEebL1B67Yzvj+cv5qh2dEhNznHVTpefz1cGfFIRgJAYNDsKl
oYBvvM0pIXkQSykPr71sUX1gg9P/ZRsjUzHqqLxASL6QG2UuoR54Hq+KxuY+e8Tw
bGIGfTxJA8ZD1AvQu9uMU1OePQgcvT9LMMZIX9as48wD2Mt6wap7yQY6MbK7x/3u
hjT5UOikqS2Uo0zGw2XXBdPRYlZx5Javq7B/CLdKYHkfRuYbXCcBtmcFTeWgl/AJ
AQ2UOE3nVXIeOMu8q+5Hqq05/CuDe8sikFcq4exV8e8c8VeHzU0EFcTgSDlTTuNl
1/vANIRDvTy0W+FKsD4giozqzBEr8e7g++7Q7j4TVEIHztoLMRd3pEorqsVFQPYP
JbOt/riPKhO+RmLqHTdgC6gEplwVc/HGlzrOzf58qFYmh+nec1UfvlRXaDoVFfIh
5vCAv4hidOKlerehDrVwyOk5tXPhAvA6gTyDNA7v7Y3bB/O2ePQLMyR6IIvqb3uM
QxEDq1QNS+mOHiLlqKivI87p44Nb2tkEy0BPAwsOxJ7QRkBerR6OfjcJZswcmqxI
gl1LJeQUJBj+Zlqk1t0JDznpL0RvVt3YyjH+e/8vKQ/2H0uXTj0b+89JTxs8dF3r
GmNRqlqcam3BIZHPTfsXPaXqSI5eZLS/34noYUfPGsjd2ybDmOASSRmJC2cnhvw0
BXWT2gvVRhCPc9LgFi74sQGVSwKKK0RcG/VeyhwvSgvaTez03U9We9levTx64fDw
wowhJpNEWWFsj0h9M2To14T9CWnGNrDoxOiwemjN3ROaw2DHJ4tU0VHdvWsGtVTP
w5ggUmaaQjfkUTQNrOmrKUXmPSsJjzTFdF8nMvrN3A9up0d65cQc7eCBWTAdA5m2
u+kKQM0Uh9GxQPo2FS94bOi5N0PGPKSVzUA+KQVKAd8MwDRBp8EwLvyKbuT3Lv2Y
T2nDjrgT/ul6h49yU8p1AEBHp/N0IA75+0qTPMSlahMgLqRsSB53FplZ48x/4iwN
ltbZ02M0Py+MXLXAtNCr/MFm0x41D3OPU6j7dpfqmlz+6nJnaRk2brEX+wevv2Vk
J15/jnkYWkcGWEcyU9Bl8TirxUdF03aaTTxe3DzU9uATSbAR5as9jLuoZjhuB5Iy
f2WC/GmjCLyG0H56R6GwDPn9ExhvmisPL/wtKpBfIJtStF6F+xOPImNVj7PQyVKc
OYm7JyxdWagnmn0kPG+vrBtV8vRm2IDfoEvYSut49kn5uVZDLcm+XZZCM1GEMSPm
yn0wcfX1ighYF83GJWWKwsnzYwVMzQCIZuXNPyArfa3g3BcCHEatpK6UGMqYxK+2
rIyc0ANSNt9Vnri4kb4Q++EXfBphoyyGD2ohEhglY2qq5nMWSDRjFO3QtVO5gCHb
elyGdiXzULhtqdg6RpGUy33nLqzRxqFWMvI+mbOWxNRpiFShzjLZP6EegFYXSfcu
UKqvBcXQ5HKtYnfBZGJDXK63hKrVkdm98ACz6PYceno+AYALlri2lOi5IFTyO1SM
KZ98EOBXvUhT81F2xS8UpvbCiLjHsLU3/I+zajpZH+vCQyq4XU8kewq35SjKUMG6
EhNXgI+Ov1EKhltjdPL9LPwK4THX2k3tFChUTr+8NEHDysPsHJEe35vmt3V6PLAB
duHd/SKK1iBIETTpzPcsXRMsprvrzzDMb/ns0I6aH/Sm8lmbHwhnoQF7MIoINiKg
+GaAidOUAt5Ky/RslAMSZ97hl6qQMkYP9Ccv/BWOkki+lAn5x6y2wiCrrVhaDlWA
0gjKWjCEksyV/nd/nH5EyYdwNxlM7vulu3QpU5bQBmRalFeeScNM6ABHZonytfVO
dmMv22ER+nYKpFOZYOqdVp1gLCuKsrrUdlQsQYxjKnlkjSjwixZUow1hj69BZ6L3
Ou1avnDiICynzy8sxmk0ShtR29+skFj+OZKEre84van6n1LS4EVqzQcGCXB0HwTS
UjIGCcHf+TE1L138KEq4swOxa9XbRIP6PY3/0s2jM3QOoUBbTVtATWW3C/x8uOEv
OieKMGbwsE43K7wlfsEcX0mDCh/U1Cj/bcNkZPJem+aNw9hJMo5r7/WB1J9eR+tw
xQW3ucrzwoJqA5VOJGhV791WQVohi041fUcTp2572T0uGzBLHeGGmJ5G0BuNqL46
EPCjSZrOjvAOot4ibYw43msHCpCLQMOasYEXGqnoVFg8ePapArhUY8tnzVWyV+6z
fJmnygtD0pHwybIg/whXt0rYrj+DMBbaN0nnVsXApQAbou4m5HMtX6JjEEE+GhQz
vmppMUufutRBJoctKuZ/69UGSI7uUnLH5oCdem93aLm0LEM8pgsuDP4bhh8pk906
Jea51QD21OFg/7FTqw3Wk88Qb96S66QY7m7e6wRCqxs6ct7E/W099QuLg0YFS6xR
4mP2gduqZJqz8GUH1rMSD0pYIZbEj8SC56yJD+5DP6XbCDPM72wP6fhBUrqzN7bD
oozrhqVLUhfU5zE/OzDJiMRNGeBuFQDqyKoPhg/arB0qlHItYVrKzkjn5ZghHJTt
cBAllcK0tfCOrYXOXfPY008aQbhv2AvPtmqph1kuC3JRYQLDtxdjt0iJ8rygu4T7
tBAtRTLMrEBiPRUsdQobKdGPeb2X0R9/lma56b1JzI+u4YlnoJyf6S/Qh7S7mFd5
zbtO7phWyEl4U0tcKo2XEpreHeOp9PN8zhOcLoxRqwpSGnwG+hKTRswiEr9quuJq
beREDLdTpt0q2kKs6roG1m21tgDMfO4Q4zQvZTv9b4h5CREb2LQmP5MGPxLXTyfy
+AIL5AK3qZhQ2cms9ajXlrq70ERJ1VuUu1QcSHWbMH0L+s6bbSsbFxTxBI30kMfv
DIgIdaKJqMMJK8cGs+3vUGLV6bWbC3J6ktsZH/u5N4vUlc/QWWc76Dng5Ifh5421
v6dive3q7ASxaaoRNjwDry7On9dL6h9jK4mIBXK3OlCj3tP6Yg15J7bcnDAVSr1H
mShY8CX/IhY95pscvD5oiyXhBvM+o2fXlaDIMRou40JcRCjg3d4iXF6Al6dWZq/t
8sb+nGPl3e+ilgLRpsdF0n4Y5y39QnkOjcHP+52urSM0xXoOvexJgZO5twoGDYzd
07ZJ1ierKmoiAfkZ4ZfNJydxG1kNCzzShM14+bO2oZaZUrUvnexoSk4nb0ybVRn9
137TuhJiBbATqZhWZa/WkRUMJouR0M4xYP+CLsF72Ap2FxmOdz5vV/hJDEdAJ0i9
cnS70/aMLAI1yZiNoj5a+6fIudqq+0AcmWP0GHj5pbD6/R8vXC0AMWJ8EkExbQi2
Gjf26h6XZoKJhk+iQY8Syzea5UzUNQSWW8vl1OPU5SMB0hfzCAR1+2iQ9y2kN7Qg
244h9K57K6VZzITDcp0fuziP/Ud8gYOBTwYDCQzHkjRHQ2mfsMeiJnWdw4igzgxh
d4zPcboQfpi9TqkmFJh66ZPoAO1TUaF3/DbGI5iFGxSMNSLGpyALHFSvqUyEGgPR
eELkmk8g4aPOeVtpTXqZu9mhElnSVv2c0JAvAqVbuyqMUI8Ac0NcnjjEk6XghHJC
R2hNASTuDqr/9X8uBXKhVxZ/THnSHX2S4JZ4GkA5i1Fs3WQSbBILs3p5HQhJolqB
cqH+kJlqiKcA6Gmb8HIfVVv3zHNS4rYVJcsRwEDbqaLNGwL0lHKLA/d10jX/D1Aj
a2jQlMaNTTsyUMa4eqJV74L32pWwzD7CrCHsRqM79kVcuwQWZ/SKnCGOCRhdiAoP
WWoSbs+OeJuWoAwdn18OncXPxIK/O2FGTjCRx13QKGwFaVxc9dchqGnt1q/iAGHm
Ahew/HND5gRPleqDz1kakXH+XnmGf1aXZFWuzUVB+qArHnFdRqCwlq+N0PwHvx5R
QYKqBZ6ghTIH1iBJBcXCJgk4Rd1YGEMWM8E5i+5P5tVgVaovXLdBv2XussYtEhzQ
ck/2B6IT8rZfvKzIBN+GbsGLXs7DsI3md193FOiT+A8SHTwfRlsi/MCbTK5gLyQb
D7P/pfE/i2xLZ7DdkV7icJsZIbwDwvv2pdQO95xV9jRGXlAIHAFAge46RoTN6VsG
lXfNm7lExV1lPOX9s98kL39SddOXcRYE7ncWHIDbEgTboYR0usBGcWIkGK3LZrz5
J53nEy0R4L/Mke0gODwOFWLZF9RmviG3q94lS5P5l0hfWXvOiq+gDOGn9gQk8B8U
wBEc36yG3aphnkCq+vp/KLq4FokW0AEZRySF+gtDyQ18U749ZwJUg4y+Xl5+Nup7
remvUFgF1qDFWn22Rd3Y+ZHkT8xQPCVhY+Q0lhpUBNbl4eqlcREwwyDgcEroqKBW
A9eO6snUVdv/QAjBuoZGz7srl51uS9657kjw0m2G6mw2QINYVmHNjwMmi7e52L3E
cA7ETyc6Q8gC2Vb+MjHFlA==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
APrAFzU2R+uIUFSzpSGt/C7k/s0JIZIKzDKFKoAOJGi0YnCZqHlSzaZ9jmcjqUPR
ARtWxtuc0omB2+SPJtegTfjedYfo7Z5aDP13i6CUmKA91Au6LSiDBNBVaTVcvqu4
gZ73+N2J6JcL2lh2B1hHmASVb6GL1LjsoCPO8C1rePVOA5rC8QI3TglOgDp8EJiG
gUwS5jo40D3ZzBQ5tom4vCU9MUSHoLqAGDvEJE3VYYECEWcMutjQi+JSR6o55hRq
CNSfreUtitrKoaaN6+qx//1E35j9wRu5z+iDtDI8ouXa0k+Re/5p860ytPhnG4P9
vPS+nZs9FquWsi9SAcSX6A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4976 )
`pragma protect data_block
SqM9LmYiB+MB5+Vyyo3Wp59XnVuERwFLdbX6nvFqaUn5qq5Qfu0gpVdqgGrcHdoR
VmBRrjRtR1iHfjAO40mbqbK3lPeQRv5I3cFezkEt4EuaKeCR0MDBW0/623k4luKN
XsPtA9DhBCqfWzMWob6NiOVXx0+oAZwkWZyYQHPbL9zZQCSprBnBDNH28RWAg3j2
xz2Tylbj7eTFW4Yl35kppleRn7dNmBYpC2zkOD2AzrBYfeqwRPARU0L7YkIoOGsW
nvknTyk78vC5bSQ87Y+Tw6hj+nEmDKdSp/OilWO3o0uWki5v0Qgv9WL0rbcU0kDA
QCAWRZmAYt/B5oqHyNilCiv+FvDWIagFOVQk+WhfAV32rGZBtUZjM+EHqXqYpDu1
LKZ1NfRwV0iqMRsp/2EvEORpoxkNrky3FAbpnIyBu+DizIjHGtgn4GskvlZiYYwm
/IhPQjg+TN1zFxZ1Pxdq1wJlpEF6aAXydYXOimZ1icrf8ioCh5uoi57fYvBWs09E
ABWGwUoi4bf07xrJDWVsGtl/oAo5M+iJT2JpxyyBJEnM53skMxpjAjhEhm06/v7i
4bTK1dmOIxeNY/UCp/18iEDYFK8kqJgnRgz3hskNvnHyd6o49GXIxSO17z39Ux4W
uDsxOcBPINWGLlsjCPORuakYqKAQtT5zaWTdUa7K77Z8CaHx6O03rPAD2QfRcndj
yT1R6LB5wzNPdmkNH8VrZuqDne4MDTH1NWXGgUieWjKbtd+jbx6kZaWBKdvkcNMW
aMiPKiCQ7oGOJyKHyVW6CLi8Gdxl39aT7/aHjoMXaMqh+ABVr95Uxv7wS1VrwI7e
Zp6md9kjVozBQZ+0VtrqAb2m9+tsb1zN6WrMIm+6cSCc8vXHw+/zhXE9HPjimBzO
aZ+m+h6nveV03zZ5iJ9ge3DCubg2imN8SM4G7JRj8k9Vn6SMYDN0Rn3nK2oopqAK
7BiXAfS4hBQgTv9jPZfHkvRYZ2dXd/UgETL2M4ln/aUZN2PFUBEIbMG9FU4A1iaY
yESTZxm2eDuoy+nYbY6zVXAEV1b49febO379TLPo9Q5CklmYMUiy5lgkOWw37HXg
MPeWPUDD/NgQ/D/3U0rgnjjrmAfYgt9IZvR5XFYOF3sNQzGcxzai2HoT0K32Ttzt
UdcVc2uuyx0RUiKLuhPWTFrZ4qakV8zoiybH0oY76QejS7f2UVW5MM0LzpnXxKoy
T9DdiBQOKoo0UVOhxeky3lvc+WDRg1NPNDAvIjhWHMpX0naooBYmLE5lcPmwzNP+
kbolA+3ggOdCcgBrejkLQGc0H6W5OQk66TD3Bc/ZuCa47+zhEkgSpVtJdVlMfqZ/
zRFsPtS2aKCPqnpu7G/VFajs3nUb1q40i2lup9+7Sh5NW06EA5cE1yW+PrL1kZ2L
XsfuUN+z+VjX0IkzTMQR8DG29NCQ85eEdQ9jRvEqBXC7EXXV5gPyXSEvTBV2yBGo
Loy6NfqkAnQz5JAiQZFGemM8TGBx35tD5T6MBJFBluag/FoMUjxokzDum2YKTVYz
ck4/tphCfrCBOfClFBl6XmSUbUNCOJ1bT2t7xahDx08e8+kqho6VhNS7lPm6Z88c
ERN0TTJUu3PNeOaJ7NsuQevBksnaqGYU/tTHGoXFTMzTjd2BIJURn2PllmAncWbZ
omHSEKBCUczDTDD4psyWlXa38Rn0ocpPTqEZlj+boCJA/w/b4XUAsP2RBYbTZKJP
d13e+qazjJ7HUiz2jnB1XrF+7cxQRuTnvH0n9xdto+e53goNFiSz8KUOp83gOsq4
X5Wn6YM5jwxpbucoVUCzqDe5Ca0Q2uhFyz+DiYtl6Kpb+jorBLHPzhhseYNutBnt
b7K57ynyZtdS1hcpzs4LxLvR+BLE41l35jv+3CEPadfNleeIgEHWM3BHUC+zi+dk
9ejjs10cfyZdNSqBHdAVkHgTOgKxvxtFzwk/qva6cXotBythkPg7nY7z4zFH9rkQ
uy71bRPi8jnEbec90OuOlYPYvepkvhNu5Wf14SrDOWW/+LYjfzBktt/XssZwwkch
pr5JpHHuXyZfW1uT41hSqA2yBnPV5dW2GatN+KRF/mtKj1+Z4FXql/qqWEADQoQ8
bRFHNDnZm1oLQvh1FLCgJ8Zs8S2fhsI1QZpCZQ811VsD7yrDCKBziWtByrzywCNE
Z4wEZG+Jfk6KH5iLKcq617HUYEfG7EcBViLSVWrwxfdPUf9qocJV/8mGdbX4tLXT
CN1G2NR3fI7JohEO0V0AJeSko87fZfIIFGvWoGRdM3yt6kif2WKlDgBKVOyGCsUL
L0MRcSCo4aZd245X2jTSX8vGkaDbHG7Sd+DyoZBcPApx/zWKQzaA8+Lj2K1drgsw
lxxloLLIn3/hSs8dB5jmWqwqnjTRoElqLhyaZUwO4bj3nbyKWTzISYsYG49m5ZCt
bo8kPGnel3YJ46tfSVcg7piJjJW2JuZGyJ6dnuelX//mHJaNg++rbOrgYxmFp/cS
VLIOtyRpkdfGTAgYlgHYA+h7k/EQmxZoEDFckOcuAmCgGwa20DUGUQlEz/ap0CjG
twzXxKK8LZppV6NiCv5L2vwht0/GNcUorblPoAiyWC3Kj4hBuZoGVGX1FFkCFHzo
l5EmB+XHR9FhePqt+sDhC2tNmd/Vgr4+z6ckMuVz4Px/wu5iO314XzIDRFhlHpq+
Mz0Ovt2+46LK8l2s+hFRQN5uHZLep6qWG8hVKdWH33Y3I1GucLiQX/iaLbPCQSUf
Aq/s9JmIy46InHVl5Ngtf2V9NfB83mjViFAfOAf3uZSjKK1rDZplwRV20gz+JjsS
jYiAYcpNFQ6bOUsc8vB8qRzuAsvwL9kCvtiVzNUTmqMSjRuD7B1EsspWLY0EmJ23
2++UxjCUSSgtz3Ty3JOIBnnwG83v0UjOub55FD8bn+nlJODl+kRgpKvJpi8XFdGz
BQODdwOyJdIYamOVIe+s2lE6D7aoxrmK2AwPa6Xzk+owTma7VZ68EbulJRrAQUb3
jwH7cXEv3kL+NvHu6jMdX2rLKgPZASlYq0cUR2sFYRiOCwcMr0+1Egp9JBJhCBuM
gT6/zSb3tl3w960DREZlRNb34ABZtUSfQzbyt8py/Cs24dqxBbAUCG/MOK3/MTyF
FuZ8CHSRmIVrTdm+pKfK6+80Ms22j/o1y7DdTZWm/4MDm5CsJy9Q4VyMEP7/l/kL
2fghCdGfgi//wwhqzfstlz5vhKPTAs/jLOjjrZQqqZF8EMT7Y7ZA5RNm4oXtGjz2
FwRQLDOjBWrMaumk5eu8AYuxtZ5eIBLFJG4xLWqOLHqtwNRzmkDfmPdJGwtHYOT8
MfWxAeUBn4hLNDJNPsGZiU2oA9BDVCKHMGzz9AAaw7Rg3T1IIupQgvmvmv+0jOcM
PTzJqDyEmMpoq5G2I1cH/D8rK/suhpDgKilCLd1prexoBT35ARPkvhvPBo83B4n4
5q1RfIX1z9EAlq392CW5XDFyd5J6I1HS6wxzwINjV5wd7vSVOxTi/LW8uBbNRBdt
YpE5/4KV8f9D7M06aZRxh4dRYwr6Js04N0SxGebWhwjbQCLpFRjUaq46wm0+RCTo
s0neJavqD1jMYgT+eg7ehBhhzPIixh8uXZ3ZL6DTiDIs4c7RAJH9TIebGOx+9uT1
88Eec3EjWCejbIxXZVQwE2asHuwccxzuhQyjQhtsfFDTt591NZj9mxcyKIvLVtJ9
/Jvw4atJemVz7mxeU7BxpsjAcW4xX1gSKWAFzbdVXBFNjyKlPxGOqIVSf+LCrjK4
cztve2HDdHOYxaf+EwF98YS+zpvFXslxeNeiDBzGxJB/kPFHKfKf49XSvOsobQNi
UapmgVfFmK+jGI9NcMFMRtd5oOC+H5ezjnz4ipBi60CKarwjXrdrRwyVMGQ4QQbr
6qEDHe8hEaGTNv98dyZs8NqU5CZCLjpo3iIUrA9JcN+YN/MSS1WPmMduPj+yUMcB
++1yCPa9w28rW8bPJIpbHM7apK9G0HClU92v2XrZ5yVbbcEbGss/lFTlx4bzRwXr
0ERaC4utjQXJyVdl/Dx0W+I+yMjgYNQfDEbPtkytFF17oKI0wmgnRsTUJzpdgGm5
s56KP66DZX4NlvgoWPfuXEUY2Rngp4vq9dItjExJj347zBGKXkKSKbmG0RPiFEZZ
+mjrJ8fO8IhoiMBcjxbP6uRnrT4P5HQY6NB6xQdKObq0TX2BEBjhueJiQ/tMSVbm
Q1ZLPMXGkV3X1is/FVKhdl/cdAAtUcVOfPSRFBBSPaHNGO1rIT3Y0mLcXaJ4Q8mT
1M9tOnrJNADXzI6UIMETwmRoifNqTGf47/H3IrRXgUeuyu8GdxiRiRJhduPPyXFr
6hnYFk4vmo3iPih0rXIqQZjOXmv0ebOK5kFAG5y322rQhSq11JtJs14lpuj7MfpN
6rWy2iBLflAoijpYonxkyZ5gMk8R5J1Cxhab+AARZ7oUnsBMtbc+dn7I09E9yY1U
Q+NracM6OgPq7rgt5qQDD3s91ZB/3+yhBfhyxs/fjvy+mpZAXwUD3zdufYDzmETJ
7zSaT2ychzcjwKssfbvGUtXEwigyHVlnM1zTSzHVpCixbU2g2yTUPtZGGCl8g/by
PbRPEoD0XarkYoxpYCw3nI/eqPHzcP9KqSSxgciZVzsnXWFgQMPKXe9J+v6NULUj
up7/vaFDQIz+u87azqaAnke5dPZZFHKCfw/UOUNB9YJCKLnu3C8VyUdmR4fj0nlI
7bfpL2VUkUXF7FYV/iMnCg4GkRqpkSuZCrMF7J7hpa+u9kv0dJs4a/R/9aH8O8bz
xYwgO0QUQPSb7cGJxiQdcTY0gIyoxfoGEqahOt12zpapM2SZUis3yOMwFhhu7ir6
YtxLiqJB6+O8ekxfcUB9T+UbnXOFxSWbZuTtrLDCrHyKlFEEbl0DScjDuYjfe6dv
4T9rCrueqspDqfm3/SDBvoY7T6SyXSo3HD/ZBKS0l8Y18NfaSG7kGElQP9QIO1O3
6rftXgLj9z/u0VxDyUNtCs2s4eI76zFqyKlUpywyzPoOgHYFiJYngcpt4KEK9EFn
5bZuySVyfVPLqym61xDgVYJeftpQuFKvvWClCMw2O8KBelvVqzBzZUgaT9Q8mgzP
GlVmogAcx6Yv5pbBAT7yXg0TuCYtoEozIVO/zrFAbGF8X9OdcR4E/+HD1L7CbZhE
C0PtvEmpaMvdY3AtevpDp/xMOdCVpK1hNpuLZZb1+HD0praiTILTHi0PDjv9Zopw
YWv059ovpA/dPzSKvu7qyR+JdlutMcIF4L92WuqZIXsnf/IsZuyF68FOwiCM493O
6BePZLk6WQhjaqwahdPq/H4cEOsSfwQqfWohTBYhjIwPcEcbyr02N9W+xjB5MMEv
IidqWgxxVxza5/fAj91EesDfkm3hQ7oWce1CODI5S9os1sZ1cZdbrsvIDKxSrhI7
2JdzqphW7pG/a3zgjfpxBdXrwPKfcAlHl38wtx0Y/0adYf2t3JH0Tc24g2Qdsi1g
cCsTh5AH65UWdYQVuyB0ksQ8G33NQjVUEP7KbFCWrpJOynJh78uuX9e1oZmPzKRl
9Y3EojRtZcbhXrf0A89d/IKGCW0r7t33eEREAELSCGj823PP8t/gN5befR9z2Odj
AaTHUL9epUosPwyDKz3UxZ8On26sISmembbMlJz64VH1gRQ9bXfWTQreUZ76ETdD
io/YAVzyopueKJ6jRj1eSb3cSWF02ojY4RWO2zJbh2n/hhwDfrlkXJ4YSFbJWgGB
wI9gB+0fu8/73J38PwrKdyZD3JmNsfveikL5j0Rzl6Sl/f5N6lfSCfHORuN6ahGg
yMWGXE/5eVeZENLug+m/Y3QNVtmcxIOISJlcZtjR4BgsnSkeK1nMdQ10CYCKY9SP
AIGBLXqVRYuAnVP7PGhZp2F6meHkvzcI5A3pi+bvZLTN3IAGGKPVQ3Lx+Zft5xeE
yJsSaQ+IdjhS3QMJD1VJooM6Dx634BAT1buB+e/I8sUIsVJKof/tbE8qgPyKeGcK
ptqt12H+m1bO/+sbcFHtY1RrWl0gBMDcXq4Q3+XA03U2ExhiVqK43RtOkFuvgHIk
5fyWyksdagZ9PI7qYNVSFes40Lp6DFsKL3B3yifBWT8m95hnsWF6wlHN0Z5LRT1i
OFtl8ucYTWz08EnM1Fhy73hCrEshSHPgkxNOyCkf4USvS4cXy4g159o7rJL/PIU0
1+9J+ZAYDV542emge2JzYfBVxI/p6iqQt3Muv3rYb9l0q6JTyFmxJUaCL3hthoLy
HoWLi+mfklFBaaUY4Mb/+o9aGNk9vQwu46N10f22+8MRLdJnoAh88wKxsWhSfd8L
0jwuhIi361dbc9US/lJqp/J6Ud5H43KWNpmccaQpED3VM0sjTtt/M/m/YpT+DC2j
/wIjuwQFNHi8CxxehrHW60o4yEdM5RiO3y9GATglizjIN9GY+q9J/Gx6dBfccYW6
aRbC/zk8Bwk4jCplIm4HRIYKa/4OrASer/iEraKRxV6zo2UczQTPI7LTmmBIVCMk
Awsn/ulDtajMHqPikUNYl62Qjm2rG5dDzFFeM2k5UnR51KDJiOGva3z1hzQHUub+
IkiYp6Jkf6Go7KrtuELtl4eWWVxgNY1adRqmr+dKLxU=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gTL34Y5KH+KOTQl8B4uU2PHjK0hKyLsljjrKFH9h684DJCoc4KfDiwqqGW+00Jp0
DGvAGNLIblT4sg4yOI9+YRHfWdIc+1OHoR9BMzEEs6LVLM9qET6/JQGx7dCh/Egl
15D6s3Zf6DFla92ae+T/JpGkmnoGwIbnY5Nr0d5Ccm5Yci1/+EBDU2juj6MK2l01
lvTvgMsBAtxaPefFayZJrdtndlGdmAM7JJ6uPTTJa3Ct/JtMaMZBeChHLq192+rz
mzLKSeJG83WjxIZhSZvW2s0Gcve1nkEPy5j2R1xTvy9B26e4J1wyqyN6zIaqBc0n
AdMpbIxMY8ALW45YJH7VOw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5344 )
`pragma protect data_block
RZX0nsFldirqJbe5USrqvGJPl6Tv7fn9Hrr/LhyRIpS9EqVL5T/Bp8Nid+d8vs5g
azSJSnIJ4Nsqr6GF1spNRB3ZpaXajDSFzs0UY1C6jXzx0xlVYMIUFbGvkhbVJe/B
TQ2Fxg2KNB/36v3DkEBDz4tXDJbdJZf32/OURlub0Awcq2dzsLQwyBUNY9Wf1VwN
OjDnoPktFj4C90JHm6deIYLY/sZdW25h95Ziun9AB9qGIZBUulgXyxbq55R1rtFt
G1Mc9t5vhv8lGQ+0LBFSGeHza3yrfKjXDViP0rQpVXCXnNhoRKBlJVne3iap/kcJ
cPTTVaIzjMfwfk57/ONRo4PZxEY6qUu3ar2PQB0wgTHrxAOAqmNjrf9AqLG+MDpB
qNyYN5FVGDPgk+v6Ga6Ymz3gK4yXtmNYfonOlBjYpd8dHVuKQk5oStGG0tE90oyV
Ur02mdQgMa8vMwx05QzFf5ggpvPnCcSlnQGewI2YNFU+GbuVW+4LAC7RhDJw22du
7hVqHzmw2y0rgTsrF5jjuhkryFmrsCddmkOLx4WnzIh7Q6y2qP87mVmHhjbyPNVk
WoTrtPDMqmAy5DB3/kIplszTx3Ru/C5xwpOiptyJitS6Mx4/0Bpnd7oEjwO6ToSt
SjY5Wt9gCiRYIRjiV2PkICIZqhKl/e3wj9lz/EfClsBmRdRbuvsj9psc2RSSCvNQ
gbue2RUyfhoJDmOnMsV8Qo6EB6TjG3hb81duh5dsZtCYd+WMAr108EWqqjoIuNCs
9UVHwnlctACtKvBP1JDrrJs/6085R/Et06ObNLRe3JDPXyyUEJvYC16weIUmhBdn
xKLc05ljW+tz0WO4tZ+jQWiW4qjJEw+RIWS0nlEpEIBkmh2TNuuo0ilmuTc6NMc7
7cfPEDGRc5jnj8tf6KdZQkLdC5bbcr+L22V/Sf5PyZLhso4qRyOJdGDjKN+e89zr
7U2BevfZD4RQiEuYjrx7UJiohUiPEbUT7rnKSZKnf9wMoMR4qjaSd0cgZFZyZm9j
1S59qbaLq0IfSdRcdrfRv//UgBilibTiwKkIkJT2+uejEDCQ+/xRIcfdXMCoum7q
xAqUlIuOGkB6v/SW+mUEO046DEREvuOa9UEXAQzJzulyE552mTYYmXKnk+Mik6nK
jgvJYjrdMuj3Ji/tHEXvRwrTK+ujA14VqrJkNVCcJgTGMc5NJxdfVtN0fGQLXSdf
5CeyN2KYjUAEXvQudMZ9VLP2fULqzplRokSACtDz6Hp2oh7/Vx9rLYWGewBctOeo
pcjnjQfzZW50HkHivApajfbrPc663tuQlPoAJKhcn0/iVwDGmEYj71clVfD/fqJz
Wi4id0j0JAM9XMwsQEgM5f9JfQ3B0AojB9BdRb6MCZkm7vWGKkQrMawMin7XompU
g9jColihs7x2ZX0UHoFk3NNz0Rbs/oSeeTyaef8pFg0fj7r8Kif58byQgYSO0KCm
NBAqGQyBNHyi0K4in9kHaE0vaDaBsJsUXaMDCg5h+422OsQdSSKbDjCWC0lx2b69
vf7CZf2JG714hra/hNL3+BbhcxndaJCMA2InlfADMRCqT7O1LIhzOHcCoxhbzb3b
NND/em6XirnWBSFfEfJEjL5SvjZPigb5ekyiF3dJ2g8p78g23/krZ9+FDQYjC0iz
RI3/cDD45slFzCaLtqqvtkci76/g25ciBBpt2o67QAXjIQ4NQ9gzc5V13iZfx8DL
LQ3OFz6xKgPiMUH4upm5trV5HEtJrHDiLlc2bzVsWndZ752il21i62huZqiQZuUH
SUTpAvVdLdLImSDDDp9JOGMX2crtJ9tfenjSYtLMOC3ZIXo18+uKyxISD54uCSrW
KvLyDPPFS081Pt9nQ7k8hYgoulLmMZSH+jnpfaooZVJ0wmoug4n+a2NdLb2RnvX9
dF8wml59MpbnI9Ty8ukTa8GykXQqa6qCK7HC+XFECNTRHoeo/r3IC0OG8nBAYGul
x2L8f83tiNACiOKbNwynsv6Ir6IEaxZ8fGrJMbJxOYGXd/siexxvx3N/K9JsOpNs
HU010jHnUTLR4cd3HUvJx3jNK/fhM46rSBuI2pxG1V0zufn8fOQeJFYXL5xAEHdf
o+10FX6R4q6eJZRNoDs92YJboXZ9LiAFrmLqyhsVT3FLn4pxKyZZ+byZwK/mTNmN
Xjeu2ROTY4hgCukgKbQcrniD/DTDFnf9cu8dCLjS9+zXSVDzb5jHERRWrXjUQaaN
z5DVxiXknmjgQWaQQzrHWWnPqCYOOUvBnPh+GZMAuvCQzmazC7rh7r22+TRg7aPM
gg4ueY5Wqz2PG4+PTWYhXRKsld1HscIf8nzRXsXty9olG5YXL7Izr35OuZBLtVjq
rTSpRu0Irx8luOlboj3SukAthW/tgY5INUA+iZwG5MVBFNFgXTz+15d/Z0ThOsy1
Og7QHxK/IpG0jpHERSegFN5wCvhH83ZDE0ql1KJw521gJ/v39+mM/Vi8C3vJSthF
aCJdfoJLn+9QGl2LgjV5p+FckBK69LzarhxcV50IrT+lErj8XSzd7B1GDTW3Sque
1G1ZsivT3nljvy8Wp4PGrcLDmqzvdt4hnP3ripATRTSkmm8orROGideshPCV0DyK
L9/wqEfnZOZIBVobikDwy2uxB0L/W7pXWFdGezlFVGN868dSsL49pkqRRSlqkpM1
r04NE0Y1M8SwwSHGvmUw5YoQdrg2Z7IIgiBLDL3JfgPC8TzJg7wMfjgW5IqrM+Pq
eVmYQOsVtb35X8xlVyT6CiuQMjawd7ymIoJQw48hPLPjRvkVqpNvuPdUtxahKJ9b
tqXXe8n8zEED6iLPJdBpZseDo7enVryO85kQdytwMTLYhExRSQUF3G6iZVz+wgf7
4S2uKWscmGaWJw2zZTEP2uW37LPiTGHXNznazMXEzQ+k+KlUhzm1AogHeJ4IUwdV
Qazdu3Y6E/GpQ9XHEALj9NFEQbpJvOsUC10T1KmNTBwE28Hq6Pe6ZxQgcMCEQH7p
z2vkMEC9wy9ZxU7oUZ/mA8SI60Z8SBw/gHyXGIwxQUthcNkEy162/+RYh5GFtR3D
L0Y0UbqoDdrsWjzkiTmVKl1nBVAwhWrb/YAToTzRYi6cacJgGWwhOZH7Rzqo8zRG
63SaZpNgpPKVptl/jMsb7uvqjGT03oMNhFvTm9W2wg41foBfzVwPiTOrMAKnCg8J
tMRb/WJ+b3I+oifLbmjygYHHsicGPFNGjdVvgvdKolpn52/C7cG0hbm5Og3n8Q3x
1vEkDGm/ZQXpVZJiqFLuC9WEYHLCcq5ue4ZtLyyZclCTLUO1RXu7656CdSyEOnXu
ZrJcC1xGZBG845qC22gTOBlxT45z9XlKPVuMPuQKFoV+PQT5+pErl7L1b2nWBfkK
vXHUNNTfXPEXgr4V44FmczTsoibjwzLvxSCjQXdazpn4nfFq4p4x6EUUCZ/eO7DB
rjnlrR11rQ/Dbgydba1DlkQkIr210EuzqOOva4/9MsLlIqhBgbhWv/rl7ZVF/BXC
m3+sWmuW73S+LGNvoMeEgQGiaM2LbtmgrP+dCv3Rj5o6KORDUe1eiDNXIKih4hhH
U+v6YqXaRu2f64omRIJ6UktHAMdMPcIvJZPAOHdPbsgrphtcFEsbX/GjnpdQEN1f
+EKuAG88AAPcD26X9P4SbuSD7u8zhZzPyJ4pKJDucn7onLlvOMZl8OvpLz4uYRMh
OliJ9ovYXJxaECDHERPaoP+1Kp6aFQHQcofYHyPQxUwquZBGqWau6bHbi3DBN8Zl
+g/7SyWanLybmkmMEoyPLr+P+ZDrN5Vks5u7/mxgS7MpDn9ttC9b6BlWF1gL8hg1
vzajAJ9VJyaKxzXqY6xHoiccWJq42P0FT7/K0w61dtkc0YWMHnZq57v0RCAYG1Zy
2ngkrD5wzuuukI/OYFNYCBBrqleDfvBOzSb1LnrzzFpm7ISfolVvkonVcLgjKBhr
IXvYH6kOMUS6EgwJYSUPTXAk1KEUmIIKVtRg0IsNT5yhoPnPohKOZtY525cAf6+4
K7UajQPBYpsBwiVWOJ5VlDdEWxb2GeHytQGgPA7zZmMBLA0uoIwojhMjzr5r6FJE
KbAfMb66hAYaG+TvQcAcKCUhY9lT5JKE3ovrdhdHfxubLDlpBsf7AASbqHEUZaoh
16R1v50z/3kYci4AyLo96rjja3XliLkhTEXn9QqYrerkndcFlI4cVAoW4u5yKKMw
g0gOIQugHif43QkAXHC+xHB4lF5UADWKxDXWvCFqAJGHRdxlAsEW7nEbE40INF2A
FW6WdgMqj4eZ3espTCjh9717dZQR2380hZPjDXPlx4BfVRnb6/T+RZN4b89UibSM
8OvJX8UIX2WyJONOLOefcdRduqBvchNX0gMPhsAdnfWmj+9H12zk1XBzGsrOUCiW
fRYRiILIH7i9ydZA3PTej8Nqmg6jSUXvyP/6ZTSJaSnCVQKySExPWkbQG/DGhmjU
z2f0aiQdTRFJBqrU2gBaLh/aEIFWJSNb1V6TL1dTR8tu61er73JxdfTdvf1r6uB+
odavjFItQUJPyAnzq9wVHtRDBRWtjSzGLsLadzRBHmpgbh0MWkqLSgezc/JB6lLK
DcyzAQ/pUhJeUFId3IFnOeKnvCRslA2TxFOOiWBTa9tKd+LEta43G7Cr03spkFQ8
YWyJCqKFqoy10KX1DHWuDWzbyAdhc2E92HGd0v8GUjVPqdX9j8bsIs1Lj+I0KDfJ
R3L/mhO+aQUGIFs6Kgu8XkvgCvRm8lqiKBuswJjJ+GevFn2EPDMMnzywhLk+8O9T
erA4zPzpHsrh6+k8W87KGNloW0ntvnmRfOQzXaX33LD6qrOaThHsRx/wNffW69L6
ltV5Z1x6MGr71O/uaek7J0ejkSIzqdfWcYgtOPOqoLpOECZdG9G98o4vx5w1W9ZX
XnTtFMwcPgHdZrB4oYZyI6JXiCzjZqmtARzc/7+UjeGL+hm+tiKhI5AX2D/JrJYY
xEzdwuAn1J2whbHiv3J70yNmCULubSWJaqSyFQ8QPbbngYZQ/6knJWYp7XoQh4dy
NYsEixLAN9Xhdutd9dnBV6uj9aRHtyvEB9uNVWtvKZ9eiy51yOuoVqiFS+MKsrnG
ZyREVkatu4iNOWZzu+DyZTzp9TpWJOYuQQmxm3Q+RlfkqSr4wEeRYxXv/YgnX+OQ
ikyanDoJ6qS8zN3fbnGPYLsKhufYAbRpMK1FiPamA8uEM8uMZb81eexMx+ow0ech
IMGEPtAJHVAOze1JWcvPvtzpuCKpbfuCfOzdJ7umh+9lhVugxxfoufC+XGrf4lUo
tQEC9Biiom2Qn3QjG2oENQtdEa2At7Th0TKHW8YOEcApIoN8Z81CitjOCoHYD6bf
6Rh3Wt67fmvgirpmOqte8t/vJ3/zIHoxZ8TB+z4CE3NW7V0auRlUbAb8LQZrezGq
f83Rx9CNrhoDZQ2a/MukcRAL+K/NZqX/eqKmuajgg4b3QnIlQU7OLTRe1gCDqgrh
3wMfXihZWqn2Jh0RDfnYz94Ir+kO6R1SmQFH1gur5HpmWMcLS20LARdpDG3z2tzw
RLb+SN8QO1Ck7JGn/XUVta3XD1LPdvPhtWwOYhqZyDx77Uz5xZrUGBim+1AL5rDi
4ZUE2C8zF5KoIjpn/jXe+p/Vtn2FlO7fe0YohKmgA/H/b4+7iPsfdo2Ox2rJE51Y
HkdgVEPU0XBPUZrqcDvcwT3rkuyuuMyyhMTTTOZgvr2i5s9qGsxIyKUPrc75Bw+B
vqgKC4KgwTC9wHiclYKJ/Hrzf/VM+jHhkm+zJgwqEdXNFQYiqzX4V97HwqG4Ou2T
1lAFKjsgzZh+8Av97XzymGRd8iMj2pOmNhnT5Sjbxt8BFShGdshDdIOpnpqxyiDF
5wyNt4IAbXUCtCptsAmHVIMzsekxiJ5Gn8TefHuiwYdx7MS5/QnzIsWo0qpWpN/h
lxomVebu01S4kpuAvCVZTlA5Z5sp9sha0gSfm+lxI6gAjitL5kWQuXt7zsuHU3ba
6ulAdMf6A5bKLsOoFb13P8Yjnvdn3njt9HLchiWEnfA6GlpgxmFWA65FulLEaat1
JRniiWeIjOdQo+wOYEHhboe3UXB+8lROWPrr3FA4h6Own4m7JpHgd41WiajoYLmk
DBt+3rIZkVTaHrglpyzjxeov4VvvnRlWmwmHvobp8RpCrCMzGs9A8r2Jzh0YQx/Z
yMc10DZtqlkF/hHTScJ6cB2oBFBAdN8OSCMwzyeUzDeiobwj6n13Mlp519H2fey8
+ROrdSJwdpsLEzjaH+WraPTtpqaB9LuZMWEiHxwzt+2/sqvKW84TMizSEVB3QdLv
IxxX2O1iX8pAcAOb3lq6+evht9qLSIJoP9ha4O3wkwFK4sBSlaadXafoI4QfFQr2
Z6Dm6ibKcywcFZabLh+41qpG/56HhUDqSRdUy+pivegMXfMI3AvGOPnR/uHk7otV
ol9chkynLKPR6QbNsiDn2YJT/Hx38wIx/NkfTVXPQfr5rneC6+pbrrth4IdtDX2n
gNDtMWvWwxdsGYMS25JaCgy/4LFYDdNa4BAtcs/5pt5hJgT/LemKj2ejiMltvULg
ZTVN8TvJmNwjrvdQVXYtFeEXEfHfSRzi5zJUcEY0Qlkmbm8vIRP4qtt1HZq5Xy7a
JcHnz+l2G4MoDrzyGj+xtwD4KgwvM5SkjVNNaTfXT+Dn/uarNpchACPr/fi9BsTF
fGISbFZNf5BfLOCWoNS5pmUzEC6RACiWwISHrYhw2FrbG8W40munYEU1KFanYj5q
HgoJAwBEeDu8II6+1PZEYs/+wzx8/vawfxJMOzyuUWBBpTHgCAu7wctEZth1FbXa
TdvAM8TTlSgi0yzbRk1UaSycricNn/eSEewnephbqtTKjhkvtsTGBE6EXqT0AgDk
SZoVpnCaqfm6J95TWx6ln9USPgB/tU6K9zRy/ThMWEe9xwhIgfu/XOpcu7vs7c5S
YD12lpVec54dSTNbaCDzWLfu5SPwCz68su8q+NAVyfBnuMFvjuBbcWINxy3IRdHG
Ny93wSx0eHoMu9xnDU90diISxXXRbCOHBGv1ccuqG1sjel8XBR+g7WR0eqAUBjwT
cwUdPADSxRxo5uVYbtRzVw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
OyhW6nXGmjmIFraOrwAD8OhcF29/XMkZzTFPD7fJ2kv+r469jZguWmbBgc6Tjwwk
CQ3MxXLGAvKNgqnpdesaxI9FJ+o+8X4Ozom+q0tYS0dIqb3DURh2SJoXl56CmDg9
s8438aQ6W5rXAtMOeaOZAo+Mi8U5WF8IS7tFUuQ1bpSaGKtbnr8mySEulqijA/Nj
ezaNa9aKQcWcO0OVCkFVEIQLbpG9n/l0HWExUg1Q0aLS/+WuT2RlBdOYMSixBL2W
3HA5q+/fdIV+cvEjwLo1cqJblgpJJLPRY2N3TBl9XQSTgaJjEOUR+kY6Iv/CnH75
0Kynx96NN/26qaQop6+X7w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 13088 )
`pragma protect data_block
U+uRtqKlrAU9qlSZfl8zpyQXUftIMwPNO6Nd5pD4tGEOIFWxR/uMMegWcMVbvMd7
WjG3SJybvApjFeRY6FFs+m+XdFrHkItFP/+OCIa3gMnOfmgTU/iK9BzEPtnQxbR+
Yt1j05T2HXhLyH3a4DnnoFp228nXnD0QXupGzP1p92yrlaV+eVBl3Ckfy3YLQSP8
zLYAiLdUN0uvGPWgsCFAr4gxCOwdjKj20VDA6gLfwwbMwNcXHM0TUi0/jh5Vr+ma
WwLNbY8GK+GSnnAvUWORSl+zU6yR9ulUGcqfS5cA4lyrorRi0zXGMFYPS94gZ+uF
sHBJL5VyjsbRAIthoESHEn36Q0/6qTqwsvuF5t2JFze8fGmwEBL4y6t3lw+h/CkC
cusfSSFcaNAVWQrZx/GUmnE4h5Wh33h/ncZcbozCwIB6LjJVBu0et18gh+isWlYl
Pa3pQSzxEhLxDN9CBAxChe/C52DxHKzrIJoLKhz10ParDDeTQ+mNBKB33EYoszZW
sOJ0pffs/QZ1j6bKLFrtJ+KyHWLNW0zoAZ5jEzupVH/mHz/OiGeFEnRe4kw2rS1I
VcnBckMYePbs4Qd+oVdX582B1DC4SYzGHg6OMncWj0eO9A2uCarjCZ5LW4YzzEoe
Non7Cv/f3LZoOcfQJCuYaugnZXWpwcXGz6A8g6UpJ6aX5SJfig+28g6QLIDaK1sj
My4CEjRZCtgr6fdeGfL5XocxVZBOlQ/JygbARoGIdWYpu3FdT2hTdtf9AgAojmJH
zC19mNjWGw35Bz2Xj2OUK3PGBsbtlkqwMispACGlo2iJ6T3APQdD2QhL+DUCzPWN
aUtbRkQZvxs7X4t428ov32zltyxp2md4YsIftpqapgQoP61OcEhviQtaFR48XRyz
neEcPjEooMxAFk28jTIp3MNSiMHuFVtuEIOPK3YxTFjKpgwa2B/MKOAsb/4/2ZHg
2IgHr6Y8+HiOxciswBKBaopWM9K2rzj8fvid2RL5fjW8g9yGSNby6l6aV9AWlhK9
SrSDlux9jfOU2hdw/h5PQqF1q1JanYOZmOXLGNgkDSt/gXUjlXCTSRxHrRXzOsOH
5DpB7s1t1L0L1qy5kytBEUruyoz2wjLzL7Y6CF41TUwxG85OwIKWp89I5thUQfjJ
q9Od6QLHZUTqzVpIPCGaz1g78Hxjaupedg5k9N+XTUtfrAaNFc2/KSQvTIFXoVaJ
wwmSi90AiZoAN+DFyKrWnchxgHIy9Kqqiq0HV7ikAvhV523cQgR8wYTSyUB81pKQ
NenpC4QtnTGN5gm0n9dtEenIdxtuwl7Ci0ZfE4x4KmW/B+jeSdooWP5JEJ4I+7Yn
MM+BywCrVJPFwUZc+dAFQkPqXdXdFF1F0Vm809teRBfvg4SxVuVXjzS7mSvYjCdt
Q2USTze2fqIiP0TlioW6o98VSqX8BE4+RlorzmBi5dNLHD8sqBHiMqVIaFbqirci
8HzkTJ1e66m9RvYc52F9Dmz1HBorKF1H7AbnHypTlxOnOLusDgji+usm1AyGVgrQ
61Es854gBbCOrn5yFg0obe4xilpePLR5zIikj6p5aAh/RUKycpnhI6bpApyTwI94
kqTghNbiWQTWnxWQRuDtRN6V7nI/dYYM/WEJP0GvVz45eqHDJXJ4p0TatuU3WpuG
Qo/kzBulUpf/zEYAEVrdnQSg2ro7n5evzfpy43Ru/7yARC7l6FJ4sBEz+bwIjfeY
MdfDyT+5wG2368tbL3a5SGV356rSwH45IinlBIjeiPNT+xonvmVOuFj/eeOcMvGt
HU8MNR1R+XuPX7Re+Je4SzAKdaym1cUm0kvem7t7W0UqTLeDuJdbctTF5a/VFbhI
SVfn1NCnNEEJw5AMF/TJKVtrfswbuIh5zPgGJcaIngWyBC+8uL7BFO/3Q28j42nx
HlaLS8NX5tO2D0cMSIHbBg9sk0MubwSzQzYXOXoAt5Iq2Gzb/cE5kqE8G+w3ByWd
mnQJgg6ZKKO6PFSdmqHco7CN8gu0Ll3DSttgeJAMygW8u91d0wcOTcsCEUnfNvu3
s19c50m2cyc5Z6dc4yDaYXOzGLtJxhjpc5BNt+RIvSvEDqUDJjf7fX01+RsVd7IC
KB3OMVKgU5pGkAvcZKu3y4ki6zH9TLJP2Su0Qn2azHISMCnRT4Oya8oJCkKJ78ki
ri3CsDTh9vn7oNosCL/DfZexrjBZx9EN1zBYWCRb/pIqYYkc4fhGWcAzaBhn7v/M
UN9zizbcIIla7DL2mqAYMYMEMHtse+kuRRbImS0VGTZ/VJhxmNHIgO8zSlwgzWps
5iqyza0EYUd+9Jcy8s+BHLxhuvQuaXSFEQqH99Lmn6GgngmZXqJ7Zu3fuzMMSU9M
ODQvUGLKmOJmSV9OFg+uiUyEvcEEkZutZNfYfze0yqCVfY0E2utUYdd6sY9xH8xA
Wf4RjjBJdv7Xn49E6ZEBkyDmCRMeg6J1JzS+jH2sSVTJ0N5J4EAXfk1mAnEaKYS/
L+15iLyp5uYZ+i+E/E8/FMhPetxtTzzAV5oqu/vI4MwS/zH7qmNTP1b1JeH0XyO7
X7ct1TEqbeTWfEKnbz/rpvwxX+9QT81fwFDPjINcvDS951rXG1OPYvggHH5rBPqA
oBdkuQ5QyXsucGGdvvddPXm4eQMutbRoyftUvFUfyqoyAwggHHsP+vNgBqwlrG7M
gBeiZCt6utc70t1z1OJTai8zjTQ5icoct/aGGDY5waLTH/7lUzK/zQB+ulU7sU81
bRxtEpdoCMy+3H5BnWFBlhneKlsUeg7oAfdT9AOBZImP7W9mlb8KKpDqUT6CMI4A
jPOXb/520nEymdu0Pr49pjG8YZep2n/WHYPqbBg/lFC5HwvF+F8vuVXnEARWEqWF
0uxKYcXeZ0VRtUZSl2Cw71n5LfbhgzQ53eRLNC1WtJSZJUGF8JJHc4AuT6vhfW2J
BcwO7vq+U709R2xkhsfNSWqTxqAnj1JNWzWGTyK1rvriqBx02gVRJutKnvVPMlTF
WfPyG+FSGq5ruH+rg0pbbqu0HV8Ohw8qgKi/sptaRBI/DOHw3hj5zf5y+TY8DmSG
oJOzmhXCXqoiO2mmIaigf+u2Ta8oRw50jfzNJzUY74DneCTnSZJXKKBX8bzS4+nk
Xk5r4xMZp0KL9ZBHp7D1D9fDeTaVQh9nSNxeHNqi1RSRSZSc8+gfiNyUn704ajyq
m9wO4Gjh4BtnJUwZDCgrQ8Q0JYuyATMPeDSPKtp+tw+L4yNY0pD7TK3QGWjNS/oV
8gAIOzoX5DspA9DtGAMLZk7iTBVysHkGoI1UM0u2agsZFcOZLLESODSib2bbmHUG
uEIwo2tfGAq5DXFJyyb4IHOCrMeCBnmnc2XaUYV+/u5kf/mO/hKm9kHhtb2bPJ3s
+ScLMDqDkIItN/Vb8XQJNtUOe5xp3XolXk+sAi5fGeO4gABUPVRNWXWXJxI2t/um
U3zVo3Dc4pMAO0f8AzQ3/8mCGbaXkZK11mam40PtHSS97Ue9lbiWBcGonSRugYbT
+QLAfXfv5eGJ4IxuLHCyIcPw1koa+oeAJ9nUINzbMX+h3Qn8vURPnJbMCn064KlP
NQQGdZoJ1gOW5P8TUqJo+K/c0+JvMcosdMmDCCDUx7CXy28qQt836oK5M+MT59Do
NwQf2UqvyZnm9RG2vWZJHPJc/GJ86Ze5uHAwo5uMWWJQh76W3dLB2Bf+/X52rGOq
VnoCAmyO9Edr4UQacoMjvGgMHG7N19HwHZ5fZ06zaUCb/VxBeIx1JGulZUVjcI1H
+l3JJj1vYMdnaVH9FTxaycb6+7LQOuAxeW/lUNM2sWRtdj/4Lb2BwuTBZHpz4k+b
mnwMPtSelDeBhmZvYgJMzwXG5JQSdfoyHWN6C5Ogrr5uUlwM1Jn4CRCZ1KHS43vv
6RefKtYMCTBG6r17Avgg1+KRmsohFI85NTOrb9A9ippSXMsc+B3aZ5ui4azT5mOW
q/TTbi4KoXnyeel4L1Y/mi0XnWQUtc6vkaFSIUmqiTX8RamLE4YorEgsIc+fOlYR
LngD9E6EXI/0Mx99lNbUOJZkkrUYi/rpLK3ud+tg2QMj7IHOuszIQta/u1yJ4Pom
tsFlNCDCurH6rGZw86/TI1h1eJLKlCvzqC4XONWeSmztcHdJ3CqAqbFblwMIy6Od
dYJQdkR5lah5KxZ+Fc5awy6ELQCajCHmb6+LBmafaanmMF2SvgMNcdoKKOUtRsgu
T5gCh/M8zf+a0wW3KsihUqftcnSNXT/e13e03xf9w7u2rpnESWq27uWaInsYtvpB
zNdMVLpRZ8v57yTrm+nRp0uTd8MnXEbxGigk7FQMqKtxH9n++NoMfQoHoAHpnhI0
1bsVPD4kT2d2LyvZLQOR+WqH5QRLoXd+sV5Lf5/ZXCunQpZxfQKBRAPM0vpC1uu3
UCD6H+5ytK3dR5t4A6d6VFFUhDrrpFRRipy7JUN1SkAemVTMVpMsE4wvTmHpZltV
e4vVAr+oNQkWi817fi6U/ZcTX/Ec/9SjLZ4vTTnCardSwrPWxGBh5mbW/D+4kaLu
d98gKxls8HQjgrFeYwghS70LfDT0MbdN5/euZUTL4Vw1otCLZYnrWqcdjWpDi6oi
LdopsA9wyY3CA/b4S6ZtjIGaKxRl5gouS4boGxXNsB5IYDWEAguR4PDX1mGuIUSX
2r3SPwFoaYVBUPy/I8VB2BGd5h4HNebFXUYjzp5wJVN7k0v11hX5Uv3evCjZFGwK
CBVJsPOzaqUb5SfTZrBRj2uSQgBq/fcJ55tgFYHcpqzFsWany+lkC6txGHmmctc/
ggVEgZjkEK++BcHPqjcS1tm8FG5BmAstLXu2T2PBHJL07C5I7iIg48Y3MezaQeQs
tNWM+rqBbzXqj4wsmnEikY2OBtp0vOJwfJu5KLP+fcnYz1MHBZGzYUlYoIavZ2zn
IFhgpHTmJgxroD579V74Of8+n+1J0m1W+457ykOHYoF6wbIvPPsImdnP44cvguaa
CH1i8M4v7kbKg5qlvKDAnqxnlP4faccAYJ7CHGRxJ1dxB+359ds1IL1kWHJVXc3E
KPu9vGfRfh8d6HDcMpkDKPSgwuqjHxXh1bkfm/dznLpxgeXQHzOSfkPDBoBxJeUM
GIq9oy0YLjBB+ZP4vyNHHkEdS/32v3pdjui/ewPDuGjKMQ0x2TY4z79gOCjd9try
0yZ3D6vuZ9n+FgjNl2RY/QyOohZ8+R/N9QEwGByQUA2wZWGBMmHsm8M0bODkd3Lx
7TjMJhUZE6AVX3QS8v4bnxH6SA4RrWSBMudVr9Lu5bEaWqIGn4Xe7Iqcm5P/qlpe
H0bGeCnnDPfonF45sns/t6M+b9iIc1LNSUPfK2Hwv03k8L+xX3gEQHcQlEVsQmrB
PGKIIOJY8TbgYHvHeNH0omIM7MqOZa0D7PoN/dqNcCfaVbszZLMKokF3sXbFoPxd
KNJJvM0i+fy51p7N/R87cqPbi5yVmSWLq20BYBqGcGncqNk6ayb9FBe7Ri0w26KK
4KrG2CBqeGX6Z11bDQRK7RIoYm4qTfXjqQkX5RSIdH2aQkBUWEsTS4Qq26VKwyq9
ct2nzATXV08aIHz5XxPfz9+ue+x/7Oxo2Kkwpqp4+eRNpgs4thKf0QVGaS8r1Ymi
WbHRQGi8n2yGu+ndGM0WBqmC6VeS5NjpcpU/91uHLXK8IoaXnz5bmYRAEnOWDEMA
pthG2bwL/+JErc0aB4waAqeJlkeqwCSOflklbjR/4d4gZKZXOS1zDXg80yqUo53O
woUFbjFcSnn4qAsSnz8cmb6BbRzxMeyIs0XSUoKlTGeAMieDlZ6zY7PoTdKxQgIl
AFp3suknKVmdwqh/PmxXE2SPPS5AWY1JGXozYFjwqi5jOx7nQJRh1FRrOeqNzN+q
3Dn9DYnq4MV7dPu8KoW7rzJuC6V1AvgVyjdjD/OrDX2kHUf4XBGDh3eTR1B27Ddd
IkEHB6Ewrj5IUTChq3xKtl7j4Ea/GDd8Z/WAcCiDt86NapaDwrf8NdyIbqGqMhOw
KO9g6nHbnY6ng+NHkQQCNxNDsPMP8NMZBYz1P2tUgF8sRSnNaBGoSuJ+CopR29BF
JGX5pn2qCQEilA2mHxiFLtS4XbTC/U4/9WmrXc5mhdJThSCpShtN8xkFlrGN2aep
c9F346nd/mqToO7EuOFvHebo+Z/dbNGHvFRYjuMg4si/Wm7ucn4aVyRmWYhGdbfu
5BbRpLCnNxXqHYVwLK2mB1dRM/G5xqB/TgtZNbvm71JQDniEjuKfwEiIMJJNGVO1
35WI0w0mGpmNSPDeLMhCpwEmwprQClPsl8cXEpUrkM79ro8fiLIgPnWWx8CwgWjW
iXKtLfAbUV1Enr3GaKjUsKSX0ioOyHG85DxxwjNMILUf8639Ii+Eo+Yo4USX/yXL
WU8hY+Lb4lCNS7Re6lSdPoj+o01MQVOMBelkFPjqdXDi6a5Nb+4OFKV8BPfrJztg
x1EWUWpM2PPvGiqdXpwj7p5FIoPwB3dUuh4oS1sZLgMxHElsWxipf0UAgQYQkEFD
c4Sxq0l03tXuA12qAwdmiNdb41C+EY3cKRMFEpOVHY89KTCE08e8JUE+RavsVRwl
Ntg9eWfldSz+QCYD52NkxSeJuzdoOBl14wQfYB2yBYeWAm9y+zThXsiJCBd9gZSU
FgEfd6ECs9wOpHtqvR6htpQISCcp3TwXjSmVrMepOWZd80FPbM1XI7v6HwrMz5hz
/BMOcozZ+vrdTvh7OKxXunpSbbTvIWOtIMVxwAbgnVT28sKeiZbZrfH2ZxD2/Xjv
Paony7HKcdS9FW4oT2UwF3uYeVJiIXJxSyD6Kdy6zhDUwWnTHU9PnMC4iKCdi3Lg
pBD1xPcXZXrhd6hZmV7r8z4wg/XdKxgJ2J9KMcPlN6zPGXKrApm/ZsgpgVs8vnsT
RY5cFRI1ZoCs8aQNTja1fKRsa+CGmtIgXSr7VKmK1CGLw1BdHWP5WJZRi+3lCTry
KYJx2VWL6Ku9/K6Vqw9BL12pSHdRgS4Yd9yxDdjZM0/ONdUOto11/HPIfbUxH32I
qPsq7+v6ArQsYdSzh2c9uxQAnecEIWMzNvhIY2ykNhJYAIu35rrDNs7I2110aky6
bjbIsnz7aRPkfU/VK56aPqlk6+TbF/1Iz2yfUQrN/DT8uEACz9oKv21nzEXSEI1k
mo1WD94u2Z5ii+b01HeThgqWwo8lzu00srENreTQGUrHCgnb7k+HMmX+XFB2iQ36
iAA3THbCkvlgfJ4ZHZmEtT/Tjl7H0LmbUpyuQhs/6omU9+dASsKaDlZLELOZFpSU
lUjnl4pxGg6RXagzq6UNE23RZht7GUFe3f0+i9JJLbcZBCoff6xddnikDUuFnhmW
CV5r07ZgJ+IFzxFoPm0KiSBbgDyTdNC7o9EdoSE0QDUJ0a8nsdFVv8SlResbDdkp
Xd6sUslud1dBsjuTSJagX/r2HmsnUXZpHuZOolT9XCr7dYGv3B3nZUgyJRc6G54z
ybph0aMzJTk6e4BFX4ZyDnHQIlwBiXYMrtL/oFhC9AA8ipjPEKVOychCSJ6BeNWy
pscvJMOqvjIVg2qUJxG6SID1VaUULni2IFd5CRiKbT4HXq63dIpb8zOGTUyWBNPD
EejgeRGEGGBn2r9ZkXD2N/xYw+0ggAoNWLU5t3ao1RgVpoFTu7dx/7Ys3Bepz5E/
HrZfuXmqP8S0Myast99RK7YPe0i3Xx/rNXgngwz4E0HxM9IryDHGxJvs7FKx/5lh
YJcAanUCOmelcPnGa5GR5iIyUtefIifYX7fh4ah36aadAePCjpcDI9N4w/P3SlpS
fJXa0mUlh+uMNW4J07NjpqeYShvPWnOGaQUNbIK6c5e5kgeNhQOrBqfrmMyCXeWK
OrSo9ZBjNdz6GsLttjs4rKLy8HwH49BtsC9pvapb3LyXarA83dk1bcM8Dwko05a6
JupjvrOCr5HldThSRnRRQxNlICJxsx91vdFnOi+DgGlij8i9d4Tp6xVgbP27EBbF
7T5BqmRmL6k+LyZVU29Eeihr2Elyj3FU+nbcrL2rc+/wF4aQjqKR1Eb37v4Kr4+N
HrkWNl59HIOdB17SpVbjsUFiO1ntFO1m3Kdde2YrDE5jYlSXOUcHYak/ILFphP0R
yUkaDZbh/1h2fMSd8Mks0Kq7JI/k6NfPlVEkrDzWLbfR+wFNSG+OftHMVyfENOq1
a95KS3UcYRzkX/9rE0helxpiU+4drmJ52iwwA9rDeeeZeo31f+40GD/hq+Phf5mI
zVGY48ZseFCqI5KWgHeRItm5wrcy/X+wpfDc5tqF48TjYn6RRZWOvWMnP4SNBnqy
SGmaE4SzU/er29CbOv+mSumlGXk7kdez6svveWhjF2ABpHYmbL6L3lQSm0i02WxY
J4MSuROIU7czQbkQXJjEpQ0/j04FWmXWy69ehZNqX981LD+ldnTad5Dvp6UlDaF1
YZ/KOMaHhcOuivyjGXKlDKtnDsZXkcPVrqGxI+kwVfreNK/bat4R/aZ6hefOxEud
vkapK6BL7f1uc+xWrx4X2COm2sg/tkGribi25OcPySD88U/Tu4F7MhETbBmsol0X
a/23x97cSNooUOZeIwhrR7rUZ5OR/XhnPmUAnWVeT5a7xlTnbyiBdJ6V9yhcpFNI
q683Ioduex8w/b5h6QsmCT/YpnmGD+B42L2YpEkOVS2aHUpYLtvLxPVV56KMYp/q
DSqE8PPodFQ5kz6jGk9YUCbOPqoVCNqr4MqkLtKikeICH4d1LieDe2h9TlHZXcjv
F3PNS32Cl2KgT5FSFStgsLp9FnXDM6GMqxyN+jQIcg17DFmWiPtbWl14JqkoGuUn
xDGimNrnuwum2FiiR5hq+AnAzrtEWp0cD8/A99nfe5fN5hlxFiU0CPqG7eiMKZDV
zY+lISTaaHwb7l/lPiBmjUGtf7RoY21yhD31MMM8nWrByj2pVwZ1ZTuN0yGeIsfA
1GjlFB2cjx6H/V9uR2q2lqfrZYREfIFMT7bl6Zlt3Mvo46+1sLRd2MCnaf76zVrL
YFvFGaXwBz8vH7779Wgu3ocodWGhx9zwA4qBY7zo/olphTESh2fbwe+63S4kossw
chKlX+29m4lPz5WnFhhpbHQMQH0CmHYK5TjCp1MUq200eLCzFTnP3a7QKTyMNPP9
PryNuXnhe5QoZoV0FH2EYAUk7jEVqNiJ2gBNnor6A8BrnDglKsgk0R21Nr6z08jx
8v0QJ263vQDdP/3hyof3lYLo83bYiuzW2kfqoQiNQNQeSRWn0IzprspvSD2L6Hy9
CLNv7++t45lQOfkhSHjNHNyzGDoWq+q1Yl9ooQGHnC6huiX3iNbB7Mz9FlDmd1bZ
1cIvRPMTGrYJbYsCi5acmcEN/khc4W1z62P77npm6tI7U2PFNXsH+Wif1UW5AvXm
B8LGElqnLjzaUtVFutoQM76Y9BRxht2p425tbs9dYRPalcsFmfyC5cktmwJZr+JK
6GWy1dzYu1OpRPGua/aAEOcK5QVpcIIA+getg/q6Xt4yXfJ5rJ6f3zbL5jEb0Tfz
XVS3PdLL44257tSkdJ6skr4iLCgsjkcausSxhZXCGsCZNoFAvENR4ckI/w9skHVs
9VgXHb5zG+nZ/NxRym1pNHZAUgxZ2YsP9I3Mp5YHKaq+muglshnaCB+ue63EgdfT
lFKuJwAl9Q7vmfh0KWlv0jq2RyKqlrcudXUcVROArf8sQ/BrbOQ/rUC5laN14e+A
l112BghcrehCYg0ZWDWXuE0U5zCqPWKIX6ZeFAYi7eAZR6+lx5w9nt70wspDw0ud
+2ljabr5nXzE/6l03w+AyyWxhbiswxjXo2+tKIb7Nt6DrR0CnYRaGc0147wvLZFR
ag93jsjTj9RvXIjAMSk/AU9wN5WMCowbwIPsM1vhAWOHTQi7MZz8VHDHlmryd7fA
E29Hv2nmqgB83RXCt5Mrh5B5Wkj9cX2UyWgZEx59l24V9/fU9Yex29/2f3R7BPik
n6AH5SogTXUpJsy8vLR2F3E4baoY39ve2wWWpKaNGr1DA9bLvMdgaw3nrpAQWO2T
jUHKaAf26abfjKT0naEG/NjYFpgUb4pAE3Bdts2Mmx4wQInVJ9KbmJL1lCbFCwN3
kmnVsCIflHffvq9PooCbp+vqtucELX47lJlkQLvHFg5a9+UKBKcd4Wx2gnbzFWJD
mwIBJbJFO+ci26CQW4NA/2kydLvxPjh2eW3gNrpVAGVAOQhAtzXGvQ9xh0Y2dtxj
yKfVmoXo74tvpcin/iqAfomYdIBRGngkTOYnCjEh9XcFI5KYTvrlFbAX+HEEPS26
tenwOGTrGf4MUv2Bvi1bhIqJY1Ja5fFslsTXrQBBBb9g7SzHB5nmtQmsK99UNCRm
7rXIBFjNqwDYle1G/120BcMtPe4g5FlRTSODQ6TCL33fMbrDddcgAZxib1IgD2Ca
+SElxsndYp8Q+HUpDEeKc/i49r3C6ZUwhWW4Wkuusc2cyV3K+eu0QuLMW4gOLvq3
Kx+dDAj7J8JW0Fym0P3pS+Oqvvu/9p3E4ibioHbEAyLbLkOt8qBArAB77DC/LNzo
lxXRbDSzUajIL7vE2PPyoVYrjEzYscWE9LeToAxPaXxrXLgEGk/Ez1MUHJ0CmL+v
Yu6U6UIIbJluS4Mbr93kOhZWR2tp7nQSBD4vJybpOKoWUN44g7qotZ1vuDNAFNoc
+P4/G6WniuQ1XXfcZJVkx+SzD9TDG0jZ4xXJC4WzOEGDpeufA51Klq+cPMe10oDI
c9oJqvaMf42+MjvgPe20sLszJB+MWSPhKx1MqzR/d9YDZEYmwsft+cHngrhN7jNZ
yd67BoT8quen+4i0jqgH3ycOP8ogl7GKMwZNYa7VuBXTILl8WulkTzBnNdkZKUay
YGpbH4uaqNOB73mj/vHrrteZ1nefHusJM2irV3WzA0i9UZeRZIgJ2d7ol6Kflb25
gXPsvFuPh5KBCACWC+EO+QW8wfgR55BZ+GOxAGmiVRAlwmJncj429hslzP8DT4yP
wkAUIkpqNr+VcxiFz5BId3CbeSraXTX3CgexYkKh1xelFmXD0F7dd0+hHQUAb6ma
/LW4CRlyXKZuZ1yAends+oY98SndCcwdmlLcHd8+rGCfMf4tmzoyWhzWX8BIugjh
4NJEtvkG6bF6SpnYLmKvZXtdHPAlDGTJe/CNxbeheaS+4JaewTZAewBLN3IwaUJK
q8qz1PZUibUZ+OWdhcqH63UFACcjCOoopzKYccMSYh9G000y9JX6aiWa8dW/9wIG
6FGM3P499GODu682FDW3fagB8LwYEV8N1eW04ZUGwMhY4YnJh5Y3KhY6WFCLyOcO
iw1liM3jK5O/ir43ZJudQA7kCMKvAKeJ2crgJ5fdplihSvqINbVB2mKdg9owtpkw
fJicQ/QN/M/N1xWcyMQCuCfwpvY6tHEcb9ys1B4WadGfeUDjqL9wP0mzBLp/+qcV
hIOD5M8baWmRS257TPL7mNJOUtZDWELF/lqDckX+ZFzZ5w29rVs1pliaHCnD0Ij3
v9RSyd5U9QdVv0H28ukv4HjaJ3aCHWgfyqMGs3Wn2aR4PLw9ugZmaXL/tI5C1lBq
K0eeoY9Fb3J5IjFRkFUQ4tXODi105BwTOpdxjGS2mCNthkJ/RkqL7km99NfVJ7YV
X6rxW5CjSFagCADkJfkl/MzxaEUuyq30WmxgsAltdOqHEn4gUKAs39kc0HrPfjk0
7O1lePpBj+RdPMRZc0J8zCAZqP+vrF6IfIZCsyHBu2ZdRSlo2bIGDm3TdNhEtM52
gv2JZQzcaT0R2CwrsyQQlfrFJIvaUjld+agyohsGdU7Ab8NXP2JCuZGjYmWvZnZm
P1h7yW9CLy8v4XzlHzfVuL/+vxvY/Kb3OJFlOE7lbJvYaWSXQmLiQD37MwL6rkoF
FraLunEe6HTccGDY8T1lYmKA7dbe89+3NruGNR9QYgLWmOoc+QLPRzSUOSIn7cNU
/rJRjIvr92GC2zzMGBewgZYsLNa/sFOCb1F3NFUqOtQA7rWMtvtMnuMmMmIcMKCS
i76bcZXVSnp4Fd2QDLBPMXQzKo4xDjLJEO3oWvN6nZ+QB//1IK8vOt/sGk4CJCWq
70gy8IuiQkDWPWaaFu5ikdVlPDZkOpWOvwqYNphCrjT7Df9c3so/ZhXPmd6rOElX
VfqlLrMySuvZeIQ9dTnUu0s1CmgnRPlT9WM1PnYwRQX7NCDplq7xRTdQc5Rs0Zxp
CA2ptPEjawaK6omUa+mfDp1bnojcdROEFvVPg+Yf5pXjtLXhTIVeZNEBANjHDdlu
sxr+UH6f2G2Bj0vyhLWMAASgohlS/IBZGj3CocWSOB0x++vRvTGmajY8XbTwnCsd
tVKYnvgnqCGfKq524F4Gj2cLYdB5d9VZHronT6Wq1e1do1UoJLg2D5pAADwHDcjJ
7RkKSJAPMikRpHHsYEvnNauaJs5J9XdFkB1PUWjXdo8qdNPjDJVWyoECF2u3t5Z5
fT5huZsIvn2x5xMpgFufh+ciaGfk/CPopHp7biYBpaKPKYUaCHwtqbKIORfE/s9B
e1ENZL+5g4GoAz/rnudkQnnAfDxYd4/Pkk4n1CIqt/7o8ebV0vbOuz7vVDcLrwXt
vftiCRSz7AUKDHbAiO7GiqXl1PWqSGySZB3DdJjDWNicGTvSNzLKONVI32LKRO3+
vKQy/KpwgYs3ca/Vttt+hAcgsS1zb8lWGboAVGJsLGyZAlwFkNylZuuipdQz3+kJ
Lq2J3viGwD9teN+peYtO+TwJxqu1xByhj/fd3c4Lu/ex4kX4oZ0r777wOXc+iJ1U
D0PqCa2AyJT8cTrydq496fsM9WtG0aUpsY1E3qMrQlqXH4ZTxUBvojMd/+7Q6faM
sbNmmvJdfFtQzQvvTYj859/3KhNHqwIvZduJBEhLpezVq/xJtpYnmm5yi7Bu7PUp
q0I3tgofISE1SZI7IdZtdJPJ76MvyjDqoIo5gkirKCRxdgb8BEMynMCXD8LAT1GC
zZLhvk1/Oaa+ANwfqbb06kc5NfX3RZrtmntEsEUyM3BHiGflFnkCqewuh8/nmzvb
kD3oZTV0cwxcuADOMe0SQ9PffG1zAqACF990c2yaPI8IELdiqENtpleLxsG4oyON
cWcrQUw77/hkgTwg8URO7Z+sgiqHG+FwaERtJwbIiQ+pYoelJsw5vho42LFKm+Gi
7WX7InczzNR68hJ6f9b4ZsKFT4GGGUhcYpdbWgzA/9jIInPZUfoFwCFLICCvxdn4
Sqz+vhkoXO1HsLPBwPaZjBzoBSozi6WESEncu/aB1ZylkADgRDPpr69m0epH4hWh
dj05zvjqdJEHSWnw+hkHKAuysBkL0quTtZSHT9CvNnI8Pd5foCLyWrh8Exsm1j2D
QDMOcqIYK72HSwQOq2+LzaIMOQN74M4NOzun00RY1X0DnuET9cKVRcTRkERBcp4q
Zjr6sHIZmcBztr1DRuLdlGdlJcNITDa7Ly2fGJzeOujU6RFCUNEbbZMAg0hldXMl
+fj47dvHknJOYT7zt70Q0G0C2VxhHjapBSsQJOu4pMlqFZUXElMuo2LhZnfazrO1
biNV5/U0ndztMWQQJcA3S7fVBHl5zb5EUxO4aPUezqhNZep9qL5mywQJRQn2WSjB
EJ8epdV6grN9+JIA0H1RoYFRUuu8KoYFomrZxH0PJApkpSKMmD5p8iHU5Jz2pBX9
A5ZIsxTq/ZCx4yYCyLqVU8PI5IkCZNJjjmGA3KIvzV5cXgU+K2XPqslP4Fv9Y5KK
Vl+McxoI3J2HaiSgCspS/GEyNjv+sNA+DlpvQGAhMNkmjwGwbToJscSq/4W0IU0i
mOOl46NfLKN93gDxrww7OpbBLBJqrTEqLG4MSE93jZOwlOLPTFgkWDFyu8wHdiIJ
51YuPvIW7DwYvZnfCkJgP1F+VDPpZRkgWsX2D5xDZRQg+4D4vfoxjSG3KD3bIhSM
mYf6ZlpJiPFhFbErJuNNycZWhYNVbi6iZBH9PoI32D0B6zv9qADggdRlyzABNLp0
Joe2qBD07RMii/27MsNShciBdoDdD8AxuvY0kgW4YutDLyXdNyxqSrRxq+z7wOnh
9wshzxzYg1p+v4XySXOJ1kX/iVcfy1yzDBQuas4TO7eLZ7Bh1zJNMPCIzEppfNBe
QUhxwWQGQ/cwiHRAdXvwK09ujeLeKON+0Y1QTZ35PfXKEz2ohyS02kVko4hek9Xr
NLd+9qS3vEJUx5ZdPNPqyxpkZmO4QjjnDTBWZ8muXjl92xuDDYUoD03CkqrgTIZq
8VxHH9+ol8NgyZvcqF7/OUYmIAcvSzGktDUa5w05yx3inXSD/uXgtfJlDmF5Gf4Z
FwmK+Gr0DuD2qvEK+ZQOOWkGV/RlqmWNTB5EzGEeYrZnv/pOFPUo+tyrojJHiOg7
sSVr/35OV0/LMdnZSsjf2uDYoSnCecUo3cvo7QhIboJ40THtXYkEjtZwhSg3UWjE
CwfalX9XWkJgui3v+uHT3t8vwrvgeBipn0Hn+0afoF4mOoKTwpnYAJux+LX/nyMZ
LlfkjTLof450FwRb5QA49bsRFsoe5rzBnfjdFa0R/nvmD2utrhMlUzsemEptQlwe
hFmx6KI1xaBpzAyb9Cben7tfnvtrfvd/2YIJXIZdfc0Hv7sLRS9IUvIx4wr4j4Bk
EJB7NRuHx06eb1JtuWGfT0vQl11SD/4aaRUCPmoMUmGBBRWObd4ZmVcYPL9M8LZz
poSn2mgW0zeTZ0htx0N+1Hug64deR82RTBGeXvoh9WsqYzHWC3AsGtkfeP8M12WX
IY+TB1Li3C4lSKC8Gl7qcNrM2598Xt9xwI4FIjezvVhT8t1sQNg5DFBpOxZVoi4Z
M2PglKivXDMrz3IuDrnDS84IoEvx0qe/2HV5CKBEdpxyFf22Tp8mnlbOl1Aie0Su
PEi7wgAl4sa87K+v7d3IMkUNJ/S/hoQOMxhsaqdkv6hQYqCEHt3nLXQT0aD4kAyE
+wKL99jaO1Sp3HiK6E2gMZIEcZB7AC0t5fkrCpQV9EpjwAYAcGyosam/IvgBitaZ
rXmWt5T6jeI68hKHJk9KWg0wnmdJPJBs9AoToEFHC+ELlw0eQr/1GJstw/mUz0Yb
OCQzk/gyMKeBn3JBMKwaLfNdmNBxm4ktU7AYrnb3XTX30bqQVXLYnKZv2VaO0mLf
/KybdO2Tearj4cRatmmOjTyCkZ7cfCiU82Mrx+QussCatykzLTejuOotIUFpaqtg
mqsflwKZb0K30H7lR9suajZ24yv+KUo1J7jZq88qOJ5V0XWplKRvY0Rz5ldPbT8T
UBOiEJ+mARztd40gbOeQMnz9XKeFtvmduFhJ3wUT5gKAK88qgYVa77eBFBA4Nc8j
+QDSYcScw8YdjfVPjXh7lvipEauMIQK0dpf9ShiLvMD8HLUeBxY18eHZhh6aQWDS
dNsELVCLBv81TLrdpbcJLh4mHbMTrI883OdjywlpZgu2biIeb4JTvyqnd6dDwuRR
YKJnfVNooHzTo89o3B39McZJElqI9/E5DfOfOytyu8/twGnRLMWXWYNNR4x219jU
ybQY0UOWjYss0YRDjDUjuRopL+yxR6qFbGbLIIXacf7xXBLHWbIDWUeLpO5OLHo0
lPP4ldqLv+jKuVKdC5c4KtYg2YXUybanQCBC2KbFY4JBNUVskeMJ+nLvJupJYsks
uFEoJAzLPJhkX25xo5b5ngs4B2lvxaN+wHSo/dkIJQQo672mWdKy2V1MwP949gqh
ldrDXRPKv6Z8fKJDa444N2d236sFoDEUKiW9d3FppnnUzqznzUFzjYE1fwtxUyD5
3EnN2dhiGux2EXH6GvCVUF6gAXPptQI/4N6lJKfoK2vtm4Jcmx6ZQ8itVsYKiGIl
6vg/nYTJcZ32d9nDpYvV9RPtH7N2808DVZyXcThIlgbrdW34xm7jdZc6F83kPPxQ
R6xqeRz76arAcNBIUYl1QdFjuVMEMgsgvB4HAFo2RSd5w/5kVrPR2Qt9A32NVSMl
YCCac85WuMz0jx1ZgAFua33OZG2P11VDtS+puZese3NV3YYRTayEYkXwAnmf4HEa
R0WzRrbz1p6mdDMgEa6Dgpg5OhRxx2yhpiyMM678lCsa/ft/meujy2m1pDfoPXPl
XHnaXQw50isW7HKcy1TDPZzB35nwo8tSmLL8qq1d1/iMSFDIO8l/7ers0nQd3SIp
UJsGaj9XBokicYjEg2tAf5z5wCW18d8X43xXGgFMAGkb9Alt6IQokBSvPfJ7wPam
IOPH32Knfw+tORbkCggqI8DwdaLnw/BPQWh2mKgMwN/ry3TmWadpfrxLHU5XwkAW
2QRsVSNMBqcim4FmyVltm39x8vfw7D4lNCjGBPzLNnxeJIJPFvOE4ms6rZBd4odj
SRyJBzmPcDw4W+vdae2OQAbgbxJv5oA0f4dG5A2uudPdA87DnHbIlJjeNb2NVp8C
D8IQjdZLNXKmGVNFg5TBISPA9sJVtRkqyDcVipHIn2L/eZ6xn1bj6J3OQcKqeAWC
b9b6x9m5hOtf9HuHuwGvPDrghgMIugi8mgHfbMid4ZFye6mPDuxmJdLLfFiJ+BC0
SublPCVdJiKrGxbw0hYQ9qkEnnWbRTBXvLNWJb9otJEmXqAn2kjkSxkCHwLdtReo
c9+B3dlK6wm8+wuHKMFoq6dnjJMgDN4sDZSwBGaArBrGShzdUwz92OlHuUqPAFsO
9ZtFjRgRXnUtqf0n6yEvruVtsmhGOyQCStJFAavXiEVkly0YwytaXHr5Q5oL99Nm
IdYxS9Y9KR+qeQPJPlhQEhfJrgXw3TZEuWE7Rfo250p4BJDK3Z51WD38A7B90hch
i/Ec93OJ4KxOA+kgK0hSjIc2hk46iZuRcn7QoWTl57hCxyJY6yYnDUm4umSXdmQS
byAvLw27+iOyhPxB1OeWtliLZB0AlSJqd3wFssCFzT8UodvSHW8gC3JJMIGIGRXZ
SxNOFxI4Q84pmJb+FUP1DQ01ifyJheuF548BZddDPgei1BTIXs3xcrrYbrA5l7qa
wviXOkzas4KHJjPtwlamiDK0gpiFjLgCA3BfRJe5LxwoMmw570HpSmlgxs8Un+2g
7x2co8Gp+HKB+5KMoWQeuBGXpZTUWtnAE2uMYdNOE2ptUNTSuJl3Iw+PlCluU0+3
DwuSIralgXl0+VlIk5NFfOT3MlWkQHeEktTpNErHGiyYWgXfNKpWSsmofGkz3qTw
DvtoTosxZg8P1ivLkPCACt92uRUuwKJwSTW19EY+o+eGowYWSGk+k9k22RfbJbCo
F5n3h4ADgZmfQbUp15sM1j7aoS90mdSNF/Z01GbrCmwt9G+i0v2PbIgXDdrfy+nt
qfcz1InJlGBjtD+UIh1Havli9IRIVuctHGTxPyIBIM8GbNEjr4BFJrdH1o8bz9Su
v3Pk0C6XyTiWHxoV0VhJNs7QVm628B2YGQ9oHPHdmYU=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
msCzV65ynbHW0gRT9nHBdUIDTWIn7Tm931B4f6Ux4n/d/jopyUKgWMcSVm/qaL9D
qUxTBuf4fI1YmYlIBTy5gCJx0iF3Hood4MQGBx2IlykmmGPSUaYuQTGU3PtJw/jY
ScmzgFTRrAUZIl4LyOMLGUecWG/63/C8JSXIQkQV0E0Vo9flKnSX0SNlqaY0Jq1M
ZMM0w5l/40d7XEkmVFinGn628kjmndpXgTkYtLPUIp6kZiiAvg4ywciN3mRC/480
o+slqEHQcROqNTGqhT0m9y6E0r34//B6vVqgfcci8sTYK06xRxyZNaLVwfuHlm7g
CzUNXF/zQU1nw9f/NLX6bg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8272 )
`pragma protect data_block
tUeIbOb9euADiBTsmrsdZ8jRmo1FA1bVxbz/FeGurDoCPDQTqDCZy0lT88Xsq2kf
NZXQPKQQrrg11XN4Zg/HtZYgZ1T2B28UwaPqL0d+SmR+rEnVinlKBmwxnWrxOAIc
BpOEQgNg342O/NJrD//fYHuv+2tPkuCJ6OgTGxq/mm+pKfxyODeLau+ALeHU34Km
YFjFIt4j1MUfe+5iF8PGlfuS7bdcu02vSxDqsrq3Symt2ZJ9QrXb55Ob+UYJNO97
adLkfNYwvlrHzmXe6X+UEmR/sPCsy/g5PswOHBzu2c2LtO3I7HLNHEvOvbXjUPAC
1H3VBXv3PEhw4Ens1LLtzZA//AJwyFPVshFh5ZRXdsy8t0JxvNFU73qGj2yyGuG5
QYd9TVKOji4zhM/IGmYibKjWd0d2oEMl2QFQUxa6+CMVPt3fSKKpwLqAIH/09zL3
DwQtCU/yoyR/f696rUBP0Fjlxv4aP+4ivi+Xq90G16+wxIp7IRe5ppXw9Ul8TCSg
AXSoA/zkIwKWhp9ReGbkDrqOkTIeAnxreSKeHbM9w+ez4NNbmtZc9Dk8DVbw23yC
oRQFkbJhYNhMqU020f0/n7ZLEBDUceTOt/NTQ1sBuxHpolRA5+pDwptoORfsuuqV
LtSPg/rGtd5Me+ewDnO6XMpW5/sC2gqFn9gzdE2X29+cLWYzHV50+qdjl160gVmS
8PgWD5tNZoXa+HPPbG4XyQ7LmCSRGZ5HHBzvgq5CGnHvasQ9Z16KkcZCKzGKE3qL
T4REnzNDr4Wp1eOgjjO+JfTU6ToRyV7Li2ZDAeOpF+PnUScghanwJ1fu+87s5MnW
+200OJ/jyeNKVK3LoWPDsNBCWltdYP/i7AWmkU291e17/Mlq3FhvHpYmcDgvbi2T
jUBLimOfUeIeuocaXOiKXuj4yEHjh6oRAbccBvKM6SplWggLfWgzYBTisunQA7VY
7w/UzSy+UJ4xPWbI6ouvXIKPHNqCWxjqUddHLi7wzfDg1kNosUJi797jWpmYN6ze
iE2vLoDxcmURv0+11f8elKqCHQ6q1+ErlK0FBK8lx0WKlrvivl2eQ3puRwk4Ztp+
mtv7u2dpbhpsgUEhbvCcZ55O7N2DYMleMJ+Iuo3sIMcJ5arY2WoKPDbmNGSF7aqo
ZSrrxtlkxNKE518MbuGlCjZpe4kR2MGUySqDtVYrklIsV74j5YZj5ToKssSFht5+
i+1eVlWLeZ64mIs/4nqw3SY89BjKtOTcMEZ5PYxIYpPEqJKRxHnOZwQlpyFZY/t2
fDVTn70RGZCtSNK9/R9BtACXTYRSoxn7aogVIKzTYDYNUm1BtexiENtJeXV0tSzD
Be8+xAzhIMNGCCfliQgxubZwU6pZL9VovzTFQCWSkUm14fLtpkYw0Tibg4FrOTTs
/2eAlFBMZ9MN7eZn3TIybAGJKI92kXr1s1EDMYFRYItEd0RNAyMJkb/IfBJispgt
4XSrqsRen25K4iF+YFv9GOdKNR5TBZdvEmdlN+xn7PKdugfGAlG+Ok4EhdFOr2id
h5YI55nTsE8efVT18rTtDMPsN+tVuo5Eb1H/1u4d03QuuwSj6mkcz4zbAru8sCP7
WQEtiQxrusrJB6l/+/MWhzknFO3RfKSs5KnYatQbu3sYQ6hDPqyvOOfoneV9OZWT
odlsVx8dTidbO7TD1bPl9sudEf7WOWz4kVDVUV1g0t7k/xRnYE+7MZLp+SGTf/+S
JWff7HBnpMCOO/4gX2dwBx+APHK83OdWr7pI269hdkmEfh/2pucGQQkneyfFSIwf
E9mYOrruBYogNA1gQ9+4OLsAKKLFKIxgXUaLRkt5x8zcvyjRCJNlC6oNCjb+ubJ3
x/CfExJF0DeDX5igrc3DgF+kZci8nH5sr9BBYsxBXIZoKSZvs31iB2Hy6F4pBe+Z
9aHLeVBMgixs4sakXM1uGjMkdgHJV//A26AGYJuuH7E97YCitTB+DTSiLku6uT+7
3EgKJDI+Ke7yOBD8UbEMtwCQNfZ1w+X0rXQcVxtkVT8lSU1sUSCRJyDh5oNLxyDM
D2Pku9WPf8FBhTMERiAn58sOajWLPtzubCI9nRd0Xkh6VotbBuYr0w5alBav5R2/
QNHP79ZPn26HWK8BimP8l+SomVxeuZSd10eSjI9Tqhdrve4Fxb67LkAA0YmwYVqU
LCzYX1tUYsA5PnlQ48RjiUvQeB0tXxvL8qlkOYoUyGvDaIJLaLwb59kM39+JuNyq
pMiOEWkoGmldsQt1XfSrcKZbDG1BVvJnnxjKrogP0p+VNiAh69kLOOchTvWF5D7Z
4VR6Q4Zp50WWEm2/RrFPemv9OiJpvJPSVARbh/RhHaDpRyDqFNqlr8RfSMVmkz2v
bnGRdaII70hTmWBsE7EL0c21hHTfiKCoCOpp7wnaAMztG0iuJJ4gdYpSgcCmgRKk
JT25/6tikJlxWAPRuGbR+YWVse0o/Fwxd0UE1TDOKJIYTxWpPgPm4ktmWvmEulTI
OmiOR03O45n+0/HCpB97V00d0rfFnzFVEZnKtwQvt4CbBRlGT8+7iL2sRBONTpTY
R4ChCqqJxdJkGY0Q/QBwtD/Ryl0gT/3mx4pSWI95O9Upsx/oUZMicfz0GHEjcU+p
u/PEVz6QBqB9Ul872y9QLW1jClN22kM6Z9CfrYVfJqjUOor0uP1kn8MJ7gbqXQYO
QFPk6iKVyhyRVImf0plDGxtf1he/ObT49OtVV9caegnZkpSgbPS0MgEFSCstme+X
BwCOraWqvTIzlVXt3Vg7oAH/odHYjE2+R8adwI7wIbXQxBkIU9Dy1Iqbga9lzFmp
Oiduw2RkL4Q592zLXzkKRezrfGuaMjzW7sTqrOunflBJ9rM2LHWUIKGNq5UOKAo9
HhFXBunimE05vyS0Y1vXa2FxVW0pTZE6X8iURndSVSGpvILw8yXYtX/QrqlA1zhW
uWZFruj7OQ0pbwPJ/xDEH4AKEy/LP0uv3A12X+MxQXHrb1IJVgQUKA/1TCEa1ezc
ic+4J6rELPbEeaQKfXVErwB3nVpXk62D8qFE/foqUPC3xqzgJi/AZYVl7G3vLHlw
RfNpKSiwATunVd/Pk2nAztRyMnP5do87qAgFqelUwQATdVjsbMfel6G6Yx5xk8Bh
lEvxhS00RvJupdpi40L4SdzVEhiZ9NWR88RYOFwj7hUdYnKt4gx/VARf/ohpzYQM
1zgGHiPlMoVSfBrEO/KQ4soRMA8HoaFF1sMyw+qK5T6PDQMBIXeGcXT9e7Y4iBhU
Ue4JFWqxkpWqVeRazaJfQQPMC1mwVByNlM6ZY2LE4tosmBcud+WW0PeW86cTSbx5
DabFsssO7w0xGW2kJk47YC5kAGCT9B43phBEWUia/5RaoOHr3vB1PjBfIKMQjy1r
TiVzG964SVNWA9OqH6/tSk2npz8+MH/506boMtJUkGCbfalDvlKXwXLXgeE3MVx7
e3DJ1RPem2WtCsC6YTVhr1Rj7ALTXMIrJ+DQE/cgh+IKUWLcS8yhxAaVIky1p/Ka
j850/HlEa5QFYjYmYWRn/CNn2hDRduPRhgk9smzHrD6ucqtZy8taDLxm2fzy/mLG
6DUb6iynm/67fhalvTX0nalTE3SV7X2pTcjZ1YYJW5Xm31PxrhVRHW4yYEMH5D4s
8pVOXy3Y8ade2YH1ZhYbHW/7Axqm/1XmCJL4yomkN1syuBVMnT1FUbex71i9I40b
PddS5aVbGoX52tvlFfxqwgOuc3fAbYuBfSswSO4+/M441cEcmweghlFqStXia8Ue
w8SYbv0xJtB1e7ZyPe6/qOZbGqSr3+Jajtc6rOuKdSaYivVg/KgJ+uVCgcSWc21H
YN0g3hKhhR/qXqScgpyLq0fIC56WMGZyBkusrscHCAhcjiYYzYVa+2Z+MSYpILmt
BOyDSVuTvGFh7z9jvur6yMOeljspuhTqajESZhK4MijtKbmsLXwHMqZ+44G9rEVC
H+sC6dkZC4CHRZzV1chilKo53vhneUtAzg8W4DxHDKYRhs+zSpmch1ur6Z3pH/N6
Ncvf3Pf9YoaBvXMPX4SgDo7dZU68rhJJgEaFssDh/kBuh8Rn/SIgFKN/KCRwpyoD
MwmJ9+en8kCEuUOMMCQIVc+CVThtnJaoMhWPnSl/dUw2MPRMmqqyz3LCm7zM/U2J
cG8+EiMXZ4kpYz+6ZIZ0oO5gQ5F7WAjvPD3WryVOQuwiUjMo0fdaSV2LaJgB2VSg
/AP+/g2ELKM+1hJl7B7WLYqO2vtXmb5OCuUfbr2J6f9ysw5FiQJX6WY4RGck+jCl
bP7XrZAho9nuj+hijNvTlcoSQHsirNjLVJLJ4LI2jd2jLCF93QbXTIoXBRn1SD+V
9BIxeprGtgXcxSNZ9IE+ACEG9IYblKWvtuMZuLl7vvFpJr5CswbcMsW3SgfmOfpM
Ys71LuuG0BsyBk+cvE6pwMkEmWT2hx5E2aVRKSfr2ZGPhCSp89f1WFPKZ3Lnq/p4
zMKiyYnKji9xMGAOviQ9gO10LH5ZF2STzyr2Kg4K91EN/UZ2SwZfgTXq/D7QDcgT
zaNnhQJhBEzkv0ltyYazg5olube/EL4zlslLm+jF3beKl4j4y6/ZT2nkwoK+HxNs
cPP61vUjURI4jaj4JhTexpa0QSmICGyEwsy3q2/jdEPNd3uVo2uiWs3ajvsBA4KC
Jfw6ImpZqLd4LrUZ3gVrAbZ8MmNDd9NU7KyjpsRIIuCWIFY2DnrShSW+qdJRPdvN
ReNVegU/obbpigLAautiRtnlN78Oq6KgYbuLs+y806dKFtXSSf0kkWWTFxu/jczp
Pmcl0NqcoWYNRuhA61nD3pe+m+2tdkxm06OQfd4Kfmcwx1RC+iYkcvJH+zNEm2xY
sN4h2iCaKMnZDaPEnOkVjFWFD81rmccMvliLa5PsAoUbzzX6AU663pvXt+gUEqC4
k7sLH1Skdge6o6d46LU3i3+UMv31t2Eg597dBtjqYnu2Ej6CCoducb6gJ7Dt90a5
QuSwUp5pJu4tt+HZckxXkY9iwx583LelcUsD40HdOluHKrUKZHKvlr3gc98IJMt5
mBGGljI/k2TnMPVanbsR4Sz7DO/nJ/TRq6XqTeeRAuq9elm7d0yVg6tpO89w17VN
goc9OXi+YAEE3ymc/mPbgfpqkiTH8qP/BgAsDpgWZRlQvHp+DNnqphOslEHV6xdX
aZ3VembOw4Jx/kmyB3Bph+/6MggFGqyFbyls3a5mL+uqPam5RZy+F6lsyw/OALrb
i79oae8agw3mBadTMoaoT/UPEW7b0pe4Rcd+G47ci57uWrho9qwuo9CY3+mMWkdG
0MFo1nymIUEhx1Q2d4JexeOHA42/FaQXLJ3EndGk+8En37rsZyOY9SiMeP4Lr+0T
1EgrjOg/KISke3HEqjU0xYYEQzvVQng+jkl7ShALa3V6RKQAOTUAvgdw0P6KIlLN
6FhZBFZGIK98/YBlya6kwKHiEGUb+AVvU+FIGcTSIMprn1QjLQ7Na3yu3rg76Cvy
RbTsdIFszgDvnvXmXhFr5eSIo+/577g9I38XB2+riDHPsQRQpL1J180oAddIniP+
4uaejU++q5VxUg7qfRHk0AaKV7WcMcs55OZGZVAqvJq7LcykcoTmyPDheMwIyvhC
yds6+aU+LFBoyN1+xWDHAdHGwA+DE/WML+q8xXtOVOg5jjTx8CuTIvssteiY4irJ
fw8AcVrfdJPqGcqUp1hfTWva9Qb+k/nAb3rxELmj40t+C/sXgEXzqCn1a/YLFkeg
tF6565mmKRK6yi07kXthoe+eI7H6BCZ05b15wGQEc1KQVLTT41aIkhtX+thb2NN/
Y3JUikPclIMJn4Rf3MCJcgVDY78p0y6Le+GycJmiVCQ1pf+XjHMCwak9vdyl5PNL
6wsJgGTuLk1WhYjG59SL27VvhUX7xYsaUt2NSooSAp0sHFClcQ/bZLsiN5JwKnJA
27YMyQr8Aj5wuPKKFm+f479LyLBZYJUjNOLTufSc0t2aAMxUfx+SBpFL18h5kx1c
gGTeMsD+bKHSNcKBAn6m37LSB4kfz0YLGm+lC/exRWz1NUo6tz1TSI7RvjQZYAPV
qsX+W5X0sE9zXPUNZmMahJQBy9+ShtBBvOWGU4e1j4n0W1oarx+WLmdqr43TYGih
/mEc0xjEyydUv6DO0HRTvNtNw+XDMqlzN8MYjyt9R5DxmFYMjb3uaYagmcvifHm4
GQaGbXz6qK9b/D2/cCHN3qrKpwVZp6Wr6zOWYavO1gQ+JxUnmioAVSkRHmYHzpxI
BKoyAwCuEnxpXO9PY2kSUq9CXWWe7nIni47yyjW4YttSH/63MtwW37ctbJGmJYeY
3mOYDUHsfsb47qdqSwqCYrYNR0JYWIaU2vZXIhJoqIGm2MgSitfg7TO8DOPzBFIh
W/GefleiQTim1+Jl1TimKKISRHNPrJqogSTR0VhXu9nv2bDdyeWPebHKsn9Hf/67
1G3HbjhXwm++CleY2fCAlIvSLyD1N3v1ng8K/A7K5DfxRMZ1IrV8qAdeBEWAWxDi
j0lboE6BKmu8dxzKJUUw+WTSr9j/q2Qf+GjX23sZt+A9YZUkITR//osGTvPJANTK
BpVNG/awUB2l16KWOL7Tf5E43/Q8Qpe5/LSurSmoh/LDgDkX23UplEX5ZSYQGqUx
F1UN5TxiZ4E6xVmGYEBTu2it0/7VKv7M09cLhCbADN55VvxMyJx25Z1is6EvgKAU
vCzOzgA/vdYFYbKHupeBa9M/rkasRybQYa4fj0oSkQ7Cpfj7zBRR0wrQKYO5ZYFQ
HEoSLttNHWUUhe/FJqgsvCQ4pj8z1RLpysp9XnCZKVB+/ssvdCV6iRGXi1fLoP6T
ji60Sgrw41if3oNQy2fr9aj+zXLPyS7629GQki9Yzf02CfCoUrXziRHqq84zc1+e
vOAfagI9KTOhBA4z73M3WYUDkjEbrntaSGHyx74VLRzDNt7kD+F4Hjr+fB6tn1mU
l3z62L082/uORCZLSrq4YNsH1R4ZhbKLvUElYP+0cyhUIzkpfLM4o6ZqVO12ilmw
FC51Z/W1QXEyXSuPCgsFZSPwE7DeWfMY3hExNjPVqzad41QMlXLZXBL04C/xAfux
Z199ISZ4EG8UaK2LH9O4u70rhop2VPbrmIvJO7r4T6cgwVvDJDoZGphU8FLIg/Nq
ZPhVrhrP4rrkOu7KstNRwHeCoVpwrrWn9NyCkGQeOtnW5pGTxQ+scBdK/CCmtmAd
SqI080TaDSdLvYyhCyr3J4yGG3b+110FQpm07y3akGV6eO1nxv5bN7Y8VqoCP1/Y
HCbK06GeXyeEG7FVygAXyrMl5WyRJ3JSHwJK3nOygVWnEDLzrU858GtQk85PHwe+
QzRpzoYmOrChOTcQgixxRMIuhEkzXdLifFsuxJWWqV0+U+AQy0GkAAa7rF5ZqKSF
HoccfhVLEZt7HkScTMzdf8UzVgPEm/MKMtPcTzBlwN84/Z3ZjRc3RXvxiBuxovOd
IGcwEDh7BPbmWoDkaWcjOljoWfryguGQlpUXHLkp2IFjqwYy6f3wzdJRsrwswvI6
RV+PAv5kdWAL18Y7iHqi1YxMichG7oSoctcqzLdIlZM7wlQlIFzgKo8rh+TFmD2B
ecOsmbQCChQlvEQcgndIjcjwOHbLU3cgrUNmZuN8iYfro9gOKylHu8yLW5ofAuE8
LnY6kjVz++jKcXkzX7SJVC9wKmm1r0eDmAiq10gvlKYpMwO9lSm4jJe43C0yDaZC
rHzZBbZ1b0nrEoIZI37J8RI6xCD5fQiOXAEMNNtsH5ds6T193nYMTcsJ6EwR+raG
cttINPMMIQOxfgeEOVcGqwsQlCaXp1e6f3gCfnLzlmvu0ce20rgo0RBRiW9JEeqw
HJmEZ/Kvsje3wOGsE0EAo26MbHbMjQqAdZSTMHDGNdOg3OlT4TzXaDuceTUjctpu
l9MaZ69lZ7G2KP1vAT3Q8a+clM93nvTCiqCqfAn6BX0uZe5E5IeRkbCEUZqVECLs
KwnNDu2XOkBQI2ilJxmvgVM0jju4+ASCfC1hUl+lZT34WoaK7jzmV1t12K/6IoQV
F2kWf2NmV8V5xKwXhukqFo/whapIybTIurm/pykjSWdoXtTJiiPqdi0R836xhaiy
zlLhlqGSRn0SoDHl37+8wo/ArgcOYHSuszgEO+NRMmmOL1tzS9nT1Z7pO5uvhLvQ
D4QfxdZ/EyzRfFuP2XgMc5SttAFLwxzN59dQRgUUX1jaxesUwdUpWWUBVW9O/HC2
Q3FUhbhg7iG3+bH83dce+cEhc5DcA0JI73Nnk7F7bR/8t1Ld4NyIv46VpbiZkLRi
yPzgu3sDv01B09r9akhnzJwmSYLw72FAxgww21Xx2f7EfP1a9u38r1NcI5yDgfCW
3KdWl/1F15bfd0GjL9dosYk+ibvCQOIc34eBiPqWNusDIas3BNY+Cx7W84RWLJqK
4js+ZN7UUopvNb3r1WTSpE6MTiWUBTdELS9nwMsTWT/4tsWzZUawc3hT9spNJfxV
ZA/zb9kBCn8j8TlqSDZqZEfoC6oV6B/MfSEWsfB9aH+9B0r55OCWu+RKNd+AooMl
OBwWcnAdgfvdrmYrdJHSGVW7gghSxBYZpdgGQ69w+CeFNsL/Oz/1Y/+xAa3jIwSH
saUs2NlMh1NIAcWT7hTCdJ6UwggsLRIqU6m0v0PRZPQLyypBDW/O0AQKc7vHTxBy
1fjDr0s+0Sk0/y8333Be5Uw8EiBdJibQUZbSEXuBP/6IAqGUvi19fp2MDSeRcu67
PFLVa1Nhd+9CkNehKGZNjVP2I9NZKH+dkGtQf4WhCF5Hqg7O4tARlqZXvmkekFZV
bDKi3XTfkgIzsl4JtG/LC43FoYgD4txDd3aobsOQEzkhlKmu6mxQu4AZhAVdQ0qH
BUqLLMThieMVLWcIqubjbf3MAXFv3ztQqfAmV/a/fkGTtBJUo1w/jE8wXiTLK5m2
jc8tBP0IdTVAutRmp2mRra4MHOfil3ofY9qaTCEejiacF7KK1UsYrKN1QtyKFLtL
MiTHnaDoC6c//YkTyyrE4rH9zLLrvttGye331m+Ki7T7bUOrLvdijToMlsPf/cGY
bPDSJNGoK5+g22/OjZf+BLmmTrPTagLHkzWw27Sc7hh+/IzhJLqrd5z3npNEit0g
jWIzFT0dJbQGdAbUxuWSxKjdmdYoT7wyy7Cv+OXEuJ+4dhtiTLj2IMsxaF63aTGZ
1bSE1f75sOmmeBEnbG80axGfdxiHlW6YY6tYuNAJmRGAW4TEJpl3WbGu4tP5qG5B
5PMwoONxohRJyHgQUcVny8rEGMs6hcy0IOABXIyaAusee/7FQWPjI53GJiTYI/U6
DDcFU/EzsYKq2i8T09W56aeMvLpIegob4utrNPrd2W/ZBDsa3AxoULXExO4DeZRi
1YbFB+w+lppHDGFG2ntj/bnfJOzynT2fFSewh6aJxF57Set04jr/iTBzQuNlxpNK
i3orJ79dPQupi/IcF4Myo/OU04cj/gUx+ntSeqvdpdSUWRSQ/yEWGNoYFup2/mPo
yha0G1omSfIR8bsV0SRdNuf/afAlnC/KWIPeJmeWzz1j0ysEqipiCm2QESG/aFxL
XLIt2R6IntWH6GQiY001xTamCDhUFiPn6DFfnrJhjOh8E9RJm0JajQurFeYbqLtx
oZ1oT3B+ZDUgWkeQE+HLUgv9dLHrXeQwrBDoc00or4eYVYwZfb7feWIbWQxuwIY9
nPWrO6AFVxwRDrDmmfrpjOfl4lj1F54lgP7ryYCc03zYzNSe4fn6vDjUnYkzIOUs
HiyQw2CNu45Ix0jmg4jqf0WP1vNuyzq0MzqkZOkWZZvOM1CcXAUq+We8Pcit3tKL
cT3JQfwoWa8cFyPnLcKoml7rGfhTYMdgS+KE2MzRpOfQuUu7gV4GksMo/jDdRHib
V7LqDl+40QiM6JiY7IM6U6t8c99YiTqsdBNuGl0u+7diMjhny/EOkhHpyd/XHcaq
EQpLTjdKM9w5FWnDP7bzJyjRVtMqUWwhtcFIIWn6jYLD1O0lKtU+pVv2rKsX8f9A
n1/2K1lHXZBM568xP4QoBr+UWb4RZNa9WdfCNljKSmkRzMEFbM6D3ccSS5GNSFs6
k73Swp7EDYXeIM23foH2maRYVno6SliCIV8oyjzJrZVrKBs1fIq+nkzOUy2vbHLM
7f2mVCRlPpy32mybX+vPxiMP9sl1yza8nURUYEExPWTuuiyVaJUdr+KnTpaXPufJ
uRmdTidZswjvOPOsPgc+p0PEQEQx1ec3RKn0EVh4g+ue0qIftKinTltOzeOIwLZq
UImqWzZthrbCRzs4wPP4ccbU3wEYnz3RDtzsjYTHp1271Nl6idLKTKimo3w+PpuJ
vYjFs3V+sU0gNdKysqvJCDdtzf/H0y3C4DTZ+i0rkH8KcDwKAG9MtPAMXL7zKMjt
rM8G30Gzl+vBQF9yG3DyCghnmlz2L8+D6Y5gJbuea6IHGdDNkMb4QPw6ngXLzMrz
seeV3vwX4AI4ELKsUmO7ljCzpGmC2yotf8i//b+cEww2ff4ghIL45VG0pQ68z0+J
xrU8vrEJAPqoN/Kz0q4EQf0YzfzF2M/jv82Kxezuky7Vp9KRteRCVU4PjMkGS8PF
ZiOVib7KABQhVr1gD/Gsy1KEqsJmINx5L+ojlm8/04pZYqITEr2Ts/niyIk0oq3C
uKSscXnPZ+sd2u1pF8j+hKGESk12R3SR6hTb7gWYFoEnAIZi6Zfv8Ha+Uf27gRfL
ILXtxiYAaSdtSaH2HA75Ahfq/Qxcp0oQBBx3N0IZRjqQppjvl4lzMqDDhtEnNbgj
DcKbn9NQdA2mHsYtgdIWFXHyb0v1bxvjJlEcVCxXnoZQvQM00rcuXnscnYohj5sN
7Za01Z8Lj/8PFYgUXuLcduMpfX6/3S8LdcBDGM3RXJQ8JGt3J7T4Z6g0PhOtR7v4
Npoth/4iqIFsATiH+AU9HThgs4Rx6zNWoIT8X+Ob+Q2MfjQaaltPLkuHJr7Ypnm7
e+drSIQ9m4CCFg+wkp3gVQ==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GIkMYrmSMCSVkIH1Ung0GxtMCMN5EzmKTaJKYf3xSJOEaAn4E2L6iD3Hb5G3lIA8
w87psYa7/09Wb705WziCsuWqULOa6UE94wE6Opjr++furfuDgz2epYvI74HP7E0p
tO8wx1uryKnswiyTD88/yq+TwiuLNEs6k0qR30GxAl1HUc0LNaFmt3uzgCFKg9zP
BRa5bp1kVThWhamDqLmMMV+XkvTg+zhZFOW8bPVLHzBBGGn9ddACoIELmfeMJ53e
ryD+eke53XApiAmdsiSy7ejp8MDKl0hbLNmxtGYpvxEw+LTefdrtWn7D1M+BkMKn
QInjLaCR3TYu9fKmg5mETQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 21232 )
`pragma protect data_block
LFno5GvdTOjNvdYiHP73FXFwf6aD6BER//Z5DPg7slH8q/TpukLiGPlMCAW6b9eI
2KTqCgHVffytniB+loTG4C/qXhUrRQQTW+cCh876RU8+bcQpltLjaYWN/vR7enfB
WTFBdgoRKlyAne/JIujF5WAls4eLNpnwC1kSceiDw13I3YBb078GOIoAKo7+GFyz
19HOIvOESdW5Wo4o9VGxTnlW8ifZQR8e6GtDSRZqWnom8IDPBzjo527nVufSMna0
2X0Bl4r7kJsTGZJRNXW4G0dVYJFJxyffWPjVliu+KHN9qAf7nY3QAfME+U/j2DuL
dYB71FmzDLimGzG1gkwzbtVmAQyMwXvrbnFxHXY0FMAMUjY5Dn3gxn4jcJImJ5Xz
19gbJvJoribY8P5Ijd9MKKK3gxj18qq4AdhJt6p9/hpN3u67Tu0kipOXeO3mPmcF
H48qsuG5CLJp0vpIxbos3K4nE8yKqrAPVX/UYEIjuLHJEuY/N+vupTtMnW/Rko5i
3GeSmwz7Lse+pIFYUgpVGJOTEA/ot7qCtX9NAsIrHZisI/89315iZMYR5CNLTjca
gIXbHBKTDyHLNh2gP1SOtFeeP590+Uj2rAY30/gIhCVVoyGw6HskTc244B4AItPr
htABr7DY4ib4PSLoP6wyFtKB+Fim8fh6bWxnr03Ji8+KwVsBoOM+vKTU8WxRSuYV
gLzlNB0H9nZT2M66rtnqYl9cjA7xHQEUjs1MxtuOiW86RilpCjGsWaMIYxVBHgq8
rb2nrPKOzpVbtHhepPMUE2P2wD3x9HE70joy7R5Qr34A9Bh9GgjRtOi7Q0eNiA+k
RE/W63EGTnuQZzyQJBBOMpjd/mQvj3ER9xNtVg2Tg9Lv33kJL/IbxVMG6VENMgBC
oJAGzL3fILp/uwZeVYrel0l5sbeTXeQCBvYMadyZyDxaKkpn4qQ0GM0+AfinouLa
um3kTSn5rQFhjXG72VBmk0/q0KFW0I4tw5hwkbCD+bZyLKVuXNAtpfwSsphvtYZi
D9vz5ctEZBYk5nqV2+HJqEKHVwGyLra11UFe8QWD6bp3q21V/jmn8I4Yyg5en3A7
Nzxhhb6HNkq6s8Se3q/KvSLdPvViXh3kVGMZiqrwGXjOfM3vCcbGRxhYbmR6ZQCq
gqAX/Jx9oLLplZFxJkMoWf9gOzTKk/7+qzV8rhRdq+np8Gk7FJJPpOkhXS3bQDdC
R/DuFBrL6dsM6G/+JM/Ubb0zIyIbRf+DNScId+IvNS7VxycoukZxFywU8qCCfOpF
8PqxTf+ci3Xw9XlRThGPgr/iSL99xj++zqadx3Oi1w9H3JW3bt9dNDytntkX119m
z3ph3zAAscsZ0UDD0rLDq9KCAy24o9DnTSS/AYci902SJRsXrLOjfQe2ihOd6XUv
PDQPsjyrr0YxbXr4fvH7tWmYPFCB+WF1ToHCiyvrICT5OFSampQkZclOMMe/4BdW
kKWk5Y5NT2LR8Hi4ooHxV9/AsofVAqDcr2ltnVOXADbomf1Wo7GKQvfcwDLRZe7P
iK/ok24GUKloxTHhioIOKsKPmXdsQwdvw4EMBrdenmtom+60Gc99utuL1vuv+nL/
EelZn08TzFRz9PPD++oclqAJ0XFZpRH1WBYh+97SBYhOibsB3mi7QHBv3PwK/H43
5KHcnvTNU99daejGjpzbBTfprqTynXw8UyOOTLw7YlxgbGlVygG2cKSeJsfjxlo0
zrtZv+56P0mk2lDLjIodHEJRSHP8ztgCEX6n4TKXs120b0iU3ZvHEoWuVf6xOd2B
IGWXsuW13cOdiedmaYwpVindZxaaL/1BAFq4x7qHpmEI8JKB+Xt71/3maI8eoAap
Mat6tCGZdsTsn1Wmp7GW76mTuYdj0xG27DuiWQGtI6I4EeU+6qstvkI7OdFmLzhv
qKHjWjylfB+LnUuGmB8UnWtyFscstn8PU4ziXVSibMsRp3QmBxQ2c87VzUH7pQmg
HljtR/ILLJJ7nQkKBwsMq5LiQU3rUow6OSuXPhUpDw0f4JV1FArwhVaIk3682ySe
xNW/NJsGwUtZw8QWG1g8mbsV6zzksYetK2T29ONHJPxdjGAWXIw+nJIBHj8CFO+Q
45GRQKpi4PeEvzHjMGXMgLv7bM89lkpfm04ac+9j3Ip5gqQj+f3Enb8A6ZR+z4sy
YpY9cImsy+oFEUhfc8HDPgN/TB3rN6h5mLWl5Ek8ytY5M61sz/HF+sA+7Bjz3eK2
TOi4yBApP1wRfAXFlM6Z1Qi4ca55qVu7cBujGt9U2I3Mi4+bSkU1Sp0c1iTMYrzr
BQ8il+CPDB1MHh9ysZiY02SgygL4b/PEXnmMcZk/aWXnYmZDJW+fW9ARIr1tRuTz
QPsdamQ4irJn3LJlB5tulL9+mhUyqPIBWRsB5Flyz5uGngjiLrWve8TfIjKkEoBX
52vvqjk7yu8hOQzmenzbH8QMAPA0LR8f4o6D4Tvo8GAq7151ChcHaGOVaR0GKMk3
p+4qrIsRyJvr9ExbUMjE7L2wpYDPAlU+VxTL39kQDQHSfXg8L6/76apU/tyhTdKg
ADvm8X9Y8f+MoAXQ1M5ck2VlSTO9Ls/mVBxgv5ZUOyeDiyllfbEYzYXujDmxOwZ7
elDgM7GSohR11NXZkQNOvzbJ68k9Du8a7Zkensb/RnRBtXvHphwJwMmCKA3RhAzD
efDOY/dQtAqU41xTsgJh2AepNmROBNmgt8yFjI7sBGyXdBzVnpuONkJhi2813syE
82eyR1DFYZiiKKTVyYzSc3u9QNvsobUz2WebyG6Xe0+d96eSDNOSXm+seI5SMTNs
lSkYXQfcPjQchy2ff5I70IXKAgcO+cYK6nrgSJLX2zpX1eMfqiikjkMcmMI2vLmw
vdZRokZGNeacx8om2++FPOJKbx69+bjfvGyANrBYc/6FTCElGETBAFp7fHzObrUE
akuvVKVbI9z2x0GPpJFEH/L8M3avGp3cbmCfa7NXETXDlUErLskWSbmAHV+J2fMH
6tHrNm2jaMKaV5iobsxuOKByBDtR4dHeVYDwTybnOE3Pjm+VyH8MdTWn8fd9dtC1
Am8nECSo7OjGFHwegCXRl6AZ8uycmIc4FPZQN8lJl9EHfWKh9//1RmjTxveB17+X
NHvdK2eMtHeL9j0TssaSfo8UvWfLx7QDFBEbOv6YsdRMBBRsviB752rwzmadMtKE
tiplOe/SbQbAhbxZIlZdyXW+x7OJgTzpPkKWeeEVvDk0vVMr0GUJZfYKvoOsgiZ8
Hn+/j+mtrc/RGSgP2ZCZr1etno9932WDdSn7K8AIj7F9X7O6awaM3hvzjnUv+66s
luvXx+wH4dFjfMVm6RD9SBwhvH6Av/MuAtMOCrlPWk36XFecPvujLkCDtzovwMHZ
pbEsF7ufe4oOuUXxThH+XxnpxFIr1cpAhJNvZFysnPxN0Maff4AgY0En476jjhzB
bMDN05l/nLa+EfhoAh1yawR6peldLs6/zrR+Q5IrGsgZFV9ix5zB/+Q9lQyS0z05
i3Z9ZqP8DjzprHTQ3sihWDXmBug3XQMJFhctdqSbFyzEOjhf5e/1U90Ui4Agg2mU
KP5tfvJXPmGOnwnKff86K2jR+pmbstpX7A6Svh9xZ92UUbsoYlP+QoiqCwo7h4KP
/gOY6WgFyhKXF0rHFgnq9HvCmNhYsD6PzIU3HwWD//IvaMJay0cTaEGuuI3NSuZ6
pPBE++iMJvmLnF6w8eflaHrcaiSeoaWE2XWmP0eHGKESP8PtxWod0bPiYvAYGHTm
B5JnGyQ2fUl2ZouR4aNyr4x6XnHAxpJZf/tE9AOH3WsdzTCU/mgl147vjakC7uF7
RQFhpMJp0PzSKphm3EjqYfOJBH0jCtIMtgQ5PE2zBgJS73/uni+zLpw4T3ZGrc8L
X0skSqoxpgG86dsQaFmRs44ckcF17v1b1brJ5K/LSo+tCKem1BBoBuR+cVOfv3mu
91KlvmXjhvkWYr4hNGeuT84kCjINvyXAGNutXqpM7Kfx1/p6AaZUW3O+OGsJJX9Z
f+VckzOW89Sv9RX1Spig23blgTtlXYIWkQRvrk+6vppAy92l/otbCuF0k3hbiaVx
6lPsikxWQRig299r+1eozhHFUhoIz4PXNuDhNRcBaEe+nedJyqQOMNw2vE8irvTo
LsQLlbnKej0J3Z7wmP1dJtrBAHtw+isfGN6o04YosQQ4QzIckCkz/JbwokJz4DT/
IH6+A3L5jbMFB32YoT7cgwfeKw+K79zPRU7zdT8dVibpBDgMWCNzFjqHlNP0HVJw
9moHULK9XMXoA8ukkw2y+rrgw/1d0ufdyRRa5wr8fo/bg9/wNyr9U61tOV/xF8QU
eKelsSjmAyB13ZTgax46zIAUF3DP40MVvTstSkUep0qfaEqxOVTFIi2H14PzIbk+
DzwcAoxKahW7vW7VPSwKEjSNvRi93cRQrf8NtzRnh9ACTsJP8hbqXiOleJI6R3/7
ZustDJnqKWcO8Mh3V4lzpcyNCkAPEQlhRgtR1E1MaCarj86C1rnJAdI/o3U9WZPX
0ZjKGVF1jYZH8TNhkdNo6bj065lhqZwEgJy5ccJnVtA//YwHK8s41p1H0wmA2/yJ
1gaJWhXINOiZhETSIwLbxsPCmzp9pags4cpyaYY7ONIxYyBt69Ig4ow7eWDVQIl6
9FzggBdbtuyTPYwMqU6MXy4uM/Jk6uxtWlGPFPw6TBGeSD3gAAY8bGsTFNx2p5Ki
WedobUsZD9gVYYRi3tGDDi0L4K4xF4wt+EIelBQJ4Rk5FwdtNLOh6FX2xunXuiZO
dJbX6BMhKw+z9ZjynDvCUu2uGseOzxaGaJa/zkGZ/1fnvCp0kiVqkYyL1vnqTIlo
rRGycX7COJnI4wH+frp5z8u9jGHHtDF7bE95Xvx9XYHnYHaYgJcmZB/Svlk/8Unn
V6iwQY25z6c9C4CeYr/O15PnotzGMDCIoaWHMXXbXdWFiNuHj1a2aZldgcTfE9Ik
Sfw5HaBlyLl8gK52QokB4JynekE2QgKzDrGd24XpbF5Ruw1Euad0p3tCzA/LmvsH
WJAJsAJR1WUGHGEsGjTKOk+iihhAE8vLnPq+EL+tq5TpqUHxBvVFULW1dIvtPi/0
LOk9AjSwPAlUZbdHD/tc/LMmt4pKsnjHSh+mLQTAP1A25iou0qdrCJpEArHUIcFq
ZBtWrWgC0NErJaoMUjIjTI2SQEoeTL4tSe7mz/ABQvOduW7mVENVHMfzBdR7g8Xs
HKRKEG4MOcBJWDnpfOtb3WeUghG4746qv8wRZOD/ZwS98oq9r/t+ABpu0tYKfK9h
Bg3wL7pnZmjuCDFt07P20QJwqamb1LV/+GD5mvrEoIqnuqQdr0Nvn7t4OWjA5AH+
UXRaEENaNHqE1o0QDRNLQVzDE4CXxp2Kxi9ciPCySz6dat4kJ7+k3tOl0SwMnLGU
+XUAdoctE6R6i35FAT43hOSIW4SJJMd6fw7nwiPW2wS7hDvprw7ixBzqSWxFEpBF
tkj5WpGuabu0CUhFMdaE3afPuT2XOOpqTBm7Nez9KacGTL+4/1WoImPKoNdRvUE3
7UFgpXdSu5TU+le+EDpDOYXO3qKjKKtwtxYwOlpMBSAfMfNrVZl/kAv+g4pPJrgc
vJpBkZGkMVqL30wDin4zBGHZwSbKVzq6f7sSFGrBghH95QMD3B6N/NvCAoVoPnq1
FbPt9U7A1xUtWG1o+LXYjVsNIqBVqp+NXDjd94XRucybDWxfLaTT29//A2Mu+B50
9SQ05iDMwtvUgh563SfvDAIbr6TIENqf3qu9opo0P+wIsEefeWVzFT3E3aEhd+hI
Lr/Ahr1CX6QnhzEW65mGKeQ3p8m18BJOFTAvZpQYyG0xqlXZjTTxoiIea+KWntj5
t8NLk/4ENKMA6sc2hLy46QBMYQXqPDlyJ3ab/A4NzuTgh0a1FrjkUHT8LlghR8zd
iUFLfxiCJCjpjvbVYxxFYqB2yAElVLST6fsL+120e27r28OIyKS8XvvNa0CqCdsE
WOz7F4nZUcFdnhKFukhjNhVBMhcbki2eg8zsHCkY4OL9REQD6VSvlpQcMOqZV1PI
s0ARFK21ry8R9lUspxLQnsnFSEOyJw+HhNXn/FWq+o+rP30XTIsg+0s+nPTPeY5d
WpOptX7zTQJb7+DTIgWkswERhk4ByyNFX1OqKZCCWONTcY1HHF6BJyURCRNyieZ9
k5tLBDjjog1V8cQlXiyB8U4lKjkIIb/CC17DoUgQYmSgnmTa94HyZjy1b1qKsK2v
EBwiNu0ApHY8mtfjdiZdbdsVwOVbjmbcSPu1OF0B4Pt6KW1Q+7Qk8W1OTv6Vp02t
1LmbgqQOpMjDyrVMYFrfN7Tcz5J6sNe93K0lE/yS0IMDupzJqU6kVk/N8IHz6zQM
rt3j8mn0BizjD1duLeVSFWLSNbbrLm3p3PpDdr6HRDwa2I65mkvw8E8NOVmuuYZg
m+FuP707gNMK7qPbJyphp/xMmUJQkM89b2hgcXrf9+M6ZPziFIYO+8VXgd7xSJAm
Mc9npfAe3blwtAHBYhergdnxps5oc2NQqmGA2cewGjES3yGdVa1EDWtg2rdU4BP/
2NaXEn+CVqU6/47MjgRazVfRiprZMBl4JP1rGmZWzdlutKl61CfY7JW3qcKKwpFL
pHDvU5RObBXJCIc7De2OUMgjzPDWE/oUfJMed4cOjitpd9vjjnGV8iibpGTqFkjQ
+/NhRR+64nez3SoA9wFx9lWDbvxA4fX2nU0RSfwqNF8RYllta+1QHP/aFuG0mrP6
DAmQNnirZO0IGD47akNHRLfPFv1g3sMcx8lxk04yIyHH5ZKbphllt8nW2HaTIgEC
9ctkbaqUAAV1KlFtAZopRBl7kXDaXOn2u829k68S1aZtDCELASH4CScVh/V3zY+A
ErhqcEliKqHkKlqfy12N+6EGCdf90ZYy/0rlQLJkZ0IfTlC2XuP0YEb14Xpj4MYq
E8G6PFT1ExINcBVKPvRMUcZJeRRQLtmzPT7UcMABv54gGVCHyNm9kWiJXBDtgWHA
4Y/0+9168NmlwPKsEBYqEkEZGZf2wmtTIxW7gCqeTIj9ZYugbtHLLL2W/yMvEwv5
Q6lKcFyZsppumg6OUzQUomY1KkVyBz7/IQcQyDMasvu3fUmEUFuin4kv3vGZ9DJA
sPlY7hzC/ujFup91PbkysBr7uJNx+Ogo9gAWAPprS2D6R3clY46rcKOkPo5mMoeD
F/YNM9wpwPsIt7ck9Bh6zNb7sFxRyzJa61eHgbowmpdv/iKF/z4/XQarD2A6SAK6
SZPx5y5acMu1I1hBWT5c13Lu37kheQciGWLBNS18akKLEKSyxzxqhLcYiXBZf45d
Kj69VBmdx+PEqEtz5b/8vOx1qjtEE1Ynynghz2VPbDhwvcxHnIrsSYKPG3STMYYX
Y9DsnHuTtKD60ku8w58Pt1IFxpJKirlbDbf0tDrvo+fZmoHe7xBdzvmwP4Ho/caZ
Q7uT47YsC/lpFtD2a3ltEJBZStWnwY4Mh/TXTMd86xd/xw7/UpplfuRcdOV4Y0GU
H7c/bjt4mk+RyozczXGuxpWJW9lg5uebNJLFE/wQ/Hiq/ISn8hunVKq0n8S9hcpx
zmeop6CQCpckKlR16x8kr0GblRwrgXPmYS8U+v2qDql3t38OxNPS1XbWttAiu4OH
BJg55utECAa2X5LpqO86MhY8CtHxp18zYnqaArl1GZgQsbGk3wtTg51jUZSjQ8wP
KSAD8zbO1NrG1kTYRVRYUZf18Jgopto7p2yBd+XE+XD7DmzfpHqHPWNAZYVs4jA/
fL9IK+apHmBvbcHifv2KKILgLMfPWF4GpT39JL8rp5sJrNeGmJOZRDZ+qtLKOY4Y
IJJ7Hvg9UZaBxvGcAJhpuRxA/++i4sg/8zsBDyK4P6HGjjEW5B/y+7lrQ0qIEs8f
I6jOfe65k1MW9ZCo5cUQo5PvYcEUhy/WmaTIt5yZ4Gp+tnwARCwAwvSeDI62KyUD
0/xeskBVu6lj543QKpl9o09BFwbtv5eUTkOuOjVAj3cM235mc1SUVEoZGWhNv5lk
jbMVYTmEHzdEu6151/BDIFlmXswFUpcYQ5x2l9/vstAdkBF+v59PIXUeaaE3GbIR
wKN0r994QqfZ7DdBA8gJs/HDSVvWXQlddXqeeojLSYwSmPVMl/MPfkQYKZo4PQiC
I2jZjDRrytxEuxwaPtvWHgd2WexRYvSBqfP+HPhsytMDv93japQg2TDODwV9Gumv
Z7tzqDFGuAm3JWyxqOrKVZRuo3HU3RzxU+t28/c2qcnBfBdim7smXht7k8A/Gk1g
irM9k8FOzB7WtVcrlwlepeQ9f7gjdC4HgHXb16qd2UEvsqPtQwe7V+jg1AzfO/aM
e5ya6a+P8WCjMenY+h5S30U4L5kD4y4NXTYJjUEk+HCgje/HlxfSMgA1O4zSooFH
DXaaJ7HM7vY0Vv9/K599ZNAZYneoXFXOOCnu2WzeFU7+OMqrcl/pPutGFjfFVEE0
qROvJte17NWEdYDXxW8vgAgWpae18JP7QdlQoOs+FufQnei83ImuVsLW8H4rU2pT
rWHgmUJb8hw5bYy7xqetBCRMBl1ikhZ0An+FUuxoQaaE01xOYPkc0RVJffJ0Vyjx
nHeevbquOBS6NN/kr4g6EaLFhXxC338AZggsaS4Gr/4FIWQy/O2BOWBuxEAUC4cv
fOvEX2WESbF4BFZAasqjw811d4yD9cjfKve8GscoLj+LOQ/ZjWq22S1U7/qKMD9T
Wq9i2D6gk9mu6FmKpmKuiQG4utCvR+lkJcz1sjth7dVFm5Ks/zS7UqbWWgMMeB4Z
ZSWaXHL+7Yjr7ncRohZX6N0TRcN3BhQDLumVuoPLisDBWb9mGkwJdKf4so4regM9
LHTH1HrmN6pYjO5MwlnEz4iiK/WWpabgVcED9ACxlrG31TwqhNa28lE9m0wC0nzc
hRZ6C9ohtG6OW8wOrjl4FnxnvEgrQ5wPhBNlOFWi9heI8Mb1wUPTgCFYFLEWLmpP
Uq91AWT3MaD6A3gFwg4UxMIuyKhbOyZ81FZZTP4QiWIrg+q9y21hgROqpCJl9/eU
xwHZRfjDx27JQxeNQnwpYgzcPc4ywYHZK+p0QtXcGFuMqyOU6iFSBipDUheTzYlm
wKs+mqGl9CU448LWRNOVn6HbrGEoZnZpVk3Tb/UYDJ2O3/QLksRiCp6qh3T9LVhL
9Elkaml2gqTL+9x5ERvaJWhOf/b4MuHLmhKZgbgfEAbZX1oYI0dh2eaTVVeawAwl
5+13mqH1lb2u17fM/UGTTq7M3D6gkKD7AMuQn/rgNkCmVH+XBq7vJhZaB/KYoqqk
xK3sLL06oWAMGCn/x/0yplqD0Xd8/RJvFRV3sIawwro+ZQpOR2Pukg7+AXswY5QI
GFN/z5sUgC9lT1lo3aOLuCH/XX3BmNGqpeHkWESbO2+fU0aWl06+dGOoIAMn79VA
LsowGo9day15YP/xkqhxzwkj+Vxd1X8Y7E4E2yw7f9ccsHoKo5xlgyNAbvaPKSxd
hvI8AytvqZvtOiue0ff3vOQC9X+2tQi1o9mP60HJ87eqJeICL/EL5OX5Zn5LF/W8
nBQOGkrkgutgfi96cuDDONxzEj35VSkB0lrYAf19xKw1i/DbzT9YIxhQ4Vq39mfL
atL02On9RPmbBUwzcIKsAhLh077KG6xzz814PK1+it7KJeW0HLmnFr5rtjc4v1X8
Bjik5JnJ/fPxFn2E18xh5k6qfo8Rh8LaACIp2m+DiBXAB+9IJM3/ft1O8fQYLV1m
E4lCjkA5+qGlmlce2sGs0u+3QIzqHLMvyFrs1zFuY3gQPte6TYN2m2LFhRWPhTtN
MCUrAfn/LThKVH9c2BuF2cILtNnGzDr7o0dWIvsSl1klzfpdIiIwwSSAGyxvDD3G
cbhuM0dn0BvP+gB2ZROXyjTuXVB59LRW5CJrywY1KWzBNujrxakqMKVZG/Bv6+2K
ZcTMUzYq14v0EuOfUkLBONK2djkiYm3Ri+osIanqhquUiQhLUCJ8XKBRXaDNwTaS
/5t/Yiqf7Aagc+6xTmrbjWbZskshMdpPmSbBOvgVD0clpD3bMrP7wBfbVzqaiaPL
P2LphKnT+1vJEMKVCyT9UC0qIyiM4fAOMsqtbwL2+GmK6Dy7luutqYM4HhVHm4OZ
bOfh+uSdX9vN1Y53gXhTVBH1+TTYZdAKI26rAJgq/QWGXEwMDbW0cuR34c8cAHBg
2JieDGdK0Mi73KZ1wwEUwRF6FV9qpX6wvLMU/7Bh1wVh/jMuS1MJniFhOfHmjBdw
lUa9ThSwaidjZ0i8tpWErbXBRcRmS+ve/2H4V2eDSK79B/j0yfnVrCOuXKVMM4gc
ifFDiW3yhoNcOJvgTuRyZa8wwjI5PPWTCnmyyE7He4J+wrJgOjM/37n9Hscg1uaL
au3sZ4l7gTcX5EoZRGxIUcB2bI47eBsZpZo3AKxht+mUCPhu288KNDCtQmdhc8Xi
uC58NFY0BvXTJtyH+xBWqLX88fgVZfO3xxS8l+BAqc6aORA7MEquVSgcuqLe1rDB
KMdexTCHWNQHyBG2EYK/KTUHlEq6w9pdOnDlKUQB++oYBVJv6AtZqdaUzD4xwIpx
P3ZY+eNBY2Upm3K3Ne++cQA5Yt12YASEBcyZwwUdsilYL2dKvhx5/7DbUojn+vah
V9b7woGiuawR2T2j5cvismJiqnz3DciwjcDSXJQ8DBKAXRJ011iRXImj1dBLh6Yx
SW29MyANecYhsRi53jVycREcdZZOs/Tk5j6MXFkN9LVQXN/QqQdYyU9d6RXn/khS
M3qUFSBiEtnHw9et7rtRGYaVRGqox7Dz/BrCRmyUJRpi78uwgbuwoCTdgu4F17XL
dt2vGi/817IrEiqyWHYLB1qTGFP0yJclic8WcahFGTecg7SF+5kbvBn7u+P6EJOf
REqmYWuwvxkubnSdULuKMg20SVPXsdkwNGqEH1Cnvj75k7t2+44ve9HkJ+RGvnHk
wGbYyzodfDX1K70ejxwMJo/X8UiEOuNJdYqBHKJqL/ckWmS/60kQ4uG2yN1efDZA
P3MuZyWdfKFOpJ8jXiiEwklZbf9jqNxvLhRIeK0Q62VEhnlDq4+zqlWoBjPkz1VN
dJY+gqUufe+0bRdAG2GonVyfSNrrfGwwL4AUN1npdvtP9fGFnTVt7xTposBy+MIN
R0VeZSXS2CWwbPf2wagHAhNtLIPOuBaDcbuhWPQXri/3VIFCkz1rXeLES5xU5jpO
zVecN6KjQeQOe/kZB72kwoDE31zo01pXYmSiFkyjs/MLZouIRVM/TdnmagEsS+fS
86/GD4m4XQWjjWn7ZjC/Z6yKEim6AHK6TAq7ZMbyHwC0vyLkWQyhCvwAmcQm9RLY
LdWRhEy32ES3+WBQc34cVUjbYxhqvU0/WmkObjepl+VFaM4e2rgWrpuEXlDwMObN
z0LipyiPb0rXV5DGZDfpZaLcZBmnE4uxJBwCS+JBkjCaSex38rQkDQiWcPpI1x1A
142O9l21KdSwtrdquzTErpwN7Q7BDuxIZ6fScMomkrh4x9+/WzGYRkkJr9TLdeEu
jq1JGCSxiNKvLVQFJz5o6+dPF/tQ+uP6wk1qIlrc2VuDOZRQqICtgh7QqzM9tDmI
Z1hgyAtp3IS6wzc89nC0G5QJiK48zGy8vMgg8mZp/CEzf+r41cQj1CXi3F7AXRly
Sy5fl+OLgAhJn+MD5PUeihzDlqQEBMHsb2m2KYq44346KmVRVzOPaFUmR5zrcLPr
9oXtyW2yjZCHgTVRRNB1QV3MLApl/VbV4gc8BBrC/ZgmMTynx9ZcM6CPV/r2Xtqj
qFUq92mLoQ/FY9a11LPDX6i8Y3Dsqppk/kuU+O1E1Ja62d6ghiZnfXmB92OBjwOU
GdY0lIfFmYJ72BfP7/heICfuhkGCnpBBdjwOukB3pM1Z0HgQkeI3NfEAqgS/Llaq
UPJaitEi67M01suHKPK6QphJePpgZnqtLURrRMf1FntPsLEGZPMrV8YslrtPDu1p
6BS5N3jw2fFIx1dqa5AX40ZYUtTKDqYKKVYhdBKZikehnkMagcPEFOL6woZh/ZqS
5qzXsFdC97qg0Dbkl6hnqiJVknkHIdx068E1H+nmVUVm60r+IKRRVe+Zt0YgcTAs
jl9ZWltSRf4z7hh4XIDDjGNhM44k+hSv16F+PpO/t6khomTQl+jLNXV3TEznqqLU
UJ/kHrnpZzXCep79NW8C9ZisOVdAHKdLmxVKTSqySUpgLGeRaPUKdu/nkL4Vf4Mx
mt78o38Xl7et0dPnBMtNStJwhBhlGqN9lM3e1IFWgBp+hv62FTjIN5/olQSU/GGz
kXIpvZ5i7JXW0OBYm9SfH08jzY7O2FTEqxapwvzP/ELv82MRY1Vha7cgEYCRrbUX
mR7ZeJrmwh7uLB8cu4FqpgXPqXjLzVlIdYD8O0N7dq+WZWaxnh2HItVmFh5mUvFs
5hj29Yhb+qr7Kw5FD3B/oHWZ8VVezR5i3ctKj+1B/VCg5svyuma0NlXV897TjaBm
DN8bcnwKo3zFOGi+fRYkiz/oouFKV0irid7K0Owm+yCE0xQzMfUeTYs69v3ffOMf
TLWhh7enTrMa6qmM9jLJRXUPOVwRM658JuMHRGaKXkveLIYPWWRMZEiUP+Wc8C71
zE2+kAlOFV06cfFei+HGhNrcIVz6vtfyaRo2T7izZMNbqUrALAJfCxSvTgT/Jwz8
S1L2asFO5HwQoz1cqPN7LkfvWYN+UyUroAtvWHd/oXaQUO7hPc+mxxcBVTcZNFeE
gfPvnCXEuRe52TQhlgGs6a6e+n6LGY2TQGD51kn08AOZxoV/pp+XaausER5dgpqn
iZYDP6mXzZbnJlYa01D5zsWB9sFj2Lwf2yvnZ863umR/lgsEIqgry7cVPODq4n+V
u+QWUhpM75ebP5UVGpJpA/vDqDWdD1/9vw/P9Sa6AXklfg8UlPRCA1dlSpkHQFwa
KX2y7EqAMNrIk07B3bg7ILgYaiPFBmyZsrhtX0ClXKio7GRc0rntu+Z/QtouDsth
5qo7JJW/AX0Yow8VW13j7ps9fr58pFCDyt7oc8fGrQG5kwjHfgl8KkLrZadU8OCe
uuHTP81hfzjc6mihOzT1/3yV0TaIlBuN3ClZ7Ejx9cYHuF7l0CE4oRr/MN+BE8CE
t9FWbahmW+SGdUSFNrFGqiazXaRy2Dq3ssq0PVWIK8xFR47lo7eWZg7DXdKxyQnP
sssuBgxAN9ipjPchIlkn+rA4r/K2tPkE8nyxtrlAp3ifTnhnMFe8/eYB8v+HOYGL
WuZyTlpDiAnQwgxID6JNNyflkNYlKyBy4OEyqG18fQrmzbs5VRfmHjr11hHQs5sr
Za6hqM4PHQe7FzbIQnCaUD9SRe469rogjOFuDvOMVpSGgAHLQVzj1WAl94uk7I3D
R2Lv014GyIhNMengl6b8/SycmGZTujdQW1mgiy76UHI2kDtBKz7L5nN/Rs1w9Had
ytwXlyMwTke+ZG8Gp4D9zQwjMIUNuH0QnPy5/C95CWuA/PCq++3rUlxuqX/56XfH
GCgnDvzPWrc3uQJeGL14OoOZMJE4mb1iETj9xXs00gm00zWF2mNuZK4u+HCjzrgz
Imk9SlLce0ldE64Aj0pssKETA615RV//8p3u5VusPWp+qmuq6ITL+L91YUkKm4k+
l5cu2XujGzVJrXxy+W0NglEbfB5SeBqq1gkhgwI3Dj3et/7GK7NVi3su1MTRVzH2
gOTi2wfzco4uX43rMeVAWAto7uGOxFymrLoSpRtvfcxqpLwSnRNtNU+Bs9dnsV2p
kPcTHnepj19wMOQU4qXtoBStiv048JYFwQZDFu81eQGojggBdLnoPG3H2JiwTMzA
OZwFuq0o+srmn2aB71dCG2zXHdo7LVfdje6UPmpyXwVBi4V61ZQAez9ZEGB8Ms3a
fAKC7cq6GbPsMKBAkZYdF+h5M8PAt4pHXVERoYJt1grav88YZcRQxgCTV4+7zpp4
f+Iki/QklqCvCp7wp+sBuOs1wd6AVr4FfF/UqKAC89gAhU9/G44pBtfCzXIQcE7g
xCAdlYHPR0RxZiiJfo0mP/2urlP4fJfXO8eWHX4k3GTIJAfcH8hjTljjXdXv8ffG
pf+JK/0tmHWn58g+R7NPT/3x4t35ylXpm9cJj3zO95cjcgs6tvpfSwHv0yjRVA+y
1NvZtXgFZr8VZThuDB6YDB4dGx0DM0AR1BK3bKBygu1sdfSrqbBAfmDJuKKBFkks
gP9h9nEhFbogcNceJMtnUiTYUIpF0irordEhwAuN9NzcsRPswXCSwhp8Ps4+2JJo
OkYWSxTBTeMtLL8b7/qNHLLiLRFa1Kjd/qYiaVxya4tyYDywPE+4QBneUnJRkK6E
JZcfMfZjwxCVZmSEaPDRTv+rVVH46qIlteLs8+1Qhy5Ph+fF/Roskr2Uzl03IcwY
vgjl+91y83xFwZdQFYjq3pl7AdOV5DV+FwoSG9BF5gaa1VMPohsq1zZnz67a854o
7q/TbEbvTJh1B/z59mjAHz9UIYOv0KAx6Hf2mT4oC6ivmVur4dvFx9h4tEj4PBvM
mAIdtlQiRGdm0JN1GJjcJ5+k0D+FcVlCfUnscHFvCcTxXbRdiKaZHZQSq4KYReXy
ad9aF/4UyszBzJRh8HSRLX6L/3PPogiF7QSdOerVTnWtJGekU4VQujmfGPvrwpG6
Ukyvai93Ao8naqkqv2QSbMxPIcmgMPsi8sjb85k+GH0Iw/9ND8UvfaSq6TtXzDlh
VS6UOJgWSttR7gTROq16lhXUeU6XhNF3FY9Yhbcv5fwl6rZ9+71VLDSzbFNYY0A9
gj8Zef/soHbN9nbTspg3inFjS5qUsdy91OgIq2/nYjnYrqrkQch3GYe672as1kBb
FA2fQ5WKd4bmmB76S1CAxJlNGsqTXSU4in216AHncLE4Wnq4uDr8/XWNYkMr3eud
Vs1gdaBCRinHzgjFtCVd0nc0GRj5QFR4QXtsRDfd0j0o/jIexrKRzI0IbL2tXKKy
Wvr9PEzMuXjzw2XuekJAmhbffjrzsBJeNuB4KpHlCnBvgyktzHezwX8OdsaDv1VA
9UoDWStiAg5yiFgUZumRAYM0hq+IGG7M45MP6ma0DadVOl+p1UtxgvShY2qUXLvX
nC1y6kxZuctdN+givMveN4MOiVPZhl+Iqf6MRKm/BVHP9Z40GVaKu55moRJ03/B/
Y23z/khvJsusxDlr3r4i3EjPaLbBe8II30HufeTapzFCsiL3UpxLeJsN/w+449Iy
9K1RbWgjjJ4be30Vt92oCKPh+XUK7sp3fKauHfGTmC493Y1B3CL7kiW0WrPKGseE
8BrtCu3+8gTAizKx8nFYQL1uVcpqUcD1qNHMtIquQELCKAwBMX5K3zbB2HW1i9ud
7WyK+Gls8EwmYFc00SKHpMTqC1C3H4dG6a2JNkLjgdn+sLXTYI3jJZwEVwXd3IMl
EHfK8TpOl8+HMmw2egTWW6qgWr9lpsELI6F2+FPNytqgfrwXljGe1pgxrs/teBjR
ENhCIX2rzhYWqXPhugRafAawMP7mfePT8jUh4QAkRTN1VaSeMArJBicViBSpkQUu
NWPghBmtf/bTJEm85fBA9tpP7/XMqA/mjv331MM7VicwRa3JoNgibA7H1QmtMj2V
XhIdR7C19MO7aoKGIFTXxe1YB6xzo9YWU5W2i/MYcaU9KIofLoDpcNUBIHT0Xzvq
0435n2OkRZrSr3s9sMXH3S5DmETmQ0xxHN4dXHI5JDgVMj/hlFNNEBy+xyOSN6+d
b5RMnf2p7Ck0siBqm1PH47d8tIEBS8yrSEAh2sdpxy82eKuwrDoNxXr9eoU4ZA2M
HM+0qldcwZgWRCAUw+uL6zMP9dFXcUAMS7d0HOUFJ23UR+sJ0MFCxjfb+1tJb2KH
fMiB/u+seWp1txXY2oFFnxxkyxJsDqrJwoJb5eGgSCQxRj7PNhd+1P4KpJPkuBCu
D6S4Ir+hTAZAXZKrUt9yXorBzfkJDa4Za3DVdkN0oJl2RbIq24jwMswAVNjFy7K4
OQf7fe7OGm9StBXph6N09AUH7MaG7fBb0nX8NMdTJ6+11WAH4jILk3NAj/CG0GPK
Vl/n2tasZcwvq2Y1MdtT8u4h2Z0wx52eS3o64zGq39yjFZJHikttER0Y47vjl18H
tXc39bF8posgk7slOY2k10NsaFElKE2Qy/4C1cvh8wt48yiZ9F+zihV3hd8rYx5S
0rEXV8TzEULi88RpEx2lPOt4wCAnnNfsu5+fsL7au6XbZ7KJ8CKGVwuSoht93Ef8
PRrQYImFmbeKOoqRqZ8j9EQtAV0JQGZ+9CiD3UnXGOs+VXv1xbkdOAmjS7EKBDdb
WDvu84yCBg/dOGRrqiKDtGfCANjcqxAaQNOqsPdBw6iKQWze7cISRe4a4NZ12xUp
F9fhVftiwV2pfD4gz6th9/FushuKY3KIQOap8miSXGErpwzz1llf4t+sSYlrAHLu
DJ4SH3AtXLQohOxlC0jRWvSEYy/P+Q2FxdBGidzPJoRNV7QQHEG5xmK2TjemTQpJ
3woIDuLtuMK2nRumw2Mj0+TXEjS3p6Ac9UTH0CjUIoPOO4Udh+t7H5APzJsQ8TPT
3mZyFamG9/kFCIK4zZqjSEB0tRf1+oWh+LGD+O1x6O3yL6t54GLHLQBs9SSe4Bn0
jTIZmlabR/UzrUlunbakR/BZIZEAFQ+hRrj2aXRrR30CkPZHks5Kjk/EuTOgDm57
TGDdpOmsWvWc+SMtSwA9RgDRsSM/FFdSd1wAffbXFdW8D2PYeths3SqNrL8x0xBT
r1JemdCT+X6jeIirqLRlOqYsDOPMsyMWlGF62OOuDABhDMHbcwm1Qj6eg5n3quDh
GjINWdl5U2aMOWEhV/YvAQwWRFft008q8q/mPmHMHdPRTessGsRsxDRtgODZvtpV
DTpnwxUDx0kn2dCnAkEd+qEV3gqLKtZxSBb2M07VRtzpd3yGNhbWKDElj9RGebOk
zZ8mabd5KHP4FGBf8VbHzLCR0/37Ys6hpj736LTrAaHYxT31IM4Z/mBIkQSWp+6m
YnAYYbCR9UbJM8sFe+wJSrpjIuA3900FAAXuvv/BlE/YjrdnoUX9W/AMZKTZBvwk
QyuunkZYf7VWWIPhvEstZLtO2xvyDGcz46vm1WDFp7jx4xKvsLpkYqKRxRoeIZEj
Ltm5/XUE9w2ehFZ9cCZ4NnuqFG0bIQ4rgDSUABrskBJVibZ+4YhuULYnu/HZjuzZ
2iQO9A6nocQHwyW/2wcjKBucel9t53uxh8uUUYudYONX/cV3dGwuPJoritHEKteU
kRL0rMWjIsbXYKDcL0AnQvSoRJ661nkzYBUU+TqopKOmWdI6svz9TsEoIpCvYk9k
/8UG/O40Jkx6DP8vKG8Yyo6E5076UuSajKTVPuoe7EEPY5H6TvrwWJHHlGa7QDAL
WyCCGQkKQqc9Q7c7r56WX/NvG+/vBxSj6ixxxeMEso5CYBmP7hUD6HwGOySpQVqC
u4PZUzH/jB1ho548CSVz5QRBDOovDVWVV3AXREwcXuCma3e3w6Ra1Oioc5cNZZc6
OeSVXTVa9FZZvOnE+YJ3DSHckYnM4uuq/llCe+kHzQOXWaIEuGE+yxY/VDk3Tx2Y
CDH9irnlOq1tSSMTvvDLqw5wY58Je/cu4Ytcv4ZD/AvEdMlTA+FVM1nx0jtGVKWD
7ttpgs3ZdJa67Gqde5ks0dzZKUoYBxkq5gfnVC9Jxrhfh0tQDkwnAFnk/KybUo1l
Qjm39MjQr8SM859aJwKfOyYrDIaCEE6+Ac17cc47+7yRs9kfYywFi7MOToQ3E2vD
G9kemjruMbdisl2YKQN+tFodoompbeAsrtHNv8cK7N00Zfe8acz/BLe63Bojgf1u
X18HEgbs7tyOcFYzFB7N1hAif2yADWQ200gucFKZgvrEiRdAwyg5B4oB3U3DmI1g
1FOWoWCmrW/M0cb6/RXlN1mvPvd2W5Z+lZJ3ll1h3/0PEt7osDAIAfPbr3SREPun
ZhptggogCPBhZqAWYR5U89NmvjLoLwy8fRKnIRVCRxsx6+G5glY2wKTjIYJuZqFc
255OfTwADP2/ctWUpSa1CvTjR+ysXUIIoOAnyrOWSelm1IWgCCFwl0gLtyzGQeDo
92+nYmAccuOxIDfYUx4uW2M4//KbcI25bLdwYDJI9q2y3yBwudkSLK6WXZsO+4HF
G8DyB67+Bn06dovQm4PpmNiwV15u2W/QlrULZwXFZ5oEv5c7dpCneqnRABxsw1E/
V/+WLcsaxyJ5qCSC8x8wSts5VqWAKcYExwj1wGlmyQCqG4tLIPrnLPPymY4lT6TH
vQrFL5y2IwdI20XMmhjFnNbfD2sgPjPpEi5dR03v4VOZJ0RdXhZ7YGSt4P2vABB7
cnmqtXGTB2AhRlw3QIGdcnDP74CLRiCrc4AVMlsw9RAbrMkdolOtyDNx1+JVmiEW
BVHtmE5Im/RtOZ/utGTJnNWYc0SSDGepvmBmbS38LKl70x1RXhVlggXfiAE4lS7w
ddbU/Uv3hT+UWucM0KbvGLyphT5IL9pjLPSK/W0EKWAXgucSHthVsTAhXDwltQj+
d1gHaXu2Uu/Mm3yiNwkucoGU1udosJQcmryf5WVpcgDnug409jImXG6KaaMvknbB
pICElZquIIA4jgG/3vvcuLX55+TcBAS2+Wk9wK72a1H74ZcEtPP6YB4BDwH/0FYn
JNGVyKkRt2iFqzTKCxMUR6laxEdo2FxWN7rNOIVnffjby07Dt8KmU+OO9EOSo+h0
oBsmZzvAnIbWSgmMr4KJvtFnofrtZilxvB2C9/WQWGXYltvQL1VewQfU6l4Ha6gJ
SU1NBk+VRiMMWT+cGo69uLkimvb/kkUtHkP3jo/hdGj3WLGICPtJwseBDNZL8Crz
3ZXnxlPfDAMot5OstfZZq2u9ADC6HmQmE8rLSdoVoqIkdMcoHIglnPAPp24PXPio
pcscSVoVw8u3TsTz+RxLWMn/jC6KUn+26nF9ZxYJaeIBzRQwekDCB0gRGv0ZXUl8
crmXFoIYynILyikgShDDtSa6+xdStKV/gSSlKxKhh2+KdwfWT288aQi69ruWGrm7
i57rojZPoRrQqYH1/IJgYO+dnXrj8HOd+x+3NBoOm6dRvf8MJMj/Kvd7JjiW50Rk
wVZ418i1rwU29msCtnSDuK1IJjmMqBZka6oFxVrE82HglBPuGdHGB0sXowFlfhKf
umbqHo79U9ZjgrP2Ts4Szk0NuUyW3vf3AeZLYamezqSzP6RUyXeOfs0siMrIbvou
iuVE5zQnXfF/J6cmiUzXaNNAZ+bBfqAtsi+OUiBvAGQ6qe4LHtZSnhcVnmkEhroV
Mqv3gxoauIwc+a3O/UMDdhbdqoH/KxNoZbM2hRomS+NK4dZItQItJdu7Nm97r2jv
iO5mDBKsWafKv4tTQVopsUygKrzSgX2Iqyt/6OidzGPn5dimYE30QgXg1AuvTgAk
qcb0+ikAuHhLJBD/qTpHWTabNvHq4xPUvw3Jig9DFJ3H4ZfETCUb3rb7UKA7LoEz
90zSKeIhP9qQI3IBjsZh0AyAyt6N1v22HfSH82uer/fQN7krT9EDlI+/UCqQrKBK
EntQA77hJgFdFgoWWUK0LUu250/03KWcwhIuyJoaNbxe0h6StUOQcRTPolxnj2Km
NJH6cKtrx0SmCoV4qH2NjoVk3uRSGlypICXRmuCHpkOxcEXahu7OeMrPF4OYzwQ9
jzY4eqD+i6S/us70eHbPZtGJpmvIAkBrKRt5vEyT+4xw3X2ODofkHu+8uCVyaFpJ
yI+lp69wvflxf6w33Rwa4ic16dwBZvSvhzZmuGqEabpHZMV1OSKJJ9TB2m3TVnGz
iPPk6Sj+LOousieVESp3P6Gr4qgvs0OA3cBDcEj7dM7/h6mqpD6V7DrLNuIsyoIr
FDwcSm/53jvQUeRFJu9AIS4OPhS34TJTgXLeCF9gwRJcxzYclK4nrgt2eFdGwxjB
m6epQp3HpwZy6mxdtPSfRp7ZiYWbKnodLD9ez1zvqVpGC3pOCQhBiWNpVag3BrZn
fhJBTeJZQzrH55j1jNKY13h5hamv5TMf4QG+Umvuv+iT6s97+qgB+7Uo0tT2Qyo6
71CEBl4cNWUrej7JeAeHwLYNmeJZ6tKy6KSBlp+itsdbu/3QKJXDRjLOQEDrGj8S
HDt+fMGCK9G5WqprokftZn4lr3sH6BiKNU5DiJSYlJR/fyJZ3M+Hj+qIlczHjfUq
AGvvhTVWaPJeWfwlf9KfR1TTGigedRP8ombHgXehe9OPvVPxgQTeu9LaTJLZ1bqO
ATcSRR+rKnzRL7EUgjdug/nmkbUbKAcKlB8a0PzHZZ/E0+E/E5cfdhI05K6aidWg
TOkpQK8fy4COpQujTaWMKs/FcXALZiP0drsR46+odCMcejxaTGL2sRzP9xtvxehy
JhuE/1O1UhmHFfDw+TGz7sePUL95oVEgDs/04ble+WBXqmT6MewqKekYPf7wfgRj
7eASVku8oNq6AUU+/je50EqxQkDEOlnlqBocppz1uIQ0tbS+K9arNmDa3hqpGRJV
ZrT9FjufSEbDtowAh+O60PQTqNAVyouxi6ell9vtGy5qKeICzMTIibM5zkH/ORck
zZ3TamisejZPs6anPw1VEGWzNNPNhJglsFlxtZqqUhVXkfzlJ34LgTmY1xEBO4eT
Iqf666+grcrwviisA3c9RzDYXI1l6nA/tjA9Z1b2LdhtLdjnD/rnfdeyl5wxjUhw
ogw7dpckAhaF5QE/pY7wAzzlYf1+4zm8cBWthFHJffDXQusamk06gRklm7sCW7PX
72oah/QkfhQwaAXQ4uffnoN0h+nQ1O1DZKEbmQxdstedCOkXM2zvn4CMjqmf0a66
lgubVQN/2yFgiQl3mUTRk+yDPl1Z8zeNtKEoQWRM/Tl/hqu5dxOHhqa4hQrqwzPt
ruLHTYZ8uUwz7ewAgW2X3HuEJDdpibM0SaydakPIE+BOyla60KFk4wNBBmxA9wkj
gxbjPL6n1dVsyEQQa/81AirvUXOFcqoB9sW7PId0+OfgSosBt8C/HBuAoRH0B9Tu
WdONr3hsxXGIdZN8pgvGQxPJBFTzBs1pNZUS+gPxAaFuEmQK3e3TvLfSEJn05o5N
760DtXhxdYuzXw3WiTFblxq55HTSGYel3vmPjoRiuPyXj2i4i8F/GO+3PMeaoHlF
F+SHbwBWy3hVs8nSnRW1CDuRXRJ9VdfYQ7QHPrIYE3ta90Ifs+5NAUqUf5XV2mKQ
va4no6TFEbcV0+DcsSLST7v3RLTdf3ykqQ6r6VgnjiYsUu5ncfVhJjpmDNhCzM9K
EJrombKP2fhPIQuTCNJGtAUPkvmJIEzRhQpJQVrt8dUZU5rTQZAhg5JxZnjLN/8W
rOVKheZX/Wh2xh9oN1McmuSYKmpXyPR5b38kc8toLKJdS8CUFIlUKOp2rIxeWLLI
rj7lCHaZhHERFltU1baxAnrjscvoPN7YxGVuhMcxRpKG334mTmFfc9KCipJ8L5RW
42BCvs0ZdVOI6Ghxj5ZRgz8+8Zlz+uLkOMl6xH+RpBIgE8PSfiBdRxrKKxUlyA/u
2ux2caNqqaduBYlZDGR7PKtkMSoWt9Vf5Sb4PmB1rKJhkZIIOATjMO2icwxDYoaO
23kIOXJJhvhzcpR+96SvWvlYN82p57ajeHfvOz5cZiKNbgNkpnSCReZemCcsbkca
ZgVMZyj/xNk6b+lI3ibMNQaPzNt+ouKQRiTNik2z/Ok9rmgX9G6MFgCYEyrBiWOs
YY9/3lZcm0PZwoqlAYne1WNQ/IP+8JYp6cu93oZVQXXXcaK0BbuTClxEwzIOcIdn
tvAgUSK4Wr70BT26IpNAl5kh0GaME1DjRU3c/857Dljz4PlE6t3mwujp+ma40gYi
fkfButQAUltUu+HbyxILwHhnIbXyPP9M0Ay1T3yGjJZUCrm+rXx7C4sN8hs5wWsO
LSjkm3hR/G+m1hB4KYAmPS3tbCgBhBf5FPwllQU8vKIdZI4OfIDDbp1A0nMKtyTb
wxGSfLkLvhcI3dKYz3WpBGfUfs91Vi65TNQw+7H+LHnHFe1tiuO+0ZybGPnYd/q3
Y1A79czyP4Gpb6PkOwCztTsR0+iz+HFSD1mxVELvG9/O+eCCvkhBtBhFbaf7PA6D
+43QOIIf1I9NI0cd6OQ5C/mWbZJ9+Lw3ThT0djZIuwBs/6qoiTi0sfS8we7tS9zw
dP8A1if6fqifMB/iRnfop2cubSbUNMW0EW4/qrcc3jlkvsEeg+Q7uM+jN8cHruVO
2qKyq6qMVWmRVzDfCaLElRL+8J9Bg+dGOk27AQuib2y33ZFIcjCfuEIn0SSFhJLu
6pSh60c+jsyrNC0k/pJObfSHb2efS1sOJrr5tc77uVGNFmRqM++nYAjCGetQ7BuF
B9m/tFPvY//kwipYh0rm/XN9PuKldzP/T1+9DwmbUs9y5IDhzkdHCMRnhbV7gQwC
czauB5ymGPBUEfES4XffH8otgIzKnYgVlvEo6m6zx37vI4baWQG/6VzAmtZpEfcG
TYIY7cPYeojeDHKE0FbNuU3UgxGf274WgaoED0RW3lwGRByQQnFRMcGR2dYCht/B
Ti6aJCiSx1ANQ59niR6LYQZUkSeTtp6jjKViWgIA2JPdmpeTIBh3rplF9eggkimB
p6CYhp3+8Z7RMesMzWPVtp8o7/SAWFoaK3aprHQBgmfXH9AnpNBZIbqeKWV9iy05
zYSRDe2VASRcCsq25Kf8Nx/t/8FpUkk4U93rb5oWuI8xZ5bMrhnzyLmM2+ZQjdv3
esMU28CazZt8Amv/gNlTsRs4pHKLZFiwEpcZsqf5bvQoAu0Ykh3F2s2TrX55QskB
BAczSaclP6Y9++vgmnaVWt3P5FAnEo3AXc+P7lGerZT87h+XgjEw9fEBBKDC7tSZ
y3qooSZnUzgUTeUZVkyH1c5oknB4LuCQNiMD2ExQLQULNasU3XsD5tcYqUHxlkUW
HcgBdyXWaJDdDWVI9VGiL5sXIDCAA18/PB8kR1hWNZ9MOfUHGhRO762xs38d8QR3
y2KdlKnPs1eyH+/7MZd0lZphBDicBLP/rihB/1fwOi9FDOxJ7K7nevaXdjW4W9Ds
T21QwkssRhfghd+AIhF1yNkvwxeU2YTimWHWXXLXMp2FY1VGsQETJX7ROlDtNtPR
pn+0hBpnQW0tZ5jlIeO/Yh4fBevz50e3pg2jlritWX8ylHI5MyFl2i5P/EZeJn4Z
K4Bv61bP1eklnkgbbMGllF8YTaacRvlO/1YriCJI7UFLZJ3jIw/r38wbP1+dRGTd
d8xy7K/ZmylsAqrusa+UnH8HuPFpy/C3hbO6Y9TVmR4TsgqN5Ny47tNxTKaeZiIM
ZGt0w8UEFNLdwsxBTlioDOYfz9e0Tkez3NkVqiPGSN/OcX1KD4AOkKFqnC6unrfI
A/0HsxURqQYR7LFOumPGIb62ga4YSEaw1A4lI7HqlcqqdTMzk8cERNoBPpXAh6ql
fA6aN6ED9lHEgZgKDd7Mjsick9r83bmWjh00l9jflghMw1kciFAHvHeGGgey08Io
ApVPaVVszin+IUj1oCqYscvVancGhVpdVk/GFLJKvWQrR8RY5kShD6vqeQtjbsL3
G1BV3seY1gFHzxQbzIU4X8xSnnSYBoakatCrzYOv045wkm1NMgw6YncWSDyrRaH/
jtDLjtnY1/LLebd2Z16a0Pxfck/CcRbQee0vIaqbAJNX57XG6UwKSEmMfUDDeKEb
s9ZPKCFHzWCnhNUQrLqho1D7M4kcISLzTiJFImJCo9oZMGbBq0N3G5pfp+P7I15O
ecJ4eeEp2VdiSkaxsZH/AmKqMlxP3CUyYXd+8pMw+NWx0FPP51uVk+xdD6KWaYbP
bq31sxzL7ayVlfssQ3bCLgAFlFT3Co5ZDNKy01o1mQCWk9RKNTGh9u+BT5mWRfLR
jQJwoOEaa/09orQSnfxxAwpJ5tgUOIsNx8qIzRzlyENE2u2fQgAx4sTxA23ao7ms
BiupzYU99sGbnoL/1g8vjoAksIdkDYUUxat32LwUyB1rxMQaFzd6cKiAO68lKoOF
e+Bqq5firxRdvil6rcSGa7H7XyS5Ej6CsiTAa7HRTUotmvUz1pQMN+NVxg+upPqk
bS0cOVfJAIEGVHbvOckpimBxxiZrn/A2LIfA26fE5++d8d++Go2LL4BO68DDqxdB
YBlzXbbNArH1xwxhmYIJz1xK66v0UD4jWHt2GkAui80FhAr3g+lVWmCyotVwrQ4p
ZIzqeMJxW3waZmUMo0l9iK+avQRjIm4m3uh1nLWiF/z5ySaP9IyHaQa4G4nqvmUm
ifPWjc6CY70uBOYYDzrWNw05cK8pX1GU0QYM8iQ+EOx7ucH3oankx/cBeVtSZLn8
RqMwFfI0793WEAD/MJhnn0nnOne1K1WoKvvaQKCxcQSqIgsvvUef1+mRAUV4v4k8
SNWpKryVCPFZCDjshPVrgjyR9opr+49H6+gyQNbRHHJCSKVM34kFefaPnXDh7ar4
KpGbeSJxbLCeWT0hk/8uL7UhpGfRsCT+DbqzbxOZ0CtDSoKGewY7IgFm2L79+n10
/cK0FLDRF2nubeffyIq0OOBa3xzvq8qva5K2xrqeBv4JM4Qk5MeIkYyo4KXwGrjW
WYs/epIXkTkHyZsHZP8lbE2CDzSbhG/Cxfem57Yj1SmgSoUl7lCv2Qshr7qpmDRU
vnWyKV0t13hd+u6oe5xmkxNmp2sEGCesbqlXeeS6fCOtZHs6arbfBIydR5LcGNRh
uBX/uAkGITeuwOf/p1zXv2wI+ryj+S45zTX3Q0Veuyf0/gr3M22yR8hlzE81eCz8
sFV5TlXmqCja3rsyal498ekOIWeDFMQsqtVJ0KuFAxp0OIE6Ve4BvKZwcpaZ69Jo
F4Tr4xuhUUAjdByu/ODFFRTEltmTeroKa6zUlhX3sa1BejWBWiuXbTyXtzWLXxzP
GLmnHa/ZYAnu6Ce3UF+fMeGrvZwRRDtJZy+QJnFU8VXzmKR8yqUArlMQCqBo7LlK
zK3/1BdLH5OmAIy1zhtOA9Zd34KLjgxgUsAkTCgo/k3mjBIaqxxt5uR3YJUS6J4U
48F4K+p8L2JOYVerEGVJ7hr1iXUZp9DEZnIKvUEo1P6r16Pd2ZrQy+f6DkCpwVcl
Tp5q8uWTGNLNpRyjH88jnx0y+3AOrs86F1ZFVssXfz3MKq3seBX46zFlPIscxlTV
H3ZnXMmB2PfVQ3zdQE+xVvg+WMailpliDw/ECVRbvZdumxGvihpLXnYS3DXr0Y1O
RgUm9s5DdCMJb1BHGExMf4P+dhZUjLg9Nku7LRlHXBzwrCMyhZ8lipjuMrX+SyIV
2bvjRP0zp7Z/pMuuuF1nh0iU4GFTaam0ioKiD3LWIKpMY/meDXggfnZBu2RhPCJ7
msS9umLzdDd16j1/V8vvGcYk5W9+RA7h8vhiUW8DmoE99S2jvALshJt2TSY4upEK
aWdPzZY9xRP6G5tJTKApeOO+MHo+ZM1LCsH6oX/tAR2C6L7vWaNjQ1X/N2PER35S
EDcbMM1XaH/2f3JfqiRjyEwaboGU2L9KXg1Ii/9MKVXBjBGnRP+qFSuik68t0rM2
zHfxfE4rCBMMe2uUVghqOwJoh25tSazNfOyO28qWyR70H1Zsaudc0TIzdjW7teSv
LlAbASO2QDaMXitavalcgvyNJsd5F5mxih6va0U+QKpHSIvzw92B6HlB0HwdZhVb
hX8R9stab4645jNjqthxMo4oGqR4TEYPqr/BTffPgerF5k/8mvvcKBv8eoYPrJ28
KMLwpTuaUimX4lnh+ZJuDKWVfR54ijKjT9v5NUAf/WvphH4ATPCXfhk67U2Q8FZu
0q/zjO6nothe3LghqxLRJz+Yhi8wotO46TR5Vanw0RYv07CxEAxtaL79Pr8d7zNV
1t0Y9eVFyzf7/ODx+QFryE1iduUTkqIaMycdcYRMIO5cB3fAHdw1CctmIuqwkL9Q
BcssOOj8SeDf7N0moQWSB7TRT8JpNPbFIW6EcWP7lU7/lMBC6xpzdRUhA75AgoTs
ccXCXPUXAkZw8MPIFwAiSRnCvwoIw+Q5jf5StnEhqBp7GFEwr5De2+1BiOr5eyHa
0PWOiU5mFRstys0Kd9q2UNZgyI7CVBD+rhBR2lROxkrHgmK7bgLCO3NSjWOh1cIQ
U5Mww3JsKGfIq7ud90zxhNQRYnCyoRhr2ENOK5hmzbHjblvM/YWakYytCeob1TQU
EgXKv2sgZqw0R4yRTbIHYytI2NGieyt3obrfgZXQXXw1quGUjPku22bvTSw/9bSi
ieyiCnTWl5EaJ5cjhCiUbK0HtnYOsLkjxQUhP79rG0ITLOprAyY0qNBoL5Mc4kzh
ciPib6SBEv3xST1BO/BO4Twz4CTDJACyR82kSpSuePzREMNb2Jg6a2E/ohe6jBZf
HltCeINA6YpCmMjlC+BikEgGSue6Q96vibaz0ClE2WYGMC8FhWUydmh+OI/Rebr6
cRbgLlsfd5Ah7RpS5r0C8pAreM/XYqgJk2SUa11orfLHIikRjOO9nSPcRzWboMkV
+TUpZMwA0wTSsAfrWV921jFTcE7ejNCd8wQ+NeXxrcNshTjIJ+tA3nAw3yRlQZjH
xPPm4m3dtSqs3cAlRKElgV9LB0dCnCQHpTQ+Oskn5LC8JI9NYGjUgseZl/TyAtX9
rrZJh1REiozhb2eTtE0RC99GmfzdQT64fIYHT9ZYoRKku6ylYR+kxRyeRkTEhAMI
lcLtDzGhIa5eAe+/VuHYlJOOHGNLwsFjvRA5F0t5eA8mrKhPjP3CFzM+MCNGPNCe
4kqZQaTov3bQCk8ZCClfogsZCvByyc927a3mAgy5UwbFalE8GlaPJMsjUQ3y9edX
xXeMzcXNhwjkrTp7KpdUG+K5djzp2LC2mESppF1z5dmb6oRHq0rcSMUvemXDDeLJ
49MuuPbNNqq7W77d1RJXJJ+OsxRvlP7TsannFDpllKfVgSuSAwX3nLXyO327c2lS
yHcdHkHRmnHeF+vMTv60/X6IXBCmRd1zLmSHMa64lLo7mFpGN4/YNYK2qGdVI8TE
Y0lJY+rrTp6Rvqkk9zBdPJuAH/tFYCY51k88GfyjDaUmo+zY+cenF75paCkDWAQ4
goj0Terd/79zIDW+gw73Vl6phqlDlXD6xZ3I94gSmGAEkyUaeAg2LCtwEux5c/if
gHUNlhXgiVriJjkigsot33kLJdu51Ut7hheRZC6Cpr4shWtbK8QJ2YdJmz0JAblC
5wNb6ddWXCsTmOJhutfGyaZS/TBUtIJV4E7gjyBKyKHdEOGGUkh2zV0xpxBnEhVm
FG15jam78g09e32ZDJvghhA6s0fdgcqJJh2C2SacOqledtQAoitwAT/RtR5oT/OG
vSr0dQ6T/xJtyOc7FReSBCaHVJU82WKc6tNuuqwWJGMjVwjEQRxd7yQ7hFUyjyEo
9Pe67VK3q95lgSkg7WzHAWRT+5AA0TjeuD0ghpxVVKgzigCfmUqLz0R+9umAFsSI
1z3rUxZaAdkRGrlVXivt/8tKIvwHSu8XDovCOt7dcZbWLfuU5mygCQyWZdotX/Jn
T8WphAPrU8jACCHMhfO9iDDIeBDtu1Z96ngC/vbN/WNnB33yFhHsiTEUciGU1gGt
avl1VWRISI0+LqUAP8sJ++RaXDZCrU9F2DJwrsH58kNGZop7dqzeVA1JnM/t2w7N
AWiWy7zLuAsydNn4aIA2Jf5I2JZbMkNtA7y2Ah6BBXQzpRC+k6oIJ8Y2UpOdB+yN
2VPrOkVe0w4i46AiJRmDbcUQEUzc59m7BHWS341Lsc22a8Nl8wpQ1U0vFlFrCgR9
sKr9FhRUzUYTYbhr8GKm4ZYEdFVw7div2ERtrZZ/zVFpuTMC1/cxD65j4TuzhA1m
I8jgHp14ACdb1fT+3ed952+neIQ070C9gfnXymzxOb0iOTSxSaWFnqX/H3Tvn6WD
7WOQwrZdcgQmg+fJcnS+ywDyOJSF8C3yb1UhkyIEgF61lefwttDeRY+CsPsk62Ot
1a+wTsuJrE/buzhtZR8k/Q3Y0zufvjcMTmQUcCnePLfj5XYsNhxh3f0ahQQaynbV
yJjYZ/3HH08iYlslbG4CsFlpFUe0SV/5vEoI3+vKYTEgngR+8vi5hoTJEhXfRq1N
v33rP7zbv2Y01tlL/5++8CWzP3NxaJAIKdjDW5CrnodpE6m2EnVFU4JPO2iDA+yg
ETd570OfYRYQxWAtznpZRw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Wqhy+esXAdfCsUzn8l89DmW2j3VbAqoCvgjwI7KtqMNmIg5dbmZKn1wWG6a0j5tu
pMA0D23vwTXqTxnq9kiMZu0amfkKAUtak04aqh32tqZ8cgw/8haHSmuWne7N5zlD
Xm0PAY6s0dgUzXeBj5S/4AMFWT4u01Ud5untu4IQKoloSSTobPzZIHIOcQpIRNaa
h557/6bdFlpddclkmGPpz164ySp5FZhg8bcyc7n9/9wwWzpIj1tmy2wUJGiBy3BF
f3CbbksHUXT8qHImsiC8a4D9aIgPtyk9gyUEDC3SLX8/q/J5MkAujMO0eJ+Tf9v6
3eSufUPFRAeqSmhngpArow==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15856 )
`pragma protect data_block
1LLluVo4etjsm0fgvIujZMu0LFKz3zQfzj8Nx/rHyYmQn1ULpa5LWyF1BWJXScSa
0Mvo4ysfupRyGmWjeAmYyPRlBlPtF/SNmGx0dxkHhcaEfKyAyjqacZg9hKwIOtc1
GOPKu/t+KpwT/OxTJHpwZ/Z4cat5dSzAQXvpST2gbAF43gHfcyM6H42eqKbnJDKO
hF6/xaUoPzSSPSAZP1L+IAKAd73SzNLQgXNi23c2f7JcRm22zmdvifGhGJT9e8Va
O65Y88R5FvQCv5HiDt8egpKqj/jTPn82yyU5nbSiFowCkMynim8FNVw0MujUt3oO
Cuc8TBrOqhTvFkesMixNVnYFIxA+rPdu94NrUyd4TsXoETClRnVzZmwlaBAZJweV
VXd/RUqijO/xDXHzgWxbWuWRzT5rl2xWqSwP1XLquu2wzogFxWnhtVzMW4L4uojg
mLkCLMDvey413U1ByO4WD56pQc0M7cXlG1SS6aPoIvlGGbeeMBp/eThWrp6J57aV
oV3vkkEAlp6JUglhYl0D8kVtPgugVf6gL+5RK1y7+32cJCBOpiq+eGBb6nJBlU3i
MzHcILoEFXTJR5jZuoEuhhhLkce8XOgpGumG/bWEzswmOnaDZYxRIAryi3lH7gwE
uHZ63UfaXVgaG8s3pOkN1HlYq9Qm+fqhB9AM0HEYkCO2G4TOkP5Hqqj9GM9bw8K2
zNu9BPH5ZEeYU09320023rfZUz4kw8Zky8KIORRrJNRHy8mIA2yI9kaIOrNweHmK
UNhl35AI4XXnZ7WqQt+gdXSlWodscRaWWJCvn68giV8V9LWC8LhJnY6cWlhA+zSa
JWQgOhNlK7WMZUsIsjY3DIYzEcbcMcJU2GlK03+zMnVQwi7yYOL5CVwSu7OZcTLx
sMXQvTrQoVspGm4fEnUBFvetP3vMnIjcgIhv7c6Ah/tMpBLsDKK7GVFoaQHOjI2B
z8xOVK3oj4dmK3eqzHZAeYfdV+OxJEX2pUzQAXo4baFwZmNWLtHkeLURAaAG/t8+
MRA1mOgzmGUeIRpS895om7IPJ/kZ68XMq7ZJy9ocEY/jArz8oPM8hjue2NyUOugY
H2V2GfuQDgCSG/NU5O6aIM4ZYVqgsqavekxPS6dLFbzMObS5+e8fB4JbQhVjL3nj
zUCNMrOGqEYyydlbw0Wsm0HGNHhKu3qdQ72ZpLa3vdGTIT3vVTsb5J2RZk2xZ+Lb
mhfIwVXEtd+u1HwgR6Q1rGPC7kXV/A6CAFWkuCBqGdG4PRnpmqnRVYavMAqxi/7X
WTQtGPzswszfXH0nKu4KNSBtS1yagzm/ymfkhqA0v2g+bW8B1mc41dfambI9247n
MmSLpxAKqL8pTDxZK49S8hmC87GH+gmFRF8QPaKQ4eu5kcFBf9Nh1kDL9Wjdh40o
se26LnMUu81u7fQgSM/Mwg+pQN5ZPzi0U9ExijM7qrIYu/Ls8ZvqGnY6bzuK2+I5
KE2sJKIQWvaFFk1foTJ2RX6ote8oAYZXwrXsvWm2vPGoYrT4a+oXmbqGFatgEa4a
Z9B79jtHluNWPQfvb0kslH9ev9bfM/O/6JsbYQMTIJN48s8iOF4OsONhmU+ADuau
s53IpJrOMILe7Z9mXOspxLXGiJdKg85qv6W9N2b6yEf+btEwwnLxbb6hn31kJa4F
4miBdJaSfgwzHiahM+o8vxaw5gJxJiqNOX+YH9t3aGlKq3ClnUsJ6o69Cve6i85x
nIkun2Br33kt2OLC7mzY+/ymUyoajCizQWo5AqL03Nqnjk/ULN0vMHwO77O1fhbr
b5zanrMf/MtUF0TxoUmmVEcTfEQfEri3WPbfRfdMQTvBBIolHu7S7PyTPbFFOdf9
u01RMOhqfzyQGxWBY2IXY8Z3JJHX2i+i1mPQEdQ8lhxWb3HFCYcrquweSwooDF/g
dT4msworDKdVMDh7fdMRVCCjQiYVffBclVsa1j6UQgDbD95oy/Q2KQmEEwtDtxBt
C2xaE3blH6Run5lUnka5u2Y8mL9PX9AK/D+jy+FaLsGXJtr9U9zJlTeMCdu96x+B
KxKh/vz3t3ncTtUUBeLrmhaJ3JH0KekHGgxc5SiXtYXU5hyY6IPTpAqB77bY4RuI
x8e0DLmIhebffqfVar7K/KHW53Nb8u58qRm2/80OBuJ7moKcxm7qdwG4aKIG69Jk
TQTtYs1GN0GQkrqESSLfcufpyDUh5GCdaf6305gNTjG72bLuboZViyUbzAnup1wJ
Rc6/08aD7hoBaLlTWCQyETzC9bpelwC3O0gg5uaAZ0/11HKza+3ji7JLsw/LjrxY
7/pORFFw4KB2W+4GdQV9aUXQU3W6XWFUsOi40YxEoaScBRdhDxVTKNTbKO0HA+wB
gZhogmLD/4Nf3S7sLN0obWLSP/wTSxlb2Ekh3aGw9moHxQomYz+Z9q/AyfYrVYB0
D9rGJgB6kjR8pFZucb6Iy0NFGSwZPMrlWJsgFOlbgwVV8pjpKzVf4S8My5jtFTLN
EkScWtf4bR4ILn7eNWHZUZS+/agzzf4TyN9TbPRsqrh5aVBJQSl4x3+5qYdZEIdt
LBBwH22sTGeWLYR7SPFostw44X2TcdLm6YeL9HsxAYg3+1KdH4yoBEqUYkDNL5Hp
Ha/GcmHsdbbunMqyP+t6bm5J/5G91j2Zgz1unLgjh3HGlT36yfGB9kMJDaC4TiZ6
QcJMINeRuzVyS3ms/hH4oh20dOlLyjjWHHvjh+dsxXMgIu8LhGOnWRj3ISJtsfcW
74qbVkrf3zRppEpwjxeTwXL7xLYalvboGX02zTaOE4CHMAdAxg1ZMaszMnAutzKY
7nNZIAFFZwYbj8SRK8kQ7HjL5/nSXEEhPsM/V4ZRZ5V6kFcMPYa1jsksNjGgCfWs
/z9eTnvGrQpZ/WMSIlnbm7hQdQndFDzkXkDGRsavlyrD1BxM1GbLwKHww/2eJHmt
aXoek9szhLDs87pmbX690y2h+2QHybg7WVT8cBSyh1T8hGyJPG2Eo7U0Q87FSrIK
z8sXr2x92WVZgjn9/JFgIUV+sCkaCQDiG95ikFwIUwiJWfSjhkcHH/P7woCmJrrs
7lNoIOW+juIFYl5uvYXfff7pzoKz7usiBSytyWn03PyzDIT2QUlDpArpS+BxNzP1
DxXyRZ+hplRUHsSUUf3f2JvIVNYVXGt6B+3+fbCUP9Uh/58JMIRaRY8GpCUdAxPA
oTsQms6sR58t+RxLeqB3K2YwbRmbBgbKHjepF4y3X+vei07EATEuYosh/X2QDb6h
JaBpZyZjxdOvbdbbP62QEJH06Nr0czfmbV7rhxporSQWWoKqNgsIB83MDHi+/toZ
pYBzs620dPdl1rQCVQBv1e3VbZ+TPSt841MFX5I6kKx+sdrwW5R1/iNELMZ+2ccl
YBX4xEAc+r/qC6pyldJjub6CXJ6l0pJ/ao/AkxhdqkWrTUvGtmuHJibSrFO2cyg0
f9LUqPh2Kuu6Ll3VvKBe6FO7cJ3LRn8Xif2r54uBodCOgqkqEarXOGbzdyDcX1fY
lYdZI/p5Pmy/OBzT2X1y5aIspoMetWQybwAK68t3Y5IH24bJQbPEoVRDPS33/nTb
RBzn9tGElBPRRSoNi0AIs9PxVWptbSetXZ76Ow1TLIzgE6chfaVmqr4dDFmSc8nv
d3iny8ONIks0geEuWclBebtRCP/pMXVruwdHuCmcXJNQEvJIbWUdHKSTsFUpq9tk
RSAtM0qUI3GVP3BOixIbgpSo+M3pzT1zJ6aTMcS2jANB7XDIUkttFkwCW2M6c9Ci
Inat7bcKR9/S0cDA2BnThYPyqByJV2M7mCRTl3J66lku9zSzwNBkOu6aogxH3DSD
3GRiJQRy9LDA4iXYN0s0qceQmwHUSQB/g/fTR2k9LYzcUk0hFMEfhN5GDlhA4fBO
Bb6sPOd7fZ3638hCLJpXfjFzX958WzqM1t9DPuu9Z2Lv6XCChFObRiVr8WKUqJ6k
M4geInv+uJqsgFK2HTcbJ4zrVYVpGA82zxxTL4mT0FvwPB4BWM8ohMgsOpnY6F5O
GoQhinmVL5R3xy37AnicmyMTmpDSs8z0eRGY2VPe6Cduqp0JbpFOru76wajdXi50
zVAiv1qEC+kgXNEX8ce6Ea3ceKhXBOKoUtMoFI/oMc+/63Kcd5zUFmyiEbuaSYuQ
+KHGAkOeG8sqJlSZBhUvf3KqJ9M/PMYoKw87UfzLRaFgQukxM8h6dGkuxD8C4SqP
JcJ5UtG0yU5XwEwDcQB/cgMOsIogVk+kN+btQWffPkwGLGWMSWmonz5VmNhI5nx4
3OurZs9ywlYvEczqDnw597+/ONJz9F5OMd2B1Je9dEXma82hUfTqPb+iv9CJIsLK
xhGxipRikLx6cFVgUes8qRF6knZEmB/UNT+Lm5XcFvdMBNur8RFuNQIKF7PFakmo
Gv4t/bvuBTHIVUaZ0wlUqq7S/VPsvCxIUlr5ioCAt3fc2brbPqbIdwKwQ2ji5S6A
1Xe63itFIKcDZavy15LuZre77Ltnpfs0vOYZImQCVTWVa9Ebbafo7IJUzPNk/gMW
nxpomPtcRK615l01DjwIn+lbJQMbpch5310CUAW3EVFwJpl7KvSBaSDnWyicHyAI
t5bd103YU0/8Y33HukkJe7ZoLKYnuya+eA/mX15iMwbyOEnilBS4ZhdyxeYazsQA
vP3sPTExFNwULsBzGSSm/mYZbwqX4lvNjLiNV7K78zfmrktrTZ4mFMSlUkATwupK
hgY4upnPoO9XDIKi3+wjPOLFCnsMkPid1YNdeNRljcvz7usssTrr39u6zq73UFsH
M+Tt/P2USz0Sh6z05bU+e7O07oIpbpnIWu1frAc06OMlwZapLeM50kuAREfGYx7X
lVIaaZWYtWF7XFiC2ks5+caAOBiZtqQPYMU033tO6kKJEUYJUnqT0UutxGBeI6x5
UgbuoafHWZhMc36ekUR6kNV+F+VHsmvXWGQgdptzKcFzr/kp2JPtAImj1/5RLZB/
QVyaoTH0nbaugzg1vh7l0vOdZnzc74mI5X2WiLT6IePGMIV9sUpKX8v0Gmw5zlT8
bEqfGx1w+CNFhHA2wyX18ky0rEOpFCHUc38CPLrHWH8UKCisyN8ltPqmesn+jsal
ks2GtGabHLdT1rY9/DZ7FlQxf0vBNErbKVHimA6IdQb3JnJhdx14SSosyPFCbF0s
5DHNf33EO69w1vssEgmUxCl79HqJpCRlXItK8rgoe4Yejk3xX2XZsKaw9GJtETK7
7cu84iVKRG/BBTVy6i2NacDnR1+oZUWgMstQG8y0geBbdTUbfUfY6BdTUZC0t4Kn
dMoEVaTGqnI/gF6j0F6h/RjrPjgSljQJcImu/RkdMdq/b1RNsNlS1raVbeeSsw/y
1K2GZOBi5URqPi5ZtpSSnby0WttYuZKTl1qA3wgPohiJsBL4QKw8b4BbFKBiny54
lwYeEKPoxeDhz2ttB+wgjVcUq+NO0S7GR5YdBnNow5vTcw3LPm5/7HjufGlQ4ADp
i4IrHLoEi74xPNo6zKnC1lXbTcWuGQ1oz/Z0QUbIkTpvOuevgahFDeE3pcjtVOG5
gSnBHURyOiNiiHTlrMv96cIU24VyhF0re1o7lLLNEkOG0u0N1xwGQmiyK2UIouLg
l/oc6jB90cR9bNZAn9mKX0MpSpXu7RTDap4GepVNyqT0aJwARA9iYsvbdfWBVA17
Yf2kEypk+zrHLve3BekyX3GO32QKs4Yhf2RM9jA4WcbzfxLF/UrJyKIsuupyKwU8
MkA+ti1OyTeOWUPpkY8GkEq7pJtrxjKtBNBzARzzF20S2Pc85d9E+3UimMxVtG4P
AhvNPTUcd6ZT8J/89zcE8zGPqRuKmREgLJ7nLbQaigdCMy9GPbp41jIbLrjVBDsI
9N21I/QiODctzvp4v3cLsLjoMDGJQ2sCwFq9mHbUIPi3CcuM/F7/gXUN3cgaGV+s
5zOh7L+aNQz/EhQ39hVlORR9Nt544i6RmCnEuRPvIn3YKkB01zbFQmz+degM5Ukd
FuJronu4W2fPChhDjlmVRooHic5+0fb0Wcm8LC17En+z/hxYHUTJXaJGMFc1rHY4
kIdurBqqRinBor1SWBP+jeLr9yhHxO+C2op7LGDHRrhaHYOA3cthXp2DSPA6dQpK
UGqYQ8UzE+t5Nj2PBZW59zrUcQqARdaq+k6CxlDc6se3bK968lhGpCqhPrVqy6Dw
e0acfQB65GokzxXW95qyfddKu+IZw/16OaejbgNYIyMdMimziTqsJ+vCHrQ8DeYR
QSbzgprpe79w4EK+euUSzyi6Tooa4zdC/mYnFhZ5WwhqERhG1vc8mKz6wHClmlYG
GRftWnzaAGnKcYIkaIQ56tg4uMnqlRGg/BXzvRTr9FkEJxfjGoUq3U7Mse1KFQjm
vYZ9IVjPuAirX9DEi7ybj4qFlBU3YTRBoc4O0vSEsG2DrIIGqMkbR0fcc6ow3vSF
kx7XQzD6rxZx+ex8V1eRzPagoc6iRR96hjRug1vSLot+uGmEGrqP5/LFxs7XU+N+
qoJT4fINF94kXcNcz0GcQa5xXmuQUM/gPStqog4xuPLqGgVmysPksTy5WQmU9g0f
OcjDIP6U5vbF7hGJbT7xpnbm3ee77aZl0BX5maZu19wa4zo4klGiv6IPnfW5TdvH
KViz75Hl4r7P4zQtaLzgoDvRJhraJKpQaKh+suXPynLw4jefmXE9T3cJE9ugb0Az
HGo16Nwdhh4S2aADMMTAa+R2WK0mzPGmRaXS3aJCTV5IDozRseqbv1MdHQ1p/RGP
/C3AfP+fDDhaEl7heNvtahqyvhsTB5XzvYRuBDGw9NO/VX74l3EEF6L/AHc0JezP
9F8iptm2tXj9aed8aen0HeImIeHcHQ2WrRHJaxXU52GIL2cLCOskaSDSygLh9yNg
gOS/AcO6qoKdtzOy/fIDTru9NFjZgwA6grpGZoOl0Ih9ysuy/+82f0Ix9JuD7sJ2
0jaLuoRy10kzxlQ7i5N7VSZPMSjiC6YBx6ZUcbxfsfgTuchUJeyOzvL8e1GF+8Me
qtD73BrhHFFP4V38NGG8a3p3h4DPj/Sp7kpj4r1GgzD1JOi7YFTY4xHPnUAsEb9O
qZS7E1/qtfzjATOOcnuYwz0mvzv1iTTF04bvd1FB2MEVpDPwXTaSXAmTuQ8GewTd
gQMBLPx8IygNBkKz/lOa66Do7YbDQIiKeWX6a9nRYkuwFx1AI08oEkS1F/tM3ikR
aaCnLxINNUyRVEzkNbA10oM6fSRch3Z3w73t5gaZV+DbL9gHlKXB4bqqPMWF4hVY
k7tguE/tNGXD6jo8Dlt8OL9KOtBtVEDdTib6ljWD5VK3LSJt2UYOZChg0HuI0nER
efUZdGQIQbAzui8yUbnfAQYA+dK7eAWVmQDknjuC1JxeZv6jcjMeGleLkxGQLQk2
wrLurug5fYkmjBtzDKLFabhjn5XsN50qqSaDlWQ5RwBqOfuxMq2khuAcGf826+e5
frKmzgfsNCcB7w75K8eiNb2sEyh76kRiNZ4xopx8vLVGmwoyR34qrZObkmSYHQMR
sIBtipTDAmYLAP85PA6+hxfg0Kyixr6NUPNC3q7ErLd33u0ZbFpGuqQaIqPZInX0
HWJ93J3Ory7zsGfJBQOj+CpZ6/VE18tgewtavE2YXGGGR1faBzhQxYeRE0nWHvGm
lXvBq9GomxECLZHLXaV3vQ0uvqwOFm4SaWNvQidpkXhyh5HcuNNK2PNiKV80x62/
LZfSwzdQxjuzHM/tmKJfAsSBe2Dbk01qV9tlmQp1mnbscacyJ38GuQFg9WWR3whe
yhaZTVaiG4/PgF4UgdKOBQ6LnOWhdcOTYIuqSyRsNPCnlOcTowwtLzjVvLWsKAku
LPzVW+9dAM9kRSNHUEUw51ySk79eApH6qYUw0g8GZ1NcitVPXmK7KzICJ6q/w6bu
ooS5nBRD5lCgkcYkhucD/Gvp9dhvS5hh0TZU8QAd/XFsrALyLdQ89scpceHFzwhG
9T1cZHIi76ZEmSePavnlKF9a/m4dPpo/qtg4NAHEMf9e8Zhn0DpGepPSOSOHziWw
Pitk5dNC+2ZARFdylfpJ88N0gQgLcjfJaBk/MHsrHbNRKlRWVy41NpEKmtxssEMS
GWMpawzTnHI5XZsZZ+LHWRYTduNzxLoPHOfLoFpy2KTipXPR/9HBCQImQy9ALbSe
d8S3oNeRw4QbLtH7LeeTFb0peI1SuoDD1Tvw0hqhqS6KfuZQgXzBRw0TQg52+K8F
Eup4rOpM1YZphkfXoNjfspYGLV12dPOaGjgPyFYoYnIzluC1LdAZLiO1FNWKQnNm
TzaIcZ1WOnwVCRTZ6KjWwgZdkhDA2FWedtFeUtR992/KXG2p/TG2ZjVr9PPUzjM+
XV3gUeScO4k/lIT6opiByB2cK15zeBwR27nhgI3Rbs/IU787O+ZFpK2BycNDs9vL
TntYnQnA3cpWarZnOEZjGXxrSBcfqjGW06F5rzqr99xD/6jLNRD7NRc0D22x781G
jpARl3FGfNjFZRZi9sg+qJKU73y1gFJrOKFfFtDHFfAvqDRh0HZVsCLW1OAMoyxp
wx4+ru/WOR3Nmm1O1bow7jTjfYivBxirjDBjEG7adRpQh4EPUNy6+8RFGs4JpaR5
ONvnrVKkY34PC3JHqNuHp6cTcvXJKzAr0W8cpyOEJhC+FkRVDKERBVrqz7pZgCHG
jhNr/M7Mq1UuOYdNr8jAh5Ct37xhoQX+uIyqB8dQjdB8kIuYSzNKu0cEqPIwrWo/
rzqQRhaRvh5JDV33JnJbPqU90QHK11s7A6JEqaGdbEX6Hkqs/6BCvaFUdB1Cc+Da
gV2JVqRVxflR6ztZFcauXCZsZKvzWx35YJfhk0vYcZN9sP2fw8b3SNKcQbWq8skY
vJkBayyDQCfY8OqsZ6UJi8h3c86rgp0XR1Cs3UWc4zRJ0ANlilzx79A4IFJKz3wb
0LDyBD09aXDdKcE9OGQqno8FsD/0Q6HL+RFW5PjLAwHdjIxkKF/wxGQ7c37Z8n0x
8c71aA3QzSJahSzp8nw7GlQBPQvWtvmPRQlh8zS1sohxh+nSsfF32dBvrbWr20tz
AbxtWmqWlgopmyBVs67BXef0W86BM0d6krw1a35QTYwXV83Z4lhb+dZOt0ApgT7C
Tm7SzROS6xb3kNyc9u2USpoMPHpq++keFQ5Yltm9dt/4wXthRuUuwHhckn4/ag/f
iCa9BtqrYwmVrr6RAEdPGooFMgyDWTbxsfmQ5E4Z9MDIzFOerkGreNO9i4PN9lXd
65XQNmvICZmHmAKUcM+r6Kp73rCfETSzeXoljD8MR0w0TxCIhKk9BVRu8vL7oXft
3uh0SCe84NrO4p7Hv++OLxtCZP3Agl66gd1vbxDscf1w1bcwDkvutkYfZ8mJgfrN
yBhRmcbLtXhIoenuNqUC5vxIUqKbRKyZHrqkfZL1wb+5Wy0+EiBTx5EgQO581VO7
JBkexDSk5I9wq+loJUUjCC16E9z3nR7hGv2YgPmllwN7slmOuEYxmyPs/8kMVG8x
VVe6LpnNzi/7tSv5ROzzzrauoBbeUFC/3ciJ2RUROyBivwdXNtgz9D4WSYu6wosv
C1YtEYZLFpYPRltbYytIDXj7Hux6p4LI1ECMo8C4DlUrw/dytJv3VFNsD40Pn+ma
mT8wLk7E7tcDcm1xfcaDzlarlvzPQGGOWNY/cgWEOiAsgvkursmwaPs/W05mlWNz
cFv66/AH8TPJufOHwGHpE6fNH/vidJl9pybHv3KNMler0UUz2Eec2+p62Fycu8SF
UAcO+hNgod9jQxvJcJPhoEc7Y6gwtFHxvteF5n8dwFx+unC35Kk5DKNMy8OsQSqa
qYLJKB5zGo2a8uV0mhdZaeSjpmiMMlz7gOZxwWb6nJmai2cbZ3cBdojF5AuDi+zc
KrOHaCQmXmAtzl27Hm6cF69yXuAcpvR9aqAmLGE21KsZi5p68sUSEHwib0tORdcy
KEoWP9VGqc8ZF/5l3DxqL57dz0hlW2A2HefBY/L8ZcMJ4VDwQkXcxBAWqwcw7tZB
r1+PXoknCPXeRs2L6gRXcBU/rSIYSDC+/xZaZ7uC+tXOVs6VBESv6w92Qgptey+W
4tipT8emtRpWiGMy2ISXOovyONMVDr7Z8ehcR+/oJh1ZAdQVS44qv0LJ2pdJPWoe
85L/8w2X9Y1FFQn9t+Krf/6J3imKIu2JMKDdJvja8RsjmynJtpnfi1u9P4zrX+SJ
a4IudAH8rSuSGZnAtFuqMBSpCxKyKt7Tzm9JUWde0HZ00kQ/4N+32uGyLUQCv+gk
o887O04skr/5Ih17jkQNgydKrfDvWYzyHU85RSKsVEwk3qa02q/G0WJE2nWDjb/d
n9Apy6Yh5FO4zDt+uodNcVMtBmzPuCiRBmK+lzBVC/TrBFaii2dkZtgp1J04AcFj
tILpFFvlygVBUfEIiwYlKgWySmxKuJmWllsxs0vp6BYzUVaWShy+jEjCNKlytcb3
UHbKaQm9XN1IqbTlIVS6fChSe3hhPY1FTGiGsnXUJYveHw5PRBMiEVXo1t046oas
7HVZ81Yqh0pCZB8EXXwgjrPyGFhZCaMq19q9C+wWfM07qjrs59gV3ewX6Utz2Ecw
xbPd05iXTwEbqIWGABqDAsTqS7lGgSKpQDXBumH7NNl96Rh+i8wChdVwVFURzQys
7FZsk7jY+211oQuaLfcwJ9t0QRnXNPq/ZbN1mRii8uJS4/66+pso4WYRrRhL15pX
ImP+TcXLTHlERl5izIukdJRuYDNvzEAliXkdm+l8d6JCbKqxkDfU7Fe6x6qsSPvM
6ZyldZM7daNPHHDO6SXsIK6cfO4nb8f0CWMjrToF7dtBHMhatLa6lOmUeoBmGqUm
HlqPWj7naZPtSBQMx4ATYy+S6N+XcygKBichm3rgBwejxwGQvLs34UJE1r2VM/he
h/+SUQA1Vpk2fQRdEvYvNzd+hF9EGF3kSVg0yYgo3F8sNwLF0pTOmUgnvEdM5W44
mmYrzx2Gh6WIpXgW62Y9MeuvBm8HI6vHA+VPW+v300qQGYVqImfynnYIj1qPhUu5
jT+TRejXE7HiLeDuEU1JMlcHddez5oqFiXKsDrj/KWncgX8rBmCxsN48ZsaXg+1e
RLcDYY3IUeqG/vXZUVGsO5hIFwht4ejYfPA9ugx1vxT9RmJ1NY/sxG1ci76WWFVp
1xi/v3hOdfwAUOUlqsXGvZnskk3CctSZATGt4W+x+eGXJnYEFJ5GgcQK+M/67WNa
h/czYfDDjKgR3tTiNKOlp7u747wyNAzvHZiocp7gRWte022U6YX/HBWErZzycRYz
6mkdyvqATeGA3UnuXxJAfoCEzx0B4HF8Fzrw407bhFKstZcaeabsDqVbG9vTeH8e
euAw2RLB0WwWU4OFBYABR9vtnLH2EsEX8rHmK4hqaBUdyCCi/lCmWaPvOpLXJvTp
qHcYjgw8Itbs0GnkaF3hPfvCUQBMy6MsW5C8g8cwE3OgaIOlUGWhhL0hzQmJ3Xc8
DpDrvnHfqbmSp4Bvc/KvMb17dydpX1wlnNAz+zcO6n0DKIwUGSazgk65EzhYCLo0
SPN4VTo3VFIK/1WP2sGmNxDS+l87O2nb79NV7wIN4CgayoUouIHvtVnLK6vd/KAg
fsP4msddZN9Jp9R6bCs+z4rL4UOZi8gDEJmA7iIJBXI6MAUnJE4MGHn/w/CGLtvR
j6DIE6U+UYaRK+amnXMN81mxh3cRYi0dfI1drXXc6AFAeI/6K1caFICzPSxjF7K3
ocno+OerlIvZarnALDBkYlrumS8Fe8HD/ycszxIT3ukp5GNgGwSJuhYRIpmYH3+U
T4/FJfmQ46Y1E21G6xjjnvRNWRqtuqv2I44HhHZQIipvPCGIxvbuYmhOE6w2Pb0h
Upp/LWidCJf9Zdgj+Dj7Fz452ZWjbNg2NLGqbTAtViXCFNfKaD8sdMW5x+wwDOEd
7BX2+fhXMhyqSQINbHGDap4QKxzXsxiWYXh9LTCnXaEE0oKLxY87wagghbDKQNae
zjj9h+hBb0+owKaJuv156lPbvN88tx6Q+tJxKmpUcePTQui3DqOE5hF2WJ+Y+kDR
Bkfe4vyDFe5wHf2szQ4E6M6iBhaY3yzq44yWFXZxsyU1tFCqvWd0hBf5A8xrAGgH
2OPSeX17LVIvBIrkzjO58u44Beh22t9toGnONotaD1xJX3yLwh9kLRMSEF12s61x
uVXs9hrBao76iNjprUv2+EzVgCNeRLOtmz2k3B9+Ky1g5faxOoYGHGvICkE1Mdyb
US0OoFUJp/Vo62r/pHcwk73i5fPMtztiE6BK7O+jPcepKfqVqzFdFwIdcqJkSrrF
518EpJEfuJCyaaTjm3K8Y2eydoKnpF9XpUbOJAaO096gcZ5S/dZVNc6MDUDvX93I
ped3MqETumAD2mR7sCPBYiZ3bC4JKk/4SfFeipqu1eR5ijYER8WpN01urGZPiM8z
dJnYjA6A+m4kYfGZ0/jlXBRds8DZzBcb/R6SCFZAmtupYRBodoFnTYd9Iob8ftww
JnO2TkUidPAhEPMRmzveZ3i/oJQcUY6VS0yq+kK1o2h9N/bOUtt+VTDTr1Pk+kWJ
yQQvWVcCz38Zx5aEZlye8Z2iy4dUbapaDvSP4hrmbaZONrQF/57upP628kcDlJNx
izKC/VvM5gyBJwVdcRkZNy4S14Vt7zbkUfxzqHKRw2Y8LR1tNbfaGlEuvn2z+zKg
Yhc4vgtCyEFWXmw+HtClUJzctDifyBT3rytl1YYcNT1D6OgU5uTctrWYDxMLKwjl
SAKo5Az2JnQobsMun6DL5qcoyvWX4uCc+O+7834crYSYLqEc0WVIy4hTemNTVoJ6
GvU3ubnwCAm1egH1wrbYHsBws2zBX7Y/uUlMEXmt5O4IhsKFa1pu0xsA2x7MR9Cx
C69XTjLQ37PCd5zNRBPatKkGED+fVhRMZ5xMDNQQ5uUpA7W+0LIzxG+OD8+FEX8w
9uskaC9iySrXZcJRlXF83g0CLS4suBGPOmR6ShoZP4/mAcWQ8L5ZAz/ka9EvvOOs
stsDD0YEaTj2tX61M8PjOwuPsNDPit31xB5sVPMCSMNUP6hWScmL3SPRTqJAnJ3L
oGwbR3e5RVwWJwGkVL0LqMoAag/kKJeF74v05d3C3V+Wf1FQUPFXMDP5RM5cjIqQ
5FYJ0jIdzDq15crnsnxsW4muJT6CV3adsOr9c21e9zHGUEHPgtd5Mqeor+1t0D2A
w3hMWQHFZ2qjr3mq3Bz6aOkKWbVWvKQle2hz/mBAFyUzHaU42704+jJx71Z0VfP8
4w9ICC+5KGpUVXv6ZyqZYGtIGy0uM7b49fJID3DLI7BlsoMvXmRoylXP4uHXip2I
q3pSskt0f3oTJo8RRFsXyHKMS9esh3lWf6eqpwolIxZY5z99KxpmBcFWeY0TCQtd
e7aBpjWq01FZEG8bzzKFMpcffMH1rfzfgd8a7ykCjGgfnQQrnuVV1YU1ZFhI7Dzr
G4WR4P+ev1KFe7/DYIl9lyU81frlvWpEOUrjCGIGbsH8fxyRptezRhnZBeGBEVma
5qVxaDDquvcADxjYV/2A4MORXb4Ckrb9wPIJYsPYXPbHrhA/biVJUmWDe2TUW3tm
1TiJgjaGWvsUNz0uf8GpqjfkzdnDNUqw/IblsswwYz9J3JDZ3iHvxitUPQVdkt8n
LG20SmhAFQsr28Tv+XVViJVkP4rk0F+RfYggf3HYDtAq6Ne4Msb2YivV8VaXtjNu
LWk22zwaix7Y4C/bhtNzVdfD6oMAm3nRhCHLtokfm+zsvCRwx0xxMRiEtoM4jg4l
ZhE/44eboBeBjg+JqaA+9dcY64ZakeS1jW2w4WzF5PuQ4vzuAfsE9g7iTdCLSati
ZADlbHRIowPH4DWJySn9mo2d5qiPuNe0Ks1C1LlGcM+RJiC0o+QaHI37eOeFesrT
vnn/eiHWTW3KQQ7T4H6bt5UTIljfgBZ5DVVoAianAGhx/YrO0e8aWoiT8FLohHMz
HEzsXF6zEHwCS6OH4YU1S5Ct5CSc/ieHIabdIlsbkNPMMdu94QiZzMF1LFtsowyG
qbQ9lCFKyCCGD4bIpE3eImOrrleMcuLrrNSVg+Ip81SmOd3nMfmg0zPsROlCZ7jo
LlVeACmeZlxk5PkGVpEcA0gwR9vA4yvFfMkuQVEQzIjKuiT70YXJXhxoehHo0J66
hLtXmJeRAZkuASWvqD8GjGniKhgQE6sekNkAQMkqixkn3w+t+MVTq7hoRjQcZgys
Vyp+yU4mmopeVmNPnHJiEUMUgE63s2UH2y94P4MEjdWPIcx1LajkZkgRtzp4FRSB
7sGY2GQBsalBzOEt54rLY5d/SsPHK5B+OcHE6SngRiap3HAcn87IfPNvMz4ixyC/
Q9Ar6ttINZPhitJUdvQOD3KILa8g/s3EuhBsh/j68lQW898dbC5NjAugtkg5/G9j
DSsxh+q9LmWxiI0zyt2spela6yyJAqwRWr/sJTIEKQxF0OWEa3N/6NTbI9glhKM3
ar8UtvTq+JPyzr8VTy8ipjTywYpABrSXQt8+TmHB9G7++ANdqDPo4ZFOZ7j3pxsD
OKOxBKp9hkbIJhiUBXtXx47S+c92SNWgA7l1b9VZwHw7XKqBbLF1qJ1dmkEjDMxb
Rs11mVWSUWfod+tBM391TsnERB+H8I09TY16d7bV5kIFJ+aPKz3kbC4QVCiiE5GX
HluVYG7EV3Ch1OXPlp1s5cEBwIyEpu98uv+8pWKX0v9jeYCp5HFqJTT69cNNZJ+C
xzXIXGWAaJ12b0nZY5fPHOSK/G9nNGpDmMMyP5UI2U5vEb/ouoA1dEm11nSFrARC
QlFWhb5wutIWgnvTuXZdTuhq+YAPs92ZIDO0avOI4zSrHU8oGdPnm1VLv/4a7r5N
tNJoyqT6waaSg5s16JUFvH3mp+UHm6txP8z6shIrd53f/udvwCwJDt+X6heGQvoL
CBF42MdKwnaFF2e9Xz3uYnHj8g2tEad4bfkZ8Ee/dsrkJhxNIVe6zdDLv+VNKZA1
olgnHT0uPGg1rdqzzZlFhXJcbOu7r6ME12dS8bbVt355YiJ9QfUHoIkw3K/09js3
CMjRDm6hE3SAQ66b2sBUQy+MtvWGK8nnuS7ftMxxJwJJzC1eFnVak1WKHqFcOjPa
Uvq7YEsjhvZ0fy4DcB7XSygIW/yRvIzOwJg9OwwsaB0GOS1XQAUeSoBA8sako7Qm
hPTYQLo0mI1IBwSojcBeD9N796K+1QEOI/KTIg+Fnd9zjXP3peTNuc0d4vVUdymT
0YZtJCJsZAir5rJwdoNhhpPwDMQ8hXDZxSJxs3LQeSlVOUK30uErlLp01Kks262x
gsclBVt0jkdzvgWMsz5bKBVMOVTuqNHYJbepOdRAoT+nLlvrbQh2mkN1zVrzfZxm
ViK4lAtxN3v7G0970Vk7ovLV85nnM56xheGCHANSdTVgGZ5JUbhSW03WrQR7MxaP
Dl+nt3Z/y+dMsJFBaYMLO7T30Xn6YbjHAXTieD7WLZAcz0JybTFl6tE0GBn8vmt5
fQr5h95eGUtfHd9pkjIuMF5ESyk62ewBzHMD6uxZJfoKKYIeNj6fa1Pspp1gMdSe
Vf3IKMc/xfUAsdarLTd8YQP7Hm4xfk6Yh6UH6K2OCT8FT4/Pvp3yq7ETlnPF3laX
uetjgsvElyaIk/L1VYP9r0SrunyUi5HUsRh5Nrt8/FGiB9Wj33D9Eg9KcWgiKk5i
qBS3lvZf8qZNzYcAt/BBQl4HlPR+u/IGT45oA6ZYzhWm/9w9420euqK6Cu4zFzLb
UUBYEyTJxDlTZZtyqsUN/bjlzjxigqBlu77Z0vup8ie/JHfFpkQitKf2bWfGVZyv
N6iBO5g3zmf8BlEHP5KSKm0953MKINStk87Rhynr3TddHrKMm+VgEQHz/mfhKwxR
2S0u303aZukmSZB3TJXlpYAgmCOFzP6BcZoc4NpCfF7MXuYNijswWefLuON79wtv
sOZy7nk6ZjFnG0/XloTbUGBeMMtYs2iDW5EWPLXiDgmeJsdPX/nXLTj4pMI9d7rK
HUuw7vHfJFxDxdMwo+9aOKm+l3JoYMtyq4QPDwJExTQklTEXjXzbf2eDmMMjR5/R
43tQoEuMNCdXtcnAClOWpZh4sPc6Btix+zcw6UozLnBwr4Z9N1xoAJEdwEImEMEl
oRiphbuVkY95l8mYVftd8FDFkukrQC8TbuxmfUKVsXFWaa5b8NDcfD91qmQ5XKG2
7ockgMpMzG2+KO0k/k/5ZB+8jilBz0rt5mN+b19SghhW+0/0Fg5cldZdtZQh4rt9
1qvZgRO7za6fwBEnusVQIm9XbaI2lQJ9aZvb0ZHOBEElyOEI9jvXIJaBepsTEV63
JQWLoUVKMozxGmzb6kl6/GohDOwhUjYp3yaaJYPGsHLYgS4izs5aLfSczKg593wf
Bl08ueCxUfnpdoYwRCgj4SyEnpxeRsyjIK3mSTIMGaqIu5drZIX40sM3pyiRy7pi
fn5SKVSKaevGeMrVeebpc+Usc9OjGwKSVfjIT9I5F3k6qVgNij4pCZnfgVlPl66t
guId8jqnVY5nQtrwV+JbepX4m7K9iKoMYQHvxogSDlgwRh8easdVRgxC9nVxqdxe
aMey13UGd72/f18pMZduR6obWh+GCXPcl13reNIq7nyFwcuk9V+mCfwpCMQkw02A
6uU5kwbz4pTpULCGToiqbHnT+x0BtUO3+Vsq7ciUlgbFNJr2mr5G3jzXtwZmsFwt
0K3tC70QdD9ycFTzApayfDV+CIr6P8ROetm5RYfWt3IEkWNSYs8y50SIbIlCF3rn
NJPNoUVx7CcVFI97FOrCjA6wpHxreEGVCzNStUm9Bpt0iFxJtCo3n9VjZoEd6ZxG
ul08Ij7droFJfuDZHODVZmQ8sf4ZKsHalZMPcNF+9sXJeIxlBf/8wgzZa1+4X9Vq
HMsGOcYyM/FLbM/pD7UUOX2YkN5Dfoe00NGHoyWQVX6vz8buVqg7etg64BrGLVav
qdiGqDojKgLPsW3EY3RqwLBjuyJQuHsDxFP1soaVHdtIhMmk6dOPYxtIhGlkpyVV
MzCK3BX0SV6CNyBDJhuR4PnCRcxxKCgcI5oJI8taC52f4ssvop55+AW4f0MxZbro
mMXX9kk8gPXwOpWIztI4wluvNXrgSo78An5Ul3Gbb2Fz0qUmC0LfNl286uHe0F1R
i1ak5PeBCOIUo74wUv6ZEEGfC/NwhI/atnqoGGbpmPC1OO0LjHN+vCDUOP/+O5+X
kWEMzrO3w3ggohrMCKEYHZW/+lrPqGBxzRCNaZmGcMH4zntUWcrpYYBpo//VHJRC
4hHrYE40bvVJ7g2rq90WyQftViu52GyWYIHFhHlZROW3EZBKObOk5HBcR7pnpGKl
ZCb71F224d/rSCh1kFLmpNikIdZz+TIrjG0cps/SmVuQ7tPP9sAhgYACZ1q1tfAK
LvjNU7YxW6DI21y/tf1jSM6gPJ9T2lta0X3QTVd9W1OA+luznZ766fU9mzAWtFGD
2OvfswasC5rtDZpm/ag9/mBfPCEeOOsUl+qtGv31SEqhZWab5v43vV5cfq1LSF2f
cuZ9KFazgc0MOBGOEpttDZ/AlClTt5QMzPSaO4tv9BXZUT/Fm9WZCSksz2YBqwmu
Kpbh4v9OoRm58xvx1Abveegq2+NunDU1pN1lP1hJDzPsQxUcIs1GqIwukWznblsn
ahBdba2fqbEV/LfaC55GjK8CFCmfNkK3WLB8QIr46pqm4mdet9rv3Hfldbh99H3W
c8NzyKtfOl4KGCA7ha98oGiOZe7jf5BmMAhacFKeneU+JRYxjBAhOTYW8f/NklVR
VHUGQJpeWN4WWS/YZ5UDKRDuJkKDZ4FWcVmxTahmK6ocUwA7o4NzWXyJisP2d5Ja
mhnoDR1rtvcXXLcQptP7kFDJuAQPqVMQMhFqoj94PatI7NQ/DUw4fM/TyeHA0lRG
Fs04NEAfEqGpTlJBgL/wttjj9aZHEZKFbYMtBVborhWqhP/MPLxBY6ZQ3ARBO3Lc
oNmGX1hDwkGXGA2Q9to6kssDfaI0Zu4qH/L/122qTK9BLSSwah60nQnQeMzRl8Q6
0Q8+5L1QkuWZvFDZpOlIN9gZ904OkMfWnSdKpEbuG2DlidRxQOjbGvM7ScTnAzzx
ptXSvy9coVcB6lTNo18QRo2fvHOvlB/alNlh948ujw+utr51RN4QuclldvjRpmSW
eAUZkIlhWrwSfT/+MEDmJh1Dh+k5NGKRNlgu6xRMAADxKyZYQjnotqi3YjDk7wxf
XK7aemBXw4EkG9zYCs6XHzbK24VYws0svBcc+OvNcpjJvFRlJ0uUGmKIiggVBLui
CP+SzoqDJ8ixfIRu91yMsf+Gn4tX4Zh1hbH0SPA0/1sIVZyjYxOR6YqzJPJbe/uS
n3FS0QTRef6OqhMH77ZnaLNPJD0MmEHZsKfFzUQ/P3YIQZZyf2qnt0KexfI5FlWM
62o53tno/NLabZLqthrmEHJOwDGGu1XDsP600EK+/2lB46UuWzkuH1NJ0YO6rrg7
j5eqHsQYsw0yx6ADaGu2GIc1vEjVedSwv3elUY2pXLQt9fcZjaJSxet9qiFWAMnL
up9mH05vmF/9PHBei/x1wvpmLtsGNshlDnil3Cw70zB2U+rAN6wTP7e9OH89cD7q
4iPMGc+0EIJsz4ccAb4B7O/cBERPM0D66gFrPIGDMAaOSdVRN1Mw7uK2tR0vgtXB
nSk+ceRiCZoy6LaH6Mr98pWJGAgXSiFj4zzaTHHeKEwZ9FSZx1aQV1vSxa+i/Zyg
fxu652HVSvMJd+L4zXz0375q1RWE8vistT5McUG//63f1XEIeboNxTSCpM+gKhps
FRjNs5smGqXBRkY6CI7vOCkf/J8Kc5rIiAeKga059GhIjAASoKUuKJMy+SpGNqdT
Bhb6CDYk+kaJPShKdIpjB/Sk7mkVfCaitTCM3hK4rcrx8GTbCUHQcpPpY487Eoy7
0SNu6eEo/d+lcYygL9fZJdxGDc77DaBtJr7eoVur1AC19IDZo6lvUNoLXA/DGw9h
85LElpUZEIUnk0hZnED76+3hn/FkceTVzUjrwLaVusfcIaB5y5+sozkX8oFY9Q3Z
cy+9dJ7NWvwbssiiG/msuEGQv8XwxQsXZe7/7kQA8MilFrdkNCAoe9BMjQdT7oGI
wCmZruoCVUuH0Fds4wJ6a05UuaPA8dYos+d+krSNsjX+31VpaTmn7SGGR+VORuyr
TtQGZKOdxqy/2RyXAqQSn5LbAYvXkGAmRQawX+UodEzgMy3cG3Cmax0W0DrFCGK2
Fso7BOX67YVLxDKeSKFP/+ViPkttUIqH1jKGm2LacZ7x04rHriq/wduPt6tv7Snd
js0KLAImfrvKjz78tpWji9UxG04Zq95DeWrkZf5lvPBSLlhvwpP3yGgQ8rwjjIY8
j3J8MK4rVxO+Erj8uM5c0uNRaGcrD/UAv0Mf6xovnSDaQFUCx7fYHMp8OqY4cx/S
rhh7EriDdob0ITnc8jlyKM0bFk6EpBnuQIDCeFf9DAy4gk7zJ/1l6iBq0XIEtDRQ
6dbphFBtgJpg9DFDpiVDYty+NPld/KHrGJZyrZw2iLUdr7aZc8Awq2MeZq03hgm4
dx9c2NXIedFPqfd/24M/aD9PP++ga23vBi1beMIwbPZ4DW2uymiop+7mB5Hh8XPa
NlCDok0rnRM/uV5ZVMaxpbVosFt9CXciqTiBKBFYxCEN1M3DRDNDWCefQNT5qSK0
pCUaE2+GYpxUxv7UH32vjcfmwmBWY3anblE9+RG51Cf70O+4Abav6ZByyJOdB93k
q8fwV0+Xv2ui20zOJNhPYS3ASY/LM4d6emDO+usPPOF82YfA+hr+806o5vCbY/cu
jM8L0ZXSPcu9AGosjO3TaklAhPPrcY3W+KWK1ZiUqZXSGPXpU3sUAJcWG6fs+Cq3
tE2bQ4X5c0bVnOSFtSnO28n5ZTtObaOUBMLGLtGnhJEZZJ0j8115fOg3V9L7ZJwI
IeoWSPKuJ9s9f6sNM7AikYqppmgA5F+pNwCDVzn/EA/lMN5yqlhs5C8EHe0UtlfC
fn7JzrKzIu2OE9NGGVG3AEaSplCkO+QnGr935fDxWZiwlxNaN+7A08b8o06Mljlu
FxjVrVuSHYEoTHawwsm/aH4qE6FklIhPsXTmHuMsmMgt/X/0YaSzx88K/IR9IaFs
adKYH5F2PQ4lKMsoi133MzNh1qdMz+WMvPmJbVgD3ThaXyoPBQ567JJPNbOhAqOe
VpUTKtbQhKltkY93EowYj8CqymcK8oL8CDvMV8cKipIHe+JXU+5BhSXPRtUu5Es8
rpLU+emTlQgit4EAnTnRv8CtWp1dWymFgpu3fdMm9P98GZu4oOq6D97W+VnbyOnf
jqFDIZZaCD4HUzKHpt0aXbzGcN82FoofDHUMmHmllOIU7LxLSqTncTXDYZSP9Dhd
7gudqaRk1kFH02f0rQVC/ZAhIe1izG22NO+epsG04QMEui0xjbuVNO7SvipJZOr4
TcxO71F+W/JSkGQlxyKSLH269KOYr9gGpdPPYazHVIrcL7r8D2mzKprSIp8MaFWi
N3RdTg7B/YXp6nVjkgutcn1Vi3ik3+fnMvzR7ROLbwwrQUBfaDhZqMkxwVlZ9s2K
qlQ3nv2dp9pFr9b0AqlP3O0yZfMecUyxnECIpbKDf+erwnz9v+HCKkppR5GB2I8f
Q5cwX4XNQ9dVO6QDjrvDW10fDl/9DcZvMLD+a0yZA4y3+/mKMeLFThLdcYM8iv8o
FCm5/zI5mA+IlpygaB5cZbPccii/2kxNyXW7Heax07IcoNCVhSbLtMyCdA6QUHEM
VDs1jMsu5zKKbIS/pDAk1uon5Jx391H2bDEPIQe3GaDWi/kcEx+yc9LZNp/hSNuG
6CM55PCuo5io0KDHjuGydptZsSbXGq29ZtdeqLnNwwgjUT9CjFCapunemOwAyT+4
R/qbUpp/TQgdRXwyJDFVhAgzrP00SCeA5PsRnRwk9U548IHcv+4D8gUSREo1Rb7q
S1xSSwUzYZjQoj8FnSICOIHB4HR58hssgh0puL5GQ9T2gkfjwYPuMXg9q6GhnjWi
u+0qTR1gCz4WofQpkSkvQg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LwBHmqZ+ga28ZBnDUFmrEw+6aTB0rU8oDmxon+fgV7fztSjI0gNnaYu+n7RsiP8X
3LzyhnL3xDautt1YT7QquG1hh2mtW0abszswhalrujbi55NeAxBUfmwA08TIHodP
fRrQDpCDXKeXq1IMTWkw319K5em7PWXohURfCVDQ8uaOvSrec1pHsIdF78hEF23t
WSqOeqQKzpx91VUzboxO3RW9hodam9lmFe8AIHid2dg1HGqpj2oP9p9ruA7qYcps
wzOg3bUBsWH+axkeITFTG+zuSdir8Prypqr/inZbHiOELSGUDUCilre5uu0U5RMO
9Lhf4f/w83NPWgVG/i9XKw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22144 )
`pragma protect data_block
5ZBggNXj0GP0Q0JvnQPZaaMNGPFmMduiUddZ710mnHRXWfm7O3/IwFHjJcBYU6GK
EwsWuXOBk5E7W4E9AKfk+5tX5WuzQj5LfhScy6DvACpc06AqM6JAfGImyR6zVCOA
cGZLxa9exDKeQLvgIRRkb5z4SWPwAxJdXmC2ZmBqc7asEJzj6Czve9ZVfCnqCcLC
urngrPOE2/Nz20paFvCtDPdexZo48XBA3+eUNJK/LTeSG1STD0R3U6dUh2Z4YkoD
HERy8CEKEPhs3gfARP3YvLIakm8oyqRL6E7hGa4hA7EAEoZxwR4/cXb1CV0gs2GC
ibdeqBYsGINfdcPUx+MsaP/cBOhgjma164DS2M3em96zSvTdq7mmSYhoQS1BjdpP
Wm02cfqqow8bZcJVw1wWmkQKPEdzVrE3tcsjTdpE2INjVaGiKTD4M00d079C2Wq0
PEA0ccb/85l63WC/caSa5O027vTCCqMsDzxD5QhCw63QtAO3lYRuurtmKII4xCJC
NPPCznQkQth4tZsQvX/8JMNOg5Hcz36wx0knmF/phc2Ku1KPQrWdnXakaUgYmhgb
q7kNk12U11lMlbd9q4aBFfWTLbN1O+1mB7BWP8cfLxzIuCVsrctnt3mHEE3UgvIl
w4TSDYAPG7YKtLBLJ3YUScgm/zPEy0qXPUQXT+DE02f4I+kg/XkzL+J/0Nz87oc0
edS87c7JgpfWY1oyiT+vceuVkyHt1N6JFeB+rFzsblh8aADre1ZCsW0512tJYzl7
V7PKdXRUVZBKg9G8vR1HM9f5ycoISnEN6i2aq3nKY/fudtwW2pWqyrgrG+6qMLxQ
ph8D8IoXGfB1XH+6IBPoM6jS3d6Pqa6VeOlLPOS4HkSi5e2SXP1AHB17cr5VjmXZ
Hb0lomvawI10oSgYqFhO2A+mscJJ5A/T8I153WqeHMVcakCZbmh3KJnv8wfiZupo
8JlZEcIlCJn1XA2oFSNKXjq2aNwDhXkrUpTa22+xvlNx1QsDDfqqoGG/pV8mrPrX
I2rj2eP1GctzvvpYWN4Yo78di00Wzo0hyVKgGg+FrX0Q3H5AfvwA2lB2TcX7/xvz
hfeHdI14RtCR0nhrsCcNrK2QUBA6XSPQhS7UI81qpMmW9TDChN3TiLeKYydS8Cve
deQZASb80VCuZ6QURSVBCSIE4pYrucfUkH10m/0WbebMZ+pGT9sTuS5apLopChez
2ezW1aI1ek98E4/KJMZWa36EiuR1VgFqIYd4sKTUNpL3crf0w/gJ482UMEm86Ds7
i7uU1SQa/4fvRYtXYhChOheVNI58/TsmT2UEQYFqoVPq8HZMFVohbnejkZSI6Ywx
VxyVRYVTp5LD/qfcdmTsege17qOchAUBbIJtClV/cLTzWS/NCXF6ORn2FO5OZfWZ
cv5axPVBnNn1l67sDUceLmVloF2vcS80yItrThDup9uvq2r0WwSHP8pG1+oo/dVO
wCF8hqGjFRLiHg9gZJ2PLqPSqE5K5f4kVUYPo5gGLgBab/e/8GTSOqGdPWTA/s+h
8vSedbNTwciCgbCP3dso2kRwXlArnx4YoSojOJ5BLxMwf5O8Uvn9WOtVDU9sXcPn
m83nQwhy5c13dca9jLpPxBiTaS2HbuWBbObW1SeXQcgYtnZq7FK5/aSj7pgwT5UZ
NrwIxws12xBAJVEfVeEhBLE9dW9sKxlbMhVG/rN1VcUmZ9QLOK4GJ3GZ8d9HLGc+
Rks2JmNZ6nS5SwcJGRyykJtfo/U6A+QffPN+Z5QD9/mH+D/eOjop4tWTfghrnxvt
H8LHdcKV+QNJAqYUT83fYDFs73QVCa07Jw1ymjku8szkSpmhaBA5hGywoQQwfeE2
z1rRZhCaOFPpnx7GAKsOqGKKQXerlv4U+RRRPjo322mtoSMrVwvsbsfrjWRXY73Y
AHlA7xRWwAy2qpPcBc953ujuVGR72xJQOjT35g1H7aR9RwindsmkWDMN/AQ9DxGt
EiWCaXOYeO1PyAQcXzBkwUQa/U7VIaXsBYR4p8VbKRKN539kRqfxadkHFZNZjL21
HsiErxRbIUALjEteDoQ8ZIe0ywW2xL9LnvsbjO6Xs8m6CyrYxubWHbnmR2Fw4K4s
7lC/XZbyvAGoSL9XJGixffNo0aw+8xAwwcodrZfiL+s9Ui6H0gZe1Dk8p3H883Qh
krdl6FlP4KNpsisIGJ2KIU9nMfIMb1UzdqtvP8FJs1uSYPZlgxEKvViZuXN+5kMh
feE07FBAKE56pRYwQztDDeDRm7S/gMA+9Gt9fj+KCUZbyrky6trdCh1xPYdCeroR
/07J+q8oq8MwM2pnqmSlt2aND/f29CCG0+pq1vUuDE8U3JxzxN+OxCE9GK4M9H/r
Xb0GNroJZdIgN4fa4uBc5siOgLjk5D6M/DiBPm+nREiqTip2FWANs3CuY50fOQQP
Ao31safD2oysiNcITC9a0Ppcmdv/af8K382IOh82OOy5N1Q12JHdiDkg0/NeqgQ4
5p9m4Et7X8FWcr5Xk3VQVw8yR0ajjM5vABNe5/O5bNRdftdkhLreK9ZuU8TFJ5u6
d5m76ur9QwrlEEYsvq3hf04Dn4SWIFGay3j+rMoH0ooQovoiHcquIDa1veT1dOw8
1TNNbJTn43im8w1wS+s9S+HraY8q/9j5zcH8sSsBYE9uJ35QPpa/tbCdzFoO14j7
UDv9Eh2wzghodrRfLFJclOpKQvcgFbgpe1ltesReNKpNPjaseprmenDiA+didnXh
rDr/SCIgru7czEUzLm66kVDqvqwRNO+0dqnFCiC/vSDeqo/ya7uxdnFLeR9tomHV
ugc6+bcKt1q0hXgz8zMZLu7chZnWDtizUaOZulKEYUwW+CVJKoLWUfTD30Rkj24Q
bp1yvpyVj6NcF1WctDWu1uhCMbtaEFcoexfKBlVMiLXYzH6ix96NQMP5dHtTAojW
asprHp2ZLI4iVrcqk08QX3EajZ7hqCkN5rt70C5pbWzS7pWdYb4aFf/8LkpUBFGw
tdfEGL8ZJATEO9QxBIK+xVWpCLUyR0JlQc/YSaNN5B6YAfeve/5GoOjYdk3uPomu
t+72Yhj7Cn8FT7fQXIvGiLgmkImvS+kCePfGBNwlcA3w55xAUFJDjH2m748Z8bjE
oaLMdr70gbvR0QjtdV38BDx+Oa1xIb6V+zir4R5D7YGJNIo8H2ilUqYKms56sFQL
fSBVyK6jL1Qhj0NbMQJJ3WGfEXuLchAZG3ZxmuuYJvf1OQ2XJjUrrruA7/IdCRG+
B2EayQqZLCSqcjyWBfoJ4Zd7FTroEKS0CkYtOMkkKDeKrXraL7DOzDY4x/Eq1Chz
HEVtpcS/XhWrCYcO4WPVp48czVZbS2D14MkOMqxhr7usOWfMQCF92YmSVBz5WqGQ
t2QkzunS2uye0YuEE61uMoR7ZYf6+AHTZqArFptEoFol0SC8Aw7zeJx9zoKyo27R
3H7ljKyoaAAc7GGQah8YAh72ep9qo2tecjWPIqFC1/rVRsChkCOKiqLsDZqoAsHk
cHhxFwLPtbeI1fgiu2EEvuCJ5wfLsqgQ8ah3UeocuicJ6kd0+5BlnZCEnn5aDSod
aZEDrIM7dzMOJjRRrHIg6tfjO9KyfSI2X/GPfCFmzlfhb6PP00DYy2w6poUix32Q
tZ8rQrtbyqeHq8zRq/Y2oT+lNDKOOYkXqwoGW0gL3J0nEWi6OWm2ATh2fgIsrgyA
F7/nD4jmbK4kcI1RBfYC9SZmo5hbJjZa77hsLOnz5rD7YQo//fPojiiZl3L6bP3z
LNqC2bEtpr+yTiJOhUaOU+WMRWo5Mj9hoby1LSqdpiPuiZs9HxD4RG7lIzMrRX4l
6y1OeAcK21TA8CSirQ8Wr70v9OdKlcj/OzEdZmhy/kjhPVJjLL955jfYK557sI6d
vVKZs0SDQM9mYbz/DAowJ5vJoXIpbU2x1lpPhpIgS0aS+tmnusyIBBu8K/6aX8xE
hVWG6XN9PaDtntuw1pmoy8YGNbehbEXVc18NtMJUOgsO6IY0XvPMgHvTK+MIqcA3
UGg+4QdcnCRJh2mp5plQtcEbvzKgwJNEQrpafMbmMMctznm5z4/3Vo4b+ww66LEk
4itFyLD5b9lU0Dgt/S/8I93NOfa0niK45VwNbMf2nvxL54B+IBbvxlVC9642u8z7
qdad4NtzZvzAEGee2Ky3QnATcHQY+UudXpm7/nALMGuaB/BO0XejlZWtZJQM2W4V
Z2Xqk5mwYSnGB9dQ2Vj1HnKM+bbMn5FIRnBV9TPLy3myPXf/we226PGTqtU00jMb
/h4pre0GreDQkGRLQ7MXax9s60xlLyf3YSdocJKmKCJxC5PEEPzYSbnyekxS/Ngq
mHAqYByzaA8Qf7hFz6pgcxVsurtc8tbt4qmEr9jwqHSLWJEMQSNcbZ6E0seQO1rE
s+kXkqd7yy4rrxqOVzEoEsgwU/tTVJIBPjbgzkeprHvCYzogPYov5yEcVYdJ/nr1
S1H7gOQCqCwbsM2dS2I+9O9nWQAjKHBYkyhwZ3qsPjGspFx/3Z3tGbILwsjJDcm0
vvBaPQUINJGH+BHzgA03yDKnP84xtCQ0LzTP9RoA9VmLAo2oKCyBy/Gp4Cp38dVR
0Oh06UrLKrGK3hG0VHrM1JzE53ul0fnTE4UU3SLhwMoOdScAhmTgva5L9mrRXkmO
TAjL2SarDekisO9K/+ZKqgLpYl4eLe1BNGlJrz4RTtpGzZXqXzrfK8kKGjmX5uUu
8ce59h4pmnZ0L8wI4AV8qnkbdM/ycHpzwSzFz2FaFYPB4bzU4EOqd9Oyj/kmXtD9
OXx0vens/Nrv7s4gJlot+ehyCpLEbB8YxYqobgA+ZDz8AQXRtQBwxOnF9mzCX15B
wUFWg5EvhIcKBKPzkyjpQRy8GCzFsxKY3hoR3jr98ntPOBmchUDSXO4FuzxzMU2B
XTV9Po4J9AS+2NT1S1TRwLOoEEDchAV6W5BiAibJLvs5UrqnuN8nDf7NLMe/hjXq
+s4pT2z/yl3DJD7czdlDGChAPMUemXepUh6OonnexN4uc23ZBAUqGJ/lyNXWDYnK
Vfe2IrOzO83Fng5o0UwM0NdW4VmSBW/y9R0xeNZ+gAe+UM+G7Gqfcs4fB/vrw58x
LWIwdEMoGYJCABD5lLBdZEzON/wP7eEpMM+JxwFPZykO0ycyyjLV6O6Ba96cDjN+
W8PSGPud25u5N03FkKggtzinhexiPxvtjpan1OPbrFRr4n94Xz1s5IuuXfLHy+SR
5xNWSjptBj8LcUffjeLKIVI2l9wJHo0VOgHEcYTer3SqknbCQfsxrwSUAhwW8EAG
6dMIGtZPeV9DeYrDSevwF6cqykxsUc+PDZkJTwXJlWCByv1giWxKEKL2HiH8siA2
XKlH7ts60eVw9nWlyIuYF0k6P4SrW7kbUmNzrwqV9hmE9tOs179bNQCQjHBtMjnq
rV1m8D5nDGO+TlIK+ZOToPrOKKCoB/oB9ku3v2V5cBb5ypt0y5dglc/kYCeud8IV
ZA1SeFTYI0MZA+iOCmMMVKqwgzjmYURuL4bO0YUpVoSevu2c6aX74/gJYMPBplbA
d+vKEiuIDYBrmh9yUoVYmSheuT5PIkgaGnZ0NzPd22iOn9AJuuFyiosnxSS8qSOV
jeMYEzqjzY/WLcr3K2aFQoNZKpSb7mWf8RSzs5LPdhAjUA569/cm8YUgHC8UkZEc
/8EaPXTBkqkE660Owc/R4t0H/tuoOmY8BERhNvSuuKyPWKbolHXENCyaNasj4UV3
Qk/g1aZhMT9LMASDo+gOxlmgNZeWudVkS7ut4H8aPcw09HvFHGunTlamHqoOZFJH
96dShejKD+Jc8fDPG1UUzaSXpRwnXO4aiRtftngJ2drPKahv0/Ykp+9xDptWA7Oc
VZn7FexoeaGu3DTiAgzxSfvQCGTsyT8kFirXCz4d/1ZNmqesB2s/lK6M+ypvfXt2
YwnfGfCcHgnT6EW2WUIDgIhP6QykyIjqWM5ZpO9PD+CigsJliUkPyR96UF+Rnnip
//yHvURTR07FYHs39PeNqFW7zK+U80y6fUsDUK0XrHwOleQ4wpN0PYZROomOKC1u
vZYOGztCiTXGngKpMlHjxj+gyk2ftV+k1Pzb0r1uIhm0yS4gFSSPkJYRNPFX4+YH
58M9RILoGbPsaeaaVQHE+WdYKz1lkHoWuUjhtgbMrWE7qLuLfy3Y7PVZ6Vn8mFjt
GcK7JDUSpSdq1OoOIgtbqZ6ixO2dc6qNaAqaOx+qWy/Wv3O8d+F8NERe5vmy+tbF
H/jsEB4qtNjiuWC6PRaHT9OKOxDVbOirpMTovlZvn46pH6jvcmtgtmQjNaGU2BEq
DwC76XcmPtNXc3C1LgEQcIJSC4R6vXQLKqHXw07ovlWfRl6nPZ7JNQJFLKo3L7On
zppykdLchmHhdHfWABAOfsiwGcGuFMs0gwSdJ/oFhX2go10LkjeLnF68bo+iWPI2
Ic/SVfNsROm8lymYfT/K0t5xZIo0oeNw5/lUQ6432Okn68FOTvcBIxDkytilg1sP
JTT8L1gLGHcA6H9Ho/LaqkqYOuHls5cNB/XmnnOC6A9vHLLreODACinzmpsYkgSY
oHoe8WAiaxx21G9/URIJjbrhFmbuQDuxDuMxIoYFfXvqHtfdpQXcCScF5GocxSBf
zhT0C1eMT8YTl2BR6E3y8iFhQjT+LKGAU1V07vrckC71DCz+JnYMKCOEpE0pcnoM
EdbDSLz8nxXW3XvOp8QwAaXlc4UBAJ6wTfYR0HMPgo56MLSqWrdpoq7xV1lUyGiU
mzeb0+K4gRcaYy9yNJZRXdetQRRMJHnt5yzghwBBqdlB3si/eHDRKJVfiQ3/McPP
xD1mYO3cbz1c0xQ2umJFqBUHFYNgZOSWaoMjiOUNGP3Q69sD9zsm/c10d0lfNMpT
q5MhNNRvIgU1bmnh4G6aBWe6fI5IqrReKG2fEgT5fANdfqE+D8zZGJiUHv7Hy164
aNrs87ATeiRF+THeahCYllMRDP+HZMRNkNLshVv5yhxGhUfIGs9geu6j0GyqWsFk
IW2+q2DBEOQzOd1z0o33pI1sDSxv13BldSk/DmIS0HRUPYYFSgp6rE1VXR03turq
aM6gt4s60hpzNXnxyqBJLeaeKKUG2/SG53GeWPUuz8U8qaxSeLkfLn3J/TZY0mJE
97IJ4WJufAC76o4t4YOSZXxaOhFSCdLmG6zZj87Z7+hh3ito0I0nkSx4+BDIwyYW
twNaXO+/hJl3I9Z0RO5LNILympB9wcd7IrTc8kg/afhsLf+IH+z9BR2Pu7yoMI8/
AlCqA4qffk+jSuCEjG8TABke9hgN++zVxPs/HYADoG85w4Z5p5sEqIMvA/QHR06q
OAeZOaJxqk998T6OU4uiwBHaZNK1JQhddtcqFRwrAq1CB7JneEbYr8CFt42Wph0A
PCmW5uiK/Hw0HlcmNlNzYh3g/dNTnEXN2nWc/lXwZOwsPZdt4kDKk7y1E0+GNpVm
Dxwcz65wIzXgGvOyvxsRk8onUiOXIlbGAaFFUhkLZL8R8eBKN+N12HhlMZMCQW/r
X2OVE98WDZTkqA2ooFT9MhUHdo4/zKoEBfi4B3nM1Zjf3Iq4DoR4WYZ+Al47PY1l
1fFGQWAGX0Ih40CxmJyDIeM2s4XUxsYNPViFc7sSVF6AZJBAC7iMe4Ii/DVlwpmE
lm7IiQGv5jf64zDXF4CINxNzrE9MpFiURIKaOaxUH74ZypgEZwWDuwfCznCdsTQv
9KxMcnl07EkAUbv8Gm4tI24k/jsFIOe5gcP3L7n72VSdk0pPwDoVX/onhEQXqX6Y
QK1xDVfshRVU43bjF5poVqwvyr0HTLYwkUK7nsNi2PO/idG7mty3yfQvXKm8+zzP
pnDaIo42LolUglg+Nsff1MlbKaQ6dOycXwx20vD4UcG8RY+ZIWGsfATrJzG5DJDt
8GJ/wltjyAyGdYEqqySRLbHs+yKDG2WOGoEm1FO1aWgraXRahPi61llNCRADxSuB
vfdi/NZeQusHhOiCIimyvALnWyvD8VoALfXywC8rRUDGDy7GeVuJyaa4WrOOr/pR
yb0WaiO/eTBgZc69oN7Hc83Wf/L7j8H1fjN+BrZum+vP9fWm8NdVjz3plI9mwHz5
ue/KdFEbg9AGnl7rfbeqhAX5zqzTqMIMth7qxU4ej1wHPn1ihSxxXNoHsswVIvYx
2Nq3+3TpRitzYlX/tbqm2ihyfC1LJuH/xO+WYVavrlcY58PHEODU+6MhS9VVE3np
78VCJhETf8enezxRhU4mxc0UQ6hnR5hQQJHGR+mBTh81dv5q3DSF1/n3+UGEWaoe
KQBj6fH+JP+B4gEWFQCLeHhe9pK6zG7zuJvEUb0i+07VaBDHPa54hNq6/SgzM+ge
Agd/Dizbwa4HGJ+jX+O/k2vkLn/Xpoh7IV7DA9N7r8gEAGJXr+vITatZmTcvuYeg
f4LxBpV6gE8zwcRtrns0yrwGPHZKWRq/oYNqRSJxsevb5kdS0ZkQUicjMSGE1CL2
j0PyWh1X/YVHKm96SGf4bVuCIyiCM+VxoHbNWAQ4j9SoM/evoXFg0RF4MdItha5m
AUv73yCDpjNifhq43YbvSQI4lolN73r6fSSv3wmY53tAA2sWQpTQp7DLMHvBKf9A
EP5poDWv8Dw4tOgUaDA7g6E2R7zQ6H3KYLmNIiNh0znEYY8ZF9Xr5Zuw4IbZYVi1
qko6HUBtdMmeGJ+7WIZ7Ubwx0TS0Cn0O25UPQDQm8i6vavm0DiG5u0GZogCxJRUi
P/0RIjcsVO7gAFLhEoBeh6PHfILGtgtudgZnxGJvECv8xpjMQgnRcj2YtXZKm5SH
Tujb4NdttaQt5TWcNApQFQOZX6wMu6HbwUdNpg4qIogEcnUgvKfHmvU9/ilnZFgr
PXr5yJ18jExsRAAUzWmwSCvUN/JzD781bgMd7QvF86ebS5kezn4EKb0mCI8BKcdH
X8z7h9ZR+7ih+X7vU/ogBXpMImAFSAniLRr62jTmAZRSm5rqAsUb1uc6OEbfuLhm
5jlJevCryDbQVKY2s2905DfCPwB9hgE1uOd1557sF+q4V/s2oqorQ+8ltlzvGP5s
X7gCg5RvzOn8yMbsM83QehOrAl2tNn1vDpE165cq5QGwAIn+l7UpOT6x22shS16c
EpWLliXSiG0HzGAf8f6YQz3T23t0EEtb8onhYMCbc0n6olVCe1r+ULjpkRQIaPC3
ttNltQKmAMNGjFlGWhYOHKaLQzCEjTl+QuxMUNBkb65QbnoZhPrmgXa9j9BoeNSr
/t10lRvgyG93WIdqF1v+9t/te2kCSXZqi62vd1Zk57eid/gMDCJw/URx6qCIOHqx
L/monbTeIGmZlwyDmRHfwA0EpCci/77DpJqBiaFS4a321U4s1Fvw6LlNaoCm57qS
8CpnQ43PK8GhSZMk/Hb8dJw1v9YiCFCIltp2GYtSHpT893txqqi/ldm/IzsoRNkY
131M8oUklPwdNwhS2HjKVGkxaq9Is4Z3a/zmBPBX1DdGsSbxv8R/7uVnKfYXLY5d
eUqEEBKb78jHyISR1YhrhBuS8zsonsqsTsuP6EumGbOFwhxqh1aHgv/wQYPIEBmm
phC/sHXimnRKS5zobjrK2Gw4I0kK7OczyKMKrz/5whNRmbW60kIVcgeHmhBMSC2U
K4FecIn2tDE79Rm2NzVmBe/hlPHl3bwEyFtteFVG9VPmc3ytNyntzY9H37vWCMzm
gOURk/CZbCCFlvXg9zw0gwFNSKFHfnhUdOP7b0BDivEMvHT31HeKP2vV5bt1Rmwq
2ZXJpRLp/NTXUesQC8/dycIqabvGnhQLdO3qBhG3GHA2tcCW5X5u3Gafkg9kgXju
ZIG1crrfn8HjBXn+Wa3KFxlhChYYSv+/FZkRX835f/9RWzuDqC2Ue4U0S2nkqUBc
AcP1qMcX/9hxQ7LAFXiMWB0yKrWy799nALWToLpRQCMwOhHfhK6FMyEle9PqrYd/
OQ+nNHvu+cX5VUwIPiHf84wYkGtoISn+QUxO0Moxx/gpX1M8l1p1KELLFb/+Pgqm
waQywrGM9o9Xl5g9mdzKWEabgzKpJC4N2BmJlKvBtZYSR7fMgEOH1dng5GNES+kp
ERxNXcV4rLZ/hC0rYeyVnjYoIU0tM5sZy+NmhHbXnwvx4ESAqIFZNBbRbZAU69f/
m9O7INesNe/UxiNqDrRxq2G+WlYSSiDmCPOqs82ntFxXJv200EI+vNi3sWOl6pRm
uQ4fS4OJHypwlua1airll2E4RPO2PW3DOR5uhY19mrH4/iHngR0vBteOTpju62h7
Ym4+QnVTz/uBAHeShT7HfNrCplIfXnB0Mivq6jP1HGqd5+37vBasnMCYc0ZV3wOb
/PTwAhYbcyucMtLlJLwDBuHU1rJWQQPYHqUdQDIJrQd1EL4W335boudIO730bTl4
kEXrNKseGRtC6ZiUVzotS/8/PAkK8bkUJDUXBzJvyThKBBofPnTT7dMk8Kg50+iC
LJiCR2YUHacb8wpVFsPBf7ocr/WLWZrkIzue5sOPjrq/sZEdbzykOqJMwXIdMemQ
w5H6AMfjjBpavTbNIS7DJ593J7xG7cQkzwwTX5C1HINCK2mBnVd3lsBvZKiH9I8y
g2aNwpqv7XMdkX7Dyj34IUc4ekINbQgYDIDlGLVfwXXRZkxzajiv9KHQHor3ZuEg
scVZKvW9EyeVJGWxt2NEqhLj4C2H0Z09eUSN/RFRuQ/eKwx56DqDX29kSqOjDp+M
A/rkKnH1I7/nZec1BUTShh6IVIU8z/4iJ1xS0uP8hyz9EVperj97MWgjIW0Mnsp1
2RtUjLOFQHYi+CCtRimwcem4iohxZnoA4GFeuki2P8P0nI4VQU+8pKs2hw+C+rtM
zQHY/c4Ul9ZIRYydnE92jw9tKljWP5tbmH2uhgnbmIUir6PUY+w0MQb3e6R8WtS5
6YzP4A/g4EjUY1Lp3+Nx2H5BrMcF47kkvvLmqxV7ztWjV6sj8kFwUYL3twZIvKAy
yvQylPQfk5NTz+EAm9Z1M/clQxd+tyrv9eD18tlkVtjkZhMPH80ZgunlWiYkb3uc
16Ea0mSXyS/pP+3BlZ35Szg1SUv+4JcwNJSW0UzV/CWHq1zwb2MBeRpyJdI6bFon
HgwOc0NldHr8HXU5JIbL6CIP/a61JgYbLLm0y7C6VbJFFwL3teRZERfA7YlZCOCQ
0NDP0tudauO9Vmqu2YVCtp2XWZNDhiK82FMH2vtEyux0rm+GihymoQBSk/3PXFxR
lqKO9iXTUOxGsvdWNmuzTUkBxO1gmZAxNDKdYfkDOi/tXCLFz/4JU6746m16DNbM
tjX+kKNCTUA6ICiYQQiHsEG3N1hab6WTqO5r2zagm0LY3kxcipvDDivKpu7ceY14
VT5OaUX7kfRfPbuX44JxSTPWi9fpNJIl/J4ju6oTWxc3E8Ivl4opmM0Fdwwk8vSG
3JFdtdXpBbmOAUznURHK9tdDZgJVwr3gjtKiCxXOP/5bWvbukYvHrjLe7cSS8KpY
vMaPJGDq4nPgMa8Jph/wwYrVXQJxYwEVmLs3sF7lQbJQh5VEU3zeeyrCWxrFyC9A
G0QpgXa/RpVHOyalgjpSDHI/lmTc8pP8DzMMTzV7IG97XBN2GWoSyqCtNeQaJMI1
V2upZH/KCBCCaowe+45CiMUWY3C5eRvwq/RcLBZvzibP9KNzfU4KkRaQU+BWCM5K
i5kFTgP7we6SYv6fFDvy64Glqmmij+Dha4C/RKoPPDmEP2wcsjoFXdd+6O57gzjg
0EUf2oJP5yEqfMy7+61RaUngPnKhDYaZ7OX9GhSNrpA8FB9y2M6EnTkAkfD5U3z9
jS21av3731BBH+1n/SyM4p1h3R/ANBcIj6SsvYaMI9oUGlO6MV5qF4otGeDQe3t2
Ql1Q9Dv2I3tb4F7j5PeT3iO6BeCDRED3v/q7kXiKle1CCddiE6jhkPSmDfdvjSjo
T62TCL0y0q8797V3BodAhVb6dchPJDrvgWzvOwsCgsDQyd/7Qt7Rq0q3MBsS6XCq
wzH1pqKYICWOKWMClTNUS9ZQkgid8KH76VO49WbZalhMW9YlQS5DoGMt0lad9b2v
2mlNixrAx3ZHI9t91x1iZFdwXEV57eeXCwEpuARAkx58fcPp/dohAK8zYQZs4k+k
WsuE79fV6d6NlKuX/AEV9MBIk0bvxeAzwARWkV6P1gVQ7PNgBwfcEtYyMyAxdvV6
KwXSUvvAEoqDK4+Ceg5f3moUL+kdrv6bMNh5RxtVLGVFK8sc3NvAmO2k2YNQu2vj
8zj6TsLCz56WCr3LmTosJUWdyWIahgU3TH/CGBHTqcDiE3aLuxtUHpr/Ny0bw2Nc
RtCFy17Lzv/pt6nGxm/sV+UbvcWWnY9mKXJENT+BqKJXOu9Lsa78BXL3FiBG1Vxb
fjQYxnmr7B+yCdOoYQRBxH91w/WzOFTxjI6831ZSiRiBkTDTvhzzgwX+wEOelixU
6DGuz/Cq33jzg3yjdWvI+lxdVaBx/pn7ahIha7WU07/aSO/Pz/pvmecTqOhCac0v
mlKUa+nk3BpCPMyxe38PILmjUASkK87xUOIQYVku92DD+QmJeMvPoapcWYv5CfLN
rk3RQWfRTTWExw6jlM7zgYXT9Q8iY5Q3O7YYVe0i8F96HG/oGX4PtK84AbbE+5nj
gOvVAlFwYxuFTp9umHd45Luvg+0Zi0yDvzW7vrvRP1yayENWV+ngZnql/HwQrKNw
GD+FyM73Pz4gJg0jWI24s7ccJcCuTsFw6Qeik/BttZVN8VUjID9Tk6IRqy5U0XdA
xR2RvPWbnMbYZ7LsAKXyN38Tcxm/QCqsO4nssylkj7uYjn/1WfqVvm06qUZdFMVk
epr0zBTuZeDaqfG7AQ03XZbr/wrGeObYsUfh0T4kSJIXFZlUGqkoBO/BceP8Kw7F
D8mtFeKZpNu3q+y0tZVcUk5wWMZeJo9LfkgqtaZiDhL3z6Fygz1w9/S0aen8KU+y
vmm5lBzRW49gc5U5CfQ8xPaxPEeVEJxOHXPzt0DBM0Zf1rVgrGX2p0lAKUu7cbxf
rGURMYrioAsr0t65WOvA69sdCsfA0fmdCd8ujVQpYhT6wvGlm1t7jdgtIfPfUMBo
nFzDzYdod2QmjCjeLJZ9M1jucgtKxxGcg4nXszKP5WL2wiSadh9nLewmm1oNSmbc
WZFpHY6FTS4MwLyWngM9yVR7RPzum+7jl5W+OWjVGpcOfylOFZroeAuOYQH1G68k
TwSdyUVAYWoSsY3YZ0QQEFmgSKFUUxC38Kgpkr7k6UBWy2+6zDbzBHGKMOhmlX21
BARYjqMsIjbMk7j1q/MS8ngGWzDvXNdKE1vKH7mHyrBlCKLEatmkq72TR4B1q7kd
7wOeAAv5gDhraDAUpqcwSXb91GFWLyVJMsNu7v8HQcWz56roe85+6osMjQYmtpsC
0sv3C89B7ijsH2mwmy+EnH32lMEOV6aK44mIHsc6a/NzwpW1n5K4EO8LiEiI33+0
06jrAgaOOfkFJrPTquAKh5FbsUh7HS73VrSAViSVrm0i0RS8ay1KguX77ZROELLz
a9RC9kypq2/4sqHGQBNXaEwc0coGj/UwoUH0o2ORDozydqiBBQ+nVDMQZzjtkSHd
ER3M9V5S9dzIyrzkAoLqmgXSVnRcfgiW4tyVboiRwCMCiR0wQmDWNF+l/SApuEGM
KVmVWBxTz05liW5zZSNM9q90LUdBA2jg/ZamLf+fZE25akH6RNDL/ELrTVGa+gyf
wogSI3s4T+7X6O6g2uGUTbcyMZjwdlqTS6bkaEBZ7ixoAC1smIgAsemfr/KHSy2n
sG+xL6Fs8M6pc8t3ixnIV2UZDVFrXR/QGfurJjc/MDZwKCwfHNbvDJFFg4KUntWB
l7Tf3PmsUWJ7HkfYdCf3EDN1W3tN1PFqmy94vp0nOpIr4R0HCcJkNNiK4ku2U2Kd
v605kT4HnKA9PocvytV6Vbk9SYypDDgvORISRoY/zBbwyrRYKbS/jByAQ7hI+0sM
Khd6yr1rBqUmcZqbZfU4lz0+H2ISmtMwf9vDHdNnemcJNxAFYxSS0PbNt3kzgbB6
oo8jVQmF8deuSgs6QqNLjILzU+51pqb0KpSoeb/hsWDJD+KH+7huBI/wilArUebn
NmA5ulgRaZOEhISj62CsT3mwby3UloIg5NXlT5YpoMcyjPyOeOdG0a5Wm+LFHYNB
Mudnk0xB4hOqq1+RLGjYJE8M3jqyh2yHmr3WRBSjIUrfyFlKqDouORezcXwUKTQo
iS63HO78lQnoO5pG0sK6ikCRcI7bAFU7axHlkI8CV3/c2wUJqz+gaG3BaTk7zVI0
X9frrsrgfGQs2B4gKbtCowUnnOdWwVMbtkJ/EeBeRCVgUvrnU/HlugU5hovBECZJ
dGpoZid57c6SzP+4HjVs/KmB5VYRJ0Zr8ohaRF6GXgcj0zx5sBJF50NimZEc7UtY
wilOF/x6B9W/0CDvSXpXQxYLicGyiNpsz44+EkKfc+GShXOVDQMsxGLwiwViKNwz
V/U+PD2vVqVBzornLOi7Vchpn0BAb5a79eNMm6gzQiT+Ljx1ELdST1mQg8F/Pw+v
jh3sg9RAlqAAHa6z5PNJQJr7nDvqRdVOdN+SwnZeCUzt1A0iiQh1wf4BDLdOZxwt
foeEmKQorCX8ujnUpHvB+Ko8MgBm50VKhBrsPSs9zNJKWsCw+4xLQ5FCxgGRWwVd
yfL5OF6AzHae5GmahBurv3QeTCB3WXzQpqCUhd7336U3duY0yLJN8Sk59XD5kEsa
nJN6/jgGxf61La8+m1ENFOjjxG1lRdKe3h5kWBRw2Ot8m/x7Y2DjziXtnLhd8zjq
elaM1dQ8031CRdM5UzsoZOw1hwtOcdYFmIQSW+2LWA039DTxIwvekcFVX6AkwJhx
TQbuwK/qYa4Vx9u/tNWqhtjVBrMI1Ifze+R6bnT/Gjz92tsdKepePywYVB4ua3RI
z6a1nht8fk7dXkg0ibCbdCU3joqSnqgLrg6F7uP2Gy9VzqywYUHWEJm3yTiLTEQX
g3dlNtf0WPlnOFAhsqRafwxw38rc7sTG8LlBXhv7zLeEOz6xiwUutvKOwR5KfXC9
TXB0TX5ET6KMyXlbt7cvZ5yKmrOL6ZuGOl+rxQu+PCc63vGnF17td8pkoYuZxg/S
jLIpwFczWncpp6EX2rBt0KX5AoY5loYhIuUZG4Xna8Aup6msn5gzaS68ydOslgMX
0lRyWFTOXUVpgYg9+Ic6I5XhzAX4Q+qIOBUlCiA8Txxc3eTsqKenEHx+YzXefyii
dzidsNmrqAtEz1bgZ0WL2KrQIMHoUCf3NLZhuFg5GhDxvxRYGt8d/28LjaCx7+sW
TlpiiryCaDCj2OfXYp1n48Uldupj+xbl5tedsfIqISnxUotjokG3l9Gunj7Zcx00
Oqi2Os8hnQbWPfsY8hv8qEfx7dFmzdCj+PPWS4bD3o9NASWZlT7amzrqYF/ik+ID
M/xhMPYTand/5MmmZ66rih5X0Vk8RDLc328vg8Jn9CP7qV63C7D4Gc1hMxCdEyza
jS+oEqSur6fdD62ZuJwxHyjb0E9kNgMW5U6hDIMhi58n/JPI5F6A3U7+77xK+QGT
kUgmW94F6JGTJenfOx2ribIa6TrqTiI+7WlQb+DjnFz217+qZ/tEO69PHl+ETf59
NDqDqHZJGdngLhh0P026fOKP3fCCGsnQJ956gYmR1+FZ1O8WUxc8HqIwjgLlMM2w
eTAVDqa4TxM592ITaTwNYhYvCXnjVAHHbB8qmU0grB+NP0tRROYODqH+jltcC1S7
TySi0vPGf2NjISXzLRkhAYTNbf9TlFBQWVoADJdgsI4PI4L8cmR5j9pRdZbH1Boz
jWaxZoszh1Kj3kpz1mLrYkzL2DEH3v+UUjdlju7fATFhh5y9pcxCMvN/6lCJxnot
RUNEZ/vOJTr4X9U9nhyrqkr+Ee9nmeS0zI/GbucE1NfuJsXCHpCiOntG0pg6+r7T
sMT3cKUPco59MXOCF1wr7SIYW/7H8Yl6xrNYGV0sQdPtphF+5baZ1oju7QzhT5kN
kQCZZEQXQgC6rgrvPqlhFgBZZM5+Mtw8m9XCpAFywal7q9HWVrp4ULJcaBa+QD9d
/8ntrLDqqHNbGYZaP3FhlK3Z3YVPTKYz20CAaIXt7n/rHo1kb3RidBYetvS9mg57
c2VeplDx0KRod1Ul6/IPFvDad1U987h/tmAwfsS19grPRIeHzyq9skYVEY3SxDpE
UfHG2K3ZuFfhlBDUEHr+b2kZDTXKBnpDuzKHzwgXi33Vz8DikVqr+xGfEhmTZG8d
dzz+HR6UMts9IHbElgvzGsJkWGj7zD1LPttzT43mcXdw7144YhmaYL1J5/TgAKOi
d/cOUYPsAqIUuyQlwJR+BFlxMXGWS52XmG9aH8f0BCC5hmVA+mcPAQQ3K38a1/yp
xGoluqhlqPZp4rHd6zg2/LH9M/7sI+BRFgWwB2WkoUHmjGGLGb7eOzt4TefT9ySr
pq3mX/UTbKDtYrY3jQnWQ7F2WxbP7MN4FPYa62+cNSV3qu5UIWOb+Zfhkm3Klsh0
SaGgmgckRSxpQeO15H4OsqKY1zhpbxEhx50uLAA3GgeFiJvjzngn1frzv0yVqWXY
hM8RAJW+YhXyvurbB2FEwZ8odgTgGElZJVTFu526bWgPDWlVSS3hySvdJK1vj6nF
RxX3NEU+s/hoY4TITqBNtqZogICLC+s2m28v+E2ZcDaQuYRgD9Ox7E1xtPBm4R2/
ZsIoYF09eIRATeZtK+IvhS1+kdD/Oh8jNryHjqVZNvYBiG5u0K+Q13e3AW/Llnkf
UWVCkLr3Visr525jERpWE77wHUMUmRQVjI4hvgTkigEC8Q6nxbiu1O7MtxXiFRN7
8cQbYDSRhG+/Y2LvQ3OBFhJPuSq66gtfhhZI1uWkYrIdeU0k287K9B+SmI82Z7la
AQF3PlLfFS0LI+Vuk3EquTIz6mHxBLww83g4LPuewHZr/wSzZO4RMKr0d2MBYvDo
voUR5LuV4QL0mUlEr1oidVxRganQOomAWGtZdsZRSTlauckN9TZdaK3u6vc77EZe
MPhy9tMD9e3mYqHTO8ngE74JPVchTpFOQhdlfJMbN638zIa75e7lISs/RUfTIKuC
nu7MmYqJZ/ULUqi4zl6u+CT6cothve0Fu6puzpUCrKAb8ulwPtegS496iWT++icc
kC3BjjHx2HQpWJtD/7srS8aMEjKpGFt84JoNKZSc30k2HQnW2aE0ZBqQ9Us7B3MO
tRoMDSaJqRjeBaK8URD8b6iIoB85yEsrWw/jNu7/8HHkhwf/kxgadRjl7ZlYeO+b
oNyZUWbRxHaZVYxWQ3hoh0ukB4qaZlJnF9xFmuYD1uEf5HY/vrG2WyryBFnG+sEn
NQSXzTQr21EoXu1T+3PcxCphnQy5XIiRnWla2ZBL4fZgIt34kwOqJpnU3MG7lA8/
cV/lSzJHext/OKvpljCHy6OnIPoUWes4gemYQ/7lJs+2QvK0qIQFUseUrrrihpO5
LlyxXP2Qq9JqCEDkH3jdoKUJFRlYPwZzCDl35OWKse/8sSczWOMoF3EGCGL2bplm
fstoBbMsnJpHeM9y7E4fTerYgxQyhwxSYMW7Qv2QS7gnmJIn1Ml0Qf9p8wnZ05I2
e7lyVitJJ3MquwFvTBOpj+tYr7XankQc1WRj7dmS/UNATZ3W1n3R/M1ZaXHOsjDd
se06yTtTgnpLddAYa3VvMjOtS//d/0xmUruEvERMFqJLkNKpLN3ZuYSQLcqdNRWB
KrSi6xNbI+TAvqOvEOjoDg3OynnuZdIy/qNjRIkfF2s/GwqPclF4/s2gD4vwTLCi
PtAXXXUbuMpUCmkuzeTwyAO7yXmUDgwjEaEE7C+H9G+BexW865L3U7eaO1snL/G2
cJeiPYQmjD2XPaattSBsic7GBqSiTLKtWusHdA5ITZ5nXUV8NHhHrMuQkAa539JP
qLPDJKf32NUTEWsyyjTqnsfg92uSyPA9VYerOOZOqR7QhsQAXlr4FL76RoqBQf97
f5ubxZY9psPetsLO+BazlNoKVH80F9ukVPuXNbuzyH49DurgQU9nGXKiT4iJWEKG
xf7hJ2IXYAxETxaUrrXP6SsNxjvo4G/Bn/54IHhUAUdyIbvjbqs2d9kVlDUzzkhS
6Dh5ERChMlCR1VqIk8fJSvmxXxXKkzq7NH+a2vpDAc5ArqA/NHafp5SMTJiN7QZD
MGXvHe4bEn4/cagCzBYAjvEw3dfY7JlYNQ/uP4sKFBY/sUEDlZT4QY6xlNNqq/gX
CmomFf5FiZBccuArRyroV+OgeuYEtbzMpowWEjddfp8c7QmREdRFx8UAwJ7bWNEi
P9jDQgf8euyeycglR+y3HixZpbCVBM3D8h53tlIrEXEmcpaEqqjdnnNxhxr097iI
EmF9KXsOcTsJKH8k8fmIZaXFg1WL2Hw0lsilFoRjvMxzKwfu2Y61R3THy7boGnPo
dFNVsGnnFfWvyQMhccRft3jPfT/YHGV/G+oUqM9eXPRHfHzpOk3CH2sl1Ozn9NIV
GRs+ZoJCQ6Ha3JlO6FHW1Nf1J+l1qdBpZbritMIVS/x+ehwV+5gXTqpfG6rY4nqn
cxf4qEW1WqQhBgaytIuH1nTsDvKpxZAHSHgRmczcA+REdyKC+xKksnBBBHYV89kc
evJfhMdm4dUrsBqoPo1JvOUXdQWD7i1UGbzLvqAM+HTROa+3w+0pY1WjBEf38Aed
UNDfqLv8oEZvu5f8b5pNI5GlOeqnB4synao3cI+ZLULcX1S2CmrY0a+A5klsZypv
foyG6c0Me7gd+11f4vgnP94uVXGJ+qMo1hKQSv6A3cY0+zqHZKkY2+6vWkfCKKaJ
yjXmQ7FdEFUkopWWyXn43x8TkYDaQmMrOQWg0XDcB6NdPGt7Vb5RLwdKALzv/x1T
URL/5LMOJpMywpiEE+R0kLYisvcr/Pq7zWaisPI7/lpDrAh/NDoxSN3kKH5qV7XQ
7fbNPeaOBeea9pcLLagnvrOnNrYTUHipcVd1bMl9Dtxo4jtn8zzGjS/fg9M6JTux
dl9UhtJmdBxtS36JZz9QFSgUWQuVKfXw1j71GqQGODCwVftQVU0O94s4i47DtSUr
E7X4a8rrtyHgqqoebumMSkPFc897yX82mJlZLywtF6oYBgdQYIZ6R+RMUDG3mSpj
wn4D+Cf0ZVNriYDH/KJ9FdxlTzkWhMYyWEqu9SSHV/332+EsZ9vXmrKuL8ngECfM
z2dCWRZnr3XCi7und5G9voZlXx+ICe3qiGBMlSAjSPwtv8jrjtbH4Xf2pUhGQsYW
OWxZmsMCOoaE3GPjC9hz5POLy6w0z+ioo5/mhXC4OlAym6XxvqglkYBNB8hsPGQL
JRt0Zu8GmVIH7ZW1GQhW4m0sLulatXSfv4mYc6Mx9fzRkPwEHzUv/QQuo2K0FcPO
jZMmdAqEwXuXpgLBLgGN9BrUm7qMq0Z7i9Z2IanuW17hdj9uP/1ART5cSpJDiS0H
IEA+GD+V6clKdXqBtXgKiyKe0CLAz5yzb2PNHY0uWkFmvF6MEZ6yS1EVRxA/H4/R
u3WtJ4zLoZL8i6SPzvtoiJaRjUp0eU+BEXA3lwCBEDU+81lIE+lCQektVPQ/AI/q
eOs9nqYLJYl+0vWc33Um2OZ3NNXj4IvB1PK7VR6Z2cIVfU7/xuoF24CLYk2U5U3A
Y8o6+z6tWicrbAN+fLcms+21ukytAUs7gtvjptoGpwjInhfSNlPXPseyEBEHCzSZ
EI/dDaD/LMWltGActA1bYnkwNdYoz/PgNkfKtbG2tU++eNBj1V/qxdhjmvFoh83N
KgTVao+QWLeJd0XLxhQMQpvue26ZKDRt4ojOg7Lf95r4bPNDD8y4Yeb56qZIVmBj
oGZGGi/iNLhj6bHZNP/HjHcHWR/C2XgyMjpBgE8ljTpfDKqws20azGoGdEo9je6S
S2OzWOTbJmZeiEvLD9H2BL0dptYG7oKJ+mLN9JS2QmRSTgXCDBJZQ6HLwBoBn0f7
zaGNTz76ZvwPu4WWInKC0UpBcxxkXIfqE6rDvEY+mN0HHOfV8H2a3R1ueG10kEhV
VWSe6mxnGPCH25t87ityxTMHTUHT+blRlJhd0S2XKrbnx7AY3leH7ly7+02A3ZK3
qrozqk4BoZxvxsci27LmJJeKXAeVLts89ZQiRpObFqxm3QkaElfcjajrPqWw7ktA
kdlp2aHWxZZD2ROYD35pJYFeF9coGwYTnhihEOolXVJaJXe2ECv7f1pFuZKULyz4
3cyiveTIVbndnuufLB9C9/wfI0/d1iZa4WiHSoGVUoMLP7o4O8ybIESIu56tfKTp
UMnCNgriXWcombEbHidC0qTyreZIKd+cLVEhyKUwX6Ipyc1HGwQsjj3R9z+BoRV0
biX+7I5CFUKpjjmXxoploI3Gj3UTUwIesIaumsGfu+izC4AVbmdKxF5HAtmDswYT
GHENCgp+BwR4jxChBaYtX+p89pu4zQtAh5CG+R6aN9Ig4d9FvfEWNLgyoHw6dbyC
2YNywg1e9PUFmOYdfON2Io4XI3GUDqJXGWshLE0q1v58EdhNhn1W4Uzp+beXgzbz
+IY80RiW281+KL9vlh/B9MZqd8nq0HCFDuN8Hj++kPGIDvLjW4vMmzXFijzJWG4u
hmG5m0iTBA/1zq5efuVUsU27CktMMSDd8W1dnKW5hiuohhxrOrlVKckRTT7SVEO2
r1vkVfLBGejdiufUIEyV68L3k/eI7sOPz/9YkUJmxRVmJ62MlytyMStTPWfr4lIy
DZ3kUAN8U7OeY5NPGo49SzlbNzGqzHKdsZvlc/NZY39ZlF2o8d/WE8e02qsH0dzx
gzp35fsbtwXPIoODuNQgRNiTR+qg87RJG3AIywFAPZtVd5f7JS/mf5LjnEVRzdoX
O1lLkNFZDylcstMlRPScFu26lwboO2a50Pi4X6TIlsZiG6wz3fgP373xw9j7kTgM
v4zswJpITE7rhjOW88lvN71kgO8yyWn3yMqMScfBIFBbmoMSJC27XJRQ6XFwwZ2b
pR9CsswzzwTEa7zQYmlAYZrvT4n9ued1bJFSGmDM2UELZ5oc5EbZ19Et3jSiayF2
fM0Nt3wKqu/KORkePdFxRWjc9Sf4bIHHQVtTtuDvu+4NiA0yp1G0/vlB5qP7PNSa
cQkZBR/NphxhCskGMsnmZ/qNsXS/5b1W3ZFnuZEEK1GDpxqGSCIeWJack+RF8k/H
cQ3D0+xEK/YE4yZTYQr6IO5h+3i10o6rJ+g5CDdTQCmIZ5rvxLH9Mf60Y8Wsnm02
LSJBUZTZqUSUN44YFXHz+OvM3dCqkm8soMV4bXm/NijZ+t2jwDbKkCEZIWE3Ecdo
FZ3RidxOst42k0eg2fMJzhEhFxHAmDrBIGoar3LP4YQBiV/34PpIM9WKecuM4MGz
NKr+Bs/7M7koEO2gT9vGc5OOCZcWLv3eCFvd8Yy6DiN6YUsoUr40xH+Ygn1M+uzO
lgKYs6Oe9HYUa7FaKhoFFVM4p3G0kI6NAtZBQ+itTSMClt9gHaGKNevhjMfS5GjA
GDqtSdM6wbnKRprTT69c7O5lAViUu+eXHd+pW3Znkm9O802gKzmmYpUn8NAeYE5H
yjPW5Ake4B7TbDA5l83JY065DTy/U6a1BaOBUlt51i6efTAKllmH222JZYsUz9Iv
klcpv5zrI5+5oFuOmxQ0cjS3QYH71pzbAJwMxKAyjXytlfnEPezlcqaVcOq1ydDa
nD8f0euT+W+1HKYHXwz18rY7s9tnnQBY2Tgxn6h+n3i+x2OrbJhVqe4YCHjTfrqP
r055BwnCrNcdS7seWVRciBwEvZL2oiJ2jJ1p/NPFWziWLrFeMgVBWwRUkWnXkX4p
LosWZAw0B7tbXUcLqCW3+T0jj5EtXcaoso+Q3VW6zT4qulUup5sbt2kUgIMPmlDM
7qStWxSO7LSndS4Zg1rwSKvQm7FzRd3NqIeoN+oM+yMVz3CkfWwrChOCt7QX9mT2
XL1LU+8C1XRrJS15CDJ9oxO5kfrmp90uJUgNZv/ow5RqBSMTBxDOXQ0oTNSUmL54
8iKiO54OxyqCzm4EiYVpqinRD8LKPoLwIs6oB6a1JJncQTQTQzEoEGOZzDqX0p3d
xv7Cr4rgbcGH/2M0pO4Cx0tp1m3PQeBiXsp03c/zaFat24zvrMy+aYpX9SUrCjgj
6n3z6Y0ixfsQdXMaAQnsNkxhO/+/MM/CF665IjfAUt40R53cKKdmZ4wJvTiBLU+m
j+elMzu75doxHAdSunJ35aOU9TLD3en/oMb3UPq8V6qudmqsvb6FFnDVmxAVajk4
wxU89vFZCjfeeiJjjoeredkGl7yzDNhR6ebmY3SslNpRxYra3vEd1aTv1ftIeJqR
1aapf8WQm0X0wotAcsy7OuTiKDYRslUiSdy5+FEq9KAMouJ5j6heOLBRT0/BYUCn
i4FlTfZIU3HawldJWIX3iR3kmCEYTkclYOMh4Tlrll2ejG3qQiAoiqPWgYwsvrQF
TFjbszATGyWL5aEBCtlhY+wTg0m0SS1YzDeA9vfH5qPLI5Td51wpzvnWUwj2J38X
1NkTPMv0tZWVVh+tbMj8YCxUZc+ttE49AK3ettL0YKAgNx8zXOYDbWXqWDcJvVpD
Emj0kaXf2N+ii89CVWJyzFOqR2Vwx7z7c04//SeKkczBA+WM7RqZBtcvL0JXwmF3
4uEFtqcqv1uJ1ZlWH7kdI11OroBYfRKPT/H8C2ycauWZaAXuCJqNJ1ycT7TG59OH
/eWfUCm8iqju2153+Pux1ZQevXG9gS3+HMcE/buFy9G1/X+Heg/+sPag2L56BXts
y4u2HC232YQ8gAASH1KCumVo8Ep8auVTowdvkdKPnDrzTuVycHDtGIifHEvuIa/I
d3Z7ShWhEQs7NR1WzKXDmPnjej7/bezIlw2atjKqj/wTp/FpNM3NOly9niTBiYO7
vtA4+PIY/wBbY6n1DMDm/e5YD0jNxj48tfW8uAy3I0p0foRb5NZqJwqv4Je76VZv
/GD8bztjb4ZK+3KySY1Mm3HPZfbamoXT0XEOyKUPnc7eTtBKPeWr7WZdHN+5red6
azcWnXEQVRiiEjbwogZ1rYduZoFhgBa6EIuQM0wBo/wEmfdx5n3hNWzBIZVwKj4G
6t3aXSc7K6MoCbjWCUks6WHZW1TL6i2iNHtoOhJ2dKpdl3003VMWKL3gqD7gazxO
51b7jaxYnr4/45iZRI1tOP1YKlLPGHTLyeBcaTGgnpSv9fBS4KvNPpLiHaFEz6hR
/1stb2FxPP9l9X1b1CQ7tF6YqIjGLO9ESLvK7zHIEcVDX5mzR2q6X4QbMKEUiZuM
lIZlwQRfFviAmUaglfgJEwAyaWel3kYhWWOcoE7sCuvIhbMDx5wbp8xfx9jXPjN0
CsOSwPGfF4jqpOtp9p/1hN9VT7dJc48pvwBgTq2cyOIgakXkL7nsYu2TIRDt8pqX
th8KsX9NRGGmFpQC7km0uAHDbww8IhmAIltJC7Y3M4clZ7MruBCEpGZqtgOCabPA
L/oG1cfD59wL4Atitom5ZU0Oh/UifctryCF7mwBIKm14Ir6HTDOjhBsnYseMnh8R
Clo6iLIHF5CjtmMkLZJW/+aMXX0tPBGdxfeGmTIHV10LyIKL+vu/irwrEgvmPV7n
6ZAxc36tTM3wXdF0yNVkUhbdCGwIqjuRsAbWHxIlzZPeOaEl/9XuvLIJ0O1oBbWf
88hBDu01KHW/ZN8uhCEeYJ4EhXcMfdtP/GJ9CC2doCghKBMTBh9dw1bg7lyDjKSp
Bj7S4qHvjK1wy8i1WwKDlffUZj5gETSW85YfdNfwhXJ3RGhF8w9sXBHbbM5/3Kon
cFOB4g93ihac6nLMLIhGJNustC8XXa9i7lIV0veLydlvQ9fsu5TXG36BXC/qf6F2
pTe4MfdC+7SDzFblFNbJl95+Yli9zxQViKkO9bJ9ozbIdh3MTntqsQbRWNAHCjwB
iBdlrfvTycKP9VDt+NDKhQDKWwgeq+zJElshzQ9zv0taj0NQ9P8ke1axsUrM/UEs
LGAdlu3Ms68k21+51SuQ4wNlFqXxrfAqYuQkv5sEDG1qe6Ec16CTOwgTQzG/dGYg
8JhI4FUK++PJ9ZY+3nZmBx9r3Sps8iRjdjeR32C0tjhsMIu+EmPVN43L9QI8jj5p
mAbTCEJAUzcHuKCfoDwQLQUdZV2GU/JSrXSC7zoadjwgXtnhGlK1gv+aAlLcZ0NA
VqoASGgbRP3epyOPWFDINl+ogGcBtj2TG5Jf+QjshVz62yVRW0dfzRRHiDKuDcga
vGRocT4mQqENor6cfXX6f8QKdtfi7tiyNPfjp5XVC/B8B4vPlLFHAmGP2e7dcUIN
aJU0ZcLHedJtvBFetzoFWOZCUWnr9fLXWjuh2r/zXccqPFLVWi4YD8kHOhwocucY
OmxVne0VKa4DkNJipEerV3Lsy8HS57yGZwlnDSHvgLbzZxMuZaelzm7FEMYgC2kD
YBhfWs+LkX9Cb+rJ0asPACiCMf7lJnKz+v397406Nkv721ARxScSx6WB14lWulI1
00O/MjZo7CTWsGn/5gH9YP5pQ9wNlME/ZgmJC3XIxnhKDDajISuTKNTGfF6R7VBv
M8/kLy8/163wJg2X5CWE9Sis/r+qb/1n7SgXyj3wdSv3VqO31XZ31B7tce68decS
npS7J0UFK5zaZ8lsglTGaG0SX4wRGM4Yf++YKk3G3ezjQYO5yx2DcgXh6lcIZkRJ
owCUjXgNZuEHRiztLRv7mlyODCg9+bCD3lmnXmJIA3Dew5Ubdpi2IMwCy2JDws6r
Y7jTagm5m0a+UrfVpA9yFy2Ygei3ndin0UiY8A5byCPht2phazQTnEuiUJc/JcK1
OURG+nhcHwwEEzVwEW5m0Y0ZQ7gz5q5yBZOjmrvww+LRXaeFvMNUCaooV8t9EIPs
c3NYk46TZmlXdnkxQ+vL3d6nmZr0DN4IjueBbc8NkyYdlJhmmbr0mn2oqe6nS+sw
jaM6iMAcILw4zSfTZkDWkmuKQyvn4WX+3d4jPFQZCBxYnk7iNx7mXvbJxVn7rvMg
Ht/xFLZaeF5YZJE++XHmK2aNymo8vYfNiVZ9/3AbKppCoM4hdigRUYKatk4S3tuw
NqpBwyqZD1yxkuO4PR5GJyAnIsb7XdOTm8HeIs3L6rIG+rX+MTqqrZtPKuEGUbAr
VNsTfNFJpknmNtqJqZcfSh7nE/N3KwIgkDcQeS9vp1tllzGPA7xmyvof31EsBYeK
koN8tO0icTvtLiketV/ZA1Vwm4I4HeYLlWiSpNivndZu294E5ptB450YrhQ28AX+
F6TC/uIlGJDHQD6PYH6Yh2UCAqA5f0pMJ7vdQaAsJGcteQ6vnHMVCTTNP6GVKgbz
gBcJ7ligTiW5pUEL2kfAL9x/fGQitxUY5/C9gJU9bmqZ9cozrRU+T1UBv+m5cZ7L
TYWvV7P5tZR8OzdFsy+SRXH2J1gvgKTX1Dz4wwLCoH+Vt2wUGUqLQsx1vt2o3qO0
KsZ1GHZQ0bqv1sfnGj44yh8jQvw3F5GFKgdRG85Y/SyC8tKpzcSan0x6K+PFcrDu
2L0mzfyuNec7DpSQttXEyT4LUUJr3lD2EIAc68Ly5/nMCO0FakelHJIlJyBw+M+B
t27svNymnrPw6WG4jO37ntb7PnrDUxSjEJHi7/asZOuqcvoDIZiszwN0r4JUq/C0
UmThxnHmy/oe4aSoJZ0JE50Bx1GtwYZvIOgvaAAhyhFJPo+8p6YXT4M+PNASJmYQ
LjB8jajM3AoA/UOrYYviGnnJHjrGTbXUKR/PBmRT+MZeCY6RTcT0AEvjEpJbDr8k
6QRV9wLFOHk/Zp517iiOFGxd0hzThScA6mr+JRZo/xi4ViHYHWwS98T1gECbPGyC
uh0SiL1ObEDamqdR3XFhl5JvekBNq1juXRXEGP2qQD9cLOsvwPyHA3k9DOEqdgbG
nXzD1iRKBQIBjkuduw0/I01GQvtXggC6SuqksqpxDbS2psI5Ab4Q37hjCfimm/2I
sUuH0poQ05HLBpDTMGSAv75/SX73cvr6308WNFeGl+XEj7sxV+FVl+mJIGFygayG
B9UyTDUy3C/HAh5Jcmm7xGvC9hGux0Kk1Fk5Whs3Ny0SLC8IOug2ln+dC6FkX1Z9
kv0LLGh1ed1s/B1derexecbFwQEAGjUpLaLeQist0mHU6u5ZC9q059Ma3T7FejQ8
j6CLHycKkQaP3O061OMeqKIyYQRmMIrcpJbCG9rXHXex4l7tZ6AswDoGyuiGYS9I
mLiJbkh+9moLgSZeYDtsMSZ+ApfIQGfsb311zU4jC1JQZ4I+iag1V7tFyiWZdG6c
C55r/bieEY99ZlIFrtoAxPX6FdTqCr+WH1s5C3iCWegbO4LkkdS6cwKUqBgY6aWg
HzJhKe46BV1MMaPOGCdvTtF9CpeI94EIebZ+n+T89G8BhyBZHmE8hssX9Otbs8CB
Hf+8WV0fg7ivqf8qPyltazZrUUlFrps6JzpsNsk/rcnxz6YFvBfX83qnR7JzRw/r
vkiC529nQTAFGM8YEPlMIEwByZosml45FsWGjftjJG4g6xCRf/2VjDDvRLj5o4cY
Ys5UTmOo+oYrMwyHl57CzW4Z8+Qld6uKyVN7kuKYOgTGFKYzrz6DXKcbx6COHiEv
IPArTbCF3AHqAcYRTL4ijZCHSl5hRwYlHVvuOHGHyaiPUvj/Y2/WG3z1V6oP4dq6
2e+ILkPYWy/gWilkHv4fSR4EULTD57WAz4ejUgP91wwbxGUXCw8NgQIJuFMaqC4q
/9cbnbTyImIAdLS9//Z85KGmPwObkuq5uYe+40Zb45/vxegWJ6L14PGUcplvlVQn
knNraG1M+EsS/T6tNGkHmFzZcIwNXm475lT5kdadnHRDyyPQa/tNZEYsWW6HUIkG
+ftZAIoPn2rA7l1UzuL9gG80rfISXoCfC+6WhQryxWPQt2oSePKa+swhWMvNUMkX
MbPxDItrAtvzntxKOv4tT/qIW3ZdcmUcnnjDnyNqSGhVBoc8sSNcVXe0gMDZ4B5S
UJVFFl2KQxL7EQIlaeCXfxxtbCRO5yYNSUtbBViiIB0nT7rflEksUSAhQEBu68CC
etMmRhRDOsnPad/vWulyEk7lnPiNavsQmSvlgzsCoXQpAw/MDUW9VzG4v6HXttht
o0T33hJxf7MDHP3i7IsxSr6JOJ/CzYj6j7tEDtyyimdku70fwk/16kDhciRsYANF
F82LUcBDdF8M3aXNQftew2OyZNikyiDCKkI6fggPUn8qjcSRRLb/siQypavqW1Pw
iOdkYWd8kGp5tMJRzwcco7TCOPEv9cQgVylcf5IAIFODB9PCPuk9aSoSd3SXO3Ea
giQBxpAkE3oaJSaekkkmOSX+YRaONz8l9ViOut1/VFuBEYqs/Y/Q6gC6XhhZrpX4
wxCDJqmttxaBgvNVFj1v1c2vjUu7+o9Jy8QJNaSilueVdcr5RWMikfd2LpSemIn2
fMHraoxNhz9oxGRp9CqUJMP3qes9dFHAylKDC2XQh1L9H/bxvdsmGxpfA25TGwWm
PgOathopK2vosDgrZEJSO1zWEYTdZoM6Zf5wISiPePCUUJXJ5eIqMqt/1d20t6Qz
7LnaQZc1HHGSraADS8DvsJUWZbyUgKOPkDy5KvrHyuUQDBcJFGPyaeLHlLESDxta
A6Vc1G+HG4P/iAHF1liN94txxm5VJNXboTZ/V3Edzh/BPy3cAMwFsH6hGo0fiTOR
ottShq64dvsqYeVR9+i1p7Wg2AVuh79edJzgw1DYWrrR9Fj/kgYrx3ZzshQuefkh
UjiqRDd8EfsQS7hlx0eJ738JramovVbu7pBVL6VebLAf+IiTCmbRU5Upp5kUNgJ3
Nc1pPdW2KIhvbqxAIBlJ05c8Nu9L6p5iup3N5om7lJsp/4mVj39zMMvLCFMcZcu3
Ozowkwbxp84fG2wZNEJm8zCTb3XLVsFAdjgDGB/tVspnjDbXInNHcSum3jNm9t41
hDWEu6I2bWA5JaAsS8a3W9fK63YkU4iaNUKjT9JycFHXiu7LqTR96+Zxs3ejSV/o
kIDtZFKEsnE1QOHFXqyILhXZ7UFstgxHR49OmURA5HqJhUMwbETIp66s84Ocre41
Dz8RZS9Ge7dL2sa/W+jGC3u6KqkiIMjFd0nw6nKDEJbGQ8sEMKK/4aZNLTctA5Fp
YqEqWg1vK6Ho2+S+cLXgTWdXGd6oOGUrj+8rYwRzSIyZimf0VRZsoOh+XxABWmUT
nMPlB9KXXH/dQkjulFOKwF6j2ChovRP7dr0AG6CwBWFejCdO/1z2JFTrtp3hzsc5
tMUbmiYGOo2DyDRzVzmU3u0LZb4lL4oJOno/8O/McXRCpevohhbMkepieXD1dii0
KsjmztIJRzAjUXGpcOPelsXiWJ8KTYrGEl1PGCbTsN9MezegjlJ1FiQ58a4P6GpL
hwOW1zA2f3z3Dis/BJIK8DsVh4/sO+NzCfMJIarltauDyGO93ru8L9C4GpJH2U1q
8RfXlOjg1HyyT16ypsZT3V/JgTM42rkvMLnPPd3U3guYbkINdAMcWgaWeiN11qad
uLVhn/4uGMYg4IZEm+P20HIZFzlO8JDweRtIHTuhmowTWVYshmSkmJ3aMMkqgBsu
iSergnrrCU5/WCM3j/XG42yuQC6GPKNmIXbWlwCSC7pQfB54klWV/KtN39l0Ajva
DYFltd+276ma8pm6Kn0wLiP2pCgwJ0AkVfSOBY/fHygiiWg556gPKWWtGUwKKHOa
xMU7jjurFG3LdwEvZc8I5mJDBc283fwJh04cyzoNvnZm+ljBTw5bMzNxzz+UMDoe
shAXuliMNPQTdBr9C1t+Uw4OE23vxG+G1O80rQmtTvCfo/AMxps66GdX3RCoVpRn
r+Tg/9Bq2X6gyfye9sjtrMc2C5sQEzWvBOcIcVAYx+DCqytWlgu4tKDUNwIECtX9
BytYFYZE+61FGLtT8mXOxc4PZrZ8Te5XRkDVEIKyzK+zv+Mi3+cv0OQ5iSvKqOHX
rFIyAV+0F+iDox9TxQwIA8AAUoi4+kqxUGgUk2aWe5rE1doKpX+CPOqqapmprz1B
l4JAEXqK2KYRuufAnliQGfjW7YK4VfofPm7YL20dRRUubyIJRnWRqjxJWSz3/WHG
UcXwXwR1T1BNULwpVHuwiXpWVwNZuwfxcu+QsanLZ66B9MqL1WuLu2NTsFqDZ4Bl
kNiRyHjgKhMKFddrAxlGmquntcED/LdI2+88ogFafvPgisnXbSZfl9slXpbc0bs2
P5Nf3VU2DAGLKKNxIBm7d3dEwZLzNWeAYgoKx5KdQCrctm3bzSunUNYMUw3bL407
/xp7jekM8XJBFokmX2r4K7k4hWmGhve7PJ4kHujWJ/Wjs+JPPJbkayrZXAPPfEnt
Vu2XrIx211EaMTDDjgB+AHX0zSlcbyGzPHtok4u1k4v/zYSbk+S53z4hwJ57jU+o
8rT8/MznXfuTs/LQSdtZvQ==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Zj5kro3/cohgWve0fmMg3sy7YCpwXZtjUsV+roEBdssP7Yb/BzoPkDJtvs0KxFld
0YtJWGu3OfpBfPojBlsnFsDDgpVzrFaWW9f+jYcb9ABXa21AYUPuNfkunWV+XLZf
q4cLQnTPPdiJZCitiw5ASntntsDHrSszwMX+XxJSXUFJDzRM9a1QYSO/40qmnyIt
BLzfi7/QMRTBrMQ/apAKLce9U5MZ/XlPRSeTUab00ICCHWVYQ9mCsZQUkI9sVeqL
r8nf/PouTCZ346jXqTyccJF0jVLSVQi4L5SB9kmFCqQQ1Em6n+CFYe0rPrFubH7z
04Szj+nGpiGld58eD2MU6A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2016 )
`pragma protect data_block
YZVF5UK6GRoItAEFSRWfG+xInhUg1ePcbz4bzc7ImQpuDmp+jKU4zdAPSn3SiDyK
FBZoTofI8NuwZ7S77h4SfR7/3TL+zSzJZHAA7lpBa3ro3mdFdmS+2R5pPGzTMRhD
pH9jUJ+oPrrWT2CplG78aMvr1Q8XVcrTiGESLxN+XVM9HrkQSDOgGNsnYlrbGszo
3fpO/tnCyJfrLEtYS8/bWhP8nXHe8dKE6MvzOm6R82YRh3ETwiL3p7YajyROuaI9
EmaQC4QmreZD0e2vJEbpHtxcHOqEqr9bXT0F7krReGE4YhlyVvwscFl7VYXaQp0f
T8SoqSd+DQsYF2ba51W6lYQFnElmPSSsR2zlWULyoBplYQaX5/WXwgts7nyfbyox
UuZMZ/kpIkbZO958pVMXYSiK3a496dmqIKscAtiSxwFoFYJ7ycOkcKXU+63jtipW
Iik1l+SFD12Pn/4EyKuAT+NU6heIR+jvst8m++iKmXf6KYpBE/bUQdrftZmqCVPM
R9XJxwCLiEnwAS6APrsiomiRKZIWQFtoZNOb0hsP3g1plAQ5DVlMGjO/XQMDDh1z
mH2Qvov6evpNXQzNi6rxojR8Cw0Oxa+0+tBlS9gWiIwADc4KemDosk5uQjAYVFC9
yIdafK0G8OLwmjAGk2t+JRi7G/rMmgIA1nBVUZ9IT3lgOGx6Pc16lvYD1J9OteAX
dZ+kEfFkASeUuVuQp383VSIBa7lCWfPGcvScug4uB2AUZlydrCFBxL+eF7E9e1xU
HCZ3dtzOG/itupj0Vh8AWbTOnKi3Hwe27SSdcfnwXd/lEFHUm0tbLUQN1ZSyzBfD
HD/rQ0/r4p/zH2e1erTz+6lTSJpntQuNpIGfHbdM/LiPnAjB1RZ5Mu34dmraHBtv
r0F1veJ9IkyUa2aXmoUMhMcU1TJVoTkf6rv3NxwxZoGkT2dxqAbDxsMRjSkj1Aie
CHDpvkkz1mtZfrnu/1j+XpK9ergWxV99dNmhx39VCK5TaMITsrc+zmcF8rkx7n4Q
9fFns0qh9y55b8yYKxs+i71eb3MB8kDfhCWU9GsBoflr/QV/Tp46fVObA0d2/TqN
jb6wBFcoY5X95nVuGPX9vl7SMuNRsURUHTK3qRwZ2YrkHRKPUwPdFLnN59Kq1Pi2
pXy9O0Dgv/WK+uA3HgClD5+pXvHyjfnmkmSgyVycVbU8BXQHwq9C0erRSWmfcnwY
2yIDFzP4NMP2fGk/oSt6IuQsBRaL0VUurfcYEhvjkQ22VKUcCcJnhH0iVgRGchOR
KBzg/vLxg2VLou3JV7yb22gZi+YChO8Hd8ljGOKmjB4kjJmvFYmz5LIMZXea+DPI
pq4dQFD3n90jUdaC1Q/zjA+98fmDk6pUHLP62Lf9GQ3FmkWcscDGk3aRlAP1FiUn
aUBE39+biwii6rOGNhQOGArxxqH5n/Euwkwfd0l4AFANUlQA4qjkPElZOQWXbCUs
XgHLHsFqG4xA/Mtya+bImxqSBfAfFTYbfpszUl2kxZxnbCYc87WOGAN6KuH8UYPA
hdYPiukxtI9dtltvR1ZCXCcgxY5XPhy/E7KFtm+qt8/8z3qpsn5aMfNk/gPHWCOC
T8nvbXng2529+tC5yTsBMTpfK616GIb4uy0oBCrqlY4TvleB/tQhnzK+7X+Ck/50
mJHH/jPSltsJC91R+Dr2Qj/FuCf+ffp0KWRkXkmgvjlmZJOggfDeqayrLOXlOp9p
RMRSk5HOrUQ20yjbGf50yiEDib4ETr63JU9+dOkx6TSO3xtpzMm9LzkXJQ/ozcYK
i17k1U3o6N9FwcEy0iyAUHZ3nk83Zmx7foYw3Lx1gL4T9hgn+85PjQNDvnz4xN0+
bHYMLHCs1og4Pf4AKIP5QAOhooi3JgdPaahQTRQz+n+4DWxCyQXROet/15tKPmxx
JOHGsCmSZtTKfGYQv9oPkgrEkT47baX3gaqAy+dJVr2oRm/pUT63RQ9MtS5x8hCN
J08GclCwhgUzPj77U4TXVNg8HOTubgv4hpStz55n0FTkKQAGkYqRPkqudSQwuYiw
nvUZX+oVU2mcX9Jz45WHOdS1He9SEemXk5TCFa9zywH2kjySPxu3nOlZbtNY8wZ+
Cy7qO6ezR0h/q1ORrvSrU0/jnCe7FhHksmG8MxcXY9qPcwKPukw9VJUDn5Xp9b3l
NpjQijC8RUbqn/g1oIViUE8zty9SKja/HZ65wvIE7+DvIsEjOfJTw+nZ3J5YZsT2
eURuunVgz1o4xegxyrs4uBqbXse1Ndypsdwb7ok528CeLb3+eOEK2r2x+2zJjbqd
u2pZsZvz6wcXIGtCffDy1snk7Q60fz1YDFHFTMU536UCvpSgx4c4tBlkGzEL8UbS
hYXSkQ8EtSvZorI4wcQWywnHGNwASJzJO03OaAEpoF2ND7oM1yye2b6bh4Gk0Ea1
c0X5VoasrzLetZLoP3MG5bELwSvMbHS8ynDHJfEAVR5zX+GVyIhsecmLyz0x5F9L
ZJyvXsv/CGLk0TjBSTk63htSPvynJQ1E/CDjXtWPwUZ2LeKb4IylKe+IGolQI139
eahEsv9B884eK+PuprRkxI4rOrORfa4CB7lW9PzTFBIp0HEhj1pGPJSHtaNSJb5P
824RctSpAFbVbKqBJJcEYHpHf0YWJtunElOoqJintseiS/V483NSDynsxh3Buy2Z
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GZq5GUgIdzbNHUvcY8Lkpm61Fs56co5GlFhCgm4vgKKvHLJAHQNkboA2wLxb0uqg
B7gu7T2xK8zGjSzhgar7UzxL+vSeULwnPskdxzcm2loxP41/+ep51wqu471oOekq
t5STJlaIH51vfwFohCbzEfuSWFi4KXwrJcvpshrG14xJreLqsL1+48UmFiUemvCT
AX3Udd2gZMER8ylSArdpSyqx6UBI1CGrVM6o0Auoap+2iRAus8ggJPNPowE++s1a
N63P2A3Sad+ckzftRl+Zj0dGTPhyPom93X9MLT5FOw36IspAyydc2PKcKT73XJhw
Se4yt6Ojwd3aHfXMrixvsA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10976 )
`pragma protect data_block
S3vbOaQZC/fwLxHr+LkWUR0rv2JXqnY+6OFZ9cdDadIfjEyVA+7w0AiX9eDwlcU1
B70osQJj4oQqbSQlDCx9LClIWiQbTX8oG/S+GwNeIV+qCBttwRfi5AIDYH8rH+1p
D5pZ2cBbXFh7m6o7ugeTgoo3IjV1xJNcD+Kz/kxGm2OOVGeltBO08PoUpCXH1UMi
MXAsn5/JWH9v7huGJrpJbhRTYOiLVD/hbI79WEfbB4GFneGe6vAUcPQkb8Z/J/g9
YHutVnKU/LaqjScPxSc/b8IxmWl8zeQAmUGn/VBRJCbFKltfsxp/bTJise8dEjxJ
5/Z2sAEjN6XYEwTaATGKQchTeIMkBfCrwgC8eAPVyLK6LrpOoVfztwv2oKGj/E0R
If0/qXZqc2YYEttsdybkS9DIyW716PJaMnDqiGYFj7mAOPrZUwUMPoxkkdgU0QB9
upJrg/6OaNCfQAaFmXCndCEwk3NuLtPChpUhRZpwbphvGriic1qJzo+ikW+4O5rH
l5tT9ChnsGUGj/uPDaM1tTb6awneei14dD8Ex9fVBpvF6DDN38YOBKaws9JA4vec
dVXXUHHOjtMThU4jaqmAw24bG+NJV351fcAxCaGXDvUN/Nl6vNin9pF0pYduUTdD
BB9gLayU+dRRKCn5HhtlVRDGbXy+c7a/h00cddLouRDj8Ds7puwSgDEJIqAiPI0j
M5LIw/p2flhhZEq+ugpdqLuMrk9hHh8x7XQ0D3ZcpG/+pf21eziAfBPVgcD4nT68
oZuDjiSFTuUNVbnsQSiU8IZpZDkWxWlzJ2Jt0z6yCjZzpaDLH4RWzzZ87z5yZBat
FnYfhcGUb+E5c5JqcbxglIOn2IJp0S12kvQRJwrRV00W9/7+DzggqPlFop7t8Uaf
8M2ppZf4sdpHbtovLNOO1NuR1/rNpZc0oQh8143nKC+6hv+/jQ5AmqFLj+jbzaaP
qUVTn/Ib2nFs7+ZAuExtFvKf+MBc7lIjCPAlFoU60shpyXOcCCPF/pjbRndfEDAz
hbfHpKw5RZsUWOjJ4f4/QAjIDtarAZECqvlfBxTDa8XgsJtZKGXKaUsDfn+2QX+f
ZIjIU1f/ay9mmcCS5J4mjb7m0qKmXuojfq/BDHYo2kKR5TkCzMDi9dflB2aSGVNG
kc+HQoQqOzlY/Xk7ZTM05lrE9K0gLp2sWrdV35QhTJMi9g0Z/9WCX1ucWY5ZbxzQ
5NKU4kHThZpHwH0hVTA1Jw7PTEcmBx4dFO1rg6AghGlmUfjsXrsQZiz+hLBB600+
NkSTHAxkudUgcgU5SF/rNtwOezOpTQFPcDJ3NVn94T4L1PC4Cw0ijk40uf9fd1Ph
svcsn1qwlVve92oTZAWw93+bdOibUuycN7A9LgzaWB1zY6eYmeYi19/S8tAKxCZq
q2HBOYCZCNjTFTBQdsL97JHqEgZIXeiczdcfUSR/WfmTqjXU4h1sXhnfIVLbRlbt
GX1ncOi3n4l3fOR/QStRi+hjjRjjv3TXVxFTr2xbarRVFYQwlb/sP+/2+K2lp8Dl
OKqxEYgA3N553o5+4BU6lkjjI4+HQWTXxqCgXEvHy7mmsHV8qZMl8Hxq1G7yZh8G
LhqREO80tovHaHPiWyGJtlw+ALao7wMnqUDycEj+lNGm0U/OKzoInS0IuI+eyEvS
cn8Ub/kI2SY9DBeOBEYBoW9KHGOACCktl7HB5iKe8TFB6y2cZju8pm2MtQeH2+cs
rSnuSa8zDcmjVOjf22lLQM7vaqFMw5H4uwwW1o3Ht4coDlUfPWIMjHalgTIb1e+F
EBTzWsHX+3i70XkormdanfRp89eDDmXGTWxRw2gQ0fq7cwRH7DD2beyQewnB4+4x
/uJUrFbjJ+LYWUkq41CoQ/7OruAwKDRvvyXBrCDUKijF68CIRUM+aZVZU8BZh0PP
ufjIdyOjqoBr2QU88l3MHciaiIDqrJuT3yC/LA9CRaqQJIq2H5oZhAXNFqHWuRJL
X1jzXygZC/lhZ92CNKaevXP3BNijfh56H0YVctiBxErCwoVvHHJZ4GNCqVchciXJ
aB2TecVfefv68kIuPw+1zCL4HPno5nYy4zyjebzkg2TmOIM+mPEYmn3STGTlV2E8
5In9n4AafCofHJjkPc21znQb2pK+2p6MMm4OLe3zPl0UkYvH6c+AKEhR7OKmJijM
rNtXBlphGD+aLg0iK/PHcjA3btRMLC9SoYFZumtQFhT3b49wvU01hJIBym98iKjH
lZ9+H7ZjCQoUi42UVzk+kHvLidl37c5j/iQsUj8GR5+a92okjb1vj2y6bEHBAd0d
s+puzG3TJrVba2snoZdbB7gqcW2OxrPOR6tfWRBj5KIR0JU3PHcwtzt5ThAD43O4
RVzjN4/i+D0GpZzujdcqTpqCb115myN3i+wH7otTqefd4FzG8P7igTVu6x289D8P
wzQ58Z+RJK/gQ6rDfQN5jdNO4vkDbF9XUT8Uc2qIbXhT7ECDgFNZpMHZ+8Sl6ds9
0zYGVaUz7Jsj/ojypp7mrlvEvrquiU1jzdkwf1Sqleo9m64XanwNgVBQP3kwMYmi
qeLcI+78HBGmvwlBtHkctj9OynNmVSYmb8xphu81otV9dwlgb5GaWGrl8qc2ev5o
0D+gWxhZ59Jp5yctH3UrLO2wTGsM5GgeQnv7uyu4FOh+cESKCKRfnxvxSWqJQq/9
IgZBfcX0SLAazvTPtknRnrD9fDHrhAMK+orAqGCUyhtS4ibWp1mKz2eNbFT6odzQ
bcJDTIjCkc1QT/JUGginQrejn4wv3u/Fvb/D8yMiwfQQ2rHZEZ7Zpz2Y5D/p28Nn
RL0oGBhXZvHGgieAkhedGLAzyrNKvhga5YeHjrnwNhuv+hXkc/2gSOC5V0xVyTyE
TOODDr8yneEpEcSTDUY8Gy7472QdBnZHafE6kry5Lg1LqNCe7kKcLZl1xw5Wx6fB
2LS6eXMglGG4qufkpW+7gQHmkNqYq2oNdqEbWXeajxwQUCUhXSrg08H1cZI8U+TA
QrVnDoypfHplMC9nEgOnFBjLpzrxeSfNotVuS2TYXpSpOl1QAxDpXJTR7E+IwLHL
Etn2QnYlv6kTE09yytyX0Q6II4PwdEuyyOIc5rDYlJzpSKO4gUYaGbLen9c8ddjM
PlEYvolYiEtY1sQzfCiFNqiL7KX9C5nJfLj9+Ht5THrfSir+4lyCCjYGYMZ/+cyQ
6gKCi3Bv6iSZ4kP3JEc24Xl92SwlVLorymukFB6i5VrqTsqo/poXMULxHzkVJAxP
zUBHhTRBQ7kx+whJ7Sp8mUH1mnJV/rWFYstpJhGiLsuYH5DASRzQ3wSo4/EV8W+m
GoQdW0jTZV+eqUlW3Ba743o4wb5xOB/ueQu7J7TBnnYNI+XhYA7cvkk3Jf1aihX6
bAmYe6SVx+ebvGFKXFyCO8IKarKQwNjETWy6sqowc6Lr9kxfby4V34kTNjq8y9hv
Ffa13asN5pA61yzAQ/6KmoxF+guHHwJDGnUu+ghR385cPFbYp/l23tCCyu0K+Idq
KgU7AIqjG3Bsu+BbnfFgBom8cg1H5nQPlShnBrXtKGulyxsjt9u0TO9S9kCqwukS
+j2L0NNx0NcLGT6bDHlGyhDVOxe5ahm0oi0JH3AILTbO3IuBIt0DlDlmU3+3d78n
8Vj+1OntwbqqoEvAW0offoOJZFpAW0oq7tl/QKEi4qBfCAoftNMrUtZPd4LbvP04
WxOqF8ycQwC/zppqXdgaC+DsuwaBWGIV7VI9TwnC6LsqLX0kVSm4Ne99KmYCe0ik
4TfHnoJ0FHokxzm3n5NkBj1zOKKdKp+Qr9KiMnPPyO0W4xifdQXgHCmiEjjSSoAY
Unu6Lf5EXKvyCKHQKy3XyXUAFepkMZRwQLgqnwlQUnOwXyTJyyBRoanpdai2y0Gy
BH817tfdV5T1QnRm00nswn6VPX4C1FE3wLGwysQSCU922IrXo9jTuysrsYdFVBIr
pV4QmjuR7nMIHysmwUPJVyNcTZViZYVblxhR0VBaf/cLFAQrsJagmBDYp5MAsMea
NnrmM/mHj9Cw0XPJs41zAYD4LXOSxK89e/+zLuR8DWZbHU4JwbPl9iX08zVQDZCm
6iQJLBhkmC+hdzpZc9h9Np7BNzf3/RWWYOYNWsEwJQ9q88V3eBQ5rg3UL/eqnqBY
TsAoTnwu3XwEQ+e53EMWpVNtwDPj6wcuekmgWV1vd4qK60Bw2Vt08ZrFE6oPG4Ke
mIxUxW/w5tXZlpFO0SudCnh9FFkjpAW2mbd8gk8tcggMbT+C9/ElweRKWgiB2DOO
Kwy7s0Kcu2bvmE0CIqUYgpaPsBs4Sp32beglLk2aCffJNy4hgIuIA+snYJSSX5aP
WbzDXdGM5sxU5Vq6sQhiZ3a8vV6QVl7hWCQ1Soe32p8p2qh/tFAr/b/rSOUTeXPm
uNXuUJDevZZQ0SpJRbdPh52IMmYkYS+AtqCLqydsZwLn7n7mCo61u2ISaiQpHgNW
3aiVn/QSM+GU9VvrU9YmW22Rb84oQIDqjQfK/ErHTj6u1/b7iU4ATANVL2XWW5NB
kUL8JeDNJwMVpZnjhRQYbX6nkzgITPgblGgkwNpwcwHhUE35akDsAO2qdyhE2IGE
sLWXUYetenroDxwqUdbsV7za7WQjChDTvF0hafZlKSB1M65CkwMWT761jJUDT6yR
Wiqe0AmkZfk+k6jiLXeJSmn75dUKKnlr5Bpu9N+Fxs7xawTYu39l0aSPzCBveRc6
AvbxnhTVCHMAGNumd5osJcSTjZ5cHsUqNmgv9N4iMh2HOUsNBelgd1mte4vKR1Bp
JPyUvkojjo1xchovOg1++Zvq303P51BjP4FBbDJaomLD9/gbRtv+cPgE9kf1jnCi
dU2K4ZvA+i+i9yeRrNnaLfzXvhfKSBs37m1MjR0yfuGQW20qOT+6XyhM6nloGXAI
SxQ7gdKXirH9Js/P3CaXx+/SEMbhc0WhyuQ2zG3+si8QofyF9iVBpVrVdbcKL23t
azsJq7tuLHUMy1GUHUlSxO4JLz2hnJoMPzBrn8g8ABp3bY4mUC+jryJHhKc9JA0e
hbU3XU+ZD4b3C64HdG7jVaF+pIx6kOvzNJnSgxTkuyoWhs7FhIUSPxz9fAihajkG
ybtRMj8FdVktpUujqElb5ss/x+s4m+HCdHS0NgNN5Oc8CMxRirZQA79Mran2JCVj
JbEgMOUfGXZnk8ISL7htWsTR/A7WUXbQ1EdI3MF9kdCzfhywxTtdJGoL+2im7jk+
lLKsUHgcIXbavmrc1F5tfERru8ENhchli4K31kPjlYSojTKpxRthwY8Klj10evev
PdsjryIecQASrfCvXjUtsbkV/XaQss4RWSTKctlJq/tuKzKcwoC1PChDDHaD3u4c
dpe64F8vsHmhMIVk5/peo2dMlY7j0ZqTn4nPvVnRAr9/6jMOemvyOeaB1h4I1SMg
egzFMtoKZgqRENfiElCMvl6S2fpaqXwmQZKCdDm3DVUg5QJqFz38nCnTlWYl2i95
deykb911NMrha1T+w4A+Bl+raMW/8TpBdIGi7S3K7T49IyRXF7SFfMVLJJA/ojB1
CsTzxFghGd+3ED6x/30mxiTs3gAWbxtyCGCdBKs4kUrZP8VeS3wnr1W+RF4Ao5IW
GxxF4gv/luot5pXu42gMftDKc3YE0nOxN43/MurrGi9mDmRQqcjTyV/7DxtxQaj2
Rbp+HeThDyJoOKXwr88IExKvflr58LrNlNfk+xYPbxBqacvIqUWFdAM8OcO1bQ8+
sy/7alj+XssNC4xHsRTlycwQRRMl3oN2JSDfMLn8/NfrHLzXnS7hthcemibqPAeI
J+scZsoeaxrtqiasiS0dqPjhWxd+a2tfGKKbBMUx7pxkZcb57mR+e9nxLymXrt3B
7h/NQuzKqOd5H6r63PM97iABdl2CqryD8e9Y40bmSLXcfSsS1IeD1xX5N0i71rB2
kGv5hopw750XBEj1h1XM/xl/e3ciLG7T12uBYGMj8W6U72X0hxb8riox0nkTKmPD
I413Q35pE6RF3MkzQDOko5+lxsz4SzFgdIrNLDgI4C7VGSjeIaC+MOiX0Nc1rlxF
ALG/OWWN4mj8k2+e5qCB4Eg3/DYHUxS4cYQDmrrQAB8pbEjhDwtsXxr0DCnhSeEx
ZkXRnlH2oDzS3OFOVwxvgQdUxqn7g8DHFNeC6KvzL/VasxQsaLTiPaxlWRKW3FMV
wIqUTn9xnzeue9GCSKiEh99iVn+9y3v/yoVgVZJGiGZkoZy50DdPQ2UDPe/Rb1y6
xWk70/3+wOEAdcimToH+pz8Y+2hF7Z+ESFlwpv2CH5VoT/8k1LExcMnYn49dlphJ
055oyVP5ueIk4ZRqCJmYRkLrSBPWuOqwP5nS90QqPWAaJt9KUe9y7mXoneuFnhIF
VKffa5WcJFX2eeVtjjAQRROTLQIZyZBYyx3CetqsK8zNp2wxG8/DgEyoyasoiNIT
7XEQAwHFH+P057i8GV2v1XQQw+lYCBKT2ZmaxxxHAhaI4hQ71TN9QpXAEwCxbgfE
Og8ef+3QBDAd3U2IFEDGaFc6DvjTROi4nhUBslG+sMk1U+bLhSYtLtQBwDMUpmdr
rfr8wWVxTilvSVxcpMvv4ZQlyRrwDzQNP7idcX0TJ1b+5eX0Bm2EclyR/1Lq29e+
Im/x/yEvxXnj0pJG4rggaFW94DMvYuYQROQDDvt1Kj9H+MVVMEFTBt6dGJU7i8lp
nlHna26Yy9pdB+OekRuNrlfBOM1zzUN0i5yoGOaoCh/MNJKlv7eqKqWPS9croZQ0
BDYY8Ra8GxQUVB1UorvxXhnfBl4v0YJS2N5RmblZzp7WUsPx46Zuqb0SFODqda3Q
ISyUOw1x2Rw9gecHwWNO4906CRViAmbkEWJi8iiNrEZ2UEnszxWoVRLzqnx6k6Kf
J+Q7EzZekWEkQNUnFdkY8hjvLLcAw5L7vp4Pwlc17hzkNBwFsG6Ays2K+WjXs439
4Ydl+juVwm1fzIzrLlfMdCmlK4KbMbto3K3/g2MJTTJdB/5vncFOtqTy5QARu0tX
6Qv3gNgTlCXV3CZ36nodt6EzzgolyHYcb9aTNafW4sQz/nu3OUNbeABrNIF/PdzR
cYPU/Zp7gOdvms8XXHkD0L/FpOIqiFssEM9u0HEGSTM5MVl2XDcfbsfoO8L5DQfO
lqz5sdMJqxNcSe7tnWSZLxami37zM9bVEzsov5Ge5U7F/Tj1j3lq+QMOGDZUe9eR
OP1yzHwhJA2Kd+q0s8JiBuu0nBHp6S6eOK0IBAgsi6Y0y7h44Vs0D2Q1g/cDblZR
0vJpJS3iyeqJirnkE77LfqY3BOwDPigf+FGVJBjKPjg3BaAlWbWKpG4/t9CiwSo2
usej0qW2Q3k3MaMCZEaUPjW2ci3qz4Pez845ZjpdKAxY4oZYhWfi4DreSnk147lG
HKZquPLQwJfCZHNGRaRPYDvIk+aHnKx/dsvfcwFRPvCbXAUvdWm9hjeVt226b2YD
7c1lIk1qEOej/JV07jlUJCHDyugPxnqRGp2yJd1bmBjkrEttY13Odyd9UNIpE/of
B48Sb0oA8YNnPYRFFE9GOENBkWvS5fEjInsFzlJf6fUJao09N6eFQu6U3YdpnMUN
QLaV1F8/piho8j1F9PctedaC66MDCPCP4NfsySgVrFx0HtNTFj4r49lCrzW04jkn
p1AfuLa3F6crBdcyyra7KeBp+3kCbi7Mj4umBO+DpuH/t92Wyis4FZFOrvafIqqu
o/qcaKSzKOyFTPK62cVxo9sroi/IpL6XkYwvRTXo7OSkfMXIi7cY8qTj4BV5PmY2
QFEH8SIb3gNMS933Hs4bcglaiwb240lbsxDxZXnoOymQTAlyjgo+CJlEzFh1M4lh
rXwUwHHbwlftnrKjxqJnctnGRcW1UWOVmk3k3JhZXV79czUC6iUPYyrAm2Cxrfv3
fa+8BmQ9IFTmG0TcK9QFubtFDPtLJ5VGLhwrRRo6xOc+lUA9JxTPnUuntMx2dI11
/3xJ0JfUCE8BJeeZ1wKNDDGU283aHJTalaPQ7TVqWnwFwNa7qTi4O0+5ibYZ/aiQ
GTwqBiaDN1YjaF6+tSBL7p/ME9PqYG2oldzbgzN4K/mvzm4H2ocb4KFs7LdfT1sQ
3E9XfaOf8Lh8a8QDOGKSn/wNlglr0mgyAzgAV5tKupxJ0DwulonBwXZL23GiDgRa
ylnyn2HOdr+KUu+p7MeGxyfmsOOP0L1pfufmRpWWWCvd1H6RB+pdp5JTvuvy2alk
io+q9iJFYW4eXgpaqH8uMWb3n3269TOb/SqWBK2NY4YIFh0c95y4UZD95ryoWggT
PrlS5jgGH7jvkVuMQkDkHkDEfAYcLeo5MEISjMpZB7/UyuvPKSpvACRPT5LY34yF
sFrL1CEMlPTA2GIMnarn185T5PcKlvuHPJKqw6AkRJQGRjkQqwdsXM5BTW4MPmbe
Cr9deEfgviV7+JZkCXThedNvBvLL7wcYUluEKNmps4sfKOHBwuz1NmrZp2AicFf/
o+0+1i1oyFUqliyBgF+ho5VJvAirYIU27+F3kdPa4ZQ7zwdplIcjsqK/ephTGV8+
KR5An6RZWetJsvIm0yu/QqLj4UR9+6HdYgk0aTI4pi5iXwbqevUBabdHJoFSKqfp
supGjakhTxpQQWMPiqZ58A9XN7Z77UiHzkVLQOEcNbhahs9ZJnuqMf8xhd84xS80
HR/izw22DqJqF6LT+Y1/khtFgsYu9AihMdoNZ7LYJsi3T+2ApcUbL4cxjEcsJZKI
dHocNhTqzjWxOghlVo8eBjo1wv52YfKurPtVIN0XJr3cGGWYfw8ztCh6lNRP5/m6
n70gHuGyZi4NVTLokL8imSiZwHRXo9T9Rarxamx5z3IOoRpwP+8ImzR1XLKbbq/I
5zHO30s/dc+cC/uwU6mHLk8NF/4j+BP+1aOkg76FrHgxE4Wfkt0TO+KE4nWAIJ6Z
rsclH03xJP80/p0fEc8G3rv+qarhT5aSMgxARo9iiamfolYOLWZmWATo2ZqVn4A1
rIEgXQAN6rcWM4LOID4jjr525yhvJKHtD1b6A5rBN/p5qaYt0mOUDJoyN6wPd+I3
ZVONO0S+HAep2EkbJUnYsJlIK/iFxYGqC9eQHpHKOvmDGwZKbzdHaJBNhuGYICas
1AGjuDZijdW4rBnWBMqYG+BU6ltuC77XXgedpPN4VIWISYajOdHjOkh6AYhrVegu
rhyziyQRS9Yhg+vSFYf0ATmBgsCXpRnKcaZYEZSzrTa6lYkTCZy+uvrPsTpgIi9B
copwot6aIf9I/gr5n/AlsOcbPaKhHkjZ0gTBcqKLcgCM/cB0nsBeQjCcLiczx4+g
ssDax/EMF7rmGDSio93faERplsV3QuHCofFRnA2HYD5i3tlgr5Tpex/bbzzLBgVa
Uxs+/SJVr2Ilcv4MhZgkiqee4WtsWEgZpHu5E+0fkQVAq/lebAqJ0m2cfRXd0vzJ
jv3sYMddSGq4PkbenwYzrW86V8M4GcxPoojgCygaKSGkshdXXNeOeLS0FiKuyJae
Ln3Stvuu/ehMWPWmPWV4azutjvbbnXbc6+xsMEEjaa85wLyWz7u9EG4CyCfo0kZI
xdoSFVA9Ai6+NHbnNgUus/vz7CmoIVj5w62OMUQdsXQsK+4dUPsWATOB0skkyG0q
jyVwS4oH+dVABxRW5NVEQudjWi3CxM7uHZXSkr3QzT60w9NjWWbWzpYOW37ntIjk
zvePPI2i/sBnka961JSBGd6o1hSbeuy43fFa2axurRudgp86/wvwxr3RYu/A5h+C
POmIt42QdtyISFyAUrCZ4C5673RDTNfQ1vXEJN4YJqruQoBhHzcr0WXnAybzSeh/
kxcGHQTAzJSlfUSygRVdPYP1+baStm/WWt2EqPOlFNMux739xIGZ6M0cC8Ik4R1L
uuz18WAJAdXTebY2VKuo2HRbJyGC13JYCBDtw5aC/GrwCLo59H3o7bJtCJrAvb5J
xqaJo2zhvT+7HgV3Nc5wpNK01eGaUJ+vFdBb87jyp4iVNIomcRhsC5HuMmoVl+iK
/ul8hBHLxzJWmscqaAUltlaN+ARAT6n5piPH6Wvp8QXLiFCZ9gG1BgpX3Pbl5jWp
7avAItLC+l2aA6XSPNsaGhr3eikeyDThXk0iuQQhP5Tosws+9CXhMFhVZVESTWvH
57sX6s4zbxKSjcfWl2DG7cIpKxkfntsX0dpXsR0Yhl3jdfg57Ui0WUK5AOll7iVz
35YTxd6ubbD4ZWGpkZPm+hEAuRWSZeqc/TwLPFTd5+VNOtYJGZ2KymcTCM/V7aWi
D8S7NXgxTyOwBzqU/9gTy8IQu7YLENG6VT2BbUdeGalhMFcVsBKvVQjMP5DYYx3P
EdV6FSydgxX65W06fAr0SrlR9er0I4rA6cjk0PA6k7IWjEEpkoCcLGOuHlFAbKnv
VgjMMYuR070BIk/ycoM7xZpOAQgIdDKktn79bGm+mYczndJCadPJeQszibM6NNy/
t5QU1UvfUQXLJ24G9CDDlryxL4zfIxoEd/L2WjjQvAwObyATPXfoFccT7Ri/Djke
Ol4B8cQggxt1v9xL1JmIJdv6K7zIerfMAke3ZrUGUSPe71eThf6PYAZMBF8U5N9h
/0ocLTNyl3E0sEFR2+EyTUWRHPtaqJZd/FJLghUHCtWadMZvzpP/aK2EMja3JGrZ
rehTKRLwJVISImDvuLiG31THLWc3ZhRTza2Hwms0sfEZFfoGgMqrqxF8X4KPX04I
ss5ywRZIZTNK6LmfcpzgSkuPh2z9CH9iyjR5fBJL5+VnfOYfnG6+ma7MDkDCnCir
+BkNTIMmQAiisFUjFiFwuWitst5XTQ6qvC2ToOJQ2FwJdOALte8wJkljuLLXmjlr
tZkgUuTtGM11o1dptK8ybPCvgrOGXgXcUQKDLr0BifTpyEq6HFx/uii42l+vFjmd
kzU0F6cgxd7uUoImnAKekNzCPgjuwi11xQ3J1F7p519yS7SWv1BMtCGY+b/mCYVy
g2Bz3Ze1VYpHnAUppHFazOQ/0X2iiDROIaaXn4sdmDMyp6wMBrtLUGPGA0XgP5U3
Kj7ZrBPN1DLjHqsmKNUIA4Pf7gJCiw8kSx0YgKMADse3l9Tc/sUJ44qoAHhajawb
Aqa0vULZ3eSZINIhbmAMMhqd7MK1+JQ0sOmUusyS3t+BhVJian3aiAUV1lEMK3lD
J12QRiSIqDw0mBcZhIzT+5ABMrbBiSRrTSw6KfZ8tgKlwYGtxtCkgqnVlj8VBE/V
lPL5Tmo7bz004Npq+HH4bPd+yh7Uc7TUt3B81ygpiYchAImaTutwXhfTSVTDjfu7
7c37WV0Yd1J4P6Vx1HIi3W7Mvn10k3vpnmJ6OWbq89kmDZDGsH7mQo2KxITup/r+
6BbqNF6gCVLQ7qMfknIchgVBUGWHBVTTVkTDSjLCgjeNRsw56QiunenSY/u8RYIW
RMFtCryvBvLg7owAethoVr2XWNJDS9VRnoj86LW+vaZakDdBGTz/MzDSxnlAusYo
hXSX6LRuqlkZEV42zEr873hqwypzbCIJqeTgw0BYs/Mnc5T7Khm4jWpSOK35686T
/75W9vn9GP2hGBskLnc1kLzn6mW5jmuYwWNd1vs9iZxJ1pHwoeoGeYf+lXONyZN3
4GS38zmVu+FKkl/lg4L/Ncr38E0CP8RynF1y2TgKuDlTJR4gDUNQx8ebhneXho8m
dLeSgrz+aN1YIBlrEK2dmAHuA6guoZ3ANSwnDgYefJLQcsNZVC2/XFr8rJwA87Te
lYuLnvzJuk+ZDJtxOTZ97VWQXcSylmMx/9YeZONb7FlmhmrXYBs1Dob10C6O3s/k
xU1AnVymoqBrJJuvsl+cK3q7tX/vUJuMBmAbTbwXcNfdoBLDxMEL3VwRMkGFHQDe
zTpvbz0SmYtviS+NcVW+36JkYbMnxYoYRJSKdz954xVITSSd7lOP07zaZrPv5s46
3fMHnDKV7Sl+UFZ8v9Zpu7bpd77l8pHdEDTx5PXNvkb1VBOEL3sDzMo9CCQ99wb6
suIAf+QLhF652/qbOIuSR2jPyg8daK8Uh+Z1ARQalopwnU4OVQINbOOG1YNVowJI
zKLeYpzZ/6M3vbi7ICn/NalwKIBlbuRZpMINL3byc0oWS9/+O8AZVKJKALLv83QR
TqPLjKQfHHnB6167k8mZhXMHDruKYpE8NJy7BW1kTAVOUuXrHDELHny8fp1dmhkC
ezZt5krYnzOtL7G/NSzUEvoQjcxY5t05PZECT6vVqsY//jRvQrG09Lqz7nmR7okH
KMJQuRc/NkoJDEJ2cvoiZiuk90kZKhim0YkO6I2jH1paBhAIVHlxIr/bpHNw+Nt7
huo32juWbRlKKbuqs9Izpko6i3Jxz+FmpTmQls+YZnS4qVas2vphYfSlaWFV3W3w
PW/C/1ebR/qbKyQSgBwp/7YKGSA8PUsvUTLfT8UFpgLtU9pnkIfkKCh0ABPHib2I
96hSccPi6ga5FDxPQ7B4SBAOdvWgSRQq1VjP/RLp0WejtHveYjTAyPPPUiFtJkAc
i55qZHA9yUkXd8XbXp3BKnJb8qvH7U688Ha47Bf6QFUXzL9G7r4QA6ft0O2QphUV
rnGfhX47qSBGfVOwFwDZX5VAU0eyuJ1r16B/eC2NSRLMh+nN9i0ILBglDZ4yWsqd
bTQnRY5K09vWACcaPtrTqTCIajEmAy5pn76nHa8bDZIVjyD/+E4Kav6ClomsEODs
znrHCUREgUjkEaC3eWYB06fIOC2RRN44YmiSql6whp+ncq93/YeyErpSJ8gCEOh2
0eo0izKnf/wXbL0+lRsuaUj69X4BuYIiFeXW4AurjXZMQnTssrgWRxwYDUPm467S
JNxdrIrW0uVe+IVUZU1NxYPp/qKfOpsxh8f5kBMeJnKqL+Dfxja8JgPPM9ViA3go
rXNIAkmjX0e4X+V/OLFBTyhyrccT6ccQv/4SDZ+CGpPqN6e6jzmZvMx7E1r8pKYF
jd5uAhEGuZ4G0QrQuDuiZ1nrHVHQmLnyCvdtz0Op3oNKQRB3cI62SkOQx+MeAJ3v
sZePKPc2SKL88IfOgln9UTOL91+RuGddWJ4LD9D/ZifE+LdQuiefrFcgR0EwF1/e
6ql/cDSHcAxR0lClyexTOAwPw9dmKNYxuKZZXezEB4ScIG/bo6i9omidNWmxqSgt
oyNZzENQtiGIqeP2Ms/HAnMwqX7iM3V0TM+KXUtHvutEtnDLv0ex3yvvm1Tw9jTg
vcTxETbshRfynq53KglWwxQxK4BndpbFedwA4JwpV7MyVuwCuxbVMIQfQGYNSPBF
eobphA0OEKTQqofC3MHbKp2wB86ExVI083ZKeQ5LBMa2WmkLXis46RrpnLIEhnZ1
3ZdCJcd+tvbU+GmJCNnIrfL3dPM01lbHGA8D2Bkx9qrfjCp1pMqRIWIBO9L5cA6x
341LpjrVWPgQGezxjm9aBPFOMV0HEW5s/G4CLwEp8HRqD8j56Qz7xk6dCb0zJKwU
xb7TNrKssTyy/JbrXAYXEr40LuUBje6X0HC1+jncppIPWFuduioD2vGVeGIt8Od5
muQXmhcVhsLAZ6MXTsZ0ZZfpFdZlvddhQANTyvNN9LaiSJUwVi2wxcVIMLMm134D
105kgkROa/uADa3gn2fjcAUewkWQuvdpv4jDfGlVv2HSswtDfNJ3kgwbXFBMorpt
LrDQdJh9DfKehyxjJzGxKgHXoaxCrjT/5bBJHaI0rScaadFbu3KS2vw0WQjK5CXI
qi5vZoUQQhYl2LTXVyk+UUbTv1hWobawD9Wgx7D8kGuRucWOghoH0vDfsEPffBdb
VLVYMqnPMo5hAvu/FxNXa99dgo1sOKlhY0LuA/vlBeR+G4718twCGqT2yQusRjA6
BeOGfbdri1cpnl1bpAGEVf+noicu+rUQ3eerBpP0flzgF00G00z6eINwzpRXkCgq
WaA/NLlZSr3fgIMRKojiIAt5MfQVlvsNNVxb1+qlYCRhY04D8zLaNvYwFg9WJMuo
pjgK0Tk2oVsAzLgRNJ309Tol/qTZoVP0kujMFWzUWD/Q4+4LhB4Wekghk2gnrhb7
6fvm7VcEd5iRu29EmIoFdPJ6lznCiy/7D1e5KTKQy0V4TRx6ij5yoxRP38/rCKc9
BZO/OSmHBWVkLWJZBcmqqTWd0LglSuor6N9/f6WStriIgSVX8ZVkUkZtKlLob8w3
1rR+cUcYThttV/cAtYJPAJzZg/bkTI5OA8VK2rpf281jkTfeiuVn8z+X9GSvrPTw
0suns5TKt5ejmMPxkpN5bgyn8lO1oN0txurzwgPmuTqzxvxB8zPuyd9I+zmqtrz2
WtBCmUPa6FSPfPX9RZOaHaN4UCC6mD2GkQaTnLE6XHYdttDSG5rgJO+IILsKqr3W
UI+kanmvxsWT92oK4geXrJPTqlCI3hwjrf0MGuf1vbIGsqcFBf3zU1hYHRCV6aNr
NsvHijcwASfpQKgj7nLhcupg9fCzi5s0eOlO3pDufwaCjDQGFFbAV+OfgHyVfmat
Hwz1s2MhvgOUYSYLXEvaZGX2YtSwNDP6dMA2p33pFYo9kz8grKsbZTOM/PGk6U++
lQsEBUYwoTTQG7LHA1Y+8syHFDrC84de+hL99dEIAHk=
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VXcH6rKxZTXoLBeDI7jo8fKdZSX4iDimPvq++GXw0K5VWoAoYyxb5VRucigO3xnG
qgbOFABFqQqP8HgwrQj3jfeXF9C+Qg9feLOTAEmhe8jL6qVzbh250JGRIjfszGYE
FuND36Qv1XZPPVBtFK0YzKEfG9hpIQGsPG9Z3829bCV6iYWm8qGojVCrXefIzaf4
sKTyMCrWOsScZeeHwBVEtQx0ody1kVyg9kAWQbU+1IECBlJuLpoTVF0ptchAE9iK
brBdL82r+Fjj0humoBRXeIMGlbKv5AGiTSBxzWCvoTZFWrwHZScONh6fEchG66E2
A4/bEybNIn4Iq5l0jBGOWg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5040 )
`pragma protect data_block
8Kkm139nL3HjVXhEg4XqBa6qHFG9uaRqKRbEZCLtRawaRnkVi0BXkfIjj/eysx3j
4aZAvQ+HO+3Cfav01kc0KEZg4+FkplNkH5EO4F1H/OG3uqXCM58QWYBRNTpBU9sZ
ZfRj+Y3Oc7st0yVa4tH5ztgwXB10JLGua8q7R2QI5NYYu+kdPVh4PNax8LOxiT9n
PnyFpkzXsJwFmsTjyoROUbR1xF5nmzqAjkpaONB3qS3iZvWZYCO5CQZ42TKyd+A0
1/nkwa2CKOdxNWBfUIp0RzUwMgaRJio3+62Gagtp4R4+osNFc1fSB8tC7uYTiQpB
GaBsgi8A3FClr02SzXWLeydaqwIGylu+0HBeE7fCtoTbOyB9rU7u/4gHTpw/1O+8
me+DQqQ+0rvg62tNmizEYyCMriAJ9K2kmcDDIWmkbsxHuFX9z4v6JBRPngfmlJys
utRRherBfOitfUe6jN/bcXinFHWjkegvMCKld8Khiu+Yoa46aVM/AroUMy0nmu2l
L/HHeaoaZ3WJWG/1RaYQDwIWmTDsgb/LFjR74GqV2+Ae0nYSW55tEPHrK4b1aQMS
GlRimuj1PVCHzT4XI1O9KvLXxWIcaiF2Knc10bNz+DwVqPipmSAsEYvHL37QBoEy
ZQf6iTwT8R6fouuySgtJV5py/FAoJ2wfxj8Spb4hF/2Cxz5PBtaEmlxg0KOWXf+M
pvWjMysYlQryYmcH4zhNGWsSFxYoS584O8Ya3FMjq+Ta+jf+0b+K8VU+D8fp7KDB
0sFTs2Ak1QKGIY4kb4KSz7pm4C2o4n96U+fIciyASLuMSLbwtnaiQW68KkdGNpV3
KwL5x3MHyM+MLP7rzmTS49sV2EYJhybUAybG9dPaNIbLUzxgc5pQT9u0fE7BdggJ
hlouE+VZPnDXt97/TKtCu22t1WMrhtAPmf7lYz1MUklnQdjHFtfh5QkOWmkKUpvw
owOCQMcj8Mwp3QLYUI1Oaw+Xn3qJ8tMp9/B0MvPnob4Co8+4tMUAhxDdzKUaTy0Z
Yr3bfU+Fswrn7JT2P8n9Abh8BwvdzckgeEnPvBcvTltb3FvD36HHLQpqmnXLVbVV
rb1BElWjPMjZwGaG5e6/sbq8qnJKSSlvCIcTsCMY88cifit/QbI4Z275I3WaPzgU
FU2bsd2xVtD7pw69uGt+pZrHhYYdpGN4g1MNv0/PYF5PpDzoWTKDfkusMYQMhfHR
ku9pijGqWcn2a6hThL8/a6I8P4FmUCQrYgnqKdww9A6d2VNd7/kWtdpEIS54EggN
sGY7Xe2Uq6toeer/hEDPIuSsxo/m/lI2jNoPkTm4N7hNmrK5oB0kOm+XOQAK9jCW
HzuAhmCYx8m9dnAZHBAursOWMXrJrv4l0NxtLEzCEBNQw+pO+ELLsj5oGFRPMwAc
dnpkyUoZcNw7DT5kdXAp8mcmTmGpFNrn9D0IXCn6rehUK164A+Nk88KPa5MC7g14
E5UwqvWLhRdy3r1k1EeQZIGpM5GV7bbrT1ts9dmYRM3Fds8mNlNZ+OwbUK2bQoDO
wjn5J7J3zPV7acRoM2v/QtUD2g+pyg3PCpohkA+tZtD/TMhzJiYHmYaVgm3xHLWQ
oRTyCwRQG6IpkEd7kjhG3F2Zg/MJA6r0GJ05eOCMG+SWyPVDwuPuH5u/mJ/AHzdg
9qF+1Wets+VzwblMRfC5Ple36tG5asghAClCyYyHyNuHR/LefmO6i8mQzQ8GdUXX
yDpgopPkC8SbjYN3Hp47wOi3iTAYBdUD/Eb/ZQHOY8pUdappDy4kjKRzi/X768NN
wtFe4H2WeLWqEtoRymKx0Tp1aoU+WNtODDQnCwqGdbfNFBe7422vyOK6ABWiJi7e
jFwfBgyqG20NRujnNSrvp5suAEbH864JF+YtCJOK0jcrMUOgZb4eBrFQzGB4IYaK
Oe94Mn6alxEvLbgoBjGpXOzWg6LL8w6mUfX1pzMzX5Ib9C3aQq9dBG9oEk5Eq078
73wObHRLw+d4qW2BwpPBmPqjUGRzjDcpGJlKAzHAhy2n7BjErQLzbW0HxTIbL+Qn
s7/UU5fKUR8KcPb5cm8FWOGGcU5TrVy9pY7i34hyQlvO/EkJifmCXkJOIj+Nknsu
fRePSHol0TjsyOBpcoTTjevtwLwqdy3v5OLxZXNz34N+KnFnPU2ILcDrFq7lRtr4
iadKOM5NflJpX8JmFuVTZl2HiU72ekP8j4s8yxBI1kM3mwLs0q53EPzvka/NU9RW
jI1IGOx+JYQPURIdqe/1XIqoMJ0/qsUT5AydbrY4LpnamaKZPCqF72lqaFzo/cWa
lRBXq+DprEc2XdYzoVJnDTV0yCOo6qgLkEjzhxxDkfXzemTt+2DvClmy9FYBYya3
IC7bvb6OfIGid+0cJPwyN3SI1E1VU1dCq6yC6TjJr+N5SzlJzSRU+d6kcx38A4wN
oaVKKSO71/PFuEduT+qFjciHeFG5QsGwJ0wxCxoOMvc3A6TCVARzuKYz0Fte8Hx1
hTqDY9KGdj9yQ0ASrON59tUgUbKMt6mlUfjSbbvhZWrUeP9vu32/mkAzYwm+Bylx
YGKv061iIJeMpv+C7HFBdb+4QE2qBbjdJUQt+CFpAU2EwkQexMyyOoVQgnxpVsyo
Ai30qEFSEgEVYbVrZyCTmIhPC6lp4jaD4wH62KaOOPg3o+K2yQ6qz2K1NG6olDq2
Dlxk25kx/eHKl2go95IqlelcqgrBhLlFVQia5kPXktIx4gvCLiacslKaY1vPX0qQ
cXtYVJBxibdagGAeYfigvIYDtTsV8B6CJhF+XZr/GI/aWDljLlk5DyzijLH9Mzcz
0r0l/qe0V+et1IwV+F1VS5cjrL6G/+FtOX27Bp/NcBnSVWRBv0ZE4fAb0xi6sFj9
MHbucXitCFy+UVf9nSU3UsH/X6cpVUzIH+AgEI/CjabF4LOmXeTPHewSWYiolfF2
0Cxfty0pSG9MQ5dDt32DHLOXJ1Hu7b1XtRWATHSyP+9ZUeTh8b4rHSEv4kwCAa8X
CYaQgXeB0uL0TqzrzIe461+fOU65rF0vpsO0bZhn2HXfWWxVzaritQQ4gGzJJxXm
rOpEFU2vhPC3Mdw0+3wUAqrkPju9tMlcxRvJAxZAVnCcLtB4AnctVqHKZ1hTF017
xUln2LHqsQWFtqO+lxZNFC+XYeg0qmURsrHzyFG93aTAANFUqus6VWTWbzA9G4D8
ohoCkoftynFXoHtqeTEoREiA0RhOHNoopEuEnksUT1icu/s7DlHvE2aEvLFWAbIc
NAOpipFDRdqVUOOhKR3owvcNRwfCprdigFMkWnuZqeBRoEyJUJ1Iem2c05ltoPAF
vxecxdyw//k5YuMZHPczpRHDlN+4bZCjfhy24Iz5woTWrZRdAVHL3e9hoMTI1YDz
+EQI6S8AbR/XktAcXxc58QjW5O9iGq/UVs6gXL9VAE+2bWp7Fto0pm33Dffns9qd
WKt//WqU6eVFKPLPSCxzT1iKZjGp+3lURCFeSzsmMVDByQmvsvjGGd0L7bo8mpOM
iR1Ty2x4okQ0w+Ki+NlNNupJ+Vw4oQPLZF/8076PxBc3WbPVGxnLSB957oV+yAGB
DhV7+v3UY/mC2J+Debycy2D9lK5qtK+v7Boqsmteq0GemgCDduIZso3mah6Kgpj/
mIAF/IpI/IM37Z04ouYkyROY1rbajqrPsBFVD1kZYGpfBM6jWOvKzksyUaEcIvnM
d+K9Ne4qbJFGpy636tW/BlEhVP6fqHhpJyqIDpRt+/eE1YequFccQhnKR8TXO3YG
6rCQOuQcYvanfFaUR/2cH28bEBYBpj+jyAJ9znT5ys1zLgZNYvhZG+3hg885YEti
Ns+uN8dZBlarAXSpru/YVxkftJsExM7w9W+wb4QNxNrIBEyv3KyIZAn1h4Ltfr0k
ncPZ1NJnDiBnM2sg23FyiRXRPsKUNZgXk+e0QHkLDqeAM7VNBScXlM+zr14n8BPD
72tS391fnk0CJoM2x7VsrPgqIzfcOnlnKRjGnrLPnvPF6dhUBRAKfu8bPbOhH9TY
ENkuduyP/xGPg4+lDbR1fxfjBZ3Xhi77jNdoiUkRBWwRt9M+uDt1ZanyYZPisZT+
pHxSzInNJLnPTtQTaIF8dwbqyQSdqHlVnnjZoiphI4wvOe3lBhh5ewg1jASpCyVd
C2CBOcZc/iqlEKlhSov6kQiSCljO+4L53Zr5ajIelIoA6Uf6IK+XrcN3S96NauxZ
DEvc+wDkWGynbKu1oNQ7wJh6lqW70r818Vl8LbeYSG9KC8KAEDLJPzXC6NiBgVMb
gudwCntoUuCMStqdLqG6DDmiDPWiTk3zl17VaJYQsyHg6tDEyUK8O6GHrlajMntB
2tdYgb0YU7l+0G0xM5rHs5jChRSdlK5d43MBFmQpdSFYJwTUGf3n+pSMzoEJ6C67
p8qp1PIY5tqXvvO3Xh74wokMm+IlvnnwwOJYKkR3XEem5ZxCzgqafb9XwrOBUnSm
OgCaJhJSc+gh+LO6wUJJp3j93F8D8CV0prZjhaQnCikIN4o+x3iPdEDhjisoIiRo
4jMLSpkZyCqR/MELqkcHkqvmo9azqsZCEkeKdi+SfkTa6XYK0+z7iW/D32fF+ZLv
1biIfldJkraWNFoQi7nM9JZAUUnfkWocfvGIkBbeJg4najtefsdsDl8MropF6zYr
8fgTFY/4Rcqd3U28sRqus6a3h9A6u9rSbfRWfFFEjBB+ybTfiisKX7i08DHCMu3e
AAUImu/rfc9Pd1j2cn/qqGmaFtWW/LRniq/GpZHlKD/qJCe6foYBXF+gWh+0FpuY
ahbfjMFWJDhtcZ+N2QGqIEHhqb0xxHOmny1eONP/MUszERTYCRKaXs/7fOcPmCOi
goSJSQ7xEZrYlxVPWkcqUtz7lspgdWNepZjMmU3kk5XXp+EHqlv1qn/aQHfIJxT6
mKckuR1WN39QE/kIu62aGiGta1H8ch84upjeYjaBI9Yr4OWszXifpa0lZzu9MdCH
Ds1c/tUoPVXalO5kFYGZy0W4aEIF6V9xmzoW4gdlPPz+jz1n6rfPdTLgmCjEpyOS
Q1xKj8BvP+ES76lxJbOjPWWx/8tFC8pil5QNZQHq0Wzgz0yl6XvVaHNiD2RqvgYg
ciQiMJ3zjVMjhB1w6fUgQo5FVqVSgC6zJStP9SUYro1dMiXEWzc107yb3znIH/IZ
31dnWs2aTiXZsAjHIlZmCxHAVdKXgvb7o3xsqfL8qrCHYQCY2uOBDtPDbUnOT5A+
9A6HQYMJptju8nMUEaobgt+rHTJpePlYoRSdJXgDdwqKuS84i7FmILuzyPEaK6ai
Ya3Bsj86f5D90O1fL9RZnRAlM/YMpHhYMX2H6872PsxfuOfe5wkXy+QgWCLmW/OW
XItDkQdgFRNkXS3W/P4/Q10BJJ12oVCq5239q8wYEZKrF0h9ZM/nTlTl6D/AJOvZ
HfwQo9xaRcOIStaGb6LAB85GOUKsUQIn7jtdnLuDJXZ71Xe/E02b01ubKYeF9XwB
LogpWfPbCJ0kpdIxjGhvVpZGTwTjemde3L5PypIcojwzMCnDyiC7fbFXA8VD8FT+
nukG5w3Q6HBwUVXAEhn06gFzAVNhN3rssq38CvlzbBZPX3XrZ0Bi8ZqTrFcbMG7P
1isMokQQ5Obh6ZQXpPMhI4fTKl4gK6A0mYwphO6aUV6tWz0QRZvKb857w3NhHV5a
RxQ57nZW0Ho7majud6kDd8DjjG7emmr+DJ2OB2r6WuxoIy1IUjIp2VRmLGNUjir+
23/Q1SIClB0Zi0bdVeQ1H+55wUvbhanO/l540LQyAqGfon6uGRAG1mUg4ivPL9Zw
PvOxP3QIf9/Cb5uYvmEhJpgwrAwjUXXNukMAp7XM0PWAjfrmqk0lTTeFTm4OKWPt
rO9Q0ynKygt8d5niDarebiiQfiMfSg2Uu7Bi4OiLNGvNKoC5M206Wbx5zyi6H8ak
huyYTieWua+EZaCuspnHgxKNvCpNfqH57FKnCWChWi3LHdVSqUIDFcWf/sU8Guxt
HThQ/jVeG/dzhj5bOQjQNu8P/V0lxELOzklcynAmojy+tdKhoVkAmUrQaRYUk5oJ
OdjZBxAFudCJ+kbjmnQBG0NfV5WN8rbyQs/+4bEuK6+wmgKy4cB/TegpCA5f89Fk
qfTbFqo8zkd9dPWVCObWUhM7ZILLiTwEwvTbGRxxGBPCt4rc298LR6htjjRuKnwr
kqTJ7hjkhegG8r5iJuSY+vwCaA58PBiN4TPYgHZeJ7Px9wuBILT8EEjcNoHZR2zq
WPkKV8wibt641n++R13xDHnJXGJ+gbI3JwPlAet8v2ifxobIBBK09yVEDr7FmSaM
enEik6eSHYlLpyPhDxT5gFWlaCStvGmrrMkhI+n6TGUNFCOT6wEsF4PL0LLPYRbS
L7RDTYmbV5TUuq6ivIGxyDz16f5W3Qcu1c4IrhzYlOgRIvHu+GUnFpo9l0cjojrN
GkRZM0TpxwO6iRm7Yq/E93TUtPtstixn1PSw2ibe6WVqrXcGmA7LPbjdsBrtDPhZ
mRFkHGPlqdTxEghnTYnRUL9FCIyEMe9QzYbGfMmL3izXcEMW+y9/Jw/6DSXNgT1q
ExKuuuRGE4P5zhFISLQAo8miUxz8Rpdbob9+ILWwRBlU+78vkdE8buG9xIgTKGma
sITuJ3HkMhIAfCZcUWEz+YHhfSo/LvLYJ3drw9XRtpq7MnBBK10xBow8xd78TQaa
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
h6wwNYUl4GA4pRXuCfkZTjH0RoQ6CVSGafwqELDWjOkcPT9BS6JPU5NVwWKgywug
qzRsnIkNBtaY2FJ5l1Sqa/jv4zzPj7w6NGdF7b2j9SN44fr6EAGh9Cy/Ul8F/zev
613qbsuZihxNIgnK9rrF0ZF1bixtcK9Lup5k95IXTOT5SQVUKnGcME0WeJvW/VI9
t4qmkmpzCoJnM1soOhh3dl01jpLjCAC8c4BXjPvDBbbviCzsT68JBxD1uopGV8Pn
DBOaz+wgKwlzsJWGuubp33l/A1inVyuheuGg0tYvo8C7cssCT+izvCrsfj7mNWQH
R20HF0IoRQwraNXpy1cpUw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1072 )
`pragma protect data_block
S+wZQd3n36/d1tZAoSjedV6MMArkEoYbc5HRwbY1ushntbGOgImho5gbSVDGRapV
HCj0N0BIOMc0yUVF41WWObBi1fNIIKK2RPRUCuHBS0wrHefDJCRhHSLi6gIG2oSq
K0sF6D075LC43oJYlnQ16uNSJLGdDpvWwzRpUc7asPHq8uwNWaHT6iWaZijh4zgs
919MBY/W2liRylyYZuCDwIl2k/Z3ZecSIrk2mUptm+sdvh0ojVxlb7u7/JADRn5w
/wjM0utFxTO7/d0EPBtzES0bpEMejkBEyHCFvcDdrTXQ2Tq1C5WeKqmyRb5izOak
rfKXOX3Cc6XzHIT7auM82/GyNMuDnCghrNYUBnvs9wjc6MYXIsOK9t7N8Y85VDbm
gvdQpIQFN41YIX2ImouSIF924rY/76XUDkPojqtoT9OX4KbxRpEiVo8g1vTG9ZoD
m+WmhQTOQJl9gRZ7fJkOfEJEOWBH5I1nu4vIgeHURg9pwjoQQkrgAurGiFZW2sSu
J19XW24bwn8ByPbAi5nR8DhH6lvRvciOyhrM09CR8mn6I/7nbgHgJeeT6vWgQOPR
DYUqATsm9QuzntzoEeummaiuhkJ7JMMYCCH2a3U8ZsbqHDTSdrExbWdJWIVutv0u
xUNVkI0U52Acr3+JgwoKI0Fx8ysVQB8DjGF1O7Sniycg7BkvglgO+VByZ9riJ4rE
aXFRD3NJ0V2mrUyQlb+wqLsMsKTbtcL8pm4xuOrj2+O6awXEDBhhMKVhAUehGXC+
GU68wtx0mEpjMxt9eRJc6uRaJgtv5WarpoQJqEggv/hPDtP70+X3kH55I02QnR+j
066M/GLc7vwdMO0mGaZQmTpaTkjoCPm7/LyN7ZVg1nmjeN2EvKsj5RDtnV1iCd5x
Sx5zs6fkZHWd2V0X4lwsLfJ2KmUDU6Pr/Ts2X+gY6lNsStCepys+r+BYOIBZ3qvs
3zfHzPeoMGjpuHnD4ntVYG5M2x9M42T5naK/1JB8AAurnOd4UnWiQsE03ZD7j7RC
6i3zykikbM1CMidhAvkIjGnJFI8Fh6YZIgracSCUJw9cOKw4K3SK/dZiz7nxpqjd
ZwkOf5yIiNKvxbvd1u5paUy+R+NyuOxOcMMNbZD+9cwWZKLXUaBMQKSbDCAebdK+
NfZ1T6TS/Q/k22OwR4E7++leocpgJ8dqww9XCOEv6ka5izsCpihG8zqx8F3sg9lN
SLegQgpgS88S//jCH223k8xEHmDvU3NnFfokglme7lm9bhZaowFfyZTELX0QWEYy
9HanI8oNC3RvbF8wdpq35QxLZyM+hKwddUG2+pC7zY81hEO6DD5oRoFEhuxqgdej
YadG67+YkjA1l/wDjb+cvV3bwEFDcjugG3VLfHigBR01VPomajdiyQ209bh2+Jb1
wzgnSkVINML9hpYv02McbA==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JUgIwFdSaeex1d6OdxT4IXQc4jQG9SB7GqNv088n/sczsV10XmStLF/pIkeOEMmj
sKHfQqXhE27OIfqibvTn0TsG9xb5Ul6K8o3i5bphxYpL1krzEp302l4b0CBpz+wL
kwEuqdA3QHA+l32wFxCHzK8+RdP69XcjdrdnZfmglpZqtHULndpKGF21t8TCDvBj
hyhj879jPjNzTy9F2d+dzsxdtzc0N29koA60MUrMUQLHp7MUZxdCwSHPC/PPD51T
Tt1SYFUXFiq2XBzON5SFIoCghfQuA5xwMNzPR1faL+UWmsBmU2kRGbm59zz/xmeX
QXEMrQuMlP/FgilHO1n5/Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 784 )
`pragma protect data_block
oHMWN62mZd9kO2O5b643YPO/LDrwlVhFkLwAtctalDEeG93NwMoHfUtW/SulZ+U5
jnWBlYu7/5ePaBCuWrHPYOJ+7nsb9ZKlhltNEh4dnNx5Vxju+ax8LIRhUlzLrJC0
XV1FhPGo6CT3kWeq5LHKcnTvjyRvb5WBjSF9JG4I6+P1ONyM0VfBOtZ7DNUyIiOE
HYT3yeFdcNapaT6nESc9QP304hNQu/LDV5RGKXHSHdBVPydb8CdsyV9sWNtN75Du
FvNDLwSU4aePHnVtQIhD6Er06BWCUs0wqiaiQjZaeR1a1ept5Rk+mHTjuBSSzx8K
aMPCi6OxCWeHG99BKAVdgywZJk400issZS66Yr25l/Tkd/+IeQ1JgQTU7iB+N2b0
RJXsrZiCXB2K708HLid0vNQtgE8a2j5Sf5SlxKYQYyF+tahmokyYTYvmlzIHTKdp
LSS6YKJva5BLLPIcMUnCq8hkMQIenE5LZiopTk0v19IQTvdJyNioiADK4yj+aqw6
k/egXpNgfscXmd/++lT9R52FRCdcHYXnRN8OPORphzr5tLM0tTs4yrkQvQpZH9mE
iERuYNEItN4b0HcpVC2AUT58SlNu/BL6+5HoCuFL+IBkX0szOzSj6zFRIGmqpnss
Y6gEwUyOt6cx42TDzii/u3FF093MWLK31BjhP8KC2TuV3mJs8L9c50MBagy4/5fF
LpdTj5Nu/XdsO1J9VQKADTA3JfxlXjGZUKHe5ynZj3Bg90wf/bpc5cryFgLwCfrO
TsjbhMDiFcqaCu1Nem+X+RxGpoTCQnp+MRVTeWvrysve5fATddCDmR3eBg7L5qzC
GqckQl+OQNJKl5LJqU/qDIhsyRuSTfaxO++lFSn7/HPkPPizE+EeOloWb3L1bAlm
APD/1d2KzuaS85YdBCPeXENYxiOTtyY+ZEidDLDjtdWbtOckyvSE+HFuDfyBxhRA
EF9Spm7OBmWNbo76EdARypmyifDtFFSVQngE5qvDolsbTh5Sz92SjwVEI5abGH0f
xW7xk0ibqHno9rL0k8CpjA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
OftXhhnW+hptdd+Br5NCjMFdtWrogjPQJEgjQzaY7LtUg3GWgK/FoqD6PATlPqrN
KA30oD11G8KU/MzsQnt06neLvrGjVAvgR7yfghLhHyUtxZBIysMUKL3B3/vGONlc
aoSUUqUEHFGsPBfXJp0qK3O3Hnr0GmJA1EqZZKNM95cnfgDBaJYjt/7NCd2F17EU
7JGcc1+vsJQuAEl4nJtS3PGJ7N9NZjwnr9TPzkVEK5vs9J9u8fxRebBwlHBnFART
zuL3NIWcfyIeNKdVOF61QXeX7snEnPXcfUIRY+JsLJovZZ5aCt5JkppTAXtuC6Vh
QIs2pESrtxVSIILeEra7aA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
3Tim9daniU2Xs7NzwYHD8sUScTYiYmDgMJ1RDgXqRhyfQ+tVwmT+vCb0yf/zq+aL
BBXdMrU9vye3+soYimTV1++TmIsfFu307FrHHA/FxKQpIR7k+2fVhP6M6dSFofae
M5gUPf7OdoITUL+pSB2nO3MyCe+rusV+XRcyqOKLGjLUiDqBOay0gH3AUnSiI4et
k+6qhTXtYgc1CrO1vpRv3V5FzJi+JgkDsUzTip/NLCsgifUQ4NkOhVJpSFLIShKi
AidOl76yqmAEPlVom5IOJjOPIddC5QccCuG26OeURpIFMx4DwKbRGh6z9Wuz6VjV
mhoh3GGPGin7B/WXih2IjX2wfzclOOzrL7p0szE4Ea67w+WIudblO877DnH70IoR
W/0Y8Fzm7/pBQxRiGv+B2z2N90bZtWunv5pCQWIc+urvIJsO4tH2uSnnhrL0+Efn
lxwpzBFnLrNosaw3TcucjbA8g1TybaWTjF/7tGCXF4lpV+YMiOXHLrwe8DXgDv0U
hp3+y3PvtS9KHKYg37QjocoBPZYLDwLMZhR9OgvsUqmQGb+5ITNrOho5AIzNQRPV
Zmfll2HusPKpt8Z9pHNUvPx4HSCOnz1iYpj9/xRdxMm610U7VDj6O3iw+Mh4GHhX
/KvS3KQaIatPrFfSYPs+MCDc4VkZMpTROK9E4dULjmm7z4T0fwExWnGO387gJ1qu
bVsAWe/qLcwuwXg+Yb17eecjbg6FKsCpZVi+PeHfCqkcCc/98LCGS01guXoSb0sm
x6Mflr057lFIMfvDwW5zNc2glNsJwKDbWKl3FuDNqf1d35Tuwn9UTVJoPhzDNBX1
HbhWMW7ZnFa0N8EvknMF4VurWL2RtYvjaSCP5Uzymj8HuuHLdT85beltT0SQSNqI
C6rAXuPM7gXOU5nezqQURnGU3dklJ7eiiLK9G1VcfS4=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bw5LYJ/F+kWktn3O/Rblf26Gf9PeUXRlMWoCyNclaFj4lQEbIZ6Lq+xOt02enDJQ
9HbwvyaqSSmugept+k/0G6glEAooqCLELRQcqIW3cdt64ZaEPe2P6cVA9KHqevk1
kvjhpkptNard32w6RDmPZQ6Z2YfSFbC/NUsAV7xWqWUO77WSJULrpaT2/a4eaQEQ
JrVlulXOev0sRNQO24fAvCFUIwJDg0kXZR/K0NLZsDkRseVZaW92c1rK2IWcpZKp
BsGTlywXEQGU0VIYx9AeHzTu+n1WcEvKw7UyggDVgTrPg4xE2iiZ8YwWVxTmTN4j
DMqqvvXScorSd60U+7dyAA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1792 )
`pragma protect data_block
ay5sl+l+vtejGBNeRlRO7t6YCvTKalaCzAs3glUp0N1HvzwR7RO/UbF3fcSQ2lNZ
Wmq4YXCnFlUqEbG4tOk+L/C8vRsrA4qbBtpKEQvH5LvPLzPoogIfJHVH9txYmG4Q
Q+PqW51SgObHUfT8eldENPK97tJ9P/V0i4Su1gjgVdv3VHxjuYo//PhwOh2RjESN
EzPR8Tzh+tAUoy4ov+WQAonZnKeXM39fZMtHlEigpYqshsxVxrOI9I7hKv4ermub
z6wbosH9oZ4hcdQGiGDFue8uaI4lQP4NooCgHqGCeFVSZuZ3zJURAPFSmVx0vHUt
i6nE0tp9DCLdZzKaViISqlTEqorkqrYoTTTo+Mhd3XQLw9hUeL1aGLG5ZgsEMzOe
dPP7aFePVCHvDYmJN2cC0hOc420pxwtuzcBB4v+0pzY2JKzlVavM9pio0JlKYTX4
K8CGKJll/QA4pg5JljrgJioaInnVd9THZhyLAond++E/9y8NqRAvwOq7YnaNSN85
O3PUXycB1t+dysPo86XVvZFMAMB86jY71eHMzPElvWOjZeGFOBS8lbrZrFvtQUJK
m5cwFN+HZ/vt0Ggz/NyFMthz5gC6t6m7IrybDdBxXYK0KHGpn1I6pDI1qaD0/lNR
QGI5HLhHf8nGscTGQJgMZQHYdbaPTFYkrPBEZyq36PbeiAwOBGVygKHfbRqkjDuL
G9pJlZBZNplo15HIumw3Wb9QNurT4RUHjG0DPt2RjtjbutbrdvgHLj7zqv7hjbV6
b5QHF3UEsnSRZ57+w8TsN7Xu2cBll+uvEbBcyFbUBWfYHSuOr5pcFJJ8MWudFtrp
+TTl1L6Ry5eln0FYbHhBaiG+Cp2Zn0txh8pqzV8PTksRo2AZw8mnq/EgHKOUQeUo
whJ7KFXVefkbAllrF87E+FU4eqPBQsIZNgwpGNXXCKVBTv6O2eiLfHC0mZIt4/2w
2E9MiYCMKiLaq89K//HB64sOHppC5q9oUmPD2JuRumXoqk0GqHDabiGd1FkO0ZVK
pzojLHkNptSmdqBLQK3RxU2tv2K+MemmXe+/AUDn2kQWJdvQeOK172I02P5UJLIo
ch55h6Pmminxd9ZY769b/hR7ROgS54xPHBFXik6Aq7/yox0kFwfdxa02v7I0q8nL
Mjz0Kp9K+C2Qu4U1KtiNmTtZFmvQzKjUCpG3MRrZMCNgJDlFvy726RvzA7Q7aYIf
VIkJBYGomAzUyYufx+1R+nOlwltd4B6gkxN3pGQM8DL0960GVls8iawHWRN+tGZR
EXW7UBDyLubvDp3W1LpnA3OKf4BKmPGM+SjFqKBEJ7mkn0KuhI8gu1sdHcPzXefe
+zERC0fr9/Qdo4O7WEZlaD6zzaKykc4wYCRhGDCPSqnZE2O5aIB34FZAWv8HCW1z
xenahDGGjGlg3H9UIFBHmbpwxYIMvAvYCsYQUa5IaHgUUERKj+h671QkZvsuR5/u
PuEU1KbjoGbof/kzZVLJ3iLjMPSoYXxLsJCl6U02FDV+GeRJeT51qElg5Gv4v3yW
X/Eri/t+K2uvJOzUbNLMy0b2j2oFsU61Pd+DoxIyRighPzcrbVd6l8QHHEj4WNpZ
WYVDjC/BPOc7bAMzB6qkxqNOAcDqpC0/ziCCddw2jL9RptWbYXFKcxyaV16ekX4E
7xVw2j1/saRcAxXIKH/F2D6b1Yr4TcQabAlRuIiQsoul9Ewj2jjtU/o8hTAaLfV0
UR04arLBq6mzd+wa/sKmLb3P0vjD6+L7mD/MHo4c0ob2QaUQileX5120XlBXwrla
VFnF7LRywt2H8lF+JFdN66KLjNMN16BVLGdrbJHwzgUaYs7FR4EJoBHMa4gt0Pvp
TbWyah+Ops0fslgQoqAFkDihWbmjz9wWvk8e7JOZpvgv2cmsUyOPUCtofgT2yx6C
ohwmR1lWWsTxMvhpgNK2wM7qUXFtZUdnwqyi3nUnBMrnqrbikhHspAczj+EdU5+H
4tXvxGuxdRTpkSDJn5eTOZ6G9PqNq5lCnPhZQY676suY3y5n3yc2JQMDriBoJ4H0
aFj33ockwhaMOCT4fsZlc8HoGuiWESRQnp6RStlYQfLfhP6BNsN1aAi1zgaXB6MQ
E2WTcvm470rqjOhkaKNAfz037vCyDdetd3P5BmSsfXsMeSONA7MkMELvnfqGc62d
PzG8U0/tF2y/QP2VVl5ijFx/R61CXu6uFjqthHyG5YSE0ZyzDBoPFyXX7mohB8aE
MB9tJkzsiuGZz4a0khJgJQSpDLp0k9xeMxARTPWKYTCquDWDdn19veNM4FIMgZ25
wyzNmRTGTFZxQ1b9ieYxKqZ1DmrWW4bA9Erndsk4BziAYk2hPfh1144pnyA5+hgJ
d032nUQdCJSJKhyp+dspNA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Z/Sa97QG1s7xdsEHm+/d4YUaqzuvMdkQspW76pycOAdsXCbeo/0SNmtTX0NvoZv2
PcohjPeTCLAW2VOkXRW0sO0HYvxnrF4E43qz/iuDgoB5HQZ14FLoqvoVRO46kgX6
Flcpf44oBKkQB4YG0zGM8a/mgzY3G8EJZeLw0yvULLVc8XFW+79+Z+xaHscuj4UM
kUABVV2G6Mc98y+TdLu/wHsY2rKadSSd8gIw6lEaz1DbuIEapFU7gIWXcbtDYmqP
qKuESfcIBKPxI0cjJivKJJnYTtXc8KT8CB/zdluOrEr5MDeMOSYRQ7SkRHiHMZ0T
4HYF87AkYz0+sCuSpN958w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 38464 )
`pragma protect data_block
LbNnT0wgS0LN9kkMAAROGHSFgjoa/H5C6mbBC/3cuZgAdP3xbFSfb7/9iMt4iZCH
y+KW5ZeW4ubbykQCZn0HA/nvWHHyLCU96qUcTAkp4VlJ45uPWAvRy+Hg/cDaJcck
RhAkOiNslUjdHnqgfgW+VVsPN9hqVA88bsuaX9KTTjBz9ZC4DgnfSLkwl1R2Iajy
PStirPE1rnft+SpZZQRY0VIlqdqCWkK9mLJ6NO0i53z3HiuKnZK+Vs3UR0ldCz/f
+LPyaVnPZDUd22JG1hF1Id7zh2p+1pcoZx4Pj5D8ZkzDc6/iWy82l9o6mZtv2c/g
uS5O8Mn7pOw6In9wersHXGLAnwCxb15jEHlHmDi3RFkaZ/d7fOgWMGqcC3bBPzyC
vbQsCa38n5z1guo6ESxVD036RTWaqpVSs3xfChT1G9YXqt0tij3IAow6c7jgqZqL
3svHau+2yzqlr7r/IGInjC6rkQX7usgXkfS/S1qvEPL/yKsltrOb2k/WUMbxXXTv
V0gp6Rfk1Y+AswQZ7T0POeu+3vOXJiPx2Kz/SkNiJE2KYg2cQTJBImNJaCQONxHS
ki3qs0zs8XCar+2LHjz/ziMWsafiDAtkEf/TKfQdYwcS7QGv+e5HtzjVRMNrkFNZ
TC+CXZQmtlmCJkHCMnsglWdN6KCXcWhYttL5AtL2R/Ez8rdykWvhg1yZv4olBd//
KPGQaC1llaSWbdG8V0Fvvy7hZYwBSWayhp0uW/W5yVbUTItJ0pXcRdqzjxo2yaOl
GslYjTNVepnMcS5gnMqy4cAdWugJFgtpUtx7lH8UDgckzB+1KNRZgir3sY4cxpsR
gdcnLxMYGaF/Y8rs2weagOePu3ClO338sN1i8bUulRCWpWBLamk4izRGnMCHciNd
5dRggnLrYH7jcK+0pvXVLy6bCeIqZneSCl2mnC5LcwF/XfWbeKySihKydy0RlkM9
pMAUsM8/bokflPUvxUSxoNiQ+mUN8H3c5U7/PkNteTvsua1+qziQTqbwL2euTwiY
LJTiTFPMk0S4f+Ma9kCxL1KNIQhJwviNCAhilbmj8QKmHCCBiy0TCEm/fQg+ivIg
R0JxWvaM/VJmXnft9DDaJIstPtv8BxUpMULlZeSgxApoibY/DxqnPa8IDlIL8VzG
Sf/4tClLzZk+g8kAuGa+isDqzPKgpUVDP4zkQxeTi+WDCuluMCBqVVXsLNcFrkq8
61BHE0Cn6FjAW2tC63bpx6xN4XzSRsBABdG3mNOUlLRw2XK1xhsXK6j9mVRkb5Pz
SVBZThbSwoU2rFuJ7eSOxbOZHoUGhN3lAhALDAUM2v/f6YOrEfFbd9V9PDeFv/kJ
3DP20m0KKvK2VuJY2LKhlZ5aBXfAmTzgD/WSR6WbGZynmGfjhajdItbfG5Pa/xfd
f+lLiPawKh9+PENzNfjOemwZZgg3sy+KhyMHhwREdTXi9Aab0OnAHtvdCvJBlxFr
vjwvDBcNYmCdCa+wNooxq/pl2RLK8ugH2E6WDn7VcyPbJfEkS3JgMQivin2wO9W1
/b2UTbRh440lqfXAkdad4zmgPVlSdNUYJT4u2gNKt7Yu8Ygj1H+NxfXgLjOGLheR
hqsHZ/inyaJxrrk0KA33M848aom6menit2pWQy7gqsdXel8Lq2C+wjQ2uLpqsUjD
kpF4HUwRS1BM5/kebjefB/qpEFXBOBw69IePjvqpmgap4JbpRA9vNPcIHNQBcBOL
setwFnWCo+HtWZGrLBMu7NwEnoeCmRNjjbrBuknfFC/fPRWLghn3jkh3VJN7TMkC
5d0wV/IR5GMA5hU3k8LMfUuWnxYTTDGcFgLvtfUZYj3ia+eEvoSSrIgcMHcNwu8o
iBvJT0Iw14OIXN54qAmxa43/Gc/W7XznNbofwmLuRQhO4Q5bW+B8eX1prico43Ee
gk7daOK2Mn0hP0qCOK+5QQnNGRrnuMIqy0CardeWwyRRvk4gMkehzQuylm6ir+1D
mlCuGC0TO9+38L0Ezks4MvJ2Eaa74sSmZU2aQJxty9YTH8EAviZJyA+Ti20bRdCl
5ATgrKNEW2MwO9PLAkf7zgtonc40NwnW7QpaoJMO7eathnuFLqxpGx2wA2bUMz0c
OgDo0oaC6ATRZFtGVS/uCyW8yLond1g1LA6kkebJpuFKNNW8c3ozaAelWBhhnYxU
dc9gHmcKpj9TnXsvIAzekqKWlupYrDr0b/aF2gnJVsqkgqEb5gVpQt1WMyNmkI2N
qd6i4IQ41RFv9ARCOOGQMqF8gNDVb2dVUWnwjCETEPMyfbKwJEifN78V2CSvbmPh
JZoEusIC3cCNw6XYstv8sO9vRRP9KftiQTLDHRYbNo6RUDSXBRZNDPlTpKw5HAdh
F4Wb8+rGXHa0q/ZXievlddHLh4ww9oJXchGGxJ3KKoWX2VBtIHqVk3FLmYmbgn2w
ZpkvLuIwFKHr1tInEXwtuCier5ZPBV5YIsxfd8XI8KH1IEM0nqKBIa+M99tKOyib
PZAGnY8/iGrFaerqS2bhP1BUZk8VXo4GCp5OiAEyUIdQ8HJRNzZ3T7EGrf2Aio4i
WoiLR/SkxS5XmGeFfVYcJdVIq5R7Tne285Y37DNTwreSToYCEosOPngTwn016pWx
bNULA9StWHZsI5Dtk7Y4JS7MrZu2M+Fda1d0yv6zFm0q8e8Y1MezvUWpq32tDZNT
6PG0ovNZVgufEz8OYHLuRjU1tdYfYjC1ZK7kO+mqSg+dUTZLyYH0QtqUEZwr7zoe
Cw37jwSV6W2mZGKmLrawz9HXWQXTXIe/XB4qXtguu9+LcvULy9IrN2DSK5HDzmtW
3Ym/gvIrs7t14+EXWRBAynLQ3DnXtNdh8fq4hGyRTTm8m0Ms8d+HzieMVXsNqP8B
GTaOUGDcFdYzn1zYMIg7n+QFgz/zcV5JLsU9C+qbCqb7b4mBPWKE4zmO9hBjQEN6
+pA8OlPRLJ+k049S58B/4+Xl/BLgs4iv5xzLYTX1ApK/zabA72jDmK+lffN4nytJ
4yIjwZJaTxu/x2B5HgjO6WwCQL+9nTM2j9McCRralp8C0lblltx8gAMSNLQePi6y
pyKLfLMhySRyBNET8NsWGhiS7l5fwmirjGqBIlDA7AS9GuzJqYQOOXqoGH/yLLAY
u36JL9cQnii3GF7IuKqn3DbWWCfukloSq+QysRjK32jjLzp6aZWR3TagiKiPl5PG
/f28kbn7i0BhL3YB57CsmOIO/27QGAWuj1TQtbHoTUIn0U99MjazWUHXBqFWHQ3y
PJ0YHJ0pExJDfry0HLbMn5XQjRnN6LqBVZhxOAq5iCSsxRCVkRhtrhMRB6rmoanm
65AqqUcgTdF4fa73L8KVk5rf4PvyAkWQGeFudvXK5hZFRJcp2IAKqA4e0ScH9lX3
Ld2DH1EJSKFYyO+yWmEgYzkuSaFGrihRBJyuQaGBsRUwzjrZdGMzVOykZapzk7Jc
2vt5zR2nEqH4TNEQUCv/0ZktDsBdkk4sEmruuuYnwvtkzskeYGmJ6abDM5NHtJ+7
OeRKctBELTJ7g0N4c/Pq+eSTUG+qgTrKPRLqknKPnf86w522M22jdjgcrXyU3ECh
vBDdcVQhpcXeIQPwXP+S0P8FLo3QJ1Apo/zcqSN9IphcoqhemFSWnYq6gic5q1BZ
AZzuGoQ5WtbICP1JSVZhJOIWiV0x97yQ6QtqKGupB4FITXJp9+h0nYdijz4Y0F4Q
a8zC7c9UpN+fZPciHnSn2Uf19pseha2AonQfoW7fKGDylSzAxe+nCzeyvPssEaWb
8ZSPnUY3PnRnH6TxCp4TMSJvizKxD0zShm66BSyTtC7mhE+3qcJamIPfsYYm+FnI
IV0jTqfi5j6GrSTz+WnutPOXJdyQY2saG52ICGUc98AsbTAhDbQE0+NvYiYXf7IF
8tey+zSZXmvdvJbY6/s9i6y9K7+01r4YU1sENOWmFBvjbwFx5MT0bu32CTF+x2th
se9hZMCAgRjTq8Al5EzIvtPZto3ANl9qtt4aG24+aAERmY7/f/sqKA3L5JWAPEKY
yyiqXMyLuOrdfKC2EAyLoCJz/6DiueTQ2gz9VPyQAzqkRcwZC4jdMhh5GznrwyLq
rqmlDkT/+P8xXjLH/5Wdrafqg7n4tSJFAyV0E/Eo0E8iTxszD/mqO89qGWNzLtVt
TIlIid5XD0oELThj0iU01FPmKzC2UAByNxKBiaFRz8Dy8R8AbBD7ErZNPxXYnMUR
6ScsJR4oO0cvNPjP/NtQMxjTp2zOknwWpv37iBUD4NKCVkV6eq2iJHJHAxGGnv0h
TPdOul/A+NLf5vensiikEf3tvcOjjeS4xLoHvf04h6HbcHl3s2sY4OvHwrHEvZu5
n+pDwmQiQrIWSyjRk1azwsG+yua/wv2fNxQ25RfWpb+pPqkephCDkZYW6+ECPtSC
uwFsZnUKrDC4Tj55SHXYz+h+5/QE9bt0Lc8ZjkuSze56ELPqrSNcbXn976I3mcJ6
km2gRnRVGSlbhpSNpDMx3ZtrWbCvZXAGF6qJsQAwVEG/qJKmw8RTqB1Y1RHhjgbP
E6s5REehL+D8kbt7aAubhHgZMxACCdBkB+FKAsDJ9n3AWBDJq1F4zDUcO2SeCTkU
wScpRuU6O9BphWsBo2wScSnpVEiZ8KmUaJbx5UuQW3xhrp+a2KCzIDRC8iDmyX6B
IHA6alr70rwT6hKockKVBi0hYf3hhATODp/fSeYzKHwwpqTM5ZNFgV3471S/7fcW
0LRudh9cQY+eiXW0aqwS+K//k0PHGEzKvnrHOoiWy1q71B/fW4Cj8ef0qX7pjZ2p
1M7OX7iPGKBdslVRXTgQFFXBXC7oZG/V7n76N+5pZB4jmESRmY8ARRg9Fk9D3Dna
XEVVueCcdo1hUdRkeLasbteu93SuhhInC9co0CLyT9fI2bAuK5SQwmFQ6+lJbTp0
MvH3WXyl6B+AzHEJDhEFZgd2OQN6SydDa/pFnU74iX2aJLpbxIWKDNJCC8C8+NKR
P80pjquZgggl5qb90faaT0z56nP/GbkNSO/VnWT7cPfsfLV09VcwiKUEzXtAf5El
/T4hT0oXoFnWYCVX2W1ZPNXQzEIos5RLjDC4Z0eZbLRETG0GZjY/2n+/2sengNsc
NHKnV2UvjrctAwYPEnfh+aNXglycTs61qoMlEaZicaf/RU78g7nDnujKDVGAtZqD
01fCQlhlRrZww8CM1/O5P+4UzgJA905Cr3tcJJxRMGlEQ+GSrA2h8llcFlqB4e1q
/eH8ktqt7XygZCgzJl3PTadBmFTfalNryJ3MUD90JJ93MHNlMaWRIIm0vYU9nMTI
U+I5HfoPKLwb5T3heVd6Abkmr8/PVQx/7Rihbgmo8O1SsxiE4jWrhHHXzHDqiLfT
g3b0msF8VUkhAObgLDf482iPllaB+RUI3QgYO0buGGvBlGDMAdzRU0fs6H0l7vPh
4Kbqgc/rJ2bQAAuwrUHq03GpWqAbOsUxv6axa/+Ru+wtw921hGe8ZFZ0Xyk/UHSD
zfcU9kHYj/k4KLqfRNizkTXHzfSqKF4UPV/+XlGTsyYkLxL6wMHAByj0g4TSyy0D
NDZainwrbUlA+eJkGuJ82txhPayTQWZNow2jbbeJShzykTnvI04mzWHbWKNaf4lS
KZv7+lIk9ytKGVVf7y32pIjJYnirYZ5U8KIMukBZ3IkCZKaengxV+/uFUscVIMKv
1EcdPfW4FNNAfNbHRA8CRVlxlhll5iJ04AVZZkb5qfWU9O4SM7N1j+/sDv+6oklD
NdQGqhG5xwPb8J1ILNa1bbXOvAFAC56MjKlclSPSBAl0bhA3tSxo1dhYkmEshvyt
dRrL4/dDZ+742fqjcIxbspMQ+hdSBaeAX642kz5NbyEJwgLlumXldJ80AMsDgw9c
rYZDhCAMu3k08CB1RU7qE8zZmiLR+OccZFN8xTKyMXLfolaT2Gy6c0m5kbT1gZaJ
WTrNAlUtxgGwYEnBMronq3BvAV9LGoF2EsShHFzkISBxSpKn+iyUF1BCqMn+ULuh
Jv57npIlFaMYfqx1N2V/yyvolKVcb29moZEBT+/0aLZ42XlKh3CgahrdMOPQMHLk
gkrqQIDsu7jIH4rVabRvJqGsixtl0wPtGOUm81GyKHdT8td+u4w+VTE3AQWwccjH
f0ztCAQhetvrNRCvmwE9At7gJNH8AEEeMY0oChVH4cKlfngcjirWo9o8VAd+2DCZ
e44sGZKU6BAKguSQunEgXgwfWgSXFgkYcMujV2Xdl6yIT8DF31Xd+0q6OlowJoSz
WsVnmISJabtdxQH4y3C+RLYXtnLDEVw+STND+5PkkY/uSwuRUcbXjBZuifTNU4kD
8kVeNQLsM3l3SvZbWIwrDTvRyNqvWCq7k4xpsZw892QN93LhiuTZ0ZQZs+aPA26n
wf+R4EDclzVU8U/5intDqnUXSQYDKF7uOoUV7L4xweOSvzi5w3zb41TIILaAcdyr
XJaDiE03TclzsfjHz0eXGnEUraed3N0ftYOzc9NKIqZGqLuqhdeAtza9M+Rsn7pv
Yq6aAy7+reUWxew7/qHO5NTVA3L05K6qneAERhQtBcnjaA4bEvje0KM6oSPmbLS8
OlPYyLl3UteEWC5A+BfEejqFNURqgvvJunot23y8AjeEtTDPC8kde97AYKd1R9Ir
7hv384NZO1wyyYPJ8JWgjKoOA42XAHqNkI29GvSarmtHMTO5P/JtqheXtSd1kRnB
xZQI0+dQJFXWm0I0Yz7BhUrncLS+HyebM7g1MD7YOeGM7XH8DZMNxcOaLeL92lNP
mf3Vaj/WJARLJgbO0n3BF1ouCSwPhOmiR+tirsyK87dBR+lB/3pQgUggRPVsQam/
MKtTAAcxRvSZhauK49gLgdRtqallBwiUHoS9WV/p2aHSmMPRVCojtXiLg0dzMvOv
1JHJifzjqrFjVM5+q6R9Y81kFTU63sgQglG3XpJmqy5rFZm1RJQi2jJO6TAscHrl
I25w0818mPreUKOosLfsu+JVAMZtptA5MHZ1q46k82FON9HJYpfABh5SMf3qjAOV
i5Nu+piIz42MUtJW2JaxsEOuj4mJm1iigP+5799FX2TDRKZZBHju4Zcn9PixOHRC
ZOJ4kEf6BbKuzjocwCEuiWVF3BX+aUs4TF5RA7iWor0IoVQ5orQLcBJSnTqFd+/D
7Er7zPUVwbsScvQqDReTBoQYQWQJlmV5LD8PlMpy3OSTlWkBk5pDv0PE7vkF//dv
5L5iB89GwOsVAYl6Ol7p439pKNw34Q6PgScM0RWvr8XA+14P/Wb5ioZAF9+eNaNK
WU+UtpuxPg5jgFzGeGi+1Kdgsa6XVvwQ2gSJHagGdPKf3EZhJ+7zAjPU8tnOrm2p
o+NalYfsu3pafCEFDwxJi59HMSJc6Soa04zQHRfq7SAGYSaZVUacdJ4Wzk9fb/Bi
LBkuNPxmzBKpGH+5ZCSs/7w+zWwThbUHyowv/XSsw6DtF5nBp4JnGiV3tn8DpTHj
SZ1V6Ap9L1TFad/PKn4QvvQg5Eoxk6Mt8Puk+Aa3nnjjVxEC9S4YjMvN6MOhBMK0
1lqfiSj+cIu0A3NOb7Ut8uo73Tm1bRGG1npt6SWor90CgbR22QR1D8FP75b8qFCb
XQZoECPCVE/iEEEfDxwgokC9ZjstY+HO/3XMmRvZCD52X4cdnZEfWrQg7tmBtewk
sqY8r097xObhI18Ug8Xq/OS+jelEqNBDU98YILlkr3x7IBNDjbNOxx8dGQfyrWqk
2BMB91ZVF5ySROJaAf4XF3LY2L43ggL1NfJ15WSgkw6u3p868KqRectI0ERim0X0
7bYlNOQy02ZL3NFwERWVhS6bugO+q0HAfVZzd1aB6kUbf8Mjtp57okcHQ27BO2f2
bN8cxE+5l4K/AOAIn1NmPW2DBymIqlEWROs6RRESThWPNwSHWl3I26MkFRIqY3TJ
YR23E9YPZ4eKtUsVx5WjwNeJYKsdPHaBXeK9EvaLyvu+ZlpXoVlHU+uz5rJibLb4
PqAzH4yNYNHDNrtnScP3c+OEhioGpMkgcJ4Z0CZzOR/qqqpKgBc0Sl283DfudDW1
ODhQkSTlUkAOCcehuRKKDUAJyo0g+7iXwtxur8x7VGQN1GcCwzgfi63PIEDtGiky
OCThRG1Ta1L18Q2QuxLYNaootwrz5U81fjfe+1T2ooMQzFp2dH6GSiA4h1SkWEbc
QkFRVZ/kgBow2ro+vwyS5reV9/hE7I37nCBL2kqnxxpkqgHwHL9Ivxr5MYusHscI
OFXazblUgAPHPUmHQe4HAfLLlJKBIa+EmfGGmC2u1LcsRKn1f41vHRuqfr8iyFTQ
U55jDIJUwuIvUqCAuyXmcR7ar1qGW1mWdZgcKcShodg5NwQZEvL/kPVEWrhi8AyG
ruAdTdI+ysBa0PK4GaaBv6AJi/sLHYN3WPfnotUEWLO21AN9khRcbDpGAo0QzlSi
/BYGyYfk6RPmPdKMqYa/tD6LmYLZmweknBwuXHDIeizIcIi6to2A+pNKdULzIFxR
P21dfbPjisQO/FR/ltXeunG3TLgsh2RDh/T25ssmrc+Ufk/5pmLzrcf5N/GxzRha
PWYH/FYx4qd+ZTO+hGBxYChAlGVgGkpYHGvdHjmq30vc0ipaCN88B9vX3iYDqLGF
Ujh9FK5IYizbBd4/sCu7YmYAcVvfMvHHRRa75QqQ3legIoSydOPOvnnNX8kFs72p
MuHPBuvw4CWhPH0y7y3OG/hk5lPjitPvnEVgRt5nVYymsiu2qLicUQFuuxHjwEf0
JGy+I9d0vRYWMo68II+xPfqfvdtyaUYj5HJxvl8auCCq92RBEkiAlRVBXvs+uRLJ
yu64RMD9moR/1c6HzazszVZ0rkkMYSfWSf0w6skAJBlH6KXQ6FYmPFJkm2INHzG3
mpiG3mtOPpbIstbzkU4pEhSkHU4CK3U8KFpdcmSAA6/UR6GUytifIa1LmkvRsgpS
H+aXV/BEIt5rWXU4RxjBVuRXAzCac0iBr8JVLHTO3RBUSZwB4In/JSbiUM+URab7
fnXMLxPJv16xU9d9h4Ovzsdcc1MqJXCtky0Uk7+hr6Jl2UmVTtStYgXq/FZJTW0t
qoB2/qqhH74M1MOkPSX2mbRR2sQwT5jJw2BoLxrvT2V/R/sir/ER3GLFE9x52uS7
T5/eiSEhNIGh6O8+DcsuuIB2ZYgK4i7VYbF7E62T4T2AcZ6r3cx5Lg3OCnseLsfT
ltL+7v0GSrsmX92HOlWgbfsvnh1IX+IMs4k1T/M85G3xICDSD5p2ZhVZjff3t77y
7VCFByWOBMm6ZZqw841e7/uT0ZluYrnCxAukiwkI1BayQrnFWh/JHVBmS7D46J8k
I4kodnhFzkoqVPMYgqhV86EVVUKGz1avuyPh+AVplZgW/KdNpsz2dUGOPXd6h/+Q
K+7cacQRYQGdB9w6KfQnPWHbh7bzL5TeF7HzqDyMSTKbcEumIrAzg5eHdhZKGXlY
hSpUKzL1VUcZkGPeaesAIPERhOOXBiHojyRPxWUry0dDdfJBZ/p7QL+1In4ixZ9p
llP3A3cjg71oUIOYge5RcdfnLiXy5V1jB/OiPcKDWkEnEsrkuqZnpkXHfoQBQBGD
4FKCe4BhmbpukFgpvJu3NUXa0kzFXwrpngl0YcmrBaLfAgHdL1yO4b1863UI57Ok
OuZ//g/R/4tHBJ7VFhcF4I1KrHUZgFj+6P34Cw3nGbOtheirnaaF1waZ/SRXdClh
Fio0Zgc2oY0vSTBZJwJ2ic73wSz8PRkpMlJNhfxG8GHCY/Ipu+tkc3846o8VstNC
ON2u5yC74GEoqw2tJDKhWdfm3RLQ3pBacPvFKQ2f0Jdy7sZpDdFQoGziFsQl1cJz
XGUSXPvx8wFCUFVUA8zgj+7Ni9VYa4OfP4ikU1/1g27Wni4LSLvEE68FuPbSy6w6
FKtZ1rAWpJ3lgig1RMYS+bFdWLs075iTDtD4t4rVJBTyAvGtQyT3D8R2tufT3hxT
fPe63OxIk+PxqmxdjZkVMtp3ofCg+97Toy2emd2V8JREhkiVSbI7AuMoZAWEj3n9
iZLWQdGcSEmyXEuIoOFJHLYVkU5ivcX0nFCmDwVuh3jeeDQIxXL/RdXBHE2E4UmR
6+GRqU1NR2xLx0sBeTSZSDK2sEaTgZy34aDmCASDBhBSKBexyd1w05dn+BPk76+i
o/SARCDtC3J9TMwD2PftxsTbluYKqil2182yzmVJ1W1ElJRQYRHZUHqf4oXgQ1tm
aU7xDdSHLGbhIoRxPEfgOh1axfU/v/KbXZw3t3hwEW55nPFJZzUpQUz2ELxmqFmy
c90XH94OE6EA8CJDNOdlSPbha7TD07E8hR7ZDh1PmnKAkuqD/4izjBm8o20zrUAb
ROJCCoEipbk7Fask82F+/HBBzMBIAB11ltpQxXRCssDnbvZcEPzl6BeubbZhZQsT
N2FFGFGmhH3sO4Kjpu5iCbhh5G8zmLxUDFql5Q6WhyPgQ81egikNpYxyyNRg/CPb
4yEXI6/tJhvQovQmRxkv19C89yZYXt9LUU53WAAo4VY1XkX1AiC/8rJONEvBf4M+
CJDdaJzmILxUjIeCqXyDrhU3jVRmMS9t+fWKxlbY3yg9SRaIfiegz6fHn7pGMLPW
O1ZdONLhu8pa0AdhLB640qQC6LtOdjg/YxpTnysZgm5ZD6APl50AlWKC20JQS2d5
W8GV/AzOqBPAqAtixk41hfqJkM4TpcaRtdSNLwo7p6QIcmyE4375ol7lKpcHF8QN
rVN/UDc0o4nePp5RWTG742W2pSjbpOQQsHebP5WRSWQU2u192amDItLYW9y1s3g4
DNFzLGFDHdNbv9cIUB58wP3kMz894MCyeadZiArzJzN+yQx+CRK1N3BVYWxx3oyL
c4esB0TViB+gQc+9zgCTQL4M2DbU8hiNNT0ZKUqdsHnPdQPyIlV6Bd3wyhtbS9Vo
3DZ5zozLdE4jlTpAne4o/tgS11ols9ACpjKD4h6sTFnUu1fNzUkLY54K7bhVt2G9
bqVFK85yRdVFWqju240C2X8d2eBki/unhBk28xVRNfTILBp16hwaAWCDcTq89O/1
ha0WRm/jMJkfyt9+8kmhlELhPEp8lpDAgcYPLULXb2MkiG6aMgOpb3gQUGMIozkz
F8tKvpzR0PKv4iJQhR1FuC8Z0bDS/6rlKJter6P3dbJDGdfTuwyS/rLvx1zZ8+UH
CBhHGJVj7QFfFRv0J2ZSkaevFfjXICKJISDIntP5gsggx/JZOdc8C6Xb9H+9IJti
w7gonDRF7F/BpYlzWOR4mg9wLZvqZOFXuWRKHukgxYmdNw/I66q/V+MiicdUiu9d
LQRd+em187BYim7dMXUz096UqKJBeCOuAEtUX2ihk3QSxD+v9v+PaKU/IOOg3i3x
SNCkGO4WiM7+vAJihBugPLKjrsbJxzWXXDAaBgSMbT71dhe25xFFAVSao+AYQSGD
GU34k2thW7jg3LHTE3eq9yUBk+wCEECpvok6Z/fM7aIz0n+EocRJJhjSU8dvUq1i
Wd4G0AVvEiWexBxfc0it5bGuvqDfi41fvcqxGBijAmX6Llj2wJkWoR+rbLn5VcmH
vvD6Vpa+CPHIESoX5mSrS2oFtzNNVHiBO/VQj0FJqN9HOFDS0DusrUBHvCOsfzrM
+fgsAJFm4BRRypehx+ovHIsa4hskIYpfL5xbM9Gwnz49kZHx0RNOKngtIaEBzHOr
ebPAErUWZ6SMt9heCO6SnzlPLAEBMxPdWaYuhXqXTA1zUEWIl43qpbtP2SnDfTlO
nr/GABhULpPNZgJqPoDXyRIkonVM9+MEl41syLeK2vAaneQ9XLf9Ba1wmkvSO9ky
69pQpQGsxon8kx526TOVL1WpRQA2yp+hT930gnyaA7p42ISYwjEfzUVKU3nJMfjN
qTFvGVXQYY8OQ3uzcO5o3t3DU438f1qC8OCLoNkgOG855r/5CvGliBqR+BtiAN5I
3tpKSd733NZ0wPaAtWsL4Bgz0vfNzfW+q7SPQ/SwLVOaQDWu2cAYSJSklgsyVydK
gJ9+YYw70MCWU+CK9SZ/ulxwkfaL6FMznQGfv6Q/el4kczBLY23Np5Rhi5eWmDIq
+bffmC1cdgAHAwUFvDN7F1XXqW+6zGdz9FisjOpgH9S8FtIqxahlA8wGJ8z2GnQK
XovftrdmKC3CPIKyqN9w259hSr7ydS0CdxdBDOeXYZnXZXCRpKWDc9uz48KAn3/p
IeHzzsBm64Hj6ob4Poo52r6I67a/qCfeB8VeIAZVcCfXDKj/cp1GcRdSg+hcGJMP
JAU7PHTX0L5mhXZiN1FWPFG9VRCQLe8r5ezkT6Diqk6m143Ubl/soBWPUrXHwA1W
E2X/IMFzjc6fW4UiH9N/ImXfzFf/02o8qnNAVJKB6JdKB9XRg7MnHzIn2upnM89I
NJ8dPYwb8bjXGqd6oBiMCHXIpmkqevv0HlmmD7PWkdz5ykoq5EUpu5xm8NtVeNZP
/MLImFy0gR327jv5Wwhgk7tc17Ri5WZq64/5qTZql2VYRiHg5jv0UAwQrdKr2vKC
Sd2CQvrXzreS2gChrqr54yGBLwEf07/wndy3vDo7u/Uy+oR9T6Jkyo1A7HopqB+p
GNstVFw+fuBNYVjmxct/EHFB64eCHephSRYVj/dqWft3ZNhFidrm7xMx685otI/y
XnOdWAYg18Fy7J0WYp86To22GqpxFZud8UpuQsG9S899cmuES+xVGIJS/XCG2pvT
7bj9/hByUp+2XffA8tA0fe2pegDqnmTu4Nprt6Dr6v3yvp9xfm3/dVIWb0UbKiAt
Fsexy5sRosJthKIr9vtlqrJpMac9GDQ1tnUC6ObtkftEgS9bhbcSZNMi8aAhbf1m
XJbqXBwWnbcL/0eJ5nD9lNBrzuKGK5dezRPxZqx4pXMrWAGW18x/p/AneovORNCx
9hynM2rOT/j3FXxo6LBE+Moz5jtSi3vIlbudRXh4IXTGoHRfVvFdwmpbrQ/MeJMu
xUxj7QPRglALZPUGKU0vcLLsR30FeH0ZH2yZNic4WCGz+UvZ7jlavk+DfzBKUYfT
acXSfvmMtmg+qpiogS68hGusITrhzgBIHtGrH0CT6R5PGT53Tmsuda0U7QKnHbI8
WkOEat/NghesqfzHU1L+SijIRltGH4KOTd7VpPfFfk7L1B6cXqzmkRBSKodvZCAQ
e+wJ0Lc6ixWomlTF5vrYuAnGqD9FoK2PmhK1qO6VqCtRZa1Zs9ProsI78IP7hDg7
Da55YftOv7ZspeN2t7rpnZGEaxwe7QFrbTGa37sUU8ONVzN0s7Xq2h6huThYwOit
AcVyedKJDmjRzVfkLyLFZ8d0opX95FKrWk8fYwdDkv+OoYrbU9gFJQ63hysDzgtz
KhCIbl6EaVIs0iIVbWrDbxw+H8XiQ1Rw101SpwASKWBGzCdWbs4uf4e47KemG8jd
tuSLYgXvzZyDtwOYLFdA+IAXHSWY//70HVoNsa6LZxoKRMEn75W6B0dQavBAqpYZ
s6aSpXy2H+0N3KojfoPOOaYFsTNUDOF+qj3cpzojlcXniWVVkn7+CmuZlMbIr61E
OGZd5vkotufgWnr4Y5HRwpSXir22jNMnQV79m2NJrAX58uqQoipSOSIlAEPUp4Pk
OajHo5Sj1jZorLq/Z+/JIdvtYChBW2NIZSVUWBmeQlFqwqk3T2B8nyB6DfLOdoym
TG2hk5tZK8S+PPuK0hxnUvl407Na43g3OTTh7ETzFpExxpyZFEHmkjNt8CYmDMB1
O6H/i8uxlaZSovwknTdsZyKkNahqetdGjU5vHxiDORWOynWRXiRyV9yNT6nej8PL
/Ia0TTKQ1yZZ/P7xQer+s4jUIJmIC4jekuS2+OG+o6NgTlFfxBxYHrp4dfzWnpzR
/bV529ppBIxRnDfg1Z+X2vB6Cna0yUB0VLfyEPqDBTqLg/bgk/m/P36CIuOBrX0Z
y8Qw3ISfpeFTkY2vlro2kQLK2+xSXwfj+cIn9XotQfS1DSTrJvOgZ6mGRdK7HG97
kJZtmmzWpKt5FO4UHP//AI5Jk4uJxFbtDjrAzaTxIen05CsJGtkJwls5KGjJARb6
aszfJNmKKJS2RcQIecFl+pAZiWLufHCopuBPdKdU3P4mtB0g9Q/abxq8KBGIaB/i
7lKRuse8+J8T0vsurdkXyPYk3bJ6G9usRAz3+Db34aeB/D10Sl1Vd792u94okz42
AoDfCYG23R9Gn3eRLhiaXF6SeaLE1CZZETeB7zgcDc8tr62SdUW4ZhwSv+jDm87Q
u2WEdbKCSA4DqNVwvk+VYy+VSJwl2HOctP24gscKf2MxsoNQltPCbP/nPgUXcLcp
6wx6Ulzin9a7mLynvqIwynq6dOnSJIy3w/9GHkZHhE2J58om1zrBLAr44uUjI0Gu
vCpDCfaHsrlfXeRdgiJOM2IR+CwN8cLIvH8zNvoLxd4KRMvxfxgp9/Q4oNMrps09
N0UdH1uLh1Viwnak1TKYvVbXqDts0pe9naxNwd3AXdZ2LGjZuIMDXdrYfkZYMvGd
CAjWVyRGfKKTreFbFk/Y3Bua6j4g5GIuXKv15B228WWD2nF60jqwhzg8oO9IWi1k
WCCkWaWMR+K2FgQjgOq7a6oVhtwNfxFGxUEX5KLyT5GI4WzQsaY96t8pZcSaGAOk
8yGzJ7Kc3IGCrOS7BpRJl9RqLqZfaeVwr/9Gd7ISJOUkA3HNhwIJwEUw8xZ5X2SE
a60V3SbwAq/6FJGa5xx2XWUBL3Qq8LCH8TWOP1xeFidulmd8RvFGUGJ48dKjjKvd
0gM+7/7YlNkIvpIe3yPvv/nUG7zKbRLIhd5WL5IRqZlGaV0VO+/hmlxLATDq5WO6
Xrkyg0PJyioLk8fbqWyOvvx0Uv2keSRjuOAZaToOJCdGjcky25rjFoq6CN9+YBUV
0aAnFJye29ZEjxOJD1erGzK/J1HSk+fr8qrQML4pr+g/r2waWBHPzD+iSCW0ep00
kSOGKy7o0j2lPqTnKifJBNkpcpeIaZJwmk01YVqD6Hanmm8TNcQ58WEA2e7bjWmP
IdVSXTjttCXZoflsHWkENLyu5JRc65v4BGz67VNAsVDXaX+uQMya0qvD+ZjOD0QG
AIhh/1B9jZzKPYetbSVE170UW8bl8w/rC+mm4GnjGCdcbLqjbpCveoLchSsvtg8B
HrLSdTWXXIH9Hf00WSdtf+3GtNgPOXvv0Zn/tVjDWXYMXi2w2Iwr5Z/3gnHMtYRi
ZLv5tk3xGxzmhbvaAgjjEzSI/4OWo/g2B3TJxYk+36rC0P4MSTGn9RYzOqNay1z4
Jq1iFnvORVbHtefi6WwX4jIdExAQilknnJ7+j0CyA4N4sqATOCd1UvE05aW+VqR3
kn7/7mYVI4jfbvskI1nuKNXvpfWU3FXBly2/S2TXsUbXtkfDQv7pnZ0abVtV/qYm
nA6bgKreI91mqMwLpfGfTrPXojTGqwZ3dU4Qg879SoWF/ehLGzlrDj7w3DYWrBk4
s43HpCAP0hqoaW35ZWF3sSf2D+f+hbkOr8HCzAFztXnO2tv1anaeUcKEGGACact5
vkk+9lbgI1KQ5rZ2xQBku9UDlFkEP+jwToCnpqmTDAYmrOuvtvfGORr2HF+UlWGz
OKmkXWjTGzJh/372lmY8SUIOzbKJIVOL9uXRdKmm2IlVw3YW1qjnQFT6Tta9nP3A
pHB200rmaR2aGYwQPytL3n5RHpgEmg+jtBH5s2IbHwVL3eg9IwDUreM+QK2eWara
5K+i8z1rOVVtT47VoF3V3qyjdZNYAslsUHBbGa888WTo6j/Mmj6RltD0ni/BV7FG
lsHlLZ1yLcj6iOl8Ei9RnEq+HQOuMgkez6AfHHadG0di1kVOWvVau9S0UqDIV/Kg
42yvx/6NRiijbYymaeHg9totFpUKgE2lS4x0xNo1CUA7qZCPCVWgdLYidzUQ8Ler
mJ/KfE6r6nTx0Ej5Z6S0W4ZYzwXZSPbJkY3EgohmjmZLV7HK/8xOeFiyoFBc7IoG
MpKIlZZNYP34xCw7T0MxB7uunTSQv1jJJPH8bDM+P80GOWFwU/P3dN4yRX/aeove
BKNiYu3OvWkS9LOwOokciBR//OyULpXH+orlUBFJ8WfKJ82u9OVaEFdAZkFxvaVF
LDAAAyqyMJv3h0/P/Du/bbj0eR9MetWcIil7HDwRXChDIJg3kCp6loJnJ4ycolKW
Eq525v9JIXTQTEaUOrfq/O4bFLXPnsQiU4VGS1HCk/edj6hf/NgxDTubG1eRAoiD
NmJHf19hR8STHhsPJBg/RVOHk5Bzz13iGX48xklTiT1r6TCS3Hdr5GkVXxy9r52T
PnS6WcufC7K2XCNoOjWldyeCWNYoEQWlveVIy9oX48bgxxllrgo9VNmKPPm7wlqq
RuqWyYBTUT15bGFra/Vo2No9vuHXSMMMtthdcw43mAILxP7uCZ9KSXbEYNTukKBR
QC95myVuVfhJYGnry9Hq2utWzI6/O326V/iVCkA+1+/OcNXf0Sa+xFe88eqcZd3Q
SqNvoz82LfcFl/TsfCmTD71SJWVnzMb0JZsFsvSpmuwB6as4Ac0Mmdn5axqs7KWp
eOmpR0OjCWylDraePA2ACrtbefMVQVzhd8+V3gevNnAGgRVmmV5Zw6IY6+2ps7zu
ttshW/28zD5i9kwfkcAubo8mFXJPWfgvi4G4g53bxN5owTzcPdPGyDX1vwWrDpqI
ikOMS25ig+GYPOQLqJDmis65BseSCn5aeUFT1iA2WhhpDzxIEikAcX6msJ6TeDj+
S53E8Kch5damIsdAJgLCZOQ5KrxiCKnTaxtFqdvnjQbAkGWKXhBkZoxFjIrInmRI
WYxxqQftjfVg18JVJtE32qxEsPBVjaXZStatqzvUTr27X32ujuug44ZgXsW3xs7N
QTp8gAReqN4ycFj05zQXhapESNpzEhLtipRhbF7s8JBR8JicGmLFIpGbnPe081R5
qdOZZHQZpXbghIG79HHpFxPzSJNLLR4b+NUkb+5HjSxmKzjuyeXKbSdIzJ3HGQDV
xsGHor9teYPnHFnH/u7+R8KyxYu+Cmnk52XUyoC/QEDkteh7OsiaoBbOm4iCPS53
B2SKMelj3alofAfQGQTwwPdb/BVKuEDfns3mIuS9NNs7H3L0WZJOrT8qyZC+xn6+
jVQhwUkKxxHW7bd6ixI9JqdxGe/p1UOm6U4M+asUtV9eYLexXIIcwGqwUvxHBcfC
nS42Ur63eLWWiYE9lf7Rs45QLToDM4plRo94YvYdN9OykGAcZ4rRcOX0U0P+pP7l
Nogk+z+clNsad665Qw2PR19JKVy56t2dTEMXRgpglo7qNhSM0gDkyz4PV1Mn7ZAA
Hgluse9s+64J2Xl54mIgLE27SenNGUTzvIHwfq528TFNkI+1qBA/ZfuV+nAtqb9D
fX1qiyG/JUYi7oGr8N+KH6zjthTKRc74ccsu/WDhTStzEQ5WwiJjh7A6IoHCXI8U
IMYYted0j2Tj6y4oh4dimB5XgHxr9PU6wAWWT/Ja1hweRA9ix20Y+Vitm2b/UUZW
88GQiA/MU/+q8yJStFElJCTyAmmxdvZI6mke8C3db8a32ySTL08nVNUbLHaNxwQK
z1RZPfGg4ki8or2ld8HBWUtmuh48EKQytn4QmLTzfDura0ar4kwQxvbSAp1VfpQU
F5ywfK8Ur4ph1nYBo1KUBZe/1D9x3U+uPJQ7ffnV6qXhsmJYPkbUQUyU7QXlst3p
WDdYIpQwb+QsJCRAyralX2+hOidRi2k+5ion0fG7byEYbsRCN/YA1yTJbnU+wRDn
NQofEA1091XrL+yXu3o2oKhu4cOGV6v5vyii1+B2CFqYtqZ+bMFBVAx5eS/a0YD/
GBRe+Tjml1w7QebdRlP7UihAZrlVybmZr9JUZ7niQpxWTv1Yu/yanhMLwFQlV1WL
cR3gXY89uuXX66HAeOW07h+9uTGeH/ExlwI2ERrWXDrFcZ3EGJoxu4Za/jeSlYuu
USFjmkyfPFVCWpUGqPclfdpp2e1haI1TKT+I+Q3NOzB2QNk0VW3aZ+sXvbKTRD+U
CU2X4c6lbnT9VbELdboS6jMDo06Zv5woeLT+j3XjKu+Rr/ZQMZIvs/w2idG51HQ7
SH0mzt7u8XAwnevWEvRE4OsrXZ5jE9E0uiK/QxGkOzngQXF5bbgHxwmFAc4LVl4V
h4bGWIYIVn2JStTxQx0mov0KU5UxZkRlORp149T0i4oJfyvlEENUkfQHQ7wfJLtM
bynbnx3oVuXb3pJTIhVru6HlXqSLLwK8a8aC/e12QU4cuOBgSyGcuue+Iiy5h31m
XxNJ+WxG228zfCOca5VMajMCNSkAuJYTN12PxBuVrqlHY5lbOqs8bN2B2FRbaOFR
282v3WBk816VeDpSctZBhvC4inj7oFLD0JtM5tkckJUvfftrbyoPjHXjLrZnkW7j
hnNBYQtWWzX1ay9B0up1BAf9qyl0rHyw/PhL6OdNewKKUNYYetAWbhn8dMlJXqNt
brUOw7SUSp5j2CDMn9NU+nx4BlSpU+3Ws45RRlu0NTK4vvjjSGN9MCltIuQoquhg
Ap2F8d9c7EytYrZLHZ8Z+C59ZHzTnytstzkE1g4Aoqpe739HUa5hEyxDSpPJEJU4
RCQjLCidEt+DEvjFiDLWXlBaWhhX2lLlAY46ZTaY5z35OIZXGwCja5D2HE2WWstZ
L1Zc4I3fRE8jVoO5RzEC7XDUbrHWvi/oX2PLJhxJOtim/Z5clsRTki0o989FVGFF
w+BbUpygJlt3sRJ/VM00Me3sBKve85HvGDx5JS3R+obC2eNnxK7ncrJP9T7Oo3d9
E+TBwuo4tMZ86wdSem52v5rhvuiWu6E2mDKLvoxt7pqyGqFfxe8d2pA+ZYp3g5EY
lTuNn8aLi5CyFfpGxPu5+tMQApxqSB9Abxx8OvPu4gkx6y/rgIwIZlf7NfXXGwBc
fjHOkrU05O5jwcv7WHpUGXZoTFhLyqNtsYXdz5CVTbpyUp52EnuwTyywA2427/Vv
VT/zXbPv5Zri3kuoRXN3D12MNF81x1CfSkpi3Z4pnZlg74js73qcSGnuoydjAtI8
YI4z/B6JRb+iwt/rc5r36BBkXKcWrOkdCNkdjLZ2AUFEoMqlVSxkLFqdd7J0CiYg
DZHOZTntNafSXuaMptOAzyK0ac3wCaIQPQJjJJHy5mbpfKvSNlGZOfkeYO62ttb1
Mh4luS+kYqzuQoZ1DEeqIsAr5QxlUolcxKjrucrfgm7ssUu9rVntl6fUgvUOdyYp
aYYRfz1QgKNzC2BJnsbfda+uVsjt/gzaaPOMIJ7Cu2woLkzjdVIMfVm01EW9CjNd
2CsjR4Q3ij46O5pXQFogNR9a+1pZH0oSm6pXr4CNrmCq5obJlIZ3rwzqaiplovAE
qWVltXtD7JTftuLKGna/CfWtQhEXZVtO4EHm6H5Kmyx6jYa3TlSiLCFQd0ZNfbrh
Fga5FNVlHnG7klVqfBG1u3YJIkgiPos+Ar9xk6sXOSxPSgE6Xyj3kQiwWH0FdD1S
GOVe4/g5U8a6fcf5kzg5+p4qc1FmRplxc75dD+l30aMyhcjnWxr23afAPgL/kf0L
+92SyiIe+O9L/w6U3KhWAW0Ypk0Lib6QlBoRMBpdXP9WFrpbUpV8R6owvrJ0jsPM
0M62vTJOYlbWIl8TKsRyYt0d88sNysx3n7YCCiEMBX/VVH8LqwSkrffBhE61SNdO
2mEATK0WKzygWRNidcRfakwKVbBT5DG0BACPWEAZlvutxPALmuG9+n7yr+zS+Bi/
ojlsOZAXIGCxcyx+Mda/PTuaffgmymtYJUOMPl27QEu+3w2BF21x7jpsV/Q3qH5c
GzcHBSSxSHEHOwkGQw+HiL82e4j+RINEFJvrNpBX4JjPP6z5eOUmT2xFZH6WdGKq
UJbrtjQLXjciCs30clU5oW3pvQPEzvT/JNTXMDKtWGhxIH6buck0QVVmCoSgMud7
zNKznNCBj1K1Z+u4yJ/r3L0moEP4vCH1rmmC7XBdCk0UUR9ncYwfdnlYD3NMSE4X
qDORXVtAfwzNuzJT8OlDiL2nq91QSvhjRN79f5DqIlfONWgs5W8ZFYHXHbJxkn9z
BoNcUrZegzwgTUIE/ijINjqZ3hEOQCpz3YlvkMeruc4wr/V/7f/SpVlsJ/g8fwHq
iwoqHvceUK9bWANDggHi0eRL1OYm0rX0bB293Y1qinMjcgJoMPvkLDx1zIZZc91+
43xvYNGa1u9C8E2/CWVqQ9v07t21lsbLOfZCLcbrXIGyOHDk/9JQbCpDxUfUE3Cu
Krf6N6UrWIlR7i1qrtD3MWZKmBvoK9xl0K9QvUn21TjkyLKgWA6SNJX6bD/hhlPw
oJFi1CF5myllSzXAe3oP03N3/Rzv227Bd86FlvcieEx6I9tfSlNXDgBVT1IgIA3I
J3n46zishzsDImoLk8FrulrDVI4yYYpihd0YuDH1AbA4MdkkbOW2A5x9Q6SOZIDh
ZKc3FnzYYQw5zWMIBcE9OaNyIO60L2gK0cJ4Pi7cvSKQRY/Wyf9hJ/tjkRGBzbhd
QBmyqFGMQ+XRFol2LgShLroKreDw1FaTGpSvUAXY7L9nVCQfFaEU6SyDQ+gt+rnF
gSUUFfXKLJJE74BoKTlSX2NWaGqN6s52qPZD1P9q0r5FjqRimBX2SpQVJE2AGfXm
j81h7eJBCB9fCzAV4uvmLgFLONRIuubRNOYmFckD9GfHk9yFuyrNg9Bf4a2DOJfE
WCMa+paPrUdfAJokj+McmVAEeIat0soin46rlN9ay1UKY4gnAUTDdbrr1j0xbCaT
4EgUJCFWLcpoXMo5SudbdihifWjAlLL8nyH4JjP61CtImAXUeJp87e6CzCjADfdt
TyXMdt4lATztPcUxXaEnZKG/dKTkj7NjrkjEI1DhZQ4THgLzE6UUhzcmZGOHE7nh
qTfuPU999idyb1BPlPCWsG3sYleESyPexhYOmGgq05jcR16QA7ppARKTefJ9sTGV
a2HEAAGI9y74M3TA13L1+iX/SfXkzBjDCxtizBdED+gF9+G3wRgNGbiwiKblQ0YD
2Xtr7EXIzL1s/Hvd4V+SZkI+TcNnqBo2NEmjZLqbDUwREViqc29KoNTKwNkrAeFv
qNfHrx2kvelzdgtD8RLQlz+G0e+BGqQUQPMK4QiAqGGAvxzkr+5TnUfxkEHP5kOt
6sFj0VMh2CylKXETGhcFMu+anVRN+RowtoDFz6anpm8Vi8NR4+HlgSmIL06QsKek
LOGcz2S2/rcA1YXiuHNmS9xWNGEDoPtE1cmcPZqfjCGrlUu4PvSytuo040Y2zPOX
Bfa85bfgH3Jh1m4I4ptBZIL3bUY5rfDJLydahbkjVp8YCve+JHe3o9cwXU9pBXXO
ydi3C1xcNqo4h9v1tgalH/gnpYlZ4M+gw3WiLuurbFLFc0GkAj5ROte/8y9PEs+K
Ue5Rf1Z1apPxOBbrAyLX+2sd17vTteytt1IJDMYzFvWUzxqo4k5Zzf9+4hx0ZLv3
aFLO1FGBcywaV09rUquQjDR+iKf0UvErlaOZqxmxT2o5unfpuREHhTGCc1srwIHd
JA+V0ZCFU6uZXKrNpCNmPcQp82wpTcCvWxrjoMY5DSl1ZeSsUSe9d7CR4uZXH/bR
f3CyLgobEONzQvzv5vw/U60ptlRTZPNOyqrDzipDI4R1AKD6ZCFZl3twwDMeFR6Z
5damzhYZm52f4GDZRwNHqWMcaKx7TbGWzeFsqB1EWWk6Ln695fJOIhmVGTFBkA3m
ylh125WEiRo49JmjH/jrUmaDmKxIbzvLOQdmqXVkWbyiZbtBGy7bMDuyhdwchM4C
wT4wX/43fi/KfpW1CgCi3vjbtseqLYN4TJDlZHCbbuxtKIMLXGg7lXZLqTNbgDhB
LQR2WE9Z/Sx47MSuOuGV9J2qTSElk2r1X6dZVq9RhA1sP4yd1t5KSJNB69wpwyGK
Z5f6Oejk0waFbqvoLIm0oDHn5j6G1EneCTin27+S9zOCyA+pbsymoyfv/CVENiq4
fGkmum9ESDRPn/y5gF3YqJu348QMcA6Rxzxs6kFzbECoeFPIhZXfKvHLVDK+ISl0
GVp/9PAQOYlYCL/rvDB2IbAfX81AbXzFbFvKvhHNf91IuP/JFeSjkvcVS5G0To7u
1lFhBv0TpkGu2c2HOcL1eerjEfrg9mmsyeRACUCb+CUCxjA28V+XMY68qB/Amzt6
uyJIyfwQMsJCaHOioPrqSOZB8RxqnhhrB1SgE3pNDAA9k7gUHdmWcnhvg6frBqOR
non0c5/9Rp2TQwiA857UiLC/I0IThTYwPUuQ1XhfDMiYvU2r8hlTzZCebv8eZju4
67KXQKeaTNzXYzHbZNVLc/1ShaGjEFDZ3IyJs7RnGfeddXZdk5W7/Q5sx8ay7BIe
b6iESzgMQyDRvvnYIjIhJdLBFD4ykB53ojk5X++/Udf8q2WLiS/31yU6u6AKt1d5
PMOiHh8OMsk50F1YKMRRDfn67isD6ohq9UWi67cYN6Lkbfvpl/XIiSbC2R3LUIVH
DsQ26K72rdwNp9KR5V3jluDX3XfKzm+kFZl8xGbPg2faFgWtpNrXu559baWmsh4S
QzJ6aP3gIx2QkLDeNTdv24RwH9lFxC4WIkwj5Nr5WjRUqSRrQ388Pd/ryxUkLrVs
FNKVxibzAu7FoSMl/DGxApcyfI53EENcHzWsVPFo4Hot7ePtsBEGeB9EgtvBWgB6
8+Ixdcs3+v1CvGBMBO5/bUztXNH8aY835Xjutv3AyyN7STbYvcr009p5fL7G5HaS
I99JFpGjZ//UW9TQm4yt8EKxsr+cE+sMo0giBbIAbYU5gBp+z0JzJVxGquXNzbcL
j8vohE0Qzhrqd6XHRXuogLLs7cluITWZZTR4VRVwx1NgIh8A1VyzaVbeLBVPF9GW
2P/aQSaVjYW+3xbYw4QBdA2Aov3+Q5JowiVf3ktIHCWHxF85LrSJ2ws5tvwQ9EZd
LbU1PBGr3yeNEkZIZVkNR/aRWdS4Sx5dBtxCBQUPugHTBX/tfsZS6wRDFPj/u4sv
JmTRbn5WVfbmLTYxmM6mho1LqvjxnLIpYWVTW1InacMABlDLPM7SqZ5vYOSXF0TK
5SaWScpu3sJEWZ9Lbyy7UXclKLRtySejPYnYlfkFun9nulDn3AhtRKXJw4utbAXC
lnGqBaBnUaqwr1r4aIfmyLatm4IWCBAyn7tZ1YftqlAde8D19y/M2MAEYpr4azi6
OBds8BnesJNLW5IE7jcg9A5nEAeXOmKcRaO9vp5urd3TwSRg0g49V0eCyv1y4J0O
rFP/XSd/A9LEDpozac+IYiK1b0ork33zUadcxJMVgtBj4w3vUZZ0GLVOQ9X1pt8E
HhNU9CQmgAWKJZoGJ3X208FuFz5ftQwufTuhXzEhr/5iyjJiRtCL4gs1iGOrY8mo
5N2tp/3UtCPxtzdxZSXYwAnVMO9A/UAjj8Z/oI76qlDnf7YRONVLmKrQN8OrZ9kU
RoIMSP44P29JUs6o1E46wnUTRSCIM0zuv+XCyayd+zdN/iJsqoZhjKFJBrmUGbbs
TF84EOBMjjaHrDCGFIQdxWkS97ymR4/d497HiGBMwn0pZpyV0eFuv2CXGM7YxL+0
lEIrfdrjE59CF0kvEtFl3qsc7glXglmlJHhxaX5NFCsg3VFp9kwDZgTHV/0FvtXV
vbUDxIJV7qQ25pYASEcqa3Wfhe0dQ5p1XQZiwaBlSePMc1ZbbVw2JDCYs1Y+G2HX
k17V3VMuRrXXGcYJePI9Kr41M74RiItpSlkwe0FOsj1lwgQholDw64jq4ZHv5RlU
GbpRJTDNg1wv36QVclWjkaY6toKsPcKYqb62teVh7+82R+9BaHyUlmBOo02TwDri
9e5CngRKinf7ZfxAyDYCRW1s0TZHFRetqM1PgQjGVutZfMSxwGcrq97vPrFmtBQb
1kCUAGzHZxhR8KQ0GZb+M49/JhyKPMn7QVerpsqSCK0fBC6kTOX3RLc3gh9DKE/e
4563jMVXl1TTKohMbpBOe0Y/jJe+03GBd4kXiXtd3Hel3+uIRteVvpOBfutVZzz4
1iVWsbgZlQbYmOWM4P9mvJEFhBSW13E9bvZtYAk3IhziNNWrH5nTVhOQYrN7oAu0
8PRNr53bTWuPRT4dWJssPYJ/ulMIki4xRi6UH3cz0K+EN2QCtvtwMB7mic+TQCim
6NnavRAIBqgWaYNR2HL1A8fbxLA4vFu5/MFeA6C7XdnPFoc55GX+JVD11F/jafD+
dKetDmFFeHkjrJx1zbm8CRxtTgmNcJMTUEyzlRh9RlkHvkZeBazsZRgPcIdTbLS3
18NdeRQl6kU18Yw1XPvXK8LhpLRlEWdfkuw8BWFcbRoswyMLtFeEg9f4GF6NYhX4
1R407H0I3SaWMrMlOrkYADNzF1R6NTxJVRe91SD42XSgHTg4KZmZ2tbN+rT51cml
zPTzH5tbDUJ0HWtr6dgJATcZyA48R2S+xTIotunBlL7lRYQnaoW3zKJZhHgV9vfE
P6eP9wKBukcaATo8GM92rjaM0SdCpF5pj0c7L/SFscuvS4gwqkcID5NISRgtPS9R
cK6Z12PZOX54gW0dUHwqVqpwsEt11dShTfk/+rNlFJz6bQBi/ewQZ15PfTkCfEqH
CkO7RYs6w9L8aGEiYZEvh+sV8iWloWL8E2i+bCsDLz0lG02oi3D60UXthKJW9Ppa
cIdEFhTP0lvhw5Sk9M1UcASkTCShCYfHpdMbAGh517RRXZyvYFn9nSxuovE43Tfh
Yye0LTwdeoJwwTaN/bNAuTnXUe/QsatSmg6Z00KUnseVQp6XjtydEQhRYotxrw7F
717AYelUkMK/ZRrlAi5g2rc7QE1reHRr83bZEhwhL4R0qdF24GByFXsy1QEYdJvU
z+lnfdUULoyEr6/frpUge3ZIOcJ49N9ehOF6POyDPLKcboL2LNgH48XOV6TwZXoO
IGltYxSWdWV4HJ1FgTffXdf2+vevj628nbua6NQeMiFf9ZQ0sgjCTwdOWl9HQn4Z
JdzNAZKdsymMJfbuYCiJ6saVxb/hCjuiM88QbTsKiloMELagXQbYKZjXencrv1op
yTrpl7z+FOanjBq1vhhu9wnf9GOmyBw5s3Gt+Ll3tdfsIeqQwHYup+z/aRF+Ck+u
Ohkq+5SRLs+tJmTjC7EX7DhJGyVYHI82JZq7JBrBiaWp5G3stSptsOwic1kH9BRc
rpF2EPkF0pSo6lEPMQYQFL+9Y1Iu8E00qeg/lMvF+4uk1AvAWygrfucSSawEOTp3
XxHpmDj+tM4CgiWNzVGtlnDXbVE83rSXHcJK10A2vYIVHBfbZWW16aDbVsZFeaaA
iVX2oQXm+cVhL9esmcvpz6xmmvI9IsQVepph0ZPowMx/0UbIjx1XfTXkPvyTXP/Y
TqVtbKpf6VlveX71OKEd5h40BjoqkIupo2SEhiJEVricbJJlj8+r4OsrYhDU2hj9
l3O56TR48g4NuybeQLhnm4gNNiLdyU0dSYF+b9OiVUfEvNOilfsffjeUPew/4jaq
Crp1WJoT51C0mCIjwYvi/VUW0aVFqzfogJswhLfU3zZAtapCnJHV2ZDfh5heJRfH
vqGsJZw/US1WC6uw4+wi4awedeqAwYzWLfV5sCh/w0/X0UMNekk86zz5qe8egJ8q
qmpX9QOIDtGfA+U9889gldwBuTu7L6BwHMY8E5lkxkGZ+0azDf46ymegu85Fa049
pGCiAG/nobisVGnkyXsbE5ZIkLB0PO8weOb1bcSlmc4/tV3UqO4dwyZwu/XoD4Fp
48oFMQ312KKA/BUyq2s3xjLi7ZqDkrkyYhKJw5XYsR9oQtgqqThUB0ggnoaWaMTG
uK4MyG8oRA9DyFG6yFzqefmVydd+yGUwGRo/Dtp+Ej1D3Yzy592aW5oU3hqlmkXN
AWtxVWH6Lde0A37PLJTu4UkCwpavvmzipr1La6Oum4FJWL+2jv8PlgYlc38MMwoS
BTc4rLdsnnQvagSP7AhbYdJqofQoIGQnmBC9dgqPkzTFzpKCA5QfVWjVaArHTpT8
3Q9UDJbJyIB853xZVVZtvq0+8T7/Yghb+gPj9PCa9ZBa8GJpXp2GbkJWje5sCiQW
Kkpzbdwj/zgOzKVgiJ9DVwuICq8b3o3TSsF6xd/nI2QftzNQ2BFeyvwIJwtIUuCh
TVfikTVjLuoFsmgzIjZ18lpIFYE2XLsMiMWbBvWlzgMtLA9Z3UgHOIJ0K+YH8XoY
3cYHl/gfDOD12HcvqAccf9/QsmIWRJsJ+C+px071J/CCHuPonqYohbJXj9aTt/q7
MWUOgKMduAjEqKUvnQpBDutlcg9sPTzoRoUbyPwJcoD3lzqFKYxIituwZjWnrnFy
JZEch4mI6Xzv/AbbWftzD66SLyzkWX7vrqUve5PMK7evyJhMJp2a7RqEeGNNQSym
cFXAViOV7P6VVT79vsExmBMHnNUJ8ba67q/SnkeGRU0DXPHTe2yp+47efMBzJ5Jw
GrQ9moF1azq2ltQNER1LL2eQJOOs0KZN5Lm4+eclvmc3hotHm9Cr/ALf4vM0dFM+
r/9glKuChsVRzEMkisyZp/sSpsJm72uAtJBoOyzhk2NGHnEQqj6V5yaWGa3y0qVr
5PXOK/kqbTQrWM1h0a5gpFQTKJa21BE5CZ1itXt2NYEtVoUupGpvFEwJhbfVma+m
Ug57iN27wwWY0dOGkDDgeN7Juplu6VZ24ojzaR5IMnalxDmGAFXwG/TVWMg/QLWL
nKojbY0lxJCrXW/m56JHAOsEZCw9TdN60MwyNefmxlJcbmwtskjZqhhAFDRKp8Qj
z+yH65b3D9NtlhcqEQkkMjRktsa7SzNRlAkHOUMMEUHdnw7k7zW8vb4tOp6DIZPh
HqISSSP7KtGIPJX2H1A4e8kC8a4Xq3SxubUS8DyDKWqrw5NNUZDpalxFmT1tDbVp
vklzXWWihM6Wc4xBCPYCcLK7ocwxAgSpmeHKHGg0NwPbSbITm0/+KUhgvM8mccUg
ESn7IJz/KcFGvSUzijAeIDpptydArcE+/oNiXEBv1/hjAPDZIodKTg5jR49azR/t
6n18Xj1SdZw98lq4xmCF7V/sOB3GSAT9dqNRnqgTH9NwLCTMYYOchP1QsybJdRZt
DQkEX3kaGOCStTrZ4o5RoyY+tMso5o/TMh3TckTaGlL7EC6XwmWGzTLuArQaOSz+
v4YeAjqTEhlNn3qdGSvuC2mLZw9fdr2J9ICZad5Z6C2BuMIvhNAj2gA9lOyEUMaQ
xU8HooLwprnkmCARu/4qP5WaXGKWpl4uw/LVVo5zAig84DA5R2Hr7ay4Ln/+CLYZ
RL0xspjPL/oXHHA5moCOxhY1q0Hd9FfacGlMyvx3y73B6jryPYTCV36Rst7LP+Z6
ZU8pDgCtttuwbTzzWzTP4PUTwuL6qXi8D1gsNrrNij+6pZ5dxbvOAtF9wgksJvRb
tLTnbqd7mt4A4nG6bMsWTcRJd69vH5kTTGRfXB7DtQyEvwrcH747LBtnPTlAbW4E
Midpf0WxDKClg7azjMzyMe+054UJSa+jsL2a71L1xIZGbllKwLPa7Pys72lnN35g
3Db3k5d4o45BPesJaKokEGRZAgkBx0pgOmkkS9HcsMzNAqMlSCFhQaEjR4+KN7ea
bcdOwQBV/9ptFeS3/R2nOTmmgKEW6v+jlIJCQcZ34cJpuXudTUMZ0u1M2C94AzDS
wjp/77J3ORKEhDUXIZdVqRdm70qHUEDbAEMJNLwAZ2OX9fYEMJIOew/xwxSM9GlP
gQ3zYbWxQ7UwZjxdplUOqAmmIBDc8p+EWVJL8Xh/Rcka6Y3jdwQoBuuQMSTKPiKj
ov7M9CzLT5l0TnlKDSm2iEQpMt8DD4+Z+6wHdiaIrJnPES78A2xlAgV4nAQaDwnq
tPmw8ZJJKVUTBBtlMu5NTNrl6QA8m6K6ue7uWdqyeL9YhQpQC3sQQl0lDamupxtM
2PQuI+hOMotQS9W877EIFEELcE/7d2iYYUxHugqn9kw2bf0NyORuXfXtSfPMmOiB
mQf2HPYnStAqKz8TKMkr+2vAZRvloBL3Ojo7L8vbcKbh3+RDh5wTS+489L8phSuo
GAceJMkqiWbtJJYYi5oZcr6d9nW9BHIg4X4fTeyb+tGAFbg3z6Ygjw6tBs9WZlH5
S2p7wRUwJO258cKIZOQS9uBGc+7919ifU629sTflIY6dG6jd3U2Es0W0qf78+ezY
/xS5sZbmlh+NIwzex/DSlBc/j9I3RbUEAaTjunHllkD/7OJXEu0j1kr94KtAhSN0
kjimXSV4gauuT0wOQXUTWUo8eefX/SP2is+pAWICO8hi4KgdQLdDWHpgQrkanPAk
ZwWn/3CiF5VBa6+9D9/T89h3er62TNiN1HmGg/ybhijoQ00STWS5idZUXZCUpIbw
f2c/XlxQXgM2fFI6wPHyogIUUGhCw56RX8B5ON+oBHWcvLAXDUF0PSvjYI0M+CSZ
p3i0Dq8YRQZ2Ad+i3RaD9VUzEV6DCA+9F+Zuw+/vdaZ1XOXf1MP4SVXK/JatsKFY
xdmjjkG+fHMU9KHfi2DNL5K7fb7cb+PxN7FXqFIYIi9acTgOihBAP6PInuKcF8yt
ixnqXp+fA8yA7WkV7OHAPc0q2GT++qCWuSsFeK4zExGNuWlquJmFnX7MUboL4Svt
48JQOJKxG7a1ZjORcqg8BBovh4rG6Nkur9rfcEySvHkQz6VmHbBSLJPtnsEVFYPj
wT96jKBgF7KcEnCf2uFaVeD8lZAOfdsNki/SLDD6hGLUidure0nQJDZyYuFfyGMm
XT45dkgatjTLDPwpYgWF4UIFmuiUHOVAaQ93XA1+EVpJy2Nwiae2fW6SAiq5Qben
Ec7Jz1SyAoiw+I+hT2DBiV3EvUC6piQvsGJ81+v8r1vMiZjYE/QFczSoN7EPWD+E
Hu07eAg5djGF7ri0k91jiDZyV/BKJuHRx6Ep6gb/XiCjq4DezoLFAqSFbbjxYIy9
syqERvHu7IBs1PrzpbVyLl+ASQwcqtDv//95PtaOztge+98ByG4gpCs8d1dFQRWs
tm3oOxb8eGKoGug2e0z8RwsFPNoV95+AjyceIhQEWd7jdsygL/BYm2ZD3O+TDVdH
y5yF1qoFEDgVTB5rb8jH0Vk/8h6Q7NMRtjwWgVWDZKn+Dq/3xNGZI1LJHeCFc6yS
C7GnP7OzBsNJMT1NFNyu0SeyWwPvXHJkuELK7QOt+g/SwHSGRdWUQBYTBJX56R4w
eafEec6+g5K+TlmeLmBLWpvTqbmS+sUsmmj/AUvDZbY8O2IjziIiUcueDDnZcJUO
Q5DezdtZhQmUqTU6CTPpMZw3rJCsm8PVV2Ancp/lDsj8D3E783QZoK+redY+gN8K
huex4e24nl9Wu8T4Vu5QKxWOV7KarjNIsk/ecfkPv9hBvhkM5Y3/yEIvnhDSMQrn
beC+YdvMQeWZYmk6VBVgTKi8UfI4Jn+vQalVM+9dnDyC+Z27aH2C+PmpPTn3Umft
e0siiVjJNwP5GkGLLn26fF8Ypxlt2E83/Vr4w7ZwkxbJXJaHC5Z7Qf17AyhJ8OGl
JJOj9kQCiSnZ2qj8MmKz6swFwaF+loA6fZ7fppIYeVrQoi0VXfb7xBCsfDWBg63v
cKiyXPvZ+8u/cD3h5dqNE1Pt7yVd29w+QQxg2ww1xoso+tC2EUYJP89Fgn7wQ0E/
nqwspY+E/EBjX6dp5b1634zq4af8wAZ7iLoAEt7jR0/OQIxlOo9jRm87fF0BiQeT
KYwRgRLG4XCvclKOEYepXZn7rxmKyHfRR7i5k8qjSVmOtxEo34lrk2NNta0da6Ra
TM0Hw0CQ5O64ZMne00aY2IAl/NXc30J5LWHyM7vnbXtTpvoSuQzVfWjtS8E0ztyX
b8xovi2F8q770tmBivpbzMbXIUpzBZIwKvTs7ZRB5VXllWQOmOQouTYu7JsY7wPZ
SnmQJ33+usBfpg9uYzYzmxQnKtWWJdm6J4INemNwXMbzI6pGFvur+V5YAXivn1TL
v0G9wpaHEL1wGVQwrCFiT2tt7CpVADBs3SqiZErh4SaVckLqVUKgURF42W0ADM87
CHOfpbg9FBoM26gJCRTKuDyq0tFkQouRUEbEBVkk9BBT9+FkBwLkA0b6oiMuH/Hj
Tl/cT4rOYjnuGwaTNyhz+OzlLtO0Kme05GizbgpDgEM69fYIMeL9jIOdycn6eaNd
dEzxbXRSCobaVZQowbxIrdrJV6mLidKq3M84AxueW8v0FxX969/sufsP57ILvabU
vPeGq4BeC3GPpq5VujPWD5mb2mENYt10YiS4VV1obFM9YV9KvhAmUPGAig/KAOS6
f44AcLzk2O9Gyy1ejJEUNHb8Zfpg6MYwu4Kq73jjvhumebuDJ/EtsG4qAhvywI5E
FtyAPZTAOI5HOWqeVogT13tG+y/8aFCcewPel+sHWruQLe2oer4+WnU0OM8MC+qW
PyTAzMPPEtZ/VRX6yxIP02oZ74qC1qVfQFNyU2vRBx/lQSO/bROKAE4ORTpEQnLE
1yS9iP5LRqzsvU0JXt82qXTfr9STZw8CXFQakvRkQCcvmAe7PzUmn81uCMX+WanC
CrjNHX1Jkm8Xn9rNoMz9m0X63icgyIPHqwIQiThP3mv6z+CPcwNxsk6gVCpLZ/2G
2R/pmH/tW/X/J3Z0rbvihMMybikkRCH/qCq0u3PyF/MOELsfKB4HgByRd+YwCzuP
gSxP/7FyAo6uTTmER+AhYAHuUZ/7IiZWpGizHBAdISSo2cQja3XUFYdGfo5CMdjU
D5PW81iTJia/dCEmT+7HRpLXRXtRceF/qCuWESFo1BYTZwF3LbXkOOi/GZ+NIeMy
uPkSxVRSIShZ5uRhG1b0KT/ZimQz9IxD6VekxltQR6A/P48xPqekE7dcUZpWUVJB
WAvIR1VaAwdyVDG/Kgn7ShnPt/HYaXnikU6BIbYtpYQBkPV40ADRmaBRm0ixw3lU
QxKK17cWWMjWVVEaSLtlMvLTnaMkZc57b/tSa/L0Tw79ih79nj3c1XjVR5D6uTgx
KebwVawMDZNMLEfzcpburWCC6cgEjK1audia7jbSi6bRDxMhL5jzmVtAtO0VM5tW
lMDhmUBVXOZuT7CdacMigk7hQXPZgDR952c0hzEB8hQJdwIhs2SNUtdvOAfbBK0U
Srjpc2Xmx6rnrJKsS/mzzXHcNvQTz3NS0W2tdQzJ81KYm6MyrQRdPIqmv8J7gMnW
0OMYtRBXdyqK12iKjoZ/4tzy+GQC6+gDM+N7sh3ft1Xg12Ceo9gBWlqKhOtPHrR2
8wHMJNk2QyBU7/DoEWVmhHgQ2+VSum5X70MrFEYNTQbsE+LbKvv7ddKDIefld+/v
ODO8+VIyGFTioW+jMOONSArJWs7Mi2Ex52ayo1PilXRCHv/c7P2cQBftaIuA8dzZ
tcgoXTHdA89drJbcqjmx9zptpmoMKVi7zrptxHbMVQVoTuowEmYAkS6e8XeBzMWt
0MCxE/t2RVLpgcKCXrZc7tRwFvA9AQ8POIuHvOOkb1CJP4E5M4lC041+rNlV8Aab
0f5iuavtuK9gfIsMjwTdSsus0az+O9ZyZsBA2ONWkEZ7RW3Uzj9uLXOk85VMqNzr
WTpiWkjr86s9PmB67KZYc/zWorz/7dCS2jQHpxfCFTbb5rn8AXCnZOkS4E68jsm7
E5k+is/HGD+iQDjBFfKYO3U+H2oykwGKLC+6qHk2eLqeeUqpUFrUQz/q4LXIvIan
9oPsyyFKgqUjWPzJC1hH7ae+Q9fteMvqW4lYTl4qAPu1kSY0OeLSKO72ZhrTC+cN
rqvOKgDuC6pCigA88CqLwO9822igi8pbhqx3zZnWMMlvnGP2FjnoL+ps6R0jXElU
E5UKZErskIF8XIt1UWbkjNHWlsZ3Ssj/fL9grTCAXGXqIHxbL9JxeQNCBbtuqoWO
0TvHHbCEbex06TqmDS86F6Cf+vLm5fcVjGvjpkgRYdaZrjAZ3QMmpbJLC33vwSeb
iyyTxo/yyUkUWhTlhphs9TOWXCzx+7+Il+4FwIWXS1qayh34Vvh23YBo55dDKMYd
yT9KsDd5+WG/LxO0yaXc/idel/c0067/Hky+w1tvtR6IhbH1ejEmPX0MgxdALB1t
Zf0Qu+vCJza8tgCKEU61Z9Oyw4+2Uj55WGtxDdUWs5L2aZ6PICIInfkaX+6Ona7o
MLgYHjFlhKT8iSCqysxMF2bUS/oVktIo1SS9FKGMRyXEGYNpfOJuDU2Q+Aoae8yA
V6okQPVxJ+IK6QGQDAEffa7m5SPzCg1T8JOTCqSglugHOglBXadapcoapF3a7Npf
jFhyH2KGvnHC6ID6TyiF6C8HKfsBg3WT3I+ETORbAsU80Qik9j6r751lsJbWsblX
ZbI9nqlUzINkb5UG4Fj7OWFMg9gIMxXuLWVv0gL4eFskiIUpVfplBOWqh8y8OEa2
HL4/4LL2icUR91NxOSsaONSbccmN833wd/Te1j3cxJEKbAIoSz/Sx/5fwI9e+qnd
CebKEGOvYySpiXHlPAItsy4lPE0TwHiCk66/2XpgS19rQYAVdINdyJ273RyLThI/
fqv2vei+1VCImCQdTb2bkB8d9DTyA+3oVYx5YPKqmsmLN8rYN8o4Jxde38qAjz1C
hEDEe5UIS/Ncw/MGjilH5ooP1bNCcoKMTxwYEfd9/7X9ItxWwvvTXLfu3pV7Vb7V
AV7N+kRidv5UOW1Np/9DETN4VBqanSmsjkTUK3fmXVr8hydaTXrQAM/ekf8lJKws
/axIfIFeROdSw/irB3NKp9P/49Vuhv2rp8mAmQOnkFyLr4zbyQ+ksBb3WBnNAMC5
aiuBZmfXL9/bkYzV53BecF5D+QYabbsAuMeVs9MIdp/S7VhGl9hWLWxOwnR315a3
R/kQ6lbJTDebeiUhrwg1mVhcZfO1ODGJ8/IyaWHDyI+8f5vHFYX9OVJrysIRLrvL
AzlAKtGf+UEgroppAq2npty6RyW2JnRT/c1795T+h0z7HKmX99epvAMXoBIvbXuQ
N+DuW9fZKr8LFf1GqaA1ahRsh33JaqULVeIdfDPFGckawJRmBN1VqSpDSA4uxLpM
GYFMqkdtwYA0UuW32jiCCSQ7duAJDruULZnlzKlrAe9DoP1+nNu/hcWqgYS9nCbo
Ag8Cc1XjLufTMYvnshIfRKglRnmcbkzl0jsbqi8s+sXYsOsCFrQi+I/TaFL3w1sE
tSmtSu6d3rhfQM/TDXYZxtD06b2/PuIbRkHZ/+L00h5mEGqZkoSxHkRLenrVYrtT
n3KSzvuBoXZ+bvChu/JLGkeTWu+Y2f8K/srfMyo5fuSgVR77IAgBv9zWi/cpccP0
P84/kusr+LrOm28llmWU/27BST7mesIMHmEckDFzQVNo5GZLrH/lw+fita7GZVNP
rJyN67u0mXrabLLp3KImwZZieRijgii3EiLhWyqZ0JUfBnqbNguTctxNUkc/c91L
mAxNsMmNogAD4LKoe05cSrNtxmjHTg7nHV8BmzuPDTPXqTkn3MTHQo5aH+rBU/gA
MCWp+flTii9M96mbGH6+gNXvgCxW3VaA9L8U+s83Mfw66EbxAEWHchUL4bdJg6a9
wRBjgF2O6heLT792Ju40HbtVDpO/rMnc0T3LqotKWMV8+LBMd4ZdOcgs5A4ZUNZT
Ckj5hk7WpSRD5yL8bKnzMuYpGFhMQAKrSTICGPWn9fkpVbMXNcqDlrr6VJdYzQOY
SCWVsUfE3wkgr2klxYyHgBs233R+/h7qdrXcklx8tZgzCtn5NUQbj/U6iy2Dr9Ha
7xj52i2Ab4v/NkNEx0kpGuyhmBA5w/bhjodWp+vcMJOrkxH90tRIDfxFQ0cAxyJf
vFHO0qE2owYsu4N5z09tKo1MRqUW+UmjHVtuDP/SgWbaOKjkzNDVO9UdSg8wXPwg
ebuZWSlAL/jg4kvu5/J0ega66ALBZ6zAD9SeMQ8Pyj1I8bfeckLiOFugNwfvB5wh
7Z/fwCNq81CeeAhdss4FhhzCvai/MsqkFN+N6KmIOOsdUtDuiejo6qJc0czF5M3I
lUFZu871xMaoMFNkX0B22tgUZivnwXqFRGb2SPksHMC3GOX8Ws9ehlHm1xWW3OiR
F/qEL2lJYGNjMSOzGtXeQZ+HLkktxWrhvT289YFvWi08D4bLyDlcjwB8vG02OkBH
kH977KbdIXJroAYWeHILODueDJBiE7IE54/SJidWKh0DzOejCoY0fSs92MY0zilQ
hrCEUvjQdj+wNjeauY1JjFj5Bfc7ShomQP+Irc2QIH3dQOMBu7OaB9erRqt1MnPL
Y+f773lz+OXOVR0Ak7zZCKvvYJYdBN9pAgE4aAgNW9rMBWfw43TO1PqwBmwNXjku
4IEYaDcqsw+6YYtYIq3lEbRz2AysEUFtSDpmlV1dNNq7O6Vzyff2+Tdw7n+j//bC
Rrw/dDu0qjsTY1fE2rWy8pPTyWhexOtI16DZASe5FhkcEe96oHRvo+NU3YX8im/O
Q+d9phYcjJE3LxlHefP9CGDsLI54dKQrqz2b7o5BsoRWZOoQX55deDTOfjNkg5r5
rWev+UhBlKfWXnDtIpS+qZ+TLzoyIY1jyngZjTPXj9r2qcrE5PB0xcC58R1iR2gL
ShSNUU+i7vhjcTZL8sUMGIiBF6uo4wKwLopl7nVZfw3AiYIe0U9Q+S/2xQ4DKnK9
pEt+PPEs9EC0QhwXzH1I8PitPtpvsm9DnNBW37+Oi6WYOqa0NRj3ZJD2PqeIPrB6
RBUwaTUUqxRmQbW3P+v69O0BieWEz1UzEBt8MUUTTfi0LrDnPDDvxJ6PFAgvodUt
4q8zL2GCGlzP0zWzvmpkA6cxjiYt0aMN9b1mgt/h4CwpK8+6CAxQPB6g+H3KiUw/
WedbaI1Fe6c3MVXqNHQLAV3DLwhFb3IUNtk/QWVg9Fh+WFvqEZLPdC2zdyH/qG2E
cQmZVsS9o56fSbMyX/+Kai9prK0sdaVbbGcTh7DhkgVeCPVtzlC5UAZ6PqbHTiJu
Iwdn88Umm9dvRZIlsZIsDw9TqjzeTWqAS8Fz7lrDD0B2qtsh5AxItJy1Cy+XEOw4
+8hlDoAydmAOymFU3JgOLVqLq6G/Su1mBfaOHQLcyzXVzmT7yeFip1VkrDC37q7a
+C0OitFk1OfJq089GI0nhI++oF6umc9WqvjWIasmCCbayi97PGWb6F5yEFrxkdMZ
JZ7ZLBCblqtwkicClP9QwrtNTgcnrP4uKo/SKzHwFXDUFBRLYsQdZ1r1L9r7htVb
bnz00bcSioc/ri7kdurHO3VrTIACeeZ7c5dOfqlhTIA2Z6xrhzVTJTUp/TQpQFDM
rvr7m1MdjNa8bmHUf3Pi2FY4NG2lkupbBBHuzQ0PBGqmtsfVJJL9vqGmlf1019fM
OFTCpgh85Ky2GBaKrHPS78H1QFCS4Uu1qFjIflGZB1xpQZXcNPvNfm1lo10GYM61
a5nUX1OT0eGx3KbzDlxoi35E/lYXXlU/InaxMoUAvB7owCRF/jQ+DHAx2dV+IrhK
TtWY10SWYG8zJo3xjYBBofwLhMS9JtLaudZczbe9kVuy0MLuynKEbfVjGbALO7dw
ZxhIHK1WkgY8LZXdv0uSM/96JJBF/WU+XS5rUtv0CA663F4Eb/+f5H08MPmI0+R2
0RJfujj4PNBBd++mztuRg88u00401Ucm7nzmi3EL+W8KhHSSayTcEWKAXP7+fYI+
0n3UZ1B6JPd9EIwugkV0nPUyOd05fP098PjzRVGrZUxpI0cY+L9Bekbt/x3KQO25
eTM3IoDfNMGiSLNTZ1ngV67+uA4/nj5Zq/ekIcDcKFSjw1z4EKqaQ/Ez44FGBo8G
E8il1p0sD2wSdA0XnrGGdsLW2SOg+5hh57x68Sb2gFBPDjTn/vNLLJbY4lR+e2ve
0SnQA+TClAYh6Si809OxXj2CipMV16LI6Xfq5Rewhaa+COQr16ovhOOktelPrwrc
FK8t7tvRk7LKlki0rKOGp53R39JtLkJX5IVAmdZrhGWG2vP4uQoGHiuSs0HOgUTO
s8cNiDSVFJy0BRA4kZXovJVwmPY++Ur+u5tDduOwan0KJzx32+qugq0BubUSQDu3
8jRYoSc5BSTuBzaH8sbbDcPrFH70ivwmRNk5UAx+HqbHWxm8DIkua+kWQG1lF4tO
YZIcLcDtjGofM17zsNSuZGq1bVS1RNBK3Ns7dG2BT2f08UH1R/Iicx4Fdfsr/T+X
Nq2msOv03scS/agedNsGF6A1E6p6Ebjx/p50A9LDfnehIsGKMJEyXiNfdrfvJfgF
maZ1DG76oOXxbvA52ry5jIS5QnBp3jW/afHNW6iOI0l86ZI76q89d3XhGJR3OlMS
cAwxFv5FSHC9Syazs+LUMMO4jWMim0whT+OhwkGdLmzgWFSz4F4OS8TkLL2jGdJS
YXvvk7UbZbQqiEFv5PCCjWP7hLA/5huImTyP5n79gNVhdVcPCZnO0vv49dWeasNi
i0SF4UR8L1y/2k5HunEsFnXPWSgMhNpKH3DrK7Un7QsUUK15T88mnYmsa9WqtSOW
foEt27xv9wMhbpFm3OorYlX73+/oDcCXrWC/QdvNMizeGSG6k+hfCvsTB1a84BBG
AIYQk9g78OSsazFP1qQZaODFKH80sus/gIEuWXxBwlvtWhVO0nPmlJqh8oRiddzD
a1ZqTOtDUoTGSzMdk7hAeZlrfU0RI5teuuKC6LXUI6AIEkoQn8Wb9PhdR2RgXffg
cVXaLaYaIhQ98lTjh9RJVIkTMk8pOmNmCHvVEK+s39mzIbj0I7Mlrbfc1or2PJTX
h9OfUdxA1sQZhVXZ/x6tmSGtKLxMbyoy4A/AA5fIvXimQM+UICmA+vuz9iLsiGUc
6BuLtAiNwlbcaJeJCcyhhId+cvqEEcHMk+u2WfIv3/S+Mks05vJW8R9kuRJJqtqd
iGlE+SWw+8Jd2EG3eG6jmD0d5LalHJXz39MAT7h//XsAfWpc+oBNwwp6CCWjDoE/
Lgj5esAtm2EeU6Q9ksa/d8ee6rzAWujg+pSaTyweZ6bQVIbMnMYnKeHST6VrcV9J
W9UmSWlX5ZLbqfiK+ILuw2pA/tKL66xVy9AsPTtscbRu4az8bAJfvaC7CSU68469
v1BNrm/UMEKWLu0N3p/LEuTFoW0NsUJn6Q7BpTmLTtkYIS5j2scRd4ZZjyY2KPIY
YumX7spgoxwk/JZdMYRcG4ydoFhrIqhPh1z83EX5vSQk/756QX8s3IL0x8uwYOem
Zct/YjQ67zz3oDqXFM1mnu7reKTrW4DNv+xPjC9gvuVn9XPaFBNb4PHOUfAJzYMZ
Jfw6ZThG6cfUIWeMTfpXt7WQNFW7JxX4IlR0Diq2vASE8OUJ1Ah+EbXidPu6ge81
cWymQTeJ/mwuAAs2Uma/IJ4LAG7jAPd2jhahYQVmykbNSEsfwTAU4lFpGN09BQYN
S5KlPzWIRYfKmsKHc5iUCuN6+les/kvwZyXfXw4JT6KvWEszel/iT/FnTHzXbZ7G
z9q1W7X/YBEbPsPt/SzXh0op1hQzhWASI1nsO183PHP/3B05gaYajqgcmtjfXMSD
DUNq0aI2lzKji2oqhiGJnYOeF0V5cCriboJI++slPY8s+gAlPgjEOA8hWd9WMe2L
s2b5a3ufn/4ISBFnkub6lOA1K3I8+nGmdSZT/bL5umxhfF1iDIrWzKwYW1SzLB69
z1gqRw9r2sJzSPjXWTg4yk5J/AlDo90aS45qiodmBHkIbD/AkaPcckSmhzRsZ2od
yQU44o+vswmUQ852PlAr3Lxp+m3wVM3AVAgG/lOAXvto87oP2OU1oUwzZnHbsAGo
e1wt1AanzRZz8L8OhDS/HoNpLVV3ywajb4KSmitO5Zrcm5xJVTU1grbgjxdSb2ar
QLbDqPHp2CcshF6Mdf0JVTgyPKpdwH/BC5TogJMv71FRWXxGuCX4ODtsD1kSZ4HL
AyjnFRfzUBmlxxZDTy4380OEBZtKNJxcOO/hjQrxNZps3HTv+L4FsMikGXjNmaKN
+nATzGdmNGssUe6gYey9QwoN8Hj1+U6971oLhe/ack5ZwoBfC58/LSay4JDNfed7
w07X/DVX+Nl3AEZTmwxR3vn24OAL7/FSCl6VWXOMwN5XGNASC1eVBLAsF2QziC5v
HFgwWUwauWxAfcGZstcAv4BuXkPyJ+5sKgVg4oqwC0bruDw9qrXkH4nxYM3Kff+w
cDZL5GRdt0ZwJmGjsGNg7kDAgervbTsMVJAvmyUpji7wBWlhak62jBg70DbzfpE6
6NGc8ATK0OXM0ASMez5yM7EX6BUkmTRTPUxTXVjhILd/RY3z8PK9ki9irNLsQg3H
7u6irIsKnWr1yVWOif8j+1SJqoNOTzhYvz/c0hAbD76O/HKiC7yp4qJw5oElMRpa
qoLqvwN0zEuwpSfObTY8RFLsTJaiuSz78lCIaOlAp82hel9n7DRxIqgOzO0zbMfj
R/xgcYX84y4b0yJaVun0bBT9xAjfmxEfsYVdex2MdhUOpXBZaU18RpWjAYhhOpio
f7Bl5RT9u1ULbykRjejVN+RTohwwI8XJHKJoEALBHxg+5GpColGH1gmhWjFJ8Vt+
9sWOIYOhmQmgHftwgBieWN1fU36qcJUGbKYu+f6P3wyUQS67zuSBiFG45CYWPGPV
ur49drcx5zH7cbl/bfmHkwAhw6KuQCNMjxDwPos3WsUkUv41yd+pi6rjWqfFlIAG
jRRaHRCHc3Xb/DWnUwXEOc79vG/bGa3ykPoYvhHtH/B94htrSGXOnH3IIKYX7HjZ
B1bEj3LqObx7uKVDi0fw3GN1qUEKz6Tm/fvvcYW+PjPXxx5tJCe/7MeIcDIXcdMf
n+XO9amzLppDo62oZcAGxuihjqo8b6MZTYLnkTpdDA1qVFl15+edvdW3SomX5S+p
Ohj/1ftJjKQDe7kb7BXP02AiTLH3tOUvUShiMabIoYnYE0wKdw8kKyvr5qqkZeSS
WLpTNEjiOoFGq57QzYUFBG9/RlXZdxXktYnaV1fmfq8/shP837Bnzm63hmk4q5hL
uWGpWASVDWfJbOnbMhShabgxRBb3o24qlAvrE3/KUYD+EDuKaKN1JEDS14D+754g
HkC6nlY+r/yl3ZTSL/J7oTzsvm1wvTdrBqLNZOxpZd26DnhAP04m/Y8U/DYDFduG
SQaWZ9OR1NWM08z3fprFejC8zoT/IG9qq4dv/ATbdUzgmyMOoAir47VZhNKfZ/q1
TtEYskGVbCCIu03Dc6feCTdQX2jpxYz4hGW8210U6S8xfF4dR3dpbsWJknm9q/eM
wJSpkpJ8uZDXjEFzTAatwEy+d0XoB3lKrpKVTjCAA2lFdSYk3+lFHam4oxwUaeTG
6GKSdxQQetIc1Jk2XET+F8b5IEiiyYHu7xfv2XHeKLKA2rK/rOZEsJMVMdUyKc0p
d7Ew+i7yTLB6c7SGFE5IJPtjAXvwsRzeRVq6rCkx0IJW3Q136qwyK3JpfsDdIJwo
/VPsil3lVNFwdzDUBOPhystrmKNg1QJt03TEGIQSpCjgNMAHz7AXi37R+1eMs3sq
0ijakDEPR1UeyxaxUyv/SqoiVBfEMdXB7OA4nSZY9eY2nTNtmhiHpOwlcDaJ866g
uSuAQUJ+DW3p5itNWPX2tZjKkFijz297IhZHG1XMsLz8C9Oz1+cDD+q/LmFMQPD0
0Uw3YWGOOgx63ajEYaVSHnju/6HwVEq8Cvqcs8TuZC0BJk7uwdIpi6zqkEn7w3ju
HT94Ju/HxW2OUyQ7l9R3Sb6ckmaj5tYRHp9HmKPe7mEhdRBNNMxaJNPUkgcuIakI
8azl3BAbiQ5t5vpDtXbQns2rOq2+rOFRIKU5Hajv9HY/eF8jgj25k/Dw5SCJdOEL
hr0imxon1aTuctC/jQMy0t5hbpoT1UWp8Z/W8nM9S2mg+eF22cyQXWydUp766CMk
k1MGGQ73LaJZ7bUOwXm49Qh44zzAJNMUY4Ik4lIhs8Ed2MpFmy1038cZJznOwYjX
uIY2AjszXknY1MXrrDRi5vMUVS1GQ0H5nZKeT63Nm7ru38KyX+y5SoQniZDkLNEj
PxtRA0FgA8ZWuDi13y1kvp031VxOckfM6Bk7ZHKFI4NUbtikOUSeXOrMne/AacKP
vDEE0CjCopDKESI+XTSQ46BJ/7ounckvV0iWd2n+1hbOjCBNjiYX8c/KSWhhSTMe
WavVVkJKod2J8w1bX9A+WPbjEwVt/dTtfXlRQhuA2OUdxHuO6/WWUhYoPjuusKq4
Q7PInAt4eXaK6M/WQFvrtLzFVlaqHuKyw7dMg3DofgxVkKflGvtT/m4cD0G6kRcg
aNjdPBQ1noBFL3yco2IjT1LWdrFxaDpBEDEk4reYGDfbmz3hoXnfleoxeodhcLC0
0MZdCtM6HCfv/Nq+0r4lBAvy49+Nnog+3JfoWTQBrGkv3aveVqqHSmaNQdQfSge5
EP0dNGJNWjHqVCFsq/U/uba/G0bRVQBVbSubbDotmNlgdJ9fBHQwYwNgROZQafz3
NYcClQYrHzCkK5o8RtiTRPOssl0AMX/cTB2xIUQL8YK/ZsIzMgM5xjr/ysu18wR3
nUxCpY8ssc45M/GjhbKFoZLfZblCf4CTWQ3sOFKMEROKTLLbd5Z3Xx8ImXk3fkGr
Gg7mvFH8KTIuGSXUpg2AjnSacRfc9rmT8EgSTmdX0YH+GGi1V1j29If+9//TLyJ3
Fu6zV9W3D1yY0Qo1S9YEmLf0ikYjay0wCuSXrYD7DAlkmULoxGWkecXzmszN5jr/
tGGr+Dv0D58UnBwIYfaYB7Od18PZuLFhmgagHQ8b6/jjxTcfGbClilY5aluOI07q
fiOxkc2ZlmCOTta+rouyrahhCpENArhTrSJmtolHUyG/zWO4hkK7tTxHfq8cfKJ2
dlu+TnBc2q+XT6b9fZevZLBl5PIFVqL73hp8tjxwsiswFGZ0DOi5CNkQ7em/Dow4
Gisz27d+H+x5d0Y3EPakEWjwioJNMABgnU/JKmYePNkXYztzHR8ZTh3QF+YrrzF5
va5/B4G8jg5Z3VyKHQYR9MFtaT6GdavWm0Waz/TC3S3i9B/oo64gpVMJ9qP7Zzce
wtVpMtyC15kkwUMNDUbqnz7fl6vx9DoHmpX0dmjJyG0l4MPKCSix+iYpsNaPbMkR
gY7iH9KceuKvi22DOHiCAVc+hM5RYxv03JlWEG6UluR5FOg4y8Viz3HMWo+qw6SB
rPMkq1Og8ttxezEsfUeMSvttxvIp5FiC7IXzPX33Zs6J5taYhxSyLsnrHk3I9vNU
/WFyIAL+u1fZXDP50KVp7Wi1LtCBx8n6U1MkNFm99+JZ7GpkRGkzoMIfybttkmR2
HlUdQkW63RapvR5S5eg6dB1udGR3mfnxCTF+kQSyBEnIHR1cHGAiXFLkld6Cq0Zn
bbpGmPkrv/CUZrTn3bDXOqfVSmaZUQGR9aZu0tTxDuFfO2AdcVxGT+yngUZIQA2t
zPU0wsz3EeXutRHQDwX0JcfMdGCzFPRqj25MxSkq02cnRI7MtziBm2xGDsdWU+/K
g2yUsawEYll1IuZ6pMJY8q0S333/q6p9FR0gXatd6ekSh66bldtXUUdojnQC4Y9y
+N96RvPuKw6kHjLgwUwaAE6ejAAiTYiZ3M8Sg/Ey3GL8kWnVbU0CTwiNs+qm5fu+
zRWOOXDUyiBnZHQHfMCMbiNZGwz0yvxBm9wQsMDlAop4YHxIzvEzJhiT5BmGgryx
46h1uNtzRrj8FX+eGeHt9D5sUOqg6oLpqx6yyUhIlwBaX9EgxrSTRmxnI0Ed0Cdx
PDx8t3twJwJJGvxRfyJiwW7ziVxBOWug3pr6ElMoKvvLagkoZCoJ+AZqZmoUxvRt
DMrRUrKDeH1Ml+MENf7aoe9M0NUmdmF455kxfNsClN2ULQIUsigAxXy9/xBOqwwF
XAa5e+Bf3oeSxi/sXMWcKffjCM+/fxbfzY1WVp4a/5jSRH9hqYmhMNAmRwje5YOs
ryEN/Jy/xV4/2P7OvctA9vpd+Su5o2mHIs5m3iXOeM1lQBQsjGuKChPJUv7i7Jf6
qos0SQ3PMlb5PJHJR1QrUi8ot0Q8j7ENl0idjM2kFkOYfgWJFHn11ip2DEfm6p8m
6HL60p7elh4cm0wS9LckNst35mo1kXa0HtufJ1N4HnZsxkuM6b81WzBH6v4TJIUC
zW0jzBlaYdiWO3Z0iKaePWm0lLl8E5lT3c2TNfPP1X3JkW76FvAGeIdg1n+95r32
aarWRbBhLitmAoKrm9CzfTIcsqEptSWTBZg5kvXGN6xflno7lAl1c3PIbw60Bfi6
t5mXtP8PGc1+rsrdN6aNwn/+NpyQuaEM5XDxQHuoshHmvi4S7jlV5N1eFlUo06JP
0Qhe7jts+dH80Pbe6HvFWI8v6MBHerJGXvy4nPVZmH40onqk/bvTlYeyZBhwnrkH
aabGaNJABBURkYq1QAqsDk/Vg6Gg4v52MOE/+6IbcwNloLtW37dXqLHyOFJsCI5q
iOgtVhVqxMhacas/qaFXghkYBhvjZXpGzHvo/2uZzOf/xG+JaX1i0mijsv88S/Ng
x6HZDofZ5U/+gqfZIRurwSrg83o2/IjtfNKIURNBY20MvyYdvWRlnk7V0L8DhYZL
CtoEtIf8gQH7lmLNd8R1U6LbwUpd/BYvJXv0lGTDkSdrbv6dzIYanDN6GfuNR4oU
3BUxafaoz4enzLahKa8K32lY0STH08/OuqSVjz+kgje+bDMhdotDHvyh4IMs5VQJ
JOnWcjU6FQkbAEZejHUT/S5JAOCYh6pNL7moFJ9gT7SoCsa4DvcqN/ZJxV8Fgszh
0XhD0b5x3A6icSKePnYcmp8n0w76Z+1HUL8LH1NrdvDrCuov0fMJdm2SMlgetf25
sjiDFc7di+g/HbFFyHYoDf+nsOhImzmS5c2Z60h+KtVVBIOBigxzG1P8gzP7PMkD
d1EUojzioJRaOZB6ToOqgK+TmxPViLevpXKRrr48ekLAcmMeJwk5ENadjIUIcVg4
kvY4+dQ8mYzMn49TacIDrnyi+2mbsSeVFSXxSugEOwehK4etzy0JUCVCQkYHWKES
nbP3SqhTPaVNYMXLlWYqHXXlmZRHVAMq+A9Czsqlrt8jLwg+esOWof4uUTkWdSlH
DFwlsPlOizDfsMFh+9s1lmjpjiVyKimciG4uZjyBkn3ACE/FTDM0B5aWjXIdK0o5
idI5vHrEvzsZ3ctoHt2dP24eqRQp8wzLyPvHuYRY4BJNaTguTaeNF7r0ojLKLWS8
CZF/VQpu1ObRHqjsCs8Z1s44/QqZMMlUIKY3PCWZrLR4q5yYrqDiHuDV7b+WBTn9
IPyqBWMjMhBWlkL5PcDIVFc87utapNCx5nfKTQ1ss80Mk8yQSrN5Zm8vtPVBokJN
K57O7uAl7dP3M9eKi5tuyObpa5ceAK70zE9zfLLSq7B+nDJ+0FzMhk7bK/fq0Ivx
sT/a25NCT5Nqk297FQmOFZARwdjWXeFMF817iUbwQD45/mA7Y4kfpgX8McPPrPqT
3YZcq0bCyh27RZ2qM9a1ksirf9xDmzXws01/jn8LbMNoVnt0mNeK/zhiOkhC2ZO1
6eJUzC0x5hFlwvpoCmezmqfGom6FkNrnKa0zZJRaz5hA0M200tGW/bRU1/YkgC3V
0pyrxzS3Ff5jbNz7ZvpoQqPDkxM7OG9FtGWNOXlh513ArDltHh0YVSSsdQtL9DRX
w4m+ct/bsjp3u+DaQbEPBVplsFT5F5KrdgeQt5odYW6QSo63T7zuIIGFk92Pf62V
3zQ/BC2uEIq7l7hoNnLKIb8MRroNoIdoycf7A3UczLDYd5C6ImOEpb9CgVMhI0rC
CI4cLls8H7cbBTeCVyatAxWH0QdRVcqWGWwIhXEa9pOHZV1UWNrH2bub8WnOc5/0
iZUkutckn/v8Ik3i7b8JuJs0Tan7Bh33Ma3ttTa/CTsZ3IHyEo62YTe/NFTlzANL
lrw3qbGLJJmLQQMPMYwp4++uQT4wYT3PBHm6VobiEymsPGJco0F5Kr9zZJsYoLMR
Ff0wRwEoyqwAb48/BXPluFjeskhWsTd3jDhEhV9Cq6oJD8eRKb13r6MRx/1WOOHV
sjCtWnbBNEKCOMqXsOP6/xslKSe3DxiqavaJK366SpRXI2bUbsuGkb+Njcz0DCQX
c3Uo87aN79mi4m3P/Op/mz80B6hiQ+Un1cq1tD1cwr6eFOSzbtH1fZNT/L/wDOVB
O/i/xTGcljwl4xDJPgnMgQi3FkrXG7aNpooeynMEdFW1ZKkemaR8rmafvEtEduM7
GsquXO+snuikD/0k+Ag4+Kq8eu0bLTM20M528Xy/shvR0Vl1VN8JvZlClB49uwo0
FpUiExisa+U2HZv8rphguAV2lpbFu3L9jgNCKSoyYYq9/dzs2189QN4/UQwgdzkf
yhagPP8X0Dlh7Ut17y1r6T21p6espR7B6sH6HoucMzJCTr1Om7f2m/NShR8ZygTZ
Y58vokvJVHBlGB/5+672dblWuMbyQTrTYprlKZM0fqABWbnWcGZrAd8B3EHCsTEt
UcNhuaafFZN8BtZNfee7MuyY72KmoGTNxezDsLUGmu+WmJF1mhdQwTK0HXEg4OdE
1vSfU0ymppe2yLT/c6glk0fanVJiU9BA3nzme01uHAtNLQshc8ZdcVXBB3JPoj38
KDTnm4dHpoW5P2HhnnT8hj1QKgNdyn9Wo0S1/rCMhplXIG0E+5IiCkm2HtCNA1hq
mZySE1ntQz9uDJycdrQb2PNwqEhsmzJiy0j30vuVX4GN6NIuXJyc2dgQRqUxegLZ
QxzMw297cmOFqzWo9+SfJzLOQT9yoDPKytuEprkMuhyE3jPZ/P4lOyDWUTgmQBX/
DCJ5ArLj16BStRsjuIHBHjmWuMyTUiIE1jo4lPQyc+jSEhLtIpjMjDxPEN6Q08uu
asIlloSeECl6Rv/hz/oH93hd0DOPzf1YM0jD9b36eVLk1KvySM5g3aSf/IuzDCxe
21VqrFX4ezUiLWWz92zRZQCz5/0hD0CbM6w/7SHIMy6CiLzXB9jDkXcXsHuUM8mH
E7F99idEC+7CbJKvq2x40zypbj8tVjUPesYPGgboUzXo6uF57lL2Pp/1JC1oeL/N
U8+PyPBPrT+d/Kcw/VRUYiFr66VeFwIOMHmJ4S2MxZzVGYw0AxFKRGvqmMeBpUQi
WocHaXQ2znDMmbZ0OHGgH2oZeYO0iL3jIirZpT/pFO6PeBDmyzNdCv03bmMzNiA6
PnHp+CGhHpbJee41ReGEe5EZVNy1WskUKUX2TCCw1bIYyDWmvA7vN8UeHj3BFROr
mgsArc9Rw7+Fk9gml+WMBYGwOlm/HnbGCHoN2dUT/VCkL5Tu/NYNslrhs2WzRyER
qqu+5SiQ/PABvLtKXDXcxquRFLOgnbLEBvapbEeV8fRxbMeNYsxmSBKrWSZ8Q796
A1iVuR3xY1xMIuLDTZDSXz32+5/B0zdQOWOseoj6dFo62YMm8LEMmF4+zgyyTkTf
AA8L+4EBr5wktzzt7T38VPfK5qzrNlRmlj8u/+WH7/zWLyvTzDlD2nfk/3D2qCSe
xG0GOd+qzONy9/KELVKjZUaXEwScQjJAe3p0xZlSJK578j6LI1dSbyOSPS+vs3Y0
3XC6dZKRsMRx8AT5BOfjd+nyVlCSevbh/ObYxStOtg9RU+XjyTBwSWLnaIieA3UW
izHhcaam2+mXazV95O8x885PGUwr/rfmKLiL0LNBhEB50ba3+xL8EUhbLuArrm6L
i9eWQW1kdGQ9ztCerWfJsR6BbIlXiKPIfFvnSAjNnlwytxwKp46Qa3F2YVM4oQjr
ukAz5A7iJ5+vlCEb9B9RhxBVxBpW3YjGtEOAXVkqSIdBa7EsarJdX2yBHdiUtnAl
EtuZ2T66+M651uKVDOOjXm7LUW5suL5VNnO1FUY9oGCpW01J6TuLnKu0XAIHCqtv
mt5G7sKesKj3grLrq6FDJDBSebhlWFQMFwsy96pyOyqAElCp0r0cCsxVTkIvyXfx
YuACT5FbWfrLUd8AfzoSax1NB1DTy5/OX6EiJsMZsO96cLYZiKqGnKDsk+Q3TQEg
MxPH4EpkwRte0Ga53Fe28HdAhExRuV66e6x2LpnD96pqR2M3C8ieM3+NjFkx4lUZ
zzRC3BoP3XdQLL0Nt6kxlLpwrguvttxcG+VIsdwDJThhFHL01AsUTMiT1hSaB+mT
huB3FgsN1CC0rUS5/nZO/t7UVD4sxu+WkGwY2ZQj/BxkXFWQktQnHQCQzcOgNHz1
9gzk1jQobJx41Tt25Gswq1XGoGs6FjwwXV38M2DzzcZ3oFjzUBM1vbUDMVKwrX7c
wSDJ6S+HlgZ1EEteAnYdzuDNV6FEZLbbBIzRGOc6E9EZ1CWfv6X7uf992fLxekCF
Nvee4DFoFMOi9zSOYY8S1lnLjZ92CHHtupN5OoFKr4pB56ZbDoul/V1Q+Ubdx8Zn
N5OYvX/GZEI3wcXKo4c2rNFJG1+H1laU58FPgCFl9dypvwKSH/LLu4slxkxvnyqJ
0lXDdkcGSbWvvVR7pzj+CJse3suoRPmzOo9JO+dX7rhYAbB5NGFi3LmOPL5clUSs
K3fQSj7GBmcqnMZdzAi29W1yM9j4JciqZNytIlyf3bMPcXJorQ3uelk+9v1UKCMA
y1E99qUnjVg5qazkhQZTmS2OzcyPHUnGSgr0fQLfogiA9aglQ6X1MbPKZyxhvSsw
R5kHXYBfILMlSq7K8qv+jSHEtkCw1eKoyl0hPDo3q3ra4hHIpCxWWTLwsrd/LU9t
xNVx7j7jbYoN22JXJvFQ6EB2TYsZEMp9V2zrwe7UlsrkUGweKmh6Svon82iTQPZC
AAJJEzufS8jQhN3Bsdkka/BywVoRQov/kOephDPftfU8zaRJBxMi1JmC2zU9kZK3
UkUrjSwrCuhy7z9Ot3ZQjiIl8CuDte2Zut/HxUdTHwMBTmi3a4OgOW5Hf8bGqLer
CXdl9sivpkAGi7HfWj6DI9Xhn8PHM8m5Af6rUc1WQwtkw/KLH+DeJUB8mxpCyI1D
7bOAb09JNG6W/xLGxRJewSleGfzXd9bimLs3F5yuY/LVf+bOTdzFom9uBbYzTF1n
BWvxgkC5xegcc7G7jwk7TkKt5B/JUrt9epXOnOtpbPfne2UzjesF7uyBNG+1Z9po
WuKhLznlV1wdULkcEyeCqAJarAo/rDw4Vc1suSOB78jPErQW4x+W/jv+XcsoAxbi
+4OsIT4vHOuBi3oayeFDB9sTyf0n4f9pa1x0Jp5geG/VPDyif9zziN/kNhLFAmX1
OlmMhzSjVpTdMOW/5L+1C5XgcRqm//ghNhBSgrM3Q5+1sXFeCZr4Et41aa4DEbgN
NXGDSoWpyKLsPMU9bB7uhtSGD03giFJ/CC727RoTUcDeVU7mhDq4WzZuXElH8nbA
TRi+fENgARQUOpOMsytgjnaoepEl+ViXyZLhBPLHhxtjvDBvW288dm328JBhucS/
xDgdLqPRQKzY77mle3qJDJb+Ny8C4/atxcL9uOlbKHVzkMZ2BJu5/JkEQyek8YQl
/yX70lpnVo3mKKLWnN9zWY6LZAsTA3+aVo7SYFJ9xwrBw6zMz8/CseSrrF4xWBrL
SiXKr2bYL4tkvV+MS9BJAk9AqMqkQt8PgG7Kr6JaofASen3kSSUN1GGAafMNBcZZ
MWN1/82mzmLIEwjFRTImpo/8laAYI6BS0fPFBOTmB9PyXRZYlvgQKY6frlcKpa1C
TFfLvwxSGnxF3TFDfWIZjSGA/ZJAyXYG5TlkjXfUSbCt4mMDVCnkP14VqUXEOhIH
HvX2KYrKLBEUZhxaNPGvEfQqIt4mBA0AGNKUO+d506Gznz0irSxv1PbmrpEPbnay
Q9XGP4gPtsgDcmgqJbSPluQQGt3/80epwgMZVupb0OiZON1VvDOT6TL9pAujdYpS
4nRv3tg1lJyufUv9VaBdJBYsDfvnbtcUxG0A1NxUCYkf9KrRzCQDhqYNqHRUdPZh
ivyvnXlsnj87QUqGI7H8zo4VueffY5c17FoGOnJ/3pABPyTwtp2I0YMB3AdozDdV
iXcqm7/LGLRjhwEcRXqGSLvx4a9cOUYOvcLyvEYo5Og8QZ/DkSUPtCsqn6+Hj8ns
MusIC4ABb/j+kV+13YOOhJKySSuKXto7VEo8g1OWPzdqfo4gsBBY9g7bF6b16KUO
2BZnTpUd0gWlgsfbuBtiA3CpVnm3heB3f/J5kwhY+d9MEQob17Cxy5k8oZyPhWr0
meOfY9sEc4556JFooc6uxQG68P4DQde3oA4CONCe634NDM8KGIEEDPhkSQOUqd3q
Z9U0DjX+UqJc4emBoZnYKRXjKSry9xv6SwLRDMmVQqMfJEIpDk48iqd3SmOsDeP5
d/5gr6UrmUB/11tFtUoT8LUtPtiNWJugPQbsJd2pxLu2D871D4qWZNzg4BVAXbrM
INhU1V8uGi5/ktMCoW6vNYxwKpSVTO+qaQA5uF+nucd47ehmiOcT2hIYadLtJZMj
vkMRglNUe8/32fl/KvUN3rxewOBc802+M6LCy0xNIK7mgfrmC3O6m5yMRKnjYyyp
DTB+ES0mGxJbyCLSsfSDvHYvLiwAJu7F3/PgSQJCRrrWNiyo2xOXRLVZ2usv2uYa
OE9ZpidcpZEHRZ+o9Mm2EvGHLripMG73+Wq4T2+1MT5nO3sZQjyxwYq1sfcSP00Q
loZ2jLJE3Lyq/Zip82PxJNtd/8H+LaXYPA7+N0QBwCtSfaF5KwsHNLLAGJtSTcHN
wt1YhqNfEBERmIQ59cjc0U/wiwKV77HdTR9PzNRBu6B3DBwsLYR6kztukIYah3bO
HUqinVIjvjic/a4aStSEZDwPGdr0xGwakiVLgzpvHp9a3CLGEMfKjmJKvMGv1Xh7
EypwjsCTINQNxh3vtCnviWAKGMuexkYK4B1NG5HpLPQqRSu2O6FFHAtHCsPbL2CZ
pjz96+UMWd75AJfxjmNwmHWOg+XdVKCuw+UjcUI8OYaqIArPtBnW6AHidfjJ3phY
JrV2UxwyWF6zH8KOYFC8R0PIL206TO/elsxJc65yahcYtWyXZUkVzIa2PjcE1yKi
Ivp1b5z17iOa0F0oUD9uePJDYXxJGznV+oexQu+4s5ZbPRUenBiX+lG55ueg6pbD
NorXKUxuTYjDGBM3klDP/QbV/8pfzCWyKRZHWqlmpgHU14NgmGXnlD/KAbj5KHhP
o5vl/bBdTyzG70mX2iA4sSzg8pQ01rIRKB+zVnafU2MW6YVeuutrhJ4qGoLHe9C8
onelHYpLlnxwPOqsXh0ayqYqBIoc7W+TNqLMyFJ75Qo7pnqyHmzJ2OFKetg27DAw
+ByDiGa4HsOGixJ709ktTFAU+0a/YBOKDBdMOowTXEf7amzrU0mBTEAgiQ8dkO8c
xUmohcLPnZVDh/6NEbtcT0X4cI0sfLturlGbuOy1eowCT3CDAlkCQoqxtHR433AA
zc4bx1d+18cVFI/e/36vmbTEjl6wp+ZP7i74cZse8ri987jTz7JdpS7f8J8PGIkn
5PnrLV+xewzly1Dreg7d4csR+eB5yj6O6ECycAm7XsL1n5Iv5CRMWS7qpNP1J7Z+
tyIMWy/7xl7BWY6LU0rhPjiB+Ue9PnYPDF3+GyhlqDpp9APHqaFnOrMg+0ime0Jv
1UvY+d9dlBMNfLT+JWs0oaXJ3hGEnR6eySciRVz5JwJkDvkE3Mv17MEta7dQZHtG
bO4o7YtUvM+QBWJDmfQi3qqr49iIX39BM0uzoceSdFECawuz1G9bcQPd8Q+DIsWb
hbsSlyeoFE4YwQr7dl9EWt5KbokRI0vPZpY8XcCXvSsoMKfa0bT3h8ve+mD6FT70
sZg7b7mNFHl6Zhsgu99Z6ea2fqbGyYBgUseo4zLkDSgNGWBddqzUIicV5l50GIok
mkUGuZTGXWtd+bwNvrYDCmpuHXC+KE2IEa6HhfJxBveNwe5WYgmefb8LoiDVHVd/
Wu7NHbp3JsgINl4EvgVh4OIl9K3lW3jV5BkXwVWKkyIxznsgkWbBiKkhxFeoKm31
Skj3Rwf+hvMezmUKP0968WyLd9/5Tpryh7T6gW68SgdicHg3NMkrFc7Ie0d1lASF
V4KgpYyTBklVVjGuj1n96Yxv0ZdDPxYxOAWgC5Rhge4oMoe1W/aM6scl6vE/laOw
V9bjBljYYLPinX7eFw/WHDbpsfBqzHyNUvTtaEYbbrkVfKm0DbvyjJmnlFYl8jOP
Fk7M16eCK/MgTNsiL49mjm+nazM2Y9yxYHBVoulUqNmFHtkcrlgj8sNuQpoyxqUn
b4C3sCFzekgaop3RJquK+iu6jO2xJfWZHpEVKB+zBy7N50A29Eem7x0Y+uVh07XG
obhBDOo9KdJ+mjsaeCTrBnVCgW3iWc16iYgT2HhOHyV05NOHZH8vvZnB2SyNcXEo
GkE4moFRtcF2MYriJvitmKRQhrDJ5VWIM8xhyBjOZl1UZP70pYsu9B4i67xpr3Cy
uSNEispsSou3FpTu4qGNMf3OLtUY6B4Z13W7k5BL1jZrXB1JMoQRgVxlniGOODnC
E1NOmqDOQ1bN8YWxouNqF4HDl1lTbOtpa1dthRT0hodqZsDRspNDgBxiv9mE3OpU
lgyFjch0XfoO5Wpgh7Stahf5Y7x4SRTVv9B2dflP8ZyCEULx02Wf5RjNqDmnQA8c
kIN8k5XG9KAnZPwy0p+oL4Rl6CL97GNjDDgKQEW1rAn5aLi9P9hPO/66LuSXoiNl
FL2e/lpfSd7hG2UCUXqdlNExXTvT8iHSKWVGO4tV4XTrxi54CzkfeYr0aUb8TNy9
nZdpfGR6utX9VGXLthdsxjdBozY/SKALpIAeLt4pjqw2y6e2FA3ZELBa7JpOksIL
6z9zshAscfbc5muRqcKzg+OYuExiwlzk5eLM5aDNliXD1SU2cwYg+BUKEpNUgBt/
oYI2VxiHzAEBNPgnJeslABZ9P2jrBqtZs/OLF57fAevswF7QjGJcf2UspCFDLL9u
cQ19bVBGJdxcbXDSVEROpc32EuMs90FH6oqjKYFzq5XhVeh0x0rTqcI8oZilVvgs
o3GksFVxksqv8cjMJoJ6TawmP3G44f5yc4YKN8bs8d6zt8yTnhSB/nPDOoxfWoa7
gAhtkk2+34dCwfUB+HNUNeSND8eZKvYnXJXUksKoiHrnfxACusc7xVHH2ZePql48
mjzQ45Ot5apwnxnqtw74rMmmGfULHLns6aT6ID2rrBXfeF2NOME/2zNqzac6RdCr
w/C7BD+33bvVqU/sWmiNfg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
l0AhF0CoFkt89t77x0PQrjBm9WAqv3e5SVhJK2ZkM09QtzvQuJt3FQeiIxfrBgzy
BrEpjn8PgOygwQeDEu013wPpf2JbpV0TwN1QJ5rCDf56Ug7WqNX0LFCd3VS5fZ11
2j7K8cHAzNcSDVqJNEN4fnXeGwnnfRDVDHu+oM0QO45EzWkZJK6vuChkir4HN3AC
tfZU/JGODniagTEQY5/y4mnfq5JQJuhAi3v7hoddHqKgjdo2h6eeJ++4bR425s9e
3e4mU+9lC3etKMbwNcmG9IjtiLkEe6G/StWbWG9nMW1H+CbrfhsCt4ziph6vMI82
6H/BOlT7ae2CCqT7cgUIVw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2864 )
`pragma protect data_block
FmCPeudzjl8rgKddnCwKIdnsSUUX/ZUuOdQyYxnhPDZWfH50Ju35YP7rdrlXyybR
9mqJU2900wqjLWo3mgHMRndJNJNRNN7cVIYgD2LP0P7zDPPy3BJINErm8Z3nUx6e
ynNBS/aPYyTK3+S2K92TwpldrmISO/gdiIpdBKbUUUxgVdzyv7IQ0KMzjdtv67DD
zwAoLZv2tem6DkDfGzPL2WHOmfToNrmCvGn7MNdjWrZAeHaMF+TGS+OE9EOxpCrg
b4Bm18sFuf8elWQwHoxSGPCJ1iC8HUkzB8tC1WOof8DVKaj4pmKzSStt72id+sld
4ITPpsyk8Ekfz3r4uZn9vLc8VNFZlORANmt4KgD084ApixMnrPZKR24HhDYXnm53
0K71/H0Wuj2abqFEywoHFEHM+jeJGrogH1EYhpcZbIRARUKx9S+4QQ8D4C5GCuGX
na8Y2Ta+1cohYhRyLXRNtcoViexhUN4zP9YgIpIEUVDDvXNose+0TNGsPVf9jeRP
My/8xQnK45fUzqkQdYwKuvmlxs9Ck8C5TJRGG0qabSIfln1IM+e9eG9U2q9kgny3
qOHOTZmoMgzIrOI3ab68tRChwXaClzeqzKYUOPGeISj7WbDQnGm6z8ipss/F+gHK
bFs70OLM7qvz0TNSHkIJyDi3K1f7h803Oa7nuCAJVfx0wfmkpdHXm0tFelyRRW+g
4kF8cUEtOs+CrYl919qz1mhu/70YJOztZbHJUF/awzogrwWB5PbiX/2/Mbp0s2vl
SCLBM9Og7ciK+G+4zDuMXNXObwrzcmsuCzOR/QkuN09xd4+5fjQlcBqxI9McA9xT
2j0ptgFjAOZ6SxmA1VsFVrkFhxlJTGR2sMH+8Qb1JiJcASa0dw1eavikKIXnDHTG
NOkd/8EQ1mHas4naNysKivT4Fof/edX3UGVNirP0NI7ursxOe4tw9uFtDH2NaWL4
/uzUKHnRUj+stD5jvB2PwitbwgVflFZhr/a6Ixc10J0GACZiTjLE1j5nkDS46uLi
QLsZiuoXjWQ63wPC9OUdbOroRR7SfvAIvqZnPeAYlTJTLFdvBzTJAUJt7DwDElFR
LGaHrmzsgn0jnkPfRZToX7qIGMXc94IqHnuRdRkquhBniweMfujfMWD0K5PsY7h4
cEQtmthHDRpUmMo1R8dnBtb1IWKbt6qZZWbyjOUK4k7qhhLo2SxkVoNvRDpZr/51
ERY3x/HDok4GZmD5xjcy0cF264u9sqn7QZ0gkm8FeSJxn63NL0R6iZvoXJ7edf/7
FjcT/COU9w2ewYksTR6XvGmo6Jkv1+HyDl1FqRoqJGuL5YZr24JzkwhjoA1gUkoM
5XoqgHPMG6kIHll4lKEcCsjH9//IJMHCFJUAsmbdZUrHlSQqjDl4s/7K2MX2nfu7
j2mvVJ52sA62e4yxkj1LnNamcA6UdQ9b0eeakk9q3v5F3z5FbHsPnmGLXBeyJK9V
JRnRjUKcq7hZh9nQQCPTJyMWGBSoNWM3+z9BcqSSLMy/bfpJkeL04gE91yEJEvJu
gZxH9SVq6uAhVSH3ni4D17WOU4QiGVG2Ak8AB8kGfQwKTOo0JLGxtrTAksAMNYIT
DpB3F58H5vgUVdfXLexrn0KLUVHF6AyhF158G48yRkkjttxuu9sFnfF2XEvTSkEo
JchVns91/LjrCX7bqPilbh2dbMtbq0WBzUgVbG6TnUTO43hrOBg6R7LP2j4EvYGp
BcyJfVoPpULLMsE3Rcr9+XdKPpoViTA2B+MI7JSuFn2X4h4pJCLbuXkiON+yUKjU
mhlvZ1rL5AXshEEfibER2KJuotivhkxmTgaseAur2633YVah0si5fbXDS0bP1RwP
k68mEZT9MZdRlBTznSE5/4WeiXFLYF4R47rXk7l4qtbizm6LPYx41S+V+O6zTEwn
SnGncXxSAVqZrSJn9APZmxDXfrSwIK6ajft9Y3zLrGN77PL1NvHjHatQyzObH3Kz
YlBwUFIZEpK0gEMxmE3H11FOd0JphOd05rJ+PCzWuSqKofNYPIggpbpdVW6HTiwm
8GQaO3cvnyTD4y0UVb6r7TrXXwqWa7yqdC/LqhSlq92ZJQI9aFWX8D97u9+c/tdN
ybk4sq3pf6ry9tEcKKsOwr3slZzv/G1DEyDnZsBxvvJYpDDpVNc99CbfxVlc/70J
CaHE6cORF3Sj7w6/oZnyK0AvTBCqE4ni7q13Uz3st++vngCjyw3VRR+Pb8vlU/bD
1j7tJIWzTAz4jZhsm7mVwvzp3a+lyTzbdSPXkiEaX8oBAfKK6smtc4Vze4DOI8/e
FurZONyMJf3NsU7ht76CoE0MOxd4/J07s08B41UTD2zjb+FtubNrIf7N+slH2cxh
RG7x2T/j65U9YhAZz7GboAobMKz8V4X9wDZ8i7znlm3F69R7RoYIcEXoxHT9+Bzg
d0jwvaoCJ5X/KB0aHEu60QPmnv8sJ1XsbiiaG+S4503WdPc80S+7/Qzg9Bgj4Q18
V4K00o7c/NuhMD4t9PeBuW0CvbGsLoV9ygKJei17xxv3CTgN7hzzcqh+rJsaI+A0
QE4c/mOXU4E1VDLmdIpUdBwtn7WQu4x19Wfo3I3303nbWEQ8VoR6OrcjIYCKYRIU
dq/F0GV98FgVlIeb3GgvHT6xUKBeToiv5D6dCzwoJ72n1nAVnbEquI48cFJPD4dZ
Dw/XKhGd9RDZyWvvhALg0ahOSQE9dVM4U6T5jagBNGj743QVqihs3+1V14iUOng0
Iz83UchehZzVImHf7KCdop7ZJjprAb236mUgCylO8XP9y8/m8fdgqrHvBXkg7qRA
BfZxdiWwKzor2B5s1fvBV8yD+5wMX3I4qQwqNW0wjg7rZ0dmt0/4ttvivHmCazWN
VlGw2ut2BB7BFBKQumn8/KTixbaQs5XBhwoRqjRAQwoLl+2fpVXwX/sLAaGenbqn
iD5eVMvwSpYUcRr5iM+BBmQmThSc6LgosGTCBVnNkbIQfl8Wu/tthFAdfYQzIPi+
GkfJg1I9jC1JHVHSHnzrZuEw686D5UjTKUcdGVGwx8Zwg/xdGwWltw7cNoP3d2I7
GnSWuxY3ZkKDxmE3rdnxnzeTtSKzXMaAYxkSYQmFFjiCxREb/2iTNjX8iNYAypa5
rxZSqeFjIKWTvf97XoQwu38a6p0UFe0rKWEwCoHerfBTk/JCCXm/CJqA5m4VSF8I
FIVtXpjtL2spkviqiwxqgDdI6wnlSTYE2eQ7pOuvMIsIxwXFExQy23Pq5f9tq/dN
e/sqDv7pJI03ffsCrFw0Wpg3ncANrso0OQ3I0RLQCzGfFNeFhDLty8kUvVaZjhed
0lGkI+8Vpasf58mf4kJ1it4FHJyjjD81iYFF0/qH3+NBfwabQ21Fmc2EIB/f5mEA
4XMX9gi7JKbLyVB5LUWwdXJTrI85SH9dfKExVzmGzdcgdXXD/6S1dMtLnR4KJWN+
8r2XDTgIp1kg3lIQGjb5gh37HBvQaRIJYTeiUGw5XdrmNKzH4Iw8rbBnnSZOzcNu
+LF1asQNkbMAZUy2qnb33zhmEM26018+S0xoQdZTZot9hfaaCBCHDxfDjR/3YPRq
npKHNfvogTnKw0x1KJKcXzCrVjUbp2N4YGgkr0Q8IoOy5mJ/a1kdrzbql+UtPfu8
BlWCQIN4Zzbr/U/h4qxzweIyCtq1/wPRieq1N14C3+pQyFL94+6NjFbIM6WMc3hP
WgKWay2m+pQpz2ys9oKT8+Cxxdt94CVAjxrceLdTyHR32C6nWXXZoysCUP4Ep7Ov
ysj0/jg8lyhM8qll/+S+PuL5kl+5nMa70CjC1uq21kE=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
XI/VsOoyZ65n+wtNS43n6+DnjbUzqXGm0YzzBQqn779jr7161dwKA8kJPWZ/ER0X
Ez21s/vRF0cr+EHVUWuR4+qlU6KSNp1SNOEOJG101tJCEG81Y7GXwW3/hvRU9Y0R
mjzlY3HPpQxCOxFdj5A2UJr2Av6ajXBJAj0K//6BiU6SjRuHElb/waR2SQeujyen
neD1fi7VAzdsV8YiR6+Jz03BIx38+1FSc9ub61/9pnU5Tly2WXLQdSMdB+bWcNt0
B6UkRC5OSh/uHpPGEpvuw3ScXiK9ehoTVKXP6m//uw0CZAHCwCIZua7IupvUTVit
E/ff/D4W5Q/t5cNO+V8fDQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8704 )
`pragma protect data_block
DWgfNb/GqaYZlIDvw+4pi1mHzaUpdZ0kv5c3uzObJBwwZcVt3nMfCZWWUAc7jvzE
s3DNVKoIdi6Dpmg/fkpph9EwIvmwL8/XEozJJwMGHDLU5yHZaiq28ISDcwzDRa/W
RJy+DAamX+3Xo6UT4LbQx62KoYOmceCJszEb3sRN/NpIcWYjxWQQou++K5QAKiiY
Mz1RW4eHKz7rlgS/LUdMtqLdbiSUhuKVeoeWVi3uRYJNQzDdxmslGP1fbOmdWZPt
SpzoGHdEhYLd0TgkmZ+ctA+GaJKPRkQHgdcLVf+3QK39NDtjWuFUzyw4en6tLuth
RgBxbRsECXQgpmV+ToThl0GhAMMqtlHSRyZUf9S0HzUcJHjhEu1P1I29VEIMBVKt
SUX/eOj7H9jemC13hWyEcuA85aAFti7VWhAAH7J4r78elHlIr7hxKNzhyvUMp/7L
SAvyBuCklKNPyhO8ALaFxu9H2dzirgfpHdaoBR4yjWhNiOfQ1tU9UsHG/PqV7R9s
3D04x+a/91zF5OmPzRC/WVsiMWHKgrzdvvJ/WFata2JNxBCPSlNdKkg0yd469vU4
VWCirD9zG7nj9BlP41S/58gCpzASL4pBaeme+V0HAH4DtlIlxl0oLCAkXSY3k2e1
F4J1RTcrJx3lvovLUN51xYGmrFAe+PLWHvgnw/Nc+s08NCCjolaXmarmm6WoMIq3
caLcK3fGQXgKhlB4HvxYZZ1wq//Iaj5EwULeorRMylru7WVPkWPenmXp+R1y98w2
f+5aGHZ2khj/X8SLSMoMAgSz2eozEkk3dtQyXKpT8kUZopkUrY7YbE013u18EHh2
DWgmCaC6CghKdjwRIY7GXuGvqTIvb5L5n5UaaaAQnpAeoLu+fUZqxaFVacg/usrE
E3Wlz8DF5AtrzrxPOY6SsJ1I9O3XTe89R13mLEX2/NUJE/0LbFi0WOqnjEO/ocbX
oT5zUoyEaDhhj/JWEeVJWoztDvAtl5c65btjwxUl46OxlG4aE2MPr9pOvY9Yv9X3
FDrW4aOkIoJXzZORg0e+tX5UTnm55u2AHLmmc5cx7a+yjbtK3g6tmQLlxMgyOV9z
cGfHjsnPGKajHolA0gGOoU8FPxb3cpBJa1ScT4YuA7Gi420C61JAXWebsALJYwlJ
ZvQcbQPDVeRfQqCGY3C8OVT213FD6JmNRPiEL9fBamrTXXb8JtoXU8FqhyOeKscq
fK6lNV3oP/J6f2TROGNbkWWj2woZcyw/2JEvnpQn5ozxKsv+al6fLNfZjS7t3ZdM
VxeuSJ5wMEG+pXn+rX+jjlwXZVzfYaeT2D8TsooU2tjR6Jdri+onyStJoriMC3UF
wAL9tR9uX3mKLQFf41kyMDJu3zf5+WzaG2EwxCdQkXgt7wopIsyZyJ+eHzq+Rj+O
kZtna8P+YCvZbsCpkZBKyaDlHQjIASW026K5RFPH0oSW8c0ICF3mokflZvLh737z
NsatRYIBj/+nK4WZoGA75PmUtAGUeo2+7zJINviUlptdjwPDCJ0p6FwpmNeoG2s3
mVNTf/bUr3IHBkr/fhXBKOCi/Ho3b/mHin2DqN13wREnN2bxdfcZrGo7x3A4KAsa
zMwX6iqpZDXixG12CN08aQy1LQtjKTgvb7VL/93XnxNjdramBHBRN4b1b8hEO2ip
avSl7vsvxxyUMyCfAcbt7+zXem9NbDlyUhFDC/s8gJc72nc8GgUAiheKLINxlxlA
p/4ygzOBbhEJEI2LUmmNfS0CHsympRLGbaoM3gSq8Sdn/hYQ5s6Y5C5D1kRh8Mui
fNG3BeYYqwrvb04F4+MoM/P1CFkUkguS2+57UjUMcPsDz232MBB2IkuNzTgNHqmv
pJTetBgydvy7enD6hHlXO2yCRP8LjRbtrtSMhFD7VfpF61+fZFrsWXSrArz5S+Ty
bbIxBCb/1WX68THL41JBV4TrvPLdDlaBYTxzCxb95BX94KGiiWnZGdFKqsEVrL+L
RRHI/yS8UvjcQwdjYvwU+YDpOb/bRBE/JKOu4Iz5pno5Fm2u7518/Tg85cFcACNl
PA1AbMamXhXcZyGbt7fg55TFYClFya/1etFngTfEl45y5dQs/0S4/5lutUdUYG4a
/4p/vXdMJEve5LLxa9SGJMMEYIAwjrLLqACUwYlUCh8vt0rcmX1kDYGQdX7odLa0
8WtsGFfcpz1fTeX8UWbQJAvnMBMKWxVV1OfB+XSzkwFkk6vAAi6Fd46/NJxrukcp
7RJSoJl7Trmt9X2fsw9nxjfXzCjokS3+TgfTxvSARSd6x91zZ3oi4Zjhddd3WRDh
ujEyZshE2TjWI4fR6bFkZ3hVhawcjYsbhGxdvEhfsAXYbIPrkFoPPL2WkGC3JNmY
7xaGD13MzFm0dihYaq8Q9MqoQ8X7J9A0IlowC34SmZnryPoRsWwt3zroiAYZU4fm
Xepc6cTA9sVu1maUT1AMdk9oNcefvpLutry2P+X2HItQlpDznIIXWzqqwOz+XPoZ
+7bsoZZzvGRun3fyaXUUhoOuFvVIflzLijJkOvxQMIu/WqVlWyg8v+4LIVDeRSp7
tYOroawCxVhPMLwMfoCy4LZ1rd6NlDZ5PIkftjCx6m70Iw4P/s5Tw5nwIOyTsTjJ
XwuWAnZu4ABA6WTEs3r/MH8UGFuFfo06uSYw1G63RcEeLtM3V3gIbk+ODqV7VraS
nA0DOqZqUVLOQ2k647bbZvVDUEAwKANOFEQ7sQ4zrXXFveKr0uNQO+Zll4gOLVk+
rmBqxUbQIoynWstohAHQAx48nrgVSqAHe/vMjAbwk2jpOy2n5IW0ZmmYSMHp+nQJ
fEQEDda4kuLMUuwaYRwAQKKLOM5qDoxXplqnCiAHVdjKUUeLBxcX3SyOYff1kXQ0
wvh9NwT+MHWQ+UyyitDjERKGd5eryeWS6R56Myqw/0f9BC8Tb2qjNylqS5AZQ+k4
yiX1bWGYV+Ec9peNEeEMTjQ5K+kZYRQW/KWCLmfbBBhnxITU+T+5JBf0d9zn6sDs
/WRePdHDfXASajSw7YRYIUzEePLVLhx1/KRe/RjFr813eTX9ARQhxzcSyF5+o9Pl
LDZkQOCfN4nUVsN8ufg0szpXZQakelnWBYD9IBiG/45fmv6f+rzumKRZjayOzVzx
/3wbCVvPyPJwmzrQLXdyT1qvNwdBZuPt7dfqS1nWzNr/9YkHM4dbY//F/ky9ivTr
o2NcVaoTde2zk0LEHOZkOTL5IxdHPF6i5+hdEqf3m9uYMdoGkz48y8MAAwlg5pwR
+qQna2hyEkNAPft34w9CM3KU+pjC98lEt4sz2g/QGVvaiSO2i0gK5c8nB8zw52n/
jPiQkaUOiu3/J/+aG24SlNiHJnoowqlw2G6btq7ssOr/lNn3tthUgruG5FRU5QOq
wdbLI3n9pLSmVHJHcGC3ZUqOb9CKsGiYa0VdTbWPmbfFZdxP6mJk5PIYek/b6Uty
96uMCaQn7H2hQcUjdohhzSbGad8DeFuOdrBcR/o7Tt6yO28XjkLLgR4v/d0G8pjm
vWBQg1WfNNtIj9qhwiLqy01ftaS0Q54WbrKO9dvfcBvsSQDsmFmOWpRT9nmgWCNy
gGLv3ErUZ41ZHzyLqFmDeEFa/3sJR7DPO9qjbhYefN0qHDcK2vgc/N+gOSmCtyY3
jfMCf5fUZEmmOQmV95S9zWpp+1MVFBPA2agf2QYt4tLjSVqMscAaEsBowRDJNwOD
dVovnK6NStkXYS3vRLa6vQK0AAGdFohihBXn3qVgNKu9MCdYgeCYepq2tchZp2nh
wQRz1XY+AD7DuTCrMDCDHvU7yYzfhbgaS+GmVbEQiwxiuQskT78/bCP4GzfoiZ+4
4HKI35vnxMf8DVNbGhL/VlwNCOIfXkTTBadxsFzvEKy/F0H2SuOh8d01p7YceKuZ
ow4K/A5ypinpqMOUMuK/k0Ft1xKGygdl7axzT6WxpQB8Ks5fyRUnlGAdNFQg5D+p
85wG/CZy/KMvMHl5WL6SpAGF7Jw5VmsizXdtwqxyUKG/dcRLpBmy3WJWCegMIDY3
zK0Wfnw5Y/UhWyMBixb0ya8D/C13DWpZ8/SKTrLf6NbTUc25tn2QcBG0nHbBn6v7
w2sIbtOaTjh4IvmG9soXmhB5CZVO5/KSeWUzFFpolWVAgFyQguRtKQuTfQ9L1Zkd
ApNAfJWLz7bkCJbcr3wwnxgkWvGa9rZn2vFosysjahWZMYMC1XUreOvS3K/m5G28
77Xj1AB7H1q6TVsf729pfN5+J0GO4BCkBY6KX/VNbMf9wsZtjjV6wtqDOsiY4IA8
VVKd2eVg0evNGQbn4hJ7gR8j6nCaFqnRRquwO15Pp6gMYvnBWuPscyWRts/QXLB8
dgLO7/a/7nnmZRcRLLJdCN5dMTyDZJv7HdV/lz+2c5KA9OtlhnPAWwyu+DMYM3/J
d+jLW4uwTBeHVTNUOfgYNKkSXt0hC1U6pps+PwwAj/kJDTB+dM1tnGhR8wtAeO+6
JKZIbxLIuFCtmumy9EQhx8oqX3quCw2mDBqA2W7CtKIEO5L8HBX2FeBjRkRCG1qV
KODWxHDJfvQthTE884AYXmc0ni2Ibw7Z6RUhb8S/UOi+x5i1N8we6JU+BKxCoNgV
WjkyMmmSYQkHrCOrSruMTW+NrYOXRaW+Ki0evo0FTShT60QXHoxVDCUNTp7K7Xvm
tXVvNfqkv/sfH8JFYjP4n95XzcgrczHHNBGZGWibyzNwa06sfFDsOzk0MSYwOjIg
guqyKJodVzvVwv0ie9z2l7YwCyenotkl6/2HZR6LI3CI/C89u8aZgLQmvpMlwE5o
VGI/8yFtoMadpssi7VZAj7mcpOIEI368bduDMPPhmLkQUIBjtDBj8ZBhrtpdLo2J
Lk/U+7UQmyrTHbsxBuOEDsEB91SHUsqyzit+z82L4kv+YSqlvfamt1r+Z8fBsNqB
A83gJI0WWDjLdJsvbbjoMk15/7PEDM/EElRTKxug+P2R1p+yK1AerqofEp6Vmxen
Hw2PUPszyRx1hPh6Vtu9pSUXkw9MtFVLFO6eNW0/yEfNzoBETl8dVWbb8YWy11sW
dw1pOS7oTuydd4mcb1dhgEQ2io+eaThdlpbnkXjPW/2ZooVX+VuMVkYbq5fkz0mh
zbE5Ot4VdXEZwaB7vnZ1MOHH7fCFnxgxIWS/pyJf8JBW0yPcLUFHUog8iBnZ3GhK
1gQaRJcec3OpORdG0Q6s4janX3qxdlne4RI+LGWyQLt7flHNJwSOf+GAk/fNPBzE
RrePSlx3Z1hBeZ7DV7xDVyaiGs7lvCcZMWX+Si2XJtm08/ZOA6E5gZKKMmL7Pob9
2YOQqx82eDy/F80Wx0XFeUC94pTDjgRP7LG8qA+JyYmkh7Khs86fuCCwq4P3GM3O
D0u9MON/zdwW0xZ1m0caiLyIIAkg76cb0JHy6LEh6Y3dCRpcyW9izZ9tKcC7ENGp
eIauL2SETyEIuV4mpZXe4bfL/+9F1id7cWTv8m7eEQthXMQhT3BjseWJTc3vBFoO
GAT/r+I4MAmkTfL4QJhpyqfqRiqdsEfUzxsnkznhbx5UsNx0bqC05oRxMCVVFB+F
KevFqqEmQ0a1S4/g9YcQD0PcueUx+hq9zUnhne+fRIID3a1N9JzETEGCZZakWZoY
ZlOPcvtIRZOgmbw5oJxExg3DYQtWDvbgKLJG7y1W86Kk8ePgBYVXPL48sG3H4FCc
IptXQ1YVgGGvup3JerjRLwf6b4Cl1Xortf+qs8lCPy8Inz5D//o/NIiy+BwGM7sm
3g9EMyTnsduPUuzLbDRODg7CHES+I2eWFWfMsJPJLpfxEFo0Rpq5yLt7u1YAd3xm
MWzkSghxcoVhhl82Wqh1svqiubw41TGIZi5HTu1/dxBJvQXg61s2qlIvPG01EPzQ
rNvxQMdtT9X+6RC9Hr60L/kBzZwd5WVpk9k9h47p1gvTca6i404NE56WEjpRBwrt
1e2tbIFtQApC/+OlwGAcfaNOduzaU1GUvrdnvY64bm9QmFLC5T7aD8HYSJBtU4pS
xz5lBzXHYE0boW3MQgAKVmW1ZQTRic36YWS5NG1vaZpyR6sjhYk9+qimMa5rOJVy
W8zwMp6wdM8o3XSPsLLCh6ThG0cntpIzAOEx/ad7GfL26aa1ysMnNF9u6ypN1tCB
BXteJ8jT9RJBc4+SJvcKoiuUt5WIs39T849F1XbI3rlruiKOgDX+688vIo6a8MzY
Co7tjxot9WtpknFps+UVVfvwdO5SBL0VA2cp3rB9UlfwEj5wjd5jQ4scInCNTUhq
nij5EKlogtETQJuMqnkKVg8fwUkrggPYtELrTBjrbsBbLWw5csCscW8V6KdcP3C0
Y5nYYjfGbGZ3pDTJO5TWP3KJ6rVaWfHBpoycXmYhc038zMdN9ja5Td20trzbZ5nK
AQwR3T7zDHNADdi4nzYodPjEWK4BTGZUj9VdSwnDpvWTDCApBR/RF/e7QnEYNIr+
sYWzFqzL7BwzE5qQYGjIvfEUj6NjrbUy1cJLgzTEUsrTm6vygK1wDud8nK7Gtrfr
4W6ckr+897qDWhWHZZRaxodGHjv0iraV8sHfkv8Ag2xvgqSyyT7aqNsRPx4AOPIW
J04yvMX0x2kVD0GYl2NlfLd/MNrN4RlOktj7pyAKGzEbRw9kpRFb5TCxd/cQszEc
doan/4DDEeMBNbqJILkAbaBA7z90647hsXYCVQeIdoYFgA+QLMpadCUlyxf38of5
3lnkdQ+9PiB0vmaziQ9aBPZbR2A2EGqYJPG12yv8v6OrNhnFcZHqoot9UV1kC7Vw
kl0JAVSyB8vBl4T2lyfhrFxEF17AopX41TB2zUSmTkQDjwsyFxze+Szj97BHX+Pi
2dt+DN9Yc8Jf3wgxaxl+k/ifUX1F9dBT4DehnBQFsujtcGjX0wU2JtC7zaIMcFr1
41wGmphYxLP4KQ2GHH7I7hpyigr3BZtn5JbwnPQ/RG3vaui7uZ+LiIxhMiHhoWXB
aHvzJe5vhPR3hwXxLoHzLjO38vNzmgo6KOwgfBttvh4ok8RqwkguMmGRj5IQA7jY
m7MotALl5sl9Ze3DMfWjuGQ1RyIr0/dQwXaUM9efKOFenKZczrHC95hj6yASLURQ
dZrTdPfDk/XAOjGby9Es+N1f64wF7HEPhhPenUKp0ZJHNGyv6glYo76yK4yYzSTE
2xtIvgTgHXwLw4TSjIU/w3YAsKBJctYQh08T2ynONPNeQbLnJ5ioMFbraimi8QzZ
2w4lSNINvHMz8FzDyrJvtcbI+yNZ7fgtV+VqyHl9+kRt7RPxMxY2c1wp7pP6qgst
U1qtW/ORlvRIBpTvMFiY9lHZXwpjXEiOZZE2vx+JF9Uv3JKZdjv0lzA8IV1/orEH
QanQ223jX6KB/JvGggihQZgUsI8V4Eq34ASPOi5ZSkC6Su2bGoWMntD59CsFhQJo
nARLiCSj2X9ZDicYy+BAzrBYD7/YofQ8s3KANCJI1/JyyD9mLdtvRMWZDQjpzOvZ
d9lS8SGicTCzAVRGQzMIISmpDWrQ23J7Y42TEKIpl+PkwEEDb/D02HFbz4kULQlN
Dpd3OgFKK08dxeSzfz4STbaSV72UDCrhfTkKv85bwcV5CDU7mD3OxA+cP0V8Ksgf
ruWeyMOeGAC5C3m4YblzfNudhSywMOj/fIfnHLBHStL8xF7Xi9FvRnkDGpZPJZH5
ZadvsjL1gWYVyNG1qe2VEq1GMmGFVPZcPWKcuBn9oTiYH/RyBjQaJ24JTZ85yjCn
ySseTHx/f9b5USAJLAwh2gSS3E76T9Q0T2/alIaB4x5K1Bot/Wc7k+EeVjW23B6m
DftXlqBn3aKYG2X4PTzZnDgoXTf0wu1Vu+70AsyG91U7PN+qi2GpOL2mf6TEkedE
Q8Nhvh8IiEZtc+9JtLYpNTObs2M7uZ+CP6JlVvsAoCy/b4Dfc5KXrjvAOXbsrFsp
A2Rt2WzUXOc3MrL6mmQpWT+ny8YfcohPtNHk9thn6ccPskTrcYmtX2RirdWe1MQc
vnHWKN9E6Mvx3CdLDReh3UDIwTUoac6kX3gu8xF0CKdSByTh2Sbxr8B3JVLVx/xp
6WgR5m/tjmS7dm3pZ1d4K1w16+7YVxc58hLZDnCJnoDFYGSc0Sj2uwSuHgbLwlHz
wGabKezA+tZSrsrYaBxIg3nqE+dhx1tKQj4LP3csOWvKCSEoSvnFJJZbf1hyq+Ak
QJmI7QPbxPe+v+g4pqgRd5sEOca/D0ZAC2HZ+Sex6256Wn6vETPKlRpNntrzEacu
bZ4R0faj4l2FNwjhiuAA1cB0NTR/Ri1s0cxK/4eQ9SRLVewklb0IcQVHWFQzJUsv
btu3gbwV3MCwGGtlW0y5XKucEzyaLeTsx1jazMYqrN3tAK5enljfqA5fes4huPmW
aiWxDDXxw+rUi7jC9X2+cTW5H6inqzPcH6s2mW++2V8RwZ5H37XSWXCfs29GYWtm
u2+g/w2MVm96++2pKOHUFSveIyA/qILArTJZaSUm5aOUVExCYHTc8DlUehg/SE16
/DRkqMyZBLk0QLrz4TcFolhM3AW1qAxgfm/cRgLgBQl4DOkTz1zQWYZf7pMVNCQ1
bC2pY1B0Chg2958tGDxhkOKntzaCb8os+V0LPDqinK2fKEeUMoH3gQU0fzOiwgFQ
EjmK+MUUaZUFjzmRk8yteYgAC30ahAJAbTfL7dq8408GJlRLps0mtad9HpIzJ8iM
Xpzl0bf78sAWVtYZQkZf5cYy+DTwKkiTl0JlIXH7mMhGb2SCUVajkcf4O4m8Y/GQ
zaYc/yhli15x0u5SXHjv6yQ369Ax/KOH2R/HSWNz/9cQDNbugi9o4niZJp8p86b3
6SARbfjWj9bj/XtkWA9xMoyBXvPIVQX/woScXRzPYDAh5DxKHbuApCLQrELiaixq
LKvg9bFX4lmREw5TvenR0vjHrHfRnvktuz5bLD60EmKSVkiz4QYvve6Sp3XpVCFz
2pJ2NSm7QZPodIwjIHhmrGvt6pAjbdqQNECVR3OIFX2T69dlgOeEAP05PtxMXtzu
Rinw2adjxK22RnD6JNTqbKLGv9MLyy4wpe1srR2zKxBy5aNrRHuuvvD0IbcDa83f
0elecgLXTiWflHqJt+AHvDnq+uGMxzKNDIw0v5NoyWHPmbzk47HN7LyIca0d7UeR
+JgQQxtdOfvzi2BZMV3/Q6BJEjtOkATJ68wanRy7EJGftt6e37+DV0RQ7IIZ1HOV
jSXmvsCeVazFAD5QSHQIySNxcOVQc+6ZjWzemSiV5ABsvoGY9oYPjGFFLpZmn+k/
gVi4VfkN6BWb3f/gp6lqLm1vJUGxkcZTnQAu9Km1NgAoEnxUlUlKgBM9r3gU3WuR
SludE7ZF0pnfcZgoIxDuG2CxRIxLLDBn6EyvAOYQHEUCt+nIpBWmgTZQLBOHb6t1
kgM/BVt0ikETr++C0BOb85tAneqX3q3M/whI1PwOkebZHRWak/YTo8s3xUAf5mgl
PZOzLH+d99/CJZr9uOQ8SUFg194YDobS9o0XhFLL5gPNAE27wWkBI75qhQij0qbc
D6JV25BALy8BU4KgIeNU+0ryu3mesrt+ATYYOoNuSbNkjqIw6OWd6NqZubEtQ5yk
CSvCqN8tlfAdd64UZZC43bI9dAfz1mk6TqhNolslFhcOpyjIQfHFH9rpdoioal0e
6MXASyjjwgzPbC8Dq1d8/XCnd139dDOvkqk5eulWwvo4j7oWpndUXbew4uitx8bR
MhsV3YwS8C5tod+lSFuowcHPer0zfyTvn71+GiO0I1I9jTIOkJHNzg8xfRFCLmdC
q4c1nDjOUQercI75bjs3lDmJT24AI5thS4b8Kd0QLQJQQsuoNLgHe1XQFcpEU2e5
evnoyUrfeXoJCom2L9jB8G9y6ITeIYrhTu3HbuRuUO15roHhtFc/aeW4RIV5SKwv
TcFureeGt4efUvTdcm6hzv0f8H/hOIbY6fyMeKJyhJR5n+smhFrK7iqV412JlISi
ckGmaE/pKTjMwjElnqmwsCa0Tb08PNb9W4cDxxy3TSn3XA8POV06fuuRvBxhUqGs
awvmL2w3mSbJaEZPO6+HT1bSVxrkzC4eAcn4ePiSzPFexAOe3kdT8XvmC0+ZLRPV
MoTn+ie4gduYxPf0sxKneVIw99Ajdfgmt4yPzBURBvQrD4OSjOpkZK7k7bBVaA7m
xAbhRYxnf7iPianPSAVD/2Aa/9WSazNGNgFZDHYDKYf8eMNui/qKYSK/iBYSW2W6
x8Exb72JduXU9rX77etoUJ+HWpfepcKGOmwPpDpTaBf6/QVf2oFpX/MEOKNbKF8F
zV0/WLmqhDw25PiV1OYSWAOcJ8gt8va+MrLC1YmpX/nd6XMMwGTW5H3kjF9Ju5y9
IBVoy+6shbkLbjPnTs9mEMDlISyZ5K8dzw8IckynA/FawpYI0JWxil0LVB47+n4b
pErnVCUTZdeg60+AoJ5sU+nrXVkwI4dJptifwXZ2Ii+2AKksjzL4t6E6EvSLdU9i
DB/y6Rw6cWlEtlShumXEtIgNNY0NrqqSYjl2aFFQ5bIMJmjcNWUUgHf+ufrlps50
JUdNdMb6nrRke4bQ0LpQJIzzRE/0kaRzvWTGIMRqA6de+JH9y9bXuctH76G7GetM
ZnmXGoeKKdiWiEDprNOYfOYxJRQaJIQ++kjml1/bq0o1ftso+SJkYN4Lt7o/g0vA
fR4mhW3CDP9j7zgEAB2cJBhYNSmuC9G6gIHPwgaH/KOjgied+5+u8Hx/r2MAwXan
e8nS54I3pUXOWj8MU+0tJJWiig9ocKQX3H2HviMtov7T9bT0JgXPhN6tBr1UxmUT
PKzXBzymF/EEuyxhuhP1/jzhvQ39qD3jLyd7ocseWcuZ0D3VoxwBQAUN52/TxDKp
w/uPpWXnu1QKYbQ5ua5byl2x//AeQjLpa+QQUzys+HKdx7gUWCk7cRZKyaTK5Q4q
OoC2gbt03or8TTIS+SJUsusYOU7Nx4mxgVqC+MnjL3klc2KwVPT5NCJkfxS3ePyP
H+QSAlnwfYQLeQ09vB1oRgQmnQ5xdvPdvYKWrQRlpfV3oFALyf99MMmlIoKmE1qo
Ea/QH+lowWFTtJNTXE1PzQ0VycIIqnhwF4G55qthBJufB/1HrNOJ5RpB/Q4mrUr/
zt7apV7TNFk0zoKAUY/XbcBoVuZvM9NXA6R/ZmhYMrXyjW6zD3OGXO7GiLUVGBaw
ZNcUKivaMRIeYmVpywtfn9CQ/U1cQY8oLyB4Lfxh2wOp3UPcHoTMRRSHnWhpJQuZ
yLty8ZJHDt/AUutACNy9ya5bmFWvuO0214PQG2gfiv7+B+AJlXY1Y1Op/sA2ic6I
rA2j16SOvr5hZNdxuUA52UjKQ55a1c7vlSi9w1oEc6WU2LSjeRQUfnvCK2SEicPL
+7rKgELJWEObnimV3gWim/9zTKBd86CpT8/BnQIyH19TvltojE3vw2PrnCu0doYI
CpdYjeqn3Hjmz6YTSKRuco7gbo2DcJiJ0MpENa6Xarvn7EejFtjnwjj3s8/6y6IR
w44ZwNEnVK6A/AbU5qXQzzO+fnOnXX7SS3P1VL/KZEDwLkMJyVpDrilw7AuTrGD3
3t3GCulk0LMyZ5Twev/dcQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GB208Tr9ObvtdlTl5Ygn76ySXaiyC3goxu8ki/cdfrmhKEUU+zBDsuFv/M7/5rn+
GXit95/mPx5udlk0PR/ngVZRTMXezeWsb3gjYxHGvuOoLGLn6KFhnUvCpoZCUQKp
amZqDeTvKA6UGZ1pm2Ai5/HmeV2y+35+KCT4bXIEdNxXKo8k9R7ti1zXdHbKPYVf
8wfH55o3sMoivQUDtf0hWiVqHhok3GOwwi6REeYDxIevByw3Umi7Fg5YBR61mQRU
QmSFRokubBNwHWqpU1Xwmt8NUINRtANOWnRE1KhTc2N6aeSY9jsunedzVJnRmY9A
cYjLmfpfAA2CJrJIWjJ6ng==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8400 )
`pragma protect data_block
lKP4gqKMhdpJrWchFxitJPqDWTyCfyzOg0Gusrkufte8ZtVgcKOYXZdE0aDq4pV2
RlYEwwRwtYBxFKWLWvwPHHgnsHDwGkgZHEqB9iUgehUdKOG4DOLqsykuPJnoaXSQ
AOGiSMxtXnT2pgLnojfI/UNApKaNyvNHoGaJamQ3sNWqtTMXPp92d75RXnWzTjrF
4RYy1OBSuTYrMMuKNlGRoQosi9jPH6N9wa14cVyBHzxAEUNAO6MsbDaMLUTM51J9
aM7re10SaZIvZZn7nAfc6+GorcPkzg1E49+Kc0SZewKFf7nv+xUNeESwQz9G6jZQ
pqPzFg150CudjQTTWIHRKpsXknZyeozomwLYa8rWugbikWn/fsOED33JJEBD6Q7i
fMnvtxzUzGCr03R0GOT5Qvb5t62CUID66gyZECjOk+3/ELl5ZnzyE6WH9cQSAdB8
6A59YZDEaYy31+0ij7Jvb9c7vyURInlv7MSU1qnROgDPGSCPXzVCqkYmGTPKDs0B
QsTpUjO/z4pgFDsPPeY3BpKvG1KqNeetU6fJIxenww+mxE44lgn1+T/OiGU7PRD3
ubRZl+RCsjAf2I/vcJf0z0PGxfeE2cmH4j1YEviyR2Ag0jgqif991YZUOLCPzdcR
pYpqqzKfP62nQq1P4HGS6+amj/dJfumYi3Nz0vH9kGVz98oy7Be+xSehtp0wO1Nj
fO4CyZXxPj3w6Og8AN6BalW+YhnJesmmpUS2CXRUXS6UVCYfi+GLi8sWVWLdAODC
ymw4QdNhEEPD8nJKIj2yrnQHMuxAHef/E/UN4hRZiMvuLznMjIGOVQcdT5H85K5T
38u/g47oyA9luq+kZ2nEvSRmvXXTxunJ3eKw+vPRqVu1YLnll6Qu0KIY4XVw2cdb
JE2PRBcCICWi3CadI1h7ydnDGCke2/w85nepmdyyfmfmzhgWENS2LFDAwwfPgGO5
CDMG9a2jtLjzit6G3LK2tRqftgekUBuYzb5s5Pwru5/ayh7FvIXImKoyStVr5Vn0
LqVM9nI7Ogh28OE/OJOZIRGlRHmXCoi81lW8I3iI/fedJ4mgyS16MjEbd6yzYvGv
Ood8RuDb9LGR4E49bPt1WOO9a4v0oX+CWf0EblBmWdEEtuDy9DVlqsrjUtyYMqGo
wHTBehuTGPFNCMr2G2viPQiX34Z97dlYyq4mE9Wjq9DKE1J0qS6z/HK+z8Tiv2Hc
aeBSkouhNu/UflyZutqbWRUxeG2vphItrHh6noq9eo6UggMGpn4cSQHMvIH9Y6Nd
Hes9FYVWmKiiD3hLRlLKibjVFe/P1nUgMFuqw/Z/XmmYz3KZ57vLmdnkJw+pbeK8
vrSo/oFNQlypClOF+6WudJPpqi9TobtfQlU8IrbiwPz8UD8LVvE2pwpN35ObWgJW
fk2U1mhcvS1Pbk393H16SIM6L8B1n7+zWnk0cFFD5RuBjg4riF9k9Yx76mqrtA8x
VRO4V7XV/xRHWdhoucl0tB5z3dTP9MQuU8d1ygn25qjKzFQBqWqmUYazMaDrH/u5
zC4srahhpGqgskvFsWj74KiGNRF9iKp1SbyuGk4NIpZNUAkVZnYTnRK4EIyaePWo
moLXLccdIiitTKDjNQWDFJRsz8RYAyXVBU8cUgrtjqkXvkmAosst6TV91PWFfiDE
Vosmw83H9c0hs43fw9jQe4Fg5/LItJtmGcTlxw02ZTo3Sxi+JH2hTyjoVVqmdRY6
JwB7jt48fpSE/tV2HL87GN06ZqkpuauTzMbHX2l3NOTkIvMd3P8HV+QrC4i1H8/6
F+gUAG9PpJNghtpCyvD+hdk/auZjOXO9Gfa5HasL/4UqEBl2IKyl1SCDnNkjdGEu
sBNGOJB9Pjmjo70hduYufSkSeFdgy9h9D2iAoUHAEOb5uT7UlOXj3VN2m7AQ4/6C
E98yL3X5U3Dh5eQfPsopVT6yigCHWt2cbwO+TyVqtFyKDWb4I7gXTpFQcs4CkdCU
MjTSS0j5Zw6tquAlDs8lW0WNkfLob1tLLmelsbVByjA37vG++iHpqZ/IYMMTBqqY
Td9X7N/TQvbU9UMY75mlfrzsyBqV6zDXLKZQneXShZUcNTcvOJ5fchzMZBTA6D6C
vS1ChpRsH6H/WhzEzA9iL4/89R3vlXXZDSzsi6n/2zHqDTK0Tz1cbOOflu+pGVNB
7XNGYJ4VcLgL2jn54Gi4zVkjV4dZLZGLYpPGnrAM2aoXzIVpGf/v9SqUKmAk6m7/
G561Fzl1MFLVDIcI4HPWmO54gyLoB1IwYFfOZ42Cr6imQBzSmzSTUmh914jDxFTa
OHVd2A/MH2VQVgBukRzOVRS+bc9xKT/fdkeFQmm0n/vi0J00HW/0MwOMFujb5odd
rZHklTQTfJUX7PXwWOHzdeBnKeLVbV9U3R1wSG8PzoKFAa1V1dVprA4a6nkgW0kc
k7WUDN+dpCI66VElQufmpslfpENEjbBaKaJGNUfZerjcTBj9ylC0HvD944Yeh/a9
NkGjOy5V5pTyEFmGCm5nzz1c8/kuAOzoY2D5r2YKNZBEXa8clxGnlwfox43woT96
j4cgEmtYQWZxaWUixjYcMDRzyXBfJGemD54UbnUfgzRDV021UgOBIwf9+oiedEGJ
uhAwXUK79k9/AFvkKYF5GZlOYJkGUYEjeQT94s9lpcigIgB6+ixc1XMizcYtA3zI
YzPwNbwvr/1DCg2WXzG3n4GYkmUQsnl33yp6aQy8c5esNf9FHC5GpdrxMyySNLlD
CNiopnN09yKiGFzFRLXj8QWOHhmvN+qR7no4YK+5eNIjml1IgqDKO72JrhKRr/Uo
vUrhLX963k/3XXO3ByB4xp40L0xNpnon4x47GEcQL493r6YTnHt/myZMwQav7HjN
MsktCQi2kPfY1mp06EV2lNbFgEQI4XyEzP6u4YyqTsYD0dIUC7jtaliqjBrCJm8Z
yuV6LyFvi7ztTSJRvD3W9qkx9nfZSITWIMq8UmWFDRFFr8S236xloAP9UT1gTzrU
vH3PHFjs8v+jXWRxRHptRyZpni7pPuwlCiSaXxtqKBi0naLJFfsV5wcR3d2yjmX5
9Jau5zCaP2Dbu4HSw/8zmESm3AFxWErIMkpA9nd4+JdMI1VQFzbpMXG1aR2qHbY0
UdY0NVuvToOw6xA5ErLZTaREaqv6eQuczNpMLT8tBYe65+Oaf53O0CK7EpKwxVYe
cQLrDBHX950O2fX7x4pqEhgoJP5UbhLKtXL5s01qO9SjqiMGryWobrH9ZX2fA3ab
LEgC9BDgjPlqgWd/rikVqfAC6dRXVPO/0lQUCXqopwJy8MXTNc4mkQ+vKdWJ1BoZ
/ctsWtI21Giy+ssmqmN6GyCwqcV9A86aSv6h2P97Cdw4fjdgv62oXhPqd4bvaWZq
XRFNAqWToeel0YUKfW0L6Xr8PfFIhbD2fnrHCIVkgGXQTCT9jxj0vsGuqXWcSoev
H5YKbCgm2n8AZtqN38nd0VRyFjSnYhXRpe0tWzAwRdEauEePqpyuQSCLnwJsHo+C
LSXCaInRRFQTqPpKxGOedxJyKVT4EY+/Rg6pbZyUH8ff+fIvgBrfHHZrOOO4Vpb5
wZ9Wkr6KdELzdi0iiFopEsmJcZHSFv5k31+JL+OBEa5R/mw8+JpDZLZeW+qMdBVD
FICJOL4U71SctiYm7bsjnkxTT1qetKEe+84o2lLDITCzVOvZ/UQBLLOCrzrYMuNU
Dp9nxW+qF3JmOzAZ0RLmJ2nSu+r0Fs2GtUnJUHqcN+YjCoQv7BCWQBcFA+PLg48c
OqyCe95N0L6x4j6meBp8V9FqiHFQ3KkIU/YtPDdxx1X1c8d5UCSKtJRZpoIvwv9K
4eRPvThDhb8MET340qbDMVKb+hoMvHAudStqFjC9C20I/+8kkK8Nbg95FVhotydM
IK1F0DAa6ZzTbmX8y/Rw+yBGykJk0JdbSNv6Nezcn5yk2+qtRcjYwMmc5x2ng2/L
Xe4RYISH3x+DtFSB4ppBVPKX/ZNQMwcNnhXIPi64msbvwld2dJL6X3+0fp6kGcX5
s/bX2wGxzDPZOjU3yWD8SyeOqtVtNj8iQ5VULn4EtOB0SH3hGZl+gqjEpOLwGRfj
6nbcw/ijccW3a/M4ur6atSEK8vpuohlVtBHdhLN5xlWftuUH5NHJYz04+zk6d9RP
w0rkeP5h48cBk7mJSwequV8HkFSqrxdZwwxslJXCrNvDBFBISGdVzCE1vsGSX8Oe
ujbnPsHIjbaXZ/BTRCGgGR5YFYMkb+9uUVytn6KIHMQWDBDQCt5Q1MDeGiNlyqoJ
EgIrqXq8oy3UsDxoIct3DcRRSarYnijKyO7RQZJ9JYl0Tq1ws93u+I5/WYt2yv3T
+Ksv9d/3SwT7nxng7LEfgX0pf7qXO2G2CYdDdBnyFGwsIuMumtki5BLcE0c307c3
gYk0FTgkX0nsywcj5toJHycLyzfNw5V2KELvjbdev7K0lu1rhKmVY2EN6FF4OmCp
GYQ6A92T49Q0UcXFsz31tQii1QwZOCFBJ8zFi+PjbMinJprfcPzsIEMjZ35XXyvK
VTr4S30ahd4wkE+I19c6y7QUD7zMJkhXuCU5EF2uBv8mdjUPjZvbyM/FE3T4XoQy
P17MJAb3Dg6zOgYl2n5rI6f7kdmh+cnXVs3jRP8S9Z53S5X4VcDRPVgR2F3Ecea/
1EMVQ8lFrGL0JsVNpih2uGnT7ma7oTk8kJygxy4C+xA+1eY+vLaWDlknGOJnlHyy
YxgMPivTkQI7B5jbq4xbMO4bV7RwjCW5B7WX1sFr7h4GpR/KCU0daCJ1c1jtzJiH
jP87/eeodiefMQttSI+SxQNhKEJkZ3WZpLiH4jlhJvOAJ9zzCFBABflqQ37LHVrQ
xEKxjMkBh19LlHLUXn8fg6Alcu3ws/EOIWcFynltUknBDDBiYcF3MXOZripJQR49
rpHW/FluRaBxb/vITt7KZQ8dj42j+eo304Ne0lYK6rFMpW3g0gQR8SyxFnj5fB4a
YzUev59wfeNF5bJguqRdShwt9pUmJmOlBCe3n5iQcxnnrIX2G197hL42aDHDt1cY
Ew50g0QJgSmCyUvgefRv9j9z2vQ+LoC28oOtUKKn/RFc09jDupAqPPOXSawnxAVJ
p4jeRIdaeDV0OiskE5rzKGq8D2nvBxZTKLD+o0qmdNCm6QbYyOZo9kcfRaHXiuIT
SgTyLE5fx2h8Geab/kEeGcMkuAEZ/+ehJhaWNkwgVQ6/f3C4/aSIOP2Pqemx1ejk
VRM+ctmPhpo7RSd/dtMd+T0frKFw542HP2/jR35kko5asNAr14qjE7P0H3SnYpBu
AShaYDu73BLnVBKrIVz7wziWsvnyBNBLKwFVAXhb3RS7IJurW0uNfF3ZM7695O9G
QdTlm1KOtL+EBvgn1x+OnseqbJQK0wrb4yvrT2zi7ooiKoQlgl1R6N5no2E5zEIs
nD7t/J7qFp+01MgqFvE4WNpahDoM3tsxXZvDAyVqy74/Q/DYpXSe5N3YqeKiiWjc
pi0htYjjNq886z9GpNMwb59hTKQP2YdhUpFUhAieijjwx/1KB/fXAKSTQksFsHLt
Bz7dfhGMspaZMBnjyQbJUmD7ykkDcacHuok19T8CA8dxrb6/mJRuooUAqVssqtsn
qenooaBQnGx/Ds4LhZsmfZ+U+I2+JElCi7xQ0KM72+yWHVrCBk5IjjFdTZYmwk6B
okXBLDVKKnkrFi02kAonuh7/G6yxrUvF3whDqhINfLqP4dcSnJou0lkDTXm/AaoB
R8SEFFfsCU/rpcxwe0ps1Cz40R7IiI0pO8ivbWETSDrmUU2YbkHplY05v93FD7db
D1jClu7dtuDisRsLZr7Sk85u+37pEOY2139GDhQwwKDYgH+e60ICkC6Z9NXSSEZG
la97QGFv3W4N9Vko1QNj1bxIV+PZy5H6ULbAjghI4gYQ2PngeZoThdsIwgL8xatE
cWnJQgvU/gaM4ZqY8Ouh6aDdqfAxTWHrHtFzfUjcc/8CxU5UzILs8NNh9e39sMSh
F//vO0rIFi7VH5nwIBIhDF8A8nbqaRFhjUMAUVrEHE2acpi5x2h+1POe9Yd3WVZB
CMp3eMBakUB74jH+59sQk/51yhWmnDVx9YkSbG9mXOi7cHA2g54OhRWYMUWVJHXg
wTqvmVqgYgT1efkb0gaSBwISLt3f2iFV07FrlfYIPByNi0TrgpvJOf8xhRpA38/V
rz0o68qARnwbK5U/imBDh0ug+YwyLA8kpPpV79AeUuJmPyJp5Sgm9uZSHx8+w2TJ
EOS0esFxTt34Rjawnhp8KtFqrlBC17ykfvOIl5r55jIrBoEUGL+W2HkYtIZCSFHB
a4cgj0HdP8xvOOh/4xaeYtDKUPQT8ZJLDQUn/5dProomgN2HsL8nyWS3nZbkR9/M
pYoiTBHn6bev9VkRdzLaRsw5d3WanXVEaj7xQv1xUSTYjP8zlYZuTaBOme9vfM4T
zMtcy4YKp9d/dGfX2wlAXnhA4ZgfTCJCNdklGj8lgKyEu7Pq0muQhXPBMOqO19OX
D3sYWFthp3LFTS9sn72UA4e/3jftbsjlUpVTRRwtWY6+lRld7pSsqR+g1zb39YEj
2Sjnxe7BBc/Ges2byJdY01UfzAlBO+TuGt2cTXZ6NOmJ0cpGvQEKnK8MNCsP7OyC
1QxoV+wn2grhoKqHSvOWvD1pQ8vkqRpoEhNerhS74cGdW/SW23a9XXK/qZJCaPSD
Ar2UnLskX/wVp3TvEZvJAK32JRWpedCdA4DAyupkkXcS4YMcMwB7xUNOwfbPw7MF
3H/goIluhh/ntFF8pJh1vw8wEsAl+H7+5HCV8MiBqfO16+2cezTQ8C/b5lP4mEFD
DtdRdhzqjIPSqhfKuSWUZEoHYLWHqp3T20rQQxID863Nsb7aVrr+JbL/R+rvfCd9
dd34BH8lJ+s5z5RfK35r8zNyp9ujLW2YiuUTNObT+jBfjVkZxrOCUGE2pp6E8G2w
cAydM2ABBGebE5KN6ZFE6x2LCrZl4/0zrq+RYiqnWgtTqB1mtT2zRK1XT7fk5Y+0
nhFZ1zxhHIdEEdNTRsoa6yqq/1R+0BXgXWufyiyteF+rxgvV/wAUrCTqc8CbIp76
nbu6wZjOw3v9qTMLiyuh9MPeoKu0roKJ+51twzQ1ALMivFkcNPWEv+h/yco+Ez5W
OFbxaEo9Sl9QrmW3xPy2+KnJzy2sWzl9rTHBRB8DjPSvErE/abo0jFbRCbNoMMYe
OxvmBeL3wYHJvOUW5Wg/3rbptAjQ1cZKZsxV3E3hh8Nvagci9rp2yNjf7e7B3ZOz
ykcP7dmBfgA8AK8/GnyGF7PfHYuxud6dY0wU2RVpT7Hwtek8KRyLGipn5CTtvgLe
jQuYA2q9KUMiW7bKJz9D7LhKkBnjUwdBcDBUxdGzuHE7zouYuNt+YxgFkRXwb+Br
KiwysPy18gfndl9xn+07PJRQ+xBbNOLo52VBLFf38oGhSiJIGEWNWeQCV36PSkLz
aqJu+k8au5FkzK+paP1KftUEvsBSQ1MKzj0xorD6zY/UduetN4puPuTWWMS1dfPc
7UT7k57d6j4lI3fIkGOvGRujo7edelBBVakx6yO3bWEsGXRjTP1gKAafzCwOj4Gf
YN233NljNcRLFXV8WmxSpYJmfUBD0uOPzrFRYSOcFdvi1tvU0MN4kVw5euBJ5XUl
WQsL4vMKMELkH2wL7OpJ27HWyymZjUwhoRt2wUUGh/UioR7vW/Ex0yzP7sL49dk+
WmiEQGMZGn0OJShJhEBORtGQcBYXHbQpQCSjWG1Ud/ari+AyTqjbqSoO/tnJbEuM
+UPkMpifFIlBhI0Hq4/VtftkA1+frAKdvdFY9Kl/Y4nnf4AqIBiVMI9Ov1E0JOFy
hxwTXleUyopSohlBI/DWbsilKxJ2NskFSjQ0aBxwtNF+rZ+2Xujep31+BeHBr4/7
o2ab/mcCun/PM+Q89TxUKIDH6Yc2zjkdKK9SC7ZSfs8duLYZlxjk6ynkDR31JBgT
nhq81oG6IyxomVYOwV1fxWMpMdZ7aeo75+Lk4vPBltk5d7Hd9HkI8gVxeogxeYt/
oM7PdnnismHUqHkBSorzGi4V+cswyyO734HmaEZjCQkZ0h9kZqCMrQ4rBHDixapA
rUl/p77DOjNdpMERA12+bElmccAyuLTniy0278DKJLHtPIM2VqQhHmKfM3PZAaNL
2voN0BRrhRf18X+XFRz3PktFZii8IzPJ/xDBn7jjqirccARtB5NeygJaK9gIw25k
k8wGaLYYbzvkTWI6BlZRISthq/EbEIjTvT4cxwRVv8vFFrMwZu72UzWkr1b9QWgS
tDy5iY5X/jAHsoC9opXoDTtnCLEOB9Zqu498s2p4mNdqJpDQ/+xCq9PFemRWp7h5
ZBMDuBxS5mazC5PQNnkr/K71Ck+8FjT0no9HWW4LZLw8th7DGsPaYufbJtNthkB3
NAkTql5X/AetYBVf5v9R8Kp+AdjZGbP7MSyFvTFQ4CpPao40J0aBdy4qEKR29Xe3
nB/vY+7/AQ4SB9XwQm1dBnQpp7TmmnGjOrNH7aqnrHqG0rMIw1NsNLhiRtzqpwlT
mF9CB9NzTi0mcXfsCD8jNPNvpKwOejdjQQQPVArQNAhZI5k4awEyyHvFUrGg7Guu
faugN7APlPW7rxhqyIkyJ5YejN1/8hsoG6lic8VHXlcB69szb27XFeKc84LxSkcM
e0ha6PRJlQ3x1/3KXWryjTaQLXoPCKgTzBBCd2F8Z2ePfLYDjAIJAe8FHOs6tS1J
+K8+N8adF/zn2xt9YGXnaFSUvbEBQLfkhHiZ0mQ9g2ZL6MxiNB4yLKplo7o1n1pE
KiS0FkJKy+pf7yqviEsznrD9YY1gi8qkBbux1pfdRikSUsNcdBMnvcLJmZbz875g
YnnoE1Ggu9YdaJDz+rJ/JgwcccXPfSvL/3qtxKAnvINjQDlNxuAmupaWJsCxsT9C
mVdaV/j1g8QTHqv0xyo4SP1aObncn62yurWHNVIW+Na+ng+HaN8mv3niXVSEznbH
UgSAQJ/wTyeILWb1aydeKYMbROIhIzcVyhMX+0oIL/lPkiTuc21oPn7xF/G4HyBD
3WBxRDqDY6C0JBNdQdvTLZXa3PWKa+sFqjQFzN2u7439dNEs+1RGCLUtUlxJiszz
e42ferFZPjkrG3l4GSxYVa+XCDHIh20qTNsM7wS68bEDRTNUAQep6k3gfqiPz+od
ps9jjgEzs7cPLFVd80Gr50O0MSxZFlDU6FuxP1DTiM7zgtGM5IlAkrFt1edkDSI+
3K6O+FrCmrFgC9CORVhwvo3fRqQuUG+7oIhY5A1kOM1tIPkEUuStA5l/2ljVpe/s
NgD2Uh3k6OxYgzN1MyN7mH2ShHZE6gA8g4u9qe3Eg7eQ281NQ7+ipSmUJC7aCqwB
mYEBObYt+//zhmmDYFqpbjKAHJL64BiP4UrwX6cOYAHjf/kxbA8Ci7QqCgUEw2cp
b+c3XxtkiMNzM2VBktzwCOdLdIi+FzZNjzn4hKg6F5htnuGn2pMhV8jLzLb+sA4t
43iEvRUyO9+5JwFnGOG/Vu/e/qp8dRZJ5n4OtvSOLPWi6K/QbfSNqH/GuoE9IwoI
pW67PMx8E4wLby//ABfo1SUol3jiLxlsYtt0voEN7kJ//lfckziwziXzlQRdM1hu
H5fMvUqQpLKYgs5R2lX42B3Z+Fm49RsJjJ+/n/ZNLVtA/GcUoTGySHN+1shYINx8
IlzPTDVnuKWB5TptI4tvG6BeeeOVQboH4pZnXb9pRE5rAG4FmRr39JdXUYMvr4qr
QBK8mZICICtrWluZBeyY5QRaqN1jLNj0ycqoZ1Vj4CAy0stdpIuUmYsNpJoe6CvD
UAU25ep1LG5dwjLGqKd/wP58mV//1l5cYthAt3R3DCGOBUyGueQabBR3ZrgF8NIT
oJb+BUPS3sFoCpuXKsQUQrufby/YDDXvQDjO9NuJxjgTY3+Ktm03q4ZYZ6+3D9iM
STeGwbI1yXCp0lwXtHzaMCNkbboIzykdoScZfZXzc8tYAegn5s5+opnAINm7PN21
gt6FKltQpbCdGXLgN6AM2MXGJPcrG1zfUo5MYHauP+jiJ7nrPra39WSDtCoWh+MG
SzKAY9SrAzb9n6kOR2jQoBxmfI6eGFZeel4UCzvo34mmNw8Ql46yl5Lenzx5TtnS
lHDuk5DNPLk54/HqRqbGlzuuIPzuTvgZZKWUnzHrf14D155D/CgDv9yOL+vBI6wb
rQV8A4Kf/m8DH7qCp7bEpgf5gBgjfs2IGvMRUIhKdjx/gTjDjfxmvS3vdT4uDkLN
nRzWCvrn1S18TAfJhjaO18S8Jl/NzoBxEW4Xh2Z/3LSO375B2miKBZnIowuxQxOq
5LJUhmP4pL6q22PUAM/nhijgNhx6R5RLmN3lm5Loil7C2DcxmcJkaPYs3VMofOYo
HiAOpPDgNqNbZp7II3AVn2TDD5cmC7GXo/NBjX2HoUDhLX0iYfPhADBXglhYeD1i
84yi183U5t2NB7utWsGLSWC3Oiggt360nSRQ1eXB9fSyew9i/gLOY6RZsvK1Yq2L
jooSn/MBbBhXo+R9FZIb0gf1nCRqsvgikjILfliS6eR5AgIxtyfhTIMNp9KIlR4e
ylbw9VuyXnOODJDqGnDQUNPIFj7tBXl1Fmuk1iRfbtm7cAgVPBk3WSLnzETtPmv+
cT33HU77aQWY/r81TV0oXhjNEHCcqAZGJh4f/M4YqGfE2fpssd1pbvvc/GZti2LZ
f9Q9pn8JsWS4ZRzZUIm8mfV4ni9DxfY3gj2ar+9AQbst8jwlsGRUt9UgpNt+yAHA
t+a2opyxInf0QbHgIOv0IHbrkbPxb7R3Nwv14D47pAD7eGs/ULUpy3jolyTuEJ5b
+QopkQe8kxPjIToHu2UPGAnzXBsgZ0aXA4FKDxwJlrvfXkSiinQNhqRINjPRzAEB
syGnkWrY+jL8dfNSQ1UjHBj/wZzDaa33jTLFWK1F3QtjPm4ZA7GhNhzcxS9XuVZ2
ZClzTVyT8DUSAm938G8RELvvmvgGnnayatSCcrodsw3KNAZ+EjDsyaEQSBJmW2kA
R0awEfNa3VymDwG7w+uFdIKSTR8ZaK3RHzmC08Gb5NTDRLOAwPUdVGr62VQRp/Zp
jUwPpQ1+kkuK0nSVZAnwEBM/OnNEAJjX/d3y1VWJwvLrL1cI/M9GDGhZcAWPtOum
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ROqXtwu799ia0dmbVw/atCTlCFAGma4c0mmYYJO/ro8+6bk941IVBE08+Qp2rYXk
t5exQe+VdwGyF6J09V7Fbl9lNsipgqZ8+vwdCuP150fq9lKNfC4W45yTIfG9KQ2+
vfsaBzcQlyijhzTpOArh5nGkSERru0RmHMSEeNnBmBR5U9E9iL6gx9zm54xEH8Ee
iMwY+OBM9wuk5gXC/hFaR0VXWSQWln70iPYs+nb1miHgx6C7NQDshSAgqWvC4acl
g+t2aFCS6eNMtd+9hQcKs1QFr94qpRD1Xx2g2Kd8Z8c07IM0RAb+SGM2bMNii7/+
pGfRSOdpL1G2ml5QNmIoyg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9840 )
`pragma protect data_block
iG4Nj03d8fOBgAEDxZMq5vbV8Prz6jjqZ4kpE8dw/LfTnTt3dhFaXQUt2ex/BSJh
Z2wXub0aS8GxY1PoTKYcGC5VYEKHRdcYC1cqu1E54SYzvRNaDc8cRvxAAJRwH3ZM
cxy38l0EUWWh6DEYFfUosmF/5PVWxKpDKohOKrDDek68zWU8Q87RUrCmFMRlw848
3/3sS6QTa/X2qyXt8Vc9e+uHo+zKFo7LUXP/2xW+YlX+OehJEPjVHU0Rdhrq0mXL
GoSxll996CS6NxAb3EsCKqHmK1918Nf6EbH0qrhTxj8BuTv2ZMFW9wHb7u341cxV
Kh+B/DozIW9nzF2lkrnvIkCoc26i2mhvfXWs/vJ6iyO1viB0o9PDFVQEP6bSftqG
Fh7JK5xhKAuaUIZt/rTqGOHMwCmRxs8n0RohRin9sgXo4xXAfWVpWlUR3NhnrLOQ
kJlI465bOgAXv87pTWgI577+nycyUkvc3gMzVY3ybOkYZJcZSqkO3xuTFCnk3bd6
V4NIs5ysQ1nZ3xrEqFh6jENfluGbkILHE+ZtE0fQSs8X7QbOIHhL+BE8CE0qvsJX
+KmxSZ5PWSkJquJWm652rs6YKIwizMk95ntjinTfVyVcnPjjGI6yfXzUWixHqLz2
fS8zbym71riQ5NBX347fg5bJ+gYObRz4YGhdSpPdBO4NTKHBW5MYLktaGqUTip7g
nS/N1aJMa3BCHAHsAvLnLTJHT+0iM26EgnXlkEEYB+jYJh+ox+s9wvq+UI5qT+Mi
OxnlVHaH4wgtaa39NET43PZdSfqDeziR5U9ejFO9OPEQMyI/D0NqMHKQG8l5tM7I
8lnOfjSRb+D5cAMxm5oEsWkIC/TiVH1e8lFtmnF0Ep1bQx+UrU2xXiKuO1i4+zvf
sKbBUGwHL6gGWez7SfNMXwfKG6Rfk4/WocVw+3DH2KfCagEQxX8GT3rHRCHHpX1t
GWwodOYYR1gV1IkRXS6wGYz3q2mf+HyD2xjOxDhi3ecB+m6YkAngiRs8IeYXVCvd
cx7Kw8MbBklZmvZ/1d0bg8K1b3ZqdLIPYFwYYwAsBULjmm6ODpKDpoyxUYP9XYTc
pkjx4JsKUOCPzGw6hdwGw8GB1JKBBg+IvWJrn8hUcsC7y8lHG1Yh9ORw5qsx++56
FP5Cu7LSSrniWg7ozMhZ/94W5IWiNTVNZXEkNtp8biZfKbPqpkMgTBao9u3e3guG
lwX9BXPStK9uUmeBn5JH89K0uwhIFrbu805X6FM1TUrz0Tgk5/ca5jKuxhDqKJdB
K1hrrGdz8+lwj/C5YX+aaRKk4PnS8mp9OqfXTxwhPdvALqPM/A6YqmoS/TA3paDd
FW8JU7x0eJYbCo57nA9syhXhukUIIjFSJaAJ/EWUqRk1GxEokBUPmxA3eanwEZ20
Jh5a6JqZjq7mKtpFL92IyByKJnYIx9L4+4LRcX0OkUhga0SaXjIZdKToQ3nFS3MO
GzrwvGUorNyApMfwk9N12HLdsBJVFaVLUBWg/ytqySASGn/Fm6Sg1s80U7c0VmZy
9aGahqMGvZXz7N4FYhhxZkRdCOr1xVBdI4GQ+X6yxjhR7eYMKsqZV/VyAGrs8iP9
t0enUgsA5tXg6G2CctGKlMPFEMEoaiTUs9Jb4TnRQb+yxRgq7+SloEY4mW+AG1MD
J4we28Ux7k6yMcK09PTtRN9YQTQprq+uRuARFJtePsa59GIU4ZKwEjhN/28Kp1fb
y7KngjVjH9V+ONmQWac1hnaOzjDBxedDtvn+KWoWFggDnVBAO+di59/lrXZ+tof6
CptcGWdQJ3xwlb0d8BAzScDssdoC4GmsFCD6VW/Of9Ym+WAu11hwhRdyVayAxbEM
RwFpEmcmgyim3JKRgrZF56qUIRBwm6Gle8MCB/kIIUcqkokIQU9ysbzvexFvgctS
Sk0zCs8+4ugKSR3HU8H2ECXKzUJrEV5B9l0Urh0Ytvao+o/eYLPeXTdp7lE3adMX
3ayWVHhyaTx92tgbhfyrik1drwF6BC4JWf9h+2QJBDnxnqhyQ/sIyh3iO2JQxcym
tlr66iuwOvAgPEZ1rKhOBAerfOwHeWj3myvNp2E8E8gEYmvtaVWg9vgLu9+x0nF3
muxuyPR1IvYjKT1zrDB/pz2WIfK5trTN5/7+sP0X0MWmnQ9lmF70mXhU44XdaAod
/MKtr66qUEFP4YOD8AYB5jjRS98rzPwHJfn83tlLW+xNihQqS2s9AdXtJ29d3mTB
sD5tpoC0+oHv6Jad0OafR5JwRvItH79YKPDdZyPSCE0ORj3/b7H3ZRBONOQKvNyT
kTuFujmU0N06JYWkzyUpVmPCrLsU1aKoM54xO0QiZoEyvfb2K6Z2GEcaVYH3hU2V
4hc0BUvYN/HuGUXk6SWLxQo3BuDqTW2goyFWk/FGllC+S1BUKcOwO/RVJo2OKpCh
IuNJ1hMcui8bV6VcTnlRRbd3SrM8WBi8fXzH/Esx4DMalFrZE4Wa/AY67295lFur
3mZXOUXgGaR7DRGhLLlU8mOfY45W231qLmifQer49RcDWZl5oamx0M659NDl5KQR
rqlSMvSCYwY4lemj204vvr2ZJqh4CUZRzXMgfxu65k8pByOD5UDyjwmPDTqlRymJ
LuondlgaYJlE/9FW7owZghYmiF5CQgs+vffADSexfhymXup1rdhe/8DyJImm+g1g
qyqCw+EL35C3mtAvsZN5SsdOVZfdSHqqekHTlhjiMrKmvHtaJ1WfOsAiHXnI6kUD
V4nKeC31NoJDQRDqzs6ZerkWu0DHb6f+IYu/EiAlOxOHeHa/AkvygPbuiHZ8+yZ4
RvusiKqOOtjZNBAQzpum6sUt09jd9g1QKSl0C+jrmhfWO361nqYYa18VNuC0DvMR
SzA1du2ETfzAghOXGwojOlZIrGu4tDP+jR0UuWANpf3pFJWocFKNR39LZoOleaNx
lt8xaijbrpDs6Zd4qHsc8qEsdW/qCk3kpT8j0ko4cho5RlN/cxRzTxSMm2GkjfAo
MOcU+k6/UGQOfiXjU0HCydyS+9iaKUF5eceWJDcsEtsfdb8xo509jpXwVbAkWdPc
CiAwuitvStBU40/LpEdoLdCdPsd1rfXCLw61XmOO2uSQ8cxXn86/QhFwYX/XKamm
b7utCOG2fZJ1TrCErIeclvmj9DQ25bus2VVBDyNzmfZgxXVt/3JDNYVfp0N4CpQc
V+fvPpN+ojigmgySV9XQA3Fzp4+GUkU/0gBYNGMjYKveIFZOCUDKPWaP3y1qUvwq
skokanHfi6NSO8aCQdzsMNJ5BxpX/EfV7not4AmGTDLgdGslgcVNl+NVilf/O3uK
g/Bg3fiT1GOGyG58FiF2JTxs+rWuiKx3u3NN0FvK8xtcwOeVpJNnromRxr5wQogH
GEilB4zKc0HqCNChZlWvcqhXOFbVcc/VjaGMudfZ/pDFva+C4JDZb4VeAhm7fBLO
Z0s+skGkCtS/2YNLexDPDLyPOfzu/DYaEikulBjYYXUXMYDqWsXDxeCfjkTPSPDD
cMWZPzcq5paxSPcBYTyGR15w4F7EhR8Yx3VK568+j7WM1L1NLZSpvGxs4VIF+FdB
kIq5arwxKCjHRXKVM+w4TZPIc98zffdyJBZudm3eCbXiHkwrZFvepXviwieOQmF5
yq3nJx1o7ec4snP8zLK9/5vpzYJppuhfmVdQ8h6HNnKy+8tWX9WV8rPtbwNdnlHN
lJSeHwnEIC+kUT9DTWkQSgoy8mrUjtUedGUT+3NcAU9ocey3anOTxX5lw+cLjD6Y
RrW3qxJVfsB8x9UKHNuK6lLUYQgnj0x21t5OzjJt1dUWaLhnIF5NmiQXO0RziEpw
ao1XQXe3LKqdlUU3D8BP79Rckd1kVQ0qBG1bav2T7Dk6UPJwqCxxCGPR7ukf6ip/
0yDiXaE1S22VRB6W3qp1J/ds8CiGCzTpl9L2bzkN/TtDDgGAwFyuSqBB6T+pWk6Y
ptD7y7c7kYIDQZFuIdlKo6iXu+hKak9RMudTF09UvaUey4QgwpDkmYe11eUUJycC
kjb7xRynmDgoa7nA92Lzl0ZqmN1UzkF+ZcX4RqFtnlOxhQU0Ck4XzCAcuRybFwWd
tNIrwPc7jpHs2Mah6JkckaQDac2v0o8g2EeZBZiJ4+g3ezqagpwhiarDKJ3Em1dd
wA1VWVYXe8F7En9U1dD8wUuKae6M+gyg9SUnSG5fzpyNt0Bph9C3cu9nYHLICsrl
gRz8pXDPoVVYmGnph3wgAeBKIvN6irg4U+W1qzx17Y/o7xO76MMNPNsA7j4TFlH0
sa5BYk+/jmPxtCKIQCAJRU9dGI4tQ9nh/bh8xuKuldjtP/OVhXxWjQ5uXMMeKb52
EoGEqmCNu8GTrubYQf/wM06RzGqoOtm7BJHXkkx2QCqrvPeOkkG4pif81ryFWk8U
u0P5++NOAhhn6Ta1jogwT7gncol4UM9I1BFhfncOMzL87eY5gcmp7KcoTkNlBkNh
5k8ruuYyXG0u19bntb8YmVTD12RbIglnGBSqxefclnGZg+y+rNM6//QgwI/8wxDy
7+1TNfs5Hjj7vbB18fQ8EhjkUSMAzHrLwALlGUJKXVe5yhvhI0998g15QtNlwovS
xArf6xMt7eTYPumBXoUO4RDqLd53ydXC2wu716iAuSp3LNprEVkl8v0dUxq9V39p
sgQXPB1ik9LZw4xSLf8D1CisZMgMOQdrMABL8HIY15FOfhSU+s/DFOUOz2VeOpUc
cMTCSkC2uO+3mOEB9N8JrEvpNa/2HD9qtw+Cq4G7xg/YuxqW7TlrYWigs7RNcUTQ
E3gMUTkuhK7Gtnn0wZV4q2z8DY80P1ycfPZbNHNHeZCsQHyq6/Rlpngo/UeUTuC/
hvXV7pE1lYyWJxA8qa7fr5aGT0VKfIxF1vygT/tTlwjJJgzjytVsQXYvZHuOhmgy
CM9ldC8i54IrfuX66UqFzbL2tA2nGoBo8ZyPOopFuB4GdMOLjNETESKteoDxd208
cMffAZ6f3AHPgJB8eyiG56rtXPMLbSwnXEd3K1uolimn7FAUSCzzfVzxyku/d11s
0E6idiSBY0XwazYwDB4lt+ktoTtaOHUMu+BitHlXKOMMzJjvV/pTeqlezlibOKZG
gNT9mEudCRUSEvfvJwd+pM97sOF2+ksrt3hXCEG1nyMV1EqN9Osf88udWItMfvgq
sZp7/+ni2u/ADVUM1Qx/v69h2FTOBwo95S3/x3TSWbxTF6VoEN8MXALjAFNmCn+t
DJRCc1uu2cXEiSxSMTotr8k7GR9wFMzQXQDpiIrRZPCbXaK8QVCfVgQBenN5jzCv
vx41o+aocvBiB8iToXHyPYN8lsvAO36ETnTwaGWn+kTBUpjRjCg9u+EMF0R7gZxa
FqLoxoGE9H9HKQkoQPdURiGZI7QBMdvUlOM55lY2YsrgXjBawcbbg8VonoldDMYa
GBto3Dr+ysHOoIG80xnhrjpa+cug3toPkep6Zx+cHEyIm+eylkLoIiSww3NNVetJ
YRarkbFKtAv82yIrGo23mMw1SI8kdwPcoiRPrjxbbk5Zh6SkC40xXUtUySc8e3tq
BxuGRWbBXKY6xjOgELLuuM3NQTRLIWwHu86kuKY5pl5yI684r6qNUr2BdE1j7PDn
y5qIZI8TbngoaweEA+dEKFU4opI0Nffacdr+vdqaBqnkAB7GCCUFbdon+Cu1Rp+w
0HsJd9Op5tQroQTg2Jby3kOX62MfZhlEUJV2KDpSReTjOJER1bxaVCNnzTYAVa/r
gMCKbMqfLneLkIUsB0TQhiMIDVQdfCPzM3Lhh1evSrwbEJuSSOHeFdBiAtMqjY9u
w8javSD5dF/g+PB7BKXmYPFqLmCU9wVNpVbWV5VngrzoFRO38ueZ7TFZJ0FLbewc
6luJYzC3LzKoo/E9TYS2RwkGANW8U5QxQ3g+57CE5hP4vGIGKX+kONdYcK5ha2AC
oKVICiXPYPzZhS5UAp6dTd2K7dPIAOHBkSuZMaLfwKpqK7aa4tm5c+0pIDzJcwNd
vBuJNwMgsTHl0Q0S8lxk7+f8GgYUpML+EqzmtYT0OSTQ3RBa/6KKC1gwyGcEmDso
YYCkF16MWAZc0SRvo2fqBGGwLwwAi53Cd5x89GWHE4fa+FRAY8DBTyfrIr/0mqfp
QLcJZxJbBqOphxNs5PfQdw9hYRFEZ19DUsJQ2o4kUbRhPyHALtQFrpwCUMfnmQZz
AVkmgXC5LItykzy+RPKxRNq+tFAt2WnvEnrvti2SZAmDG8QTeTByMmFOb5sq22IZ
QDYCkZbJ+DikvywoADgsVnm9QzMr26pu8kf9ctmBUn+4Ax8vW6CC2a5NdTqyzbEu
w8wifm4JjYOdUZWvCUQC4c+Q00d2XPFd7uFaT8eRxstpBlN304R7udPINATKUi7y
8g47OtHF963sjswvw5b6SmU9dPS5rJ98qB9zz8EdGoSGNpzrQFObAPF1z2BRDe/m
l/tjeeg03ixjFCAeq6ZXlXe1JTmNHVvjIBCqbmRVEJXHzjJgnwsK5Ib48M2kTXlN
uTHV0ksmXLEKgtQG5XLOO0WsbO2zddmbd5ydMsdgsGhplE5wg30481b3s211aAtR
LRO1B+47QvvTyAVLptPd6b6dBj+yMTrQzJEI94dG/xaHgLM9JHVrtRGWTd3VxVg1
VHsz49pOdsKF3qmSinbNLIZx0z2Wm2SqR3fCE+VkrsLnBN1NpVYujfpYNtApdjuK
cVbdoa0UAuAmsAsEFuYzL7B3rXF1PJ/8K2MhAvNYwX1bjkdewAarMJCk29t/YgBb
zwk1BQ9nnknymj57RltiROuSujtJsn+aPBm2PKn3bPwilzTA7RxCjnkyLIpXzacv
2shmKaNjPLXfOBvQPItvGMh8QyJjUgtWkJ4PekvJwC0iHvWV9Nf7m5M79Gp1pfng
xim6mAENO6g/pD/eisB0yXfOIJ305fz+wRLmOpc7B7kowWZ74YVQodNbSwS4CCVa
yINcg5giZm5wNUGe/tZ9aWCLostnVYVh++WZg3RdazaCVwRly8RC11ITnqvYu//l
K65wt2bbMEcGKLXU8NcImIVa+9M+eFlEOgMDDbPg6JH0mNeJ5lZbPuI6EoWJD5j+
bG+d2fBPsNEz7fMVdaUSui2+y95SYIEYD9DpOVg+rp0agulzdsfGye88CFfygvNN
AUXVrHW8wzNKDGnhEFn+96i/iqO+GX4K7qrV7OrZaX2UcleINs7hr33NWvBxgSB8
2WCrZlg8dJMu8CX9uvADMiCqmnpPdmwRh19sEeTS/vQwTTSsNm5uojNMRUV7kNSH
nPir2m2c6tAMDxhLNU9/ODobdxEk8XMDoC1tWHe0LFVFUIJGV5vvyxVOapbfjRQg
+nY1jo/0NqCslZLfOTYaeuLL1CXLLiLuhso0RmZlro0xj2cwbbF09ETY1KANlAS/
lRTIDQBOrSgfLEmzRxLoBbTh6Jw1sMgfxCNALI0xid8pNaRkNOX+YK3Pvi0KJOiv
5vrasH7uWDVbH0EySp19sB2UYYr16tT7Z3qdQ80rMmYh2djmXrArkObDnPmyQ2hX
vXr5CHLMzpDjzOlsejGflKqO2VJlLvqpHTwnsm4X0I1MN+Jn6MFScyAD/M7Qjy9x
Mfeht2UxerNr+aZfMPrUi38swDUvFyXwfkhHgrfLtfaNeJEf1OkKRe09qKlLvLHw
QUtKuXwHZLPhHcV5CoYS85MC6XwcViq0tPr17zXFHgzieckASfwgZIZtILrBOpo2
CkY34TF7+PCAPL0pENytecgqUx1UBodu3brhQNtulv/vYeV2vMy9qaRTMcunl6Rp
rnHgXpdpcbRAcYDbiU6nJoLREelJRaTsl5urPRydhx4tCAC11RSt01k3OnU5PtAw
O7dHj0E8kSys/CiVmA8vqu9+vlcxw5qf6n3hPh2eFso8yZlzjWGzqNvLlKHEilv0
TLAb/pu+K3kKn5m65kJYWRuFduTiqYDOcM0SDbia8BiZvEvIXUryElGiecnDaYVJ
iyVPa1hB5XE9fKtf3+7BDv0SJZaQu2x5cxH1M1x9VcvfCP4hW97uum7e9EgzmKaz
HsdGke0F0TNiKrnjjOy2SifD5rpxgSy/+QlltRFeOXx8008QYK7oVAGyBparuyDe
qrpcFjNrIp9DENfRtKwv03dVq+EBF+a9da6UvaaHKya6lxolUItKo6DKVFjJR3Na
c8nj22BWpCB0iOsTFrusTHnPC/wMJSQgr+PxdvmQ/qcqIPbJyFmmIBFZu0heZfbi
O+wTa8l9ddTp5avwiOFZ5nA096ZMyALCzIS9sQZDosj6kOAM+GZNm2FNrvgNoLER
lR6hM4Rujkgn6akuLw+OuIRO99sv9sFukyeWdsepuY9qCl9fWGYJm8AMdhPifafn
P5wwactHy9o9g0JApYkiDgiILcYYmmMgeQ4ZzcQbXn5uT/LowXAmhGbv8NEozOdN
PHF+LnmgIzqyU/nWTzMqfVcS0bNIs8kD0QLqvsIBLT1GdSRKiIOSKMQgLOln8SlS
Swz1F5KtksnPyU0++yk94iaub979/KltxWhth33VI7pXBG7uCXDRHbWC2Ib9xOk2
iuMRQcdh1yl9RTHxLSp/NkXuprJLl6BM1ojuCTgxnNpBc1TuRBbqwj5niBNXnTtJ
TRq1mJjYlzjq1Ca4g8JxBbvGpQhmGtIAyveTIKhCws40sHllx3LUAYLVKqCy6em4
TnOuij9/ZJB1qDBkaziJRQoJ/7uISe1J0qe9d98hr5sy/8ELp/4LczEnl3WBcrIZ
T16MNwAUmMlpqLd51f193qe9bGhG0lMI4m8na1yGxzEp3vwAKX7qt/OdQrRTjP6/
6fCuGeKCHrMvy/dK14nnCQ69xhD2fo/RFcf13sY4zG06kbJaZCUbBOD3bAeUj6G3
qqrsS7JTLOGFX6SzetlARP9sg0H+BzanxoENPpzr1LZL/HFbxtrCb6TBdTH6fGrM
/QvrRqHyAEjxS+Wka9/w3si6ndLFj6PuHIaWye6rFkYfqrVdcGyzRnDy2ziYMQKP
gGgof+9QkVQHrKO3cQC+S8olQ844ua4Jyc0T62lZSzzN1BWH5GyFfMigK+BA8URE
fpK4363Rhh15mrNiPpBSgcCW6tbc2WFZEnqfvroEmZfemkCMu2BBnOQ1mksYM04a
7G/jawKED6JJTGDyEqhcdYTw11YNeKK4+1jD5Lbhh3xZUcuj5iP+mHH7ujuI5RJJ
tYvlrO+7EnlZS40R/K0v63E7+Ri1kOIRtJyYjdl6bUTcPZk2PpEYsSrnwOAbuUUE
6w4bNzGrcwXLlukONoKLFg5sa5kvFPtWB7f9PMvnxpSp0l+Cgk0ha4tMLlyjtsQR
lmI9Eom15+6T/rFaQOWhCyEa5m9KhknH83gFA8I9kAudpxMhgEui/D0G+cyPKfiY
hf35IcPlXA3soIOS2CHXGx5XAwdCwAAvH4DnCFHUWwzwSBW9xfXq6Fg6s9U7aq0e
WlFx9S7R1JjxS87Dlfapl4B39B0Ryh1a2h6T6dYDjP0YhQdJqeicuYsKFU4XWLNd
vJeqFmooXPc4Rod04yijiG+l7kVUgQW/X0oej+4GTeIwx8xZP3++zP5kG8CtPexa
G7c/Rf0Q0OhWUf420LZZoa1eR88LLzFfP2/yKgFFQuaSxRAWv7uIVHTbP72o7Zum
1uAJJQ0M0Bq+QCMKmh1Gc9iUpLMYXcmMu+1IadX4ueGWMbb5YJurbQ41oU60jJ8r
O0r4s/3xBTOlozSv5FZ3jh4E/JbjUX652OpvAaoAdEEqdLWVDaHD6cNV061JHU4c
otrzFCZ+RibhzYgZljLnfYkgSvlFq06ZP6O8p3uozOmOakoG0dSLAwmQAY8uqw52
OeHE0+DGJANVWX1bnVf/9aNpfy1ZmCkZ5u6n3KWDA1B0cK/BBGBF2tXJcBC1DoYO
v11/H/GtDQQin3fgAJ1y8obdofsqEpn626/WTdKHCYXGusVnz8YqACFD4bXNqv/P
r0wkOkgT3O/zrxiJr0HT+0XjBauZjTFN6+zeHZ0VZRevVIkgeeskyb675fg76PmM
xDlD4DxnfZ44dCbfBWGOQA+3/Et0+KpAgrCjghLwGVVDxTqM1yLzCglpUHt1JCF3
fuOKMEL4q10d+P+Vi3ubPJDVJa/Nru1FHngyj9OrERXelfb22NfV4w9O/vBAvRCy
UfVHH2B7mN8MOJv0gINMw1tK4yfK+GGel3P796waeukxVDvkuEjG1O69BL7kFp30
JN9cLK+ROoKlZEIhEyrySlM7Qc2FpszxcyeuPB8Dr73E+Mul9kk5mXbr4S1dNytt
9D3+6BGMlZbZZCyDRIo5DVilrBvn5n7nI/Pe6El0p8CScm7f1/X3o/QCLn0PZuZk
kW/u+0va/8ywKJ/JPdSxsaF2APfkn9GVXLEDPaxJlK5wa6LoFV5KwDLRwFhE7inc
q4oQhG7aunOdNIRy4/tGMlZdtZo+vDshHW2GePcr66yZ9yD2lwtxsw4lVuw4X5Mw
8AB0cnQqBzjca7SDL488Ug0qmhWrOL/kv1PaPC3TtVoxUqKseVH8P4LTJkWIdjHR
4XnS/NP+idNXgVT92+p6DilhNuD4kQiLzLLtiLu8Sug1LhX+2LXzohcF4Ej2xn7C
doQNJCRVSf3wgrz7Z7gSj9EnzcLeL3cqJE2b5bE4XXFbgtAhFGc58ixQ3ciwe0UK
4hSDib9vOZWmQnfBX6PBRDgSOzqHApXhvv3udDyH3nimmwMdKqPlUzhYB6uhnQFn
TrHujy7kD3+UZZ9zQ1q/WMuLJVZ8PgOJFakio7xIVEEgBX4+RIi4uw0Ww42NpiBT
FmWtKimQnnLdu+XduiWgoPaeY315J08IAh2btMc2wnW7zrU4Fe21wWz2EqpPLD0u
a6sP60+K58bQgHy4/dloa/jFFIzqg/KEpOypA4XXStsZ1kEuB3FL9xn0ECnqmfCn
jQKFCpKal4uEApAKxswDoXTRWFXpjrCBOjoNeXl+EMufvopPSeaLH59zCv/06QBz
5NP6Ah8YaPJQ/SQleabWb7TEHJOU39VAJAwhORY1Ujx9slcaOdLYGxjyzhmqzHGZ
oFZ8TxN3yk9oQCUBHs4WaqV5xoYPJy/019ZNjiUP665NBSVG73aJHYodPN4TzQJI
KP+Bcb/uk2tK62X8g+BnQjalDdDm8T5lSMziI+0eitfe2Ly7h+ZIEZQ0fj9bIW64
pe7KwB6natVflahatLQTGBegM7XK4G4g2NHaOy1EjRVINIQUdOxfcb865mh18xho
a09tbHCO/urziq99K1aEOnj027dE6UNIKkyAXihmrUYaJHgp3joP311mUM+u1ywG
ip32cUwZcaFCQsl7mVVAG/UWjO3HlgplJ/shuUCHVAPEDcBZH8Wh8EqKYb9k7K6h
GsPtfrAUia9bEgAYAM+IShX9kkAFLghxfCjMjyUN08KS+LE8eL5YVng3oP3cFML4
rINYHg5pEMdf0PfYtEOwMVJxTZIM3fxAslWEWOKv7xBKCWMRwOokociJC17yMns2
cz/Ii3GFYmN1UrdQwEnOFpPWyUuuBQlx2mviL7NDneLcW0UACvrhWpn0E8jdR0iS
lAoFuPBTyyxUFOWD8aEHfMtZz1ySJ7SemTrGcPlchfueGUp0WXZZfoziBDjS8AYE
FOgDZROCBsItvD06vtb4NLSW5yBu3V9iy6BdZx8s2RzUwOX8ZdBuCrTkeIu1BRv+
BHl0AU3umfb9VgNoaeiqCGP8GKwz6A6ZQaRo/r6wqLj3CJD6P8ggQsIqV7LEPXAG
CgX4lC18ybrrX0nD7h4GMJn+NrsGfVHEi65n72gD1Eu2FUqNKiv37nX9uiozfJ36
BNuLKXp63doCHuzwhkf1nR5XUx640r5qb93RfB4iTH0hkV1PD4H785Z8GKmolNjz
b6eUl6kvffGkR1DCOD38q7mA9zQCok+5eXPDOjSxzAGgQeFKwRE7pNLFPBqgCbOq
vxVtkA4kdSR2+J14PYf02v1WfbxnMlt/rSyetmqXm+8Gzsz28MNIiu79GIuBQBUK
ur9GwyoF8DYfaU4UsDv+/DJeY6YMrXXc45UobAdYL+wkHfNBm6Y/O/IKuEmI0Png
3BknlA9KRWPxBhMWs3PyR1qTuEqDO0KhuCOSuOi+UE/kGhZq0/s5VHb2YMy1DWLh
17MIKIA7HRpDKN5Xd3qpnCdT/xixU8V8MICqhBbjFaewYBwfbZXODxSYY/xsr6Ut
vG+RILZvgzi1oJDixLu/jvqiRMPPIa4UgtLBdMYRltatwbfX3EujHZiPYBD/xWvQ
oKgBILA2TBxXpoKzXLTu11lL9mD3aQKFTqBQFZMpkTDsIKr6+CX9Y8q6w8QtRfu+
i92yKi37vXtkiAOnZBpM1YxBcWkrU6I8PBJU1NK0xwS8nGEOiIYaVeo3dk3qqH60
oI4Ss+j7baUpgFI040N46MRBiCopKMdyTEWumFRTXhc4ky92zqXdZr5TfEjX0nNC
2ZPdMkHzQB92bseP/fY60bTIdYmK052sTBi4Bt0MOw6TzhXJmitv/zfcQdjv/2Ms
PqScJs/ccHxFL6LWUKXDLd4rhEpbYLYJAuGu9WuuuuITbzvD0qotI6/wh/K/JmWB
g1Qu3kAGiCvSI9AqRpsuFWH2CmVarrnEvcSKbViPmJB98OIMVbOOWXjTMhRRW+sY
bgp2punwRKAhZQqFg9k0NFH2+oXlytIQmOLEsbByyVIFM7dc6Ct9zwq12ORSyIaE
GeyUnq7Pj7NkZczPLcaR1INeaYbPdyWtm1lNhSnXtlgRJOGzNijWoMqOAF3CUPmF
AvrYKlj6oBsOqbm+CNgAcHH1su5sTEl1nCH3jkQsrRI8R8hZLxe9da45gSKrSlk3
mXyBHmHHy7CdZaBEDnCHS8DrSqEgUIPA27jb307V6Milwg2D3it5p+S6kJlpVS7y
vtndeG9cJZ7be59+YJF33chJ3HZY9OxzfIW4OLRHkElZtsLHMMKxHI56cTm7u0Ek
Hj4WSBgRfIlFfE+ttXdOzgthYWPGUiPm3isSvCBm1yNpleKt+G1dFUqlxiHPWYBE
5hFDZ/OOMkLwBcqrdJtSofHrkjlCRcNdhPIMLl9liDijD+1b5bxXb81gVihtHOBp
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bxmvSUTcf9vOrlX0QWiaMs+3pa89rWVWZuPtDXf3nOsyKMeaf73RyEVUU4jVtre+
SwCf8OW5fGha5DNl6J1j/z29OL9ULHO5ohcRaPjKFW4PvBiVZWQBWs5yZ5KrYmMW
7icgTGLv3dGcZrJaHv2xCbZy6f6sWdrPsolQGXYH4gPnZOLq76DVYeUQW9MC6+PE
2kwVhLAULSWA+MRxbETnowm+7Bl441znWQR2mJMjqBYhKf/4J0Wv8+BVGuqYtT2A
F4ESvcYXNxEn9yL/MTZnem+KfwTZLlt5ch2ZdvyELsoV4MFm6pc+66Xnud2pKwbG
7qTlur1YVqTLiYXASSx8pg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8608 )
`pragma protect data_block
tHtcn1/zLNrE4Gl7om+xGd2ABvdeND7wEsJNGLpi3AdjyU20Cuqx5eFTailPzeg9
o6kL6OkTRr/nbAD+io9fGroIe8dEsUqbmLa4BDmZTkc9dbgxDW3URMdrDq3SoGSm
BZwxjLRlE/Zhpzv6yR1TtlMRA0ggxDI8KSl9XZhZ3vRIwmndTjI6r3E/8C2DcDtt
+pnyQ7xJtEI0mj7VXubk9DEYlpSTFWApa6jmCpziuZ/UpQdElsh/E8hscQd29XzW
TqyRHPrCP85SKpSN1tkVuhafgSLIytB8BL1Z994gdWXN7Cl6oCBeMQGQVqLL61cD
9Ag/efqCn0dICOn3j7tQ0hfY/m99rsgVCEltbdqMXO86UqAQ3TWxPmvERpMLgZY8
5sBb6A7+qtjMfb6Fp9eXaKjooeKDIn4fd+/neFf4TVVX8ePIS7syk5UjcEiaHwsb
Rg5R9bCbX/XBCI9Ip159rITXfFEAO3IVico8FamcfadNcNg1Q790VlBVjKFNa813
6JXN2bhvmuZ/Eht+DexIA1Vhh0Zd00+RMIKd8KaTGWd9b0I3HA237zxzYBMCB/1F
dMJwSWnfN5X+CuDkfUeUSfXh4mebVUX3U8pqvP2H8BAW3UpdeDJekUYdCoCnGn32
q6uPOhHkAC0FlsXksZzjjIMQkSysH5K+AQPHi3geKCHd6QGlAfBvMqOVE9E+w7Cv
/zO7CycszQXFFb8c10bsxtu08y21qUHOC2qnqqEozDF2Sri/4xGgOYmpO//7dpYL
bwl+zTN+7yAq52GwnI5VxBJ1m0AOr//5f1JBgTp1dJSjFVwqp/8LbXo58mhwKFMo
vD5TzjXei8B2pmU/joy7sqKwc8mCdjuJYcIrarnWXnIoA5cZmm0n2xqd2739w7D5
cqL4xyKomUbotuik5lcaAO/wxvdC1zcPKhRv+GIaGi3ilwL8EoOEGAnJKbHg5bhv
EZZLENRz8zh4vfSIfcoW1NCoa6NtWoyqFUaCfkj+SQTOTgmdeJ/L4lnZiF+Y81XG
D1momVZDgC/LTi7rLcW3RgGtsEGNHerxV6zswCCtECK34gtyBD0ZOfs5d6dTAaH+
WkKpW0iMagQ4Jyh0dZexaeGlDnlYm3Si4iynFnOOfmTaZGnpLTXg3bby7EvzFvzF
cy6Y5va4hLO8c5ZdwKhBm1gqPxOZEJAYUYJf8G8oFSzLGHP54h+MbNvsSVgBkFQG
PkY2qq5mcY1gPnNcfLDP84pMoCh1HeRtJRrGJlt8wy+1KBMxiOSlhPk7DD8P6Aqu
nyayBiwcg1DaZLZiEqXcznkNfUO7GOhOUBOeMdqSLZaK/PGZHDuCfepozF4ZGeP5
SGg6jvvhLQARblWmJCFr5ReUb0Ej8kFkf6fI738NG5xQMfgCdeAKq4+KisX1FU9a
dw3lPFnQn7e6LtfeXQ1yTjOZrOYdYslEBXRxeZBDj2Liu6n5ICNRTZOtbhnD7LVv
5ZTPzHBHwHYbOGUe4VlA7nrktlUM87K4Ptx+SwPlljZl2Hn987S+xJ6P2BIXR0U7
9DmyYhm8LA895tb4x8cIh4El7dlTtMcIKHUF8iX81cB5q92rrof1Zsmxn0p10JV9
JHPLxsmHsNETbNI5FID5B6ojMlTkGFra/EAhT7Tzjy4yww9nw4mS1mN3DDmxylUU
BU5oqjKV8iSdGf4OaD07QwOtqc/F/C9U0CVZn2UJI5T4cGC/H8BxrylDB8RlWt/e
xxXdXcBJkBoQ3shwZox8crZ8/djga6Iw4wFZqst/eF45Jagc6CtmEXG85weHwL8P
d9ahtTIzzR5DqIIi5sl86WbvOO+CvFm1p8kgpwvmE8yWYWaJ3UDjg5sK/jXnc9Xc
ZGq8tfP09ejfBPQk7CZk21EK9n0F9JZ6GBh8h1+nqCqgMllhCWMn1n+ms+kpUThH
4G6ip7AQohm5mus/M92E6nJtsMAwLXU5l59/K6EPM+MDhjDuYQCTJNrsZqJq3PV0
O8UXkkIQt5az2Q7MoFZcbKfDJ2Ig74t9VeHZHZthDLNK167OIILH1lfYR/HpSbby
3jF7VEt+RSHoCXxUvF4VC4w+prQ7+Jl7pdmyb+GLIAvUH+1jshmAWseOVcVOSoel
OscVXh8lvHXhyMBdh5ivaZTwisgsKz2PnMLdwa1XJ87IUCWaHYARM0D9uO1n6apV
UULeat40WKWCMMd+EK8tSv5Z2HSxvcpDNzOK3tn3b65CuiCoqktypLYqyeq5pBgQ
OB0ht3oQ8WYpCdFQKoVmSq5D5EcZTW+bxKfrvTK1ftiMUrM11KZcMLq76uHpzvxf
h4Hk0uQtrBosxE14RpEHdtzDYk2KsivBqW0qPib5t7blyqspFngDDtCx1LnA/Mtn
SHSeYCpWsjKVYVvdz8xlKQhaEPpnFyIjmquxuWnFkKkdyJbJf6XMSPySz8Nu6nHE
1cSBBU/33ugHQEYfq77Pkt4XZU1sYuRPouyoGkMZtmpOyRQ3BbKhN+okTMnP5UJb
fuxvTMGe4xnU0mIh644vkomXNxKwFm9AxGTG5ZIDbahTkcX8bGKMulbRvX/udtHb
ybb6iQaEiyRMGYKz1HuY2j4UtOIiZhN36d3Vfk/gAu1Up4NIUPTaYtL1GebMZM5M
V6uju7kfc4alg6p67sMm4a2NIcS6iAH4S8JDyGMvVlfkjoLV/H2QxKJOe92HGIX2
Gq8XXEbMLsvHyL7YWqts+wqQ4snQPGQK+rDPNRHKrnnV9ITsUXBj9UgVEbWjwJgw
bCY0p4UNEjClQoTW0DW6HIJpBylrlyCc8lTTeGMxhyxGYw5BHknvB3/bTGEL4skT
xNc8jxTzVr4rEFciHNkbP4o2kyTwvNBPiFYFGz6Msc+vJbYYR8JfpwaBBLkxIWlK
c/ARsrWwcV3PMwTFmR7v8dMwzJsFe2lLD1kh0MSbgXZHxY7c4eh22qOxk9ghGmOZ
xQe26c/SXIw4cNLO+vod3rlrLz9rnsccBMhoR9Xzsx+rknn6Woiplj+G8izg/esB
wnN/B+6iMnKlbEn4c7jdxBWOaYm51S0rvLbgxBeNXUr38VGTL0heXNJQltePFcae
CH0eN5iWdCZyVLsOd5kXo2HJ7eX1hOkw37wFe36ICk55raXs0RJWBHYHWdauJKW5
j/KMMO8PJ27jK/NU3KlKOfOEPsc5ni+C05B8cd5pFo79ph2T+pujz3PUjZ63FLht
K0H/Z0r0RAp2k6Fna0COFiTgpDkCbB8eRz5kwbhxevr9nP1RSM5Gl1+Kr9pejCzK
+DR3B9EB0ZyFBDt0MsIMKzmQN8G+E8ITQ91PJ+O4CxEesH+Pxns/GYA3s24q8s/c
cfzHm/5TBMYa2ww8EOhu1QBTMgwL4gI98BgIxRbs5QmKfQXDe0fafQyt/r+ddjrZ
gVJIT4aeEo7HN9WWJ+XtZ50iwKn62quZ2l5p5pIYOWxffTwU+Bb7peKxaxXDbvcY
CVGDJW97kPtXPKkt3wyI7q9xaDy/tVldXn1hMWFizvDQZ4aufnt6Xdo3+EiAJSKT
DicVB3DAFL0Ui1vm0FxSTzyKMH5QFugmmqQXAHxiAjKMlZ31x2ao/4hB2MzSOXDT
xA2suUVwTCDn7kkhfnqZe1X2/bEpHTSISlP1+tafRqoep07sCSK92hO/Op84+4zV
qqFY+QJ3+JDXGOg3cmiSkbBs1zwuhfRyCzSAEVE1uwuoZX6fsY4eESHVbK3d+aW2
ClM6u5r9vtpnz/rLfu6KrBAl1srDvynzh9p8+qZ959rmvfTmMNH8jHyxaAm4fRlO
6J7pOy+HzKA0AZtx6FlNl75IzFkzh3QMsmH6EZzLC9jWxBP12HTIqQ/lOQyT59VO
yA2BVrGBBEBF7RM3Bm553v1o6xF0t0p68zYp1FqM+3huWUSE99DoP9PwrDbBQo89
FVLhMddMdjQA2g+U1mOkFu0rNYugKT+zpxwdJ0kgvLU6ftknuF2ri3NpbVyUrbNG
1ucrj+86gCnIIDnkSVI9AAe7HevSawgdJxUIhICFAZO5htsnWNCXOs4vDfYR9e7X
HIuR1cBM0pHDFUfzQAVDwc6Bh/IrTVVLqp8+3qPZUPnF3BxYcGBmiQADw7kmZN8W
SsLzrNE6Io8A2MAue6LChBrRq29b6L7xGxtREX4TDKk+eCdWYwlc13B3Wc5dRPuN
9oIRZPHX2UELIKVIzYdVdL6MYcLQN+U2RtjueIECfAJNndTfGJLdGURcylETNNZz
kctrhbF45sTirxGdaN1ZaDpJp6K2qhFxcLmYpwQ/0xZ/Sv/lN9Zu/BWZrlbJwi7U
DPDDT8mnW1/A6/83FS40ssaZq3br9jSFQOQjsKxGl2sVZCSZ91uB3APmOK47SBFX
6lD9PzFeuZLeQFflyzAqf8hV+m9ei3qnboaCEGucodrPUibOrGzSrL5leOqjWOKR
wMg4XGi0FGhGUQIGtEFdZsqjHWxD1cneYs9BsUhVeji/JXUPp212ZlsutUpo4tOC
Hf3c36e7Ev4eNi3WxKqDoLeu4+0KA58GiLtCZD1R82RYO/kzrojdigbzrGSRJcfd
RXjPq7ZRWLBLja3D3gJWZWqleDPfgFc7ilXZBThHOlmND5ZI7mJxXW4JCETXZ/jD
sQToLRHKiCCRmxNPF0ZpIbh7l/WJLnSQptbUKT4NG2niPPB3bgqEOUBq0AqaElHU
FMbTtphGd/C/e1L0hDxvpIY8rDy/I6QK5nqZj3Q28hbIb7eE6wbox+peSznt3pGn
PVjrb5XYp2h4978eXmeE85xDGi/6CPYArEaok4HfyyzyZoh9hK4cqzQAOY9o3W9F
/+6Xbsq/9eWngUIz3oB86ogcAflPklBTlKq4CL3aDzzn+BcG6Fe7b7TYNTpCIq0i
aI5avGuHkrjV34eKxAsT8UCKOsou4F5JfvZWcEW4voM0jvCsHNNOqURVK0nQPxhC
QEZlpUpnUHtmuXreZgeocsk4U9byXC0vCBtDfqtwRWymvm1zCuAHq4No+RyYFzGL
bZfqLEMJYDdXqRSm7VZNKrSfnVaaGjBWANk2GI21K38dWyrw+WlWb2EKalQEx3Vz
tkbCkK54CLo7U8aAb8qZwPE9ghUI/OplOQhSs5agVsh19JVKd4WXI+40cZebmd+L
VVedTOQTQZgnRIRFcReaSvQsCdpVw2D9XEBlJFnWrS7harzMDKH+gnPezntugqd/
O9GkQFMh+SUwZKVZJmBESFA7D8UZbhYlQDeTOZimcxdxOpD3VoBEluQ26AfQLHpv
PEZsAWqyvqM56Pghlyn6CyPjyVfiCOD1qxxzdcnaofHBd1ZvLEWFBSQcQ1h9EnQe
vTKZu0fScHeuE6DLVU8LWD5jDbIcOuqApVNmGP4sEceXJHei9PIz3WQfyH27zpSr
EXPkr9OIdqLwkD2b7mVlAeN1CTbOYyb7PPaKFR6FKZBjRZNqAKluOkECYDm2yCEe
UPmBc9HAA49udakZ1Jr20Be102gOKtmMlIig28YJBeDUKY8qjxOdntB0KIGQtUcP
tU6QGrIqwnViP8pYP/kg8yXLksXOZQFbsFLzY0MLyc62aT07zjZ1RBLTO5eX8lpq
uwJzcPeDj4/o0glMtZJWVGVuxdkkQ3heU4w7ilxJeqBK8Sm4DjHPRFG7A5/5zb43
cwCCKFHLr9MovrkvNhdlXyy2etDFJt6yAzhflv3SaGduJ4KzTmarrIWln7urmhW9
aI/89mh3BzweRawgsJq1CXrSMDrAlvQm+cG0yD//1571PuUUWKGpqoBgLfvJgiB2
/VxEPU5FavyaY2wqfbRjwV0uQJwooUx7JAxsQbPJwiC+EfONmmHT0qedtmXGunJ+
Kpo9XZzi2y2pfCYJtqIHXbhmyJlCPZDNK0O9MrhnwqL97tFCbIl6IW/z7abM6ltD
gdnsu5N9RdHm4nfZEXZy2mYvkYX1QgLmFVXrBId2zZtIc84yDGnPHBEbsAVyBDpz
jY13Zn+b0C97N5obdYjyFDcYnfAlC5PRuR34lBox0sYbmtEkI+ylRPCufI3uTVom
2VZoQnIV6h2P8rU4jfo3CEp8R4qObFn/b+RDmcXFQGmHMeGT1vDoZIAF1qR4OUwI
zcN61Qxw2wwebKYWEHb1LdiK+H+58d8kKcxs70e9RL0/Oti5Zj8ETnXH19Z/KawR
U9/kw3vFQBXH0mddl/8Jt+MdVjwH+42hplc3E4nxp88MhO06ryqaQh3Z1krvnQJm
qRegaebqI581p91Fxx6/zGiVRq5BBPm3BheBx0Jz2Z4E1YzflN6Han2mtqv5X9CI
KarLZICM6EtIJkObt5U2hrcti6+uP3TTFurEyxRu0mQ4MySZk56EAJA+HvgYDr1n
UaTLTmU3IMqgK+2+ERs9kRH+/K6EoSs7Iw/ZiAuHhOjmhW/rM/hWRYUWJZFR4bNw
AGKJi+KjKfsTarfbncWbYGJgUoWD+PP8cidUKUUOvo2cE3g6KZYGYFInlhWiCRPo
CNu+rWBTINPMt6EZBDNXLMzhU5BxvXTDGtrRlAkS/ZX7SniHzinMnZFACIXz7QCP
DmSAT3Ae9WNECi3Wwxq+Z+x3kgrSoEUcKAS+IQt+4GqzMhxQ42/xvBfeJk4DiQlV
KqyMTn/rqVOSqe8JpjwuJdeXSaR+/kgZmbQVbb6fd+f5guMjhV48rrGyHa5VrTqG
OCN1+AcKC/9553dFCvi7ifoIsPYJQBsppR1bOZFF8ZmBK1pR+PFiNLTB53mUYR8k
eEk0g/6YHtl/xxSl6c+NbEY5chkvPCp8gw/SUcGRnZHo+8+ZRM6Gj6vci0G6Vg+/
8c8+GbERzOtUT4TnSVbMh5sesaodrol1FlFBGTLQespSZ2jdDJH1PAhUYOv4CtJ4
248y0DmJMUZgs9mD0Y7Ibw648il/ANm/aHJ81sDwpkrrpV1gb/BLD6jid421WcO9
cEyhnNSyY+Sg7+/bXiLKme3/6e1Qo+PDl+QQLiQ7SsoS+QgvRctJlRPlceyXhRPo
YILvHOeoKNvBJI8ntffwzfFjud7pzQJEr/dRQ849Wwc9m8ACiNLZJu258wQCyrwu
ds7+MIRpOOd7a9NozkVhz6C7CNyxE/EPp9pMyXHv+Q/TFJ5l8j68B5qq5hBrItGp
RXIJZZsEiZwW/+5MUaqP3VGC2vDDpkKqwfWqJSBLURUHsn/fWe0fJ6kIU3dUtWHu
3NPAWM0vVIYa9t+nWjU2RSo4Zsu0wfrCCbcsn1UqKrbdFQlvU/Quih5n1/CKzLs8
hy94zFpwvWb7GPLAw97O/Fyq3YRZtk+BVFfAAGFe7feyUyOgV7yraADUilSfyF+Y
mtEOf3Y2Eeg0mATaZMsQzP/1grABGF9uy0FJ93zn1hQu6eEqVzU3al3XxP7kqnOc
7sL2gsMWcpUPYFwmJLit65X9mwHm1tbcYv81FuziMhICXiFJKK0lQxsvf1gaaI8r
qHzc1ev39DcWof8ALFTqrFfW94aWP+1knvM/VBEfjVhYbwxMuCCHES0qCefmpVy5
WSFxExF4GPmzCBB739csoxs+byYyruVnNJqF93QFLa/Gmv7F2cG1TMaiApWAz932
MuelMaUWeQwmxe5U/jRX52EVfz/x85nF38l8sBg07De3im2MNjSdJE91CJjnfZRE
b6yuk51ObSFmT7p038OXUofGeONTyah3FtYOibPRzz19H+WBGWO1/AWQFJ4WcRNh
TtBaAAEzYXx5tc5CiM13CHqCLbUlApFAfrCBw0rT1NxHKfwkrpvteUJ9GjBUbt+n
Oy+W/MSck17gtCWQDVHbzvBM33j+F5Slo/QdQ6LrL2xLb/0Lp7JGRhBTK5Xu2r+9
qNEH7Yj9ZT1VgWKhlG3oFmrMkrQaRA5vYMCV2ndL2ei6gQtDYZm6REkB4cctRC8G
H3Y64Se+HFr0f+qW6K/XVJDvkAtdvIdwMZGCs/kQ2YjurlSFctVYrfLSzHhaX48z
oZjiHMt/lLg0LVuASt9v/OONnkKz9JFY2sDOfYM+1VMKg2lBrLZHjIkQZoeDqXIo
3luUdcZcWNibhqgAoSc3LQyM6XHYi7B8YNlTtmuZwk1Dmfkas+tyZAeEVmu3RoJC
8g1a7SzJK47tP7aaj8g7pbRVmKm9t//8rptcAtGe0CQjVJPVsIROdFe+fffDyLXe
cvqAhJ+n7MRV2QULzEeNWSCzR6dEH79oE4R6LsLV9W6GmSzqcvAZEQEyj6kXDXWB
xPYa7IDpT5h3KBjXU+Kt7FSDQU2/DCt4rsDh9wKpwOEKOR6OlxQH3DEVtdabo7ao
DyLFcqtat1YELbrNBBBt4B/M4THFbbdgWfULxEX4ZQAH8ZMY66Y0NNsemoVXXm2a
wrCN7UImRqv7HL/ecineXzz+vkgA9qmZMi6p8ozqzotr4NbdAxyyVBwYehxIWq0L
DzcgHFZOar1vk0rVMubUtTbq4HzZgJ8PfhTuvSqqyOLbmSLnVMoYfJdbi6u0P0+I
PobVcsyJFrlUA08mUf1nWKSt9d+RmCaxdtxBM2HKEdeTM8pwm+CZzQhhER3TFdv1
Pn4f77uXb6rSxxZvc34iR78vJzLAnQz/iAq0ecfbbJ19ScSJDQcKwguXi9JDilXH
AQ4LtWZosc/tpAFq7Dmlhwzl5IleELJSCCMD70pk29RY3Sq62pQi1Dp3CTX1gAEd
EE076nozKOMWayliE8tr4vHgU8lVqCHGq+KZydR+1seJdl4lfczoo159WKSIG160
GRmFwmrvfIMJGnx8gXguqcPixXmAM+BsF61bpLDHmodkrRlm9iU2ZfR6OBv77Pzd
cfS4sKRZ2zBn2igcwyGR8ZlDN8Av+VATJe1VRWOnbAwR4BihoYJEdyp7UzAXMG4d
Kd4gY6g6Sj/vfqGvwrw2XMRY0fhNqN3RX8Wi7TemJrKdZm0aPPrSjzqGevreSDp+
/70swPsKbN9jRCRhMNALJcMCJ0SECqKV2lvmpLHTuY6oxX15UDLobsATPdPZkhrs
aAO0YYZFL3lBCCYDzUfg9qn1MTOkIcTNNEpnlnl0MRN7PZJUe4iwXYdP0M2yAh5J
0YvFDwB5QsBu0mPUUZ8JuuESyKEpdKjHlreHJN3bPC5wv9Xb+Mljv+0E+22UkoiN
wah20hK4Gi6LewvdCZgje7ssCkSP3tOb9jXEANG7PrVzLFPPGbE/yWYSeUzFevVi
O6ttTyQg0c7XB1dNcCo2yxU62bl7jIuMpL2p0bmenXnhrtF9XfotBChLC4m2tHxO
x9oSprDvnS6sn6CQZjZVrbhD9ipkj/nxV9B/iXS32LDB3jK+8hpv5eQl8MbSVK2j
ReONxychbeUfWPKsFYjHS78HW/+Qha9c36QASJ7HNrhgKW5uzO1tV8SLe6LsNoUA
chpghvgkeSx2kna/VR3Xoc1nvpC9KBDpE9oAuOHfaQtZ9zbGT8DBwc3T46XqjTHB
FyyIE+CXQjdxe/QHhYxAkdIzEgUZPt3IocbXkEp6Xn3YB2Mrqbw54tAPlOPP0C1V
BB9v8MMv0CiWhBtrdPuTqEABq3u8a7c1KXhZFspGzlROkQomnAlhQVb+SpW/EyPs
sEGg2EYnboDLQL3JknlcDAc9kEVVc7pp0KMQANin3nOj49KpvgABIFZreQ+6nIed
jscR98H8DO35LBwPq19wtfN22093P0uNObQY4lqVe96PpFm3mcvjKPPqz0fZpIzr
LQvo+wZFyGZqsFkLYSxLheCj3wabRhRrfBpHUZrWERG7tamUDALyyGgVvbdHBzly
fb4wLapORsn+tuwPcjPJG6DSnE1lvlL8jMUHTAnb87MqoP+H9iYep7w5n1rpMNxp
C+uAMbc40VeOJ8ZZeMW1INMbCDQEThRigXLsxEwIm1sKxcY/guQdn8QePmUSupZh
p5kXf2iMUPgMxzrpKCjJlMkJy+chGbnYck1sUTlW/nFdajdR3+cKqJxrEDKWcUZF
UI1mqqOcGUjWCbGOlmOlTPB/ENqww9lnxo5icOAMfS01WUoiaXcOU3bpAN7Dn2IH
O+etV6cvjN9PHHoReHi9oGVOdlpZvNM48q8Y7mHAKJAx0RZ3BojW8/PxYZhmhSDN
ahcQ3Fijg+yxHyfCOs6qNATG9YQoO4c8nspo4Xwz1C3FEe0ewel57BKBMIvVi3WC
GQ2JE/dqffuRpLz5CuZ8pD/T8k21nX1Gdla+hwuKz1jCYkrwGVvRToAH2VaC2URy
MpntLg+g5BngThKhf9CITj41lSiR2e0cfNBqGm6YtC5BjWoxZOhnHlpxaJSbCg/H
lwdy+fQePJaW7+NcjBSL5NxSCLt78i2leOn01NJKszb4Ok4V+nQwfYMYPE1B4ipx
n8+uZWPfes0UBsrjZ3EO4pTJ+woVAFODpwnNLrFodLQdmnNpBV4hYca1y2Q+ftXZ
XFLxKpx+Dp2TbGYr0jWJZs/Mgs9g0b0iL25Vd+7VY8HceWZOf7knu+lZho57t8t1
1Op0SRDawjH8J54qGHgR2Vluixs3cUczrUae4bbe1KzvxANKmqXdwZexbdRNz/3J
KaKMjw/ud/4APU9dxemQBuTl99YrF5mMZFmX0PdeqowqQ3inxGmiOixNKt6FL5yz
SQ6QwES+/to5rAzq62nZELRRmqkoaSeQY4ekhIUa104uIRsaUVQePxqsTE27yeep
0MtIikv8SnBfuZyjMClrcOVFYWaK6Ur/GMFbijY/RZ34z63lk9UEq6xKA7NsxaxT
cEFBJTIDbRzbTOy1s2ZlQ5/4ahvYVkviS2G5gAfA7tYGXbtET+mZMQdVLIX24NUi
TgnoWhA4p4TyaZGZ9d4RtL7YbTlnPQjyFPzD2cL+hKWmJrPLkZo1cF6DYahwKtl9
6cp1tlBZA4AkFHJ18goOa4HdksWPMZZmpgGYltFX1/+0EuFRA+pyuXsSDTC5m/5b
uzzZn7HVWRrWHhJ4Of4Sv9fx7oPPxCDazz7zPowS4IFDh92TE+xP9+GgG/Izt8k/
KydWnHQwMQ5FT5FBpQ/LgbK769nhNdhskL1e7jCDWLM2Xu4abxmysmzhqhbTYh8l
GCcX1vgkiupU9zJLZHgI0MnFLK+yAAwzffyZAgmY3cTgL42UVET2Fg89CiYk57iR
POGDbzWKJS8h5xOUjWIZIybuCVRHC2Bn7U56ymzFJZhbOxRFxprYq/daQB6ez2KU
Ip37LNHZFXUh5FwRrIczGjIyS8YyyczrWvX/Z3T2PO6Drn989EFsirdxV2HupyRV
RE92J2IU3RbHgNfYwX7F+2ySZSO3PNVhlWVhKS3kpPfM48bBzw/cfbP7rXcbBxhk
ZPH7HeJCz85BmtSG9Ixj9a87zomvmcYLh14LQO987bp96aiziEQEM6y7Czkyw48V
wJTZ2AZba1lTEjqmCblJilQBE/ccLLmCOkQJE+OINdE4vw6+7frEaNtAMRYZrXis
pvGlhnEQzPBxtopqlDqDp5DqffuEGM+a+yAJwsq+veI92Vi5FM9pRm3nx7bNTpsV
BwlG/ynNrRdmHhfwtec9WQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
e4kH9ekt5lZWleHbD+diYzA7+breQAgrLuTv3fM476XhCCxI3+RC10e4jHRKuQcO
AtqkmDa/NCo2mUNoDYWMeUHOT4LrsyOSLL45UxBkBMf2JgNEjpcUSK/hm/Pf2gZG
P37YgpQ9pecYnMEUi+T5RQLrOVNBIIDKb/yQkHYuTBNuDYdrRZmwzHbE5dJu1cTX
7mt7PfhcMp/OdR9zZDrAjLt1c/7251u9577Vu6re2je9l7NGiCHJSlw9/bEkEuOt
5TmH8Sx7Uj5+4Lnzb3SIzhqoBRpl0cpVm37F3c/8RgDtQjXls+aVUA4kqUlbwj8A
mDUkkaX1TprcLkofwRkNHg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 28736 )
`pragma protect data_block
S/BE0xRF8cZqgblCw9uYA0yLKSsFvNtOr0O8yKKbTouzlP4zAirK98cMyfecn0lj
9EfGJEfUyuEGeJni5Ja+jC5KGhaOJV8v3vWTKYryd4mK+P3q7QXag3h9EyNvvic9
YvTmXqi//uwVz6sBGovPqZPZDGK0mvp6p6yg/17jOqwz7mQ8IBFb3oxLp8WtOZQ4
WzungX3m8rdKuogosH8yCmAv8tlFQJw1JjKhTAegUoe/R6SVHbGbuzAGFLbbxG1W
Fln9TOcmO7ciZRfRPmXDfLyOywOgYRNP8yvtoNiE+Znh4h4MFP0QAikb9uomLhsA
RllTAKbHS8DPNsZxgTyNYEtgZ47twFcIGeAUVo3Pk1C1j8MEJS6vWRAUDEYXUUQR
2A4bRrK7C83ZMygevjz7tWJwPNScM+yoB5kYg535FlwQd1Oxi8XxdmWAH5RhqCjA
YAWLq69NEfZNGy6KvUgytFFZvIN3h3mVd7hl1CeRivYnL8pP2l/OBcKSAwyxqYsc
K2jfJBCUAURxJEERZ/IjX5a1eurHESB54iWht0Mn+GHK1+co0+ABr+/qv37wX/VN
8rXLBwBYVdpsHXQ/KgscrR7MvAyNufNYD2CkymYRMM057TqLhB2ge+OnkVM3gbRq
OVnzhB4sjgjsBv/UOxoDvDqBox6vaR6QQmtQZNe65n+O/LVThvL5Xc+3SRi8wc74
4vBl4EeyelTc1Y8j+Et+vGgUmR0PrjeGhOgVacx/LKaPMgE9C5J+nR1X8dYlOUD2
n0m+rEgqPvb+HBiafwqLhkC8COt/2KTREOQJs46LS2doX9tj/05K3TyavYZsvn5t
QOGRBKH0LS74fyuT9e9arKpTOLQNoTYMsYof7i0wFsa81O3yb6qPwbpzKoz+faOD
T62prkhB3KX22wRYgLhK3rnRC3EbTJ073pS5wyl5WY5atykFLs7tiwnUjdzNNo+b
HGEWGgL5Vpu0UypzpxG+h0zDCbnhP8tZNJxNptiMLq8yMvoQnYQGex8dmk38x3oR
vR+cjCF15aUIcskhGLbozsTxOaTky6SHs+hLzTz2AM5BXKC4RbTp/7AxI6AQFm9M
6BpoKVfb5Ao/tBpuYBrM0NWxdfxn9lHizVIGWQ5PldUb2rureMrEhTnEmusLXkHO
WULhxny4ZJIPoP3J2hvjlgO/+ADPuS5lJzxwL9Vo7H/zkSEUQrsreMVByT1nB5rA
VK5/Y93tCc7kavvVn3u85UaP2RQ29SVWjBlRJOnqXMqT/pvtyYAVOi5QtKdCscUz
xYTSG5Qfn/V5xd0YwMZ4pWJ0R7yF+sxQXltOsOOCFiVNFF3blpnXWBI+Hinqj91W
3idiRxRYK5W3PyuEA1Zpw4ma4MxdBNOGObbaW8UImpKmx8CvM4qaOsxjklYZkVU2
Clo1Y2FT3U0rpYE/gu299Rh/X1lpO8KArGMZbaA3XYlfY7tXtKCma3WF3NM9VBnJ
2ndC5OFrfJrwuUTit0yDf4KeiLfJFNmnd9r2GMFM995XA+ciYPcotzM871i+waIv
CmT8cgJkt7LHRMv+tEmcIYh2fkhS79IqKWQkUFSJq3QRdbASuyENBbyRZ8BHY1qY
x4QM8OzXe2MdM6GzqqwuEaINlgYwWMbp+kVSGFWu9/7txZPUF/5Ub6674dlThOEf
5gegr5sB2gSdIxFEvXaPVpVinJ5UONWYPA3YBRlT2F4U6rv+0qH2l6m5WvlpcXz3
YhOlNAXfPYULse4FxdNXFT2+/gQ8ItR0zHbngc177HFST/UyO98Mcs/pcBGqC9fT
EYrkyUnbA9+F48pMlgX+uQ++2joNPkiEBjiXFTqLWwz+9WUGj4Cz1VVKzQi5qde8
eDvRt76OUVrKlw9D7/As3UH90KNs2GiY1Fg6W3Ssxa8lXNgezrFouDXNI1p4FYth
Yha1MFoH3bFa1ec/i/513zNJlZidvzHTjj6ae0huyRVw2LbHHAeiYjxZB1iGtMlf
hDN1K1x8rYeIANvRVqHL4kWlptNSx8pf7HzEEyBhJVs+dU3Gsl4casq61/T5Oh70
jbnFMQdfVWVRZS+GOY8EW1wewYLpFYl2Mhg93SJCfzIMAcn48c3n92iBHNbEyqkY
zWfunXXtrRATlfnfzfjnUPLFfNd2bR6egiYKY70vEwzQJZmhuJPwTS78IE89ugQA
qF1QtkHGnZCxuD3d8zhesLz2cN52HWM7nO2/5kBjEZXJ0nlMQmb5+k9j9mgZpmJM
O9NM9qRhAOkfBxvxuLkV/84OldUi1CvU4ci7QjBjAK+XKHNCIb7ViTrRAaeV5q9Z
05pT3WmVYo/ON+u2Fkh2+Uwp4TfIeiqspByKnZiAwy1Mr4HaYAj5MV7zU9rJoVR0
3CJZ2SIloAbkP3TZfPUHvmAR31yVY4qDo4J8VOZTuqPc1I3M3ijyowkaAPMUfQV4
1+LGfxDc7BoAa5uNI2J8PuVSG62kZOTkkmWcJqM6GrNL2l1ViVp9vUnUxhyfPH9L
XR+Fi9uUM4ihjzKKcOJ+7Y0gZTT4Ypfdzk1QiMdwo4DRIovbHEAoOrb0g2T1RKzg
C9I/qQqmNtXNOhKnnmDYnTSAnbDLD/VDyuEr7OKKIB1hEVGe9tWN32fuHpPJn9fY
BN9+u3UpHOiaEvn+p1JzK/YqddfE1pMKrhs7K/SbqQkjYPZGDPJPL1nhHHrjCLND
TFChS0zd6WPKSHAjg8/9P3wcFodqDJ2grxuOesvyYvbaLxGeFVtBm4X2KaiDoDTT
yi8LBTFVCXEMFvnY1B4lGDbIvCspQec83oMJ2SKgPsJO+od8qgnmMx0PjlOcALfv
e8dfoV0SDLMNYfaIjwx1A0tBOny9tEHajQnv7U4PaDJAj6gI3Ke1GAPsHZvLqMoR
deXV3PgsACBH7Ma5BuWF9pQiXXqQEkc6+nknIGVk72QwMTWiDYt2kZenG4kFxoc8
8ho9u9vXjy3iXp1G2/k6ph3pKFrk+L4jG535DIJP31VEwOD+cOxV2rTT+pbpjnRW
NRy8o/yl6cPVCpmQRuwHbPdfkwdl32szi/PyTPu5ikf50zb4RIpUnLfUNsFCf9JQ
R0/9ls9JwXFqpZLjlzFYnLltPKb4rBYy+xCRq+xEgynzt/XnG67Ts9eDlXHJFxjZ
V7oT6Az9hDt0HOG+8kch1tN5lwYEjQuFzDR/05XiH57NoG1q7h4YBTaKg2+rcddn
bF29zmTKEYeFLbXzI0nuFYD2Ng86td6PeIlNxwFDvpOJuH0MH90pdN3XehtkwGm5
9EU5HBti6hpTPfjtvBZNemjj7ka0aVDvjBPNibG37DuLRoDD10IOOKusEZ/wEGle
Cq3BsF73GsT17iuUmwx0P3pTIb7JUtwZxFWypAlviLahAiJO7pyzwewgAsFiNPKW
a/ACa9ha/PjWOfzykfFJ7ZJ9rQJjSzJEPPRs8o+GbV4O00Hzvq1sTsHDK/6l/3GL
4xb7wd5Ls6xX3BOfdy6dYsf+fuy/EIdiZ4ExaaApXxBoAGXptgcy9wrQa9aUTBDk
lQDhHBMDLT4TiTa7udk99oyScVAlortoZQKjH+TJRH6cnBPQehQDgdLq6wlwaf8v
uo7tpHUCe/pL/gq8wqINDuR2FRyzmTdDrVY1y5eHWyxB34Sv8ICubwT6HG/1BtfF
H2O+9PGI4QsXJGLR2xbAlloF/tBMoG53FM4YX6rmu0UeIRa1970sIQMfkjDBzlpv
sIsudbaYDOOvZ+DcOgO98W1ppcJgw1SNGhaEVmSkKquicR4JQhHOh1n9swgCpvYe
xQBlRIm/lEL790mNlfMZc/H6Kz8Du7rxfJTUbfXfTJZ4B+j87cIUKKX740TK1DL3
MDDu9oQM7intfvAzJLYG1yImafH7k6tHCWGc00gz+tNN2n/zKcoCVETu3Uh2M98E
FIZcoKsurGHTgXR4QohVgoMihl5p6nsUvwpv4c361pT4oysI4jT7C5SEKOIJNv7X
15aZzXwHeazsiOYxzv9MpkLnAgMFa2lL2Ooxt3wqYtK2teWVjpOTsdxoKF0ioCUh
9+pTM5I5LEFRiX9JIJwFA3yPMb7A51HMQ5e0WX0WHXIbNxEkEbHrkVj3bafJ9h2s
v8i4wd25QM0/O3JUJKMOq1OAJ7cMB9+mVUFk91D/SoZDIhY0zwzVXX8vWWp705sA
m7JGjt1hnkTCssAlFSRZEAt+qGxlyThlyJ01Ydo7pSDvICtq0d/fG1MLidveJ0nB
DxlYwBvsICWg60FfRITiLUVSbrmL0zzMQHCqS4apyiSUOFbPCZt3vUm1nAklofYW
VoAfupspsoPPEbk+EokU5N128n6Z5HSILmhJth0o9vTCPxXN+QpbOiq37aDn1tP7
yxrzxafS3H480TpkaF3MKiI1rcRQ/Up4seXN7U7h32531a4HBVOPOV9MbJHD6rOH
La/TseE64vxuCTLxeam04jHZh+aAPrpvdEzDvk3qhAF1+xJKiji6Yp72J5OZpSGP
LKO8V9h0hfV1ZjnJU6xQVbqyqbhQA+v50m/mrAS7QLj6CHtllcxyhQAdqpK4UqbS
WyfEfDknsrZ/enj8SQmfttQsDL4HxfmqHLjM4XoiWjBr0RiV6enDg8G0Sa6Jr6Fr
PvdbrNeQHz4ok1jDijlS97wLt/awtswZGSeMiwOWO6Azt1nqPkz2EvNNiG7NbsCV
+3cwAissTJdwgjynxzK7+qIKFSQ+XeA2zkEzkCFCGtqKcXhwnaAkoxxU2TFWyTCO
ggzdSUkfPJ/WdAJyvXGxVsMW6T5KeOV7LVQ5DDHrP+GNZhew6ZgX7UyzewuXygEE
Zz9MECH4+Iav9Naab1xoMROtYuXA2NpvW1tnboh9aUmahVpekR0cOAZo+0ZWeixp
Z9byUkul2zYhhhJvHqLNLP11sCiJw9ta4GgY/DgnkLZMH/WbaIJ80wpklav/nvpW
5k4XcAUB0d/s3Jh6z3iLT1ucB3ou8p5jRg2xpNtuzAI/4eJxXIf9x71AQSqu3jsb
pwuYy2/lzFbl6k47JuAMP50KnXUyjU8O7RrJpQ8UNJ7uT2JxwADP5VcNIi4PBtUZ
F2iS3X75l9de8rePz7mbwEFxP4I0gSTsfoX1RFXpF/VhhWqjdhQwMeFjNbBrn7LF
IRdR2gcY3JEQw2Mt60qWFI5ssG7jz8zUYcGXuDwS3tnlkUqeXK+/+owB+Zrb6iJw
Ha18mdCMMYkye+jOYSAKu8E5WYpijBoJiCdBLsz+X4LE56jOb4rUuxRPtXKae76E
p1PDixxDA+Y6qKuPJniV21+YKNrdbQEJVW91bMgmq36LqQhtkjMEAnZRei6teXBC
eUME3opPE8xcBI6GqywTJrrhDUGr1a+x/F6M3yF6sAgTbNbXu77c4c2+67O8RMCh
/71MhuzK7rTR49bBG+rk4TKrdyEA9OqSR4HBLt3MnVL1TY+jM4XiBsQqzUuIGmVm
jYR12xU9t3STA/EFl+bUJWkClzboiWxNRJR9W+L+4LYXeFLrR63Y02FHT/X53qPS
Ez6qYpLyCpGdAr/Gyi7pCtjpWoHfTbxVwcYDEGa703tU7wMTtG1lxrdiAuwlHNH7
hLb6nM6HkCUEJuuXMsOStwRs2+URIKWVRyDWhQU69YKyxCy9HYORBYcvedcJ49zj
wD6gr1Tpqff50rd1P3lFq8gTpx2Qv89aZG1C3MKXOi+ZGdqOX/3wTbIpoSK4g29e
Lhr23OSwwNjy6GBCrIVF4p2pXk5wIPZ1ZeOMp4rS8uWdI6vYhZSbMVT/akrS//Rt
cvWI7XsdTLyYD4svbHMu7zlkkJCUJNE7zK73yVZMbY8/0vmnyY7L+1lcjwUtFK6w
zx0NJ3Sy5M+DijiN2IE2XUcba/QTrY/gDDML4oRJbTWhHV31v+paYoTS3YYu1PmB
Nfz55DHJA2kAL6gtNJ2ZAld9qBPm7t+fvSkaqloqANsuoUKvYG+CZiQkILGzrUCq
ej2F4/3bmBwuFzQ4w98EXJn8r3NzxbdTH1vJpFs9mYaoH2dhDKNmQIOWCLlM7kmB
d9RXrTiCCJkznbHUafmvKd+FsuOmFgXe8o1FOhqRY/rSHNuvwYReZT3Dylpq4rtj
z5PAUduLr3yVsZVTS2TAGdoLPNfP+300epW140LjC4vRv+tTJnu9bAVW0ySE5JcG
/ynyQVUDkw2T8u+UOSE3FL8dSgXzUUQrP5s4I0jptus1zZrz4fr7JNY1qg71D03F
qvseY+SJY0fPJ3eykwxq4HSBM2KoFtMN23M1D5OzQyUjH4W5AywrYrQ7frHIlZY9
31XcZzc+SmbOJW4k8Mdf8R8J8c4FAs+1mFkesv+idbCKr7I3RrFvBphg66KuFrrH
TE7wdZ1t4oLsdnmO/mMWspMUgOPs39Tjv0Jnlwj/PfT/U4kg96dwuBfkkDDYVQ6e
NERPwxz3oWoNUYPxPoBFy62beh0cp4N3J1nSchzDDN5zCftRd4dAR+nLu9vOyE1E
ykl2Qd26XVjjKd14AfiXbTmu05ETocJphKqjqLDnzhr/EXNf/ZBoK2xU0PNESL9c
gOVRDeqyzcNctmQ3vBSVRj7M4S/pQSyVuT9/nm+SyxVZXHcmRHJA7zhAXUkge/te
Cln32ifexmlM8vUIjy+ib6zKCX7xGUnLCmgrhfsRLxvpqXPlJlOQWGN+EPiJDBJr
Tygfe97OQrRXelb5mBQwg18WaNXPV0WRCSmI3xeGL7U57NLL5VYVNGLyiicCKgzT
G6DuXK9A/Ret+cVqCKBA52hLtaWC+3LK7KRlDJekibOgXA+g3eSQ8Obz/tLxVbru
NNT8A0Ek1a5dh151Ov6/JyhxGHuf2M2yI7mlmUXFNT7WDLl4dpN/nefIs26EU517
IMCyuFf3/32qaBi1am0gh9So+lPpbKLo2oddtkbTB814F7PMT8rfr9ZiTTc6z6q7
UTnTxENJNxOfOjs3viEcmPmqNj41fMdvkZtv9gV21HG6L807x5402XLEKTwPMPeu
NPprCGzymRHMjrXcoaeNoqjVSyVBMRJMQY6lSSRzqr/I+SJYBMDc4G/wAbC1bmTm
eSIskyPlubq6uuBanPkLx13q3x+kEXfvbMzlcnrnmkQVAWzUM5bGawvEmnLLbDlF
zij8O9ZGhlspjAQKa9/EUgV4TB8/kHOuFtX6qibiMEOJYviWe/JPsu3ovXs7POnW
J93/k8DdkoD8Zk3uCnaFDA1MIR2fbQcP/LC1OMb2z1VJwHpwCOXLY/uYo3JikQ2b
lKc/J8PNBiExp0U+Bz4pVwX1MD/e7Y+x+xZo9zwAO+HM3C86W+bRyIMq4a4Hn6fZ
edGRYEcLLqwdATngPm2n5EM8RyyANiKk4MJgBf+GusG/9BHKOBlWQJ8p2nn7tzBQ
teoWwjQxgFpGi324YVbycV4O+onhSYqoh5DxLdQg6WHErYyawM2HCZmMzylcHZkK
j3CZ+Ztj19laEKQLjNW1Rq2fpF7oKNVPiCbFddv4LyUUnJGZoQSq/Q3iu+DmMvE2
Vz38i+lE4lx6SXLaatVkoafQdWi+5OoInyt+bpRHKFh+BeytIJzvBiadLtct6vrX
q2etpmcEIyzvQs/vx9nKkMVJwYq6LWNWEsNGAK5BH7bKuzpikel/1abeCsjGTRAc
vvW054VWcjv5VeE0ylC7qdRmUTMKrRVJKMJ8/C4tvrZCwlSN40PoxNcX5xhjMJ4t
xy5+Ss38hv6V4NaLGlmbnC3TNP7gBLJFgV8PqYYeLWKaDRRdJqnHPuhmnZODo+en
63bU5XGkPL9A/boe23wtAiwOs23LAKiUOQ6B2NmiE+KsYmy/l1XcaCqUKhs77vhj
FIejQwrMDzJDPlrnF3BRcy7ZfHHqr2rjDBrac59Qw5ntkK9coWIAN+0TZhikf8BD
xM7/KmES7ks+L+NVJuIeFeUnqLaGmdDrX4MQ1qV0N1vTHurYt8MZxMiM+v0zo0OX
EF3VE5rnUS4nZ4BL5wLDvieqhEYOHOdw3BX3RcmX71HsU0cVUfdubzY3mUs6SYAi
UfiFJExW4g2SP8leYVaDIEDVzYeoNRIkCY3G9KPHzCSUoh10w0mCccS850k2Ptww
Qu994B4dm+H6ZL8IuSut0VGir35FEqOY08QkwYoiGiWSKFvwtWJLcNy4Z6HE8fjm
TFq+j1Xt5Ws+epc005mMmjd/gdWxMj60kYJE1ofUdHAsM/AC+Ut187I7cTOlUHKC
JfJCkocTmLTcpoCqlX6gk4x20rjuPePro5pydaYP3aYjez9hdtXZI8NwaFIZWzDG
Y/GsKWAH66aqS7hq0iNJyHySOEY0ZENATQ2y+62Acu1DgbXzwKOhNNvF0OtuPedk
OgNu5/J0ExFkuH4NpWkmSATt/3aF7IKaKbdS32hphhJeQBruzcc8PbkwvW1c9UCG
V7FKfOTqM5oky2vb/QdiezVY1uwvpAAnrUFYysU2PubvgDVGzmHnJgjUuOytKOL8
EH1zI1C3G79cehdxG6dAZdSQ0nGnxq8/kY/Zj94qNgD4GC4mw+ZoOEVO7TD+ciZl
AG3nIUM/xjnLjSgyTZ59GaVF7LWfxUE55CzhORrjpgNItu0jWjG9zm5w4Y2iryVN
PD3pA1JnTVihH0rp95NPTxV72SGIZrmWU/bWYrs7d5V+88ApHOM85gr/WrPjUX3k
l2axdEPechP/KuhqlnytR3DCsdyLWVuVX8aAqso2LVNmfhdOCuHxEKj5BiIXhOkm
WiwPVnIBNfjjwNSy2GJwkS8Nk2rsbkm1wkEFvFylQ1r7f+PIrTBDJojYNHV1qpKv
pwhu7u+os2tDSO68sD6zaIshXOcawH90aH2Ukn5OyX8HCORshnxkpiyJp26u/6nB
i9L+iw/fqt5Y9ZQ1o1HGD10JjMvCcr6oKiAkjFg034Ri4GoCHqcccQTC9jrW/rrm
4IyIImKw3ct1cNjbaVarX+7lDmSMzSD+FycE4h+2XhwcO4OOao5Ud7pWeU5oxtK+
4XoBKXdoCuvKXczvtD+L006u1dPuuGINqATniHqNUOZWWsh31ryRqRW9CirHN2U8
eApDwODHZAMF+srso1TqpOft2lHREjhD1nEclJhU3cSNgXCPFiqGsCCf9i8r/Bxt
vp447Pd91jmJibvC0E0lT36v1bRNyU68ilwYFgkXY5S4faw4QfX4q6r3LfdxD1Ma
kcQ5eJ0VOdJFvEuKAzb5uKOs1BcrgCc4x6a8nyEGGr165FNI+4//QkkObsBqWV0O
BypHo+QpT3A+AblHYreR9Zf1/tMXibRy4paVaq0wM+A2uVxQapVgYiKM+Nhrn9MV
IRwcZiz5lWuLUfbe5mY5bjcwTesu9eLMtiNdZaLt5xcIs6sk/YrkidmXv5VDXY42
F+NGDJiS9zMkvG76x+MVfEOV02uJ/Ql96DS3j8MkqP96+AmGWpSSKeXcidUrBePr
mRoC23BzPbhFHPLgemHB3crevrYjI5PQxT2dHEY+r91yTDOKahY2iE9+qQjUcN/3
FbwC3iARyICq3cQ2POHq/8AhbpvBA0suz5GbOunKpw5Fc1o5BZ+79Aza9NT4ok5b
GYbAF3PJ2fjPxUC35IGqtFgRVgLE2YIWqhrqzSE2p+dpXJ8G7+L1HtgvFOY01VI7
sJpngZPoQEukl8Qiq9lH7+W6u1y8+BICtMSiuhK4OPzL7y5bGUApEIqSZFciN8rD
UWjPv/H8xyOyrVJqxIziHpkPZaoU7ktHP4moDaVSBeL9X443v8nT+21ZOUzEPFT9
vKa2wYfYfyixBx3w5miBLaYWkc4z9KApuyPx31aMI21btaIlUFmF4Zce2prEMX7/
COQcZCRO05oz3rQalxfASd7kzPMGZnNMHYjMnzteiKlXnRlo1P2/3ofAQfOe40b9
I6pk2cRKejjWIto0SipufbckYQdhlFnALChDOsm3zHfxQe6BBsH820OCO2XmYxMw
KrCV5nF4IqxxudSrLICNduh7Iy/jzgDbTortXCUbc1ohWdFFoV3PwIi9qD1SWobT
tTU6Kn80zR69vnnIdzpc6HXONabVoicNh/pl5EZ7LckHHYSWB6sJp5X3XwjbaBpb
2sqGF0X0LXkn4SXRW7J7Y6xvuRfCmEI36bZSm8HzxwC3qgVLqCZvCZsMAXIJSgH+
tIUyQ4f5DABOLBuUmRiIcWbb35+GJUB0xz9YQ5A7LmIQJ/WnzoVIzAEdxwaa3Sf9
K7d/DU0vsgoHxR+HlsZyfrif/uLXIa7cQnv+JhAQLHNCnvePh1/4IVdc2n78cHzB
uBm68Tj9kXUn8Wr5CAzZGnv4pUTEPHU5h/wS1fkaFJpboRQuv+MbNnnghKoz3SUm
L5/au+DOQRTvnlhcBc34ysKndKy7yRh8In2d0E32BFA0XadNyNdo2uHTeDaDb/Z+
Y3eP8PmCXtOEYhv1UEL6g8a6ViXJRkq93O8FVNyGwQ9PX42LlGm3ZuSCubfsAEBU
XGUSj14cpkY0Pmzf7C0u27z/t5tqhPAdpo3rWMtDaTfxWn1B/DKwLsqUuwGBEPRq
tX4ZuoH9Y2wRRRiEaHpRIrfk+9M/ne55SXdlY2RyIK17jH+AFWOdjVVoGBex3VNG
sr6Edunvadzfhdw5P+Akiwz4EybKyp7VILWUX83dIHnT6eQ7Mn2Csy9U56/oP5e5
03gA9WnsY8Dr7crtVmQaURSVZbkcBy65DbPvYQ9owjVe+NczoeoB7uUExiQzWqfC
VDTsjiwAr8ocAdVsG+t/I2ywRq8h8ajok19/7d+0nrxxL53tBazDOZuQR2QuBrgV
PVPXqtyMVW4FI9ZzVjt/Vd4qCHVj7WDWDkuONy/ukl+rViqSZD/rE1JaJ+b5MVv7
Vm74kFMd18vGsztoLkUojPxCfbV96Wq0fJ7YNbhZZSo3eauqJBaFAs6SuRSvPhz+
ct/n5v33yMW6UbSiCQhREUoPn6cR4H/ei3NvRqPZMOs/xEGhuH3dyayj53O4KsFI
rrTWmu/Uqz6PVeMpMAaiAX74f4k7NNsf9uBzabPwfb/pCxrA6jd3Pg/J+pensXV0
EoV7srq1xFnkqbNcKSwxtnSKlRKdsLHiy/gDPOb/ww3LVcgckRDaq7c8kcxuvDgl
ciA/TWHxcdtHLFzTFCxxNSwnWcoIb4u5xYPD/NMRuAYbfS0WVQWPAR0bQhakTLde
bDF36y0PrfLRRNUx7P6MImcCJDqDFixJOc+Td4MBrmVoN9sHpMb/zl/31bdYk4Q+
MkaXQAoAEo0AORhHGYG6QlFUNPcU5uZlGxSJ3ay4QwIolzFhDXF2NHweh5dRiox8
72jDoROzZ+5f/QoZL2zrtDkbQ7Jmk1WqYIH5ZYKacJWI5pxYSEXQhFvCCN/X2wCg
9jV4tgF0P1J1Z9AYJZYy30dEvRD9fUs/+aaFuaVi/U/aDIQA6AKKcL9pZGsCnfhk
1Ht67Ybf6iNh3he/vL+uK7Vm4I2rYz1n8NxEdSpjZo8Ih2DpV/RsvoXKYKDiuHvE
t2KapKA3mplDWDGy8j6jZjVmh/aQA3K0EnBfZ4lou/6PRIvllO48O/ARF0G/o8zt
Le/nQjNDbu+NQmqCUk2+ebFh0FtAfRiHehwccdheOyXVFtlxm3yQSWH1OC737tnG
mTx8gAj4gGxR0MsSlBOO9mrlLFYo6eY9KDf/963FyroDAARyRnOHtXXtZkSesVZf
fUsIAkBf8yVrile7rtkmObVY3vf6zAgfrKdKXwpde4pR3BMbPSK+GM3JW2JXLaGB
YJ+R5+UXDzfUMNeQUsoF89D/Fs8Ilyv516oBm7fI38u9Uw7MFH5ajmUX3ZbflIY5
9IqilwLcp41rCjTddFE55z2DU+C1UgxAL1ftruZldD0JkhBf85EoOne/ges9EViq
NbY5Sj4K90jboSq7YXtAxKMKgyiAPieaS6WtAmyF5mQuB2zRdl3o3mgjW6GJbx1Q
/doGAkyhdolLJIiOkE2XiFDNLUu23kAGshUKsfxtRHydQexmyleV5TF93HCwzWF+
JRDik5YlbooKb+NZCXC3D8zVbPNvbARAIDbMKUdPxE3D4TllRxAkUfn8BVY0fKUJ
XkY7CP+InvMp9sXnNolnju+KLWvHO5ixcAzSpty0ON0z69+48gD/3IKKy3G2cwfb
gyKKfq7AbA5Gl6GVIV0J2H0fqZZS9OZlmo6+bDCMzENsLaulpUS7+loG2pHiK+jc
9mLAJPXVojXenjIFCZCxXq9lRkD8wVpYu1EPfXaST3Z4Lrwin5Yyu5DUTyK0frUY
7DVuXp2MsmNowWhvmF1LFfj17S5ghmGeN0+4H+1zxo2Yr6JQVLUQWv1AIPRDku4u
fJrllW26U9Pr9DULy0rJvrnIME42/WZ/PZzwa7hdhcf1EPwXG4g19x6ZeZpqdXAq
JWLjzHE4Aaxbi5vbi7ocX8yaXWiG0zAI3xSWzHcC0iv6K1ELXHepJIsAi2LEA9+S
jr38gCRupSZT8gtxWfCWa+nboApFzb7ENUDbaKNfgf4tVGdzDxcpY8ThYdBpQeLV
xUqtdzM0W7ZAsJ6pGt0fVZcX/7xS/EmFSws39n0NG7H4CitY+r7ILHRt3gvBrlYk
BgZ5pgrRMB/jR+jNI629Cn2W3wVDyqccrV48bRm7d5aM2oM+zr0n8M5fq7kxbSWR
UEgvuARCiqw5vWywT5BdW4/AvoiNxJSdju/CDR7RaaDKwnz4rW7gbFawsJu+K5/2
8QXKkXslu+Sik0sb6dFWWXz+3MFIK/wu4gQ7vgJnCXEPf8Y7WJPxJdSUa7oUI/i7
E5JwCBdqE0VUMXLxzM9lLq1Mw3JBIdeJ3t2EAuBnwSyS3YfY4+TsbX+XKgSp7KTv
bfxd0AEiSDbKNM1OHLfi7IbYTJqQ1h+MI3giQN8trvxi5YYlakVvibsgY0j7Unu5
fD3tAqWdGxZ/whXI2gPBHdsgF7AxIu/dZS0d1jRFsv+Fg08//5pXbmT55SyuvSEl
00cbrgArENzboIjkvDKhF1HIN4rv3yMzjhtuHXoavlAxT6LLIZs9TBnJ839kG5rG
EVceKwdTMAh3PBokraaMikbNTPLW2GO2L1ZNxAZoKhtFqc/7lhJUzMLsAPh3wuEV
LRyhJNO2OAuwQpW5Lyhk6hxlkSdR0/QjH42h5IpxhajT3RG+LHk5jxH3878roneK
ef+ggnBrucs6t7hXWS9DmMQ28hRJwKovHhSk/HFZY/UgwGKvRw3XEXEutqdN+FDY
S6b5kQ27PZfmpIL/CAy7j+ScgjvHTid+sCrw6Qfe8XXqHOHGEvCTM0P+5sSB+V4u
WHde2HmkI3Y4bfop2C/aRczpxM6fF7FO+qE+lzJZnohGvk8DMOXOksu9Y4j+pBjk
RDEjjzw4CUmeF4CHQueFpFYNqxyLyPcBK0fWLr5AjP9VAsgy4tBrGG5iRP5XN9ag
9SET69W0HEgzs4nXDCvQ7aX5r8Aw4Y7wae7Gx1LDfdImNlDo0KvFhO7CkLHyaRP9
yvzSKKrNgSlTHRDjpAc7VM5T0usU1XYZ1wyYPpvoQR93COjW6IrZx02/2n7lqrx6
4CXHhhXSeeYacHJBs5KCz55tqZoyqX3cApepl4wK2gPjRm7H0lT3Hsa6Ogww3pLS
38OKoNBpGki4DOGmx2Age/7dwbpJruyQDbHGcZkGbKpZPRaUx+a3m5Emm9bXl/4Y
OOKU0UwsQxx2bHVs0zRZoj1xivAn8b0TWfb6FV4ddWadkzs00Y9YSDJ9J5S0Kn0U
wp9oUQlIWW+nWGoDlFNiJ1HxmAWX60kAeNkmZYZOSCCReqveJ6aA9Nsp7VVfH3Ue
hzmoVj2Hvd0DENc8QY17bU1dh5cUqQpIj68EbbDDCZ9TxPHXQ4r1woevzZYDW8DU
fFajccORcyNWfPu5xEt+4L8H5Pne81WnO1mfaRRo5lWzXNRJ2nKcIYkpMliEO3a3
JHGdegTcqvd+xPSkGoji3nxAs/6feBFmK6FN+MnuMf79srkhdpZylWrkwjSOJaNI
i+PCGdONikaDEVetb6t+nANXTwzvlzmLz2Xgs4zzhOuMGJbD549ehBL6Hp8iaW2a
8/Oier4VthQfK2HNo+IPuusdnttb1Qrycyh7cGHqoCE/R5PAdT6v7/L34Rx1ZP+b
HA+/YuIUPuC9C7k2fEP+K/dCDb8sc96AMR/yiTXs/2Dob6N5PtZMfYYFwEz1Pu4w
8ELD9/XBYLdf889p6mg4DcmvXYphcyqsdoXbhEyUGkyk5fVtDHjh+UDaNbxS1Z3w
MphisXx2sJonuVNDQuPclJxTQDQOOe1BMPAeTmwH3hIxAO6gJZrJCO8xj2CkwoCp
QyVJwB3s0pzdwsQenJzRDav8+vbFWZfMK5qC+xys86hGzNBSVG+ttTE+B4Y0/ucU
H2dnO1zXQDi6ZY9RvhPC1+9AzNm6OS8bMTFBh5J7T+xlkl/V2yJpjtFLILa0Li9F
fGIxv1pDsZK3/jQrDik+quuUYIySDBl5p7Cx/cInUEGSoJs50ozk27+LUgNFHGiu
fVeHE/DpogjfiTlt4iV1h/jONmWhUZpY/HnQScY6pM1KLK7E6w/tRbbZbiwgZ1Dq
llm25/9Q2UKvSISOMwOS36z/aX4EvqOMxW2TRLLnnWtSuiL5/HAti1GNKz9g6CA5
hWUtUlwh6NHG1SI8JRL/sIPj21zCT+egXUYP3Ay5oPHdc9C+QDPZxCp8nMR9Wari
HK7hZ7dk+DCKZanC0LU8FLX1rhNSCvg/gdhPceeErdq0Kb8lmWVgvfNerhr92q2M
YqdZLcNaUnaiFnZg4RIg5B/LYn4CvGc693zPToVBdQe1TKcKfmah91AaHf7MnUrt
keHev4woIpAneob0I0pvQdcGbWuvAYT2idSxV+NEyYL/W9ml4EfHSthDRfApNp3V
LdTgYfSivY/KLVnNLoORDVmR3Vi2dKxH8U1/sgR95n/gmNNLw4MD8x/nuWN29frp
NyINVw/7dug1frMVeUgSpJjGBKAuUjIy9kC0s+8CBTVhNGqjsbIh3WGVCrZhRo5J
OdtEgqMF+XBbqQohl03pPdBa3J9gzERsrV8wYJXGPhewqM7Eb791OuHK6hZ6vz1Y
qwPbUb52/ope/hH0toer3fonnFMTEVP5QvsbrrSKrch7uNqRiEkHOXF3k561BB3A
cSXc6EJXTus7JJMV04pALw02T9xaDcd9ouQGI1ydD/rRWvaDBOvaARmSOcaQJw+E
JnTJvSWqwHA3JqqrIlYHvku3L4ZOUAITPeRgqwO96B2ipPaCl/fbApLmew69Dhat
J1VA2OrjSwVYkG/F9qBHDry1LOdD0L+gQOZiLkc6xzCV+HeUA+FhBwfuiXrMbowG
my4YWUYuaWgwr/qgkf2pT1JZ3Fs8L+dj+aUWp1EazxfkZGxVhGmymHNTl4YQNKtm
/6O0S+NCSp/mIALyh9IdbwSRgSDvAgJupcu33c/xaNskZqdeUWM9HhQMUY1EvHNF
AgWyslU4J7sMI2RHznTvumgQbRQhsmZvLTlEshg1V2keuhZR5H/XYzYG8tNnX3Cy
OFZH5msPgZQqeRNVceH5L6Jgm7nJUSEqYGt8ZhUjO305zUnHGz/MCDaWVtb2sVkv
5Dbqs3cVS/GwRfqLoBK9VSWjIfnzSDDeUtWHOYYCpKIKMV0cCcOyYd4m75l4nQmi
BS1xawySvUtxf2teFtUrISrstXBoUNDW8mEbOA8qFykjdYGWVIqHIqBiBqM7EQTX
RjPRQ7zWuIbSLd1x2urpxBbNow/y3KBsACm9XmBonPsoNkmNY9EGl080Aooj5jgr
SqRdzMH482qzFJyZgP6lkCvN20g0uxUYZVce2S4lMa62oI/0uhtlhAoJsi073eZA
eDvl9F0gbDVHvXr5/XrUJgjp0fYEcCE6TfXWDiceUnkRPBXpVMGEhTA3wbD3joMi
7i6e00J6zVDwTbNFAevWHtQAYkCBTyOrgWxoOzIzXQnswvAcrp8+rn0aJ2B2mLpR
hzogMWP1I++rApKInUFYzS/RMss75fH7KNYAc//LEXxdC2eYMHueyfIsxvAunO3w
5F45hk7Y9+oRFpIUODBOocrNmNldYpF1nhtL7hzKEd17NAkzGdM/rWTCVEco5IBT
FFYEf/Wp0Vf2gPgLFpHzL+eu0oZ2uhgeviZln14k3KzRg4A52ZURJ3IBNBRLvRgL
PxHGvaLR3+j5eWkoj0E0q5vnvlGYg3kLRmk5hNGLod/nsflrJPxP0GFiqIdwRR+h
65fpxgj5jXR/UtF9wR0n3KDBPH1X2CD1uAKFXLGJQkzHh0WCCaKb+97YdhHDGR2i
OENNyNSaJ/SIvVoOTIPsQp35ZRB0YO7ap5BwW+dPA25lDc33kdSn5l4J5nTw/i+v
7JFsCB/xWLbn6a1A7VFHpgJnnD58DJIBRztbQWEDcAxb8i2bFCdMXDuvK/4hifC0
6nYKt0/JS+hZuX4VbxcT2UTXT4wad9rCznE4zSZsUXg/zRJ+l5MqsIOnYcHQThtv
n2uc2cSO4I5NgE9RNYitNLJt4TcUHWfSFYoRXNI1lxpq3w1qNe2JCeLWmOKz+wWs
xFWX3txaC5rTYUFODfkykxblPoCHkquZAtxlLuJCGJaA127jOtGm44eqUO5Rx9fX
lXngqN+sPFk0NHqUXqdCpR1PAPqFtbCoGWLgwyqNnPCQwtRKkYd1D98dblwg/wTW
v6kq21HO4Zfez8QK3j6a6RM4dWL8QFETfsDWmyUfYEkr/l8kIdnPEPE7ooLq1TCS
QVUW4WhDgPi1looSK/WqnpYIBhY/E+yuBrflcUsRHKymsLUMQII1w1yXmaDybyUb
W3+gKpQ9Rb7RsI7w6ZcLd0n0I1huscVL7X6i2J2Asbws+68dYGCFSghpCBaAmI7q
8DXQAP4tIXaHWpoNA2ic68Hl5Lz/+NG4gvKYeityIPiFZm2NmJiTUg5A56pGPUIq
evjljlTIWpEfDOdJujwyt2WgtxP8ts+9NCJ8j6jVSUfr0H3puTmXlXlcj98Cll+C
oY8AlPTWqJprasOUUndNvMGE6z4dyQbw96GyUpaaHV8jzJlA5FzpsUPnaDJpIZpr
zP0o2z6D8l/s59E8I7BDa7QdmeOlA1lrMBySBiWiQXKW2VK4gXGVux8dINWKuYLO
lTgAf+UGXsCNGxfN/+zZONNPD05TaZrJoqUpcqmdLp4DLi2jPmvbatQ/xLqPVth+
x5fYEnasMP/TQ77MmWvxhLj9gnmrH+urJE7xCOjgSHSpu4YO1f41XX2H5K4jBxMw
IydWfXX3Zy3zSPwRTnrivGlQhoS5NS85ckZ0x9kN+29dvK2f3djFq5/AgIV6IPjn
GTX2RPftWgEx4nUYN4o6JGxupfygGaZyueAOIMGMXuRdkvLGcrAnYxeAKshOPEDF
rNNWwmjWoyFxbZ6uKRvk9/JC1WH6fr/GGi7frg1JxTGIpx11BiG7SENbVUy3mE+n
3vT9a+TgrnKzKm2BUlCRL5SH2p0rXmc4+gf1kvEoe+CmY33l/Eqmgcf3jWrYR7rF
svpzWP8P2AfbSiutCoymGUV6wKZg427DnjVe7/jsjtjGEU9ADghlxq1S7975j4hm
7EgPFtVQoRsPCMnJG5fE2IEpmmBXPKwM+Hq9VUITVv9/Capv+7xEY/89vQtGbV51
WMYU+k6tuSlL5O0lnfdqOMJoWhxAvj2VnZf13SqqV+z2FZGHf5Wo6t4g8oVXehUk
9Wml1TsFC88n+9b3ykBTFhhSysbH4MExHCLJlwfjd9Jz4wc3h3fSFIn+BGbaGE9F
F5Nd8yzHtA9HIioUmejPVnN6CfhMN8gw5wPrmtJII6z5a9T0A8l3EiiAcRe1PBF3
nx1XZuDr1+ONHNh4GY0+lf9o5Iw0t5s5dkOl8qprFNTwTprdyFoXZG77Ts7q4xjV
JVMv5PsEEqlMpMNMG3OtJjI0aqFm8GIKhEVbhF3JldKZY0elOcL0Hf8KAAtDG02q
Jni98sfWFzINuuGXKRl9gWWsKbi/eNzC741ymIs7j968obavZ+Bf9sTwVlQMADHy
1WU9hMY5DEyh1b0mp6FjSGc4OyNGgjELYKDqTZxwFvPoWIjW9cKsngDlhxkfrodt
gTTKWGwws1veM4EM8X5O36GVBidf6jTaCxNWCZ4BkrMRZm1MuG+cADGq44pSE2IA
INZE+AE2bDUqCLJmVG5Mlq3pRzJj/uz6ESyvsHxwlWt2pjr0tVUCadnwvuf7dNDh
cssBx+Kg8+WbdBPsphhC5UzILK/QDQwa6DcJSiF42DsZBX7m8pRT6WDpmiW5BxeH
35y7tyO8N1CZ0JO5VWWKrmz4SlM6t7MUgbgO+Eo3dh3NvWozB+QWFxxJp0b+RpGd
WGCh9ayucGvKDynrktypc5piDFfA2xevo/p7KLPgSPhMV788IJHrT1JqZXWoJuDX
LfAxFiwHzyG/Krbs1ASNOEzA3oCUWFFqNWilJ7SmJJWeBeDJcArhqURR6HasUrR7
9TdEFjO2DZLNkciA4wcOe5nvF4xxzvtwA1L8LN09eQt9hyy68bB4anTpt85zORJ1
sg5tPL+PSUnItrR0HsZTbQ3Zzb9arPGSVQpdLk2SKtoBODCkBHSH0OfWct2tLpn8
59N4uroCm2joqtusfeQ3KTnCykXcqoYXuBfrotE7KzDKEXID+5hMYw6IbVALZnxH
Tt2gFMIEkC/awvHOpszXpQRhH1+OGPAN0cprJM7AJEnnf+xIH92SwOTONpnl5KJ3
NlNqsjuSmy0RL18L0+G16+owOzRQywehLcLvZcwrQ5bBwj11p8weDonCeghjrZcc
BRGkKdkG6h/x3Eh/KXTVYwk7qyji+OmpfwlYsH9B+b34RRXrIeUdF6iuUM+0c1nd
zMOkNk1SJPnnyDtajMab37lMEAkAMlF9Ql1ldmmiZQBH4yzG8sFB4TCEs+dgnEff
ToadIOnHF5vAJDKkKS2B/vqiTuCs845hKP+1zvfGezMk4DofJlR1JwBHiLabhiQ5
0hPn9bRaYFx8s/Ry7WS/mBAyF16KTg7EpGJSoMSJigcqxOxckaBePnZ9vuB1klH2
1IF68NWVzU7oVo51cNU85z4aKpybILfafMT37Ee3RGuHi8/Q4s8L8xsunLIOwj5u
cZl/z4viUeyHoBQCj+QW/Ihpnx5phW2lhk0j991Lies4v/A2nPUJxE1qb7SRL8O7
c0F6sgTB11feuTtXHDP1HlljL2K54QDXQolhFKta4ZFcDenBZSLddRB5vsHsLO+X
t2Bm4qbwh3WoQLRfFvbFTtEibxvspQu7JwvoCpJcpR1JHyW6X+aTZ/zBP4G26EAD
F+sj6y6StmqweyI709KZFGnmlhkPEmfP29r0Dh3RWWwpfwDtlIaekP/ffL8/JeVp
mcMPDt6CZZYY3qSQkcRet0REIF718ZfjfBktFJv9lEoX6t7SZeoVvPK70QC77P9O
rymKG55xOEK29t/5ZY/BgO5bE/MttqGEWVCXa43KoGVUaN1EnCLRtzPdSayb+NGN
ur+8VnBOo3jw4NmG9KU9mDft7evTEqMuzcJVqKz6Y+vMM7hCHi5dTzFNsCr/Oygz
mdviwOKCKv3w0nWq7jWqHdQW1gi4vBZ/Jz6neC6x25APbwOUQyWdclevriA8P4Ut
sTe1WgdVpVu28jItOnxy9lXTdlHk20rogVOBPNhU7q7sGGq06ACqH02i3M0H7riS
77stftbkiBdNdxunDL0L52zEW8oia1EbTKDbdCf3K9tM115oJbY8eP7L+U36GXQB
FpLwPJIE6JyBJn4KhELXnMYlnyqoz/Uk/xYBV9KoAcCBNOEMjoY+rqcRKzRLtLUB
AEcUFqzCdMeSvMDmYUx6k8KV08aAYdcqR5UtrYykyi5Oga3/7DrXfgZX8yX95JqX
Mhlk6XuG8OIvPIRlEHIwcCLNW5xNJDghjtzS+YgtVk7DVOEQLNaW6/Z54QMezveO
HNqE75McE0ci1UH4xI56v1EymXDRACwGz6gRSUJeyb9P7nZWLQ8iEy4QtQKx9E20
7FyafqcofzCDj8lBlM1rmh+sb3iYwIEURuSUYji1HlPnF0ys4KkB2h+e1oUhI5YP
NRy5z8nkyOGVTCCYYoQf3sIsPc7Y7yuTaUUmif8q9tivi+O+xvMI8gGTeUWrLSZ0
NdIAuFxVYXUmPrSeC/mKZaNbZIOmOrFsh82UFYfmTO16kkZclHm4XAK3gJ4WQ3wf
2uRt5fokyY0d8Tu+miKAum2UVshzKuGu3C0p8++MgzLPZxV5/gIpgjKxLFDzymF8
e4OAjFMwNJQG+5+q+VE5Hy4bHBH/bfxW38MZTbjSh4Yqmc/NjR2apuYEOBjeRDVw
mrrGruRpwn1ZfWLRfSsjHXxzuRWZrsEy/hQdoatYHt+KwdaA966GTnGxnG4mOp4A
p78bipwJRRFclifqIU4sqFh5+I5DfETL6xwz1Sdau+0VBZc3XCmabZKU8s62W85h
fSkQioi9EXu6Km3Myb0Dh6PVeP0fQdd8dFqRP5PNdOoz5W8jn7QTH9GkpG3YRLmt
0UqA5yb6exci3/4XzZCGU2KUm+084QlM54Agnycgzb3TCSR4Hx07yWPr0QUK4sgd
GJxyO2oaJxWCTx/NzXxGRcB6N0CPtNgUn84kMg59phMhtrf7oD9hXA1xeXRlZWIM
XAWMQJVQEnXMw+2eA7E9h0pZnUXZ6o9PmTeQjMqPu+5LngEteo0lUGSYDtc1wSmm
0tWnHjdNq7LggbQ3OEk58qkfAao8LVncq4QS2XNneAi/QjGAHd7P1n+ZfJW9i0kW
b55whomKrxIfCcBckhABA0uTTTUsFpnOpzRMWI3aUY3w7dBZcQlO+Jy1UeshkB2w
g+UP9RTQGAUcC7jBkGQpMeZeWaFWv/6YlSKR+RnwbWoC+K82nIt3cA+x7ym3HdOd
dHP4QOcSigtmcA/qujSPMy09UKJcKzO7Yf/Mobfo0k8UDtN0KnAuMyn9C+4EoyNU
3eLhEb/pwVYLprfz0BA8YRTgwobK36bPLbnu7y9fdCFavcrSviR/brPc5CmN8oPi
eu9fVO7KXX1XrQ7pCPOZYtWW5sJ6dYKFmBTsd3bpTujR4Yrx9bKSrt23OG2jc/Ml
kliwuzh6i0ixtR6jIZh9eTr1MxjGnCcF9U9ScNBVAIpVbdfyuCqzMoTva1yPTbYx
qSnf2CUmUvCCoe2QNWoEkMPtf5VBKlnrrBFG3ph693k6fjRVyRqyVjvHnyiERDS0
FQW8gAeA6x/EuwkVCNAr4cGLT+Woj3l37XmohemzTK4M8xcJVYi6I0tPG5nma0gm
vt7l1YKKMdu9dithqGcx5kgUvs2ycARqGNyOtzcwmK8p+NOheQt6oC+Coud5y1TB
fBb7P6VV6akFGbKCaI6QwT4bbYE6cDvJa+VBMaAAO/uKVhksbddLBvAiC8xNg8A4
3/gtyfD4vJ0o3KjI6SLeFDlh8YDVdWlQ7GObuxI2K0XVVuphf8WqKQlHO0RGbv2z
eS1QFzbZAtLzrVySQIcRCwAqkY4OD8X8ianciGu6cvSDUJEAYlBFoBehr3sO8AhA
7Jgr8wrRTinYdktfyfMHoxs85//LvM1at+/42cBaIg+AFX/A/fEV9/pE/of1Ki/q
dwphDLTQXL1s0JISnfeGbab3DZiAtb8WqcXmg2JXxG6WjYTOs4/tGrsLqPbf5qR5
zFi7jTmIvD165JN4tT5p++gST44gwFmZtNlHZfEFEUGkTVjF3qMzVpMjKDTYnzaL
rYn/MVlk9ZenuUNpqNv7OSsQxXberH4cWfL3fD2sW0i7O2oy7gQBYETPBKsUw7Ac
k3A3OWEcdSJNy8fu0RsD3BJ4LP/x3penhEH5rSlzYSQyXiqMjz9PtNceqZVwKd/F
na7iCxdhJIgUkG0CCIJQRFvrs5HmiboQdRL/ocgpD9LA7FMqxtZU9b/q/xNKyAjH
FPEj0X5t4RWtQUbQ+2LRzWyOKufzUV2qYB4Rjx5fJcsudpIKs89yCMlGYU0Eprjb
RkuvvqFmEZUo8ulJsvqiNtWGsjB20dcsrsFEFZDx0wyLsBY92BUaZMr+M3xrtFbd
IMFGul4jnggXZqYEwild5493PQ8IzvA/jP8BrdaLYTL18+myDJLEzk5LbU5qOSj1
DYEFRBOAp9208o0WShf33EA6xVWGIfFMjqINYfsZtd+UpYz+haf0W3MMKYh/9SoM
ri6A+mio2bv7nsuLzpLvK5JlkZctJkyYdaW+Q7Xubf8MdeXz6xsO6+lSCnBkuH0A
dbdl03L9jLccYakif/qpRHJA1qPu/vsAHNZxrwbdZ/aESLjH3cSjEvEV1Q06Nern
dBfcp7Id9h/mPEaHMcrBZANzDYrn4J4NzjCu5npynEZnNvubOtsQfUH9Fsixil1e
9UF+pu8RvsGoF2SQsQpHuIqitYcYXGrCIWW9e+JjBVT4Htl4O6qYmxefwAsByHTv
zPWkY8jZub1Ssb4+VWx1DIRMazbCmFa8uuMEoYIBBLk1zhwgvn9rosP0w22lLkFK
x3VdN/yhvYP+w2k2PtXnQleY2cK6Ad4ryeHku9SI2aRY8mYlVjXCGuC8lFvKA/81
FBympWl76K4XaS3mh6bFaclgEr6+psxv+1+OyTVM5hkA4ObhSPn6mOCrHerCyMWc
ye76cPUrcGMzlpWdqSXhXsWCkoRzC13kQI+FOujT8dI/7OW27ks/h21LDej5/8Uc
MSVCHgWWqGtDRbiYGRnJUX0iHN5yYxli884/wdVZ3+he1E/z56RV998RHMhFG9bw
gRbKZP2j1pZbQy9ng3yOxZ4tnNyWHCR9hpICTxG3eghtE0XATI/+flO0/OpWt6kg
wCI89YnrMs7ebYPtt1PtoURXyTdtKNuKLUJn8mn+iTmwZSJvYcu2T166HBmYs5QN
dDCT3XZLbZjccvihNEnJ3CB2b7Tl8+/tgJ0f28o6kJ4Ps8Ot1CQr8ClJFuf0VvUD
SBdhKFHSKfLrXZOddWQqnUWDg+VIEq4f5aTyhPu34ICZYO17e1oImRCFvL0aGnXz
lQMGla75HvbnYAvcYipJQlInRrlQBBb593xPuW614kK/5JFmz9j5ex30b6JVfUUT
6OyBDSJH/2aamGSW2RQEjBqis3RDX1YQXVODjtCXvf/awypQZuOB4iyea3pigzHh
MRYPGvT80HrWWFWNV23Yv5/EMlnblsN6+Qgw1RmNSoRlJmJ0nX/PbnclKLS37VhF
HuKFNSk2AKuNvLBLL+CiROcM1MgvIW+b2LOhKuVbhE7iWerjwAiPPTLRI49MluRs
f+9gjAArFlryhBegd/L+WKWJUqyMPRRBSdpkLbmL2NoTxgf8jywYjN0u8nfg0guQ
dm0qkUyRsTHqy4didWXdXlU9+3a20VVRo234fg+lAzTF6/VtFHJEIepOruqCsSHs
8Dr+d6rP6auMQKba6xfh5atYtE3tu/X8jq/ORxmYFGf4GImk7OCPOKNiQkJvHNxZ
0IyVQz/VQs81JxV2HXQYhGTsiXSrkMWc3Dr88jVVpHQzyJQn0MF45ODaCfrCU/or
sbgEXEvwALxo4ZywWbsm3p7lu8s7h3VMKx7bQobzJ7YSaUiiaZi+b9PqSRZBdeB3
5c2MsSoWtwoyP1xV9Xa4yPmYgflWuZ6b0fBKlE6++kaGlxUEvG1t2Ha0Kcp+SVyc
Eaf6X9oynJrktXunBkEIecS4DJLZ43Ay2tfwmbiXJVOZTUJuEFlTp6lSXkbl77EV
Hs3wfjui4HElD083lyayEGgTkL0KcLktEK/sAyUAKiCpTMCaIWHtVNO7RXhxHYbf
1gTiw9QwuU09tARascpW0uKgfacpy5TZyXNB9NbNes1gJMbXJW7G0+VgiVBVUGYa
9Dtk51PJqNWCqCdIHUxih93cuUwlZEK8sW4ZGsUDMr+vgvNKupLE0o7/6GLCwfYC
06vjZX91jgh0H8+Rf9fZAJKncBQLKIGnrBW/CS4unq+J7rFLlvqsR/HCic6X3ALK
QkbK2/TyiGQLuXfl2bg0npALdxTwwGdPdV+LxrAen0bJfo0EFEdOJ16B1edcDNOp
LAHnqcVXsB9/nqRguzK/LakTpGqJ4MgIEqM6XPjFG0UcbvambqQ5GTvzraGo6VhL
51tI6ktODx1OJgLfXeOdIhdZBRLG7NDcIUIGkJv++6XMpnVJVM8psKWBwdi53oT/
0VkSUGiutYyMIeJ+OuoKMGIPFrXsfqH+EMIn0dC5Dj33m4MTBk1LhJKot1fjPYzT
fpeloV5+vX7XftiqD4cdakmZDl6IGSNDyOqz8EH8EukB/iK8WPfVeXsUUVedJDLL
Q/LBdB3v0mqHXTlcUtkqmIzA2jG3IMZe4wFlXMeOFe6QnTdWX5ucvzyl5FBUGaHd
Q0kmTh0Wyt6SxGXbtPYUelNFrlvCrVHxgvBlplVzgxJaZuzHJwz6Z3+UOUBw58aH
mNg1vjbWfnvjJGUXQbN/6OmLrvNzFVNdVSInTtYNyWmQI8sREmzfdaHGjttPPTXB
C/v/XB9kIYsFiO6L0NFItmxaeGHcNSvVrtmjge7kEHZLf7MiXI/lbyVOIiDGCJzn
HeOGS1gRqcpJM8PTcMx8+jXbVI61s06qycBgF8jb+WxxMERboyol1bPzrLMsZtaF
OGNQ7f9PUVm2caAXbvDREbOaaZjB3ZUH8hP7izvthCVkBLkzIhnjFBQs/qGaTpCs
PpW4N2h5zZoQ38ygBHu33ZHRyofp16rqSXNj8eHgvA3Kv3eqDBfPeXxXZ2TYYgkB
csFFvLfpgf/TfXSkkkmgXcYzlJEKimsKvoFUIRumnHQ2yuW1AEEqw2t9Gl/CrmsH
+X9+zc0XTw6SrfMFRXLixh5nEQyxAhTlBDfxz0Y1rogtVgFo46fMbC4X1MSZpXdt
6y8rkU0/mlOQJEsFBYOEZpk2m5s5OeBQXKj4VKaH8Xt/duzkvxeTqp6281P2KwXJ
b+EfepW1M1s+3ViHce+cQXyEGVRNtlwCgYthENBpSqWFmD1e+zoVyQ13Eadx8oJw
YSnUBE43XAvrCWEY2+lKhD7ebTshXQWygoX/U8aduE5xsy36zvnM6cU1O67Qw3h9
pwXtfoFLdO+3jeF/wDWZfBaIGI3XPiozyZrUL7dWgsXPzhaCYyKluU7nKw9z/Z59
6IH4+ft4xp9ct+46SQhOumLrObDQsUU0jPNsv0Qy0N8hXHuydE7rFtWVB0wCjoGO
+d4X0CilbsRxINZDKYX5yn6JjARtBmCXkx26a1NQC1FWLcqxrafMy++bZljrSoEE
eRO6pyq0L6/G+a7rw3Qmn9ldVfHOv9STzba8Ww2ItP8RsI7D1otuxZuB/lZgExnv
6tvXenFXm2DtncjYz6MVMSUB9kZKBexo33JlZBLgQsaCdnxU7bkF+EEiX15h2Vxl
AvbmHmvrn/Gf312QyBO+dxnOp2Ebp20YMcvQRtZH+UoY5WhkUEbUlsJ1l8/V2I6A
ybQly9oZhFgoCDz02m7B6bDO2Ny96vWhtg5V4yQZHvoXaAuDsi+z5spoC7gSuedK
E8WqmJIjyGbHAN4M7wDUAJwHXHPUJiLcmq1Qi/4wjNcar+2ctUa0UMX56KS5VqqD
P2aZOPJ93o5MqvymiqkGDTgGOB9LxuXEqAJCD+2/+LkglCzdX0FiMjnJM1xXWZJG
5UXVgExhY1QJaEZ4r0w0K+FDYJgr3P8nJyCMW55Y2mNEZHp8zMCgrADd6XJ6ZjI9
5LVEbZpM0DM4kdZqpa2rOHy/RZG6L/gk8Z06rLguNEdqbWqqWMtt0q+iUVA4biC5
kImg9BornbdAv1R+oG52/evmI8tifCJxVkjnndY15V4bA+au+rKI26xLeDTRnmTY
HrnVLeIZ6xDFRzfJxgjETgkVq0foDfssA8Bwn7/SwYM/fCCoSaFIMVS0tXgPw+g3
Gcvk62uIz4LMCkVwXyV1BOBgcxvBTq8ReWm3kw02Awgd0wFJWMY8Nvrl0F5Zu94h
QAK0d1acGqGUFMqtRXodv0dsUOtpNB3z3vEzH4gqo/4+svHFNOZRf+HuiAEW/AOO
4V6btp15Kr2Xv2r14GnCiicvSeigjPwPWPMpKUsoqyjs8yS5MwpqPAPVVGnHoup/
Mc878U9LNjfTKDkzjaXijkrLX+ciIIvgFTV86iqWRWz2Sw6sFq6lQyruqyiacoTj
ibXxCYaUzEUgt4aRaq0JCMtDXHG+seCCC8FQuXmKHJ1ZI4pd4H65vS0grJO7qyyM
EtlvTPc7saeda4tNLP+5KDLw3fUMu47ayiGgk484wc77j9y30D1boZDIU6Wonr8G
S6+pU+amheK8KPbH//Cev2K4iso0jWujFy593mdf3igiQRDC+2pGA8YW1kqOJZw1
cvBEJDwNoJp/N19fzTkBPawSL+Ac7IniexTocWS8AqhONXDOnj26VljTSy+PDZP5
BPuPuwtu6rtJrW46si/IGI9IFh811yhVrYc1vL+AhI8yTnRy1xGzmXy2dmUcDv5h
6YRnBmto5md9hhzHMpqQQY7gmt/yT6ETtPLwTRwiyAoa+AGp+34EMuCgpN4JOhwH
xJcfZnwd4EI+lC3pCvBQqSFToeM0crm53EOk0uPOFrB4eTMON12VnMU7JUfg44jR
G/t6nuyHUG4cWn271Jxc+k8mWAdZqPAq7Y6JXGiosZEt1OvrB1585U8ldi5aGP9Z
IPylUntT82VED/Pcqkok1FNYXiF0p81nkIodRY00gDUs2QJZIDaHc8XX+el2aDQM
3wu6o2Rh4w/s0bjGuzJ2/3D6bTH22tBQvRGjO5JCtFhTt3syv1qrx1IEWw0cD0HL
Py62dEYINll3+yHBa1RrYHNuOtDT+QIc1UePb/JXc4BfHjPnB1sbEgiTreuATEyX
ciTNjx4NCKouMpkw4211/upzt2vPPCjk5JEXVzU3MBPb1s58F7IuHoeQl8jggiy+
j3S0ltiTiPpE5zg4TKh301lJCaTbVi4NkqZncgzjxrE+FOe1v5pJqkUrBEpCF/w+
GuCH6mPUMrRi/DO4HuKSfp57M1i1GAU5rJlNLz7fnM++sTImavY/A586R+K9PY1+
XQBOyTk2EqnKqQeS0pvBkzdl/jIyhEpuqGwQ96Ng9YPPd2lYwNB3uKkRpSCcgMpt
XkUYxGFJPSFyExY+4pvabS3GHG7WUGxE36vf+EpmxqvYBWFPWxTjWDLHrue5Wbuq
zIAvzNUpsB8bl0s/KwcHlloaawQ6KuAL8/K9ErNJR71o9+4avBI4Y8srC16QK8Vy
ZGzh8Ig8hOLfToqbHAy9591aoKV142fcatgHfLVI27fqM/qswtxZOLkG2IU9a9mY
VL4WUrCrrZLipVR6gmG7rjjlGLCmYni1GO0Ji5finXfcmOpqdby5ZgQIf5loL8xk
qQOFD69T6rdGnKcjEWk/sWvgZGlhIyJpeacUGg16EJHIgXKlbSHLAoduYdSMg9L0
wSc4GkL0rga291KMcyyJnWzyZq01FzDLfLM6Q3g3s6yPmUfX3cdmt5vhROazmNpn
DqFk4fTvfaru9di+bHnRrhTHOlUh5R7Hhtkf7dG3gOstT7szWGrILDMQV8ucrb8J
RHySXsNVLxnYU7zCscDOKB2kRdSueudN8Hu3T2+zanpeaaHl8r3BSbj5lk+KKYBn
ONarMBmI4z33AqP1rP+7EuSCNjSwaCuDQJNnzlZjnojkOE4NTGpY/q71ddZpoKOs
SZA3s8iAwga+2/T1WHj+cTWP2vzUIAKaN+qHeZhV38L4+xfkf/zbuGGXUjXch47Q
3lDhjYx8c71cMa9yN4RFvHz+8uH65KG8wODqckXwGUBj5FTeTxnZhcIjTbmFdsEC
+wqUgV6794PRkIQ3b4L+6j8trBBx7mgzTT2a08HciDO/SIFJLH504Iat0kbUjrcn
sTXm59yjSLsHCZ3ap31Ii8fPig5Or1Vuueg7xtjTm1g+vKE8ogZ5PFTATlqmxC/V
rS/Jzy1ODrSWd1YAQGMD7v3Qk8BQgAqdVhnway2IBx03ijwvTAz87/lCQBr0EVNn
NA3DOG1CppkEI5iQtljbKLz/dOYKyDqmlwza/bZ0ySXEOSIFYXXZIsx/FYqm2tY8
5UFYrclQ4/GnyrfiYZLPK6fDcYZtMShUsWZhxdg6DmKva1W8bNhHE1TZIK9XJvBU
xOkMu+Fbl2TYY3GYPRDTfu9Uuxzl5319inczIqTajpi7EtrNTb7CCVwt9OgXxX1H
wpWtacVrW9m1qiiOnm9MSR4dbx5Hsqk+KuSltL25DWeD6cp+Vw/HTDP0Z0ZlWcpq
d7lT3oxKoxKPIWMpegmpAYsuCD4PMhVvY3i1W3z/SJmrwxR/gddJzaVCfUFi7TP0
tWZ6nqMPuQFCumqB8dzS7AQptNIexPuBT2uGiE1+EBlAPDx9dDS8IYYuNkJwgslO
srdanVSqrkpRSupbOrPvyPcy+lXi7ifSTUlDY5d5k5LtuGMpiSH5ByTQBLfyzySg
4xT3CqQXr+wweHBg9X6nzhbgCk7l7NWaMW1T6qgXBwTOjiZ4vC6OkjJaelJtxO2M
44JJKBQTju9MvtUSaocOyjjEk0Xl11YAXJv44J8kWL3Y91k4sMsvM6B42KeAOXAM
csINvV8gmaoMV5IUN/6JFr44nBvl/oQCcYGQK7ZUellKEOB1DHEyF9NzfY9bXJM/
SPKGKhWKY8R7uo8oSwIcGCIbOfAGDwYDaMjlRGlIJkxQtrjANbvCqjw017eFnUhX
TDieoUTpBN+cQuAanHhwtCF1ZDAGzcdbPnskNwM8k7UFa1iLDMMFWFVV0WxCb4B7
NFSC3N8ZRJE8BTLn/VxZg10Y+BGVI6YjcNfg0JqI1wA8TLPK2H14UqF/V5cqVNPW
h3WR7Bg3hm62GL7lp9/iE7fc3Gg+/CSFG/9sjG8v/1J84/Y+ox3p5lb07QLmGThn
dhmatU1XxmE34InWfFQ3hMNMeGLJzTGFdbdexx8XnYzHe2k32UjKWk3gSa/PJogX
0z/e8jFQoXMhUmIrBBSNQPxs4VGnKZ16kXLcyp4AB4ZFAP2W6HWa+Z7AIi0id0MS
jG0BAE44x9OZRg30KusVxj13uwdJevzbisQVoq919Eb5yLKrVSgrG2BDbIf8IY3W
FHTRmEqbeezYOpV8LLegW/QCSHsb2f1qRbC0l5O4/sFfqfKjngAmBCfHgeW2Elb2
eStrRPSQFUIbyPGG6ywc673O1EElRsI/rVGfVdzdUvbzBYWqjLs+bcrrlO5y0Q9G
gqsbaz03K5PlQsDl2lRghDWxd+ZhXaX4wt6jJ+eZG9jBRKDkFJqFi6fwPzdJLMni
F0QXTKe4tpBTbksc8wXuD2hOlo2a5Af+qlyRloPGSn9RC30W2NwltR08YSOetHc+
T9zbVI009lFeCWFs1RoTqKFFSVeTOfzQeElGRvIvZCD/lE24zQbNo5o2YxCg8WXe
u8Oq334RvyZxqOVI1mh21T+81YFDTal5qG6YkZbP9/xoNUyIcWtaNHZ6Y5hR/sT5
CSHGRxhPlFFomFFChFzbJICg6WCxDcdMJGGR2c5eyQEbzQbg9pZR/i5pF/p7kNkL
MWTG2NbCZ1p9PzuiDS0iRtv5pkP1WrMTpdnD0dQJ7THMgl2jPQciEWGYTnrSrKPf
7G8k7/SYL8ScG0Sxe78/UQXx6ZUFuzOWHHhO2Izk7R0f8Xx0aOl4WTN6xNJ265YI
YT6nWmYG68K1HeFFrFS1E7inzveDFx+aJqo0EQq1m5VaFPCFtQM6iWHpznTX45NF
Qf5t9Ja/vNrq8czjTxaImzkMpEJqFz6gBObXaYh8myshEtzNmqDQfmnASZdwcgbJ
9+vecP6+24ApwmptgHPuMq6BDIOupIx9k7W6SQmqIgMQoVR8lfCEQG6Hnj9cvP4n
YDBf8ZR7Er+HC9GvVHMQHceifHZFTNRLn0RqlDqfspZ2dUcEZUTTr2HXxpQreSoj
YofXF/npvu0qStJsq97EzzVoASV2GSQhkhiJX277d/jxZhfvoEAgtGpmbu3sPS2c
gwZLPUD+ofgfikcZaOZX39tB593LNzruhxiqkxY+g3z+gYK2VAYko/GsJ3S9TdQ3
9dfdahCZDWm8+bisAXVYBdI+7qdnQ2Nj9kokByHdIODuFmSPz4rEvPNDbZOk7ifk
hm8Eedtxczn3vNMT98hpW7hi8t+YGSAESO8FcmS/c7XBa2/uz249B4RE9Jg2nkiY
f0H/3kj7jJQ43TeQZAAxt/FWg6nC1ndd/kigWWuQ69NOHwl0uczbyUfJbrW3kR1p
btJHQW86va3kr12TpkfYFlS9V7F2L1munbnnVNdgjlvIxmG1wsBXmid+L84G9cEl
juA1MaHigqqX36lhMLzaH/B3WGbcu0bwPr60u3WEDaEQin8Leo0hTWJccxHqk2Bv
TeEudpmNAkwJWq80jp+o1ppXcQjr7UiNFXSDOZmPutmiAeoz4Uce5T2UNBA3sdQ7
rOmi9sKghuc42EubJpon4KZNwCtteqXJVuUd1z99/5MCSi/SKot8K2tLlFIIJt/e
KXTvXic8Nfhus+odoQSpXou67QjLryECqK+dP2xKM5cGBNo94yJKU/51h8hTtFFV
K4+6vUDCTkOGE1fKawYWczJVrS9OyBXJMblvL3m8o1Pda7bhYORzD3KpUD24RMYe
NnCyNA9f69BGdVW/pehg+jIG9uXeS8oPNx5/WB5dIQdYFy+mOcTs9BQHT2IvoRxH
LFISiyj1ZmkGKf3PZ34fGeZtw62I9lb4mtsNctJDSzIU+AFUPtiS5QJwscUqFp+G
qzk1/fTgh702H1w8Q07epN+oWCfv00MikRARlxdZytVmgS/QQwsB5ql60z93E4Wd
s2EPFhSQ3XWKAeCQaHTTAryTeoRdwuYLdYVsdzt1uAkIVC0xiSin+2xZiHicXH1W
YiR93vJrHFDt0xPKpfDZP5o9A+8adFSxtMnRPMMdQlu4wcuzy3UYfIOw2YrVKsVn
Hg2D0vBkX9F37vid15GfssC/c9W9mnipXrLv22kc2i3l7t/NYpUgC13FtmQOm+Le
8jr0s+xOwqUQc2iAniTMqhRykmtN1um1KFvtq4wlSS3bj+ZDQNdW5Ju2ychVZ4j1
VFFv6WyVKjI7XceBHxdt4OKh7hJSHu7j9IIXkYrAlBJdjn4CVIkoT+xrk2akNaet
BA8szi/M59aQn0nhZu9eJGCO2UHNAcEr+P/nCC7COmMg7KLfRl+V1DAs6paN9Y0O
pfVw4CbftVTrxzSiLKBSVXpHtPR4q3f3hAGvESq5c55/RPhuqWkS/8c2qztNBppY
Wff8q4QCqcfFR0aBypryKlkKoiFcn5rWlSI5lxQYJILL7mrSZi1uNBGxE/9ZyfFE
4AWMvAWDfPu13PAACAA76D8UMb7Re1O991Wx36hkRwig6vsG+nTa1d5EN3IsWO5J
lBswiEafkO4EINys+0esN9FcWqypjb2VtTfvje7xayMQe0qrvhSXmvdDEgGC46i4
Oe1XcuiX7C/zT+zF63OnI4K0kj+IsEC5JGA9MkT8OPvELz/onfOIjxHGJVmuI5ZD
BgwboKAZIcMkoGck7OoiHyHLlCTQ6q3lsEDBUmFCcB6B7iNT9C3hnUhNkZsJ/fIn
Mi0xCfQ6Yq7vWU/yfYx5/cnYIyhSMv64e5V+agjmtbTL1LpxKyPOsU0Z2NHltQ9u
ZzFDm9GY102I6xwO1NvQlDej+QZQrSK0jx6L13H4wTELcSr1yH1Rtca34WWTaSK3
TKbqvxOhFjOEV2nAjYaO/SXXdsSiulNK/cOvrXiaqhhdc1X0A3rXROolbRDEJWa7
DIHCwiXVd956SPbpLZsqOTlEMd2NPMjccvdxllsPpaj9ycON6HGfnHn5MCOLuRf/
v614TpIxA7pHq2Iqhb4iLf0TDL0nK5A1hOqnQpGPeP/qXaMU7cIT23vwTGSpdWqi
3cIPVlOZr8eS4f3R2BPGhayyixfw2gIWcBS/6QH2S7zT8knSF8BJVrQFecyniYmc
zOX50UqPUR/ohsmDublCQ5LOtnbOkxl0E6UUjfufwgnvJbOtFxHDUn+o4xZ2GDqZ
UR7KHQ6tNl6EruM7mxBeo87N4/F2D0AAvl2qWUd0fS8h+5DAJH7bvD9l12p5e0CX
+rtwcpMiJ4zLytrXUgFKeWlfVzcNQY4uEjTeZi2sjh/1WwlbMccMixN214Y+AbP0
+JsqqPRoIxrlhVEOTT0T1EgZctf9fbXJnBdglkXY4H5PcHqMYhzCEsLxoD+fjAh7
7jYhtFxTVmUPC2w0Pdl+bYA+LOch1ZSDc3bDSb6mAjJsGCYukHnKlRZyiy623dQd
IigE84OtV7dlrfMoD1rIIBm8rVm965qq/R9Jvsmpv2PO6hETUVoWv8m4SP00GrE4
zvdarSmikHutbvbt9kT/+GcPQnli8XBVlDTLfOOeoX9l2bQCDkx5tDpfNXLJXu02
ou05yry8NA7tPEOMjPD3auuBNKRVelR58up25SCBqPhvHCmNXRS27t4s40jMTgq5
4rF/yhgWeV8jrbg87xmky1hz4o6U8usEX0drXKaKOC8Qj0tVWE8k/YxL+EOcdIkc
0HdzQKjWuHcVliAE488YjTQL42kCAeF1qH5CYrtcaDf9o3lLMLD+2o2H3j7Y+QGb
PLXsKlt0QZLuin1tTNgmkbIekgveREN9Zt5QM6MqpXm3+4In90OwBTZEoQ8Orx/X
nLRJQU1P3sq5yTF9jQYmXEAVBjF387tUA6Gvk9phQolQmpk6N9XDk4xCHwolD2/A
A1fEgfY04ThTEe3d9ZTjZb+P6yeDVnYAQtVUyDxrB6tMoUwWFaItKiDvNG147qPR
2sv1kpbsWl7J2KcjpArJ3Npgacj1NxNB9KN4aZlRJRHRzw6Nmm/GjVQv8Bd1GUtw
j9KW3aR2gpWr7Jp6c9jIOWvM8NzuFX96sNgh8Azj7TYlIoQUCsOQ2ZztaD6f3ROj
FpgVR/wcLCxxd6yEE8XpF+nOB8+VzvTo6M2gPyqpfY4dcrNS/Vn8GrjSGdav4Ur5
sC28lLDkPifzpx95H+JUqnPdXW8Ao3rpTvMZJJlHPYRgNMOL3JnWGc5xhrX8hzLT
rt5O6xQjvFpcD9MQu/igctEwS9zdjpeBi0RWZI5BFDWMTLf+kRrjpKkXkRt0bO5+
lf7a6i2YK6SJksLmlwGfC1rvn61IhX9wHLiVoGGWUk40Qwt1objPUOeiVKOdM2aF
rh2nZ+hJBA4sAOO9pDE/F3yjvEkQbfRZYoH4EG7aDcKkmovVl0qjzjSQbziZNQs0
n21VsvGehi7ndo6HP2pxlX2WYCLQOEWMv9HMNK8DaVTg7saEDIHVrLqG7OwhImwO
EJLWtNK8cKjaliJYnj356pImsegl537M8icG4JNQpdA6iZ+f+4K63buLBJiYNvq8
ZMyBoXDS+mYOYSsecVpLmMKVl5KbXWF0ZR+PVbdgsh0XizIPVgKEmQV/JNIxzDJg
1FwdNn4KRkaPsGOwRt/aOzLuD/YAEb2QFBIKts9puY2rsoeyxIQn4Q5z6fBVfFqQ
3mEoQikFP1bq6jIf+pp+nnuezsTJ5+6lkqBEvatgB+ymNYsh8ToBO7OZ47y62WuY
uVp/60TDsf7NIdywzg6iCCB2OWuwJRAhAg45S0y6QtDU2/NHfchO2vfM/jQm1GkQ
nWEzh6ZcF9l9YFizC92J6FZwtbvGiriLDwcx1/enjPgSRs4tOjtQ86Dvo4U5qiWB
V37btUiWjOzfc7LsjD4EG9G2h3BZoiqHQsQaVwsU17vuCJalNsxalA+I9oiIDFVN
Nz8nRALNDBW6EArXwUHHqVW8qU1y5sSWT/xekodB9sPq/4RXrUL+QRh1rzjPIlCZ
/27BF4sZE903JgEwZ8r/BnLt9UAvINsIPs7gDZJdJ9xnDyjb+IUiCz2FNcQnZ5Ln
nD+C++qbfmJqZDeZrd/Bl7bKN+IgWoQJxzZQgZC5xA1U+eUAF6YHPT8nKn8OnVWr
0/VxqxYBtY1WZ0VHMSFPs5ngnabErGyhZhj/8BSADgqsv6wuHDPp8kWvXA9n2dkL
8C+ZzGUa3S2lsHlqogQ7wS/BPHUH4BckwzBFVR3/u6rn4YSDm/DCymH3xVmb3aY8
VNh7ZsBNHQkmyitjga/y5dqFTCEJdgCbOAUaZe7p5PH+MoKHCGCRmjxqxLikpnhr
Y9OmBjT/kn3gLW1tWXrvSyqgSNdP/RDO64B8J5AuGYeIJdmXDR4FMp/TMbSy/7de
WSRBTvSLEwJZKheVbDvT1k5COPikhWDnNe9j13iOqW13mhUjH60RJK/Mvb63juud
A9Uklgg1OOaQ0E5i1hkb58PmS4EABSoMFB6jF7/GYKO5+UUjGVte9zVVphCbvtXl
iGxLqn5bHJvU+L+JOvq2qccEnGQMoRVexqyTl43mjUIFJtItxLkmbNcacqB3Wd/A
UBtA6lGjAmrPucUghDo3J25jF/KZiy79pyGyeiDzAuFzRDOMV+ANrzARmVW6nkwn
0aoxdrrYxVIR8KxeFonZALOz1j6zDDw36aYT8mtmG4G1pMv/rn7zmAyA7Ptpkgfs
VU9zDngM5N+IlzR8sfaxkLrjjVTvM/9Yfw0d4AxUf5OM3O5oB+gsPVKPCn2HlODD
1SYgYUWentyGOkYdFFUe98W03dvBQk6DteiiArdH6Ejqt10LCLU501CWYAefLFJe
ureRJTLIfEt7DVeZPZnVTpR22JBKMk7nemSFHzn/hbw/K3kETwGaXcmRxHg1BuhN
4VSwlFvozIGgdOeWDdigEyUa/uOMjsQwUZVwiGHCs0u/Be9T4rhQCqXKtYvODx/B
E95Px/1nslkfQ2KAAVWQi5y6K2Y1ammHWtIvGy3HvpIMiLNTDaHj/CLmAc7CSoR0
5Vxy5m2lWBf/tKRM6jGuYjqRBzL0GBLLycydEJ9hAgHorg5AVUr1EkDHHkOYQ2OF
RlhGcb+lQAg2cB0IBk5G5bezy0RPVjTGqb7Gfje44xT+FnZsz6n/cIe/dL+E69YY
JtNxbA9mlgIxhTGz5eTg8Y50mvjRHspuG3Yl6k4PpSuS0yEV/vC5MgHli/VrlDmf
nel57mjNuj2mUA3eRsX9xFr/A+gQowGw2mvbcIrkY/StSpX0TmFdwOg+rM2ER9aO
KcR2lx1PPr1uNiq3stzRMYAtcxXJiWIVW6zkE+iddOo/CjfQtlNW5m3rX6/r2uEr
8VgwAa1cfdIxLWLsZDIsl44C3ffMp6ZUAS2zMzTSMFxNYm1A0NYVqAXmYK6C+hbE
pJX7jFGTpIh9JGIMlOyABshKSHlClWZXngeHqhrDi+7eOgntKNnQODWpoVlPOkTi
ZljmXm4SyzpAXxr61kcUvqMkGQGUw89frYj00zCY4HUL8RdummFj/NbiifrFW6+w
EELez+y1zcBzTLF9Yu4E7TEUPZpARkK9gP7OLau2VfoHWx92bpxQC1s2VxXjPIDj
c9ub18xgvvLun4byzjclrr8wJtGUxm4L2ZtEEoxcVa9GjsyB63Ruf7osXefvXKOO
mhj86IXLAxsMi9Fk1u2VPttfkoQnYSnk7Cg3bGDZiId/RT5pR8/j/g7OzYpwcAJ9
0/UWXoami6Q9PyjcOBd+9WpLSaiCWPHYDSHq+Gm7CCX1nfujNwAQlufM29JdrZ8Q
T47px6en4f+jkKF6uDrMRIjWOVBbhOGWG4kHjh+besvGNLgl00TSVZv9XPAR7fSw
GVnfG03DL32A0IyN1UDeCI+g7lmMm2BPIyusk4hXWdQ2fsVdvELEeHgFTrmf00TM
8tKq1iAgU+xn9uW0ULE4ApA1DjhBRzhaqvO0cucjEuJYUg7W3LyPpwAkFyFPIvwA
ucgx62hedrFPoXu9DzKSyCiKD5hOhkV41wfrpFB+yPGnqBWrw43Eo8fNczhE3oJk
8W0Bnd0EUZ7GupHg94lx0Km0RVXVUJs8AohyKb0YddRFyO6Hign9dCMUeNMmvG8g
m2ljcyvBUZSllwo1qphAHttOvIbePT07clrqRl7E7gF1maGW5OKlVXKxMQHTxHrK
89T6xf9LtZEdcjpfHKuXJ/EKwE0GJ7R6HWC68rbxSzOW7Aj/uTsYXm9cbEMGgDDH
Re8JNbUjBkjD+EmyyHnEocQ/OenAFHh8DFlEkMRqoAMVD0XV5VhL2xz0GSsnmCwB
JZCL1E48OTL+nlb6yclBDVHD4b9Gij+N5gGUdW3JwqXXBLdval0WzuYA2INgcuER
9qQT2h6aMpPey4DZ5hHE8XGZaURjoYWOFo28BBQ0Ypl5uIxujCHxgjaIjC0E7jrT
tfod9inOuHSfrLdaEdR56adP9TNAWEiz2/NUavEQ06DM3Q10Vys7fC6taTaxp+ZO
003wK5BiOva3V1cTcWg41+9TCt3TiR8Fj/zT5HqmTqCgAaKRwOdr9BNuJrxy4o+9
K6D8mZKtOiMpvSxH88LGk0lrN+3yhyfLg/uMoExB8u8weqBxWqzJvKU72NSAkZmQ
C6Qv6UtM7g6slFcTR2HDTiI7b9yS5wbKXU1lI5F2jrZF63r9aHJg7CKz/Jl6g9jY
0sxHYAXuCrD+RbsKZLt6zH8hBUjbT0AI769/I8FaYDDbSvQFhgAQ/ED7vapAakxK
buhYlzeMaSJO6yHIlmCzoPv7DHc0sD/3HaUQq2+/ty8Mwb+/skhixZOGWiAyawm0
4Snl/zQbtVahNbO9iFT1d6+diK4h9NNEUZX90Mo7TL29vcZyUx4K8N2yO81WGavE
Ubh02Gq+m7RyQtBzUwNpcTFdZfNDw6XlsFVC+16v8655wbPvSXTa+oybxW0M5Mm5
KPvcCg8PriKhM6cm3p0yLDKa/36ywSuJO8R4NYlbqR+Ng3WLdLxa6Ijjyh8DJNRs
8/ZtwI9flxDl2AM36F8KcoqTkaB+Ji0Yy0ZECQ8psdbQc1sRLZuzv8K0x5CDakJ5
8EQ80TnLkCSoLF2pqjWyhHclbNqHm6kim9mgF66mHu0ks8+d5jGDpaIxqxpPce5K
zDqUqXzvxdGLGEK9fcMeEVrj7OuKcoY/NWx2l6MoGXp7k9IqjsnjfuakK9Gd384u
bN+wG35HXBl+Xz4m1rYAt2C1/cqEYnP5xFhd6R16/9CN9w5AZlZi+juYVZnFhlJo
L4fZ/qrVnzEGhjXAkIM1PJibs+eCChFBEoLkcWzt+o+6qxPrSDIacnUXE4Q6Rppa
CjqWN7Ioey9egqI3JJIPURdD3IkmPAVf53G9pfflxaER2h9MO9ttYl8vrGXZ6dZM
plcYD51T7rLux+8+zvxrHO+M+7xMZN1GV5TFnOi6pf0A3XBLrvxAIuApIiX65q2r
bgvN98B+cjWJD9fBpsE+l9SFtdsVhYhEuHR7J/tDGU7t8MntKxX8jz/T6ddr0qpJ
J3QLfzomcYcKncE1I0V5Ou6SH6+rNEZQdbGDviygySVZMpRA6XQ6JJpQ+cv2OU55
hMhFikGOEBBPuwMnNdatLXEGi2+pO47ueirKn6xhAUYalabmzyWhRlbhWV30cooC
/KZQFnjgmf3HYl6vQ6/JsWd64ekLQjjBKullW8NTXTi+05/msNGl2HzMFBT55QrU
Ti2+tHSlXycxgxAnpGyOJ7g/hdFMBcAO3p8tQK3364rcxOkE7jiN2z+EQj2Qo4bd
lUJlTrRzezSQwyIHvkEEc9ZRBMVZs9pjOTj/yRdXg7s7S7okkcoRKodJyj0ScbYD
au5igAyWMqYF/8eSmfxiGEWCFYPb0sySv0MS05SdiWEtFez9ZPyMO9R51SRf6Uzz
NmwIBG1jQlxEX9Z6f9A4/QZ6J2i37lDuf7O+d5pDi9lubQCLrqN+3Z6gDnJTBuBU
231JTV9ji429+fUbcimenLJc1U2jraV++MXRcw6OPW/6lDFt9pMQLCEXJIYQEs2Y
00hHiKEBgJHP9m7pFaZEoQRLX/sVqs65ECaAFJ9FT4cjTivOPZ0DL9HOt2pU7dBi
D0dSVglUUzVGUTzBla7lHajnA79SFh3vXVpOGsKMf5raY/MDyqxsF1xY1zKOtjyK
x2kk5N9Jq8/ML9mhoXfX0CS9HslXNFr8SILSOODoS8GNPxcmnq/AWawDsldEVPVp
ykBevmKMuQhqHklvdawYLkqbRyI25e8LdvhyJ1go7irXm2+eBXVzb+TJwZ5lM706
6bTKRaZ8a7UHlHuKC/fmDIgARkgma2mOVeaBM99ixTvkgwDh3ImegQy4kC6mj9Yg
V+O4dDO3ML0jDmFqmy0KhGYKNnEFvQUsER1S9NlyrgG6InFyCJ2Iam/HVeO/yWfi
jELb9Ccv2s+md6t7bGxIcr4m4/1raRpjiV0vPVIENerZFsHei7vezTSLBylebpgm
2ZBH32TV7t7pTo1v9OoUIrC0LRiiwoRaohgXNG3iP0o=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UU5f8Bto8FbjKrbPzds0x9GfOqD81dEa5FZNdx0APjRBEaRhzsmfE/W/dv3PZjuq
G/BK/eVnPKJB3hHnDwzJrZTisfKSeSPXnkg+udu2faFTd3xW/0muLl/ehPoG0/UE
Zmw4tY6o1RLEF+sxNqM0eQ+AlgdMianwh7QsZQWYyrekBgAbA50sl2i/t1HBPY4Y
GKbnrDDAIJT7mtFPeBbbPmq8LQA1dYdEn9DuuhYyd+TSYp1NZw+A47j2UnAkK53Q
anKHWE/CQ9DwK58fEU1/5SfsFgAAEWKNdT2XXNY2VSmty1sPRZ50fXBOht1H5kvr
ArtBuxV5ck9NXW9q2C6f7A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9232 )
`pragma protect data_block
2rl6HYFAkhvMXUQl0XnHErJX7rAGF+EjqvGK/j2Wu7MZq1VJz+uk/Iq6ivNzmqMI
cZ5xiBPaXFDq2Cekoz5YU+njVVhZyI0zb03t1hl41YllePsdFITazHAnjudHB+mY
PavGzeMIVuFRBG7b2MY4prcbQsBeMv8VEYcZZMqXNxS4BypQQRvWAQbpIwZ66+yB
3mLXFBhABPkGkEOYma/wS3UYcmSsBjjOydhe8MKOBcrsTR27skbK6lmc3L0pOEwm
diXMK6cNFpnlhVMyGh+x7LgbIIPTqyhTNdQWMG934y38xNTr6MzBfPCeT/KkteED
+0sXUANsOf7BsJMRBVo3lWGz29A1dOGZHpeVO6FWt8QjWrybdBmWSONH/X6vRU9l
Yzw4Qp4HWiWesnF1yA0RDSmi5NER3C+URkZLpLak3onJABthSjVc1ThArO4/v9Lw
xeW5blUfnCZ3uaSfwZCYMgT2bfh2mMSBfDA6W5vH4RxQiiTOrQaT0x+ACEqGuHrc
xI1Zh+Gh/NIeu38eq6jMfbb7QQXy2TyCXZsAvyHsRFq10EUWz+XbmjjtTT+0BrPO
sRLvdH4AT9trVgEzcCgCgDjZOo5+0GipqC2I0oCfLoUvJ5mrI94kIdhRiXdmMQrQ
3Hr25D9KCiJh/HZ9KdbOt/UxK/5scpxeJVDH3BV/atpt8I7HVkc4nQogzyssgURT
uDe5mqr8ouYLEmeFBgeSZAKury/MYEFeCD7he+bbVnBjcgZk9KErnzjr7hWpJv8y
maEiwQrMUbA/VdiOwL8pgHIIWgMq0raDOQ1lQm6m7zRtDByp3bmBc+Zub1kfYcZi
DM9ClVVDUjCpXaB7YjMThWAHvvVTu4lVNulnpAiuqf27bfcSMEWFfz7MLHMHYbOG
p/7x24mRlmMA2IV9kBhGkXgbvFFLCzZAn/H1HuSziMaNcwB7LQ/XKmz1ThXBKYc4
iI3uEx8S0t0wfmNMQ2SqvT60bv9q2AD5Ct5Ph5ERu7oy6rkNDbL0JZbPb04kI6l7
BQfg8cfwbFZEwUdmIeV8cU3Uc309zlDVin0bvcIbcPFGuE33pITnftDgEJ8hZE2p
LLF4pE/9dDIYJsye4+afVqPq0YZDLQEDQ0UXCgqkpZWiVczZnB9u9zf65g+MKG+T
XGVxT+6QzYF2h65pCeXo9IhoVS3hMCFYBray2qNxv6xebUUT935kHNtzp5kBBr7O
XfTHj6QR+4lzEGRCnlI4upSkligryDF4XDqee/1L4Ef7Z+NbH57Tnolw2QQG8THH
JnQacngYJ8s8Q9TKpUaIhc9AUzwwSb74mveoyPY2+Bj+/mn7BIGQawJc66XNR5f8
1yrvW7iKL1EKGDtYeRYNemyI/1KEzy5p02XSTjlcRh41oapdTvZuGWBYzQgqKEvL
9eYF8xW5VAVgoucq0jGcFvmdcZA7qmShwk1dQF/NVsnzHHJbGVpERDX+0CWsl8k3
3cybsEKu4Nb1i0IWtw2nGz2bZebtlitngGu87MSCDevLy2jOF9oliMIYw/v6Qd5M
5ZdjjgLr9lPmGapySkvjpQuWv5PVWVp6mIRAvbF8/sFwLn7ZGsXcEKkqRg4tbf3z
UVxmloau2ouxrji69+24521Rx/CZWoFI1HwO7CG+dLmkKTUS3srPMWUXbE7D9ceN
i2IVFuem6jwLtyfQYNPk+BlpnoyAxuTNY6kMsPrtGyOgezzBuG9VOMR+fDvkwUOo
a+eqCXIQYthlPuleEToKnVJvLhLSzxrgceGZZqfkLPAfQiBiBjsN9LKly1Erkx4V
HmNRPAjcqAcUUFUWsUyM7GJW2/1Uv1NqX1aptwfs8T8tZfoSGjtUM/lWllOgcyLY
1pAQVQdPP6pWwbqjfo34A1KgxTefBJaIUaGxbRBiW0D8aVe5NN9m4SIkeTnmxnqs
byz8HCZrYODh8pnG/fXIMjP5jGVQpFjVWpbuTilVPDucdwZfhxPy6RokpyJ95Qvi
e/T2pibaDr1QGM3Xgf9vf3Gc6e/s5z9oDvAnlijWPDezmisLyBUaIKSHdIx2YWbX
snbxyexB1y/SSdVODoliBHrfxWOl5MfOnpMGrcxHnLAJ7N5l4GF77PcssA4nm9a4
zL5N+7PAlNuvwq8w+UDYMqLmBVfB6+L4IQs6itOsw6YfgW3OmQlF6OVMgZ3fY+hy
waRGnxR1nCQ53YCrUN5/todttAt1hxY2BZKZwU/5/wRYMZUUCBa1u09gHk8I88ZA
QbXpu07jZlyhuWPhEO63Uy7VX00E0KRZliX9FkteqRvmCzmzT/mDAy8gh1LKqaeE
rZAEVRsgvlLK4YBHQwohpFCHeCsupSSIGiWzTo8TETPBVJm+TkQ5f4lmOZZlDnbg
nmoiBOZ57NnN3qHrPuQyxczsdHh1t1cLRIVQ8yixw5MLpsue4zVisdSSTqMXvZ5Q
zSRPpk6tG/o192wYAn22SOmXHHwjeo5N98zoQ/FDmfjPl4kWJ8k0LYekBHVCj+Hq
lnukfSD1f6SwOkwSgPonkl+P2emhnNhy3R8QV7nDGUlpd123hWrgIqPYwaEN6yBi
dW36q3Vl46mWfwOPbHiOg+SR/ppCIoV52DvVL37aZHNDktirbbqxsmflkB26s/Ij
WnB2grPrmUYJIOpKEFqmNM+r3TkPT3i33GZkWbtN2btfh8QChRIslIKig4Hp3Lwa
wkySwGgXKeXxqF55/tsf6jkFLXDvPdNN9FGArvwP9RkLV9Tr25oAZjnCEQpMPFeJ
dA66Hqx3Oh79OQhyRp31Zs2iB+88wj6iazI1gsHGxKdOPsMBMnGpVKJ1ImVAwvNQ
/RTr6IBn+cSPOoss27Pg2dvvLqMhHqkE+jiNb4SHHw+cz/qA8XC5uQZj8Y3CCnre
vm7cdosRYh2ChkEoyllggx6v+6fAkSsQ5ofh9a6F6VNmOaDkttt/yPdFhJOCqK2F
e6zLwow039Bn9/6Ob82Dcnun2kdwLPo2LphmjJwCa32tgCgDi56aUIbbOyGMcUBe
vbsMNL6fIR9iX6tPC0DLi5pdXJOkH2v/9sJS7SyT2nxtA30aaqz/dd+BTUvju46e
P/MNDevt23osMEayoa73E9XDHt0h9S6ALNi/npA3isfKmAlsrdzvo0XIdoBP9Ekz
6AmHclVAEv2L8lw+ycKKWONVRbKvHEoHFX3UTwIKPIf0iLyLZIEVCnNwgPnv6D6E
Tn8DMFRfVcqw9GNq0E2D8CH4jr0X5bqcfiHKnAFomJm9WWvIWOvuAKkhuSTGnlea
pDUoxAyw1MyQj33E2KE0lc8Mq06WThN08/6kZApw6U9uQXBIs+DuIRwnToGrtU/m
wc84+qRWZ4f422cha1bHoS3lIOaRUD/C7stCRCM+nGgPr0A38nWqSlVXzy33TOLP
qQtLJvAejQnr3rtFw9OlMSuBlk0c9H0w+JIt8yeEuGVBH5Okev7E3z9mNO9BQwvu
vMT4mWfIm75ZiFuMXZFKdHfHT+L1vdzYo5wMO+hpluVEX9B3ykJJIetBpYN7YNuq
y8LyHnpuGc3bQMVc62r4+miHqOCTCIqkpTLP35d7CXyO9EwkXPGtbfz/ViipEIHF
cw5K7X3aeSgB8zAze6+16wTAE1N4euVaw24N9oIIzsHF99XA7Lo8UsIwQiUxBUYZ
7pcYTS0wKC8ViNysGyi0S/yvi9Yrfcdd93pBShTjJF8hgwhZ7ISddc/czo9fRljR
PprLDc6ajU3u9k7r8fNxxc49jWkYZmjwQmLUYLDLdw1kbVP9amaSX9eEtxH4mj/w
U3uU6ENAnZgqgLT/QQdM9zwnJ3h/uovSbJNwg0J4xUusxJ9uqUClOzqTolIKrU6x
CUyxUU2wVNLyrqJS7ykNdHqKFLxmwNJsKy2Di55AbaUm9aEPMMWQd+jy/S1pPEye
rhD2GNhrJJsuz9k753uIYpBOTQN/MzEDy3dpvfG2XKomECa/7RTPGD2WepgTSHWg
LeGGHaYpFg+1Ujtv7v6sDLcM79QTVl2aku5huxVel7eaOOUeJNA5L2hd9sVFe7iJ
yAQ/U50J3okeqjOz2nv5PQTaDP1hKALwc8zvCbtwYP9VEwiL/xuhvzshQk4SOuYH
A6UplG6wHI9Ozt2pDExBJOPcgr3PW8Ul7SEbZr2ei2HWqED0O4pz4NjKUDxH2KMz
Ui89S94Ti9WgsmLCkKeRSwU2UwwBCm+oPKx9xujjitrgC+1ghwXSNj7NPOW3ucOU
fGpIvET69+Cw7Zp0BiuyWxVgUNFHWDZ2xlZWjY1VbUQLJxhVzTiqNeeXKpGiaDjI
pm/xFcS11IPekS9tm0+tfsX8f9tgG9KFLD9L5mH67k8i0gEtpaWbhIlkEFNrVrsQ
rJUaJfazs6Sm1/jgXk4dsszTpm8M053sWY5oR8sNu55bhs8r1pqbV0RWTX1xouNU
PoyVTV2tp2ynsmVPZkNExavDi2YQr62KIZtuG8Sio+mB0P6adkCubrqyDZL2v6w5
O4Q+ro9sk7YSvXkxtI/36RDW2jJhRsudao7nUjyTN25QPdHL5LPLPdN5Y8mQ4g83
z3tMIZjuX+y7B0djIxKZ1AdzUzq1xKpyNqVl26Dp7IHWYmkM66P5EmP9IOxffiwn
3FrimTwxJI2QNg0t0pZoOOgAfs1znSTXr4EF/GzTKqNZZknoacoBUdabwJWxbg86
gxZvJ67kmE9FrdYxSfU1uMOe7TJ1dUgJs5xAC2fg1OpHrlB2JpZjOd8vqZg/brt3
dGqz/NnyaczqfyXhSfxux0QMd3DKbXcb9v7TLDfoqAg1XV0/uOsCvfw8TxyGszCT
MAXV/Ilvs0M9+A4ZEYwDSaOW6wIayGLavDMGe4f/CO38abB7AqxybgRlH72Qj7Jr
uwNilK+qiqhbqMmXAodVrIjxOkJ82erRfuyjVjtAIAH46c2cAD7MX7exNSrFoa/d
BgvCnEW1eEgtSWWjzZc3F08OI2KKDqgBGZSQ/SxPZWSali+KY+cQoQ3kXZvVMX3E
0knTHh1MFANwzyVRSgbaYfJReDBKFWh6iiuMoqWxIVJvsKp6AMc4s+7Ewb/kQEzn
14Ai01f0DX6pWzjDt7Z8tv11+Q9hGzVud/OiF+k7utd7NnmzDWGujJuZXLPudVxH
peXgIlkNIBwijiBcNcnAALI1dFmJmuWIuUIQcfCgv/+pxuusUh94PjzezOctZKCS
i7o69P9Oox0NejiTnWPaNJM1e5O+B2/NAm0J8pKpi4v4fr216bxJP1qYoMFO54OG
KOLWm/WHFVeWBTbzo59In3UIDHH3BS5YFsDFSbbW05IRo5WLYlBDQ1X5QjGq3CFX
CI/YWdbncp+OzDOxNkmIia1SmSI2FGq7lw5wR7UCuS5JFijPquKwt8Q4v1zmPPqQ
F90DX9+eoAGtikF1MmSx0YzTROU14pcHvMlfUvDKGuyipFPoMMxebtwAm4LbHmKf
KLjpm3FLBCBiSFb7xiVkLLJ6rpS8mgpYGxzVhDZfbtok4TbtO5CdsnAIDHijIM2x
Jtn01MMjVrdmEN6OMTNABnmkp0W8W49PBImB/j68YTYXu0y7nsv4I32Q0+nDPcqG
0HEMZyBO08vqpIqBzMvdvc6QRXD+eOZMylDnh8GGnJb+48o3WOwYLNCsZWP/coZ4
jPYE2TMxmWlRfGeaFy5mgeVgMDrRLC5iVYnbU7jZhjclOD6N7+3jTMirXfw7sNGv
Dkfl0AwsydDb8Fdks8ebslvQURQS8FuCX3BzVQw+7mev5cM2XfKoHsKUlqfvxxJH
Y6WCEREHp0g3rrWDntoyCUdUg9EzgodEaf+cZXqMaAfrS1qw25EjR/yHHNWXwa98
CY1lDAT4Fhs0ZVg0igVvrzl3Yx3bTMOGw6nQJCPSRExuQ6qa5flQitvOq0Tp6F+K
dU8wK/JndIeMW9FKAnB2XBmqC6zzAsTPTF5oPpNVF5FkKwD817n8N0ILfyclqMJI
LrKqBxPfFSjoiyaxeUw7/DwRyKnoJZxnQtUIKbEwLVdle2o1rc8+O750lh7Anq1B
Nb+PSfa91qnUA5802YIV2lG+sCqgzPqnUurWzuVCDSYWoRF+k7T813qi2b2thtBJ
fKcaocNyl1w6gyIcWq6VwuMKV10dgcny/+t0do032IDtJ686HZzP9md4IGH/b6wn
XkH83ahcj830kp6s8Qd3Rdd/C0JYYlZ3mIbCPP1UHPzE/HEt6B7gp31AA+DRvW3V
UqUJ0H6CO99bjtgY2pJeHDZ96P3g/OLJtLMkUh8fiTDb8Kor5ccGR9tgtfijBNvU
YsBPal3gDCFHn0ugs2fA8f+yMqtOhkEUOYW+IdColNg0nfvET38lXthFPuxLNsBM
K0oiNq2RnI7gAJHaJFCCrjWLWlM5oWZcdSsGzhf359Bb1scvaXsr6vVLJN75S+w7
i2T8282ehanPilJYqtM6WR/yeJiupRbtt2FDyQ+R/zJwpEnQMLH+0JHtjEZOVKrO
vATIW0a7+7baMNq1qofCkCk5L02ciAv+Sd8XZIq4/jz6Ziw98kVgOQzfyIAT9MZ0
eSrfjqTDN2b2LB/G8BV+Nyz08IqehSSIE5FJTwYwwjOR7C+FG5J8lJFsRv6c4xu4
NGcVCtPTiIUK5AiZ5d+UNc5C4ly7BweA9G9fWUNtJA47m2Uqt/a/Hv1jwrrmGk/0
CXGAsoNyjHZQlIHejUPgINYizERCQrN2GJeBBaFJYHjCuYEOTvI7k2OhmKVraE2D
nArMkwOqpa6oNmJMAZhBFjf21bRgPQHnvr6+O3v+KFNxmGDw3kKh8k2mLfsBf2aL
SBeUPR0895w+lx6OC6qfEKzwlo1DLa6JmJygmY/XFY2aspucWfyIxxfiuAtcIMMr
1HmJDX9P3FnuE46D8GqrYielgZrQRTXDmGwVQt6qrB+xZQ/MQH2JbUvQCVtiXEHf
n0gcaqjKFyPj/A4ijQB4y608oFUNMI1DWAggfXROpNzUSsoD8PvOr/VBhP0ljaMP
OASIA6g+R9oOHKBP2Nsh0RBxPcJKqALp4p4y5GmoiTOIwZ2Cf1k1PJb4ngGgwDzC
X8CFgfvU4ClzYmEJ1/fQX/7gGnyxjrhXfwku8FPkWkmy+GABPJKhiSOaVHlIn+8G
QYrcjFDCQKEbkCDohK6mYN/2PdXTHv/r/CY9MjbPXAcQUDh+maDtco+4PqvTquP+
12hdeli37GveP+wzg1zvPkQQdqdUq+FEemNUXw7hVsIzUi5IazFDa1SOBqwp9Ngd
NpDovpgILfSQOtsy+p33UeId3f8RrTXSzq6Pex1MhI/WaC3gbC2LEDtbd6Sauaxu
ffGLCJa2UaTS2JTpZ8t/xllo9+8EN0PabvIhiBk3eDyLwtRKKtZVsI55+CTfiGu4
MDV4zn7UKmmu9OCNZureEyBlIbP8Ir7tYthw7a8R8PqgIirpeHiA8vVOVZIxYbfv
W0mx06U48yCXW6UPYnRDfuE7He1oTmZpeb3S+a59pkDFSyGVQvSbNT1OXybCotsw
59NzPUxhUsBntbbWqmvsB4dnt2YBpuXUVxkydcDy8En0i5KvH0yzeqrNr8Kmyhxn
UYOi23yVbNkUfttod9iJq4pIVwqDA7q7N+eBepYdO/6PKf410x7y+JJrAaq2t9jM
Q7DS8jkica8VTuumNN4qrbs1UV+HfUYDIhG8R2Qgd/VKMPOp2EreEVywB4DnBv3s
g8DykIvup6rAGIGEJN6sXG7AzzjNdL+W3CI/h2SVCaB0/L5rrEddfM+DJkp8Eq8F
zrvOHTcGfs7qQQ3QkG8lZykbik1+E0ylZx5eVRleV3AS9rkCJZ/XcnEVvEUJufbc
oISPA8Rk4QMtCZC2tR8hLjhUWhxa8WOeOhG8RHemiRFmLm31PzVKraqEA9H/DKS6
7lnNBmE2tuqEDIwZdp3rhBWe76FyxGHu4N3QaAJaeg1YJ1aDlMjM4pPKWr7kUOI6
x47o58TxtFdopb6p4SIOmmiiwpNIFmyTCWq8Sxc8Q55okOFbP175XyM83ajFZeEo
eMClYDB6i8oS8sa3foVdMAq6ESIMpYrwIBRWVGCbh20mtbpptGae3r5rhcegXaj/
FBV0zWphJKf/ST9TvfAKqKq8uFpm5dsbQCEZkqz16D2wbVPADqTH9h9g+lsdMysD
hgBngyNHA8PCIiPgrbuWeHnnfya+WT0NEEDzqcTrIJDA22sppW0l/wCAT5B8zHBK
L8v2fHZBVK8NWJK10EKM0OuxRH3YqZmomCG5GO4xQ8ThjjIhCWvQRdYpMf45dgTC
5bVtrFbWpGeLkEmJk1R6g5v7rbovPl9Miu6CMep1ISzB47GqhwtLSC8yvHglabxd
WbRB1NVPts7wFv7tO1FTbLjvpUqe07k+rexZarIjCOCil+mARLnouwgwseSrkKEs
YfhJ9LtSiUuPI28NsBnKaQNTr83frC9Q3B+AKrVofFTmsOhFNqgwPa1wri1xTfv+
QORa3g1Ulh22uLotUaLAcFWtUreMFWIgTajF4/vX6UZK5UCPOQb3jvXsY6bScitc
pDuxnI4AvTTh/doUJ2ldi8xdKhoz4yObVuGjPKPZRog14OzN4FNEye583YadQ14H
VK61hUTeFn/NBhZNC62Cth0kCRoE7cf4pc79wTNyAnQ17CmYphGkSrPE4B7dVXRG
XvnTLf+RE1pk7zpy5Qa2YbnDqnCEq9Od/jX+FzrR4fxEdimpUJbQ9TisEUkczPTt
g/+sGK9axK2SN+MZi3zRmBbfAQ1XCJjkxK2WvAvtC12rfZpJUtDC4CiDr3otH6xH
JrzMOoP97BiLJQayApPLE3JdTq5aA8rySaMgbdGrC+QPAet0fTIPBrIIdOCNstOZ
o7gujS18IDixqp13HyPvuKVzPOhAWDzLclfsMMp6oPnGXhH+byi5z+f/YmE2IE1f
aivzoG535ybPjn+jvaQ1VjOUMopsfYvqiDbm38NmzMNw2nO9pEi5fUYaWVJCae9A
3PsCTkqgglMnini7T6AcdF6kLZn70dt24/gNchxJn7JTnkJmqv/ci37AR+ifGtVo
67Fk0K2nQA+ecqhHvbTwj9RvlSJ6uMFY046hc0KCccHSTSrCY/+a3wylUPxvSCqd
vtWoNpMrsuPHsM2ep8E9UYnoHF44MIA7U9bc1wS3GSq6Bc52etmlhWLHa/Jth3+i
7Ch4rm/6h757v9aIjGym7bMZH6xhKRMX/RUYqR1p0F3XOLpkTR6ix4loK9mf9rXs
8w2UOnrDaHb7y4hHpR+TolAyWFVSFdwh0OFDaEa8mNivrTBmzefIExv+Pmk5E7Y5
xTdnoKrDdmOLABNPypumMxBg2zY+vGs/rKILqGctNwklYPXbT+D7C3fzX8Bir9ay
LDGDSj266BwzeHWIldv9Ne83txaE8tUt5EBubc3xR1bZ6NbQFgQQqGux8ztIWRdO
Covj3ujjD4KGGefpbfq9iel3cmQO4QmY3VQ8bfLrDk0d2YQEIAZDyxPK1iLYUNcR
0pKQ+3GqeL3UriP80CO8M/rtFAOaa/eA39e7eXp+HnRg68Lrp/x7/9+R//h5q35c
fErrH2IsJf4zcg2Dg5Rb87pQMz89oX0K63MOvNQqEUXbmZ5v6Y7gjfrQ5MS339jH
DIEZy3qfrQ/ueqJ+zqby2v9ZY5ulRnvp9Vd0T6PQJrLX3CN01N4zPtybZmH7Q5EU
eoCcYZCs3Ka2kyizJ6plLacoAPSBKy4FgI7EC8B0kM1bNVEunenLJXMABmzR2AiE
6CwGer5Zhok2reYz/q894vPF3n2J2iK2jyAsXcwF/H4LtvEL2HxS8Cyw3lWS6d0l
8Vm65SiELOqfPDIVzc8yac/HRVLN70BBFYnwlxWOKjqZqVjC3nrDe+UcVJ5h5zaI
EPRnZBVtcxq0OPqQDlg51YOqczQ9ba3QCGZgiL32sPl+hK1iW4hZjd1/mm2FCfdy
lh47I5a6c+ZCCyYaSod3FzqXfYbRf/e29+iZg6n2Od51muP8o8PkWd5pUp1FOsz2
tZfprop8oWdVIZjXv0b40tr+ipHH/8S2sVNSqe7q9Po51l9mGR9s5CdL4Dc+Q8qk
I0HuBteUManogL5h24BPfcLB+/82N4yFTNQJ5qAAX0xOG1AonPL3gE627YkSOZGp
Trh+v2JIPsCLqzdBlZcT76VozMgMI8z/NeBWXrtFFiNcDKZ+dNDMyrsyUi8EqE9a
qbM2pcYEiMME4fOUq85h4Jx5/Eq8N4HtBU8lrpigv03N1Lv9AFJlM15lrxltaIdQ
QvJR3NSZ1LU1Z8v5RyF01ceGUkL6C5gXEOjJ7q7DV4tzNmBoNpYWfJZTCdJltRis
Ub6JTv9dGPagGjsH4pIlSgUEIV3puBEHlmYtQzDfP4e566hJRJI5t2PrjeaMLVFO
a4frcNEbHQpAwmmGkYe2KpJEpQBVzRHPz4+dfPt3dW+kxWsVpnClDyFJp031bP3W
3JoZSDUJLCKUrc2rz+q2Fs0XRdFGw2aBLx7vNGMsBNo5KTOAoLSkwTks2IJvvLN1
XhPwie6rJYnT7syxR6fjqb5W9YyAKBJPy3jajSlCqRTXOAHpt4+qI6/aVOVXy5W9
WA9PndGx7JQT4GMInYOHFJpFMeyv7coVs2yCsok5X0T5ZunfMlym79dXCjacMkku
kX4Mwa1D7e5O8fKEr/TE7F1w63paKk1nIyefJlyT90EoXynH9lnXbybzg8XAofzG
3dwJE4ltBb+4CG4qyZuFb5wv0isWK7WCAXCgPbt0D8ayaGqyK1jib/vHG8la9WGx
w0l6cRtcsujXqThvSfvxz3waQMU+1fhBEyHGaV0MSfgOOKZMF2uLj9twWijT9Qqi
WDbvNOobIUas6wIWShiC9XdPhUtUr+scAYXrQUtp3kd0BEvdYShxcQAaPMy1SwCT
0QeJrOaUAdPWpxldUzY9gveTuxvzjbtWr23CToac5P/DXW79kqZD+01jS4+NBwbP
av2i8VGI4yKAt0Whtkm6NqalQE2SJf2Iyq9lKor8sa9dYwv+hYPjGon/HK1PzO9u
kT0nAG7KdmPeYonrqoqhwiQ8GUFXLCH7gMc/bfaSt6pJo9g966VfkwT65YMl9NGG
r7mD8M4oCXpTuugTjVZVuJ1d62+UuuISoWZgSLDy3cuwchuBkNdM/+aaDofCgXjv
CV+g8SPWBKBfxW2D1SAADI96bAPH6rNJ/9I2010XSLaLStFV8jF8SGZjVanrgHh6
Pu0zAo4vDjt0+qevM1WUPayKrocHK9t3mmOtUwvjeVQ9SW6PpZN9XPZ5/EuHfCDQ
uzqLvkqIzLAKE1+XvPf8Bk514HDwIMmEcPfCENmLuAz1qV1kBWY5BUfKiSOeCapO
dgKl9WLOhAE8RWaQLMOdTqHOCFVQMwBk/CvIC4YB5S/JOrVWrO4cF/4db11v31tR
rKcUEYdhbhDO8sPmByRPpe+/wyeyDtFOjvUPrWyty4J1rhX8yYKsobhu4IpeWLX4
mIiw9GAiJnk4wv7ZpuIQchcTq4+KkRQNcFTOBS6sj6oc8R+2/91kwdUnmMb7MJU7
MjBelkV7plG1d52i0JGd7j0/qqXyKbyOeGcEy4FbW7TEjafIjPmVN1ScRTf43DiJ
SEW5seVrOkdZU0u7X6a4lwmGSFL/DLvLnm39xndqsE7en7VktPVdocG02XFQTF9V
zbUhwImYnZAm9Rna5BU4U5bZyYmlYT+OiKEyE1/kpEq71eANkV+gdIC4dRVCTi6I
Sdk0ikaoo5F738tmWmJfNmJQT+iq/PHPllZ+z4BEWY9L+U+qh6Kwnss6FOkzk/w6
J9S8xf7LoqC++JZDuPM5Tsq2e3w9qfRuffShB0tGTeCzt06gxuXiBmwCe3Pyoc06
5x0YqOuTfhih0IQRSBW+70PEjFxoOjTG9i8/nRHa/Hk1L5T/B/WAIxuh8YZjjg8V
vmTbCMsNYnZskOd332lQ1W3l0IDlvtSLAcyz+EGX4Hp8ytVF83fi88IAtlTVdycH
l3OQvJF97o1mqQO+RkiEghksvIEz9zO/TD69dKHm3T04tm5Q4b/bcBpODIhgCadH
teMkklnFR0kH0DMAx6Ffol/XdjkNLv3bpqRO7SxOguIiGWdK7XhLlX35+9t4q+9B
kbAMy+YgCP6wLQbgHxJ9v/1+PIjyFDRIRlmotAYYCOcsM0YQ4bSt/QwAWSYfpZWr
LjXYJ4tOks6fdChLzsgAq/9UinCq9rBGcTeeglIUXmRl0kVzAy/fexi/vG5I8kZK
8PDVV9KfUkYJVFjXiR3kl//gHLrFO4Xd5xGnvFA/EX/4iutroJd0qb+M+Yn8zLZ8
KK+j+vtqZ7my6NxrpTFuhw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
YeDJJQ3+0pvrtGbaYamee78SmKsdmG2kPUmDDwR9LfNbfsD2cxTy4UB7SVh4GppG
Ot81wojXnPSqFBzRWaRM4bJBN3EZdD3Zw2IoDHVwEgcwgXPpyKLsD68Y3S5cMaq5
3bnhSoxb4UvlG1uzBhsDPeWk7upokblyp2AGSRIDn8HEIfQyOXvXGRSjFWfEQuET
DNIauWrZM/ia8baEiS+0E0M7/aGdR0ng2m0OHUrs2U9JEpsY+WLL3a1Y+aolH3A7
L2kGfcJJ4qS/H/7mErYKpBnpAXDDgpXASLiagIT6Bf05zOc1t6E6vKRyfySVLCQP
HxgnVOggmS2niewyJssZUw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 15248 )
`pragma protect data_block
SQd/rWNXEdiOzgivB3vbU7BBEH9JlLZz28idVvpKv0Vz7dFl4ZcioBiXH1uURQuk
/SS3+CD/FH/HavFrQgkpv/zBVm9Mdx0Y7LjRmgSRIy1Vt6zoLXu+GnDviuQG6ZA9
DwWki+c4F/CGOOAClmWFrw/OlVsKyfJo+1/8puCuWXt2tBR553gLLbaxp0f8joND
z3cpnUIT9U6kE2XWiAuPNKDxVZRiVOD/ucHSCHjpOAdvGz6b4RFoalAs3oL1Plaj
iRhZPPV/a572idh/z67YRRkbMYludpns91j3oKyGBNIcjRtj4YZjGa30dlPbOzRb
oMwhRHe2i17DOU2I5jS1SdzIS7lqmJ0Ne7efprtfkLioBlqLSkML1aE2TXIlxvs9
yWMAo8086j3ZtL7I44twAUlyT3XdnIBkO8NF29efvlEl0VT5f+X8LIcU8avhAseB
BHAycqukff7HXbkvJMXD0/ViLaLwTOqwzxVp+TcuzM0x2rFzwj2WCoP8AHQIlROK
R+EmXaBxx37dIzJV3TwLoA/+xFJ6RIlhTseoNoXCUokeiSAZCtMdfJuYbBotGNmJ
d1VHDhGf27TcZeIa/ZgIbRN2q9s1xKGCoUY36jPnNoKgy0hxk6hSQClkLPDeamZS
PIXTpZG5eGcyUmPqe9r9H2CBxnPD13GZ5J3j7bdadSDuh9vI+lj5Ax9gF/vozIYC
DminW+NAXoQbsyUT8SfNLV1wCeNMUi/CvJ5gA9hiFP6wbSmd9164k6yZA5DZjxiB
xf9T0vy9w/AUJiLUA4ZsslpAMoGziZAkgoQ6y0GttoJE3j9zfdmuACWx9ObJSqEh
GIdcpkEjwO1iuwynMsyZwWX1cm3yDCtmcUT40VylfZRJGKAwzmof0yz3aFN0aOPe
vdfuVGZicxmIyYtEom3HhlN/tE4R1X/0qN0oJqHLhZVB7ptemnQ2PmkupjXH0/BC
WWeQK5JN1pwWVEIqHVXcD1GJpe+dKA/adJMLGJleGK5UKRcqNzsvzZlknhlD1+x4
oHTbkHBE85K3pl+3W/E2BVJumblkdVL01VnXbSFaxAoQH9gArjGWSypx0oHlW95O
Z+k8+2Ex09GVmjeTA2j1xbRr29YbCShHAKK95QC+kmfT21AU/lzFmtNcOcNZInL3
gK0VghVDw2HtKWCA/gFtcmrXCGq3vMqZd9rkAOiQoMXLBTdd50Fnd0/Wu8EvRVt6
En8EpZigWnNLsexkocQ7zrbTJ75hIicK0ZuiWQWXve+yPwEMAJPUuVmYFM7zdR/e
GxUQAjsLwFsAzH4cqz6pIqmk3a8DzWoB36OkSXGusZ4jis1PQU+IpJ5JOhGBy/af
gR9EQhEYH6dIjEg8P1H5FzD9uqiCQ+QABAHUYkvZlgTxDH8QT2V4pTLReVCXcE0J
3MAvTs8Vqr0/wCZHDQXTptt/DOtxo232/tn3sTwt5i2CMj/cuZwVdCtFkJl0F9wS
siYGthXQzDr3unCZwdxjaj9qCELb5Dc2diPnP9T/fX+OV3rTWs41xuFvm6U1hRDq
IfOBc+mkHRTwHN6GUbwGxPn/v/MqBj7ObAGp6t0ZFXXSBk1NQ/yptNCte2y5KW+M
TDv3OYdSikfB6aWScJcITAGABehrLWo+VylC+zJsyWUAfnWu9jcpX6ajseYfr2CX
l+vccoiamXcOeUJsov51SnRxkpgz4l0Mynvou8npHHgAWMGWAleU5KtcTyZSfWpD
yWWU/hyKIb+byCzh502hP2P+wSE3v5/zCKu20FS+prvlScZE48syGI/g+JinNsRf
XoSgha7ipqJTFs9GXkZO/B1k2dzcJ4HdPwmIflGOaTAlmoGrhXMYCSJFVnrqdF4+
Q95deNI0tmXcL/xeunEWn2Vzp+Xq4fgES1NFr0+xUz9GdDtOALsetK+4G8nJNYFo
bDw/UIDnhV6Ls3cBmpSFT2y7JwL3fb/2pXnUh493eRx4CE93oPAR+yJjuziB0tmC
8K+3xVO0Z9EmTOxlJJsb/6Cv6wOsGuVK2xfF0Qcn2sSje/pD5RBAzxm/bUS0xoeE
7EkI6DT8dToE+CNK5axmK3pUXk1hLV9XpBgHK8Zi71diLfAwDotKe38N33/xkjB+
JQGjW9woWhNbl84Polc8weUUYDhftgAiQ9eKF+99hkHRkbDWHUXl42cTDqI6aMU1
w0mHUOGVFDuRLBbomxLiKO+TlJEZA1scrgY/9nWH+/bW0iYyDUNLtGeui45o9qhi
xDPIrn3dbnV1t9wfGcwGJeg7sbMXyUCu4cM0+o5vawmF5MabV1WxGVjFBcOtp35J
q2zv+xtqUiG3xHUXrc0BAQNAQwclh77hz4YWRzO5y8GmPyWG4QyoWFmI6+eZ7yGP
/rBLyPOaiTGU/iouPWfultGk8zK0VuBWZwl4kyQJwzK3X7Drpd33HxnrYHJwKvIt
ASZFp8AESgH6vikgYNzASy3Odc0ZALI3DvhviqXGCnuX2tX5FKTv5N6WmUCqDUIG
pACR5gOiG6EWpfAeZZJgaOqv+VYgIaAqRwd1OQzU26V1ILLahyaS2P/bdycaJDyv
wA6gavxbrlhgSRHGZd/fIpYLqrSKFvoMn0Xz22eNWOUR0wXnrCaI+nnpOBJlDdUs
uvG6Fk3i2YVrZOLcUh0nZlNINidL0agLyGwRLteGucSa12zZwIOxbc+3cLHSM7m4
XZhsMXaaNwCy+KnPbMV8HoMzeozQHhVPb1nSh/tKXWemyePZIjn4Euk8u2Sk32bI
wgYuBGBXTqu4svfQZQa3eFjla9xvsz2bJRxLSKvAobg/wgIJAwFajFvEoLEtzVzP
a9HHhdbnMiRO5LNkja1PmDrN10vnC6hjB9scciELvCwQQQoWf5n2W1uxgltTtKn2
36qvmAcNATmuYVrwiFW2rauSZ1uC9VIS4y6gi2jldFbOL0wmr0dhaGJFP3Rxmrjk
SgWOseCXqGW+uVQzuYzhDYOoKt48dbrtWBpHAJIjMZd5IYrZwlcyjZ+4mQNB2h9I
TS+/AV4nm6pr4ZOGFyH1dcEwz5QPGUY+as39+f8/t+iLowUUWCVh8lP94MpOXICN
pzG01wDIXlqDLTtbPKbfhOv2Jry4WTLIj9b0XvoEC4O9//wyQJPPmju8e6Whx9pn
ahw9UtijrfmcnkxznvUj9VAGZ7fbdw4uYp50w1/bhuRSRJD3LHiU8GuU49BHuYdn
9y45V21ClP+wM2nShZv220/fHT4CQ6mH8SsqJrbX5W1NP+8Z9zMKOkQv3ZjCwMI+
tk+PM6YjtcpShPALQ3ShNrsh+f/Ag/NsmzaUCSahGyCSatAMclfnrhQX30xxQjCq
a9fYbJrOJmnuJFuoRVx8DkE1Az24NQ/CiaeJqLQG/1O+UAgpu7RJJ8XAj+51Fg4R
AOI7nkDsQt29L3RiQuoUhkPjqSqENllwO6BJDDSCC/xvY9/f8JtduIB57WQzPx/L
zGQAb1Xz0HQ3MJzuMRy3Z+ka16laCIXdzNZ5gtZ6K9bwK7SpZ22qCvxvThAtf4a6
mHAp5khStYQSQ7QxofnxxCS7iUAd5Qse2xdnd2kRD04/n1DR6K4BSaodmpAkBWt2
RwlaA4G4N1A2QXEL776DGSyIzHyqT1jmHyUy4hk040fZb50zYJVcL30M/O56rdZ1
6VUsY/YHl3YYSaBDBLkXQHHy50VabWK82Mrx3OSRqkCYrHvtJ24CDswd8sdAIVtq
NF3jK+6SCnwC3XXu99ii6lrHm5C0VTMckCoPIH0nOeuYadysP5cFzO+SYccOpUKr
W4VvP+wg9H4tCWm2K7puqhvWbi3T5P40Is0vfqRBuXBj1NY9ZSBlssaFd/jv/jc+
GTdiAP3wrH7BLVt42X+UqZSS4jxWeLIpuAeIJBTgm1Mmruf56BiTvb2XyWyR/Cx+
gUReIoBbMVUXhqMh1N3WPeVP2+bDfDiuoEKmLv+aMuqpz23tuGZM1BHRwIwSGTw9
0OI3VrLTyvqjwaFPc+15zjyg/h18w7PxFbtvh/jMuqSUdL7xIN2ZxxbzuZchZy7o
WOeaAKoUsd+mYx0jQ1yXqpZ5cuxFU5ww892WnlLPjJ8mictGMfBkkq1d+qZ/Bxsp
YIKHLsEFP3j2sRtyo7ENENkzdiMZtKMaz9sT9BCli6jyGFNarZU0v0SKKTad1Lwy
1tRZbaZ31QXtVA5xr1QYVueoUTyXJ5QcI7vn3tBAnjU4hfUX2uk5jwNGfuaFzD4J
++DJ8eTeq8raB0Xv7nSxSULDiVdoLTSYwYtDbr2TbcfgTKrgNHijkZnuRdzZEMcn
NUo3fHY1VuIHRqAvFu+zfTftkCLD5PcZceP2Tpie1D5ko6vjevEdxduthYLrPLiZ
8mWiB45AT1wBZgERy7nrOQWabA/3+MqbI7Yda1jgxq0rih9PK3gPh3WKXUO6lBJ9
fF984a5hkV3G4IQV3XQS8WOrWIctPMd3HcIN496us76wtlCPosY6ghWiOnvITm9s
gnwb1NYJmgMZHfRQBB1KG90SIUggcS25CyohUaHuo+x882CNJdfzERSE8Kg8HrBN
MG78F2OeM1JT6sHzpwglIqW7gd+Gbo3tk35RR6SlRx7Vh0q/t2DCTFcU5Ft393Al
PGj/W2lOzhogW8/l9b75A0xTv2TzAOj6U85s1UKLaKkipgkcCdGC9+uOhmZ1BGbk
290rGUFCplHMGNI33l6WJx64Klb5F1t6XAfO1eSm5eM7nlvnpQowzjIUJE3vMlWf
llXW2TX8WZwklwVHk+XN2cKnhfqNxC2fHfE5hYQ1lr8n9mc7VGqxvPFU3Yu0/7rw
F/eGyy/w/VkB/r9q20jbKkDw2ZF5+kNbtohF/yoNhvmfh38sh5jot4G3PlR2Gj0/
sGgF0d6wvpM999UxW4Qtsyt+5A8kYDNFUf08iIiPgifjkS3ddeYYINDBv9/8BATj
tiQFSBIu4tLsDdhXxrL0OZMQNTBL6DYKsYXizLZkkabh5CoNhh0/TUqZ5t0dF6L4
H+UfqeVRSsNnyIvkbvJ5dKF3MpIPlvvoqnq0g0c6aXit0B4OjGmvcExsJovVaVYP
VDv4J4FhyyiiIpuCQpBZSIkHJ7wo9pjp0J/FOElu3kgaDfaFHG1Nnhg5mREYPElg
EVRHlmXmubQe3jJYrRlXoHxpzMvUIdwkR54tlfpOvX0hbqgtAa5iolmyTa++4gAu
2VLMLBtGZYoE6DYEhk9atGjVwvHIWHDZ2gU13zKQpFVzY4jzqWJCzbiAW4HNQCyi
0AK5Xro+z/YVbyVjQaO0a4gExnal2C3fDctcH0gTjUiT4uXgl13kf6I5aYB+sLpS
shO6F36V8cNZvfotQJjkqtZb5cRMDY5oxbhiepDyP9aczBxNtGGcfjECsa1W5CJV
4Df99fpa26XBFChzw11vXTYVuJM4GGa1m8080+VJD/GxBUOmNKVMSi8isZbtU+Yx
yOjlFRSsaIzHuSHiUdGT+0tfKP5Jfcr30AoP3XgTnc8AiH6S/ZYkYiWGup0SFQK5
bz1aZjCAcAMmY8XC4yhxh3cxPbP3PX6wlnMOhOq/3s3xOEpv+NBYJt7BbGTVVOOC
x9C7DgmD/vpzq8WqmmstSfUWGYvtxQrOoOs9g/oM+AI0BmDB6h7G7CvF5o38+Dgf
mSive8ZEhJAhCmf/eYOEmgRkSWYAZYesdPRJFhKdRxpN1U3ZXnkDtfhZMPLIMpaJ
YPdqHo2EtySXzQZqCBWvKanqzS83TqBnlwrjXw0N2IEVYNDEN8HTqQIb8O4rkmVN
t17mu9cXvG6oLV3a/z9trSLEkEUqChz++HbEjGHSb828xnegh7lMhccPa318McTw
5yc6CoG0GVgx6btJS8nZIH7+89H3YPvceE1MG3K913UOZ08HKKOslODqQ/Yly97f
vCIfV/0Omo+faqnkZx0pnDE24PEU+bqbvcq28iSyMxm0a1fiQzt3lflV6qHHO7Nr
Y+xOpWClnoyONSLHG5phgYODaXHjHmWgAyeSl+yvh2jD6aQ9XG5kmFPnjH6SVPKl
oXZRIoVWV1vGbqQvK3tSgV50RA+ruAlRrhBIuyNhRBkTvIxCA42Gz8DMbHxU/4aC
uJwDkB+SLGV3TnOInvuLXe76Y0dN4YrK8lGkmb7W61hdj6yXXHfTG3M4TV0vCMdy
90LQCGERID90c02mywEcgVWOfkwPjba0670tUmIPE487pQ+MWVxG8fGZBEQfvOyJ
cKH1smsZwy1/PfSEBY1ruzhvO5P7Abj/vQxdvON271tXTl9kHz2/E37FX6xlHav3
g+GWjoFA/1pTFBdlQAdqGwJ2X7XpRND2aRBBf4aS3vRe+KDZdR8yO+amBO2morI7
eQakwNpQC97HiUsYyaFLTdajceBo3NWTe/C9zcSvTTd5pGiDOpKiaNmirzCtTGKO
hVU4aAhV5z9cQvA89dxMqAcntbYCqeE0NwEGwQ6BhQEg9aprXWV4VrTKZ8mqa8mc
lgV+bNNbbYpRqG7vZmdzy6/QOxZu5sR566XCynkJglwHvYgwd5s7iiS5ee5U9gt+
gY5yTiUJoZNl9kqpcLHvhPBflC8r6YirFrOY42qlUFq90H6+mMEdnzP13hs2CPkS
1coK6tggrwsbyQZ3MA6IpwcL54a6HgNxhmACkQOyHO+MdT5ZRts00/zB6w0Xttob
Y3rbgp+GAtIxlZNKNrqHjymJkn2q372G/rx4JtK0E5A2KpxEZeTFo9ynA0VfhLC3
qYpq/Jy5TodjWnvXsO/FqF4uw3aKIoZQ24DsB2WJKIcDkNrxgpY3Uf1koCl9vwGS
9HNf1qZrDGTcge1xo+vYsPkXmFVoPLg2i/qRzRvkOU1b9ZyaQsS88ca3jejTrVn0
Sh66fMH3+0BSsY5NjM9Bw/UFD6GPqlIwR7JEAkLaM7cFzirfKnCkPJtCX51yJzlO
90WFS2Vbb130wBJ0ILXTtp0E+YJe52eNROssnd7/7T3sEw1/YMmWR9Vrt0wLBK06
IUr0QrdqYkmdFX3vfQ9k7GgglZsb4Q4ZMpJLMG6lcl7jwOmDA9VNDouJBUiPXwit
U+bomLOABvpdYho4RicKg8GVSCgicjoDAqtbhKHGYxntOyY5eanJaUNtRv6HfHzo
KOs4zpC5fP/I/02xzpa3TuZQs24zASO4iwHnXqtHmfKvAFDga74ktxbMxV1KaImi
kAXs9yb94fBx6FnBWZ4XKxcFm/uJMn2F52FBQxB+QahkOFehMAQQUarbkANqzykp
IsSdbsj8SHCn0wWB9VqNJ7y9wYw5kpm46AJfQAmP+frwtJTl5O3hDj9S5fuYjm3F
gzEBhnOY7wIebaGkq8Y48d5wP2NGej31PnaZOtC7NvzKdDOXwIRg4ThFJvvFimqZ
aaXaBenYNsK+Y1OPDnR3pYHt5PMHZOUeIcnaE0xGr7JTYFQYwvPYdOcArhe41R4M
H3c7q9Oe39V3PzSFQEdcJN1ulwFN5B1sT5Sewc33ImZ8FJpOw8SeSITWjnwKsapq
GMvqYUkxJp+azgAsWrJlYZfFdQBuDYZgtko+cgzOzcJ7HImhpVPUyKhXUiCotMiJ
MyVACQ7pKaqKk2Hw5udVCDF1ZPxnUnpXyRwFR8VRoum52r505JXIBDPzwwUOFXLc
J7Zli6v8rAJkHG1rbvLSuljxcyg+z+2cDrhNGfbpIYZ7POdG5HUYc5qj6NiaXO2m
AXt2+jDDV2AjcMIWqSEdQ1QAXbua/AibIovenTwWM1RbB6JJ2kJVX/VqLeCmLYZ3
pGeSLGOAqRK4CPervcSHNtjqwb3fmz2Mtt5FBh0TYF1dUvil7XLBBL0tNx6riqpV
ffdTnjpPE1s6DdYqHi+v097NL/vWGDAB55xl48RPpruzYwv/kQ0RO4n5BPaVvlOd
8OpEJJMlUh0pRvYp9W74xkcPZWEyYNQkpUXei147YDZU0No0qxQ+JruCecOgBFES
3uiwdgSTRK+jUtOXFGGqWjU0mJed1RPO6MkdaJlNvHkx95FbkEvwEEAvQpZTzGnz
3yWv8iab+poyEMFr1Q21Ltr+IuRSeWrl30cFi72c2oTJlKch3RcLT0uB37y6NBCr
raCLo/jcVeAaVUik5vcr7wIf9VBc/T6ltkB5e2SHOBhC6PVu+7vOlw9tBSmfi49q
7+zyB2mj3wffIfrxmACmchxQvIr0ElaSQPADhDiFQE83yqPi9jN8JWo+lbhSLX1T
HGFa+20slAEpzKnnYjdZMpaMxE2RUCcjzsuX9dzTcE4K4onlIk4jqwukPXRf/dTK
C/xlguKOzdknX++oia05ru2aWcvJXf7NKG9s76r4ERDzjzdUpLo4zk52Boh7r2E6
XQs1w2WbX2cHQyc8cQ6PkBJ36lFBq8B1+79Zq4oiOMWWqfSNq/IcO5o8nBaLusRL
+uWiZD18rOd2fIKu/qeUHGy9hPgZyLgGx9qG3Vui7LzgWh67MzvkRGRJJVgY/ewF
oXQvz8WOQyWZ8n2IS6oYy4GlLV0Q/t8v2SnhQhLWn1QXnrFr+if6tEI9+ZY/nDGB
jCH81FWoSqXm2keJA4Kfnd75SIMu/OvzJKmjMy504g8Q+ztTruC/r1Bcgjow/iGC
s9niCPQuFgJ8YWIuV2guWY4D4qZ2cnn8XA3CBBLhIVm5Zx8l40HGD5rO+cFnti+k
R6fy7hLtZPI4PNs2jTf+ahOb0pULIlQcPN/kScF5VWjSUOFlgBG48PtzohWIqi/X
SPhDSHCLc8YlU3NCQljslSvwFtTQkqBKjYFzKVS84S1JhpCMM1QKwLqbYgJdiJ3D
mAGOsAgIE/hBXLR2ggNKvXXeiuQU6wRCVFMkE/gItLnpBjGOuUWSo8VN4d0nMhwD
gl3uzkYd2pZwEMQ5vRoTF6hzkbDQ8J8GxVDVnwoWGQKF24HdEK0heXQa5qsMdk2D
UUIiE3eOhFy/9Mz7sv+CCmclKGyq/LQjO5DtOq1kiDJSKLQg7OigWkK5WPMPkC8i
ycoJdNt1WXmOsZJuDmh/moUmaTXjy+/rpI1lZEb1Y1209OzBUf1iMaOMI6RNluNf
eMxTPKlybzf2PavgThfrqYaazyRqsPkiOUqYCSL6ZZoCZZheJcyQskR3kQHbOP4s
2ANHHul5te0Vsjo9j9inR/p5ODhSuu6NKRbwT618EVuq/q4tjqaB8dgeef5Rk8qK
Jy0ox7X5vECRNmVHJBe+cnYQEOmlAvHxxzULLg/rdoY7RU9jLGuVs/BWiAMv/V/Y
1SZA0iKHqaswnDuTxwpRL4oRwP7rZBtKwE0Zwxey0eZR0RMmJfb7CWOUumPWf/HK
MD2w1R/C7rnGsIZNeZc9u456M2mB6Q21sSIt3YcRDFTDTsb/gsOMQW9dWp42y/ep
ieBOxx0j60pHSQ/fa7/l1S1WfgP0fhdlQ7fWqDpGQ92MbHZTI0VvHqSJu6cLOc2J
FBXGQsJAyL1KiEtRvUybzwyUxTX/KC5xlXk8dRpiCAuR5a/ZMx8ulrW2fl8MOFn8
IgObZDRQuJlC8oOnTodNKaVwPLS7krtd22jnNES6HZ8BiOYBqSEnKvyQahH0pLrm
w+QAgNI2EXULBLdLqvuGvPJjkU2XS/wc06WPlUkojRAppRiSDqzJtqABvM6n0Fk8
z0mgizqxJkMN80EgUGbKQXuDkzZhVdN0k5wUwwReqe9qPKZaPbChjvPTA1Gyub9N
/5I9T3pcpB2QiT+FmDF2emZVsmMzBjIfCXuPM9/lxqkErZbkiePtcDDmBRir2d8S
Ql9hToLCRS/FiJYSTR6EnzG6u+PkTmhmUx0ubSFmF7DagNQjwYj647/wCl5gbOqv
BWEPgCcpLVldk4AJ0zr86WBnjm2nhikjaQHCdONx1HpYgC6hmBqE9TG7HxRoTvb8
i5yDNxom4qArsLk7S0VFbBQ2FJ53qM+QJqvZDFrQONknVlv0TWy/xUPN3RRELqpO
y+OXxYb8dUtjvI7s3HOaLEa0yCS7Q435lnm4t1Hxi0L4xT0gvAdVVvNmT/08+86E
3JK3PA1ra+89Yh+L6X47SRJPud1ZY6XQwmm90X9wpgkh/d8kBN9Y+KIAIWcOjSF+
6hcSBe63fCc4JTFhNLMwgj37oAacq8NctMm0tx46lsCbmDWmgjDR3Pxpf+rbPd+C
v6+ZF28oxlly7SDRjiBUC2FNxQ1bNj/5OH/CmE9vGSExOMARQTmjn5afApPpcbrb
Tgwv10e4MTouU5siHHRIOEAkzCRCc4ffhv+aR26hmjhmYzbP1svxDtLHwF1+32JN
jFaMdkf81/GdjctdrEGbHV/uUMaoiEM+dP1TE6+sGuIZGzZr6q99iJurGEu4mxm4
BV1JaYErqykTOqAyZrn8Ow+hdUEcO3AzT4G/vmiNtMnbfn9w5a1COU34c0zU4f6u
CfAf3E/buo4PBR2LDJhZM3KrR6tmb3H7RMEgfV42IRx/S5jwdKkNqfI3desqqpPU
ykAOF3MMBdbPccC88d5zdeV9SPaIPpYxkWHVLLxXUml5WPq1gie7VPEFq3zpW33M
Sb5L5V6z5IMiYqEg3GIAdmLRm8hbshw3j5bTUR7KV9rAOS5C4zARhgBteezlSpJx
/w2ICHCruvke7wWHDY6qccmsVVCC5++LYldK7XBHcMRdZECLY4ObV1EjgG09UTXO
ets0WqCAypFJBDMg4ij8g4hD7hTjoEFlcOPy66zFRCjPO7X5zWWiSesl5OZR6tHh
anIz/HpfB2Miq3o9oUIOjB5F57D2YKznQME2buRxFoFpbf2Oi7Hy8+/SH8izlWlb
Z9RwKcQm1tw0+H9E9B37a5C5NXVWXvgNjDCDxp12RY1FBGtNao4LelHbGATpyyAn
N1txJoLHFn5IIZBg1ED5SfkVu/NcYTsSYUdn1KAITrQEDEYAzw8HXY5nOht5V6Id
elSWgF7mUDbAGZv9pExsdT+YMqkM0QEcfXxi3HmGfYndN60WXHQbqLGvdvQ9Mr8R
mruNdEKRVTEZuRDRHANEV3N6Xbjq72FUdNQXMn+bJeQc8StYxJqkMzf01JranlRZ
yZP7TONHdyFoZ+W3P6YbyEohjFV/d6mOLHJFUgq2wdf+Y2z8GG6x5g85k91Z+GFJ
iDygGVWS7G3htuynD2PEMqfpXp7XrGmtOcDwcp1StQJkFO08QTl/zYYoYkYcW/VJ
4sOXjAgzqKxuOWY11eFLjhiVp7NUAI16vvsofBfEbURcra5yHfBc9YSyVKm2xPNk
nAAbFaGH9rQzZfyeU0CiVheOmYq6XKBnNCBfycmekVUU6RYwI9jjbK4vOJtz/fdm
5/JCJ+17N2jhij/gt0Afzh+bGJmtKBWz+cyhyjHift7fmFRdDJjeV7SKOIpSLAIG
8D9OzX3pw5AyXDbJiazckevlBP6XJVCpQdmd2vwSAqsuw+t6+kDv8FlF5ZHtgN4y
pGAMM6gD44juyrzCdZU6vAsV+cfXE1aOY65EglDhGsW0rpzrECg76Cieobnc1V5l
HRNOcwGM6xFT8wEDqfLpay79IoawDtx/Imu4n7AaN5n+kR0LMaSmf+DtJdEwz/2W
4SUdrHvylqEY04Y0rxFJNWf55LvrPwAaNnsKN8Kj8zV+tsxMHuIS+8i6WLJ4cgly
N+Ru3HIVarFp4ktD9ihWjh20owhHzCtoCM7Cy5CyOnY5UzVAMoChzD2//TxLDylU
g2zgJBxQVaZ/oDq/taR7uPMUD+u52TpNvHokH+eT1/uLXRVWNTE7QVg7SEg5PpGJ
Xh+VgW1b3UDPllxjhpX3c6x/n72KrjcAjOVYE/qV5A81y0zPe2qzWzV4RYWt5RmU
CW+XM3BxGz1i2I/REG7tputgEFVdk/+GeD29EToMUGM2Wuo3huivtXu6x1GnokHO
YA3QcOynv6+GMRNTWzkD+1lM9bJH/pXT2wMWYoDRlUwFlMn5hHjFda0qrmgjOgLY
65dzLUhflSfxCqhyvSOrJ7I6YwOH3ZstGLko6d6SNEIiEckiI2v6+5FvXTOzCuOQ
ztll4cCC7U6MPhcB8dwzevtP6YN/osdyV7FBcwKu4bltKaPNh43zYzIVn4dwMMVC
i9VHe7dMbHDCU5F7lE70J080JU/Efck0yfV0UE+0WESgEkv8A+fz7YAwbSEkRHKz
nN6YJsZ1XoJy/PcbHNO7vr/4LLjKrul5t65LvQXeji3jDe6ORK5xViuZjpeTDN52
txwYzBhpyeuR6krxAgc/vXvgepS01eo7iMM141hQw5DLnE4vXN6xhFQ0Xfr8P2d5
qNxfDVjMQdQ8SoQ8g0Fm66bvmy5/9p2d/SrxV/G00Sb+IZgjUJFynt3FvJ2Zq5VV
hiD8ooT6wJSs9bFBb6tORoFfQnxTCwJeGDN4vIVDK/Xz97TiPzkbrynPeTlS1R1J
ev0s3W/hzch1c5MgsPS7P4Jsq63Cjv0zA1URnFgS6NRit8RmebifNnLWg5CV4KzQ
ra+twYvmsh8zlCgtRwh7f3PmaRzMBZ07Iz5pPxy6qM+xA1w/+unM13+70Vt8nXhS
fh1ejat2fkT+oZ+HCtINfwjKXnXuX0liB92C0Owvzz3e/gpwsM6gmQ+p7powWtg3
MfRp02+ywx62YDNvue5x1oXwcCNQFF+g1LHkXa9iGq6jP/OqVj269dUdgOCD2ygO
nT4K0P1vD1hVhU7OVKB4khOj407lA8T+wFh7LfEaSZtctxlOhESWKl9km5rfVE97
NOdjlz5jCoUWwSJOyJDf3iiwGsaD5mm1kgPLL4FK+lmb1nZ70T0/nanya3owueZb
cx5B4TX+gHh2ltsj+rYzqtb7m27H603+ziIdJFGAoBKA7WAp3tG2hYPSHtB1VmL6
ZNW7qL+wure+9jVuoom/IVDX5F3ubaIKw8UvclwwEfISLx5FKW4Gy8v1V/rs3O6v
a67LQE2Q4Pb0dYRF95CB27qTD6ygYHgUFMC5Y0goTpIUtvVgohf4ta355c7EgDOt
1itSxZ9IIWUmq75V0IzfAil3Fv3vEjunNjBVMREpD3JWBcyNhwsaETy3ZAtxUKOe
9FMHh1iVtbexvZl3O9Unr2KktxpQEC7ils8KWxWOTOWP8x0SPlroRjBuzBf1u+ry
yY06jB3Odi2IZtAUwTE0ZTdBT0/OWPmTg2fTgmx7Btb/Fruv4tBTXceWqq4ekEKc
Qnu8hAd3gNWFf6F9U2FB6yf2uwLaJci4+6oc0cA3EsRkkYofNC61XlwY4pgg101W
YcZS/uCYcxKbogmf71i+130IXl6lWY88puWE9dtY0su1kHxInClJ8e5OeOEtjrlB
RfG4tIlve6yJ+G1nwQSMAcmkSgVByX0hlcdxmNssys0YHtacnKqIblxxyOgZQ1Lc
R9oFOW4qrNWz+o6L+3EHRRnm0Ui8W3L64tzD/xu1h1foN5x1q9Q8uXimxs8MjvEk
G6TeblMoaXJPQJ90MsO4/b55CmNWeA679jKHSjdlS8Ggt/SVDrQI99PAHnFWKTOG
FXeJKIb3PdNZ+CEVW38dBClxV5uxrK2rKzvLx4RvcvjRWxq93K3J0CbIGDZ0m3dR
a0veLk6aUcXN+0hJKDBfvzaoVzR6V8qPlT+w74ecE9XQHQgMSG5Tq2fki9ea6k41
PTwaQd+DiO+ki04GUSPUyOD4regGlhjBBdvhdpzIuXaCUyHO+P6HxVRD4XWpcekf
5/njet0a+f8d/bCFFo3+pZiRjRQpjUAggJ79sIra7iPW0tmg0kTmcqYSlcHZKgii
iG3gUr77Yozlxlv/q2RcndrGUsMgg0lJXt+mqYKz3MBCYAQf8Sj3TDNhOMhRD7+4
qUFIBoq1ySs6XqF/K3VAnoygsKa1HCM+bre5kGMX/AzO4Dq/fPby8WYqLOO+TpZm
aCvPnfnIP3OAnjQwaLgAuPTnDGxPdOYzpsuT7lLDSZgTGt6w3PUwGxuQfBa1yKew
Q1aHeS9ZdTm4dOOPF6viokHnF+nFLi1NkLCsPU/IUgj9hsZOnzUT5NJWChKfwWmu
yvKAmYA1pD/clRjxmrzVlz3pcXOxBK0U9d/Q7DZ4sbQxmaz9yr4zHvwENv+yx2Ja
Lt2AxLhA+s4VjuJKJHXSRCSisTwjGeDocsMybztZNoYAE1+ABTRhIeXfCEuUEyeQ
0jMQ5Ol7Wo9sCiAxCCEJyTf9IH4l6/QSOu4vyVjwOLmTB9RkPhYzk5V+veCjPQLA
F4j1+Qr0sHQNuU/G8bchoT25cTuHyBRQpxSEbrxYnIHoWT0FEUa0w8Z+qOtlqMNi
nqlXE/hPSNYtEF8cjOhwJVYvSkYAEkjk+aaymeecLCOMPXc7cedOXcrC45S9sjxz
lNF92NaoLPk0+YPbnPcNAGvoVc8nwGUQRXaqnFKml0Q2baA4yRIAAsohFbRCLB9X
fZoygI2cq4LoviKImnWefOHYBRZZDqYa5FL2K2m7didQE5o6dfOpj+FdlgxJatPE
yoJImv/kIQ/HBEQRxSVo+cc37jVfVYfOSziqY0k9wM7JimK+i6McSASri+3dgjEN
xu1JwzvF/i+myD7zA0fp/3WK1URQcyvTWmPvvnBlPv+45DLMHfBNnki5r4jenfqr
+hbsMD2qW8MpjtDbgu5dqDnzcZA7QmjieqdkOVbp2PTWY/1lSEMCig1XAWuZpt4B
UN9glTCz7VtkrmX0P9q6StaEbhzQGk5Fl4hgIR2k0xzDUqWTYENL73ZDSkdc3Uiu
9GzRP633PxU0uGmO2Cy8KgV3y59MbqJsbY4/djNZztOl5lEkmfoZYcWYKawUiH11
OP2j4VLP7ghK8MYy+HfISYumtuhwofcOn5PFn+5BESujJJkze54KY3gaU+IDCMx/
kRvM8cpT+XoCo0Q4Y2RZLY8qSPB/w1gTUeRLVUPEPD3Bs3zEXHvCPLoTUbH7nQLU
NJmJbJjg45965PyZ6fP9sh0HY9dPJfIV7YYGax76/BqpcvogjeTY1976Fb5VTl+B
81r6VNDASs81Uea5iCq+2+A5JTqosxeg05VhfZ4F2Eld2gc6efL5UybyKaLAAFSN
8q9PRvli1qnku0Qh/1dVb5V33C2QvpOGS9nNeYgS2BO5//OG3tX1BrzTUnx6x/+N
lGLz74AYH0lDuaCPG3B4N7d9vexE5u9/ht50sBCvK9Q4fxgd6ztbv0uqLVEbDTEh
VZUHDx9cuhxLsF0G3sqGHup6WEKfm8bCZ9YI5X51RDXOI7pa/KfcMGHhJIJkmIBb
kiHNK/T8LAroMueoHknvHhal1DpX548Q2JC53o64D9xtsjYh6x/25Ut/F7CxcPxq
cIca77i0RNymElEWbSAD3Q41xkQ7RYCEucrkup5A0UyH0PYrOaB+/ybWQkmLW667
V4XKDtkJsSM+Lqvz0reZnxLTrRefaPTl2rwN79P/qV1sNo0smM9XXcPEYdpdJMA3
+Z4TqlG5gpM8e1urBqaPK5XNiTJFdzKqkrObVYEXm7VwM3x5q4sW46t2RLDGvRNb
6yIu3wgU4XHIDtUIhBcCiYTn56WgH9FW4ugfY29Zkfw5Y3z5rWuDUeXWGqIL6O7p
iaf34yxftVvDT440S5OrZheIp7zjakmNef58wBhv2m+M7dmYddkCX+rRpWsd/p29
PEQ/fV9DGmYChMP9YQRNX/KeFh90vsPlFHmKE0KNC9PIhr0bSeHk5NboClkIAj1m
irzmibxueJO7Ruys8vkjwIwE298tcIZs5clW/OM+bp7PMGnxAaBCWJ+6ISS9lRkM
BsaPqNfHY7cDd+ALAwc3/1U6eJv0B2Sq2LW2GxG8prEQinP05wNbyutSlNg+6/Z+
HHM6MEwYZ3z5ZFtsA3sfQQq+JMV6jHIS1lRRFAO/wYwc/6AOQ1opTwDa4dbFowN8
EgHToOHj8pu+EeQXK6NE3oagenmtIPqGidXRmxJPMdhdtm9k+xLSJ4gnZ5xdLvng
8xBq+BUqgazYk4j4ghMHuCnPzOHqcw2SDObUH6RPfd1P6WU5DfjMAdufmh8M5tkU
+2gqLlYlOPE6okySfOb3u1+scz9qd3SSwiArL2zTlTnIoQ2eVbHeI0CgNKG1eo+J
V00eDOM/1tQj0mGMutW8FScThzzNkNgO7z8fE02O925TpOWFtujMOeOeJZ9xnkKZ
IymxaVpicfZ4SInynUhhHeJq+x5sf5M/nITMRRpIV7VfDO6uH6O/Zj5HGLNuYxIB
1rLuT7hA4jPk5ByUZG7aPlqMJjxSzlipSvGSBAMqmavfQ8bvkXfYpXfehLftinbt
vlDru0spFkc3UHTI9DuTGUmexaxBl1MkVd0eWmZOzjMQ5qVYG37cufROL2XLmoiw
vHcKK6dz1kunoM0L68RrDfW6yv+Ukj0gdYTpDSL8PpW2YtKhOYn6ywHcmPhqtBCt
TRdI735ifXa4e9AvnslIVDrJMqnbWAMOIxBfBwSJ5JIyhn2ojCq+mx60eK6y3eLp
1z5YiPj7vViYOgNEfWEIWLJNexveqcOou4oWH2Ei9nqfeZxRBA1YguGwks+nOgiR
aGjof+1PFt/SosCprT4Xg+Rrcw3T0phKGB/HoSKIIHAhaes4/tS/kvhoT46LCsKk
RswiAPuXUzDG8L2dqwG3z1qzlyWMQvqryE8VaIOeqYAG6eHW7uWRGozM+7oUR8ID
Png/KD0pNz5KDjGjIousTUnQIAlfpRidO1mJXdqJWMoXHkWYZCNHPdxl5EbfxXtY
5hcy68HTiJm04JMy9r9LkCAlu96DU9dQ6m3pivijniCDAhHL35IMzD+3iz8VOTJ6
ec2eVudGDQZsDTKhTMyKTltjIMWbbIssLbHJZkuHSfNYCESCOMqVSYKQ2qMNCf4Q
u6iuhfCiXyYh1tj2TF8WH/yYtR1lprEICedL8XvuL+LGWvFSfq4oGlA0b6V5I08I
wZhSa8uaEetOwNYlwSxm8OC1qFYlchP350HKIJ341GncLLTdvvCWyF1bUjbHq9rR
yfmX8gye1cKTXOkLdtxuvp/omNITnW65PZUd/b3twGZtHkE4U+l800G8BTswrIjN
k660JKkY5dOqCvO4IOQT9TmpRioZVSw3QC4L3qwUuetO0ojNRjVx14KEwtxEB45M
33Bg4+tXvdXLtC78lo2uN4EPc8AMmMaoLDVRC1VFY19c8bzeJcaNiCP8cpzuzgFK
vXLQfSlcfewEG0nGXrZyyStFQPtVMuch//HlHQdioGUnGfEbBbrxoA1BmvPwajuB
oOhzpBwD69JmfIpHs0stRPaWXNIP+5jyPEuYSYc74oR6B3n63mh6wQHI/XOlwN9R
caLdMnen3BZIc86dffwAAbJy9v80q3QwGcSiPOKGcEAEnklQyIZLw38vzJCGzUhW
p8xX2ccQ38kGfueInEMSvd2P6KcZNuXzRGFLiznMpwepiIsszCmrCvxjk9CStUjX
5Boo3nwuFOtv2iHVk3yJmW9mRrTdk3Mvlrtv/XXQcVisab6z7j76pjKkLGukA5oA
fq371WR1Nb1tJxP+dQ1N6nqXwl3KAWrK34+dXMggXET4IVJw9lx7ndnb0yB7YXgr
UzM8PAR+2LoRIasFT28aAMArEM42OJcyiEnDJWAZEr3q9NuM6k+lpKeXFr896jwQ
slUITcNOIBV+7LTtokzCMJzc60JljS4duOziE79q4FHNvt25Mc9iE+s6Ft0fe5UI
e7UEdeSsqgHsWSauXqmbI3WOqFHWKVyoEe1aHfukIgqqco0bJlj4oKk2M5wxtytL
rS6hs9I3ShspkaxzmkyycPQMx3B4WN/rYN4AhyM6Wfnr4zETJBS2ZiCjRjhW9ILE
2DVl2B7sEkwogbGfIwKR5UNf7ASRVbkE9uo1CnoRaK4UP9SL7G/5EYV38YwTuw1J
9NNPmtc0pvNNZ/Kn5MIc9SO9YuNDRTwr9nEFbzO3iHbh0ZFvdN6o28uMyPPy6qMc
NFQwqVTW1cjhx6StN3J4a4xtMYqGEsYGnxCuTutQ/SaoWdAgyHOGlnA43LPql2RJ
cGC9UWUxpxNV2FdcfoNe/0+iXgEy621+szQOim6n0iKIeD4kQ2c/RtpggOjTog9g
7aM+u2Kn9Csor+nGF+BCOcc80EJewX9L5E8R07/2V7TLJRkU4P1HaxdOOr5tntCw
cccJ9iVrLv7SGHOOqpkBgC2zgFXASVhlqLtlO2Fasq83NZZbUX/U3Yt2L0ksPY18
3zAoVYOfgbYYcMPouf5Cromv5S8frS6ekub/MSm4grhyHeOj+iYvYxkOb8oxoCC+
SxLGpsttiDVS1RJS3ow54G5d+tst5/ZY1sDzWNURwX3KMOtVGmBtN3b885vaDxRI
KZNKXKJRUMn7SHFgOKnNi4ETijslxGo5s1SkeohiwxZmdu6lW7wjZuSDsDWEZ5gz
rpTA43QIdpn/o6WaKI25ZyRkrOZydFQLF9VNIPHoUSik6owzz05U3hGDr16TLYcT
kBS9Z3WGekyYZFDyn2DVS4VTuzE23Ej/iAOJb+CLhrS+bmASfRUHR/AQzsD/JDBO
pNCRFbal2f7eYHVjzVXPZUt+jrREpPOK1vMlk63VSnn4WbK0mwuTuqiq2rRQKDmZ
94Ud+nGzhHqBKU2hzzMajRCWN/0yb+EBxFCX/TLsHjfZK98XsMn6lKXGFAc8pa3Y
McWlI308BZ+YpLwVBqAIk7yIJ0p+4pQAJ4PbMssowRhK3c9q9+4Zbw5bSg7K4+LL
GVl7pPxh4SZ8yFhikWY66/aIgOEjVn8WdZ1nEaSQUTrzhOITEIfmldziHl+ALC8i
oOYUKeT+2eJgzClyUj0Io6qzDWCGpySYQlomMu6mjp3CHlsbAKKZmNozhb1PDdbl
qn5iUEEK99BkVgBi0GZzX7agkei/6LiK3dDAseb+WoOF8zNUXMjTXq7iagDMWDAx
4U3p/S8Jh1fe62jt7RRpx+pYSNBdNsxPuTypRWAgZv4//buycXM5ZT1cQgk+Rkxq
WcNKljXmEt4Ad1SbNEhmTxUcTKpKlNm8pS3uufyDLguDWLdEe0zmJMthJf2RiyAd
pnb3v3yzaLn/s4A5KjdgPy+qrhSlUSnh/eo+g9XQW1eg4CHuzJLwTEAdHjQgkzzl
mD6yC6CRAScbo7g3D1pPT/gNDUWGnmmwD1hJ56ZpTS0JLdrxs8nVk7DyeXxqTIZd
NbP9FDN9eo+Hqo5PPfJJKyRG83SF/Pm0ik/rEUjjgqENHGSKoif1cfv49RS3I2wA
KSGn3OFo6sWagojbMRsSp8du0qHWoIikKvg5ndBDv6nBG32Ely2knLfyVzQU7nHt
LujX2SxxOSOJSN6n4ijzPPaTO1R0123VaHtE57A3/NUsdNiSsEQLzoIxV/JaK5OJ
tUFq/ONIsqun9ad2iaISwpCVzvNwDqM5ZchMQS9nzI0db1h3nyoeat7aJiBikCbd
hY3Mr5AR0xERw5yR+o5g9NYJxZrOedm2D3QKAg5rmqj17waUCZeGBC6W7TUu+k/a
xpt1qmRg7BCNBTacXqxHtGpP4gOH5z/U7IC1It4Hog0nTGtw0q04lkYPjWaYK6J9
PZvXFybksf0gIc2yoVCiSOHndBN7afHanHV8igQA78BoOqUGxLmmL8bcx/FqtuUj
V/YD5rnPM+605S65wBsNOTUL945HcOGJay+XB9LJYjR1ouoCVkV0A3RuJnk+e+KC
B99tizFMvHBw0jEaH0MFffaPy4XrQEYiweQ4b4LObeBGW1lhZRgPqJaB9BDLPouY
nFNLCIWSZqE+K9g+70Pv7+Gyj+PoDDlwOpmfxyuJ9jStmk2KtTI8qyIggL/Oqxnt
dbeprzcuDUY8PNEZ4Dd09IbrdP23lf62CaBtcRnQlJGX+A0Mpya4GV2gO6TIGKmq
g/5rR6gqG1vIEGx6Q0w3SoU+xNiV/CF05q1OXcMQywuB/n8tpJ861Xj0bXGacaTq
W0myAGBdUaJHYpekUiHZH9GXR8l/SGLpzRnDHnNCc3TcEpYQ+IjbaEU8ROsfF/3Y
DbfEVHH7/qeaZOOBJt4BCCLdLholJxWzaQfUg5lCylnEvbig2Haf48z2Dkqh0bEv
S51lRAmRmYzrqfTGonMTmEXKGwO7Gx150yIPF9AUHxdPF1E7FtXd2z4/hZRTQ8t1
BcH/80WGL5V1z5sWYwBgLdWy9eZaWFTm6mkebcB7fc263A2iMCHHfViI79OgzT4F
zMw3NaHUivFIWEpG9P8be42OXvKT7WMnNbc4yY7NHNqfCVqFRu0vlQIba9aXmsGO
gVMbDLfLbr0e7r6yx2VPgkag/dcNKe/FJnziuim6R8NI3orMQhGc1vBpzPUYJyxH
GYJvEmNqFnFFr26asTAmhhZt6IitGSG0wJGR8USjM6gFrwKLKNL8UpugJz3urNBs
dZdzTlFckNSn9GbIR2djl5mE6lb17GLdGkjtvKaHLNw=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HXYoKDvyBZFMiBZfgav0KJ73qYEDWxcTjvJN9voFEdFT1Px1iNER1SN0XE2lrjN2
ClU+Q3BtEemRriz7A28BKQTfBYDw1D/Aopy2LLlD2h4f/AHh7ppWCHzoCNSzsvk3
W/xkFve9r5t7f5IvUFtJ2VexC5DVdGX49l3JRARKueYQq61SX7EIoEfC94z3CTgo
CjxU9i7pnv/vZ0Pwry8GQ13H1GvY7CGm3/es/OEsM90d9hUmoRr9UVUyYEOUR8Cb
jMR74cv0vq90j9ck0ZSROau11uU03qDNt8q2UCIO2tdZxyfspuY2IRF7+46ciIad
6T+PjPC8g6ERT3eaDoEAlQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22512 )
`pragma protect data_block
Z5y0vpo0gFen+rTDULhm0XJ/jIbC591jvMAhFR9k9RKi0TyvMlNwpfh3ZqPFDKEh
XvVbX7c1FFVfQnHaLJW4OO7ci6k8SXUfW0FQ67D0l1RUl8ow7SexXFPrGdkTimfB
oezxrMXix9vv6WUMSwpPYSNoOqXjfkHxORDjhpaPAaTpttgImK51eavY19X59MGn
kLcmyx3j8qYte86VIsW/3lc7d+haD8eST/ABb4u9RCUDF+M9VHrNeISuSgESthz/
at8zOxHc998YSzYlAnKQHigpe9TLXwG7C412I1ZlhopyXlJgC89rF9xUR5WJzKo8
1v5EagDoXpkxyEGzX8ddtTzQez3N3Gore0HwDW8lP0njQovs/PvUdInW8BM/8uH0
18EBaWIq7rvtQaEDs6BCSQ5dKbF5nALByUXHmESj2seOlbuLsCwKykVPffpPlv8S
C62pX7+roRRnK63JXjPSJ+Asi4HotyWoRWuHt8LLgsQ+H3KLjD1yi8Sh1SMOJDGA
19wh3a0pFJlWeBXS5Co/L84+psaAhGOt2xllvxvvzVYJS8lNVXAMwCxU+o/xpdQd
c487iSiHq4WDwuznb87GMOuuNVfTWWH+fYPHItsFZh0R1/YZvgXBoYBocLvJCrQF
MhfyJ2slM9qR5rot4jsf+pCvHupIoEazTfpjm66gK0Tw5NzDIxYMIQ7XALpqpDVT
0lQvYl4PLFJJCjK7+c11KNhucfW/Fgkl2LGd6icxFnjddIGjPpzvx0oKogEash6c
Lf7GCJX+Zl9qqGkB0Qjv1kEeSBHP8zred1vxY6V+zGMvlehCrc6AgYrU77MvswnB
AQ7lk1BH5eKZpx86Yg1cIbCULeo6vU1OHJN6PBcE/40i3qgp376i5yl58BSRNBn2
tvSabKq+QxzQTGpUvmaVPkKb9hEonMf2pgDhKR57WaiyC1ELvTI94RjJhkVSiTSv
onAiHs/w77GA+lUwBZAwMK3B1C5+z6ZYVCP+Y2BxhmRZtbjKeUmPfiPG9zNtAdG/
e9Ut5Kf8qUPLm1udqdM6G17VcvDmQWLhMNZ1gDY1J9offbg1/HGNA+bO8NNiab8k
i9LTXsnc7vr8aPq8pMsh8j2pReFAMBZaIwElLs/HXEFH30WC5HYhWDENJ9k1kqbu
vOEM9H4nI2amQ744UrxHbN37c7sFm5iXhAXQrSunzaSMsf4RWYpH3ajSSdm8iZfu
ESwxgXnFpNdx9jtfNluvrWR+/Hw6moOTzcjBD3WSOVsch8VEMppg5UBPXvarCG5r
aJXxL+DyQ9bvcl5+SsIoXM++WalrQhUGGgzhhh2faeobJRtHWI1/sExFb0hGWwnH
gToZJtz9zGfFO+udZfQYgE3hsQkwvrvjCkcvwBlPjPHClCpmLrHdMzeMJmL2gmiL
jXLKx1PO7m8BFBOH/x7DNTiyJMlNPW7WjpnN6dxX3Yd1z0M4lfxTQLJh7eZzGZrw
AWikA8FRfh6+nrMPvZQWQ1d0Y6nmw+1jqIBHta48p5nEN9K6KdtSDf9DI76FrCe6
tciu6BlYyW/T/bCPNfmYQw2q48BLIsbm51B/ZIsY1TVmJWzmmAMAUik8oq9x0yjj
7J6NzC3hYaKBZYlmya+0+6xcoGfJoawJlv3pexoipD9ln3ZMUWdjDRuGc8Q4vnIg
xbkX0X47t8vqKnH5CtWFoGoRrMAJYq0cBKGfMo3wDxzAZkZVhbU/8Tj/y+rCUqtT
B3pKhXBkgBTvPGurR1zGGId7lnQto5W9DZrqjpmw16IHB7Td07HDVrNvF7LVElYY
YMfF/M6raF2GrGkldqKvUe4JxnCtLcSspOTblehVZnYJQrjUDCHGiq6l6qIaqNpk
S5RUdA8poSUmvCqayb78EQtSAgfEodi2cRdXzNBSmaj5YAdVUjz+dFYDFAQr/uBI
syoec9IZbdHpNDm3rKVH0A1HmZQVdAr/ySCrEgvB8em8fzhqAZiPjv8fm3/jV1sW
xxUwINZeyROWIQAIGXYXPAEFDBSW/MXnuXYOm2XMEuThDef84eXqzag4yUKcZepH
AhFGz0rEg4lnWznZ3B1HZj6PL8suVNc07BOfMwJvJOpcRW4DF+8fAEsTMZcCk+3r
z/8Gnz2x2+XnalEkdJ7i5Zsx5EvFONPrqZBTh8Zju7y18YvGSSZxEQKGqeHZTsS7
0154OkxHz18CuilLE60ci3g0YXeJNXnKhN9KnJqZkksdC/jDn8L/3P+dUtHDyFT/
rQYNLFenP1iB2IgM2QOVQiAup87lsYFepOIY7qp36Pi7mFufq7q920d7NKYvHe6t
LDOE0zb+vJpZ0OE/QtbGk/NdsaPyEsp9LnDjIOVx/m3RegzvjqHbBDIDy7K608In
9/gcniFYf2/bZGMGSZbPkCEbjcAYb0jxsJKY0hl7CnT4EUzx/7UcN/DlnMgLIFzc
FrBId0ei3P0r8SzA6Cb1Qoe4Rak0DU7sNz8aM68GqFCXEy2Qhn0IJ32gs7xohtAP
gWaaIiApxN86xrofGHwBxqeBYc46F/ZhfCJrDzq7IUPv/qVgKS4AI4VnAlBqdK1N
lyEow7hThVQ9p6XA3BSODaIJzHU053EKav4C4CtnVL5Jzm9bTBa1Z0aLM/7NCuoO
RnGSe+WGth8OIKVtSCiXvNAhhwr7ChvyK4roMPkx/YeoD2YZwAgUXmMWMlRQ3S57
aEuwWVwdKi6xxfq9ES/xuj2RiUjYygFxt4/UP0w2HDH5sI4BeIc5FMNCUuaddrh+
9eEhQcpn4xFGmHdKXOZ2P0Y8LPIO8wgAddCSDuMWEx5HcmfiOdbS7Ld8mpZrIQZD
ppACrj61cY2UV7hOmVATpohR1uJ0q7klVDZoI+UdSwSbwPL2c76SbK3EnkI+p4CJ
iHKsiGg1uarqlvUGwS7n44E2Ile8dx9vuRPjN1El0LUnT2MdRd54VKMQ+If94yYp
l9h2GJoRK4ngGu/5FQKbjQr7qpcGlgFSWv7/ekJZUUuep/bb5TvFAUJPjSms9yKs
NTJpnS7t1VmlprXOrVfdMNDN+UPgf6JUc+pzjsUBdDL82raeMxlwmpX6fm86XOT4
eK9HKkUkZiCffGbmCm9Nd8MyuENR7jwnYfWUoe24tzyauNFux16Q9bbjSM4Oelmv
GJHXoq08t8VTe/YgRDGmA/GwvtXBRINt3SmV/96hOODZ3RMFFlFTnG6HK7ZyR/ml
Z/rBDLwjtLr/gj4E0ML1pRrt5znBgtD1lGB665GZ91Xjq5KDFvKsE+WyB6eeVVsb
VTLBgLeUKxS8CWBiU773yvKA/AxJc09NGcuP0XCKbNnEK4+NHZv+bFqQt5OQk+cS
KDCNhypK6XR3I9/tmpQesQcnqvZfW6lr0HVuY5dhsp26s158IoFgbBagZZa87Ha8
DS+PXZB5Ch+GyRm9X8pd7S8d1glSsAbruvp2B4xVlUxe3nZJ1BZ9lZ8qdng6GpK1
aO8LoUmHoh8htgRecf3IJE95rtrmbH62FpJdsnP/Czw4d7Hob887GBkAIZJZPhcj
9WBqpTUHZb8dbJJop1AtwycISEpr6iJSyCPmqSBwXDMR0wdqE6tRYIDDRmIqmoUX
h3zeZ3UwYuL/BgTHJwQ8mqxWtaWN8K3ultawUAZxkjEb8uQh98huu8DPM4ge8bqG
sVAIobXtqXT8yLKAjXPVmfNfciX7tPh9Vcv8Cqa0h07Ig7LyOIfyn7y+zZOnfI7j
QIYFBTowX+Gnre37/GoZAMacOqPyoBUvXl/kryLIQdzDuhEm9mAlTz5kcJYrqGX9
+gm3xGucf2Wy1ehZO0aUQpjIIm8GiWF5KfIn6ROyDVBA2SmkwECOFVcXLrPCan+2
sLfdEoamyj8UB2Kk60hftyx774ayGRVdelCIpXK2Up460FhfCaLRtIuj4vmx7L46
BSPJVgTFse5dLy80ABvJ/F0hCMRU/H31EcanUTLtfQxZF/GBw4GOvMZlDHH2lfgn
0gAvhkd2weJLlgBCVzX8YSHbvfuwWPoFH6UGVputOzBD13vDwLuVEUiXaBQ1Ly4h
kr5fKZ5+x7HlrZdsLd2E+ZaFhDwSwTa6p+KEoK0JUMefojMgx59gZEDkmiEgcrzV
61d6vQWndBfX3zE9r4ILc734TPAdkQ1Zv5PuoZia+mMY6OYhuoFRDlxWEsf0WHSH
IOjAA6JCpC9ZYkcFcwoRbp1vmTLkygg6A98mndFzCKTSsWiFxZI8/n3RAX9xrMN9
DOP14VgAdioD1tIQ8vC/iOx1xR8hiPMjlyj4Me5zpwHSBh6+c/4xc3OotKXt1+fI
htMPnF6ATUBkkLhaRONeggNLJT9NKAId5uS4QT1b76u7vtBtn3+vnrRQIoWpp0M4
Je/yW3x200Lh4LXiFBZbQXtZYpvyVKuiPopiBD+FQjrBJDuOpXY1mm95QVpuoBPV
TLgrsM/w+Gqlv62B2yKW6rcNpJyRF/jiUFvyKSDU4nOrUoY3RRT4NYoxWeOCmWks
PdlC2F8DTX2QYe92Gj8Xy4cyfbaSnVlJTVBBJv0rcFKTMXSEClIrvMJEYWsKV3Oq
WgqbzpKNg/ZVB2bGdLUIVmVabWTVmrf/n1xXGmzT0wpMVmdI15ZTiOzYb3krIuz1
HBfgZHI0DNX+hoU9wVrlRTGoKVsXdkJvLywltV/EtalHVorcpFk/q4eUtO4fx6Pq
oWs5Kk9wpDNp0uOhwR0a98avoSarc6fPzrEfAfF7kj1XL+KWiXqSerQuCI0czeC6
xAcAx9fy5JTuDbqSvnbnrR9Lj1k/fqZKRzQ8Mo5NtmBD+CObbCQt62YODWQhjuQf
AobjDZP0+1muj/Rki69ez3Trq57TTPpyOXLO1JWWj2UcNsUXdkN9mCDrqdtpsbSA
kYrpkzbDUt4AxmM+y1cU6DnSiH7w7GgTvAQm7+2nMRlekIsv7tN3bPdF27tKA/rr
T3hUL1wxiilgkEWnSwGBOYA+etvz9ya06a1UofbO0LsN/LeyOTkwjBOmv4zuwgiO
wZ2+/GQfabfWVvSEGABWqFrdm5kTnTRndAbkxg2FysI+MWn9POrt6l3MKHRbyoBR
YmKLSnQ6t0byEW0hq7gIQqIc9OBWGLB1vd09EPfLIecSvigZ9wGle1CT33XUKXsZ
5snWzbajFrVgsGibYTM4bxmdAdivrwReGncD9gxlmqMJwgDmD9xNXhsaGpXqhRg/
ivZfqxrGlrBKSQZDQx8yf/lQWdQ+cZA4mUV4pX7hM/5ZI7RZtUtAY2a+vjKDQjnD
gRXt5SjGq95IwJ8fy9ugaqD3nO/76O8qAJmWV1oJTpuiSXQOj+FTZMB3ao6Kn+uq
uEqSPAWIoBnRk4Ey3ONgYXb3fBA2yYhO4TjH1NTPAB4NatETTyr8VL7dIgiFrR/i
rTU9rfbLDUEG4OJHBiDRkkSE5+ZH5aivvsoe5VO26T8RxlK4VjRDxPNt9BnzxPtR
TrLg0BtDNkQc4UgammMPhY+/E+jGfmGRofPkKQcSIz869z2PIzkga8CzIsiED24G
/qw0Av8q04bcnwX8d8bq67ixUIO3p8iK2Mkb6Vo1T7ybqYIRUrnxz04bqQTqaTB7
xjBUUE2LW+YpsSDUtjIyfv0ZC3mGr9P3BI/5OxMJ+54MdYSddyQhCCVqw6wXfeBx
7DVk3ce4E+FKVOHy90TMe4dBaoF6MnfZvFf+BHYCDPWpgz9882roBiWbEK9hZlie
n7uVoJfRFPBlaHyglT6h1nWX9rJonbuveBosZjc06B5uZSkRGc3iIkYdCcQKCDiM
wFrXi5exhiJCa4o6jzZmGO1u40IQz4NGCJEoap6Q/aCRJeQwSJJUswfSoGgCK7h1
Yeimjjx6kO3oPkumk8JzIVdTNvoYiwcS2m3OL4Mav2Nn4XujPAbh8Htue8bqji4r
qYtwYeQdDUaEQARRdj2J4rR7LTtynyRgBmz9ONdptWIc3HSlMk2pmJLNvlsBcqAV
DIsgaQzXi1siNMR5OsnLAkYs119iatCpi8mEP44/r26mrss6IWvaHjzBO18eNKor
V4ThlMryecQUtaoaATvZZdo3SGfwD/2pNR2BIfc596qvBf0Q/r6QufE5v5DnMKSs
M2Py0/OEF4BvxKCbHkMc2yZoxPd8ZgyAQ6V8jVdU+kZ5IsHhyVmm5MrNKwAyI5CO
dW9Sy8YB7gPyNhGN/7/ftRIlNRp8Y7O/et9joRqhTYKR7ekJ+bkMJPRM84m/LcpL
xnIaSb4kfkWWbMvMmEGjCs6ZCHCjZR+jDa8W9YB2zfz5njUDQsQlVRK8F3gEve58
w9Swl0uc+EWxFv+JlrAIHwln1vDjdudCAiCwm6z73rAdR7X7L2WmWpSpNYp8RjPI
OUu32kMmuV7Dc2Pa4ZLkFbclDUpQuOtgX9HoApMf2jx7+ei6wNXjip43ACXtVtR2
Ng6AVdPVD6+cJDoSh5LoMcEMPcJ5L0czmFTHPortgz7uhcskoUVKW1w/ZGaRa59u
nFVZcMPWcKARLka9wBLdD2VoZVXVglsdycGhe3wVZKOVLwSpagVNa4kkNll0egbY
H+LhT8/tQ4V3mirtHL7YrfwXj5a0OST2k/9PMCVtAQGttoxAwxZf1Mr0FTl3Ab/p
rJ+zmPNXa3V763nztqAA1kctva/jNQ6D3BZ+7p+c28aNKSox8jAZ7zkY99Oed5yv
plnA3sxLUY4CVepHz6eA6UGxrBZjPgkKnoD85zs6jaa8bewUqnwh/UIL64r1mTzD
PR6gOJfCCcL/g4ZlJ8gzsrM9QmbEer3e9g8/8keA2JosoR9m1IF5hGL1PdKbxal3
QEFOPudg4wV7Imh5j0Bt3SXVAuz5HOkn36b9CAkm5ZsbCpEdC3sBQxDqY+dkj+Yo
6huNSTS/O8PhiVcf8cOvPwZsRBiAnd9SfYUpwSlENJOdZQ9QltsRheGxW2ZW9q4T
aaoo3elnmIotf5OvIMq4Ult6Y/xYcD+JdtIpJs7OrTt6iJ+6Y0FtlMdPYmYib8Hg
/kTYW+eUkHCM7igJOEZFqy9M3CtkNHIM+71P0Kvd8mBD8d1qwxo9xV/PTTxthIeq
hP0gp253mFs5w2OapTSLY7e5R2rVp6JtmiKaokrdthSP+b+0+zbjvvfg61evqUiJ
CwhwTnzY/Jr4nQyP5Qy6KslHZQUhLVivV++EZMWJwV7/2YOzIiq6n0ocRrHQqUAz
AQFCcmW/iP1S76kRoLB9ywtw3C1lLdOViccMZIVbKmF5GzwNikmDDCs/KgYxpO09
RsoZC0w170twWsGy4PPhpApI6PwO0bB2cBVij74i1Da2CVJfdBfQm78RiHusOQiw
uKwWSPnbazhwOaqxvFOeOccwvWmwMMNZHLLvRUp8TbNrZ4Jbvt2DEfmbAkUvJGG1
TaUTtiKZy2oqtNegYbaiQhpWpcnIEpK6V98oNtR5obX6lEeuArnoKWeMEoMSO0vZ
ZsS+ja9rCGCXNVgLitGF9MRzk2yhf6bKneCWuGj5XorWoINbX4k6YYOxa44zjwF4
gq3/1HMuRkfBZbbApaB2984ehT4E573kp+K36mHDVOcHMNBzQVbHXyAACu2o7gcI
6uWXJznJ7YZRfy4gJnkH7vaNKhw8eAFARBawCIsHBbPpkzkpOXdzYyjjtrcLJT5f
HqmqHVbVE7b0dO5S4DJ4XI1xX0J/VeMObqUkAjYR361A78pNE3fu08ZWazEhU8NZ
II8w2ahLUVJHnNSDJSILMdCBtofceeOGfOGYWu1X7tJwpbomxscmGg0LxxmzcT5V
FTuplZ9O98S0hck+1Dse5AxMhg03aVG8Z4r+VjiWhYI6cIkq43LpfypqMh12eQWH
SWdqKlqFsW5kaQxHFnVeAmQaRl+iABL+p3+CKkwuoVoPNdrxeCopH8DUTSGlQZkY
ew89EZPa+l1KS1NDo0duouLuycdK3Irsh/r+IFzfjG8cfrl/kqqq/vWPaTpb73N9
dHRU1E79ZVp/RYN72QRDyM5VsI6f486PQv9oS9YSVn/f45UC3hg+POzc2dDyVud7
OBkKTc7fXuUBB5dN6o+Xha8WGLL8aiGHmer5HJhTDNVhBRe8EpLs/e3d3DX3hPtV
/paRE94vM+aH+oARjIMFLnLV4Ul8SB3kq+KAeywLe1b9KF64DEobY3asfTCnBXX2
dXl3eGn/F+QSGGaAzTAX63ju2d1gjI5lQpSuuPwUmazGU9TVbL22SHf0PVcj1k/y
yMQ0ZegynO3yHtERTqTuH8DlmssPHs8Kjo4/elolW0Tmn4+S0ntOZMM9GEGDxPWX
msxGdXzhJJKB7xsgUq7pm7Ro4PkQuuJgvSDCE7BEmGJwhDdIg56Hes5ark3hiRYW
YBIJUAEAJ7ogl/EZ3YVAQ8MNkM9k9tXNhKv+qTBW0R70Z7xK8HCAdnbq59OrVzCo
Q4T+JRZyJNyvTdxsoMzkDnLNQ5G6dGVRxl9ui1e4aOveAlPKIuoZBtsGU9PFW3E/
UM4ba8B00iUt/nvxsvoHqfnEJElTz/h1Zv9JM0wzcbBab4cmauo39GAxu66QmHXG
ZALDNmIH1JbXY7YzqEc4PzkU7ti6EMBht6l8d1MYuu7V+N44MxweWfWjjpmcxP62
ejziJeSYhG7LeCNaYfBFb29/qiqScmsCjOB/sIhWczTzy1dvIhLkYYqxlpDs/9Xa
9809wSEYAFvrL5vBL2qYCrdJsaXuGgLGtj17rfFUmNh3qnZiyhwvfj+WxQpCTZGi
SJPDPJ+9Jyisqaae5BJouNvmhB+ddcPV6YX6yB+OVy7s5XN8Ca7oMy+6ojphPcoj
9wrUIKv4x8PL4i5otOjEZ9GReNLWvyHWE7aw28mdbfVlZjTSAeg9RehYWfmJnUC/
2WqL8Axl9gmNFCkVBtW6sgk0yoWWkO1i3Ugrs/aNQ5xG/D1cBCYKBx737bxXk5Vl
D3jFVRBv7DwufLVKFU7wLeRTIUN/KNgoAnXU+LJjVyzQ57Fg2Qguxh2DuHkJ6CQm
L57BZ7YPIi0R3k4krsuPwc/9Ptx4mKii/LrwP8xQiUeDhaA0m1J4/BV59gE519nr
p6/clrYPx0Qk4hFtKHeYY1ytHKiLd0py/BCeutke1FpYSf5fcJ/8StI+Z8hSfvan
tMRzqTOk/f4SaMa2XyYPf6f/anolS4ChPFVWDENZ1eLaVXaTtAwmGjpWxeyClc6d
vmXCxTNuiojpcY7twGVzOgvcruyPaakDxBsn5jJ2qjTpR/HIVrRJAf7Ah6HZsxDi
0Vr82oboQFH/2AoD60AzwpP+koPDhONKEB5MvToJOcgLiFMTQ33T1UtuFgFlALWf
54RK4Q18ophpV+SgtGJM6JLw5eK1wO9luXWGb6M6O8bOaJP/m7eey1GPdtgUO5lU
vSXONd0aqnePhEWGHY4nfr4rla0rvuRz53rNOrd9pXC8dyca2Yx+KnfJ40we58RH
0K2/Df1jIL/EpozfppXLurD7U8qudCXS+1/spTJRdtFtbkq7+GJo1ZEeIqVEMHhH
0A+p/an8cwry3Oirv6i6fKBkIadBDKJ9nsEJUuM0OX1DeRQOQO1WAg+0d9+AYgDE
rZBJXoDzSgU8vFl02b2gkOVhI9LADXL+3mhRz44yuHFYzV3waZaKHqlwOaIb5d0u
wsTNJskg/JfO7R17mUeQbAZ6tqxh3HrF65VTs6+6d5my9QO9fvqEywOIeNFsYvYH
JDavuh25Fs+/bTjKXcrorXkclxmxgShAKsnp/wMZ4rmuJx5huCqKNEizYW6RL17k
8+GNfTf37WAyieOMI0MOCl5Pu+tcyrw78whwUvhcSG5K4Lc+HSWWI3MNAwxiHgvK
FmdQyLPMf1gC8vOfKBqWUuJ130JyvEUha/RVpsKL6F84Z2w/tPNZe1ejs4S7xV2d
HJlVYWl36xisDRG6fdnShnotKtA7iRtagYJpUWJZEB8YmhMY8pQxJcZ5+ygmHuBB
b9Qpc0wkpqBBko15v4ILC16bhXSyUf0YxvO+YWPFXY1A6sEE/J2UmNgs8/xg5G3n
le/lJ7w+Pe2hyzxHya3TDfabh/W8JOE2DAoByEnzIzy9TRDrpEXu+qll5uKNwUlQ
elYIAcSt1Q+AiD9rCr0SeSLwNVNHexUxTn4X2zF77lwVpGaMUpMyFomcrxUPJME/
PceSV0rXm9RgTv6uewR70JaOoeJr0udVOH1K8jpj5upfNvHT61Bs6dViyUbk5wNO
+s5Awz4Sv4KeBebAvqGKOAsgrDCHniBTCNOW0utEVUrVKWcycxIt9WQe7EL0GU2m
8o094n5vG5cML1rZ3Iev8IjXTY7iMm9VWpdCxLydr+kkzP3KsSJ6pFWCAoDKDf+T
BPlL/8QkXYYuB1ZVwqUWsoFNWPhjPxGgZDAXgvIFEnFyB6VEXe/mTmk8BZzqousa
kkPBxU/z5mx5iUwYxH0qRdvbkh81H5NKuZoOMeFARDgi075O6qVzgLQqVwfmJNLt
z/4LWNoROFsM8BzLQUCC2Qw+5MgIgDiJyHPwX0IPsp7VN0I7aepaZihaC7VcgVV2
PpOJXqEIj27E8CjxPiQjGuT1SLY2ZbihUHfmD6+34hbhHwXOuLTiZJymXI1yZEtf
m5eJRXN0qcLeVhHzGGDyCzunJTFaOrQyNFAidkDlkWXw8ntfflr+veVPs8ibaZCE
KRb+eniIN1cBqUIbo87eiWakys2fZrZKcyAtFYXtK7eLp7BbQlem3B8K9czt2lz+
MlMlN1iqbObUtN5JIAxCXOwvBDHMhhzhdfJf0ugnGbjm1BVfhT7mZlkiwheTTSkK
SnyFZ1FyzbKR1XGz0928BfHw4XinyOSCdwJ4OAlMChX6Yf+KgcUVAnxz5YNrJ/HS
Ij9f9mj6ObtleaqHvLdZUoh0HIJ9TkAnk3pMAtpX1uUEny62ZofnIVRaodul72zs
UYytMHqIUZVlAkRV8RIy3NVcg1eiwqK29+ygRShEja7ZOD1z2mz4k/M5aB6bGTYx
0977+c9qm8NEG2nD45cDQUzXkVu+/7mKXHnIrIlqwkomWCSapR2GmwPxa+2tY+Ug
ZB6c2paDjjZwRuDcuBOj0RKU95CWK9v48d3m3tFxAYWOqN4vbfkAzMW0vEsmFbJK
Ns6aAX51++el2SAoRiCSVGeTgnsywXpocpkATrL8SYWDk4ZBBLji39O/Yfm06V+O
fHF8S3Vm54FqlJbmql7W7r9QuDtbK80vCB70OtgdZMD862GZnPCisTxBi/0dhgCi
kFIb6Mg8Tkm1t9GRHPom0+qlmpqqyOq5pKfgpD2EnCcqJpGtMZokdA8kiqIKMNmS
Fmtu0E1QbHivx1mKQ5Ltj7Iz37nJxCeV48JBdOwfianURvtK8SBQO6tpVd9ZE4jv
Oa59njUC36Ztv3AN9MvPit9ouTCH8CZWUJJFL3JObUl9AtsXtyqK1T4uOjb2cVmC
5+lmkf8ZrbcYHAUwuVpV95VOrOwzBudZ6ju7PuS4AziDPOV4FUuJfmye0mGfgMLS
aU1xfeuA2NtsbaxAuPYWZGWtyvqZpjWPanJw/6PqUbJ6dbQdwWdKrA1i/HU3hRyg
2WEwzq3JjsAI3KsvJZTT8XOw/lnBfoOMO3f70QLGJtHiZH6r7qE7i/YPhW9wLIg4
6AHhjmVQpNBBIj7L6FbuDcC48kAuITAnDsgACT+uWJSR9LibXWMKV5FawfJp1DFs
Q0IYdmZaD07pQ3Eq7BTzdCtISHLOQJuAhhM6ZOeoQirwtkvkoTc8FRMp/+3qEc8J
7DNqRvyApS6oX01UQ78VjOUkebycVSwtqz/fvaSLNa7zhA3xumNZupAaGkdTaJpy
jI+bdkT1OkzlnLQ2Im+mdqv+A8pvVuT1nraWLUniETSe7sw7qmZ9scryq2MnC23F
IDrqM/QZw20iBwA4dLGJ7I464mxGhoIUgASgxZ/N0e2Hdj7DKXt8fkNmXP62d1uH
K1mopf8BxFKJKTkEMfKzgJNxsqqgU+FEiagUIxbnTyUX1hjc35RKFr3Vcgtkxe+d
NjAnWhMxvElCSUyHOmyykLKp8yKBTwkHieYyOahXOITKO4FMdEl4zUV00jlymohh
rgNox1bBiDdI60pFNLCK1WroAETtKbEZ4dbgEItLSIt9AAraEKDJ0wa26zm9mT0z
rMu3iaNJoryYuv1IncAdKLNM/DJsvWK4P5GM5laLdgI253Pk/f+tXyIj8BKgbYdt
691i5Moe67EMNBCF5iM+tvawj5QaAO/L2uiRE4NnI4bhQo0bqWNC4BpeJ0K4OYZw
gISCD/0IGTbbGy3Re0nTcVyeiclJkhk6bfG2JPSxD/rlgslCi/XvHddgZkdttBDL
MWW+t10ii52bYBIAQRp71kZGeNS0LrZ7Ha3cKOeFonNWmugqWzXwlFgII50seXrt
0mnxuy29bUSctsp83nYzLm0iL0nziyJwBJk984JBrKptLuNcekpPrk4RMq2y08bo
ywfTVPm+20vej7loaZqHGmbfxT041WEe3isXTB3nrj5QYeqgjUCx3sfJqIxaphx8
sOHUU+UDhocCg1GM0vXWU3pTnvh6VuXu06CSTwNoPqBS8TwZ60RRJIQ5JvlnLsAB
EwNRBBO/os9EFVFYMAps3BsWhDoU2hL9mJEzBXoFUhLaxikutYrW4b5tVHoHVHnV
QinpK7a4ZQnw/UeEx/4iycjqu8AiZAC8k0amu/nv9K7gD6BjcQ/Zo+P3OgQJvEd9
GMKlpEg+rU/Wc3dVnpn9Mfg7nDuQxqWs+eXhF6rxuh+Y0AsEwK+7VgT5JCYwtvk6
DBkQpwaF77kSIcsHtXtFR6LGf3ahi2JQN4tLjMfFTWV9uuYYcg+veF6G+YVLKgvH
8au3wU6bHIU3d4NT80pgSbw+gR+UKpiy1fS44tDOpt/1v61Sq8KF7G6UCsfn0ch7
RUKEpWG+lQAgLhVNXE1dQyQpNH38nX+AI6tZikY0nJJJ4Dqbqt00y4AeXxcKFb+k
UK/x6QMSnldSiYFwQEA1KouTfdCPNQQX7OPw16KKUvk8m/AW6TyMJFJLmlGPnzrd
ouiTt6Sfd7vMHcgHMkFowWbBhqTzQ/x0Tbpu7tOCnIlatSiiEibTWLMbUrw09lT6
/vNjDn+bFyGV5OzoUe954C8qrHg+3d6KGp6c/vdu6zaesoWc2n9tzFCaKwAqtc2K
DvP1+cjcnqWzUD19LVEIB2u/T3Q53yshYLPA4O9WGC9EYWrpqFth2LuOy5qOSc6a
hpuipMW94oRumnr2gd2sKQOQhdMmsrBDXh/tkiaiIyemYit+XibeCgj+a0MWrdHQ
UEsI9tJ8G8wMb7VNXy8d3knjCmZImNI0FZirtWedQQnvE8TL3byT1JsV7kemi2fb
9ugfPBiHSRf3ScmoarfRBq/scr5WnFaLTC6BuQQmLWva5pD4dMn/Hw8nW7N6e7a2
J0vJ37rSgnh5X4ONgTL59hxtci/w6cwfV7sm4ymPtRxCJPT7kPZTZMMgEmahwe3T
sBgM5QLAiClDqAUrC1Fz+jbJ6snh4o+4zY/+EZJpUXTDUx3JEOdRUW/g3/JpAeMS
3Zi/3y+n53/mVBa7MZrNohip0BaSrJjvg+QPOVsYCb+3ZIDJKarsU1oJQhgDMa6J
vlhL/rC0DFCmqWYRB+T3FLT65/v4YG+40XDQt+uhw8iHLxffhsGzjIuAzE8spIn9
5TP21TRwkxM0kPeQpH2an2iR+qT/fupsgI88AzUymwf8Gfnrqze4t24rh1YNhlwS
D/h1qO9gnn1uwf2b/fV5B8ExJWdlaIEwTsB5znXeT5jgnLGewWMjP95ZGnEbiufS
f4AOA69qD6k46x7REZ5kVSNQ8a1x8xVlr1IsB0qmvSTckjidhpPdFqd1g1Fh1CxN
tgR2mmIpTXP2Tcw20f3hFjBOFgCh55yE8X2yu8a09fFovFTsobT8MIe+TTtZIiuL
E+LZSaJl1RYKqrxC4PU0KAVq8lfUmQgYYvu18Cat5NxiUq6BIipwLVMSsWOnkaLM
Ue40Nr+vG7Bp0l4NV5LG1aJgsuJD0YhjVcy6i60+yvA0VMKKrwz2yiMIpdFLH6Kt
RQJ3Fr5SqeLZJLAEW3BCdMYtsDSGDUQb3TWlMvs4rEmuNbHSkfLhmpCN26y8hUil
nd+HP1fXD6FXpZK/dAuAfT+QAgBEkXwmZs6hvyjEyuQ4dXnu6eRhvnI5R8pwhAUQ
3uriGk2PcRMNUyLsm393F6BtQYXlbkZoZH0OH26IDJzyju7Nl+LnyiI1oAu5NvOl
NEiYI1QBOqtQ778ABBZPlYPG83XomHfCrmA2oKN9DvmcVUlkZ+yDFDVy+iXLN2zi
NqH9YfHnIxYYOyi1Qn2o0SufZcuwMbVEnFq133OSpF4StnCa7NZZX5ufmT4CBBYU
Qqd/tyQ5llpXLezE5R+pjjoByAngE3TZMsscaQ619KiGzM4H+cwryPe7j+8tdSMz
Pv6xHO3eWSP27T50NLqCgOo1s/aNgkj9AmoT9A9libAUcjJ4ujfXMycBf30ggM0O
60E83X9imDvpzJaQC6cDOpypqpr4Ja8JbuIARvl85w1V6wGmM3/k8ASLF4y/lT2n
Wvw0Ig+pckFmFVsVcaInlRECW86oVMVvMq/0xQGbmbjab8Frj3qHl40RG2pMWoMO
uYvMfoNeWABxjqSOZN9eXwYb41U6g5HmeMPnyFQ2L62Ydmg3ZW+5rHPU9oa8vXMy
vR9ylVSDg5k6uvPFMJGDusn82bnhmh46kZF1SkvfZbJYPTZbHvcfCuhCaKq0jMRh
W7RLjedrPKzO9LwyMFInVsSepjT8/EfntgUENq+y1QfeKgFqcODNn/SmWJkBXNW+
ULTTLjSMCquppKI9bBK8BWJ/nrkLnhrGhRqbD5QMDHK6l6fXTvphm8WtxwJ555Oe
YM/q064eaXIVpLtancE6b5ao8fi0AnJ2HT+gWh4mc7RZlD95OrUa4maUI7fLePVG
YNa0Ztfgh5P9shGKvuX12Wr6QQS1ci2itXte2QYgIGybpJOPgETfJBZV4PHtpeHK
OdvDambEGnDqRNOZALTSkWceq88M3bVWjeUsTX77H7JwJeCfLVN9hY0XBY6srreX
zChu8LE7OAAPL3ApnEDjHCn1UIBiCnDRjczeSmpTlkHJihWQ5gFWUFicn33GGujF
Y/HSZN08ThPsaGAiK0cNioA5+foD3aOl2yhq6RXwTJdPchc+dDO/r2fL9D9IFkUN
WXoDUG8jv6Nb+hGIrpA1yCoZFumr4e6wj42fxp0fLWAkbbArEfOznVsm0Evmqj3x
49OXEjNQwgTzPIZrm1Xf+CkWpkb2HpBrlyjsr4MwP6TbjoKHZe1o8RJ7oCuWMRF5
E1fC+b6Dsi0c0kFJByBeIRJr+58ru/fhEuhq7tSvvg4lUyEE53hlkI0ZrijnGL+B
LZVU1CuQr+gB6iiTmUhlJ8k3nDLm6oNrmJ6Rv4BtZryGxjN8HAzS575kTnWb5ULE
diazsz571J1qDB5M0QiBtVmBuMNU8PalnMSDR54O6Ix5nJKxd4urejHV6mMS54r+
8w5kWx1NYOdXwHn91RmcBSLElSoI6HPodYhXP5ASeEKNPWKPBus6fgJtZxpDBGmN
mHXi/uoXyZ4nPKS6FZ6m7cYQmJElqLsQmInw0650ekjkjKtAj4pUPTrHX+yjzAZr
4uCLI4XCyhUlt1vzX/lFCSOGIH/GuGPTaqjjztNEk1bUBXRLJH3C+pc7yubnegQV
wVhBexuNcrLZee0yU0seUH8nfy4U34IlcFpqCQZk/rBXCGkaZcs4bqopZ4Ns1DGP
3AGTA9n2NWXojlj++NM8HZ4pE8WVVuAioNmOxJQ5/T+CGsL3gckAoPlUPfP0BFSR
7IgVHIGERd2P4Z/TG8Fj+SJoPcobeZ4EHguli5t2nr4BbyJq07VQ07ocNUU4eaKT
mRhcCiW3zzGhumOD+8/uurgG2o1NXtchOfyAl2RcFgAmtXRQzBLJY10lvE/BGPaO
Z8fqq0QiB3jcXDcrWwWSdoJWSUtdn+GY74llvvvOSqqLnXJMs5Ip+me8lPl0gLFI
rvjTw6WY91fG62njhR/0unTgpe1Zoj7ghhWiM2w3dXc4NUdIKdfGIzXRj8wOd61n
irS1hJBFqRq8SB6oBBeVmbutjmg7IQ/gq7VM53nRUPlwPcHa3iGypP1Vjs24iflN
Kbj1EV9xF43bi97BpBdFR9pOquwxF6UJwR7gyYXWXwLrvzWWP9DUgRW3L749zNuL
x3sOUA7ZPqTrgM7LngiAE1LGiLV7HzavXe6G1JGihVN6GK2N80sIM30Gjjthk+j8
Nrlf/3Lbx0zLEz2UTRoZr0tZjA4c2ctAVdU5E/vTeTDxF73GIOW5VfZNpQciat/t
4D99IcXO96xTKEy5n/WnfXk9I0jhLmkLzzA4I0rxdEAnDo3OE6Z5E0VD4Upvf/eO
z8tzUTY7Lbr6o5SnBurDx6bOAMDmeSAkDDHN74lNFI6laDOM2+SVzkzmRs7AKF6o
s+E6j2GPgko+jdk50XKxAWiOZKRvKkZGJotGAGhmYSEftbc6VivLR0QDodIMosKg
l1SumFkJJMgvLT+yXEfbTZlnW7kwKGfXeQHiPEMdTkW5rI3EgTbUQapu/UoMCV10
B6TLCwGuN/vxV0oWygliITUoPQLPk3YCUzRRrOTCX1Z3Iq3frrTfpU9UETxMDq80
VTK3c31XrLnBQvmCkJmW9ToqJY8phh9HDsKtOEoSpoxPbF4ZG9e6hjuPD3O1hqkR
9y8wmBIlZkFXOUxnM7MdCQcQ5Nnt6LMwD4dQoL4dtyOqXuS/ktazVaCWjZF6jbr2
voQWwQrwbl3K7LooX1BVV6xogpI0vJof7f2lKFWWz8VA/2obtKntj192ySsU2E+e
j4dU8e8JQCBT2jB6qvyPAEwf3FB3i1PALNX+2kPsuZqY3+pdIHKKySCA1D9KpDr0
oZEo622NbDzjSRLEPU3AhuTB7XzhQnyZO7UevHeiVh+ZTFq2iU2hqN28P9G2FKiZ
i5pb5h8JOFrsr85cLqKkuQfXjpDcQRw4A7LXfI9OLre0MN2Q0UoUGJEOYtzxLjH0
LQevry+FFCqrDfK0z7N2b2mv8WbUWPmLsi9OjsQZKoYS27r20pH1QPh20t2eyDSt
NNa8uqUqO4FmEFRMykVMFpOLDzbTSCqfSj5YbabxSJcnJNr17LlEzbyZQX2mo/CS
6jAXvhDOxHB7MaqDgjOWqpvPllRJSOYAO8XnjInsSDR43FrSbYJwFuvfpZF6ACpq
fZa3qFIDAdD1OOPEAk0rAGrl83KDySVAQqxC2Pp18E+wW5T18Twy9JSNzcKSbO91
CHt9yyMZko7aZstAnS6wdq4E+Xl+shfqlXE7UnKuHkHwMMPnO003nJDMPwez7o91
XT7xVdKqjjapua5BKJNet2KWbr+hQQTUJJo3itiRvhUkl/IXArzBkpH+ScDUkJJp
4iZ9cepVSXwRFdZEilSRWoL4AL+17CzWJPbmWt/+ReY+9NSImEB4RLihA0FfOnrN
r9c9H3SywsUvMyZBl/LHnvRhL0uRKECok8y//InnG1NCIbmDsU8sjjxZmKhHPhkA
95EOJAAhb/f/tHxImpz3oKAiCrQ9q/xCc13mI+EliNoXIlAk3N+w6z32cydQSGlK
K/OynC51NdoeTZVIjYwaDBHt8Ngz0t8yAA+J03IcAestiDc4erRX/F0JDSDgsCrV
ZSoAE1WMW8lTvnlqps9R+viTibTl4e59uXcapnsZ4U8YyFFY4Q1Y3Zyc0iSvIUnP
pe40GxbA0b8fiHfWuPBDCOW5CqKy8XMHKN8VhhIsn78qXVWuKkrXiU9C3lFm6GK5
MaFs7H82pdYCiBzE1LyNMosZcdC477vXimCLbpw1cUWTJVW4oeIHX7PCEOuiO15J
dJmdBYBSDyn/JcgUPqdUxwHWq/hDVLJ7gzFNlUDpaZ00ZBYKDPtfI/YUfrvJpaka
TcGENzku2MHoqZndr6tyzhLpeOp5PjngULRlFZzLjJPEaOjcZTit43lk5CMSeJMV
6REWZnG0QrtOfGgFJu9Z7rxqRObRrwdm/zzM24tjbw6tuNF9EgvePkafz1zzcYm1
i8++wcAfTMG/jQFgFY2K3ZNPSg5WB7VebbxVAoMwwEO+nfALo5Ln9aUZR03YS7br
SNxAP5veoiunlwa7Gg/DCRDi74Cbi/3HBlchW4R/CHsGUSf+D2Ici/DnONPMNOMf
5OWbIoK9OOMnKcE+8SoP6uaw1UBluxx245MxYPNCIj2W6XW4VjQBv/xTXyiPOw4D
/eZ+cRDVvR/PtMPZx8/MVP7yzY8l/5J5j+hr5R7PlFuT5UxSBYwMpJk9vOZbmBwx
sahRuTzW+LKypsQ4reS4huBnkyyurVM0FTIkyC+BO6QLT1vFiCE98VyEnR5ihL6l
w3lVtrZwNpNvDFjtYGO/6uz20GilPpedhg8WgD28TRV8dIZ8L7VPdQ7YMxBidW0M
ABuYxa72HMPehHE6MP9J0jF1ropHMeOQofkeuq6CLyhMdb25uiQ5NoWuIPNjvFDO
4SymiAcgGWNJ6jEe6Z4xBJp7u8Kq1/cfuWV0ze+462JPKPiYLXXNv4N+AV4EM02s
ow3OBq6uGDv61Y6gk1Edn6sT6lONJuk5ef28McM1ZPGAU4gi4NPgSvOhglFrL21M
VvVa5eS+9TdRXec02wwotaVYzzq3uNajKQaniNfxCwTxz9evV83+K9guuaVeGo9t
x2b1Xo5V+u6rmCTjPOkGLazRUte2erxoyS0JL0pwmJ8BGVyH5ePSy1KrbTdpLx8K
37Pb70H5oNekVe4+8XcU7aPPqMvYBNlOJr2qr0hqyeNEhueg424Qa8dVOtsJUpsI
ng3B6G7AZQJIBvn3gP65quBVb/IaKnztjQgk2hoOJ+KCxkmkNMMYf7AHftlG1RUP
ZBGMu6dn0DRpTqywQ/eBGVukE2pPCSTHIdka+ro/qfCQCKDIT8ThBJ6ezcVJvHXe
8egSr0I7TwGWvMzYSUO3TLr0pv9Alum9wbbw6QrrPxCZzJsh5/sNHRC2Sb+J8Bxj
904KCQPuKuQHJ8XKN9Qq+ijsviV8517Jvo2Tp1zRyD++vnqzK6WoHGh8e58xy8c4
NzxLlLRKUeXvX6GY7bory65YTGtSrzrqws5S1kL3/jbodkUt9Bqy1YPN66F8mtpW
W7+hBakVlnwPlRdOdBUBa7NQ0h9dlJUw/+N5lqkfa7nwF3Dtq7c3G7gM4LowrrFz
2Ur/XB6/efyzlXMEfGXdNoiCtzPiQm8mxOcL/c+eQefqFG0Aro9xBuOisvWUhlje
GBzqbiCpwruWCbkVGw7ApuGSn6X4/wNiZ347N8sykqGIugJEAf0vb/CostsTRD4J
b3uZaQdDfyFn5rTP6SYZ3EbGjGvSny3hsKOce5i3BO1ZiA06vqDGkr5dHmLrLqDN
984nciAdN6rgu5EImdFt0XgQFEE5FsQIFyBC8V7kde1IzLCDqUWPGVvgh3wPFJIp
ehvlYr3nV27nRk9iRzm9rvtu69mAbpa2asNxZ0RMjiwwsJp2Y3IkM9dQ2QmL9xie
eXhEknZF6l3Aq4HM8Eql13gqbqKcyDUod1hIbu5GvK8r//m04kjubemE+UrPE44a
+zcmH82+X08+bK20UdkCWc+59C0HxNavQFkURE3e+wObU05YHsksxvpRYveawNLI
SNYy19f8x+YjQ7RkOXOfRJkjS8+OwyWsoePRiyL0/9dha5ArbFNyl3Ozka/VvOSr
OBV+YwpFJRMjipzpaaymEeuvEytk1Rni9OIC7O88//G+uYlNc8XgZTaHOzfIOd2t
LKuPqKnxjwdW3LUVUYjE0FJX28MSRAysBKrCwm91094dii8aXPoWK8J7nZkO89Ha
MctxM3cP3XBx8ojBBkbSuw1V9ccPqb+Z7Wg3/FoQKOceimWdbc52vCWgpVAyrGMW
QIgzPwGX5HPJftxLl/2j0Ia1kqAt5Qweb9dwGjCuMfKKGF0oZGItdvVkD47frRcJ
0Dl7Th9N7lzVOkP0napikUM85Ldy7V5Sg2gH7u5xYoSVrgxzLcVHoHuaGFS7Wx4w
j+ponuBRBUN85MteCNMlmfVOwpYRF+2MkBgl52C6aKuglGFBKogOSrdefrBibTwS
O5Q7i7sMsTAWxMewHKWSN0HdyoPB5Fz1vcum29hfU90hSZfz1WIMZyxW/M8cjS/K
RNyP4cqzVZlggzVYmy358JttlHcTF9Gf00GeLgKQrpeNKquF2kG55E8vmg1YTYLF
lVpEEvAjRMxspk9ctqpqNAWeKZJb+Hkk7YDmiKGhOqJGFmayeHQY7fVqYLIdZ68C
2/G6QnHXqViargQCk8tSgRCZf22R1bwOltq+/2J5LdptXNsIPiPmVQUlesrabY8p
iVtOKLbd7DsEX4jKw0O79RGcKZd/OLLhUoc1ndrAXYFBRPHOHcQxc2SMhvOdCXrE
P3AhxMWf/+JgZM8hiBLDvJoZSKlYm9Mec2CD2+GegY6LZMjrjI5YzaEHDogKgrGX
GAQqnKsbsEhClw1zHzvuHm9R0ddfKmHmEU7qrKGBplohSh81s+MgOb2lvwrBKzP6
OyZ9kTEAf1rgINLiyx/1/tkL3nIIOsIjNjgdjt+akyfwK9GtOi08gRgyCLJ43uaB
xufkxtZcEk7pGwkdBV5EjNtUVsE/fRK5pVmMkUPHiBm4wNE4pSH+LIU3uXur6zHv
ysX59j7wBNoWS1iyuqt955vwkUJo8SI/MSMeCL9X3DDuM3kIXW526dnbwqY9YgUF
Ud1u90bVJB8L9sWF48TEeqgw0EDznJ/hyAZPTjpNrKCz0N0oHEZaW8wbiOteprfM
AhcCmp5WZR6FmEcDxwTJQ3tTYont739YCQhdqEOqSJRc8+Erqmay48USqiaVfX2v
1bLXvMZYT8c7uTg+oCMgSJ9SR72KZWV3ObwaZpAKJhGLyoBQgHFKjAorDxMxU8P2
skgL9m0c7XF68yTRKhk9dOIj2KZVtU4deE4GHTdzxhJYfVD1Za8Fjrrz4mlQO506
+s5Q6Nq9vvCQBgbZWBRCryBySBHAN+xSmCQRZ7REKACgQslJ6tt9tfGEcrJcNWqU
VM26mK308vUzU4vZb8myHgLSvAvU7d5z2Z4Z3b8gwuHQ2zzlDDJlwvpt3BhyBh8i
0I/O+BrYk4BwbytP1E0uI7hoIybS2Hst8xg7XVtf79szBd9AxevWDMchnono0HHw
WpIey1873vm/hhIxiYFJE69UXV+7DsTCnf0VXBTZ4spFhxs4X9zxskPbugQ/mXuk
tpAo63L2d4w6IgGDE4PmXW98uB1abDA1miMgBcvt03OkqJLCYkoMGPdjmKtBRJR4
MHbTPC9o5bVvzVc6RWbKbA91hY78bfs2aZIhB+qm/4ud1hqJNa2SaS5P3+Vz1Vjk
M69UVu6NgI0DAjRRhfBhaviTyghKBXBlRuvYuFBaRQK3e2gKpJNGx0P8bJpR27Yu
UhyNEWlaUuZEq4kAtPB8ElSMBPh7uR/LopnaGvImnD32IHLhu93zHA9K7OWsqmBJ
3L8G3OiU62BDvBjA6mnaciltjoBNi6T8PPhiBsSoJq7vrYdeNQRwS8hmhZqZ+KP/
H/yRl3kAmCZkNx7mzFOkskV+TU8DAmSRDM7n7sQozEa/jcVB4/xB024cjEISTMM5
SIGcYWOrT/S+5Ak/ADuDlMDMBYYCEZlEoXKNtSJPn5KiyGb/82okXBXSBZ87Ff2s
AXcWolXjLAVaXWpBWduuwmluWJ9nvi8JXSabt8LrSuZ6IYvDw2L6XRasPYh1nsl9
9VRPk4whVBcjoNgw8nuURFknab9pHtDdKnwc/hVVPNThIghiF6jN3ItsXMqyNOXO
I341D0SmyBxGGxbELt8KAlInVNhZA4Oya+vV0cOeUlulRoH8ff5dN8lJpYkCYB+u
jB6qA+vzb3/W146dKxcU/UfKAo6KFVi760SazwQbHAGw8Uib1bklG5jwQpYbkxq3
lI/u0vOTA4fwL1UoQZ9WcYCUX9BDA8JNplXPZNekzwiY9bqgQGQiOrPITo2YJrQj
ZB+xaP6soDdK1ZxvJBYn1t8Io+n9caVfhmZetnDu+KUwvz8/XIHQO4lwq4Pvq8qx
MkB5wFDocF7iWaptw/ruw+kUqHCy32+22baD6PMCu39mRwv3WL6jFYgp6Q/FwmhP
bsJGvs8SKT3pNVvdQTelpe5Wod3Djqkk8dCjDTCiy4F6RR11gEBQPn9xamJ0yFUW
wLQkMa3rT03oFN/ffkuJ1HeLhQBZKpwPLZLU7iB5fnwzsth59vDGjJzpPPwiKB3h
Haql11LGorqGpRaV99AJzMF6+qXnw1xAAK5dHTlZn5gjKpqoVE1wXfENQ00RGE/y
vZiBimyO3FFseYz6qXf4G6gmpTdr7h41g+hk+IeI9QIwK5zwI8Wa8vxfhHopeTQ7
gZCuvIQHrMQUxDfwp1H+sCkLUUUlcJpxIYbo6xz68NXMeqbRvNTb4JNT7UmvrtoL
fCdyfRKmc5qjOCN9/2X88ZF7elu6uZscQ/GKHY5U+vsvEDer3tCWWwZvok6CiQKA
b0+uUVJ/huq8qa6kv2WYwRv5dsFpy69RyjPesywi07VeIFC7gwA9w3vXroG5lJt0
s7Yca3oINZrwtQdeTWmLzSkXphXrLyyt38EqyvI8XLsNa+4CzbT1Vz4QvQR6gA2Q
EFycjr93YFm9nP/vWv++jxdpoOj8JQXgtftj+Mjb81wEBA+C1c2XaBJihpiDXRje
BJJYp7q46Qbqu/4XD8buZzDk+GwQvkb+4sOi0gfo8FUM0PvXnJcKjL/CR2qc3De4
VM95eZd3bzA1vFa3QIZXbwnLuDJqXggNyJTwEiJtejFIt9Dy7i76eZPwly5lJSH6
N2QrD8L7htR6Jd2bHVHAPrM1OZW6jSVKzSTNWKsoIbdOCWansKE93iOJsr05WRQV
u/1sbZM6+lObgS63mQiRTa2+p9lkBhAwlUnLMIoDAN7SYA3vmctpbRZ4Gskcp3kX
Nsg0wNST/Ac1lgx9r8hK5qLtVMc6MZSzSdbGIAxO4gX1luZEOTBeCMCO4FZWKBGj
T6fRL8945/OcUf8mI1uFfdqTOy2Nfupj+eBshxQEfiVgzG2pFmR/nvRbz9+kRazb
4vD5TOISYMWdcI4Q8WSvSJp/XNnBrorWO71j/3L84vZszULmk4qeljsm867Okx2E
z5o8x4yz1HH2bQ5Swtrxes0U4N6IwPux4Kh2LV4YeJkBcxFwSdPYNIPhNRiQDg3W
lCMCHijG+4HT+PtwRvgPGGvAWZdfSytUOGTB97yYxD5xgSfuFpMbbzgT0PINoTGL
bZpVVShCuQM08WAiBbB57omAczSE5KdjzCiZ2CqmEk1a+qvj59FKT3vVTwLdx4dh
5ZJVTChfuSSK/eHRWZnaMTG2J+ulBReQhF/HbhYXB6hbKWP+ncDzeGVR4UZcjixC
XcSd9vmoxKA76Y/KQWz/G3mLEOyJyXUyHL7yYshy3Pl/vVJWpTzuAOSjuosEjhqR
dDJKLFmO2AJVbDc+IsYUA9Qvv5DjU4Ao9fWe+Pzn7Vk6JSyM2rLmRoBRfbltGmuL
WvcsgpsYfyKLUx4T67HIwE1OUyqtlolv8akIEhMOBe+nnJF6r5X8wUnvQ3qbxT61
6o0nQQ+VaH+eO4ORZM9lf4JfCC6Qo5k7QgV2ckVXsBh2KXzumUc7nQrST03UKBCa
JXDSwgADZIXYALFxXy/U38tq5sY2J7fi16HHNoK1fK5BRSKLfPl+nirLGtonoj21
zOMEJIbZs7zmVng+cdTeo9rDT93fRkjw0zI546T2E4asuRMrNcSMd303WEmevFiW
2f3Ve5JI7atf5HZt4fsGkpFcaJdmfWHPNAxhz6vGxfBEgB8qSUaiUXmHD90EdbK6
JLToCUlny0GyDC9MmZiLjsj6Aqkl5oNBJ4Xkl/ffUzC8ZWJ+Zm8/HC84ItbcUK8r
sCJ+QANRQUgbqbvp6BzJsnFWfO6bIu9IpC74GLUxRJ9GDvfnWr23ZXvGtJFSCG6n
KLNEEBROwFYJWVoLefOXd78sD1Wfj4wygMJ4jrjtTfe8QySKmoU+pF1DZVUIgnCl
ZvDDZa0W5hb11VbOCcitBESWrIvEksvsVUCUcipW3i7YcauZoCTFgwkjQqwC7ErF
ySXUnGWPNDDWYwUGUIOvhCIdBR7NPkJ32++BQcFJhnJw/ehbYoMd5l875KV9fhvI
64mD487s1hUW9u2cEH3hk3vnASUUaKT9rIeGcEjKoyxyWYGofRySHMuMjnxJ1wwh
pIqRYZYZH7wIbm9p7L+fZ40leOabeGFnR8sPA+CPqvVUxteLCuzLO6pNh1S2mxoA
oPmNlt/E4t70PRaFXpPdfd5YJFiBcw8ONTJGWItJDCziH8zXe8a2pomfN+sOmDnV
izSXHvm/tlwurO+VnS0pF2K3AXfaSQLcgyXgiUjiHCZCu+IuB8Rw54RRKdwaOoJL
pYQdNuKf8zEGOGp8MrLzRwWxz15smdN2/DTYxMtNMVeioGUE1XRSQCDERBf/Vb6+
HHLYmYmtzCbfvgnqOjc9/81OgqRDdaJDhmeL8iccdcj8WV0X6oxlNRJKL/LVL3An
DKlHLzgn1ui03qgRWiZLZzYO1uMjBBa4QeO6+II695toigzYWphTvBDEirxxtSPd
HTl/hraFjYZjZJJ5xYybCbNfDEt5ODdz0BbUFYortqb9U95qT99Rdg4cC9hS+aYq
cDF2YvzBjjUuTszzzeNBI3uwAr3k7PWFofZ5WZF9AnSQ89Cb+ro/+Sm9nyx73TPd
zP67BpRPKddkDdmiv9S9iRCPBXW/LDNWLUXJGwy5skaimbqmC27JjK6GS5RdeE+H
MsvlT66ehAzRcFuyY/MUUxprPNm0md4gZmGEu0aIHM7KvTjJ58SqBU6YCLFVUSdD
dVbD+G7X4UoCtS2wfgsWnXwbdYkN/YkcIIKqRSiGNQH/I1GX5jveMKnJQDq9L7qa
LqqlKCQUq8tZ3PCTUtn1IsrjGdRQHuCCYvhdpodFqIbXCqnI53T5eVTPd4cXsDjx
frikUFOrhbo1KHSut/rc8II2KlpumdUg2flEE8W5yZ9EtF32WnnNRl6hcPeojLem
giGWyHGKSm71840aXhkRByMFM41swALDw+vnHpJ21n4DDIX11nJQjbLBpmRAaYEy
tJ+j5GCcev5rK/uzu+Tq/SmztIDnCtWSAvDfwk1PvmlYpy6idxhbeRCe4AvwL2+z
MdNlaeH0MIw4x/P9Ws0Vxo/N/ne2+2vw3o7Uvy0rkUrgjNUtsFm8sIMoPNiN5Lfc
yvzazBzfmgErFF9wfe967omXw/NhkHz0ZLaSbxf1MnjeBTXp7BLMhE1bL8DkVJiO
8qj8JS9BveDWZcV34KeVTt3R0nPj8HAN0Eqe283+btLL04JD/wUunR6Th8F7/Xj6
o5JWKsvTjTtKbqSe6sCHp/9RrUvP2yFgLcgKTVKCyZ/EP+1DqG1DXu3Z+WP8VxEx
XMAzVnPN3isuWqX+VhxAFITkwShwDyjatbZuyF9904r7uST9XYIrrX+ZsN/4g/7w
ZNoPvkAg5yjoQuVmgCXEDENyGZOiS5X1GWnSxfN5grbqe6FrgS8bexiBalWZHh5w
CTNn3HycbWN19kGk+9G4iMBQ5LLQ+AQo93Ps9PJ9pVpfh7kRfLiDszuTATIH0p7R
QF/DdolZKYdxK0/FIPiSi36O1YKtE2fsJuJ36PTczmJCGp1utThusNxtP8G2hEEF
nj76zP1phwul5X8pbe+iG25OARribmGIU2+vODD0WAFdZXx6tXdpT9RybBxxeUrC
uu3vVAojva6DRPlEEVcEucatIzfQwBqSTjaCFR64SIXYboHIq65h6J5lh80cLYMe
7k1XgaCODELaEcd7q36hzGlx4VYBgI4IPLxk4oZMLAmqiDmJEYSym0lDbQQb/7lb
Bra0K/8QUHXxelEuZ7rh8HREERPlicbiclegdsF1uQQlWwd/XdaGyHT14CCpLpek
RaR+2BxEajHe4wvLYXzx2MEvk3lLjleV8I4eZCieSAunedeTmOzI7CTgwMptS+nY
7llKg4Jv2t+kVO3pFThcqb2eNeKZU4roYVDM5N5nd9LUhu7V6WpgHsY47PXI+L6N
RVRW7ZWBZ4CHjYHFg2aBxRFLZGceFXPe+faSq04p8WWG5Rdw98iQL0fESNZ0uTWU
WNE6M7TR5VRNIx6RrxR0CfAlvZOvinh/D5+1EDlsxiPXQ+jMLnkAeI2fBq0pYcIH
Tuq5Bv3mAjw46tND+nAR19klsuMyJ1DyhrnXGnPfUOATx44Bkse6e7AA81wIIikM
USAIU0CAgYjq/3ubx/uNbOPmgSxliq/BpjLoZu4BD2YEuJ5cdgH+Z67m/bG7IleN
SSa89mYg8O4Bs9mABNjhllyU7X8L0e+9tRKPfSzTX5lIZUQ+V0GYTidvrvRIMCtc
wUmzwTzYoGUQrTv/FhoagwMvfZYrgu+SO6TU2O30yX/Y+u7HFmJkvEDfX13nhOhq
HiM0MXdAN138G+p0o8OkLOxjJTnf3P+cq2p2iGqdDfknh03doFVb+liTQq9qe87E
NTnZkUpIJ/61kKlXjeo64mEiiWzmPDK/kYsP+irzJa+nEXvPuhkk6e6I22R/swmF
RCLLeTLzmcIJVqn7ocIULpfyNaQGJLH/6aMkl0ibglGbrsyxsiufhoidNcuSm83x
Qq9WmeKyZJ02By3Qx4EHnzLuL4eIOzsxKyOkDbfoUfIa4b7Xz4N4kctTbd0mhnxK
9SV1frd6QHF5EORoy6pb26IZGabTaOf+KbJTasoDfh87SZQnq0caAQC58fGfr+Aa
mxCUvOtDcPZXKtSgEZdAYccdh1RfcR3Gl0z0wRx8VqZ1avqsnKSeSJB7XIRyclRB
tJHQPmgLw67wMqmqiR9s2Td1M1KLXAVf50g+r+RLPn+PLbcnUoyK80VScEDr6Npy
+pTniEB7L6cnP/HjixbcggsVa/Bgrbkpl8KqbHz/ZZS40fA6pBehtg+kZTxl2m8I
ZadCNOv4JbN9usy14h9YV66nkLzsoFDg5GRVi1STs78quq8jilhgqTkWPeasapnS
a2kNnk+LAg4RnohGgNGpsYlGK3IPJB+9QXnkrVmTsPTBmv6B3JGfI/r9Q+5FWvX5
cC6xhDzQt/dkUkcvvk1rCd2yQ7IiUVRPpITu/pUejihKus3giEDw9lbx7spsW9/g
Bms+Rzao0SFZY2tXvnb0RfsrWO5Scrwdd7dA8njTaXkWuAuL/thZgUkz4bIFdv7y
igkkdN4nRx4ueC6uCfYI/NpnuXWcGbXHmrlhPoz+BCQKedQkx7VCpVB1GtFW34CH
vvA11V/KjEanu9s+CeJ0PDRH7GlUcjR/p3Bka/j2EYwCGx1uirfyTmo0F12MgVz5
XsypIP31gFY9/gHoggnHMwHRYmQKQEqFJOuQ4q4RUMidjyKNbZWoHk2ytL2IS+vL
JG/DIg4pUY78XT+d6LnIsbPy4ROS3S33h6qDfYz6x/5qajmcgb2Uwn/hWAMMjyXS
Zxvk1Ab0SEIhNKh6snZWutArTyxkW4tb7A7784s6fM0SFf14/qVNzemDN2JLRXlh
LIF/jEOefmu3c2sd0KMeolBu/zzxiaoRK3mO0YswJQWwFcN64V1EjYo6forBrNPy
KBkMuA2Qra48pbwMnZfQ7Z6zXfB/12uXSTVh5g//AbhUSVI2qfjox7Zp92ZU9Olv
2jk+kCmUvJj6ibSowpAQDkApZLbZiP/aMu2+9urjfjO46OPcx89dG0lzjYa1m0RY
fJyoydWkBbiOyv5AfrWpe/nzy9fgIA5ENJ0S7Z1Pe/JrF07ffI6vLFSKCpmPifyk
hoEbOlFxApgBdqya/rXGMHEJnS/ez2iGmGaC4U+QtiDkdruh4FzawRhwjCkUFSsI
Itt7hm8uldjD7lAEzNijkakptiSD5zntc4vnrLDXdJygfmoA2FdTy/OTR0LiLHpM
rV0ZGWtNBzk6NW4OrY1L1R5emQJjc0YavY1lzAYDt9E8H8LBjUJq8Jsf3GSQtOUU
pyXkHbMygCvfXIX4bYTPFUhsFXCLHAx1/BM9rp9n48mGFIR/X+BQnYHXyQw0EMVP
rAXQh7c6x0dIBhIxAUv3zILtHVXr59PmNnR+OXSvJSTdz8efp1nOgLckHFKlR7iB
r4/iDmyRnHABef8sGaGa/wXKeehMQ7RtU+Rldhgie2bf4spBN+xH5hS7RuwM3kza
7caogLpMT0BvmMKMGpvwVg8aNdj8ygCpaiGZ1nStIGZ7MFsVnDy1EgzwUX9B5BFq
4YPSBr50Au1kCLZEyCafUs1IxASvYrO29Ad31hG3sADwLRB4FWRe5nJleppGezmZ
KQQNwbPIqUESdZHz96J0+o53uBc7hDdozP/BcpiCFYZ4e7XXW4cNiNfx19cx2AyX
LoDRHDg1jlupmk6w9ATf7S3871oOKeOtIJl7DVly7d/XmNhWd6iZBjItjW4V3KtJ
BNeyKlN1jjxnVx5t1ZBgjZDIeCjKIMCcjcITAgRSPRUf5W583wOCOCSlAJ5s3keA
a5YbwrA7X2m402Z/MyVh2TI00dYJRatu/EUG1g3VszpfOfdvCwA3VIAqH9TZcMhR
+v+e1G3L8aJ0t2WJh7GadjBB4DC4HTSO9des0miq3WwQpGMsDa2ZFQzqPJExt5rd
F25JbW/FoEhqFa8s2tTOlHXxMwByL1ujCnZSH5431ZZoKM+rKV24+iAn+Bpd6wOB
PLiw1SeAn9aenOVT59IiArI7/A8Luaa0Wp1SwL/GeuB4WUPxvWhFJT522Fzi1x0r
s/v12zQCW07meKOrVOqGqWgsMacbwOBYtJ0n0GFVqIrEkVWGCzjPQyIen6SV0qAV
9VS+jCppwhlFhswei2lVhSzT6eLeFjxWFhS66ldotwLHXvMs0CbWujB5U9EtA2jE
1MTqHJEv+ueg6NNpJS/lC1YzB24bbU0TO0DSaJYT7QHBklCxvDxI7L/bC8PIpJWz
A75fi+zrwOlMjvPrVKpE2f8jlLzoUWJrNHE3iP3Uv7GGct8chKEH1jXGg1KkCU3M
m8uK8lalM6Qbk6O628hC2r8YfG1ECwrOdUborPVLw39vmp/rmnlhUDuRTAqtNYX8
Jt3vbeGMKyFuWMAHGZUYfmwDNqAEUcQPcm+pccdv7O1ZeGtU8XSmmPomJHpMTjIB
Kzy5FVS7cNwbNkWzH3945ilwKaRSz/pV5giyE66ZyHc7C+6obsIeSH/+nEyXbtXQ
Jf/0/qegAIpp+77QDshAZ3DAJRvoXxR81jukgNOgnno/+mnlD1HSPC8/g5T7pQYO
gsTMiLT4i5uDy7r23wUpXvoxYK94OT6hKuSQjvIA0doldpvqhFNKoYA5oyRaaBcQ
rT+F7WbXHXA9w7wkJmkxjWzdoafhWwCzFVVPJ4rKhZmFRIStQT96wcDyffIW4F5z
aHCgD8d8gIH6fljiHBkuBhdH3noaLZs8s5zI9qhPzg0G/6piV+h/ktmjmqq8DhEs
aUehkVWgvfCHlQzTj+UTvCwUnOmGLjPnmUL3Acjo7ajAwtWhGlBw5+k1VqEgWLTv
jjsd2NWM6r8l7Okozvwp4za1iiAzOQFyBiIMHG6RkUkL9m6ZkRxZMX2hKEDsEb/o
5CplQH/0CQ4OK5WzcswDI00chqVDOUrV2lTxXiOMpOPguDUrUenYkjrNB3o+NMZk
rvWE/PdiXbG6M9B6CV1JnM77aF8+S1PBMREBP9o9uSWa61ytCQJoA1dmaqiwg7Yh
dzGokDF/MCMXdNDHxDg/wxsCNECzDVZGRDHeMGwYHHs56eyHVpgWRvBw/f4nXbKV
M6xwJGGcntJouUBTUn0AiPyMzcj+lPF87K1eF1nYzacaWJrWFealBk0PqLLfRxfr
u5+pdNk4xgm/QqRh+ZP6KZs3RmQ+UU/ZDmrz76Mo4Gg9uxeQfxyYw6KXVzU+XnQ/
Fy5BHXO6IwXIu2+36CSzfPg33mmkwYm+9TVXlzYNeCzQniHyh6/s82hgqvQetBOk
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cMfPjlbsjkUvpRasSNlBw+I7FRk3WUXzYjbiaFUdBrL3l2xMJ/ZMJQs65ZggsLUP
7IsyoqtWbPJSxF0N4We4iE63W1pSyWyg4afLDxC5sseyaILw83DsAbMtzwvz/iPz
vvx/Ccaplq0q61FDDEr0+3u1lDHoQCuSC+n4YSAJSGq4TuCrZiEnezzOrNYWbIlT
4eL65pDJBOT9gnOYpicwtuXB4KYN8vYZEiBh0ojl2ay3kVA7TFc44vta6X6GAjDB
/qQeK5eLOQiDhRkZaf9Gkd95C5j9SbajcEL5jhwfA31qCm14425ohLpNJPfodEo1
TVJjhN4EWEt4DIHNjpJnag==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6496 )
`pragma protect data_block
bsgD6ZxXuND8l6iJru8Tn/LxkIO8qJvqI9V31Vsp/8qBIBpLxZBtogDPVO2qywPY
a3g5oDSybJtN08ie9jLTYfBfoVguLPMfHJakDWJO5S3ZHLgsauaWqbuY3de4Ni3Z
c06DpVUx3A/Al/J8Um2gUompuaaK2HjVhIRzrKkniqvDKdhdffD7q/2pV6Eg0eDP
yP/K9xpfA5buSiljedZYlPlslwy3DpPTFAmr7U4z84jFYqk9nOYEqIAC45vtHhM0
UNZk4mHkPLcjoKEaFf9/KrJ8HzLALawx542CH3rm/Pi18eC1FFdZR1bxjHXd7g8Q
IwEV5mXZkCo7QXoqF8FSwoL0vBwpjbAT4xJ1rtgpeDnGNdS4tjRY7KSzq41zk1oq
L8jpgZm39QWDtuEn2R206RACJU+F8ipLmG4DNBnh/XZVPLm5ZzlxyZ0eFc5b/C1G
YsP/UTQdOknvduKn6VxnTxHDBrO+n2GiEzKGFMem8rq8sa9BMmIr0S6yafVcI6Qk
jZsgcLKD6s2MG/VTlm+IhxKpyc17yyIk1IszEhOvrEFO9XLNkItuGJuSKvECpeUT
7ZJNWl+Y9UlZZEnI6VopmV8PMGehZPSHioEabhjuAMgQA5NfNeUP/oM4JlbnMNZ5
sdJSKyVc8N31xHuRZcxkz+cbzVU9oELObvcOhEerSHVPGPbRLBahAjs1AnfQ9i3R
48pG7QIXdngdEAbCm5jSP2oDKdUS1uaa56fpXtnAozFvYM8hwz9xalYtYm1PkGIY
RQKW9qII6Ywx2Kg7mIADg4Div2jO4yy123eRD2zepfZqHDGUOPWvodXIPo6O2c/q
vupMdBCMp3KhJHnv59vy9oWaomeXpsSToHGNkF6HBjIpIG+VhXCefYFN71uFCp0z
IJDfwOa6Qaw8AVQl0ts8vcOR1Jq0yrjx0loQKVDTNzKxk11Ea2fbkblFqjadEZ1b
8Sxs8llOIdubXArPzGJlAF25BvvWEwhX2flBFUs6MuGdRgB3kfxHVZq5QfSr5FJf
bngtlZubgDOugYMdRLP+A4Gazz38nNWLXoHc+2Zbkh4X8dBqMCXX0rjr3CBDAp65
ydFqC5ZiXhHmVSolZgn+J1iMilw1HN5xq//4DBEoaepFeJpQHHNrz4mEx7rIyuNa
oEnYbh5wu9ExpwaB9tGNZEoyvGOwtss24L5LW1VLgctPbY6flyDUMPhx8pOwblCo
P6VY0dZb/H3RQkLU+GjOdnfFFB3tzOMWOYFXXTEgjRf98hg3nkN9FSPp+QBvuppW
Fsol5sgGKB4k5kV1yAvAgiFxCVkB5o5nlXEnK2dRfMqzNYlJJYL+nfXpJO8uRfA7
b68CX0TKPucUzNsRQ1t3YmdFLqMb02isMuE9Do2wZ4MO3HKsi7uMcFKTch5+CDh9
QnDIqs4nN53Z7C+Wz8bxQ54sa41yD6u3tUj3gZg7Sjo+LJDFOYih1uJX9lXh5wIG
NBJu4wcby4xasqPr4dL+uT5MFuaVo0d2l19hRdZYLT4WvLjmonCtUifR/CndP7Fr
xmLyeEdkLp8lVrbuaRfUY6gooCbdbb/DQy2ugQ2xYCCsBO07gLEq8a3CiJrxAQ0P
dKW6NcLxuRb2yZCgpzeg+auvWr2Tp8H7L47IMdjBDJbu5JmdSfuISHLt+R4yMoIP
j0hHEkiP3L+QaB4GQXXU0YkR7VVt82UhPC88DpZXuPvGNwB3Ix4BBh8UesIRgDTU
1if+xvpKzZvloS1waeNwJn8D/XZJ7BJOlNr+4Jgm/bArR+qaAY1mV+EnDABWLuEi
ohFv/P2y/sK8VNGItmMtvXIXOFxVKCeTyR/B8N3iu5TVCfo00zE0AwOJpOP74eDR
vp1/uXEa+9mOSScI4PqjNg6b3qptF990GnwR/ayIvP0JBgFCQOF64qzTiaisWHeV
GrSre9ePFD+lvSumkxe2wUeRA9X0xwLfB3Tfig1d9ELKzVlp8Hz7erlXD+AwdgU5
khVgXoZR7mToTSI24yU8Yz6ouGHBCggxYCKE/InX0gpAWEX/c/wLNMIl0+dnAHcg
cE3h9UCe7yXcklvi8gYPdimVSivD6XDHP2/+DAkpsphDzzdi52dGdCGcrsnvQKSS
ob+lCd4zQWDEA2PoJSLs54D8PcQjuJn/VM7pepHsch0MUrKrYsPxCacRkw4Z/Xl/
4yE1thGxJrn/D1OA9viFNa5X/nWxLntlXQYHE96H1QFrvSS9lQHH67RtKDGxADbE
ILgApDQM6MtPgKsDW/wv5z+X6e35jvPoVcB3iYCAdYjfvJKbdpNTrrVwBSclppCv
HcBI5gRfAPAfySALPy7z5mUcK/7K5Rfig4NTk7Bkdm5D6Jj1zIM7XKpTfzMe/uGN
dC88s3aZ9ldVFed/yRY8eNsVJmGyx+pD+2CP0fi2rWycWIVRhf5sweD1s/QBs6lP
pc8kxkntMQRZcblhlqPDbBE1uLxakfbvuv7/yDWDqiG5bDhN4bj/Oh6fziW4oXF0
oOW90Q42/RJzndFyflylEbEDBD0yUEwVxL8AAw2KHMY7/UlCJ0we2uqsveO0M/AF
rKUG9n/N8s7zXJwShFSZ3+JrkObXwl95qu37Edt43a0+Mo38+deSpiNL+VaTz1ZJ
zawdUdwKDxRke90GXohjbJF9alSn2T56PighHrtq9IMyyPGegBFqiqohQ0p/veim
iY7xJVAnkE7552rbZTypOHZM19mTnJQkxCdq0gI+Owj3DGkPS2x4wc5Ix1IFJjFy
8O3fJ8IAk9E+YJhsnBkXYeH296puCQXZnTWq/lRD8crdXd9ZZouGNXUO24HSHifN
uSvKqFdNiVi2vPS4EKO2rNDAmHO1NJHLNx6uR+HUbE4vphUm8SFeuuaSElPD0uao
AhhMxLnHVKgvD6KmpkHJkYvXPKRuBiW1UiN3QwHFWbYaLA+fwOfDTBbzL7CzjeLT
+i8jp7gvPK5nZGcTSPxfoxBWAl0rkFUR5Q06tpnZ43LXAEvQUP8yn1y+sj2s6axQ
XndR2rNKaAbmUkPMXYS5iFVB7xwLbk/J+RsrACvYxga6AchO5L8JOorsSVUib7xa
ROF8zaIWSBUEAAi59cy77K/rK/HK0sH2j+nd8ZOqoL9ZuPLbk7ff65z92i7Ms00n
8uQaZW3ZzkbNRD48znnPAVe+ex4FPaYeI3sUrjSJDDqu0782SVKcSC3ZLw5ulC3W
gAIP7pC8dArbHxjOIRjOX+5UARxbkeMSl0JoML4+Yf1198sRvJ6EsZlqZoxXe1cT
gruYI7Yklft64gRtaGXI6Ls8eObXJeTPeYCuSdKbEVimpHvlPkHQY4L/muPKAtq6
8xkpYWYphjI1p0C2PUJQ6mnTBF2b4PaPMO63yz3XBhbjiO4+XbHGsBHiPSlDkt8y
6Vy0XwhV3FZZ9fQ0ytH4cIGppGOEbJgi99F1HfQaqCtLZ3mdwJNwMCAQVn0Fz+Vr
/SP/8f4aEgfTVkiTVOqAqbtJJvwmncw+Pph62KLBaLjOfiouRDGt7HL3tRHsOyd1
JgjwDR/pXvIvfsdFJf4x5qGYHaITuo8WNWUHCz/VwajvBFT1r7goL6iNC4otiMYY
KFbu1FllW92Napy2aUxHj/oxNXZwtiph2GJD84gg3k6MOM0eJX+K533oLZhQeIPI
RNl5MSE7h4lFD+BcLDr/8TT4rij1R7t/oLK88NU5jpa/eaEhTtDUX+sfhxejcBFd
B8cMbf9oADG5g8mhrW2l04tfUTrZcxiYAJeIWjLjv6TtvvDgt6TPrpyA3e8XMalI
o0JYsSyKc3cjodlzmlPNBPTz2B+mZH2wfGHVLb+WVbLaDQL6mGSYwWDYX0hgCpvY
06Zi+vkvcuLQ86TrEgpcq+mLCR9vEuT9uV54eSeaWIGAiLuglYvTv7o+J0Y7diqp
LEcameIJF9si8ah6IA30HxV0zrDeLkPVR5d6svUdD4oPcCCgavqcdRjqx7Okt2iL
3OrpdPdYSBF+RuL15ZZQd6zrM5b+IfLmc1vAkADUNNXcLZVSiwCK5Xg6GN8zk3wU
JxhX2VS59OUuaTaA7tGxsPSdHNOfTJvQ/TA5GBrr/4cqHTXIqg9kTbspUuRMScgH
UJbdP4fv2kLNk78VeMx035lGXOL0FDZurIB/YgT+7uQDlm6p9cHDECoGlfaiCsM+
x8tTn3HyFsd19IVZP0vYG1qEI3YP2p8TVFMmijbe1wdjm6ySLbloFxafme5fuV7L
4WmO1Fkm4kFRSo/fGKdIgUxK1xX7Q8O7/ZvQ6JQi1woXMSn/FA09eRK8HbXEYVwS
tUF7loCtclcqr8o7QKeOKcXDkdIHzEhfFR2mguqwIXAfK21wwpKzkvBaunlhKCkn
eXEnLleDwDjNZbzrd6LkieJEVSrR38lmcV9p1Q2MLXT8acAFdUt+EpwEqrVPX+m/
wtCREFzercr6+Kjz+XbeSQy6ctz4LnKNJHJUjnccAR+WxXQykvPi9J7Fn0JzLb8C
uAVQ+PHXN4gTt56h840dxwukLTailA3/MfTgwlXFpgPwK9uyq1/UIbQo+XwGcMbP
+7XoOIFze3zSJMTD72MagnJbWPIS2IaOUr42V/7anecqtAmeH/BcES8LOufNaSDv
Nj/XHivXlQCQLlk6LQqj3TGzCwmrNBbzuaaGgPI0AQvgn51yAbIZ3FsbziEpgKho
OTt8amgIS6eLQsXQpiOIXKU285JfDP7H8rsIomPQCpJ49PLtbJ989/ozMJ6g96BM
Ys94NaORzL9sLJ5bIhimr2xtPJnUe1JFKxN0qs09B4AVwKIETjZi+SNKuktfXCmo
aCJaUMBAkv2R/JJ8AbqNyh6PzP1EshvV2kMb9316v0lojwX1L0DvpRhULyljrZrj
CvV1H7x9p4ztyCUC3zTwy9ylpLf3ZtOQjAcpZRa3JDfOYmYY2IVp5RL94k8uvcck
lJCxAiN502VvDVtl21gANUT+qSwUehgNq5TdoVO02fVzMcov8k30VjbO3FppSvHk
VMV//npb/bzJA4bS2BWuOEHLDeeKjyIpnC32PrWfD/mHx7K6PNTb2bHnEIlm2Lov
y92Srm/o5WOb2cHNiFyHQK6BKT+oq41WfyjE5SFyr/Cy5ErndNRtf/zsKwwmCC2G
TPzIbFadHlByokmY2DQ5B0OJXDRFAKdt/Zud6I0DIXlb16zFqthJqZKXEYF198in
RZaAhqH08h2yPJW6kgQtRdrXlhEvZHH8UN/P7lfX/9MZO8qI+BZWw4lShiYDpPiq
h+qXGmtMCxcXmOxvRr3t/oT1cvvgC80FffSK3VYptvxEk5rH7jDzzj+SumcqEL7K
KQYHdp38H514BtDBE9ZfD5nsFumI3ke262ykfB72S4/PozKPG/cpBD7m7s/XdIaW
iNpFLbz62WE++1xyINDPlXnda9YANLxwe3yw6xh5Ukrkm7PRxoFpL1Hzf8rnCry3
mpJ99dMU00VNpZaM3lSPqDqyVMFhuFiC1t4owXOxFJW2i5F9+HaWtMmb05YdS03k
8Tf0kNP5UCXd6RmKr8JLjenr7SYPXiAW//LedK0gHzl56RGCq4ASjielLaC3DaEk
jVVuB9kXP/ig33Tt/5h5p1f19v4lzzn2kFq5c2DmzLSRmaUP+4rnFdHudSrIQiuS
hXUNq5YywR+hX6XX+RN9ln/P/bN+3kHT+zVyfTXxEtcnZrULBNl2t51ziQQ2/O/3
0I2rnLI4bcXz+QWprR0y/i+DFoiD5ilDa7WcSCf8+zoqraaSPyHQXU/dchV7f+5Z
BY001kfrjqu5n0S9SmGVq900R3SwueH2Wlm00LVk8zL0qWv7qiuuBlOBYf+KqUEX
otATmgk4k8LMC4XhvHEG9+k0o4n6NkShQSQn9l0Rmbwh3ekcH7+H36HhnnOX3yM3
kr5yzrxUTKOwSsQ/6nJqf1v/kI86AX6he+1u/ozSUfwVxMKBUaZxLhAIoLd9kmXD
CoFs6cUjcQKo6su6nb5PNRahVgE3w0UXQw/qVXAbcQcxg0k99E3Kg56Xq+bIB9jZ
RAZ9oUQMY3cD20VIa8QdztUyS/ptIClJVpZ4yaNHrOuKC9Ax2NcWPUvIPuz9BKVI
CObbyqac262k3wCAjnSc8Y96o/zOLbrlq9IKuMnCiz0ZGHA1CMY2fXIJIT0Zpq61
8XR8Bta+CuZmU6xFKGFjVgqVGy8A+mU7AxmmwMq80qgv9tyrspeQoM8w23aq9b5y
zqIQ0ZZx2+0GbiC/CA3KD20bHO6Kd0+9iYn1ARRk2wPbvSMW/aORS2SZiq3z3qbq
mCEI71s6CONJyjS8nBgWPeWzWeMdE/nIdtHLNlS9YeOoSltGybBdS6BQPoy36+YB
XybHOxvHrHukCW/SGK5IYCWmZALZ3wFa/ERiBQp13CBd8yf5NEsRZnSaVuqmlYSb
s00wK7ll8yvzq9e4pu2jwihvj+ppbXiJCbZ4KPizxVI2jsic0zsAd7hSXSSXi61Q
LsiuXRh+Emdyp3lIvzSAwT8TfKL2ssDGGxZbuadBdyrZ/Vk5V8XRShs3ICATDNbP
onrz/3Si/4lBYtXzxxXGil2Il3St6aSSQvHLo697ynulacCru522lQnldSBJtmrI
xQI6id41OVElKjohUsOhGWW1mQ26GmXy3BRYUZacWqmh8vQN3emVu90Ivj6otosN
s4/KuHVQ2oebDYP788v/rwd6VtgUQ8UI7OxgQ1bkYAyhQZp+G8Xpaqp1D5LxlMwe
IyIZO8AbUXy7UPXkhy4cnNWpJvKaZxhfIS1NuoHm3ZMl16eroCHpVAdtd5ymI+hF
3BDeKUw2L6q+M5iHo2lB4Wi/4N4qagW13iyO4F4UROaipDQ3h95RTSimwJou1NQJ
R79Bp0FCHsmAQ7Gy+x9U0ypTq0fbks/WoP4KTv5YQmRrvLU59kG7RA6QGqY+6GQG
AzF0XciuxtQR/5+WfFZy2nUzBrtxR6sQFEdKZRIBg+pwA0mY1Sx06A9mVkr9JMLo
DtPiTB5Bij/03v3nfE/0SNDg65OsPUxe2m/376to+hT8xrD4dpYNneWc9YRQJA6p
t02DlQuB438+YDSrjKCyum5NVK8jL2r3CmJ1pVQYbyasmAqAoEbwDf2SsGFUST2b
ZzFSyDKCCInegJ3DaYuVfnif8zPqFthwhOitTMzBPz8LiDQe9g/DARVYNt1rojOg
V6F1iPGhq54R+PpquRfDcee4Uw7HgB/pGTVXlz7puKM3qTFSVJs9c8B4TpXJo7sR
RXVS9OkNlSJUGY+IdmNVJB6kEE/vms3NGZpNVTf8T/MR6a0RmdjNxqRCyV8AKzjF
ffTF86h3zBOHFDHenh0xNyW0krnGyVgaGBqtHQVG30AC3C9ouAlNuNPOhb9K7hDy
hifGGFlWM85B1bgmU9Q0zcHJZ6f8OoQIS/ECxb6FT1pLzJpk0vAyNNvPljtjsIGb
jFVFjUEbBnv6779nSkzehcgsjQnIIw7VLXz2bXBtCqxhRXLSQC2xTu4X+uSpmnoI
9k3IZaY4iPsYs1+3KLx2+xgLOHfsDAfCx3hfZB8oPTrbmehTvGxuC3tbNR7E7IxY
dVGBaEfEp7myLthJpCm/O1pQCsWbjt4N6I9qJhVleXv60qHTX7hUZFqV87n6r+tM
PuXL1PXMKVJulraf8+QVbJoonAF8YSXZsyJT/IFlzQvw5As/B9mKhfZdFcWBC7WM
WG7egXkN5OdFX+gYgEvtYQZz84KI5QSBqvlN+/d+Y2ruzQqXgS+DqQoiE+o8LMt+
IYjnoerQkF+SAORTk0YskT4mBSVnNjzakndu8s4edSnV6fX6r0F0qDQfxziKTGo5
ARB8Ya3eodK22Z1uvY77Y+AY7zL4aj+Nv98UxejSWa6MqBaBYug6VmehqN3WgT06
QnVw6gDJ7YtOQ6U9L32ig5o+ppXU8JJXzwDLOKI1kj2766hOhU5l3a/EzYcEhmwq
QyduqP880ZVJ9/l3kr35J1x4bURttQ4i4uj3znFZd8WlqvlLn7qQiorD0NTMpPq7
gCpQaJpkG3tEWuJAa7k8sqdx+7bngnIfEGpLU2TDab1Cr+o9Qa0FuL9PZcigM5pg
Nw0TIZY/KF3c5wdBNoA/Q1r5LTKWEDSY8wmEDhe0CBsW/uXRoKu9lIPwA191LRdS
Nfyt9SctB8yxIZkN4plbpGnZ0kt0jaXzhF2UZZsiI+6PjNFQuKBsGVK0C5TA3UT/
hhBhDSu9HBo+8ywW9aVUBMyM0Ayk2Wgr0E4MG38q6LHAPHarJNMBqTVvHsIDLKGp
6m8ktJa+7MM7LkIICufjARFSV5b//iOVnyMEfhh/JgON07kSZyggdtM5txDMSDF+
7EdqF7GPEH5Rq+yVoWef1r5AEIRsW6IWCXquI7P8BsvkMULjnTrpX2rcWEZohbzm
136F8ODgh04+BHGomhFv1klkYFU9hjMGHk5HMzgxKAATe68wqMzIYFu/0TBP3EBb
FIza6ToJrb5CLLi4TXraOAw2qREgN3p8fq4PjonI3fNOK5lxPu+U9sSwUSNj3U/p
pNy53BCB20iueCHoVNyn8nZ4X938/1J/z5BBQvqKPVAErhqzJyripjgd9l9MVrPL
j7lyCaFwQdRV+i6Gi63V9zCtYjZmpt0/clpWb2EI0z5eQlfORrvdpa24ouiaT0rC
LO2kjyYV/hqBY/jjKRSGpw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
m51uu9EppGfFY5gWx++7CVw3AQpOAzGnI0ncBiF0MJQSvvdcYh3Oft9Tl9qVhDkP
kiPldZ5Ix/C42CwVHMCDPwdrPZPdjwETgQ0e1h1nEa2p6BqameEAoL6oq9qttwC+
7K0SiLfF7Sr5BFxIo28H4D2rbFiERBn0WJ8fLx5tFcg+iYyMUXhiQWch2yIILIU/
0cfc4t35UqbcuMJYhBLfPlk0ZLunOqG4lIRC17g/vrbwAFpRKRxZonPSgz4Ng+fs
9qX9wUBsBjj/1kGdYS7aRPPjeW0cYrbK7JsojkNkfVblwQYTJE9fmAKux+WT8jbe
6eowZUXew1FqKzUt+Lwmog==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 23728 )
`pragma protect data_block
9mHsIxNZHU1ZkJEFgYtv8aSl8/4QokCZxIq3IB5bAAgoTfXTuHBkbHP8PeqyNyfU
5PdUn9E5w/fmJnE4An3yfgcX1fZxE/yPoleA87sg/e4oTsYW7BT67EOYnoM8jPt2
Vs/xb99fhPbbm5DDJn9dXNfoTrCIibuLXgXIgbb0G0/uXKOLX+9vqulMqUAj1ZqV
TSRrqT7xGNd+2BzOzGlH/wgRji/vVMljFa/nAazyxVqS5Y6xYKvWrzatUGdXJQyG
jJphogR7fMV4w6sl1jbfQT6UfSzLpQCfDzoqchJiF1bDcLCyUTpZOw0ui9FDuDBb
sd3JNSqCkoJ3kKK7gBlImk1oEZ4PG4WIm6oueE2gHDtkTGfYROFQAvSyslSkvSFj
kPT1xkMlLiSExRCTR2lHhX6DX4eQjlU05JxxHntakJeDCv8ZkjbIldmpzdBA1LC8
4Rf1x0ORCXQTVGv0kaKUSWrQWzDC3O057rMP3RnSnMtTWXls7jsYCw42IDvUFn90
ydnN/2CXdqUlb8bj4hAdi3Aqrtl4AXWOgBlVJvIBhrToHcScaXWsmK7qNB9iNOUV
hS5B+ZUId8QYsKX37kdfP2dfVBCdNeotJBM7gL/kzjBTC2Vt/GKBpzfsQWt3KVpQ
j5zDZlWqRZuYI3/d3w4SNfLqQsvZPN3+M211IJt8TgWfYo29hnqpQYhKjctPyLcG
3x8Tsk0wUejOA4uvdtX/A/dph3Rh1s/VqNp6TnppiJHq3fnaMzZHcdPYYcbF/rwy
lJqtJzATdzyYy+I4GlavnM7wqdLbbME0SKjd1K73BEeGhO1ry58cGyLdBB656mel
kox4fsW1Dar0vpKaduFB4HvdiRSrxlrspF0V93uu0aQKSqtxjUf651HmIa1LWJ4x
xvDqNqj7LvXItP7ZN/231Jm1q8XautG9ssjHUINGi3d0xhYzVaag42DeixQ33lW4
LztLtOMXtG37R3vHDUtYOgI/hY9TyHZb1ggavkw3shdtFO9SS5dwXHYqZb4wDdj6
u8Lnv0tLkkLg9uveP5aXDgPQCggtBd+phntpVjMVmCaOYvM6ECYeJueZ10i7a8iQ
RDERP1ldVwigp6Aj+eigdlJPZAqsia29Bv05GAc4Nc+71UcNVC+Emeex8uYM5NLL
njaU044HC/9mcH7X40ycm1f/6/BnJWV4+J7WOynQjMWJ65NnJBLa95Fk23wIQHNX
VlmQo4pXdFLpQKriweQYvc04eLwkQ+uYEHQGbkFCmYa0y4Xk/m9H+MvqPQP4M0bJ
DD6kswmMHn3XIkYbv+eL0zWMo5Kc6W1whdSSGOro1xtsaIcLLxYcLAq4fH4LmtPd
P2hYKj7WeTrb+EAAZyD21PFGsVB7zTV46q/D7f3sZfTd0OolDeiq2KeFR+v3pdHc
sW82FGi94T6ZhfVoMn5LjEya1NAdI/ikyeec3TcCKTNll6Ta6FZ3EXYfgdjfv6dN
fX402gzmrI7/DLNQxVQAuliweeRe5Cyr08lcQnfy7edc9sIEnUTRlLEnd/M/SuJ9
nAmuoiPfccZBjJ3GFMWwIy6G6GGCRuWYwE7D0N6UkL9M34LW++ll4I8PYn5MaYhJ
OMMGwqrb+kgb4WcWIS/lmJjydDq4b2km09+Q43CP+u3A2LS8K3/hI4LbxVXxX4Hh
Pwnt6YpkLsBZwoBgUY0O7LK0TSaTIkOfbNZukJ+9gRfU8YuIx3rUK1qVzB4ktmmW
CZi9H9unFWoaJICKidDdHh979+GRlS2StGw4VxgXZI5U36iwAmB8RJjMNQiqlUlg
76iQHdkcFRkld1fjBMC09VV31pgKkM0t32j13C5wW+d5dFB+6dKt5n/oQTPEbszt
fDuxtXfD1bFkOWQ1jtG77txJPfvj1/ounXrr067JhFe/FmQyDLmITtb0inFs0SmH
q6jqRWJv+R+Z3sINtms5SJoCWsQNrIUmDXFXO3xE+ce0YLFlEYYkJAw1KbSvdPnV
UM4XL810G89Ox/oE5r17SyM9SphtV9Nd6pPqaH5Mqrv1prZavWn3ICCObMgdg385
su9pYzYKw5PfJyjHKaf7BUI8C/r+KhSJ6g3wQHtTdol1ObDXLYfJpEQ+0SNVUZUh
BBGGR+A8NwBRufvH4/sYhZppB5Ya67drNb8xpTwfy6xHDgtVETquW1bL1R2LEeE7
XSljMmNWxsR+mqHQx21LGqB8Jnj4wZFXzFBLd6w5YgsrQnXX2jW/32QQxOlRMsqb
s79WFq7EGCxVZeHr/b2sAi6ONHcnzIbYFDtFK1XOymTMT3xZULABY4xkzawix5hs
W/Y+nifked7nSaYsT7SFdGasGS49+8cZkLFRwSlLQXP1kKQQVW4wwRkItSu6BHyp
xOfd7V1bnrFcm+Yq6h+ffj4qEBSdJud1njOA3pY/S10gZNlxF5AkFWw81bBHrtCn
0PvNE61JEw5nrXM6uwH2dYJmDF8sZ2ZO8lfOwl+M3j4W/SyYvVk4xzlIs/EVF5GU
FLvLM+I/DatBAYIh1ABGW4g+HCpEXsCB0gXsr442Y0gd5mJnEnwQRb014NAEgswN
Avbn0lA5cosN+JBfbqNO5sEA+JkAMj+40SXMPSxFcP0OGg5aCyt/01U2OyY6ZBRB
C3t/tDFPeLnL6j5xaCKoXrumNwjkDi0PuhAGiFdSel9/iP+UgS0zyZshP0t5a2Tp
Ey7avE1s4nvoENcuGurBvzTMCdBTw60rfZryVyYFkqaguF6wBmjunfMmtbuwjoG3
meX6afbgvoGLcUkcPeDaRzDVjL/6iTNvJzJyqzoiANLOhm7RHOLc2DZJEpVHx9X4
r3gF2bhGxo+xn+uF7K8ootzFy5uIwhJlaX0fOf6uGoEw61OAv/AwMcB5x0qVqpRa
vaPl+rSOFnk37aQA1JshZMG2YvO3jzrON6B6C0oXdgfGOS0U1FrUSVlXqoR3ycmi
zvtQdkJEEceXOMD65fzch6v7bXqQB8HaReMtrSj85UIKeEwfCU5+t3/RNIAPGnsD
2mxeIaZK4Vk+G5U0tYmI8S3m+K6ZEqAi9djqLCFwyHkK8pk9DRGoErIHj/27Y8Rj
AYfBdFLlMWAWR4Jkft9MVztefCIZ+rpKWBwOvgAJFAoxdnrRsgaSIi5/pN1SAVGr
MIJEuZiOsmhHtN2Rl1qu06Obyo4Dhg7OHOt8DB4h0QSRs2LBSayqgqQ31JHBgtYz
H8GdjxiWGiYFgCpUb+gW1kH0w6Y+9nwhw3QU1M6771euvNYCCFwzGrWTE0OtB9fi
VZdWuz9QejRDizgJxgX2kuqkGcEELglQ+SPQF331ZsxWplWjVeth5PprAICAwhru
AtStUjgS8vX84HSbTRLOtXzaVQfWo3o1Po9cK3JaOaoFzgHU2x32q2qIpcWpp54r
dpYE6AN/5UIHW7tAS9Nbr7HmGLgK1bvwFZecScuE4TgWAYa9Ie9WDBi71+1sEUjN
5c7aQKdn6/DCWdD+PomQkyvsHa7iCThiKz5zpG1/eqiJaABoYVahMBZOICAU8gC6
KmJCy+CIS/DZiNGVyIw3vfCDV1+B2bBzyp+PItGE//GqWz2TGfVpKiBNoprcfQt4
JZ08gYi8nHNXEWHuDEuJFCnoWVWMyOP18DdFwEM4ehSbQ/wA11tZAdI87DOXqhw9
g/XKlPwVwXUwPThKcKsUZW2OZreJuR1aaPXA1ghkCgCwhp78hMj4QU/XnwTmgEdY
jJZJ8oFYclrCJoyu7+BfpbNd3HilQzy/qtOBIrVcudr53NaCV8qxqIZoynPpCKms
4FIQ3v7dnta3NXCJ2swcXqDefVYXzCXgoVBjfaKclXawCVjBIaLfqFR0qMdgxMBi
Wv0TPKhcveFbpQ+vYZneT392glvzlC8D6+wUWltokygX/SvEZ6gW9f5XlwJ1quMX
K8v2u1//+jSkvQhV7k2GoJ+ehhG+dP3qZ4HwvI63HsiMq9JqbEIrZBv6K2nGNkD1
XPH/HcqTBlE32dU9trhJnhhIBHU0JEjGEUo24HOl1Xs9JQxI+Y4i6+1GNBS5fhF6
lveK+0XI8RRPWTWaNoiaqV2IOQOEvrsIgduQU/uA3PY5hxtUDPk9ZHSCZ7ylArXq
2TYvA/OhSNkYA6v4CX9SW2cfkDw62IbWUGKKxxcYdN1zOm0Q3q0OfkIvxZA1lRc1
GYIheJFwCoXf2mRirJ/35hLlMXsh/oFt40v6tV6/cLypBWprMo7lQ3HNkO6HIY4s
ziyGKVG5e8Y0VQCnKQHlrQboWs2+6rKrJOk+FEzCGArJSh9AYC/x863Q63aJwNZx
eub1sI3Q+67R4HRVy1mVvQ3c0H04Vg5HthlCzLv+8vkgQsu2dcQjaeLwqvs15y+z
hdTP4vMKAw1qMZKm/B2e3U3GWiZXfQVl6DaeH7Mc1vSdinC81CWvJxGeEOdH0Lxy
SS/+SH3A3yC5268eLJcJ6KcZM1Zy8ref90hpS5cgpY2vkFW3imsBVUk1XKFvGX3k
Fgw6v+EX4mL04tvnjb4jM6Ap6DdCwUKwe1b0YLxX9oxSLR74smvH/NVsUWCRBA9/
cIR9IZSULjrGCUwatu0jTGm23w6zyO7CqzqTk1I2TRWYVat7EByjkHfiqfCN5YGD
/gXi9vV7g9OvrLhPI2TQjw757Qk1uktbRTUxPkhOrDdsyt+WIzLrHI4N19RI0Fou
Lc43xyyWqdPlF51UiA/stUVqLfg3UErEHwX0iXyikOv7SbcxACHvd9JlOXbYEbfQ
M1B89jIFsS9zvcwM41hfw7mrygsAcG4mMrfIXzOLvmp2xo/nHI8/vgTUljfrWrdH
LacM28zrI4AVnZBthZidhoiW6UzxMufAQUZ0aL6M6ACXBjOdfgjRF/rQSOYSxd5Q
wZn362RaHQaIYG1eW6tQTxz+5iF29L7Rn6bxHVkfQf/Ecv6csQUB9y7l3mEgYn44
Pbl636UK0BCZpTJecU7KL33aHi1YyNor8kuEqsgWgdL9dYpyymS6oRLMGaQpcyfy
xMCXwa1cqNXt+cFheznfX90/Bm9P0/y3zvrYllKLys/FkITWR6VdnbWlCOar07OF
s5Y0n8QO2/7IyhxTNGWDKwmlnPVDCteMS1NKdLGz1t2MeF5zeOKeUP7jd6ZbVGP1
8dvb13iBokbb3UleFVrjx2qn2K4K0CtVfnzEPzjCa0MovUt3RW/Os6LYT1Vx85xM
ZR+FsrJKbm7qjvkNZHtYkKXznQFv2OLD3djG+eP1jFyMKu33t6auPabwaYp3n0W1
4qIIT2WlboM95XghmQVYcBB4LpSQniV1qlh+adGUpmDC6UaCWLLk1VUBnsSvFQA4
14hvWvZhg+xQXypdcvHbiUXx6rcB/Oj9b4RLzFeJLcB/oSK31xiNhPatPr8O3rlW
ZZ083xwmPX05IJjFZQ8YXUdeBEwmkaqWg7kRUz1OMcFHoi2iz8hyRQ06jyUJ6uRv
QdrVU148Nm36GpyqUIw2LmxbD2rhk74fXCfVGGUwo2ZWQux36yeBhK+nb1HaOqzs
4PzQ8OZmW10i9pJkJSuV1aGgDN75AvXaNSrkqeMx45SN3bD3tPKYSg+OkgUoNZmx
rc++1yv+lZMf3kgDRPAowB8m5Z9/hDTqnQW4QirjyeFZ8bagZSwUtJi0CQ3w17CQ
35JCdQVk9NNtilISEC5s1T7T/DJu2JcUdec/OZ7nEr5TACwyZRL9UcLuzzL4aOIj
m9k8FYZT+AdOdhns76IdgxwQ4GOL4cp25A2mBcizkGCKz8cH2FZgw16TUTWOhoYw
Vn1+OAi1bqMyErRIGF8ns5cUB4dDwR8tMFP2LiOQlJohbmeqNmuvBHYMMYPDpYac
EWYe64OYiHED8C8IplYBSyQKn0p2AITPrZyj1ngXlQKRlmPWYzJFRP0XdkRmNxEq
lOYCSR25xmLXFOfhvaIFcoY2E8tllYqhlLrGmwDKieOcEZIbIewngalUICc83zKh
YtpIrHzkH9ysY7qiZ7d6Rp9CHpBX1cT3+aN7hB1EZldioezYCHwBiHspx4ckrwxP
Y1rM+ixOLJz9gJ3LNVchSGDHJwsyyhItMhGVNWv5gVzf/eG9A1YMOqWv0B+wOTQv
YTjJU++o1kvZ1HC5ER3KAgjzmU28Wg0AjZ6Lcy21FCK4r+mBPKkDHOGz0pNtK6iU
xeoWx0oB8NwNXIzdoy3x34Xl/5cSDNY/jGzbIf3eO2cI6n9ZV9E/6PgwtUATkBBg
LWaOpY7AiPoHjJLvVtvhA0el9r9kyzVO5Wh33hFSkDTnxPbtAa8SKKD0EelH006g
Wgjnt5bbNPnXe4t1Hgtad5Ywp0xZ3Zx7DHEWcFScSEOglLLSAfGMjieXIHlbPxlh
JAKNxboiOpvLMQYU3TqdiDvhEWh1LepEUNv1pDFyQEHU/G6undoay8EPH5rfhEBO
DoU4NJvIo/NBQ9pl1xo3S3FkcNtk7JZ4TrhDCIGzvH7xjHw1JVddfwEv+LKxl5m0
BOJGUM4gJPpmWtvrSEmYCtE2lqACBURh/Gwaqb78Q3a3uuRndtKVUb+oTDwjCSkJ
pwKEYSVM0ZpeMvB3j6L9WkneCrXkE9UfivytjPQsh7mjQZ6alX7NaFGsB6MPBZU8
01f3XeUZ9YRkhFxF26CzMJYc/fgwbOw60KrF0ubURCsqzTsTi1yOzwenIq+pWFJT
Rmlu+WQSqP1LR+TzYrG+lY6t6en2dY+Smoq7Ivwk0weQYVgH17zcKPBeGF7VmT1F
BxxmFsN4DpusLSu2rtZeN/ZGy0dTIlh1Hi1Hzkt+xWKl+AGb9W5e9MWtEqFrSOaN
i8lov6i5rq17/4BNqNHeFs6d7N8xnOrKZ02yOtCqp/Ovdy4NgeIVi0pgRRfa6wih
Qhk35rQG5+1GDTmppWMzIJgyWXFsrJWGDItvNaNc80Wr5hDqC9BRyB3klmtjsXJ9
rmKS6hTrZLn12gC+hmJoNMc0u6si5BJcAZJuSjhBkYzhMJvKjRjzdyuq/J1w9AU/
Go7jaaXuPPqYZpgg2LM4Zuy5M/tYbyopzghkZegoAPrOlq8xn7AcxkI31XXttap3
vB+1epHGxG2hJJ9UqZQrTNHS3acLvJbsS4wIt9jNhspLjqBbnF0PH3G3PcYF5kaP
5hdBbhfANzFjcEojxyYJG5POXDfu6iSL8vTFdxnWLid1DxhDr8VFLhnmAfl9BXQU
woTcMMpvfDKrOytf2/3C0W9grM6T3DPQyq7+eXXxsfHhSJZzNurrWHrRMdhgdw3G
f8pB8iAe/bi/cNff3FF/PUXg4T4YtEg4M9t53oqPtp+crAJKk+TOJbXkq0x9CT61
LvaeOU09d2RW6VSt4Oa8v+QibfwLy19gbyJan0PNYbWtIuK+HSarQ06zdqxvp2fg
cQlTRAS1Y1JTAV7KZOCqApgBttSycJyD5iInOOhbh9szyBxXvRGhe3+BxWqoXfsk
nFcGSK0jyOgJfvZSu3MIAseBeiTbJNaEEGN6OxBNSXcj0Yh37G26t2iRWr3z40s/
BYbpn0Jd4bIxJIiWGejnzToE+lJY5UEx3Se50rG102CFWWgNK8NlaQJ052GdR7Kw
pnJ0r8ksIrVCJX5OhF5aDu6ira0xO+MpOMHuo0wTCNjM7C+WuoQQL4ms7YEKRhBF
Y5ZJSz3uYmEFBHhwFdaFL/xGSrx6CXJD+9BYuinIdLApwtxE6FGc3xqlG/6qarc9
ep8vPe5dQ/CWHrKIp568kFuudRUio0BBkYacTwsDB+R0DdRMHlQYIiejKErn4U3L
Vwql2i33h7RnSWqPpgyD657zAKPQOx5vwsyEuncNJW1MNvcpQXWqlfer+3GAEqTR
sk61uAXYPJX91jWx/5mUMeUQZIDXLavBXNsDi5XSIpnzGDIU/+Iy/a0lHO3r/hU/
FsdhfyGnotJZ/KBKr1TV6UImyE8PZgm6QFpZld0jxljCKrN1YO0MXIZl5IILOjpU
nhl2fgYicR1zht1veR6l6GDT1J7MceSiTIEjfosO8LbqK592MihYcpk5usOybxTt
Nq/K91jPQQ910N8rOMTpCZJcfgeVVuSdXiBiCjIL6GFF3vshz7++28e2QYolYgru
nPkx/6ednvv1yLENAJPsCjj8Lgwy0peBPiF/dQehd91wTN8MirTn9X+bmq+ZMM2k
qmy5Z2Lxn4JbkeznXgtV5CxcE+Xh1mFVAi/zePplEuwd90U9KFoDezlA/u1rpkal
5dAOnYy5vb7cY3jeD8mKkUYvK/wxCFY83w5Qq2fiJKSF6qQnsd4rU06u5j0cfdiP
K2kHTn6a/az+FFAil2y6t4bTnEL1HbpAQhXFD2NACQP/wpmMJJVlQgDDPAk6kbVp
NgAvcAo4DXGspvCQ746x+ssDkQe2g+Ux//Vdmy/jYqFFm7AK7AFK2tByxhTY5/2t
9U4YM8dOQEQ/3MQ2nkOzZUaHbJmM2NOCbddTPfdFYpE/3OyQ6gg/xXRX9n0QVjVC
tA3bDEPjrlyFkz96VLGBVOvfL9pNUX6xnBdDgoVoLvx9z1Y9EQG2Iy4xjQT6vq9+
2IZdv36LQI4GlkcJrQ27rnwZZ5/KiDI+A303hI2Z8spK8r/QwC8RTlKD2aDowxrm
lGqc013+jGsdjdTBZfl/1Gll1smVBr+tEIU4L488l8Iz8OIWQDJfbx/Kxzs36FQ8
LO1sMhyA19ydo7oe0eENkU3PjNbcT1qrnRt/mwhp8kKbMJf+jo77i11x4zCxh7+W
U+COZlpL504ryPD/Iw4tu/gattrhguBFmbqEu2zDepSDpX7kR2WeOg1isTXGWTTL
6VoV1xUS8bf1WpCIjuOpEId8oXCBgSL4HPE6X3OIxBZ/IGTP3mPXlpe2MtUC+qmp
BLF30KtnUAUwBUeSvnoU0/l9lVrew6DKfyUQxGN8m+IJGT5Ozfg4ewxajv8xFHXu
UUyf4gA2YKfty9xo3vQlXLhRxJFFln6LlE1i1g3xBXNDdeTMQx44912/15Do5ErN
lnZf1c9eOw5RlkKGDWIYsyr/Hv8gCsFUsysjqSeMBZm2Xi8aRVQrl2b7nStckcB4
nLKFtDNvT5CwYX2mkWTpcnchYWASVAmOT61s/otBgtWIAaHDksgDWLEH5glLOqo7
osAZLfdhJ/ObWoT38TfY2xxcj404dHCk0n6s393g50+ZZvPFb4Z392LO+vnZm7rr
qRni0+v/abaS6uxemLgqTpyfJZKRH2Ra3C8rkpbb6chnpvROHw4L9wJUCYKNhznB
ATBsGqYdCgBe3DT5MXyMxc0mweguuFgpjbUySbeAHaBrPYW7SFtDm4tFzsL+pMI5
RTAkpDwIhn+QdMMMMCOXM6BcgAgb/mhw0sLA3HSu4nvu520gJ359TFyaao2rJI9w
2dRRRCKOs42uN90PATKbgWQfrQJfoi+/XWfT8qqwVe0XXwtywrr5isV1LPOfneIW
hSviZr3Wm9kAJjPPEYi4ARMyOa1axwRUm71VojLlCxncAVVytGl1ptysuAm1Pl+K
0aU4dytAz9cuXykWLzJZEDbrdqXjRg9F34TqDfN05Qx+p6QWVba0CrpZAMwmtKOD
r407DqP24dDzvUvyk+04VtabkBYlOhCT2rhytwux7w5ZQzf4S3pDiCpVObScjngW
5SXBCnOPQacBfrcBcKURIVUoEc5/LraFbCsmDGO+7SOv82/ozlMGoizC5A2rIK4Z
bLH+QeJ1WMOm3pvGaaUrH77+2jdy7UP++vDhRPTqEbsha0x1dkndvmWlGPbzo6K/
cssUqPO+SdGlXoV+pc8h7VesCfKJ019u4vSslyNM/OriUzuRBSv3j93P8kRbW2IE
4jCDBSUQmQGtgf7t7jdaub3263QauM11BaKwBLebvuOzqH8jw4eeexAWqaxu9Lxo
M+CD5/D2GQDLGStuuj3KCmuVUAz2mT0jy6HTbqAiSNBC+rsCD6CXwejMn3BudI6M
6lQEnBNH2wZU99R19LWxlHDB3MDaQRsSVZIK77J1LqG54EhFzhbw7BlZt09G3Hyt
NNWeebvJzp0GzI6J/Bm4oMCQt3q6mB6KSRukAQzo3cJ0xFg+JV2IEuuTgPuNIu3Q
Igr99fFpMedL0EC61DkkjqAOgZEPvVS8adJS1dWrtsSovH648ORm8nPQ08lzEMdV
u9lEPlgSP4e7PmlrxC4m7WMlVbeMmWAl2UpS7QWEoUN8+pj5/lyPHXYARtG4FsB2
tfnEM3AQTpmkueHzggTe+IYxhQiS3Wh2/0ArnSXxM9g9yNDcvsLiHikaBD19W2dY
1L4vhBhmVdIajHS646dANc8fKbmXLHfdz2kwBK7VoGCyHM54/mj7Foq5QOhE9D2s
FsO4ee+o7SA3u5tqDEj/qfrx0nRV8VuBNIl9GLbQ3ngKcIacK3qPfgRHodqox7DD
IMXfGvXfIkAW7/+rD4EWTVa7VhOkoN3HV+3KOBw0Wirh3CqZTIsQ0C3kYtjSFGqv
7UGujkBxyTwqWEe8sK0HWOrL8+vYxN6A7HHXPxCPDHQZes0y+ichdG2b9MY+shzk
W4a8NivNqccpg7BkhddH7MYdtbzO9M6yMrKaB4FZg9TH8egL92OuQmb4AxISPB9C
YdyjuySQYdzlzbneS2/kod9xAoYubRDhAC76q5b+M0Ui4ctEu7Ppcdx84RL09Mk+
sgIIQfiqgnRV10Ok4+qUxjOu9zW3R3SnJe/wmAe33K97DXNosv1Voq+qGoIMq7JK
9hyt5/vlY/K6C6Dj2SbbWo7z/20gkND55nk0OXbmoZVp44QFHSebF9iyAQLnOUL4
b6FktICkQGLZSH83cixNf55JUUp9qeBYOfEPaQbZSRdRUrvsaUJPLpYBkIhd04Fk
W+Vu+7GD5Ev81dwLGCbYHkpkhk3r4gozDzwfVwUT6mLngfbUzaq6VuFUGlxNMZ6j
k/y7381/mOopp1THEXj8fTkCAtrfjJYTVcMwahKB2DrGIZcr0y6T8luiE8vkj71G
FUd5vE0UwOXJbqyWwBW40CVo9gZ56Ndu6T61vgG/yiDFo3V+oiYqi/rdOvW+52Cn
KCCGk2Can2VB8Cqq+pcDJ2SCN8u9WE4imORAaeyoejXdNRd41azvvRqjLtYhLOTG
UKvE/ZLAck5mcX29qY4WEVGheFl4wCWIxpVFIplC5hrDjN6WIJE9PEgPURKYacEL
2z9av9fhkFXxVxZufGVVLYGVopgHOAKNayPPOp0wEOPjo1OtT0BrXZyYz2APf2RF
y4X8gjFySN1UdkY6pbboFQvmadDX/n7pNPZHnfE4XbOeL9sGC0nc0Tem2viQAX33
BLKVV9zkbPSYgQuWP2rE8uwlR3GFMcdxDynxE/mwFmEBz14aWP36kwEUTqrpN9LO
OpHuQvwM0Jo3fk+WgWGQ1mbxxdBaXV7RAbA7uYOoe6UZ/7jhp062d2C40wGAkiSh
Z9QVLEuX0YoPxRpmKa0f0aV9ExZfPW1Cx76WeUO6v8RPlwe1a9I0afAeKgQVHAbK
0iVNthhF2DeBOu3fwZiwCX2rTph7yjmx9YpCRHUCJW7toJatUoOfiB28Z5FWa/wi
ygXYVG/GNLvGxaiWah23G8PHlWxTeqIKYL4K6Y6re85Sn7/OQ88ugwudiPN0Ose+
p2gvtJOUkPJEiBn1378OeY+FDVWssIIZUxkLZbxXs9z4Zn/Nn5dqg05Q0SCTRYam
11QNNiF2eYOSqsWWQDNhc9m8E/L2j43uy8Y+Fsv2qEjkeCrF49vD1bj7kTI5juSO
MTFRdZcolzLY73EBlonhmvX0EAqtHQn6qck+iJyXOobKSxTNN/4iViRMta1TeWWa
egPLbUH00TVhxp11kJVh1hAQGPWC6ACwjJZwCEd3KIjdLwIaVsmP79z9fbQzZqy2
+5tcTbNaJ7XVUUnni03ZivIE7MPpurHdXCo2tHiBpyjBpGU/HsdkfIg8LBfiY8sQ
wFOu5zUJ+Ceztn/mzrfiQzIzHFmdbSUSr4Vqe26kAWnslrP62pKyUaFZEG26pmKK
85MUlJzPaz5bb+i7Yf2xEfl5mC4x7h1kZeDorUzWru5vj0eMAuN19F1Y6JURRO4F
U/aJyYDGrgcoBYzj3ppebaPklfr8xrfJwiyJBtKicMa4qiRv1XQIJ+ZFCctVT8mE
MzHdi4Z5A8woGufblIh0k6IHt/UQsWX2CiHHkevUTUEbzYR5LGiboIfsalGO0oe5
Lxy7X72u8CJ5MVs7jMzmj8uaLEtWa4jNlj3qJq11/yNDxhW9jVJ4XG2rruODII21
YedD0uTO9/6g6Nq+Zr+RugVBaGLT6bZ3WpB+EM0e6CcbdH8/trxu+9BM5ZVSBHhp
40CHEvJpoFpwwHhxzjrLjbOZAbTN6QC9oGGYgv/wxpD8ybGi2IO6SjM/X1CRwF7Y
ENQLsVwnK+tVClMxKli0vh310lROBq4VdESMLH8UCh4qX30ZZJV9mu12UGFzArzv
h7oJkQQ6sc/NqMGPM/UibMt9HpJErjnqsKobhjoM5otMxM5eEQ9VpGl3Lj+YCG9j
HPeWRRuIkfG4sUnHNxJnKpNJZqGtXMWiyeZqCZdrcTE5MNtCkEf236Tyn1iyV9b6
+3L2PwAeXMV1vuUdrZVgeTq3Ejeo8G0Z7Uzof+JB8Dh476O8lJpkpwmCfNk7/V7L
ofOLUr4TxmjW7Bl5RJq0W14ag9iT2/6pD/xNomg5uwxsIRhUvd5ilHykMyiqDjVl
xzBB/8EcZQ3+SXlHfICMmYO8Zr5/8+6VmrgBpkLVr9mbsnK+3dLP1tBTnVLrB3+2
o9rCGmZa4HbwLX4NQUHqvCTsjJch+AONd+YozQGOXYggVd2kmEeYqsU2WuFx5g8x
rZqa4I9vzOTNhT1XNr1WFlw0f+qxBosQ+Y+BgMYn7cu1EQRhQQn/PrULY2XZgT5L
0YBMOImcHULFJV4v2mxkhp7z2wbsWHAaFnqwMKWWtxDR9oMzddd5ziIWID77TP04
nV7Z9oi9Jo7ZcHhnSrMU6iY+K1yEx0BST8oCXPSXe5cTjzUEbdhe6fXZQwf2hu1K
TA6FH0rfSQxXVSujeN7G7Wmbu/dQbJ1Obv2TZ46jz4JWI78oENFlx3gPXcQDUy9b
DpIh8yBeC33JsCkeoam7I4on3RpSREBUy35rpefFjEu5Jskm03Mcj7JxA4OLg2rq
nraeEU1Pxv722jwTh7m0NmT5HIEuKkz1eOflZsXkFHFzEe5Ji/9nXFjfkB/MC2cM
VKLJFOh4KQpytSBYoEj+jNW4+4Yrae9B/USnko/2vCQ+G3U16SmVmmg+m+djZgS+
4h83+tNKBLbd/03qeP0LZi6qRTAfaw8OT85qq40/d7T9syaB4GXG0VVC3l+DCpXX
8xJ40ECDGbpbQmzQWeb0xChfnlSburiomuU4y/MVBvqr1qLO9lB9R9d0nelgf9NS
wqb6UWDtHtKO7o7b9wtU4+ONs6LStafgEUPYX2KzSaEgz+kAdzNXDSCso7QkNr2+
H2cHkN6qCb09ZqxffhUW514ciWa90o390ZIG5K4eEaToYLXNQVuoIlZ1L9+jvbig
oEAjm9i3ZvTeOm2KQoazbug/SkPaMvm9JAZruCdUgh2KNBGxOsEDjQ0LG9mq4szJ
/TrY/ML9w4kqxbrWzbDMhkUD8SmtCHkLOSVd7XIYu+7OUGhbevHDtxjz+8q94g51
oLf19yeFWE4qr2m1a28/gBxZ8sI6pNzUXIUUiM+hZjw1NFxayBmTGlUeBchM1zan
zMVf28gaauro/cAA9eTWi+VBLuB0FzUNGSqzXVCDTZwGopUPBo+7CPFzgDLLpg6G
GUN4XGfnXJpettqUUbHJ7GkXcQnojOO6S1vssMw651hAOZPrNvZ/jmE+QEo8FkAn
EJcFG/eJybAvm2IfH7kD1JGib1J182g4+Yr0gQPpOAJq0/XQ2RJnNWKDk+3XlIzZ
ELv3LvyTxceKJPKzal6orER82XgJknkiMx4vHwpM6YncOW74snaXz8BsNDfuAduq
eMFTfptU3jzuvA8ZAdcGF4+pyeMSQz0V5q8ozSfpadv/2sBwTTQlt4H+v5/Llq+m
4NDdOqgzTT+L4Pl7KuTWFmmOLwXN7IRTNQnRVTbE+Q46/A2M/Jpi/2INX6bW4JEC
4/VRVW7kFRaYNU/hDhDw13kVnaW/ZZvxzH0tnAXqrynrFRCyK9l8Go5ShoK3GK8o
JehZ+W41+vFRaP2hoQ239YYYWFqEFA9jEGrc/bZQQO2u3lFNkE6P6/TscBM9DMuf
eLZyPtBULWgVrFqcuDmWPhcqrqWCaILz+ZteFucD/h0IsyjwqdZOzU/A8K6QWJ4f
Sb99tU5HJKox0ycjHcVQfkg/ja1nKJIhBiHACCfzEMx5cTCrZ/sp/vRpujaRs6mQ
hpeUwLM8HDSbM0BTxhyvDidkfX1fXNvIYkxEvd327LhEmp2/MqMGAyA9ZuTu8v/v
8lA45M0yRvjo/sGgLpVC75vXON+tmvIAVq+7zvK3EYMnHsEKftsO8zezDuQKRYmF
zblKnuo07w9hAmIx+Nkf/fJHrvvz/a4mi/1dS8+2Za4riqnK0yzJqzZt8GtpNg9l
A6goqWU91Z9davfw/UZvzPedQg3mPzY+qJ+lF4R+ZET6op8oVQxVjtMLvimjaTSA
DiHZxDekXgy+prZ2SFXXv+QpDtlONMCSxB4L0Pf7R9JxV2hcSLkY0jvYlsj70uUt
kVALW65Nvl0WYbNdygUSxZp9vtjAtUCbrAyZdAsUAOm6r4ib5Pevi9M7Hi5XGYyI
kWF5aJsl5mms17oeKT/WLY8hvAZ4c4+996T8Fyxa3h+4TRsax5+e+S8AU+C4fUBY
Y0Cprf4vYJOzD6uhpScLP51OVpFcY6I8rmp9b/tM+CHpYwJLMakE1eb8ZNXYv/lx
HXBnzZWthslRvQ4t8c2eLdpGaCqdEUSQrgM1r1aqIb7i95giOpA3BFicGpDFpZZg
3uxwrr/swWFxnqaPDwACybHTrS69hK2//4TjUeT0C39B+nnOpOxN4keBzJEuMh50
LUpEAcAIJiyfENlwUD4QkUonqhyz1RH1lOIS5KT2dSWVlLP07EYMTUj3lAMHvokt
KG1LboqOe8FP3e8S3/LERrKWIyo0Qv0p3w8ni3/7y/k7bp5zg4eMzSUI5vZr/koK
8PP8psHbmr/y2bwRd2q5ktNhS+bBIqoNubJBJnK8RYr4a8a7UqhbNw8vx2etl243
iPTIQ2sFXJFOCR8HcM9BkgpOgOsyClSLwvpzCas/cqKVan+LQWBs398i1Rigu8Kt
GMFHl4R7kQ9Mlv0b16iIKs7oOKlv77ojJcwGfK2wzy384lQiPVvpZBRg56LCaQC2
bSihlLDI5qTpB2cktxxoN7rYHTC9Zcb5u5xPQ4z4CYk1HgItkOZhRh6wb9x+QJKK
7gHU1O18Z9PNeFimDCG0iHu4GnVOnx02RcuUUC7AjWf2y6R8E17SMjglqK7pQ6Fh
u9nPqjS9T+pCpdSQB6b7V/M5vlHu2RYrRpRiHVjR4ITiJpPymflGSuD5iCUqhsu9
AoUAwG252vtyYwsexgPj3GHWfkmoMWhpcd9O9bOK+qQPHewAXxMQVpmeA23gjUEp
4EscugWc54Ny6wBi6JfGDlRFWa5ilCmlYJpEwOGUSU093166ap+sWOj+tCagtSre
IVKVwIAzR2YaJqflci0wSgGo5vdt0++QHAejTj9JHnSrLPuweFFETfcsGVlsCvhR
JdFnPqCIuvvh9NssbKuKyQ431DmCOmrrRuofIioZNfqHu0zeKRCQ2R4k2vVWdaTl
8KjILjlI1pqc/mt8g4Y5+oNb/ARshgtbiTBdxC4JARcWx62pETYBRxqSBgupEAy0
o2+VPpfP436WbkxLmd7zWbUVw3Qfxw/p6cUi7UkPqEzs6N6RrJ7gu8x4e4vO4e5i
iynXiPAgcDNc+/4jICfysZQUNsBwNk+kFydoXMXwue8EttBZfnn0G/2rk/90Od6u
VwO1urikQGHjv+njc5z4EJ++h4MAkicY9zAdWrzDB7QTS6EWWqVKBASvbz3Q2Uwj
Yi0w4tj83UepExlDmtXvlLZPUkBpKb9spCLckSuOVDybVUobvfOMOErVXTXV0wnM
aTQGeB0A6cRir9dkkCm95xDCjWsRYpnnvw0mqc4NV5tcERAsxl3WM6Bm+49Sjpyq
2OPOh1Opqd4gXvxSyPpdRTjuXgambIdDn6QV8W9xo+KOIQTG8+L9IdvNiePBxDko
g39P0VZ73xDACNbKPkjH4VvzKCtj4JUvDgic8sCb0J842M2qu3Nfvbyb4dNDyycr
1eEniSz4zlizlWn2Qv6i8brkAqwsm/FY3/uX6tpY49SUA9z/XiztYVF+Y0Ymxhn9
NVSjlQ7IOVkH6xVYGewksxC2R+VtTrk6poKFrqkWgDTT5ca9bEr2pkAbuCt5Kvcg
+C/0nzt94aUmJeq1rCvLfhhG/J3Io9ox4kfrx1RvmzROJoKa5fGqlW0HNy4k/BGS
I4O8g0qtU1RmzHqj9hghYJ2aVuR7CoTjAKoj9lVs6/kb/P7LZRaXnkle8BTNMq4L
s0QmGqBcBIQ8lE3RXAuBkC2N8RIW2GnSmuWF3L9eK7T2LM2qLYIj/tL18BFr9T67
EK75AAG1TNzLbTd5GC44W0ImXiv85jAoxuPeOXwNBR/Yce8rmOY5mz/h8kKNbk/S
dSCZgV5yMg25Fa2M2JMq/KeDuEfUQCzzeaHDavPj6gqCD9QoZUIQ/S6CQHcQCxVv
+dlOAQH01peoDCrfpWfcxjnJKpZW+slHQMscCsbLIjjuGOfFee/1iGy0k394GXt6
tvKmZT6dgeRyCn1Igb5tw+p8COYnWVkgoVXaSR+ZIGhfXSKqi+hofNepUg5Lyr1f
+g79R5jJBqE6qS3veOBdbWxzbJn+5S0ZG3YVVpw5br+Fk1r4aj7tJaGCQCSoOrA5
Fbk3yXXcvX2/QaPj3+4/FXIzckn1U/LKhOAWk3jnpnHvI5y6wOeSv/LdY9h/tStA
LdTVzPBNbZO23+ZWOelHc+Jq+FcMY4pyo5io34FWhSTs99Gu1T5F0ptBX0d9Nqh7
XDaMslTa16Cx5K6+rXY8sKtmJ/UHZOjxNNSc9+N/WOqH19GgLKBYMv555wx6AJYq
h6W6h9+SR070ajknfUlAnhZGlYhmMm6ZoM9Vs7Usrpg+zcJuHHasgrBhONGavioY
8nNz6qHyd+Xypd1GBF6v9Gmoao4c2RSIw7GmpbGAN0dUNH7Ij1e+H/rt85bbklPU
FKDJWpCyyu9eIayA411tNIbdpCfWGh3VWfbIi4/PkPb+1CsVL7ELgFUJ/qplMhmd
1GLMwFd6n78mK5qtoY4p7HPrnrcBDCmNPLw80IEJgl+8BCgNztOg1JH1dBjr7IQ0
acjEoY4JX4kAnTkDThAqNJW6PgcsdY/zlZ58EjU7S6k77XYu4kev5ywOwkApHoT4
z79GaPt9aFJbidtHlOrsVLRUI4n7lADZ/i9u0w0Ckq4fFFh9fnschkYmrXwlvCgE
mTyRHV5PNJLG/Gfr8tVaM4ojvWMX7y7Os1C/68YWAG9mPB/riibzg9IQszCtBHZr
NwVNn0Dmv7VJml7w5jlQdRuElHErhBTTV4YygvJOCcsSlH0KxmCTXvYHSj4dEQoa
INfXCK2bjFiSpr1sgeqrQF4sEzqjIxTl4Jk/rUr6DIKHrt+SsFJqKn4WgHroQL4Y
G/nytubJ+X04y6Srb1oTaB46CGJD8cWXdQxSIWspWZN+wX6TlhG151lOhvoWSlFg
2KuLluek67voEyL9JL1OAmq5DxljKoC1LjRC0h+50bIWKmVr9aoVcSLeWIMuMZeL
X44AzmSDO0SaUldzDmpIyxo+4/OLtNPk5bbFbQ4nJnUvIzH3oTGMjYgG7Q5+NTeD
OmONnClURmPTbS8EB5hjwzEHoC9dSM1G3n0wAw0LwxlAKxiXSJY3RWDQP1OnF339
mSuWQ45Lee15OSP1GYZsQCYU2wvP4U0ojqQQLErCJ7mzKnM3WObdZt/SL6FHoEse
yXskFcyMXa3L9Dubs3U3uKp/dHBGeitiOr2g8PsrDe7TQZRbA4V+79cEZy342MJJ
UOvqp6TvlJZsEiqy6fuPjOGgjGoeArh9h7TDmEuzDdiJE2C1fOtY7iSch4D1oaEx
It5E1ny0uvlzj85g0OvyxRjHpdvRr/f2+5S8+AlHZStqP5uswUdcFMgFsUCPCP+Y
ic62YMsWps9Ec9jjvl9bmsGxR06eFBM9Gutw3pnEEON6nWNCkXT967f5uEJfnPwt
9QxH5/r3yxkyx0F0gQ1SoQuQQhjRNeBfVMgq4FoLJw57/9MJW25U9PnO4I88u8ud
TfnDXXw1YRrherMeE6koTqr/ep2j4Us2s+NM+UeeoWn+qpfkGD5c0/SQJKbXuPtZ
UdhPv47/2PcF62C/8vufpC15yqAh+aGR6B5mFRbDLf6wlIBcmfoHT0KXf+8IItKZ
xv35gr5yWwMw8OfAfcpMwBSJOyZnptKm7IZdx3bGqkBu9QejZpu3++jeSE1jmQLc
cVOvTvdBH0Nla2nwoc1J1LQcbJ9vvqR/z1xovKhSlTBc8ULi0Um7qqBEFbEPYSfq
hYyufBLuKkkHeqhqtJjiDgVI8os2NAa2UTNTNmByv5naVpXYSq+gpwacik3FbB+1
ow7tlz69Ay9FEXPZ6bdBvip6001mZhzjgU/kK+/YWK0reof1xcOPfZXWl555zeda
2rURcWmQwu6BlyRDM71VU64x9yTq82H2943ekHm8Mgbzh7IHfdW2SHbuNKfYb5+C
Y7rmqM9cU22WHWtm24AvODKP9BahNY1XxZ13zAUaEMbYjF6E+Q/2RfpmDwK6ccTZ
5YCs5WgypH9PL7KYiJmI+tWSh3/Wt7tkrKGZ1gcOoouZnqCkqzcFPi2ZtHkirni1
AyyaAGOzPovAdLUjwcWPDCpknNRlAD4fggvJMKTAfRxl0kyU8WmfOKmN8eQA7nZ0
TKeajctWd9vaglji/Px64uMkAYDmanC/siZxXGvjtu1UYX3revP3TCORj/YB1NFC
b+X9Z2haNy4ua0UlFEJYpjykn/vJn3zBQu4pBCYUymKuZgWBWMqbr/VP/uRlx5zp
oElUFA00TWqxOSXHuCxyLRAPDSFM1h+l//vmbI3ww+MLWdEnRWhhCljOx793FPU2
9XPCxyXY5hNrK+YtfpGOD2ifCxBQWA0jSm5JE4vc0XIEzayAxJxSTWWw0t4Ricuu
ag+9RH2Z60FTLxy71sF5m5IRpFS0PqyhI9VyvGJZu74VPmQ8QWYNocFLdp1vIwmx
Rgk7YQCQCb9Q4itmfRxjeW/4Jc6LHtDKrJeIgsaQDXwfP1tYZJ2YQ/oNyqDQd9wf
IOEE/Mfj9iWpYpaWT95KlD7uCxptP7YXKiO6qgES/Goufc+JrRPZqV0qxLnYSqpL
x+ghniTBredz3nHlzlrJuedRs3GI2v9pnobGEhakIRgEgEtCvR5hSjb8DBqWDSbf
yU1QNJOyCP2xOwxBZVOQWpd7U3bWM+/TqJu6nvPL6UwiSr+CvZ53kgfNUoskKxKI
Qqq0yWwDppoZKbECvo8n7qOFDpFzmu1SJ1T59lOzWOtIjWlshtTvvwy++hxN1FO3
8XWOoFp86CcFYiRu4aAEivRzxqs6VIl570dzl8BTWE01WVFd6zgpnFFwrZzT+Etk
TdbgosOJ7vPD8RP0scY8iy7R0fAtE0q7B1owShDJn5EbU/Hp37dPYz4h0H4cd9r6
mxlq6iIOFOiP4riWIgLCf0djXMpERpXir4mPAY2poJhEAdD8nWL20EqAFZWtgqM1
0w6NsChJKqOmNvdwbbLhyo07txoDCEBpgXYyklULHKVLStGctfIqMRNyz+eTjhvz
62wtYUyI37lSiOrorGLxfZCiRQ0n11/cRXB82lNS1TeKteR+GcGZZfp2Ztaxr9Eh
3YtOvCTVk9ZslZknJoobWtjgbIPmXcWYYvedI7jbSqqwA7dqMjPd0Va8hJuGdxeA
YQlXcpXwzzQGIDYIwvgYOWeb+LHM3AhzJkmEBhMTz8ahFn9iqrDOYDRwfJE28JyC
DMikkM6XmGlBJrpR53Dm65NMrFFRSTqgNMJJAoD5tDVm7R/a7HGXbogyk52kkwc7
ARtHlQu73s8zsEUjIRURFF/6V/A2I1nWghArZqXXV+hOIMGi4UHVi9uAt8/CZHdz
A9aCbTijz1tbntMKZ6OoR4YYu7KXesQJdHeDv3vx8119VrS6wkLLISU1lObMrvtS
1iELZjQj1Yiy8jLX/l1OS8ii7dpSdCj44zzAr1C+yXJwlUPktRtW3GQW8cgpNkLI
5KbiIcRT5lKrN/1cKvRdv83P7bsB2gSYYVug6+EzQTf0d6TXQtQO+yTvn0sIwolP
wALcOCIFYnlQ/jNMtxJXHPRq33Nyn/KH8DKpTI9a6oUYFmtWL7F27lo0pJxOUNgt
sg5fh8tnYawU3gD3R6CWFa+0GiFDEEXhD7LKFF9fUSZd8PeuHuJoMypm74guD+W2
HFPjgbf3oQVaAicw8ewFfo0qDKFJ34qv9gMvTIljtQRZk8ojOQB3+wdSmrjLOnDY
wQohDvwhircVsFoHRo7qk3WlZBN/a68+Uh3UAv9d8dtEpHWkj93LY5G37R5ILbfr
NIX4an4nWtKyiamE6wPXCLOOh45lgO9AmlOV+yjmdu5Mw/UnE2hfj9JDBhVYSubH
qBeGHMWQIAOgCmB6LqhFPzz1jLyNUjC4tqUFpUut46PrtL/gCFfa4+ZJOIRXO14V
ysXc/0gOhOoli10+wjB9HSNPkb9laG/apCesldgfpo8Cf8dMblCEj6EybVLMe/aC
8zlw1vd/PjlLfpgqXhj0k14B6crdy4DT6sTC/pJmCwxhdLQbPwzJlsFtXeg+T3Sz
LSLpP9u6+a9MeUZ0FQUNp639jsh0cFr1iYolZZ7pJmmRTXTp2BjAMZdR5oOf5Fks
QtrQU6Qce6cB/Eu8ZR7zXUO9frSPySj7roGM1KrkPhqNtxxF/II5g1OlO0yfrJcO
HfKGfno6CQe6M1+PzAqyWrKa1MlAKc2yi+oyBpuI+ub929/F6T55zaXGvtwKNrDL
lN+1UGDykWjySVpgFVB0ubVBT5Wawav5I9AjUc/1wiZl3ntqJo9d6rvMG9OmS/cb
UT1ZaAai8vGmp2+Xi5UkeJYWtpAoUvimgPxZXav6uSZsxEln1E/bMN4f/M1sngOV
DhIf+9gYtcXV2j8Uz05erOthyCaYmoSXdfL5fZ5Obc1a++hA8v6G34cUoJCMWv4O
6FVLSFwf6bIIAO/uClI4zW3DJuULp3eqv5bBPsJnNL+o26w/emZZGGqSu2gbJcEt
l12IsLh/Q5HvzsdVqMBxp1NdIstB4DX79ERzWxYxyLjQPOwVwJLvBmuwxgBhqFS2
LWQTzKCPWbg0Iqp6Ser8QVPtC2ApxmXD5LHh0DWqe0EZH/QBNusrIE0I5dzduvZ5
csdnQE57LCkT2kv2H5p6h6jMzMKBrcgTaT76UFnpckIQtEM/+3v5UuYJ4ZR0JSTr
21QyN28UsAJcPc6noENbcSXnU/wTIH5fjfHCbbMqPT1uUJA1idfyjz9WQds/19As
9iiJjiywjwg8s1MV8vM/MrxZC418tkx0izPvUBaQmdJie1uC2kdR9kBAMSZv8fGy
g5kWcjuaPauQDXSVsn25XbDatTcpSSSlLgXcgmLyTqcX9QzXPgnA/V07iqhRri7o
gvq41jILjmafp0CA2mxZw4iGn2Px/rACwNNZx6jSHPevdjtEOscoUvODK7l5BPtK
zwP2KBwksr7WJhB7w2cpnRPVBfcgwPvQhixZA8Sgyq3jmiS53AchEAhdxpGB1oU3
g8q4Kefy2zc+B4OZ3dqFnnWq829hOzhIvlJQvSs+ojT6nYIx+IKZ3CKJhqi9jAtB
if/o75Igi8ddBgfi6IR31rmgsC2RJSAvP2ZRRbM3s6BQOW/i9mLvtFZR5TrRldiG
rSPSFjyqdnFD8sfk+Tl4PR64lXd3ePKg+2iO2ANidrRbMRTiuy0qpNHsbYpOCz29
eaHB4LdOqruiovraxh23E2WQ6HI676PxBl3BxWzMUoNgqhShijbniHT09ybOT8nN
gKqrdukan1gQf3lt5BU9YZdDx0IxOTlotmFxlyr6dW8FFnbt3qECOdBIcbSipFQx
QkKpzDBrncdPJfz9+g7s9B2mPEQ6gbuzQ8s4wdLDchoDUsg/+UKYhdHlEiL2DFXX
MAns72XTGx+F+Z8TW2q4gia7k+Eu1VXEIHxwImIIAX9lU1Yx8omfk1sBlxoTCRy1
kmFa2iwUGnrHr/yBOXBdNtc8d0B1CGaXaCI/7UC1T7QoPQ3lBfvvWzKRvDm5X1jH
vGwPa4udq4vm7kCwbuCFYTm4eZglTnU2UkIZFnlUv1BPvOz8GYwS/URuuullqRUl
wVnrFRJzncbUypKwDKRnOEIGRxdFp19syworNaF4WrRklMHcCsdqCw6DU21Vw+6I
bj7h/4yKZVz0tRqaXUEBgUjZbQ05dpm6tF0KCIUhW0rgHyIt4R69qt66U/kojqtZ
plKKVsnm4sM5Jqf6YPo2bRy1YbVLyktxeAwmSep++IQyFR/zgZud6jF6Qs25ydku
YjULVs1f086jKznpTAalA8PfcJCxCSvUOX8MInB8RcwUogrFVh1FAvA/7AclxRQ/
VSfXbEjWCDiFTxSgHlB88BLj1aZ0rcXsous3dUsBae0Q9EO/T+rMts7Mi0R1SxZv
IA72G3bhoqShMf3lrvJGwyMpNfr19Wd++r1eCmf3tpNesjBAZukIvk6yA3sz/2Uj
tLukU9vMBG9qrI6W1EIkTi9XU3HyY32dSz4iFkOe91jwxpSE4iJGQ54eiTRmOvnZ
s+Shes8pCa5e43ZkTUWPeohFIw5pm/Fk6YWTlCbtednzZSiSu5jahkuDsNlOIQx0
L2nn/ZQSJZXdRJrcBviT6xlNRmVTLyP6FBKK3aser5GdpL3o3sGvniBp/rGcCuZk
s+pdgr+T+ixd27mEvCZPM7BQvs71pCHXcE4C4fXeFXwrhUKsD/jwoqaobJBSGRhh
+Wmz7UNRfjA0++TPfzCO5tYVln1CEESxGFfz2AGP8GzLy5pWfC45QyERNHIQLNuc
JXrToOB8coNn32mbFZPeBpsXX38IbU3XbJbvMYZqrH+GGQYsCKfXETpZJ7V1ZZu/
eMFUZ4xZzUdNowv/r4XEAyw2SYOZr4JkuY1E5jodOzavnrV/oG8dKTlcjpsHvc0z
6jbyPxuwWGJUYKBNKzupwFO9LSJD9xIfMpmCYbQVj0tf5/pDptlaKQlxO6blXoXz
mtT44Z6shc1atAZTEdS1cf4aPEvublQnFZ/m2VyY+oIlFuyd3zh1aknRhrPGjGEl
n5NhFyPiNXJsQH9CUgvboXmbUT9FFfC0DmTb1WduyV7PKGzEDFoQUh8H4w6mEs6g
+x+YmisE3p1yM3piBTEc5hb+F6pTx/DodlZP8p/8pKxRWArUTAe4VSqVBEcqzc0G
lUPw0j42F977EqdbYLwt4gxjoK4md+l6IDfstWxFTSub4z/CH96517qpRCMK0rcQ
LGKQjZKUCJbfOyv6FjBQCl0HkvU6VQUlLVXMXhihOMAgAVgmY37Vfo080qAGLGlO
hVlZNZc1/DMaZHQkUjVSxf5fudOinPb5MNwHLEHe0B3J/z+qNGLG8v7rRWHfZD4g
vgrMH9F5k1g4a9oHc0/rsq6kwFEM4Ixk79uR5LN/jNb2RIOu4Opesw43SIFK8N2c
xyp/t35hxLWAkcJhq/a2DGoLOuoGlx067LWyXzCa8u0t/m1a7k8QFNDRo10EIqPz
EsdSLEZ9N2bHHO+wZx0S+FVitd7heNXAABcqMDwohO+5XULEmACv9jjvRvEvP5g2
FmaeYQV8S64LtP/TFFVHzrUYIC0oQpk8emUsc2vwuUAEmNIdb20aCDQchCsza5jL
gAWx07BW27BcaWwQinJU3Rd3XG+8LNKPJaigA+WzrZH4driscuHb86ptiOkHHA3m
qQ1Y0P7MS7GdSgGXKmoBS++cg6mNVpz68m9+EFFnAdHucBwtwlSkiYyyolsnxAk/
62yD1wKrQ7v95ttF6ZSkGqkJUmZKQ/nyFo6AjtjDovVuxPSvGTz/vooBvBCOUQfd
TRNXd8PczmHeLGsCsXrt63tLERn+Qaw08m9BzA+9L8wIVVSNyfQMX1vD/ke4kfwT
wT3hEZ/OJVK1GffIuFlfwd5hYOJvYd3jfymufhAieFP4nw4aB3X2uzanPwdSYrHS
TzVviEFzbmf8gPABZY3BIvKbmuQDIq2fovYEAZXzF9dIEupZCsotWzL4Cy4l59zU
CT/7nonpGIqpSn+oRf88t8JOrnoGFko8HcelaOvy3F97+VH86nD+Ngb1Vf+Y+kP/
qbeM+PvVWeVnrbh+dvfPVjO7QaDq8lOH5JOk/6ll0IJMbgynrqjsrEMhWazGI4Xd
XeHLal3iZteJjTGzIqvIKkQO/+4fzsZ78dAfMOrvviC/P7U7QGKLF9cRxkPn4YT9
GO6Mr6/rLVOEqLGo/6W9TonQSNRK3d2+xs3N1w6J2GQRSAcng+DbTEnllYH1VT8P
APlaRX4sB928+TUAPw78OxVnsarEgvgrCUHXljxtKfZRRNCOVCTUJpBFrAF9opnT
M2hdptscM4G/1cdzk6pMEt4vw9qvl3Twb9F/L3Nr7dKjNBthBJl4RTTj7q3GaoNy
NqiiEKlhqhSSKAdTU3ooFk1b23kaHv+hxUyRIJ356RyZga68z2sX0LlgNDSEA6dI
4793SOc9O5yvSUZYChDw6SDOU1Np1dnyYbfU8lqU8zGOQsd7CUuIfwalD+8VPZO+
xxu/8V5YOT0EhClPrez90glZpS1dfV3Y4PMcyacyCcS10BUPpTwAILdPz+3ILuwT
Ro/X7Z9qnc/ShyDloTQwSVg6OZJXm3qWSa4xzVi502+1yqi2Xe+A6RcRg5jAuHfq
K1+HwvXh8hRm9hTkH8m1gXOxGytRyWTe5bfrxJC1ILWLCC/9rIuF5f7BdxZSsvhs
zKnxIYEqwpCsfZiV3fku1uyiPx1tAk+tspRv+XAHf73YVBgfwHVRc0ltsc9llPXC
rcVg4Uji2hK4ieLJjj7Cyu20M+AIWJmFhHzBR9LKR4GzHbOD8YzFgIi0LxTic/K9
iMETsm1hrRX2ZMKPTV+ob3pMWJLgyiMe981AS5sEjI9boQtWGdEkcLYGzXES+DA4
IOjuKlvLmv1uepbjr+rQVcVZle3IQiAcmILF85L4hOYCurFaza5wYPuiepCsREe/
ZkKn9bb93xEOB4Bafhr9uy71apj6zQ5Uc2UgJaJlTl9l0HjmJ82e6iTNI3eUMCTY
wRXVQgQA24J8kOsyi7kh2fDbbDfM6zUtQQv9O45yJVwPAatl4EvoPq81Y9Dd+t/m
Hd3njCUriKqFSezoaNEs/TGLMAA3YJPNJIp7VbRBD0Y0mDskeuiYQzWst7pQE+p2
79h4VilhpQiuPY/s35gP7TO0b0Bwu4uUOmtuBGjBxdPHgKeV5DxUiGK9hgFoK7jf
ROGGydn+Pov7qFUZcjBa52VNn3fR2VwF1sNQslKMkann6DEllcJ2pO3im8w40bW+
+dKvWCBDWoIwNJgh4mTdvvksVyKealPpUyyAyLZuU6tzclf1j5coDOZZBvJ1Pe8Z
sP5yY05LoHIUzJl+RYQHpPLskESxcTmHlGtk0X0C5lcd18xkZ07ZPlIHcJ5A1C15
7btuiYudKciVeTSPruKgfA63hgpfzdVnJ0yHrhGr17LgXf0x7bLul4oEq3YlJUmR
CWe2au3uFu6HBSRv++/LEDnSKnXl7VAACxj8dyzQsAE6dRCt9HCejIzTMOmN2HS7
QflH39iDpc3/o4m256DwzMPvI6JDuR0GXjpNZeP4lmPfeQoPyWJJtij3I5tgty+J
aOMel5au6iWDOK7MrI0Xhg78SaWzg5uw+sD31trIlzKNXlMxdjDS/VG2GxxUcKSS
ColPhBA+8NpFohEv8ONguokveGfwU1Q8BAqmGDyv5wynX6IuiFEwwmURw3lNMu3Q
90830iesNNcRqW/V6RHkhdN+RrsYHHdeUby+jNaI0pgECJBgsL3ikh7x35fIeuuw
GlHdeRoFtYwU599XRV1EkhlrJDCqXs+O0lKF2+2BWfva5PYxVBxVnnciiQv50V4C
/8PekPAsMtmc1Mk+V03YKkAtE48Jd7aqdvPFgmW8NaVAQ1QIbLHULl3xYZI1cjY0
jCpw1YbeYCYbm5sUknV+bhZQy/pJofn40znqfrUpsMHcYPC911S9xEHhOulCLDSi
PWJUSYyoUErOQRB8ad9K5gLfPvUCCCxV1NmtU3E9M0nBpxYhu4jiigwcVXv+uR2y
4urR2GMB6YoRa/pa4QGqhaWeLltyzVInSvTksDeiokcM4L+0zOYy9PiGmQ+yKbNa
ckPVeaTbtMyQ+aZ4W43jcm7K/Gwfm1Mqvl9/4fDU1K7CPV5S/BhNmK0hgjwGhI8D
lkCHo3RfLqLjgKzx4Nsp75/sPe9WIyr2SHTIGQP6Ve9bAx2fa/A/MEtalVskT7QR
J4Y3Qa9tobYGMAn+PN8xP7nVXpGmYyMMdu8Syk0uONRkxWjFR+ZaXH/EKjS0PPPP
f0XuusR+z5MJoyjunjj3bBYSv74kRSandb9GThRMmmhirTVexRqwAMfGPra+WbEM
0L1R8qg/n5LoBcoiManQd/z1//gpnssYk6zAgCD+hwDJtaYkDUckn0zqm0iR632+
1y8q37lApmiCAWjdwiRunCrr2uTeUaizE1TntO5DviGk5bd/XCvHqJuuEv84vkjG
6HudKw0+TqryV5oVYq3F15t1FqzzrMYeS89N37+Jg2DRMnxVBLrh3eiFvnrPQa9w
HmnNIDBA1zrVBgI8PvLTOYlq2Qk2p8g0207jQZwLo2IOHJVSKHSYJQ4jGaCz+W+L
FtcLM5E1CTFP9WQbhfUAbgN2WGdxuSkVMecKaSU2CvSFVno7CdEjiXWNv6hgTwL+
Mscd4vthAXDfMXlj8eE38uDDjwQRkDG7wIFmtIGzNetlA3uEZUTm+EUjfFKdU47g
BXDIhU/gT24NxTyiGBePNid+kSIHMTZJuz+/HHraGX+izCCqSl8e62TmiOi16OKo
3737bjxV525DEfbxxEbVSJGRQH/xEOvl40k0aeA7h4cv9AquWkvylUjx5XqgsBi7
5tWxZ6QOTNLhtGoB0pSDOeslM1QA+30agGoIcVlhaX/Mf9D5UzLufhYugTQxqTOh
hXlquVchlYdrgsrYhOXeuOThJU34GakTMTjwue7gbU+tGYH5KxtTfsVBWD8BoKDu
IWeT045+oR6g//hXU62o3owGH+nM5tqVh688RKpIbMD5qaTkg81vfr8ikx3pJdV4
o9BtEOMUP6HudXO9s39PHJ+u1oSnbMtcbHutpLUR+ygrGpT8lPCrT2g6fslChK86
KcpbTLE/jHvTb5IzuMadufp0pHCSdii/vWLKxykTl7FEXx05xnXm1xrzCYyrcz9+
demwlq2JfyLkWkF4m1sCEKCL19SzWHfHtfaEcZab/o+F9JYQuKNvAw2HBKY3VtSN
826e3WUsNxngg11172sb16MlR424fOyGj0vhKLWKtd5T2gHoIhdYncJDshfxQwop
DR+DtyS1oaxrPgagxRK4epd9XIKizSK1HefrlsSsXde36tQMpbv47wQM05yl7aME
/Qi+IP8LTTA8DzoAEicsgAu/o7byPj42oyTJbOBX4kUDzgB5V5oSYCxYQwPfU/wS
3n8g00MRy+MS7MQ9bCXS8YEtwJqni2q2CJTadAI6VzBG7EXbZRD9uhN9hvOukdvV
fcCtpCy/Qn+Bok3rLm68h84y8PlweWxxBiRqgU9qjv1EcSzSZqFSxbCQVE9ilZES
69sypzjhG+SqO0CT2p2Gad0cYgtCuYxAHqEWMb872wSyy+WI/W2AVgHBvWsLj8JO
jYWswP7ZyNd1+DwUIjRjGXj9VGv2+mKRZ7ztlcW7fMaFiyXxAG689+LqAl65H3We
yj95ztkhlRkkX2c5gDdjDKVA4lbLewyU3TNp+FEe1Iy4k1buGSEuXHpKalGWl1HG
qnfH90M74XdQUc7/+sw2JSgLweMemj5gmQv1y5d+nhHBZrTRsKj0W/7pcMSMW77Y
k8x2L5dIBzp6CH9l9ARLFNUema5l+5Bghcb8DYwiZ+qkraTCfvN8E7zosiEPZkGr
iWuQNZRqY3zzQPts77Fc1CBoZToNTFMdiv7UpAuOkTxsz2W/0Ryy7pm5Fs/+0/mR
HNwTLm14RClV3nMD5nc9wb9eDp5JNjqKVGRvHuN9sUr6crbRIglC4YC5rtbZ4ON2
M/IM8yXtCOGE6019oILIHWHbMt0cjTGKwOqqF4UeMYQiRY+rOL7nJsocYM1ZkETM
ZO0RyP2TrejOUjEdMq25614pJsl76oTL4GXaLL1wURSxZNf2Xr5wu81ERtMifTMh
Spa3koOFsV36BFL6tkE+OU/f3KccViD7/jxc7qX/BpgsjyJV+iHeIwe048iAZxga
wBk7C/vFQPlYwq7OqSFLsV8PnpFQJmoibEry1EgLKsbv/pZUecVVdoGaXaUzGwl0
F7iSvGjpyQwh/sRSysnfIYS7Ra4nKrndoEzDxIDOmidzHewTVzbNB0CUsQrrVeCV
UwLuRsLltIHRGKn2pkabTiSKG0OMelzXHhDVNyQLcpPZ++KVgj+ClZKVrDFq7LmG
ybtgGvOfDd+pYd08aupChGoOSAQbL6WlY34pxol+cSyxaRIKivddJZ+SF2yGIe0n
CZLKcVYB7h0e1UszXGIzFHkf6gsPlliWEk7Z7/aeiEEqEMpekv6HoY9iifjMnQGb
5LIBTzhVdjXeQQNz99PoE0VdfU7IFCE75XJzuWaD8qxHmwA1FFBRjFnHLK/7ZUY/
p8FUFuMIkxdTj8pVN8NqJKaTltbEuQAKxT2rtP2DJJj8Rj5ssfmmKKjDwqUTnjBR
DAR9hvA9wN3nzRrMett/Vj0U0GloMiS6ao+iZhY+a0CdvBgeg/1yVtNETr2P2Xo4
BaTJT3zgxKAiY5rQOaC86Yhpd2QJ9/O+a5hfbsRj3LiUNIC52QbgXdzQeH0PseHQ
BLJSAmm7YA1rUOueMK4rSOUqXtgk36jdU8efSAhOIW1EEcMIdocXIfsNUqxX0caV
Wj3SMiYiHmbkS25vFHGuWUFcXBJmmajSxa2aPGBsXWfP2a8QsAT7eQWhXs+dnSBC
aVjAjhFFMbmAWN0KUwIo5xfETzQj2Y3696SXhGZRi5XfTnPfxsFCd5BREegFAs3F
kG60GNOg24XQQrRNJiOfA7OAAsmnVbqT8VLvahPxVGj70/H3qjFTas+bjeGcKat1
b0ThuNiWYuhxjv1gVQqz/xYY6mQp5TAUFxydEKTQUNLPKaPtCFt1yDy9jsoqbDPh
IW9AI/nxNfd3hLVWM9AlJxFjYQ8+FAujfiUz/uwszLPXaHhtT/MmDcsxplefI0hq
yjbRmP7OF3enJVfRQbRruV6idZRMuaUGlsCiGE5QpsbcxxrDR+T3BZ00JpHhmWmX
h/NckHjNvcnrYhLNvaDZ9WacnATHGQWN/IPlqn0NpikgMX/rcm9JDWuzoBaa+AJF
7Zyo6YgKDIppShC+nevyIG1lUhcYj3He0cuvL7AadZFytqK7nKIUTUk9o2xN4afG
L2X3Zxdx14Pn9SGn59ZA7uAn5Vv+ddgtqSjXKbDAV6nqqIY2+ddL9xkAYdm+M8vq
lBRvtJm5SPYYud5UkX7SJC3u4HlkgTjQZR4zoJJAIt910LJ5FsEAEwnuo+q7Yaxb
Iaa43/RR/dOJNAnDJSAvJLy6SeoucF+MGi/ZUe2uKAAqQic0aWVUm3XDdZVoSB37
HsgVDuZqE3S2IB07TzESkn8MsS4nvZVbNQfnQBxjngf4Vkc1bFz8ySGZQzWhwyBe
fltN15IMvGoXGvnNajVFWc04wclF/qTE72tjreNFavdyiGb1R+BWaFHH57+je6zm
11MBho5oS5eGtxFO9o+GQ8Q8iiz+kPHwphhV+7fuO21WVKKicajbruwPwdrUmVXP
5va+WQDTCvlhiT/KpwhJtlEJJRlYF3YQUkGqmEA2jmnzMkA5JhUaYc0tscty9wJI
+hIIbj02Dy2xODp+6Ann5jniYjmU/IVOLelfHa1zVh32RVV0nLUmC9al2gANu8jw
jLT76W5VWylFjFTBAXqY4vjU+vr4HvBh62IxCMasjNryRRAD1xVrui98gXdDhc8R
QO97peCHaICsN17qukNPL1SnIAXx6KGtAcngxqzkA95uz3ebBjl7R/yNDB6X3Bc6
iUQD2KvhWssyeLumTZ0CQ/Qk2t6Im15XoGyEM6TldN7k4jXkf8lnA25FMh5oHTez
4yae1Sy2uzq/iaSy3yE5dmtRQ6b4iWkzQ03pJxhwc1okKLNF9X7W/pOcWDB2xkb4
tMARG+uQeUtgXUeSfdKDqhQHnkgvWDoybNEDxdupti7i7phzi94NQ+4zX/RREiXF
b6UmCA+Vc7IZbcTtzJN0Vg59gehxRQpDXJlcg5WUJQ90SAg4g8cIYM47aMCJpuA3
kC/EKhq9qOykI0jT0SLGx+WEJ5yM1+zeeDurrwV/7g1DxKFcmNBgXD0WH5qFxebA
48Z8hsKq3eKwIme/3O6v4DFGPUGWoWkmuK2yHniMJE1RgoJjtqUbmFTMSY8RIfs5
PBhqy4AvUk1WfdTKXcULCvEOKQaRPcuAm0oLQ/ZpWK8kNw0qJ6bdPcCkD0xlP7MO
ybJsE+mweivRjtankuLEFB3Mf5LeqG1LQkp0cZ7nHRJQDwh3c7JPYdJox6lVX66K
P1OeIhbQA+rOYkoKVKTKriZH8YbxnxVQbEPd1D4w71/tnQX9Ms6td6L+5qfVZ0jk
Vamky63Gr9JJZNX+Y4HWm1xc9R9DkmRtp6G1QSUdwTXcgiSCjhAgLE+H4WPGt1VL
z92JCmumbYCh5YWx28qBj3PvqVmuljN1wzTp5orYgx3inOSE+wi0Xpnh+TN58zTX
8wgOkI3caZW7ySDpHKkYxfGJejJnM30YyiqLz7pDCPU0LQvzNXrNDsvRkXL5dNrJ
kcqPt/lLXBrFqJYuJ7RNM1VGzqv8WUAGE0NGzOKKdP6GzjSSBVm0VdkKiMZxdxmT
QRnI5hf7/JfBREShl/YmkA2J4wJnVmJpvaXj3c5EI2PKAaQQ+VvBTQ7r6A7Hm1jC
FQI+l2gQqpM+3EPU33gFdWNfenirELw5f9vZ1BXtQQJ2TzUuVy2MbXUj2WZv6rp3
3IztKIbmOFu/4B7qImNwm8+9ZtO1/F3vGX9sq4Uzn2UOvaRBac3o8DsUdLy033mU
mXwO0RGPfcfmnc7pnn//8rbktdvBiQVxeMn7VgnchP59jc/kxxZB07R3x8uXqy1z
OMdYQbSTueyXgE4hwmM28DEc7qUrpb/GKXrb8U+vKk1AOoBCS6WCXks4b5bHCpTe
itRPzddYmEpIZVdlyBYeEbuMBp0OVrwogqQWWQ9R4UXRbeLeGTcnOjWSPeJXI7Ry
Xhf9F0+l+TmWyLBxws/+PDhHcIJrjCZbXcDK8LXvIWra9DAzwp/x4V3J1s/wLwS7
V/Iqv738xsRjz72UYp2faw==
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
AGfdWbD4bxDTsj5h1ehLk4Ej09x1AdOEsoQ1+52vxhDG734CYvlY0sLLGAVRb23d
I8Cny46J2XDxcJpWWA+5uyQc5RiYn8JQGGSG31ayPsg9mo1A3+iguKIvlwNN5NKc
I1FgXyHoQN3TmiYG7rS9hxOCDCExdbFSFmHgafITiOWYyXmCp8Fs4A9fw1MU7sbM
wgqM9PHQ603pz9jyAWTh+ZXck23sfZgEV/jyp5AvMfe8oDOh3CQ8/3HYAlg3cshy
0csUvBlVO7LGhH0wOniV9t8SYHeg3TGNuLNsdLNAUQW3QaNEX8ytPQ0VKNzh66ZU
X7PIiqJK09EKW3zYYuMFIQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5104 )
`pragma protect data_block
3rtt/dgYltxSG+RqvKKszguXCZPBtD8v7D+pYAIAhtItCUZnEthHbu3X7EF2b0oc
mTITxepPJNGb24sXgoj7bWUKuvanSmlPn9KkzRNWX6lPktepceYFNsy93KWFqiTQ
SS7qwl0qt49+p9WX3iduEzhcOMaSgXSOtPxEV2aBstfvW5A5N9p09WwUIx/eCPgV
dCyU9jsGXpGPS9YARY3Pz32Sgk2e3LEG1YjFExRxN+7cE2BIEHanbKSLnX/koAa9
R3bd8KZFJKjQg6POT6LdVbKL3kTLqteG15IzFaXgwtA22LgcdmngxSDuG03YZyIQ
xEgm+USuJZQqk+SXIe98ynv/5MaUS4UqURN9L4UZL08ZFWn8xL15AmfuHMN8IpX3
ooDIOBml3qsS18lc9m1KZftdy9oXpTvptFJ+j5MVcYj3w4UboN0hgL3IV/G7OTaA
5Bet4eD7usamDf0w4KagR0mVlS+xVgnctbW6NTom3xTshJz5qfA+FSq5+cMH5NAB
F2joJe/mlU+zVRQ+emI7MZBn4aTzzTf3HmMDVCdeWyLOyYjXvghQlgK2k6pL3gNe
nBoR+dzsp+tWLr6zttK5FHNvZE4PRbo+fB7artuPxxUjiKyune6lyIcg2ynUyM4v
pad4ie1qpwcivKlcS3e6331EMM3Fh6pzCp4BurTrjmaDLVanWgOndK5Wt5zrusAx
QlHcaLOjODxO4lvaAomNyTS2RMiRrHFRMIvPGh2gTNxDxB+s5M6MYNRd589fcsBy
DqNlnBlkt/QkLKLUJTNbbfW/d013+dWeZvjVgg7Cc/agFPmr9w6T5Vw6CcRHUp11
2UTV4YZkKXfRc+zeY7faRGXWNSKYypHrQWhut/3P1p0o9s4MNUd/XghCHvOqgblE
cuGPyT33OLrBETZ6zpea7NBZFiupqq1+eiRf6mfowOR6xmDb7FcMK3Y3ZqswWAPO
rUKdRiWshixkHRoW0Y+5Qt8jCvSExt9h/5Vpq2cfWOTYzbk3YlqqJ6cz6erQYFkM
1su2GN6Zd5xREiOcV4jcVB3hbq0yPoIojSme80UbiKI7oRcfwyhUBjrZJjawo8Fo
HzMn623lc+BV/rQxkq+UZhui5Ed6AZmO2H2NQqFp8jddPxgw/Z23gXE+ywk4CFA8
pA97FWh1mjWh90F4yP1oZeuZLyTSej4lnZo08gQ6jrDZ4RTzLDBe7cklylsU5eMo
LmBDcY8rg1iGhbpV1Zc8v2GcjemUGJxjElj2RptkpU0yaWCY9haHNsD4DoEh+Rxa
urC/l7Q7y+7Ahoh3ux423/k/kH65rfoI1aVXLglAicS8PmK+xVu/7Oyh5tvtEuvU
+JItuoc11rlNKJ8LA1N9J5nMluMxUExXf0gp8sU7L6hd5KusCv0hxt5EbAB96cuF
C9Sqhz9jya0YSFCOdFb+ohN0PeeD4dlWFbnnK0GvZEp6ppmkhJqu7fAdaYZkmnq6
KxnLnMU8ahgFIvmYGtFk5+Gue1lxclW/1SZcC/+sOpoKrpmPf2qJoPuYFNv/jVmr
NoEpqGW7to1vD84GXGvLVwaGS0+AE2g6mOKNjteDvwZjk2qVqrGBh2mIxExbPX20
lRL06keSAZR6mXjIHc3pnJz5GacxEuPMPeLBh3NIC1tjfv+sCn2o6Q2J/PwimOBR
egmrm8zDZAvl3skTt5+GkPyXUY+uWbXnc1RQUruB0Q8jxsdH96kSYsU7CJKDyunL
U60CLykNO4oWxLYjqcshziUnywh1LnfZO/ciaw/Z/Lq+25HOxkKaFAcTsCdclKZj
WHr2JBeaONsLmxXXlmNlA75imFA35Epa2fzbh0Um7DldaC+CIrYhYBPel6PB2DST
LO0+rYk4l7pSbcFhE+XY1Sg4Xl8aZj4WUwi2eglnlJCZvjunaeGmWX5+HaHois5G
mSS73JgCyiMg/w3vde/FyZinUZC+FeaOhK8kBRBwG7Uu3C8u1NrJQJE6uuPk52te
M7sDLm3IVA51nmAp2JqVgNRgwJ3+ylDmsu3ACRib/eGt6Pc5E95usUPCFl04rQtL
LIFL2ERxEDu5Qd7WdcW3dOGxN9zAuF49tzI8lvuIDIWOK43/70e5AMRO4BYlxfSU
sDjXGqCXcFZkFSppi0WYA7sHDN4US8euv5vMbLkZS4ZoSrbEa/ruUWV50Se+hF0M
U/hrBwN+14gPHH5wemT/sSdaN+ipEpffgcYSOQK+ugPnJ3GYN35zONLIZEK1k9Di
svfEQ9hdJd1D02SB66+aUsw7cjY33FEOsKjfe1B6ReCdAAP92t87l1LcpdIaHzLp
Nz6Mvn4mXN/UzaUUKtOXHQtAwsEzZNiAEdDm579ne20vrgqGc8d0V3+OPucc18uN
3g2FbZa6B4kZK9SZxKBh2wg94cScWBu6MeZi33rxJ0Guyqyui9BJ1T2mF70zIi8l
7RmkCNYnLLRPOYL21wkIwWSLtGG0ewWdZ+yWIoj3ow2HZaAmbAbprTfzSwAgT3GP
K1mnqzi13jHShbqjOvQLCQsk40zOfLgxj2K34I6WwBJdfk6HSv49FGHcABFuPstt
yTRZ9amk8GYKpmkOI65tc1iiJdXrtE0q6JUhQ7qVylFMJ6KjP0eo0+4LoPjp30I6
ZHJ8+bL29yVJ9xPErFX09pxQpPkVg82i1Z9LGoijL9sjBi+mvxNvyT65CVxA7Nl+
xRlDJ0XLaVsHGoV5NPnHhuWlWd3YRhdTuZ95iOkXHMRx7DvzhB8PTgZeQdjdf/7W
KgZHjxzNJ6jSw+7kcudwYB8/53VNwGnYPlqBB9gGEPIDM8BA4IhG2Z217yNhLTf9
7e2IOQJduK5f0lwCuIeIm6ooG0RFxc6QWFzYrCLBsDw4nJUzm1VlQUV18FRa2AE7
2aJi9VyrOdJo6+On4NUWYsPe6GSWnDo+peAFzL7KEQCmpMdD0K44DIENi5P7VFYu
DDH5RnTxxDu/Tz17WR5IG+M+S/rClBeNLkOQ7sLtWU6PE+c3FDw78+LmNc/ntSCS
dztQ7EgdtzVQQJtyPAXdWLEmZnaPXzeOWA5xX0aH3crT6lwFz5/0xJesyofDDln4
KUbfAKFetNmH34au2v0Jxp8nl+Smx5rCYg2Ffa7/ouibU/f2BH3jvZ0BRcKjwkpU
4WKxdyRwzFnaWLmIudRB6LXLnotn6uHUjB+VcWOTr4Eyeej3ML4UddFI4PbujDmY
Aa/up/i4/qzVrPSt6OhChXc0K9fvPywDFUGkgsCrtWsb5HJv0p6HSvDCyLkSQzkg
mvCVoTD/jX0Xys4eZZAhUkMrNFEgnCKL6sW2PYL1DHXUX/vAoDeCIH3+A6Bk44Dh
YMqvhZ98YWRaIKdauSI9YrrhBar1fAKLT7ADS+PgixgzUsMoChZAgx+rAJHsoBiE
yHWJTq7oZoqkreNu4PIHFpM9RgKLoHoxiOXJD5Vx0FlhAtVOSrPd7Dx6/8DH112h
M8bCjNbWdF+TZ330gOjercIeHNqjAMc87xxVa4BWya+dK2htqv7Tcr4HHOJTU8Oe
Kb8djzi6DSYTMsM6YP8iF8xSkKKQN8IFgK8EOua8b1q5VSh4xHEWNhL6dX9cRkHJ
DBMghuBiZdfboF73BTHRj5EgqCqJh4YyPOzWXS8/I+ud+oUZJi+U2jwtc4lVORTF
2j12QBtXpn6xHqY+VUOQE0SUcy+4pD1bVgfO0058/m8pi0w0+YjfBRIk/ZFv1VM4
RrbRXqeCyNJ8VkDGclYrTmNP7etXKWieZvUp8Eo6owqdg7j5VKmB4dLcDsgUyrRn
fmmH7aPAINHc9eE0ZDOqJJXGtdeBmLR3G6c/LQlQEBWbW2rPJyarRwXRki+VF8AP
abh/n+PNlLUSiHDk1OYt2Xp1Ztkl4WY5CIO1lnj5mQR857b+0PMTIg8LvRhkZdZL
BMkJ+JkiA8KCIxyWRq+GEnhF6hwaE3+n+SCd96PPZl1Qsp1dddIPa+Ox4DqPsk4U
V+tJFufypf9Qv9zTQ2mMBicviI2CjJXQbcwLLhpuBGG4//O/lsSVkA2/aJtb6R5B
PGpclSht4t4H//3n5+g/N7lc9NgAT26Jy+TZtmGmd1IiHH1kJUXARzSHCgDiEeof
vHhu9ziCctfpy4wW7gq2Luz1ITVKZm7vFNZXN/NzogUlPjKJaK5OJ6xu7hlObN4f
VO6MkvXeNDgyn5Y6iOc+BEkZcJjj2IYpOOcqnQmnS8aK4HGachUfyTERiRbwZbm7
XQJmjN82c7VztqXsC9GSa5gUJiiG8JMFCp2hhwMa+S1Q5ViCFbyS2B7w8dDmr3Na
ANYRwcy9fAs8Nyf9XlDYSrToaMq6Hf4GdOkrGaPsjBAa71l3vPvWzUGGaL8z4gmz
kSTSn8zxBTgx4/sVb19NCQV4jqyMispDf9biEBdc2ybiYriPwyZLsxa9aVX3cxuj
Xz2c8GRQS+bGTNBKCirZbu5Xoh+roZ3VjGYsthO+9mO/ov/AlOuNXgOTITQdLim6
+IG3nds1isQvRlBXDwyLWgD3ajBLH3pkO1/xsXwlJQLLUf4FLev5L57atAY4KhB5
nzsMhJPne+AuiZtMHipENoKGJFQVi31G/JE2RL/3DgUiKS5INFGaHijJayB87US0
qO3iqAzLMroMg+92n2v50OQydxqvZJE8TXUFVzdMZyEgpvlNBu8rbS1fbJ2L7r1l
GbF2nF8L+Ybox0LOmNDDz1g5ksWZjfSktXWQczwEC1vW18livwh3qtNk5JM8FULf
SzZxzAHS2J///VT88VWtg7OADYtikSvIcwCuVTS8KhQ813UeNAebqDCoTVWUTVuI
DaYX1DR6V6s9ltk8K9QqqEtA6UC413nOKijHF5ul0dqlb0jxxTja4fPWJbyot3cW
A5n3SiIMH/J4wyL0aPQQ4wJ4aP5PHkcAf8BduXssWX7u3uZbiDTZCSfhX1phZjck
YBW033p62hz8KzYNkp6VmspgKG5uVDFuZkLwWCx3yLmHQyY6uHojHpAVzzFE6uT9
GggBfOJFCTnRGJ83sZxCr0EcABjFNy7290LQ5EktymE9v8ZGIaDDWPt+JM1qxQV5
4GrJxHrEcJp4Mc1fdfuU/Q6lRq6LkM7OnqkwiQlNicLAO9yN/cI36riGSWo3OApq
0VXZjtwjA55gWUhAk/WzFh21U65O/iK8Q9RrQkDNZx8hhx9Gnq0JztcOljckJ2kx
KVYttQfHkgRRjH9rTxzBQNBcPdIuo1sQHxNsd5uNIh0/AlwOuKC/jsjyDLd10lk9
EPGaLbEA3jkdSVChgXSpPgNKpfGZK7kbJPGY7/Y4u70SKNgvtW+4Bq/5F+SmkyyP
0m21v9qiW1QiFIFD8NxwY0yogaOPiz2VAvsCKgOnQRVMdLU2rOgDo90oPO3kRS4y
Z+/lNfqcq9DsVR2tS0ag3UdvVY6ydcWXu4jXq4pAZtZE2lWBd7w5Ld9lRrjlrBnH
L85k3E94lsetqYW/UL1+NtEsLz/u16QcOzDsslvNtpppvYqMl8PNXPgkVZF0PYZo
mB75H3bhG6D/pr6gOjbxNBqXoFVkiehQ0YQdGcLsq2+lHo7mNlVOmn1Vefv9ThqI
6iLLhVB/AGSKPMDWwSlQ7wJ5K8IMX9oET3VtE22WFkRkW6/db0aPrSZ44Alb2QZo
Yhi8OAqVHj6L5lOKOkkt+arOJ5kyf7uGr33XNESQR00fc7i1sz4hEUey94949H5E
Gl0gE2uhvhjEpSlNjdIsqK8WwpxykSJV3RheJ8Vo+wDtFTIZxhRUY5v1CfYAFpNc
CcqzPpfzgn5i2SuksUzYL7bL3V5BrrT5MsySTzlgbyCLD+C3Zbllo+W44d8Kwux7
GOFzOEOSaBLusDOh1pn9noGLar6KdA3Env3XLuqHHIRvBZ1aDwPkBhA6MqK3dE3S
C+mNbm4Fz4oG/Qn+EZW4OMFQyGTk6BRLERYKHo7g0v4yyhdtyDWRnjsqHoRC9Sd+
pW3z5ncZwoAkUrrHDSTaERTiiakhuaDr/rlisBPsLIq2X3dgp+pgJ3qCD1mGQSFP
UOHQ07kYCw8fHBMC6QpBW4JNVS/LyTqMZiilT/Ld/At570eC6QpHLk6FprehyTcV
LLiY0W/9gT7r1oh87dGzAC4sR43lepjPQS9Tj5gTBD6rfyn5ilw0b5rq6VbB3ug/
VZRtC5swpleAGnvB+gBimXOqOl6+tk4K3WgQVbPeNrzG3ExwMISTiaHiPSzmMNN+
rnzgp2ExxKTYbL+2QhpI0iAIlMsCK0ON2NRbtVcqFI4MZjE+fRB2BGZBs0UCaSBu
VKbO9doP0lItNlYv7SssMRt8GuYOHbF5b4LYvG7gNX4/gLz++cgZGCq0ndseD/cl
bK6b70LtloREY792b3ZeJELF6WxutwzCvnxS0sXr5WF7M6XHpLsxvGDq7DEjJhwD
o0xkRBVof/BOPbIoL1T4rnJU0eFFGjBMYhn727LH/H+mNjrhMaTLAlOEGI/DvYJ7
TPmJZ0oe2hpDP8P+HqxIDZ+U0TjcDvQveVoiQGFMnpev0hE6eflJpNQLT8zhqW/I
nd4P70iD9HDiU3KKgaS30k3uliHqTpH/A3SwqVkxvsDtkE88JrttXrHWuK42svtx
dQnm8OZCjdeiaxz6+FZLUIdB6uGd0KphJbqUqzXLKE/9OwIYO6t5aB73F4WKiQ4g
UlPbP3p/NN6mX24V2BnxNnvQggMqGfu5oD8J1PLeul6Hs0aLumviBVJ6Rldh6rRc
4//tPKZImKqejj1bJss+ELSf6LEUt1PD8VaZwA7qV7JsszMydY8NkwheZit46mj/
rXZiReo668SuxBZaK/kPuA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
axLReZ78g+iRnCA4w9H0QLjxiVIz77jGybAB292ymVuS9sZMAy4lxrix75ZS5rrq
k9EBsDvNrx2jq8z9e8EzokZfqpWQHLWQJmuo/vRpu3qs1CGCKjAKmyg4AzMR4sUU
up8rXvAjExqBXzkziLO+UDMKb2y6ap7YceZrlvbzgkXH9J/izr2bX8O0AVLRbsl6
bQZJBj0eqBSBKG5AuE2qzW0dsucdF1un7y+Hc0biFLtnFFtfFWodfUMhldjY9TTL
biaAbMAffcIp2aTGB2rBsJMgYAYjjqQW1y08vwGgcs2NU6C0JNtYQRbI+Zbtce2v
Vh+T5oQ7EbNpLG5AZmiJ7w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2624 )
`pragma protect data_block
ahsRUsmzmw4vqfz1OgyqPoqB5IyJIA8FR7YceyH3EDc6spz97NGBljmvalrOnP8m
GLFBVyIauR3HiPl+cuzLKHGCVP7usYNT4KJEmgwunuZ3XYkfLuF3tL3yTlY25CPv
lftwiOhvpUxuyvDPuCXQH4FL04VGUqrBsI5kQJK8hMgZl+n777ei5EgBtZp3UQEA
bX9b/kDSIdcyCwaFnoTfwH8DiX/01ag+XSEeBn3375c71XxSmeXA0fr52Z2xC90F
lttPZpeJZ45sv+tsj9fpJzZWa/H+OG8vkYrH/ZuHoUh+a8rmbV+t6qRQttsGWFH8
3bw7Hlojhz+gqmIvlZGnb6AqGoYQy5ioF/Pu3CpywaovSDoDMykooTtKUo/z3gtW
aPfy8/Yz93GWMqsto4Acj6gbw4crF9QLRDQcDAL8qd8DHC1wvTffO2AagWLN3hWp
1nBw0BGZOv1a1HMM3ghb50wCi0nFQnoPs5Hn2ZcgT0IWgTqTQtlM/zLm8knXx2lC
PMhyub6mKLl2tghg9pr60rXPE38tsEXuSAO61olU8yK4qgW7W6J3knLCYQafQvav
5T59V79BUkXOAkTGvtWtR07vePlegRwHWU+C5vDCE/DagpN3Y9BIzg4jCXsVPXi0
EWQJeMxxRnU8y7hZBKkvOyXd/CVNZoaLOQpqpropZlL5u6Bg7V27HrhR0/6vWI2L
7l9KDtQ9GMJU+6DdXOstTuVYrW/YxqbJo0IKyHJMWbeHIZxhXKhMjAONKT+lnd4U
Pgm0sm7/ExgF3Ko88Cebj+4QKgQY+msxYHcCISS+o5E4gLmqslERyZ5N20R45Rn/
Xw2tGHDE30Nqa7NAbv0pscfeLq/gWc6NoeIQByIogItjAdH8hIWnlhqxA2UuGcBm
wPBzjIvBqWHHycP3+I45Sk5MkMb6q06pw1eOHCSusuniMtsRWBWvxDjBd58ZmXzO
9XgGuCYXNfnwUncNhrabzl89Sg3uv9ndmMsCCjhOcl+xrZArfff2ZUUOx+bgqRDm
f/O5fANBgpXJd27VMvHCskr0QyxMdP/DufJzil1YVctcSL0CY840TkBTOz/9xoHf
D5mjV4T6eHmAAOf9eRQLmBAy9uqkijwr5rNqYNneqqsozjDzFxwxIG3FIwUn1PY7
MCI4mdxeXpfodyJuYW5CZen7hgqtIog+sDaLI+jhEtfQfWaC0Y83+dukZGzhxwZY
ZzsbvmOIlkCw5inCViuJct+uMlaWvLVecQCdAEuJ/rSKxRGI9XyOc7907WOud8qk
BkfzFhMgy94J6S9gfM+VnLe6cDLpDlyDzo00qGnmIzH4nHuDHpLoKk+g0N/zgN/3
JHYVCIOj83e8olEGVTZ1JNIk8xSCFzJ/P1TKD3blzF04VzaUHDJpV2vWurSnu4Wj
SL1BgWF7v9DIgR+UAIPraASG4+TNX/Pjkq1KNjGZdtdmk0uQpWMKQP35VM95hHDb
+KJBxel8UMe7sw3m9Vek2tHRErYMArG7OqXQC60GI43YZFQL0fJg5njwZPANDIh2
3dVhRtLJ9Ai0WfI6C6YxNs8gJOZ9Nf5B8mXwe9p9CYT/+vGA2VzOO9pDmlNW7PpJ
PbS5ysYwAap7omoMt7TJVEcNRGojXeX9KHdkA/RBfS5n2vvVH8FfNF21oZfSQWw5
ktxqmIkH1t9nFysOG9OyXxuf48j4hN9jjZSwZJNTTZhJ1M8dbKerh1SSng4vC6o2
DaLflLgOw7ICa2MOGMPTmcQPp37wBuYUJU90byynNsDFD3+swu/dTH6ET/UDA1VN
7iFXLe68OgyRW+auRmt3vFYyh3kYljKgO+x1u48kE48umAj6SzfS17ntBunLg2Nn
vD8qpBB9wqJ19REZKl38eTJTt0PUhxgR6SASdNE8FZ+mGfIjTIEVo588bZ470kHV
breKpOcKbZudlT6MYTsVlSA9SA7AJZKYeGXu9iPnMzaXQETlZ32BjnbxqTU38BJT
5V2JRVSbXYv8ENiN+vWwC0wTBDBtlvhPuEkfP9Z1fZMY+GK4Z9txfdv7AjGDUO59
moMKo09A/K1dXEVlbGDfsADw08+XAjmqPsG5rXD4v2TyHUWF+PhcetIJnSRejNAO
TXiLCP8/i0N7EB9cFj2+bXACnt0+uEjmr+Hm9hILzp7P3iVBttnFEruxcTZcSfy9
QPzuR3S6SeZuoSc4b6jSHP68i9fcBUR8JnKXic0PIoXPtQdozrc/0iZj1UsQuvPb
bwg9AmpqQW9COnRm635DzX02K0FY1sy4SGp8TPgd2aJJkj6s37hdjfVB1/pHZkHK
40KEghbW8HcWARw08J6nmE7jWrcLKjFKp5TagCX0J/FGWBKjF1HWVSfGmJKkaLAq
+UGYci/ZepEXJhfDZs5s2OD4kuiBrTYYB1zFeP0mC5WMY0BZwM0j41VDkhT8S+Le
ppKC3QZ3egXzxbUG7hBsRTrbYvsVWFbajZyi1xwyxarfIu4PMG0o4/29etYX+KLY
Jz0QlWtT7o4yEwGja+MLM0rk8a5ckFqHs0GL20WyZrjuN31dLORiM2RLYdTCgSIw
0JLrBj5/hFB2KhKaYYjJ78SGTOd94PbNvpz8POYaeyn83IvlfyyIURwIJmjBgdEB
XdMDRP6NUnBO94lVxhD12DL+ghnDg+6wIQuV6QxaGjgTw0K85EnsvjXv7co7A728
JwXUVtouEqsEdPYXf9BfUrU/gU/RgqCXtWLvYoG+Ddly0PNAKv3HByqtN/9qiHbO
tVJ6wbjJdMv6N6vVSb+EytxII/oM2MbCAXXwNHJbme8GByzZ6tj5Ix19cKxvv4u6
7OeS3xbyHo3KFUsfIMWzZvR6FP7EHsPVGuFcDNFkye6KGmKlG5JkuNHSGHjLqXNe
9zayV2csHjEsQ+d6PZL5u8PjyOGZtqq5tClWK+V7mINN9ctCU/ae+iRyOnQjNTvU
huAD8RlhBhulpVuVrF2NrFu1Mq6zNLOLUaV2lgrzIjLISte5Ygjb7VWmuVF25+uo
M+BIxuk91JTldEsb/UEJByveJEQUSlwbtaGujdItkbiOCpMz+kxL2y0Aa9lvlKKD
E7Og628TkMCc7CzWRyiRO5rUuYBOeJpCtkPIFXgEMFbxLN+Q13GXZA2/OFWPqDHk
eLbTiKNw9oXPs4SIkOlvWRVcrIJk5gFenCu48YYq/QXX3S4ECdcfmuPj5N60dZKy
5l6itmt9qHrEzmvXMocWTG31iIGi+3Mwad+OJcTd6mVMiUQn1/Uq86JRD8kmLjvA
GuisreyZJToaBBlowz0KVhhuTXKDGFrJyGJZjIkCpd9uBboNvRrA4ATt6TJxSUPA
eLz67nHJ+PQyKma+VU1W6iBs+UoWpnmdoMmTMcY9MuwACHPojW5qDS6y7QkFzsGE
AbdLt/jRQl+jBYK0hx/EDrfbEQFP6Pzxz4aBHMDq5GCP57jrLOuHSXrjG4rsqnv4
jqStl7gNZhPI1IGU4Ki1M1rUuojhI8bEJMdkB7RB3s4=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
kcJUbujCkEMLkRdSZaXbciiBpVOSjc1fbF1fyry2ythqKUOjB/7qBVG+lo4j1eJU
/GVXymZllvNNz0A2E8sob3S/8CVakTuqmVRdPDWZQlFH7JWDfwZ8SVd4Zw0/rxnD
YIuBqB890lrgzdR0uItB9q5qyZL73M87Le9Cum4xUYkopgcGCNUohNv2QfP3vJ21
sr1wO/jSDk3xFy3f4NWfj8n3yJxjJPjy25Ekcs+TiWZ2OS+2mwa05sWIGTvP7MT4
v+bbiD//BC62dA0n95K+SupCYcGDFuKQbQywOe9K3OI7K13LAs0ceqayZoG2E/P/
QAc4pyz8RW3wzw6hODRZ8g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 18528 )
`pragma protect data_block
yfJ/XczEjc8dIs+HXqAuC2laFvot5x5zPAZnxNVHcC7hUCu6yJ3sir1zzM1k7TuI
kTMfBsWJpKI08OxLZQitBuYbuqTxax9/ww7mtkd7yoon5Qnye1guJKwlCSqgcvnH
y71zVGx9+kNorh2PFACk3V5VDdr37c8Wl+qgf8yWvor8leHnKo6Ib2pcl5uhqnzN
fjob2mUkTYs/Eyxy2Us6EIMgh0jQ5EIp5kKXF8FBSdk+EQTqJYoEmstxBEpkQfDH
jwLvhsjNYkz3yHDFT0jxRFWYMPKJyIwOEazj6rvfCN1/KpKHkBWTOuyWONoQvop0
/X/iCPLkuPURVMxTC5G1JeBPq9xxzeA4vlL5xfndjb/PffmEEYjE/J8CDITeJvMA
VxPg5izP4mOCN0XsXkOGqHW06War3VgYw1nA3EYJOliUtEzksgIFMqswS75H457u
emeM8JEFyv2fCfaHw5k20VbkOD+P9OW0uv5WX15EnqD0ceESC3z9xLPkCNOBPd4q
TsvU7fQOGDUGXSqZTxslXpyaos1d0S9CGoVY1HEb4H/0hKw2BVImMkf2o22RZ3tz
oLdujGXEaWWyXrUAgAUy7LB6Rn2rXopIYQVFrtioGo+bBNe39xrt34ri3YcHOboi
NNBfQun3e3eVd4OQIdPobeRG3NclpUopqjvElmYWhWlUkK9uCX6wM83fdvj+nFod
3mioXSDTh6YaDpk31/CoMih9OcnsMpdJwyrDceKpkwjMCn5Ys/buN0lgoALrwIsM
zkWlj5VplXYQ0quTYS127SdZjDT6ZhNn4ZA1zMycHUpswQ07u5/yaKvzFbxdJknE
MkQSp0OsJzP24rgyiaw005ratFyApqyRlrmzccYNL1q69Vm77W6XroTlj3AweQjT
YmRnmvSUMLXC1I2vF8T1yBidSRhV30LPLBe8WECtZqTiuIbjbwtZgcmnGCNZc2uf
IeNPVUlxMiaUWYKPfy0TEZSPkQPzoy6yNi0Xhn04fQyQzpEUhxd7sGDq32meYXRV
lDP3OWs6W0D3BlBeUcv4qLNswx2/jMkOGL7dydeqljuWhu/jm47KIamBxWWyeI5/
48YZtvz30P4BsvMOyjipzZiHLiR6l6Avo3sh46qHjJVuyi7b39nbz0zTgsZMBLuW
y5RSOrveRd2YLZ5i4Sc/vWp2s69DO9Oyx5gKKgfaSjjq/nI8ZR1w9Vv6BdJx1EHR
i2c/787wmCg257MNfQ7B2QfQkVD6qSqs1xO79jIkNxHq2UHrpR4J0bwWz/VOgtsL
QDgHSdrLhEPX82SfF/rmEppzyHFAGGXo79UhZcBgt6h39xIXW3YohDjrIrpEkagk
WQHEhBgrZOgOkkSHlFSbtOtdV+OyJbZxfthu5GzKFiyxf08xAaocWFDOg7JZPl5p
dyz1hfy8/obNzE5ke4gluJXgukPHiRl1I49t6mYGer5xe+JQ8vP6AKMREfhzA2yn
hhhTnmxhve1rpIDvH67ezTNOBoFWoI1/+GSdz++39qF8GEo35u4csK6XpU8FCl4S
o+iwy5DuAudYkQBhKkTYD+P0pO1EK/r7/4dYblz9F1yWVrEsbyaqDnxm3iB8rOh8
Yt9x9qK0dgubLjetPU64uR/6Ae5Btxa/ZFYR9bV/8igbHwf0RtNBr85uQiSWOkRL
+Dq3V6nZyStpMtkentZwHPQJxSg7xyG3Q/dJfNewNdRy+zHxxtkDvot0Qqr3awzn
xALo8GyC1nMNbSgbIi4e+wP8pwVwFaWEdaIHF+eGKPJuci0zHo1QqJY8oEva7EMk
ZGdllyrt7c2868Blnt1RNjHxT9OdYdFuIhpTCDoIBInnoJVJJ7eGsLB+LUGXxhon
Q8mEezzpZvwXjgO+s3/V1MYjXrjx3jntz4dNYgldeRUxjftet9qn0SVwF30AnSaW
Ex+IZeHxowuSh/vEF7Smx+DtyuyMzaEpo5DN97gvUhmnTqoUw5z7emDK0w+DRma7
213FmWY4ec740qVtl0x6UF386Q2OGTxsxAkelG+G7dgFn5gJdWjwEbSN/Z7Aj10U
D9S+cfIaKUMtOf5ahWzlk9t0VDN3H+V52hGYX0UtKcae1rsevM7jE7gIQepbIFvf
5v/N04KvucebgNHmsP8XvcqcH2tgKu0lEwaogCXF1DpbfVILsUSy0daEniw9aREZ
SV5TUeDU/1rnJKN6/V6ofr54GeVL8bLEfBjKeQWP+J4lQZxEZ0lZ+dxhQGXcR+SR
t1aGxuJ2JVdIfA39TLZAH5XQJjyh0fqy/mFqUtR+DXhrUh4hYJEAL22K8e9h6ADO
N50qphnvFP2EuYi0N5q90fDaYv7cHKrz77+XpQBHCbRdE1ARTd+NrQqpXgaV8J2D
yeubzzHR7ZfcWNWzOWqjMBlmESuzZLIIvGsGNhu4/MPJLiiFamWweVRXGWdhsmJK
/EO4HRp7Ll0Gru8+RdOndddM2evV2k5Z+Rrh7OWkab9506Hbl6G5qAmb48hp1vjr
siQpmKWiRRNt/4B68OD2V8rMknniLZBICo/kGT7eA0Weskj4evHMHL/1FwnfB0js
wf26JP0aYElOAbttLZbMGrVAbQSt9w+qlVtRB1sqh9ojq0lmnhVSwXhYOfcUmUtN
od25qoF0KgOzRq5jR0iwtR3tj2VIG9CQ38TzyvQhYaHoIrTsXfkNpUx8c6lowEoH
mVNgJqAhvK7BWPvLJU8UMS5W1OmX5TBXQO30KeKgO+21fqzkCSPppMc0PePq562o
PXLm7TOSUrmhT0ZuAQexbGuRlvuf7PFr7fsytNhdvmpNKkbYNBHQwMH7g2vs+KtI
wOghanxu4CsDWnAVwmkv68mD+FIZJt+2PYJh7JYc1238FSaqcnK0A7UD1blxbLlF
zQYw5BJi1c8Tfi6qFL9omlrreJk1QBJfcfkPjR0mizD5EmVYKFvxTBmv+2cchSjY
bbwNJ4euql/hSrHaHE7ULjq8cD+Und0SFP2MdKlaFVGHOb5Bzm08+Z3uncqRqO0J
Bv7nMdCpGICPVZlIe8AsxwrU1aMfqn0eyPl16dBMRrubxc5cSywaj9DWAgu8Txxz
tPsMiB6H6EI8kFhcmSgWzNZ0Cor1fCxRad3ddoxRnC4fVVUvfpOHVjapAejeI7LP
3t1dDf6yMoz3v1sibzKknvnAbnMExK/S+HUOSi1Y/Hs5p2vwdKI03el4bRJR0eAs
s70X2oQGaKtdSu0qmpsfizxbu4+cusgCUVbxCSDYYadS4lk7rY8ZcriUhTCRGjDu
qnPg2Iss03ZW4JxcUnI7tG6KQaxcNISzUS12nn+Sb7U0ygqQ2GtIJ/5+m76GVpio
wpCInzqMfwhd8qvN3nYuHbT4qY7HUHcTCkLrMNGe1TlJY5C6/nmI84fh1qf8WeKS
NQJBpEcx1kwjnyVb+7hyw5kpPMV4Zg2TdA0OHsujy0foBPO4r+ss/h2qA8PXtBf+
O9ANlRfRgzJWUumlYlWqObw2ERN+gFzY2B7KGk/iRQrQG0Moo7jvoFM1QY+q/HlS
pseYbJJzw1uN4UQB/ZjWg1K4BcdhuWQaJToBozZf3gByol1YNpBMLrLuX3t8twfs
X9OjJOoKuC0ynVy3o7W0VbB6A/pMtLfyC3CafCcZoKJQcXgd9NHw7WJ9kmcujFx6
KAgezmooxqDD9WlGpVBwoAbrbGuG4/ZT80BbFPHvuOJL9ALblnjNozRGKWgXIuIY
5AqC+FypXWWcnv47zpOG/Bcz7t35xA0+0ccRqBXjXL/m4RZcPupi6jZsJxO6jmYu
1DDBLOCsWPrtO2QhNdXhqp37gRnVqRzVP3rC8GnFyH7CntbzYzFqXIcL2396Ukbv
RmpQNPpgK+OLS4UKYF7hjJM4DGcvVfiat+KhiKAXHmmxseS2Vpb7qGTYPDUNlvs4
MIbbgTLAWqt0o9KEJWMmhy2sKMPm6rTdiqSP3rPgVPTkYK+b4p+lnp/3BzX2VomL
I1CPdtQGVbZ0dyjTipGPgK65JvWJazzbf5CzlOeRNOj2oTZl49IjpKYL2CoyuD+I
SRxdnuPvjT5w3LgfiZsNI+OcgCddL/IeYVX6hvVG2p86RRJRy0i6CmUUbeR6nVdv
9asFItHFGvV8JlcqmPCA2+eTUBi0w4fAiUuZZzDuKbVxQ760XpesdBHpcuNgL50H
0ct6lJBFOnHM56W8OB4zde0EBF+t3+uYCn3dOomI8kzVQjNHKnM++R9l1nX+libc
d8x5AQUYebbv3l0jwfUn+vaSKLzjS9h2OeiTvgQmXgfE2N6WQ/bc0+d25cKrXmlb
9egsUEd/Frz6eCtJNqu1ohzDcaeuaTsdv0u2panNLbpkIsYgSY6bTtcIjBkenCaF
ZQvKg67JzLqzi+LDF6ghGIabgrWC+qrMUJw1Aw0XZOKIvMmWX9yGyV3Ki+ZWrKCC
Q23MsVAQEVYT995+NBuNAfEvyNE0dWbGUljL2lV6NW87V0wkO6vDGKthXLRZAVw4
eE+OW0KyQDQrub0tC1gfoJrsthOp5Hicz6wmfXr4V/Fk53bu9ZNATwNmvUAgSlBD
jXybYHylunD/hhA1qc27GmCCTZBW6YsW/pTXFrw0Aci5Mjxb7or2hbyQFziqnN0f
RuqpYt+y7ZoFN0ua8sjCGnHo3Q4Gyfcvcp16xXk0Er9vER51xlSsnLxRsZQjCF5z
1h074wTftQrlVjvuF4SO/tpCRcgbpBdc5bX07NF/zrl5AfB95WtkzLlzl1/vtXsQ
ke/PuHzyEVKpvcO9z7B9Z8a0dKvE0pvL5UjswEudzIwffvB5hWilmc7VPzWsEKRz
fYq+xDitxdOl6znAnvsRvrjq7yk7sNFUiAhzofDEXix5rbxulWuoz8d85XTIqX9F
h4ifKwiw8/xd4yVGUSfgTm8wpjLk7Om/yl/oLm+v3cCWMpE9HY+D462CozcDujtK
vUl4Pm/JnhidP7KdwcWSEjeFA3QUjtSOAk/JBcAl/OWzKXwuiROvivSHrDC3lK6o
n5bxexQ8wzZX/Ku73tyhfUU0XHw6YJ1uQfaXBwuSEnkU/kHSmnoAcTFEiPjKvLnE
U5TU7qS3p6Qa2xw5uXCBzVb1DCq8kZGKS3Oh0IsulcKqahXg3Q/6WyNIJUaMOejb
ZHPgY2bjICvywgp8B3pTkSnkyTa2AhebUcxRj0cr63opGu+hOCn1H6aP/fRP3Hhh
lp3iogXrLbl+SMO/oSNo4HanyZM5LUP2rBe/1Is/FoXmq/7D6W7n/dOim3Rz7DXM
7TPaXhSJRwFk9D7YvjwWohZl2IbYt4zeNuUGu+W+tayJLNwkM+WG4qWu6Ht4hUD8
7DYV8haCnWGBm67vQBMsxxL2dx8OUZxEX8M4cOvB0MAWUKxiFH6QfIyjEAlEPWUK
Ke2/47ajCdpl6JGh0OjfyP1i2aXVCJ57ZQfbB53eSZ0XQVBjSvUejTHAxSVK5+tr
b0XR+WozboF37wMyylMfmGdgVkfu8I2HfmSxD/kY1G+G3kJyk7JHFavuvUKzskvt
rg+k5POuy3HmlfGhlzZyNx8yp4PZ40yOsDoxGPDHrTQLpL0539qMN9JP2vEtl6QQ
9RwuuggcDE7AlJbZeXPsazKVCTo1OItm0r4+SuX+9cED1e3wFiK8bO95RodbaKUv
roLS8lvFk6qbj2FS3mAzDJII8OTDnkLbgl8mAHkK5I74DDhyC0trMCshOIeSeex5
HgDfiNZWFlt+L5S96FTWZgUZmcvNcHJmmrD1FXqDdOUVl/hw6kaEdPxKIaExoiCW
7VM+aRr64WS9VsRSdA0p1GEPuFZx8YZOf1KZWIjgaLY6qjvE5YQnkLsYtO0EG+v7
+GAgOBtWGPSUm/q9cduNdhVqcOvPlHg71UPpoX6TkUBSXGqjyeI5ocZfDOv+7Vng
ZdkI7C/8hBoljoGhp5+40zcjjN/lSUqXEaKZJfSFpYo8UpBerymz/eAb3oS1yun8
Eu8//RJuYKgUZXkbi7nOHn0YxMZ9jz6BQ5V/EoReU96A6clEh21MIs/ik+ar0LDO
KpaBFLbJstGJcu8i+H0mVLwmQOyIKs3GIlzaKmtUyAMsq3P4+icmX1DNSF7smrlI
kUOXvxNW9PBsMvC1sEhasHugKA7G+MBdZtP+se1DiPDUjr3F2ah3wI8pzDgjhvmw
hDILFs5CKcxuja45RnmznmsGIODdY6wgZ3CbF2h58VxrKR6GlluSmdkssiT4sQlb
ks8TR46BcYZjWCsbS/EwfIu85aelg7oTZYPocJEWBXcibZiHoAp4Jzup99wOHeD2
FIDQlb/Ld8jPYXBVO0x/WIuwY+CDCYe/lEo8Q/pNQHoMFf6HYakpgNjdOuiFRq3x
AxjR2Zs9mnEJdhxTViyB1qFn+5WWqCfnhq4Mv71H98XNDzqiKyjCMexSmzX3KZ8+
fUJ+4hC7kktcy1oM8OqvK51YquHh3CkEA+5ailOBo+Miry7zGaWBBMP6lQgtItvV
i+6daAj1NVAjKQCANi0wStJEwigy0JD7A1oVz+P9QHJN1WDLlQ4lNDJcO+mEamTD
eLNoouIuK6SpfVx0QvI7N/kcTkmOAYQV1oTQ3msVSHRIeUG/aMI7Zi8J66BqMhve
WZn0QvQckM49yzUt0kqCODMDLnYvQsJzjYfQhQL5hzcss35T7lDVrMxaY2l948mD
XIsUaJ8WO5Y0VbdDU+Rbra6ZtDl78PIFMWJmSTcXQ7IzdpZ2Krv+Nzag7ooaWVH0
WxPWYUUVHrJ0LWByEJ8eEOcMApXp2mMN9RQ1UrfW2Vx2bBlC4NxP7iRvz4LF+Noq
V5ZM47U+MDGLlWd/qG5ccI4oT4ZHtHjKi7odXA8fuVnwIGZ8e7UM2+mHq6njzV19
aLtE0IYGWWwyLh+KysjV7FOvw5X2+cPbHHJF6ANRwooGQ+pwCzLRTn22jmav3PTJ
UFkhnqGX8RSjecI0KhXmLjEZB+vJGdD3y5MwzgI7Y2cQmqHgwUiSNgx31QhoEkQW
EkpzIHAeDnRQVfPYQ8ydkZsWz02akohkwsKjVszOn3TiQSBbIP8wrTD1NJn22HdR
N7HDNbtuvyrqBsVw/Sm9HU4OrCgF6j3KvxcyOTmDkULd4dC3nyxfjDhvWalIsyJp
tiBt8vEHwd7H8P9KMwTFIB+/D0Zyu6aNbAD+5S1DZ7QpaL3NXU4uxpHNrQ0NJcQh
xpz8qoWUw8peCJDJwQ3QPRhYP9ULl/v9BTuj+4LqZo6wA3A4xreLTBu2HlD4K1ua
Ba+tWJR11+4gcO+wQ7wtwW5075e2i2Gnt1Oohp+fwxizOe2K9ogi7BHCtyOZAQVe
QUk9zKwme58J0Fyo9HeMC50sZk5iwr+y5S9oCXohK/c9+pY2eZSxJmXFQatJ5ztj
Cz/l98Ul2aA+j9xUppLBFmy64i6TPr2O3VIrIVXfb2mr/H8mvcCx0uLqhJvKWS26
R6y8LOTAQcr9xI1vfdVPoQHVU56CgO2x0NmFFnvEhVTwsOy4FV1vCGhLllKYD8Qm
Rg62IBx5oiiSvPQ1KulsskD6dr8lAwuaW7N3hCZ3ZFZGvJeH++ccKSHtyID4+c5P
8JtADXSbQvhwMKouA3Am27qLZm6P9VJDN0ioDfA49E8wTvm18a/q5NvQf9QmUskL
qGdu9oI6JMPITjLqAucAbp/FmqUswb0dAkzG78wmF1gU+VdSTFfqkibqWRh+Iraf
ksIBK5lDqbWU6LGIOoAoeCAhyWLC8GrSsL+tTznRV95nYa0Wemc4vNh085ykMxwv
mBEMBnGaMfn6HKoE9YfHg/fPzM5+jtyn8tn8PE9i9IsE9jGniO817PGZlNUPSHIk
qpkZvnHCAbs8MmlO6cXz/jZwGhV0JUbpY+vC0yeQ3baPb6QPVMk8dvdeSYyabIEC
0LamsTTbzM5+BBTeW01qBAM/fS2BdekiFtOHAJXilDLrqXVqSmciLYfs7tMVm3Jl
lUhIVA+gSyPQBYVITlfq20E8JKw0iMXiH6TI+skFHX2wWfB+Rcn1n8tZDxIM6s0D
YG1LRfUIokVcHk6bvzHlvUAe9nhVX33vUOLbMhqblE3Ay5KTaMruBM8k6xTpe6Qe
IrtHC970wM3KbMRz8uXS+yCH+Ep2QAb5APmWRjlyKegRSB+y49u1JFlkd6v4z1tC
0qsASTc4UmFQ+NTmXfoXgXvHC4NG9sbdI+R2HNXa17jwH4UstHeTm36vFUxT/04m
+aEBN9J+VNAKiU07ofLx6HwUg4w3h3aZPsSlAsIwofYWEIQ/eX9gqgAnC531FWjJ
8FENAiRWEPcRGXclSymrlOZu0QuxtXFDl3eGwc6LW7MrUUEQ4XAN0UKeYVHtndee
oLX4z3mR8k5f4tO4xcRE1z3qAfJCWHh4X1GXR3ogc7wps77uKGvBz6GTjz7gXJQ4
mQJ6Zd7iI4eQ7kyvJzYyg0dcT03UweNwPTDNFqnKCh7fXKrFeBspYv2xgi7g38s6
ogVzDqorfkUqT21m7Li1guUBzulYbZz0tKF3xXkABUZjCqPkN+H9CSGjnn/QC4gh
sQz8RwwKrcOdPASoqWe4e7p4Q6YWDega8W5qJWp0jVY2CqAJsHIB/30r5wdYKf+k
HonLKrEOu+p0m/3yhQfMyCvIZqe2rITP8N1+8orIldNY/1LNY6LKptQ7X73+LkqT
yF7qCgXpRHIG8ResgGWvSx2Z/PKfZCbRhHwMpznXJ2HZ8XLoyYw/AutLUJmoaPs2
fEtG45ec2IyTESBEwdrwm/AgKy+RchNFPrKtCGNsEEJ/iJbJdBdsznWUq665G3Ce
Ou1svN/ngY+3PcdEHKaQIFfD4+vPfwZrwkT3StgWB6LKk+qozg8eo7hlzHcNJ2rR
AA88inBN4XBVHSuyTtlZfFqfn0uM2Uua9uOBaj03HjsonNiKsDVBiABTLI0XhLly
3lp6dcDgnkXBQXHyJVXKeEwK5DyBTW9mBC28qlcT8TdlALRHc4G9fPokixrZK0UH
GkjnWZSFmAUrodqsxMPVcHJlu1BbyMmA/7ribycjO9YQFaexH4z9FxN0tlI/2X6M
dhu9Rz8mosQ0MkRx/sep0+zWRrICpt2mdKlrqfJVXW05RrZy5O5hQOPDvxrh3sSJ
ysB489eKHzEzAuI9NvYy1CLu+1u6m0Li7uvuWOX1s9KLfSj/VwxxOu2s+CfbDCYt
iaxyrs7yj5sxSV3phgTqZJefxuXPdYFVVEEuXJq51rZpNBCkd+gNmQAd49Xdo1vF
6l6+trVd24KuGH8BKyusyLz9ACdMFXvc1iBClkjmLLNNyF0knq9fg5ch3iHdqV6M
5kmx/GifWd6bOS2LsL1P9n20+PJ4BZF7OtuPaKxqYPCzqay51mMuf6v2MiF3Y8Yu
Fu4WvDwto3FYD+RAIVyODZ0Ls4iNcEKHzUl9Wx/CdguEOYDPVPbg9iMZACX2bI4M
cTYmvy8JUlYT+bbnujSAYKU1VycRHOxx6MbUWh8R2qqiIf8u8EAwC557pqFf89M1
v/IWHhbtnlL2wCkjntqtSBnO+MNTT2pve3+3Q09JXbaKUkHgqeMV5OkA78lnRSNU
TyjZM5yKC0HluI7zbrUgCtGyXeDGSZHYq2fHx9FJI7on6Edry6y0BonYReD7lL1e
s7uNT3zdhpSY8GsAovgUDAyO//1mEJuC1CBXDlbW6PfG2MnVw9zuvOedtTuszbX3
MfecEiNDRRTsZuqcrnfopCEcUya/XkYwZd+T+yFrmRA+NjK0aGJz7nMWKm/aO9p7
VOMs6MlD8+/KrgcWNWnNJJdY1ykXFOH58/bJgj2gD94dcQ/aTecnqDH6ri6CbKj1
n3xXhYJS1/OYOiM6/shtSeNSO/7pzHt45Sj0Hcebu9jNPPfMWbg9GpXTFaEJ0DVQ
0ddOQs6ubP9oSCGuGxhW2Bsv/Ti8Dywk5ZNClNewVFwZA1nxBEAwN80jq54DpWh6
lVnS+prYkke1wUXWrOceDiIFi15dEcH/xxzE44GY4PGZCqnaZ43Hz8X2dckebcZH
QRRfm7BLo9XN7KDUi6jgqj0QvvX76XwpPHnSdHHSBfc1ujgtb6TyMk55RfcZVMMB
1i3N+jh2daNEPqSfVvXuAY73aiSd4bSb1DxVtU/zotmcuGz45+y3c5gF1TDGvXmY
uYQf2Ih3AOX7bh3uO8j1UACAuJsdMSc0hZ9M6cURA+rqQRfhDogpxeR3w2cTtb/r
/GlVZHlRvFiu/6gXgKULVFOrrj91NqfXL7jajPknHT4mrA9YBjtw7Pcho7yr6lkF
E6Tby9AoUKxJdca1KdpEPNONO6XqK6Ac5VYeviDNMkXeBIFMRtZTJsrNQGWmtKqp
ir7tuH3eQt4quJJaJwYeTxYNyEN1MBYSuW9/rmNSulHZ5o1GZbamCgDZnKxLK2pt
2EhPRwEtKTGSEotynsG18vYri2XFZ4kzbFlN8p9nyb/oNXGBxhfeZTo/YQWqs+od
2WzyI3FskS1AVdQgrVuuLJ4KRvD6xuo4g192WjrP5RinJ9IFgbERBNiwOyVg4ipf
/stcxezR6ewu6azBaq/KIUP3sc5oT+OZBXlCPe8yu82+40wE1IderBaS7PNDsikI
Ihac4JwXnFmYRYtlZ/diwEKgFVMM7nJmiALWVzHl553y4c3XkGqKDSg41cBYvDnZ
TLlx8fzewJpUQ9sxJQnfDmAg/ngEipuO/m57GrmrB0uZ0gRCJiqjsOXsJ6/6ATn7
wvOvU3uZ4IY4Bf+QG9gl4j1cJCe7NlNp0QR+eozEsnyB4PNH4L/6wwHKr5UKCVXG
mqrBrHGe6TssY1leBidEhCWgS/QEiWC8tjJeJe7IbB9H00UwEjlhONz2TElkTbJt
p0m1SDB9c/tjrSihQFRW3Q56N68aJGoQQOsmbC0eSb1srnpBGjgqO4Dv1hpvcCTI
Lx/WsOV7TeC6yFsnSLUJcGXOiVZ1lk/6kzRMC1nUfzVyAXn2N2iGe79+MIkFO3IA
8B60frFwjX6JmXvYZHGc7JV8ECiUOJY4OaEwwUGcausAsnyDi7BZiGnu3Onx7TDt
+Z1TjWRiOCNgtZP/BgLSeWm3iIeNWfzOujwgakfVrRdVn1eDjWbvaXKtH23UnPBW
OQc85gEpYC1agvP/gWr+iH9m3C5x72cZSzoJ/FNQmKmmr6WTEZsL3cYa+ZoS88n0
QFsZF+bdPRE9Cs9FaB5JuscObju1j9ZcvfD5bjMcfWN9izUbG5D0djd3oAhS5hWD
nxyaB/Ud52btPMFV6JTnhKc1XUXpY7qQ7fpi0xRil6E5GIRu9kU9Wv9yMWXOaFhH
iD7OBjYk5R3hv6Irm93MZTb4IGGbn+6ObAJAl/GQqwftwdQAI0YWBvbjVej+kLNZ
IVydJKoI1z9o0BEHuG06lsc//lxV08Q/eiQyBnnQ5mW+PHVsd5mdi8AE7RMYZK/C
bvRVG5agQf4XKJ9cvGVtHkDCTtta0bvcOZdyXiPjSU4+L9ulqDFslCxkOzjJt8JH
JiyVI8zxemYUtvZ8r/bq07T9EeW0xYcDVaj2g5XMCh2YQMeheqV8cRgWhgwFwV36
ZgewLdFdCNBcB6frkjT6lCc4opoueeCEpTHaklvLar12/VWwPPrNRbHzEpCn2xhI
/rzzvnkDpVdHROAhGmj1kdH0dIh8/WUs1MadnAJ3+YOeJgg8Wewv3/HhLMWvhbPX
i3ivyA+uXBaYFOB6zyhRKoMy0Kuan+QL2gGwkvEjs81CD3LWy24ihuSPsuRrbwEF
1y+7wuAsmn+YirjIZTwKxlP72YLy7MMC5U6cNA2ymVoxDVAGLjmozkCeZMGVf+x8
BDHIkdKeaLfLBG2IuxZHj+5FvnzY0NLkdkM/rNs331DjqFUGUKgTRXx9ZGK5kO9N
6krOeH9mqBxSu4CJqF7fp1RudPuX88Xx9DLYBVCO5I4CPvCDH/ek1MYAu0QqBRD1
8IcqErDBpbxpFeXnoRADc6H+Lj81hiGY/ESBpXd1KkjLdhKjbuelV9Yb1zrPa4Jl
8pWR9Oog0XyembjYgYdefgK+innf32C9ZGnJte3kjQw7QUOPGT5NuPFYtQT2mUXs
8q4ZI/hLuPn5tCXXo5HQpYzUQpXbA/gnJGkVbY6+1dytDvtD1jlQIISQuFDM1BKZ
MjMg8c2RS0DN7fRSzU019uGvW2u5uyCgw54ANFll06UATfZbGrOK7p1/inDCsEu6
/aVUCq5kXFpFciyE0qKOWQtQW530Dg0MG1mgENJ5lSrMKS+2xHUmCwyg1SIG7Te3
Yce+PYVEXZywXQWyZES4ZrElf9lsEO29YMnnHjePkM2fTHQB2LYbYC3DwAXq7/87
/LAPE20ZiLhS2EyAfoK73cL4yCwh3DYZaPVeEJqDsjM3ilkIr23e3Ibh+nZ8tvZf
i8nWeSsnErQ6Bw2vvojTu7Nv3AKBw8VzGfqcEhaA+5WrkXVwOcYOX8MC51KJqwRY
ShkfxNGLEa/9r2H4Iwr8qhGe8/EltIWbl1MQImytDUr9QpVa2L2aoWjn9egZ/5Ie
uPkSUbL//6hdIAueZm8NE1h77OnZR918Eq6Dv3tuWME2j+2QGyRMDb3ZlEE/JElH
fNC949m3CBzF8s2TB+WHOyt/9hQZ7zkBaGwE9cMqhdjKVwlzGw9FrolsrYKsz2nm
B25Bm6nn9HsqB34bVhFhz2R70rH8v9VoB1s6lEIKUgghiGR4EcSIIP/upCucAj04
aMePoeH4XfzWVPeE9MTyfaPQ+GvMhbGAopSIT5TRj9kL+mMboQotqp2TCuIxnWsn
k39qZuJRpl0cosFRRki2dEFY7o/RTBKZHNaiH1AbWHqApLd5Cm7w5ThzDoqmflay
SKGUf/4OIEc9nAuxdwRwd+GGaxjUU06kIYBr7iYu04dTZdS3wL7755yaxLiXskX1
76uDabisBb+OMpB35HBVQhrpBFsH5pbUc5OgK8uu53551JKsYacbk2CIzcNP43S0
HgvKRfFEk2whQl8bonKNXiuY2zR+XCNOLw05/bFl99PZ4wBDLZQA+5CBxR4NnsnM
hh2GyRpF4sKoh4zEk5lKavGavaONvqED4PhecBz47GpMoOKTaZ0lgoel7dRSJC6C
kRN9sv3iDggTcLbwl9ULuzpqZ3dQuYKc61Wc81++Rn7y6/i6dqYgQAP5TL+jjeIJ
CHi84SNtzkoyWrOBtuRCJy/uONKvnBzmRXQmzaveCubwju4/ZV3QnUVYsR0+Q8Z4
OCEat608eDOQwUz51I4dlOGKF7h5/a4X5K+eVsK4Pt335bQvainY8xH19b3XeFjd
OminjPNATKZ3c6viBr7sEPHedJyqQxEYyqTIielCH4PzUcbugZTFhY+8/ivGnxtW
pgrbWJ/SrGRKFvrdxEOkxPi1Mt8Wqu5OmtL4lidUO5VAlCUOi2mkeCg3rIKXuVrs
ZaT+qXR9FQoCuengMV0YijEn2a5LiuPSBk1vFgJDSY721BP0cl726AspfuIauHpD
gEdt2eyDvnnc2VAiSwcFuGd/FN2agWp+hrH6Dtet0bLDGCzw4j83rQLHqSHeJagk
vz2c82kQWlVC1AmORYC+uwI1vBQfJ98afoK4eVS2GHsEIVBklr4k1wKEZplUzQwG
2tOJTGaP0cuIxTZK32yQKXlz7e7ZK2GxlPDPtJi9AR4emL+EA2oIfuYeYqtu5sf6
x9vBFxlY1N6uMkHBcv9iqKlIOs+rkq76/R+h8+0H8ND7S9OEzsyKS5Xo6LNakBio
KuKgnUgosUVD007Dx9h5vOrNnwSg+2e7Uw1eDYvEUl2jXStks5EP15NdwlEj9O/N
1tiIK1Sgfy/acqZ53BD/VH4awdpVyn7bFPxzcQR5spDnkxQgcyHKuoOv5tu6aT3Y
JAt6OPlovN/nxkBGf46ju5rC0jI9Z97aSREITJPR4vjpdTbwh7odbQn8lzvT6pKY
p43tCDiNc7ey4pLFzadIYgRp10Iipr+kXmbpzVTeZMhIgrQkyTslZ54XlO4MUssq
M3h0clAMyGN1b3Ll41cZSTiI2geYIxjP4ZVXHsNDBLSCh+FxYjIEJFqS+n0c0TcI
j7BpfwyRqK9TSIsfEQ/KcyOWaoGJZ324tyiA7G/Wi8x0S2q1zvbKrdnu5+DyKeZG
8egIwviJ2mVIsjAeJgXEZFZJdS6hzhyTfMoYtv66kbazylpUF/OhD5WqUiPsVA9o
LPGYQEWKUuUK2QB/wZ029dijblI0aCSapn5LrzLmz6aWAOOxg7xANk9qli0F3gxt
mcCsB5z6uHpSpXNpa1lOFr9XVJbqow/AedWLSiNglVhuaKewQZzVSx9W3jnnepJZ
U0+FSpwyPUme1x7buiMUXR9ecEn2R4YtZQK9JG3+0aNCXTejkhzzwLY7Nie3sgK/
wg43I+IE/zUrPaXm6vgQ9/D5rMssJmjKIHJNe8Y9Mhqn8THYKYEOnP9GzI9MURRF
utg9r2c3FVw9e6ohaDacDnXtyYfARDU9hzYiy0I6yiK5bK1BU8uonMfgbfl8k34X
a12woEbnPCVVteRD3UB2dSE04oHj/OU8zNJ76fS0AAReVjxMWndg643IBABNlZw+
quhy+6etbT5C33553Kmzi9jYxRwDR6EhHqQya1bH67o2DVRsDyNufD1hDbc+L5d9
Qeji4zq72i6FYzyoDY2OjjxLsVBNYSDUsGIoQGbqziSTqV68l/9UcrNfClqsh1vz
o1q0wc65/tOhVUPlH8S3eyN+nG6J+P1atMYpeeAB5YrlzEpgjKa2DN44L6oMtaLz
mwCaiqC9+551UrUZTty0fgS9ddpJMas3xkgNfTwNr/yNK0yyu5ublPvYZO6gRMHp
8K4opABCG4k8tg5AZeCqP2rCZD1kYYqLvkQgVbhy6MHI9kgrabx995LDvkc6I61p
2zluUNfvRDTS6CumhTbFoyKESlFDKfOBQzDc6+Xur6ojmaJ0vB6u+6Na7etB+xUw
wQaFUVXTGV9Z0ZHpigFvZdNc1yTilkb1E3zvc4GzG5Fmr/6cJtQfFcKEr+XXIdRm
XTGxItpfWuYS++9+sTPuugHGKuTp9n0cj6DvCY5J1Ap9Uyw18GbNaZpL9vVlbfY+
XMO1QPofQKk6K9X7lz7g5/M2bDiiqSHAOJTC9c8XHz3YLbLMBYPVTd3O7KpwHJxQ
x7ZnG2uoaMhy1n2OTU2YSLxpGL/K/q+WoCFzJMU5DfbQnCbjKhAZLxj7kQipzxTY
sEnle3CACi2JDKOUkDQYc9FMAitZx7X68dwEy3a6nGz6zEbCpTFKSWdvyBbHmqfq
v8eCl0qQnRYtH6+U4F1JiWO1zsUTQpE/rKaFBPm7zEGkeeqMlkacnjZjyj7u1FIP
syJoFNj7qSKsWqPSRjoXSe+8QatepVuWKuyUhb5lM2ipTRYvvgHloljIdr7Do5U0
RduVKw/0nRWW1QC2R6TYt5AnavsE3yAg7Jw29VG88x5ZHOBgK7lw77QEFn68LCwa
NvDh1Z+Xu8+M4C3P9S7I7cUr5r4I6tWLWuuQzqIWAFReNZPCPEq1cRyIX0q4UxHH
lYwQgEAyXGJ0DA8bysBDmb36wUMX4la6M/gSr+VbnD68Y/EC05wjOFdrMJO4fEZt
UUVTJyR0NQh9zL5tjOEff1ydwYy46XFK86JQ0H5PEvciRoW32RXbRRW7siNeGPdb
CZ0BtyypV7hqfao4ZDzBZNiXpMdcWOfkEXueygqVV7Vc/kYpM6BG1u4f2BVjovjB
CF1ZRgeSFaRJy/9FtotjYqPplwBAIGwF06bBBV++4b0bQBUZfc+L4CT2gsjuei5m
7moNghT7idPdfkBcYRdN/5Y5pDOpUKZn9Dk+c6PXDMEs+OzwzUM5KHQeIE71T9lq
OMWc6rvZx7FcF5IWnUhPPFGfL8V4kIDpCOT3HmuPwqjN+M75LqyBHfl7lPCqRCeU
eHICSn04ZMmCqDA3LRsRIzYzPTUkdYJcI3rucCdSfU5cMZxA1DZlUhcRnp+WyHjn
wDwlkcRloXsRUokQV36rp8foPexGP+WjwHoSwLMwKmEjakWSiMgfkn6EBCy9xHiM
tYFZxn8vzwKLLJZHlWjae0L5l600EBsaNfdzr7QZNToiPW9rrxlL2piomsGweVZG
qlJQ2ZEZok4nAZERAecu6GRn+dh9Hh2HkNXHdyLl2+rt5kF+yEmEgkDv9goEt4Sn
5X56PRQ8L/4djUR2p5BGIinqhEyZl0CgT0NAJKoV+D0A/Rqm98BLUFAQUqxnDnLD
opPMD664b+CRbnYASV9+MfAJvp5GpkNaz0hlYUhea73HwzGCDlvpssEEzg1Mp7ME
1rr2VWa6op5hjzBQEL1iOSj1N6zCZPlrcawzx9EwPjSIi6yMALm97MaCGLDNREDq
lsBgjF/v2TGjbHXkQM2CGKt1BpxDBRXTJrLDfLvLA0jp+zQbWYswYeWzG64F0JCI
2dQG3lkyINFD/v/meWHLx+OENBg3IUU5GsX2IlO/65AWtuEJMdS4MOWBvRJcqp8l
qPKkT/G73+NagUXQ2a/meS0h70OCDEcJ20BnXYTA8yVenrI1DFV+aJfLv1TLq2xO
ManubSOtSmTR0oNS9PKsykYkNDOvmNPNcggv0t4iY+swObesQcbt8Lufor48QZ6e
xcDDKpTXuL2jQwsztlq+8QE57hE4h39xxDWVtBFa8Y9arbFEozQm3/dCVgKSl7iG
Jc4+DM6FXYKwRo/rqQDOlfcC1VmPf6HEj8IIgbeFhxuW+qJo4dYz6HR89UD86IMC
SlT7jA0h3ZCngz5MiIYS5pE6b4JElgI01trxBnZb/UKbLft0tJs8mnHTzd9fO9YU
Z3NJ/9ZwwU0xP64f/Qde+8FJSCk5rmI0kZQDS5f8/b1eWASacDxlIcU/fRGY9eDt
lQuCliLtYc4a4/XBgBDqOf/oJ0A4s/iMPX8OexA6qAIym31+sIpifBNwsrd0qzKh
T80tCOM8ivqs2g4G9SH64I8MQJo5YVk3YBW+dufI3TB/zd5j7k2tiShyMGevDpAn
T+xRs+Mwly8j4N26foQUJp/aFewm3WB9M4TPGnup4XqJtzT4sdfqXhCVUCL0+YUj
lcSkBDKxURqPzOe0Cw/tJsOqitXlvc9GQqf0pefQKic9AOYjZNL8k1nzZFVKoziJ
YWPZR2jJ4yw5aAmyQmwXBezPJcXyoN6xlpvYyIhl5s0jYGW62BxCcyLhLP4te4f3
fe97fPUcPH5MSYWdyG9QSXmlgYLtv6Q1utuXE6IENCP+o/wwL7+t6zH3WOFlbUzr
MQEifBLCgJhYFfy9xAigRYsXnjDni2QEJ8uGFA63GhfbC6UdeH6zp9OxrUhAIGoX
XbBTWf3z/ghMSWgC4EfIdbBZIVdx9hlDZyHfaKIlewyNo0nhDD83u2ZB53GWVAUs
TKZjNTmVRGh6ieXUDJ1D8zsyHCGQLGE7oKoHVEBQnCEZJoIOrTJDklvCHSPeyf9P
WLfxa6G873aoi/8JefONB4VV/Qeogd094TFd3RBWf1lSB5IaXevmW5UZE8sMqfkU
hFiJonXKPTiZMVvNaxmGaWBSJVKRue1LZ9A6jG0t12a7dhXk7gehrSbBBVjBXDZu
YUUOzVgkDa6Yf9TIAIVpfQ8hNFJdJlhbTAlM9Q+Cg45E0yDl9bHB3BA209SqZHhW
ZiUhiWeDPKmg8DwS8hS8KoN1jvM2GLRPe2xi/KS5V2mX9Aw8/bqtF96+AoC4qxuz
whEz7cfJIXALDjpsN2JTgYnZyNjLi/LCE5agD73+dmERA2RHnIZntiueJkT7TBv8
FOBxrEinh17bzmCCZQ7MKKPkKJaOArd9SOT1XsXqIDVXLzkc2c73gdcfyz9m913/
KmCaGbxYAOmnLJ9ateViOql9g2EjjfDyWSpAKYsVJ3ZQQqhThvIbpyoSwIIPN/zi
CZz3tgiHTxkvWU0R3puDnflt4nX2sDaZYpnZvkLTYd3Q1wXxunPHc0cgwPSWgDMl
tj7ROW/Zg67eVg5tkI5n2suknT4bs7M0+yvzxHvyt3wFGnbpSVEv/kMZ/uffYQX/
/GWoILg1sFaKYdFqqBNGaWCAn7walUuD80lGXHFhA9hxrMZ7jBJn3Nd+Xv654hd2
fE0U8UNic+poZHIs/ikafzZsHn9nzx1e4gQQQaxrGhImhAUtxuEnB+TJSh8wkdeg
+NAfQyGMScKXlJ3bk+eU6onFNbWF1GZYwRNffX0OWafhMiII0I9K2TijvholaOeM
RpEbpPkb5mWo4J6ZnF4nDW5LgLcjLjM/LSn6zC8JPI6IrcfLpPGEN9u6K1TFaI/o
bC0pVLvroDWGM6VpLAiSNv3s8mv2aw5NCKX/Fey7WrevorIBIKb04FtD/3yzKxpc
VvU+puoSoU4h3n2PIAGDO8sIuyOR5RWb/I+9M+RDUlvI6WRLceT7Aei0jL9odQ+Y
KueqyY4dNQhSrEbM97q0c6eJOaFcUcOu6CqAnr0m8wNi0Azuwdxumsj2BHYg2Wlc
/7Kz+gOb0mrzEsRsN0MocJGkmS0GVi4uFu4l9nd6T6Hzf26Itc0EOvpIuB5JOH0E
QMn7gOc97vLTokBzCK+wYSFY4wHmQjFL+KwE1jjN5vWHO+fSiKS87tHm8q4FGjba
rYycY46uapoXzr7vPe8wkOqFIniVdT94yqFjqBs8j4+3NaYRMeG7PkHFj2XYyUIU
7pWfkXx4ydF6dOpoLzJtL0IiSBJL0rY9w254l4Z1/vnLBoXhdl2RJfvtHeOAL6Fv
CDRc1stk/Da2vz9hQKZTE56sCcw7rFhjM1+Ppry8aMVtwbzUCD6HMbBdV4NdIdK4
+Ick2sq6xRwO83tqDp4rlINys37uVVyu36vyFCH/R/xcxkNxgkz8D8mQCHGnVXhQ
RlIjT7lF9o+hRXjebrszi7ZTj/IJh8vEH1mpHbZLXSn8E5wp8XvoND+DkDqeqtVF
JunlRI7qn5XzjaPYHjHP2OrsObHlCp+1N8U0lCkKRJWKW0EWPmSlRsuWfbZppjbl
zeLLjfbaleoEGu2VZEyQso/diUsXi+hsHAB5z0gXhOF1lPHNwOaFixe9t2IWnvez
WTxRMdRANepNkS3M2Ymg19k8GuvZVVXVy+s8TTc3bDeEl/+jxW8NWzRl5eZ7JGBA
TgAbHzobpw8AVWqZfhom4M3t5hnKLWJT64D0psndmIub9ZPuNAgF5vf4GkyeuvaZ
0mQGJavlrIjbbGcP5UyR9/Fu94uXS1z062A6WoJrwnbTDx3t8xI9ioVVpp9wHDVN
B03+kmgXHkFOVG7l9yFpAy78vKLyQ+EIhK6l46U2STS62sHGLBQRKJuIqUMgFsa+
5+xVzN0djCZqK6hGjE9bLIbA4JR2Oqj0qJ+L1JQeajmLMckpNBMzNcu097fItkeK
ULdAsyhP+af9vTxnSkwvh2dzX3UYPMubyPZsb31yknRMDsLK6emDe81/8pDmroo4
EhChr3BtLqqECZmvv8+yPUM2jpqzpykBor4Vi48KLBX0b3sbrSB9Xr5suzYF2GVT
QapzdytMO3z2altTGp2g4lrefg5jKFpDvRlGoi4RQE29Gw3hQgsNoxbC2sCOCFAO
Z4V4Aa85NrXECV+QYFP6I0qewaDsLSnuraqRwGuizGdYgfgBXoenuyXzkyxeCEwi
IEpoqV+gEITfzMQCWfTcT2pCJ3KvUvTydrSQDXwZPttE7R61yXPKiOCiZ2iArf+8
zEzCqHDpekr4fDvv+Oy5y5+TIhdCLrz2BrLCn9B4YS8grjdPEjv7X/kdXdd1fhhT
OXfewNamrrgEWFX3l31Ep5QRFj3wEBbRvvVt4zM+fwA6IQsYdp/720/zIcPsS8Os
EdR2105mfl7TCyswB1dsL521LC2CXOQAdJxSBgh/nSy9sqBFiosjXZ9d8hVLuCYN
KX/MJ8YVU0lllVEsSEB7Xqoozj0FY2RxZ2j9KQe0SS/Lg01aOKRqquYt2gTYhuvt
2qhBCqAqZMNEd08/DBTwg3c0Ni0nJKQs1pX0aw0i0F1NieHqionuhz3Kw1BnxWGq
RrEEkJj7T0MiiMrhdncUXlj0c7Xu00yiRw0U09zaOZpVk/ooLBrMKETktAVN1GjL
Pa8qThTGEST6Edy9QK3U08iRhSvvv5X7hJP9iBltyxQ2DZ/4w2n9OyTGYmr8DtqW
1Kt4J+u521TR/Psk4VF5EQiaPHJeWovVILhxZRM5B6Plx9SZ7P5eTM7pHQNzu824
yY7dZeyb3UlaNrn3m09/MQODH2hIdYl2+nFu1Nj8hFOCiE9wXm+RCbBxq4goFeTW
zOJBWMdMIzWM4I9i5ljZTj3yQ1MHTaI05OMzXVtsQNI8fhTlfBY+L0dkWoSyW1vz
ly8BmdqPWoCxm/+WVXon2r7VfAxEYVHUgQ1tbVzunJyCcMVC1cZj1bTZvTAYJjtf
Dhun7ixgkFdXDXYWEx4yHehJWcWNr9XpvxKbFzjhJdSNuatjlrTUbDEx1v+P4le7
fKMKSEBqOkXrkfGCWFDaI4jreehvDHH4Mw0O/OWfDVw7zKNS6k11BZr1STQTUO0h
JIwl/vuDSjfcqFq51o3MTan/klarnGb9FFCe8xLppk7vKnKZZwDO14JSiJatVZBW
ZQQ1E/snEfSbkGM1iqK6hHvJ+R6/Xvr6Ii17ItbGWP4mL6cUT9agZtKDrWP8FcIE
3Zm4vmSZPp0q0mdrEznp+XUS6OGhlDLZI5PwQahLOnksE0UQLVOWsCloKpIGGnAa
FOXAshT+x7RQIoNThVWifW6tBWhkP/D4dOffuQshEKNqzwRDZlehHPFfaxfdLO1u
QQTb7OQ4dms/EZ7kzQZ+HHD/zWbMtSV0VoMuToZY++dPqOnnHtp5ZfD0VD+kmqk7
y2Bz3uO6rZ1K+VdxaTz988EyWiOSy/yx7hL1XrC2R8ymJPyTmexQncadqmUYw6H9
PDtlo96drTbPMOd0/BYMtY2vJRTlEzM37lUvtD/MZzckbojuxEBb2xi2O5dN8xcz
/Auz/LKNrY1V7VfyVf4lbdv7gGoxEI+boWxgQskw4TIWerGX7qftHpLwjxOsOvgE
j5XDRsRYJHWXpuXJmVFHw3T5dSx58Ym96YstBc2MygCWZrzkafTukICMvN9ViniB
6+1t6IpX08cRbA1D0T/aobNrKbXTYWnpBTaCpZ7sr9jdoiEvYAb2F5GcbMdFfIkJ
ImRUqLJ/BNP8MxS7oUivyTdv3ezOcP0RBKOq9sxUBHAu4T2nZOaS8QaSUEsT5Ncf
03TtYIf0dh9saJf9OKBeNcSQ4LRZxROevM7dfCeMFLIrxZZuUZAgSUWmiwmhzOwr
p9sveC74CqSUclyhzDCy6Fd7P6SHmzYluRFiRYY7RQi9THI+gxmrcL1ZD1IvZeTW
0OQAf8Lr1fWm495t6GG1dpu8XjNaQmf0vTFYv6SXeQDDow7ULCJuEef7Hzd8OaMu
SmgHM2aPVtH4dzv2ieUFUbf/faS1oSCROpvWVPqNXB9dneZT5nng1jQQ+9GpzdnC
AoEoHvESwVEINYkCm7aUNwvM8dBGJLqqVDwNoqtCYZU9qOMUoSIHtIWrtSgdUiLh
F5AwCHp0ptgE/eFDWIsrjP6pMbVE13VQ6O7uZdBB5hPIpqoEJQS4gUiSLAmsLQen
9kXYjJ6QRENNgXPXxuFq/cRHTuknoFUhOmrTb7xMj5DtOoJbsU4Y97QN22ViilDe
h0AwJQqKI3MaQd6/9AtAHkX4HpEYnTV0VQ9ILMl4hJmM5Asin6PrSoaX03gGgazF
rB7yNoGNbFnljKHIq4TT/OOQQPhjwlDYbDDc6miGVP4vPb6EP5+GN8v7K4xkReTm
0YqDPpNUzdCzRdCHKrsUct4NVgjd13xXFq/wxB4PgHeSiJhdhaKpm8kQXwXMp06u
6GGL62+12fZOqIuje5MuuPNsf/72Su9MzZm90UlsbgFNXWkq+3lkICxNpoDYvZGt
6/pIaqyXEhY42K8CXvd4aT7X4pIF6Oq1h2JUnbGvdR6FbRI51B+RYeJYa9pX+5kk
yUvZMyku+D6M0r+lek3/+ekIA2aGLHux9WGsrAKMX8mUgOiFMCmsP+NfC6KtWGjI
C5nRl+FxhfaHKorxnei8RJf4ucesJrHnM5cRxhTKonI9wvCLYqM19FYjqSKPjguO
tz31Q2mZT8KF0i7mNWePtWstIHpfx0EggqTsL+TX42FE4cdd+nvRvMSq57Cy8bDk
Nc4iFf9ninRzzk1jpvS4hBxZvv0UU9gWDza2k0Y3NEoTRQrvTrbPgOt4jtSysHUr
G5EUqk9JGl/CgJjIGxA0rKudp8lhyS29Dx0If+zUAHoNXhszxzYLv20GnQ7asZIG
Mz51QadcDQoDFqDUkVF4ev3gw+r+CIzTRrq+rEDiY2Bb4VMXKmT1Ycs0tckKIxqe
/91zz9S2+wyRKtXG11N3Yp3erkEdQiinGtCDFivl09Zqp2vI3JJ+5qZPCfp6Rpmv
DYxasj2Z73PyyB46md55kX7oX0IKUsD0BE9fpFNZ4Q4YxHVF98uwwSAEsonrAnxh
caKoWG8jL92fUAMU/mvRSG0uSo+Z7xKhRC0da399XzMT9HmJHngULr72S8PJPHUv
g0dxixk30hRvJ8fWjpiAPJPGPijCkrKXuEdf6GHD5eesMRR9nqFZQoyijpCPcgxR
Vg5mRDDSVkyR5JzusOqPsZ/NQEwaKyDKHiGor6x91lgCRwL+w6sYmEltohtLVh6U
TVm5F6Ckqj9oF4GFz+qiPfidSqcNOTfVsiXuFxXEZo/A46gG1St8v1hap/ZVNhNU
Okmq2rO7eC8qZa78I/fWYgkN5LsOBTjOeZh1hHock8pU4QgcOaVWQF+CjVpxsmMD
9PwWRMaCW3fQ/MyBkkqQw7o46TWJv25ampvWP1TK5oamDd9EnXZ4uGQCEVPk9Qqt
Z7tmOKL6qVSYL1JBsqYsAYIhrW2DK9iM2vjae1Rnc36QVU/qsjp5z2y2CsT+GNXl
AOvVAs+2WWRHmxw2QANbKpaspP67p4cfcGOx7lsGubh6A9sONPZTX620rQuXsvuL
oqUZrOMvJX+eaLth3cmOEpS/igHt2cSl8ZrF4FKyvlevlefBGGL/7ww4SsXW+Ku+
Rep9+pbRm6FElMbn5DKWM7HwLqOfM70j6L+AwVIgba59+MWN6zFpunM8tfPtMnm5
uCBMMghIlAZ0YWz1tP+KVc20ymZ1DE3Z8GJll1b4zADvUZs+bt0+iBV6G8LOoHb0
Im7+aAm/d2KETCrKZyyYHdgsM0Al4IFWut9vxjzL8NCkYKJxsPEegVK2oShTTXvu
lWrHGYDS9kS3PtLqw8dbcuRcycujF8yTrFVU+Mxksu5RBmeOaKXNmVvoArekyaph
JStYR8heNPj7RJ3hNWeTZcN8wHL3HlzTslKaJejzQlCCJrnDkcF1mtLPp6/5cplA
UAf96r36qZSvZk/6JlsCKmi0Y64akXuaeWaXko4Mnj0LJLt7IV9hRanESWOC+6iC
T09Jr1w4PaMk5u88C5HNS3sEVRsijdQF/xXX6fqvs2T7rmpXNCjP0xHdGbnpCFo1
1sLlyzRLOdtMdb3DTqiiJzMD8YFUOX+Wy8a7GPf68btEpgpnxtBHXy0ucbUleE3o
dtFEji76ZlWWlVemt1iNL/BWdk5ijPgs/+aoP1gTNIGyEZ+OSEz3ReO5VrKTEk/5
gBDi4wxyC0dr6ea8d3jX1tELFmZ/U4fEVQEKI80k9QNbWirMHEGiA5sb5qaDWL9J
vjYXalnCJy/vO2B9TNmr/ikUqAES1J2pAa/zSfJiUtouBvhzKdOjmMkrCnsMPyr0
brC8V9cbPc6z/yyDEog0sHUDewlBKH/bvPmQeaCZ+2qQv1G41qG2RUz8jaCi4Zmt
UTbHGa8HINmqZXsveZEzUviy5gsjKgnpQ+q1K5WcZLHxPdMJM2KGn1xkbok6gc5G
wZriwUM4eZvaH5xvuDAVeF1hrQxZlMvI8gJ+4KXMA8bafVxaxS24bZmJZf0GF3TB
WuSJRibLfnHb5K9QKPQ+71LlnR7xFKqsC96bnRVev0INzQseOtMUZ/k9UZ97jyZ1
f0Z1NDh9YVLHVEXcuUomGZZrFe/7UaFHY1vKtsGCghzB+G3l0OGhVjEX8Zmm0Icj
WG+1mM47ji2jR9l89UFq4dbMOq9t4mStJHC8sLACuEWHAXYKrNA62e//NILAB3PA
y30WNE6YaNfUI7pLgrYLM90XIo5AgU/4XEw5sr1qNjZ5sEyopIWJAcHxd23o02K/
UkeLbtPfIi1iA7wOabSSwG/ebxB5Jog1xcRELlqH5bPdVg4BFY3LxMtEKEkvYzdE
jibMnxAIs+OGrUznjP0Et785AgXF6KjXpuVgEXPG5LXZqK5+1lMNjyFFWMKtxnEP
Fsepa/CLGCP3PIElXqU/9clm5guw4ODrhIoSdO+Vu3gbnS6Eyoo7FDyVsV7pRPy3
L6P13EHEpeu3LFg4TsYSMV/s0DFrCHfmUrhmHnwho1GW2oOGAgTsN3uqeNzZV29K
UBKjP3lxkDw2vew5bsewELNq2H1b6lQ2gZ++lWMxPQoRuqzvp0MHaBJ4MzhYv5o4
Wpe2bImldtsYFZ5KGrj2RqUoC27xDnw0FbAfA7PVpGS96O+gWdXJ924RLefP6OmN
zm7EogxVLsTGD0nhhfDBoIB5Tny4l9jjQZxR28nv3FfUt79b/bi39ti8UvMpkaAr
qlngLG+/1qKO5aWeFBUmCVrI+96dQKIbvp7EvpySB/LtbS7y0ihtq2x67FcyHZHO
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
M/Id6n1kscpMYwNzcHO02GXGDumeephJCqUZsMORBt38Qx5SK3mfGb2PpTV0xBWz
ohj2/Dj4sfe7d0N8i+0sSyYowf0vCDBBPO2QDqAEYPEYqAWIMEXxlxo2EefoG1Ha
y7pcx4Jp9TMzhzpA/3/cBoRU/ECoocjvXRNTMUDAhTwU8CFd2NQZ1vICzyCYGyZL
RDGAjI7IvXfN+hbbFcJUo2A9Aw3d0UVqY2r1dwdJNMvoT4zkUFPpODiWOr5J++58
VJWQmMjQ7YfakJ2nZNJMi3uQEcPbARor4eDSgMPzWnKSId/J80G94fUy406xbVWR
Tn2+HRjMPg/KNF/pUg6mvw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10416 )
`pragma protect data_block
rdEXVnjEn3xRKX+mKfsGwDUdigkVHr2zBOC+t/kl9vnYheGkF3Wno1YHX4fYQHhr
zeSvBafH6mfv94a4NPzRezruKa2QkayMhPDzdTXrKY00ICTXtf7usnF/HIoJyAIG
51uSGm8rRk/bRGfjXqRnnfJvlZBJDX41aVqm+j9hpQ86ECXOIO+D3WGsZDFnip/p
+IVLWbd75+fuYXLcjn7lMAeKpU886lZ074V06BgmJECbC+A4k0AIwxaBl42TGGGq
H6SJlH6Kap3Qd6RrwFtf9SZKVxv0/poNPDrI39tEGB4Vn5zWCvSBEhQM1zvINA2P
Uc89ekyL3tPB2Wkg2wRTONny/NOY5DSwzwTMs2HW5iTLa+fZhJPnENe5GKcOUHYX
7JBskjlFbMbXbQskCl4cNOEc7iJwrgyhCMCIjQ9B/qLXWGNY8/fzKu0+XAauVBTu
RjSlfuUAjHUDFocAs5IIPFUQkgfidGbAATh7568v+HP6Oztv3h+Lw0TWAxqzlOF8
dH/GuJU82f+mpqJ7bIqSOfuotbK/OdfaIipoqt7PK/t4MEqfkFY2pVXPLcWKCB/O
XckDOds7MMIncmII7Al35ae1TEuT+PRV5xvlwtCfzJ5JpfaKchbYXwpmzyTcggyh
bEy+EiR1BX7rNBUV/LZSc9vM6WT2a36zMoToAYf+bsWHibDZRDw2S/MSTj6HUlyw
prU7tOuespy9qYJ2pFuuvGq4QOdXLiGMDlvVn9dN2/Sbmg5A2Dq69HvbUi608hg+
NTSKJX7UXUm8yrR/xvWNDFcC2WIHR0yAuRDf2JoTza/Ato2FqzC54C9J+XONu2Wq
XbGpTmhgEvMQ9MV0ormnWz5PLCiMfE3cAANZ3ioWzWmTQoPvZxby3SCz2MfeuJM9
HjkyrL7FC96jzJ0+6BK0Yd5WDRd/Cf/zkwCSCpr8PMVe2V1T3PnKIwTKHGMtFUUh
qxMcRk5r78fdJrPM3xYfMRxpocrD0aDajUXjjApclEgd5hazSsCFtJNJsRZ6+0rI
DjKz14mNaYfL1H4PBS6ANiTaKJUAnBnKxf/GomIeqex8gRNYi8Z3QYamyxd6gsOU
22AKWbLzeUYA6807v0GaIzKRiZnNEK0/uxCSVAKV8LaEnOXG/nrbn4d/CmzZS72Q
/QSbF5REl3FhwxoA3hDMV0SeevRGd8mQnWasXJ0MkysOr/1r8ASmJU4frv/Yh3+U
HxUURVjRoa+a1p7LvvDYiLYY3JNypIGE9d2ZOJyQ5+NAeUfL4oJscvaT4AsrUWEC
87lXT2dwPKMyIJu4ydZ9LgQvit8O1m8KF8az85x9+wDZWhKc51tjuAIpf7qzGPS/
cwnuv9yWjAayqL+ZD+4FpOjID5V8MMsANvFDEMV/gOrit/wvqFdQ1bR4RPga8znL
UU+2h/xEPf0xw1HK9qTI3wGY4ptFqyc9RB1kAHP7H7PtQKwVSn/5cnq6s3ForMgk
FTY80Fo6PYDxmqfqL3zB/qO33rytaU2m1QoX41hjAxYxK2zKGrZVQ0JT0PzO4bqJ
R991/2qxXEqse3roVccdBUIlmn0a+4SyA8uvktE38sv8vvFWIj24j8TDo5YxrYCW
RoNF2/JD5hlUYFTIYyUBjrGxwHCBq+1RGeQZ3Jvi+/CYDE+u6P5xNKnoSHczFq51
N067kMERLHS+p+5IMFwUpXcOyNv+FVTthCyci2oA08PnivssduPff58NrQYPSp2+
EFyv5G0sU37ZifglXRdlIqt7XLeGxaFGVZnVuSUzFipONtdlyYV8rMNck8HoDQya
imRmTH/inp74UPIxwWBLVXcPJTRqmV8y0SKm44ZtFBmUiA34HsnUWQT0LFWnQxdd
bsh+jvNM39texd5/FkJmUFRZ9MYMCCgV5NBpjPjbAUV9NFdn6EJ+9juLDTsI6Oo8
uuZ4+yetcALf7CruYK8zXKt6pg1YVghf0T8v7QHp78y4dqZQukCWlvXXst0e9QcW
HpNoT7b65iG0fUwCQqKfRc+4L8gCp3hz4TQ6ELdKLqnpiiKaVXcBrfT38jpLQSMC
U0Ay/Yi5ijVXwsKBRhvN8QWwqfG5heqocrAE4WW/6wVGT9oMS1CO9NM3B8UEv4Ry
xKFpRHiZQ8OC8qtPQ+LopkiNJWTZtsmmtz+fTnbeZJSJCKA603laZf6M8aRcMRBH
l8Cajo6dBhrCivW4+T9GDmTKqBsXQ1LCMhrae0zkpQoj2zn1loQisCumGjQ6tTF5
gGnj4zAUqjoGWa/QNnIKoj416thTeUnkdj6pwPLjP1P06DcxAJWT7FhTn/xHqwSw
8wDYc4j6qiLRSfVqBp/3p3RqTLkI0CvTrI+WteoVJmNG9LeMilW3JkNPgom6jQEo
F9vT9qLDbHA741BJQwKoAbQYGN5uD5OptI5iufT74GdbEMfzAOJFTFGKhp1PNqfT
3Sm8alliYAXU06OqF8aBDKr4ZgCyB1BIL4sBePVmCDMGdgI62z+VqBcBVQeIIi00
qn5fmSitpZabXPAb9nlN/DcnJKXLxLovQhv0Ay/YcO6Hv/NqjnE96fwAttv43Odo
5KPHfmg7bqeUDwDH61uJ0zWH2mvmEVAvaWjlVlcHVVCR+V0eRiwSypdV3kRsh949
2wNShRKqd25SZmnwnIlVPnTauxgycKJbHmqBLzu4MUYFfoo7IryllqnF8g6A0j/D
pHHGklODou/R8fRZs3lg/3UVT6jw8VmtjOOGxondkG/UiFx+Ka/Tu4x9AOGw+Ps2
9lE72jj0DOub4AQqbCpSNXejB2N3TZzkDpPyfES/5gecT5LMZb+jJ6z3o6N8mFf7
MBUUGE2sAWg0AXTbbhzU9KXdQ+re2iYc7sze8IWrv4qgLCDzk+d/fuC7o/yHgTgG
8d9UG8RZCatyWfN+FvbPJGxR+NVAue7cl/U92H58zia5t/m7uR8obJxYU0TLtl7D
APhM8rPZfRxZRTePk8bfZP1oEjVivTpsKOR6HKdv7fJMT0YXAfTsS68fp45EP+uy
o8fkWVQH0w5T+apPy2t+/ixNtqfT/QcuqelE+CmpUeg7KL6+4gvcC/TxYq24BI8t
yi1T4ERNPI4zHJ5m84ze9/GjB0UrP8pVEwKjtaFN2BaZsLb/YFRDhIVGUivtsq8G
2h4t2RmGyR1Yd9XI4CQ6lD3niEYWtPXKphLbglKVPAqd/8km0KuThDJoAc1HFskC
vTxSVtZpFz2EUTEsbZAjosP4m/kvO4HXNm9EvCYXZp9RXIwEDXo8PMLRlgt0t3+n
k2YsoBhQsaYTIqNYSektTO3OuPsQWEgO4uP2Hf6idwB39Jf9gCU3mtQyWrlIjttX
3dHruYyXDB0di/TvAxQp59l/g8M+ZLy5SK5C/8tqM4q/L5MDrHZTU5vyhFVhUrlq
rfMYWieIdhIg7bN6mHf3CMJIV7Jsz+wpKFAc6CfCN1agbC5B4Vb+q1j4HvPa9zWY
D9/mqhFEIoy/7EQzrO6mW/qSpEbQ/GKC9ZuyOy6vnNPufZchmx8sAQ9Hsct7jGBr
1u8Ux+yMtHaaXpQhFUQgp/TRisNxdabuyFi8IgwyjJWdnvRIOvXWAQE3V1KliInX
IkkoPjyeuW5VGbj4C39+FKSCU1iBKrkR/s/W5yV0zeDa3PQpVYualHpTwXOR2W/Y
bOOld4m3L9PppXK+FzfoyxHcDFlX2w5JBapjrNRlBOy9g3i42jC4nZEkskkbXI+F
sE8vFsCMmqcWHPsEgNCbHVp7JZY7tK0G79+sNDnW5dMjs10ePRxK9z95NmJLNFGh
9dOSUFwHuZzMwFpcqDNXkBrx+GEMapUiop1zXVRudgDbuEYFqxODJBda4csFHIsb
KZiTw+M0b/Q1Y8b6nZEzwdaj5JHYbtSOloJ5PZ50nHE5mueNBl8FaHxSKXRbnEM/
2U5+Q98/WAO4HgBTkyodfiFj3caBf7Jtpy6OhvZHLM0ZZy4qZCxrGkkE0SAaIaoP
832bs7dbMLn7aOQ8oOjsaN7R4zSYjKpEICJLFJ5OWnwYH2MPcCU7o1NqtverBWZo
QmZlfoJSmq5kCywqDfxNm9n75R2kQIzHd/RLQhCr+I/+PRBVEPk5FiriS5bQ1gcl
2pz8IoX7YmeW+mMMFkLn08JWeoUeVnBZyQuAj+1IE7cwBIpZlX7kyc/x8WSMK5QA
qz0GDGsl4XEFMJJtmCqge6rL8HYKDxZzuggIvYJ+bYg0rLF8GG0M8xC/7PsByQSz
78Zgrrb4so5vDlChFekSt0KcGCHyXMGAOAkM9d3J3NIumZvCanLvAeY1Z1/cDcrA
9ALboF2cwBZ4Rdn2tR8dMmBSuAg8cHlD50wFoUFNHVsOR+8H2Ugyjf7Xla3+/VBR
kXYM7cBVkjBFlxE9HsA30q60Msa3PgdIPdnqCSNECzCzsBP7xedkybFuZFLAWtpz
o010jWH9uKJiEImk5uKFCEb2f76/KYr6Unj8mMfYS1nukKR/FWiyjbhqBDSNr5KG
LHtRw3pRm2MRoDX4RV+obUJGPu7e36nIFy4/NXNBlxKzj7CUDSrWI0Bq162IX0Px
vZPiUfAuy2hNfjZIKtWhJ9nLxvPIfrDueXF+M37/ETLasBRkAbudVIoGduwpdzwe
0Tn81WxcLJYhPvowUDwv0FFPU0QecZ1oQ8pekhhaTGZL9G/Yv9gEvnkuReSukfrn
F61v8CklnnZE1JbQtqyYwWCnuaVWwBMX6EQq9QGUNFRy9c69nvR0ZHxwoiURZDfP
PpoMs34Pd4pSSQpU2/FOtZUXySweV1ZiSaEOqpSYeON2EzPZtiGy10AAEybEizwn
B74tHpm+8n3cVg5AsZekzGgkyhs0v4Z2PLII7tce8SMPF+/8pMfCIx4+pTfcThPj
/CMxn80/FeeDkwMMaY3rOLCoSZXsWOoxVO09nDMS03A3mAJjDVFV1Hssldh1RfTz
5rdjh6/o4QqCHXTy36u6ZWkJeyqFo0PIoVPIWYeasI+w8sLg1GiU/cPxK0CJOQQ7
4mLI9YmYUSxUta5fywmUkp7ou9KFEGzwpNe820KcnbzRXCN7TI8riY9T5nsMal80
zOpiqs1oAYWLW5IzzowPqjtkpC5E4koV7o3QTkpkuBatHOp59eE7TBzpvG7/m+3V
NBIkhaKAbtE4H02uYUVTRdviUq2M6PjG7qykkKYu8IX8oHEjP7U6UiP5UiRzYUDT
plMG0FdhFJYyBx4SC7nlCCO0krD6I95LE/FccMu7ksmdxv4w7rsUGr/GsWfvIXZb
kZp34+BC7SKY0SjPMx2OCElaREdWgWbWYn2DQkWbPyKypLH+Ve5Bb5GBt8xooqnD
kXFKFXW1oezEmYnVz/QooIiA9qi+PDl9iTsuV1h4IQPNiVvHF6U617vIndjYcIs5
dwNxG6xN3Yt6KkMJtFlUC7o84gVfXf6fKcaI22JHPf113xCPO5wSt/BUTz7aUBCw
oBe+pEdT5We0xyaqB/LSGBwzxf1zDsnuBeRwnFL9W/g9Ulej9IstQBuVrBLlqNpA
Vhw5pdKbvfIXSdIr4DR/iF7xfECVhk13CzIHdr+y71D3k9E155yhjBSwkW41QhEj
ZsR9INnVCqorwzkLhw+IxMpmE8LBiNAjlU1Tgaqqlg5G9+Ys6lMUUAMd+todeKut
w3w46pMRkrvlNnvVDNYPGX5Cvm8xJ9vI6BN/asS7fHq0AGud1S7GFmSjLeQOBMRs
2OE06OdSwY2fyOisHzCD05+Yh7Kr7idct35PU2R6/OQCX8Dc+3VO7/vajpEVWX65
buvbnpD40iN9v4MgroHPzOor8x2BscETs+D2JpTAmmbMIlX6fGwr6xP+qk3tANaD
qXmA9NRZ3jefPorsJo4bd8Dtq0WoAERFopO6w/8FSvpX9akEEmLbctDFj0cDnbgl
LCqwhSb5RdGUL6f9fM3Jey3OKgsaKGJn8kOZ/5Y7i6Ww22hGhfZVMDkBCVwkY/u6
JiEz8xh0x54LVSMTy8THnrGK9imojLcpnWcx41FezE9vldx5vkj+PlI9syqzXPZe
U9U3+lH/pQvsiCMa779iVJFbsdxDpKVm8bfS44TIrvbN5SfS8s7RE7A+LAmAP+sw
OvD1f4+8z1XfRYMAeTDBQwQni1QCbum9e7U7hobeW8WH5bLKR2ngRqS3DTDrFYUv
o1Ya/uG+5Z0FsSLHdZFoLI5QiUnNlsAyfufotrJqjdWLUSmJTV/X8Y6iPVfTm48g
gq1A5gdz/Krfps/7ubMiK59jL/wBLE+7zK9/sEVu+jnjlvzuXQkIAhjxhjmCgLuB
jHflRVMzadgeLTl6nirm7xekZQuHdm/RihBB5+hVBt6VTFWT3I/QtvAWpqcb5P1V
usEgiU3cc8c+k5F9CbzfWp3ysgm5+qNgOISJWHsbMBw7bj9eo8k8cRyEoCdTscAU
mJ7O90ucoiPK3nEFGynUG2A42vgxwz/HLlZwcddf5YnUd+tDYHRnZUKUfThlfjzf
skFl0khgwmgsSd4SwD+P9c2WpzwpYr0STDog/a6YrnyoitJzYiuJDetsTRFu/Xh5
7ZnmHfVCvb0HO4k/OPVOjL9nfJNDS5n+NnWUZsiDWJS0Xtx96BhqKSpEhmrzRKMT
Pmv2b5BOdAxTnlmVIuCu1KPGRjbqgvx94+25LEE8GTORw74h+zx3e79mlHUWQQhj
qoSbwdqYeU0VdFdtkjb5aoYK4cFzc3wzSKO0VyUU4RkFtiSm2AXd5aufugCIm8py
HQ9fgYtdcFExqg4eLzXI/QZYkbpVyiumfRsOLNuAPSMsucRts0mW9DO7WS/73P6B
hr0i2kfyszV7UAy9tcohIIhkb9ngvweOl58XCpPWY2XQwn4pkC0a3l92Y6PmySJw
6X12Ca2WHrYmD4vFr9qOknxbnVJ/Rp2StDxX7KRd0nTn9+26roLtLEBqDvBDVsra
NlNivAaI+UcxVhtKXj1gXiGUDswOyI76shd5Oa9G9aLmarX3Pp3AChowve/TnOf2
T99r9T9z/H1m8kkWEOp0hjhvEAQxcbmpht+Y3xKHNTKWa0YKQcnKwtFVFyeHW3RM
eijSHdITE+Z+HhDGPvE+pkg7NVm8Kwi3zaPp+OypRIWUSvk4ylRcZq6/Oc5eIcf2
rN4BnVDuXiY/bQCtAu3t6W6Xq3PSxzQH7f/sghdup1kd+197rQXjAO1Byve+vQ84
LpSolzkR/xFqxdAWUZSgaS/rL+/HjSMeTs8p8ECD4c7GtJT67X0tFixGXCw+3eEi
Bpy6jnO8H10wXIeXE2zjIJtoBFjVUpQ7p3GJ9DqdSu2JtvqGL6XvapxhrWLCi0d+
qMmSdy0btis97mow9c0X9sDOUfRbT5wjJ8TIxJ/YCRgiMvTnrSNoGqxhSDmyX6pc
sl0i3lLATcjVcebpFAS/lNYdzDT+vv+6cI+1y3xPyIhW/XtozWgaNoVl/IVflyL2
h57JRZ/rtRypIrnkfQltXGalfm+MAxVHH/1Mg8xQeJXHjm721ZA1XMi4Xm8tiY+P
fiLnRYyUYI98LldFMfY1BVZR9xMxz6zkDDoPU5/1JhRo3klTwGr+HlX8RtcjgGA9
yuSNJTBe3QqBIhjKTxngAlvqkt1YFQB3DcWCmxs7qmCYcyor4sv+WPw/xFvqyaZB
lKn13Xv/OxYHy0gsPw0HXAy+Yq6wXV53/pdmUHy9A3akjzd+RkR92DnCukx8joos
WNoKfKYmaI/N7euKcOzuGtOFCvdNLwQgIafLWg5Zew/P2zURlOy0dbDk1j0bErRo
Do2mzp9yTmFuEs0fwcb6LZV8wyJaDOlb8qxTJ9O7S2g0WBF028N9yFlSWTQ3hsps
36BBxeGYQC+faUkXTDzQmuZvuIoL7Tt9tSjCU2gG4lWyqKk6ZLFtfg/RtHxFtEy/
MObGN25GpS3uu5Gx9ivkRWtA91mfeYaA+Bs+WMVpXsqIoHczNXahY+iQNbdm9+EW
p2mSXY/jvLK6vVyomqrsl7nc94YUHTOvzy2d4K5Zlg0hJVKUqP8tWbre9jp71iKW
Vffe9rpEG+yilD2bgqYqr+H9+02Jf+ZPufqn/E7XnlR66wvi2Zupd094Bgq8vHNo
12TBRcfnjKnKG6DV26Fn+MH6HtHkMBqhg0n/rlpSjklbz0MWCqKuKtc4MjR2VcWG
DtzGQWkHMYeNvs3ADqTvlF4bB0Bc6ctBfDNAFc0DyvDoorJTWkNbd/qtOEAbNbPD
zsCLtbC1nZ2oXS+8W0DZFJuQKIhwEoW50ze9SkTrWofdHlvf1xxU+k0QmZxkFcIi
MXJVcWjT0ZT4A4hZHJ6s4u+cIpLLFM9qBr3sxdKqt139gfgyBwYnYDXGJpbau9AU
05PUA99G/FfjXrKGO1Ey1oTwh2TCaz+adc/BqBJ72lC8SCUkStro8NukV2cJ5rbv
KbS03hlFYeGSOzxUJOncaRP5U0K2N3LHs2s+k+O++THq3nEYFrmAZa/RPJqsShn9
zGmNNqnG05IdxQH7/iSAU6cLJXBjEPfQjcpuXIFhPwYkzffuB62ireI2Nu0euz4u
Uz1VB4ICwfEB/ZN+CUOUH9riDxXSMhwn+KdBz8XR76BAfRW+adF6jUCJPQMCpVZ+
gB4kFz+cMwNhAhJ5WTghqx/ZmyLUClhjUZrab2MBENFFjbDwl4LjoqL9SK51KadO
ZphzNszcvbVt4AiGFIykEG90EUojQm/+nerBdx5Qad8oCjhk07wWIyhHws0GEeGb
RiXMXmPqBOOeDCt1SyhuZdI2bpOTheejDANY6tvyOQARZz5/pzrH56n0EPKHAG0a
WX7WujuHg6AA+c8iobaA6q7mL+bDWsXqjTdCqb+iRavtNHt86L3Jhfzwy5lt8bUl
Y/u0MAQwa1v0AF/8qaT4UmafKTqA4P/SLBSHj9jFXwU/arDImgKVWjsBQNk1d4y3
MHgOhEXoXiArdfuYeRo1ZVTCM1+1ZVFAkS3yVgf8etyvHMhiFzMUg+XZaZbyMa5u
ftWc+34p8KX+F4ELdGQzdB38rN8W+TjuW7xah1OqYTKrtQXGl5IuUiPCi4Du6DMj
0fvMhmON9tq6eWRjZg0D5+FzDwBCR/cuUl83sYHvLv+gs/atKXklvDMe/W5/fYod
kn5uqGCUm/IgfuSbNkXRGOn+YCt+SeJRjR2kxj3tQyVyWUXLD/+xL3CQSo4tUMyP
mTFviOGXfGf1456R4pVbT8+2e0uo+jXXExG1akTSvA4b8A56V7IJx900bx+6xArd
PIgya5isSztuCVmsWrI+z16g+PlTtvn+4Wcsz7jcwLR+ZlLGw+zY6mZAR8mFqKzu
YgCDCD5S+5mnLKOhY1bohDTIjEjrL3cYOzKsH+A/7ZftuWtVeT4NdD8jChfYc8hi
n6UMF/qNHAAUF1rLfMkyoxYU+mfW2d0lV1z1RdpkLIShquchhX1W9jExMLF+9MjL
gzilAsWNw12BHfc5+FpTtAVUKzXEudq9F+abCUC3tvsAkoMeq3AoKFJw5vdQst1r
Ut6YwgivMKUgL9fgfT1jc53lfJt/DVLLCi7Jaow8guKkzfVKFUddQMAumZJGtPpI
OnEuBZvinq16V92pBOp3LFQZMByuVIXxYPSKiPTKQJs9Xh+FKvGLanciwcoaL2Bv
iTVRJ1aPRNa3O7rOh6Li8yw9iwqkVT7kquQlQvamamjUCngT1T4FDd+gKN0OPxS4
5mHQylrv4gIXDdb6xM/XlmvyL+GjtA0Pp62dCfdp0Zf3M09pU8qYBwW23Q5sO6jT
AB+e51+tq7JT3jEb/0Hchb3uvAZmoHPL4u2uKyb57VaO/mJCTBJBXnc9zLzpAuU+
K4Rb38DxQCkymJoR9H0hAyXv8XmJc0wCog2mUuJnur1emrkMIyuDpnEL/1q5VEUv
8VgA4HcwWksLrs8tAYJrEZzS3SytzDwmwSZ/G1mP4H1mjxo/197AAlWVwesJAGO3
NkUHStoYgTbKtnQJxXFzdFqBt4TMzYiwne+zsKtFB5BHqDwUQb99blNzDCcA6PdY
HxXfjmeRIHZiVX8RO/942rtcE1JyjCT6+tqZsrRWAOinkVzfw1Ku7NnChCwPWEaB
Xzhge39htpbD8cd3tTycIagQqPrJqV7j45VVeuOfODyy23Wak79Ws7yRkvjqF5Pz
VJOiuTJaicuLY1EY9VXrhjvM6K364/vGla+3GE+iedzeHx4CAg5YLpChv18r28Ht
ebqSV51G+VyFZ8pmw7iw64nlvCklUqqA0NRZ+25bYHNpMNEyA4KT/ehjOGVzrlLP
2oq9qM+Z65uJCLIbVCi+L9pCw4vm/pHlTIvrRtJb5I9PUVNXUzUY9pfNoLOjjE+h
eTUqSfVoxGj40lCeFONWowgw/n28Rh/rY7X+lylWlq73RHSRnRFG2Bfym/EzciVk
qiiPRZw/pPLqXL1MUguMLT3vqaQ2M7lw1W0HMysx9qAj0ZpBGCrAyNYGXGg+Y2sV
FIMCZlZaFvuiJKnIpW0S1hyClP48tFIpwtgyZeGccG0k9lISbM1biK4UIk2jXeM3
Ow0M++91TlqiHnwQQxXjIUGdRUXvCrHpxSMQ84RPcbumrYt5wcEbdYCkDlq+eSBK
37YgcAZnBIprUoz29uep++SeCh0NAWIZjcAqZFSxhv8oWBu9fpVGEtm2Vm2+/scN
EFqy0uBKABkc/ScZ2Q0xn3+UFA5N3W7IE4VrjC7ae9BvkZVSGTUbnDhu1vNCty4X
RxzvmNXSL7dN9HLSOb8ybk6Zx0SKdY+/Mq8PLj7CNrZ28qTFRwkL/NS0+WhTqtUI
ER1kIXzeFD4FAPbWeXhsqMZdnNeuVWqfJ5aamLRIytPu0Grt6h3qMe17MP1JS3Ko
64rp60gv92NAx6/baGWKELFBj9avYGJ2CSebhbrkc9W5oDwnxyc3doCY8yuiTAZc
D715t4xj6QhHWbs5n0O/hn+s7w7zv8g6RbgA3ppftP5HndTZA1JaJoPnfFiJ0pDB
YT/KHH2zkLXTxXc9/N2E/016vwUiWL9MIn/LIciwk8gFrQLX0L3M++xVgvH2h/8n
QMvCWMet5/KsqvJ+qWmRvNuhI7e8xV9rDudYD92GNy8vcKzc95s7+YkAqrL3GSBh
n7T2OX53W03J/vOGcLuhSa5sw2OyQkbO1lkZ9+7vK4RlDR0PkuwWOuzSh5dTeIKC
RAMnmkAsJkRKl+BiPmdO9m+sypkZxeO8iBssr0yN7oIr0d+xP+YLM0HHyCBLZaZH
wsvX/ixqh+poF+BabkADHgTMMElo4cALX5Xe7qyeucFHPgbhKcVImy+ZcgGVl48r
Lk+XU4AyTrqNaB89wdsCAcQhXE4whmBewZS4ADOeylM80yvia9B9Ktn2oBWYK73G
yROa5qHu3Y6Pf1wYUorKmOLjllGywWiDG3wi1Sjg/mJEHxZnD6z77dM6meSxg2ve
Wvecfbx29LEX8XnVO5aeOdZ8vXBsozF3CJaYlqIkqobAf2KmqMjCF2cBw83139jY
4N9u//+vyWI7m2Got9ogKJH/km2v1KKGTTvBqomTLTkZQGkQJatV0gGo/L+dNOoj
csXXBh1zKZpPn1vNsfJRjrmB+KIk5oMtLN/E6Ui4KgVhnkDtaGvWyneqGMl0WRsF
w3RVgzk37jJsDIi6uIiW0YWE9Rq5/Zj4sqwXpxmCkGkqLItqDUMr6gVAK/XFkUDn
ewHSVjs4yqr4vYdVVIgoWcud/nXmNx+7NkuLoA9zsJWJE0e+zc+r7PdAcG+dhqTW
iGs0lnkR+He6eO9jIhzMOs3iQaQSlHbnYfyFY1McpN4G5Ht3dQHKST/XO+vn7EN2
PR1c+PvJqancf8Ge25Iokky9sepuglMznCrXX8tI4w+NzmCyMZ6znzAnHuTYUbXf
OplLv5l06H7MWjgRuvUOtcoRTmFV+CR3QN61IgTrvCQG0P5PA6AqNuF0XIAByaR9
mMb9As2vJ2Y7g6Yw5OSxzGpxmC/FWarqnfORlyE+/+PHjuQfBFaxYnfI77h+85Xv
Usvpj59oXeK5B6mM+fTA2cauSTUq8tz4rZl2FCoE/ZGBAaMeALQFK0y53MlXjZfi
x4TpLckk8rBPCUEAn8eVPJVJUS+BBRtrvyYwmDvYz9trXzvYVjbpd18yN6dKlTaj
/yxerLo7gSspP46dgPtVrLXeKs3t6t7bdq0u1BVGqezrrfC1NzewsACNruL8U0LF
kNz7R+CxT+L1pw2Y+yDaPEz8t6MLXDqjWWCTWMQxLQHc9Cnq/BI641wOQ0BNkw51
g5/8ONw7+W4iG/3DAJMOMFf/UlgZrxKgKGYFBCuV98BU7hf4gvUVlwEzcH0ZLGtA
OO2JnYtTR05/oWuteJJrpjQ4Sz5gCmlQBoMMbr7i4dTzr+2ZEu/tBwKb9qnUdYRe
ZUinZkB/Q2xpM4bVQsL/fh6P2N6e5S7ltTKRgsX1OarbaGq/J92+KxLd/cRAXycA
gdMVe2xQwlQXGcb9ebUQXh2x8p7Zv0+ZRSNj4kaNr7IfOWC76Qcy5QxLpcuq0OHp
wlv9trHcAA5mNpMPVLazzQ9UKYDA+Wl6+xWjh4PomVsGSAU978rct/x/DTypOtKM
753FYmv+hWYo/5QfEDxRukOoLo5gZsZx3cRulIWp3zOLigvr/VplQruU8WZr9H+1
02wIYy36qd0IOoPs+MKUInMIUNmZOiW448fsmaewMcwPdfN6lhgSSZp/cCXyDNda
zFS4PPpBH1xzet0rj/b8OzUWbc3ngT1oyaC8CPQa4aRO2jWk1TWY5FQsWg6K0mgD
9/nsNclF1r8F26ft+MUiu09nJBvfruX6pc6pOKjoVoto4hZyeKHhnX7BI9djND7e
FOm8ibQKwwn7pWL3whvGbBGZOjrvJreItPWlwzd4zEjwC/bA6Fki9oQ0k34dOdT9
abmFZDG8W7+2oQ2L2FIMaM4ANbZha5yVqL8kkr4x+WrpAKZIE2cWjXMFwfrsvw5h
lJ/B/Ys2YMzEwxNWdCaYWEEBKDpXGJiZzmeXCq09iEySddiW19Wm0Fix5sdg9k/F
w2aTd8ob6UGt6k51315NAc3Yoo0rScXXtx+wTMRTWhFol2kNGoqvfbu8+N22X9HT
GtfAUSDsgqZIrEGf0YIw04+odiUcili/aN/jdufE1gaU/SCTSq/aVAMLZh4mFpDC
vxFZMYyTzU5vO29+Nnme10IqNao0HBvbLqDjyMSDBA+OI4S2IaA/bCcgvW2ee6JK
hcsSVsdQFag+QTPODVLNjFcaUZ9lqEvYksH8+SdsIpuG5Eo8C/XUkeYPjyMHP1I0
48YuyqoHXZauMT15doQIdQ5E5/gZvD91lO0r97mN4qPLmayklkQepFGKIVh4OyEv
Frl98KjRsDVn0joJB96gNZT/JFUpFMiG+G48U6/RItkxrxWfBWHO1QhO/8/VwCDP
yxDae9RhTM3NpVPkacIdVZNikDIutkEHFZSgYVgeI+EKRq/ah7sxilAM7/86Gs/S
BjW53CnrLfMVw/Wo8itIQ6j50/efFUiHQdrsl+jLeMXoxHI38AsMU6f4dJoIDmMT
wDWoqcpuFo34Yn1FL5HVscnJ8i8tXdJStd3AOTW7ccTyHQ6rO+qclWOoJ5Vxnw6R
Lorz4e1pX0fT84SoT/gBBq2Ela/AFi3eQRnZq2gw4VnPW+8whcBWYDemDyqH9LND
35/Jur0+ITpSWpIOfRRmUQBshUOjYcPP0o/Mu9AiRktQm57JVNO0pntIohWfWXjQ
7sLIwVOrGV0sTQPqk3YAO354wGQOZgAhzu6bnLVJ33hqNb1uhgSvJLmZZ+VsDOOh
SyTgM6Loj7wVWLgzjf0sWTMHWWwYaSZj/tHi8eaqanwjlknmlGfB/55N/6JLYbqP
5siy6FgbXWefxQKz6QGPmJN4KyT89DSx8sn+xQv+6Qjq5ZpgpmbhhCDVY4VGSTxc
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
PFlN6sNE0pKT68cjUjEGYuXacqDf3BrE4qkAt3GvLEJRgJ0mLqjeBMnXW6lhmeKn
BZ2pe+/qVTWXN4JvCatdfiAANQgd6edMUN5eTRVp8rz4OhkMrSk+g0EjFRQ+nLi8
c3Tv1rbvUTq3AtTbnOO0iz2r63Pb0Y7WK2vdkQFfKF+ovjLET2yf/B47pNlKxt2a
KI5lLWNe2Bse7irWdqj3Lcr5j3tdyJ5AhpRFC8hNGcuiZrbr0iu7Be5OCuBFSYIT
yTgZIM+SihpzlxCV/LjpkwwR8DWvosOSpnuXuABK7Yc0fAP5Nx04JwmUBeKfqOqP
7eo00o2A/JJnMptYPWYxng==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
f9RJKQDte60j7ImCEWn7OZyVww6Imu+8USdFYHsIycJuZ26lqsab1jX4i8g6i52Z
BDrpaiwOSnBmLdAblloUoQzFcuEJRxC72yclo2NYwRq5VlNPR0LFyRyPuTQPeA5E
br19cOhJPjCsSRKGs5ExydCB3tP4vkyCZbYAhyO30e24tHEmc+d+DIo5wvMsePCi
XM8XduHvQ/xsn6Abd29IfNv0D8Cg8Vj/OmrbiAyfSWz37QRRqlx43xwdEIGHdZvI
D79ZgBgsVm528RYkjWQy7HQFqfL8QB74Rb5KhLyVKGeStcnUBw92S8FgmPKeg7Fg
d2JXM7vAVa9vXpqj/Rt5amhEWv/82Wjc/H06xuapDRkgoFt+3WET7nchwU5uJ4Ds
OPco8nQaMD6MuKs7y3q0r4tRC4ZiV+sbnBter+0vLRy3ZnQX3BckXRXpBkchvh6+
qOvW7ewUcxMKrTwzORj+UUaRXpxLOmxhBZj+pvonreZTByxxxlCmdjzI5IgtBY4c
0Y11G9N3/yGjzBXepAR63pGN9MHg/7HlDioLx/ETZbVzf8OoKbzcXdZunpC7EtE3
tVP5Vji+yf34WINjBqg4hOv0qIa/THG05OxCs9ZyERmWr3Th55c2Nfot58zeJSgd
paze+OMi8GrySr41goedxfml83H5Bi7O2Kru+uS5TSEjRgRfsGTKeKw8xWxxYpR+
sZvV4uj7eJabo31WKxvmgTCn98yQCtDS9ALR66tT3QZmjNBZqKA46Es0ajnE0oAw
LN+b/+4s5w/p6Zmuuag+yViDHzMI8T9+RLm8OO2sQKRFnVjSfVB07rAJ2FZGuq0o
mCXCloQRooQm16cMWl9KdHG8WcgiWRmcFeQq+K2EnwEJkdmGq1TYiHmjuLKLSl2E
x92gHL+/Bpbv6WUtoGVW56cunDLkS6rcnGNZ/BcJg1xu9ga7IU8HWn7IYVJGiSCy
5Agsk/iSYkhplfRL1pt9NnuZq5aCZ6rTDCnP68NsDkmOzCsWbLkV/x3kPqsWNFg+
KWsUAe4FlhQuWIExoDR6i6p0sLUiIt0Jg3xtkevFoGi1UVGL4H4wDqAeEXFTPIBF
1/jcQpP/opNup2DDTmqH74pe5i1fnlE4rQhk1bVCKukw94Z/cBJzhvKlJtmwStPv
nXpEMLahlkU5jPW7hgKWi7HAW0KeswJFVEeJ2lQHYMsTZApagz8VNhtQ9iv9dgUl
aPPmDwoaJHMWUZoObhPFejg9WVSn2/X8QnK/08vMpj/tngerZ8Yrr1RRH74gy1BL
p4DOZBQaNbiseQxX3EuaJcWpG5nfcbm1EhqUTQDYlCV0IeTczw1D7bJeNaMmNtu1
VNUgTzk11YYcMNkaudiOmCcP5/FWvu83kCJwnFP93bcy7bEPsITPrP/fw7ZNJQE/
INPJjKMUSEAdu4Q21CJme1/glhAQsoRcIhpirfzB1pCgs3fen4gAxVDp0vnB0aOf
Nz6aj2wtruwA2PJ5C52SaTxKhMzeQkVEJCOuL9N01j97PIcH6pjigqKU1Q3I6i2Y
pFQYw3Vv59tg4jx9ikkJpyvgJ9h7tvtLwkLsni397HXCS6ME8wPjbhsO9huv+9W5
4fzlVEKvXTADFlJSnwCM3aNkNYCXhQLSgUGdB+MS1s0vzTUg/xxZMvBl7VvtLb6g
nFdCSufe9FSUgh3/sxGzRT7UcCPTg3760Ox0ZXEOl2KyZTsSCBd3pSpVrTvl5VVT
+v8jC2vMs3/3ByGUO66De8r0ejpyttfzo5SpY0qZsRDFDed6aCdU/uDfhjeTbtFL
/9ofF5ybRYdt0mQ7+X6LOar9v8WXSVVnqj16EfRaTUfwPIKRH6Emm6Xjm8NU/E6N
C9pnq2mBWr5UXP4VyM/HS7Uq+ON8Fpc1173y5WA1hhkQBhI2BGCD0grGDST7CMiS
LqrKfu6Cjl1T1E7bVHTRs9RExEsBzeujxWUfZ6fmS+fI/do1zS2s+/WdYvUIKBSU
ggcRQ0C0uQ4ST0yamTAu13lJiWemueNAy17BmEzi58WuLW48JdiFEIRFzmSptg6D
wy+xCe7iHbU6AUHPelLlAVOsrekRHlyUHwv2aDc9k4jaAtv3UKSPU4C9q/7XDSvb
dPZTEOTN2yzMNoDOIkhXJK/j2BLPEvRu10D9U1ZKoNs1t8L25HD3p06fy+AmHGuM
LLG2KXVkyE79KJsgwDY1bAJl81zQxjva/aTEXdPx2wEI9DM6bOOQ/QWjOg1VPL8h
GMG2IroRKE+8yGcwtz94LotZSrAvZ3KoK9eWcIRF7FKkZRjeBjHnLS5g7ZoZHxlH
4sGNOASRRXWH4zYrfUGNvxWHJ3mjJqo7aVGxUPn/b/gdXq0Jn2Qrrd24YaIWVeXH
njQTvr83Yw6FJbL8OtLrza4cijXE2Z7OKT64g5WxkcZczcNShaStlhlgBs3y8xFm
O7o13iDGx1FXBvZRkIomXUjUS6p4jIDWjwF+/mgD/ud/4XMCl9bVxF2Dfayh0Ie2
NV77iCWNcwpdR78GUKpY1wW2FuF9/4stu1ixXYSMUaGA0BJZdTcnnM2wZDAn828O
kE6YjiwtBUdx3G8KikOyds3ZgrGPhVlUzmNR8yn/KE0HwmeY9Lpvoes9PnXViCQW
ptkIWrGo9Dyn+AN8frESN75C6ec1735bt5M3OiumaSzVmzFSFVLb+qrOe+abEW67
7AlNtjcePL1mtgGtyTNqIbFlQrCX/R+Ugek+iLr4TF8YMwrW6QsMG8Awpc2P7DUh
SRtpD67VtadA/bHRy2ExawpujQuc7WTSDrPeL9V0oNdnB7vMdsKtwNydVQleTW/p
VYJIXc+uMD/rqIT+tMsfCCN5CdxfqzLdsrhjVGWIRB6s/+1p/rHX3Zj2UiGZ19eZ
xvlmJxy/aj2L/htou+7wCqzxJ6VV6ZUcwJ4xV8dSfN8djlk188FctbLVJnxgWsRb
Y86MdNcsq5aXRSzwweI9FUZlF/abwGkCU65EEAy92lIhD+FGVYbmT/YLpYTL75eL
0rBu1copsceQsr9+s69XKtd74O+D+9/L+4Wl3h9xgvfhGHWuOLPyufYr3SaXwUMk
a7fm91A4obZ7y2shRIXruDeLYIHnowUj3l6qexJ40OUTLZt440lr1GxRemTEuHqf
FSF14xbAtSI2OHqZyUuIRXwIXu2TSUH2PQfdCRGeoSsUa1EPcXI3lzICxN8zcAGL
JOZ61DhrRSOVLAqas4804Xm8ClcvpU4Q5mot0ok33wqKJs7HWrdRvxxjWLkBw48i
Is9g302L77d4YCmxqywpSIGfFZcTP/hf2yeVqm1jgEK6t5aBXJZ07+e4xOogMFEY
JAswUbh/kA2jti5tV18O+K2R/b0VvDHcMxzGg1jC1idkMjjqA6Nptv5GRV12Zbsq
Ij46mmfodeeMFm6v+m9LDu4EXpQErrSPt5bMtUvYPoHt29u0m58D4savhNuoy0jg
iP/FkNJXTdxF/TweQL5TUoqluQZVUWujEshPfrdLvvUTN0JLowUgRZ4PvvcBTy78
fLzRTk4yoSmXVO3MW3BQsDR+q5MMpa1tkKT7TnpPxBknbJ39y8Hdii8n4agNfj7c
KesN2CUF/7XV5/DSuf2CERrjwF4RQLOr2Q82hh251fgJABEN7yDvDWBJIlKhWna8
8RsY2aUhf8cWX++hoYyaZd+JAxau13I4JKygRVKtsNmqqnd6UKOv/zpkFX9Cd6pg
cIXtg/bU9nFMwL6X9zCYzXsep2iEcSgKTSVtE8GonKhuWwS354QMNVi96vXUB95x
RN2ozc0S2c6SwP/FZe+ImEeGAjvE9KgcO7yN84jsn3GNw0VE1X6aRs6ecFYXerKe
fmUC/Y2Kvgh2gRc7NPECzBmGjaQzazzGH8NFHRliND2/i0sJB4yZXKOl0jDOZ6IF
Wy1B1vrD7imF+aDBC5zlTI9Kq37CWiIiojMXNrQyonTumkq2elDDJ+TtJ5D5UpB7
CKE71lqGPPdWHm02nQ2XMwjQmRhsLAap/LTQbFfR+qx/A2HEGxeldNVv+GBX5n5I
4sCZcFe8rFsyULDKYzhxU4BMbnQDx74HrKVgpMK9u+U+5I73SI6e90wuGuVpXXaK
7BFQ+FKNtFLzCMthKCpDQiGWwdpNxuo1Q79XkpKdhWxmp3LYiQoMR7fcTLlFRpMT
ixbaMnkoOxvUUVg/YBCHQ/IsKeVC3bYG+N9ItLqNJJhqad1Xn/J3Rk43h/lwYoX4
9D7AMKfIPgzFQvaZupdBiRaD4Tc+fq5UdmZgKLXDF0zH33quJXW0FA9qg4EWf85H
7ItR+4All+Tab3WXdqC0puM814ZlOa12KiAAJcHvWR/+Ah+KJdYlQbQfrURjLJjj
ksFk3ij0BbKMKCqvU+iBX7CMvMs8MK3X4dq4F8saTDKbS3fKExhMunh2oB/hK183
2kxuY9DSKl4SRBCn02+Wk2a1S5blWKC/E8BraCL9ptcIFz/5EK9YsviFcGMXG9aM
NkTcXPAoiYzd/HFHComXykEm6U/9cEwn1TPTt5RTI+CAHe5H3T9V340QyMbLKtFg
ihFOYSIdFrDfUYujLkeM/5zRuQAq1vc+5NwcSYHj3nB/1Y0x0Wm4bSokWAkDk4pA
2cMxOO2U5FZimq82K6MhdAbc43x93iY0GMIGScykJEVoaa2QNLlMMcb4RnMB7YIr
kt2j3zBmUrmCsUN2TdCTYw+lqRydH/iObP6wG/S2Y4D+Bd/BSwQHwa0tX9orviu0
3dUHaJrJx+I4ahqXlO9nNbq+FXUDIJQ0dofTAmeKLrIxC8LN7e0jj/+dRM1921Xy
O374dXByF7avfGX5OKJkT2GKHRhpc43Gd1NpQaWzIYDnKTQAjw4IBIZM2pJKxI8W
1FJvMVAiW8ESSZbAEw/cmvwGaqh0IkDKtCfIxpop1w1+2eb//VSFvSxLDdQZvGG1
VGNzv6up40XDPvA5q2fiF/GCnxZSANHZm8iLLN5tw1TXu2eNy+PSJqIb8WdEPFiR
npx43zgWNuWV2PhKRFJMM7BHGUx4ywEXkzPqqEF8JMR4RdpvbQ4eaofosSbeC1t1
CetKpN7eUS3yeSaW7YnR8Lx8wtnTBNDsWOy6Sg0T1WJp7C7WPHsQ1nGMXNhw89qJ
nu4maKjubblRxx17VWSG1vjvSL+ynF4fYhm2TB/noa49gFZRKVBhQdYPwORSOGJa
vJSlvCPRVqWE554eNXrxgJe7/dxSkdYEAdNmfzoHdmKB/jlH+gIPVrGO0CLNJrcp
8LJ7Qg6R4oLtHhANG1X9nTdGU3D55c+tQEk5Ewroiocty7QBCy6+vvKMhUfQAIce
9KEMoVbHjeE4YNuhw9WdtPJJAVTBoS/NmGV9wkuHJc2B7417T31hAaqVwZbyqxUN
KxmXMDTBy2sRmJf4RxOXxtqUIwRqrQhZZ2+pYj/0C8po2KYQsZPEnAkJ/Ui2ocvQ
5ae9W9yGB7iBH8Gl/vpAuSTAShy5JLHHhh6/W5sdY2M4uD35B8LJLI5Tl1yweiKb
k07RVT/Tm2Z8BHKW6OKJHXF39lPPmDBIIIugM3FDHjlKzTRMISWJf0zg4EcWFcrN
KVsCABaQkOspcJ+Ss1E/Y8q5buK2utRZKOPfumhO0NRajFN5duUgfUGhBtZfylpN
uCC5oyk5cc7lxH9KIFxcXZjIuw6nlFXD3AD4Ut+s+So72vtQJUqJkzqRp8O/ISzl
TxxBvzC0FHQ5zF0exWBGP5WTQ46C+A246nyWaX1isWqv/Aix+4EDbj9q9wvXbSC3
zDE8w8Bc0mn8RRiHSMWn97TKo8QHbm1raGE2xHX0DGqaL+0VS+Q9WEwA/vQUVDpG
9pXAOJr5fHpkG7ggAzS6N1qQ7HPC8xssSH9RbCv2EWCnWyymxNRFi9b/DNpI2EB2
Zx0Qky4/I9QqP+genxr+CVKiS7T2R+6WFhaPDloyAg0F/H1U+6MmjIr++eMtGmXn
We0Dq2tjfoAbLGY6osOTD/kQfMtm4rSi1//Udab7MRWS9Ng4gzCifzSA8Kk2mu+t
IY0oj58jaQJsettbLJi7EjAb3PQR7MylmJB2LOZnUJWJE7eD95l6GvdbL574LrW9
hQi4x9p/EELxkYklSSu+SBmgVHp/rFwg83hKvdx28AATeM4r6ayTwQyZc+5tBlcQ
VbQk1EPZSbq9vWfry9rVW0Sif3iQ+XAHnym0hc9Nkl7W4k/8PlhayEoc1BG3R2f3
dy2BnegGo1e1mIhqHk72sq4QtkoHilYhQYPA62Vl8McGZDn1DUc+3FlHiWF9AJsn
a+pVyhXACvE3cPnWHubZ60KsRhyEgUhK62ZrVAIQjXlPckDAbGrt38eN1gzRGyTS
BQLxwHbzOu+RSKVZGNE3R6z8+kAwagZAGOPhWx0afv0PH+GdWYITJGnTgnq8QLVi
HCMwbiIH4lgTSOpSVdee4USDtl5NYUM1EtcQi2is1Pu/w7RPMWtsqNaCHIWn3+UN
G1Q+IccV6P8HUwpaT9vkgkJz31JzJcJGQ0U6XNCZBF78yUdFDtHE1NMc3VXVngr9
L+/4Jyc2qBkaA4Go5kzrgIO874cPpK6doKpQdcjjZ7WNu4ZbW/adG2cREreH6ANx
GbDqPFnqPxiYxjoHDhWPJxSyzJEMFe/sHI128gF3l/ZdTJEgURu64blOMR5lTnYU
/J5jZ7dNPjEMwtY9PoE3K5pZXafLNB00LoXVeChCLkLp2iMOb9MaPUBl4P/2F/wL
MTq55k0rcXEktw9ZpAQimVXKCgwnWDktkt5dogpjAMTeBQSCY1WWHoICrh7A/fJR
UcYm7ya8mfbdVySO37yIyKSwYLVsfJudrLObXLCr/eUtPy/pIQlWqqSzOTifM9ky
ZrCZk3+dtdiMht2xh+ojWqCM983Bp6IMMRBxjTvd6Ta8hD8oVDAzBuX00TR6h2Cv
Pglzq7tnqckT+fjPtKGh5HgZfO4vROCXhkXymhAA2SjmKmecF1ndRV9L/l5y9VWj
2O1GYw4kboW+F3ryizSkPnK5Ass8GygS6AUMGGgfA5CYNkEyZxKNVuWqYGWrZExJ
qQklNb76uClR4adnTchaeBfekIMz0HrxtUa92QzqOu7sRGKY+l7yGWP9wfWoWLIA
zFv/p3Uqnq0vQTDvMiA47KGEyKF1475yKM1yTlLugOcPRaiwruYrpex5KkcDtJdT
fmzxD2Q3Qrl+zXFsKFaKS4E5mXXqiJi+lcvqowhfgJUHAz1jV2kJoPe5h/K/+Ik1
zr/qtOtZg9d4x+XQeXE3tGGfCqf4YMhHIcjmC76iJGTighy2QPJO3uKXYLv3Zp2B
cpST3ZBYve6GAt3ac61IMcF8l0RGs7b/RZdE7AzxJMuRxbu9w366BzP3Rt9Y6CJ+
HjCD11PRABS8KsTTsLjE3DtUa15Cca+BAxSDndz2AG+09V8uAbH0grZAicc+z+VS
wJmjp7nl+ErP2ZqmsEcwywquc1SeS6V2F1hKZj+pRPJKx5Dq6Twe1nfdfQys6ghV
Vs2vFZKyXSuGBDR/oQrCOqhwlo+2R8Y5LQqXE7aSqxiOSrPzusCTewPyiGhagh+x
R6YmQGGFXownrfZq4xnLumWWum+9tzQVqcyeRsmVcQLyQZO5NY6miQORQ2asT9Vb
hj8qkw14e7a9DlzCPweqpqdgMPYQeCaJRVrUn+CATCkbqh3Q5bvrjHMC74qWmT9R
OtkM9zD8WTpn4gtKPzIECUyHhJ5c/bDbzUFY6IQ4raW5YoccU/dWBzxGiMlFVAbZ
lr6bGL5VuMk6INKRw8ladFjJN1HSjMRznGiXefbNM5ky5cbKmbUYn3cCNC7v1j6b
JkX+v8rp4XwEJx6v4A/56YwHFI0dQ8o3Yb9P/L7c83kTcIHixg6AuwVnjxq2SSN9
+1yf4sGTAr6wiNvpekOA25eN9gGvz/n41dM9PuwXgD7CU+1IbeQuDnicFuEd6qsU
+dcnqZYrZ3loMnooyQsatieS86qzQCokgIrSUKEEduAAKK0qnED/14UPuRUE3rmH
t7Np4786k28knG+pop6Ehw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Du+XFQLC6nx9kaju3tgvqH5rzmLCvMVbcgGo4CD52heWMMqRG9i7varUrI4T5eRn
9YVRu75aXy2E4hJ9Byubr41ZzrlhQ6YopYK5hC5aDq3Y7icabxe1QYHTKOus7nev
G4BrE6UX8PMhMKfKHAe/L1UlAiaaSrH7343VLLEy2riKVJ9xg1ANJBlFpHGe3szl
lp0HuHXpvfVQiupz07SU6GD/RlkgbkF1pUbkS6kEL6Kriker1Oa7dPk/01J5O4mZ
1fbC/+iVbH9n5iGV8HEMsShJfQt2ynwadLuOgAaLNsXz9d90ozkQE+MFin6UprIe
CCcZsTkJDJKkVR7ct/4grg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14480 )
`pragma protect data_block
lWqvGuG2VoKHAPdhRVzopHcvP7eMwM4p0K2no04u7S/8KSDz1CvFDHcmFgJSnvvr
Iua7d114vQlkwJZeVOcsSHGyEzPYMooqHINBCP+QpIMt84sjusCS3uEvpwLajty1
Uv+pZPraSBCkKYtZXQBKd93WbhEj6DKIfr8+NuZjNofrW6NB07CyEy7fB6RkiWo1
BJvenGSbiVYYO1Eqmvd9SYJKUnwregWMLTxBSWSbGmF0bqFTAkTEnZRVr1BtasqP
Pxv7OJuDOvq8nasfm34n5Np1Kgn2iEYvHWnK6YYyl5e47gLGNegcK8oAwlZGhIw+
FApHTx29WZtAtxgq1U+DBgWrmZIgftgbe13vTCXApr01dO+pZMToa8Q4kaViKodL
pqD9nI5bcBavTFjIHmC2Bm5xjgQdyUuGVba38MGCsBBLqB0SEBsa7eIyEA/CCJ89
RDdYP+islhC8JF+Vt3WnAmRgbDN6SOE9kv4SgBbu7F9F986BQr6RMwHjQdd60Dtu
UZNfzdjHUKjhD990pxlP345GXZZYFxJn0jVG3/TF1xX8/mFLyDgOsA0GegtFUdTR
A2gjrByPVx6iZ5sWGA6CxNyRCJX1NMBfe1qWsZ7zgeXVd+WlF/YjnIB/Nqk3oEhy
v1AzA/n0diGrXO+HUut5iDr66U8NVenFR4FauQx8GGYjjMKCd3xJElZQJw+w618B
22UY+L4gsCYtoPAIKWX5Z9KnRQ1U6zLnYi7zbZk/8ZgzlSdmnouAZwAGgvuwC/Q6
0cv75Ku5Btrw2LB5zG7CSDZ2cRo3JqbeclrMeMg5zDUjGnoIjNDSOsYtlIGH1CIi
Y4N1xUBT1J3750Mm3fH34Mr9zf/Br6nFI4R5DlOojfI+zIeZOyAvNANqkJ9hRJl9
m2JO4qu94xi+d6QKD5+Xk+ypWCkznenPxxquqtb59Y8vhrIHTACqyuACxx5GO99X
NZiQGcj+x/4mIt6BCXMVcrIsHthF/Lp/Qj81Ye0fVCrtjDDR4Z3MRoGUlCfJqIvM
ja5rPnEs+wpSdBFaIeyNICNk1MRYFD7svPb5sAce1xbZb3nU9hlqAJ0Ou13XbS58
1xXNvmAHCqeIBs9NMu/cTANXNFNLR2gA0dAcbYPPdHHkLyCj1PH7QrO+JooqWH6j
OFpAox7Vdw2xgU/NBC03PZ83Ym0pAnHW22zEsTI7+RoZfnwKqWkwCoo+dlPt0BIG
UpdoFg0ESiRU0CK8+LWXc9I5dT6z3vR3PvGcEZkdH20mYusKjpvR7GPmfYqxXT8e
Z0abcnM85uUZ6SSq4CPjJdyH7D0GsU5N7Cg/PKCnppfbSEJ62ShgSAJYNKauAfAY
FhuoV5eGUKMgkfb3ZxUTSDLzs1kdKWu8WFtvcGxK74C0o3yV1FMc483pYT8BRczf
miwvKIzBGoW6aq/UyBO+d+96aSsy9GdoWg09eK9GOiRzTUB2R1anQIz8TtHmmtvO
1PP4XzKgVEyInggg+xeC54CA/a/KLhAT9ZICJ8Y4xehcyBcwp7UU4oE/ZZ7c0xFj
Vojkg0JPFh44YYKN/kF19D4trbW0bgreSnWlLEZRMenbuAtzyEi6NmcsrmQgPt0T
5HYfVdz/OjJu92St0vnxWBjS0bJ6H2e7CZPFvzSq9VavhpYhEEqZixE50b0gILrs
1gmSR+u6pFheWkrQkdUa6OBZawcaC8M4sTaFyBbeAT4Km5ZtdbPJnqz+RHGX3CH+
InpwupoMo6yI9FmMzWLPmhObNfk259pwl5M+7ke/Wqmm2wn4KAEnaE8KXWh0pQjX
0vNGjsDkt9Z3PExSfLxNKYJaL6o/IncBebbDw/tfJrjTpzwFskmra4u/SlPGySk/
hA7xYIhfNE6DC51MPt96152R6S9qFHzpxPsNoDIy6xXlYclkVgPdqfdAIgMnV5dE
GcG0kQTbPTEJYUA+s5GN+bkJYoXf1i9tbEex5T9o3FWByKem1ly0SyaKXxV05qlj
E/Z8k+QlL4cgAt3zOE0CbLf8xHcG3r11NYicsVK4joh0jACOajIpeIGueu/czMLF
nLw2VNd2GGrd2fbBNeWtoscSPXkw/xCW3S85KUY0cETfdV58hjs3Q/LkxKdYyk93
PjQjKK19xJYamLaSQRtpw1ejaBh81pHGe1fz4NnsCXgQVXjv15zwag3WV4g/NLST
dleJy+ICRwszlEcuW0QXSvs9AX/3Vq8ZvUD9LK9apsfxsh8c2wbkGpJUWxAECw/a
Q/kUYp8r2cQUlIhpz6phDi3SIU5g/6SfusG+RfB5ZMxf1A0bZQXANbS9IOumrREh
kcCr5H68EaIxOiiMw89xMUqhFyAc1+UFW3iywpLkP9cy6L3ATdWA3uI7bMtlzdCZ
zrxnQ9D3ZKjiSnI2VrERftyLPTRnMYULQCbpNa2jQgL4tu+wNnD4qWjenn4L4XmU
Kjh4FWKpWSqvWsvHkx0uHPxxX6Uw8/cXtn2Dr/2rbxack3rA97R4Pd+q17SBfocw
TfZfHddUGzvE+5dOKp0d1Jwbmd79kihKn1S5TyF/mH0Yt3LWvF9U/EUclzUZvi1T
PXHw4vRpB8ysHim3W4BgMK/m7XCRi8esw53Y9Df4k6RpT2FBwvZeh2xRsRW+MtlP
WanETSHzc4y1vBxQ1KVTZtIkC+QMYRmpB/qeEi/WxZLrS1jNtxhAx8YcjWCi7Nqb
3IPPy34UgGgp9QPmQtBY6dqozYFC99sjVxGwaS7ywIjU7KKvmRBFE0jvQK7ziYWO
vBfrzvlHHhVaYO1Nuv/Kp+N5kLTUxe7IpUkMQpUFWZGOkrV8irOSolKWrtQBTEpF
C/OPG5uVDn8Wf426aVBkahoSFVQ1SryZgO1sH7ee3bMY6zdN6DCenPGM2ofyB+eg
C/Ay8hbloypptNkMDj+fFO6P2EqiAXEW6nqN+u2aFbpiHBRPZkfCnHZPi1lMqWBx
pR1nERjwSux12sCbekuYg+e6VFK4/wwHwboIEFkCHpvzVVIFBc++g8NeIBYARtl1
6eMC5KZd9hFQRKjwGvU1nEAIsu3hkLk65p3YP86Vvgvhz+UU0ZEBgIce7fpvMyvf
VTL3tKKXqFpsyNyoeqfFSZ7ewX2DTbyn2MzDQYHAqpG2JuRGrRoLj3luOocWW+rh
hwVPshGKSIIILF/akOUZsmP8hgma3zcFd3JgAzi7ECTdZ1Y1U1iCdTYNUmH+A1Pe
FcFgQZIJNK4v/y2HFuL/BDCpIJKPvlHIFcUrXgZ/cVTonkifQwnx8ToI/f7FlEU9
xoInGx2iu1hUgZLDSWL0MHA1u9jfTkgNfyY6VoGbB8/U5ruv+BVU6wMkM7N+Hl5I
07GinHCGK5YUiylPko/yVu/AlIu+YT5Cos2aYHO69qDi32XDe3v7spHC7vf6lrzv
/2lV2xwK3+NIy7v1XtwRb4xl3HyKP6e9sQpfXXHxfglmwgzU0X+mhL0e04N39ItV
0OEePpp9zwma5krwALFBovZEOhJot8cdNjkwNWeR+wAAhi3KU6oN3728ZgYxPXzP
abCKWBVgRazLhJRbdLxMgjQWN3QJZuJ83sieEnxftZNqQgf2LSI/OJEriro+wfpl
CG/506jnuj550DmJvzEBta2AQjwwAdEoGaVgsxWyq+6vZtBWaj+YlTn+wEdHuNF0
0EdbGvAYzv/tUXmFPz5BkBNynVrqpBuDjlKskdv1CWli5kIgCPDzrjSBuCs+cpUH
QeF2vzevcNt5fkH1NtD06utahxP47vSBq7uJX4JVGrW/QPUlcdAxpDBasCgx+tTP
5PKL7vHlz5K9XuRoE68zxFfq/2f7DW/r4CgON2aoTn+l2FIEL+sfdvPMLAXDe4Td
O88TQD9JH8JSqit2+IodBsPAGZx81LqsaSEiM6BXnAqU4s1Ir/YRgY3y7nzZpORV
axUX1Jb5ChimApux0PdIOO5eI68aeazmsyPppIDmYP3Rx6e1uDexXW2OFQgTlg/V
iNs9PfU6HJWYbu8tbdE///MxRcqC0GNSMWjWrrF/fR2gfMjodKFoZlU4yipcQKv+
gidOMntQmnZhUnj7Fek4mFHiEM1dU5POoeGl+zFIbM5X3OG0qfXzcOz5dMjs52SB
3fjZz8n/DqtI8TMz0k7t6q/2h+1os/9MqagljpPTYzIEim1scIJ1bVMJ4USlku2l
kWvZ8t8N5A0Q/DHKELikS4lTESad5z6ob9C3In/sFnQ/T43gvEA/BHx8W3jYWwsO
80GMF6fEnpS0HPesfNLQB2YiNTCfd8n+59N9mX8f2Ngcuu3uF87/gH+/CdaBkI29
nSnMOkUD27tSo7icV3a3o2tyXYjibyoBc2jX7noNOF0Ptz5GM2F7C4bRH50rQ/Lq
+1QFc3uTVbNdt9q6yS1D6iWdSXUYxLLK6GRIEOvAQ7Z3Fi/z+vfRJb1aiGjkrfaW
xQPSyWBAWJfwDMsH4DnDS7bS7YdIFut7cEAsoCuoOxNW7r8bwCIwCGGuyxWWKeRp
9r+ZGCj6QIPm/ACKBBku4whiOO/5WJJxGNq/epzbskcIsxe83IyfyLoZqWGwPJK7
4Di+OI+Fo0dxYy1HKO1AIJfh4CZYtGYp647DLrDJFW4pIWAi1ushkoyWz8tUYIAx
hdIrBJWEa4Mjk6r9X5bAZpg0ponktHX16whyqxWf924GOuv8AbCS4x9+N06YkWdq
ei9hRXdjyrJDKItaM/w+3t7HgtzFI9SnYgyjt2WWOBsbs4MJdr8Tjgcg4NI2EIgu
LMNUDwc53nbXrXGNKQ7MSmLsXv2QX3IlVjYYP/2hN8VQYFNNOTdsmlKX6vO+ilih
bSWBiECVQ0jGKTbm1dYpxjLGCu+7p+AzKmZ5WBK/dPB0szYKlG6c1wBp3VwbxR5X
L2RPyOxvysTMWI1tvljZ1c+jJ6Ymks6kPNMT3I7uDv1a6HzMtm4oIUKFNoGjPWDM
o/jBgLEiixGbmnBjNiCG+SgeyO7NNKnr9z1lGKAAMea9E4SR6207zh52Finaqo/Y
9ju7r4fId4POV27lU0E76LfcC2MR+1dgKGHLNjVfw+jaK5DFrp9vog+ry4f0672y
RdyjdYmX4BxREL4U6rE6abJKKw4QkmB8NPHqxIFIcAHiGq3E6q3U950h4dIsxv+P
hYpHnJlduP2m3ZDxB/bhi31nw+lZ0DsySVGWLX5myNq/dB9PBHOwjhF3rVZBKacp
5ZIzPmlnnBZbdSYssabN7kNQQ1VNeIJK1WH+HE79xo9eqsUeVQ+qru6286nWzR+t
a3D1UfGxCsXwiUdzjdn8PX8VzmCMlJZN0heT/XnJiu+ikhLn5dKnK9Wp36SvONGM
1RuT6DQL6+wlPLztea6LwXf7wlEjRo2Ov6AbxoTIJT+CcUZ83IO4yGhPN5iRIS0c
NIxKckb1uq1iCgP3niQqpsDh0eZt4B9h/dWPPtq2clLOdXSGgIGWoAt8a3gmjptP
Bv9EMlZbD07T+h8lTPjA/I/UJnD35/kPrCSAlnY+mMN+OZRUZdWAnmqCl0LBjVOj
TvER0/IH4ZslvkzfFz7F2TeumRlwpdaDrwC1+AutsAeKDWV3vZj/b9f36Knb2JSx
pcYl5KJuylR9Af2ab1dCX1JlwsxihHW8Hqp29cCuKPsWskb+oGQJjrYfzQDrtVwV
l8cwLwerk5xz1wikliceqV9qtZLSHfcYDktddfIqFhqzcsmu02J0yaVZICKSfpz8
i0/zaRG5tXraKxdAGW7xRgXnWX1Aii++WKsq9ZipS57SozbntfVUMIEnNJLMLO0q
0CBKZkiJuM7iJ2CQMngBoE5aBoW3hyOIh7aoPQLYkQZHMaB4XlDjr96BLaiPI0h8
Q8Qy8wTN11ubd+5HCHhsBjk7d9+5VYOkHUeOEimKz+ItOVRxPvqc67g8i17GJed+
4MQ8ZRYclGe1UP9sIu1fySq2RWpHy5sh97QQkngW+Vr5eJU+e/vCHw3XZLn+bkUg
+7CevFeLWsK3xuMI1a8B182tkfgC4g3OW0/uWi2ErnAqlG59FpoEqzICBBBLG3ll
mBHi1yNCHgjV1EkelGU7SWYzGCqdo+jf+R8FQZNWXy1+hzhn5Yozw94nzZx39VIQ
0o5zLuHjLKiYb1KTcpK4TFK7QJgObl2Ih3PMsn7c0CKpdcwmf4RhMJEgiVisnB07
uG1bdaXCcN00euSSfYlJLBHLmHUylh/c6azuVjZMw5a2jCfFHRLOo83fbA5x52Zh
xy6eOPL3QdrY36kGPJkzcYV2nMMqpRYMe8H0JJFSjYVfzoVh5lyI4XiPxRiDLCEJ
6bFm3G9U0P8O919lqwlIdQgO0LlitXRTdE9kMu5qd4gCwfhw17ylaR+URLSNqHfF
l+NP/n4qmiwHcIpBiiXYdsvOzvLtEenOpW+ga6wOuBUZPouXMR+G58q8IE6xCEUX
LEMUA7cKRLqILt2Rd+Hp/wh/ZW2E6y5wTajVzthdH7IqUsSovUQeLvF4G2nGLNn+
KHieHpHptCjrD3A9Z1BnHGoU2m89YSAmncilfNOmsLi9elsTjmONdlu4RcMCXkuw
pEDVQDbdirdBthLJKr+yjRyi4WaeAm72Um58hTbSTpNzPBfn+vjnoYwojesdQUct
ljW63wfk82yUfM0TFNzI42gj92qO3PnldzF7Ubve4SZDO2BLUwhj2WonY+0cpwHS
wbB4auyWVIzzdodjbsuVPd/bH/JjcluDiFndQzj1LnBL801/QkiWJbyZckQrl8Pd
choGoEAglB1wvNkzqxk/OwHyfC0VSeNNe1aeOockueyKJq3y5mlAEnsfB9iKeqiq
FYI8DmCfbI6Fzo23y6nVzLlIhV51NTRmC1+DQMb8tyItrI6VWS/Hzg8oZH7RaxEn
WRgqodb4KKekOpxB9gQnkbWWlZVHFlp1ik5n706Y2JgemE+ShP8Z8nL3ZVT9wnvz
JM7eJUxtE3sIsni9HRSdhqf2c4n5vopVvNaFMmyQ2wcOxMTnfkT9wQMsCJaO7hPm
hYHIxx8q142LSjW1okvwASZf+ILVvffDpgaqVCVJtAEZnTbGBcwb6ntqqC2CfXpy
EaVSDIcNZcmqI2TCsmnn3M+9XCA1Ms7HF0Ugw22e5AakZZJFc4R7ATsQ2CQr9m1L
rnX7pqT8nzce7qc1Clr5uw5odI8hAipzqkXnXAwvSnYnWSUgHvupny1zUVRolyE9
e6Vma8Dqsy+Sb5BsaemIwQmRPpeiyPy1U8OYMl7rQh1c68ZRXiP8oBNFlp0S0fdu
VxkYuXv2lDNAIYxgjNXUSL2zP8F+E6uciqnndQYdbvIY77m9AXSXxe7yLNz/57hS
jG6azK4kAxVqf2qlBWt+GKb8iZ2HSzKJWhLHqzXjMjz5krJD6t7GSjTOnaCtZsBk
DQylPLJaIxG229tiDVfAdxGeLrdw6RtH6CNK/+jimHbhfa3X7ogCoCm3Mz9VnkdB
uINGNdiygRFzVR+FG6jP5Mvtztai7NMMfapyH3pJaoBhZx+Q8twPXDeiSy+UmTyi
lvyYYO42Ltk0WMSXXkQRM2S9E3xS4Kw/oVmrvXu5LARE0m1ebTN7V8xKQwNYT+qu
X1xJGnC0g85+/C5gFtk8tlBCM8f6em5QTmM2IrWAVfBhRcarfVt19w+3MNyIhFf6
zifT2OxQViBUMbDAtM5gQDB8D1dZZqUqHkcO8uiZjJ8ora3Ww9aGNX5rr0rPaG0M
JAvckVziokUiIXw4Hgn6MbkxkHyT/zD4BMQd9oiRqn98pLjgAj+GpskHTPbO+3U9
9yAwDybkysQ2rmRwpAVIowdq7izkJDSCc/rn2pVih8AfJxZgmaosgdTOIddL+WlM
1TXlyk5KvNXKa67Optmc1u/hv3QIJtOgG3c3H6bHLxTTQfP2SYxBXu6zjj59KiBX
Rn4JadG91NghKNCqYtMg3O+FJi//VnK3WLWd2OAy387OAy7szwiIeJPlh7jQ4mT8
Gg9ObEgRExLxiMkBC2p9CKUamp6BISks4oODuFRb64NNgihWcqlOzjA/+49/xL9O
BGbkxiJ9HlwBRbk1RL/2lvVi8j9OzZZnDK5EKT7FLnru3/T611TjcBfx19rDOAf4
/PdbB2yMIP+jtdRLqSSPZqnIPnc7luSdqgLEpywAGQN4Tq0eaekPgFJFGHQOp6oj
YVVMaLxNcsDHxF4xOYtamUyvrLjZP4P9QhVlB59KzrUz7qP+r1Uiv0f+WZdjVyPY
N5yeQ5jNc7ePyHd5c4I/fAaGd1Ql/Qd27L6PeKAdhNoRDGgJSCdyesgwdMkxSH0t
Y5+7PI9F+8PPsbeImutM3uhDYWZKjO2yrNJ94KCW4DUfrJR4VygK14lGzfvCYApq
UgBDr6YoMmTv2MFyeBH8uO0ejM6TsutcEvEW+lbCewirnd9GPA5HZV2sBceyb0Hi
ouhUxB9d0g+YhEGCOPkpyc4iBNSNjxCNIbKc9GTcNQY8AMY2NhIyU8K4Ea38VOE4
q3jqI7iHIwOLRZXUEkYU1dv22ePEpM3Mkgh111GACsGFxsQqI36YcIWReZDqtnsi
RZVSJNcx14czE1h0TpjfpTWVyIkvDWGehhvkVMdIkKiJtphsG68OuLVBWHGFDmZI
r5sOMteEaWeG8Bc+ghLREp0dYOXuMjI6MH5svIWimcaaN1buqHOGkrlrdnqQnQeG
lQoyk8O82MK+1Mx3Z//6SlAbnvFKEfUc4H3w2YKf8ownEUh0xj2sXJt+wit/aIMT
jawm9PRlm5mZ42+8V7FXljEvGQBJnaZISWzxF6a7g+tnzwFM4i3b9ZWddLNyzo1r
jhX8Y4eJ94gZAtcz0lpoMSt9QT7zD/b8zIs+cxlAJl+uZr7RtwyTyHvk/PnxRY75
uKGPIvqt41lPdeijCjsum9I0UDWLO7GfsL1MyqVZ5Xay4Lm6x9cbeqqVkhDUFmj/
QTzWRb+61Q9uxNHuYgl2fB9IvP41mrPb5q4WzcJk5jyZhPlCY0A1/hPEk1yOfcOt
RvyX/d7Bp/M6YDFc7Zz9rx9gljyN7k57VQwi3EBjOPpVPV7oZtsR0Y3pig/OKI08
CJzGvIcGJzyEjLJhOrkJG14CNOIjtaVcqVTixuq6o1QAYLgtNCNYJ39elw0DH/vH
ud7H6sJXKJYcK69SbGEN+yHn7Qi5VBAF912IFoXCFpTCfF0ofGh1LRZKK3ENfovB
KuA3zeV6zLb0FtqSmv0c0kDQy8uvoRsFVjJTjRcxQX0q5fcflReTFpysa/MOjEXK
57WVTlDBGtYtSczFaSPS/55TsyhATUsgR0jTNJaoaDleBxx/F41gfXYF4jT0Ccr+
vAEv0is5krvYkCYDKGLMlC28LOOipJCRn3a/OqFSg7YVwW8z4qtGfJCKgG8aqFh/
cX815mU3u7f9dxA/is3guqgocLdydlhlXVobhqZUSxhkS/oIn1KMTvH34wp8LJbS
0ah9k92SjxbINvd1oYtGj2PsaxhtFUQ86CFk50rnMORZWotBscBxnKxonxiTDDby
hbJMXZcQ4n3MLZJBUsV7MRAi9Omarg6D+vlbXQWWrER1bFVxVn+tZ2i3qMNqzbYf
37tPYvW52js9ZAy3Dx6Nzq6wp3/+X7eftM2d6xR5jT8T8wQO/G47AOPnD4Srr8U4
lZ8saZAS8QZHePht2xpzIhnfSFtGfYeRvNKLcfTEuT+tGw/xTGoy7qebmajBkxgZ
ov1xgYrxZKyk9202Qytgl1jAtQZsEY7ruWipsqAzDXry8eS6eh0OvDlqJtRmd1U+
dqwznQ4zcR8Zv5g3EdLWuMEWzOwyh71brgBu55FSa49It98o/LmA3eu2UQeqD30J
ofgGwYNDxAdhlGTAi37Ilr1g5OKSxQ6ZhoMFO/qia0kXEuMh/9/dYT28j8N7Yfyk
e1xDoaLigANeaoOGFsMkld36/UQoiebHpgupr89oJbgOiiSX19KJywxbWxmmqw2J
Zbz2H9AxLK+vXkXw63vNa/BTsPiys1+eySljGPW6+x//8poLMNz31Cu7VafM/t+s
XIkNtgZg0qSGKapCj8HwXd9VDBXAunkjO+RdnN1A5DNB1b+z2aDjRn2tw7naMomE
ek/fLzjj7WLG2B1q0fOfSszQksNxw6Mg9/9M4a7VpxF9PSJgLoKadezRx4M6H1d+
UbULe1X5vuBEmA+Q61bpTxX8+m7pm6Hjb+h3vBg/dV+kPpiay7/sQDcBuOeHQcDW
RxDwaaRAfHx+4KMjEbnVi7TsxOxeVfHwFjZg5lDZ4C4pOevuc8bx1yPdM4Ac4bxt
O2c0XXO3FTBs/VShgucEe14i3P+80VFpHyKFJOcnG3D1c6EUUsWA4vrmA18ARZSu
NkNv890IaSKyKebinLeAz1Gj+30C+GqWnjvW+uQCPOnFkHbLhIYuTXcytEIrN2GL
q94Vcr2r5dKaFq8gf2iSbwikZhCa1O9Z+OxeoHUdamPH+uxQBpt8alr4NsbjnnLV
ONwjimmA4ObYD1eRdRY6rjYI2lv0YN0/uAZujeTxKCLdrh4hzPyGb28zrw17/0yf
SC8yEeyuZY7MU3Cg5C47hTfbI9tsZsHphTIVD7iihsJeV8VwbshUfYNUPZBan0qP
o6Fw9VHRic+LdxYFcNVwWG9ZxEsZ+pNXptXATzTbt4T4XA9085bAgkrrTCY/QeR7
XKtgr+ld1GEX6urTAIUnOIhW4hfTICoMDhOo51HmMfze8AjqrTnnOvTHsFLUvANy
ZHlHJZzdxBCPLiCaqYqTb4HYIiawUJz25x+ngTvHdf1XoHJJ6xRuLs2INoNwu4Nr
f+17lAIjH949BKs2xaw8EBAs5s2fE3iS+4dgMuK8tUVDa/Vi4VRYZ7cppgIVbs9n
Hm5u2MVWTj32sP5DbJ8kygPxpvV4z87YxNIfRdkmh7bspUFX5C0aOMopMlM3+BkT
G5GrNI6I0KDURz/wDtYhz2ZTWqFKyZhjxRH9t57thdhP65uXUIwAKRYpIycUfvw8
bLAGUI8mY+XdGpbTIRoEQTMB1EtSISU9T5CclYRCkM+ReqfJwOTpTIgekTpo7csY
dkL/GQAD9M0x710CPDwEVp99cgB8YptyG/E10RK1WbbQXOl5IaBLfcBM6a+cOiFF
Pg1a51IstFIsBIRtIMYPRACFCUcUWL56cTurg3DFyveJQU4VyrWL36eiB+okTXLE
CZh4v7SrjZtY3Dejpn8KZ5TwMgIJDd7GBVtT2YGdLWCWakfQM4FirSfs6Wixl6xV
6fGgaD9SbyIT5LAV5PP9S39Zgs6HKrQoPwJaUikPtH3vyl7L4wbzdv6gANvMIj+S
mLp7kaBGOfcbrfckW0EtUhdCYscjeSAmPXRsEAC7xNOzKuf+oTuMsS32ZFUW56E6
LcikpWRa+JoqXeo3FktTatHhpYqv8jims5E1Uw/Fe8XcaKWvZN7ySWUJPQry0WJd
6kzJ27Bl4DQ/5iY57jYuek+9fviIBAhfzxoDdNsPtvQtyPHw/Oyig/K/be47tnPe
6vYi7uIvsUJJHSlQBFlPTA2flxttZVXEY/KLgWu89j0ZR8jXPZJDVRSm+T9SPs+C
z9igk9Rf/ytXZG/IbVqGKIDXaPwun0E/eaBF0HVIt245eUnjCWm5BBtMbgiZrlBD
I9QZezW0jthVxutKTlNuYHqCWYMT+vGVg8Umf1nJMIH5PL1y19pCdv69GgIkavgw
ksIDXJaWfKBL0VItYi0H0XkDlbJ6PHSBq05NcUDIzD77uyGsuKO+ELWG68JxOjy+
na4w/o+CI/vF2Axg//H2teyY8i8aLCZUWCuH3mOtk/SaQgjtM2POiLPA5yVSxke3
sYyL3ciDSrvTbZsgFzzSaMcZgXIGwhRF6wsoc9Em5IES2wb+E+cYuRN0YC0a5EI2
q2qP/IWVVW7IVACLq4DseeKS7nsfQIdeAxA8cMgGQ0mDZQNWufeCOE74NTaTnsJO
7Q8pj74YyIJcCqp+usZkGYDGjTk6avFeMARdw1MQotjN0W6/Rm+Bkyio6Kgbm65g
E6RH+LowTVHf8BOn5qThx4QjlcIg7Ie1wCxSeqRzqcHZJW34nDtZaJVPCdwk5sG8
Psj4wRNYCdLgvEyZxHuisz8VJGMjf58vJT8pc/+G7vnCDl00oIMZyyciXrKNDdSp
HgBmTcIihL6+OmcZ96vkDkW2YHX1cWs456+V5zRdUQF6lC57b+S2Jw9mxccuQnma
ozfNSNqlmC00ekcQMVegiq9TgTfAmJoQ2jaSrXIwOQRaHzdPc4STPzPpwHxSs6+K
maaMwKx+wNu0ulGqjvd7xWldNLHDGgVV3DFY+Oj6WuTj0XAJr5/OU8rXj8vu3iWK
900JjRTiElGxDzjGInhOj8bbpu5fvTMqigbC5dSEgQfUIt+Dw7zbTgyS3pcguOTk
TysIRoAg1cLu+rOh4J0s20R+KrkJtJrfeeLnBAJ+Dk3RZDQVSGsN0OWkB564S/Dz
s8L5H3slizYZ92gjrpm8gYt2ilaW10SolMnOX76o/TweMrTAlDqpfUYDfDoQD59m
l3VAAdVpNvx1FqPdj5O2UEBzLJ97iWBIYBeaGtHhlvDVTmuvVARuzNCWKfYW8gRf
PJYw4Fw+e+vrJBFfq/4MfaEKdurz1H34UpJPXsz5QX1riPMQDQRV6bCPXfLsEuB1
20xBHQoXpYN52ARDya4aOvV3ZfRDDm6k6N8UYahwCUuS3mwS+sl/n4KmbTGVL48Z
ETTAmOHbMbHAP6xsjgZEe+93ncqgGeBzb9WP1y3UXQLuX8LCUCUNVrsvP0P+CxOy
9iVy0qPZ8l3NZoGhKEP87ArAMv1Y+Ima0v29OPeM53oN8Ldw6bmwIm6Uf37FuIaI
EWNST756aouOmB9DsbwgT7pUXJDsLqPdVcillp3C+QPnrqWvw14mAfjFUiS38fD+
33ezIdZQSLPTOGuPS3lF3Pc1hts++4GmuICTGI91Is9xARr7fqLqMaMu+dk3FDiT
JJEGWR1oNcL1bc8by8TIoVownUCyzf8Y9oMQASwiS//5/a3LXUF5ZYMqfKc8NzO5
olxnCm9O1v5Yv7tnNJLkVtgSy9/Z68PsljDfoamHYpHOWYaroXddpyrlr08siirG
l00rR/FQ0aBo1cfPQ6LVTh8uexaNVuEZ9P4+5qjtRCItCMngb3iYhwz5w+D1xVV/
TgSwnq1lrPmqT28XBh/XBSvctZyOmd2b+WbZeU90ffPBpcZcn3x4Jm5jEEZ1kSls
uPE/Deyjs/5zYdub2+tM8LCNjFH5RA7s0vHgimgVRIUKB8qUNyKJPXIdxl5ECJdl
Q5Q1wR0XDT6D3CeKpfOoveVox3QDrl8xV3hTHo1wBuQLhR1pZtTnQzxIqLiI1dgj
anTUpBwwzfJ33nPorNa0gYNPjDdSd0A8WF2bcO40U8/ssP49sIJhTzNScZlEWxx5
8Wttv+K5M1jVL6/jbxp8mQCFBZQ01btgIVvtX6X/s7Mg1Op5o4bDDw1HcGDVljxW
Nv8mRXuW7mKO4iYNcSVCgAvZlWkQgiIcVIQDtHY1KaRB5trtjQdRfFvpBfe/OAXL
q5lF6fTK1kbErb8sAWlMl3UPHkqBs6KHEAHUDVjkQkxhqhZvmer74+CrPbS7fdie
8Zm1FD061NUBtjAjqCqRdguNDWL+gp+XFqHyPPmNkRjEaEmOHJ/4GMFjgAC+MJDL
Xq8fKuHW8ttgPOJTFxoUMNp4AaX2ghaMWz+fAuM8D+7kTf5vIx8SSVyki3PzReAG
3mLQmgs9fJqOQk7xCXGI4O06TSWEGnwHl+eOOVUA5eYk+wkMCBsopf8hrocGgJK7
rx4B5jf3Ds99ERCc88NSv1FmRZLVsKUjXHnxoOib2HRXq7sqHORwpunUC82vBGIQ
l0qqVlN33tlLcMA7uNbBuK7wt54/XYWAQ7Bw78DI4NSjZwKQQFO6cOfRjWkOvhgd
fH7AmQrgcNjSfPI53rnV9L9hQSmFOIDcimMuqz+A9gXzhELV+dwy7zsHfsSIsU4p
oxR5Y6dOYgm/e6KJ39M5P6RoU3BrHBeVhaSuU2LKjXPt+LOKw84rZwYLjAE/0JFJ
e+djtHpXZUaohE53M99VAHKTJZOb8QpW8MNTfLxVZ4MpW/pS4aUgtRlLgnYzZXm0
tD8uzQCuTi9OHI7q4Ta9H916qRaEpKfodPwtE/9e0Nj6wMG9p797VU8ql0cPn4oB
jVtxcAqdR+zHpComKbiF5ps0RYK3xQURt7u5X47IFbss1+alEANAk59piP4AzoaL
tKlf2Hhn6BORGqrGnJCrfkXrmq/16foAT8EpqwP8XSLED6x+5H7kp3cTGtuAVK7r
8QU/DxpXZcs5nyoG0j8ljH2/22M8DjqVP4PCd3kAHKFqUYPKiZbErcHkU1M94hO7
+V9Ff0gIO9sfgC4OYc7nnH2wl4K9yPIMsZn7wkkJRV7C7xL6S6HRAYtDKVafvPBN
s0fQFlmHFwpEbR9uRu5fl7QKahmitp+xr2PhVszAP0X2Q8Dwx7S0O5txMyOiDR4y
N7uVfLneGUNeHYIY2oUpnr1hhMpMxfbWGzR7FxzNVdXbJSudsOgQrxCdmkzX+2Lc
/F2tsHVx45ANdaVNG3DBVEF2pgmAOhyeAxqFyfdmUFh+TvaAI+4Yq0ZpKW+ceF77
WFxpLtk7N9TSVYxPOMtBtdoARSyXPeBvfmT7XAtEo7uiBBNcGcxSohVEihi6bhg1
NsDgmlw9/+BxLgPHL3uJvbBjfwj0qohMD6jsMYNayexBeexMhMRvFZWBRsdPlWaO
Do0r3NO4S9Z3WbXv5bbG0XsmvlNVumbVLrmWD82hwCDfTB8+O38dodpsWbXfY+EO
tBoCLNGLTwjq7mN5ZVgRTe1HHIYtDNXBgsNU+SjOhVLhgdSNB+1yxWEVWRCm4f0A
vUiEdt9+pNXonuqt39b4z+p2YKZcm4XqedckpQ7XEi3b8W9tjKJx+sq4xBpN6E28
tMRHqUfeyBGRXtED8w/BoTaKUHN3vy0gDsyIdYMsQ1v586nCCiVDNftzzhXRuKWA
lBWRuDKqSKXaNlqWdcADZR3J6YkekR2JbLWq/kkGrq35wPrqozXFbHELDNsjBX4m
CWyw02/qafsjGUV2nzcdzkCJVwjbdxoSEDEivdxAYVYLGx9+o5f3DuNFSPjiuWN2
Ggv+4qCBujBeQNQq01qVnXI6q/JQ3iGZO67oZYZp7ip+BUMPWIq7VYlVvg3purOl
rPrc2+LCrocuOB5Rq1iSS6Zkq0QpifBLVOFByzhmZAYDCvK4hnFCScnt7BdWaeq3
vJ6l3eQlLX90P5n1qaIR7YEnvGONknoCkKV1WvgPnSBhvYeXu8FDRAmOAvvws+OQ
uPBKN2r4JHO8nMsuR7DsqtH+3WWdi6pXcDhz63XiVoLCUYi305UJUFmpZO/IZCoY
mhtl2CEDDEiG2jqEjZ4bqO7UfuO/7kQOJDqWqw+rTjNazI8yleMyy7yeso34NE1Z
Jyqj8x6PRKGlSNeVt1JoNRH5AlCqzokekq+Jd9L7r+nJlPckomFa5dehJuaUSti2
/2tEfrOOA4k4NQvya56phMiEL8Q5usMhtF3AkrvfC7yQgTYMmmS0tO1DprdwUpFg
YmcNheaJJkaRs7Xo6YoGREfXiuKtO+QPO1/nWmooHYuYo4sF5Fsscrp2VtZBCqsK
8DgoKvTFvUDT+EZpXRlqJvDVvPPkdLIHZz5+cA0lc/wmAO7acBXyKUG+XiL5klxX
YoUHs0LtwMXXIiSwQ5xO0S7RKtY767Q2vOJp0hwKOmbt8r74NJAC82LXI/ppTKAB
rmAwSXuj0RFcJxc/oNKuFlhV1gpcqJDFyCEh8dheKX8aMuZCdmA8ORlcmyGy82g2
BwTA0hq78GNQymxoeEokhJmwUqyesf2MXmOZG3aMmaz/0L+CgIkIgk84t6RT2Ich
HlY0LYQMkdj4v4B3ULYIZDC8+2r29pJPjHCWm7H2vk7ahqqZ11TDCoRGkWnDV4DJ
D+muLvI6hpZ8cznK+QJ05CtWebtVPBZIkgq3f/fl+S7pTGr71tecDvJdA1k6SP/Z
JIo8VngZcHU5yjtrep2ENArlFLmwHLaMUs4uU3am+Z+Mk13fkCH8vMl+NUAJYVAB
tH2ftTQklNOqoNUcxjng/0TZNXFxF2uIaRa7sICkbP4Isj5kbV5WctuONb1suklW
0K8mGMLjb47CW8dFQp7I+7NqZYfFE6UYzpwBC6aYMpPLpixNI0AePxZQiegQ2Byh
3uSUHaXlcEymtn48wOg3cfVR9itdEn8L2Ts3nHcozKJx48rY9i3PuT3W1Vdkr5Dw
hhveLkUOsLj3Zct+0NQpwJB3xc3EQbthbj9SFgb3slXksFD2ehk2pUGy5GDOGaw4
an11RgKT4J4XSZbcN3jG96hdH1Ep2Qh9k/sUV7VCoZy++ip7LwqiX9rJuoixJjmQ
ljx7+D211FEvXAXtjvZBDtCuEweYKdSyN43A224I4bjsQ3M4e1+obfP+UzthosE3
GUPN1/7VyRo9y2sTpBiuPftaYfwqoRE11HnoIQq4G19qaCUef8tBvf57Rm8D9iic
SP6dUhlovf/dr4qImTEBsiNOtu3S/lAM/GZRZDsGjOjAnqC9g0qO6s4ZLfc2Jhj9
TB/5SlToq7iYJdazsOW3iiUv6UYg3EWSpmI6Ky2no9S6+NFV2cCOza3kcKLsMojA
Z4b9M3pg08sQjJeXNntinBab1iGC7hzeqSV8NL7nt79HhNWqeZYqTpDy1HZqmw7f
wX/5vAyBeMyNyBvnYzoa9fYyAGNwuHYv5if2msnbZqO/yAszZIyxNf9JI8/LlDpV
PJ1/3ewDQ3HiTLBJK/6tRaF3kWrSM3N+Ihicifd9u0ai7IIcke5YqVu6LhWqP3Zs
poEXP4uHaQie9bzkYdMiljSm5t8SUM57M2bX6XUI3Sxd84dLip59MrFOkaVa1Vb3
F5sctiz2Z/DHIioHNz1P1rKQ+7pfH1zJz6/xKR9zy1FJ2/gUiUDe50MZITqCAJJo
YogNWV9Oy+C/KqTiZjVwpzlWCQ8vXhYlvKur+ImC8j6BU/PBPUNuLPl8DNMlAKUa
tnD9F9xX/k9NRXWxbN7hYhY6FJjew+6hoUlPbF9iUCdOhpLMbG+CcmztcUgfrXIh
p4PkR6g2ooUGurlVOkGjqeYDa8ViDuF8oH+qIhxygxuXqN5rJLdv7B09+wVXUtSl
cQYF0DiPvlen6PJVvvDXC9xzMm8zTVx8YOdQFRlQuoXd5V3dtxXwrHduzs9hwfMD
b+f9+KfUAjAEeCxf9xG6d0oTXx5JpNUJHAmYBn/KspisxmXzzoCYxvmGXcsIzCCy
H93heqDlwao9VpnamIXSpF7noY0jeYBNQP4tTNNkN39+Vm9uEK43cXlhQV+gkBuH
SNSoGfMHgZbfX97Am7we1UZDCMZyfmtc/rQ/gLBU/08cPzezsndHE8n6wGc4wkBO
PsPlr5i1fp7i4N8taK+dbY+gfwgt0XVhy1pRjTcPg1nXnmiDBemrmlN1qSUdbku9
S8cCCcuuw9E+myHpCCVN6+Kr/o2nKrtFckUFQd+vKRfzi91sFa1s5MdzoQ0S2LOD
1ATKt7R/Y+kFRxdm3vbLrX2I/sNVGDDkrF14bhZGx4YOgq3MlGGS342pww8rkkqy
ngDbw29X085jMBK/DFM9O2gK14wcs5tpbpQ3HXnlhlQDWZ3omznQqjDO5H83s8jK
IGW3wgLy8vdk7pbYNmX+KxvySctByZD/WSsDFPEg3BswruOJhHOsBHd1DfpD5QxW
j4iiouycluGw41kgsve3+PmwZrqH8NDiHKBEw2okpGR0Lv5oB8m7MGyStsYOJg+R
lilLXK9r8TBSNggFfdiV6x1wdXfamcsmoc0WWSlt70tZmGkX4kSajb6UzsJlUL+h
pJR9J2EUmg1uTVgdiYkUapA7OKI7rm68I55PlkGfkCssdN2snWpuX/+HqeIvLVnB
lh1gnTE2wGaoEL2GRuCleguwBAQKsyOVZmTK9/4ippxJj8MUfnWwYUuyiymW+MW/
IUJeOwu9xe1B4TVOjMOHimtxPA+EL9tGyDEfHxL5vDDdEpPDJnDban43kDge2bXt
i59sIbTJTVK93UY2n3B0hVKYrlgNMKwFiIVyG0WaOLPRNtI4W0PTE/ejsuCeqCvl
XQf3pqK/mKzZVazUXYHY8lBcZm06hr1UsmBkkYpY+yaD/KNU156+bP8EvTlin8PR
9dk4UDMQnDUjoAXFGxYX6tE6KuSD3RoNgMh5GKwhwLcBZPYfofBh9+lUgKo8MN4q
GDkyHaQLejmKhmPMsbL+jf9ISUN65R8748sYqwfL0baWp5DdWXk2oGefE+o3CPHM
WCY1BjY7BfRApGW5Rzqlu8QneP0Q8V2aA0Y6zg1e1zglGlqRnWENLu/WlXmv7+4p
QL9BdiW+3JSFvgY37dxdZjG73k3tWFjGNKiDSR43hwuEnysvQuaUc3k87hR38pAF
Y0S71NEIdb2ySCCa2lVB9tfvrtbuLZTihzvpsmceFQE/U+oD4jIP0YSGtG0MSquk
6f9h+YPxjkaI4l+xmgPPazm0W3X7Ohy+wWwjSbZUcrX+w/zbDyM+knZXKsnU9tGo
uD5sQyJjVmX4N5ZJjW6hPpCvmU/QigVKKguyV9BxKgyC9T6vUIHpqhLzWt0AAn8M
FMowhQ7S6kQbSz2W+oZDpxZkGrZr4ElXtXlwz9oTxPml6iIMAgBUFlU6RF4gJJ6A
tyis0KyA9l+2eDUQGBaGj6+BicK4W/gJWfAuU/lzUQbHpTb6ZZXEdizGPBWEyTDT
Gj7gkimksmm/RBhnmuvMPLS3rJ8GH37WEysypVFQjnr42cQMRFaHjTGN+b4zNAdj
MAvfDOBiyH8uXlAOqpwEBXB9N2NrftwfRHQOIQnH/HaBeleyQuE6i/Fsvpvr6j/l
drTj06x/Kf2H4qn/dkfqP0qeDqK2QGSUI0jABybNsgAEoNLOPCEvd8Q33nyRShmQ
U6dT1mkjSaY1YKJyOaVa/b7A+oI35NZ67ANJIuEFpV04rlegxkuJ4F7E3fQsthcl
XLqv/BRodOlqFC+iIJI3BAgPhxbfzQzZmt+en7E0KYadsi/VLcxekvXYmXJlIzoE
rNQUb/cEHNNbJlQF85knUuppommmgVm0c4F95G50+/CnxQSvdjtbH7SYfDk6IBbN
i+hU10AaHpktCCtywApGin3xitbdaUsjBYxew3uKhXTjLBfjPCWah2+IRVHrj7GB
w5pYxgfPWUplh12ocq4UC6yQbPKG0XiV1wROHGilXxMTdNsyc0Dp8vkPSVqiy/8y
qiYvRrhxTEDGhVD0dVC6PEV3RriRANQ188jyMvJE8ZQ=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Zcv07OBA9KDlEjhRzh9czuKeg9YhWyCyWYpm4gZv4x+iDyOlWvIoWhEuw8kIAe3B
f7Ps/7bs37ksVgkcDgX7dDjpHObJa6jMeqDqd8xqCrNc37ZHU+fOQBAEZqC3yX8Q
HhBC4bo4LExyxZxadW6TyvaqTV13FWvqTTFq7YKrFK8AnN9ox9NkI57zErB5sZPa
H2UWHyeHZs3+kNZXKWxxMc+eVO0HM6ey8fZeluRbDhQrJLoTpG4oBlHYwu6Q+ta8
WBYV+TLuVDpSNnSD004v6uvAeq6RaWYpMUAuIs+uI2MtdKudTpZidWE/pWSXPYbw
Gzda38Jj9wHkHZMb+M38fA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7632 )
`pragma protect data_block
/Aphog5ZRnYOtv33OW00YjsfQqRleyUrluyQIUlHtGkHuE3JEbzw3QGIkdlCuJK7
aJD9oBIaYvTf4hxc2LIeM+IuT0+lsQGLepDaWZ0sIZdvL01+mudMqqVn6IRsVa/y
BI6FVtQwKF3eorzwKp5W+2NjnOZUmnKUZYo2hD1jKUUxCXq03Vz/WumT32d2Ekoj
WT3OJY/7mulCvvFIfWqnak9E/YoBnUtxfXHMONc7ckz89xMwDPOP5Znu+wJsP+Xm
DwENYjsF0dRPIVhhMJIIyKhBsVQS9M6xeKA4ut2Muh6KXNjQXerpFUlteel8vbGd
1gSZMmCr6GMvKtyxaQxm4Fi2emxgl+c3FJLvuwMjIgD4xyvrtOiQ/I/Jpw+rgIxv
o47rtNlcit3EnmFgj8+BsIQuBLBZXRrRxJc0i7YDz6vjn6zdfFo/6OBYrag46NS/
D3UBhfzqwBhxVwBgeV9dFtquyz5ngeZtt8acHnqKMyaSzBGZWnHT130wT3Oxwm9t
MRmWVdyYawyO3bc4YAGHwXHdUvNHKMIkRwVX2w7a6NZFJ7RR+vpHcnsfPMBWU90d
IrRAw/BUnguWi8an0FQNGwNTb+xdq/X3NgwmMfcJHZ6kaNDj024C9b6AWfgywVEJ
lHYNC294DmMsvC1lAwejzANViD6Fn+7SeAPygDx0BDDWGHqH8GSpV6Km8yZBco/o
RAuyGhQyCh5ygypnJFXpqw6esOI0HntWM/R/0kXzlfyDX/Ru/XceuuhkD4zBcWcp
FDOVZfnuR29AO4t2RloV+lL6A56CBEgify9KWzkDGAP5by6DJvqWiJ0C/HBiGJHN
Jeu5YqJDHgAJjGjpr9fdiuDXDfjk4/YFAqOjAoXNehBFZj31SY2NQIMLNtBzlw7X
XIfj34mmm5kE4mVdlTwtAD2DSq7ZFv+ciSZ25Fv0KxLq//MhaEJhO035CwHY287T
tv1T/DzVGGNMGuSIKahf90XFF1VIQsxJJV4AMAaeIgVOPE/gAE3B6M5jPDHOSJJA
s/bO3T7VBRe9zvwwOUnpg/IGkHKg+JTrvB++A3burNzvKolWSTuZfI2Ly9kNK+Mc
oIMDxluYdzvn1c0XWf+VCNuxIwMaGb9Aa5GMUypDxD2ut9iiQ0+Kti0c/eiEFfRJ
IP2vY3Jcflf7XdgmF7NNhxT6QBRljVHNYerItqXeJ4h9w3o9RA4cNgaN3FAsmwV7
B6GHnqE80VxKF5HBiGg3+Jt4tHt1BO3Au8mEO3G89WRwc8RaWc7rpgfQvBIv+R4a
9FJc+gnLim3oCJzi9+v4gH/iI02X8Ahj5bLkovGtT5fUWry51fxd8Mwo7ws4Yqr8
TFP+5zTpZ3fsUl89/IDtrgGTk2F0N81yAr+TGB0paBuTW8CeOXjTGlzuwjEWpneK
Q0yvs3bPyZY7MrPX5DeBJ50eEQfR91zK/q/2Py+9esyW8KegPuNxL9gMywcYf8UN
YMFHBG2FVR0MMv6nhgHa3GuPPPg6U1bre1R9to3M9ISF55QcJB3gh9YEfa+KwYF/
PLsBgR4Xw/dcLmd2Y1JrMGKVfAQN0nFXU647EZ4JVmJpE+AzJ+Mi/3RcDClNgjhv
dYkHFU6pflL7fc6EuMUehNI4yBlziXAJ5if2gFgNQueHNXMBurszT+eKQPzPOs5U
E1/Lmo3grhMvCLjSo8aVOL7PrSTOrsbybhssmlWaQhHTRs3/rg70lbHXV9lxtMpp
axrFaNiE2ROOWOLkS/e883+zz95kILz7MXnGljydAVnGZ0jzTKG5YWZSsM0nmNU0
vQ+1YNTZhWb68gNiBbeR1NHQ2KLQR0wa1PT/fQ2OX0YLr7Dtzi+wZAMk/s4a3QKK
au9nLxAd5YOmjXsUqF6O6Vto3AWkc2jy9bIkikR7/0IweQnY+4Jg+zoS5Gw8OgbG
zOp2pzAeKvzfHjJWj1UmYCKLuNNe0rcCXFuObFXpb7Gmhej2TSjULfAwBVslT35v
HkrBliPsklgbUjAcJE/+kGLjIO+sV7LNNEcRXWy6lNKAJtYbeLmST6nq+/m5lZ+/
h+GLG4L6QsUBvFNvXyGbPe3r5OSrLHzwkLXOfyQm+EKHK0M5LZmOJS4pNSmowSyL
aTkO3Y15+idBIwMvKFxhL5X2dY3I2zY8rE+RMOw4O6YWZHXfSeSPy24r3z2eN4qm
Y3roajgVcKmSkIPZ8M/JJOnTqIQggqHphZ8ESQ/l2T+duyFuvTVwXN01P/se8vfo
nR8Xqo1BY9qx8y9+PHVrXOcLzBOAsKPctU11reH1Hnsj7A9C6/oPifHyeN6BnBRP
n+JWDP5ik5TXJTgTALUovzirWjQHOlJp4u4BqXSW6L3YWHL8bcM+H+R+M2bqiaTI
gdNjFfklbgcwKI6G/pCH+3i6CbcGKymGlJjEEAaKEuSwDCfJmgc1GVSfx+heCJvj
e7zrYDbD2N7fLeXyWbicT9vnIyUvkLOM/5lXt6h9MvE208u8yY/Krt3LZkAqfRp7
FZMQmgksjg8lZHRmpYdohVdEDM4aIM0qsvo/2yk3EAb7OMcn0BvoXeeN4XvE+PUG
6GgGnVEAZBs2NJMTdwQj5asmqR+6kIdjksJEPETp1TjGKk4Ocal1kQ8ibgvW7Ep7
wcWSw8wVcsuu14xynTHIqbxoNqL6Vl59Fekss3XBp+QMXRWTcU2i2uUVuT6poRgP
ZDePviYmhhaD6IZGs5fCXPsiFzSTBp3kS5WJKuIuP5Fdlmch3lP1y93NMQED7oES
yj/NWJp8i6HYwaxZjF/Ub9PTlnp+wJhPzzi5kPhYFrdeYAqZeFMlc/WSC6cK1Wvw
7s37bFAGek05QLaySopMQ3JOBPjJtZf2G0bFemDiDUYG8TFcvtVt67/T8h90neMy
PpHhR8Qb863Q/bxWyffUIIxfF9I+cv75ZeSBBcIx98+W6ONdVOUoM4z5MObn+ZJK
pYywm+swjFGOSW6xSVrAqQFqQEnItVdQH4AaikhM+bf4q4D++GUstScoGnQ8lfB2
bQ+WGapEPkPjSx2BpFGHwYpLy3BLK+1WBR6Anmw+GzTMIKZtGDRG2fq7PWw0nxWH
t4cSekT8dspQCsyZ9noE/UrZRDlOGaCUJEAFR0kSRvenwgpvpjchQNx0U048ZRrI
rvXXMYSK3K4x0Nvbv03MsCXU/3SV9sE91j+/yCMh7yFg76AM/H/xSaQ1U9c15p5n
u41EjPIqIKIEPclN7OxE5zqvOVZgMydhTsHuQ8RWpbXbmD6gtAQP9YkswsE2eUy9
zln7hs6QloCW8n0J7tk70ZEmIvTwleiTNK6mjbFN74R5pIMCwSp6fGVYZavKHJBw
KMYeupz0JVsXdDvp0RTf+wpEi14GfLJa5v984C531XN0QJgMv8yOBEJ+pn2CJKYk
G9ebA06HA/mEI+6MCJLlcaSjLw2A/CGGn85OsIrJneUE2dG1jfdRJZqgbgB3PuD1
B8dEflFBvy/tfu2+JikIQhE6XQkV3+UC6WR2gIceKlsjUFVHKYi/jLjjRY5PVow0
E/50WkaqyqYZKg9I2YmzQH8JEKa3mVSw3t1VMoz26QWbF/0zIHNHtpXNWbqAZg0M
XwBQl5kPrJkoiAKpb8LJrahTFn/DU24zIPWKGFjBnJcJM9lhjeQnaewsTtC3jM1D
bc4EKXR2MnB95eQ0XOANkr/jDKOq6WkPX9XzL+EJ3u3UsYYiwWbkhQFLBEerFj37
bnQPrFnk/CI054dlQQrEJzpJH7Khl+N1at0hmgsYnuC09JohY38u1FrHAeZARxX/
qKESrTFAFa4TXKO6mApLYCa0WkzXyKGkFzlKr2b5lmYaeZYUS+UHR9wXyMgkES5D
CANI+6N93SJQX0uXJRNxvIygHuTuy+70qYXk2iyXy+QRODbTMbVRtZkzsY+g+opj
az2Tq6zvSaPRdIXUoQ59/Z2f/hup8RygwrgfBpFaCs6sAInixm37g0fhgANth/Iu
dWpDsT5ErSDfBEc8POmG/v5rQTmqUSNd5i6hMU5hceAtlO5LH2xs5OsEk+QT46jo
4iaWbpGjQFJ9olcNcUc5GjphwOCWoIvoEpclDVfpFbTDQ/O5eJ7cbyui5mzO9NuB
tUKtgLY5hp6z9ALIdTnVM/DQV119BbKXMrPwK/A0lN1PWUhUOFuwXwpX9usjol5n
0cjV4RppGaA3LT5fU82XWNjsj9djYiSXMtNhykIrok8M9rgJms8e/Yxu3s2/3BKX
Jr5hfsJ31fqmmCmzWASgrewsXbFZtP7ufiYyMHZt5LGQyenHFzH47o8V32ElEzDj
naQixdA8OaK8I99y6cyg0m7ws8J2Dz/drG7KMw2B1xnCbVixWghJl+qKAAzuOeVr
optdaPQecXY3YroH/rUshulNdGISyj+2aSiG6/5NTKl1Kth1z+Z6YvcLeV9Kf+Dv
r6zanvVgx+gGQNGbVBrCF1a0oYZP4iGcx0+jtGFnqAOrwbZ6zpjp176VhbZCnUyq
4gQ12zzR5G8OdqBWoUKM0qI/EcY+DVBZZ25F/Vz7gkGVqGlGeia9wh35ubZBu8rI
dDRx9hAVKCbxgZAR3Gyxh19eTHIihu/vrqHyAH9F6afAlc2kqRI0hb8J33kt1vg1
695p/SWswT9s8jKaKnMky32xhJrN+idPaUYxCaNjuyeBjPOeCiRgBeAiC6cQbPnh
xhKluF8mLRjsuGG8WMBmRY6EjAn4JWORg/eryZQvdKIgvITg/7l8m4T9dunlz/6e
ovHcKPmXFTGQu3XOBJQZZzSlFkt0GX25//JpwI/hUdGfAoY2vwFFz7EcsuzdRp2g
Qr+PJFytTsY7g8E8PI5QdYd8mHwFe5UdocyZlWipRtxK9huGtgdmtsmRWPcJyl0j
fty2mZUZyLskk5d0okoxMMsMsD93bdDMM9U9Dy+ODLGIYILSeqmOFD3XvnO2yURH
uG8upuLwUAOsrUYw9rbPrt2UH5OFTIfmjKAyx8OkE1/SQ0oR+NJ/hnjZkBHHAOQe
S25usDG8k2NdaI06JhOK+6pSZT+eB4o0R6PizaaA681v25C75Z50jmyBVRObxFpz
7Q4jwnFxusV8yihQneurZD3UK4WuAi6FuLkzdbOeY2iqA0fU3kKGrK5WSzGjfmB+
wpVdOjpTA6eigvWUGwjiwx3eZwgTc825PyDQvFm/77QL6utU2UXWFkx5uAQgQZGS
sEIruYrfo5knem1r8Cz5NaUO6YQFY8WtA8OGPfPEczsqCCSdmy1mYvdO9awJ1ZFV
zeQ0D4BucpQtkOgfohaIpGH50U+oc8xcKsjhIakLdaJwVRiduNTHNMWEvG40VkYr
HKuhsHwujdP5V9aylehyvvJNKYIXYvsa5XZsnQ4OtsTGiQLbXfyNPQ+sLoycFFNf
9HgvtErgtl+Dgjo1l6l0vG92Z449LgaUhuOs6XTe6VnzkvClqlAPVtII6elUn54X
SuoC46A/ip+wYjhdXr1a93S5MJdJpMS+XT/GwA7Um0fyRC7kxeBV65tr2i5U9Ty6
vcX85o3Iwb/1eLUoOmbHRME96XnvyMGX7+nzZSNLHITSIH5V6pLK389oO+a1MVKv
dr591yPRynYln28D6xiJUfzOeos6hYcXVYG212l9fTpj0V2NxZIfFrLKTWgmtEhq
Mrb5jjuKcBR88v1A+RR0Vc9MbdXYBoTf9uA71dOPjqsYBPijBccxxQXXsf4FPPeZ
wgTl86tZAwvT82USGqlhHXiKligjxvM8OOWToPlI21799qpmCfGT/Zl23cpKdZbx
YMRELkTvl06XSIhalYRbHvt2nKitE8MB+3eqRDdPB6n36dvhwj6yrsXf+Aw2qzOX
HQCcQErQ18jK/KmWiw5G+BiSxAavOQDYbgEZjIdsEJiWdSOUwegvvF3NVuuRzQd8
myQiEkwv+wXKJyhAHglGnQ8XK6fo3K3R4YwGZobAp5W43qtMtKTIFGymWB5enQaK
HAG0vlqD/6tBpiJUR+o1blOv594r0AHP4Q7UjN1i2cU1zS0ftbnwYSwkdMkeIwrH
L29guLvOHLPHYooSs90T7Ij4aFQOqAGwvXJRd3HDGDyKYxzg2ULyub7ZbhtR/4XJ
2xYJ0UMMt0/dcRJ9q+zTfjoAHsxYZE/2voYxCkC+P3UYoWAmBOzDypUctHBowL0i
gZu2YibZQywVxF7yNbBx6yxEehP4rTEtb0D0OJbd85zt+pUUTGpwCDtEczhBjTsm
helC8dds8+POYEnZgxkDEYC4/u1CtZZC8RU+L3sMxXEGiK1td3jYuqKpM3p51cL/
iZJD+o6f0rzOoN1fiDtKG56SGYv8C5m8HqDyOcZ5Ou3wgL4H5v/fzCGyWgFzRr2b
sYOdZ7FsrrPPyQxJ2fCS3txiPydAf87YKq2zaDnEk11Hm/so0zmUx3Vq02POMqDH
ybU7n+1cLsyDl+EKQL3JbnYSRqs+XWcT9J1CNHSLRxorrrekrS6zCychHKuZjRTC
eenRfgLUF1mIzLza3eyylSbmpAaW/VSAes/A2eh14tVgv3EJvJy6m5uuTbPHrxhT
fufHUtDAFfi4/5Z6wfj5WpcQ2eKiPibkn1HzbTQWDngLEa4bzPCxlcx6Pk6lA7jY
HDJEOy/yxS5Qca57s1IWEe3EWE0CekVkqJhhNGJ3E9/pE2gyKlqz6OVmp6QCjCgn
QMqFaUwyhV0rIVr/gIZckAd/o9zD+aUV/GP7o+t2gTd7Zv2JIvhVd2NRbeWG3PJI
iTm/wXsi8XYQmocfnA42KeDrtowP2S+KxXvbuwTZOWcTE8Wev3L1F1h0eqykk/jq
onx4s2WX9dxuq/RNG3W0vh4d6rx2rhH4xJB7oFOUPpdbMToQa3+ms6Rd4SpVb96o
XXUQJX080ZF8ttfh+MviLzsZ+Z9sZ6I3dCa2lFg7dQwRqnlmpjtKT6ZBHWJTcIb9
Gt0EKCwDVtgVv25oc5Py6XRxRJ8uLyMI9LnICZjipzPSxSi4xmxc5LiEM+0CWQ4N
M7PHFOkP5SMMIbFYIbW3i6mW4G5hmIe+UHqDa4+RjOBCISmHlNzAl3AnEZQtKTis
AtWP5Endn+/tVRUp5XZbcn4Y1RF4GpvNC79xSmYNLDudwQenjSLZBzwgDvFLF3rZ
Z9hh+HI5tlGztPC7MK0/i6o/LRq6Xn8TTb+7X9qTz6MTNdy+cS9GRM6R3oMLDN74
C+bbq4vZt1D7h1Gd3QSyv2sYbiZVtEiHGF0fVy9lC6Wmf263WRNFDg9Pr6l04D4N
iGZbh27TOwF8PxbmMfBSXs96zCxZqot2xZFw26d2gn5TctGfPf9by3c+Gse9wdHp
eprx5NZLpGUhmwN88wGW7G0wjC6ENlp/hT3CSpFGP2xQpdEWWcAuy/WsfAV/dRGK
VD9DI0LaWjV4xtilgpHAnIiVaY8T1qBEgjAOkCW9moXJDQld7v93MMXewX8rsEZi
xmWDyPhr8z5l5gDMYfibNwIwB0La9/8EMih3oq2DOnXkHy8XOdb6LOs5Af6wXtJr
Orw8fCOyIdymh+A9Vyh/qv123+rTXiwhzrZBNIl9IIh91aG59aSf2iLlSQx3BZBp
CHe3RvrXo85fuvkpUyZCBlfGe9TG9yHWZ3/G4VQxxFqPhfvPK4lOLLT5TmSRTPE3
m4duD79Tl1wwQidYXwguRAxSvXtxhlkKfXt92lpD44+1NPHT7IREJZXRIVJClANA
la5NKTGEkWrlb9K3nfcwBSm+39OAZ3RXvayuHo7SVkSK0QUyuyX5BtPIe2p+dbUq
CdhWGaCInCvMFM19hEFWS0ocotbl2nHaUkTcMGhz8vrQp3kbK0CBOyReHtreMxVj
mKkZzpPTVzHZPaPx0T4xq289y5/yGBncKWgur12vHPpLge4iVgoNUx1TeZ5eEcqo
K4qi+tArHz9Fis53JITQHtgpHpWF9Yj9IMQKZJ+3PV438N/admNdzEQgh+iELa9a
D/uQzKwrKCiC1VoyX0cT49BpiQMUl0/v/TPCIxQMb+B+OgdzqQ9cEL3nf27V+MoO
RMsTvLq5pzLEC44ndIHSJfnSErNmrcAH2CWanDwVWB2PhziP6ytIgnZ2ygpCbaIk
qvR4XWMWyg7zDoKeb5l8G9xST1nMFwZgKVnBvc9BuC463T9iW00zw+T/iLQVgrZZ
yoREPKbW3UU5QVYskLuXUWhaJLripXqE7F3sCN00bgzVEo5V/9rIPhc/M0tjZZmA
3K1q+/LNIbegoh59Xk03ygGLC2so2YpKgACOjhjO8gbkh/WvyPqbkI4kpxXYO4gd
eYnBR4/++sBa846NLBwBBFdHr/neNm2EZ7cnPoh4wXd6yo6Yu16moV2kbJ+FrbU3
gDUJRA3Hkq+dP2slYLi0WiqtRUEMyb8QzW2oIEaa9BNY536qyN5ODhAxwKgNjFru
ammh6Qd0mpSsLPGadZtvBVUFAqhVusmRwYGgvIVCKKMB6X48i+/M8JSfeTkuCLn/
CMYvj74tBW6Gg/hL6zGeS6n7gcU8fVH2ZWmuUuJ4nywaefuBR7IUdPRUoY2HcI9X
w9IWbTz0k/ICrpdhnvx+1bEVsYtJxS9ywiIp8mInypzX14Uh9iKi4s9A6l67Io6x
W0nPm8nfXQu+WNvuCZ1xsFYZsHbP/3ByM9mSjqIBJZPl8FeZCqmZRWXpB5jDBKjg
tkDccsMf01LgRWDMF+d2r37DRCijUTf6fclDS7wzTgc+FJpXjT1bdg+qJ+iPzP3P
x4bv8IsQJ5Sdyt2b4Etva/Rir2n+ifgfDWp1XVPfVQJEsXwSvEsPLRWqOjA5JDdA
syIb5RDK1dBuenPPkwvr9LqQUYJ3IKc7732Ws/F83E7/JZr4oDwhWtRi8SmfJEsG
n5kQUuLEWUZt2GbxwSVGfkemudeMT1QKi3NpOIIx1cdI2hqHWqD0q0lqS6QR0WiW
1wjVf66T8eTeOEFd6p/qacypwqb0f8dH7fFf9XNUMRW0sywEbTAv01AC7R4cHdya
MJkKIxFb2ggrbfZAMIeAIS0aOxt52x8MkwtAa2z47/BgjO+gsxjSdoTNETZBEswi
w/oxugWQdhLLxcz34cHixhkGUAi5Baz5q0l3KT7RbWXTeNDbN9sn8dv+lO7TBqgn
S4TbOQyQm5ztcSMpelbLQJHFhUpNJJl6CkM2R8UPoUWiFdkh13vhKTYgsMY1pFgE
pmftoDKujAKQyTZNAbP90cFrBvy4jveAydH+MS+pRiank8ourk61xj8LABOxVJpy
2F5wMqzc2FgjORDGy5PSNdjMA11xSTc2jxzaBOmom/A7P95xlGamolzWajoY9pKD
4pVCehv17tbiiKY5fScQw+0pErYy5QhogUa63Fh+gkS7F1ewDoTcFMHqwGQHaOeE
nZWmsiI/N9wuD39rrbrWRgCmhGhx6v4y+1a8sucitEjIhGc2bOCkeKXjAR1x9oRI
rFHrZDZ8XQzqHmIoP2ZteJdOjA3kxILwJ0Z75jjaGSM2gZAUoJcIJfhaGPljD17M
uTgUTnqLsg2hTV3+BeOf6odFj8PjFl7F30PRVhn1Zp8ZZHh4/eS4YCswFwmQVgPi
5X55pK802vLmcSHEO3rEgnl3pSlVOi02ctxlKZUjHn9wvxgfwf5uIVbWc8N73Ijz
SVBEWer8QFRgN1HLHr/U5lOnT9gbi34YKWDcYnAZD5yVotQ8C8lGHHjNr53Hl+Xm
M1+LUSYhGhU1sM8+8USI+ES++1adRMqqHvUp2NYmIGXaqQuz1vjzT8/EICWOBEUS
rsB7nkImYwDCMBbQTnOUlpASZUIo1w6Fs/GOR9/3/m6FCc4TddYzGIy01bg/1+3n
dfqlub7dvs07ZJFf6UCLput2igJHh0vZA6Ds9L6QykslfGQxx7CxgHAY8U9xuUhL
h6XLT0jrGBVumku6y17MwCN/TANIocxBpRdTXwY+l3GzpRuPLrLG39ICxRYQFXfr
IrsZIqeQVH8q5TpJRgxJjbgtMTurKumQUFg9uIQDUKQ14RfNe2YLZ8y2O1ixyzdl
Vur1k75j3MIV4jhRZnvYa0ugAz43Or4yZSDrxH6YvN9vp6Pbkb+HcRwUfFjFpRX+
Dz3KZdQqlls4Ybq6dUPEM6l0zm1b7+3yiT/8XdXDtYeJr1FfawYQn10eEtIQ+R1Y
jKiJfrMeEt3Tv5FuDQ7zF3VoPg0DM7FcPnaGlv5++12YB0H2nA32UiUZK7q20NMn
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VDsLADZa3GAUGe5SW2qiDpugBw+sZMg7e9dnzQKl9p27OsLZ4r9O/aC8FOzE0LHS
DlI4Uho6gqyw7RR4m4M6EBtTj8IZVgeUOFV7tAe66ND8bKAMQYHDO1WDaBZeqyDf
pk5MAt7arFCe+a8Stj7JzWqIa8BQWgk1ctSvRrUzMdARE44v7qDaF+o3HnF76tlr
5QPU8V9EUSwmLeOKnY5g5buBUpm9qZDry0nWX4+qjLUeovMOAdgCw/QhehelSD1i
MJ02Y9HSMKbj2r6hdoF7xLDRZt1F2fWqSko8yNgdm5ayJ8PMsHhxO66rHizIzPQr
qP42cHLft6W0cdxYbG3qjg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4768 )
`pragma protect data_block
3BkNK7630wx+4qyqRSDAvRK7mFV8oD36+nfMhWlGdarhI+Dsemh69GmBk9pcBRCs
t+bBNWMle5JbAEY8jWORbMQiElq4Tia5cEQ7CjfLCF6dWJk/AglQ5Cdz5gGz8GBE
qMXrTT1CUEmp3qqwTBIBNtCeQ+TpwH0l9jtBe88SBKohob88TqG7fpROJJxaGk99
KkVel5E1MZZdBlwVv4fgptTWhWKmI8zLF5BbK4GY4wrH1Htvz1J2VPq6HA/ukeqc
HOka+5cuycUrVhDW02jsZAY0Y7D/M0d6+gH8hJ8WeeiE+ftjwhFKkrv3GM2yBzTq
UOZJloK2gUnOfcq2xoW09AVisSlQ1TjbrP39n6w2YSkEaKDtb4YmjdacNv82Ncm+
CAKC5D4L6qC4uzBHtujD38Cs9tsvTJD4HAG8VRWdJNXhu9Yr7tIEDpVmD6iI7u84
ZLNV9T7xQRCcakDfeLSZeGaOA46I7TQip9hFz1v4SOj+eaQNAEHtYzqB7Ih/r7kp
S2zsomq3J7P8kN7dv8I+5r0EvNCg2IXbw77ypLq7jPVR59so9Ml2xBpYZ6hBKu7d
Dfa5JiqXa/dBDGbY5wOaAIRDC6UMGPCWUrggESCXc4MrGL4tXhfY1bzsZWoTrFKm
Ldr7QxlCW979aMtl5evNSDQARF27dBcTTJXR8ihSC8dlXZXLzKu6B4V65JcUpQqH
wv0E7OEqRYwrYV/iOBZUMbsbgaMJK5SIP/8Dozb7WmwR9c2JFnU0sBBDj09MGm+l
J1bTN/TNKM+cb0iNcjPmPZg2kKuMLi4X00m1gv3K0lw3GzwHNuJ72soSlNuHh4bf
7/VvNUd1YH/jTvtp0UUD5n/2eR027XJ9ynWfVFCOc4UpMluXe8JQuMCzW1l+MNfw
7vy0M4Da+nUkOLY+KdCsv1YR4FrE1U3KtJE7n83KzZnQQzHQOUtrNfhU7KebOARV
cMOb63B6QxVdrzOC+RQdD55bA6ZfEJgdIPLPv+cswNu3Wt0w6WNks9KZ8WF3CBwg
aVYDD3MoX8sKF/ERESAzWW60I7XgSIzvNjteDW0vHCzqoRM7hWouruFYodsg9J+L
VtunZT6a9rFFdXHN7dACHgKEhqFmuTnHD3zlQjAKj0UU4ouffKReRRY3H6Y0Neo4
7QtgQ5dJfXRCE1JBPrykdHiDMonyJfzHYDCNTKrjz+cQ9wnCAoepuf/6+3y1PVD3
aSG+J+eSC3RDR5fjb2+2N26eCPM/KPYRJ+h3QouL0OUQJNCyV8UeuTIxBoHGp7g/
xha319kqGGV3ck55qYkczV3TQl+zzhvUhMA1JOeCrB95s3PqqPwsQdQwqQVs4+gS
U/hOziw6AQvlWRY2Zi3SZPQfoc2wwtQQ8yTVjvyr+fyuCk5r4+ZDVzRCQW97aOb+
fPKE2jRXGavKKqSQr28PVppGHvDbysJnT/H7b4nln9XAaXTAubA4+CbYyjTIC714
f2458Cfl87dZF0FsdcEl/zRnsQFwW1z25X4hqxQGTHjHp70sAUiUKqfZFNFK+l6Q
Gq8A0pJJLJbA63ELQu9ZqumuDTVtkjueuW7G6ls+HKis79aFJXNV/otVwPFas4tk
E7M4Lo0rEyh1vzIitanK5dkxpzLCnydyGsh0Ce+gj8BUBWhrjiYzAOP4ybZ/vYEF
Zs58w7PvNPAFLxdroZipYswEO31XwhYyCTchcIWp+ylGNjTsT0j594emJ5STIFnA
viRHFcRhQ9e0s3poMWTKoFlsjrSOjjHIaaWbyxim++vpj3plBbCOXD31HCre6E7C
8daFFlrjN/MU6PyhpobEFEzVgIYTS59vpIPcYRHjmAckAzAsHWIqSRfi/IpyaHlL
vkD0TmCw6HVEEiMkIL/xN4MdeE5RQLQjx/kU+eNT9uN+TgbiAVe7CtSa6rQgdY25
ouNKg+uYC4Rty41hpJCH+LvvoRYh4Bf6EGsXxeAjF/Ki6wqg9z3/WD2w7vgIFXLg
qh9JSunBYGEPWfUm13P3bonr7gorkxyVPchOnUNGSIsQKFJCdcO5CfzFpEP2Ysvj
WbfKmBsxAA3nbe4/cCZMeRuSVXTGhOYnD26wAVf/ztjVkwegW9q3RON+ePIDK34d
ufMAU859xArtdf8pD8TRYogO7Z2LEhBkAb6XXTgRI+H0l8TYhByKh9fzNvzJFxl7
/fhQ0IEhz7i+62H3mYOA4sL8a4dpV5xkPwmpEhcO+wbe1ENEOHDJrjdSMUqHabmK
LdR6I6n0IjpMmUlr5bWBwPRgIllmUrlCEWNCOROt/VfdVxyHFOnoNPfJTuHN8K+w
HHtPMzcIVn9rC6TzTHZTMCDkhuwZaf936VHQSwy2sakpEBImoNC7WClo8VF/bTgu
hdTI+d+zTxvkumZP1QcpKCQrreElESTkcfBg/bO0d8CJYILfRLJ6P7dIG081dQS2
XEt7P/DYHyFoPF2HndjhK24LnsPMs0I41nCsJ06ZOwqZg/7+eOaFcV1nuVmMGV+j
PnFswBDxd9dH9LCdEn3pX0AOqQ9qrgvCZLoPzXTYI8xLkw5Qd4T71KyhsQdvFprx
vUCNlcEs0df1CfKC8ZCJWiOSv52PUAp0+Q2Ohzytlfy3/sG00KNq6w3na3GQxQ+k
u1PejtBxHNJKXHhI/pkFV1yF2Z3yhMA0QwZUP6zUm6sSbg6xxGQEKihaLhecdapw
pSbVC7TxQtArCp97T6U9hP+kTFOImjQ7Mc9P0DgOUOMNW/bIPaKx8jpnQI/4iLyN
c0QufeMvhFT+oU6KjILpCDmr4rGBq3AKOD4X07ScgL4RSQ5cpOkw0Kt7oye7dYm2
dK23Ia5Bc03YosD/X/i+gDAtdEUrpYDurUs2ulM9KfylieUCAvbsqfnYql17ro4+
mtxtvkWPM5UAa4c86fBPjFby49cZImV02iu4zeT0QerRqxF889Ae89XWaJ/9c5ub
5WqcoW6W/br9yGwFdrJyv7UGuaXxvxdLSDOeRckjgIJNg+0KFQXI12XQIbt8kwJG
LNwHcYfj7UvtFOkhEcGZaBaXS9uwowBy2gkADHfNdsrt9NF2J/Dz2v1gc6M4ARB7
+Y4qyqKI098atsR9AbNP178WDPsEdVI7w42xR5hD0Qt85R4RZoplnlKFwTOZW1RR
QqT6QvF3/Ax8FnMsSMdPSqLvlbqepp9aXcJ/jHw0Kfg3Hj3LN1ZQ7U/wij3gr+HL
L8eIBnvhmedHFSCzFRQB+zkLqsF4lrYvqk1OFFUT2Tks3jCNeWzOd6pqK2LJAlji
xJf8vzYebeenmjJ3Fy9x4QBH8dAvqkmZXM7/PoZcJ+m7lLSzcy2HdDwKhqzKBnGM
wOlqtw30KJ5uzvYUuwUZTesnjq8tzyZJBa5oCrpO7LANMDVrlhWzmpuIT6IEiMsd
4Pwew8buXa0pUQN1YOyhCGx4BWckBt5vAYneyW2d1owW46APAoz6cO2vTECfV7bP
uBaMIQeeLwul2Hnd6QvvDSY7+09wuW1C9PweenMmhnmE0vds7ppnU1pGrodGO7Ug
h6IkPur1j6q1xPMJtlcDh2LoXvF21p1kwzmOhnzEew+8AgFCqMdwMtKU6TxnGfyP
Kz7KI3SIrXwSwqy1w60AQGkL8Iw234yLB4apWZ7bbmceLVxo0gUFUWk1YIM4Cn47
w3xtJYjLK1Gqnr3obWbmaLKF/qeAzO/T/lfExDA/L7pRB6Td5WgqC0QYihdaO3wS
eE0wLh3fTCQ0iIlntEaBO5AmudI+iCbsBM+6PkfioRehKvBJnR9QyonVjZPgbB/3
/4uzDjXS3zkQYQ/g5RYTVGFP19D+1b7r11DwyPtQfsE9qoUuD/FslrNPz/LGjXA8
bixUSJQjOJEE+KyA4OQ21/Q6BnUkNntaRfcTp4ZULCMFVniKT322UbeUmDCptY0J
iKiHn7tqUIpae5uEXpoGO947EyH4nVkCL+XjEU9BAEFE/7UBOMKhgJyzq9hNTyY6
m2cMcHjI6E/oi1juC7GSkDsdSO2bmLzNCN3nGJLuamibc7Qwn2ynsf08CZO5i+xI
8l9G/mUDM2Gs+EIWi/o227bPvwe/Wxsy14eZEC6+kBMZrkwgeqATH4sJ96KV6Pv2
eqGQF5twuNO6QTX7hp6wSiZKzQYTTkoJJtmg4e2HyjyKgJqnapmSlSkeUdSwS24V
TR6j7kBu7/LrYS7Rgv/n2FNCI83D9MZwZ+ZdXgxK5Wp+CBgDyhOVz6pXbIZn0g8v
ZbKL8CSLqYoqbXfT2Sc9SDPb/+w56sURQKq4JvBu8y3rA2bdV5lRMZYejEBzh4z5
70K0aa7X20g6l/6bbel1CSGsRyFtk7ozUy12R6S8B8wh50oLYplfGwqtDavEWbaz
V8GRoJ1qi0LL+kQ3k7fqyvmwigBIMVPYE6i/ZJKuGXCIQvles6l5XCDzYjCbbciu
rucYXnmShTwoBBSkTKCDhrnC8U61KNr5+dHd/ufxdE1+owl7bfGSiXL89fT1+WP/
/9EMA26dIEovSxceoXn+vzb9QA5PKszkB/eW93UETK59XIBa1HvY3dl9pWynUMZ1
migjHLS5uxQuHHp4Un6IkPjVt2WEQYA2ErSKDqa0OSR/z1mkpbF5eEYXtr2aZXIv
v5Bm3FiP3ckOP32N9pIAcyZI6kr8jPGzgL7TjBRER04PkdNya98lgWs40IJJRFkg
M1QRHrj8oIoKrnyQBgrNmqBskGJe9Yxg76UeDwSFwTplq/ZJkyc88o06oX0o8tuQ
hlxzTUfAupvzcMxmaY2OyCA/pDz0fNzHB607aDa/g79XOGnFRC1DS8aQC7Qj0tJ+
e3PN9UopuhPXTy5LhbqCY03IS0KDGUNgkh7TV7ls/fuTZkYjDRcTPMMB4qLrx+je
Fd0eDGwwCRwiv7X0G2WBifetx8JGl7l06u9eYW0gFGTEtoV+2BzUfipeaHnH6q7B
JBVhNR0RTMbIUO1/vaB9Vb52N3MIDy1NyUYfMETpjGVolkWl+xdjI7/N0QKYS2aF
P+WukdxTQFL0FhmEwnD529Dj1cI3WAfbtlXsGWCV9fwpfTKWPtXZj8VqPP3pls92
zvgXRGHccrbbVCeap+FLtzF6MAHLvzDJPRHaKTmwfKS5uJrPcwTL1LxduOHLWcTY
Neu0IGwn8jOQ4lXzGVcxvklRxrV8isjeqziNmU8rjrlWDnycVaQvtK4W7WFQO9b3
vTU52q8pEyHfBrnDe5Vw72SAtg5QBa59EFDt7+He+OlmOyvf0rYpHyqpVPJgfljd
nk58111s4c8hfb1PBI6Fr5b8EzazqQYIYdKnJmHf3/MG0YR5oR68sNcH7rhZ0Uqp
liUttAEpUT2yERNLbRs359TlyonqFzylsuK7Lf77qy0zyC7QSpDD0eWI1EwmGs2d
XSEAiDlNz4jYzifQyYUGbW7IBPBXtj22LkPh29tx++KA2/+dMJSMvVlAqVv5eKTT
i2nUfDbf+j11YRFTFwHn+PcrKjDR6SIDfh3zCP6DCazg+hshi/Axoo7NZNL4xUUg
R0BVJnwBJ6jJBOq79CTt3hw1r5TVJgySVPdiK+ZOI/3dXhB4slEuUpAHvU00bRZE
UC/9KbmnSv4nIyeaUGHP509TkGJNvYPUo9njf0NugRe1W5lqYUPQroqHyP8iXdBY
K1CB9CLTsTNGm6RVUWbXt+hVkTlUWAUM1YZFu+mAZjhXpPLsA6oDsisRrPGyyHDX
b8QPSDDQOi3aLD5NpAXmCHxLyY1qfVBdPUIcGzNZub2Xu8mTRYWz6fzhXS0kcqos
C6ZFqqKTBqYrEgzsnQL0NoSx4/y+pJ0XqJogmltPu5d/OmBP0TYsuRJIDXqZwrEa
8H73CWkVmG4Fdr3zkdAWvPenaET7HXpo7/LTMl9QooZBp4LNTZjLWmof8Ez6MV8T
GzBt/c96i9aHvDmItjeLcXDqLIISYjR/2eoaZOSnmylOkjJdvWH0EzJq78YFaqrz
rlYRhdNTjjwlwTMa2qKAV7FSyc/VQ6DDWAPgsmkYnM115fgRWCLjCzkoysXpaoFE
qXd1LUUgaWwCNlhxBrboSIfSO+fYgFKScMsI+xx9MWbQ6IyrMdZsl2XtjDQdEg3T
/nid0RxWWy/8YZhl4+kGLbqyke8xC1p2+YKto5JlvE1zATRsbXprG09gnxmrWcUI
dKrPZl+NA0veHq7l472+Fej7Gw5zvYmoDMk2uyXuXy3pMomSz/9akL3kj1CtlIEw
zb7AmiN5+F/cc4+2aEjo8CyUvnacFuKNGX3uriQuz/7gP+xYeN/VDSlkfFEZJuQq
GMFCCdKHj3V17c2gI2I/LotVG80HTeakNSOCRe1gwYjrTNScTVFbimevMYMrsGMS
rJ4na36HM9D3+7fsYG8/QA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
l1Nm6/XONpooZJ6coT8GtlE49tODSHm6Zra/6YlUICx3KLjY7pR5hwaVj5UGTko/
QA4lrH39qVbbUHZramQC2xh5PjR30bp7wurJhvq688B+zkiMGlApOQtvSLTLkPnn
KxPu+GICL1t/hyBs2nkQHA/qABRg/N38J+yuItImrc121vZCQ8DBcuZpQkEJTU+Q
dcBQCSkzpteDmqhQ/Yq2MO1+XY2DMzcjuruKqta/EGLMObem9yNpOAmEXPS291Lr
kosYL5qKV3AQI0ZE4MFoOjCxWhlv75GQ3zfbVUh5VWW5cbIP1KEc2PmwZFCw0VXr
XG+lz/NmqfG91roY+gwD0g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8720 )
`pragma protect data_block
HMilHNN8Bdy1cTFPCF5aMoqXuv+WO+XUBH+qv7r4hDLymFDIJ7At8fXgPkuyfDV3
5pCbDUn+t47R7wfv2S3vH7f7qXkuwss9zIYuDM4QEMw6VPlOxNuhw87VUd+lNPPn
rvazeq9wH/YWKR9izeKPQkhIDc5xI0zT4agCVkUAocZRq4plVyptOtWzL4aJPxzf
VEek4wMzZWDEu7eJabYGHVnO3DfQfzFTa0TamPHOmfnYIz0VCoELPkB4qvwpGO+x
Lf1icEpDPyWarcY+Wex58t/w9oZAYxfeElFdM9ACDf65T4q008Dt9J1g7Tzj3fiS
8qgKSVhlvm/m2sVJrScSZLV7eO8BcClBf3LVOWocTY6KtbXUnp1fV5rZM/F7mR6H
Y0ymhZDYPB7HaFmTq0dAxpgXniu2lKj8X8Ty73n/ir/enKaXnhOhct8y/HUoaqi2
sIGajijXu8h8KhYzZ4biFMPRKzNhlOGEyHbYu7ug2S4QI3APOiyNRX3Lv1sn2OPl
6BhAbPlDMHt3tUkj1kVDHVwJpIWChrVkDOpdIYtQd/f6n8OXxfWAq4H0h68glDlm
WfNuEpwqmb7yOIjld+kE4xiadmU5duacodUS2Fm7hA8vD98Z9GXXKwrL6eOy5pTC
5LLjyAv454fDMm8SGZMooXIHe+8osnrJ5f1khUE+YAVLX0fDBFfVHP4+gXWDmy2i
TvRRIVn589d/6GO5XWBFqK9058Q0yKAQxz5MORPfs52VtT9QD5aUiEuReZJKNI9d
s+L0Uq0+r7xzZ8BVZ3P3aPCL9rgNjKqWl5/789t+WdNcDJAv+6az5vBBb8TfjZ5t
U/h6UJUkb0gMG6Yd7nsk6EMq1kWxZs6F0oyhk3THyZ0eNsujE0oTLVExIUqjFZnT
HPzsv5wcZWiTrWRUehp6dcjI8ro2z2aMH8kJ+u3tv6i/sV4B3fjhTT1vboBqfa75
RM0iL7F71KY58yr66va20uIPu0puTU0mUAnXZFXaJhpeTppDUc/xDTgdeAnyAnKy
FxN6wYoxAz9tHpx0e+OyLKzvY+YktmOW6T+yAGOtY8Y4oPkt+K6M9IqwnmQ51q9L
8BgaO/vacdVVGkazmKHEh6Cblwrq3/ZIafSIMO9a0aWZLXH/So2EuCzS7/f/TKy5
E2RgHPzG5SBMVbdixzQgkD2nlqSBPqvrOQe0kzbcQoE/CMbHE/7OUz+yM7Z/xhYd
bugG2Jac+AiJSygDxnlN6w8dBntuTdaKQjD2ii3QECgrAmMTKeiKQLZ/SQNVW4xl
nAYgGjrVvJH7wEiwKnIAuL+NZ0HAHSslYXr7eRAQme3dLE8gT+rjN8qPoMAMOxDG
FEt7IQFHSRouNw4RG6+0gUElEEXkx+6I0XQYLgdTrMW7AiPL+wqK5inLwwyfwa/h
uaFYAwfyQdQpSsLqo0Bw7REhYKMKpjGuHU+nAo/CK1Ik4+eXMF8V/9CVxRQrWJps
Iw49cMAF5a8VP1B+BOKKCalBZ8hJCZvGjIFdWmDiW0/G0Z4tF/4YXBk59kpR+ioP
uf5YyR9PDfrKX10E7E6e78u4Aw3PusROz8+8o9oUdBp4oJ9NAzxFFEwcjnU6+eBu
erXHM3igVzMCFFu81rrHpjYZUU1oZBkVAUVXainMfqwzk/427RZJhlWf1ddlcTXf
4r742lEtUKGC3aWO3eZJv+bSzqMrxPEEZmTX47RejrSMy53kCPHKcUaBvhHgbAfr
UiigqB65wXWZ1D/bdqmz5zAunXpP/9wZaVRr3X7KW84SBgQKuHQvKcD+QsoF+tOI
CfFsBnqwIrakSzj8KBnIFudoAPKD3GN8OHA0iDvCjiziISJPvCqsMa64f32+rCus
RLCgdao0Y2VUj701WLo0o5HUO9iWGStJSlL9w3jFbzIlLcjUf364AB+y23E0YnLv
PASXFFddDqaXzbsec8NOn+dghkqcRA/j2K5iLnEDGCirOTkq+dqQOruEHKaK4Ksk
QjUXBVqXejh1C6kP0Q7tHC2Td32lJtrJfg5iRgg+iQKQ28UVXWCBKvY5Q1Y0kx9e
SGbIq0C26qA8O8ruTinF9VYOhiX0q1PKtMattFz3nApDd10LQHpu+KN9zlrSr04U
DcQu5xleNahdNUHMTn3DE8ZyIo4jQLRq+FAogkrsVa3X5j9WZR2Ro2L4YGkZiAtB
TsXnZe+gaXpSUGY/tks+q/VpHLLBzw7h9ieu7h2vdZrFok6GtYP+6XtNvzpEvfIh
xVWvsMpvInkU3o18+YrI2pQwdvbwdyGDi0/8L1LBOk2uxJ/dW/H8ri3G+jgnlJkL
yofIVkErYm2Y4YeXKw63l2jGW6fOo3fzhc4Du6RkEpyDtacNDu8MTpwdVI7A5xX7
e4REYiSiAcuTaQslqiVS3kMn0U7QaTbXx11NnWPoPQIL3hZ95f9I/qvv+cTVRxZQ
JaIz4wz2o8Rh7TP8dPhgCoQwWIsM8Ehzp6+ifd5PjnUfBsIIEy5raxLnDP9k5Lrw
ycsCxriPoewOKdf/ic51jddT2NeGwskRXwzT0XEqi20pdzCpRdyuDRnn9NahYOKu
f04o6kzUml4SvU6lRLrb34HfPXwbSARplkzfc745H2GBk9/aG6Wo/1qgkSDAwbm6
rl2oRZhv12IqL5fRpvMLlhnIhg3QeU8DDLaIVqbkby/i3BraTxHQAWjg68jHSI4Q
yIpPimayg1iPqwLM4zQSSuieOhCNYc1yAicdBuW8gh5Q2VqdkGICvKxoPnA/PaQ5
4CtqciiZbFgSesRYn/dB0OatJgNBwQDnv8w0w98I6QlUhyF9HHdygFewbBU3ToVu
UA9Iq9ijTjahoGEHZBPTw25Z4pgZUWOzvWJbwAsd9jfB/74V+xG2pOa+RybCPumq
gSle0CbFPVTdNBAnqVDsnkkqDgf0ned3mT16wEryJTx1uct1J2bNdJvvyq9iH99f
CGLwzIZL1s3pibhQB2hSPO9J1fZvAAE+9w5uBGUsfzhdf1r/GtXvtU+KOvP+6X9h
W4mFKRUx3gCFSDIFwBPHs8WLpI3ICs6cc4At8Utd5Y8ITP9UhSQa9hMek6yZs7pq
M6BWzPVAYuinyuR4RtJyerL4MCXYyH/3lZQifUvDZEKycGJbDmJTmYFZ0oOZKugc
4CU6rBRA5ydXTtUWGBJbgRvvC0Jnk0hIA30aaRA3nu0Dz1xw5LsAgLjVdnws0xD7
EKbOYCjWIychlcnjekYXQvkM9tJLHnsmEkQt3ZO8Fu3gdoGim266/dV+rmlKB6rf
diDZLYeGcgup0bp89oM2nkMF/jNo2O9gq6xXeChJ5f7JDNQCXAQTCKOHu+5skhnB
VGVlGEAmVx5tIWiO2CtK6WPIiXQ3mMKQoefsmmMLpV0MyCfEJ+rseTt71K91y/tE
LDGzeOGr9C5ZV14H+AG4PQpYWw+lrwyxE8Vw3wenUTPaqQSrihtRvzBR51R1+Fbq
TrmRR4n2htetW4VS/0LKjEvtzb8s1aRcD7Uh5VTE/oVmESLrXAh0crUVUgd7ZP9L
wAealRs4hHoPq/Qm03lhbWuxXwUR5PwP3iDBc5mfN+Fx72p7hEgIThQXfuFojsGg
EO7Xr0hflCyJaGL9mEwf3ETDsAgNfB17xkThbe1HYvzqITlkDMDzsGiuJvQ3eQ58
LDRIiznGIBJRkugRqiVeTfIps3gyHPvPSo0yk47+jPumY9uMqXTDq1lPelAKp/n8
4fzs6L1pnWjVc7yUV011pkDSVa0mzM4AUvY6VtwJNjnOj9rKXM0UPrjzzDcp25oT
oYqXUzYzDYvFLFlPj+FS2pK9Icoev1AiXJESNQAH0SQkIg/zlPKHEavSdODsyBkA
qMHvyF4PQ5nJ0n+IeubyNZqSdTeivOm/wRogDK4kLP5Yr2GCjHZ1ZqSvf6l2K9+a
5iRJpra/ivlTZ4kx/NtYI5WywEPQWf5mmN+TbiyaIR1iv+UKYlSLJecE/hSFOAeb
Uw793rvDflmp97u8/Q02CVOpisGJbzeNsc2mD4F2M1ySZgFc47EG0i4aDXSXwGn3
kO4PBS37V3x27JPpX5pmhOnPbTJHp6WKtTPJTEBn1zng6Z9x+/r7Y2rwtodsuc3J
d0O0qLqi+zfUI8jTvIqB76q4OH8Gz0aW5QwLJ5tUzolMjLyY9R5v6H5JuiFVyq6X
D5k5qp3hw6lD5a639tLZsqyN0JfKHvmk4nEtX8OLvDvDfB8sOo68nHh3QtMfefsl
GywIQdcAtTw0jMj27AfxyE2+Hu3Ksa3BSRW8JAkMkNh/QRyXYlC/1nPntom8tpb/
S36kBTFztvvtB+nxynNgrsTGgJLQ91CuFkPrZ4XHmG2uDZofzRptQGPKPHdAjcRE
nymDLgSF/xw1DnQNcXy9Gx54vnHj0DjbGLbf3JEHCJEQwbDnW0U2fWFYoxOCosAE
uu0lo6MPM3CtpMvxS+9+8WA2g9TgQ3Nc3oyKE3boGKUDk6eK33oR8JkWgQvrrlZA
Gu1q/AqYTeAWBvC20jFfEW48s2dAbVqQGXNBDxRJ0q3INTp0kYKpXmB0jqg1C2Ym
WGEszAOsyIpqWPKfl1D3uc175xHo18q4a75y+Jvmb6UKOh/TOHaFn3yiMkPgx1Wa
7z+z+1y4osTpF6CKe9ddiFOQCOoz81mRIYlNDrhyZbDODdbFXS2TNydh5HQojBHd
K2hqIlGJ05k9ZXxFwAw74SKWwANAbnOvgKqAIND3gXiACc9zyznJVDQ4THLI8Yam
aDIP7Dgf2aAjW2mm40GrHKpAjEzz6IQxSgZr1wTfpAQbbZQEwb8+2T/Uk5f285YK
3sEMzP0AN9J4guLLbRaJ6afoKuX87Hl8APvdrcG5YMAJGTnAPO/2NCRObGUGPeHk
hJm+ocKce+58skR9epIR7FuJlgHeaTtG2s1E3tfmhTUF7TvRNdiWXXPXk+fo2/tk
dHO+IJ9Or/iwZ7Ja+7MZ3MBi0yBkuLSiXzrgEqldjcGKo7zHGMrreAcRLsF5Nx6I
K86e2AaLveoViANIhvkPjXsC/XD/WScpSyxdmHeqoqeQcrxFGw3tXvlOPnhObwfk
B60gLz9CDWB9JElTZxHOyQeTiJSzRdOhj4d7xYVd6IlTfEeb2/FbGgsrIabMnVFE
mOdFvbj0xFrYlxx7NxMwO0eT5j0yEZFfvPOrfcnMabs6t5xaFdH1v9KYST1Y6McX
89lHylzjfD4MNAeimYBwRk7Bw4pvceVosgsXLuuIdcjBXI1521ynacQ/kTQ2JDbn
LMoIwSjmq3Z0IJrBX2CMPv/T5e6WUsURGSEfi02+LqrmAHnB4zGjX4v/5SlOeoHM
xXO56qIfqtqFAAPS5JrBQGDpMDbiAS69jMMtCHyUFQ3b8ZQh8JYH/X9BHcGUmq4j
xuvjUNiBkA7gMg6HaMXmmSIQRKGAAP/v/8QZa2GCvuY0gUTX+dA6kUoC8zLkHic6
lTq1x1PEU0zBGdYyM0ktaMpGbuv8gAB+Koi4w8X92bD0AsRuQZzAoM9AQQvj07sC
eRT29kwF4GYs832QqZV8S/duRB5mOXUvwBhnJZy3qxMs6Y6917affn3uMD2qFNSn
kfSRIzPUxiGeUB5g5MMYfA/39DdbRAWPrky4WG3uPl7s+7r1XvtSS+LSo/LGvbjh
fy8LdDHRirVptSqTyL5ndWRvDBQkc5+CM9Tq+VAcOWJPJZvqPqTaoXlzAnJNambn
CtnPUGHKvksUlpukMVUNuwJ02FTu0Q2ZIbLxxq1nuxg0AHJUTGnlFTrVX8eVB9h3
X/uRuxKvpJ2XBcDlNCXNRfZDZ1weykRANMmqvcX7CYEgt9fFvpza1ljWcU7epAKl
d2N/tvNg7RNFLiGlkucyaZvCqFy5BWUDICDE03SKL0W0BHTm04mXIe2UaU4u2511
7VhnDzly5MX5TkPBBFIJxcnNkHwiaA8y19jtDcgD8aG1UoI4d9W+Rpi+ykatJWHY
n9mFitVlsLRt+koYPlbdkwsOffjOlGiqmFneKTmRaDOe1fSIetqO8e1MsNthkZYq
8uW+NZ23A/YpocJXOp73UmJ0m3ARCNNz5BxG1HW7FxuwcxVietkYcnTDnzFVL3e1
sqACTK6FiTenNGjrjlENoKgtyyK1og8e+IH3bVh+W3SGj7R/XjuUvtVdGm0ZJNl2
b54SFMTKYwMRM0U3dDt6sIICYznnAguqj0Kbv0Um+MGmey9KzxkK1JQmCLuScK+H
nZXPz8wtOl5dCoYU+S4oWJv2jHQGNURqnmq1NNGeikRUb5o4kPu5IX7TSPt+tPxa
Xjl0F8tiXLcuZDCNhdrZC1bnJJpTYE4wqctqtboTLEuIK0VKLuYPHeayeySZE21W
vOWloFXfKvue5+fVvfHZa5Vblj/hXOw3Kh4kOMNnv9RPLwPZlvzUB1PqpW9sdzeQ
ENhXMQLGXP5V8u2gLBC8kJsh6kR7wt5vrku8mqr8epETUH548+W3gkjZsD/SnyZz
mPd1lQbif+Q4pAydhByPCD5W1gHN3FG/FJKk02zBmB+17FzMCg8Tey/xH6j83wE2
TKOL88Zb+pYTRhntVJ8Lhvtjx6tPhLaSOMm+R0xPW3ttC9Nyez9c157jZCw0dGso
HX2YtXOjeUk0+zDf8TYdWxIg4+twqafY6i4rfx+ls1fD+W27yBeMfjYARtfk1Her
P1Tn2IOcbSNdg84aZfOvWDefzTItemL1twKrG/e/oEYXv0NNd8FDoZGsmOD/gHFo
xWZVqpOXR7BCTzrPEIdqek+klq6UxF1wHdpXs6S4ag0iT5jX9vBrNWvPG3jhk6XC
6co9jdcSwzSio6LEgI/VWHcbA+i9YdMCSWg//YKVXh23UNUnSc2AzKETy3hSVyON
5Auojtsuf/orUeY5mYUlsc6PiIksMpmjczoI1CxiIm5WArdBllY68EOF1OjzhV7s
pLu+H4advqaLBpShEZpwfcY0wCKptuXPZGwj8dLneYDXDKSZ/qJm9Y4g1oU1OMB3
zwqPdF3hJir8cg+n/me7ufjLT4WPxh81Xz8mnhQ+OzuIzfFa0z4zMPnpQAz6s66V
vqDP9Eme7TcxffpaWrt4Mt1wixzsCP9GhtiaBEQ3oxHUST5+i3xkYn2kzsN4EX0I
Ydzx9fXSPM/8sfkgSfmLkJxd1dfDbI+vLNLkrLRKJJerkkqFqcO1hHKZHvoSyK5S
pMT/p5fqZJCppNbofYId8klTwoJ5uTOrsk7XdoRXPA1jyBq3IUY1X6in9ns0e1+X
8+ByoCi3BMceIGsW0wxLdq3nS1GmAXY3lsuVLQaDCXGBhHHJTxhIF+SKKEvLVhP0
0+ZAQj8IkOQIdpOl5BRZI12ScG7h1mluTAOZVJAtbqCzfvl9zOBJD9JnEP5hJBl5
BPHK5pIt4w1JOXjgNemFqahYgQ9X1EnUzczBW4ELblrFWaF1XBFcgnzUPyDSZrSC
Xgw2YsgeCZkOHF1EZecW86ogVc+la9OY8bXNPsvpIKnYfRkkTQbRxzxg7nEGOqr/
CfKcWb2h/LWFNzL5EZn2i6/nLZUq8StjGsEEuebfd4+zkqdYSIptZER3pxLmer6w
+djK2dZHcYEbAQZRVVf2oUp2vhmVZ+i70WQIP1/Jht6nRC2Tom7uLbJ3OWQuK6CQ
1sLiYTGQwIsnb5rzehKamLh5XY2RGGsCBDARGc6LlZV0FwWszeYLzJCimBTIJoDf
bvWRQUsU4Ajk5SYpQ9v4u6/Y0T7MpiaxTpBez0OVHENxEDxA7+cFRAMXRDoiAvQz
UiqfjDHuQShLY3OBeM1X54DeKYse7Q+oGU6GMIMj03zVYDNwW7F81cyUPG3Cf+v0
pO5K725IPAQoSl991l45TCsW3HrL0fE+mU1Hq6s5pmaqgbw42uakRGvhbaR50pAE
Rh7HG67LroshvkQ6oZgG9g9eYxdoK/QqDvbfNU867fx6g2fHdFwPf70vAbAVdddy
PQ5yWNwUSHqqIJzPxph4QvjPRH9NGBnH/SCF36z8TKIghLCnPUl+6oKVzIBMhp2M
oYEkqBnA0P4hJ8dvx+fGYYET+Nu3M3RNbD6hamRCKhNLan99FiUGEUTqghaaER2Z
FWtHSVsN5ixMzWXGC4BSK8SMMF7zQkDG4iFQmrcyyXeE2l4LUMSsVM+kBWVaZAlR
t9/0eY6X7B1GHhOnTeLJjUwNo9DklLdFKRNgDlCnkHWw1qMaT52HYTHX8VVoRZPP
3UWZyF7TiqNfVrv8xRw+UGkWK3Q8s6BL7cHqXT5h7G8FCif/ZP10q6cTe59TxgTW
ugs+wXSED12XmeBDPCaZ/mIPFx5XW4QkPpnApkrnocJYpjAjpZHmb6UGVTHT5aqw
hf9C5TEmVLJpGsP6VdNxhGDl62Ep1bZdYe9ONVqVUUjKBdiHIwEzY74KDHj78Nz1
YXWV6W8KgIniaKwrxHU7C3LeB3mp/iYuZtFDamdTlLdiFPAJc0Eb5ArxII41dNE/
oTfILvvPeJEfzRPXokHjb5pTN9D7kbO8beLmNDTZaQAHZDI34+diTinqNxdy+6P4
RTBFMZQwhUsAdVYtbMXYInzduiVbmD9AV9HOKGFql0Y5/yBgS6E6Qu+qUrhof/Lt
jVTgDhA1RG76oIlvPCtZdj0i/eE/itAF5V2l9FLOOpKWOXx/uLfdnJwMYk9qgVBO
N7bWB6uokwAz5nvaNvxlenzWqndFf24msgkBoI7aMwFRkIj6gh1ZQhAiNqZ+6FwW
6lIwHkXyQMyVA1vWninqE1c/ZhH1t9tVisKXuYYI/H+owIM34PdVSVXrCSlbv50i
4+dFZPgryLrzB3PYX69HAWrUfgFaaDyHCnoFpdcNv01piJYSZ4kDUEr8a2H3Qbk+
/Qpt4OH2JpBPIsSxI9DVJSZbZAVm5coRgWSaOdykP2oG1TeVRzucywalbgqr+G9r
MLf6esXcHmLMgWMToX5I/3I2YPH3X6VXRjEU4mxQs3rxOTnPuj6RVyIrJSs+k413
Nv4DMdDFAH47ORY32IyLjCvlFPLsrdJmwzvyC40K8H3aOYqz1rcI1wViYF447Uzf
bhTeRMHnnQDLfgyWDtWjaFspKF3yVTMqMAZATArxqBm+H2EkBGBDrSR1Uj9lo1xB
oPAksgEim2PIAq78N9I5pkFY72JRWnhDnPUY7yxQs1Jxt3UzeZ8O1CkkE1PHJnQY
a5G8WgwjNWXBjJrrihLeu0R+V9PUeLy9QY1dCnPmbaGrRXn5JuE1ujD27AfgIzh8
2ttDz7KzVySR5qAB4cRKHE2CtYGdM91A10dFcdoDOtFcLZ0EdJbwu44VF5qMPbgQ
7d+4DbF7bsCzydSJ6DGkQnMNIe3/ZKigNRgsPVVfwdpATEo0ed73cViCxjbDBZs7
/xxIqs0dQBExu8laUrNH3Ut0l4v5HCJIkpDcZCJZtbrl3CYAAxepZPo+8ALRvKIg
7mnwVDlomYw0DyFtFao0F4c8R1aDhWN55mf1sMQ4Unn7RhMKQJ8vQkD9eielqhhP
72Bsq9ps7Pb+d4kijaxtj51IC4rQNIuw2JQPRa/PyfNv5o/be7Fxw5sDklAV0A8s
F1sd7sU66dxb3BFxcoRIHzfkCmho3qUNnxbuKMtWrF8GYw0Pswh//vrItLsOKgvh
a0CF/8PX+tM6Zswr49LenaKL5Zfh2Y0V3UA8kE+PC31J9kYYm2QylNVtvpQk91ub
NN0KrVlUbq0z1/brI7ASV3XrBF+/jXk85jFO9XV3YuRt18arZbiHRBuOojiKyX2O
9fN8qUjQoWtVSZmf200VO1zpOyf3iF8JpblbM1e/M0dGHk4MVQipnId40y7oJUm1
rPxQKbj5/5+F0tQCp/Bo7DTRXGP3T6WTa7umfGY1nZbrlhjzAjHdyvNCWvi02I8C
dfWNNlrAJtSvJz4sZazTHcubUai9By5xHoo6NbGFsJOXaAAoRfTosnhaN/5A0jmS
T9hruqXBiG9jKTneYSGu4L+lYvRvB3J+gY5gIAIpAv8Ks+TQ0+c4kfGhCUPkHSaW
uR9cCUgE3euJQN9YaD4a9Ln17xXTAZ3+EBoAaM3FJyZ4dkydjBgclQyV/fX2bscN
hdPCF+RAquH0zqtJVeiWGPHFmi1qRN/RjVW/F+dK3stkQfK3+Tph7P5AENsLExeL
0CrhOcGm9z2VhAghmGuh1jsPVLFLvh0iTINNy44VNlUgw3YhpVA5RcjLP5/xzyyi
m+LAh7UvCMwaoQlEg2czH/ODRD63OYfbk/Rdk7x4rGWBBQbtb0MW61epDaFbj81J
fJ4P5ebRbIriwqQVD9z/ouL9sb3FCLQ1Vmp06lIs02jlU3zki17892icawnIT7k7
oy1ipUXAOkZ4RJm8p2VZEyur9nmcQ8cPBMTqiqq4cup1z/l9BFHm7IOatjk+JT7Q
TumuFQxiD+a+UnKX5LRxXpdDhZD8OimMSM18kfmBUoN41b9HrJK9YYHMcf74jcoA
Ub5saqlgxzE42NoqFeTvL6gkOWGNFIVVksOqEC9XFDYlqQ3WheYnLHzlLj9Lu3pO
dMtuPbRvF8dyzVXLEqeC8UGPNjJvzJLQzN4vWqbjI27ivHeSYSI3tU6aE0gCPt6L
1D1e9r0wL8s4wjhvB36J0ASlJiuR2g1X7gDYGvog4NSg1/axA3iqdTY7gV8KGSHP
ftb1SNLn4rKhKHOsbKIvUKOO4kxkBe934up7TZntH3dPCc5BQ+NEm8ewAFeqzHHU
G8q/QEZz2gg07/7PonTea86c2wYAJuHbPn/l/k0kuGahKpmMFoE6GO0SNUOa6/+1
nyevQADOVKAffWM7Xbzc4aS0GErGIwP6eZ9djJx5Xc7I7LQtp5XL+r1eypDhPPVW
BllL1qntQH/ovo43iZhvPtFL7htvbRhbeh3nVT0XzMv9fpEbHvc8SACye9lZS1H5
Ing+3wz5xHwwtvbY3MRxQZeRzs4KyOe/3GrVIgkHtYRf3uPOsXQOD0U9xaUYuQW8
OEdGE4eAOE9Ka7eznlMiEaANxhEtfii9CxsqvktTAIk+Z86q4Dut5sMqKmLDMsDp
J49ntzSSp41HGfW6NaCDSb5Z8G55Xi4lOX6/E316A7UE/SYPE00k/hSdWdefOnjV
V6BXX6ObsH+kGHV/PPcgxsYUfZzW57UHnnvuMVfJS7Vs67cuAlPUGEGtQ1s2YtOh
Vt0irs8n6FTdlPU6MV6EnEHrOVKWYsGxzKroCICRKB8MdhjCxgN/enhIyFVQiuyn
BHLuv86hPXWcOojkbGYwB7nVnrbjDmZB0c8UenvsRBWnkvGgutYXgE9XP915Yz8+
uCSuChK24ExnKtfXUcHqZT2xV2/GzSNFD5XerulVxGOZR0TIK5Dr6xjKd34z7/6U
KcMbtNTh0OX5zuzou8TD1LglojtxTptdLKLnk3v7SSwMxjDqmJRbUafNVC2AIdQ/
FJ4Sc/PEj7n5GBpqoUIKNZD8j/TbkO5A3Yb7PcaH1JNUfHzTj5Tz6le9OfChSV3M
i1Hc+5NRnGr2FLW2sOlDw0GnQbrOdes+9SxY1xpnBBT+WYtKdtg37aKtU3IBxMZ4
zCFtcyKY4q39bd0Xin9pq/VCgAd3LXMgSfp+aa/ctorximoZq/5UtHEBHJQpZRhi
op7sTnWGppiFiYhDSC+COwuWY5YANxZmVAf725cOPXE=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
YtJzAfwvQxEAqheFvvhosOhH+Gx3evXf7jowxPS9FeoczMrOfRPII3VdwQPjd8Sr
y/g81gxPAlSI1t4SXS+zQyBjt7xwBPdQqqh+Jh/xduwsOCqmGdQu8nacX1BVaulm
bxuQxkraQtw7K1w9VbwCWvPePmFWIZ7bW4MvvTH3uSntL7HRpZ9jJ7uxDc5sh4lj
opU1nBBzf8WkWRjkQ1QizxRzC20JCXq+HsoklacaivhNg/Cir6N7vGLQQjsOuLdw
aJ8YJWmxZVMVzJvKhOQmmeDpYSqa+Jj8mafJD0Tjo7Hd/6BGv0XV30gPaPmQheJE
z1vqNHhUibuuCPLIA/OJlg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4336 )
`pragma protect data_block
8HqSAHhDL6FeavLeSExLCyCmkgSIiV1NSkdOx0uBny0bHd9mi65CtIvI+jZrQyAm
NKwCEmKzgjDG5LusVzHILVGOE08fCPdTnQG4tFpIENtdZ6QsUzuaKRAx0n/Ni76j
UC7ECRgf0IM3ZIKHcc1ohf94lkL27jUkNygfTBeQ3tK+fyt3s++QkhsQX3PFZa86
DmT4hG6tNhc1vvwXQN1VIQTwFAdfkg67cgkkEHvfz6o2bHKQ6n4my8mZVA11Ncl0
XICKbki5OmNpH3QCO2ch9KFRSfBlVpsNACGIfGBFK1GPip0RJHl0FFoR5RaRrxlu
MRhamj7uw26i/oPf9dD99AIYhSGRb1DCA294v1KpYluTftqMbFfvcCAVysnxaxjh
Rhdt0aFR7gc8idT3sM298VsUPr4u6GcDoqlZJFg9v5GS2yBX1N2mHyZsjjkBAeNI
QZlhavFyLRok09MHUxmTOyOlNpafMpCcx17B/bpHzpJF4T3AA0fodn7WBUAi7psg
lXV3Qqg9pbPL/GOTLQETekPbXAvaffiijTSIuOEExQCqDtU7M0dFFmvtSOon882m
FcRW5f9VgQ1NaTM27IoIlJDLvwq16M5Vatu37dUYWSizhsj1gnUbhsIFR2AAYKvP
Um4vsY8a1B9iYIiSJsLSnKTOLydP56oT34GssPXB6U4y2kAs//9elYJhUzJano6X
ipDuuo68XHBFufg4xZeDmXdSjvJYedZ2oFL5JRTaYjmUxAoh4IFexMjQSI5oe+sf
ruiRPBRPbwjMzjO7WWhXaQsz/evT4GAnVkNnYJ65oQxdONKXtGuW0xi0bvPH4qWL
v2P26mtcwPDRkvaRg5o9ar4hX9W4RRSzvawJrmWpGQxSlG5wUaMr5KEIesqYwdqv
v2Fn4tOuIz0GrRBQSNyjoLhx7mJ8nugc45sklcP3vwu3stuvSupKpIEy8Pc2s6j5
kEjRony2ehs+aKP2IO+Vzyu8QlfVlLvCNZA0wvByHNI8NdFGyk6N2uuyllW9Xn6S
Z2ZpELB3msWit/RS4pUiWc2mssb7TrGY0BJhIWpr2X4nt4245RSZUrJMZ7ylx2PV
U/Nmlv8F7VrJfu1+87rAa7/VBFvThFOASgZ07PnBvYDpbs/Jd0X35rU4TZe3VIck
D3qBBIeRFyzQ7G9XmexLEpwPG6AKDSNXTf22pXGaBehvV9Z1CNjrtkUIoIXIowvw
40w/ivndTHrTI8yg9G+4uyOoYM559CdqVOxEUzbtWrCRbG0LIW2Eii/+CVLyvfV0
FapW44Z/CAHvXaHc4EzPchZbHMS62rD922UdA4aDE94zy3iqZgSn54RSRxqYrANr
wh2XATqPwCj7qdeFPGeFt6uFaE+1CtFUeZmGI5UgbsNdq5BHpTkk5EvKzHHxUIFV
LQOvoWhkJv7V/CYVbhWDdnMiKZa5iH8yAsdpyjQW3Z7T+JcuSALP91hzEWYQGW4P
d3Feg08ZAfN3FGC8irfZjMqUFjUBeCmfdFRtD2CXOAg1wM1C4COuJ6g4oZdzXrLG
0+12TGA+ZUvCdnFmNRNiF4gGRwKd8U/c1k0lzeEHnvfvIGq58PM5EjjMW+FJD9a4
wrAswovXJLFZOq6BKsTw+bQ7gPAsHgGfb0oEZoxNGiMtebV3lTW9uPRn5a1sUAgJ
oGuDNvByg81h/mqTgTKTzkh811GbIkwI5dUCqhk/OgaIBmN64Z9rRAC3H3hmwWwl
XlYA5eJsxnVIuXAcYhaacbVJhFwXxEwFlaJuvtRrxFO6bFulhvJevVbfmihRnzgW
br752qMb34XmVQUJ7G3Rs5sY+Nd1ls3y7IKrtnYU2L7TIrZpLchg+a4mmJ06kymZ
qd2L5xnmAs/n6seZcrP/yM2ak2fswTmCbz+G0+1H3g5cl70WV8mPoq1PZqyFx/Zp
ETan/ebPus2MrHZQNr1g5QUQDSUspYN27nz/tu0BYq71zk+En6zt5FdjRduM1WkT
StOiEFbQwRWeqjsP5lEU1mE05MI+zWzhXP36E6IzdirxGzeHhQ3ras2vYjnInnaF
hERXOhK08fWHLCuFduTzs4t9uO6tIRs7QMuyaglb4sGHBy7VhTCVUhnBBEDpwkcH
1Q+0KSIS+Jq0Bt89ndtXqazt+vPn1BvC3ysMop+jeURPO1Ig/wQ/6XzFl5vl02w+
V75f9LYKh5oCl3OilbJlMKHEEm1BBWFDXqYC5uhSAuNFQ63q4oj+5hxMtHhoMb8a
03jWi8zbh4KMSw+G29ywa2E+HTsAwee78O6S7yYnnDHzYTu2yAuVJQ+5e7JxsAcm
4pAgLXOUx9Duhg5Ov5BtFCQCOkD4sw2NtoiDyQqUxfEU/q60189Gndb5Zm51XN1+
cbr2PFQqMGzReDGEAL8O3N6vnAmIdPmreBzSO76q/U0ASMvxwGQ1TaWizQs2vwsv
cQB0i031eJeMhNQ9i4ckibRqZSSUzQqXxMcucESKhaMmNMrD8kYtbTUQbHaQKxdI
6Rev/Z81wtDhy2j4gnFIqC1tOT1Btz7yB1uzKRDiS+KTKIR06qbQmzW9Ep/bvpZ4
wqvmz+JFgNzKqY3UwVdCHSdJJxH1ma3drHNplN4NW3u/T87J7DZgvSH6FAvtuYUV
/tKKP8vqhk7U79n1ufeQCtU2IaLDlJ2f119BIYlfTnv/xUSlABESLJTyyPR1vHBq
mG1vciSklnTIDIMCg1HRzwlAjL8BCaSiXvUvCeVWRk1UtYapzrtzOL9eFrocASgN
JDLZPZeTiOCinoszABnXIPUVScGXciJRCWhG5M4HqiLCnOblGH5OgthUf02JCLg6
wtkyWM6g6TZsNAvqB2fSC7lRWsI87c3XyIP9nGfQjkttA5cBU6hyjrZ7RhS9zVla
4ZIBUBO1IuJEOSy/pkwSn0N1povJuZc74ASNip3xMMsr7XIfZdS5kvwOXnLgpgiq
BoE5HasiP3HBswhW9xrGC2P7OpurX58QSmZRAu6kmhXhYe6HX47JFhebmv+4kdNe
g3F3X3J3Pha9KxFj+GRanCWvbh65acE/d2EQk/ba3WzPNjmWfli8A47U25zU7Xnp
ft5LQOq/t/moobE5qN0uBJPyFnA02z1v5ZpTvb4ipuEMGCvzLVol/2CHKhGsTpGm
1J88SAl/OwXchyHrCmDA6xTX+dOrRQkn6SEd1IzrXr7REP8negt2eLLpXj9dQwcu
sbVoron3FvehcFdvLYds5w7YXOWpJIyT1ZquVnmr38VGTCHUJHWnkOPh8XVDMZ0u
x0XJiAOWC0w5cwm61BUOtUEGVUjldlWTmaF1P17cIfSM+UWG8GXpP/kNUT/kbcLj
SdO2JgbJHZeUTDFkfZC+gPwr2tfaOeuigZtCgL0OHnANh1qwRgn9Tm94zOcbCT1x
Xy+fK6xqSGOMDKKwjjuk/Vr+vFV74eQwEUb/5ejVjo2zX6lE2eJo2TBbMdcD+jYu
WIenJVJ3AWAfE01qvPRnNP05U3nbj/Rq3mvEliY3KykbjP4Q+aAXThJWdL5edBHU
aafRXHcD55eMq8DLhzsQnweGkatXEtK9TpOv60ecrUhCOSTx1mVGck4cezGf+Dwi
vPRwvsdkFsUeyYARfdiJ2zrgDOCYqCPYrXrw/Iza1ELc9KX5p2SJpfPTNp1foOw4
4UNYnDDRzKT2Iz78HNRV1dPynOP2RPYBgLQEQXsCCg4irkPX2f1IoIBVVwvb6ZCS
FgfbrDa1tAs39IMVOXjdusp7oGp97QiOTk5lC3YU0QqQPQvkkF429COwvI1l6hOF
tj9ybKBDTG/05W7cuQLiNGuCiADqteRp7RyByM9MG7WzrBdK9SU9Jcu9VvAQBNft
yeeifcAMIkEU5XBkjp/5IMoaBjpgKcGvRnMk+K1HiHRQWpn3un7DUOn5lr7Ux6iT
VViScXzn7YTeY0xOiBmFL+KDIexlH8iAUaYqHB9jN1Ou/AXEYCP+bOLIEKY1V6zI
isB+ytOA7QU5IzkiNsvGBO/6pcfcbolfSYbkhPJ2YHgNfesYWmq8r+6vbyg7OMeP
TynAHvLIujrona0vxseDX6sM/3V5EQ3B6W+j0bfEOnkMJ/oGWh8Kj7OJqHZlLwXx
ykpHK3xOTQmdSle9+UojKKOztuJrv10YYZa1BcNC5d0IBpwY8kiQ8QC6cMy9KYLn
wETJvKj7eYLJuVLEqDphqiAYLMAiM0+gmz8BzrXSRzHwRG4MAPJvMg07gEA8l0XR
dC+awAz1ABykjdfG46ah9aCeLfoRhHbPsQ1YVvy4rjR59kc3Kp3xP02qUzjtCLFu
KaqDYMF9pgc8L74GBuo8+Jy8Cz3FJPo/rfQpoorMKEzZjCU68HPKL2Vs/CualUDe
YNEtsH5RNjsZ98NJ2+dAvZiMpqdtHFvV20HV2VXgucSNx+lUrSa47NUI7ZHDAQaw
Jb1XOUs6UquKy81+x04mghZ6rUDwz7SZP0v9LTOhtf4OUBbsW8QxyIrafZ41qdnb
tk9vnzGQXdOa4omOjznF5MzAHLKf8cdRgINAxKjBzFkqrZF+wLEyXSgQvdtLH40N
XQtK2NW3xZYj/w2jf56sWPsbwqs/52VzxZuCXBfJzVf5uj/ncRihirjnF5T7MhEQ
U5lvKl/sgPPIyC3oQXWT1LJ+XXkkNrD2UScBHFGW+NRrMHFnFKLP/23nHi7XYDQH
yTEym3kDPu+6fIzXPV6o0jFlPWo+KX2cUItfTrpdPSfHnFlgscur83w+nLi8KvoH
a16QQCyXg3ROoHocrY4RXfDL1poo4nDgcqkmAFO4qTDPkxdD3LXT6gNB6b53CXOt
lMTgVOVI9iX/k+ymSTLUs2kT0z9CHhXpacS2BKUURdelfzy4oLrTi4d6mA7/3tri
Atyd04MjyAOlIS/dQwtgWQ1gd1ml6xdp8DZ6FXi3qtN55L9qbUn4vQPltpSzH2NW
JedJ4ihESqGg+DV32jKNDKfGhSPAvKLbWI7ZlGh54tIhUuRkMhpjKf5MYNnh12Pk
OxcKpz3xXPm9Po+nsdBNmYvGFmiKXK/IxQx3HYiKzKCVUw/Z0vB2JSJGz8pnhvVK
BKIdbqT7lbhg0m3uPn482A1c8A9jmojQb8sI5KVd+j5YUDcsqquUTbMbALZ3FNKu
/mlcYG7A6YnHWEloJ4dJes0lKRWtQMbsUIJdosMEMaQ6Jxh93cMixGVlY1fTPa/C
oUHuLhof0lD09s89krejg5bVU8URABth9Iyb3isyw70Kkzbhb6kViXHT6jW/Z89e
/p0/xX+dNonMUi4pUtOHrPe/tvVVvAmaliNkBg4FtNZ24EbPM9xi+gvApxCRWmYr
ssMP0Q6rY4DB1BB5Fw53NfhgVF8+TIEnnoyFgG2oBFi2yYk75en78qKaagIG5NyN
dciKpvUAGywWqowUZc4E10jLEPLfyUdm+Ft6B1vFbZmJOMeaThG9ksJNpbd6tCJY
7PlIjU8lz7bgEC52kxQrK5d8tdY2E0JniZi0jO1Fnh1jGqeEZcF31bMaT8khAmiD
h7oTB6P2FQUQzl3MEqKrOujLv/lEh6hFpnMV/8YJvOBxEDT81HzctPhBZQOG4O+A
dvkelw/7hyV/lwM2hgrb8NcL4iSfkJepeIrFqATSyl2O9kEDrrBScl8B2kfWNmdi
O3OxnhIJw7Q0ZTqGheVvAE4fU42sayUopaU4h4YSmNqvW22Y7CmYdrjjthVNI5FD
NB3gpCWMvRAT0+BW2Vp0cmzZHpB7eewx4ZzyIdk+f4/+YS4sI17wIcUqqiyIIGhS
JNuuolk1qIF4A7xMboQ8qw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
T9BMVgBRZi3ovDEcNyCeNpuRUld58bnwUEtmCaO933PMyq/9zyq/HbtLGz0UcNYx
23doFCaTdeIujiK6B2yBZJbqSpuoCZomdxMWOlN8wdLaCGiv1ns4gAaDBCxaT/8N
iWJWHE241WKsGftpujQYm/MCeCt0hzhWMNdAcwVUwhKsGsmP+Km5WeZh68UJ9UpS
ioLD0PXl7R31oyQx5FrOuiVhTVMPyYWPtkmt6XBycLArWrJlpbBCHlDhM7k+37Kc
6tFxjt3LdRII+I/zX89rVU0ge4R03qzBnxAhQzk+KNut9w04cwWOOZlHFQMrRqT0
NhU3EPiW5sarBN0jVTMG+Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6560 )
`pragma protect data_block
xaIPZWet/kRWeQIZc/gQRjwYBoUSTjQ3YW6poWZcClTjE2V6molGC5LWj3B7Io0N
5flWc+RmGX7z9UpQ4yzwouq9fwv/RztL6qhxo0GSF3KwBWL5BMNEBLlo4eEBPKwM
m7I1A0S6/sBHyR1TBYzIr+RTZmGmq2D8htJByszFBbcgN+p3t/jmymH+n/qMfrhz
YCRxbSDSTXmrr2LtlURyFSUosa2+2Ngg3BGk1zN/1f4R4HQPKmS/egvNy4xjRrp2
PNJCAP+MgLsmGMYrDM5fAXY3XxezZMVPB8nunZHTi7uvYdJin5yY3MkBD3Dyio7E
Y6ktm4unUhOUsN7zR3zGmbG7b0fUQ4eyFFNedJMa9EaaEdGcSe16Rv+E+TsWlWE7
JLswyiybs4J4x7VkglDEknhZn1c6n55Jd3VhZvPseZcZQZeSDnHzamKBUx0ppYEg
0O0opNr1GbCzyw0t9IYKBMxdGjhfRiXi4uDDBJ39w91NB5wPIosNMTlgNt+bCuRf
REXjVO7c6kbpSHkO9KThgBNF5sUj2iRymXnEWfPtu2ZT72tsMVRO+Yx/NjcnPvoT
VKkA2ozX2i3dlijpW5V6IbdOlAGoaRBFoJ9egjUryxO/3nh9CPAMQpinAc8M+CEc
38alFuba/UIiv9okq+y4fUF26G14PfX90Rs8HdxvV4r/WWbKJygD0jRiG+YaU6rf
F1tbeR0y1rVp2QPULmMTGUXuKqREOTrway6w7CMIvIi6+ffP4kGnNrqdrLOyrYt9
h4xyd497ddupAoYZ5gv4/4CB4GgcEl+J3O2YIHN+oERBdlvm0OtWIcepwaK/+hAQ
srL8tmG6zvZla1+gkZVkBJ/669QhcqIU6o5kusw0dIzkWFEzaG13jgMB8BDQ8wxt
lAe/Q3/DbNg7Kukr+vVj+b2ilEvg/7YNXKwgdJOUw3NzUaC9USzIvZqchMhHA+FK
EP/zbBzFlEwy2yWT5NoTc2v77UuJZh6smGos50qd14wEPYRIaBIwfyMiHxQ9pawK
FHw7b4I8LdlbBjT0uPLIVCOfC9Pmty5lVeUBeojvH3J1kQj3Pggv26ofPfiGY5fM
M6f+d9hrdjy9qWPo4tJTqHpKNQflDfF3gO/RK9tlCODIKHJItDAUN99BnuLCZ5ie
4/w+xxdblzjV6dyZ4jMED6tP3TYyE4CfLyGjby+93/KVvweDX/fKonP1RxxZgHXk
k8SNc5vrZ9zqeExQAeSYYkYsjvw1AaakPeWfKLdFcdXVn2v/MsabW1/bWOxYD8zT
Tebmbs4+r68SaLZBj+w87qlN7wCwfBz8XaNzJ++WfCTa69RuJmVbyq3n73g0iiDf
S/H1sRyDDmtqgPXpI8bNKXuoKagGSCQB6DKFSSv36GUm0pRoAxb3HxlA4HZncQqb
iltfV+ZgdqEwa4vnooHnjKW2mzI1X6nIVDWTmoB0EERBw82yiZPs9gLA2lrTrAbu
s9DjPMZcrrVDY+oY0Q3bMvBCcPVC81twONHchOxoQhEmK2lShyOft/mhF+Y0GvjL
tZRVwtuJutqMymrMah7t2pT8Gdr/TT34uUTBZHEffUS9mdsSDD+a8UyAVkYntqTX
21jnZ8qKlhDWmgHDF+D9e8xPzBqpBTwYcJH/NBG0o5Ctg0G7GUyY0QVOsuUdMGVF
ZxLo3jJLuqnVFgrF4rfC4TNoxKnPC7FCV08mfA66OL4LeC/nch/RtXhiIvR2UmGI
mEwDU/J1Yvw46Cc7tY8cdub1P0g4cFW8+PCDXCUPnQGvKJawFX+epOZES4eLJN0K
NQ/uFIGRNz0ceCA49LMPbz/kCzgdx9plydDj5buy1H8dBDRycqC99gnwTjhAv/+W
8IOyZ18HhvZ688fgwtJOtrhRMO2oePV6etoDK8kPw6c36vOe7JDnzA/xtB5NCNGL
7BHPsQ+xGP9KgsF6xh+mShArJ3dJZajHaGIHYdtipJtsNaRvLYtsgRERdgab3C6C
7RcQKueOjQqhpKIRoM+ZTG4u4zJmvNgKDgrqWZZObctrAexJo/hrLT5jP/J6/Mwl
aBAzwI8+BV2JDJG+tzwUPAM+GRu1u1UNMdLFemsLJM1O2pTuO+58rxoYXnG8z3DZ
iwi0UfIARyOQNJq/SdJeHVJpaa8r/cpLGSAMt+qMSobzZA8n5CL3cQKEytoBnPHN
Cz7LHygfUPhm/YGuwwyl6/28snAIt9c/zr1s4MbXEvxAMewaaiq3CsnqddNsXqAU
z1gVQdHW5NHrVzJ49VkJc9CQkfukCcphyGnz7d64Or7adkz1MEyd6+ihZxGiVqa2
6zpOT47UDfDgXZzHWB2MIqbNXVQrj7VqTRLmqE7q0eOF+vZeN5kKsoWLtiIXU8t6
wKp5ExtjAyoo7HxIUAqmVIgYrRXa7lHXy4haiiveWGXjMEd8nopI4ezxbS8i60of
npSZMlWHlKukW0YDfEUzulQHJW+GaO/c2WfNp5271XkbqIQ+GBIPVPhTo8qLqKkI
4V+5y9nRJEKn/qNUfkz6me5Za4cJ9dd/qJKJz8z1M9phHds+/WVPLD4Cq3yTxXWM
ow6V63owEoXhudLEWMJYXpYmJDrDeWUcZIYS9Scv54UuxciWl3XE99VBiX7xDy5N
qMKWuOh+SdRsq+OmFddbZLpNXevet2c/UyPWadPyrghAnmO4GE4apvQwPnIOwwhl
pDGFNBFcdf/IFb3lNXDhFLZN5EO1C5Y9KZ1lAhXXrcRz+7ZyN4GOzQdg/TTTxP6j
7+0E88ZuKsFX9Opw2CWiyopA/ZpeDMX7jueo1ok+7xjUolwf+Nbk8qgCuH8TFdGG
CY/gKYSTQU5Rzxo0kIexGdwjqUFWi1EQrKI24jKfE6cMMMNDF4TXQ/MfiHUF4+YL
Dp4r4ysJBRqeUs1r706HuHTdnMnZv/iHAmrrNyl7NE2TcAx1Sv1lXiShVNwYJ47X
M7Yd2SsCkWml6Hae7eMKubc4n13tPCAk7oO7stPwMmO4a5i8xsZi5JSqhBZoe2Gu
LoTqZQGLmqzZHelZFniiSST75QQZreDMpAc1JsDzgTMOXlwtGdkUf8/5lz/MUviI
yS6CyLv2pAZlq5ujWxhb3OU+KJB7qo5j4SrsZBFy0xMDpimnRZYI3T/Tbc7JyJPP
RGCMFQXrS++Pmz8lDWPiGvCs8S0h29Vc6gCUHju0SOmwkC168gT4MiU5qNfMLZQz
Ddois07Zi8cQqLrIw3qo2L+2MnFjJTqb2Eh6VltTCZHWh1q8n2jm2AFWPUgO5fP6
nbfeMDe9/RN5BN5xTOAYWXGqGAXIoWnS4daRf8SUtzeWGTJZkidEpv859oW68L4v
mLYAPlZ1pkEARt40DiwQHdJ7rjyM8GNubNkZVmMcd2ERGumzll6MS0OU4ciCMfLA
u6gy8svn5Y77PEYv1UPWlDUtfeAbBNew0qLr1ZEJLoZN0FBSeVCZs1+Km6uVRT6e
mcGx4bMAaaCZ+JVbfID7/Vxjw3f74Ybh3BoAfZrbf1mRniE6s5lDul5YuFhrpidA
J6LjG8ZBBTDHqaShywPd0Fnl4fyE9KHhDyCMUqCoxwKTGhY/I6qRfv0kzd7xynt8
gxDW4ok0ZfBoin59nS1W7SHjQ5+j6VRw46mNXL3fSPADk5JhDzJlmIpywYbQB3v/
ixPCn8VbOJe4kG6kNtMZE8n3+RMTBwh/8By8st4NlIfgfP3HFy/zu+8ofiFqYjwS
uZpb7BDKb46BLCe/8z5qXCYuIxAgLs4MFo1M3O7sjPsEUyw69YM30FxN0FrM/P0D
95qDLpfntVW8uyGVhNH0WN9x/FZM7PzC8yejZPNQbt6FV/c5h3fTRUbANRf9Q5o2
+gHW4bnsnGCCs35Yr2SAxyfnHC/PIU9vU4LVB46aHqIPjx1vcPPrfVscrev+O19e
djgYEo6TCkS4yAqLo50vl0dmZzm2cnNBs47O0T+tzFHl59UJ1XYgZetjxh3Z+4FW
YLSIcYd74cTDo3gmRuDaXSQN4w3UK2wRrtq3iqgY1lKbxMbWE0kWDqgjx5ea6ytk
c4blhaFz2uEAutMoRKwv+ED0rZqSX4IFzOnLuavqEkIRbqIWUMhyiDKBIVJWv4uv
urfV0v6pPA2fUL+XPZSMpQ4F8n+Wct+rnDpZaeflpfLilCSdm9YHF1gCCrh+v3Qj
aI/RMZboXSOtj1IFz0Gw2b2zO9PihfaqD4Hm6F8owNk2p4Y0NOUSgJJp32BmBo7L
K9iWF/RMsPGSk78n7+LeOSRxX6qJYffAYUuskjIXtyU5pPBP2utl7fFrNlFqFw2C
Z6fel+wVEZ9s8p7JQLoqYSZrSJkcssY2g43Fn/HA9sBhLy/81zUiuR/PWiqxhpWH
Wy2BmDyT2L/RDO/sCrKiZTb4Az6qp3VR0hz+Ek6aDcx7dUPUMGJ+VFTGRYq96rcs
riIcRya1Lfmwot4QSv+ewNX+qUsth12k0jCcFlSnft5rDXx+qDQcwjpM0HGU7I3l
BwwckfNtoL/1yNv8pS9KQ4Wrx9Xg4i35gvZBBqW5/X5XihFtVESGj2H1x1XcJSVf
Pjhg8qgkIryY1TeChkbNjiY/AcNLbAzvUOhuw8idiVmAZc9+9i6xnYJqmOPQ4u5e
r6b1bEAiYmoI6/dT41XBbrbQ9Rzs4aLXIrQ2xfp/FPRowM37FIwtz1+ZGB6xZ2ks
XNuOzUkALLYcTzeKS5QLLyREeRFQ9wJOz+Dj7+s850JbRIwOxsa5Za7ppgEtfs5v
rxAUuBima8k/aOWF16Tpo6U2hAYWnUzzn182tv4wJlUIq8f+8sxSevk93IVJLPLr
Le1exCUT1k3xAIepB1D8d0kH/rgg1jMXg+zjrU44pGWlfuScllAAZ8wLrdhTfE7I
gthB5M7BjvcAvIRfJADxyS2JDMFDrXBHwz2FijvLtqns/j44CgmYKyoDtdgFEp6C
optK0b/q3qS814DpGbGxrgnXlGvU7oDC/rKgaHRT0+zohSKWnlOHKB/G9Unc1MbT
J/KsDEm5xWGHXhUD+Zr4gxdnOZMqFMfR/ZOxZi45FVx6OYsG2R3t2XVrTMrTeeZG
UjTsNpyoFUoxL0YRKl2nEe6JVEEh9IudTPMv8ukaBGD+2NSTlnTG7l8ek1pWHwTw
oKvgrEnHD6UhHlZd82lawSwjUH7C/xlkqe+WIUuSkgUTXudkMJj5Jhn4uVXTjTvT
fQCXx6QWfc7QtHCDn9u+f8PIW/nWs2irgMeukmKhJg61YC/TCh7xXPu4mcJq+ynL
xsOOoQBfzUDhLa0T0noIxAesEr1MJuaMovYpD0XhsYEErdkx54kh73cGqI7RII4L
8CEZ9PXCJiVRr1CA7O6KhormMCC2vwUgsYtTrqU37q0K5XIYf7HQJmYQlTw0RUqy
Im0KU8uDPQejrVML5z2b7p6JJe7EZ25J3oXfOI92GlxqHvrTlvE4X8/b9Yo3yYhi
cMJWaXtBTR8OahcHtVWl0PyP20eSw4wKJQaTF6N4V5pEwHyN2501hwd6TFmFL0DK
cFikuzw2D8/2rohe2UguYACtNe6gHfMKKH3unn0y2uKmacGS+s/49QdDPo4qGZyZ
VFbIJRpY/kG1Xgsh59LUm9fTocUetSTpLiBPExn4ZXOYhzNAuF8/8Atjhc0BkzHC
lOgl8SMGrXx6fmhtiUNiMKJBbXG7qvAC59bXEryMuB8qmeW9b0FVddYvKdssk+Hn
hIikRkH+6wCr4dcSpkqsV6DgjmZwWKCEG27c+r8b15ridyYwUX25pnAuW6AY8VeY
V73D/YCfl8NUrcpcTD994U5g15j6+miOtjQz290E8v6wBtWl5hd/aVnfm1FbqUGo
rYnpL6nY8Fe8JEx4AqPRy9tAtNw3aKpBjimGyZHDn5utvBN5JHUYBfdF0HcKXNOR
whh5Ruv7sYvvDITaOcLPpJxvmyvXKukIOAajK7HE9a3qfI3fcKr7P5G8dfYfA8DS
OF08j3oVbFL6LAfC+li1EETs00PV6zdYPU9HAlBklK+F1EJjORfhhTvgHXvpJOd6
Vrr9FfJe5PYvrU/ooDgzzDyTnMb6KH1lhb4Klx2S5U9xJNMDrdFgza5CC37XhSMg
nz1dIBE6nQBOh/w6YWRAQaTzOtJixYrfS+uFw1g8XEEOrxJLJGuZug1Z/vM5P7HD
rV7LSmYXhDUZ7uP+6NxEmSXjsnVM3mydfrsDNdBeOaCvyNZk79xwtk8sSHgtgopj
XSM0VR47ZBGZItOCE5kEI4gXjAZAsevazxHtar0UhSTWnO84STMn5xcvGHdU4jUf
Qy5D3bdELo1thOC6xCWVpdOAeu76NGDbZHJhiNflk1zS1DJDqZ/A9/YZPr5IQYZB
aYOkExHzrwUJmlm+73pEztjNvvBvtMsBiqYOteSb+xaNnTal2EpvlQn2MTrKHP3K
MV38+vyXPeOqtLTjlG1PC5FOmPa0kKGT1XTAGHFVW+IyAK4px3GMEU4Swq/wvQX4
w4E5s04TEfjZMlO57TiLjYNPhu2a3Q6mwIziyKOOpRERx0vV2lKQBoX+9T9rpBuw
o3IFULQwY0kmz24oXNxLCJvala38pQwy8qq02NmTiS/c/GHOBw42APaSUQ22z+Q6
VEubv+M+beU++jCvGpa8NKAbQxsXomVoGTUtVv6vVSoQsJx5jJcaN/Wx1EHpntzS
h53NVL77gVZOE4bjikX03BfN7WxBAbe0sEg/DmGMiy0FGqJE6VsyOVNwsst/k613
qhVCHb97iIXD+v0/XTi9cSg+6hPQETd6lOIEt8O+8slzsIe5EhD1lLsaFTFHdiIo
gNghduuUEodX7KLddXCfegC0QpVTNkWg2wVJDR2UNghl+6eDb2uvSOX6067/FoV1
eXuSWr3UUAlghwvDH6zn8NtgXSp+0I7+ZpFFMP9WO94rk+M+PPNRXsAp1Klk+coR
aLrjDxSl/114SDFCwI5DPV3yhFdspGz7DBecvLoZwgaJHmgQOMBbevG+fRWD9D52
oUqsLjQK8lIxIzmvbSJFcClGI6sxZd1cX7qdPhvXGVqIkuHYcTmnhuQNW/WSevcq
TnP9gaJ91uRvWLQAMP8TPcn6jR8nS3tLbEMypGZsWdjmFQ4nVzA8cCVmuq1FCTBW
0Ki4lQxHWN6wt1DlLM5qBgHsgvIe2dw7cIPpQJXqqYeh5uZdU5l4c3lG5ZCvrTsu
83yDoDXD0X/lUHRycQfxHO02Gaadau+8jDis2GIF710lwLeYACEnqxSr515OfsBJ
fS6bUpaQeEXkkZaUfrRI2azfHJX5sZ4F857gednRCuOe2A3DoENoEyaCJ1OumsG0
Vk0FT+xUGng0CEC6y8LuN+fwwrp8DNl8YZbbiskC93/MPEOyOmswxK3prKXZVHlS
/HQZEO/aahwIhMFC55+CviERDZ0SG3sloRB+kXRkItUyqIOqeV7ee+hLmnwK5+9Y
wUEpLTeUXknepuSQEBfgAF1Wsfn/JKapJl35txUY83Gf3BUS7+VCpJNJRqKHZeFN
L++1Xm2poUz8lKCXbmcQvlqbrsEmgHZQn6Iiue+zVGAISL9+FwzQir9yAgxccATd
XCaO7EjDK6tR3ScsaTasGZLXMlbqmHjUwjIP/p9j1VkOo/HefvJ2SqerLw/K36/k
DTqP6GFfY+idXyu6T/HZJK3rlVtj5ITdxFfAkt6jKKpppNqNVxieX3FKWI00bsfN
j6poAu94ow9u1Fe/Mjr1a6JRgMspEbd+SYzBhN5D1ztasopX+p+guJWyrQ+tl5Wb
vviX9gdpTZYoNrZPSTM5wOTjoYNHhloU8ObdOZSXvz5NC6yeBxhATwdoZstmemJh
KaSfzmRFg036QxcLpcLadS+AJ4rljvNOORwAQg1P60B9nKQfszpF7/3/Xr3qJr0W
92d5+xar/TXFZNMlvAZ7cVbZE6yofBrwaQLzUW8B3nOSS8dppLQYwlINacR+qsXy
JZi4pXN4TMkzTPUlcMrMHqgZClQxMnnjG3Qc6EWzyVR0474YGJHwrfCCrXdISPvM
3MXwVvya/6YikX+VvYfcOhSDvYqQosnQsEuURukGQDb+LeIiuipwaXu2//qU97k0
6CB82uT1KZOFvNr07IzF0UHxHXEdlP2GMIDl4qsbQ3LtMdecmj7kOmm2R6/rH3C/
MhJfKfpwQ9AU9jaLFfO/zs3R7c/CEhcxatBPXEHLJLjswT14FzyttdiwpGJVgXxC
n3ylg9EikBGRrXaBv7oVazPHYbFR+Ll3ZNjfZ+9KIEkLtOIlj5jeX7hEFanwscnG
tcjxFnUjQTlJ4baYhkDY+uLkMk3nQGES/PV6JCWsuV6uOQdjjInbwAum0m3DHPoM
JH8DSyEKKd6juPAyL4RoRM78vE9OxlBflFJd5lgif2ARjbfissAXNxjO4krXJVhb
oU/yD0329jSQE5SH+sIZYscAHl7Yus6CJ+kW4lHW9VtOwCwy1Nv7f1x5zJvFZrr8
mJDrxHJLcjRrY5NRREqqUmzI9ZOM4iQpett9b4LEvhZ/0RifOgRU3/1nWvlxIFcW
TJh1Q3Gu/uNjsa867JKb4xYmAeYPW7LJ4tUBMcaKAZgDD52389aL6WNJJk3MriYw
K20dtALiJnu5SurB1q5VlaV/aL9OMxyRCOVVhEboNC2MUGdLWRID39G10nzXTlJu
DI0QPclTEKbbu/dRPpY4KY6rZMzhzwjtg5vNivbkK5PWOs9S8/NeInO1LxreWwNh
QCSpw4An0qhCs0UMJvcN0Ws6r8QPKFYj5QY6c/qxVFI=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
VVpcslns9Ei17EyqnVWqBXZYET0mczcqCfLGhVbmDFQkWYqIlVQeG0kSpc8YoU/t
uLnbhUJbyXApLWsli5P5V1B3HGFl85K3xJup/venuQBw1Tnv1W5U95aEkKO3iD/S
WOoKLe7RxTlXvBAxPi/j3W6KDTV3MgjLtmupmR1ol5XiiEX0NNABsEkQf+61DuEh
3r7+yrQ3eAKwnTDXvEB92IF4JPtlkPG7oL2kjvD9C0F2y+koDvFTcEUh0eCwIzg/
DNUfq80zxKKQQTo+Nylk0eHitXJTgdbVJBdsrJdxxRXsKwDE5png/1iCoxEl1RRF
i+POxoFyZOL/lfJ/fU+Ulw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8928 )
`pragma protect data_block
tcmQ8x6SdBPORmLVket8Dw3POXO+1rxzEbnbJ++OsHc9xw5rl4ZCu/DOoUj1+nIk
lWVzFKcNZWU6eU8FNA3VavnergZ60tmWgzjNabXnbkAgiQ23GUP8wY4+JYUokkFt
bFOvJZ2TkMPMLGmyfFqM78q9rQtGtuproAcQ7kvt2MgkV+imFPzVtK5u5U7gM0ID
5r4/pFDDOC3trYf01pmtjtF9x/eR/Sk3Laxg1I+iekimGz7QQoVV5AvTjE3PZjTV
H0lHUpKfxLkm4dcdQiUTPu2vPfrsEOCgRIYRrWX22p1G04TeEy/bO+AkQNVxYxbc
RbgaaIKP5ubvhZgyYNFUa0GTSmM3mtr6jpOA8OeiEzI1RtcryFE5g0lXuKLa8IeS
IJgfR/+5cw+mQErfBhvwA6KisvC/NCpbDciz+71ZNXYZxl+bkZoyMIwklSRzAVBA
WmmltGfXAW2GQzYTmr3Lky5/PRyrp1iLQ5ptMpeQ91+/6S0HLqNGhXfYT3UZciEl
B4UooiqX86RbJqYb4F0OJ6QN1C+Dlz0YUgwmOXGl1cKVG7rGp3jGMLNyBMcooZrv
gUTNoW7nXJK3DNtZJZn12rJXeILOrUpR8lZcNvapLF0CH7gykyhteR5L5y2Nqkxe
xzWNqJ0xUPDWnDnzTm8+TK5+YoyKVC/9Kc2nuBFBQ2nwNNsI7tvskdOUzcqa1Bzu
VxEBDU7z37nf4Wy9ucFzNO//yyIppEEX7CeAjoo1cjabc8M63Qm1jq/nPWEiGL3V
JUQzVdcuOZxzmPDRAdhu3OP4Qf/j95Tig2GCu/+eArWPhkXYMPs2f0j1rcr5DXjj
CVxeqz2b75wBi9T3k2044XlXFS1TIvLDir4rtXXdYm/VoDX+sX36Vsy1ZdkJUO3D
/etC4mcdNgvK3wnRStBDPafP9EKzPwD+hjy9Qkv+woHRnxEXUcf0fGHBgBQ38lpE
QbGghMLs/ANBvF7LCWlKyYVVfIXsEk98CpIKPA031KpRFBRrGcEVtuBnV0ddXzKp
f8Wo6chO/sXUGk+6nO/dG9PsBGj9T0S93+IlLuGrKT7NtO6mg6k6eN9yhEP/d6++
PbKQqItbcDviSCB4wmlAJ0zt7/x3PunfQqo+bveYH0nCr8qaBZjwTjH73glEU0HB
8HnvoihhLuN/D2biJj9kgHW+jgcyqgt6YtoqW0b59xw6IcPWMH4FIZYvpzuyINiF
nQBD/z5xg7YvDfQgfOG51zW3jnQSGBR7bPMM4qgh6M+WrxKSfesUaiVTnuZ7mzwk
EHSVrGGG350EUkkyr69xAs0KqTaE8g/QteOq44lVn5Z0reIyhn7yGMn1Gg6ML/U1
0go9i9rxZXNAx9Di9XVYIoMGCvctQNyGEFdyrgU4kpilmhCvZerUgLwv0CUY+WbR
8qkjnG0C9cpjVkjZaxm3hHe3B0NoceV0IpPISgLT/BnqVcJQLMiVlkrWLvPjAJ9d
HV4BelhwdSL6q2u0QoaHn1YgWF1LLOcYLtQA/M7WQqyZQ4QtYDi6PY1zpHy3yBwl
WiCHZfyqS66sc5upRi/Hoi5TDh28zhhyHsRLjoQz33D2TP9dRaYm6NNPluk3CxCX
/vp8buekgjlyaqiYxmmAHN4A6YP/R51Z6PnWm5arDucgBqR8OP2Z/gGt5vlpSjej
GHEnT1Xx9KOEmVR4f4Usp4f3rvAoh6lP2z8/cR4eoEwvRPn2HH5EKi0fH3f7mDrs
5gacS8I+UqHv+41+MUnTIiwlm5EkS/UFevOZZnxFbzSxEji4cGqF0TAXW3dZxEbN
Ii0An1VNr3RJaF+6hcTPuv/GUiLaOUIeYVVbUzC4ek3d4Oi/Xn2RVClVeM+wJKwi
owN1w3FJknfZB5IBa3IyoYbs4HRM0whFVBbpeXb7s56qbMKYRzIDs/i8L+jv8cC4
mykaw9AsIi7WUn+dgdPSj6clI8QiFJVwQ/7y1kFPNUjd8Ro8ChAK+PbG2K4t34OX
xrwmjEb391zPyhHOx841NDxUrvT41OYHD2fqUM0/L081I6ALhWgZFd31W7oXt6vc
sSOyhiPsOfVmnJkd6hhnokRFG29vB/PJtktMnMbjR1IeyxVt8YZqQG43CVeNYYGT
3wJmqU4IdsCBOehR/p8ChNrf9pCs51C1DA0gb1HY2RctW35gSdI0zAncBEFgeKhv
GKefgwJ4DRAlwoI/lA5AEvSQYGt2IdYOg0GqLXwtMy3biYPBwhmja+2PwhJQMYGK
i331TX+2uiFygUWg9OkEazUSHKQgitqIGLR71eI2EKhUuwuq3K7H1ZcgW3KZ7AOz
tmuH+SF87DzpPbbU9zAeZtyL/sbaV7BFWC1IxekedzTon6BPU4WwxMiJU5snDFlE
dvPH84ZM6SCbvALLQmFMv+lMqtwhKzJBDiobI/p42UW9iTyjh0PYqNr5e7JBBMiu
/Kfc6Qd8BkdIs0KHKdQU7XpYo/I4IHQYnoKlfIFazrX6HUFbfwQ0Sp9NweiHm9JR
nkbVX6Im/YBXHq+T81y/iDnxluqv6cOLbLm24bEnsWG7aTZGrRy2RqSO3i0Lb529
PK7OaUUMFmcebW7Mv3vNuOgG0wB8FaTpsGfTUJgqvbKTkDPGBtek/7KsVuYIn0s2
CmRZRyF33AMWHEY2gDZEkvgz9tJIN9/BrhjNxoN+Pz0MTXodRxECmE3SthchOXZS
stJFf4JpDjEIGbkER7WyY7AvqwDTYxw945u++wgsoVHM/53uvCIfwo8zCzH8r0jb
aWN2aVkovg6K7NtZop2ECUz/Z3HHAb1wKw/fQojvlUgbud5Rb5uH1LL6mF/9H3NS
l+nJk06GoCbAJ+1Hnj+nIKi4WUPGhAOEVIHRkaLQWArW09LhT3mCfQtpz4UPF9qS
f4GDD8IBoapmiuMYDKlL0Eio6ijbMh0bO8IbcZsPQGUGrIsKHB1XcABrx84HhlUM
GA6qPp54Nme17TEL6NkL/x57kryT5k0InnvLjBtoe9vZcbsFpLk8S5CI/Yv3PbZi
xqNT/TW8cahdir2OljsDeUkNmTfySANeoF///BGtPHro+SnnphEJCle7B1Ooz9v5
dS4Flyu87Z16JXNrgKa+4pNboEftx8Sd2NHxyeEBEz8BDiXHZL4czA9o8fzc/oz6
xynacjEi5E3OMXLTWJtBphTFELcyRQ+dSNKEKCjTW+w2TEz7H2viSyf8Gheqelb6
T1UqnqPs8cuGT76NCAuPIiC8wpvjRWos2HME7zhzIa0TBCFYyGqDIDX2e34C8Aej
uXxWMzG8WYZjCVm77yIW4b1KCU3CyCPcUYBLhDCHyRZVn3m7qOwcCXB4FACTxlsb
9WqQSC37lUqHqlL/1q6GNS8vtQIYqgGB2GN72edaJg94oMv9YAy8ZyEL7e9iuDKP
SrckSwNPaM4+xi4IlqPIcEmFfJvYfknDGu9NYnUR3aNcRHBXjGMRV7s7WgJ8DdB4
Pt8U+OPe2R94p7n6ZVCPpXsEk2up3mxYb0K8acTNbokQvM25fS7oi7VDfvF6+IGN
tgoyUtb4K6pet7M+nsb7ithFaEky+CTApSgWVA0USwBDnqaFCw+eg8XyB+bO8fXP
8rpL4v84Uh4UFGQCm2c3ht2Ie9+dPFarWK008Is148hHCxxLEd4wEYqzIRuzjvuv
9eMhwbXPc49FXjQXIcb3khm61jUIpK7LlDdag2EuUCoqZMMdijyH0ag/23qB+kdG
6CGK/wdQ/6T7h465mJiKXmLgCER5N/DTPb1VmShhg87bXRCLGBakd6wI+8NKVPw8
aytJWcF13L7uCxTW3wrXOfMxmEVA7JXq4HIznoPnBOaQPoRTjZHyIjw0vYGzWdrk
LONTiLb+d6BUC3FQQD4lJLCWsJs66EpMGQ2PKWbAdrLFfCf/TXVlfWxIpID8oW4N
kfvTdjXwOu2xy713PYyrcaRoU4aWgH/G0879RDHfZYN8QLKE+u9A/lunPpE/QaI0
U1LPtm0OrnIsDtVddmNICuG/kqV36JtNMALgiui0kbKGJHdQNz1b2ZlRxyGfhiQt
a+tTwxZK2vYZLwb2a8b0tiMatpwFEXy1BiPI3QnRxFCr5KXYC0UtPb2WLEY00/N/
7qk/8M8uQEFGcuGb7/+z3nhU+s/Mdbtzq7jlw5IVF6hxQ5k9lQ5mKw7c67hwAjz7
mIsGzyqgrwtNLoyTPore+Jp3say9jnV5GkVIVhF7Bgo0/S9cWHvjNcxsMBpdXJri
5aI6gGnjZdVlv7Yi7FvBtY/8EcW2VYFuLKUZb8lfpG/tKLSS6gcHH+JZsvO8MeYI
pCyNJWm1ZSX9usNs0EWE0aNtSxyCv5FbiodPfY48g5rZDETGFk7p4pVimnanB1fm
yguJUw0FKSOr0ByviJkawK6V+FfE23j2K/5EwY6wxMuPdTvm/BDsG3joXzhCNW/Z
STpB4S1cePpk4VWeXiyUyxBpMdqlalpSjvNhvtk8KMbuUy2RjTNi1o0FD/uhyA2f
ygvZOzW2GMkc6YDRvx3gHSWhPQ2ATVQgAiPjXzPIYk26PKU9fPeunm4Q8RdlpD+b
Vn26pkEkQ3MEm9dDoeXX53OfmMJAZS4jP4BXMeNWTRDoEOXZ1594pfQposgSi+cu
y6oHkJkBS4OrmE+v+8Ap47nL9jjenKMJHll2o2allM0T9KxaPs9ctojeT51wDSFO
Bgg9Rd3hWS6RYbYvYb5xAto4hocl9UTl+L4VCrhik7hiQrr//XCduHlH67kM6osx
bRq87uND5oT7QNA/sJdlgsdKedwEndmwYQMN1tGbMwoC3KCIO0Z2icKxfCEGdhJc
2sS/oOagy7BcvIbm1SQu1RfeCaoJlKb3or6J+jFG/03SqfRjhlnw2k1iApGrn0ag
WIGBLRNwS1cif8P3N+7REBsRMDV7w6u+W7SVkao7PcUrlf3YVtsal22bEhaggOSe
Qlm0Pc1B5Wj1bjklooygGjjnasWfoABU7kXVA3mkkMx0fmWSUd0pehDpTboXvsIZ
bLUe4B3swbwlr9CkvVRijRjnLclbJqAva7K8bpEkDm62bAA4YubMo9fzAKodHy1F
4t06swPvZ7BDSNp9jj/tiV6OJGtbTllneU7f9WT4zetR4KDraojvFTaOE5IHi6ex
0Ct+tfJmH2fx4FF8Z5VtGeIj4cpzAJhg/iXIAXWSqdu4zZJVomgMCyRqCZBgRdW0
V7DOM0sMPZTqAKvNqeaZkxErYPhjiL8p758x7itIlZttwkTMsTaNqhWO8G6tBCO9
2W/wZhnwE7bAchoxBcV/1ock6Io8wJY4/4h+s0SVvrteaoztWHqJdN6Ee/DwjPZ8
qCJKx+ZZNPC9w8rnCnvtyF3q/daHGnpJvBP5woePMOyG46ydtVdqEQ/BmjQ8mAz1
aNH08ELpxNiehgEo4OBHu+K6S0U/+uZqECXE6tUyRoM1kdETwDEPo4Fc05kEir3J
ACjuvFOpFDuPUewE1ygyxixQYqpSbASawfnJ8deLFWtliWyWYb2oVjxG1GuCNg6x
D/PNHO4LvppfNadRMNWPgM1lLi9C7SUXogt0O+Wxg6JnXNpeGR+4ZrO0mSccG41i
Jnw2gKxnAIF+R4SFbCzvAF4ShBtwIAnfgBvel83v19JZbDg0hbZkC8cfFM+eYDY4
ucltSVLKTWpA9oSBdf+MJ0LFgI/rJAl62padZizp/W3YeIzlN0hMiL99HnloTYH5
IT2VMu+sGJKqsBj9A6+9L6ZTmOfFb0D/CrmNAxKCxGvYMWIeXYRyey0SDgXmIdu3
dhYdTlRMfeJA4POlQZ1hUt5eY5DgPH3V40gDMsq2wKuwNAZcnNTt7RLh74DQ5EFr
P2Br9t+YsxAFtLquHs8nsY7DyOOAzo+6EOq242p8nKG8jChVHTfNsWcIONmKyb2j
TMx8s53hSO5IGyUCaQXYyYiImQ1HKmwQwHorOKmA3S1MuhwRK5chu+UAyf6WnSWB
/N/yjcv+zb0kZuH6dEGTg/WOLNG+XTAo2ClFJA1uBDlvkG/u5uPgXRamkNIZbokB
PM+Q/VesfPwOZrXEh3y7QIJ5vewY7YbEc09bNVq+HL48PW9Tt6LBwU3BR0NuQxSn
4/GKTMj8ZYVzgtymlXh5o7wGHFe44CPmt+bANoACfkDLnLKip1xnOYF1tWIlXbKK
z79i/mFyzADEmvg2MmD1++t8xAZPJcTyjMMOFl8xaqSrVS3mi5dywS8GcmgbS4fR
ue1o3rEzKw8QRS7PU8bx8EyWtbklZCqvrAHib4TylVRtxdcn7e1l3oEwfFvJnsyy
Y+5z3kcGU3+UUDHH/L6l+d2ZuA38Go3kD29XqfQ3g5jWSpxJCAKOygmHccZMLHLA
8dwkue/olomN2+y2utRMBrQGAOmKrquwJAP+j4fRzUscFda72owZ6iD/HPZ0YqMg
iooqU7e2HOsPj8UPU9WHKxZdzRWaxOCs4j0v/11HrsHtzxqRVeAoTHswaySaAL1q
buRKAECEpkfpGCmqG4AmO2kjyAb2BVAj0Av+OCU6QgCaumpz+Q/4Vnl6Yf5+oNIf
yCeQ3KM6wTaZ3KXA9DWfZRcI5X0e5DPDzwKuyTokI0xkAp5LLBlxvNNm1eYBk7l1
QiNrv6ZdoBtxwMv7weTVn518wkf9bY+c2sBe2ZwoBFO7uv0sSoyZ/XF7B1Tkxl9i
uASXQK6fYwlnFsmWZvCVkSzodUAwBLRwwwSTmusnatCOTG48jdO+5dTDZ/DW/q70
Q2eccwGFf18XbCYzvZheC0OmzGz8BKijf8Vffu1+YEPlA/1iKahTNadMluxOGtpP
EJzSdvnRxdxgGaRAYuSZMpFWQgl9F3PADAjwCtCeL97c+Rg8981ps+5bKInlOCSO
s/ZzUBelDDXh8lUd0QUXUG80Sc0OAYwz8bwvBHaU0I9P9NUqVysH+NXeRLB7schN
So5mwPgEBS2QS3J86gYq4MN/Ae+TK4qCyxYd1dstvVjnC5uZQjOhx2fVPKa90phb
4lsDbmLW/QWTjKivRMgRTuN7fem5r/eiS8RhEmj7TKOLHMsT1mvmgG7SQQeYLYpU
597vzlH9gi6DAOdcrX8LvBfANwjzeOV8yFqAUYfmDATQf2kmCh351kD39kQdzPaL
bIj7DKiv//fL8K7DYABN8EUqsBnp2ZXa37sOfVYyA/R+najB3in66/Xi4F7ZGhVm
HobCcQIgnWRDQc3sK2R407T1oUhP7C62ggVjCQ+kR1/WstwY8kZ51WwOY7aH/Csy
Zcj0ExGHjjtP5JQc8IHn3E1GGuR7nRLX1ZYqb/GP7xcaft5Lxfl5O5GL3Qu+9eTF
ZSy4eJrsB0Do16SfeywrEBlfrwL/uSqrqTf+UpR58mN1ybRrIEZGyLLKb46EeNqd
jiYJI8HX9a5LIpzxVx04H5g1YFlbodq/zYCgIonai4dkCY12Zyt1c/7X7iGp0x0v
Dx8iMpCzw35Ls6srBUX53hUsBLR6wTM+vjzkPdnC/jOki0B87S0A94NvBNw2qJYi
2e0SayWHdtDDb3WBhgfJljhc5nGqWDS+x7TjPTm30bUC6Ukjytw72Zthz6FopJh3
4NMhaA10bVD6nuwW/XJGMiljQvNcTXl4UIDXZmRwH7Kcl2G7kQQJJ4L0uuWufs96
uapKm/L21Avnhy3iwb9OmbGjA4J1+dubx1jEJfj6Y4TxZU5dc7KiDSNdBAse5KB+
25s3eTieU6ZHufncnTmQ6Ke8u8W4uogTwT1TeIX+9LUcjVapZhOF1aFniv2iB+9+
L8BjXtTOAQdf0HXvY9lUsH+98MqS3McTwyTLhPG97VcEVrAmcjkeSuCqg4rPHodp
rf51KMpVWXIbEmqmga4s94iQyHL1d/v1ebqNYzl+LAn1K6Yp1eihnOQnX0e69utx
Fo6lo/tMOqpqb61GevopU52cLV/5gMz9Yn+MUWV5k5qofWgxO8B1NqziodrFxsMq
r/HePQUw1DuLRiyVj/V9loZHVEWYO5luLEn4IJ7FmpYHLZ6zDMRAgpb/+PGvFCjt
ZOU1q7Ip9U/cjLgV76JdP08kqnvdwHtzd+rQ/RqAV2Qq1rIOOTJ/GAHy28NPw1J8
CEvZLCcDfdYN5B24KypPXb9IMjpRrvVVMr5XHEr96jfj2632uEyOxL2GgbZ9VhuV
1HssVwn7LVxfMUMvYHHt46JjxgQyvnHHWMejpBRWC93pk3kM0fsFb8tm19XccRs9
wGY+Xgs/7T74oHe/lNyro95SRxu1UEInJegokZgsMhhTrR4C45t8Tfg0qrDnBtQa
DvqMBaJ0HvG9Pw0wVFfC/lFr9MUGIkx2PmeNTF4C/h0ahTE/DUljimBpJR3ouY8I
IOV49R4syJ0TCIay0tevYglWvzQtKWrLcKsDCVpeI8YIsEHP9/u0MMJ+TeRY1Qze
rp6io1MQHz/bV1Inz/SbYbXbdaWl21RnWrdTX4nnSIUgMj1qTytb8IzN/+/1d2wn
CIHUTZ1IQA1EiJt/A5RyaDCxwuTw9cP8nBKaI7Ft6avNvKjnwCZvGAMWg8STXob5
twScjvVg/DEr9DxdnmCUGVaiFEBqmZDffQ/6Rd1sW9XT+WnvQO7lDkJkKwV8Q/a1
JaqFH0sPqQAlCWrr9jVpUsOTFeMw4bLFBDNClI/wIAYp1QGT4yVmS03fjrTIn6Fk
s9GWCaRmrPM8kC2G9yFdMm3uDfsmoOBDGYrgDEAw6EmS1asnRi3KAw+cZ3WZ5n1+
yVHGwCdSX3ao+cXIb0ACMtTuktOWKW+gDpTy86BjfmKjHIfNA0LDCX3OXPkTGAP8
cnrNw4RySxtI0quim6pttCbY6IoyZqPutajGszec00nR6FirvO3A8+E4py3/MTai
X+bTC4ZBwtqpOH9ycAlxN/BlYXUqE2AdFEU52gBogKg4jJhxQiGr3wGuWtWCL8RO
Ogy07/YxbWiwA8tDuompav9NABXaRQZ7JNn8OjoQaU5vYpHIxPM62oPBXXpvgmA6
yVdnjnnd2wzGIGvDQaUmnxE6TEhMz42Z94NvHl4jD65MvBGKDpWMSEtFsiTXS0Kk
2Yvixx89dCVOeNANwYeeRsv2JShU7YkXajPn5xOwoWE6wxvVUhgRjiG1E5jKwgSh
ocZ5wMWYkwTmIyLq3Z0pkGYMFNiqjThbavP2v57v18v9FWPvT2323Mw/u3iLw4f0
D7tpXbYy4/o3HMRbYSZTxuJgx4yVYZSH4xB/RP6/gndtOb1GJ5Gg++7s7yrmTZfK
qS5Z7zThrZsZHjsFSb07jDNRcklHVX+0XeJ8qdAQ0SNhVqy48CZfaH7wgOjdZxVk
CZQ8IiWtaNCI682iw99G1bwNsusVaqddUIwhvH3qfr5jlUUKUvUNPQuT8LWJQbiY
DtKCD0+kXOCX/5iT9TfsdizD9YBt5d1dq6SxTfGO14/KadIi/zjblW5w4EzOWuej
Bju29TRAlCXqs/SM7Pvkkrhdg/BhjU1kADQVouijR8xxfNKQnaqTKWAwIvWhsfje
oyPGyYQUjuU5O5aWiHxS0mVmSha0H+0+3qPcES+/JyDfbEoRsj2EtVbRDsdYAE5t
LNP0k+yDPBzh8ASkxG2niZI2IhdZzXHg6IiD/hmL8wViiclGaXs7KGQi45Pm96BP
EYvIS9J9XIsCHJrNU6dHa3KpCuL059bZMUNOeaCPM/sflhKC4+CVIyLWmpW65wqr
amNkA3L7Ov1tPtM3KVBt6v9l1owwJq8eXJrbWINkoSPEFILFPKvafxzVdOSY3Jvi
1Hxvf8/FHKeamaWqlZyvV2D0kFLhwMHC7uAtKpOZoyY+UcskKUsOKm+NhnTJ+i8o
+LmMjUbAmH32BLMpHQwXMqjnrCqVJO3BHveLyui7nITb6Ate8u5r+K2G+JkkqGTx
mhH9SVrmMFudJhmmOZHTgn3jsR9zEvdYqr/28TyYFrod1aLY60fBfvwrRUhNBl+j
qOVXSqday2VedFlaC6+nsmDxOPSWs7MGWl3IVXQ5CTYuSwXC5EKysvjDOafStcNG
XBU5sn6IgGKg+3W06aq2T+YC1SUpbdbQxfvV6+m6qQN2r1Fl9Z4ilNaDDikoTG9R
zRTD4yD+e3fwxPPLYKcPiuKeGKs3JHvwU4G1/HsE8AxNiS25kLAaJZAF5IPOsJFJ
4PAmOrN7xnzqAKby95VFKTVKnXRluik1Z1Qd3qU9DcOIRXcZoOdN8Vm3oBJFAbpk
dDhl08qfSJSzy7ipjzngz+LiYDS8ojAViScZWFBOKcwIdQBqqKaXU/E8vWk0Yy9v
oYa48mN4j5jDz+ZJCOdEATpM8OYhl+ZIVY/vbADJvgtoWQIjlkrNuQDWHdt1BGjq
zBsXEi4BBDP0gdD7ZJ0pWndeJw44BkQtgECa4aIysxPyjb+CsUcZtZs40j+PJ0is
s9ZkFrobvbpscrvw1Jrb8l1ZFKBmRLVBoUJtjrMnSbtubiXqKUybl1OHb642gNGV
eyf43ixh93xRBCwlv8XKa1n5zVLDrAUlWwtpj+ahCYwBFSSwy0Lw5IgR8SY4BTiW
hDQ6/ZnVRY0VwVJTO4W0sSyfsZGVXCVxnWQYpzjIdWO3GjEiQfbYRUAkQNZ1/L21
w8aDbcYbelYHsHqKSkhCPVVKTjTX7q1BbRptNX63bA1hKApXFhQM0hvmUd+upZIR
ask+veYCMFHNiHzobJJA7yasBeDjTbAN+39kfGtV9T9m82iMaLgd0lEuPsTsOuJH
wy1ISvmKqpZKyirQjnqJKlyRZR0Hkc3d68gK8m1lSin1Q7vBj2cgRwgFEPE+YQDW
aVW6cyMh2C9ENUgojOmKhWi5Vgx6yBkgh11YOjSTfO23fUjf+1rfSr2SxR8pxPhp
wy6DwcSfctLYkxXdVZI0cOr6W2ZcgcgTI17mXzidQL33hDaBgurGkkvlpIQ8qjpq
5xVQ8A2oIlOjnLtdkyrNnQw9B5QQbR4AkenKzvVKrMYfX1gqJUWS3mti0xVcGJsD
Fzj3MOrAW1teK4zGY+z97pAzDkVDQYD62ZBf/8EiLOlPy/mJOe3BUHInDY6nlx/h
ngSgBGscOcYe/BY/8KY/02NPNivqBwr1E+7vX6gSjHwbgEGReinjYxhnBa9w5wDF
KyKM4esG/siheyKyOmct7QHVW9ZQ4hHlY3LN/VfkhiTn9XDjaUZR23db0egR7NcW
tjHvLRpYVqvlOJE43xEf1pgqMb0VNwGP/pdS5HtkyZiKSpayQ9YXTputyFN3/0uQ
9r7AbiEt0aU0shCqBFsvemlSULPLmU5kvzHBwR5FHBrB3+a8pEE3RK4EwgQ44rQg
SzKtdxG3JRsSrDjdoau3S8rJjtujw6QaHzPcAR/5xRBcnW7lsmkQfNZnTnyNsJy7
VF2ybA3lYZpnzLJFlUJaPvYfMfrWy7M8W2A5/h4n1uSpM3znEL72O/cXy16xtt3h
edNlUeJrtJY254+9MCSkU3mWFgJuYrvDESDZYS5X38CNjuUoq2p9SILli7nn/Gzi
5IbGF0wwFeQrlgZd2ok024sUTrFBZG7kP2vQAfxyLi6tDi2x/y+6Biz60Z//d17G
I35CofKIl+FEFDPF6bEeOMcocwoXJv+v6sCA4T3SgIb8MEDvmbAmRv2vAfpeG8cK
1sNbrrnWRqRRlPPhVFcJEMnYwq0LvBqwAmUGreOIKyFccKGmR5XbBulscH6R9obP
LZWWKA46PhACk1KUqQlDrmoJ18yW9taWRSPwquViZK7n8PyNCMrq8XTIdJuV5WYq
U6R5pBGlSlxTFrjudfcLYyTro2oh2SVBpY5myRP6MuspHw2EkgA3UFFnYM/1Blw7
1Tvo7b8jkeSaKfvj7avah+FptMxzNFYIumTtcbko2UfLg1sbVUhe2M5qUwySsYke
OK/UDSrAoLwpiba7vZmmbiuTHD3HFe3fYlwTaJD3dx8d2cWMVoyb6CYjCkPoVwf7
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
gR6sDqfRgUZjH53+FzrxRjtsh4IjFmT2oCyyYuAZzUex7GSMAoHeAqsJEHYSOvL1
hiC/SMzJHorqPehgJZHUaw00ZOshvDsCreVnmqebVDzZjv0ltFMKfDtPwwT+0+v9
dhGkYjm0E1f9ojws9KNCtaxwPHVrA+7wkWB17C4S1S7OpWznk37MJmsYRgv3LviK
goQ88Sj0QZjKGFdQc8JfauWp/3vWQHrXcB0JiEe8OZ9K2V9RTado8PS9P9a0hwIa
MgcIBi+ahG7/iUZLPBeeDvZa/lOo3K2nmEGXA/Itu3kH8RXo5qPSrrNb6GwRoN3t
wNFLkRSQKbeMi5Jf6c3Exg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2912 )
`pragma protect data_block
dZDv0kh133rdf/C1+0jz5hVlJ5Ca9fKPDQLHZyH5XMCP/v4jZczkklPPohwPZJ9B
9hvQ6S9TUz0zGLTawtzwuviU7WlmyFDbJOZU5gfE/v6Nsn/8R4fAcax14BXzThpz
dOkyNFDUe7wHIXJRpP3QiIS63vv7tCMT7U2jAgq38fXSRmyoFaLQlKTMUuZdZK4m
StqHZoR+KkZ/uEF8DBSCBLQkbcLZ2X4uZ7LqQ3W12JDMO5t1spXBdSno1Q+Ugv1l
0vI4hI0lYsdrokrO7gjnmAq1bAzj4ZbioUhkcZAbdWJa5OLm+35osTzi64r60lEF
r9oKChtMNup5LgxNNMSOFGH299APS1uPi3kNNXHEYzFzJRflt6T1YP/CxKvfJaJz
SphmWuE7wezgX+VzY9qQd6yeJX+msS/qPDXXSUkWGbsCqPlxvJSB+FMbMRzhxnpg
/EOszwclcHbgYmbMoJ5tJjsKWpWx1iUeeZQf5aKC+bFVQAlAfcPr4OFetfON8Huz
Zl+npGFA8xSD7CKTSLGJmdkn558ZcbC+uHdI1BzdCODA0bUtSZwSppfb6i5Wt+QJ
4mmNLHVwUO+1/YhwGWW7ejkaKwihk3GbiMmCfG4QhWaAr2gGIPBXJm3ZL4gfVf/R
Vttzssir5VrCaue0ePDahW0wUOcNsJHF8bIJ+XDZiADETW85zQadawRBCKPEXRq8
L0klyBdsy0wQICUBrz07ibhB/omz+JkVGa4mtdwF/omzHZr+zf8gf6Fw9xMWmmUg
KpYlPscK+Aq2tywA0nKGg1FAkDwyx9N51M2QBa6LI4xRFobTo+Fp/P1lebbTetsz
R5qQW58rl6/WqCuCV+Ob91OLfe096e15KGZ6Jq89Gx2qjwXxTd9xxjTgDaCymlMg
6ADklQpzarW/TPod8+uGUD8creyFMB0qcChcqoOYVNIejDjS/txVauWGcW9fFekJ
nn6ts4HlDCGwSWvXfrPIWlS7wJkT7NtowXtV5TiWQrKXp49tEUHetH3FgID47b1o
vz8XCHRGxlXn4/sUohs2BEABUP49wTzo8lJgJZ8b6ciXG0WoqMUK4fnnBpG25RkD
qAkqnkVH8jGPwK/le4Whd0Cr1vNyWM7MUiYrLkVp5Dz5Ouz/sdU78EKHDQFZESar
jVIap43dvfnWEMAanI12afYD4Ue9DmZCZyP4plNjuQPGAru94cw6u25Z2WnGLm3F
enAfKGIP+uF9riijnSwdvef2ezr+WDPGvsqBNjz2ukeiSIBTm4TOGyVa3Zi2BKZv
a48NF735979TmKnnNmz7ObGseWrmfsLZu0J1SEb98QlIC3qyxShax9/dWh193uPb
1KlojCX87uHTOD+KWmC68Xv1LAGjRWQH6MFsoSTPY9yDYjvxn8RAmPL7C8E8NdTH
qsa5bs7v4WNoSoiprAizlO2ohQ3CNdDypufPHOL+fg90t5BPWm5VtOER5yytJ2aZ
ezDMosCVm7LunzSHNqGT0SR6t42wQ84qlaW/ev0fR/n32Vf7EkokxSrvS+InH6of
hGTnyd8DapPLWzteAOYvHC0Hx+WArcoJ417RZwtruw5wdV8WSIFigfDN6hTir3HB
mEWlj4qHTYPyNXE9Q3j3yMvWdPibTAkfgB2H8VrwG3x4EXQ9rEVGJZSNcZHG1Ccn
nXIKpZcgryW7zy8iPQWFKPrD6xR5vKy5vefX3F77I82VuiFkkekYFOqSl85mnsfI
zuXfmsEXDUEbL4Prt7tWxpjYksJcI03ZAHntE1fN+EAbYcr5Jy2lNaYlAYCNCpVm
xh3co0c2ugdm26cm+aoCa80w8JsnsmOrhDbOhsqUGMzVGybMYf67D7SElxvNb7P5
5P0858AAnenM7IJa/k8g7HvdBHhFhhlf7ZWWH2jiZwsYjDWqiTn9BWknje2LmKlE
d5USMis4FKfZ5HsSohMmnXRLUYvmiVETIJbY+kLJYcRb/J+FjHB746iuyTebPWcK
5XelqliaZFQ4lxbMBLMVGqaOqOiQ8js0ljoWE2MkAQ/DOyEybS9jqteXKZz4Lymr
kz+b3tvjAE97iPYnyzy+DDVuICcLTlYFib3mlqtnMd7urXX5ziX/qGhiUKAJb0eI
6UCA/7d0Qm3Go7NfkglV3urxvuI8EGxiQBO3m6+1KPLhJAH4u+zkaWUp7G7AD+O1
jHUv+HqtG2EySKJWbilIWdhXxA7exqg40cxrELVIkOed44aDpV8zi5CsqRzHzgk1
04S4W7k40Q1oRJey9LvFiNLCiSoKQB83MKUM66a5HJTSrcfothwLeaWpu8redxJE
H+nTy97eSnGQ6bPyRhYgyvN6wnntEYAgBVcSH0/eQvAGqpgnwF2MvOPWbJveMJQY
ToF3fz71+umjtgciUMlf6eBDD8OLLOwW71PTbGzk3TD/CyeON2KUs7enZnTO+tlx
RPZ72b6JdPN6/BMEkL2KvPBI0EwyqbPsiN9GP8djDeTldlKkeYLDskap6d2/a91A
f0A7wCo0WP6hFygqG+SyvGdbgxxT+AWnJncNYGmtQj4yAITsWQDwkj+tZMURDqfO
bGVpFa/SxPIxI1FEqY0C7d8RwO7RutTETgmhzM1IW48dFi32gG7h5c22vgyyw9ja
DI47Tcs31M68NwKzrd1dMGjfTK4ya61ffWCiShPQ58XU+VsqYjyzskfIOJ929K45
h0WliBk99dUhDoHW94E9jJ94n7inSUTWw1/Smyae9ngdbxoh+9s0NQDy1o/K/GCa
ScEvZJqU+vTKKciBS1mBNfKw3USzzWl3je/NnGJet9h2D/dAQfzlidMTGeXwib4s
p1HoVdoYNAgYU1GK1ehOpLT+Iu5Wshoq5mWMhDoQbX9rvYdEQAisNy2TWPfZT2eg
3+HWUkqa9aj+CnXYyWTe6CQsxU1NgA5bJfDQAkyWyYA0d5y/zn8B8q0vNh+tXkIt
XZEHWhVfHrxjVSTI9sElzuFNfwr8/G3bOYl9mk7vzOocgaFG03adBuHb/8tIN6eu
1UucG5N5fkAj1cW56vBajz5ziNJ0ntvNRTYpV0S0pZMDbgCHCVGYKaBknWMIp9I5
BR2KNptLGLwrNE9n9ULQb9AMd+99fRgcxMsKy3RBVLT2UdG+1fKWmusVkLcp4AYa
rrhfftop5TtcVtd2lVDWN49Pg5B/Sq3QKz3X2sNMzT5iLEwtfVn4cVfT/iMP+3+p
VBXD51MkqRzxeXHFSY1eY7NZZq6ozfGC+d7BUZOUdKiPakc8gE0mHLzM+WMmnxXl
p/gVqw09KiowhD3dn7lrbh1Vug60gFZB3hbj2pTavb3qstmR8DteCq9U6iBfvO+C
9BluYo4COY4+CSFZqUC3VBknqFS4vGXj/4XUnkMgPtWGzs2PqnR4vv7JpwUJCzBQ
NO0Yp0AK9zVmHgVgKMumv60KIruxbV0E3uKkK+UIbDJvVxE29UKO4fJAPNJpVphU
r/A0hhl+apOn3y9oVqERQodgML/dnIXzH0Ex8uty6yBRsW2wZ2KJ0oupXcEPqR4k
uk1q2oxl7W1W/xYXiGgdETy6CgSnH5h0k+14H0fbO7kuD5/7+3o0NOcOPrjBPPlS
mHKOt+exlW1TrJcAKYRJCXj0BCLBfxLmVaDjaCu2W5ckr2fFN2jhu5u6PipZ6BhW
G5SZvwTv7xcW9AXQ08Aw+hoQQAY/uPW0qO8INwpjdckidF9blhUYEZZGIsvVmV23
cXeHK0SPeNQzc5zzgxISy7Rye8n4cH759AFkD/NshwX5MhCkDCgmKggB9ZAPozK2
vhbxwRTnWZJ0+Yb3l4iJLnAabvhaI16/zKgxBcYd5ZzC2zlz+/VfK+cYTdbkFj53
VgtbsAddRUHJqhTRJTROXuRIcyAnrfneliebOHp17dY=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Ufhgq/WNQ8JXLsl/UsQDZ/DSM0/VlOqCmCYb9EHAi3xvV64ePfVa0PTuMxaMIvMV
wSjWNWEStWxwRjrjHgGTwJRUTwtCwhoO+3CSFsQLJvIhYNj30D+HnUItFjhOrZyc
IM48xYHTHTbmRIor65jr0Mf3j/PCu/Kvd26Cw2Ztm9CAVehEAcxvlMMcH+2RtFas
WX+7irdysfUkz7OtIgH9YL8aB3kdp5W4AdyhE1QXn4dkHKuyqJ31ZMNa0OOooTWp
PSpICk6eXOTNuk46GmvaPOpvYZP3vGo6UWvTPBcpY0z5XAnqRNsk5DSkSRBgjsBa
rldwi/INWtI8oojGBPb5fw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8016 )
`pragma protect data_block
0iEVq6XkX4IMkNGloW2i05LcZNWlSvi2Dbs3yfpHEirTISPCzgeT82KKlkp5s4tv
M+iBpRKnEgYt3OfBOcU9d1WVovgoByz0x0VnBX1wme7XYUxZb7uDcWPbCKF2uMec
NvkamB1uqQkgQ7M1alqQ67jwhRurRM4g4WFGaQMO0Z94ipaGIUmroyO37edFzYf8
NhvJH3KAYLSwIF9XI1NmQi8zcxzyHPI1VjUXt1HEFVpeuEWvGjJ+F3aYp2+JqS26
fffY4iW1LdsPnpIlZyRlQp+wVhk7OHqX0XhjZOXvxFH7VCtXGfAw+lRb2HJHLonh
4HtBIiZOiyLdc8LL/VtL4EqpJg2EUdrIYQ1Kv6Qtw2tI3/7tt1ymf2suqtQoZ+DW
g1PNL8z049W5Zkwgb6ugNBBtvKYZFPi6dBF5Qj8Ol/SiMxb+V0Y6kxCkyttHjdHp
N5HyUkwBDfeHfZmLqnjdiBHo7xu9IzwjB0ayqEf+1vx4LRr/cmPNYE0cWuaTdgz+
3ov6ylnHjcC7F7v0kboST9oRYam4ZP1xa0Dz7GxBQ97YCfF+0vitrhpIsIQdQSqR
3VWxq7x7D8RN8OWMJMqz2UaH/ay52KCxAJU+DGenr40ip33OkqeItLOsVhhzetm3
1IGqLSt71CRHFUxoH8wzzn6sbhmTIlKRrSAW15a+9XDZXc5BIOhCKs4A99FC1Wbn
zj3+aqNvdloxjFDnqpKvrgBN96+plXNwJjM3hyiEBRzIwQJj0WFuqNfBK2B3XSQW
cNnYqwsQIToytjX7gBZL6F3gUgbooOxdqU2KQJiO6gdnXfGxAH6wh4FvJxxqqDSZ
Q5U7yEcDiy8U/A1XFLCKKqU/qKSACCUbiqG24jE9qj6sYziS2PU9UDsHfge3kg+x
BiCWiKglf1Az8Yi/8LCavz432Fj+uT6MzlUzMFa1bcepreLNuAL7Cf6DZsy86AHm
7AknZSr4DTB5OsEVpPQFINQli6PjjrB0J5JRjXxSQb2gwy5/ZHeP6odo8VvXLu9N
WpKW5YmC9XvD3SxUAmT11JnCopu/Q3LnVQm8ZZuc3uocPP5HARx0pX1W+nyK7yup
Hcza9M6g04/Igt4peBUKRISeFDDK7u9YovAi7hBIA0z/qohgIwhhVaQJiKTmw5dd
4Sd0CUmYLy5cBmxOZpqJ/P4toc03FrH2A2dKFu7rLfIFdq+kkbHCdsD7/KFK7emN
QxF/KFE0JaIhGfti0AGBOmMt6qazouU7MDzNIUXOoj8TXYcDICov+VjC2VgUQXPI
whY5/X1Cv0ZyN6x44m1yKn38q1f7VcfSPwosr3MRAnztLqWEIHkZQAWcpM6TKPQ5
qJxR973NHHC9KboffcCDxJBHJofGM70wikWZxTyH/I7LyGUtpiRicwv91Ge96sGT
+0UzCPxxoZnR4lB6Uj5dZuk/K2rQZxY55z88NGVYuSU3eQnbjKdqPamtT26rnKCT
F5N6zLNiSQAzv4wPk6WFOFb3ttd0xj0mMeLUuhyXyeZ7sXdnbxcfBEa5tjKnUe5s
Xfr3KuX7GXBGZTM9YivUXIchkpxSBU1vDucfqTNi2Hqz/Bv/JBQrryVrSCGr2TCt
soSO/A3+/EUtEQCKHN0Fqdn71zbO8A6TXQhdKmSF9m/d/IwHq0YV4oD+hv1iBpkn
zVq7717u3U4vhgWY8QUf5/RJPplUhAhV5x7DHjja+wQufCJetvJSgvu6eSge1szJ
knISakLSKJGwaMp58MlFIO0EIKM6EMkZlLKx2pv0fcZdSSM2ZTAfPs+stbZghw2l
/7gxKG7HdZSQ2mPqEZzS752YDy589NdlLdGFGPSExTc94XO1RWqKyGrx8T5/CcRY
L1ys0rw9Br6kn9WdJxD8wYMlgAxqKzBgulRHIqrxtYJjKvxo2qYy7S3x4ZrJ2ZmL
B7p5ztxU44E5l2++0exZhYbBHG9ouDul5R8F44xREdvMLs/rDzzGQ03WWHTXb7kx
BJ5CQ8aMSQSfFff/xOb49xMSs6JiyFVDD1mol2NB4FGyyT9Iq1/8PQ0DKCd7Bpbk
+k8vM5ySrf41hb1fW1v/yexzDcrsO/n0/ktoNXDOduC3/++KrwDrtrX8q7FO3ILu
v2N3iZwNP0CzBZZtTggNHjCaTg+s6pCt9EDajxcpDeUKEjMGTaWwTu8Sc2gopNml
e0mTC7NEAlo3UHLKR0ismKjrLAaG4OfGEEpKUU0jSUlbqHLZ9Ee53Pf0A1U1op1Z
130en9VeKGy1HNlP2RFhgN/TdkxhnMg4mtcH1ig3TBS011vTnGb89RK+JnqZ267u
K+PoPPf7ou8fuFYA/2GcDlLDgrTJMVSE73uskhiWerbX/tV/B5fX5VdHHpXM3kjS
hICwVEGQjYL7FZZfrn7pUjqmI2MFjhDUTxDcXmjZe9f4nLVABGNd+mBRGQy944Rj
DZdXxdE+AHVYazJFWka/bAHrG51fVU6p3cMTPLfEkGkWrkZjfqb2uesR5nYGNWmS
K1XmPifLaPAm2L09G/ODsmrC87Wk5RPWkadDas+C1bUZdeuh9LPA9ILFg4whWE9h
who/s0F40t97HKMBXKIqoSJac24Zhbqz52nr7JqiYtpCJzu1fU0ZcK7Ng2uEroMm
1r0jpEV2TZZyzckrKdn9IyZk2wgk/EmORchVpTarwUmIXuGO4Le/U8jvY2j+jXFB
zGNtkEVaHq44peQnQ8DrApzr1lENOOlUFVD/3JPJesgybwm0Jox9RthATnMuDaiC
ABqwPJZVK2qwss+kq9Sww5yO1jvCDTOg8fxEL/fXvTOwhyEmmp0gaM81NLt31m1G
8KWJzwH1s72T/AZBqLUgabx4EYOS8vVIhhTsWznM2a93+WhhsbVQJYy4uegFPPxz
Wgw8VCezE/7BUjeW3DBqAYyhtx2xaC9YLLIoI9gHaBDWHGvCAqgaalbtRmWbklBH
3ulYAdRs5QSAllRZl8/axWRByp4Bd+roHl/vlLUbFHX4YYKGASA14ff9/S3HJKx+
EEA0Ec490mB4W36t3NQ5IVSZnvxP3iFCGVL5lAjA8rLmRFsXSksiVAsFkWp1nC4m
V+PrNpnC3Xu4u1ydUca2fBUN+R7CiCo/maOv1m0YmPYonWdpsfxC3wuLDjZ2p+qt
cVya2vx2VM5qUIjWDGvlzNho5xxCbu/HBjnRaoA3FFde19yr6YXlMUcPSvsY4NV5
WpEEc7HOkzlGn0JgZ+mXwqHUct680UVvsO6VtxnfJkz2PU5eHSBI9QhY/KzSMqBp
2uX85Wxw5aMhzkDsdk+3BTL/vFz/No82xTo3TGw6Y+pBZCeJ5BQSk6Rj+uWYpvLb
1OMRigQf8ai0hIOPdI33kMc07LJk4J83jLLHWRCDDUS3brI6Pv5SlHCW9IJmGmXp
bRLEwtdAxIRKhZ2sbxIZR+L6lTMRF9HtrNm3RNzV4t4bzYtvSGQdewz94CTzbHhh
RKPr9M+UIlWfoKJn3/+F0/3NgxjBIlWrr2SAtQjPMFNRyW1PsCQyeIM+WgeHxM3I
YGAgCw2O1SLcB0Jzxt1eca/eiOAmeksebRbu6qz131YEF4t4rQFqraLnE0uH/jlA
V7fsvE5c2MayItIHuZs2IYOUG0OuBXJx52a2lg/AIlCV1u/bGn6NvgZ2tx6fsbcW
i2PNK2iFo512wuPuohulqaYi3pFEXIUym1t++I1LnnWTnEx0uXjrFvWDpKmG1iLH
Cg7Eyq5TOB5amhMh0Brkjm3YWDhbkTwHxPWAPt8xTL+W+u9tsNXkoxK9AiRd9CNh
aUHoBuEt96AkMgdKKyPlh2Dhim9GDuV4U931stPam0FkCVE687NCQvBiPvsHo73a
MQ66NupQP8HI4hdtvc31l1PoJV3qMvFXZVJWCeqLmSBn2Z6DuhBB0IgLZSCbHrTq
h/1TUgpOKvFKQrnixmzworE0vRUQ9FSDxWfVYiL+BSFSxfdQK+Hqr2Kur8kUtk3G
veU5Um0aRbtoowD+1SnWWdBjBeojGuUiXubz8LrhzDJN37aUHLWAqoD6w4i5jVPM
/n3hxeoNDQR5FNSnikE5tkNFWsk4BOKtOYUUJbE8O/n2uXsrHbCsNTKzZj6PO+lx
jww49A6M5p+iZ5Z4iKK5jeyRIP68moni3eTN/XyhxI5b9rB4HoM+MXJwg6AwG3i/
cc1J5HUPu6ULGMAb0iHUA9ClsvG/BLBFKLyhyuuQjXXP0kMk3b3e+btE2eBgPH5A
igAYeYjtXwJQlEllnymrNG5BVzxBFSTM53YtFhlqJxSQZIi7mHoZI4+qnLzzhC7N
SIirZAcndqGKMAiziA5dkb8VEX1/kQTDggnR2Zswtfh7B4uHpxy6PV9Fx9CHDneR
qbN1b34wgg82tU88Elcw5CgRyxPdlipKe9fL4xMw3bSaIyu3m/dn7hORiRrNi5wx
iUF2R/1xcG9fC4O8vR0xY7atBP9HqFV1uxWSl03/FYn13jA4lfJf5MVccJ8sdYiO
UBFMzW+98meLFVLagFitM4qtXyrmFRktyJ9CBOexu8DeC+hO59yS00c6yNFMZ+b6
rP7oQMVmqgSMTKm7vLb+mgc1+nxKMt8B/5xzfbsWdljKcjTQdcfSAsXQo/FWGP5K
x0eNK83JYhzxgaaQK5XrcrMlxIYmruWJv+85Y/q7miIslnxVm80H8iVTtid2OkKa
qXQfUeYScbDP1x0kdMC3tJDeJjxvkZlMbz7yKCX9lmUxCwu7cDsCiU+fMOqZk4fm
+FKFBam8yC31e6bj43Xrbn3jY+Scd8JtRi8de/+ynf7V5trsFtupijzzly9KtUKj
40FFdrvvzx5Xl/OBZL8bJoUpUsZZ81Mujf815dhhHV/ZeaxkjABpgax6HVm81r1v
ymjKKMAMT9norEoM3RGvnrvXNL2+zv1CbPl/E7wUKwh2bB42j+UqO71ih4EcEcUt
txJK4U/pwsw0YSoiQVVqQW5DnPgi1IU4Fssa1815zbyOqFlDPkhCFyJxIWkpWmLb
vuYcjexn13eYuOzdKZEN5n5sUpgAtGXi631k/QDURjUjhrDFIg0ioooG06Li+V0s
RGOWkq5isbZ1ySXkAsfmyfI4cqAysu4AEZ2O/X7YqkEMV9dach6Ln4Oot+WN1Xdm
N+B8zovuqUYbIrSXvhnQKWGJln+5ckt0fmAw4k2BPoPPce9MxOUUROZ2pPvCuUlG
kFspuGbUevSmeGKuwwrt2JhpjCAax+/cNmiEyQ9+HJSY40i5SQFSKeaiBJE5DosC
vsuCfTBkvnGA8763rlxyKeeYh+GuICeod/avvqSLw5S0e4aEL3ENDVIgGWc0LIW+
nqNQ/TO3MvAr71Ws3KEjF/b4oG6nI1SwZMattveTyqq7POjuW9M2p2Unr8Ba38yb
l582FIMb8zLmyEFYWCGJTMtQyhVEcIxYpu3LP4YCaADxCF3rcsAS3jqMX/h3xS6K
9jvdpKr+XlwferoVpdnLE1C5ZzWqugDqfFmn/WbaI3PUh05BYiiXkiSZMZwQABg7
lGaD1hAlOFBhS5UgcstB2dPOv6N8rtTxZF1tyHS6gVH62ZvDewVln0c09cpeUz8E
+O3W0/SVLpzrDVRDTSsaH+kN0ZLU6NMMFpxHsE8lE8nO8UXVAgvhJ7pmtZwEtXbV
pPCdd95gryFHyIpoA/Ym9M2d4Csh1ZW1pKoqtvCpVKkl8s69MdUkpdbSz8Qsgwdl
dZ0tpF0KbJkeuxOJSqXUqVEN3Ib8lfkQxo19vcsBZcRkYrfQm9qca89AhXRPbsMi
/3EEzhkOOwb41zwAho7RX+XFu7cE99xpFvYrygJBHcEbxucEXSenjbJkqE7ZkVgp
NSWaK4gc37c/7yrckFti2Q9DkRQhY8nQF7SJcWOXwCXRh5EXYPUU1i2/EC0MJpbs
ryLQTX3CkX/4DhEXRsvxmRZUjMBzKKuJa9SlYitAO8rH6Hy63N21iqqu6ZxH8wtf
6ODTP0tZj81vnQzuXK1iSsvdqUJprBx4jF/UAyRv2hy3CWJdxciCuv9NrjmK3Fmy
AQqSmR8BZhc5WItU7YefEBuHPdcRfnriA89MuZpfjnVUF3dzfRGQ72Jla3xgKfXB
Z9G0ZKQGc9nm+FyUUJlKXVblc5wRc8ggzsh63SM+OgktK7MZq7bAuJ7ZM0zJlN1T
fp8P3ab70vI1+VlJrAArD6eAl5WJYE7mcK3o/7ZgfnCMPdWtlHnripAbRBVPrRoM
bq6+2egnciTM4OTHwGeb4W1+jSbRz5MwhvHFJhmdS9Rw2SNWBdfVVgz4mHDJBeZH
TyElpkw/LO6hEtwfQLaHVzbfouC6I6jjOQO9SExTG0eXbRLmwxg3+o8wTFh1OUNy
93tZdMczP69muKSumqXVmQPjqO1lq0OeEHnFpJmY1Q1Wp8fvq4cAwWDeyAmlD0XZ
Y8cKirQ+lSnoQ55CFEGPXbimsV27CoO1DeufaiE3q+3tGGEUsw+NKoiTjmc9urVZ
8kNpBeEtgLAG8dMGMQcnBtAplxshrH7SVHcoh+PC+i6LglyNH9gihGgbFkKQulJI
s3KrxoiuhlJquBSnZHda+8K8zwe1ekBAfFG30yb5nG2NFkt3Vpbpmr7lF8GJ1fza
n0mlDV3ke4JcMh3RME0Dn3h2lTGPSFH5mPINjf+PDVhv8wfVeaPPiF1gCeAiUecZ
Q0mapLWfcHlM5mDcc5kHfsuNLeCk0JtcS2O50yrtIB1+dg2PynQ+6LrM0MfVzKW1
kuP24euHeGR7j5praja9UsS4LKhSavwRSWPvbAk2/UI47yY4uYi8L36pYygOV+6t
JL1gV98SoPPg5CexWSP64iqkB0WtSbNFR8rdps4s1BQplOVddHccumEM8t0GQDWW
UuPZ1H3uxetMF0ANc9Wr+G4L3ZpFXlUQ58pAGHQQFv3aqJQBM0alyOOLPfuDIcWR
w/LRfqwtTBtcGwz9esyMbGh9IHEujZgULAHo1w+mHpPJxcizzXBc/z7xP+vpP+jg
zf1Qtybjtsf8pSciPo3c4Oay4rg0X8e594ESUj/Q8j6AZi5RbK4AkaCm9tOO8KPc
c57lRPriklJVqJNLC1sVfzgoDD4eYBE6zlmx16YNJkV9tSSerB8z4TZJNYUDIHUx
mKnUdjFmKaKhSXYByTJCLkvOcFb0iTeyGOlTZJ6juyCmUDEd0wQsP2TdDw++Imc1
Cz4umDCpyF6OqQ7UI1gx+A6IC0D0asimD/uv0qoLm2iMpGL+Rx5IJTgM7B+Pklcs
DyNQCIjvs/ibHs0hholqvJ9GC9HNoqD/CfdxgXfwPXzMWtGvCOLlaHtg0H0DhFAD
TXxRo8cT4kKAGWad70ttMCIOOaSHawnHJ540HCxw6drqY/J/fqSJ8upvxOPU1dhH
CA1EgySA3zV2N+tATAwDVKbjedThsevj/ZKUnQa79zD0qa6IVhgl2CKczh4LHknv
m5X3aTgTARJfpaNa2ALvjqz0RyICX6mPIjGy9oTW6vS0aUZ0oLVpKl57Azce10gU
TP/lkyQ4f15vRlvx3F9d2CYa18fhfs0LYPygJ4MaqB4o5O/tE59dyeaKWM0X7yQ4
URDl8ovQqYHURf/ECZJQJ8rAyt+JrtuIVlrYkEJcPmTUX2OGkIVVlUL0oQ5oE6wP
PryyMzeSJ+UUIYYP1gJLVu5RY7yZW31Y8fySc5TvBfYdhY+evTsia5qglOmjAxcK
XW9nWSxhLiVQwSLwDVwEWB+NHUHruQcnJ7rBE7o+H6SLV2WDRuKJ1W52L2w7Q75b
fLG/OJf5AQd4mPhp5+nUG59ftSLBcsHRUxB+l3J/kp3IBcAXq8dY38gEwSU8PSIh
VP4wkRNtg9+xUA9rl6HNMHiKVQ5VpnMZbJL5kka0pgHoBADODhmdlVJ9A1WGRkhk
Q62ZIIQrIQKgPF1kAXAzmnusPaDrLTtbk7j3yDLs0SFfmI1r2OvsAbtO6ynaDGB2
9oDWCvB6Vr0n20V/i5JNEDmrh6LYfRj0WE6DzBD7nhm8q/ZZNtHv+HarfYU6Fjb8
WOTAjrah7pzznIeCqOkjregihBoP3deT6+mNNHAiOiBGm9NM0wowaivUvapPz53M
yljeKLOMqDx0EFUF1VNbTbpd24rBjvXHycZHSI4Y18eBVfC2FmdQn1GvT11KgE5D
IgVqRii+Q8vsQCU2bG80nSn+IIMaIlQaScduvzClwBq1eqg/SFk0ghBOIT0u9Qj1
6Zr4p5EtiyGrSvQytC2zztYg4AqkJXYj6z9+sZKFcg9ZoB7/UvBz3IhKPFpP3I94
cPW0cj81xddfsi0Y1DojvH3kO12CRDS5IOc8tEArCaZPL8w0oeS3tKGlHUUSVkSv
m/I5GSt82OylrL7fJAO6/7Ebm0Oro14rHfNg32Y7B2dr/9qG0Z6a4tNrJUMcgtEK
KI6ZsOzr+hz1Mq32H+/G+GwSbgMsnnPgX1/F7Oh6UuG5R8TXjvvilI3sJHkSA1Tc
REog0DvWHpezz4ivktCHi9Yc49NiyiP/QMgoU8Q+cLKzhVJ4XlqBAhoVoe64kwG5
5+ULQ/vSAqUrZIWNmaFWyMX686PyR5T4pWPqU/9yR1IpdQsPFjRQIjix4JDIcrfQ
O6TUnSZg9Wf3QHJpk7ZBWrKRcmRfg/F9SFx901db5hrxeEcoa5I3mZLBYvwaanam
fROPgjx+ATXhRVbJbgK96R82aHiY91uGp3Doyb0zdaU5dBqMMwGe2r5tRMRGzjiq
T0xtpzuRxItGK+Iz2nByJDMLTKY1e+KRQ0pFxNc7cXbB0QxYIvSe7w0gnwXvHhWU
zmLZ2oGHKZNk6/amyzV+i7MIRSy/mJRqupvNnkwBw/fEZkak07UdGmoEDftDUrnn
0CCMo6bJRbLIDSF37AIBtrtgdzD76i7ZaQ04vRB55xXuVUsB2cxntkdIQJSQVsC+
33f+OrOVgZafK35jUrEKwJXbVtGzJhHsykqwfAA1aVjw6KtaWzRxqwYvAxYhwLok
CqJIEnJYoc/EKFEkjDCzjTZfSRwRkI2rZrI7+3yBkve/kOy26/apaMawm3T4fbmo
Lw0fpk1xG3k7e8FNT58bJtxEokHs1bzyPbfL9CDnwJkWv0wYnk1Ep423gHJFz0xj
sfFzlRSXl+YUnsB78E1Lot7CWtaWH3/Psk6D9CB5Hy4gVABdAWbex+mMD2vfp3Ic
0GHpksa0uB1Xfx0PzKVQjTHrqHibskPGYd4foRWW93XB+pUzvdUZDk8cKuYQpGRx
7s6MNlkal2p7nS65M9KMxJmCxHG8A03re+5Isu2RoIQB1L2t9xcv3P14Kzy8XfC7
vJby9Noys2B+hUDQGG9Ps+QI1k1slU5j/syqGP7hfSNOGnYOrr419n+HuOGoFMwR
59Gyu03WpY8GI+EOeaBN37U7PXS7dt8ChZMT8kbw2cT4gWlHEZgjaDEuAO+NtWN2
JIshdqdzTTxAeqaRIXBPLVQsWA3uJr2DDtnkCLxzCr2aUjRthRA5Bxrn7cgdmESh
UFvzRRYG1zpyUgtr7Jm5NiPhnkB9k+8IPRVzFmp2B84bIg/gUQxgPaSkBPypuyOX
hq3Mx5MBvj9doqBdGWwpkE06iLCSrqm7lJWYggX/Z9MRG/Rk1A16DkTsRTtnrw+C
ZzpwCJq+hfT2IJLl5VOfDIkpwowmsz1ETb2+MXth4zJao3fXJuur8y1ky25/njy4
aeRBCn+FSCg99iDRgegdOcxzK+m+og8pJX10fH2ZekghjIFOGpVekdtIPt8YoKpf
4jrh2Vrzj8GLYBRY05EIw5eQi/KW9MbG93KM9GDrK8jGn29LxZQoHcIOyKE+ZRQu
2kAjyjWE2NBQcOUfS+djyWUGtI0MfetZN0ntvRs7o1+aU+YDYSQ7Qayd4AKrexcn
VPutONpcQbS50hgd/49VEJIVxg5jan5TJwwWANtB3P2OJ+KLH1G22Wh8O0wSiStZ
RLDL8pXXWxTeEfx/InRz3XViGh36KWKYxYfqxpAnUVx566Y+LQ6T0TuaBWbPGmuK
JhEJH3q4pFtG4G8Y0YkaiBqPoKEcHcprZgQRrAc0kt5lMvNDG+fSSu6CiqP/ilyZ
MMJeTu5BkzzT8bcWMBgm3Aoqz1DcZ0vc1VHQtuMwALrZmu6dBNWifCkR2jZQKGPZ
EGxZUA8YaKObSEOAL18TWgAa3KsPRyHKOfkyqhfzFo33s1H5KlQlsOiaAffWOKLp
1ulzDN/aBaVg34fDV3vUPcAMmSMDfL2lgsVTQ04rGdf4CAsLPNbzvWDpQ3JY6QsU
a2OxgtNaLqyEZhN8LA30VtDcIZGKkHcyNt8PQGwAb+pvvnbdl3BPtqkHsdK8amEJ
lCUnabGY/Vs8OB2vJ6nIqYhCkoIc/1xWYxzFAbxXsrcDPXD/85Tzki2F0z38I9yb
pGx2codglb9R2LYOJVmoG1KE1aqRkplLNndrWPSYllc3W8SND6sfuQRtjXyQOhMv
FT1t53PZe1DycQPyUfLzLruJn/GUIVOATDk1vD7ur6ffHeUqZpkjpryC3mLTR6Vm
fVDy52TksAaOINGWXGNjUMxnFKM5vOJzWhC3tMrjgR3XUvKPjxsErF6oDUXi0Uqh
90NeC7umsJIBeQ2PNz5DZp5sMHJMgTRb6sn+z7/3l7x2XEUtVGcP2QltQfcbxZKu
Zbn02g4iewbQNF7mEF3sjL0RwaIH/4QwVxf9MT3u0A5xRHHxRusp2yDKlheeaTwR
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UtswwrPjr2VNxYKqrUnnwpue0fVsBSXRd7f4TkgmcgFiNljUOOL+clD1J2ecUqZ4
JDvDXUx+wCgAqOMu8kio4VeALqQv9haHBrYJ5qLTLn+yPLNmNGZtj07FQiQrf6An
rB3doW5GRLD/uYNEgTnJW7oQNJ0mKtxZOTZF3ybmH2hj9rnSKRQ5s3Ic595EjCCl
ifdegJARE25aU+q3lLs1l0aSeUcOxAwwnIdR4WNjijHwNtZyxdsIHju3CLWKmCOd
XoqSDz/j1eWxPJNRkmHB+3lFx/8VHugsvswCtjoZwyt4oVYhhPpcteKQ8OxKub6N
iVpaK60Pgd5YEOKCthEsBA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5392 )
`pragma protect data_block
aokaQn6Z1t7oBEVzO+ORowZ1qrv3oOeGXfpNSkFsXerqHP97igz39jpbN9Xae8EL
iZ/FqJXXRAA2NMDovrzZ8ki/ZFE1+J5KmJGwAaSH7XWnOOQAjm/OpRzK2tcnNRib
oy8hJmcHAQjsYBhk1qIPLLyE68wlN6X3voGlm6cY2coMrQNXuJrMwvr52f9pNBaa
1autLnmSeEGknXWkfyew2D3VKYTz3xXe/gjXvRb9LaAkD7jjSjm6J9cXIPeY0PtR
sOhbj3tw18ZjsQwrQnCLENQOhFeZM3SLE8jbcFW693YJxVSGNXPqH+eJIzOX4w/t
G4CJZpHUMuPuO/9BTJRcCTkUHVF8UPQEZKaka/gqtt5rowGmV/92TmyreHNNhxh2
rqsmEGii8m1n40JIL1a65Ex2T8jWDXrh6QFwXYNKpKQnV8hRTUY4mRHxvllwm3Zs
jrsR6VTaSW62t7D+lHwZ8awnTVEEV9KkuevCE3Q3pWdPjxmT4p/HkFKAvPp+mBht
Ze4KB/Zv4jv1SgSBIgsmtRZWFRarRQlx/dBOT6axRpMZPI3N9gAFSySrlkKfLUQi
PEafvi9KcXIN6npcFb8OrMxV/U/8T1eldrg4LmPs7I5LyH0U2zAQGBsmblLN4D5A
K8d8moid5u6PDxODsPZdw1phxKU+yenqf45MyTylhu/xPHg4EuVQbd69Cx0dnfUR
R7WGzaq0lUJSbJ1KQD/NtJbZJ+u2QzDZoJieLTyA2TvQ1EVUucPOXHjKZ611V6eT
FLDgAzAKwZktMIxmLJcmrRF+xZVgR5mpTT+2DCK1XmzFkt7hQppuVN5WCRmWHhE2
zleUAqPD1yrR2uHCBu9BKg1wvx3NKLi+SADLbMYfSGPlzfY0ByHXRgCnCGHgAfAL
LnqscUDUx/gyNIUX7V1cdlVvuiJKAZytP5i5mFBMHS2/Qzk8uyjWZNhOvomviWvq
7BDr3L1EvuyCrqk0tecAcn0x8RhFrgnvqJ/cZ9XRV1xR0wTuaPjafbLdJ9wxKpZa
iTDvUttpCBOLMmvuxxTxqbZqMo0Kqm9tBxTNvQ1Q0Jh5bhGiyZV2Mk2wcK3qF5GP
J0AzVchsuwhFf94M/PoGtB1hSp7SRyaU4kOWF7CJf+iY95utLuX/q8ptVGcj7Iel
2v+w3vB+hr2/KUXwKu4HNS58cA4/44oH3WRtIFZMkBBudyKuY0O1lX96EwnVCXTH
xbP7HyTR+0sGIXgq8fxjdyRir8MO+TsqZYiwPaEJ5C17KR0i74h6ijC7chfj33Em
p00pHFr42LZ7cWs/wjHexUcIXvMjcKjzWrt2P+X2iNr/XxmaeuCDp3Gxr05TIYZU
0G9L/nv9T+FJ2I+TzbsCwKD2YXqm+QTR0z7kFxszW23QSSmoyg7RdaO8gAVF5JL5
M4GbRigXyzyP5UjQRSiMTmXRjkxTeJb3Lh8LZkueimD78mKlYpJAJiN0sqbkioad
bjewllBUfXKGHaeD2viyZG/MOLP34U6uYw3bGokPSTkyPsxubcn5tcGiJ1Kvfc3K
r0xOcvjLCfb9TxxDmeUOTqN9OIyCZUqb8qRuLmC03TCIH/1zLO9uSue1Lmc+p0yi
hu98XB2pwdYcEZVFjloP9Y4nOJExdKCiB2cNfabLgOtAtKODouHahmoPnEh6jtFo
uyq2KFTraXj+ig/FJMVV9TsOGeQzGdHoaWKLm3FJhh6pLqahPom0Cq2ZYBkPk/+t
X4+1nTlvZoV2fmE0AIZgziv5uvah9YoTVYzdAh9a3KEgQAgamSfAUxDAxlenWZ3K
vYNchYB5LwjxRqGhJa8mOuaUgfO63uS4JaAVc/Sb8xg49D+UFv36pVXRj3YoauZc
R/QEw8atoKVc0xXHHNNAE+hN+uoW3gB9MDAp3lbA5uY+vQoO+5vA9dyLkuxnBT9K
2+AjJ1OIMldir7uf2Sy7YtSkMMrGCGhnq+QgnP7YkDwLCunMqxEbhIEhAInhtQei
dbjxt+masB56BCSxZ097qXbjFmYwP2iFua2CZnpulWEoPq4KMn59XFP+ghqj8DoT
LYic5gkQEh0fDwOOFBh7TYxU9n07FPSstXQtoNHbqzf+9N/oSWrlqS1WHDXX2dNa
6PHbhq/pZ9W6VjDutOjz55e0ujb+DZUrARcJ9sRVKvAqha5dDssyWJpIiefhXFRw
xY+HtdXATEnZu7u63uNXPjUbhL+2pr0Wb703yRFOKaiAfzgxcpUUbLhHTce4LdAJ
560boN9M8/PknClGtHvR/G35r9QHDT7dFWTyBEImRoft0Omgipazg97LmcCEceQt
QMAqDlXX3qeJeS41GGOa6xKTa9m/IRe4sQtRp+u/nbIdgOLbmrA/fS49NFEG25Vx
FDhA1KizAcdP0v/inkvrLPvzy/XtJ0MppMEY9/HEtKe3kqiCA6T/1Ge8IkQQO1Pp
oKbDYyH96oqE/310aIxK8O2Ky19ihfqKlA/IUwJzFCetFARgvH8SvhAU/Mpz9PDu
c2b8VB2jCJ+MgzWG9vUznoZf7ONmfMOxQAr7grNZpnHMPPRc+bhZ2P0dR2yhDc0g
Q8YuZiRANs6WEFDocDmZCzTycR4EC6N73moGLcO55VgY/UjdQoW0FmHB2kCyYvHU
7593gme0sAfFc0vYEr/GiSwvjgmkXUFrEdInXwKIocPpWe2oMIQF6K+yRCC1TnVS
vIRuPccP+dJuD0xYRwQLOrb49HwDqdCNIx+VsKaOyUfw9DPZAMIi2kIDHSPa+H3F
GZ7jEYVK2GHvxkhoIQlAhAYDLSbA/RgpajE100XhdMjoCNQdIFb9eJ241DS68nyw
zpeKtW9Xy3tDNdqOVzv/wuE3k6hFRFgF8ND/rL6IGM/Gp82Q68As4CmhD23ZN+Y8
m0P+fCyrmc1F2Ar0wlG0vbSyqIfHAy0koc5VTUZT/vt1BGkc/MjPckIDAqtmW5ua
HUpeAgN79YhBquzYH0oelOZf/fxkcUO7bHlAdHdoGe65i8VYeaITMDpfHLV2lbzc
tS2DkNW2aZ88FtzS3PIPvjA4yefBxsdz/ENmyH5VaFaqL3oV/zSAw/Ogg8cP0UeA
ZjVqyMrP7pF9buNG3f1m7PDAt0ewZjyrVSHL+MuPFw6Ws5kQ9LrjZFurtdNVOPzW
K/jvf46LbHTQbCYVpYybjBZILOVrg46ljOnqc17KJoce8XdrEbPL/lBg+8/RZUwX
ZaTMhqjwrAyiQlffLALIjQ6EFiW3FZrn0Fe9eB5y2wei3XO6iCckAUmQGbZ8iY0C
VrIIIATMVdcH5JndLsbgTgTPLE3P9Ezrx9PmXRnNjW39HpoghkKEx70seaZlzzKL
lp6QOsWtaQDtONAuBRDuQlXBKTw/c8uS5/JkQe0BW3HSBTSi2R3YwUNv92CePTro
ASuJNKvZiaUUP6FxKvwgTVFxBF4M2Co5cmCMNsYczQrnfgN14TtlkUX5hb3h+v3m
ka/Vldaimf0fhYfZUk3adCSgNEU+9ETz5FAMdYE2/bxXfBvJmlkLPl0/70h8VAi1
WgV14MslGZprUbZEE1NPB7McFDgLyxd/gkSnwjbVL6uGFoX/oytE1li2gAg9fjtG
GBiMdrIIZys6mu1DiCrOky7TzA2SRseK/FOg6zWtmGMc0N0d7UG7xI0Ht7xf1Vdd
hDjrY724JlpJG5keqOt9VTngb3XYyVrlAdDKREYFmWfHAz2XqlNArAK8j+ere+Zn
RIDfWNDEwKMRgNW65eIw1dVScwCEC5NVGPqEV7c4XU5fYIZ6GXrfti2TmhP7YkY4
g3dNOmfHcWyoIxJo1Ug1Ipdm71NmmAneyTNeqTglxVEhpH0QlParbSEWpUvpJH9I
wbfr9uQyEVoQa/aAhmFpbRUbNrvYkJ6XpiOPfzNMQxEi1rfrpC/7M0BN/Umh0cp4
cMND/xL2wXsjbo77n4SBMaDC0YWJ+RKh3aN6JMYA9CrLmqamnb7KeEf3BZTDfMt/
EHNpPmCZ1+VeP6FdnQ8P0JcGQP522tdcdPOCWFPgrbrp+6kFsJU6YT/Odv0fXY2W
aLZ5Wf6/y1EPN3tz/0Fn4XnyZ+cVD8ovnuIKgrzHpqiJ6IJJDtCYC7FpAQAzOgog
B0JPkpBOCFaoxcVGLAUokjood4ZIzNShWrfdGSTqmSv5I2b+bRamcGB8J158gGTd
Dz8jIeWJBsiKape04RltHQUtesclRT9buFNSw7Kyv4VAjb9FJEZGTwoOwtpS2RLA
fuk2G7TEiowr4KlWDBwEZQy+zGC3bk0t+i0a/Gn+KKyG2O7tN9+2sfKIdOUBjVzp
13Po7gtrk9MlqQ8QOcJsi33m9O+qkQD00WOAoUjnQs32vXtJiqohjxtOf3o/vcZd
ETmrMibM1p0hy7fPo/A4WN2n0i4hjpBo4gE5I33cwoqtlwUWnb4MHSADczmfrn2z
OrWw/763VGSpEJXzpJ7FiIbNrDyQqDMlSSYTYwhec79ZZpvEPKVGTtHTXHIEjXM/
q6dNpzAheKq0RZXrkcQfxzhyqxEamYzAVVN8Id+rioTSlter0sK3imq9J0sJaHFk
BULjqAtYzvO9dSJxl6bPOLlwMoiu5XSIGA1wvedMyTYbrqN6gG59AsVt1JrIROZf
aoGipbuTceMDIvbDFrQq8hFKw25G9bEIX9KAiInCzhoqR7miIx5KCgpInQRkebkj
DpKOXrdbnHpLR4df0cfcZI4t0rdOhUDrH7YMVuVXvyuzCwQtV5fGeW4ZgbaXaRXP
S1lNeqInBiKqLw7l8JSEEUTve3vldcIeKT3bAnhBAo8kb31QulA6JvqEJ3i9Inln
9JK/pF3wQ+Dd9fp/xn++lsV5v9Cg4B4+qqzjZBtl3yxXFgZ8N3EWrhiMPbx8UFz7
AvFuqoy/BEEY9rerXygWFKh8UmQWsVXmY+DZFdKYPCXQGJto5tUdtUDfDa5LZhZk
4NMr9dCwcjD0qWRiwLIRTIC8KkILZbPsGEREuAE5CxfQA+yH/ECi+zR853a/8ypI
N4aArkwiKfHax/J3vwpOovNn9AHJy4gsVeVqWX6cnkHPa0wCDFGRc+M7GFBJYa92
gWONGGNPwUxJpXII4g6N5BFVnF/v9D/HpvVKu9pSDNNJJ+DzetTzq0aoo131UNx6
kAIWsI63h3SLYul+mhZberkltk/MIS1aQqiWeunIxlqUMnTz6kYiYPgox0AeEUnq
Xep32VEefKH2hmD3ZxMPTyLZcLyx7gHz8vmfz4CTRxB4+/2Yx138rdh35ytOCRfg
KEgjBDKdIkFHThNVF4OEhiDWAlw9czHd5NNo5UNQz3iXoajlsj5LKk41r80xSB/P
JnA/JKJ/NvZKVfjieWLfa1mmFGYaaUQFaJ14y4xi4iWuREo0CfhVEay9iEeKoqQQ
UZJzLbKjLrmmAYWwHkewNqu+ZUsujoW+T1FozijF6/gCgShSrg3G6yGmMVbRpZ+o
DLsRXsKUlF92+m5uCWcq0SoUBSctXWrItplzlaxzXH7Fry0iJbezanJOxoD30NcH
vX8Nkvmp1mIBh+b9NBfLl+aZVPMx2Tf2WTsj/KNGvBdzCjlmiUG91KjLIWAcXPSU
nONyfs3UBSzkNP9lorcIKwwVLdA/A5SeOZIFUVi6aOL8Ou803lLpq+78k83N3a7M
cuOCy41pMO1rwbn/+JopXaBklaNPSWnrBLkoIM1DO0/3HgpLhTGnqU/ZY5Gjj5x6
4VmsosZrhVBktGqc2+dZK2WYRYIxa73nalrIV+RoHIZsDw6N/jApZmUoPqAllqiW
P61bu0FLTmRC1V7BcY3G2aiycB8a550kLwpsXEooWq9dZeCtKHk756h+0PsDQUBE
60mkIx+Uf85FD4c5TxQmEZH6fDBgUQzKU5Z8FwLnbY2rFCxvGtnEUZSK4tg4OTEX
Xe6/Zmbb/k6uy1TOSwgipI3ieUy3CtT13PJQLlTdg3cl1m815ob6Qx+HGGKkPQ94
nO9BDE6WzI/bK69mINOZMHwSoGMfZdpztDPS9a1o8TdcwkfOWfxk6QGzS3mS7OHi
9Xw5orRrvoBTakxY0/uzhKFgQRV4KTzhd42x6ei1EHbG9uFI5QOeGDMPjmmUaSO/
EnBc+bmwyDmJJl6Tukr++l0qDXT5VFuT7xOdxowGNoY5OsZDvpteuMVE99HxZwxF
imsmM/D+HS8CFpRcwaXD2mSgjDEHvxemOr1u7/2x2OCyUPG5G8XjC+BZEZIFwPFi
OEK8wLUOijwVBVtyZHeXcTSDVKifQ3/iTFUP3oRxucdYdxUYY9Xp/lrEdBfNVobX
HrwsYOBTdMYVWQ7jJdhPtHlnKJyB2vUVWQS+FhEF4zoZMT57XdCAsO/DFZqYoj5A
yYUC2J1X+AwtXRKS8j9Eva2zCBnJmTXbwwVBtwrYbJizJl7j/W/ALBqPhw6dYqQ3
ljItA1w0oq3+g93FXAEXwwGBkJp/z0oZwn7eynl+r3Jd9PFVYwphwEhqx39DqqYJ
VIw0ImPC9XRoKZ+FzuVEVOA4aZEvQsMBmGqvQcN21VaJ/OAoG0xWse3USTOyNPAZ
AOkF5WgBMtGiyO0IazHlm5yph7Kl3g5889W4mrueYUoWXDjy1fjI2shCypK61bqw
aT2HJX/XjAIRRb/ap/hMYL7753vb+sLPHIQZSuvKlj6DWWtUMuqMwKoSs/NZo1ej
qrH4D0e1gpLDSVkhd6vK1RD6eaOYJUJ8Ng058q0OTndF85k4zRNGiG1QX/of8xRn
LX72w4WMSa3Kcskz0lmv2sMfmqbXQlr8n+L/GQWSnc6nlHoctCrsJAPBjY2nXOa4
earGU3EhVp8Oa00YIvpUyzjicdvY14IL6BVP1M8ZBkMzTlMQfRXLzK/uMjUbTvye
C4y1wGqTQZjoIkBJiY/KyDjx1N5EKzK0dGzCcuNiQo4tC0LdjesySq05FrwljUu1
N03k22j8kdFkmjL01Pl1ehpiD12lkCloPPebTb1UvYTVORLEIfw6XE80gw0PLwWK
oseL7vFk9npzh28FeGXJToLh629bnMJWMexPumX48K1f9FTcXbGcX/jPIAhVbLIN
Vy7BrtAHtqIi8EFxhG7kAE/ruh9om1LqRDXwT7oFjpUkTiIB5pi187WlNU0Dzcgn
Uev72C6VJQv5iN9FGP+/vPXTL/Y39Bi9aRi/qNv7Yri/3z4CHfbRbUmm9xI+tTyz
v3aN4aKsQIiSdhPfqoWGkw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nDBulu8u4Fhu/MpyA5sWIO86Eua2Oy22/F1Zi0P3kBqASaYZAQB18t2VfvL/nlnx
Tv+QH4rXlacuyvr9gG4pTlp+vVROlLlak4mqV3e007kf4gSDU9CoZ8Uj9uGcLymO
TS/33KgC+Xs6z68j17Kdyk1ENbCcijYNxjYZAdQz4KYFERkeNYNjc/WBuvxCEbjO
M5gE2bX8om/CL/G+Zio12261N5O0H+WaREqGeV8njOEt0E0wyX2TAnndaE5NM8p3
/m4Bh5STVin1rYyzyVDSuEKno4na+Yg5IRvgfQPoF910Z21w9N9zrgNIkdjMiBkr
OU+Dc6Frd5kpZZ0JELzM5A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8864 )
`pragma protect data_block
UAt9v5KqwNbu+7RGAzbzx1GxiOpon20ZNyV1EQTArfBdjxfI0Q1WJRGQ2hnw+/Ud
NHlDUKW4QhtG65sX9s4NIyzr5KW5ft9YpSUOI5kICjd40klIpCkgexXKBq5L/VNH
IYOIs/WrSxAFrPkPvmkLToR1znPL1PS8m25AjumYxBoB5D8Cw+5EKldD6i2fhHpS
h/IyK2WDyx0fh85A4e+WWwifHhtMoiFSHqKLED6AEEZudjoSkAI/yprcn3dIt9ov
LrvIvocyKpjVdVQYwbMAnvKdm/kAdrLRZN/KB7ILwzWgiAYb/NnIWvRh9X/atXAK
jlCBYYevC+YGu1XHos9Ho6JMskZjhNRZsmV1mzia5vqCXGoP68nPdCulJQ3hPTfD
PF6BFry6+17QAfDGhWHzts7jwGOi6ReIbFafw80n218M+aQS+Dknxsdqeg0NBR2O
ZHs34gMM1qjRd0SD788Iu0ER7AhZVjVYy6zhdM37mlVYP6yxJySf6Ltpw1Jc4vAg
R8Ssqc169lK60ZwoD2K4XvBS8PN3/Q2LnEi0nkSs+vZaVfi6uknec6c9xsOMqhzF
4aoD2pAb3GxZjNSFIXLmmOkhJ+bmesOYc7MPealNeccZr6MHZj1o0y+7q/QCOJhl
J4VXGVnuHJXuS93gvQABCJTWKjru8dlXspkFIalDTY5vfttskWRHjW4C098dCBto
TPFHcJcqVcbaRAwdJDY+I2Xzol1GyqZYuJJSYXuUGeXf2ze2tC9sW1BXepQEo0xE
J3GUTwyr+s4ioWwlErh1eVjM1qyOJWeqQnZ1ttz+1LuHfI3ExCmp9bNqCLq5vvTf
UeeXGMdnpTvdaAt7WZ8RW/LzSxns8h0JvQMeAFDWWoc1+DM5ygXblMWpiC6amm9A
Wwz37cqQb4U6W8vQXlCHiCpwltQJpCoZBYmxd2i5rPMnsDXZ5PHJqVbVllKVpa7S
cB57ud3Qb1Yz0kc/2y7KbQyql6yqv2UHgYYqy/froS2UtQeYp3ytHNwu781rCy7X
cI1+DymkrgOx50FKv7t4DA378y6owgdRnmISzzPJ2/VKQ0mHKd1cjOpncrjd4Y/6
VqPqklzHv+oDHwTjCv3SUyAIqV3rHgthWURa6a+n6gw4Zmrwfmos1O+C+NEeZs2Z
nBfdUHTbnCUITsD0w0NM1haY8UO7wCHHusgcfHySX1/GeKpIvZSVOaffif7W4thG
elMQQwJMibFwSaweP+nkBpqXxa/Xd8sJUdqYkbvMxg6HTTPo7RK63WVOCWdpvdTI
ylSXrkJwLq+oqb8EzMiCve7t+h3BGwkLlq92KFIQ4xeqVIFTPS+u0Zz38jgJ//mC
Sg7dalM0GdHX9FzTq+ODnFtV5qKYhV2ub5JdCpuVPhRUH1cf4okj7CyPtxjxKK0q
N8bC0sFr00BiEWsoQ6qDsh2cV8k3c8qFvkLK5rDfJhKZiOHnUITtSHhJpfuagqc/
VQ9oAGnFMXE3vJIY3B6DQoTCDP2I1vd6ul4CWkYaNMxy7d4AzJnk84veBMNTUhyj
HUbf3ZWjbhLwI2G50vkTHf0rsXSjoEIqxbUqwNS9LZdg3mMW/A+A5MGshK9c2NkV
FB3vgemdtEAfNZzc3JI3j2a89rQeXU8Z4kPaT8XXddDTfzyGAyrbBCdAGDWCx2e+
mgUF5OB5vBuKXUT2rlN82SXDc8fE5J3r7qbISqe0WQ0DdPTVogCWPQoRYq01POYO
xRLKza17stV8WnoQZNsxNxrDm8UjNC6ffww00JOAvfYkGyeptnkgO4j2xu7AloxM
4j1PR8gi1NtDJcQ8EvJ8253qGbj7CS3ksnIXOCCd/CGvhdwCshLmnAuNmoQDIbAa
QsBn5nKsaQENibUxzlvcw0Y90Ivq6kmRVVoLDfiSp4i4BoyYbwpCDfAoCLQ53+Fj
5V3xj1GKbkE/u+OSQ74zIEgez9rLLwxVn+Mirj5ED033lUX/HwwXqp1rYjsbdHAc
O/04Es/5QmTsjW6FEWsBHAg8KwawX3wf44x6jNoIjwnac5siokb8bJIrnXBY8yNG
UI5E6PG0HXoNSrkUKTNJQBIu4c90TJ8pQIfOhkQmgaUyfshWBJ0sqLxKGJIUVC7s
zkAm0DuEmxVkT2RYd6r1s3zSxpBjgglt7o9weiUZGeAzeymyeX0AtO1ulRHzX07A
l7gM09ZXBMLjTaBa+hQxHHjTAJc4c+kAtVsSM3YGdnNOgK8+3+QQJAiu+UJX46vj
joGr8Jf2CLx3Xx6uYKAoUcwLznu2FQmyTsRsu+oXDjtTqUTVRnKGqfU3fNj/Chjw
8eVetl84kBFnftLHJUmadLo79GgLgNXSJAFkzz+iCTpDZhu5j1g6spaWL54jMQQT
LD6dE4+0WmXjGQ2n6/IiM4X8bSqhM/metz44A1Zbxz5zwqYQuoNS06/vqNlNj6Df
b2BvQBuZZJj+RtdVi171q5cWO0EjzDCOaq9+wAaGDFNp/LDwoXWfxjpTz+8aYcbX
W27ayf8Z1lkahjxZKXwxUMFC+Y3A8d7pllqlMZuo9p3UTR4ZnY5BqJeTsU/acIqa
Ya5Fz+1p98j1RSVsGRrtZ4qNKZUrxDNA2hYq0tfmQYNKmrMPgPSfSdvTKwD62hAP
Z4sLDQ9Uu97No58UtMIZCK/Oo15U6wsY+inzqwLfE2sUyh67vsdIA1sfg6mHM6D/
MKU3xCMTJQUj3H+qZGC0BNb9UAWhYqa98dAQxmGJ6Olg4GMojTjqRhut+qvd2MLq
q+xQjjfYOGPFRQ90rZyO1g1MGBOZ0vKo8qqmKb2AyzEI0KeqmlNOeyIm9I9X7GuE
PvuFfyOa4e3fNVfVbEk/AnuQfMnHgf5kKULXzsFFLm5354q9tISBui9KFO3okVCs
GbfqoGFzqPPEyXpCt+978YP7lnZ1Uq1NlV8u8HCpfVb4Gt8kvKD8/plUOnY6NgAz
imSez+qcm9kU5rt0+PzcxZDQxU8s/pv/dn8mg5sTIsfZha9sQ9VA63SPOLn5yIfB
JJXah8KCRQIIlMd9YfgD7CZzmfl4DL6rimQJisi7d3F6nkuyd4TMb98BMA7wqwk5
mFD8+BxQ+fcqbLXFwJoiu582gQJu7/9tXrBW49f8Rdh4ghmq00rjP/aLOeL+4ipl
G5vi3oXscIj5xp9sf3S24auERp8Gnpft3jh/NJcXRP17doGzLkXzae1IRQ/0NQ4S
NNSZxXz/R7b63jGCPtu0bP2kHXMJ4Pj74JKpzdCDvJFVp4bODrns4p0l4Lvu8rJu
nZ1Qo62iGZwF59Z56RKf+4LbbEmPyzWU7woBycLgwH+Q1ljeqZL3C+6mS1H2+MLB
B2A69fvM38jgyF3Pud5uvb0thmM7xJxcZ4/jX8Uc+OqIPsdwvsoFa0v/0CmJQqXC
/gC4dnHOIN2BLAzkJdTEmUuSHC/XtCMHqzHTwXSj6Pw8wbhAcBfA1zMtb4eBpX4g
GSJYA7SHA8qnhOA+DfN3mCyZv3GbfRKtWFBhZWMCFt1LQqrgQdwtNl5CdyE419Bw
RaZ7MwH5KAHnj7y6eU4d8INgKucSyv29CtYPErgQJf80gfYunnbD9aNZ6bPdxoVa
fdU7e8vfXjXznXgUq9nNreBWHPEVtiryviYeUoLI5wQiyPp6M6XNoQroWXXCIvJp
fYKDDcbYQI25yDSi2GuW6U1cNl8OziIZiZHW0VEiR1nu4jXGCqO2rk+ouEI7GD/6
oNhBBnFqW4qmliWK8xU9/MpLVr84yLzqmcQmjtNPHjPG9QCkIlWXEcyJ/VBGsvcO
SSvrw1Sg9gQ8ZJZF43dw7l4PdInmLPGWOS1VKez8BbF9ZMHa2aKykx+lV3zO8gbF
T5Yu2NWq6R66vrSwEGwHAjRkZnlJv/+ldYGTlBZwmqGHOz+GXhETVBFcgal7y5s+
O8scToSdQOhaaJgWQYEVLUsBv3UQz6daOMi0a+VKEM6tKQhzG9Q42C9ZnZLf+ilv
DDql9vG09k0hqjgLnsO1oJzuC0afwLhdQzFGnhvQRo0KUdbnaNkgY9BLY9jEf7QZ
tPsm+uvsRznz/FDTFJvGbeLB6oHO+242n50y+mD6o1NQnwNW00jRKhikP/0lyMcA
S8KYFF1jJlCGAALqzdsHtXTiy2gDHAz7Xw6e/6NtUeErWhU1fnyK+uazBRPy/cji
9OQPpRF757XuGn7OeoAtIaW04DetFA7tjVkqtaxqwcAeZ0Lzj2qbY7OvUA59mdkd
ZhvkOiz6GJmZnriQ4Qacb+p7s6Yho7WjHzKkHFaD5DB/Y3GmtKQisA7zxvHq0OTN
tBaXEXOKDWkJUyW2KSx/Klpvlo3OSbnn5pnrtiGVRyGsu0f66GrSPwgsEzHLTvqz
tkn8S4+a1UG1YjAw3rO+1P+9j5FOrrSEc36vVX0ss4GxuWTXPMfAGGqN0c6XKjTh
Egbb3NPxXlEvOtGFiAWHvvw5NAY2F9PNqySqyOcKpwyJzNeYwULpwntsw2YJcdoO
RD9KLtgN1roA+E0voDS9mNPDwppivNKbA3dvY/G+jZMDtEkzA+IAL2e8AhJOwkWM
yn13znBktN4cezO+yVhX7bpZTCLArGgTRHuSFk9qjHDlSshQYsTTvq7ctotRKLvY
nFyr7mmk+QfIQXeV9eovCzuWBU0sHW+D3E4jm74+eZra+1z1dko3MvO6h37Kvctu
cwlzSDk7ZWIZZ2anw19ng8GaZVF0oFlikQe3EMwMGvVRW5GysqvxAE5TiGJKDOfk
Sh+MzACBj8B8tHN49pEoz9xTQv+h8wpxMf3o4mefbUB9bG+rVLFjIBesdmKIOFol
/7oJIw4OnLN9bcN4yvxQBEFCVB9ghkDWqIjUu3jaRNhLRQ8qFdEr2HL0UwLBWEbe
bnGvXQVMWHcr/UadInzZjTfmleWmOeez6DUGpo1W17OD2CpscPwu5iYE19n8WBxQ
jYqQBZtScp9l5/HLyZM3GtWlWwMHw8iI/ffEdhkqi63Eb/ZXp7c6pbqYnnkMZu34
s2GZHRWMDsG5DmmyLLLKywcsZNVsbjcWxLtWqXbHRSJDdhTAkaRtHF4jsL/9BYa3
iw0DofOOcWbrnoKyJNixw4FRgCHh4zoaXgFQj4o6PNlePwdjXgLt7S63nizss7Wu
IESGhBL83/cQ5FWXXRwkdp5eNK6adh0EA0L+Qy5s+DSiMuirGGhvMfhvrCOhLVS1
CvCUPgFX9imny1VVU8OcxHMrPSoqWukHwXePW3Sr+BiZIdOMlJz23zOuy9QPYpbw
e3GfBmipY1EmoQuqZxh9srSTB0rYijvIOLAyX8TAg38csyP+sT0fa/Le8/MqExre
tICWG5+EWjmo4eLmP9Ueo0g4yukaHJI9k+KLyJJ5MGXCQOndRYZFRMBUFyLzwl4m
K56H4OOc7gquCvUk4XCwLr9ooDlSPxZUuI4tojU5up6lMsoBuuRaROkQtuC0XGER
ookWQ0DKx4CwT3GOSyMwuqDoVbAIMHDqe0/sILiIWFI8GjoNZQMafB69Ieayr0O1
js3P+XtYQmpAp2QuoCb1PLKmsmtkkvrnSjNiHOLnPuCoi4oP2B1rmmTz1+Fq69LW
OVyKoae8tbXrphUOT7+sLEB5Y/ooV0X9TxnD9+0Cxvt/1bzIG5zCMwcKNVnGuPFA
goihSdVSdGIjfAGp2LRGSC/ieRuSvatupr8xj+ufo7AaVu1pMsb2WuEQ+JG22h27
DGfkoUoFzeyiR/R104/OTRLpMteCQZZcFAUc7GlmWUPm6VnKngYgfTcWjG6N2SIZ
fBeVOdHjZDU7zIYDvFeafL5LYILNI3iCYpUmbIqvKe5CD3JOIp6YODs3Yow7uwqM
5egcN65JegZ9SCb5S0x1edBfmL8mAAoep9cHxzdVEdNhoTl/NYJoQ+i1GSKLKE+J
nHniOgCXIZ7jQ7fJcBXQrX3ClTm6MUHIy8pqmJ9Gi4gcIGrZIIXneMaFx8XXMn82
AANAK8bcbWmMnQpnnamEU9DRmCgp6qjTxa1y0C1EMkxpNGL3UEYlfH+OEsV7+8ug
CFGAwXY5YdkE81IfiwifHSIX6tS0RxzwROc2VrtF5OZvrsDDtAca5Zss6GmLHhWN
lnOv4CfQHn7Zjj3UTfCJXhDCCfeMxiyZ1FHW7yV8G9zYT8Dag9bcjNOWElh+GDnU
Y5VV6ua035mVI3oJ+bz1/oTapGYAU97biqIqwDRf9cgQAUjSGCAq72T8rPaOJHFX
JWzjJ+8N8gK3jjAUlLzEG3aXjMjo3zcRcmrZC3HRdvC9BZKKCU/clMO2P7ptzpco
NjX6Un4AL9ocRW/Y1Tu5QeFcJOD6XcHVoUo6rCM8/QakB7Kp1EEfry4xQN19ATq6
Hk//PHO8YlXr6CiXkeinQU3BteS26vRcBvDx5feDb5caOZYaFoBPMnpb7Tfmk2cD
qdmVYJbSid/QnxVGXqJyYnSH53cYeWDmZhe8qgtMyMDRiQyTLwSP0TBeNawxdvDA
oRYt4BhmOouqRHJJdyuDVX5/6EYqElv3pLsnWLGK1HO/tv6rgovWthaaCzCz3xOm
oO26gALkRqXogGErScjVLjhTd7DyujuqoJaXSQnKoZmmeSIqOzJX3txy2vv8CF7P
Gio1xfyukcPEtuTPJ7mNpLKz134dOU5FMVjq/+eCtuyOtmv6yyjpSdyZ4fOcpQNm
9tjEqh/v0JKn8zvyZa54oFs1Qc/EwXa41Fjefbt6pXwlTz89eawl/VgY6LKYPmmq
FZW47fopxTcjFJRxcqgaaeanm6Y4Yv4VAbWV7eoSAinhu3kvx2WnLw78K+5CIMgD
xh7d9hp3Qn8AG6VMP+tegY3PrRw1ZqSOrP4VY6Pjb44BYIe5rcMJFlU5UstFyMs8
yed0/RBqbAX+I/c68nuBim/c0tTTcvREFlq0mA66FV6XdYVHT+tXZNsIJGugSQ8G
yrYjUhOOA+vIag4E3uVysUmLjxrIN3nHSyOTfXl26YtHm7naU2QDL+kmjhujw1Mf
qyJ2MNrgx3H0Yr4yheLQAR5n40F//ojdPH97OGU+TS04OgdSDlUsEQwugRJwJmyO
TVqdrOvqQkHd97ycmE0UOSNyMFdyqdVm8bX4rnJtCCMNtSKXG07JRRbUxgBrEC6F
fp2iLpWtnvUZpLYILtitcgw3mnuJOftfRrgyzmTuwKwmu9wONV1AmJJs28Q9Z7V1
9BxRKxeAjc6kyo15bdhKeDfhSVEv2dQMoL98uHUHjvAGu6uBvSVuvv9v48/0AbAc
XqtuZJG7kxudtwr6DCFGCur+Su0COF02jQYx3UIe0xoH2ojfFDMqanTYAmRsZYM+
d0ET0WqliuP+xstdNrolyw2+PsYFbaz6JOhwg2Rr8U0Wu+I2wzEV2wKZgpUfyIsP
1XnpTQUn1F5VOlYbYSn8xs7/WaSBFZCjfHCXnK+l0J2xm3rXTq/No9jJWc80TCab
BlRWbBrqEn/YChoDG4oYn6KYHVnF3sJA8KFhZx3O/Ipos5U27E/6106slyx/WvPf
qGtOaxMSseiHNWQvfY2cGIk8eJrp5NrZ4ddNerNz4kIP9919g7We+nESzKOuiSAl
0ZtW3mQRlZt/Ze3Drg+x9SAF3+Be/Mrmcm+vf72+VWGvuliUk9ODj1zlHjmzMqNT
/WC8h3Bv12luoJT6CTxVQ4/pLCQfpmCL2GSlLOd9Q8luc0HfH9f7SN2emVKvUfNr
fy2cLEY5mdg5yLa0OLQOPcOp2XbmjtGoo8LMGhxIFofShiayxJugGkGo//rjckfD
2YxfAvJ6UNF/TIXn71a5a9gcZKkU8toCUoSiGcwPhY5hOBMSu1n5yDWcM7Xz1pI4
nriIFJo3MX7rSOr0KiWhVC/NsccQB6Jt+I10lzk/zPDsJ6mds/If74hChiLN13tH
VBZiENkyoX+XADvfcfUecAMuv3zdmS0XpTlGsleCR0APkn02Ii43IHGtBv0ZrBUV
Ms602WUA+fyF2XeK1D1Yd+kcVvH+eoOXo0e0xmrRTcm5q3+9s7vCvgt9DIzL4Nhq
VCTu+vvpplCLf8I8zux3q2GtaW8ltPBiHO1o9SzuyVbOuezMRp0xerC7YAHYO1BX
WbdN6HHceyKZao05gIhZN/dKJ6vPXsDlP7uVHQmeXDWrHAEs3FpnBCxpUAfNUhsd
1klraNEzmJR3tW4lGS2viZ9wY3acNsnwjjpLPUfzFcqWlgFsJ0CJTUlEVBZxSAq3
qtCXMw2eIrE0Xibnq7fa9lJLueyvB1sFkjerWNumP4AdRmN0Edy54Un0rYu4e/HM
2uTRv7ArfH9oPHW0X7Iypw3XAtaJh/9OcPIPsAh1P+CvZtwu1cSV7ZGVCsDf3xyq
xAGlVJ9VJv78EkvKCcwhOrCejLD1iKr9khp0n5CO38pPriPG4KLXRKxFDx8uqJK5
mFMQXT1/owZsNv6sODkPtSugUPjaKBBI4DYY8IXmqBl5nPKT/XUu5iup5IlXOFDX
PL7mtrsvZf2OmtrSAHYAR2MEmhORdEM/jy9ecG3NiQ4Cyyt5mUVfDT3KTCoq1Z/X
93Yc1+QdAmL6P9RrT3e14/GHiZoE93BisT9YZR1wYpmqjXYfdAq/dl+v30IeR9Kq
NQRSsRxaBrfSxyBPIvCyXBznZJt3oVILni5GRWw2dHYo1atDx27O+MKGq+Y6KZF5
IIlLGvQtq6a2GgZ/C53r62MecHL83TI/0Rp8Ux5yHpCKolBzBmCBZVqNTPz7BSNj
oA27fI+UB0RRyyx+HI3zgqOp4A7wpfBDIr0o8W41dHIzqjP70cMBw75FiyHCcuGI
19Jg5inrVsg7cd/ll899eyJJDG8fRNWwitGbNcVztq9strZJeVtj0pqzZJnHcehe
ozke1SFs80TX4Y0iHfhR4GcuYFVlvQPHId6hQ49/v9op5B6DWwo6IQIKT75eKs7p
FlWbARdIaXxBkm3+nWaOrE9jVx3RzObrC2THqc2ySabNabVKDIJ925JjtKOI9sA7
6ugNkqMIUToDVCjCO2hcvnmvFBdOLPkvbv3XIbBICtvcOuSRb50rM83+4aBLn5Fg
RmrdTgb/b0huKBjFz1dQpg1WybZ2x8wt1Ogmqc4EEDkXM+jJQOSGDjhCsC3cFkaD
uwO2cVKYEsZEXPuSFouIOTe+8RP3xxiybD7UHBnjYQg+QDwQ3IDeLV/BAaZcHfM1
+VrbXUjhNEdgggR4jPJH81PjpSGTzsVgoWtJXrm185askwhWsPNLTTm5bx/cPbrf
SiKUpbW2SeWfFJzaZh8F6tuNcbtHgEFQHlWwBvACzkbqgJFg1FUWNHRe0Z+8qpVr
/ex0PRFykkqci3KhGCNUER4iocsabqqUvstGckVZlER6DyeAhnbc180aAVPF0J4V
Lsnh+8zseZi5kwjjonOH39ugIigj7lJhv10ZWjnTSutG1BkcOmJB56fjl7Cj1SRe
KBMTl0oJSWh6Zr0MScS9fNsh7zKPcoNLVg9ePy/hJBJ/2+r1i28sKxWHN9yL0jN8
XtOSyUDy/y0yj6M2xHstTqp7tBTNbGUjf423WjFH+B1brWEzRA4WL/sa4LIEY9lV
/rkSesPJONi04ysLqlu7ur2ja73J3A5M9MjniZxxEALG0S0mbcBC69xtDrXqVJ1j
soRhe0BdqqLaeiH2pTe10t/Kp2gDR1zAPW/jvyXc//yS2AkmZ7Yt9VlJvcxQct/N
ArtuNmv+haFr2n50ziiA1exD5qDgE17P/mDahOW5CudycQ//3pH6kRZH/1uQRRSa
wA0o8mv9CG9A8icBsRaZITHvFQhZdUK7AIZDmtgGydrQ746HFS+SfQAZ/eWJHCRj
r+Pzph196ga4qbd+4a3ahVzkmhO8G+jTLBOqnYQfKw9jMejNjCu/AdfEkGD066a1
c5vEsCBTHzUEnpcY8wEjTh4nY0YZzkNsie0qcwjDw1UVa3CDG8937NTFd3oDypXj
c8bunxs7kB+hwZxX7/cFZQ1kx2OsM3knJ8gW8LdwTG9Y3M7mzYuKVKxPVkGBl9nd
lyg8DNTuTrHMeAVYU5eCWVfgrUG/+ceyYI0dvgniDJjXY8jEbFKcO5MsieRrxpIH
Tc1XmtAwiZ+3nBXC3WQ8O3BfvVPjewLQZczE5DLjvGVvKL3RiXXdCEmBY4cIPAa5
08VIYoxE6Oq6+nOrhZzTyuL6jb4d+o8sL/fP+P9k4odBxy02jDuDzBytWhDIl7S7
WSr6djHXZU8E1VjXA4rqVJvbtxoThQbd/u940kBt+GgDbSLjdr2H3pSAS07QDPEP
PXMAzymgD4ich57MUnP1OXkn3eLwS+wF1zrpI2oyrDYsfqSHl6eBw3rM4gl8206O
DTNIPh12I511Il0D9RaSMHNBd1BaD7WoNVf7IINp7obPCfO63BMqnPJthr3ftlgg
m3Z/UD2L9Lh0NJiHWlUUYnwDjvEmXm7AubrtPiCND8m+B1BMJX/cuMg2fBqzrSFF
SAsclJQl8nBNaSIBAaQE3R1etWjDyWbUwO61Vv02HWop2I9RApOFBX1YiLh15p6H
Bld909EldyqX4LO2seXH3aNX5ujXIb+mRykwCOes/O70WZg53pQstH0Z+h+DDQgI
Jhu2rU31ZStVz5mcyK8UcOpyUcuBGtWAususXwUfMEGHW1f3I25wVuDn4kToFsMS
kdK9XdWIheDkXLDZRveASrPwOBINcIoecYfXnNikhVoku15dugKJHk6y7bp3EpIB
UDZVWFizImnFGIUkzczvTzK0mdOTUi+ueYks8v25bRjntEvNmAG4bXfmKe5f1NN+
kxY9XiAVXW5NpMA6cwXVyQSPW+L23L55+ijXNatHf10KCA8pe86UP38MPU2bVzcX
Cen1xgePWIjL3/WTQ2sIbAPeXwRQkVGC4fVDKZoS3h+oEdyvaW+tnd+/3P/LWsye
gaE/SZRZyNEHOFLUQDWorRx4W7xulq9nOTmDDThMVmEkFB1sB3UMLWZDs2IGU3XD
2YO7zkbIpVXUVxUJCEtXvhzjKJ46+kufec2yMKf427ykCrLTetfa1DR4LNA3iIRH
GSkvomt32OcwhV/a/VSQ2FfLaoNGFZKT2MlFXlTtMWlX1ADqcixB6dga+YTeBSCW
d+pxfeLhSxJ5BlV17E54Bt/C/cqRIK8V07ttBwM8W5olFL4qVLnR39diTCFulvDb
qAQg/Zx4PQVfnHA4IMnI7N4fBCk0UvcQyr1eyXemp0zpfTcFpf9MFyxQ5kceow/j
wT0hkEoT/1VbX9MCKsXJVbcRjypYBzOXXIg5ulNTexI2+JR3oX1vkBkIHMNkU1Pp
X17xladxferdUbbZOrBrNoQ9/Mt47ME/EJcQxJw2uKcxHvyyc6M7PrbEKPefpTXj
xQx2dZXdMudx0qPw2xLcob7CQdBrM6OvYTy8+odtnRSvsJE3JUnMNnwIl7L3LLQl
6EZfT1EeDj0t81CEKaeQv7E4cPXae0oTYZE4fxMLB/TdSjR/py9ds73vlfxzD7ed
qkR3i3kcgw6Zojgm7oIIXOzgNonQ9JEdMTXgD/KWUXf1mApNC0Z2igkEFpnnZpZj
EnMivlRAe8TIaQONAWlsNUX8aqUzQRBIKTS3WM52w1SSYHHX0/l/GQFeb7E513VR
sdUP83i5V83RhT5z7ra5xB2umS891D530lE3fwYsmi4vbwEcCo6dG2vCOGbyfJBL
T3ZQakzvcv6zeIfTjEgcK+UXT3DTiU6mjGaPSjYan2Lnqikw6xpw+fAOVxKYBKhU
zF0S58gAhZpGQ/7+u8S6hmRfVYTfonfhfFiiXXyHCrCLid7JYligrzOv3HPyQKhh
+hbIn+29iOhS6CpT8RpgyxLcd2RQ+Rx6bjTNRCJfeSk=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
iHvBjbtZbaNvkSGABjBOv+GbvJneyyrs4zNhqLZUorjzxUhq9woszIVm/UFjEl+Z
+093aYukdytfu8KypUUjIOKE8U/UvZ5uB6sJsJc2IUX0Yb7wAJWNDEg+ugOUuTqd
y4T1mln+Dnn4KFJiJHBMEAWGso3F5oSZPGspqCcClXlHRcE9l3uG7ru//ra3exTi
teWOA25oUxPy90LtB1HdsV4iCCHWrns/nuxWuQDl33t231OLN7Ff2I0CTBPfuO4l
4Kd4OROqpFLtjLQV65psx3DyqAhpfVEFVvutYgDA4kU3Fkm4HQexHtO5dAyelFts
rkieyGJW29d+d1V1bpl8ew==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6272 )
`pragma protect data_block
9njyl5DwmYTdhmWiVsPfgpJscUvUJRBdAXjLqGzYXs4fRi++VVfn326TvczRtG6W
62EBpKaEqvPOZg6aiFQkAy3kEdPd8h/s4J9T9ZUwddmeoxhzBm3BiezvAGHUdeUW
fq+Ddt+Hm7CafclCOx5Yi5s6f5oCYTz1Mm/rqJWyyUD0lW0K39osr+BZjpaA3GGp
4oI+BkKYZSqsuRrQshBPe6dHxlBUzELbi/N+rVHKLhU34N6eumeTlgf0E7LpfbT9
KLAMAGcKWxsCpl1AcyL9dzcxK20910kbo6/Q4ivJmbPacDCRQHPt33nLGpeCnN+W
kAY4Bw7Hb5+3cMemDspH/u6X5WV0QaLrQ7QS75vGTBRjHe3EiA/dfYDfbcEsq1T0
kSJnnuAv8fxGWG9q64sKML/mEmkkaDzQaKohOuwXUKGSzjbrlKE/Y1DRJ0Kq/w+g
9opBv0kPoKNobi7vGhkUfMDq4oRRcbht3xdPZMb3F2Bw96W/5/XEt0yaLyVUhAGq
VzqWky4p90nizaAI7F35xbFJuWx5eFyu8mAiQ7NaZuOJ+p2FloYA8moP3tbykGka
r+IXEcRuNMpU09u3QanpDUZaltpSdykPHSFE94SIcBhjf0fegrZmWTYOa+5WzQlC
8xjwspSgmO08Sq2+w3HO8wa2AZHfxxfpFyPwGPaRXoOLY9v8cBwcMhAWu32h/IUj
WhiCPUFbmZuAv0i2fndVxLeHwIJCp3t1TcaFIMFaNRLio+NABRaCAQQM/L3tgmVd
sRxgtIZweolvEiGHB0yGnkhST9CXXKbnI1DmIabG9Bmc6oNIudv0/66hzlNHhiXD
4xSXfd/TC+yY8NXhfHmIILwOIixv07tcFm1g1o0+PG5LY4jnVdaGclSBWH12iLpM
4JWVATOEESUHcKALDKFrQJAz4y43jEv2vlIaVMi0UbIrE8ofMsqt8CCR8cVwYWHI
VGLOEHMxjFLcvpOS/O8ljLlPqR/PQkaNuRXPeSWwur316e5N9PS/4m1PamMDPSOs
PYTgIOVe907US9htjeCrpAwnNIOPvTAR6hFSlnfqwExKkcHAHL5NPZPpQQg4B4d0
sptJICjwy1+J0z19gpC2idU3GVXfPthJOhEd5Pehrd6s3kPNy1Yrj15MJOriP/eY
gkMe76ir5j+YIJwFTBf4+8ych1chTXD3oVZNq5L+aWgzLJ9MOr5+JwfzvZu7mF8r
RhXuUs9EXz2c0LTqfl2akyGfsE4bofmNmh/1nW8iLJKnHfBvcA+xbuAlFNSjkBWo
A3OcNo+COVaFC2h2p/bUVl87gUJw/o1a5pC5P8pjZk0Kxsld0+vm7xLDGkeH/ds2
Pq2dCPPTobLZNhIzpHUenHIpEJWkkUeJGa88mOobFVyalowjdOyyLsr2ecu1ZdNR
wckcswVwkWKUA0WoIpkN47DdMPEpEgsxXqPNrrv/9erqS9olcH6kgvCOQhxtRwkS
cMgsxxcWLsUZkf90AFYV0Wv8r/4QWL1+cNtoPr4mi51dQ+6WW9DbTksXq6wHwuV2
UG6tddmaOqSAogrEZx83n+1X5Hrw25X+qjekZ7ldhUxCvShN+6I3R6SZnFXZ8XKz
5LaVg9Xv6tsuOo9PCqIVlQCFKLgQ9sNUFnvRJlvpgts4rn8gIhyKOLLcox+td6IU
//+rzcK45vNyPS8FIXLyCVnqGHp00KgtcAree4KUgvH6ZE4sYub2M+XUy3+KVWuL
fGUgKkLKkTpR8zKE6ah2IMOs6+nLpQi3POD5wuFodYPvzWcrNmoxdKw8N36ibxsI
iJwFCtXQN5gUIkaeQOC2a2LwB/pRmugbFHoBOSzlfRnFj3IcawZnl7Snp4OgKZOm
kTiPxA2Sx/2UQI6OCLEzbi9UFesHDJCqe3qbfaBb6lqN0sq7PNqudOIeUq+xJ1QG
aiXjkTSFS7JMIW9Nwsgg95p5MiwWF11QbP6X0XFlRVQ4jvyclMaQKz328DP8QUy4
8P6c3th6LleYfDbogKz4HBD/WeBq8WvEnV1DWjEgO71YqfnEuPZ44qGAU+1GqRXe
mpJrq2XyHrxJJHc77mwaTHC5QrvVtBjXmJ3RlRBvX1eJvR8kTkPxaGpHd4VDFlEU
82ykNlqj1jHGZ0kj4Fb85hiShZJxmre1wI1qjIM8pfDqhqfG/EMK3UEeunSOgGjf
Spl+KTxUJOBDQ06x41nYl3Wm5+PYOY89d6HP1WsI76hzZS28eBPoqQgVdvwV/uEg
PfqYygxvsBNdznrmF44tcY4PreWKHWcmVxKl288gDyZf26vKADUBmQ4JYp2VhNff
wyZBOQA2nA8+R53D6S5m9+cRBlKbw5wrqS9fxAzcxBUCb3Vq4fCD3c/OsMVepSJ8
Og5ng0H+LrE1xEbsZl1KIAfH/D5DWchwPueMVD3hDAfwcLA89ZnK1mbRyvTmmBOy
iX5uSvwuwcLgpkfuOP0/LLGutDU/Y8edxxqJGSxUxw0ipEB7b0M2JuFlrGTKrlc8
9B236PzN6qkeU+aH8Imc7DkDxvXbf8qYndwofd6VN+paaoprOlVCVlTVT1/5gbVn
uAWkW6ed5Ns9f2AJ9EMIvBUEG6SFpYUEoBSL1Dn/5TLvmp64FDxcHsRCOzpwpAIU
bAtszQN/41xR69Qlr/witnnsKJfoQSm4SgZny4Td3SeLYN05zeNrw45InDaT6rhK
/glAGLEfovqmSCspnOuvD1iK1K583kKP0xJFrkvk8XwnVeWD9GLw3T8oQVwEO5xS
jiDrp4BW81ERkpF1YA1ZkxQ2h+AXFk9jxMbutEdSEGi/GJpo0OgH+3sERcjSYK5I
GbcldVtNd9ICnD9SkSiIapFCGzPrVCtqVRm3rCKUdFOZV0BTTYDsH4nG5G9i8/uq
gdypGTzAxxa2Iy0ZD9tdJNERn+vZF7L5+uPsit5fEFboSnRqFABaF2ccVaOZC+dx
JJ5eOiVI31oVEueb+cZ4mULaOnu8e5VRv2Vyn48eGbLoqfEPacCxwwjTrdJO4h9O
xzvS7f0eZ0M6yB9RHsf0wmDKow6KO+DIa8/Nu/u0R7S++MAZuDEUwW9ihCVMBI4B
gDEbIa54cemOuL15Adi3JKuf9/rLHBEL2Ti+U2j0I0oGSsjPoePWURJFf9N7rP+y
D04mBvt7/hABebpC5PkYEIUYyVoIV1AdkIagYi6prHjGc5GhBSxVOOVEWYVFg+Xw
QFV+FUJ2C744oKqFJHqnEFvu+SmKukwj5y3qdBIYqLZFn3ZEQgpxH8gRpo6joQ1v
xjNxirXTK2wMlPOKwJf6Tbhybu3zD5I88wmRw4xkuhRLlbh74TX9FUOjZFaflQkl
Uv1edNwz83fF7V+pzJMZleM+j+35hynXHIz2ffx3xjNy0EcD1REvFIdqRqh3GIg9
7qr160lz7nwxqDQd0t5jJIr686cDlMaMa/1aQo8d4slsAtbmKUZuKxmEtE989pIp
vKVnB1I834bRFc1VlHDdXU4DiGEubP0JmGLbyXN7VA3WH1AXzgOJHLf5wmJ7C6vc
2sw0UtwAm5udhrxei7dJRTDqEPqdIDCSL/YqU9EZT8OEUgy4JouwJOu1SUFqYtKh
xlQaYMrdMrvlJ+Soy+jO/CLyfXV1PFtmgNy5P52D9ATVuVbmdK2OZ1LxzwTm1Bwc
3BJkCoG6m8XPwdHPJGcSxd+0xq30qUXM2EtlnGaRETqWY9Y8UJi4PSY8mvJBqpXW
u9FFCm1ds9s4LI6jPf7BSHjmS6mImeYzB+ogecPXcEqyfT8jZKkMi6FAClDIQHBd
egLH+RMMwiFLTwVnyCVdz8YQJDcG48KO/ocE2aT1ldFXaj7qRbPy7wpzh8fxDzbx
KIMFfArWL/ndUvpB+tkgroNLgAo7kp1ppmObaK/H0ZWlthoho17YcVR5JqRNA4wB
Rbqm36xzfIv9nmZC4AwyGvS4RLbhVbj7k0xPvUunNLo1UBuR+05LOLues+VWBMkm
WTu/QaPiwzB6udmgZlohl9LEQ7JL/Hgt0Z7X4UPyNHynOxlsE3GOjuMffvcUupRq
LcIoEN1yzVUsGqeGhiKrb7K22ibwP6487R0kD0FkmvCfZgbC+82ol1UeqaPhjhyT
8vUy6n9MWU1N2kIb7qEd4o4QrKSQVq97MttGX8Vh6eHLEnePtoEq3OzX8Y+DzZxD
CjMNUjgDwKgNavyYPQ97W3Lbib97BZ/CGqg5B7o02w4m42G16Kae7oRU5xdzU1Cq
y4e/gSdnZjVTuNuu/zqRXe8kJqkbNZfiT5KmwLQFr6DI51+kNHZg2aXR7RLSTp9M
uRFEPqqZFaSGJHQD3QcXtHPGua+f+01m3V54/QQKG7IlYbfk2E4EPoRAPi7wDVxG
ML9G0iOiipPUkESncK8ZA/TKVvYXaYczLdvBJqV53bEC5GqMH+t614JKY0QmM9Ju
vUF+w3C/OX71RpaHvO+rMFehnSMsY3MR9pfn1eqTKnkGAPfxmRwir7XPLuFW2TJ1
zY2hpUSWUm3wcU3Jj9kN6ueY88JA8mXH4j/mOKHh1bDd7vF6NbLeJ8XMeJd3uHqW
DT+KJp41hb+ted1NVUFwNHw/Qs4m0E/K8UECF2PtYlUuFgVfBmAB4AjWYkOHRMlu
7wy2YTKlFAslqboGFT6PYVEFHHDqHNFd/eXDwFy6MPWfFAzSw+ykefUNOpkFEQr5
tVaFzaAQHH4VSNcigj+0TIMtBVyQJo9P1ov386MitIqcASlzZijiGC3Zp8wXqYtC
YSvCnkkcgknWXitaQcewAQWrqx1BfLPuvgJSPtLzBbbgiLT/5zssFiqnEtqO9WNn
YfQhWJPwC4agoPrNRU1XsXVz7SFyC1/OKfbll/JlSAVPViHvo1/qqDx6ms81HPHl
3hop9sOuU4EG4hfffoXlGpMquMIb00k48r1vggF6Gq0+c4MCZ83gxxrWLq1WLDBo
22fHi9yc4DwWKsY0+lr85ydqCYagLVydn6QpkysRYndrao4nBn3LomyMGi13RcGx
BxEstImWu8TbOzhJ1DJ1OYAuAG1JMKzZiyCnt8/T9jDal0Ix3t0VoGwFJtxxB2rc
3kluiw7gUdNc/G3iev58CeM80T59MR5jSFIUvBiOmlv0tRuy4KV19pFvppLCNFqa
wdtwqcFzr0S9Ct7Gm5EDxa3gDShiOS0EXkLzaVbcaE6t0rzFpFiOizibvFd/5W7V
x7f0rfcINHOb0KmSYStrUUNzX8mpUgrYX1b0e0sDZCctCWvTcSnxEeDzV+s14bd4
XtxcJUx0jsnNK5mI+Elet2V/ycMTFzE06I5AlZDQenaRu4au/ngVusYK+CJaTlpd
vVcgIpdIbWaO7IT2aMUxmkRTR/aUliiYQqeqrKqPuxN315VXj4+ANC0XjrgIqAD1
ApXp9O8IJ7tlMNpINXhcuFKG9qP+1lbftSL45UfI7H6N5fudWBWXmoIrEuEYqFde
yYgiAbWj7Bncjc03hfxw+BLG9K/HIoMUfD66VjOIVrZZykQ8SnvJ2fJkzY0iL2uz
Ss0OAEM0lcXPc2JFbuQRTdYnJHLbSzM0kUttOJcmXaKjHuHota7/T9DYaF62Gfup
AToh9Enjy1naps3EBDTUiXu4hununeNHZIrLbLUeAIFd40gy4ZDznUPIYryQ2pfE
tqRZSKyowN1hf7hgYj2/6PTJhGdSvudQj8Avg3RnHd9btQ3y0VDMKD6IbbGRuHFk
SuFl6Wp5Q85Zj1RRhGQwSpo2IM2oGFiyi0RIQEhQQej8vP5q7nQuVdXL6bZZWCQ/
lCR4Oa8ZcqhG3XZ5BWBNHR+UZNoUS90j39KRhE5rGnNb3JxpP5pT/m4gEsmdPsXg
xAek5JCEf/Bj/VJJikxNiy3C/9hLuvE1O5FJ6X8S2cq3fbNZH6TJTxiluLj458+6
SetHkIjAtaojNb3TLOKt4ax6kXzMKl3dK6i5a0H808CIMIZyEkwInwQutQuPY3PW
6kVlg84gv/rMwkVq1+4y98W0cFPilEuZMDGdiFPPDmEci3CAD4tvJ0RkhpRYiOK4
2fbeWvtNXNARjIR3WfaHqK2nfxLmRMFQUrmSSMfCDQe4x+Sl5n3kKyXH6/dp6jAm
Yw7D0UJ8w35i5ojppw0rKCHACVyfWOqXGk6qK/DKyt4j6DRV3H0LddM/wSQQ2RQl
mIZw+B5JY8ndE6Po5H2HcGCgipmHfEw2jkLM5b0sV8fIK6GdmI84Acjq6ZpgJ4OU
57OsU91tJVN9T6r+yGLk7R7ozm2o3W8G8QVz0J8dBP3+yVrkgmtMFVALyfm2H95y
W1xcBLYXmumjGcZhh/3Z68QKVl7guae25GDEh+NVstFBSwfbnfQXIQOYdGtQ1P1C
ssfoZhdkZehfyNdTuBlbG7OQvvPvqQ5xQ4e//A28/1umT6gKbj2lC59SbPbvcZyt
eRVsP8JGiDqNZSzHSshgPc748JiKTYItLA8sqjGWkfsOJRJTxnlqoUnjpTXYJxP5
xOWuNnnMeWG1qiReKQ3sURwJTBDUIVTVYJajKbIWqFaL7FG5ttb5Z/gVn3we1wIj
mINmKnWme+NM/slyhLNTli43g2RN4wFxLAr2oPFk8+3zd6uZqcr0u4hsYptXQY34
2z+23TYkuwq8052pLfKkmozDXwZ0UQ37Kdyn4RObTsnRVSiPMG0XHiVACdxzPWzr
ds/RlkGdhKK1vkYwWCT4XxADTgpUlgvm95FOFTlIP7BMmpMSBBOCV9GRZWv3ZVyk
DRq7ohdWIDqODuoxANjcxlLtkqTvktVvailTwnBihE0puu1AYftI5f1koRjTzyYq
qhkfmRrVSC3+43rRlOKey90anoEXyd+cjx8M8iC3EttJzgOVE+n0zqmFEPhLDiTJ
SbU1r6POY3cj5zKPRc0l+sHuFSICkj7m7JpuklJGmqWkqBzv81lAL2JUz/5kn47I
0JiYy7GTyiQ+XqtxvaaYGTT7is0S6D1r7JyjU69Si+puWBEM++zTNGdY4uS98v9H
UGN5TtIgPlVQqNPOn9IUsI3c5z1r0LtiLQ6VAfsvqzpmCjqc25iocOfsIJH0a00T
hs6q/MsLIINX5p8XlT3scAmm/adq5a7n/KRK7UU3NKauXNp7sboEOkwDHv/puIxv
5A4SnnW9/iq9EhqBY6l6HaqC7yqIyzviMzAdI1fYY+F/wmZl3tEnj7snK4/haTbI
/eFEJq9WjeKuj6lUJ636yTm8WNEgt7FvATZPiQ7oSpgkYKE5FsJyGG31OpqbtjAW
9QZXXmzIv0Rq1A/NLm856IEG8krN7K8rx6ncBBaK8oiXTWtLUbH8nqQnD/iZR/Wu
eHst7rZp90kh4Df8zPeDCbc7mOqpCrVkBglOnC0EHQGLsqhs9n/1IHedj/a2Ns/o
NySzKlQue2ZMcYRD5wlmoDqrHIsnlQeuaQarlcdQs0tX1/EN3JuMMEoXvNigoW9K
qb0eD7HtpS+QRlONy7IiJFv5RsP6dIZfskUEPgxR/AOXhhM8dq+e2VZRx3o4d207
EpwdeWyooopy0QPjtkF8DV+XlxXGfuIphiv+IS8oBP92Wgg8x01W5DxHSLtzPcos
OUJd3Gb0DmDo72XrT1KAtEE5a96L1I6BzJzux9SFbgIXJQ/SzvnkbF8p+vgnh2Bd
u1ywMcDrU/+zWxNYgS81HlYZLbTaiBqFzB4kMJh4SrTrUe5hwVALrhdFduP48rpj
bpLrlzMUjQX06hL5v0cgCvkMU4zp9pBLZ4hOucrgMzgVi0/kf4+r0tPuuRLu9949
TQbMVURhBcO15XVc0qOMgm0wIfDCc5rbhNBGvC6dtP80tpfmTDmiyBXC7YSa7Rxf
uQh1iSyn1p4ci/IZPmEp4ncPJZ/74ewbp9ZsTu3F35fmho1zqfENztHLSfwvxOLt
Q88LalbSgBs1Mn74BSAKHhqVeCxQ85zpodjBVzuz8mfMIzKCyXCEpjKgLXRtiA/s
sDx5/fZCGZyntS8R0Wr8lPUUq1md2DrAWkUVvAXBLoR+PT5IWHIxOre7+fvHeDQS
vlEY9eV43wZ/ngbWu0Q62vY0FYzEloISDK6xrZBB/wBKUn7q13uYC9W3mTxcdwoq
rOYQAMuR0pjTPV4265w0fOUzakwvBsBhp8oPoERbsYn+qijgW8bUmQgGAJn+eBYQ
vvzD/MpYdC+W5nBWVwXoeszh/nD/Wa0spc9QsAYP2IgO797Cv2S4p4AVS+HsjHyx
8Q2ryWvAJ+LU5i4wp7NqKCM3ofQCF9m2H4slrcxi1aERCG0qYsj6wu1Lc/YlWGLe
R8cO4pmd0P08PmtV9gmilIs1gTOR4tu+JMfSF0t6lEwI4uw5AeIeZVpDaE1b01VI
25kYKwnhmZ6NdtWowRLJ0JykGQITKHppuKLry4YCBgs=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
geFjVMslQ+LP/1tyD0Dqg8bgeN98EGQwvnR4/xFEWtbv540LRaWkxyZGHbofhNSn
NMmQ+bP54srRv9+DxRKWlZhIc1m0X1UwDc6fFPmM6C5S4eLuQVdIgSEDj2txSSGn
a+mmLd25bFWmcekSZ+iJDEhRe49+lzlr+vS6ikqrdGJ5vq68qdnTT0dw864GeyBD
Kj/ZUhxug3/um/0NoCA2MkHX6p4/PbhUGWVy5DatEI5ejNDrpoP2FgVov1grgcrh
hpdSFDEr/ohIcj5KUQ4IHNqedMM2J11BpRPjhDtQAr2MprqqX3iIyLgqoqiMtfpm
+NZlgPNyVMYp03W5stPMaA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5424 )
`pragma protect data_block
dKD7u0oMOZNUdkea449oFhO8/DiFYHV1qx2Ee4WR7z6+7S/rPFHuck77wXMScYge
xnuiwdDd+STO4xNw/5NyjovXSG1NIJ0x5fDC3/nZWnr6oCJBrqx8V92KgWtphZsK
F7pqUbiAteiwBcA4MToh9QJHrUF7ht5pxKx/aHR2pSCmowAeE/6Zmc25HtrTITKB
ymnKssad81AEWs49YH6xH3wM34jTXnmRGik+ioizVXW/q9wI2Vx6SrOhuDmCS8RY
VtaTwybKFVLbbH77h90/LAtnCDFOcTCi/76+H4yQmA0p5eSj2mzwUHVt8LVbHZ8u
1fb0KdnfGmIZFeWca80MenatJsELawO9L92v6kNiQeCjDiWEoC5md07Jq/8zOLx8
PxZJGDYAF6l8FqQehA/wp0KH5g7nwq4AgfVSQVyQj6kU/T0n6ZAShm0P1TReuQNd
yiT3ANCUfw1ezozy4hwcnFz59VlDPH4oel2pmhvRihZqU9PHizMWLUgmNy1JRj1K
C8+tch+narKQXS1wCRS70GYOXbZeQUQmDo4HWEAF3khRGjgrSNz84GPk1VmSR3Ad
nPsol51Jo8PHRBYI+i4BN0UTOBQqQIbxk2txj3NvV4P8oYqYlmAAgElZhbnpb3wg
jIBi0DFJzxOjjdvyAGAh1AHovowVdMVQADfhYw0rjb/oA4sxyAzkmBNHiN6wS0jZ
0I6Kn67EDGiPsNH/XU39ihieKT3bSzSZYanjmCF3LBA563bgOcNwipFrVocKQEpy
eNKxsAs8vVhl4M+XCb5j9Zf7j6/srY+P3GAkvgeQ1NSFPepWZD3Gz7wvSTPu1k+0
vb5yQNHi6AcNg2JJbsqolQM8sENvPZEHmrMVTM4zn4mYR1PLHiPiZZAXYM5aHeYo
BqAt4QD5XW0XTpGQTfaLMqFLl1yKttXBUNJJ0tuhFCcPuFmAvMq3XENojZ52X4Ek
eF/slJsl0P8eRXIj9W6Blzkb0R10Y6zhF0Ty9sTcv7+Cjx1VXqmLiLNmZ/8Gl5kC
yFAbesgJ+sQRP69Fb5Isovc70CMTNzDAfTB4AH4FOhVT0LD/v4vqLdYehdlF9RJ5
6RY94UtTDFXB3DOIQs6BZktWGLgaSZF8lgxtsWiOO0Ynwxhdzy7vFzfBINUnh6Gk
SPgSUkJ7eRQebnTdcxc4G4mmZI1t+tvNfT0TufDo/XWCLgN/qTfNNBeYVHFX0iKJ
IVe5co1K4DQmc/uB7DUwx0r9PUXFpK7I3gySU0ioXxGIqodCvMnabYopIX997yBI
S06yTtjkI/5iU1dJpOVfNAKqAhBNkO/jYb6HaAYgjT3zDupr8sKH+d5f6z+3nRGG
CUVGUp+1u5aIXlsDCjWRXq5vf0JzE5BFuefY0I98t5nkuw+75zVI24u37rJaqfhY
Pl/804xm5Bj//MQlESteTM7fJUDXx6PVEZ/Q+1WQsHRAYn8xMi1/ukTjuIbhJfy/
l5S+yfYN+0eJh5N4rCF67KIRKVDRH7cHbAonp9lCdUaPpiVYjcLIBHZDVriL5YeK
pZdF4fjki35iYq8d67bG4mhlbOwroFcM/G1+PbuyBBxtBmnMNaWMpPS6OACgW1M7
Fs8RfYUTRPf0UYpmrtS7H7G9cI4oP5s7pY0Wr+ZscFBCEIwlKVQYd19E+oOFy273
xAlPk0Gaktp+HfaBJv1wqbHnssmgNz+XibnsArbZdxI4GRGAO+7nbnF2yfKYuCLC
/9eYElodxWVsFwM0snNsllMHMNPx/JTbgdE0MQsUXpRsnaZVfGfEvC2kSNeaNht7
xdV+xbTrQ18fUyVGRZ6f2lB4MQ84d3C7SSwOJ2egyTg5t9vphgN6V0Ei7o7jL55J
wp9M+bjfWClb+2ZWME0D2N1EQXzoKFZ1WB4UOFX16TeFdEWUFntP6wPNDdyLOitR
Vg0vQuE01eAEiQU8GlWmjhNpAS2SwVw9m5Jas6SjVCtSjsaDvfyZglaYr+hc3yZL
wq+k829sG2zdWNr1vz35Oa7vy833qkvWifgWo3gAwadrMgdtwWI2zZNiJybda458
FlwUY8yAXJ3QQ0r6rDW1VvOZg68VFmYPOi+643dG4qiWMmLtoyZARPQ+cEtO5cV+
oHYNl9hmeW1lvWMcakOnQhwkPQ61iArxrJUyqzehdJfMCLpPYMXpDOcnfl5HBWW2
ibOXM0S2jodJN6XHJ4xUFv+C1uMNpaEiN0GWiaOb1pC//umSd8p0Q3dDyI7Kic83
pSDbre6Tv4OM6VFxRugjoaUK3TMiv8YmGA3MT3soCbdl5niaCx6s/bzH5vIemWhB
sjxb1qot0mjzk+IkNpSoPsPzaedNpy/PF14/GRozB8nhQ0YyFsaiG9kLp6DI5v86
gzg3gbd6G2Uso+g97VPJJHJoa60Lzf0HGTmzu9UjYh11rlsHW7dinNppwb36mABS
7f8vcb969ntXaqUXGLFVubhkDH2IzgQuHd+vwKJqI2QeyBbP5tsTLEYeer0vIRO+
oxFw991HaHTWJcrtTr1slrF1tCjSF08k3qoWE/ECcZUfFoTA21Yn9prjn9MG9qwP
RcNqTTVcbx6QVHW02nZMo4sg/VzmLKRO9/8RPBilk/qf+Pzv9TDUxd9+6WQu8uMM
/fREqwxa76hJgkCaLjAS7kriC3PC9Ni6gpKO3YwLzZa1KHdS7z+cKkejju9vCkPM
edZNAeyDJnK711nDLtJugRGfhouAqGT2VzCOSL00KkTRfduK41v7uL2Lvi7bW30I
8oDyspxwCd13Jef6Ian+YE2wBi9rCKNjq8LB33c4sgp1Uhwz4kMLHFFcIoxRYJe1
GJaLTLM//VacdTKsRpgwTm2O0B1MFA/b6wkap/vByCHdZtj24cPTFqX4Ux9naQQ6
arAa0X0k9Ipqk2hKYI6nNku79gh1B12hp9HFFZO7ez5RXEEccsmtHYeWXbMMPLcs
OD6mgJOxRZNP3IF8lFoIIeLtu//16xS4YStqPqL62c3ay4QLMtdoGwF/Zxrdg9Ik
9AHX5WQfqeg5PnEcEp9ho2twjqVAua0BHwwAmOWTD/4M7ET+xKbu5C3/KldQUK8F
qfSs3fNbHtkiTYD2/wgqaHjcr3zxvl/QLxmu//xgOMzN0N40wQbX1Gu4MCngsEsZ
nd0giDAzO7UO3YYOa47v2y1seGPd6EwbDkGVF2W2mVATBWTqsOcVIQEb48jUJrWq
N9MUniZJeW7RBPVUTP6G2vYc9NEIvRVBNWAYRg+fd8hE09C0iU/rKPs7Zwz4EvFl
biEyzpUKbPx2cIkcZ0AT8g8vLkesqkClT/UKDlvUMFGQMXMtpSsKJQvnU59qXf/E
0aCs/culNbL/WebrUz+VS9NmfiQc/iJPIu9qBtWrHDVE9IU8yNspb+A4h31AQxSd
6+o6UwXsuUKu0qgo5Z/72a1OleigOZ0nQRELqTBM/yf8pDmkTK6fJQ+Z554UADQE
9FRe6cOqL5eVIf31nQ5Gv/FYuaAM/v7olPluKQg7rtnGqhetqqVby/MJVA4fQEJz
2W+ygQrlJ92ebSLJTNyUeBkELZEgHGT/UIUXDhlj7eMxCg6XSSnK8LFiV8tHMrWW
eGwp9vkFgHSY1nom9/kw647NrXu+ouEQCeIQkXxBBU4CidZ6i7H4P3E+3Un6wXHR
G9M7m8jAQDwWDfikaWgdD0NsVhMD1fjQXlmpR8+5yvOsIY0ey0VHyz160/2KhuWF
VudqJu6eUvo5QXjrzavj6gICfjW1Qovp+O9n0lkW7PUwCLXitc8pd4PykabY6TKU
tZnuIHw6eDi0Q5+Ne+OdH06y5YfdNAIaRZ3diQg5KxUL3HlKZQZfywMKGeoU9K1T
8Wr/KeHIp1WHwK9+qnXtPKCl0YMuvGS3bv52KTwJUkjc93TTgrC50VhE54d7EgJ/
GONbPmV9R/7bVd0bElTjW0tG8ILO3TGPUaF9u9LUjPUY701JkEebrYFYPR0UHisc
13sbLXg8v/ujZlhZyTF+PRvzgNuASvdAnhSq8CWCiFiB6n8UBCdGBV0xsi/Fwywn
tugVH85a2v+G5hxoscIWUhv8btljhGjNqe0wqtt0SukyCjivflPHfJAyZ/gOVfAL
YPU8WFjFrVcMjS41V3E5QI7dGIkRUL5n2ML0xjjJm0w3FQ+xU4f1n/EB5P8nZDJX
dIVFRqCpdPUQ8b+c1E6q+kGXIPgcuPB8uSbsK6YEFzS1d49TZgzJvXqJ2uVudgcL
wgNX5+E4By9A0EwOmo0JWi2bSVlWvBhIylmH8EvN7/AJCzickxoUyFEqzkTg5HQz
8TZ5zG4J2In6kqwkhUgXFMGrZPoLe7Hb1wCQaFkCXglwe+9ulMVXjq4SXTZnLi6r
/MjVbR2GEM3TQabvsTqGoUvcKY9n/RJ5cPcqwQQFxe1lxr3Z1RNC+HZksJBahIpT
YbI9EdxDT/lB2uJNCkzAE96AQ3uqTnjvnFK1+jRt/0urPRHCqkqNUarlKXDusyxG
VU46XtMh0uPeWEHeR6i6I0RgmHzXrguj0lVR59+0w32chskGNzrCFQi2KJfSES4x
2GF0OcG9g5t2GPdoPjdUwwbvCKxxqGJ4NMfGRGfkRMEYwRZG5U15pgIhRFFdsTaG
nZp+vN0Tg6XAogGQU5IMZPeAUBhFViMaa7xRz4fiwFmVw/agIGheyJ4GXFW9+LPs
xIWioUkINCO9Q10QGu9Or4drJZ5vesUA34H73Yw5K7NYgejkrujIhbeLidhy6s2V
zZ5s/XL1QrIW0sHr4egddlR+pHvsW0R1WG5hhSicu4k2/N6Hnr5E1SM6XvsMxKGa
2IJs+cwTYEGi/DkWCmxSAgnub5MJ3EpAcP7YW4iQmpH54uPG1GhXdyl7iN4NwdSF
wZ16ga2aHI3uLV6PDzOM0yH+164X3w38x77K1LhqlmKMg+y0fq0h8I7HP68L60ax
Hc2AvC/bAaes1uyRDscUOyVOGiGio5lCUky8HppXbWN06htxknGy4WwbkQTtHsSJ
agjYYwgaohEgFtJ8/r+S70O7P6lcqiRoAAKDz9294o+Ez/9zHjd+BF5dWx6Hj39F
JGi88huJkeWTtFHXXdSWUPcKi0YhqFNqlKyE34QwMXJ0JipT6o0lE4LW9euiydll
rwTZpaJSBxNBDeIWRZ0orwBUCoKjYLQTQ6PQjP8dIKr1L/znn6IwloQZPcgVQwhm
4grIFKJxxYF9jR2GbWRabkFhxL0rGqnqxsYoZEqM9XVIo2/KMTaehjBAgd1tfVvk
zt2zFWo97T0Tyo6ZZIGvTw7pAehv22W6mIXbCefIYcA6/Ais8iOJyEVRQiQhDmLH
bMm0I8VEdrucpEGRDR+4OXwY3+Z9paiYZgGhHGGF5Qx/0uOXCjYzHHI5lJqsDckn
YcCcEzFBDMIpELKfPLg8X85ef6JB5k9V2rZhseo2/QZZr+GjVBWarKtBd4s+YS/s
kWtO7HQ/xDqMN+v/JXPqK80HoSV/UDK4xYvIp7PXz8BIp1uQ+KAZR9jni3ltJon9
64PzRTY2iuQb6a7Ml9tkvnpx2/tfucaUrH67nzRoSDx4hi4PPujyHT5Ut5fpwjCH
c2Uiq2pCIMk6KunKEYP2bKUWUcq6XBm/SkzW817OCDDMBgFK9W73PJbtZb2mi6EL
qzZNZZQHUbDx/OUkvGVbyOPtT0vQwd2JDSFsBSjtVikUpPiubcyRghvE3cf+QMV5
YCdRG8tgDINDlKh/54T71KhIQA0Ok+lcl81Ps9KTFSOvxAqqStA2oVzN0wZGh0PW
E3OGqyPI+W7KJHrbId6C8Rt0y2zoN+08+HjwbuCXDWa79YinQh1rDBVEm4HK8xoz
SaK7nDWQ8OtgNY/1MkEGgkqurdtGxEU+IPyPmGkE4xSACSXeGxgYchxfZYAecI9T
JfrAjY4EunidQiZER0yMuhy2bcP868XxYVNOYSFku3+Ivhe4Ozd4cIXj8sV/Wc9w
Wrq4Dmep57jEL52ZrdAC2Q5AqQDs7mncJHOv3GDL2qY5zs//ug7Oq+pYdiQM1P+M
F5DkOVoL+jeoMnoAyMI3wiD2/voVCU3SjqFEd6Xc++APdYRHvnQxYpVrASmyDYFv
8dQy5rxCwSywUoo/h+Ekym45NmebSyYim6hwErpXZ6FngfiB0CKA/K90pFLFmKMK
FOK0zZsb0pq35XZPkQkr/ifaZzxKY7XvQlL3KtTzZ1m1em8/AdQ9KrC6saJUaJI3
xKAbc/kqsmPBzoUEneG5eBepmwlc5gm0c7NpVbnPt4RKlVubTZcRKgJ3nw5lqn1F
0CDRqB8UhaUisaiFDojnZ7zOX3pfgoaHm6vmT5mgLPqEczY6oj2oyvgOl9pqLDSJ
KPpVf6xw9LUYPEybM1eg7HfGlBUiSfiaruvboSA375bSCje2gA75FIwefhpA/vwo
GzTpTWWbV/4OdcRRQabFI9wvViRLfexSclaDiGtupdlMZf877G4nVuasuZ7tKEny
2Ch+wJ6VGpjxLNGjLpY0j8AZG9ETG9YMDoYGoRtBLZBS8Sr6S24BwSd1wVJgHx2a
BUrebp1Kc1YHCum7RUXuPHHyTqh4NEl0yWyyrasCReWAPf8x4+Kt9CtpS+LSlg2m
LIzCtSRHTOZpZW0O3JCy5epKqh/QOBPK8155uSCXy8kHRH7PPB5U+GuJO90x23kK
4VPVI3TbjVCt+b+sP/+DyJ3vXN5nhNwYm61ZeXsAJH3FU4A//E8Jn9aLVdu8UtjL
zQL8u/IODlhkK+IYqSHwqCD7b3RDeYuQYpgQs6rm8v96nWejxArsPAzdjNaj3f7V
GZDjq6+aOwJEKT4ngegtmDxWwVRJYDgpJGZBGWZHKArue/aul3N3aJ2bvTzc4zZ3
rJVhpkTsOkO/2rrhUU4gx+hWA5CNqWJG56KZuIbjXJdqxAECJ/0Z3wMEUlFuINny
sejXAe/MUGgb8h9lKu7AI2AuJ0qMZycqQv+jEmwKPWBY6J41qBQceWQH6VO7/vAJ
/Q+992DFQMVcVw24Rr3kqwFWgOEs32a6mKqb/hXYOMFnQSKdLX74N52JoPFKR+Ho
rT6dCNZ+3J2jslylbdT9vlkFtsokuj8PaYEIEt8V321Ln89VD9MV/VDPjF/IMrwj
IoJZdnqRgp/LnLd6dYWc6C7cdcQqrKQbAYwN31ps1SDSCwFvdaApsNuzfofsqw1U
ZlpNUNJ0vGxuqI4ybQBuLMIxxS29cBo2sbZ6IB4J2qR+QizoaC49DRVH5zJE+MDG
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Dj6ARVLMhu7OIIq4oBVYMkb3hN2u1VNhB8XhsIvaKLd+VPCnHagcnba8OjXyyVcL
uYOji2xX5NNn78j0OCH43N7Ka1OKwiuGk12Lo3GCUSYY5AF4MBwqKpASUo0wN+s4
gMzUByOzDd0zCasw+qcB+aaRrxe7syptGNiHVX9Hh0w5+uXNsnjUbz+rJmi1aBwn
biH13A90L0qFQUjJ7hsp30YvbdqjlLTzI9s5wNVmAynSeXywUSLVv3/Wahn1LwEm
Oq2pTDAtu0p+01TArHoSWbx6zdZb0GAOML4sNmwPxui062B8gRwo94Xc9gtUOQWu
pN96xOrnUM5l4hGDVKqTQg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5664 )
`pragma protect data_block
kpFSOQB/WHNXLf9r/XA5R2Kg8QmAyetvzzfz9fTWBuUt561Gy+qXSKVbEc0FROOr
VHElFjx+F0c7XusBCgXtOhz/Qs+3ERIqbHMZKMRKImMSbuWHbxPbdK1QQ5M3F1NS
BgUU2KKGooeD1g2p3kV0eQdyjAjlNYyPzVjQMar+eti8XMXcP/uU6pGxPSQGiNnL
gRiL5DUbAekFXXTpSxQ4RUH2OtOnSpKqLzYOPvhXtizXicmXIv1jHcw15NYMmr43
DYN4iTVRY4vbZA7yayTO9xSUsFumKjuvpLzJLDrv7fAkiS3I1pAIPMocHXpa6CGM
1Q3Kf6vStbVjSBcoWQOJKGmcFV6as7eaqnu40M9ZWfpHBJCVW7ucBKEyfTAXSIM9
DuSuubaaawy4E+oZsj6mchmCAibZEHbMNOLtsBCgfwRRVvHvVtCo/Jg1kt9Bz5a9
FjrdB6fPLFX/DWnhoHKulWBmZoWFsI6RfP1AdON/jLBNQpvD0IGOy+aLcSy54yXP
66g6tdjq6jHq5PMq6KaQaUQ9lhy02NhARALBiqnIPEQ42UvPrgUVnAQfsc4TiiRl
FgO/xtoRgHjz4db/t2OfdYM23byGZsf85ro5xlCuNkg7iQbWbgzjlM2PF8f8g43+
A2He8ZbuCvr1gJ2NwxxhCnnEiReDF4RK4VEQ2yNP7lszOqcmuGQK1Ugr0xu7k2f7
Zjc333eZaYhirBfYCRouhdPqgbjK+HaAcaE17bBXytcAVQaF7ae/pw901XoLJb6D
5m0yj24r9NW8PWJSPMe5F0wVkGtUrh5NoTjSK8Xu9m+yReXxPAWRC05JtuoIsMyv
mSvurZXHDuLpFD/SnCc9JSVB2YcTWODPcCZNkB+cksh6cZmYX9jJyEAzPH2QoY2O
4sffjGFa8G96S+/J6IJIaZH6D7/L2ZidCw77d2BvvVkl+ipcGODMq0xKUaAahD4N
3CVISIJKaPhtpGseTjx2ntxa74B86+7OERZ692NzX7yLLogC5SiU7ToItU433c8d
Qw+J8Wq1bZPo0EulW2XuYFxCb47xopH83v5dW8BGIMV7H33TR+wDCYxhmraheZDx
1lKdnUgFm8cMs4/eVWw8CCtd+7IL9Sp/Dbq3y4JmJxSYr1Hc9e/3lopCLCwGXe75
P3Bcl/UQbGnkdUCgKWaUeT6sqLAAwV2nnLHr6OWgeVOf6/w9QBq82hZtxQF85q6C
HwqVNiuOE/K0OKA4+2uVqr8G/pb9EVkC/h6u/IEL7RDixb/OVxy+081oWCfxJhiz
7suruhTAmGyna3huN5HlY38uZB8d3JKG2hm5f22asAxHB/NAlnNOEUlvHRLIO5us
zJlejP2yibHwS1VMOtb5apTqr93MWtvrtuatnIu4dDHgakSQM4IlH4vIu5VQgymT
IxGG2ahPpTqn5HcIo/rnkmhxnEXFb1ZcFLcx254HxSoC+yWY1BNsyi1XQvBMbHuH
2skP5U0fehpJPKDsxgkJbjvT8Tbw3eSBetppQPuFh2dK3uBu5ZByD56/E5oBFdNe
IoEXhqfdm9z0iW3XF01pHbTZNo/JwwwdtrZ8R1g/Sd0sp6/FS69+oVSYGfZkp6bC
K/q0786zMXEHP0+l8kOMYJ6e+Pg+9MeS1sYgoAnERqHsw+Pqc3RgVK6b3K/lOmE4
84Xy20u1oXephNTzqq6N3VaG9cMVM01rIrPQzk2jeuqMRuUdtOAya0FkZYzLX2E9
sPgC3HZtE+xREwJzja+OAabAK6EZMiDBEe0OZ5FpQENEg3f8FyKNDvIKn56D/fJm
+UibnJKfTBNQvuJP9Dzhx3WH4coSFdQoNSX1l64XQ1re6TfkpGmDrZtxQjCYpePJ
KC7nUhlo75dU3TQQ1sOrVU0XngRzugPeA2zMCtxjChOC4fGZGD+EDCi2rPsVxg5k
6FL47MiG39i1Y0FcfpXrETb+rnrOogye2YSiPDRMWQsJLx8ocBg5xXnQ9BqvFUnZ
Jym7nHGirWNJKICRNcv51eBDDdO3bAbFw4VYliWe/kXzVqwxJtJ+ubgy3KJDZdPs
dem9aC6jI7BkxSrhloeGXNiKssfG7O6qqH5pjgXKF+VFatgohxGyzEvKzpafNawq
wpWwy97KbdG+4ZUjsSOdB94uHIwwf1KYtyIHu7QUKoLqIhTcW9Zzh+7TY6k0QveF
4Ek+WSb5UWNXDBUOiUF+pqFZlIyVUbxI0k+hHEVnPIkACvCA/nRRPkw9tJnEAWaF
hh41ajr2njcXpjP1cngZ7Xex75t2JkHjv/q+Hn7ImqUhCLai5eOu3tjvNRfBd1PS
UySrNdaptxDMU3EiLB8AihF3v+IssA283h7QqYFjze4op19uk/eEBkKPTVtpODIi
GQBmGF8hDQuoSXyRkyFLsPwvnzqOcDsg1q4EplZxcd2AYXQaxNzd/hH9ZM/8/MSj
7LnpTLe+GlDmdKqasZfUjRj2T1nDVBSEnpGwy/3IMqliF0cIA8216jcgUoi20XGM
zNo5tSpd7Q0R+L2hjXlcMpSTeCJoRWFgfWLkuVf5YqGj8qFZVDhibxvu1X2use1M
CR8syz9FUevu335UkHKE6Qgla4KvVAOz1Sw5tq+bzxoFVGRpboqf0voDm/GzFhXw
reSN441z0RzXcyDu3x3ytKpQGggQ6BiLDmyjll4xes8S2kAZlWkap8kQOsMQc1ZC
p7hHNwW54tm22lrIysYV6UUhdkwf5fqkRB19xNb1R5ORbLpFEdQfz1XJOBi4R+2u
sY1WOa7sKa6pT6AkiDvp8rDig19t9I2/89QJ+kGTj/XqvPgRloZL1QES3NLpz+X/
Rk3aB31MMjWzU5RvpQS2hHSaDyYSjt2OH/PxZHmMRgdPEuG4yQJgboU2mm/+zbD+
AE1gKj3SQm7h5upXM3Qep9TdArGPZW6CEX6Zut2+HiKl6fTVaK7iNSzdF+4dpVYO
bQ2DsKa2fzOmz7/OTURbKeB36XGzDBtWPNrglXpfuaO2n72HJbyexsxnS/FTld1Y
arPw/JwKF6DSJH7EJRaf/IVTQsWtvOg3Jjyt1VJGAxriEWDL5HlM56g1qJtV3uG9
2vyNGfbNjFKAhFUnH6HFeqqBKkPJLskV2IGAIk2/E0Y6EzdoaPodr12ynjPf66wo
l6b+/FYdRpKLdkIroxVzRw1q/a+p+hBqkBKj0Ze77EXyJqA8HIXU9j0B3zw8oX/5
hMSTGGOkRqQdXtSc09mwlUGOknboz+5dzIBZQL4MXRuXmqu9nHUZS9FF30Y38Qfh
0dqhHWd0lMRk/88y3Xbume/xQYATeF9iT4ydpMIhsAWrhZjbTGgif940aCSfvLVr
kCYabCs4sJwW4jpxjt/edT+GPkHc2xfGYQZxl7R/C4DbcSurGIKRlH5nHwn9hV82
MmqnGesGq7fx2LjjIHrn/WDm5vIzpe5NlTc9Kao+smOnM7YkchnE3q4D4QgH0qFq
EcVRko+cxuyNilPtOorPKkNtzF4kkWY9Ssm/KLpiD3poOpyrlOuhHsHeGN0LgcI7
xYSpQZgIvtQ3ezvEFDDI/dd5lHG9legwYlfTecT8sqhr5UDlGMlROjXeV8Q1U7z6
4eoGpD0WMccJbAs8ULHiw+9jJTBDc7LxAKRaAL8zZ5yeq/n+Tw1pLkj/W2Bn3DCk
ylnP+h5tmihxBalgTdJONZKiHCC5VuKNaBOkdyJa1jlEH0lqq4Gw8IkOgK6vmWbq
RdTtCQtTkIiRtr0LC8rorR2TNpw7dcC7iOm1XtnUREVcXZeEhOX/zsYsbjWABhbp
ARmvCsfgzLSnFLBHc48W8AlWB2JydPFC76Vn6tiz1iDPAKGlneB6iob2Jv3aJ8gX
oDfLjyqi6wNdA/Th3eXP/24SB4NfmibMqkKWG0EgHjCc4PvbXNYUA6YAvEkVZb6C
AJdhSWi3aCRtD6Xi1BR4KT10SaIalc2RBiOduz9faFqrrE+5NrY3qoMORNWogher
ptasDYgyfHih/XatR2ITHCAfmhw2YIByOPtxhSpFo44rXK6PF1/LYvLc3UZ3mXVa
o6FTQTAE+esI9et1gLUdG+ebvTfhOTn0SxkU2ILG7WfItezsS6MXlb54uMPAB/1z
AXHqV6Acm9uPgHyxZfKdSty1GKDBhiljkI0Uv8ES9vk/x6Nl1wAGkOBsKHqh8m4G
/YV7Q7vMc3omT7QG2Dr/siyP5cVcCCk0EYy4zQtvqgdJN+K1OYc+ZwNHCwTH1Ixi
BaZifqNBik6QoH1tK0QMM03o08NlzXDMxhiCbPxXJ4Y07nAeNqCIBo/BV86+us0V
7JLLklcAAcKhR3mxyVxO3q60kqng3rr+THq0Cx0W/LU/Tie9+Upn071FakyKMef8
9JufNYTywbZHM5mPLebpU95ZwKNA7HwnuGCHKiGIJ6K2fpRNQ6i/wk1t4fcYhmZq
jz2J6xchYUb2MlafiC3bVVZGWCj8xT4xn2jFAcTtwQg6g2rQo9df8Pv8xaqUePhI
auKkWE7e8Hw+pbgmySvpskodsJkYmmWdtttHhZ+WygR3xXXgsOsEBdQG4ObvvzGW
GBTu5NAuv9am1kfvb75hYvZCYxcvBFouTZ/2AbxE7PJEnmEmUw9v6m86h0BdSlMG
ugve6oUJva+nAyXTQAf1x6IwyMymP9eyiUd445HDO2guSLuEQbjsE0lNkqqW0Cmo
V28UniUattbwDKWEE1UmLo2NDfAQ+0gx46rPyQJPPMKl3W5JnCuarrHBZozjtMim
V+4GeA3H5Yj52+Lj/z2DdSkHKDnvqTnassXkQT0aace/IDIx6mm8gGNwaG+RScgI
zW0o/t0hmkSQMPt1vWH2YEHW+j6iDJEjYhOiIB0iDYGGcT6ZCcfEl6BJGZ72PIP3
aXnpUbwNgdfNpoKMWC+X+hYZyRqsw62a5RTNzqqvHa7ZZea94FNE5qlIe248EfT7
ixyBzBldZbpYoVAzBL0sLjSEOgEe1UwKxiRaGkkAt25ArcjTxq40CQ7urJJKKR68
bOfuCRY+LlMwJE+kFU6yPQ3qC1jrmcEnxinKkx9Uj/5Q4W4dKJ2gAFNBcRDm55X4
iJD5UDPvpgeG1g2W42hG+ZvUrIMb5fooOZuZ5IqygiWrGo5uzgn661r0/AM4PHwF
uug1Y81Jm6XAW+a73Sq49p9Xn1rI6SKNj1Y50aeU4RxhdQHmBWRYSbb1ruvEb5Dy
B7mlJydhsXYIZFviHkVP+7D+DSnBJzkVa86xivfsgkp8yMkrqSBzSOWRi0Pl9XU/
dmnc8QnALJVHNcp0rLkpDsjRK3gH+0kvxhd3Uz6Cl+Kzw7vBBqa2wyWzhWA6YhsH
EbsAtmvblTV1Gu6UQZBfKqqTS6OO23Fv4QUxUNx8s2eWXKMqGbjeYlDU3d0Hn7by
Bap9/G5hmkhfEvfCRaSw9qETUo99rmoEZdq8weVRbJ41qLn0J6yhXI413dztUAi7
l+t7lmwi9YZYSdl3oRkasDqndPxoOgmE0j8xM8PSN0nB35sdRvAkVH7MzXhEihTa
8pKxVbdWXEXO3fk0B3e3snj1jq+xBHoiGWd1vv4FSQZOSkshafgVPTmWjpWkc/qD
tiJmeXNZEVhNlj8OszW0xT/ggAYbUVJk2cn0mVP20SV/JbdPWVfLb0DXvQUblXys
nNefa/3CDTHPI9u3FBaN2z+lx6NKHhLOxfmIiRpznC8j2D0q15r1KJzx5TXr8rM/
DolF4vpfQgk37XIFSfqM4qRO0HZuhL9HFXQmErjSigOevbs4agqltoWt2zksDnhq
ehY7hzY9pLc1lizOoJvoSz55R+S1dU3GnLWenbcCK6T+CnifqdILetnX9JrsNncX
GlT0MbjMFrlqbpoptajxoH0bnmdW1ouk1pwdZlk7dfnCZnam+pL3VuENyHzM6UBD
pGA2bccglQ/msVKnckINAxLubCzugFgqcAHyPW1HmC7yjE8WN3Gg6Pu2Os3CevKl
CR4QqVkSiBH+pk4c2NEbeTJwywhREEgv8uxP3IS/i7PUUWiXORPACdFKSzgthMoy
Qaa5QTZOH0v9TXvT2k7yFh6fG15PSRdfNTsOTr2WmDT66A4RqelCUtMugbSfkhSr
wP2SbYggC1tBuozDsqB2CtwYZU3zxhmOgrzC5DIrgSLNrRnIdnEy4NzJbH8iYgEX
ivYxfyXz2KGs3cH9wDThFR/wB86PoDinBI9gMBo2IAlflNvABb1EUPP2VsFMBCaA
IjOj4DD/nIs963JfhsApOUbnbLgU3Jwmq/UyLm6p98CgduPcQNi2MDxHOfj5NfoV
xQVFyhISeE/6hsvA1r1BYjYGeci6B2/EV3HcW47Qk6zCeisMY4VAI2ZJ2S6zSRrk
xF5kQiRfHl9WZZP0qM1qDuUs1FO8w9Xu8r/LZtqX9S99wLoq9hC5dF45883j7+md
Nb8GAASMxirpQsBs4MikiMCMfVIMpmq9iV4l2Nv5AF+J+H3iOlprg1PZV8WUZjzx
izvyD6ofOuxE0nhoumxEtrLcILlZuqRBpdJ+zOsmvK49V6obg3YsRwFzzmS+H/Ox
krzG5AbGE0EYo2R9sJHdb0w2Ohrn5DvDLaf++XaL/MKPZMQVWY33a4Gui13E/J60
WlIEpJ1Am0zGVaxri6ON//CMQjyJ2NIfcbFRqOtMsyySSpOJENQMPmx6Div4Ds2R
iLqCmMvnBRbYON+hhV0XZr5Ukek/t/j5qccahXU7kzBXSBUIFVxxPOYxS73HUnPf
szRaK7z3lFSH/+JiFD6bcPLu9UbK6poLFgwn5ymTYxMbuzHDUpZQ1/UKobojEBlU
POiT8yvTUf2POjzi3fBX44dOnu45FXKaQxK3WpJkC0yXA2xOTkng4vo6Sf9/kloq
wadD8L1+6XN/lqpwcHumTbSBpRV6/snBBw7s3tpNiWOhcv8Zo2OWS8NKI8TCZ+qH
eaVQXJAsrWlWWD6leC0sZL5KNAzORQWYhXL72K8ioulS8Rgxs9pWer607UAw6/dl
X0qPspB4ccFDMBMpzBVK0slYKTR1bd78Zt9pliZK6dw9xLb1+H2x/6u1tvwFj91A
ppDol1pzALQAyAqwtA0qOlgcnagQtr87qHYqpFL0No9gVhKa4gq+WLz0p5ozxsqT
6jA8vxLcPF4xfWRRHgEiD9VtaeCOnTP+DZk7LK4UfQd1MXJPi8hY0MMnZ0KdetPh
gvbUQR5A4iga1tbUgOt3CAO+KoGqCROEW85h0cwPXCgg1BETsKl9oqUt7ya29hks
rHr4YVZw9Vo5dQ+0LPFOpG5ClI0NA3HERkBth5ld9DA3gj00uiZSkY9VhWwW10Xy
bQvzvTE9Cly/+uGAinzVkbIdUAVuG+w8sjywpNRy+RBLFjwiaseWtUBmkx2w3OQA
/lzvREys35qGMtWwf+RxYnA5J8KVMKvj+JSOJtMD2gAzFnlSgYC8wFYujIux2t4P
Q8gA14ZT9cSG4NCy0halfkjCNgTOOtXKuzKLFoYOJUkmebo6hZ0Atqs/dQrYeSO8
XtJVvkpjxLZ2E5APFXhnTE6bomGvXu7JJc8s7VT0uX7FLYHG20pHIqHjiVY0ReRZ
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
O9JvEnn9GqFNIGJZ3p6n2W0jMle+zOUAP0NDfd5UONIZKdx/ER2HWLU1fV6z1jjM
aJvrClDs4UumrBagwfZOvVkOhB2lKPq+32ZYrkLwS1zH/aJe0julK3B7EUgwDI5l
c/El1FVSg0nJcaZ0G5beB4+AsTdltC2pNI9/ioZyQ+Pcl8aBihXTlUiXOlF467sm
VU9WLjOxEEw04QS4MhgaHOz5HvhAU8TnsCH3nYbmLz9uTfNnus4fKXtIAXfru9Yu
RzD75YmS7kJAMUgbOk0LYJZRtsEStphmd5+3rH+6No41CNaa4IzERZ3glb9mJi8R
ZQoMORMQFVuMDLs3NtTiUQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4720 )
`pragma protect data_block
Zvb40ahLkDR9OeCV3rmCIGdNvoHJK48Hwopc2kvQxzLdgf6nI8M3CsChEj67imqj
Z3x2az/rslTfzbw+aTe513eIbSewq82xESBxA+8JfR3dDOLkQjllBk5t2XOkgDEP
C+HKsHx60Uu1t+D+13VkcWf71NC1smtiWkhTVSyYxTgXbFosVnKlknBis6yHByMm
p4ZSD/6EV/7RVZ1Bd9bJEKUBGFUauRy71GLWZb8qoKbHz7NgVNyyrVB0gakypd30
xPuKZk9jOQZ/WksKZamDkYRK+npJUIigrLlIhJHIfJ+UoAUUKNif4UXjGPMrr98t
/SP7aj/nbJyjDzjFTOeXUigxI/LhMUJAFKjKiYWM/jD3368/kU+zONaxhZeGlRRd
ER2axHAct10oHQcdoUpdRFdFOjHsOVUZUa9RvgMpsd1+A0Hllcf28XXMYokumnwY
hWJWnP6VmX8MieHaVmD6CA7lCV8++F+wPjsL0yYtHkN+F8qvfHIQpb7XwGDcEMbj
lZYFtao3Z0uebqY7kUpMHqYk82Op49Ana+YXzU2rs/PYl2Qw6HfWc2oL1EU6S4nf
3Cfvda5QY6D18QAyDs0ylQyehJ2H+ZVJXPJD7hWsARqQDDqQFfErYkKyapEhL013
PxLNiqQlPijkjCm1cws3fSoaEXoeMaY0WBwTQ1QArAcEQPNOzhGQF+6GewfRb5Wm
K0gUMOXyHCkw1HMfUoxk02J01oAxs94yPKfbOcjm3m3vhcCIrFT72XHmv4JPnEhl
oEHOz69ONMBAIrDoLnj7irUQbQqIugwlP9cm539487bPQqD1WsFatsLARz8lWSaZ
RWcNwl29a6hgvp7OVaZsuUss6NklRNco2NBDX4L49ExrZzJuzZMU77NI0P7MFpJm
HcXWrCVJoicj2rbe8JBJ0cpke8SRhyDFBJsf0gCRB2Uh/OS3r70hWZuSOVA0PTeJ
JujhXK+28dEJVl/5fJ3d/5165GzSFEi5yQ+cP7q+LgO1idhbjiQRePZRVYwAGgQf
hxZXUKnx1EQO2Ee0StqG+Rtl8aDMyPFjbe2nE81US4JWeon0asUZQbmj8wGWpNMi
OHsvz6dim44qktIbjL+t19Q2t4ilta6er5NM4iKO7HH8yWXELRCOE+3UDAfpd51F
0IcwoNLhliq6PQDCMYIaovYAH91ZQshMKdh+wyFRRiEHob/y9toTna0t3D0d2l1H
R8IPY/c49x5MufsTBKqJj1ZI27U0OCmhuynkJwDiFKLGD7jjpBXBKfLPXXVA0Qhc
pL38CkafjUeIzo0gYro0NzTdGULSX8WiYaV5yu8MNz3e7/lP86aVbyZ8Fl4PZ3B+
uw26jhxPiQ/vEmKNS7G/Hemw4OLJHlSBYlQn223ihGSFMQ+tfKgaPBNT2y4HM4s3
uHN8A0s8loiqqK6/HFGxQumLcFZFfs6nWM0Dhajm/a3DyExCZ3bAJrr78nLetxbo
zUltoV2IhF4X1SVKgU1iR033pN7Oqg05jfTMzsp8/UhD8ASg9tMP87OWOm/AyGyi
t6L6AOQFwsowi7KEHgD4UKKj2gy1rNjMUi+8whPimr+0TmY/3DSiTyo8fvi/RbQE
CUSZ4qFyoRtjLs8c5PC6xxk12EqMqNmnsQ2+EhbGUwMsCZ1d7CcgF5i0uBgmjtqn
x8osQ5C//a6zEDXRBNV1NVa7ZgougcjUty42bjANRx+3xfMVifw5Ah+s383vd6C9
ICUXkJtsXkrqU3E/GH47cBoUx0EI9W5Y0bV0qKfPPgDoPKjIgB9QekuWEJbGGwOC
yOTKHtrol0mZL6TbQTcYMqpae+jKv6Iuk1TB//XgAIDobI4AtXeiD6Gpvs4DUEBy
SQCq98zrsTEBg21xfzeH77N7j7xQs9rgVsGoaf3HXiE79M3qVjs1HbD3om/m274/
sxT+Rb8Lv5Y59k09SwY8izzK8YVXpZprETwydFf2y8o/cxPlVoHfdsUlxsiujaLc
rLvTWvsKflwj0AJzi+enmJvZdc2W0FNXRysSDX0vCkOdwl6XiG3mg7R39A6a2BX4
reB3yjhIsqbpRELqEtN/ans3R0n8KylO0dL+cY9IiTR5Hl4hD9re7hP3g0kCQJPZ
mCwPyUGhGOd9LiXooOkyaE12Yadau2cQuiRzb9RX8Tu+QqoqJEjqrywEHmHL8q7y
MNv3PcQvdg2+lusV3z+IBmz6PDYvMZcEdSYpkU2qoP2WzN97g57VrNmtleVt60nC
OcSmn24hViX8UCrcLBLu6Tu5A/ohN5KtYxFjSdUE02wGpiJs63/ddpyTYNfkdeJD
I/sU4aMuGV6s1BM0vawQqDS9J8J90Tv6y7hrfShRCiNbagjKNkIdrory+jJIzLK3
esPb5EMwroSFl2DkqhJD+BXRehVPVz9o5zBuN/ZsFT4ON0uq3lca8aeuN5Sq1/f7
yT4JraQyfx2+rrTaum7loyPBbtEN9EIXcFFrfJiiVzkVso7bk6NvIfpQPTZqZU2o
kGxxJLyfBeLV/Wav29sItmKeZVChszLstCwML+EZgzYcwprR2nHVJRG302da3ZO2
ZsBOnbtwoqQuJb4Ugt1D1T6GzDaqmchzB+5IcFoA3uwME8HUVxsRrYvY9wlIG8KZ
3hlvN7LqiZoKDs77aGdTFUoKcXm2vNUEmnnP0BlX1VwdPLvE04UFm8ZsQ7mc1CLY
kRZulpYxvMCgJIBnTP84XBuTTJKDwNeSrmtGbQXX1JlETeWhSgYJdcYGTld6YFoS
GFABLvRa4SyMCpOvPYJ2uEtpUv78nCLzMRt1KO5FrC/kTurZvFlLjxfVflRa6FAq
68+kOU4iQMXmnpaMPkhjz3qtLxhURuhKjbud3MDqFdTamgQuf/Y9NxnYWvqvHzPD
b5yYktd5S+VKEwYFB1k9o57b7v5kVGywXyYEjbIu62vw01zNQdBYkpf3+Hul6K80
Itqj7AY2HM3ges5RuqC6zkSb01VINcikWGj+sGf2Vpa2w+4/K9obo7y6z90ofKlr
88Wnnj7Ae5k/zK83g4kL7Maqt2uqUePjDuH1k1Rsxx64qA00S9Xo4alKGbwKj2ke
1e7k5YvNoQjv5W65DgxXiRKVvE2zQReu2kETv6axoXl2MtlxBjaA3bvkxLH6STrI
AmoA6wFjyhxK9Shl3BP0L7tgqqcA3YMOfjsVHl0rECxhDEff7i85NwOpR9IM/iwD
aI1MLT7MZmTSs/Qh6z8390xyHXoEvYoQk4KACNQshh08PacgEHkE9COVihnqIH7G
X0C7ZVjXw4+PO+8pB+yN1kwvxs3Ih18pcDAOq+effDD5UijrzrctwgM03BMKooy0
5rLUcDdBZaHVqCAnVDmNNJAl515mQ19oT1axctiC0UFdaSMfPk8MVaCcPcM96XrI
x2ZLjqTfH1JT+eEmC8nWPbKwIaZ1kJWDNILbZK8qJ4Of/xBfToteI9WCHm3PigBJ
9Qpt6/Z9gkm/MUtp3rwkcOrLNlfkHuD5BO8r7AH+wzChBNfI6RTvMQ6I7eEgZ5q3
si4uMgclK0Msb+6P+QoQy1W40ygFonGkVQm/8oSWLqTWT7zMFtla/bvNtjoE6jMv
nACy4AppW97NZKB5/HxEdagv5iGMwl2KtiC9XlxggAazPhnaLQGYEc3q9YaXd5DT
OcoMOHrCZjZ4NrIlNtEWaZO3hIvVCl1zOfdB2tPY2rt1HCQl4/0LIe/1uBFUETKv
UUEZDuK2nVBNGAty8J3trajPHYMg3J9MKnFS01Qv0jFTX3A64qJBPdh61vpfTcH7
WuMd1TPOXvbgBJVfSymB/NXvIR5KeQD9QI1XA7e+F+S9u0hVoRLXR5TuOAMjjgQx
rZr5PRdTLcFvt+TlM02Ls3nsJgBPwcz1MUndbyITNSLGzJ2+9U6jvJDPh6GmWK21
lRMzjHplklXCoB/ATb10kq0eNljqRsEyFqvlNBphJyoI9RLcypIzrN3rpZCKqnxk
NcCgrHxvn6ixVVtdPtSsPrVaL5sZDTwEaCbwVsePvo3KLzu8v+aDC2+v63ezCBpE
KnFTXkIT2rJHWYRwunR4/yrFmDB3bHK1cTtZU78NBVR6wEuCVWcRZDzwVKXsYxZB
hRYjQ9oQtXfTvAwDRka9i+YvDXuHWdE10d11jMNhZlzmHjrZyJXpBuXq5Cy3/XNA
JS00JQUgd4iLt06bl5aGjbQ1aO2tzNRENagiABPa3XC6MxRaaynWahwciqUrvkFC
BL/D+xafFFJIxeKGytYXIt8iIW8uc8x4AupEJ7mTwUjCKJy1ivI9tl/Tm0ZxvInm
9s6cIGBo0VRz1uQAxJfSvHd/cEUehOM+RcCr5qK1BgeqEYiBhSYT9/CjRZDlqbUG
oIxWX6K0qQWwcuUdthIH/vnkGLXfPkRlKk5tcvMhKpDkOnOl/U+QlbaBSJzHOPFb
qHKYjjUlyZoM7HOYq6P7cs9MWhKd9YFalhMDnctWJ2nYitmG0KQqp8W6n2Wts8SS
9ayiUavKWAUvqpd78hnnICmriQHHgEJozIyQ9/mjyMN+oQtBHr5fOb0PAk8kSKLm
sWGRSQBWqi+7soX/E+s34MtSUo1+3xEtDtOREepzgbNUGIKD5p4w7oaZ0X7u9G1/
t9H+QEOmHmwnE1Q8aRxDPlpnLEElwYowCKujIAe1MmfzU3Gipv8872DkM407nT56
Qnw4Tm/k7LJ+1Fa7e7ANduttbNZQWmz3YiQuYqmj5BhKlpWtnR17EB2UfMj9R5Fv
u/DnBoZj+rzEm65mWgceq4dzPhTjHKBLrGBWyRetkAL0p+TcJ3aQL/ZwaBZQAKsp
bcivV85TRI0nrC3YkKxgtiLwFTotkOI4PTCkv1Saql0OX/ZJnLKusWSHkmg4BP8/
wpERxKPTktp5jzi7uXFadSI9GwDD9nR4EQipDhhGt4DRdn4+u5NGS4XQGkBDUJgm
2+bG5ygo3z4nNZS5W+ZGVzXV5TKEkrmlIKsrvbU6stflI5HVms1g+qNvdnZzSGwo
gh/vYHnN1Hk58HLncRW/lFpPKPxubttQu3x4ZoqBk6NqP+Uqrm0qGeAThwp+SpEe
HciSRNBR5QuZSj3gLDRd6mfHaVww2/2eJcmzXBxZR8N3eoiJ2OBXH7Dlzrt7kLYs
JoOWsIUfbeMUOzDuoHfHewgtfSBDjb+moLgPTS5qnb8tJnzUOQKj1Z+EBBqR8j93
Nu57xr6P2f7JU6YxxQhCFwycdwNooNmZstvAu0ud3ws3V21Eh/firo+tFxEqJAEB
bdNrCdygOIgKKWmQONp007iMVvVm0YSto3oZ4keturgiZMIOQ/Ait3BN+btJL+Xn
7b6dXB5T6zdt7QZVSeyOqSXhpE1O2Yj4Ekx6UCqz1tjtRew0unI0Tc56qXoOsMrz
GBUwJzWulHsirApHRIJXHcjE1d84sCfRG6b4oyCFOaEGYrRnSI+ycECaidDUwbAs
ZORS/AlVrZ0DOhTZvzFTiYKCUFzAU91IHEvNBbxPGA63fYfRTNHOZytr/hHjcv/Q
mJp0NvlrkStTmB2tBPQHg8SkA9p3Ru5aH1IUvAy8Mhk9pBtEN0Dro5eFGm1ScaEm
shZzg5LRtA49f5PLraVSoXMfIqRUlOwjXhgfe7j14bQzc34o0p8YVchBd4BpEuKo
ckJ+0E8pOgCEutLzxrq1t2RHQEuewezrrAtq2Rvf7nKzjqw0bHonMwwnrOcYQr1d
FsgT3F0T8EmlOpU57hh+Gtfiul6SQ9ATssTNf0gDTe3a5G7/096I/E/PI9Vw94xP
C/xa7mJfWKZ9W7TrINlNA6LnUaQcqW3aFyQ1SVBhWxweFF6o7wj4qFVLNEWJhVCj
J5CEEZsAWk+YHlFk03hxQbelckGEJMWda1nJiPY6DdynxAq9LTHAIz1dAzhXjkEX
Jh5DGY4qJJzNaOoVaoEuJHv/r9s5+5JTMK/EWmiSuxq8ewuVHC/K7DVOXqjkeLQy
Y/KF+MWg1Wdu8KrFbQuSgCis8RANxjmfzVZXMh2iko4KHFMtv61gVVLOEVHwqoB3
EjpIV+bNJxVi38gGlfZOQXumqmckch78Vo4zlWtehnIRCw42AJM8WSNSnEvbipqB
dZuayR5bWzTVfGCkQul7YFqBCCh4PTwTFzK2AFmF03hbSfe1jbu0GBTbRZ3ydLuU
D38QbBkSWBtrwifGZTEqXrwNxMUNOpseEw4XA48nNfjr2YG2Uhi1zxDB8cHjmVrR
Y48At2phn+UD56CPDStcLMZSGYcpx9/gAtYVe+5U3WjXtxmSebIrVuQQzheycawr
Ed86GjWBT8QkW0WW5UkqiA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LNqZ6+Q4ZLsYRY1nA7OuiePZ4QWFIxguxO5tPoJsvpjP+DPiK51X/2d9GDIOyl01
83wT2PFfHQTWWjHeuKUL1Q+9EkQjOQlMF+UcLd7B22QV7DQoLnIA1JWgZjiIHEhh
hso4Xzi61T8P9qAu44Ps+b7YceJcp+xKC1GilVwIfF7ReMDkZvO+0iJOVzY0tYY9
KCQzBeqyh1ObBz4EuhqRu116sDiXgD8rs66XoD/vkXJ5NbfxdB5GAbtTFTebPqwz
0ENFRy0Ig0ZkgsvosrdsaMgSEVhb8yIspk9JPVaBhmSbjHdmzb72pChMrNcjZKE4
4Jf772YPWSZCpuiywAaPtw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4288 )
`pragma protect data_block
Zt6BXotb4aHIpzM+rL2swX/dlcZf0Y8L5y6l277SRGQQtIAkS6Wm7C/bK3ZfelOT
q6i17bd8W7a4MO5N6IMqk1RTaS2NJKY1Z6noAGeWdXmUwBsssX78NOYYHivg7JWQ
B5+1dR/g54ZgmpjE4qi3Wi+9JewsHA+UAqkB1dmq8cSf7vkyAmQJZNQNyUxY2uNS
W2yk/ESA5w5cvfHkJ++NTBNoQShOd2khcxUHtXoVweV/aBQa/+94vzG6V9gOhL0I
08Rlv2eW0Yiy3f3ZS1hqWwacLrvIHBrB32/KKJiHHbiIMdefaNt3KDi+vaJ/C7Jh
vW0NNcww7SU/oQJmXR4tRK3RPfa177qwblBORPuNjvRV9vh7w0jTYVgXscHqEElV
Z/zv2O6pODE3ZkNt4rrc1xYhNQV85taji90+qQREje3BjTycrliKGbLxuIrDoKsM
ck/1JfL8C+rnRXcV/6wHaJWrPtPg5HL/qic5ihaLesYITZ5/wgYfEnzdRa7NcKBm
txmbN4llGVuruS8GPGiIehkDryBa9dGhOgoRJAfjfcNgOVI8s1Rs4xSnwG5k3Lzj
422CzHITDh4pH8h55EObtBkhWjz21Y2oLB5UGrBjW4zvf43AxsCtb8UrY6/VYNkE
WZZDbZdklGUkKpBUt8PEMm3LKs3hQ4dtmfj8yQUraS29g6LWbvPKkaxY1vXb7Ldp
8IYlLILdHTZKGVlpp3UV02ch8Vd0/RdrOVQLvw0aVDq/YIroZPNNWCNGAADIbjXu
h1O5RVlGtzCE1gwsD/5/4ePzZTseb7iInOYmKW69NwrluAD2XpxsZUIogVXx0oLh
qDWFHWMhEVFhicmiPLN+/KVoZtD9fmc7VgHYy+aM5UezRKv2bze6s3aKaHrNGrxC
E/TDWbwmdpzOBA0uX5H8pk7gleTGO+ZkWrxMOdeUnE7ee5HqzOo6NuhNbY0m3Qrm
GqX2qAFjQibO28PEN4gU/z2D/BgTlWIe7KVt3F7lGEmB32sx/RauonwTGXJ9l0uP
syil2sjyCwevWy8YXF9THqJ9w2Tsy2sBUj0VLSt31cF0gqkjYyU3dwHPHDPAEuVG
Pc7obS0+xgN8zB6lsU0Iu4UwHcno/yUTTps9b+QYzli3EoIeqzQIawxXiEI9/U6E
tLGlsKcJfj4BK/cCGaSXFDFkvrL+JdgkzI9ZEjNfGGUhH7/5BLjn8JgC5OJ3FKYv
Kvz43P1aKcDMPA7btoA8GZ99qTy3uqF6zu56Kg71DSk+UysDMzFUk8x7OChD2xlC
idm0L1/Kg+/RALQr5525/fiz2elj05OkUTIsAm8sq28I4v6tWUovclR5UYIeS4V7
T3hvdcZw8rWe0KECmkdixNyqGU8k/D6R8Rhf0r2FJLYqIZUNueqgIQ55KTL9TddE
aPfaNpJOjufge0sCfKVQxAHcG0BJUfWFUsi0xP4wTtVh9XhfgzoZDguYHRwXuHZ3
2M+0HVEQWQyoNgOyPBGaD48K7lCVGGFBvBKgTp1TTr6vTCjYBKGG/NrevSzCUrhu
kaN1o0HpAE+gnb1dmaYACwp8DqKkOYNebJGRtsSeTuGTMxy9h4foc3zXFunNJyJC
N3qeKnFmFYlB/0E08mrowiGlYjNZnN0yNPM5J+XTH8s31STKbDnlEIeXqyz66yEu
KocXd1mxZQdx6xLTBTBwi8eWvqNYYJCkxh/ragq8EV/x8Vuesi4SizA57RaYtQBZ
ZPa2CNuwFfDWX4z5m1wBWI+sbpRCvZtj7MmAzi+Xcth769BBnVyxDATpWlJ1keQ1
XXRg1rE5RG9QM8+JV/pki/qDDjxyfil6uNdVtklkzvmKoTFdmf+G8CdJgK98me3t
ZVNoWm3L2PMyZQ9+fUEA0icbcMFSNPs94mQH5S0CskgwIJt+V+cEEB2uInsKkUOZ
s20W64oT8Mf6we9HTMgYUOUSxzOojQNMsHcWNmRIkoi6TRwtKrM2Im8e0QQWsbsf
oVIplxJjragHEXr1emrx/FPa6h2GqbEzuqaSi6UKpYtg4EovESVCS1qjtcGolkDr
/UIjwK8k7QLl1nMd+5PeM6P+Itiks6z0dwAlOPf87j9dIrx/L5qmlRgiL9TfFjT6
jurqaXPNp1NduTStjXIYWKElG6wCWs8AZPTlcpy5pYmQ+tzp7zwx2iFF2zk+nGk5
qDa3RnN3f8wGDpy/AYiD94PkKtMoMAB5oGgmRDBf305GmBvyeOl8j2EGtcY7Vtwg
vOYpI7hu/snXZLQhDbfty8ln5HwRy+Yo4PqOsm6T4gVL4GWbwb2WzWmFYAoohfGJ
at4YQiOSNG1AqmbRIEJRPI8E0EnGDnqMGYFtp5vgaCUXdlwrkKKJB55Iu5gRx8Qz
LPb0tjTU2WGBof2aCvdWba80DG14WfDjVELPDoa329GZWGFMQVrvBSOgKs6qVZDB
mE624TCT2NMVqv7p4Cks6cdQfT61BJvCbuGA/xeVQrdT8E/8FgdLokN9gWNzyJSF
d7QlhtJ5G3zmvYsOvnI0Bfn0QrfrgdDZcfbOShF9Qi9IHKv8IwzEIVmqsvI75Huc
80FKWgdyZh0OBNC5dk3EfBk05vqHssknzQbtJzLg1hKQkoqKp+hgcmFUOwziWWf5
3Onw+ttmwlSe5sRdORypBqUjVGNqgZnU1I5oc6ejlHdLzbj4PU/giQqs13TYRhoR
myk9ezL17X6umwxgRTC0Xxjkst09KjI6UT6sMya9LNrFqgIkzyxAlLl9aF9i5gyl
AwB25gvOoIqOJDtNOyBNNAWwZ7yXb8I0BxccJ3VvMgJtR4qWWDtJQ7qTB60qgmai
2F5O9uXYgf5/XGWNvsD2zwQJKsir4dELZ86a2v9EA3bsdXxxT/LjuPYnGOK2YL+h
nnIJD0ChH23vBtJKfzNmOfaQZg9E+T3lyHC8QP3FLC3mo2CdQBPDNy94axZpVitE
TrZozbtQINvtPhOv77HiWjOivSDrHagX4eU71W6oAlgi1B2tkiN70E3UGqXF8pXi
CyFdEOcx30twACXtZLsXcIKcPW7gCqIy6rFiPs5UD5jsEFGcFbbo4kkAVyLXLi6R
FOUpIvXbAvnca3fHGsBudr9Cjg0+2BvJJuXWDXE83hJFgu/JF4+FUGS6Nyr77v+Q
N10lCZUXgB7/ADt2+LuxBRfVYEpXxSm5UyqSy3fmrlqAhELYWntI1irim2ifmxme
DL9EK+6mo6NEJVWK5E/4qr5Vvx/zIEVkbEfTw7BP23SArm+l4VD3IBFX/gSbb5z0
rd57swxV5Os/z2fti9GcRF2Nt8TC+lgs9xdogX8B1OsOkByavDNXLA6dKPmGshss
IkI7rsHOswYzJ5sqByGhRBoEL7u+oJLWu/akOhZubDa1Ed+ariwtrRHVs5Wo8jxa
qtWQD5fy5oC4+gM8NUy5NdiMxijVpnP+UBenbLqynqV43UqGk12JXobNF7NRb0+E
U+K8amGEKwQxFFoQOfw3gwxETl+d8m2f4FQFsgQu71jatLDXxllo4L7nzcydwZ4/
ob+K9dcF0ip6AKlwbqm7oOPEWA6iqJmty9wAppm8U87xnqbTctUNJIjkRgCF6Niy
zSixoE9OtBeaby43gMbPOUyqDbJibZEJU/fCMnrrLW/8Pue8tAIRgvrgw9XaeIIM
68whCFZuRlYR8uNaasS4GlOvhUPpOhzVrdDbXKOaKb1WVKlJo9OEQnp6cwB3nWUH
QmzpYZ4bTTTk/Zu2DTUJoTeDbOaObC867EeYnpTLQdUfDS9m3DEiVfoWha8dRXv5
dZJN4W92BpnsZVthroyu39nCzYKDYZHvIQzj3jitnqRUPIsPB57bmBU23I0NzgHG
G2R9J/99pVjG9ykv9NokbmwD0PmbicTBwUYDdYb8rtVPeLm3VKEx73dal1jQb8eo
V3mzzZhVM/ZXdRV1FUoam0EmkQMzc62BvfVlRxPugzBA/rBzOtaEX3S1vq3LiEzc
eZceJSdFOjRkdCSDv0uw5EM499WgRz0oKM7H0mNJXDR/163EnnUgtkwnMxS3v9T0
GSCi8cXvfXyAW9dC21QPn4ixOk+5PkaQGlb/fid+Lqmv4sqLCjcpiPdosUBZ71ly
Ih+6qVZDZNMzZUJNMssGn3lK9Jk/ZeB1fnI+Ciw3G+nbhtLfFci1n5X4T/Yg33HH
T+UHdhhm5wduOY3wdFgwrc1nBo/dT7Zejc8VUvm+d4bzf+J8TTAVVG3807hsAyCO
16ALAb6WprdYYuESFeUKXv8cguhNQH050lgWU1NfuY5IEEy3VxEmIuSBmuOci/D8
uTTP0v36QjaH0TgsQafClQ7svbj0QEXw4ucKFueQyZMvKJ2P7wM29Lr2Kn6BNc99
uY+guP115a1XbeqmeqmWnkDCKgHkElBscGHoeH5oqdXKMIQn7ee1d+tU6Hvhdnvc
5vX+dZL8OY2oWJkPvB2h63daBjut170u8nEJ2HSDzd3RDLJE/ZDB990791Zv4Trd
bHgB8vtdWEaMCy/Zccku5KdhUM5upagTdMMARM6HcGWxP19+jQrW3QQ20Qi9zquX
UOOpyfekrGyDXL211rCm3WLzkWJK8vGrhVHnjFkXTbI4Fma5OdOe1+fSqFbGxRHy
CIztR5ERKzQRHAN9tCrYNp78SJV8O/sSOoLGv9FAE866VKnm9tiVzNv/cPKWrGll
7AbxW9wbpkLYVwU+TWRsByqeavZ60zwQVYxCXn9NZwIXWSH8DDY5m/O2FSgaC3Xb
yfdZCqZTHMt58luVUnVbQrsnGd/loLB9IXgRPV2NtVj+qQd8MWFotQCsqi+7m18h
Zk7jg4mlthnUqYnRpDpciL7kT0Is8pWRu03FKDUzXicoWIOt1oh/sElQdv0k6sRZ
EnmqXJQtoSoBAcLXOJ0WjOry5LdZMXHifoKa1RwCo38MZj7CM6R5AHhzlj2XLq02
ffipFf9Mxl/6irBCPlMTFqGFASXbxguavwL6Gu5tneDTzGkXxly5UptBWHEWpXUn
8lNtH1xG7bx6HZ0bNUo5HpBJrwK+6rEJikptm1fRLqj9sLzRYVW7Mt4DPa0w2U9E
+j1v0jlMR3pavTprR6FqMiiHmY9gaGYlP4knAtFXOm1X37cmW+K7qL0YzF8lqOtv
pIlgnNjsDXemz3dBJJ55B6d/FMj1CukvjsCsPmydxY33/6rgvOqVkkXXkLxGECuR
n9G7ie8XVJOSiKYRDmKJ5BlJq4uFFC/l86AITyxhni8tvguIPu4vdYZ0S/td+7Jk
MRoq/Z6pxpsy8iRfkMkzU2gVA2QVvpRfyXEcY9kSLEio0IWDJWkMsqpv+2bKtD0V
NGPLNVxnPskp+G2xJTUmX8QbwoS9ZYykm56vIUdZFncI1kHWinEy9rSwA2p/XpYq
PsQjGB306jmwCDckvUSwiuHiDrNnBwLb+/b4O1HUf3jOZTMZve8crHNj86D5mYNm
34O+6ZkRyl/iMy5v9FFO54KuBUEI4o0sI9tPDaar2NLZOqYG0pEUYAM5jIlsqdNY
3iVhNYaV5J5B8NAxusP/OgxvYguWMMRsNfPaOAqtDo4bmSuWD7G3rJaaEqp/Kh2i
VgaOLTn5ll+4HB29wIeQaZ+gFWLWka/RqGGBJ6FDeuQr4J8qiFyOQZ3SrjabQwc8
iyyaJJnNt45TGNuG9rJ7N1pjDF21ZJ7vmrgecneI9l8OUrhIsHpozFx4zwAwmVl8
bRoBOAabFLDkm2N/8E1bIA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nZeRp+OHgCHI/4FXHqsbt7nEBwkaXeymMS3dmr8pBdQW8VtBZUzKeCurBtuZbr1I
f+Uo6vPaNm0r0Y7lp40rD0xs6E2sa34vYev9V44VL776dqayxG9i8OuMvjw0llwN
EmLQ6kT2l9F5ZYbRhwX1tcuipwHneaMcAmmLiuUrWK6O5xtFCAwVCutvvxASixrc
OH3S0zNUi4JZPMl/FAtDUCNJbzERzZ3z9YbiE7ib5H0jaQsAnnwlWNpY/ixANCLg
NqTp5UFa/WE4J7QxAlfMK43lKWXuOhZ4OuZu07KTF0YXLm132WiC2e3/6gPPCEOH
QOaUoOuWDP7wFVTGBmSb7g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
/rtDJsOK5wvRrmOlS1Y2Ax/DIal0rCs1U4CIXAseUGjZu/eGurJuCRMEN29wub69
mXoSgmLvkiQSvWhan6kG6w+fbavsAUeQ0IC0FRGhC9EAEHWY6oFJoMBD68XNqh14
tyQ+08KrLqoBmtJt8cQpxUGAm6mwYKMM6yg0isyhfAmEcfloS15ljfyztIJURPSi
DABP9xTxLYV5jNiYt69k4GCbBOPwoxxQYwSbJhRgZqRTxAfEKmh/EMjUyuyxUDRY
Ta7B0yNTsQEgoOl63FU9m6RqE18LlvebhNp4VZ7OmiLEgJ9UMM8KtEvHdVy2ApGR
jf0ZAZ5oZLgY7I1xt+RmMb2iaotpo+Bg+hfJ7TpPxBPLhwEQq/CkrRuMSgttb4nS
iR3jxDaTKXfKYV0qjtYOfdtJAiT+DW5FV7njHrTU8sV4sWJ9UF0CNyF8x85Hu2rz
pArEdZpKGkVpj6j88qi8r98l7TpLjB6YDI23JQL4NAAOuS05HKCCF8DltN7wHwjt
YUa/7a+GIn5ehmcVOe6UZFybT9dGbeCJNTJmSinLds5bijQxpfZYat1Jth9R5cG6
pALaIY5La5fM0PXf8kTPnONftAIj0/DHR1JlHEfoFvda1RKhn0gG/wCnaezVNApb
oJS7ioNBvZRcTydSJ6jXMV71fqe3VgHtTJAt+yG/AdmRiKEtSXYBCXPllEfpu63n
ESiPPW7Umd/FO2f2l+Q0vaGSj46HquERbp1G0DJile4fFUBfNRveNPexQ/+PuFPI
WWuADnP4e5E34lxhyD1LqOEhYXtdphZK1bJdcK1Udb1Ktj3644V0n8h6iNqNG81x
MIbPSXq/KaCy6aKLOhVUE3C4+KGBiQJaOFlaJtbIa3netAJE9IPfMC4U18AsDrOR
cI7aUJIsY3V+qw/E3keWGkKyXkvIpiStlLAzd4LqndMxjkMP5Fgqj1CDS8B5IdSG
G5OyQLAvyXtcuPYBD3PTlsXwczFCB4Rvv7E25/Lq/qPbtU7emHcR9F2UfBMi5jXg
oj4j2XonlbG8ueoeI2fL7QTV2X/C67lxb2qnkolzKW5NK2yUojgqQLCYadbabwCa
2F5f6o80P/YjCPxAj7YxJOi1m/JFxRFptk5k2oA3gRd3Q8VdeGyKbYnoq1PxoZs6
muI2HQaMmdrqpHPAgrepNUS/4ZLopIICSo5/T5/IpyzagkKN/+Zt1eUK6NEj/73q
mGxLtdk1erCfeyhKYLDtWXdTKkqvoegiwsfoDai4v+ZL8swxFLdZKL1SQ2B0ONsY
VZAUjwmBNrXjFPkH4n1PIuKPPHqtswMzYPFF+FXrSXNW+miz8xpwjzKy4aYosoZI
1OuRVGRmPnSO6qQVnlZwoZbKN0q1Z/RyL0rUpkqRIU5rrfAaAvsOMJ8fkCJPNNu4
cLduxsEP9vBKFnMKHnW/mz/bn7ixUB8ICN6WJpXuhajLpHnu0xsDBgCbz6TOfu38
0Ce/A+mBTmyiPSVc8FjqgI2gmip5ng2eohicW2Pm9tjxaVdgitzQ3v1yYQmUT7mD
Ei4cVftTWBv9dQFweidLfre7v8zHg6rdT3paQyQgq685XmGgA3lxm2cwj9wuj1hP
N1nCeEn0mcTErDCaWmNQdS66VN0Jc2xYQG0sUbvL3VlK//V7lED23/wXHT6gTPKU
ZamckqhGUWAY9rn2RVkeZINv0q5dIe7QWLf7nrm+Z6xUMD9fTOCEHQv6SOm9joNw
2WKrcrtcgdQGPbwVgZ0VkUnGxwj8woEtIQwXY445S+I+oSfawrn9SEaeAW+0n2pM
6usm+5/fI4914lTVLKp0fh5Ghd+ydeupE7dHUScWPotz7ymi8Qf949VSQYE4hQlS
TYIhsWYjoS4ID31pDqmIS8DJCbUpG84kvhHJ3lK5VKl5nUt0DiRcRZF4rhR254N8
tssSE+rgeJn1dUs0RBGJll0b8FN2u9/dwlPEP72jv0gIRMIvyZPYHnSE0Hn91a0k
CwAbbqg3aCCyTyPczqB6bagnWTHcWaiRTABtcPjHD98SSkxVdO8TYRiZZHm13Ov4
HYg2LlgrryvtJlnBVKRqQs1lvV0y+qLMe8W+WA2IGL8vsMgNrTxxMeRdUKwYnOnW
OYb+nwu6baDi/47nleOrEg0UwQqM8+3vyPcoG7vqehz/lQU6UrM6wVA+umcRvU3n
HZPelAodTi4VWK9jrQFU202lIgf6T3Alm9owDrjtS2jvf7kItKEOueK9gifeRr5L
ORc+ZC2hLbta6x4W5zrqIF03C9QJWy018Ujs7wZFOvSjM3ImCCh/RyGdZCJP9Om8
WZhUz0xmJUGW+G7kPmXWctthCHMdYAByjv35RBvy2HK64I0LnjnlEm2Cn3dU11Gi
kfbRmbHefRW94mhtc4eNCty3kMElPv0+lABiqIXOxG/cRdzTSDA9iKYqqJnnuDtS
t5EcSvtNjKbi8binZvWr2aOQGajKimnr/XoMUZE5A833zGzvFXcPfTJHNGTzHW5e
Uy+p3Hz7XXXZ1c/WD5xD5bx3pwCymVHi0VhzeizEVqi3Mh8QurdOohTvy90VoQTQ
ZwQzmnVt3Zxc7pTxbeeh7xs7lQphHUASsghlmqNiE2EIyGAE+h5yU36zT3MdGVvB
rr6V4EZOXfd48O2U+XqRfhrDTZ3Nkx/uU9hz6GbhQi9m1pj+mB8gWZHYeplv9fw1
qDEu6xbbw6FpkpAV1TAnCLH6nrRfebJ2JBUBSygzireVLFz5Yf79cuuMe1M6kjLG
dbdPrL8Bp4+eg0PmBVNQ7fZ8QTiTFqe4Qv1jHcRb57DkNdLSk9W+xGsSS7tXkSk0
PlJUFfkd1TBxLLJL2OOA6ypUNHAFHK9e3iqNBEVthrkHwzIeiZyUZIaF2m628Wh+
VVfsRVylzEZCjv0RfqKObZDQPIp3HH5Nz/gjhHnKKlxnxwbhawj0/8bvkOqxf9lm
TZkJ+NJwLsCxrXaucbHcP/hukzVTObsZ8yyfbeD+E80etem9odn0/crrWlwp7cZd
AQVXmU11JH/YqppfodWaLobklGkZFEaYOQBBJjvQ4jLZhDajPeFOE/OsTY4tycPd
//ch7h9Dcm0BLII0o3wQpiOc8Cf5UdtdLoNEZwfepUdEg9aymmAaUskYwxC0yJkA
VH7BjdgIFYRPfdZmGPhLQRa6xAJaCQMGAjrpYnIyG7XlfGSGPvqV0OzzoowuxZQL
WuwibIyx/5mL8ycJj8kCYJTHES/InwIvMRLk0clxK8BFmN8MHmqlnMBlSvmQvCBr
DyZxzZ2YgTIXUZejo+ob6vgA/juvhK8v3BJKaM2FzhtwmIhP2JJr39grlg9bbJ8f
L8+IXJCi85ZFpyGNv7+DWG8efF6uNtsM1I+bk4vPqShXbwx8InvDglcegoLw67MG
N2Mvb5nIO803pfW795wiwhx06FwDKuSJb+6P0wIhpCovRheT4PlLEG/ZiTW0Pp0n
6bHpnjhn86dh42UIGiCSaBRjQqkN6egE18RW1nIGeA8E7sU6DssrGCSOz4LvqgHu
7crttn8lz59C63fW44tJlBZmd6FtiSAh7OGQbCI9u7y0OXyzRPwTnHn40ZdLC4ju
CdLOdlFbg/OHG3FYNHCvaStn98AS8e7cLfSj288fnFbQAtc7YutOdh4kpjuMpjgM
EnUyN7pCuiP6cabuNS6tDfgQK6bmqbWyqSmmdkLH1gSRT8/ICGXGiiE4Jgizqz6p
iIEb6WKmMOVwQrACYJV7u/ZNXiEUTNtT03d/d0tbH8/8SB2XzLp6H+oOhFyykLBh
vuf4TbI4pKJddUnqWxCzHEIh6aJlE9YIPLMi4DdsvHfjkj1g/LeDuIM+9WvddwZ4
d9gkTyt3fbCr2Jc6q7WwgFRg5MdhCuhyPPsyghFQE2Iayi/Rb875IO+sDhWs/iP/
a6LBR4z6PApHpDEqmj0IofcQcJe+r0+63QqhwbHhQ0cV8e9jf7uYcdAf2gHrFw03
rbvmjsotdwh0mbl9gTmBauLSGr0KYJbKCqHGgyhkKygwEw6GbMmuWsz6hLE0ae7G
B99jcuE31Bll6JAv6gpj0VDXOcIMJDqSnOcQm6Z2c+fp7LIHW7xdsEPLGVGP9Kyr
CxCCbX+Zwnh++c4kXZ3pbj2QiiTAGRZ4O4ap2myt6xBTNol1MYal//a+iohH+YnV
Daf3fu2gFq2y6l3Ucb/HGeP3kvzZhZ2I0+8OTfkuNGzQF7B8DSDw32YSNBb0pGcp
M1old3GP0Yamp6pqVeQ9xOTsDtN88rPKZjslWPi5Qx2pcwOFIdZLD1oY4Xejw0I+
iqXpTQUMrEEGLd5d/BQbtWrhynay9vvrS3A3WPMb72MF8wULRmEFrTR6bTVKFYgO
4/Ydmw3wO8ukvsYJHkSdIrOpoLHMMxwkB7o40vBvNNkqzBRXoG4fyB2rGtEFvtA7
SXgCt4YxfEDu/IOwhQsBGqLQGsEqu3SOXitX7aKvqy9MoTbFSkjbL/HKFTdT2hwD
+CqKTrMzRXfzCwqxrauaG0mK13uu1cpgkr+nIYdsbqkSZSnkGPAHnggzGTxVbK8Z
7k6nFzXD1+xDiJ3+UsQ33AhdtQ06sYI+scWNfuARDy8O47RrhzUldOJjrrVTzjfA
R9SW1MsFxcrb6udYYqIO/Ea26XpDk5YWfsNX3aakJEuj0ZvMCLo/4JD3gjX+IqBL
yK7pW+fOYwvadnO+bgydxNY/Bggx2w/0GUW3AGXaLlvWEbW3YidCqgEsulfTF47J
kIFwGnnvPUmBhby99vjRYBKO+Qes1uEdV7gaqXSebPdnPH5yy5KCJ+bBM6T/pdv6
9s7sR6uS/7DRohYD145jXgrl+1oMbNbAtG/DdCsYhljh6SbU1zGAbFv9wO0ZOrIT
hlA+rvS/t7vmvLyt64L/csQ0eQDmYV8VwmOhGLvPqPEdtO5VPvvgM7DAESAkiRCO
BGYh1qTyHnL+w/29Oq8NAl0vbbYAxzEfhXT+WIvLrAl/O3Ba/9M6UFOviToKOPB7
duvoQHWD/EhTUfoeX7eQj6FeR+OFAAWWyqpH5J1g2ZhyFXNAAlHnQiYXjGFsJ6+/
4vj3IvB078DtZfVXMFoQkAW3VMK2/wMM9ql8GIz/QFI0EA354L8oPe+xDg+I5FC9
1IlShVOJzGqAxhcX/Pl1KGIX5XJoqE+Zl15zySAeVws=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FGx19uN4KiSfc6GA5MRfMh5h0soJcVN2tGDhas9rupbnHS1HSEiU5FsEZx7VKlpL
DVlQ+HqxcuuJUf0qckXVzABR0vWdwnSA53M4LvGVDkn8FW+CHs2XvhHm0TEf9PSj
YJr0gIAHCi59Zpfa2bEcqaFEFryu6Lpq9IiQNJDqY5TUOd0cfhl+1r72sSFOyShp
AjyUJ4+d4fcBDmcTe5CESZHszQTToj7L8lqQOeQku1iYNO/0xn6+oyihULeXLmN+
soCDuQPVjKRgtvBYC2ncHIwIT8GWtq4UsCkbxUqdj63PJhA01cL0+eWqx3U0XRCp
dbTxD/NU/FPGOiJS/GDKvg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6880 )
`pragma protect data_block
Ey4aGeHjtzQ4IA7fb47eYeCTJJWTbBwOlvf3oe23Y/yXepKsHxGUKhNviyP+Xjf6
DeEh8wPeTUvP6hvk4K9iddsh+Ntg9VvpQ4WjDld6sUVRf3YKbrIDTGb4y+ZN6dty
pWB/UHU+YULrxUc4ScyN4ocB64TCURR3+Q+9iG8rPH/x3Mtxlq6GQHfA+BIIBg7S
vSy8RuFRbpjQMz3cz19U1yNy+f3GQJDtsEoCzDNq9n8ytqUAoQFVpL07ZhgjeOse
e8LmQsY+aybQHJkG+IXLuqe0H5lNhpJjtBbpXJLAYgLGK5OQQTZcCTdzzpWynAol
CT4V2S98J+aRiGFWk1FThsrHRDybMW1w5PPho6uxUeNuI+jZ43G88l7JT92GeZSy
OSBi+G18PSDLxjKxttk1mR8ey6CMNL50XcQX14Xnu4ko1DsVPPEUoLlXOawnE0Dd
zqe98NUUc655uAIJmEuHLMdZCAtWgrRMvPH6IXsK5hrIpzbYiaBGd0RzQWpSTUb9
GXqN9hxTdx7w7OmQTHuGZBKpJdEd2DttR+0rJzTDLlBZdwQ0itq9R9ZSRmszVqlk
69Xh4IThvAJRZICtT89Xs361/4mM4QzTKtP0jkLrO+YcSy/rF/7Ylp+c9XB6zV5e
V/JkECMRsZG+Bn78Gfpaa+IgLUcunGaR3KOsg0CS4LNOqKq7izgtS9OL5UY71+DC
/ZnYwNDOu+dRgh1YeEu29dKvq5RgYYMEHJAKBidlokPLUmkr9ALtsr2IljM5xDvX
Oo0yGGPC49Z7/ECI+4avSOs49t7T9ucUKt1EMJQ3btM9H8tPPui0De1U76YzDV+s
osKspO7weaKHpCm5x/bSJbLRfUI04XYpdN0I+NykvAr/gZ0usFdH3MYyzvqR/Lxt
h65srcTxggOaxkWvqEY3LsFY0Bf+q8GkJ49JTshuoLUx+FWckvHwCkKS+qYqsoJO
BuPAC1TQAkERy9UVfh4djVEufB5p+JgFOmGLFu22PRahn6lh0vyjs1Yab2QLGNY4
04bg06WDBsSin26RgAigSaa24WDwOvDtcEb5g8e+I0hVZCNpil9Fz/PIuP30eQPY
JAZ0yLH1pdyioL9MR5G3Vs9XaFtY18ioQcrm0u68LTQf2j/4M0RSSHihqWOfdKfl
32u41H2yzrDMUhoE9Cktnr/3oUq/nK1N0PS2ox8E2XPvYlTDxBiY5npIRrM9E8Q2
vm3EwnKaabVsvIDf5HA4jORzZHSTRhCckkuhPXFCI0LNuEqGUzyVdA7Kd9BDjdHN
gQlUx1m2rpdzXWdNima2T7Kb7noTRgZzvk6H4f6KLOPNLA/XqtSQQjxy2Axz18Ci
LcWVS0brIkA5dYqsFq6oR65SSUvrFFhfFBXpW8zcCP2TX75wvd4YDQTpdWdHyZOV
lpKJkJ36lhWaou2G2beI6f/34SA1YDlBjbK4RfDDa6hl2QTtMWyS87nenoeAZV3P
AtwgOAxGK5NSANImTS3WrggW3uR8+EtN0WfH9MCp28YLiYsOffx9rPhzbWn65MV1
EIo6QKPWWOrbn+4Xlg6zur3N60gjghW3vCSxlQj5Q2iRw3VCD+U0L9rggHqxQGWd
VsY/848rvJYrMGfHpJy0mXtdUKav9qySYwhatybxGF+4diqbrU0wFtnldbo/EvCH
sQF0e2NRQF5KkfzVO0qNm/d/eAkmwrOZFkzaNCm4DTrwPX6RpCMNIvt+yiuO1DiA
5np/Qb/kNOGenxUA/AleuSxFnxaY9c6q/IMLZ9+ajTQVhYaqWSRaW+j1XTqGu9fp
dUyXi/7l8QrwkQKblSdLY8UEalWcqz7x3vu/6L4tYq7AyPpumLWb1ULKTlCZORGi
5DEVFt5UBT6NPMTrCi1HrtNwIwce8ijKxJS0a7e9h4WKJ4+rFcwv3I6oN8l1XB44
jaf/rMyAr+Trm9FoH594nQT7cv05ReXiGXYQOLRsuonutxKJIgRQnDhXQjCpS5Fm
eX+ccO0b/Vn2x6pE1gWgEdzJdW6bnMtSP0O4WCFQtp9MxkILDy+yAQwrJMrB3/My
g7aRq5NQ10mfL3BFZAHRsSi0RmLD7J96qT1IrXJEWzIfS+ZIUKHyJON5XJXYNZpO
Sr4/WITDGCZCd7x+udJEsnltWbJ7bsXyZAj95Nywnph5xDBgnlUWeeEdHRpEDxmM
XGlbwQUUHYcnxRB10OrfZ6SHOz6EAVU4MtS2uQxcfGweVRyWT/HDQM+S6hPiod1y
1nd2XClwxz4Qw3yRJQjW3UywUjOaZcQpSyo22d6hoI3U7Kcm2k4pk1obKtZTAdFy
suyQW+VUotcqaJ3jhQOM5jcolib+C9GVbaqCcvbEgr6mnPlgB1ehf1IyG8MQrsTE
j4p8hpWB1QdkS/47q8/WnIgUO16I4sGoHcRdQxqCPjXBG0Jl3pkucHURf3fpu+6K
ActdcG+9BXwE0NIU1UC0xAjNgXlGKQJeL9EWHWpnL1rkXWxRv5cII3c+sHJ0G7XI
vSg/XNhP7O26qPoAfml/PzQt/DUBaqZBUVMHBeETuogM2pV5dRpxK/UzRAi/4cqa
LKLXII9OMqr0W4V4bwSZc8/ndmF7gTAVamwS/elTPgI48iJx9rKcbqw91h+eHg4U
GjusquzBqe68vJDAE7agf2t/bgOIIjmTuEFUxiFagpTOwQuKdqHnMf1hXYf5faxo
5O2TixJS7j+lW3MrljanJQeTt07Err8GWql+MyXZN0LrjaZFGO/QrVd1i/pScYYY
KPVs/Te6KaH2qqSkZdkaTEAoyWAWlLIJf57cw0t8GI6vlL+G6e8JIp5e/6IiBdlD
mM1cL3qAdI5Ku98p9ws9DHrW+V2qLJMyMIxC6RAprjaE0hwHx4kU4rnh3RxbICYX
DaQNe1txQj6SJXbclVBHFHJO67UIfbnqOlUkjnZJKLwjAqspPlmTup87Cc+7Aye1
KGBUAjb/nL1ojwIOiEg+sd35O2i19vfGRit178GIOy+miQoOX7j9cfBcoQoFks61
SOL4oJnZ4fd1H6y5XPEjKRvEm+xFHY7w/WXrxAmmjHEPgRjNtAMjUVLqzppPt3nm
39o4NBC7o+yYa3KqrtxJoy200GX/CTBf4wutNnmNxpw4zj0ylLocvq/oo5WoZlAt
GmUmzIsFEVfA/UfBhatVlnTb5LPYnLmcfiCb+z75HIIskgPr3UShobgGnL2g+eIU
VzYNxtmkJE/x3UqOzalqEot85HiiTbU562nMqMKKlhHai24ZWm3vYth9NhEjLoVh
tthDnV92oULkoJIUJwoSGRuzEpT+BGyd4lfoKshcVoWLfb1r9nHypd772uC6K46/
DNQGczR/Wky9eplKS7fE9dmr1YhrTzv4oy1MQzGHEm21OPpRgW7L1ZRBeYsFyuVJ
V0Cb7+7Qaiy/5Mbd2jL/BoLFxYAkiB6O/ModVL6UbaAvwu+w4IS4n3V+n2v5vrFS
+q6XvGknCPaUO7AxOQZcar718NlUD3cffjQyyF2OEhL1my9LuebIpi6uteWBcrB6
3by49J2apY0hp4OtpU3r5/k12nfJeJyMQORk0MZBcrzf0hcuaDiH0T+MCOUE277j
ald0jV9gPO1qZVwcNz3FjnufhtbBHEwm/L71ae/UZPZtzkIXxjn5iLlcfVZvT8IQ
cdkeIofLby+9FYmzrepfiB97IkMXANbXQLmwODJB1oDDkxqBq4mXsT2pByI/W196
S/+sXubOJsSIYX090pC6YP8zRu/milq7aiEKnKEt4GOoN/i+amLZhxp0ZrhAlWrZ
8GAfZBPAD4u9xHPNA9XCf4VQ90zAVJNrIzJddEvIzkH7liEWg0SxpQ0RShuOe7HH
QwSdLf5t0q+61gvwuwNA6rXekCO3N2sa+R8llNkzNZLMEDSA9wQOl7sGXK2Ah1S/
GWaANHhHHAU4zLuYOInNJVZY+899EsaD4072YTnUC0EtXi9hR/8Qjf+akW1C1zR3
gTAbi2847r9e7lUeH5S1ksRMz+eGRiURmnT76KUhqJAuSbB06pitk5qpqUySGhER
/1jKk4EVWlTeF6ObrBFsjo+UcxZUZk+ZgGUlFrgwrKCtozYgXUTn8XlTR/wOXktF
zdhQo6bQj2Mxn6rT/eV6GMamxEkm2w2ehyRScb9diEqFJwpYLBnFKoaAaHmVv/le
RZtpKkc7mEErY8rEQB5kP2sBCtEQtOEbxH/cqfDDuexw9OEQsY+vUzUM6K1SpHSg
h7leN5h/5iMZ/GW8duzT8azTpDmm4d/+2PalwmkdmagCbAO88Xfi9x1oXdEWdidP
6RaBkP36qFWHHeoC5O/Z2q1m6+vppH7Hvfq/EhmgHEE0s7WqhfJObOepnxxcLo4s
xSrilRyu+ZIMqSjrZTPLjb/+YNI7iJXHgkBxzhUhJqes7QjlKQX32A7NfixwGkg6
ZRRtlfUjwkswmcgMPByWQNN0i/C7gC8tKA+GCYkj3FJbUEqcne6DVc9DQG0lyPSJ
ReUz584mk1QqTGXo+Z1fC4PCrqUW6WOIsmycmbKVmptSmol7AcRS2FwfwZR4oGTf
ztsyIVhUo4SjcqW8w1ByjAEL14U+mTKzmOW1RpPHC2YrAWba6Oa1kfdHLNkEYhWT
pM5FW1eRS4gd3g1Om0UGRCrEybv4bNFvoaB+qy/vacYCoZvZIUTWfhk6tZ6eVoNa
aOcB1fi3+o7UnI8TxeNByJFbJvHM+OlBrVBkJPpDeZ0wIcA1Ts/f4Wu6fwKTz3yF
5joAtb1GoAMgc0TzLOduq7lyYr803Hvc0+/t3geO4/7u0PlV81zHMUz2w4+Wf2gK
oLZkOW2EkysSivER4ATt55oYPIS9LZOsM4wHQf/XpXJ1+eUEHl6CZpw5kr37hEQb
OsRG8enC2NGu42S3LQ10+nmRK1RN5ANnGsEDXsssXxfR+h9vKfzC+/we2QvdDQok
JMPLXdVrWQB88RIriKAdI7FDZu0GOUC82cG3/ItONo1T+2jxErzQMFIBMCOMG/QL
Z8t0gZ/b4QNqc5GWKxOdQ/wZmk5/m1H/gbd2BIO+27iDGXZ1W/CAEO3Ni5qDmLri
t4LRo7etqo7gFGA+PF48AZyeMqK9FvY4MT0RTg2SfRPpuwEc6crRpKXQ0ufdNUHr
pZCnEk68N05WVv1f4haBTnOe74MQkzOmRoA1lpIAij7cBvY6Ca+fda03dxb6caBo
gG2HPgcqLT7W67R+vsAq/zwaOUJ9xn69Rdc+qU/btcYuW0RHxyO88ha8VSOyaJAD
WTXY07eWPbC6Z2euB7DXMmCfPZQ+hdP+FsFqa+b1KrrDuoggb4IbJ+JybU9IV/w+
y2p3wZoOmvFbmWwyX8R99NLhKdWV5QbMAhjivMqf0HykkmdMYc7TDP0XGuCV+uDk
MXEmpvx7yZr8lHdib76hngu/w+3FoHSRg1ksLiU5u3UZeyj+DKHf/4mFHzDl9SBM
9H0mO67Ak7T5B64/ZF7CY+fxZJTDni7pQ0RHmixmn5dt76/iByxCTaQR1H1oSE27
7UDByCzSrLl8viKSX8Eewy5WX1zlQ8lUx8F4eupdqroSBuOWJAoWglR9t+TQdgfH
vebgT5d0euiiRoMenvycuB7We57hB5L+3lE1hjbn8gnAMgN3e0vazhRgSYJfcvqm
8lmO/Viua/e883fHAgYYspNF/jWvGI/si+ICPegGUWib0oIy3AOfCZRZV/i73B2F
wegZ3m8P+Rj4pVZRJ0SvMPRKYGvQKd6lbD7wUdLn5fs4DdPNWW5JPEgaoeaiYQJh
BUAN0JCCdDr1uGQ8cn4BNB7FV32ER6/llWPdutlnGDb4ApCWXWffD+TNYdvThNf4
z2I4hCJV8O359SWVmQGfDLgC4VrCG9MUIUXrcLkxkexPnTkq4JIhF+FdWRtG+7hW
o/ElJFuC1pfWbGUmBvDBaFyDlTXVJpkZj2r3EA0wSlOuEqSH/52z4irlzUtZQLD6
QdCD05J13OvgKnf0fweGIqrt5yOI1kMp04XgmVqgpxEM05fL6TAjAb2rUdDil3OC
JMKVU6rO3zJtAQ7Bey9pP4HbuwJcsmHIEsYrTpDixxbGqdZ6SmDhfLWKJkt2l1OA
mjjL8H/kjs5puORodv0pO0Wumj5QRF+JqKrEDUjSiLl/Sd6VObcMuEquIlaDObN/
AtZExpHeleBEf16JyDpzqybEAxNZ5i4uo0zJ3gxeBW3nrPaDXnXSEDNI3MRTDdm7
6QMPAPS1nVSVwQrJ9dutn+ZnC+mtr4DxMUdzuvbKM6jSE9DdxFctAatHyozSqWH2
DkXey0zkOaom27nOXQn/chDMWc8Rs3FgSEPOa34U2COGB6IcGtg4Rad2dXd35qlM
Ty2QIVo6wHWET0g5IaJNwZVS1gpJs+YphfaW2uBS9nHQfLIe9K0G/4hNdPUqonrR
MfrehmJWd5u77ze34GLAlwSV8yD+NFLNn+ux8Qj0ltRCWYfIIU+DwNIql1VymVsL
0yoqdc9R56kqAhMRX1fr59OAAxdsQ6UocNLsvNnXBv1yLiVuPBxe3sPn9jf0o0RQ
gPItiNvWvyVaW6N2MOSHkpPLKzY6VVnDQkRygxUJmhYYFlJoC+fAmT/0I+8oj7RP
4vaRmtfiQadgnjYFkOGh7pBEAfCiK4iHkqBA+90GDAp1Pq0AzmrU/PQMErgzCDrZ
jTxooHcD6RjjFEaIvxizJpftpn1++4+bevsk93uhMLBYlSIwHnzTeN9COhtKDm1F
YrrpbV1FVJBfF452n6glwgPgczzb26VM+/KTt3134s5qrfMq8i6TAePjIDKe1N/1
nFgoNSZmkivPhhBY/w3zbda2uGvZRupkAP4s9upZSB4MF6ehOdJ+ueWDMTKKLHeq
9kamqzCcHEVDiK/EhUrOQtsi2F4GaouR8WGTfpQ3T7vFORNp74aEFDGEAcgkRnnt
XLo6+ZjeMLSfnpZALKVg8rH3wrbTIMY82U2gPLzcwctCOXWtXj3uS2fIOAwWkq+8
A0aofH4Ux4ns4FtMfnHdVopa9NcjoW12XfQ6IukfIbL9pg/ND/vaLT8lKA+n75n/
FXZeRB6UUH9cM8VXrHihprKmEeghNeGXO1kbtzWUUAgKhB2c4aZmB2OlirY9zEo6
WknmZLL6g8W2d06mUb/XDSmyFgo7j9B2iRj1/tzcEbKLBSSELuyCePGfXy8pGkol
RyZoku4bBCWFlMf6KkYemlrNK2bDDPMyCKkRfkQZGRUqJ5YXW4TTPBtVXEpSWift
OD7SYfS4v85nzbmpYGm9XwQn0cuoShD40XWBQqTn+v4tIq8O2um7fkX5ZqyGqoqH
OikWLRzyplSwxfKdhOmcWyIJBQFcCGlUI4FXTdbaTFqRjhDu9CRHgfZVJOoSPtoL
QZt1yWmEv8yC1L680JHQub2/fP9P9K5zLeNi0vR3dGcMA6sQ7v6JV+ocHz59+3Xy
X+Ja7bqWpOXdcuBqSeVs1buvLJs9rAUlR4HX6cP1poCp9olgpUhApiRGJo0Q5nIX
Z2tfxFMLcxNdt+Zyw5gvj+qnYlW+s+j86dpbliBsqVkIC+cNy8sC2HHHPa4GrfBB
2YJSVnZnVSrfdEyCF1LDQlZ1yaJQJm0OciW5IIpkEVhZHy7KGUR1HCeibkRCsMCu
psLjg9PgU6aWAaK6SbtMJ8tUVulSplZIZPMbfhbYHL1oi/8UDXqVsuUmyUKBXRJU
rHOGWMIBpnos07Kb9c09huakmaXMjVMbZAME0iUnkDI23LbadiiM39We2upSnWkm
5+H6epkMEQOmamNy16QF7EHqyU+8z0BWvpwTB715qHQA4L4UuM+9+mY+S+feQ5/3
MMGMfwJsBFRj6fLAAIEIAcrcalwmO0BJ/EIYBSAoqy4lpH7NCjLjZdtIdAYGQyFr
A0sdG6Cdy5672ddV4zAo7WfQdVkLoLALPNEz9XSfGWyEllvuVi7bn0l70h4uvV+t
bP/Wmk6tWBsFHCcn27Zn++LdMyWAVGAIEgZcn6OHnTcXhPa/acQLd/wk10cifZPG
JkoBNS54rvbrDUkTHUJ8UMmihuFGRy6BuTSM3AyJyK7RwxQcssVqlWwV2E7jJGTh
8ZUuvC86tNIQVoqk9VGnGI2WzdjOT7w7eovfxwaDdMj87PpADSpUKzH0dIpRVTK0
4EuEQCmAV3OvEbQ1hm/dQdP7c1JyIzd28G9s6YyBQEcFTndHpQWq+FdkaSP4rwdu
GFnBRS9y4CNavxD51GXPEBd7993Vc9+5OPvplfM2Z0Ei3SaqBMe3U1LdndyedDj9
X48dDX63PsyRz8/WrK1mNnhh/fgUI54PEK5H+gAvaPbM1lN3EUQPAJ34p5/xBU9y
Gqu9I81s4+ozjPWZP8dCl8rTayP08H87WbcP6O4SLp+Alh7Y9/Lj542nqWTyHHAl
0W/V/+ztuRlXwEqdWkU1/bKrkcHFDaRGNefzxSCjqh8NPbyOodwq9E3y0Jmzc7t4
ppObN1lLZLXdUGT/Z/9awq7AV8ImtszewHOiLtFEw0zF0GuCcxtzvBM1Qx/FriTa
ANOe5GzRURXsFAmYFdhntoxG7d/V4xsC3pv7fqc0H8SOBixvlnBz9QkdM+soN/gs
At7+48KleobHiKHithpK3nK6CsoIhTXEh0pbOctXy4geDhVGB2RptSpUgJsC351/
RViMiY8Wl6ZDRi3w4ZJbIqeqjtKYE/oxXYrmXpo65Qr1/yBIZgKFmaS+yJTk57JU
fupoWHMXo0ocO53VIiRhKrwVk0ucFr9ZN8VL47syHRuewBVr0kkLhcsH6pv/+QxS
D8OCBmCfspX3LuPHkwgHA+4KkAW3ZUSipKcds7lZSC6TVXI7F/vQHSXefxgPrN5F
jlqVWbk6O27kV6oCIxAveX7h3b5lSBxpxHnj9+o/20/y9TB+sejadVO92jR7d1pn
YnXtlIlpFsOR8c2GCJ4iPhOl5L4T5WeylZ2V3orNFirq/goS50XNEdUYMuc3J8/U
EIvERwwVh3ZnNPIpNSD25AGpaJi4Z9Rjg+tNm+l2ZyEGVJzXvFr6tAzBx+FRO9JD
kKyozcQcqCZhfXRho7On8PGinOgMIBVxPTAuSVOaQe+6K/FSO9qXUGyzJ1D0V4Co
TkvQp35kBZOC9ru7tvH4Pqu+i2UlhJPLiVe7Pmnk5OczSmnejMERKAtPq5hdgjb2
AWuZptd/mLVS7mpCoW4nVQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
NKbBo/IdPeH7q/Qfr3hdXskkHPixpvqk66Ej5+35E0kpcKisLEkxovivRu5jBOWD
nit13il6KQIXMNkil2aeXqdThliN/8K8wud3Q10WywCWWhJyQR5gDJbtPz5kRncO
kak1nDIZA5yIrffXgTVkdbr7tQRVvYXyT9gcMhmb6Ont0XFs2g4Lpf6h6Z6Yfvqo
p55iLIzQ++1DJU6mDMGdXtK+zymGXEEReLNSNDFQn+IQZp47GhvXqViIOzBJpQFe
w94gHKxUPt8yM2rMuwY87InJcQ9jhaL12nx1vH+WqjkR+qzmNsRcLeEaS1T2YN4q
aAO0+BdSTCJr3lLCWRhwrw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4880 )
`pragma protect data_block
E1Q+AD36wjhkclQylh9juaEcLWagxGSrTWxd6AxuhMBi/EQ/UKJj4Q1Y49wgpr/w
rXNn5VTlhATF1NUDuzNRB5sDLRsR+LqGp7zmCoQciHavJi1OPE52jWM9VGubpNhF
NGuUlRToD6f7umES9/tf4t8Pj0F31fOKxfNbPXc5uLIVFB/xjtKDOE5BhUfsZajE
lHBQz440ezCUyiu4XkIkDhw/WCaRfLubIJS1cojw04TgVs4HavUXos/X3mtTL0SS
SWQlpA6JRr/0xRQYEipZgBMWnpS9StshItLWBQ7io8bYaibVUbTa0I+8HMGbQTql
SpK6uZJTGgkSIdQyOz/EJWpuHwoZOONgEw6VJ4tAq/1wUK3aZ5fTCXdcCTx9+rJB
5GXDS7RTR6X2vFC/Lb7Q7wxnLF0/Sp5OlJQl4Wf5H2/tH2dcG7VfM/A/S0sMkJaD
0I1KvP8BkMCuYhuh1pr9odudEKwOY9tpx8emUGatWEzoxW7HYPraiBZ1YCKNXTc5
v6NcDDjZpPG3edK9293+DXtGsc8AQS5vuEaC8jI0vfjfebLzUXMxexWFDB6VJwXo
mybrnTN3+bnTCcptltTyUc43MUWqTzN5ibcxAoH1LozPBGZU8NPOSsWXGoU6wXZv
gmqAMos2+x+elohzLnPnI89PYYIdbVJO+DwprLQUKcJAgPbXmIi1fKTWv9uZzsFw
Ggm8KB99i1F+otbWhcIDWncnsy/xqsdnuvN78x6xsf8kJnI9xq+3bjkKlETqqVaZ
beQKfj/sxrlznmEvUTR22JDYZa8lD57xwYcnAwbSyFi3Xefle8kHoUdObbcfDzcm
lhy5R8LYiReOTq7uDW2N61h+3aMWW9OAW9ZjQx8/mjYpZE/TjJ6yUmtPoZqA1Myr
drmXh0EVXFz1mJ+eK7PEXbKKrv8HxdbLeSwlhRFfyP8aZXvUWywyKqJmHw7U7y+2
96T1AMa00pY6rTU2Rf4uYtvGs7eYSI9OvEuP3L/Ih5wvWdx8f3bH1Bqngd99gYJJ
Fy5grW1z32fJHTsdG17KazsLY9MCiUhCbva4dV23eovBXzkl0vg/tP1uayZTEReV
RQuJMvaTqYL3T5u8LV0i9lN4JjqK6DYA7hN1yfrnfv/AQRL42/RL98QH9lcMVd6a
RbyaU6YnJFhIBPjxspJV1pUnwbyHs7yb5aJpv5wsEf+29X/RFniPCjbMZGatTeoK
hPzK47xwkVXjUiMWxe6uxGwJX5oguprEMkibxSZ7E3wF0DXrc5b+eUDPOY/O94Lg
8DfRHnU63U1tKOxZoRtVJ419qnprqWn2K5pH+Q4WxNvuEbKHZ01ThEpEu+pEpimm
dCBV88vB18U+qa1j0ZLaXKSny1WiV3BFBzl9ToAZ8rWSAfvqYoy/Pni9JZl6VhG7
uz+NYBdyZnLDX/Eb7fKKh9z6lInsknfIFVUXd2r/Gy3TtWndRvfARlyJrElpYaAx
5ZtQEI0iDDuQ4mpmWUStNpEF8p9akBhs0HlOlC8f1LT27T74LIS2hgGgzQ634ufu
mc2ZTzRowGl8z5aab98V91JCvjm6aBSs+fKGFzcK66oMLqR+geFcYDcC/j6/ge0m
6i8MQbEwy2opG4HWxmiDZN7nu1IiStGIuxmUmnvVd7Obx/VfW+dndt6F9Mc41SEF
LTYzHemcVpmqKsgaV+NbXuC0VFslL0pOdEkK3BcIlnbWAZGvdvrPY+Omu7SS/aJd
5UZe8FGAbhI5r2UhAtK+lU8sWAeNUEB5RDaq/MpITehDvCG0fsMHubI6SRDPuHe3
BDl6Hla4UyqKhg5oRFL3lDsy24UiKYMG1N+K7LRy9FtWJGxPD7qnNGCkmwM6fuv2
SSiFVuuEQy+r2RhoTFVZ1uZY8JMTstGlaoxMrP6a5hjsWoA759EIyFcDWJq8aO7a
5zcW3TefyV0cjqO3eLG3z93FKatqfgUEUNzySE831IDL9stWkB5ZoqPjAxG+Kv2l
FKrjcvVTclLcFEnBBScsWXJkrDbpgpMQxfHeegfxqtWSkUxat8M93bC4itTVmt/H
x2kPtqMxKcmeClaiIo43CsY8KiM3PtrQWkkf+uD3/sKa3ykw2jG/ydKEzVDFdzJ2
FxPx/Nu05QFquivOmXOPIemq0fNuJV02lEdEzQ9ouTMhe65JNn+Fc+TRqLJxDkbE
KFF13MmGSToA62n6Q3yG4vQ4YofuyAinMEvkuIG0iwU0l4g4c+D1tcJrx2zAzCVy
8QlUAzc8s/y1HR6mJJiqIHqGpUeTrgu0AXW1Pty9LMRc0lXu5J/DNQ2IIms7XuLd
uwPuZfbFxUo4HJYBAA1fVURnG/pPghb2CPjQjLPcfWXtJ6lmuHdQFIs/UBz86AXl
hg3/cPphRUId1EvfFUI5YlNQSrdOJHN/PcQERVNUgDM+xdzQVMh2j8JzRzAi8Ehb
RUqoiucuajIel6HR2AZx0DwFjciwNYsUT+Z4KPrLzBBIgFwKdHlqT+ELllRFtGOC
0qHgXrDc70Cm8Q1+cE/FuaxOCf3VSNi3dJrTpE1u9+WIOAYxTkoBAOOR41KRHpMf
2XY3lXu6HpFUWvz+pkS+lVKEFcMCT87sRbqsxIFNsruUaHCNljTTNMI09JFyX2WE
uIifhEhs0qEDikslb/uw1COTU+HLI0CdMX3wd++Z36UGdzgU5+ezeBahBP4w5ggO
8BXbcVejQjb3mWWSv+01d1bkEw/a648K2ByRvQlVU3+Q2KbtxPZqg12l+k03EUkb
SSzUckURTYMJuJLHd6ub/jCN3nLYTInNuI8CpTiccBjoiyusDSK+8mZ/8VebO3Xp
77WA3PAjFdOWKhTC96mIe8ITIVERfFBtyULiD7V8d4U75IBSfJzKotgQBmp5IQiM
mxU527Qp+t+2qQxpQ6ClbTVp7uHRVupoyeFjPYcAJJ8uWN+YCrnUTj2j+60neade
ZOEn5/MD41fcepgCQlRQ2YKvZ9u3zxQsvvCFzjfFLh5ydfWBQx+CxAYJv9PAtZvR
Ow6lb+SaRB4pNhMj1OzPO76TBAqqqO1acFc+SQQzzTB8KleM87bcXKCyMelSwMSP
+WqI2BVYayBYnp3prT7tJRftnfE1tNjvRlyiQb+LFGD8HyHNJELI7wxHFhydNbMV
ketyGWETQ3u5xFd4J8zH90U9NOJFdh77UPap0i6bLfRTmo2KoaYWzBRNEHuocLi0
Nq3Sc08He9I2Yln/56Kp0+jn7DwLdN+bVQkZHuG88edaSr5vRTyBCTPGOvRE4kUc
4P4p2t385xrjQE/R5laY3WobSqAUqf8KIHgTS+X5Cjc2+cAlqtD6GsCpU2RIedkk
KdQnBWcni6np+9uBA6Ok+e2fArtGv1lkLm9X1NbkPucotu3TG+BPRPoBsyjnAC9c
U9eX1Yesl/JWQFk6agPPPd9iEUCJ+rCwoPKpLiwIeaJf8TnpQExEN84R1LpseeRk
NnV5xuKuWKh07WFaRenmsnxihbXNhz1ZsNKQ3/aectFECzOLJu/ayul3zul04Nja
/A4ttIrHiJ2HugIXruasEd4Sg9DWD8te03JqLehB3Er8R+tU+4TT2GNTWxm8Lp29
g1TwDG8gvz+/pD/2VoH13hyKf8dKzIQe40Tb5lTKqxCh9VmW5BPjW2JrfiFVnAcF
s/EJQMSaGlS2jHCyIR4gChkWxqicdeUfzR0HT8XLM59bRzDBwTWPT0znCA+8yQZ2
ZTAwAEdKsNuAQ2fkhl/bM8JUbnIvXguDwSJTGaUEX5sLrATCdcgsjfEm5XkjL8JH
zR1lmt3Yy0hl63iJJ/WC4T1LPmK1xr8r52BQFGG39iJfLW93RoFbXP/MZcUOBiMD
dy8A9Jnek6at4FWjfeGmtD85i9+aGyBk4cThpojzcT+76tOXjQVSgx37j/uXYBEb
nAvFSGN+ispUcpOLaEoLwBXfTReH6SsLcNJUbJ2oVMH4wOKrZL6uWKcWvf58tZGj
6nsd/FkpaWQDQMfT8KNCjSbc/S83v6VzF0Bw5bGG26c9no7i4Ql6akV6+pU4U6sr
sYx2VX6CNTDwdXAXM6r8ggXqh5VSvWcUW/ktGMEZpi9rglP7Amtu71PkYekrdQAu
cyjTk5l2/9iUNbHJQVRD3tIWxU11+yiJ0sZwvayDb19NH9cORDAO4dnqJEq6neMC
TVwc47UfzcB+mN+FJLgE42sHSwWvtF8e87RT21bPJ0la+LugXSBMclrrtM4WScN/
ce1XGPEaKoGY3szfU3FF7ipW11t/2aZKoUCm/ixFwiDMTrMGJ1idaofdY5B+qNI9
4vSjpH+zMzkybtAVq2bRWdyh9bI0hyvmogJoI01Rorej+fjy6DxzRNmq+apQ01ab
ERYG9zO2VmpBPSK8oT2qsrP++OVqVJJi/fhn8AxR9X9/sOo/qSI2rl/chUMNhvDY
IrEqzICExJyEdQbU6tQrs6cL1cqTl3U4BuGD4GuGcVlt9fPscn31x9PzjL7LLXOs
xJ3M/6B1V7UH7LYLD/sWUN+AmvjDG8EAQUkDkeRfoKp7yrInNH8fXQ0LaI0qQwT8
5ba7mEsk6V7aocbClhp5vIbXimhIWxBpuXip0Xp/XcZ2u9a3PhUYMZ535ZzLlPYH
yZ5yUFhQ+Bu9fTy4Mfcif0hacQX+UHYela4nzFggLJduPlU8wJZHvpCGPQjPrSn8
2hgq96q46shhCqkkc0cr8bcAm0ZeYBUNMCrl1QWmGFZhBU2YGFEEKiVtwPdznf4D
Ibn/XAAaz3qIxDU8XjzjSdbYAnE5k+6cSL+xwdC/sTdzi6C+juUQ86fbUpaaR5It
Rv3fAuVhpdtEwP58EKbY0t9vxzxvx3K6qmcWyIt+IsZJLHAsY9bOr8SfwxAG3m7H
fpTPcY7u4lHyH+7TWKLvV0VG/MoVEWPayI1eU+m1HqzoH5de8wbn+fJxtt6uDiG1
kbwhiEVaAjEAHwo/CVxjoo4ROzQkYL0b4f7G5e6tEXstSYCavlNMLTqsF2MlehcQ
WH/yh4W/U0MK770XEMj3fr1LA23QaDdGbPRRhd2IY1VqT/09ooIIoSySyXMacRPl
MjXVwbhf/g90a3cav5q03xIPSHuqoWZrpQ4L591Wfpw0l222AZl5H8Jx15/GCXqb
txpDikyKrl4U94omcG7xBQvUkOqTAsna1zbtXdTIHrnlwBO1YwMNn4DpgCGXEe7y
2sSZOo95hswOlu72agxk3IANBkywhF8oz39gTDr2QKEJgVM6wbyS5Sf5hBEpjeGJ
7P4QjMQe4CmpOp1TulfIAU5XpUnra6/pOd/iF7LeckPDEH//CNoovcnKvB4lV4lD
t0+SjgRhX6txFZ/gVftiAEwUVDC3svwi0fi6JsFoe4DQEpn9fe+v9KFqeTj/fVnl
HELR/mOW9aEUB7F9WnhYlzSUU/9DtiBWaOZVMyqdbD0js7Nh140IveVbz+/AZbcy
WvICC4HU5RvkQZDs3E5/7ZzH/ji6yOiCj7NdPYdGa2txHhRZf/vnZI9/HpVKFpL9
MnR56v8ETO0ZbiOJLhEOpoNiv3+ws/kdEhksboHK3rxa6u/rf8K47w2/NjncKsnO
mPqUUrOgemuxgkwdb8jKlvtt4GhPvrhNPL9w/9B09XdOgJQu7q7irJIOEfThT5Kw
KT5RxmTxK970ZBgSIvMJiM+LfuhRMCrmhf9B6NUkf92CDDy2zp453xoowrnoqiNK
AGIV+Ao7z3BX0PD2MGY56a68P7A7eqHGLZzsRGtHzTFbDVT9V/78E/mHtS8GPxif
bKmIZZHppXK6zMsFYFbAn/EXpxNimfCfyEJuibl3j8JbPxto/8rvZF4VQc9GrKcD
iQoiLSAxbIExA/gtZE0NZMAJxDDwHXt8I5mhGTPVs2DexySxtz32hVrTIeQF3mQp
2pMv9ev8al/FQZQ3V8ZLPhuguMj9aw+OJZOdk/Y/0jzTC+cvJHBz8MX9VgFOnSOS
PRvE2qp20/A7BuA141nsmevH7D6se+0wRJu+EonPngcNu1W/13xxDssCMWi268gL
/xdEGC3f6RmU0M63bBCGqaRFh4xmVH2k+N0OluJb46IFS7km0R8zboRPefI+aTiR
yiXK6q3kpJR0RFqBbc74nb1qmj/0ao7YVugSgkrd3iMetfdH8S/HK9Zc+V6jraIM
qyfkX1ncQ2tPsG+IfaVdAl8mPdVkuxby3ySTEhenHhUcOpXRJiX+NwZz5GFBkbSI
Z02134z10E+v9bpZF+zRr40tHDTqdHxoIuifqY+W1CK49157tuJ2M5XmlNo94Wd2
svBkCPqr7TIyEK/Oi/ffxlMsDVuvQK4vc3V08tEPka//VQJzp6bU9Ql2l/G2p2WR
cfTfyOyjEerWenZRu/jqPg559w26aTyjme53TRKl3MdC28YaQbtQUOk7fWHAVy0w
/JcKiKV80liW54cyV7dpC+9jY5PQwzinZahjatO3hkvd6CeHD2XTZiO0GbLYKqRY
+2a7CpTHA6bui6QL3vZf5Wat21LGqUrkfoFEQxI7M2k=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Z/fkAfZ/60Gj97M0qCbAYTxFbtmmS/C+ZMInx2qMh24h+S/dBgujWlK7BJ04WP6z
vUnd/cQPVvf0tQ3Tje4gtepFIrdXjZ+aJsKKBNjaabd7qSRSlFlJd3UgsPDa4HOs
P8iDUz6hcgA9st8lHWKvlatwsgKP5Ldv4Tg6bCIxEBrhfuY+EY5n/UDe4h36Wdtx
/tCixyaayCbZvgp1vJDH7vGpiTC4uZUm5n2xu5bMXZMim1viAufOPEfEAty3q7Gg
JrWlZwq6SKTBK9Hd2AQL4S0Qs/aZxRW4RP+VnKbvyDD7qRubZw4iA1oJr21iYSn2
ekmyUzMArZoVqBXSQmbTBg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8992 )
`pragma protect data_block
1LW2mo/ynfEvPNWfw6QtxWkmXpGDgzcceIaCHMrYdeG76c/QMY7WdMLC8LCEAQr9
/0qbc4DmzIz+6nC59kHgwhelxEZ5u9CTMKH0DhNG7l03hLmIClGIITwPWq6DS2zl
0XaKL6y+K5mAiKxTST+XTM5XrNxRBBiWYaqbYG0/hxFVToQgkzyAoIATWeSyUTc+
v3MlyteIqRWacUIsPBls0mja5eGfoJpxgcRcjiquq3jUhhyxSZHUIA9j8GwL4n6d
dkiEYxQUaiLks6HK+H50PKCZ82BYnve2BFFRXuv9Q5ApbmXYlGawoJwbEgaIKqgs
jgEHarMCzy0Rj8jq61EWZFEOKh98e/hoJ2BiP7YlquKj8iTni105755ENV6Qj4Lr
h/1VOTyAT6qZclGp+tQ4i5iQKLWWbtknHXXGIMkCqYHQgoIcIDFvox5DEYdsSeGG
7ERwMY2r8UB0xH/LzJGlLkdic9xvvCReaqEv0zTLrN3CXJ+MMzFZF9/cKeq6TxkB
79djQZfK9DN8n2yrYA6FFX4kaEm3hKwPWlRMBz9f3fBtF1qkoU2aj+PUvS7KNHZF
Ucc3HEswHWbZsYwSXoAKIzJyjxYjKT91DhZFE1OiaXWFsQuYzyLCzSTnI/MXCmQO
E6ROcMQ+PYbNM6QO+zAgHBBZIIcD+tPwnr0VgZ8U05HSG6Bor+lduSvWq8upyJv4
k66mfycevzagJAGY4aekIHXnGlD9DbanSmKxlHqDdUb6nGrpvhx+9DLaip2zwnoc
1p+FpvFvOQXlyNcpFm6RqrbV630zRt0JdtA9YtTFEOuW0OmeYG/G1R1k7kVx30mb
e82/cYpzI0fDZBCBbfzo9f1SwhDNbxvm32xTpVk/rXgjW6mDVufjH8ze2Oy0+dia
hIF3LjWK68OGRUaJgaaiNTfO2VFm4VFY2T5AXK2t2nD46ayVC0rdM3GNsHeYujXB
OxBXcbErPavdMZvZ47oM0We3LzoyODuBEU2s+6wia094SKto62RNvYEPYzlWG83d
7Mu+Yg5iAFFFcfPAUTuGxHJz2YR899cy5bGatJOtF0ykBHLA90wOx78++AhqqW5h
UiUigPGC7WUAMoD3ZfxfXlOj40NKFw9JqUph+/KLdYMHV6SH00N8goEyoo0zJeFU
XYzcNEztD9a/h6rOd5Gy+I+mV4emv64OjbX0Vjs3/vgxitUGHFMbOkByN0JdqDVe
dGJ1Dd+R1I+lRZqaiocqT94uMHnQcLfWd20+3Fn3WKa7oRFjzQpJbhM5jTdiIce9
C8AuGi85Anr14hbu6xFZ4GKOkYisgeJ9rKZUM1bqhPOsqxZh72ZoGrVRl19UkHAq
dK2j3jVNzByLa4e8eTOgrssnuq55oRRkMZFNe6w6ST1Lx7Cvyfwk576Z0mI57dvG
fvVAkklox92VdCtszDxSh7EIdJIhbdR+/Ewdi/7zTpmlheTYlwql3eSj6YUcf3z6
2irj+kSpp2zyvSw1tY8buVmYefogI5dZ12AG6v4DIwWMUPO4McoNzKgvia/NQxI7
fifRWdHDSD0Bu03fA70af3hm7S51zE6Gu0D1LcN3xcLVxgAZGpf700wsrUAm5XN0
/MZfGb3xL8pXDFsIiyfSqSzoqf9L2C0/bIfKkwYVOVrlXnteCohj9UHCkVlEB4Tu
nTFzAqR0MafF48TkTav3cg9JoudBGYpP/Yx3p4zCjyYT0rTWHbMtDJ/8FCzodKu9
tPSJeZv0W5QIuhHFsQ16Gj/U69/ouzdsz4nMURHUmpY927Iof3r4x3sb/SPdQuEz
40s3Os61p2GxsUb0RIvliXp6hhRdy9xTZAGY1RTdjlk6Xr8m2oB7QBrX/J53m0Cx
Br28D69xWf8INcMIJCBKLHP1MzuYwDzlEcqc0b6BSHPbgJVv2ChSct+Khhi+aZfA
MQ4X6+r2ASsIiRar3KpgX5QDDArb+nHogeFYIAb/1LpUmoTUOcRIvV6akoy9THUV
kzDd97iblDUfsgd8+q67ZBSyPrkWTLiD+IWRxI+rMAi95k+a4n7rm9hrVPCUeeus
bOISPhfuO/XM902wm9sD6oTY3Er8iwBMFajFtcX+383FFx3pvS1R3aBKlERSCfTj
Zt8ngjARIE9r0CT81cy9QsfRxRJDEglG+1qw1FVAjhjeJM0grmoxY5nnlHhI97Pm
TcAuexACI3LIde+CIWwCRj5geMtvs7BIzezXPelBxMLYmpI7b05W5ayeWJrelHup
Uc+sL7yrI6fKpLvmCom6TAyPA+OBQTjgXFmcC41q/noBkI4SCB2IQDhB4H0FKWl2
lzm0ip5NQzWf+rYu9PmQrdehpxpF22NOYPqOPp5qZlQwIIvUR/8pV4PaFkn7Kgvt
eggY9yiOCgHWYVnz+NHf+YMw/1rVdQW8rY+pf0nbg3jhUW5vWoAmsEfwGsXkB3vu
2fK9wMEpkaZGHnrduoWR4ddIz4oBLpue0WRR+FLOCvl42AHifIwcq6Jmz13ZUXJq
RQRqXtHRGizBylNCjIQeKJM1ubwK0wWsPZFRrX4NQg0cW4Q1wsIe8HtqJ8CeJFDg
WuXBIAewgemd784n6LZh/aKyaNQ/SWLDyuNM8Jd1G0ep1Q1CsvL67vbVAt3JQaAx
PPwHYyrjFTospfa/n9NgHCekG9Pi7I74cke7VwJRaz0M6KeTygEDg0sk2Q7ObQju
yutbMV9VMEet6NjDUla4BQhV5g1wHDuzdmRLJamCv6MGWrjOOZlbYnw4+AhLfFrC
c8Uy4JkBBoCrxp0D/hZBGHBMkuAujl4rgOV778/gBOLqK5J8BRYnk9sNrEZcDVF3
D0XG3/Y4NYx7c3ehdag7M7Y43Oc/oNp9Zt8HmEBRoEF15mV/pNTNtXErZADT+In7
M8U7Gb1kNcBWMvy6zYjwYzVjvqaJBRpXG459aqmB4PuEp+pHvSIjR0ZcYS2sb5lR
ZISm6yTV8nB+2dwG71Wj8Is6WLsaIor2NnLCiXmGikzpslvCeR35HUSBT/7CSkg3
dJFxocPHVq8SOfo0qHVJ0RLlDC1PFmSXEvYAeHLWaJ4adDdIZDjpPu7xT4E6BFsv
VHjbqnY/6PhB/2N/yVJsDRM0wKtGLRb/srMOAWiXRhL0W1qFOSO+eIRoo0t0bVPh
Y7napGifkzbZDxosdEUS/LCHkqwviSol6r+s/1ThpGBeGYZAwvFQbJjbrXGH4qLg
6upxPdU+VlLS2ZuNWd0B3zY+Afi8tqCJR3zNwsHqc7JMACP/HUck523je/j1qYqA
UzWSQKl8QYlIS4a6WTBlfYpP/FTgUJNc4VBRQT0HSJDaGqLu0vzfIB6lGyYcLUsK
yM36sK7Gr7JzIYcU4+fHJwVOd6GCBlAiOhVsq68pJNpDDVK+vga5u2z1CHYzfiB7
TQMXvTlziqDF/btl0IizyPLS2jkQmD507Yw9Y/OcjEDYcj2mzZUa8DZaAaX/i/u7
vi4SwcU/ZTj0zVIHcyPOlGR+jMG76I4xuQk9xopCoTcSG+pzQgkM/tv0gxlDqiPu
wYPZ7kgUf5E5nyrKjT80VmPIK3sKRKNN/2MPclxfMjZ/bBn+sxhJfB4GOzasyuYW
i9XiHbvx0fImknO8vTANa48iLNO1bAvGS85E4SWhQ8o7oxYc+zQyVXBAQqf//z7Z
4QAshpKLWhQQIj0KSNhVNCki4wG2RgrllW0UfWBn8QTYjGt2nJ91TOZpISjFyD20
GBGXANj69xeyp94CnX4HykZUrOdPmtIuG5chmmAVd/wxvuQhFJWpZibT5fN6XSTk
n2yWCtCoghqWhWwjGPt0y1zo/4NBBLDtJ4qNTofZzbZxKUYEXApUEkPXXS4quY96
IPvsEPJuHWdP9JNqOgApVE1RmeXgFrqsBDEVpr13Ogr8YBnvEMb34mkC/FNbI4Hb
5i9Qwhd3ZOqxNnXjZanMaFTMTiBsryp2FATTnZl+eZRFqgYSWDrSL39Gt22nvU0R
QeH0DwLEykjzkOSZiCgUwOl/WkwoAxY3GozIYSeqQlYXFcbpaeGQO+KmRB3ELBno
NDXCsiNelt0qSNVwc9rsMIFKMhTs+LV3ZFR9JJYFzrvTlIGJAbSAmVNt7uZNuvd1
RZItUKnjbhibztnVaaw3rrld+qLcZnmxb/AlOJ8ZNcnnvjNQIjQRE3drSsCbvr9B
9gc/4A6v1/RD70ixWlokSJlBgPuirpXIqZzPee7IhAvEgPQ/rpYSNGU2TuFE1YLH
nKSJ4xxZ+VxzYqOP6DBudXWsLH/o3ey5ebpdcQ/Btkq+MmZ/rwVnnGfaUSrgRT8g
itlw688dp79B5YNmmDIQqNdsv1005sKwN4G4aCTw3NXcf6iE0KrM5GpXKim8/SfC
FmmfA4d92p8I+m8tatjHqVmkcdZ7TIYj4tZvdRXbTZ+k59frdTldGPKtkIdxslSB
xs++535B1Hb5FYWfgQqX8FWHx+xLqNQDMwaxJF4OGT/CstoxHT4khZv85xz3HYeT
k2aA10ojaeOdgkbZIW/E7W8yCkgGcBnopqk8cNW4lmLydQoKWVhBYg/ed3Gbm5iA
ewVb6zDuDZXvv47eiHk1PKXnAbfeD7JItYJ1elOmca0hyLZo2eBBTYsxs9lZT9Ln
CXntYdDCxDV5LrLoL7X9ZisatgyBoSbmHNAc8+y2JUSMQc5lB8A/zXVip5b3S4J9
hn/3ugIS5ItxKE9xdxm4yAQWA/gKHEk6/TzDR8QQrxD7KOBwmVIQe8b4ugo5YPn/
G/QUVH9O2nGRfkxqWjtMhdWvVZWGmAsdKgibuQRTniJ0lbwkjv/BmZLmVW4Kvj80
F5JGfsGJEPzIt2ienbdQlmxTifqmOfKoEtnzIRa28XcycF9mAEZRB3OtTy/zYEwI
o/O+at9xTEsicCxOTjdsDtYKNLHFKvjB0ZB1QnN6LtL9rI2fohnhCz1vx4MFQRDI
0xvSHpaseRhCGCioUQNQGfyNXeflfKXVBD3EeHOwycScASEP2uAzWzPV71A7XzQo
OWMqg7AFrmnYBE+4EKUJz+FOE7dtXxHklKmZIA4ZbiEciUtcAZoTC772XPHv82Ch
cO59r2nyDC6RrHqGl8dbptjoGE0EtV/5C6Ll/0uUAqUCyJ9lGFc8IoqBS31MJcAL
NZ3XXBYwu95jkFfVLOKVflzs2ciM4E0opYHDgzSjeuHIivSHRevIgT1JP1lwNjmZ
tQTClilTwDrLs0ZqSdxRV9lRbWDR8jNxVAJNpEe0D8tXz99J29P5kdfe6bYOk4cy
Uc5DFUq285/CKJkg3hLxm4Rc3EKm8MzCyL3wYIsxpJ2b1TlAJ6dDIn8+mKqF/zTR
vuGUesslipo3KqPlX0NVgv8AHr/8UO7qCOFBpg3I0Xv/r2XSVoJyFlsrooKMlfBP
42dD2njRxFUsr/9tr2jf89eXec+Si/ABDjQNJ6ScQCZlX8lEyF0Bn2Hf4TldRWDe
ZOCHM/5LbIEDdUm/6rbhjb2xNcwOcwXPOaVsqDiIUvUQY18Pfp2rzR0fXurMBn41
uUfxKHAaO5OOHBWEcBz5CesUpQDQcuW1n+vcJBU/wM061CaYMPj3EgwmgQNvksPs
wEgCVvekWW2I6fDTgzdkFvc08IWktMTjWjrOEaC4fnxzZPDBFUjhP/Mf3jdghgjb
8vwZ+ylKYsquh2AfcZXRowFFpJPZ/x7f+hS//InglpmqqnBmzb6HZpWQDMOqnxMy
35BDcsQTOf9qLYdyatFJd2SpPhrjRATvESdUYP+pq9Xov/aY/Nfy73hRH3HW/4ys
yomgsVaLFG/tDCnAno2YGQKhniaMcQrO9A1NC0f+uUhWasZj5JYyb4innUF2tIV6
U51KfYM95pLnlNMg1xP43Y+14bmznmu8LKfsmQ344n044GrfoSJVhzcjLoeO2yoP
GvPozyudowlsgQN1aNVSzF1KPA1or9RWZgMp8D9VYk+iIg1Dp/5nMV4gV6Mk5Gei
+uwubSJjz9iuye4eIiQleZDP7oAXYqK0/OlqwDMHPQWxImXFqdg/xVjioGhsRyP0
s3kaVIl6xH7Xb+vG2nziKX1MqTUs/O+7q2u5KV/DZnICOWrmJz9vixN1JSHH0+m1
Zp9DQzbUQa+wkB01ayAN7mTaYrIKbyoIf2k4ssCzI9qGhqOZMtHXZAQNdjRO2x21
b3rhvr6lII3FTXg82gezSVh1v4hsG3Z0Mcf2hJDhJntKxPgUVbby6gPUByisvnZ1
0KvuEL3YNM0DZcr2B1PKxTJpWNAwmK6DMCrzxZVJikT9PJJf7DvFUL9lh9Ko0fgI
FRRHHTm3as9WQE0x0kaBhjnEHSODrEbXfh+TxRrj4/6C+gA9A5eGFIJH7WBloXOU
rRCvgmUcWqbsq1funsCf1FqcLjhDmOBv6xnKgVzGYtBttIDuhfz/jKCUgb8cKsl4
LItjNPNapDGyXXvzyb+Kjnjs1c6/4c7qtP43TYrYSTamkUbPsC1nwbqACknp5g5V
Dg5EuZ8ShKV1r8B7ijrYmEjPpgnCMM71z5oZr3ft+FC2Ard49t29So//u91TcPsB
IHhmZX6NY4BBf/cCqY97aWC3DPHd61MmqJR980Np199lkbd9zh2kfPKw6ieaywYh
VWHdfNtKzWD9qu/z3rfAsu7gyOJw9/geJNYCG3dqjt3vl2L7F3LjucYr1L7lMep5
x7QVFCrEYD34hMnRP5hHZ7eXXxRzaSaEFiIZh7sgPn5BlDSS7C/PQFSF5fzXkiwz
v4RjmNRB6+XgcM3ScTU1/OIP+R4n/kQXjer5LPrKwa4mMmrQiBpQKEkuzQovW6pR
2yqeXPP47pBjOuerV1BSYWlypCbpamoVa8hDnwf/PAkbZF5LOVHM6wM5QE3yjOn/
0MmhixbVpBR9Jx7qN9I7E1h5ICV4gbRbBZ4liLpPKoCQ2a81JVtzR393/eGHjIiW
w2lcwGW3qiKXhmw6MJ+dWc4ePt1fUzVxhJGBR/q/ddaAzOvn81SJpTSbEbo6ED0B
cXhRh6IMiLH8QIkB6zLKFbBgGxlaINutgeWqf9gF+jiguysGceaUahV7jOjw6yhs
GiJviBvw1aiAUmwx9t7nznaio69yawmhVib5UOTJlc09Q4PDSpRmBNIYAJS9fdFw
0Xgf+EttZGWbpNi98rXD+kmMvnJhgGW+BuQOeLKRvc/VMrqPYzvoK0UNH53MJXTX
dykbtU6TN8/3KD75nxTByvFL4AsRMWSYIx0KJ4/Q0F+XfrrucfTf6pDmPIgZl4mZ
6wxswQav4RcJ+1HwsNn23DfrYF1U7IdPYUN6qdf4C5s53hChnQqGgPa+kosI1lfY
XARVPchcae6IvESBzc8RqXGZt+oTaCKg6qv7mxW441XDtIuLer61Vsrq3nxYE62a
PfQI632KKcsLZ/VZaMkSweT2gla45Ny/+Bgkrc0M/KmAphy+9ZUYvwxaF9+pW7Ar
8zRDF08JwUFwJK0HXjEnf+pcaxjnRbk+bVUSiAj6RMaxjQ2OlL/nQ4N2gkf1WAqQ
AG7Yk12VfraHiwhRLZhEG7dqCimMS0T0O9e2rVu3ihwtwQC5d4C92lr0YyNAlP61
SdM7/wPMkrfEAka4hANY7yFFwR7XUkI5ulGr3AHZKO7tQM73cZd2FCGpdzE6CLcl
+fP3lmIUfEOkKwCWOgVGc3dla5n07oRE1rEbZgRrxpMGqI/b3YfPxWI6jS6aFM60
w3pXDcK0bXbJiR/mJixef4f1GmhiUv6N07B3hZSAtO6MfPCX2fHXyV4KyP4Vun6w
sin8WS3wbmsuX9/HRoBJIcbi2/EhTupbSt01ywXZsQd8zW58fC1xHwFFHpInplo1
GOD5ETZ0Zi0mipcu6U4t11h0IjXDz/7DoevKOQl/XQ2aLmnV7Aebw0a0StQ1somk
rZ9VKVBvcCWLx8qpFORWyAtxK73mZ5Mwt3yauISCCj+QTLDlymViGIe5TIP16GO4
MWCogOotDGrXRJohPWhDtmu2sbBRtsGDhDFkRk7QG8QscJgP8+iNNDGcYT1vOdMZ
1P+1WpqqcvFZszY7hlekbX1k4m+4BCRt1Mu1rNkEgSKCOBbkEdjH9GMhzn65d6j0
Pnlf4a3oyFmeA8e4rfM6P/L4PIFMk2fOT9szWdvrc+hTQ11dO8+ZBb9L0ggsicpl
rdt5KcYZrlsu/nNZhgYs9jmkkbAys/Vmx7LqspuG/Bp7S7Rwc9KRlNEuP/ZhHVUv
hEbsxa42q06TKzESoVR3jm66mDkQiySWDaNTSWEr5hRSEEN7zQrwy8+Jx9Sxgh6o
MQAiDiMeAsBZE8lKSDV4CAkSipF17hvfkrDwzD7s2DBsW+yEI9kpwDHhPD9SSNy6
aiJ8WA2gjcOmpV/s+xlXN3STtTGJKDYV6Gnu93Gy43bAmcomQVH0IKznt1FSwikR
EcWH7Ze10WL8IkTbGjW6tstRQ1ojO1lwmMwjVdehBzbevTlJeT+tXF1k3bHXxeq6
YQjgCZkyWr8JSy2mVBb8fGU4LBcU9e3BUT7FWABZBo5BRxl+yfIkY9WSw2xS6/k2
bERSnFVqX+P5pzA24yTbMsntmUB7wuz9zWCRWwxghlz8Q4+Htd7FHqm3diiFbIAj
DgxDyrl9wgycSJGfyvGBHJM+nHr3Ovu1oRL4qLkhy8cWopU/ChmKSZckHMk9hFJ6
m03lHeSiEaAQ0d94SbEsJOqkPYQBuQ7cWLj94XbeEgw1oRkNVflZniE1bccZ+jlq
D5e9bHfo36aBclL2JdXLzaGfzE6eE00ahRAOI3aCGTU0eMdZjFbDVUyjXHqQyt2v
EXDwn/oWFMdqP8I5WXm9g2am1xwbovQMd5rQR/6SwXyCYiM/nxNrtX2U9McCcuLE
7PoXjgwqbgULzJodb+0LW6EhiKuAwMVSh77R7vXnzvchMlLFsMOiuiS3XzVMKYUK
MzRFyJslyIRuKJK+PmB8uZniyOsgm5W4XzdleuTbbafkpjKkiGe0/gV1fRaUoGBm
OMETyb1xYVDJFN1OoS1KWRoBRZUg2m+TBMY+mfctQ82R/n142BEcjutii9m29htJ
Gw53qYrCQUEoKk8xweX+aEV0thSIJXzYyPF4PISZ2M5F+PBmjJtAx67eCG2UHdra
hiEYlMqkV5FlcY00yz4Lp/iYTlpVqnVrGrL6ZMtPiqCQh/MEqNCn8s7IBr2mLv0a
r6y0B3A+/H3FVRTve1QuW6mQmlw64T5Uasnb1uyVARxjF+Qn6j63/rVU/veMN/gW
sjZm6qoX7Hjyv5fVmS0Ex1EYTk2tJv51zgtrrEIKvU1Itie8IyqOKd6SwRfmJZXn
T2bpIjD3FapabMN1kAiE/SMKgy8NfTaGaaMUtI4zy+v9tZMM+lK1StHFY0l7DhUk
MV1gnj7bpRHLkxfpDc67HbznkTnnnlZNmBqNB5ZYFwOnn/0a8FfzRzuxVfDgTsVV
bROKTOyzasb7/Xp9/Pp7EgugGoo9lxaAq30yY/qdfhfXcKphyMrk9hIFBMGJjthN
bXPqwvViuIlYtXh+dt2JbnAzhItl+rxlKq0V7ZLkaM237QwY3T7HeP6DwEAwQ9KV
EMOMV4EpjHO8AFMvwXv4MkHgodzd8wS7LMzMk8o7f6Ic+sixy2+YPtm+LdvgIHPf
i1IsQWkv3R0kgBdlXchtx7MG5xKk3LjeQmCzJz3npMWL1ZMTDEekRGACSQ6z2Z8+
WgvOH2KI/QYnOT28a6BGd0UPRCVMJC6eXskbcnfrr67CnkP1N2VmxzrCZJOyeDcL
83til318P8jMKsy6qvUStEg1EiDA4TRJlYRPpTu1jXAAIKorohuZEs0+Hx1HyBh6
gvy4X6qKdf4pWSXN+xg6puj9GOACQJb89WMz3bTRMvekdX0kocYYFUE3tL+JxPOq
RjmKVRvilfYOOf0lt3sxrWFNZqBO+KsGs3uIGRV+eYUS0q7xEZlJk8wVbr/aDEDo
qj32sOMZMaKLRlTfEwXGh/cKzw8gOGh0szko60+2Dw4zOvQnYQAGMi1Uj4+XqKCS
YdCTxUdZGXQk709+kfOWt+/Aca8fjM2PtYcUidLrDD/IOoUfXi8vJzPYbbN/ed5P
JFBmLnyGVT2ClGO84eGqU2DMYhMKX9Ss+HhDHN9SbcCnLLkz4EleWUqMl8QBPgvB
9eBL3cImFPn9HmW9Bepi3X6kFGf3L8qzdAK8P5+w/G6JuETno4G0q66QInISvW3b
0rtvaIy/SYGIA14NAV2NN7z/J2SZoSXeShZLXskpTlPqgziMUrliuVmjF40GR6v+
8WiKYTHxqvqUX3OBz9xjNv/99qz4eVgGYU6zwigw7aNIMxjfUi0MzGDGfrFsbOek
v1Ah56Ykmw4Wm48Iq2KR5TlDPmiNH7LpEoH5e3SJdVlmhz7rz1LRXOJEMn5G+/4w
OPcGMabii8WlFQVRTozPITv2hNby8CNxbL34r3dBlNzlPv6RCxHJf3tVpVjG3gOD
8SHpklOPx588cPHTqx+LobNG0nd4RPWV7ZIEdW4cLZMbN6cMmTX/yyS8mVwo6BYu
n2NwGNOGRrtembs0O1bdfUVc/9D4dwla+fvlG91iBh1LZLDLi3yQrcvUr6W7ejfD
uBKyB0yTRs6sQdtk4O0IuvCitEA5E2Uq7vC1lqH2tq8AXSMimeJTANstOJVdWanH
s6Rq1RdY3e7wBVI8chEQnCrM2zASSMa5Koe88ChacYQ4+59ZlTLRJzV3MhxgnSK2
ovlFYKiXHuUpWtT1UuyJS72aMaVAJ06rx2NZf5CTMOndpUjQ/aGy7RrxtUg9h9Mg
tcJf4kxMRyJ9bIIcHSs866i9ZooSrRdvWX0xYXuv6hmMqaLk3ulkSs8/4uiwbnWn
tfvhcBwERb4fcf9zmQ48+4xqKfscAlZq2HdD+zc8Q2D+KBHRxusxb3ZC6e0vI+wN
So+2fl+IsA0NcVucOTFyLDdO6W8rkm+J1wlT3CVZ73MmhbdzSr4ddbS62pEqa/Nm
tbeVTRPPW+UX/KDe/Ryb1+Uc4zUe2sOjgVqYUdelafNVV7HZMF0B1mziHLBoRf75
UImNeUDDqSMqU4auDa4w4KxYofaddMyf6tcbs7Ou/PGwKou86Fw6ONgQJ4ld7Cna
hVKvyonZnwYnmj0/14oF5KwU9HMqC9bFSaxZk8xgh2z6geu1/nJVbyQR65RSFEF+
QX+1vDeJT9Mld1ldxjJdhExnje40x7nAkd80lT6PDH9t0NQgDM6dd5bA01wYjDD8
VdWYxSbGjqh3UnnzxN9lnlDrJISluzJ2br+/aeGnk8YV+GSLdlXMim4nVyj2Kplh
iiHux2nYKErh1v+1/F2J2xG+g/xv4XWUHmcYVz1wgXexSUFP8NKT9bcqlSlYyaSY
o1Az+Ik5LuUjWLVzH2midVa7o4+lJkeo26GmBClYlSDl9ugI7QGBsd1i7Gy5ydnk
KqsApXPQasZSES9zNk7rIJzMBNvHRmzTwwGlyFrLQKT9wFNbvOJkO8q34VER4tIm
QQ8Ttf0V5k9NSX7Hgl6M3HmmLnw89nH5MnIr6DahC7IrQLURDCtIcDG8y4rNAuBN
WL2GxPy/9nT2xDdX3P2O07bqgd/1Jrg+NMUdmXvSqK/Spt6gSDDQM5ysFRWrl+HQ
hhxDCjVNPtV902ty4jtkBi1WC/DXhiDGtSJo7FL5jtt1aP59mMeYVMoQVQ6XurMh
C5eNplhogah8pGGCAQEmdGU1I2hReq420CDkTXQU1cxd2KMmtMg2Gj7TnwHfQp5+
KQH99qqVAOrIFBuPDqI1bNhbhc4FRCMz4ZiZcXxi7Is1uE30+INAZgyJ+DbBLI9U
b1o19eDL2xbwTxP/xrWW3ANp8q98F1dbDhSRpfUALCZ+HunhmZJm8p3vfeHU2z8Q
PbcH/Vv/Vz4MQ6pV9LGtZi5vnW3QC+5Yk6IfLcW1Dr8eA55RrlnlakqsWWdGpe8l
WsUiAXAdwVa0zDb+GxWE7nzViKuQoH9VBfiUoQ0IaMiSsgSkdQbgwAXkDqrIR8YY
06PgiWJXL/0j84ztwyvEaw==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lpBeM3blZZZQDG4fKDGqC0DvdlPxyEna2X8tL+SfyjQLu1ldhg8TU2Wy3N/uRnU2
AFNCXY8PAhVSi0vpykZWuPVp4rRKhBMxeLM0S+z0KtyrNK9wrb46dN57/e2S72fu
aOiwpS2ZKacgriY8NjbXumH1jQDm+Sr8+UNGEGVOMeNruEbuU1Dggv7yhIyW+7Mr
aVHI1cZIByIKRi8Io2KDjt3iDoGBU7oXguxnXN0a+qSTDL9xY2YylGK8AKC7AlEl
WWw4WGJmldZdpx/GEC2clVvFEb8ggBRMOwM8vl5iDc5gTRG6XNLjvVoH0UJHJKsR
RdcquWDsYIBMyvfDQFT35g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
ULk6X6o5o1RGFBVPKnCDc8U9a/2nFB7L+iY9r7yRlyy4IZKhjWCg620AOvac0Mga
MnAojlq/Y1DsSF0mXR2woZQKfKk6nRGNQ8Ms4Fm+DhoeTfatE586Hee/2F9uXMBv
ZrOgwgthv7Qb1Pg4LSJvUL68xRiYI4YSMyEda5jLcgsIK/GoL7JVPDNWYjUdLCnV
93FFYyP8vGqMxxwP5awOpXTiSwqr3W2iwxZ+POfmk9z5Rm4NuBMAQ087WQGgJUUk
QYXWkLUvCKLQwtGfx1RphsrjDpq3GyHNqhJHMfJuW7AUv2zkhIVBx9ixh6agsoZM
uzyaYLM04sPzgcO5Dku2QlUwSNlxr7cgTkv7AbtbpRU07SDJt5U0PmjhIxUU0dwX
kW7SrPRxjJz/68xXQ/v3U0ykSYdVDwkUmJNDFN29LNdCf31EsKCR0KUyKNECkNUR
s1tl4Ew45a3gFDTvFom1+xkF7F5z+OlYYfLZ0q5Ke54CyDGGqqrLLA1D0vUMuRm7
6zZiP3Bf63zIbrSNCBhhiafAMbU0krHoGMcV3RRi8A0gqKpisa58uxYj1Puk/61f
66EgvqAPI78FYocMMsmds2JFD7bMy1X4O6c1yx+quThTZaiiZry62co7mYOrWTmF
s4yukE4OJYDyMMseJXyacilMWoRiV1ehgRXjrFqundC2r7X6EH4+yduDRTb8+uVm
+I3ZdvCpygoW3/7LtDfcjICA11wLB/3R9zwvlCeF3Y666WXYOWFHhyGMEcJzBGf6
MU85+BX2RPDMQYN6yFDWJHoIfD9Dy6E26/iwTinhQGIQDkdTpjNqN3KqXO8SVuic
ZdXV/cVc8WvpQYqxLq2epDOLKrKniiSJb8E9ji0hLFUKF0j2A9J7rgh8qxUTgl6I
jYkxj3oeCYmiYp8jc4d2dplHlLR7NXm1ngE8qsUYIHyA5HeR84ZVlo3GZaThDZcb
PXT6IGlQ5EGvCT1hihbajxVQvabjm/6Da3bw5p4cV3/m1QTc2VaFjBpmN2jXpOIK
hXiBlujw2GCI3k/IFsmfGcRmyYiHKJA2sIH+ELm8MH3WMuk+VCRPfSmQdpTq6sKG
Ip+/rRdmho7v+pExgpXs/yS8YKqSpfPrTciwsCfFtC4vYAK5fm3suuW37bd9BIYf
KsI9yH+l7JG+jXOa78xVsIoeWByJeBCMqes6gZSmXS0JVYRu89dw46sJ8kFc4VWk
M7uSDTT1EQ2q+BmS8GDL8ThTcjiZa3zASqjNicM90nvW4KORKjUKeOfF/v3MrPY+
uADUndCuH7UfdJIoVksdemqvfJv4YKxRWev6O+q43hRer1YZ7lAfMnYMcfDJsYPb
upGYnxZzPkkKtn+W9lK6ZLuHQKsWCcOzxNb7dEkXfXGcXkEcHeHvqm0UlTQRLTfJ
uUX4orS53nsrghQO7/yUHG3a6dZVAcq+bUiGLsMoAVBxSi3dYdFApwNrLAXt6i2b
UaZVyjdLRewxqyOkloXnzUulS7a037kq6FBx+EPN3FB2tJQLErY53jP31ps1KTwO
veXeW7OgfNzAD8IZpZsvfpTaux3QdHw6KyyUaI/gZZrBHRxvkXt8i54LeaJDmxwe
3vachvLukPizEYlQwTjhNSi2yz9ZiSejyBvPEtWUYQ/Vf/tc354VxMOz2Y7AYm4b
kgTwVr1OdzAUz8/f+6/9S31BGsOzJzKry0pIMzIQUFMJ0XLruekjaPmpKMMnv5Td
EuqVQf4QCEy2pIfm3pVHgyvGsTj7RS9ltNKLtxTJspJXls9O0kH0ohJHbPKCnjxj
ZB4xTJhnc9SAqp+QmQqhrafFlv6bgvpLb3uJwUYKENmlTMmM7yac/ZB4rw/T4NMZ
J1J1k2tXlMUUitlsENOy3DSFUN8tllyToPODQUR68OthQroQnYa+lfJZ3JCAawXY
EyZTSXfuyCpoxOgJFJOZPEXUzhtX0xiNwfPgIzjUPWWoO1TDs2zX9ikXZJ2afAbW
jl3WMjXDP3WF+mq4fyybZ31QLIVq70oneFVFk5qo3l6ifA5i1wGxHf6lcK5b6N+S
SLpkFuMLTyoBO1VAfDBLIoEQHISwJRAJaYy7A1rGou3jAiXjtv3RK2KXfwqXxFez
VECqW3tbBQYlRIY+DqgRu5YOJlybgsyCd5g3MsuJfe3B46PI8bHJhTCjiGYSsgsq
TagNvOrgfH3ygr1DS5RG5zIQg0wipilTFrosJJG0qzrEUfJWalYNMVuwGkEalko5
rHzOfSXS6sTJZvs08Q5g0TnP2yXo/EKgDnamNt4Hmm5jrU1R84qAOHEm3zwJzCxi
7PosmwN8OhN1/y717kjHPxC3Gr+/dd3EEaIfBj1QHMJrvHGvYPG6Jb7YId7EVLFS
285fRvminrfGjL1wgzRIlPSMENZQ++OO2C+D2oJ9IIpTZbGvP0UFUyefrkEfvuiX
inFyZPsLK+SZ5NkleGSwWEi9FX2/14txnrg5x9uAPjBR0sk7PQBC8icg48QK3cef
o0kW245OqbGhKgrtY5E3TzU3iJ2Mq8VwaNRrM02DPYL1dxMiqbibXBbbDVyOjE6/
BcR1O8D5Vn2J/Ye5gg7Hs8RrXuoh0OVyj4Gdk/994P1tfE1Xx8gJAfrlb9Fu8Wfe
lqlf/N8vAb537tLBfv27jE3gJLDY3FSI9ym2WD64u6NCAy8Q8X2W6iPXBIKL5uAF
DrQJb5R3ujwdaJ3AXsAVwdCX9Qv/pjtFOnLnF+lB2/i7cgJhZDL8O4g+noyoq7AM
FSxaQnK8wayQKi7+aJd4jR5VRK4jjzyRQRESdRh0cgiydZTnX4Fo2dgAiOZfS27g
sbg6l3DuRXclHrDDjFamoWjos652pmffD/YgWpJoXvfeLnbb/dxG9s0nhgAGazdD
3Ec4hNiKeOuaMaY0LRsPXLpGTvXvRKOVs/8BUCfH3ildXm7j9uaZsDgiJOFI1TKF
D9uwnQRHnEW+mKT7He8vDmc1V7N5pBlWmV+rJyyz9NUpSp30UlS85WsvpMy/OBaZ
CJR66L1EIQ+beKAZh5SZuW4KXBzusalO0LH8fS9tsBnuMc3RskxsNJXIGbMrJ6QD
o7V3uwXPZMrOLtlgimVAnQcrKcUA567+XEhLag9SUgnsatGQhX80HYh57iCbxmMd
ZL2gJyWk7fkqFsAMzl7Pp7JkIQSCReNFpmsYXOozuN49eYN97p8clW4ZgzFlY7cd
bku5l1OepIjV3lkDNeiNfE8/3AZV8gyM2dKaFewBvaJnBx0+HxNPglnIop+7Qp53
4vbIONfr6VIymJacgphJpJHG5acWec3yPWGkQXlZsL0W+GTnNKsaGdHQPEuZ2FR0
BIsUk56fsrm+tp1gKuAPXbVL4D1IQdy9r38kaKBqe3W9S/Z97qmxEsqGZl+AnNg7
zzSIYmPWqa7B8chfRBzOe52lcWTOEtaZ59xyfy12QNdOFyN0TvU2dZrXWRlVK6PS
YvOg7XIF/fdveyLBFgCr1lm3KDADfoMYSeud4/JkpwLP0RQSFNlJ7Entjif9bOfn
3JI/9CXjWKBXhAGawj6sXPbwUAeM11uqwK3yW/27b429pLCoeng4DqLeLc6QIOGD
wM7BVGBc0AwlXmeR1NBi0hOSNOZE22iGO0uwh95xKPb+SknaXB+slvcJ3pc7IyXr
OMWYZnCBlEjWfofdA1ADmCFunPHdEp9QWIvPyte83ZRuEqWmSd38M3xiZ/FFVRX/
7zoZELCNZv61Ee8732K0jUPb3hWlsTlK20H+Y4AXWBV4FOa2Ch04hP7M/+o1QZ6X
CzaS6KQzkOs/4/qjdDMHADbHyku0fXktpNGdBFoY2uu2cXykNWxXKh4npWCWz/V7
5ZHfXz0PBzgkzey84FAChS/WZcmKp1CDBULlxVCj2oTFva/qOH8Ak9Xo282QrWUu
Ogud4C3eS19StwWMw3OLRCKB5TQeFo1xqGcLN4M4rM4HWHzWhHIKHXWTFdD1iRPd
674ISb+iEzIi1YPO05e4xoHrmQ9RJszosCuZVeeGbB6dIMgP1GX4Gbe1rj+JGUuC
WzxFqZCByZnXVBIibch+c3lEfRdavFyrUhGdluo0h92wSE5N29CX++PBhAGGUjka
u4fjjJlDx1pcRuVrKXdUBlK3NqOh790n/UXyfGUxfa1B8yT+/KW/YhLg9JZeQ+Uv
yI2JTEe9yQmEtGm5A8azLz+gS4/49rc9cus82Wd/HM85wbHuyYWTzwM+F2NnASC6
Y1tpR7S9GwmdRvRRyPM9qDbnK3tqSqq3uv+7MvVLelYahe2VIsut0p66T9bmwGLX
A11uW3exqgSDRQ8GRUkPrtTpu6r0u1ya85qwnZzryknfVLlytVxGGoSOFuFHIpBP
SxkL9s5Fcqbq/fk9VJg1h5fDUleAD2x6RATeVKPG7iNU9yPPqxV1GeMeLlygeQNC
sNMbUvyclT5L8LUKoLkV28GK7r0EIULKhXpG89/fdjnUvznmfUOF9LvqTwD2MHK6
Tow5TYYD7JjSYYYAmUOewJcFnvRIEAnJ0r/0TryPGbcKZN6U/IFwyOinIy+d1l9Z
2vYQ8dgAp3UFAsHPKShcemHtOa44hyI6JxrRvlgeppgyySBKfSXpYKW8Tt1SASC5
GDj710OcAUkm5IaXosCYIjQJ0mPJRlh7ML+vwoar22wKUTVFmWbCoQ6qn0Il9igz
yll3MhTfEN6Foav29KFRd/EoM17XAs0DzlVeC+q2xGQxL5oamPtg/umogqdGGkay
dTj1GqxpM0OdzaPHCnYC/+a3thyUokbJ3VyUtRI0TCNzUoDQr/B1iR3/1R5Q2k98
yjh0916AAXwFFuwLWngb50i2oEKC8OsWWnk8dZPZ2q2PBOBwEDuQaAQD3YMB3OOQ
eMPwRwvQqtcfKndQrOUYEdErbUFlWRQaZ6pNMFfIPMdX91KyWGEhmEnx3Hpx3dK/
yjn/JPOQWxXYmDTaYv5JWDccgtaoz12U2YMLrwaMTwBgfiabmJfSBLaUvwdm60eX
ywysnQyJtByuVxVj2ssBvpYXxrbv3VirZrbGUEtubxjUUAldc1K2PFnfuEdbvZKQ
PvZaj4s5qePpc0X3uCLEopABbSzkqdMV+z1Bd5zt+am0ScqcdWaW2mBFtqK8pFKX
VfjPhVNLYOn9GGvNHKo9yn4xHXyxRkcD2klyQ9s2OLA=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
b0oLyWxudE3VMfxCs2wUd7CPkd26BMcYBK2AqmHhYmzWKkT3y09ET9bXuEEeHWNE
seszGFvOFBQuyrGa39gLtHREOUGBORyp3Ljokjo2lWyNo34/2RsuDGojOshg8lRU
RUJidlPjgSiOoURJEpk9dDYI9lI5jDUoY25I5g6tPQMcfruOxQPo9NaGi7Zoxc25
TTxKdm1OBDZfnwlbs0qQ9E24ODmCjE6ciXQd38X7TqbL8Xl69esGz4P4wAEJ3aUm
rayAtGHtBTMPC7j6U/cFuNqvkeqlP+rtuWfvU6qrXwxUdZ+vAAebZNAeKCJczvzJ
pnAkxFiXX2g9W7nWjLU7jA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
i/bVMlOLC7JqYZE5d1FTXPYixdIOqrRCa8bKyvaiveQAdzRV0EC7lJWBlTmebNwn
/S/LMkz0gxyqShM0x27phLGNFGJJIaVfhOhSVbhEz/fWxZzoTxAX5y74IGujD4uE
SLHEWu7in5Z3x96FJck7zSBcUvK2AdasPCvDs396wvbKJjQAQn+0gD31eNwaOYPE
L5CxFLTGxlP/49Wt4ZtfkxcmHNQsR4+csowS93PO0VtY9vADcEsscByahCrFSm+r
cyED0U2T83zLgDSGj7UiA5mSxQ0dXNZ4uXStX4UTzUomyf6Wh2QvSGh9v1R9Mq5f
hPNe4Zj43SD+C5ePM+lZte0T1ORHehZhSG1PIlwWPnJSp5TpYbRGR3QcxSoZVD+t
tfr/NPA1z4OFDOidw4IRWQKFTFoJ/Esd1JRjH9jxz+uxR0GUXElOUTEwjpE4fSjO
C8WFcWlZE/m1/NGo/nDYDODQAWRiZTF7uz3UWH21h/GUTAeTSQ42fam7OYuPLJ8u
uuSZtBU0zloMd2VJHgQy3HfDkvYnPDLUPS+PBtKGJbxfvtBnQPLC/NwnRjIgfJFS
HjdqKEmnARKz/+ePeIcA/60YgF0cgGO0bFUhootTMOMwd9vHkSrsRpnJ8wH+MFjh
WCKX17gjXhACWdkUU7MdCHQJtGlBi+p4fpk/Te8vAs6YM2RLR32YDWsMDt7Gm7eY
KsC/pKIUib1qAkrD0f9v6aKp20Kokh6W926Knrunt8ORgpcVKLyU44jsrSHLqOyx
iMEt3mzanQ3ZTXsNACYluQjDRq1a+psCjP7TF+Xy+1q1T4uuAtJVqSyrdLqPj/A8
yHRk84Z8GpXX+og93XfUn6YVi2omUN5hv8mrYnhN0Hm90VDsPhp5LK10shrSmpKh
7awC0q1KPfhb7VJHlNcQl7iMOJnSMCXdzt1USsXI1HkANww2eWvcSoKVXAzh6mR6
ntDxUfSQecKXx9hvKmH2CKGqKNkltVFMlz3YNMnlpveT6DDfpS6BC7Mt134jfT/p
XAAHDZ7fa5BrGWnfiWwLJ0ldj46ISydcYRd/Gn5YZ7aZMsYqW/Ch5bnE/fyKKvTb
pzZrWwBI6dA4I2kGX5qvre0dXPKhM5HKpnYu0nZtzfFKT7hfteAERlMmPHmuXNaT
PDUrs+vzSyjB3e8gL2FIKgBfGVgeU2+qm49mh+l2tnpq8CzifVU5YjuqRPueKcON
PfHe5DyrR8m+vDO4F0bqEILGRpb+Dc4qJfCx6poVLKmN2qJsOVPZzkMUQaRrRsHk
wMg5tRWbXxLOWg2V4lZGe/4FC8JNBggEUGl9OZTraiHcqKeKTWhrD7ZLt54nxMsu
I3IDYbdyxpHtQ2ShjgE6VcCk3vkekb3a+88oNw4BsP9NpfVCeBqhUwyBrPPZrDZM
+vnhV3vAUv9yrSNwAN3RjzahRjn27hlB/sK/dz58dmlevB3FhftPWqF1K3YqPeFV
rTlQHx/i9IuTx8dHDPCW7KusaFNfCqZvHOMNaMDiJuvdv2sD2YHznrp1rZtLUBJS
jVNl8qM/efAGmfRnjj5lUMWtpVjFMLfXDXrSM2sB9FgXWWotznFuI6t1xL2TE/aT
ma2ar/eEzejI6ooIeECcRzNsl3bJTo/f/Q8v+cmR9FEid47Z8nWQMeTrawBJo1hY
gCu2ATqcaHMwQVV6zUjnViFWjFy4e7G//yVDUE2LlCc+l4vm4EUNmiZ2fSAk5O0E
6RJsBIgrU1UO+ub5ASksJFLX6zbWy1A+d4LHufLAmzKo6osqZOrEo4+cv8EmM7gp
NYESnEgby/vD9mF4vLbRr9KCjl/5lfyMn2/U2PCTFe9dY/YVXXZSR+usNFJR1Cpz
JYuwvJgfHJg5OkRGF3rqeWsfutlPLLvvRb3if65Y4HTMV00o3mIv8iLXn5vGdUYR
fwm2gyv9E9zO5Fp+FypvI3gzWtRP48gJyFV6ebfINGDbLtuxpn3U1fvi4TVLZlnu
+hQyCewvOB75qzCXwqses12ynkjV5fJcI8KdiQftAygSzUcKOykRbAqeyPLkpTt6
26iBzYCtNIcjRG3Ypn+Casqk+v4MRBqKDyTjL34UzS19a9Z2504YQLVhhXT84+A5
kf3AJ3k5LcsjHKU/KvFCuAb6EXC0mVmkZgrpCKwe77jUurIEUPDoDmCyoIAD/mdm
slPUNrp9cQhkWTDaBBS6YHA9HCx7sxLh0r3TSo3h5mSitVREauBU/ZMLgpTzCLI+
TLOuxYUK6UmkVOsVwZwk+pxoeU1jxdDTS7J+1+UdcG21SpyjNmZDFKlZ/Jk6762P
JY82kFDwQnmlpgTZDcmTMHg68jqn63m8yNEcOIHOoc9Rrtdw+Hldn65GVYEzAwkT
QaZXr1BDR8QuDxHlUC5QnQM1LYYyLBHlX/miEd6Gv9Q2uNV2Y1BPs1QX2GB4KyfG
7iIq08GZSHTeEC5EAAsrABbKsj88N/bHT5jBP9kyYFil/rFCEAFJIJppxdLO3NYU
fHUQJkI1SlijnAdlbe0Ys8yiNmmwmVJ0Yj1iZFP39ATRrsSsfdwGCkaiYpX78nXr
gPD7DDksJYpnkQFV5zfko6DbCL+VhluQoZ1E7S7c4DNhP34glWkaLlxACkSq6+NC
3JS0xRO+f8SGa6cnWVk/vaPGjkP15YQ9ROR3E+FOWZ8Yyilk92wV5b5V2dS+aB15
apDrQkpLeZVC25gkEr3OOBd7Q5jIwdQvSaxupaMrCar1iC55rsaGEuKpTkCwJDpU
56IovXlfoVtfIlCggAvnUDLWFPJWVofj88YywRgaPxPHXGmNo+QHrFsoeWD1VJN5
xUOmCnWcGCwVDXugPbAv7DJo1xb9B/uCECOQI9G3yyHV+msAB52BHJi0CW5Q/rsY
Z5sRmzNlz+dKx9OOtnATXAE39+8Yf2TeZ2uyCozz+hJdBDVRVjime4ytbc4wW5Si
UO+gjFqv8ghOSXLeWpy6q6bZQjJ8S0GXg1uOlqkf+SV8jnRuXy6vBhabigpu7LTL
nV8sv1MLysrODfGpxIpBifUdnrO6WvLi2Pnt66Oo0PG2ieymf0nHH6f4sgJvvSbP
/gu5iE6jDktYenvAicNcpBOBieXQWS4nuapZRjo5E8cXBDSO/VdIoTAPtk4/VD6Z
FlmfHYpbuVfJ4sUuh5MTC5H0Svuv1RcpiFyBLU12p0bHKaA3sydBXULfwTLt2rM8
QJNYWbNv+nlFcv2EGRcA+nhDpEtMdxMqIQ41O2TXB4exCUWqOHPZCoaIY54jxmhg
m0rbDim6sY4vy41mQWOTUHMQd3FlnvcMs5K1xm/P2h97yqvB5sSaXw73WwUmKs0P
AL7+giHxFfilLrvoI7vqDSaCgQApC2lxlQn6QcZiXrWcIQaePrDSfPtKQzs70SwC
NhD8gC57iOYXAXVbBQYpvevhN7cYyk3umCBBLm2L3lQRy+/SdEod219ByDayIktv
jFZPOND6Fp6vkeolF0F7oVPId4CBssQqLSh36einGH7gpS9xUZGl+XbKGb5w6yiB
EvGGdkLiN8qUrYhSyw17+sDcq3AIpDGEQISGkY2H2euHcEorddYXHT/0Ybyco2nh
oIwI0jzIc8sJAi2R9i7J+qmGmAWMcUCs4o+/ka82k+fmtckHJeQTMAE4C8LU6IIA
nf63PI9l4zo+XAhA8Q0NVYVkrf9m4t6/iDM2KfTwz1RQsr7g1mep4dvwYyVoI1k3
d3qD/a1u7vDtlhksnhW7OKwTlHO+WlBD8drQPcuiLoIqMcfLUcH/wz5N34z3TO4t
0Tk1V6YveGsgQ7IN8CP8LZGXw65ffxQVtPBVriNFss3CEuJpDSdzZ+RbWUqrwct7
lBfJKI+XvnrSXI4GvVvXFGP+kMJijK5VkwR9d1l7BGk3uLImK+uWBHPWu+yq/ozK
aKgubvmMC3zs93CKf5FdwGaurquDXH6egfXx8ag1zsxV+z+GPWq6g61gK7M0CYm0
h+FYzkg40v/LrjUe/MsGNVTe97/G76ieYj0/KGjWR95+PEK6CQX/BWwz8r/LwH9s
qMAdlCS9L8IVBTR2P0z/9SZo2uv6xyu1MPVACaVN4qljNYY0huB8vrGPXSvN8CdH
ld48NrndCckcll4RIQ20b2kzMOWn23LYD/YWlJ518DEZI0JOzxief6/LJ0D5gkKI
mJEZU0RvW8HHvXQByo0lS8AfEOMYRTkrC6pPNhhiPb7hNtpzilZrlSBI9RWw6jCT
bU88zKZ/9XDfwr9W8UNCoUAWxx6q6kuNuLiy+XDR2ciaFGU8qhvhFNTDXMLkNP/l
YP0PI67VIHqPYSh9o0vKy8w6KYvhgr512Uo+OfTJL563UvI17sPfY3n1RFTCoTCZ
lCl+j0PHcLTuOobrRKxqbRDifOIfMRYs0j1nFlTHCC5YVr3t+/CwJQ+0kr5bGYKZ
yUQ76PtVb18j81PeNKQQGr5unOFOgFuIRAxnfo8snDmC4j3RAdm+rJt87ML6I261
iJD3r0HmUC4oSpsWYNqlb09khBtSsYcRZMR3YtBVQb/F/aZ78AeAp4XExcXKsoRg
q0dxxg9E2h1ECl2wZXopV4jPmGsPKgaENJFu2MoP5EciSvmaLo6/bXN7/UaNYo5j
R5KdrI1mdRUdXyPfT9PankFdxLra0IOvx8H7h80cWycnKbl5Br5jBbo19YbormiR
ORL6LZadxjHI3liwBsIGrOnTkOGhtBNMwPSP6JM+FWTVWrrIRh5SVyobUKXVP6KT
hlPN+w6KRUs4+SMYmoHnNioR3Wp0jIT8EcgrvAfpso+P1HpCVf3rIIKEbIjdi9r/
sb4OYJeyXF0pCfBBqPebar96MVGrglEOBhX0KoOJw86is5rrqWVbAtUsbrzS0T+r
6mOLV+RBzdyjakICqZ1gcrMLgnZEsqtWckSY/JuDqtZLv9ZG8ehm6/Jlk9kT8M+0
pbvFVml2/vPNzqAMZnRTM4XNHZsEYtGQtS7cBWdrT735/MUaC5k/ywIEDcrTy+y/
nrUkmm8KJ0QS9lZWazduWlKz2Y73FbfSObhL1r2eX1Dbkf5j8c2Et9wMaE5fmIjA
gwWqqrVTp0y/wqNtfEjaBBeXnKRTrLWZaS7Ch+L5R4NCgPg40CHuIMKyAaN2uNBK
v2obPELrWhAfv7FmjVV+edRXyIg2B2dcea/wg7XSRLv4yQOVl3klj/wNhOHEBKCy
j09xLYuxQEJWrFxKPvvU9gp2f4d7EJk/XuTs/OgbRORpw214J1nXt+HHJIwiPrW/
UEvjYaMfVM9KZpFrFo2j+roc25j7rLVTEAJ8/hOu/xezmEcpLVtdxHYcThtmhmLZ
LhsRR2He5x932osgAxVh2LW4Qa91KXMMe5zDYbKDkSGtTOjn8aKal/2x0ygkXo89
0q63pzZQdnrV7otrvjxuKcVJ3GHAd8szuVzhDuaJlvmsV0bK/jnd8fw28kxUFyA3
eYmt3PER+PlQNcYBIwRsxRBZwZE+FfdYg7qeJIwPGMLiCx1wF9yTF0Ywzt/UXZTz
jWgk5Ok0h7tBgSp2b1JvF+BBTNazDdsncGMT80IHDlYb57rvidPQ/TwJkDTnEBfY
BsecbJaRFPBlWOlM1UsdzNd78uSHchJvUvu9N/poLhNL7MzgODSaJOp88A31pE36
FyUs0FCz3KDL6Tr6VM0qixdo5dVDuk4Pbqc0GcTqtGqwpINIpmMZHfKxu7hnMTJe
+VJ1Rf8RwsopMBX2H6hR6A4d2ALrg80p8XOGv20u8Nq7rIn4n7/OM/k323uw75uF
6ifJyjs5IePaCNkcrhWvWzAG6KkOQHYQ47Z1ONvLdXvQfgYDf0gUOHeRiZak0e7Z
KZDtLncbxAjNe3KKf0aEG/vqpg5eUJdwB42jmK2mjM+Zf6P+vr/TOo2ymK4PkDVz
ce+bkLrokDD8AhcRDe4iRPAdNg/zn/PfyO5Llo5/YBYkUYBWBo+aViyv6+rafOOR
mz5fAzwXs0y5H8l097Y4Q+ibj9+SkGKFG/UOkNaAKPEbxx6ZJ5nSeH4JnxN+uT/x
Ai2MCFf244y26Mcu6s3T0QGFVRr4P6tcwyFoATkU0oXn56yFReSx6x07FPJ1IGBT
os9dxtSJ+NU83e/0Hg6HUMizkSKhdhOf8iprAb2Bu1ArcVNtZ4LGRCQ8dSCVUBdL
tuHBpLelLU43meWbS1ySzGPKoPvIsAP76JtAn6z3VnzZniVxs2RBgywLu5YnsE4b
cHMQL1I2+MIYE5yCX5x71Ru4N3DHCcZ73Ns3bri/BPGepchQmIUiuxJRxaznSUdG
5ZKm741Gbbp+KjqcUrYEav+YG2QZ+wjTI1XO0czNRmwk5xtpvWNZN3DR2tiUOkUE
oIywT/OEuFksjizdEwYIC5pLzEsLmA3E+4NUssEUL3hWqprsLDgIrn+/BggRlhyT
0e+PGepktgJtuaJoxIZwT2KMaD3lHet/tIQXGgKBIsvuwIjUMOxqkB2s0C7A8OCm
Dg3wgOpKnNEbANWn1MfKEZsyTVxGn8Rlj5bqBZldgXvbhiTatvivMmH+eHlE3aVG
IhB6tpmbDRs/rdK4RgXlkfCBHi0/SCdyXRAyTtfwsmU3mx8kebCRM5u+P5SY5aQh
A4Hcue1VBg8n3hlwvaBJaFipGiAngDLEePW2qwEpJQL1Eh2gZ5U6ZDdiwERv+GP0
FYZu5f5SoNkAu9uaubBx+hqXFvXSugCmuyNF8Y76s7lMQieZ9leCDChvYdB4QNum
q0ojGfkk6SFsCa4470n+4mRqVEpgYOkdWdWSNrjNJbBQ81jltpbja2rc8aWoKcas
tgp6TPqX/nUCt6Q3vUPy+BsedKhMXM+QVRipVxWxDbz/g9pdV51t0W2F8ZjRdLKX
MDV694xWC94B2T7Em58YYyzmVYVWWK65nhpariU68pnorwHkbq0yCol/y8M12jdP
zHsEwnXtyQfJqoucf9q9dEANF37oiCdXQAqHnQkoi6wHX9AFwtC7yGBfjYrSF+qX
KbnkqBZNaMvFUfLbExiV93W0a8YgimKN4AXcRXW6i0QxLV40atJL0YQ1D+PJeiLy
k/ZC4dEm57sEHnC8AZy2dzgLjqHPBMyOHeDNGd16j4YZqHb0IwUx4ZW78DaByX20
nvtC0iJDALIlHSA0IX0FwrOVXz9dYnuoy7a3d57+cEImkqFvSk3ugjhPEFoB2Npl
SdJcdtqVjojz7b6uVh3hht13m4PVITWn/GV636aYTxytIA3vXPs0QnG58tAkQhYW
q7uocsDhNGK9DqdN8LXKcgMFKYmfIwObeRIyAElfHjnizwIMZOCinB4ICUBzghRu
8REl2wyCT8BNzIZ/sx1ZFlaDlkS2BN4V+8MFBWqX8SxJTORvvsrLD6gw3Oo4qI62
0CfFqWiLrH2sBwGPkOINbcNy4s1gN76kcfJDADCtuL5s2EHEOMayHpAEAIZYXDSJ
Jwg4TCYM9kXNpE+o5ly+cOzV+/PqgS63ooQ4SD41Q0WVudkf42Pz0dUdwxOoOoTR
P0+pye2aaavIZbW4UFLB40lxsqgLmlHNg1ETWal7kVs/lRVLo7/JcrPUHJI+PWvh
xr2+tWf7kLZ3LH3vzQoxlBC8ELZFcAJhDH0pia3dXfo/uQKAjwqK2SKaAVTocWpK
+AAI3bua1xCX0lDkNvCjMUj53DmXvEozxgJ7Y7jUEADUEnCTThflCnweqeALp0wI
O6KQ5S5sV3M5Qj3DsMTAhxsEymV6ECTD7EYS0DhIXTqZ9mNQdIEF9+8kdkFOdPd2
zC8ppYaJdOnOxOx9btGpbUTQdigIJI1zKszRu2pDkWM1TOo6NKsKapuvcu04y3Md
DsfSjsv0kEPLOzqXQlopKkbvV6uEH+tOV2523zg15B15UT6S70b8sAPAobzAnUV0
PxpwhJjnDISvkUMiv6gZ5+mpwP3pmoO5QH4dOuw6o/UcwgMNb90zc+oUj6qCVzX1
S0Age9X76i/+jLpcwkvP5Fx3Rl6gBe2UsxBzWPHMA91HbUy9ZFyZ7eU1fpWdSpmz
RmBY6uxUzYcKdcIR1ghQDbN1lXyJg8iIoY3FF3LaqJoEXT/z4TMCiFopfNAwUpxi
P1zfUjKBjYR6xZH2qdhRyGDDIBUs10gPLVAyPCBE6ZfXwtSfI3swOB4Fmd1P7Nfw
4g3sapKS/wvLypSm9LGI0AUwDy7eLbUSdXmSuoIRu7HQNCIgtkZyY/vMgESAGuB0
2KnoHWJz6WMm+s28Ey4UfUAMuUAqW3+ELj3VirsHF9e26HO5UVb/MPIXCcxklEps
P5Jmx9C9u0qRqrtku/6MeovV3dvDtg71WW408XFpfW6whQ5VVGPFsSqJy9dIjEN0
QpGHJUTUmLv1/UM/rx/8KPo/el/KvQ2JqPZqfyJhPkEKxYvhwL1Ve65Y1XqsDbSx
+Th3AAGRQUgPwi60denfynElXUVHP+gDHe+2BLTwLStZNPHAEuT/NmnZwW/T5fXk
aEflcw6X0qVDzx+AwMCgS+GyoLoFQXmY3zOu3nvWYPl5RXTXbY2cbj4z5UMGd+cW
skl04pD7vkcSoWAIwdLrXJ0j74APF2JBGgbjKT84ed6hCud7KYDibKpKY6MmI50A
oeruHqBWiZbDmYYpU2H93uFVZFRCPwU8HGQmiCuWKwXt6ROS3qlMJ/7SkrUeoFzV
YUp0TKu4XzLDe+7UgQ4ZcUj15YFeLC5hUYbpj7R1yL0ko6YALgrk+rRbWJUgkKE/
1orqfxJacbkEpf7bengLNGbrS/Ou58TK8qK+GQBOSAB5PTnAY0c2/y+gxHxkpBKV
f1+CYx2kzPjNXfuNUo9AOxyc6XoZRaSvXNcIkLXJd/cxW/eiMoHj7nSB23bclg72
vTauP4b6JCddItZ/m/qt4VpqUZCesw1dqzUJ191OqDIYKInFiJKNwKckOZLeMHlD
iTc0R4mlcggNu11tkRCgjeEqVBOirQRM6PijobGLNfYtuMtX1KrC2vWYvDZkIaYh
ed2B00Gp46KU/BOryp21YbTsePHTFEEewGGYDQqdGUkCTU9hCWZTYduKrSFHw8GQ
SLvyWKNsL0XYPr9U3N2Kik96b7SLjDMC8EjH1Z72kKtq1bhU8wq5XdWD1GJlabFG
VzQTdWeeDlQOa8t7LfYjjatj/lBw45qjtw+qcFr+3HtOTzO13oftZ+CdDLkBrgZM
YQXUumO7HnNLzlB3z9+SmHRgKlzHD8Q0JN1pos4aNny7NbaMUjvXdiKuMdgIg6s2
ys9ctqs4mFNLaY65g1ykWlnWwKoc5sBNi66L4aHXFK8m5hJtgz+ly3UFDKYcKk98
85Xtp/k8B795vQLGZsh3LnFNS7NA7OueLH8d6M0ZCJJmOMnRdhgPZUyeOEaMc0v9
xCLgQsORtpY6uWzwJBEy3Kv+pW0fmt6lATd8urChdLkVNICWjDNdEIEToL34YyoM
O+6dGim3Y3oKz7bsu+g2hqga/xaKuO2HRmvn6xPGQ6QGkPJffI9T8/zTt7HKYF5V
vDABLHpq2q2yNU7GolsHh3N9w7/hwEmeGjBYzouR3vNpXiaaPdp0ivhy5Ze7XDrF
ymOlwp5WGSsFGq6txves81JBVFS6fS2y3H6Sy7qU2kNjVvsErnv1rcF/vmrR2YHq
dgF1MtyH2IlaaTECNf0ttac86gbjp8tIrbp6iHZ7daAhJsDOac43UaWID7mg29RR
DtlE1jL1MB1pyoSbcK+1e3LXzhOIf0fLxu/hamAGuGu/kj5rxjpZLpjv2ZF5oXn7
1TYmGxX1nF/RzdgJANjQBzn/9eaSEqIT6fLDfALGMoGb/T/mqOeW2Dc8Yg2Ax7wT
VYVuQzWZnjGlaJN4B2P6DFvibJGqYO74Yn2LWxTaZ5RoYlN9BOc8wmgibtH1r8N4
4HHPXCWLZanm8APRzBUZ6J81qDi3l9sGUk8ZXa1hnKzUYAnhJGTQC+7XEhoHf606
07Qb7JnIZBQiRkzZGM3QHhChD0jPUp3xGhDtiQRXgF9CaCuvpddMuZ96aHw90kK3
1boyY+R7hD4Pe1DBsCS8KwViU3kDFoX+FBp80pSA1v4Jarg5AOcuUkIUiBCe9iBR
4FDQFIT76sVn102inKXxsvYaJ1bAP/lfcsFfa25reZqNBigNu2gXfRAlVxwRh6pi
oogexETcZWVKW0ynPqZUHvfxmIu+sZdG2yiZ2huIlLZEpwqLgeumG1XL5lDTzR1t
NuRM2bZkm9bdHN5AK3n0afqMwOFBJffoql2ZUlGM1M+29RogydZBXzUxzsP+54C+
Gt1bIfuuCxUTZdDC5ZAcwymVwc14cbTQYwJPQ/lLC6OgSOPn4oNHbXoxbC0Hb/aO
CW5uXClsMATqp5VfCCr3FB5bNrBQ64HHX2l5NTW8oI8DNp8vURMeGgW2kIB5XHIh
FuFn+a0HDvOEPQM6RhiPnoRS8aRHH45WTYxO6/v0hku64KDpY6K3r1Luc8SOu42X
qWZ5JF4/Kbp1a/em5RqKyb/EpukJLtHcyC0mA5Freb3NxNW9ydYMGt9Fn+nxynmz
JwPRkW8TausdeSdoDYwU0ew8sVOg6bU/wxA07XNoOOuifdYM35NP5t0qRLlSfVNl
yqz+uP8jB5kMKx74H9U2TgLIMnfEQ90knMGEQ5QO0Sq/wJJQwe6h73/m2BQFN2j+
A3hO90YeANaCVgmefH5yQY/LkCCH4oa6d538fMshjf9u0JOIlivwV7STB6GFiuTF
syDxOgFrxNeJrqI2bsZsCG/L8fPdD/WJeFHkxYxk7X8+wLX3XLxmeI9QB+YbX6bf
cX5RnT+jpeWaI1DTKkgkJsoEyV4ucAnP9/XE11MJbDNngzpWradC/3TU3vOmouK0
tBb8ZA2C3IHZf5KBVHY5csZcrtrMOLSRNyIwFz76VbFLfzQvHmxPkBo9QVbAJzgj
fwRhgwrrjOMYoQZAybHBeyl9uVhDSHTAktIX81zgeDoZurjASk1ikROs79w6BKUG
Zah5iD7AgmMxIK+siaGsDDwclI/g3nn2TUpvRVjmPcNur3J54lejR6SwGcqop6Uj
5shl5jCP0lbyZ9WIDVnfIN19hrTD3oTf+t1uWsal3JFbFxxRvxyrsZ//TkGh/iU0
IJu4Q5opva9LC0lAoQkOjocP/02gJtBp9LbP+4qshWT+a4plzFg9wvZxZpgE0x5E
KyD+AvpSE/HjW+xLKut9lw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ECnA2Y7fJK7DufxLfL2y0+BsSOgA8l4kJkdtumSBbs5gLx0net1F6epqBywPBMsi
zV1ea+XNJXDfQOtxiFTMyY4wneim37ejqFTWb8eEK5/6f6kWVYqApNyiXSkQnZRj
LcbWRefMcuM+VOXf+92R8alpL3YQIbP86uGD58DM3PFIAIvnnOcLkZiA69SZSD1H
hV9Q/NcDODAASsztbuffcSfi8n6Ogor81tq8dPfi989wrIYlUSM9M9yteHrspLgx
siHRSgO34uqaEHSMG/cLjNzMCQ7tqz+DivLgOZUTH/jy+bufD7qHDdTO7/fEPaEc
h68L5dnbkkP9kN7ZYgeB3A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10640 )
`pragma protect data_block
5wDydGWZfwAgIIxTQYqF/14C89ZsCP5o1H5jdYC0oQIwWw2ZiifUJgyEAW0n95ST
MRrsyN7sNiV322iZXmDTvgXp0GMHc6VOVSCO3nh2nX+gk1sOvMJesnZZZRiWwSTz
qhK7+LgzwRb7Oi7zdV1dMOz1xjqQhitQaGRPD1tPVjiTCVBtmWk43VXzyOO0NfX1
cErOJYyDOHzzeAQ0dBScx9cU9A+f4XEYnTjFShDYHHUYuxieeMw+HzjNCyPXdMNQ
U1n1IXCeecHEgzvEnjjM49/bC4RXoIREslCTMDbrJ50eBedrt/yjCqlywEwen/Qg
f0A0T4GWq4LceOa0wd1/eX01y8wdRrYKEeoO2ZtRcz6dN9HNV0JDwIIXuo8ycbRs
4GBSqE4X43Dtb7ZUUmWAsDdFdq5NqTiEbPrMr6mT2fym1It3KER03GxJhK6Ow9e5
C41yLDfh4uuHeFZAPK1aj04D9ViYKYvWVr7BxswdHlquWSLtnwLpCPAFLEFeOTRo
JLdZzhUMXJGY8wQmhvH/+mXbytQptGTiVCdP3pGRJ3X6X203MzN/eL2MlWZ1uBjR
iK3ytiyq5kEjp93QlcGWefkF5K4hVJmuqQGiscGxLlO+fs/DawupOCxCaA4sJXe8
h3ZjYQ725MieI1Kc0hgv5BWX0En9R1f02RKVlG2z5mGFTNbUDi5CUeG7QqJDjY+8
/+ukaG+idSrvY5Rmxwn4gnobc0Iote8cfAOxVf7v/tfFgq0018jKNPrDPc4Ogyue
t6TIPTYSkqUh0yMJwbPY5QRsd0YY46ruw65SNkExwzapPTja1l9+ONAfKGsqQBBI
ypsv1zXVGQGm+Ir2kHxmMUx4goT0TvVaUq/pXwqAxTXl+zgLtD5oWZgWgSPR+Gdl
xSUOfXTNR1KzTeSH21hdwCJ4CwgxnqmwUdewyIakXZu+sk9TiuVqgFXJgiQPGzgk
ApmHtfWcNeXzFrr8Ryi8xbsQqE1q1NK4bJh2TFGpEIqJ1Mv5/xoBa5KGdTg+GEgD
ZpQjxvzUMNzT5bYyD2H7oowY9WXN+qpjagNTWBvSvrqNsZ8NEoF4BzMx5+UT48m+
xNOjVA4pAWXU9tHB8S8hjEGafr0KHGCjsxqID8b9sKHuo1UMnlaPVOqZXgaHFYtK
TTAciPjytWl239Pt7yOakRap6s7ipm8jBgMIfOTu1gv1ghBOlIKrI3Ptopsxl718
6e0O3Gi7PTOCSiGExQuLCmXeRkIh2DJqJvzHTzYcRBj8jUI1OebnheD6tPBQgFPl
2tAo+oh+akIAyQQ5yFH0TgbBNzJ0jyQnGLrM6E7i/jGy+89UZSRdpValGMFH57vE
/huxOFp/o0qxxSvqELfuGC1y/DaaBv/+or157ASyK9nxx38AaEMJPNRlhVxiwE79
uNrQMVMA8PSCTz8UFir0ibXZolZhk7r5RNc4mks3qKafvX9pdFFOwC+dbLK/VH7i
utCCysXPB7VPe1IF8jQGSNp8Pm2FjsWl90HNT2Jx06mP3rin0psdP+d0McBrC1Lq
2pxDA/o0JtO/6lILjq9lB8rNP2YvnW+HnCHUigrWP7SyJO6p3JZPzvaJVKfkLiYl
lEBpU8gXU/JIbAy8Fw1WRVlsCgHIUHo0cq5zJwWudAFBo90N2AVQVWxUQBTGGASo
61d40mIVia+xuXaf2yTHz/gA6EiHmSyxvGCcHWKqfQxhWkrtlUf8oqAqFl+r4r/o
C0FcxOL4ZruSl/k5mBGPtjgcZ/LWLcuaHWJAH7bCNFbDFtjkx1r5Hz0vn19JvnmF
aCgBUCwwuHwTybsvT3Foaryv+BHz0zdg+iYP8rbr9Fq8Q3csrJ7jfU8WnFvSdRkP
ZlVNIraHF3Jma4+YZ089DeqQeDLMwTxkeEtbeSxHpBf1lnezog3Chf6P92S6UDlH
lmWFvdoDQPXzlfLEQB6UR7qMtNWfwICsdOVv2R2rsVK7uJaFMhVeFktlG/9BRfHd
aMtShq4YSdNKJXu0aLssHZXaEKNflM3XTWx3rHfGQz2m0JlDPXvggjP6UpMLONvy
sjrhaaHxyKNEEnkx5jC2IEYqXZhid/HuHhD4COUjZxxMulmlMGCqHCUgoWxOKxih
s1AeO5Omksp+Y5dm3UwwshGPihfhW/Sgpyvyt2WT8QN+6aptdw0eerJQAa/93uDO
AgNqL7rVCjxS0YVjsn9ywl/IzqEZ3sjpdj9w9MxfwfCYDfCg4eZCNScdi85Yr+l0
9HUb1yp0lIKaGGZZIptbYNWmTXdltTxrED0IvsD9vg+9BqaNLGYVqKM0oe+cykDR
s3h5zGdDYuphmdlP1bIC/lQ6mp559POmamO/iqILNXq70YFXYVAJ3UNGOC7SNQuW
VmL89zSz/QBD1fPF7QtCFoEnalOttQJVO3nuwrI2FElh9pa+zwgtymBq8fCuZZuf
+usdEHIYGNTwytphfc5ImkTNlxdtFUV8jhmWEBpEHNC/V44U7ln6HCnwyck0wBzP
zWbd68fZ90YXWtuD7VLAVIWtrD1SyK/jF4WX0VnjjgCj8AfV4LbWUfo7NCDKC9k3
yHOLrogdmU/Ez8/zZPUD9UfwvXWLT58P6NNX7K2BPAj4APRAsuUuhaSGcGHJjNkp
5RGWNoceiQJwHfujuL43ynpBTtygslLLfpzWIcmZf5Mm7MtMM23vnf45dDPvpsGQ
C3ZKMKW+8rG0tVvSKZ6QP6gme4ASla3CHHCranZWmQh6GudzY4JTk0ihEeTLcm9X
b05Yf9ea6JLSIHWjQfoJoF5PMKkIsHcqim93lf5wYGnmeek6g8/LnW9+9LYhv1Ww
ikZEecCS9v6In0MQqjjj8Vuzko2lAXeKinDQtAE4+bA445qNEA98SKofRxee53fN
DZOtwVGUt58+vDdLsu6kC42qVHNDe/wDY8BnTPlNl7fC+bKBTwe7CAtPxgnCLxhh
Dc2pmrJQnR5fQwl7+9nM7z3cKvU0vePkwj5/Umwyzhp+0ecm32eGelyBJHYREGFj
0JMTevzn9rbFnBHCXVsFwZCh+SaHfM3buRb3VgJljELEMgGUVbpypdc/QTUkkxoH
MncVPOzltnVQmPX9XrEx+RMuqpRZY/sLHFgiQzA+M6r5+kRklj5I8Y95LvZaXGOo
zQnSGapUeWNT64YO9gk3lt7DY9yJsL99vKll6D143oJAOPtT2bji8PO0vyiTTSWZ
9HJZnv1fY8MlqahPsdWa25Dh2zw8BAqP2YR9M0+xs+i/l3b+kE3rAf4Q1Wlz7JRS
FCp7qDd0vAmj5mOshndsk3VcgdNXvl1Tv88WmKQxqw3UEmVD5xgU447K6Ziv4x5m
tAvI797gtYybDdQRbhIgckecyS10eo6RSwS7ENFuv0ftkczwCZWAz6SK61B1M5po
2RHCcdI7qB+HQ4fgaugVvhZYUUEsO60ZuyZ9so0XKA3ueMlQWcHY6nO0dZdqkTlH
ZoSy/lv7Rz56XuXUrjHqj3JkrUhAthgadPtMJc1BFx+Pbfot7PioWTa6qh0FraRK
S8BUeMo2FJmZyxGpLAU8QLA50jVlH9Nu132Eo7nUzECXmyxNXKFzWdRKApbnBclQ
UBg0agg73b41blPtX7QhuiREjiviAeX51b4K2CbdIs1H1y6e+5fbc3VpfZuH7gUM
FnBGzys9/HGUv2wtB6f8HQDmKD89mwm3vCws2iyZiwHBDaUraxX8V59spxkyaDAY
rZwuCirkY2IYv9IroLCtmDronPiE8AocdI9e5W7c6byr3VVwfAUNwjtx0hDvRcf5
+jnOZ5+wuw7i/e2GvTi1utkg1TDZlyaVAPFKFpnewtEbQp7aQy0mWOmPDW+T5S1L
lWMpPK5Yl15Q3qCZFHM+A/ZDu3XM1SoK8ndk70qekuaW4cwJyfYxrg/GrPZK5O2a
swQrpOeKVNe7585TbXShEJqRem88DxyY5z78dtoBnK/svRMpaKYMYHYcRjU5eOuv
i6EDFWjVJs5A5YPMkqdmHAZugEn72qd6puYNHgG77RlxBwbrmlpb8NsCJA5dLMfL
MYpsLxTIbTbBB5QKhAaxAv+P3XtSf5QJBlOi1mR6pAjygg3hc+wxzMjBhum8GWgz
LJYJ0JK/ORqmplYsAUfqowFlAGWnYQsLxK+G1abMtdvoVeaw6OpkcDzWN4FTDrOn
BVLlG+YRAeCEj0oV2UocJh/gLnVg5p2wcSXHq7EB55iUsrD74tDcFMsPk/dLqitz
ElUF2PTveSpqqF6v1jWTL9A9NmT7jf03rlJOwx/fFqO89crCDKkKOV4fqa/l5n+m
KzNrxea21nekuVZs/p6Fh2Sm6Q9Ras78c0oxIOjUCviD6zGszo/7lWnogssyFEWk
kbugIiXD+c0ePOpUajiPe/7N4lwMXsLjy1m204lhszdTkiwNsHBxVJCGmpr/Z8c1
3KGXQmEMcYqmmiWpYL8Dw9mELky2y6She4iDGppFLwjeWyhWwomOw2Kq09UJyhnI
Ym16DiVy627dmxDE1OLGdN9oaUChdmVC2fPb7aSEXkJb0c8i70d4BAL6T3uLvE7k
BXe0xqse0A85HVCM3nlszO+EE36mz9tVWxLsW4slc9tdl2Xo8lCbhEggelyP7iMY
2iC/yLqD4a/xG/MbV+/FVe87vtgAPlE+AS3vo14f0E50bkOGLQeDkcCbPsODbW/7
BNu/c++MIZaH6k0pnbTJ/nhvNkjNXKXy0u+FmQT8neKMAPAvX/K1gVVVnnQTPuf9
8wrMgBKputLpLCQd8sF7KnmyZwCFaef3tXOt/BUjuKsAhIQA+RCaZwO35ivE8fRT
zeaa8Z71kJtU5/uANQ7c1O38LR1NEgV/A8KIJ94o2eGtnyCRX90cMwSMdfuPEPA4
k925cCQOesE3qcafcULvqyyxnAaurJnTzObHWX7VRXQE6Q/zxX9h+sbAw1/OigPy
YvKBz5ePMYvLf4KY4mMEC8fgu8s3C91gMbdk1vUtOqC+MWdt6MybOwdDaav/dXjc
OZFWs2clCQ7tSoywrEu2hIN5GgL3+T+Jk4dpwCd9lxjdQPPk4Da/9QDkusRRD1FV
QqGJvUdi6fd1tvEKukHFeFqxk2CsSyKUqfh6EzFkn1m4jB38YSuz1Pf6dEHfpKIA
UtT71y2Ac2geX7GrFIJ1FbkpcZMOofR+DzJypYMajbgldNr89pWmyCkk6CPZeSfB
VxTM6WYUo6lpulxJbSy2us6l44oeO2zqkvByGQ2jBVDSSOwakgOIwrilt16ReyBG
qqBqUrCFtrd/2BsOsQQhGakrOsyycgK9mdGDHDDTV+7SVH9//gLo7pStHRomOBhN
CNItUMihs2ZhOViHrh0m3z/Yaqi9VidjIRSnFe81QFs0JjReRvdLSelXFnBItO7M
UgaUuR4I7Of0jn9RGjDKRvzs3IDDn+RPWrfyxeAc4WMSHrOhm/zW8NxOf0THdt1y
OUGbHrQZMp3KYjHjMdnj/aYhsrIoUeB4KXRobVxAACN1F4neXun0z8xLkAm0p/Ey
Wp3sNmoCqCy+2+PvIPgocwtr2pfbvy/0BxD5whr4U8FAtrdV3/y+I+AdsXa6m++S
6socMMf/Y10GrtUpAfmLXCdZKUsc7CNi7m4/PmdKmvizTCqzFMCgBedsVZuvhViR
2ccYVV9xhgWxqUuiJ+CvfHfkwZFuo+Idzzjrh7whfWsJd9HdlmBtiArSVgGXUL4i
GhUHDRHdl7Hh+HcOeATO+6Juwsy++q4o8UGLchQyjlEWbh3r+nMslxH2GdUV1f9p
qpySzPyl2AiITtEXueaU8fq/B0E4OO1FBErWdvZGVo3Ru47WF00w83FLEO0B9dyq
+xQmclq8aZTs8tEDtxwM/Ji5jXIV5isl0dxlelWDRqXZHCvQFakuZwQrw3czE7Sl
ABN1cSlfWnISZkHOt3wZQ2hcDfqYVZrnzjstgmmj0wUiUcg+sBiYCo2Uemint/Yy
N5Ljgw03yYURiJthncSoRXCtb6dxAYK/Dd35NEyNrKz88kwh7X4qsf9V9+BJtrEe
qRG/wyz7eKPO7qBAh/otk159FO/QLFAz4KD/d7zWwkaKXRd8Rsh3dCW3zKORgXF8
qErC3eFsi856CQArrIcneu4+9UBgqCEfsGUQqXDwbzkcsv/T03ZFXm06Kkol/O8y
XqZRF77/N09kwrhUQMveQfQUJCCXL+U4yN6voIsNHrQ0DdIHxh4xE73VVBpXgWLs
UgF2EflxMJYYqeNmKcumVo191KellyjeAXRx+D8zkkTn/M3V6HL5oATTZdqCBEjL
0LqBEpab9P2CYOLv8lya4cp2RDg0SVwNZ1iEm7A3diqZr5gEguraHiuEmam/LhVp
b1nim2rR4UVUHhZhdpk+1yYBmGnq+xwPk43UEOthCQ8AIX+IeDSCypA92E4TnFB9
/qfvDOobipc4LGo2sGS1goQDJQyHDT3JdoZW/msCeLwVmTBRucCepT3QeCjrXrJR
MumUodqXUNIednGZpbCorNzfpLMhnqLn+Jf6QXLGPbMY6BexjVHCDDmzd1/2xsgC
qiQZH50mEwk4v/fFBA4z0ksfvC3nq+FQnIsfz4hk6iL3jj4DYyh1k5mSJB2i/BsP
wTtWcotjYOPJcnWnw5Q/gRdxQ8iPNALyX9gO5biB1Qe40P+PnKIgQ3ymGPXp0vtL
KDxlioYQ/ayw/yiVXtRvM+5EDdZy4j5hRhfTjuIMVuLuFia6JTHTDLYD5eQGb3wC
E2R5teCtWf0gYTX3XEhZ9ulm4ObWYWfNx4rTY2/EZP8qMA8iUy8h2hf6KeXKp8Wi
yUCPdJgh0idHI+TmeYEwMMEpYS8f3ekpH3k8OkdNQfd11RLJxKqm6/hTrdwBLRMi
RdFkT8cvtKZvd42AUf7w68kpuyJRg66iL4Q6cOEOsHiFajmCCQr5PaV2iJSCjp0s
iXcMaBf3B5eX6Ud/a1Ssf6NYz72EPCJpe4RXh2LgvrdvPgu6+TGzOqzGBIPeotST
15QsRX/eNFRsop8Yiz/RZX/xIrVOzD2AfZM22PyhjPFcy/d0cOE05wZ1PnXr194/
+lwTj91n1oPb0N+JT5hy+L4CpJUEU0Uy9/o2rJkP0ENb7OW/xwQguJ/hcZvcpl21
m1ds2y9lyU13mWoTK8cHdyMgcCaa0iR9HCKPRh2PtaJK0zvfaP36TiLeVBoUfzoH
f+qu6VgkP+QYRhcuLMb9QMY/0GGqHxN/filBrGgHpPvzaT8k4twqZ+mrPjT4vgb5
AfeIfffXaByGtZ2QCmp5RJcWPUos/olqyIDm2S1GgvFFkkw9V9BUEyf4KVCALy64
iQHt/KjM2uIhvy29SoOOTEQ85AHC7eD5FfQCh2BsPiydy4AI7DZzts7cqlG5v6Vc
U7KQCEfInxlSvOKqM5m8yDerI4iwKWv7r+SqeRbes2oPq6liVgtvUT2m5VCmri1W
LSNl7Gpe8kAFVzpbeHTfnfSOtp+TUSTOqj9Z0OVRZ7lWECGNxTdzW7UB97tznLIV
xe9gXTOaEp8U2mL0HiUyl6SvHteP1DGC8zT8tvMaMl7yWbLcdQyHgtirLaw1L0KZ
MAij2q/v/HfBG7m9DzgxpMz4PIISsZk7WdSJRsEMSd0pd4x/PxnaSbk6lrr/uiLs
Ym1p/OfveWUZHiY8zKlf8dWxvY9SfdhmB4CsAOOxAIEOTNfmV6Y3O+XKLHLzWCuP
aM/jLkZSfM3BREqGwLeawI614jk1RF0mH+pTj2T04w3zHhE9F1wysyrlrSVesL60
gyF2htNEKyDrTmH015VLTGYXezn8qlMEhdB27qxOwksZqruyb0LN7IxOd+Z1b0Ba
7Q2AnSzF6+USjhQZ3+jvK7DasUwrQ/fg+PKzqkoM8DE/chQdJ3S61SBHakVFmUKI
aY84riAkgnQ0rnpEmPb7MVDzlnDNTjdE+7VjLHz0kveD9wdiTY6lpicaNTQniS9R
Xft1CbNwjhq+CgHIZ9q9KZEG0onrBCwT5xjtmbryHGajOyNyYcE4cY/TgLdDG+vU
Igp4Jsu4nmowcL9dc5S3GLcso2dRsS9t58pTMEyMouawqNmV1GjOLxMFVyMam/iu
scAd7B6lzLFtIWpshLBccrSw16n9AmVunkFK7xGuLjTqlfe4HVfjhK9BINn0md3I
mRSIxaomHgV9jNUGCkLJt5ZN50DF+IFDub0Xp4pQBrNh+XGRVtLpMfj2UyAtYMqp
PL4ptn63p5s1Z9Dtms7TUXk1MPUQFUJSIvrAMyRvWfAe+f1lPqBEr5ffYgL5DLYM
wF0Baq417TwhiUe64XsVCF0PvB8TWa/azzcMTdY/VdvbOvrUIBIz1I0C2/cLUVei
OWYpakWC00Z32w70kpCIvF/h+xJAZRrvU4BGxl0gRsrMThGdAYdUIHCIMNw1nyvg
qYZu1spBGPGu/jfyOvhw6cI38kDD5ZWye3qdHZT4XYhN1o8ydoGbq+PjHWKnOCI4
knfiB5RsjyxOnJEeTT5O0PiWIyyzTdIa8inWKrRRck+NdNdsBL1nbPjVTcNCzgnT
qjMRQVgFdnXAdytu0BmyUcUIruqP3uV42gi8rrhaAXeDEYub4wZ7f0cdmhUw9efX
uyDBusPPIT6QAm1i0itwE00omSAZ3aAJ1TAoGoV1GRcGFw9XZ7pcCvuXnDbxRqvU
TQRbEw7h7yaSv/pfxFa/DY1/HUDRGnER+GLT8om3Dhn/5O+UWpn2f2mcpNbS1gJt
R29rMW+icISq4njC+uD5M9Yn99bJlh+Wtapuc+ZgvsFCfe7bRcoos7q58RoNpZMb
ih39sCXBVHPLH4oSaQlyRPs600n5Er+8IFN/1kKf+eTwgbH5wrc5J5rj/X9G2V/y
xzsUEsX1VdidiJ9bqiolpW1EdoeK6gkGynTVqWiT7EdziGjG2mHs61XT4sU+UtwJ
eTdtlRhdKb4pxNZcJLB2oREbPyYFcdpga1Fvj3DKAyT30trEhKc+m4y2VSr9+uPk
S3d7CO+kL0tV4UfKbtFu4ahGIeZ9Nuoku06ue4nSwmSM2iTho0cnI/bPuBEcT2OY
n7o7VtXz05vhnjv9pCLrat7f/fTUDgNbxyaSr6E0NjGrhSZq/thLWCSIiiUPEgmT
eo98BjJJ5bkPF9o5ubZ+6vvGmGdc3JmKjvd5yf6z+PpgN9qlnjFNZQZrhdoV1/DV
GVMHgel8Yr+SrY3tH7wnDVCcgPen18IJUuKsQPVQM+PPQZpNEW23TAxhaOj7htm3
3bjCfNiZD7T539jMHpKMdmgECChx9TwYVnIX5ibfSu4N4r6/PpY9500P6x2bJq6f
KCm2L/Tod3YZfQbOs4ZW7TrLQivVC/Nv3tO6eWaMz4pjkukBj2UgvccKq7sfe7OI
Y1a+XcNEubKhrp1RoSe3xWKLQBA5lspj/DZi3FlNUlZORCKGAU1WyZ/RBs4BKZhP
rwBA+SzUWKWxTCZL3SMx6LJ8NsOmO4ZNYJhxnAWWABoisiWaeuZwP8H3A7tCGEyh
qowniW9FkR1fHAlaO5qp1pSgp7QfTZz0K/rsO6PlDj98gIzAWytKmGwREksNhBd5
NT/Z09IlzrDRZoA9NK/14+jQq/VZPVNNBlMl/FRsibv5Dr/PUycogCUpUkMCMLC/
qGb4ChoFdzdiayRFr8amlxpba1adLNBiEhTdkTQZ+0ZVoP5dTJkpLv50KkdUMMBT
Bs+tZjF9y/3GVCjXgREWj6SjzFkK7Ek1LJY4K2W8+Hvg6wPZOTTi5IxmXq0+Hur/
TC0wqNrLoqA8tKW1yAlFOJcjOsMuwDWDriMNCDlFXQok8eOno2UZEMC3TuZB22zl
y3znIKZD33vKRoKxX372DDHtULj4RNKrnn41raF0X1bfaqa0G/4UrQA8P9DWqYZn
NTjP5e5lUaI1efU/HUD+Pb5ZSZFCWlQoOKb8jztwtZ4gvuH+/TEtsgqbbaAVrDqS
EWTWqHTg0wLJa2ILDvX3YGsP9PHft04VnJdpRwfWPdCUilJhvDYUlHtym5jfTCG9
9ItSqgtCJg91/SGi2kL6uI2e478zeNCk+q2HmGpNIiCHRTeQDArVsXcgvD2LayVW
Sv4SGD5wo1NS/2VzOLvvDivtWWibyBhmXeDoAPP01XewlambX5X9kgryU+LEEsMn
O7KTuj8xjiWD4p6XCunZN6t22xyrSUsdhlCqnOcDnijAPCdFEqZyX3eAj17EON2U
wEU6RIK71W0Kq1KTdjXvlrBeVuK310EoNzKtIXiRTBo49g0nXAQ7Z9B8DSVW11m/
ch3lQzSE1ocPmBI3TfcbsAeC+9mBC3OYh0nyWhdDcDOGA/ZO8h9G7HMFwKbNFB4A
RyTmOImI06jwkiotmYx+5bQBNzxLF1Kuf699SXV/8IH/Es41/r1ZSvcXnBsmreT/
MC+EqtyfWZxGv8n13/YiRUzPSa8Ve5fx55OGyB5Hu7Fyx9+ZkZbA8tyHUKzStZSp
XdPkLOo4BmJKGBzMK4HAOon3NiIa8HBzUlvJUpGGT4aTS/mWRwUkpIGP5Y5++Ylo
zEXZq3A5TutvWHjqsozd7aqMoh7nnIcZ4QGOwCkbXUC8Up8ZF54HTCRptLGvd67/
UMkQn+i9C5AcBrH6GARvQ2OLhGNH1xqpVBkftvt9U8qJ6Tj6+eYOAGHGn6+5zQB7
6aNUysJR1018gC6rIeu96XlP9v+u6AylDyfz812JlRVRRfoluRKLWZA4GafQpPh+
2gOAfrocCJZ4YsZFT8rh2EdsdMI1bHpF/EYz6EMhyettwwagfN4ZxYlDsDmrauAK
bBFh6vLw24s7moxHTrvaPx9FDLDCb2CV3q6i9uObNlC1Bs7/JXs5ujo7aFRmuyq8
66W+wG20/qPSb03stFpE9VHhxyApNBHr+3cTiiQJMQKOVaBeV59xhKqn1zhmHxJy
vDEmH+7ySTs+tutPtD0HSNaGU8/iSGCxKB+q94p6LbXpEdVHVL39feX/1f/XeYPI
IBLzZbPqr9WE0vGiD8o2wCHVXddkbrt2y3FlB94s2E7onpGHbRQpI8m+vpE7lnOD
96w3dL+KAQDOS/gmuKKmi33Y+QydhZRdJXFjtoEMm+T1505o2mXMzuf3QH2pqhq7
AKuOgsvPnB5KNkC+yoSq5rjZZ7+6JSANdhPoRSH+OpxdjR9mjA48U8tiDZCa/CuE
4ihcXNM15UUEzJeyF1a/9rnQx4GNOhUaTLbd2ucYThn8FWeQo1XopwoWvNakaIEM
/MbaVmUEhEZr2T9XDSvxLmP56+132YP4W/oSMN4ot01p+SD1tzdefkegQ0nGkE5d
Vcmeb2TrxvV0UZXbX9moSx+AHFtO8LwPxeNqYNScRIUM2zt/zVcifyZdjGg7vsl+
f6iRLGoeLBcmXsDj1/36rvbTpdwDmFpcXAKzOpJb3+RiYjROpAE/9W9avrjmuzU/
a7kNftgahBoBQ5LZjxx33LfhCwoX/2R9rtqY7fjnzQwCltjX+cFGZxd04PlvoSjb
olUjRdPkL4BOWvREWmnnNKKFJQuby6w7n39K4sR9OlBzpsfNKGfNE5Nr7RFEbM7Q
PQj5ux57gb6o/Ez2WWW9jABdsRqobVuguoRamsRSsmFrEsTY6POXB81yoHJAes/I
NJo673EsChc728a04jf+QsBIt0Uhd82gqZxKdjQP25XKk0ycgKIYdgonIK1xt9ba
vi2D/vneMU3xc1y/O5sKutAta/WhYEE0+lT3BEHnpEIN94S2Rx6gCJvXSZUFuOtV
jZX2ZhdaF2Y4HooC1j3XQeYwTDTjSDCL5b/ELo1WNabIFTIZkA6/swKATbJvne0B
GvMtUO565e4Ci2Kg8FevqmRPH4r6YPfROXaAzUixMEInox/TWcBatOF75wLY2IuZ
ZqifTumWqhmrd8ffq/XZ/9llDNAxMjYoGF+J7vVxBd4HhdBzuPsI9wOfBtHU0yDj
VXlkTT+avIFxVx+DxFiWcPo5qaExYVMNqvYbxNZeFVR66WsrxAadqdw/qacrKhP9
KBuz35JrMf9ww+QHNa2duTPFCQLDLTk1B2LqyYTtPyKK0QCijYGdZD/hbPAC9Xsa
7nu7CMRxHuLL4KUTnWS6evd5GYb6cvHK7919sG+cTVadCLiRxecA2S4x4QZ+DaYO
7IW03ayo1b0W70o8rNRfmCLfAd4Ik1Ox+pH3bMo79Vcosp401328KuuD3NRyTanC
XNChRzguga3eSMQ9DBBVMlh9ysrUjm/S826i6NpJ+Gsv0qBEVxK7pYAAr7NTi++O
xVWthRiAHphcFa052Tbc/GcTkQG2tGWSlURxyNQrTxD8TbQxNENFxuZGb0fl4RTW
/4fX5txzPAkcLVnbJM8CnRltkbsIwHlAcd1RC2Id/G+XArxl4TeqdyVec5M0CK8n
lCAkxXq6t97jlu/srNfSYrJ28NIgZ35BuN4deRg/MYFE47jZ7FPVFJJFWXZZUi1u
h2zn7xjUr+Z6BGGtweoT1uxk4vrmmSoKYT0Vwf78hOfpVzmDnIuVMR/JmvhwdoaC
zbzcs1X/BydyXhQEd7AEFdsgBW69V7vPX3Uk7geICW36JQsjMBxupCUL9dJt6ET5
SgzeQwyPnrwzQrkI3nLjq8/ndiduYKxwHotSs/MyrkYKQSgz6j8sXRNoqGoyiTCl
GaWZKTl/FLpGH3bY84YM7eoS5APm7rSpyU0DeVOIt6jqzlnCrPy0KgLV2gtMWd+/
VSbyeBtiNe728AcV5MnmbzhHaJvvMXTvqNZtg9GipngBv1eXc6LJx2aWFK3anYyB
Lc+xm/5vGlZR7ReyFlwvK3MXAUIuHXKbfCbu65+uGCKW57Nx8i+DmhcBH5zTVXK0
MRAqDMGDlSDs8YBhxaOf4H5UTIylqkDJV1ek2vDu5zRihj1tdMUpEfgeMXiazwN0
6F2i8+fX9OKN/PQ+Rp2b/MHh0414EdCro8k/7d/XxFSQhj/cbB9tuhuaqX2bugtA
BxirzlmAxy2j1Z0J+2m/xESX546ggZdvl0EKsXutY4/2IzRFP4WnFBSFkWB8zOL0
2la3AXbKdPT8Dhs0xiNwfZ5VaEUAVznLf53j7GHrDEdYXPODd7JzzDk+6ygYeFOX
hOEUTeT1X3Ct9SoVhJHrGGyRiBg1hIco1KYizF8RGtnowCbNI5OvAfVE7jzK4sLJ
ezLd0HluBtAfmH37Q6lA+vYr4dEBdp104+08LS6uhzjPfKkFd/G+30briSRiqn6r
H60EWV1RQsPz6OzqxAvPQvUVVNsRetum2XGstSpncGykvrVn44wZhOLaRLiGyJEv
fxWNHxo7iTr91GvG97O8Na39w47Sya3FPNDviEMArkedSUJ8rtkSBH8upiI3Wi1h
V4qfIGCloZCLRL9S7vRBOJjdcrU4dFXYI28s8844/hgepj5V/QTobTmYZLOzh7HD
Fi+jKL3yGe8Vsmjn4i55Hm1OQ7COerPCXDmLaCZbJeRjJd3MuojWmHmOdWnOS0oh
1YZTm8Uu0/Bs2i6S7kbJ5MsoOWhjGjgTjwM2gX1BoG2o+j3r3A34oggL4Uhz6Qm7
7II5wG4xLRDNNWJBZ4dZ04ruBPaR3s4npjVz8rFGZ+8dKTpVZ7dd/thxClmk7h5J
XI6KSsJ/5/DtkbzZnoUrT5KqKuQvQvgtXhRcFmDK8Pv0xqDMzigbxBNDDYJ6xMsx
gNHsVZM6jFch61GYazvOZmYYqQjDtSg1e6Y0q/Kv4jh8ZbPcnVdLDM/wxvtw5JYj
WkAh3B6Ha/cHonms+kZYNKF4kwGreBQiZrXzdRoGOmLqDuxSNG+50qO8WDjhKmSN
9948x1sNEXlcLtZigya3vmReYMYMlPoOg9rU2qeh7JDeQdCcjZeE+JHsmngpjFx0
Q2IRROBjZm4kucxpELkfQ4AXJUDr7g891WrHfDPNT6KBVAWpQ+AuwdvjoFl9SMfF
UoWSfmdjuq9kMLWWbJR0yjHO6Fv/1tuZ7kSApnnGJXmHc6I3waAmsYcE7m5NdjDD
Api0/bLE2U6iX0OltoCvNMXExJp5fSoIcFUM/tBaN8bu36w8qZmiPRPMU1dSvYFR
rDJ4eCre693u1CXtK8RGhOJZA3s9u08TRCCGh8uDwSnNu2tJmd354dw6CGi87gDj
8dNBa1UC3DQRtsLztKMfiLKgTVY/6PU2cgCsrkU5tb5fc67kADVfqFayyz6DtbOg
CMpPv0s6Z+DS6jPERnca/D8VRUi2Mhe5oV1c7q8HdyU=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
DxLBV/CG9WTUrX85UsGgyu0FQrs9qqpYHtML1dfnRRvl83v+1gpeTKlAS41XniRK
nFkdsaDIWiD4dmwetXdAPtqbjTfyZQlOTpnS8nqPJXVPD5KN7tFSjE5JW3FXZMry
yQbFWXNBZpUPNTq3IeI9brx0aHN8yRygMLDTMkVNcsRTeWw5xeZY7tZYY14dUSS/
MYA4FgJ0ou5xS/7EGqt9yhX/LKjNUXw52c80g2/yp3Pco2hcZZL/xT6s33EVatSL
BEF3pSFmqQyjuxi6lM9N3/iw3bdJgZyjm+DjbkmEvMX07pPi2OvAI6uWpR/GreZk
evPE1c28gN+091bVTIsq9g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2704 )
`pragma protect data_block
fh7cjNZWDOcP7OhIBvU28VLaDl3Z0Ntw9yof8YwWy8Bli+U1Y0fVW6Kp4elThR8g
BEIVmf8zu56jui/kWwSz184Zp77izevXJq217BQWJn6Ynmlx0kfujPUmqSACaNQ8
HCYbt5evXo46TGBp3rb7BpWk7xIuRnEtk9hYUcxIKPgXfHms7fcQl6KSmbVxoWUO
dxE9DPBfA5NLBpc89d/xtHyDDr6jn/kEBSvq/kEIdAZMLCbU8zkYZx9Cs/2yv3AQ
6QsGGDm7MwMiYOXzrPe8RcItXVkl154496BdJQxgxfxaaSYo5iHaMdswqG1MSL07
auMWCcG1QnicuYvrdixH0nZOzGJnwDORDxAZWxhqj4nCwHp8c2IkWIY3Nzrz0fox
p18yPWs84wwpuqahxSC4H4021INte7ohrcOv1m8k4ZJmrdnrS/TF/DVAYCGFU90I
75Sgx9SSBdvr4kkKcU30mlxXcJTvfQzgIZKj0uN06U/ItS6KoTigKBlkGey1WPLL
ec50HtAqOtIEtYwv9ntUD20DEbjGAaX8lwtmMpuec1FlnKenZB0ITKhspQODROki
D3TPaMVA2c41yOcF2q0ILpZA8J2b6b02y4oHZ1vxtgeVqcwq1aeiz5S3XzdCts4f
V97KMOVWOTDCmiQEF4gAzuAqIcxhoCvhF2vXtkFVDQz2bstdDSy0HnOp9QjtiCKJ
bFvzr9yWhx0qkVvrQer5B0ADsfj1o7Vh/7Mn4uaLcYgCrw6TLCL2rMfTk/Y3JRLk
E+Eh8LtiiFfcV63FbfRfLAQMUk/0JjcRa2mHHJTkKqpVWt9PATe6FrSZPZzR/hjF
eIy/tgJKSGQc3od8QAmYYKgaFI42pJoK6Wm0e2yIoFq3EjXGi4yxmTQfEmk6xxoG
++QQcuYNfy02gtRHOksFsuhOIHyERGDZHMNhvfmBhsgsicAAQWe/1I0k7/C212T+
diLjKdyxV2hQ1ckz3c4QRf6hvO+mQ+Rj0M2k5RTjWUP11t6ivACj0Vrz5Ihhwg27
MBDjjUeYUCujdj3XeBUwp4cKb041FQ0lCi3cXDL5TCrSj/N9V/UhPvBR1XtHAeJ2
vA92QPwyK7dAjcVVE2QnRl4jEA62QT3aB0MDbVZ6vaRjh3P64qBxkdXsK8HhFqfQ
fn3WaEhQ4BrVOOUnkzxnydEBv6c2oFMotSHi670dlIlrDEDJQu9zDX4Dmyw+0byr
N+F1xXQ0qDP96X5YM1wYwVmWOlufhyNaxCiKeL2cbV1C3Rx2EP60P6bJRRbuUCV/
av8wRqwIVpXCROJJA/KAx9YJyOk1MN37PudqxDcUmAzOS0Yl1BOxlRlWwAf6hAtk
DQSxC8fifxVsZhFw2I9dRWKGF8dYj8SbexYDgKUbsn9iifeQuJD3plDUs5lporTZ
j3nEfw4fR7DJhrlhzrOxSvr66ASUmlBtNdFcqS4C8u29UYDYr1dAwMyr2UMxmZUS
tArtkeHr4zSwjM7LPVGkwdXO+47oHUB4rrjfMb1H+3SdzebgrLDTzELfiqv+E4pE
csjGFJ4tpBDqK6ZhZyE969NeVKnMFU410ciZY3kgrAatIBNUBKnAabXPD2KvNOk/
ghVfIwVHl/iU89dpkr0EQbJhibyV6WhRYSWuCYCgYDxn1okfWyg82LgOsG+3bVDS
/ryTzDFev966FIhhqHhShSlJby+kzec67s9Sx1t1VsFyVLG7OXLZ0SJ7whoVZYhl
2ESwO1oRI4EvHlY7FXbrq6DmGMpO/INrhXFBqOvpKEixHQE/dBLvsSxbnHX5YDdF
rviM/l3pXC3ZmfJAxKByI54uoO3JkXfcfcRIZ3AxYOB0nna9Cd5VJ4BuEK2/dQ/R
qfhSjeDtGd8DzEg63TzWswum00roqNW4WjKsEHmxAS9//2P+ZNXhm0SeTG0Em6Ja
VbsYZkCkL9hEQ9fiYTkBqaRtYDJYK4ZLPgxaIISYs3Hnph7TGgL1wFqfKW9HEeCX
635jeo+uhQKYuIyir/Jw55RVn2Pho9StxfU0TPLzwrSj4ywr8NpewdNn/Sr05no+
KOdzkpDzXp48Ton3rrXRERUpeGHvcq94yAjG7J2q1dpyTV0FxkJMNJ3XK0llyNDo
0IzlmFgZkChtyEBhnwd5UxXTnN2XajxmqXIy5f6Kf6N+XPTkDb9oiah4TGgUe1bF
p1YYRXOTBw5LpDAQ/Di8CSA2Yr8m8QmdGo+/HikuUl/ZgL8d+qgx4L+vNHgZWsl0
QSAXWUwzLF4ft80pUS8x7pV9H6R0dNlJgD6M9uufC0jLVbNRAVl/dsfbuYpxoLIW
M6AnJy18AzUjLpeXtmtgb/RfrPasBDL1ZRxVWPMTv6I+berTATD9b9I3CuEyQ7eM
VMF8s5jJ+kecHuIvn7TET6SzWnsFr9aYB8C7WCIDcXhyiKwm/qqJF4j+0ZmM/bTw
N7Gfv1aCKpd9PlSzkCf60K10z3sp8xEPRzB4K/+pmaI9Ju+z7Oyc6YgdDxnIHml3
VxqpzIHUUwKPDt4eVdq+p4FRstul2mPDBJQjGo3y5UFehMmtBTD7p0cHiwUG+YtP
QYrgw6SZhPKm9Ob96Ra0Muh5uwyg9QsrEGRRkekame5TCj6COQeGcxtwIIfZE056
L20RWEDrc3RJwjuI3myG1CFFL6ZGuuUmRI83p4S1wrREHLz956KyGjRQPDBKGb1H
FHGn7W/3lFBEop+zyarm7h47BdevsZaXe4bP2ovd58lWAlHahSA+8Q8yE+ewKCzy
2I84caG6Saw3ZI+VmxqV1hUsKD3fqMR+xejsxXsBL5ERNOZmz3BJ6UiGspneuE21
bwZbTEylNZ6Z1MgLSrvzXYCFa4/5tAwA2m/n9axStlD11A6LRN7PU/4SZmdugnoi
NtrFe2zsMwFomYYNVDel1qw3zylAjqR7SxhZYF9oAA6pjmld/S7YV/0mcWN2BJmv
rpVDU5kJ0Fo7iaSvMUVq1dxNq/UXnASr59XaG32R2Zim/AjtNR3TdAJhkwJ4gXxN
AcLOmbdHtwrBVT07ObU53IrqRswFQsEeNc+FjQD7BL+uEgJYyZPN82EtU8G/4OtF
5hCs4XDdGzI+yNR/gLPyZ11QkWfmPaQFF/lywB8NRj44qLnxvKkSMb9CpfYnWLS7
iE/B+Z+5QN9ekMGVaaQeLluBvlflSBxEB4hTkFdkiP5+K6mLi1Q/uUglmvyvuddT
Jgj473zru3kYdx4HqHYBZJKE7RmZzUwoVK6XsY5LGi3deW9E1YjSGPsxYUPAutHF
IjzT/uVV4wiJX7BwEbV3CkFH1ogUzwAqFLiBqBdQOwZxu8NsoBJxqOa2jvR9RMNp
SOtNjtn3HQGB/+d1t8wSYjAx0ilqg+iLR9YgZGZbpyiTWzko3/OKX5mQ/Hyh6ylu
A1qqsTLrrClbq7MQ+8Mtovd6oL768KWKoYld7PaUQzrs18BlYTCZTMVHhPCZ2b1y
bMSlVI4c1LUPJ7FnFguccj6EbCpdNBhoopSA3zBQEKJDs4K4LlhgEbjx6ucNXbN/
QbZdfYnF4V594c8G3w+E5honpGIaRjdeMiVSzSiNqKfDRr5wUPNHLlCJHZnS4sfu
wNp8F1fu++0Fkaj8g4uvaA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
l8YCT6Ub8oAa9YAWAGMU6Y1HA/iCLl3z6FMHceCCJHPhbzJ9AR60tO7Ef0s+FK4j
wnTYzn16GIsW6cDXloTGf6bBRe6GCblzwk6g1owhWFvHwj/KzYpmQ/ZIYuIBOvRP
R00RrSdpNjpdVJtR4ITqV+VlRs3/0km3JXd7e8BrUHPQaYvidIZwMVJXi9jwar80
BpziZhmUsjrtOZQoES6kAoCfsZbMaGTNgWFSGc+VHabVh5PpXdeEMt3bo/rmmeOD
seBV8MOFBoIFOoHlYpttJeP8/nF+iRCl407Y1HsLXPvhHvZWfb8mJ5zjYyfNLYvO
gsb9Bdw4bYsZcba8vbtipg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8048 )
`pragma protect data_block
eMg3mdbg2rUMaDJtTfLTde2YVOaNI51JWMLTs8ZxmIlTrEsyD7vc7CkHWMnv44oW
FSCXnSBoI3o+722mUUWEzLQT5CTBbzWJpozZvKF752p3ReB/dEwwBjHtHA7pHUwE
kDaFL6ZJ5Pzuqzu5FY7ruIssgepIjrfeID+BVVpN1pymLOeJyq+C3ga+oEY46TVq
ohmo0XkAh6SUnbAhQROduWg8xWx0ivjOQ23+APFdbJVHVHwaJxv0D1Pifb1b6V52
RbRH1IsQgVlD8bCrj8UZ16wlOSvs3aW8e0+1w7tQKj6zZkRWh3+Y6Edme7nBo31W
kWXTqStXQaFIv7ejEay6Gh7+13sP9xMH0SBKXLZXriIfmkw1wzTNKgF6wGZ+SqXJ
B0QBOQUgH4In8pc3EYzC/6FMur/w0akQkKSYjjYypye5MG6/SdtsyJaSfpHxAY0a
hsl+lHJ9R7WQ8xpDG9JZ3azcrPZQaIjW+6BBBk2vk7fkqN6F7PrNrZ1Mgku3FGLn
Xvrc5kWQQM/+cGzKWvKAw5UIkfBg7h39XWTqUG9QqyHw3ISpV0FPeQWHngZeyB8I
1Hn9cyz1qkEXXQeaacozYTIAffOm75A34bh6ekDHGZVI853dk1OqGFgzzJkVjeSn
7mqxQgIYze2oaxI07PoGoMdB+398lbRblTVRYb4hQHF4m2mZAKIGQjLlkvWJa364
kJtQuqbB80u5+hvObRm/RTI3ekyWr6aV86Qp7eRwvOcIMdbsVBCK85aDq6SHkjTR
No3aryMS8Gmyi3B644bL8lUxlzcd5k3HabhN2fD1AJ71hDkmDy64KSnyQa5iuMT3
xTt+fe3Mt8eR6wrYFWPI8yj6+az+cJWv2oo85Tppb0gM7U7h4Ou8OPSoVipbtOlv
ctvjVc+/C3s1Cg3e79B+8j/MszB+je5nxTRho+rEh9SVKAcFt9BvnWe8MpTbDk6j
OCw7P47Xw9zWcmH58n+cTQTLyjSuSijAyNpS9F7ks8yH6yrHA1vLUgWbCIKSVhF3
Z/zijZyTDeoFdmAYJvL7udsVePCJOm4tqH9Rq1jPakOOSnquK1/uVBK9eay7QrNj
LuU2Ghz1vZLfyT6y9mU7ugM3omKxR1/qh7E+uObi2fqqSeXZ53aWDjWqgocelOKy
mdDijzKAKbp+Fb4pJD7U9hupizNitUzM9oBkmiQ5oJmk+Y8CQuB/MIL5osynwb0r
9EozWkkphCXSUGqvdw4CFxR9cYvHvLNpARZ3yalQ1gf4Sp2s+JegUdyWwCCfovLg
OormlTBx5NnBO67c8U7a9IlKn9a1glDstcM1owhvzEPIOUTtABr3ZcZNzBg17NDq
u+cVsT/5BW9tkqQ2Qs9WEg1HduKRhnUpU3igmWfYn7S4aONaArNM6pCgVmqNng8r
bBDrZswLheVq6sbcf899iPcoeKpznTryTLqftk/ggA3oL4nRkHnS3yMDkCNPv8PY
cyWNsgyjUt3zsYHzigzCsDcDMXOfyKG4sWk5qiQmGWAaJDNTVYAzpnEIsvjizFpx
Kz5JeTrN+L8OHqbHfdPSWg65ivL7MIDZ38J0S3XNvNtiloQ7y39rxbxajnTDIAHR
Qzic1qKXNNC77ZgN2sKISBuC4ktDxvvsxYrGCj/RqqiHDedBBjr7w40vFIXTe26J
5voKDqM0AdG98G9VcvO9r1dxqxdVvKm+PrNEBv2aJT1jMz5V5XJtbk2IeqNzJ7ZD
zRqPi2aLDShoAMpg5dhA2zB38ZUDfKVuwG2C6ViSS4ffK8qOtSio7aFKP3pPBnsn
dvgexcA/CH5zZk0Ue5Ns2qIm65cEyTCq2rzosfNtK3qzXa+lqNMPIrAdUdCoobwN
CPVvxjK1LR1GGHHmxjHkqaLLVw+lMaCoXl/eqhaa1CYnyLV1MH0JK/f3cHzKzWFP
gP16qJJL10pckDLpOA89SAM8BeW2pY41So8Y9YwwQpzMkIrsRujxy5RtNrDE62mk
cdoZrkzYzdx2g1PqNzYFHydsqXfGQjMjM85Wl/WH6s0JiUi07N8sl69SQ1i2mI7j
ygkzZfLaWbgP+4ff//oEox753O23nclLE8N72HUHexxTC6wLTpDF/kFEl46WUvxY
DFqyE7hNuD7wmPLx1K9/D4mYNXBUzWB4LJ9BXP4BWRnMujYiBVGvfGZn+pZvoFpw
50V92AO4RSaZyu13Hhydn5nHixCdevxHE9pF8x6siBV4gqYWR7U47QBIRoHvnndV
1uzkej4VIysHu+6GUpzRI4XTVQlrq4UIetqraTGr4edVhuraVmuhRRHPGYbtRYaq
o2Vi8UG0gmCmH/MzEu3I8zR2V+HR8Y1Ty0Ig/Q1xgN7zZ4WCineKbo+wfw1E+kuF
L1xUxYt3dWtgbn1ygo7XR42qmdatb4AhWJ3UEyy47Lh5nCESGeBP+KmrDOMEXwKB
zJK58m+ULGXIJ7wVpSfEWW3ckYgBU9iAqLCbO+NGdJzzFijOcy5Vkm7wIEvJbqPH
JqS53Hg2azy8OMzFi7jXbpMFC+TLnnkVoMiH3/bwopDo4czgozd7Mb/UOdIXheEf
PXTevDv3uCKbYdPJgFNIaAxPLackpFkskj2r9gQeCM22AIYA4nKHDHII9F0xxEfO
iWOP3TbS7xMVL8E9mBTCN1rCqI9FM++KeN21EjSOLttWMFuUNdluHnvUXRfENGtb
J+06D+AvOOcvPNnYXmd4QlwqmO+1jKZy0Y8sM/uXFWItGAvbZrcMOhIiJMcKTsYD
s7rFcqKJzgH4iDiRR3+q5p1WlNDMNSdf3oV3oIwjxVkp+I8Lz8k0mWPqb8QX/6rB
5DDRF9X+Fj+/0WZo8+/zwwWm1Kp3XGKs0g9q4HGcvV0mBkz0qpV5hxr6hw1MLnyv
C8Dh77eDKbll0xSOo2dlAJqkD/BBgE5PDjXPDhbrmJudUpubQ6mjAgI/SvKh6JKz
QNWW+pgB91453p1hSiouUkAHBydyJ3/rnnVJi5l3+8DZJzvxIGfQ9+QCW/pOCNtC
XX9eRk87YMr41zCUKIdbijQdKIO+VOzZX2bFzTmLtzIhIwfzyMIuS7RWtFNK9axG
U/kPK0xjtoZ/1EQolMYxVLZ0jxhrYs5fdpgZ8lk6moQ2nTP42sruViPi0DgtqRMW
iQCb22j+KbuS7tuEPVndut8vKme0M92qz0d/EglXY77TBQ8Nl4GkP5RoL8zhrK9l
kwtPmJe8JEJTmP96dZ7D+F+fapMFBIN3x0o9ufVUoWtZtoJzkwRkdPy3fQl/oBIl
YvSfVsdBupiTlObEeb9s0kDIZhnYDFrttHYKteUV+TCRuzN73NPRiYxsOqI2a0fE
CSOPtD1RaM14/EsITERhpBuBVRjCTkNom3+HyxdWY8J4L/fR1f5fuqWeRW0xt/OF
SwxpL32pTYgxCf1hy9YezZUMAY0XVxyQPPaP0Dp1NrdN/mhsW1HmagXXAu2pVg3i
DkYU5lsBK7SICXjj/zbVLW8owic/7Bio/QkEOqKD/ZJTMeV1kNUqOYFbTH7kaS5y
H1GNNGpXsLGD7TeHQLbdeUDBx7lRz8m4pXn/tFvi42YcP+NbZ/3hG0LZULZTpxCs
5EoF1Rg06QjQWhAO7i5OEKQyaEQuLEMC1cjXnxgY3X/V8Ja2VwvrmY3m7wVgBecB
t835kzadil0lznh6P9l/ZVqD0aBPItEEulSE/ZpwUgre7xRyfxkdgqpCkxa7Of1V
G4Y70MoekGRgJA2+PWtGKWrtBgL6NzG+9ZJeD6T7PeVIdX4O0eD6N+JU/T1H8Xe9
NiGMuY2dO1reOMAU7aEAgTy9UCk85lqvJwYEWwUqRmh+2XSiT41OVzeBCuBb8Rsz
cwAIyG3PpH7HVxbnNORNrkugysGojnr27Bqi2EF1cqx0exz0S+1OA2qXkWsjr/3k
hhbVNYbbt9pS20KlA2ldCR7ioTHpu333L60DWChsKeoTfVa7ap/gUAd2CRo1+s7W
fPTB27WvwP5BME4fgluryGjoNkbBM1OXv/IeSvdmjlHgYNDUwS4yqsqd785j3wbr
ZX2PgbSY8gMcAJ2X0hSiay1dvaGsWNLr4+Akrd8sb7dXCQQXv0XxVMT0ml/GfjlU
QE5+PE8R9w/hntpODJ7OaMFaCj5Yh2K5+sPnY1tOsNFMjF6ThNQM04tAGGxMOKHG
Cfw5IAputUS2FA+S+vZbrb/PwlGtQp2cSQzPi6mImYRSm29ZQ7Xaiatutsjyu/Ze
uLqzNOVbzG1oyehxtiTDYJ3oxetLjYWK5TVpkHPRc5XpDSQxj4r0BGauwkSjsCL0
A4Czi3FafAt3DvRRWL5J8bGItjDUVycbLbJVaQlsLUq+ktgl9N8qvYZZUyt//z9R
gkCzqYdcNL9/gigAC2pVjJCC0DcBLavL+GeC7fuNmBhs7Zu1DlFdc/zS5x463jwd
0LsMSYB4cHSY8TWRXVnlY63fEBmmSTShVYLaIxBSMKYuTdbYOQ6rNj/DfiERnmrR
RWsw4dcm4PH6Z441UAD7M6nx8oQynUhk+wUUlaek3UO+QXi8SFTccNUv8CQSWkwc
LO2es8uOfFzWNj9p7SQNoFP28epcvTDch0hxg5TTi5BwMqtPW/DFRilhQ6EAppet
S+xMimWH6nGQCmxbMLr7l3FdaNC6MguA6YipulJJTqBFRWBkCZ1XJEY/sxUrhDRz
HmThI2kQvBMtlFZEApIAA70RVZ3KYGXIlsamV4Sj0rRj4Wqz1g4Zzi0Mkc90GUuq
XEsVI1Jv1HQ0W1CZQkqA2NYlKrHmyun+Yyubu4dWCJoBocki/5Y9sUKAhwIrRQmd
dBPcNj3P9KXmO8lLdYA2xZ7Y/2+er9jJyr0T3oMQ4LnvtEhPK+ZxiZYFmvmtMOf4
aHWR0goi3BB+bBiYPCvlSOPDv5DFK9kBWY39q2mInXvWatN/9euZI9mm4JFjUpKg
k+AklsymAOlRnVSYlH1n1rQiqhkilagXSIPvqHkLKLPnIsEysjn+xB02len6WEmX
h7WdFeed0+8zvqE96R7qm+h7ShSyhwDpaD50qpBv4JgOlnKXu5KStyDM1bF9ZMtJ
YOL71nmYlgFQzq5Nibn1w1PPuJ4hAZB7LIfulou2hGp/PFZj29G8Vx8upJ10/rl3
R9PmzeQHNAIIoN7AqGUFDDqDHn4oXVNldUTFlrMNx7kHF4m7b02ouTqay5ZtFn5/
Zb33Ls5l604SccSbPJ9rqpc1wA+LyMdAanRbDwn/mm6akcJuPRU1n+RpwLUoZY0W
JVK/Cas0dSId9vNq0P1TEwKQvdnH5uvp/1nCL40o8D4fTWMgfaG6dh6JqJDFC01w
s/FwaN+MRMMO0mwOQlSRr+0RAdU+biR2vLnuHrmAyMsRQMXxkkQbV0uL0y9sO677
B+27AuLfzoPsqjO404KoRANJj9/XLMd9sLgBcKgFc5bWbenyddfBuieZb/g5F4Zb
1gl6Au9nhNk5YIz9Z3CDHum7sETneIoOiZJ30/lPl2EnTVhn+fUizAVF1CY0rRwV
NfKe1UaXX6Zm6WaHEhleFXU5nHSz4g8V3EnE+nMt09aW/SK/DvLPFrjKuGK2bqqM
7uD6SZyi6wqpQFJl38+wFS5wxkg9jgyMiLJuvOEd5ZI/sGeHD1gPqZ/Kjhevznk9
aVVzoeFEgF07XD0H41qLiQT8FjsYcdx1z9ydycpNSah6jRYSWOSy142q/QjAy6sl
1/0fivERnJdY/YX+V616xU9Je5tVlPMR9PYbeulPf+V15DSufd+v/uwSB/d1O/t+
H7pY0MjIVGcM1NYwU4KmBKLy1jm+QPkXrjBS1fpaZEnhoolhxhj3MJ19PxOjSokN
dw41WMQYRg7oZt/djmMKqTv+RA2WGlaonwViD47Civ7obbsPCY/kKKAx+/fjPK2m
/BZcWqjW5VLZyHJVm3oY0gVDJsESHz55B4UDGdSg8vMeKjtjmZ9JnVi6hIS8T9+H
d2YeTFjhxhBYom3J2RRDbXd5qa1cTF/4qfUb3XnoH/Om2Mn4WKztNgFC4T5rL62Z
hNhjijuPEsjq1RN9VYuBKWTt5TsSy+EkFK4Gbs9uSPilZzTmmaLMi0s8lBn+0nxH
J5nGNKMx2wKyUvM4TTaVWVHE0Ebvyt4B6ixx8u13grdytGdxwIsNu11U5b/MTCvc
cPb7oF3fUJ3ZXiNfq8yVliih6wNUzLwhiEDMMb7V4kx9FbUuXLjB9S4520rxbf2n
2bwa/vRSFPwosyEokR4pzXPjkP3J6pTXq7oZm0DShca4M6+bWKVyJI4HXiLuGtFE
q82iHMuK1xpAgXLeSyr3iKHsysz67vYjdReV8FLWYaJScmUqiSROLNNG4Jczxedh
i60XVK4LON3nqSQZ99OIuWkCxs0ClFeiNJFweKO8ALYbd09z9Z1PtAIYQkQFl+Sz
tiauPUYlwb7iYkAgmzrbFlrHLkEAOcg6Eu93TcztNJo63jzT+mDA8lCRSFUHiQo9
2WnnT+IbMZSO3xSOw4QLyFJBjZWwqTFo5Jx6VXmNrWOV2bj3+fZ9led3tY3LtxPC
eQ0py+u8G9gOMtnJ1St528wIUfF/oNLnXZPiICIKLw8veQ7t17r6BolW0yIODd40
ChXhZ2C6T4a3cjbe4Qk7eIgpx+tckOez3XK7SxNb/8q9yUCBxgLqDOGRWHQIfMKh
KlvylIqQXIp+MXGqOEy1hUe+rm6KcY+du4LvNJFlr5fHybfxZUrqBsgLuhyssmt9
9YwT0FkWwd+mB6us/xiWb5DY5mXLS+yv1mWvnOAVbeYtBWsUQ4A7l6eKvyw7l9hb
f8/xAIaO4s0Tc1pe7xWM/Zwl+uK8rpkHfcn/osRHAEmTGK32vTxhLfCvT5VaUNOL
mgxTcqK4T+1lkRwnL7cWxvzrpVHYdsCCcHDPYp5SPST7NdQ5aYjR4gOqzANCTWDY
LWjM9HCPnfpo5IERxgDtyqLujO5T3/vZVEy1uVJUnFieG14m/YiKiEEuo2WTpB5X
Mq6mO8T7lKZ7y5CNYqViX6G5S4rGaXE2RjrQ7vXgbUCpnLagZ1ZRhyBBIAeFPLy2
/crENyjDiraO9Uoi1OZ3/BSIetunkimOlqyajCUZ/KbdaU2n8BoInZiE3pC5ZPVo
aJIHjexvyXK+em5X+2TSaj4el5OOaMfURmkNPUnFRCuX2CuCm6buU02FyL4VifmN
M9uviqKlTfd55KbmL8Y4Yw5ejQ+O+uQ6023AzNfZNgMF/iAM9gMLSymBbKZ9fOXA
kK6wsU+jHE0m9jcGQne9MLf5h/jp5I4samgU0Vw2sxs4QUHqiMfyPD/KPKL2Num7
oMYmeGf0UtNvdPMR93D5PIygobrcPubsuc4xmyLdEw7RNiCU5v+iWEdGbOCEv6eH
cHN1s32wBR7LFCEvOrTsU/s7EgM9x6SJjo+AOeyuotk6q2CWKm8YvfnMoOUU8OeD
ogDfUaTMd07yO3NT3sWUmBo7xx0rnX4D8mbYsJrPat909RK563x+q67RBCEiNIED
tfv3dpoar6Bc9TN6SE0ogNTST4Jn2+M28NjY86fBmmt75pYscBwVnctryz58ZaK1
Fs6I3mMFlX5ch3c3ZSY6ChR5NLwCFwWoquT/4UOSf5SiXD1kt7zjT3qy2LXWjxmB
v7qvHeh1jBi50/E6dqHgOGJiliRxQqrivU1IVX75cV0btek82I09KiSI6AY52VP5
Lz8Y2yJGFhWV+u4xOcYrwIs3QhByawrC8/zeIKJePlUJsfh91kNiExxqVqmjqEvF
/5fsf7Q9rlK65cR897psvWuzUFZ7hIpezqdDg98KleR0jsXfgwBD5yHgfbLlOQ0P
Shb8YN7dGLBfXKlq+WLmkNVsaElOZzWuKWaVVN55x7ETauPgkmjpur17SR9YUBia
uuFORHuM0OPbsqediFkdvWUYkWxCIUykuv7yHPryr9pvuZvihmPZU85fOkLDEmSO
hGdU35vHxu7US3IggW6QK/0iSvPgFmaBgEAVirFtT2JrnGdxkL+UWj/x1XhAUmND
37fF4zyGDy+s+zsfoUKwWSrj5ZBS7EgK4m4BXTik3OL/XNQ0gHR16f633A8pwMOB
f/d49LJzaaOnWB5ee7c7DC37vcxasOdg0OVGw0c4NelP1J0T5new0uB3qAtKvDLM
OSzSeuAR3DCyksVeMxu1Ds1L1QjaUUUB1b96wPBl03+eTGsTZSxqiXh24AcsvEUX
ID7wcVAcA917O+PF9dtwxiq6I8zv6iCsuy3+84Jag5WLk8owAz3VymdJC395I2Lh
7/9CcxM9Y+TeA3iU9jc8UDUSPAm13cWVBnXEidQC3qOjjzNtXaTpoLlOspzlqdmv
zlYDQ6rDuxr+bdenQfpDw2dP2j8aohjHbNIu79tDJFErIxggA40hk2L6NZYNvyPs
LRRiHfWCar6cN1cF1DRnPkApgL30XBbSKO5yIKADqTMbUweuPSaNe6QvP89rweS9
4bOtOC6JLdGa/YROYzXrW45n+wslIqU2xV46/7NsDuQJXUmvqMI+juEMwC1phiXg
wTZzGR5E60qc6mZEuEUfLPQTryahpaiDAiBp4HN+xopFE2hnMJbXpQ8w12U8XK3f
XmHcIKoeXcN/78VzO6mbZf1996KEC6aPmVW2D5s40PoXl/tlRlMvwxQEo5/O8Pge
QNc983M/oikmSWz4tssijUyJMHrpdUjymCwrx2FzLH/DGt/zpHapd7O2VhPxwHSA
8K1vTdJBHA5Csf644s74grdBxgnYvhcuVgjfas/cav79qrV6MLFvuFOkrPxEGhkB
CoSNOGrlRNLML0rufigwNzURyvAbMWhVN3nrzVXJ9Bl4Dw7DW2/cchUBEINEeufx
ovKjJKYJl7mDKB6S84A1rQHXrls8DjRcx/vEMzKFS5iHGtxuzadjr6afqEM5cU/P
LXYJco/gvvnAIz2WFkBkAYL+JGd3oa01Y8Ii7bo87j7UNqABy0wqMLB4XlAisoXi
X3/3VpaFp2hgiEM8maszeM/Gzzxo8r+U57iUkhAMLlpIcS91x6ys2ZFnlto36Z0F
6ZkbntBe3nsha8xV8T/WtLRAm7RlmM0Dw0J/8QzcBPeX5cJhmMLmMzLEK1B7QkcG
AzSNKkuNHR06XA/Whv3PI4F1aOsruta31ft06lxUPD/xGg2b10txKlEi8rZ/Kk18
Vx8rxTsf2CqO6TBXmwR6e7PgsWwgsP/zb4tOxb6KeDGmV/XxZLJ1CCvpz6BZmHZa
2JAYbNrKgyIW3MGfO+bQ4k6Co8/emppTFEBYz0zRF48NNWzQjrKtdEpxLBAswYNO
Ix7cK6AQDi3KAYsg2rA8LmAt4dETvoP9A+839qtVWGfciZvrgM9WQgNoNF6rm1zL
ESU6JbVoIRsiKa0ocFbizF8GVMx72hcVhZUasc5wCZ5SEsm0CcBERdDVFOc+M2nX
ErcgM7c2E6sKp0WNWE7EWCcx7wpSTjgCO2DS+TCILub2XvOhxJfT+8uhufvKnjbo
9TS4lwFVP8SQHbzzOs1VpXLnhh1GL4qAo9cA1e+amys3C+Qx6NrlITznlBuqFiC2
k4s8sS0R6Ann+zHWg1d1LwGAje8y9lF7YvYdXwQmnnYgj7YEbywXOvr7wU0pj9fq
s8upQu2cFANhJWX7ufbhwppEDbf6ZQpaE9uxuFuYYKC+QmdfOyS1yvkVxbPUZZOc
Cd0Fy/xKGMac7aEMVnsH3qGO6C0wUsB+6mlZ9p+jb30Ak4Kb0Gdm1HobgF/KffcL
Cr4gr6b+dbJ51dA4rjcFPfKqEl6IncL24WVqP3MxpuX7e8GYZSoRMN/yfwGvQm6o
7AidX0h4rOlt2yjM0esB7zLlVgqWBHlEZNkib283Io/1JbODBblP3CoxYLHdtvL2
eUw2hmHDwLwydlhXT8z7RdBXCn7w9qknjTAFoUbGH4IbudQC0WBXhvSHHLdYaz0R
0o6uMWNmrSCy1k6tgufzb1oacdQnuv6nCjnk+kGpc+ADOH/ytFjySUMKt4eoURp7
fUjOalf9g2KLPjet7W7h6LrLPfwWFGfmYqfcwfPZu4mbFPQAekFrA8CBty2WlGtv
HTxyL7zn+3bQhp9V91MbOk69qnw1gG3ZjGbTahrgFLDQoT/Yhn2hDUIVnZ717C2d
O4ilGAEPtsXtcqnxpZsGXeeSs/3WHW872teQQApnQ1t67FPEWHrt6WB2Tpz1xFNm
V/RQ+NxmtGK9cjFyqsHSRTCJXA68cR1yVSqXbhRp1yb8D20DT9e71XX0hiRoN4wD
lsVy1uVTWFSABAlzvq0xanPqvgDGFecaMLE4VjL+5GTUG8nh4pEcu9Imqzg1ihUq
SAHPOnxXVr2RA1eQtSPp6F6REhVXi9pQefAiPQoUvB09GWUbMyk02Pc4IgvK2r3R
Y2KrX3CHyasjIGROKiKlG6QdxUsTDdF6NP5R8djp5JhtiVF1BFeZ/6rj3Ex5iaE8
DJyh1Rd08hGmDwOmkFn3sziFIpEQcdfMvbV6mFzg5l51UMS0jPgpg82NOpBoU8UP
2EEtnGoCKw9dX5JKgDugrM0zeCm/waLiAAbAIxNCVyfSPH0MVhJhQjj/9OVWcHVD
PGiP5NIs4DCk9Q/Yicexm8iUcbkQdXo7ssrfs3uQvx/ugeX29xMnDsoA0arXPZsk
KRNZ00u+NVEz4aLEQ+B09UPzZjOVINUu8MFYywM26f6Jyiy7ZnwwRR+BImvZMEPB
xWMoghkxul5ps52LxN03qER34Ralmf+K4Wwmqq5CUDo=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
XWV8yK0YjlsQOTaPc/w61sscragbwDHctnrH/miqdPkk2GcqYtsXpneLEHQiSP4O
wCSMRrt/fgdndG0RRT9nq+XIr95kI8DIFm/wALKR41Fel9V6+iwppIAmFv8MmUgc
a/N6l4ox3lE52/5Now9znSIrwJFvGOJlXdqTPugR+mM/ny1Ds0h0Des472WBoOXR
sC1EXHot5EweLY/zOHeqGYjAfIloe8r5Bnxan1+Shc78n1uLD/ZWsHfEWgcNgl+g
RB5l8h9JIrROlxLUAVOzoUddwojmaU3fXH6UY+KRjomOJJUUMcd0NW8DWzOt2q2A
Ct4kXF31zNBppuPjM6KepA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5360 )
`pragma protect data_block
IzSwzlsyrk0+jrEgaPQmrMQvWr1BUidTyHR3m4JyOpgl4JPDfS1dlNzHY0jA49DU
CMUGL3c70UJ0bdimqm/NlBHonzyf84zDzC1HNE7aWTgS/DgjIJPDRuP8bSFUGW9c
Xi0dLQjagYULpS6eRBGffOBC0oodvR1qZ9Iic0AtTJXECnC0rAof2tgzIZw7x/5d
hgKsKRz28ZHrGT6NFq+4PJrTH8wiSPfpUYgFidboA3SApfUN4eEYumn+uA28IyEC
vANeFU3hE4Hw+RJkmdHGDNCWPJNrGhZuVJiHXGBf2Kfm8GDiAXIeg2YCrt2Zx+oA
C1JFeQnfYzX1dGYfc2vMZV5mifaxrc1PIoGrcyNn4fTxtx/TE8/M3xmkfVsZQGXV
vVorJzCNzKBPb0htvHnHYzLMrKT6A3pjyvyKdtlO+p4PyaTGZYVL883Ud14y7HdV
ZQl7BqEZ/JBMoV0EsbatWd1lQEbXao7ZPRzrs5O14+LWhbkm6LfUOX+uDYrzahgC
KsAoFTLPH8WHRtJMCHMFY990km+TmoCZz6gVcb3i0GLK0EIRfK78G1G+0xJoxQWk
g9umMceY37yctBM6BX1JIZKg4aN1z+WiI1NcoNodwqCVr6yOkuyCcmb08+izByCU
u/adfIlfwhnR32zYvt/fO9zdLgLdBEJKDxz/Xo4spc/B6cT70L2XpbycsCZ/rcM2
c8Euyhak7tu3FwtTTdCGNOdOea53p+2BJz9/FWgWhmfKXIrL97HQvmCvvG1/udhp
g08Q5j2JW6KWzcwzdMK/lc2CxLvIse0iB+CzRWWALj/fuT3ddjaUHfXJ8zBRni+E
P2qKVZFvYNSNHh8eUceyjlfAO89P5RGnWK652Wq5kSAgjo4YLeH9hszk6QZ/lAG/
jl6KSeom0eoXYXfipMasWCsjmCdDw7WNsG21jy01fIB1tZ6KwggevrWeJX7xe0QF
5mkH8PY9btkAB9J5vY0tJIvYeS9eSvNbzt0A9WtRatxBSB0ilc30l3YGpvMRDtJK
SXHR886nQrETrzevC0rSsavawpdBsCFYJHpy7MlLQPwzKI7uhnc4RKIZqzhZZcwy
vMKIpiZMtgnfIMTXmJ2pbWQb8HQhRmv9ne+eFhXyRPcAP/7014Ilq8SAxboC/OY0
vkzuaYBKV5LKHrfJ6Yoh3O9AbBfZ2ckL6Swh0xqIBzXkQ2ZfGxRHtSJNNJmvbB5b
pP+R6vaazTBoNByINdhLl68Z0b6CD20/rsfKr82kLWD5B6mG33OzRPDMeFdSZVz9
1d0izVmTUkc1WvTAKA1Cq3aQpEgr5JWO9w31SzYz7cp+7K+f5ED4m2sJ6sjdF15N
lEV3tnuzkGXU1ybE0Zfr6Js5b7FsCvDkCKyDbS72TuOb56fieDR+0xpkv3diSKCt
soMfDcNdqqIvMTabZ5gaMDInHUdbz182fLcKKvIcgsQVtqDsfsdCVJddIZVJHCfv
TK8uQYbdG4NXiQhst1NTr2yoMIT9s5FDHiHmOtT/szcfIo9pyrL1Cd3IiNwdlm/K
p+AmT+2F6QNJ9AsmJarNnLLXfO5a93uxHfv1qq1wi9f1TSBkE8IAONLSZvVtBz/b
NgSuMtB6NPLSOLfCBmWoBn5wA/y9udiLb1j+yNydVwYE8pdZACBwJpUf6Vt1ICZp
iBqG2Xyf4V039ozaHHGjo1DON6wYbssvTm0LcdokVKu72oq8nyO55H0tgSEOEuBK
lJBgCLImMzsdTobvgAcPU4ix2cVOK4Lc6bv1xGwaCfQvkq5Kb+7itNISLdJSdV52
tb4gSmBZsc39SZ9GRlhcUm9rt4OFLxzL5XER7/ndif3WhNYEm+Z88ASYb3Csewp6
l2FXXocU6IERIO9DCpHICDsr9PjxMUDW5F5FZBESfmT2q+JqEUTF6OI/es76JJ19
F0LAzSJpjsFyrX85ovm/2yFJCZnPufdHkCDDhOJAvnB2yN6GXHxlFA40OFoyjA+y
XH4yakZ/oZFf4J7XG9PUcn9VIjhlubA3zGdhKhw+vWpRydRBXXhDxdfQ3Q6buhF5
R2klEHtRRTXLhz4iAOaBqhZ3NSTF1XbvV9dWsOMOB1kuDnuE4t5mGV+3itiekcBN
w17cmNaLxaIswfjMzRynbgicfn03Tt9Ws1i9c3rdHWELV0l+Qw+kAFr/SWxKH3K1
JdJ3hlhzyi+SRt8cELUjjbFZEe2VvGARuUhu2UTYfIlpUibn5l+Jq1XCcIY+vQkz
fXpIH1dQTYTO73m6HQxmg8D6fdhBs7cfeqPK2jMeVFCQ6NmOBPrBijKTpL96cvOj
2ioNDBFhbeA/+/atxVpotfMyaVtI0xtGWbpDinSup/A4n1Yj82wXR2ud8QOoAeEq
cHbLlFMlz5QItOd+3huuyGyni/UOyHH8wg2uP1jCb9Pd/VLmTWtkzfEOWi3eOg+2
lTfKUKfisFIzvj7TW7EyIrUYM4IMfp93f9NQIJMeWswuDmAA1rD9fSmiSbJCRAGg
btQtD7vUTA8iwrCCaBBqLtCb07uGtFUNbAOddigrkhi7FN+MfJMGob/B/HQniNNl
J1i4G2tae8IypKRCXrkM2ZmCivT4VgtXJIBpSV0EfULNmv0442KPjn1ArUO3rOO6
iWUm0c/D0zi8BCgqvu5ctex+sAU0sNJHY4jhaU/sfG2yV+6Q8Due42tZMUfEE2kE
lN9TcN0o4XiD92gad2+IJxZ5Iqs1aLPHbeetiXRvtMiJnM5fGllq6R+ktkI7A8ce
8Auk+axVLvzMZno+8Jb7gQdNLjW2tmYgO9KcUpyc9w8PSd2ZfPkLLZNbWf2LoaE8
ohikE+7zOHv532zfEBfufdHmBivMUmcwM1Y2uW17eD3MW3/w2uzIf3Pf3y4DGF08
u2lmUNMf08rfoG27JU1VvS44jbTjWhel/78z6c0r9bqTTyw7+7faGn2aQPc/ZENw
C5KHbmw+8OmpcwA1p94RbvcRPM0+60g7PW1mxI94c8fZQ099OpmBeZfqDGgzjO3j
g9hIJhfsiq1zJTQ9DtvSq/nwSwMXQPIt5IgLTKv+n6ikTV5RPLZ95R7bowKTgvet
Ws6HUzAM9yKBqwXkQjhxSlpztfniE542lk23ZrwbnbS2tmxSVn/f0sF2yXO7sSV0
B+jHiMo7/iedWc+ZJbmSJzxto15L9vYNvWdXZrH/o+mwtylHYfA7ictQl2MaxaZb
i4Cj9oMg607+QMB5LuSMkaljWvGro7WuPiGSbOkou0SemiUAeGWxh3YTz52uzPsH
rI1WYyBJLgxLLvyxtzCKubqyWE7nFr8nVIwqU9iuQlYsxq19NJvt7i6kE4BDKUfS
8ovYRHkqzUw9ut2OUANNvp4YBXfJJsjk3L3XeQfR8MGCFiazH1S+udhORlS2MJgQ
04sQGJ74fnyDbcek8i74cMMJpOhtmp4979G3EhKeBNVY4p4xnRTGemIWu7dxhRx7
TkqggCrG44XU8O3oEIufhwH5ylCtxb1DGAGHFU/6idWVifO3P8jOThhSfycXCRjB
jEx4dBrbTSMranbLRkP2teSo6HHD8joz/XlapqQCkEzPwJwDO7id9glAa2rLhhZD
0f5FqdYHl9GHb8vz/UC7qHopX2FjQa7wOyGMMjWqzmUVm/iICnOgA5x+m2eZqeGX
Xw+lbrbCz8GRLCqWbC8HoZbhijXoyGb4Jhlis1taD2bi/H0D6Xqfc+uY65hnzhOV
Is5hGTpKPp1rzRzdSnrPu1ekIjYat4IWJ0YAoyXZO8NIfwtMq3LD6TshzVdqM7Xx
ZR2NARNw7+rFJr9f/VnQ6vaEOwQw7ic14iE4wpcw/4J30x4nOoxcNa0bcXmQLTHd
zJpmpz0b2hRI6j34jxLPv0MJYZ7dY86mK4sq2OAnR4FsIU2E54yg99DDkjUsfLBz
iXPrAqZL2arib3kNHUz/nfCB/ij8YeH+OYpYekhM+8ZfNIqwmN5SJjWIQm0/z6M/
SD7daa6hrBQUlpK+mUFRfnDHNYCx2+uFbWujqmoU5bO+KknjY4RvntPJgVnULKBD
ApPSdMdKd9ky6dWJOitJNUstfBESEG289iFRPMIomJFsAMMmK7lhqIBT4iAlwGUv
uP3i2bmc9xoc1aqasWX0P+LKWlf8Ljs2nJ2AJSDyKdQmm6xt2hxehfk6APG5OeNU
lYBsFfdA6hPGSp4pMS7Hd9Hs42GTO0FOr7u/5t7cDRe0OMfCKG4Hjn6U4AIim3TE
3Edik6JWwozqvo3LcUKZDcoQyAvF9Mwrrvtkaqy+ZhN4Vd2WOC7TJnwJ/WBTAfQ+
DQ/UNYAN+E0UmCCZjugCu7OhcTxgGPK8IJv2UJ+ZGMvJmZ5f63nTTpoDVKfL91S3
t3zrszQ/E0YfTK4uPIiHyXf/xY+7mpTtZJB39xm9pqJvGSgIGXCWKDpE7Z3/M82w
YjuRA/WrAh1gcKGlNCRjEPvmvhPsSIqVlZ26fAxYbahDt9OfnqGo27rYbsdRuzrS
5o1i9/ZAhGIhhck0fCGomybUdJm3JCSU+ovj1AeXLif2ezRVkRi73EpKO+xyWAL9
NWGViTeMQJBFTNAPU8RX40BaaU0kUynGf7hGW5v59admZcZ9kgATdwuModxETBto
UzqJYiSrZsPY6blTtXSmRQWVgtE7DzcBBbxdlZEkHBGH86BaqXD1GOo7TAKlv7bW
knho6zuPs2l+QCvkNJc+17DVqPdwj/sTYEC+93sqnWk/sZM/0rZ4jhbRLygwUSsX
TZhikkmITXEmnPV8JrLJ90HxnJQTtAV/TC72ts/yccJkfusdo7uY0a6PGWfJ/YPU
1/xUJeD0miUZZY8fNSo6BKGogjvguP9j+p8shNzxYuXM9V3wA+0gvjC1L8kwSwjQ
Fengtu3C5tUAijM9eThdJjyTR67OzW4rd/BUxdFQAnTWDK23AobATKRTPt0qKi+u
c9V9pc9O78RYr86DZgWLdAMFShI4rKP+NO3lLBzJ1xtFX0/kMJkApTQ81vlxY4ko
5NjnwoGS+eG2dN6CVUToFe9ootDCk8VPvatYLuo0qGwWRD97ZJbYlxxxakqRwPR/
8FwdbE46lZnLgbauDlZacC0aLrZLxZbzYimGSOAmgtY8eDcM4nVXDEUJKroMF0lf
kL1tHKT2cpK7qVGQR5mAR972cndYb6uUxW4prSEX5B0946rbwzH5+llFfD+FZbNo
AexIH//dZmaiDz/+lEfjkgA03lY4KcChE+Zu9AGaVGkNLCIKzfaI24b/0n3imSfs
HTQTGdWbDLtP7phLuYLiB6XLzDsv+oSaE98nFwMPdSATyahWE5XX51hPANOMiR35
j4qyqWIG72FYfxsdn2YIsdidgv3DXMS+YmEDcjzMtrPU0rGyRtP7rTlFtH6fs1cx
R8YuFYtjArRiy4+Y2JSwXIjxo4kxg/4jvlMc9yeOa0Vd0QAPCAquL7eZqZKtNszV
1/9D9IsWIII97AtyqcVaekIO+giDa+/8lQF/PwjAAWMyqXMgGCdIG79x0mWpUBsY
eG96EzrCue98adI1jAdxoarf1oTgvyauEIj++5M3UI3gNcbQaZRzvsPDSGxfzT5+
sRs8s5Hznw8QA/ZZ2W4MoU30AG55aSIDCTtieYcQi8u/+sU2cnb6hJ035T6Z3cZ4
5pD5zQjQIEPTjdwTUgD4PB7qXkT5UZOKcWsD8Du7zdTjD5ia8Dig566/K90UQHyX
/uSsAO8LEVKuLdaKYJ2RJkPfAURepfUJSNtb6E3+q80r+q5XuvpUkKmkn84Ri6Nx
MRYZ0fBIAoc5+fLTk5xfBeDOCJVeHyRxiwQdMqlFBpmycSZH5ps3ToVXDdAbvpQE
LDoMcZqNWo2BPenEjNr3ZWsNdwSojoqVuI2ZOtJTZ1GjISbZ2hYbo1lYvXRsc0/6
kDUCwxQDTyOmWc1BmnE1EHprbRbEOkoqau90dpQEkVvajc05lftyqJhyR1rI0DwS
tIkn/DOYx3AtAaHMjxBBwUSH9uYxaiYdG4fU2o6Ep3k6GKLkBKhYhbaTINdp5MhX
wm2Gd32+Anb3nSrE7VDLZgcYIcvFtVsUU3wY/2+O3oqvevAzuTPmLndBhTHv5Swr
af1kY3fCSZAxFm1RfBLXFoaSPq9ug2f0dl3c5nzyA9X9SpuCbnWxwRY7NeFisf7W
Nq5YokVVrAnCDfDkqxy0XxjxVz4xyfV9qxx97VGopuRmjHUp8T1KnxN4xtYvhVYb
nCzzoOfK01/7RPCQqi10XsNws8MRnLemzX/ujLmtiX5JnOv02+pkGA3Ct/aFDR/N
wrHOlGS1OIpz2SWFDmuEG4Dfdi7qyKu5q9sZKQrYiXirFagEpHreuEIOBdbhL298
70AfUMBN9JwSMa8oEiwuXLXkqPkv41kIHWhhl6IzoJoTTEyOJaMPMCRpPxkpBETS
OLgRpJaNgDGVNOowDHX3NRCYc9xSJ4CQWQqgYVLZg2eZH+tkMYtkFlz73a19V7rw
AG7G31+k7aNu2Sc6nLL9k38W82mxbs1CqJpZENOCCSgd7K+hj1rz+WnzdX4ynnRs
z5rnwtR1hqG1mStXayerD4J6BvT30hn8TAELzsp9Hb5PWy8LQnxdFzGFJxUFicKY
E/nyqz6nQrv+f7pturzBQ2h09hYuz4yPojm+owq34N+AegQ6kmzM8fENbr1a506l
TpofguHZl1mZSaqCYtDhuLrDW+ApUxmO1/GixuHaO+XBX5BVr7Mmt5e0RbD8XxWr
Iz8qL9OaKcj5l5lx4ag62V6UkabvPoCn2vkh483xinLEPpGChy/pjZ6eZQFMBOgp
GW5kJX++n9TnzpVNUk96aA8ZK9CABOKvZORHSNl/B77W0UWJXUXz40ExrLmfnT3A
JTJMdVEBfRiyKKtjtUOV4gqXiRFL1pRNHnWhHHlF/KxMNlSxNVFwlrvb1wend5aI
oeBhE6xtJRUL00LnMnOCNDiCxLKRpMovlr2sXJKx9ElhVIeY3gBmyVuPduYHRyom
pe84tLvMbIHydvgelZMyxpvKgHIMhA6JWmelE+M8J8Esk3XQkgrqlgaus/a/Zga0
u+ZmzoARL4nsgP+CwsJWA1HQFbJkf221BmzJumqpEFMq/SVHd5RrcLcY8dbC39pM
gatiHeSxC5Cf82/AcPZlc8z/fZy5rkLIQaE/drHIxE4=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cE2oRtHuSb7yFLVebdaDJuh5QoesMSFkZo7v96BD9za/tzyJsnh+3T0vOJ5R+LHi
RdUnYXMBeJ9+hN0up/brHaawi+M4skNl71iLS82X5i2tA+MvUWKBlBd83IskP7GE
RTc31TWkePxKd1oO6HYX8X/jO8ZObbPrLz8UyIulWLSGZgoej+T3jZ30JG0JGiKC
BK9HvX2NCUrkGXcGV76zQq7jXF/adkAttUOAtHAPgyKHWu02Cbg/F9L2dLzgTaNG
J9n57G0ZTOKLrkSKKqPcT9JKF2vXQOY4FEJAwQJSjE2bHexT26SB1X41OX7iNL2H
rzEeaJqrUTcifWT1CI1AzQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5904 )
`pragma protect data_block
s8M7hgxbx78v4+bMnsRSGYE0HYXyLv3IWEHaQvKbxqJqt7BPD7eO+DJwsMVVQrmI
8lDyaGdm4mNQGU2YjBezRLsje5orh/dx4cw2hTcPc7aytn2KnckBrhyNGVp2Q9ZQ
kkodBL5u4vLzJNOcG1fwI6l5UA7VVRyPkLivSUDHs7FozWglRlfVX2foF00bLO6O
A6CtFUIZbnKD7BeRAdy/6XX4J5+zSXeVGmSHQCAo0e+iGodsj38FeV0wLfVoxQkY
6Trhu89X5zXyM9BEAQetio6elN4z4NUd21kXX0SknQy7LpkyAgTuNhSFmAMOLmD9
tDDfFMmohetken0O+DM3YL9ItblfIcf5SY6T+lnM5ZFA3i+qZjR1OHwq5m9fwLHa
0Z+iiTQiyLsa31cFpwXO/QVpj2b71v+ECXE59+yZjbpbtfrFYcF1WsrtsCBJlmHs
6AZ8ILM6KAKp963KyJngOf5W99jfQV2I5i8JvQTj238L/JdL+jwU7j5MAOVbvZNA
VbI0iUddaghvFOiKq3dA2W/c26CG1scyW4Qbo7Kuopw7toMcnqTlrMqbgY9+JOqs
ZvVLKaUoVHNyysNmRYkWRHF7Ql2GehgXfyS39P8xDqAfiKDuglgfAkCW0jeivN4h
WaHMWX13lnx+Vswb0oOL8MKSP57P2sKLdX6XUU7z3MGuIwkZ+uhZC9sDFxzxZ2bH
+wwpMBG6QuVvEIqOqPR8hQCHLLYxNccBWulINku3gEGYi0hSPRY4wcUDtVTOVWQd
XpTHl7x2SsCuXHjnLBfWMOH/+OLzjgp60SkuvvIMIaNfhnAaBXMYWSZ7MlOEA+QO
dyuR4UuOJNksknVPeePH93MKlOc9XFBQAuQGo137zQuwA7tUmVN1hrEbZAtDVr/M
xZhjkyL0vFkwv3RLvPGZiRzkUuR1aBu3QE8dXkkqZN5ip3PasCwLK2cQ+MT87s1s
P4uvMJm097wkPFcqpEYy6f/PyHTOr0tE1+qGCxuf/aWme9unttW+U+vme6tfxmW6
U3ZmlhHW7wG6VEemPlvM+ggP2uxQUGGCMHd0tpjTRkJpmS6oQ8G+NhkQdYWXojv1
87LTyC2tCQpBSSIgFZ45tvmmoeOLJZAiixwHPFdQkOPT6E+6MFoDqzZ/evBNX7Ae
ES+6aY+UEqy0i1a6flYALMETv5jF5G9oDZPzQ2McPtriaN/zsSIz/a0xxuHDIwuw
MkDEEvWFlP2zLj48EMm3wtmsnVu5sonqE9kzhnhNkbfW1j+v72hFy8FHnoKhagWw
Zq2txsPX72tLttZGBEA23e9nhNGrI+Boouik3YYL3bnroZnv7RELYrZyk5tuRp/v
avig0GrgeeK564PV4m8RABLj7HQJ7llEksFShDvq7T26MF+r43ICPRPUopOfhDG9
mTj93Sk+LfOiIb7QtjvlPGFSjTTZN4rmHk+0xJB26sntqzEV7iQK0adBXJl7z/bx
Wha6wiZ9LEJr6zYzATKAJ5GhEvybtKqDz6+dSfge4w8HLJGvIfIB69c6oxT6HUye
ZHoUZD7R7aXOwZa23rXgCjIP9+o/P99KrVPbyEnQMFxwW+xIY01sZ1Tv8tvgkHXe
VYYoc8h926biu9nHqn13LKr0CiTlqvlBEYGMr/18OyFzbMlBQtibPTUWNuuGal6u
GqZjtZkTR9L+NmxkJGnIqNsuaIgnG8nRfEaNctqJy73oY+r0JuozKrLqXXFass66
3no/FoK2Y10Zrd2tpsB/1TMnc7cnmtf68cXM7xeRPzgoOZcyhFR1R65PFB197LTV
jlJLAPAmXiLftyas9DkMD063MUSRQPG6dJ1ALJaWEchAW1QuZve9l/aVq60Lww+W
6Bmxb5It7jLlccbPcrjgS+MbQ3D8oUkLFcp40zvugiEldmietC7RWfyl6elnjEzU
SXMcQi+0S/JMCe3l6mROqctz5Obg7Ugq/qwNVorxlfvPbpTckesd0s0dCBw0+kJ8
8DuoNq2gMsUzHh6HyIcFcRmMMNOLOvQFraXAWTzVN+Rwcyx5JnoRXlOsOtY+DbRz
4rjH43VFuSiBxcqOe09JyTN+xzdyedYAP3ZELWNmB0AhUatoP4y5D2yOHrbfJy5Z
jFBwFvZwxup2KGDq8pesAfGKNIKqVj58KRxgPoY0UZZmrlQzn/Kgtv6b6f6Ysw7r
iBTlBrozTgMmmUXHD5tc/kvtz30aPm9jOMbJtMtoa7OFFXsxeqvXLVgqEeQyyqk1
ULCYOqjofN8gXKk8gheAsSDwJ2ti/hz7EJqcyx+rUROdZx5gTk4ZdJZ4l+gN7iCH
zx6H0/RHAASQDY0cOHmB74Nse1B60o8lO9OziORJb3gV6XEXByyUyV1JvYtjOZTx
r1vUuu4b9QMBNQEFpuHS/ks6V8n3cLQVjG89x05kqnbO9sg2LFIwDEKIYv1OHb3v
aWTgtxncTDUOHK5fYIyhTNX9NKuAFbk76WUDpxIuCa7IWDMqhWDfuKyj2YNfZr2P
Yzy35a3WkOiNDcGQyp/JM09MApG6QSa+2zeSxV5/MLYj6XS2RZqZHfGoHvUaCpC+
3qqDGGhqhIDO7zi8+2FE0TTpKXRymbofv0N3bFY/+r6FrO9gK8cjpiaakcy/UHvQ
tkLb6Hql1Xts3f6wNhXSltqX7XDWfqnKbmQ0m+ffAozGleGLgGLpeUHRzHuTRdOT
tpJzkrqCi96DnNCHTMxz0KBB1Q+1NeDlnAGT7pgUBkbguH09MMrRBQep79PX6QBV
jv5SOwyUgyU/K5pqmPMrCzFLroaD2+WJYmV+60/7Xw5LLifnzOQo4Kb94UefH6fF
ooUiTCRbJjzSCjHtVeMMK5jhtNnzRyS3DY6fb6BHQb+GrmbP3GynOb1pAzUcdXVl
BDBUd0AL/Q2aV+PYDJ4Xz91oANe5jeniTPXKHc+1+PRaOppjo0OgTiMTZQ4VsNBq
EJJ8kFtGnhmAlVGDATtQtdsNlKyFLVBqOt9dqK+VxN+2XMqZPWAnmBFjRYwyr3+A
HGbk2lsl9S4bj89z2yYdWdXdd+/TDYrxws4nXwzgDVV0QP3TwSotg7xqelWnuQ+r
7rzwweNxcrbRbO1ajRkCHuG8woTz6HjRcuEcE83KAFASrKeAC7DJ9CciHk+ErK4Q
umIt8bE/FpOmrz2pRUHjg6o6h+SQ+zOno4DBEIDJ7AaJTxoarqHpS6B8VBDLZQ3N
phxr047cjDMyzsNnOrsWyB8iHokXBzvbFSTUCwlvq9LCzbA2dDLJ+1iphnBPk+aS
cTRPKjrB/Vrf1tGge8eZsUo8ZTnsEXVdWqMxRCRC9WLB5qc/CAK4e3a3zsOptBDe
Sz+2M1dwIIA1tz27nVt0AiXwH7EjOmNfJ0i+jjreKdWJS4FYIbg1U8R6+PPqA/Mi
almMRBnZZjrLdfvDnYkuTHJSdugAjEQSxhmbuUE8ylApUMNk5L4eTAdigFY/7D4g
mTbMfPGhM1I7235Wwm49Ay8CkqOvWPCzXJBdiIJs3oQ5tWw3sRo/LFY4KfOw/r/3
4vYQ5ja9evyQCtij5aHWcRdIgDsOMfUmk3b1Mk0ZwWRynL3r7WvWX++G9skqS37+
DJacKdDPLZIlFxWb/awP6U07V/B0HEwNiIgv+zqVciW5IOJsRkKYzxrrHSX5NCYb
ZaxwXzICg68Ha/d8pGno6fY90uZff85zXbmURopbpHs4qsUIBgIXEeUDlCu6dPtp
WZjmk47OvzCD8Y7JB/d1/86b/o3fdcomshqiiD2GlZtXDqdrJauh2L/sTRaf/PY3
I/hB2BvL/Vvowf0rl2yzK9h3116R7NvMHwjvsWZPjkAwJQiStG4G1KhDGAtDOgAQ
lxc1Jx7m3iYp0e4hrij5bmwJHIpzgDXTn9JxR7ihW+oce8WxYjoS6KQh6bRCqhKh
RaOT2Y5lY4J9b3Qb/z8A4n2hygK1i0FyhQvefJgpkORhCJK0NjHB6n6Q+NsvCJiL
cxNktOkhexHJMWeJByloPltIHPgeF0INlQFnmKhHCXKEPhXhvuCB/lCJw9F2R/jM
KnvC9R5n55zVB9RyxmHA3UV94XU1MTkicJMISkxwwZXHd/Dy2GYEAGrkB1CQhy3e
Lp+Bjviw+dzcV0Hcms5msbK8dVrymVAAHmTCFCtB7APwdE6NBK2Z6jrVmB+EYj6y
D9OdoTMknpfBZoULx9+TzgnX47AsBh0cA60H/vYM6rVwI/ZMWfJX1uDdvA3/KbNw
3l9utkMB7hStlHpVhok6ggLPrrGoxEl+oKU7nRGtv/+anNv1dubA4yJZA8YmjDRy
3ydbMYEkICO9vDxvUmktHzkD0/AvL0DI7dOLWGKcLxUQM5SBZpcLr15jtxACStMi
FbNb099WNyhpyYqK9SzdOA+h0g0P9l30eWqEwcQVZUXkl5zCTDacjqjLYNnRcTSe
5F7+usZNFQRZop9i8fjGk3oMTzF5wyfTulWZgSC22lhROEUDnZkKVsD2DR/4CntS
73HwCapKaYbIZsB2GdSXLSlSMw8AzQrW7Qqc0zhuKvdRMdRqopESpHlWIv3FEW73
r6yF3fKfQsuDAX8l3OC6lmiZxR3qtxf6wy5Bxg7xkUOvnO9GymID6p61rVYGY9As
msZvh9eGMpV/oGxhTjnx3JXsm2v/vEhTlKkamrakcWapm4mJ8EBt2ihzHkl6xXTd
kSCI63CCCg917YdQThFWsrxEqeIRvCcYZU2lwMCPi5mcmVLkiA5/I2VSPEVUkvdP
sXD/PTh2bKpGbqhYixEFOc6eyQ7ETjRYogFT6/9muF74QRBgQRypoWVGiRXKkGAG
XihrSG/Xht1FPHkHQTQgNYP1juArJE83XFv+cEb1JZcxTxL2w0rQVAlo61wYzioq
mx5OlxUNgHnbam6Y/Ua6ft9E8DpEIHIXhQel68FcKR5hKAd6yukaW7AsnnxxXd4u
Wk86Wxm2eIK6IzCQg2Cvr3d7wgqFV4fbgzp22cXrpULqSjeoYlUNn+WZ0w66NSRE
9fMsRNXmS4dRLxaikaX5n2Mg9yCSynXZfBe7t0uBu6xJmBl0NQw9Fk+CaM9E/NqA
jOhWZs1I/Q0222td7ITylRV7ejNkIWgATRVUeqWnJdYmIfIpj/ULiPvhoPDhUor6
x9vh/BdPgwxIvslGlsHucCKeCA2ZfDLmxGbz2RuiVVkEEIeDVKqgJ/gcEBgXrcef
Yzp1tRd+uN65t5++0k84ZRzpuQcUPIYg4vp6ixFx7D/mqCVPF3tYXZWGNn1z4NDx
0IYLbf+sGPIFQoh3UpgKAEkgnZ0p+Rg0emuABrI3JqWSkrXV8Ogy0ZnDvTo6fORj
0z7Hy5n8uFKbYTSjs1XXeczJ/Nh5daZPpQYikTzXi7R0WJhnYV9qtVBharfCJIHk
Vbvc/GQ63zUKBqzyOYZ2it/RFq3b6pOSwAhCX8wHwNWsKhtQvR1tnPjWnQsARw2e
/5gKYAQ7K4qgOSzBk6C1/d9q2UMuppDnLsN0+UE2II0/sdA/SJN2BFfafDFSvkXi
/fs/7Cwgmq2GYpUx32eJL7A7O3Z4sArJ9kwV6CXn3mFneRDp35SyZptdmI6ttG4S
leNIzS1A5DzwgU1mbWOMkZ93ZE/Iefrfyyr/62qlWJWRorqS+vX7GzyhKdRTK5/S
/vWs4ZS4XvfIl/MmwlXtYQnEeP0J90HNvtJty+6TDclHK0OYQZEfqZdcC04JApcc
GucFNvuEG9vmS8qwcpyIfhxKEJ8pbReKA3TC4UW1nfSLvI7DXYxUiZxkQ6SIaDeP
S8wfdFybJWh0LbBJ3SZzVRtu+zAJdcsFd/ArTz4YjmFgKUQkShf4MLhPG43tNpLY
sdQfae9lrpi3db0iKqAA0pijy6mDbKbnQxUARG/mB2CCojGzYe4YFmDji9Kw7I1h
2ctxQxBjlKm6v4phmEnF6Q3roxTt24AFxnMyKVY9oSQ9ycjHkik4xFQmydXprGox
+81WxhCGdZP+RXADLzZS+TiVNOBvPm+Gb5CNQ8qkv5Z2Tqd86I0TvDX5CGoxs/2t
m33Eq2pdQ1L6ksTLVS9mOwhYU8d0Bvx8sP0ODMtFC5HQ2BxRHDKB4jXbfi9VBVlD
p9xVpUKcLHniGAAv2Yb/TRvLw6N3lcU21Kt1aODmkSRe8aZve3OS60SpVoNpWWv/
7vd4/bN2zOBJbAHK8k7w/vJJ7Y60+2cxMRIpZYauTpq586hUpU1MZKOtp/yJYE/J
97qPMDvSrPsFORTwoUctIPUQiUAo4OlGqf7RQn3TckGV8l3r2t8K8el2sMy/RkqQ
K/SWIfzxwCT/Y38xbvczpQI2c0os8mbBDJXf9HnhNs36ABEXfGrsrbmPoTDadPfJ
vWWko44i041YVqQwaIfd2MfSSgAygXdw67UAr+CqvgkK3UA7myHKGNHh31mNGlg+
gDsLbGsRZmuIw5R+y34tqK48nEbCUd2+Y5wjkaZhjsG8TwK5p8Pv7lbabTzqoiuy
jzP7us+AhtRW+FzC38NeGVfceMvQ3OCeyEp0FTFc062JWcDfBhXwRoCbKLOEOp9l
OkAR87eN18v9pq07djxMSsNlTFVrK3A1dXxXZe9bei9KMytyExBw1YVjAc6Jv7Ei
qrEtM47y2lZ+UrPB6bpfMmj0z64oVbpMnKpS+BHAPoDHNJaJo6vTxsgAPcc3d6Kw
Q+Y8PGdxd9iPzbxG/ktfB2BAKBZ5XVQKjUExvhpxV1qqZ6qHvoBMmAoAGhYvraeV
noJuxXJ5rxj6HZN542etkgYiUzz6Ymxn4guPqBU+4BA9Vy1w4mZOvo8dqRyPNFNc
1jPFB2SJjNoknW6EHKHm3BqzvEeUWChSnrN2BemYz/l6kcooZ5UxTGTty+Q9e2Cw
2bTj3YIrdMjzE26s5BZMk39lZtOZOdQaRVW8dOy0pOZd9izFIK2JYF73tIfQ9FxH
OPts9cBSFiKJ7YjCDoLd9UUnkCsLtcrtZcLrtX7MhORW6vcQFsJYE5jiv5parbvO
96RjQO1/91UZiwgbkkHQyun8uwZAYwk80LLd4uxT/ctUtly/RRQl8Gv9WLVCRmsZ
9fdkEjDJVFuB+HifdtwgReNSYTT85Gf477sULM+rmf+KuDRWReFUXkmBjg6pXxs5
ugAUfXC3vV0o0/RhKKWiS55ZeLlMRv1QIun0dT+06M/i/2/VT/Iz52cEtSZh4OPW
cEKYBp63KkfmymAOUFmXg2k0jLzvMpOUZ1tYb2IGYgFQcMOG7WVnAl41DP0oCCSs
dCrZJCGRyHjctL87VUitkB2EVk0Ta9sVaLm471DMQqU+1JhekOYBTxaeJ8Kh8KOB
G7MdXS84czXyfFUmHcQ4tl7a1wGnq5rzy3FVuik+yNw7SPTVxgVegbpHJecNLfge
G/5KTBGursG8DCX3IAmPFb8EsJKcmWCTmVbn/Q8fkUbXaOkqCZ+UhvKqITTzp1Z9
549XGNegBdZOJ5VI+/CNk+l7tyVyiXBKkWf8vgwYT2GuQZ662cVI7I8vuFbDln3z
i1tJfsd/9RxWcBmzgbJiKA7wGxkyz3pDtTEXWYYsFM0XHcG+YXbBI7QRFaYTqjFU
/CYRzp973vdCik+XQpi9rIHqzeqhYmxAnfMjmeKzuBUGG2mxvARd1w8zHnqir05B
3EFTCKYW8Oz0Il03hqVDmlekj0hx1ejvaUZNaaFXfMRoLXtB/uA9wb9l52/1NBc0
YRI+Hk4a10w66MEtt4fvugXhLao9SAycXSCHdn9ZVlz+Z+njvWs8JlOXL6QzzbtH
TcKPnfi+BWq0jSZCeHt0auFAVC0vEmxLKR4a1MUtphuxOEXl1pEO5fBMjpFQOt2A
F/rII8ty5RlYxKfxoU7v/4kO7a1bpAO9rfGlT4cEl+eMJsf3ZXdOl9wdck77ccfn
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
oAJTKcTcJ9ktq+u5DGxn9W0qchgqxtecxNbbG15DgeYRz8H7CyW9u/3wfdBNBqQf
E+rAp1eSV58YSUcgZMMFLy5mF6HdLe1j6rIu9ycIkDeJNmimVoYovH51UByJw++D
j06gY261mYIwhxGTaABbfvwGpekE0sQ/C4fOix4JkOWsw6ltEq8640aiCQctlxSM
y3aUbXAKPNi25sOtjDikZ8fC0cqSQqBZRWelqqV5hXHdvh2UuvbdryEhYIB/CiHh
/YYuvKLPeHWVUIXAmwda0Q5SxqN84Ujmc4Y5xia83Z0h4Dj0+OssblBD+t2n8gGq
AVDBSZMMxi4yQI5azGlvSQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7648 )
`pragma protect data_block
/X8gJQnH6VAZUXA8ZEpu7tw4AQeiQ3pF928J9O+dxdXsQjhZIC7HI4nOiY5VeLbV
SStTffUq07PLFu6eD3Vxt9d/+L/imytRYn5AlP/6DzgBGHi63FHZqQpE4QGPfBMG
SJkfpS/cRW/F611+fTTpC9LGuHJBdgpVpuLZIOMzjmDFmfPCDDKgsqw43eXuBmp3
7u1NxWaZtBfgsVMnPAIUWPWqFI0is164l80o7PCZss1c9qqQ1heFobgLICVg4tbv
WISOD8vuglFqtBI7O2DGUpcwc98ohEMc6rV2urwodYSuA/zBtbuHEO0SeVTZ1qEo
SYzrqRQQBnYh7qotEjCw6WAGfUqGJA3AVOETO02pcP9QZfNYkkGkziVztNe8fTBx
Zc7+b/aLjfK2gY3DZAv+JiBQPROEpJqyJNAo3cnlVqCqPViI8CISB66ngJj+mlrE
qWjjrehhCZQFovQVN/N2qjzsWQ+wRFhGmunb9UCTgWBmX6J0x22HxkORffPp2mKn
Af4sNw10iw1AyILOLlIiNs3I+lbzDicRdHUZ+VMin7eZDuo45amtKDkWPLwAixFG
CTw/81Xw4U4g0Uu0pNibc7H0Qjoqk9AIN2E5IkH9RMYiMbBwzMCK5SZQ6Byg5ee/
hfmo5x4LYTjQ0R6tdHgLHTDNq7shU7KIV9pEsqGgK3bjesleHX1xp/5K42NJsRKr
p6okyji+kkU/mKD9PG0y1LxIX9Zh1bQyWB4Z7LFCqBa+AJ7BMszPsjv1+wSwX//0
RU8g8w39+L12V3mI1yKSxOf+OqTLjcofzzJ/XU/++LNsVNI3uodwdudeytUWB80y
E39RzLIxSK0n0V7OcxsJcP+NFxPYAiU622quNr2sK76KDf3gj4D5rJg4NN/DrEU0
secAUaiAnFy07JJt0VI2w9UHFdmaRichD8c0QXjqnmQykN+ZRw/Om21BHrLqr6r7
mhzza9n/EvTNIRKlMSe3zULavcUKT+N7HB6Dd+Hus6f9l0Q5Xf+CcUVuMWeOm1ly
QyBlybcS8PjH3zdrJSe8EYUuiOS5yFmW0iDYLht63NmzmtGdp7LLeOEGhRxDsa36
9R0zGOLShQGKb2YXXXZgtSEPxNH171gPajkgfBN7R09BPW4HnbNJPEEOvwYCOVqJ
Ukf6Fh5Hrr+Qv4FieaSZPaj57pdBRp+Ro0M9wZqg7cVUoNAd1NDVuWoDLbpPMMqR
CjecRVOzZ2EUOtADJGyP6eH5GHjzLaYfHVJGxHV/2SxWn26X3UvrAR2x8OW9M6R7
4xs0uXXKwh2JGCRoYPTGEVD8Mi+1b0SqIBNYyboVxvD5mbutiRLGdo8ueSCEaXku
YZlC1uK4y1hc1KfFiN7ZLeJC4jaNmMVoJoJW7SEdyJM5p7A47TgThtt2fuW1ZAgB
2owg+GuG7kV/BU2WgyKMf4W1gM4zmDvplKyMlwXpVrp/8pG8cWYP8DPhHlumhFbh
7dCup7a7r7OtEt3oAsVSsSjJvIO5EbbED75RCJZtdwcPnKQQjXXAP1PL+U1IBvf6
iTH2Bzt7ah7EYOKe0Y20f28OcDG+KxE1YdGOJJEgNs3NlRLrN1XGjTOvuK1wpoow
d0nVQJS6CmRcfsbCa4GiJcf0oZeqkKrgXiFMxtn6ST80GQY5uZILTYWfYOrfcoX6
HNj6E7Ybsjiq1F3IFbrTnYMn3xam5CNwv8/8uAEgP9HNBp9vWCEgvmOjJ3kzwwU4
m0KJrWVlH/Tfew81jwpcVvsy1REvEQvIbPubAqnfj8PBDsT4D1L6OW8lTCur9Y0h
BUD7OWvA+31riWsocvKjgqvA6gMcN0ZBCn2hewqEFo+sIRW9IT0UNgaHmcAg08Ic
Dy1PVEHXZzLNkYopnZTrZw2L1J/CMpAr9dsUNElNNPRpfGBXqFRvtHOtb4kHKbh9
SbWdAvMm/aMF5dPdB3EAyrVEhN+Vy1MYJ36WjKVZXiTO+M32x5Eu4LZiJ7/ws1WI
4WCEOK5aQk9uBMH+PbVUndqBwwOoYVXFp42P0pTwNnYtfm4VP5/721UzPbHlPJZs
Db2B1Ad2TKsYyID5+/nLwjf6HinUE+40ysmcoMi6709LuWSwlgVWd5XJ0c1X9RZM
G9MZDvyG/PrEj1xYqNIDowUrqx8uZo3+jVlJ+rAltU+UODZaBIidGWB5Gc8NrVub
e4QHH8F25zrlbdtFEtfA+ulNvat/fiTr6jKs+RoiWq7oMOkhtxqfsIT5qGVv/NXp
Di7afR6IwdsN9sbn+BDRTrfVm9oKmr0VbpgCNkkgPsrTyUpBfwBY9kFzgynn5F4+
hV+HaK8Zrgw800l1WSMg2a9JbrpAZLmt1MYtZmzi+oRfH+bZBNTWjqY21fJzPURz
nURM1uNRSNuxQwWtlQrNPNtpR6MWAnarREfmWySuoVVVSVw7huSk7fY4o9282RJZ
+1bRbs1YMjlFRIqqyy9Tw4XV1t+KASDbtiPXz1ANB2zDibVzyuKhDw28WFmKyVNm
2qcs8owsSjPuoiy+HXX6o246YjPitZqkYDBehqySTkWInMy1thyXc9GAfi5ew1sj
iRlM5g08l1e+M1BG7XrEe2Cg+nNGF0OLHCq/VeSSOsWVNo/UQvkky315Q+UBnfsB
TyDyJIJvgAYKXaNW/ITPix86XkVG6fvGtS628HZjeIPLmGWwPTjUWlZOXj305RFF
8UELRJ/G4qDjk/EUoymC12LUzjyRlTVEXR0Ul+5NALsMCmtejr1TNtCVVqyzZcEq
adtr88prkYy378DLDzzV2W8OrgdlYG+McYfjN88ed4y/RTtBvq85isMqBqvWGNNG
2hIZMNfZYhDC39yPh6T3wgT7mgvIZdwfqX2aIoPCLWN5f+V5ilunHxE1UKnvteSB
UzCcN4ybRM+Lz31emtGKuXus9AI0x518yZq2qiFSGRmSxsuuh9QAGhjx7n4S0Ob6
7lNfuKxUyt+ZtNZa9thLcswVPUXAaUvxVzt+oHE98Zhs9D6QUIuD1i4prQhiUehW
/lY3mvg21FDzgMZdCagFqyyK6TvlBizBNOgCElaQ+No90pdLuK3OWKCb2E/XiM61
1dD7VnyrykkCkA6//3d5wJfsBXNOcBJmWr8SF4AiLaMIvYFjc/8zuKdiJte+PQSx
29+MakZYIrZxZLU3llXeggtbWWmIO7qbqkGoLNYJtozdJbvJP0so6Cx98B2uN9BM
Kgx1cMteeZfk9FKJiRzE/GqErdnl8SRtIwvZNSFKrQWWvS0fkbvg7n9cD3qO7x1/
qKwg8S7A2B6i6vEHxqxhhebbdYtWdMZ7OmCOpFf/TrRHR2ctjwtpQFm4lBOaZbFr
XSgEkmCoKHYglANv+M9JbnULJQiKS1iZIEe2MkHzk26uNCYFCYULe62+F/jXHbiv
fhFuQDK9/TeNXsYRz8PIftvi2mJkq8GDNSOa8QRre7YCcV0OScrQuhSMp2ijvrxH
JNAixYnlCwRGu/woPfJy1JqCdsW1HCSLuyMjG1AAuBOOF5z7tL5NTXZYSuBztpCy
XWET0AxlPA2xVjzby/a8VCaOAQPjjK28wQn+OwxM8nP4iRi1rl6Zo2DQC+jJH2ub
hI7BloejVRN8ZogUvOTddqHYJipfOR1Bx2H0SQsMUyIv33W9l2FI0PgZDlVSXzqq
Fe8COwTiHrOlxN0VppvsezQ8PlwyZt7+oGROmtCCjDWNaOYZxv3ziLYiY01HnU08
/5F7mFJKX9P3S+40dqGaCVSygwcbJ/1PeBDpup+WAzbwavWeGeqeIXrU1Ye0SkKS
e9yaBi6EEt5Gfru3lGVehyI8kawd+DPZ5qMNo71GS4Db1SDJ1XwJrfRavHvgyJj1
wqtKnsVfHYm9CqGrlEHMnAN6HyZZdpezn2ye+Kg5mwS2jL6lyvGnIkqGRWgbUEh2
AhRAa60jh6nl3R36nMV8fCP/dcjPCxwA5XjUZYcw0HBK6dt/8wR0yzJQu+LhNkSf
WMfAAGUfc6GV2b0uKHKggVXERLDzYinrYzvbu33F0cVTJ6O/06uTnot6zErKYhTw
7+aRtn7GSe9HBrjw85lTkSNEJvlZ+OZGrU/tzX6wBtutsOKzvp6tfYW9HEccS0y3
EIqr6Gxn7x9PFQW3tQfwY5qBOldADCZQDWs/WZcIw3chjc4tlYcercCHNVVIgWs9
1n04LPWgpCI9re1iz850lqJ/VeBmtMX4giw/lk9ViIiHjazfEoifXt9mgLjGg7ft
q/QSaCiF1zH6FwTSHswOf3vKGKgC+nFpdTNg87wlTXU1/BobUQtwP6zW2oX3c1SV
1vglADFXtCFc90/Cc8X1bR96mLug3EIoCCaN/nGcHlUoRKNlrqKhEJn/Ds97LytV
Jj9cT22XpJQr3SZzK4waJsMb4o8+9qBjEmAWGfLb4W8sU2p6A9WPLpd0mw36T7kC
/Lao/p2xInen7oVj1bJ+6KJDcERNwkPCPjmk3+O81ls5Dw6nw0OTlHGtb5TiGeMq
18iyKwuxIrwzpoLuVatulG9bwRFZERjseI23yYgmEAHTMpzbKg09/xvPnCBaJUU/
WwIJc9IMK3SIzmFgYyV8Krkg32LIhB5hM32ifbYu9JUnZACjYxlZirmRsawQa0jV
tRgKjzCiJ5sfnx9MwY8W93zTZrcDISBDtn0Ecz1oBtnR8pI8zwOZqPP+KGbHYEi1
u0/OYnPDYX4Zj243k0QA84yRJzYA+c+YlpsUtJf/f/Lb5uyH1xq6SAQO7oUzuPqy
yC6j4r9zT9vWw/D4knWK1emT7vFqBD3zfRhle2XXTpgWCh9+gY+nM4FlPiY5nq6R
chNLKviY/pgR2dTgxdlU4vB7KN51Fmdmh6fKX+uOETxR3lLrGEAP++WCVNltAU+W
UE8do1Zu9iycejSY75jYYHhHZqflZNQW4M80qzaDnYbVlfI0GDneaBjNftGHdUNZ
tNyq9yftJZGcjGdU8rYbg1tQ/3R2EFXQsMkRrZmnKv/8a5tKDkWu/qKG0DG1zYGc
o+CGrxCN1zF8qw45Lp5LpmYtphl8yeykk/2BoHzKnY0faJrFGj4fqqflzDtEFlCQ
pNIoZI2dUG6PyartGqwL7ZaqWS45/psWjCqDKOGxoYm94FA2u97roVI/h3TDH/2X
KfSEmq6Ebncjib4zvrFGoV4+PbOcc8j0/mWBxhfL9gKRvO8cF7vi4+v//FAU65Zw
2TDnYas/IH3qOsrkJimVQ0EW8kUGCEbAo/zKYhn69AmYjK7i80glH46JU5oBC+m5
AjGgJ3Hh7Amm89HRgoqFLkY5052swGDyNrGkjapV26E7+Ysy5lmBgD8CunkiIRQ0
WSbVy6uPBevHHic3YGjKy1ABVS+fYj096O+MVnXvJw6RJVyQNslKGUQn+QgagmJN
BwsLhfU6jbwChW6pWYClt8xhD318FIN079D0YgNyAKb0jyxWIsvmg1NsxVVqBVBn
KB1A6kHN5JY4o8XDg085TPenqGHQTmIkX2lAeYfDG+N2OzGWONGjFOptJRl2prnY
SG48R+qjijIF9h5/B/Z9jKKhxLiWI8jo9tCOU98ZeZ03Y6KSBC1j7NDuFWw3ZPhj
LYMPmqTAPCKh3yhdvfkOG9jl2n4Vf7Y1LpbSXi7vW7B3KgdnDnLvTvDfH8V8+LFy
sGu8zrmZkgNCA2X/61ia/toWRN+558SPlWLBnmWfBRyq9vG32hT8R1LmTShSVfN1
t/FGOH2zf2h4FF2Jo7N1XPHBEXl0WXQY6tp0SqrbDCEus4WI+phqUv+f00UV73ow
7vH7cKcYEP0jUvORJ29WKWSmnxAtgK/l3dDcXGpSBG60g6uG65VOfwtGeOGEzAap
P/KGBN12YQ24vkpHyNCMsWaszJRKAGMH5WiUXgHh7vJwV25GJVhS3BhEw/+mJK8j
6uCPtCraUTRmHLq200DGs3pSy37Va9dXXOC2sd5QWtHdy1ej/orNMR0MJ/c05Nd3
sD4k79Hdi7HHiBd/E4srw6EnEuc7zBq0Xlcn8AdTX2KbAlLnGaTLezpePRi6hX3q
sihNDhpFRnsPAdOhuRbgMlgwi+LJLm7s7/racd/IY4y9pxOcCX7Lh7r8Ng6+H2Tb
laoIBVNFZlK3k4UvYxfR+IOsm1byRrBdjqYdVf2YF1D7crjfoZ6elUXC0LIq8byf
jfidzaOylZaBgHMRtu1valXj1aqadtaZyf4o4cmqheh8ZzQ50u9H2U+5LDchuu5C
36JWVLz5PLc/SAzJAY5Yz5X7Om1qrFwYtA9YRBN6TNBc20tS3w/HeRU+gf0mQBUR
QV7Uxhg8yTArtLFb32NmkFWFIGJPilfpvh96bFNzhmZc0zhlwvYfyCemZ4Gyf/9g
CjzRKmJLMZdIHYEqKbJ2s300Hp6JgZ14q+lovBE0WN+d1ySO+oecw5nUmOE33bUs
V3WHpL5IcvzTKN/4agLV11xzmvbdcPo+SN4rH1yc38WuSdPxBPW1cPlSviHXS0uU
HKYrzz/qYTesP/YeORn5lWBtKn2ru4KQJ+D5778CAw6ZBoXoYnCvPp7GJc4BuvRA
dQPrM0Xp1+OMO/M3L+oHsLTkOt09l5K5eTt70JYqV5W3MguYZc5eG84GIcumu8TX
n9DCIZn8IAJsLHqLRCdjv164YyV+9zc+ymYgFzy6GJrZpNdkiwdhof9Gm/hFp18c
Lu7d8sUI/1gntM3PKiTJ7Im4l8IVFBPCjleIXuhFTI5R5Dmu9DSS6B5cYPwlkXfx
DEmfky9AGjpKHJWJ+rZFgiWf8Hylkab2d0DlGzNi0fzu4/Br3hX9TuK1gq9CNE10
Ri19riN8YM0q/fxC5l3uRspNauh66nbIetW7Iu07z2zTULSrpVSMx4R+1v4TG0mA
SXOcB8ukZmyAXaMueRTy0s/xcVTIYnNcbL6QqGlxvaPItPWCCdSTDwKUNdtW9Pfa
/HrrWV7NjQ9YylLWxaIyi/lUuFrc74/QhqEKcAAmccjvii8UKBEgdV7wtQ5eUd8F
eCUksXioi4GAy485PwPRwUw2XrVdm4JZH+mIuMlWzj9f52oWcYbib7tu1/gEhvd3
vnaRW2EA1eNjnKNNvutzipWDbMqc2zS/kc87HjRfh/kQW1ZUp22vaY+5N3kvFcp6
NZX5wYEotbg1JaFUqCBM4s9PLVcBSm+NxGMz512wP1l/b9ho81h/eg07GSjmuRyN
N/YPcOdl6yhPmoSMHLzyW/j6vEEU6JYJCssSU/cJ7oGgefpFMRI9XJffvNUW1Pga
6GMyE/tD5HoE35UeLpIu7AgLre1hPzmmLVvT0GiJcl46uytQXtP+xDcH1lVaeAs1
Ln9KbfhPNf932HFfK2E/1SCQxLnsJ41H9xPYB6pLyuinxPO+j9FkstTjtam67mYx
kzeWhEPDiREyeoyT9cBAdXiwg4vr2GTY5iIaKua+U0MCv5RvwWcVZDuL3g2MYnMg
aUn0nli66/ZtuxVEhYr3VWm3ceYzSbFyzRwyFZryGgyhUDL5iquyOe8cvCXdbqcw
SbdTXX2iYEFNo8iRvrlxut20GECIDsd/CWRs/BRCES4Us3GUZ5hHwQq7BMVDvA4V
RKXCCkaWf5KL1dmsryLRQPUENNvmMvGLrfh5tMabXp8i8IAbqjLUzwjMIDRYb42D
pG/hBJa3BXfuaKncc7AlkHhlUPYcPJHi/MRK+kepQTvVgYgg6jdKeNn7LhCkPLdk
d/swbORWXWKv2j528NQCh1vyVMIewKQMEfKSgvW14ab59Ft51ZUZ40on+WCfUAxI
mGg5eqwEjIcbbOdTfscxLSgiherKEJ85DpUQJqxV241THeTZxjNWihmNS9J20IZe
hR5jgageyVMA8asZ7UL+Gl51uXuRgZkeNT4XIzR61rExLJNuMOwsPkJQ8oXb58yv
sy4YheewUeB909/ZTpU9FVICLw6jGtktSrNtywsC4IphyChDwS0MY5dt/eeVZ427
ch1j6/Q1j1VatYmj7Tfo1RVRaDzVMM59yABeUgUKLb3KcHamTS/pfWjZpGS1AnBG
FBa03T1ijeaO0MSSTfIBPenh2ziTW7cKpoIo63ijWmNLAyKlf5SMVQ/noICpyIjl
G3E9Vi17ea+HNw4IYn12yLf+9xMNZoed5CTpRncpdcqHVsymyoJ7TuL/O14214O6
BlyzLeO0IoAKXbDy4ae/8P8zC803d5Wn2LjApwOj8//tpr2hDoMW4mgdicljGk3E
LafpvVxKmSO2tJhrbM+z/jC1n0an3r7sHYpV9KaZNOAvY9TOR/nJWxmdl2LISFd1
sugYMomemUfFDN2ExjwaASFeGACB3UikEH4eZ9JsQq+HPnuuZy8yPSLmm8vRb5ic
GMvl2BA3HODEKUF2TaBRB91j3Uo3DOM1VGRWSFZrBsN9d0SXHJAVlhQ3w98r3Pl2
Y6oIOoy15NwYKc25lNyE0VbJFJplm24WKw+CGt13BKRPqLjAlLbsBfQrA2vKcPCf
dE5euO/eP11ew+FFzmVpxlnKLBDzElCeErmsnAeLw9P+LboiygJtPa8TNTKD3rn1
BJQmv45ZZ7HfUX94MM/C0Smoe6efNTkMfwIzZpu4drnrufRO8OALSoHNbAWW1e1o
Xm9tPgdQGTNvaQJetUUtezEm+71uWbgh/qzc4tpMyQ1LxjiQu3FIG1WKqrOHUbNZ
jtWiotpbb7xPx+u6iFccI/DcWpKFz+ymJIu3uCTEF8HAe5xN/WVOUUBqyMvrzH5M
1Lv2jeCpLxGjGVA0wyvZVZCxozoC9qJYHWLwsCX2t+zCHwdhG02gpN3RxdeS6F72
8LxaK2KBwbSW6cWv4zRheVuS8C/OXfVzJ7+DqUkHn9CVALU+ikwJNsnxUkl4+nvC
BBGE+TkNlvDDxhYDg3LZjPECIBVkf3qxcCVNF1Jn2sYPTvj21fLH9nOoiLcFBcdJ
X+QbdqrkKy1lrOwIQEHdOHyPReRUAjJ8QS/uJ/Qj7fZrtgvOSXp/9NiRzlZMxSG5
tRRsKUI7iqJW1Q4ApVwhtqYpLvbjLKu0/G62DngRVXiLVm1y5i4j9kYhpMS+12Cx
obSfj306LonfeZPeqZNssQrqyNKt6RuE0dEK1GEsGrOQvnaPVm7WQT2fAehyd8+p
OSS4mVRr+aP4GLPBL9t6k3Wb88yuM6SlMC8q2Z6A92qnwhgJTT6J805Y5GpwpcE7
aKEo876/T7tleJI4WFezgwzy5DlhQrUzM0whQgKPcEE4ptMlvU9VxWnFxyilm0AT
K4Mim18aoXe5EzX5X2MaAVvOKG29IeBWaHs2uaCTFg8QPOJu87yfZWtub2mu1Pqx
HuH9HmnkKDHrsLEbpLlDs/gfQrQy+Uy/Cj2Rwoijp4MBlDXeKt/KV3YRHGTG1hrj
IeoZpPRBJEeRRJGwxFE8niMYX3YmKfg8tVMbzU9DhYd0tZPhOOKY8qGIXuhRwM1W
wfEmizwlVzXsoFjl76rRlD0cLyuR32c8p97JJ3ZWAdL3rainh9rggJ9HiJoNvTvy
0uyHpxSfSKsYW7GfZxGHEOPMefhgbQPPtq5vKgHD36dUxC9ciDGNo7m7uyE2ZGg+
cdj6cuPk24lZBiw89GH7nS7r9VKZW9khjdT6JqtOfYAxi5W1F5LfItTZcn69I3vz
GboVz1WO8r6CvpN76CMPMKbP9V7nFu+MvW8uCKZ7AbtmeIwQDAPFCbEzcuPNujB7
N+LWLRGIb4P51pUgyXVr0Plwv0s+U7jy82e/XnyGYdIWTqdAY0739RFXLV50ekjn
KoquKPtZj8X4Fkb0D88RhUvAnpNTW78Lw1iBebrajubn8znGlMPF/9PSc+QH146H
1/jHauLLMjDQLCNak1xPj1wBuDe0VNxfOvZS2NGoqFQ3PWtZoTN7tp2MV57DOXS7
gwuLu46mQ7Iib8AI3tzWaSepuMYdH40bmat8PiKpEB9JbEWzNdgrNunjxyxLsqUZ
3VcqvHGKllFibHPq5Usoe/ykcmoUZC1bwGfYih/0++Vhg7swBuX1zobQauvLxu8n
mejQ3gQhNNKteg/dWpn/CKmHVI9Oc6lYSy7ZD2JH0GDIich+pffqH+BrcQHZ7vWI
xDM/tkReMwHKPV1x/pGt5k0FHH5wbDcHLBISTv5czT+WnPHlYctHRU1AdFydU6KQ
iiLPkrUbX4GnSANwsXYeB68rPCyZlAIvyZ/gdsRt+Z0H542yxpZYKrfRFTiCcBDu
+6oL5D/ed9B0j5AfMZcdRQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jMZcA7J1Dm8sUR2TYX/9AqARR87bVq1cv3uc6tD4YJ5kN2kuikAzoWLptXfBNRqR
+UQfxNSDGUY/502sapJDYeO76/7I1HQTXStKIGqeMfI9QcSq8TghOK6BmLJSiHOQ
/a4+AguJODOYPXCHJ+nyWrHUTh8ML8o4tRe0tA5bmkDneNZ3Gm3JRyUve8ib814y
ojw/Kccm10CqgnpHE9o/PDA72H0fseBgw1T1jgAebtifsF8XWPDGhGF9lBBdRYfz
cYHwVYp3yWLnqh3ia1SkAID1Tf5QoRiT573NWfnpXAHoTzrS8TFUt8TDHIqWCDfC
kqKYhnB1/HdmzGfAKwEKLw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5632 )
`pragma protect data_block
yBA34urxq31sjHH5foFdQohzsXxY+ai/B+vib8Vqbq3k23WQVLEWCypPijbccJz/
yJ1SUiAEow540r0gix2Bp6gM7wuFsv4i40q4thgFeeJeenMss4zNQEYX0MWGAZS5
JPdLNj3wPnIwoTVckmHN0L4lDIukhXRUcO7RDXSw6JFFU0EcOvmZQzeQhfJdndtO
hy9re1T+PpeXRAn/k0AjiaEHXsgfHWsbXnpxntYEy2LBxfnJl93Z3rRePgnoo/z1
I5js9M62hPKX5xPHxdkxCjorFA9PjVmtFMTd4NNoTD8ax3wvxNMwadF8SMdW8TR3
z4dnwmljc3OX5sPyw0QGpYVQ4X1bnQc4Pf71ERQ3FPBm7oyia65/1sHW5egSE1NI
WyumBYeARaXsE1tBSFPoC1v2vUyO8EBi9TdkViCmdx4rI9j4uXRQ7o4HA2p6IV0g
u7H81Q3QOd5HFgNoP2sLQ1wikGj2PU0lYRhNKf+or925Ehs8KfbZ59YVXQhrZQw9
WUfUWue007DrdUFkwug8dwgznzpszh+E+QaH+sUy92rqLkh2AKCp4Da1diLAeaLV
Gf6wrGn1mL/mgoD9IgoGhzvDt45Lld8bMIuGm/e4FT9HPCoh0JM6Q0bUSBBiQTSJ
6CmImMu+mXWYtyQq1iAz34kwmvn4V+vfvgd3SXajTdbVayBVhk5TCjBcefeuBggY
UoAV2MSEP3vVK6+/sCMmSrP+6D+z/SeFgMsRV6LeOVpjJ8DHsdsmS5JRcly4g8bP
O1PWCP0XorVSLing67hIDk5K6DuA8mWTd3nOptaHBpD0j1zzBNGh8sKLMnIyQis1
AWl3B70iMVxdGolKaWMnNfftUw95O7z99HSHovYOsjaqiGTY6fMdDrycKz0/GUDQ
hIlRRtGPvs67FHDI8J1DU2xtWt6NgRbqV4dQ2tG4WXrZviI3y8iJKw2rgzNXNyoX
kWaWrCXK71guRpP2mjqXGjaRUDF/hw0K3M2aibvK8zRwZ5Gcuk3qAJx6UwDKD+sG
AaV9C1XPsYco2bmf07W+SGcWN/VyxPHF4X7wCsyy7t3l7YI/opL4VopPU+zq9gdl
Ysat5BdTGIuMu7pMMXCXKlx48t4R9qh7egcE17Ux5K806lUC+Qwz/sjqCHzMqop0
X1x8l2y5v8uZkhWZua5/wT34dSMjxJHQJZ9itGnsKJDXBmFOTTXSneyG0NAigvlU
kiA8w8/Sf/RUugp0zospQPvlwEpBa+YIpGZ8D+mw1eyZpMgKajPxGh4R9cIGI3lQ
V62yi/zRV3unj0JW5He8cfcV5CZprkqItmZSoyhTCqz7AJoN22OqxsVdmevewPBk
ODvdS4w9Um/vn5uEzTsR+GTyouY0hGhgsnlHDGpc/6AS1MuQxvMETMRpnEVGS2Lv
+8YXqa/kYSshIKsEYWmxXQv+bPu2djYu5ms/+XS/UbJabcYikEF++/gSDLTNBTkf
IrcFHvS6DHpNX0kNa/wWgEoTXn0r3JzyLydJbdluf2E2dSPYQKDsb41syNC6CwYw
DPSwU2OM+r36ny3mujx0dS7A4303pRC4YrLZhQ9eCuNSA2fhRo569OK3088JShAY
Uj1Ql4nnExsQ4Lm6AI4dXc9P2GGwtwH/VqpAz4+63BlnNuYfRCUZKTk1cXMloytE
AsT0kvrb1ULT2ykMwlLjX0x19EDey9n+sav8ML4GbybXkj4P5LmELiZN5p34dMGV
6JywQBiEZP0EBUzszMznBXuoi00+M8FlKtOfXk+8zEwQuRzg5aIrWmngqf3ufOx3
hbdXt8dTeSbdnE96iR/p4wpTqlUAu7lXLMpsxnFL3lQTT0pM/TCUx5biccaeyOqg
5GVf0iXm2RcDpFvXliOIATOlSrm9DzaUR+e56JlMsTpfez+a4CV80q09OnC99oPZ
uv/MgMUde0mKmnxM5+Gz44N5LpnLVsHNLPoDfXfWbghbF8CaaoXWE6hxMnsa4fk5
4XALwgikoWg96GH+pnj8XWg2yiNhzmK8WecvUbYvh3Ocn/GQbSZZhfo45gtycICf
KCIflxzQDuB/gvBUPXrP65Pdc1bshy3DszD+oeUZwMtIJCZa++r8H6e7r/29q+63
iJGxl6l2hKvjSZhwkrnfWmUVVeEx4uu3nDHoRKj9Zw0aGRux9Y3YKqq9cHVh/yEp
nMk11xNmntWjwCrCeCoRNPlIYM4q9B9rJvG9fjvFwsLOpkUOvxZnw+Y6Za4QRbn5
BVKXVNjLs0MSLddjhD6IJqkUtYF/SjyNySND1nZxy9+jsMnp1HPnQru2u5MfY36D
2nalbB1yq9We1e1EwepFZZecK9FLDp0BRRqg+HR8RLuHGw96kY0fEPTZKU+jw6Aa
NYDdo0CGkXB/rf874MkIfC49FQNOanBiv4btF9UHXe8U67qsB/vhCGFh/tkCqsOQ
lF+BUAtZNOgRtoJW93afqGqOvP9a2RDEV6PKRiRFugXRUhKDVc040mcsKlXQkPk1
yUNtYfN6xkUjPl49/5zSz7b/Efukz97GDyO4F9/7gvxCb21Ixm9+ynkfW1Aqpgo9
Xd5W5d0DTzNiDU/BrhZ63XZ5iy/9uwMxAM6BFKMu3mIc+sDwBj+xa/JbWvcHBuuz
Y8+lZO5OXSZq4aay7lJl05GaTyG5mSZH9JkkTksfNnQ3EkVxxPVCyU1II+/6yuKp
Gz98fyiu45O8eKaQ+1FbnNpWHis6zHJiKbqrl3PI75yTIj0KOAkoxBo5/tL+D5uT
kVr0sSXRau5+7H46RwlFuXcm311kbhOqeaLoPh48Mba1FCiS0CfAxzUWigL13fk0
Nw0TpxUfyOCGGa2NYAAg6DK4K6XHcjH+HFbi4Kc1znYM7FKlgJrAcMhv1ss6nkN9
eQClrMy4VxXi9iqvin4hQPc0Qav2hJIu1J0hT3DolKoNU3ov0W/JZLo44MDkAGFt
VZpUcLX9CJ4cEiLuM35Fx9RSdCiUqvG9+k2mK+L5N0pwxK4jQSUoQDgUnAcc+oLw
0Zga1ae5HJKlGrJXYPYtPeaDPiOkMprNWKwJ26fmVhPx9vqlPNqz3fxuw0AxhY5e
7xXF5cHvtLIFoHLBVEjY3wdug11VzBSI8+XpN+1W3nqEAqAQIUcuxhGsP3sZKW7b
kojxO5OX8zHwU6KhJgoSbTgADIvpZvTgAbFtg0gJrjeOlLARBUZu7TAbwHnTK8YE
rB3ly0IAO1ndJUrlrg1/hYKoPV58rWePb18/8atcY46FCNaEF1wjKQNjkNL/dM16
d8Q397geXjMb/a5HwshlJqi3J1Su2CNf0SQGwiTiHw1nnby0y2BAmurwMLZ3cqOp
jW6dJwx34ioE0WH9C2nH9/WSMPj65TQjzG2Nt/esm7e1RnsrYEULN0Ug7/PNBZIx
doQC2ZcjZYryDNeoBwXrnYTge0pyLKWnqzHtH4hedShrrXY6k9qNw3nUxstyqgI0
SD1q/Xzo+H0aODiJqMm4Tfy7fNIcox3x26FMJaKzb5vhQOESzBeYnrX6lCkTm3wu
qXV58AX0U3Y0uG2daW0pK0GH54ZK3jBjxo+ff/57bGGZjCBCppfnCpYES4iYPOyj
nSMWFxzzIkTE3mDpyFSc3PZCR+UUcjcOQRnVOeWRqvyOqmRXXrm79YWhawzYHvMf
vyNHKjb9llRqXqCkpNRMXRO103poP13j0+2HRgCZHlu2W5M+KCc58VzeuBVEl1/d
3JNOxzC2YUa5lD2wSy2LXLgTJv8OgHeMpEJDVB9QWI+RCAR6nGfAVcOeRM7fYFlx
BItyaCCPRHnqLDEgmcJFacknOmmb5G02IzmtD1Weo2XPewyE+BOmdkAl3CfjnFze
pTXv2rIUGtCmm/GkSRfZk0wxD96ffs2PRnEuSg4muHlj3eDWGXMzvkDwFvEiqGi4
l5bI2tixzGRI/+VCwHwS9Htf9X3iTaLeVMhuOHgvBStzd/xi8ICJd//biBC/oJUB
98wsdgjl0y0gZmpReGJO8zjb9HfQXIg6x06XZbCEdM30Ufl1z1CMgcbA1ABr+qjb
7rXwC0+uPGthtg1d2fXV41MTN2xO2nguuJ3EwDaBohixJdBhxidKWM+F/xN+Fmfy
T+qWgfBkbCKNweTMwEn7dN2AS+HEWVDyZgyc/8C6QFDfCZ8QxChbUPbIi4uCy0Nq
xqam4QYKqosuzuoc8GWUCNuHHOKxRSBWexZ+Vimwyuh6WE+8n6lGjxHJkIjk04tb
cLfAadVtwmDOgppnOgESX4JA5KnQg+MHtrHjqYwHkddqRNeZyAI1o1oTkSwFdRRM
LOtXkNvAxtpOWN6XTQU9jbg8C3IOSaZRRwOSENPzqw+5nBY9TZ76A9lCVNgmnz7j
VkdIYZUywfbhvRQkvjrTDtA/1gEbhZjRTnMJK0LfnTqTsFoE5cggJ7GP9Xeee/fA
8KYzSUowWJr5nk5qOTNCIvnbmQC7IwuZiB+UX1vcRAalzzn/qI6vQn8PH15fzdO2
gl5q7d4I1y0LOoeQ+Cz4l1p0xONMGD3dFZ1fPAUmEaHqt/7Kbnbx6omgQxMdMAvV
rqOzc949aXlPyvWMckkws4HOxz0SnW/MAe2tjdN6Qy5P0JsFxoEWJvC6Rta+Q4Fm
lCdTJwN+Yaa9p5QjkGiS3kD5P+NnzNl7gRpJ1KDs0NQCzqEvpfCeloFxFjCNS5Q3
5iZt2a9KYEETWPSPhWMuTIKmmKu5/k/v8lP14BT27BiLaMDurMN1PATbvv22pUie
TrztDzH2+DZSf2r71s/SLmOWbLsCi023PeLWpXCAS1p0PLgE38vo0VfveKE+g5xS
Rv7IBCLC21eD0lALVIuX8QVSLrBLjsWRaX9+Jm1J+UtAacuPdLGKN0IZfCxWHLNj
eB9Tw2cOpYV1BawZfD/tJju2bDt/B1zvKlT/aqqLhdTB/5WCp80oP2EsagBP+lTE
/8MVgM59baugq1CIc9UqCATmpFMO6HrVc/7Z6MIzYGoo5T31kY7SB+SIID20knOH
9dpgM+a3m3p8xODe4EYi07LwOO0sHRsiaJmU6eKkaDRr17VGEbHg+bZ2vSBGhT/p
vyXcnnIHsT7Fv4UgI/BIZnT0JgBtKv9CEM567nVV6vh7P/iF4RcSlBNYopXCPrZs
KcvGnYrQ1wlfiWkwKBpJJ/aPIHo59StlzImQlctALTt80Sxh1CecD9MjGdIwR+5u
kMZpIUEF0PgLlHN2SiEXceAlp/bHAocRL0yCjpyuzpS0GuOUKZwFjpaJfOgBPrKY
aguRQxX/izc1YRSdnPkcuPYy9/FXLWceZITTxfVSsQdO9uzPkoQ7aZEl1/3dH66/
fEEfR0q/sngw5U0Gus/fuoeyZ99BrRpY/PEPOmpHuAVv2wHvZPmoSigAc12x7xqt
d8QPPwTdkI6swpl5+l+2KS58h9KOFUiQAyZwD49U/yXSWkllkEMKEoy1v2egM7cq
xHNBe97Hmbpwam7XgREwW833Jj0ZXI1kiqIGDBO7OJdU39sTiG2jxvcwyFtiSLfD
Kf/TNU6tR86kwaTHa0lVKM8EdsCU4olgUvgYGtwktZT6Y4ZPsHuwkHf+3ySBSsKj
QPzMfZQOd9EP+pxRZ/pN9lv+6z59xokZRnKap6n2zhi0nM7zkhz82Zy8iqgMkLCZ
8wHmz9i8bvY9GxYIx+vkRfO6uC0IE8cU7dwazj47XQZQSqvVF6Q0hewL/aaATu7l
mVCeZtn1v9m5ybioKN145fvlPM4t7HKczOHk0OSMj3Y/nFcpD8OgxxCXPC8guXzR
yD2KaG4tkukMDus9ATkVVgd8b/syMg7P83kRJ7lHg1bdVfinQd9NUxYw1ghi0c+6
YzKAsoqwsA/aGoODHzoCH3bNaDZ85T7YRJ/w+5AGifbuCMNELMPuS4aMVJeNCTL6
XuMz33Xy9w7LUR3bMyka2aF9hcmviQdNxOvrYgwK5RDjTBmzaEdq4BnBqRRUYvcT
zgmTOO+kOLXwRelCtJDlYf/a2IH9HFziEaz2hM+8VpKKMwVzV0wvwDp29uVcUbY2
HbUKXr5UQJiCiHHcuSlh804zg9Z79nVlmWZ/3vRwU2KoOG68u20ryEap9q7zGsOz
PR/Y6QGQTaI1I2mqQWEb8GkVs14FOFCxOZQBfIuyQpSXJoAVTvseyG20+Iu75fY6
Td8JEnln9n9PRd/+yrROAs+fclIxN7Ow8Z7VJMv5u+pgZDG5MqM4zup9ZUFnXWZl
++cTn4/9x5bSGln8h/5g/pA+gH2WzKD5Hd7qCLweFKrpROtEh0hZvUbXN34H3nMc
Qg62OFi6osnRRli0IbvJpB+znfsxiWCHhvfww8b+4OiWRXdyL1vp1BtxzgMAqp3/
4ofO8cKjgH+J67hrq0o83PhPCfH19TKMDJA73uOdS0yQHSmbN2iN7XiJm9mcmcAT
18l5dU6QwijtwG7vgClircALeXm5jmb+yAYisdDofdY4JGmOj6v20A3br8PZwLJJ
Vrx67dr2k9VAWYG+1QcB9V7W9FvUuXJawxSbqG/qv1bv3dfwbyVL+VAyTYM6/XnR
o6YCLOlOK1+5sHpW/oLINmwzg+exeloNQc4ZpLtvgv554vMo4y8PXMRplD0puNBJ
G2zaNNBh0nxdQwlp5eSfGHZxWawX9NajxIA+CPO9UdjHqcz2FvWWnXiicOMZ/Z13
qhkf2LB+CP/Qm9SKfc6RLdPBmKbYE4BVjXdDj8aG9fdnAGbGVBORJPrBm6LBiwmv
IeBz3ZSLfbqNYZAYcVChDi/SVlyWo9sAgKEPESahZoyWrZQNODj7yKCgQLQKVRjH
nwrzTCxjVGbk1iVMmsA207Yv6A4BiX3C4pKNCm+FBlexB8Y5oKb9uHBvS7qOeDus
26lNghIzLBBXQUPCvK0Whnb0L8vw5qgWNe6pNrfY6dMeUO/k8oY2RrqeLSMrFUJw
+ZvvCjbxf8qNeyriqwO3zicQ4RI5kGhRk3aS9OU6q/U1n4kbWoyDDe1fshsYWVfz
tcG0LkMgk3p1w/6TRnG0PNeJQJegqVCnvONnL9CLI9F0tkikBKsdiRHL6ndb+KCC
Kmxm8b74NC+9o4rUgzl7WdRmfviVY6YvK+Z6GM97rPniejBRUA/EjDP0ZUlMFII4
KA8sHCbNI6XUZSp6AYLWS2J4PhOxk8ICn+unymqsq82t98Kkr23qnAsPni0cVgTY
r5SUUV4vzFXiYBs6msG9ayRfK4Mb3KSTEK4d/jTR6wt+yw7+QixN3ioDhUthTuyJ
UZXIm5O22nPBSa1JFbN/JeeKqjBoMq+6gB2P7uzPSaM+OOaGX0/afzA/Szrm/JBO
Ss3CBG+G61PEyDyP9vwCz+XAeJdNX7oVqLiAYuJcJKrVOatOeVizHkEu53bHiJ3C
8s5mXzkEF4wSlMWbYy4K9rVgJeurH++ijVDFfTqg/nOlRUBJmDPt+Gg1mOnsEOSd
76O9m5uohu1oi9ChDe2li/JFnuUmy4j6TIM8TwJDt9ihnaVD8V8lE5ik/61e4VZO
pLOeTAkhCerLQ0oFOkRZdg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
C8k3+wi1DXHRQG6ZpbITmsIPcQQsN3nLhYKloCq7WjNXqoYTffXVj6Fm5MdY3Etw
lAAkTeY9xAB8HWM4J304Dxkq+AZFjJuZnsW1aC6AGCsXqpfmJ1dnEYunVPL1Qssb
2kQ0tB2Ekyj9i8YZxVXn8h/NK1F8fwlZAP+0CXviyOrL4uqmAazC0snUREDj5LOt
F13q3s3h5kVUl/UNIQg7Mu330zi3O0vhmNakqTHAVvqnVDdMqKOA3zUmWK1qpbW/
CDi2sAy+cuB8GrqyAY5qZpq68+ybFTUOOpdpyRl+X0Sc4AzFvShTvlkGvD6ytkKC
A9Kw34qAcILLaQB0YQ8Lpg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4928 )
`pragma protect data_block
g+6DGKHZGcQN5xRvGf5+v7hXWTDSdfUKZC+uPnWFA+iP647VsCvYTsb0PhAkMuNG
kqLRayt1WAE2K42liPG12vwnAk/jjDrgMA7Cp/dwV0dPh+ghSU6gjVpUbmYge7hj
EehDFgUgeuKMW857DFjqcP/eXnefDpMhMAEuuFSfYipmOKjIWSleZRJOuKg3ZhhU
1GsLQ+mMIe8YmOCRhXeIl/poNWewM/liou5MqXfPLaoslepf9oHN3xkxoUtiax3E
bGHoGRNuoMLFeIDevkZJJqCx4yNCjjcLtdhzXho2DXbpoy61rZOq5Ft84YvnbVV6
TcW+MNkU5sQ/5xACTZ/tvE9vWPy9wJZyaXuACralUwB3OdQ+1OjLmk5kgBiYkbbu
BmOlKS4COdvAwy5vFKKz7Gj0jelMrpF3G4Fk0KvJjsfQZwg7r/euPqReVWREKg9Y
+8zWA9/fPxl/wI9S1vwoo+l0CJQWDhXauAc74O4wVj1MBos0wfp+PRPB6F7Hd/mK
6gZEGFKKHgLQPZ7aVUwcF+Xpb5keRkzTALLZY117SQSxFzocivEaGSpc9DVWthEG
JizTqUGuOuRb3vBWVOpjbC1dfOmyJJZTCGWedgMFil8FKCCVQYX1m7VBzz1nNb6q
Q75PBou5tsVJp7JKPBWAXpUC/PlU5ZuI4JIWort1RvywnHc5/T6ZwbJ9HPGqek65
IzwqPrRqQpyptUnXBpBCfL1R/7LmU20NvCuCckyJxh/oKnA9dySXFTzUHvKBPfvm
hoqrUIv3olAlvc+iCFEgl6BkQIuReBpTpCkG+63ZPMrHMWYhZgRi3rY6b0QpeAo4
7osszhter3HnVsz1wB/fcmCYuz9Js9Wwmgik1thSKPqYAOxnWIxVlKp8j5kbRSCO
FTBK4GdaNG3qxJG2C82ZRdEiHznqNVWbOS3q01GiSPTPJXXgXdLwb4mwUkVp64LX
tVoQJMRyfeq6Ew7RBCwCg1S7379oQPLCJz4qXsiBYaTmnM6tQIGsgEPhmwRWh0bs
84KAyImbyLnZLHsK6siyL0kSDawXrKMYh3TvJRyjUTWEAeGvMEUXgEeFgymdKQRM
9A1pB9CV2j50EFIRqUKt/jduEksfDLqd2pvtxmyJ4EVZECyxTcgoKK75AOfOCMcl
edIJpPcLss50EkHSlJxuaHh+cAOR6qUjpbUGg1llnq/AXqw56BfTzxwX9XKnBSFt
/SxMDwR1dQoTzPcruEXzkYz2k/SCkydKfGHdOgyJXfKKU4jfPdxfUpOHBE7Cs5HH
1XL0tfnc98+WKTUUICpAnI0vHmPNwKnEultNurqhdD9l/y7wevb3nTOG3fhtDJ6u
/oEBB1E8SrBOKfwQj0oxWQHiDSI8kosSvsWLJQPT1SEf8/uGMGNb9nroPyLzsL+1
xFTOgZeCXxkRvrLsbzBw/lyvZTTQOcWmDnbStFGzRY/wxr4grkDt7d1bNIUIbRBe
oUUdF5BkSv7e35mG/kI5TvmuD+6l4mZIJxZzz1W11vY9wKnocuZj18+pgyoFIiRa
mNrbZ0C5o5aqZJsk7IJCSBJI70B1oDIWm4ec8q17Y4DU2o9oafeOkZErltifr1nz
IHzm7mdEOrYs+8UzUDSmPybSX3ZBxVPL5p5PzQfLaIDQ/7welE/iFgMFzRRnXI6C
VRx08aQLTg3XOIG0kj8+1gG3IzsJBayoG4D8zITiDIxAJ7nh1X4y8xBmYrHXgG/V
KDgfPwIKd96NIYmPlcJE+oFk7I5PfRsNjKkqPugLW4KkazD9XYxJyNb3frsmKJ5a
M06m+JzyMKggurn2NPatf9Yn+XX6k+4dxzrbhcZ2FHit2uOMtQ3+os+eliW4Kbuc
pi24PXyVDGBUkTHXXXEPJtufNWq3RHTMHI+N4i4vwHjIEKtOlOfe14Pl6tXlsmy2
7tn0OO+9rMY+rl4Nfy7oAwE8MjyEP1tNet9IPUWWiDlRX744GvibgyyELfVCc9oe
RqS3QFhfJCQgamN5+Km1HEEJ115HrUJRO9NnIspCR+3qBTgU/PefJK/JDS0KYo3U
5VEE7pA2bxiKve6/kWDSEFGgB9muyPoyZrsdFxRsmTJlAc6fCA8geklRPkAQuXSS
dRJUuFYFgYTzEwERWPv9ICtjC4F3Z+TqFzxUzodI5Vx8Yk2oHgSnsELLo65GUvcx
T9lLYKv3pqTNfFhWv4ZHD2FOg2AUjTQGqEZ+nFVUYC9mjklhuGFDjaLa6k5AuJdI
B1Cwo6vA4Q7jPH2SkedNIqko+qs2FM2SVCxh8FFPBHChy/r829F4ouaiNBbY6aVe
Yu2bOfaxiUHs6mydVi0zediovkvoLpbmAa6BeVmo32GiSKQ79rls1cw8ZGViLfNV
kLWVxC7ZeYOA31spRNklA6HK0nQqv2WJ+rJanjeNu0XgZ7FP+iiPreddJxYKXm7E
rUut0sSpeYLMIzv4XfmKBM9tL6Lgaj89hzQaS8cOy3ZF1g74v7dxKTXc7SnN4Wgq
gMCdKsMNWkZzrY5m/BzOqR8qP5QzlBPFCv+qLobqnKR4RhHQKM8sfoIHNJnFThl5
iL6sauuqRYRXtV2MuAtTuRe9oKpEXQdXffCHQk+knvjgCYWz/3Us9TfiOA/6xGTU
2cY5Qn6A4/NOYHvJnEbjhLumbKY2cx0em0LU/681sHP1WP1I413HfK+C9sfHRuno
zbdunsAh509QQQ9VEIhGVncAQQSIy8Wuj++oYl0XpbpdQtUNuRdJQuI/GmWDFa27
vvHgdOmHnAe9+GZzdUB8qV9pQnk0OAn5UPuSCS46v26UEOA0uB3JHzx9YxcjSLBB
3qf1vSXZAIdr8iqHu0ynK10LihOleUEFg/hR2IUAWw6Zm3ob6HSUMyaREIYxBbPg
doyOQ/Be3Fpb/uoFINGLdy6SmpwQY57Nt19vlHLLp4gsYrjL/gRx1ROrK4LcQ677
Wu9XpfGq4XHLyZhyT9T/8wV5V7J+CeBz/N47ydsTCgbHR+hAjYOTQOhKnhFtRoM4
paHUtFjOD2TRDBCWii/B2QoctY6uYBEGGKIpHdkJeq4LXpJAHlZzLO2CFZEHRM5Z
BhNyCULFECTdITIB5NJE+Q2Y3hCjkd7uVFunCO4ICswfkBU162wU3ZlC8D/4yEHt
m+0kbp8k1XQuahoXyaoycPcMYvxo+zl6DT5pivh9T54+/0pWp6ZHerfBKlaakL94
wAWLQrh/1mH8P+EE+DXFX1/4QG3M1xCzYE9URRLQY86BUyKj1nNct70rs+vKgJhj
I86GYhqJBxo0xs0LgJG1n4XbtsKWg4CxpOjtaa95gLRSeEnPuV12TSNqGUZWNTC1
t4M+bHbOu9GJLN93uYRug8LRatMiPYMIx/TSUZd1hfyMObcuSpwM20TVousLvtLf
fYS98ES8cRjDfZO98S+sjJvNEvSvriGp+7RdhU8zw/+MnS6tvZ6zbW3YexgbVkXM
lQxQZEQeNQ+o2rSuidW9S+PEyG1wxe0IPdiSr2eXVZKlARuf7EnyZ4CO2iPCn+Ct
N0fXLeGsUpK0C/xYUk+bJaFfphk74Zz6pAwDTA0s7m+RtYRORYvCs00HzUHRupV9
w2T87k24I84sUL61kAp9gdKe6x4661nCscQd4I/l8ibim/SMaCjTBZGwQw/YnsXs
ApTfd4IRcp1Ct9o/3lsTfx3DgFdrgKRfO0JiIklxeVBPQixZx41HsAVIhD/oSwYy
rhxurO0uqU+wBn1/0BsCRIvnCPNy3cXojPWMVUVlfNbJrsBAgh+8g+oYf0319YKy
A/CJS9fSm5BnZ645OEy/lL0QBn0hjHndokzQUIRGXYPB7mTtj9llac96pp1wNIGA
zMj+s5kwCahe3sKg74LqWwdiieGXQY8ho49Zaob9IUp62vbh60rjJnr06jmu87ss
DCa2wthrwVi0bskKWhsGNQfaqvqug8UxYjSOaeFVJ575GUtrXTA9vQjWHqlC5YNe
RutO1NXLyDhaceX8AXh1okXjDKW3VCUZqV4Gc0Jhu+YXJecjENzr+gvavWeXhGEH
YNBGVSLhPS7KjNMJQIn1mqxgjr6oZciUs6CHmmg3tOMn8GOv+hQqxdDBd1/Oupxm
bJyfC3ttxr00K3HNKt2dhJyfExCRTc/NLGNdrTlKbISggNrXfmWZ+ma1zM64j9wM
ZvCjBPLjn0ffYMPLy4YnhdsyC1tgQ+HUeihnpzdZlXnXRKCR+emVcddHPHgbyZPQ
r6eqoEH2pmLzwczRSu1IhQIhV/aL873FDvD/Fx7aM08OL/tQfB5V0yOaVi/Mty3i
Hl10xxgl0JSq1kHgkJLEcCxXrH+yB3qdiWdF972Xw7oixWikYTdox2Wu6ZeoR96r
2f61GqmPHBU8KICCyca/3GqUgY0Z86XT7cJ2zIcCls44qILwBROFj230LT4ypUh/
rdEiifBZUe7GfCFUzUQ8GsLfUypsgk0hi6Go1TkRuQKhFc7kOwUQUmsmkaSf1UL5
mor32qrp96bkgd6Fdz2ty0VUBsxEHzFT/UBmXGUcL4G4ybgoWe9EIruZA9Py8hR0
SX82NYcppw4UQo3keXDAfp80D3lOp4+U2mGysbRtyZI45Y9M7yd29xQaNRry96M6
HllKrt/epxEiAR7UjzX4e3pnGwDR4/2tvedSnfk0m+0oPFAJnsL0JQgx4ws3ECHR
T1la/2cMa8MVuLHBgQjU4BOkOOyydnV3oF/CvLlRHnoryEXTAj8slCa6oXsNsX0m
Hjzk4oa0JIJbqLM6UrgYNKXa+0ETPlGF1TNy+hY8RMUwmoFKFjEd8P+YuXf/dj3+
RiFp1eWPjOS1yn5wN6heDZR80bMuYKGXjuYYhekRxWrl9HKZzyNeiKFqdE1DYztK
wbI6wFAtAOArazXKWJUru2DFJ9KTtLYMz6DO18v6c1GjmcI441nSLSzHSbz3nH7p
Dud2eBwQS3WsF7Zv5QT5ZC1YBwxseC85zSMUaEaGAPoWEt94eSSzECDp0Blf049Q
GLUChXIAnY/fzu3aDVopj++jlFCIGpkfivQMf7smiuzDyhFupUd9Ds6k0odGr5Xn
vlE8VCkY12UjnhM9+Xmd7C3le40O+vvAiodZ0Hptobuk3XrA6V0Z5uHgHll1eL/6
tFIwEqdFu5yufYoDT1620NmUSKJXA+AXtpOAEzL5p3LzdQqGC2MV48WeD/O2LRjd
xa2mTWOF1pXxZdSHbmXdpkeXa8ZlebFUT4N6Rty6vyfvtRsAxQVqJoFRRbE4vcq3
m4bvaLgeBK9GXwblaUusBQ3PVAERX7ZBkPL8/c8Q5gj0ZXFMQ3/3hSMXVvj6rSHB
c35WH4y5vGKMctz97id6UsewxfdvF6RYOlTcobKITJTTnrj4li+WBHKp8vS5uCnK
A8EJa5Auvl5HXUf1PILePAsdo+SSj6NUP3S20pp+LG7f3AybUFN6EUxPMhJxsYKr
rEZ47EeMf+TG+xC88kzZwKxUkZgAKVTRXYflrsjWFLmeEFjPUAaxNenDwJjKUAV8
F5cWnTpoIOx0Fz18VhO2jkuNWYpMe7wxPxydfKfdVRPyHM+e8dr/2orEemneKkZ0
xxSIUNJnLclRYtDDUm+KSg1X5Uk/rzzGBBPsa5a+IAnEjb1tN4JGohcVLHuPm3wU
8z5Zg2TvHj43pzg1NnaIxSPr+f2nqWfs5KQjJdibSGgVLt1heVbXTuP+8EoWFXNH
cnWfabqbomhjdWSCOLurrkhKoD5rFllV+oYLjlqtPOSfTJilcIdFPB5DB+FbwHW8
KtTEBUY4CmNOzLnjw6OmSImuKTETAon4Sr0RnqustPIA7AesrYADHEsOODZFlK3K
Vx+VwjzPJMIlD+R3TbM+R6oitb7U0CWs39LnkHGSPPmEqF9sVLwQQmPt7NZW6l2c
GH5vJFPTiipawedor8LjW0AsotfcffN6wy2CkKCDrsFu9VrEQC08vmjLSA5yQRyV
0DFTUK+yHPdBJH+gdAJZpiEnXEQfzDzmI4faU9L2ODR1SM4Gf4jpnb6HwEX/98lk
/YtAmxxqHocotrt5SBazvfJsavBdF68lPkyYVvRAU949P/ZTctCXYgpDBAUbjj8x
1M0gFR4PP4GtfpZh5DujS3ZmM8lI3STsSqUQuYUoK4l4OIS7pntLTUDZv4odNLA5
w13pkRQakLME6ws0tx1rwjBY9+5aWJ66omwUt7EXFo4RBE87KOgqGBFJhyePoNH+
oSMy0EVtOuKKps+4dkgZL9IOruQlsbhScLskdzzkY3ey2coEjqy4R8VdHEJR4zjp
lkf1iYQR2tQsmCjsXdoC4Uuqkf18c/TmUMXo5F5oCZD4lax4WtM72l+Y7tMV8faE
UgS0Zn5gXM5gfo0OSq5Yb3q0+jO2OHTlI+jJF1rzHDnM+nvI3N6GDYB4GAPjHb1i
UOLuxtlx0AaMCjmJfSWYMeeyTQkS1be/zmosr1k/7KxP8zNmp4kdcTzScswwv4rn
nrOwQGJmZRwCKuIJ75j9KivXpiv8pErgqyplN9+0Yc4st17hsbIgsfYPcU6KK7ED
ZDjmy7Zw8Lhf6iFjNVuphfutyObnJH7u+tnCGDpfac0=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
G5yZHKcJWNIM8TauDJd1Mb5J6og3l/wjdh+VMgeO2+vvYXdZQU0hs4GbZdENo/B5
/LL554Xz+/BuEbdU6wLbUe3ZHxcWHkbB226hyJP9/lCgzOMqqSt/Mt6iIwJUg3c9
lW2X2XXCR9dgsSJQdqU2EPPsKEyvWD09BWR6CV3rjPK+AEBGBNlIgEZSY5v2rcHV
S7mOyNlJ+gQPqvkwArYJllHRdSD0FZJFcs+DEvn1bffQiRAaEqr3faxetaxcsJZM
lUn3jQZ5L++E9gbuSUMXrKRf8iN79otW8D3TkXAECuU4gvyLlh96NOGwuVUo/LYS
+BJT7ajaf4e9btf04gLmPQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9792 )
`pragma protect data_block
YYRD5NhnJkM8Nh3ozifkNXsYMNmw7IImxv4O52z5uL6L44WpDFJ6EC3NJtawoaii
sd12SKVFcqHO+AhAJUWpGQLA9Ob3iuzG7t8r3biYwWw/QuSHwBr1bzEaJ162NFpW
w1a+prlXzPY9skwXjBS4pB1WDNGBemDMRFaIihSg/6UnMVvB1wM/bHsj68ZqAX4l
KgXL5My9tdMVtErzH6p6ZLCc7gthexKOJU6f6daWd1u7mfUsGKNCQZURKVp58OD1
hGP/BAuSLkXXIPFlWctTyy9Cic5I6vVOrDYtyR6TrNTs1iw/bMYr91HYnYMqCOJJ
73AZRyexwWQZaDMPfONxjced2EqpdxAb3ZTQhJN9H7/t/dnVRaVfEBTNz3cNlrvt
Rlu8UQ6CnKFogNn+O15C25RNqNmJ2yrEuaWM4SJMwWuByADZmJeYEWMTNO+RYUkL
Tu3GQ6NpFBdEOGNQ0Q056DSiClqaIE6R+ZiW8FQN9sLF+90KJowwr4unjd/Y6094
y6T6TT6yBwnI12x/Wklu+WcfMknvveNVyl9HrB2xF96qCxsyBRKlSDSxRC+yP7Sv
VrYcbCHbfwoEQTS0PS8EwGljLBbXvjY/lVFFNCNqQsNM0/jzpjeaNua990PeCp6O
sZUgkRu5nTBKQ1Efaq1hsxD8p+hkFRNleWVdohpS9Lhh5konQnTv+jQ+nsUvqUOJ
HMxM4uHdHaiZdDN11ly86UJgWzlY/PbzNQ3y42nCdnDSZUiKo9dy3dYqdo6A/77v
6VoYwDD//77mPTpaP1AiVurUZ3wKNOWYXn/9SLWaFen2KWF6XjeV6tESaLlpELQC
Hk6kB9jKDQ9LBFHnzuUB1hRpmUDr+CNFQ9khqxFYoGQWPA4kseGyJoJLRXZ9Ftjg
e5QlSeEONhD5QDWkWuOjmlb7Rfn4kpbZ/PZHibgOofByKdzsNQtlhXJXG+/AsrqQ
gEJzyp3l+GhHrXDH+JxTWXzO8t6txwbq1GiB59EAgrY0LNU/rweI4tQLZHGAeSDN
F10B/oVzegyqEvrX4xT/KUys/2N71Lg3+edkp1KZagL+w3fRga17WOQywh5aBDBv
jngQ9IiQbruicuevDvSZlklZsppdpfq94UIPrfE0c1e757k+o7/tsjqnsuxlAlJR
jSnn3A0Xm1chrS602+ktYCPZJymtrYCY6RUJFR/y3WdGdmNZghv52/odDydwBJuu
cd/v2zamfATOHe8VAP5j3TioRk3zGjMDGUnt9PnJNH5v/kURsUEemall2QTEdvgr
/7xPd2dhwmqzltAzy4KPpfSSm45HMQu1giw2yivPaaoYTrAP3p06WtnzHgtTgN/8
6YJ8qYiMXywAe0siWkQ9jlTRPNLGkWEERQDKsvCIwv/Nro9upTHNOypg9beNVJ5Q
dqlo0ufwhG6Haol9cLqZSqZrA8L8Wlc7LQfDdQLLcXUgvCJRLdUELLIoT3ESWfSR
TWrQCBaRnGP9aqgR3YmnONPwgD28z2blJeRIVUeZ1iyl25b5PUEsH8gSdvM1BoyY
pjXaVxhdXBFwJL1LXvIiBWE2Dx0bF1HbrKEeaayluG+tlts+pgN7zpY7xFK2ghAY
5P79t5VpZvCwg1QVhl2Rv8Ywwh927J8qG6WvAtLnvTkyjZL79xJhHNwYRELwnfw5
6OI6Ymu1HvxT/GuSiG+4P1bCarztsJNtkT9jS/K5Ma2RTPnyhRNq1noAYk/zqFNY
mEN6Y9qhW2sJbLFxXokfgVTLxQxIdIDLZJUFaDKlL+KYHh7hfsiJVq9IBgLMRErC
KDX1JQdEHPyiUufDLV469nH8jYprVHpMOSdr1e0VJSTq4SKyxuDPhtaxmQNZDwjB
jePksSsPQU7NZf9ctnAbbFifDeU6oZsu0COhrkqmYmxuXkjBldGBu+aAtmMBVlB3
ynRlvaX2mYTuM5bp4/8ntP0dFYiGx4QOTFGpgAJScQCkCwfxx6xrMon6RlHpsZ0v
yGTC6tUsNFvsSUc+THkB7OfFfXruwRMMcB8tMcAmRhgPhAQMKLfypVnlcRZg9Xmr
thwERkEfemwafkp/Ae7SF5V7nquLiWJ5XtBwr3vV3Uti6ytUC8vWvbkXkba9oy0Y
0ebLL5SSZTMOxr+8wOkNjsyFX+6dzKzj/S8fV1yOEPOJXu1NW5hhr68VFOMr3D2t
vxZgv4ahyyZIPMLqmGHwFWh1P9u/dxJg9mL+WFHjBOq0sIZoSoaCZACNIyDeggr5
0Yc4m/2YU7zrsL7yh4KGwApcJ3IfoRdHRhN8NYHUB0bDnaM9p3HCqA45Qx/JhOnm
K/NnlSOWkXb6vN9+uo8/kQ19YM5fPygiIqgo9ePTDOK6f6XWsZ69sI7Ap4yHQdIh
bJfpvTXsIbOHllKjZ3FLfuc7NSMozmhfI+dFDPzPM1JpE3uu86eAfRiAvpfwgHnD
NmyqQGY4/Rw4ucqzCSoESjawwP9wB7GAijWdvF/Gz3rMRi/xJiRRkCEFEutYJ5Eg
6gW6CGEYxfypyXscqgK4pDgu9mVBV5g1FzVsj5TNRRDUBz2avQrbni8JtiI26qaU
rX2qyqsytBHcAzxOu/kdVoM4s+CHZcfAGLS3ISaO7FGLPwvWbDKg3eWw6f05ov6t
h8VMYAEBinv4JELovnyeBBgKIW89B5RJstADzQqbRDgk8lt+3KfWnTr50CYpjr2G
u4LzR6tSJVe+jiqSr8jwPNUhcHmMWkeMYmon60Rzz3HxByKw2xjmtF2w8WhhRwtV
FIvUiiINTebGonmh5CADjiwAeaMAv3w5UbnEIwxv5v/InBVc+K0JIYkiBlMZUMhf
A2mofF5I4FoaHYhr/i+2xE4wagFSHo2RcoxQQcby2JvGQNLjbYlq4mYDDiXUl0eG
zQQl/ZHgWSx2ZkAfbfD1kTJqxUfeUax7zrTNSQqd81Ki11JgYC1+dy9vKNCpoY8z
GFYW4PamMuK1uPaAUQ+LcFsxskVkF/Hq9vE8D0OIQGRm4/mFX/Pwwuy1FM2smMOf
bG7gYjT5CsKmP9Efha32/d17Jt5F+lcotKXd8lIbmWvLO8K3TWIyj3nx3ZBa6oc/
Adrnis7aY77D2xzEucC5Qo95dqkjpHsi59VJ0rMhmn6LEO7qpGTRDtc4W+JBQGUW
Z/e0Tj8kkJfLheHoZDS9vMilpOzYo1O0t9UfGWeE/vaHqgdzw3pPyjmbjWTqEl/k
DtlRR/ajUaFTjRuHDsjUqaWcuEiqYr1I9X1OdWezBV5Xw2oapHAqr7aXEjl40QlN
T21VNMqLKDQ4pu0CiKAHndWSOWoe5gbaF+0Kl+2CO2RzpzVr9it9oVeiz8xJCz6a
NPRsh1kqugJ3kxYUs9ebHA+ChYm2n773evYmKOtmNr57A53hPUt86QpAKn3Prpwr
gbDaKwS52SMuGv4QsGlXXq8pkeG7tP6lv9vbE0CaFtsIkFyCaLQSrCNCKa/T8s3e
mCR+h9LNJBD7dgBu6QiqA3K3Eq1MIajuNTpFQx3F8y9OeyNGPvPs7Gh9pAAmdq+I
3bNf37HJFhwrEwOWguxnsbiOnmv6j1k3fdrX0dJQvbCP8o7/rc4dHZP/Q2FoQmy+
Jplg9xN0WTejkogHNjmYoQ0l22EQMNaHIi03GqQzXTkbRwq2OEO0jWCTcsYD26+i
4l8WFo9mBnB3nNvW1zvY4eU6X+/W3r4sPpXZ0PP2j8m0qSKsJZVMTrKa6vlosOSC
EyVeBp5nexMqqsxOvzfB2S/UM28Fdl7z8Qt4tZM1uo6Dfj5j1I4yjDbm3rgM34AR
iupwZ2C8Pg8p6lvUdw4ZjAgTwWsq+aIUCkqgqWJcs6krLWFsGNgtnovuPKhXUUsR
LYh//v5KfF+r4uRBjb/tqVDMPmAJzoNO1eUhD7XdXEDR8blYjYTe3KlS1IXlyql4
hgXHzfBOij0QfwaABkoL1wQ+Ouo5pXKari9aSyRC53aFxXoiiPxLxJD7HAJjuhAH
5jlwVNfbgr/MDasZpZiLXeXjoaFUBs2m+7LSfaccPCjCk26nhYKmeJS9/5sh4V23
Nm9Kw1Y72chgA4j3+LyAsM4u0yhkYfsPLWVXvqF0oqn2OlkAlaFRGhM+tg6TyRd1
FNyrGjLnn75p2cKOXMaS0BCa7W+w694qk30G9Fs2xrbIqmFRNlGNONQNRx6+EFWB
+dY6dJhnsh2piyyz/R1uckW7OQP36enMQVxpmSx4NpxB+tTpIlopxJ8ovuWL/5lS
BEIZBhVOFDs2n+VYQxWDTzdyVghODFAsxD7IkEtNQPqMfw7X5na/I0QhNaJbIBHh
AcOjSnuszYhids+mdTKn0r7QAENf1wL2v0yjADr1mBPjF3Z9GP7HM0DZL79bSCO7
DsnS+h0f3qELsYEa5KnXxoaVCk7h6i73dlmeID6rlBuIvY1xScH4DczUb9Hj0BXz
VaW88c6Bg48uLVDo+2t0xoAUMkzP9g4U9DT7DKJmSjNTjThYfmixfl1udwlAY9Nv
VPNaXSKXVaCag6LztGk/CW8gxMrvHeWUzpQM1eLLpXnGiyZZ6KHQQ6bWyXI/r7qk
Vi/Eake3ma0oobZS/khGs6bn+Pcu8RNFubXfJBxm4O6J76m+4Clg/6LJ2ObFYeyT
jbwsR5NHw6RQY/v/QncXu5bCDg5G0v9cxsiI+o38MOXX2JidRw2hCfeZTc/h2HBl
QCXbrJTAwBMpwPDkwueRU+K67NaPKxIdTL8m0GcHeFr1GBbVMdTVZ3vv4DoNurHI
AE6Euny07oJkopA8RYMMWb2AmTZS6JpFRven/PUOPkNmRG9Vw6W39m4E9Crtg/pT
iLPctQUUzAHvk195+pRSct57Sf68tmWlogwojZ+N6Pbi9Gjyb6ZQ1FkS4SCZwzea
oi///Cvcmu1Z/2+OK/fTvk8w2L3YiwWyjHKM+jU0vnsX8/ocfytJoclG0q6nWLhu
ZLt+PnH6bf24ycsaqV6w/pYJNwM076JVbjLX9SZZiu4TcK34tcCInLnrLHDltS34
oI2P15kgRoOwy0n1Me6xq8XJuluf1P6v2Ogg14W5nAHnTrICxP0LexhxXMA8e8w+
+IyEzMu2UIQmyKWw/6aGMbvHwURPRVykd7CPNZAdEKZFOBxahOPwO6zCYFVNgh+l
l0LWewKtYia809NssUGdAXkFPhMHNSa/2pL0bJavW3Lhja9UiSoclYWbGEAjZGGL
wHl6CqmlmbMQHhAvSyqxizTCvQ1bT/OVT1qvOQ2FZ97IUdLPhHXedG5y4g1IllSU
AUwOkBCRD5JApfL4uv9IlKEZ83i0XUUpNlAZZfNRCgFXg70Zkkp4xOwCAww6ZciO
hn2Wj3KJrSvFjHZzKGg8LH2Bxu4XydNM7nwLDOt8beBrWTJw5RjHgKrB/CcL6WhY
7Sl72g5fSQ8G6U/rzoLfIb4YilfzGxoR4aA7f74y3StHmKPGCwFcTNtUgNro5nRl
H7aDYxwz3RWSwwIZZpZBFHxEU2soG1eWPsysacqVd6QsQGtFqPUABCzoVWeCs/xA
Xd1HR3JLOdWLH0MRusVVj+2cOjXv7qJzhmmb/q1geMATwRBof4UN8+D5ssE0EXjH
UA8wuBvdFXWZPZHaTVdVi6qkgn/+vNU39B85bLA1yuujbx+tAAY2yKbg8Dy+QNGw
T9KyjZcKbU/Z4mPo9ytkH7kJgiaDXbmP8oOnmO95mJwR16CKJbMpQIcDNtFHKGDV
wthjFyhpDejlstYMHtCEl+fGJcUjyngiR1i6B6rO0ZrFxP4k8eifdfNOmMzjw7l5
6NhWuupyo4BoMwfLJDZxDw+uoc9vGG/oczmrrzt/OHLL7L3QGrL8wy6aVOGHpBPt
8Z+o9uC7GHLtP1wJCNLQBidg7IyqeZs8Tm0xXDJBke8NCucSgaz/ZhtBbYTVv47P
WR7DjXxzCvZXpQzqER/qOvmk16DLcQWvfKGC0iq9fb/qLJ7tRaRhxWi5Ew/w4w01
E9aXHzgzmlgk3cPoG2xfjQ9A0BYEOo3SsegbEVUWDKl9HStMVYWFwqz30sw5L/gu
U7Yn5lWrxWvKniRooGEwqDWKKFdq5nefqkcg9+4xFEX/JwS0Tm6J2bBoco33oAaK
M7COSYQ37Mw7zbz78DChWNCny0SQP3X4Xpsi9iwItVUf/PDiMnmGjbP8UfT+6uWe
2S22LIR7JTuR/vpzie6DLr1e855VIWABmWq2vAY7J3A35sk5gbfbWZftGHXy1y5M
lYXu/+wy1jHHOhAM8hF7uEtjkWTAlXyQiMqboEmgE5e71/T0tpH6UHMNCaNhK1ze
bgpbk/H6IxWVrUM7tKTLGmzT1nEc+dgXkGCYLo7ZyZjU5cAnUneabDgELvDmTghV
PPZzv1YSbbikYc/XGXxBv3uEZIj+nwvi750SBhUI3kvDwmluU14bgBEDLSsvcYQE
vvipnQ8ggx2yWpSdFcmBkZKHxPY8dBjdj4712x1Pof7FgzwXVx5F6wWpva8BPJ6U
QnMkV16IfoImvznCnf21FIgh1xBdy5YWNh3i6PciP4Ico3QkM6402AjyHNSobC+D
ZrFsuGVTS4ftCX63gZs5NQ12TXuj8NSv+Xr/jQALq7d1USJD1CMXWXeDT5TE/Ll+
O2fKLsIxDVyJuaxWCjXgVjuvbw2uaM8rW4scYc+KG9mNk7jCyZVyY9xVeZdVFrMd
4Yq4rbxUNsRYok8Y0sslDMIQuGoWrJfelF5aDpOXhHD51JVOndVHl073nwiJuvPg
tE73tBn0ArReOV8MsQQC1S6mk/hlajR9kyY9yANmUC7fnvTY9WB41I4hpOTcLYe1
04aTGfRnV9btc5BWUQTyQnvxr+sxSMghv3vRLrccLRfsmsvvx6RFCd764/CPHYsq
rpvb0DTuZt9GbY5yenmAuQ94sOeq9xmqZhvweRYOFeaEiIazkz8MA6LY6y8o+KM/
Mf4MKP2P1rFn93kOvBJkH9xyl3/lmI4jOw/dAQTs9tG9Ob5Ci8W5yLXF7kMgRYuv
WhkKzd9I2sMakRteeGWPS/PT8ZGxPMOJRzqVOfqdq9GSQ6JyBBsO7iPM3L9bW3OH
J/GEtO4oEA1++aC81cNeguzZsv/laLUMyfB9lxCiHTIEtiFF3GEodapEkhgASHfd
AwgQLGNPmrXCUPaNTi2jrIH7k9+KLY1I2VzHLJTniNfYCnfnnV+i6qEmIRZtiWuS
cuOIym1R0088MaglWUhayEpiZWLzh6jhd7nGwXhPJIdJAj6CXZNQV7QDwDMcC2B/
l4r1YCqj8PUIj0E9r7r+m6wX7najnh24G9Ol2CZTu1qx4wuRyLYewhRrpi3cAabu
5Uca9WhN2/nEa10ChqJfB8OtNH+4l/J2YaSX23kNXXUIdwzl8Kly9vxwCmVbYRdZ
c7Uy+c/uUK/qnkrBWFdnjQx2vGkWoSZlRVKezQJNKrs5TRA5jVZ1DPC8ir+vZ11d
gAXpodNkDbcuPe/i8VmlyrCEl0aRC0kRzVbrOLNfy0/aIujX+4n96BXBilxXSatP
oEuZbtAus2nu0iVh1JaIy+pdGCzPJZ6c7Mi7YTk8ABWqds6ezmJnov+owHq5NyM7
8DF8wNaMcPoVxM/jx2FZ4h+MkQzTZjhnSBygmnssvYznQcOvuOXcdeVZEvFtPjwl
DtkRCyOG9PQ3y3ShqX9SiM8iR4kyvW4papPsRFitMfgftly25676vKxPQA2KVoma
27QSWj8Q+q1UAxPMuBmodWbpYlFMi28QWmlMl1KKUp1evmy9yXt0MqfM6KZqJpF3
TUJYLanZHBqsyGcLMOp5K075Tmc5Dkvk5nT89f8sEupo+2kwIsA5Bcpjw5HWSQKu
ErhLCwfHIKKx0U1ximsdblvta/m3XRINwxAN0Qd9snqe/BprQLHyy+l6neh/lrsf
lyz1paxBMAN1TVzoCIa4gHrKtuw9DtCh7TpQprWNkg0TH9pQ3JrC6gIfgWkG0hvo
kL3oshnAqbrdMELuZa8OzcLq61JYOHHypY34+YaPn7q9kiwaeUna/QO3S82PBOT6
StHusFjgvBtCjWHyM9Em+ooReNMlDg0zWEGeZaZMOUr5q9jsZpwKXdRzVjD3P7CG
xK8El8a1FkRDiGjNZcIymd85u+eMIeypUrbwx3tg3+vTmFxQuJwt0uCLiMDBBPbm
vddzb55jutKOoRIcfZVHScnW24b7okFqfgTTsWZN50YUzUROaFxWzN5jmW3cTTTJ
TkHzXNzuwlRY9ijDdagNyW9jgoR2qp2VE44+QjcHtY2siXMIKx0tvl/hVqyQGWLf
y8A2OkDk5OHIwl24twZP6bjcY38nNhfqpyI2oX8Ti1K3QgsdDM342FsVgeqYW7X4
i5t6+JgKrMA6na6pXV38LWL+uyhyFuhS1zmSapFcebwrp7OXajAakXRIyI/4SS8G
BOyEJaPggSXI1qIY7sMOgQOb4D2abiyrQYCtZKTqAYRzYkry7E5HHs4Qk4CfuU9t
6lctvZd1Fr9eoWT7V+m2IsyPYivhoTlD8tp3mnrm716vBME4Fc0M0MV+3v5IUvJ/
ye2OX3inCyGUR3JckdX+pLNdVXS8iBytgOnS2YDV6gIJAPvWtcO0C/SxFRqXkSTC
v0EpzlmJlbcLfzf+3kgZbFV/i5qhIBnCxQMyC5W5bZO4hdWCNB0O4XVgafl1HG+a
yD2ocBvwVGjyj6RLWJYqCbBGDdi9BHDlv1L1k3kaVr2aImGRc3v3WS6agWIB4gIo
WTeWK+bHhi9CevN1hBlcT/u1XMcdK1jme+ibfNxaRk9QaMfHrUCqMKgy0ZCX4TJe
CJpcArhXPnxgqih8gN610ee8jFR+cr9H8+SYBm48VdyKPSaTyZcRjxqoom1/lDOt
njhMp4xYjJqza+dsTGzIiwJW9ByAYUlbT/Nos42DXZuQreR8rt2TOMBhvbKqoIRz
bVvv1XbIFMK6H5SZVG6KyNTUXQgB/5jAR3dizZWMYaRmS7XA3KwryUzEPJ7+4xqQ
UX7FGZJJkb06NWSf372zzlreHr4IMTzS4lqIEay4tQODnt7uVWJ/k7LgC5VszGX6
GClQUTl3M1ps8z66GCd/Y3Q+XNRfNF7iSsi1nSuvF5XnviuhW7DhNs7IVd1Q4jAU
PQXhRcyYpe44TRUuJoiSX41vfoOaGYfie5PQXslyJ9fOmESjy6gZwiyAmOW3DoUM
nA7fChXM0gr66uyomuQ7IDpt3OkbUllm8UvQuay5+g3VY0lNN7mAvjgWTeITfHEE
u84pe7ipppwQW2cviXZVH/0hapLcH2wiIWYUq9u9CjoWliBRaKYlNjJKerPjbbWu
+AP02RtwIfeIe4lMMx3PsKixIW7Vid4l0MMQ9KuW+qjF6eYTwhxic1lSPRubMBkD
+JsBaWd5RXnGA2pfewc6PbXa2eL4NQZdqfXRaLOmw1eYsfIh69MY49s9PASonA8v
0Ne/DPR2x2oLBQ3vDM6WNT9XgHeB0irZTKlWNFxwBhNjSuoQMUH0iipBssS0SRVi
1DqvA56UJizbGzW2Q0iSsIhv0Mln7wj2fy1//XvWr1tLxPzQS3aBGx2vV2If5inX
D7P0BUlEt29Ehnly1al+Ul8yi7+memybYxlESaLlyvrw7aLcdYGekK94f33wb5kH
elR3wsdGmpDrjbaR1q8xsplk4ACy/6KtnIXWpahsy8l0Z+mE1cX+jDtXyp3R0RLb
0PoJ9cMe/HJ/aPI8s9z8xhLvguwCocBgKk/H00jBKIQuJAWOQGf2FB8TWpz7tj4g
PDYSgc18+vNtxSsbAEcgDUuezQC1NJ/CGiIO7MXXvitDuFlagdSH8OEHItFKo3xm
MtXEBE3dbmFT5PkkxjeIRTKgwojGmUfUlUxkrNVu6QGv4VVfZQOw5EbwPGbEbgqx
nITS6xbwg909s3yQyUe6OyfUldBMm/wkGUAARcy51K5jLsA1Ub7MZXyIe14AJd/v
4l9PaL8atUamOMC4toap9rS+Jn0YyfK4J7qrhk77qrgm1wJv3Y0mV8U1hcynzXSO
AIgJLruEZML0vxahz2azzojfskhPO4xLGP5T5i6pZQdDBvnVpvMQrN/SrxOwVmxT
dSw18IwL/9hCNd9rqQW3PBPk7dLseoK8BvPhttBuN3mStNc0ryTJIs6FgyFKKkEK
VT1CUrEbhLs8zfVFP7zZwIObWluI6WjGlU2WjajcmV5DpNI3+Yx71T9hAHwYpISM
TGNKw2O2r37Vc7zV0RKV4RYU9/GID6WPtLpPXzKMD0NzeCZFD5ThjMmHwEj1gjct
DL5volzdWP00FKiAziSQ+k6lMMCiHOKzZv4cYQIy/5L/3hz6Jhb7m8PdoSjWPsT7
fn24r80YSwjISRt3ESEsOzvgypEQh7yOh9jS6Q+fKjXMqRAudLMGrpbEphEAdAqV
JUoj28VEcVVPOMAUHq/MIU3vXfEffX7b2CHsXgVCb33KjLiWL65lsD3cHBYHXCZD
FoUs+sOqDymC1Cpfh43uLaam5MNbc7D1eshmergBgIvYmvaf1N7SN1I8PUuhnE/h
FDq5uIljzLLhCOQ15L+Rz2rgoByPyjLnpf0DSb2HyjP9TjC31hzanWfmGXN420u/
QeJDhxibD0NZNaC7T+Bd9vUc59UezE+WxAQxSWDNiHlihBxZKT7MPQKUrYNy3S3W
62JkD/gYrbrcalua4TtHo8VKLT6qCiZmR4P1li/c7UG2zd5A0teH6d8cGtkaoIk/
h+P+cTIoj5lEiBj//SF3BzoCrkQvbmuk21bg/entBDQuQQAZsyf/Gbc7QuVvJrUk
wITMIwC4E0o2lcQJw57YuXCCnC3T8UiQUfsZ6CT17gYEg7NbTWezy7W5WIKRC05f
yJ6aw8N4LIMOKgm18ZDGNspeilyOwfq+75GVdRR2TPabJ0Yc1G0W5NpFc0KMt1u8
wBdAjuLH5aJ0tfsggobOjGxH7uHq/c4AYCagAPrXJKYSDxo+wHDzolRrsP5J75r1
qNwL7bwkcHGRubzxYpMuDOyqQ0uFKm1U5KIEw01Hnh54EnJ4jKPx73RXVI6fDiz+
Py014+NoefLz1oK3cYzuAxv5FQ9XJtpcqFnz7GGIaFRPT2Ai3PaqTVaZlJGS7xLM
08av/21WvrHPYb6Lr1hODf7SiNac1HwbPqA0chaw0Wf+TX9DCK+DylA3rdUfWJH0
sAew32sO0b7+i+2uPkTNV4N6miRNjkqBCvBeLkDFs/MJVYM+Y8oQV3VILzx/N3AX
uZrRkhm/mhbS4uiUaA6/9+oKT3zAzSZZhb953iu7O3Gx3RepvihXm2QC6Oyr+kY3
aHHPOCTiF5lK2um9EjP5LfYUV/PQhrTG7X6H7uM7fFUsZi+/e9pOrWtnXXx6huS/
LT4Kq9aBbvfzCqE82yBCLw3XNTJx2J2Ugk80yfjWdmE+DYRTqRzxJfzyQM8O/AUj
SirA6lzR0Y39UNWJQOzJ3BXRKsTI+giKYJGqfWXHTNORLcqbCfbYRs866kADEny3
5VSbSVwbFFMMFLLVxTBKw+YxxhzUPiDFbQEXOnPQ7vO0qN4dXE8ZdgqwYR+ai0Hj
C7+3Df3SCwmDKEla7VqK0EG6k/D1D9OuZ1+hlHxrsi/hrn3BPDbFYRDyhwguqpKC
y76IJIfv50/2a2zlTnvtcIQLXfKtc9Np0EB4z4J1WAzUtlTdVHQbMCkGrwOKWXFe
OaczzLdq30QZLQ4r5gQ0heCc9nn7ZhPyM4aOuz8vgKTEyVyTaxdqOTacnPBUF1eN
9Sqp0gohu8vmpbqCJOw6e3G8A9mOrFCoSQD5eq8nsi2sGZEHb9WiwKv7QjGebtCJ
RSyn47Iy2UvtO+0OF9s3VJWHvKVx6CCtC0AJO7YUGkjafaAplH7WjnHGSXvALVH8
B3FoGbM7k8pjvLvFCUzCKyILUQ4Y/ipcmf4r4ouuIuHr3u4nJ5Kwa0f7QCvEGQNl
tSLOEkcIVuqg9bGQ7sHu5K2GcQa3gzQ5Gzh+fs3MtxYYcY2Zb94zoxUjuaRk3yH4
idtxkv0izFzj7kJQwR1jRSjJ8Un7LdIU7gWd3La8Mh+WhoePK5ut2KHNJ4v3z0iv
wzuJg0VAmv41PN8rcCqbm43sQIH1gVp4suS9AU/A44XlYcSdW81P+16Ykn8UeHK9
dgsKKj4hUS49SyJ5OpXW5saCiLm3yyflrQ8FolI8ZLLoSrxi7m8cvhxN7+aEAIea
YDJTATgyFJjgDHh9HSUq2fpAgJu9gL2g8lxKpYhvCGa2NV8G28avjbHiCQ3IieFI
4Nax1ZdRrZj+rQGdD5tVERI4ed9MpMwI3DNL09Y/qkdPw1kL2NfD6Moa8lea2ioO
mlDEqVM8hNrq586+v2z/ddvdUxO1OP4RQKcGjHgk2PippvaJGXS9Dzxa0phOeeIi
rPyTTIKUwwK5dfWEgUuaV8HbsLLfYB7refiCEeezTgKcEO6KwMz2FHvUkLJpBcfC
XOqLZ4QUr6N15xARXRtu36SDCpbe0hUa9VxKM3LPdkQqXoAqXa1BfuKZqYWL0IBg
8Sm+vB5ZmtpguXjakkwnTm08MR62LddPr0MtGR8Ymfb1v4b15fSWvuV/iR1iuWh/
AFcqx2TEC0QjxAwjeE3JIk5StV3Vv+cgOKElHkTsMCc0HBcB7LN1Dz3YoqMvGhtR
0p21rQzD2zPEbjlqteWeUvGayZamjaTU+k3eF+ZO7OnZpDT/SMqcqMjtuX9uYgX6
N1i8w3QqR45cABO3p7FkCykufgI6YyUNGPBpYpI61yxFN2B3sVeRgE4zsghcinoz
8I4b0HWnINdfDXHldoZGnz25x4spX6u2ZHT3IKO3kRxNQv+EPT++yclZ6AdzKY8J
fJmNkAnS8Ci9lh7ANKpR+pCGadhMoJRk/tQMFaAhmZ+8bR4nj3nWISWN5Uf7DAtx
nroNhCFInlyrVQofFU5DOhAh9bcbwLbYkFZbITrJq4DaX24nLCtPX9iICafWJ3Ip
043S7ifieryhPkBiGrFwRPmaec1v95A1a6noabLXiqRpm9L164leZARfvUHby5IR
unaHoxsIX0dRe4WYG5VgU3VJcAl1Kp2QQeb6dhs3DM//80w2X2WbLTZk+kw0X/az
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
TNGn++9nS0Bo6C+3n5ZMaEvW8+3CD58K6GA3VTL7wRAcNc0OyArAIhgDiGYwWPIw
1mnLjwR8kjrniSa+OyPNPKxnQmldu3PDzD/QnUHwhBvK99D2x7da3vlm6KpigtDa
pgbULZMy7ye188BdHUXAJHY7/YqDbVDfzygctW3Uwpmf/N3VUs6DCMv46yDdtRru
fraOYEAATDkZA5ZWvuHrXzIkxNUTY5pTq7J5FFO5MxX+PSiQpt7PmsCc6vj7f7i4
ZN0GnQw+eb8qzIlZzD4OlJP10k7tVLu1JLkhMH6dNflsaxrloVxnc0gDj8L396a2
C1fFlv9MhMO+3lZg4MZ1Eg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6256 )
`pragma protect data_block
9oB9PvblYSbilOsTCFyqYYcxaOBCGIqUKzSQO1ONQWTQWgqbpT6/cJ29yd2T47tg
4QBatibEp6mR925fZMdnC69MAmfjInZd+0H+IW6i+4jDXTFaHUr33Vo2DzFWR2Oa
78YPD/yNGnhW9BCv68kpeFo9wEAzI6+597Kd5G7E+YD+jOL8clvwnJiBabTyhcyB
JZee6+jnyeba0ojuW5RCKWNJuLFzI2HDZUVr6BlOpO1tEE9Cr4QW9C90SD6/gTNb
NwgsyLK+gMnv/NKUTK3NTMc1YLAlj55gjY6HMv9qtPb4yaGnNlNbc29uebvjOd48
ojBcSiZdTPYZLCmkVCxiaKaBfoBjM9ewCTcDwiyAxgUzH4BHBn4nGHtCLolIc9Z2
3YOP3Qbu5Tyj0YuExlwsdB6OAIGpwF0kWkxcpGPDmzfzPEqk0QK9Tr94NRvz5SLh
RdKtTcQfhsL21z2DRUOHfkicoULrfXmu5ZbydDbHCfMIvs/PF5SKDci1+T1VBlUl
DuH7q0inl7+Qx1WfNIlLV6eGAzeLp5y0CIgZMF5PHCpQnCRkdUD79k6bQxiSeOSC
zqPlNJ+Dpi+3DCVkU0Ph9oMjAK2sS//8vMw6LDPGz36laG6ueKCa4N87LNPlxHyZ
dfJvK/y9MFTMf1bbIQd6TI7EgOvf293tcjjeDQaAxagQwhZgY+xtOy2CALOMTQHG
4vEamUrSGfFqMPZtyblBHfyKKvQnmfasd2LqMW69Exe1EpPnfUlVl8UqH0zzQEpS
vzoBy0kPe5eNvq9gohwUD5ZdLjB1hBg1OSNOwLZaTBeDkWJx9Chd+UxuV2ReTL7J
c5bUVsMYZt4gqr3W5EkUErmraVSUYJfp/TyF2Lw23u78mS9kMUKJRRMcgdxB92jN
aLEwOTbazu19Jw65MV8Rva7Ks+pWnp1bMVeOL/P44DSyKKNvYZ3174+el5uY4Yq4
nAXxGUHQcOgYo9GbemcRSWFrA4xtqQOxSwKc1R+z7ZS1VzNrQhWIqevbgiZnCbRN
DXKDtKXUpeEdYx8pJBJllct57081pajlwaTghOZmkZ2ttvOxvNqNDQ1plSTi3j4G
+3rIDS4+2ptRfFSlpxPmoXHAfvVLtO/CPj7yKmGbt6dFUV/YX1mKIkJtK3zpgLJh
OpupzModJmibXFuBrdUFerEBJGlOjPUmQeQ5lnaHGgbrFODXA0vfLhfTtr9cs4HN
ZSM2lHPBzrBiK713W59P1D4fCVHHugoN1tVg0IzzvOkx1Lt4PX4lVUt1Z59k+GqD
MQbze/8AF+SXNRkjxMyFcyl6TK/KCVWQqvqq6xjrjeTuUBanO4weboYeOVlLYOOG
c+erNBSN5bYPlYB857uTXidDglygOmJZGbR+0hp8KdJctXXll/OLYYk1+jicEqLs
Kw00sZpxhvIVF7Uuxt6PvwnzEj46SdqgsdRnm0+/hkXmZyMVV4+zDhwU2dHPIbIC
Qv6UbTWwcgbWvwnNcfZ/uFr4pV1RFBel5ErxQ1It8PC8a884gHCJR9LtsEKiezgd
Fj+oW+MGsItJlX9KV47eIBwbLK+gyvFzyrbXjB4ouImcqR+FiI7Ddppj8x6J7CMG
bt2sqL8AiO/RGhsFrAuRCR3dm+Ijdny5iKd2Wphdl+1TFZLEQk2gvLzs98Gb4zU4
80n1q06EMLp+54bZbOvFWCXYMy1zfeu5OzO1Es/bWtrfCOpOSvle8aeOyuDmlHgY
fJ7/2MRtWA++XlF/jg83Jbg5XBynp/Vbu46qxmSIwVffnQcHYJTHUPsCtsYK8n9x
C4v8Jd/ai/dqb2nTVO6/GVQ0slSbHGogCaqTKaSVslzd8exiAuYvwaaLTDGvsTri
1cdeGi3bzAxD/O6uaCUK9HuyrbLq24SY5IxbXWS0lrU5y+kWgD0MYwkYkDQcBdes
A5F22pi+ao6wAKdr5B5WbqpQ66bxG4UViIT479d7QMzI4fRSeSz1o0P8jKF1fVzt
gq4iQRqIzEoOKuR7S17FMJVcQg9e3WQNuCuiOgV6jIjMa88HYiRQCHosQ/nFD2Og
GfFADXekhsDxUsdwrY6+eOlLP/Od4UsAXqHt57obr3yYHl9G0HxrhxewvzXdPSRC
BKgampzY5dYjDgiIWZgvFjD1DGIXYfK4C+SI1SGadFak7aS6ADJJymb556vi11SO
934PRJbLrv942mkV2cuWZ83L7wuCTCP78f+O0OcXg/8Q+5URAAT1GPFxeiXZ4WUh
BpC73adPWFk0To85Q4phR+eyHcy9uwBWlI39x46S8v9wU+SrkCz91HV4Sf6GS49+
5GcfAvc42Vrr3Tcrb+phylUXQY7m9IohPDT+QMC5OWM+WL3PHqXIYsxENytYVwtq
Jn/aTjs5wAZzaW88CxBNG7dJCSnetnGKhHyd+wKmUTCeguQ63Oge8s7B68eVLzdL
vFFPRBoVekz4ZDKcFlPgeeJXIRF8YrA81taTanI6lYuisFE9GTgLNxz0hN4LwGDn
c/zhZArd+/yiy8XYSm7FNeBK2KNMcnHHDfMCrPcTKsZGI/x8VmAII4kDwN5HxKkW
SqGJiZ+/2g/tqjCE1tjHCiiye0AskpKU8BuYJpYGD5UG/eAAIpQ+aHO/Hm/zvI9R
Ka5pOca8lpYUKDhKatQSuNllywdeJyC2zWUGpBCPmGJFqk29WC7XOV3rH4fk0PFx
zog1pBxJe9K6E8w0FPQCr68CAFL2f+c5h4o8Fb/Aw0MNoq8WsfNLwathR5gybADR
oEKMZft2OGqRoOpTAUWjBNGbvyUSI5xNQ4TqPH9jmUMXgL/xOe7aarkVlMfRR8tU
gV/xyI+lLldUatRDrkLfNCJ48ytzP1nYQ/VObzVaV74Yb2Oiz/kWkWp61pIsouF8
ASBneT6ORpZN0+Bph3mZ6bH/WnU0fmrtdexlH4/jgI8QhD/D19tKxNIy2DoLEDgp
WScMPB20vHPUt8WH+raVCeL8ZtkYPH8ZUQsCtkwkVxulRrmJXuFTMYYCc9Jd118f
mqjvXOsVdz5MHtjC5/h6nxSKKkX+z/r3bi+seoHtIDaC0SKi/fLdtDLEGQ5tzWXB
Dp1Z+LSZqgyEDg2yrQNzTKoW6wKMlz1bMe0HlayScad7Oo9JGO0Ri12Clid0PT2O
1hsh29BrokeFE7sBXrHKxKXMJEDsfQZaysORJySyig7OSo0cDvjSMk5o85iBmdGf
HFeFgvP04ioNfJhLILpjkCuyUJk6bdw8e4cKbwXPGRur9a885vtRqO9sVx/iuhM0
A25dgLuANO0Rkaob7BXSCGJ75DrEZFAzhgraa9a6k9noC9LNVhNOOmg65HHucqca
8LLw3UdctTp2svcuKvD5DQDzLxWQKB5Cg19uk6GULQdTGLXqKaY+672NL3N5I5/g
6WCfm/q6ES6EcWWFlhcbD5UI9bIxgMtpL+Qndk1Ogu4Wg5dDx0yGLdtIQzDvoc2n
n4H3az7pKhZRFZQAinMRNNUwinDjPihrQf/19W6Po5mmskEhzGvLvqwp5L45y1nJ
JCtifx0CCJt0AB55iEueBMleHwBQdm/YlhwwfLhbB4byPYBh9Sanwn+Ka1N9G0e0
7iAQqrDG7q39pjqB+zBgVjl4fXHop2x0pf/UFuPxmdkOgY/o4vm7WWEO+BFr6aww
PQNSUPuIJKPDvqxCWL/kM65VCsC4/9JS6BQ9ySYgCYRtHZrZbeAVluoxhaEVYNK2
THEpa7pnFPo5qdQRnihz4O2z+mEJSriupLRAW11XvOCiUB8XnVV8pUQwoLhbZhS/
kXKfq/4nEeNQUPDJEtkMXaR1buCeP/xu98A2PFRqqG7JEw3TPg/csN8Ur3ryFoRd
1QS10BibrD1P/ysqfiok0KtliRMB2FMtmZjWSRx1jm330n11scKaBHAvrI+j+vf0
2i8PHd7MZJp/CJb6QQ8Mafw+c9BHVVSshw/y1vmhrmHuD08NUN4I3zY3KHIXjGXx
cLyQ8guUEedNQ2CIta+4Zb8RMsMQ9MDc348rfr03wvr2rDHkS8ltKlR8vGQ0nn/K
PPsjGzjvEPXKZQTOasPtVOHzcw37GHQFTZCWsHAS1T4pybsfCQ5CUpt7y7S3gYNN
4ih8FQIHyOitdDSa+8AGo9KJITdQQea7YrPy56awPQpJCQAyGSR4xO3N/vWXJ/8P
sc+XwmIX6TM10CkzW0E841QG6Mdpwr9Lzer2hp4KBzdNQ8wxLTgg06CrGGuajq6C
h0/zmcV5BBh39tvPjd17dsCq0AeDejjlQOPLxOOMtqGhyoruSXjA0Q/XPJqc9Uu+
o9Z/xbqICXCMsMiI6Vl7lFxLZX5SZ9bAHLXzXrYrjvgRbFe1m6lYUaxQsn1wOZo+
s74+8lc317FyFsWJknbrTHRk1LD/OOJ+gT9GBODEtMqhYxFB2qpEKrqUHcwHC9rk
DeENMd004y36m6V3bGW81Ib7hGZFIMdQyz414sc+lUBbBVtra3IQE4mfntcv8O/w
ezjnWb08ZpjUGLcf42cxjqop5lnVioWek6JVYYkJUmtqpZ+iMoh7P9OwjsOOgkvI
Npe/47ZIEFzqvFFunrJ44Ezw9kFGx//TySUyEkUtMNroY8e3/AU4XtBOaIoXoZEt
+D4Ujbbbr4xfINNufsbhVhPKJo3bujHxxkwrzck1EGR84k0exblHr+ctuyB+QU/K
cCEScST6jgGDzxEvtloUJ2MW7CVgT3atnANyOm9dEczg6ocDNCadoQ7IF9KhxWM0
mMSDFMinFYIbc2r08IL++WVB3I4607qGEg7v/bj8THShau13bkoRLKIERuRJ0rpj
WAJc+iu2Jy0yWtU5AebCO9PFPdDParasNsxJuzV6hzR6MZfS1W2O8jpdKgU9Pkih
e1eqIlaF18dBGxiPiS0e9hHVUv3TBh/0mzj8TE7mZAz5TL+aXCQaVnAfIW1IefM6
8XVoSFgjRcyeFxb7lnDjKX7NL1JBYI5MBVmJ5F9YCWxNDXjai6Cmqq+axol/eF1j
kEttghq9JzHqWNW6KhkeGpf3w98+Y1tKS586riy1pxOGgxMxuwrX4XuylUQh/5Ch
mxMt0L9pBG0HGeISLv9PFRDh9UTL+SgwDf0PXA9+lwY9LAVhUMgcXwRdLK+2HYyw
0fXNxBasEsP/6S9J7UP2WavLWkch1W5hpyDycBXDplpQk3ZMmdkNt6LbV+VqPR2K
83PZsXdQSf7tDcc8jZ/orNI0QuNEkrvJyt9eIxpOlKD/zT9abTGxAQ7o+A/sMZe3
tl3arWSBF2SCnDULOmhIQ6RtUxYnCOIwdrzAJK2pSMfVjXg1RQDMNfxWrOscGOQV
yfjLK+qE4rR8ccIswi8n0Xg4i4mG0WoBnOa7zdWB6svDyMqFJP4DH0kOY5V2WYWN
v8AyEBr6geei2AdhYXr9jK8wzmTt+G9fbsf1fsB5rGGld1B1qYYiANHpSl+P9Q9t
FGnP92JdmfpaTCF1BFMOvlYTDyQqWOgZdMjB+jgWpzBd5mM0/KoJOfPeCccfnyMV
JmEYr8Lqc9fDDc9zfkK+ApCAllkZP2JE2MGC/VvOW88Z82e+wbXcUZPEHhsuRgZH
LQn2hMjitwcJzwkIKVo1i7dIze7DZ6iPWkKkcGN1qnMNrxVrCOM2DNw7OEG+HFF3
V4FU8XWMCTExPSwQeqqzv9H/i1QvUYiD0b1xzJ29+R02XKBcr8WxtAaisebx6L55
iEds9XKBh45ppZbZIt27XMHEVIjr+KZceONcrgwwuan0MD2I9Ed4+xg1gIh5+lRU
61KuU07OW4IJG+lBQzyweyEf5bKsARbkZj8VFdr2dyKx+dRirh11wvTaZSWa4sq3
S6JxmFc/kBJ+ipRUDLcIsEtAqANfCv6JND8moi61ugEvz4gmK/PQ8pAP6L4Z28UN
TUlHKsyNLkke6Kjxk62q9mOKrHFjv8hMsPV8DbVZG/Ac2LNxpqDqBoZ7FjuCmvsT
0dC4RxhNWBvf5K2SOMqHWRIsXv3Dic+Cf2rqOiYGz3wXxqYiOjLoWdScI/mLZeru
n2VmsYHCaBxmSsa7Jhg+bslZ9tS1ZtdL8T/7Yx9uJ67Z2Qh7GXchhoVQxL1+VOO6
7tqIo8mPZBbHp5M8/E4dCcvL3sOGRY0khyN04BcrXnTETmgIFSLwc+oz9Q9uUFxV
hZdJnAJq095wdE2CnM/ESmUMsxSySvLtPbDlvyImFTMf574ADerOjXBQYbVtqhTn
+gwL5SfZBXLcdUkJmgFhFdjJBaKqxGO7vs7PAnCof3YArYtPpS/+q9hBA57XCU93
HpCl2he9REqsuHbfWG6d6IhV35EEOgOZd2oaqEqFjRH68tnbXm7f2rfCGlaukN27
Ul8aYlKldVaquU3UN57KTKM+SeLfPSvyTpUpGvzYAR5XYreDXHAsuC4/3Eb9Liiu
8uZS72WWhnsGN6aVerzgorHmanF8GqbcKF+WV/ZE8M5a82WCir+2dfJw34A10ab8
Eqj5NUAA7D8St4cZJRAKX7Drjo9XP5GU5MeyobOzDxbQc5isYUsktyKY/BKwwmgo
0uA2e1uhTog2G38Hq8/ReGQMGz6kkKeQaINTemyvVe2mr/lTJhVkpVSIYEQyq7+0
fx7/A/wadqf3ogBoLGS6FFSxmkbqiYMdaa9kUva0AHzj5ojE09mZZhyrkifoGT/N
X8ym9MsSBeC0D4hdyi5JXUjqi2PtF6pfBXnEYEwtIaEje2SezNddjp8+KZd0wYDZ
XSaJ3GR4QJNswTBwNNOUmyrR8JVqeVTgNfDPdyUmvDqhk7V8ccwJDo6yaRlBWWmw
+lYrihT9mrCRxV7HT05JurBpLAHJZtNw62j20e6fV0cA50nVSQQ+EN1hpNbkDpI+
lvT6Q6kDwMxlext9JKAMYM89P+tr8dUpX26H++Iwyujc7dQwygyJCxQ8mOypOl/o
GUuNSb4hjv29G2MyGil6uaa5wAUdp0DrDiCM4gfeB4KZ6jjMF09BT46lGFWyO1gv
GQlZHR0jDkAZnSHvlYFBFGSCPhAOeYG0TcJrNGI1k21HgKMIcEkuEAFIWRPJ4IGN
iZyYaSNqYLbe5Y4J4RIg2qh6Yb1kVcZoKjZN/QNyvu0abR4SmSWslzZnnU3Fgx8w
bCKeSIR3nP9GVCheqgiVRBxEOup1fxkKD9r9m4ZqUJUiYojYHXI84NFB7LVP+VXP
2FjdoYr4PWnZKxSh8Gi258JbK3tHKOwOLEDQuqrnxla8lN0GYHs3I/WuxaH/jPBM
1pPJ/DksZ8mbx8dAeeuHczD6wTDhJEZI3odBg3rdq8d8vW1s1pwwz+HIOy2AexKa
x6i/C5GkMoU1k6UBb6RJC+nMJJu42lfuD6xu/FaUsHyGMtcpq7Yhi56Vds+HXllb
9LwSxq/HLthDXliBLoTNFMkDjEhODpEZK9g/JKcSQSwLgOcihndDvfwJNTOtnb6Q
Wlvs6qQyzUPcq1XEfykNqlTNPiK9CjkZSG9cIqpcFMgTedKxlTGcakEl78iVWh3U
uiUyTWY0vu6GJpZhAPwEpv8CgF1e1TFSojqgohlvFj4szXC27MNoqpX7KdrkdGZi
3zufJqcGO6dMYgHLD7z2y0qqvVHTzcLOmoVOMSFnsEyEKlPITZsjRQ5zNIZMfJu0
86DgnAXS/cWodh0WOhR2/8tK0oelWgoCl+q+4YfoKJMXSmpMEDinZ7iCAnZu9AVW
cfYM68uMr4aRdGK68MRLwolDtVlhwrhMRLiIDpQ2Nx9nJz6I89mes8YswZwEDzcF
nCvNw9gR9DdrN/O7Vq4mxBb0lWAkiDRDxKHK/1efYSEJm9IahT/d2bmPi+sWayMX
2zIkPGaO+0KT9Dm7FISZm60OP3iksMQYVpv0ebgaLTVpycTf91ijOzoBr2UBUTwY
S+dN9iGMD2TRWOgYLrN/3v6BYZ8yY8IlmNk/07TJi9EvVOeITzUNtD0kYiYonLQf
cH9UUJElay7xvhp/syek1DUl/Ivu5kcRXCeQl3exgquegvJeD30jE5FAQPlLArQJ
DbQi77ZRgeRDS2LxKt9OX6LGzRR2rj5IfY3SIx6033/cJsUK3KnJ9NnfxVMbDPJ1
dEtMSgSCXKTyQXaK/75TWMBv/mzUEZVz42zYdIU+2Q/JsSHznYxDSKk0yZV120h8
lCEs3kB9MIlzGVSX0PO3QywprUo4nWflzLdJfYSgmzZuz0OMmNpYWOPmxGn5kDXf
ZTHw85SOhUc7IJLeO1mb+TNXLoQOWICwY4EYcAcSXn/NK/zVEUJh7OZXbPr9hzVn
cFc3lJFYG/weBJX5kCssPpuvUh8w9p8RjmcSD0ybe2U2jIfUI08y62z9zz8uw/4e
/x1jHMt3t+SR67fu9p/yGg==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
kQLY5GaDlX8ajf+WJo5J+MtpZKiZDU11H6C+GwcPcQ/kmqfjuXBsb4IfMq8aHGXS
Oh+wouWmC5yq4llHQ4ppbDPMLiVYF+2jMSWGn13sgja+iOtimNqnQd7/RuOlgIKY
IKpQJKmCzK3NdwQ4YQftV9N0trRT4g5zSSGUu/sJxTj2nBpG/f45PWKjif4fNdOv
Qlk1tv/OxnMuZ2lNPJlIyGcOtm3j7URoniPYQKICQQjBhktE7Qr0ghv82c0o20f/
qhGjjaLh0KDILqWamy6hV/hME9RyqAvwVBGx2rkNl6QGZhbLgmm4hurL7UZ6TA/e
XGrwUr3xjX5/6c+g22sPGQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9456 )
`pragma protect data_block
rct/jQhF2eQi+3Oi6Clh5LS8ZRGMdgnNiDI9Z2ad6hy9TbIHnHXaGeBaSncA95S2
X+JH+lcj/q/bFgNxTOj/DvbH31HkI8VUG+4S2Q+btU8sgufEGQ0BARaeuo5RjLS7
sg2GQxKei9InhoYoflijHQWMoo0AFcWN8yqbTFjm17Zt9EzhCAO4OclMeAd1Togz
W5r1oJsyRMk4Ala8NnZL4SJ4c0OPf/DaFg3xa0cNfhMWYVTAZrn+NLwIv0YwOv1f
LRHqJF95tUZVqQy9+9MWqz1KME400RskyEHz2bprPqsFptarAcq2eMnxopXAebur
YD6OMRz7sxVKshClJo6iKzVxejPH6yrAOJ8c6OG762aYPTknKi9uLWsOkWVoBpGz
7okuvz1mjrvbAVmFJuoHieDjRVWe9Jxr3E1/d+dK981lT/GrihFQ3o7zFm2wyF+6
7xrz/v4dV2HuRzO6yhonEUQmU1ITeQ4znE3XneJTWgHRJjkw8YwUdqHQIWb0d6M8
ERnG0n0j9il9rbV3keRBZbSl1+H+pahmot+Pq+whtdNR6kEbskuLyPHTUHGbUjas
HSXTK7wupM6Fc1KN5E0SM3wYg2+HhIyEHKhRnpbnk0WvBo4afM2yIqsb26AJ3bKy
WYpRLmP3F6lzeGtxzBJ2T+G8M8pM+8YArcMG2Hy125sa8ZpqNSzvuUmjAsMCAWUf
3ZxKVYIltdJkHBhyv8T4R5N+AhDNUvPHBGoY35BjW/TpSi/9DGBAIQKknnfqJNKA
KyeCmLpvxNBV6cifyiKPEG276wkqm7iXo/y6ep5WEVvEwk1CwHm4lZDabnVOKB5O
3AkgofjvtQzowReSZg1Mm3YYOkm8r7SE6LYa5/hUSNH+nJtYpT5574iB9iyHkNaN
rK6obkTMvOD3mXtBxEYxO3XK5NaRYTpHeCP3k+lfDKQfNrUyCtUkZdG0Wra069Lj
mRVDPsfd84vCPXvDYmTCybQ1nfbJZY/4xfKtux70RXxeMrdGksC5xByaU5A7fv9a
6TXSGBd3+SemQ7obl0l9gETsiveXnWsvCa1G1vhms6cv2zwmyCEeFN3lO8z8emIL
ELnaZqbdPn0TL6/Ho1yT575XAzey+N4q8F5l3EWMtgR3e5XqBoieuLfkoNqxzoFP
ENGv3iAPxXPPg6AuSkpXAjhUPHm/DpHdmb1ia3S6JgO6Wt+UBPYs/e+eQj2HDeLC
Ms3dXx9SrH9geJRkYK6k2TiGcwCjdxBn5M/kUpZ/Oj4t24F76WqYC4x77igmUTXW
gkjxdDgJo/ucFpwOY82em37WA3n/TiVLuFJEft+hsEA5CYcRhqD+M0mk310hgKyd
74pvUvH/7tFaH2QM25cPOFQ/ojMG7rhiX+YmSqR/z1rJ77wOOogM20xXMtuuXqUI
fOSlnj/TFGwidyVLi+Q5WvbmnO7MrBPtlLkuaNydLhJfbpVgoL/uoGJDVXQCJSQh
TxrLIYuz4Nuh7Hzi1orzwYXwWbEpYZ5XEQzz7Riz11+fg82xyTegzfCRgll0c3Z0
Jnj3XBY5Htp9j2yb0dRtkggxCSVEtUZ0gXijpJE60pyElnTFTBogLfs8h8pVflcU
O79Ey9QlDpVQ+rRgq0lFTcdCmNPXTqFxE4I2UlxjmPekdTcVftro1XiQ14YlXQFn
OXaVApknlio8t7G/A3QCA0NAOqbCJuT0F2/YJzwVhyRTQLt9f3RFH3gWaHlccauE
uLFIvCrWLLPi4w8XcuMQEeifvc68sqJoQmp5Ojw9GXquflVU8GNJC9FVsLyQPseA
sqCkRbhpB0q+LMkO5VoDK/YGULf8XnNJKe40dHkPctF8Zm09x49mfCWCzMijLcT6
/mwWbPi/c5316paHBSL4Ww7lQWmIY6fOMm0CMw9ZrXFtkW9YB/0LPt5H1xk1mKXg
46lOVkmt62l/RrMOibVDoU2XIy2MDEh0XwSUc8j7i6A8WGpPmdTfOdDlu2jUEUg2
n+w0ITg/AspcndDOPQeJHJXR+kwpy06j+RCw1yqLl/mDNXpBmYgg/k+lIGgrWGBw
H6iaUbO9mr1xGbkIi3Jex8bpI+hsbYqlQn8KVjYtUuAKOydjp/VU3WOrwcSzpoUp
TYTLZNwcMzQz17fALnFRKLqitwr1Bxc3uNNLXGi/tRx6y7GVvIqLOE+965iFlkWt
IYnlekGWpH+faj2neNoT1TWYiOmtPasKwdWLZgUhd/2wqDCtaHdwylahvhZKLM/0
1lBaILs/EoXokIF3GYgMymQrPUy2Et3ouCPs1B4EskLesBxHDHE7myH88RvfTMCu
wUparSACI8yvoRnenqA3p2SGHE3SKNWA7JiGYF8VLX/NJJrdU/7sjlinBm85KQCi
5kHZH0oXUASZAVUEjvoG0MnfTk/GLlL6RpvZystByJ2tftYL4ToQ1iVw6Gk0Mk25
HFoQOzkVeumrX/mFBk+G7PNrctKtkJYlTfCS46JABUQK1zjpLdaOdhVMOtD18pWa
4oTDHKiAV+TpWN7DZOJh78wtLmxOjqen0RzM9I2+SWTRe5QswX0SFEU4qA3nH91p
bjoYwF+YAFVWqiX5+CBU5+Kqgx8pnOZ0A42jJXg254mIjaRjMdgh+9jSMmICfDPC
NZsQx/nWzkLEKiI9WgXqfTVMRrxHoeMzQumHWWSlAe0zA3nPgbk5zdc6cM1VasP8
P1itVZ9QFBEp3UAkR9dKZuRtlPDu7eZ8fu3++sU8JMnqEAsPOcyb08wQtqV7emwG
dnksFA8gej0l5uhxix2jurgbK2TG0vVke2OdeNOLHFQxQkxXJ+57IPKuFhJ/ZI1N
V0Q7E8ulZbbG3Uw/0Ir35B09bkou6Yt/4ihxb2j8OD/TTezjVn/PcxS60WGwjPgr
X/3Y/hN5KQInqFGoQ5W6BccqolEWNIsvu71En7Bzq6MAfNu8Se9f5O1OafSyFswe
YL75XKmBbG68IqYSsQr1gnl2wjcCTcXV3BAIoMMzrOX7uKxjapIZwCEc1IrlQY0o
uOBVM+ha1uHhVOXfv8ZZNVn3ON/xWs8KgVNUzw123jq2PQ8NBn1H8IfnzS7p/i/9
vt0Ow4p3RjCIr3O2jdk52ujBxrhfEj7qBzxU0aQ6S4WDckMOjbxA9eTXoPEcXRQU
ywGKvlcJOb2Bnuh3ul7l+/iZ8jbYXd/+wM75Fscn9HEPDkZROfh9fuH+dbo9NgL2
8GHGsz6KPmaJsevcVn07kO8LO7wjl6wp2HSWyjpLuCOqqmHGmW/FAl0QClwKF8dt
0WdCV6Rms28ZqknMTPvuCky0vqQoEfPlkt1F4YfrYtO0HJIlaFGiuHe5thReBJbf
s/Jn++DJ6EpF5kPq+ScV8dmaPrG+mD/OrsZSzVNIJvN8fwJ4RfQBK3l+yQnMZqrg
RDAblaDvhYebAKO4KDt0bZeZR3yItf6+NjlcDaAJa7ozOa9syFv/u9Bz3tQVqY6X
whIA0rAzQIbCqfn0uKJlYnKtkiqS3TkH4d/o2Qaz+VFDFh0VCH9WjZ6sGc6mjHuH
2CgsjWYzxaUEeXm/uttkT1vc4qUtM4hG4dcpCYyQAlQweW37iGiIhMmD699S9T8l
8p+MG2NUUhY1Bbfxi6bz9+QWQDPE47H9rEs3mqN7pxQJCxQG0PcNsEqWPZ9ZVBW0
5YUVu4nc1jze/TKxnf+VPa8uvtN4M0FXmFNUvbnV+EGXhu11Mh6PfCVLIRL4E1PR
O4SvBKsjUd7x5WL2TOy2ewrnmZF7eJ/F64plcG3Ss04sZ8fPgw7fu21PJ2XuuEvp
qiO31DjgwsYG2T2WS6emnfX8usmOrO2xtOg/R2iyUZVXiIRcKjXx89v6oA7u+kQN
K3LN8Xsl0YVEoUiEocUHxKdYuQOKQmHkY5PDXQJJCZozfXtFqXlnB5QAuUXzdZWB
qU2G/rN2oz4WV9USMWdmp1jYiF3/Qj4fGCNVqem4m4kJ63J2EWkoqZ1+zK7dY3tp
ONV8YbBqAlRuox/E+YrQNVcWgAE0KxLiG2R+kb/CmDn/RUvUEPjHI6OJO3mzkzHZ
qGCkMoQfmhyW+IfzMGaUIjL6iw8aQJrn+SDexzAJJ+lwKHfEuK8xXlP0EC52ArD6
arpbmRpVAhOu+AHTbFS2H3xbtZcodKPB/OMNYL2Z6a7bi+0KHFS+R0wCqfD/OOP5
sCwbRKJnGlXjPVOxJDloT+wvwppA+qbBbtYPQqbmRJmp4yliadgfPXpwS9y50i3V
z1rmk+Ih05lq/6LlUhbsd2rAt0GQhaTm6EecZxWw3+pwj9V4dmqhPar1+HVB8om4
PxMRG+/BOvtwbJTo0rhWk0oEFm1Opu1PvChHmL65d73INlsQCG76v3vuLhUqy+r2
fRTClSjWNy0JhKAXDYSvok1DMb5fazt98Ok8RrxMMV6mcIoUQSpwdhCXSx8hj2EL
cwFZ7VLCCDzKalspXe8c3WmsyFlr6mN0x/BxNrIJ2DcpVRuQky90VSERWH7RkCTs
0V10+1+Lnx/fL3dbqkD3irGYgBSSnfCNz8TQGXOQNuX9hBVtaxgHfpzoi5eRFwyc
oDVjftTlUiRqmycICTvAQhlp5M+ZwYohnpD4hU5eNGRIHACVQDivDJo8bGzgfR9Z
Fjlym2m3WnxoSlD8QR1A/KDnkClVYO3cCvYeG/qfH7qYNF+NBvyrQswsWWIa3tM9
Z8+0MBCm8EY/Q7+rCSQBNYVO+Qca9QcRRryrlJrsVBwRqPYe78taAAAzscC/8YWl
ceZJVeR/RD6oWW4PRXbJyoz6yNSqUVu4PFuDxKuRXXqxWnyVIu5lIuwpf2zaTMwC
63XUFg+X18Armi4uiq6HJRwIOCvNbxfgnRGxNg+QsZkHsYlFmDHica2wIDiF03WZ
uqBYTj5k/5lsSeAAx2UTCffIQ+0cOBxtWcLaX0AEQBpfvhmhGoJ2uJw+Onniju+J
q0k9lNf3CjnaLEC2PLSOVu19hJquSPd0yfPjAa/j+dt3kuuGwWWyLyxVqMQjk36W
9DeJx9oO4h5GKwEQsU0jcqltUUDEJo5f5T686sB7DTfdeHe1YIdWaQkqEwv0H0Vd
n65MZ/o8zrOkJgCsiBIu3qwJ6ipKdX1nuz4r80Da04NhcSvLKmk/QvWCYAOAFxNI
/MHavyM8VXBlYQG7PwkDbl6zWjKM0ThUu7X+zZ1T/TmZTxYGFWHN3hOGuw2cSvHu
2HPwtcWq/ZdOMY9BI+7OobI4L0IijuvdTu4EY5bSweLKQtp9cFFdaqTIZaprMbMc
t+iUUbb075eK3Bnd4woemB/ahGaazMRGnzPoLQ8qTJj3ZioopHPgzxAUj8r0uneR
7cYbSHDpLVmfz1srRYWK082iBlfA47kK2yxNM6S5Em/gkETUkWK+cF051noGJgO/
+ducLsuMNths3NT6SiBC32ob08EYS2+FmA0pLwL+YqJzeLZGlyPmNunOVcuV9lD/
TGDQEN6MDnuGG6UvYFtQ7ym280zO3j1gqbR6QUIvRKB/mOjF0jLq+NiCySTSneVr
vgTN89oUr2trOv/pbMCtX6DioFL46RdGborWIiPLg/fa4/6YlnMX93WPP5eV/n9C
mSs8Jz/PTaOkmyT/+Gf1U68NbzpAGrHWXBy7x8oGo3e1Kt7xTVCIWqQBGIPmzcoz
vtyzcZay21UqlpWjDFOKFVn+CuMWogzfo30o2rbbjufUE8X14RI1x85eK4d4F+Ex
oR3tsL4HrgOyKvqTDHrg6wuA+zpy4+tnoOcWP//kCVyHJ4sHV64FlxHV4rm8OjZ6
grdJdHeiZKU4zsvG4I4gRJqbgSGIg8DKheCe7LIWyJjwcjWJ0j0h86jOcdZYTCns
rFZhBkiY6gMgqG5GmA59DkrRXQKdaPSGnrvmJ9X2PDUdXWCw7BnFYdxzXEsqRqfW
FTkCKRxYmUIGq3d53F8zK6zErkiAGnotvtVjBrYy5PFVwBIC07V28SEUr3Mg0YmQ
0awUahAGHGbB+KBsLrJCErKW4MuwZBoxF+VFB1NoFoHcMEEsmW7QDfpRjfgGBXmN
uhvwh7GBJw2WGZuaLdONvmGL+mT30tEV+KCYuPDUOMip1g4Ko6xCVkbM16ofVQRq
HS5yfs/38H35J3znySOLrOKvNxd4YKYu4nM/J8WU2bcLzGtghCgHZAmGIop8OvWV
x8M7AVXd6EXP7QA5S2Jpv6oK/2JD7f0bQHN7EtJTQpP/0eJyBuP7LYiItkvoZH9Z
PiTro8zcS/OPUYzorGoyQbAMrp0UzMWxJudy9eIMESeh3iApICZwiubA3siw8Bbu
MdU8isFURLHRDUPU1qewYElmZyy+AAYXNSvY+Q/jrc18nf8KksrLjZgG1MYNkXI7
s7pV35OG+OhdU061RQYRf7Yt7O8FCyfIiBzzuGPW4F/MSvoXS24YDqrPdYBD/HU3
MpkJ7yTEN4WJxKc84Zwa+d48vq8Yuc3zltAyathXJVAcffkUBJZsGL5LfSiSk7RT
1pPXe4tcJBdt5DKFS4+bV4Ap/hVRzenF9yCPkFSOn7llfo396jHPG6BHJm3Wx+et
C/ZLuP43D/hLbY98fmK3zuD+RVP/jYzDH0e3mJapDPIrWgLIeyYXYId20B7LWzB9
HkXOWiH0DBl/6YtKsdggxeY/XJnUYWaFibsz/iRO+QsKmii4Isc5yRbjr0Rbwh+E
uPCGXAnyAbANIQIA2vHob5cEaP212L3Zl/7m7SX2J4r6pAOGcLcaYTwEBHlvqway
w8s1jHZzAp/sHbVVPngyIYk1MqmNZbhptNghd/OHKFxXq7UU3SbJ7VYVTJ/DWN74
poJmqkaMynh6Ur2x7PdxoXpt4fDvUxkuveCLoAbViQNIC9D/RbDNzTvLyx+2+6iy
qI+hKk8wSP2jX9BLJ2WK/zeN6Rdqt+44GIXkLi4oRVD6T+YlCGMcQSiukqTNZ+xh
zuddplMU+K1C4W+nY6crp3fa3WwB5tC9b9GmeFJipEcd2lq3njN2LsYQgxXKdPm6
MsCs4jPcUmHSWRCLOKn5ECRvbErbOtCSLC0P5jhje9+wZkl+lZf4XBqRcDWlxvS9
tAWXZDSIwk5zKf4QGma5opn4NwDW3DSR9a7W87JrZ11EEp/EvMsdy9nCqxxXURgY
TLA1ddDA94Vj3ahXt9rawOvmchDTZq2OHS53sMNrEj3D+fP3tMmUZxXFgZ1sQBVy
knlYZQzIHQYK3vwhAGCqXOiKOLc3x2zdsZJ0/MPWvUh6SoHqbhBhMfAp9cbs1FBm
jZWKWpRKqb6k8fol4r4kJ8M5i5IN+C1vFvVTCaKW7y/TXVEbX8i06FgZ6xgGjesg
EYk7AkUfRjdRMh2IKG98cOl4gyf2H5IhnVDVVAHqhon/Ep/FrfbtpQc2eNhd3K6C
DCkOjzbWmRYoLxoxC+HquBafbMfI5lyqCKiVnIkKpVbOnzVWs5GzmpRXCqI04rMa
k8MrfcvTSE3B0H+8JDkong6fyicR2SOpPJCMJecqUh6VD11o3gRv/dewmt3gkMlI
gKfPW/CaYy1f3pUIKhxgYEVgjSJWyf5aEOYjBbR2Gw8k4zloybJvbXh1bTM8lPWs
k2cEKCT+RXTl+4pUcA1KkMyDwp+0Tcj1cQvL4gqCxGzmr0GMc4NAj01Iw5I2Kyh9
cXIe5YamScoSn882aZSrbKuFGqmYHOYvDA+hW9zebwVfZTYbapb2CXSfmKca0WgB
LiYVbBawKQfWEl5VUfMygYEJOfByj9kGwOxfwOt9rRS0538TkQoRdEgf0U7YBD0U
IOh74QiyYCYsu+Jhua7fZutYTq3BqwY+RmOCetMUQrV9JivjMfw5Y3SDLDLcpjx1
e5aasLnyvia+d5OrvX7mbmwaBO1r6v+rDiA7y6jTaFSsYcw4JmahPvHzom6Ar2Ys
6FTL1UxqE2aS66sPdgE8HENNJ4VyPUO6x7cUq1uF4tT/EOXm4q/7cpn9oPqvQYQP
0TwKVT1aI1xT01HymwqIeL4xCVBdVkBvS4+0qSqbV92yTgCTct7abe9F67iuyINp
8iiQtZ9hNJ/VKjkaI41NY/peh5+rC/QmbRT2YRbp54Fa42vN0lFz5bjeysUhbL/d
f3OWUmaaIVKu0qJaPgEHYoHu8n3P/ygjcnZqEj4VEnf21uLhOuQ7xJTZk62FG3bK
hGAieFMno4M3SDbMcLrYAFBJ0t+FruEs9G6NnRRI0mn9kxH57HIOsQTd3/itCigL
sm5VTuXezhKEpLfmyxXvTb9kXKvWqLtG4iNmLBUJMCmqqFfHXze3/sq/cVuZHMNj
YpCUSmfDUdgIAGqNTaQPNGosDFqmdevAv29Xn+bUZktqAUBtJqHBAJKFhK4Alv2B
uJgjkknZ0LbfyYCSVyures19jwmP7yQWby9p6S/WxIKcYHm4OoXvbRxXY78CL5++
g9uQVVrbZlECSV77BdhUtfCHmGkwsnZqU/EtAiBh2eGRSJoUidDYeaIKllYnEjxX
TnK4AfUcU0b8H5xvIVqdcg4Ntk/S3G93oFJ6MEXRPzPM8/zxAtEu6pKZaa2q8Qr2
P2bdJwfk3lPy6ytU7AI+E5toNZ07D21kG0LHTxNVdPj6PGZuDNOmpGasLlLxp2ow
1WLrRSVN++erOZm5xMt0bxZ0IXYHpfQlSe9NYrB3MzodJbdLlcicndL8KcbvLb7G
SBuLO7Mgsy16Knr7vUzXKgFE5eA0gVl0r4dHYJUbfpJhTVvc4MZdqMKhPaqzmiNI
BxO7UhSSa4Talps8f5zMKkEu+J+Jxmc4MQECbQ2NP0bLRGdRWcQ7AmtLjzSzHTBR
PxRi3mJWHpymsYV0O8alp4ud8N23nFRSuS6+jM35XF65O9dXiDsT1qGbEL8KPIpP
+qoS0j37LW04SjHhQ7DThAMHehQquTKZXXlZDr5KROtgGsdmNMUPynbuBhwldhmr
Cr9vvClXW1Y/TafJ5OzMkrWI3oZPydpiu6S5qGiUa0kEcK/5FGdQht6OVD47+ZzQ
t8B6dFsGTYE+t/Qe54KPRLdouTyvt7ieiFHnvdSfJSVPZRdfMRWSijD7O7XgL8bV
ha4xIaM8ytxJAxLWMbvliZ5RXevpgBi8k3mhPZKcZI4bc18WzEJODpZ62UdGkXJH
JnPs2+WzG6ZfzPQh+9KD4YZb462PjA6721vZj/W+K1e/f31t2zo5RgusP4CSr4AF
JjOTWaAYka1wX8RJ0+AN27AF+i34hflnxDb51eIqqYybfiwRCmHa2fOAPgiMZ3dY
0pSrdBLo7CKan0oibQ7NCXiPmVEzGTt3+ELDqguetU8Tzovmm0W6ysUnFTbDKenM
FBoG1mKKup8Rkfga5+yHHhSdz9EsTzAa74SYwu4OJSjBisIUgDTlMY/hw33GuLEv
glG45RbJk9B7WxjUxxLxfZdISYqkDaliX0K7rD8xcxUk+a+adoGJmyobHjcIwSCA
QBruOBoDfaehX+m0Pk1J9JzGA66D7nlfOyUgGrDgC68nMwG6LIKVpA8oGwiQDfR1
M50eIA7XQ9+kfiwJ302DJ5VQ0G76pWQKLIoyfcpBROu+pKCxVnfYmeje3NOGzleV
UaYbw22Xlu7OeDIqMbSaW1NShecR3hHlP6vlGfwOIfkWXvg2vup+j/v9ukyLqOdz
3LpoBsujbd6C7E/KhaYlV21nt6e5OkQ8yyft54QJbKRN85eJaS4tesYgdZH35TTw
0P6UhsIi3qbGvddZ5wLNjmvMME6T35Oqgck6kh7NQFTrVldMBj22/A6Qi5Jrk350
2jzMTN5JFu+H7Wams0vvha7P6kytKo0HQL3cR1/KvvAuhVhTXDzmpT8NEPlf32Y2
23pTdJxRdGwpLfMYp5Zyp6jusVd8nNmNNfJX06wTZ8iFa2NcBfNGDqfh9eT8Yk8i
kkZAujZYcmJrP9FNXEsFy67RkyYcyPYD6NISzd/5hpAm+G852YLcmzoe4lsRWcJJ
VdKB8ailHW51XhEZOMcxvfnZkDbMNMY/MdpNp8/+pgqpxxskega2b546juxr3xvK
F18InGxFGm3ewhAeji7K8DkHlXewO/GzWgov47fLEPvfV9wXbF2AtbBl/EOlTJE2
ppCG5ML4MxUhjyMs47xYmkmQvRAadOTA0CZKwkGT9F8QtLdvIOLmEJ3iTOZyZVjF
SqOrZQEXAe5e3Ep38KrlQfMfCvJ7mz0DdgTZ+BXM4vcpFQix4gMEIYYcJs+nv7jW
zv2Jkt2s4A3CbG10MWSnWsK6U3qmEHlytqjviIx+E6OibdhsO4qDx+nuPQoEEWiJ
F4rFttV1KyP+zGj04g34ANrUv0UdNunQKDfd2zQOHp1Mq+WGY0SCMZbr1r1OO8yO
hmTa0Co7TyKMtnghgv5Ere7iedkGqmM7U3ts31t7VmWAKKslYWnP4BmFYZfUwdvA
uoga4IeZBqB2awAiT3pADxgQIjVgJezLQxrk17rRhZU4SApbVebXpOWAHMs7kcCu
cWaQ9RaiD72mxpt678Sg+5xVg7C7hCA8ex+t3sIZbO9Wvj4C3S++KwJHIUNC19Wp
u+vaMx+43IIo7yU2KqiO5uc/PBO4FyXfG3r8cZHAhHcnt3EL6KEvIcJg1vvBlfR7
wL/H0cKPUpHTejad0EyfnBEGp4F0lyJY0KIx4PjRU1GbTc4z23b1KCmykZnOtkXC
u9ytwNXvu7QVmX3IU/uaB4i6Gv0DuS1o6vYtHc/Qq2IJ0RlHMxbGdQoPFMp6AA6W
eNnjcpQRTb2kRIOBsYLqnkKhlZxF6oM4ep7BfahSrr2lNWpqgzaCuK99tpLbfQ1O
TgRVau4P2msDIKL1WUOeP/J6broVYbhjf5Z6Oh+sUF1t1uG3XkeW3yOhFLtfhHMW
woZwqcDyJ81UkC0EgaGY+fn9nUa1AlLNsjFM4gNXYk35AAEW2oEBpGe6RH0GSjPq
kIk+uoLiquZ1eAaupJMFyWJyQqSVVYoh5rO2FeZ/pd3ytmcmGcw9LL+Si1azssNz
0VCMIxEC0iPsCxskbHEMCz4eKMsNZxOKyiGipJYhc42LeDmkHAgeP8uZiSPOTBEK
3tKISx4YeB2sUnNUUicJoFlCZ1vNgResRMO65Qa7zdvo6Lo4nfBMLYl87ExA5eFv
UbM5i+SCNRUdb4lnxPdJ1Aq+OLYdRpC1fWDLW9Plr3nTLLe/RQHao3X1E0Qn+LJJ
zpIcUkti1LOiiRAPY6QZli+uB1sYhxO6EWSl6IpUlX/rYwh1Li33xhvU/AFzir6D
vFEDqL9jRRy5UJqMU/yDgmblH7YV6UStlji2cRaKBxZF66rfRcTo8gvP5TiMQaWN
UWfh5pqDtRhxtp3bclcvn3qS9UF/P12KAox6dw2qfWS8FkNM/pGafAXd4w5TfaWc
PDleUwBirHj8U34/pdD4PvlHvN29shmn2h7Vl7cte4RXM95Z+N2nACD4G9VQ6MTf
fuZ5kvTggjtaubuWx3e4dX2/c5SLnt0wa2RgRun5YH65+cxNbGdCs6yaFkl7AqlY
PEKpHroFeoBzaATbfBnZgK4w02peQOkhCJHrMUWKKkd34/Q1kFYSkuB3LkCjYkQX
aEFN5Ocy3Ja8LTKtWI3pS6K7/yQbVXdL+olivVyopYtz3WqOQpcUm2HVs9hGLceY
0YeR4N93jbsTAcWolQh1Pf29yDK6JXnFcsv7vsN73wYgzYcgG4Boa4Bi4H9mgj+q
DkwrZC9IB8DJRKuC5vLTz+dQ2wVfy1+UwMIot3Zdp6ulcCWcD7As9wz8xFHt0dD+
0s3ptCKcIy85Zpv+wopRr4ufeoo/vzoWbMYcQRtJ4w5Jjwswe7q3ElF+kb03RSkf
S7xvqlkRTQ5mXef2S6309ErhP0zbAgg+83xrt9t8CmS89w+6dfZNRD4tUuIIzaPI
PIHyMKElsiRtUC2y0up/uR10VVr1dHZwxPbbqavETsjL6HKXuhG62u2sDFJsaoYY
iag1LssWrjGD1zyb4K+XNFvoqpSqN4SUXz/C2drh3lvcFdOriLivBmVZ3XyGN/g6
ObJZ2lHtEAoUEOUeeEkWrGRVCd6VEq7+6xDZo08VqCG2JfjIHhvdemkUv9i99HIN
pZIVQz78X9+PvxgKEHfhobQndrb/ISOh5f0Ac+kSh/9BSlzarrQVJwYv9FBJGkpx
ZRXZxP4UzrCcDENx9EvQzm3k1rKI75YlfQicb7hd498JBqRKICTDN061R0+os3r+
X0m59gxpdsY6HWGlmCn0IBwe/zvdto02Z+ROtC73/pc1qIhAYC3hD4hI5yz5bEEM
bsfC1U+UfQ6NtV9kPo1wXB6r8DerXyJ/pM2Ez7nA4mTLGPFJDi7gR3Qpt9WlFoYo
5erFmrQ2rm0kiXroNSfdcUELz9/oNjIUIqrLMWjPpXcNG7PFqQXjubPsvod+3lTt
0DoX5I805aajFQe++6Lzf27AaWFSEQ/4y7fo0unZiYYwHcvIaFEFat1n7f9VNteJ
cY0bK2ve8Z+omaE56Ta8blfgOVmt6CnFuHjEdi+eGID9KzrjUuIs2RyXfAzRQni8
EESm8SEkYq9vEysIhqfXixrkIRMa1LSsa9Aw2p6aFUAwwGpgJC9dH1RcoOJS10e7
8YXJRz0SmENn/TrIR6v0TZCIk2t8/ag9q5RxINWDP0KV2QVP//z6m1MLYBWyeI6k
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SVU9ts6/K9sY3P4VBK7CqpGcoWXPwcEXJqcvsvke+UntwUEDkKz7gZk0SfS1Rknj
5T2ekimpegUPnvAxX8NhHiK1/xceBbuvBkBdJABetCP/y8qa1iu6mdOYKRT+iEkB
5Nh/SZK0tpVAhg6jNBMolK9FKUKmWhXkE9NwB/mT+C+yCRc0cqEz4vOAnRqSHg5s
GBrb3/QhZBEZ795Mf9wL0nfXwpiZ7FBhmaOaF/NcARpmvW4bZ1MYdsKGDx6wAvmX
vllML+GvTCBn3MA96rDYoXLDuQ3vOhQQ2LTdUlKM3PuadnOaXRt68WU3zjEtWUC0
RKw5GNqEQWNbCNk/rX/0KQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2672 )
`pragma protect data_block
bdX58E4EMrwT2WvRn4b3FOHRYXy/aOskLGSkOrIljU0oVysdr+lZDAS0cax4HUWz
s8qS+c3YVOeFuUVDVlvPOPj8YShH/gB0qf4WkxGS7TKEUkDEzsQAJbemH4nSxva3
uYyXn3Wi3cqKgZ1pQ5+3vaBklL6MUAG/rVhMBIvm36fHyRTjqx4b7eOlFpXVdbiO
FO230x6805HKclwrAr88aGSUK9j5w6FknmBBCygFye2/rCDdb/dm+DPxDDEE1lLn
YyuR9thdTQd0X5Fcn+ZGjDRQnRVTotqfsCgFtyos7XJtLDZJXVReSf9ECUNScjWP
D2qXDWl2UlAIXpcNM4V/bSm2543BwdAoPNb6/C9ppyrBzXOntCfEYVGTOr3VRxHj
LiKUtMKkw2bx++onAlOMFU1hJylElLzBEuHUdnIatxdGpOuIhvGjzEqkHB4eHJql
OKbl1XERLqC0UKFwpTYu9VU2sVs3ghaYMDrpYN4CiWoziTGBaOYo0O8paS1tgawL
Eh1dkXP9nWsr6aDGdI3DlfRRStXeubKjerdaTm5BJ/IXmy65xhDS540IbUBeABvL
791lRGUWJqttQAW5RflYT923MMP6Guty+Zdjwk8mypUgawUffo6eQTBiS0p6wCwv
lmDK4livXs2OmGNKdFSjSot33KHhPG4wrbbgFojTkFL3ii9VU3nckdCYajMJL5gZ
NiUj/PP2tVibnuR/L29/5YiCoBZqy852hVPi+7aJtfdvBFjSvORlZ4pxfM/lbDcm
FPaXC8nIO0In7T9VnGmAn0foZChNuhwNp3QF3bOekTm1JN7Zosc/WsQND0dZ4+q7
undRdCGfozG6dp4QeEaQIpfOgqGPBf59OBkGoUtnFzFKG9Xmprm8btq1K2ynE8Wu
wjnvGosbIs3xipSc/Wkjzc8h9edI/fcHQZKscrvIwgW3GRSpQR1oDUm+MRtwTabq
CB84rGOyje7hlU4dSLxnIo5MomaC8dUtY5kBorMCV/xuMGLtPmckdohU4cMrpHHR
Rt/B5/PWxZK+CIb0NUR9AXkI8eV1bdWHQj/bfMmViGw+ja52ylnhAJpAXuMRh+YE
a5oMxB0OFoWEGA8G0/Ke1OV+8oFGPoYCpjVZVSF/+iFhlvSHCtJ9z4evogQ/xWWQ
uWEpvHdhnwRigdez+Hkby4YfjsOAja46i4OydpQL39XGl4l/RV8UohiBrSQK4c9y
eGaaDrjY9HO4E56okKKjyhKXV3eIQpipMOe5aGDqAnVAffJ/02fcBzmVtMy3JsFI
Gb0yS9GaudAhm1yWlqFlJu3uPsvgDesEyJQBml0HdFBK9bsr34taJxaH3d2h4k7n
X0K4Jd+cwg3iEwOOs6R/+M6UkGpxBeIapYwfE4ByBnbNW0ERgkwB4lBxZfz+d9ts
revgwnz3bgpbV6YKjd9InNyX3Gja/lca81pFSZSQEFvst5qynT1rFuKw5lhPCB6v
SMi43DwCkdRhYjxKRKs/4v+u/b2eaTVCsB+pbZcYCxk8PJs92ilsiCzopmfr+1f0
4zr9IZdNrOq/RYUEl+aVT2cYG2XRCI/34w+GSR+xXJ03UfYviGI8u6/tgKgGo5E+
gdz7H6ywXJpRIwW9hAEYoTTSrp2/JLYv13kerEOPVh2s64l2tNCUoTCbGZDWpmTs
yW3ScEIEwanFM8tCnDrrQJzU/wOnbwIq59wFjAgdwNZhCX8LrkuUfmq7NXs+IzoD
l3AZacFR+QW8hgV6XRUfYo6S31wbhWiEOv5WwWXnn4QFoSVnMVDNtQH4te4MEK8W
C9hsxoMSdqSqAJPkOUwZNZ96ru5EMpYgC0RZoDzyW7ot6W4xikyh1uehivPwl3Iv
2E/3ep9lctI2g+IwCiy6rxzGlhPaK40nf+++h+Dp6n094vc8jUTwZIC2JVADWvif
H39CmvjVMENVsA6SZ15cE2l8E7cXXOyfQ1N4qOu94dF177vEzGtilfT7AiMZm362
GKGNFjNLpALxMC6zdgkWUKOoU6WGNST2CpZuKBAdazWJjmJPM8KjmLMF8J/Ury/T
dd0XHlpuE97f5bIAH/lRVtB5xup9yhq4xHij8+WRWspb7C2WfqgoTJy9lgEIB8tp
889bQ/Xp6C4VZkOPfCLbxC0lTSV66UgYXhcsA/19iZozL5rCodceXzGreaT1usme
qY4paa4Vxis6fRPfRzP2BsUjEbomD8/+rXLXJoCmGf7JQmnuzrc9r6yyZeEIpFCj
/MZUauD3aRsKSfyfXVNZODrSLDSx1HszQYIhvGEHXZqqGrIAmqgPMoxjYmquBqiG
+ih9w98ghXsWIi7yOqw1ftjIov938+aAuWuqRFVLrBswJkF4FO0lwzvQouKpua8V
4UHT3AMZxAH0EgK7vRIDiA8ihmfnwfQXf/fndteIuyFfb/GkGd1BqsIQp96vuXFf
hH2PM+eFz4kDI6XDRhxRUIpeVx3GYQFWZ6ZKIFKHVNPdoCkawDxrMVL4pNkSX0mb
EuTY6ArqFaS0bNQ2JhzIAxwk4b646X7gQO54N2jtwNihrUo/JyX6kHcdccTffwNH
byHj6SARrklWz0ACiyHeLfG0EybCN4zdxPftZB39uIrbigv1CoT/EXKIGXR7iBwY
7ZQ9+IibuZ0enbXIz50CqB0hv9ULjU7se71w+VZ5tfUsvXRJqpthJ0tNIrvcu5mS
fbk50DomyDSscXf+CTccPBUruNBwFJd3943/fxEWsb+cZIiRyvdE6htrMXpGaX/Q
irN/GDMQZNYXngY6RuRZ/QBGDW+89ecICTTTKOKVJHrgyZNnT/C84G2UqVgyb1yt
9gG8mOZleYocJIiGpcCGGiFjI1Le0b/sHLxe6pAjb1W8+dkoUhJLo/ztAI3pf5L/
cozLXXkWSd1owkDBToSx7wLARw5pGcKYBZpXLx6ysxXrPTECrIskOqRiVvkFF8w4
ca+WnsbXksvA6YVeKPt611S2MS3X9DW5y9rcAeNUDaS4ELrlF4ssejFBrITEUStm
vC7YInoH7MZZb93o0LNP47RL0JiOyBBpUhyeGiXHTbU8IbtxFVwlswuh58JfCIFV
cGg+7jVtEDyurECK7ftvqP8s229J3tSjeRZW1LDvUI7UEZkN9PemRi8eT5GlTyNG
Che31yGu3EKIzVEJOV+Y7iqtYXnvpUzAjWwlEU1K+7l7c8le+NVsXPuwN8nk2PO0
x7mvfzzhvUOd9Yff3PIzru+EG7jjTgMRItZHhK2XaORp8Y7Dt2VVuEWLVLw3M2Qu
KiBdW2bkV+XarwdCXOoZUs3b+YZt4zp02IdPVFDQvg54oZHJqfMHHvDevdp+Zs6b
bj1d/bDSXw3gMy9rzrse0MJySWDSQx2UX6EHLw/P4r1UIaPApIHNqF5sLBD2X5r8
HSxyQ3fHGMDiRFuA8IRT/uyjmvMPF+9DPKrDBXo02FFwQUJs226bJ0hkd6l68r/F
yqoGV5bKaHFHoB0hP8ZcKgk2rJTQHZxEME6VVlS5URWORifZVKY1fpHtKBziS2Yh
+JRGULxMDE9ovMgD9DhYPDmeycD+VuO2G1eKferLEE0=
`pragma protect end_protected

//pragma protect end
