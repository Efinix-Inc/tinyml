///////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2024 github-efx
// 
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
///////////////////////////////////////////////////////////////////////////////////

`define DEBUG   
`timescale 1ns / 1ns
 
module master_coupler#(
    parameter                       CB_DW    = 128, 
    parameter                       M_AXI_DW = 128, 
    parameter                       DEPTH    = 3,
    parameter                       AXI_WR_FIFO_RAM_STYLE   = "block_ram"
    
)
(
input                           clk,
input                           rstn,
//Slave Local Bus Interface
//--Slave Local Bus Write/Read Address 
input                           s_lb_arw,
input                           s_lb_avalid,
output  wire                    s_lb_aready,
input           [31:0]          s_lb_aaddr,
input           [7:0]           s_lb_alen,
//--Slave Local Bus Write Data 
input                           s_lb_wvalid,
output  wire                    s_lb_wready,
input           [CB_DW-1:0]     s_lb_wdata,
input           [CB_DW/8-1:0]   s_lb_wstrb,
input                           s_lb_wlast,
//--Slave Local Bus Read Data
output  wire                    s_lb_rvalid,
input                           s_lb_rready,
output  wire    [CB_DW-1:0]     s_lb_rdata,
output  wire                    s_lb_rlast,
//Master AXI4 Bus Interface
//--Master AXI4 Write
output  wire                    m_axi_awvalid,
input                           m_axi_awready,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [7:0]           m_axi_awid,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
output  wire    [2:0]           m_axi_awprot,

output  wire                    m_axi_wvalid,
input                           m_axi_wready,
output  wire    [M_AXI_DW-1:0]  m_axi_wdata,
output  wire    [M_AXI_DW/8-1:0]m_axi_wstrb,
output  wire                    m_axi_wlast,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
input           [1:0]           m_axi_bresp,
//--Master AXI4 Read
output  wire                    m_axi_arvalid,
input                           m_axi_arready,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [7:0]           m_axi_arid,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
output  wire    [2:0]           m_axi_arprot,
input                           m_axi_rvalid,
output  wire                    m_axi_rready,
input           [M_AXI_DW-1:0]  m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp
);

//Parameter Define
parameter                       aw_State_idle = 3'd0;
parameter                       aw_State_aw   = 3'd1;
parameter                       aw_State_cmd  = 3'd2;
parameter                       aw_State_data = 3'd3;
parameter                       aw_State_done = 3'd4;

parameter                       ar_State_idle = 3'd0;
parameter                       ar_State_ar   = 3'd1;
parameter                       ar_State_cmd  = 3'd2;
parameter                       ar_State_data = 3'd3;
parameter                       ar_State_done = 3'd4;

localparam  S_LB_BURST_DATA_NUM_WTH  = $clog2((CB_DW/8)*256);
localparam  M_LB_FULL_BURST_DATA_NUM = (M_AXI_DW/8)*256;

localparam  S_LB_ADDR_OFFSET_WTH     = $clog2(CB_DW/8);
localparam  M_LB_ADDR_OFFSET_WTH     = $clog2(M_AXI_DW/8);

//Register Define
reg                             s_a_busy;
reg                             m_r_busy;

//Wire Define
wire                            u1_wen;
wire    [CB_DW-1:0]             u1_wdata;
wire    [CB_DW/8-1:0]           u1_wstrb;
wire                            u1_wlast;
wire                            u1_almfull;
wire                            u1_ren;
wire    [M_AXI_DW-1:0]          u1_rdata;
wire    [M_AXI_DW/8-1:0]        u1_rstrb;
wire                            u1_rlast;
wire                            u1_empty;

wire                            u2_wen;
wire    [M_AXI_DW-1:0]          u2_wdata;
wire                            u2_wlast;
wire                            u2_almfull;
wire                            u2_ren;

wire    [CB_DW-1:0]             u2_rdata;
wire                            u2_rlast;
wire                            u2_empty;

wire                            m_lb_arw;
wire                            m_lb_avalid;
wire                            m_lb_aready;
wire    [31:0]                  m_lb_aaddr;
wire    [7:0]                   m_lb_alen;
wire                            m_lb_wvalid;
wire                            m_lb_wready;
wire    [M_AXI_DW-1:0]          m_lb_wdata;
wire    [M_AXI_DW/8-1:0]        m_lb_wstrb;
wire                            m_lb_wlast;
wire                            m_lb_rvalid;
wire                            m_lb_rready;
wire    [M_AXI_DW-1:0]          m_lb_rdata;
wire                            m_lb_rlast;

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="ipecrypt"
`pragma protect encrypt_agent_info="http://ipencrypter.com Version: 20.0.8"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"

`pragma protect key_keyowner="Efinix Inc."
`pragma protect key_keyname="EFX_K01"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_block
YzB/f3oZpLyRTJpEiM7+zo2xESiZvYJFHQJ/XLQAFiC4+RcYCzx22Ut4hbzpYmbj
EmmgwNd0bD6aDarVq9nU10JEU4RGzZbe1YFkYhokVj9v5jIG8VJX0oco+rk5m2PY
FzbUqJUg+vWLSj5KcmtHKNt7wnch6jh3j2VikftAQLPtiKhIFBq4OayJn8O9c3g9
Vi71QbQ4Ai1/5nTJVMhGbtkxJ2ZnvIbkR9qdp2HrKHrUNOwoaCpIl8uDswlZilRD
m5vDdZ2z6+7b1VT3g0cQUGskO5DLCmnvhL6rJj6sHg97p5PmRebbVGheu+UgT8Ow
+uWdML9FpShZBtjacgMccQ==
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_block
a4BoAN0DLu4GnDONbRq3wah3cKyoI2hkjQ7dnxljaYU3i/PNlTXFLNyr6Rp9pSzJ
p+01ijxCchmRtQfU/CD1fAtMw99O5SDlWEPnAWzBtLYrx6/msVYKOOEAn1PbUvQP
3J0cFSYSI7wOXActl+EJWn+17+PmtcgaPW7FFvqqkn8=
`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=33472)
`pragma protect data_block
7zB6120vnEh6oYAZAMOHWiJVA4n60R4YJ12KrnNzri9SKm5ZgddhMH42dccNgRpe
dtgzkgznFaD7emTXYkqeVQKHGgtiLJIIt/weCwFJv7AsoesKG4pLnxdqsghtooym
X+YEA3ktVzKQQiakzyCZbNKQr0NImHI4IhuuH7gZOSdwlhXb5YdqbK5Xe3Ge9u4o
U1S5DCiPyUkQj0kJvmDR53aeRgEybT0xxKSHDs7Iw53WMrZRIfr2mgfnJTj8esdh
7VC/hxJH30fpo+FzzsvZS68kWIaxHZ/QZwCKcUJqz7yDSkVeLo50ljncsjXFWk4E
b+JQWXwQKvMGOEhrXyHnZk+jJx++mAomHsiUMavyLlF/gI7ZR7uOyO6iidlHy5YM
xALoliE/9tVxAwUT3BnYKR+bQz6HLp488FflM/2M95fEF+539vCiYTSyooTXJx5e
80q/dSwPHjY0b4TvMSL8S4wA6BInQIJp050Zw80I/z21owWnHjsKAHOlbuVy9U1a
R8D91hgZ13svpw5g1kzd+f8cllkTWhfUwpSwBS/krL/VhYNVfBDdl7mXyqKijkR2
eBFVcT8VN3Yfyq2dY0jv+V97OMRlX68UeOn6edXmngH9rM8EaFLYnUZIPb4yL6pc
QzvzUb3pK8cjGbVZMAP3rAl5JtxZXH3/t/RyYbRKkNWn4MUzx/ZaZcGyQx4Us+FA
0ABvJ5T8J0htYexyOaajEkRtrXep6LlYQI2ovDZH0Wz+o/L187Oia3XdZxsqLKoj
5r1K3Ju+qZNriu+MOb4BjjUmNz1ePE3VmdsPwxNfT1WXaACNvPG0X6CcAU5zMEBJ
zJeDF4En/BzfGCSHe2/yYcVVfc2gaJVe0c1No9Sel26JzPJCxAma3nF/5VqdATlU
scLS2CK9+NwKZiLPOxbaINPPLLks8e6bh7M5ZH/i589adIyIZIoBGyTLWJP4+cDa
Cre1FaHikLEYFYh6N/2sUqmo/R58p3iufOlDZ+ZsUzf9BXDAJEKizG0rmzNIfivA
aKaFH3e1biywpFTeBq3ynetiOEMqKKGga5RKJ9H2YxL5E5TCLQX1sLi1CTrQ2J8L
JjrO6maLhcRtgQtYETBboBXnS7IaN2Psg9mX+kzo3cq0qJlik/r+62W74BgOuivJ
/ZeEuX3sberuWHzXWbQSwCGWoHjYgd9Uee2nfAssQ9YsL60xxA7Jqdg1NqvjoVgY
Yt5rnOnbEKaHOPLGNukWBr6WTqvDLG3Gsuc0zQENyVa6wkZ81YtTPfxaOEgXrziH
n531lt7TRk34r8vYWs/Po4UP99Lklfv2RHA0nq2tgrZ2lxCi1zWmnsO0+EMmJ3oN
Bq4lNVqkLmJl+hJMMx9JVXGEbummiRJpfbLtYtH29NTr5XCff55XzZIEqGZV1A5A
Ax0/gg5QXwRAkfG4vPdrcxyK5NwLGynQWrhnrP7HrxxnSQ7pqrBMzg6cq1P/PGNQ
FJtAQyByM0sEaD81WwV53RPzGOBnN+dy27N8Qdsf/tfQU04Vlm93Y2ap7vYg4xgs
4xAFWNhj+YWCkq+wZuQ4lI3U7hWGSsCjRfG2sM5EOXToQzP/Qr/j7C6RHGJMYDUR
Aorzuhxe+gXfGmN5S37Dk5marAdQeH6oIq3HkMPFIygebUMfqjb3N5KsDBw+VmUW
l3xZWHs/Lr+ov3qmTz/n0O0E0fBrzQPIyNTiWVYZu3IPPAJN369afbS0JpkN0g4G
JiFRkEoFsfVG4ORtIJM4HncXL/JoBiXVrJiZLo64X9Z49jnGu9u8Fncmqtnd6By3
B8FI/y+YSfzFj+5yG/zTaPQ7CASEFHcJvdExuZ512ImGAvNAAFx6DeKv1HR/pkgy
t6eUygFMBBA278KbGrzN+UfC9fkT7jBiTj/eS5yt1KpX4WJbJXl2aUpWN0AJtRVY
Sc1pUP8g+NWaAfJudb9XfEzZ8qEHz/xj4Ju/LlWxSv7vdmZKVjWH81J2iNpoOvwc
40lih2OvvPnsnggymcJVC9jzug1Jyl/uSWoEJjHVEANs5jcysJabJEhq8S2NBRUR
k+APYTUSHg2GrnnA/oPbMqlsmT67N42hUC50HzreJ+Tg8gMNL7fQcs0JVJ/Q1PBn
uCZ+5+VAtE1B6Fq2QHcJM/yOdAKP8+0t+YTD7JnbVL3ZYDSX9w/6lDC4L6Vpzo8Z
TV2yHgoQhU4jI1NKZjVKHhRn/YKAvJcm4hEC6SIK6nPcOWq9uyfk1EuFquy97bVY
Fy8vZM8X0HtNXd+Rp7ahMT1mdBhYSQzYNWqZDa6jtGkukmPnBGdThhpb8ohr6Owi
q4AAIRg99mK2kPFGBbC/EiAQQwnAxojS4AYEeyAWlNRQe8FXZNaCOW1ADsMfTDHg
4MFRCf0PkTs0BPclVK8Ste1spdpFFUVO6xnfRLzQVSkMsPzx2fYkNjdMlCJreiRz
y3bC+j0FY72LYrevSLt7O47t6RLhhM4iTrBX5VPcLHHcywRVo8+1fpPcpvPqYqxC
ZS/7EWYxiZaqe2PONV0wTB23FmibrLgGPitJBdfC969ueMunzSc9JwvImQ4K5MAN
tle0SplQkg7Cm08pbtf2OAQsobs6nFLx3Js5tGCrf+g6yVWaszS4pgvxR2aTdX+u
FzPik6d57DH9NbrmyGR2S2ZWb/LBXzdXNQeaBybAphs5ahWEZ/HI4b4OjSpDG0ES
8MVT0rXcogaRgPMDWVKKXHx6rX4JSM/eBjk9Kz+BqS5mKuvvuMGN4hq3e9h+F7qf
Bqw/3Dnpic+xW+7kw9M543FEgUtJa5NWvEIyOYOxkrt474kUv07hKMb8/e3jWZ9R
fhStQMrscI3L8/gTcMQhD5oPTD8ZHb0ccKXEWnDgnZ16qSaqcdxavpP2IQDewni4
nfTQili2uO6HWMgqOV7Q1c3NhoNwyNv4lJ47tlD99QUht8SLLdWnhYoho5m8FDtN
yZC8xrwac0VLy34I2KqucFo0U33PEz1ZvMw8VUzEaY5bLvcEY9rEUc7eLEhTQ7c7
B8vRzgfur1h+RsneMKYFY0ihRAk9jENYymh83HynSHvU4tGcNfAdNKl+ghXYZkUm
5pYMcE5czlSfNagjqdATXdoP8fSMfFcsib1bZ/useCZTozgJ/XhxWWc1DOVCz1JY
eimtDp8MNMrITJwyN+XFjQJ7wiKGXbq0+TnHFz1ZkJkrJbunLb0MUsZJH5oPsTuJ
ZDEa06uRy8uvd04oZBeQdTg9NlC8vd/ABpkwwxMCN0Dz1bg0LcQZnKVjTDZVr20P
baZwPoymBN+b2AnDfsR7Q/mvld+FimOfSSm69g5ymhdAsAHtC3SbPLMODLtbfR+n
eljRGmMBZgWSape9FZGrcn5eERF9imAVp3V6uYi/CGhzjainN0dqDZxaOqa4w9QD
XPaTgImUJ1PhWrRyBfxWqm14mGJKFR53yVBdAEuL7TILer8FW4Od3125cN6EGEUD
IGEzALL82vue2erQnyhknodbbAl26GybDImNWqKlFi8pv/HDlMAAPqOEBk6xX1EG
jPMtPrvxVETxnXFMcLV113GUljW9qd9pxFEkDLVuW5nGQPWf/rZfqEKnkFGGRMvl
HiFpHACpSHI9FQt/TkGs0XFmRFySdp3HRmx9POu9uuR50RwyhuFBc0pgBYQnGIC+
FzGNKNjRaGwQxKBlkhWpsbIwrGotRUurjH+A6Boyla7IvZbebrq3we87byJ96Vu0
QFdRR8DlqcHsThSyE+golTnb1ovQ/aLyJrf7XTLjH2rjZiS+tbOzM7lbLrAzQeGi
vn/TSigJbfyIgYv0ukK8I9mgasZXdijsMxHxZFg1Z9/Tp8cd38ILe96bhwlRSHyp
GaqBnmlFbPK2v5dEnUGS384lNMmJ8O8Sme1IHdfRDtdfv+qSnIhgNKUV/g9NZq++
Kk5nuS7nEJZUAmOPKk0YOO3vX+XjsEhZaNNxGi1DkB8qI152hEei9vjYMkeHNQda
ZJAjin09ZfRa4UzJrBSmZOADcHcy0riCfE97oEP8p0biZJA7Qr++j39wwQAm7UPh
/mL3zhR9ELV4JZAU6ZlKUbQABBNZBNVu4RQX+Yd/2A5u/1JNx9yuiRSLLrRHWOla
k0n3XhyepRnL9KXaQVs908/mXoZhIdf9M898iIi0vxfkd4su9JO1/e3rede3tVi2
gW4zf+FVcQ/gNZnDRgadAMYXaiBpuX4h1gaOSPFvriom9ATWnwxSEwMDp55xQQE0
FalaT/vcuD3wTbgdiBVUGhJRkThWQR3rVyarhDc0yAxIUIblp4rC/NZJG+dSFQS1
UngSiCSuWws2agtpUXuN1Tt6vTAxLp3ow36NALuH7tyiFBo/+QIlZICquT8E5nqd
/uM/j6P4ASUnsUkEeG2HaXowLjNCua74kgg4HCKFqcYNH4iJ5zkIZJPOXT/CVGqK
DnMpwFm9LyctFithcV26ehgnv/+lyyrB7UE94YLr1y0TN5+VIrPp9V08lcmIsmLa
HBW/68dAhdtYVZuWtGYpMLr+4/HyZbkm4H5EqpUpIR4a0R3TZI6vt88a7EOERLQ6
RPaM6YLOgOeGR25M7fEX43Hz2or49R8DCXvOlHwNdHcK0xN70dgunLAAgxsW9GmP
2ctLjrR019IXwyeXck5RxkNi5X+iBsYXDgVLlsoDwUSZunQXh5ruUiP7K9u7cMA+
hfWTfjRcw2pyFV+nEID6PdNdpgAAk2uXL0jalhegmxpxNZ2sA+yQ2ZmaQ+86os/K
+2Cul8JzlhCtXhfvUWIOL+b2zsnzkTCqEj2229BWF/+Nsd/NbD3kY41a20sQJoXV
OP1bZPJs4tarFQF2uzfVoEcHHNrGTs1iyjyvWvxY2Mru74K00D57q0ClRQiIIt20
mzuNKbpM+BLV2ruaLdnst2Tdp69n6xN59Ym7BvGFeI0wA2Fjm/cOIDPYYexUU8aX
dNf0a8gIapjicxiB5j1YqlSXTP27sF94Qhx+aKhFabYKcjZ/WIQJPOqeJvOm7cut
RCGMHO4PIUmWL40nG+N7cx5kk0fwdOLFuKIGGwAMuRnTMnbE1+bOLUjPY9vUPAaG
AZUXr1WIPPbLVzEuoD8HxgMnAD6/H4mKIDX+dUmwZLXJ8mPJDwpHSefSZUEObbV7
C8Uwrs4LJen+4DSXZRSVD8XJ+RzLLUZSGOkCRL0wjIehF9RxKpcsgcYCVvlu35Uv
XwofAPqIx/5fXC7NVSixjFSfjDXLixXgBPfHzPGxs7NL7CJNuPgmeBgf8cjJD6Bh
XrnHpZLwLllRYkR+imY6vANP5BFV/9eQunwf+jyGmfC59svsFIu81AeIAzJjM7r+
WjGSsKsY8l2Egjp0u4E3Ax9i1Fg7WRmNmzs2jG4EIs5foe9jl0AjQOk+f3a9m9FW
Xk5n4InkMAtbAJ9Whx46GyZY5K8+InO8sdykfbpyu05c/uo3EIK8zcufkhomBIu5
ngEWBnEB3oMxRaQeFAUm9WlOFDdd884k9PTuuyvWD25JYNHf9GL5hhzlOPeScP0w
MWJ27p9a92gYq7GRbu9YxsCF1pgC6GzmF4TX484LMgX2ylsMF5zms2phgH1puU7w
ZlbUN7uZ+o9wAvP5G3AgUQmE5+7+1wiX8lhBt5ITJht896ky0ZIOn1KmU9SKwNCw
hWYmzCubtiL4KhjbbYr/AN6zBUEWMH4aNx7q3i5AmyZHBANvSbu0+E4z5dyx64Y+
Qx4sMFg1ueCPImJeRA32DwkC9a3xMbBLB7TtUT0o+iDfepnDcH331UwoCudQWWth
Rm7gFCgh1/w1R9JbVNuKkR1XifpJgOVzuvH292q1bStm9/IO3lD7MlLSI6OKJmqY
o/JoVFGXZ4TKQHJWudlIHjANU3+5hjGRtfb0rjN5jVXqLiTRiTl8fdGjxaH00so0
ufXkbDYXyvELHycAmRUft8Owsd/VHdl3pL5JnmT4LHG1QDPYgqkfmEKfhiAJmfNv
hnbYZj1eD7OPQywUCZtaedk0GsLE87p6JGXZqnZh4x7fZ1GZJ/F2c7gQrOVLxgn8
2HAm1FtSwvsjg8A6yt51yrS+xPNxg/VpNc+8EZzpvUmu+vg2EQwOWbUrv5TSSEXB
DvUXK5hT7Ir1v7013F+CQFG2R5Avhn8kw6yMqBKQ98RjBofNp4sCybFPpQtikSBE
6xVkhe1gFbJ9TUUkg6nXehDCCg+fYq2ygucGBako30ut751Y8dgwbxwbnZ4YN+UC
1KUo6FmVgRY2X1z17JAmf232FG4VTzkitNnC+9FPRKj0EoFR2x/mTQE+kjHgOIhN
dGE9WUHoCvh+CDk24JkkmjXXL5WGm7DF5qZSkT/toBqUt50nbhsoEY6IvAe8TxwV
oa1cy4gpGZa0rsimOR+rxQwKX2oQqj77gRbPgQgSVyN/dPCbJHygx+HfBe76vNkG
uBVwa625/DJZSrgTwpBvR7+oa8oz81FBM1vGy00VI1MzS9JtQTuXX8mBU+gFSfWO
z77smQ1boN3k7OsmRH7f363O2Mh3xTW/uf0GVw+L84TDOsg6JwZX+ynzLRhr1ccl
jlI8T8Er89kv7954x+M6CDKSxMSvQwtVfmUHNAlU/B7mDUaa4zCt6f/LEhK2DE3o
0hY/n96zoqRaTkCPru8WOncF3fTeDW57fWxkepl1mX3xfaGfA3uIBR7rqJ0dV20F
qPcpDbs7SbkR4eW72ZpPEDWsLxjOjn43T/OUHc3QGSn6EDojkPVEfeLq6WDvKwXT
MxhUZlvO5vcFSa23wGbvS0D6AnaVA1x5840XbDPU1Dq5sM9M1zUvVOWQqD5bWfye
FwiUSjxBDQt3nqbRdZpNnoATrcXZGuS9jabJmQL33uCDWk0alp/nG2OmaRLwTPwp
AHCQRDxqtkjnPRzqGvIV2uAshkSAFSn0JZaknXRatNtZ0DSjTrq7V7fLe5wJOzzk
HZpgfhR9OuDZgb7ut25y+zE8yqz9EYf2JkajA6qXEjV6bosAYR6cTpCzW88BY6By
rP9SVoqPKxibTgEh0mIh2uFMSK80aCDWLZkHI8PpljeR/k54aXxfesRQZwzjfQLy
A/JOrEGbu2QhUXDwaWlZ97/Wa6BX55RXCg9XuGaXRiQBRgKtoDmxM6m3/CpAO2sV
CJFtQGwSUet0lHX2DxRrZppfdvmWtmrmEFS5w9Kv5DJxy69WKOqPqBd5nBCs6sAP
7rgWn87kU7IjoX1i7CLHqb+G+4IZQPMRaptIeuI4byBTEG741sAIO/1lc0dWaGO5
EBLRRXyL3HCMnxRdkC8zTW5vB9vOwT1LKpRlyfg81POefoNN1Z+5ApWMMYsphtP+
WtDEzpsrvu7aUQhjALtulkt6NinqqhZ3VH9ipInox+KfU67GTH66uFawsAyowXpV
MyQHkif9OwbbSJV5WUMq5FQJ0QSJDvmtZWc+FJK00g29YYyLRKUyOEcU/5v0pdK5
XZs0LLZzKK7I3HpE9zqe2OoTfX7xZo/FaaOzO57Hf1lJOPYTe0UCLgg29Al3nA/o
sy7FL+cjStf9nohLPtTbRIaPyau1OR60KRGavEF6KxOg9tMRO3IPI+XOkzKBIrTO
EUCqWs/9EHOO5bY0IilT94l2WA/JGJ01dMyscuWx4tXTrk52gxIJPGirsLYteIou
FIN2FDPSe0x+8l684ijUiiDKVK14zFUJ6ZYLH+OQGusrL2XCHlapXK0Uynlk5nqy
WWw0gob2kPoPClRnhrBD4CnsslbMyaTwTYlrLrQFAn6vSO6rPmXjfAV200UW7nxy
+q55eH3YLwtwtm1blHDmM85IuEajfOI+SQJ+R7IlSS6N7N5uPIb8XtG9b3+zwKGG
WlUSRsNup8QT8P8MBEoRE4mkeHVmUYrL3GVqZbTw0I2lx3JBpFbg41rALq48aTCf
wQKguFjCCQXPjX8hrkyv29TFWeLSVFhbZ0hIMWtUP+48/ief4QigBcGoP61+FXzs
+XI9zC0O/2PoHtZDgU8BSMKuKWHGTcplLCymptau46/4VWLE+Xvg4wsCjBliMVOB
etYjHo+MswLbxRoZw2bezMnZQyLaxwwN+3hgS/nfvgky5uJoZ8LamD/YrgdzK3Kv
dIOQFKrTU5c/keKlZo85wE+xtAbNnh7+GcC0miZxK0oeKp0D4MtI9l9wSFEWeUnP
udo+j9iYytd88omaAUWcRJXRHKmxBywZnrPre9yK9egynl55uSalDrC1Kze9cCeY
q21oPPtoVYCsf9jvgyad1+//sJqDFZUrn20PCL8Tt7L9sno2jJL/Yqozo6LLUjR8
IFPqjv30mpurYZD3QVIjpCHq42bD8AbnwuUK2UsAPXfmUWTjOauOnHWIECI92yDc
ytQlvymKy7PyTKJwCnDFn/pzXLdbi1c7okNLJb8Q5qgkK9f53PotQQqRtWoi/oUB
5SMsls5wn+tcJGGwncIEfw1WKS/4Kcq68n9Niiuc5Wjw7RYJdzjc1ue9xvU8gmTb
e/0CCFnyqE1mPJRC6kLvOvAlcFbpq03DOJlSuHuOlhNIqcSWHN9iTAUZRvG5GvkT
gi3ubVVU0Pbsd02Ak6RXV8BrPS8NQjRyS9ItzzQ6fdxtKrWBswelZx6XGObLwTLR
f/GJWXQRlrOHz3igcvUOzFLqHz0xxO30ubh/lvriHKgozP3SBIudQxrq3JB4vb95
D7Mbj8Kt+JcyE54MmtegQkQvj8+A+/Ns+11VVxo7HDZVn0hBwjp9IBYNjI7IDH45
dD14RjikzQy2ZvNPUshDnxMGWbsI9SuehiOC5bkiMFnIebvxFSmpFHcQVBbGPrCI
tpoq3Te5BgJnjLG/Ibu+4PKuN7JMG2/dKb+FHy9tP+wtVDmL6DxNJ+5PyYZKkfxK
Xfr2QJa5sFB/2+B5sNYLFuPs6O5i93YyO8TtlJt47bXJ37afDEV1tGQP4JKOrWeB
+XmqqkzoaN5rSMUzuCm7BMapHTh4aPG9TPCo6+XpCWFi2uEXWC6By6SAP799NaDv
qcosvvKxqGVF/UMyUq7Fscs4KAWD9uNZL8lQvENqjKM6HkpGG5j7cWdAqXCzIUZv
7LGARu53P5+YSsVLSBXYO73w2RpAjTX9Vo+SrUbEfd3PID3rAdQxqDfIpvzIuJsL
syPut0+KLP0x+Y2B6FdjZxMqe5g6cYCJXmCuf/oEVg9bbtcj8SLkSHzmgRnIhJD9
zsxQsBW3vcwBQra+yUgZqjmPoeGHVCrQbtlRTtL4pw0kYXGQtlps8/MCcvXiCPD0
8YxPqj2vfXl1wjWGKr36t/AHkwd8oLUEIe0Yf0zN8d6bbcvsy+0fRtiJgEcRBhiM
xTSM/UTwdaR0r20VMFH837sw/2r8WX7pfm7fUhZKDi8Wxv9U+F2DabUUZvrUfaGw
OoaZyDtKOwbnHtOqbi5DX0Z1qcfq9v7h22Bo3mHQZvA3roHabtUfiC8lc81meSH0
LZGGkfo6HEW7EY6tj6PnytMc8GqYnqkilnCk40mKpPHT+oKR+67uqoF+Wd0WHAas
VRRiITxytXrLTlz9TGW+R4ehYCwVb2p2/xRTbuxXukDA0akVapjAZI0NT/bpxqZI
NT2Iokiy4xFpqps4NY7zBOuk++LGbwMsHjT5qvvBRd1C1W1A/pUF+sR1TxRHyNvz
a5LVFnkvDrPlAS7xZvEeU7TsmHUOaNS54mHDMrrM+GgjjR/eiq5RQx4M92bARCTH
3F8YkZlYMI9A2eQYSeT5TdKXDw1pJ7buO629VpVRcsaRWBLDrClRso+a5tJVwmED
MRlfunnZ/caoRfpOIA92tsNMc2nwc2fAiY0SRU5mL12xaqg2pSwd4nyMZMX0P7ia
N8cTA4F2kolYOFRdfZTu42rNbOSWcmMzrWTuSFrx8Hdpyvpw3X/+2IIu/HEx83+s
kw9+FN7kwYZXXRIOLXrvi13qsvbEiP51MJk+l77oiien3RdW1Cu5J/chExy9OCma
wOXtngPQ+lFkrQPLL2ys/bSA6ro6pyI4Z0ARliZmmSg7jm9NWh5Rg+PZNBGX/ifF
wvMq8Rgatgxbq3a2uQauoB8YknVqPEbq1P2r3atl8puDGY1ayappCHnsISidt35/
W5C7kRzaDaSzgeZ/lL7gkMMVUQV321niYroUHU0oyfUNgt5Ht+9a5QH3CiRNGKwf
onZcMNMISHlBhhsZZ4AqWIAu5YczY1XJxvZY8oFLjhEOmbtEPT5ONJxzNiQjmqbh
uW4K4vwVENH9wt57LBQs2AyNiA2rkJyCv07uz4H+983B4AZY5YFJ4mL//8xyk+6b
M0bWsgVp7P+HtLtncfRU2PJDenZLWMKCuDjEeZcTLkjEbk8JFNzZamKpts9UGmVR
KoBhYwppOZ7zYEL5aWt+hdv6kbmN2Vj4GVcsgooLwSyrNhkZ8gQ/i3BHsQ+carVD
rIC8cEtibJRuOHLClXNVrnlSaXENNC2sZiK1uEHjW/Pm7t8GbQx2lUhOGbw+LgtL
7aod1GChqnMk1Y9mcS/s/Is3Nh0dvG4jrF+9HsqRKsS6iqqGjwpmN2BYszJq0wbY
xBcXpn3AkKiwFRbjHCLT4OowgljNAkZceYiCMDeCeDdc5BudeqiXLn29w9gq+6Hf
xMx7/tKEf0EZla2R9HXBNzK+bHdzf08kE41KPwIM0XU+SCjFS+eLMitYI6PB5Sv6
djQpW730rBHAkkMRGZtyoQx6BO1L1KcPZ4hq6g/DPCFUFJfLjxWUtUKIBdVa+Dzx
LN7mwMQChYpQ3V/T83wpGW/eHNyJQMwD1KT4PEwJcvTFqx/AEpbXEsflvLKO52Xs
gwgpXWZyqQlE/uXjgZ44QUP8Hev5lUgGW33j73uDFt5VngU8eEEY1HHOlJVAI7c8
CFSXrjYB0FF4v1ieAgUl95QZKPpdtzLUYy/3nh17t33IPu7t9vnXf9lzPlmYJr4l
pe6HmyyhhLuYnBuT/PCpH+46nzk/yFaWJLMPAE9lSR9oBItuOKrYRkLeXwNZdTlx
gMFCBOHi82kJQ/ciHaPTFj7B+4lNXh/5ZIF5j3FDNhAlKYQAIMy8nPzqnpaMyK6b
rhC8sMDtJ2WbLpBssFRwgGiyI/XZp6oDWPAmEYSmcAOs+z/8n7rEcjyA3sFH6hMU
3YjW1oYupCmxVAHRxgyD4UDjcbvGrNOSHusnh8cw8Qdb36r+idw1f97JItVbPZIV
0usHj0hIsbyBsg5DAoSnIznZzThcVBCxtXYA88kTgrttzwUheKhziOXg7tUYztqb
KGiBd26gpVmOXkcQqJRmCC+wG8V2xI1iw5gu7fJDiF3opnQJNv8nwslPAI0wJoy6
OaFdM1U8cHZxlgWlYoSsHpIzuT84wpvPbOaE5dD+tpJWamB/KakwuJLmaNTJH/7y
VTMgtZFzz8JBnvrK4FgwlkEARx9upOE0TqmXsOBeIXNGMbW261rT1RlkWpcidwAe
ry8lSbmncx+IP84vqG+iXxCvVIf6V3K7r/LDnLoljrTjlF0EDLMwBffu9Swm822/
I417cNGZkhuxeq4lM639snJDJWQRGB4WiWbidqPjrnONJiVGgC+nhip1409argBA
J6QFwwlmBRql+19NU5WeMUEX/Xwvw3lQ97AdbcibKtFRflw33f76MlnJSr/KTEit
0J+C06SmAxU3EAdUam5DR+7B3oJbYqd/s/yULq3IatVL4juHgpnHBfobLbaUydWw
QTcWTmIGRL+CzG6f6eO54LvLalCiNlE/ABsUVW+mPnfeNyrJOQgCcXxxzxP6r7Bl
U0WtLQ2N+rP7lXUhP89vAepH0xolfgCgb4Dc2l9FHccTQMo8zeuMWuEYgAuOJV40
MPWD0ue7e8gLOxxzXFFP+fKMMZsSNmfLL9yEu20rib0v79pmDnU+JMDZ06A4X70U
E2wCBinlNf/APZqHHzgUyvfe0CH/OYQa58SG2z8ezgiP1oVta8hTykJeOPQ1UAiP
7HujBYXqQadU3+GGmmgUJb9aaoG11oOP8syPaPAe8NqPHLGW+y7BZ/Jfl89dOf+V
P4tQsVmEMOYDD1x2JSB6AE7Q8v6BXyAymYKL7JWC+Z7bpUj7/VuT+wQkWtjnkYd2
F6AMO+s0QNe6caC22jdPx/CQ45DYvQyhfXlLs9rRtlXzSAySp1MD+isYLso0+OQj
mLRJUNleGp/65QSh+MeuMRtrGo49zv0/BRpGTr1qY3FNEtrRkI52Mw+F95LfEOGj
dr0H1FYiBzCpXefZduPw8WsulnIj/MTuy2uYRUhk0P0yQyKghcYnx1lO+UR4+pYF
n+xdvbhTbqsKpVDGmh/Fna0zZYeAyIRZy3IMwm7Q4MdBtmuCM3dbQvcfWO0l4TRH
24xojLAv36tc1pJS+7J8KNwcKsWkELflGE6ds9DtDyfJaGTMeRsbsX4d9ZKDvDwM
xS+CiekqOJbxox4+Vc2nX2hebVG0T7slS++aF24E617KKCu9AojnWPbrLrNh69yF
9DQhteKj0FQt5f6301o4oLEF7x1QNJJP0TqVLCt29IDN3RukejUN5/b5qzd/Og5G
Er6Dj6uugTyjEH5YqYO2nMqKBZcx555/uHaGgUsBNWN+ZsNEmphuiysKZ5AOxCDR
Yc2Cfz7zeV6bPZi7IhZ3WllO007J53Z+qjhH1vKpD7JxEApFDSsL4zBjT5rfSTb4
SH9a8/ZvBFjOGgLHLydups7VQM8rO242tnwrZzfez2jGAhd58z6I8k5Hu7SCsXLI
Sjlc4mBuIMFYje/8NBFkld/wWZKRvFVYKxoe78IG1fKM8YrLAChtKIAVEPC4OYZq
Qpl/hkqNp1KnlssXvjmdTkxjqieSoCybtJw58HJoeQY9QX1FoD67IV1quZrrdO6i
gDSBbKAyWatcga6IsRWE6UGae7m0duDUPzKBfXpGt7FDd9+xShV0LvK9pDHC3ws5
88xVTuFdXGFjl6msVABBvWg1QRFL6GY1FhiKzgag8iNIJaoi48Tsowyw40hvlbW7
z6yNSBgdhRTr29IdZ0Lxm+UpPAkLPvLsNFgsr6Mpe5w/TihdO/gd4uMhXGb7FbDA
1w1ECq5CdZRZsTWLNM0l5GARFEjGvr2HDfvq8AXvkYDoUrl9YZPXprG4QDPQ3Joj
1OcbWAitGXfi6LhLW0B2Fw5o4ls9Qu3CX3Mr72fMfFQ173Ykkc0cW3SVRCV+ZAUK
x+F3zAwSU4wylcD/vFl4lc9b9WEV/0GOLKlWq+3Pb204lssopJ1nz2jK79Cb28nQ
gdbURIcE9nLP+fBhurh31h+tI853y2/m4dCPBYjYEppTkObJc+7RVE5hSVPxsLOZ
DIA1fn4hqIG6EI6eMaM02hpLz1X4ZykNRsTuws957xcP1QhG64nizie6Yx/aEzQK
sktTqahuLebbSTHnn7vgohbLe0WixUcH8kNZQjUwFkOZ4hrAzQUBt+pX6r6ANlpB
lZbeZyPKZ7RMFTWmRuhHe9WpVmJM+bHqt95EuM0VuY92dOqkuI6r5gtIB6gbXz+o
M26j/ObmVYRrcB6BwK47CUC4aYxmwllNpnnVK7hQxGRCxdYK2p/tfMced+nQV5xY
xhWPSSYkV/gvQQQiIr7RenocMeIKY40FJH9J9yz26ThPlWoAdNNTGxw25ZX+exHq
4wASKhWVRIPDpg7JIS1eLbF7TRiGOp5NfABMVXRs9QZq/uagKRae7gJ9XNFAriBL
TIgrzgjadAmFyDJhWMMcSolx4JvbYYSCDOuemjaQm936vX6xdD6fq/CwGe1hqOfZ
+wamMWmrthWNAPWbdVVUgXsqdnElnPijRdml8fiWDh2nZTUGDHoB3HsxQjOSSdjg
Ue+ZQSgNoq51dIsUQWEscwHMWPGiun1PMPc3UAqpRValwd32IC/0nERHvqwH46tT
if9TOe/V6gpqMVlxTWYyTB31QSkgTYlfWRvnRqcJsa0VbYLfPBLbwH9OBVtl9S78
9W83+n+0eqxRc6eyIuJWG++tuRLWRfcHexxIdwspLTAoxoTyrDiemTqj7ryoUIY/
lrLdcFLOQn3AaIJyDQgbEVMyMoivkPV9R4kVmAmpoOtp3rvquAMWwO0SdH6NiIs5
GU5LVwNiAUO2YAZz7RFWOMgcm6Ar6pj9QQdKmXbZNEfqPx/3ZbJS3wle7/i4wkDx
o4AQW80XIN+mQwkm5lfE17SXTHDfe64dpbFi1eZV7LLXzgIdI7TtEtybFC4Sr9jQ
Bbz7zaGwqQKiwDpNytSIpDQrCB8CZkk7b1qdrTBTzyDUyw5NBCdEBdFeuNa6lun1
dLxBieA6ZgiJoNNWfRsNIkQwHv5NTgTnITqDS3n+FnqDe83+/+NYhS7eTCwLXj6l
SBec0qkGuWc237+bDdi5uxpxK8K8DlFhvKVtScSeJfR7JouUv4fQlpjpoHdmxocv
xoar4gzRdJoPsgvwUjZewXDMvAz0VcE/i2MAc64uGg19kRWAM6V42XKpfBL05M1I
3qTIaOxGK2OMElKk4PhB98H2RM+QguTG0fre+0hYIIOPKijRdu9NZ0sC8ySTKmIO
oSKyeU0UCgLuAXuMGsP/PZ9kPwYfKhtDc9/de1Q9JZDgTEtW3OyBwWN/zOUgslWn
6/vVHcj/jbXOmk20ARn9FQJ5s+BSH3Tty7znj4aC+/0nstF05X2qzItwtnpdMs9j
FVhW7RqIWrLo35lZAqrQNzkcJiJIHQAhSAJs5uq+GMeE/Or8fWxraxHn1eV9BaSN
jdOks1i/OWOgmHtgPpbShFmeT2YQ3tF2w47dtGg0j2LMysIQeRaH/QtNcLt8KIfT
sAGKp8W6HlH/b6dgRxDgR1nvi/Ev8KI4v9gX2OiNqRVy96ddGAs4ack4aYxQzIDG
3YjdqM20F3cYgp029FE4bE8hS7lw47wI8HdFCdPNnyTHIPIG376SWb8tBayGMwRv
Y7Otx6IDwcKlnKW/y/bukicFUIXD0cKXkj/AhvT25apL9F8nlTihPfDQGnddHeLE
85xITHAYECIyGJdnPsmegvwYQpaElKCd7P+FDP0e5o4/piFzjJdevJJyf17Gdamu
sf17l+WGGdQfZ4pWhLtR3piWuUm7C1rnOFk2uaQ0sXAxfjlmQGZQNpCXtiUUbCT4
qW8NJojFK4/0/vzDa1kKGvRMkgVceQR01+IqRq1utq98nMcwPjcLSI+xL55NYYsY
E4sOHabImvIvL/FLQ8G383LuC7xgePg6M+3MtJqg7kpIFlx2ayPibdoMzAxgpySz
vxRMrZfJK4kTzM4huTLKxrUg8kX8cUXgPp3wBsc1XQq15txm9HzjT/3+Om4lz1BR
4C+2GQ2LptFEAQDXAcEhYCLEhEw3E4gc2f4ZySPg9UK5lmATwoHoRQ9MyAcT+9ZU
vLZbsYlFsGTIg+eHKGOzP9bxYQAQUNCoXZNHY77rTBMfFH739xDFAmuo3kaHTIVp
5gwlNwjcDmZWsD9zrJ1vHVUtpxCM7aJAt2AilaUxSMIta1F7sHfloc0JrbMPlOZP
flNBw3d7DLyrwhXrYUvQYHJjEGvsG/94LnSX5gMuej67CCy7pMbOdummLU+Q7Og1
miR3dB1lrthBlDhjhoMxFc/OrZyWhYH3GaDgVROUWikoZ+x3otK27te9QBrW9UCe
pRSZKGL4Zp4RDbUkfI69FPpAYmCPkDOLwrGk03SE0JnTXKiKadXVAeL9oY4/U0eT
+LfFBUCLiVzVkrm8nlvvZGmvWG5RLJ/33uOf5CzcEU8Er2NERkCPgzHxpux72K1f
NBHpv/5PP8S2DKQivU1ILQAR1Oi2rXZpUekTFnFVK6qgICtUjhcaVv84Z0LdG/7M
5zx9Ce6z6irwLFx/ZjSLM+GGoY9dW3GyQ8FNFa2zwqNkcAHbKxH7Ee/skeN+1EwV
pf1+iD3I0BgqEyoumKgQ2slyJ8NLTikBXJjnWXe3flKsYOXJSz1xx5AhnoANES1n
bEpIIX1HJeLOqYGfsg9QfbsR38gLwpDYA6txU2dEndCRRSIXNmney13NQs9LR2/m
n4fyiHb+m4gEDPNAhAXC8RN9uLQj4G9tjl3Nzdp0rLfDzloDLlyKc3hKb7DZ2OVg
X7VhLu3mmQyMPx2CGi6xt5bqJP9NkjoJpODtUCxn8UMOrbRiYt8rKe49UBAwP+xj
VO98sLwOfd0bQUwCv5HkBhAjBGk8BOSj209ELrdnCrK76n6dSpX++mpDVfo5UxEI
sVB1cfdNMrnCvoReA0wW9Vsy68NdEU6ve/NEhYKBK4HPqdrWZTBKo6k0u5EZGOzv
+cEXFP+izY0FYYWQ1SS5SBjcoOP0STXa7esZVeh48t3ZBO+ui77LCymWZAuVomLl
+TouBASOWp8KbSdWV1yOEHVhiHeZ6h1UUAQyCrQhnW98ehw32qTyGKak9xLh7Ci8
JCkzva70lEhzKsvR9C7Inga2/dPrxCjZRvRUV9jM9TJzBdkI6xhrPvfCkLp3vcXL
QMRWZpyl8UXs/HFuIm4wGhuqOk0mFtVMa34KpDLmQz0zlJd+BA5fxs2vJGbnvGme
RNWIbHnp0RLPHM1WRR/NX0vbH3Zap/Iw5+WXERP7YIkhWcZv3Hm1am7NGsSG60py
aUVdtbw+blSEaDV0BhdLzb5rxq6br47E3ZFAmPAfFQaIDMzGSB/G2RPU/Uu6kxKM
cUPUleeVu26uRs4j2WGaiL2ghQ/1YqWoxe8yfeguIS+1OYo7COSXKjIgZxbYHCkP
JCDIubIHXPoFBKdrwrhl+hTJG7p8uLLwaVucUYJl6j7rTWyT1/I+Mwk9HxeVrEtV
SoYfmGobUPqquZ3p4EYHlqGhmQY94dFPa+wkPvpSF0nxo9Lsf+7JfnK2d70Igc08
Fg/Rnky1u/4C/uRkdeaytrcGc8pWmCMq8qOkJENm41eEnHIbzS/kCYUd0dCQpa5N
iFWgUnmcPjH2COZDv0nNmCZOihCDp8aYBqC7RDjbZeGkuqmyk3ewhjGrfVFcRoPq
+kirdBODoR3ckB/G9iYApxsK7iIhSULVk64fb/gSOYe5+vIfLMr5vglvvBH3hwvx
jedDugU8IZk2Frdwxv+77ysPKxGraFD2cU25NTjJuI2fkeYC9N/t45qcuqKQ8Cce
1Zt0L3+QMST25J10q0YBPfYBc+im06vvpbcR3HsL/TIxZdp8HUBnHQpBnCwpwHGF
zFc6dpz34hGMKyzqcVd+61ZP4eiRl3vd61kF35n2SCsMEbJNTTiWPoFLZZDkgPCI
aPTAD4RA8BIIwNlVs9ugx+I+mesQwlwncAQTXoaT5ojHaoZnuWGxiug4okONCSwJ
DRPICMDo3cg4PeYjvuPdAglMjB2kuK9H5tvYYMbuIauOiTDNM6iALxzEfN503ZQZ
GTg9h/zsyA8sit3Uy8v5yGu7/ggDHcTu+7w00FLvnq+hGHZg6sncCZnkEZb9noUF
ohj0Pwg90MR7zdhY0DZ6IhVHu5042pAFlHi2mmJABEb05kNrwrYFeUF4xBLtGIqF
oP7mVVrbQAP6sCgD6vNrvN4+63b4Yw0o16kEptn3d9zUlXRnpDmhfWkl/pC5TRqX
AoNWS40Zkkhl/buB7j+2Go6x4lD3ZqTLkSruuGkPWsJyh2iQ5EZ/Tfg3toD3gG4x
yGqu12TERSNOkaoy/W3ipsjf2B9JCD6DaO5Vkzf6fsnNwVzjUE2U1uV5bweAXX7w
7+Cddy2oFjvpXjDHIjck1sm2B7bU49ZvEIoB8APqa31qCVFuoVzYQReI57pgdJfZ
CHIo/PwDUruobB9TR9H5q5gN7Cv058GuSW0o33AC6SSIJUb0fWjAAhUpeXun9vRW
Ek4Jhk6m6kKuW+XVhFsNPBszRTMG4DRJVnXRcF9B50a2+23ajXDA6Y3GlCPHBMeD
SjqqhcHIbJcIOHuft7NaCeLxZ/qSUdmRYreio1rNYYI0R/Lkq7BK5i0BnDtTsLar
jWD1fDMyDeSwfqa4webbBrOqTDD1VNj4gO2qBBMCRmsbi1Udvw6KD0z0XIL3Z7vv
+iqx0YjcmHBz2vD99cMAJ6t9MdbPNr6fVS0TimI8+t5cf6DCq48ojttetUqbX3vK
ZISpBxu9Rb8D2AvjcJOMrspS2xBUn1pRDGb7NV+3bwAQVwT7QdUKaGh7P7420dt8
3CG1rTwCQVNLaGao/0rtFVgH3lPzh9135b+WWspcvQn2+IOsULbKgnJNltUkMKGJ
r6mvzJvjLMK28bEdUSFDfXI3xvQUFPXVkZHBiyNA+hbKICNU3SxWidONs3nUZIyC
rOvRhn81SJLNZeMTy0e9Fj1iRvftXO/rgbiggnLRLQ842y+rttQzciCiKyzInZmJ
AIppr8SBf7Otfycs7HEsoRfr/vgDdGENdKLgqq0Lbvo8B7yEgvVo5vhdp6xDeIgs
SD1+ISZDpLjNQ9x9yBbWYL6TBMdQoBfTjIdP9CmjTNRGaei3YZcrspydJ8pe/waZ
OEp+kHIeMKSdPJ2mK2kAYVYlqD/qqJCZGD4hgxP8kdxsmkwY66yHBv7IaiUBWeTv
vJ5vTyF+BAe97bhqYOgJPKFcI8KySTlBXGEfgg+I7hwky9ATZDWhk6sMU+5SuZMs
1ebjglpuawaK5qOar4kg2XWbuZbst4y6S0yuDK4kocFpN8kuTAhojH76x0CHiDTF
LmuoGJbqwxo2WpgpiWIEtOm28ifVl/QCEovC1BYqhvG59geeqo8lapBjWSmFG1Lt
DCguZj02dyYmQHMIXzHbSc5t+b3PrKbiyN1G3KBZ9xqSKbV7pjtRJw+5QrXvHHfo
6p5shkynMHPvI0J3IigVIG0nX9MX/Xr9q+6PhUceYI3DPBUtzBteN7DUaRXDg2dP
y9pXHT4szQzvT5VbeD0rDZeAMVFC1MYiDsFrkEoCLp6CS18VwyqSUz5rK62FKmAm
nXRBj7Moc8O5VcN4kHsWzSJ1OzFmENl7zcGzpnlmYal5uAFb2vRLM4fUoSc/Id18
4Ng7acVAIRj8IQfGlpZoz3W3Rsu5rj0dfeYGK+PcAC2q2xAa6Uujy1dAcDY6mVQd
wHK5pWOaRkdFubIu/+z6utUvs88YKXwat55QN8yrnC1R5mwJxkAJMPsxhbYeZzr6
Vo9dvPZz4Ouc6UqEtiNWW/KTWlncCsnYaEhICh6OdAcBGYfSkQ5+uiVvKdSGhQnC
kwT6KjOk0IscmY+Plkt33+qcL+DZPkM1dESBTI/H0oD1OQa/37OFOsS2OMkfagow
JBdjtFPzYQg4dFUUiGDXQSXinFc/b9l3BJOrgOBsqq/WMYWWChNBkq6ZscRDMVKF
x6NKPYMpfR1dwP3ErZKLmO0UEt94ocDVhHuQPs7v1hzpse7ceX5iRbt1WNXwbbX1
pv6UgHXhTkkZG2iRK9U0BHiB9EYP3zeD1aDRFU8q9o7lMjIOpHlVxVqYj2kXQws/
tyeX08yhBLixW9ag66EODkdCMqzJedf+bJhbuKxUF6EYbLmXzjJ7OpCyt/o0va7e
k364cre+ufHs1ud774GTUoTjaBAmtyPxJXRW5onzboIYs7/m4ZH3pi77CxUBO7mk
bedXCewTbdkvI8DV9i22Ba88xMz/xPTPulGAybJEh9ojrGkV7gIAfBq6mkZ5G9J6
u5EhKQPb9nKwO3lEcsZI2HNG1MnmKM9EC3tTz0PDGWA5liJq8QSJ0+uhyiHewZs6
VwYdVpVzDh5jqR84KxDmAS/GnL6FuXIJfaXXCPt07pnn9VOZKauouYA66QN/ND7H
XWxP4JVHRvAlJmSISMW53aO/coUBkCjI8ioQ5fhaqRjmiQeNs3jxQEgKxhbQPhjg
k3mLzI7MbGKYsmtJcHjKuuv/l082/J/R1/h1GlJFxo0zAwmE6bOk9zokTW2gUCL3
7yCWA13gurwDzweeGEYxoYy7njStZKEnAHfs0dY12ChqzsdSSPXRpvWiiOdRu9ie
iMxO3vB13O2z8tQOWQvHiQX4TRiHSwpC2g/qTiQskfYUhvZDNP6IaGzPdmhjC/ZI
GsdE4VpOA/8jYsojSvmb/yCwURalRohQike/nMFB4tcRu/waabXZPgsy9wSbfv9g
6l2J5SoYkHAF5AXs3/ZXn9Sq024MpuHUtip54sbZbhZpOOTSKXc2AijGdVsyHUFn
jJFMzdpvdKcTPf6C4nje73KDexoVN5Pt55RbT/FK46WPKKKjPfFBKqkb0ewAfWG+
ubsvSoNt8rtzPK1r0ooE+wJvF70VRPMJl5klfvsZ88W/jiQbV3PQ2AUxoTUH5om5
V+x6wSaNGhQIU1I/Bg57sVa5+xGknmE7CLPfZ5VX8hFTm3sAJSkGsLfLwR3rFrLw
INUQiE/gtPl5Qm8w3wK2rvckQ94P9mPv1KMtywQBNNKw82WgkguDNelbhoaNfMXy
eJu3P6y60y0XgPQDqTy15Vf6okxLEW23wECAsERtXMFZf5M907wsd13bl/SVMyIy
CRQOg2HrHmGx8pCbv3yaIlQWG2Cwovdb8e5S8nbzkT24k7R2/eXWOBcyUXaZ8tae
8LYabOitoE6iW+DPH3FlOl5jByp5oPunxOa/Ef0mrdylpoP4Fcak/bkVQZMReufn
fDsrExMHQKujKGhp99RJSg3l3rrEYXlkKuM+kxdWcY2XzT3C9G7DblmcvJFJDcy7
TNWZbCjb5uLIVnsmfL3TUsqjoH2h/eMxjMGe/GDZmcTdPWm4yXaCzoKy0JXv7Y42
rds9Xwxp7zL7D7ogVPnDGiPQh7ynohicwygV2CUqdAgQCaJFFfNp08PSBBPAHvGE
5TuipC14m/lAeWflq5TH5mgX/kl6bGihOEhemmhvuMLFfRnqrxgcPHLWcWd064gs
WhFxgbau58Bg2ofjfUqxD+i1E/Xr8Ua1EC2pl6AtkKcApyUcUkR5W97NgMge7jHy
k0LOcQzHXQRbnIxwyiwK2yDUS/TFjvxBKeGQkiJO2LfSiKxZtBYPdES2GzOB/HXK
92twbqL8F/M3J9/Kozv8opUkp02ObzrzrNwZzL9uwlCqKPEU3qu2EY9xxF6JYclZ
eYmeQM5WjoqqbgVScNDb0Fun9lbzMZke8YcuudL1Hyz/3i+W4wOzXwF24EOUVzfM
pI1EVq1G9I9KBHn4x8dvMqFkbAGXc4U6UrKIspRP6j6TAW/kzb19Vm8rKyYtaUaQ
RRGjRgZjcOMCujxPVpmdCZuMC0VneG45UfcFhAdL7Lk34NBv1Wi76hjEcJcxgei9
+joyFlM5w8O+uOVrj4f5fOvWiLK52b6Fxonyn3OsrPVT680E7g1QpegI13awcd0N
N+A0pE7PRVrj/AoJAWoNZ3yFlWN1K4xF0l2xETgiXRlq0btfoeH3xcGptmXndm3m
G1jbJDgYXVYtxV2FSzdnb2GrWfcnDqoVw0LOeSZbcToliAUwdz4CSWI4xAy92AbC
JoX45YgCG/psBbhCL1/sn/IgI3eW6tc03IYu3p4dTXXoL0n4wjN0DEXJue+Juu5N
ubS9Di9RlzTM6hizrRp/aLoOpvNkYZ4fxoqofAdtMOUC/urQmgnQ0I0oYju9efnQ
yMVpgOh7fs5i2W/4yfsA9+AjxnPZrIVFdPW/YaA1ZX1pfJP2kmwOm0AF7YG5K6C1
G1QQTj4i2lr2xFp/Up0d5ksUHftUFkxlXU20p/oGsyOdmuok14Q+jwSPQdj/Zukd
Ak00izWDD6vPds0lSHgDE+dfb27TPw0qn/8FNykE/Jk95b1kKbqZbpgDAUfRErhn
xsQdEGsbTVNnozR7IN+O9qYLLWiv8HOTwtYEAoi0NsQDja4KY47nLgVKR4X1Z4jA
Cp1tirYp+F8+ZrkXRKX8dJUaE+LkXX2aVgXWZ4sgushu/vDvq0zag0zaflGF2EZ5
VvjnTeR2PmFoAxutrUHdlicaAnIUZaK2IVZ8wqm7d6yw5V4msxB7hCiyvvvhEIKh
fcgPSoSIR7yyq0cHrrxDgTRy6C437CzwLy6xL6OeJta37J7s8WvDvQIxOO3QAyuk
h/TmoPnCmUhGClCVmqSspTDNa/cBXjjGDVOVla8t2GU9hVQHkV5C8Yctl6z4Htgs
tDQu9FvVJRWDbqLabaKskR0rhPQTKBI88dtbLeGb1b7FAGLRrRvBbn93v5lCoSIL
yjePO6VrdorpKjaWIeZj9aXtOBZ849EIxnrBdxSOmTUeEu0Ux86gKv2F3rK6AYJz
qB1+YXvi4kw+uiXoRSuyHNaiAo5lsZESgrb+WQJFJtQCQxdu4dS1BSQ3uMHMSw2G
/glYjIH31rN0fFZap1vWY8yyACo68FN0P/KY6LLebgohiaIQaeJguwml7OGOhBiZ
PlgeOw0S8iV0mgMdsFK5/wsoUmFPNWGzP7rMiDpaZPbwFGYJp0Phq2/C62KNCMBq
ZCkVq2b6bTQEr9MAyg8xCtYfePvQ9WaARi/5ELjA7qEyvzL9rYGdc3M18Mq3BRm2
I2WzFvHI1bd8zhmmtmJ57YtnPn5GaBQwkNw69KmcXj4r4FQFibxZLNGXU9Jq2oSE
OrJQ7Gb0RJMSDEz6MyLyK4ThliMvjp7AuFIEs2FcHx7h3Lixt+loZuD8EQLt1JyF
UwlsQbfzPIJ1U9qXvp5FdE5vTqvug+ravIBullpdamMRkHJnEeTAeihJedhEYhSV
8+kr0/5an8P+UCp+kTBurF6FTZ+t6/sfCEiAHMAKZAqUUnEfipSJtKQt6dclsaTX
2yauZMAy50AWo3GgUKL3cjoH3NFDYaM83SDzxMYQjf1+m84/tsIqwgOfsOZjYoW+
0XcGOp0puO7Xa/56rydKeNzWHaz3aQYBq+NLlpldLKe1cxxZ1Djo1/08c+g4pZqJ
5bqpde/70uH0G0XD/UdMNr+3EM9fEDIidduv7ki1DdcV62yyA4b2F+4btzzZMm/o
OUZEYOpSpyt4EOq3GHxn51X2Qftl+iN7g0UkIKAX1vfqyezvwsr50ewoLRHDJEWl
FgoQiKHy1fqrP7YCa9KGpQyLu0gRW+Kxi6hekZfKEqpHKNvqawraH1lHs29pwhck
ZGlFTc/uHSBN9BJ2kjWhSDn0sgTB6h+CUzUSo9Fkyc0qTuusGNPhUNq9BuC5620i
RSsewD21DRVmz8mPr0HdOwtxCNJY46+HCB48nvdyDZn0a0616ZglOKk8WXBTf+9X
kJ20UCaqLxihx1FAt3w4APAVXlZ9SAFJOxPJmJJ0UlgSFRXIADNr8jwv8+5qxEvS
80gOTantEJv5AR66QhHaedc6H/fXbehdzPbCTuosmLlpVXU4ABDYJo+7cOxtsZJt
vnKWbPIBQq+wtJmKDUW80ajsVw8epqaJPm0xLxj6ynDaUDCIvl4U0XD0fXMaXPfX
bfNtvyQL08LMYFJjoWzw9CzmarckkYzwTKzetDGYPWyzFZ6Sph2NNPMBQy8wL4I7
3OkINr+8RzixM1xLO3EAUyVrpGy4mtepLfNz+JRvKrrDV3kl83FBX2oQXzK/j/U8
eL1JNewjOxxn5hHCFidtatjjFwZKKgLoDNjnp7+LpEUVqpbDXO6JA/GmLmJ2d7gE
Hw2vWHVfL2IIIiZ4iH2xzrNRqDZSHrkjL24jMr2xTGZX6xH7PD/btYJXWiLBB5Ln
7L2ZeLbtiwJVWC3zpqWUyrxXrNBLq55fIv7Ai21sPUbvp3YruBejgF0GKGZlabiE
geSoOCc7iVZ2NTq5q/T5gwWcsvD45RiNIQv3dEYr11QHe8WE2VgUaw9Txxe6vJhv
96nONgfUEJxXdAOJ4774VvpT3xhYMLP9c1syLihzWPwehkbNaHwfTeyq94skItFF
YiMmgfWINbN42jMPigz8R0dUNNbxN8btNtprPMpgsrllzqffoaWSCNFkDfo/gP6l
tZ0ieohM3u9YSJU1cOc7BuLH2rT/BtaekX7vmtb/2cEEKbvHIq+0TksHikeZlr/S
Y2jUJ/duyaT/SrQX5Dc+sIkRIp/+Ym/dEGgSixjFFjJGY5dtmiPSkBQXt9B1DoQs
7E8jnhR3/qJB6JUSncwQ6oXyyQ0VzcoC68h4VpcztJ2ZF44reRgTiaaoafmTICG2
Jv9jr8PPdzEX8YMrMkekyMF7glZz7rNGuy0tKYy6yP/besRb6ZdrQ9rg1wh98cRt
aPWH7loxmdYPoJQTOmmur8dmakU9FYCjriqGXrFHHb3aL6Un7dYqSJ1kphUQ8br1
n7YhB5zrc+PFSnuouqzjRgDIOrHB7NxrXLPNOzpvB1Ze70GwIzLLDXdIk/BIBzvd
mrgxiA+Vt/AcScFTAU4/DnzTbAUbFcqT2NHuO+MG6u7DgSK8/FNzQf5w3ljV7eao
SjL/Pl/4H//9YYt1Df4xDy3VYffvGrAhYecSLIGIeMzLnYf1owbJKh3RXDwOtUX/
huuvMvDMMlTh42WFja8CVbBTjbaM3jjsE5mFzPTbvmsWPRT2pzOvoyMxM/XZfvMt
UvPSUT6/Xk8T4QRKz+VILiJWK4juhU0T+UmSlM1u0iHJh2R+2augdc1Jf8yEcvTl
gqwEtR9IvEAX/JsYdXVDVbrUZ7OrF5EqJpgCLWiUCPFZBbnaNLylXxOEEX7dMdLp
a/lU6A6qpvViY3j8q/ngbjnOPnYdO5ol1xyrw/Ewf8gxTJoUB8fmHgkxG30VyHM0
3oXw1tR9+Tp68kpWWMKP8CNElS3lMyrX9De1r/+/kKGjJz89wk6Gil8Z71pgCMO4
RNHyt9n128XpqECkqTl3m6BzOoTXV0FPGoxijyg0XOp0Ik/ubuJiiBbp+JBFZE3/
/fl9fuTSvrzqwfzTDbLsXvzRQQ9Fldz5iuRB7lQSONJc2HKH7B0VjNFAs5EMbWzA
m6xoO1082uFJBx7Koz+9NZavgqHZQuJFQJIA+2IlxyyS4bLeIJ1+3zth7RlomQjT
SGUYtT8lbJNldecCMMCDXZahfFXr/r765UoBYhnH9oXQLCA9dBC8Qj+sItbGmmms
7wWFanLq7s30pH+w8AxRdVWoQLtXZDfn96+sIO38aLJp/CWJ9fm2ORi1WLdOIJGi
dVjgzMHmT0lF91suIROdDDP7vrHhXihgAKY1vz2n8vf8dD3DZiX9NAOqswuRuk7y
KjhN45cTbtBklmI5BUQ9TxNmtl2xtKLiYXjup0b9ufO5c+mCb20f2HiliJOX123s
WjSC3NmIFHap89GXE6QrpBdpAXV6I2azC42SjEIIbd6/AYx+Rugs1Iy8rfF9985b
1nfjjoKqk1XP/ebRWMIqfrJE9WOiPLqWB9RaPVC6AAuFpAWYm6WrjCINf84XwWWa
ZLBx4+VkUgNgbdfLRp8s3xNO2vtleXDBQWldbzLPMNffFttTwMQRqDTHVQZZBZgs
V7mfIZuoSLXN6Z0WcoDW6VRn283+sPQ6Dxo35sBea3qSUWD87hWgml0d6FVB33dj
h0l2AEDFVTuy0ZwFylHAq82t+xUwLjz3YR5KlDzA5rbDnFUHUnMWBsWJfbdbtZJ6
x98NxwfEeL1thXcWWfpv64CZ/ZKQY7V2YmP2K3duJ4onwILdwFnGdON2Yht6YSAq
NlfG7PoT+fQjoFElD36EY5vFAPAfVoi2JPeuNt8GrkmNCVSYLRIYtXKE9hRozOVG
z5vm50I5a4Iidc5f8pfz+GmTC4SHHWtljbRg2AwHWuCcvPLp/NkCUqzM8YbvF054
O0z0A/U9m0C7wUXcNc96LM+QWVzWsuA4M/xl1xTFHM+Cd9F8TZOI0gQjD7Vjh63w
UWUvK1C9OVdXAywFi1CWGtUXltAy81q/CAjHT81HJsC0+25fZucTY1R6IfSuZ0Hx
woMEDaAnZxGyOJW/9Xbz4sUAhsRN23y9dovhFQVdj+ci2QHMTFmn98fyQaa5uCdt
1bSM1xEESweO7Ef/MIrQd2JhSAcs2AV1Oim9KY35ROl3TGe+EmtwlaHeX3CF9fp3
X5VvrbE+PS6p/5nKabsEsA5Ev3u+Pj1GcFYoqJH1Wl/PPpMw6r3/JnjmbYs5XPF4
aTbxW7C2duhZ7hQYEYbu36mwplJ4F8T3xFv22OvlsHc2zmEsEqiycLvG6mhpespo
tNbjl4mtvDndkQw4T4+dRsoLGlaZElG1nKJsZYgSP6ZXDt9bl2ImFfewRfmDLyIO
lWAOFedISOOAqge2cel6qLwtpXr8wtzo3xfgLdD3PPxUvfzvMDZJiX221VRRIOo7
Z7KgaZCuCxEixQ7mUz0jpy8DA3qCq70lbZ/Vyb6QvCISR4a5ZvezRTbgHhQzfvui
3IpBEpblXzvc8+4X0SH9B9mUw9Y5u5i/kvhmuvJMbrg07DvPREiIQx8+X1FJS9lj
qe/Uy//Ezb5O2Wi4cwEEjGuFquwtRmjkTH9v8NKXVlM5Z6MSSEyyqhc0dn/cubKY
gpXPqdcykXY8zQKzfRvF8MMfK7p4LDMGKAs/MQ0Rbh1rImPuR+qmlpJs7UFzVZEl
f5XKOrITI8yo0v0lzbtgL/kcvMpkW+epFJRRfg9GEajM2/Eq/qjhDD0ozeT9ldt3
1vcDPBwPViEF6LZNsbTKyLz9NZ5S+z08QwheR6xVrJEK8o8gq6rPp6/WMmCmDMN4
Ot+5VqmYEuaV/7senM8Ah63uhK911ax36xyEG/Vok1yL7k5YyfS/UsI5erlvnp8R
aJ3YwNBMQYluY0ezR/Ai+gW33o1UrVuTXQ+n26LA6gz2C4L0hvTWhRJIMNBzoZlt
Cfe2TAXS1U1nUGx6/8LerW4aBkG99rshP7VVEMCjuJKERt0MxGkWObCq5AKhhEMA
aCPRXDDyCy7CGCqK9Nym2oWCJn+khFfZYTOljhlTMC0g2uBmVfkV3n3vryGbXKCc
vp6wCymDSeVTotMqd0I5RPscLOgKPFnPPp8Z35HZdjzZ7dUjCgn81yrRM3kmurgb
264YLwhPKq+nhGPcad0nwD4fgkkWlP90sQGbs0zGM8T0CqOzP+1vjNZ6Ew14Oj9m
hG2UwTRZloqgV0Ylq/RuCAzbSrrDhLX30YzC7crYlG3Cf2xbf49F0rNsedNq4WJm
UHQ039EPso46jnzBxUcp7HrdKbHNAXeUX9BuOBIzpR/5fSjiG6D47q8+Z919oLRG
pXcBlsfGQLFvUTrLWdzKKL/cAwi8pLSIt8s/otkOWhat+4x3Vow3BFOtzO1W2mmo
N14oDvQ/ViRZD5HtnHmUYO0EFD9iV4qaFDEKefdHWVpHKrh+rwi81TkQqAqOASIR
HwcqVuM1MyWh5z4D85sMGSv+F2YFX3z83rd+g4CC2bP0dXacHGmlXUWNMJfYMCL5
VYmzoN0A9NeLbrKjI/fjVfLlx0WlWFJmHhQINNMqhguLoTe4QkEpf+Xwl/M0A/O+
On3EDrm5GSKc369PIy5+0rrJ5ldarAr0bZkC3siqNEl9qYs3sadkc70bIZdWuq71
NHIL5YtDMvxaessRPVEg5zTn9+WHhE23FlJAcZq+KFsOW8VKfvooT2whEOcH6glA
nKR45t1UFG/l9CObswTS2D9RaXNnF8LEmap260f332+WG0C7tIhdTSL6QqXtSqeL
ozivViRg6dj1NFNXNDNg1jrmIgWgFSl3kR7YMU5WJ1Gn8gFx8MYOELgXu7IibQuf
HvaOV5yJ7RwrhLRMFcLn0MAt9YLBgdxqpD1Xg3LldnLMHf7fAVdaGL2lj7f59B53
I8nQjgtQe70iyhVFX217Ut/c5x8Qx4KnZo754J0DJ5SXq1NK8a9FUlWOcGHJDSGj
/5YI19MAuIxBFaNeIhyYcrk+aEuHyno+TSRiWhzsLf0v/yLD/rGG8z6CUJks5k71
QZVWG2LYcjVT/KurVPJ2hsxsrel3ulTEfjS2vyHdImBAcRPMwhCVYueoe12E9iil
hSFQKnkIPBbdQjjOUdZmKg+KRC5TeWzTL6N+IrrWEwuaHVMKuqEvT/fS2cDt13k+
e5qgvW8rVFgHntUM3aqduKNrsiPW6s2O4I4piDzpHcaUzcW1J3I0D74BsxopTZRJ
OhyCzs/u0P7jBrXvJPSj2fDzf6ltBT+ETwfvLvVbTS08W7YUeqDdvFOgGKv3dLwT
uU5uOewt846pCgIp0KfjUXhnmKQuQRzo23DoWHPXvQi78rK3ORX7yXyk53tO35Qb
EjhSAV7AR/bQP61vSJNgMcfksb7UZjR9OG2rGFn4DYOslHe7XezLS4qnpJnWci9z
O4/kGuNCfCUMxidA/iHUCTmcE0XLY8+jvvQvoPQOjGmvH/vXR9YOozlJ71N8AuEJ
Jss6YXqQ2kmXJN6UDgd6LmGzFGc6gOaQgD9yeUj36yxpxhzzi/vwrcWBIZIQU05i
xRhOI+T3h9EWhDoqSLgQHZ9EFFiUSCoYS/ua84jqvjCIP9vn2HbFPvwrfD+JBqf0
4/VuP3Rb2CDseYNL9MfoLF1DmrxqnacvmR/6JnYjvkEUROja0q4D8D4oLKDYFkHs
JEQujxW628evJ72LB134+Vcuo/j4j6becjnIkBtWvC9gLjvyd/HFelgSfjjKehtS
c7Ts+kAqt3bdjd1sxA84U4uThFqHLQUL2A9/M4rzLMocKhSjvZmnR+GyRw+2F/Pc
6Uce7XEprxyZOhEVyk7AxcOeAw9/1SRRLv4yBp5vA/pvy0zeYIkiPF8LoAKef6x6
oXpuIcJWXy4PStCh6uk2nsTIpZLJxiJtakCDL+yKrRjCwbCOHrHqIgUPNvAB986n
KlCn1+mrlNpZf3kWify5LEuHr+PdzbK94+wQ3YCgcw5exVVsQXGC4DrZT7IqYtbu
Vgu/bjUmFTZxrgPpbowTEwj9KSOhlIR8A6RYk5/dnDBUDk6pDw8wO3RfUSfMaO7f
1wo9nyF6AkiF9PUL8i0ds8AaquWfrcdZIvxcxEJtMhj3pTBoLu82KP2YUvTiFlZz
YWUO1g95V3cOK+D7n82dF2ORCG9txwwjRMOxgjD0q2hCLqu5QIkLJj/zhM7ofP6j
4dp4Uswr1hEuJCBX/vtwTXjYIhXYTekwgM7BpdnTIv4Nbz4363yA5xI1D1RjniGt
/1xrC/qfcYAWV7TzhFrnnL83UulnIMlNxKIdeKUQjuxzS7Jjsg36Z3w/NRYeiJDh
NFcAKttj8feSfcR6nBKzkVPDtINCubox0pQgb7Qi34s+ZaT1rgCqZgnUT5vBqmja
q8PvkVfu1thIObpx2Vb08UjS4/Q6rSmEHxqyXak6h6QWVTrk3Yd4K3ZngIwIcy02
9iQ8iX72sbhC+ATW2rH8e659rhjGg3v4ixpF8zwjJzJhnQweIQeiuagsCxF97HqS
7CX0ZX4LPzyxz+ZGnvYzFy7RmLpfWgF1nhYaPo3MFIx+Md5jX3DgDG9zcQYTpACA
SusqORW1ajli/78uYGNSjZLstsD4pf0APQRrpiEGxwXn/C8DyvRoqLKrxZ6M03Hm
iJtf1NZ0KLQcsM2DcsBtarzKwC1ZITuuQ+6QnpPLThr/OqioPEf1SicF3nnR4JS+
PcGr9Wf8S8Ts9wOs+gcqPKYZFSDPbrAXnyAaHa7v7BD01pkQJooaIakROzKpyaST
Hj5z4TIMFVdV8GQwWaiufacjogAMqH+tf8wvMDoIWDC6XQCcgvNoECuX+1uz/zkX
lwSQdrYtrlD14qkoue/jPRMKZAHPv6J2TFFG5wWZ9HuNAjeaqCU6hY2H9syPvNLh
caJR9Pu7RMw7Uaw509bJL3CQ4FkjhVAuCNmfY4jjVpXESFQQ8SYXqDfDt/u7lsTV
t1x5KRjE75FNGt5YZKTcREgJXn0E1VvVaiUzBXRh10Gyw3THPmgP8krVnOkRFRuN
F1LyMopzLuZsdzi3hKdyAlOsZ64aM021duyZ7SQM+SHY9hDfC9bFVtyxPYO67W33
mREAAcM8RFbA/01LvkFc2ElQOyvb3FjljyvhhUmFC0csztb4yk0kHGnTgrDG9G1M
5ijBG/XwxgSSLRCZ+Q+ZnJ0JOMwlw1ce9ATbdruGBpXuux1SalSX2zRn6hpystd7
YOBhLo10NroUgtVWGuYnVJqXgpiGEV1mPeb7C18yv+LVWHDlU9EZV6C0OFqLnbV/
NpOoIg8bMUfPQJNcJW1bowG4w8MhzdqUcIFMrsIJhbpD6c8N55wBsRRux4bS0+xS
qN6FkKIhX06oWT9zits0OMunq935m7rKLgGAJ5y58FemBTsy/8UWqcsA100uGL3h
NX5WFjzpm9qzrVMl8ECMXp0ohq0X9zycQxMvyi7uZOoE/5NIbvA/MZfMbHw2o7ta
4af8l9BbTlnOdKFCy5P1tgwM/IRw2WoVwVV4LOIks0BznG0MOx4uiMQvP6QjICfk
a8xDnBeI6OyqgrPVswk9Y0W1rIcRbLHajZ2afBqgUln5AUT24YCBahGan91a3cZE
s6k0sejEH5+AcgTwWjJv8EuWywXetpIEnNb89XYo2dXUCW+85hBowAh4UwHK18Ga
lsA32lh4ji12e8rVnJcwg5MoAYRc5yQXjSa0ACPGqy6KIXgTIXhCTFxi7e84ESar
6WTJta15Vr2RWUZvDD3U4crRCQ4re5SZdmv9GpmxgYBRt4sbfqO48k7uF0XRlBdT
VYA+KhomkqoOYkjAB8gXdKaX/J/NRTs91arOwJhBkbf6QHBfXLtfwwhzd1g0yCvB
1JBT56lzeS+zypbraIZCmwC55rm3SjJuZFykEwXF4XOqW/tPij7FJcKWlsNXajHP
5c93yeKuhYQjqcwlT7yMymYtxpMyiZLefsOuf+SXRA752wa3i0veh5Efhr3HkF5A
a4BsV3rWknd50D2AzMdiMVYgVEfw9jGZI9wEThWr+OAMHY1c9zPovRiq6KlwXS11
DnUUxTfRNaNjWBWhw2L0aDPojbUKGGDx0cTJMpYVs41ggl3yy0dLV6EbRNWU+G63
EdpTJZsEF6tCUDp09aAR7BMREqeT8jStRTF3tbIGqavteMmiJxr4t9uY/4obCzHF
hVV/QXz9ZV+ZVDDFv2jJUYvu20NlY1nHC/YqvhpkPR/0qJKMJi3zOQj4tgmy4BHA
S8QwlgNvHrUgW/7DyxnLgBzC2zPvTvK28I62gIs4+TOdLrw0vi3QdD92UwwPaF+o
EqNmFLN09zVXuaPK4ZJr1VgVEQslDk44vlKRWC4ULqQRItAA70bQTrotI2+K4Sr7
W9ATRXKYS0IBlSiTVDCGdg/Fbul7lrg2aW5X7/vC8O7vf/ZSkDlTEDT/k8fKd7aH
/nWNudeqeeeuqHWcAuMz63Hhb1/ptIicNKROsTC7sauYwFMTKeH1+8Nw4+gTqJA4
6pkIPvJ3nuo4gzdC1DQhYeeDF6TLMIShjeaKJ6ggYpavC8ahi2WNnubGm8o59VHj
S5LsSMw78LTuSf07MN0vJg7/ii/7wIt5qwSAUmiWIIBo0fsqBLI6MzlylLRunCMu
yRiGcvUt6vfmYsgmSGxIww+OUwwX60+PQSb8xQ1LBpLctbviXVVdzFnlvHkV2esT
8q7zEj2RTdlS+ayhcWdoWFWntV/6SKtQZFEnUnHML4IB+ESdHWR/FxCgg5uCwmUW
ZDf9iaUB8I9CJ4GKI/f3wenjLD9LAgu0JTyW2FUdzS0WBqVKug95LxbYtGBHpEuT
qns4f/5QS3lspBi0XBF79ZW9zfaiHkY/LFqV5g8NgEl+Hllk6xykgEr5cS6B6t7u
Msp5n9xoSFcd6QCoTWSlOxQ8BD/vN/3MqLcy79wwsCQQMhzmrI7DEHoEM9hUMNmE
cOoFg3IE0I3xnIj4DapwQcc0Pvwy1JMu6ZI9nlQqMiZgcEq6YppNMeNvZENni4ML
LtFdTxa9rYy2sTiBKqrFeAoxA6wfuVF8vUEZDslVk1XrEmcLYH3Ikr2A/RgGnjlF
RXyxbcOtaF2udtqhGZxE6c2LUErsZt7n6AWEU/IIKE9vrlQslfW+NE6Pem9uSO2/
+YdT18Q4PAOnLrSMDTC5NixRds/6IV5dxvlN8aoAg5x8UIjCgaHskTvabH7esERx
rz55JnMkLjLpQW58cVhj2HXIXFL7xkSr2N2Yfsaqz489U6Mfuzk3cW6VnX4itq43
18gU0PqRe4HJn9iyowZults4i1MoZpAd+cDKJ2M0kmQJgGPl1Hsr3s3bf5DbXknc
cdnQpalx+oDH7skVK6h29Qy83a0U1ekUar9qYah6YIpfH3YfquClm0pEx/Ub6X4p
icLrEDi5+lriOGY84qCow0N9pZq6ECFmcWmHk+BtqyxWEA2w7PghpopudKm5xgB8
uhaJGw7OZGedHHed7ar0aNQNUt7BGNf6rBxzmfVjwpkvzpUkXvdhWT7l8qxgEFGt
8wcSwLrT65RPGkG/WdY/x+kQdq8AFgbS5iutvi46nUxxC/BUxCpBcVLGChUkWj7I
AyqjPSXMgrPlKNc+kcIp07B+G5rOPTx+bvXvxV2S5UNxdDZ4M7PiIlI6QuNaxWHa
3KgtnEklxKa+VQUkfk2PtZfvO5KP84SVFtvRH598FbWX1d1NkXcfUhOPMBt9rnEQ
Ts02uClU6o2M9mIRWJDATSwMwTYY+elSiWOFSI0+1jYHKVFacoRGA0Un1ghEdmB/
unAW8ELwwRasaSdVQCLJYf3Oz84tY0TQNXnQEyM5ZR4Q1DteaeI9yuqN4DiUzos2
zczjQb7YbJxad/BS6t/o68nTpy/gQ1l9kNO/P291YIwm+yEVIV/9WNLVep91YPOm
L4cCjlulTQOsaLBm+SG+jlvaO0NAeuWqdftpQxRCZIz1f/a23Wv9kfF5FrIti8t9
PwX2+PR2aK4JIZgWDTfV2DJ+PBTCWMggLIGkhYxHLFj+mloS3yhWvxzI8P3o8kfz
2e+z03jAZ6XWh++L+56pnDDJyG7r9dxK6R3Qs/DWlfS/bU8IZnb5GcWQII2RQjHU
qpcK30cg84yaRKmbzsI5SPXcHhzwkwucRb1aZRP2T0oYneAYBf32YDjpffd5kfto
tup+2C0Co7zp0BThB8AhhnEdsgEsBXsLkIf7glZtlP3q58SEGUJG/aB8vwcEaU2r
/x3p+Z+Sw9GC95ZkYeKSPdmr4f+O03fEfNTjvjxe1PVwFbfszE30Kgd7+Gp4LADZ
FKj6eGhc+6OaRv9a0jqvJ63KoTOMsepwiYkfyuh8I/gSLwP8qopVMURGY8rrtJDj
r2/rGXtuiWBrmgyokjGuNKXMUAO7LgQIiM512GKJ/anIDy4wJbfSxrvmd75mUVSC
MdPLkk+b0bWjomDK+CSr/0AJLB6j3/IZP5elfajKy1nH3hndDoc/UFrjc/lbpH6x
2SLoqoLrVnb+6sgEIITBjAwFWfMF13L7Zhp5ikeCarDgop7+xyN3JBMaaZhcbp4L
WO6n6qnbx5Y3BCGZ3aAfsAQLJI/iz3BxLJ3SN78icgdFHLWCy+2YODQZWe3nH7TN
cCYdaIsM5QdkLKXM3kRkVijspAPAsF7soUgh8ZGs1/ibglpOz2BUt73WbqIKgnZt
zjJqDbQ4XcMdIAnCMX3WYnd9oW9ViWUE0TcKAPGJuFfm9kfMUP32PWppByb2XZgH
VJahUHdx+lSVZd3fVx4ieLCmQ9Gk0ZH2iInjQbAjk7qADlP87UAv4l1u054vcw0l
eD1GJ0OW6zI2LnvEwjPMiQz859Dl1DooGWh+gvzpFVxGFzoJbjMyLuup8icisem2
gGtHmikxJd0S0m7PQ+1/+A+iQZYcyLKhGhfWGyCl0afjg4x4tYLQUQ3FlkGKGHER
vcD/7AmEuEeJz+ydvcxkSOhQbx9YbSxkD14aOsHQ0JAgCXPtHMbUFinrJebe5Xdv
jpRhnv6ddbymcgMQLyBYyFnG4jSyg1HHj+XE4YsYXmWE/IcgpBzLrw8gcRy+1Y9b
xrzWkdXUKPstViDwI3s49lteCRLFJUtrbVX5qzoqD937tUpQYLATVkMxqO9JSXoz
QNccuegWMqjd7YrFfmHTPbVz+MIGIQOJ9j2SlcTW4WCsyrPbEP4dLcMujdoY9lS7
5tcf5yZOWfsXfeJCyrQW2qKdnWJNBzkpHkV5M53tIvgaeGZOuxohKrmmw/ZU/YVC
D+/VZ8/CNEvtV60FsKogee+ViVAFW4zSDryL78gH8dO/umjR5qpKGr8Qtjit3Br9
QLbIK5/P5O3/a/dg/lJVzg1wl9CDcUGo6Bq+Ihr1mZdRN14heXXwiwd4Aw2FGIMq
207P2kixSQwNizMDHWvy+FZm9GMAAoL5Ds8VCWsXwu3DibYVVsyKDVIBf73KhMYs
w15vLPsvblbfY4pIGE/gyPTj/V/hzk7n1x3IbNDzSJcj3aXz69FJfwV3joVGQezy
4uHkE7sxbwj22x/r8mg5xIh1AsBbBfiLwojPTTpJjoHbucqM3Xcq1nvsvx+yPqXX
+EKJbDTdewZobriSqgKunlnyW5DdXfX2D9kqzlGFmsW2mCMeed27Y624JvHwKtI5
1FSjDf8traGPx1m3nU+hhtTUReFqu3YV23hw6BzoGlYxg5l+enclR2Xak/wVHR6P
snKrpWgTlp12eFrrNe/GGUYN5W9qzXSo5R6mpInYtVn/KFx3gNeas/xwFRMimuNL
/WnABDILvGL874RSl7uzeIaAtm7Q4KQHvPWXnpcJD+H9fEPzd/Zafhnfw2Dj1tlL
okRl4h12X5fj0ErETuUCPgR8dbUyYccoTavBgRhDMlCAzEYI81lOpvtQ7QZOvniA
aYl0KE+DmLjg2gPsEGzG9qZBugPP7rwZjYVCclDPDFUYdqbsEUYtLFcvWhX43DY/
dkwqU6UEIEwkcxnojRmH9Sxe+sbJpxi9wDheyH3gxuoW4pDapI1bN6A3gpRqEUgU
Yp3W7tlysHNEh50+5WEVKV4174X9iTzauOBoIRemNKAyY6c0J6iuOpoAuvcOukRn
FdrzQDrQ6NNHzyx9qjXID164ozFk+ePNCe24KeYSQBTKAJd5v3XJLobT2JwEfSbv
QzUNAmw5KuJ/QcpeL63DTbGhr275lDP/3Ge+XOXCNd+9mRDO7jljyduUbT2HpwX6
k59uTpNrGAYQpVsoKtrzX9IRpHxKbDzxX7/mPLUEE+HT0bisf+kHL+7wcmhxiaB9
dXGZO1xpJqq1inQVo7GnkNkciHu6ZiOfh+Wi8yEwatz0UJuzGSrjo8RCwh6EXAW7
ma1jhh9M79QKM54bzx/SDbTw3PVzwLvkQ+JxxHvt1Q9biCt4sVcdfogcdiFP8VMi
HtUpye+ca/x38eyWohLGUXr8E6112hLyig+PPXwuULMZfPqGzGotCH0AXfF86KCh
T2FPZQWgP3D90hGtXgEyCch54HP5SDZ6ge1CEMa9vlV5tP0qXYdTQ2k+R1NSTA2S
+0xofEKpehDczYxVHsM2yqX7jiPc2gXXwKMhIVO8L+ZRGAnK/yJwnsx8o3Hpiehd
uzM025VHPNlfwwfOjAeA5E+dGYRugIZt9+BiN/VxDJ3M2D256arq6gpcj06mIXzL
GZqC+lWO+WBY32JJK+UQtiBOlLTkV9qO9Z/uZRO03DIr4m6pJElJfFKP3K84HzHQ
duDCP9j8ooUcdsYn7nH9as9LfG9qNEVd0TP0zvmQjLHNs6deHHRzpNKsMVrIYwxA
Wo5dIDHheC4+De1Cgwo3PE4LMGzIZtWswydI6Mo/htx42SwFBKDOJWTfgE/yD1VJ
SfP4kb6yBGHic8p/xSrbtorW/zZBMAkDg3leKT3uyp8CYKIO+eQ6BAzFid+VmwGv
5KCXjjiRg5JfFCqX2ORAPKNyG37tgKeLTq9rAPZHfxQjBRw+mm6pF6298ZaSmq/q
42ZWVdlmEdR/4BuQc55QbXA0lTwlPOAE8CbqFUz95Mmnh26WMfgLfzDOmXhE6Sz7
DwcpoR3yAiUDiK7bLJSHsIvASKC1lavrXJx+gJ0Pff67CmYH2Gp+S63NXWNZSg0P
yYjdV1VFEBJrluUnOB4I7YcqaI3Un5zMyHPBcTz5BujtZja9+NZLumAsca377o8V
9EiuEPmVUpFLYp5Su5dSRLPYwm/PPoXkZovpf9a2FbTjG3P13gqjzm+XKwhhHf06
HBHh9m9FoMH3V3Ztxh9E9MsFDzbVB1NBEcEbq4li3UCSFNVhjNQGfpPeATIgFMDw
h+BolSGfhygQC9UjjyMSQHKtdT50jC0YOl3TZ3rbXAXABXCTjfrDEw/h/T9R0WyD
IBVmm08a/ks46BXU8Mqp9FvC1XQxrvwjmESGXU0QtPhQev1w8JUtg9Xb7sNcr/P2
/EQFgf99uQPCt4isaD5dEZLhs8aMyQmnG/SFeeDJy32JmmTuG1Cd0EZ0JXblXs+A
yJbUEmyl5NsQU0B6WUI7lyWZ+2gKuF6UCS5kn67l7mtSrJXJu4vCom8nAi5oITUA
OE6QAXjzaPoKghCmlS1PVBpUr2O6k43KLzP+1DbG8xGJMS8bqspK0lSDT9jPIQzV
9kMSSMavpBAH0EOXv7sGriRXbv/SsxRTezq3ZXJkxwJljDtqIsd8zJuIW0kSihJ9
OxfRY6RgyG4eKr9/TJjFdfX35hs1l0gMCfW63NEGZ9aOfvR8oMBIDwLe98HJC+qh
xBtQDpz+jYp14M2r9JDPyychplamkNri+JkQN2R1I/QoZOzS94/1WxDHCnqelwJK
d0+6TXYv0C0mpMDbBhBJPUV8GOeLytL5vmxQLlFqHfN+/d3TOdf2kSJsubVsACPZ
FNSmv3tb0sInDPuTd1wuBUOmKUTclIK/+N9cpbxhIzOlE+7dxX028ehWCZH+UFfh
1E/8uGG4aT6ns0jdcYxla4EUk3t69kfCj6IF2Q7uIXOZ3GpOEhPcQo3SqOfmS0Gr
0Sfa3xeyD2+6NdjJIM8oHxzYq80SpP2rOPnYsbvbpT/vJaHAf4MnMt1qrtZCjCiS
mn3TAySolVh7S+nCQZm8eHQwoYGCZEUqJEOrwvio+ivqk7BvKVuqnKgbyNHfdaS0
7Ii6sYTLEBrij6jHj+DvI1mN9nCQRB0ZEnVUiQDZHgvve8kF/YWidqM50iD9s4Ez
jkXXADvj9PQ0hdeQ9ITTbVUVAVSBfAQWvTpUC56Ju29fKPRa6c17T/I3VLf9BHFK
Cn23AJYtyIhEChT8a2a30KbhInsu8D8SbBj/nHO+ue+RgmHfJRQROJBY1dD8XNGM
GJqJ6U8GJ1Nqgn+SmUjQk0jruuOkAfaTOocOsZRDS/tlrvg97WaJnxTrTwV5hfI4
yXSNCGWN5Rf12xUsnqeG3NJcKhymR5UOqbJZfQ6ELvwMQviWrBbbxwDtrl0tU6w7
Uc1BHtF5INc5TQptpgpelYj87HFwS9As8k1/2VE5gLI5G2AMVIO5nAdF4V4u3vj1
pnRR2gqZgUs+5cQkiDOQmUjK/exOf8Zp5M06bbUei2yBSQoiLjCq3cPWJzUG/LOl
IUt4UrITvnpasAHzZcgAkwxQrxv4f4fCEI1Ck+1JzWGblhWdygF5kprX0uF1hBLj
D25P29Ukx7D4Z9p+KMuXWjgviHJlN3jVXlBO7lloMf4fp5xL2kKHsKuOw36vF1pJ
B+Vs3+ixpQyO1SBqyi1oZe6ZQ1A8uVzXhN5tAiR/tTrr2oDyClKdr4cKIjMTq1a2
OSn4MqvO2DdFgZtBURZctm0m6K2WiPFFekvEkSYUNo2hp4T4VAqlzU/aeMQoJqio
Za96/CByQVaKTj+nr+MoeVD5vnRHonuoBSqhfisLlwN4WO0XpmOLPyboaZ+VTGCD
Iad8oE8EFeQFsP0UKgU1qu0/XWH5bSTy6P4L4wpjovOE8bmz4W13zP/XhpbjO9QK
QSjYJqP6slxgwiJ0JTt50b9gqTg2ArGCPWEzxv9HkpJocpAr2pdqm8fsXLetGoSk
74od8eSelgYlBCozjgP4FUfSyWqxVC+j3HdYZmamqplB9uasbooa+w+nbjez72nR
piQCcf++D5LMRaSzj880Pz8UrmDnsVge3pn1NYX2K9yO4RfnK4N3AJXZALHPa5KB
PTHfiFPZ8FBGDMJkyvLu78e3aC99g35Sp06riCpRdUibZdReNOp1xQxQvYgS1Sxy
g7rSvEmterNmnjgBQ+sanBa/kgPLKgUvJGVn0kbEp78U+VaBSa/5+s7JO7VPYFYm
L0vBsWeCoNuse3RMKRvkyDjNNzR44Eum/uVEn9fJ0n3eaTZ7jHVgAPsS6ncRujSh
TuKd+b/djghSMte/KwAxxjTkLJYEPrvDVUfFdPj0mbD2ZbYCWS8Vw7WT4deRgj1Q
Ep+X1TPUCXmjWBbnX3XwowOR6FBQE06zYRD3H9SYA4aoddnznlTm/jr8RAvm4VRb
LTrmcyiDFluWvCzNWrqOZgvJzk3p8atVA3Vgdt3ggDkHqRrUmquwpENHndirjfRW
4NrCXsC8T+THNxTm53wVvjnrhG+nTf4tze9a+UhGKWOMmANa7d6XQFAV3/jigAJA
+EiuobNSHiLlzlTaienvmVdoZkk28OplbWUiBFToZ+x1Ha8TA5E0wZ3LiXXAQ7Jh
cA2KEDv7lbc7DnXUpfj4ssnXjryElY7LLlm7Eiqy4dvrhCBNWw6lnHFOk9PoCdnf
2JjZ/GzM4JTg7ik71QfuAGA6X8DBmcQjdB3Bv5duyUo5uxUOLTvVmJYV2xGu+Ez9
3y03Uiqsm57hJBez99D8TWEAtsC9g1KRwCnr6dAdMEhU58xfIfrFAxIV79J5nT2p
sFLzbArCKdsMX82lSHir2cnOk2LJqUg4i7gJoSfbuAEsiN9cNsXyUR7Z2in/ZVb7
fulk2pUuQcjondbQcffnDDQcCawto9gkNrSP5I1gj/2lhsQeM1dx/fL0VJa3lkpF
44+EKiJG94V5Qb1e4k5tbeC0cquUo23HMVpsrUV1u0qbvQ3OcvHHhTrxHVy1LdSy
bplGD8smB972NmxJC6zaAbDkuw3nGDgZmKwwSyfrrLng7x7SihUJBhInrk8NWFy5
bxZDGS6vDHsKcjHHHR8588a3uajVvNcQnF8OUc9QbE1cZtlkbRlkLz1TfxcwtHNK
ai0cIap2cyu4yq141cCehVNeGMahP0SD+MogClKJZH6Dt0hCYLCCYcoKxTfwCnLn
RLW3bA7um2di+LLy5eTDzLPN85cxkToKZIZ8zsVdgBDR8+L8bx7dzC+zmg2yCTRz
9dKdP74qxf31UJdA7d/0T2DFmas3LinZyNCS8WZI50kKJXIqpcOOYrz/gO5M9ij+
1rxNyKSGwdpCjZbwSruBkXcyHR84PR8x/T2Mmp1UhSqF0DzzjNGyfTmscI7W9c0o
lPBDn2gt+PicGQj4gPRUlKR/oEZ9nOIPSbMwlJukM8fHNKvdea9RCFHWvjHZa7e0
LzjyxM/27imuOlXaaB4xA1uQJvClaJW6aQRpOfuCXq3NU3XQXKTgmtLJCpFFQ0O9
tzJXnD0MHZlDGFZZXWBZQeiJtS8YlXdLmSVcv9IZ44mfWoBGfG3hpIG1vtvGvu5p
2I7gkiWT1QGNZQROn71It+ORynCzoL6x0g4gRqb6uV7HMDhQ0i1OEHaVctOj9iWi
X0cMy8eLkqeEFM6QT8+wnMrlRoHZbUdlYsjxN1ygtEvM0AM+IgipARZgWUIiqMr3
5MJM3T+2Zgasw6a9aK6rmFjiPCLGfzYRp48Zuyn6jebOh3IffCFygn8xuzV3vSil
rDB5x2oWGqa5M0R21Y97xElROg4benGk8WOY0vL6rLDasIhjiakTDY8TddDj5Ks0
rwVdyZMlJqzyOZ2jm79LeZUDEwxqPUSxMEbI7V0ZtDjdNwH6yQVGNtcivXB5iA/W
JRugFylKj5XG0k16h1uOt96WW8byy+3GxoyqcKHN96cnEpRd3Ti5iHiUo+65/9N2
ZFIeu1pazQp03AeFFzlNz1m4coOkTqY7m9QxJPuT0DFXtamjRNw0WC3mp1ecUgNS
Z29hRZ6g7LcB4EVTqRYSBnrrbTLT1CMQ1TA/MiZfTsmEdqlSyhR0uBqSpdxpXe+P
HmFanpGVVojMBYXxEAbkyP6DyiF4ijDqS5wgSm6S+gj+h/RClUfQoyomFt0EJnIN
sBhfA6Qg+g5UQa6KBLnmeSvFOc7MfPA5RJr3AZGBh1Yk0Wqo4Z5H8ZvFuqdANjXe
+G6b39EmlxezAJZ7tEdv+R/I/ej84DyHBW7GPQ+3miqvKdyw7StGv2Mq2cIu0Eco
/WZggSCiUaSXCBhh9Z+vneEf2AfEFPix4z86+qm564NBKBqNpAsXFCcbb6mSpYtR
h3nnrY/WJzqqwPAy5qx0zsvbs6hDo7b/lmrYw+aQ1yz4yvypAxKFxO9v5PEUB7HC
RukWmsLmWO0ZvesjZ5tdGMxAjlPvaXl9hGzBSsroVpWoxsl1SFOFMWCHv2GIToxM
lnyCY7PdIoSBBNwxZ+bIWMZtC1+WWD1rAFIjIzF7rZHTKbQhT1cXmcv5B0CV/0Uh
sqpcN9pj6/3uGaAYZVcg59BiLpjL+IqMquhaS7QxoO/xXMF4QXLQUwKbGstQPHx4
dbcymlBPJAvs54ZyEjzEYjlsrNfECvFRO29aO9m8F1PvgxXq5jypZ6cupCUtGbdU
rGZCBjlwX6r3vr226rQkUDb3BFqos+q0D2Ojzd2uNzyM7NucMfkG5agn1j/vB3F8
1tQGMgtpV2de1EEM3VVscBzOPIPwKqAehf+nYIg55swH3G1TKIicmzbncsMiTyT0
KDaeECWDpA+TbR/w8bZY83z05noVma/2PSW1RPAhSLj9JqpuXnTzEQAmI/zEin03
1JnNlJ6heG8/rA9/Lev2vfaaYtac0kLEV6kI0YdIFumivptxMjz713OOP0738tu+
fpIaHslCyq2/pJaCl0qnb/a2x6CjD+d+kO3y+4LZoRz7XD1iXvPX2c0PKrUB2jwq
EWK/ce5fvHSEG4GYLPPqgJJFtwyOxPf/ieLfaVSdN3tcDrgwIAAXSo/4KIwtgOH0
2AXRQxwqk302lQg3g9NCVBFMMsxxt1swcMsnBwqmBZ2wl6D+55NklPUnwjU62sOy
5rJmMYRlQ73U0SCnj5kzbuw5goMAew9jyDp4LspjU3HuZKNCx2Q+Cfyh+vduJniN
qgPBTAa3Yfn63v7i1loGwMk7BfDNtQFRBkrcxJ0DEK1zLueKpcMD99giRyyoV9Xx
F7t5IW9CsfUpdTa1f9hhJaS2GAyFX52VVCTLPRB+EpmgaF3XP0j11j9MpZcFGkTf
crN1TYlZ19YAIrXqEX4s8B/ZxWpCxxSkzzI3RZjg8x07xUBIgZKkW+qGj/86kPmg
er/ORuKkIILXhqIIIwF9Y06TdVX2E8g5otiv9Ueo4hC3EIDYbQoDeOi1OxI3I5L5
WHReza2ovuOygyWnp+yUen74gfHUV2wQWlFiLTMiUCOgt1l+f/yG/4YMM2O7P7Xl
hJV3/lwUMKIPob/Qm/V6shHN3EdwJq/XH4uaRs92AlvyX4iB+rwkEgSAoJd87JHq
/kzuDd0dtaLwFHAzkh+tWLyof4R5n1X4flc5CCXTfH01TfawAl5WuJGWsNjLbb6J
xlOtJRdpQEbcAcwAA+cSWgvugelv8QijTNdIa49JZmSzTw5Af7QURWKA/yP2nrbG
ki+Vkm+jVlG2hrc3tChbNUP5n6Us2PLCDybpVtUjv23YdCAdcymLPm/meEZ6GgnS
1nBp07H2Mt1wKNNHVSHNFHLFRu7+mTCJkSG8I8Q+pTgJF8SLaRck3Xi6UtCwv7mM
RPUyL887iGwy/FBVO7Dx6Kcq4V+7968ohsPLViX7naCHlYMUI5aYbb40/Zfvsddc
ODpkNlfvgzEB/IFTEXeRgbZomsEDYwuvzz/Hv1pa3Siv+oWjShSfCLoFIaiCJF11
flkBQDWdEBKNFNZDUihLfC2Mio40re197zXzhG5qCAuQgHZeyMJYReO2j+8u9Bgf
uNznIE5V51c11/XEwloUHb/pB3ZfAuu/4CLuMK44Bq80MBjSpvVSPb5rjObV5HhY
8h025KwehtbDDnHxwdQCp8+7r0KYVMA8ND0+6YhMWAQbWRE5GzLsNwc4aTOUUx5P
oWzGlFJH6pNl8VNuoX5JZw8ewPISAp0f+932CxCYurOi2dthMDdDsPNRj3elOAkn
VK2cfryf5dhnJE9ON3wk4WKEB2M44q0hazJ3VSsmowxoV+xihDw5Tir/EgCkQvnX
K/vU/0h1KpYDNeWEWsp1ie4ACJwbBJp+ev3kHYIOC86vhdu8iIOwsvMF2zZWBr6s
Leb0Vl2HicN6UE2aC3CIDcn5PJWb9JVn6t3gded8334/+CPUhRU6G0lQabaVlpeX
ukBOF8MlIi17B23icjB4duuzCZE21A8M/X56x0RjjJ9Zil7pswpkXGOvDKytkGD0
08JPVOz7naFRyjtPGnwd2qCkNWkw2VTKrs0G2/7PhEWauOhtWi1P391oY05ELtM8
vGXh4FQHNY+GiiJBznWOlYNrQ0+5V04CTcCUqjRn9w4ZXEY5+UXLQ33YkWcZyvd3
R02nwEBy9PbkY2kaYBTVw0JS8gWXipxuX5/D6kY18aMx/8dyoGWPbfHneQ4lgZml
Y5mzG3Vnl6oF+MLJGQDJR6mxfRQW0V7vtn6qVhL7Ve3KXDr4T6cCi3cA0UPjT0bR
2UUkM7nnh5nnljeWYGEol8F49vmR9eBcKQUoliajU08f9O5ehNSt2971PUyDXsSG
nzP0biDJiAO6qRjGm5Etd+YlKASCN4Uji1zC/nbuv+g072XJUDTDseaZ/FN4qOCz
VvpvMlATaTnLdyeDJSrrGgXL+M4z9u1l0SXSENoeOJYbvJvphpbUJqxQSu4G2L+q
85yRor92F8a56qPvKQsieuzmdvoqmQdPBZQY8Xwrm2DcjaQzJrXMZ+A8RLfO9lgg
qPsimKLEnksghP5PszYKgraVtybSDAnpgBEhKB0MvogAcdERM78nPyndz5EFBZqH
7iStSRFnPt9Y3TBgoUorSyvflpD9NZZxICNnROl7K8trPuYR+CVOWkcAcFIFGsS2
p1ELR+VCflzKLGm3sL1ypP+Le3KIfwsYTc84SsbT6LSBG8E6d3jX47r4welzH1o9
fKbQohGRAV5dLOCJlHLDHL8wsvYxp3HvjJ4emeVwIHOedGfRyqf9gKSSuWUskiSy
UlolbyEqwDFaPilc1J+8JWjgqk+8VaYJ6awaLEzT8pS2RptG6HQwRK7xqI/PNmsN
6OwkF2aPR2Qmsdz3WAloNW/F2jFNy0O7MDNiFxRDY0TWe/OSN829E1conVlOJVg3
J70gIUhlnjvPrmgDWbd8KQJPH1bukClKmJ3kfV+uJPcVCbl9EzFOK6gAb688q42X
Z5o/1971Izxv+anOn93GZE69C3yW+H33NT/zxxSkIXFRJao6wDccHi77rcFuokrr
7Ii3tVDmUqVjlAL2N/YOrqdV8xV1zMAMTSgsPljz4lkliSNYqevEm0yi7IbaKu1K
3zDztXLfuZqX2a7pTHyI975CIES8HiJDpOGNmSvMcrftXEV4FNtJLCHCITBcjbq4
OBSNfgMnFV3dtBrpC591opWCGaOVca0UPxomqZiRaElJPLWyXbgWAszp7lor17FB
rQay/mFNg/nOLW+cgZ4FH218gQjjQEUXk+iW9NCMdJt0ZwlgzVNvuGQzktHi2a0R
gpwiIOfosIWpHYplT7wvo4oBRIaVS0CmE7P8WGKH/TiuWOOA5OmZ6DrlvuZupeoe
ofu9XDopJEB3MVrEWhDJpGXkYSSfDvXWCvXtNXivma6rToyQz/dt7pspPq096eRN
hhajDpQ+BmrBXBND38Zv7ulx5VgItzAjTHj5hBUIqjToJKybiK6JOkqwMto/R9vQ
9DvvDvkfxLu1O+jOYMHVe5wRW+w9rvTnvLwBEXhRFraxHq/gsAEFXTBCGDnlba/8
fM3HXkuEFKfS9t+ojUd4fcMhhjVsvE7+XT0S9jyRRviD5r6rgpvA5gkoJJKfkCGk
8ddfT1ix8l0RgmeqrcgLC/08XgpPgT171woN8i4PLhZJSt2G9eDIOq4kODVeQnUZ
gN8Ck+PORPWLNgwPFjKJoUbwuYk9zZ9Lod2TDHRwAuBq68TyRQ2uNCi9J4JtfPkc
/bYB+mahCrJod0+qwQszPoH3Qz2YnAixlcSiT6bZB70WgYHqUi2dvO+w8TIpCyTI
aFmiyzwJDMP3uSV/KGzoTdrWNqCVcwJQkhIq2NjsgnGR+K0Jg6gLE7NUv6gKr2pB
RcBtDbDQ5ppS2TO8O57dMNWe6Ll6cMmp2CrIuntXQpMhDBkmT3zBm87Bqus6ROSl
Oxm7UURxSYPDNU9On45mLn6TImaRhl0NQ6GhAp5mOvFjoA3sSRG1vwUtog4O2dDQ
ACemGJOkAZyOxKcdnBkX9AQS8EKyEj+Uu+eYHBL7J9QYmJNzQH0E1Z2oEleDvGUa
6ojPzyyHvT25hl4mOngaJD12epHWrk+4OUvow6hVqtqI3HZMlhKOJc5GJQ8WFzSa
sdqOkaxUNLJFMhPIuvaA61sl/ki1LzQfzjahRJZOPdZKhMB9ROStkUv+U53HvtX0
kVXiRtFid7sVXraQnxT5ygmTTMGMF7XnOKkc+b9eVNtyK3bE3xdPqO8MLL8gv69u
y5i7KCNfY3Esm704+J8J8A9PE0bmM4zMw9f91yNAXh+3tKordS+lgBaukwjf88Z1
9tdfNMBnynfX9FrNlJqXB1oY1wpTDAW/yTvCHTByw1YqNRaJDhTCXsnefJ42JhC/
MWb1XKN4/1oM+bccK505o+pxZtKBJ4UKeYKlYg04hOdAK2szNLK73NNt4bPbIskr
VYMRezA7uXHxSpgfTshAQ9XtaEvj8d1KzYw3b+B+9OdOr57qy9FOGDfKxYBfYlmL
lfiyAz6KfKzStxJNMK9AjA==
`pragma protect end_protected
endmodule
