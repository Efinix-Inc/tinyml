module common_ti180_ddr_config (
    // Clk
    input   i_sys_clk,
    
    // Reset
    input   io_memoryReset,
    input   io_asyncResetn,

    //DDR AXI 0
    output ddr_inst_ARST_0,
    output  [32:0] ddr_inst_ARADDR_0,   //Read address. It gives the address of the first transfer in a burst transaction.
    output  [5:0] ddr_inst_ARID_0,      //Address ID. This signal identifies the group of address signals.
    output  ddr_inst_ARAPCMD_0,         //Read auto-precharge.
    
    //DDR AXI 0 Wrtie Response Channel
    input   [5:0]ddr_inst_BID_0,        //Response ID tag. This signal is the ID tag of the write response.
    
    //DDR AXI 0 Read Data Channel
    input   [5:0] ddr_inst_RID_0,                       //Read ID tag. This signal is the identification tag for the read data group of signals generated by the slave.
    
    //DDR AXI 0 Wrtie Address Channel
    output  [32:0] ddr_inst_AWADDR_0,   //Write address. It gives the address of the first transfer in a burst transaction.
    output  [5:0] ddr_inst_AWID_0,      //Address ID. This signal identifies the group of address signals.
    output  ddr_inst_AWAPCMD_0,         //Write auto-precharge.
    output  ddr_inst_AWALLSTRB_0,       //Write all strobes asserted.
    output  ddr_inst_AWCOBUF_0,         //Write coherent bufferable selection.
    
    //DDR AXI 1 Read Address Channel
    output  ddr_inst_ARST_1,
    output	[32:0] ddr_inst_ARADDR_1,   //Read address. It gives the address of the first transfer in a burst transaction.
    output	[5:0] ddr_inst_ARID_1,      //Address ID. This signal identifies the group of address signals.
    output	ddr_inst_ARAPCMD_1,         //Read auto-precharge.
    
    //DDR AXI 1 Wrtie Address Channel
    output  [32:0] ddr_inst_AWADDR_1,       //Write address. It gives the address of the first transfer in a burst transaction.
    output  [5:0] ddr_inst_AWID_1,          //Address ID. This signal identifies the group of address signals.
    output  ddr_inst_AWAPCMD_1,             //Write auto-precharge.
    output  ddr_inst_AWALLSTRB_1,           //Write all strobes asserted.
    output  ddr_inst_AWCOBUF_1,             //Write coherent bufferable selection.
    
    //Startup Sequencer Signals
    output  ddr_inst_CFG_RST,   //Active-high DDR configuration controller reset.
    output  ddr_inst_CFG_START, //Start the DDR configuration controller.
    input   ddr_inst_CFG_DONE,  //Indicates the controller configuration is done
    output  ddr_inst_CFG_SEL,   //To select whether to use internal DDR configuration controller or user register ports for configuration:
                                //0: Use internal configuration controller.
                                //1: Use register configuration ports (cfg_rst, cfg_start, cfg_done will be disabled).

    // DDR to SOC
    input   [31:0] io_ddrA_ar_payload_addr_i,
    input   [31:0] io_ddrA_aw_payload_addr_i,
    input   [7:0]  io_ddrA_ar_payload_id_i,
    input   [7:0]  io_ddrA_aw_payload_id_i,
    output  [7:0]  io_ddrA_b_payload_id_i,
    output  [7:0]  io_ddrA_r_payload_id_i,
    
    output  ddr_cfg_ok
);


assign ddr_inst_ARID_0  = {io_ddrA_ar_payload_id_i[7:6], io_ddrA_ar_payload_id_i[3:0]};
assign ddr_inst_AWID_0  = {io_ddrA_aw_payload_id_i[7:6], io_ddrA_aw_payload_id_i[3:0]};
assign io_ddrA_b_payload_id_i = {ddr_inst_BID_0[5:4], 2'b00, ddr_inst_BID_0[3:0]};
assign io_ddrA_r_payload_id_i = {ddr_inst_RID_0[5:4], 2'b00, ddr_inst_RID_0[3:0]};

assign ddr_inst_ARST_0 =    ddr_cfg_ok;
assign ddr_inst_ARAPCMD_0 = 1'b0;
assign ddr_inst_AWALLSTRB_0 = 1'b0;
assign ddr_inst_AWAPCMD_0 = 1'b0;
assign ddr_inst_AWCOBUF_0 = 1'b0;
assign ddr_inst_ARADDR_0= {1'b0, io_ddrA_ar_payload_addr_i};
assign ddr_inst_AWADDR_0= {1'b0, io_ddrA_aw_payload_addr_i};

wire [7:0] dma_arid;
wire [7:0] dma_awid;

assign dma_arid = 8'hE0;
assign dma_awid = 8'hE1;

assign ddr_inst_ARID_1 = {dma_arid[7:6], dma_arid[3:0]};
assign ddr_inst_AWID_1 = {dma_awid[7:6], dma_awid[3:0]};

assign ddr_inst_ARADDR_1[32] = 1'b0;
assign ddr_inst_AWADDR_1[32] = 1'b0;

assign ddr_inst_AWAPCMD_1 = 1'b0;
assign ddr_inst_ARAPCMD_1 = 1'b0;
assign ddr_inst_AWALLSTRB_1 = 1'b0;
assign ddr_inst_AWCOBUF_1   = 1'b0;

wire ddr_cfg_ok;

assign ddr_inst_ARST_1 = ddr_cfg_ok;

localparam [1:0]    IDLE        = 2'b00,
                    CFG_START   = 2'b01,
                    CFG_DONE    = 2'b11;



reg [1:0]   cfg_st, cfg_next;
reg [7:0]   cfg_count;
reg         r_DDR_Reset;

always@(posedge i_sys_clk or negedge io_asyncResetn) begin
    if(!io_asyncResetn) begin
        cfg_st <= IDLE;
        cfg_count <= 'h0;
        r_DDR_Reset <= 1'b0;
    end else begin
        r_DDR_Reset <= io_memoryReset;
        if (r_DDR_Reset) begin
            cfg_st <= IDLE;
            cfg_count <= 'h0;
        end else begin

            cfg_st <= cfg_next;

            if (cfg_st == IDLE)
                cfg_count <= cfg_count + 1'b1;
            else
                cfg_count <= 'h0;
        end
    end

end

always@(*) begin
    cfg_next = cfg_st;
    case(cfg_st)
        IDLE:   begin
                    if(cfg_count == 'hff)
                        cfg_next = CFG_START;
                    else
                        cfg_next = IDLE;
                end

    CFG_START:  begin
                    if(ddr_inst_CFG_DONE)
                        cfg_next = CFG_DONE;
                    else
                        cfg_next = CFG_START;
                end
    CFG_DONE:   begin
                    cfg_next = CFG_DONE;
                end
    default:    begin
                    cfg_next = IDLE;
                end
    endcase
end

assign ddr_inst_CFG_START   = (cfg_st != IDLE);
assign ddr_cfg_ok           = (cfg_st == CFG_DONE);
assign ddr_inst_CFG_RST     = (cfg_st == IDLE);
assign ddr_inst_CFG_SEL     = 1'b0;

endmodule