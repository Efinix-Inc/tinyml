///////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2024 github-efx
// 
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
///////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ns

module axi_interconnect_beta#(
    parameter                       S_COUNT                       = 3, 
    parameter     reg               SLAVE_ASYN_ARRAY[S_COUNT-1:0] = '{1'b1,1'b1,1'b1},
    parameter     int               S_AXI_DW_ARRAY[S_COUNT-1:0]   = '{128 ,64 ,32}, 
    parameter                       CB_DW                         = 64,
    parameter                       M_AXI_DW                      = 64,
    parameter                       ARB_MODE                      = 1, 
    parameter                       FAMILY                        = "TRION",
    parameter                       RD_QUEUE_FIFO_RAM_STYLE       = "block_ram", 
    parameter                       RD_QUEUE_FIFO_DEPTH           = 8  
)
(

//Slave AXI4 Bus Interface
//--Global Signals
input           [S_COUNT*1-1:0] s_axi_clk,
input           [S_COUNT*1-1:0] s_axi_rstn,
//--Slave AXI4 Write
input           [S_COUNT*1-1:0] s_axi_awvalid,
output  wire    [S_COUNT*1-1:0] s_axi_awready,
input           [S_COUNT*32-1:0]s_axi_awaddr,
input           [S_COUNT*8-1:0] s_axi_awlen,
input           [S_COUNT*1-1:0] s_axi_wvalid,
output  wire    [S_COUNT*1-1:0] s_axi_wready,

input           [bit_width_sum(S_COUNT)-1:0]     
                                s_axi_wdata,
input           [bit_width_sum(S_COUNT)/8-1:0]     
                                s_axi_wstrb,
input           [S_COUNT*1-1:0] s_axi_wlast,
output  wire    [S_COUNT*1-1:0] s_axi_bvalid,
input           [S_COUNT*1-1:0] s_axi_bready,
output  wire    [S_COUNT*2-1:0] s_axi_bresp,
//--Slave AXI4 Read
input           [S_COUNT*1-1:0] s_axi_arvalid,
output  wire    [S_COUNT*1-1:0] s_axi_arready,
input           [S_COUNT*32-1:0]s_axi_araddr,
input           [S_COUNT*8-1:0] s_axi_arlen,
output  wire    [S_COUNT*1-1:0] s_axi_rvalid,
input           [S_COUNT*1-1:0] s_axi_rready,
output  wire    [bit_width_sum(S_COUNT)-1:0]       
                                s_axi_rdata,
output  wire    [S_COUNT*1-1:0] s_axi_rlast,
output  wire    [S_COUNT*2-1:0] s_axi_rresp,

//Master AXI4 Bus Interface
//--Global Signals
input                           m_axi_clk,
input                           m_axi_rstn,
//--Master AXI4 Write
output  wire                    m_axi_awvalid,
input                           m_axi_awready,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [7:0]           m_axi_awid,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [0:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
output  wire    [2:0]           m_axi_awprot,

output  wire                    m_axi_wvalid,
input                           m_axi_wready,
output  wire    [M_AXI_DW-1:0]  m_axi_wdata,
output  wire    [M_AXI_DW/8-1:0]m_axi_wstrb,
output  wire                    m_axi_wlast,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
input           [1:0]           m_axi_bresp,
//--Master AXI4 Read
output  wire                    m_axi_arvalid,
input                           m_axi_arready,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [7:0]           m_axi_arid,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [0:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
output  wire    [2:0]           m_axi_arprot,
input                           m_axi_rvalid,
output  wire                    m_axi_rready,
input           [M_AXI_DW-1:0]  m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp

);

//Parameter Define
parameter                       DEPTH = 3;

//Register Define
 
//Wire Define
wire    [S_COUNT*1-1:0]         s_lb_arw;
wire    [S_COUNT*1-1:0]         s_lb_avalid;
wire    [S_COUNT*1-1:0]         s_lb_aready;
wire    [S_COUNT*32-1:0]        s_lb_aaddr;
wire    [S_COUNT*8-1:0]         s_lb_alen;
wire    [S_COUNT*1-1:0]         s_lb_wvalid;
wire    [S_COUNT*1-1:0]         s_lb_wready;
wire    [S_COUNT*1-1:0]         s_lb_wlast;
wire    [S_COUNT*1-1:0]         s_lb_rvalid;
wire    [S_COUNT*1-1:0]         s_lb_rready;
wire    [S_COUNT*1-1:0]         s_lb_rlast;

wire                            m_lb_arw;
wire                            m_lb_avalid;
wire                            m_lb_aready;
wire    [31:0]                  m_lb_aaddr;
wire    [7:0]                   m_lb_alen;
wire                            m_lb_wvalid;
wire                            m_lb_wready;
wire    [CB_DW-1:0]             m_lb_wdata;
wire    [CB_DW/8-1:0]           m_lb_wstrb;
wire                            m_lb_wlast;
wire                            m_lb_rvalid;
wire                            m_lb_rready;
wire    [CB_DW-1:0]             m_lb_rdata;
wire                            m_lb_rlast;


`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="ipecrypt"
`pragma protect encrypt_agent_info="http://ipencrypter.com Version: 20.0.8"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"

`pragma protect key_keyowner="Efinix Inc."
`pragma protect key_keyname="EFX_K01"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_block
aLGMEOXskW3vMi11+2marfIbswuOaWn5lyluxhRdPbXe7hpbIAi5vH3JBHImykys
TAz5LVEHVVyWzV9J7wc0/Ihe/7WhJNSNcKeKnuTVcwiE9AkIqlTKfvMCvPsXf7Xz
8EqAfdCnU6wqjrVmafHg3Z4JaMiUD0ZFvBolWG0gOmbzRdTmOeOb1cpy5CaDulOU
yLMdfnULBbhKfjUuVmZrPUBKrYaDF7juB7ijqZjkgINfC5Ivw7IHP7W0PDQvlX0q
SCNR1l/mpQB31TlzO8TapLzHMvpsRZ0qVkq+xxhEOdc/HLK9FF7MXPRFtbj25OhO
6tdzgTczPJsQCxrS8W24vA==
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_block
RkqCl1xdMtIcP0wjALJvqyTtlQvr8WynQHBmvEiiL7HaTh82l8Od9PHHg3T4nfrp
by7JTlLBvW52VnkBGGVVKlDuzc6U6mB1PWTxPs48DFfevDzuuh6TD+379T4xgT8R
giuK9FzUdSMhuRHLphlxNCKqVtEEn0AuUrPkbahPtSE=
`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=19456)
`pragma protect data_block
eB47qOTJDM+fdV2b4ke/bYEiV/yY/U6WxWgWACpFHOYMOEx2mbCp+qJfUf/qV4a6
hxUy4KNyPStbsyxZiWMmzGqZc4M3C6MmIjz9z7ZpG0HZ0oxfOov8VoYvI/hO6Jqk
z9E+03HwnN1IDE/4RSxHsBZJXmkxaGBxSwj8sLa+jT+YAkuoUemiIeC7ZgIAPABd
Pe6tzhgtcnBomYPb1YgXplcLxZdfUPZ5Cu3DKnH1CmQv6N+xj65Lb86+9bAbcefq
XA97LRchTcz4fMhSJaIe1PKroDqhRkyHYqVoNUcr0R8cs0l8irAnyq36BlKzplKB
32LQTbH4OvRhT3C2BJiW+kEf2W/lgc8sK22qcf0v2nMN+GhdklcVnGLAZlqDMTY8
lHzlYuy/NilB5jd+KnqqH6WgLgXZ51578DsuKnCSFAWW4KDKVuaILfBtXEllhYis
pvyVuy+Z0rsCK5/Z/xyPdep0Z7lK0+VwyprwOAgtvyIA30zUQndOvfo8/1xY519t
5eO6s2aCeclurKAc1byZLU+C48bNUQpaOzuBSx0hzwE1rYcYuGxuDh3Vg0cPR4co
GmKbZYfOUt6lMMoodDMRm7GZbNwNQcFa0n4oZsJmnJpEJnaFxK8ZsFkpn3GVCS/A
rrqn/sd3+HsYtUKhOFuo+OeBgcshJ+PWrkfN3QT1ukBMnRoZZWs8MFd26SFHxZW5
PFbx+tsAYM3cyTuW+y4a6He0lWmlXtlFjiYF76Un7k/q4wB2KQTAQNfiA+09ImV3
v5xeGdman9mAgibSnaSf2XpCybcp4u3U8vulVA9fOa+9YGiEa8fakxWhpe6Lki2a
dr2RxemQlOHc2lzgMO6RcTVVRoCM5Pqfgy3Dwbr40SHIqV+CqAqJw7G69HKm9Sh2
EXLAUbTin4GHm18Fzx+z0PRdL+7v5qHz1Mo1sbUjdrJgc3s/KOY/g0PWBvUT8nmb
URI+AuY5xvoNA4j0WhCr/GntEurHeuBX34lk2PwXnHlhWvcs071lveeyBhrJyJiR
iIIf9XfN0/3YAcBPhjTXw9OszMa6rx74K/G48WcgRmILjwGYrgZZtXGYkPg/vDTQ
BAyn30QAsipaWSgocXJDh5r6kNkCHMhddeziQRyysorUjHnSsIttfh33DZGt3tu7
YuO27YVo6OXpS/XJPA3Lkn9ezBYfORzIoETpxkw/PytaWz8hEmG0CupSxufSLb8g
M1ByVAlmgH1FEt6euGVUQnqn3K/d9DK97nwBKLPGuF4q8Gu86NEYHiXpJkU2nS2E
ekIgqVvrbFTsMR8md1uMcj3Mii7fZ8+cfpXwH7Ms0jzB2X4egUjKQ+cDWeQh5e3W
lhqohJ3xKbzE+kj4tqSNjlFBSEEJgBAMFeIWEeTRLi542i8oVMI3WIBBdaphsjMT
vBdJGt7Bx+SsN2i6RkT0FIinD5a3Tl1OVxA1YyIoVhSizbzphVzDXudpkf/rGaxW
NEiyHhkVyIfVkUrWMRaNG6wkcW9QHXbC3Gt8KpVDhMeV+kyFkLn0uQX+mYqkxp99
b8oM0eLfeVa3Wk+MQwgrCDoV00mVToBKMH+bJ9AzJCyOHWps+IMtKcwGvI0XvMZ8
5wUgFnihIWXAZg/pisC3Csq2jGeNugjUAKjIMkLZHTsv7hMhZev11OpIbskMtr/a
YbEVFEh7l31emI/O0HqhOt8d+ninjYnjEt9YT6LT0eE/+ph93DAPxrP33d++2mqk
resmJFb217E9QZoWlDLVnr2W6FeJo1fa/CbsKMOEAaIKbA4MvuDA6Fj70ED7KAwJ
uQDYvVG8F2KjZ0vDPA+V+3lNiP/DbfARr7UATjdzuGGhSPOZG0rHQ8UfzbdoOrQD
wn8FQjXxR+GGX8qwAB9b1+Jkwzzb1qXRe22WWYwuGMoYhKWxZDk6i2imao2hwo6s
MEXghvizP6HkOKathz776BwQKPFrj+0ahrWxzkOH5bFrzCS3wTUPBhIOQJj+icz1
8yQii/Yz0E8zG4FCxUz82y8b4Lg3qjvWqVsGWkSdcE6GeimN1XHVqTlWd1zKeI6r
31w1KJc2tjYb0YsxOX09HlvqJkgcJz9+PSIjMD/D36XHaLnDuYXXwrie1Z3ytcv1
h9QAvArbiBdX2OQsr8EvyPKVLIUOtSYUaZcXwG1Sg96AbsCAvc6pE53Q2gch/oE1
43Te+QamUMDqeZj1mLF5YGHYmJx9QZPAE5gSfjdl4I6xP/DtocGk1AzEj+gjYYUk
L19gx1lRYTAIIT1EZZ6QQ0BYpx1mVTnioNLXxG89P8M2G8faqMaB2NtUofv1PPFT
d8hMQENmlvt5cS3hxE9nyyBxtam4nB9lbV0v/c0EeOyTOqKS/k0ofANvORcoTFYJ
X1/hrMybt4MRAy4clJ1pdmrRNMmalb7A44EYqnqSYTr+xnpj5EztqpjIh9CQrM/s
yN1ZaFLEF4vtKj1NFPf9aRuqQB4BET/o0unUc0EudDLG8sDsVB3JEGVo1YwG4xVF
Y12bv2RV+S34gUehdelKw2v9ryUp8vruvGB6hZFcdsiYWr+cQzF7f93qV+5lRqMj
G7i96IVJzmvDYHTH8JM+/Xs1GysEsB6QkfE+l1fcTG5cNXZNqPBT+gxPmvuGJHve
vDTw1IITx0LCfnkF/HGsdtm14VKtrOUH1K2BDkRFbO/Q9KlxjGeC5UXqo9YXNCbE
tCPVYPjDxe75CLLLAtbkkYH7QWmLHsOtJjGv7Szg1Q8shSxc6C+79sbIfuX9u/2D
1S4osHwQlRF58fy9oBxw2k4mxxuRb0aOPG54hNsgfsz9hsH3JBfFaV8OowzzNjeN
QvqSB5sGqJTlTHg5NHngDCOqvJBbuoNmby/0Oc5Zq+2iVgr2zaOBGjAULOF3dO2N
Suq5GlT1kUAxiuokALt7H5v1mPzn88/UYrAK9WNFOKji6/n9/GxjVLCFLuBSKihc
048FIn0OVhNu8AhQV54i/9SBLfbkhPhRqge1N4LlsrdaUTFL7AcYvDNJxrx0/h94
eS0e8izA+plDLiYW90SwD0GxZi00zSCdZYxVFNHXTWY35gZQbkHTkvOoBIMzyT52
pGDLlUhHrreUWJoyxCQIkMiLAEyZChGNsFrbQOm7M34Jdxfy5u4uiGTQC1aN9rLO
4BdNaSyWc7oKOYNpKMgZ9xH/KPgTUY9EZH6F1lbnPAKorOh07PB1hrKofwm83EVz
OFRCJ+wVak6zFWsQmk2x5WpUd7LSygWHbShFxBdMAEzGD0AvdLvmyKeNR2HJcOI0
ycQ9YntZKzsOibl+k/rrHxBf+qsb+mZW7po1Dye3UGW25ptEP7FH2vXp0MWbdIPi
LJlL1A/Hu9TTPLoFag+A9T0mniaSsEpnnNJ6lDFoN+C0yyBR6hUXpkj7CU/5PMlb
khYT+YjPuotbqBhJv8dORVyvHo1ic1BgVNxAJslPbv/TINMkPdMR+YIK9Y63k5xV
4tNKgiosWNCz+/BzswI1mIAwP3k4CEJ4hCaJ/tEnGA+o6ys7Ml3Wucvekh71Gdp6
NRSJfLLetMzSvlbNx70k4BAEbkTyo+ldI7tTV761sk+f+Zlq2kKB1k4zOczzGerA
Tw+uXuo8WuCpwXG6A1U0MhhPpXJAomS1OTMxEyhhIbODitSr6lrtci2+oZbUrmmx
NBiAdrejQP/5M7Sb7HJE9n9MD8MPAX/xWLRoJ09FJMJpLPNXOZIwNOYGnPfDrK09
RgwgEM6ukkphikwtS9qDRyyYBSzxZnMn8K0pPuvrD7QovQ3t1Hgebszte/SChKWw
I29Y22moyOv+p8llm/lVASej8OayNvDzQg1NpFeVix2bNfE87FzIZCVPHG6WPd4g
mkg7ljNrwFuvq6gG5uEyv7L/g7KTbgHQvFnddU/o5tL20HzHSjN8W6qhytsw5uS/
bRhv6O/TAUFzvr8pZK3/da45yDETYYM/1miTN5199+mZLp1crWuh2hRKxaL24WKO
2i+U3bvjClwtGSMHTE5ckErKHPOjZYaQ8PmkME8zRxUfWbv68iIJ8wEHmO4FvLAK
S9+uWGp3FCCBsgNWqZnBpugcxvP9wVCWWCKaAlvRPuU5/0Qu/OuP0VvczfrdYHtx
eJyi1QMxg/YyaPDzYbVqGOmVQv0MPo9epI5JHdPb0QK7nHYeWKMKAgm3EVwI/3J2
pfDGGx5oHLc2AHk5P70ydwOj8GBCzZzVd9q7/l376/S5AvG8/zRlxCDGHznu6pgL
CqmgolF8OydpBhDeXTL3fh1/E7zff8UXqQZNUgdUK5YMlYG7KCzr1akiO/zH4Kt/
6CaN2ZMjL7itAWGjPIIQ4SfwAq/DGoqGHcEDg19YirqPKjgq3vp6Ns0rzBU9nLYd
8rJWGFESp1CLah3pIVj7dRVYWmk/6/OOmLS//h6w1PEmiCT2Bo5WJrhxz/ToSihN
7X/Xr6HoJNwZUD0KSNWFQm7bmZyy2axD2zzKhQ5bomjllf7Bpm/Ce1JHzWHd8NNg
1shfgrJX1dZ7ezWW7vNl4ayygugZdSy/3f0GviHPX+gvAnOvhpjb1FJyysWBoH6P
e3AIDCOOpJQmD3oXuWZKN5f3CEB99tba6bLJWiPsnQfF9Gh8QMTH2EaJHDZe1WIu
TviDsLcHM22QTcRFsLQYjfN7b9bA/XIEFK4+ZFlBibx36cS0A+WbZXJ2Gwb/MKpB
+03ArpZa4Fjofh2zSGG6XZilxBMmAMFcyYZu8n7TJS7tJyZg6OelPXlNDox+ymes
M3Qi8KfdL5NsHw8wnZFkdOi1/kXueimSbM+inACeoAmiJZ3TJxIBlaPhTbCv7XoU
6+vy/lMw8hKX0f0fU8KXrQDFs6lJ1cr318EFJkOEhZVIABy4ba8QPcEF+7JS7LbP
neAfrZG4x+Go93sgUSSvUnOeFOeK1Z8Gwqlvb+hYLSbAPPyCa4eN0Ay0C0JGbiPu
qag4b5qBeavqwXtVgUu02kYgYpzSUGCGpmDiNBGzsQcz15N2YHHPmrrTHHTmEroY
sx3Wnw4lmUl063WrkabxtRrlywog7ISzv3JdRUxq+xZb+mIk1SEq78PEbOTDXXXh
7fiGRK/Y3wsi7pDeLhCxMR09a8T0j/D6l+r0u0WnROrLXMkHIgnO6yuqI5DyLL1Z
L5tsNwEP59yP42JIhtXBE0RJSuO6K80p1K5gmXg3nYR5oiIa4BvTTGYchA9Ta4B/
l7TirvmyVCZjip8LxrFBzDY/4nVs285HX5eDUdaaIN5oxndhRJYZ+NRgJVxzsVVQ
gSOiYAAIM/zxfNpP6RXK40L3Q8lkS+K4A1umbS08gTdqm9MdoMGhOV0m/ZXxYzsf
euzpNNgQTNDB1kt2BlL5oTZv4vWUqZGb4xO2UZQjlZTmp84uJSvJPCYA3zsbpTIE
tu4FmBQaQHsaXmGg7x6vNkhawa4rKOAMtky2C72RL2aAc6lejIptMsQA91VqFDpk
dQRq985li4AHfy9Vqy6xBMD1cCbAmDQgI2VBYtlT7WXzZElAyQP6/GhXKmI5fUc1
ps8Y8YL9EupKLFXJJljutUwK2/FfDQvU6wiLVelEJ2IPf++PUPCAYFcGk7AkyzGm
cKzaQXGKGBpcKxk3u/s7N7ujufT+12bnsoL+J5WjfVoPtwIwp1OOuLBmFSPtnwSF
y4oG9I4oLQSP+OwvSHwemiLxD8VhtILnZrVMeSbmK4dKHnyDNNihes+twhKMsn2u
9vjKUwVHlFYNwa1T/TuSYQmXGGepXLMIDvjumGiVKRO74SHJc6BN8bkChj62v7oz
edWabMwuABfbkRkFspdCQpn06rqWPK1NSTCiqBQ+X2IavEFtiwTI7nQXtHsQMmdB
gbmlj6PqXlYkFpb4CViU5zMcdvdglQVhO7SE3Lou1fy+ptJ8u+HyHcDe7TxasIhY
SIwI4TKg2KVDFFed5MLh6FcixmMRJ0hcuwcFQPR3hrG10rb5X41MI/KdpNW2CoVs
uLIIZA4zXYu9mlavXjPqRNUrhPL6u4lGYtt6syPI1WiyJjVj8RHou5odN8l5pgrm
ruBauoRTdHvZlGe06Ll7ByCvPakUWO4O6kY1WoVT1JNOSChkIUEkPI+p7W4lba0d
jlSBvwS4Z7Urfcv5hr+21rNpbWCJZH7gqelj4vGDB0PrezRDJpPMTuPOuh6pogHP
tLXZNRsE9wvyTClKOkauOlBI9llRJj9CquisMSVHHOfdUf4SSkjMJOxvKWOnry9f
P6eRwAtROVpdb0v7+BcTXhHsi+/qUBoFZRjYkQS9dHBzPevzNLLQDOvM4ENCUmYC
zk+55wMKsrVfct2OrtNUFdAN5PS0w8XajLzkaOK1b2n8TpWET6Afmnj6Zkgp2Wfq
dPBezSTUT2AnVmQMtXExbRB+zlBME7O757gnxTGgx7WiwSns9WwhIJO687HFAG+b
lT4Ru9jhPESKzEz9rfQodrsSA5G8Qh8kLmRbfb3LmKYqSnS/Q/MVDENlfezHeMlv
c7u0Z2d8uCt7hQHv/9DjSHKJ2nQvWFfjKgjUxA2WV3sLXV63k599545z3tlE+cjE
NuklID3nu5XGeZDJsG1iFK1WQ7XgBsmYMrtZ8W4JRS1CiLJEW3mQIc2Doz06jY4J
whCI1bsEWDJ256zELLLbZZgLztqhy2T2/Eqhjw04kiq+oCEMuaTEillAU3JJx/mm
Hy5nT1oeH89Or4eIOIYL4D1L4e2MxVu4pCwSwA+eJDxkJdy74hNxlCGFYDvEj7t8
WjdqdWl9TfBmjQXzVJQRy/gUBnH6eWdGMoc0uC1bkczDxwHQ3PUCrys8Wm9oqG29
Ywo0md53LBnFAvaZiTppGvL3OGr4+d35qUCgtdSWRCmc5fCMhOsRcuNxBMuro4Ub
wS4B+jQr5HzOcX8YtvZ9mD7rdpaK9C1GoYZLkVs2wtFNjKDG0SQL7m0DB6cpUiMW
wwvm2FppLQEXvjvIh2i/tkVj+bTxSy0aDU/iHxeTzydq5YkvoLmqIOVBe5me2DZp
1rouXfyso94HXBPpTEWd2Wg8BV5nT7SJUxRkFpD59H3PZHqWO7l6QB3zR/8M9WBL
G2fC9gdFM71AlJDAuOlVuAFvjNB5DRGK/tsITSIBkq5ZeZKbMgJHFZ5Ooc9jM1gt
8a/O0RRaRhmEKv2jAm5TjkdY/sjn9BunJfNCkeLulgRGM/yFxW2+2L8y3QRaxjnK
wEE2n21rfmghzVO3fV9kR14038UqgYPMq1Qdzohe7OD2/buO/t37McWNHbeu1V9g
OsiG/vlWWVy8EJSwUfqSDNi+HbPYVN1mLw2U6EywoFn0X2eqZtjm/goxS64LCode
ryTZZXTH6WRMgEEGLeNSPE7Ylo2TvTNQTU5zpyHjpyYLPgRz4Z5aSworYfCALwOb
EEL25XGnnxGB+9DQ900VQdfoVXZvZWMoTJzhjwPUnqLZkXqR04WpPEOPw0ENd3LC
c4lGWm6QRzLpMt5X3xpTt2E28J7oWYPszONNqoKpE51cd5Spymt4B6KDtzWTaOgr
IFoRG8UIzfemg38hgON0aQ9D37+ZWiEFoFKsWWEdnjlEds5Yzu6HMAI/bDD6Wi6y
gLhgkdEIjVXvFOsu36bl7/oEf9WrupxKtM6vHpXpF5zODR1LIA4ZQaFGD69Xsed8
ugdgRj6l406yD9WxnJuhyqBjMgaQKYtJUmVczd88khIneqAyeWWn/TIGj5gteO84
pRSBkeY890DKP85aRNCIsi/Bg5UOhNniVpMKqXWwO0I8irtkpV1rEQDL0xRfxTgZ
pGLcx3wVQMyax0L9CGUx4AdyMesjxv5WQTtPMsrISUzpNgx7fS6AKeFKUPq1NKmE
LzvhqIAGPNz1+ujaFJdmNrzsouX6/CQ8HUFcqAvNGNLK/5PRcJqPvXc7p3+7sI6j
0kFKwNfPsUwKGmpePnLvPegf5BsmHGV/DzkGYuPBZZ3eXYKjL2GL3MJoO/hFr0Eg
VQIFNjThFXP7nW1Q8aaFu8fMUkxC7A4ssxqO6vYxq1CRUrxMh5nrJ8skWIXXBhvo
p0cy6Mcen05oZ6gPdU75tx4dXJcc8YFCdp2SwJ+x81Uj1zc6OY/aHn6fdduelSJr
ep49KaKKyF0fx5Q95mipURSYITVIrAWmzEZ1/o+n+GK7W3ZlqQYEJ0dQH6hxjj5b
X/js/lCpSsbyMmFUrn3bum0GLr3vggni9qp/bkfXFhfnzwCYROHKYWFm7Z3rA6DP
gjTfW5Ne67vTL3hnS14fM8nGVkp214We+UqtYcOpqG5dPGssszgUHJTrDp6hllO+
0vrJU3c5BO0zMHeKg4Q0GFdY+2SqgBj+jTmxEPc6HbWYywECuQG50r3YYRMdl8+e
OLxaviDDWGW9TDkaSlwQek2bEGMoQiwpyh+00F8YWikXolfWOQI4b4xZ61TPmDYr
nagJkxHkcuCEFmmxOurelDP/+IeIB+vDFaVIe+DngEDKzaUZnne6dsqXBzGC6amK
HUZJdt+wtjEDWFhy8/bNvZnOPg14cYhoDixdQsvH2NR/y83ByJXCcIG7nnj509br
uLP3EijVt05MWqjbHOdxTMP04jAoIQV0GTuuus3+h3ua9eF0HxJdt99/uZaZo4sH
Ffl009+25UWaXhxz2sOJV+dnvl8yOi7wQc3LcGc+6kDYB6G8goizrjdvOfsn1ZK3
+PKhtnm+3lwpwK4lNb7mUni6LXidD6lEDq+zCCUBxUhUHFl2aBKdm2TcN3wraHQ5
BhkxoM3bqHS3OtomdhdYpQNFB6Yzl7F62l2bm7sJl1l8srErQvR5SBGsQ0pzBR+T
4BqpUeu0iFyCgBgxDhbir7TJYb2sR0fjm6V2RiSxm6AYo/gkYSaAT+W/D9CZhVI0
loZukwjcOQTu86LfSpWp7+2ps8EJGlx6TvyHquzEM/41NOymnlSdpSUeXD7ypAex
RUJRPawdRMQ+toeNRnZkK4ncTbscHQ24eSbvjTZEDLXlUMFmI/qqS/ydULbls9yd
oxgMAhDkwl8yShw7cUfUhvlUW+XfgchRiqxSVoLTwVNiLgnWr1zNxQnij3HcLyCo
X0x4dJNqYBQSniwq09dCjlC3IVB3UkF0uA47kh5qwCRZo8FU/lVt1p7TgHLo2Gl2
XlD8SpDtEy5VRQLjvSzRaGXcZfbgWfhaPxS9kO6ips8DoSWSG1pg5vRT6MMrSqv4
fwSCXcAyCbDtytsL1h5TcIs4zXra+dyIBHes+vBZ/906DJNt5OQK1SM1NkksbTu8
iLuw1fG5CbCst5uVZFZpa1wZE5EbJTX4X/Y2AcaDJ9v+QBcwB3KvaZuBfcptQdcO
ZKEbPY1Lo1f9Z3Sj9kr3RysWAALJ9uS71f/VtCY8yQCUBEGOJgxB0GymvlPWvqjc
D+XPXX6m1r8UN0Rx7BkiIppsVy73f4/5ulbaWJ6svgF4M2KvTJgECdJH8ljvKfnn
LRhk9m58+fYWLIhTWy/312h0WgpIIpHJvIyUJOVkhoK3bo+kAgJVpzYKqXON6VRA
tf8fqK4/7lO2SaJvm4P9D5Gs6/32sC9YkfHcap+KD6jL6X7Mz8q6g7+HG1ZHrvfS
uGBF6tLAnnKhFgDOUi/N8sct7zjy043oDgjo0T2MB20HLIeQO+5eLRUPTJ6ibQbq
GltD2j6Gsq7B2oj2Tj451WP3RjQBfB2QCgdkAJddenymA3VPWxtlP18lpEHTIXQL
bCioiwdvXziJfcWr4dbzrKs4t7WFl+1JokPkN+BLqwMs386aIfU7/VjPTFRTxIUs
NfecPnbmNe/HfQ1yzL9jJCUptCataCAKbG2GhE/0X/ssd8ZfCLnchJJsXsShG2yG
ckPIpAApXjzUbrOPdaJaHYbCzvfpKemd44ndSYMkTX/DWTSwVde4rM0BqC8KX8xg
tm4QWVel+JaghaA0c6VnmEs0noGHubeGH8osgkcYrJKpdACh77Th0/I2beoQRz53
TE27VSyGi4yLJr3OrmYMLKx0G3MdY7H4PwKDiORZG1KxxG/NyhmIeguqCiTfdcMr
wG1K1qlr8PrfvuynIASpl5aZ9ZxH8nLR6+g5TGQC4p6PYdeCUQBcN4hrPXQZsdIz
AGZ88VrE+XgB9ia1ridygZg0OUD98DDLVA1N1TEriwiZbp1rqyBP2ksbkIYrPDPU
r2Yh+5mEigXV9mjpGuKDr+1yTFRXUHy8FdlXByMCQDGgCj0Z9TTZLY9AJEJwYVsA
/tpNEYxOIooxWAxh9ihSniksAsYx3iT87Z+aMB1CfBc4XiG8CWxOFEyP+4rul3sZ
xqX6VSDQJL1QikY1N53KZ14zXwXRM1+4dS6/t4WXUSxpSgFSdvAmV647UrqONahx
kgioFzdedpWjiBC9J/3iriRhuthpvsYC6b+bY8dR1Lp5G65jmImpTWgOdDLA0zE5
65q/3DDp8uG24bbbjHGa2HWftOFx4COESxTkaktXQewTKfpkeIrz+GeJF+A6HkaJ
XKhCEnogzICYph6DD3KvRF4W+vDb/a11Nwfz6EmgQ++rnnmA+dG86/EsVs3uX243
iZL02RZyxQEH8w67WXATDxxE/rehLucTWRAvNHFa0eHsmz+j6gpzw/mc3dUZLzAZ
4dgDnLGKPvqgxMiKlaQT7E/tu1AtAwAXaBIk0xpMlmc/mpf5s3+wW9yO/beaW8wo
cjMiKNMUEfYjqu4+9yE27xSEWi6NgyX5YztnOYMZvil5kcngqi/hIYTMDeVQB/ry
zTNyb/vTQAgunUuwayc36HuDqTu4EfJ7PHNF2HkQR0DplBjCWqFAXCcIyF/F+A6L
fnocNW/oYXNImm8K0rizBSao/utFlLOT2fOLdIvHev6fB6IdezFsnLG5wsUNeVaD
w2G7xWFfQj11dEGSFtNwrbc9I+k6s8LymmSf77xKRRf1xKZLlpRtiZMQQW6VkRFt
T78yb4Et3RVB1C2ckCCpCsxfNyvNQJPVulEXDfbSDo/hDFzCOTvpJRRLCkPv10pQ
48Id0gCgkXxkzp/s+cGoqhQJ1GfEcenXLk4IbixiLMD0k5qw/Fi5Fcuc7w5bPHY5
gPHPixIsajhEvJo7z9v8UMfmEoQIktbdd5kSlqCbWSjdEHsSgdmjdkZuw6UrvLBG
kmII4u0WIuxD9ob8ucfL8PujYN5oJLiLYx4YfORgxD33FfkWphqhn+UTYxyiAkKB
F9C9dn+2RqWvi17weWAxE4NBXkgE2DhMcTrJEnV1HnMqh7g9pTytZtA9RQ7/JVqx
zqADPNSc67n3JBJik+zgvYYoGd6UhYW0p1nMtIiureqCgM9OWzs3+0sW/rHPRdxk
exx+Tszzu8pFp7oTGxh3uh0ow90qOiqJE12T65T964WJ33hXTiHu+03DKXtxoALo
os9RgqxnPjDIWXjFBNdbt9fgisPdFuQvgTe//i+D4m1AhC+ZLfi4dLRFX5aEKR4V
Km/AA5tvDh8fJft+v/psejjdO57FUsZKepsjtCE6aEMaGTRnHFUA/zObtMfQV1pv
I+UAPdAqoDYkzbGCk9oJxyR0Eey0MqGAiRrYrBbj00jmcAem16B6gMhsi/jSf2aI
kbTtXgBzYOXcEjQkXulSQzB0ngqlY93F8BgLqh4APHjrKBCmM8Oqavh9QzRp1q79
ElIYXwkt5tuQitdY3EEjLD39tLWw0sy2l4ugPAwd6LZc+lFX4mT16jT9NL7lH0ig
aGFiuvjNvExszPGQwh4bVUL42P6YOVk6zImkGCZWORu6dFNCaN1vcuMPZd8Uisg+
HLjKtqnayoqR08Oc1O7iv6EcUUwL4zNckAxY9MOcXpnd3Robd8MES+pGyyMDFNT3
Qc78tOP9F84PJGL+rh1I5ua/OJKrDQlQbjhG961E2VHqp8xaGQezKekTjrEEy6Th
D3U6r9Zh30xMW6ZlzN3CZJBGswuT3MfkPWE6hm/cCVbW5UWfbQv5dTnTpTQtRrUj
knRDV7FPnAA/PRag77MosG7Gdp5ZYfG35l7Snj5ENmAFbTiJ3QAtOSDh+Y8/lmF2
Qu8uOVxvBgLCAMzVFYh9EmCFeyyAZe+OKPZ5522Cj4kT59QLPb3Y5scZyIJ2wVc3
nWX8zNBdqzdeUIcLy38DgKD/VEtqQbS1ZrfY2u/csi4HckoMtRTPwgK028JCIDpr
pOuhxrG0O/5DW8o7cj3K1pqNILYJBY2Z5HS4CxOm0rTOByxdoEdb5yxHTCyQBXTR
T35RWBPGPT9P9S/dAgRWUSdcUrAPvcda2/QkM9NTmUiG1uB/BSd5bpQjyc/XPVSU
WBBY7KBWi8qhZMbGBNo0w+qd92kwuk/+nU6/dPIkGkEuGsoqTu7X5bUNGDosszZD
X3AOKuMoZwwP+6VKjEmT4TkVXd+FmvhH1yttFvJ9YWj3j8IWihgy/+LLLbBc20DD
LDJm2i56ydK9ps4d29dJCEoYGNoHvJyKl36Tz4sYrv3miBj4210wA92ip+HIbDUn
lawu7gctnMw6ttsa0vPfxhxiWqTghfBijc8k/yVunJNIqyjEDiLrN9OGnb3cQm3c
wxUbsOkl6OWO5G6f96OFSQSt0mIyvqrOtkdngJ99q78r6h4XGGw1WyFOlI0xpMJF
rNf/NyHWMa82GZWRodG2gVDbMCQnTFB3dL/e8SPM2rtbe4KkHFxRnBUZXuvCXj5/
fIbVCSejOQjyXVgbFP9iwCMSVd3IL/iw1trm2DHE/fjaWmJumTmibY7IJ1KVqjDm
vWAnL4mKsaOhwLB6kvSnbXnoL5QdWtFGq4UIVoBUP75bTKl+ftmgCaMibzeAUETs
jVeJ0W6GkX31DMJWbnVnPtVHNdgOckiqSXGw7eLl634CayJXEMqXvHW/R4GSlal5
p5+Q3DFwP9iX2M4tIjMxz8lXoHFwvCfIT7NS8msySMv6TzLxuvA9osFdpib2aNbJ
brkgZQ/Vl+89GS3OMQxHKfN4mnG5GA/kHoTgLHkXU/nzfcEO3Hp2hkd4cOe+J5MU
MTwwCluKSZIbVqRNpikpROwxr6+q9g5VV+TTjM++QaY9EJNTrYk8zDXZZ4QbuZEo
2x7cZmZoBeVnxHUZlzSJuJ1UytCVKYHXblR6YsqooJ8B5XF7JYmPg1h4qgMI7Aie
iFO30bBGvvLd/tyXVCZ7xoAMjsdIvAl/sq13qfdMAaK8jkbWYGu7YsqNnYbjVa0X
VbHdDgWGWcmCnBj71dmYa6qQ1FYPxAG18LDNM473Ic5g7dL8Te+XlJbsOInh8lyh
rdUV9Lp5LNUmjTxnjNV3TAm9ur5Px1nt/zv5DoornUxB/4reQkQ8jAQACBcOekAB
Z9vW4QbAIXk3veQ89R0AA29GfnWFQSQ2CUMT8oygUSudk4mKIFL6+Ta7hosDQ4SP
V4fJBIrl1tDc1SSvCkYfxd0nwiMQyGvPJ5WasF6v9z7sPZp4kWFt3bFnV488LASr
ZSpJQdh4HXlOo3g5BUxkdwpGkrGqMvFpnVvTdhfwILsq+7udAvjMRewF7Krluy6+
jlCuKI1doBNoZvXTITKcdxITOj5iq82NqUt0Sz5el7ztneSQ7mx0Sf/lAPvM80Lu
b39HFZ1WpNgrcvi6Y3k/IMQEOdcV3D9UMdiV/7Tmnnd3C9Jk2/tVWAsZw7620Idq
sUvBvhsScyGJc3+RNHQyxdM29YB4Gj1KUujl6iVeAMAXBI0wdGXhuM6IpKjb8YGK
PWSencUlTDkZpN9O5JnTM7Ai+Hw70nMelBiX1T93uOV5AZLvfjJzfGos5Boq06iS
jTyPUGLOhDo6P9ADWh9focavOGZ/cdfeLWEwlGmPs/aT53DD/5rPY72jB+6fToUK
zQjIgvF0dpIGqW9QlwBOQgz53J5nDF3mTAIQxQUuy4q+brp2pO+MMC1lBZG5qasV
nNWBxk53lytR2QcYt1uRX0QOwICMm7N8V/aFDHQ8BGjA05BwEl+2+ISm9DEmzUnK
15xjXpKwGZQlI0uAqXTShaAmLLnZGjLz1aatT3WvlDVtS8NkVb5Ac1p7OMmTJz+G
3PJEh1PvT1nQLD2dMA7/WvvCehOcr2fs1AM0HLKlB4lpWTxCoIMkewi7ndTkrEjP
v90ZIhR+N2nHKYf2zEj/Bz6rEj+09q1DUHYR4E18YYZvOT1hh5pkJsdQajwP1yrx
QT0HDMvFNTaZR9hzhs3zSqzNzwtEALhyXOjBRij4Kc/P+9qKXqfWnOpg9DIkKlaS
qb7JcqN+kV+hKi+aANp6TqheOhZu3AfkTqNQpSrYAyhr3yln56HKdtsHduuInYc+
LqLhMbKNkbG4+++lGb9fEa/HonIgXjuwQhUpqPp85O49nHMRV8kiwS4itV3FM3Dx
kjdvHYUAat2qX3gqTYozuovTdo0hywHVx/3pJ0pJ/OiyPOuIOUOG3n6SCcq78FqH
h1UntVmm8fdyfKJHHDWtVu5Yd4p5tNRJ90q8A4RHgeV/89NOZqyINdJ9qRlYEHh5
UmYpEG120VG9OFyDsUr0c+P77DA3Zo/luLmN4mnD90XuXSSa/j1sfS6smrKbOiRO
lwPwPgeYUYUDanxg7APaFxos9DTjXQCY0Q/FlOTa15WL5qNXUSTWXFkrb4M9JRkA
T9c8UBidpFZzzJm2OcAOeFd4NpiA7xRUGSYph8sTxatECzYA9F8Cceeaj64e936G
c2QhpjuwuxdH/eixXFHFNSaNGRsM8XAL1AkMU4bSVeXu/9zXQabDFgSB59WTfkfN
5O2NHm21enj/QTT0VPrOQnektxuHpgcKaorybIduXk3SlC/3R+kGSCQEvmc6I60j
jZqFsiqWtFIhfC+tDbJPB5t7fd/IMcEcIVzNQrydohGnRDTPbzyA27a3g3M9NeU7
O177LFe3eGJThLCsUOXCqLMvxO/zSh2cVUq5PgzibvkG6B3b4h6e7FHprEpE9+w7
bN1q6N2DS+Q1lEPLf6TDl8XxiymuBVCozcLs2r5oYtL7PNAxA3xsnB+hsHv3zhCe
8Zx7kTkGtWJLxFDU5HVhaDwWtFEp6nTg8/fSBC3L6qYOycms7pJljXJOmVSqbSuE
jpWQtiVJOvaPFW2aSYo6UikQHWvEbV/nNAg+8U8LsyBY1xA/UmOXYSMAt50UKWJo
P+h/UcI7dmLMsDfAHaki0nNWKcvh4SikznJDW3x+cMhzqQNomFyzzEza3SuTalFx
BgCnXfMqwvOxj4BCZS5udyRiZ0jVZdql1OQRryQQfYU3zkzTMD51vT0ensYzDzbm
fr9NLVs+I/B1cyR+bFJ4ieCSkPq5eL8IwDVQot90TDLyye9UcZYwRJokTrm+anY1
lLnp4fnvWbBiYv+K+lHfJzdt7Jf+Sdk/hpU/OH82Q8SJRmWJf+e93fIUCTrT90Jr
PpHiJ6iogku/2MrCoOXrM311FfR++3kvBjlPZxsed26DLXfDWihyL5OHwMfGO5Qu
7JD8Ife8PNZWHr9JYXBYznO9iA1TmJtrMZJq9Uacw/UNvUwr5dEQoxMDdzNFsLZy
GasmtzdwuQSjURrQ/0JidM0x3wc/r7nao2nWzDccLRxZWEzinAx+A9sHldNDj3GS
gW157ao0q+MzALZkmDoFMHkF9NGH/6NCKekIFB7SnAKkohd93oIEWagjNAh+HZwl
LrCqeeKboqsRpW+6b/w1RDxO0PZoM40lMlmQuZDiMvisT2KOGgVB8pWwq3HCpGVY
+vQJ4Oqzy/MNOtS9pdVfw5/+BmAzOM9PYToVGAwzCnatbjNcDYC72IEoTJhZzSdJ
XgkPySBGgr2AmvBRjpQXWIsj9yXnCvtyI6f80/ntv22mAQ1tpGoTpAIAO42zlyWW
6pKT/nVp2TyxWlMduID7VkmOa9zY4BxnrC+CWt+qwiZwG8LFnbbhI72apMnwkqQy
fC7YS7IJS2L3qfpuTsXJJZLy3NoABMOwH3c52fUpN55oKc0n2OjxH3GC+rJLE0Vr
Y9PHk/D4bpphT7Mz+h5HGOwroIlYqQW6otpLliUKznrjHNCt4GcWPTyBCGC1UmN4
i4HyDsi+g74aHaSZ3OAsTNRuDsUzSDKzclBsO0GPSBbsayBOWmtqrNBk0jyUaFe6
aPXCkqPtETsNQlpV4S75dXVXP9/PukKEXV/VHKIxX7GgXL+9cbrguYtn19VS0aH2
/bgB8lDJUMDHY4BOBvwEjddSwbS/+eB3X+HTrtJ0YOycLqkf3biiPN5ANZoBhe9m
Rfrm6w8vvKdeJzSH3LkJ+1yrPxdFzrV29C2e19k6VQECrnxu+uDzt62BRp9mnNNx
dZ6Dj0R6DYcweI13SnAJXwVo6WohnR/tySXj01tpzQhaM5NhsyU/YdcLuikgsrD6
R4ZB6te6ah6ThKAwU2sA0Rovd9uKeBMpPwPvkC2h6CHMrZnO8ucaSudbgsSl0LJc
03fJDlbkuabqkFG3vb0CNTd3cvqm50Kz2Pf4rNgerJFWK+yyVjlY8I2Mcc5juZZJ
x8F6zTrJy34rSO+UzJlrb2yTOOgFRvN3Vi9Bi9ujHQViIfffOGtOzJpqovUgeG+S
4ld8eOvsInG3VCEIsTgBvHvMOP8b99wzVWtW3g+xn49Im09KwuvX3hkrAYemXVc6
0ighp5rI72xUGwjCSYdsIS7fkZo5En0Zhyp3Hbqd4Czp0awpyEbM76PCB9MO62Y4
1DMlNpDwQrfLSYC02GK40WYrwNO7JPqi+RyURzkEeNH+Z7Ad3qXiUQYYIhGV/V3R
aNgs6ze7tIDLoq1+gq52fgT6F2VSqatSvJnFUeuavw9CCOWsZsXXpzvpcico4Rue
k2TrJxNGkIiz2YlWHActcJElEbgwEKjO9PM+kPC/a13/Xcg5tEHc0JvkgMFz9Ia8
StjBSR8tQ4FFxCyMkVeZHAGfIisTeKINIQ8hG37lA5UZW8o1C24hnUezMWonMCIo
WbFrDZnLAp3qB6d0CwvhgZekOyVBGMogmF4QyBTvBhGHu5O5GeQMzo0h0doCePkf
FX0HCmc9j0AHxMbWkhzYCl+NA+zwrDaiyjl+4KlvyMXXQ4bLTCb2eFfcMxXJVBhA
H74mDRkwSNbPp31aniqvT0SVkDeSpBwoTZ39aMfEsBEjNjx2kRJrOus+uqMdZ2XS
/3g3HQWTf1IDstJQezSB3H0y3WmH12F2aeJ7/sqYQijeMwACDENucPUB06NLWOnp
QMWHAsQKAyr/5w0vDlLmJAh1qYGU4uAP8d6RX6ltfcZVpTgS4CCdvO5kuSaFtD5+
jlr6XRTKLjkUEY35D6EtJYIOuy5Ph1up5WsSaxGnyp6Q1k/jX517p9MqVpUraixD
Fnolc3M82BOmC/MbhYm26RsQyRhakHPcXNWQrPM7AABP8AvD3Zkl3VfT5scLl++p
MKaj6BQXjvMiG8NJsqZ6in+C3BLHjo6JqECbN2UjJ2qTCZ9l9I+QCBRE049h7na/
GnBN4EKOOWJc0XkCE9VutfiTFF0EgdI7Drd1yiYfiweFufxrqyJjv3P5oNWqcQGm
ObtWNoHTDRjnf46pdwxLetAArZAgE37Ij6XNrrlazb+VpdjVo123jX/Qlc+1wYNx
xA8Nxi++WDtCfqxOpEG7vR2VmMoZ0xwbpSisoqGUj99NWWEfUyD377JfnPNTr25o
qLTQa1TEYGYCun70f5erS1GEL+K3TYPm0cOsERjmOyxPf0vMwJO7vnjMXFUfzmBM
Dq4P2DoSh6CA4z4HFHDu9qXlAVstHUElzYw2Oog94F6A7XGDCQZlHTjOkle5qDKy
zLsS13C2fx5Xqmay8/RcdyvdF0YB3tT1Npc39SEu0V6lM4kmhXqOJ1gmBhJGozhJ
aPOk9HynbTZXx7Vdt8hX62UbjIYaX8KqL7pRpUr2i90VoiEEFLzZ9glxnRbhMCvW
Tn8Xpm6JBf0Eaq5RGdZcIuUyXel2cDjfC4EmaLjhzXOLRsZGLKqzZytdkrMVfeqF
NJHfSg07UtL8vf5EhDhzJlkEzR7z/EfDPo3yKOsMAK0d9B8e+AVS6m1Xmh1cU9S9
DpwzlU+0k480uh6jqSEPy4zghttM3BjxDzLAF5c+e8Mug7XT35WbOW2vqdWSXpYM
2ilXsBvOmjwc2Csi08WjLQw3KVoJ11W8P/vO+oE71QuyAWF96jDHnsvWdSsVbxHt
KglTZGnw3J82xNEasYg/ZHnHIaJJ4pjKdMTVyespI/WZ+47Cq93/b4Rzj+Oe0E8X
MVSngsT/+hoTGHqECx1eA2zeROlkpbCzOua9PblH0WM7W+k44VWTW+SMLPI5imfl
mRw2nsdRNBiZVDKggIAR/Z/f3BFU4k1GbxJ6AxSh3G9UPrw74lugPGOmJ8J8mO4h
LqVf88c3BuEctFuxeIaoT/daXCHIQZ0wM5qwcT5PLaf7NSdTf105PyJ3yzvVAT7U
RqM8LNL++gZbwNuS/6Oqnkq8NgNqHCqTDS3VMS2CBmFUOxBY1wSldx51ioUfT+aG
4ZBk8fU3g4W67VH4bKqXHHVgeJlZm9wzjUUewLvkL7Dh9YlWiRv5fkttN1qkDD/9
16RYyESxTaCY72lPME3WsiJL3+k4w4XWWUTvjQiHDkrTZZuvc+fRrND0nL7b7TdO
VTnC09jP/DDBcACWr75/n+EQBsqwltFIQNg49fg6fbV+tovILy9Ium6bYyBmDYjw
g2Y90IjiGQsGW7Gj7o3otL9o9GLY5lIAUCx9XX0Kjfj4N6obgusng7De7YkbO6PR
Cgjmo9KKJh3LPr7olCl54lS/87Y0xwLJRt1dI9twnWbIUsfdzzyLGD2wnD7wJ7Jn
IvBhVG+FYjcELSsdMjcq49TJMeygL3esNnvscxuj7uYLiKknLBnfGZVi93h9bAQP
YudED7NcaNro8iZvpMuxGIXgiJ8pbyOyNsJhZIMKKTH9zFA4ZiV1ADaQARv2JEaz
EOpvkMGRF1o64dmzwocMFuhf+UdoO2YSQIi5G1Z5HjOTqKqxdicFav4kNBWqWrby
wNVI4NHaryHzm56Q7QNl2N5a4oB24DYXX8NxoYZjwcxINZP/ezwHCCVj05oluX2X
JOrfS80OYYY5jRctWzHz5FW3rA8ybI3twufcwGNTquiIpEsqTmryNJZGxkphf3jn
D2p89MIPdOg9yhbTg2rYgXTj+ZJmB/O4toitPrzh4U4gF0tAK1DOuxa+PTXSwAgv
icMnBbt5NXtFCJYxAPhO6HEB8do6af+FojaiRjEgCbtbtvBmrER/6FLKUDbMFpUz
Y9tTmFGFiZOXaxUQJtoRYybkJajHz5T+eDnEOuyGF/k0armugyyJXtbGlgbq0HkD
u0LMxWUCbyQvwZneNQRVkcnWkyVvqG+rrbLFbRObxQGX+Ru/vt87OWeZrMAj1hmy
DLuS+Qlf77ACCGbbayK7TEjgmPIuWuiyFaRaiCVchctbXJ4RLFyBOB82yv01CRGA
Ne1YHsBmWeejEGDJTptvzn3piRO5+k/V0iLUao52QKad/e6+0e90OgJKqcWJ9Yti
k/iGVGIwBsTxkSK7gfgJDMs8rDFLmwxbrYW5BQu3k4BngJVQe1MNqa027j+YcKQk
zF6L1mX4CW7m81RjHspTvCG+qnbtr7eJVzeX4AgDdRyhYQ7weBG0Ukx08JabGTV9
I2LaFaQbyt6YiJZKGFq20k7VGpEjw9lelj+gBssFVegJ4CAKZEACHZwlUDgq5E1O
LmbRM3vlBMb+VkU6e4gKzeQqXQ8lNGIDNGFYFj5Xp3bYaM3cfem0joRubyjUKYaU
/y2OKjGf1oSJ23w45yWPABzLsX+DWKiHGtJYTGSjWtStwEBc4gThDWz8KOwahEh5
E74lQXNwT3eae7kzw20L5QGYG1b1xfTm/IRXxRItu87dbOo244KQLuTil9BGsC6P
JOT0XBdBIZ7NqsyCTFbcrQS1URgEKb8ulrdgC3S8tuemY6jLukIu4U+x2KiVlkam
9a2vaNyXaPaNNAyLJpHIL73/0TU0bsb5xtMVsnlab7mQqY96Pqkw59WJHOKOWk6l
q1MhWezOL/7JSpa2bB9hOMOEqK0gwNjrapTrt2Av+ni/+efnBQL4EpgYl0cu7qnm
2phb26IRBchRFfTnC0C5lrq+DNJFsc/o+EV+HzR7/0mUJ/LKLog78aZFB6pjcOiH
qUjRiNgn6djKPR6O6R4j6zx20wNK5s1SUDkOChTBLzq+LExJz1KF8WMRTqIHZcVX
x20mSUEY0ihE3usXJSvF5t/5bkrTvs1DROneQXIApeRQvEe2aXmj9y8mMQSRKakL
RVuEwK+PchcoD6RgeSEncdddXOgduXvFrEQIkuQZcM+0PoxYvdTpZfpEU6sOIfsw
FiW8oeXR+hw2gs6sHM8yjVcfzWHtOFBVK4tzx7XzAoF+BJ1/EfpD2P4BBssNU3Cz
KEilMnakT/1o1ooMsWXDAojMMBrTT8FPfJjFyBz57F5TIjjhvmfPFcRNaAxhq+/v
x4VEeMuX8xpOE2fO7JTYYIEkbmadCY5jpo9/8ChCDZOxn/K0KUeC90o4UjhPqUXT
W0obGG5kH3cWg68Q/GFy7fvw4utXqL6DawctimuKUd265kSQ3Q31yWfSe0YD6xPp
CRGKswol8/CGjJKGOksH9tSevycKgQyahuY11fkFmAfg8C6mxi8lWMbDmiJhKylz
mXN7M6ahY8pmn8JKP8sdRf/jQsaLni+eMKi3Ic6Uar76muYtnWHNz6jgAZVVxDQG
/tELBKtRyGYaQsfZjSTVZu7RUtmv45r4CrMHpfZ+YTgDaFKpv5JQ7lcMb9DbP2LW
pssKZqlTM7/SztziANLzvUeTyLLd1TNfZLbTJ6B+Cj+3O68geuzKizh5w2aqvA/A
YxCV1Nn59u9LmkStGfNWs2HZ4b55J6/BnKL3PC3BV7KhIZP4k3o0gS3iFAGaIU2q
rNlW6fWDWD6ICqYEfhxaEs3IP3okgrRbM+G02SeU6y+atkO518JgLI0sO/YVXXCh
wCq9I75jXIWVtjMaIUC+AEHOsasbyArfSUjL+cf+RPazOmgLNYTtQeYOJM3soRFa
I7oy5C5sfA5yr24+jLcWykM+KvqcKr+ewky8cddAp4LwhEuMvYNH9YKXd++Jqvw7
koEUpFD87Z6D603Nwet5ahLZaqs57ihcUwhq1i1dR8bu+cNvFQAvL2vEW5+zawQz
mNQVz5uAmkM2J7ZIoUxUA0rvXps+vShY0ykuwKFPjA634Yp1NeIGUVlR11rljO8A
IlJLn3XBhy+4pgKWZl9Epc1L9GJZbzuSFGrnnaQwa7nVL348676Xa6MGJdhM7ue2
WPEBbXb1+p3+T+8rmdjzotS8WPtpg81koyhIEYM0d2JaXHX8Fo5wSoeLZPWhDV3X
E+8WK2mqMJmYO94iYSE5HkeFPE2N43oYU5pE1NAPpfPQp2qIFp9i1ILFC20fP/aC
joPtiOjg7umRnM/oRU+7eJRtmHLyqj3V/Sa2Ab7LzXBpq3wpyoSBZN2oLq5UEoWY
M2oG/OamwhY6zr8RBReFO67HCuTjLi1U9znhMVmroAOTaA6h60fX96w9aYeN+mSe
+B0L6yXaOpaYqI42lk6xaV2HZKHz4SrFPpPFk0+VLwA0yiYl+mCSaYkSS6qAdJ2g
n1VrP0tDmQlUjy2vf4V4nAxA+4GeNBKTGdNPMbLblrUpkLIG+K2ccbzi9FSzIVjY
CYXN48dP2bu2QP4/bwmYrNXgMQFfGLUxkl9dblLpsX324ldDRUG4JjWs5nHFb1/c
zMlOfqflkPvgHJNnmaGvz6Fg/Q++k+dJ7wKAydzTBI90lvkx6SjV1NfyX2k9eK0B
oHCjyhVzjSGgxiYkD+sS0KxW1GnNOUOYNAgpfZPRhHlAHtdHF+0WK+fkXhIRXTrz
B2fsxBLtmLTV/E471kQaxMWHt/6s1jrFFT8eQhyAgFf/zpqHleCVcL861YSzoWSE
6aYh69rPRodF9X4R8Tp/RaVbbty1r2v02Zc/oKo14rk40M0Pw1ZZvxBl9ZycCqB9
3HfQ+eQN5NtCe4Uc+Ojc4y+o2+lAc0R2mEcy4oPpKyuUCDWdRYm5aQTCOF/o2DiK
q50yBC5ENFrV5UTv6MG50fCaum8ACzO8QD/RScdeDdzKoLOA9a8zy+6I8aUDD0RJ
40efsUchGAUYRaMmWqWY8TPoPdyMRPaIIRh6qynQzjuKiQoE3wryfZzAeHArAvIt
wqLhGvkVRvIyHwi6XJFcRyoSzFYBYlDFaVN6UnCGsDxPFRxDZ2q10kuqsodTFJsy
sBICLc0VowD3eHX8YiAfs6ycf/8ZcegnRTIWEXdQY8GqeEHkODJ1d26QLnl6Kj4w
1v27QZYXnINYPBdvT8sHwuIMevILktrWe569awo5vi1G5n0U9UWexoy8Mw9i2gf8
UgHZ6NaYnVRrxgBliWNbl67F6QWgToDOYfU1aycYGiASJ0lmJHJQ8KQz9eHzMyzK
9KUWFEc15whlOBeci+h1XkxctOpAbXove1r9fmwR4y/Ki9EKnFsgCVlzRAebBn+q
Pm+0JMLsh92J02bA7BFNJ6a8Q6XMwRYp9C6RSXbOOXl6gJ8EdAH5rEaH8TwGOR4J
ttoH5RPbnQSlJLxcAytF1q1mO31N+MuXK5hV9Q9EOoph3Kby8L4IUwXy6izKTDbk
MdGfYQAtEWwlE+A/x5hfL5Y52YlJDP1rP02PqcqPTOy5sGLn40RAhTATVyOaB4gC
OqV3rSUzCJGFvDIwGwe6m7GO8YI02VlhGoVMapZ1d+Xmuv9/kWM0jwsvGaiMemrK
nyPbc9rVCL1nWkrilsZmNk1njSjKEW8It8HvDE24aMBKoXo7bMTWhKfEmzi96y6Z
DLQ22aJj+9BeuZjS43ppwlX7tiHBjV8364YBor0dMi4QSFNRJq6QSrPnUxADhc1l
AV3/iHGwjTtA51D3CT1kVrbT+RFihS26rquUlGU1ciEIUqZcOpRvsWofTrxxttKm
R40gqvd4+zwh0TJ+vB1yh7CQFh0y/apZY4CezSi93Cv4hD7bbXzoFVR5Isua35le
wreIaXquU8/Vegh3etar8GgmZpoajC7oIIbkcfB5dcaaOiePu2hqEeY7sY0Uj7en
p7VEkBlDXGbOzexyzF7KC+OiL0ybnZcI0DkBxtuZDR/4gImCKUoSlwicKPCUH5ib
TPB+ZlZ6MklA4HKOLXuN//eP/c+r7ajyYWYNxYaAf5O8AOemh+SokzbW60q4LAea
SI7fzW/SQsyskap76mz/Udc5ByFZyae6dJefML9DSDbknGSCXyxB8kPVfxZaD8Bd
s8smdZ1ILViaJJjmnbvV3BM/s48zVwxRigbFolw+oOTF9D0CjjIgUuEB2G0BcRt7
LLEDeNI7kGdRxMDke3vW55r/MV1sDyWeECn8AHvkH1xxWhTBR52WgUWEVkGgfkHK
Dpntpn8o8iEQwjhqFSkhNHfX6YiGxvpNvfVUxnDN8ig22a+NdMC0f++w76CNegMv
WwZKJsE+5s/OM/Tv3Z2m+iT68WXYgDpmEt/PqUgsTGNCmHrnCey+Pz0EUex5L1Ae
Mx8ey6s4Icsbr0A4jvzHX8PHVkS/UC0dno5UhFevvP1WnHb3FjYNIlz7LOk36rEh
OKNbPC5IrtdpxTsEDNspGsKU1Vt4tWMHiASPZSI64r41K6ILxnx79PolVE1qWIs1
8R/4ESmTMOMuabTVpRKiBPUjCJN8DqCUvh4UKgPqx1cnmSSGsEDfZFSKOV0FIF+6
n0BaIJxIOBAqz4GRAOqADrSm980H2bai8BIHhMoNeKMhWK0kjSeXk8Pl9z8fQqMe
xGlt1BFWkXDXZikV7kDte6kOnqTEO55Rbhthi9eHGrJKEH5zVp7tGd62k1+a5a3W
qHowKak1BqN3d8yKuGr0DW6srCHmR8y7nO7SYKYM+7FXB8x4dJNSynsLSbsonQBK
rT7EZAhHsDKw6ZORcW8fFiI0UQja11uqXKmn6hGZnuu9RMx73wD/2AB2R5AdRO3K
9e+J1ZUDE9vtyUul+T/OBthd+lzKLY6VR7+W/bbSkJZChmrpozGvRdzGjPb3gUjD
79txRT6BcMV64TPAbIF4Bbpo3nXPx8KO4Vuv194xY9pCpwTLQGPoyWT0tLjYdVZi
VbM4d2nkpKs9hOgv3Q9tc8pritszSqETG1vL1YNGc4HL5PZTN0AzKdwBBToj7TJ5
I/qA4DmSMV1Rsk+7JWx0N3EyPr0DDr+wNR81NqrWYvJ0VObMoLpAEGUmUT2vHJhI
p4JLCPGceU5s7oeVLdYIBfDmR8wRB1mNJNCdj2H/Etke8EEv65Co21TAx3d/HTL3
P2lzeAXo2b1UBQkkUe3wxcx6eznfvqozzd2XnXalQIhmfPmE6/4NUu/cTfBbKbW6
O+lezVZYAMnQKIxY/XCjfmcwdd3YDrkHo4uWR824ytJdxbwbvG+PHw0Y+1+WJ0dQ
jOO0evtnb6qGuz1HvePmFE96JgfKLOgmhqyu16tWztiF4UJsPu3M1KpbtghbSl7+
zwwZnMqU9NtSLRQxonVljwiwP2LO9So62k/thWHxD+ssC4WaV1YMzpaYp1GtDzop
bVaWAzf0ySp3pJ5fnFRoStYynNao6X4z1Ln7x/onQU9PurcRtPp+BHy8ou1Il9JQ
qrmt+EfvEpdcaN6IyF+qDhuqYqnGyhhX3XJ5H5bau3zskDXNCBKvPz1PTq6+eEht
a7VnoN393bCSsOVzsuCK7jIJX+Cc7ivhj2BcwlBQeIO4tGVKanqAH/C92M2BGhPn
xgiMKaQtrfillEqiCdTwx2o9kiE2Z/7PSZ7qnGJb/fzry27dNwiP5DTV/s8bRNtn
xFEmTBnZp550/bekeTg0jibbfUMhxQpM6+iKIbEzTvCl6Yo/tHGO0LhULTK6lj/V
h21fBrjOpsikVfY52PWZ0EqmhmbM1wjpc90/0ok/QMFxSvTCmFzRIlGGaGR13S3f
L8oLnQpz6vWaD11JbScaWc78lRgLvFdFvLpE40+MEPqpJEz5Djo3Cq54qRJBPL7n
x5Q9RSA9TyKnFWnO/TIL/Mn4BCh39La9b0k31L3bd5JRsZYWGG0VmZoR+pEGWPJ9
Uag0k7PZaJK+NYhQJ3zTZI/mPu6gpR7Snsg05f0uuykJGg96VkRuWs1D6Wb5L9xs
w2ECilExwA7u2FuKIJRbL+iiDTNiN8yapX6NyJAlYHfEOL1R8Zmb6i2ximbp8ua4
wVTS/W5CzZWoNY8BbrNCmMXyGsVeQfr/OMIROvssYhz1UOA7TluzzghRJz4a4lQe
uzVg+IMYwd5DNenFTZZmQpFjsB416LEraux0f5sk5jL42g1f5E6K7K/sQ4gs8SvL
PixLve8k60ZI2oprDPEjUPtIzcUTxSv4SgvfhzGp5MbzW+aTK38kuqasu6VQuNTd
GriX5svbMiJR702sOQzBIZJOMzk3EdC8kzZkBv4S+kBZJHoLDVOndr3CshBHiUMY
CTBpW9xCJaNXefVoHPQTAdl+u35Q+6hUuCBuF9tM+aLLxF1T4q+KfejRxMbnscaC
SNADb/uetcLEYB91wn+4m3qQSgs8827WnjmEBr7KhJPwFMpAkpJpjsK2foYkcf5u
bKdf0v1Znu8J+5qqZFlS/319syc/rwV2ftc5Xl1fZu5Rfw84vYL7T/apV1A89+xN
FoIbinSYWgNTqoo3OA/BSF3MWK0hgECT8V8vGFTV+3CW6RqEkqkQAa0yB3Ug0Yhm
VZYZzUGRCntBntfdMXfS0xVvTWA3bVIxK204TOoXaDVYAFLIprZM4E1opQd1z33q
Wlo3Tlo6w1r7V+YFuQfprBa2SWrCEO/c+cBf28KKiAOy4PtO+UJIheF75UX6n69d
WkSM1h22GNYnok7RbZiPZyEXH3l3J83vVcaqFaSJfC57X6CXfLItmo3FWqsSmVj/
oqG6giALXhmkodGjl/0kHcMc5TXqnXR801qEq9vrRm08AJ8IFLg0BbOnoQ+bkyTF
s8Pk1cUXw4rvyfZ3+ioehCw2sS3hatUmIZtNukUTri9ZFPl4P5pzjOt4VFzbT5YK
FQ1fXgDE6LIOISWw4LhTIQ==
`pragma protect end_protected
endmodule
