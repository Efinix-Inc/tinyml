//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2023 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = tinyml_accelerator
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Mon Oct  9 16:24:47 2023
// ***************************************************************************************

`define IP_UUID _30aa6c7c6224453eb5782dcbe16593dc9d52aa7c
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)

`include "defines.v"

module tinyml_accelerator #(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 6,
    parameter                       ADD_MODE                        = `ADD_MODE,
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,
    parameter                       MUL_MODE                        = `MUL_MODE,
    parameter                       FC_MODE                         = `FC_MODE,
    parameter                       LR_MODE                         = `LR_MODE,
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    //Convolution & Depthwise Convolution OP Parameter          
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,    
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,        
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,        
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,        
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    //FC OP Parameter         
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,  
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE      
)
(
//Global Signals
input                           clk,
input                           rstn,
//Custom Instruction
//--Command Interface
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
//--Response Interface
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
//DMA Master AXI4 Bus Interface
input                           m_axi_clk,
input                           m_axi_rstn,
//DMA Master AXI4 Write Bus Interface
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
//DMA Master AXI4 Read Bus Interface
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);

`IP_MODULE_NAME(tinyml_accelerator_int) #(
    .AXI_DW                          (AXI_DW),
    .OP_CNT                          (OP_CNT),
    .ADD_MODE                        (ADD_MODE),
    .MIN_MAX_MODE                    (MIN_MAX_MODE),
    .MUL_MODE                        (MUL_MODE),
    .FC_MODE                         (FC_MODE),
    .LR_MODE                         (LR_MODE),
    .TINYML_CACHE                    (TINYML_CACHE),
    .CACHE_DEPTH                     (CACHE_DEPTH),
    .CONV_DEPTHW_MODE                (CONV_DEPTHW_MODE),
    .CONV_DEPTHW_LITE_PARALLEL       (CONV_DEPTHW_LITE_PARALLEL),
    .CONV_DEPTHW_LITE_AW             (CONV_DEPTHW_LITE_AW),
    .CONV_DEPTHW_STD_IN_PARALLEL     (CONV_DEPTHW_STD_IN_PARALLEL),
    .CONV_DEPTHW_STD_OUT_PARALLEL    (CONV_DEPTHW_STD_OUT_PARALLEL),
    .CONV_DEPTHW_STD_OUT_CH_FIFO_A   (CONV_DEPTHW_STD_OUT_CH_FIFO_A),
    .CONV_DEPTHW_STD_FILTER_FIFO_A   (CONV_DEPTHW_STD_FILTER_FIFO_A),
    .CONV_DEPTHW_STD_CNT_DTH         (CONV_DEPTHW_STD_CNT_DTH),
    .FC_MAX_IN_NODE                  (FC_MAX_IN_NODE),
    .FC_MAX_OUT_NODE                 (FC_MAX_OUT_NODE)
) u_tinyml_accelerator_int (
    .clk(clk),
    .rstn(rstn),
    .cmd_valid(cmd_valid),
    .cmd_function_id(cmd_function_id),
    .cmd_inputs_0(cmd_inputs_0),
    .cmd_inputs_1(cmd_inputs_1),
    .cmd_ready(cmd_ready),
    .cmd_int(cmd_int),
    .rsp_valid(rsp_valid),
    .rsp_outputs_0(rsp_outputs_0),
    .rsp_ready(rsp_ready),
    .m_axi_clk(m_axi_clk),
    .m_axi_rstn(m_axi_rstn),
    .m_axi_awvalid(m_axi_awvalid),
    .m_axi_awaddr(m_axi_awaddr),
    .m_axi_awlen(m_axi_awlen),
    .m_axi_awsize(m_axi_awsize),
    .m_axi_awburst(m_axi_awburst),
    .m_axi_awprot(m_axi_awprot),
    .m_axi_awlock(m_axi_awlock),
    .m_axi_awcache(m_axi_awcache),
    .m_axi_awready(m_axi_awready),
    .m_axi_wdata(m_axi_wdata),
    .m_axi_wstrb(m_axi_wstrb),
    .m_axi_wlast(m_axi_wlast),
    .m_axi_wvalid(m_axi_wvalid),
    .m_axi_wready(m_axi_wready),
    .m_axi_bresp(m_axi_bresp),
    .m_axi_bvalid(m_axi_bvalid),
    .m_axi_bready(m_axi_bready),
    .m_axi_arvalid(m_axi_arvalid),
    .m_axi_araddr(m_axi_araddr),
    .m_axi_arlen(m_axi_arlen),
    .m_axi_arsize(m_axi_arsize),
    .m_axi_arburst(m_axi_arburst),
    .m_axi_arprot(m_axi_arprot),
    .m_axi_arlock(m_axi_arlock),
    .m_axi_arcache(m_axi_arcache),
    .m_axi_arready(m_axi_arready),
    .m_axi_rvalid(m_axi_rvalid),
    .m_axi_rdata(m_axi_rdata),
    .m_axi_rlast(m_axi_rlast),
    .m_axi_rresp(m_axi_rresp),
    .m_axi_rready(m_axi_rready)
);

endmodule

`include "defines.v"
`timescale 1 ns / 1 ns
module `IP_MODULE_NAME(tinyml_accelerator_int)#(
    parameter                       AXI_DW                          = `AXI_DW,
    parameter                       OP_CNT                          = 6,
    parameter                       ADD_MODE                        = `ADD_MODE,          
    parameter                       MIN_MAX_MODE                    = `MIN_MAX_MODE,      
    parameter                       MUL_MODE                        = `MUL_MODE,          
    parameter                       FC_MODE                         = `FC_MODE,           
    parameter                       LR_MODE                         = `LR_MODE,           
    parameter                       TINYML_CACHE                    = `TINYML_CACHE,
    parameter                       CACHE_DEPTH                     = `CACHE_DEPTH,
    parameter                       CONV_DEPTHW_MODE                = `CONV_DEPTHW_MODE,  
    parameter                       CONV_DEPTHW_LITE_PARALLEL       = `CONV_DEPTHW_LITE_PARALLEL,
    parameter                       CONV_DEPTHW_LITE_AW             = `CONV_DEPTHW_LITE_AW,
    parameter                       CONV_DEPTHW_STD_IN_PARALLEL     = `CONV_DEPTHW_STD_IN_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_PARALLEL    = `CONV_DEPTHW_STD_OUT_PARALLEL,
    parameter                       CONV_DEPTHW_STD_OUT_CH_FIFO_A   = `CONV_DEPTHW_STD_OUT_CH_FIFO_A,
    parameter                       CONV_DEPTHW_STD_FILTER_FIFO_A   = `CONV_DEPTHW_STD_FILTER_FIFO_A,
    parameter                       CONV_DEPTHW_STD_CNT_DTH         = `CONV_DEPTHW_STD_CNT_DTH,
    parameter                       FC_MAX_IN_NODE                  = `FC_MAX_IN_NODE,
    parameter                       FC_MAX_OUT_NODE                 = `FC_MAX_OUT_NODE
)
(
input                           clk,
input                           rstn,
input                           cmd_valid,
input           [9:0]           cmd_function_id,
input           [31:0]          cmd_inputs_0,
input           [31:0]          cmd_inputs_1,
output  wire                    cmd_ready,
output  wire                    cmd_int,
output  wire                    rsp_valid,
output  wire    [31:0]          rsp_outputs_0,
input                           rsp_ready,
input                           m_axi_clk,
input                           m_axi_rstn,
output  wire                    m_axi_awvalid,
output  wire    [31:0]          m_axi_awaddr,
output  wire    [7:0]           m_axi_awlen,
output  wire    [2:0]           m_axi_awsize,
output  wire    [1:0]           m_axi_awburst,
output  wire    [2:0]           m_axi_awprot,
output  wire    [1:0]           m_axi_awlock,
output  wire    [3:0]           m_axi_awcache,
input                           m_axi_awready,
output  wire    [AXI_DW-1:0]    m_axi_wdata,
output  wire    [AXI_DW/8-1:0]  m_axi_wstrb,
output  wire                    m_axi_wlast,
output  wire                    m_axi_wvalid,
input                           m_axi_wready,
input           [1:0]           m_axi_bresp,
input                           m_axi_bvalid,
output  wire                    m_axi_bready,
output  wire                    m_axi_arvalid,
output  wire    [31:0]          m_axi_araddr,
output  wire    [7:0]           m_axi_arlen,
output  wire    [2:0]           m_axi_arsize,
output  wire    [1:0]           m_axi_arburst,
output  wire    [2:0]           m_axi_arprot,
output  wire    [1:0]           m_axi_arlock,
output  wire    [3:0]           m_axi_arcache,
input                           m_axi_arready,
input                           m_axi_rvalid,
input           [AXI_DW-1:0]    m_axi_rdata,
input                           m_axi_rlast,
input           [1:0]           m_axi_rresp,
output  wire                    m_axi_rready
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
oHvqb1SH7/LZ0uzlO/XyeN/DEDAW2I4uasQ4DaEkDjFsDNCUUzA1zY2tyzTrdzLY
Tz6NDV3WNRefUdX6Xt2FkCouIks7ySCdD/x/ybRyCkEQ8DDJvQl6LoS1SfBUl+Ok
EHdm0A+VUpmdwGqQbCF1H+7qZqZ1LUGDrHx6mtVd98snfeAGMR37Wql6zQRWjAnK
TXQWfhN2aMC6u9+A7YhVKOl+S5/9lxPksSHEsghiOp5tJXc/oy67PnZK/2L3Jw6I
i2ODKuglTjjp8mTlR1dRdfCeriZcfK0caEEDU9zdyR6EIEXrLlxB4r08+glzMHr2
FxpR+tjuylI0AyEOKa2ABg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 56016 )
`pragma protect data_block
jNyHL/rturF/cu2VKtQGCSKcRoKvjxul3ZSHtky3BmEmqgxgCYyLnkInhUvEFjYc
uOt3sxSt+eOTegFrRpcufNPZE3mY+ycO0hbIAa5ROyYKq7mDNwFEMqj/QeRwNMC2
Mb7XHA+tl9E3AVkCXWPggNksALXxVuZsoNQ0clZT/7A7e5APMNWNcqdAog06RERa
VRosIFwDHJeofBc1WXYsOfdm9fUIYy87/jBEehwT2Ceff1FobP+jvf68+wbfspuA
2XayRyqIIHnZ3Tgf8rlpJZpEh9O7i2xDJdTDKgwg+V5c2mxTTS/cPZF2c99RWgRU
GzbxzTykqE8UoklwuMvGZ6WDX3MmlYt47WOuYJJ0S0xLzxal0ZjH3qw+XYcjfIEL
Agpcc21Uaa3pPZIRsbk8IR/QUeT0uSb0C4Yb+qMSUE5lysfbizh8AmKy+pyUVxjz
O+1Hy0TMYZw+0LexzZGVONd1vYhv3ATdTQVUKx78QwGkEIyT8XtoeDAr9xrUDLwM
98GiaY1gvLfkoDsEHbfQkktero6jDP4VUPbdxFeLst5LMlk+EBPfvqTFQzOrZbvM
Wb11lwUlUAubJlEuVgqFyC+h/PBXlOYMo3rvMCb4mI7MQ0DdbhfcuE7i5cmXsPMF
UwlCQKo6Ng9yoGA8seycdSem7YqgRX6lNfoJckgLW+KJswYqw1W7EHMblAyavFBX
b/XxuEwnrXsS/9x99ZqtUK/T6DoNu2k8vLvnH0rup7y3PTQp0VfhMfpy7KesKDyR
UbfUcr9xdvI4m4/uxSf0DBQbl7cOSQQPSodb/iN2uZNQ6RNYApbF31wQTnH+QhjU
BBasN9GjqVmQl146Bj7mSScyy0LZf/32ml35FBJBdWQVYba8gic3Oq39vYku0soI
CnfGJLXUyFvzgW7RF6T+gKzpWlPXGCJZ3HXjgieLmrqaTMzliazq8X0RRq29e7HC
jCVC/FMjHek8merZzgS6yONXpI5Q0TXxXcDPIKXFVlCaCkKyXCbjkT3lbyTIQ070
cPKf0gm3ofXx+f2LpcjyST0X/yqDW27aOqne5S7BPxc13mAySZe+I5FMS7CdaGNp
rynuIZ9wo5bLdaSNTAzi5elsLxNgkCFmngNVSob6haz3JHWP+V1xP7JChEHsXCGo
ZcAg31ef1cFGN3nqA5qv/VFH3QXp6wCMtV/KbZnMJbCSnZPFLZR2n1PQQv5Gt5b/
myCtIQh3a+i6vfash/tPiZZg5HF0q1y9UccRWQBIz8EGxU8rb1eZ0Mw6l2Ojccle
yIKrDncPZk+xE0z8dnTVezbhywZc18y9W+wxfF8wsKdfHuxwtxM5bOJOIXbCpLoO
ID7HnVdUrmDej7KWX3AbZjt45d25kdCDMCqm0ua+ET4JbXSDjVgmTSrjGBw5hlrW
F+zZxR7i9w3spsoDD6bdckbl6wRQioCHgSAa96ZZSkdWtFxt92tw67yBvfChSxZb
NkIZIi2bFeQFNTyUwoQft23VXqAasxVbjowvV5MeND1oByYsS4qSu63hL++r+e49
hK9hPDcPPFZwTGv5EGX7LqKFoW1BnK2hti+lPI8ydI54huYhumarIUEnzwCyoNfQ
NHmsRvcVJvtWjhfHxtn7xdnlju6CJq49gVsSQD2PJDjrzhWmWtgheYEUtgUIdH7R
xpiSwuV/O9lYamoFvaS4ROBRg7VBEMaPtE0Fe+wl7+yP+ZsIMoHbQfzBPTQwCZAL
RX6AwmW0l2ZjMmOqYBBuwlFTfiFLjupHZUOJICCN1T6MXxG20dQch1KoYXvo7Cw8
+2kc4UoJ9vdA4+5iUY31XLGRLJjUROd0zlxZ/MTwEjw9tUBhIYEQeoizeGGxn2Dq
vjlydYWq7jytogYvTEes+g5pkp1OARTLGOrevDjCScQHrmCkCmd38FLWGE6Ph2W7
nm4Snx2dyx+y2QJ/ia3lgZGtmNynOLQPnPtxbAei7dZq0VBJ0p+xtFxv42s9g44l
D3lsi2lY0vMqLQcOgrxoF8ZUPRxnr92+EbxGDnivRdCofT0zgTEPmR0swKyG8di4
G1ANOig7mk6jDPNcTlGc8yGuQCt0BUkFADCxNNDWGWT8tB5wKqzbjlPbGdlwOS/N
4cxSxY7W7iRXZ1RAdEj0wIht3zeFl4NpEhwBIaFxGzNyQwy/tnk0UmfmPZbCNyKM
ulPfXjKVgSe8eYYqtNSBeI26019S4+AjGMwgIarIEAB6SIDdnMi4BXWj6ETIxTVK
iKQtbgXC42nEutm9lA7Byr1B2XASCkKbeFObz+pIpaMRtnJPJXixS2RSq3F3o3Zv
w4G5GIrR6mysavhUqXM13wDXPrl6wAC4cRtk52b4J9Dexi7KC5BIZDrfvzVgkodf
CdyaNntpTvduUgSHxl7QkMntRl6GV0v/uxMscqmOipOUekXc5G5DtiNmTBqyobnj
ut8dSdGt7lRghbi8le92Lh3Iub7AvZSHtoTvE8jFkf6LzDUJDt0J5ih07FO84evL
AX0YyfJeOaHxIkZSwRjPEfgGJ6wBbMb3tMRumRiSdlWgttCoQXF8H1z4ky3VR9Ez
F9/ja+bC9l6wIiqiQknGhHuYy2rCYisV9vr0z81hrDpC5KaspkgSythIU95M4hFS
wy+zG8X/DY/CF9me20ugWW1JomcqCVq4Nm/3CcpPMV72TbWqLZc9DUz/YNnOZnah
233Aqm0jy61iwSbQcZCrYNPedeKbuEatOLqhOrK46CxtRfu+bKBRFiUBsiqzR+AG
5F80nqPrH+dQWmGANyiOaBlzuGWUzMYE2XqXoocGTiitnmPkZzgOLS+g0DtcEsLW
RGV67j3VyihA+cmZgv/QzreSefk2L3gun0ALZYhAORv7uoPTIe22tGopPadeHcO9
FAaX+DbJaYYtAqKjru0obGmffwsr705FJrBmDs/y0ryB8qRUrSubJnpAqeHbbyXy
rTR2JWkB6rAcS4GjFj+alHi6LLqDO/t7NRLrX422ipSPRSVqGNtcMHQCN884fFkB
uvzZwSAMX3+4kv4iHj807k7xV8sp4v7UwJKaczpSVOLrhoPejRBX8RX9MzXX+D4y
LvI5/CBudLK2hIiCKYcQbgcpzNO8cgj/q10NIrycbvc+0eHDOl7yFNixYLAoil1W
u2ODa6oHvXLMvlAVawZI48nrWJIHZ1PUUOw3Coi2jbTMUmRUL1t5i7TDPIdQFRSB
KgQpICDNc2xH8RjU/u4AizyFDcHf4sJnQkRom41PZECybNDTc4+/JdYgLlqIbrEO
d+TDTjOmGF4uioCVOb2ICeg2c9uvjBixHclKisSns2RdO9J1KHyG/1bktOSL0X8a
rcISTKcEpZR3iV56r1lJMogNNdX5Izib4I7iJ4l+Jk5infEAFMF8J5E2a6L6ARua
LIGZnEWbwahDSIKTRKrzto/untKKRezoUslmlHHwFabfZAcC+wXaDUUiqWlKDbNp
UNHRJo9bbSqQSWY5X2YKe2sBA5549XNVNooFZXYdnvZQCoICWDuQK0aB/q192owb
uDDx3+yyFdTxScjHf7ZmrtqwrCtjyz9d2YM1Uw7omCxtxdNeX599i3HkVf/3c/pX
05qZpiOZix2ikt2d+rrKWACwqFKZtdsKpkEOGQm9yct7YDZ3gMWyzFOBmWXeVQBL
uV9warXJyqIsPsst8repDK3e4j9oBc33mJar85DsT+WWoSsWRji62auM/TKbd4K0
GJTxLCjLW7fvnFBJm9ipn10b3oVAJORg+Xl9seAnFI8DAXWsgz/f/uVavR2I9jGw
WsQHQghDG2EyYhjzBbN7+w9grgY7+baCnafHULhvuW/DRtbXUMwTsk+oA8e6MoyT
lyV1BCAhxrBxHxcu6HH+Bw4TWo0C+VKFIixRMS7nHftEp2Cq15MDx2on9gQQlJl6
wAbP+cOcHh6cbRLJ9XZKU6BB2iGzVLQoCdBiaXZf1sfBz5Ebfn2ckldDaZF5nnqL
8B9o3tblBqXNn27OTIqJ3Axz+24t28y8McmaYh/HT+FErLrea8IpV16SLCfn5lQ4
5iQl9elCHaMT0yTUFpGIxtekLheZFKSSpDVjNjsKs0e/KZVFbcqTJOyxDORQbubW
5JpRB79CZD/2lchFxxeZe2a+wboV2PfEUBUhCXlwRqmUDL+XaCb6FHFjizgUTQBj
AGpvPZhjiA7P59OvBtdSJ0fXxxt3FzQm+RQkOyf8vOZJ79kOe6MQwMec1TIl8bnG
von0BWp1wN4GXYr2TmNuISe+m+CvpJAir0P6HO0d079R5XGVp2UCXC31LGovqM5n
v3QoKQ5e+FzE8svXjFTj1svlDwDoSVFeGnX0x2nLV0aHY3sejPVbNat+tMQ8lHPR
pzNwHdP0uwxnYL1Afh6aCcRuHBKtwDWYPddr3T6RSiOX4ECSMX9Z0mSIIC2Vl1QN
0jJH8Y9QTkeidhrJmkYIRRj5j8W/02bMZUk+5cUlUuylL3DKA/FkvCDcpWAA2xaW
PfBQaOwc2+OYgSP/7vbyn1n28EvO1w88Mf14PUoR06gFCsP8DP//UXqBEACI7tvt
zNYbvRCTnwT4bNxKqhxeKY8W/KHNfP7kbpbi1iEi+OetVx2dEzVG5R13RHaggz95
tagTVw8azR2F7rpKOmD7eOAtTEnedykTXJiwK984IbTF4mrjili7mrlaXeu7JL95
Be6GBidMXLIKwmaxs6WWC4z6z73kr3r3P6tzMO8YeeO1l1U1LuMB6MNdIlBVX1og
SC1MAA1hx7fX7ZCigj4GDfa0RLd3DbSVqut+LC9SxHwbWuJcrglQQoHmw4D7Ndww
7DwHZFd9W4ysVsJo5/IhW2mY8WqF+1Z+9v3lvQ2ACJ5wxhk30RZ8mEn6YQitBOuf
IQh3ViWCwZVE1h0KY+e1lGAach6zvUevozNs1xCsez61Dtwqf8TZ+KCOWJOv6y9K
pCeEsijNy8I3EvOyf5Nc1Lxm5MzUwoD8iFgp1MqepmK4yqiqOryPx59uv4GNcUAH
2k0hAKLNWKqW/2FY0cCWUlWP1kP+PYGX1dc4gnHRbBiVOMEI2a+D4spY9Sva2qkM
0uQ8essBoR1/BjcJ9O7zWp/wMuxq8y39IJ19jbmVnfFV+StHeaZii84KQW1egA/Q
jEYR6RhYqAKV81eGgQGnOuiC+yC23ubYhUKa4rzMS4qLfaoVO6LjB9aEf0mkMpop
t78r7UWfedrFLDVkL2jI7aRu/jpfufpkdHh5SSXqR3Q7DKnJh9vn4PGCYuEL2PuG
9yjRas8JvCEJX/UjxUjvy8Dvi/ciY4BpQYsJQ+IdD6h5t3vUEj43MAI8ka974N1I
1FfVw3gpbbyGc3c4R/FVT9K/AOLPhzingo7yDoZ7+Qd6Gek1xt33+qfaWijqEIOO
YJk/0pWy3fHKfHo0Xw14NfYQ/Gd30+W7nsFKooJJJQb4c0HCE0LyMA9eWp/nSJdy
SMzhi+ESQLwCPsneT7sVjGB/rQ4db8vrcPkWUcTpW6iGAx1mcKKBp8l8GY4Xa+nF
4Gov1jyA18BcDDXx8yqvjtL9uKCTk/GuFaaU9egHJ/kVj2N64UQm3f4L0tvYzJL3
PeRGRJ6an8S+e3pnzAYtqfX8Aw8Oa7lTDALFooAnNzli3XwFAbzLfl7XMUaO02CB
yu91zHWII0teSC1JzarVEzkdCYDJBkEcE4qzhwoewV7fBrrkGP6Tbp1pTrHbPaEq
E+ohoF+gUsCV0F0q9ySTkf8cwY+LZzfsHBSC/13xhwvLGQJy6HMSIEKhGJhYmU4f
7j/uc4X1mlqYep6ONOb33/dqIZaTJTUq1a3TbIHyx3KuvePAaZz3wTNWakFykNKS
DYY9TaiPoTh8FFMHgqy0kXibTh5rNS2RL+4jXP1rMbfTR5CXhFJTnRw177VukY67
MVX7z8mO6qR7zUODQGbdzLYtK3NdTpSACe9KgAwIla4xPAWZCboWmDQo2hHgKuyt
v0ZpP/U8ZY8FlDn/ygE/umRHafcCgysjmhe0QaJphQ26tBZXAVPFd2qOo5IzPTSf
A2RhvYIoxLb7IG0GybMl9O5yrOVoaorobJAd/5XYB+iuKuTWzazNBT7gmoFy0x/d
ycAj3xdCX6CsAnyTpw4E8iz3vV7RaaTvDbyzvhDub1nwqjRdSGFJ4zgAUWdkKq9J
HO+0BagQ0Fb0MuxSd0NYuRAXVNVtSlOBSzyJBP20l9c9en0zl7gYNx9wxkB+e5hx
fVG8XBgNVRoNlmnxIred1HgWsMm/TG1QSSUBXMuNK2wNBoA7Q4KH+M+hT4+FcaZE
h6KXPigwrB7eUm9uKFXa2Z8ZHRpuhfkxIi+BVshyZlh7KlWHpiSODpoQEjxUmWYJ
29HznSVGN+jvByoMLjnmsSci+Y/KFaZIB7Rc/uHN3uubAzCEm1ymTH9aRQ4Uu8/n
fAs6gWk6qtTx5ZChEeVU+78R/fClG1x0K7Na/2VKA4k/xVEqSD+x8b/0p6eC3rdv
5oMekLWNuiTqLXqNoPNO1VjLn+u5cJ4MQDrr/vGTLcOt4YFZ9D9JcC9ZIyQ5hgWl
krpXOXOplg+o/5BSu7WaCIoKIy6LtTr1Yx0l9j0GeBfJVgsPo6GrMwFw0+Q38kri
EanzQPKpw/jsFzPKNebXAVBKOYgJuN6+snKsBRXF6ZPZes+MyZCE98AxZ58FhZ/N
E/18bkFkl5J1Y1ugc/lSyyczlMJbQyIoZYYpGkbuAZCAU66dKz1c/ufuxg76FuRf
EQTPnu33lUpJityvtg9jZCioZSoWzWYG9FuLem7OdPNlWuk1AfkFhgWMZQJwW5GK
vQNd3ECoMre+D6Oo8PELUDpI3E2bhJ8HRrxg+af5nR/covcZFuZKkRCVFxoU0iy9
Ob5btA1q7CC2e3cqgBc5kAh28yrwo30DiRQIwy6gdq+60Od4FZ7tL6AG8mNuAfsY
SokQku6n4ZdbDbMkjaqvRLANWP4hCj7/qF93nbdZo0kAnTrW3IEZLmiaqevn/8MI
eVqxpYImuMgl2bduHnwd5TFM2IVWxMnUVDT78TuRRSzkhfSMT98x0JhMLPU3SVGY
CXSp/z7fHtEl2w7jWCKp9Kks5CiZ1gW0oLvswmhVKSFcSzj0PYonz9v3NrKDMcur
YIl9zUUVU9VOaQE1AL+sq9h4E6UFH94c+j7/L0jRmquyGcRO/qBAIiJHxceBXl4A
liRQwDxZbLoPOmM7erqlBXZaKq3AUmHrNnY4txxQ/AA4NGiHkwhSgUtWUglVAhnp
uUq6KHbWqGtPqhO8H5gT+73zSe0wg8yD9Hc7e6eM3jxPxsMyJf8DPl+SIfs/o9O5
x4HwVEqmnBIdA5ycwzLHFAIXTEf27qMUBhA+RlEQ5Ijr7CUiW+H0rKsYdlKv60/T
Qb8bn/Pe9Jn+vvJ4JeVSez+7MU3XBCnwnUUoz+BA6qDb0IDUbr1tfLYey0JSgCff
mRAPoZ3ZZ3iDDol8+x6K9Oj9zkFujCztHTdtteH0V2XtWEXxXlzrwtUaBmbMBCyA
795X5TJfYcjq0kcWn/wYC4Sbi5+XMP8NrGQD5Gm4aCyMwae529T94Sq5If+JUuC4
2G5GkZuKuucavBP68evitBTKg7p310BbPuhMPz1Q/BrqsukdSBK9dc1JuTkL5tZ8
tA8tVLgf7CjwsS39NJ1No6+ymCZvxuTYCRH74DHWl91POcNucC8LBUo4N36S6gEt
DNMEl84XPMRIaS3HFVlJr1VUZqg/pGFFgpii99tBEu40F1APxnLfSz+FqCHEyBmF
+hd/j5dC6rOU6gdElo4Wsi4NZfBuSf7uldPiYlyleQ/o2UNwn7aWcrVZjhGDO9CO
Y8NFxFcD9PZoQlSYwFiqgAbJodJjUGWRZbbeWuvjNqJBcaQG2jibsvUfOLOX/A53
aR320QrbZi91Z9/E7Q8JHPqhIOFPh1rI4/s9bH3m2NnN7hqSGo5SHdWJcKFwFd+I
4WM4c91ZfNQAkEPlP2rkodBPDMQ9/PXl/apc+nV2GPRiES4Tn8N0FyMNkrxEQkxp
x1ceaX/Aa9iWiuSWJGnO2meRxPXXyIJlJLRBPdQ6XCJ8oToRxQbkHY+bkRjhF3bH
D4y9Qfx0pkE9LXEcIVEIjCIlTzQI0e0c56xWr61/L0Ly2xa9tVKtwhFJHB3EgC45
J7DLIK8nm5X6dVXn/Fh00QlQBilbCjswyKVVGXyh4ItXqVLQBHq/5nVg3D4LIGcj
vAVDOQqE5/uiF04YM5+XJ9S5TeyQZB1NP6yZHyxbCWXru+me2E0soPUKyHqlDQz4
PhWTe/0bqGY2VL21Xwt3v/kVr3RfkYSYMMssE8jiWfNkldV5cM+JykZoYnNySMwe
Teyhyr2ZUQwrRzUmKOqk/0wAL9uxkG32rDc2vKsQEhiY+46nu+mpa5fAufXSChC3
6S4FmeYJz65PW5dT5hiiPnj2nXq7jEVeRtc7s34pRZBMhtnfPMsDgQPtbPhH1FRA
oF6onoR1S/hpfgQ/3fTw2Y+1AZaWstxDf+UHftnE3PDd+KC/I1nbJjb6TZMb7X4J
Qwnm/klls+0rZ49ri9T7JYjN5I8Qen7PlsZaohcxnvXVK/3xaX14biNbvoak+87L
KH24wWZlawVq7fht8ERoBDJy6gEdqlfVk+HQZcrSQ1z5Y8Cj57u43wDccWFERy6G
fY7OjXkYDAIOu5z8CYEdTu33JzheCvEoYEY20T1xhkC2Aww2s79eC3J/yOYDV2ku
Ke6Mb8418VpxOCBqj2JZKNpGxQKZwPnMsspxo2O3d00UoReEkImAMuDT862sGEEI
OLSazjrLZWTzZqyJcSRv+M4yN+JAptBEEl3YE2Dp9g63cnNIL9siRZLq5x7JreyL
pXw2ZRQNybi2veDMe9MFivqtIqS0qSoUUMNC4eTiNAEh9eVPYTBGIKkxrQ0QSTxo
6P4Wkz7d9P23s67M+QP/GYGU6T1WhuZwWrutegDjyTBTKQdMAVN/iDKcAoITuAa4
QkX/cszdZt/Leppkj1H52eOBs4tSadfbqJlscAeD3HmeeOppWZOzDWVbVAh1Xxs0
pEst53GYtl5tSDyxJMoGKRdTZyNLZSt4SSu30gDfZyivy6ytCP7C4ATzbi1LRrVE
IUkaihp4G0Cv5xLT4b+52Armrf1NyeDEUlOBufJvc/zT/TlkOTuplAjHa95ZL2R7
0Ylb3/aCdcMZ2WHZVLJlB3zKKvzoqEdKjmRPr2UKQV9vqHR+w1Ym3/EaVOldnRlg
GzNnQPr6DsVbvyaV+XShhMnABtwHKlWWA7s7r7rFdjMp9FBLOg+ls2QlW8knjSoJ
nYx28Ax0mRAumYaI9EIC3c+0Zxog1diZeaOud7emncrL6YI+EWGZpDkIoLbyK3XA
ipozwTI4iqFPcSdoG+uVDuhGgMrQdsro3y3zxQFeOvV8/sUJ+PMK5+oNbYNdyyPG
NL1o43r4aS6i5YNaeGea1TLbg7jakndizZc7A4cySpKLJW9duR+o/OC2j43UTFpI
2PrLcKuH4zKOWqTpuesePjpzyUFI/H0QCHpPU1+lMd7DzI1MrVMLx1Jhy87GrmQj
ijP50iIeodJnSkgcAuRrMsfBmneOjWWD1/emb81Kn9pX0VfvxXePG7fUALat84ud
mZmYRGFxHf5YaaHAfErufKbQerXggR7X4PxOkY2U9zpSD+bmqYVvde20+EHtHJBT
ukj14xa961BqeOHdOjAJ+bOVNcd158R6C5Ysr27vQcaLKCxbHwGdvUaGswBEojh0
JLJM1/72VQL+4LzM3rAgMUT3H6Yad68o1ZiIE2G0XU7ajTcsggCySf4tQHCkjyky
O6r0TlZMlIpiVwocmAYJks8FK+YvSjduRXkItm8Etu/vs29zI2mvVV7YOt2UgZD3
kEPQ+ZC1iB3UZUevxJyvM7qA2H1QrC6CdSM12xxKiOulH30oacH9pnkLqVW8FouD
cDGtwVsNtHeXAMlAOo3Fp0gahemUoyFhCikYaiXVsI/whN4jCkT1gu2/oj8JrE/w
Z5rXBvFFbQ4DuyutMQjpJQsruSKO7O4ao6VCuP6/Jt8P307qB43euRWAfp8lNZ8p
cl6sYb6hN9gr0bUyAanad5/tO41cDbF/9VoO51qQOCVH0Jr0J/sodpbVLpEVpb5t
zElLt2FD0HO68Y0uSsPi2qeCmZYsnsrieTJ8ijakWPKKpiohDRG8bJ7JmbjiL0wB
IZp6J5gC/Q5UvtSIvv1vEKB0ONLqIgq3AvtrSkzE+wLPcCOWS13z5migKNyZLcdw
lVBRBJdVt+BWRBkF0PEcnDPkxU2KvQ6RRxUKPdTdAF22hvSult6SkSTGGLy376zZ
KKqFRyDzFts9WbxX4GDnKo9rYM+nsbgOLJHqwh39GoH8916GMIqCfkIV+WcMmOD2
/AuEPXresqNVIfu24mc2h9nxbqqOH3JgZui4+wuXPkehSt4AQ9ffQu/3jdJBGNVC
0nnnVqHQ/uMihkWuDqrXUOZzpx421qSdnECtzsO5aXXG12sHNs+Yu54h+Y+BmPSO
DtXSfIt5V6gLf7GHqjeSJEFycQvIQPoqmgengOBomMHCDR+iF/Zh+xu3xv0FqQ3f
IUbUUwubcQmknDmLY8lGarvHNz2FBupjHt7XlChhzmmrjdEvnqx3AWenlUvgXxbJ
4TR9t/bMhCNTlccicDfe05vC7q6A+wlxYPfRJIOMy1/6X5qEhbBIOzPzOpIydUtq
Vr8nkxUx2uI1oA42IaiFzaSsLQZhjcgplrD5Hg1kQ9EOhinc0f50pSuJOMpxZZb0
Jub4IN94Wi4E1sOD8oSlbMb7UgepF1I0oSRLmrHrBdEs9VVpm2PDPK/h5H7YkPDY
qv85pbqZ4KhePGo7lA1meFVWwSej6Cqp5TjctOZnnpfHYQZFt1jLY9tTj2do4imZ
TTYU+9mslqRa1k3FJzaSBqaTCOVh/zpAPbuXoJEZgV+abidpWWFijdlGHvNWHLGH
Ts1ByM8tVXqqP0947pIdnKKYGbJcupfqmLoLeK2lJJZDT4QVk8DmUyV0rZDg5o8K
jruBwDhLwOAa7344R0udOMZvDuJ0diTTE37p4mlXijalC0mCT5di169QPpX/w1hM
OS3ZuVKhNvvta5GCAbjTevpxti5jJjnL8jZxg5T2od91soJn+NqL/WY88IvY+y6G
5gp7TqNF2ut5xiGK2yHhCx8V+0hXnlYZj5dHOkw+l3f5SUdbe6hFyGdsRfSgGGQ8
KKoPF8Fj1c5icNDWr4FHJv74/f8SDFePI3P5yxV+8kDAkAaRqzoO17/1kmb8urUS
Z/y7AJwdVdL47FEY8VhZUZlg7tr45FuOztEsqPoJrr1AlOyeKp1q6tevkkRkrOvN
IbZBP5uR3R3bme1ylTKHQcbYj/pxhtWkmpBQSrw1GW3Reou6OyJXEhlXIP5Jc8/D
wvxWykqbG4oKVXCAuMPo0hslvGx/Gfj7bKTh61csSB9WuUoFYhE1jXy+hw1RQS6m
oOQCxb5LjpRtrg++xrw72TqMU4h/NZYCziJugJaIBbNl5HXNZXOYv0cKw3GRpeM9
yZ484h2IJ83I7jQJOdbVkU23J2CzEXNIv25e+XIlU/mTZFTndXb5qqWwCAWXqu3Z
3xxAN8nGQzx8d/a8yRiMVUUNn1Rxf11BUtYizRT4yu/UryjSKGbvuj3WyITBQNbN
X5J7UzMZho1ccvWbEAj84+USoXXdnvz9UtpLVpzG2xl6+JFk2qN4S8svcO4euIyZ
0rI0AybiMhPLou9OKcRQnQjmWbKFHL8vyp2YcnzhF0LV0fviIVMwxoK+sO3zZ8uE
3tiqZNcsLxTPegwgq2+OCWnC1ivKsF2jjf7u1laRQxwFjkyoBzYxwg8XdtJG2LMA
/fUQSR46x/zeM6KkgsCFTuGYN1cPR/EeLmUSFfgNu32/0VmM9eO5DLo+tvo1ZNK/
u1MHLTcnvMaWIFdFuI4EXkUxbA2qq1CYA5QVT7OWVpdsyMgvsEVjvovJw1KxNnXo
YQCjMsVznayCFVpXRBbr3bNtFUL5Ty2/W4w2EnQSplazEFhHT8u6Fl/rM+s5gXu8
KCoejXKq0K6BpmRZFbpoV4m11Tx16LPEuxNKYuFO0ghnPtu0etqqFAklB48bAcEq
NgYkDWKGPIGxdLw6DnE11S4e98bXBwqh/cM/UmVBolXgz0Xx63DAGeoff6ldic4Q
VS5lBelZ4Rcsi/eebfr1MQM55Odas7jVfAg/ArbabNSfa7htyxklGSOpCp+MWI2S
e+/QWGaGEuqL9zT219z69bvmbX4Odcy9En8LlB3L3dUDdl852oIKggoVi7QvVZNh
3T0vcatdbyrYW1dhkmCUYsdIe0U0mbUNRg0li/jb08EO3+vNq1FXrUGo1O3SZ+R3
Y4hWFZR4qjvy+wwzFGYcgRx5HU9WVoAkKrGr05FrQuuolcXWS6YtUPFC+c+xnNMJ
RO9ZqsBA4W76XAnh47mwCXhNPd6jTvfcTcx0QsODPu57ri6Z9KZnjKA72QOod9Rf
0ppfYW0YAx99Pbih5W1KEi/15m2xx719+CRQRWgi3e1OjfRnOdm1W+QHO/HFo8Dm
t9TUVyV8ku42Ljpo/cFeleBWbVZpYtMtM+t2Vc4DnUOcUw4yNv5ccp4dujaVB9Ke
dAvhqF2ac+4Fje3bAGQJPiEj3Ss3iNKQJhbjF+IWuOkYz4BZiFNFo1/fvj9LQjC3
17ngn5mAowT47DUy5g/dpkBpf1LGL4V5n4unTT0pOuqfRUviYyzAoDgAyKDmcovW
I6PsyHEwdcMvuuYUY5YiJCcSwWO1FMU1AjiHLc53RixhqPhBpfP4s611P/ip/Xrr
EaTs7gJZIxSyYt8RMdYV/bzPJZ8hCs/xLSffaTLtWyjiB/kjHaQ+/pcYOLkW00o3
La01FvLTUXR4bYyOTN3YyhUWzNjY5/splQLhODQIwr0ORJgpd3++dYRLzM1pvbT2
S0rkESX2CUksW2Tg0yax6kf41zHTywm2aay/t5BaXIfhGAVF4y3rsst+i9Awf5kn
7uqUtULhIzCI3NPyHrv7cQ203NW/5nijwZoeYqRhUFuB9juXY0sPblaGMdu0K6gX
ePsDAqGp726Cgsv7STtjXkk3e7Slnnofc8+KK4XDEBxVDHnWkJ4ZkVZGdMvVExeQ
TeiEhBytbsug4km3jlMyI4O8BccTADKRuOv3oO4G0bkLN7cfUDZ9QA8PW71rlT6Y
0Iv+pj0Nnr3GMlP9DXTv04L47Li46P/ob8p1Xhr+UCKE67Da0nq5mZHvYrjkr15i
9iUqHJLKwGwN1WC+xu6CQ/+LmU3bmv6tP39w7m0w3aJrYqMXWZpI3o17cd+HISov
2g3LP4DTjswVmCL1ZXT+e+qIL8W2CJfClNf4wIZke+pwJIN2OLba9xljfKpHWwn4
RXpD6JWC0XSuOt7gqYBzPiMHZeZPe5StCguZ53myX1OeidiAuVH9ir6c7kCCf7MD
+Mgj7wtkocM3sFBvetP7K/cfryX8/Uwpydf72ke9eu0f28KkCDZgT608WU4YPKz+
5EPi8UMx6AiUE01sPNFDTjecT5Ar1mlTkLFjnhcU4P52KCgAmbgwHx2twuHsMEd7
K1E0fWyEE2Htl8FuccGlrx9mPB+9cwxy95cd3ni0LiZtnDPm02gGmIDm4RrQykub
C8lg+RDUXkVifm/AHF95sZ6nKcX2JNApKPGdyPoqlDlftNaLPoZVE1MvyuSbzxAR
Uau+2Q0gKTku3HHgMbYOHUAZlRTijCuK9JPkXA71ULU7Joxn1clyAz29PsBMdpiZ
w29PDtkHw14I/75TXvpzqKF8kKEEsRDHpZqavwnvAE9zHcQDBWZdmuSEepy43EPM
Im1Lb1JJsvTd2W02EiQj7Qd8Q23vYA7HxBbZURoOcgCu5QLpH51F0RzKlh4/rWCy
eYqsSseQohxCv8qWMhskRac2PGVLJPr4ggnV/zKPr0VLWTaWgu5wQ1r1rdQX5Xcz
8fl0Xzia8f9rL4GjmzXe2wUN5mmQjTyKr45mT4zJALnlfaAmEILviHOrFpfKLbda
vFupTGIZL0tei340Le6JDaR3qdg5gMTjsppZtsunfTfXBQLOQPqWiZwUSZA91akm
0xa0bGiC1yblTcYXAyYeryniLWepTYSeZlMtbKg1qUTA1m2cyMG/DtY/DnPiRbPJ
9fmSPyYCyQ5fGrYb+pYlhr2WrbUvNzvqw4a/gBAn9M/QrRpormpxHyOoOsXuQqQ8
RIy5KyyF52nnP4JbinutDd8HVUwb48VLG21Z8X0ZrjFy4NmRL2XHB8rDOabex9ML
f0iVxhUSjdva1+oMTe81SKjQsH3QtF/etsPGKm2lGZ2OchdX3t4bbrdrhzHxiTvu
Z3P2F45nDWT8ejy17YaNAbhldow/w2yIjG3+8UOXf/kiF0+9h87YnasZ/xqXGxBG
jE3ryyPvxAojXHXzTC3zshp9xFYa9OZcxRkfWFigUhjE5xJVzSd6q1+W+ExF4BL7
EL86NgFfpHSP2Vu2/uoyJKrwdyMlOuYnkp3tWuaoclm/KGv7SYZGye88G61npfrB
ngR6w5ixDWO77Ie/vmUqL/WkV3zjPKEEVSB551yhGSoDlTvke9BzJWUUFsNzi63o
o8p/eCIlXM+FWdQu9whgw899wExKnQpwN0uqf1TsCUncJAbTTnLaVOt2rE3ULZp8
ba1PRi9wciCja9YXncNr55BISSOxEGPaAiOsU8U33mm9gSW+/dNQCHQN47EB7f0O
4Y7nVRRXC63GqYhCFXqH+orPUguc5UZIBqcp5PC23NA2ui2sJZJ/t0yUnLMPKEsp
mSfFIdAKiyoF4RdvjLPteO1aVSvQrUbAMZtzBkPezJIZ0yeeUyu6GhA8S2CdGxj6
fZj3RMj9zFS9uJmiN+k7U66k3PEvzRN8pg9OS5rLVJ9XGRnIN3m2uSzTOGo+PyvJ
mRrCPOOgqDCX9Z3OzHp7ttXbibkOMvcsQ2boBnqIIO9VcEQ7UqXSxfvUTJjFlTVX
GJMHEEoR2MCKBMnvfnbIDYNEHZpySTUpb6wubv25HcTIGe2iyl3EF02oRTn2krDK
1LMSYg1qYhUxC9v3NC/ubAi6A1T/+jtNHudXtnMdAhbHtMTpmraqEPWgwBeLhjmM
29Hsyi0yPDqOtxTyIuiVta1MoOCiTbYvz5foSuAZayLzSw6thJQGU2AytpqZfCrM
7HwkgYhCuCbNRZah/2G9XkAXYSrCBweK02dWMMpy2u4//jT42zKql5YCWbm0xcD0
UFNGXN0eBBBZeUX7dAr7y3KGvSLV8973AKZl37nfuSgr4v1+HgQmZ10DpcftYnkF
YtsHkTJEt3TYFNysD/UKm59r9fIvhCvDlCNtLctNJmwQgDtm2OMNAbOW4HvQpKwR
bYB+mEbD+6MCNiY1DQeUUMyvvIhYakuIxzPDz46Y7UYnXCPMZ4D3Oaw7s2kIs98w
udHwiorUuG73MhOrglJp7kuINSOFmQTO5sbLMaN7yLHVneR9fGXAKNBqVr/hJ+J/
OTGmb1x3Q+gcDQi8SdeNxscKTjWunwT2mNXRSiyakQDFVOF6pYoP6LuPfNnbAVjx
eFEngKc7laMrHhhyGlsfh/O6ULE1HZ762krHuc0uSq5PFuThyo4HFVNOEtcTXyAI
92K2fAQcQClAJJ29EnMYWCtYy8CMmpHVReYEb4qZQMUlhWdys8ChmyBVsm2m8WKL
rsHBxmXmQmylQdkJcm1697lzAXBH+GMpRLjfgCNuqEEUoOCbAvYf/+we2lQEiLcY
dvS9U9N4Nz8WkesdozyZxXptS1H8DJRjsBCH7N744OfKLVZCmCgbXG1aSpcl5lvn
oAY34b8rh27+PTO5hYmK9MHZwZDZqiTULzXtMMUdMFLw/58e6PdmoRUthJYeysN4
hbpHLElfym67VRKrLNDE/NAtmoqN7et1vNCj4/X3LVrchh0UiJBBPRdhZ3IiCONP
nP3HV3q40AAOVLkDWCxO9T5t3GiP/An44GaNjLKiDYuto2cZQNuMmSLFoKq471VE
dK3uF0zW9H/kBkIarIZfxdtBHLKFapL5dKESTVB+Wtb6r8F9gFsTJOQeH1Nwre51
wEmDKdZJXrKp2Q9dmWxh8H2di7PL6eZa/8mxd366kZ1U9dhUKOcNPHs+u9oxcHnZ
O6Nm6+wPIxG2+iRKSNO02zkoNAkf19pI1oalu9XcBR8hwn2dq4DVit738398hj1I
shKnj/MwZn5kEfqtgwnjqd1ExRRjFyuOFeokpCmd27g6DLHgymvtZKPdQyRUK6dh
mUnlz0suODFXQl702PO11SKngVxAmEDDBCIr8t3Rb6wKA6F03CxNdyAufcSnNQHs
N8AfkmUgpJjofoa6yIVKD6rih9BCoqNByhD7mzf0r3/UA0vU1XfIlybVFQIf71v4
QoDPJa3a2elpUN/Z9OO9PFL516vjjRfm+oQRC63T/My1FGTKZLTauYL7y3tNry/Q
d3VS4LqavIa/H1DucteuuBwsjkDXwRtAh8rgDQTlxUp+8kZOIQdvm/LtUcBVx7az
413kStWk2NJLA4gOa0YPf1YnT81Ve93jVf0AQVscegrHrp8sL442VsNlrm7kLzpr
LK8vt5ohEJszFUPx8JkHONufg7dpQdjCQPpCoS2AqK1hsUoxdLueQipkHLGifA5a
FaBMU/ZDPSJdlf3ODBUaCxp1F+Lx9RHo5glG85/COIG1HPe4Q5UQu5vGzjrxIyUM
G1RfH31VeQfY8D60pWckD4ENE5pNysS6zD3uWj5xFGQVw6qlD6Che8Q5OD0CSnHM
7HlJ4CL2cOIg7iN8nZxvcLmFX9CHkzb5yd7VBi2icn7DIhMxTUOmI05GcGGC2pG5
NsvKBF5gnhuwizRT13cJwgXLmfB4nNxB1Lw/MX7Uh+vdKN0FpSv8+Q7i6mOs3MnF
hf4V36aHKit5nQT3kxwX8JZi1P2BZPqNsDz5YmoezY+2vwPIt0E5+YwEp9RKhrpP
1OgomjOUMxImRRPpA3nVBBBO8NWY0oTeTLSnrXHnBt46b8xEhxzAbrZsHZJcTr6v
l2wXX1l8oMiTk7PX2/QYCDkzCzHgTeZey8vaPSSEXOGtcyxQKsUb1Y36Ofb/W7Tt
JxLEcwbV6GGfHo+9P2GysVsK7nZDPcrc1s/i+19MFaNZl4VC0ZSwXCLUR1YCwJTX
pmIjYnMXdnrtrR11HwNZniKILGefqNscO6zljLbVeb8E8a7JZm9F0x/If32fkSOR
0whlKTLX/HArdir60eZLeFWQGQISrdRxpTMQLlYc0HjYUxrUNJdatiyvvNXLTsoN
DagVyUfhsfn/qmLtHrgw8+9a5aB7k4p4QaNlPdjuIBr2xEDb5WqQK7dV2rlZw6VQ
mo+kTTsDjm+JtsHTFI98oVlM8AzTn38Fr6N1xv6P3Xal054F0Z8EmjC4ywbrkhoF
keW0MZOY3VAv4YBTSCmdf7Abt5GsD7Qz/HibXbl+YjeNVY/99ipUeZ4JfFDAZTum
ovkVnBD7TuftbyK9W6hbtAd+ReQ3aENS42rGm3qaX9Gnz3YfjcJZlnNsbo8/T3Ku
nNzWVHCNuuW+G6qgj/NghysJx9ZMLsf7U33rdV91qfjnqfMnbhTutufdv8Xx1avc
Hj3zNjgbqEoX5v8Arlvwt+9lORjP1dNzY+aeoOvWz9qXMckAkr2u4JBXbG+PjBvA
QEFMyRFG2xRg1YPMG/BsmXYbPsolSfbwj41ok5nDwZ/MpYtqSBQ8iuuplCfcnl4m
lx4NRsnrWD+EZ2bhnBQVIzBsrU/bac24xXMNXm4lBqIwfKAADryquIxQDzCJ+XTl
MYYe9RZ00/JDYxydNS+NlWUQFcMmnzq0mf/9qDwjTSkhCUVVTTHfO9EP8SMSCIIS
mE5CDKxmSlxpQdklpPkjrXwtIA7nr8n+yqkCWbKy9hbZ0z4+bhGK9OAXMAmGYCqt
YuwdbMz7DUE7YYMcO66Rf5G2ZPMaJrGKSqbgbAfzDWIlikkaLCdT0kFiG0tfsEBG
BxsIvhvaiAmE9qTOICgtvKdM1tEvOkMOidACYhnukgi/XjRlJ/Hg+F3n5BLGEjQX
cmDANzSysW0jwzFy+L6khUxKXroj4B+PTX0U0E+K7q1QgC+EtRS3iTXLQK4RwSea
os9GeeLt6QtgifQS8pLk8yar4aVKZrjzKe8wBbw2GEWCV7w2J3J7va0VjzAKTY/N
xno4kU69cIeq56fWuLmTcf4CyJ/b5lp/XW6lTwfyZbngYp81O0q1bxWMLjmc8U5A
Wf3ymnjHLmDEnF1opWIAGi1yQlPkZwkF7kz8Ww2J+4QztIIjUkoGZL8p6wgDzkqM
ksWFuWUnFxFu0TIIovzltnwu2eo9fvbT2udVO0XXF3+HuYqr1F6271MTKuuQIafk
kC17YFq9f301wUCLcAsmI9gUkaFMi949dWWEfiDYgkM1LWQgR6LaobHiqK+34kGW
R9oCi7sfqnYimlaB4iJN+tbEhXfE7WJdH0r+qT5pWqDWlWua6qYLngMKcj6i9QoE
80p9yyFidXCwirMTZxhisbT4S5Iw7JfTKJcYGrp1JE0qsGR+EC1SfLMMMpMZ7hRv
bwYJV+cjUpYHjdMh7e2iITeNpLE0apAvjJywV/qRK5kNnspPTXJJgFh3t1XXDhWE
+GqumMhAVn7c7COQIYkorl+d9QoHjx1WBFvJPVe5Vj2pjl5Iu8zUbCZPeg20XQa6
7CcftUp2aCMsQIUSK5YAp4fIf1iFwGSIVp7ILwT/07MyiToLnO7U171w4dRkqJ98
IFXq1OujYFrsRzhPHxqszgNoanVA0eB30c0X94PuZlMVI3WkzMu+S1y5TOyKXGfv
5hOcLHWRw30H9rRh5NuqvtSmmMt1Ogp8rEIJjfsHbiCYH7pnz5Yw3gyF2xy9cqG0
RGTABBRLBNn2ey9KYrXU53z12yNF3fOEAxRRHmsVcugSYCKXH3ND/qbAum8Dq+f5
XL4DXFuWLMDl+kzznxqe+fLMjLoAKj/5pn9w8qzjPxnI4S+fkbphS9IBiNS6vDld
TKMg6bgs/KnpuKQIxWN6p+ixCU3JvVRCpxdiIEztvaVNW4xORXfV1o2FV4HGO6Cq
0zpT/vWE5OP/inZL0C9nSZJWfzEffNDwPVnBLJNtxNpFK1VhtN1RxVFb5o72r1Hj
Yd7gA742mhI7bmsJuyeDspiX2yEURTIg14PFmsmiqCvXqn80CxuyXM55WQsYXgx1
NCSddPg0tqFKis/UM3/G5KVyCtT/sD8UGfLNtxK84SKxKAiV19+u/yZpOzp8JAb2
fe2YhKflI32XqW4j/Yoihz7zS95oSNQoMk9dQeTqMzI9iI0oI7+zFTYIkwP5zLnu
NKCOfqnCxiSerJhk5NuYZbHbkgHDTKfZ1piB0i+LDH7bsi5f9ScJA/DQ0IoIM4Wx
0vi1HBF4dMXz8eA31VlGMkACtFHYyfPffOr2vSyLlr9eIZORcMauJOMjIUlqp42i
PcXV7Jbqlyl0K1QygEp+ZAIS4lHSqlq2E8DHD7ByrhitjECkJMedKmWzipbVed6C
NJ1axwkMqr+7qrRAd10/2fA+12q7KXNPOkFSN/4lGj/Mc0JVLhdEpN35hBt7rxW2
pQVwMvEIR7Bid3z/HyS600vmOGbjHr48jIULW4W1ViwwxwpwpLY2KbsRrUyB1gxl
3fyEoqi+IBfO4AIYTqbVxl0uINkNvSaXr5ZoGMzD6y9ltqQ8L1eNwGkgItQ/S/x6
sU55tZzr1HNB/NciEjn8ME7U//2LixVIkLybdjwYVFq0oFMqtAOvp9vLsfnGYGOQ
rIrqXNt9mzHZk6BE7J4HN1GeRKNEIjv/jPi5fMJZEx5h4tx5kmPfIqZiUka+xtpL
mtBNAx/ImIYAMhOJiYTbbWaSFsh7hVHmYB2B/NoEtPzMVOUZrH0r3xCy69U8Uyst
M46k93InYGzEwZ7g8EpliNp8hkpQ6hKzYoK91YNSWEvppOMYp5lVEvi9NOzdT/QA
8XTMtPC7iNEiZ7Z2kGy+lcYKOBHm/2xFPIkfSaqX5Eo8F2iKPTG++NQb9RjpZW8k
85MK8DzuktCh3uaPdMytif/j5Cv+Ko4eYTDdT1jaXFvaRHSJp5Aq4Y90S8N/jXBG
F+1BMxbpxNiNOyTPxSsc3Y0Jj79XsnJ81TlUBpzCeWO8rXBCcn2m9WqaamtrU7W0
pjEkpokta6ujerqYnzr7mjz0xt6BZMoZIUbBEvVDMZJ8eq2BviI4r3wtO+6T6Qrm
D9IKksgEv/bQtXCBVsH23S2P20JDUOhXbqUMQ5A7QAH7HNeUsyadv/SLnTZuX9AI
wAcsp77DVoxRRavHP7dzclvU/7v5i+UTG+/WGKYPHEfxQeLzMSUBB/EKpmKz9GoU
mS7XJ4Jq1eDWrSNzfX3FPmNdlq9Qu49KZ7yV8qmZbRsB8PWB6BRXiBwayaa3Nt6U
X6QWlRZciH1dPeRecXF6pKJ5+9mok9ch6aaS+h5BqUcgxcm4R1ec96lXAP3pjAIb
intOlHbaNKofTf6fUX3aHGGPCqXxzzm7dNhrhHPz6+msgvBXQZvEYNY0NVJM45Mx
seTEAAvkb6PqwrqLCYaHg2wLogrRwBzp5SO2bbMpGCHKBbUBwjs24pG7i9RPqb2E
rISnfEPmTTvbGSsB0k5g7gfHyMJb8BG0FP+p7GQT745q1DjaYOGwlW3XCUuBWyo0
6QLL8cUVNoyIBVhMTZzcFNUFZed6ADs/O5G5IoCAWRbJu11Q0hP+5fTiM6R2KnUP
bQIY/mRO0ef50bS/cXO56wrp/yuZaPs2ncN2UCia8xYL4yZb9itp5eNFurxnketQ
E7esUbM03mQdgVXiE2I38rYdEQDMABMUDdsjDADoN9+tlpgM5ampmzTzP7wY9Uj7
Ujgcbg+bVLjiKk7mjv6fX0TZexd1XtZOHAJQuV/ktv4UTQ3Ca5aKCc8SyTGF80mN
TJAr6Bw3Sz1in18Sald+xh7/kq2GAe3iEaSSUZVO2t65b9s5js5M+wx5sXuN6o5z
MuO2lCvg0ASsDKHLjdSNmGrELc0ynjymiuxc/BZS/0Z7tJaExIruMLDxg120Hu2U
D+Zs0tBL28Z5WUoFD1UC9uJak1w0Vy+DMW14zOPTXqvEy39z8UVd2cswuDaUpIgn
xi9SJdSM4EqQNidVXTL2FXsa17hlyEb1tobTfAaAvqcyVTz1JWU7wYt4i41dDYpN
+CJMk816F0Uumu0WOy8ZYPd21+QXa/eC0OL2ZL1vS38OKaBy5a53p8TyrOr+S4Jn
yspTzboI1bJMe570Gck9kkn7/rtxL54qceGm7uzhE+tKbKgkM/cdTc20+gRTbsR4
vm9N6BR3zqudCBleee83z8AiEmbQN+fcWal58PqfL6iZOWG5E6ilF3QkgnaeRsZB
DUC/FdAUHg4N1PiJ8aDmzyQ7JMURr3m8+7AN7prHmIeEPhpC7MqG4y7gI8zmfvPl
E6ofGxATuAus2v1NC5fe9bS00go952pNhry+EOB57ESJKzU1eWEpLi2CRbOdA8cQ
TQLBvNi2f2pDP2h/0QJbUWzma4ICv9QggU4BikrzoJWHCcAcmtdlKNThGg8fav0i
rH/g2YJIES/m8KtVSgueMFSciPlf/W8RJXy+43//hR3MPw3mGQmcx8dY1NJavkoZ
3zQfzCEDpxKqpfbGFVEbpQ7RedV9NWV6ezHQDBEanqJMzBow5+HM0J9Smw1aPRG/
eHhpO0PzI8T/w4j4srH09u7FU2leOP05XfpHA4h52gkV7d2/Sj2S2iSyqWfu614n
QEsdoiHqLzcM/cjrGtqzK2Z3Xs2smSknurxCya5plDROgssuEoNxzLAl1+6I6j3h
KhhB/5469NjskNv0ADGn+D/UXpp5aHuKRMBiho8F4MQqROZKGATo7+fUb+GmL785
1KnyEChCM2o56LG5baE3LkajnYqgp2Vbnnh76hh6ejIPuhOOTeol9oi7GunXyBpG
KNXum2OofIglDWMGrcCA1pOSRs8ufARBJs2KqlNvJ2aVDI8sGhL2ITuYnNT9MepA
riUsBBYh9Ed+HX7wRJOpFEKZoxxZbnG400GWXJGa3/d+6mocAZe4xeTYy3Iwxjrd
U536hWEZ4R13hYFNuK4F1/zLdTGrqXGy8ECyC9q5DC0rv58ACq4bm+Ac//7iIFDH
iUYKN1KgVZRJlVOtClkP/Qz0XGTGn5s6FzoIme9r6ZwwZY/gXPdJdheAbP8A3QFI
zbPdutnkhdQIXmfZRTBJW2838aWJgT9EHslWLUm86U0n+ge+qz5Qywejaq3tzjgC
oRO44d430xfX5g/bKovO0Jywjkh10Zdw9NI7TutGXUADDdS7G0cuiSLt5FWcsGcn
1NwpyR9Onqzu/KubiHPhUEX3brQSpMhs1j5lRk/oDMWLjErni8rdN6xavtx6RCkL
sULreEII+7nG5QeW9DCJDlGJrwmk3Ts3jjSfWdqWfygcMCeaiuSAJu2X93eNqMcR
WeVBrxjH4yJ6FCYNo9bY1nCLxAhD7OILJ4brDoaXDJQpuqc1VASNHtU0V44Pky2a
wIbqAyKZBP55HIysGcosa8joYFouQfkSs+q1DHEjCSLdkdLz2EvaQZOqEUVPdx4t
huWgwvn11yRH9EbZXh6UsToX6OM8o/A7ENLLCqb6Gv4RlLGtLVoSicSd7clsZJbm
o6dslJkc3wO+FKANT4SYQG8sdWxtecBwMdIIkldpg7LpZpM/YUxZa5FRo6CXYy3f
LHUsqVMMRP1YVn8KAdIBqeuWqH4fw7k02KQbEAjiOq6/e4DKcwJoM7MA6+8A5T3j
krEq3SZlFhDJT82nByZRsruKSCno87T6/FnNMuWv9RItSYeaHS0z7Q9cgCxA9n1n
VwOeBvz+BhK3GJ/nCYbMJddZB9SS8dS96arb39rJcqkpzyVHMXZ8egaCGau1lLt/
zyJWK6BrTYJ1zpdK66KN5qmfE9zLxasMgji2OUqrREdG3lk9XmtUxXLvX/hqh3nO
8vujrvpwnD7Vcsz+eYnM8TTLoCcvPFxFfOvlnWy6Ev7+09+YErtkpaCu0h5Ckq18
Wm52hTQCk9RsqGuix/SHBqz+VfX8o7u3eSxUDgCo0u5OCByJWqOOoQf8GSTQp6Tv
DzaTJ8SRbvnU8dkoPBGCQid0gZgB3dlw6Y1O/zB28Xuqorxo13FMM0nh0vMKiRAa
JE9mbtTVEtmN79NJD5PboINk3xCqYvHInajLE7p8t3kSAYeQphg/Vy4lvb80MlGv
daDZneHulkQeZ29o/zKM2lbqyQn9CJg8MJ9nf1vcSUvLNG0oCvbNQNH4bzIfJIlI
rq0PfBZCwOa2kpi3f8Scr2W8EtB3XZli7al1kN+ZndH9dR35IJlWBSwJfBstR2jm
p6zhjUD5zwOOTIv7f//pyiln5KqAoNwXxloeCSPv7KPwHH5rtB+2pBDf5lqcvGQV
3ACTG2nE41NjUwEl3udNIvKobvHg7eZc/Ry6rR9defxWbX1UIbTmwv9WzPT8URAc
4/dWGf+uv/cM+jKu+2vnsYKB+dO8RibGrss3iZLy2Eqk3Hrosvzvsmzu4k1fTBs6
NGXFqU5MkuJqbqAVmHuRKz1wuegkU6sZdCNtqttCqDPBUuvUndkp8TZNBuVk83lK
e2Duebr3/JefNm8wdYlzLjXHLMP1qikootoJ5jcyjhF09jpbA1uuiAvLtfBhRunz
4fIr3D/iW503YqJ040ARvUiSpdTMLtrWa5JEE5okU62qjSSChv2Idaf+dT/ShNBw
PuLIqd2qvOWPI+eyrYHuIrIKWla+xtJV1IoMB6JvL98ey361UXXOWys/9nbQg70f
L64rI8YM07KlfvkIHk12omD0FVIiphNhvzSt/k60gAV3sG8YWvptEogSOdDwxT3K
+bTenCWDMQoiI5cqYQ1dulv1s9RmQf8Vw2MIp1lL18Nz0DOomn8Un6Nng1bo16OQ
Ckj7Nb026GjOFq252KpIA4lC7aYxhubYiQKMCD0Ok8EyqvrJ88GN4dj0P4A6bUlY
JW/UMNLfXI1+ufz6Qg3DP3n/FUnPWqr2mHHhgCoda16flFv1M6LIj+jyLgHY2H9o
2LaNy38mmwVyWt/9miCuqXOobURQOatNSta9hUWlWn89Svrz1eV9D7UxrCRB/FGn
mY+P736ymvtqSpmG9zKk8kwPLuiBK6sa2io2yhLh0QzEIzAg4GawASS4ci/6h9pu
HLkRXLYpEQ6hTUpNqCoskX7KcU2zC+5WZ8rvr3RLpZDU/AYrRQLON6zdFbas56mF
8Xz+Zeq86q7w7pxASQyqzHtHMaq15oQFdL5E4xHExAXhMR0D8YiJZnu3INmi1q1f
jW0KeWbiZUsCaw+6+6l9GCjzNHjw/BioBMZB3Jcbynv30p8bLG/M6EYL3Xc7u2sx
WsqhpYXRegdkb2LOJmQGis2/i0uwUZA5LBnzCOezfJghO1ljvvZ3aMiC5YXll3gL
xAQNfbOsNSXcz/5mfPa9a4QfFKKIlohxFglKHpC1ylEqAUEHWK5y3yprxwWU1h2Z
7UZ7ojgLJYS7eXy1zOQEOG2cfVbLADjQzehegO2N19O8oz/rlUPXN0z0TGwzsMv+
49wfRBKWIPhZgnO9M1ykIHH69Pfw8duiHGMPQ4uYrzGYihtT0KYe0w5nYYO3pRGr
/8XbmrxjMVrCgJza7OTTSrnWhWD0TekAHXZ2FQkhgPEqAaT1oBj7XUdT/jPp5KuE
ZXQ4k8fGF+zTFr3P+RuQeDS3UIGDT+DQ2DBd9HNPWA87MhDAH943kcvv6jRsnzj3
1vDLXblsv2YduGmJsfnY8cGjHvHG2zNz3YVD9VDuVJDZ9MdLY5S8UKmHpXYN/cCR
ifL/xvjoufhCR4LotFwu3w892oe75S3zs9cqsbamko4g0nIainnOF7TR4gnD8pYp
uVNoCPW+vhve3aJABjFKiCmwGytsrmWqI/mPhScNsSgZc3dCX/2UaipUHMxA6N1B
oq4VB4jEpMsYDYq5x0M5X/uafLU/+1Hsk151eGDMdz/9kF0kxEqAA1eG1VS/XA2H
lUTpNtbwVWo+0YgBVFUjs/kAUcfnzJnFtNUJJ9zX39u7W2i69N76FNYRNTnweNIS
NhZTS7m7u0/HEKQORahwNIeUwGUz5QwQDx7wT9s978mp7rEjmpKqTqSrbM6ajmJw
dHTqdt+QTUvhg/UL9q/3UvOevjiQrxzJtFFMIweZGxYhjQ7T5oljcF3m8ciqewWP
vqHh8BnutW9fr3cq+L8ZumlCDiKG/ULacBxLf6Bo2PoDECs/l7v6zQmzWnRVykhG
HaWcE1/s+bo4iRO/2ejSjvKdkA6x3Lwj2SWt9tNhCxzaVirsieAh6gkNQwNurszx
kfIzfQL3b9/9yoHmsfANKcrZkoJ5K37RScuGshlU5wHSkgJfiDuyL2CKgYtQy3I3
Y2dg0alBCM3PSDBpn4M9NSThSgT7XOYSh9QJg18vB1w43W5aXU8b0HNFi+l4wmbM
BL1AleMY4qAKFzQHFCALCKFtt9aS9ndXks8GfPXnJXOech2SP+LxOdppe4udFEHn
vwl8HDodyogwq8UlpfHon2gF+ke+lI9yxm7v7jsYtDIch2d8+rAZaWA4DLoPUNzq
NNkJAa0T45dUdH7d6RWSi+IKn+DDnd/bVhqWdDlmfms4sTZ4JtBGr9OHIzaaTeZ0
wJ1Mgd50ZsxMsVDKxzbUa4tlh52jiBcjgfPUIynWrFCiJiFjFK9lKOCMRYtyTl0a
dAmFffQiOYlw7fP2rix0a54PXOsPB1bVNbRZAMYC0K3nW4OKqPUjAfs4Dg0lNUlV
OHJDO/glSXoB0CAPkxncWwHcb1QGuNstbSH3rP8R1UA9cdQO1X8ZLxa1kl2KlKf+
0EOHrZE9Ph0eqsd7uqQdfKdJDqGL5AGJYz6Q6VDTBvN6VoUTookljCz74XBUYU+8
SoIcGy+hhcbPbCeGBijAw2NGGPwhKMxUavhMJQu5b5Lh2AWKc9E4QFhZPPIVoi0V
eRjASRaT4gN9v4e2WcWFi309qXDe0P7uyDpAo4iSxNpXC5hq7Qa+YwgJiEdr0yzi
uqAspiHN4On1nUaF+te8Jqu8wUpp+jjNkBqRYF6FvTVa6x5Yi1SQq43ieOXa/VCu
wS3vCELaMD5Ak6IvvbfSr1CeAp5zELjT+GVHDSo3Zap/h6/stsSCPRcPU8ft7BwX
6eygPzhPjHbCdnV84XlmLEUKcf3GuDZzv3/lODIuqr1Q6f3qTCrZTFWu9Wvzb7kE
o4PqQgsGSL4x7wHz9QPuwleNhTOlRsJzx3vwLqXGuc17lfEiu+kbKyBK677nKVHD
ybRdfRYJ/1nwfZNumbqZMqZSq1TdSzUdEerN82dwWIqcQgOYtbPgz+F/wpZJgh/G
J5yQ5PWjAFcEly69E0gpA0gOkNFjVZX05TsQF32h3Kj7T0B4DSiMpL8pQ9EbA8BQ
eM2NOjh9JaVYrLqG0uCoF69IQy+pa0RKpUxPqJbxuVR0bR+scJ/lrp74no1ryeOL
44MnAPiwE8qZOz0VaSlCasjCcfU2o5oiDrExt/CUBatHvidc0DyUEI9xjGXPbRzV
u/Wmh/ef2X+4QMu6TLSOKdyXI562aJSBWPoSe9FculTjJhEwMxbi2mM47LFj8TJZ
ADBD8WJB8RJtHKcB/AD8IjDUKPPMSZgxn0GEC8cnI54BDYw4pcUv+pp79TDZjYa4
+taeoPP407xAx61rbDVbAF7STHuALYqrtRM4JQFqOidhs7Gq8oCzD8SBD0rHddev
+TUqi7heZoK2q8sXAp0ThMojuJ0dAWVn3PVcajaaD0YRI267JqxAloOPFErPbWs9
af5W2X4gRM6rruUW6t1fbrN8cd4RTOclK7DXaDSQ1W1nSwcsvB47VhfE2HxfNGXw
j4/g48Us3yqOiG/tBCNbTF1AVh+P2sje8lizpp/IbjdEAV6T8brNMsoH5U28NIht
R9k97mjzQst2SjWxbKY+aduedghr/VNN3JUomqPNkd6ZpFikEU5b1zSLi96YhT/K
WoJLlpRI9e4fHgyt+LPMbVvCgUAK/NujHHXOUvrHcJevR5JJuvcFP3GwnfFepSW4
c+u4jazmuE1rDwXiRmXIG2nKPNIxrnXN0JS7bykAfQThFAu04AmyCxj5qX7nCfUi
Tlv5CfgbxhLTOhKaGp5sW+HMPTiY8NjKVep7aRMKUKh9s3U+njXWsPXp6VhTaba2
b4W6vLAy3X6FCtqhMbSrKlPwBh9xepT6RyFn09StyjI2bdIwKvl9dLwOrEELlReq
g4+oWsBDmeQMgyx60bjHp4f/YC/GU3qLJqhlknCjaIWpWzM8efpHmcjC7vuMhtiC
Llk18JnYvCMlSRHrDCZUb2/6wmuCgjTnMgZ84DI/ZwxB0FFyvVRfIBp/pq6/9XZ+
GxAvyelrWSidzA/bTumX/UnkMyP9gPJnbQWJlF2L26u56zusaQxfI6OkeLX0dZZG
Lg9vhRBIO4xzFyD1CERVfTW7euZ7VldxaCuAsBxks40jurLK3fwYWfQlRm2tRpiN
oCYyU9fs225I7OBR1SVagr9Xnb+jfWi1uLXWQyVyuxr/vnTaApMR88JX7Pj7sZTp
CKaYyz9ZcT6bVuXX5hEa6VOcITsL8xbHGLEeeSOkYiztoXe95JUHAl2X4yTGzD3R
DRjVOTZADzB2sHGSazRQRSvPz56zBT2HajZd6iLtzn7o4JnKZ35NQeoDuaaBwl6z
p47Nu0adOiKhk53bREMMyl5jhv+Q3k1h5Lg3rPMMiJyt8TIPEa06qL2CjDuzfAPE
PkdSp5mnoUgxvjaOPdZjOq9YYjpOYmtRbe1kB1LOZZ7+f2/vveIydgN+1868Yzu4
KpDO6YSf7yZTICbaGq9N4E1mbWfyqF7DBFACYjyb6J0lUykDeflVIMllRzn+5btW
UVuxsRTLcAclcLoEOeTKka/5DC1OaW95o+oTG4QCxnXzHfzN4E4vaUFhpFF9klSk
LPXjr/yCJB7df9NBDodln2+ZhZH0tzHOlWFy7yPBGB7/ar5YF+vU/S9snAx4hbNT
a092m80B09sbH1p+C7z0lvwN69OCov6mI3WwAyuuG8p8hiUUInHOfNS9szZ0pcXT
JOe3NrKRzN0hpAW0/1MlZfYcvrljxFuTnGUk+UpgkbtViqgk6CdMWbYTre+3VOi2
8wIp3g7NEgvorPtMr86ofQjxcCHFa8cSFPudTh3mDSJQE+bitSFA8Ch0MXkV8Dz0
JhXuuTcrda96T2q2tmHonrHXVVc8obUzoJM7kfLIzV7278sJnWLC6LB5FpVP3bjd
lRyfWx3yeCf/g3E3nihN42hUvrF/KU389SKr1BYGdPUf96NCid6vi9FAvPLqif1k
noGQagOAQdY2vBcNzEzXrGuZqLCNj13Ii7lujAh53eYR7ihGkeuwel+Bzmj4TV3H
WqGxqcmFKE8ahPAd8dGCCZXmB5IUBAp05NKHYAa5TSbiZRfb+z8T/cldy5e8OY58
ZL6PdH/FkrvGueOsXE5FnKpy+Sly1/661h6pBPQgveZ/3boSkV2vSmxvPO2k46i9
ucIZa2kEwTKlzePj+i888eFTN6gJdPnZFZZHFXCOboim0zt44pYYBrPVYHmF6clo
hqu23IVOlUjuPGchHdKsbaq0BFyf24Io3wMn2ENVGXWaAVFTKniPa8Qmugp250yG
sA496IFp28twTkHHxdKkjUvubN78lUEdL3frqkZtgE9xoz1qtpH7xnOfOK+L6LhE
AmqlqWKLULOMS0pE1e1deESS7bIWIGWsLr0VkokSWF1l9m74s/Qmnf8E4BDyzAFF
eS/Xz5B2gf4N806lxxxN4ktCJV0ZFUrAC6odjog+LpPj8GT9OhgV77P0dUqksErV
/xxmJOlf25iK7Hnoq5C7D00JxQCdPwf3yQaFFJzhW46B0ATEMgIPTzlGl62m0ojP
E9MmRlobeUtlWtONQzhVMUeO5IBfCDGI7HEc1l/PxnAyLxtyPYpdPn6q/FmzRYvW
xoSGn38p1brquLuIjmnjrDTrlIPTwIXvMlV8194GJTqLisq1gzAEaCD7mle6wQXd
8Z1xWwwq+XdukqeJK1VWh/mMQxp+76tHjisr8ENx8vfpygYyPK5oQHSDeIXPoMng
yGM3mG6T+xXdInCcuH4d23Zq/dzlmagV2OcwMpQHuZgnYxdIxvzdd5LZKYFz1DR+
+jDHgxEKtLIY96UXMXAizqoypLSvZhsRB+qSaZb31bqG09H2HAVu0dHfihKcJlqR
UbpMaaut+G6zNSn/3CHt0AjvVSft9Faxd9sAVxCs/yjxR/weIgzRnh1cD6uxF/lC
cn8EwM4EP5PaZoa3xHvPY0UV9pi12Abg0cVTL6ZfuaoXhT9H5s2SE8uwqB97LowD
WMFTsJApeFNzmayb6ak058GDv4kMJ8fMpiBXnOXV/aFAB5pbcRtbtiVLFvuAbLWn
U3gqtB3QBzQEJyM9tAnHlqWDn9kgJWtCgW9Eixc2D6FT9NRuvCnzm+wR0baXLvZX
GlNAtWnzGHIGQsdSUs6TISpzsHWhos7xOFe3k1Oe5S7bJSzt3KfMJKpLhyN3QQGt
771VW7yOs5D5ZGyiZ79s2XkUvSUQNfBFTF9bjDALtiICpjZ7UkYRXpZwhcCMJbsF
IfG4P7v54RqINc0iPQd8eXYNy1sBfumtB5KV8KXE5JL+oHffsq8yDAMPO1pqfqTH
FRqpdwrvnh4k0LAP8et10LAk16ZC5aHmqXMQF9Zto5LEGTqUrTU7gmtW8vPcRSwZ
C5Ed/o2DB1v4RdywMkQ6KJYuADiQdY68DTrQuIY762/KoPmkkgy0k6pjktWtgBXV
pv5xh+zanMzwvZAwr51g5uB7md0ZiBAvOTf3wY8U7oVo1eJgiXRliWRjW/zrsHA0
d/FT5avoVgFoAyETUGusJd0bhOCAk2PC/clsaTu03Hoi28h+foFjLJHmJ/B/qpn9
lZyt6ZElkr5jWdGuIEK0GcdfdxNknepqxgjFUo0gVN7vQbDvniQf8F2Gjiln77x4
PHftwDloVGn6zIaHlBj0JNBTgHdRL81XaeWbjHIillBHXTprWoEtqYvPlUrqKA1N
ytsuEw7ZLV0pJIuXYuMUiowEo2SQmxKvvmeWumytGzLPV2AzS4891qptyuN/z3e2
FOEokEh2aWGTnzXARDuPU5ITMWdgZ2DLW5tH4HzZloFlTgT3NymicN0QZk7y6yY1
dQCmZlWkLUSfmj9ASW8ZRdEinlutcciClwoBj5ffBYksT8ww9tj0I3iuVK9dMCkH
yy93Y9CYWxn5Gy2N4TsyFsMHgAzs6dAUIazNr52h2ZfhdemSCHxPbYXcwpjzSSbd
jm8YlyBRzNjhLfNW6cna7Fpyme+1Vcla3LfHn0ooU7pFsqAvf/wE+cLA46QTVA0K
gukJARnpfk166IDqu2hVHqiXjc7YbV+NLN7SznK2UOQUoXpcw0eV0vNVeEZ17XGP
x1DhQgP8jSyDfem5/5ftAB9ahpdhNbUKM/JM3jcDDKfLJbXcZd2P4X4C40nYbcLM
06W7+abd30xrCJsjEBeQ60dFhGr1OpmpMzFatw6R40xrlZGfAe1cp66A97M7HiO7
egbm7SddNhRzXcNhayseiW4CiIFL4IPnaS6HvdLbojkJS4M8lojBXja+iizAwVM1
httWUgdpgHvn8TGgVn3/kC+8RNu57DKANERW8dD53Zes8CR8IgDU5eHBcXW9VWjN
2wYkDBi1UM/OGs/QG8dqc49lIFXOfK3gUQK+Kyty7v2Ranx3Odc20tYymQHluWy4
CV3nBxb2kA/G0aICZP3k9oO62ZxE847WJeJRmsBxeFfZiaI3AfO9a2oH7fEHxVDY
E3oBdpMjrABh6dZHig6tS9LpHdgFGY4cYJo8Y/4DaLZj+i9Elu5KXPAw9hA7Zk1f
5E7pZAZ3eUbMgCe+7tiQRCEArUXGILQoPcWYZaUdJFLeNHBdhEVt/w2RZODiIWqe
zs1ngZRSzqpYNEoHo27JgPxTiHm8GqaMG7ELfzrGG2F+zYQob4xza53qmR8qgfw3
e6u6IKQli0fOa97gjwqMSMYFj6bC+wIikxvPJCZDHwSFKk+YJQSmqTRMR+7ZZddE
WuAoTCGO+A6BKsguH49727fMIH1s2d+WQFwxh4GN/a2q3rkDP7URjRawwqgoxLUK
tdn/YZ9WanKO33pa7mrf0wSbAek1sxJTKyOglCdrYSxEpI0vnl6s85k9e1K0/3Xz
yxXK5vCtHB/V9yrRDmeqQXla2PZWlZYUTQNlqTHhsCC/rAjfbyQEYGy4UG1lgKGl
eMiRK5D3wSMUaufYZWogtitrWKESV9mEifGKP328CsCy7NcO/DHMlll6gdsGffqg
JAC8gBP40aEl7GtxZWV91+XbuIxQWxzkI5euhKrCIqa0osihG66ToYZLkmP+oYUq
OKUw44++TuL7X8YVWGQD8bSwgXG0iUyTT1uDxERGC8Up8bShmpwxvRwfF87JYyIH
e5n9jvgC1clm+orCCgo+H04FqEEU503a6HtMMDK+aaXZMLeHlXLU5MYNnEEl7N31
50i91ahCqf+5KWpRt2F5Ly+nS/7y5Zl8hu3ZkSFVXLKnuatY/Jv1goqRM28gCQYe
/9WleaUuutmHqU2FTg8rV+4HjSnIIcCFW2Hw6offR3avfqFyRCwDIGyMVYWjT9rV
kUcqr9yqhXLs0ZxFULBMYbEKDB+MvutPavKm24jbJG5hW/fkydfHT4UQfwFgLUV6
FWWqZPdCC8YAeLSBEwW3itC7vNDrWuuUOY2dzEiDcGDEThLbRzzYU530CdZack3k
AF2Bpl+3LJRtJkX+xtjHn+Olg4qCOdg/O6BxaAR74bDlVIwIK/MnoumObNkaNWMW
V49EJGVrDLf5lYx5YW/Cw0meuERuQdW0qWpIr7PaNBXG9affKMvFUkQOcau9YooW
0GCgu+ZPawmuHXYCGoJJyIDMetqd5bnt8why3SV5xEsnpl+QsaOu4V4sj59PRVTX
d6fmHQ9yIG8Zxp33YEbYdBBsN7aGPkTxw5ZyhoiNzFUAdOvRjs+4A7RbF/3bOVG5
QOy6w4uP7DZWt0BiXgJPoClQzdQdYcqi7F6JZPNjgHXQrc85bgu32zcd4jaRMSdn
xl6km51p/GV/fzL3MrEeECH13Lmw9YQZfR577cJdNRHqZj3vF+1n1FgyZ79vElKy
tXb0jX8mrhK3wPetcfYinbOUeUsm6d6k25gXus6F7r+f+5Uo0koMwek6HaMDLSRf
KAcAiVcmatr13ipKifPczATEpw47UEOqOusIRT4T1OXbAqt+YoDw9mPAxoISEDQo
laXDA0Ijpab5zO1XROYOGPQLPJ/09TUdEAqb8CT5OrJL9QhcOAFv9XSQKYBImLq3
7g/ue5Q9Mmcd5+e3F10xljuw3uG4TIrCV8LUR63Xh0R2uXPav1AObd0p3AzCiXmm
ybY+vy6XDQn5XlhtpdrxW+5DF2ezjOpAQ8T15oPU4njuD6ciauFMRdqcc4ZeXSWu
TaJwVVRnkn61Z6sU/ntKB3kJZp2O5zdBGIOOPmyBqDylXO4QjbcxVdaBrCChrCSa
8RQmZ9O6p78SnanlBsw/IsAf6OKS7F2VB2YTFM7vcteB78biJrgsfiT4jWpWU8FW
8YxdZR9xHHDOLcZBhAtPo7GOMxMw3Bn+kWe2xKXAPhydyLx1R7/8o9ZLQt1EpndT
ySFoMKcFZDqb7KNlpJIHzKyDZkUkFZq2+nVFS7hUolpCLTbrn5ETyAjUjKtaL9bO
oXEVbiM/izJYs02i3FCVCGUxLdBBBTCqYOlMrlE+4vH/bpGFelIiPYOOZKlIkxwh
jOkWoHyR+AZhO3KYF6V79lftMwGzV3J5cvmFuL79XdNxr1yj92YJ8KDO/iJFYxkb
0Xfk/NVZvclkiJ8tRGN8uh4OCiaD/xZ39kdCgousY+h5s5NzOCaV03zJiUwmFW0R
aVhxzqxofQ/JP3rKTXI1JW9l8sDp8yvU8T9zUBP2TxRBW/dvOtsyv2pYyF9a0jBc
rc2T1ViNyDQb23UMiNtqPPVELPeHgLqdQOfCnSTPvwGyeS/aedWqLkfh7deQNgtm
Nr4PzjLgzYg6xrRl5ZNPAXvZDy3DSJihTXwjQSoXTFz6jq24Oo4giy3R/t6BYB+E
3OMw0jn3FDVc4orf+fb4D79Yz950Bync5lMBwZp7w2dqNQ1jkRnbMoOVEdDVTsC/
p4eFB1Uqzzlyo8pZr3bawnwvRPIQyiQ+v0c+AotqU27296OyUQxtaCn20dBX42Ms
fePoFCUdWxQKkjjt356LCltWX/afq7ohg3p7j5m4CvJ+kqDZKVuluv+Z64BLqNbq
X065uCBOBbctZqLyqWV4rStJ4Odp6Ulhsf8PexiWRA+HLdvcKZCk4ysqDOWvQX4K
Hs/hyAutA7oAa1pGDvoThfpsNFKiVUyoLzmP5Q1IBK++aMjU58OFqgV0l0pDSqsB
MS6URv4zSCjiJgOg1+ScpUhls7EYgzJI88UlGm9u+2Jbjh5QGq7qHnd3nBfyt4qm
WTjwM5AZhWfaXymnB0Zmt9/L9BH5A5mlDmy13cEqlHkyYUeSZC/nNRUtv7GgyjGf
0csgVF+MwFVSlLz1nMPk/Z5Fk+W0m6osJ1ANyfZMDb6R7h55rpu0I1iIOmB0rSc/
EU1aDUbgrmplV8D7uiTV4wOsNj6RRSuoC1Z2uOaQhCWryKJB3rnfBAlKqV7NUEwp
pRBz3EseG/tlq24I8krl2s487ZeAufM4fi1FkrlVFNwu1qWCaKE3lBoF5kS1PixS
Ti2QoZW2TdDcLrWdSBfNxA3yHpi88je25/heR2JMlZPKjZiB8hyzb+y+AzS6jhmp
ULbG4q/WUgos/RULItuwBO/CxZWmtJ2s6e6cP4RyJt+iHg+3/MCuyQvbJScng5mE
RhDAL8wX0SX9DzEet27u0Z1plbojRP1PNcPGPRWdg3k/OWiMMKePGA11caxRhL2l
pceeiRpYHavVVfmn7aEdlTGSo9lY17yF8kVOWSbtNQXaXIFSIJ65Xq0aP4RK/MQ7
jg9geB6qKfX8K6aHXkgBUSavMoaZ8xTqkPiM1bHPIv0LTi2MAl9X+vDKE+8vP6Ja
wvMktsGAbvkfMsB6vOA3fEWSBwGzogf/94xfqy71qGIJIpb9PwPBliex/nensOL+
VdDIs42/ZVKZJNjWDkzA15WPuJEFtw8bGNnyy3cnFSlvRrit3IhRV86PaQVNW+OX
EWjQIjDgq2NgTlZwaCI21nww7z3UceHlbFZsj+uxtRVq1Du03Qybn4t+h+8oH07J
Tkm5tecndU/Z4f3m6+AxFPQ1hCUeUArIR22cKvr1UP4fddc9Z003idGf5H8tTZ45
r99MchqWEEyPALU3WRsDEJM4CxmqeKovau3rTgRZPwC6iSmJR8/c+VMAjA3IDI5c
Fv4HXyeDqatO6Hcirgk/Yi2rAW9g9aeDNNZCHEsahLiVK9+mHI7hkAUOEY+EnkIn
Mr4D24u9IpDXWVfzw0eMIKpsiJgEO+JhiSJK2uVhlJx227IJeQu4lt23dbx49c+E
/W6lbB33wdTao4h17dXcQHG125YfBrpmuPyPiG9tt8OetOrf5gGK/kfs4Xp4Vvea
uINeb9xp8HNUV468Z0j26COsXSTrJG/mi29525u/Cx4pPtntNPLOKNd3NBH3z2zw
SVZc3y4Rtai8rx6i93CoP7dGMdzKhCWzi+zzuzrxug7h3KFQdFd1gQ/9ujN7e87A
AltgOuMLikR9QOvKHgEFLcVABUn+VKizHm5rNwzD5L8UKIeHiM6BofjYgzunCdIS
9LOHt5oBUObP09EkY+D+RQtEsL7Oj2yVh5iNf/3TNYMHOzE1FfDYgOWDg1YJXNC4
3Tpv+3BQdXhS1k1bLm2sYAWB85V7Y0JCXC/YoSbysuybz20vusMGKNaTZ00+jMdy
teWaIn+Or8tFqCqy4F8W/S+y6WrsQmuUFup104DE46RLfFgw9lutQo9BNC7bDZS9
rFheXAYk8ejbDLk/srU5My+YBCWtUwdinDisAJmzyI8+pYbY8yASBMOwRGkfBVvj
c/eNN/3/db60tqHidTJZv+KR7IrnVDdcSDiF+JPMHH6ay16HP9XS9GCzOX7UEaPb
ogh9dDWKVGR46B/8VAOtjJCSTlexGORbW+8gh/eolf7qPF7kI70wvDTAZA7IfK1f
soL78mUJcI/MmxsiyXFJEo3Sf1Y1pFFykOjRCUSn2w+RcwkMdKTdvv8emEcPN72+
6TNTDY0b3SsTYpbfWLsW1DYVQNHYHCJIy59oqVAuTYYLuCm8PC+4HN/AMtlc8Gdc
MxXlfso+S+obX2GigDMoV0qo/pGeVxN1rpKMFQ1YJfVUnSBpVXYD4yQZePxrHWbM
7JLh/QFmvnZwR4frUMGcZzJGosvlJVW29oG6+2nfsjEFUTu0Gvf52nxhUKG1/YlJ
6LexkXfQ5oSrGGvPrsGNG/9Mj+wBU3JcZ4swl7ggI3LTRdd087ug5AosMOruXanG
6ObaIF2Si7MWFz6k4XaNF/gF319010q8Bv/+GFW5uW3O3jq4u/2hTy0ZKlZyGnkn
5q3JiXLCJQ5BdzAWgMaAr/dOAXLlcg2NtZFRzRtl5wRDwbb8niMG14P8imTMxGpV
2zgH7x6Sd80jNIfZmPgqhQMqmpw2snzIuOat87yvN21+2Xg+eYXV+GuQ19azLD9e
Xc2g88P3CWf8rtYmxEMC+QvLBnaS6YXz/T0pG6pz9W8dg/LwUW0GOwF7IQ9hXIW7
ERls5kNbxJ1qAn2dKz8kmyj6O4ep5zMGzrWrBaFfR1tetewiHRf/uuisyRgLrqHX
HIkRVYqDXv3yiYBG4oCp128KG5Ph2FUyusPHwLaoPeBOWYU3NieGDZx5SIxm/jsB
ATUp0+hPRfEoktTUSW1HtubMqLA39N1AKXOPhT6GDAg4Ibo3cJKCnS5+WpeT93YG
5r+5kGvqTV7xvD8iqggKOv9/X2aaU2cZIFD/OAb8th9nZZGqW9VsZT4ow70DcVsZ
t7ANZ9NodPyvsWKKVThKRQSYezQxPQ/vvNfE4stGaOemLQGC38L2DLheWKUF02jv
6j7l7Akm+WyN9Y/h8Bb7Z+R/w5y9fvBdcQScPrE93R37dj5woinKTtqPnfY+s0kd
CIEn/NJxjymsvpKDLUhjYSLgXUMDSLw75ze2WXz38pxChcG+xj7EdbJyMDPf/0M2
3LVL2eTfUkuQnNpeF5GXzhcr5aPFKxJTVpukWPevBQN6xKAiT0uKfZhZvLkpHQvq
abBNTZiJ1QBeLcZN9fXniKZXH+C7j0TJNvRccufrfKUcFyRnqa9hzNo2pvqnXuc7
bhhKuW5Rsif6aRfaDrc5tbbs3Txlu3NCTRrUFkaPGhYqXxuk1mCUK7xLrap+su01
ziI//lH4j+LpprpQEMy9MRUE5Wm/O5zVwyJFcq5BjHv08KGdPMOL+jgO6qJqLg1d
63CnKdsiwPyG94wHnZVLv9f9I++nywoCEnzBcsFNKB1RvPl2n2i994kIsreMmPpx
R3dUXANfngDBgGpeJ3Nk9rG6Oq+iDR+jzxkwiruyms1dtd4IhWMlCdshnePSKaVO
jwQfYjJ7q66ISdm5M90Tf6T3cya68IiDzQCERDjT6JV2SgmxS2AS58tGzRvqohAw
6ZpUTVFmJHZN/c7vSGRFY6myROmvjabK6X8rcob6YFu3We6p0g9Pce3l5bxQ88Km
dClWh6nnA5QJZxCVgiarIMXBwd94CIFSPn3oS6rHM8ig6Hkcg7rny+8GaAUhPFEr
2BxYmP/HWTaywf3uhqTzO1/wdKRfZ0Y8PleBNncClCcawVCWnfYkOu6thdVatjlY
WvZy2hoZb1Xgxle3wT9E3Xz1ENsiqtVEiGfuatdM27jqAGfIkaRZMogVZYHj4dah
/zfcQYFgWS5DAfVb+zqqaLQHyhoYi9ycb4fBgmI6BrGzqm8mPA5RBHJbI01mLVJ+
Ioin/vuSLwnZCXnon8bP5qdBtD1uAQfIZBnPxNtg6ks9s6oJwMOwOlEaEqlRCiS9
rQ+a2kMGmAdWN5ex54ItsjXRoxhuqpBaCOoIpdvikI8BJ2l3G0xSfFj+kHDcUw1N
fHYV1aWd+a8szrTijb3CHdIUGYJaUmHyvczFUAwkUue0yKB1KSroFtQaKUXhOz+3
E+W4zpxyDNQgPM9uiASMOsYxaG3i7w7zgYkYTM/sIwlJAn8sOwPAKaQrrqAWwENb
GdX7aPJOCe7XDqLeEOodbbxUO7b1cS3Sm3VC1yK2QLsMUyO3KukQfU2OSXRJMt8e
1O0i/3wDaAAliHd13U3Ho75EnVBm9LvzoFy5v/r53klm4TKxCeJF5XRGqywgYoMb
WQSPfKfKNNpUTq4NBRkwYqvdUZPc1idvzn5WWcJTtOuV4ruXB+eGZoejS92896aU
zCSl4kBOd410TnulMiReVndw1HlNteZVAREJ0JTYHn741Lxb7/Ini10i8xbxt3SV
yDZkhVCwH36wBvTkvaIUacwVBJ1y7EQrLfZRdkoEdX0IYC13RDpRaona0Ijq0wrX
dsHgqa7LraO1zbh3LG3Hpx298Yp5R9VyVUeQvgMTRU91iitmRlf9SNraAzIEQIyB
je+FrQYHeDRFgUvI4NQSRZUVeNzyZwSyItEnAuR2S6Yl/hURmAef3F1m0kN4aows
vxE85bJt5tnct0iv+vOIcXMBDgSRcOqk1A+mXjADcDZM+Jt9hmV81jjko0g+hzqV
8smAC/6rifBARTsruzgI0rWaJ2Exk8ddo7/utbY+KaQ8OsGRKJcDXRKtyjx5clQD
gJetvkrT8kXWBBBpkyGMVozmgDa3txbpjoGaSiMgu+8cQxw+hxIXDPyO1OWG/7Ly
w+zr4uZcp1uCyaN8UPXZg5OvfbMDjGKC/0N6LBMAth5KhsTZ48V6MeGbodHT/f7I
NQlD4hzndQfWSXmBlAxRw4JskFJT87iMBSYyN8m2PHp2YwlH9/rv2UO21Uaos+f2
XLBpapfCY9lmKjxRw8h5vss6m+sCQDBbahM6vmw+B8h+XdIDkwVkANJOti7uZIQc
CYw0k4K4tXUhl7iqOaWTE81pQIEMCmCIu7BSckQ4gv4koZn+dQv/leFQFMZY5GBc
rUbeUm+xjE1ZzUiivqfeNSENTTprPM3L9+19xd64hC6BnZd9PebcBLOKg6wokWJF
19ji1oG78QN9Wwn8GISkRCZDs7qJXe37C2jvG5A4WKNpIPcTvuXoXs2IffUY5GH9
e91Pz1WJVB6nTPdO6LBITO3uRAPRX80xsNu6OUl9klgvLnFErvFkJV8raOYdRsCL
7OQz21hcMcr0axtZWJxLwwfOUJVAz1XwYQt6AD1ZTFrXP8LwVFG800ODB0tSMM1+
FQ+G/ERpp3CC6UMgF9Gg+hU0HmyhKfX4lCg3aUu95QJ8rufrmUGYdsgWmHUgMwtn
dUjqpZ/SW7fAI0Sq+4iQMjv/jVOZtrWTRCppfR+gcBi166vW9/WWkhYEJewHQkWT
xvqocs1zjm2wQD1RPdTGIBfAk6RiW+s79W0Ux+UHu5Lr6dpinMQQuGGnwanuzjL8
JvCAk2NdYRQjvmZ7qgVuXsQDE9KnRu66kUbagIdJKJzCZ19tUnj7HQlbDGb9aI8z
fD0eCVThPSlM/fziUNNvGS480cqpS5NsGs65gwjDFE4jjhj0i1P5K/FoHHWIMIj9
oCOG4CxSYNUL1Gm01AlfsaQf7Kvc25z4SmKl1yBnE50eld4aGdb4cvAtHBw1fPx8
Nzp54ST0O+uCdUimhZ+YszCuibao/ZiEKCsofelasK6kBYUAfU83czamGPm98ocm
VtAtP1Nx3t6NuNGi/3vNDQqeu4QyTBL3VuId76GcEKxoszAf5WE4WQrNFMC7xg/6
GXC2BR5bMhCj8xQ6EXdrAmbmaZ+FLkIGo0+SPs0zyxVL9po+APZlTfY5LS7F+eJP
pIpFjRtKzqPRGi09w5rJ4AfmvwrPcNVqAfU8+xvxosVImNnw9K5R4Jgm1FFIfjLk
gImG8M2NRtnH5TUQKtEzS3RKVDwP+9szL4bQKgCZtBiEeW6pwjJLT6g4oae6fniT
m6CS26GiS99AXQMhCYEIHDudRgsJ+qAIkvjTGgJW1K/FiUPBZGcgDiKTEA8xGICv
Par8uuSbbZfpO/i0EdqRRLh0qHFFnb8a62m3QnL0WU4NogToN619HLtU25iNjZiJ
L4AO1yCZ+FoCY8Z9rxdy9GUA83VBx+KhUIi0Xl8iIHlDYhGss8aO994Tppp92s01
M4Lhzkqy6BAJGGygp/HAA4kOremwDRawFDaWgngcEg4ZGohy4Hlym/qBUvJjPs3W
6rod+5l/7uMauw95hsdcIrcBA8UgFgOQZjhT1dr7gzB0bi1/scXBKvDauM3bT4CI
ZPsmFeriOZx2kSv6eSFSlgFQB68Qldz4xFGRm3bQg9tj3voprcmHnGLalU0emVvw
/WSSgDPPMWXlom7/smAyhuLQko4eUbZHBz8uXE067pHNjCl3Q+YIAFvh68QPRlmx
FNuQbkn8rbLPsNuW0AkcI6JswPVRI0TNjSBQK18YMVXH2g8jT6lHd5+7y7lZqzu5
oiDEFqZJ+Jik/6SZSSwgj1CPCnnlvVPO8oZoNYLxAXvS95Zro0URwW9lukQOqcBW
s3jTTjyHeSzazwP8Sq9aNomZiIVupQLQJD9yFwZKyzs9xPhG+kHKl7D1qtoYTTrG
NAYrczZHEvvmcIF1rXcKicbL15qWCO+X2+FBBELgAAfCRvhr3GH5mZiWvOXq1wln
MPg8rfO3xMMErMZOzY8uh7dUsEMa0e8tFIp569WamIXaPJgVXVeAxyshHOQqQi/v
SY/hEpbYWqF+Oo5U6XgalUzCnKDLhMnO8uMSl8UMzRnHt9pe4FWjtgs7VcAjGr1M
KHBZc5h/In2r6kFsSNK5tbWbklqGh2h5CjAKkRl5h6ixonLvDncH7k4PrmxEPokZ
YQrn+M7ugt9buEMe9oFrdhAUjOFd4XmxtM8ShdspQPevwRCht9cokfho8YMZ/Bpj
Hem0Rllyt45mS4+gpTShZpBDUGKNQpemDcdfTG9+OCXtiboPyYdIPcCJ6AvZrM3V
+xjhPdf6zqIiPqI6jWi4MSg6lj5GflgN0bRYJqIx/SvD5Evu+V4eC4MVkRzbD7/1
QuY30LfEGUxea4g0C82vKnANOyTnprAnKHeJejNf0IoYWsN3yKyoX1V8WsYF00nq
FlKdI2ulZ/wTY5vOmxMR1fnfATuylw9M/ryubZRoZKWge2a7Nub6kNc998lcO5j2
FEYhRravTA1kGi1shk1H+HMxdno0vn5tuLbBh6ODWArGqTCXZRTZ+HOtCZflMbcL
dtSmDi5iyrDf/qTCFNKytqBVGJ1LwLy3NurM+dU5xSnFx6LPFiihPveFr7LEzhvp
oiDiuuPELjP0xfOCRO+jSaoz/lycKldZ9UWUIQc9ejxtN1JeT7VOYWuHwUDSe8SQ
+xI9hH5Jc/OCCl9y5p9FPzM/TZP7ThPNJMjMVDAmk1uiUlsc2sbcRJTrpoxysz5q
eqI+gb+5e27xA0voBERdU5DXtcmlwdQ17q9c8ZTJQLp7K3x8rrrvtjkloe80sidq
C3mw/MgmF1uNtAOefll2yedAl2iQuNJN6MGxsAx91WtrBTTClALcBKihDaXOuVsF
sy/VnP9/4ZnhW/Ee7BgKjNJGjhsGnjtM2/urSNuXP1EEZhzm+laP/Ae7pebBEQdG
eb/mEVKdIRWZ7RNF5MadsE5FJ5657Jn1lqBVqn/ejrhy5H3j/1mqTWGlotTCWRds
3gK/G0dmdFhlpdFaaxvI5Qf+oyTifteCpG80oLywo9ZXY1D0IhlmsIHCy4oj1pJy
AnpXG7J5mf+vI6bRsOr8da8BhxZeLNc/3xiL9IIGhvMM3U8276Yrc19tawp1j4ov
pi/cHbSduJ42GVJk9tjbJk1dK14LIYyh0O09nJqas+JukpwhAK9ieevNxd6sOqDb
YdD8B9p/5ZyCGUStzEMUY7kkmrwiN/lp7bcMhhMstQ4vBEcR8lLkwY7jTyrWt0Ay
bYaCsTceBBMbg5PRxoGlG29ZsdSKLxTIumo5eR7qT7M4TTkr4b126WgVaq5OKI7e
iCB2iH0k77uLDZYA+MUL6o6/y93ssQocMjICLnKHVSk5jcr5QmC4bWB1gKsRmyiM
8WE9/54WzfDXWQwMYAvF9TVbcjb0CgsIeuQXAoCwHVCospEfasbp19RtQ17s/3Vy
o3/9xcpdzRY/8F5m9vym9QzbBsgSVuN/fu/PEh5pX9gv2nPK2Q/76De/pnjveUrQ
jacT2J0we5Rdm0mhVkLDqoqdeoCEjtiUTVnq/4tZ3hafpJc16/ttUXZU5uw2FM7Q
JLEst4D0HNRvkFD0ESsPPx3ymA1f2v9WDjlHyf8wOCA/YoxD2XXse7E1KZj0/Qyz
CNnt39D340mIj8am6rHVBeoH+ou32lmiWV2uAAjzTBiLELwukJDPkahAUnl8tq0j
w09nI9N1JEhCSI18wq51Uox3Jz76UVz4OS5qClGMVIxiiWZFOujdX0gsBLWo0xe4
rF4QgLiD2ytu4oLZOxsfs61PlrwkWAXxy5GPza42xDv5LSYJZC/cqBA3AKL4yhRN
y+On6ZnCGvFqLumxKi1IRIVfeyzzsxInk5BRcoTHTnbqCSLnrpd7Ga5Osuc7KSZL
CR7HzO7YRvmN0QyfzyjJSl3zUan3Qse4QGzs9sSb+pnlflZkhMpAFL6gAPJrhM5P
CoxFQyNE3N0apFhJe40MPxSlb+Lp42MAi2iUUHc2R7vGowqnn1hK43kka5JYK5Yk
rBDqNi1MZ5JOVeW1RsmeMbkNQLAc1yBKONcBa4YVGJ/A2HQfp4QgW6lYJpbx+5W7
3tMg3j+D7sDMtWpiKuLSwL0rBMKnnJKXOZSjtrq/xdv+6AfUJFfHnpx9pNuo/0qO
AZoYRIqgD3FJ4xMoI72MW3eI/uLrGzc1B/q4DJ5/to7WbjTla+m2JGzi+S7ud9PA
1SwWzLi6DY8HWqZ7OTVxU4wz31vn9mbEcLISCaLaICef1+NhfEnM0V6KtNa0LVd2
ifY5jKvykaT0Diq8u7rKBI4O6dymM2gfVjkiwt6BBlQtbzuXrt5LTLP6H388d/xY
eHxA3FOabj8OG19Dy0ZK1oqEZZ65+HXujTQYOUdBwEYaRwRXHHnJjg+a8VSznIdo
Nx9ikSkshFHkL9PFYqydjbJr7dPLIf12H6plkCZjMEibKmuyO6hNE5Hx0ef1oVdT
M+b5+H8K/y43JfMfTGoOME2KMupl81QA7eo8r3Twke9L4I6kyHWTuS1Lcgl+21sd
4nCiekmCzkJFvy3HRZGu8vKYvZ3UKepuvQfOfLOVcmR3HehA6aS36dyzdqMhnU3p
UzEeuufcYcIa8a6hGYrfb+xL/NlZb4v6s1zZFmurbSAWZB8jKtET/+xFmVozc5ir
Cl2bd063Tu5qLQZxT+PD49U7XdIauxRGaunMptf5LpLNrunu/m7pmzIKcZNA0RLz
LDPB9bYfjrlPNOn6YewjBeaGXxpX04FVvi2DK4uBO3yWoOh0HAyxILxO6uWsX3bF
EiVcUPzYmUf3BkKuLfD9FzRKP5BiXWzt/Xu+WeTiC4eFI0n3qgjDdCZdQpyMB5AT
zSheCW0kBSFOi9X8W11nnjz6a7R5E0EoFfnI3AplCRV5e5dZFnqsSGQ/phjBG1ai
fJMUeVNAYtLVpfuuD1SjVb/N/c2FQFHNl2YpvIxTAQsh1uomp1vHl2f6BhlhmKZX
iXvkWlgl9F1tRx9IL25RTRinKENfuK+sjncRclfXWcAX2Duwo913RxDKd5eQDhsE
PqZIfU3xXlaDjtdATwQVwdA6c+3oi33/JYNhfom1JhGijFsrY9HPkYy50EFWb1VY
h1D0CdiWREcqZXZvvpyVmXRaYr019LTZ3AgGgremumaBj9DAyJMD1brDFXy0Kgkv
AYhkuMReWkDWFQITxjf63r6WGwk13TSgWcL3Y9LNMAO4sGd6ne3T7TRkr0elNN8Z
+HnWYLOu/tkijxe7eHJEdnymCXkH7v+CzUk/cj2JvYCmodPYlHCdxK5zuXibPxO9
/iiwfu47tkI1f1BD4xIoDZhHL2vH1CZZcPcriIy/QYpr+v/lR2BjOLv95fZb8KNa
75J/LuB+Y49EGzmKy96m27dj7i/1dJ5YVb82PlCi6ean2L8KEVtkHkiVbwyyRBe5
YUWvHxNBysWE2OJl13FQzHpez3F+DW6vrdFP53CSH/A6mq9KBsWyT1Th0uQbe7O4
ojFYQVHkAvju0bbXPGRn3DayDmQuU1+j5XgpFuFPK1xKtP8mzFw9zUeJgKZsuZk7
fEQcWGV66gsk2+0SvazW8SDnRNmsNYpLOMORWxWPUh/JWA8P+/6wBKHNpnQSx/c4
Fz4Uhs59jOAt+y8c2tOJHygQNIGt6GYGqasX0qZPSjkmZdpalW+R8vNrus58EBlV
o4qYNXZDn0aiLGq0XhrmzsjYpWdsQHJ0gI+IeZqsEsGzPGQXj7U0lZpuqai4FgsO
r0GBJRBimdr7n86ykYAjQF7FLlZU+qDAPJ+oNSGFqLIhArYiAwmXKwkM5IviNCnn
jZ/ixmapY8XUHtIDWs/Z0Cp78/rLX8QnoH9N6pm4oTOJezhwrWLw1s+HDNyM9Vt3
62fZy8aKSonqbaKg+31Jo6amZYsAv7um5hy16COL/3AQKvARY2bVrCk9SNymp10u
6LCB25CPYazyl5tcApD0zQiM5bBGtIyb/bkEPlZJEidO3CaPTHNoNpFbzQQ4Rr93
APt28/cmjzvUkyvqDoTKygRX5dFNphYF3lZCM8qt3hBjqcrb0yiH1w3O5FdhLurU
kEIGMpifxSaL0zuBO/73qMEwpM4PRJTL+eILPoTmUOEZ3Pkz2nC50Tl45Cm/f0eP
D5xEOJoRmFAdpO/dBeC+B6QbFQJJlOsNdGDbooOZFoy9hMi9pnAfhfW2kHtk5uIG
8yYrIUjb7FCAwEmS270uPt82x3LyqN+jDhTVlVENv0lKj0wQdP1Q1t+zU89aZbur
dwkv3DzOyoB1rWVp4KbEojkrugNsd2v++M5Jgd1ph7YkMGHigrJ5s9WjmvA60kSS
Ui7QAAMgbiL3Y5xwr6ybCi+qfA+I+hlQsQ/FgKCT7sAOv8+OXzB10KfO3gxbgNVz
hbKYtF/64/KsePSVE5oXEPBnw+Os4RMBxgXEFuxN3d92WSCGOIdA0v6Gybw26PAR
4DY06c4G1huqTVlqpFpH00LQ9mG4klUOL/bSKPR1HWKkbCEjw2nNIZERO9vjaTTH
Li+ePwfFHmnWivpoTBjGhv7ylEA6rxP9BvDDncfqEKEVWiCxrBJKd9cgxl/nDQux
N9741X1k68X5jUEKBrHxMJ4CE2QuQjSD/eIxxcA6YrGfLqiit1dkgZM25bcdBZHW
jiuxhOxNTJtIF5xTIDdlD388Q0CvaHXoQCqfLJk2yqWC4iaXxHw47tMBJzeEuVYa
qf8EmSRFLbI5H+YYGjJT7Kb9n9wGY0/p3zvWgfcXcLfTYiLzJPLtJevHpsWlsRn1
I4uDj5qli8M2Gj07ZXsV1Ly9Nbd3MybDMVbUivJu2GLp6iJ5J2j8t+s9YUjb6Ubs
nTIXQ4+2RWQAE1BMG73/sVVq7RRm/KBfDmTFzYMsMkAQMIzbRc1yQ6aqZCQR7XdV
pC2Ix4PM43fqE/IkiVaniwlynx9w6KmdJuCVnfGNNaXj5Yqzt+4BJQ+baa0D1X3w
Tj+5r3VbAzxl0quqdywfjc9zXMuZUVjmWDqM307MbfV+GdMlu/Opa9btLt/UbWqy
s16qatRDLW5nlzUgTZhC0wp+r0Wt1Pxvxrxro6qnmUkEgM+EGHTOLR84Pabf0hB8
h7UekTxdCSpJp95cw7JGepgXbRp5fFu3rpo9/MFVNE6IaGe2wF09u9zaBd47S2Qv
oCLPGlMw51Lz/SRHKqwaBX/qk7fCowYj5tkArqAFEZ2iZkVKboQ1sqCkNq5AVeam
82JyHWvNKsFR5+3mB/a/aoaqLw0dJr+7RqSkVCCJT+kBhV+irbZdMOO0dNgnjUFa
qXJO4wIGvFuOkNvjmSCXNauBvMF7q/LY9lYqVAuw+my+1kufO2+mGG8p2JGRMYoC
5cuyTGutqp5em1tlKPfLPvUFWiTIkk9B7NuvlPCmDiXiQ8hXbTM3DPLQR0VCoJIz
rnG8lNsSAdgF9tqQXzmcytLQaHcFAmBgnMKF0mdEYyLh2N+zfln0kmFOnxSAjKz/
TgeOkWxa7D+ji10EcgP/e83zvpQl8AiJD7vbuJt7JCwWxjKrRbqSDWMjqWU99pWN
4A5VRdcHygczEvkIBdP8hzVxLWKejzJ4Db5FuxYYBJFGwfEP1ldKlrS6ZuBoUZcM
aeGa223Iz54C2cWdQNgW0kCY1VlcPwa6zcNxZPU5u/s9C9n74ZL2ROT/hh7ZWM5i
3nhyKG8LOwWSREqrtfIIIF22+h6OWlrxELQkfpX7dqwqWBPUoNk7isoC3WAEc8hk
Xpwxr5ZUlmYAvF/HmiKyAEJPwAJCxftAeblS2zOf3Yzzni0PMMWEAS4F1Js/Zi5k
UYKtklbtezm45E4FEdtxBbatd4bVUNqKrX7oOUeWsogbWCvG/22WOgeOqFFGvSia
MwtcVqdKkNQdJ2w3Zz81EP0LXDAVcHVRees0NjXmbnkfAxzU90WLwmR+LGK05g1P
mUjrBCyNMzpCckomsrNX7rdZjkhEBMbIYFl48KH7tBqKFuohbsMBT9YuWVxgJtE4
efWiiiMR5TPHjw4jgBREvtb8PRJqf3ourZGL0tkFRQzKjepG4ZP813z71+OfSqDk
cbp0uFJhtSpGkSKVAxCC8XtOcBCdt0E+QEK/fQS4SX4fO16YXyl1jAso+PLcgeO8
b0xZeWzBsGqNeWNdVepmC8mMUzzhzgFIkccYFk7T8cdivrBatsTVPG5Lc+5Th/tw
9g+StCRxlg7m7ULlPxuRdvFU+l9FFh39myOJR3WA8d9wMA6pa6X5xrtfkdyag4/i
gjWab5iFL9GjfbaryXSWNX9968LPEf0CLVVPr5QmB+Myf2bP204yPwwrQGNkw5pL
kv98YEe5Rg1184HOoCRpCxYB0f8srZBYJccHHLCcb7Uv/EMDlFZzTqLpqU9vFWmp
zd4V3mbVUUaaJvOrQk+ckea9h8itbUmiAQRwwvzw9UPkNxsiA/vTkLVHQFzV0sZA
nzBT4egSot2ZpZdB+ZmMbjz61eXDOoFw2st1b9Mniw0myPeSpuAQV6QKuUb+trtV
ko9ZJ5B2kPdYb2hRSafRyMBW48ALiIUiUolMIa/yOu0rOCmfs6cWjx/kVWKNpi3t
Nhb3QgursaFwnq4WViTyjepzxyGGjk+NqcWb1qFKAAjsULC8AYhxYSEj4SLtkh/Z
vsR17TVACrB+AveZfJpOZou2X7msQvDITVgKAA04Vp/68r+z2L3xqkkxBAYV/nz0
NbzjDY2yRm0CA+4HIT5RL3yzbrk9lgVDrI9TrXyTjmxGxG4SL9EY9xRF3qii9hCa
+BmmB3rI4loVseB6nAVNwzzKKB5pXgJt0hXlOGz3z6YnfJMVtS4am7upl/52C+rD
babXL0SFLnWpJ5ojukAJbrv26MSPNLjNjDVac5vzXZUFBWfJfMIFkWM8S1UsVr+X
cUDCCaC/L7dzqA86Nh2Ow/LZEaHGRzwhCShE7GbOB9AeyNoFrRp5jZz29PlgqOl0
Vr/hvgE8cOOZP+xJZyNJkhCuprnAl4Qy9DBSIALsCuchD3FZVkYuQgIve3EVxOvb
yYXPerbLZWKUwS6ILqqSXzycWzG0AUudIWd3NdraFQlmONQqQugychjfOldq3YAf
QwYLTeCI63ghzG1bN3vfzqEstrRo9kjyFsGRGofdtL5RSwDoIFCl/M73i4CKCoUK
Zuc7hSkIFRj7LyH3eh0XgWopoI7a86Evn6L3J937eLKXAV1Sic5IwpCGpikR/vAz
tcWHTyQOzO2+LrdgeXwOpCiW5amIk9X76dJIWHXXeWNm9EIwdlJQIYsiOumeL0cJ
EIR7Mrrbk9rtlz5V+l/7RT507VowsB6HleNj3BD8tNG+aASJBV1tw++aVuaMpmW5
ukc0uR5kU7DFYACnkc9EH1GvvVx46mS9c00Z5F+nV6PI+yVtM13upVTyIONB/DTO
jOOpQ/jqJaKdLg/SvhtZX5y+m/ExJZSJGvf6Q7sQcMMe8YBk3EK60a0wXVtPEbAr
zuaaWvkZUS8hYhIYjCI8NrOSK8BuqVQujEHOKx9NaxB3RHpfr2i2BDTTUR6TGEGT
4qyS5JmUo/Wlo1gxfsyUILevPwcd52QaBRy93XhUTV9+KZzVarUDU34P13b7gmRA
fJBtEeVJ5QUaXQBPC5N+kgSTEkvS3u7lfXusWw/jcBLw3V7i9PPD5FXcNHhc0UoA
hwG5j2VdK3hOO/5LAda+2uQynG3gE7rHOER+lufIND519R+/kS/iUHfCsXPMgtqY
8VzthA3E7UcU7LgmGREsEAAHT9mX924GH7t/R+cqNFec3064IMBli4l2WEp2xSnn
nGaxmhsAfhAPXI7edQeI5ld2d8Sik8fPEMKC/Z7u/x2LO6b5S07Q5UOr4UVihL0f
EysAiDtlEfVcP29I1bQI5UG27quF4fchGYTcRgiFS0o8w4uXZTDleLIGr8NN/XF3
WqT5B+lY/5I16suc4rO/NuFWHiZz1/ouyYyjHW1/HQnqvcfz7GTgEnr7GmX5CnxS
sLALOK6NBWxzYg7A0IfRKJZHFVWJP7deX31U3PFwGMCYQL5lZ50JRHfDRKwt9dAX
C5KYs1Qm/Y3jr23Si8jDVYK73kUUpsxa9oT/Owm78jsFWfEMbVeDFFC3UCKiKN/l
NeTg/gIPZgxP7MH2ifAhlzfD9DiMLzEDcHdC4yjNDyRuJi7ELbX8Pnn7y3MEdf/y
5kQCyqJoQTkuNi/LEbMWScWWu1MyLor+WyLdP3ca22zI5ZGVTT+uWuT9CXFm4frJ
8djlNQws2V/f7Tl32FfzRmtA83NsJC30GWXANES8E7KrbDI5DxMLod1tEwR2vJ97
nkZ0g/YvoQQSk3waAWvCT216926Q2hhGfjLFs0+3SUpAx1IR15RMxa1SrRcphOaH
HsACqJqUl7rlqIbdfHfi/HuOx4v42zBApJXmBc4Pu99blrMld1Sb1onp0g4AvKlg
l10mkEnBTjx8htKB70VYReAjqDzpJogrzA5qLQnPaoE7dpfQl3yH4RtW7mjtjrjB
JoCuh1LrVqQPEoEojgTfob/MULNyA05z9cp9/07YPWQXHEhAvNSCrw6bEgcWv10F
hAZitqcBh9FgMMP69uMay+jTot5U4XT4HGCKztr72lWLuGQSCq8dIoMrrvceuO8D
lDmDEc//47W8VAhHRa33DBWKu8vhi/zC2bWBKhBzfHhgnLCQSyQokMXwYHL3kVNO
AfbNtcTdlhgWwVShJzbWqxLmAnYzxzMFxeo7xXkjNmu23q3FUlS1pF7tVSsIRBDH
DFyaPG3sgaCaMM/17PcSYhbr42jYNcHnquvteYa6IKy3sGcgo0ktpYNszfVm+hle
57Ju5KXW2qeBG2l+X2H8ElUXRcEFKtqpXO96fxtb5Jk/yB2l/KJU76wLexyAPgCT
me91IPgnBG15s+r3xaepZgBtTOV83i+u8tS9LhB/lW7rXgcv2so3KsyfnW8eX1WV
Mxmv5icLHsJwctGLF2FnrQEFtjgLyZe0hVUwCr7xTo+sqNxee/RuSE0nR/lepioC
rXDoY7Ok0K6A2PEg7svZUFk8hvpJq7tLIZ1JuFoZqGjjoIVr46ihfXNYHU96aXNb
Wb5UoucdTWvrYVELgPUPnqp5kzI+m76z/mrbADS9PzpSQSNBSg9JvAomV0SxvvhL
7eFpJXVIzHFZiaaDzpDmNXHBsXd0cewYRSU9ubnv/UIb5q1h56iKxvVbflw+X2fS
pbMaBxNeygA18XUYmJYmdkcpa7NYqUQYR1Dz1F+UTkazMXScOyxx/UaxQ5BUQ1t1
+3dyxw7rXL2OIG8z9kCbg/1HlQgtXGvyf7VtHJlKgSWgxIMwzyQbW7jL6RlxuqH1
wSyco5eXGVFVY6VpMlJKxAmN2wWl/47hTMggayB+OxGpyB73/dzYQYoLavJj95Gw
GhuilnuwWqtwygCPCSsf3EaWHSu/c+8/JUukAybJ4u77c1kveh6FDrYyaAljARhx
FGkwbRiHhOnNuFKDQ8EOorDTSC11JY5tNIKbSnBvU+dP6B/E/ba9GVuEvz7KqFmr
tiFc3nRg54W84f/ZmvnDEf4XkCDbpHmgbrKr3c+58lM9UjdmbKbOa3HW25+nUwFA
GIkP8uiMOj04pBAsPQ4m2rEGx5S2r53DWqdA47DBWeHUFKtsBq6BV9+S2GVwjktF
lZCCw2nB3V5mHhF89UtBTptJ7zo4WoPbl5jTOh0I+5yb48mJTn9ZLS6VnWdLmwO1
42oxAtoLnD9BsR5ORGgOrs1u6iaHM342x283cf1z/+XjRJQyLd8Djkp0gfRHskcz
qRrWeyq34UfGG3AmpiofiRxg099CXYoPxEz2ab95UfXfcgJ4oe0LGT3/ViXS3kOf
1J20QxkAOOWMp2Vg+tsB0Tq+vjCZhME7huG0rA8P8kttV2kwcUfYinJZr9LYmLqX
NrPmshAnaA+xNLkTMeHbvAryTI2lkZRWKHlNlPFRHpyjOSKx1k7dr/d7+YUhpNfi
QFC9YD8GGcwJ1nl6Z79Lr3uJMkVEnsYEI8MhaLeKOB3wWsiVRQ/JW3McXrxKcuVN
Sg+tlLuDt+Kxwf54QggtoTzvadpj7fDY7pjIBnFEl5Fwth5qhxtzeEHacbFtpNBo
OMPJKRKOt+9GYLxRaLw0lfPzmxtbSeyTIvEVP5LQKkkei6A+DzghPoFKF7mVX6yr
mIVWOXN8ycOQ4EI0O8506i1eJE+hBlxqC9ZcgZ9j0Th9a9J253gUDF2YpFb1HT8o
38lsuvHsyAqvDgcX0ZJM7oZQfL6JM2CstFsv6NPMWwulpUsrVGLIeKvsIiZYMsfP
0w6ah2sfkP6P0E2ziVuuXLWOIQvXmTwiHxJitV943DkLPDih88haCbIie/3zBXVZ
GVxiVG/9K1ZouYhmcgC9ZctLnHwRXJQ1/Z1UJuxVY+VM2usbRVXZp1GrMRWfz1HO
QsEnWKD+hPHy7WitU9hs+AYFj2twftxPIa7vaX3YLzyWjMyOhj+vh70vLoMJ624q
w44BS+7MVsPpq618TpzQNAGUBW0+a3tvBZFXWU/kKO/1ZNRm4r8FexRXh2YUYan8
Xp9Qk6JDDl/wrpQylzHwDb/7e4+qCkf1F0q8XCXN+KTa+VYBWz6FvnNRPMOm06Hm
rzus367Z/bTEmCloOG89y2iCtPgoWJlS+xWLfYvg6FlhKX34iJwV2V0yqa+Q81Nb
+1oNrtFavmi6DBYy6IpUrR7ut/vbcoHjHx5zI8kJyWClPCoP7tTmrqERbShXZUHS
JZLxf0NXR4DOnmuXoMb9I0qidHZxbHWTtVzbb4HzEc0jzbR2wHoZVbKaQwdN2hEI
CgDYLWAkpDq1fI399iDg+FuR6or4pPfxBfKAQPAokMcP7njLIQ0VMTvZlYrYSRyg
lfclW3bLkiwhzqfKt669StpSt5xy34HSDanOs3gCGwf6gngRJgMtfEH6iVatGCQ5
AfSv73Rv2ujKF+mGshyT7CPUoDTKwwlH+OnGCSSDYhYURFojDvIWvO2ImxiqBBU2
atSYtG9tapxJosSxvrmgYJ/4bZrVxI2rceQhB+H6eYiBtWlToMIDO6qedjQEz7TR
iHj7P/CLVDXBfKVmp3Zh02BRHekKmQJ9RnSy54TJ9YCD4FBedzgKYkT1LCW37K36
huUdx9vKyLf3Om92Jz2QBR5ixzF9ZMwOJrQOZojx9SoIivyFhwo1q2AUF4Hq7SIw
NvY+7WL0ltH0lhkwbwYtdQp0nsfQ5F0m6VyNe2poxnC1TeuATXMV0OvSce/Q/TG7
A128MR4JAFryQggZXtZAu0z2YsTkw22iIp7F6KoJdJManVeqMjODZs6Pn7YQHbQ3
gPm9/QmbGhnZBG63qhk/UlhWwTvJ6baOjJEfoeA9uAUCzB90p23R9fTFEb7p8GxN
hNkk5FEB0bw5MOmXNVqJRbcGAm72lKl7EsyA32h9rUStoCl9OozxHBA/g1NzNSFd
ZHuIDkp3dI0YmJjFFzEm3v1cbGaF+obcsZluAJowu1kjHh6Hm2qO8vgXAnMIGb94
03Om02pILbEqRWzEx8gnxVyBJsTR7bZG9flrbtcqqBAlW3ccqw83pwlmI5SiDFjj
IAVchtasmOGHB4U3U08z1R0BhuDKc+FF6y/qxoZBdxI4D2/n0ZZGYttQdYSwJfzt
CXp5tLd5F7Kg1exJLfBB51xrqjES1SKYUbf/UERTiNOFAdXCUQIDX6X1h9Es0yzl
GJKSCj04SbK/WUNVRE9JowHDOsJmOFPQpiNKLVIT3nFQACpc8IQKmePkHOgdTkND
2SoLGn0aOUBwVBZULM1YNAG8+G1O3dn6dx6rOSBPM3d095Dp67GZFoeV5/J5h4Fi
OJv7dEkVVQ4uQcvWOIFbDQBy5GFzEFwBLN/rbtHxzYsyfMtE//x2QakZT3T4WbqI
kKOO/WQ6aYQgNWP3CwE4cvavYBmggYJ6PC9GnCKCeTjgLwZe6uEIEm774r4qUWHE
By0HhhqKYeDzA8FwD8Dyw2uBTi/Lz+iAKDhjxER4oZvbG4BRtb8/uEkkuHtQY4+a
Hq1HJpQA8v263GYW49Gm2BUbyt6X+PYoj4KjHPibP92B9APD2OvtD+UFqar84Jdw
0TZLHXmcQThodKHiGv9hfLcMpAFslyUt/tjcIspJpEez3BJ+H+peyVYcDtbRIBXH
cD5QXXmu3byHcWBBDZdNlJI6DNrX80Xx6SaY3ShRUqkA0vKEU959iTp8996i2FgU
BxX8Q75gutQ7f8vxMpCTK/2F+zUtyWpAiRr8RAWxYf2MEUL7ZrvrfVEiJqsEg6eu
Rx1lEK27roB/pmF0fwmIHWPseL5r/4m4FBThX5KkTyTiJILslBVhPZzTQwwcd/b5
i7sVxqocF7YaGcV0dewXzssyz6NjY6eCmnPGSJLdcbb0Oc8xU7ahFn8ICLX1VNJJ
KFTnUJrorciEJTGSO4zh67D3n2Px9nEec1qiF/WD+1M8dI7APmy/CBIQNTayH97Z
YyC+Vv1HAQfH1zeez0Sk8kuU54PSMSjFa1cGHLFj0a19x+zMGwwjapcTPUe8U0Z6
rgIuaDzFfpaK7iUUfRqVUz+epy4TJItODvZVGtCcj5e5G9y1pFL99pMKy3w2Rb/5
bMunKJGkXG6RQdZWBECp5OFxADJdGkxUGKuCMh01qkhMvvf6/2whk7JmSIPGrkvJ
UeRvpplPv+LKPY96Ppwt0H3vs5CS0IzH2hxiy31l6h51bS24wl88OQuaCA/kxxFI
c4SE2MKoMXxuNKzEuCi/DhfaymM7g8xNqQeVg8J/AFTV892zpWX6ZpwwNPxw03jy
FfGcoYxawT1/XM3S+dBNDKNkKcZzGjk4ZmLq+XvUVS3Km73WTnpXwmhlWVtI7Op2
HnzWQLmYfHH+H9kIggZpIur/KhyOq/gvR/W6e+bIWGsV8wO9ikEAvZddm2K5PQwl
EQcHgJZrgrrYa1pTJGOup3n7/vAgyH4VyfrwG2rR4LqhwEHj/VTM8gQtE3FhxIEp
q9kzExShSx7YuYa9PwSvtvQSfACTLYjHot1GTVjpDM31lG3BhfbqLFVEWjjwcQYB
gIeEn2Qjbe0rMNCkJzpMmtJw7udLYD7YYyNCuOZxrO/UV4/CMt3mdOzuoiiz+fa1
q/tw4BJVecl5zjFSqQ7Sj+XXi0f0tjbB428XvuzD3MaVENhyPNpz21JBCFywDTy5
OhG9VcFvhmSdbtJgd37HCqv8urPBw2uRqXvyQl5Cr2YN0vrT+J/B3HbS0r3rX0Jj
fDfBxekdbe/yCjKsVR4KNLbhEAG8TpZCVDjg9qwyOapGwLP7VIYcnhkxIYKQmqce
XUZucLI0cZZvbRLpS77J+AUNE+DKls21bptecESX3Z4Yp/8JrMyb5h+E6ZTz/Wjv
yIzZ3Z9E95eJ/PJLTFvbQ2Zfdixpj7PbG3Z7a9shBPNoG07MeFhS943aOWoeG5dR
EM8g515EYRxc8QoZf6tOlMpDuxU58ugTrh8bOpUJLkYwG6UisTnZURTH5PQd/l3u
WUo2rADWvYy/cLxjfA0IwJC1guwm5mmue/NbnYJaM9vqpyZxVbD/iIc/Mq5683uv
qwv4Hqavbr7yfsk6VUR5a7C3oCaVbe0Y4q+Ir94aavrlKlFPvlUKiOscJgz7ANBW
+D8uMat2McHZsGSlwrUTRZd1rDOWs4CexgWLuckpBRnnNCWI1Wd28zkTRJZrXQHN
T3ce8p361bAQgzzYlZf0fkNnLnE+LtqHS3mDV8NxV9t0FnMJqm/4pjkTRFD3/2Lu
h4exJ4nJfHR5tQATgaFHGajSXFzH7DxRUDxK3FtfJUfFu8aOkTG196csgyrs19uU
U9+NPJ0EJE5sL0RYCizhbOP75PhV/tNjpjHMfRszv6sjVAiM4h+dYCSo81M6HQ+p
naQTeD9dnXLUzBxtunwkyKEQIdCYofTFBLKDimEAayETwiw90x6fupkBsQl4HwfY
lMy3B/xSBRFq7YhkQtD0ZMa0JGQAZik1Tsn63/bUfvPq9GKmJ1NmycYrJ2DCRiUU
c4v7vUbxztc7PitsO9J5sZC1YPTKfxdW+XZMQFHLbqs7FYEKj2u7aLTdxtyCBcTA
7FBjV/1InJHcr6xhENfZ1o8cyrpRqLM7yE7PfuawZGG7GaxOBau/M0iynpMNJQO1
73oHWLcUaziqZi9++Dv+lt2EpFkp3nxkAlya+mt0JC8aGSuXjY7FF+9N/ULwYmXU
ssPEuYE+3rB606mTjDvm68tAIzzRQ1zB7urm+8rmnhz2qJB/9aexV9BaNZHFHijZ
4xxtO1ks82BsKVHLOYOgM/68woEmd0P88Lb4rDXNflD2QjW9Ain4g2ICgbc5FSds
o1B4LzDsX9f0tO+GhjVjrdU1WV10o2KXp1Nm4Y9oAWSOtulmI6+cSFi0RSSNSNJ8
0T+cW6+2nfTSsr/ybueHyETPiuY87C7PFaRaO/vsv7wwywHTLqs3h95qd1itSz4D
qZhnWHZ/+8fTnPEg02rMiJOuYzo4zXVYh/fo72k66z6X7l4BbdVqvwN9LPGy7HT5
xd8f3NkvOIcUG8buBK11CgSJM3G/gFBuM7eWuHzf/TIoSNwbvxk7OIvgV23conRP
GlxJbNpZvG+lWyt1IFq4h5OKxBR0qFRuV+M7NUxDhNOqeFehTgvCzDFWfpNxZbV/
Ia5ABGJdoqHbCmJSyHQ5QyyPPYkMIV2gAcIo7DOPDBr7uku1x8eLbBv7wbgBaEN0
7kuWVp8JQH5VeoHnMZ9VXu+njvlasIgG4yb9kJBv0bNIM1R8/WDeBTWaXQUe9Mce
moTVyojqyfktTjL1howCAPE3CPR+IkfH1YiWw7xVmgE+CNWR9of4x347XNj5tgVT
PfoUfaxInGGvDAWIWvWsTBGiIW5bwEgm6Vdxejjw00DyNR/sBBk5c+xtfyE2Ba7M
LQUrbu63n1rOMshbveGZ7YlHR58C793LwZq7WRuHQrD3qPUUTbEluMV8s91rUoni
u+LFjRTcAyGfyketViMDYQwu4YLuZpTjHzR5/D+tKTU6bwhOU+kplmgXVb2zGFad
tHkrZc4oQJtCpdmvFP+jV6paTG1qSRG2UrB0hGj9aL5yx96NqBvxWbodgdL9IDIr
uNPjEg/q52CmipFrhln1fNJDnR+D4DqDVRdJV9uqXFTYqO02VSocV+2wpyYtm/Hc
lZdQn+UXRoaO0i0boPuWr4qeC6hIZECiyeJ9tBFQXp/FZKbY+B5JzHqYYDDKUFAB
swW+jI4c7VVVt3U+2hixW77T0oUQPZxcuujVpXrnYP+a3Ehe5AsZlRQmRNALB/h2
kUZITBkZhuDXgI52JgQ/7IyhHb0zwy4IVh6Llccgtao1yLBzhEmK+/PteSHHn+Cl
FWmtcWqf/doUkVqDput8ZTD3K5tDTR4rqYUqfQSR7/NjCJcpt5mo3/w0NGkk/JMk
grbQtw33lQgSjN/W+zscxTvlgbb41Lidt4cHILaGATvsw0D+9Ogfje5G6JTNzMM9
6E6Q+j3FoBswEKy3gtp0rzOKPtDpO4gk5A4fSFJ3rXx6cuq39fH5GtVg0EQoPHA8
zHTLhzfJan7ozxBjla91uxvE8F4AMyT4+oHgoj6rzImB7/Wi8r1jbLMJuz5iHGA1
nd4WDCqw/y1fdJ3fswG1MUsHLkBRv4vttBfni58bDNwIMlsa86ngdMq9Ovqm1diP
HIzmn0s6IZPEBrtl5aaInqACgKcJSBeXxXUY6Kn8cFNHqWlARmNVLdk4gS6cozAK
xz61vqkh6s0P+ZQ3O6Ry25CJAPQ00IqNWnvFkDNA0NIGwsasU7/55FmUWtpNwK5/
QtWpqHkXHn73/tfvsRI2kgGD1uXhI/mjc/6ZnnTP/KbPIIV6vsOO3J52FLujTR/x
EnzHEdVdtvV91wA+ffdw8XR1nUAss4de+rWuDky2++9gYMcLVX3RypgvKQm2jwxO
Zw5p+IQxzsQ3Zo6GuUD/Wnm9Gs3va+R+6mAskg0+SXcE/kdDfxozoKj7HKAmPCBI
JuKugVPVGoAkTqwK6NNdBwTYdMSNhDjVSIwizI6UMmCtJwvi0wU3KTqPVR4azui+
179k5mqzZmQxOMEmPQpIQZUq1QOHt30VTWeMAqOvsVwpAkATLMPdzP4rJJr9qWTA
RyX4ERSCeADOuyJ9KQsu9FWbS2WRe5225rF0aHfRDqql6lgc+rmCMIP6yjMFyePb
0fqwHF7oTyoFRhFNwZ1S/TU50mCqcUm360WCWQvaFGCyER0R5RunWnjSaTSfdKCE
qw1QW5gvZLFCC7xuEm3HzVM2DYz13H48/fsnXk4NiuJdVEWF/s/uryLSWFEM2dpr
U1bEvwoZ0fkt6XVeiDu6M8MA1kAYEDpeYnSlh3NquyA6M8TsGefwaMeTBEa8oQ/S
6hLmrk14XKqGhFRMbg3Ohm/hEbapiW1yDQXkFz56kIcj4u+lqeqhJeqj7vu/jOEU
BDN8xswfWgk9ngKQvWVB0OYeQ++b5dFsJOBSFj26MU8CTmE5i6se93JyRr3arDJX
WFzz5avjkis3gd1Yy4fDrWkFj1pSJTyh9qMw4YFoQ52nW7PPcdZgS3hBwbSUTjzy
B6hQmmQk77fcKUZqozlMjhcpmLa9u0d4rq2kOp/Dp1Sy63ShSEQMXkbUzipxveCx
mixyxBFpICKe0rL7bNahGMgpCQOIRCJ3U96ox5VAtA2Xa/7JKoJl4tcTBWN5oLhp
9mQ8rb5n3lzTZV2n3Wk+Lv7+C6VvWzEhM4VvhyWxG6vvTYQfJskoE+/FHCcdA1VH
+O+rDmxLiKvjOe7ncTWALIVkcKxtOkmJbtJlMhffmrIxjmmLE3NdTYE7R70rwB/e
8LUTXmb55X6/G8mbhBWDqpj/bw4ed0bz3HLJ4aV0PRCSZ8iWgNyNTsAmDM7Tzqkf
THrEilk2UZVu8o/EYuaw1ucPClLjjjeGf4cVnyhI6VUONYNhBTSfw4QYRafOKs/V
nxUXzkfZ58R4WjCSLO7Ha9Ur6HqxkNJ7PULZ0fAX3DcEUnFIuOh3MtUTscDP7vCT
8Y0hGJHslE+T9PafW3E69FzdvE7WoqAeDWdvjOlQD/xlj65uqbx2QKs7SGnMw0pa
pZBMUNaXuQ9m5pv4BVauHbUXDLcJhUT9KwYXms6SkkEPVKBar4oRXAOGfp/KWAJ9
feJ5QprAs9hbQVwEMxY8R+Ts+KB+iKlMYHa1QMhTGRXuaVPxJCp9buMs2fzmUVf7
VL90y9GPHiSb9vu98iA2v/q+LjLR4m5xGj5Qz+V2tbGgCaMA1NkjW9El+hI6dNWI
R7LTkgqFVWxDsbiyfaxay/vVQnt00+RXE9/5rZmEnc4ivBpCP4fx3RxopD4rDoyq
6BFrzNvBakQrfGQBLTE8V2O08rx6YJ/tgzQfyPiNxYodjGJLHwx3vqwzfoztRRfx
a1DYjEJxgnOdmfD+H1Du2528WoYFe5deklDaJr0rbRQFKguwi5Ostln0tCQ04OPL
aqaIK0dXKBRf6iE+05QONFoIibO8iaZT112SkwUPaVL01q1SKlmiMvc9Lc9tmx2n
C7q+ZmnBBUrlTY9EMqIOjMnOfyGt2dt6wOUDJdWQbB4CjqmJw4XxpZy4PHeSiGw8
XdH1QKUPg3GFIxA2i6PTVxQge3TWw6oOVm2IFX8DRoxRnOwRD442suzG/tB4hJ+U
JA7wn5PR7w1ObWpzIm0CO2PqezmCxaoSyVnbo/MeRcBMydZpromY8mz6sB/F4cet
2Kkl6RlW5v2s+l4N5ufqqIsgnBOG3tmUcWy1zG/rwW69ZQzWxMMu6mHm4YZ9Vx2l
CRguudg678XUXPBR7oZje0RzhUoMC0oe8VHBe6IiBwuNb/zD5BXhTx2cCly9VFdt
OLCF5O7oqGZ247RewbAJxyX3csdvkt3SHQK5RCG3Z089jzKodPRg0pBCYFUNd9IR
8+VPcEB0cJlqKpjSKpP19A1q3FdfLf4KVDhb2jELbvVnKw89uoPuKP4+tI7H5Y6B
xuVgXHI4lgFwOMna4JmtMc+cBSpElc3XnwVN/RqlehdUyG+WtDwGwHWtosuXHdVB
8G/opvebUBjeJ/71XCQ1yK6PtKEqdxsdExq9rp/8Bmlkp1yDpIB5y+gpKFT07s6T
ewekhXBMeYdeAfcHikaIdYbot+t/9+oK8YCqCO+wIubX/Udg21dOQoiy+3eW4zxp
srpPH+bJMIFi026yN0+ZAONauzJ6UdNRvhsKBK6AQI0eOTqSLW//qOJN3q0PONk4
t9dWxU0D/pACZQwY1r1bCcdL9FCOhIQRSz+YNw/jScAZUkMm0wKJdV1VEfNnAEMn
zd1DmdPqRoBYsr26NPbe/cXM8bCxXMb1pzu7FlPX5/FEtJcwOPoA0V803LbTOMOf
b98b/97nbX7poeoNLcb1EtKGYgecxv+//K+Mbm2pUxZ3uIvib8EXohPw3YOSROQX
77jVkiWKOvHrakZKfGz+8vfpsSjpm6iO0b9QET21lT/ls7PQyioUt0j6yhaT8MI7
eD+5Cbovkpob4cgkyDaLhy795xR3cJbpuN5p6wCwXc0zpyIVvCWA46WOlReqw+0j
66QT08cFZqom9kY3pjmynAU6fNn5Nhc2QRQaDZS6TwAvCyeCNNqx7+ICHB8+usSt
5p7r8w88VUYQb1uOpoYND8CWbOzMYT2wwCWcbRCN9xmQCvusAE1sBc/8BfNnd40F
A0w3ALoungy/gnOzMm/5dIG/sU+IjoPBGv244OPG7U0l5W4fkKFEoWaNCaUCcgXB
PR7MF7N/jUvnzwUySLOwJ/dmwlc/wdwBDuHFkBW3p/jFzAPz5XUinDg0KOqRN1Z2
jc8lqSbmDrzK7Nh1mByY+Gj1wyxU7PBP/m2nqryRYzr7JdoRl25/9Nbdb1kIZO6t
8NxF0tBC0k7QL2j0nSX1VPrKyw5N8bhRBYlEmnbg0NgDf/3MAxpVcQUhqVtAhdK/
2Z6iM09fM6AZ1+tGoZbQkUtMdmGcJCKMHbOH+GrZo5bUVj2a0Luqbi+ZkmuWF+dR
kaLHS9gfnln/GIWt5S9UD8wX/zqhw009ABsMfceiiVoN7J8ZaSn7nh7UOD/El829
MjKP0+w4T23uy2TA05j2XokxPu1LRnnAAQCvvqgHMDTNxTCQ2kjT/gFKqcDGHf6m
/gkqgd9jQF0ga3y9YR6PklSbmeP8EqAF53tZ1mlYfd0Ck/7hUAseYRvmvONOzU8x
j9PueNqeRpUhEFXzU5QBIuLm+PvjqN8ybAysqjTuuNcpwL3I0GfhfJnf1DhAC3EE
kYhtOssbHOEOCkgRQ2z6BJduo/C2XCTKlY7hZLnp7Kvgmqw9X1UX0InCUYA2zJJt
HWa10MvR2+nKiRb9I7CcokUi2SzpkZl39etwzxinr6fCqYUK0/KYUP+/hiIb5JWC
YyLwpQrFLyAKVDYdJ3sBg1lJhvW/fxlKvr/X8aRwdJ+m5Des5lQkbPomZ7kqsPxl
joUyBezi8Ff5bfCAqZ9JirDTsOqEaFyvaYzGZAC4x/iqTXsHTFZlm92zJtvpskIi
O0iWH2zjTcOn7o/+rQu9LrEgf++xNXSSwMq2TSEVKMN/nN+XeJbLnDDzwYuu+RkP
jnS4stVjRjbYZ+jSCeWfGg5U84hyR528W/lyJ0p1ntQxyuevJ1RI/e1MUBWIxE8L
wOprbjHSV8E0dzixS4luAXpBssS8EKKyDlE+zlitwK+nZuZGVgEyraeBdFmrvhbt
llGApAdC277jsyKQYr7rX8Q/eRqZu5TDp+xC8ob3iMhaSik9azFSUlxb2E5Wk1p3
az6ajWxyJCZcnhF1EhI0vfyuH9nRaADNZ7SP3NvMSi8GoJKFlFPimF/rGPrfi5Ob
gLY18Mt38jiUCzLk1cfjR5JiTJzSdeW+9dn/xWC28oxM0iruVBHmJ5f+I7zzwmgT
7hfAxuzQcY/KPtod6vwCquZ73v49zCm20yCn19QfnURm/hjfC7Pb5fT8idHRbrr7
TloMjAxY7w2vk9oBDTelRx3wAheIvHW3Ix3aW3si3pgY2rVJU6sLZf/Ol0y5reqW
MjVvk6LRclN/sod+U4ixQVI9ukjcn4S80FdxvOWN5ijYmBd528kKDOwsLZ9eLeq4
KcB5jWgX9CF1+H3yTBh885HFDqbE1YyVEktzqpwjj2jtizgsDz7lwJUbeYIB/SCl
yNeIT07EwO3nU2UuB/IDb62VXSpl5EiajoXKWkaRqu/m7MC3khRsBSX1AUCwEOKa
yE8UzwaRHavM816RCbS1hXx4K+w+bO5AMWjFfw8wFH6afL0f0zF4gToC6daz53A9
GCoGHZQn63YH2g9gHyP0eUL+a7EWiGElaEdZ1GmlVGJUNBYUEHaH88KInje92XXQ
eHp1+jUwGDSVdGd2Y1sFjfrVKDzfJ2Vdr5p3WC9CI+0sOndJn//yFnd2M7HCzfzZ
9qbfORz30+vXErTisBNUXum6EYuxsTvGD6tnyHj4gdOfL5sD5vKt3LLe2qJHxQqB
1GUPBf3ogCVU/O6h869gL812kYA9jOgqSAlsUwTd6jDUxciB+JD07Q/jOQFt9zRZ
P9JxL7LIN/xLedEB0CBDWlOchdWPDck9sXWmDW4BOJNTiF2U+prQq4kMi2r/zn4R
Oj6kfi4FRyYVvG1Vwit+2IgU/pfb5ti2zYxw20lSekWgXTgKAAe0A7pt0R9Rg6d+
5uh+CSGEi7nBqGTXrWEW2X0hBPZ1qAFAUNjbYI26ruBXZpn45nWRsF4PNuR4O5xv
NYGHGsxwvo/zf+3057FNu9V3mTyTcRRvOkARWbqSzcjkdxHHMGHMgYgywNCF7vxh
ZHM9SD/LtbYubZ/IrJXaMsNU11bPwR2L2PiExourEGtsykexGXq7ct1UOxfiANvV
ZNGyfCwqldkXOrQmGXN/HButHt5HuE+6iB/UNQ/YCwGqzlt3JjeTzFlIgOIIXsLc
reI4F7/sk+BXhF9BSNcLGuui28lfgOp/TyCGEBwWVH4UblYW2ucQ6g6g06fgLXV5
LmDaaIwBI5+9OeHUvX+/KBo65azF1KNLjIj6GvEmEjSiDElA5/l4UsyBD5IUqzYl
+ydKblZvaeAUP8hfxFy1pUafJkBGX7B7k045PjNr7c0YPP/7hVfETuAqTDwcDVl9
efmZGa5yoq5nmh5RzIQC2EYXM8cUD2eUinSV2QcNGXoNcvMDEWnm+16zI5WMF8vj
m+5OaN1Do4fhvdEZ77v0PwMgSe36Y4VaRY/xc1B4Jqwt930pbt8O8KKu7IHyu5Hn
p1PX1az+uAfwKprGHsDzClAaPVgTrQE/RU3Q7lgA82qe+P2zr+daX2pU7DathKbP
QUuy1cxJUd8zBYZHn+9yUcN7Tamymg9t0Wj+AcdPHjT+ArhpGyUEnOaDPvSVKeYy
BVauNjWuEGsHvwxA/Y6h/IknwQhf84gcHac7t6EHAiQ4knolDt+stJb0x6d3LO5w
bduUjuFwj0hMetYWn/uK5lQmPQsEaezACR5tChEtGz+yRRflbumbsVKcL6hsOcep
JTmp+Yholh+sRASAQ+xYBXsT3QEaCBAADzfUGhRSIQxHa8pzQepulFkIWUd5tfHA
Tl0V8UmxRzc9X8R7EEGUolzsyV7zZhd1mCL9A0h/RB4HKlDWsM4JQnPlrdK4u3hC
GksGWnOzWwcksdb2GSuiPOOWm0++JyrJMTyNyCgmfKSRHTm2pZYKEqgoJmNa2LC1
N4WTJY72YwiEw6iymWCySsOlMPxmnFBZr/9ljLt06qrBkJI5ON8vp84fYI6wTCsK
S803i110AU+ztGgSRlvmmvs2diBDlaU4Yy5mDZjLybMGqlkQmOjF9JVUZ9Q5RbiU
w71T3vnIZGJJQZjKUVXvctdy8d0WjjE6xyGisuBuz9qDl1/tG4W48Q0h0Lt1PVz3
WdaJMYFvSZWnWNSwRN9oGbPQz3WFvSTLq3VkoAknOLsS4nY9B1CGQb156rPDKJBY
IpMf1BIzQfVhBLrFTM2VBt5869QNX5PiD8hklTAXxQ9nmuF8bt05w4lPgCGQ0/KN
Mf9AMIcq4+M6IbYfRZ1nFM4FVsw3IEd3A6Y8oRMAdx0H6dnvd1CoxZ3B4v7ntUFr
8ikqXqcrI/XVLC6rjQqbbswjkCSpEliogXx2+v5+XqEDzMG7Axx6bl8uRaVHOx44
5WLiREv6lZHK5kl2jfLzZQTzgJYgYaihT1KoOsohpNgcG+qbd8dtG8LQvftkU5ms
lcg1DHpcP2gTZ+bmOZksffwijPuUY0FcJ8gO/0RJkAAjtn3ErejhlbFgvFHe84FZ
Y3Q3W1P9n93XFO88xiMyagH/hOFPZqwGbuyP137kclFN2R9Z+dZrRswUbiMOXE8u
TAC19JclhJsYJxGl+HRzKcdW0qdKRon4Eq2PZXFpUYEbrA+CTXROgK2cY3dbO+M6
O8ay3YeGAnQr+AaaGxtqP5AuY0Rjl69ccxCetUoL29CZIVUB1eu+1UWSjyOI4y8o
bZVX76yOUK4mhQEFHOMMFemX+EHHKH0iZeE6KwPmTmtZgfy0bTGkq4W2jYUw1pPJ
7AjAboy4WH1ffLCUb1toe2WMl22d+62vKYGTdJ1U12Y9LNPhxQcNJxLIj2Tm6BqT
Tzi4xCnWfpwkkMAgnnFexNBmTiHZohCXvRB8RX0US86P5AXb80nafmCxBsYfOC3l
Vrpt6odDK3Bx0LQGD49WmaxqKIHh/FIieaLn8WmEo/W++s3dHmG4SmO7e9yqofda
q8KTn6iJ4kR3M9pfF56Hj5Uo47kSHSmQFS62A7hkga9rUag824t8cspdQPCHOrUt
IF1rGkmQxPsBirlJT6Q2ZduCPenK4EpFa0RzNjsbm1TxA7Se1abR1LV3HXb4EltS
4NsjdZNEvybuJ6iOV7BHRA5/nDBvUgSdGtrf7/u7oiLn2rhbPmjVaG5D+rFb6R3G
nMCtoqqFpnl16iB+CSkgbl9+EtVUCzVdm0sw9eUsaqv3EJrpTev+Nm8pJRhuAHN6
N687fAg+BIm3Dihmaa6BRMmVqNRuT0WGheunTJhjj/nPayLFshTtrtyaWqjSyWLV
mS0OXQZBw73wq7t6OzhZ9ZwxzRYPHS0pDWvamLdkyrszGxG17mVofts25ZQBkjgX
FH3bKHD8tEdqG5bAkXYoabsLIVcqX6G0MofYOpZ+F/tcbtWX2BKtASJkm5bJBViY
85CVGyrwVCgz5L585XIqdOUazB4ltkKJHSmHPjLWx0nJtLRJ4JWWswV4S3kHmztz
aEtK2Z2QPYq4fZZovpDLreDmPmbVh91aC8OgTSxBhvDX0TlrMXvbRKh5C9DaeUHB
pTblBP1a11fh9e0qpY4sCKm0NEukPsfYu3BjHiyDgY995Vmzph5zxIJ828AjVWmq
yvDD0zo8asP2g5VEDq6kId3E+8cpsMJ4a0qH3s2c/A2oMXsIz5L+oHn63AYoQEHo
LLeniidpyYx7eexRbPRO+/BelyNxXWOwua/dBYcp97Yx/fxvpeG4eCwTlHE8hr6Q
LBmFqk0GAvLHoNFVxBwnrJqsWqy4qCROIglH8ugG3Q3xz8PmC5K9fmGAIqUJm+FU
Josc41yMoY8qG8zvqkIP7ZfBYpCc0dLwnE0waXrkoa8hAhf6D7zQ70e8uiOlUjJ+
reWPq8997Bts+xUYYfYVI0HhKT+an/FYR8lu7Wr6TXHrJyLQrythHjhDuQ0eNrn4
rgKYCcSEE1RkS1yfFBx/3UfiHRWOwjvkZLVbfZwzGkwWjLt0vOvleLmnCwJo2mEQ
evwM5dj0Z1wI4MbztccctvnkxtE7lZHsT9efjPaA52lx1WwHLaQ093t8JGZGwDdN
cfb/+JCGR+JXdEmLwkrZoVxVd8Jf6qC5AY1ZzL025QyRZ8xJIr/p7qzKBc3lCkhP
RA4lphjXh3PnrK594uThIZChspLVC9gOAjq9NsKGGQToGMkJ7W3v9qh4uWcNvi0X
8EHvJ99MmQNQbzKY2VkYyHMyOFF0JASRg4ChtVWHj9oBLGj+4WVgtJG126MlrrcU
GT4S6+DeOmrlTGxBcNqXkaeCjIFcFYy4y9JR731CXFLT/UCfRF8K2KzzgDLg+Dom
mZgw9TbuDSaG9FGCbFqz2pNy9SIdRhof1E07QS/4TFVtg7dnQcvcFfUVeOCTNj02
wFCRXXzmoEmELEY5yo+WutPMFWuCelO2+mkzCWTCpWshnQTNfOwVwTellGCVn6Yt
Zbp5IAU81v10T9rUY9AZrHqFa8E0MNI1PybEWkjm2xDekv83lk2idEwLc9TYsJPJ
6l094Ug+M8MDhLyDw5YGJy48e97mUHWVA1TqcvEBD0bMgt+EM4ITLn27SBjVc0ed
VO2dFft4b+Um11KZQPNfFSI7gbehMkPmJzjUHiAT9saeqYrwl2t6iVz3Y69wxM+H
qXbt30kmAPe3MC2RwwdUH2+T5a88VlmGY2pATuXkarsbjG74Z6Na8cWQjJjVC0A2
bXNqk3hnAAm/YPrwSTWJBLq4YMufP6obz6G6bD0xw1L/Q19k+OFEFbby89jByhQ1
9ZYtXH2pwLOa66UvsInUDQvZisvD8DwWjNMc7V+UjhH/tuo+LutXEj0FD/8hGdjq
cMKIwo2ReufWHPSDm3dzsVhg9XIyaLGfTQ0SOJsVsFmXYbhgcFk4ZrOItq/F3dRP
kI8EcxIhPw18pWtqZD6Q54u/+UODV4lY9ImF+1E8ckA0TftDQCEwLDNFAX/oFMEN
o1QmoG94b62zHPvLmHAZB1jv0ZJDsdWTj0tSIbQQZRStXaJwMnNnmdJD1ryNJWuH
mP+Zp9pnEu8rk52Ccyd9kK56GgTQofW/lu5wo7jZ8eHeftDxnp17aG3273vn/zob
/mBPNZn1CaFPYrbnPXgR8C6kRdfArAL47+25KjKN2OmqRb9CubyQOE8NEctNVdkx
MHBGguIt3kNVs1t8lw2VoWwA2mZLI0B08NUf82VWVe7ag/rYZV/vKeIr9kptzCN/
nt1VcHlMvAP9VrQ5uw+skkTPlxOCf8Dk4/uQ0I1FraQk1WwmtpYUUv4mVXQ1kV3h
mly+De84S60K0g/ERt7t7AmkfxsEZe1bpWQ9zqnHrBjLNjnT0knIqm9zkzgSS7oR
Kd9uZsH4uN1uyIvXoj4oxqquxh8FxLla3PuDM8yqKPtdj/GJZ9iitvjZ237xF2jH
HDhMlZcFMwK+4LmkaI7dXsVQDwZM3HSN1eAEE63W1E9WFCrwxMuq0yzwKtiHQp+2
kFvgXCPMJD3kOZ5QAypEAiYNpc9cNVsFPs9kzfi5EsmBgh9AYPRsFqBSng5uslJ1
UK9PQJcoYqfQ1VQKKBCoOxa4ANc9o5Cs9ooVeM44O19x7QhT8bGDn39IDoFt8G+P
yiXF7MWcfu1ThHC+M9jM5Km9MB10+OYLyAVcGWRIhIZOVwtyy+ac2X/YshHY0XrK
JHIoHGIUacqI353dE/1ybk186dMLAyiw9AE/QtHsDmKas2GMg1ZfMXbvn7JnAEc8
qOY5a+16JNiFH2LMgl4bGt/EJ0jYRr+P3btRzUn2hGWjyLVq11ysF7ChbIbvKfew
BmZA1wZN0E0umqkS8x7q+fFIssfzRBRrMcSKxsoj5uEgfdgboYJsA6N6G4UQ9wVg
Icp4ANUARbxrMCEFRMPBURCE8vlLdxTUB+tRfSSMG5lmPjlf2QimQ7bdSwvLiAtv
xYR+TDPvuqOMNJYkDyqxFan5nHLsX6ntPvbtTd4Ky1+BVBC7pe3MbQfcK+S6bZlN
kXZOx4r6hY4N2Pn4liwaEHnYX3+RAlNeVS78AHlLGHIVIFdWNbzWWa6en4sDp6Be
9pq1X8RULR36KgVrbXIrb3YBxss1YTGeVEvcaFWL+7F046jgglbEG9nboooYBupA
ivyC/asB1IXGdrYpn0xWgewiy7xuEMUiKnPXTuWTZNGmajxHkIgqQpW+Ky4Z/k6F
aypH5oVTLSbA9q5AYNUScneTu1ANwuSvcVgdfCSByyo3Vr702xKBpRvbjwdOLa3e
aeu+rQv1s31IRcLx2TJM7ac82nX6jNJ1yd3tQUWloikw7u5rd3ducLQ7kqKt9IAn
ehJ7aKGCjM0DqXg30KMPgCDkK1Ho2mUf6xK7dRYaOGdKoR23tG2wvUE7h/Hmxyg0
poUXhPFcnp9fp8GVEZTbCutP+aldkySyN83dMsgMsQEiY31NUlLYMah1UjF/6k4S
XqnExb0UgihbBPnYomnffJ99x2VV2Fk6jxQD2yM6MNlhzVtSCXdMsZ9yn7vpKJhM
QaXXxW6DViTcCL1StJsE6qKZ+u500guHOO+Lpd9vg8vtlCgRGAEsVas3gs1oF/nh
D2+pfstW9m47mVYVlp0ZdBHgbY0aehUS3/lxQz42U1vcofHQpOzViNyiL3qHiCGt
5PGgkPQ4rLoj7vVxRnfPk/uga4FEdaeq7Fn1wrS8aP88kHKkzVPz6Onhha3YrpHq
mgKY5+eQ4O+vP2wojQu2Yz6ukTaGiI5keoDXAGIXccaoKHaE/96CH/x8DGICNctq
lQ8k2yKwk7RKGu+JuWAZdG60gMw6PclJ+nst88NWsVKd/R1wQyX4ZgOhEMhoFCT4
SsL6ES8wwibwmP5jW7BQFVFWSLGo5oHi49sEmtkwgK541H5vBzTFgMiE5uqBq64S
NKoLnJuKOFmmgwgDggbRmdHsEg2aJiFCYFHabfp+omqnVS5dDlGyLAPOFJ4Uco1q
QO9X55x2XKB1CLqPhCyMqkLdwXPpN1zMmBat4VNUhsQ9iuxZUipajEYpMeGxttwz
k3tioYGj2M3ZGyWNYRGidXA+Agx25kQw9fDZMehDGoM4/inY0T0L3rg+6ohFzHAc
Zb3CrTJtg2oq7DjVyq4JCQsgin2D0y3CzTGcoctobxEy4xBL0r1uncehtM4I7r1E
s0lE8k+nNt2XLFKrOkCaH4JjJLYgtthZFy9B7+e4/ajaddiEDMn9N3M2XtE3+Nc2
ikPtWWMdcVUyCMvB0O83Ew02MpO/vI1PrS2Pe/MV/l6e/JnKYEJqsHIwWPTjf2xo
zxO/C/DWTOrBBM2XCvBSxVYXQVo1WMhLCjFInyvho2AuXIcBrXI6X4p2XZFlAple
mmrRPJ2chnpb09rkUebhlTlKUhhme9trRt4d/hme4R5X3ZhVr9pnKJ65F7LSMCtj
J41Ehcza7Y5TIBuKrZj1SafGVcw9PtybPmE3LkAM117TioERoGv/8eqnNKthlzXi
56Fa6zGaB3Zn2zEUhBymrlT5TAH7t9xNhDAOMdp6TGaCjxxAytKJwlLm7NambH2/
B4kP/fTuUnLA5Ys+wMqG3W/LnirZXv4PATyH9LB2E1k6/ZZPfH4CRrSkYl5SA5DQ
9YXiM5BVy/UuSaIfKiG7UBF/J3naf6HbfwkmXvckNul19kNtDAXS6bNE0pOvH4iy
fbRFw1t/s+F+t7RPmwfy9mGzx43FgUex45maWbnEnXhar+HWBkXX4RijAMmaQXW0
vpDxp9rmOC+1M48pZHJCkieRhkwYGP5R6qd5tubqOhUMxSaiBciud9VdzrT884gN
YvLhpmmiY1jE7rbXFH/++b1/Ujn5hXDxzbLM2892XBbdW5mVy7x81FX3IUalPQCE
QHbA4Xoq6XfcglkEcNy2LTCGMB9KtF6p0Ucn2cMVw22EBcw8slfslS1r6nBmxnFH
ywFQRzlEgKjP5Pw5Y0YzvICwLiJ7VRr/KuJWj1EXBKmPSvG3E9b/HdtbD6jS5CEG
qJDLeNo/LliyfhSV2O1i5VxLjMwYE6uSjB4boVu4GaS1o6/cxo2JmSk6HQYUcbUZ
p0O9ulzWkjYH7uqvEFEcoHSoyASjKa/PQqjA1ltQQTInlGwswHzq7wTF6xKVNZ++
v2jYdPzQpCqoYgoyzMVCEnmUqgAtuS6EjSO7ctCvbse8RzRWYltwPeZprf9f2KpP
MRkTat3ny8oF5EotNOMF63902r4cLx3GDBwVUwtxKBrz4CPqRjFzRClyqOxuDCLd
eKZaT+YuX8k65tQlUwR9ZcTz18xLzxl3l6VlvQoa7hlT1QH/9Mld8cy35mKkvxEZ
L4B8qDoaCRocegmQcsQtS2GWBjKFC1pjXHdOR6yQeFMJ7E852xDIwNnSUcbo4Bd+
3CL0MPtQHKJIV5duEzKsOcroCdzu4gwqivlGhAWYoAF8r5rrjrC1drb/BwZGjUZc
Z7t5tq2EufMUGoCO6n6NS8OuPeGc8JSuqBCqy3E+HD8be/88UkkBdT0FCd695R8m
ZbifkWtc65LA6gj5Sv3ke8sOn19s/H1xOl/hsZYfliuUgP+Ez5/IhpDyRGHgwVCE
5g2ksXVzzLE9l2PJ2gHoU9hzpXAIIDybEP6PrdILvCZBg984RRSSBAS5wcjVU6iT
Bod/OUUPkc73AB7IX+UPYLA2xYLC2YQWwFjiAnMEpQw/f5sPQnZxGm7jJHOmJuCs
xgMZWTcnxXnWfvKKrgrB75/wkhztbOfMA/0KRfdIfAQWdJ/RRz+0lVoXPOC5vMFr
5SbRWtPJx9JtwCk8+H4nekd3EXuJtivoKujGpXVJ8XXCCJPcfPQxlsMDu/ggA/k2
Vhqn2g4FmOLoc8+GfyemKk4qDDrN5fUyQ+VYxZbT77/JgXgtP7l+Pih1txNnm2JV
82zLDWJstCPln96gLVPerPiRxJcIAoCEjP/6CXmidxdhsgcJHOIrNJBVOyGq6TeC
xGTSKTZQOmeTvfTrh1hrNCt/HrvFTYQKahnCVHHXF8EjU5HONnto4soFkPNfoftE
3pepMiRS4G1YveJ0Vl41yzReiI6WlqxB1+9Uufs0HeT5xO8viNEkqF4YkWsmJqQo
0GSkXpiOT9f9M99uS6Pl3wB2BzQS2dd5NA+E6ki5D3hwL/AxIRDch2+tVY67/l5s
c1ngxCV7fwstakU3tox9mzYVsPFquisgzoJzAX1YDbrKe7EacZczHQGmatMofBqQ
x+abCSgv0aKfZlaFRcHVbk53ShVWGFS1k1tsXTuJ8YXMlygld1daPYjUmhDcWLSD
nY7J6t7KdhrLVjg0qSVV5LyvtX+4Cv/emWJcgwe/ymeJRZDLym55BgXA2t/no+hD
14rwjmFoWxtlRfdQwpRfc0a5YJ5Gj9GBUFhFkdAlptjiMC+8wA3d0RdLimb5adX9
J2X2Ys+aeLMPy3c3QHlSB5jhATUyCt7H8+IHoIqmFW/5UxF5mVGepNWN4jRsO4eZ
HOQ2XFBmnbaEoHyIVpG/f/pX0ZCeA4gR+jigiRjzyPpXVj6fl8/ev8h0V514EIzt
1pPWZTcbWEQlSX7zjJ+iXXQlgiXK3OBkBkWJAbYG7TQi9zy3HKrkFhzkW6NBf91n
OuNqVDV9R27tHLgFabp1Os5z3VbCz+uV3QVxTgZD476QQNio59OnPHJIiHrQdLV5
nOyKojWCqsxS4RXY39mLGhUHRHVCojrgLVegRNF9BInHCk/DN04K94fDNniHxVLH
8/dxAH5JpZX2r4h0AOLqsgBQqsOGyr5SaZwBvMUGZRrbUesVRJYXF2Qg2IhA6QoB
3cT3uxXa7H3eG3R6cbriLudgBfZNo5GfBnXkuRGbZHBtNY4A4XZWNCocz7PgHcqq
gNz+JvnqOwBkq6R0T/HKdXKnZYWLe+v7+4QTuSD+JubummqqVO73YI541p4nxIn9
2FFizloOzVOpXfsUq1mpPyLPu7EEvzAud7nMClTU9iuU+tcSN3i91IASn91FLVKr
HLsX7PX1TRyQULxUh4MURXYH3Lb5Ipr6EkvkgSu4Z3lBhXItArgr6lIezy8HKZhS
yPUTi5lphdb9NJKoICe0smx35kbBmNa+IFpP6t+wqsdkMAOu4F0C5XSopkWmj4dA
4zVoRZ4LEgRL8u2GgmzFf6fKZf9HHyrq3mZ+PGxwe788AS7shPBjLfSpmJ8w+k0t
s6pkbe3cw2N/jcaPCfpS/IK+d+hZg2pv1IvnEX3cy4mGI6Cs1D88xlJ2qea58PS3
3urQRnGfuMBHSWPZtZxYvDMiYaYoXbuWTKWeCZPcUzB4ThynOIuHliMjIDOwIUkz
dBv4WIiBct1ozAy3mWc6EsdxG6HJFjl+qF8ZEQRAE7jnH02TT5rYSKI1DM+AXBM3
cePw5UdVrVe3Yyg8/puckVdx2hCQwR914tgQxjXhUdFHBUgSqIF8SQMCuoe2cnYd
xX1ob1rtMmbnFAJMjLUazCtyhMTQyW2QuPb6Fg+tt5zOXyUfWu16QFmzHR9UdE8d
wcGqdy/cfjo/csaA4DwEKhgzk6HVEZVMV7xVpobzee3VGwVy5SqOlRkzWeqbogbZ
49uD1UwwmbxbexJczHl00xp7iYxXgzdFSu7RKR/ChGmW1fHS43eyuVMTFNxY+R3d
oB41xizEXWfDK5r1aAlYN6RGeyYkNRtVjIDcb2OICF+keZsnN35R6JPVlcNSvZYx
b0Gt4V1w61uRA3XoZwJi4HNAqNkvctiKozs/GtAKHwsc6DCBcpRT3vYYu4sWITFn
VVQb2FaLZGXe5alhvkR5b12Tmd8qdz8f/SbIeRGubMv15DcxqCvVh9I0F1uY+et6
MVC6SkI4NaeYij4QrvpA1OAiOfgdptXSC+XtvFATr1RoskxtolUTzCxS2EdbAV02
T7X7WDF1P7hoYQ5SQAYdd7c6J5TFRPVQ0MLL+dMJW3aBGHXK+QI+f5HT3yqo3Uma
XArNCCvjAWZIuFKaRIWMoCuxf38aLaYqTq3UcWqZ/5ctxzsb7ibbwr9JHttiHSC2
4aSfG/uEuVMdl0Fta+BtHvuW/tzSpgQAptBo3Rw/2lIOj/CXYNABsgTYG3/ofr0P
h9MgjZbe2y7nr+jhISk+3RRuJoFCj/Vdc6DArzDbqsLFJOySb5myOD4WHIu7RZJt
T5+xZKtohAeIqyjSBfKmOcGjko4VAxhXqPn2XdPQM0DmtIC+9t++3baWdQsKL3LS
S6jeaOqN1Z94yVZriQWzsCdm2NolYzAJSV0IT+bt16flUUoz4M/aVsU5HeGIzqsT
iX0GgfYKasjR4hhCxd+wZmfwZ9X1H9BJbIPVEpZ/znSw/yh5nQ0D2KgGmaf4Mwvn
HFO8zLtHgnRrPFhgJyzokNrjQWmQdDauiJUXL6Ky3IOsbllyOaZ1UVqysHxzxR5W
409FWz7FnpBswIrgH64Uh2Nzcf3wzt1BMDisZ1o9j9fLCCGD2QRBT0p6S2fiUPKN
7+Y0TYr9KQ5yv78hzgtADgHb4+MymQBZ1209qUcsHwL1WLLehB8zSCDvtiSfcaBj
B47+O+6huFDoNQTzPb8HiarZXblDGHkJmCx+R1QJxw4SNfcUDrUHlap/sh90cYUE
IKAUjmDat9/fiIVSdjxV7B0UefD1hFZZaKu++tBSTBiCLVMHZ78Ac6p2jNKdb8lA
uEcFORPZO6m2PqvsDCAHmsFjgeVMjJvRpCf1B1DdBIQjmaavMHOgaWVPBiJ1y03O
+DC5MsoKxDFfqq5j0lNKJTT2nmTmv4s28+n0fMuGfqASaj9qs4u77h68dHYxrwel
V8XpJ6o53y/O2ANCjsneA04qORY+svpFC8PvjeilBXV9yNcNqMHkjeWCjisRru+Q
gvvdQeCCd4hhvKrSYsosz2gV+saY9ejsG5Nr9g4vtde3JgZAi2rWzP5x7QKxUhh5
sTc3B0PIj41gufUskS1CgMxCDXzLIGsO29u/PYLiA7yC2WJBC4AInhn26aAlVt7T
cy8BETeiQkkxBn0ticZVrcN41uVhVX1wJqaMZi3prsb4LmOdQdp5EtmXlMn6wqMf
nEf9X83JApSJbHKpel9zkyedLmxtohp+4v0b2myFHsFKO0q+3sbxNV8O6yVcOuQL
zHq1d4P50LuDij6/xC9DaotcF6ppCTqW2Aoq3tUiXwE8T09z0qRAQXsIvUB0eNyI
CSrQnf/8gZCetKjVZ/xN3XrSljRCgho1/ymW1MAlt03TcZSSkJG9d8GaCtzdHUIA
UF181Sx8lCsS58QDvdEZAj+2DV7OaVGsIHSOsHppASVpQ1e/4YcI7SRyzUj8zMwi
vBxG4FBVqkXBrKDUniiRiHr5PFpMagL1HHkyEs05NbL33ul608ceK+t+7ukxiXDB
KFPDiWqBoetefhFDUzOpTCnZqd4f8LtHuiZCvEdR/8llqprKv8iWNReWko4gIuHz
Bkz3Em1F8zdHsYtr4cSjbAdLG4Z1hDu/QPbLl3gWwx369CyDs0Q4N6ZRvfO0sY/s
NmS79xuj+LqDFWWftFS4MkeyWbrmOgw7eJmpv9CLAs5tO3EvPoiiWLStop0mZeYE
ImYaZjohumz8NQBAOpiotX2ZyvIWcHAgMqqBsrvesi0d34k8TptldkFBTjqxkavt
FWH6Cwh5Fws022/f8cYkzym9kDj2CK8+U8Oaht5h77KyWwsgDd/+ZCZsBINjr+jn
JggK9/XeY7d2bQkJKKH6u8hn1haqeQzxTNKBIw4kfIo65wyEsnVMZtdMddXGlG2f
D7Hzu0Cfd5YO+Yh+TiqEo2gSwYyDRq0q4osNm9HkBiLi8Gk1w8EA0XiYjWMm0On4
vgP9c8VItngLKBrolUfr0iaizXHL63Ol6NpXS2HwJn3Rvo0Dt0XKc0HFePLx82I+
m9g8jGqi+ZjR2CdaM46rhxSqByiWLpCiPQu19GxBf3SyeaF+Btjw5hXU1G7vLO5h
548Xyu3fqQfCvOOqFlieoVjwBbfKxPXhzebl+Y29KS+5IPUAfRczW9OgIe4Pjp1w
o/cVeEkRLxUmBpqmdjP1088EY0m3uzQZAetRyCDgqlKB4qAprTB3jeV5MYxLl6ip
lg612QaReg2d6s+9b4in1RtR99RnRyTk+5SxyQKhUNmCPZ2392xa30quzHadxGN0
2hiLpCpLayAoyZnTjzNizJX0hfTGbNQhWd4IT7Nba6pF+ZrNEE9qFR+4+l5/LReU
9xcpQh2OAg/l1dFWuZVXlzwamBlDvqoTSyBa0P8GAdi5hMRfJNaxtGhUO88hpiKf
gzcm3URQrlXsx3ToLHfDzRNEcNYjK94Lfi/B8WKViemhzWgrOc7+LFPIXumgjCFW
YLfLj5rrbHYyD+bZP3euxBmPJcjjC/3TowU7HwXP8j01JwxaL7nn9xpAhAXpWY4T
hAh/+rdO1+FK1cyCzrCcHnizg7U1LsJTT7uRImKyxhkvuMq805LogCGBJyniJ1XS
qcAO3QLPxp5lILoPxdE2ywGL5fW13aOXpY/wAqEsqDH7qAuLMDowNGBwzocqqAJA
Yj8IIMwtn7IJbkdL4fKgmN7JpOr4v6cDwYCTbteOcxa6H6a1ocX1BFKWjWiTLfxa
8I+kSeo/hhxMRGiXOm+GOUu/LGPaH77pQr+lLUZ79fQFzI7oQMLaO2SKt8rMpQXh
jKz1m8CkGl/O0VwOPl+eiuqIrwhkC7eONaUGRY0JMjnjuqdvkXVyJowxHxLCOEJa
uDxHzmP/BEkAw71iEjgxjVTdBIF8My3ygYMOjtN1wsL/jv+LoaXl1EqjeJyq3SYg
pPTqxoavdhkPNfL0zeMxwwdrxR2HSWBdOx2FHRPKzK16oouSRH81OZohbiWOExQ9
qKPqwAVyC3xwVCVrC2fwWsmm++q3vs9kB2Xg/jvj+QlSBw3PAl2+zoceeGRpxNwL
kcRcuUdS5M/lTa5b8Mds1xT5bfClue2JO5/0GyLqpSImp7ProO3/vGcsXJynsrTw
KYIKBGHnW3fMZq7mmd+aVPNuC6+Ql1GUCCnpCIMucWvuCdpfJ78/oseX9FaV9cSl
jRNqsSZOT8P/dwkVtNEGAi4gheg7IYwAhVuvM96ExBySyWErvbx9THlXXPWUv4mU
pm7STgH5WCzbaIGhC53yXqP1LCo04QHCDCXjTYjG30FQOzVU40jyuK4NkN/0rAQh
cPTdOStCEonyiHJs4PgE2ZvoxLV2VyEP8dUdm7ZwQfdy8f7ygKGMGzEKmfIyB0hw
HEKTjC/CWwfXyN2R7e6CXDN0El7jMsxUKZltMeiEUuq/Kc2HuNDgVFR/OCR+cTRh
ECgMASJ6fiqpXNfPCMQp/AXevaA3y8qghSTthBR4LNYDhB1HvFKeX2NTsTnVfA3X
5LyF/rfuixVO4ocntWV0nnvR33dt4pvLDN+BgGZbxt80mpNDVjqYivdjC9w5kWOO
ZMCZlVA5gPglhHpC1PSGgIOq0rE6JJfpxevV3sl4s+BfwKxP5vZ7bs8KXTQr+4c2
neqEFkJwo1cg/FLEE2q0o5LkBh5Nkp0Kh7qFJWc2mFmjQc772sKnPw84OQXAYStA
mpHYlt665AIizmXGlxZarUMeOSTqsXG+Swg9nxoMQcLElqIl3jVpKUXqQ8gcdada
fNrSYeGIgyeVYlLw6hhn2kvOYFNkqkz38WZFmLZ+/G5k7q49UpGAtg2tc53oXh6K
X/sh29e+xV/r0Z3QZtGVgTy6+N8VMv76qPxq31UVv4Gd2OEtL+yylw5mUPqbGANY
tZo1VtyNbs6LrCY81un13gMGh3zrWdHPcw4QVo5tws9NeZbQqs7+cYLoxrI54IN3
qgxnCU8atMSJPDh9KAK+ugYdo0WpfBQ/DdGHGVmivqc/wkAJkW3rb2Vp0UbMrwo8
OIwNVeHwjcFMCbDUeQENNrMai3aJgTLCwhyXwV1nBfvq+WFgonkmScikeRkNSRBa
1dvuyodboH0Y/hfgXjWgGmUqk7HbaJ7B5GMnQEw3WEyY5xF5Gtz5mv+aabmi1wQj
RUGVVWT93TcEBnSYKHdruys9p6dC1jAEgBZgCnNu8iccHLsDciiPRPC3RK3T6Db0
OJ3pGm76igopUIOREByxTIIdO/zfWD3T7tMt5JMtFZ3t2j7R2hv08h9O0cQET8F1
7eZKYvKl+3dDaAJFR6p+o3sBEVV8p1Szb6qTcf18bjiKSLoNB2NO0895UIWnBGvg
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
CSThiVodmwfch8nDqLnt+Uelhw079wPux/aGov81YRJJu+WCd49VbdnCAS+vuUmU
H2Q/BHCEXXioXzZIYYzoW+bBsgHiaQMEv+sAOX7lTjs1IZExNFDKDYjh+WL+dY4S
VTSLKcpVlHAmLOKvojGKxFQs7oneGbe5LuJl/rnPP+BseAZ4E6whmZ0zsWLTWcK0
AtiPJ1RbfWSJ5yh5f5jvZOXSwcRPDhs433nIn1JrhxH8yl0QTgXCDBfUBI7Ug+Cb
kNJymG8KC2M4SvDdVp4gnuRjRkOEsysxA2K3xe3BD5jIRrguJnHyp2/1hXj7UROs
/zLWdxuCtqLlzJFjNyck0w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1200 )
`pragma protect data_block
NZKR6cN685zr/pY2WXJshUNTLbcsxejAd5XWuChbnnpUtkXSQBbLyVPZi+wfCTGZ
f/bE71761JkX/x39cJU5TJC01XbwwwwkzDkLW0NOB3g+YGzFKT0EgecGQ5jtE8IK
EvXedDJGgQj6Q7Zy/XQJlcch6F21KRITMWlJbV2Rwo3t6k4FEzvkLpjDP10v9MMV
67Wzimhp+T0c/OzsRCA0mgn/krLSBjAoojbgv2+yVPG0IOQuy4zMrgkiU/XrBA5i
mVfBiXqjXtXsMYxtS/Rjnmfn4nMyHVKdyrAbqtd/2VGC0gEqy93x9wFe1f3r+jq9
2f1oTFb6Nqry06g11cTIborElkbOPEqOj30KkpRqzRokYU3RzDcFuHXI5Ko6eGiv
xpCRDA932av8D2BDgmNrg/vee+bJqMTw4LSpChDUs1DdsCsVwgRIvaAUCxQkuYWd
X8o71ZnzyyrU7+TRqglmTPDpinHf03l5UvjwgSqk8DH96bK5Gvdocn410P8niNgs
QWD6enF4g/+8QlT9UeA7fp74RKroc1QgOTda16T2oZoieuIlkQetrKHP1SgVsMAt
avSQHEx19n+sYklfwE+FFkt0MY62NscFXilj5eEHp/q6wWr4kkSesUjR03BT889B
5/R/fItm6bxTop5cXYrtfSFtnZI4ztrP244C1CjxamchChv0CqOzDHT0XUErAsP2
HeJmodHMGzrWWiAEXq4jg6+I/8w7zXGM33VYcsY5yZRr0aEk3TjNgcN+E9D7x+d7
YUYwqo/Er77jKO7Evb3ATBOjm6oeEQENHK5eSXvgyH2CDSJjMfEUwmHJlSWsVRGs
2gRCqkNkA/1vhEiImyh5QX7h+MOeeWPTYM0ZCEUBgswB4ZWQT/js3DdBaVKsgvr+
h+nN9G1p+ThvIRRsHvI1aVWVkSaoBw9844bhlDL16xCRtrlVEF4MBuVPFpKSuAgD
jnzAg8ia0uGOKtUCxmMpD+QWh9bTeE+KKTQTLBCpK7cQemIX4vjBuNN1UC/SmaBn
Zfc0TlrQnSG7X77oVBSwdAJZSfD+hgbDBE1D9HXZPSngORA01rBvsHoryJPoYcfP
1p5siq484AMc/+iprRDTxT7/Kl54f3aSjzxfW1hlNRrNVIY96E6GRkei8CqMPs1F
auBvBf9Eownm1SpAW9zeeHtfbZGKgYZOiUOFZtsYIwFK7Eh9WptkDIrS/1MMkvKk
cK2nhf4CiFIiPTrlDBqf+PTF0f/iu+WzLeMwd6q8miYU+WqNB2v+t5mKxCh2kbmP
9KzGeUCh9imauyXdXjl22XO4Z07biexzGEbmbuWNKgBvXVASVy/8T29yJ3GwxjKe
nnN7MxzfaB3eNe2zIZphNwaRYTYaUyilkUgnyqYq5y3+GQUn+MGMFY2BGf1RhK2F
1xn5N39v+932tVSK4JXvYfJjLyVsKVbBkW/foJLY6WPB7TL4YchU3pkVj2yIpPWl
Y3gtGZpfkskvGxtEYZNUayHF6cb+OgJ39sZSM9mmVTGF+HIttT2+vPLcT2Fvx4Ax
OuY5U072iDxyz2Sg3T+y+xQG0fg9gB9A+rBs7yHYCkwWsP4zbxjewTD0lnzF2dYN
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Pxgkn6aOMcuGAlw3myFIhgXpRSvzuyQwWekGMXKsRWYyNOXe/pcc834iZT7cxOzx
UslFj2OPXILTIVO5VPuEZjdlStARC8QSEfiEytSsG1bnd9bUMjTtWFg9ZPW+MCB3
f/reJKx67Gtyt6FBVQMA2120rOPXpKbTC+tCa+VIOD3W+6gc9tx5nQ5Js/Hf1dkf
c+VpXV+tE2YkN2BptKjJr+tKOskBeP1lyyvAvzQAeoLmiKJ7XMBQ+zGp7GXEnPeB
uZFsuIwBn9Ai/UqJmOnH3fhwJ5lEb0V4pyA+LJc0ffvt05wDNELpWWKr0VDpV1Qt
hYW76TkvTr4fSRa9AUHblw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4672 )
`pragma protect data_block
h4o640YNrYmiWmrU2wpCwFXrb13Lr9ZU6yQ1n2M+sFcKC7J38uQYrDn7sQNMOTVL
TZgB1QGsI57Yu6W6OZ6MNG2wzRrHcQdKD5SyOGssB+mOijpBI1Yhj6uF+JmRfjwd
wiBf7W1D8cHQsdKxe7Hs/FYlTiiBgGlEyGJetZNkYJ2eI2LP6Kx+/9EvGO1SG2tg
LU0UDVc3bUF23+LohgwPm/IdUQ63mjP8nCgZ/mGiNmmwT6SWDFE+g++Wfs/cKbK0
NcAS8ZBLIBlsLSuFJ9dbkuLHWvu+ibAJZNsal1wlVh4dekL0UvYPCBpdJ5kgmInu
M7wWP1/SA9UVtlU6zNA43vLI0Sc2EdZBwASelfF6lZoSnVWWxk90nbiPwibWrrQ6
bOKnNKtnUh2AYbHESVHdsQzCv5AfWXq5NxDaUBicw8isDcjTRhHiNhvR7TKcY4Qp
TzzFQ4QwRWnplEFH1GfeUqm3GigXOfevxt0wOjGQ6PKxEOpgAtOYIDGljkdd9/h5
70CKaSMHItGd/hRFQEgoG+RhRnmKZXCwSu1lmtD1S883peCm0Jsc1wK48YMczd15
24yNKYGxERRwPwM4YjOdJBd/SK62UrVKX7cIkZb7D285Pb186qmmXGqbcRnm+Ycn
qNZylQo/4WNW5Bup3RGSLSF5WlvbPc+mbFPxFJGAvMseV7ghX2mOuM1wybk+8cjx
ZI/TLaWL7T0ZysC34GRBKqr4Q6WgUkmPxhA52ILCVpgCfXlJHLC5G7WBJGauAo1a
aFr2G6SCRQS+frTCqEc0Cf1vR8+PJZf9Dmi4Z+tN/fw+7JkzMTSA2Oc2hApn1q/R
nJdkUK6O54aTgyUki1OEj5SnJWmR2zzlkZLy41Y91+U9YYd8gTli8ZxZVezpJ5Dz
A+hzAiu8bBAxR3tntrvY5lbP4lyw/YJMr9z8qP8FeoAaF4g5NK5iRTDXObjZHdCF
3tjEBXrcAiM8xgswQ8xojoCSdiO6Oickuse89L3pPy3olXW89sl+A4L/mUoON9E6
fQtbrmTxM5qTB9is3vmFlKmGVr6rUn+xagfbOPWEqxS2FPAssZjY1MmDetaivAFZ
JooWph1c4ZqoKYH5oEuLggVz6pVUbaie/KS+DIhvi9jVxz375Qz+YIPmYpo4N+9k
LX8q/Z6oNUudbFYIaieZmB1c5Z+jh7GZF4BXRArmWqYN2rO3cXtWIqheDJwsPIpJ
pWznjjB2ZI24UyZvOWcV8n3yaXQlzD0ZAe15leEwkDWJJ0FjoT69X8y7SGVGzqUI
Sw/F+BXaRmAcfUZOkIXWGFuOwS6Q8t7hc5z6Jeob3BbeMrOrUaMvddfzKnITZqES
QiMFgKrrCbbIHizLq+Kjm6A2I9OHFuoxmnrrCfw1STPQfM5sahkSuZ0YYz982SN7
ZZ3gfLJ29ZdfYqUN0gA092T8t/VUz2sEsq7YR3YkpKGhj3aQZCwug4eb4plXoEVB
hFv6Kdk7IIb3kvc4Eiks1t1ch3/2BGZaBpun95x/lO8d+vMiUpTrcrz3XPgCvzWv
WnCqLBZGAeLcIP53VnQdOey4Wak5BSdPf3IcuEDILGu1WUDhQruvaV6arNjCm5iM
W0RCyoChvl3H0Qkimi9IqPA247w5+21OK4eG0M8AYzEiaH0R1aZkd7Tio+GLQL6F
P319VukkXACZDlbxvLDYuVy3zCzTpZwwdiA63fp/vCStMlhJezPYZw1LWOJp8M7p
ElEtRuzhVlYs9lCuYNB3fEc26VFnEbMI6yhbBt6DgEUKtYRTuLbsOhv66NLLxb5K
jHxHIDHWRrSm0gUedhhM1qiaBb3mRSUB1ldJ1cdqG9V/rfMgFzBZZzyuF69+yuYW
SHU4a9Bd/lDejCIgMljxBZ2ASKLLsXR7MAnb9/97AoLBJKm940Y9xaGqmgSzh1Cs
60nF1P4gjvCJMqJJ4G5buJVlNfo51pTw0ObQYBxIHs5SEdqdlkVhVKo/+E7Zrl3o
jF/9+PLF2CT3FalL+G3oeqZN/6vRMXZK+wBjVIm6MP9hGCd/e/ko1qefOUvh870F
5OAG6xn6dB01geGnbQ3Ntye2qbTl2x0O8+OQH9YJ8o6gBN1GLkk93rljJTtVnVmY
GWU+SXHyyyx1Ii6OaftNhl/rV8VKxutsTCOVccuabAP4YK2/ZLyKWd6oXuWuTNiq
/Wg+44GEvCH3+P0KHfzckaHwWlFzOQJX2jFj3L8U5mLVgzTn0/BBpiZ58HD4bcx3
xgFSbY4cfo36nDN+5KtqhL4nQ11cJ3r4u+kXODZHFDwAsXbc5TqhmoyvOh9OAtxX
GGu3U4AzQvlrG8tNN0eCEjq5NjZZfQwzm5r5bY6AVtI656U1B6PFQnVA0iv07jhC
McKO3+Wjocd755SQMiKYP1FhkK7PqlnM/5xR1R2jN7Zg+eIW/sXI03v7noFTVvAm
j5Myu9/8lIUdNCfVffwGqFMEBaXHszVe3D5Iz7y7VWJUTrQu/2hzzpJNSPgAB2GB
mTc1xUKPjf+f9IHHAyiWpniipwe3IokeUeubSxmSxio4x0kVRqBr4u6vGvBa8pIh
k4zHkJDqppEd/PrjQneOAeDoD2YfvhsBu3TQNs2s9WhM2RZ7fFfuUcWtdh5P4+Ed
NcYEbQo1FNzhXbV1SUJ+6Df9XcAIK2G/2BSNk9ZxIo0UE/h8YL6qJ8Oi5wOC0OlZ
GaFL75X7FaqyfdLgYtlzc2VoEcVNulenkuE5hRi4acV4nvO+TgF9ewx0Q+MSuGJ6
CzR9kAaDMRKZJt8NCRwz7lZLk0m7dssdF8eAYRfIxH1ceGlH5hOevegVsCtat3zU
HWktTtPRNjhvSDMqns+5Zn9t2KNy0L0LKVp39rPxbYvBM2yABtS6Sr07tsoPhpr0
i70QpoB2FP0jDFU3+G2A9iUMrXb6aO/d5NXG2GXzn6xXQ57d/HWTwz7uVbsc1zdX
vzmmsmkKrra/5w8GHpbyjC1lS87mDGv6Sq4RSwJqGCcHhpCmLCWwU9JLNnzXaZBD
oXZceCGxYgEZgFzzDmCdTf9Tgj3LDW2ZI0ZroLJQff/XPkK1MpIIl88nmSLq/uPZ
V6ASfCSH6vtDbtVHd1DgytFpAPeckk3YpjUCi9Q9wiYwP4tsORb7JNf5mKJvK1ya
dgsV4KHEJbXR0c/fElcrQZLgWXcVCKp5/hE1C+vbG3dkawIPlNkn+o7lTS9e6TDM
TZaXDep4uxUL6CYac0iYStxVQrE1w+/iBkX3lLXFBadWZfHOtvQ1NObX43rVEYRQ
f56jY8p+Bl1OtJnxRt3WuvLzwizuP9WByFhGnQQ7XpKhuCT2dkUFFz1gXttfzhX5
HUiP21n2yxGFm8cs2sCphvAbUyJ38ijs3IsfTZJjHQr4RKUzQ4PFn3y6ItHVM9Yd
ebzhqjln3NT0Z/9HUOI4W5AMMjcB2jIFpBanMNAZdo/nSJrWdyT1CFRGDYwm+e/E
sdKKcUm/gewgsywK+bfUwc539A9PEwhAwF57xjdESRBtOw3BzWnQjWjW1Y3IHF2Z
WinkBw3fqOtpVagzKKpckKYRFJLIORPEH6e0UbvH6xNeDyDh6b2kwssMxbK4bqIC
y6i9NXzVnOyIeT0zyZ5PjUT+dWDngeHMtk4O2ljupJ+TwS+GUe3CG/0KkgHs+WA7
3owPjOmDqTo2e19QgezS4VPraABQHKBFyK/KILD1sfP3bLYqgarkXh52Gver9fIF
eHxM3srwriuQ0Df5uxsXtP2gbkZ/oxPZfDklkdlLigaLIRtYa38/oShHvBlQZhXU
EPQrhLuaQlQsRBKofpcBnpj4DDxwAqKNUkCbsVyjhofg7Cft/g0cKoSyfZLCwo2o
TCT03cs/+U86peZV6hCqvnidmfF1ykKXUbfvuT8E1r0ID++tvvkWR4LlaG5h464S
bvn7DgU0aArc1fYp2Zw7DLqUUvXHed1uqhvzkxlc1Xj9b6HG6vjmwHLiCwDoQaJ2
40S7JTHeAZQnGrKUnA3Hwx0ixuWHP1+8CMN/OVD8MVbUbBUo2/Lh3881oSdT+I9O
uh/NhV+7hqyRj3ltNnOKUIpXfTeZ8/S62OuuL4jYEzCEMWYHXAbO8WnmxZv7TSpA
yB6E1lH53/o44H4PWURTSxl/9UhBvHUqZBhnw0fLKZAy8r3HUNxIWV1jPyl4brJf
HK9/2IUxq2OyJoE/eGvAC9JnBZyAp7Ua8S3K7dIjdZMVRiA/7Xlq33c8Mny/SdUb
rGH+xd0akzNTEZcy5rFq14qJMwlQvgQmYugW5JZE+IVb+ACJJH6Mbb1BkaBnOQI8
hWAWCjJ4L+mU1DIMAWu1NtKugGKgP433BNkD6iOm35zJnxRjmAJBHGnnCRRJEyEH
HqMEhgnGeQ8SjcOXA/FUSgL9NAQOO2bu5xEEgR5x7xdlRbhC4DrJRJAiiO72jbWM
HQF1LPcI1Rp8lvFtYd1kTNNKLHwWGAfVl960wOvWJEimh+yuNdU9Q/yQvDKg/Tlm
AXIjHMP/wEvFE+aFq9220ck1xH6yBnBEe+pLN/YetXdIDjwd7ifDf33l9xxwL2Zw
AJUiUrr0A/bbbFg9QGUG1aGryYhl9nb4udqjlZf8LEx040PY59i8eTQkQugy/FCr
N2GkZ/CrzgNXoGcMR8mSatM4rQt96bjUwMTnvXPZTXnWAR+sNWh6oVqD1KAujTQN
OtjRmwP9zP0olV0ZnI+39KMi9lpgQ7E0M9WTpcSHqGuvB6fm7qbZ/NAd1XyT337o
tmuMWN71WiJeFwMxd0BISuf9AkXJU8P5HeE88n5CH2C5BzseZhUDHIQmVRAv3cvk
OySTFdcVJ4Ag9sz6jGSbB4kMdUwzFEs+9fEJXxpokAYDfWqBr2kKnVMsa578s42w
ZoypWY/GzZOwrOyeEUPL2LjQ7H39HHKI9K6OxjRFqs8xuq5zN2O+auyQE3JT4981
8uIRnhjY+Yf9xL0CqsnSus5rekHncAuSzz+oeNV80AlAIPJ4cVczgu0yy2aKjVKR
BmCGL904/Ek79SCAhiCsnYpJfeFkU1IWVCUKCfET62Xmxm5LvUgONi4GD5m/bfqN
h9ekedWIOwhC4pZnY6V00sKSpfXXbZTANKd8NtOXE+kd/hqep/ms76oiDtNH8ZU8
3eFWkxuki4qym5dYm4sg99d7TSZ6pYE1E2u2pVFwqZIdeaVy53VF30XnIYma1M20
5ws1uDxQsDsWmqpuzCk8y6n/BT/ck7z0MxiGwgTMlrjPdfVe5j5kjNN5HwLWQUeJ
gH2rHRpKU+22SniAtw6Umuf12uuAuUj0gP6o4QK5xo8L3k3FySskJarK/WiGdjDD
P4lAAUjHiyFXeAEXl149RAVCS20JrfGlXWRlpTNFofxH8sQRB4ol6dFIiAfSUp31
eRhD07QQegH4nI+9WcDcXDkH7cF71BzYe5X0Z5uk2Wt6Rs5W+hhz+Wtyvqdv6752
YKYL7ocGLYCUjDbcV8hB5s2VUgenHPFyoOx4cF3GouJEXJjV3jx03o3pISfmqFaH
5/POvtB48ouM0w8vnCqPebpBpamyij5u33khM0iZ4NDXtVPsfmCOVBgXShmMsX8e
1VeLzOa7NuZkVhgBzXJB+DRnuE7U4oWD8C5acaqFW+uQHAHI8AJUoYRjKd+SEwkZ
NEA2Sx6uqJgcKuDIiano+uCt1TGku/xikOHmTjQYXeF+jxTYoBjMZxUgG5579+6q
cBZhULN1QIILw8i8vy8VrI28L6Gik1pONuLRbiflOdlIrBQlk5Ij1FGTSEosb/2/
sxn+4xhn4+z06Dv67YZ0lFpFrylQdkOZheYM9pefziygqiXHq8YJHXEa1inMR1cJ
XV27bhEOU3/3K4uJEVGZC979gXf4/rmn4PVqqu0IBhsfJffPpRY5ewBA1fZd+cL6
rYCfilgey5Ctzw//Z44Kmq1cHUx9d8vDXBDpILAq26q1nlnTbNkDF+frtHfVdrRY
vyETiySxN327IOckAIZUG2iYY9GxClZA0ZkIDCi/C2ZpbmTuzYOrymH337zy13gN
bfikzZe4RxIvRORXnMUdNuiVTGPXl6vcr62A/caCCw1xJKF0uUSy3+FYTPmpVwFA
VyNHE1iXmu97quaTp53jJWPgCrF5YECA6gnmAo3IRdW/7CjSfJUDzoQSGAFgW28Z
I4ZqTR8BsSNQHVIU7TOyKXproyBosXTpvuH79PGes056i7Q5bgDyOeUWj0AjZh/+
cbUojlgzNRnUszHsga3tZw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
apblSJ6YBRU9rmOsVn5+u4HyYOW8oD4mNp00oLMHJiyk2QU9kTR/cWtyczKK5CA9
Xcp6vK9K+Z0mMyKUngTLH/v06tdMo0+OuJODxclnnt3UDVDRJtNdUtMoIOyZK79A
K08xd1ahy0M8bbgg5K7KV2KN1wOD5FgP8llzEOCC196RkWAtmBa/gw/aOuRGazoU
fxaIrxF0Jv//qVgBaln7dMMbuB0DguwtagYCZscl4vJhQ+PiD2C9th4VQyEcIYJu
ZdPqb6tmUg+hNZ5kjqYJgE0V8UArJ6KuvNNBt/fy6iuiIwj+IifQUKW9a6J60GSR
V6EgsgwUrR3K9XR+E3oaTA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9344 )
`pragma protect data_block
fpqePilvPxdMVyVOyYQFkc+nTSYIf8tltNItuIHkygE614zKG7piuEOoFV+Kn7uH
rjhoXPNzB41TbZNeaeCNSrtGgsXn//HkpbWzN+dYLpOaNgWiuwCzBlmE7IDcfs4l
xabGO5mcAf7gGr+JkNIHIU0KXLOSjAIcWBarGH4aptz5OFjDNCT9+MpfI7xpwtM/
16QuoBjCOZ4C3ia5q2Pd9Ec6ggmrNyHR1WmzDrihxSTO9CCkScVoHZXtwX1RGCl6
7vEZuNbHKljvVoly/5E/bRIPQOIli5m2oInLVUBCrs/uXj8Dkb9GEQDqI+JAmSeV
M/b6zwFznE2NQeghJW7SR/ECDgIaMBpY1vveut8MgX2CaIv6yHu6KLs2jskawggH
Mso4WeU+UtPxKz9x71Hk+vxuzUQbL74cWlXTWTLahCH4IAurCQTiLL3nYuLg0SPZ
erjrLi29GZhRrMsihkkbaPAiUT0zAvRvJkHize/+7rUKxbFLG81R87ff0H6f5C4B
gWBjgUsefPrbzTt8C2bTje/JvhbfrKhe9jdb00ioaAX5MpFTVpK1bxjb++A+Rt5s
T+mkCpuOHbP9MBUd5J06eke7XkS+Eo+syuJoQZg4gxnGuoP8ubjbYr5CuhG4EWAC
d0e6B318k+SsR9sSjtyAIUf0q32AWebZe+L197RisAW0Ban1ERyJ1GwiL/UM5fn3
sQ6oFxccIUBAgoiIk6vRk8dWQL9/u7LvBNz5NXdhB0usQ5w9Ht7UNLI8DCxXbqdR
5RhZNbhP37wrerH4CpwitMIEV0etBkEzcYPEVyVTiS0e5r/k/50crCN7ZZJ0siO8
cTBMrv/hRO3jmDkTBhs38qn746Z5h5fzZu7oESd0zHh3PeZFj0aSpQcWHYxTkV8P
wOUvkBsCRomHIbXsbKtuUrtAGTx6eU6rzzU1sB1ttpPmCHB7ZJHhkyLSseaDrrLd
NrLPU8ChUb4FVxMV/0WOE0Hd87h3zQ+uQvyf1sx6JPzz8Qe5wm1847YG5f/hnphJ
CRsd7xoHfVjYdEETtXSamvt+FIwDP2RHNBN0wSuVjwnjC7hV9uj65fSVrWg47bib
euRGA6I4ztXeN+VrpSN8eJrNYttZfip39EJxlPDtIGYsPQ3l06YF5l3Fg3Q1oXne
pfpaoRlViz/i+ghAg8mfE58i/NFtbDKx4NBjOQsqxtd8zdY4guATGI8nBGKe6hLJ
UnPlLexPVSSblZVxxuXyidtOursjNqltHOkR1jCdbnmt4bmuWO7AhqiIildMzXch
bncG7vpeRG8ZnN+A9LZbOOanCut9m8tUeHjr43ufftVKNBlLkz6HsBulbyDFTZ7Y
d7ie727uL2rGnQQq/flw8Tp7WTKzgAylV04H36bBhiKxMCZbbE0ucXgCt0yKxuCx
lN1Vm+T0D4GpqbQjIY0RxUjqEqbL77gQk2OoNRfc4HXyG8arzKFyc0lRDXBQcfyP
EIWLKDShU12hw13egeObiA8+WnpbKxKgPeg+XjNoJYJ4FjCqGWVLadzUowcA20aw
ql7j43RtSIUJbbCxdcFaORNudQDUoH4ZXahg/0bsDH9qm/WxdHz1KVtK00iqXx3m
kml7uDNXYD7ZIlz2yz6dGcy2WZuEuvLetrVztG875Admf9kRSYwpPqzD3L4CPFQW
+jnt/pFcBjt7iAE2kGRhKAEL9h3UOjGxQSEXiIbG/SLS6b+U6rbc7J2DdLxkSKqD
QD1yyJjWPPcGVgYic6VKq29a63VAsovaPCAM3Xf6UBNQ4kDbeiZeshlODnNUhi5I
FmdASwDCc72yW0NMCNa7M0YqoWRa5UkWl5tQAB6v1LGe3hhLPA5Xn73uwgZfawMO
EREH+f2WR6WZB3F1dF0G881suD1es6dZ7O4TOBajr+P1lzZ1fPIJJW70tDEaxdDJ
Gv9aCMcVYZlVv2OO1hCkcwe6z2bqB6pHdXQIS5979Ek+DQANFLWm4F13Xj+bcCCS
4TpSQmx0i65VdrJtK8mhyh8J9JSK1m8ynq/NYa+VX8n41DTxGYeSoHjK9bOhmlao
1mhnvXKr4Mr57fYib3gsC8J/eaMXDCfmnpwAme3is8wXgLHh4WyZ1jK6x/stFCpz
AVTgjfqm+2pIky9WZsPL4RPrvYOj3HPIxOxDFH7YyUe+FrhfAlWjp9ZUmnf8c7Oe
tLTMBhZLAUZTgRbvpyApQazhwp8w0ZvYFFUZJx9VYMij+nMYmdLQJOLNMVLOtgob
VkSADdbpiqpZdQ9YP/RSXad1xUbcjtmgT3KMXhjk975bCvAKDCW8pU+euP2O6wSQ
b39ArBEIsoZDXxGjupwWe5DG/FWMDgeIstzWph45z3KEAB/AAc2prhP1Qnrhcpjz
BeM82YxP4o+lkPP9qhc9VH41k4xDh1N35XWFaCu48QHJBuvI2neBTq3WUmf3OzWz
A3QL/m9kim5Q2aEM0mAxYx5shThY+aQ9wfCj+KUmKLnBcyXZLwc9g4GKoY2yhVEH
QclcsdKr3IKfvf+gZBhqNtNJnnD6pDK2MTa921hXpoe+/d7GNwoBHhFUmJc24N+D
czSf9l26sJS+rcQV5p8h2FLY6pihs9qvdLzVPGjBahWhLc3NV6x0A2p/EgNPPPsc
KeHxGOdaldYHsNVgE8y3KnXQaYkaU77gxId3JgPqjRScU9kKLMeLbOy/LCXveBkH
xR8cGabsLanEabM/ujavrq0UUS8wU6fRaA1ddhMDjxFM4oiWeibBGV1gVdx8zYXv
dbwQ+ZCVwXcEgdTZa0zSR7Uo9L3XkulTbH08EmDavocI8XUlKHRPEqaGJTigGTCy
kOXiZoC+CjobRGoX3wU0ceP3bjw3j1yqTjSVyZ+sKC/NFuV/2E39hQByF9qH1xx5
Mk/ZmRooSD6s5mfCO/mYkJREk8uFrtj6dKYzEcgnWoIu62RNAAMQafVPovbVZhFh
DFNFgv7wiNFlbYgfdR+vAPsP8De/PfnJaTmVdvZDE13Gy3CiBTx06vESRJX75158
5XYviT/KeyhgKaM5slhxSiIdeWK9Xcylqp76v8LLl5rRMQLOkZRtGgms3p+7hFNx
GX3isEo1WnSs2fD2NFS67GTU5KQdmEafEenL0XQzjuQV0U76Ttfirya3PiEFRg98
+l1TMo5CSLgM3EiEs9ukTqKi9fw4dHMeyW9fUK8g75GA/ABoed5vqIXfYnlbex4W
5SsMKYhxlXRHlV1Afk+wtUOuuE/VGvWNcLfT5Uhi8AxHP/BIxLSgCag1YgMRMcHK
yP70PbgzogIgc0WlTOp3lrYsxSpye7T+Leb2gygKcMm8qU3c7c0QxT8GuPjtumKo
cHSI66BtZ3v9XOkayzxzBxutA3DWJF+ZTsZoqeOP2MZLN1z++gSvfbrmgtMoBHF1
4jO/HhkYbJ3fDQbwiGRMwFMVPex7ij4cZvtrepIygkOWFYTP9ADGCUoPwgwXgwmv
4tQbyMxGmFyZnZRUG75j6sSjc02k7WABCpahtivFeDaLVykxf67H8rD+CB25spSg
hH307BtvUPCpgU8c9ygtlhv8AsV9qjaTpZXZOWENAUZsvhKah/fhEpC6fYlWlZvi
TVmj7myxf16xxmOCzEQq+OQ7h87DRgYIZT0Dt5j5jjk+q43zLp08GX3PC4iCTlY7
zfiX8+bbq2DE67TEceAslzjr2Lr0f2xUMxS2E9QpR3ZBQ5apogcpepc19GI2X0Oj
Fnk0/9bE6ja6rFCRhfmt88u9Pv5ArCtxIA4Z3O4UV1/nx3bz2744Wf5VLM7wuP2l
iKo1WNih8vtyw96NtHy4mmszm5FVLJicq38po6XEDjbwBWxd0l6Qq/fFKN+vqZYm
ZL+FOkj+mRIWXryd0eONTWnmcMzX62EwpaQHPYKTC64/1D7KaqlAvsUUI8Swv40z
7kMR97AdaW5YZrFauQJnV0p4zR/PkAsoznVG3Ff2mzy89ceU0YMX+t7EHwnovMlp
bG4SQdHx4yKzIpY/HZOclq0qUSewMCI3dLtRWZm9DWArWBsO+/BNmy9T9OyaBfwb
XennFRbWaprUXMJoBxo/gkAqgTdk4C3Q/tMVxyBQB60t1Fw+YwBku7yCuYc+iPfR
oiuSqcn8uu7ag3qXDHglBrIyqPebXuZp6bqSJobMh0XBxcaEFaJhujC4mJSbtShk
TF1suZi1T50gL/4izjPq7k9o3UtTfweI3leK/WcMgH6VIvpInTeAKykD5lSFqssv
zuC5zJEWDFa/Wa3iGdMjBRVZbdgf45+RoH3kkFrrIa4inC3b+pjbZul6OxA6bIfX
ocf1kX0R3jfBPq2iodz+mulmIjEeCaUnSsJPMFa+bVb/EfxGQ6UE/G2gvPNnwuFV
G7uDbWhNo5+aCJAwy1+kBex8wY7VqWm8lGmOzuTNFwh/fxXbWkWs77LpcPdeGY5Q
q4ZHMV5r2jQ3Atc2l857MlVzSPg4vxtF8LLQjXnkSf/pgRajnd+PBKfDRNCn5arG
YiyG+boJnGsOrh5/tAc0yKus6vcqXMOgE02XJmPquGcW5nK9Y8Xg6HVrzMPXADza
N8+MJLymOsfq9H2bhiju8ErXFxcRn8b8h6ZcuspXWPloQyAEVEefUgyAyLhR8Lvb
pzB/5TaAfVmTIuthQgjkqIslyAQE/GItRzxIq+nyiDWyQyB44N4Ib3errEIZw/w8
HpgZubnqrE7IBhQDE41M3c9n1S+2AlVt1sQgLKv2IPWmI/k6KiaSpDIg7rSNGguZ
x6xwPIQM0DRQCBbpdfLGHSpAl4HSbGtHFXFGtFeTTm1H7DZ3G3Lfb9xWm0kLSnny
wOrM2wKNmJspjNxVYri1bd7jRcj/lwJDk7IWgmWAns+FlejbHDcLntpTEf7bC+XY
y2lZsPp7V7GgnA0oB6159GANC9DLcnAY5GyIav99GhKDIXRYgFl8BrUz1285sUPY
rNm8MUvk8AGd3WKlVcPLBLS/OHdZDvH8di8AYWFcWIXZ6Keu9D+aBLh7fmrFbdds
fuvB7mlNFY6xPmr8QMXLsInsAuzTGg13zMxV1i+kdJDoahyYtWbzhmsHOHEuW55h
UEOOt67J5Hez9HXziKMsrHU3x0FHy3CLZLFcrf6rxdVAuvT2EX3neidUIpaDbZNC
SOhx386tNmJwp0y5j85kLtm/OCKYOCgKutxcSwkM+IZSvZ15AHpfRR0dxzyHAyDH
u8xSPwAtaGM8XP9YBPYZJy11HDePvwjy/JjP/tF17BnpioeXN0AxQQdj+DX2Q+ru
B8E62yKI5pCHTkwiRkxAszF7t8FEWBkJ47UjqSR2u/wjSHE8Run27CgE1YdZFGKq
/laDs1S54rF9wL7ve+xw2Wt5JnhoN7oL01QsDCLA/CqSv0N5LGAdtiOURFXsHw+X
v0B/+Ckqe+mrCwAFOVkpTZrUK53OztD3D5ouR3o4TPa6KELqmMMHO1L25VaxBRBl
tD79mdjxQdEGnvX0eBmFk2ou7GCdJzDcxkdTI5cPt+Bztv5gfXv1N6D6B9dIkKsV
Xp32aX6d0amk6UNsvzN8DiKCyOpBHeGaNTwvzolYdjd9cBstmZJpB9MbkETeQTnH
kEa8IYX/ImBnwZbJcnoqRup1yvMTbaeo76tbgDUzMhzsFE4M9y8Yzp3vdzQHMb+C
mrfl+IrA9Zm1iuN4G4/VZe1XCJrNCmXlEjTdVmoE8pzVNTyqgVf+QYz+/qWUiyD0
A8oXtqn626GlqV2H3pbOrKEVN04pnNmk3Q//+pYlzaP0npbnEH5RkGXCqGzDBnzh
1528DSA+VWHn4E73jPI0lR4fUumzQf7gnawyTV0B9goodxh8B4wrd5njrgGaLk20
cXKc396KSHDpl2zEob0wPGGwlTLJsqt9N38kJFdECU53efRRfxp9A8hDDaGuDuQC
zdCjLFIYSXVK8jJahmEkHJ6onAjP8qj1XQ+BiJHlsVe0jAwuH8ILG2niEme+4Wu1
Sjdz2MddHCIzVJwtluiEWdF157EP+/VgcBQBLfubA3bWDoroFhb/i+Ek0gP4lHNc
M31dm+Q9g5sd7Q+iGeGM08l92EN+ZGUTKy8n9Q+OP9OmADB0LWvLY1kBeGtY0zmE
rITFMQtpWq8ix4/R5Tj+MI4VCiGk8DlqP3kREXsrsmt11ME5eLALbmLUnL03Q2tj
LWpQzAhEXY5KoP9T5qcXa8ZMQdi6L6qtegUkgeR9/8H+cj4bXTRlJ60dxbN1K7Js
l5nLT3idj7XayJdQjcGha0l53AkWFR1NvDjOifRtWaqjSlmv+BObEe+qIfmM4qqm
pxf5t7mAeNiz1ggOSmLy2nm8JC1qzI43gvOlnggtQjTuU9pSWvYzZL2AQpVgco1S
aznwygV9Fe1/tBewjCWDFUxEgC0lJ8ZiLOl0VTz8kspS5LKfJojwopOjABD2+YVy
YIGrZAPPWvQE7/l4um9/5udMO32KwXcdN06IOugyWd/NnG4UWqzPrTPdi+lV83QU
NMd6i3u9eAilaQ+e2w6IdBt0B3cAH8J0C54jRv+StOWo2epRP6jVgPc7SBR9GuLt
7tPHF6abS24/XTuTfqxIGToIcy6bBc+btn7mPRRrSPmZOKGKUuf0vw9Lys6Itd3i
IGqn7FjxQEIFIwwopk6Tai3XdbmI5P+2b56xfUiL73U9yCs6Cv1wLxN/FPRfDyx6
ppeTF239515Al17VZ3+pRxtBfzK8c6AuakaLiN38+CwRyNBxmqySV2O2R+d8xfFj
WrJWsiAlGW4DdNaT2AIp0Nj9Wvj3Su75AoTEESRSO8KrwQr1fIQq81fqYa7EHvQi
3Ka7/WJqaopFtAPlc3TylM1vjD/VrGPeLlPzrJIohwdP9ffqF1c3t9eSu/adyweC
E8eYsd4rr7i5aDQNIba+9EX/TtCpNBhnAEgZKMgGapIUSVg9vWDuYpcIfjyU8mxq
NvzjYsBC8IYF7HxmoiVhe2BeHGK5gRx1r355U/0zkPi3IP5wL9Ju+lV0A+ITS04E
/W3HVc+8Oz8A8n5dwo+P5XYENMGKAq9yXjnvTKjobxjirwyJK7r4JbRbYnYZAYeB
FN5f+kZ7Zpp71zEHzNEMeGQsId9KUKLreQUSwvfJ3zPRipHcqKBp4hgDiPBgcVnw
znW9s4qwUuHVMJ6/Euym41NfIWBC+5mQoiqq9p9dOOnzPcnbDWSnuRqYhDfVLRTo
ke4q3IgQIaPjXucAt1qie91bQsvzVRw1AHNaiqeUPxNokSGKb6y7pxvgJyiPUL6p
DuwTZfYpnzy9o4qOEwo0NISD2vljnesKvUPe740XJRXK8scfhVbW9ouDlnLOXSpT
kOyJ3NiKcqVXhOii2vqN58zlfGcJrtsDsmwgblclUfQFug0Ya8IYzobDCmX9glc2
L7o8XgxIDPtu1b7W+wiaRb+ueX3O5qKrScWWo/YRDw1WWEoRz7nRKFfa0PUAwtlo
aM9cUkQA4JCNO+AH69/4T8lPYXdk7LdlW03FI5+JDFZlcSP4SlUYmIJsZIJ2Jw88
qaAeHWawYmIld8UpLLIIRM0OGi3UZkqGjV//KUbEFnIuZt/tUTsYxCdQ5LqV3JvM
xRrpAnP7PA++zW9j0WgPFawrJkR6sjh8Fm1Oiw4LefK+UWYfgSYxIHhwpjsilYwz
ANR1Yxc73E4YDaYVFYkDEgHXiqa9eEB0OeIQepfGMymzqb2NGM4XZ7aBjKE3RG1T
UbMrwGwb092vvoFUrzta2iCQVCsVM8L0FLW+55jieJASWfmduN2uwt9XWvx+xppB
Pl6zVJSPkV5FY1WpP4aqnbp5uIB0nOSykynAlelBAs5LLPZ3zB/OvMPq3FRjgHIj
6sQh7WSQ+Z2PFCjtmzeMWbkXgmT1TVGhTQL5HsUSXrDLA7DKI4wITpSBe0ktAuFD
06+vUWHiDMNKXQD+fOP/btrcmGTw2fKe7UfmLxD2vPmPxxX7PGGLA/1sz1bsO4he
FFItSLKyPF0Xc0nAIbGyB6ZnPlC2/hXAp5m9fCxNpmHc3yPEl/7NnLFyqh2bOuZZ
bvxZzHaZS+fEEFj1pfNziZ9YdfM2cbf9kmDO6HiuI9kSQrtUmT4MGJW6CBKkTcl0
f35ensq1X44aFWhyPnpFdhsAMMP8jyipz43mxSyFFA92OzJ52V6uxw2by0y8Ru3N
kr3YbGU9n8tDZ/Rj7b1oo32Q653isokyfrJXy/jvlP35DlDW83BDQICGSitNSsjD
t9ObiLQ9HB/fNOEzoMq9uhvDpzBfPuO0OuUehrk6G39ffpjn8jto6WBtr+KqMISF
fN4u8yYDTSoizdNzlOnPvgOjA9SKkn2lInqcC+2tSiZvOSph4fB2K9BltLAblmZo
q5dlXcFPhHxgNrke0FjxXYHTxnO8VSkwfGVOdbdCO0rTURnbf77rsW1RO07ar9IV
jRMfWcL/ZQvnCq8cRiCsV9V88H9mBV9+v4RLB6Vbs5UBB2EUf5rBiWf1UA7Q8Ti3
oVzMHDbmWBxOakZmh3pkay19dXMJggHynyycACgHCXgV0/i1bHGVuIdYdVp14EKN
e7K2gImmvcGS58sJefVmBQ6bEjdoawUI4wRjsTV6U01UmG/iWN/y/JQLI7hg0rrJ
8KQeY2oQjw24AnzyZMQnw/8rtMyWNNrk+nsfJcVi2F23QnQixLuGcPmI3JSmjsyk
6KIHeoMhtPwQxTLPUeu6FlLsNVyzt8rmULHPnRxPkpQTloeBhpZTSNDEdhq2XJw4
vLSLqWqhW9MIvm4tOFUwalPNHEMQf2oxlEaIv8VN1wd15fRiWN/ma+LTBT+eGbyy
i4QtUCVLDF7bs1sG53Rx6WRY6a4OuNfHpGimu2w/6mMlE3y7dIzudrB9SfRCCRLw
aXRIWql8eXidi54smZy1RcP805Y7tGTjRezQ8d72JmiMUNLSJZN4UDv52o9+Pln5
Gi6qDixfzFHOSB+2wPuBjsefzVGeli6MFo9p6tcI5c731O2XjiDe6TKA3x/NOPa2
a2Y/UeSWv+Oob4fxXrgU4Ho7aVylbZsGlwrkIDiuQyVkhXFkYuMSeNAHqMqMZ059
+eVnphEohoQjTWRBA4ZtzQ7HcVzOSu3YBOZTz2lu/0+U5cJOB7DIqVwgmylf+ZE1
CBiag0W4u2IQxYNNTxq809Lcj3RFdO7MiFaAz6+FEMtl1Axc5eMdcpU7PQY8ZjRH
oeBRFHo+qa77cwoa3d2TAGwNH4fsIkgZvq7IP9nt1bChO07ZuM8fvgPc90/PvV2F
LH0HkzMMpmUnSIQnrMTxxcaktu2fqaTB4LT2Xc3YkV5ST7DRGNzJtUCQRI+czRmE
v9F/Jf//mLGOoTvDSY37/PpUE2MgQQgGPRZBvZc4E7VyVIMXe14Mn++jIOquqj1m
/oxgHm+IaEwjhZWgLNYqqVlJJZjUQDV3Zya6i2MvOj2sinmCdRPOXVighab56zqL
GJ8Nir7TRq2eeyjDszUQw/Xh+AMacam3X+nDaGKn70K2RLK7IVgJF16wmVAafKT8
OR4v/0axXH79BiCFu8CzQ/CSdB/w7n78CPQzQO1mIeg9a4huWr85w6QwOwTT7VkR
9jzvfPGQpd1jkXaXlFLuI4uIYGPK6FrCnx0QFJ67kXyCxDVoYF6ihiAJAUO7yC6k
47sB1f/iYjztNHcxBqbLjDU+rUj5dxie03KKo9WCvon+eLhb32V/QFN3N5Jzd+UH
U5XuISJwgcehYHyi+m6bDz+g3FxZSPQj1GIQSlQLA+1mL+A73AvPwnenklRzbWgn
p+zrLrag2bERiauICQkF/SVh+O55jRY5L8XYQUPYYPHb426AXxG9jdKJW7DgHGsU
5q8pUn582OMoHDPYhCrr+XDseKMDImYmcM6qMfHIcB3Fk25uAdRJjXKAvnnkOgD6
78F9Fhjucdbg11bBWLwFMP2Dd5PWKVHFyAr29g4WYckLxXXfWJOvB5Zi6vyv9Y1O
z1fuzAALUglW4muub0HN+oXtR7fU1kybzbEvP0xyJbNXENfXSGRahMj5cF0MbLcW
E1apAzlFKJRr+3xFapGlPSerbqUiwopQyJS7+JSZo3+51MJxBI1g8uBvbOabsF0d
KO+LF3vruj1IYlsAPyLGFgw3KZZlcJEEqSt5+nXL5QLHObTvjivJB+VlE8D+PjjV
2KQQCWPk+4rTEpN/pjoOf18dFfO/fLNYumNNTFYwaVMNigAeryb7djioc/m2WGgH
vUL4hppX2WqYUBhk1aREkvCqWeHXth8668m9juBgqbZo59D7F9tX2ecfldCkY2fD
TWmchIK15qxtCySqax2YpY4iqq9ISIL6sLak8YUOWFz/5iHlQkC3mKjlyiCgNVuT
Wpyy4ot0UY+CARppOBwdioMUEf8byrOh/yYa+7OJjPtM6zld7SFlYTIuolcw0GxK
znrjwuUpkCd9lfGbBSlEf28T4zZLzgk9wt+VoIsGYLA/KZkpVSYlUkF2a4BHk4rD
seCPaPqQfCARfStYim8G7ASNrzavePDxsXIvtCKB/IZIbUbnVi0msCPQMsG6XqL2
vMgcijKMABlahxfTawTPlCVgBXyLj4qHdpjFMvUSUxwu3ZaxnL8CLzWCszRnel27
AenUSwmEj5mUIQ8QT/iym6lBJ+1zAO7YodSfRpOluTF/Mxla+CIeOr6VHznxgblz
GJJQkImPPFYd+PgNFKXS4TINx0mTA6mOVsGNG0uSGpZ6pMtXNf3quip8is98MB+Q
FKEBQVuOpGdQYEzxtwuVFZHpdb8HkPbCD70LCx+xQwwcbRNCOYDauWvpOKVFSdqv
WF7VYffKsa8QYg24NvMilGhXF0mahOf5RP0jrlTHKKRSKgKMZFihsFPMZsTf1mMi
TP7Khxf5VaRcaj0vw4+ikEsGZeAba4J4ByazNNim8niHuKQPkcFydTA+PUYMX4vR
G82JPPhG8RCZaDw5AZdiNr6pIt9++9Y54UYNvvB1BnDShnUTaeJ4NhNXLcvfziUl
G1LwNpgy/bnOLl+rHuhvDfM1e6fdLoqPjGLT7uqVGb1nWPPjOPRHW7p1J1y3x7NQ
Q9KytGXmkl8Z+16EO/wW/NjsTYvG7+KMXqWeO72XFtSn+AATqQKr0p85kv+nfz/L
jVVS26CQi/Bg4DmOot0tL4e+o0dt0RW5WuVebAUVDunzrmjaHEYd8wUHb600iEfG
QRyMunoO1cELE1/y+SNx1Z9MVWNGQ1c+OlkFl+f6d8GMDjA14Ul6rEyBVBfvOi/C
Lz/QZBKUTRWFN0WfW++qCcpn+lW67HHnAX4riVn3UuNRlc2GdXyuADBiEHRptlOJ
IRLnGdcf63TqoJcUETP8nk5ij4fbM1+1qn2O3msR49gEcKOFJgSEMgPc95xNiZJa
5gLmjyfgSe/vlmOW56pQJ2bdWi5Nt2D5hvE7DHvPaofOEmhFqCAwkgF+jn+h9phy
g4vaP8oK84+T6KS9wLLPOF5vp8svuA6YAOIyObbSJHS6fRbuYMUNvm8GL5d8vBMg
v8OI7mcrw/XARx/i69hdx7S/ORlc1QB5dLUFH1RZok89AhZaaxgsUpFdHVooJXNW
SzXYp7+ERZEb8YW01VXx0rUMyqbka8bL2uccKIK+jmDOQ6MbIJXpFYlHiVi0typC
Lptlf7smc+L9Okm1D2YW47yRJlK7lsSqpsH4KCVKCJpLlOMEmGk0ueqVWfP8qEu6
b0Fug5qgqcxBnvT3/FFjZ8AgQkNICcSM2h6XoYyAq3yaruX79iRb0o4vX2LyokCR
FfvQL3nSSVPPMOTa+zC8ytjiSuCbIBi1EQyr762Rwt06j/K59qh6EZbIr0q0K8rJ
TgOs2WK1troM28OpSKVrTOlYzdD/bRUpyCRGSDstFEb+nNIT3eS1IqK+r02ikf5v
1iqP29kNPHZvcJ6YsoubJ4k7Kb2eNRm+f4bsTvGiC5QxH7nojYOHmCDRFDiZszdv
4AK9w9vdwR/QUHc55pdO0s5Luc5c/DtOBKVBRtF7hbEzlItluRAAkFUxVetUnhf8
VfkRqBum9E2c1d7aLdspBpF8YLLlcdXfjUVVIWCUamKHdBPqfaOs7Flchot37H9l
JgzpHltVfbUeV5OtzPZjIFfiDioeqz5J9/h4AneEk6V6EqQwwDF889Cf+QYNHy6U
MpqQuLKHw1LoM1sn+QUYxggP8Mf62GgTMz+YsRrTA2McD1PP4vBt9G+wJ4vvlGfB
KFta89ARuLbfUAjlal7duXTKJSOUIwff092rf7emyLjIThG+Mr1GThV2D5uuq+LX
JHALH2HBubQlbyclD/8+lOrD4voa5GBHCv6aEuhQNkHziTWaB3bZLKT7KPt+VBE6
oNYiSM6+6+vN9UOmUNL7ojA3s8xTNj3edMrDdDCqPayuxXOQSQNWjELc2GFdJpHb
0ADHVqXid+Aq6PkxoJUzrCtUHmLMsVtRHnYFxKlg6H5Efp/cope+FuL6hENicn6Q
uC6PRopSwafNb+/Cs+cNFIwDHv3ZAincb0SNdssD7Fw=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ckD9jtVzdk/7qlGsx6ho57eiJrpk1dQZtGfVu4WhRH1pl5GMWcqeo+3UMOxbe0/Y
t2YoLOstOOJmYZ27NyY7mNHjsFbPSyvHSq/my1lzEQ+Z5o88ejUyns5U56C2Ap1D
+iM4LHpwCBq0D2t7vLMdB4la8gG2xQvKOOIayPuV1rvAKSf5uBvwHfCqdaXBfW7G
nGkeLF9Ll49FSJGFdA9djTqA/GbScyMmbrv/g+HaQrzX7VzXwTH88GBmj0VdsMXq
Ng8Mvsb3EzONh1bCwY/sKvlkzKTsMorVKrDt4YQBL5HBC3N8JutUYvkfOcmrxuAL
cZq1vHWaR7SOg/uvCruVXA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
liZlkVKma93Ea1ZuojeG7STBjKYvaPGxFGLI0/Q3Il1oFoImPEFqedMgnQcCSDTr
3akLSPJ9YSZQKOGN5ryN6ZVNhGONMT08ZlYpbXHY1KjmIvUETmFmm1UgtFcx71bT
gcYtxRjb6btOxPMrNtQC9DOGavvgBeFoRz2vSURHWSu2A4+Z5iHG5tuoFUzXa+oc
c1fX33JYBmIcX98IEu/lbxDl949SYu+aWPKVx4s/X8IBQnHrwVP/g1CkZg9iINaL
Lk/NnHQfC9Pdo01B10yoiru2oBpO9wWj5NK832AK4thQQpTvHSDO8/lqIM8fDRG4
rqhj/HZekFHbyXOQIkEuPnfvoioaeDl9/wVxVqKPRv588yqbdomDFWx80+JFSh6n
q+XnrJiOjCLdbFBCbVrlzaIesxtrS1k8XVTv4y56tQfjn4823ioKdB6A15CpOAHA
Fd8/kacp9UoSPKsolEzz/E8kl594jtMnY1Itp8cbk2xeNeWS9pCKjB8ezh4cvVHG
JFp3LIwmS78+TTseK6QQ2yvxBy+mFNd1x6IKbtc9NdANqBtTa8RCVtxrWHMV/X4z
3TYk3Zwu6b0J7KMs3I/SlhDmjmYgiHpNXpxodRtmuxsYGAq7YIc2f4qjBNd2qfVT
SHOplae31DG9hmy1CIjLctUKWKK+hazTEQj1gyEF15XqPMI8v90xCQZ39or9FwEH
XrN8roGiFUNQ74aVVE3gZ9UCbfWKgEbTF8xSaji1Xdbxr7T27CzOgBolWBRCY4s6
CGpCVuUlwpHwU9QQZvAWu0S96cQyvvmkWdEswqArnAQsvcPQ0tofmMXfpYCnXyg8
OoM5FJvwR8UI6A5mNn2S3upF0VRump+4n8mHmoBy1tstt2BNPNSrQ7G/4vv7qbyS
NTpe0ckdNth2/vNaQ0NwIF2oFpDbtdYmVBhPJIHFwFEO9D3pGdfG2+wL4NxzhiXp
51bb0yLn4LfWJt+tnVikpbgcjDQylqyhXL2DNLHIo3MnN6aQgLoMFK0hygzujPdB
VHoa2edMiM0GSGHh/CiX7NPWr/7Ao2qhf7v6uZdSSXeIVt0ECtHYtYWIuFQNlCkG
0gRiJSwSODb6J6WpXBhXcR4k8ZOoNmuuhl1zMnfsaZ5c0l8YL5OotDpbMXviEruU
7iwh4teZdp0yXIKof+kUBBD5lJxn2yO4YuDuOvrMH+ZEEtEvFltdMUiEDQX2QFqV
qWmX1UCeyQuj8ZRDroqhKm5Tfk1j3tBN3bv61OjVS4SFl1d5IPHgj+dwG+IoXVA8
m27/hBdocY/GFsnF6dS59X1HVIXg0ZgVyVuRYJHSsDWjV5XDEqJu9UFnZzEFT0uX
3zRxDtzdU3XosoNAes/YQ87USBLOjQMUGRCM0uV4AdR2nvjuhV+zC3igW8sWq6mK
Zp/R2vbmXXX0Of51xe7G0VRT4wtlfWZeETk/1DRu1MuFl1Ei7TMSy06rP1qdy+CL
YJrK/YXKcIAngER6Er7iKaBjX8ODwIQ5Cl1CAWlS2ojGZZOnCs1qRqsfFGJCq+Da
ajxrs6mgh8M2sI4uYOAQ1wqW14BVzUU4MDzuviZMuLFtCsFwOqY+HA3ZanmW1NNN
nG87LtIg6XqqRMSTEn/rHTySq2E5jdYHMLjSPmnb1DI9+dj6MnCKWh+/zm1tKn3w
OPNIPiCpaKVYO0Aqvk6TLGs1NpXNXVKWUoOC9o7zhXNMhZVYFtFiQ/0FU3zCxHsg
HAHkD+xd5RYiTi0IcBz9fU6XXe7ck3+72YYygYDkU4qTXgAInrfSPRBJCEHlGdac
uTNn5jW89LA6Y5HsZZahWpTCE7hfNm1gnZeEzLhzxw0BH3NG0vmgkXoneC0XzBA7
quZf5mVCXbz9F7vYBjQFhlONGYQoFDSHFROT7X3DUN8+R9FipBNtpFcRas5oFJoe
sMyLRvZt607PvmStmIwYZQtnTerXpU+wli1buRjbkN0EZloDDx03OXg/PCSbHHke
88Q91ZaI0eEERCBgm10ZBbfzXPYDDrkjQSoPfHSNwpm6i1HQlkxhQe+rnx/TjKdi
g1Bc5BGEUaxlty26G5/nxhqIyE/x4vvFjTrzOYHBgK1Tli+bdsOAtyN0AAQ0ZX+H
TJkf1/aofKtwo+pYDUTsj1ADWJGtNFjOuRN68POgdC1Y/XCrRj+7sKb3aj2p0kpb
cHvcu/PCsXMx2EtuljfRQXSR1Cvy4nB4a4psAFhTv2rsDwgt1l+XgTTs4WciDomi
/UpRQbvrMZoO0eFVkyEN6zRohhk23DkGakIKCcy5yOMQ2XZaiyIeFfC75ETSnYZ3
eQ6vpmhPIotXewXLRp7LWOeAUYR3sTymkHuGQmFmsTAcz2isJ/QpzIEhHsXq99yj
EoMxgZeyxUXPTXYDi2hmouSe+aViSwDrmAlVMqiy1z/2P7XLgozHRKlCHM/acFHT
lLvB+LwS1P3ow/Ul42lhUcW3cyaLUJFjNcDaMNOcpJdakMz6SJDYoZzksosJeZTm
JCWqCk9rI3x6CyGF9AWFvMc+S2e188AofOsS9zhC2UQzQs711oAp39mXlVUrPD7V
Q9nh9SqE7K23+I68OecczHfwVw7QwfTbxNdTamIlmA6HyezLuqXHLaLVbjILel5J
PK9fb2TW33jSkRkj/eMzRH/bz9LFtMyvQRsyurd3+GNfxcU0bDWrgJ/d0lV8uUTr
syKKNF4X9KujHf9J9A8GnwFQnY9qx+lToz4NhkvH941gr2DJMzCY21BdLvIJQNbW
Xu9i6g+lBm6dq5gTZUZLtNkEThuSo6P0xl9RPDnLIyJYuitApoYJcAF1McbEEZDv
KZvTA2cntYQ1mojqR6GuBotA1HLpPGeXQXk1bikuD6YGGcvhuOCxLxTOCIS2A7zQ
Fu54uGM4hDbBSv3OoGr2bQs4EvVe9XBa6lRDdN77kKRjiji+pOAkBZLPpCK88E9i
47m2Z/i7tUe6bkqIsNpbaPl2TisKIQG9AF8w7M43iqsO11mu8B97ziUm6UlC0tGr
F3TCnOd209MJu4r6sj3u8AIO8vU6uz3Ivrojvyod9TxaDweXG+XrWiF2+diaQr+N
br7r0K5UD9uKKxTPE1cXLdOg0I6bvxcSiUwhvU7JAfDIiLbrupr4qcKAEJg/clR8
bSQxVZK19QT8NGm6j4i4u2YOHLndRMWz3vAjd4sFyM5XAd053VDdhG9InxccGHtw
gACj/B1nYxEtnVnnISgynDl80IDy7kJ/4AzcXJMgKZZk4HihkkzAj1oke/hxmV0a
mDlN2SCpVz9v5Ig7Cx7zNa4Aw2zSktcUepbGD1y6a83XwlKXjI0gMjm6ehYbMLJQ
vgysUN3/upsCbRebnGi7yBthFeotMEtrNNrE9pia9UbC1IiuuKV0mClLtg9Ajg44
/+BemJQAeGi26wnvcoNPn7+Whxa4+kR8XQ5QUlYPFik5Tx8urT6jKdwKjm/zroTl
jJoPxZo535VtO/hkM9yRBzKYDeOnUSSPtc3L+9nCdGPIS2yZ34j0bMIpBinR37gu
xw6DLdkRlisKcHiJecG8MhN6epa9ZHKvcB5OXIZ993HS8bVlHjTkcqCj6/eBUSoV
S/elwY/XGMRosQB9nVRaGdfm+q+02VncDG5llqAR6aFPB1ixLdBjO7t1kvNoHyWj
YjDk/oFXeudp2MEdobS6+SFW6CI8JXmr5xQOyFqHqbqBSMNrnEgQdftIRU+pRaYI
7vm/6T30wAanFgK1sbCbggOW3Bfy08Ot28ZaaqCyeFpBe/HD3kLdcXUQtGTlp6Ht
PAvjq542MeiWGEtKCN1EYPCXnaPanAvNE9fovkJADSBPX5UPSYNENuI/Q+795V7v
9L/J7WgVCjFp1peIQ5GTxVqS1vvxc9kUo8DzH5Ea78R1qxDU75xYQWGu8WehJpT7
PpXEt+L3qwYDu9F8evdaZhJQ2Ad06Hy2S4vmEdRtqgcoCOSGeOTsuc31uYtePRs8
0pg56y/4D4Ou4LUMSCZYSK9XtEtgwczyJu45P92kWiebsD87T3mGBXuVn4TJTrK5
V21ZBLbdD2XvzMgEigNsrafXUKiX9rH5mC1bTj0xKp68Z/6h2YcjqxqDlRGPCtZk
Xo6re3JXG8VTdzR/0jQOyTPOvFfqryU/fuLYlu0cYJOC9GyOoSCmfBueDxjc0wt4
H9UixZ7RrPdnjIK/BI22T/ESYpEbgiym2PB+BciaFvXq2He/y5hRbYeYG8nWBIVp
oywk6s0IzeYLzgMgzOJaYiVuXHyWKCmuG0aqImQb6JF0MksFMwkYgnxT6BfKnh63
Y/BUwL8qObzo6TIRTFYdToD2lDWE5mZNipdKY/qPPnkFQc4cAWKcTH3wk/W8zzzz
A7r1g4otfWdUCKA0snqEMx9OzpqLAR1XsrM0vyyEE1s5h31drg1lnyDDSSkNDxvl
LVauEExA0s9c7deQGHID/8RUu4aao1xt1xo86ls5NYF5x16yIcHkKKNfTuWcpJJH
VNPKvzGoFP/+surekqn1/bIqVOTq0goGBgrEJiQS2XPcIsSlY28ryMnhCtzX1fks
OtccuUTvY7bixDfySwQ2c0q+Dg2Jc82tR0QDegkfUkh+6YWSMTKta7DBa/2Sd85m
EVmlqmsoJcjt2UlyAhmI5HTjlmfjGhBDAXgKnainMMGE4z7EWbtzqQZFjds4zj9y
BFVvmgps5nKqMOYH5tv9x9CZjqhPXhgw1N+8AZ2PJdoiA9tl2SH9CMNWbRlhRECI
K21ydr1wsljuWiIjym9OqG/7oFg3445HKSTZdQGvTTZxWfOHWQTd18T00epgbX9+
rjRxIN9FnqRQpyeK0RwrpzGJqX4ObW1ONF2qxUTnWh9kEFkHjJ87sfoiXKnniNQ7
oUMS9gJ4z6Vk6l+UpliQC9Y2g+MakGX2megQ4s319tp2ODmzJ3urqGgUDPHeY1F/
0hNu/b5/mfKGpgC5DtcRE6A6hZw0DTiaCu3rZuZbGVbHy0YTcJDOJ0lNjgZmTST3
C3C/lhjNAB9ADbzz8bPeoQO4L1V1LKxu6vVviDT/b5g5BtykvnJxfoM+BmpaONtU
quqUyx0M6OiPBjbNmf7ziiVFWO66OJQVkKChSz+TFQIWQXFwL0tsSt5QjFltkWxI
7TNWxMN/VaTYDpzw8HuAT28S+MrKl2wGa+bA+6MZBBqroJLb45qPP4JX0GvvRgVy
q8qnqPHz4uoRzi/cTR2gE+YJu3j+ZzOnZbLqFUe+bvz2nu+4a2PfRhdm/dvXaXzE
Ck1p625wiaTXBPoLHbMQ6yYxiCHlI+zxmXEx5b9LcnDDtM97e8UPR3q6YbJ91KSM
1w0y1QQnsR3klmVTB6Tt/5wAWRq9aoRU0j1fxQKK1mO0uOJ84gAUEmN9bePmc3sT
7Jw9HwVK934uTOtXH1LXRJnvnysdrJ0Jy4dcyyiNyiBa2VKudEjCZnlcYSsRsHdL
Tnl2fj1mcT6IJFZhVrN9TCXUSYNUft8+qPPyfz20JputNsjcXLubYfTvTIiPznYJ
un1g1orGvKKIewJIpdUHxMoxGtSAsg5oTA6a57I0oDgVt75Y1tLLIXyBf7UTnxCx
fTJGRB5JXfXexWw/t95ugrjEX7IXpm9wmW1N4UGCuuuQJcuQM6jnd6+L2hzMpITu
071+7LgmshZpKM4wu7ij2woYtd/KlGY0Of+ABvnm4v3r3a9N7WtdTmXaeRs0k7XH
dg4jK2MS/bw2nabUmncm56YhPMLu9BspWS8SduEwMkz22tMR3RDPxdeoflV891lJ
qRVUfDneYluWrwhbL+HQNs9eL9000izU4zTRTym2p4qzjIOdU5F8QihFw3ykf89U
ZoJrerRWgDpaH4E6DbTtVI2NXJdK/3ltR8ctek4cYlYWKSuhCEYjd6XvAx5UAl/H
c4hu0nEqtKoSjQ7ls8R4qmpsicVIkLzX0EJOpc1lLz9Rcady6TMETKdcc5QRXOD9
9Zl4fqx1FLGuNfaecHRYj6yRnneUC4nxZ9EujGrtFKrNN6vHxbyh8RpSkrkutFY2
65BtG7jG1YCVPopi3LWHD5njsjNRzmRUEqAUFpvrBwDbnnpYmv7uQeK9Ky6i2I2z
c6V+4saEnbi5L11Fz6w8QJfRIK9XppsaRaqSdpaXMdOInZFriuNNGtpYPhWGY61N
hKUdf8FwST9cL7GWMKwifyIrM4FPq6jNub2k0kyoj+AyrFc11+oB/pblkWKuOAUA
Zo/TiQHtMCxb+U6D8TS0MKXjYV6EofFX/vhgPZquMQIzORrP6MlGgRhSEKq0VdSv
1dSLhGfwVKN5DZ/BNGKl0XLtRSW2pI8lSOmLGBhTRltGtSqCgYUIpe03XDW4VBZS
blVtydUdcvVq1G2wCQ84MXqyjM4fXgnfroT8kexNenf3CN+SDBbsXV8qps7UgWiE
h1ONrtzCuQFIwCdfuJ6JAik2NEtd7oJAYxqDMSaU4t1RoHXwNIi6/6n9ID0ROaTs
55/TZCBL6S/UCwqRpHuVhmZ/2GDL8FJJ7Tzqos+CYUFwZ9ExrJdKsdeOalmPW9v0
nbi2d8QOkH/KvAA+5yZa6WIOJ6bbIqMcaoNp3MLsZIa7vVmFS+vGoj91Hf5LNvsg
U5euCgowZte2WxNjHRP+Bi3/s5wy0nOL7FkfHJSa4/bu5MTaMCgpIYpwSYTHJOHb
BDldLn9CS6T5F7z4qT5A0ylWHx+u7oG/BvcnFzK4EB32CuqJB6WP96hDlzoVvO9y
NdLFTU00ytcKI8SF0nTpm/7Az8ymifxg9fwdwirUuiPiueRjxvsGYq798zjBQgnc
EagQBLQPqAXdUCdc/f6vTXM3ZF26532V/KihvZ/P5Wgcs0WdmQJZ9Nc2sCCM1j9r
4jm+SeQyjwX6TkAHPv/MJP4FmK+KzS8GXpJ68MSTcrS57fzsAuXhizhT/qKMOK1Z
kcmJMql5NvidsALU7ndnxgzLyz4RPzZa8FLQmH5znD/GHUReOaFVmSTQHsMx2YWm
dnFIlk/WsZ7HqQ8BWx6Bd0/zqaCpXQ39z6cPBNfD0BYbIamczS/8iPHGHffCO0F5
TqRWjAXTG6x2Ibjuxri6BYgS1Omj9iQuG2ozXEvdFgRsOZ/r0DO/LESk+0wUqX5X
lYZ0wXWRw8SheY2VWzG6YKDCackoTcdAC8U0K+YUumwNDPBSswsBqMZ6PgNB34q2
LzDwhaKcNqtHRAIXXX3kSkuvZR7UlysfHyYz9kBg49/kkrOvXPrcDVfb2fjAP6Oo
vputM0nf6ilOlOJLl3CEPIk5wYSejHFFNWlXC7xtmM5w/ghxmpdbS6037953s6X5
Q0DjTcCTXLUruQH5ootQZGX010kFnv4hq8c08RvmYoMzOsE3WwbboiftLXdgPqlK
xHhPtF9zBEqpId5EadMnoH0T0PaR09FUNYgGL2TB/C1ZHnoMRbICo+Y9IVWhIOJ/
i7BVJGjMZfc3UOcmDi/dDIuprWqZb51vRHXkgcjee8hlkGy1WEzT952q4eq1Zd+3
mqwWuK1kc8sH7aCYY9ZnMXvLVi3/QGeVFd5YsFBZS5jjtWsud9fex9ay4epCuV16
5ni3LroSl8FBm3BijbVsjdgaic9Dvq4o3HxYX2hnNFC2gsonrEWu2AdbJlA7fQ/q
/kRXa/hYq2Mxcssm4eFpWuhCg7dIXI1wz/znHc9UkfUh6N/xHVky/SDbiqlFxD+l
3Ay0M15QL9ZDtJn7HXtBmWT1JbMNH9Y3AT2oSnYtCmEuQwT5VfoqZrxyomEmqC+j
t+br6RnoJVaxhABo832ytzN0nco1nn9zqe0NXfSYDiq0NNfHs41cTt2hZIK2g6pM
BxAHcKKXLp/V9vi7fOftRIQWDrsIpBDNwkhHRXhalY3ytDOaklXCxe6XABFF4yQv
ZNEsHgRkMgXUlhj78RtZ60cArKZUMJhpu0nSzgq5kBm8o5tCYrgX65EWimP4o9VU
VVWHqZNnenQwiCpsWTV9GZIj5+0+QJM3Lt6doOzA8I+0el1/UwVRZzax+iZir4NK
UVyTD+BNlj/mjM5w5F64RzV2IwKFuJkDHJFJ3WRk8qf0zJO6vhCGYF39/xImC6ON
NsuhgKt8Z90iil0ePE/D11bRn40RSB0zw+lUiBdEXoHo5bEL8lClIOpXN4Fbwlb1
UYMntdadv83F0vnEGlubZUOQINDocLpWzi1499mWmg7pPtaFu/i3EZefBdyvImIb
9rCwdtHl2khSmzrVZBfgQr5Af7h+E5b4FlL7U6KvCWPufkf+2V7dpxxHEQ1R++7Z
fsehXTtOD5+d7g5pQSR0C+FYeKhwE0AyXRUo/XbFdE+jg1Sj7kKGnTs0cOLpxfRU
beE8qQPjsC6PXKCQ4ja6kSLeLhPmSx7ie+629FBLrzNwum9t+H6DHJICpzY1RzWf
IjolRiZPqoMZSnD1FLlAOHhRBklrBfXxkjtbjBeE2rdXRr7JCkFnaSop2534pvGm
8tSm7N1GduiJCpbHk1Gi4BwIUm0isM4TgIkxDPJLDlvk4tisEUQSFl6SdySDq36+
iNr3/u9aObsVElWQGg31ZK3//U/lkfbH2AY2TE0qcD3RMCVaBqG0x3KOho6tXKub
mFc7vMBC3zqcOWllbWDhFkhrbRKpB1VNVs8XwQbo0vecllUj27bmDGOdIMVCwgVC
LbI9PfYetQdv0/A+hQ3prGWsaIUYmpwSREqdtRRRTWvJvyV5K7OB2Z5/26MCl8jz
0kb2o6FTVwqDoEQ/BRh/RXhVjyoPT9sQJYq/P7JXGjsUaQ3QcREiPJ3vy4S0vs8v
m7YO5H2lz98zLPigByPPlrqqTrMzL60pS75sTCCbuNSa9WE4p5RFT2eSVIHW/Elf
e/6Nh1+QwJzIGA2a1dDBaYAXKHi+VI/5rc08hAkD8U14mXLWXOAcos50vN/Zu6c3
7oNvcw/6ToN1W/iNU+IKSj13yN54y0g8eHlPCEOgL1R0+t9Qtbwv2CLq7ySOhWJ6
S7wAGp+KCepypuab2P7iay0WeTCrLc+5EX4zHl/wbuEO8B9XKRIKWlmQLLiaUoKx
lIMYcQbbW9vZwvuMvBI35qrE9mj2/DWEtXeWH1OH4Yh5DGB44CUWToBKBKUaRA6k
VS2Qy2D9zZpZVp5tuNt0KGkSWLgpBwaTOeoHVv1f3tTCOV0BNdthbt/MCywIQ6t/
x2SN6rJcFeo6Dnm9MMlEP67PFWv4Su7/gWdTdAtVph3ihtXgWyWHXDscXvuHbG64
HND/DE2DacwrXb4NJt0GfNujeC3ssdCqM4xJCgHuvkaYfJblf4Tr/7DF+Rk/rZpo
tH79PALSOyDuVZx09m0DvNT1tKrn7Sgg8LqBPhSYaKU4kvyrbZY+TqxB2vzajrxY
lUsT1FAWrZVhBUd5w20oaD96Bc4EBHhaldVws/SusMV/FtjE7FOpM7Xh8+b0jfgM
CMMsM0C4oP4iZ5fjoYQJFar14R0KK4/xGxtqlnNpxk9nFVUuvHlxIvKsKH2jaZ2p
fALord+YIWMlTNqftd+LcAkrbkvh+u5ulx+xNguKCHzHqZMpb/LHjcv3KlvMFCmo
IImPluYc0ppeQow9lR+gOEVGMt4uUCHE5t6Ac/oej9y5bhJgKbrZ24FHcKiu7hrA
lZqkPVrINoi5vXXNZCQj+s0mwEpVgDPIwU9O2zOlxOqkT+XZmABsPvpfHoWJDgc0
sImN0VOdA8Kc+GAy1A89EVPxMVW5XiRc2EEQB2c80WTAMPxKK3Ya7o2l22WpJQwc
9Jxro2quD6Ns1iqXgfxOqlHuo8geTcXT2NzHswLIcw0XFWKe6lCcKmY1TpduWnnI
6zI2WhQ4pnmM3kHwDHzUS/uDCm+AoMeZYwsu4MK/b+dV6iqgqoJVLw8Jh2RIvQMr
ih408/Sd2C/TyxV0XFti34zqP+wD7aREcdYhoXe8rp2BJIOyf5WudfwthxXi3TCk
v52p42ChBgxL0WLE3L9yVKk+1Hg9qX/svaVMZGL7pzQXtR1yttJ2vVHn27m02hOg
57m6IrB82ftSlMvjDP7A4m7QHCjt8AWHICq8geQQToBsJQ3h6amrojn8LobAbgfI
xqc9SPl8aw2+0S36pVIViBUqSHUnFdz8F4JENl06BZmeDlQuRSOPe8pAWkMXrZhR
p11b/rWSJC5nBn1dJ2JhZhmbcMcq1hopWhuJXjIr0obu2kCDIX/pl4LPcgXzYY6N
GDIbWWUz9KRVPIt7poh3HT+OFQHidj87GyJJxVooyzyONrj9MZ/Cy+QJjqwq5ULe
6z2SV8EXvGOYqEkkTDsLoxDKs4EIfxmKXxYv+7jQgcFXbE5HAFQDVSt551zbn654
pNp5T8UNLDtxN/BjvZrxdJ5mZ86rSsQ1HO8CbXIv1uUrFcI+b393VNTlFL6PNiDd
eYo6wFDhFEtjBqY3Bi1dxVYuDbFE2G1xoKZJ9Qz8rv2RI3uXHoG7XN7i196aavzW
aO2D00dLnnMVjwvrybCrr9nqpxh0lwfRm5+BFGMkIA0GZal5IP3NU/ucipwNoZJ2
QJs8HmKbmNa61rb7h7jEQs+FUmcHC3ROtSh67Ck2sAHjarMRmANbOjiysA5+FON3
EmcOqivcCAkGEtBvNoO6ayRTkgwj6Vr6brxM3yA7ZaaGfNW2frXZ8PnNkxvxvF/V
n/IK23R1dfng2/fc2zESVIUyINTVubW1UeWERc3d2/qAmmoj/IRbxKOlTTCOF/EN
kLqpwPRv98i33Y+MPbWF/CVQ3OntQ7T4vadShK5OOEnB/QrDQgoww5QZNYVN0UZQ
tRfsP5GVHkOGv3R5NpwGJr+RhTZ8/JeHajvjkH20UNHogC+OaXJwz0+ctsX8YEWk
Lboi4Vxx/ISKR0Cpf9LV1PRD7FFC/BaesOFXhKgUzK6ay6A7t7CBXoWCXYIvBuPC
F717NxsO9cTbgRvEAMt90zFfw6dgGLZScO+rsy5aw9klZFFoHmRkyNvdILh/hSH6
QzeHWbu5c2vfwQJlM792O54bA9bcXdwsnZmp06EKkm1emosewfSZEJ5+/yp506IY
QpkOivah/nwB5zBCIwuZcmwXq8P+OU8YXRaYoFtC+/vDbqtR0nncalaYgxkOV/Lw
QBEismY08VeO9smVjRqvIO5oRMjQMYNiUIoc6PboHdmBsOTSCCln//JQuwWdwPeA
a1AFrLiB98pRhSoxRyatfA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
W2aEH6uAiJOPFir/V4eL05r9hJ51145V8R3ZCH5aMFh2RZD12nJEwZvh5PwHoMfs
x4wCiUJkx9W9kL+2jEWN502qKxIUv3kM9lEdBy/j6pxMuPpxiRxlIJT3tJWEGXz0
Kcf4AWe3QOQq+RgKjSFwtpmw4nZZNHYUNdSP7cbGCPUGqp+KBbG8XyEcMp1hL8Wo
9hjAal3D18Hf5erZYZcazML8rB+N+Hzbwtftt9b5vNGc9xJRYSMBI21Xc/yrqFu1
D8jrsdt4ByTYz0AyJ7wPnR9C2XfJjiTyh9arF0Xo9iquL9OzJz3hAc7UItL1rwzr
/KvzVjVmtUUepLuYqDB7jA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11952 )
`pragma protect data_block
kLRu3e4188Nqk5VqxtpBfygmJ+KOkw2wC5jtS7/9tDuUlMp4n2NZfuA7FwGNP06u
NJC44+Y/trI725d+IR+QVBCAbj1xFc37QKEOEwKz8QIw6lIvr5WMi/TWxbr/28L8
MvNBe/pQ3y19eMHa4EjdgoFTt6Rr4anPXMcS89csPXxA4OX/1Ok/9Cf5p6LSqmrS
KqIkgYXTGySR32epOXTLQ//zBVQrLkRuVb+crA3ax3NcU2FD2mk1gd07OXaeufpI
ESzgsaBlh4QyGImCGtSDHFWxAS3cWauCt3S0z/1l1sR15JXLBitNkObto6cadhDu
bSVwaKKshxb0O2iaEXxsNUQLRmpMK0wRohFhYi2xkMJJM0uFL88SdudSCK2PWGu8
ZH2Toc/79w4Xo3CnjxpeojiS/PbxuhlfuA5ihxAYdyen5dGI7PV7vx8k+YPWGrDw
SNjAmsRc809nc/qDO2jUBB8hYgywBOmmilTHJjpZrF9zi6mehJrCSWNOGsHztFVy
EGa9ixDZz5UsyRG5BBFKZRwpKf+X4e0kjDlUYkJ+TYCgcSJYarMXrhnBiV1svoj4
HCPpP02NX2eCcDj6tzsuCtsk/FUw5wySaIS/2h+DByl5akHRV8eA2ZCQBvI0JutE
KCqQ39wRho4gSY7K1vDCGrb5Vm0VgZzPa4vQPmVQzXXJTXMtgdWdMNLsoTRAD3cG
2+7UH7t2LYgiKIdQyzaiwVcO77PBMcosD85U6mLu1qrFmMbTkBsvOTnHzAhx5BiY
xAUgc1I4170I27TcWjXmlExToJjH5+6CbcInPP+mLMkA16S13k1fvslgbhahkD3t
tio4bT03y1jOpYg+9O2cwF0ZhCtST3/p9dl12y/QZbtk4RJs3oNiBhdesy1Hazx0
fBMpnDUEbLNcRX1U/6TdDKW/Q7ftx2jKxgbrADCahJr2y6xUWUOH4UyptHGIh7Pk
+vqCRaiyuoMZ4fpBdt+bbpCctRGam8WEc45In3OpwcUGgZd3WuSOOEflR6cnuz1m
yFw6buuxjqibNCNV4PFgaPz0wovX9t15JcpkLHVzVJiDFYmVxLoZJhMUVS4uuCkY
IEhLqDamiF2+Y9up8DvHTFM0GoJ/lGEAesYuakqfUklMoi9g5atKIllFOnvP11t+
l+3UxxS5eK9BFQWjYIxQmN/pbIFjXDgev1/ZWeZ29Z8CZhgnsrVv3TltVYcvo1ED
2A1/27X8eko/0nNGkeBmSenVh8wWes+yFuVi7EIhQRgE3OzanrP3j6CqmDdQDaxU
GhpE6tZOtXgeHbKdcUJBSVTGQ3uzDo/Cq414ExS19lEXBBWPurm4n+pkH9VgYE01
ootYgBKpeg+vhs4vYnBsY7gKoPjARt6H96J8re5vwm41gOPkhF2TdymfrHqOxVg0
hj9nc4HBgBew7i+vDqfqyuaVli7qxxpWUAFsiVFhxka2pxv7Tt+CJSniJ48gJUHH
blXF+SREwQHuqYi7h5rmU/lPfVIXyhQtIdh83apVdsltjMJejl7jWyVXHHTEjXKh
ugKGa+CNddF5/rGzKfW0FLF98zYD4IezesLZxt1XgHfxhr28xX26qj4NM6SoKzD1
pjP+Yf8gHlyxZFBaqRB48dczrdizMNE0MD8XJ3yZeJ19886UJz7FLFyM5e3g/7CB
JMGOqQ9fgpGCdfwyTfI9PTLydCET4ZkapSLVpJ8yz6U3ETiFQKMBbNH+1h08NMLu
fYxMlD5MdFPAvVagiHSEbQ58hAsKRoFkH9atC4QwyscC8f95w5sMvIpLS/ZAf1MC
46nXl38rMgyfhG5MKAQXsMbBhmvKtkMzZsRYOuZhRlwEiL9c6vJS4/4iPrZS3PTn
sjjjYvsBvYD9GMkdwJtjGETNy0LHg8n/b9TDArNYsD1FTqW+sWZ5e04Xq/PD4Wli
BEmUy6Ie9QOJ/tSD1ZLTb1CZ7H2m2E6WOa0cmswBDj948fk/xhixIQH4HM6MiKgA
IFPIpathPfbGFRBNa9LhawSaMKFGRzykfiCEY/47OTskJ7rEeacd6m+MVgMDYMR6
sVpKEdCsgjsBHgXCkGEd8R19csccQJVBo5oyGALZzh8OYA7eMvtBvrrUoUWvqXD3
mdZDbPS5unPmtdXhZKRaFc5UvZSYe9By2UkygBfWEuJanAlzi0wk1hZyb6ni/0W4
Uhecb0ZmDijKRDtZOO9svCciDNLY99avehlaWAYVTNjs9P585eVqX0VnDAJFtSW0
fQ4Tr16HBTXc809+Dl0oZgeSMCND3g/vlF4Xh9VuU3lc+5jhPXEhVLN8eOrMtTiG
yARl+FSJ2WdHL98Xxa/VgngfqPxKYOtxVLv8MVJLQ79qPvtc5qNVIjmRzG+OmfuT
6nuVHQviOGACQVLhIPmveLYCh/h2omGI4eQuUbOCsZXq3ekq/wL+KTWJPGLBaGt0
t9QTxXDu0ENVzxCrgIcnHzq9OxVsxWI4rogSLwlrqc1tfhM/8GfLbduBfZGgB83I
kDJa0Hcn0ZXG9YT45NYcKH124SgMbZNVNNV11Uc0DkSt3ZLnLwmMUFNIUKOMPyY6
WxTcO7a67OPn9qR+/9qrLX/3U+bAxnpjN/fIztIqWaUi1tze9odO1gplzB0CnPiG
nSrg1VLcgmKD5Nx2Aau3QR91doKZpU3JOGjkhJQwCknv8km8W8+XHHzewCgNQCBu
WJF7VWxkHUiXOu91+C4S0sTlIWNOs+YqgyJ92TX/AfkW+Buer7auc/Z3LaYVlc1B
ridTJoUb5P2ZjLEgKBM8548H6XAKvLyomvXmVjPsH73k2CBfDJdzZ1PlORr1Lroa
GG2bMI5Qs2qqJe3OmFNNTtF532FQmNeZPaKVMqCWZ/+jsHxmiJ2XvjDjJEXshSwb
7zFEpbNEIICrjmvJ7MHhiCeUMJJM1gIN1NHG4/oSx/SPw+MyPM2Uld7TMZsrFYTA
YzsVXAQOZUZuO3+Nqx6rcvdxe7TjioXK0JcSeb5owWq7hzvaYylAvcZdHB3rLaxJ
/ZjhrJvxYFRgKhVPdWGH6uyjtyje/Njeee28EZAE7md2Ru9hNVEKrE72kip4hO21
ZT6akkHjySKTyHil2A1+PvH1tRXY52k8QmXYE47WFIHSOS6M3WB+mIIXDszZEfNn
c6e2H1tqCFbRn6K53k9W5g/0SrNMWpSdJNS237Ll/dAAG9cnuMsLA4g5FP1Ik1/r
gYQSgewrHLmAUssTDjPyvVyXH45bfW5D/ijou8EJtTYuM6es2yC27RTijIq6/dee
vZHMIuSM2GbWrPCUHDdg8cixL8TD+cKSEGFMTg9+2gAJn/zA+fuw82hOGbayAOGB
7C15kpQFm8amfgWKPUYYF7Q01GOOesZ9ZGTbnZoDdI/UllnQPDHGmdzvDKJ9OKzk
6yJ7O5QuBKxsN3ifBXp+BZLmobVdIgDKLSD8OuJS+A6GyzFAYlBLEu2ZvQUAIFdw
B9n9a+dx70EJc0RP7OGaJBzxdQyO5od3aW8FmEA/Amgxb1IlKpd2nVrSJMicYEJB
8Gpu74QbQwNxHKSD7ULok78WnmZLFbDfvFKAM/srR9Z7o09hepouDokPtJRXpkIJ
q2HXAGW65hLi0KXCdtEkDc8jJm8KnUnc3B8hbdcVKNDgqrt/QO5EvMe+x3biuduy
bktpUOOdETqVCN2kzbLutGHCCCJb1OyRG9chOHUQTMrPzSaLgto+aBxPUARqUesB
JHJ7Maoeuuc7RWAVoG7bbeyGBpzzsUvSSn2cLShAZj/L8EiSyWwl/Fzch804l7E6
8v/o56Kzy6mZzxjHaAf4CQJXgZszQDc6ovIFEO23Eoakdw37Imh8hIvD9Qy2u+pJ
WYNtivt+CcO6lmkpZhf0ddB3jnLU91PkesoC46O6GyQkJCI+Uv8u18ZLVF/CJnIG
JyIpVh3PxGit90PbQWb8gxP8Z0NJy2gx7HWrFhnW/cRXCr5WXqnJmt/XP6NxpRyA
fYLPfzJvOT8JtT53MJ4hC6xx0DKmSCMw7X8K4q//fOKo4955odi6Bv1gKNLrJ8EE
sXjCNE4gPd7T/MtWzh1TTo7uPZ+XrB8Ikv0hKpvoXRXAVQWcwnMbeHXhmy/m9rha
o0VzoDbSYTLg/XGIg6x5gLojj60OHZBMz5exi/FyuySIhC8FV5kPCouhwe9a1tAY
n/7q78GhEnxcB76ytRAWpXnSi7AzTWxJ/rOI8VtlMJo3nft6sCWROvOfa5GdX2nj
VZDHiDQX1NxdTf/7qTUX4u2RqHCvwRyzrlGB2zs1nrFwli9kO5Gb25LuHtOiUhuQ
4Cv0vgnD59vWvv2n1kXUQ3O/YoM8msOXMF4YshBWaNSSAUTXAs/j7w4L4TR9c5lh
O9mzgt3w+uM+jesiUX0mPMwTHG4wb8aIFZvCiFAbCBMdQq6wsW1+DVP+9cxRMGvl
dna0TFgDphuP10JFx7Xg92QGjI3KEOQ3h28gPputNO9iHb6P6H4AeozkLtPh0YNg
kJzeQYK2tHINpE1Zq1jqIqvABGQueDyWsXUjmMjx6VvWuthiQvc84/kx528d2uoK
Imn7EpD6iOkRP7YsO7jEkwH8NbfXXkhKroHZIsNIlkbARiCBRoFhuwf/tjx3Umqu
c2dACUspJJ7kpKlRQYDu3RhtrUFjpJfFIn+ZX2AE62EgFFVx6m3dXr+W0yBRFAgM
qCLJkSdW6t74FZWtL/FQbpWx6R1sZKYZmz3nOlh1YRBn3VKEIO+mz6lKEW5NEyI9
yqaVA7xZl8uegCrVl51PbLpcV1fK7WQ2ic8Iflic4nq0rIJgKK/Iq1T/KzMmWWQ/
3s70em8CmgXCMyr6aY5AOOe1U0F1nGbMEixxsI9zQ53v8foqthQMU4vIzORGvKQB
UG8kINz2KL2WYDHzrGFKOS6KUIOU1H/9OAaOhgtz/qP0VDwxROkWivoPWMXHVQjm
tM9I2JZDCOXf9v40z5qlOTmJjf7MlpF1xWSonYfuTzK2uzy6EZW1jLiYgzb1qhUg
a2yMCyuRsUhcFDfKuXd6lS4P8nVtqaGWIYK+L++VjxE7o6vW8sY6coJsVPkcpPcQ
SFh1qm4NLYDfGFr+/VO6lCjvSvmxlsfHqXGhKkHTweiINOElgxnKIi9KMIcX0gsM
Gjj7qAbKBv2MryIaAuCun0qIvjFREMZWSNEPeRiKiMIt7ZsIuJAWtlH3LPao8Sg+
6U6lbXza9LbavD5c1cpb2/MA9ovd1EXc3yDW/kt0WBEI7vuPACgqi/zDi6dz7IzB
AtQwIBlqjPKOd0J0NvKZEgclHItabR8zlJb+O76GA0sCX/T/xOMAaG86jNQs00UC
kZkQumXk9L/M+Wt5aPybj5UK4fLHDGjQnf3yO1aFEbWLgKIkdGHyySY9g/JwTgoE
Kz4qcCRMtxAtOQCLZIXnvealQtRR43sjN0T6EwXTCzbOnthGtqI2ZazqzBm5pkT0
VlBCjBWgpsTDOTdGigKO5Nl0KRXWqhjZtiPMoIVij7nKRZcek5upqYX6P5IPoL55
HGtJnKtYXa+1GqelpaeElFlDF/6VDs1UB4qCP01E0KCYQAC3lZ5efit/0wyHZFrE
UEWgpXt7PGeIIVtjaPoWOD/Cbk4NkQhxSQ9L2STdKZ2vwGEs2yvjLyFyiEnSu3ty
CDYm4St3F99rLjajtIWV5u9yR13sJ48AaNV9aMhjnpx8yMcOeEH7R0aCc+FEQP/F
PoT7G1cZehAnqcz9ysANv7RL0UOEnKTwpHQUhgwExFWisU1F3tLhI16vws2DnZwL
sfrezdk55i49qB8vdmF8lSuDuV2tDq3OqY3XesTFdpra2XqIn8JccjR7qiff3ft6
aEpS36YLRRTa/GJpKaS2g9k0VzIBy0Ql5HJwaN9GTtOl0tBnc+BMLisETpUZRWZc
uGjg4rkl2rDhAre5IoLVECoPil3GXUWH7uXIrYw3YUYG778kV9YeXCGASHyNxI13
EOfaMF9I8OlX/AgGhFx29jQLppS0a10vdCpEqGDhLwgBj9XtPvvoau15YjAyKvgP
kDyivsDKvHtIiyc2AZYpsAOS3T+moLPiZl0ObObHof5zm1gowHCY8Q7jA0j3tvL2
d9WUujHbx3Xs/GnNDEAFDZIBKa0Plitr1eH3ZiQ+jQE5Wxg/qOyEfPtPZQWOz9mH
XStHsZq+n9rulIvJWr3ZQ4QGDxFhJDyKMlO7vCeYIHzn3DsQmUdg76oKdr12fUjq
uQnr7HEiFPyonIdE88Mtakjg+IwEEkdeBEYIWaSYKfxB14d1wty8vZzh47r/DvN8
rr9NY9E/LOjQ3VI7xhUm6xXwrUt81s0D2SEFHfJLjcTTU4dT2us6ibnYAkFzB/rH
cYMQqE8WlvB+LBz6DLMzcgwhGmqQLpwkMkQCfizAfJoNH6LPm9Uha1yE4yfhniHG
vXaOpNu+rc97Eay1WVjv5ztM6i0YFvBCvKBJPUG+r5sBWQGOi/hik7vuTEoz6H4F
6lD8g3tNu68oOq4bdmDUnxsnQ0WgaaXF4RNieGTLgtxhKjB4NCxu0BXNGQsIki0I
nitwOi9D3K+nuD+HKttHycUgJ7Wu0F4FI7welqWqaRaw6mS3PQQDBnu/kp05+hM3
OlvIaeAOCbT1GvKujGnKrBrmgyfdxiqQp1/I5BTmQcH5XUilC8aa7Qk5W9xQ4KhF
fkTrvL3lSReG3RnrMpy6T/jMNBRP6ZAPwex7jVCzcSSDKLbf4gTa0pgPF1lwuTKD
Vc0VkPjGLZUZeoV8DmSenUNnPjet3lLb1DXFgJX1JLpxr9xdNR0ahizJFoMGt3/a
9T5Dwd6dpzHA4NQVjSfOgJq1DMLmhmw6/MIMyR+Y4aLeRUOH/sg5kZIC6TZqZz/T
8U9Tp1cjkSfTImzVXaY/UUapFvQ89ySPu+47jcBzMHea5k2K6aBbk4xJe0ttdoWI
U5cMmmetypUiXBStKo34JwfyC0CS0tDh1XVy8hX/Y+K3uwmeAfD1z4piZaf/7RHC
p9VUoxcv6eO73IvyIHqMp6ChtbONAdYCnSpUgnxrFFUyFsPd4STj54mqH8lwFw+X
HU/ztEV4uN+C2ERqhy+4Z5CtEHO2weXUKExgKdS3pg26zpcj+S9jLSLpD+Kw9CFT
edYaAmOIaJFz0aJbQ3UpGqoymvAEfLlXPGpl7TZ0mGhoAICg/XG9k5c7VUpVwsBq
lVYGorH5fJ1aaBlodFwUJ1nmCFULHjYseyZkpzldZYVJWN1hD9gsirAdKe1Wt36V
8so5wIUBlKEUcJq98rYrnmsuym8pn04H5kk0cl7ih0QvVMSKBCG7deJ7aqBEau21
gUsmuB3TK5h3VmTIuZgR9oMGzF3yqFbC6MIzqoTdPSTqKkrWoI4m2OvPlwenqNdt
hcCwJ8Ch63FiESKoSXureWvD/loEJ90AfIhV5KAzyr6tVIBjiYwMAIeVP3bfPdo6
+kYaF+d5uZCKs1PggcMpAqUmzRSM05GNnUT0SxcoReXJU4dpYKSg53o1HXKdYkve
E5wWlA4gDrEuwicThZplnRR0vQoz34BTDsVgMobG+Kc3OWae7S7C860dFmnj97bt
SK3nXmsNcLJQMFfWFB0zUmPI7ZqHQyXNG2mamllyzY7LTTN2fpBLZnLQWpo+9XGL
dk7v99RyGqW/u7kw8yYz5uN/2xo8gQq81KY85Uuq+t97ZKsvM0+G1JORMg4GVaum
q6jCsCJrCqUUDCSifusszwflKQkk0R1JAdeYAh7XZBRe6nNTGlMAmjhCJajNQrbV
SRmzR3aHLcCq03YMEa9Y6YGpcQj+Lb/QYI3Tq0U/aAKIZUWKsW/Zp3upsILkG/dL
GGzyI46+cz4TbHwCHA2LVFPi0xg7A9u0xQ+UxU/UZZGIQGGZH41zQZS4xL3Fm61r
7eWpse207v8ZYMa6zcaiq3Pw6wA+u1B54AX1LUuetkHQ3sB6rlmSCqkiaIPbI/DA
HgEWF1ZUqCFwfzF+/26b/nFytTzO0rQhYXuK+N2W2JG27rukWORr5vYCsPYU+mcv
nlSfWxW7RbFPQ9WuvIWz6KM2Ojb337t9OtU/Fvf2ovZFR0FbPYkr+rdPQMsO7S3X
ecfUlv5HSuq00Q95o91g3UdAverdYgTYWhF6gk8sbgk0RWZV1XS/OGeIPBfPeAmJ
uUpEXloRxT79GZMaf8MX4r1CKf9HhU8854x8kzr9LY5+GIzDaTgqODIWDFFWLkBy
aX3Eqc1enJulM6drNSOdzT8Jjn/8zJYY6ai2kKdkDZ+RIFYBXoEnEcxN7SDmMjsv
dZ5Yd5Ck2YKvGbWwXinF4hfo5GF3vt1D6d8UDkk7Mimn18dNyGPt7ZvxZDsAcHoO
SO1c/4K0vtLEO5iqhGIKJgrQWBdCR6ABM1GfWYmGYxzargrDliwwLUJ6fF/l/sCR
SqB3L4Um4Lh7V6uDpjdUAJHXTa4yqea5rmWWsa2VlQC1hNZHTI+1F/3IVBgVwLfj
0bmFEWmnV8SMqHZZH9CziFlAd72EOxl1/CMlqgH6sL6TW8fcfRRt9sDphNW1hCJv
PGwrGdCY+gVXGNXh3FEa0tVfvMe1P44CcB7ryVJraHfmXfVzALzROozsx8m6AjqM
+PZFPGZHaHq1PuQ9uNwKB7XPRBgjz0fPYgyrbdkcH7P42RziLynyA4DRW7qEt5VO
7uLxLt9gm8flDjh4UrWL6+AhuG86z05FOH5nobzAM6h4M7XAsMTvtRavCkgsn7HM
JrG7zDiN/utGIhrOlRAPneaKaUKDFdRL+g3P1dioc58VbdRNUySs+LXaBbpAS7pE
etlaoMupU+W3QGVVHCL00Vzhpwb/y+xyXTyDOIkfHiBRoqwbGLh2dm4fRDgpsJX+
9PFUGj8ZV4dMgqapDiA/ZerfUZ/DHvE29AG84tklmc8Vic77BAQ1yMx48nXewGfb
RD8f2E0iGuThCyiuu+F2DZj7JTG6dOchAz8s5hc+yhQQ+8dXnR0Y8VmiKudTtMlm
pZ5qpDJvk9/Co0ca7MN+NIBGYBqRdciEjyfnlzcE0kQH7U3S7/SuRQliouHV9XKH
cHKiyTYY03s5X1l7UNjgsc1mrtf+W6XFrHNa92pY49uk2SethushcLNwuNfbISFP
g2/oFmOKa2z72iNthZmYgjDeFj2itBsPVDy6pIyqSw4v/PxTUpvJQuAkJ4YzHwea
yKoeQPlAFf8H2/PUoLRFx1StYZI4RbPhjUB1XZLr0fp05ju2el6zMQj2qekpajjQ
KZh9UWPGf4Z4rRJEbrEzJChL26ex9AO3Ju2bNW32Tz94mnfSFAZhAjkPttUJemqL
5gMOKxaUg7A1YNjMrDAvMqC0TS3KEO1wRneEkWa5ev3zvMhda61JIYVI6ukbq3cc
bjBa54LievDAHDwfoQdGvb5xoVVNuRNMY9d0VgPrtJ2dmYCEHF1L8Aa2x4b9SouS
fB7JUQYvwk/3yJuP7AA25dEDcDAqinDI38ZPkEBltlxXMtYZVtbfk2xZwODH2e1f
FxN/ag0PPcRKn38AYIcVyyOB5jR+9Gu1UYndUgB975WIclsXCi1E9Cgv1nRPI2q7
rtLUz86tP+zeC6hph0x7t92s63s7JKKLLCluLDV1jDnkV0g3HQnwPZwCz5Df+jKE
XsmjfSAxV+/x9Bln72wQEJSlAHU74Mqxp3EYaY+liuACNB9lJd37d/kT939oJBkE
IyzG+oMPYu2S/dgHaNeghrmw7+fT7FD0WksI/B4wOrazG97AfvsgnF0J0D6W+zdt
7KeOUJqtW979ie4OgJvJ+CVTPSIP3Ia00MVtuEorSG991kE/Ds0OYWWcPWKMSgx6
2+QlcqV50WoeYpTI9KiDV76dKFT1d1XQldS68lyhOkELD97pHeDkYnqrOk4oe9+i
/lMvbtVqyfuy5mpd3r3mNtJAwblO8SdR00MN0qWbz9sB269OjcPRO3KHl8h3m02x
ZRuVdhuCJwF1ZC8zeWpZwpaGwQgjPb3H9dtYI83Q+FH2FL8MlNLVep5mMFmetJk5
1+bbosLLsJKxqEgK3j/wDUvDzxLKHpFxCPvdK91RHgWvmJBit7hES0l8IBghGu73
SrZn9NUWm4JNQgqNTsAn2oNn2QoKf6sg3XInXQoOSUPh2Ei2kO7iq+sTYDgDgv+N
/7IBcnhsg15ezoumGrvWkH5MxQ3ieBEXFaVcGKSAWOFavpOvjpa7lEaXamrthsJ6
Rmf5xNnAwuITvM2ykSM4wOvdO1vt8cMum63kt/EQuFsPG7vFH0ipGLwiqZlveRYh
IESSy77RAiA1ntg7c57h6yWneUs4iHTxH6RJqnpI7HiKjjZciRUYgk1Qwl9zvWDq
StsV6LyrdGImE4n6tCYeNZugudw3DpsfLs3vyq3BW7vxB0JtImSp5B/8p1mLv4nj
iDMPG4jGjbyeYpsklZvwlyP7RnaxQY5BIm6zhv+k+klfyn3CoglK3zILo7cDwyjj
4Iqv7HKiHmgkbCV7vkCk8Gn1mv6Ls9hxVMG24urx/MT9gaBjhXZjWJtIKiXwlB5D
wTMupe21x07DHQO8SiQhV9r5F5vibUHll81jg9RZuwcFrDO/HygSsS2Sp/Cfr8D1
pbkv7hqu4bqv0YLZdH+A4x7/9MguOL6sSraIcjR/AWcILR1qfSFNAygy5EVPab62
asHmjpo+BQZAGiNx0/ZeFlHzgTt4O8eUgKhlmCJGjBOddEk+Mo2y/gpTc9YXiSQp
beEWnBhaTJZcCy6Ejp6t4MKlC9UeVWhjTIFmB8JRyHH+wtj91V4JZtxSYaenCyhP
8xIv4VLpAQTLVOfO1z4GFSfO3C/01mKh9q+UTIlCAY7QFjQKU0Wr6JddBjXXtiI8
ngtp4VOWrgetCPF0RHTLsw2LLMPwFpuAxxUMllUBKiDmb+bXeck68yTlYeWs9sbL
t9+0c/0N3LlJqwyvDI/ZRIpgn7IsKWbxEfR8mpSDjnR0HPjKWozAD+M5zJrETSvq
30Gr41YqZB2xgfMd+qqPvVXZP47BgtTwVMBesTIdCQlUz+YZg7gq/0qKK7NlrMmf
14U0lLxJG/pZeq6fmc2ggQhw+q/92fx6KWKGVNke84eoazHbyWr/aVtivdxUryLJ
65I6GqQoLEqoH2OEPSXi8MLaWtAxynGrtfqhlYaT7izJ+/cRp4lIpGRJAXcUWOuA
FzRO33/AuXtfc7SSu2kQ/qUadVeO4lfKnCFL9xeZCm9x7zOLADhiz4QcqEzLOHir
FxObz48YWtmKQCVAA2xpZJ0Q19z/i23SW5Cz2j7y8qnP9AK/8oM8CNXT9Hs2gyrr
7toot3DA8noTZ4CI8PvmRI6LdjNN/JaWH8MjNU99mJMhdgkSxqNZeUk+Kfio/HLn
9vibHZnAzjaro7IN6AUF150QSokH6uZA7Vy349Zwl7zJ80SPYAVJ92kjkpj0Qj9r
MC/HTXOYAxht2dXbxy+VKPIqg2hnMDCE/2RTvOKxfFxYm6V176pd4XBBD5OZ4ADh
5i7ZKCKCZqBZ9Rk1X674tGDIPtVRlz1VWM+zO6Y8stF0DTcd1IdFWyJV14B4baCX
j25g4AMrkBWwPksxPpRiyrC6YPvWAPXOQfa483hAPGJ8xIXYouLhL5jA6GgSZ7KI
D0fIN43bB8jPXVNwZEhCS/zLRwNq2zBb/lDVrT5xcktRGjQMtvJWR93QQwE4fI3R
ZcCV2frOHeOGwx03PxkrGsGqsqBkmDTeDsgfFEfcakySqzJGDR1oVUkvAga0aFas
GsjbZt5hqcOoZTnHbMGBdl581ANmq4NmyRx6W6OCViztWu7ipGqmen8NkgXGzyY3
JUBO7sD9W0762B5ctR3Q8RcJT7BUxjDxbpwRoz63mF0MQbq8wb5OWM1jmHd2WGyF
yQSX2FNFNiPcpCsfJGvoGSj+75t5iffXg+30FTia+/wVAqoZk+Msfg71OXKUbBH1
b6bAructuNuASltQQ6SqA+WB8uSSzVYAj3ecmskBcyiq7lv4ZUI92U9AhBJr3EDT
lUauE9vfk3i12GLexXdV1LAFc2G3ZEBVsl2dJ01cU9RP7f79GG861WWto4he7G+g
8LdqX8fPll/a9yKLT5MWTQQHwLTxUzbcGpSQrJ+weNFUegfTa3TqC4Z/o3g4r08J
6A455qoIXXgGbBkBjtT3ONH+xyTBTfFRG0yv64F5Bg4WQSvZWJOM0N9T6WADjE7i
Nos47kWs8PHmfIzn2UGFlaNGQ/NyH4+YRjRlI7PIRHQycXpWTgDjPwGsK56KLQ3I
Z9Q87oVWeZIyWwpYZitpRX7Bdh5E4Se1GSaRroaqV8Vvs6B7EFV3NqOTbz3kx5TI
CwnmNYE1+DZIxCRnyLujQFeAm+dvrDTzLepedxRnalz2bmayDHZlqVH9Nf22g4ZU
lEIMdLXSjtiI7td2GH1K0AFyF7KRT8Q/xTGQG7fEhKMZtRR+w4n4pVEed/LP6SC+
RqsUbxa3v4JkGAKzFCe4qNf30odpN3HSK7q/8hpKEj3PK976U2PdAXcnRit/8uiy
blwa82PUnEUrp8btpBBPtOZDCy8aTFmncAG8dXo4DwQEP9pL+yq43NBtzDjGOi9n
YHkKne/4fg5mP7hORjRu9UhsLp29uqWdO9RpGg9YIBfvVFjXc4wtZlMwEsOJiXwb
1/6+XFIcImQPXYsIlFslqfa8e61MREGbcR7XKevjfzF4PnSYd/vXqfodMGZm01B7
JfFZY51CMcFlGQuEgO5T1s8Wz+ODsbYEbYqFlMz1DfwC6XyLIsxu5bzje+c1r19F
Tg9UeWkMQ30rWVc/8e8P2NmSt300lnF4/z0ZoTC2r1Ti0EdgjyLVPUDxQaiB32aL
sDZJMH9Un8xLCk4TnM/PArSnPbvW7aS67aAe4mnsZj5lh0/odxOWhhWCeNilG20F
rMEPbXCeSQWLc1xt7McSD/lYO3f0DKD5x61ZpSIOTDJ3vIQ2jLIGyaimuthKGmqd
GTxHphVdaJW+9G998TtA+gDJyk+Go2JFQnevo+ZH+T3gWBmL9XoFAiFb9ivtBjnA
O26ph3NJH0cfkVWhTn0D7vym7sQ6WjvgAZUbVi1b2BxVHXYcmWQuijGVrrtx1jbn
gD6mphgq7yvvj9jGqfusRZ9vQja3NbQ9glA3F+ZCFQQl9e1T36PU4+4Gi4Igcs/p
V9uUgvUD5856bv/MiKB+DwGgopuFDBFeKpOK4qjJg9mlN/vsvBDbNgo2E7ibGWV/
JT6MisjCdOOWiUJYH3eU1CUcuMkK2zmZmgVs0GKX+Jtg0RlgcD/OQwv1w/7FDw0b
qrlloacoxjg3KTdAI77HGEiHbLn3IZd2qkjmzSntHbLcErVLwDA6c97cGL3nY2ua
Qrui3R9DHjhgPBbgu2JOJHB6rtdMMvuiUA23Unh1odGsvaUn7XagusbxUl35QwZi
U96PWbvTn+RFuUaPLWvsA1Q3ieXSwYIcIXsST29O9AVdbRwVBQKRwl30cj3qMM6I
dBwrN/XRIRcLC50vrUGb3c6txqgNIk8EqnWO8Np1Xmn0VQ8Ug/2ykOES0Uv59UmL
riaeqVfCv7lPrQ2LBh1ctQL63GmukzRxEpizHUVW6kE+1KfOwkH8XvcThu9Yv4cu
rm+WTMvK2/TbYYoRRajV+8zvB0XPRibZ4lQ7yrEvoHt48GRSoYaYs9cNRGHLg0D1
oMPhTemvgA5hoNQ366q3CdsEAogQRZzN9wcUg/BijUCYZNLlsJytO5/6SSwXS/D9
vtNY7DOr8d4diBzyKkn+Uod4ZSNUjmqc/Rr97Vc+O/Q3Xx3HpOaC5aHuuDiaDWtX
ccYnfVDsbW84wPEDuBnTyEiOT2Fd/hhbV4bmgjUjN4abr0kC/mvRGRHBhkIViRRr
23Hdo6b1mhi95LSLrgwNvHTli3Vn9mVrqa39Qop2frEXx86xkutsxSK0vXH5MWoD
VamPAjySAWn5ryMXXN7FfGUHrKHV6EJh0b17w/FnnzJbqH5EjYNbtgN6WYl7+ZQb
0RbLVJTp1n1TrdzC08tjH+uz1IBAm7djRTyuq4NPRc5Tr2vn/oG/ioupe5OvUxRL
WB5gohyO1Vp01qa51skscLykMiJ/Y09OmjnL9noKp76mi6cNI6fftKpWmgHWmwu6
0m8/vH1C47PEYM6rAzaf/M1EgFHZZ1hUgb0Nw3ZH2s9lthcvt07UDp4eYc7nMp9U
zd7FFcMCt0Znj9n4gOrm3K+jCOJE+pyhx5knKpc7yqk5jBCznYTVRN0aWEs9MUMY
Xhw2zsAOCQewwCiSsr2eKq6lh9P7LZrYCBZiAnpkZDthxDbgdwZguvlnjMYcmy6+
OlwfPMYyHfQ18UWWd4Hfhz7CG/vTao4R+161aRRS4eC2ebIBbmQpINLx5H9SbjuK
nzuHvgE1EdcwD6KTR/25uhPSKAJj9ZDZegpgn6Buj8kIkuDMXcuxPyQfdA44RtWd
EjltwOaXus7hQ51KP0LDI6rSJ0/9qWPasXdcmKf5/le03z7bzCHexhr8oFhbrDpO
iGTTnyGJC6jhQ62RTarmLdc+CHjisrPl84fYjRbkXnNN3pzzHiikP/T9JOjq12dw
KmJPi0XtX4khQAzh//79CG6jL7Ntzvq88YyTt50RaTJrV+gTk6WtHo8yWYyfDiTX
HBSYcydvPPQJGlT+Plz+kKxiq8zoBW/WvSdjLMPNz9L0Th+LkTwJBUVjofDr75Q8
vmlENQXkZ9PQOd0g8RP9UON4M36wllTHLiWXOD9De3sS45c8wYQg5mhJcoTNsMZu
pmkrmpkt9xLF2GPWzvoE8YZ2YL2JvjjlYMMSMxgABidNCYAXz5Oq3gD0OWDqkpA2
owB1PMxzuxTLcYp4jh6Jw8/vqE3tuNK/D0eEfL3c3iUkiuKdZLFKw6gamrfV4Afm
/3xZpt9FAmokMa+8fd3t+CXFP73ywbDzwlL4t1wqK6sGnNxIMb2jnSqNFsqkl3YR
D0R3lL3uV4H9uKm5KjrKqV/eC+/Ha70lWIoAsFSEiB9LgxKOtnT7iAStnyVPduLm
Uc2W6DmlAwlQkYbM/sciMn+fHtrJHEopl2IX5DppKu2ADxXIVWbWtGOn8RBAn+8S
ezTIIqtYQs6Ea3kxQuaX2Eq43nWlSVYMnYKBXTaXXIclmDZp/xENBcWnZxrKHx68
8eBbzFQIlIseDxwZWyQ67cCCCOUcStALe5mqfTARRzCuEAUQbdcQoei381Ank6u4
hJeOavFR2/sZfNq9kKKPJpE42Z7212igvz2NdADswZlNdr/ERseX6A4m6AK1Q9ec
5AdbPuDzDyp31Lc4XwYbLuTEhp4dOP5tcNxEGXGBQBmbLX66W/+alXpT10UvU7+I
bj6u2UvAb7Srt6RZxrAHd5rdSAak3/JRf/wzOXz6J0PWYulYaqq8Qx/a6Vw4czQB
n4tR6sf4Cr4LK9/L7PXa4OWL+cnBsTP+eUOQ3jtmMbBUJ8c/x05FySE5qxGo+sK0
48XZ+SzUjal0P/11Zfoxc0BEAB713q8cgwRP7gC2+pWJXdDKO53xZofS8xx2h2YX
fPR1L7H0ZMAjM1yKKaTujqn9i1zrds5Ng9acxPEl+/sHiUU1rLhSukKaBv/sKTuE
GD2TrA0xDOOXs0uZjs90jFTyp0nr3Kf/ZAFO0sd6lC7u/nOJg64BclaogQJF7kIf
SelZXj983/A65ZHhk9cA2ytIrF89biCKsAdj0SYxEpasC/kW0ENFbLDeO7hhEj3V
sGcI2zhScRVlRUU72QsjS338noS4fVbLas86wR6T1X91P8/CcWlcxpGC8ytfh7D7
ELHxyWB5WBz9ClW3onx40yb/sUU8NjIirZEX8DwXFAe03Vrhr1KcJA911f8bCoJX
LejbIGHlOZ89pk512wXch4ZuWYv6y3bPWMzkXSzL2hmabvWv98OWXE25B89M46eC
hKsZJMTS+pmSzcUSiF/tKWUQ6u0+3+jcQRXU4sKa7WO7L3p84KoPSQKj1TUOMFjH
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
O1DWG1mISaNc09wQ+MgMW2ROHwK+kr2ryrJ8dc1Gzn8ZnX6HVs9doS07f85AG0kn
EUEbz4mDxS/17MYYzevY/GSHsNEyKqzl2LUQyBXpFyA8YarNvhk2XZTATVym4IEk
47YHKaq5ZpurX9VsdtAXjhg8+ADYzQy6hQ22AS0xwLVAVFJDRKBV/kjlG/vuBurS
LC2tEvWjKSpuDQZ46kn7r9TI7FJI47OyeGAngu+Sc7HOe6osllHo7Iv22fSbDGMw
irbvthY2QEKZ34wenRC4+tnR1G7jd2AqfGkknBr0tyvO0EJHRi2aMKHpievotXtI
wGQgiFUEZ709ZbEMSBbI3w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17376 )
`pragma protect data_block
mXB3mfeMsA3nmIG8rBdYY0tAw+rSD4lyXWg8MJ7BK6haeerVEskLw3WcPjI2HYOk
nDDa3xk0LY5u8S2LPfLPhED2ydXaCWJAqNCMAz7qwy5U2/lFkFYd9lrYS6OmUO/q
8fwkLEWs1WAHYUyjv0C4ZlSYk2oGTd5FZADGHoaSabURjOvDvqLU4oKAQ0uBYj3w
90QtQhV+x2ir4N6WOJYk2r6bxd6p4rKQYHJwRkugLTp5xp1J5eAz6gpPEFTRTZHZ
uxl3ijeEr044CT5vaR/8O8h7Czps2a98P1RB0utlxnq2rxCiobjPp3ZQr7yUVEl+
PO3v1zURCup8bRVSiTkvaMpq6ax5BFyeyVkFyGtzF+DF1AYkgu/ok/KGqn0TTpCq
Ubi2wi2lTp/WENyyCAE8zi/ejbfPKdnkKl6PXSpbHrLgIqrxXK1veHfedR8DPlbW
nEyI3neaxiFQNUt9tO3KdXBHa1Xd9XuvpZJnofPoVqgyUEa64L2sdKcTwWap1nsj
ibWTyepu/OVz7mcW+eTLfnrZCIlOsEu8BetcMgixVV+HzCzsoevNK3ApRQNy8l5S
aOMA3BRF5rxdUGFqWyDjNrR+yQt1qb23dRTkxgv3akYo2beWV9FqmLvx6UO+/nKl
/22HdsuaL1VAnUHBCNgoZlZa1aOpkIVdm0zMssbxjkCIOv6/A9zY6dWAFPF22nOR
5pNzPmECO7XNTyD3e3VYlvMnMRpxTlrfF/Y5O/MrdCumGKqN4ddhIe5QdZjLl+Cb
C9/kVI56lkXT47zp8DoAjE4SvHoJuCmBm2w5OzIA7/D0vYIB7BA+x/SYDilhpC5L
AoRNFIL+UMif6Gu0zblulpfWUcHgt9V8ZSVxNQ9p1aW3I98fIHINn6mr8UKGeHHf
j1eAOucD3MhvF6dEzaCkD6TsVlbOWnlFhB/IoxQrn37+4Cu1WI/1HR7plliTh4Y5
6D8ytE0hZgRxKrEPWXJ1H4SUwYT/Ok6EOuqHpjvAGimzU6FRN0s+Gez6bk2GyZwB
poNXBhM8d0QBIpMmJBA8D/rIc1tfw3IF6H++5Z3MgP5PZMAXD3HkiV1FrW/cD+9v
yz8HBwi/+Ncvclzfhz4YPjw4iGssEwQoklfIjjNm5ojCjynne49YBgK3KZcxhX7w
GDxAPf8Hk/dApwvzvU0Z0A8JZmGKa6dUCWF8F4Ex+UdcPiH0csTkwwAqGl4wHtXN
qBn+5TQFxwlNRRWoTocxbjOW7xVcBegnQfa7tM2QL1skAMrqEjvfviq7SlhzMMZW
KAcojoCbb+JIICguXdjYikzYRvTvnmMVKpJoXpWz8fV2RDpJSqQgzuF0ZsKJYrWW
WL5ya8gmBSk5VNY6LifZCmkRG9mG3GxlOF8/gwBmLGCtzOzQq9NDhvDPy2eXOthG
u51iXJuWXYEMdxS936kTsm6vccrm7sXjI8HwOyg1jjgSSbjENTavXC8o/L6Sp6kQ
Aq9S5lGWYA3Yhyk+LSIhJfcT8Nre/WolrNIS+8/BNQfZYXfGYIKixNg6Krzhf2gY
g6Njvi57bfC6P/12zozPQxVLEtp9ovtVuuF25j20VJoTH5+b2y42jiwGLQw+g/py
Q0lryqHjvfezyTPML+35K2+qoJExAmJKhlDhKN2xhBhlzOt8uC4zJsIJr9dgofLK
gsYSRfxAwR8O9jvSdZ65t+OMIbZAQsBu6TW3CEtGt1CmMuZJKASQT+jDpEXAkDGH
315ZobaRr+0YHGut9v/Y11V7Afcn8lchHzy/utOstQRtrMa4xAdGImvmJq+o0PVU
GN3V4rHqcLw364fVULIBFQwXcdVxVHk78NYFalHCPimOiKl+fboHN5FbDt/CnzgO
9EcrzRXs1u2mNWdVp9MJooD3aEpTL8sYUzXmsbOlsAfrDBC7UOkPWmDbhRxflgTT
5uYvjzX9z+gB3L49pYGFHRfDhR52OlE2yT/J16eyFNnnRhtd+QgUSYRTtU+UXaLO
5AJHfhfH4sAmKR89PZLBLGwSiVp4PlyMjacgpqcaWFKwHK104duzjqBgvOZffaW0
hhzmUAwDB19fY9NtAwz78aEZQ7nlClk32iOgUimGpubkMLATIIwMqqI1bnv19G4M
2eRe4LMw7Hf1diM3Q0RJyUXsH6+xhwcIkSiWuwXqByTadPqRvV5hEUQPv7fbJKtx
LsMA5Q2R6UWdkzwoVx7V71GU1XCWOTjuRu9rf8ylNYIoJXftWz8+ByWRXjNPlpHu
PVzoa455oARzVi5kkhz5AznTFp6A88JFBCbA5ToVSbmwOQAzO3FV0FCUSKZV72rh
y0srdHD3Yd9Qqv0nMd6tfwJ7nL57dUJpOVaAfCQGr6//M14/Z4WClT9RWde8ixWF
IDjhrBsNO/xFPop2V2A0YG9RWj2TQ2qMf0CFUIl4Q9gvL65BjfquVbJ3b7T8mnJA
FS/iBN23XAvOcl5DfactyCcS/pyyNOVw9ZV8MGUwJOcv2FPIqrkzkDOCMB1BvFgQ
POLJ7WwKZ0v98UPwi9YKZiLtf1d0/OGA0FgBgOStjWJraKBph6nDufXwdFqj8tdF
Rl6V8Tyn5O+h9RQbhN8qVhHI7tRm2nhojqO9NbFho3uaMr7jASbe/8yNgN/x8JOH
+VaOXgNTV3L455b16E1lrY0votagpI6pANA49z9e97DurnuB+HouEcMDvvgXv5hd
dar8xr3z6OEEAbb7g/e7L1RxcbBtJ7iL7kQr/xLrWFsHwDeJQ8mVUyJnQF5uF2dx
t0KEMs8w5xcIumhmQfxJ2J/z4bVcOKnCIht2m54fFSw6O1Ip0FO3S7hgdr/vwdzL
avS5uYZXhJ6AgeFA8xE+GZvpP2pt6Wj+6SJUD+0Ex/y2EhQ1T403YYSlhOGrLIfV
8fwAuj1d76oBpOSu51xMUNwrPyiO4ah8MhZivQW1r4i3+tbhYjNF1FNzEvgAQzBR
FZaCvpmVUJQgAOYBgDUQeoIFfFLmJA4QomrbKT3ekp4omX+rAR6IIVLfzySJmG+C
DAb3g2b0qXhOkQZjqjQMdI4Dn/uevgZUYEUQfnWo2whdcdJzQ4IL7uvhX9JwtUM0
tZoUKFf4LlqPFPeWrxEKaFtuEegNt+Nqgct/hPVbQKhnByTKCQBRK4QzgnOoeLop
xijgklb5yQ0u86tr+PHgxUZy2x/dFIu+8L5lBzCctinAtjBh6IgizSWrjRQalYKI
8B/zYH70PKFGuX1r0zVnpNYls16XE+QWoMAaPE4KOPVtdHkSi58JS62IjXHFwcVV
7xmAH/YoWy0kgXlYMGm3xHWj99lMCS7Yu2P/r1Ohwu7oWkzAjJsBQe11+TUW9DXZ
5g3Kh6FLx9A2ZKzLGOIiJH5EuIAR0CIqZwora+15pijKSo8zFvQLlYvaFgwkh5j+
9wWNUacefBJCbb/AX5Wq8+L6vYDVETU4eVCj9mNRgy5AVFWkX/PFQR2NP+IUgf4y
2cmHS0McUqDDEWkyGWTetePc2n7dGUGGaAZvPp/H5y9o9yici6Zn1sqTbkCSLEfb
SA9Qda+hfj79mU5o/FO0x6JTJKtykshWb6u/c8j0yoiERi1sFWp3XpdAHC+et1WC
3mreYzc942Omf6/d2oT6OiAK9IpVqdiRl8EjO4ockzOW57oeIRmQgSsoc2MolG7b
DuABRXU2bOBXOVs0SfUrRaJCg3gungi2ClZ5oiw412S8tby8TOqTup8KnFBgaAq0
ECJRzRrbxqAfUhFXiODqPVbWEr2YeUOiuiAZvZ7MgivQ6wv0iLw2azPrjyiCIJMz
OegYP2OLoLxYm40HXkV6F+vnRMMPhIK1uYqJgnF+xSLXAdBL/cv/rxrhA4seKsfM
IJfzpBLBRqHkpJDB6oQlo+7SImWG11WosyaBEVwgKAsjuqcru2CHyJMi24IQI7Ed
xTnortow68LzCeFlX2rOdzWtDwcNgij3Hwnq9IV0QTgst56U5S3t0Dx8s2EbKRjj
ykiYaAH1GAIO5iKmMeixUqaP0wdCp85Be446UoFXXOIzBt8gRx5jTYZezUWXEuug
FO/wUWu+OrWNPw2kdvLedf+8ZetriJaEtmKFaX2gG503XuZbRbXQtuUh9PbcDbRG
FBpkkee+tZTQTUbyFAImZultAN8lH9AlnLTH/CMyBCKjnSBH+pyjquslErGVQtf2
Cst0fYLPpyITnMJW1k87wJgEGXxmPf21HtRkbzD66STb5Qlt6DqmF0hRYjK/vayz
i56BBZ7HoN2361UYdNFeIqQMTpo8lnFHo7JRnPVgGJFMnJsYoq2Njmh6gy06vsRe
yde3MN5iPj5GAvh6GTKZdlkxluklk+nCiucKw+ytq7Njl4cr/QKICZpsNI3wcwsS
xmxHt7i0MglJgfVvVY3xFS6UxCGqR+ga9BBWmriX+5Td9nP2rQ6KP2jdSgoQ69XZ
AS/XWElq0Xny8vQOLyPdUX9QhMH4pAhST93Fep2MT/E658tBVwVm+odRdeAx8uE1
pBbaPVDBG6/dYUOVnCOquOzMpzbUr8X+UfQiETiSvFE0Ube0HMmmLBmh09csqeeq
bBIN6L5OrUKnMy+9qXYHbMSxIeJZ92nLIu1+2NZZOPJRqx2uNvW8CyX86t334YAo
ye+Lmj5tuEIUrOAy4BX2wXNhpmJUWRKLFIwC/o9kVr0fbtFUEUuEH/Y3MNp9GMaw
sU3zfBAFc5ykVS/qOx7K2q2Z9lUcraXz2Wnflq3cqDHQ8lQdDShtfH6G0q/+Q0jF
4USfsbFFIvKEYuhohTDAixpi5RkChwNB6UfPq+SvAr1ka8eiw3eANkAjGcfPE9O1
HWWpLGs6uM6MnJarJhERsOMviOdeRnR5VFqx0oZ3IP8gP5YCQKhBDO3DoJ9HJZ8Q
mSwxI6HsIYyT6k+o/HtR54diDP3XSG6Ukp5j1hBJO0iju/YP/9KSRJ1oZm/LTWBN
CjQNbok4xqCk2RLhVkKKu4LBVze/MQc54uiIktE57bFizBydnovDcjbJtmjI30et
4kp3Z9u2pkdivIsx72yXG4zC2j305FNUYSBYR2ZDzWsPiFv0NYJSggKADXLA8d//
RFVuUtkW+HR8/Xa8YpOJVNSrZUhHh3pNkPm5qQo7uei2+e4n/X4EHSbFNYAMUEVA
P9AWvEutfgfH9FXHabGkjGjk0O8wXoRUgrOVFFRxucG1Wj7SUs12vDLwTxYbu2qq
tV2/IgghEAq0n8/ozicD4II1mSGkQto5gDKIZL0zX5QM3tMzpCP/pbTmUAeYEJiY
atwfLRLjGmIoYbGIxpdCjIb6g3ZCERVWes6A+VqY7+NSWXq1HG/O/7PGs3jBWFgi
Ye0WSz0N6xn2TJuMQasaYFlZMBCESZYI0tWHN0Zm8oaoof67T9A6swoO6voY9bfs
CUJZWcROS/OP+PejKOOAAsiLI1rj9pCNPeYjsGRmiAQ64QnELTU9s6O9rsraSAy+
heNWvVmh4Z8CYKOu27eg2O0tYeWeOsCoYuDcRAkhqEkRhGHXSNAvSIB8+/iIcsr2
u3wpOgV7tm18A70IVMiD+KA0I19pQIOliADHcVWvCMr8si+2bV7p4ol6wwRu3B3J
XZHINDzJfqz6mR3qn/TlpihQfIsbvqduBzRSuSClRpdSoUDyzRUW+G82q4BOo8ru
hzgIjm5WdT9LRD5EjdUfd+MUAT9f1H/tVJF0hGpZVNelz8cN9YXfsxJbw0YCUFua
PsGwh6uK1mVcuuImptLYoSVqJLVRkXaJe+oATBAryQFJ57XXC4NgUf4q5qEeKqru
8CCh+eoYDoCguJ0LmwngvBjsjFLv4W2r7Q1T/cHKR1xibAsNxIFh9q5dyDOxcRZ8
hXnTBNWJ5YTmXoDtzKihtyb39HqY0YqzyQ+RteGSvj/9nt1+zbgYdKJH7D200NgG
KscrcIkQtB+5J7t68LvXA1JqLu0TZH5zcL5Ymwih5ynUBXuUODYeqP8GK9fBzYRX
IoUTn/TLeD2kc76JUNCmOyqUJ6Wm1TEhOaWjcNQ5/zEHP8jivhlakO/RFRMspSiA
16h7vss/UgumDuXHf2tKice/K6MElROgKsjOGJf9tsv8mvuxctIKw5VJ3juVTukj
hc9y2nObhTK/kjCFxQ1mLnKPXXb6nrwdErud1QccsG7cTq6yW0GAP7mNL9JOEMVg
YjuYbGBMdt2fETPirCpMFd+f0bQLIBgOKkildWyNm1tefHquMjL50V3stAE1GYE9
5ayfZIN3pRmRUDkkRgbK1ZXrQQ4UbHv5ZpZxpw0b1bMhqt+iVmFzoizPKgupgkuD
OX9uio/T5EksKoVO/BEqOgT24V0j9VSwN3xniV7kMQaMfWD2GFggq4Cr6GA8W5mK
F6lZ3tPsWMDtTG4yaPyjXx4gLkFFk/jqNnZT/aQIp+4ghUMOuzhFGea8CUIduPr8
2a/3GyMtu+i3Wc/3UGLfR/QPY/YHcDUufdVH8PzxE+jzxucJ6qcTvMPzMzJ8FBvi
dgeMQwC2mEaZSjCqtp2IKStFFBKdpKwCCza3311Pcx+n4mwa42k+zCIPaYsSNY95
oLeJdyH6XCunuaR2T95tX4z47c6xu9iNG9zjNPEQve4ueF98wClRpeyG7U2kDgnb
1M9dQWkcXI/yZXWGcmiqBRADcb6kRj7SnsL3MN44I0kzPU6vNbVd8Mh4fDMAcpzB
TtD/oydX7HYcmroz0vOwa78HgmRndWAAsGEmBP044DssBciiuyP87nzde7LpboHT
ZQCdQg6sc3C/yWnxY4TuFR0g59wAPHGqE3kHKpExTZBji75SA5itHV717CKnDmzS
ZccFUjq2xi4gxP8hKeHo6eJxImRFpCOj1xyBgJQ62MHneWM5ey/7wBq+MrVlZNry
ZIj9hn2vZq/p/EuDuPDNm42N6NlVcwwoTJeNfDCaSEkUUFYRv1SOUmEumLE9zrwl
GZRFQkTVSU9LqVA4DIItqQZSFAw4Y/gey3uqVPdkI8FPCou1KS4ASEhTRbdO2BwX
58xntMEDjy29rlVs+Pk/9kCxoG3AOvy1sUbQrAfH6yOtC81+wHGoA7O/ooLfH17l
Q77r7a7yCxeNEnyt6gB/o95BZifJp+WQxxqLnzCx2Ty7ZJrpssSOI3MY+BHOSNVX
kbdYta3soSLUn1fLW7l9jCgyFUro3s45qDfHoVlyfEgXpjbxt8UiPi8Fi5xtRK7n
9SHuyorbW3oRd23IKU1jhykv7xTKb7xHZTB7PNrCHXnWRdkNMY4OXAW5kND6cc+2
I3DnS+31Mr2NgtmNBPUkquqXnw2Rja/f29xX68SZ8wcDEkCQNkXDY72CITawDNk2
99MKdu48TGDIG8vH9RxM9en1rmQZiNcXJr9nErdxozCnrzTJV2r+VVlA/FMT3i9u
0U5dSQ0Fw4Oh/ekUxn/Cm30oRzkWRxFg7pVwUv0pVeYuF5H1vTAKQDNjvvqip1Aj
w0KR1tWgyEtwT/smDL7GJH+MhW0v0Whzea9JV9tHkkP7OcONqU4qrbJq9FPVC7MM
qoihs3u/yEatsGnO51CbKq+EsgPfqrJAYkwKt8MvZOP7DyQPM8YgOM5+l0VTr7gl
ZHMrk+Vl8RhUoIg1w3s1c/sCpm3ZKDqrbdkCsUJbRLUnjgzSTrsdPU9dKH6frhBt
ucNjWImP6t5da7l5n3p+zZTOPF30ONzD5eKcYb75Wdb+XEuI18zW3Y1s5ikU5wbx
4ajLCMpfCNHFbET13SQutziw8oybp+nJ3Ilofil1LAEBhD/x7HgW3iBaFRSCHf9m
qo6fwDaA6u/ycgbolrqClDWRsD99qIrQOJrLA9juZ547fvejdziQ03kNto8Ewzfl
YPaYUpUYoWhKUwmuX3H8zuuqPWeW7qeZ6iD+zGBotb0P7/iRYjhUUI9NcUuxJ2vc
nHxnrqQhgyVZ9sZXL0RziwUKnAt/PEcihXiUZ7vKIlV2HTiaQKSCACbqdXJWt93j
U8+xg/dWXpUMjHtG+8Ju8xVEUXQMRlC0E9KP6dBIMz1qOBHMIlJJ+duOS+xXZOkM
ZeaXN9etaQX2ej39lbSnFQMoKLCDE4hWvxvOTmGepAxKmSLXl3mN7gpt86yqTjCn
nERKw54cbJm+lz6IGFvu6+5mpL7bPxY2Z63U3f0VqNTYmerU8+7yyi7IEUTi7/LF
Q+oygmoiV7cSwXpFx1lkqtLM7r50flczJsja3HtxjLhslzwpsGFcQxS6yaxuzuEO
dYtUHNUxJh6U4OG1UiSqymP+1sKgBheJVAZKcn7O0Y2uw0K9rt2QJxb2vpW7HSXb
pwSeZJkpOgzGOJRUJmjqcbWPgVXMp1fG8iW+0f3GNICzn8/ybu42Pb36XWT+ICIg
Jq1/sPkQSvEOE2RGgOCrtygcH7+Prb+FnySMSOLsLaO5h6p9rt9n/H/ISh+7WCUd
o80WNWvvuhcR83cfIgfDpMFNuw078+rP0Ct2NiMDT8K+IC/dP4nByJDwJu2wdRIQ
Y3OhQthu9Q6vrnmRJeBPqoPTQvzq2tH+CmMnOf6GlnpLnBP1D+JOqseeJxTQSLpo
6ke3cYUYUkzfLIXGLZTZic+L3OXYpheCxoxa4AT/NkbmODi0pb/IFV3jP/jc7kbh
519OOxGJKCQ6BObfI/mnpulbTyJ7uyyp/NUm1QQZCweE/d9b4A58Q+hbJjxnexbd
pFH2dzE8l2nKuibHklxoRA6Mf9JZfWbwexirB1eqW9GOEw+rqSB4pbQ583GX3KFH
Z8MCX2ue1xutTEyXa4z+iYXHuVw5j1FUsYVUqTNaQjnYW1eIKTeGZgk7AYDiM6cg
E0yOmwSWgd+LA9yv69XLeykAOmIO67JIzFDrMd6yMg0dDKyMPCNivsZPEaoygpTQ
wwJQJ0C4AOTDJeLAwAwd+DmFxWCLovSIVcOTQ43nJCPg56iCVCngartLjlXEgxF6
+HF54RFhsKOFVeXDYKhWWLrY7JEH+1lPZLUA4va859Lia+ntmEzRcRZ2cQ1IhPnf
00acgcZzK0HAMirc3gLQmTs9UjGF5d8y9o3CVYNPCTTUJSO+oOcm3+2YB0OaTFBi
aKhoQopdYSANH7ZkFSa2bAJHDdtN/ZXMzDBP1l/UfJKSlyBP5bJTTSoUnLSnCcd0
pOPi6wirTF6kb1Vk4Ukl4Eqvy4m/tl1A09O3TN9ztl6ZEiKBD5BVIveHuqkk//FS
E4uFPqIMxSkG/D2BWJDfckGsr4mliiKgY4Z0o2xbI0kjlfXzf1n9VAnsGRWRp3Wr
MnRFo/UBFMcchDIfeQKwaD1hwjlYwffL7+7afZid6ofxwTZ53MOupypA67O+gcJx
bFaxp9KgPWJNbpNwvWFw0olmH7fCRnImgZt9RX2Eg6HJohvNVGEncgJ8k2LHMi/T
lwruML6oF5NgZbLCJseYfabgMRE3g+9CBZ92exz82vSPFJNDB9KEUaTiju8PNwMM
5ZXp1rEGZHYZDSIbtGyrAAACocIsmCuJZ1MF1I1QoCHMezNeAZWpLQjsRTZZMZoE
qDUCEDOND17bm6KmSVHKef40TaRu/JdaLywumF4PDIIIn64kqfBjoax6MdPmRZ+u
6Plg7s6KqNJyIIEMDaR4euyi4Qn/nEWBsD0512CuChMInKLYJOfBR7cD1B/kNg/v
a15uwsZYn306snMQeoilXJlT6RWpqrnakGC6tm8Y/OWZTaTTMSHfCXm+7PSlTCU8
vPv862raVJ7T/UqTs9oAXTX6v9HnS29GFNLT8LsK8V1mxT/Ma96mi/almMKfhFYa
2TD11z690cnP8XkErsWdbP96ehoUyloZ6zI95XwkqVftlIGuLslhTfqPHMFZELkU
NO0EEHB3684UfRP4td6MZkiS35IiqLNm6O7cO10Mo6pFwIHrIqmzBgLeNnpG+Nn5
NldMcLFbQsHvfN9cHOJ2GtBXlmZ1/OjQaVudUfnYUBsKiVOCR0ETMT5fh2l8bxuz
io2FDXbEILVSRxoo8jq5vet6Y+vQnVP3+HreMg25PNZwnpCjSecUbFDTxEV4as0O
CqCYftA0sy3kQrn+qMgqunlsj/1MjafzOJcq4WBlK3ui/jcAbIKMp9nxm9EfBXDq
GiDpHPwXHUcE1+/ZlC6w4DZ9iMiCShxHCREcTGoQIoGmK7UztP7fN6w4PaNmnqfA
HqK59ReTpz/cVChUD75Ti7En+xTHvkys7plUQBrxU2ws9XNvLBKbWmj3eOilD/x9
Wbjin+e9fyaJZ6I4WznYzFjkCdw9CgiLMPHYKkDnzVGpqqENBqniW611pJPe06JO
vz7984iY/5Fvyed14gmV20weJOBqvwNn0PdkOHx1e9o1M5+nEkd9SItM66W4iqRp
ddhXRuwKTF4zI5mkwg01qT8GDmr8+3UXSu5Ek4rnwav7ATCKVqcGmWYGTSwLHx2E
XMF9liQuoQ6gHiW+iX3Neplxlyn3QcRi1anwb9l0lD/HNjZ5fNnnsrEPS2ujmFso
H0W4asipVmvMiZSqlgeahK+H3leJEYMuf+N2TZzVHt0rDHbTgpw2q3iibutRA3xt
uUN9bCHq43tnL1zr6HhsGlkBd4QxjzY6VCr2Hrm/wYJCwz54h3epTXp8+0MNE5da
n9ZHpLjQgSd9i76TAerkw6dzhIZpiEI/nqvxJdFu9cdSmE0ScwfwNOc/W4fshYdl
1hqQeeg3d7ZaSUxN1MyKDa+UUgtdT6bFsOWtbOkRq0jDrJuDnzhmXzIXtsln76o2
0pww6NfA0vH0ucRo3k3odlpEs4CcsiCfYRtLGPNFS/lJhpd1wCCMzuuDXMcRF6tj
9ywO3FiWc3ATWOZo2Tv7395Y8Ib3MYSrVnSb9UDXIK4VF7k+i1Uc4s4AC4LTZiOx
y9mGzJzKUj2CosjYz4NUZG5V9yZLeQMvdciRD50cC37cct6RoVyDnU20QYbCniww
ngW/e7DfH/DNBhnB8lNLKmXYuiqwDT2eiZjl3b155jvj1RNYdOWdPCs6/N6m5YN7
XWbsFRjEwqeVgQnV5wKlDBzB/2ypu23Coz9JmB0NlgSXw4teeU3AbnGjoEo7Usrf
/HiUPbgDByW8O/vynfHW9yNPwK9Pi0eEFiL8gBjjtGwrhccISIopkxz+rlZGUvZ5
trsGKO8FWm3Eo915CkISqu3f/gpcTckpxLH6AQyGrKqEgh7lVFWaGzvWEwjddRbj
fxgII+bcxlEqADPtlLWZsh4mE6J91g9RtfJHiIn7ZYX4wV+6l4h5rXrbifcY/wiI
cf7auGGDrbeCHYTuJiteGNG/Bx+WsdkcBpj3MFF72gza44qrNR9NlKwhprWh5UaK
gXu7C3am0NEaR36dtCPRMtJwxyAVv522xyk8+S8B+gh7RyPQp8rgV1r/m6G3TZcp
RXialbV1368dlWF6ntidsekWwVqSo6v3BSls69UjXcdKyvorFID0oAPjrEB0Sx8q
arz6ke+0aKpEf+LZwwxxLcGfqUBwkuoEZdK5dxU/1HSN7XgO735kW0INC4frxl8h
i6wusDBz2TyGKGbjNCdRv1Rdv4DIR5+mQMh6ibP8evlndWFoebrgLXOyz95EZUtt
RiK5SDLni1X3la4DUcD3I1ukJToC7Aph8o1b54g4auMLFcU91NO1v5IHTrp0h1kZ
nVzPy83vXAoeWThzsJKI23/EPDwRkl7dYpm1f1efsquvjFm6xPWpFbBaK+VF5eYH
kxd5Fvd26vjH9JMzzULiEnYOza0KgGmWY4YstF2/IgHILcMp7050XsjkW7qMUI3e
a7ZozRNJn5iFqCMgTKgbxlz76SwFOeMVc66KhgflbbJzemwqcMCzWi95vJwKGyhi
Zt55ViE/wNCVlssUmubniHd6UV0IbfKKfbNz6TggSF7O6V/7isA894KKecdXOwZt
RE8T1pU63C2cO0HMqUKsbAIX7bCS+jUPtjbTSUNa0fKgxqCKFRDVVf2lROFIYrR9
Xcf82FwbVcquWhl1831r+aZAWmWpU3RdA1u0sZMfGByFGT/KPJts6qPVsc/qyX05
mj9ZPr1KSlGbUEZFGq1ASc2Ib8H4Vdc7nr8zvC8AiptUcDTXIMFXMhxrQvPDMEI8
JGYQb3fviWkPSMkruQlAcS5DyeBuZUuUHS3VUlDfbtTWqXG5X1eVMRVqEf+QMTBt
RYJnONSvk4zisxv/L1KCN41huEk0PRfB4k3fs9S3WW2+y7Yy34fzU6DdogEfRyfq
/zD/+AFVlL9Rq3DEWwyR4O6PhFiY19u8hE1T2uUgpUcX0oTZq0xhCFm28+l7O6/C
C2fn/TJ3U1Lgl/c7yQlPDO7Rc8h+FIOgODNUdOo/KTgpU+vRZn4Q3+liXf1cJ6v+
hn8SXGpUy+xpq3SUG0kJ2td0a2dakJab+O3pmoLcl7SVqu4660GtTbqXlcrEt/6V
WhX8RXqVvpq5RyM197o3srIA5vdQPwTzzQYFnNUPY3ZjyS86QTJ9eCNjLXzQFQ7S
dalx7QvivWR/qBaK/94rznHVijrFrHmXZ+mtMPmeK6EzDo8wO5QbsGUR9jYF3qz1
+Dri2+pGNE6xGRzyN9PgkXlI15dhxWfDdCK0iZfNI/XjeFzrfm5Acx1PZV8nXOS0
leD31hRGZa+xonnJeYlpRuWc0SZfdOWUrpnjiPsDmCxPfXquiW+U7kJkpHvh330L
2Yc9Los6tibIqhqt07Rlf3d+tvlzuynTqyX6JOa3caIwO11o4SDp8Iwojst7rinr
izb7nnt43DkByfl0OtaM/ri0qqgnJTA1vMoz8D4vUNskw8azbMY9Y4WdOfKl1LoQ
H7UOBDmig1MF8F1HOPRNldigyldVJDXSItcEPvD54Sjn2ze9NMUgGftPFy07tPxE
SNztnRpeQBMeNDP2pW1mRUAlEROGs0m/4qOMfWjkRDQaHdSN8/n1FaLJsUq+3U65
cRmcqjkHH4XEnKgTnJELO1FL53iS+fe4rMu+AT0jB4BWJtWO2C0UF+aL6DFJPRAn
CAyfBMO1rMD5Ao6iLH5WuDPUKAV1D5fQvA2MgcdbPN52UBy2Q5a4efcWk42/bLj7
2VqDV3KZBSjaj8N4AgzZAseO5/QV3AJG3fAE3Q2XzhKCtlkbR8VXjMKzHJGBgacB
aVu6rhYQ2EvO0EGkDuvKT58T1l8FoBnSDqeGdgFtxnWftE3agWWowzzdywpSbTcj
0bokhTzIpX60jaGpzZsO8fa0L8o6swHzOM4EdLnCDqXpq/QN3q6CqT2G2St4ETq4
eoilmGEs/vxW7NEMM5YAmhW6162i2LsmmpY+fzuqVqvzRLmL43VIiuGC0m5gJsGR
n8bDdEbzppZ2tTroyskYL8wFKEeXfcUSZdkS333dvSqr0ElUOMviun+/molyGfX0
S2H1E8zr5ZUTGKd12ed5cmYTdlGj8H4RSgoPn7ycNhablhhD1Zx/vGh9msKYoFxs
wQR0cslYiNHd2weRqHh1ia1Qq+VbvIwyYHAxelOrp+1iEgunMdtnT4GAjOw8J4aS
MOOrMKwZDdnS6CVJ7sdYtcZYyk8Y/y8278VUH2BTtpmrMj7mT3xLISvcYFuQEpGg
09y31P70w2MPcEFyJZrtpAqnyJNmmihN25kbXJ/Se5P2aB6yZuCAhQcbDgqETdvT
4isYnkf4cDzjdKNE7Nww9s/4nrGgCbulOtesyvJ5N2dnARQ09uFG7HJeKq1pXaLM
3Y+z19+sTs/NbxesS6UhFZOG5+zxvU97RYhd/KmRnno/hLWNyqsW7tnggzz6VY8+
MAqroDD/zYoO8vhcJcQKDf3zDrzxD6ekyQjRz8TJ9itxM/D2wzug2tnF1G8nFBZY
cmPpJIkPPYBJn+hTsXaYZn+0i5H89sY62OJjQi2/8ISE68XT1kOIAkU8zHFQizzy
lHYrzCcwHeaxvFuYKG3gIqi1fkpgojOs98Vu4ws3jdvi9R9cGH3kAzXZiUkk+0Ut
UblOYUj5Rp9GUT43NRUQxXeLB0OiY6XtkzhNuaUnGq4tqO/7I75GZXDHCDabaxht
Gjj+y21MkiwMc6uyxwBbE9ueYm0aWeHOvYhEP/nNVz8ZAgsaA65CxkNZoNUt2208
xibZcVPZCAubrX64VSAqs54RXH5vkcOeKEvxR6lgOh7qQV2EwMeWJtVG/Pq259p6
oE+6YeoJ+o/LIVXptrcBDim/OBoi2MMBtZ01oh7LpITkVoFWODNDEtB7ZJyuKFXg
+LlQZWt8pQKvrz/ZjmceQ2zMKa7QuknLQR18G0t65btKFWECX0MpmPhn9PXOYsqF
jqRYDNGlZbhHh4lGMvdFoTxbY1pz14xR1bAiNZbkTdfUCaNh6BQ1GOpQq0CAYMSa
2nqqaArTR6b1b3qnoe2MID2du4f18XxnhBnBs8zVplIs/7Rhbu0vnzMJsvyXLqeq
7kt26aVItYP2F9qDyJ/CiERSModYr9mFkj1km7GgIAGSaZcFgRTzdahqiTon+GiW
J9ELKYu8Hk2+yUBIGZkVDWXQJsRPR3mNAF4jXlOXqEhQQyuSmu4qM2BO8GKuZ1FP
Tuq/i5sFw02W+YNKuusbaT+AvuTuem5s1sdkNnIfrhKjaUmEx/FXzzqNjlvd89P+
2pJWiRHbY2sPkWFWPs4hT5TxWzGCBotlsVy751BinyZt5rQi7R57xXfeRtZ3lrMv
G56ALN+68/VmrijHbPN+Mpd0qn36aZ9yYKsSPpnndMCb5NbHCJ8uEQEca3IKkeS1
nS8AvUq6RWPWHca1g5dSGRrz82Vx+rmkp33HQSpyz2ee93LeqTtYKTDzBhJZi7JB
KPyHKqGBJYTgJJy5GrqxdKbdVUeEEz/mABIKHHuZtq+QknJD9u2STe6jb0Iw2kil
92LgfgldwHOiS8OXkG3BXUGs62ZaOqXob7lSAgCrIvgPRGj3CiO5oJkWPd+iTE++
V1Zy0V3apVVKcVKp5Ge4zlq3cRrF0S5OVE6EB6giEqtb//YtxepCiFubZK68Br+l
TA5a1scNNrXKlo0m+scvCOJUwF0GhX0VnZAddlqmkG01I7W8lbmt1mNZ1UAAAY0F
vHtwMp1BBLLjzMYRI5npo2xSkEP0d6zNGtrKYtJ+yYK+kAbPaP3e0SVKjlMBzOap
aqTUIQwN1LXmtU7JGViIiyV5le2TKt+yZiaPwdkURl/Z3BDUNOidnDglG+jJRvJx
G3uQjH7nOcrgImp15rskOS5xjDo38csVVwvPNMgOs02EQR1hBvkxBBuwP3EXmN1Q
5vlWcD4z+AV8qrd+mH0XlJnVwmpzjabYpY18/dm/jRwLtmltniWFtviV6LabhMpB
4UXYB58+csmE6H5Imcy2CGv1UMspCKtvgXOGIj/9JIVeT+nVtzvm4j6FcU8eCAlO
Tz6eRB8NRDOduxcQFvPSYaXsDaLlTXIaL2ikntTgfXP3W0P7Y6zJEJCfZo7gDTsd
0eb2VqjaT5FuvVGQZdfAORhteG/+BRQ7dr2psdBWpKzRztrThfB0oqkEMKNfk5/9
/NrF9SakuXANQqxdb7Vq6EHiLf8PhqUNqQk/a3r2/7hLLUUun7lZudIz3UOQlL95
4pnYlY6YINfzUaku0junP8cJn27pYNWtlMwK9HKcmLu8rSdiY4q+Lhm/q5jUIpIg
WscXynW7R7MEjC9mxQek2Ea7FJeWmh2i6/0ysgj6vzwoCcZhLZ2pcszRnap9E5pv
1lZMjs0ht/ailBfAZGa9KTFlflgmtrg1TgUONavASg3/C+fEeJt32H12JwMxQWXQ
VUEzFWeZMnDWdfiloPfo1uCTjgzJWXE4b3YWzNWIml8GdRW5T0PVThqmQRbgUdc2
tMZ6d+es74a9Zb/Ff/kIzBaOkw7E6n0BUBZUe4yZaKobBeeEwYU4KlNp9b4ZXgEX
lk3JJunJvwNLP8RMfuZph1CMZbCUv90xa8XyfAR227leiHVIYkxdTqGuizEgJ/Pw
Q0cpqR9d9qdgyJJVr4e8IkWb9gft+dVcVwJsQJs4RARtooWfn/QU4g61p6SWQ74m
DxC/R3hf7Z5piYdkpghQDflS0HIi915hNxG8mJQTxUAOG+OhcCgGBW0GiEJPF3by
0lWkCWDd9uxv/dNTgcy1+Ms5m3SSOU9YjFGwv9hN4epNERRkYh1/CWZacpTuHx2R
XGiEJ//qg4d6nZIN2wbHSu4lWGEOR9hm10wzAUTzOryD8GM+ppKtjQ+kIvwMjoe3
h4EhwGHS4T/fTFDnq9j1KPFDNXmHUDXdFmx/lNE4mvgG3iCv5eCgJVGvC8WO8DAb
WfWDJ04wtjqctEcNJ458M5CD/D2Xfl5+qlN5CrzLx4J2XqvSSoLdRqPqYqOTqXfg
LKrQpxjoJHQz3EHDVwKSl3Q2QF2QRiU/ICrvYPhfOsmXC0d08jR8Bd4j00ib9af9
3RDfFDicuqPEOX+7U1ZrRqPvUr5YBOSxsyDl5fB2A5pu5PkKFFJOlv3CzOGrp2cB
iXlsk00NSzOHrFwsyJvBjIAtpVCBD6pLAMR3Tq+HfENpTEDAhGCIlqyEpQv91Bsd
plbCcm8pvuReTD0xeqHSZCTfPnJg7niOaeNb14ZR+YrdBF509CZfaODdZB6EubAC
CQBIqmfcD51rd164LZCcAtztpJqV0DcXiW/YZQ7T6UmvGuWQYuNHfA7D5iwBfZUu
nyoLdg7WYOvlecbjsThcWVNN9uDeWqfo7RojeDZgEtwHf8HMeFy2dWFAX4j7Ct5A
j2KMKWohU1ecKNXcjX8b2pMXmzVEyw00TXTUbNBMmoN1oZdQDeydCfN3/UtpIDVJ
M4gOqBhE4tnPJ6VTdfuEnBwKK1tSXYoUMClFaHUl+XeynOUiQqj1zXYePF0caBaw
EcUxAqaxqAmqP7PBudvwn9KbJ8FVRLh2maMN7jucotMinFnZNC/7ibwC3xNxw+PA
xwP9lzE9kIWOPu4IFp1itsmrQVAq8u81zZJNFv7TS9gOUxmk5YxQeN7QvGcNycQk
mqm6CX2lCdwsWCY2eO2NDxwv6gMVbIGgy+CGyYEe/dSCOb/LUXHX9X1yoOwc3St5
sK4Mo294Th6S4+FPilMkdrlYtLms/3rVerK4JmvMinipRP2+A3U6wgJ+iW76UctV
LGTnk2OWyMsm4HISlrr+XQe9l0r/piRPFNaoGab5hS0zbPB42C9O048oQuSgWTqe
rhW0qwy2KFGxlGjLzD+dAIgFL2Xhm4SUPV3/Tg2G6HELJF5JMDdQwwug2InJc3WP
DrM1iwG5vOo6B6n9zPBarudoHieo9ATtSmjDdMKGCBGsQ5PCKjx9F1cYyBN3xKL1
wfWTai6kvrEwOA3UWtpgROQNYaQSXfr+DnvBqQSJ8m3e9EGDLbJALyz1jxvf3ayj
NiYJV+tGceshx6SktKAv6DaviLuZ5GnNVnvT5213Y5Ya6AypJQqS7eN+dG12cyfq
nGowt61dgw0+uvrmgdhWtaJa5HZ12nRXDx2A0uLWgD5JHnPX1KEULO8zyFQD+pU7
sAY18ZjPaAElMTv5uQ5nh0qrIsmZD2ca7R2Qp61+FKVmacOk2eXOuIwoF0NsyH3b
2FBoSGFzcInPPSvkqwhttdqKKwiqSTZnlhNM6VGrHyQ/20UQL3Iv0qR3/LWGFXc3
wswQUrIOTsH8gxEAzWF3yUadTtWNO1pRd1cY6ht91j46Fw91/04xUMRzWZsXcCC0
KjFcCq5fEbQk3Er9cUfQgkYwXBhym//2Ef6i9LNX3PplQwJ5mJ41YDzgmm2F0BYg
XZNQciG76PXng6wylkD8eNssU7dgrqKloaSfpJIaa/KjNoU8EK9l3Arf7BbxPBEB
J3cCApFuIyX5rUiWYVjWf31BHQlG3jhUnQQOdmj/r5PIzBYRYDY3iqzpVIS+R5sG
qMMWTDGi6CyFOzuyuVgOjxPwm6dSQxnhwKq5mqqjv1d762J7neCVTXu5R+htuZ4k
TItTk0UyyCjKcoaN1RC/1vqguY3k7Jdlvf0+ROeyziYLq9hO1fRVH9uFk/HXjGJE
VqvXso6u0pr4sqsomeRKmn+9QS5CR8574V0HG+Em7C9YocuShPE0RNM55zOi+AZ0
pRk2lrmFeCWFYpb9RODGmexxVOfF59EjEwiXFquZQFIBkaTf8R72YsmqxdjPbpb1
auj4eIbmtO1qDNLjOc0VK0DS+cKYxFk7pwXKz7Oi+GEf7lnzmQ17EK2mjl4AJMvf
su1zVxsRIgfEpYNoI3WdZp32b/zvamzy4Bqy4k6BOK/X4bTUj8IQJtSmR5GI3Bbr
UDPutN4JTEFvxs0KppjIp4Tr1batqO721alvVheZzaWJ8Q4G2ZMyYfpmMzwLiyIJ
lee5VAJKccNQnDrcIw4qJWzBxx+OstLD7IR6x1QzWDvnXPJWfW9CpAMRRQWecd0W
YAJm4Kr9rqnSuyHVWOvW0T/DATlEEa0aonN9/BMnKQ1pi4VPNPgrsp5kgd6g/DUA
/Ouix2nBVmWadprPndf+lresO0868bfEXBO9fTbsR1mOTlNm6cTxxTC1F6TPMSeW
lK8CcrYuhBKVy4NR9dDFtRWvMVnopbfPboqXqagA2aN9Y3K3sYizwx6Qs1lRVAVx
Tnf/nPdaX+ygNQ9IVpc7IeMNrlk1ZVUHRPpHuoSQpF7K437t8tBub/1V1xPjISVp
ZNwii9FGgbs36+0sLwhfMiilocIBPURzR4kWD9VO5nzHeLELNjM8be1b/nJdOnhQ
dla/XjMM5DS920eSjxlG0op4Q/rXsjkDAHRoWoozEbpULVZYLLowYazeO8kIM3u1
elb23md90LScJL923bJ64T+gL2GV5QCWEKR7b8v+BnN79swFjmfM+NRJIMLFzlcz
625//zJX9Di10tDMojO49kgqXoOiFM+YDnb67q8bAMfGeLyQXxCDoGAga1f1pjj1
yGX/YyEaeFTsRePeAg8cISCOijfDPpoi2GFMEYVOqsakFBYpvViD9w/4gDbmxM4f
eosyyU8GE3e8JrkNY6APxSbaVmjua0VCitaoa6SJ/pSTv11DWdwN2PXtKpqdRYcF
16dg3ui+kDkCcBV0E3Nu7hP5Ul2VSMJKFACO0nkqkSMknOkP5OzqK/5DcDCD0vo8
lq/EbDLVaRC0AKFoexPX2/JiOtX5KDJUD1Wy76uCQgH549BKVyukxqPVrCm3tCJL
kjTqZ0avt6+O/LMllig40wn6NywDEVug24733XZ2nfqcRnTWyuqjr1tRgIRp42qp
GYqSiivd5NL7oKo+HmJVTEWdeEoIWiubycoDP/URZVBP6qhHm/wSrLEM4LR/7jAs
RxaSfTi+1neq2ZEMtSUw1iTQLJ5Hr6KQ1TdLIUqZcP0Px0JCJS5Kl0FeaG9NiZrb
CGM9dowrSbkrU1GCDerV1cKE0q2r9dFHEJI4xYGVyBzvwYVFaT0GtTKszvVrCp+F
FkKCazKNguvXobQ2t1hb2TNsBXDLKYClm1pukQjWTavwXN/JSdq697xX/bnRFPy3
/UimR0SEMmlfe+YDBIlkuRXKonZpzJh+GdFNEmdIcEP3I4NaVmVEnB6uxgotg1Ux
3kkyATDm8fTPvzZ6uRtOwiAz15/Fs5C9MxvnLKdjFMCRZ3YZHePYs2kdhgXrIRpo
Azd0H370T02ggjMg5XtW3RGUIwjHfjyNvjwAcjE4Ul6HE3qEoSXRrJZjSIwzlmkt
brzx4bNDELhEToL7antpbZx9nuHmajeOu0p8vIBp9F8mSmK5BsUZzFgC1yDZQEyu
QSsrGFM9HFZGG8+OHj/Ul4MfvDSw3b/Wh846CPotmn2rw2G7J0gXsmo0bU1lrNcO
bXFxUgbCN3v6EqJ3yeWIaN6j/X+T3epDECP84LJ49kM5adDa2ksIK9MG/hRBl9j+
4Xd1fFo27JB7fUn/ol07I8hSh/5Lr1XAjpvca+SWi4YS5syNViNPnMw53RXNgj3q
2krtaqU8uLq1RHuzNoexpKbuHLL/qyvrmdMn+jYDm7PQ2ewv4lYOYpr/tLiQtL0y
fQ2jH4g55mJTKmqaQJq5bE7Dvaz6/TZvC7MpnYNBOgBBfc3gZ7cR5lW2aZTL+36C
PaJaUWeub0awFYmY3rb+5bwouaKwFeglvIqEZPAIdrtJD/f5hsMwUtLVf58dt2T7
k0CzAsGjs44qL97MNQslVLtX/j3dqCMm/EdV4jrC9YDuUTXuzvGO0NRC26/1OYzV
l7jbtgKvt+JVgDuJyZUbvfKjjAnaF7MnNoltawJKSJLAmjgGidv6e/tBXtNoW1sx
Ws1Upu8jFA+i3FZnagGqGOkAMyeZLGuqGh7hFH6VBJ4bVp+vm/SqvwIOHPtPYV1A
9B8JQUdqcVPiomsq7M3lj9EcY26mt8wfKb4JF353q7rwOfiOSrQ5fvNhvVbnN4F6
XPRQbymTFUlDB8BrDSYncstjq0A/A73dOS0pLkz0JVmTgLrIcnbjZuufsNbwIHLT
zM0rybtyfUtVJDHvZb8WMZWchytPeDJzxxOIF3ouQUFFpShuR7098ejVjM7osZuq
rw5KxrG1cg6uAQbzQg4NIfNGJlmhH602oRh6Ze30bRApMOL1Xs1QIeYw/hXDowMW
LcFFHMsMvYL7+VZYN37ENslOPsxUJU2UixAJ2cSg0qJhrz8hpchKCNDUEt8UB3AY
+EYYOaxvD5PXt2VlAKp2YP/M221CYjImV76VjOPAK0vGXZzXEGp1dok4Wn5X/mPD
J3mWZJNsDmVY4yLykgVmpM1gUTnWcDl1YMfTr4XLn6V2GoLh1PU+z2VgW/o88omu
Q9aJ5HgNBgSulsYfgH5FGjxScENlH3rbrq0UvcafKgy1tmr33hAK98bUetwZwPDJ
ycTLpMKcvZ10wf4owfuq9ki9OCwtQdAJX9b/XE+JYZ+7AZLKfn/hiZZMAIkYdSfn
XMNS1C43+PFb6MC34Dv0cv1hN1KiitRsBBcGM/iS3xNT52rsK4TBOWbXLmhj7pvq
uc3rWaD77S+ZDWNDg6jPHP940x5lHBrlw+JaO4VTKzOZVodkwvD9ufc4BTktaeaQ
qiRUpolznUWVKw6lX+JvqNuJH8uL0nd0E9XLjifjZtYy7hyIQ5E3bjWh60RaMcHy
KhSIfyotZFLRey9Oj39lW3x3vJy6uVX5pvsMXHYUgMfJYxIZL1A46KIfq4gHj7Ba
VKkdZCo/AYzTXV0Jg4BcczsK5+TELZlORvyNnsZ3A2h3wzlOvaESibK6TUYoo6aN
Gwfs3F5Leb4GKU1usX+cCbM/W4aTkDdiyoiidT1RqeVnnhhuZmCWjMeoGR+tHokE
m27VdUD/wi0RfTke5chfPlE6mQze9FHtE2cUR7AiZdatl4V6cupWGGEwdX+2br9D
vCoYzyTUZt8YZQwE0alfpa4FJWijO2+3lkiNjz0CCXJHIOrwU830gR22ijXsxn0Q
lVFfJ7M0ckAXAHpC6taHvpmM915IG8SdSgICyVHSnJZ+tlyg1FgJ4Pd/gUk9+pH8
fDcDZ7fA5UXpRkUl6xgDiKkaPXcP9jZSC8qv+w89e0rftUNol6CqLLdV5S5PIlrR
L1pcjko4ebuv9agNY4EFQSnkoP1qqzRESLG2Pusx1XdGAYdFOUreI1FyLr3lQmM/
IQ49bqTlurxYnUOXp+yXvEGDBabwwQ27KJNgNdLP27jT7Uskf+wm1V317B/arq0J
wOycQYfFju4q7b2wPyWT24SpV0Q3oe7W68S2qKozfWYUXpbx49Wp5XIQfg4ZnOBs
XnLokF2D6/k2MITw8do9unA1bMSBaw7Yx3Xg2B+zYKG4JZjAlPxxamoLs/ysJevz
jwl4M00qPWI1sJ1GtnHtaVYRVz2/uGlZYqfTmzZacY+1ipCsinLeyCVBmTGQIyWI
BbJb2gPHo0G6GRuutCDGErJQHrnz5qk4H0o6ZD+S6gWvjVP4I8i3xSL59G/P4adC
QHqicD1V4lqoxae/v/5MB3lYOSRrmDdep+8UzanNNQet5DdjWDQnhc6NlXHapevJ
CDW2AGnUFtbAevXFCzNy3qpm7qdLyeAfjthKqSKR4UYP9LqciYNysJ9Z+8OyolL/
nD7ikAKe3WYlv9vPHhdbgPkK89J4oJICWsvpjE1xm/B6PIs7NgnOuReNpj/aMkuw
ooDtSAGmdBrlx3lSoGOKKxDs1SUev8/FVETq+JcU5zWFSQdUecfMurpAGnOCFwYI
DaaKq9EbQpLGnDTRU8CCpr+tm11IDXtYFJbxoUnLtvNrhnTE2gLgVctxqK9+nGy+
8MJ7WZ1DsQ83maMfv24e9ZSDqkQ0VlaSH1/1jWjwiub1gCI3wESVm7UvM0y/H404
uIyB9KtTTbrPvwQPaJMrRB180ApSB7bEXb4Oem04OkkfCNsqTDZ2rGKxoyUbUd72
+Kz42cL6OWmtKWWG0pdaYNGON8CRNAVdeewXPjX6W0S8MvzRjFBNN+XnZ05eqThP
1f8hksohLaPTWCP3Uri6ISgSZOabIx4YQeKfT5+DW6oyRLObzPrWwCv66WJNcK1T
V2PQUhf5uTSslqiY0X3fDcN/WbaQ1zQ+JIzOJm8nYKU9qjKvMKoi8tLnWlnOfe2C
rbGeJ3lQEN8Eg3DMaBcrhXa+xHotmhonJcKFPmPkfD/rGM4RfIdy1o+vLAvo39Ol
RYFcrFv1zYhyAAildWG2ET33e4P1LmsCSa0aWB/uSX+CUsGq9sbSrP1Udyk8lAoZ
7956Ei/Cc0gEpxUnbU8oLV9ZhItR1ItOC5L5A9PueRs5U3afJbWT2WkVcI9CWxvp
JPGNQQAKrydGtcoLpwGtGGX2syXAT6ku70K1aeOp35QHylPOoGfcyWgmh0V7NJL6
9qttLMIJtuvpGnu4Jk0pVJfU1xezPvlA2vi7wLsCBP682u3ScWtlI+aiavfZBdcv
vblZVkU7Kvt6ys7J3nAGsW5pwG58AueSVKWaKHIMshjFiHTnMlbJ76ONDSn4ltpB
xSUnd88Css9KpfeMNrjqdETMmnepRvczQ1vIj67QvvT8ESEYxXhcSxUyv0xchq8G
6ERl8uSseUQJwWdQKdYwco0NMd4Ys2sUfb+/rvlNF2Ym+bBFMN861vi/rEF6BvKY
lJh9Cs8sfxKJe/8e31WTuPRogAaT014NQT+whZKkhaJfbB6LSk37VlNODqKisTTr
nfPfHJc3FF2JuNpDhj718DcOwdToJU9Ir00rFr2/G4GpEIQ0tf4aXPKgtlbpNyGQ
rfnvVa4BgmR8GIhP0Ug+66Ri5bRPqt/e73TF8dsBHRl+5dChQ7N6NUBDD6XpKX/j
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SvnTkHman6YMTnk+cBDV1xU4d33T+0XWh8nuD258zoG1ArJRDncI5o3IylD9SLts
hY3VGXMoRp4J8tR+5FXn9BI+LvvqFMsLPKVFZ2jhGZEGrWJHMgGBe1w5bk0cpcjv
twEv3Mlxc9qgBD+IZrgMMGc/BzFL8Kjyhf+QSz1XxLc0cB/cO8WrVVNfSErmEWIK
ufbrTNV+SGumQMtUS4dlaPhVFO3/h/TSthRHSGjvLQj3c8YT3PVk8EEd3PF+6woy
YnOdhI+z+WOMfJEoQjITp42RO/CpCu9/e3N7z1VeZwYgy0cFQunKbKcvI0OHfoNc
jbJIfwmJFaw4fuw89Pp7Ag==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1232 )
`pragma protect data_block
+TrGvGv3asTxSHkVmATQCgJyOTrAx0iooc2ry0fV1JBzp5WQ6u+bHYFjl+V9wktl
ieAafsxlw1XhEcLLeoBV9ROgyv28cBKc3JB8rRa/I0EeJaG6vGx41yCHoGYk81fZ
R5oanLB4IZB3fR97d9WmrJXrPFn0CCddzWUF38zdCX/1g+v+kSpbkU9Bi04bXYqg
URcB5kJQAg2zps1SFQgiEJf//8luA31pnZJQ2QNK7sYZt5v087zem/YE2CwBhXpM
ajVeNZpfbBa+zfjXWhzg8mOzjUXZ1s7ciJkgHfjPpLCg4vtmRyc+Fha35ri4OQdX
oCa3BpssJ/sgP5TnHSLsxtKUAXcz13sirgRyLVowcGDZ1HegJMkOwLhGnGtjZOs7
ZDhRpmKeRpkkO3HaApmZJ8bQwDkcWE6W1hB7bcQKipd7rAxUG/4iZw7Gd4SJIRSr
BC+FEDgqcS8DgsSPwF+liSXF7tyO3aQXZdUXac+b/UvOIPr3Bh/DAwDOxJ2Q+ZYP
LJihKWSORvjM99Wu7kzOS1YNmkWQuj7CNRPKZ85Zfh4LB8KPiSCwVG6vzT1/bN9G
cV6DcNHFHzzsmSliHIq/5rj7uW65lSVNr8ru4C5r1z+EFb9eJPS8KScx3QadMakn
V49yNhN7PEosAq/l8H6cq4NzXImApa0+xbWka4AAaVJFoeRQ3tdu75sNeuchAvV2
EsfkEJRaYPI6fzrjpyDSoiXb3t945sebNE750kp3Dh2QxO8pDwStuZg937la2WE1
YAzqtcJu9c5Ud+EhKM0VZdeC7T7tNVRkcBDN78kXRwioCXRmlB92b/dx5F6GlG0l
ms8Z+Eq2PjU7PDXyj3BGjbtLzVLzcQWrGxC81jtsQBRA8adgbjTtFm3nJT0qLRLt
OyU5YNTAcSIVY5ROyBkvKlBJHXYcnkXDBilcuyALZvyBzSf8ynHDiUhqpUo/3svj
dfsOzXPTxiDagYWMXNvHbliI4t1VL4OsZUNU7wSnMlBGd2T9Z66txojNPNLwXNQf
+jfInA7zWbe274EWJheoD0dDro+YIVPOdLbRFAIwD6gjrlW5Oq2ALFaIL5zddiOV
PKFHfKXAgnhtDAtjdBX5JzrXVtsIOyqYNi1XunuezHV39T/7HJHX1SyShbD1JdAh
S3ti8hx+kmO0fx2ct2V9hlNBk070TVQtdLCMV7UjTMNTwevR/35xBeXhTPkbDHtK
VEZwIf+EwUhdxSlxSV2yGPXNvp7cXUsmY7Am3uyhvt39aLeDSaGAy1Nwxf7N+HZg
wqJnndhN7b0x+NQ0PZOQF1zM4y2f0tSQ9DtXGar4E6xLRW3lkpzv12cqwrvr/bo2
0Yb/GLc4qMnCqtp1Vv1JqtQJ4sysRns9Z4Cp0M89yOQQp4O8lekYUVFcP9k78isP
VdBwQuAG0LlrC7/S6fa+so+lKonvUgqqJfX/QWil411DQfVWOiwcfri15uz/v6Wa
+G+zxPfKM/QnGNtCx1Pw02DSeLoVbBXZahkNNgzl9Aadoefm3nNNYAxa7Afdpiw7
d7svfm4OI4k7g0oJNe2pMbYC5M+/tzLYmHNlcKXfmI3N2g04TLX7Opqfy1ZdvEq1
uQkZudpkyVTWZAhgS0V2L04TwUc/BvFVGF0BKj4S6w8=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
mFqy6QSGhPPI95Khu89/LfmJs7YJZ9HwXqm2ezPOl6jemtpJrj1lSp9ZQREi7wxo
K4yfqal8tk9Hgxr32yu600AuDWuqGbsIHFMmBWr2FTA7RFncRM7tkd/NxR5CWaWO
PHFuwgzKqcOi0/7uzqJBAMKWnY9aqQIJ5PdzMR3zGgz4r2O2WOXzhn+3bAa4Q4Pp
dPduqU0gvVnj6IbUkTgK19lQdn1uWrMiib4O0ZdsITdCv+K+guJdsb83p5eVAcYW
Fy6Fhm5fcY7KzaI28suQcW8KSEX/dgL1f9nUf82ABk58Q6MVouU6MoxiXaRnRqv9
+cDqDNMLItq+6BdjrujWMA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 12144 )
`pragma protect data_block
kypcH62lcbBiXO9ut/2/KSfkEgIFiyb6ScLA+9hIZeXOgBjAoDtfcil3t0/VCwiZ
dBjTK0dipEulCR/FCfMikHOHqNZn9aA7vMQMS7DOq/5Fw72IAOYPPvytDvD942GB
cUg5MY7dBa4KYPQ893NhSULv0ZZ+NCzRJctEjd/m52pjnOVWFU0ci7frsM8bDPw8
nzAk/EhVMj9TNqfucDSlxAZXNcOOVlWdRkOhIvzqKUCxQfRYmTE0bBqZmH++pFTB
1nV88OcOFCIYnWcsbd2rGnlHSjlDjkUHF7pRybUObHTjgq4uezYYuG5hprcYAHmb
XokaFyoBNKV3IHlX0NS3655dIf8dzghsF6J1T9clnKcwGUqIPbUrsDrXUbcbSRmj
1gFWjU4zoyT1QoTXkQYMz38QEllbmhtb9UC1lBn86EMue7sl0mygwmjsszgZ853C
RwBLTwJxb0X0EflceJk3C+XwJfUGKjzEJj6iivnnJKOPSh9QmYFsMwqON40G5rRZ
6z4NV5rdLvXRQv5A3HOTVf+c3kT9RwdvadjO35gzWdGh0OAZI0TFBfEqTmYsOe5X
CJCfsE4mrNFQweuR0uPpssvuYomcSb7kbW40gclMHrrZMYChuVhEB/8SYs3MADvB
pR6Rhg0FkFeKrg7Oa5PyeGI1Rr7pVUHAMGpp+/SYrJliFFIjoqbIO72geUU6rnH9
qmvQLsdr2oC9K5q2NaTp8VEGaSOXBUJtakU01hzGL5cIuDUpvpLTfc2DQp1xi0YU
iJzQcKkATvAloeebFAgOqMXZXbWdrKfufSuCH7+t9xab7jCjFfRDE0o+lWT3jYlO
TCKpAHpXvTugcL8QoPJ+qsx54Z5jOKl/rgZrNAbKtq8kRM+ENKmUAn3pcZliUIVA
2Sjrjfk68wQXbUs4nmw1aCLW+iOoym3DNdQts6+XcyuRkW/bzvdylsmoIQnnHTzO
6NCaueNZyLBygTInWmthD3S6zZ/5+XjYadT7D/GjZ0RkI+aR+OxOgG8njI+zhbI4
3cb3WtWD89Cd2oLwj9g0J9SSaSaRNEH9eBToWC8s+VDyrH0l2VnKHFLYBWpN6P7u
TL4vSwZaKP02rkDwX7FRN/sorI4ky4IAVC4vWuyuyF0bvp5IZITF4L0J46oQ8O5Z
hkjPwNKGPye2DZktZE/6ocDSYKZugOwE63lf/N2jD0/STdOngqixrWecc1yGy0Gs
h9BscrkOLZ8PhguoGQGB4lHIaubKOr3xhwbhp0DNAbhe0W675f1v3tiZ9Zd+EZn4
WWmK16kxMCLf8rMVVwHcpGKzWJ4d+OSJlTNlQEIfjy+R2cUL5/zvtsQzD+tF20lf
EZmy2kQOc4OUobVd1hXX0IRy8cu8II/zSQKvsjLJlWvKDXWbFCKEzCZQ+bZT9Z0Q
VRx9fTcKBI8Jik6tfiP+rmloSR1Giv+MFYG9ttYUO7pp/HlQQCA0C1+tNFJxMK38
Kr4zw1AhaXhW21thl3kP+4Dw7X3fSkMBZKsgSb9yP4Byqsa83JbnNQXpzQq5w9yL
5dHxdClPWtXKdfx1FBVc69wYIsXn+MiEr4jDuvXf4V+rmXJy7SlsxFLfyy5wMliH
8d/EUa67s/aBKljtuuGj0EsnCTuk+9NPPc61IJ822vVpLrAM7VwpDasXVRnQQZQ2
sVgiGA6uEz4ls2DehpUPeBZXlaGDZ1HD/zMOreeoFjxXuzxe/MdDOZQmX6Lx+yRj
Mai05v72WYyjAjC5xI9h/kBOuVF71gNzvxn8lLB6yfoGB/WTwOifH6+lpIRHb6Xm
xD98j2xuszpW3DwVggT5DW2MM+aTs2UjHXPEJ3u00Z/D0F2qNIlXWfwWYkjLZIDZ
B/1wENAuOGAJPVwC8XgPDCroR/c/ARVRl10MwJzdms+nf/AR0DYoqzfME5V1qaMb
pX6CCZarflfclpqQ4Wgp/5LXaBx/fQD5BipwUIE3zbdrD4e/wf+CVi5fZ8cVzsUS
98edZuBAOmhi31kAbh3636kyEwhT/qwYtf44OPorXkplVVjMvxKDG5I5Q2ieU6b0
R/Xj/EdNZP49isMIw4xEO6uu5ecK8i6vwzzzi0l1cLTikHHTHrsiQxeYPgNuVReu
n8R6Lrg3MEEJ6PbbJT6ylfgvgim5RbTSuOiIg51Pg09xBWr538yd70auZB5ql2L1
sUl7g0XwkmgeN9Eutbr7wt18HJhYO6h/eChWLO2NtIG1DO+osUGp+psVGsxMoeIy
mggeB+58TDQUXaPO9cEw8YEEuWWvh5dkAy/S7aAeGwkeTjQkMekyy6nepRifZM55
T3V02PeaQ4LCosHX2eC4rw/iuINKX1/Ns2hL4u1TvOYgg5VYfnOZZfWC+ODmyEMM
vHY4RcGL44DPM8v1YKMjyEcrsBsOA2dKSIqCjwBxA5E3uiX/fzRljUt+Er9zaqeM
n9gudtbqS7fG5Wps2IVCJoiySclmsjYidNgvw0vMK8fQbPQfxyTnKhlEEss/cO4e
dTEh6u8A1QrE1wluUNINr/uSVsgd32UPKJ1pSE0La4Uq+nsWYzU1ywOJvPY2l29b
vyCLGdv4F2+bilzskNkdcxStQ8PvD11lr+ONwCz+K/Ss1V1RtoEceoboHp3yxv5o
bMGp3boAf2/KCgCN4bW94fsByOKkbteghkFhl10ZlpbUBHNvaIjymrClayvVqz2G
yNR1u0oOc3Dz1O5BnNVqidndxxE/8AmXSYgjFBUnboSQeguIpNotSMnTCDCfVG6O
JzA78XDbvxDBSZTpBb8Ds0ozmdPT/KS0oG/Gdx5VvbePH0mLlWP7LcOo74auzsjp
wEGxxv+wGrsyYLaBwAKgsu7y0PARYDKa+YAwwwP8NMsqO0lXgOVNOPvk6Xe4E46X
+/hy+dlm4Lib7kpQBsN2d8ucdYF1PdH0tAmkjap+aevQiLJJc8dkwJ+2zFd3UQDM
ivaegclXtSVA445VtRL0gjeLBe2yEGKb0rbvnlHLDEzzyFxEw3HrUxcSb7WZMVb2
aDppTi8OpBpwZOXgC1qOf5uknxAPbMap+iyrAOFBlkC2rk6wqwTORBcMTapItZJj
Xwu5rzGGwjRl0GQlLHcSveFEEd3GhjspGRy8VQyOle3zFAGEc9LyV2+xqCdhwI3n
vWKXO5vM2W41uf1OIhHW6IA0ID1YEBJ8tin6YJC9QbEqOCjvYoFSqBXKpCSBq7+G
LYVpA0YWFDfRlZoS9zJlMt6onQScf3BO7o9G09w+IiVzMcX2kAy2hI44QMUJAEy2
SelkOx9ZI5fuNQXAjR6EQBlvFq8kKFRyT5WeWleI6huMqdOjEXHZnec8k8LMcNUY
xs6PV/DfnzrtvMYv/VH1Nv4EXbSjRQb1pBgfN+NCWZmMf2XsM+uZDCrB3vRt96vz
06N/bbtW9pFcAdKAPPduyDwYlAZBpTIgeNPugDI2DB5k1XW6pEMy/464rZWu1Cp4
Nm2r735sUGQKu2WkHxsonUSM9qOaHPQ0D1BGvAhQxPUb5+5E3CiiUJYMKrJfhUFZ
a9yOAN37S0dPZRYaOchxTrKYOiK+oDtY4DRP+T+gFeuIqnfkfuGB8q3YaWDB56jk
lWrtPFHrA6hKt5WLrHy6oaXI7UpJUnEc3I5WEdnyJdGyzkYSTdmhcGAnouk+F6Hr
WTR/FYdnW/EQyAEz5v/+yR5xSeaykKaiwWX0YeDH55YXFGoU81dLwJDk3WhqAizR
bwAYojF930or4UrzSxMGDkPOQdzcSrDCoeCxT9CeaJKtOyma3MXJRv0PbT7r3/Uv
1vH9273UExFoVD72mpbYlFYrq09iC4YIV4goP/8l0vf0fM6VL4JGLmmAhKrFubr4
7Ons7eH249ByRfXbZkCGmECt/dYXzEoloNyE72qIMIUkrx6ROcMc7pUdiNm+Jedm
Dmn7gA5SvuahtqEN9WK5T0epFpME9trNvk6mMc4zDvFojcg2yBrGDq2TxLssbnR8
zJehkSCgh77MBEcrn/FqhKlEsfp3sPy0M+8k+RkN3TdueW2Mw/E9ZY8lr9SCkpc9
sBLFzE94EuWIjSvnMmwxzYPV1JKUa4fFpoPalYG2FmnPtw6l4OkuIvbVzS+w6sIN
IoesQshHRBK/cWcAiqgkgp2hnIpcOboS7GMYNzAzetBuLJX3CCjuzqVVwS9vVaOf
ouw7Iiuuhqrm572DqPcGMw+jHyEgEPab0Yz+jUhs9axAQ3iFB2CsAN1c9vHL4531
FVOR0LmkTfiD3TzaGgq8VMVPfKPdpr/YEWbisoQIi7R6n69s3NsAyxzqm2XpmCxD
PBNBNaD9cM7YyZyVxzfK1N0q79kPrC6C1jNymqzxRZhFagZM4LtLw9VMtCNpZynp
LvUQlc6rtVT/qW3OGblEtua+rYnLPF5q1dJW5TmSWqp74gwI1+Os+Gx6ary4JiIL
0NbgwkhwWgQvFOFaFBPzoFKaVj0vs07XrNF6DL/cIEwoh3L2NEeDOPYNcbrEZxuH
Hdnz9Z9ZCZUM23KD0ngvryWCgHe9J3678Y4ebAVomXwAyjWV4SzLd77IIKeVxD5d
Z1L44xZi+lMUabK02TSe9y7PCcnOTC1FD4b2t9XIQ86tMJP1UcwJskJNWlhcJSN5
8rEiRuLM1zqH4RZhaHRgRiNfteyUN3CapZYSI1nqEiFnOatrwiQyph15MWURrPD6
dVTrC9H635wC3FdY1G5/9FtFfzmQYXaIqI96YWlseTCV4a5RaE2lPfrQSTJd/L1f
4C3Uzp/IVf4ShvzMl5rPg3KzarSRooozdZmLnmf5NTzeFZ14PwRhT7EGHHp0AbuA
jNB4xlVSlUOS2VzK1C4bRiY4MyFZQZZCHxQD8h3uKw4b82JrYYxXT5nraWjtI4Xy
iFDnM0WOrlVtQ/WKW2R3v1JUS8m4aGUuDSFloA5DNBTunriPzm1j+VzI1EBlnCuQ
Rlro+UrMopUJ2z0q4IL5xa6GA8p4wlNr3HqVlGXQOb0mbEGt4mcYIuo4AriGZRkL
dOdge2vyzSwjXHwF+H2TKJtourhfc+MGUP+M6cIadLVddaQT122n8Nk4FIVrUXcB
PARMNPKO3qwv9h8f0ttAWuc2N6Btzbaj7RRt8B8p29hYQUvnxx74dd4sKS8QKG0l
6lyYr45OKIsqr7m7/8gKBjXXwdXOBzCcbCpd4MiX5iSMCFU2m29o0XmiBGTlIhR9
rleE6GOCd6HppsOnqIbHlxkmk5Bpp8DZtLqO6I2oMCdiEw6wTzVYiGH7UkzyAauX
OttOPWYB1I/sLoq7nXDA6QEqiKi8N2Unn5huxW33Xnpp05wcwBNQLn1BukHySAhs
rGNPIC1uBdU0/CAkA9EQ8D1Cr3FuZCBB86CqpC047oDRJ1ILCjnBe1rkzVTuKg/W
Cj2/IW3wHUKdY1YQVQctj15lzlZrXi5PE9uOziAp296IKb7j6DAxiFDidADJOv+8
JI9W6XfwNI/NGr3hKSTHxiH1ngvI4uZ3nqm/IbjMSS0s+H01QPgD1PE+PwAKtyvj
TjoFqEg2zQ6MIBpErsZ8TovwN5z3MT5T8ZQO3ERLNHTj7U/M3z1p0OtyXQmKBOUF
foj5CGs7giq9jQob+Mgj/9amrpz8dN0VX8gpcPF1qVJ8qd4gyYXWc7BEH1c8Xiho
pPGS+VPdA3piLwzGc90fb7U99nnKXXldIGJv8cGPb47K3X8cJf4ILaPX+Z5hxfXs
97w4cZD7QtxruAFK+XFUb1jZABNF0lfDNLtitFERXz6rN/iGCp4gGO8PgFq2+4eB
YMZ1f2Vke/TvV3cFRYnirqBgiXB6wsAR0l8VSh4JCXjPYPGgwZD00gE9ifedP586
QyYgyd7m4BVZCJBg41g4/It3UhSi/EgtBdXRSgRpNieeI8WBEYkoliSEEhpRPNJS
HungPBBoO30CWgbJK5ufq7e0cZH02u2MEIpN5Tuw32ax+nx9Uj05lfYz6qqUXGOB
uY5WTuqbX+z+ZDbCewMOAcTdjd2PVS7cIxT8/b/096X3GPU6Z3TAHCD0HBzdTt2j
gKACnVQpnLh63Auxy8UqtmG5cPxHBP4I3XXqGXfmjzTpdRh/CqzDuOJhM28Oq+8+
LNVg0MWTvMh3QNyPAZMHuxkzrk+62QSbjug/uQO5Y2TuS48EwXN7w3Ij1z03Y3tG
O3SG380geX3MlygVfp80rMNG0LKlg9UIhi49AuqXyUkz5wN9A7z+JLC/F0MlEEYF
PcmENmjS5v+uqUEGl2KASqftD9C/To/JueGbU4cVl17bvx6cJsriFjou/J7diPcM
vWUawhbBmvdUoiNzO8iCWwun1PSaH3aiK7OsJbH3RT/bVAiwcTVefPllXQ6w8pNo
2t9FL1ecrh/Coz5Fm/IX9WMKj7+l4HW07353lbcavI7usHDU4ORfhfzghhUS69P3
wcrwk7qZBWycviq8tM/CK7wvOhr27diC0dxAp8b+bBjTtNrzD10BZIfFiCyjOD7g
7DIZJa12G3VOFPste3TwhLW7BPhbHpIG4Gqw9aaV9zyYD7B5ygtwNmdDgQtpNJNa
C9kqZW56hQMNPhdc7ImE9TLlO7aqG0oCwswfCZ2rWGHjSX2fPxyhgfUNqp9pY58b
RCieV1V/EB75tDGaxBfHPoLU+mDMw86FgzKKaSPWd16NQ86COTixYbiZoGfSWgq5
L2aofjLuaxrT7dZs4p/df+5vABX1LEbDeyjjap6ROIZWZMH2Has6J62GUQ6wcoN6
8IdN+EmVCGnCMHOZnamTEEDsTKJ1uZbJZApxgPMSqVJz4Cw64JfQMttzxJrj3v4B
zSJ87dM3PmKYIw4asg3c4fLj7rEQdOUQ0zlM+sXCjem4c1T8prmMfV4C7KC9gqC7
C0d3IoMfKwna/sfcwoBtM2pnkFKp9jHXiYOZ1HMT7oCefYpEtrFDZh9N1ea2wx3d
PcmVGgvoN/Yqamng3jnoVh1ETKewP31AEdvELHap/9VfprLdw0cjCLHKPS1HH3cG
Q2vFIsd7f0uJ+UJEicyeiUdlWyytjFrlmwAwnQjrD+GPSICu/LGL/ExqauCkFOC+
rRTpuP09joMRKuHDjfaj3mbXJo3sL0v+S+FH4pKMy6W9ipmO8QfRwoJnW+8MrvjT
2hP7GE5T2GrJfyylaBAbrSBrEiCFLAw57M5cBHEfbvvOEscrpyATSkVrJ9fF2U6p
sZZs/okIwFF0JB8GE4I2WJcRNCQXIWwCsC4xkzoC5Dy5o/EhZOrISLl9ywaq097C
6bEuXdyk4bGjQ8ckey3bFzRtT8YwoICnqtnoE9BMj2Au3Cd7wijBMiHqJ4Bu77ue
hfxYoGDv70R58ozEP5pohVkZcUIH83PXvoqjMEhq4Y1ft9/wvVkL/5Y+8l2S4y7a
7Kn8Rz1iwtC51MNaYyKjFikDkigY7ZWtYwUMqha81uPBl8ZTu19+KtvT3QhlqdKn
qL51F70kiMl3PqVtU/X/k0FhxZZ2ABLfd4pRZnz4Cp3dp0PaDNA1WjnG95G8LkZO
EfQM8hJYzHsNRIfaUuFpHMwq6gMuz9RWGXU3LsFdIQe15INI5/hFIeI9EqdeIc1/
nKKbEUzP2J8aP1A1pSG0YM/n+cmr1cdkRb2LMMNa++8UPlYg2H4K30QzgiSIVXWL
hR9N6P2A1G5dX+I5dY1B1XZCQ1F4qLoRBM3xa5YD4d08flSX6uQMhJmr36tuyUag
1bQIUoXXy5NTVy+zyS3YiIRuGJ+9j0SOP37qCx1nj3pzHeGRPC2L3PFI+uNRZL2a
Ql3M1gjH92tfJPFvmmpjLxqMUIaIJcMk0zuBOFwu1Dagzr/a9u37aJIJv6aDfqc0
3/Knh5YnniwM5fP/CagL7BKDIqSsmB+x2WyyU2zUzykRZq3ggZMgwDSWRge3It+X
V9d8Kh5RIBvbYmKWSUnv9VFDfIyIYoPB5NwSAl9XqKFwVgha5QobTLR4q6u4sIZ7
wmQvbJbTgMXQ9BLvsm4UdUvjw4l4rv8eJrQgd2/LEbSM/5czYy+zBVje7cwmelnv
wXoK4nbkRuUeJtNY2g/KpnrW0Y0PE6SWkHFJ03C9/j+ApMrmzvv8DqaWl9cOH5GV
SqlOU7uMITd9ntp5tthpLtNz/MitKTRzeH5v/PkVArMF0uo75T3NyHT+vGSn+Pi4
FVx1vVdOUe+L1p8EHDx1SmM6xkqklTzZ4DB24A36JEIZ3/UdujxeV8L2LZLES2VT
HNM79owlVTM0dAt7u3wE4XgxsUOICV2MUYqpF8LaSzgzqUfhGoJVGs0tq7tdXRGg
HFVnpyhHxQf0i65RrWm4ebWDMZhxiwAQ6xFUix7HN57UrSnPztRYIef6BT8jMKxp
LNlleE0NiZTy5BBxluEw177tMabEUcLyKMdbhGhgtprqIJeuB+Hk6CUwzAjWp/Zo
gjpC6cW9zEJ4ZaEPyyeZQhxXrZZpVl/PpEZuA2srr3oyjpIx8ZyfSAbizcQ/yEEx
/YG9Lpc0jl7a6k/thO9eOh04BzLrjkE/RQqbv7Bp26DxwUpcpsIhdw7DOE/LuezC
SA57eY0FcC2siZhYpxKFFm9tSgtqwB7fd0OluBnAQJZFL8VdXfdOIxsfjadH3vXO
EeUinqS6RWddBhIIcHWCQ6m0F3JOc1t6Sew9DnR+2+Al7VOmk97QpZYBA1G2G/wL
w3hpNAsiZeXVUwJfEgYDg5SqHfdPNSSttTQIQkmCeyYn86ZXuJLbHN8NMecsONYE
3ESLXh3Ddrs/81A6PG2V11XZ/3k9c7Z8kUP5SRLX3/pjp0ZBZjWlAN89LBqsmbUq
h+O+vxPiujtn73E+rW6dGk+6DFVkBZeSQJgZtpucs4w+dG3fWcPqIj7Nieh8Xcif
EMCoNoxkCJNA3d0qdP6i+NJzEgQ4HyxPwRxlueGU/l1GbGPVImMKbpvaoTvsj0MC
dy0q8R8eVIs8oQhD2oTvlDnex4Wg1z4lVDdj2HYcwkanum69ylfXRem8HGDDiks3
41ZQMrI1IuQ50SLyokQfv4AhLoyoCAfUaLPmvbGKXRU5RxNCJH/gr8x1Qz8Xe+c1
bleno1bIqU3ejPYh/vsoFJSlmrIao7sSHFfb+GcZORL/QVe9L5edMUPghQZ56YvQ
2F4M4P2cYfGthZ657fck1/dEvCHnCNfC8f0SdFMl/aNB4j7JkZZfghHPQ04Nwx9R
ScIt5XJXox6uUKg+10onivI6kAIF7PJOTwesaNF94WvcM/LxHhSYWgVNpRs4ks7D
TMG5nY6UPStwV/yAdBwuLQEwYIo2sOt/rQqGHYkgjcK7rOvV6lv3jNLXE5ZReqnH
Og4IHi9/y0zIzuYH+3Jh7rrDAyw6lIL96hX61ozgw+3iiHWoF2m++eFb6g4ctSFx
6B2f60rKaXCVV1qVZ5ZZ5wr28DAbAvGRAj5kXL9nYvunxYGybdsfYQ2u8skMYBVD
rjOvQSNt57C3I6MjXqrTd3fao+uc3sXQWj0SO/KhEcWisyvxolgwZx5i8NWUnKa9
qiUSJgPBkSXkoJzpLJmfEcQNY+EMOX/vYiY8ByA+29C247SU0zxTtpUH441Ja3wq
XhKvBh5tXr1TXlzVHwGHUlWLn+mV8PVatEDG96vji3KbmI8gkpiXNfga/OqXjWTG
CB1C8Ivc+GgjQzWlMeE54Xcqbwk4uMl0h1y3m3/Ec8T/Pf/rwK6Np9+dlnZ+o/vX
HNFAupA9CcutAxp4jqhJ40YOwfrOyhXH7rdm0R6qgZjGItkc8nmTpsYZItbJ8vI3
VDMzkbfPGIIq0LXmnn8Cck1MLJNFJ07wakZ+zMDNhrSpxcVwEuRZ8x6aSo4jAsHH
AEzNZ1NSNw4COQwJMVsjB8XgY2gGCXuwK82c/pyEl1V5EReIZL9S6dwpbQYtiDcz
6PgHd6zAOvcL5wJ4MCku/X3HkFD4H1KA2U29ubo09k7McUmxBoU5QBiIi0Q46Olk
I51C9dl6DdJMc7AbCedk7IolJbuK9+xa3ZGNg4OvNvrTau0vg42FCMr2/kwam6bz
Q6TWRwoAkPYbQfXQaeh8wT0sOicTl9xI/6fPGjTVX0NpN9Eif2jQg/iWQpbCT/P4
L+lptxbDhebldD71s//4xM0Hte45h6jIaQzTHVUgqlpqd4bifQ8/DCoblnvzEwVT
80HDpypQomtmraxQr+jOLkChWYb31ATVi7yzj+/d4GvDJYtgDC8OLQnGWSnJsRg1
8I9pmuAqIAxvQjVocCpycY2oyCl4HARQz5Fh1B+mlrCgmoaDnJbCmfVGloyFamDE
9YfbQXZeBCL8fsDu+NltiyIQBpQDLt+FOqdXunsNL6i+l9rjQWYWS35MY5iHugDq
5Xw2vSk4mHyZMnB2D3BuXivIZmK/q2mmp1uU54z5CZQbPmJHU+0wtCwOanFISLxM
Qyj8whGXF/EYIRmz6PlDbk4h2xZmt7N7bC/Y1c5kaQWllWEkKnUm5MZo8CYX8KUl
PQ9OcxyN3SGeQr7SIqb/WpJ4/9LoTsyRyZ57GsB1tzHRlknfRkc/JQdziWWOOizN
6M8ITiAKbx/Z8z8rQbXoDtOuDgAQCXlwtX7BNJUALDAh8+G7Q7COiqJgfhi0ksvM
nK+jUMeUdAl7skjQphYxeEMH2B/gfLxEuSlvyMTqqghvS4fVP0rMi/EGOkOXsYZR
/eWJX/FkBuKBk5g9EwxNkRenK8av5UbgSJ0FdaRF07VpUxey/uCdYIeZYaXz4MnG
WoKezsWoxTExgkTiJ3aTB5ZjXRHuhivjXEVdbhCd90c+vNcfvgfSpxOaCmU6IO7x
8lJXESsL8Y4hoKTO6cPs63wTaPmFUZVsbZ42W7Wz2Ug6vK7GYaub4FFf1lgQkzKu
ezgvPrmfmM6vCoetOunaLAQZHSZZMuwJV15/Lf95mEIzvu7G1sl6yGp5tb+hcElN
RYeqtTJr2L2RO8GARsaJ1wzm3M9jMNniAzuhG8VQLLQnAP2WyfOij55nCPKyIKLf
t7nMO1wQt3BIrophghdjtTQGMcohAUiy3U5ZsCuypoYGPQeTZsGD9YWRLVlnXHvl
ROnLI/7Hnzl2PKuRwYblq1jenOZb7cHlZBhQzq/Jta2zORry3MBUVUNYYHsw8qya
9iaO/vW1r2uh0OqWhtYwwUmXptGnSlhV5O6blygsnaj5CQDYDkLqRMv53c+5XDvo
GFHJs0Y7REwy535dMi3K3FRtMY7s3ixgyYu7u8AxyL5H3/FumMlSI+wUBDN8Gx3Y
zCsgn+zJOOxQMZ4AwTDz1ay+x05xyEdMX+DNOKQY1IgJBfWH1pLtUVcGqUG/NOAt
c/S/w55yLTmrmsQQsQhhBh8uoU6xLSqxZxPjG1//wtbyYtJCY6FvOcQTDGh3SBOI
Qa6ZIU/YY6BSrBZUt5tNCPcUhLbp2lJ7zAEo4HDEBRfbmo6SN3ADN9TvhM0NN95J
KlqMe9ZVHfM1105gSBgyOGqKu8DH6BNz+Jn5Hn4ILeXPS48HhcgZTjyAUrSxai0D
xgU2cvaOWAkKwEZmgiW/Cqw+TqHCuqQOzzHO1YTOwkU2C3+EsQtzGfU2PvZxrNiP
oI1m6ZQL3rKy8s0OnYgGRQX/taWCIFhdQELAdGwbZ4XrWkc6F8xdktcrlluV1TVN
aXSSohwWQrzvhw2JBHl+oJhC6U+rkHK7AoB8PzJvkGauqcAFoyZLVcmHUtK9iZ56
2Yxae9Tb74Ux3A/bPX43VA02xZsbvjWoLusFPHa6/C5r3jmPDKI7a6uULeS71QTS
HvUxcHYOaL/PbJWu6aPbga8jyWDT/ye14NZLLJ4eHLpzvxWMNc7IHJ/X1eyBJND7
GGTsYXWDUntFPs1Q+lXwOLfyod+7TP+m3SRY5AFi/9+1LAsRgUHeYfICRzO2+1i5
+w/y383GImwFXekFw78wtLRR0CDNKa3Itj8PLLSR1MXMe1FQ5mDOaxWJzFLl5ost
JAS04Mqub/lHVAW4EA4e9DH0Y67iUWje0pKrUeDAYE35FAjVvhm9G3l5Yrivi2hx
YY973TIxrB/mIaUbDbJaQWNuA8l2+1Y5i0kKABYKoMYuJbJcDQ2uY139YrOggT4X
9XQLkm2LqcxKSWfGSU7QlpWJsLEFqk/ISMJ5GyBSaeFQCEPV3WVUfsS/5X0RqEYh
UCfd7ul1mi47HszPVQOJrMOJEKdc02fH7LoWEZBckGtIC6IkmC5vVWWSMeniHX3x
IgjZMZSBmAaStgUkEgx1JPYQCMdYaTlJ66qbQsvJa58f6ddFndLV04FWzp8kWtqh
EwetuVIcp+s+smwAdi+E40tJKSvPfAoEDhr4SiEF3Pv1XSb/575wsQln+jfdhAwN
A61SXnCT3AKZYvDzDJ7fQ92dWUAicu54brw4figg2c6/Z3PcPSVvR6qWkg6MoyDF
SYv3nb3AQRjp4l+/WXzOVG9zf/baQeszxfUcmHVM1O/YPpbAytOxjEHZlF4kAOdb
3nWNZ928Bdy1ETOvL7Q4+lkUV5N98QKCRUFXjQXTVu0vOXu9nqE9wdgwGtByLts7
sY6qNVEDSbfX4Pz9BiiCp/nnFTG4adNXCHaWhNk1jbdFiegOebc04Es18Mx7K+ah
GnB26JXuwlulQopiAaR0AEiGISTEFN0J2D5KDViCGbQMp9s1cBd8BexSU81mOX7E
GbV4fJzaNftc8Guvp0r6fSH2KRXINU2mZoTcN+6eigAHSL+q2EFSEprtm7Gavlgt
CCvte04+NGFPXQhvXCj2qOgX7kR/CFpbCaphI+eciTDdhzCen8lSuwynw+585o8I
u/NbofnQeIBE7E0o/9JNO3xsMwO4spdFYj7ZfrCxi4F62KglsvaZhO8LsYl8+ilV
vmtiPnn4yPNRJTytYkPF9EgsHyRCepbNHFMebsJawFTJ9fkqmklbvSV4lPA5Pz6E
9+FM8EpYYRN3KxVM5vhyyjv9QmBA5QFuRm0FcSq8JmmplZwA3OwHgXaVyK105ATq
ojGTqQ4aPVL83A6ePfwPo9FBbMJgvyb+O7YQCEMipcisccFtlPcez417F6EE7trt
SrLIryIUhr9Akx7h7hzUc7hvBeY8Ms5Bx3lMZo5dP73S77Z2S2C8L2s3Og0Gyz4X
hGYypHbIQ3AhP2I0TeF5DT6+I0gz486yQwtPUOdW6Tt4jsrCQ35GtRq2go+b2qMs
UmSzAXPZqEmfuSsnkpXbh3ZxXpFd5pD8YegP4LqMJXnuMlUjHwgtL0F52Z2kvHDR
C1/FWBxS6MxO8s9GR05JKeRASIzNan8x526xr3djpGYZZhCwb+JPIdU48d7t1Mxv
ntQXcTWFXz+MG35up5tUDe9LcM7/wFBtFQGAsCdaG2dgDnBTlvzAbHDhOtFMCMwX
0M7dpqveZGiMSjdarv99D0ehu7bjKiaE6fPB1mCWvq6UOU/gJ4qsoRvQCY28IpPY
U/e92sgnWa7l9vJbg5G0K6830sdB0doXgnn31byB6VVy5euehXBhb2id3OsAPwRx
RaZtO/bCtna15h/Ux8/DhfUSvTsaD8yK3DI8CEhU0cOEY/TbBbDMT6t8Psk3Ohy4
7VKtLt5l2pkqtK9U5Ht0DMQPzfAcQNVDhLB4FWCWE0MGVKAqrnn8gRV/lM4VU1tz
1hfUmcK2z4GgT5j2adjwgGGU8uheNpkKa6sPPPHHyaOQE0/N2Jyg1kvZ/hgvb24D
LvA55VdekLjadY4JdUQ5mfH8OUs4r/Ig+FUVd/J+mzqGvFjVktBdcEf7/VqsRyI7
JrMxz6HnalOla9nMa1bG55MRgFJuL+URc3Bsm1TUbUKDo2au6Bu68wcMG+4rEfGH
DBtSODUWWJ0HccAdnhh0kz1gJnU//S/4QBaWwjtqd1bTXsI2JVnd9I3VOL8tS0Ni
1f0xL5LxxRJFlzAvqEzi4B2MTw2/iD6UF/PmLt3nRon8V44B2wRY8XnVmGa4e6qn
RluzIzuklPkmpI7KyLnes8qGpt29okYRPPbtwLc3tKXi9EClVeB0t0T9GP/EcWU9
UW1Sv+290dbQnsbFS+mUF3ckvPVIbBG+GzqutZRT4fCszy7yq3RRr79d8vM4JJc9
p/4osYIIdiA4vumG+8dXYampFrnVIHPnizuktToROuksN95gKpBjd8x+LYisn+72
toyBk/gh/a+urv8aN4qUxO7Ei7qRBqi69nMrHr/1VtjJ8P/tUawEK9Fgtp6FfRca
VGhi25gbpnQxi40bJGIPi4b49crUHZjpebhA5lH8m/Ff4twrTNuILVrYIImnARTP
xMHScsyIU/g7mLlL/v4cnzNxN1PCwdkpnMglSAap/mTcVCF0BcLQXDCFEHFG23DR
gnseBcWDc0WQ7Qs7ZGcy0RHUkgal4+gTjJ6KWxXek0ZIHmd6kZRLHD3zHOx60r6G
F3OBAVRMVD02B4lJkv2zxPyc6X7Yubo6ZwA3WlpuwLiscd4ztWB6sCGAsmma+q9r
ZJENK4+6+j7KWTRHcow0hIiWBXpihwFP89YfiLWDC+DUvLNeSF7NT/rgPvhntVhg
woEvHxNFpquRDN2d4cnr9qjcHZMISVmcdfiNNy35WBOELhW8gV08U0mOm49oiArn
vcdqnKfM6mT9SqkJw4b2vkyM2vEtqdmnEL6LVIB7g5Z1H4Vlzzjg6xDMW5JS7/TT
VdWAULXs7+Q4pDMmNrcFQzjJZd4koPf5LgVXa/EK4bcHZPV+dMrk1hBbJ4Ef8xEC
K6jZSkWiUPtnrbGqZ9/7DWgvmw5r4XFQ8TvJy21dKmebxBkOMoXn+IDu/0H7bAE6
ct5PZslHKthbYoW7ke6Drh518I4Wt8nUj3emVz/rsug4k2KwBmqJTAyruImVTDDK
lcyzYboqeSNhKkfjLq/4ibI5zMCZ9bWtc8B1S18rYd3uz+TlyXo1CBmrjGYyhgyU
Wund/rHhMx7YGr+JldqMpG/7PLmAjUtfAoJj4CXLL2VCcojmWA6TZENMWPKG7zt9
SwevuAHxuQVYyo8zaUA5h29w35HVvqypzSNayfZXq/mtcN7rRG1EototaLBqcRPp
AtQkEdRvElagtyX118t1lkwyWVYE2iziM/Bai/I6ecm9VQMlonBnjiHLNWXVArI+
XCWsklB2ZWBqNTVhG62bTZ/ILIz2RKTqlVHDL6yPne1Xk16JNvhwQjUpu2oqVwvt
B+AyuIrwyHPZnVZlu4vlt6IuhZMGIxn9svTY0yWd0r3HJq4q3UkPs4/DVsH34VAz
iuoq5+u8Mv4Wyx6bV5ePJOl7aq42OG+iJiph2p7TGxi883rSES/BftwQn8QhE790
V8jOC3bmNDiSf9LqXCJKu7jpi0WjxLiKGIC7YxFtWBp8W36poI4ezDVrHyL8gHG6
UDYRuazsmjClCkIbGJ/Iaq+MvWEsXO1N6W89Zw85Leq/9e5HkiY+XRkU3bEBS45z
G/mQodnmqPlND8i46sQP44Abcw8PwFqk47DI2bY0uhiwcYdG6Y249+OeJSbYgwwK
S/tFzvujxZDObH0c+I8PMzhypcea5cxUe68T1moYVBx2/FLzqAN4MqcFCxunKXW2
WLVSmgpM5BNTr3XUhtuzkGP1IC+o0AghE+QUn90oA/TBqzTO95yXw+kyhCaC2me4
TrnR82d306oL0uYPsc3fpsyS16vKLRIxyzJfz67ECvjc4Ib3dlfr+O27ho2eJSTo
Y3pjqYAROZqTg+gRE2hw0po4cjIhm2PoUIz9Y6FNASjx4VueuBzXC0qKOYh6z24O
S8PCN7bWS1HEKC6ALqCJfeByGppqkqaQyXLXUfNnUNGPi7PUPxoM1U7/PheeRbmd
bnctuPgPn3zN1TeZz2EOZD/a4VO47bAIROrpzGDDT3lFiTo0l1bnBd3SLwQ/B+uT
MW78Y4ifa6y6ZNfDCAU2kZ2k1kwFaEg1Sv4BUMbzHJ9EKKqFNC0CLskAKR49Ux5B
ZtRnW7tVd42tsP2nB0nvEkUT5ohdJFhQFIgRCwCgYFurncPuhJU3gjYTwVQ8bhin
YEvdqt4dNE9ENLIf/BWuv3iTRCL0n9Vn7osPCJfsxqNzdyYnANVHJICAv0q5rzU3
Fx4HuePd95ZxCMUM6nxW6TcZVTvNnT6OZ3lxv5yUcjD+8ZROXTJDjatyQbwsjn7R
GWzJa3ziXtjLCkeVcf6jFEt2i/tKZd5FndOW0wZ3PHXKRjXXr9BFOEe8vgQs8JpF
nykz8ZNx/vgZTbOsF5OjsjvXt5xi9C0ZM9YVv926OVQgIQdRQKXnyJmTn+I5XCfe
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
iHsAQ4c+Yc03praDkDn9CGEbxBOpVq5eLOgjQidG5S7vYlxIZ3CdaxZVYJ3LAEPT
sqbi9duOYCZANd6nHycjv4x0FEZ63BATC07E+oo4trBs31kNPyCeoOIPRA/+EK3J
LtvGRiJ6LVV2pmmhDLN0W956BGsv4xjy1DzdI7v1qK8EjbyU6WlEfZaNP9ClXyIY
z/6ScAk9J53yBusySmWXMenf6S9eBYSHfn4D2H6RpgPtI6F7FtKxhQNekZYJdD1r
UVbv3uQdwkGkVE+BdPoheQb09V0OAKIbyWuawbBBuUk5xQLgzO7mdNrLqS4UnC0r
PXj6ESHmPjRCWWNFQAdreA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4528 )
`pragma protect data_block
+aXtq4yNq4crE9hzz3uG+Kh6BNG5t8LUqz1ZF0YqewqjaMnCgU9CzE6x96abrjb0
2XwEuG33Qff5OHb3vDjFvQ5oQcgkhNX2X1yyIwyoL5Qpi4AUGjqsDKNcrcfnt/+r
jgvkoumyKeN9PDnxnDFxIFbecctBvmILaIwk8dmXsxkOFYSeRwM3tCRMzYRL/TEq
A/QDwMOpEpR/ieuS8cM5zplEnW53dLdwiuq9g9J5DX+k900gzHaxT2GGwGA+gKKk
BQ/SceOyQST+BkgH26r5GP4hHgezUf3XSlTuBpc+ITLH79FpPXzxVYdiqOYYcOip
P0YhxfQnoT1imZ0dnEdrJ8YSi+qeMVCVDmeXbdK0TRHgImbh7cVJ3etd51RSfINP
jTE3l36cobbOu3hi4YiNq2vP0P+cApirJFCEKCTOjZ5PDrdkSAKPE9m11h3z2q67
ZAr0bLTFbRvIAIBMudMuoaRDVSnpz0hGLF11CBziTzRI3j2YNhqKT2UP2yUpi0bt
IzKo/Oj81qQq+/Bw0LXxJz2I+8ZDjZK/yednAZGs8tVBlhrcjoXYczi1EwmaZg/4
oTYxmBJJxgZ7Iv0TumEpxPkYIv5xBIZ06Cx+vd5lWOkZcAczbv5Yj6qAf2qkOdcn
+VgoL48xPJE5Zrt2x1z5TFbaKKLfwoKQTrBOigmz8w4BsbcJsx3WGY8HlnXtBmtA
l7NA/gohHkCxDrdITOV/DYXZ7VzT30akfRA0Jg/dtP2HYQn218ePAAMxXGZOTOz8
NyXpyTfFNANW3AF5b1EH0ZkV+hBmDcLhS+TrpmRYYzd1jS7c8VMXou6HIGuQsFvK
hHqdIgRY113uP1D3Od42LN2IPsMzEfPGPobLKoEUEXQeLAugSDIbvThYSg6WlplB
3cJXFCYC+VExNru2InkD+8H3RAAUqa0VLXvwdDG3rbOhBMmU9T9DiYPIUSzGcx93
sBi/5GQ2Z48hrbAbUUg5OcuuZxosPN3Mk3izO9vFJDdOcIuUPkjj86m8NJjMS15g
O20xHFAilh9jkbXq/QfXfou96FvJfHk3+c79NsSYZw7TNtBo7LBLc89xIwi/riSS
kMPHys/Ieu9xNQIHSED+KiDPjjJlsPkYn3hJ8+AvTmuSdJxNxg6h4yiNXpwhBFme
MSThZR+YZi8uvF+4v/gSBv2TCBlUhhbBmxytZe0UlF5YK4X53Y7nJ2eYlChIfazy
+AzFO9PFqh7B5VJ+fAJUzGBGRtqUuKphA8yRh+6qcCdIaLjcY/bQQ1YZ9RDWJagF
PMV1pp5Mpdw1e++RP7dM1Wjl1QIGLCU3XvivhKYWtjoKrwcFPKN2J4NUAnCqlqa2
5axjg430ZQ97mn/JdZ+MewYxrtb58tsU8/yJki/5oxmpVBN2EL+CmLmtmF6CTe7/
PbEyESweFJ+UC6aSBVbAJtuiaCUgT1Yim1dZ4UtSIm28BRsZQ1Gq2t9oWcS7ZiPu
QZUnP2OBH01Hh86jnefJijzHIkmhVxFKDbVImWpJw+sgebA4bRPRD0PO6NJA2nj0
Y4ulmCGbEDoPIf4i/S7TMn4Oxg8Og3kwN+4d0O/8+J3jp6mfmALRRGXSGmn8OHQW
Yb5WvdozPFLCetYzQthhEbWm8tJClKcP/CTNl/QLDueFOkeceQNAAgQkRCXjAMNy
zIc4M48vUitcrrs+Jt1s1CcnlwPvSiAGCL1f1NCaeA3mGtDbsUSTi2JmJZsUcQQo
Ylz6LaP7GKavEnGkSGD8hSHiHVfMEbgIvyH1CzvMKNmXG2XDx4lI33tTRoiIrQb3
8kemfZ/wBObUF9NmF7L0pH8ZD9uBfyJSaLJUDqNhNvPKccE/QBK6Irr0Bu7QrxV/
7CrdXQMu9iMa9vygCvY2GEWWCxzzY+i9fjopE+KMTFefp4Eo7rrYh1I4KcLO65HZ
TKanoO3eulfbCAC1Yh2NkZAU588KVgEgq0rWmqdLW99LFhKqs1OpD/1GPu5Uzllh
vOJSpRHTYJOUuor7gsXEPjKYtHSXfZ6IjGkY7FRqortl8LqYn4u37pn2MW6u0KxH
37RXOeyY4AonHyHYr/qSkxiE+qh/fl0QNi91Xel880eTpqsojBHxKJvDUvIwGAQp
QBBXreUT5MtxAwyK6oJGlNev1WRPoGHAy4UX7KSPfnUpnrKS0nt9HN5DiRrOWHJK
FAmKYccDbt4WLRQOMyxFJKp5xxu3+/s/5IJcLeSWSLmyZw78ju9H5PLwVRhFNmKF
C3VKFfTx8TvctXW7NUJLglkPx9UouONU8a6nwnFkz8vt28Yy4RHoiWhTSbiXpys0
/BFBDHJXisaHTHFDiZdhmU4W1Fg2Wi7fLDlPZDsAJp47BLXBtOuFWy9YqtDeXJ2p
m0o0fZpFs8LoY1pk2knOH6HHsgCOcqSKP2nk/p1RXysQOSE8LEcItpSvn6P3Y8q2
dtiSagoZJrEt13KOyZDMEz6ilqqTm0nq8M8x3XA1GduCgYVVxNlbooYiDOEvxsTo
0dVmVmwnERdECVuz76dTaptHbKSuU1OHdcihZGeD+/jnJUDuqdssukJrxHcIJwxP
J5Z9gq1UYG5L+do/Z8jx9T58KoCY4bmPsAbtycpU2C4v5Nro/LsY1xeDUN3mBDHD
uHbA9ssP+tdSfSrpPhozS72hsI0ph3udPBR0v7gYIFGOgGh/1IHXzpY8NFHSRGQE
ubt7DKgY6+wIym6nfOi4ZunhdIMMLAdoP4PC04YErTJLnntk9lbnV7lMCpdpi9tb
XAwIApLK0EjJsAqpGKEs2ErIMrSjXjQ5yJnMpvfoWHdHi5/F4ZuXvs3+SwCFF7fS
jOSDkAHD2ISa6aMi/LlDi4sHOmaIP4Ns1XN6i3Q7Z3CgH2Z2v271JUy9Ft+3LvJA
jHUmWefqgEHgAbB0imRFld4nfBKBih2pSsa4JcPjIDAVTvlkUKADfRC7nW+EqH7X
iFnooDXMp57G7YQM2tMzWXHb4p07Kbq6AG9fEwYvcV14pjtSLD8CQ7/18l9elL4r
refBKREHfGS6wTDRPrWQq5ylcYgbRa94S8rxvBJsdjCjU9EHjJASlWECOC6ZcKHM
QW47FW0blFcLiX/yzpWBZVJe7/kbMTJ0Li3aemTKZ31GaURPWpONpdG0twCcbsjv
o9QYNmxi9v8ymP4Mex1bnog1poSIXXd56lY1F/9JMuQsWjC6N9DuD9gMXiQ4VXQb
0GFG/ogeLNfNOHNJ3/p9Z400n723uBOt/18L6l872gI9o+WNIAxFMInTBEvmQf1a
2tkL658//9SHBXzGMxdgEupA5ybAJg1B3Oe3FOpiW8I8MxVfg+h8eyHaAGxyOK9U
SeKW8NBu00zOqctQAuB6kEredlbs46VHfH6+x/OQoKB6GGWFeRvV3IRdBrMWlD45
QpGtEg/V0lxC82qg2J6fEIseAeDhATwCtycBTINOV2G2nra3Ya1DCqvpe2/mwK2I
811N3uinyXNr6b9Hpl3U4IfLYqSeP+e6t3ia+9WlQqPHteDG7h0mCQA6JRTKkC2N
+Qu8Si6RUiwsQ7vwQNQEuS/Dn0MefCgyyq+ZQqWxgPfdzf1Yjm/8bisbFwoUn1A6
nEaABkNJQ1JNeL7Aa9lg57MFUHK9ikBwZ+d1eXDgOg5jHqB11bL+za0GAfc2Y30d
qGXnXz5QKxOvU34Q7XeZIEKdNfdo36L3LxH8AJ17xaZxkF12dMoxZmB8RZT3j9T5
DZQa7qmiMVPccqwhG52WoJnkY1/CKxpG1IwnaUwQY41tBBmkxqhugv2vbxQSmtwf
ouWZhhUio5gmTFFHxrIuYZRf0nOMyTj9BM9POo2Q2ygVzcUSnZJiZizoZRViHwa8
NrQUsSTlC4s/8Ziro1dOLvBmQY5c52VyokMHEeFgNRS9B0/S8balqIDkXUOmZDxm
kjNAGY+C0M5Ephla2/HBT8STvpSwatoVj5Z58BiJXxuTvzQh+toJ1en/kCoaLsaw
y7XUaH9HAayROpa1Ll6QvqCiOEAvEgzu8n51MMfn646lQFjsYakz6Fq2Vc5TsifR
m8Z8BuDLrbwj01ne1kRcplKa8EOXrYMDLwzX4SJortV4JA0DLklVopDSdOfzxiMw
Q/7/lvtlDGX4G8QpnUibINqmALBzF99/RZeCjIWwJpbhJFLIBhvnZDzaASy7ki+d
ebnzozAL0s/du4WIKWqiD0F/Cze7Q+K8VCwDbgm7bcDlk0IuSQyquwitvMPsAgRY
lv8ziHgNPdFjnN99UQlRrI4y0k6ArxNXVncNpN1555iEP4KDrh8jqxgoU0vev6vA
00zf5NYCIUycpfk2GyzsDKB+jWXHiCI2ntjnW/4MeP1LM5BRHxAxvSqaDrsaCPIC
SIP11EvNnNl+XqENJMsJIo3Hszoz5DDsUbBoWEXw2f7K1psyjMcAt4pkq8YkslqV
NoN0o5vLV41hq/C0RntEkJT7DFCN1P8oLgl+ogZBbUSe05n1keMPQFYcEeeVOhnm
2FV/DnKM4k2qxKgvN72LBZdVj1bTQI9oEI6iZraMKIqg8IadG72QMu5Gqj3/Ib77
i+9s71D1ijCeYeUujTSIyVdPIw9jfgOyF9gnkCZK+4AnnNx38URzZsb233fd0Atl
nVTebHkRGgikh/Hpjh5NPBdwVRkvWo581MhBHjR53ueOMnJTeeajvC7POYwkJjsD
26rYsBRawGD6KZ0T9+P2WoCJqCrzxn+l9qht3onzeCL0o1jXyZZ1Ozhz//nVqRJw
pRy7tjbn23lOrqou69tf+Wl6IuHhq7InGBeG9UTxsDurinAXpBJLRQB7yM1Emg85
aIQENL4jWJf7P8JRA+CH5cJXGIw27MsKFiQAVeJ5MAOCN/sAKpZtuWdgZDTIpxYL
2bm0mFLEZmiRhUPtj/nFH5qqYjgevYt1jEXwzJZYfb5muiRY7sMJMmaHkDd09fdP
tX6h8feAVMlQJVyNfUNYL78DCSlJp0gMUGuQYT1Qv2tcVsAFgkRhp7gzmF8UCEsp
t/ROFE72HlNotkfsD3R1s2nBRkHQNiMoGOan4mIZHt8uSeD022ymVLgAGrWMRhAW
bJEOXaYXTuQLF7gNxNif1hbySLgfTyZ9lWnhHb7aMApfBTlp2ei/2uFjQBhZ/x+6
3Zf7voClWiHQJmNJtI2A3ihJ3mE0Rkc0jDKIZO+eaRWsYFNJ4OUsjBjjZfL4ABKI
W9ox1agUrxQ75dtNuPF233XbdRTlNTQ3XzUxUB52aGKtL3+GcIRWtfA9pQIeHToo
s2QwbUf2s6cYZYMMIUzDFS23KTBwOxNMLMxpr0BNHQZ/RZtJHa2jXpCxb3vHzZ+6
WYOylmWxNIdEYcE9bIR7BVBSN0jNeczRB2l1lx0FLABP/SrWgjp+KlZHdBp/XX0k
gda2WB6uPOyh4UEFaDHJRpap7JIhN87OSiab09yAy42JxTKA2NHvTovhbfhoeGMD
SnPNt7+kQu9jSLxOUDZ1ZIjcCQkmWZ8aC1YXBK0Tb6HEFz8A54RwG8pArUN/tRQv
GEZAwyaRd/rMwNlH5zRbaZlOdrXEFSCNBs2Aa+nJPfv1vgc3g2NIvuNJV5KdjThG
lqLUF3hRQE/6uSCCPayvCeatskwDfNTS1LdWtVqjPPwjRfP+p0N2gbmdHc24ncML
FdsKI/tNedZz77A0Co1lI10jB8yRcjz2s3rqJupmZ7sYFu9UU60NYdl5vw7pkkNu
MQvq2Pja7UwVQ0yRC8pfN2ukiGA0jKsPvZVA/6SnDszfZozELwUvbu4vLCHRY9er
SWxUvP//5sUvh+sOgGSBJWWUCK+9RSH3dPWxNvlYUHljU7D20Rp/qG7SS33OFBXK
AEmJCggdWBbT8Mrcrnq/kI0KPZz6BCuzLqG84LTCtMqB3Av0hC2RgfRi9Gi/EBQT
Sj9OE73rQ2ouIcrPVvlIQVH/xyNweLcTymApfmF6ZATY/H4w8jjrZTKxdeh7l1vy
ozBNOfPOEAOmkeD4wS7FlR+vQewJrak5OuC1qQ6SFrllx+Ji0oATfw/34kVBrM+N
+UqCiCmOri0GcAhM4gAhgg==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
I7BhjIYbBBYfqlqrsp7PnFfEczQRKJVkDBZoaZ7yrphAxlZg76VBSlOwbS0PDKAI
zvMmuOx3vQnoDGCEo0PHWAKjIMTFiZgV/+mTe99Nn528e7ufT+p4v8EWiWQm9XJC
09GGZTQh6elFuo+XmCpGcjuuvgSxMdIkgYFu/cnWcI5Jyq+mY71NilQ5ey8DKU78
DX0Qki5xisgpd3hjM9HcmsyjWsuIyonvOoStc72u3F4MBf8q7odYgVjf8hND9nbi
qHIb+qJwOX9GaBMOMxGXTp0dRXLuNGlCqGwOwRiPL/duXanUqisbsw3UZ7yEtkT6
qgGr+NaOfCTV0nQUfH8b5w==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9584 )
`pragma protect data_block
9fCv9KvTA0jsaaeCBlfu4jxvK6gpF3BXxPCbJod+TcS1AsoxuPK7FrfHkXoOuVyG
kZgJz5OqooNn7COe7fCvWA4CZPLTt9oN5z/viWjqmN5PBhIm1xL0UYg3xhKjg1jx
LYvmSBfIguK+qfvXCPIwO+Uf41LTaRU4l0a6oCA/f5EZMMan6MXnayFwQ15x2W4J
RhT2YShq504ueSbCH6NRGUlsyi9/3ORTDcBy5NEZl3ffCbLgeTCUjlLlVeczVOia
+wEVuC8NuExsqUOcZTYM6MTMNUsYkYTLzwPYgLSX9S+kNqcGK+QUiFbMXkb/DAxY
iDvL0qhM9NAL6qpnSwHSr+3EQGyb/6NKgyfd0KmEWbL8ytRjwSAx9PK59vS3cm9b
sUU7AkPkwzxs69yYI470eGNi6EDSNzg3qomoNkDBuiq7FUPExBwpi3h8PeVn6nVH
cUbtJk9VSohmxhJUeZweH9tXMTVCXFx5id0X1ygPvGF9huxtYK/gZOWTWY09XDYF
De76WjKcfunrxDKXaqWEwMolLr3OFCgVS035Gh+yAzOt2tHz1+qF16d60AfpmD9j
hAPdeI5hSfECGuNUlfYu49pIZc5eas5X4Uf5pQGoZXCVp2VUUdBha0qTmQAyM/va
ixETBnHHKOpi+uY8A8H5UhgVzsCZFd5rUU1+yi26BKXDIc6v4qNuLsbTPZ4jTxOI
5wAOLRf3uxpX7812qiHOH7b9nn1ZzzzLi6R3uXaAa5rWYVBojdYCToyMqS3OD74F
4CWceOJos33at9X7xKnKPcs7zL/jykTh7zstJzEBPcEwtUAhYpjR7gGDIVNRzzd7
DKOL7vpGtzntHqZFgJF5QOljgqfe7zWw1TyFldL/tJ2nMHlj+50vHwRxI3Y0TQwD
cliXiUSPtj6KlMongaIdtznOPzuYAkQwzi6jmkqRU3wGFfxMNYX2NBd/kXUZr+K5
mOT8OObZ5UY2qLq10GrEkV4HjefRHKK773rYv1fP5se28xjtrhs0ElToJaCNUk2d
rbaQEHZpIeoSg4oxTjBEkhEkUiBjYyJ/AOiOpRXpKW/NgW2aVYqwnzR6XOxo99du
XNbUvdJUjkFu13eUoKE9+RnvTV8Q/OYw1Mn9SgIBTj8PVBae9oHH9yh9Av+qsRaj
/uK5vHxBV1tXg2Y9sC92HJ1CSEeNYlhtK1WI1wZ2IeSmqxz4uclyKq4OSehJCcyh
XhYsNfDTP/82IL+U6n1xPPlJmN+sedK7gGfD5w44//cgnk/BEquFkw9xzDf6mAX0
uKenm+zC8eKAGgyt0BXf/oFOtczrYgsi3rlE4cjIX1uIDhEzwgoEuR+SQ0a0zlFH
TwWBKDao59wV9vMFal93JnVwYCvTjWYWcpTVG7cJlw928Sx6lW7dWo14Aab6FeRZ
wvAv4Uw8aJLfipmXgspweR5njITa2zFnqda02I7QnpHPgsZS617cznL8TOEtr+CK
/qP0nZwhvBx4YkH68VYKkOYrWyNXs79udnXoseosv3z60XkGDSPAhSuBcXatvq0a
j+Yy5uR3m2ZGyma7eZQhAiMF2HZrGDGtxbgXKQoFO0vbqDFf8AOaYUOUJKhj68AN
Zd4PmW1umwH0Nz864oHcMXC7wQy4X8skX5AoHeBb1FECn7ZAGpDTMAzXbBjDuqqf
jvBxA3jp6XFYn1TZm5LWy1Rt12eYO+MqS9sUZHEcRXJ7/yyAn/0vYB6hcbMZRayP
UUGZIKP76W4kYlku02+bNWj6QPVjwMdv/emoq11jZPO1CLB/goY6QYmoph6bTOoD
GkbtQhmRLCOm5HuzqZ1jCsTbIjZIUlALNojh8snH+bYHp36kvTcuFQXalnhEryWI
SXNrqZVunN8qesjJYTbfXw8WSTlf+lVSuaTKYl+p2oQqRnEmXXt0atX7TGT/xykA
qNC27w2TGzS4VdJenv3Fy2e9FwLpJTCqqwrJ98wtwVopVKpTgOxRW0M7s/edAAyd
0da1cx0zVJc5regWrFeqkkwH/wTZcTnoEq2XOARrFnFZfYpLEU/gSKAJ45s0gdOJ
WCIv6cZanfv7f4tfw+OSPibwcOA/xkRPgybdF2Th7QxK18IMak6BiNNMe2mjgmGK
5MVeU1SlNueblE2Ox17Qg4k03LAACw9BV/J80E+vPr/ay1MhYp/wiHzDXz1t03gv
Jb1m+vt4LUnNyCmk2+IIoc6RqrDnE0+tfBk0pisu8eTbY514z9fZep5gASaloUBi
XYSPvpd4lPq3bzJoAXJ20HBp2cUfJv8Ews7jEF5Cia6WWGdiEo9O7rnpzxrUm6Lb
mNzJuWXTjBwtsRggkmpNlE47+lKuaHTh0hmDd3nV3T5wIfcep+t6nlcBbQSQw+TV
D/x+G8Hvckos5y7zxRtJdowU4l4lxPFj/bQGGjbmFfTUBbSmvWIsz1+Y5Vd3An6b
lyQ0X60tm98w0rXhi0iF0mk0iVG1JPi/cEzb6cL3HC5FhKGfWYrxDSzI1tJD4yXb
uusiwgAzR3sc5jlndHo9154xVv06sTZyYaCVhUsb+nqhLzxBGTdrIjKHM0YYJr5+
GdN5PljolpoRP+UDhe8XBYb2g1ZCsQNletU6o1wv4RVXrHlfUzcsFKOeA/njd6O5
LetHapUm+ZI7TfhtTBwfnOGxM5p61Z6B8Xq0wdCIf1cRgxAQfpr0d8a9wf2XH7Vm
w7frMRGl+xZVe0IPfUfnUeWlrtPdY0UqksKdxeKmX3TgTD/msluX/hFo5DnCXTjB
tW9CU0n2SLqzVkiW7MITzNijol9CNXCh7QqHwf7w56n2i9TrUc1lvB0+MqFIoJ9a
kyeVNWS0cPAJrd/9kOqiuhej9aRGsDlBih7M0vuINr42xfJ+949yeZkbJJJ+W7gE
SKsZiv8hOA0c+oQKRPc4lxlV5a5ljZ0MUCvigw115QK/Tk402AeUilymDuKrYNtn
veFCNcDjhZWO4xbhVXC+7lbqV73Bp2avQaHHhEardLxpFZz9FbEzdFC48sddf34U
J5oLhOMmAba7p+tTF+pfEn5ojx+pwadWWSbaNEx41jpXyjINqQXlgrB9lUF23y7B
Q1BFaxf48ZfWRwW5T+/R5t71LkPJrr7awAAFRsoms8ABacxkFJFk5YjskoFXEEnl
L22fMUh8D+eX88iTLvdwXsjfSZaBGAlYm2jyt5FZ6efUjllfbtU+fqwe7xCpnDUq
ACn6QrniMWzlIfAq+xe06xi0wChD88EBLpHdzy3Itl/2c3LiKCtJwkdgkfGpwHY4
ML5D8wPYuGpjMOjfS7xULNI7vmwpGC5pxniZf81CgUjTEk1cGi+EFVUsXF2aDMjP
lQpPMeJgzGkjG2fKmCuq3gYLIttKlu2ErMkV0Xj9foQnyaWUjGVnKYAm923lfCJ7
ijG+Ll5wrfA09+Hzy6PQ4opOnRMD61G0hRme5472kstkUiNr5x/F5rdfKowFRT3z
fdb4vqOaZioeho5XnB28STHMDSbifq4LPLPERkfx5xdM3OQ2UxGAZHqroClr2QHf
3jJJd6qzK6kWvRbmVO9NObo7ILpl9j6O7SD7hZy/KFjZafXYLRWk0kTF5ac0NtSB
SlTY0iGNpnwGn4bAty9AItSQMBNeeo2m2B+sXJcY14AehgykDpVkAvPEez25WFdQ
BObXN6jU6mbpAVUQLFLd7qIZM3AqUa4LMFKnTtaVBQYoccpguAtcclbj2opZz2Gx
KuCo2CYCG6jx9KiCKTXTOSsRLSfoqfaBcCKytjWuBxj70GnYuuFT+UV+DHNUkObK
UKx0pXq6KecxloViKWdtkR/kYsVdIrn8AXN6+Uw+sjK7ctJUAQXBGx0KFimzLFfl
CZoY0rHrpqXTIt/N0rLWoAprqXUjYgmyujYCPtyS3nyGmwSh0TeuAZ1OKBAIMQEL
XMRJYYSLf3PSok4SKGlhj5YZYXzygZWnnbzAhTeWPBTn7cjBhVMxX+pexLGH4bTG
M6m5PegsoSnEfYnzZJZanYhWIMdjpHU/Jbou8fb3Avx/aWgAeeleximm8TyncEQK
CaMpCxboskUp9IurFLR6l4x3NomSdGvrY2tcCUumTQOIwI6wD6sDjd41cvUW5cy2
3ApxT3sRFDIhysrOc5DOY2opJURjTndXqEB2okRcU9y3tF5qdGw5BGVXAGnQmeqE
ykU+eYnGW5jcsZFv9v5wA6vbR/dNYT6ZvhnfPjt1E9wX5qkxvB8PMPeOrQkV/XA4
UKMaWmaleqsMgYk6aF0RtofoKF8afPUWekGeuI8AlrFkRUTb43j7f4Fwg+5GfmEz
QB8px5c7bQn3U4l2ZnCP+yszW3coqccZusAHBjTXAlV9zM2OAwJPsvbTTrdPMZ/z
gEFURGMvKaIYD2mqrqgvPWfqzluAJFbZ7fKg5/Q20vW1I3/Vp3tsqosNJGDH67c1
Yz16FFvx9jWGfv+Q4sBRCkKUttUxnARJJUs5ZtUKr7heqiHLl/YTmVCri8GU4A1r
dSScHv1Hk0B9yNtemmnUje3Ud0186K+G/XOldcJ3sh0nqa5FAMuaNsfxSMWsFNhj
nTv8Bby0CUxNNwjd50hW7k7uVh3Gc5wX7rLrhbmE/usMfeNNI3Z3USnS7D4MpWeL
HTSrXM94+k32liqC7JG3jbGTgbl9g3WAOPoy3WDc8OW4TT4Vwf5wpWxI4BoL+fgj
obu+F0w0sSuTTRMBCvRNvQCLnUOOy2CfBkaI1Hf/lWDXtOvBLY8lmduMqodjW+M6
pFnYCuOiw5cLgK9NyJcJj7Vs8LPSbHAKlllExZ4b9yTFPpDjdK5m0uN2oH2IjB1c
BYJrHGpsnplS9OoJIAoSsdJwClrQsbC0hxeIAM8P4nreo1EnCnHpYveP5+K/eKWD
sPXxKgJ6JQX9GUCPFsIvUQM8jbxtTSPWHrbf8LqqLENK0eXjFgi50X4PsKrHtSUc
7fMX99FWPtRGWqDDMcP1nSRDn3RL4+PLcAISs6Bkhz8MWQxKOdqk+qq2GBn2Ydbm
Df5kke8Dpuf/UoUrowq3IxfptrRBEbahJQBAp/ENBggvE/pEd+UbcVQPvqPgF6b3
pkgzbtHvPwm30nKhBrk8nKVz1yDl7EcGkJy/foazFUoPFqvC7rodnyK0SYKezwE4
3P5GBI+CCKkrb3AdlAvi2Ik3fkJbBwz+E+vsvHKxLn8W/ecH1Q2rIrxK8r73GpTB
lxd22J+f7U1RWnx01ocoApYYazvICLYNVNTK653mg6CwRciRJgebv2++yakipN3B
LHfvylymGZEV5XSOjlRIj1fD7I21vbkva+buaN6hsoqHYp0xqkAvQLkAZ4vcimAs
Vs4T3Oxwx4KA2Zho6WYsvpDoBJyUSUNUcTvixJ9nTqo74OR9yq9l7o5S7VPbVy30
JIe4AE8CBoe3FM4NKgs6W7lpFL7eyBO2vLN3nfr+wgpK1JoPdsJduL/Z3elIwi/K
NIhEV2BEs+KrlMiauy6tIjEHQ4/pt/ZK2vUzBqMNsUfNlPuN+jzhe4Dv4fAy17CX
UP1g1gZ4EOvEQ1WUlYq7umLkkyop2lkYNpga7q9y3YWR8/BheS7VGVgyqLRDt/16
1MLjRJTdisAGqjEqEiPk5QvWNGIu7jG5aaqrWh6Lf9tDafe3sUCkjd7jidBqrvmf
AqdtcIkEGbLnJmvRYXyVJL3Dlo6ctCdr31/oaG2S8Ikwl2xSn/QjORsIKnJLLFnj
2Hlu54ICA38rVfoLXs/BTM3tJvPBBWC1bDoZahQDUEtf6NjfmU8BW2lGFIsQLQju
PPD9t3omEBt/lkCUT4p49wctDpN7oMplXPw2lDK/KPdHvVOXrBLmBwByNanQX0ny
4+vllBa3X4b7AuWuUK/t1B51HGn7ic50/WvgjEJ+GaY/j82ObLICI355DeWEmR5t
qGUAtHQvcpctK9oY9ZfRAY8V1kzdYiBIK0y1Ev96J+fQiCMW5IAENtBccIM8IZDT
w71bWr3YBut5ibCuCBsMnp5pSqdY0TI3wjO5L9ru4/isTvUd9C0U0mYSBHEwq8U+
pzDqQ38dnXZ96udUrGMLr1HPfAVrij21va6BeOBDq/eIsi+7rBHz5CBDmhbc/9LD
cm6HJk0EWnPoyeO24Q1PJERaoRE/vmbH56adsZggNQCe8k9Q3T48pgnXLAIVxLT1
zE/13+BE/xceHdNsVfqxpGdgaaVHWWHaNANHEeGD1K4FVhCAL1DuIDb+lfE4sB5F
XrMRQjFMZmJS2gsbW+8nyxvXveCKS3TK95BXDaI/C7Bbx1KXMC98iUNmypb5OQre
KRMlz0a0W5qIFPgsAyxyUjhSrMtCslEnPB7GshI8MvD8tFmHSF1v4QEULIBxLwje
0oL9x5VexD7Z4urGxuR0JsDfUVe4KAX0LUQjZVV8BtZqIrDOdiepaUhrQZB4HkYj
qUCU9xL7lbgndbsGPQMzijFIb1BVMVISuTxP8LeH566fEvDyNMXU818e3hCItX4k
Zj1uKarzSs2MIaDaeWcf97r8oX3aOkuSER3dqroF5de/MBFMsOzzvZAaeIHgr7FB
npCeuOWQnghQMzruneyncjdanHcXUevveTqImBBmS7K9bYPMqfadvptPQjPdM+3e
zf+AZxE0uslTwmm6To1+FGeIryJof1u3by4e+JiCne0oXbyi+kEag5Yh45EqRZ1D
to4b3AL1hFVvdbNgEWzsvmev2Gil6GNRIRfYF3WBNG2Q9Kz5DQ67OocL2qSj9fu6
/50GB/u5G/Gf7bb9ykKs8jR5yXoAu8qvWVD91f9Yo1M2iMTpDg7F6lIgU6Z65lZI
k89OwqKdCkT5AugzhQF3xJvYuCi/P4AjeuUq0Hu9ESOEjlIxb5H4mNf0Bf9Mlifn
6IE9xRV8drP80I3vIyjTr0R6SJ/ES6P8fYCLylDRtfdz0IwlW9nPNRwxN+X3Dq/D
rIP0wYPg/cFJ9jAqQqaEplmJASDWev0gNRiDvwyWm5ZXWGLOcFl9IQEVwuyOWWb6
tx+AMszSVg3P4LuNtvR0Lo/kfGD8/9yt8+EkV/vNMYuNQKaeVkIaYccl9mvwcTSv
jSEAj6gYgB0rF1SCbGLe+rHnGaegwf+jAwrzsArVGyQDJbADi1jewPugQhW+AY4o
qcpdypY4iAQVUvSqPH3mclU06z0+byX29S4gDj3d+JBea4YOE+oxdaUcA0QJk8J7
f2O0RKcAUa/EC+WUk89eD2hwxK8mQ6jwJCiMWyoQV+bK92evBEI1WJA/1DzGNYdJ
RnPndc3clSdq+iDCrYWCgoCaQd4qaq7mQ273Lr9YS4bzTw/lqmPPo5I3nuLoPPzP
wpE332YRScE//dvuZuzOtNH0/9F8rxbbc3uY5A/T/GXq1qZy06dHmRIQuhe6f6bl
hJS2pbJho/PMW8hdkpLVQ+C3YL50XDBeJ7/uK5m8m//9gxx1lAqGfIlQZajBN4fl
R3YIf4h9nTq72Lgk2Vdm9yhxHdOL1zYV+gxW4zFltF57FAEievtiZGHAuQg5J9FM
HfNHaKzG3XVWqrzPso/AyrmqY553Jvg0jnS9DJ2Goa+3W+Q5WQoQ/fBmsgbiTGqY
i/1SeUnfK/0Z5COq8TC+LsnhvlVYsdRN9Jqg1Vn2JwW8CbOCYrdaA8O2nVXPYQq9
Qo0ryJ2PICv3x/MHZWZYHn6kjNeYI5/Glc8ULmq1CwKJ+XbgvogLDdepqQWRpDBj
Hr+jUogjkM0Q4Vvt4GOu2OPX9b6aVNU1gOXQKUYBZt7S4Os2h1JJqMhKhnXbeMBG
luIIye1d3mjZvrOCs0I4WnxegX2jT4W39mNuwGLN6eJ4+QLmcIJJWJhnwcOcekfK
h5RxvR3JsB78uaSngk/KKmIP7QdChidLQ9BkGgpLXf9E2PBFGZfxjXnKpVfbfLfn
yIqbPAtEziLRr1DOmtRs7Gf0rZcLaWX6Bl9zHWLiANIhMw7CGXaer5IbMxa92Mzm
wX2bNwGDrCJaGcvnDqAHcjNwn5N227wq1uWXh6QVbBzM3xm3ekVazLhfh42GuUrx
QEsueLwJ3mO6+5Olk5nV33g09iD/bhsBA3mdTlCKoUSfdJ9xEgn6XnymMSRZdJeH
MybMot3i4iBphbzjQpNJCyHsj1JRjQjkZO/h7o1fLf4+hPAw/fxJHgSNdS9XwF5N
cM4Vnr4h96dz7de8oSs5BT6ovPsW6qZEJav9nanr/icMW/P8OBCq7TdujmTFg/Ma
Qet5DbY99/jNmZ4+KRa76UFcagPocAx6+EnU0S7Pctb9JbGVW8vSLXroEnRfY2kE
IsUFCIlcSBHR+M4iHPPJkN+pgXfnOkvpAAbsa+0Sn96F6O3WbyWUiRq5C52fUefK
DG4ovyve61TayQGONGp62YiUJsUxPbAJHPUb2rGQEyefqZxSRUlwpOIUoiH0WABK
sFOV262od8fLsL3V2Gxr8sirSK62zfNvkFX2CYEf+6vAiMGMeX09hYcPAFS/18hT
Ss7kovQwKNQB4U2ZeVf75zlQfm34eza4IW0RA23ezgSgPFzpx8Lygi/LWAeBaDUG
JyZYDi4lHFhwqSF29g3mfXTZIkyW200gwlg6/6iv+A9RtghyNO/jW/5ckslgSYhw
BkuPCi8SpR9g2zrn2K8mHim+twQcNQREQJ9xnHODUdEB8W8WTiKWykvWf7otfZtX
XZnEC/K9vKAO7+P2yY1IYSsfrOWN8mDxQeikvIfg5OeJ5m6dPSzdcsxrKtVKKp7j
1fE2Xr6LWHJMjafQC7PadYO+Jem0zAGsR9kIHqAdll8H45JN8Num3PpQbJ4MlroH
2Il0ievZz7M/nRNigPaX88kFWHawSwOnrY/HuLNuuj7/Cd9J7kt80qJcRqWu40xz
LbppZyZg71n9nePucHiZNBNK8RUToQpW/W5CFWpuw/H9lr/+OWX8gyvb1Uf005cp
uTzaYNm/bwFBcPGnv1bn8789T9eM5rPVP5EfVzO3fTOGF7ch+j37TFxmoHfc1xe6
cb0GRcXkLXBXZTUr/dFUxYFGJsgwl9uzf4H+QqjIrPL4OvwQog9w+i4gSW+APVz0
WEBk81DneX7d4TyAtL8Glzqtpsc8Tj1RalmuhRoy7DTYW88ezkAb/JCtGCoF3hK8
gOQ+b6KpKdm6Q6Dc1VwNugeKenyoGHPFR8BOEDmJsnmcGgFCPZ0mGlIzp4hU9zDX
amlZUSZBBdX7PwzpQcWzBeMTt4991bddFtT+dOzoVqOt2wyj2n/u3CLBH8m/WuTd
3Auh8GhHrEtLf7ThyddQCkdhzlA07iGw836TIbkR2/jnz5wV/wgotiIOxPeiqfsP
kz3XrywDma/b6QiLu0nrUWFT2m7z0FZzGHy6ZQC4hzZVPRLerZiy8W5nDKfiQf5r
l7dNhuRHtPlZqjOK2SAmsG8O8pE1WIpnHk28l3Les0cDfwWErV3TjfC1U22pkMrr
4skCMV3omg3HG0U2P/VLfzsPAlN1kiVa8ddqxmu5niBLn7geD0oo4TGoJTRlqo42
gIj5O3Q4PhPARncb9v/a3jLQRM/nHcPjibKCMk2JYiYvc0A61i+RaZEgbTe2VfSu
VL5KD90B024yb++a62M19U8507fG4a80YmXr7UfiwEiEm0hY3OInLrpb5qHxudLR
tatgcBOZR+M4athesjI373nm9nMdV3VeK/aPiKnTfRH92isreF4nUz6PkAiAh9dg
vqGxHpYJTG/p5PU+DDoWerD5FnijTU6xiRS89/u9zMq7mAs0jmgn796kyjfLBCqh
yym/sPK6d3K7MIDgCUzXwISyUsHaC5jrp6TchSCVrIMm37LaVXYM/+KYGl2HeJKx
W8c9Ou9qGmkoGdIc/ei46TECplzJKTWd3X4FjBqclCOFhNz+5leQmKAlVvqN/kF+
QdZ+tMUWNyFWJoFc+rSTaUJrT1Vfst98tG/ZuQaNSMDhjgeQe+MM/cqQU44xKyak
W3r7U7C5KURUGog2ysoDp5Du03Z02C0R8JTEpS6fkP6g3mt7FHiIL32VPBeFOGTR
lbz2W7MVtZVFiGNS1z1wk7qiEtsV0NundyQApN4YY+6kw/vRmW8BmaN2qM9X3CMy
sXbmfJJWQe0o/USq9DMrj4FYeZfMJeg5KMCYFgKCH47GvGpD4Khhqxb0ZVl8wXY2
eC9KAsNXl1XOyIL68SvnTbpkQq5VrXVOKizloNZh/1n4ZhpIB+2td2RmyEpYsKLN
JG77TvwZjAGl16EV0P8q+FwtlFHIpgIjWxLyhajUuORo7sh2W42+HEpNJvPUnUEo
sjLeNhLR58en74/c9+UrinPgasDb4105uz6PBPp5UH2SqZsr0B9nl5Jv4sb1RD3A
CkWQuJJJE+K21i9o5CHcBX2qhL2kwuj+Jx4A/T8T6WwgVaFkWOyshUXAadAL0V8J
oGEE5N8kPyw1kG04pzMXNsp5gsvbRn7W/KFqHB+rtia6+vu9z9CutfiofSU+1Q6/
JTyRdRFzQt8Zx14gt5JlrQLYHAuNtWSDNmjNh3HAYq9fC/6LED88xiBAsyzeoukv
KDL1SeP+rN2fHYhUOl/4Viu2MED2CTyTFROOVm+oEW1DFxoxZaBQGd8F0/FaZiZM
RyTWL8Aiy+tnefqkCycqiU7DKTk0wpEvjiSatJ4H50vZBYTktydmyEFBdOSco07h
xZ3DE5oAMH3AHWF6hJHLV3d75xAheR+IaeNsC84pjfP474T+F5AnLoJS0vqRXZGU
h1mSM8cw7f/OrZTFL5jjzTfYsmZgn0xLB3hPWccotom7RMyr4MVjuF9qBGm6laHs
JVbfpi+vOuUNbcqXZI3mdIeDR1oQNf5iTPN5h1d0SujCJ2xBShnv2NH+l13drqLj
d8Im8VZ6BufzNr4KceJfJhblM4yNmbbTBvNO++W7z7F2lx17JdjcfCFLWKBG4uRY
nnf7CvhPhgh1j22joaEsCqSM4oSIIJn2v9fIx14OLK4c7Z06rpGrxwJ/5+puajx6
Nj0rOgobAeilZbQOuqenqWvStLL+gck/GnDvXMhQgMBEOSN2eZBXRliriH2Qb0XG
qVttudCQXeU8QITuYpi9Ku58XzKhwt2JB8v57qwsny59qTXBfauIPmqTbR4xitc8
1hi+Rlh7U8t/xZwDzAp7cg2PxEE5sETCOo6/DtX74WrHXweOrZ9wWhbZbBU8tSOP
JIwcFuhSczmnA4/LrR06i9xlbYZRHklI8yDYADLfup7KUnHZXsn6g2R5zwRv72AI
WKORES/OwkmgaXLmVFKuhZPVWhNQL8waOQ4LvE/1r33/wGtEOA5yWrJJAlN7N4ZX
YnJ0SgJWYyXNmOqhpRqggtsop+x1sH32T7ElaD2EFzxKn7tUhtUoOS1nVtpS1pR2
8g+LKRZb+4EdqE177joMFi/QMc6Rh+F1R1gBVJHpZcxDwCXAylEgjfh1Rwf2Y9+G
DfSN4jNxP7c3EjAHUjz84DVpuR2TCdkjU+1OnGKyKUzyWgCM4/1ki2qFpMIeM5d6
RFElzQwn/gs8SLAzomWNMv2Gu6APO0OUHx8qefRg1kWhPXEZb4r94oXwy8H3fy8H
MYyrIDRwou+6ezFC+IECWvpCib5F9cMEWynMzhKmqa0515Z1Jtr47tOy0sb6OMNW
ADb3yhWXV5B/1g3CfTTGtJN0VwE7kapUYSOPpSX5wYZ+/QWiwEQ62/omwrD7eo2E
6uObNvQIIlREdDzgrWb5UubU/zFuIxl+0ByESeNe58TAV79ydhVzSiQ/adVJN2uh
mhhs9q5lB0hfTmyuSiUTxTumAPEOyO/O2kukLh/xGyLXklT/Un4bFuUtyUCx8dPW
ZJi22H/MUZZdveLjMzjZmkqoKh5D48NNekX5mDbPLTqCpYWFODDanwjIk9izxxRQ
mgSwebO8jqvfb6S1GL3CUxVKwu8fA5Gr98d4iDZR5dpcWPbJ8Em3fQT28ztlbhPt
GgWuXlLC8jsgJAy4GP1jLhzFNysX67JVJ8uu9pEpZsC6coBYHZzGy0L5Pi4tfEXV
dFJuPSZzY9c2qLNlS1hOxDl5WPA+4kVOjL6W/IdQmO45jjzgsX/k8Fz0zGn0461u
UPlUd/fvO9WiDxNo7/yG3gNtEDObU7TXU5+O+5D4UcXW6EtMH4D7FqNi4ztW92h+
ju0mJ8i5B3kaSl7SrwXiRSJPgEXj6y4gMzqCXKPFwgRylMc1fqDTIFh6txY9pNsp
9mWMein6a7l5tF9ObHBk01XvrGAgK9lAmR9Vp6cwpbUMADyns42H0OcQjZseQ+Td
cr7BrMhQL6XGiBcv+IkFYZIU+gzTj/SrK38ZjxQKfr0M7W1WGv7nVnW/76LTenyi
vAk06Wsg30UZ+RHkB4/1gWmc0PnAZ4B4cFjP3uFmBLj8bOoFndg+NkclUAXD6Uh5
3WGyowTAhYbScr7M0z516hYY0fG5GnKhLIO4G5Ghq9vfxeTUQOVBeH1pai1KVPlK
Mx/3o6v7kD9W/i81vF2iHd31VsSJTP7Z1tkMg8kL58h3LLYv/jQxBDlniR6x8v/M
d3oylrVQBOX/byIBJumBt9sVSjpcBa7RrJeMzdE/NEN3vlWdJyDkYZtCaNYGA8N1
DmT01FgFfcJpF2w/xMsRHPnR4e70OBk4wTuCJntDN1zxtZlzvH0X/8FkMNhmdbPx
g7zfBIF9hhEEAk8XsM0dW8L2M1fb1O1OXB+0WNih+41B132yRwZueuZv1RV+Dedd
1fFFmdjITNxVUYdVmj8q6hKZu66v5w26CaelrIUcwQ3bQnfAtWQLs2aTfB3AvJS5
H/QUS9LgKblEc8NUo/FpLaJcRL0rdJoN849kaVYAVUw=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GOilS93iPC+m7wfyKYlz9SzML4pjcO+5OcxIS0iYCxutPMpmCAeREoWzX13oZ3qV
HGZRA689xOnv7+n91qEPK8e5eBAKlCHISCOK3GTG9fUGlS+C6Hh3noU7EaduozSb
QF/upg+A08tsvxesfbcij9eWolZUyute1WR4+2anDblYiQlNQHH81WuAg2+jqx/W
h4vtfzo/9zr1McrKeADQs+ZLYhfVAV1pgCq4Zhs4OrKpUxsMIcptKysbe9JhVzwV
RSlyCzLLR9Ly4jBfb36tR80w5BoGDLfM324XQ0BLllxGIM92aSHXMQ+L9dbSyHWa
+aNXkYltm76DVf0EAx6RoQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8096 )
`pragma protect data_block
Go3+wSA0LAqciuN4QGbQ+B0OZ071/+WR3jwnzXDAgJuJrrN6zd55lHmSinKAz9X+
pvyccpofvUanTz8pALdAPvyFZgGd+fVUMPguTbMxzcRYDofeKhStFBwJNK8dwhwb
Kx5dZfxEinfy8fFJ6oSGSFf4RSBzUbUshs0wIEmTonFT6NCt83UbBdzq74QwDv1s
D8YK4lGnG1EKlASQUMs/j2SAXVa61kpJefn6SmKO9dhVlnI1FaQ42jetvSFNfL/2
awKyaPULpeKl7kGi6JcumcV5GQ/u4BgJERu4Cbrx8mJXFXVe/FyloHNPrBJ/MDg/
S4D3PwSmCHR+IBlcupr/MWAG6TeXUzyCoLzcXSQ3tua+WCAz9R6kcAhzaa2rlWn+
uxnH35qwN4DBZ/s5cz9qJe7puVYBJv5i2DkWDh1V/YYBHgfn4aHh4tXkVqLBVsL0
vAqnwl0A2dzISt4rI5nAU0EbbZpSwkwFILgSjASnZhLrRqXL/0Xc/x+LHtAcOcnY
AEjJEMAqu4ZG4MrGfTosG1hVrm+cWZNFq9VnZZ28b/fi22iuim2c9xAjBiEVLg52
ghece535I4pmKRgNtv9hiqAWSmWJXML3SZ7Mb7c+0ZXeZw2SonQLfvMNqYkwYG64
Gi++TFqPk1ePn18PVGYGmeeH5uPyBaJ172D7xjgXwuot4OTREt1efnznPxsunxGT
RFDTVOwMJ9Fvsx/NZlny3VwqsSUCGClkNz10brs9mrbEEMfBcZchkePmGaSOZJhJ
BYeFvuowB0NVwn38lcD0Za8WCUwGT+SHxnz2iR5lAiJG3Nkwv8dkCjElwZK9kGDX
Lg2Utc5vwoZfFJzdYsBj9Lf74r7KxhM2KaGQbwuMJC0r4lV8kAuJ2BlZ8LxBG3xw
3NpdofHmnFSp1V0ppXnGYBPViSU5WQFDNMS2vZ3+ugtQyrnRN0Pic7ll6+QJUSCG
LCoJVyVu0x+Q2Dml0TuWzgCpue7qCmFQgLXTjP52cZTmJhbVJAcm9Nn7VERIhg4H
J2on1mmj9VRAl/7lICphomJ0s08ohxgumvb+AhdTQjCj7HwMV8PkD8LzLY5z0yb3
Q4j2bKx7pxE4D4QlBu1dJB0CJ4o52p8gjvoX9trqWJkfVUgBWQ354BKjMi5Ab0Qt
QvvFnWjXz732HBddMupDS8Lp8wQqjztdrhb5PFSbcChWBzg+edKeWC8wS0Iap5ME
gMD3rI5UPSbS5LL9amFbq6huHK1CkgsDeiW0w3ldpkuA3nAKor7yvWkYlfNtxZD6
sR+FMOt+TBSz8r0DcWtk+8B/qCakyUHk/H34Qo5RwVcFfW2VcoqKI//Zl+p7EjzT
kAXfhJAkCh9uGB7pOxCHCp7dYw7NLvTbBtrhAaJaGDUaUwVC+sM5aCIzCwY0Gq8+
0daynd4RJqsBc2+9FSo8oow9F3qH/uz9OyPRbOOncPqmpUYahEE31QM3iiE4nblP
xRYcWWxJpiIHcxWhxrnoq4rUSIvNo17W7oWbNemJIys3c8ar/ADr5H4xiN3S89nm
s7RkgpA2QwYCOgk0P+KxxaNy6DBNOdgNKKTB2CoZplgArPK0RoFMjihLzW3H2eXq
v387sHCurt6gMJmxReBjaspO/30MOxVMRg1MgqrQJHfr2JttfK/XfL34iHOTMzLW
/fNH6Wp+5ghYdf4sQBMkQHQ3/A377omu2efBZIMxdFz9aJUc85rDIax0OBdhNAEB
b8XXBoAx4gS/htdihWpklZ5vftcH0Xc59+xG5JK4Y1rHgYVriEKbq/3v09W7seTp
it+pr82HmeAU1QhKGRP8eslgKjFKePIw8Z+wuqgZ2Q0iO0dzkZeWEMPypx+79a04
Y0vLgvWFdHzWtC1DsxJKPpRBW/p8BYycd6gdMaIPbA7FiSz8vsRqcJ3tYphXyUzD
yxbpfSA82UXFpV8HlWzWEzywJ95Pj9Hw8t/+JHzFsv2vu1niZRCFFRbH3ZUK2ux/
g+IrdxJKIK5wfUrOCtNBdwJ+8UwKhXYf8YkGFus0H5GvvRKqSjgx0ELKPOu3XXav
XI4Fe7YStxpodu+opf/iDkw4nUfi4G/vECVk7Wd4o4ApJVrubEq/TfeZREdn0y6n
Zwgims2RrN12eVfldmZeTldbTojOENUWIwn0cPQwypW2W62CIesQpueRvPs4tbLV
yhTBSx1brKGFVwJYATltJz8JzvRnuzVSnGW3P/+DwO1TabNhInp/ZPTiyxrpjKiq
kZiTleL5SGZTacd88nEGCuweUWVZBBZ9SRvOdjWiTiNUtU0LcBTr77uKstHaIxkc
dcTHZcyUUMM2EcsxmBh7zB1eenavESIgV8kH/otiRSUuckyJI6ByyxtGk25/tzqR
WsBUSTwEoKkbtK9fIVg25QQBZdFYHHGsBF01npK9uC4KTdcLzcDH6dLbGEwU+t8y
tJsrFQ1O1Zd68WzDR5DzOGxDC3uU/DwxwOW28ONLlEFNHRcz30OFvr3Sw50enQdH
yohTzRGKS1kXX+zn8RC4fKxqrnx7kp8nxA/niMSvbKFZGsuHlc3VcwaftXYQOteb
2DvrUketJL7y1MtcRRLORD+ysIAb2P2gkiMSiTmFx/0VpkP+w6zHWEsfv8XOcwwh
JqwStKFrS6KY2cDO72AgmwelmJqc3AcPm1OyvX/gz/3VtSPC23ifG7HbQroTqLDU
YsNdnKt8DJ+xsSB5WV4cPizjMMfhgRV8kFImaNDDlUz5GqPH/3l6Mh91+KZC7sv+
/7mlJrNQ4EmkH5N7JzX+nV3yTyBVi2hAFoXOZh81zVtDbKysp8uaMycC/8c98QQq
Fv7GAYJW0AEdK4jSj40gtwZXxszzhwIct4767pdj+2zebqb6ZIurPiyP/VzRqRZu
UgsE1Mb1+YDBtBYbevQ+DFdPTZUQNDJ4h1WBcwJP0mI4LXUcyNCHOFNgc1z967W4
5GzQZzleULVGDN3gH7g/fhL5OccQk0PtdKO0lWwdyw6Zx/hiDK48GS5AGMyKFQLC
h+4fKsD1OyRVOAF09DpbLepGtXy3KHYnvkCmz/ar9jIQQag4TdjJZovmJ8nMROh/
uV8vX5DncZuTRk0btBpMwEiUwiPCzbB0+0PAHsH3MMQIx+63B7neHFcoG3FB7kXK
4pkXBNgNATkyykzus0J/hr6yGjZ3BCbs6tCNx6fmX7+CzNc5z5DNKKIjv3da+rFS
/5KmBdiPNugHm6Vga5Kx/CbPAoq3TVhvkefeXMnGeqB+7+ZpFuFV2dgfN/B9zvcC
EWGhd1AhhXld/DfFAukPFaETsT0mcqBAmh5WPc0E64a0hKsdcicGM7osluj6QGtO
4IY8nNH2S6n0+mc8A3j2PDSThNvGkS4ENy8/yANLaE6satqWH28XWgGwT0+47M8P
QlKoX2q0P0GyZzpcXrq1ugGmchEM8PfYBAycrvqiXFdqlzaB9318HibC9abJh5OM
D8URCXOnKCtUr4+rP+zBJ8T7Ds+gsua0Vbfd41aPBqrAUkvqb2caxFrOANt3DuBS
9JkAxb7EO0AwkxduMFQ88ylbDdM9U1q62ulKqA2W1Ea0GeULgu1V+MyToieS8w5k
uGlLVLfqkTIwEjp6SaLeAVYe9zwjCippE6Js07HOFBFJ5/+5LsvpCtV7w0uJ/q+x
7plO7DDZnuM42if3Cv2nTM3M/UCv/h9K9agdiJrIAneO0/kqfdRqqWDouS3NFMzr
+EFQFFbGMFm2rtLb+UeIzVrtoaRiUArSnBfiSP+uZcdhHVrfhy9k8tfpS8FHNIRb
gtf0FD/YXA+2ULGdB3gg4/obK5BiywZp+oaKFbhbVeYY5KNYhWWYM0Ug3t91HqLb
m3Gigge9Ijo/p6hO+R4GWI7Yw+SJDPKomHZ5W3CzNeF0t5WWJge/IwOyz2mjMwpV
1IRv8cVok4fZrGYcd2KahKyHHnyzgXAHeuSlA/V5ra5nLZnxH0wJ6JFqr2lDEGw1
mfXLBDzB1eKKBAaaLTtbEivNwVU8h5N2gVrseQTuGeRypEZmGpjuhzGFW4GH1+rj
LvrqcL2R59An+nUdEKBjc4606cXZCUKVEe9rhxQR1tyjGzFtYDCwH9JxhdiFP7I0
6HXxux4yw0kQKxyqS/hU1kCKkDumSfawAHXnMTBZN3ianqzd8qKkCEjzjHof42kf
gzPAnALsYiDK9wgC/prOPlFtlrs0vg7aK4c6Oyy+w4CcsauObSJlC30Mbg/HdPT/
DNUlJRybr9hVQiNt1ea3/w7r/rPNUR9+tElIC9cnubTd4v1bdpZ13ETSetoz/xWQ
qG11no9PSkuua2Kc+YkPgAztxmvxrCE2O6inQeOnBvHhVatATklpjNtUbVUPD9qB
aOo+uDgNdwknbOsXN9oCyQi6pXWjstKwspiV/a4mnDQOjlx4qkXDutrLzIRgVu4o
8iIl9fDvUpnGSkxASU4n5MRFdQBWC5kj52Mv2brlF4OdLWntkrv1ejyQDtKWWNfS
obZxCYlj2EJaim+dPyKqapBSqpY/ylK7KQwaZ+5WVEGMbOG9HKyAJXnJCKw+qS/X
YJt8M/SvFR18KNC4GX5rrime9YF0aMoGsL4MAGYf+hFhyMSOnLkNsCLhg3pKR+Xx
btkaMs6AR7BWVr6yjRP3xCAnen8BbZNV6rbOs8lfciujXN9CAPFigR6Cv0UoDNK7
KCLYnXOyIf0gGfizsGguvzRu2PF9mrXjND7m7Mmvc5NPAMxVJMuBs0zgJrlitAPT
Oq5FwaVudkMOWxhgcEmWwrQ2PxxpEOHWaeHGDeYUVrMS1Pcz7EoqixGEuwyXYjeO
OQSi89clv8bnLPs7+DQaTbGwKQZGYvpuERAB0aT10eWR1glIgiYxjUSF9gALVTUw
lkp2i70rpAG5VdC77mkGY2WJVmOoiRrf8nVUYaogiYc5uolQygMSBRixYgBBUfDu
9indYXkVktQ5DiD4CRlEyTnCKjvRKJh7oJqthztmt2DnKCTLwqXDDcku0NqnkpWM
RTcEhuCiStAqhxyCmTuUKnDRYIBwzqOI5TG4pmzgjRqGokdyk9DQIsz3Tejm4iZ2
q09nSirw/ACIY1qM7zNgpX/9/w7c8lpg4qccP8agXHbfrzKkLLIa4k8JTRC65jw/
0lhd2NfF8IJfhaJoMH359DlN2LeXKhHPEXB8iSj4zIfbJePzLoFcJn+jMfwQM8fe
EF5ndA+3urI9lcyqrwoCcIrj+986KAN92qvqiqhfpSvr6s5v30Xm2RGH+uRqLJIA
n3Ao7qceP/Rjbw8rnSI2FvECOPmBq1FFTPlcAEVw+Itiei3BkDhM7Ap2iJUEX48T
qgOkQywlvOAtO40bQWPfgXmRA1gmqowviYkRehhhalG/8j9jKscLzARUBuqqp2+D
5WkbntnCeWAZ/fveHh2lJmemmmSPjjGxecgIE9heZstmPkBPvtpzePoZy9x0eZet
ZNvyasVMcbcGVlI5udBl+oBnCN8RRyYBylk71pyQXHeLrvSEsFJpsH12hEB3UA/5
jnVwPTfDt6PM0mld/AfjKpEA6CVtHLIUJ9CzJrVwb7rqvy31je9GPl2a14E+Qtxx
nZ1Pj43Trbo4e3+37o7lk0R4EqBPQ9Wi9lIm6dZ/+MuyITXkMJTF4KKfuvfupVfW
f0VSD1AX0MH9y89wU4vCi+8R/MCDz/ojUmGFz3YrhnQ3j0bCberDdMah35UUS7+F
nh4a0Vjiv32k5n6d1pWAJfgdU1QTsi9QjRGfmcDvNhCjzBGZWqSgu8pzxyuf2TGz
LTSHrvvJ9rVqqxRJZVrz8L2iWX5oegRNgylaBtnCmL2g+RF914OFDGg/DxGc163+
DYTqWaj5f+6xZattXFuC0KR4ZadXZlE2YR6msUzLpOa6McuWJ68H9bioEFfGFhlu
budmNYff7V96kQUsxbcoIcQQBVInxZUJX92kWPcznIqGdExWUkdb1OvkiJ764z/G
rAb4QfwPb5LtmBnfro/WzS2nAsMSiBrQPSCsGYFpfaWXSmYPnrxRfUGpZOWslSVb
dd6xJfOXGjssoT2BE2RKxpJ0SFJguf4MuKaehZLwxsXMWL/j/PhXR5ZV74PSFFVo
I3ao2iToh+yuZkQ1K6/MAEuPqJmQ6ETCBAz+YY0/ZqIP4Ep8zz1c1ccg+Vmgzm5a
XKpfW7nqDYSjwQjYpfqslECGUhBM3HprtRk+ODOkxegqGAgWMhpnlz7q8M8S9asT
O870AHFNHtLXhRebnA0oNZTXTl+4SUQlxnfQCHDXTLORGL+Ii+7VfKo5ggie9rGg
7/kU4ryRttoHUqN1bQ8RNG2VzcWKhJcQvf7uqer5aQiwOxOAoZe+y/KxSTHyphGQ
0zXBGJF9hwXZuGO8voCEDwsoFfPQmuTdU5YwE/B5BpYqWxqO84uITngqzBi6Yg4U
Zhu+nHxJMUi7cn5aOy8GAR895kJ1TeBsUs9+6oRscQgrIJ2vMeXb/wzXTCo9J6Gy
ovvPfmgjnZzzdMp5hUBWGclQ8oop9inofJysVLrJqR2/ikR51VRqC+AHkhQ5DzA2
a7p3LrSIajHD0MVyMM7TmdleEqBAac2wsZyIm83ZwaZscGxLBmX+JU+qI7yTD4Xj
ntfWvL1b1dPMb4dJUOvQoKqZJ3aST8xEYi+tNEzV322LsC3PyojGR/RNJrBJxQZ4
JKaq2+oWaSd8MqI4YY+9YFFWNuBPEGkFgY5KSC6KC5nB2zKo6JPZEHooxCUGcVP1
L0V9fXwWGEONpqkMetSVXLd6U/oaGNqdHI3ZKaIqqxPcvHMncNu38oOrMOZK6zV3
NbSmjtFSgmTM+vAPmfGn5DwY9e/zlOsSVJAR2eHISd5U7i5ylCNsFViUi5+gHGRK
VL2QgkMMyegvu3vxDu7HMs13X2T/q0op+peWiO/BZmikSYQF1vh65/VHRVsh3OqL
rySexZ/8v8+CzMCAyyLPWu+mQNFW/gbFoo9pFYq84+qTqSVFLiAD6rM2vkJl93QX
CV/ZRETOU3JOLu1tq7vw8nFWdmT4YNWitPi6n9/z0g0NAquGi6LZjPB7Xis3tC7Q
2AEtiO0Utj2L0TqIdTREmKUh/qH6nmUzrFrccqyimcUH1px941U0rcGh8kP65IuL
NnWubnTVkEbUK2xU8cflcIYxgkfTHjFPjzhxxaXPRBfH4f1ur/l6MWBB6QdLCGZb
iW+pT+x1WzF8QPTzcc1mxSK06fXnwhLoE1Sp5eXiHbMeLAEWm7++cz2Bv1sy2lrW
dfaFyG5WqwFem2HBQZu4TDQ30bZGPwf2TD+zosVN6+z+7bsHYDtLXozmfZhwTcaa
I/pwVaEHGApEzeZuWzCxPQzgkzjGuJC0J8F91rn8RuovkgyZcl7bYVH66k6z8Y5e
12ii5IHGpBr/sNYpcW+gP5CMRhtOnnEIjavwuyDxS5/yTZNgJUgS+htIR65mUAO2
fHCZZmBvmj1EtiOH6OCwjQZo/Zz4kSt2CzPzZWuSQGfkqU+xDhCB58l5vgy8mNKX
yguCsUWd/q55TA80TJL9WT22DM9xtEVtzYt2934XiI23QGMYQDALon8kYC9Nux5v
EZCGmXX5zij2GUEyJQ70CMdniMqpTfUsxFd4QAzH9CU++V3T3Ao1xLpOL+uTy2es
aTgYRbOjB03b++f3qYL6XVJqVmlqCtGxly7cRp/xnpAuhyw1ERQBU6KkZwsa9Rzq
UoLmnaBk7yjyV02gLtTNwhBdW6Ej9o0E5bp8elo2aI4MkSs3FDGd+kq2AN3VNfUr
fPpK9fkF20sfL3XFkqgNRrjJA6QUTCKTfXGydA+kLjaYbm2g8iOvy6e22uHjsJuZ
XCCVkH60q8bObPfa5b2h8qOBInhQ0a6uUFnHKuDsRdfSlQkOMudPc8MJtpYe/X5h
T5OjDCT1CUb5D+m3rki5mYkObTiELSElfaMpdojofXbwpubijiFr/n94lodYv6RZ
aHGpdzY6cgFrUeNgBea+EUQk6x4MwqrnWjwt+FJj1dZvOwW25QR14FXIZNuvijMd
i6kFDsIxhogdxTKzW/HNJ/raG0YbE0k4QdIxxt2EA1uM/SBSL8pllBGcGMPXZLVU
KuAmesbmZFylXfT6AmdUvN34YPu+g+WsaecPlHlNqcNfGLcJ8QysTV2Kiquf91eW
+IYNMpOF0A1kGOe4NDd3IUN0//n7UUJpGExkSlZKjs/ED7ZX07NztPAbtxcQLcwX
hVcV1Sh0VfFtRwKXe8rRR2VoYIFJmLL93HruQ2FQqBbpbc+1m/D9IqLRUu0ZxOep
WYYn64vWkZZyw+kXTLb0xMGxkwXx0Z+zy6CyFHbrk9g8NAxFsEpOlsqnnTk9A19+
1zVvdFpT5IE1j3O/o+Fh5T17AKa/G7NTlRoG1JcRQCfSbLnvMojiU2AbycOiaJFY
iHbjKHg6ppVvieJTliRoQtu5RmClUJ/xUYzxuDu0sKd9Ecg/3rUN2CndmMXaPhDT
O3oHmbzFGTWpvwdEUs+xHm5qeYaVR4AIQKPSc7hq5wudnPcws0AoKzJ6fvdGGbC6
vPHVz9V7anXRy3rNW3xM0GIyHIIo/OirVTSPdS4iOuw01H62PBT15PK7tv2k5rtr
2ZervEg5z2UNQKpOu+k7/LXvWbl25pMTU8R0AWSC6eukJIYA6H8iRF2uYAtE6w40
tfItH4P1XmDs71aSkmAdV9EEC23rxCqqvKiqtErcUEI6sK2+K3lAQLLZu33fvqvP
2yo3hht+I3NqM4f7xJuW0DKJhC6tN6cLEJE7eORDJ2mjNOmlA5tqSvWBgSyGlOUI
tWt5V5x1GX7oVHpf7EH622yTHlSVoXdtIDMY4wq4RkhyhzHyW8u6RFXYzQPoGWYU
JoboedgvDLEHrfuxkUX4uIgrpk9S4G50+RdAX+tM/1SiZU6jKEC9pfEAfTpU/OdE
M+JlHwZWk1wKxdcqAIB1wmGZZ8VUPJASIfCZAM6snQq6reXL0KOZ2I54LrFmONvr
wDdb+B2u0/meZZeMk9bJv5hvdGbCC6R5DqzWO6/fvug4/yKsCRQ2VaEKVJ+OlptY
gs6rCP/VzOG3MjQAyhW1QB2hs5Qx7RkQetw/p/VKcyn4U8XO5urtI+Pqo8f83Sos
rv8E4ebcL70zVzXZI1buY+XoqpGGIvtYF4zXaFqQ6eSu35YtXi+6CxdSqeRwaw+1
B2l51w+uz13GOt2kwP9w0Cf3Q8CIRdwPOHAHUzVtUbYlRBOXYYMClWXlC/M+3Apm
bVJPeN2hD5w8ALllxIcgjuBuJ9a7LnMCECeI/cqf083JH6PLyT4kWTkYWPSjLx2b
evzSsHN/FEmYAX6G2vdsJ2NScbRWINeQSNgQzRlnDkLMt2a206d0vQuzmLJbfO9I
v7n1llPNypPhPPQP2gs1pWJGYm4xFIj3EwwgTlu58dAB/dBUBZeqczHjZVFjzyfo
pDgnTyTHFo2dbp9Hw5+08GRts3pRr8yKk/xjEZNRUUq33Sb66phTTMLS4OXBiGKM
oxeXpOYOaAbe/KvHCrVVIdciFcl5MGE3XUW4Q1XtQCjEPrsmxYAf0QTBTRUJu2Uw
7hy8Wi2cvlqAyWd17y6QQ230/l0GZrdfjs8jUiE/UtMQBTO5eMV1THGEaSINE1Q+
h7rAk0Uc47SnBslCnhm+waW8VjEmsWwStFPhxEMWE02dhVB5sa8vHwJH5SRy2PcQ
i5YpXq6W5SAM301TWy2w2vQJGarfYtW5/pBbaTaLSB+gTLzS9kQjp8q3OI5pazNr
aPawr1JfromjMrO+ZqpYEBfwf7Xm3CatBHAJ/BA+HdB6Fv0AXKX4qlGhXjMCPNd6
BxKeUyk3QPD6ZEaIou38LMW54p0RSSX5LTxwt8ckD8e4PZc8Bh/0v2iAL4spjLss
/goqUBzMq0V0IylA8L4PeZAlZOFm4f9sUUjj8BpyKn+ML5MUg1gLPnz8KsPldGvp
cZTC7YD+ToJalErLw95z9ojM73feGOZZPPevYSNf0qhjG1yXwl0j72b1N+mOSL17
G295n9+YG71atGWlyAsvKQ2ujAOX82Ql2NgXRVFJxzqNpmisl3roy1AD/kWGY91/
PWl5WEOGGS24HUk/Vww474qo0EDEICF8TbLW4XIA8kVzPkJEDqtEA2D9qphTVK+V
xAkhMnK4pmt6chH5Tn6/LcfQ+S1kfmBLWsSlfgCEY76OY4Ngj+I0DajGhC5763QV
LsAiCY4G7WnRt4cPT3u9GuJq86xuk8kXe78eL2g+xh7WopqZ1I9fUxHJaRjkoDzZ
CQ0r1snSrnheH4DcWkOVpSVB5kq5xqB9NE3tk13uatiMkU30UTyKbt012l79rm8D
DBqra2YuZ8uPxsrvG/24SqF6Tgsv3AbP1qKcCDphQFgfsSOT36A9F3imAn8Bg9Dw
hy1bkfcb4IU+Hn6b/IqqG/WcE1UjwLkMHIbLXg7rgl7J1PVBm+IonHXMWV/J38xn
gjIp+o1dPg08nfTt29i4vogABlFYA23fk5PZ/QBGFV92y9QMdLKvY8y3yeRaUtOV
s9YV12NlvKS+5urIhn59+d7tS5169z8HvlmoS1wymgQTqHa24zyY7yDSxj87g6Uu
hXHBkcf8loLmqG6cs70dx2+QOxZGndjZpL66b4crHboCPNTRWTYc2z7v5Og7F7Ex
uv0AFLRyusV0UPeqAcWTms+wK5qxpvHqibRofHqivVU7qtj3U2T0qY7103/aNf4T
Wx3MTuRb96vxb4Vo6ZENyOpKF7z6M/3xQaPicZZDdOKlXSe6cnMjTdAHk0mK4mGo
/A1wlsqxZg60QsKoBVX2K3Nwzia8gH4YDbgk4460fWU=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
I261BiEKOyZ14zGgqbK6wUpnuEIOi/ezJiGibnCIOhxoxRhGxBCEEAeJk2T3QRQO
Tg7U5MyGJwgdR2gjZ/uXGrnuMEPoYeVk4r8KoH6tD8Krcx7ltHEnluN+7NchJvIG
X2CRZOb8bgxiTInckMyLMCRlSMW1PPlVaOvoE1BdBJ5NFmb2rUaABBYsOfpeecHN
3m3gz/5D4kb6EMzvwuFxlQVZ9DUzNPfxaCUKxUDljQRfrVnFbQj8kET8v7phDvy2
fqab8+6302rU9pNRxGj1c6s4OaQy7zeBfRRAxQj7YUtK7mWmRQmlgi7vgDY+L1L3
bgyTWUTqjiLv6ouEvhTcLQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 20288 )
`pragma protect data_block
exJgMhAk8m7YfZAv6rev44KgumvEUD+uKcqPaNIfLCFlqcLFBI+4BA2I/CkSpg8H
y6HjUyIjfllfLFBTQACwdhRIGV3wsnWUxNzGZlqqijulb/7/65RRjyu1F8eSH+K2
5DlwSjvsGpiiKXWzUm9CqEZG9ziJFn7E+Lc+HpKRKS1FM0bOA4VE7Y26CORYY8PZ
6ZwBsflURazGjxThdDxy+VWC05RKelX4vjRdSMo8ZAYhuczlfqfcijJ+QUrdihml
3C0vyuNSokt950yngI6AEJ7sGhxyZxBa41Uxg1lbBB5ueTRZp5Rqmq3TQf4GGLkS
3DPiPlWTX2AMTrx+Arki0NtuvZGf7262m6/bKQVnT4iu6PrPxIqyArV9OaRZmFhQ
mNOg9qulubeimEeORwBzW0LLmp7OPLvRAvrQlDBwWMlrlvga7/sbcEKnNfdTUZO1
+NGfcPKDuY6XkWtJ2AkQ0CKVNsnRn/8Mvproo8A7/caLfUC9OyK4rlVqSj7miarP
LQcW17D9XMETdJwDXwjsniw9MZy7SlVX9mxDbiHdwNb3MN1LYPZ+cGvJkAlfPGSH
TyiOlQCGJk1ixmDcRZOdL9G+YRdSXOVdYiKuBXcdbu6UMt59lj55rNtZ1dh5C2pk
snqS+aUfhXYz1onfv5qZ4ZeJ1ze5mq84FBt7uN1pJDTz2jdw/gE4Gx2qgXvcUhBs
hF6IfhChLM8dV2ERk3tmqRh5HCRrmIAbl4rMBq/HKnFX7KdiWQgxKmZNAQPNLQZ+
hXgG0nn3tVw86wq9D6jTCS85R7l1GIGzqdng8L+hu6FZwUrWzv7BdbHcgsXWJU9A
SbZ65mCsOVkX5MTnm6xBrtmKTNYiF3dayHCq03Un0Qw5cyme58N3KsID0xAPK/fV
PIoWjWp3CIML5x4AAS6NIt3EN+H6sil3lPtsjejMRu44vy9ssLozga4QuS3wqnKP
CWgVyjAK+pqEkDmR8rHR9G+lfuwoBXRIrPjZ+xyVb2eYObkzL0PltTuWniknwPEi
PpWs3ZhmTby1os96D36j9SqDHjVy3fgHLF0sYFtHJm4e9wgqqKeweIAM4tCb4EX5
lerjdOeVMMAW60JF5FadYLQ2NEtqKi3bbhdHLQHmffCJBtR1riJF/mJdS1OM0HLz
Yhp8Zmbp9gkljMmHK7vYMCmlWXU6kh5vwTo/gVVN5EXgDHFumcFTFiTfED4YcKbq
PevCJ4t6MB8cARWwEnlHCVezzRZ5uQQDoap+jMhv5Tyjtk9+tAXsjXNWtdmyHLRQ
T4pD5fPKSsL7Gh1BOndE/vkoTHyzb7VtRAloPoEOsHC9XEmEbdMJ2LaoeekBKbUp
oSWm2yNjkILTQO7STeHGRlor/3hOtD//zmQ1lhrbCFlYHhYM413imvbOG5kDizot
hw5hB8gKXWeDzUwq2Qsp7hRchzlHpY12kxsIik46QBFxoNBM22dsSB5bju0KRNOP
5RGSoV5jJuN9Dq9nRgoxvs4MG1n1zSLKLHZHfVL7/PJevIN9T82bqcRfvWnN6cdx
4pDJyZKeRJZ4KMoDZf5HOeLaCJT68OsuGMbiXGKLGSy5pJ1CkoiR04lA16UN9BZk
cv+mODszWXTEqNRZ3w2OqMjco+IiYxeIh/VGUOdRMqjWp3sf2OnM4vCyH1VnNkPm
YUKigCaNMWIlP5FJxxbLYz2cpIIR8+rXl9pmaazLafK2xe9JfuXXnMTo6DpOwCFt
y8wZlAhQx6nWWTUTzCGE0z85PV5d2g+ijEwXoUy4m07zyYxgMtCUyiv2ERfneABG
NnLstXEKD1Y44Il1FwdYmnQsZGkahpsafGLO8nJ975hOQCN6wn66dvXde03cGanE
wK9gAIqIKoSeXEeTjXhRzRhQtPDBrRrDJO1yE7l+Xp8u6g4xI+9xM/iYNAUarkPv
U9jkn6WJDRdXkpohv2OWk91mDW1MHRbdcI3xyEzEpAD7m9sxyfKgsrDZ4Wt/Mc2B
GnIUK/DCU80XhfD3fQxTaqeRlQ123Sq3HFcwc3a6xCLUobGbIKBSMVdrSra411v9
F8e3qPoPFxjB8BWmIyj2SgkfbGkmfQRrRFIOLREHuJlvmlxyI76gj1zP8ieZ6M3L
NpXA/y4VFSBNMy1Lg+MEUUWVGvGMp6HqmzG0flpwB2S80qRAnXnH4DHbmvdWK5c/
3Wo0XclUbA/mrlmAPE50ymQdpfOzFU0W7H6r6h9wwJMH1//UjsJIHcUyRAqzP6qs
LS7b+YkH5TmpfFvVC0HLuJrIkzNk8EeNP316TH6DLepxdJeOeS0mtTR/EyfvSSxF
s5p963+FcJyKE+90oGHCdTUmDZonhgX1xk0HO5ohjrkEKOEvYXq4b0ZYUGGWC7HC
p3ngvg1Royiw9F/Hcbjs48LRfJlUwKWrn20PmWwWb3xCBOzaJZtE/RhntCACmXXt
uwMZ0BUHuYF9iI2UKQ/btfDOYWsBWCTebed+VCahvEfJ+9RUnRnpcQy8r5zEUIfn
fYqvAhfOPh9RU9oXSRNICS/d7ZJ+w9cv98F1pwTSCRRhF0JgRz10P4/oLpx6Uxof
eBcgLsMu4hwNjvkylqSvLdXYEDyqsgw+o5SxYWzBFtcfQnudVdsCol0dIiNvNVdx
fyOfZYmV5bajh4YOH32Powfq+qjaRAHHMggB+VqVtIvwBQaYbfqZNNY5D6H9Cyaj
nRFDxfTxxirQv4POC17ZV49O10NAEZupAAFXLcqxnrtvEwLzvKOwmmGCQSg3cvcO
K+CdcOMTju0WHcp0ETSjyuq5DaFi+//b57C1uwUIEjeOHsgz/v+FPofBBjbjRU4O
ZuDhkX38oEz6n0ogNgWt3FZDG6sFpNBKqGG6fhZafA6K2kTAkk9AXKak8qfWbvYW
E7h2tuh45eFN5Eh6Gdwfc5Nw2HWiaoRsrvzFYc9/K9QNBMWNSQzl5qa22Rekfi3Y
5c5ptvNjrlX+WPvAasuadmFd6CEtXfz3tlOu7B8aj5wr2FGuhc2Ik7bgrkYbn4dd
7edXJr5AQ+haMIIxQgXBn6KXEsxeSMCS+jyozIjCbZ3Vx6bFfAr0tLRPyGTfVgGc
He75ntP/Ubl4f61O+vG3yRl+0o09FwVmgyBoKkwQriG3oX866CzKGuzKd/9Uxde9
L2Nu+4MtvnvAycLahjDf7/YKq7MwE/y8WcS5NoxNrKdjCmUyqoYwVBHdctFvlOxl
1g4DhLiW2YBRzdGEu5U/zz4/S1MAQDCX4BIfWe0rK0y724kqBklSysCWpyj/0+k+
n8EzUvVXBLgXFboQVRcRBDW4oM82ovBy+XsFoROCzDa3ITkz19VWMWP9Qq97WHKJ
3WRLvZZez4+KVCL8plNOKdvaqmVH9dywiJPvKIfdYUadU7EsgCkNOz+oVffSpDHZ
+SFkR+l5gmDXL+V2u5t+epCk17RsrTZno9k5hRQfBGHiZ2WruWRjbh6EveJFW2Qo
HZSntuataSoiu0ShzobOueuGGx7Bv8VxmjEryXGNI1I0yL0fjxUXhEev0gpGf5+D
1u8j9h15cciVlCdx22W47iFNUgQcYnWLV3fF60uUa5iScifRP4RtwjdaboyLmIPh
EANQc+4PiToUOYS0DJaFISqHazJeR0XhQlnHSsV6bIkUsURhvtBSxl0nG7wnrw+n
M4NqlbjRhiUv+XBYqOkwUxb6W4QHgkPPu3SQKKsV6ZI+v8qkfGB4oWXpE3Vvo5RG
evN3DC73pb1W8tgpcvhiI1bsJ1Z50elwp4VmApFl1nBQiJkHioafTIgJ7FHkcRl2
IYeVroVrIATJE3BysdC+ziQTaHTHBxm1U+ezfSvvlvUB5pt6Dgk71pg2uloc4GP5
iafmv4gj5izEJ260eLIDe6qNu492tSG0uOmDuNH3S8CAfz5rt8Rrd3oKqDMgwJ93
NYOTEsWXUwOMLvGb9B8BWAjZSkMLSmKJqyLcyUyYRTBD1YSV4bE+ChfAX7ltzkaK
auF75rDOXxT9TrowqNYuHCSuhK4eOGKpA0/HuCqjsMnF8X+Q2gkvkiRjEyQpZ0et
X8rOuTaLh/sDcl+yR0fjD7FmCn+7RkRkmNDk2vObb6+Hi+csEytIkt3fTC7ET9xA
H87CpJjOAY2NnsBOgp9PuqdZI6Whz7J7bBKQZr0cLeePsLnAf/liDeam9xcxhxjM
Y6mRbI4dA4RFoANDeW0p1G1rMi4gFZ34JrAi/dx8mJYF6VwqDST1fHsulzMrxAJC
/qruSdfF45fvY4XNBU8wHUjF6APwBboLCQ56towFhY1Iz4a3OtfRcu6Lr3RH1Ffx
ucyERqfdV/ivz7wucLzwoIYLyuq7jTn9/RTmy21LAYTwDRFkGez3c0h2ZPaeqw2f
GJxY6BppoMVNngEjSMh7SWmXcSyAXmqqlNc3na1u+oqcHAAZAYkSGd4Rs8JLaol1
Z+oVfckkPtpvn/KvatqH/cqYnrKtmzUavoDG4tNoh7EJCnR043H69ZfB2RSByjUb
u616BTJGlL6VBNBtX8/8sokDRMeYftmtnlvHf1AoD4S9oHNU2Sj4U+MMG4EJIE2K
pJ7j/hnMRtrIut5b9wHNTwd7iYNqDv2WMAX3pY24LCvONwB0ca+9DWRHSyES2Ty4
5H1iJpiePejc6/n2fpTzhPM8Sgg1WE48vTRGGCopB2jbBeRJ7vukyuD2+zryef6s
vgk9IW4s1KJRhyF02Sx/CzL/m78TkwDQGPiBKlbjxU+Oz0egNBepLTr/05YH0cGm
N95qKrKOktdE9Ic9+S+0FW7yXWEG4LS3ocaXUokF5kf40TS2HDLCBXSaceSf2V/5
qXqvMZtRUGa2YTkWfarBIWy3sPsAs1oY3dkOCh69XUAN+VJvhdoeyGVh6FV+tiuq
0dVOzJrH/kxnImaN00bki+4KkKZEVeBD3Esx85lMIrsry79eWtvn0oDpRfE7i6a3
Ymg4eNwE4IMknWmBwHJ3I/j/C0RYbv3+sseLSv2pjOB4NjiiZ/n5A9gWScDa96jx
ujYeQigH+erPUwLbi3PSx8mik7pTVVIa/SyW9Ge9H3ygUk9H3n5v9YAnPiXZRxV4
ESIdnF5xcYQWrNMDOIajfcDxdb+0AfkBKl1GPmtOPuJ90+WU+hBtxbML3GAsrRjF
w/YrEj+GAi6ISPJpb+LnwxdpQQoi5OEVXjWgcTGbOBx+r/k1wuygfvq1gsY1H8dY
g7qrCRVvh2pI3/8DilK5u24LMq0Ul0RZpRDsa3g2S37LflyQX2DdbnK2vm/WscgB
91micVpYyQKUechI+bKa/dXeSUisCYr8GMWdwdqNklhI+t+1QSvlZ5eMUEQ7VaaJ
NHTAYTX+PPauBjlOTvplrMt/bGH3UDTidqDNY7pRj6r8W7MqVY7uTnKADwj7Tf6z
MLUStv+W8YDYcINAmph5WlTAML1wNGKBQiEVaBzgJFjOtCSavws4uUhhrKoacPw0
4yru70jfbM15kJlkzMEDy7hI6OxSImegTSOmxvV1UBjK1GEZlNFQClwh5di7UlQc
ois5NdxciuuvVNSSGZt2gnXfHb+fEtvZYYfkuKIdDRKx5HYN1gm7jdTTc/gzcl26
pZc9SRrV70EqaIOOoOJUOLUJs4xFwSqurvyGgT/pTaN+FzASuFz3pO1DV4inYUEi
oPaFJiDz2WEpmPq6uKVlUyKWW33gZ/HP9AyEwwmN3W7QH7QMh/XWIV8PEOmqclSX
DUs9R3ipAhkeVOioLykOcVr1oacPHKDEjDtQX3AhWRvr6pFTwmyE0d7a/BNDGft7
Ahy2dU+9VeO0ZGbGiCvd5EmO+qo6MfZK7xmdq7Nhc9tZZcQJO/r7RACbFLVPvnXX
oYXcwHrTuljMxXFclA8ARNK11/qZQHB/CP6qvWqqvkPArIiToZj2AMSqvQAN40oy
Tc0QkLKEHwvHtvkMD0+cPkiyqTDbC9wSwEMEovAR8UNLveGAbbeu346Y6CNfICEG
tO+m1FmUixW+0gDmFECFa4I/jiBBbj4zPhUpUu1pfjUHIq2n8UzK91xu4w22mIjo
vv0gPclR3w4xpGXvuqgU+HBNOuwYCD3U2NfgZ1RCBZ94Sw5iYnpix9wTofkloenV
1tz1i4t0VQDmLujDZ8SaqV73Aw2jL/uarAPN/QJ/HvblnIMII/kIQxXcVF5MrHIe
dMcHXdNrs2Lw834JjIifTNapXlL3DlqxJdWWzSFYf/0TFposuixvSOrBTtgYd+U9
zniXOPxtJkAuUNEH5b2Dqljkm/Ur7UgqmcSlVqjrFn9m6tHPZxyxP3gQleMVFrHE
k3ghZa7NQ1MvAkwBurMfO7xmZaMvlIn3LNQsGcrZ8F8d/mjiBaMpxEAgehAWWStK
jbwpnjKxoUFNjMCZJmEx9DnKHUa2nnS+hP9880b3cNWiNKT0ZldpUh3mhoAjp3Ox
KFzmn5Lu2V9Epypmil6LmhMBXIXQLllD8sgUOrdyjwy4suKZh7EdGuvfMBYv5ByS
tf9Z6ZM54lmd9VpihZ2cpZltTeTlGTdjx1xEvA/CBbBnNaF0paaS2NlEODhL/TyQ
WbTMDgz98a8EZkVvKtMsGHVT5X5fXgVcff5frEU52mPVoAJLVmOx+Gm0xpGR45tk
WLi6UXckCZVopb6p8v745jEkIp+fQ71y4oy6VaKzb0rubCNVBXcjzLiaT8E01Ano
nGSgfH9iGmH8KlPD/SVn44Wz5hL/xAplsIFhh08Q95w/8MTUGX8bcc7U9g/T2Veo
HmMuM9TnP+cfU0oq048FRaAKAxW4DHTmJI4UL6+Q2fSIKPFqK0uU3Ykf+aUSY+aI
M4CEzDHSSldfX7vEge5mR89llwAggq0pD3I4z1y6NjAiYAGp+tVJapKH9b3HHwBJ
WFo0SEFpSMypRs6PbJA6/Crrw9F2E0dbDBSeZF1OYsJfHlo6p+5+zbb9ZUg2PP/C
hC+zaEa2njL+KgggQzizlH55v5bfUO/N5KeImcYLsIlO2Z226CiNN5wEM4XIGQtc
NpzG5wbDDl5E61i0TkAYzomFtwS5j9NeS1lyv8J+ol2SAFeG1Db1hoDDWJok1pQh
iUi1cz3CLQLgFCBXfhbQ91J2cpth9Av6gx79oRRjiyCRyIlXPk1j43bkapdaMEq/
k92wc3zpmrDG2SDMuwkP8nqqJ4rSVIP9TFMSZYwAKiGavxVLILNM5VBTxxQ3j/QS
MX3f7s2C7LO278457pQLC/EAdNYjZoTSiU61MGwfkHtZmfT3rJSRBb1t0aIeGR0j
DY92CvU5ICY6E+rzhwAexziJJiiZyj0ZCNdPrCFTxuR//Ttgl20UJ15rj7CE0RWU
ZhKsUoMgGUknhEt7+thXbq4shK+E1jCNbOvQJ08QHKvqZ6sbXlV51Uo4HoE/2NRU
EDSn4NaYbvOFvCtzMnPEqZ3/Vvd1VOFKXcfMxLGqQmeuq/8I34PGd6TFFzeeWxl0
Wb0F1+PzHPKTk8I5BRipCvvh7a1YWYb4ufWAvByLF9mnGFR9TE0g21scmwiwr4sx
9eJr/tzg2s/S/N9qNgkI6K0J01qeaPIwAgF1fZJKZyQM2tKmVEkPhzguf96ztN7l
Y0CMR32LAB1f3QDzLwdUhdRtBSMq2TQ/6CNGrybJ2FFFQDkMPBJCaargebgoji0K
r3knJFIy1l4Nap3qh7NNjE1G3jFsx09lI7kZ3OZxshpDzb9F9JKT7lrtR6eLpMzG
dlHbNdVmpVbkmr54r/UTPUnZr+P/6kSDrwP6fRVwuPMTT8cQoqRS2/khL7apSRqk
tXqWpnOsc9L9gLRQaFLYvZtpijEgF/08JuHS9heq4UJgd6kUyYUVqLVKbNBDvHox
nPW6D6/CZCqvVHc4quQ0s8vOcZ+TybtC+I3eLR+QZnU+kLm5w8GJLjkdh6ie1zic
bKyCoHRLbct+YbWW0kktIzWOnDq0YEK0D4hlzA0AcSWKshpZTQBugaB6jfrkKgD1
zgwXYfeluLep0B6WEL5Ae08hESNEjsk9gmcVhAZ0pSdEfY/iwfr8sOz0Y7PdboZv
Vc6Pq20nqpP0OykZZGnzcM8GFYBqqbwAR3xvuYPX8QIeK9Sdr941Io2Amg2qpuL0
QpV3Z3zLkj5MJMM76V7pQk4mfDBClWzAnPJthEC8SQ5U0BS6wx9FtIdjPVCaTXya
zFwJftjOfEsVxktdE7+d6GC85E8rNU7fCUqKJ3FEFkP3E/FVJNXocQFZOF1Pc5lj
8zmcGdPUAspA91/dft+bdHp8h8HUElPlmEW8vcfbsvgAFMjd5leMCJttDS2DTSqo
Dx8PpJTnYchEqci0eRQxKr2XReQLm8Bvteosgj/SzrZUAXegqUUYTI/WccjDWJuV
Tkxv1vCV7SBrwSU/M03e8y7DGfc/kYqXwh/LKkrPKjy+7kJdcHxOf/QqKFpBA5Ky
QrJB2Bc6yEOqzobYqklZHQe4I7VJTZl0EqJoUJmHJzEtCl6EmqA54f/XtOfx3Lms
Kc2pPj++xnwxm16hNB/K18+8Wp1rgyqJOlI50Fic5XHBai3QYXxSN7zUIQmkctw+
8YbszOFi/7/vx4+11wlJccN0zPRMRlOswvA22a9SBF41/nmvtaTyL2ZT1UVG89nj
4q96fMALwQmhPCSguEwdyghpBC4lXAwiGlY40nBCJ6GdMnxa5diCMat3KmyVIHQZ
orRg/HD9OvVTtQj/sNTQFNhkCcFg04lWXLKZ5cofqpiKA2DNAjU6F5vS4RQPpMXa
GntoBsYgsEgvnHIuuZNYAVEHBxI0QcL8zVsDXS+bGkiqAjStuu/kmtfuvFIZNUJ7
AHv8V5ZFnrphzQ0rXhCuSRFHo1Dr9o0NKEvQIMO5zMOlQOuvzECk3ITkUgIxx8lG
92aQ7o4SLFe4vr88m4cdGBwLNCjLkHKritDKKe+AJ1AepI579RDahO03QaQZMgEd
mSJPacAzSTp7neUmzhtSxhDTSsoLWIQ/axrIAE1AvRdv1weeT7y2/6Ls7gkghxzU
HxtZBzCpHqtFOvesOM9I9cd2YVvgais7M+9tg21uKAylrfNAR+52y70TFqFDWt7r
XBVIRRXDp7nkUdDXTxaeyE9C1Qs8XhLOlag4U+koX5xaaGnTYJr8tXAnblbPh11r
TK9fD630ISOKdmglH7iRgCRrJ/kZybuLYCXUG1iL+VWoMc/4n8fG926Vb2YXulRn
FvQpfs3as+1+1zrvjtJYpUX1mn1IBFRQgSGKR83I2Qw++qQYlul7qg3UGvVzzkj8
/HQDpcj3NsWmxG46aLTH/gBukUDlamyPlaqRZbc5FBfykkbYPZit9m+YKkwVIpkt
mkAUd0hrgSqHcAK4Lfe0ukSCmiKzE6RsD0EKY4fO2qTv77K4gLgsqRBBOG2FG5WP
bSHVCJZvyMs+vL0gyeX3pKwk/rEIXjCYkDwhgSJ01+cptkRZO3VqhBj3A5UgXaat
OI4Q/OtnofgxXdcyUnwjcb5RlDX4DFEpC1p500wNhsV9ZFWMPoXF3isUz/AYSWPH
uBToRTQWrjBHQVAA5gv0pNkWp8C5HjpCNfCxI9x1Z0LrYC+Cqvz3wQeDKgVv/S2e
zRmAEvGltEedY32RmeaF/SnKfCKeTmUfcftEQOGQO4Tuaa0mt/WgcMuHl4Ma+v+4
6rxK2c7a5pGS7DDZGSwnMy8PkdIlKppl8lEom121Oi5ImOMf2IUg3f9Zg78vLeP9
qPufL81d65ecaWrdl4gDSBcge83/WMuM7aBOHUU+iJ/xYxXmste1iY95tsIbP6Ga
x/UEVelDm+N+DTD3QkhWfLdqBK420wX5OgQX2dBQQxMcNRtlRT1DK5HMyYjRkWay
FxPupSHP7ako2kYH3A8IPN9gVfGbkulae7gEDZe2HBsQqNGxeUQA2Z0GjGLepUEW
7D1o8z8ptVbAsyYc53koZW/33noAkUtJmDMDDrCNew6bx1Ufwo4bYLNM2+j8cudr
BAzvGv6W9GnlLMABXhlGbxFRL2aoZNTUEuAGDqzAnUP4BzunitlLjTwdHRZSw7Sn
rrh1/RtBpeSu1uIdbQQ/VLjMcB5FWVbI2/JOEaYeGrH2/fbvYA7PlsGSvdYMCjda
Kue8Ugfxtt8bK6m+L5pS+8eB6Tx0hi5XiSV+/PdQpQdZINVsApFeVlosJEmqRHNi
Lbjflwp9/ab4AlR0m0Qd1qFduT8iTavwEm/yFP5b440U5lc9ZdQOAaVIqd8ymGIk
87BaOOQE/U4zw+57+80vylAh0QSPvHjG3s94sFckGo7RlxSw0LJBXBYPmEmQ4Tv8
82J3o22hNrCwO9LYpk/3oelq28LGvOdBXtBfv3uJwIiKeKf+DmQIkcT7CoCDafyE
hL4tkU5E9IgRsDWgomFeviulScpWsZV8sr5lQTOaEqOPjOkxQ2sF8w9HLKOBL4eF
jElBm1nJck1uBX6/Ihrsqe3GVhnYCHe7vGKLp79jhnaMHmVGyM/uAMZioklCqpRJ
sFMkGwvIEh6/JlIPmdAEyoPwrE49UCnM94KtBuUrKfKnoJTcv+aE2UJfO0nUV+nk
lvm8WhuzKsvV8QNcPcGZYRSaWrIMnla/tiDs0LDoG0PcHa5Yd2P9jOXMxG/2TMZX
/d+Hoxbpm/zXn3eiB6OmlPFuuWpgAhN9pzb0m68ctwOB2RZT4alGbxrboeNHICFD
umN9ECMFrTygDWXr9W8YJT8/VwLYEuqSTcPxwwIkE0j0VhgubNAxD2y5OtSzlK38
LW9TorskYsT+j7pLwpZ+JCDdBMkwmwpAve8xKg0FDl6cryowvd7Wqi8d7lR/w5j5
Rt3PfYWAAedfo/E9J+MC6jQQ6j575BlW84/y4Fwl+0xEi9DsbtoLPxSw0Lu7rCzK
85mNeoGPInkfAOPx4Qei11yEmpTk7DqB8kLqrJ1lWf5ZwlD+ApbnDIv+bGhPmp+E
y/51B60nGs3NYZphuJn5y3BcZ+voSi6SF7okVfca8fo001uB5mBv1SswD83lAqUK
6hzh7fVnNL9AgQC6azQzXFFz5P7bghm4M2KaqhCGVwpaZ4OwymbDWnzpPC4Nz23E
vE2c7ih5gu45sen+7iHGA9HqzSaYs+kHUT71BLhJmxzsbbm8v2t4VvKw9bjLobQP
HfkNtC3cFcfDddUJugL26TzvhHra6IfkQVmG9+HNa/W9VRR27hGw83D1aK54HHP6
S7yD7SUqO7Yb1Yyh8bJIZTM0RivrxWUxmTjd8UuEoetx6VhwNKxlJZ8OVgiyeV/P
fdGNy+mSAUNeTXXx9n8b4AxTbvUFEZhM23dTUNSFXQ8/mJcxnWSfQviy1FJjvMEz
KrbIyCeYGUdeZZpUhjuuBE7EkucMZdcqgrsJR96FP/uoG9fiYO6V0iZ0BtWHHiHV
WQATlqydeQGna7Nw4qT8Ump41ebn9KG1fx8mja8P3VWoBjCrn+6NY/AAAQP0k72F
xtBLeOp+0755zGKr5XNHzCmJ8DbokNl9lXrjT2Fv9cwIpD/OJTXnDssLjbQTkf6E
wUGkQARlktZJZvXCVX3eRB/6Fx93oQoJ+pdbRb2BGrv+jRy81mWcyyluaHcj4HZN
uMgkEmaTzfo0PYBZwzXFK5/hU+XBb5B6fglyv4Esl87T74/xfviFirVg5Fnyfq+t
iRTNjVDKpJU6oNoOq/OFeIOgUApqggDPebuZ70B4rE8FjnY7ZDPbAeahIrColrIR
Sij4l1e3V0mfrwW0wJVrJZ8DRhKZlZ0grkvrc6qQfBoPq+I3QuJf91h5Y32t+Xrf
TmZIDEAP/ru4IRzqjcR5LHoNYHJx1fy6Hlg5JNkf710+acpfJmZnTdvtdz5OUSkX
GRaP9nRvLWnRERae1xydGurIZoRKli/XeZVx2wo/0hOcy8XJIPyiolYtgMxIAOpw
7hJ1MKvaWn77ku7K3ywXXASwNq59xLeGbsKoEcUOYPUSp+zSEjVXv7MxhltPEuL+
JP1XzO9vcPf/taZXZHTfxeuEwCpn2sukYNMi61/4TH/Af0XXMgLFXVXvVynJGD7E
ceftEb2yA5d7UBYl4WmGq4O8k3qGgqn5wpI4reW6Vx2TfjxUhHpp8DJxPqSdHmQr
BDFg6oIDhae6Fg4qDIOQEQ3ZzaGwnvKoKb2kXbe053d6S5Swep5lErXb/eH6Zx5r
mHmoew6D1XcgwhQ1PzxWsORC2ZD+ttJ0lxG+J/6iZsWa8w8E+PubgcLnMqU3C9q2
KIuHj2eoBpzAm12QhM8WAjWsOLyvJvARKaE8TtUMleiSo+gauki4mrlXjtqus8HM
iTrAqTtyqOP0xmSGgpeH9gZf4hiqM6qJe0NWHWDl/PoTwNTD6b3zVx9KOAlD4h3m
yFJsvIkoj67z8wGKsmV+3vogCEDXdror42zJzNbciY4lZUtFY/+MW/nFSM4+mOlO
Ykwh5V3jXEINLy6uz3jHCuHICpQJKHm2El472li05jIP3uo3jY5VrVabUGTvCz4t
1Z5BnkLCMHk0urZceRI95TK6+rhy1jB9Be4Q2YgvKEeK5EajGVENeGYk76ObY5Hv
hNZG9ZszIRzlgsRFiB4Q0ECYs2KJrrsfHLvmiEyfynRui/I0QNUfULgETeXLXRVW
euF63Q1CnVyJce4qOoFt10xy7jr6tmO+b8/s6FAuKoUd4jiRgkh99pW2TJR8S8eI
uvEeATeBBJ0iWv8epvD/BJOiqOr0pSPsGvhgmfIeSo8fISG6CtI8/uBvFXIMmJzj
p3nV8es0hS5qeIfD6B+wEDKjCCN2SuLK6Tn4urlFABvfyZDTqiYcEmeqq2x+10E4
GcXW+RKMpPZ84WBuXMEAfPmCjLC4yf/XmdK9fO01pM/MOC+vsStH3ezXutWiu6lG
lDy6iF3HqNhdhG0iJLyRjI2+FCfa8ICCmvjB6L37YlGedYnXyrmGslPOgxuWlvAu
rD2AINDLhHLX/OUnB3yc2DxCy39fSzfdTD5A5+yE/5NjNcHUJZewRD22nt/8xmQP
RsW+3jT7aqKkUX9rAKy1L16pJjHoLo1A82Pvgy7a9igg2SsP7JsRidJtn1IM+U9t
xOBuIk+4xCk6l5Basd7Ya87qbdOta8fk6oZ6jVdghTR/yq4CluHr2uPUodeaXD9W
dr4KsUkVVMC/tjnHNu4m52ulXKUkgNMPBt0j6e0lg/owkciTpHd09NYlcbudEjsw
gCV6Y2mvr5bU6Vge6DyTXqyuZ5B4zGIuv4v3eN6iF+Hagk6f429J+6tulG4Ctui+
L1bK6H0IzGzfIIeg3BaX1/wH71MazK0vRRImAlOqwAohxYuWFUwhvtRwQWCDKuqH
SS1MH7qEVzt84Kxib6JgBywoKvXe4zHSf1OHycCtU6MQfa88ivBIlc2XdEibHbWt
7WXWeo+GCacZx+8Ag3gUEVMFa0q9saZ0UrNvgHNkBw9UsXHRxYX25vnjhY26G0h5
ByMuCnZRinZHGd2H7MDaO9nPCAKgiAKcKVJORo/Jg8XtxHysdV75e2hifflZG2DQ
fxtrNjK/e3MK5B/4oVFarqkrgQ78egwOLNaNkl2Croi9kBb9Pw9pwn6+W2+mZy/y
G38lZrDL4EVOMHXszEUbY25dyTgw2ZmsBrsOUJgK58kHiesZheoD9OqAUIcvEaUn
hasHmprVH2ReHlzpb/ZBngSpuZpdJ6pG+XjtGEfQylw2XLUq8b0OOImgbIjQG67m
I5f9JTBKeilrIzBqgoZt3CxfFQOhtPDeeKtv9WXMUMOCFwKBfPnqddxqkyjRdOtn
mllQli9l2SxBQajdfICGd3DYTKCR9jkNEYyR2cI+L+utV1zSPR19WuvkhXHQKASP
LWYpWd0pn1fuArBBt253ddULffaqRr8lGOlQZ1DDo9+l8uZYbjM7Ms02gNY/HtmH
R0iT47GdMYOAW6+dQ81a3IQWi1HQCwnrZR8Cs+tLkLzOCtreg4ObaYJK472JAVDF
i8/W6gE2fscwgq6DFkMsrQsxpuLUrDQBA4kYbx9cRX9DUrG9yle1u0OdL9Yb9szf
Dim3E8gcQfm30l+S5A2VPRhudI3T+oEpoy/rEOg6KJJ3JrhyHd48lV5fH0llf7e0
+ihh1Y72BWrZxAvtim8O9+hTT7E16lLqI8fLq+cCAKGI30GNrTWsBg5+5cyz+EgJ
ahe1nwrk+lgo2V+1ndnOMEqYo0npqQpWKC5srbGXgzJqQ6+TuuJc8EmnC81mZfhT
5lXAReMYdcZ3DH1uFVTUaV7V5Z7Gl8kdAo6ROZzqFQGaRJIGydWt2d2YTIFizt+k
Dr3GcY4GxVkteFLtySZ1gUFgtCLLbpkHwYyt7d77VGCcWMCW/pgTY9VuaD7Bnyqa
VuDXOPCfrN3h2aVCNhaAZxlZlwn+kaioe3FBPVVb0t8vADlen+UPf3fpl4dC+184
nyv0wh2njYMSm/kLfZ30Bxuhc5Q+ZA/OHy+3amiMsulhWYYGv1g458Jx9zJMqvgC
H2raIgw478XS6s1KKpZtcebjMRDrhedD+na08ueIE917QtICqLhwzEKkQJcpAitB
x1vx0V9y9dqB8DSQ47M8I4QQyKLNUi4/PZZsOg1msJjKzvcxS09y5U1s9NXLuntf
93kKsI7MP1/XNMmYgbyWpmc5qm4nK6phClOk3w2v6fifRMYcVbO8qY165gF/egb7
xtUZO9+Bll/0EZAaKZP7HFBuGE+H7UNfb6w8qhhdegyWLqUm8ROehv1E4Zm7ZAZm
PxpDlZ+kUMXjUCkkFHP66qcjRfzUDrRUxXbDEK32lyoJTfkbDSu3V+hJj2OdybRf
RL5KdkSHBnqBk6gpievlAN6lhBBofTIQYw7NeoNQF4yQsZVXjlN51Q2C9SoAvidZ
0VnaDK6TEbq4wUHKr+YBT8rthL/2gxkKKTpZ5QmrQG5EA3rm1P+AKfwH4X3b03Yn
PscnvKUj6duBle4rVJ2dFdAgxAavVOxxYSWz0Bx7kXKnpbkwsFuq4IAlCsEngtOy
8JT8bqYLM1lLBgZbUffkW7mOQN4Zb1pXfI0uSsTmsXEJH0sdaNJAacYXSxRtTSNf
WpzRlLOkM8BtTuXjjie4kNGmcpH7VCOdFMpeG7hcHtWNfhcWoNbkNH+TQqhG1YM6
RxO+pdaAJkML6uvtNHjkcX636T8XGRwEB/fdrzpSeWijI8lIlptkIYA22g3TWReb
vt9WxrJpEDmYiLFnHetqNtbVpQ3Cqw8QwRh13gX5uDqcYrSyvm91W0Mq7/IiDa0e
X+aMfKQd4gDhjSxTgrUTbg/EvaZwx1BLMPylOSZAJn3jG4u8Ic7Si/F0e1cXold0
qLxqgQjmEGV/WheyrFlWy2m7fDXK9t/ni/IFK6gEiLrHWpUsx18izPhkI4loIOl2
ePDYoM0DBhioASkNU/aD1iHZlFzYrCT9ho9/Hz+AWU1c9v4hSkpalrtUeprusHUC
HkXYbhlHVPZp2QilBkgrdRJZfWT1vc15ozYdNlclEzCWjSBGBrlL+fzlxW9XnzKi
M16hL9Ci775UWurtwJxf8s0M2/wj9D7gN1o8hIVhAYPRN7szXsvbIFCGTu+su8rk
s6t2mLa4YQ/Uz0Fp1t3bBYTWWVfdGJufsADjHQh8TFJ+RUmptiDX60R8pukHmX+e
6gJtqbMxNleFSd6nrZRl0Gd/KPBDccaLyHnHeyg/OwTAcfOWksYf0XHvV5Y7hKQO
D2hP0Z6O4AyVOCmo9CW7y3qzBVqyrlCy8WaXhyUXguLKF7WxX4def6BXqVrGzSb5
kd0FaC00Tc3GL11Eenh6oJvzFPG4o/f1vM8cOQ4c4p5udkSXAC7hsdCH7XzY69gl
v7FP57YUlmcN4Uk30QNR511sOpkKM9GfSrHHVrcsUxAW06LaT+XRfcpb30UJuV0X
8XU38FD/bBiZmlWRIYBM7RzET5UlPwTSpzqRRJALOzIely9NFtIHy6NHKXvSfc0F
YNYovIfUtxmoRmPv1PDMd+8Ts8VQmDivMWYvZSqUgJfT6c6XzgirZ7N54MtoV8FU
cbXw46Z/M6CkgFGqgFY5cSaxinxZsI5BT0DA5AxjMEKmU18t/IMddX6awGo2K+JR
KKTxvUu3y2RBo33KnVWQl94bOn8llLLsl8DoQNzRZVrbf1dAhhw+p8rNaDW11Sc0
7kZFuB4EOtwmViUnXQMxKozb3InD5NS8HF9Dqb767dLwGGwp23PKy/Ie2FvIoflX
Dj444pXR2pGOybpdC1MQypjJ+iDmrYQvp9ziA7Jdwp6j9hCjOcj+dOkS6lphitBZ
PgYwkqauOdzwsJHEKCLqC+EUYiTyIyl5E+A60M6AVkZrO49vU6tp8yQZZNibik5h
xBUCHnMp8TICQ82DYeZUTY3XvlhmSVxhYl1AcTRTlPufg7k9lYcStjbFZZIw7W3a
TQ3o9A8wn8JkAHmJeN6y2FVVQfzdD20PfdTwS66QlIb8RZoNa4devB79H8CrWrYb
gRryNcECg/Aji8+mxqX/RYdfV51cAvmhRCuIxRNXJOHJlm13p/fLhbXQRM98Ei8M
lmkyylCWYsME6ymOF1h3JdygPMxzzBhUqepRbnjcuzpg8iLOusJ1lsco2ITrtV21
+DbKWCBW3XXercD1Nchsmy5alefhxFURntn0tHNItDiMCwIkScgSDM8NFa8oZSJw
eoJkHUCibc+yoELEnHZAUg/rs0uTdPLSE9XJDmAQDgwsAScMA/6SIxgAJ3g6rM35
DhjV7/MUgoILzA/XtuBTRx4J/tqlW658lj7SUW6AhKdYaJC0KknMGiBbt5sDZReu
CwDB3B8RfiMIGDLvSGcf7dsAWhexGychNGm12Da5w1T8q8Y38JJGc3136ZLDP6us
GDfUtF/KZwFYvTLKm03rmUE9+BIOIuRQjLSHbK92r8u0JFhg4s8hoUl66PplUcPP
JmaZNpZZD8X4fodt6wcQvNpqb6LVFatwIpw+9iIy9rNVOMsgJ3SOueQbxAMMYBzk
xbdlvVqjg9C9Rvo3JX/uCVmJvTJY0nMlzrJ1zFNX500M8bgBcR4CvitvP3/Lyu4E
zvp4doUb4qij6ZWi9IdCPKCzGrkJZR0FvVbBTk+7iilCC1xu/5xR41qzvo+4HKYD
ADauiAmU991kCFaDooY21BINZO/hlWftJM/qefGKtZpx8G8yvkbW3oj+KC25FWTX
lguXgqmve/qT6G/IsCaPK5X3cZj1f+Rv8vNQz94UcyXjyBGya5DdXcFhZvHeYJyo
TgzAvxxETLSPxZkbigph5Z+V7tcExLzuF1iHQDdKOZGGFX2I3CRjAcvJmlV+63S6
nJjNRF1mloa9TYBlw3a/JWrPdDuRA2Gudx22hp1tewxs2Ub35yxPLvnCKghTGf/b
OQgwzHLDcGW7IroMx0sSWEsUa7Wgq5XktN7A1JF9klrYUkIJl69FV5Ga6inpmAoQ
cFAi1DxTylEstF/1mu8MVC21SVG75A/qymxvDP88LltkH+IhGmg7hhKrmtxmT23Y
9pGGwDIAMPVpLIlBZIEQaH90mpX5QsxCj5M7FiCTzDKeE6k60wxWdZduAvjrAtbc
o+z2ETxH/J75KHxr8HzmFCaPj/LxNh0dhtU4mUR1VCXSDa1eloQIoSvaXlUKZUYt
a/s+4ZgkkIaJMILe+rrajyVafNjf9vF7S8rr0zRRk96ZZ6jVVschQnHCx2x8LzqM
QRFsw/yn8/eWYuuDwOQzWEq6TsWRmDnZNph8gWaMNZH0dtnd4Ye1CbyKboW5lPO2
ILHkEsl54xQISAUkg8s6er0AWAQfABkDZIjhze6jSqpDlM+JCp30mJ0QOLP7tGQb
LQrA+8ztCBLti2OITKSuPLMIaVeN8LBWokUmZqNU65isU1aSqtGSS1/Kt64puQ80
6ythxvnDAWlF/b9lZ0K0b3R0gwpl62wrlyHsgW91rhR7nG5WZjtB2Li/0F2gPi2o
THCC3+27abCUR9Yymxd253ZDO8JYKYrRz77G4kUOBKkTZs2M4oXMIF5raMMdY4LF
Ff6afsUqDDgGNRxD5plp6eTTRP0WHxJtGXWAtQJkNsIglNj84u0naHIV2UvBorp+
g5fSN8eUcsRnGMQ5Eh6tvJKunXjI8Kdx4jyijnUrcYH+zsigpOsob+pIZQVu0Flf
iD3NLFZi98Kk7tgUNYDeYqO6UfMayW5NuAwkgI89DolJIxDqQJNhXg1ySk4PTaJD
XFTLelBqxLz7lZAFWywVTFVSguDciJ18owXs+BJOz5bS6XhGzbw9g8shLxBCBdk9
5l+eB640qnVfEVSysdi/OrSKfawlEDPYTQcqxZy7a5caVkAgk2JWtDB/qZIls1zb
8dq7o4AZeSHeGvbTyzSqfBHefjoQnKjjDf05HNlf2csaNsjQ+ztSzR036Cb0KUlL
wEmxDrlAc22xwtg5hVdzgBQB9szHYqurCYENHXrWE2hf1hQXI0ZLw53+tLZ55NfM
mWfYQDUMjyt/Y1LCMZ6WQtC1Br3sh5UNzUqx8zngJZ6WsajUqRFq9AlX9AkEuPkc
TDyuDjIml9ZOijb09sSdvaft9qlx7VvrnynMaXPlR+UCjeUwEiS9RfUdATWRV8tS
VYLFq2Qu6+rm2VHan4/kS7ON2m4rD5glVv7rDYCiZTlj60x/f8HYxfIpj7JZSx0Q
XRIlnaTGL51AET0BiGDpNY/j4PkOGYSkfu4QqqZV6nXIJggPIjfOg0RmH3se9Ie/
W5uLjGuawDRUIDyk6etoWX7QNVkMGNLfI21XD38Ly90IRu+Zq/uFBUYAm1QSbL0h
ypl1F77X5y2c4Yu0R2r00Bv4+NAb2mnQymsS1p9XEfznU1deQLv5FwQoprvx4DCe
jt+gLvBEwZOBoJkhUiHWSjwV8cqssztvftvNRI0GhnZt6H1xyQBYiZECEepAelPZ
lMMRZezEhjhCWZI4/UgNoygsngkQTPJW9PE3qAvt1aEkRpbMH+eAcYk/a8E11jUh
6s276Fun9XvdOHP+ofDvs0jJ2wwZkjG+vThcesRHmOpwROYMUO+WE+lQcUy5SLpr
0gPG4TqKitXU9Cdy5dKL872ZA3JgorqDtMCCrP36L/dnAFq9JM63Lv+bmyO+9Gea
/Il2k8RI7hvwf9x4vMNqhteL8Q2IxSLJKEUOBTWOgFaGyJnEL/WY8fwZKYiHQeZ+
1sGBTKE39zfsf+fiRPnlsvENvru0hUQJF8QRw9mdyObuQXtuLwOFy9lCUqFdKfj4
CfZx98sq+jAPCpcfhxVbwF+obEdfuaL0dXck0vMN6aFfpoNk02DHkezNElTRg3A5
dtE7UEm7HDet3YrcpzfvNjgt7ToBcbn/fk0XKmnEOseS3fsY7pARZp1kotgAXSDt
LlWmSkkEwD07oaV8CqjAPUO0lMBq1phetO1gGB9k/oRF4XFvJ+N2k94ITSTvw2ur
4NcFu+bZUJre3MHcePgX3kwkOtYCCjDv0+1dYuU7orcd/op3fgb0CkY+MMaHUAwh
NVj9JBxpqzkDcr4LtLNTgYN2Nf9M0BQ7wyNJWO6NVRjERh0Xt3Azt/CamKwUFPVg
mUs0fNOx8aghS583Zk4o20iP7Czd9dhukNH9pG+IMdoFmXkmhUrDhUIvULHqcOx8
4iTEcKMVX12IhMSL2rABcpuiz+AJqgdC7jwsikJIzly3BPdjcfWOM6mB/sx22jPk
UWoeMKV8p2o7aLPG8eqpgLv+itvassmYooIlsKqVVO4npyLzkvkerDe9q9fwppIl
WnzgRHrXbqpd4D3Y0Q01Hqta3D8NQCpefn+BGhvAtZQeVhNB/suYRZx9Q9jdRifQ
yEfpXw5pzrreTGi+sIlXupM8+7dxxL1oxQ1sa/UvYM2GmcuZZL/vbh4i5GAQzEhR
yPP4z3An+fSuZuXawx4tTWHsWy2hGh/tIMeVaQlVVy1+tVTLQGaV8nZpDUOIggLv
7Q0EGsEivhiNh+m3loyIplpMCkiKznz97mr4dYV4PsxE7vhB+fg/CP1UQ3EnJ5h/
cV4KFiyFC8G74K1GRQuBP3aDjtf044eekcckRxjNZvTShHYZkduvslddZNIQ4USt
7a9g0tGX9r0OamKqYbOUz5BA3ivo8zWSVM/IXlG2QAE1PdJPD3aA5undg/ppla7v
c8LAamnaPUWaOguoE9QAwbz6AFsbQxw4kNgbzz9WIu4WqcgJ0TcMrDxLm/D4z0aD
Ry1/PY1x1WKhhQB9Kx1YfiAyWTTr+sKgBEgf4stKn/pXrH/+oB0ELmvNGhXafVta
lwLyHf4ctjB9fYYF4Tz6Z9aQjvnlZWzhPCLZBk/YIzM0tOKAHcWouP8bJuXlGwh0
3ieg0Lh+zO6PlREo7RQett5QvCC+FTnOSvCKWKVMdH6JOL8A0y2wow1Oj4UijogZ
KjVMLEnwb7wWY0cFxTKbTkBNESxQ7Szkke1W2ZUyBSZ+48YtIr39+2NmpBVq7P39
ME/KpCC+mF2Mi7UscdP0GV5FNnBBt7vgV78voXSEqYAZ2/LQWvBtlZDWbDMUsYgP
ymSNqSZ3rgWc3SktKDPrrWSGEmAvy01i8J8aXfzCc1/O+HAq3iwcUYXXerD+msFi
v3OkT6+daOcGOiWnMvjeRL8Gsh0G5xmQk9PRopNG8PQWfeCG0ySQHaSA0eCj3gha
pyICerqu5IrUjIEt4RNx6x+Y+HFllc5w9C2tqUB98TNsGfSSI/+cGIz/ugf9iKQe
gp7+WQqG3FOy9moE3kFXnnzJFiCBIVIFv2n/YQaMXn6cRlklU15rDUV/YWtJZI3b
6t2ShKGxLBSc/7b2vKOJ13UWdoPTo5j1ikdVauP7yuo71FLP984MJTiahI3f1+jk
kwLxvUGH25BtFcn3/1S6fkfcm2eomNjLl00xSNhMYHnec1EEbFrV1R19HXwboVrT
8XB3YXASJms9sF3A8BHWmZ3kwZKAyR893GrBwWu/KPeuEtk4RHUi3iPQR8losO5+
1ctjMFTT9Lwr0BSJi+InvTTEV2bFcQsYQ86tzyG+s7DxsrvBx9hLKd53dqukFDbQ
axYI1bI3H32qYj6ImSC0nSonnzYoXDEi9WoZZTKgSvjyR3Ct57OZUqdZFlafjyrg
dsicqi6tNURBYDsQHH7qWGBk4KdgstsRSNtm6WelLZa9l8S0pcP+Nh4CO6Ftc8Sd
X8ut35Rt2nEKBzT76YkYockO3fnD4k8gmLqoQt2OXCmRXwdvpTlK3OXS0ZiyMgFd
u34AmOTeTObsHR6AkQynisig4xawIqsPszOWFZIsaJU7nXxDZJZ+5A3aMMJ8iBqF
7MZwlUuibQIV0skFMxYFwqSWteO2ERpBegjx7SC2OV+T5/tghR3B2+4+T5EHU4cd
+ebEh0iq4AyNsIBlPfFKfwQCLH5YEudhB43NobnC1FFw6aBf+ajjV4bbH9mOcW8P
MdszD5MN+xRsfQigVyhAeiAY0FV6JvNwGBO8GZCnqkQ3raUOB10k8Z6gk3AazBMr
LHQna0YnQItNywh+B1qAqlkugun+EFBEmNELjbJFGxVZU2hoPYCkqOyy6tmqJHoW
dvYCq4/bZtLK1MnQF6lz4owcW/QaMj7PGrk4Vd8nSdLNcYvc+PDH+8O/K6jlVTDB
yM344b2PIPo8/xgDQfpKeJegTqQcinI1ntl/jJa/XgXw69FZlvJ0/BOP5dWukEpq
WB+8Qr8iY25QHZEte4VBkZzr/Ym+VU6C3SKIZ+LfLBZEVxcPKYnLrFB9rEX07A2s
pRHjnLnyujJyPd5czIsO0VNcCbGkPPR1GyRVFZUUaC+aBgqPJ34aTSfPlw0sqV5L
pWiQYIcohkCWBkYRl11sr8mt9zlNmj7HigdsbXSQBun64Vbw9NiKZ8VR475WrAVY
cBo5UGlVAp6lO6h2myTjq96mAdCo4Gjurkqj/zCQFYt9ODhdvdadS9a/NELZvB3a
Pifd+d7kVBRB74xCZJyWCTixlrj2FDfEDrwx3UcMVWTKnPZyys5n12LQf/Do2qob
MFp5A5b/BORiWz3PFOnCoM2eZX+0/d5HhiLjNTt/qbbpWLaH9lfzYc3Am6SByYfy
sn1TFdTFIEQZDhT2F8WAm/B/dl5hhxwID13XANLJA03Uoay5/wGJMlf6hXjgT8EM
USkg2EAjbzpOFmoO0ljwM7I826Vm+/C69NRMdEDs0oe70UQVbKJlD6/Mzy162HGT
ehaiFMQWA9HQ+z2La82P3J6Z5LCY4ZrI/ub52YlqUsXFst9dNJleJC5Rx8aZAmPq
HKavfdSoGg3F5ENSHJ1cQlzUWKYjFWZ3kdN0yboKYtRty0q/9217kdys46q1TCP6
cBPtwMuPU8lYbKrAfEebNdQTE2UB3/amnDqV3ABP/K/s3jwZioLmG4mykAVbABhB
evl6v2QtVEqbhofsj172TgKck/LcaKGvOXkF72utkEJYyBg2N9T9NiBeYx9A7Sjd
XXYUtAtYiB/KX2kzGQQEGaIOVOELtfEybeIh2vgecJrrFQiF67ARfdaIM8OpanFG
YmqSjh+i++mkWuU9UiqO7zZ2kBdjbwP35uTDIv6+rlyfWNSkfAJF4eVlM1yr5QXr
yldIKxypGVXvhxVyHUQU5eE6qGKWUFD/UN8fkhq2Me+Lgt8gRhUDgc1KoKmGQBEN
IuDkHj5Eis/6/ypUqbC1PBgP5EZDR19AclFMrv2DqkB23DHik3szgPq2wvIRJ+HU
CbfJwrENXuy9yo67+Hw08j3TvDyjdUjqRYOSopDNJNoeqXYuDZsU9xYYz5T0vCxB
wV4aCbPHXP4Q1hO2m9hm2NVWPyaqPNO+2CsVSWvQnYmIIF5psdIpLqkMqhifEyZ+
T2P+LZ9BC/DDpsTnYxN3IR3Q6utUEKBh6RhpP7XUSEXbMIfz0GN0DzPHn+tCJT8r
c5G/SnWYgMKXjDWRQz1La65ML9kjX3G7y4/tBnYU49EOEUrSh6IL+OkXsUW5XDBV
1wC1f4S938diAIK7cfz8Iux3ESQ5JHzYXj8goFo+aCmZhozJ1tZtn2Kzp5GLKqI2
ox7NrCCnlx3V2w+ZkKay+MqCEPB6MDvfHnJQcrRIFPipAzuH7+5XIqqWEzAL/LIa
pATBaupChLYHv221De+5CI76gSsT8UhUwsy4Brmw1SxWDPdJppKJIyAU/IhZLeEo
umEiUGGm7H7GYwTpnNAX7msGT1R91yayW4uiaG16SDlZzHsy7Q0uCe81VNRwNjQi
NSDbxZ17BNZNAY0YFHPJvV4z6Ii+uUtxbLdbXP4eQKPiYNuDWJmqRCcv4qC4Wvk9
TN3Mohx8uCflh69cIDoi/Ho1rdTtJEz+pGMzUr5lM597HZ9kZra9Cd2p/tq0jddS
hQyNJSviGPNTfIBwWMhRALlcgQ0YhiE5vCac7b935LDrEVrYx2gPpqAH3ybvhycn
gtehwj3Eq+YD6e9ZEaarSAmWSjbTdyvoVp4jcY/GGtVxZUzOxXRj928/2bUv4L1J
4HGUxOdGAwOoO6OZJRp91SSEHx3XwOz9ObTVMzTCRr0KDiInfSdQ4icBkFCJdJZR
z6lGAlR/K4vNkTHvICCfEpr15dkREeNqPeO3FGlKBNJxCYoUNUHxrLXT0dCPPz8v
mL3UCDRMCTomaNEB4aIewL60TTgwTrYYhBrFi2kXdMZBIOTbSaanaVtT03NaFnkQ
JubadQZW0ZX33dPGrOJoYfc2cEExebKf6MFo+99Xrg9BGUFF4iJ38+vHw6gW4sU6
KBciargjaL5it8L539W7+Y93/Cz0YdhobU9QPAYAk3qEtQPSI6hVA4WjWjxZgBAI
4tHqtArBfO0Rzsn7XtrkTlzHynpOWTQkzOGJGjNT8799B3jel5mj3SeuOmrTn9ne
+UY7PJD9o+ek8Ot5Fzhwo75jbSQ5MLYTpRBWS9xKqNSH+LICzOO0bGFzHt0LZkxk
tkiUVMl9v4HDBsHNrKjT80YrZZ+6FG0GO5fS0ttus7I8MuXcLSI23GWYQ+89Ty/h
mMB5MLcgcew0opC5YBoMTqsNJL2Flf03USGbVe0sfBiJBUo/IQrznGzxFMSJXauy
2kwZr+E8iCuKpqbCweNXPrA8LNRnIGdq6JVScltBUQO2sxeC2Z3CPziGvHtyMjON
mxvsdj2FeIZQO1CL9DBw07Bav1kqdqdjVgeDSjzsNBPNaXwWvqnoBz0jLuMbE863
FNteebIcDqdmYRuWZhVKAlXVqS9iFUz4NLAf3tHWslQirWslTNZfGjL72hpnAH6z
d2V7eTHpWBUy82k79eKIT9aBZ+y/yebdO3sXUGlza+h3fYQ7BKv4EaDDZWQObyY2
X2IlO7osRhv6E73xtJlXo1pP3c9Xg+eG7J6p3ywlWV2tbnRB2Oqf23smxxP00DPo
kxG1VK1sRJhGejwkdMr3EfonNrhTkvvO9pDKwa6lNgjevfsjkf8L07wKcaxFqwSz
0zSxYJ+T9owBZXTV2Tf1D1VKWSFl4o4PlHIpRGwpk75QAypy9oc7YknQNHHJfkYI
d6Z3rMk0K8i136VpjVw5/WBHpyq0CexflaGF8AYcLuPN5KFcZBA1Gtao6jT2nlTV
clAUUo4LoW2Ccpxtxj2LQpSnl14EtEdlKmcLvVfpNK5M6inMkdt2AvYMad23xNuJ
bICTbLdXcpbtmiVovz9IIiDUllzJEVemSFnkYt0Ag/aB3QbHVituH6YQvcyy6TTs
Ip+cnu70wc3AjlW6vXGlnOsgF52kSgXyKmD21UnHv+jeeMfDObbsWKJOLZA7ySZc
hDGbxUswssbZCwNBoX2vmARzb4T3h+kdooK5I0AkN2PCPABxj7Ze+wI9ckOwAuMu
SlpBQWPlEJLxZQIF2PCX4oiXyyHxDLVApqqx3LDfw67HrHhJS4gNcZ+LMZge3zPN
KMgzz/S1QTnMT65DUFJwBSDw7p/y81qDPgwT/eQa6VNfhOIHrhfvv06TrE7TsPmB
pHNWw9naIy9kRSm1LOCdvBKbKvYaTV9vHrtWxoYbYA51mtGxk4b3VHS2X8tZlGH9
3iL7JPPrTVlcV3raVLE6AZF21e5M4WBKUj8oHhQZ1R9FSRzoKdBNZ92apE8NHO4p
uiGF3jIBxqt26ud68Gx7zVmHEj5z59OAkDdcRFxFcEnrAp3u5wK8xidfU0Mb4YhA
7HfM+OThwZwOwuolN/oFYBwLdbTSeylhXbwmlfmvQhL8WkqGVk8V9dKYgHX7NWEu
JqgUvxdlaEoAUcL08mmAIURLWmEYu1xAUVJROLTeBsrrvoE+f4LXuCtEGDXIZRuA
YcQ/uf2S5HgVsZohQPrSInebbjqNATZgfynrGi4r9vSvG2eHU0kpV8a++vLK/tXE
7DQ5V1ZU0E5XPEZBXLU+YfjpHneh7B4CHi/QICiH6V67EzKs7C/2YHMGwhoJOYdk
G0SUHZ5HyrwldfQKQ0BXEt0Vvld7kZvD+goI9mHKSEPNtC3HYSKbhDiUAyFQTIv/
wp5rCoOk73U1xZi5Ht4zMfFq8/zITPyZCbRV2p8WgcOuj/5rO/5U2UrJfHDv4pnc
TX3xXNXNwarOKYCh1cfanhbV4519fMTWpp9mnOl2sKoqBLhQRBv7c4uKCw2k0+Yu
0Z1kUiQxYhmrB6O69Xz25/e1TcWagLk36HZkvfIK2jqcQnjwx5EHCzwhWkydFhae
Xe6nC7vSLEL1sPlQNvz8ClVrWfoziGyaMgRCdXK3KYnUNi7aKSh58NlYIxPxmMjZ
u702IVACnRK8/IyN3Fros0RW7LoJD52z4odtl7EqIdRTNyPSv20f4sxZxnUaPJJD
UplvQQKVyeUQOTRxdeSHTKzmuBwO3xMsUG2roi5W4fawKAfwEGZwFR8U7WTnNjzf
qVex5rjWaYRLDUyCc5WLXyvoZy+gi9YBIWWii7ayebwFWI+Mb31hnkgQPptRUGwb
A8KVYAIprd8C16m0K89OKc1cDWQ0jy+LOIf5mHIWKnjoQuCDQpCztfuuUxt8y0LK
k0+AhquKiZhSElzvP4yQPAX64Dq3AJlSdvtWS3SErY5igX9H8u4xM+wVwrP4WFD5
Z8vXrerWYdBe0R7JVDWdrHmbQdc0zJw0HCoJ/2T4kTBlrWNK8DMKfk7qqnWA0V8V
TvtSQNXwkt/TwLm7IzDqApG9wh4CidZiWxVIxOJhP1qsiMWEgWVWg37PxMoiXMQ7
UMHCRk94dScOV+PYd+yONIsnfYhhm59qagdZNbwNhduhXG/nG2u9tNLY/YHVIGN3
ApTICGRY7kFv1M5F4c7UqZtvLof4yPPTWCqQAJx9LUD2BwyR2ZNf/kst3NiU3Kpg
6ebeY9fcj0ayjs45iNeo1JeyyDTJ0hWhM9/Y/a6svANo60Knx/uEZwKIvgn2M6bz
F1+5vpIqMbzR7NCfsMLDiIxj6Pnyfa2GkPFCssF/wM7I3Z4M3ljEnRuwd/o/0MCt
ZVqDdGLoVmuDbQKuLJ6LQdmIAqj0oO3DFnrg7NC6OrSzokueZQtMjDNNul1qDs5W
ml1YRC3P0jckH3AYSn0uyMmPvMfwxkdkC7sQcxuF/etVH1tBwK7Gc2KaNDYEX9e6
us2E/p/0nslnyuh0nN6wxW8UUtBG26Nu5AbZ46UJoUhIYdQ1Zh6+yjjQZ1/JoL0F
Dhn/rPmEnDneqcnkPE0XBrOaHCHzzWq/iNKQgdg+3jcLjLohPmuNyGnn4LqM7mQG
OzPllgR6arFFz7hOf2WaUrPUEGHL/m02yBX6KPqKRPuEFvJ4YO89V78RroEgCMBh
mjpcr8UDljO9xIr4dwjOoV0HvWizxKjJVI9qO0INGqnndPNjOFP2rMwwtf3HWbLu
AAi7hcN5BwdbgC+H8+pNcCYqTIN0/wHWdJam0gM9ZV1uFLQpJF/1ZcDBzWXLJT2h
JeFdqfILU9ifowGH2/wbErVmhQpe5GZKTivhNh6FaT9ovqvBkcumROEqHBfk6O19
Rq2/Sby5ApysuE2R9cMn2gLqbtMPRCIIn1ec/lsAvpoTtgJI6ThMm14EYDkn6DYx
nLJR00aXQ5TOxI4RXzxzwaswh4HtGsKwkUXTalKWQFVC5NH99A+HLIV1Sppi1puB
hKoxsB4Dx45S4U1asF/Twsr/nW0xtBCQtNiMA2UfwVOOnQ585VVV+YWYUEV4xp+w
prN+QpqveyzD6dHkR+921uWK19YOh9Is2KnWZVAYVCE=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jr7BfUUvlDpGDzxFKniJyqUoJPFn3pIxvTvvYQjzyCRvBiMF7lUPOWrdGN5nJumQ
RGIEZO1/8YyzEngYsIbZfhjvl/iirbeUEAh/S9ldApJNUbN+j5Ln35FDiTZZUR1R
Dm/6TQMKtdJnKBw0vljEPNK3E2lOLImchzZm6TvaHMB1I+FQRENfB1HtuLej0ZFc
batyd/aUL7btf1o4L25DC59blCHKwH0Y/MotItVSp9Q0f2+aqNIPZv+ZFQXUkVeA
mWKDoyr3bcilg+j4Sgm5mtov9PrSt9L7dHMA/sxw7cqOATXea8J+j0lxaMX9+lWj
3SZpneat7krD+Ck3Ld1NuQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 22144 )
`pragma protect data_block
Sn+goc6HImISjaIA8+czxfqJWQlMfB/ibVRBdWEGUIvUJ1BX45C31S0Q2LhQAwL7
hASVaPZqDmh23G1FbViDRx6dFrVj0GdXijNLDoE4w0eqML7FDTHYolXomloyJo7k
mwNI6WFJKSeJYLCrpZjbKLhmKvm0SN+vz/xYhVdeMD8eka8Q4m6YRvnmjIq6Mc3N
AI4ksODU24bLkmFfbHHxs1L54OtXbuUk0RmBAbwfvkOxjPK4OwRmLlQo+q4STg5o
EGCyiK75Bf0dtjbk1d7AQhIrFnEuKFnHfhhisI8lu3bmV5M/Gn8e29p7U0VJ9LdJ
QJzPTKomWka13eQiHIE60GVNPAnaik93QWMma7u3GTd+9kqeoVHYeRvGaAHW9IgT
97VQc3xEmANX6CIGbfkHA7Osf/414yd/PBfhnUAen8e7KHXCMd/9Q9iGW52Q6aVh
FodVfD+g4yE8z0+yzq7LVF+5kseq3r17Wpx8E9I64It5kvm4Q0UrWZ/Gb5JlJoZB
RnZU35eKUxQsenRTg0j66geM3thF5QuUxTd6G7qF4HxYisGU6Cuyo8zePk9FW/iI
Q5cJsioB6Qi9mSsnzUNNLg7+Jy5oZiRyBiGjvyuBhmuoDI9JcjMTMZF3SgEZIhmt
IhE8FgWNSgjNTNzgtzdOY18Yka5xMAvYov4Q+7kGrkfLG6g8mznqzzqs330SMi2j
ubOTj8EFwcC0D/Zq6N6oGx8FPK2O+Y2zkyuCOkd2zI5MII6g53N/hGqEIv42br3+
u0Pak3/E6nUn07UtJUSqM1KfOaYdsTm0Yi7VC3mF3o0/u+ukxFz8x4JzRLD60JH8
GtbaR88f85hi6sXMuytUFbEjyJAYzcRixtuoSMKbqPydoZolx0yRiPjE5CWnUJ91
mT9nXWp7PzbopttUx5q+7WiWz0oFRxwmSk5Bj0dg/GC2dvFVeLPorRBJCnAUFYEU
/sECAW2vFkoDG08b3MmurvEbtpedPg4ujRlQXnzOj/uxpWqP8zOytxFe2I0UpcmF
sW4CgLuQl/UDaLotL07ziWWuycaVk/sDkOyH7bumiyNRH7gQV/ic0bk2ZYxSmkrq
a9ec4OTvhWF33QK6Z7Xshj5XylaIGhARNiX3RZxAI9495mwz5nyAi6GKx21kG6MU
H6RG34dbB5tsMBP059y/yn89cOhjr7L1R4biQUF2J262ioLcuKEdNDP938QUF/Xb
IddLEQ3QNt29yny46dkRAofQy0ugZaD5wfTfOCWB1FxnIejwG2OR9iU+g0+LiA1L
PQI7ctJEJbG5muXUgsRdAQvdv6+53cylD0mqshNeh4aRQ01rvXCnN76lhAocc4fM
ijV9/QXpEpagAMjNzEFTbcnUOUu6M+GtYyaqIv6lRJfFUb6TNdNyZ27M4zMIwPMn
6b3iZPSr9ayJqQIKYLZ/rCba96khNYhPhzjbcRZvAuyQGvH9q6TjasXBtZkECent
fhpmvQNk9jHo1V+0el35G/LUZxCnPk0zGFW03nJKS/qmcFUNJAD91Q+g7DmGq2/d
lbnRYp5zNEY0GTm8PJko1FCriXjlqecUKHPU+Tj9QR3IHaLspFbkUDRnfmLBfNvx
b6CfqcTgTv/YqsSdoL8P+AKAbIXdMcb8tdGPcF/XgAoPf54btqm/s4UIuu4vyKUQ
Z35db5U2FoEXgTlcFwbpFcp7V2ivAPn03VrvHJvEb/IzkaRtuOlLDKRXCT9gD7u8
RYs+Zjn564cq0fOJ+6cdH4Xea9xxPMmkIyYZc6H2G0jiA3uOdPhdwRQv6aDK2IbJ
3iAkhj4oXOlDqVB4Mh1YGzZg0u2fscpIA/kGUX/yrvgiCeavLfXHJEX5E29BtI4M
P2SvOTIAiWYEwZrwFILshm0jQfOxM6d/pgv8XP/QQ+DVcmylcOByCSDO2pf5XtsP
Fu7G7RHsI6aFvgmpVmB1rTWIV0yhWgMNn2VbzL7/4f3JmsfpC0YSOSh+eVjxbNy6
PD8EUxleXZQJCa6GrrH8j2HQJgobQgcDxevejR7YeSvSu+VrAi48t/Q2w4d1x7v0
cqv5gXuQji+n/Tja5+T3O4/qsM+7Cy0a7e06O04DcZRuSbzzistCzFXZ7c9zuFZP
qPfX0oS1xhxm+AVnRwP6zge8Cg9dfAP8vZORO2/EO9jq65ibdHLrEPlPAnMJDvDu
rOxTUfO+fEtiv0gZfWgCJ0Sik4LOvctfEyciFJE9Fvnu8rn3mc85yqn5goaZJ4U/
Iyzm2RdhPkBy6vshj2w+lV+7bADOIpXcbwJD/7vcEcnnH2rO2C+dF4bju79vd68A
9WMsfaNbcYBB2vmqNjhT8MfnIjruokbZ9IYs8Sc+5Jh4CK6tomWVIonMAXUog68V
6T1R1uMgAZ6qGfJU+9gy+tS60LtOKuKGfK7kxF738UvsTjRGuCWXqILXJ1e44XJ8
UrTzefjhKewUzOwiIulq7RAvCujsoc0Yb19oSb3NyDZF9RLVE7PnUkb4HYa21Mzt
GDzEoO2xvK9B0ovr1f0V8+j5TYfrJHW+nlRfFyi2zZ9RipFKy/J3KeE1dHvA7ClU
7TrCoD24H3g3tAWmmlmUm3vU1bYTWBbCmrhHA0yqHRbOVQGBTRtGxf17A7LkoJCu
1V4Lquzb3dB7OoI0LJe1Rnf/nTZr4/LBOIzwO6LnJxbGGYr1lVmGlTO0bSLJtwgo
rKcdwQzSEhVcOkj+9HA3QHIGvDW+KtMOQ1hUrNWzKrWA6Krk0FNUnAgVgVprfTLo
cMCFk+0kkzdEvMKUsuV3E0xLnRlIcRqEgnYGwsfzqSIz+9FZPD42Mvq1OxZfg7H6
6Fa88zF2D2a+o3/+c5CY8gD3+E9byKRM3hP94sBxkeTfr1Gbs8SI0SXOYGpd9pGA
GqfhM6vMyqZjZUBXmspQqWpNj85VNAFwGW+aEGGFk65dSsEowK8Vc0bV7tou2Awf
+kpeYTMSy03khiOLszrkK98Lf1K5Cm8ZhSTEFJem5+uUNzbpmO9VphKa/u1HM7Qx
cM9t5nTlDnks53NU2nbosWLl5+RduCBSXEsNLhIP8P9NZztPasuYMSkxwxh8gomv
LXe0Dfwr8KLtDNPrSyDANHGOKqJw14XdWpwQboVZ5pwm7eMBItSbqUCMZW/77aIT
F1TJ0xnCHsuP0fNZlP09vBR/CorijUGpk+ihJfwxFxKum2qMur+gtd34uEI+W4xe
cjsHQVL7MCMEzqfVtDoojPlmWnM+xOBOgxjGUcktvB4nJkmqAPjWSCyBUbtXxx1g
S06qu/JQ/Xc7NLN0MeB7kSFlPN8+DTZKAR2Z9CbvERJ6Ynt/1OMLnHKTo693XCDQ
YqLo/2R0h60rFzrwb+pMhL/LNvmo29ybj66dcYZEsEMcl9WrYWmzVvEX1E5G6PiX
RABEB/POmVtJzTgAvrpMY+o6HSvkTpBDzpswkVyx1qC7f86ClYSDB5B5BQQoEcyj
U0+2+WGVTGIxET4QDGKgDObnKu5E81qxgZ6+jf1z3t2C7Ny5+BChjCTDNjGQ8ZlC
X37FNGZlz0K8rrcyv1Ee5a2KTrbDuEXuR8xi5N7+IEerygG/nGpce0m9se5WHUjm
vAwtN86P3tbbaE+z7EezF0vHBScJqRe8kXhb0cerNVzdt0jczckrfE8bdJvjwCtg
iZ6y7xF975v92Pk53/OXYoAaTnxr/r4LLb6dTeEyxuATzEp19vSaIuHGd6rQPQ9a
Sezld5vj0bw62yfhXxZY/Q0eeS0LfywT1+FnQsA/nxMmJudU70MNiLHLAA8umEKR
i+XC504VrX4HDWkmoV82C6/rJTvScwT2sEW1oioER0qD7jeiHr5pBHHi6tBL+XSA
cR+OQnp5qiXLjWA7vMXwkUNAPtsjxYVvPcQxcnFkWmX84XM4UX6FOVTUziLTMCPu
L4BZWoRKxaUGQu9mPxeb7mylEjivkzIQ/JrybsKfFMp2bEa6NMXfCF+6ct/4YWof
Qnj1xpiSrgT8bbrnZwspYP6W225ApNq3Vn4q1YChGNCXtLrB/DUxAtKVpcXluNsF
axhsDCehJ7ySHJN9/8Hb2HPC+ZG9JnG76C1Xll5gkmeHBpF1RcaZJgiXcupgOmbl
8EnZF41rbLCh46DLrBtZOPfba375ZweIbHv0zliZaqp81XLSH7+zFBuL0FzlhvKn
4PmvZASR2GwIODQFoY8hoqUdKBw5fAjCz4Lh/+JS0dOzmvCEbYMDxkqZ8ICgSt47
N+Hff7l4Yu46OF+qlqNXq8/DYeYXEYdArK2Wyun/XxyXgjS8qebV52BwaurVPQ+W
/q9yb5Pzi7MDcddOI8CcPI3u8+RR+ZQs4QbM82TgP2lnQ8/lbDH2BCSm9tUi0k8R
7CPYr6zUZdHymqJMP7mw6JjfIDvkEo+tdxhvXyeLmsZkGIi7MvFCeoi6s6YJ59Yp
jyMgguWa5M1Hy4Sw/v8QNL53BI5GPbi4YCuF+iFvoiFu1WWOge4Ew6r80qihl9yP
HjR0PcDWqcLP1WjmIKUpK9OSeHHTLHEHTwB04j2nN6KfKTs2LjjHqM2DLk0z8a5W
g1ukKCicEPxYXXxSvJabp3uV4Eil3npxM7gc2PjP2mD9PFGwd8aC8ebhVvfolkZu
UlK8XisyQ+a1ws50oCI2Uu2xnxEQP1//mWOREX0SP/L4iWxthmSD8TxRA754gVuP
CdWeVrmG5onyWAgJStrFnjwTZ76JVIqVnNVhX/VehXRn2q8yM2szRXG0AEYXt5RG
VqVU8UWOqaES0zXiUnJCFCFI7jebXK8dui6Zls1oZFZCSu5RWj9hsKHbJ43uYXXu
9e99h6tlu9WTSj4+IpsIdLZv8e/345l7O7CD18TVBgu2QPKcb0TRKBX+7FMkSHT2
8NAY0b3WYmFi7L+FhDmvj/YaOgZmKgz4rnrwyPBpEW1nPKYDQ6roXj29va+TyKGR
piIX8pfhQAeVBfllFr9VdV78MziZnBkEIJLxE1OD6PbhfFRTrLTnowc3MRQWTA+z
7Ji8YjWh/Lfp++XmIiDMWIvNmweBSh8whaikjWg5v0G0amxrswoK9r80Ygj1ybiU
9hqaQZZn7IkNxm8WgPCJphIKtpTH0rJ5crFjf+TvoZ3MI598MiFZhnLnYL8Fw4F9
aAZjyYjaL8z/dk/gdSTjD81DKjNSNak2Wv0VWRDQp8MtC3baUxQllRTfoOOpKDHe
FVOtarENVh571w5E/0L9Bv3BlmJUTJRm65puoefb6hAGNsoCm9dTWgV91xW/vxJv
ex5Z7SXi6xrptS9sXGPjXrFjRIu/5Th00svFhcTrXwHoi8rSKWyKaSJUei65dIlS
6QG5/rHDhEeghtrgEx1q1HEwUEUJV9F/qWepqEVZkum7penHacVVqgWiFpuQano4
V2JdcgmOcGUp/yC47QIqt+FZqhz7MEeRMFpuQKwzFncJ1pbrdiHCg7MjGFvOCYJK
SxuVvySpZu1MgMmo6mY+KfyMfBbsXfCrscqTXrjhCZ9cm27YCsv6IducE0KqOY7+
6xbahBr1e+LKKGQJAOBpMUegt+SCq4+y3UUi6/LCPwEiQSGdoVedEGm5JCKTjx6j
GqZguIPpQ1x4AOOufu0/rs/hkvfCjKyi3H2jFT6+3/CvVgzww4ClddybEp9qM8Jh
jpux95L/Xty+RbK5flMOi0On0lipxIoXtXV8FpJsmbhOqF1YbJuhPyrcD+znNyYt
B4yRBJ4xfOTcS0FmvXzv/X83f3HRu/S8IHbAtoBJfsEE1rJ2AnVBReFNz/SVed9u
KA3QFrt0d9u4bwTvTJaM+y8BNSrP0Qk8EvJRdsTHN6XVGwbHP3EFZXb/LRHb/7Zs
gsjWsAIdpdEJ8VaY0JuHKcxvTEO1Ac/zbxk5bvLm96hEt9EF/20x+G4dpuJKup2m
nv/59wrhIrhlHMDFpf46F6Cj0/CIoWOnuMhE68RmObv5kTCWV7VbzMynxRZ2a2DW
ZCVyDAxsRw5VshmaCwjucTkXkz3xYcRlreU4YK/3hX/5imFUS1n3qBXfQ+Vew3uc
ORLxHRWj9D4CioLqzWDgUrms1J0Ck1f3ccxpqwsqHW0sVU5+8O6qB5kxQ/RuwKro
VkHJzdUBNn9Ep17BcBnaFTkm/NUHSAqSUNc6GHLQgrUD97VGupKvgzjJ2GV/nRPW
Cxria6954OSPqQAm3igdpEUpGDW/FShDETINoTTuOOPRmjTc9O+19FzfHT5pJ4+r
pj3DUISRDFk20dy8DmLysH4No08TpgImpxdn6Ujx5Rg4LX9n+l1VNEWbjfW5njVC
hRwDgGa8zTX+bBNDH6g+/HDXdJw1aaMbomM8/oY4a2jElNODH1I6nRLLLJScrTt4
OYuKgAYndDzZhETER/3x9BS7QWxfiNMQVLmyxFIBprDqjp9rugyqHf1/Wi0p+Z8c
B3u/1ijRHRacA4Rlnd/oZDJvL9ggECHT8WhD1L6ofy9D5O84SFKWklLVozZJtVVa
Qr3ZbJDHHyNi9q8M+ay+orXwFXNWrrAnDn7lh3y2t+8/ltaIYmNXf3acPrsPvTt6
Ap9zAhh3VP/yaPrJkYnvR4IvZ0O0vPIWeBWbIZc0xjA6SuEcsMZjzi0pxYtN1jcJ
eEGhNxRNcC2W7tg0TMb+4xNzmpfQQBu8JhhVdnYIQonl+GDwGtjc8EZ93LXDotn0
LwU0Cfa4RNYyOrhfpoqKBkJ79y7VCo/TOfD+a2KwYS+Oma4WMsdAF0Be9O8PZtRg
hfQrhs8WSzL3oeZfVMGa++z0Juw8dCkMgitnfznuap8zhfQO+sfICC5viuQyjdtv
uIUxC7F7pWL4rNWyo0ZTp9LNpYOB9/ruZnTDkusFhQeFqklnD5wEr3qSvIAXRWbV
SBJ3xZB+ZgmOfqOlY++836xu6N79krS2yhFZYLipD7FZcroE1gEdDchf9K5Pfo6Q
cOgDVzIFiTCAecllGsoKXXSJAiBkIxoxiGpDr0C2VJuArGQFcZpenjlkCpYLjpnk
rl4mX/zcCQ1nwouyunrGlwvlzYAu383c5yTydyqau/P8MDvWLNRkWzpe5r2NpP4z
+qBpbxV4WFKuUai2KdRRlYKNOkbXZUbC4kt1kkRBXxQ73+Cu6QxIjWxASGsIx1Uc
XoWgdBrkACOR2TirFnnaiOKWyKedtWoh+/x9A6sn2znPSrSEPKXMDPy61V7neGH3
w6ucnDhMFydin9Fw0vGZK7lu4HZ7iieYcY8DhoIlw0gEgTDjikcduECPoAcZl7eJ
4UiHmguMrpKcjYoxAijBDWu1pdAoZ/N/8jd7mzay4pXYNiC20QICt824IrwG3s2N
Q1vY14xLPVlFZdu8Ak8a3n1o1nEiHXbgrRdf3A2cVqDDcGnyBcQPK+/8TOpYEOx9
KCMhu8CUSCvfDosJPmirBxXLa4x1JzItuFixYPI1cqwNZWFRBAZaMaYKHOgG+tHL
Er0hk0cu4bzNlqFar2jaHbt6e6wPjnVwMQToJe23TOwk6yQ5mudCgGBJkaG499ix
Hfv6tVr5nAV58pNi7quoMbcpVkNW7lCz2K94OsLc6nEUMx5atJ4OVPLVt4UPgRDC
RX1tlPURRjN3kiPUAN6oJhYAqFR4dYnKZ5zc/R6P+41Dimjjn/RHk5AP10gAgRgk
y1Z04/PF4zyt+wtL4FMde8oyKilcyCbO+rdd0II4XHVtXWg5+v25724iYz6qgN34
aeMhL17KFw/ulwXLcOpNapQLadZfuloF1/ICAR+ygLYqDgx+MA0T0JbENPA29gUO
l7V0MPOieUlGpi3TUOxKVyyQjZ4lbmONKiEShylfF7irj4XLMx+peeqcBFmZJUk9
oV6OUpgP6CBe/h2xUb+FaiOgY/GSFc4X9Ut2EjlUpbh9Z2NpkHWsn7NvKzoNJ6ke
jK3RSfgBwTCfxOu1VdK9ToskyVlrQZ5TeTLIkAe2VqluLAlQIq3Hg09/YRVWnhRk
BXZBz6YWDkIMzIUp1QvNwxV0S7jDUU8t9jo0wfs3dmd8ku774MZx2oyfDaCI6FkJ
PGtR3OWRartUDEQCs4IxEXoGgh0HPoR2fSx6uWDRz2EG0TWlrqWkmYbbp72YRLlv
YgoK7smzP+i69NwemUfzduNomvMyOyL3ie6/hFnvQaVkOS/FUbC3i3ApiPLYaLM6
rcC+Enw2RmSVctq9/UWrvOjv63QCk1nFaYHMzHO6Uz9vl0ff+St03LMoUiAFobLj
YPjfNnkDXUOQFvPbbX2Lnaw7dic5y3nj1eXpXh7TUFueChWhEgnaB/tgftgnJbNH
Rzv6jxWOgP8HKfhhVs/Smh9GzWIgOS6wBEVDpsjFpm/mQ1CY1qhJ+jbbL4LZRMnA
A7zPjPbrcLaTglS8XUAfbUJOeK6xEv2+9K2/YA+9P1T6nIEBPrWzNpZ03vQlP+eH
KpNIRpFUKNjNjCMqpMWtNvuJOKPuWMlXICEB4QNu0Fd29PJ1vAIYZbGO2w02DXXi
k4ib47WM4yXEL5ti8Z82U2JSNNbvI4y8mou0G1IorkdQc6FA+/mD0WNPPeShJDlW
3ldY05eudrGPyiCf+/dThCz/X4d9jm8KoBHk9IApgsWPHU8ixCtyY/O0bay9Ssql
tF8HQb6mqirCLnKjcwUMinnCVh7GOmSef1TygTnnwx5dDMO8F4PkrVN/CAvyfxNO
yS4hcYv8ajAOolAu6GWwHu6mRB8FSuBLf3sbaf5B1nvSd/nhT6BUTpcdNqymhcZD
KPveZk0bP3jjmNSN0u2jjWjybgaKAR288YV5tGEuneq3xRsQQDgLGqg9PsbhjHqd
1ooh2mbEzCZJeZyx6yOc7Ruyoi7kiGJnzjm3xxV0OhKcA6MbmX2FDstf8cMKKPZR
TuTipC0C5ctqfBRnGQqeNsVSYTt8mj5tIt8KWsEOY8h382HvqjObUPYpUOmeMzY0
kDdyuHcFTJrFkK6X7C/vu8RHSK1/tQWv+SnAbPZD2C2AlcEr9rznPzngX24Dk8n5
q+N/AFsUbIzE9SCnx7Q14CkSHLbAq8evAGSPBqwJz9jGlPw0oqYgHg/tBZzoMPJr
1+m94HeipaGRSaT3QY/eSNwSxQdFdgjlrsRcUkbnX6B13ZDCx9rI0Q+/z6MSx94J
deamJpsYOEkyGFifCJ+/M+PDGCB0+k9Tr5pUpriJir79qc6MPdQu/s21RyeOsyKE
69etj+D2a7LjCmBA7GJYvCJ3TwM5gk2LJz8WRrm8TQG3lQtuKoMdEzduhPaAlNBD
nWoy3GKS7yVb6y9np+1cIMDjtCT8icVt9YUI8+x5Xl6MAESYJX6qrp5XxTIZswIw
UaoWCPWlrWAX5Vd69WNjTqToSjzkMMs0S6ytyXG9+oVbp02rPT4u1JUJaraiIhr4
uxZdXteUwydbEKtdNdyIwPHIvgqLpu04vSt2McDBfbf6wfvJd17mqvK5CNKtOOkY
aXXD8bH7ZiPlBV7XN3SwmNpn7DPEeWWrhK8xsoNuK/LBFtSRw9b4mYLbNWqta7Vn
gRxBwXAUQGMAB/oPGVs44UCJOlDtqNa2hsqL5YeB8ESSH75XS4f+9pCZRU63Z/vU
wyZ9yH7u305acWHFDwG3TArt4TNnTPNkP4PIowMAl9UcWwASsfVc/f/nQ/ls5jk/
+6qFCePlMI0YmcO8pJHjSXx4ICDjQ6sW+no+OqCSaRBDts/0KG656Gdd3A+RyyOn
rEz+q5qjMtVKlKQpzl51aCa7tkt5k6IIK0AzEUhjhg/+rGylSHlaaS2yoX17CsfE
gUqVmroLjHAKtwEDa7TKwCIympTVq1GhaDS5Ce0aum4uUGioeNldJ7eBl3tQmqlk
11vfS0dIVKcOvQbZYBlEBth6MkiG0x8DXFljCtXX4UbMWyLtnaX5UNUfH0U1xtcq
Euxp8oxXvd55cjtzK+F6x5o9iZWqP5ikUNLpAyNpO8wCgaGhLvU5mGVfQHuhJs9g
2NsOgkWs/WLW5sajCHHMrfVCPUJUBA6BufcsguXvUuwpDJNjmyoSzWunomWAFzgJ
pQDWoJcGIIXbK+mbJoJ2RoQKQrsSvrS23WnqWOqTm4s/M3gB9elyltbvJ9wa9m7O
2akR6lMIrAAqfhxV2ccPAiOuVcCp3v0dVKnHAnPATVQdeAfIHg9RVfA0NlwR5153
zyWLYyImUU7hbLiE1/U2bxmk4MEY5x1pfMnhwGEfjwwRThe7rMVhWOUa/FQPJhnh
pQIpr5IcI5rG/qCWuMse6HjFH9FXJu49NPWKAu8k7jcDm04yxZLUmPdYqBvF0KRu
hXUGd7hNczHoF4a8Vk/JbE96SVmva0Lvx8WCENbmjNvAnHtp65yUPNwxYjFKlCXS
tvTEMaMkh51A9cMCda+cIQQlgBb7F+bn9EJEiqVTy8CIPbY+f+NW6oVJSLzTxaB2
/PWrMX6JNTL8gE9sAxqYqQLvRWQHXN5SVFydepYthMqA1deIqQ1ri5axxgoLgM2Q
M+CQS2QYdxD6y783KUun6MxBl5YWe9DFN+VxnL4IMDe2ppzjaoPpSdl2WzBWeuMq
nDlpNQ4QV7MgJ/yiECMocjkf6NbT66js3ELY4Ug19aAFQVhEVSdQd9otKgBSpnaX
rgar1dGmJNrDz8iKFlYD+zxME8QzpZxdhmBx9M/jMaLi95tHOEvFtMElRfcncdtY
F5VSKpy2iy83IgM3+yqDGrKOSNP7BPId0QfronUINfvFoHXp42v5AAvpiM5sqCfY
yAWDVaatxc9ttnEboDMagU+MU/JFCo4wWji6+Yw82mNvNgIHK/eA44EhH2GIO2V0
RnhVADNzWTmit0YO/+RqOYRAorfjMyalxqAwAIdisMY/UnC/PRfoNkE2UqFYrM8o
UssBLolK8lXFtD6HDPRBkHZcDd6GXhgj12vN7zL5KMfy8m3Lr0QN0hhES7RXZmXk
qOOYlZ+kWwsqxI8XnKCUpe7+tlZNr36O4RkgAI6ty5rDgSTC8K7ClCCYB5gYyWCn
YtKEN6OUCK3wGL5rdSZmyYfeebHQ8bM2rVck81hG2cDmKElsCG7PruTsxoQytLe9
jDV6QOlP9jIpuVsP0zMDvrf+H20lW+X+N6JpONgNChGFgJHQoVwKDZ2x14A6sMZq
SsQc59qW9mzratqpXeQ++ckLHKsn0/tpMxCq9Kb5dLw8sUeeK784jS+AMg6MR2R+
iEFsyc3sppqXn2MPBOrhaWi37dsl3HPOEtHz5ngiOJ5o4FHh4IIhGMfV98J6/3MG
Wl7sazyBoYbI45nH72Tsfi1RWf8i58rrhzGiY4OlfiZdsRKkPTF4l1KqiTtYsnwb
P2NHQf8v76qskt9P6RcpurO2aAf/ejPWILLzvYVLVkCIApJe6P4aGt8uei8Gayjd
Ski3vPBQJ6lVDi845poehzC+Z2PlQXiJGCCDjqh/s/ZstlqzfIlcuDBIxynUzPT5
17JnQkP+7MuE54diYvUd/tzYitxOSdQHFk3Phst0KiljUudyzxGkjW/Q7rspjNpP
UM5rfP40NhjUoO66ZiD0ajuU7flHUKqiTHsltMu/syyiRNY0Ghpn7YzcOJ/7uOnc
LBSIYcyuGjcqcRtEi0QUUs8y0f8x29O241hjY+4G4/HktzcfQnzFcTJ03eKyfLfK
/nIBvOuaZH5c7Un4ri8nVxcICRCFe9SfduwBVUkcnsiyWh6LOlWAODxbcTZvAodn
bV93Q8W0pH8/YCuBWBftbR9UfHv6eGXRN5i+GuDgJ8YFiryqfJh2Soz38C3EBNvs
OkV6nlkhKYKGbiG3wy9Q9NREVbSf3ZKDvIAv0PKQzmHSajRqe3KB/67vjQXCWkA6
17sKOmGwemcrVESHCiDNta1U7EdYvgMHdS7uFzGQpxWnok1NWp2HFQDtU1a5hAfI
xVawT+1kR91uEkFqiptN7ryxEp1NlxQS9UydsQe2ShXv7uFlYrExPtIMOLNvCltB
dyPziNXQfPG1zCQHex3z6I5fF7aC8GyIM6HwOmIUNrxbGtKi0KzTCSHfbEyYM6Kq
m4YboA/xF4h06KFDiT2v4tP8U9UtPlbqyFuK2Vfng5bh5OnBxRHZSyEFyUsEKB5x
atqcpap7fzY3VGvbo1gC8J1SfpWGqqmPlAlbU7/MGCbkDMmlJvWdObv1g1i2Tzqb
XMDV8Ir3VLTKv/pdc+Y0bhwiARY453BybkmuycNAmr8x33o4khYte5o22DUMp4iU
vVIKlyxMV7mZUMZzzetaQ+rOBYqktEb4ZvMegyif/zNF1bsRkabY7TSI9fixw2EA
/zJLTPsatz70qwKyO3rM0ESlSNkUpYBsEogOUfJLj83nJht4ozttrhszd+sKgkKr
JxqVA0Z3H06M1PTTqsyQp1BpvZaJ9z1m/u+Nw+u+CkKE5xkEgdzm5uMXxK9NLmcT
e+jJHxzqVf7wQlUMAcfYYhDvRpAk3clIxjJ4baOhgKAYnZJmnqXKSOTgcq0+6KhM
KrvkfqKUM3M0RIrb0kFXtICjvri8WcVRgNjbvJWnKICKH/FMFqk/9ag0Bffp9xlG
f33AlRbENiH3io3lhDEa8gxUi7by+n5YDb3/VyBT/rlPz94NSlI4LXf7AyA67/Ye
ImN19fYFSOVIy5cH85kv0XFNNUfhjQsdBtn/MQDZE5K/QLhvyLRzgqwr4XoXQ+Xl
mq+hnM4bzx82t+PM0wCQwZP0g7e/1saEVe3vK4z/ol1RK1O85oGKBvMF3rRq/m/D
toZC/cA0nQmz6vw0jy86CuIy2MnpWmrmoQGq1B/3/OO/AEnJpLXxkyiIfYYH0NTX
dS68Cbx2g48PYJ7RC+0YEkbipL5JMASWHY9NbOMNm1irmc4Os9DboRgtNxIV5TXT
3DGMyY2dtBMA/vtEf6zJTkMi34euMtSZXwORpIS1mdIiy4YA/CjRlcykqO7J9hUR
dCdK7+1fAs1VcifuQQfHHnQ17wWJ7t+3wgqXSeAiSQFzk/H6txyid2+6uGmmKIYF
ugKeFr1eU50I5NttT7mHwdqKitS/rMV4RZLjITpBi1T9/11Bx1diBObQtb9VGyo2
DR/Z0XSLf3tBhrGsRvLnWYZEIZSmz1O79OdTPTaspcySVdq4wZyxScFyc17Oc75j
rBfddY5jgciZ+TQ3N7XFHI7eWsLrUIsz7Fof3Ck1zgOzPXEAJ0ICjHkk0r7NoDFN
Je9R6ZuKK5EY2AnXSuE3m1Q6aAqpAhEt4cHBMMbsq4VMbuFR+8Xj5vTYH1oXP3FF
2h1VKhek8gDC/lKqA2Q1DersUh8jHeHoaeAH6z7dIzyy28JJ/i6cxSFUv8YSiVDZ
4+95fARQ56qNDlBvvfDwReCrh7Ljv1KaQOr57L4iZYTFPk9Dwb+GiQpGgTCxFH/1
rVWh7yDXGnErHay8xqVLdQaAnXDX44f0s761b6gg9nSt4r/aPAPmO3AIurULetoI
jz1HqMqJ4ypdGAnUdZZkrB3QARek4sLzY/gJ8EQMjkG/7s7WfwfwbsYO0v3irL76
DQ1NeMtQpsAFk5ikuxVOct/5AoVJ8UR0a0YtqI/bDuYk0ZfnlIa9yUEj7R+ZWvgK
vkmaZQhkX2DsqOE0hJg5BJVbETyzZ7prJz+4WTEat8BWNctIZ9okGJ6Ss9SUOJBv
51m9gghSxOb46mLCPzVw5Xmd7boPLdc2pfuEmKbpCmwUEK84MjtfQtur0jyBZWeB
OYSIbPPGmrb9/kZnUo8q0UDmaQzHyjQ1spaoqvN9kL5YCH7Qp9XaLy4eROEW8DvC
cJgycpLqjDHmkBkV3L4zWq8r7SGk4BF1B/sC15wSBZ16bQXi9mntXEXBQeYgH5Y0
34VZi9d8dGg+CC40orVSvoSdKlHMyUB8UxV+pHl0mcDfRQlmZsvUH25vzmkex2wV
uXt3Vs44GyFDufpRq8eUgqqL2T31ORyJVjKZKKMJHK3LlHRxy6E+aHpY+NB5pjAS
rWWTJHbwqgThYJ+GBe0M85j0ZCYhYLZlHJOfXL5Z3Vk9gK0G2MWIQNU2DjcepGc5
FICBP40zajPPtqC2/HndPmlxgBkSH8KQF4BY+DfJk2kI+dC1WUSOIIam9ieI7B3I
ynA1D6COskGaLQ8p0FI7Zf/Kb9aQ0y2z0dDrdGlsdjnF8Z5WzNz5EIUTKGqnJWcE
B1lWuiWX+8eXgpU12FJmCVawpfdNDVX1KvMmyhuh6Xwvs1gJWg6vrBqecBp5xco4
7ifYe0gku6pHvN5J+3t0z+MOqI5rtzZH3vVfUKgCNWjx4ykjyZnjzm0U9TrzrCN0
EoKI2IuzQ2wiBt/+fLdFYGmcVJtVmohjDftopkYkkKqgWJUCad3eSs4egXfhSxjS
zx6ZnkPd9Lm6FxANj69WA9i/wk75WC4atTPwUsAd31Q2LIheF0o7OIxSbb1MtlFk
mW8FWqH8K5vyFUgFhUJZ6cIEHY7mk+U7FiNAJ82j/ij/m/5LV4OI5s0oYU7jZhDJ
/Rl6Q17XuC2ogzDzyuz8kGa0doM2DacD+K/00wO/Wsetuql//WuRmSJ292V6qPaC
7sJyiq/ZP+5tXF7aCWFQVuPb2EsKcrvUzjrUvLbvjEyN9wdQnY9ueLpFEo/a33Ys
1eSYWq+Fw2TPdGq4frLFpTyXQXOdFq4ajyjG0Z/O/JdkZgkJTBBx9Jps9OU4pQhG
1N2xqpfcKORzq6yp9kol0IL8/SKrW/bkmh7+YMkdvB3AUHijCYNcvOQuPx91/8Nu
rbtckrl6l/nMCWdnYrhBmet99CDcIj0zvtOqGXsVwjUnrire0abCYTlnMhycKzOg
hZ10ofUHs46V1iJTrOVl+irakd+XqBUBWAEOgDpb3lGljK5Z2ttQ16pBu1TPYi2u
U7vWrrBi8bt2LzFOTd6Gnk4fLHTzXwQ9WGPdV1gPWFKOKnYvCO26gFXc/W28Lq4U
8PaH4neEL6jTBhxQfvHfDlLjOJBNtEW3sIVxR8XZ1GNXh2T6vocwOzzlYoIoOqxL
+plex+BMu/7BqLaxa3Y4jrKMTmC0hJphHleRZhXTXWbs+3/syUz8iiEv+lS8RLDc
tyUf5P6Mm/iUuWAfTC2ox2cxPljMbg7RRGeOjVxY4T/NdFQnEAozdB+VoEOikyo7
iZi1IGIYh7zrxuHRLuzmcq3HG+fcZdmaNA7m4ZX9OcfV+9ZvahFBxUUO3x5aqsMs
cWiP6tKRWzWm1DATBo2CkLhJW3C5vHMzFGuQfeyzFmIiiG0PG+MwvaRIJeTYgF+F
bWgVlCP0kEFMDheY92tJNToHYVlROU9hhecof7YE9g/oip1CsvGC9eteDQH58jqF
JdhDKvFJcBK1W4fHFa49BlqBsVVELcu5aOAQ/2dAZBgy29zs5DtSfM7oDFkGYrVx
Ce3WnjuwIumtvmdYhi275qN1+gRLjkjW2OWKdXdYpQmPUk/MS50PWf0qOWineeLM
nrLmNG/SQO5DfsoP2+ucP5dHnquCwL3xANdHakx+wotBLIK4KScnDGJl95y9wK71
ASReoW58uJ9mNu3zudMIZNdOfSEZMpWvhjd8CIfqpPswYk74z6uzUG9KfGqNDhIM
rqB/t+EvcvYo5sQSDRXuwKgjeCIuhGw1pd3QpTuc7gQdkClNK3iFpRuyZWHMoMLj
BLq9UTC8QCpxRCW+2HxldELY65qyVBo1E3yEk1fGgd7LegaJ3CbSf71YblFNzyAL
csoeVEhgLtptmH85UPu6qLFILvzgyfEbJvS/xIElzzZtcfE/7GeGPX/u9PHZQ1Gc
0sxVAOdrmK3WYQyf0Yw97BuaBahWrCJ1DMgExJlR6l56toIu0ENcO/eV4T3BA+1f
J42UkYrs+LDxA5oDDsgi+NyQdGCjYiUk/CvvHTXc2kevkmJOTqaa+HNhRHLfTYyI
xdcy+tnsoTcvY41A1LnZGoGmtLG4O2dC9fBOPeFQS0lpy343D7ukCJA/BNM+dw6j
w/BGaubHqHUnlfWK/xjiMzdWpXZGlRQF4wOj992kauZREWRVvONM/qq8+dLm3qEH
ITYhkTz4o8ijl1Gpahd9K6Sb7oIjfGtJ2vbvSp49QDqiBOLFFY4+fRuMHM9Jgb0m
SrzYW970ZCTS/zf0QzFX2szlAiGLorHnO55jythwMe8fyso9GkQKnvpjXFAx0s2T
Cg7JY8SIJgfj23HcQttm6ToVD/gaa4dPM/z4ctHe8rxUe1hlu0C2v+t5d/Lludbm
tqFtuSUQtK3EF6GqkDIYrQdq+DhFm3TUDvMgA8Fp2jYAxxY25AEjD99tVCe1qYtb
OrnQpYD8pYYdHUVP0/QgO8ihejNYCKs93MnHvQEU08zlXucYkBwpeo/oHRCc4IR2
bowP0A1qRtkN8Adb68y5V7a9RiNNI1upUK6SqvPnCdfd0+LmFx60GQgY0OFPalKY
YVh6xVD3+w0dhGpgosVDN69tEI9eorfDjbszHRSIUUl13+1DfljJf0+YGW2eXE1U
S+EzhiqtprZq7WnJA6qTwYTncdbd7Z6Wynk/B3WxkvGouF6dPIGQ5otXVsw7y7SJ
7fK58w5oeVnDBDWJVfwfe9edzU84TAGJ8MrTgns/vYry9xoachrypA6C35d/L7+y
nJHccov1S8ihdJfVCxQqUhdzPj/QpytXOitI64Tgsi9nkNGYNyiX2vxoC3u6tGei
IOxXqmDxM+OONc/wcZwZwJEHE7xXsZHcgGpUQqUKHPvmfKl205PLRHeXBV+XqfPw
FRI7LDFX2o02turGpGwlyDydoIcahjFpF4FWcDo5HUMWipDiI3nSZbU9qanmDPHl
ycIxrnkk/1EHG5xiesBXHzpH+lH7CKXNURG66NW//mPXA7iiT76d+B5d+2mDvNvY
l7lyC/IwOocJFu+KNW/tqZGCyV9GDoYjhU5sbYiKdDyA6I1K/eIILW7dyKcmkOmm
3OpaZ8x2GSVp/zWyxbGGpzVj3orOYzx5T81opE1N/u9qPLGmyPWs48rNUh5D3chC
DA4XiJQZVNHD/Uo4bepOTA6l2BM1yU7lV+49r014FkGyR/ZS8qRUaRX/ntDuxLGE
Tjdzrv218Mg5PsThm8nQtP3fme3u+lY7ztFNd547a3r418xo/N3RbqXNn6uWqVLg
jGHl6VOAtXyCMvI2c/JQmKMwvKUYf3/+7LkLrL+OjFriEheixXn7sPFg1wJ2xIct
jyW0KWziiSjIs81q7csMAzADS5S1W7flErywRc/Mav4Xl7GhHZd8aAWVrFUuJKsk
01o+Gv4dgpzXoEJIV0zkVk8ycz6tEZQRsWyaOchf3W+NCCYak8RZX/HZ0u67mPL0
DlMsE+nL60ZWOZyOSE5FLO+4PL2G7UCQXElEl1kuwRrGVHju+l7DeQCUED7meX9s
78tLiNpsreTt8f/CmrozbUOTWUvzlsRffuWhKQ928FgcJJfV/7fu4NZKQdnzrjXi
prXlrgwSQn1W+ICxm1yOHtZ5QHpFoCRqQ5xK+vkIIlrVOtMpcmsxBVHxVEI8zVpI
Urs7vIW4iUYMDinyZ3OslJZf8iAZyHdMmyz20ncbi4Ajrj4p0CHG0l3qjIFpO+dz
Vls3baouOvlP7CgByr6xeopBn7Z6psOckUr6FwRJl44VgeSv8g8TjBO+zHI2G7cc
z4i+CBhCoLp6GefZesXgyiZ47r07lyGo0EEeGh3sm2zmZAA4hLPyXbGb+MYJJJ7U
E8nLEF810LOZrHVq5XEOKjNf/yWFC3YbOmvLqad6i1P+/ompbnBWUYQOpcSZmLFe
m7UTlciNfXeZ+c9+LZt3hmpSud2VHg/ft04I+LGC05J/jEZAyYxBeLvLySt+Ojk9
dHtclYFEsOQrwDSADHJBhc3KV8a/fokzzR0IEOi59vVRbGUG/g16yr4jxSMz9AAS
0VtTasEFDdCerJiz5FvA+5COs4kZBqNoTzXEOyPuhmU+BgMZIH9VsmOhxVeinBvQ
9rc45UHpnvBRyd4CEbOdj49z87mJ5K5ICYqnp1D/kI7Oj46yp07JgqB72K28oQFd
gqAb/Ytf/yp6IOKer70CdD9P42nLi2F6nHrW/iYrOfLBfQL9ijOivIRYuVIZZ2wv
7kCqrKeyumVIYPvm/yfLHGMp1u9aq4pxHh6AOTfZv1Nn4lyRvL446RK2dzz+iJUu
ZGAkya2QKOmUDZ68h/+nBL55IwMwHkhL+34R5ZGy4Poc7/xPqoCJhD77e4SeoWzq
sHCRc04HyBOSgr0ltc5lJRkx46h5ZPRY+wyVIJr75vzkVkvyjIszXcC8alsGdPLU
uDxLGKCH054XapVSBUZNO7Tb81rs7Mi+qkE/8NMUGadtJ95Wy+RMvpBYj4NjstA6
wDyBDsOCNcQlgasdVLp/cdi/57lwkJhmTnk9OQTdtcXhCttpkAVm7jjTthzdAq1z
Lkewu+DhZgIv27UEvoIscM8XQbM8OYcUGWf6b3RecTK2vccdWjiWgO+zUcP6WsD1
xJjnCFYVTye+hWI4yJ+nOcythdVlzj4kKJ5/4hgedztQLGz4ijx3G0a274AawZvy
lufREcsPDgrvC2Zu3xAknGPKCwwTBZVBMXppwvzzs9+Nh0U3ezkFnLazWKwPEuzi
ENtmML8uJ2frT7c+EtMgqYUuoomY0WyvXRAUPjzkfMLEReL2dElJZWwTZa5+tcj4
S1MBraanLl+XGb7/7+ShLQwr7TSGP1McMl954H//6+1Bwr1K8ZpumlbaNF4rT17L
0JNJqzn4XKWxOdKfWvded/HQFKs4IQBu5WxWtWpi1lBQOHCSRcgBQmB1D+PjvSPE
KPNuwKrQc/VIWw5s2JFaiPWGRkV8wzegs9bWORi3IzyfXobjb/Q563fxHtIucliU
GiwYtYVtunwbOPU61LoJCPACYinvkL9PIKF1DySbJ3HmCK6QaIgmj+uMGXYfDnqW
eW6LUHDE2/OEHNE+gDr9ivKKMfIBWGfSKXDixxsbVxmbbZR+P3TZv1LgSO+TrwbV
G2nQ2ByJFgapYLoJIzkyqJiYN/b/AoTG2GpgNsDqNy4YZcqyBO+hLn7v9cdLsKrP
MEeyKs0bn1y1ACBl1M7lOyj97cNzeRB/zGy6UUT/LfXlnp99r9+PzisZOdw7brO8
GTLd7b8xOzW62MVLgB1JoR5uA/BfI0a5WZSsEiKkKmdhlCPrFOuOUlDBT0n+noPL
JA8zCKd0r8MY9wbDHu3h2oeuiHFspD+PoXo6xuOYNvvNNvho+JDeIDdgtCIpsB/G
mY2Ichk14eAcwY3Oxkx6BJzhwgG5Jjh129Z5B+SyhSE4TwVo2ypnZs4pF7z9TGFE
Cz0hFevOSaB8UJECBWmzCfKxIjIk6AF4aFc7A0ck/+a2etS6Rrex18eI4ngE8cR0
R9WXCjocoTWXpY6LdyGhG3pKUPbG5bxXwmRavGm4xSH4nOIj+R9beCDZWJEkN7ys
WyG9Zi0g0v1zVrCRBxW7xVxMGUak2HgFjkE7o1YP7YIMGfeUa1xIRWs39dafkO1w
5oVPb6I071gENYqAh77SuxFgMYavrv2W0MH3Z17CBqvJ9Ox17Atir4jjUlRrjcEe
ZX4FEN2miaPrHbqxPNOQOZJJaJOJTW1UV5inoa4mpDSnphBHoYwtcju637JmQJ2w
TrHtZx839UAclVn6lOw8QJPeOY6/2UYnBljAOaFRXwcPH01E2mfwxbkn+odO/dWF
kCCCtRghZqoonR6lJ+6MSAAd+oLs2p/pPwUeASvXQ1nQfWB4oghQOqzLxIUoaR2n
pEZvisdjDkwNfJ1WviCrafgRzqhQdyu9ZbVyZr6cBLy2RbKskkP2MiH5bZ9uqo5q
uIC+c/eeLKd8YSZEC7ERXYlLN4W6isKXGjGrVwp23RtECLg8ikCH6qfqU6ZmmcVh
3o0pFDFMaN4fKEkWpjdrWfmev6xuRg19RWPHNbq8XaheXChFNTnu69TN+43s2Mdt
qVKp1b7zPY/S0G39eoOQ9N7LK3czMefe91+MqlPRsG8wIp5UC/NqmMQtvOeN0N13
kRSUMYRvKQvWnQcu4361K47rndUi8BIHmFQhAJUjH2cVghnVPg6OMvZ9M3245qd6
4uhHlQDFo4by7mWy91hCvYFyq0fcBNK63O31jrGwBZp23TSakK80sBLVqiWgxRGj
7AUb9ypB9REM4E4c4Y4xt8fPv5j2sgJlBFOO9dPBR2UDOfbTciel7T75bK9FaJm5
QfMO+TZTNEQ4qbawt1s2OLL0HdX9h65WRwHb+LgmK7Qvb4F79XCq6GGvzWr3FIg4
AzxKZxBpSWIwt9qbrt9QqNq1q0UjZB10DLnH5e+0LoQXEqAkLoXFayVdA8zW80eY
NmqMO7vSXplG9eC1PNwYBzMvzJ/AoYVzyDfocMXR4/sUqiWrm6Ww767QJvcYZenf
fw5WmKreT81ZS9Fd20WnsW/VRCy/UfEQdEdWWndWEKCMkKGeA/QFi3uY7z5Pwmyc
9upKzD84rLQUItBWvK5JmVovTu7v0sKrlno42NtVSOz/3UBwNNNlJY3EpG3yGVUp
5PcZIjf7kgNxS+P3VAloKRIFUCA5nIYtSDEQNZODhFiC7KbjcusRudD+SVeTwCMq
K5sAodtpiRm4bKmHnWcEx3rfUBM17QffHelZ08sx+BiDWm4k/D1Tp4R8LortNnye
/t1JklYnnJYWoLV/HHW/VsP683mpULxydBz2VBAN33NnIuAqSbjkk7Y5QpCV9G2u
L84LRkidDdHFa3BBx2PQnXWbpxhQ7KjY6WJ5B2i4zmcjo71SlUMYN4fw1CGliTRN
g2BNOzylqTrbH+LruvvbRmQoOXoviD7IvMf+e2RlvItNP4Wf23uUv8ZH7k5VNZlz
UJd6QhZlLgEmbab7ErnZI7LTmTCXC+HpnYLCZCZYt5fShZBM66W+PufHfM6KZP0u
jSAr2RJ0002wERY5JJb11mNJ3VJk9YqzAHSQGIHRM3V9j/qyUO34FONPPFJlnOt4
PTY2nHp9GbP6rWKgwfaadMSMsi2goLzNqVcY8Sm2naIhOlR/W7opiIa3itQQCMEV
xj6XIim2JMLaeS8Ov8g7KX+D29hMvkUlsfbJlt8S1H/GcYpgAaTgJeKuKAVFZ1e6
0KfLrOHHENEPHNptmvjQC7C1xzM7cSFeryLtEsvnTS4zhrwBk1atelCDTQ9Pd4jk
I5iXthxSyv2gAVrYbDzWB1ZSZCVHVIytGvwZqbDXsYH2r+LVCXi4/GWKxGEPzfnP
UIrMH7drsRcVnP60/0unm0ukqwR9xN+dWKJBAbtSRZq4Auvosn2CuByr+RxfG2iF
G7NobFLvRlB7mTpMwBhQPMgIeEoZ956FSdUtSvnSGKqXeZx8R3CK1KDi3//x72xb
p2uLWnwW6YXtOZvyzxjC0raG0CvZOw309WLxGD9aXZoeF7EuFwm31JDc1+TVvOB6
8YmX+TKP4jy0UiEOcasQPwsx+Po28KuFnKs051sYXY6QdxJME9TrMbhpDaszz/ty
Ak0AtXqyQmAesc/dSuiK81JWCcU2W850kgZXDJ7y753p6I7nvZoYMhxImlCJLkkT
VxydHnNX4XyMD87tNU7rVOV65yA9ffXU9osnX3oaPukAv8Zh9ENgPqo+EKJ8AjHK
39CKsHMYY2l93PBRu5ai/SvF93v33U3CRdAGQEGBFkNd813YNuRpz7ze76PdCJ6F
VdUQbV2ZPhC2LdFKUvkcULhivGge1kjX8xsPNIMwa5E/qk5y+KE1QLgGrki4ewXB
g3NN6ip1w5A70ynEcYdymBWgI6c59RoZOmIkjsee/dPFAPPmqI7EicuhTO7JAOmO
PiPlujtmiekR/CapCQILOe4wvI+s2xqGdU+tC2ycqAfHo1D7ldbg/1yCRI2KGdN0
C77EGoblkKOEJrZbQx+LEGg1IAZV5eYHWlCInV//Mh79v3kzIlFBiklUkvNQrekJ
GYdi0zguwYoqzhM31pISxpPymTgtEaHve+fA//MfnAmxTjOPkF6+hd4s2OhCmhmo
biP4dKRJJG8wazD6LRiy9VVCcB+MSmcMbnx2SBtBHS6Sc6zzggXRH7DbzOM3wssO
F14A5mGcqGho1m/Y9DLi7OHnJDgGhWxYa0K9Jbvy9B/H968S1s3AoDBcH8I0EeCe
9xLdmKK0L5Dtk/h+jrLar/P1mSaODAsEiTriF5551DiZAW0GJ4zKs4YEaNQsLinv
mYHiHXSQD9ayoTrZ3/YYasiJEP7bxVAd8AOE8Qb0roUSkiikDjwZbxs2nQLi4ha/
jkNuvrGYs2KA90vmA0RvUhd0mkohDO4czm//bGBYPmgc7bDZmhy23W48jCgEy7/1
2iAvkfQccscz6Qox5IHm7uS+EG8R+niOvcvcY4CI8CMcqSXQbXOHd6Ct3V2NxI5z
TquCml2THN3Kj1oNFCDBprhgJfrE0zd/YluVrnBXlfeDrXiq5a7MqsuYQNvLY2AZ
aSe74rkvcZSclbvkS9Ci4xmo2uQkfojcF33UILEP11MlIZxUoZDiabOLb56hdFlL
0n844QU1p3RBf43Fb88HiH3ylxIZtuAPB3YBJ6VzNRoV11zM8oZp6RPCGp+l2RyE
78hRANq0VjAyewjokrQqtDc+tDWf2AJwkDjNq12gd2Spr5DheXqM0OhJUA5MNcn2
jUSnjIOI0oV/CQDXvzgUstGokr03qVS9IA7fcViMWfhuiJEH/kANYn4bUoNOSSfn
6IruL8oyP9BYR5U24cj+DfmwhdfK66Py9MYSDGwtmJ9hsSPBfqlpknYCZtDQS5fx
yncRFfFLVm1FXtO4j2IHlJ4RIAY5TztP8fDBjuAgHjbdxJmjSwJmK51EyNeU3j54
PUqXDSwUdbiLVEQjX/8mmsMM9Y+iLiRBp8tUeyC6MgG6vYgt00uvVIhbEzE5Iawv
zXWWMS+tcW3h87drZfxw4VHw4Mr++789QQY0nSYRHpY3zh2A15T/UKL5KZ4ri2fF
hJCNdWMWgBMFonUxgxhfsuUuJ9nUDPq7GSiapFA+3uTGCeS4Ki+6mKUZvY5GkpqI
ICxWvRLZzUGKCHM+4Amj6CoL2oeuxfSTUppzoZKda8q3K9iy9LwBABZsvq8Ghc7i
7qDAku0+5AKMpZ54ujMU4VNzLLQRVUH6U5fdliYL+lFm2pfC2ov3Ar+BiXoBPh8G
SfZhj6ifq6g+vQxaEkX2MOPSeNyvn38n3F5zpHLm/yUBkQfPgzFhctHynhMEpa7F
jUToZv8Rm3a2M1nGuFyICCcZ9q8vTQAPFfjb0njPjC0FyoLxVPMOnE6goOm+uDy0
QlGlxrTOLWz31SWFBDa1QrcNeV4OKg1KwHgpaRnzWay4XRHggJMTcvFCefc0NaPI
pkfnQ7cSiOYgh3VDBENGIuLKyTjmC+Uw1LMhzPFGWxPenXdlJeCxW78B6Motkuhv
QR33phUvh9AygOpO0/iimK6Ue8uIK1r952X29Yt29fcdpEChzj/9NgoynFXSCaSk
lBoTug7K5YazeraSUxv+pyu1Fdv+S4thLvlCoAF5SMWsmf7pKcMxg5wLo7bkHFmS
GjcR2zrALnUweJI3o3mF/Wg0Y6081zFfNG8HDRi4FR/1C2A3lV5UzpWmHuodPu25
6oGwhwOMANx8ykLw2vJ3qo4aeXFoJlr/z9/3sbK+2rpOc368n8Siq3S+8Sixgt2W
5rNcqkrKsZmD9xGokYiVm2k+a0BQKJz+z/Rg/BeaSYbkmmAnqcE0CfiDhlhvLaLD
qSsONHI+Lga2WIOUD4ec3CLDkEn0gRJotVmoif/Xl6WtpZTtLlJkZ/1uVHmyXleK
tkBKfAWmxSm+VNksFSYJwUY6gmBsU3lmb2zji+q371hkkBiXJryFUypwDzvn9AjC
PkM8+eGH7hUCkCwTtzqEMW8RuPPTn98OV2+BSPE4ChQtRmI2AT4Z7nh3nmK0IfrQ
vWFuHYTDy1UHDyb9s/CCFJAAJ99leqKu/Y/cPup7o15tBFadL1s2HeU5luMTr5aF
qw4EK/4TBzalOXJ7xuRqBZGeiGe5JbbrfqIXzIc/Fsbn5osmru1MfLN6lsCTWK2k
M9Tc+0DqWw0xiiRIFkpK262m5+Vwx9e73QenQGHz1KDiJSa1lTlWGX6+/Kdkgcml
NavYlQFnSrqJVqjHRaRUJLa9iEqaFrIvYA3J74Y01JGwyAlJPtcj+9sfX+CctyBn
0T/fmpuAYPPVIWBneXm14wl+hnYf0DTJTP2D1UcrKdMJiyPvoPBXUqRZJn+Aujln
EU1VodDHHcZqkCW1Zerree1n/p5p1zcDCXVseEypwSAE/Cyl83UEriGcLKw2fueh
mEZQnrE241aU3ZoOmSc0JPXjg9oBlp1oRNWMkXExooGL6hKJkuluJ7e498rKlIXI
bO1giyWscFhzqhrqeVqqf2IG2F2bnp3n7fE24yfnK3ZrT3tQA2DYtzuf941CzViw
EywTHZNlC1ql+uAbXNwt5mLrkvm6IMrMUKplinvR0CeWQeOKeq6lUpInG9t4SqJI
HMBwmCtNva9/rrZoXyKbljilbk8c4Oo1z0KMlxBEVdXdBk0UvuxYvFHYKPEDLmeC
poOWD3vQeQ3mZHSnnIbqk/LNhAbsKENQtIVPPJjsgUEXMj0eK37wl94pJz+txR9k
+BZAO6QQ1lNcaYrHU2C4FC4qE4c4CIAeaW4daXB1S2BFmC67TyKMURCbX2UIwWhs
sHPfPtXX0vUtah4iawDPMjrcoJd+7oe3bRfxkK2foMZPbcjtCCb/yUwGAjWR9p2W
zx1QyoeT6vw2z6VFaxWhOck4yvax+4/cSu/jp5cpQJDOpUFDreOA1EBuyxi10ju8
ic1it6n7ahq6JvMrjtk2oVi6PHdVzlQg1jILMqNEKlQYxYH690wJFSIqqtUwqAFr
/tuKhVAvtOuVh439AbujuZhwydH3hSMg9/zis3pfLCUUHxEnczGWoZg7UPhxW4ex
AUezJ4Gqga/BJkPh2PehJU0sAex+hfx5UGcHQ+ItTEmmNTdJN+55BLW4FDhbDCAR
SxrLhhzGqKC/mvPrfKE8l7zK52CDCf4HeR4P5rf9C3q7S11bFMIGSFaQTuYSQKFV
Tr5nqp+hiLaLw8UoKsU2XGIPxyZxSYZwKtPQDfi2YcyEaUM2tV1s5pxgyUJPOyAl
hW+Y4dLsxG2IzsiIuZK9fWX41zcf3oITBqUSBWQRxv/AGKOI5StZIaeSz5Lw4br2
76AckwB5vffeD+FDlZ7QbS+bHowUQm7fqF0Xd0lcAyBcRrvN5Um44Whms7KpDTZc
Nb1H7Zxiqa9Q+TgJCi8iIqoMG1+TUEHwXdyAhpUgr3a+ow44YaLwJ9cnfa9i1DsK
pEfyBlN9yXW+I7fUUFK+BgTN614Sx/Hhpb3vyb9PfMPFncsWITHEuH7a9fHodFEy
ridkZqbGCdOkpc+Td3BB/9Z7ifIyyWp+u7hNKnlYbZrRa4onK79bkRNRttH0ixRU
lDcr8yx1Mpy7lnwgBz3X8JQAKXZqIaMAtbwhBNrNKw3+Er0Y8oYglb64+sHxQT7/
MgcxkdkTIDLKU0LL/w/ToGi0M+FzZK+1OcMNdi6eMuXVukGchmNKzdT8X/kE5x7+
AGmERvt4w3j1H7LcwrD2XpQexvgLbzn+Zm4L54xzzRliLunD5OuNVErurJX91W3a
qiCpZJe2CUP6tex8PF+22lqX1fozWJ/JivKRkzJD+csqS3aK2ZPsFfLPtf728FnX
TQJXmsuPOg68xw2Fod07BEZ/gLqlJ6x6atefrw0vUW35djZXkkvDpK1ka6XBBBim
ufaAlIOPYiUfM4JyDoIB19PVsVtiLqeacOU63H0BuYYnfs4kjpvmYtQMllexEwf5
m9UvoElx8o8bar1P3eVn+K1L5BNKDQweJusAh8ieUwzkQgXfGeXosRCmr9DSlbtm
MHW+csmAbTK7YCGNj3LKQM/lNwWC+C2YmpSPrNwvllnplhvWIApPHmtHI4HyPDUv
KgWszCJ33aU1BDVu/koHgZX7g0Lc0sbMkw/+6k5gVxFRWaY3PPa/3tjEKoHtFcjI
6fZx2V30QEnIYlz9hzEkTn6WARg1oKpwBImrQCFtleSzOmq882852rgYuFX1T7Wf
gqGRqZX3/4dFcup8TskDaw8v0BBIEJHPLOYMuG2FfBRDZEJRKvocnE3/trd6pyDT
PwmZQQCOZGVN8QGHvlp27Qbs+i+LWrnGe0cYDPVc3CO6bh8Q6ChJjz32BnReAj7N
A4KXPijEs6/LItMMYj1kXFVmuTFcrCq1dtAQAK0Jf+yK17dLYhMo8UjYUKi4CAc2
bpkAYjZac/d4A60kuPtlG5FzOw6iTzmocpZ3gkTr029vbLArNpeyVmGlHGrpYXLJ
VZ3nuSYKDy0v/SzmHAe/Szk0AkRwFwuu8Rdr1QQasa5kb1v9e9F+sTk+7OzRnZUR
dtMkMYT4sAVLYq69B2TGKMpdHJ1s+N+TrxwGVtfnQSqQjsuaNavF+msB5LUlp3/W
oTqHGlgaLtYb0Uru3i0EB/ESGUknG6y+FRpE1SE82iRVi0hCjr9y3sm/YCPByAI/
RgQulcYSGUSmPSu6fhIlVqg7J3QH1Vf/RiIsv24DQWpH1aM8D1wrANp9kgpYIBDV
AZNsVzkBfm76/bY3cvecvu2UMSZrHEhkPNWmhxxTRMe2o1DdcPeFiVL3ZrN49huD
aD9ihWVjCYiLXJs+Ih/ug47dy22vvymiejCkU2gK5m5XaNdJDLgmpLF9wzCSHqjC
0J+6B/QtRnlmmvMANdNy3yxyksvZj1hy/B755C0d0sh7a5JMiaIeYb12MQechs1D
QdPHCvU8GJl+4KeN+ymIezbEu5mP0PJMxe/qgezPTPt92c5zg3KJ/RqTo+hEnHc9
2KTAB/iHRrKnaa63e89cr7Cx76ksY5JxA56dbKf4XwbP3NfnfVSF3Vf/JXzDyrjA
AqW2XBpgpmYHAiPeMcF2r5sD4MUGZEFBRLFO62EXEv9A8n7JBFjN0YXcjliCPamj
YIAGrSQfZlaztQWxjZA9kk3BlCo3mTMzcPwhPDVoV99FJNiZD4cai216MJLyMXEo
u0hRlBDyQdjfaEV1l0aLJYAu+oQ8e5XapDwBgI7oIcV4kgCNsprjz/Vc9x4VQWRk
I64iq0EWyAt4jCulpca40IuNyHh4IwOzh/UIIrlycE/WHG47PR6CDqsNnn1O6oVu
YRUCkY8vDtT26yrkdVck/Zo30Ti+9vImmMRYrjO/0z1bSpQROwtQMrLvnuVXrak9
WiwjXhROZ1gEeQLrpCdnUhK7hB5hrj2I/dx/6NMbekSHiKi/rig/hzZ4V7ON83nt
BXQR8D0yJujrPxt2MZCwr7+EvftFgCYC3Omd5hiWPNcY9p6PJVIVOMXy48LDdl5C
qGLzB/CwAo09Cp+rtgowDtY0rvjbHlw8kgY+Zl4aMf31P5fjYEsBG75hbDxfRnBI
EDaZ+mVH1z1uR7or0wek5akl56sA4spjxDpsMvCLwXsxQZXQPpTUHIjWLHbfUL3l
bE2oFxy5s7OdovQL1FrknrH9UHoJU96U0SdZMi8pUtfpOjLSXV07gldr7HC1aAxo
St9ODdwOpvAzMxWr2EEuV6WV3TTTvAz7N3IEfrogHyow/CX0OQ2mGuusqh9f6h48
SmNNewe+GEG1JI3imYj1Ui53Q5JznF9Hy0vNZyfcmt3uGLdqsr72BuS88WN6cUeh
DRy7Uy8jLeARf/FNfjXtdTeeObU7gcK8gPflv2fS3H0pFiEm3RVSs9M99mDN5Xqt
STXeQyqXyZJceEbFJfsOeG+StrC0YXFZFN/ky6W+9lQaRGaF1dwNLPzwWUR5gnad
aj2NzveBEOtYICA6c5B0VA6fcQQ+AWt16QynSt/IrBXgyCtyDdNn5IvA0iT/Ytew
8948i/LMhBJmztnCOxxvC0BGFIeIp7VvmGySFmsylQ3zfYDkx6ge5a1xQSyQ34NW
XawME0n7a1dIBHahxvTS/ho978pea+lNhx5lci6y5SDFqrgHJcL7hXJHAfqQx2Pr
Rff3NrYuR7yF4gGYtqxbdrNPdsofhOz5hLgFViLhX95hkMBsgzLdoD3WXgOzv1jH
f8jcHegpQs55tb5K6lxu1Nv1Cb+4U7dB3xneJaH6KYNqxBPhx9eHUJSetr5Q3/to
jU6Z2vcc3nvw0YF2EhmjxA54QEpKp4EMJ0bkqREkNlK39aPzC9q1n+u88vL59lkT
xqv0cA8vefgVpkm/LCTekCwwHXgqqXbUpk8nLpvSBKBdwWSs7cGxxAICY+o7Ar+p
SehNyP5LMthM3SCkoUxX2F6lS1r6cGCqcYfwOHbmSZF7YKBpU1DRKdglJ/cZJqR5
Lf28r9FBrDmo6UawO2yIR6HmZNC1teHiKgho4kYqe/gSENKnP6Oer1ZWSmWxWsm8
k6c89HoNCqoq3QBB+M747V94+J1w9SpwxiqQeREyF/owESlp7gD2m/j/1g3FstGA
unXwJqle3R6ec4RN9waB7ox2/O9IcgburHQaW7ZsSuC4B+rhd57lSdpRp1I2OgJY
Wa+bh6S0pkk2c/+H2HJJzBnqD3X2+9mfOLwOSL2geVTXDy82ViYHPbSKDY5+3KX6
9EngDYm3LsSrv4iyG/C8FFOJWS6l2eKJy9+0xIuwZbQUojp1MdQPRclSVgrrKGb9
MN2H9pkiEyt7SLTqjteXfzKtjxrsmGw0ekugRr9x5xwgGL/KJdvcp948/4vhWXKR
JJzMBQgQNMBcTM+B/XEfBCB2Z+K9err/UOGmXMS/2abfsJOO2jgK+etdM2asGUAB
B9MJ3/H5qTR6SdW39LS5/7kbbcMGZnnSx0kGcXvxfdnsrm1nxIHdGJJzyQTgBHxg
mGAhkrYhCpZkvNKVww9zrgMoO8u/XaN07/u5bk+29SWmbj2sv2tpB162/ED0MEL+
0887vWg1ycRoLaHPSIw8t0FH8IUhuOduqFJZZmaCZJidisqL4rsagYfrXgjjYkf7
TddfCaoZHwnXnYvWmtMoOtQCNxywoIUXVxLtY7tCKLN2/GqydFi+Xp15Zva9AmA3
CxvtqaBlbfANiT+F077ljnqoJCJgPnloXBiv7qzPlOEmmneSQucqr2cJi4hnoIre
zVKASvI6+M9/YpISwFAANZTkiBMnR5xX56HhldIL56pYRhGI+BcICojara8SEyG4
SZ/qnct5B+hw/y5HMUnRAZg10rD6xIpy/sYuLM7oxFJ7p/chWB2LQmjyJvTFcqp+
WTrppjQJoVxAY6BLSvoa6/mN+wHkAPM1IXj3OChOkCwoiw9/ekZwSjmiz7RC1MgU
nv/BbrZNLRdesQ13wghnZ22SFh3R8MzZ0s9KrEtk2TRiQLGLAVIC32Hjf+hpuEKe
/tHsrhS8h/t6qwoP4AR4QQ7TNJ6UGKUkeGjNCJO9+5KBjjFsPlaB3HgRYA+41LSF
sjGZvaeYenlyp0Wyay8oVxmsik3HmdCLFY0pPaYD3LtGNO/IpI2GK2R7cznk8Oc1
5r2ccLDlvV5mod760JMZSDEB7R5kSwfOqc0x7IXiK3XOjow1h/Sct/nKC88HdxWX
vM17C/4i+AyAOc/g6yPtxaHK9EF+XwWn0SUN/lezgNVtKN6MZcYdrryKiK2uRHzS
Aaq3f1/X7qF43z7NEtV+nQ==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
P7geeci5s50VxcVi29ULLpX/tRJzLA2jVWUKimoCFhr6+Bftg3BZic0nZeTT9pbu
hPF2+ecy+uVWCdiM8PJyEM1NHWHJGqoBrhLnXgGsR5MDS8CcxjBsPiXonKQg8GGV
6uZWWJWJLi6reY+TCj4eAC5KzS6cSaxn3rnZEhh+DmpbPiQYvLwzccIIvJ5DELfa
d3b5mBmHmc5o5YFYBjcUkLMmgBa5KvxaOBbAouyYoIefeN+USNDdajggpQW3Q+2i
FHH0tnWidd5pjPqphRNjMeIVAEYBM+PLEEJdx1c385WIlGrYx5Y2xvi3ANqh7Txx
RTvZxuKghNFCrrQyUqMGFQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2016 )
`pragma protect data_block
/CA6HlvmmT6bJB+tZcOZkMshYbGu60+2i6jvA6IVtfQdDafZPLT3OOtf3KRBwMet
yqL4fJSfqPArXVNxeB3+o0us2hZIFktS/JBvZN3QwfcjCoaUD53jls9GhLS9WBMn
RhyMDTWstNTMhhovwTzRY9dhfnjHEchrsCAXJNTMY/nc1e3kTXh7z+8R4ic031gd
PqI0QKThlhh6NsJl44rVKq2yZnBN9Naq5Dk2SQbsw2Ll2Vj5E+XX3Osu16d+admt
YllgMM+gWO8M2GLX2bNLmsDtQ1fPgY0P2/mL0SDNzc3UAzhF2M516vSwLxF/NYy1
m34t5NArVb+ct4fexva4nxMhIi05IZiq1ta5d9absPcj6g/bD89IvgWX8YTayYE+
e+0kaSKHrC0TnF1bONjyEjNdra8UmvKjWhzaaP/u3D0Ym8yX2EOZR+w8Qm+zfhy8
e8iTLX9bykzuLJmn6nvR/pnCsIKgbBdO2wXQOscgZQF2SNv94nGKQgI6ZcjYA/6l
5vD6auYtmngBPDo40qfX5V2u13WofVgy8Rx2NivCYckn/LOKuOzOVFytKwJc9Ixi
9Bo2J6vfZ5a6Ph/MvTMiDAub2xCk7BnBubTEc71S89ff0oQ5h9RFKPnw4J41VYDw
EddWYnJDdttvwONaR/nnVECKkQuTpVEpSMY1DJ35n+32yzayFEFcFDbxgG3uQsSd
wGkAKc6kdVD1exmo8O0OtwDt/t0vsseswVJgFiondjr++BA8omtKUMeeUjSN0i5V
EqMJQ0uwWUJEyrrxDBM1uAKSocCWs6vuyW8Vg4pUDBVUnZpt0nQmPc3OQnI9qMHY
87QzxpylEEtjbZiESvv2JzEfjGuCJ6WL5fd6zLoncZoaFZllUvpfX2aor/CT9iOg
jIBUFk6885igqPfLbpOrR8W2erp+e/GdmhPmUNFLJHPCuqhgx1R0N5i+uvPSSV3t
pmlj05WLNATQxSobbOALw5XiNoFAwghv/XS71Q0Ro3IBbNf6gnz6IDGUPhpqYxZg
1/aH/Zm2WYOYI6dTGNIGBSOUFjM7veA0ILP5E4Mlhf9sagPoUmgLHiDSo3IkqTx7
INaEtnWod//52PFAyME2MgUijTMx2JeZ1IWiUtYEt9jrt/YZjMknueyFJh00ssQS
3RrpJOusD6n4c1q9nrsbsaB427A2Qn1yicgyQFeA2MaA65ylKYGOc0jaQzFguJau
9bHRLNi84r3i7w+HTfdBqRISYRzvmLMx/TKuWwG7VnKGZGrXpKL2UoD4YK/9Jwzv
/fGja3mE4D1MpgPqgBD1AloA2e5YxHDhGG5WLvjkVGzNRBIUXf9Yw2A7gUTnLJTi
QUeR+fm4CT2dLt6pjCg3yg5IWfrI97844xvddr2yeyulCrCkdyQoKH6EeyCFmDsh
SoH9tFiLPRkinCsOX+TiEbGEI4MYywNdn+g/K/hBFYQ7p1TH0Y+TYupu/6V5a0Fq
oBmQxsizGur+reqlu5d6Rs648yCfaytCkhIy3OfqLh4AgLR6JNCGbuAo4+OYcmf5
1WSnD78EQfeUjbK545KGwm612ugx3+9iJE4mepx6wtlvW2YuHtf78oFxN1CxYxyn
wSIwLQI1lnFsfNVaP+NusT3rY0T5ulG442Q5pxvxEV9wjMyOd3yEH0P7jUGBRv/1
o8V+bFtKD5ZD/Yts4z1/OrCJy6EDiTBQ8HG+fRBMLaWlpwdMU7h0W9iZfAZs46yH
nziqudL3IecLz87X6sZZJulzp79Q1Pi278+cPk4M3FykMCuwwea6KX2VtUMCEsP6
nXxE1t6plOw79aOvH0uooWjV8ytpb/je6AKbjcFO2LXEea2KqVomHEXEgLdxQ75j
W4xZ4qXtLlGjyG8dMXSF7aQZRmbEpLoJYUSXlIYl506BKNPCXZ9k5El+dZ7paWwJ
LYChiAv/QhtJ2QGnaXpFlqhz2KQL6ToRuPPjsWGnPcx8TSP4Ao2+onTNBrQDIUKb
x01kntYQLK5qtm4QzkvnoDwavPuaMjNkiZgTmJ0OX+lt8Lki3tz7bwE00s2qLKG3
Nct9YzfRGbT/oBL8ne9pPN5SgftYYUggSCdlI8wGQ45sYw6YXdASnh/+JKFUbmx0
RDLxfXU3Ml6Q6GThOwo29vkYUdDpQKsqzBof8RsjbAkzeaPHnMeMdIjccag8h0FX
g06p1+fk9HOGVoKOdEZxE1WiIJSolDIKrezZs5S5wdO4QvvTPdkhjFUBsuNRpd2F
iUPJxduOii0HY6RjHM9gG8xyZN5mL7JPQ/DHmjcVzApJtWhvAQQXe+SU9VI/eZG4
oKemL20LD3dvizVMbH2+rpc4dSJTs9JG6da2A4uE8BDbWudC1BGlsksuU1kNpvU3
/E6NX6mZ/9pNEMcrm+hSKJeiqFqujkr6vXTzSJD5qMrQ19TVhyJZNyr1m2Dc0XMX
2o3NWxux9NnG/OtT1+vU3BsUy6yL3kRCThHnmi509G/LlSgPR3oC+e1uK5PbVaPd
/7+6jF7SQrj+hBYmkWzTm4TQYcad+5fkbFHsOTkTG+DelHn0NJc5jd/fDSphXjLb
xFjnyDkI226naqmUMxnomxWb123TF+L9HqfeLv2ysihhwGuqSTvNU9EwIt9gKRUy
xpLDLhJ96PhwYvvIh3ZjUYtTMP8uYPiABe4FFQNVssssqoNJHF6PiV+h3SV9O3si
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
DqGrbyvn+RdFAQbmXR6UuSV4Rjsf6vyuekfmFCtlUUbe8VaGe14xJoipeQ1fNvFQ
ujCQxjxGGi2BYwswPPz+8M2mt+EM6iGOI4o7pKd7fYaOMxoX2O1mawMYLnW+UyFh
94Vyj1v0TIlQdsdnStQtaJ0LiVMIKHO0BpXjJkctllqu+Tyb7AP8B7OV1mUcypQ1
D7Eb4UmanSP5YZhzn2lc9EFSpSbUn6075g9bl5nO3iKhksBkRRXqx/WVVBzrlWM2
o7qjQqRtN5A7XTF9F0oEgC1hV+yvzgsKLVOWdecMfYLnLU611r0yDbTJXCSCQeOr
cZAOvXCPlckCom68fB6NcA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10976 )
`pragma protect data_block
w+gKnEftKMrcoRP6s6HT/P8rCvJBiFZdfFYPlqCyAV6L6KftMK6LBjk/vdnJ7kMb
XwiBICTVY1mAfKg1RFz2bx54T18FvoTQ4O5NrDWAnq97bYM68OWDMIurRSSm4koz
38xI7HgvcJkV0D15tEDMjL/MUncv7N64lsxE1/LXQxt9vkSUYbXPEfOVgxJtNdf/
kG5DHDCvFDOfyCuWVpcaB38DikTUBye2iVRUT92JTgJf6/u+T06qicu7m4YxG6RD
nZ5ViwKGqWjrHy5poqR3AXJT4JOaH6P0/K/poZLFuNoC/4DN5chff6yvU7t6jSan
sJHSX/jiCVe89kve5eT2p//6T1FgzGN247ClDj3RqZC0vVnsglhCtACTixsVkjS3
D5G7YkwwU7EZ+foeFfvXmvQowGuC8ei10XPVqD5nGBbVxfo5tKh8R+QKq6H7YH6Q
vLxPN0d78jpQzsgsJbrIPc99fuaoSDnmcrVSDj99zUHxgvioLDH9o3zDB08wHEDc
kbDpWEp2ibLZcuxCrbkvFqjanQM0xaiYgBg958xGocIaxTu/o0wSrqACc2WuKWDw
HG1Dyc3CTbKGXnjVblsMr8UFHagnxXItdBV9wRsu5lu4DzSFqWJKLOjzdDwc9VDI
Ysr3pX2S3Fzzpl4o064Gm4DgF0cyvCpoy+s4Aibcrwj5OUJ7akSmLUWOodLFN271
LN+m1M+wW4nXlUs7NAIL+l8iHBAgPV7oQw/6Tgsm7dZJlNwh1nPTJ1tIe6E5GfaT
aOZL/Muz2xiNb/KB90Y3qN52Mus+NduEa548Jej1nqMQAWwExjVxvjC2Q6/7h8lL
o0MBcQ0JmLChI/yCN3w5C8VRs/86IR+IQsYztPhtfcA23D4YX8KVhKoXN+oShgCN
yA8cIM91dbDrGr7mH1rsDbUpRphlfya3hupV/6+fSup+OiS8M35NeZDxVgskysYp
h2KznITTVEFe6HiDH2yaP7mdaOCPx8mbbC6hw9RAJ6W0pabyOpv/O3NLvZzeEgTR
t+Ht/8Wz3TzylAvUuYVDiO1Xjqg/FYS2CMFSFJKqYaMO+Gm12ma4qLjS51xYwuCl
7na7QPvryLFjHZIFJuf7a7brZ3rI0CzBNkARP87+VpJKxKhMDVM47JsV9sOajMup
MWJ8GlUcUBSnInnUwcxew6hnNvC/FcWRTjFugB8EtoqMMTl7nncnZoLM+7yvlEgr
/m+AyRW0VIoVJro6cHElMJp4kQqIyUTIE5YTvFy/qlK6XSJRhZUHHLtxcg+J0OzW
a9cOf/2DogAIgFsEwr7vHpmQJF+hwy0z1AMaLxJMSMowFXMMC9e5KzM/isW6Ogh0
Ix53PIl6lQJzmBKEmKwXPZIiZFej6jSq4FQxLxkPf1KCsGbYXrCXm4X2k1XCY3uF
IuXLs+YTqmvkLm/Y+TMDZ9OmfxydJ20HDF22cGIBzwdBe/GAiwKuRT+/Xy6OVPO5
niGNw8Aba21VrsH/ndLXsT/QY9FMtE5vrd+FUEHE66bgghuVzpDussJlL6L+i2sI
iM+OXFmfYHHjZT4p+tYzj3qWZfBdsU2mD6jcNlBS/in7sN7qqXbxTHecoOAZWuwY
fx4lxwhIZT5YsOQr9sqcQBmcVquF2hqO1LRm4kPQot0VIacCFhF4cO/DYtwGj+a3
+/9IQBE0fVPtMylzz71tDzUI4wuGXT6UGLUabj2GDJFKrV1lfBVrtLQ/4FNuYdJO
zn/FG6XfGo7mc4Z8U1u/ySkMgk8YfcIAQszC408SMWJlqcsL4G5hBMwiufQlb39m
8UKZUnbORQwCC1F9Vti1DxGFHIU90QKxVsBZ+FIcoEupe1QY3vMQWH/gV5dWc9Zq
OVEXboZ6d63x8ootflMHYiU0krbMQVq3jaJx0w+wIQMRxWMNcB5OA1/Yv9aYZ3Am
rXSUUQnolJyZf5evNcmSw17S6iRpkR1f6tX+37snO6VQPv+3AJcCCT7jysn4arhC
BJMtSwK4lqk4hlQ7YajhB2TQLeolfjOcWl0mnfFRBzanwwZ3tMAeKHfiSUiQBa9g
anOD9IWZYJlPaLNQWzsy2JylGw8yNym2NM3XoZ4w8YURKE/mXe4c1HtmIyLbGyXy
3bBmMV1sAKbk1cSyOo+o6PVhPpFSdkY4AtL/52YobRNkYy6zKYz0SYhmcjZaYuEK
1NBR1jI6/yBbiazEYBsPHoiCBIl24JeqIOOM2BNEfIbgwxkF40EeSfHRHgUXp7cu
DqfGJ1sVTGwt5KEwjBK31plvvpu5MGqe/TM++e8N0eFpLOL1nc8v0KHx/FP+ReQp
DZs4xMMBVdgwFG2Bfaog5SItpaiApBENKomPFiyCUJ7MmPjixwIk35EwL/p6L8K+
xnJkMDRUuIigzBN44WjmzAIxISA8RH3NDMoBI0akW526qbK9Q9bgv1DPNphbn0T4
OARYXanQ1iKcowRYq+nyg7PyMJ/kUsNJcJiWpAno2r/xTsuwc2CJvN+PIDXUqSKY
t65aJP6du2ahhSstIH8jCsc2BqCKP8nTo7ECj3L/gE7EvbQdpon7s+qPzsKexdW2
yHn6BOosyIutU8ZOxSdo32tRgQPlmmCIjfxEtacIHPlDlcmWVbBnBD76nkkZu+ot
xqaK0BFvoyObTZc3g7pHL13pCFrb4denUrJj21cXxBa4rg9Wle5C3lOPLJzGjsj2
0fiSZS7FgwUYrb/u9bDOlknArVeCHTPeTk99lNSWYQamRVw/NVflVzJ6uzCu0V0g
lSEOfOChZUibiuNN1k9D9EGdDR4Y1ZCIDV/njtncFkpkDXa1atvsMfKLlSabndqX
ZiQtBXkZTJ2k2LvSQBGYND48+b3JdbgGahDlLOXUNgASKQLQa8JOlx/jJH+EyTY5
QppqxbN873/X3xAhNruzJRJ8IEr3iSEaLGLxn6BSgV1VtunkI3pq2r7NtFYcJrAF
GkBvYD8Xc0omFccs9ajWBYCHifLCrR0eMCc8aRH/hAEp540QcqNooGjgTPvy2+HR
PSJX8MT7JaB9uf591AoqAqseRt+3yLbfGjbh7wo9zH8eyFXYgQooYQvOU06IMbx7
nFdkF+Fb8KZi4WT3ysMyn7jAY12alNWHXBIOveLQ+I9LAabgYIJK7dgJ5L07fHBY
4bVSFDkh3RESGcUm78SSTcb3xsF+p8Al2HXyx276gI+JnFZlapuE+rG8Ax9Izymk
ymUIvMtn0BTNcR2j6eSXVeFKnB8j7JR288xduErsTGfEPog9r9uiGyP6x5SCvut+
mugXGB9Ia8xvZ6R/OY7E+cl1JlmWQpWiTqCKi+FaZUG/9dUVIkooQYPaNlj+hdyX
TAHsR0i80nvMlP74dV5Xk/5BpwhffyuVXrJu8z9p6HuDwPqaRK1TZdyHW447tabL
dvKN4JkHT3+EV/1tH8K3C0mEc07GOUdwHTY6atNQEh70IJXW1BSTBJ0w3dFc2r+N
um5mi8bYDwSDGh8kx3l34Tmft/m9r1WmnxSHbJ6SMWqr2xPJuLQewinGMLM/ZgwO
0rNZ2kf51Qbxubf1MyXU9P/BcdEvw0AB5cFHCo0PKIs7lU1tlsAeTJIfBv1VcumB
p2FZ2IJIBwk2I/KxLZ/IdGgVSQVymH4EDTWuvFKMNhNxTZSceCVrz/b3gNuh2AR6
2BZdYIlEh7rBERfFK9H0nH4lLr7FKwFw3xJG+CT0tGcbuSOvIpuyPrPDGSnpgCAC
BuUTtIOmrNL/9ngatuEssU/Jh6iRfTZk3erebbktO/kHE7GcdJ0dKwGfWFG2fnXh
xisjmHUC77tVYphZzh4dKnwSwlvncz6T7JVjW+EghDOjwgxngg2ZKdZPgi//I/Zf
S6TeOKl+li4LpYnVQ/gO4i+ve3ujuhMlxsGBRfa1rPSFP1BeAfb5Yg66Izllzjos
ZkUzpN+HCAbJ3np4YFPWX1gOrhc6LFlMnm+g1Y4Ggb+Pauz21G60emVmgUEmBsCM
KYg3Crb4GdQx4YRiLYOyjxTkU/b+ZDAM6EjYsaxY5FJKXvOZDvLyHsU+2/mUGQQh
PgFTPmLJh9zvTmVvQ+TOcOW72c/K5rGIU7SzuIqyIr5dU5rHdZzp+EGiI4Un4Tns
hhgywTrdwbwK5ZQn8tPurerFOzGVTR9v4u/gKXQnzh+YbTmkPGEOBJdpUYLhEuyM
zbZxl8ffbOXhJMaZSDEBl1emJCScUqcaqRwz/JGNgWuHp+ZPg2/9ADC1ZusMU2bA
U5pckzOiGIePAMHY0qiipTXPiRtuoRjfRYakASf88wbveSwNkgbtaRFHKUL4LFmm
HUfXN6MCVj+WiVCMEGaUVZDuMxhZzL3TvWPZimaJMGv07yGwYlnAXqONANEVhU5t
smsUxxO3zfXRSjAtrpZt8K6yW4cWkbg4XyXtg6wsX/hEEZDwMb64zF/UDqsfPiQo
+ZFOlEWEwHDNoPABHESU4KSfcEijTWI77cd+rwlqaIh+m9H3hU3wjDdmMhVPr6lk
hHopum7TXqP/k2HaI2iS4zD0Qms7KOmaxLNVHM3mVXiWn0E1s+PFbs/TxV9eJGQ+
9+s9VIm8mOEOogixzMohD29UhaxnBWkTcHQhAz/lgkiumPY1Sqj79aJJbe3AODem
lKB+AX4VOVyGm0hf7ULafmQt+Um0AlATpmxRRykmFYo3/CoK0c4Oio71iKp+vVCN
Sw7m+S8iDPT6xiaQPkFsL42TfINvC73YvKhVASnfZs28QLVuNbZq7B1uvJxQGqiO
5sHI89R/ZLGlMKupQoZPxO1t7T7Ogt6Oa4a8GEa6yw59IGr1yXPsnv6WB5fj+9su
DeGVHuQg5lNGwODL5iJn95IuOd675EVfiaewFAWW3YgO11bV3ciFYH7oUGUrdNOi
IqXj1+SDdhGomP25KYXswa7MZ03a3Rq44KJlcEvAfmPfOF9ygtJeBcsq+a/GQCZ8
nRc6tboNXrrhsZU4xJgCfc2+P9tYTMeBoXopkmBxYidZ0xQn1rvlNCjbprNdpGoV
e8KEEKfpY6pDDqYvmimC9mrXe4Wm4+rCxCOv7KhmkaXzLFhjbPlnGKtqVUr+DUJM
KA/umC/fS6UjsIxMzxTma5GchmfR8LQaDRUNceLceKCgdvV15LBdkgLj5Rv3rajz
U9nRNNzbJ14IGJ3v+10idoWWvNXOkdJkCWrYv9vrcLFD2y7KB5+3LMRwIzMRA2iW
1tzqwsQFj/LHMWrWgV0rj/4KaRDQk6eeTUQ+ORGHcgnGzi3l/rNYNFnvGJzkrODP
CYy4mRNhYxH5jQzGqYgANAGXQl8co7XCpKmHpz89k0WmW3KGwuxI+gFztu2Yn3md
hrHNLDrf16I5qbnm4pK0rR0tMlgASX8/ItAWxKdzzWdqbz0o/6w7iRM3gDWWArnl
d0oDMHnGzSAuSQm/PrkPdvUDvezl7PcAZsc2P5YnBpGks4+2ZZoqOenK0ay10UKc
F7JnFvzHEgrhKaEG3aJ1KaXwPJAh0kzg+Bo68RTnKstjbpgvnqVt3qesjvMqKS0w
Fyu+UvMRxR1TVCdCGvGoeEvvjR1msfnrTVXwyXTh/oQOvLuHIbx/xIM5b0SHUuvC
bxU9hBBA27JrElWICZHnOS4AMUqqBdg+clvHQdnraXHVirowBI1+k+QML+t3yQoC
L99Hfk+wU3jLdojTnN5ZuPFcDItcodDi5QgMbh3B/bwYGiCFZufi8r2HNNGFKbJr
jLM2aR9xiBpkOYIUfUfNG0pyMlqev8z4l0gAd+opZ/eRWp4aq+9WNJZ5iWvHqQOP
DQI8ZVPUrfizxzRaR4ozPj2Bo8Gu69g/EPIbhKgEYAgx/+r/izIe/nHF3cTpeliT
dkCf9K8+gtsYtG22puD0MQJHAp+wRnUxWcF6pRfDRO7zP3CXH/a2odR+psmV4pss
N4NuxkSVaB/tWhJEPm80g/XMnYoWwO95hapq/JbkWKXt/xA6Iji3rtLmIo407mbH
edKDms2JLFERHXZpsMcWh+XMXH/BrUGHUhohkQGaUDhM1zPPxr6kvLTU9o65H9DZ
YdsE/vD+tXQ+8VLxXdXluzvi99hIdt6Fgsy/gbCA+Ekua8IdJ2vp2JoVdetIkznp
BXAqHywBkOtIZF1MeLPpmrxuFuQnC6+IYkmkxky3/O1AUvtCkXbH3xtteiDztJmS
lvQYAAzGyxrc3QNsZWQha66h4+s9bznCir4QIdwwkAcG3MF0WKiEYPBoH8PxxN64
nGpahsUySVySRMx4/UtYmVxQyODbzjeboHOee/BtQq+KT3wPBBUxfR3+YXxw/tOH
dZjMXu3YY+jQAKTo9EVXv2qQ/Hilj12X4FhYABKPoBdQBaGlJItJbbz09oHRZkzZ
SLohTaMouOdFF8C0kgDwkBqUV1BOcE7J1SwuA3Av2Ahn6MhFV9wHaix/hjTflVBc
wb2ENyfq5smkWgb0KYV4Av2Z9mtoHM7QBm/4ZBZKPaUbc/9vKaneq93d8wVLrK2Q
OhTSND/N4NaSMIfKxfMHLTMsVsPT2rsQEjLmsp+nTFHncQOzprBYTXjMboDMMDrB
dckse27IQwoyF2lzrKt7M/nC4ZtKooF8dciELnfeKs+2ii6KFmJSSbqqqaw6eoFa
hdCbIypi0Dd4wU+/ToblWz6Jxv443hNQ+Wgseam2C9oovBLKq1dMouYCPT6e4Hrz
gbxvSGUFwTwy2YQT0DwnbA4cJ1//aVM1viAELpJtPqwHwNTMdoXaKfAOwpvquCXP
O6WvAIvRGR4wnb3cgJmwx7KW9UvpFfZRH7IGTEOddlD1eXgg8zYqVKbWAUUjY4OS
WLuEtiuT+z+BwA6DtaLrjRdoKc4NlexMNqh2uLo0ii6IpqV5jLmyG/6b6qTUlLNx
fRP3Vn6PW7yi99QdOc1H3xH+YaKrnVH1aep/tUXzDz0nKSDPbAlt7PZRnGEJKDRe
sMu5gi6SRWXb+DDnGEdiRc4HB4Rn8/+f2kgpwVfaCa8HZvddvRs8PVS+vIzXfo8P
L1iyaUtwhbC0S/nbv8UXaJwx/A+qm2vjcU4sYuNujKTygBpDJLcKtFDtrRxUPzTV
Ft2Q5EravR4Ef2pCrDuA3RxFv4Dm7zcjc5WXb+96WcpOR1bo+gxXMewZ1VbTMnF+
AUc/hKSmQkWNV3O6qlECDB36eXZYCsz0MmVRbYt3kQ9fiLWMIbhDmgn7JzvxecJl
X4OEHw5PPEOl1LgwDzEFN/mEfyTu0Zsq844lDUdQGZ1OgV/jzWnONE/gBeMT6AA5
32qRaYSuWtrvH3h7ZJNpo/WBZZG0w8ayXo60MJEvYt5sXEKGY3CjWD4pAaOl8qun
/hZI+r0nRz2AF5q+NWwFprdxuH0EXHcqQ9yj7WKnTjfhx7GyjrkhhMANpJBSxsVy
OifJSoybiLbxPVeIz5wCq+McHYb8EKYEy+OEzb8B2egq44Z6dAwj+uLj5JzRQsTW
rSyfLrDyhMT388gYyXCIsvTt3PLp87YmhMbg+K32j8Fg8IQhBqP4/SuRfSUGXkPi
g4y15htP0Rsl1kxTB4XATQdmCWSJ4VN4fMuORGWLiA2PBHYW7UkwqHdWBfOYtGtJ
Mfufgj1H5fMB07jiewsEvNPnfd0TvodNssJdxSZ+68dy2T2xumeAst2EM0/1rcvg
LKgyjHm+Ek1DrAbyloaw8czLl8cOXk7el9CVVHy5DpnEonb/a2epoOl7DIDyAloa
HMYglwIjI5QG7b5i7Trn1V+Krg9iq+2gbbsXNiLf3/j2vwWwZBMI+wBftKjs23QS
McAYNWP/yEMxnBH6Y25faN2yAZco7pTOx4uDalqICBmRAfRpJ7DSHl8KVT8KXilr
b8kyBIbIlHw6Gb/ohPx0Vl40kbkU/SRYjx++kMudH6p/BA6iIN6X8p9/45DYJJdK
wQpE7g6YQDfC1twPTnM8asDRhDnFg7hyhkTeM7UjnT3qm6Im9CCvbJTPkNlXDqG9
cYFwFMOl09A5oWsHk6b8HPZUqeYt/+yv/zy2oPuvL+q/Z/zVB/UIPRfUa00nePSY
fOl2Bup7KXLYSr1f9T14QKS6I3gw5WtjGuJB2BPhXK3TpXXxMlsaCLQQyWnRqk/+
zV8wiOxFi+d/dwuNDpxhNEEn3F6oOmkdpBkPbOyMm2TW1RJq1R+c1gNEdDvl1d79
OpnvijA57uLeMQhSiWq7Cnh4l5JZNs3I86DKLCLtxnJwSylmFQY2nNE+Y9V0bJA1
DG7tk5H+n6qKVw83KWGSvjmWqkplDcahi7WKqnBkSA/7aKQfYX1/lRp1uhqG7XtI
m78oXo8bklVPVbMfXL078bknkCWC4hb685D4k2zIx+51Cd+Bb34lYD7WiJQvbeSq
MrbzTAynI37l0KK3D4w8jybQRZxkujtJDoLN2mRRmSgn+SpjJBswF67lgpZ59Hw5
gOQsSETXOVfBNu8sm3i0qBUpjPCYZN0DstEYW7jT1OgrD1Okeh1PLwSP8AA9apUg
AwvD1OimIjw57idnAxnFeXBtdp6VVzQnU9TmTYg9LNbUfTbbJmNyZvo4g8nZ7YD4
QxlDB147hZl4Tsl8Ji0xzSoqBZUfHqACqrG2tGNcD5uU0OdlAOpjsizjTqdDJShd
EwM3JenOqb96FIsBVGTLdAdtGxcjo9jtWlD9/hYilwppGI9P50TJEJrjwxWfteam
gVWtoE+NeXPREMWfiYBYkKcW/x/qcPT8GtNNjDpKKBjvDxUPiyQHiQH5ZDh7env9
yU6m4NX/dDKRKSbecLInLJ5S9XGN1Bbt8SVKRYuqjeexauIfo35jbckgaCTPlL/b
v50kLwjCk0bKMFDMa2x6CD7m3AkWRjiKRIzQHLVW411FLnyhq1HprgI1oq33g4JF
vOD4NN/1Gi0cVxYZf5l4+CcBL5qhuoUfscICt0gxK1TzBhvVmpfqdHz29Fa/lqXh
LnwfYrWJQ6ElLMTgAowIrB6Uj0JweQYjjYcWnKi8iT/eqijaJK/+EqeowBKVWeIJ
rFM3oyHICuXv3Cd5fVr0KFVkzK98fg35HFfk6jokR25TAmfzj0qLFm9oB29tk33M
pt8b4w6muAFqMFjs7zq9MJ1kospftf4L2VaF4OOTxP3W1T7Cx4yID64nZgkFLYBr
dStmIMoLMOaiM7KNWp79wK34AHri5E7qPdJCiF8bLih2CD4pny2cnTNKStAGlyKI
RWKXAKftCdSCIJY+7376IoSsNXmaSLoUggwWUpXLmVo4kC8BFv0cTHyA7mrXxYs7
+Md3V3x9WE9Hniwh4XyBKpyXmBtYvUcx5vnL7rpHPEUvEzqbZMMZil2C/JxF7Ieu
OGEaE9+webI9r25Pg2bcFS3NAlo4yvGoGHFpDfX82KZFVq7Ga4wOtab264KAWHBB
EAth5FkgMEajTGyCk4a44lZTEJM+wprvCFSBniAnoLtwQSdxWiRmqny504QyJuAs
xLmcL+LuZuOjKNyBRq0GtKln5v/urz/7CMrAxzdkl9KZiGrG/OoSgJ2gjUYPtoTp
/d2hEof0fZalSb4cv/GOElg/yKp0mws8tcG7WjxSLkkNu2tzb3h3V2/p8DU6ABf+
tO+PDX3v4tufrTQSzkporcgAg1GSxHgYXv3fP9djWXtHC6u8nZLANrsy+rmEPUla
2faeLv1YA0nbHbRn2NTo9OjNVg0XKrXjJXZwttiobqtT1JrcMZ9SomTA2EC/Fs4u
QpvdDUm9gZ9P/+xRCyTSJWLlD+22CNoBQTCG4XkREvJ+UKfGyFsCxDKxlSWhy76z
8vnusttRojZAThHPFKtkgZRf5O6sci1FUEuEcnPE/EuavPu3oNvNbMdEdCmQF5Cp
/ROkDPTtdYMpgaIhOkLpl8ZDOZ7YWhTBVu/6znbhgJnS4M6ltaRdGuAi0RreC819
6Sq+9C9R+GSKyH++VqM2u3phdNMESdzrBhb4StbrfESSkHf6rGmmd7pKasS/Bj1B
GMhvPxkiFE2gVVaV0F+BKzO3C0bCWLiFKdU+UWTubuwPJI5cKX3at0I8t0j8jdCO
DMIt8fSWjDfVzZrSyiHlkKRvox/nR727iJLGKbieUGiR7zyuC8fMKlLv8Gyloivo
k4yA5RcOPltVMiJB8OdZvdyPVAX51LtuCapzQ8pazikq/hIs0tgIFoVmsIDzCf9K
7fS0wIQwxkxxSpdHs6MRyaLRkyAyqJJvdoc13M8hsM4w5EnzRScG5a6dNqaPL4tu
9lL+CCcvvIuE4sNw1uTQ64yZDfZ6FzBDSyj3x7GW7r4uPpspZAyQWMYZvqmCfBtu
rIrOK0Uk8zK8yv6cr1IDoAVeN/f2y1tskNWBUaeeutHRcurj9CZDewp3a/MTi7za
/2yqkBvHgjkhs6GkIosgszsz+a+3fmTX+u/r2PMsR+EkH18tiXi6pdv71Jqys/WK
+iwPWL7dYU49sBvqR9agcAIW+t7lb7swte3jtDd+ZQEZUku3n9QXstjOITk8uUCl
+p5G2wvRksNsgW1ZX5UWyn5V1Fmy2DWo09klwmD/mZ6GRhbMMstTCnP7P0KkfJ3N
eOBLQjFl4U9mlXW+2hZfbDvHhR7BazafMdZyvPpJf6tHu2vea0gErBEGHm7G2RP3
2gKrd0PM6NUUgDh5EH0FXtNa0LyIJ7z6c9GBX2OX/9ffnJP5DzaVkkmsE+cTk5fv
HYM21MGY298wnFIWCM/eQ1dWEpfrDKfL4TQlXigN59Rq600vLQmh3+oxoFMJnkZN
I6S1LemaXYYe3gNyRqsKpfZKfsmUIO+wB6Uo5tGV49CY5PRMyYyjKs3oe5qB5L6k
7RlhJH5TapFkE8aHX8tI59Oaaeh0gGUwre+MUc7D4Us52IJs7IVlII7JHXOSBYgq
9RkkXFYBY+LKGLRn/ge3IBegDNk4+lHYlf7dyUTjnYKoRrMH3U+k/qpDSVBdD14l
Aurj0CuZdNy5CdWRHLq0JrnQ3M1Kj4dx5R6L1TCcKiJqa4HuXmK0Gpx52TRHunPm
ApbwNdkBGZWjp1okuQwM6TRoyY5pmmalkZ7zxrQm9LetXuZ8bq7qLrGniyP9HAlt
qOw0InyJUb41W2b1zn/xJiRz3qSYih0Tw3Wry2YfRWkmJUMjt008/Cx7C15Pmn8m
HM91sZxvN9EFk318GQP5+ZFy2XmLVDRh5l88oNjgshWo1YtmqIKT1ufxOihkK+Io
BKfjSoEjCjTZ1noFuLKgy6Oa8v1vVYsy5W41xPMHdBkJG8m/GKJ509ve76V0H536
2jOzxeyMHchOuRBz91KzZgyoFNXiHBwU7KIPMt3T//U395MHGjkObXDVHR1efKdc
ny3Uf9WWtLqfdW9k3E4JTxtwQkLEQrvg3EyPuSRCu9nH1kzviJzzDPO/21rWZ+Is
ktkIqPkdBGSpeMKe/Y4Cu1rGjjVmKINz22nXq4shy7KFsNZoe2znk0eDwJTwjHdI
rHkYhzW/YGA9tIJDV8VYuxmpGdMe/PZcDsQXp1BbaPjmtg5uR3O5ZQq3Yy23A8BK
b3Bp8z1HoSVKtAPRTqqomM2kPnLfMhRAA9MZPd3Si2U1qTIYWwdsFAMhDOt5nHif
0mPqduYtp6sM+wvocC6n5UsNT9dbckXVhei15yBpDSsmhEkJiTY4BrVcHN0ZUF6T
Vq0MipMUYScvXILyxOuNLWGsv+vocfThONbmsImrDNDUR3r6yp088zPCnZAbONU1
pxIYNzNM7lB/3p/AelAzcfq5JYyHzXlmZEiJ4uSkDzxJVwkEs+1iXtt8+8bFuBc4
o8RkmGTF4WrXqH/NVL2Wd68DmFTiwieC0QjNZt0NUvkPpPdRqh6Bz0SgFlX9BBYr
HDjJC5DkzcDFeM3d0dwgQXM2yFgszANv5jw+OCWh4+/Mg21/wTMshJymH96S2DRu
h6j2m4vbNWsyZi7DDQBcWhXRwNpKhERQzhCi5Q89BWnRQN+afYum0ew3NOTjDvVl
WNebkfy3uydcKbUnIFgGJyW64dTNC9DhFkspH+tBJHEHgOTnWPf4rERk2fTbdJAJ
N2AFgr212EYdl+46mAd1lE+YnUSHslGx6kFDKNezk/kpxLiqiL0idSA5TsKZqRTx
jYqnkKEjgeDseJ1geUkeql8SX4rJsLnYQAg2ni1Oh67VzYnjcrs2aVniX+hN6jLQ
y1e2FB81VvTj95y+JUYKkO0TFczwTz2BO8ItISKPY+q3VFlAAdnqxLwJF7TjVfz/
8CXiovzUkyyBwJInx4lIGNGelu0TAxUAn1ngcDnlbDR+QYSaRgV7+4/BXb6bTEAx
6ay8vIdcKpFpumqBW5MnWH3UKe6BkN2up/Xz9BzkeUmuK8b6TYYNTGRkkF+GE3gp
3YtvVUkbQ1hZx89osJqSAP6TtQulPsMKDn2lrZowhqplWabTv9gsSngX0pdiIPoX
Ti0/hr1Q/5WiOV6p2mtuGxe7mfyrWLTjDLjVHSxpL+nyug56OlWWTDXqyFFYk9lL
j92QNfAND8guMlqzYs7KN4GrXvDNX2Rn+1OZzlCLSEzuQmDtfnZ81M4JFdAYXuzW
kPJ3DWs4D/S9KlwkZhVsSTqHN9P+RrzIZM6qX4vK5CyrEHcO/zP25TI8a4PB1O8V
me1UzP8VI2SBpSbozpy2vX1QYxstH4Dic8y2jdf/YabXIzIHV+qS71OgOv47X9Jo
lgyjL0Rcnn3jMeAFs1r/23/rlCyDxuTx95JT6ipCuAGoDeNas/yLvDydK6sxRemI
1xmafJjN7GGy3ZwS908rxk5biYm05LnHCxwA0ssMBa0eM21ra+wh2YdD++P8x6O0
RO6tNk1g9t9gHy0UxqLa2Z62UT2dk95SSMoQz296X0MQCUJs1LX4AXh/3LtCGd1c
2rVdaEQ+V3jMcEK6oATbU1uCXSdE2VBllUy53yx2EosR+iOKGGtqGLdtFrOAFU9+
l6/YttNCbvyLH4deDtMP0IUCeprrMDqy2kKRRF3L4cCmHX+G8rZnHlKo9fvveO49
HdnCZMu/OMN+9wBjSqSNT56qYBjWgwdr+bAgU/MonsIgP8Ft7BMzNYkCPguUOJuF
hz0V0oADOmV2HWIK/0uTkxsbTxMV3mpzIJNVu2IG0zjNuD60STY59vTAW8OZ6AxO
+IvbFhturkT2mTUw7NX7JL1v/aS6vFpLwvPVqpYGywUYCGIrsaPU3Pi9+o24iRGd
d2ywsNlcNeQLAzsAZK+hRDiWd4wSYmZngjRrsPgOimN//KbXKIm5KU8r9ngnY146
k0IxyZ+iU4MMg6DGoOpGQM3T2lWKuxtUJhEyiT/SwCnzUgiqliHxwiXk6Kp+IkLF
+KnRT5tMvm2Ybm1lRIsr0oukr61soCax8ngN/yV52YpRdIOp5SCxNG+t3TG6HOo0
mUchUUoeY4IBXfYjlfcGzrQGBus5C9YczuYIROcKoAHbWUHJEx/GmDuaZneZlXt3
/KVHRE2vWT5e9jlRW6g+JjibHFk9AabOIRuMSZ2I/PoXJHYIw2JZhFVw6fx+ra+f
v+OJTy30oJxR+KXDItC+18sP5X80CbvVHaCjZlI/qQTP6aEN0y16O0rjZmjl8w/t
ygB5x1VL9UyB20b1XfCQUbCUuXeMis/5PJ5P2TftEexDXj3oeEJu2EfNaEf+64ga
Ivcu+jNKjqr95jsywbM8oEnKm114NM0YNspvRqBAujHORPKtCrZohq3k6AfX7Vaw
J5IJEoKAiVck9wtNeqiqQG/dTSaqdWE6d+QhS68RGLwNqe8BK/SUKIYUmUgk+qwG
3nH0JALbettm0QxzqXNiyH9jb3UyJsIX5Ia/i3HwrexDzUMKHpY/kJeo69sSfqrP
KLr20Fgtcy/srclwNz9DkCr2EuMQIvkvDmUIK31iq8VDdypifR1dNg4CZR2uYCeg
CXw2Z8XD1sbsMFR7bdOM6UHccPl1ePA9yhZ0rRvcL3sahajNi2HQaEr7ShLxCm1M
DtZP4qAhhZ0UnbkO87f5bi42bYEuRmcxKtAOzYunstdiK1LUUVxFftJK9zUDvO25
nBFTMPklWAfheH579weOboKXWUIWn9szi5qpduHepK/V8tTmAWzL/brMISrcb+Uc
0t+ENTpbNlcNX6F69raTpBvwo7FHqm+LEvastIEAT3QvpOfRwZNmulUDwCXV5/9D
17FIg8aWNsRiQLo+fCtGFnAggzTo+DKidUTORy5suBEXrMpfLzUV+e0TsE1qSvqY
MlG51Pr68wJD0cv/ZFosSF/mTBnOh1GUjnCsVtPSTBhSv+TTRTJqiJKv9sn5r9xH
NaO5UEBZoc0IEz5FTxh9EfXyJVO4Ea3usQ7eCRNsnO8byCsoF7TJtItu6VQaCL4E
8PlO3CHpNoXs8jdcWox/l99kVixdyp2liBJYN7/NonmVrleRejvGH9VirUKDxI8p
sOjRnAilVGTvhnQPRmyTou3PuQrMD2oCO8natVKvGhyTKS15oxcIxtvbTfcj8RYD
YBLl/K/YfYIt5rRCRb80jqA94laElT+454QE4alW83z6iCfoEiquvFwNm7wJK7Kr
yMhMJDaCkCyKr/JIOn71ht7UvKtgDwwvCgU3dEoCib3f/+XTC81kTyNCmPHWJ0kX
PY+KteL4PH2s9DL6CUnNLmvQofd6kuFGOW2Gymv8Qq6pVuKgPlC4ddb2R4ab0RAj
IZaXNao5NSATyxiUfMq/i2jLYxfG3qGGCNFqW1JIGr8=
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
PFMRH5xeRmPnKtBZK2UnScsJp27+dgsWUC36n7O6qk2X10txWJfvLNOOenGRQntf
fy1rEa9OAiZPFfApIb9m947nLlXG/oJioDP1FYLb1mO9+jV/rqgwbL5LNxAv9z9P
DFRtQ9C51y0vfKjD6PwySJfB0ibGR5s4qqOzgcOP5ngV5HTnEX0RsgWAqf9QqpIc
AKwKYlayM7NuS1HtS0kZ737cC8+GBqgARRioiYSaz8kEk9LXcBEp9fNENMGxnnY8
eiLWaBz3OJc/ZiiR1olX2+dI6eILG3nl1kdzh2Za//0v6KAchFqwO7hWAetvUkza
tPTWx+wazn+s8CoLtItZRg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5040 )
`pragma protect data_block
u8Sj5/b1jKALvlRTRTzrgp/K2JR1Bw4eNlGkg37Rf9+XIkcaZQs2Z5JO0aywpp7y
ZTRI3QcOvFRsK+LIdIIqrAgI28FLkCBjuIUTr4yNCHcbSvKw36Q1HgcopGXzAExe
4dsa7JP5D25d3XnOo9qxbPQxrbqWvyRNygkKWBYo++dxOD8SZgQQTEpZDiXkmhTv
ZPlNWdindh1Xixugx6laWXKO4oyaNSIAJ1V6vXy61UOjiuas4LwDRMzbjpfHrguC
zE+KNmoVdIdC9tEL1ZHmjJFP1msurHW1jNgZnUawlrX16vCwGuwKm2CfSGLEvRxX
qjPitTccs3uA9XrAMkoKdhGkya13sIG9qEpt/NALmAJ12yKAMSSUOp1zPKxkZR34
o8v4O8twwRufzgNmTD8M9gSJA/Ov0rpRuMKcSZOo2SL6vfMN7pPhnYoJb8Tg1zqI
NIDm94kFII+6+1KBp9KP1SqAM0eH4t3e8tDd3rNaAQZUE17OI0t6LScQ3k5WE80c
HFkDhFWl5D4wf2mBaQvvs2AOn4FqvwxgwAF/mAvGjUjJ6+CTIUn8cKmq0nyJ+3OK
Mr0oYElQerYSwm7ZmWdk7tnolbvYcCzumreDxDMa3FGl/wpH4oGSBkw/MoLed4OT
N/TbiPsXtdS/8YeBxdvvCZiN+tBCXJPmY5D5XJOpF6iNj2lz7bcvnaD638R+bi/Q
mpcds88n+lmnjtIokYUl+CCE47n3KSmQ24UamYL+uAf6tDB+fqUScshm0P21wgHw
2TRIWSYYE/lz3l1gCCkyhHtZbwK5eb+iI1gIwzcdoCRx7Z1OqfBaPpCEahwtWS3t
v++hvYd7vxRs3B6XW9DRssAFjST9Ve1dWfRWtpd1jk1iPWSdFdeysrNyv/fB8cNb
+9FgMg5cycnujGrHu0xRBMrISdIqPLb/g1ttfbE6XvYxBvrm0+b2qWkJkA3DzRHc
d7U42TOt3zeZ8JppIfsdXYmHINoaYN52gJoiIfR8n7B+RON9wEswxi/c0diYFI6K
4QZoa70zxSIWruAi0wwciqugGBYH4kjmgrkE1yXI69tyIf/59yZx4xhA8r1UMeT5
SQSctvv60gn96sBqojS26YMb9a3hwOytZeAW3NNdRd66MndiEO4CB2bz2qJoOofh
F9Kakl9CX32zkLj+myTcBB5+3OHQLPi39jjLxaynue4gtvIGUpUOIfDYZ43payNk
dA4hRxXUiVcH+1OKEnWVRNOd9k0B48xHihrwpwpB17V4j8zB4kxcjaT2YKPxzHoV
A6GxcZsQuWy448qVhldcJq/8ENv0hQpvC+wnOmnHtk8r1Qhu5jUjI6jPc9jZAe7M
gjVC764zDB7ZzEm3V1nrRZy0pRWvI62M5JlIkOeAzVpbtvGJMdZ6afV9IW/oI/nT
JHZkfp0PcMeYkobCNghaYgl7I9oEcuMmPoRPoKMZBG1JDvSeaA0sQJyrFB/BW2jn
/uKQjaMYjKw+InVJALai653y2HoHMBX5/wg74bZJK4acVec5P5Nt/wvV6speP7MI
q+utIRNWnO9WtUkObpRenGsKwhFE73G63MKeYZ5GFf0Pi/wVBlVUORORHyjphBLV
jwny8bXues7OEsBWzfkklgi3kGD6jo3rTbGrEOOgBvsvumTCzjbnhIHj2h8wdBH+
7Ct29mNpXzF2i2EzJoA+VYoP4zVnRwBYz69v1ggFPzkYhRLV0/OLGm7ScTwVjWIX
rEOvSbpHQnklG+rX8iSx0giGH7Q7BMwGuvgxY2rB2jJdPXZHC1752fhXRJdiUVLN
ZbjtlFVxb8ot4SkFIfHYEWmBWrlwtvsdkVzYNi5igynsPmw92H/4kyhjU7q+RIJk
YNeNgTyqCCGrfxbQROyM3jQdKde72fUZpKZowtGPTgTDBNeSNBTpZLDwvh1LjP0O
EWYPXFMhN6CvVA9qO6wElQLaJyUKR1N4oeIpAlHvCD1+h8Lkp86ns5lDvj3OvwYw
ZCuU0WnNTinXJa2j2ZQ42LefQDMxgQrQgpFQE6R6NWLiemtmS0DOyw2pyLg2OA7K
xmWfaOZYfDgewGsKcYFUQH7Zl3dH+VDEol5nMNJeJhTydJnFvbkBA43n+zYwgIdz
0bVfrLdkH5VibNeHkFBGwMgzMdy8xBy1/FJ1/kbKkxg/4D0nTEC1HiOI06qT9vgH
a/L6sdTI8COl5voI9riG2q2CeQM33R6LIEPbkZN0aooz1UwMsuWRmTikv9lCvRLk
q2jftfv3l7POvfvCLGkfkNDpEHpMlNkIhVO+9ZEsOXDlEQ8sPWEjKYNEgmosNf2u
EKYJHAO/EY4Xe0NGpxZdF4kWVKr1Uo/2IjQhtGfag9wKEUha1zWX4FNJhqpRIgQE
PXRlorvHFMJ4/1IK9AKFxHgkiAxVJGhJVg8slfdyw4a8lUJsFZy6OLlmStrTs57W
l+Z/cfokMpfB5s8CctI5AE7oZESDaFZ9mR8HsMnge+RM9tuJx6C+jq8VQJDFmzYw
NZw7H67GxXjU2/cjWxreO5BqNWI4sGkTUz6dmAj4EIlRvJB8Z2k9q0xu7AMkNevI
QKitaOvc6j2YgZRYa2ptEwJLOWVJyv/ERasgA1XhFSwIPgPrrviFF4qUjaJSeFJV
V+jM6CUGMUl4FT1+c7lGL5mxUt06u372787zAx7j0nhjENvb4sN/2ak/YQSeQA2v
qGlh9yBH1RnjhBxl9DYMJlxZEo4SImlQqP9NpwlSTF2x3/zam5QaFP9Sh7EONqJL
+v0da/iI4fiWfBm6WVLRauSGmfK/w3X6FJ8iO/Cv/savDvn4FkB5RiwJga+PAAOy
HQJWCb8r5evTZc7GRXFLLaMbiNWYi5JfEo5cZW/NteJqBeim6r1+xu9PXJ+UyDZu
NZetzMwx6CrVq7ZwOkqKzxoZ9Qle05VX1EO87CCHqNgdy6Y7dGaelwnVaaNICxWg
jYcrhkQHj9f6cju3RxJpUjvuV2f2VEejsjxWuB06qrfRRKdw7OYWFW7gmTKEHaPW
+SOIuUZzuAWY2KRlakhqq2N156PrekVuBDlF4KF48upJhLZtYqpGQoUiOkxmfVw4
G4gNFYG8dBsVo6EFqY7awls2FCYPlQl+3ofkrTbVTVEfDWFc/YVvpH58qtLxjTC2
4eTMxGz2/RTx1f1h92R1nkTlzvPbtzNhi9mHOR9zE79Q0wSR0UCzEE1E9xyp1sy7
oI4z2tFlEQEfYR2qTw74UAs/S9kc7sP4THG81LIJQc/1iK4TMVquJOu7vVmT+LkE
i2kYEqc43KV1H9sc2IiWOBMyFpl18Ypq3KPy1fvw3GjqCrKaEaT5fvSnBxypnHhj
MrKHxc0LqlYpiWiDBaQw+3296B/Z/UJ6X4VKxbK6ju9o9ms57ktMcQQU8qq8OkTE
9Vn0Gb4yUsoBlS1iRF/L1IGCxPF4DK04BXC2daY7uHYHvBpPcAoXU5tX+v92nJsF
fxD8Sr38US0dV8s12IAHQB6lTumRmgzbhaP/FN6C8XQxdf4ei38jchEyXCLOFheG
dBI18TLl9BaXhPqWV9Jcfn6YkFy9xXj6sbGtvcNXkvSnUaeVuZJDznTpZs5SEWlU
wg5XwjLSs9zrpeq0lLlBil3db7RtJj2ZoCDqrkpoid9MXC5sSz1u6uFbVIwVO+Eb
Yiw8Taub8167cr7kf8MmocAJsB9q/kOWUSi6gQAXytfG3pRbKjG3dULse3pDn/75
qCfUZ4ZUlqfbAUTjjNkTsqMx4PPv1JE48LSJJh2igL4LX2aajg5eNZksdkVt/pSu
A/cy4xYWQnfwMhPQCmNNMarncQhshzna72fGPTDAHnJeFOkqIuC0SGCe/0VUM79e
3ln4E+laeA8Z+XHLxswL5LvoYtRBcJh4ne/GZGfCo6AOVO1r/IKUc+AxAZeGES2i
+BdjMLjROpO1yeBka/FVJ3Q7AWpgvfoT+VMp9HBETcM+gcFbeC+nc1uZ3SBuMePd
cQ6ULQ4IZExABnX58CLsM/E8UHiuv7ITByPekWrAsTBWt/pvEQwkeskDzYc9pGu6
NmFvYMB8bomg94QnoFDpw8HiOByqMl9v6Mi6vYrPC41VamBzAwf8ZlQYI/BHZy7k
7mF6pOuvupF0OVjDvSRKhsBsAKjVjdTTCNgDVaVDKT551k3nGPazJCDxug/P7Z2m
iOTpjOy0sLk91ARMSbiFFTJmdt4Kg8iDVcGSVXw/Eup6Lg7zDE+wFEEmBN3NsjV5
RoXhlo9QhJek1hqqp7k40YdE88LjCxKA1ub+ZXRnKYSZKWqxDcw8FLPY7dkVKHrM
HBG0OHBVEuZMLfHRc+1LZReUb85LHAG0yrqvjMc5t7+NyStU6VZwBHtAx98YGSxz
GS0l//Ay2HgPWAe5DQVjMyysWDEBcYPUJSKogA4Pu9bTzEYkAhPzZilzo30uJsrU
TrSDT0LsArNiFfAGgmomlNPm+mDrtuoNj9c1r4jWwl3On/x89K1JCsCPaObFspG5
Jo616cMjBhhJeVlxju4cmDo1QWZtnytTnUOQNJ7cFJTN94/kGebJEoROCPyzHpfh
4cYhKEawnFtnXdm+L/YM8VBrpJ5o0waTwS41YRaaoLJr7ZD92ICUEqPuGUdQEXBw
/d7Q+/bgesnosC46qn5Z7IHrhagX1eY20UB/XXKOFhu62eSvXouHLoBahfJ+4PHP
M8xEvuohTlbKHQe2bM613HcTxfooTpC0JC20zLNwFOJdX80IszQst2iNhgGMbXSN
EzSyycLumhQ86NwtCpOI0jAUv77M33yTyf9/m0q4BA5IwsBRaNz0xI8F7JKd9KCD
GF/m/tdUXvKLnYyy8q61dpWbyxbVByKhHHaC2D2gxskEuixG27SF5Lxo7IQL9+db
Olbufd43FOUOlzBKGoEMFoQrHMl5e4YAaNj0jd022VPBMQ1es/sYMOiIj5nLCY03
uVcR/LdHmkSH5E6dym697ZTaRd876TBX5Uk+2AONkeMY05P2jssNE2FpJzoScwJ3
8pPoKyu1ZvzU/g7uAI5J8YYuv6pRSTpufoSgyWeqFYRd/HYG9VMPSik1mtPaBFfQ
bSd3xMY4g2Z+2vGLn5i6ahOgXtAq5l/IafSLkpI+gs5Iy+uad7cUhtAV3ugR6CoY
AMIUm3Mu74G/S8rh6kdWG+maGZOOO1EiP+8Fdwz978FM1vdkflFzxTfL196p9L1B
MSv9GlSficZif7NQxLInhZgz/qzsWC+4auI9eSPLFSBkgbQnKVTSD7yDEhX8wtzS
LtPKjH+XSVMid7J6th7RS+j3PBTz3joxA3Ub5C4XAW6UqW1s39GMacU8rSnJJ8kr
cWUNkFmSAwE3dGSPUq+4t5+CjkeXDRLnle2KIs7wGdiCRhYaEtlewpCrgYpjd5B4
uMTnmSDZh8Vys++oWhzWlA3msaKdsBGeIlVINnN5IeJtW1v+8F53dw8mabZYfufX
b+ZdihJAWljilPiDqK3W0jqx1EkuiyxELT0AXt/T6ruLHbLbcADiNorZWb2hMR28
iB+SIkcffqdqOf9EMPvYYdzdCFp6znzmcxgLue3epE1iefvKaKYb5l1FRrRUgZVy
p3KzqHPdRHoqzf+J8V+bsWeed+1RwGsnsCDuitiDmQIje/9dDfMs50Hxpo4DiORJ
Dw4ORd34yJ2+fhjIUz9vG5sCEB+8Oh5IkfTULm7tyzhlQrfJG+gFGlyROYz7H+Rl
Po7OYoZ5VytgvA40132vTOwLdyR+Ewe0r1HfeZ5SuZhVTMdpp0/cpjKzDYHhtXWA
A3e0mzm6imSFmpKHBHK/o0zdcNq2OcErBnyu0i7a4pntsbPqESdIGWM+lob2Z6mf
O7Vf/vTZrVjDNXgBSICtQie6y/ad/yGCC7o076DboVDO5pGL5sCEUqFOVmKBWVKu
ikypN6VKvNZxQJYqwAuWIdIGjco1VSMh6ZjtWcgC4ZIpm3yaR1PKL3iUatCD+Pgt
sOWdx7OAexP92ab4Lufssv4Ypo8yYVzwPJoHx8g2v7PGSnypeNHqvZVqEUdT7ja7
Fr+9+gKU349umo6YpE+tiFx+2wOk4J6Qz/919kjdSQcFzvZOrGCejU+ALa6T65SH
rEgh8GkatABBJmiYEI8sAtXBqPg6MRVTagA67+yysl2qyeLdvUXXBVEIl/EcEJCo
90O9B4v2vjdF+ci5FbQ4kIBPdXyt4lqAIJBLrLGAEVXoVxtIBkT+gWblXajHTPwV
NO3LxcsbtHurC1w1hnQNx/+zjVgc109B+Cxrhr9rJ7GcgWWQsBhaqPMtaEUIZjng
hf2RT2yz1umrgZwnA3NnDsQN/tuWi5t3w7X90M6w/Y8RntReMLrCHZEyZFiYj6rQ
igbNqZJbIJ0eSavisHFXr78nAnUc31Y+EgHyNF7Qx04UDtGjnNxot/fE0N4T4EUz
2dbOdetmZF3Npxhv+WptjHhOcRJys7qPnfib2sefiR3QhKXSYbpR2n54KMyXOi93
ZVNYP81zanQvG8/YKhW9JzcicTQFHJ01FT3SVrfTABUd2CtL9jVfvwoClRMOvkJc
XKd4bX+eWSISGwORlV5Ynie99fr4y/wXgRnwjaTj3bxl+cbp+gzhlBXzmQOE6uXb
l7bGkq00LXRa0sVcNWFJTmOe01mYIFXjH1vqfGtnLJJojbMK55bd8oK71Zu9D7qf
5p20zRkPSIFwdhUoijv0DPntG5dlxm0xZQ2yX3oVCk4vtx3sgqS50xmpEpsog2PY
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jXfSq1ZXPxDmCThaEl4tNdKE5bLOwsWTaej6LeZWlGgBOf1fVmLLTPccZqEkHhE8
eP6Ocmalzuw2puso6hhEvw4VZxofOoYOvsaWe1iQYS5+FrX+0b+WHcMx3VygBFbG
zC9sL3kCN831a5Cj7VmtdOjjJBcan+hArOW0L8XnlB+tvE80k4++IhJAlIQUEfgo
sJwu96Q1n3nXBIcqQqgEATuA4IIdMkBX2hesnSuIiWi+rKN+KZoM5OuhtZ+kr6qY
5eUmXg5bn16hxPU1AZHNet03zhuZeA0ecI6kj/IPNaqSuM+/h1KNtXIvcKwroJtS
6Wf1IVKjsg9e7a078eGmVg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
3/mslXMwx3dgs1To+2QexY4CYcxOG5ukMzkOdjzJcklI0k+sLUnHDN5MJYhimNDn
ShLC4xJzJjb1oYbqMCvdx7Dkv8xRTBEFZ29eLADZi5NVrR2W5R15KlXAB1MM6DUI
uDX3s5zfaxRdmknl4d66cDrKKf0nlBy9Q3+sWALPTLOympPfCvtzEuf3DpP2IRY3
m1Ku7wb0X0yFHJMDIcegkJXY7Qcw4qXvwtC0b+iIfzM1ZTgz3SI+OFezekKq+hIq
VGeGXmjt19NwkgxrBAxtUoh9HoEDdJWSGKP16Y5T7jzxP9KcdJSCVg0VqAcAj9mn
gwQLgVzNvQg2SXWbAmKdM7ci3hvEZUkDNmtqBsqCzlRsTQg8at4cE7r94HgTy7Oz
M50zouYN+1JKJE336tWWGk/fCInL2V6K4pTFNTz6gx4NU1FDHeI4cqQQqm031EOb
0OEMhkOcu0bGzy2UGuMEsMT1UkMJKVSWscedNpFDMH/UiSMyNIzdYHNIKnQwMcVP
oo+GEa3n88VUnlxBF/i/PMSCYy1Qec47KVQXQFPuyclvTRaHgTbAw6mscH0+XUFc
R12b457DNrCrtpcjyRni3nR2knXQfXBNBm0xx9YQfkBYNSeqsAJtKgwG+xmL3k3P
mou8t5a8fpTFkOH8Pcz+9YtEgvE4VVdK+qEmAGb/S1dW+pEW5PRXxinEog1bgqGh
Tlpxww059FS+PPWeAlVzEqpGLPWouOSF9+XPeIVj/tsVpOsV2p9UdcuScgSumJ6B
dkbflqXuJgS3pv49yX7bVaRPRkGqfD/eJnUlLGKoaY+IRfN0DzK2pJNLD+xiJBNN
IBwAurYnLHeN0nEj5lU+j8tsmCPREhY0QHUzzU3mFW+SkvQTLBnwKVZjh3weg1HA
fkairiQour4oktMD6/V6i4cue3vmZOyK7Ny8YiWZx+4=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ZK3etp2+HrNQ0xHNxFpS5jNuAl6UWFF4T1eTiNGFB8ev27JkkbXnc9D+VOWAKc04
TpRx83Ti63DUwgAdbNOJhDltF8oI/+kw27dBwKOGL4ycoALOtnYCFERIPLpDQ94f
PA444zeIbk6mgp05IgtK7DOfioaQLgh/t1DRps1/HPrQ1l/GHTowttEhCRsStp7N
k9BD+QHk+UWvoJbtF+StX16nRDHET47CTehVl0BEUT1yZ3ORA5ubc/68fEW1QWEM
NyYHTiRBSRiWzHoyrs/jXgwzFB0OrrnVj939nyCNXU7mMglKHnwe9ao1izpsQSEF
y6UQiHhg7gLM+0j3Rd6edA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1792 )
`pragma protect data_block
qsGlUVacXT+fpGgFs00n9mQAXgfhoJVR2W0stXyGHLq2sCm6ddUkyNNcenQqwUkH
p0prOy1q8wqikYyHS5gKNTtTtnpZNp5cLYfEBBMOfqinrWWNGLMuNHMWNHbduoGt
E12p/1+UQ2pqd2ya9PHH87oNEXTNDNcnMLWLK++EEyZ9P39VxpyMYdmRodZJIeHU
y+hAWJejbwxqh+bXnXETwtUs/zX+JbpgqK8C7nKW5hDMp5ok+k2+jA8+s52/XBFW
vKMHn2qy/3Bh7YaZuj7bpoXt1KQ/5ICvjRvT5DSgdSvcMy0s6r5+kc2j1wba3fZP
hbSqcxnq/zc8WyJPhjecqLVyFpMN0djbkcUvodZhYcRP4K81U9MqhLtB15DciRef
ht04aySzX93Vr5PRKM80XJG3oWQQuTQLR1XvcyOlnkeC3elEOa4Bk6L5p4J/IcqH
zA11oHB366fDSLhyaq5bYoVChcgjMEaQhKRRKjB3y6butappqa1ZvLzbZ469+5R3
mE1ruFIdOOWRxhi922AZZ3S7DuFVk9OYW77zrZPc4bMz76ONCkpJHutGTo0xXaD3
1JEWFDsAlV5P3q6wj4ErNTmiRvMvRKbQEgwJ14Gg0MJ+A2MLMGpbW6quzzqa3p9p
ijD2aaMgyAspaGkhUI4E1vyIw7C2fgGQWreFcXtmaQzd3+TgkTqrl2pKIfRtCVRG
hlRu2RaZ4eXut7SBTCeDfqOGHIY8eZmkokJNrhCEcd/FlHsJ5116CLTSpkvG1Sfe
Yku93I65TOns9OofhwmxdUKa+aEs2RHaTVmL8vHVnivtwzaw6r172LWX4HoBC+0b
4lFZUWxySUOw3Qri/Heuu6B1F4x1Hc5TEx9ye7WZoZ+tRxLmnL6LYLBERn4SLWY+
AUO3+Km6dY1p/Z1IeXCSlOX0e4diBupyX6sfLTnRJjnaRT38lLMClTpco9EaEg7X
xquRL1aX23kiVpGpEBDTbX7EAfk53H+osyHFYx7+XwUnNbON7sQIN/My0iBvuEXs
YH1mnu6vkq588iBSMIkDfF1qNGQpZo8KE9gKTEJDPXFNgMGzkdTrGWvWv1nr8zx0
ngPZzYrQD28rS/Gaz6bBSk0XP4W75l0cYXV5xgjybVn86JZhC7nem5OULySR80mJ
gqwcpZJpZ8wsu3L/bA3+vCVfAQbl76jw9wNVHMPovtaF+i6dbmmsKyu1KOERDWnR
17MaCYo5LK7b/7+8mhFbv+CgFzClLJcOmXlQDM8xxeI86nMmke/03U242VSLPFNQ
i7dYxsmvg3vUQDUJiz0XCIwRcUuVLacynjUppcyqj1j+Ab/PRcVpybMDhHDRXO0S
BIx+0BA6r1v90ExflrIxXvCdC4i84io2uA5dmjEAg3LHvNOrKBBTn25gkYT5YS2h
O7jIQXq7VySV35/jlDhYLGsdrD2B+xtKgMCp/63Fy0e5z/+k5wQhSTwSGqmgmDJT
OLmDeiJaBeu4+XkV7jTphuvVyOB6h3OYhUO13MOYIVsEonCWKr1Ed3YGxhSmpKPa
OckaSbdeE1I+/6hKru5KVdCz9SkmQSrYml2nM5KTDRvpNl4bHN/uAUbwbaPaoKI2
1UERU9R6TBUKACko4tAZjIiak2ctxvSqDOIZJp9+fjhaClmFgU+hYjCAWrpzZMmn
ZSHPUOJ++G+BmXnn5zwO8uPioz5n6zs42jMwRGn2vOAxMxFJaEDd43UsQseBN+ZE
9f41T/1+JYlNsPL4pPbAdQJDHdiLzb/yc6ss6SiXe9jm9pe4Gv2kQj1NBTgdedNE
BYeM2kW+3/PjasJDj0OPAsioNRaV1YfrhoD7+w/WqoUd+CsI4yjLApZqSdg3HytZ
xKNncawOeauVMjugZbC7lqBrngIJUgdwcpzUyoK8c9vuv3tm7Fyt2K6NdAWeMhxV
TPRgGCVa77MHBmJGea6r/kruLh/CeecC5MB8nzAee821O9QhrULh3HKZLmw52jNt
CyTLm1AXVYTsl2WzVdXE05oVepq9vWbUWeyMLVLoCg0UMVyvisrZC4wrNuH4D1Q+
/klAXNH/O5TuWOKxux/JSAbjw2iVf+f1hfsh2TcDnh55D4+AH+6tSEPieKGi03RR
tEPzgCRYbkSOg8F6pjfNRBkS01VRkDVVc79zcbvACiBUYY/3e3wDUDTjYcJRMvNb
nLAOUK8iMQvAygi5q1tMqET2yIpOVJu7tzXaWsE6csNfADcKy6lTgbtwIMhWX3KR
ibrY0h+dWuDusjLW05XTcByJ4qiOIfo9aJ2uD3vt6U+DKfqzPCCgYhumbWQTYKN9
lDsGmqkSY4WZTJ3zk9IL21qeqKbVteGLpbhi9xVUs46sXg6ksBNbzWB9U04zq+E0
t12o4rGS80sihNlza5wiSg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
DMwMkjjNfkuraKa6a01RihYad4UVOSPF9UAnFHH+stiyn548W+ZzFaHMQEJup1GI
iiZjj8mE6m8Ps8X6p7wn+mBbfB11pP0kx/rFpO2PqbY5zLaEcS9R6Rbd4lxKrYqn
K8Cm4jv93u4BNcrS6qFh/ZVNx8S7wD8ubyOsL0O+t/voWqlYtHBM6zFVTJY02IS1
z+P80oxVbFiPGcx/TgfRxc8lM7SJYMZI5UuboZpq6rS7LXXH+YKvxd5wN7naaVMD
hmfVZuwFMeJ0vxpQ/EfJetdf3O9NL9KTZ192Jo1+d+BJL19VUbZs06dO6vuQ+SWW
3idBwgl9IreMd0IYAv0lxg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 30960 )
`pragma protect data_block
PwtGar+QJgdbX+yItKf9GqTs7TyfMTmuelXOPxOq0wrjbZ0sXJwPQN9LcQAUPIb9
eNWgD14dn/NRQW2T3r3AdOQ3HFGrR59Igm4VLLE5Pu+s6gtv7oc9GLNQyXOs1QQx
RhmekhooMc9fPA0FIJoFS122BMOb02zbOZAqUs/Yn1z+sgPnmCVZBdEPBNVWV10b
vnTUWx9osYhXjXsofQEANbIy1co0EdNvg9y0njs0BFWRJO3wHxEbBhbsNzFSlMBu
/YYSrlUwPfnNqcW9Ks4hc4ZVwl4gKT3AK+6xcV/Iqth5gMvWocsmHoitSrAxLRo6
2x/k4OTaCrcta4WCFgvNmeZOSKfV/N1MwrYlvgsyi1t7Tmo3/LMQ2AuN2sLkj8Gn
JdOmisAnIVaCMO0P4ZwsY6zY9jaVqHgv1GupDntcU2KXESLn1bmASVr8DP/Mvs95
dj1BpOVdALULzj1Q9XADHEUxTcqfHIav0CiYzUO6D3cRG0dmbUC64PgJufm8uWHh
1J8MnynJyPvc2gs9dIorxHq85huQ3OUnPgylfSXFbqfXRCpS3SkNL/VaINfbNMWl
u3E3O97cWw9HnkkfYUa+vBWMv8RQCM1ZJw8RqfxlgN0EpReYDfhyMKIgztozAkJX
FOBB25KbTwhonD+BDwQgW+yFJ0h1WMkjB2/MH2ogOePS0zbqPKzsKh4cnjs1ifq3
3PN28td5gGvQPZ9K9kdCNKt6VR+xaSEe9iolwMic0xlcz2rO4l+zm2k/KgfQ03bK
WQ50X7HTaZmMCKD/2LhiPgNMeUUQIh6lf4m+VMfg1IfuFpOFF9Q9n2E7PKNbyZj+
Wp4Z4dAnP4s/HReDmJLyP+7+uL+4vbTGOObtQejVxDiuyLt7PfVTsGV+ixdTy/lI
WKgLV6RyxyxxsiCgI+M39PHKEacn4xFog+cm46cL4ug7PsxXRD6nos+Vn+PyouZK
NlThjZ7V+dFLxy26pFgSCjS3WgN3SXrMADyDoi35HslYWeqV5b53AMBKgGSHE454
dTleBRmZ8+F3AEOiE0Wmp5esNZeq2aXITjPe2Zxk/1scGg/CAteOUx6KE5tPHU9r
p0Vj8Otwb18E0tlNTLeijur8oxrehher7LoQ2YgP2v/qfiR+vmY5YzGUQp3DagNB
GPDyN4ZcIrNynGl0c61Bwybq5LIGyVsVjURe/V97RrqsumW+5+SFO8OnWOiraUkq
cA+LuWbWjEKTuKafhzj00fqnNrcowCMpNf3dlzxm/dpZNFcQQWldwMIevgPSAJby
f24CHPYGxjJRAKquHmvewIGJHCf8QsIlfwqlRRabAqqJ7p583aeTm7v+EXZNqc7w
LhTc58lK8povABaQSIuAfhTW7T/sfSqpe3NIJvQ6NRF3D0TFUBiRAWNeEw4xp2Rn
G4N6Yw6KfPk9UFr+865rhNsNS6gaJBSumF+aKwznPlOF+T8sKo+YMNtCVRi3jBBY
0LMgvzPRhTIFpNT/1gWVRMhxu9CHng7HFjvcFpnUUFHKHW4iYCZ6uI6Tnl5IS1sl
eQB9XmZ66LMYty1I4zLNI5JnVhFrfnih9BhiEGH0gvNR9SBws/Fw0+ueMzIbQySr
FWejIpY469H9Rg9KsiD/XgDvJZQojW7Ts2uyPOKUQdKd1UFusOU4alvFC+l5PbGZ
rZubywcoXiTS4tLd1sWVYetswBSuZSDyj+nntui2T13+E+YeQVOHjtj7JupdEn2l
s6keet8mmuz/8t10kYGIjspiCJkzPff471hCTON+aOb6ldAiMPQq2UA/zGdA8Gci
3v2kq5phbzFcIpL01NrkkZKTbwpMdz6jqghgnr6JxVsOAxCR1EroyoF/DqKFPFWj
2D9M+E6hrk7l7olV0vYeBLXZb8CiMMHqKr0PgCp6wCed5DlxWvGXROXPRzylplyf
1tyZ6BeFeOPp4kkk0q63yt78RSzlieUM0vs1OsXo5ajpXXLsL3p3MMnl2PzhLbmP
xfp5hrIGbfJFXKjx2QguPm6Ea85FU0V3940XtLXDdDpX9x8qM9/BVt2lM7QeA1hU
5tGSQulLN+HdBOMRQPMaA8UD39F3+jv465+lOIbXNJmfv4lMIXDZGrP3FiYObxWR
wJ0XmMYlgaShMCxYfyNpr/dlypk5TcISHxRpeJcbTf1YM6C/BWJULsmbjnz5XHgp
iK+rrVMJXJ4pQNpUJAq2zAem4cDh2FI5QfjTb/JM9NVUxUQswUFdpz6ZJUDaQftp
G2zPAVInBa+wCbq1mu1yf40b/RSSEBH4J1RMxda0z6NuyIjjywuAf4gngr2qFM3y
3TU+1hEf8lfaGuNa8cpnbWuX/QVo1dKryvFjAN+jflllgo3GNt4h3O2QZfYkreO6
WyBLFqSXACcX7I6493N4w9vyG6y3TJylCdzWuWAisbpJQmI8lveDTubYwHII92fQ
elMnE/35gKUOEh/UV636ezVg3EkY3bq5EE99jjgu09fCttEZInTgR2EmbSmMdiX8
cAIY3boRUGc6IgC5qt0BjqdFiKf0XB7vqSZV4K6Auf/A4VewwTAizm8G+vNsD3n5
DeBujm2YDjlVN2fY2AvsLqsBp7IAlILEQw+XGrafxorMxHWrVTTetAIFFnO/kn04
L88bDZueGGtBgCDyu6I/cyeuxkNFwf93yzk7A2emN5sYLxUYjc8qF0oGd0ITJjoz
9V0UW1zfrKNhomNSeO4GCxyZAoTcAm7ueMGNaxJkPfIGPDNMB013SpBY38EbrxnK
A5jbC3monULlMh9PivW6MLZKF0/Eca0HGNXFUYaF9nsYh9pAbwLyuXHeWB7G6NQi
quynbv3Ky38cE1QFRfSocDCBmgq5HMyztk9bpWHJF4JgP00TjMFSqr7HMKBbOSUe
9t2nR2UFV9FPP/abc6d9Z8qZh8+VCMZWa2drx8uaQ/8QOHfXvM5umGsN5iCWMz/d
mK2bhK4tZItMzFmHGSc8yAFBog90N5SS92KjKZf75QSzqu7FDhk9hNr3VnD0bX7M
Ra7x0uXwIN8aj/nT77R5rxmYgUic2XCjSiodfT1ouPQnQoeJmyEGJN3b9WKD0dyR
0QW7eHoxkxxgsqiM4ddUbDlKt2D2SZ5K75o2bMXPf2xKvcRpL9PoJfdsMWMi8nNy
E8kE/a80Bhpm2AApgdXn/ELn6rvta0ZZFvC6Dbs8xYhyTJemQiTe+tmgexN6I8RR
wV43vfdgLrrP4Qlo/Ap1tZEkGSBesz/7sAtT4gewpsPVVogiVSdx29eZIAgNwm0E
O5+aMQ8ji5U6j056iWLXnSySRY796djrJ9poElz/rsYnlAX8sAyDS4cZdA3+h3Dh
7LlLV8qpt2B9deagsQ5wD9SlQ4ZOW5oP5K4dwWOmh6KYaUKzobX+UojGuryxUEaE
Addy+ne8GXhivzNvD5sQQBBEvnDoBZGpy8o/ERVYWPfVsZa42KN+kWVGyqiD5zln
ynuIXfxfVCPcBAQcag+DNqbMruf7v3bPvESqfOZ68VaFEQiOaYT6mvJ33giJEEHa
urwTkcnu8WGOPboGGXEYV8L6+yGu9msKrabD2OncXfYZxk87MpiwHINpfLL9Qxnt
n1snQiQ2XKKvbhyBVIcPaRjlB1IWSmDKruBcQmF3Mw5GJv34yrgXdprPqaNSx9Ku
PRwU+5g+P/+QJcDJamEhL5OPdsO06SFNRJNd1rRfYFV4QzpZVTUqjM9QJ8YF/saf
frBs/RBsZwZyRfq9xOZ/I8pfIvi9Hj3tX8G8A5KnaoIYhf06/BaIaYGQOl3TJE8i
3a13LxgHutntM+XaQzANJaxsZktIUdQNyDl5Xdm854l0Wyjs1GbfWB1luFb5MjAC
SxGMJUtMyGQXQJf9r2UhfHRS9JaG9smJZekY7Gm2bQFof26WmyHyzaWXNxThh9J0
dTjVOubMqxe/Apw/Tn7F61CiiwYHyCNTiZU4ncGEE2pFGTtCW2+8fZSrAhoDdAFG
UPK4nxtUPGJnaDZlw8e0B3mYN9OXUXsYiy9+pAnwdgflgrkSoDaRGJMDmO/dSAs+
N94j0F1Wl9JJiQsAK/o8vqykSwFY43NXxix+7cpD95l8fQ7+YkktfxlbgXgj4q8f
+vbo85/p6olAWkcFwu8yQ4hYT+v0e0vEYXKw8tCihziBbmHIxPdzMZ0vKvs1AwK3
REfc2R5kZl43e8exPj3V5ODchcuI09mEyW8S/wPoy+aGF+cI2Hza6K09Me8zN0JZ
WdBDmczHD914rU0SUgHfpRMbZCJjFGxXoAndgkJLYC9r/fEdq+FS1X8xfeK9qhAs
+jAy9rvFzhQPUcSKRvX6NUDBnIHYc1kLP1V//zLq8kwZnEcU7DhIjPU1Qe89Lwn4
R+bz8GPMlUdrhS1nSsu0yvd/nzcl7SjeY/CIYm0fUyQRmZ1A9Ymsal+NZtpIkCd9
G7ec3+2+I1+bTNTpQFVn4PEZ5yvlZ+WO+vDOeCFHlg4y294Pw9rQ2GDjQ47yq6Qi
w+9IHdBJaTUk9m/iV8cw09XnA9XDra68/VBWQ1geY7D52m5qZ35CR+Ft56c2H80q
0j0amIiYSwct8yWE3CcjvtzIJlcPaCMlFYlcuEUwbpVnL4IWchg1apvIXkRnJp/l
KuU4jS1UQ1HvYUZTyZaNwjNOHH40AP9qvag2y7oQ6qqvslra87nckKnFkoPDwoz7
OOzAnU3XWUcXhtgcBBEk52pdxv8WQTiDVnva/3Fcg4p2hyKz60LwlQRimGSB2ajz
3troMV7sf2Q907q0lYsqGgmSmoLXSNu+0oD4wXA/KzgB6/+pC+rUW8HRZSopiYQY
nS6jgM60K23oxlo3e6N9N10aBQX2DUVOeVR4v1P0LHe79d8nci+vd0bjDYFBz+AJ
kTptQjVqOIi+l+h0984TnmF7cloJbOOkSel1jUWBqIcdAtXQQJvSBlaKW5nvJYUH
b/4MwWsokw0REy9LGb9Obo9XFPvsSD4D8dP/C2bjlKcQ8O9K4gxQBh6g6YnhlDUN
bpMB5nFMa2smAC2ewdhsLia5u9kYfi4MJGcg5cBNzCKijKxiYkk5p9/921/kYjwY
CNRmdVdgMronjowPSybwCfvqCNMEhGthXgRyAVulwKYhBfDXPbn/pV4BBqqIQj5h
05NGEadyK9PtJq6bDvUBmSgRSMs4XQ8QzRKODu05DVltx8ikggzGJAq9fnTjZXUm
tfw4CBR4HVaJkfGQFhoSuEXWaiYQy5xBhWrirUOqOLT+ppKVolAmilQUUXI/xebo
CpB15q1n01ZyWn/vaVM6544HhBeWu+dHXnw7Mlx1lXph/UzF4KbNKE3xNLJNkz6D
71sJo2eW+Nvqz+4zkIrzFWlEJCt6UkjSB2Uzu5GTzIw8AUNMGZKd7jPoPRBc/V+s
EdO1TIGl9zzWYU+00N9TQKH1PrDcp3HdX6txgxlPbRjEpfwvnO+f6toZ0KN39IhV
q4ouoWvrbT0DQKhdo4PLWlSawBlgVuCIW9aQdhL6BQSigwTDaSVCiKCcO0uTIt2G
Y+zW+kAuMZuPc5acXfK3ngTphrOnUeDXcSTALdoKoTZbKx4At7C9ItvgG6NkgQ8a
ThPBn3oSJ1QW/0iCDw5ClJAtYesz++LNBTmDQI3LaqwxQIzR2EfAd07YHpAL5Xkb
8NAYEoUB6gqSKiYoqezGWd5rWZYTpVEB7PpITZmTVqnPrqa0eJaGJlRu7tGCUYXH
IqqtH0aLuQBFxeqbrmooXbYGV2Swl54BGSs1vpUw4jvmI1blZGKqPGZkwlA38Fmy
zdLhIVjolivLM6e9sQt3IqcJLQe3ReiLNBS14s/nqxJJt7k+frhOgR0SPD+a3sBD
2Yt+6SOrP78F5+mOr08p4eh3LRqY0wwEIh0CcyCXa5kLp0R8VYj7f/3wt3X0weDH
JDBydDfAPbGGPxWKc8QCjMgTlLaok8kVR8DhbP1evjkXOw7LzmrTUx2s+7+tGK83
0bggZWArh8KZgAvvP63yvTaJz3IIL6SLDbbJvWYEhel/EwT9yNcWICa7+4sQn8+1
BqFVAaHB7j5c3gWvN4xwDbbp5SQAUiafNVgUPeygm8Q6MfoGIKNKfVTYU+aDhXxN
Q2ZxkG7wn9xqWLR3nJBk9cNXKHpeO6ClnofpKqEHwjbkwAPVT+lQFqqzzQnS/xz2
t6mysfIEGTJXtLNGcovCGFJmDV/A8az2tSSWTW7HPHaD0b50hf8b++18kjwh6xwz
es1dgeTkD50mwfsCXDPOvJXrJEm/+hMD1jmDEPZVxgQlOPnhROsrq0CWFfk2wTRX
MWUJ8sEtrN3i1bUNXXQoP45CXIbsWZewtG42PBwOUL3TsA55iF1sRRlFqa7r23wR
lxuvdY/Y4+iEJJsRclSGycEXFOvQ+4nEm1xnMRFerv3miadTMo2FgK/wNMKx2M3M
Bz9Dpp3hOwS+EJCPXF8desVEJyKLexvfM9LbzP/1jneNigDVWwZntP5GJ6emy4d2
aS598Ij8XxQ90h13N2QHOYDAQN0k/pSFadpByn2KA0I9XbZSlDH4i3RZnptN0/4o
SaBDrDSSY4sYJr/ZYBtrEuoqG41ozDJ/MZVUAsAiYnbn0DpypU4ocHM2lm2DoTVt
jpioAOBRk+w5wIUzlK+uww3zhWuH/ya0pDkclYNPTb2kPVvUkee2OARiY9xhWBe1
Yfe0GlPDhVdk1Sbf7v7tpu4zTAPgny78cKQKm72JKwExJMga+HrovGD/XhBapS05
poNep/Dg4Ht4U56XHgVomULVwBnLkr9sPQOpolyHscN8e8I3JgP+fiuWBA9tKVGV
tp/3G+URA8vaAb7+Q28qr+XSjsXjuR3jitqVhOjQBAhv9diCVkRM07NcJ3wz9vuU
QJFcKgG6e+1POvKJReSRIZ/7IcZwxN/qLd1SVCcgFx8sPq/8AoTGqwuwSAf351Vk
mtOTQbWuNkMZw8v1DuJKBekPnIGpJUvgMtuUYpbddeBKkaCwMmJfxE+OqOP05kxP
jbZKPFNN6k8v40osNQvSPRZ0AUcTyi+55gKe9dp1hFtjX1/KYU8Mx/LKiYRw7flJ
39/umdQg3Awg65tXzvfubc1o0gHPZK9NlPbfYgXvNqoSU5Cj36ZMtyOe/gVJVHJ2
nnz5aygT8xXlXTEvEdEkovlA2+IdIEy45pEvwy5DwuwTcrHlE9KVcV0iIlh2r6GV
oC/fZs/NIristqXUBoST5erUE55TJwbOWJlXxJrTo7pSkAiI6nPU7GyXhXsPToUi
cLUAVJ9ow9w3dWH8hI+q2AycDD86ghylPu7lx7tA9yBiQ9RRZph69okykHiM4McW
Y54+h6rpz7nyHfNXV/1Xl9vGnXzlC0L3UW5JgUY2nNeKp83ZV2lfAbMuvRLVwUT6
2orzlahbKK2hmV6UfbpLyi9oEuBLoIIRzqKcymYh3JCnnjdP3dwKt5kPLOeERs6J
JmPhkHhjG11wbMZFa3iLjqdRBIvMXQpX9P9VzviHwCP+T0SKraY41sWfD9MhxoU1
FEqdqvJttT7oiTAYS1MmZEq9FJnyWEeCQQv05pBnayxfZA9JXMYDhCjMJzjSCkXv
WagqkmvT8KZ7AiYtDD4XewZsvCtFOQU7lzJBQxt0Qimn82kgbrV8lZwgVM93P4pz
5/RlGKfVgGb7uf7Pe6tE4HEdVCZP53se0JXMHzK6gu95Tc+aHayXwPeGgY8TyeNk
PiKpw+8eYx5W5SpbJR6i1kPxwKfBTJz6/6ks2+1B4jFqqxU95U/aFR0mrgozB9Sq
OPzslV+OzU/Xo4KYH4OUhgCbU7OrXyi4O6wF+u2itdUEa3bgfnQnLuDC6dfVmeVI
GgAeO4WCKc5tVep3I/RNsB+DF4BsDjM+VLe3CzBlvE827ydDjzIGtDmsEzTancEV
R2UI4NG56cJXsZjjm/PdfcimKCJb1kXlzsMn0S0MBs6HP8pnWZNC7YooDcsag+nw
3SkyQ1k6UF8iLBnuJEZNLBf9GEBO85ysJfr3XrVJvT5UR5MDUSYuZfsd8eH0GOuw
9oVeiXuuJ/4VOCdtJvMwAL4Jy/22OAm2KD8ZZLUCjzqZSp3pf8OmpCILMdzIepzm
2bEWV4/8gjn6WYFX5wK5kfeermyP/BxSv8MZm+crEYvsDGriWYXz6ju9bicr61ag
fd99sPoKnQgYStPrlh9O/130upk11BHYIAD+JPPuWtRaFSqjWwCAeFT9qL2aSQjk
2W0YOs2msBxXcD+PVqs87BecrwH/kRfsFj8vYQv+lTGnLEcPK3uCpCWBqDUPmq5K
AnTDV1V2t2dk8CtrXV4wFVIqDm6oFm5XYLSI5CjeRMn9YoHd1EN2Ohfey3wvCc3R
kuClVZ5+Znvk9stPleVfhFUbQYUgqiKSjOuKmHb3iM0roytE2Or2os9U9jw9igHD
9SmuffeFPTli60Exhq8QyQyj48n3Jdb6SAtF4fsh0ViPDdHyKn/9fAaVV+dstT4k
ynGJ16cVzPKQZ8wmCSrWIHuN2iqq4qdKgoZAfiNUT+QxAMtcVm4oBHQwJJF3+Oql
WAd07+Vj0hq/+DJMTGA3gQfqTFs2bFfoL/gN4yBP9j/pOKeKdhbHMqQaX7aBiPic
2MZrO319bxIv25+Gh9Xfn3o3Qwj4m0uifd8hOgLOE3A7XrfLMo+AKwrUGB7hX181
k14iStt7N2b4GiB78q7KjwJ+q5cRekAXEdQtB5JGyOf60RVBUYZKDhkhoCjgVwoG
CnFqY2hwCDR2Ot6C7qd/7fTWE7zn3g36IxLuwsCSwBcprUnqXFvYyyWvdZby/42X
r2MKzz+XgN6QG7GRCpdCIeCMEc91jL83WkJCmQY1VETLxX+2mB690dtzj3SgeP3t
f7MhFj8KpnZUi1b3nUOaAjhskbGVP9I4zGiLfDVYfvQ8p7NzuJE9ahLR/JJtB5gc
CFL5+TXEIF9oV280+RHqEjrkyjzj25OAJzi10/AKS0AfgBOMv3p50Jv1tS4aqPFk
5Jd7iRgAHqsK2j1K72gyaY6ruhhmnCWaA0KiwBimpXX2KcMYQsU2y770EJepQyDv
BazaceYpnIUpbNlYFAyUtfsnFvWLrvS6uLEPvH23PGyR0xLoP4T34H0hJZdlLBCZ
JaugIV6ZcE3ZEv0tOxd55slixfiAwlxa8HhD3fgiukStcPk0/z2rLpBMnDm7mMkD
t7z5NraoYM4Pzb0hRMkq+kDX1rM/47ytLhFAb2Gi4ZYr9X/TqOH/hkvXPTy/zJBW
F05nWGUKU8Z1C9kstGkKMjESiCkNjV0e0Wwgb1R4iRPf2Gz2dmw2172oQaCUE5yp
epey31lAL2SOq2bLfV+vLkRlkrafZiQf5LTsdoehArzfuleuHcC8k+jE3yemiKW4
kWNOFDmh6fHRgJxgjIqR6vOiRuX/LfjKoH/CrRhdk6c3SWnzIojhY2dmrhYCiV5a
wGIuxJBLICNg7zWCruCJbDZf3/CcL33Q6jG69JGM0futufJ80KBYwMcDy3bkW25G
V6jyKDV9y5UztFZerKAyShl5WuckAlQd6W16KF8L6Rr2b2Gd6Zbnju+I1S4yJdHt
QReLPGVrLBPL5iC8uHMxvaz2aboSETvAn0sDLVXlqBUzPZrHElkzC9L4+IDMLJ8u
Qa9FaSSb/OhxMrkY3GC7X5OIyNJlj9ssV5ka1a4EpuxUmQc8J2YGLYDNQ11X2EcG
6z9xPo09WJS2sLdEAVHvhr7rcjse9qoutzqmP923fq1+YaabWrTuiYKB74VcAkXC
KvlDyBIgHX5sdabTzrAvcm3mrwA7pG6rAilsiAYWVuMuW0mvE7eTZL8zb2JYNCbP
0D9vvOCfWGHp7uoBNOmMl+iNmFglXxoKt3FWHveLtUjV1wS2mwR+ymZp//rnx3/R
fqBLE5Z6RSu6p6+kyRXjdEB2LJxW0JjY0gFMoTkO6NigN7d0iJUN5BZtIfAJAglf
Fx6ISIY7C+sz3nS3yVLuJjhEvCOGtxHHtabDVimv22rtgU7ekOoAtGd6qzp3x4hO
0hxRTkE1KWFfl2JO0TjHbxy0Sew8ngVETMTPBhaxICQABKVfWIvIGkoq3RRl7pCI
Ah8M5Lnzog1U41O7eyy2KK1Ar3dW2RvmZQQTAr8anV17rrGFS+Z58ga4cjl45Xwp
lm9aKO1TaRj5DNaefH14NC6nZqyMFh7MmFRlypFV8NXElfnZ0wJ12TdR+i55OHDV
J3FC0Yc/i8AExf9MNIbyx75na9qr1xp+s9DGJeaAfv/1+YEs+eFiZzKgXwi4kE9B
CbWmi7dYeRKSE8iLBCJY+r/jtgbGhySstTRoGbTXITj+vwX4HnzkjAO/B6J159+r
tDrlx/fb3yoVkRjabdTigAN+I1AM/ImJIc5YZC3AHguhNOhKtqIOAyhKfJGgCRIC
C1/zLVp/ddZlKH3SyxhEaZHIurqFGCbmgjqhatYBFcXMayfwLbzNuzibXxColU5q
GL7DweadcZK9oTY+U54nyaXwWPqmP36VdWMmjUxVHJU1DdidFa7nQxH8ONlWR2kK
nwQIAQAWT41B3EgPkwqgaEt0Cyme/A79Htkkysiu0Hkem36i9vGYLRjglWbEAQgO
uSSppQLN4okH1T554Kqb0ykT0U9e+tsN1Pl8NUCInazQP5rHeV8i7+s8npg9hKT1
5JAknnhCum8O/HZfbYQTHdKjbJqhpHkjkz+Br0MoTQETs+2QI9ChJjrghtUNzPMQ
LHXzuC+eWbx881zktnoSO7gU20KCp2wB3G7wkTKd2eAkstayFWPAgxjkG4OZzbOV
ASyA4Piew00UC4+6qUKfD4CZzISUshpiAMTHn0QO5MmY3yPKQ0guwY5mbVw6/ZE2
a7PjZHz32O+BMRcu6zC1RYQZNjrEpWi9IeWLATpCbxjzONz2GPp93y594mFviiKH
RHmKwl0yVhqlSfnBI8EBABcvqUptHs4vBuwGwqrk/AAdfyB6rad623b/pYWZaFZW
PZ8O5xHFCBCiU00+XZ55+/FlR8ngvXFA1xV3snoS12uzl73+jGFacfPQWG/eFnLF
qsplA/spVWN0e/RYcRCAGjeljYTa3FmAcWG2tG0noF8T+ALpGd37ExQAcnsj0TfB
Zs8aQHYYHulowI/pH2f1veK4cBjuG3eR/P6XYS/tuY6dEHHvrgchODpi39as0MYG
hbDUWqetSV8SehOl7xAbY9yM9d6unuXSxXEalYFqSyG9J0bBKTM0JJ3kIiqqUSzK
ugSCGs7YIkZIK+ly+PSLIjNTR+6ApozLq6qYwcCAlgexHHY/dISbJDPTaydxIwBH
z6cFslRO2yuFrQcVL2S5p2iwlIE9YDidzIFkKM6X1EvGrubP5cWOLsJbRt5hGmkY
lnUEyCghfcltyLQohHqMIXOA7o5Iq8QFy5qBWoZnsqgNuun90XSmqf+Tx52K6+EH
PaF5RjyXGiYwmrAwWg1Ypuxt9onlPs1UuAjypaCvrE21DWVkqALm2/57aZa7Mfpa
pWR9IpUhdQq5OtOCcBF8N8fjHyjr/DZ33NExgjhd+2GCO0HCS1wl0sjGtPaJ4SHP
5+EGQ1HP8WyStLcKERC5SO3ALEDNVpIYmtI+lezppOpkqRewZArqLmhswsVcThqw
WHw/ZEgVU7dUWseDPRYTMAIV0ISG/YfXlFmk0EhVwzDdZlQfuSSwLelIqH/Qx7n1
u7AYcM7pyZcicjGfjXE20evKCCF5DIP8UG2B64fnpedFcmEZAT4S7QNoL4EZvBBq
qhFF0O+3rAS0+HbgRDTbCtliiyiVn9dfJKxgCTEqPYFKiqemFZTIEwKXaFWzpOSr
wBbV6FnyK/gak4POsBwc9KzybB1ax22nFlpFf/0823nifxBHVklPWy2LHdcw/8W3
SJJ6ofs3NRGdHAFHcPskMvg8alRh2d+Mwsx26ciwBf26MPaM4ZKg6BAP7jrEE6dy
6mM7LG4++J+/UIcnIVIsRNSL/cb3Ue2YyRRaU/PjOcdVjqzLbA+aExD0nCM8O9yj
xg6R5JhMMs9+xebrqjtDNT/quHXJogbjbHA+XKfPvqbGVp62uyb8kdD9e0bosbD7
X5FTxNy8KSpKwLWAkqu9/InkX79DyS7gvlY2N/R4n4YCBWVuHDg6WI3T5CHStTPJ
Eo+pd+ndCY0KsnXpyAYLI5oqTdD//cDOmCaAzduVvO8cUFgF42uluLRBCO1vj8X0
M7YBHQ/s36+DcvFCaH3uPX9zQMNIPXAVu/FvN9AzoJr0zRBMiZf68hIk2N4Cylyu
cg8eNPJQ0VP8F6OamA289IA+u7PWEiR9AAv2rjKCC+EM027xVcVj3rnFaFG+D2r2
8GyiyVNnkoxgVOH2hyUGVBYqROsEV/eK40f4cVqn7++9YMRONO2mNwx++CSHRfXq
d9S/LS3JU8WCMamHHRJsbtcrGp7nxOy7ng07T+IqxAV4vlfFvsjpbByCAZ6H9iuu
ZJAb9XF/Ed0IfC36xJWw5JX92r9qilsMctMgWT5rLos/qXEYUyjTUFpTVdzrOhyM
Wb5MTPQ13k+wzX6WLjhJZnwKS9LAyUq+HQGHKFEPrS9djhAosupKhn5OAMsvUtKA
qI35XzrMuoczHQCp/QbN6WN02A0JlQhhvK/Sur6YICDW2Yz/QGj8t3IteVhXa3A9
/1BNEc6ST7veu1GXj5MBxqNQlARtU2UYY7xT+6U5bxLXi/xPJw5G1aVPai1iTZgC
E1ACB1coZkZmK9bQdkpdz6mBT6WsphaaT+rhpvCnF64chinEwGniiZGnjSdpYfEh
+G7JdwNnuq25J+2hMvC4qUMiDPWPduwgSDGe3pIQX3oNACCdurBTk8qJyKRlwk0+
yDwwTguLLtSSIURHtMS0nvp2HPnZef6OpP66d1rN0o8lENS+LOL1UfUiY9Iv+Jub
OjekM2bFHU3rrF0dsc91lMeBtfojB6nuyTxSqmBezq5TyyCgZ7CDzW3StaFnkEed
8KdbZWGa7Pk38AsUfL6DBasW3ccldWNFT/sG/KKvEolGNQ5WSx7HG2031Ivv/Rdk
pNVVH2MRxrTsPzKw1PRWEn/VPlErR0fagEDj6N19TI2MYVW/X0cr/NkPS9ouggHv
91CfC3neOQfHeTOCrSxANKYGWQL3y9lBdvAEG39gFmKcGSiZjRCJjOjNfBpZHKn2
Ex+0IQjxc0pa62O3UMquBKKnCahhoNYaY9XZdUt44JS+JracQJq90GFRH6vDkMTT
x760sJcjrLzJ3H4BaaMWR46JUtyfSx7cI1N0eLNotumsSBVAmia5KSQKwx/CtiOM
2QYU5qlTLovI2K40yIMAq4dasltgT5YMfpSKyfZiurcSG48n61RzP78MbYbd2Wq1
Qqpwq5O+vz5k9muDxAhffNB8fdXEQmtIFFdCp8vZGmsGsknZAVQuAPavVvUZ8KMC
Xdx+3eca4StGAWSPprvD7NChqpxAYNZ2GGB222c3GV6bJKOxiWQdUuJRP3sJxVqe
NrB2fP6mlbEKOcVTfpkuL+3ndgGk3St4MYSdSf+g3KzHLoA99MxwWrE66wQLUgEZ
cWDs25+3dEF7cYybDyylm/QVRJcweSSE3zfLnFknEDmXy9TZt79BSkHZw4Wv37+9
YAgbKeQydmTnBvTn6Gz15nF8DWuOrBS0SJYIpqV5rL1TV3B4KSV/9tiMhDmy8ZgX
pYqfZKqEf7hbxc5C8Jxjcm4m5JMwhxxrf4rCIWDgzdDItBFn7vdPhiEBcF+9qpIf
YeaY4DizHkhLglJf90vghFwmR9G513TM8ZTXbKK3xJVTI+9ynDOM96lA+IkRCUUA
TeROFTkqsEG2+1pSm6L4eGGE1uHZqxF30DBQXBWZf9ofCOpvWMbGkaB9ney+CA+8
oE0HCQCtHXBTw/o5dPVs5ZTBDo8wSs0jlNFNrBoNy5ihB4mfQ91IUGVmZAakve11
8z9PGs1E9T94RvDp7XJ5FpByMDi+DnGeheCNgt0vtVjkXO0uLu0ahp9jNy1YbWYa
eiK0c6YRpflyi5XpOVQuMMeMgyZpAVdFqq1XiQEE6/6Dic25NSU+RnebR4zpOn1M
VrmUi7pd8iPudm4Vr//9l0iLw1Y/wZY3Dd4rLUTXyiTNepu+JMrY6LM2ou9eU1vb
rnoM4jLkHqUwsKb/1K5a+Hgw4M4aYeu+YgZ53r7Rvs6Wtcl6YsUnknDcwg6wKozA
5CAB1DGKO69UCDUERjV09D1HOiTlM41TrAaxzOSaiSR0rOdKSX3eeeWWIWNeNASr
sjcdAHCwbCmUbORhTqt4PB/I7cNXJTqtWvlGIt/eHRRDPnNuSz/N+O9QTCklJg7a
mEAWAJ+jyeJ5oVtGtFgvXz2RS73ARpA+JY2ahSMlJ07dETiWGaDEuJhxToTwppQ2
sS4eCGZT09iy5u8IKyylUr49e6/hUYXHbTq5QY3aHT1zjr365obpzT+9fAsJ3LR2
J0E/GNZRUcFKs4y6smOcxI3QotREQo5v2g2OfQh1sjAPE15zqqIUF+b/hwv3tOym
eEvNZoIGJkrXgUrN6gg1ythbvjLHXkuEgbWXBr1E99N8OmUjIxZlv3AbSx1xCwDZ
207ZpwseMIVBOxQkLd9mb+UB7OTgd7E6tYhE0dF1bcYkfDfqH7Ga6+qWkNlniO5A
lZoVNmqvgwiqalDTYY2GzW5ZCU+gGSxRUEnu1GzM/DMt23sZBD2tfqHxchYLdFkS
uZkzbMH6kttHqmA+K/na8+bb7dU7STyJYb9KEtql88+HGLYuomWTJwvi/M+Hh3eY
C5LnMZsRRrnOtEiC+GE0/jm/koUeYbmqUMQW++dOA1kh7OSu6BaUX1WCeTbGiVaN
/XXTwyco4owK5kEASCuXNYsvwswOF1Wc+r5FUDzCg6RauHAFJuVO5Rq4QzftNUtR
uE5ynNO2+ky4Rn6xkqO6/+ADvZw2y2ks3kKSPrrOATE8AKtB5qCJCrXlPFdgwfBN
6a4zgLLQGZV9Lo/elEXn/bo2vE+4bdDfHhYabL0N9rlvFLt8YkYb/WvVD8rlkR+D
KawALxAorsVV+Tv/4BbfLQZuNCAyQ5l4zscVu5Do+LjsFTAT6onAcGDdgk9BQw1f
Hf0R9JKh/pqy4vpygz6ZZg+KJkcGgPEu+2eANzNN0gGgChNMBb78dl6z8tvHYaYo
JURmqXDHh+HISIHiY277SUrbTFYt/zryLfo3DXP/axXmhqrMpuAxyrpGM3CmJ43M
tnMLkFlO8izyfz0P4kSQNTQq9DLnanwt2/wUPdNbvjS9Gdj6KkJjZ57ae0ieW3qH
h3AH1uo/P/C/rNBk/BPoQJ6oUSzw2lMicfQh8N1Kx4u8Etg5CdEgcp+MXvN1XM9k
nQPpqUHnjiD/sHlMKeNgkD+Zwwnt482sq5t8yf3qfzOmFxIWiLH39Cep2pSqBXzA
mPzq9sD4kid41451QunnsNVnrBUuHBIsmEFfxgR51OsCE2phKW0VHCp+UN9cH5rB
T6ZMtbbOujl4RkBc7Xo/IR8y+xfe6PQKgkNc+S3i/hFbq4bltisqQrUv8pyMApWs
dxvX2evTnnyAAY5/GTGZn97nSPW9DaZL6YOcc1bvNS7QGm0mqgIX9/5NagABM1aO
y4pvR0UKdqgmVcxEK8Y+zKKUAf1GT2retvZ9O2oNHN3K5UWtoOjNzilFPA6N1O8F
RmFWJ497Ll7aPLl23/KITAEsLo/CRJTKRLbHuVKFMEFuXm4WCunKZeTWz2Ong3Ou
k10UCcVHcIT56FlUfUD5YzYh+RknKtbhT08h+d/bfSbT7tPFoUeKie5HLSikvTTV
LNp7WZn+4yTrPgIQV5DROvIjBUdO7kMp43evr8kBxZ9Z8NoTr0CpvS0nYsdQVtzm
76RZJhE/x3tVgUmkyjngz9aZhUJLhPUJVNmA1PQTjedC5dnxbFal6WwnGj+XI8nc
6lPfzuNLWe+hoBCHYuj6SIc9hDtBGcqzpcUpzE3z+g33DwcpHKHyyMSxMssBSXWd
UUlqO3hR4XGJoHNMLjVFKObj2pQr/Ow8ux8smiYi7Seyp1Gh0r/XZhnteKd+pR8Y
S/b5734qAIy+PR3WDbw/6mecxNrzcbajaL0jIAzIWtIgYXH+CS5fLEXzprtBEfrt
/5I1vju6csSk1mUavAI5ri3CwMFVM/24rtThMecSqENatyCTvC1ag/nr2LNwNiri
wd6SyoVyoCdjW8YFrekdn9CWciCWO0D5+mHRuaobAUzuLCWjNNu6wx1hM1Goc4cu
Qg5sR8KsvLIIC5N7vygzxl2FbofCuKG1JLczACVjaCCV864yh4eF6xgMLGrWGrGr
t/8kZx02I7UNnwfelgL9/WOIvu9OpCvio9apsalaZnoMMsHpNUoOge2bRCPyklFO
a+fv00b/774K7q1rJV7mqUDtlwf2ni6srnuNC/fsintskOKiv0bJW128urc9OV3O
ioyp/XE8a6T/YhFsYH17MpVKEApc+1BeGHxBex+ihRm4e94Rf0M/3DLkI71mrWhj
YO1hcH/QG5SzT5ZCJfP0qW5ewKRWEVWhJohkkQ/HJB6k2MW1VPdwYCKrw+EtwZXC
L5voKT1KfR8AURtZKNNAi4EJzaTwNxZpiP8qAKDXp04DnhYAhofO/TNbjZVitRc3
R51RbnwYbpPgLYe3oQsbWJnNhSyPEGx9lwmcVqHWuMOcFbTN9YqG8QNnqRhJLFEe
q8ohJe/IGlXiPUBFzA5R2lOdRBtQf+4OAEgBqRvXRbab4e+y5AofxjDtzm22MJi7
PbdVM9ltrZ1D8U1b3vhcCgtEdiH/3/KxOOq3DTgWpyguv3HcdDaBJ57UNvR77H2Z
0F2mqaL7ighHchVAmyY8Na72J/JsJHtIYZBL2GEy/jPSGWpSV2Vl2gZRaCPIr5x4
4mid8wpa+49d5dSqXsJylrgv2ErM+BgClPalAO4uHaiHUj34zOD1qQOgeZClx3dX
qOTWExJZmohgUgwlpuVL8uPUHKtWMoq93DPNN3I4CTgiqyV5/ZwORSI5B5tklgYY
dFueVSUbyy3+Xd3KbJwxyn4VQdgBkY34GDfgWNfJovkhLRxKnkjcOvpj03jpxLee
pxh/SbZSmslLZqhQEpXu2GGNb6bb1jhYJH2dKyRKDyjUoo0Hc76+/4dkehlWOmxC
+FhKjOrrT8kGN3CnJrlocRGqLEX0fB/kqB0aFlmA7OW/2lFrnYov10c3PCHa9HoZ
Drm66hQShnBDaFNcqW78le0ixkAz3y3cmAdvasjZcb1mJFxojxhPjuq6s6yStXzB
jFVyX9NJPZz6pEZALQBaNz8aXDi2QyFWTY6YV0hiPOyqD1U/rUJAaRUFP4n4L7YH
jiXIWZ+dOqIhnPy2QPEnOPvZA9iqFWhnE07xXWN9D7o3jM9268qzYQzqOssL5MC3
V+S4s2F9vU6PidUkmVNFVhlErqoLD6tzGbS9Egm8BNKmOG6QV0AgU7ZLZZ+OQgyz
6Vbrrsw+g9W/NPXWX52KNmjmhHk8ZeckR4HO8L6URQx62MFnt/fRYbfao+EpWoZj
8EOG0uPNcdQVhrA0YC3f78czFtrMbmcu9CkTZxZ4eIAYC/T5FhLO54Cz1fShCXiN
fSEd29tUoLijp60jdg2KtOfrVkQqANqk668y9mAhBQ5b4MMDn5Z4buJ/cAcCt/La
dKlglCnpl9Xa6UzqH5uJQQF0vQiungQk9iCTckR2IytuId2KFBzK1G4Q7T/wLAue
Ukby0kArs55dC9v1lYQIN19Y+RvMT+q+WCuELZusaqqNqMO5HSLffZOceueJO4hi
Q5Q6D8kURpRIy/7s30hK1UhoDB51Rc+LUaH3FLovxA9/s7J3l+6J4Tv2o6Cyi4xR
bP2QeiprIMK/Lur1x8vetWgDOGtC7c7WUuxhineqRgg/JcC2iiNSK39SeB7yiGW5
f0q5DvqK3SsYxod25v3e4QPhPFi0N/SM+XuBVwJCREEOLhsWMOGC1KcDURwLZyC0
osW3to2zLa1UtIYBUfKeiYIzcy8ZwntzKYTojPROoOtnTPoBD5ujJXVEAJBqxqyB
7RfVr6INKAjjPPh64hGNbkAz+TvTXs5cc7ygcFTOHDu1a1JvZRBFjakGqda9eUXk
EJOTVSwN28gMG9rcZ00E08zbA2prpgSnCXF3uxQp1IFIxuAdGvEVKpDblFVxBurn
LyroFWPLzj1SvhTZIFoGwlBem1LbZu2JAOePw0dlPqWokTXUHldDx5bCf6RqV+7x
agAnLN73U9wH71cNjj1HAJyqhUOEWT6DxFg3fPT+AXNxIgluh9JINcOMkLKXfBG8
uWqh+1xtrg4+jn7slATl9IY6H7yTuApcQTwPRjOZhtSBFvfy2TgIH5kOAChOLnh0
ORd0Va2R+cUp/RFQomVbeyMu3T+Cq2ebPTOlAe5kwzlJ9jtjAHYYXsDdqopT/Twe
FJuzHFGwbPIU7AwtjOcTMtO/lp+rnKWeBZKiygLk/ofnjPcBtozvKwO5KaQecf3U
f+XlsEkgDJPqz0Kqz7GchxPDkJ5D+ad2V+0KgseN3+qXlnG+huOZRhqQtufaH2Of
J6Orq6PeETQMd6rQ+A0vSWoBkIwL8imTBLxUaVzBNKJ5xLMmMh3EA4cmVfD+Qrcf
EDLQO4GzSW4HpQ+PNeVHn8g8mGI6+pslQAebxhx1bEIHm1Zu2LY6ao2hAltPhF/g
YCOg78vHKVUgXN5KhW5nCLI+e7Z0pq5xzG/mAxi3busImY9wquO7hNKEpQPaGIgz
81tpssiZUEvahUPkN43Z4bjPOz39vqjwtyQLj0UXWWOsd4ZsRwWlO/39VMyPIwEF
LkJAva+AIOZksWZgVLm1+GSGZmgIiK0d4I6JHmMJcgiA6X+VJuD4ZN+LyzpLt+MQ
qh6njoixB2GiwvA7vp2m4mmbmsgecjBtu2g5yzwK8vJG7YjQyXLGYejcwDjU7fwL
YPZ8dMv+7GhORMxfHKKI3BhfPyCSrIGkcp07EqsoIF/VcjZBrCAjAJsjCuu3WP+R
CfL47Objmo0srShh2Bnp5mROjSAFtuhbWvQLtyLg8gREiYxN3mfK8MAoMVw8PDCT
CJ9gzCnSMqsGygkhNCRScijydvg9sBf+izxYOQF+YmJrQYT7hH0bOy4AEB8IlQbP
8/18HA5yPm9ZIL3u/iVrKzsy3+5dlsacIn/UHxS9WkKrN24mec3e9f82QI2ni6UE
KQymWXm513cux/FkK5An2jdf6BElim5KNbYOFL7s+ExmbXHTGMyCOjvc6LBmXDI4
eyH99LMFmHoSneCHfN0FU8mqDN3cpkgZaqcQU4g4AZS/mLnhiOXWqR9b5usQrA2l
AdvcTj1cPwPONmjNRgTlQbDafTgOFG7GsmHFnRcYcvfdP6k5NR9BXHDtwoTLPzf9
y224HNdhENBAavxLllz1aDiaUZKeD5yRWVy/mayI1Oyzw1jc+If8uGcGNpjDx6GO
XhXBGBthesnx4HcJJG0nkrIzQFuCTAwdT34zdGWsQhkQ4iz74XVCr0Db/1zn5sYR
fSvbNt4Tq41P6K+gV0wIJe8IRQbXPExRwA54spCtS0wdMEsNZwdyhVvRAoJpCu+p
AUlob3Pwy6ffl5DwUi4nuGIexSjWybIcgMpRg0QHWRloslamN1yDjj/smeeeNC7x
Y/RM96rYsM9Rk7Mb8NLJZ5mxBIbS3g1DbHMcscsOQ2JAO642JO5FMykZwfMtbqaJ
O0rKzmCzdfYFFzYKsCGp6uqoU22IJbDdGE6F6fEDa3ZtGaLDozG0SrPhRakOkh11
V5May3inpp4i2oJLa+iLo6toEIVJXcZ9pD1in7gK+FLzlTmvW415fzfyLRkwANCn
P4pb4oA3FppjPUp8Hro5J+rM+CAuYEsRzqTis8CsrCWj9WmqSeCQ+8siK2tlt2NV
hdLWIY+ekbYh5vdDlg3+mrCblWjGQWwije5M1ChtUjjXAGasFv9iHLjj25cKhyO5
pGaS6Okv4rX08G0AXSWcfe4uj4+k91pcJi8/lc/9ePv2zwsG1Htd4oerFBrYxOSO
CVyahi+wb8exZ9yGgTphv2RGyJVmbeVeQZKCwHOXCn2UyQ0v0caKawElW6NvxsFA
fysN5fznbEL0vl09nrdUOkRJpOzAvDg7oXUD+N/8moQNV9qazL9LCMN6a5WvNqV/
0jTdmyjhanfejYh5BofI23BCFS42624LAxRbgsuVaaGLoW/xk9NqJQOT4Q69gBz7
DhWrgZKVIE2/Newzqbh3lChz9tYlza9GTBMzrGtrd08NFWfTD4AKhHoNoVjObnSA
nqiww9A/N+OEiv9nA2DaWiAbF6OLO2qAM92sshzX+0Jzb6imtKWEads7M98lTe09
dczFhB2BXvY+Q80l2WMaLXwZXjFDbsF2cD3jw5Zs30dVpo6vG2SmMqjzK+1qbZXV
r53lRovFlPvtv02cLvwEyoIq4YiJnbTDCAV/jxKdDcqjg/Y7sSCGJ2y++h5itEJP
AM925eEH2XshV0MhkvxJD77TebgjTU1dOfmSIMatx1kn/zLcQUEhCYs8eddWgB3H
ypjtavIXlaR8U9LNmppDySmIiKsD+9hurD7Rq36uxU7ciB4MSExjP9/GOr0KFgY5
cSd+RdKdRwR89W5bDxLSX/Xy1b+AZJQodhWLOdQNJtJZamoresCEaBcistOY45TG
JM1C91i6WhbjlWXncnKKU4uCxn1EG35JbKlL8XJIBuoewDzKKDBzBcBhcLd74WIg
9LHvZRxZx94eFWcRtS9opsckycG1sZjukUG3Xa7XrqRAiQvmE29/sU2IigZ6q8u4
z8wYuMQHNN9u++X1Q9oNjZ7dUnE0OHYVmvbx/XVgjuX8I5sSvJ8oZOPea7ja0Iwi
dXJmH6UzFFnpJ4A9tae7VehShH0laFnAzhqNA9HGYT6XOGIcydjMqqnyA7JJnmxR
hhZRVSm6X/AEyRTcfRqO3AEjcPVFLx22+YRQFrxocR3sVPVuT6pJxrDgpJ4Pafjj
Cen9oxub2RDDv7ku4POnVU+9Q18nVkJ50CfMBnkQJjP2Lz/FuQszD85+bxyUvMam
WDFY2wEy1vX9CFDkNwD4GKfx78S7ctO7G7GoIA+mxvifjjihk3V+OSkQQCMnYsDs
bXkIQW9BlyiVCmDdkd9aEE/o6IVFqd4ObEFRRg5MSVntPYAmYIgigVxc+VH3nse9
0/hJnKSegdNrtDqTHUfwB4sM4ugbMQ/5umSTyhHkRKPJemljxwkWIg0zzqy8O/K9
P4AQPBWUcOQ9yDFBPUWozlbcGlRqKrWLhBNNiT1slJw9aHKbzltX7buTCINaq9fF
bh/Gpmt/lLnju0UiXLMRwtbY0VG8L3Aqzj7rmuJujJh5QxKa8ccgEZ/y6T8Jy3vb
WvhY1dYO8Fj7ElOoQQl2IaU80byiD0cSexYmTu2lJcio3DHECzFHqvq5IbXtZqDj
CbUgqAigFjBE+qmWrJ/lQGCYv/m3NZCveLJknP5u9uxjAt8d/3sUs4isPiHi8Yhz
A8nYmF4DIbELic7F0qPhwGj/c7IxrR9AjuT7Rx78F4S0vt09A/fPDSWk96sYf5VW
MLLPVrEnDsYx2bIsSpUDFNE4MeCOKFpIcwUGc75teU5brtxixDlEwwJN1SbQaFOg
wUIJ0M/WAwZqZjV5SktlRHO+T3Mur7gVL4ubqomraWUhUIM1chY4jTwGYesgTSfK
iCs3VUsUQZCA4angnpURYMwC772+JZoTtBAeC3GaXeFfzcaxPn3kt/R4lQ6FEkWs
7I3HqE/QyMrZbjOHQAvEwXAk9LwiBZgT8EkuXvY9d9qGyqwPlxjAGe3qbk4bDFGM
WIhBKn2VlvQKnAV4crJNQmfwsXZPaTKsB30id4bbvX8pfZUz0IkCnnWq952h3qug
PkwGu0QrKM3sId9lHuFy1T28vI6Dskv46+zWtZZaZAkeTuDAfAv3ZEZVAbqAKJ6W
JXaA7Ea16HuS6fNraSFQCU6io9KEAHqq0jy0XDOrFSeaLUmAljz8BdRE7ur7Y4Mf
Afa5/Ll2zk1/L60dJHdzODetXANxl94wIsWnWs/wK4I19pm2QTNUMOnIDIpnWwRo
BvzVXBC2JwTiwy7mPEmx+af1aeUtQeliayi1BLXq15o9Efo/Qcy40B1bWyOR36cg
UM6JnqhTD3mOW4LYUKlOsXK44rMpf04/XsAN2oF71+ZdUQVTMmDwcsyVEy0UG3NZ
/BNZC5SRTP/uVM722oH5zZFHEjxlEyKsn1baBQw3k2+lwrPRc/bH2XAWFJ8TlMwA
NBnfgmcNcx9SK0m+PD4p5SxcEIfNXsNttwAJR/+4uHqZzXuCMeU5SFe1jpWfecV9
3W9qVUWJdXSyCX1sF7w5zGDuughCEzJ0y8ZPbfHWG8rqkGlEbOlrnhY158DfpAsh
wAxrNbB60EU3VLg6TKIuuFSCppztE4fD1Ky3pdhrvCgBpwomaLnmoBM6S7BnIYyW
+temqBOTTuVqgZ62P8DaEcJnPtRuJCx3PvLSP5mqUa5X5XQzTSl+/bhOYuBT7XmO
PYYDVQgiESIuWxYS8mWyxCdleJtSakZWsmyKyi/vnHTH+2hQu02iZAin9NbjjxaG
WXbqibqrq2mJDMAYXlySKkNFtiadMBSj4yhOl6oT0lvP/9kngvQ89rwklw5nh7qO
gvfNi2+aeqDtvwaps9b7R5NjsANL+scdZBwNXDgp5+vE/SLEfPPyKJK2YNO5HoJg
Q0GvBFAGCrKZFms48Mh7lJchrjT7xIZ4b4MJwgbydvqupyJ70J8K5h6dI4c0hfPX
O6rTIf6sUd0X63/WZ5F5nVCvImR98qaN/nUE7o0Gm3ezktUaBDCS1lh46CiBgY4F
nktqGsMEogj2nxN5rbDscCgUhCKdh84oYkzkcMvgbhsblaW9DzpOP3TiCt20yGD9
yDqHtUpz8WDLNWhw8tHV8mG1jQbHpWfyLwPWhHsL86WIloZip2JQBzdhRYgQhtyn
huQu+zLWwjXY0IQljemsZFvT4R+4atDPDUr9+bU/XxQLZTlJFLIpq/GYNE5Z5+gr
hTki4sHlQi7q7+VglYayj7OL5OnX78FBqhrVoJH/d8/K285gT2Ti+2Bt+S8PUoEn
+oCj5JdJYD3F6MguzM50yncAU3gqZGuS5neED9i49ihGiu8Ioi+wC4XvIZdfTUKD
Ki9bcNNQeefSsy1E4EHHs+ac3WRpGZqn9IUOid4bsadJVJKnObBuuB4hGFHLVXpO
jY4UfEOOb/me95EjIFUlvuxCBYmOYnhpmK9RFf06HzYk+4mdivHaLaxUeLH+W6G3
i90oACMs1wWk/V0zm8KtazUD+aYpmcBU2ZvJw8fncSBEOfzDWkDESzI2RaoI1du3
2w2scLFn94l3/rHHyC6V+n/pvqEl3tkzpHJH59KN8vYv2CjU5lbMAl018Y5Bv0qV
J2yMuTs466sWFsV3fiTxe3v9KjorqrN6yi5X+xK34Z90Lhgr3iXeuginptv8vuBE
va6Qz+7wiocNlOqniN+dEi3BYmF3Ksy5ynR4viYXarT8oPQd1CGjt8Skdx1Q1qKv
y4xF5P1rhp+t33dOxxguGapEFRmo8WFraKVAldUI+xK4DcB4Sh1fssjBRqoDzQ9D
2/g6xrDUn4CjpXHyYqamZc59zZ8O9TUo4lDZuR+eCoACYKvY9rQqBLioirgnhecn
Z8azvQ0G7ZqSXtDwJpJOVnB7TujDMz4wcccHhK3pRP+2QW5qs956qr3SXwR+KKP7
T2dI3AiVtm7aEG1Gpm+pRND6mqjBW/jCAxdH1JIfd54OH6jgekiftFgGfqLOq6hT
0xdDI2GAfnD83Ed0oFpkTwfJMvGSIa2Iwq1JkJdO8iu+3GK18dIaqsvt12LCAE4b
CC1eMx6EI/lS8s4bIiWvNfFah193qykb0k7sHL7WjUYlwWG4i3KvrmIRZ2cAQAor
I1dvLaL8jbZFf8MfTio9ybAEmhIq4ZKx+54bTMI+SMru3kCaAMD+VicIZhgp6pjA
7qqngZnzFPbr8siPxJyGwdZp48P2cVfeC7t/0QhwV4es47pxSOwfyLvAFYDApiw8
dtMY4eZ6y6tltESSFKx0fdIwHBKsgVh8Qe9nkWri6LiGTj1MWnd1G0j3VXlVTB2C
ejNFThFp8CK5SMo9XarrL1fpHb0IAJfwA25jgvb0018FMitfydrD+cc9XGdm3lwQ
aWkqvgHmA8QhJFkvCwn3/pGbhljSpTx5W3aiQO+zUkfr3y55ZzN70Amni4bsoGPQ
HXgAw0RlQLjMb0YHrXvAZWhTzBgl2tmXIllrEtYVapqsP6Tyyip/pKuax8LrY1PU
3o5xgJnrCSP7HmJna7JBka+ZwY/+suZMHsteIaUamRZl0EewH2t3gYwYt1GmVLvr
RqEw59sUVGDuHPHLPKd8jB0pgAwrmVftsjtvW2dTAI9rqeqGZmGVNkTM99GCqyWI
JxW6ICIwGfQF0taHUEC9O13MYKFyriRUM+7MCnC8NilKMKxWReZbIsONaaj3x22b
M9b3+zQuLyCdX+6CnLrunlhArigtARlwkKUMgZSGMwG47MYVZH9JBB93KsswhfTR
IibMtZI3cjUpXoR6Qym+LTSKqiVTjEhAAZgDRlZ/TmIzcKFai5GQdURJf3zuSY9R
YfzkUKcBqsjKfDcsWy7B7XSbzOeBzxWBnfgjXk+4YrqdtExz8L/2xoEN/+4VlnlV
vnxXk1LtzpVVSTh7HxcOiG/93kqPsS9ge8j3BS4vfqRDk1mNRXiSjR7iBwWj60WI
8olfXB119OzMYeqz99lnA+I9cxCyE8yyGtk2csVWjUL5A823MZiwieHLSQ32qNyE
GBZjS8/j6kb8Zs8gSL3CcV/Y4tIM8rXgsYz0ehk2jL83lcZgA2qvGEnVCSzeDhgU
zp4lISiC3eMqsN8i46q50Pu5yF5ILh1POMDi7aycH3vBgkmpLRDCs5kcvvyIuZwa
IFmLMWobOLnDLIW/Lv9gMuOh8yqUPqUHNYoBoNcFM8lQYspEJhXoCk5ZQqwxC6I4
2Lxl99XP1ObTrXQPELBopcYlN8Zehyps7xl2QBJxY5F3S0BnrsAtnM3OzqZcgM2X
WesNyC6DOAssqFUC9+Sm2B88Beteu+WGKgT33UM32NabtsLtR6WRO8vcNJ3Yz93B
aTQsuIer0Atw6vYqydUQGLuVmE/ZJ8DS/4o9dwvBpYEPip67DJsRgYvol1RGcNjE
q1iRJR2TXqUTA5hzGyOIAGL1mdqAxwdhGwGijqlBXmgwXDdeWvijbcR5U7rVT5su
yFHAraN/3cpLNDTex6R8bRs/yo50GSLII7JiHVDZGbSAvSq5TfCkPpG11pkpweUI
MjmEnK8dDxTxYHmXEMTQd6YhHRN4kZ495X3YWxOKNgiTilD1aZFt8l29KFIc9rKd
cmLe9zs+QqiIT7HIriQBVi5D7nCXFUX6F1AqXi4Duh489H48j2JzgtyNBffQlOC9
Iqd2Hn1WRx9lh/+iEQ8/PU5STVVrHAu/i0FTa3a50MEKbUkkyfO0SNljpi47IxOO
XyB0lVv5yTXsYZFNSesups+1bmbibhCfepxq8widcGqZRyhfgf31N/9a2uWFk36c
zMm46iylyXx1ixgSjC9aGHWmZLfgWwEMAWyxR27YMDjLflxWDB//9k7BMmR9Jd1t
BFmgJLGoantX014HH4BkeoumXG19DeBUhPTydZ5ZlGFLKV5EKUAp3PszigO0OS4f
ymsqFBQ4NYne0MvBjj3ggNqGPdDQZNRHqBEh7QDZFABeUqTKRiFAF+ndbTvIvX4/
jG3L/0MqCF/Sk1JkJJKSUhoDiD+ZL4lffU2fyJP+pR0BdOdyXFUaukRYaKIYMTwt
ZruFxFaGBV2NXNTyL/YyVB6mZC780Rv5ePaTXHA6ERNVbhaZkrrvEKC0V3r1nb51
doypZoHkKc5SD7LdLHoItGs8R/w/pm8PsU24xXbnkRVyrpPDiwuRd4e/knilF7OX
cBTyspmWAaeQuVs+Dyshpu1MK3QWzhV18yoqUF1kMeUi+1xxThIlEi8V9hQWDf07
h6LFJSy6DRs/6FU+Ts1GtVPbceNXA93wnC95j53sxqG7Wxl7vHzuAY8aouYx24CO
BoI1BclA3iO+iwsKoR4CKfD172rCpUWeXAO+zV2FTl81PAHcmUHagjTboMu/LDX5
sG/94RG9hpnuY6OEfg2krKYPon4nMMiAOTIQNsidasUk8D9bFJfaBK3N8iB/etHw
WOVWe52yFWZwU+Ex0gO9Uvi7sSF+sX17cobcuYAoTMjBJxemJHl2mY5Vb2V2jbZv
Pn4vvcR20o4l8NqH8tuP2fYP9/ufBK8LMA9HUONVgAYnJCKZKcCu+1imP9QBmNVU
PK1RI+2XD6TBnD9DqqP+PAatmYTfalTe854fU1fOD/+gbp4k6NkZ7+iSsnRZb/Ei
6OADd6sh0YlbRJuWaXe2P3wP4sfHHNQIQ/pGO6KkFD4o+9ICFzDzGLjqGhsTUz7e
rLIh4uwAtn4PIhTDryWynCAZM0b45Okljx7So0/HlLJcb3A/ZklGYReqDzAeZySq
/X0zmxK1dFL9GFexwS1kgDS9seiQlhcVCc5ID0qRi+JgsrSZJutdSxWJmoMYBkDi
dvNJ0VkGWFdNs4dai4YXePCGRXqgkA02ev26Qn6axeBfE8LKyaThxb/mD/CpAp/b
HS+efwk0A/Z83Q6DGwrLukpAx6pCOWjT3D68qWPq3nsdy6sqyDI8XCdKHHZDFnt8
xe08BUNFNeYhWY87ig+ytLTtxRl+8Kk0YHlQCXzS0MpZs7tMaExxqMJmNhSMcA83
NEmZhSMS9gEM06nV9w5riCfsj5ke/SQwlAWTMo5fyc94TJ73bs7NzGHBtrOPaTfg
daigO2bCfCr/59w0LjlEFiBmOyE+xzbNXodVMYcjxNe43J9gjceOH02K9H5/BXyU
vczOx9xDcfAlGLrI+1+YO8p7DisaHdnEAoKz2sEffL3QAC8zSwNv3WUwFXhXoQDp
pY4q6L9+GB9niVDsNAsw48zhQhGxijzvyixlhXiomPHfxd0NaP80vAyhB0xki9Cx
0dScM9h/Tjr6nlOIRujYZjO99dqD7WHKV7nCVRg621LNC2mCrUXg0X0dwmAvBgTb
wh1YsmR16W3SbLMDc8ZcyP5ZnjeN5gQQkkbSc04WAwXOnyBorFpYwxbFsa7rFlaf
vLQl8o/NzjOcvXIuypMsoRDonNGy29JjdY1ar6RRsBdveNHv93DRYASdu0Z0pYXY
LobbI8EbAg922O9Y6DQi5oa4jEJc/Tu747CB/cdjyizB8Dnv0r2wLcXMq277aXoh
K62/TyNHX+R6W0ifY5HUOtG4Cilc9CcHYJTHCVXQer0KZHUb84rroBH0k2Js5j1l
4i17kNkEZvn2M3e/xZ9Kb9gIPhZHRERE30T3/+ravlCDTmwvM3P9eFDOA843y/fm
ZDwh6NheoleVjSQgWRlbVGvv3/PvNlTUsmWIPZcrDYoMtw3CKV2gYF0SbzMowp2f
BTgn26rIHi07Bu/QKjUlnoszIT173147HGHFaLAeOShfTjuWdlW6TF1hgyLUHdp4
9ZbZqMNe+Lh7VIP6+rlZwA0Cw0gxw+NcEfBQh60y9Jo+o+B8+52v4/0U/6yLx9NF
yKlA9hXdNkRPxUV6QC/gXgW4nIjuauGEcxmB7pmUWlQWnNw7NoI8JrDyBVq8OOra
c519RyVh/n8nnPRoywGggP7q/PtqJpvw9GWVmqOa5mCzr1QOZR83FLn4ngGJY/11
sT6xBoLl+9fvNxTJB0QlT5VhS5cLoNwj2SQjUT20FVOAqjrh7brWpku/DegfIW99
F7mXIx4ZPk2pHkB9iw2t9Tprwn4dDaWdQASMcbB1W2iIF33nd+A1xkEm7WRDW4sM
79JlpPIJqgYWd6QsquXLbcPeCYv/k+RgrtzvQnwxVC0NGr9WqoGDjcmR7GQP2mzl
8yKwUWxkaX61PCo15rL/2NCcrsRz1PDRL+vfnFw66ix+Hvnt4PuWZuuguEWJJaQ+
Q4B0obBd9/jTVMXJyfxI7TbSGyYLQqgUJsh2j1kQhBGDgFJbrIuS/fCtLK5TSUET
LSaLSgDcOkYo0sNW5QTBJPUCbrENJsoMCpKsxTQuVBgyE+mEUHO5jbkRhwdLQ9vr
Bw4T9YVeqzUeJao8hjr68n/6nq66HsBk7J+Ch6Evz3WlMQFlhYcx4530XiT7mdrF
W6DfC2taS2xSVqfMnIGtlfKWPxNf7U9kRb4STeiL5wuld55/sQlAr8nLCxO6NGBd
W6FSfFQb50kFOsgO0rSO1ECOlewlFJyxZoWjH+06LbQ0JlzzZp1jB/U9EdSLsojM
kGmNXzwvQ6yS+yVOHOchHpbW0NdDmoywKPeRpk6k6oyz3+S/TUUHjzVvCoxto56U
JbkuBvB2PRljLaEoxubuceysWsUyqayAsgXBlGR3hromkbRDGw3i4FrXOWkT4ygX
a+ZBRruEy7BJk1RgX+P9uzZ5ZPgpKSyiHlm9YVHir5usBqRM2h9RIukQY4L4r4q5
eC6pPRYC07OWxj3FuO4gxZwE3soryR9vtG6RF8/dOF8mV69M2N1N/MN8+uruz6yx
rZLH0GYQUzzLRXAxQHVN5rlwoG9Ns9SlKzBhZe6+ruO8UziUGu/lSDUlOF8GaPUW
NfiaptB8885ISImgzf7ybcXEYYIsCDdGx07uOTDn3ZAUe8v928YR2HJrxg1SB9+j
sP5ZZNitALB1jT+IOGiZfn5IdbX6zp7uqt7fZugHyfLWW+YiLhw38i7mlyfOE3Om
GFzR6qIoLB1skzbqo9Z03cuTkpfjlDfoWKM9Xn29VLhCk/YHCPNLvE/w9t6BRWVI
Lk9/6XLb62ryktfPbC+9VW2NdSIq5NCPcjf4y1LtS+uLKugb9WbXq1oLXsNQj9lD
DWHTkET90dV/bEuji7LiVmzIFDou6vUkimPhUgye7MdQoGmUu0qkVSEuWuLI+NiI
L9OrmGhQSnSS+S6jHVCUM115wJssr3QbdHKlZG/wyY1t5drJP7r0PjhBM15H9CkR
zpp00X83RcubgXgm5hMnb/DM3aM98tK1tVRlxtdanfnzZjjm1P39yLb9r+zcIESD
0HGQLOUfFcqheSx/QRq3vbnZ/ipKnTq2QI0nLXpyeDhQYY5hSIk0fG8PUuaMkawx
wWDV3wayT7Z7ywLmFelQ5YhF30d59MVhi7rPnKOVAliMVstj9M7lAfvphJgJSlX5
HfrDe6oFULS2XH2/mA4wENSWgz15AtaIoKe85GrH8G5CW3IAWw9IdJx9/50ZnwQZ
7ve29RSmh05B4aPw0d/w5y8Vq/HdRMBx213oiEhxqFPPF/p4HuN4CbEb+hQL4A0E
Igkdvn47TFbt8XM5T2xYIKyqXh73terJ+jb8SGk6qSyR7pDtry5uqwF72L93BMOz
C/mDktXXWuuqQC/EW4so+golaG68htXGz61eyHUYQ67InmtNrb/Vd1V/Py1psReL
oxh5GxtgxImFhQongSZVojicOsQu+hL9u3o6tPF8lNOWObE0ALI9s07dhJdBub76
Ptjb+0VCBwC6W6EhcR7u3gTReRJkEM0mJd4SWw0ePKdNXa1rXgCpjJTx7tMBV/Kq
P5G/mKPyZUg56izG37Z0g2oNFozIu1aYIji80qBjLKPIH6lwGiWbLrpAv3pvpy1f
9AekKNRVyfYkeULTdT8dYFUYKU+OUTEzQtOASHoB/Ce6e3U3T5DKPXBnejqHa8Ya
PSo4zDaeMi/+PUUqXVPgbE3lQ7J1vkojaRiV9yYSGeZHu3J5bvRojwQdpbdlUuS3
fAm/ZAbN8sxqS/dnZw0UMda9MykjRy+ulJGcdwYx12Em+cyMvmcAriQFxr7njrQv
Ga4+67348lFjjV25gN126F179mxHD2u8fZRxPFRk3n9cY2RkCAu/KlFkYbWIQU40
6i5Xt/kNPHUvqg/fhmu8xOvRkVB0yP6t+E5WnIAlL+W1Q8X++gyUs7Icp3CFl0qk
NULrZ4sIYne3eyyQUQ+znWhpBeVijdUNNkeTbBxCgf03VnUg9hMcmnWMukmL3Ztn
noT40/gf84X/uduWYkSJD6AOrJ2cA9YpzP6uLTq5Cv3sIrt9Sxype5HLUgvH2qdl
h0f1aSnXYA6OPE8eoA6tT37UaAxp+1o7ZbjA4qTbAGT4zNIFYWf8IpfhqMwZt7U+
guliJSsjuqHHsyXGhhjKii0ZsiPizBkym+GGcd4Fn53PoD6YRidF70xd/x/dvx3J
un3HsLkHPHV55ECzkOCFFRhjY/yqbFAoTGcrXQyqFwqcBFMGIyQ5QuNx3BO/jrsG
7hTBEOkdcfkdFcKKljmBymvWfm9kiYu04gwgPBfIBxYU8LzmiQdNyFaCev/OJnza
Q9zYdDjUPYJE8c2jfSowtTsWp2poGbqcI6d53E50OlI5bzR9/1pg27+AakdOwXSK
Mel+anqGByOdrgCBN9gHjxeF35JFgL1hMYWxieV77/Rz1qRt4d22nHbP/TS9htcY
C3dTyYEJhG2o3sc5cZadQGy42mjQE9nba9k0AOkFUIHa1qb+FW/L1ce0hiCLOVyB
dnx/nk87wr+lVV6H/JHfDH+9MGVjVkbD/LcPVkeGJtullrMPugfYxaoeefNte3zf
Zq652nPFzDyJhrU01rs/PN4DI5xEUG7ilnLIsqU4l+nR++Afolj1z1KJCjzcHK7L
DE4CP5d4APNmiEPYzfmTSu6Ye7DNpR4ZHiO3yzu4GmRl6ZTutATFy+Weq7tKwh9H
3a7kldKB5BPKNMk4ElT/w4Iu4okbOvzVGWnAaBgBOGEBqEUF/36kd6Se9r7Gvg4S
3l3UqtBqtj37upoz7tTlkJNQHyniBEOl/ZdGPfQi09ihElTFO6gwPTC5DyFVfcSD
f1M2epm7L2/GIC9jQgHQPX/KgCwqhwNsCC3jw8B9x5S23p+tMMpRcM28FTFI/oew
CcSYsrY127rRrz1P1ak+o+z17Y/EiB11IRjj7uNKwfIJ3m1IDiNkulcpH/FKa3vu
P75KlPCerpRUznNS8MWfKhUV1XFG19mZ7a819FiVJ4uyC3jKOURk0Na6eiHzzpc5
Yt5oisy3WoXNtjhOEnh5a0E5HJ/evk2kVFRDsK+7U4kM/bVOR8btS0CrzsMVdXtu
/XT6s57oQIrAJnchQA6kiB4Hdag71+sAI51jKgdk1vkC1Ep3jW3R4Fps8MDu7sBp
cFYnKjv6AGk8axGUkpZRpWksghULkOuyxa01xndlhOUWG591QB6u3d74y0WF7Sa9
9ivtzeRMKzKfa7RM8YNie9F0Rd1Q0Zb5tAy230E3GjH0D+F/qQbRn08x82PLFkkB
64wsTAiinpCeBI98sPT77uxHJKy/422TB0A8WtNg+uxHJSUjFLnS2hcjXyRVonWJ
E1TXg5pF99nAk9cTDU8OZJY/L/ZVh7ksH9mGmlVqI27mp7tdeFGmYrav2bKlUVoj
ZqGMPK5sCmg+V/nzIDs3szHmKIz0VHEuJ0aQzN8nk7jtHpg/Urr+vngcoEKOke0X
5q03f31APzgwOADJJ8Q9Y8y4CDxQh7h+Bpfzn2Aw5AyQZBB/PR3lhSCAamRTKDHu
XFXJy0kRsu5CWLveu9191SKZOFNzCsllwixO1qRHSv+mR0vAP/k8SDR+D54EQ/So
234JTL7t+rm2YO3CsydDUmYQsfXvgT4ntPWNJMQnbgPPoFM62wrIzSB+LG5CexiI
rITSjmucNOMT/1bHORjOajzzpHQAEowTR/nUS+QqIwv13Fq/66wYkTIXpu35JLbu
7PL2tUTwtDY0KHsvj+8W1+fDcsViITGQ7q7B41AE6zAsqYEcIi/N823gBw7SnhUj
9l8eEssShH4eZ25MkH4YqU4ZfGFgD3XaOd+MxzSDwH6fSQuABtn4PaxYn8334u0x
gDIVTcnE8TYwhyoHS1ACQO4ogaf1MTmtnZp9fAw/Y61LCrpONvQM+6Zoj/QG7doN
FASPXuBZSez+A97SWiNfaq43hV4Fxni+bRj7EtlvQl8ZUvu1DkRjydShckKzqkqU
DgxRuEt7pUbV3XcYYrguSEWQyd1BuJW5PQ47lA86LNvecnq3NRvWPPjBGyingpeo
f9cM5e8Gg6ZsTryy6CJWnR7QreVQMy4oB4/U4TYmL1/aUgaIv87SkLXz/P6Ale7S
Bt8CDVFuVafzUcETXLdwnei2yyhIqR0rUG2jY+mskY0pinc58HfNCVFGlcHURivy
ijYqozQLyeaZ925b4amefsCSJJHlhWO8NB0qnbzXDOEsNdHOiv12JswUcG9JDEFG
IQTFNa8cHP1mM9+DFxrcDKPtdgXMTsAHBNKgQ4lGlCd+f7ljiR1euE1TR0esbiuo
Kmn1co7EeEqCMTqsZ4S9p2NsfCqvR4wJo7Gd3tuONBnrlmDTmLjkfMen/qagJ9J3
l+i9B10dyjMLlH0tOmz1mVjjK/1h4kjXz0DRYFT+BQj++N/VSqoy3kcwemZ/4mU/
MdSMkzVkqb799oe3bKyacyP3VzTxA2hbsOgrGG5ot1xGZaIR+2nBY+3LVaus0l4H
smbNWshijrjkwXTvw0SvzeHRYHDTEeC5u5T8cpsgaAy3FZeRcObox2c9NMUR1CH8
MRu3MYzOij56X8joCL6NvjaOrLuMyx2BXsUMYEhVileZh2DeIuLaKatHBoqCYn7P
0t/W/dQIF39tOajPvjTSKQW5DmtZwE0jDkr+++yMzxxjqFoEkGzoc3tXETZkFKo/
GetwwzA28H8t/MZgcoM4iBvug4/i9CPwtt+dnC5WYp8CMVZ4eBNzp201EVX0egYF
1KpdTl8zLelqt3uX3R+Ew9f20V6q9MmeU84VhnQ7uS8OQEmhD0rCYqk7dwAZffvM
T0t2xQnjtfDn3Nc2X1IGgDzsatBLkm6wAQ4dcuCZwjbtji8i2fWCqfplpZcTW6uA
oFgrppDphCfR09zS4q3dT67Ii47A16gVF7HpCOQ7bqsKryL0R08QaqbzQFQLRCCV
TuMfpuXrfVjVMl77sdskc/i9yCUoRQ5/mH2HkEXDyXiKbAbnPKjNvg9Y/W3UPpJY
UgJ/eYMOV1DhDuscCH3L+b3m0QoczemegtIxPdJygb+psQWzyPxMZ/lysKdzimZn
MrocLdgjdRquPz+rXNszFh+4AtoIL2SvFcC7bkEdCoKWSbY10/kM6N0thGMQjW6X
Fxl92FFGzBbtc34Xs4Tyh3aZ4cQeHQqD7ChDI65K4jxjTXFt3eG8MEC4ZSTt7+gf
Bqoiwff+uRYH1rht22ZnrgDRK93j8itYe9hjQefZOBcsQQmY1fnUdAbGoC/Fjivy
1Cvl9Vtt9YKkSRsQPHfiUBQX5lLPPrpRpL0MAtbrX5zyKZEsCJzL/UUFwTWIGo0p
oSYRf4yUM/YoKDZEb0W1d+l1fR934lrFo7nmJsaZRPMrqsbsD414AFNtn62aoLxx
FcGCaPRxpth7FYWRkauZTPSulfks1WZro8aGV8U3hvs9xAAn8eD8/S+V4mWdCUpf
LQEO5XXO1PA/OyjgLk3UL4mZYDpipiqGwbWnz7yGXTlK7r6+0KuoCnw2bW7Op+1R
uwbLkUqyRXsqXMrOPkDnWdwWTimaxQ25Slt1wcZYU7ugUmZstZQjn4JPGcYfV5Z5
plEnSGeLjpb521AKoL1yQcf3BDtqCFbtMJuTtllDzrSaIRnfBUtSwpPUG4qJ6Iym
kJOqj2Kjv+7jEix6jIm7e/X49FQd7S/3KuusOxGHB0+ELvvuWUuvb3n1ZPpcTRNW
9V+WNmG8UMXi4kTBPtpuUp+KcFvsWwj2Lb3BA1yboQAkdf4zpGKbWwjGDA56cW22
bmQpph35OgFTbam3ynF8O+e6Ex+5MI92+N/uCNy6s49ldLHGM677XWcNvtZUlvO8
0CKJql7IqsNh4tHTBXWTRhfuvKLXF8JBL+GFnhu2UM9QchUBXYksWUWCUqOnX8b1
+hwBBdp5giSWjVzFHdP9KVvLOZ8/1m+/bUtfrmFx/GT0RYW5CDZoGFf0PMx48wK3
l3cagdMLBTgz1ZC5YhGMch1YfLPgIE843AWkxarm89ZLM1FsrEaMIUCnqL6CMkj9
iaS4Hrgf/YdoKZUKTi6eFF2vmMTD0SBBJN+C2kKupM1O1YryVZ33TS0HehrIkO00
R++Eo6jOjd2aWFHIAtqnkPlihdABOMNM7HM5LQNhOguISHhTBKzpUk7IDUIsB4E1
2k2Vw3XoGXbfJzY5BhFrV6zPirudd6/w22TKReygOI5cSmEtX2vgT7o1nW9XWFhD
bWadvRDeKNjx/oSJY/nyM9gqmemOD+lHkT7QNDM4N36DwlINL4GLhdqEvCI8HhLP
14mc1nGk7Uof5aTFetkCaB8XQ7mpc86WU7Q7Qv5wJb0hK1FkoKlF/tJaX5EKmxBr
jj7Dt5JwJu3AUKRSqjv6sP1G5s/TynBzLejaMrTOpXK6gOCeeHfBt8j4ok5iCBrY
k52LZRL/aBfa8td5vJzRt/xuZVeKoVL6Nu1qeBVP9js9EzIs4USChYBry0CDcoeU
s+j3uE6NvYE1q/NRxqtQpTS4rv/3fj/2Cwy41b54XiUTYLdTjF8OjF9DrM/DCLsl
y63QUm7dn7EwA+MOUed+JOZ9XK4llf1/cAdjmcKZXBn6O453KjrCZrYop1siym54
0wxDk61m7u9CjUtXfb56p2oJOf76AoVYbbZc7nujjfR5Yn51By9e9Ms86oh1ZQAn
1SGf0bLVDzs0epilKJYUDDU2bdzPGIwuAe4wWQE0/f97mzu2yYLi5nKsm7vHPXJK
5leqns1Tgd/j0MWcS5qw03u1tTijGV3nGu9Bx3Pw2+AKS15uC8GqbKAI0xXaBwT9
AWW5fH3UFVwTO/as2r7HLn2phvCS0nvtG3Ey7Rh12syEw7aFAlR3ipyo/s0lrkyA
ldKCWYRK047w0R2Ao0lM9F5yjfUPqPCtlK5hjY0HMtO4mH7K5JaVsdYzyTtqhRtZ
JGcmCONNF9QHz1AkRz+JbsZ4yyQJoG0CgrJplHwXqrAz2pxQ21qxmoPlKVqHsChU
IXF6QO704jNSXAnwONH1+RE3Li2EeO0fdg/6wG0hllSQOmtSpmeUufC19xH7uKOX
LKnBOmKtZjz4N3Qn1/w/87Mj7qQ23KgQ2XNOGUF7qw1C6Sw3q+dTieOB+Yh4HSft
6WvVfrxovZKEapIKxHydnPOwuvsxmOjJ1Bz7gb/e++zEBxg74pv3IQFWA/XMm2wW
HspwmbKqy7gFG6HlGFDWUcogOjC0bx/D/+GoR4tdUlqwylhC4+TW+cp2En5C4icJ
eqXgnZvBD2ReOORQTdu6OzGi0Cp4i9dVg18twxIU0cARs0aYsq9uc4VJG836SW2O
bNgSqbnCDnB4mpupOq31maiueojIeskS3BngsWERjl3J2GAz46Ofe+cy5CsmO1S4
6v4WVrxkvbMiRHqHWlSJySY5+OXrPw3eVqzNlFigXY08ERkCsUZsklQx1VvbksD/
K4t6sdpGwfKWZb8HekrYtCXlHTvd6TAX3fnJo+zsxG9+DjidoMmGi/1zpTlIFe+v
TxR3ZiNyz44jxNROIE3hvu2G9vfx8jgbldOZhCnVSLN44r8dZiI5/Kj657iG6sJ0
LeZ9vXgb5mfhfH5lc5b5xjpvHaJR+hOTpG6HuA0dIgaq8ne89rO739FaQOY2mHFK
mJ3OeFXp73GmPQtFltnSTsEo6BmV7Zf+1G9amaJzcHYI/oNgXAgKRqdbmGiU0dMi
2N23s7W1SUKPJ1gHaRnl+5LXumB4L3J6SQ0akB9COglSoxEBjR7TqFeg9SwfCnRQ
iMVxkSyUnAuW9tmorbPp318eAUsMT7e5hLAEnpERcGZhHtdGnPUNt13KoZo6DxnF
BrXldiSg51ctocpz7lk57zYx7Nb7BFHS9iw3h+jp8AXAWhfSazXUJZa0K6SKLobu
k/QyFv4GJZLSS/44uSmDnSpGhn+hiCSpksqZQKjyigX43QWS2PFoQtE4nSZIRBvz
UOiXOoXTUc6uA9WWAa02cDs2E4cozYGzxbNjOgslO3KQAbOeQepfZ26hH+8W9GDc
rYFVldUdvsfQtpLaNF+otUueBvBR6dFzFZUfOOzY1o4eDWxKcqXUmDBuo/gluK2T
liz+YLe2ED/hmYwiC7PoDDSrWAQmYsX1ErHdBTqRjjfNgP09QTl0XNN30bmJ/+Dn
jmx7kSObySCGRwhtuSs71EYNh2/alHfzTdRwsFZRCGsZc9Ux3MFV3GFN3ff9CJK1
NHUKoKSMVTOfuuk09yhf/TKzuw3A934Wi1cbAcxsjiBhoTSSYn+HSJbGotmwSFSv
Yg+vwFW5ZDWkFt5E+p4d+MM4ZN6C5ycYZnTws0RtE9AfCFmeE21iYk+nOKnl9ZAN
6F+MELnG3p2JBATHjYW+OYkuVjB1IZc/8BFrhKEP10LiwVjLYiDGI4Ajvg2T8qWm
MVG8hMmxMhD4OE64mhqc0FuOOH/ufV3gCY5rrGDHC+BMsnggPGaZ3SBcHtad1cFL
FIngz43lJZBZ8S3SIZzr5ib3Wxmg7rRcaMbUw5emOnBNZdOF+5mQdkb2gIBh0fn7
AxW6bmsQRpRkT7zGQfniLAtlJ9d4MJXn0BO6RhQVIIVNJ7JRQHoheRs3kLLXe6+S
QuHquUL/Fhhh9Ru0p2gggElumgFWmJrMbYIIPIQP37u5T2JiF1KrN5qMkfRPpJnH
ZINLG8K4ARei0AGIUe9ULckxeDgsT+lVWVyOd1SumHGKB9SnqxsYNhZME0hWLjOB
C4cmZs2clFdOtbGS+K00ICQNACqN7FR0h3fYpckIe+tIiBC2/ZDtYgbUIGwHHxbc
5GqBP2xoCRIlEG2YBeH497LzpmMYJ4JmJyVc6Wqbpbh3a7dfvjsPLLOQ7UFkMftP
d7JAncLA4GoSjwhdoLeQZXIj8EWrPLSwYr0waZhuPZs/8AfXKRY9H8V8A4ZINAsR
lS8fzWqxvfrYXSevnYcpL1e/fRHXPy2Z40st5aI0txDkx03uOhHT0swLenF7GJqT
R+Kj9ia42EbbC84bzXC3wUF2By9gDBOvr/EmTRUZXzb1S6gMlSwXNfUdwaQq6a2F
P06C7a6YfplbSR5u0ANYJrjAniFRJ9d8rEMZYxDV49xdbAdojXVqsB4k0jsQvZjM
E5I8VJb0gU4MNayZV4gAf5kUYDbpG+mgmp6avlfNXDuHMnExa50Q6m+ep07bKCD4
MGELIXoYfzAtOBlOO8p0SkqFrPQwy1zObJBw1OAao5OPXtvcPSwt5YzrhJK2EQdj
KkFD+MyeIYKfqh7gIoXrwV8/nBQmqUNSyBJ+MjIksRTuHSXE9Zfj5Yc05zZiW8cc
kwbHTNUvRRepVisywCHAZGDnRSgbNPjZ7cUtnxVoRHNvSAYBXtKSKzCOFDbQOS6b
7JKQ+SM3UHyVsKymW/5L00dMyf1PNRA0uldpnzStGXnQHrfm7SV8hnmKoNd1pKdJ
LbMPntsYbaS7JJ6v+9e48jXhv1pxBJLqn9Fl0EzVR2N69guEMe1WwZQR37yH2VQk
Z5W7WoOFiACm/H39HQDxaJx9Swc1dbsh1PZpGANggNvzIrK8cdWc1epWIOKUOzvd
cqYe4XdP7QbVo9njzCNVFV2H56GyQg4BJZ1kHMSxb0YiZJbrX2Sqoae2/Y/Jwzg3
LFclqu+ax1v96zrUjzqmKEVLjqP2AT5DUFG2VSDbvdoaQ5Siu18j3PqNvr/wxRNH
kDLkkJOzoe8yipa1MKE1Z8vII9nMSUiVsicO9CKjBK3pIo1UZtL2SD5UtWuFB/Wm
hSHmQAYdXUwhoRyLintVdy90Nf3J+1jR15YHKhu4moRsL+zvVS9e/y90n3+ytphe
WGsl0dhl9cO2yCnf71gAPD6lsd+1fRv+aSFORwhk5W1g7jKfWxyezBUMUmPg1reL
3iaW1hsxwGfCKYdiM2uUHmOtj/5iiuqcqNFubnGF31PZmrTEpLlmEpFf7AuSFSgH
nCscjGBdy7mSvQlCos1wxovbB9+AavdvmJV+i6Gsqb6INp2GEy/COfIAWtn2KgH3
ie9CbCsTRqO0gMRwgSkWXLit3k0K78t3gEmPQ8cMKYMv14s4BbAv7kCxDnkavxBS
VMbOMCwtbU5Tix3/XNW1GKubrBgbM9AF6QGEyUVLosJ8gFp8+xZj82UjAPJgEnmN
S/u3vrv6t/MJtCXaN728+aQbUx0BvEiv/rSOCfKoLrldh9axHKI6ABWFXpFW4evb
efDmNScWvDlUp4YBZGDyXv65QcVYsyNspP57Wd1bRodry7XhD/teZl9WgCIn32Y3
x4UEfOX9fQPI3DrnikEX7lEi18E+GY4wAEPvZEIp/yhxplN1i9HxwE0W/SbWY3iu
KvmHIDJeYiGJkIcZL+DaRU7CCZ535eDSuTCQ5SmcTNRMpZuM/5gklh2wAdd2av3I
CJBYqqq5SNUaHMO+tUfD1Suq/6jF/NmmN+RImqgDkkHbKHCWNQEPqjo2lW+O2XjY
tkVNjXeoMsO5kWHpmzkFjv39OZSUyYca0Jq/eCyvtkwHS6akKZeeIhwLJ2W2zExs
2HnPdSBuIN11dEw2AbqH78CoCXONkybj+dazEocXmIV23mkxK4uy8j7FTfmjlEXW
lYD8JPuU//dsB4hKFdq0/CBlCGFVfkXP/OrTgeqQcLEebxAfnzk+aL8VLi69mQHe
Y1BctXjspdPcbOd08DVkCxUNTypxh+MO2pDc8bAeV6Dji8jqJQMLKehF8RftGyvu
pJ2klOYTcFAHQEb9Xpfqp9Wjr00B0gPSNKdN+NmIBPwi3Op6mJjtrdC7CGHjBAaw
YPT+ZXIH1XV7efXGR8q0K6a+f5SOAKRcOerDLRr/WxgU8P9L6O+odlUWEuBce1nM
n8j8iXxENgF5CcTDdvtygxxZ3u/ovfFEFrtit/Gfx7ZS7z0lOvK0yZYAGARNLcr3
W3XTc3L94u0qxclKuHL5+HbX7+h5g4KSEUISuRx/QQTOlEkwnO5oc3W1nVUcN7OW
pT+60wTkTcM0SWnNGxVA313sN09RtVTMyRRxA84e6oHJLNQm95PB4L8VzJWpHEEy
JzvoiqaGhgu8mhIfpPkLsDBKasHu7g0xaCF8gkV1Xf/zvkQSAGdHk41AAXjVKI08
QKQ/Td1lKo99rEWogbgPgeu7mVMDl4iTo5p/Ab9LDQnh/WlfCZJDOuQR/N6hFBmm
sBfpAjMP4A3Pem/4QXpMVH7OWXzTs5hghdJ2+afMh5Kkrmg0nElW3698CnkoCwp/
a18JQb/rtDnEJUmocgrm4jDLWsBMbrXMRpzk0XDBVJp5aYAtovpxFARyRjvBG+Lk
I4Qg6dequXH42kcY0uw0TkQ9R5DBS1WTwHPETnrkQHOFGaw9GUbFhs/W1brb1y0v
mrZuIs13zBP7mneBcWDXeBTsl8495uttw02q48/36uSG9FSK28X/3UT4ASCnnI4E
pNzkopy1M5li5LP5aTd0/7UCmm6ZnJmZ7CFrpQRUSOdGEtLlu6E4BW8H3AR7OTYS
G3f1SFuZBYFgJXVi5S2hzrWANzcHAT/l5zjopvtX84neYr9jUIICAHQBrov0ztmC
VuYl+3JC6Lne6+7wRBipD8mkwldHKyupY0BvGh915NaTdMom8aIHadmBF7KZseIz
gJknWCue1uGNqLHTWT7Z76rMRHyb+yQJUWzrSk1SdD9cS57PMxhX3VI3S2mDbFg8
gXg3qecqoOmmxxVdVAwi4JNYQM7PlXyimZ3a0L6eWklhR1jeEhCApPlPs6GSCel/
8n0Qk0b7oy/eV0tBKniKBkBNdckiZo0D2CADmFkI4jNQKt6Qrp/05tpHO5VzJb1K
mrPGVgjmuCA7xR1sB8oVmKf8v/dCP2grQDIaXuCbIR+azIqDsIKQLjnGdstB7Ume
3SZ8hJTMwkP2SdgdbPDzdnQQwnWpyetu3DmZ/pbgHE9O/4fY2r8XvJIBD4X8CSpD
+w2VlTH23GdiZCB53GrOzEH3maHxOcKgboJLujD4Ww6fRt9zLjy2AQCaki0uskbb
WL4CKFp0M1nVykmV2bW5KZqAN6o4A6j4XT+0btBHrNCNELR7FM45lwm63KsTWfRS
Gx0RLMETIswALy8RInGcqbzcuFXSHLTEo1Pu3jtU0Cmvv+jTMmMhtlxnrGscDdgn
AaAqzh4jeaq1QR86lmIOyXutPc09XhMU4E4zFGpCKqEFIgkOWNFMGMS94b3jwv/d
V2Qu+/YFkqjKOzrz4Z9QuRw8i90r0VHvA6b+bGW8/Sje++Iy7mS1eRDyQi0a8gC2
zA2arEebLm1gUCit2EBD2Wd0QkZV3pt5H3jaPrl+ZLVWKOCYoBeg0st8hU/dY/Fh
VM1cOPYIOWAw0Ffbnyn5jQir7WI6Sb05+uhsJPAqQRcGrRnri0LnWjnSasnYMXZW
nEVSyQNRE0b0Hr9TOK6jDB684RC0dwk4Ur/cdKi8epmFrWMRF+XsSW9u4LCSf6Nr
35Hq30H6YsEekV9H6JUrYxRUehw4ZSbB5riZmkue8chZUeW0bMy26vALQ/qkOcYa
tAr22/v5WTo41rsseHyyABGyy3Oh7X3qXO4gfa3ylzzlKzcg2u10zfnXiH5An3AF
tnzMoYNOpqlQikvNskWid6l12Tv5Lxput4MUZHq1hDJS0OR2ue5S2AjwTDX2zf8R
bhvxLve+Wz/jjzgK8oZTDbliv3V9jghOr5f2PszGTiSkJv45YW09I6m5SNyZQJAN
XhEWy6ai1Y5rtLYG2oHdZApHusFLXGfjDEeOkNL7jpUdnHaeIASFpFHCxlEBh9q3
ItQMGwL+cL7vStKqmPVwXcHSj1LGFmWJiPI3h+bLNFp0YqHNh4HcdbifXia4hDYB
Xd5D8nsgNJ9riOlDvJIqzaZTZs53Owz/yOjEPeZQWJoJFDoFAoV8udYY8p5O12OZ
PR0mF4t4P4WjpcXE6VeSXIpYHBA9puEWhCfRsNy37wPZLb7zrxLreYvO1EYxhMAn
bBhN86v1aUykS3vRuqvDNeBeDvu1qzTqXK0Bx0ypjdVjJMb+2rajtpqYCoEnP0f6
pxnKMzeKasadC0RN47eXsrD1KCYOjbmnUyQAPCHZXse6UxRVnGJkmnrApNYzdD0i
bGQazPf2BOCQTOY4CLcMQoQQq4+etl/soP9waIJcYhxH2AUeENLJ9PIK7gpzUsSY
93li+cOk1RtcASyI60xZ6X12wB2CYgS3tsHNT5Isi4OoloFhrjHnN1pUu9AXI0DJ
VMB2wtw0cpYX59cBNb00KqUcLIHTypVTfcYWZwehZfg5rAzRdJNcrjmjHlFKHmAd
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BXGqDCtxIx7pLHG6UbzJKIsWfTJpFWVoDJl2PwK70iCSSH6IqIyyDlmArAQdGSjJ
lXM3xvB/3NuPHJos48b4J606V1CY+MQnmBrdB9qRQGY1diHYhpqzeS7rVAwCtdu0
Es31TMoSreQkLvvyb6KXmq3bOoGgHeU2VuReT+Dk0dbUF8YklOQMg0zokem5RtSM
bpwFWpV0J4YVTzIRWBoAqEcynAysw8yI+Pv1dpjTCP9bKJIAnZC1c6BNNHNqajbb
B+YXPqUXbSWVLunc2lsPVJXjggo9Jp4I2ze6s8N858cVgFdyYp0nQggCoVpW6rFe
5EfxCdgMr9bbI8XW1l5sXQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2864 )
`pragma protect data_block
M0OB7VLmazW1c8sfT1ZygoAt1vTQqKsLOR8vfdWA3PwPITX2ex1X+bRoGnzRIyyf
WOnOe/KMV5vxomKSyWrzEtdpZsuqbNiEsAMiE8eW8vdWMw8W9Q9cPpenRwKuB1N3
qck6kk/7/NC+38deaWAiz4kytbAQnl0Jaoeb63Tyz77h4fFbQ0j4Ut//sxNFjcIW
MUzmAHdU1aZ9AQgRrSZp3vsiwUt3734k+cFh/jQ58V3G49oSbI36xqJMVFxj84EH
dq2UOJb4seFego86C9mkEmqJGuNW2a6/Xu6JmKhAXaGyZ85a/QHeWGEi5IO1fADN
OBvI06XWg8kiSWplKIUrsG1hvKF4kJYOorl9ejPQQxzUWLwoij8h7PEpUGiteCZZ
s+QGeDYj8cXLPbaEIEQbzbD6IE+c/ZhQ3a0ZWhToGVWiFXKp9LGNwZoTLjQRVDDA
9gMzRPNCskikSCUCQqOR2tPVNNaos474Ury9FU5RAeFahhxkpqdNbxyg4BQIWxqv
fUZ26jMQZKT1Qp0knCtvR515IJ3wEUQnLMqcYCpH2kmS9YBx/x4azQQmW4oNdwaD
D2iZdLMfwxG7k/GalY37GrOsHVCm0riN4aJEQCS9yDR7mFHIwwErmZlrpjhxICcZ
Oc5S9TBBczbB8gHfDMuL2qSVOr7SH1BHSwkuGcd6TvMBrqLxP9nF7BZj9mdsd/Fm
ZoIwrK2yw4G9sw8biTVv5UONeyhKpu5GSX6j4jQe9Xp+gK+1SdhacRDRp36ZMNuT
dGTj8hN5XAGyCPBZ3ZRQEDYPXZOrsPZvMoDsvUUTqnZZXn/TWfxIpYIYgwSpyhqr
BUfXT/K9FafwrxIKZfz/kPRzwuY9Fk39n4M5UUz80quIc+lJdfZ6LErtgzVv736P
bURu0cB8EtbwH+xXoGZo/9NUv7cv5HJuSjfI2TGLaSbuc/4kDlhwkeEtF2oz3Wz2
N999T63Fc4s0xP9cdPw9E3lSPpz0pjaFMlhqJb6zLJzQVgWKblhrLZiTfjgLEhoI
ZQNvtSuS6VqhAhFltU/xXb8w8KJhuB9sHpnfNeOep/hluIwNMUhZT4e5szcbPlOH
eh1osEQHqKf1MUUfAqvjSkYcmyWOjhT126NKT7ny+/TTTBR5PXgx/aYM7b0r3J20
gyDTfQiYcstiLxS+O5XCXqemfN8k2btN02pVYpD6fLryxYrV4/BWyXMArU+A8Jdv
Czcj58/UqA5vV6Lf00JsVcjlNX0ie5LokgwJ8IeLEV+ejNtEPbfsN7d53+chjLmQ
VImW+CBBj8X7yRnd7srIxs+kT9h+/ISqaZcEAAuYTq11SPPGNhKpHvfJTRF9oB1G
qfTviV6i/NohK7veeBemVV/uF26PX0SknKwGnqx/OoDO9G73U1cG17+iSQ6PpTEZ
wiK+4wzdmVSmj8omnSzSTcQvK2Bvu5zpWSij0uHDNmcnxurrNR/SJ/MP7v+rth87
jvvZUUW3XLuSiD/fFl9PyFgGYqmEP3elzESUwAQO2NFgZMvKHW14W64YjHypxFp6
QGTfq5jVTMKZ8xM1ZBfoIJcThcGSMx/mE7JJJI77kS2H9nPefvqBIibggIVmR0cL
t9UFr4q64PczGDLoRD/6JTlQd8TlUS4p3FQ3NQNbzAKB/o6nz7cW88BCDWJb8nKm
QfDFf2cgFrwCyEvMzy0p+FO6CC6tZmAAag+SWykOGl1a4dGO0Kf0mV6D8MHuhdKY
2XQVv06hOQnTACcZUtW//k5XHH4+ohjQenjnRh/HS7PCk+DgPEBEl7vOWEUHopCU
m+4eqLtJ51364EB9HoFkuJNo/ECGYdoKP3G5/x3X8165/qlYjl5LCv5anO6j5paX
mVEPpJE/IBKRfyaQmWfzs/Sg1ZIK+bTfLKmujTptzjrjZCtEpgxBoMwx2IQKFaOu
+x792Yp5N1IL4eMC46tOjvqk3KQLmviJ8ZuR47XshRZM6WZsFk9A3vtW7MFWUuFz
cBHPoxR/jDByE/P3ySo3IRfXENJMFWzkYYkx4dJ63PQTwnthxzNHv8dPlggEGVvd
ljG1mq5mjTMjyA3Z9I5g01rXBX/dhGpqPzOfLxhMeN0J5pPhZBGIctSy7S735apN
Foalt4Ii0ZdetJGskcUuTIfRpdXzjIu68nWdKBVbajzam4eRCKv3PzRzXzPRYXi6
IW5DSYDBvTSpwM1R0oIKgEC0h30WfTJ1U47KvC81d8UFwtHjOSgP66mc408ZsJlc
L8ArtWxpE6qWVyKyGxLWsqC8Iah6+/iF5Ht+SZPZ3cjzednp9kTiwqdc0Qa/X1tn
g4K1OAHaDAnnuUcZsFLROiJDub4gGlypSpNV0esALw/P8RiK6SWVX1s6vGR/WlhU
3HgijHlo5s521e7wY/MqrTTZpr383Vh1SL/fg/NyWE0G/Jae8EXMuI7v8m2LmkX5
cPOJ2TDOrqRbPqt3AjfrMbYDAhWS3gblVHC1WRNdznfAzAc1SB9fR+U3T/hOv59e
cLu6jdmWYyQdVagNSFYpS0dfKDmYusdV/1Z+sOukKSFc6XQFqd64OxmN6me7K7pv
iu0CSMyi2M2g0SMMy08fRsxpbicLhWNgW7Oxrav1sHu5X4xdP7YyuSRj0v0BZ0Yx
hKW2b0TrvJIAKrukDTqidhDLQqKwXtbgOayX3SUxB1hJ2qS8EdzSBzJ136/UQbS3
sYJCLqVq/Qck75mtx7dJkP/BujvyxfdauZ+VBQQxgJGUap5CvjdL7afZBTo0MO7e
2lT0um4OCARZfHHZRmld/7ksU7PhQFVdSNZa/GBKMKOkvCvIvzf4pp3oS7fwJcZQ
M//sF/WaOXIe5QRHCTKOgC0MUDacsPuKS95f8Kd+Or5baaxrhBlzz9zVO95jXoME
Wak2qfQzo2ODINEwdcAbPZd+SPnNiTtoGagxyjVxsf0Dj7jTQwpaks6lYLGhCAor
UbRaGx+fZ1Pf9l167gYfA5i5IWkf4fViEwGW2XNOnpjpn4TbcGShZvEQdEmPLLxe
JMmMLp/jjSgKQSaw4OA6dteAK4zzWUsCPg5NnmQRia+VpSmhA9m5sE4obQKM49J5
GtNPFU0ZzpdB1/1XxG0YaTsBDkiD7cDzSrpp4rOMaR3JyqYcxbB0DSNvUI1z8HaS
5jKWjXfDp3kn7Z33vUj9LD415YcyAYhTcrUBfRnEht0syddnYl/sOPyQWb85QVDn
018J8GdiFTLlb1ZVtJjfsbs83LGe6PvqC2iJpAzM5qFolT/2smrtWCHiQ1AmOud8
bqss/RQIvIMG0yo6rwaAqva6Y90seofno3X33paIUcUBC8gA5k7ZAhXaC/dd9ZNx
bdv7zx+ujuxy3NTF45dPwn+N/lijiI9FuVR2EYwHsKGYStktkLjivouE6KsGdNV5
KeKDqyQrYglvZ8R8XdlS9NzchY92eeiYC5TBg36AYtGPNdZFFof2GHqPjGB6veBE
QK+Pvf5YTqlIHFME5Sh94YYsXqrBoylOXlnau6QGQy8ttJzCIM2JaEPWcE4FwCqr
Ewt9WcigOqWTrsFlNH6LZqOTOwDLLS2nqZLPf+bfLWEGhhFChQ87cbsiNgv0PLjt
IzvCbVVLpcNiCMnjENA1Zv2uG+HsbtfUSJWmT8zytZgxyK0hXeC511LVvkJRjRPp
pDR+CgcLgkybN6WN2VdehprW89pZwHXbMWPCx4fD0csh/Cgnp1ytjrv8mfB/AhFU
I9ERKi7oU4fYDGf+1dCjzOG47XFWP/1HkEYEu3o8AOUAPDbQ/naHtkcbY6EicnMJ
26CiVVjHd8VYGiICbcdmwIvqCwKio0W+0arD52xWM9E=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
OZYLzJD+qvzx3vHepntvrRoqonhbcjn+GKg79WlZjuCYok0mm17cdNnMoRKJOQkg
6fYJ67n7iXNyiM7nP897mWmIISL4kfftFwMAVQEPu8dn070MBHAxuEGVigKMXsyK
HvHg7Lw7QINb+JhhbIaTd3ba7in9LcVt+b5CT1R7Ij4wbB+RR/fecot28TjGRPvL
1DMYuQ+ZRRjLGqZfgGlx+8Bs+DteQ/TFHzeZCDGIQCaUWEnu+TfZGluruRQ7Cv+T
RQDV/DHILL8V9v5hVgq75GSLvpOXVHBVXITUfpP7miuRjNDHyTQ+Ga7O+O0S+UvS
wmghth0v6dHs9/elTnU0FA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8704 )
`pragma protect data_block
OoJwlmmpoER6JeBM8RSKWkSdaDlvcfmISHGM7TQCf3Ltb9bIblDokm/FS1si79ry
IzvaWfVBkK3AFOkMt/CXRHkdz0IjjmFg+E+tHJme6ynzFtq+dij6fVzNkFJAqmAX
mdtZDfw0xs6fsOdUl0cKiNZtQrPu7i5cuC4N21mGnrlmzsPBUt7kMhdfNyIh5ZCl
MhnSBPyfMPhseisMF9RbgDPPxQUKG0wDrJ+ULy0WuUy95q57G0321CPySa52268H
V5AmZRdtLHk/RkbWFNo4rJ9td8wmbd4nEpOOxojlv8G/HmFnh0I+KFC6Z5/cKZYr
NYfE28vnRKI7GRYUTSu/uhLIxtjyhHRWMUhy0LMKjYiP52Tw7uhgBnmKy9RXSZT4
KZP+0RsDtLBbMdHfnjznNMvf5IRViVBTpjxd2sqwyXPeg1M5siBi6DugS4/TvHbd
Of8B51mYgadwaUdsHtcHxAviekLBA9sEOsPNHZFCBdhnug5tWqpWP0dVFZ8I1mPo
1sZCgF870OHMXnV0SJ3IU8hdqbXBIS59LrdpBcjMIc7LbFxTMgGDBff80XkTO7i3
DUBMMJXyCS48zUExtKVeFf72frOHaberI83UVQhSp1Kspaz6yY16QrjGm/EZHssD
a4gS8ab/hmRuegWmKuD3HXae4mHQplE93MuUKJqfSRa4WqOEHMeG5D8PxiSjWZ/0
R8W3lDatIdOGribOK5lLjClGzviuafgdWgxEBudE45WGsWDE8fDm4w4TsbyHP1WC
2HlU8RkOavVUgbDfUjNjgLbZ2RmGHPgYnALk88W4GCGNNuTwagIwuP1UpZlG7F/a
OhYb2UxnMXjo78aLwE7MrTbYd00rX+GVufqhOz0UJynxIwYOLzF34E0yZTe2qyNU
IE8rNoxyJcy7vGH+lnBpCPLJ0S2BjWTt9LuCxsliUtikLEu2pjvyWgbOz7m0gxfc
kNPp7OSPLLY9PEqvjzDemFI+kCoCLjR6u+zLxSE4qA/9rsVBsO5o3Qd7WHyT2Rn3
VXpGcfgUJzNtJBNoCmzj3F0jDKW2eVi0lIinFp76wfVxIctAcgP/u8HgGAnGcD+D
4jfhWkAj67JqqOprAT00Y/1xK9gHL2fLODKwGgD0nQg6ZorDJUw8EVe8x+3mGBC8
Xc6/bA4ubaGeXqohHu1mZzmBU2hIHSZxG0vbNU400VhtK9uufNbLzq6/vD3ZalAc
JmewdDZC/WJLsA2Gu8vpaO3oBXMzbWswHS3GJGjZjTt/xuVWXfrkQW9JdYHjZyVn
pn4gzP3YqVAVHRvOF3d1xTKP44dX8RwlTHtlnMXU2vWW/srZ8oXRDb+PJThJBnuM
o9RFtQmKAwN4ZMbxfKpDfO/AgVw0TE5qhM8ueH0rSfp4bK0Pi/kJzpPeHTjq6FmR
NKYx12OtM8lDdrhaLgVq8BOO+LlQnX8oM8jRQJiCQ5puvgS36zohN+1+38YgcvsO
izH++O3C0xEq1ARaCDGUcBZvsyKo2zjSIeJTVVIOBB/lIV6FgzJ19QrC+BD9JLEE
79gUnWD7ygnRk0R5vlloXoLC9GTvs4cQ8w8LJbh3yYNu3qPeHWGRrlSdFBrhMR8X
T7KYSLn25xVapTvdOmHPduZ/5BmSDj1l8IRR+1BG4Rmnk2iKU8EDnTec6SoiGHxm
p9GikojPC8W4crCH3Y6gfBbWBr2z6q3GywbUH1P+PvbYljseBY2FZmQIn6UJraMF
YUk1VwDp0SYNVYSn+BcpUsfNhZqAwCfJA6WXgkiG4x+rHyAqsYaLKuiwrWFLUFxu
o+4g5wQS8iZBx7LUfCFolXxKyqfUU1XNU2m/MNSBbL4IEvLL/1DALK+Pxy66UJ3b
r3RYxpB9Hv1nwQSLUFAp8dSIjkXDSm5sfCoWhAdjjRqGE2Gf0O2l3cpKTvdmG1TL
f4jsbmFXpk305i9fRVju8Z4Tn6zNY5n3nN8w92KqMxYrWs/scItuYbmIXuceaB2F
E6oGtn6cYFRXvXvvg78C8vkViNxQUFX5rCon+8iPWrS4IPgnHQRBTlarqcmf7AGv
IGTZV9ELqAznTfSzF7oPSmkAi7lbSIbQnXGSoB5/GGjTCyya19J1qUQMOudeLrNw
7xtDsAqj07bswEWQRUAZKlxULpoVbpkAU3LTb7TX1ihwvOevyvQAlkn2I7j+/KA4
J1+aYpTncrb0TzRCMhgbHc6+Wzn9bOAnykx4L+qIoTXQrTs0FHoAoFZlelrGDfk2
nsSI3vxL7Mr2TLEUBeP7EsDwnT8J2USRfakpfWfAxHHLKINXiX1fqAwK/VzbI/z/
tBhXZKPhlHiIsXKIM4maC9mlE6qo5A5mFGVZ9FodzPJ74w+SkZqTnEIJIA6fTSp6
vbCqfMtwIR7D4vsMfkJBhE09VnpRkZFV5BH1DnxOLT2bOG8tXL6Xnle8l13P/obP
UchuCtJVUS4BM5Phbhm65ORA7JOEOh5sGbbafFQyLdqW3mTuBlqNcCkM702pKtFF
8amyXAaYgYkcmvSQN6F78E79rO97uxVKJYzQVaZreSju4eMuJJLkcEwkpwRvBoA3
0HvnqQJ1mmYMZuB5+FGYSp2JYtvZq8XaH1PXG9Gk9RXTyUz4Cin8D17Vo6QUju2v
VpBgr5D9Mw8sYZTg7hhaKS0vcdaHBadEC8xiaCTJzSOshpISWmpmcU3VP1+IAZwn
l2+zQSaKNUk+WLgi2mUx2P8++fr5eG8tFRscGr9lvhtzIwjWooqAwDIX9VflhCTc
3jROllXiuYJbS9pGGdF4UCu/DD3tdvOZLhHTqbJpw+6WJCg/BUk7muUhouP1b0rv
g2VQ0kUBu9cgQelBNL7BehpvaWqdlWPTkw4OYpbOuUiUR01bYrfnA/fvXuYTjW+/
INGVDa0k+UJY0fiX06KdBlawbT1VsOU8PyWgWKuBkWM9fNUhHvQ3KzP+vWMYiSmd
5Kaza9GBJ9NKPUtqzH4syxzPcmEd01+7/We2Pr0bAM9Gf1vq8Uvj4wTt5UN8ObFE
F9d418R3gSzUByQ55538jsMU+YJYT8Q1jMaeY6iq4rrTK8q7oqBJGG50ERiwUhDq
oi7etqc8RcC4ES9kXgAqUf+tE2fevFeguZS8T6gUcOFBPlePIjR9owQXMkBi6C58
JDF3jNYSzF0VVLCCt8wB1oKnzZPbpKzha7S2dOK/InhAuYlVRTjrmImuKz898R/o
1y6jkBg1U4vIDFsl0AiPg4b16FiFJ6vUWFWl0JqTpVrdnfL0BCmaulZpQFLXUYD2
GIX5WbYRo/Na3JClAs4eAdqMtZlVN+KNJMSItR/UuZYM9TRgGo5DrQLGFQFBfX6i
DFIgpD/wLy20hHEO2YQyYzzxjRWo9kALEEFEwlEpsGeYpHG9stWsnkE1Httw9JMx
Y+4YZDuW+OBIm140+eIjh9LtASJ3jnUfzKr1M+xdT25UI3qJSjNI3nl8iYZfeB0A
dnAmaEUsJeshVq5n/0hLE7x8vl5sSQC8uxG/c2IaYGlVXDY54oBG9ZLcRHjWObVe
LP1n6jdpZGpZ73WSJ97NaO6DvAuEP1cRELV0x0kpk0DziiFub26tqHOUwJEgW66G
kE87qxf5kIJ+l1tz+74hjakVDroU3eheP89MfX829m0T4d5AwoX05r97VXgaj2fp
El9zooWlkcgj1tQ3yQgN+UhRRXv/dLvLcelRFClbqJX8p+/U1XRkcjmz1DFkKb1Z
OFYNADho7aEumbn5UnI4L3lV4BVz2Vp1uLHgiUUN5D2QCR7hdPiJ41qzEuzaQmEF
9uGOP50etuCAEH0LH5AKvV5uYjDKtzbVwRAY3G7EaUdp9P7R3Mu7qfKGOxZhlIFH
KJffNGYYuGNQ7QzE+DCJ7R2EBZd8uTNCY5iUo2aq+rTKQjf4PTQ0o5kcwoaN7eWm
NwPNvT689xl4m5idq2m2xt6SqdGQgsyseu+ZBlZSh4ewWTWMP0IngwVBuSxIUG8X
Nm1BKgknQroMNe8mOjqAqUq6UzMGFZng6USq//YLnJZrAPrhBUIdsGgIXRXUN1r5
FDUEkA4Q8qFINLAbezjk7bIFfJWzpdVvTcW1wnq/8P44GTGlbbciqFxTpopxAK1N
anSP9pbiaAL1GhNxYBrtjp0ExOSxjxOhSIY66GC6K7vHglEiuBV28R+zqMbbcY++
fQrX/MOsP37VaLKKoOzzc8JiPXxIqhKyu1mXAnuM2aKRtE5cKkCYo3kqn1SpwnjF
rCWhGXMF+Ay3mcssiZmkajgKVhA4+nzVOAXvCPOT7tBF5SZ7fzb4xhDd0RT+qSAh
fd++7Ktu5UDtaeDGdhNIHP0Arv5XTlwHcTAi/QmbofzUo7BQYV3j4h3oyUN0e3PT
FP/m9h1STJz84GaejQMYIC+ZAPhzBb98RokQiVrXr//3tfkzxrkLIldEy4Zl7fKD
vckJNg/ceaNLdj9LR0pf+Uos4lHNZGrGlONYnXLuXERaHelBlGJy+XUieujMcR6d
k1QLY1Iwk4XP0LsjfSIcMPHRQB5k94Wxc2BfezicMcGzhNeL/2WQxd3P3nsyTiwG
5ovBSNWG9cZL3MAmg1gGXvQIijM2CJeR6v4lNsgT/fzde1JESIQv8JyX9JIChBxr
xhaPVzUaNR9v5HRAhLTEW58A3e6bH+ABHYVlHnPnS5qlxM2WXqqkWQnyoyKVrTFy
CR2WCruaPoccALhPhSvAdDUC9BzK6oHIpgCUAQ+K0WyrJN0DSHUGVnvDpouiEcI2
43eTxNMl/BdHtYkiklp153ZQ5GYiDf+OQjQEizLZGrCmLSOiUZZC7ufzpB2OcXFH
ITb2rOJ2OqryPiUvrwTqMgtRyP/Fj/LAtO0mfJXmih61hXRDGnd9Q9sYN8z9apqS
syK1r1ytek+4jy94+YpKvmho+hgDPqI9SH/sM9xtRZ3n6hQNjRPD6CjQG4Nr2u9B
c+cE1DsSCClAcJ3K7UPxkvVi/+97QTqU0HRL3ikYwxLWmEa8k3AKjQKuLbrfHhxP
w2uPdNAqBzwj982o6+j34dgngQ0Io7NHMI17WAKTvVFn/dpl2sHn5e2ws4ti1+IT
07LuXTdhUIdbmbw7MoS0MdA4932szr9tvatKUNV5QJrTvqvCn3ixO/EFtndLH4g/
KWqCF3WgLsT8NaOxn/IUXckMoDPzxs37CzpUssLsg7VcCl09MXQNvzcch1CCumId
71J2UoUPxsYAm/3E81HNkTbdy7ffodt/y+39tdc0+Z1sJIMF7uFg1arOjHexSCUv
B70bONUEGh69sukuvS5rw/JalgKAZWteMsQIk0b3h8EzxsrxkgIsuDh8evtXT5nb
TeCA+OvNxPeLnfeULvfH0NO1x1jzPxDUMo2S4/UWWWjAAhhcXTuB0SWXiFmf4QS8
t5egy3jtRstkTwXvm2HwLagYSxdIu1u4MrX+jGbHghCnnzzDTFqmD9OV6s3nwaqP
w/EhvyZb1fUJxPkur1SPC0u+J7BtTQt3Os8kTgcnaYfMI1fjb+ILZFjQ5HkwwvHd
obtwDKpGbLFNK3MvrVJ6IiAZHM5xkp1dgEKgg6R+aRe4MM2f+LIsz+Ju1z6ejk2X
g6njSEDCJDBxPNpvKsAwKTnsj1ex4E2HVgXHe23QAxAAH6UuGAfs2HQOITcRPO+Z
6lWxuwO49qUyehStGlBzhAyF3IbNqMw7sVjmqczMEXGt9wiS4Ul7MaR+TrgRwT07
NzmoLaLEeXyfbfjG4Z+if4ih4JnAQJF31/jcMnoA5GWQwzQw+cy4GQEex+sr3/43
grWHSxH5H2kv0l4ZPxv0mdMOfsPkM9KbO5HxlfJ7+pkPgwcTGk0/3LVoOfWkNL0M
LSOSd0DOBidcHG5M3sRBQYvo3tkxSLGoZMEj/8Z+ZfI9dGqujoahMXSYf1SD+fxo
JmYuX0Zu1BItsIjO7YvriJW7QdNdM1xZo4BccX9rK4Ib/J3ns2idPMfuN4oMh8Jo
pQ2xT5dsA8OzVO020DBIzz0HpZ3J0WgdaA7ZNfyRxRWzOB+TELOZa5943D1c7OW7
RDbYcOcpMkRBxJiF5FDJ4sLlDPAg1Pa07ggO1XLeoFVuYmHvhII9mn8MvQASsfsx
ztneP+C4RIfMcMp+MuwPpN2wOZMws66VaLkVsuMAarCaJQCL+RjsJ7DlI63NbCg+
7PGZVB1TC8HiROkfvMguBdPs35LCxvgKUJRqatXpmgvj2U1fge9k+KtOTtTfkXN+
41tTlFESx4Ws6iqqfJlWYWbm7ZMPkm7I/wIL/0s28YAXV5fDJ6XxiEoNcAuTL6yX
cRSzdAOlAuS4of0WOFDcd563JKbS44R6yCzJLudOevtdWTa5aJsvrR8HwV7+72yM
f1Z57hosHZScT5QNR29nOgApVE+B+IbDKHuJ+sZAP0PYnc7t0MYxGt+jfBE6ZM9f
PkkCPkcwk5EZMp+0n+jG/KbhiRG5AJSpw9UhN1hEQ+J60FoGqVXP2O0jCfofGT2R
i054QXI+Bj9ABMhXj1LWuGc+eSF3LyepLwv+S8CyB6VsFGv9S9Ao4Yqrx8VDx5nQ
zMIGTBj6fteFRNDrmL31pFaGFx3VCcAT2YKGyJ0/wv2mMI8ktIi+32zCce3e+da5
FfIcWG9kEaPQhStBTnkRb7qrDyzjGVhr2QClpTec/VfTMBpQxHsg8W0V/VYlvhrH
gVJLP1Hfm20He5XPFrEu+uaUs22NAepXab+T+38BdSLG40j2Ufaea0uX6TqO9e/4
Rf4Lo9VIQ2k9Uk4GmuQ9TTQxqFZFWI1Okt8phpaE1K3YSC4jxrMTGLs0ka5kid7C
xcDMnhmEjCb9kiD77wvxy8FIEYQn0iiHOZbO7HPZQrl9v7w3OZA6Agikkx25mJRF
XRIqraF5r8jq2dKhgh3oe5ablOUGttyHb6Pn1jOH5uvevmpdGgWP8f0yOMkE7zXu
V3+eGKdcmV3d3bqpvfnv7n0LLYjTAhmh8p9kRwHyT1UGHWU+oZdxkXnEpt/6RRoz
NghPXQmT6t8shes0bDFf+WTzi7GfZaHfX8HL60GTD/T07VhTytC/hGg2I4qviyrY
eipf1ujfJKLGx+hXe1lxHpENu10bcVrN5Lb9D177DHKIGjhak1EBd9IISK5Sgm7q
1WFuo5+YMDPEAmSUNcLDCYHi0CpE4bJYLaUVLsoSVeq9jO768DAIE9NgLzo1jeZ6
E5dlPgm6132yoTONR/opv2rTf1yAYe4cN0CUiLsPm0Y32PtiuGQleKmChzUT1sx2
bzn+KKrp+JKeWyEkF3CJa5BepCeGRdvJKrCZ8NWRdOVErYgE+quKSA1Ry+HVRl5Q
WHwnVG6p2DxKy+/xOQwhjEcmEIdW2UzaX5oD6Fud3m61zgGNGQWTlSiopXvLrFgx
Ojq1yuxCLvSW7uUCVAfkxExBzK4bjIZEj7PzZMmlzNTEJfggaNq717wDECrXJeBE
R0zXjMq97tiJ+buN/7Qlll5Vb+iyewQj/qEhqqi3dy7CfL65CNapqvXy+mqLwmkM
v90QY3oUHVr0WMM7odHCKXMstOOwxWIIDcjfyhQ1dlrgcb6SVoM28b5m7yvxhYoI
8t4RcbBD0fu44bHVD7IM4UUdIZPyJiYtDQI2nu8PbxRwH2fGUap+Hjhs9ACnxXq5
MmMS+Y9TtWZ4cdas4gHNzhTvo2db+7i/7vpI5O9xi/kNij1rqc736r4DsVij/c3X
VEINH9AwVbBUOfmNRqd8+eAvvB15eT1yyoofX5MqlSkPu7tsdtF6Qm/xHJs1V3oT
TjAAUwpmam/2naGVnJGW+IT7koJfp+avPVX2LUUq6PHnrv2aXREGRjDs4ApiQUv0
lUhx8xAT9d9EK5ASkgp54/AfKHfIGd7NPhc0PwcfbzI1PqaIXPa/0IvE1KB1ENoX
A29fyFaYc80nwjFpVJS8zddzGKoYM0Sdx/c0kAHbjM4z01jMIP4TP6b49jEUmRDu
5A6hksSTTHEn4A7FgPc3IPQ24/5K5jTH0KbwSpM7HeAQDI/GaK5ARN8ggtJmE6m7
b4C2iaPt65MuCyTUgPqflUKZReBQ8ImReIIE6wtyKQyqKTrHy0VbfMxpPWZa9coa
ET3uCTMfOlUIi1bCZMJBBkRi2s/7lu112obOfQpVXq5++QDf9xiuZvztEF1Obi10
CYzucGAHnYdGQGOwYXZncfB+AkwNsGA1DBPKCv4fYN9rx6zMMqkWYdieRVIBwNZX
x1FDczeIEQe6ZiOQrYPBqa36JQ3In/Lm2NcscQbuwNbpJo53JcsofdTpAXtN3hvR
AJJuNQQ8MrQIayJF7lokNU22+Y7M4GZmQUP128Mh/WblJvZcJUgtF4qr/2Uoz22L
pp/quXrbGoNDTrwm/8kE3IwTi2DraTZ41zJC6L2qMLqj9cIBR0oi+RN53EOuqn70
roWzRlaWOIPaQqyVvlk/wyGqZILc9WPFN+PWrL4cc4glNvsEAbowiIiTmNFWE/+j
sUc4u1+SwEjEhICYhD+/5ar4UF0wd2amWB9Om3h2Pl6+2JQgYzwdXhz6BHlu1gpr
uf0EI7HoY8b+I6xOjQPCrgvTIUB608UsZmkDvbMDUABAHPUtvJpE2a7OmBOwPTL/
+ssaz2N9HnnFruXjGRgRMQ+yY97SSFVLkDL10YnbgqsMbpi5LoW0AyI7VZmv1bBB
M7PFKH+qq8j12R5zYR2uJyZ5x5vYbcO0ZMyAy3X502lMtFPjGn9fJ0MheyECO/4m
F2Uo9sfPwjnDbrZQbAu1PbOCMYlQtb/5KwPkX+v/NTFgfdbO6o+O2Gq4+jkHgTIh
JPRyGxMX9HWJ8wJJD3+Ks9wNl4J4c3EH65HMMeQgTVuf4k2QIqF3NUTySBmd1laD
IbZ/VhPxnJhA1rha0bSsNb3aS1ybZ7M2BVp8Myn413KPI1nhQ2A1giTQK2wFH3x5
uznvIXF1vqdWt9mhUCZO5SEgiqKi9Jo/9DZceGhsMbP5k+zghWx8m3RIx8wrJRrE
8ztjSNXcmnulRh7kCx1kzUfxOIEQ/jiYu5B/SZj2nKuhaREB/6MRmcBw5OCv6+/p
YzcTa2mnLoy6AvfF4UtSEDjdZtO4XFRoMB6kNLiRoazQcJvxAWDTNATpbCadTWyu
bLIEGLPU6lEL88WtRamnrk8vyNLCqoefJ9XtgjUh9RoLLhyR9u3lddFp6NXhgV1F
I1DXj02g/A0j+2If7GjYEmsBVb7wJFvKYf78FGfSIKKPbgd3YSgGPSvQWmeORVRo
w+03hE8t8ku9aFbmgV/9doEXoD8Dv5YBUGXws+ED7LJKq/LkyMO2xuscGEaGwQlo
0N9hDwRT9cvqNgoY/PMtz+WG5sE4GjdI/pZJ0Xd5H7VR+mMf141Kgt40+9US42ru
ZYn9M1zr5hQBUPuJ7oZoird/DQl2LEsbw4spWg6liBYLilbbQgpySfxk/2RUkop8
6HsL2AKEg5ryHV7yI8e+EeQpwAA4qZhr6ZeZ9DmGVvXF3v/iMZ6p+s69B9LH50Wq
TWlXzfZAFfUWeVODTmdt4vxr3c0euUOGoZ+gdpcVXUAkLYUq2ijwrzkO1d2GTjs/
tQxAA4nnMPgO6bjqCT5FEsavgVcFNYaq1gggYTvq5wz5Y13iJpGyWDY/lmuAgJsr
wtG07b30S0FKTYgz+T+5YHTdCGtYpBof/lZFvyxMqM4Y4406LBQnbLJgJN11C3OJ
InDhXYxTewcx8wpR1BYQOdTFFNp0QcB+PI+0BTkI3x1rWBuNzkbfrEPzM2JeS7rt
YtIdFWXEkgoC63FIy2P1TUAGdzR2ISJKr/1nB3CfDrHIMzQO8PAgaobN0bhVQwsG
nOLkQJR2wZMrbJECTn/3U+jOSpL9RFEAYMatmTT0mb15EqFScR61FOwWxm5SEeQ5
yEwkf0AavGkqDEUYJ2bb025o5t3rXK+oexZ7AckQaP3osq4XmHRSf1l6Gthniy+H
5GbE3blawd7FqVdNpfCoB38EImQ7SBMXKMcd3V1qLWCnnoTjb8ZtV4PSVojJkGey
dkrnv0XN1PNjLFI+7VmF/tIKa9mRcUx6qMsO1yA9i4AD/SmhymCh2+cTh9MCBQsD
NLnk9DF/a6w1JO5gidpRsEsFknF8fbhutNgmJ7TKjIzMUBrzMYE0ZQLHBdLRtCkR
iDoISKTnoCKXJPfcf5OmrbbSeeyU3hMuoTB8SCYTDQdVo5ICxKdkaHMe98Q4Pfuf
g3WZfqYgIVSB0Q9ySZX/obOnnkuws0FaS1ofCI35YNv7PopbW6ZWpNWq1hWrQAyB
DsmaDOxSehv+Lmmx3y50hv4LCYm6cqy2xOxfZEYgSGV9KqinWyZfag3jIZpO3CbA
/zLprTkrB9kTEOX07KKCdmAB3b04hQLXB4cgQkvGRahWhaQd6Ba0LMrfkP2m6JJA
TufK8jOEzB4CzZ0rI5+lU7EUTWYhVXbVgZ6MeoEZLms67oHy578CGgKUUnApcs4X
ONNHgcZvPElIwW2xVMaJhOQwsaNnkE2Sp+OVDuzTTmpildSGAexw14BokJD7SzsF
+l+J+/d3pYmkL70jVSvgauKrgkuvW/k/ppkswiWuGo1v1N7HD9URR0nnppc+uZUX
QYg8E9V795RPFTVGvppG3LfaEuoxrm+g6o5tn6mKsTj/4G83d5fBlUA1uT3za+K9
avG0kpZMsO19+Qwcn24Ih3fBvMnX7pGh7yEEnHgW3TRnDc2L7OfHq8u9tQpFDv2Y
50yiyA/BNI8iGMXTG6DPHO86JQJCVc3fS2meEGXcH5ZyPWYN42np3JCqGtD6eKwC
LJWmPOotBhYXTJXrRtTbsFoIyw00010qdLH7StTQ+2QsSgangxLtSUWkS0mttP/Z
pVPZX3YPt54F08tlaNDVeSZ2IMTMq0dG/TZHA8yj+9PyqeQ6BK5ZTVg8QEfCygUV
vPMECMg2IklgGbP5hLuSgHeImD31rGuM7IxQzuVcY4Ec+GKMbkC/3WEComyDFv7G
DEIIISYOHx6IeFKlgpTtIzoXlKqsiWgP+hUqPMgUjYVwpnRmV2SMCnLzlhyjdkXV
bvyVYDSfZ6LDKtbWJaNR8hnRSCSIvRo0kqiJMqZcRlfG50P8FgeM7iPMzbJodjVt
NH+SP9tKs9rhZz8LI5lRqg/q4M748TJqwdvzUm1Eadkt1fXKVZIsiLb58LYpBxRy
hY7+xoICHBxBCrCoyvSjhuon3+H1LAVka8dAjMau+ne5xepwIT81kBr5yAyS66DQ
f0R09libSzUnqeoa+ejXk0OVz6Cd105ArcBaJrA0Fgy0wQFeCDhj3RfnT/RIAGmc
xLxNvZ7artU1Zf9dJawMhHBMKdIux06NF6s8sbIz2hHJpSblWVVKNqL02N0WY66b
/1xtEn6Mbp6PaC5cOFaqcGJW3+AYbxU5PvIIednK/cxukAMlab5pZANczR+08te6
1/mv+8nfuQl+yeOPCFCPr0tWqGTu5ftt+wZyZy9D7IummrOHGGL09NctDxfeHtQt
uvZ9GI26x+kRcXfe1kCeuaGsKE2RdK3Lkb0KsBEuNt4uVgM8m9kMtdQxvUAlPs61
hwfSIo+pDEKCZcl2x/us60m5OQI5UKcblE/MRgwujLDvcFV9Q27JHw93mKOI0iYP
obhLOgZksRzQ1ZDsrDZC9w==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
M+Nfd8w79VBEUi+/jElTEV0EEVvF3ychWeoK7kaK+1M8EiYqmv3sLRxYUp1vc4IX
cLuJOcWrYnMJ+HOwBSzRKhbChuiI56GCcSRIDotFrjm1gTbABfRByvu+H4QVdiVY
uyt8xdOg+huE55K2ZdhZPp/8fVcy4a5lQPX2eSmatHQBpAT2ViUYAvCl1jNAtzyk
nyjNY2NDhGEOUM1c3Gxi0KFc6l/if0LYVPYRIcHH8DJBeZajCZZOdXr3LgliMhCv
BYxPphAZ3paEwdDXJuZOA6Dhhcc+S0Vm1nJzZy+6L9Ld/6kFPMdu+IcgubiXOlyf
/PWxxEAjtvO0vhZi7Ty5Fg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8400 )
`pragma protect data_block
xH7GoCsNFGVBtHr6Y956mIql2PnEur3hzhK/XtQfxXARUWev7UBOabVFf8xxGL9Z
ah9wrbKnlyR4WbmotAXtkB6SMXW3gZiqw0fZnXCY2E1yrJwWfCvCTrdDA7LxzQSG
ieeA1pecmR/QDxrJY/e0ylKkw5jgd+7vxgszV/7CfykCVlZrtwHlsvRdG8LOUZiQ
asUBv1UaiBPa397ME9xG8iPTjUQlDUchuhBFvnQfgkB1LDOblzZDQg8M2Zyh14MB
Ridss4/aMLA2xnFXHqunAE36Mv8+ktju2OI9AVq50iqH+CtWzZq6Zs47xPZnQsip
6SG/9l3v5w0aGAfsj+GXRnLz+6IpNdZCETMioVgX9XQVHsoeE23VyIDYqx0Viwyg
fssu45tQmaW53io8hZ2le0yLIWa7ndHndbcrm3TEDiLsMQOy9ev3fyIAmUKpkzza
nMVfJOyd/TM+WEl9PvMdiHumaEoecZ+I6nb4vp+VBAGjYA1pwnufPRc2WJp2n4eM
c5XVW15mjWvLpCrTSZYK4R5CkxZbV9g4zRD7OKhI1C0Y25Wh8PuXAxKCnjgFCefc
7O9RHYRmYnAzjZsb5QCAx1Ncps+OMxx4a0iOHDSojh34t3Bwpd2TnxLkDQY2147a
N/O4BG3zl6gVeI4Lu1f1GZtZ4//v8w1TDHhM16PkNVyUrYVbVk49ml1azDLFuJT+
zNC+gOMucdAMdGtr/aEBPuXoQf2hfTbypW/iVr1XRoPava3BFhDpVfcUfk+jfS2F
4RFwgbtNWok2Dvu6uELAcMnPcKPpylPFuseUQvGWGZQd+ij2S64ByuffQbHVT92v
MojqUqK1TDuQhefRszMkGfuqLw2B/EsOFe3ZjhuiuT09nCsviRBQIj7/l+glZgFz
Z/0l1H7Ug8vROxBDj6uAwigGtjdZID4B1Cgf+Bj/HQWmap2BMYbhenVIPCnCpt4g
oIl8vko7mL4pA76fJ+DqWVKAC3uTgsjljCmaO1I+irJJg86RyGtk5R7jQVsjlRCF
xsQKlMbSa77vjlkXDHh+8qURGwsubQQbC3nUcOCkCVMoer958KhXGC519rh1ucqO
tG1ni7E3WXR6pWSDAGMO6jL1L4N6uOUsOL5ZUa5cQS5Joct2qTDHPdQy8v8WcAjv
tVw7dgjyg0FtPPv/LLELEEPpBs5Q7E4ZUu/8CbWHKl1HReswGZjScXioRvi+cHSa
ZVzKy4+ImBR968nzfzh45pedOpuN29qfK/qOFb4ko+fo/cHeh7dgBWxxZ7TsvOt9
sidIS+Zp8gUr9Bocp17xgfSd57K6PQKdApx9uYi/tXsGLWXbxe4vVtr/VS+Dny4s
n1MVYWigIXFykYG7dP30n/JZHlY71gjsx6B+pYyMkZF9kKJqKNHki6SKI20MXtIH
taCO8ES82foYOgfNtUgFGdJhBaWHv7X1NVFiBf3uC0WvL6OqJRcJNvQ2E9gHXAC/
8tjr7hgJv67zz1FWSlv0naYrq9LsB8x4wHGKYbt0UgOS1pQ7hpiQMjevb/LEC9cm
QBwifLbA7DkVyyS2bXr+Z30KkHxQMSjCgB01XGGHiy5gzLJAfIo0NhQ5XJo2w1ow
AgxuJTEeXzxFGkOvh+sVca+cZA+mj/B0wrwfkws7IDnqqfFbi1nnZi2OFNpw8cPH
Y3+rSKx5n9G0Evg0TCg/mC4Y0YYWNgCw2w5sJX9lCA7PM8LyHCSia0TuDc7TNETj
FuI7GPWa2QX1Cbj57qqUK6LGfQ5IcpYRbTMOxEqfOqEI0W0CmoWpxjQ1ylhRbKJd
EOuh+tt/yeCdHn7urqFplVzLrvQeAmnSvSh8BxWf1PncFoFkOFYqX/ofbNgmSC80
XOTuW3ldo+BizDM9O5ntvOu4ccr8LleZellWJmsWJwqLaQTNjbQnfBDe24w1G3DV
UPnJ2XIzsG0EhpXX+t0irAHpoYBSXBir2FNPOO7t7d5/fbxkJ3JYQ0PAWgvu2vBv
b6VJECizXveasY5XpJ/Qw14cnxkYJmeFPxhZelY82jfcYLdFtmineWusBtzL35BJ
uqbvbqTIUPsAF2jo8jGq1v7uY2dOFovQzINa1lE927mJmSe2up2F+StFHsl+RtOb
0I2I6+aT1eyrc7YIFTI9pRly4cSXPjLyFPmf9HE0nJ3C7o/Akt5jpQW2zZ+wVJEa
utQwMEtbq8BC/YicDy82TEzacHFSq7HwKjbWF34bqf+opRhL1J5t/cT24qqw6ztv
tVk2dI8oEnMya4U7aJebAZz3aKRfWUvWMHq1sW2GGw/Ekp/r0AqEnR5o6JOGpPCO
+tIVpCzXK7PQjAuyPwqvI4LAKEknTA5B57rC8OTOnefSkdIKKk3A31ut+OKoCpg4
foDG7eekB2LUNOQc/0+rz+spFimR+lMH0VIkNKsz0cF47c8agp93UXKTambQiuGt
7kcbfkE3rdtLuhFcKfxe9xkY9vD4OHG5rNPbA+S0pte9FfUMI3SylG8SXOAoCioj
+IG8XZdyVMhQ+dy4neQXD5CktRWDbw3wvBSOy2Or9mjrQpWG6730P+FFtpZ0VI4l
6off9t8Z+OnuGTiG9cHNVug/4MlUojnpkR3wlDVWdW1FNtwwrH7aPCGNXVFpwP+O
rGMZ80Y9FEgAVXgsZkmvrJOSAC81hsTealPTWzu2SkZH0ODj7oaUPeyCebCPBpp3
3GSrirCOO/wJpyVnaEGbPaj0SSFl2sBwbpv766as9I9DWFtGnqa3E3FiZdqnaJuu
Cm80H8iXzcFI8RXp28N4gndSfvestfS0iHSabE8QipOwO+yVIkhtZ+uxGTbvUOQS
M9tiiMMP1jqbflEppaUwT0bmqw2J+x+iqwBFYdjhiN9gE5gHz5FRYfVXpZEDwX0K
perfctSDpqxWOThFGwszp1nl6YJS6RX/N41ekD6USOCUmNkaOVCWf+PTARHVgXYa
gCAAhmLIgGBN1VXF0zAK+ZDJU7s2V9LhUTwH9hoBCRNumIKzcXz6+9YMVY73n8LZ
3lb01UqE2km2LqdTQCJMNUaK2fIcbRJMcXmLZHnA3B4zLEC+7nlt+k9GjzO12wLI
53B9OIJ+/Q9q+IJQZG1NvPyWQDBuguOjEHo0xx5AORPcv4aJvdv8T5zywA94h658
kaMhYpqct7RFM18d66gq90DdVt+3eoCv+PT68iiKyHzlV2/cMQOOcjPw4/oaJZP1
NCPbX9k8s0r+rT+gxl/P5yY52959du9Al3Co87TZCWqP0a1YKsS+FruK8FyPp2AZ
mPegpK/I+DqLYwMN1tRrTwGTX0Qujvgpw8BynKGJfOiOBjhYwt6VZI0CGKZWCIl0
3mU6Ixy8UBMiffQpsFhqYUWoLOneJJZA9JEeQ0RALrm3sgATgybqi02a1hmzqgl9
G9k7fwxY+yySyIJR5ozXGO5bK/qZUyW5bMAVmLjzF7XTJ8P5QABwy4brmAulix2r
cA6qavSsKSk8cUn8na0KcYICESPoyRRmi4ASgrEzwMHu+gGsZjS2Gr+2i3Ab1nNX
y50SF1JLNos5B/UUfIY3UKk7VFbBr2RGN4uAYcvURLAmfbJ3Ez7zCJGyma6cHAUi
V6BEtnY3jIxavKyor+sxaoxryypNgHkJ17kTPnP9V1UqOe2VlKeQBtWVMdq9/Nr2
DNoNjN9vmadOW/CXzsQKPeBo4mmAvCC22j411bR1fHZIeOR0bfFg8LSavkD+8evH
1tiPPAu9xhEK0ioD7qZioCY+oW6x99aUaylmGSX49/pStY/29WM47GR2T4GRiCZo
OKOE+qm7LLTeC+sBCC2wSX5+KLm41ZZD0AKzf4PzRf4H6l+nQT1PoR1dg/WCOTat
eDbHvqW176wIniYbmvd3oFQpOLWPvwYPugMPepxYrmj/QODoIkKfXCIKCKqs/TD3
ui1/4ABRHjN/GjcPJHUQ46Hpb2i7smPoHATB8d5/B/vj/1N03M6WcnnJWGQ9x8hE
HALso6Vt2fZhp9+kZqSQnGINeR3roX8JIzQnMAcl8NrHXM8QXYq5IgwVXnneuy3Y
1nPdft7SSGbXsd3RDKekb3B5mcWOrDxLXJHJzM+oEmXuEZ+ik44Cky4Brew4rTkJ
dAv9C/Tg/neUbZeI6e5hxS8rXcXfYhsnHrn2y/Tgt9Wes2xk3QJGGJQJQMonCH+1
9ARYXVXQtwgnDZaTDn5nkhZD/LcStGQvTmwql0V73FbHWo/cIQf0JLkLU7PZlf7Q
JsjuBg/Vyh1DndgbtYOR4ULTRIrSCx6jOqf9lRW7Ps4FlS68hiYpi2BELKP8m5yv
SpbPykVszK85oEcFeGOlCo2pQn4UGcM+I7ZJcxHM5TaRNuC15q45odsbyScCZvs+
fKRL6e80m8N6JxyF8j2efwondbNsczjOx8p3nPs3nfV2q45bjKtUYUB36nd1qBgM
b5OWvHPfDr5+EAz9B1azRAFlLJInDVoCH1L4vrTwbO8gtvChDyb1qDt5jpb1AtHC
5VOdiR3Ymhc2QlaMQRsci09/SVgeyT1DXh5xzRhhzTVfPSQZOww546isUVNF6Rz2
X9MjD8bX4opMaFIC1yRDjZclsDFUYkpvvgNa5A7iH7Uu/GH6agX5K52nN6i0GfRj
vTlORQHCuBpNQw9VLWIQJRoQ1IriRMeJ/SQ7seJ7eFMhQjUERK0Bx+eteltx85lr
yW0n43vkYgE/IWsyyP7MAShmrj4Jj4aV7W9stV34gRLDf8kqxhYrkRusqK/fmkFv
9Tat8ExCQBW+XJ/BGNa2gK+z+TaZeb71lIpYazBLsr2pQKEBZf9JhnEal6jTE3xD
g2ZK1i0ceEb9JwgCzINGNJVuJ+BEltA8no0XBM383Oam/Q1+HJCSKDrBZED9bcgv
IZYblwxQDNhoT4EpvZ+7vs9Htb1HunxfUq167uuDEtGD8+KDNxig3sZBdFR5Z+J6
VWUX7ljA1gi2KEfxE9eom29AQ8QBjYkLs35RKjnFuAAgj4oNT73BN+KqMQZHhAe3
/f1KpUvz5ppAiBjxNzf4K3Tszuueb3V5RAkKhuPPAkjMqzXBzF4y0W5AGq4qRwnr
Slw5yInrw2yLIEMtuZlE8NYVGE6ZIES5V6Dv9mqrCO+aIx6qp7EF4FiYnPtDLwoe
6L1rjuycJOyK9N0CEtftThEWPbspClsfrmg4Lk7Ucvx/ugN9Se8RXc/8dP8hwF3o
KF4EBGPNZTTrA7gmXA0CeXmkJptpP/4N2ixyqZbEzFQc7xt3FzXCW1S15nGEVN6I
Ipyy2RmTggSDRSZyDZnzgSZAAN9ldLSSvGnOP7l/OEMicJe0D/uk2DKISvkGsBF0
OkVx+gn35xTRyoSwXgdHt0lphmnDK14INnInZNZoofd3xdUr9fYYeqHQX0CO0ds3
h5cwIH8l4Utuz1Mn9+f9kkJMMc+dKn9BP3XvZ3WyOWL5WIsDOCgWqlYbRj/2N4uk
ZVLIz843g49qHWRnD+shtTEPJyaL3Ijh3d7ELar3d0gbaGevpAxBwbHntCAMeAwG
EU9Uv6P1CT/MTVP3Rv2URLF5cl5fL9J/coC/6LWVymaJYxTGOm6yBJ4oKcdDoqBF
nzNOKkK1iUje5Z4prVRzKgZIbIQxHZyzqmY3suDvbhVPx6+hwo92dydjxKF6eOwJ
zJ7bdX1HKrfDOZ9+cW5qNP5NHyAAP7aodppjMxtzPzJvt2W0u83/YrGEZz2/UwCP
DOCvt43I6x7QCfWAElV098eocFv9Vqsaifzi5pTWke5gsym6xEKCkd9J4uSSRR2J
b9Y0nbBhG/HLDruE6hwZmrNxKyhg/qbonmSoQlD7Fls7j/5vF+LZeVbITyQrM1q+
5i78rp1w63xzyYpdqVYT7fzxrQbcBUxclzFvTLi8hxwNSdi5bet5P9b2nfl340Ff
MmgNVJNe1veDIxhs8c9a84jacaGywnR6/Jx5/QVdQhgDXud29AYornieUBANN7IU
KdKSC+viqdIqdIpONhyrycc9cPs4TJafcLke4zmcrFohh1WL7ON9p2JmbYDva/fH
RIE2V+WU4BfvztcWHHG/KeDb2P4trfZUEDLjG9A8OmPy6usUMUpr0ZRy7oEiwYUq
5Z1K+XNlZNElwnfEJo0jcu/jC7i5Fw6DsL8nMSBinmtPfA4TExp7Ss40gAxDkHSU
a63tpJEybeNj5tQ4yccU3ejQW6XlJe/thmeef2/2XPBPRdoI9pMjz3Jt7LXT0iOe
YQyX4VCQDIkBVpXZXS2eIv6G/JYJIPdxQlIFp0XEdFY3jrikyVmtfmni0GGatZYT
RwpCpm+0Vf7FyZVzW3yb90esrmuDNuz0ce3d/hv13MV1g0DmOCpQa4b35k6JBIIr
DO4BOFlf0Ln9g5fuZjFlrpe7denTChsbpN2+1frScIrCw5SsPxBmkFaiYnK2YHd4
Qgmgg7TaImGdNovvPjlTEPrpbOJ6ds7X6RKLD3xSGPQBK85n4bWbevoRYTpDO+AI
IxMy2BEQU7T3Yr5VBR2zYGb5W7y0yNWW3vBUBdQmFWxkOSUMnJ2mH0P5dxKU6o8I
mrG89hyRGlR42cHSl5ao+k/4dBRAifJ1vrzFUX2FNbgLAs6gEef84H93ynE8iAMz
zr0/mprZHQuZn9+0SZIM/69UBsnt3AG5rEVOa6mYr3ECys3lAQs5wa862nQQ8Lww
JTw79Mz4kdK0JomQlbrNm4JH2QjAWcXvc/Q8+rBNgKlDVSgnOUp5mqNOQnJX3wA4
7IB/a1K5jYO/nFmWWnW2+L2SDxG/nThxY80a9mJZV/ZN6blV7qptmSMBACCaKvgg
WCudXzC+7AVWUot8gxL1YcQCXGiORUn+NBY7HTyEfsqJ1luAydqhKYu32jAwaP6r
vpww6L36zaE57HQToZCV+GzgwCkzId1bxA+Jh20PkU1Lq1bfY+y9OUapTI37Y34x
Wr9QlA2Uiomnc47UH62YNRRpdVVqwfI7NuXz3plXNvIvis2ec/IttaP0lh7nZDBU
lhdgMlBNg1y25jOAzVIxNv2N3iehW4AAF+Ao7032g8ZV6QduKCo14aaz6d7TuphG
Dr+xpS9gGacRCVNT6RNYsRkV5OIuYBFMCM1dtpaMeGJDBGt3lLUFTXBgD12xOysF
k8/Rp0brbMmAbHjiM0QwXgD9LDwfgIvpH4eb3/CVpZ3ayP03xT2rNizc+DxrBtL3
KbEedevGgzdPgAdL68246zq6dlvkaGCKFptTdzg62IEONufifq0uGcrtlvRG8/jz
koK//29fjAjV5/DQuS4d6X9GzLRapa4KWw+hEhvzW6JEM9toj2pz3MZ7Hsjear96
j5xzufxZ75HvXiBMgUfvV6ulESwNi5MObGd4z/PCcuRtkbXcEIc5iQwY8SBsRuKs
MeARhTOdFaiT+rZvGto5mY9BBYQ4ysUoTE2PyXDga2nDPBR3dM7KDvGTifSFjSkh
Rn5KTwAYG1qGJLTOCHhvIzJ6Ec7O0esA9INF6U8a7Jh2ebmbOKDoDnhZplv6dcwf
E1Jg3i+Je9K/faaT7moOzsBZDoBfpzjCQnI4hlw8txXAiTTFXeDr4RBH4SoEh4ud
nAWkX8q+8I/jlYoaDNmeZcg6uD9wshNAp5Dfri6/liGllCG7BV3XAqvrBGBsr7Wl
LRpmc9jnx0E20tSKzKv390CHFUrO6GBUdMUW6Ux+QgCFmLDxjKN2dWS3LBmviPiN
k5kUzKJA4NqQ+EZFL9P+idEiR0Lr0UW9EE4W7NyN9AzxHKR5ABQGcs8yMilxhtwk
ZqOIzRXscyeZqSUNU+1PplZkbmUMI8d4Bogvy4JxmFYA4Gfa3AYTcUXPcAC5SXis
N0qpDWCVkaYYxkJN8WU1UFw3KGPfGe8oWV8nkKLiUyE1Cr36PLqgOl4GGMjJYlve
7WZ9f1ZG4KoSGFySqNQa4XYHwgpLgsRnaUQcM0e3iEr3983Vfpgls7POMhw0m5w2
IiHVDguV5gEFs3xthXDXkagRAAucDcMhg7Lx9ZiCuRvQMCtuKsP9BYCrdfRnnwTX
LKpTO7jmViEbWqCJI0yXxuaQKhp7IaB9SUKPR5Sz98C58XN9NpiZsMuPBjz9RUY1
4D2ZEADUTVLpZPQjdzcxAUM0jMGonZAxbgKTl/bvJL3pnd7DrSFB3lqXsFcqtJII
JaF20qY+/pUfm/tL6gc9XoPMdM+8xRJsgiRMT9WwRAdoTFzUzKsE24Ydxl0jr5Yb
vIbIGxJoQMnD0VefQcHJkZghqJKLEuhrgq3cegWCIluiEkIfLkg0fJdESNNjJ+4b
K7w+w2uuduZdkv/gYCvhOvDMvpDWAjpRyNjIax82U7tnVBWMpa9xAI0N1jbV/PuN
V2bFeaLKkE4PocuUo+DvC9VmV5UvIGyQJa7XDR94xA9sr6MnXww/ti+WhN+Fxqal
+U5i1hMWZP9KdUESwQSk7eQa2j51pZKVg3fNtIHCgRkIMKSCbqSQg1WKEoxNI6mw
5gM4gqi10ZEiBoMl1u6e8Fw0hRIqZ4XUAOQOlejA2DMEP0LUD1+B34GdDs6VqIGs
mMKhcXbStBBPrJCf1OPEH/Mrp/GKQtTBARbWyBjVYHSvNyuyHRs1GvIeoEzhi9B/
M6qvgiC6qqggDwW3aNjiWCjvhYjH86AuLCOYJqs2Fi94GJ9ykY/AYZK16Wpy6hkC
IM8Rdqyt9d6rtJUmXAVas07qYpRCkdc/skevcOpdwFQKtJcft7av6n6IpyOvj+zH
cEuLTfRLJpSrB93+mbb24qlgVeW1Btmil3KgxjR38TmSMtjxSIYITRwpmLub4evD
/CnEVyhqjVCILdmcsI/dUJe9AqC5IO5n7iTgoY2DdAvHJpMzbj4zlozt7oLPWLvf
ap71eiCKe40ekSVQY58vD6ATnpfMZsb6iDC55KfWVoyGESe+SUCYAUbpOyWIoR2B
92pkw8EcU66iSwZSwZKyT0fA/JvIWNNmHTe5J82cfEyRqwDC+qT0qd7zhvphsiLB
v353UGVFeim28M7x2QuitHtsv6JNZ0gvN4o89utyj6BfrOgHEUJgq/dX//SYcM84
2Yh1bhNUMwy7W563hYAgO6ytggDFPMZdzmp8hwrYi6V3XSrjDXchYA9jpnSq7uIo
dmxPMXLcXKG1fsf4MiJksMKmhM3h86Nf1+LwKl+efdyW75Y/nveCCChz5uyZyzfL
/1lPGxmFiV9o7Sex1Aat68on2aHJ57esM+IEcaVZfeuUiLOO8C8otBV5w6ya3ukX
WeW30LhoV2ixFfaTYEDBjyEETdonQT1wxQcWG28uO0dSQIVDr+UPAY8X+OoK0ehL
5b3eTDWUZOHau+03RBMkEareV4Lluq6OVV/y/0LWuYgoYPW+/CSg2fX8/noLF7Mb
3ipc8Rx+g9nh3aQBQUX9w2Iqa3Z6o4O9xeD4Rj9aAi4UVfJPfz2CNxxuE6+9U7JP
7SkD2IBDi7AohcCkAxyY8ptS2DBUBNhLEr2TfSPusrNnXOZSVBQhzrcQzTpUGZV2
LlihjNh3pMxTZww/VrzSB28bNTdpaDcON6oPat5mRnCf6kCw+CACk9IBMl4tx46C
6ei5WeIfNB2Pr8r//2oyr3YYYa1p9Qh+8aUvokz7LvQY6ZZXOe9bI3oT7gNjoR8V
TTWsTjwkdhf5cat83bmgIo+XpTpurUEY+iX6dIxJPe6ig7pb9L+qtVL9x7jD2Wam
vC5Q+B0d0zVEXKwSmVU9TadwFrhqr4DoP+VvYbRmFvpZ96fSXqUBe4wcIjK/8xof
mS1MJWOkpaOFyXIu3DWmaxRb94vdDDVTRAUTerYQ4TUW94QoGeErMtbKkwS3HEDA
1C9OSxhBxw1dQbISEdGrGT3g9a1wjlLMIccrN9RoQ+YhKF4ZxYkDpOerKawRLVS/
zt8eV7TSlhdvVVAx2KSRWCEn2DtNUdF9frxJK6QNKtAvAL+I/p//wqLMg+5scFnJ
2w731QQEfHGFFguouWs69hq4Z7/k6jHqFHi3IfuaZzHfNPDalbCRBTD1odJ6ZEpx
Cc3aUipDQliShWGNLFleyRZMz/CZQSDNshbZAZFNw9+rwglfn3nVci/qDoKNRwrA
IzvPuQWugK9pJSoluW9VRsb/Z4F87veGdk6dlshSYX4G370lxByW22QY0fonQtUv
9r3Ds/Qhn+Ze2fPTef0/l2Gdf0kyRaw6IsE1+Y0XsYnICKfPlxiCZaMYgizar9sW
8ablrUqhHhUur//U7KN30a6+36zUE4aOSiKu+9py8u7CWaEYfkxj6QxMNt8g0lxe
HaA+/Crra1ldZhcG139WXQ5ElQeFgerTBl42K0Lh/bHl9sUNou5w+9XHrFL8dvCk
u8NHAPCYGiaB1B6cLHplAgQxfKL5HpJwx2LE3tDT5BrnQLeuK+CPeSmc5uubNqPE
9I/3oHexhCiRAEjNEYW/ZNTQk1D6+VL/6D3o1daYUyiyZleYnuE8dZ+ophn5MDBg
PIph72v2U1VaWkd36EDWGUVnlzIl0KdmzD4WPYv1mTHyBmJATj2OfD/6/8MqR1RS
XVlPVYIB7lq72apH9pi6Y0iT17vKGF19xnynQx3U4Tj3btVHdfFiWKNcC9z73YbI
nshmRW+nSnFwThDTBluXI+9QCLPf8HOnq9LZ5OOFLkPNtKsE6hiTZZMLAwwU/E4a
SUZKrE5NtKG4O8P6ouZWeSpPJw33nonp4A2iXt48T1qEU3qROwxBdZlNfeKC23XY
wdCOoI9eeDgLWTtWclZaFvAiDOkvpderxgHaN4Q7cCn3jgSHdJc1V/2og+6k1M1j
veuul9A0b/9v0t9QfaElTsgqcZmytUuvYDlTX5MT90OInJ8fb0egGCLdtz4fnhOO
lYnB60Nc5whXKCnqQFSGUM61LUECMyttzYXVGYDp4EOMW5l5sFMimsHW5W1nhLYn
aM/en1C7eTAgQEfhpgaTtNT5Zz2YR0WDWHkOlZ9JgaQqi2e5pJGB4epzd1ENJEsV
jCc/ezZYF3XjVTGIWmXbv/6Eua7Ts4I5L7gqH1wH72uAtlhBAGLtvUcNncBR2tDY
6gL6LInuhXx9c7cR0i46UUQcRrh4XFO1tgVgGQprRrLyW0FD1gddaaFGRAEXVhuI
SjjDhYL5qLA01RWqWI6rU2Z+p4KjeQoVFQK+ik/Kc6cwwV/gdDbuK42mdhv8j+oU
Q4ACWDeVqnhjOFdlK5YGLlbp9Rib3Fqf3UAd8u/YpwOBAdddXMJCUDeKzBD8xkYR
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
FDK82Pl74m6I27ibLHWE6Y04Lq2DWWTvHZL8KZmyFxRBdSzO68T35N2O46nVH9ET
QdPkEPrGZ3ouHZaA6nKvpQF9sj/57ayzJwwp9PFdl68VpWpDMz8LEdbPbq/a6l03
JYr8an5np2ZzJ5RFbyBQNKprd/hGhT7aCF4suIRg0JafCJaVgnCaVr47yIqa8A5J
HpLO8pUc07FvePGyvSMoZbO9PJZ7+U4x/qV0XlgPvp5DrS89ASLCk9R0xozx39hz
72bGddg6b+knEJJHwkXrOzqX68V9momdJ/NG8uNLEkJBYZOON2lVjo3ZrgRlu8rL
1qEUvL+wq9IICD7EpjkH3Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9280 )
`pragma protect data_block
8/aPDE+7o5t7yyNCySOVOFPCKv0raPyyepbbVWDBEDG1I9vMrXzPg+Q4HU3XUv9G
WOUOrxWPh124gC/RZkrtIgkWyflwwiJgp7JdDkRkLit4mhJNdk2mLfLsW9oANiRL
T2n7yZjO8lWvbLui8MUjHLX4i3T7RJ5w2FawQmvf49qRczsM4HIw2Ip1fnsl5MbK
RmxQczNCcaVjelPoh1D0nsTk08t0f+Nb9FU6cI8q9f/4YbRbFdy82yO40BmXS2pX
RibIHUn+zE03IOCBgTt2mnwAOw3hhkh1zuEAWkXgiEHFbK1bp2HyfDDDtwtUFyQ2
DfPMiHiZqfRmjbEqV3NZ+xYaPuaEPpGBECtkLkpS0JPUUwCMK1VG/KeZ4ShG4VA1
g4YXn/vSE2bzRTPNfpdquJMihFJhXluJxk7YDC4BBRHg2inQNiajdlnZaJkPQTj1
SZ/A9W0gZkth7osCkU/pp0kh7ah9RYLlIi5dIMFfhTl/ZWhBj2RCfpMPgnyxxG7X
LmN+ieEU63EU/q8mW3yyggZ4kM0yLQ5eNEQB6iafczuc4PO5FWtZz0lSe2t4brdB
7DVv8ArNNE+XQA9mT6PskycRJ0Ok+avREV0AQP1mW3kqNu2G11YyZyoTd19Nmthj
a7KUricTYbLfj1DKvKWkvzEqzEBF4oSF685slcPYSmpujVuAZb69lH2J+EkvGzBm
fX/5ST/GZqvWNOToFbwiuVStBiDC47xbAJ76+Lq2tNe1iY/kCNtIJn7EJx6lLsx+
yuAjtfn4ruZpgqv0Vl+DMJ6vkNNDsnmyJBHn1e46lu7Q7j9XXZpt5y39Hv0Ol46w
s6kx2JDLoLxYWKUSvkVgEKhlIjZT+eO2PzwjiO1TDipxbYikxLOIxGyihmQBqcwi
UvmtLbWGWJdumAc7OZRIXc8P/O1NbeNhKcS+3JY1ydCLmi3TXKGUCcCfKrvuILMP
Js5p39SVsulEXG8mA6UwlXgRgqKi7udNkzUn3VkYkWgO9opfosujWI/O34yFMEmR
w+VDbwmXBsakG4CX94BWaANtDfAnWCct3o4ayfXs/Qb6hcKPpCpwX8AZ3C9pZw8v
DekuSOWV+tcM0lbqZti3JXyqPQP8AI/DiSrQALXzbDbSf5BDgnOXRqcI9RgVWRmP
TTwVp4usy5yuh5dndrj2RdMwNYIId9LoVb9NBnIE4jSr3KQH2myrySrdwsaxh6r6
rJXSM1YdG1MfOHVpSq9B6hcl+hm3sY+PJisJ7VJclYmpYc8oKnRjovYZFiDVB3SR
roEnh/2axFmrSBKTXCSFIQCZCoJ/5JSvLwg2VLcYfp8Ej1NAuEOy1f5tZCUQuf4p
rWT3ijhnv+RURNfyqsOiFJzLKtNKAvYiLHSMNYh7rThTKEsMds/MdVp4c/YIBPYt
N19AYtrkJEfIG25WhjYxdBUhRaT36o/Ty1VXY5uCH0fBiLtBxdbXRpU7ToVEHgY6
qjRWp2U9wA8Kqn/ZoGoH9jquzkAfKzVxPAA0RJ0lLbVRdteqKglqQ3gjq04HuQnS
XXV+CGY//tzThhdr4Niw571sjzzHHx6RswNC/KEkvW6Djb5bx3WeW8QUGtentOir
GOIo3K4pJCOKIpBeHt5ucRD47xSrELTHBK+ooigT9RunwyYb8wcF00ilfzC4PuI8
tPUfsHIG3R1Khs9O0MGmPf7SPgCjT1dq6JcwW54QC7GbluTkf/BCW9IVWNbgd9kj
2/iGpnUqNnfZ69OPRyRz5wS0YgWR8AGiU7IusAEAvsSy6HejTxy6DWytbYZduH/Y
RXORis1uGniIMbsY/HTiC+qNF4UldlN03nIFlkZHTP04vYpG2KyMRd0z1b/NGexn
GE17nO+xXi3vs8FgKtA2086JAWO+77IaALnXY/VhHpS2Q1Qj/mYbgZEWfKRjPhE2
wdecMiA/x8zI9utiy8eN8qEqV7/hPw4n2hHCoZWN+k3V9d6puaMWCadikMbOWrLi
KXQl7r1E2c8OPSMo1Xyse1SgiXN0P+t35/w/p+ukfVfvtGSQJK5hjscru4ahlk/7
8K3aNzsOs7hec6vO1B6fyc2JnbxYfemv7dX7CnTvx3OsTFWABQl95GYXQ6I37Rlt
W8kacJk+LnWhK8fPK8XjtRBKvAZVaCKd0OApoO/rrfhZ7vDa4f3J2s7tflpCVixk
z2P734voJiIxudBr90jbbMXP+inrkM1bwhJWelSVJOVzWNueAevyE9Akp5nsqpIz
DzEf63I8aW47a8fqB56CLN/M/T61inqgU95dXWZocrhUn4JhLwxZgWa+eV9+gBN8
14rN2+BzaDelIfjPcEv9GPVtTH9t0z77YtBH7KtgFpio81u5cQUHfoFt852PJc3Y
SWn7tBSUILw4/Ba7Q4VBXpFxnpcrJMYTrWpyh8f5KsET8AaanCVuHXCBAIuSi3ic
f9O+kMI4SE4qaJbC+xsJIZS59ba43YJqWsHKxZAn96uo44y4kdWPZ/u8ENgIkU9r
ftAgVgSTnBZXlkq6+kWfK0MJAV5KYgxUc/22dlkShaMTbvw2ud01RPnYtIiCad6W
CWBBBiDc+7rdVGKY/Rh347+98kXpuod7f4kt+Cz8geHrYovE0qQVz9daCiAGepDE
8/OHoUp6tqG3rkdP9sDoFlUELUiH+0jhR//PC81He7Q2YiPRwIUnPp5/hPlVqkM+
EZ/4e2+zGAOck+KNGB6zpmrZMA0RQuGMoDeLn1fq/b+/o8zwNOGdtAg1biuMaptg
qD2JVzZ4jfviCbNkrrPOcivB6IJC6v/GfNFx78ZahyyrlRsAms7ibpV4YwCPo+Kg
OCmO/Ayu8l7YoDSPx6w0LQIKJdm6vxgDibJSli6nKyTvIxJjFkLQX130bjdh7Wtd
FtMXpw9EQDAmd5AK+5+onh5SdWiuIIM5VwhR96bxyNIHDBDRXNiJ5eMwTfvlCvi6
6Fr6qr0Ye2PrDsC9WDOC1KsRxGiVr9/IdWKfMlIzLLDoIFl8Fu/chF1hhWDluPv3
/lnYYtf0YL8WLJuHOdwv/mOmuGBsWR1m/e5s6YGAg/RIoYSIYNpAbYfND4u4K/0S
V5Wgka1Tn3mcJ8Uq0gK9PjIai3SLuZ+Ya/8zW0X682jIu2DBM75+0JE+W+SbI2V8
qNaNAOs/3nWnK6ydVbmCeGH5zCQWqGDpLZdX0o6VVgsVToo9D+8/QlU7UjLNvmPo
DAL6n/tiT3BEh9aVVOzFc1/1gpMtd54gcgvBDqACyJHh9MEf1fFgeTsu5RoN7FQ5
l97yDWYdGs5aFSPi8I0oRBI9pfGojAgW4cl4nwv51Tb0Io1/t8xfVL104NSKgiKU
viExUGlECT3r+kfvVLTW1WvhLmlkHHlR+bY51z494pZgG+gN4JhqVlWlBnTU4h09
CLOSJVpi5lzSce+Nr/FACjEi9oiFvtoWEaqHOIOaJKrcyiQc1q1PBWvXYKzb5o+b
ovNsilHkk3G3D52X3TgT4ws/15mtBkOgDr4EWPuFEtJNvia163wyweskg2MArHxE
UN8hAW9VGrmo5uR3XcwOyfwHOsQwftixaoVqDk8gastsCoeSQdt0lTHI60scK5Ow
Jw6xAtdu/+AUaYGysBZ7GLKJg2ZptTzbw0pUf8tmqmMiVlH7L9BI5UHNbFaaeLsw
ufsuL/r3pHxr8L+ivZnBL4wl29L+99u8QkCffXot0DuRs2IiuM8Yd/21qyu/0HFm
VucGnYSPsZmVBIttqR9i7dNDoEjtWk+8FQXWzawe8F5aQmaT5r6VIVjHUCLL4Yax
q5Vm/WlOf+n6kH9A+bq/2du2uEajgqhXatkJvDSeMUZ2fHUUyAKD2WLC+hC9s6sW
pKcHfmaLoXMuMEDbi6t7060MzVJtV98w8OQboUzNEPMLnGQlRlRN3N4EwskJqGun
LcxYA2Sq6kIZ7chgcWNfW4akbgjg3GL6CZLyoi3sMpVjtDh3eJ8NXblpESie/ksX
Is3gKD2qu9MKB8nikoYiDFmm6uw+paTRZumBD/VVSreB8YJPhow+x3IrzlXtVErI
hKcbq50aVULim6Hz9RsemuMKusFSqV6Y70QqniGJ8x/dU9pDls/f1WU3i4asG9qH
AhmxbRmlqVsYM6DFQ3MMxiwnEY7ijldfSs/sbRST5LcQ2yk2FZNhDlwrVBBtieax
EJsZtJVw6a0IAm6TfeJwqbkk7NZLkiot8XHOn5AgO27xxqJ4KlCBwIDrI+bVgkdd
k9xay1Ng6bdOBIIACGdOjRZScgAtp+2ZjZ0fbl/g16+PE9r9T2iLFZZbZLqv/1Ab
C1tcG00ExQSIu/U+p+1pMU0kVtfhjeMy6T2fyp//+oCwhD9E0HrZ14TfT2LdsTSV
XhDqH0pHYZvL7rYrfkwXPO7URKcrGUAP5s7w8Ss9gHMSiNl1erFzrBj3PBxfvqln
/3+d21AOmQoCdxz7w85Wgvc97ci8VJY6Fg6wm03w0u2JLb4fwVmdes/8lGK+3rOc
48IWIWam1YLNwxuwJ3wCNSh4HmCi24TqJml1b/gdy77CZns8Ka5yQrzri7/9Y0SH
hBTbCP+S7ZpXnvavgepIfYKM6jj2YlTmedDQVZ6qCDVloBmmpA++iyJgWxyK+E4X
6g3t5l0QLkJn+NlW0o+kX1NB2AIM4dh2M00WClfE4VictRR2JbHDvXr+Ytd3nnqZ
Kd2OpIESUrqyLEVfxT0KQjolrLgOSUVpPqilPN5zvFOVkDmexZ4u5jrvxv4E1lY1
3p2+Xcb3i8STHdg3LMKCHp/OtcBv+it1XJR5F2fYj+PWa2CfDeKftOP4lLStu1na
iedkNuqfs5FnZu1tXm31KDM6A7Zrz76oiUQguz2xxd2ZWcd/R38RrSFkZaUTzbiD
l4lvJEgTbnYcLtjGeGf7sLcWu9tPz+l1vdhfZFsTaYEuUAg/QuggO04D05J7frjz
VlksT2XnlkFbKiDD4FazOce20zZfzoPks7QEDYutJrAIEvTNROg5m8ClLvcr95kd
X0wctm7M55aWqAiOtYGoX3eK/CBKhoUtdtVjxSyZ7oLtO5CTnLn0Zv9t0Xo01CGL
HSge6KilnuYjhZFekH6GPQkAeRg+pwMLiTUP2QTEFWsv3pdO2cZvA+H6SwAcRf1M
TOmGcVBFhUJybTgKRSS8b3BYVj0NJ4LjTlL/n9ElWK8tzxdWSvhrkxiKBngZDuFR
JrA4l0QGpDTlenrt9teHHWLZ6sQJSAENwEq5vwOjUUkgwsa53dS9fhprsqkQ6xSn
M0eZGxb/0KXjKJlqZW5U0mkFmkhlDxqEaHGZx+DXXJo9UtQamlksV5deUzz6W7QN
v1MFgWxs8rRaTtrKSb72T0FB5rKpH8EXzzZ2WFdz3V8tlqzj/np4Pf+ALDTBcd0k
S8t9or6sLj5lh9QBIHk9OfeJg3V2nt8fxAynH8qWttbMD16TOf8ISEaGqg+lnPNc
+Bmj4b3jSP2g45MizUAZmn63VQ2vCjHwYNvrTJykhKzDQp8yo4vZBeM2sMS8/s9b
aO6eBaOf3+B/jYj7VHeWl5PWtoz9WplfSp0C7c0atQnd7UspMoUodm0izUozYM6T
n0cOykfd3pkl9RscWBiZ6xVT5y1CCBnK98lhKvDhLvaGIYdykx4eIjxCrEAW1dKL
DArecev64VismJJDq3LZGdrrVGBEybOurg6Eyyl4LBPvd27wVXMopkVoU/QHuyBp
hKaofVBGOwXFK3a825Lr9vlCynJf6+VQGuxyu9ED4I8d5qheySRwjQrOgFy4LyiH
SxF1QWszN7wUPQ3FRIvQ12dNi9DYYuMOjCIeUxCzsYVXmXNt6smrC220AMK75bmx
uOy8ymYDRXQmgCIU3NHs2gXP4zHlB3b1kEPoD3kRj5Hc6R9JNuJxSe1zOw1lcguM
LTz+JrGfBuEicyGYtkpI7F/puLCfjDLpzX6KLU5qFAA6PFXhIZdhpZlFkvGy9bAQ
IXSaKPoxM/reEkS5Ntdgume2EVlaf7660hJbg3azIc4Fk96fzI0rK+qab+KoyECD
zqyjnBM7dRfA1sICJ8vRu8TMhTUpBYQas35k6ItqLVclDQIIDrirnHEJSi1eE5C/
T7pFusRH6yDQr7SpWSWpHizaQxrvrktT/pSkxwwierGkID+PVjuzFFHyeXl0Fudu
G06kCmqRuw8evVxjS3z+3QnAhbL2MLNMXHsnPnjqETwtERXFizrg7M6W9mwlGXqp
L739hqVD+wXpNnMTk8ftoMUGHHrnh0jfP1r49qu+Qd3T7olGP+fz9B5d8MMFi9go
3wpgHi7gkQK0YXxxN11Jp9i6iCYzZHGGNeLlTZ7u5b9FVLUj+EBRY3lyk94onWfa
0s4I2cdI5No/f0X2s+uI2HlK/fXXWyQSJUyJc1kwrfEQrJNFtiEG/Ql2rOdwMLCP
NqcwHxDGC5N475MlSidDPpwuNyFjzocuQ/oOt8R2el3RmS7QUz6tRYgA8ca4F7If
kjjPf1WcUjfWE41Yo93Xn3lFpzD0qj5vPeZNwp3mgcv50dDc7vdBitBXjBYbxMBb
ofA6Pn5lU4a6KRn9B9jyTCTeFf+NZlltsR82hjsc0pylWYRfRFEFyn0bwBvRm2Z9
YFwd3UKfdhuh4NBF3RWKU8XpUsWLtyV7oZ7rWn+3Guv5nK25sAEBUgHb9dt3AoyT
1pZ/vCFIawpf5mTz++c0n7MRskQYF6ncLVi9rJRmsadobiV8YhuOseC2bfG5/tYp
coK7nS9J6Eo+A6flL4nIhFOqRzQUekfg/FWncD6fA/m4WDAtev9eFtZKeCoJiNQg
SIc8l2ZB3o1X1rGbtc5g7NLCGn8AqqKsyvIqiayYNqj9QJ27SBRMhc69nAeG7gKX
nj+ZmBvtcWblkO229t33PCHUwinHYbUPEyTyC7RhBejAxgmztloboWNqjfkaa5oh
ajKoLtG+Tsw5xhbiGs4iOvsSs3f4x1EoMdH8YvXMjhHAiwYYFzGQZhsnDED83290
PDVi0RXaRomSqjdt3rG9RheX1Ch+upaB6sbBcZ2F3/l20dkV95IlicHQuB3zPw23
qX6gUFrp+gusRVgXMEucW0If27CEV3GQZANK2VuuWCUcYslxRmAzp7xfXQCeBZY4
hg3aYqAqnT1U5X3dUtLWvuyryTj03pfr6K1DA5zWGPdGzLdt6uxiGWvOqFstZ76W
gHNeknYvuEKGJhP5lq7WQX9MyZ3yTqfRJb9AHt2yUdkM5gbck5mffU6p/9mPwpbd
lPVnyLZYL/KpxgvqshunUV+RNMp+ySnxYbiQ/cJPtfUJrsN1JbwBkICT9y8gLi3B
JCK0GO/PwqEiYdEY8r7eD7ZrZBoUCkoB+XPWf46rSAR8KHrZwjKUaqnJqIXsa4Mr
uXB1In3wsM17MM7PZK+FhETORQmViLjwPKL4dP5BAwOmyP1pebpyeGPtj5n1bdDF
4gg/t02GKSyZeWqf+c/u5kAT2PoIGqwmA4Ip6lt+KMOy1A7rsTHYz7/uirXpnfNf
KPtfD1KQse3XBOJy45lhJo5KfiaWO1R2/C3vhW4ycREBcadQh4qrF5rU9eVXlBck
zZTSY5eqh/UyeZVxa5dNGQlAYVB9AxQ3jkiQVTi61BvClSZBN/Pea26+y9KeyEBm
vrQfpPOZf7ScosL0U/eikaSrI2Exu3593LPDtwJoSaQq+52eKQgdC5nx1KXIb6jb
Ed5TKDSG1g0Efg5mYgeekjPxsZ3/OVdZE7roT4y+1g1uVpYM+1gENHzB8oD84yPL
DPDTCA9AmqldyjQr8+6y/PXukO8C8BUmUT7+m8+45vh9iTY5H/RvwG7xy8syVLWz
ZY1JZ/c1Gjn1ZE2irnzm3qIegR0Oh9pgj9+4VRP5jLI5JoVXdG0o7QWOLyTlOJXK
fxGrxAXn2BAye8FNiybAGFRwnBa69Sf0XOUwBZMtW0S+f2yiRHQUUFy4fTnlGfgk
k2iAEER5QhPpNvldtDwK/LlWzSJ35vOcPnZVgj8vu8JErGw78yMX923YPi1p3bbX
iBbl6YNr1KBfuaXQGwfHnCUNE+NekQLQRQ4RyAf+fs4Muk5PEoShJuvPWk4/sF+o
y8TiVGOqqsV8X3OHoGzbNKjzgu9anzJwLH6vaGo1gTKMqa6v4fJisL5wusA2jZVy
Ca2LLT0KOW1FqV+6lgW0iDowGb5+w83cn6zsKiTub1Mjga2/1RUZsR0WJ4vSlw2W
TY+EcC5eZ1eD85/cfDbgq6vDc5jtcI3mItCHyFhQ5sk+5XxMtfYK/fI+/XtXm8lx
L+vZKYxjsuFE4Cw9kl55Vim0Gb2kZ3vn+On9/5zS5FK+H1XGPXlkfg7OQKIisBI0
9mQcXLV/d7iiPgN1sWkrBLprGYHs9G16leC+2tTyhzjpqfFg886hnPm/l8cgfyRQ
eFReH+ofyrm+MAPq0VIgAVS+fUZ5n6lWsC8usUK/gK0kxehiUkbfQtujJql0yj4x
R2L4W0wZIpAdNLlya46anwkObgaeqfqxfjbvSrlzxLVPWTeDDCrZ7kzi8nWemjoB
V38uLkfxgnqbSWrN0byV5v4IUQU5mJgihdjWXmJ19QpM8CfU8yeQPutN1OSsd8+m
FkameTtrAt6BNqk3aNPlxS0lWgTkEgdc+kuWJ4weG0QPWUdFWYhKt6q3fCskLf+U
ayYN45UM68tfHwETEVM/Tt4jgtwaaNKviCEJdW6JO/BogTrnuan49FO8X47+G6Cd
zhufrX/UK8wK//8KYklehBDg67utzucyaDDwC9Ab2snXc81q81tSE7DBW2Y7UVQF
dDi6uMInCCOdqNGt0kvQxcX9RSgVxPs9y4/8Nsu7/AcyEePIxAKeiArtbAVcImFP
flJIMmCotianTFVUta6D14CDNkfIsVk6T01mHQ5G/dsZa5jrNE8PWiXcnERJMbQA
hYrJj9ANtbhffUPFeFwWsU9LJSpYfuimdeUjD/HcmTlP7AYtC5aFqBESxWEc6x24
mb6Cqu1RAq+Dg0K057I3c25oYjWYdT40T1b7j3H/0XvNuVUlYdibgBXyi2ehHYWN
1UaO+5145/uRXU5RFA7P52kjQKD/fjSUptlzVHHcoxR5r1nrdJZDt1fHmIf85PbS
q9xdyl8deyE1Km6MV5q4qkwkUOlVCzrLCnD4UGPTsoFNZdnJ80NeCJhsUTWjBoVl
ZtbTtJbrn66i4e99Rd0XwmOXtzP7G3LUaqbbQ10tu/lQjuFpwEmeojpT4U2gCq/t
+N5zaRx9VTungTRX/SxqFSCeNorHDQaY5oVvpAcwUAcQQdfCLxwT2uqQFtVEGFc1
hMP+07bzYXH4iCujPw8gTCfqUrEns2pFpB9hReH2nkp7kL1S36i1awoFhM7acDbc
rXOnccLavZdlhdhieoz3G2R+XOSNcc2qkZg+6LV7nBzqTK7lSFuSKv+6/F/cRkw4
4e1HzXCP5vL+ntVEHfzIPZw9/vpCqgNnbWxnm/SdXpeCcKIZHUioQWvxhoSLv+G8
RgfDHJdfFp1GHIDhBe5lZEl2pyyxETrOtJyjqSXodhYCE16u22i8X9fd2Ffddj3v
om99X1qDlElWgwckrUndqvqT0g5OxB4x4mwBB3a5KrjbUTAVk4aAPpT1eEy5syfF
k8oEKIAEb4+43LIGFVRJvYuQ5AEso+v9yaHGhT3cc/qCTk0TROOFTMHYomuK/yGW
k/HUgUkbVG+iwnF40YjSeAdbUhmEsPnDCg6OR65yARNJpNJ1YxXwm6fgribkpxc8
ArJnRdFD2BukF4CmpOj3UWhxvU5bktkyXbChaLXJboZoXFIgQeclXuZKBXqHM+f6
VSBB3V1jCMMnrgxVEplxaiz9dlUR6x9M/1g8MFeHUiuigIbhIRx5/xCHyquRsi6F
gWNWDlAKtRFq7qHHPBPwpDoU9rkbPNWuRZEOqw8ynstgvIbDJl68pFmpwHOTQKyv
dcxj+z2WtsAnn5RwIwDd05aJt0V3hL2yQYiTt5QDTm3qkFbQ/y67T0uWABmBFmeo
PGUdqy5vP6fIB8djvHKrOCx5GLaw9IHRWjz17DoJH3wCaKrLmCmlTSrGz37DZQvm
zIHyISKxxK8sQTXm208asFVejR9DSx1jKWdNXYCQcEh9zQy7cLp5dU+9TWcFq7H5
vw8YivYDJeR7MlzsQTpKibUZaPVyrJ7pLRi5xUqo6S8O3imcX7po4uv2TKtBZK6N
vE8WDp/XQ38pYxx8yOaBw1oFqFBGnW1RaBJHdrTgheH+04aR/tJd+zC4KdGepk7o
jhvt+b7eHcnzXb0SuNn34D06WreWdu5dPsgzBmTpaKbdCNzS952UZFcQlpqXTOQO
LTE5qRuDlwP1S66AQPb7EB4XOCbtQ2uwOgnn4R+obW8Nncv18uDkc1VXTV+LxnrA
klvbPRrXsmLQZ9bs/v5rtKnUkjDvDGcPZCgjCBW1LfJk/QqaXdTDpr7L/c1E+sTZ
ZOS1YVHCI0MMuRKnpQAbK4f0bZfqyRk+q20SxVIswDsXBklLrqiSe79PTlEB5hqB
EF4UhGf+rI9v8qs4fL5vbueSY7y1SvLNeWt9Y5Aqpuw2r4LmHVMWN/AEjEZ7uA7T
K4B38lTp9nuMCMrTkFlJY7Je62tX7nHAhu6La94dW7DMHG883xYDmsY3lsBikja2
KZSBp9FF/fGKJJ680olmDoDOEwLED+0rKqHlnEsIClhngWsZEniFYhgiuoYI+bo9
1ZM4jr9rdfMZ9uF2G6l/FdBUcF+QrteUCsd4pI7JQG9UC/yp/SuYik+py9lUCBov
EmDcXpMNhnKrsl7p3DXIOqCOQJ6QwUU/1khgt5NK94ryNy4u+JRuSUbdSIrftSlK
hBQsnnybmsV06Tfi2dMBWDP05rx29JJap4j0SDit9QspFU3yb3exsi6f+ufN/1pH
TovP7mBUUa/z55eW2npQh4a8MRHEXlQkYRp6zPwzweJ09r3L5U4n3EI3UPWQUs1Y
7J2cyvP4KYpVeaTwQRCyzUwJaWLEVOlvbdp+/J02SD1AvBVLJKCshdZwc0SNyJg/
XNY3tMbyT4iwRNsvxWaF37uoNaK64/blq3Qg54qjQ2YkiRFJswDtuyUNeCX2HIAQ
HNh0pYcpoJYzeYVQuXDja0K07DEr7N/b1AqZX+CXQnkb0jOUmZOQ1cfpE7hKrJIP
PyvyUGvXMxXmMugq4H71RpFOt5Z1A92BnIeSGOhGSNHs9REyL/mn5YUDMNT7Qrli
BpULcr0m7QwwuYrrVi6m6bgfls5+uYRuRC1jO5hhSZftzxcV/PxJJDN2ujyKPHd0
NjVLt+TSc0VRNZMvYPSOBokTOEEJO/4jRqlCgTyVSj5erzpHXGHJGQ/cRl8B5kVn
EYCwtvJ40N3GogKiK434YzaEmOxEfgQU8OGl47jQNbfUkIvnNdC7sOdJZf/GTAzW
SlZyoX1+xUBtToDlfzxrzmCwTXjai+P63+mLZeo5eOI60O+8B9mV4fKMSYLFOaeB
Knzdgwzr9Ztb9O+PMKiJwo8AkDsbJrqs1S2A38iRaqs+sqesiDdzORgMxWFMZbAR
8W+wy0JuSg+ezqnjCNqdEwskYSTpKTgPp0xji5egHJCK/tOse+Sjgsjv9h2Fe/PL
hyHsZB/yQBcHdUEG4T2Ec1NmOZjFeiv0jXxTN5w+vRkhNjht3EikpoKBzHOVm2OX
XfTgxONvgQdG/UMXm31cRCR0irN6bQri8hbF1nvYpRewC9VvrElFX28rWBtuz4On
XIiR91IVli7S2tHp16HeZa92ygx7xFO9RVV9mQfH9aJF9tuMblK9nsy6KTwH6N42
UH38UwG0XYS0X5otLcydS5CkYYmNM7mkRIzeDSj2E8gLNmaV2/Y4VaWI9ckxEj4H
L/HWPIq+fkDj6e5yGbc8vUjEARHVIDPpXdCdxtAQTLY/5cG3G5B7klQjNBuJoR93
/uGauOg1c2d3kAg4n1uSlrWmgFLg/j42y8CiekMuBfp9U/5oVVHr0l5X0tlh95Lv
EZkfpnYYvW7VxdoOSeHIhj2Rf9aBkJWdJpzHIoa1iTycRnAQBrJY/rMFhywIQhqG
Ep5fI/12N2DyqaXtMnl8vFVKLPuJaFjAd7FdgnAID8uX+KGLVEBWnc0Cm8MOFCa3
/SKdm2WfGq6DpJWz27zr0ICh4CwXRxFON8RnMEYBf5+JE2uTn4eg5jsIf09B8HFP
zuTRYw6xjTsAKdFJ/1ff7kXhmG9DRSr9GqSRFMdeWpejXjJB3MW4qu/q31FXxb+k
1E9VDhRiDzgR48FC6NZmJduCyuBXAAYa0NIVpAewo10958yQ1/Dl80PC+A9XhQdf
36j2IelmmbS10EHJgMfRfUlaaTIbuEnNPPTWJZmC/9M3h1x5mp1xsi4h6EuhT8in
dSmZ8IS1wSIzaIRzeU5zrA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Uw9bXwyEaLUGd+9nO36gfLy36mlyvqoFdKw3fys8NtU/gLziRXiQieF0COMHo5k3
4/cuEmemQOY1pnYu5OAmdMu02S5lg38C2VgCAK6EPR1cnQPB+Cot6Ht1aaDeb6Dj
YPJMX1WsqxxIE2/M3tFn7yuPHc57UTO2mAg0XRvO3TezWakotcTF2cvmUTuX3zdo
Q4pOcVMQ5rKPVV58wllp5Y4GEuQiYFwrHZwr0h762rguvhoSAVgOabSVz1Mc/8mR
7dglODnAZQv7yqdGuRhuJqXNG9fMR2hUBEOgbZN+7GiuWuzbbx3XNutU+xKHl0hx
iCdZ3BqI3/NUA9MStvhHdA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8416 )
`pragma protect data_block
D0BlfkMTm9Vfb9RfG+MvwrnpzP/2uTRVWXjVoasuI9tyXxx0TAFOsjVt/4PhWu0l
N8XszV7+8e38gplAS+du3gG0TAyD0EP5uCOcquTmE/xuf/YX+vphOCzOdvh2AELu
HB9UUL1ekWpEx7DSFSYnyYDAaP7IKPxx/SPNs4l1q5rsPQMRUNHgj0kl/CmBJe3G
MUyeZnkD9T/zAqmK2PlCVpGhlrjPec++f4yvwGBOZZ1Z/f4vrIJUwIihYcVkml3D
ipXF+KXkdiBuNzSck2oTHmVcSAKe8zVt2mMfX56A2YeTP7wdeU73q/RMJ2EyB0Pn
Chx//wIDPgwaU3XJRRWOqUoUFJ93KQwZTHCC71CHxvGjSSAwWqiOnHQijC2U+8He
zwzn7cE1qa9Gci/VRauU3xkAyL774g5qHHk7r6DULT9+IrQqKSY+UEpP2V9fY2Nj
yOfgyAi1fj9RaHFcDKENiGHnQfEINYgoppFrv+TZXdEOos1eX6ydqp6nL5M0Ha2N
IWRtsKnyj7xfbaXAqPG70BYq/jXE2kpgxiNKPsw5PW6LSRGXLUwXtmMA2O+crJan
YTGTFpxKT63huNWssfjcGhmYwzqATJFbi6yA+VkMELDSUxYIkJaCV1+HamuXcNPP
z90rSQBvE0xUA7Bb9Dc1NsR8tpZxIy492ZOuh+2eDGF62pu6KKTjewpYgwejC1Ds
J1ZPXSRIxtNkcvwzPA+4slPtASABAlGpoJUcU/74BkA6V9ASXSVv/imw0spKHpZu
ryTP5CiYCtE5jIl3yAj5cBk7V76Z+2eMvMTFkKQqHEtDNwadOxPfBKv/xzc4fbSv
qG4aKT9nM7IHuWSeXLFfKZH2AeiznV5maxajtkqEOguv77r2Udn3tbczPhIDrtJ9
V9BqLHyFpFIBZVqAcy4NVoSCcfB0GvV7Y+o8th7P9ot5KpYQK6fD3v+RWozoJ3xP
DJUN52gTXUttVSGLs4kp2xs3yYQqDWybpmvBkYdb/vF9vVZixZJXmPUhbSpJFHtT
TUdvuQ1hE2/MtiUTemmZUKJ4oggqCWpTSmz+N5vlqEJRwC1fcAljNfs2Yz3P/lPF
9SVT3ESIsdwSF7cbxF/bsyNOc1L4Qhfq9eMzULVHfkqOuHwRHQqcu4FTVCc9iWnZ
pI/FIONVGXm5ohnDSzI1sh6IxOGfFKJD8IF4bbJHDHTmmcUkCuQtf5REgeJaxmHF
Jd7rwNcD8GkwVdbFPZtsyT+myRHYvY6qHj/bQxTCg8zA2PBAu88sW5a9MLGt79uZ
1jeq+W+BFPv3AWtujjbOD5u6rSqHar7oetjY50GYY/z6IQJ6HnqgRfslJYeNcegF
JEL9ACopN8B8lraSfThtO8VtUaiG2L67KZKp+QuA9cw6dMCxCwzeB7CUvXFk9z05
gr1irMzHPzJySQXNngCIW7VzL/gtMDrnJscQAwuIw60LqtIj8R8RQL1s7oFwy9dO
+mzBdR7AbBOGL54TGfTvh8r5VplAYvuBAW6DsY4zVqYqHH4DUZyoD5J82z6dFpw2
asWfEzwFtwwX9NGlvejmbjqsdV+up7rDgv3AI+eIaTHht8e6XAM9PsL3HdiMht1N
SpBCt6BhsmP4jP0WOIV+5CItSM2kHkDY6HxDnMyjqr7inebKsC2R711o7DKwxSoN
WNT3207RWSF95emkN7oAbhToxD5Jr1CRzVZ9c3/MuV6c9KgTIyQCCWIJgfFLYQZe
Q6rfHRGKhjmYJ5Ft9wm96WW0602mMabCxqigw30xfTXqmB5XOKbNTFg+kubhZp/y
s4mG0EW7FiF0X5DYa+r5WIotTJ4jcy055pZcBKzKDywgy9QBO7Pv3H62PBi3dncv
GUlArHhGMR8338CnGn+Vp9dYKX2F11FAbekUgSyPaVC7+hPVkS77tkenJ4ATz5eA
+qCwFly4ykHUsgB5iSF7Nl+BczWW4a+zk/DAlZj/Wagv52Zv99VrWPixy7v16sGK
XoVMqsjpIpGPMDGY2w3yryAGymewmUPvT6fKu4FUkOA+XwlKuamY1oDLk5fMkBv+
B2mZQY0uD+ibVFmozGjVX4fnr7OY+64YXlcxLys3ZoUgwCdtdSMHAtIZAWzyrq/5
3low07uAP/cokT+6zl2iLrUGkTGbu1nzO6CZz5R5wMNySV8Hsc02uavVlUaz3uCJ
PCSa2WJGne2TX9hTNgxRk7QS2YPY0mVtJ0XpEK1ZoI9laWrpE4+pDwgQxSR+ocSn
WcyDmmawJ+3/tAjTEGSo6VCyVkWi3Z9t86nzpWU9ZMnGdL11LsRRL7UEDhTc7Dva
XkrF8DYib7zmDbHK2KEJaJFz7G7Fkuzp4GyVd5qHd00FkcRi74zfzjw/NKygpGcO
5Cs2UyuDCxvVV3JLeYaHA4Zh9lXsHtWWrBZE5R71YnIT18p5G1CSK/OVSY1FR1Kc
9trT2o5mWIXuZpxAtTm3lCyl5cdJ2C0WXzBb1gBWKLUkG9jlaLaMsgCtLFUWsPjh
3DXtFijm+eYDTriSUrX4tNBHBTbwt/hw72Tw66MeyIGYbNNYurzJlj/jT6XxHjb3
oDs5U/tlLa4FjLnj0P03SSOMhn8dGeQNXhKfbYQteyoFqgbBJ/2Nc1ar/tkSw6/e
Ug/DQ8110e4RFo0hGp2EE5wS64Aqr8GtfN/O+OQFfnrMZ8K3JxjIUY++qUMp7nGO
CWCZ5OAZFzCRlEvrqDAW7WQ9QJXbVJC8ijpwF0Y/ungkpwM9bEmpRT7pO6aLtEEd
TaBE2kFU7ws+m95JcMCAuFfnUQBMtMaxJAYv/JQRIDAHP8MqHwHdZ3P5hYZ6qJ6W
Otf5PZZlXdX6f9ffVMRgTNZNJD5w0dJ4drMO8qtm4UfcEcgcfMPEMHatm4ImYz6D
OBZ/Med+36lnC6/3e4atFPM8hwoBtsDUlwc1P40Y884DnVr3y6BeeteWpqN59iMO
vQgbzt97fRdazkTMxkPIvbJOwPcowR9ewzvsi8vGEqJ8GTPpQQ/t/z5iuhktQ0W2
TiItynS4qtj/8236446SaLBNYR9s6EY2fSvT1xoTv9aepEk9UlUmauiUXAYIRj3r
kLSojm8jYg69mFlSfQdgSwSj/YqRMK9qfIppUinBgDQcP3a1J7Q+FohkML7tPuyU
EUdOcG7vcmSi3rXeFm8UuOY4Pi6W4G4WeSFOsU85AhB0WZCdpCgefKpnA7J4uXWc
NFHf1FagbGqHWGleF3OK83qCMzZDbvDaQU93gwn0x//wgbc6baVxrLJyV8J73Jp3
m8M5o9s72gloVXHYsfmDWgjCCIztvpeH6B/Q+mNVgf2Oxoab5y1qb1sBvmeAO2iB
8ksVTHe/r7L/0x49ixxbl25afiiK225/GRqQjAapA4zGaLOZsrIqNIz0VrEprdLD
yx5d9vMqqzeLPPnFvw1WOmyqlRlTM4529C7qyGphqAb7QJuglEIuge/2PQqOLkZW
kSNtjTtuHz6BK85i44TT6Jp+ObQEO6W/6daMigg8yPrtyQr33XrCYwiaLRvZVbF2
Q0HK+nn+f+4jLMzdZ0IfYt7vj4Qkm1bb1XZbwe3anQOX3x/ykf2i0bqc7uScKbwv
u9J9VbV/skPiwB8aw+sBqsqU5yuuiDzJQNONTDT7TA08awb9YGBKhGnz/hH78164
KSAd7fuvlSrEWhbs/ahYZdglibTqHt0MzEG3lDDyjoCZBGKp3UUJea85XdxqxiUi
E4Z93XblhWWpD6QlA4MJGsyqtKb49xLE9p+bKfI0qYlpza0yCjjhaN9r1N8QCkGb
CMWQm7C+9HD4l4zh62ZFQc29FeOQiIFr7R/UthGWGZBNljIRsd9zfl3w+3P18jGX
DXy21eb8SUHFJpDbAZVrFvji95zuZ7D+MDn9ogYZW7YOAj80zJqkRaBPKXDssb/J
CR+tsHN4kf3UZnF/Egjf/CJic0JI2rGwc5kBTatisSU1sZDzi8qNNemw4PRAspTZ
uGl0Bd+UqBxZkW2cFKmFZ1W2246OAWwcOgSsUearPkuhBIkNodfglmZUsJynoyoO
GWEzDrmpBcRHkvl9yxPoveyv0jWjnJICDJFLLxrOpX/IVKA9YufyFYlaUTXRJwXa
0SV6JcnbQa39rmDkx3b9R/Z3hR5HHxRhKCxz+qSPPHv963L7rR8075lv2AycBKyt
/KieFeZKC+ov+dUmg2vcErwTXxyVPoeMfEfAHZD9Ck1Qw4oNrRKXZlQ3ivOhJWHY
3JRdTOkUvT9B35iwU/Wisuqv4exYbVEvI1jrq5ad4Dt7Z2FZYH21gRs7dve+Cs5R
3WtQ1U5uHzX7LUCmAbokk0utG4VgeWYhRdC8mKRWjDIa/CKEcI2NVDSiyC8UmiCW
tgYsiPQh7nKDojLEi+oHcwUrPGpeqiOrx8vlJtoSYo8D+xPwtifz4mRW7cQK6Qhz
buD3keLw1CWBsepDl7GN0blThmplVZ2g2xwiRv3WQVRUaBCjfMn67iiwujaPldTf
/mHK093kXGPihS3cnHFbB/RpP7ISx/Pfg1NkYe0u0MXIgubB4/BYsSFULB9QXSrV
iDZTTDrL89+T2ft5qd1GsxS0jUzRiRFoFFv3xvREH5H4+wvrRS8Ayjo1ZvN8o1vW
Jxx5o7jkyXk+fEd0H20HVlOQmwNjX67aNLLFO3/f71o5FR+pBGDN0VqgUJ6qmLb9
FB1zYyHRswO5XWo6gKX5mOobyTu9HViFat5eQgsx2rdPtVzMP7c9FEXZtkLSVdts
VhKFYRULVHWJWuqLJigsrSCEomll/6ajAyAzcsznJDWfYo9rkjLCF5LiMTJg6RRk
ToD/oxahUdKJzU9wmxOx4IY7po2YkOcluesjkRHHYhXtqZj6v/q36gP/Y3pTLMC0
pAu14hCUIghaYBrLKJcKoYNKLTI8AmsvUshu+g1MWSTYb6Y/x7vSKgoF6ivk/oxg
lUmw9nNJ+BEU85kaLi0PK4LIiQrUiLfjzHvPt/dT01a5O/vGO6+vzBx27lpFjTBQ
gL2NAMGKOIfZzEIYHBFTCXm62AsvfyTt16NznSWfQtFNU2ugi1B+8ujb0uOJZ4ec
mUV3EnZY8p51EJawNlRz0dxsjSE7b4HnueYUU/8LO63BbDEJvRUu+QT5zo7zCXgk
xP0TH+siswPfI0l+GxHFLovxnRe9v7fhaMxQ9/4PY72VhAVGjBEAAk/MsLfyBw3k
C2D2BehB8QyGlKuSGzbr2Ci5zAWULm70UuBIEidgLlFcOsp6yPp/nx9wcUCGl1Yy
rzIN0MABJ3un4erGzUS2aZyli8hO7B5HG0iRqYGMjtBanzpx7Z5B79xTyM6js1om
I9tT73gnZe0uZyNHtrkdMrITZ/EGV9tPAKXPD0fxlQ4UsKhGLzOQ/AEu7PEZflVn
yRm6JEajzfd62u2xu7YNRR76KMFE2CfOSI3Yhuo572qpUVnPpt1Uz6ZbeNrDeSvO
K+RzwfKUJjOcxIJ01BblAdNcDpXRFu7HH52HCLjXccGsTX/cqp8lIqhGRcTw/GbO
+pApNV9FMpeP2LiuMJDDe/2It3WbyJKNrVyKj8T8oHIfDPh2gtZ4v88ISibPzAT8
LTZWL/Xoax2snj9D6VY3a2gvhUU3tPyWK9VNUMLqQWWnyZyTd819RvHFlrDMc4aw
2hVOh5DiDP7OPEpAJ2RlG1bDKpHh+7uPUgA2IB1zRZmYi4E/1JRFurcMcHg7vN4+
hc/A0yj+G/frzreKI0nGJeSg4Z5PC8eppfuswgpYBgzwESoQZCikFGtcARzelKRK
EpCj4cttBQXLueelcN5vhYoue2MAgiM6qfZ0b7nuM3aEDucpvBMyB92+MZ4Rk/0M
Wfhm0iAZGVrYYqT/MPTTXGUL31863bPike0AACk1Y9AKmavB7PREkxGc04xDCL4i
NHpKu+cnxHutxJSKq1WZ/hAu8gASSh10ll0eUGtVAvKUJWgN0441+VSVksgxK43W
/BsTx3IRpvM45tqdWtT6/kHPpcJMPYzHEttynR9MKctDM8GBzhabl1DkJTmUeJcz
yuS5vY9PnWK8vpavadMBmSK5z4PiFltmyL5JEaBT9tRdi7pMWOTavyzOAOY2rM1p
TdkgN2MGTOneRUyO13bceoYV8+GQSBHUPcbvks9r21dXZLzPSeELzeE4s/XVkUwy
tU5bpQ59cR54yQrvw2DD8fC0THrJjUV1G6t2jus+AS77uld2TA3jW/zI8amlhZ1q
6Vz1oMnoSgp3QL0B+c4zVa81GqfL4Z1aTfLa2BPFJrLgcFM4MWi1TnlyDoEbxDcP
GFL+RUJ/ay9BNt3x2FxsS8nu9IzVcqwdJOB3KF070yljzJzt4XTVCKC/TODFuqUC
OHzomSvStsNlAa1gBo6ib8dTvNHGn3SbSrGqcKzKKd8VRgS2l2VgSwoVAXvEC9d7
rBwX0J8MRXF1GD5sHQYIxE74BqL3rhY9ol+EjkEK02ELZn9/rLEvg68RFDMftspB
u9Pnb8f68altr4rNtwiQ3Y033Vn5te/I7Rv7tql+48XX395uivTVPOdQsUO3pblJ
uPuG/61XupRECX1jzhJPWIIa+BhrWfZDKLxKeShVdPQb96wgvA7236ykwYW81PsS
CFvfIpabQ41jFblwyWJ0LB4zT4Hl9Li7WiuBQVp+MHSUlVNArlu4JG6tXak9iQjA
R1Tc+AOdFOt2xnSfHyoPrARtFfx+OUKiRpbm29YBhmR+wwQ3cjwmX2E387wBN2/5
JLWleFLy+RNSUXQHA8uo1b6PMxcVdu5o/wmwRRv/Vk9E9LWKTgjiDhKxkXaKtkuj
eVXC9bXeCgJ6K11TVCRlYF3B4XdwX9hB5SlVK0SSyq1WHhGeJ/t0/rQky0MHPIKF
XlgNl1GYF77psJcxUXFO6C8jScdG619xoiKSV4Noi7EJu3wRNzYN16mnNrk8Lv9q
a3DU2HsMEQGE9BD03cvum3bNyPtUAPed1/Gb/563E2HfgArr5a+OwZ+p/OHoWdTS
DGTKWt+xGNpeGZccyoyV+hMRiCc0X4cpNC9aXvINcNVmaqjtVCOllE6GKWouR84P
VEFlDy1Naw7mukKGRFxLiRKRU5QverhFyetbzYSjOkfzJ3NafcqxUSHulFgIFIK+
/KW8/RQZDsafMXY77Fo5/xAzwn4qAkhw0BFSpc3ZetQqn/dfE+APQ7eNNXAeZ1RY
iWHQNqurU0OosjVuv13S+vAVK7O3wQCXBf5oc82/XnQnGxLtjaLrEveAvt7TrB+k
ULnV37LlX/d/lzKjIFzw+yXopZMpGbVUjlc39dC9lxr2h29kgeFasS0F6AK8j8Fe
66KTeUqJ7+RHZCtbrmDd1ls5kzQbSmx4p6qbf9+XzcOoEKH0iYaEInLbyKfew8kl
Cg6kuGDS2fg3ZaMYOV2NdATppy8TdSDiPr9AwBssgwqHt6Toec41qOuS/0eypSzV
/nEnziUYOKZMLlcP6Zqf1ZWFW64eQUG9/3D4FdscZLb9NfuUyvaI6aCuXpIalKRk
1oL2YXMGR6be6sxRkMZ+BodPnazNFu0H2aqr55tynGzIq1gsMZz9rNG84/PhjERi
SptWJq6MBygqz+Ed9FXCSE13cWzDs3ZVMS5H6x8Y74rxdrQsAcbFVptPD3MEMyZS
Gt24+G2fuy2iAmbKJyZxhnUhlqWC88JMQotTfNRLqsoIApIqay0FZ/8evXdgVhkh
ZIAEmnCwk+dUvkinFNJMYKpWTxXbPBE7RU8foRRe9QhSirRd9tdjJjJqEGICMDT8
Sh44Jehlri10gbEreujRY8teosjAxh2rhU61B8UMHJCPAVzRy+8jfupBg/qQIkd9
LVqcYJ6yt/xZulQkWcEb67j8eOShvLULI6dj1F0DvVzTVqzDJ5nStJmZ1NWYMinH
dQFsT9I9/4Xh73iyvtehhHepoodZpmBSVRpLr1ys9n8s1t0sARJyEgmWT2SQn7gz
+oVvw7dioigDIaDtDtj2r8m6rc/Fr+QXMT6S1+xHvrUeBSHK3uQL9GYaG0nQsP4R
Q913H2GdUVNRfxUFc2TXjS9nhQWYTfrznMsMuufuNS5xQMfuPXxRIQJcF3XuNueR
HlUZ6UrypGxUdYwBxiccGXF/LLSHJBjMQVEUYRTOOG7I28evMIGUteYkG3OyPZdF
LbiVg+yJkclsu9MrHLRpbq/CqK0MqYkHD5j0zZYSFVS5YpTc2arzZ3C89df+yRWA
56hnY4MCzlaqrzO6oyzjwgyb7gbv6YLWXJ8JDKsF7YKxYh2NZWqiZtDMCuAjYxVQ
oMv0sDrOYaof6YF20ayzIbiNGk6CHiYP8Wuod6R/krvq9ifz1fT6Hm4Wg3JWSWIe
tiHBYJJunv2Q/eW8x26e3fa99cIqXuJq2ekasuiwSG+o2kd179jbxWylo9YeoiGa
QpzfGC+exZasgm0M9oIOTO38rLkpCaOiUCEGeuG6IqD8DfVUHVUw4e9ok7Im7w0V
wugGn1cNhHCWC2ByLZ3s7I35wGlM89yqcol5t8zsBmB6FBIWDvHyOMxFZLaPPcFg
DOkI8APtHq3kc/lC+opQl8YVNdf2cIpaO/LaesWJxVMr/FYEh7HcE+kxrP2AWHYM
9ta3kXmrX4RksxQylCrPtkwbc88l+h5FPlCYmiQRepT4GjHBEUe/YZ+ftqfV7T/M
68nds/eOKAm+mcpb9lHANnhpB7OGviAdBc9HzvgDTxkvlQtl82g3FOvdXVQZsd3u
3+lHiURRHDFrGuAe29E1z0qQxvpmDa5M81XDgqafhRtV1Sx1oTALwyDSSArCVK1D
O4aiGGICbfAW0y+4hDNSrSh5L+glK8nO93mIIOAvpPVej7FnDWihjs9TlybUoa9j
CAkqaP6Ek8gdwpfPT2NS2Gz2thwzBWnN4LSV5Vp8+958MpdtkyiRKNydtSFVnCfY
1n4GDvPMvY/NfcF4/oy4gEJB8lR5xmkOkM2eNXT4suMGzddM/Oj9lwv75guc0ExF
xtWZGZrdmMq+8+7WPilg+7C0EMcoI5FCDyBJJV/4mvLTcoydmErCnKVi2KUG96Wi
Nha9/ibLQGppkUQqZ+76gNUpRJJgPoLJWLfYBIETaogKzxZ/B191nupJT3cvDEYO
BFSAA+jJdhTbJQd4tCAnLNkLqwl2s2BhA/x9s+4e26CD4CGDX5c74QyPaY0xGHCT
getdgREOKgB/M332Vy/RIx6VGlFsdokw/bwBFxt+pWhCW1z602h8TwgzofjwsrJc
Sy5HRUrhL2KLOb9FIYVVqlh5cWMkgeZLHitlxUnBXWQKVmEFD4pmwTKLsF9z0L+D
hDjrrmqoSyGGH0dqZitthoKd9AXAoGvpEQntLF0pcIM8jSexEL/gDiUmg+RuCtV6
Z2ABd+6Wfy6sKPba4T3EjaUoifxxA2PybY3gSfauAgQadpKK3tzBr/0I9GzIKXeT
DziBPswPJE4jPRCzj0hcSK83GmTKp+5wqDxRy+OVY6SZCX9wIw+hPNOLqNbuKV01
S3XK0M2IsJYbRHYJ8iC9Bd16oYh1qn+KGR6DAJ4TfCh1Q8j0fU2OaygVNJ9EA17p
ung5YpJaqjGtZ40AVP26uSb6cR2PN162qT8jBpPAG6X28nUn9kx1LyoZYVixfBSS
gv79yfT0ErSpgI/WrzlxRYCrPhMlHu4cLI5k0LLWRiB/7+hd/5Z69+U+Bo4tyUA2
xHCsdZ92h0+aDQNoJnJs/ne8v9nbAiYGNLqZQumvHETtpZcoYuV4Rm60B2KzgKDL
Jb5kY5cWjB5w73EnU4dJOQGigoSYkFkAoRUeQ6s9vWGjvpRJYoO/HeOd82BACXlp
lfLO0Zxz7KHm9ZqrG7U59LWUS58RB7TiCWI5c6yEURld5osmyLrrP5OM97l6OR5T
7i9YmxhdPjF+/kpUiOZpz9s+DxVic72udb2DHOPz7OO0ilYhQBvAF4Tiu7emebQW
+jCxf4RXvW7pycaoiMIPPFBFGbr2aMigDUqrnLzQXXTscW9M4zK0qit/ZRx3iWoA
MAeYwbgtx55AqJKWVZnT1dJ7lGl7H7BHGPXTS9Oa/HdBe7paO6f2mr92B4B9WPfR
NBB7wv5KQO6SK77NPyjcSF18hO/0F8WZ3pL8KST+uYKD5UktRkqVWZrxO/0hu5GU
oTabQfpuwM16hgZLl41nS220WYYYxukNNj/7XKy1WszCMPP2N8hxqMmqSizB714H
1y4xoIsEgDAfThzpbjJr6868rlAGZbHK4shbqllN5R2PcCG3jW4IgT75RfY57d/h
J6nvLIvWLODqiuldNo0V06KIbqcWgXNBzVN1NJ/1jXAVHtYG9StF/o+fO++vq18t
+KEpwLWsjzTkX48IK3pHFTL8BgDZcAV6BDeNRm4E1XHvdeinnsPWBaeH2ESCQuq0
t6N9P7lKsnzdH/yfTKcvHKt3roO+Pd2UjEFdl4STufxxhCiMSuGCe3rtCGFYySci
zwrvwtDop+Zng1LQZXV1vW4ZgaUrMQinsp1WvgqHVROMEXYU9iczstgprLlUuY+L
/wNuCHMszj+weKo3oTRV1v/pTQEaXVVbAwoeJnYVfnDPAcL6qviRr7fs5VJGSKdF
Lh1T1w+9Ys/rFyL0UwIF5EDK7B48/rMAZCvMJJCSjWxvzttSiNBfCyzQjgegvCJO
+mFiIBbi/qHg8vKzHkY70eIRD0FpOfvybBn81ut1JI1O5A13mDy8tK98jTlq1XUD
hypSAGxfK/Ex/5tl8Bi2x1z8nv4Yu5mARt5RwRO40cyoqVmLs14847I8qs2MD1Ds
ONCeg0ImQGJHlX9j5WN4wD8ECC+7jbe2a3nFAJu3qGL/EkMRp7NVNd6hXkv9TQy2
ZHNKcG1E2k+mD1eGBPljhoKx068QT/RnNS/1yZ9u6QwuCRYh8Cw8Vv1pu2ZEMPqG
nZBKHx0sbeNY3b/ogV9eK/ZEzHlGqc9+rXhMT4iWLDdJ/32LWQzlamzA0U0xr12l
8V7M780q2hVUNEcRozj9Qx3VTg68yqz1duy54OjyH3DzC+8YeJefzmHJWTRgn9nK
k2pNX3vmOJejr5IF3TPFxyEyEsxK4+kealUHZDbpLCm2ZOCMTQa5S+TkbFZcw3Ra
XvkLYpSu2nY913zcle2z6VrhCCYdtJy7rpxu1OQph2Qvs1L2QHJPIeACx1/2fk3U
7Nx4qjNET3k96KO0B47uTApttWoDJ/9iuBGDbMdrUOI/xePA8zrskRT1uk2Dpmxn
gBDfCGYkTdblQifyvPrLyQ==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hPQqFSQa/mRXEPV/HOnoVzycrnLZ0liw8++yRODGF8mEOusrUxgtvxHY+WmV+9+d
1ShRzST+NVQSakKfzI/2I6jzc2hFF/ENOqtoGD8lE1v39xQbz5pmo7RUeKF+3Jsr
j0x8liUrMk4nibimUIhx+yBuFOKaF/pQYZ6k2rVFU4vRTF5dHuaaRzXJdvjC3kET
Y8Za4VSVjt0la0yj6RnDleyfX25n3YpU6oHJLs4gjGXlrh5GprHyRfqpqevegJMp
MpQfVl4yfPsxfAkFZWnH6po7rIylCdlwtWi71zbTMidA5o7qAaU2PZY9LnukqitA
SAx+Y8THLL+X6zJ5M1+Ycg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 27200 )
`pragma protect data_block
iY+u8QQK1rQ+vRC4OVxXrSCuBecClFt0gdn9S9SAY4m4Mr/jhv5SdbMkTzCRuHk+
20XQxbPK3YS257daBAomnsvm1/fa9UaGdygs54pIf0BYzBKC7h46eYcRRhgkgb1t
Fr83nxOnY57vVdx82hykdCT+bfAlrEwTM2JedHWXNrcRNW2e50STq0ofPrnDPOgA
XCMP9zAmpqyWkIuc0Qd8lfizVOgQjHL/nGNyUDSHX62XEGIIzsNTL00xsUmfd6Yb
w2GCw8sKyqD7sH4kEpaj7rxGahcTzB2lTYz7I+YkYIL5iWgirW805wpdqm46w8mu
7IHc6PiU4PdWUFWh2tHWm6b82fmneXb28R8YwNQiatfsW29ScXTyF0ub50craBz0
9zWqRzPyKnTXy1meGA5CG7jpvoq5mZWuxc54mb5wVQGM2ZLZVK5X+f+wQgQ2UJoj
Et9Lu613NwweeEwLNR/uWne6e01Iv/C3N+rdzq5JY75OgJYsP0lkfjs7BxBROrk9
G5hlscS9LTgEi+Q6IWUfLQvgkM1UvzVBfRVvu7Nn26nXihy2+taszgjtUoZm/JFi
dYoqAs+t0Ai5ajs73KtRLBRjJLRcubwS2heomn6I3uqMYTV/hd7LmvEl2vG1YGms
wEEvmuUwM3Dw//BXI5wuOdpupR5VS+cmIEdN67t818O7nr2AaE2so+dMlwUz4RMf
xEWagvojQxPfgI7VYPw2AgbXRia4EjUuoF4guhS5nbUrcWaEo5kVgn/jy6YNYf2l
VilAP0vAyeRxMxD4pjT0I7ZgWWJ8ghWFaRW074VLNUA5NxBF/WGuhFakvMJuIopo
ZhKIOnxDbe7N17lZup1AGAYahyQjGtkg+gbKu/nO0/1Pb9qFW2Abg4546VGcxVQU
yjw48ug152YAsuyxBEX4fXwU7AiFOtMl/HYYLE73Ktu9uwS7Hw3+uWzY/8/3Aus6
cbi02D9dGd1IFRPnzOS6KIQEB92ZumKCCJyu0PPe98tiLNE285mzNQbr2d2UrESS
RUNR0nuFHBewakqLHMKtbRA9cnO6C2nlx55fQFAlnqBa1fehQ4wxcBiscDtfAF+2
77IN4t6wP4u2QyRrvfl+ocGDsG+ahCupcIrnBIxCAAtA0oJ99SGVeuRm55FP+Xj1
CAHqlTpK9arsDZfWYiRhcOcGu4rvgYYGbRdOKPAGnNRpXTDT6GX6wTseglnM4aYT
wKxs8ja1x/HC7ZMZbeZ/U02KVN2DSxzEzKt6EjzUrUy2pGNI3kqWgqM0KylEIs0M
1bWhGJ6pu5qRCiGHwscN3gwJnbh1gXn1cVwH2z/EiX0MhY96abbXEUjxg7kBv3A0
g3zEidgCNxSbkhgPAu37kxbcsfbCeKslpZOXT7rUyE+l09HNTkFrMMvj30HXOd2V
3PiFQqCHqKn/2vSmtxJwbL+A7CUz2/4UJ8qkluG1kD02diqF4GZGIh6GrP0r4/B4
JoaVhXRdGL8jKGyJuisT36nIgYliIDRrJrguUVC6EabRI/fRKjJVGeIEXv6IsWoX
BNkH4mlXAUslbfEAzYexbXOO1P662QOJS84gUO+VfPFjHgBsyBrLYuWmgHOmLtCP
EZmFXjHtSqO1Pfn8qVdLueDKyI75MItPDK0nxTeFi3/2KL14bGxGNkoB8R0KACgj
dnkIyASDyKsXs5vybZ+ztdfHxFBtYNzZ7EBLfUvgaXyesWj7StsIxbUGe25Zkrx9
cGdg9okYUzs2rYne3IU39boFqv3jACwJy/mgEMvARKLyY18wLUVx5trJ9vBei5D6
TIMGw5NInlBI0HBagCHm9aFCp+xfzT0CpgS4k4J2kdRK38Z8m1p0bD+rQIBAVB+n
JNtbzvveNQ/zh9KOgRO4zFS0e1saTRx/lLYpWWnUYEjQD/cX98jxVvpQkwYpUSfO
4hdkVghu/hPvZY4w5LpSIGQeMgyDYZA4aB6w0hOl2nzRkFj5djciokjV33PcFZ0C
LEVmRZe9UdUecE0dyRmYKLx3S3Gh4xE5W8fIUr/Chdq5tijM9kOOiK0mJ6jbfBBL
TlSdqSkpePHkVFrfXe3phUT4n363WtwR8clcuL69plax9uy86SaotC76USH9oFdx
W67DYMC+KrYieFJ/TbhdYS+8rPuSqG/+VBvAbhoYrvbqnD0AZpebhlCiK+C4U6y5
hZI0RZmbmiBOKZHEQtTmVVSI0Emcxiie1CuhFWh8rL2p95likliHevduGCzwIUr5
T8yWERLNy4rFpKWd2mwxgYg3di1KrHUUwQONXDObGi0Ntt1Bk7mpnl1IiFoPA8Xk
+cyEc5KxQzCV4D9WA3CxojMfWZ9u8hCvKfVe6USBOhs4C7+BP9f0mMu/pE6q3LX2
Ks+uzv7XhyanASStAt9rX2Os0j1eVltFVLDc53eUidfWtg/dEn0WLk4h/aTaF6/z
Oz7Ddu3X3xn5SDLlJjzslQkTgBbTlhTehyzXtTAb2gv8msoikshi1h1FUIBsjyCC
5BOspa454E6Z7ZFunZ5CbMFQAx+wAoT0woObfJcGfcpUNY2NKMDhG+TSAo+lZEB7
/QpPXUHDWG7+B98dkC2ibj+C7nzIBhHOslteR3HYl2IlabZnBuAYVB5TRXvyPtM1
FRbxrSLHBz4739LOO1QYsNYK+W5T3XXQnpKawNOka/0JXii/YKoTNXMg0yU71T13
5K80dDW4wDEbiyMCxBYCwhtVV+tHoJpDutN/nXToFodHqTTkjBJk7FtUiuqpzVLe
Uv6xSRvocaIr5yiJLXCPkvMvE9CzSnvXP61HyUL7yM4SvHgwxCIo4bTYaAp51kpx
GJ/mhXjZG4nF2Gy+/c+o5JVI3KQ8A8swPB4yxsaGWA2wYdza2NLrndab25+lAaVZ
Y41rHVQhG8kcIabV6o9G/4/wVu44+DBnaqZKEwEuR1byiShGJmVK6+6YKd97LzWA
8GhkFDYx8cKLbODojqlZM89r+58oSQwMT1trzxJhhcY6YCAOXXVrawZbELZ2gldS
4oDac1DilztP3fEYYy77h9kvXk/ms7t9ADIsGqiAFwu5K7ER4daNJOHjq+g0MGid
WhV9CwdhsgghMGGXKSfZaVmgZzx2t7JrfoATm4DBqReowf9hASIFRvExsvpQKR8q
T+aWPf1Eox/RunhQYvltZ6lYOPSjnsvLjZMvn5ALHm8CLEqFdw/t9l3kN6bF1oeR
HYHavuoOfgCIqWfxn6p/oAlI2pyVklK5nEce/B56qcAEiwzAbuK5mtcfeUgP0JD2
saReRM780xIjR/SbrMiMTnyC12UnWolByVkHRGUaaxQcvFTwbvG3mWH+rP/QG++b
qHHNCv3nOvPFESnF/pz9FPNMDMeuruBqX1TfYZ0UNng8NNsNRAtDhG38PKXqwFwC
ExDlwkpxV3prBG/Ts9W97rsB0q3lZlA721nZ6cxrOXLegSgWvifpBY4jB3QDuk7I
Z9tyLs5RF991MYBdsFcycF5NnUysYfd2mWODy7qTlmDePR83KWbLq29gqPB3Eu+9
jNKpIU6yxCwSh68KnQLMBz3lQz+k6/P2IdEXMFZB1N7vjcnZH4zdRTCfQr6dsE6k
G0L7XBQEDmJe55B+xmlU4w+PP/vhCXq6Md/1PJBYX0qyPuNVmLYunJIXunQ6TRvc
RyxEd6ZWiLxPojuPF+L20Zz0o7G68a/BP5utXqZgR9JhkKAZGPXmqDGf1jcmzbNS
rSuFrrmMFtmh7Uz4cydHOS8KM7WpEOWOBYdHH2uvGyAr8ihnopgGBj9uJkXnD01A
Lxvm5yQuLpHlslbAIVQkxVk3M+Kp3yyX2DL3hh5ddmYGVyT7edFwJ4FfQXzYK9uE
Ilrd2YgzL2Amo+KujiAS9/NasOQJ0cVReja8SMHaB0Gt/tca7oRcZFk0CYfFD8nT
IOs9ETZyt0OTqbiM5XpiYkcDr1pQgQSTQw/cx1awbwUwKQBTI2L54Q6OiKPJd74S
r4Du1l8UUiSp/MWIiSiU0otJDEn+WvEl9vijsfW94VlhxLspaEUYNzEUlPOXKXAb
cEfnr0xwFuBXklGzWKmZyLm1uShGn5+UK4USq4Ra+UnG2cNOJetyaBBB+Yi9kkfP
vRheaVgAlD4SM7pXOTFOTfzSZcEkz7igKQ5StZzO/YV+9Cf8OLCZB1aoNODdU2Fr
VQP7j0Gr2rTrjT+aBiTXRGeoPBxoJYcUoHYDBjpAU3cONrdA8uljuDcalw5AUmSU
T376Jn2bVWvTY7FqALZaA0cP4/qREs9zGZQmoMz1BB2I47LQt2AeQmCW5DgFGB67
bq75UZWFGGoYhG9vzHtrekcoupG08ZsMcIqy8k4iW3Db8nSu12gC/Pg2ghs6EHEw
95WEiWpDBsBzTys3vtaqFHeQPWLhTJCgxzPwABx8QqzkZEVvyY+uQqoG4+Jgsqiu
6wVI2RUCMVlVW9jPL5q9dxMYusivrF1kBYg09CGupqFqtYuCSP4JNbXFjk3wdCzO
XXRjMuSbOSGW1l7hlzZTmCKmPwokd+AogCPZbigO7MFWX/CryctSoB3az3oo2RF3
f+HXl7X0AK1pbb9NpuZH8ukY1mzrS7WNpT+/yGLAvciwzBg2uJPdxLCjHyNpE1/U
D2J96CvYfoXFYEH1WtOU+7LqNvji+d0mcG+jK3c3uEdAJsG19TwDqWopfivpMZdw
icPnCsAne1wMCP6DxqwTCNpV4VnIShRBHSfi3CZ8bAK7DDNkF41dB+YPuS64IqG7
Fcj/0jD8Ova0bMUPgFNGoYXynsJqcizAyJQSKYm7+qYCwuG5i7YCLOuhFTLIZ37B
L/klsQXOOV/eOo5ReD243oJ+zvX36VYg9YQCZ5flJgw/08ctIbgdKyHTBlNoDylA
nZ0mdsa0ETeIvNoSGJFvv8ddZGopm8daQfGvP36ii8MWXtlnv1cQM0qntUNbn++c
IJn9i9Rp78whqeNSAB3Os6HH1iDrXRExuO1T0Gtn7wFXaWIeEKjp+3HZuA9aVaGd
fUchDD6Zfht1kDqDvCCF5/ujUzujJ+b4eKjXoTTn5QEdYabb9c+WO6skAbgzKaDc
n7slj9FCMnskr6tm3LCTBO2GuHkXoEhdo1MjDJ6rULZwbU1wl4ARd16bVeSbd5Y4
0YpNNiWkdW4KSxBX4TSmjOvld3Zc5IMnnlXl5k27hm3UGbYn4uWy8Vy8/GVCFjS2
uin0MHuBxY7ed5Ynz09NYcPJ+WN0/ZzlJc5MUXfrO3m2B0xKG0kY4tjSZKZm6UlZ
B/ca9EoQ2f6WeVUtBI1wPYKegFjZHDY5kQyCuOTwVVZKqujVaO8FdbCBHb1dNzOc
KGWK5mpOTzMd6oxkrkRv7sJVO5L9lsrdnYdP5ALnsiSUeIk7uguBLQIx5fxLGxNx
6jnGNm0SFMkD0t4Q0SOMCuNzJAiY4jKR5UGf6T54VFEClBwai/08MPGcOVjA+e33
udEqheKdrMq7LA6WOaOOqsKAIcQ7mDzFdJL8GIsq3gknRz5gvTiRbN8kWGboPcbL
XLM23tOxobXJwycpHhfxMMuwANmDkaIiwhHHZLRaqanRIBEnJveaVCNiB4ZWA7bB
BqXtdQZ84LMR9245g0jUi9A3XVjwoc5Hyx4KD+tAoCw4GabU68TKOHmjy8bdrrh3
wmCuVQjw1WrPWuDfoP5O6K/jyeltbp9G82m2K+csr1b2kzMUBJyTbLQZ9osy4GcY
/ASnDk9rstSAQlNYpTx+pM5BUCiFkpdM26SQHrgRmoUGxQn8IfT9kXk+cY5tNnO6
/fb5QOOtKbYJIL+o0ZvGqlfe8gZEe3fqdol+nowZqABpcbD5UgHuIPhE156e7xIG
FEdH1CLTI4Z+EvzlzGUocOEMP44O0pgIBaIuJ3yzyLQIxoLqBR3eVD1KUTVokdpv
LDaq3pS51giH2Ph9cX+uiq1qjWk7rxp16LMgyH/CEeSznzkfIaaUChTa/kDSNhIg
MACBgXEQXoMXbJyOcCPn4GvIPgoQ6OiVvv2e++pm1y5F7hvSEqP5sWhWwjJ9FRTD
mt2JGMWl8n560FUS1Atfejxbj43D1cr55Fcf9OyXh2a6aeEraEL02oWLdjdmesSG
IN2KuIZ0B2cJ4rVnr5LZV/yCftUzNcpUUObgUOeVH+apDc8LJvQyxj+PtJ1hZY0y
7aA6FoDN44vwEEdvtXPgIqW/IQqSfLDAgseq2Qwg7lNRcgaEVH/sYieV5ChKcz6E
F6cnGjhi29mOoHyIUv1s6qQg1e4Y+I0TiBgYJt/C+ruWugtKs9FcIwbouTu4Eyuc
RThfWbo3FRti0ABOrYAzQvm95lUFWEgm9WJiZsxQdPnEctLcFCLE7O7UA+rsGbBu
fG7lMQuh5Qkh6hFpeOYYvM1YsLzMpEJbjdODa+wkuhEWUCC7JtmZioX+uJYtQ7qS
IWdkR9JEAlaWD2j9EnfhT4UAcSkvtplu7JEPo5hC30FTylBRCDlsRXULiVMPHelA
Jxc9vyvtr4hgqxEWCTyEs/owjUdNehFYID7pgZ27Y0aRR1rB2g/VY9kNtzDMnGnz
Z4SfzyYVFosUBOG/VsGSHPbh2kIDcPSbh1nLX5OvFGpC4I1HVqWnmB5C8HbukJhV
qCGG1klqGIioqXx/Q/lnbObldPazEXr9eDzdcGpMtgKUrFU/G30IlMRH9KpMkbzN
nIUGKWlyKbEdYVc03aym2D/od3BMGTl0pYveap9noPMY6DmksGzmZGBeMFCqAA+U
ZcqkEeWxvzL8f7482iYKeZs5dj4PmyIzgzkCheuvg4xpjyLNp3b6SC4zmWeYrgWu
+6Pm2MFgsr73WAy0cnahABinPJ5VTkPq05ydaU2MClwQtDgYE2HGL8q9/+k2QTeP
gZYKJ2Fin+9bM/KepuVMyDlfedEZQe6YAFm3GNL4ersvV5edjs74SW3MymWOb/mx
n8gos8EaWxSVvHw1fSojnsqdWdibCOs96QW6+jvAVAnx8jTleeyYDSucMgANHpk8
938vD+b9Mj6301pFuezR7hATuiemiABS6Hqdn2N6UaVxqnhsOyyC336Mbdde2DDR
cp8dc+VCgEnKPPA2Bw5ML6TiLeXRqi6znDT31V/XXkGxahK8tvuBpGMC5HJFXiTn
noIKYbw7HRtaVIm7cWImZ2HJerf+kdOS3GN5VhrBy9yfT1aa8vR4/Lw/0ZS4KmhT
jnrh9ZbB07jslEBmB8iPYwnAjHKlDqZ/7i3bm8KozfNj/L6Zto7uTvwp6UG97YKV
mwEEGYzRbEWfUZ8aj3Zfr0inM8fzUvmKfRIAwoD/HeFmgPCKIw1lkzANfObqnuuT
jhb+iOcditV6/ogdCh6TvGznCmlOOeQRc2ZGVYWb2dA6WxPOcHuJer3wSXtb1weU
cGRMNhUZm3lSBMhQ7TnuzI053WGUJW1+t/WFXtV5+ZF/ZfP77UkxGsH1/E0Ezs2A
MDvwP/WXcsEaCb4zOZUvx6WT+bNeWwwDzKZAflmRXuVYzJoZ4hDYo2xWfpuPZNHF
jsHwPZVPX8nqGU9OUf/ADzjhhv6PXPI+bLSuxwrkcODgwZR78gJ0Bcuc3G2PM+wh
+09ozKe4rnU0+2uh9uZWr8qdVNA6VE/pPWn6T5AwnWBLlZvVbbSd0y40sIReS1BS
z4lgf1aIOY+si/z1hNnQdKjx8D47nDQVWXL0ylw4fhcmCYUUug/zN1uWfm4sNCFZ
N9M7LHECaNGW2KPBijm4N4d18dpBAUFrZF81xoSuwLoDZ8150hdNlYaUo1RW9Fx+
FB+vJE07QCurSXAfeVHb/mrN3GVM2DYrjbD8JvSq7WjhNkHFvwiHvDeU8ZrNeemX
89foDlJT/sZk0Ejgd8Dkjx5upT8ATMgo7rdOzSzDFdImcrdlYpX/9/D3THNJsy0i
HDMTv+sJCadQAtlCDnXlap7i9j1lBW0dYuEUxvvhEN1SJYzHbMg4xzxHaqkIY9Kz
y2nMXqZjYFDU2G62jmSr7fa4Ka4okSF8rJI9iC8MscuYrUttBUJHMo7VIGVDreLw
eKEiGkaLlZ1i5zAwFtZmUgPHE52Vy13/7FtkoYT+z/kBCfcgiXwGePEZ8pfT7Nty
hJdigN+fFXUh3ejdZvci40pueek2qOqZUtpb7nfSdn5cGG0JS+RY2P+qJzqSszhC
s9OvYtbQEgrTN7PtnFbmNMzNvWKMOPO6TW3Dwh0d+vJewEKl4f3snNYHkN1DmEv7
Rm2J9vW7jFR+QeqArMUL+lvO0U9of8GFD56XpNF94nBTEae/YvS2S3lZI7JR3cNw
Guggj2MAY+GKRtX742uW9tNKr7LQTDagxpNhceJ58EZUpOF7LH3XOc24BC3S8yPv
o+KTQRFOQuzersj2kXUE155x1qXXEjTzN6NUwaH8eXZTn4eRyDZj4vpKeCUN70Be
KuY3wkLaTk74sSsMACATY5fLDC/FDN4hP/ZK33efLID5OXbAGNUoKF4CBmwbgG0l
AZYNQuyg3tEiYvOXDghQZppXWMvXlItFGvDNIZOvMuiAU2pECkVv5Qo6pXCaLOEC
VjND0JXrwKpNX1Qiw4RLs+DHKSMv3YUbHtlfWNRntJsTcqaRxRdpJZvWS7gu1ksu
vCIMJwEpi3qhuV9AoIZQVgIvvsxfBpaidzT/HUOnCXTPj7HptU+zjPXoysfRBeeg
gUEhsnR+kL/mufhWPqh/zQMTaJCUrGH3jAYHYTeT1HRyD6liWZbZ51jjDRNbB/pn
1AqXP9NKWf3iSwEItWq4/85l5PXPnnZnBByCYgKgPKzwmCXf2Q+2ZXYBRIoCSsLG
w+6pOKREVoQWkziGoVgEDxIicg9acmz/LNcFyXmP4bbNeG3txVS2GzBi6yXcUozJ
YdMEWNv+AEblgJEps7g92Gtd5lem/H4uGGyTJfZnSx0xgJenMvjQbmRdS+pLyY2b
7W2VqY4emr6Sitg3vUWuHmFsP0zhBjZT8DcI3z/83yTyYypv3Ozp0RjMY01UdxkP
17CQDsK/c52CYv3nzvDdFSXZMfEj3qJzz6KB2IBY21uxhQ+M77BzVv4KjzIjdN1B
JdeDxckbL4HfM3Jg9x30k8hcFCjNxrYOcgDPd4CxsilFoEqpRD9w0mqpJF7k4UyY
ItA9anFrKsQBhfFQUDufRjBqNvnPDNmWB369YXH3hsJcydi2dTM9OQonCUbUQCpb
cXrYDyc3bcOKMaK1p0jJ2k3KhgDVvcsUxt6GAERin0U5elIvkgBGnGnGWwcyETrn
hObrSlXdPw1VKF2Kfl4T3uxZYtMpGNqXKUxpwlvbDrYHQ0sRc3el7YCTU69JdMBe
ZbZ/CNugjVnPVWhM2Iit2veA+Tu6TsWiezJ8Ji3qCnVmJ6KT6w9g9r/byvZmhjmD
fxiIcqhv06bVKcRqwqPG0whiYts/VjN40OW38Pr0gk7q1eBAWDrxS0Y7uuuFIc0y
rDNmZB0qo4vrnaZYli2+QoN03+KJwUDcu75nhjyP6aafiM3dDJXu96dwzUW6zRZ4
i0MnbfatRIJ47GCZZkruL2Fc7FoQ49LmVi9wsdK/gbYKnF7Zcqk44wXSrqq/lf0q
ERCCNz4v8JiaWGlI8rW0hY5cRQeNK+0fa1lrOHY8rv3S+3+OV5ddbgkfS3EecJ+P
HnkMTcIvuuIvkKrrx6pJGlv+hebQS7yX7mHpLzdsJHHE0yVuVx4gp+M2Z+3SNuKm
y4nysLQ9Pzo3Rvb3JB61ieVBdzdVbXoDrs44U92cuT3+KVC1mO7QQz1ImJUnwR1P
EWO4J/zVLiVMCM8WWIFXKA8CwmAqf0dtEgY+uzKx2ci7XU3Bgf61XQuWB1oyrO6C
oWN1JVFukgEf+bV8h2WpLhvCSN+w4+I1UQiLi6GFCt4hL3jJDxLB4psCQrv+N2nP
jvlMr7ddSEglEiCPvfwI4CFHJzaoTbmWuYBQ0H/488dO27V9Zc8NSeYBVt4zYsmv
l7AiJG4u5oSnZkjXdPGsTdMIy8H+uyv35ZiBZY1dI5kTN+yfhi8NBW9F+4mIE55c
2AMUowOYOQArzbS1D57bvXmrupqwKZi1+QHZYGPdpxpYSG5b0TzHgtuswqlbkOg6
aVbVhidfG7mg78obgFTt7H7BJ81GjkHC3q/anUP1s/jlo5smjyuDLRex4FjK5EkH
sYS3aLSSH0ttzK263uYH3nJvHrjHv5lD4P2Xz70b4FOtjOuTCanKNX1MoOBpE/OE
/SBdDTGV3AXv5VqUDR7DclLzohdcP4jgDwS0dqiQLLxsl/FLrjBwd0h4jjsClWpn
Czs6/+kUe5EjvPlBQT1/E+c0Upw0XCkuGxqCIxoHuq0JW5s8W9ZsAqLANMtV77pA
LS1dUXnAJ5st61PliGsh1wOvFxs53dFI/lk6+j7NmVB76P5+s38eAfcNWK13J2+W
FqAa+IxtCem0aQp/OP6/4uBiGxs0E/tRJR+Iz73zjEBdBMlUEcroDBCUWFBI7dpI
wtC5wIjk5S7cSwDav3XSYh1GJFvWI4rYJZnrabmNOcPmiPXDdStVZhlxEBAvIB4A
2pi44ZHGOyiVU7m/ihCpMd8kClblwBQGFbA/b3a8xuFtzy0ArjHdxgeQCxn3z1Ty
Y8CiVZf4oORCIhFsasVIGEm17/RcNykv+bmpgXFqW2VS6CwA2E2tqqf7o5V18wZT
KElyT7srN41G0dVPZagcqIuhr1ymvVsEhBt7PGUL0llH+0ov0kYlw2TWvtoHK2D8
m26wVryjUfbxLvQxXOJwmRlq0J+j9ecATrrm2lWBbIIfdrb51huALlPbNN2BRm73
teHmi2KEii0WxNxwr32JSxe8J0G0EduWx7QsWhlIbfywcXhZeBpKttBrulyleNa8
Zuy0Woo56znLVX0K5vZc0kx0EkfSLhu2De0lrt6aowrdUa+/2glQRlwU2QsjOk8V
CoW3vqS6azXThFbHM+wYGx0YGS/uDEzgTEh17Km2bjcU+eaKNaAXrpawp0jCYWI1
XlsXJmWc+Zw6SgfWO3K2FJZZPGp/iVBrcsUJ7oWbWXU+i0P/iwlYy34wQHBzntfe
tP/jLe9OtN84btImT6co/ewN70gSVHfD2X5DzZ23s8x6TSoBZhCM3fklHVnNVSvv
saAje+YVyh8REUSDpvVH+2263pKrxUuBvCME68OvsL/h77gGcXDtbpYjD6TFqcFy
Ptl2cHnffd+mxRJT96QexnT3OiuqTEsQ/yqdVdkumAp/oOTg34rIWNk/Ze8lbFg/
BYVCZCUzamlhrbjHvuFZtsiTnm5Q/h7YFx2b6qSOI06808ZXqD+1UJ0X21gacXQS
wi7EUXo6qWp+jlN5b8K0bMBZMDYFox9hnKZIqNxM+5+S0la7vNYfpYFBIg/eBHo+
Ds5c0wLi4Ik7aLJl20wQUA7eBpuAJxzrhTCObdhh8m+azZ+J8USqI45TL8jf7DXm
ar+8YKzJGC4jdPdOOHkffOqtC+UJX/9fm9FRpwkozY3Aqo7E6tqu71gWcJxjnf1X
9DohTv3RIZQWTXpjxkgQ1VATKUyzsoWtGQRt9aJFn6qKUhjqsz9Oy+GXXTYyzYeN
iYIu5JAf/hJfGR1AM+SJjsefzaVDfPRLG3zYwwrQTS2bOZTMrgYG08G+Z9puMC+7
ozq4gA5BZ3SHUWM8Uev2c9Oc5UrhPoJXHtXQp1B7TVZxE54lRHeNHS1YWLL3+v+4
qn2f8IDPgy+ICcyb0Lls4JinKzZdmfrHrJx+8e+8j3QUC8Lka1StlTt7PX6az9sO
sN1MIUMbpKoa5MqB2OgTYclylh2pgFEEJMR99XxQG0jHXPCH1BAe5K5jgbd/y8TP
gURn3YGe4OKVS3CPdflL0BUg6IFu+UVQlBz6zJ96DJ7yyF9BBMTqxVvrd6W7hAN5
AVydF53/+mOHCnD/N+Yq/KzVVgLR8CFWNtTeYvNtm5XXyCbNajr6Oa53g7BdtjqY
hkhvOD1yu9ez5T3RwR+6Fdl/OL4zqBUxDfxVo2YdqUzZGWvWcPL+dXkUbeqMUdV+
bXl4XJTVrB7mqE62qyAOVZuZDqrZ+4qP9qRmQnRwpBZ0IvSYgk3DRSAQOeXp+GG0
hR1FOsm31Yh6q76/7lKiHmfRha/DommB3uvsKTJjTP8Z4nIJd/L0u4DfSOKVgDvR
tfBtY2jro2NFaMG33pUcZ5qgHTCix2+fuWvYFOcN5T+odsjvVMdTroz3d4slU15I
ilZ7kfbbedhb1x8WIw9tOz3YvEcb2/43rA2SYvr48QlPekb8/gnf5ndYWqHENj17
o8lnuruwNuPEDpvve7yiWH1IWxsKVPTYdYywJA619WdAJIWgofXCUNjKJyobw4I6
FmuXycpHGlpHHv101Bc+r+AttU43OOz0aXVXA1kvZdklz6RYBwS+C8ti5knuMWZH
aGfGshAFzV2+6EUy753R5vUduiZBAW+V1252QxshYDEhpOZkkig2qKvdScl8r4sW
rt+4CUJSP5hwVFuR5OMeIp1+YM4szU7BZPoD6IuKZ0ZzaYPtx3QnSSTLgYvFEEJb
4owD/fWJIF5xTZJID1+zJdDNv5XfCrdA6HhwRdPOLy/FVeNYXrgjfYLqQckHXjXr
2elj5enoW1DDu3gxzBQKa1MsU16MingrEKNhfzFJEoXJgT8K9DQtWI79RxahGbn2
ATDi1/RIxauLcc5i12gcTZtQ01oPuxM8RuAILXkym8z4gYSF75UfIAscCAfavxzq
Q/6U0BR07SqCw9DTT8BjNDrgcTo6f6VC5djckySPoJOMy4j6y4Bm4xYLOYHz3lq5
Xn0Tcgg0NBxosen0aR16kTvdC+U2OlKuBc3oL32/1IHZYq9Dco4ecwdpy2BdPWwk
G2HT8nkr+ZGpfEbiMiwtWKjRzwkMRkmjhd73E6bNFlY7+qSHwBnBZLrdT/alSvva
SlnWUAIU+ZFaQG36YKtrt2AjV8Lqu5kLU2e9a4LQdX5FViI0K6qHsiWXMgtk4sxA
UNGR7dbORktfMzgMIO7q2+qE6xzpzgp1AMDDPEdgWeIab/yZ3iBbPYvj+03yviEA
oHDwlyXApFrqeNn538Ght79RVDqsGQARhjzBSAHSK4onZjS1r6zc0A4nCaQ7SSEm
jduWXEG2KXfaeB3r08aVLiIiYEw109SmVJQ4C/cOJHG6yyEdyzcmikCDLUgrKjpA
TEFnxY/9AMZuKZZg1UQ5kONp3Dt7vnZwYoagGxcM5v7dCVvn+vNytNfa1R/iWqZM
eX/GbbPe35Ow+FEqOmm8KSDmqdbiOUDoGB6WMuqxuAIAkyQre/Wqzj4qzE3pwBP2
IUawQlEFDGgQcGlstOD1rrjTDrQMfOHgc0FgIIeEfxM+NneZwXDQ5zu8p7fxwL45
YvfH6r8uGkl6KK3xTz6hOoK2gFdh4U3AZYmGfCfxV+AwP8yQQtWQ9twlOg1yWClT
s9xBHIS28fnGxcdvHogJYOKv4am00b6/4ahCunMnxyS8Sr9PtLgK4fVtsru1dhFB
CaygFGjtyzo7NV+kcFN1HditFL+0khhE5Ps3pEnZI8DbFJmr09TqGPF3+7IPQz9B
xSWxDyTYYV9YE2jaqQbyM6UYtrKHh582svRsAtYH7GDhunGP/mYemtGce7R7Krt1
1ARulRiq4MAXA+svXIkB5P/QS/5mLS0RAC6AuXmNGsIUndI3sUh6+yuS5g4ZPkCs
dc5OKS6kH8OatpEpJ4piNRST4oiiKRP+YYx48NDDQCfS3WXD/9Iz7hG6JhP0kgOD
UXgDYSW1YIs5oaq1sjdfGUbcmisSGRX0UAHImF9ZGs5tbB4nyx+9SB9Zn05LrrB8
DNmtMDMC+8GGJnnO6jX5BUbWEwWheEZbZL1Fd76t6y36FdZUz8E7/l02RHv07Bx0
uaV8tK0GGmMsnonym2sIUKFr1GTyIK+hUsNk8GBDmVMMFKVBfsMrxzdMd4LGpw6A
pLeNHIdDBCiO7EPuYjoE3q6QlDOWDgsAkDkeYtEDBb+Mi8iESCgNovWE/tv1nmds
9SPQVKujZhb0Jyd00nwG54y0spnC4gtbM1P94Qgrh4GzOpx/hIllZSDeS2dZXUQn
5/Q/pZjckkYbRavNBpv//Gtl4zd5yaZVmnandX8d7HRlzM7R9r1GRcdKC8H/+n8h
tDgi1hLsz7YNMoqmHq71Mp0hvXexgZbXB/9RYI2FJiH3+L19igwyNh8280IqaNPh
TO/V/DPfnbrFFactHTVP+dl39v5rHQ/l1KpC2hRvOJumgKycoWhU/pKJCPQuOuG9
LS5W5vtwt31dx3D3pEQvc3meI2GKz065ERc9OB+Z7IGaXP5EjxaxCFpFxadC0fDn
trF77duVkyoqi4RQ1msUEdfSq3D2qTDINIerflRTsQlnbKTyPNn6UCCvVINb8zpo
sMq28qMaRxRwSZ5b+dv/fqmgfOg9d1oqUdMUUxRAYcy2rgPK/zYf5k/4GiSmD2RO
Vu8JjWs/HKokICJriKwLKc8BXHWdOj3CM0OEaoV3/wbzn8MMvx6gGFjK+DCzX3qW
kl0s6vGj8B1Jbmo1WLCcmBsRitVzb1ocninDNvQXeej3f3dwBd6x1KI4Gqr7ZHkT
oCOL+zjs6SPHZV+ddbXeiWpXYWrWIpmsSYksk70yCOPbGHFksZ2Lshtr1dA/DdAo
GDV3LtNEfwJH1wKMRrvU66zBQqfxRVY0jILhfsJAsKGsSL0ExQVvOkDAe7aQMj1m
S1LCRkaqOl/GbGSVqKKD/cGg0fFqRuM5UJwSuoACVj8TctJvhpU48gDNs81usEyx
gzetyOpFOupJ8FmWJXsSjOhXPb9dVO0A2NpigYAjeZ/hELD+UbnU7Sp7Eb9gOmtO
GJSH7hC+ASzInlp+vjqcC3XBcPAT22p84cuuKgQdWgslbdeRKtpPiWWwMHGhDifT
tko7Lwo3x0HQKmXEzShfHK/6D6Kvb/XxoARcfHgRV4G4xpGmVTT1FwFQNuAakbOF
N2wgfBVmpdQKuufqhLV+nPt+URkwNbHvz3utdHoQ4L+2xtdcTVne5/rPP/zCWZdi
xbCOAVwhVx7qCFCDqFjtoePI65PqRB/D12nBh0bda8wn1QiFDyUmbd+oDJmVhf7n
E58XO4l5sj90DAzJKVe+sNzPhJLSE1wcemwkECmO2tr62xgi741h1BpIwS7DC0tI
QhUH2LepTmF3Hc0QJSb8B9cGCc4YOGxXlpmy6LmX2imKDohnGJv7Mql3DnWfFZJR
Ds9CfrVsVfU29y9GQfOOSym+BbBUivd1C1lamV5+RYmGE5VEPEjdH6ZhkXXtQzpJ
dr8AhVPgPeokOq8mvlSqJ324VnF4k+d0q5IWuamY0mkoqDkezufTDYHXPp+DKoZr
cErDaxtiNYouzOoHBLDjupu6Ek7v38y1WkZjl3qTeMC/nlwRpAjQq+80E+DngGL8
yENURBHXkySXfNgxXO0oU0yNH2tp2Yv+vHMbS0Wwr46z1amWFlSkUkb0AC4D/VsX
zcTxM/X/XmF8x+5z8jJYNDFs2qryEpBhrXMhaqmEhscwuL2tnoqXUM36HQDouHqv
6AXtyBY2p4yhKUYSNFUX5vH25CN3fIHfIfUld0U+tLULgpy0vAI/WHsgmm5LuTdH
AbbqDeQ3m1wRdDsn8TG53+s1j2U3O6hgnrtQzTYicfwGp6UaGrvpguxoHDTtYu2S
7Acs3RXuFYd6qJSdYvuVKIhm9jIueRKSo6yhiu8PadLm/U4fYjV5zD1vOH6EgwLp
k4AvY5T/qYVOJvzvTpTgylQDYZxbg63tBh1yrzCLK1TjmaS2MxiT6Y1rjn4gK8VY
YUg3DOQ4Q+4Ri1mBJzv2tY3nLRaYEpv15HYF2bZk+FbCAVaFTTx4IkT7HG9sAn+M
2hskP1VcYqP65zSlKjDDboQoSL5Zk8+d490sY50XNm66MnIriaEfyodUydgtmy9x
RYtojVbAzBdI4c6Vhi+2qgWhS58DG7OpXS4DejH6J2T2b8CRht/jlNrrpBjaPTmh
+W6d4H6zTlJEMWsD0BB758nc3OEbjHlKc8CiPCXxAryEEbFqJZhWNbCrdxvADiJn
d8+G0KcvFRJ6TTErTrTk/Fe5ZbBUQoSZoKx3p+NW2zXSWUDVJfct6nXvkN6BW3qW
lJ3tfKHVTiEyU+ugtIg9R0xU/GF7KcT+1u0/Jtuw4V2crf2NyRoxTfMeWf7v2+uy
yeUNJkZ/N2w4taJtXd+B6cjIfm8kF2gmVvKC47QydRLd37XoVk7t03mrGWjrlOBw
9Zp3yZqpIdej8GmoKwLnifIvahHBMTy6tqNiZ7yHDz5TX/sqrePFE8pMaX3azMiC
nD4v9KVY2/IEK5nJky2Q0Z4Ue6bYJbbDsrANPCFI6PsV9LlSgsK1fekb5wTbbRaS
BdQjGycEXC4ImfTZDMuYq8BwrLQBwbw59PVIpk4TrCIT2ab/w23bh5sLLpo047Gu
WyjWq22ZUa3GBqyoYM00Kcqpqpivwwrg1Fqku1M8aDDxYFzBAAPmqdGkRVCyVzmG
0PHwnH8drkxB70yEUSod4agyMQ3nJ8PS1efp5rOE4Pv7raNuoKmLtwZo0WccKPmc
N6syYnP5e/l6G+AGqlDBCgVDKAP4irBm2TjwT3wb7n5Y/ykcRipC1YGptuT5TWYX
NWNbf3ybKTeXumNTpDnnL9ISeJkTsS10NbvOzqUC1quOMpuh4YCtp/tinVz50AOu
DEwUcEtctpg9tWjImFEhzxWa9zTOhWn9rT+vr0gfAVRYCQgawQYxgGSccNMvUItH
Sqt5Q2HqZNxQUrex1Oo5VacPwsHje76L2gkLWGzfrkEzqHucanXQPtiPUmrPnUTD
63JKyT+VjKHOW9WS7wMMh8pSuU7G3/bz0z3iCu29/5zzRce9i8krrbBqVyInq/6v
spM1fKP8gmUKHAhipJCLB3+V/iML9o/f3i9zNTdX/SiK3XJqrhXFOke3WBFt+o6x
QaEBgOwDtgvUsEY76Tvy+VPlsKqGfhAoZiL15W7yvIeZz0vYn0FXPvYLIi8fcRSn
EFeTBOdu3IcJjUDzsk19WQF7KBID1X0gkFWiNSMpXJPaKCFTd6N0ZiOK8f3YDTbB
oQzzKHk1n/3BSIcDC7OS8/m81DD5GEJOQzGmea1NSmiO1AO2hzVZGNu+QBEpla+U
sPZ+bxSHTYxBDNYJp2E+gcx/ShHVSqZWf5IZh93KJQYYM3cTEa0DMohbsKeOLlVx
9XB0cxO7IBTY7pOJk+quVcg0fL9Csi0QpIuztpq9UlPf2FB5mPjN6iUp1fJPu7ki
XfbBPL9oHY2X8PaEZeUk/TfF1yjudTCGqP9SEoolr4D8UBvJk3VZVM99CRWkLDCJ
ubDoPRbDxw2Ka1hPEf6VLAAfoIj8zxvhO7uLXJksuPiN+DFWvqsBv4c8mBftRWkg
J+cc4Os2O313rjSzWbUX/R7LjhGNFsnS5H49BTOcTWwvEQaCr0daTV8Cc9rp//lS
iwm2gKRVsSRQE5i+j8MKeWBm9VuVxf87ElxO+rc7RuL6D7lfJnKsQ5KRMCNMpE2B
VeuOX0ZaGjFBFpQ7CEpg6Xb4Htu0UkbhE0xrUio11wejO7pVDJVCemqD+4vcsiDB
d5ch2RXaWGIaosPsM2OsncWC+ZsggIbHe6II1C8H4dXgemcatIe3gxy4C8eemrPK
bhsnXLMbl3FUhMhT9T08Fo/7VmW7CV9UZ25bYlldXQAfZMRiHs04PhFaIIzcYdQ8
Ah4zZFxik69wceQqQl+4DNB2VCjBQ+HCAcNac+q+pfAUl1B5LvQB+oUw1ZNEY9TN
SKM7DCz68DNWNMGGo5dOdjoYPSWpEzR7tfvNz1OoR/yzzCOweFMwhYzmUfhCxiUJ
5CYEmLEG+VcPfmI5b890Eooz7GQ8lXpmdug1aMOXdh4h2F9z1H6vsVLcj91x4phQ
s5njxHKZdOZz3mLFMD6jsebSD5/yl67eupurIzSkWM+nQ52xo3sXU+98nGoS5Qpd
LnknaxfsQ7ZvhOWPmaPYogMgzdY4WPsygp5wr3BZ+6ODuXnAyxfrODy/++y44cdM
L+Ug0+BhqY/HVlSul8o/hYlA4w//w3Xrl6bDeL6y+FYPHiQsXhvVR1jie7mvtzaM
MGazwJyBRaQvx1lBZrhbdeTRSGdBUKOhoUpNannV4lD4mN6SCOdLBBZ1yJ4jxJV0
2dpMui13Bo4+Gv3jpE3Mzwos0w7d1dTcKRxF1UroALsuwAAqLxQMVImWfq9OlqkH
dHEW/XuFrY9mfcb50jQmFq1UbZDSt4ZLAXKqezUPdLeBLNtWTICYfsDhro8q/Pjk
xrBPz67Yz6HIjJplt1PteY6rXjrBjjyq3jP3oBSFwVVxGKMKgyAZCtf1LJLmmKM0
xfuDP/bpe92LtYJ28U9gkfbTPUwwea/aP7nBdMPrKkcZyI/cR6iERHfm5HKDONuX
T4WjThnAjhT7rvAjyawdABSddV489Kf9/p11tc015SR9lTnJYsLoifS4LGENXAmx
KXOGq7xOQhAj4mCFAYvc5Q7WBol2P0H2jVkL8FN8HX48R8be96O10zC48MkXB90s
xFbTh5v1gxTu5Y6awrJgQHIkto94sImWwixmqcmwxMwbT4npKeoEl+g8+h8f75cg
1/7jgTzkS7y7L39UHkrtfQfEnZO72a1j2O1QfMWfD0EnjeHREHB5/jcQGxBxsQJO
3Lc25l4C7QRMc7scWEL3mEdITtWk2w+lwOwgQsr9g2L3fv/MbOWmi1ZxAm14Tleo
owf19I0dc5U7sDDC07ZOYivx21n0ej6qqj6oc58uPbPNhks5c+ipvzGjAlDgYt8N
/jrVUXa7MvSRfrXLige9bNHX7KPELvXfqBt+KhEvPW6z8NYBbxHrL9ykhFE65DTi
4O1YxB7ftIalODYyvZyrwWP2uPXq+Y5JYoAbP3fM+8eD2h5iqDQdG3OIid5X0/lA
K0oZHrAo65TXHU5T7qAnXhqzxTQicALjOe2+BsUB9AIgR204TkWV/5PkYCL3CDxO
m6BrZmqVVmfU4pD/iwx9ASTKcIcuYRboGNc+LIkQ80fCz8zpyfsbc5fg8hWlSA6U
anDApc3LpdWW3WC1+hhQ1a6jiI+NlmR5vEqJuVn81FWYYTXOXk2DipZygkqag2JQ
JG9kuUBQbikSa9hPFIuUW4hPk4PLNjkxZS3Clll9MjuRuajcwxJXbIvu8C3Q4+zM
SwrM21B7S1K2UdtlaWAVz4EDVC3JmBjNnRYWGSN3v15iUUuV5k170X9vfMGBtQK9
4T3gt+YsFeMrTATq77bJ+DjBTEXK6PAUnXYTWeJw5bWYSqddShrWzuDpbTuNsvis
eL9YW+nniAl8sWzp82/DFQ7nKGiqtSH28OnEQ04JECiMDtZ90Co0iN61QnhlnhtR
MCjTmQY+O7CxcV9G4aMGoPFX7yHTThVVWStuQphGNKzH9WxyOItYue+YcDMb/elU
O4Yl0O+f6+8eAy4Xf7HuMBoX/ls3zRO0HogHDAxt/I6/m4ViQZjMSaVxmvtPPfxy
rv0ctADbuZgZ5B/fxcFZ1JUrda/TWZmbmefVJQ2rnGyD5sBmNI8pmW78QiUbt5jx
ctjQwb+mIYIIpgVh3XHkUq+elSBPsTm6XyMFy6nQSrMn5UgAZ5uTfTdUgi4LNE3H
3+pTpW8xFN5SaHMOPTPjpWr3jYIbVE9AOv6Jix+qE7YIu6iJnSFkFoiwtYwAEZZN
XfQN+RYXRd7CKuuS2B8EvvIRdq9URhWD9XDjE/gb7vZH6mYeSAHSi2enosOU7sOV
xOtyV4yXiaOCFL1oGycNkYWT4VKCV80tlOk0DJJDQi/2IIOJzJWa2t50iB2t58HL
OOpaA+tPuUuiEcVUOYjKUjyMF8jvTWtuJp8K6IFXVPM6oBTpUWZI0T9A/8DBNRAB
hdqcnGMBS9G7hyYQ8DPxTtexYZ75jXMvB5jNHTLyaQ3pc9++cLJVDFGFxvkbRa01
iO6nWU0Ky9S5ayQFOe4xitZCsadn1YAT7mDbGqon55BcaoiKoYphhE1vTdJt1MXK
fjQNc1sOAWOk+t2RoarELnIfspkE1CKUzGZ+4L9hhMncPfE3q56iiN2yJb8t3eeu
6kFOBJLzTVP0xFRMILOTZJ1EPHRp/CLILuFqbg/CUFqsDoR3SrG1OXCZ+/RU5Yjo
yvATAsxAcSUwEFwQdjeg8E9vumuoWYMn/RQao8ouW7RYGViuZoXyE9nG0Pb/DqxZ
S9N3SFtOtrAn6WYGJOphr3Dt1wsVX2lLooigxklFVAJQ0Njy9lBI38yanFxJudWt
1nWxb56et+PwPClVy7h/VhubncnBoMYD/BOg9p4AVIDU1RgoLUQN+37OA63pmn8L
IhyA8gYyc+OPANEMeSAlqkkpPALFjFgyjiTfiDx6KuPPo0wYXknV75F4wbC/LA5f
1A7+LNroRQ5SqANPcsHyAtlHoYiFcZledScdXXVTsiyy89yirwVjJQtQ10l+xfow
ufCROYlIckjr7lDfL8zbPHA89OGUtRvycuBTt4pyE78OKLmrf7kicAeNcpzyzpve
9UTKbuxEpX99RdpDamTBxu2xK+gt1ubltZM5hl4m1CS9Lkg8lPnCur3pBGIaUIRr
J5tsGF3PgEgshBzJYLUy+e3N+ZILHFaG/XhmEw9LbuF78RqVSlMP8IYu9fi2D74A
pQgCppERMIzks7xn7nLGkiAl7MOyV4WjtCoq/N19KFQrFgTCIKTRk2p+iAnWDAGb
s+PV7rvfa2vBLil0Cy38mR43ZyCCfAQO/bA9fs5rOTs3kfCpIvgx1RUoDhs/wp2w
xAUhlfNKQjcqRtpIsyX8F+KU/5z1XTuGg4+lQsZY+urfhxi8+27Y5iHyyCf7BuGw
DYUkw39Fw/QzMqSCeAIQuXeu3geKgnPxtdrtDtrSXHBPJ0TGxSxiXV36AhN4/muh
JiH16Cg3nJbsF517048hPm2xOUvY4MOeWqE9MQO0Xj7+MNM+Ij1ORWkmfFqSF4SF
qZoNuP6uWMKHFzQfTdOxCU2vFzLkXAZR755kgBdGz15p2wnZZ99k8vmqyKYDaOSD
VaVEO5UAJ8Oin7FZZKwbQ1rPZIIop1Ubyb+DMa5FaDwyTV2ETqOFqxx9pumoDot5
/23tjAZpWQfWyMsoI2XBycm/9QAk81TzMStDeW9wJ5AlsuL3Hrgv2NWUbExaVKgS
Jnna+Il8NCEyC5tJaJqUD59X1PikucUdB7sNnCqpcNE6vds4FnOwqvV9nF3EQtVh
cLYHZ2P32r6He+FBek6DydmMgOekoBkJbunRAPYBXfdvCZujz7Qty3g/nxswAEIF
hYBS3wfCp7q/jD7sVK6IufLL7mmnQgXlxdQ/eFRjgPqjZzJ/Pfq0qpWuiVe7L6vR
Al3H15qt5vYyxQWUEFc+SHD/edEnf+V9xZUkmPl00tB4S3F0NC6T+vE2M+4I3NNZ
fdavF4axtYOiUDxwblKGaCtopWzlnYvReSK8jI4vuO437ib6iLnjKNzrMBqvwz9m
H6sf/TfhwHl9j+5RwYIXBhMeDV1auVwS7vlMJ/XkcQDb4qqIdU5HPs9lLOTt9wb0
ij4/bo6I/qVgmiLqwJsQwP6UQdxD0GxFVaCK+yDxEG9WiTROWDVojgta9I52NoSk
Af21dJ4iboMARegSgS6dj7iVgZHyfwa5Mv/g65TRfBblETSlLi88xZDUd7LYxGDp
TfqWPOtPOe1+LsOyWPfSIDuy/Y2sIddCVCODz+HFL7LskWjp7iCMMSKCbNx+bUsf
oz/1eLChYnDMqmzDQjnS40Fp8/L58Ub+s4BCB7baE7jfp/lMYDuR+gh8ClefQMTB
OOhLoZEvlugHWBGDNfuhWFG/guh1MpdFfia+LTliLqgJDaHBcBRq7ZCVL+xw+U2Q
ELGAHnJNjA3Cx3KWAAUf3xJR8KQJSLJyHrIHHfsaIUfN0bfoUDIEzIEJNHUNp68G
b/F7Z9Sz83YngclOKcaPiCElvYjmKhVKYutIdCfJEOc/IONS87AFPa/23Ps+4So+
8m9O1RL80wU1aVv4tAfSJVJqZHuA/wnCNmd+/Wby6Kp5uRdBD3i0wCQe8mBwrPkA
lGzQ88WbsoeOAryWQOFu1ehVJM/rviHaDtUr03B/8OHS+1tdXHIcdvl7hAWwee97
De+kAB4Qm1FaG4rJdyyMXIPEubINwaWxPs2Oi9wGCcPyVJLPOUZw+JkFNKzx/fFR
HAvb92kPnycGZoIwZhIdzlQ+u4D7qISI0Ng+yO/+6WG1MZxQscWvuoRc9rgrCaui
IV+UQsfs6PCIvDU1MDrjO3eDJFxd0nDosClgJFkbdQs7s0UQnKQRkwNOqGCT1+Af
JsaStE6NYP8Ud7JYnpjufWYLBl2IYaVXgwRgehcFJiY6kzqve06cGn9SpLS5lOkR
iJBdQ4i+fpupANtYa/HsScYZo2DpGa/oolpPqLacgx/nLGv0yHLWdDDcOU0HL/Qw
QBL1IQ8geQVFucV1zQ/Ul4XIhrJCIOc8F/+mJFKZayIv3Nt0RZJW/a4H8Zez/fJh
0tzbxCUr7g7/zz/T4P5QPDLFw/OmQYrY8VvGlXj4/keyLeqSk3HYesGNLlgR2u9S
4heci9kcVrOhNJ/DMJuDmRs8Xx8KUAvhHJbDgwaD4Qwnct6FqEskJ97rjsCrIR03
yjCNqUdkcBsetSWDzZMSqEydcK2WV6dh6Mog7B6OUHfNZeNjHWckDFzRxkhRgHgq
65Yhc15sHgdQuM1Ez2bQI6SkHQWYC5OZV2MDoqxn9MhxC9DTLGG6LBu6NeP7MzJ4
ARjQ2m6n/i2J5QfysR3cODSN+W4HS1oDDPY8InNHvOOB0iLDA2sWHwXXiCCstPmE
i+i8pD1lK24IqhLk12icjg2GirJx/t/3hLtmIsfSzoSSaAQq2pqGtlL+sImjCYDK
Ox42jxmNUqT1kzckKioZCoUbHVsy/GhDv8bym7/KefMavdqKeqd5SLrUzR2JZ6cB
GaoBwzj8TYKAWz083Qt39TJ49Yoo+wsLGuAmkintJm+NfkZ8jZV77U+RoEO97MUX
O9EPrzRe//HlytBA5BinkAkSbSu6PJuVl16HO8TY/j4gdRsLt4NSNtT7ISwVKLIJ
zHlOEIpwEerzL6hcdbzAu6hC6Z9BjPHUBR58yWDT9mtNdUref5S81vzK/E6wfvxd
e6uSZmg+t2SuWPgXpkDXlOjfnXvwi9VxdijWmeoh+NAf8dMSw0LFq1zCmEVSJCn+
wy+OXu2hp5YGfMLHgEHlt0s/Tx+82bhASXdnx8Ns0Cn0CcZXpod9ZDxeaQzLXPe0
WC9OfAFayhYMn0VtyFjjUuJESBwJyhuLaVHe7USTu+htc7tbFbSSeS5bugErUfIY
AjIPhF4TtxhBbh7jYg9qzHyyCmk4s0vpMrBtu4IxIM5RkI1pTBlT0+XP+RVrDO+u
D78rkC8T41dlVFGWS4454bl7RmzP2PLzC3DvXCCBQhIhNYEVaxFSdz1akHIq603T
n8o0tDv2wezarVRHWtdGg+qIwZYPDFT9sX+RRAY2a1fRuLRWZ4Bgn0LltHrHFxt5
TNnC9AnTxRMIVQxQQUE76t5pRd0ZP+KyXu/QmiGd6yKQZIhp6IJ5TSuMGBqLk2q6
QPZNRk0UkDI7ttuBIpb2WSSOJIxVZDYBocnXtot9ZZ3SIoXg1wuRV2pEeuKxv2G6
ylOo0vnsENUEkAoxEq4AfHS6BVT1NwbemB56omppplDFcG1F2RNyTLQMnt+hBnBQ
WHlOWHnmV2SNnUD545vrsMvQD17uGukaNp7H3SAqdJdmUKd8iDXgHqzXMtg/Cyz0
K86TvWNJjDzaMAZwVJzPSAzTPvih6R6qSGWB3p4CjtqJ5cdxH7okRVrj6uq1qWDv
+KwGMBWOuGIVXJK1gRfy/3hETHaIHkkvghGhLcM6t1OTgFFK0vG8P6UCDpICcRN3
nzurkWECBJKVRVXU3lzL1DnIdiZcPagswoJF8Aq9r5WUsAgKarRoVE6XHzOChivB
tKnsLF63nUahxnom5JJFAnWralJxOyRuSWAHKyrSN6qc29ImECnsfIKZ43sEA+x7
x7YgL8SPeZMl2YLJ7Ik6eZBACud7gKx5R4oroWUtEAwfQOqBum53A/iUY+e4Ques
pFM5+L3Pe+0wkTl9dh/RcU2fs2u6IheCIm/zIEa8D5H1HH0Z23S3fpg6m1B3M7p1
IrbepbJJruJIrO60XOq9IAjFzITCDWTGSWKrC96Qi0LKlE8/bW1sppbWWX6kToS9
QpxQJiSrQPIqMnSUDOp8dprzj2JSOoItlMKPRTE++ERyAOtgoiYLz/2S8GAW7mKK
xQitnHATZEAs65So9l7dIUxp4LNvFd7O2LG0s7gjpNGSro0LZf8nnwjJWa89D7YE
Oh2GsRPGybiNtQpctpMd9GJMTJD8kuyPUsxAqdiP+iQ4/x/7nK+uuFBQgEKo433P
/kLhSeQi3wn/GptaZstGIR+JD2iihJzVn/KLg8UFuBqBEbDe0rWRpTIPRbfQFwnk
yLUfBBynSHVAeBtfJ4sDwvec5kFK/cYoSCnQON+ecL+PRqipg58HHrinSU7C2Kqp
3rpO2hlv2oetpaKoQdvl1CP1t8AdOdPshMiVViBMXF+QtE/uPry9qqPqntpLdDls
XWuAgMBeSGk9CNgiafBwZyhiBFObxMA5clLSxwBwFVCDgriD0s8uPj/Nn2mXX3FR
kokcirojKyKy5mraPBMJI53JVX3jkQLjhCvqRn80Di7dZFmnBwJIluSM2ujlGL8C
7UlNHNciL3aoASZ1DDAD6ch/UXu4mKrzzky4LMTWqN7GJuSDNUl8LXaCLmHO4NsG
JSWdw6l7ZLJs9V+MNz4sxxIYhARXFztvs52090jxwaSSxf5Mo56FJu3G/hTqjPyT
DKFpG2NSBlNJHofLj6xG6GCrSaNLzKkvBdeH/EDL2cL8HZ4HiChH5N9H/TLVaecF
+kZ+ST2AhhK2oVHEKmn93OeK9SK7XMpX03zCJfbGHjIKr6q/HjFPqIO77pyYWezY
Zfmx/43bROoaBlDTYt8+B/G7sPVv9BAFG4G4sM9Q2StfX7rz0yrQ6xX+UCCPov4W
8/j0C0AJyCJM/Ja+50Mt0NWlSlmklZWE774a2ONunX6s4DrNW+tZdlDrHtYA+pYN
wMwg+BWNcOpJaiPXfqDW2bEOyEGLgREUjv5sm+DudbfCVel9U7ULyngDXCci/Cph
JF5+la2yN2pyNJMlIftPMCDdarkdzQWnv+aBLBfV71Kr7olSUC/DU3i5Zsb4yA1L
AFbKKg3ww1K6nu7m4OKLWV3qib1t+W3/0LH6PtVUNmKHPesafumRL67N/fHV+4NR
oP3hScwHfMeJQFX+WvHapcQrk9mcnQQ7AR2m4Rm+fEH6MLcgSmjW6Z5NSa+K8Rx+
mXImrDoPJFWEDPv3rY/GfdugOsZEEP9tTzh760sZFu3bSFNXfI/A1vCDYifQwDOk
B4vtT9l3nky5R9srVfRoeZ/hESGHOMINDp+7IunmqRrZKiEPQmcXn0/9p82ihYDT
3rI1zNsXT60wrFTcP+Ikhf1ZIMiBYjR5san+uGMdSSV/8NAkJB1RUr57+7bR/qN2
pu/IG87P75V2SI9ox4t4UgeSDhU6YBm/PMYcuuQmbcqadeQmT9MoZNkHVerms7p0
lmCq1FfQQuPVNW1bhMP42J0N5ZXP7xcS+PUBylYMyt5jcLd/Hucb/sOMv9Ei1oJD
OAhQjzLsyPzoAaYP9+nGkTigoNy5B2/mh9o1OJSnagSeLW87eEe44opw3n9op+bw
uUls6mNP1mgDRRVj1FHw0/FXeXgG5m/rW/eUP8StHYixPGXpD8mM3Pk0mR00YEjA
7ZTh6UkFXPx3gINwz3u5R0cAlKT6YxoQK6x60Q3e/fNGjlWlNBzkw3oCzyc2F8b/
69nnGAbDVeBtvf58n8p3QeV++JABOy5toOzNdPhxRXJoU3ayQPues5AdtZKTmsIj
6b/Bpr/pMOR7zAH867Ns/WDwszJxmtFN9ghfWCsve3Hw8Uj6iXe1yGtNpFNNYtku
vbXvvALQdNSCMM3nFD+i2szEULcQ2a+XhI5jwqvAOIrWmsOIqs5l2ym6hjRlIc6G
TLk4dAvrm+z2AO/ksyPKYIoRqoV2BP7rfU937cSYhsjfnNDEgsa/CeFJ+khNhTCb
pzlSaedNAT1PKq9wRm39QiBOpY+IcLXmZTLxO0z1LG2BekEL79qoVf7iISMdYlXV
FlwnU7m5L3G5n6TbO40yMVvEATEbZlPVeHrTDxyNYtrjq5HNm8B3GWKIxzGMPXG0
GRRO4T6e83F/H9LHpgaIcsbR+byOk+yoWJ+ltbkarCrgV1Ti6CnICTlgN9Lbp1V4
Os1wgoXj6JPMnhUAi7wabB6LPW0v2UGp1gCJXoPVwEwaAlczR0kOxbf1zDueGCj+
k9ysuSyrGoQQsy7jLaf54rTFJsjeaajanwViNrF4fWaUD9xPi+KUGYJ23WuZUsnD
OIhUDtDTuns33BxwSKnEf4J3WoVgie11cE6L8O0az+tgBO6QnEz5g+s2cUiRNouN
Mb4YnM3bWIYtIvfPf7NJWYudfDOz+v6j23MkNZ6GeqC1btdQvm5KI5o+Kwy7GAKP
t1he8KVVe4VD+IgyZsmQhD3BwNw7KnKoZSKFngEWtvDmyzhZDef3BVOfZn9V7wYt
1DsdUJruFS4fwqRaWsNznHV+Q4pthB2GNvnYPkqGZd1bfcADLZE5XkHJXRr44eax
D8Oxts2sV51K9L6lV06VebuxU7S8cKmeTcrs/m0j7a8akNdzo6R9+sRDPEsAtCWc
mmOEnwjyQVVbk6W6MOvL9pIjZYIIONly0sNIhZk1QCmKYYbRYtf71nAL9kMn/jU9
21JcIWQZad2hpEv/OkhJwQyAUj4ggkgI12irpgCezprIAwuzMl2JXbo89xVH8h22
mvkAf82mTDAczhOog1RLlsDEpY3TQTzkKO1/alPQhPpQKsR+u0O04IuIAO7Kr/pc
0gjzvv+hd6zRuI0FrJqyhukuiwiYrG0iJZTtk8sRBa8tIVz2DecJU+GyzFurPyMI
an6EpuqEGwhlF260gTFnLLZO8TK+uHfINTo/lbqcblthU2K/PIYYJ8IHYBb7Il0P
jDbpiNgsJRoO1/LLVRl+GSSlFE9NNWzyx225+v+3i5F3g72B41kd+zbxS+1JQ1nu
Sx4NZeIpBXezUB6nW0fInpnhwOA0SRzACnBKz4ky0LoJBMtaFTQFNAg4mBlEonDg
o9XxjOyHEsspiAUVfoMjuhzK0nRSrEZ3KXJpdXZbdCAKeCiMpTQ6vUOIy9ElLRtk
xNwifDowEkyzWqHRoElmwlvv2OQmAHFuNvgEuI7L7q0cLlYrUDuCcRyEJverD9S1
sQ5mjT/Utz5BDkFyl2fyO1Y9C5b8mqi26RSRcUnGexr6Gh627uygbmyo4wk/XDly
GS6WLmaFIz5t83fY9R5jSVEDRHyN6SNIO/E05q69G96ZPrHFqpQyBsMqf7dwz/cd
g3gkesuOoNLdlzDjw0XAlzgVQCegV9DF1H/Qgmniyv+cNbYqrQ0CP66J6WjaHquO
BKKAyP0KriZsHXusGS02oLKTrKj7FkLedIGVHyzgHGa3uPGf6WlXjukW955PizME
WaANCCgsudWAZ1x7heGrLQ1T1BMGhT2bMSslpd8yZ2TTJZqFOwWftT1Vb1hMvQA7
tDSBXME7rfSQBuJjajeAhdiPFM2JOqd92lzuAYEInpu1lAqGaOkRErTFeI3cJjn9
IkekYUuFSJuHGJSn4WkSMkv3Ymw1VA+qifYqB9FuX5OWUpWciXdhxoz8EN+XBXI8
I1jJnL9RczXqKMa+SmVHA/Si4dAw//1gfmmLskA/LMbSfVjujpFqcDI/0gpoVSmL
hZKebUMide2MULXbq55shQJByCtSMHiRe3RKNiBkMsWSYPegB68BZe+2KwKQRGIL
cDAm3ECcGnESpzrCI5DkX93rBahX/82HS3GTwa1Tk9d0ZFj7TNkNcxvxr1zomIWN
fVM2nR2HDMbhMsvJdYWx/aqSZmHmdv30HKHLeVsErlglR12a2ag1DKoVfrymwhAA
hf/oL7H7zsa9MksDY+tzh84rTFqeef4jRwmdcdXnOcaxbyCxDaASw9whIDo9349M
cfAslu95/5y9uHiMSGr8Xuamodm8MgtPM2lzs6u4O411HwbWiyt2G8WMRwdQ+9Uh
vIkWtkKAHnc3bWe8Y6CuGcjrF41FYPR+Ol2LKFyFYxzrHPYaMjicVjRkcpYrl9ZA
nZ+Qn6wGVkJcQJ989dkI5W48WF7GJW7J6HBrgcYTCoog/lvaKBiA4MIUH8XIgXh5
CrVQLpUH66+cWwdTCORqNiNyF72j9OaOTV5YiK3h2UnGO++rR7vSlpXC5HCF+2tP
NiNXDeDHsSRB1J3xanjU9vKwkakPip8FquEcWScodh7foysXgXZaMK8AWIB63xpA
KD0m1tcIkQpvGXi8aibDa6T4GgbQ4qHswQFa366TJVCrcXQYh6AP4lcsj41Eb22b
n1kX7NeJIoqTAoOnZ+WpftzwhVJNsRvecBqu2AE+edCHSwDUCZocLlZs16nZN5jz
qb0l+K3LMW4QMsXqYgMYidDCMuuJO8x3vVgBdlR4OCqSEDn4w5k4DLuO4FgR6WSo
w7+rQ7kNrpZV/haM1ueT+JLgVhW82CV4ZyaPhRpy4oN2NrBEvemosXTERJ/9hu8e
DxtWXWcI+ZMScU77J5IhI4F32vFT9z/9bkhupmNNzH2rTcAsfVOhRLG4h2NtF6pU
rWKXiSbYWypVInkpcH3g1LAD/FsEjVkGAeDO3zwf/tpjpLMG2UrWjn60yJpHl6Cw
9uS627yx7Wj3/dEddPEk+ZJ6+EgxPlQ1NY247H9SpQexfxCIbJNbtRqlxmUXBvdh
TmgBVMxGtIZEbMR+7xHDFrQpbcic5mudkDoo+W2yYXEy70vK9FbCuNbf+7o/x2BB
BpC+LJ+F2lAQT3WZNUgMcKwe/CoBzzigt50ArIUIm43qxk9BD9lf69r5MHldhrhv
BLqaSZ3aLgM4VyA0Vv6QFZk96uLIT8Bh46sNZnGGOitvhiyXV6IPwDcKWZyCXX9x
M51krjF3fzgLWzpqcuL6I1foVQLH2d1h8OviBSCUvXIUWmHoUEQyv8WebgB+97ML
q8VW66zIhwptGPkPJToH8FcoLjw2e6UKDeyiwO0QYJjINFNvelTefnsoH2W8TF7X
looYqAz6aCB+rl3jsNG4O6XqVT04GndmCdbZEMtug6hTw/dIGG6qEszS70aCeqMa
fs6TYNZBZyVshj3WsQxb5MJtMMoSmeXnojGMJW9twKXeBayrsMO8rF/AEjLD0iIn
b3oTHCPOAyv/d9dKoelb2fQJNzhhPfjjONwUtH44quEONn7L4o1NScJ5maGTNI0I
FPgZQ/FWhHEIr6oXRxNXUIJwKwfLWx7O73nYzF2W1FJZWfQ2g4rzPoNw9+Sv0AqY
uJZ8z4cTQ4Jrx6NrDrOG1/j9bjosf0IzQ4HV3zyO7TkK86avbIDnxclhN0gct+2S
YPrjqBaayNm+XBbypzIgmYJtZxyAJYNC6F5p2ySBDrB7JoLLy8HV72AtpVfSLiQc
N8NcVah8RdVcvapqkPDVpSSekeh2AFSE/JjA3Hk5mFpD3kGdcUlWVVAwpegcIbdh
yin1bkxcZsiW5Pu9qkymHkeibSrsvGWhLTIqnOXkmMF4euA54BTPPt1WtujZeoS0
BeW+VGjy3fRNsk7sWiOCsDsAkzCe17lu+n//jfP3z64APdaehRXAlIJKJ4kSlCRI
bTFQwkygeYyw7Iqq+i+A25+pIoBgXKg2bQpGkfwBRY5UnEDnL/vYbI+pYU7P6Ju4
f4YUolgax/R3zRkdIjnC75xXgdllgYNstS+etT8AcdLUIdEKNwxn8Mpfmh+rUkMt
+gLmxLtyesBhaXNYmNQL63IOCCV5baRny/ZMcZhjNDkbRedt8sCS3RuCZkji3UnE
oCOWMrdK9t+jEEhYx9szo30cMlGdxiw0215NX0xT0E9YSgXaYyBCewmhqJ6mQnGs
dqi3aUQYm9I2RQ2gErDeFg9KDjbrf7d1O7Ullyh0G8N/SaIBipKpH+KG3PEGqPJg
Wv9KyIk9UCF62BMoy0LMKIRaZQoZE7m5aIAQXcBkdAgay17vKDsbxHJwyQDrKc9b
i1vOdHtN1O1Zc5hyKfNlH/cAwlBLNknFnt5vxVrlyqWDHyVrKbaOd6V6P58yV4xz
J/9SKh60nigJkyRxz/aHQIiTmI2bI2oEJItXl93a2RE8RskB67IiaGZBycKmRR3e
Ck2vPr0aw91Jvh7q1/H+CpixphX678olIcPb/xTjtTWKXMpAzMAz18L1Y+NpH31c
p+GV51P3Yrya7+w6uoGJshL7OIlInpqgRHGfcxP/XevS5uLgHSfbkD6X7PuVeEg1
8HPo6qN3nVD1AOK8BKbEA8OQkVDBgumap+iOZHBQt78to7oBQmkdaFjfNrXupc9k
CmAOzH+hvVS5AJFDhRYQggP5GUTkUYK81KPNBJ2CSezDMyCGHEhzmEJ0NRNSVaaU
YQ1M8yqldsPyGkPxmBafoEizXaDuH+8JytWV4SLL0kKTa8tueqVw1604kt43UXM6
P/TPsGviU5gpUbqi9pp/oF+D5R1fLxPGqSKnh6DoyEetS4ATVyd8f/U4+xq4TgLU
O+bOZ+TrrFnsPoE7fFsOXQSIUsfJB4yfIKkE7XlnlfYdgErolnC6b3kBnqMeh3KP
OKTfW6UGzElhXRva2INKU/DN8RT+WtAn/cFLojBaAB5s/qUjra/J/+DVextZG1Co
/Ik3M3tEoCeAq7uLrem9pQ/3pr775nMteG1I95/cHOuwRffy/lJebGuhcl1VnP9R
Swa0UOdjYsmS37OlP6qcgVN8A7GI8cqcMitxLeAu+nkG/DKAKCGaKf3M1efw4HHU
i6JmgZu1ME0MDn9c0TmdkcWy0A0wa7qYNg2Icl/gVBkqxgvOi0lJqLXugJTXyGB7
aSTH+jDCoAi2rj5+phy/V09Q9JnEE5sph2NdmEtigcvIwz1mjVijZ1/kq6mGOa5T
giDgbXdvcvJE+lOnUOZk4DuCELq3serGodmBWWwuYPUsUFHAIoR5sR1d7R9h0rg4
WlbFHT49epIOvTXyzfMeYHndjhGcrJy5+AJsii4EnA5Lzql1Uvm7Hb6b8zw6lkeK
AVk9uw6zM3qX+9+VUdo3W+9v65iGpOGc3m6mimxMx9siDeIdGljvNWI6eZ06rrav
aWORDLZsxY7WhOw3TxEnDwkCRhg6ACqRJv8yhNe/d1QexM1cLbE5oTf5mAkz5z13
U83m8Tq7fKyo/GsqtU4iieAM8ebKehNh3VHCjnFJR2cZi1GBprPay1gwZ/0rF10X
XYSI+eN2dD7Hi2nLkkUwy6Zo+1+f7wTymDfy8V3Jyi+ELPG+2fhftoYUkxr0lU23
lJJvaimzL3al2DkL34cykMKopkU5BvQV+kMeuml3UE3vbCzCkKnre3lQvIRjL32D
v1Bn20XOfzfwlb0ZGvTdMCadTRANivDJ3AeTiC0poVmcXFLG7ac2NRPsCWaFZJTe
jIw5IdtGAjxi8sOzPGics/iBn0FfCREEPEKVkF8G0QYebCMQdzkWCdpk3gm8URrx
5jHXR2p85rZjLlb/3EhdDb5yXbcpvMhf4TAp1tV8skig8j9Fpv+g1bHUPWk/3DRt
SDswsgQaWnAgs9OlJpbd2LmS+WkpSGY8HLnYPuTJjaOOxVPbkEE+BOJxchkRHhH4
2J3I240Gx5DSke9PH5k0oKCZ4XCWglGiQRt6Mdu/iZ+PQkOcVI8fwwj4U+8PisqS
iograxf2+rsTAK9vY8rNBoPyvxNH3kmf3/VgeywHabtpd+euae8bTU3S/CReIlTz
8l4ml/pHaROH3VPCoAi3M2GCNAuAbcZycNAOKDkvBajwwfkqqAb2qfGMUXrCsA+G
iIZ58wsKOwo/YVZpKhRDXffvXOf6tiC4EPn41zmYbj5EkHRJvxto+k+aW9WXpCdN
KgSNOqIXGhFUs+3SRJNFXqFDFx63j0Upg1A5zBxvSJWH3RfJT5CbcVdADu7he3WA
yV+TvnFoH4KVXoXqIc95++5mHjEB2FeIjPnfwvTc7FP3HwBRraOCorcat/Ae0C9p
9NHVizAnB6jwJpLoSf1ghekQhIGNoYtidhDnUd9ChJPk0pCUosqB99Lg0iAfrUb8
+ip6jr9PwuYaLgYk66zpuAUlxPw3ZliUo71qu8M8xhCDo2uze1mn9H/WgB/GC1R5
i0zMuPACLhs9DM5mseipj5pqQ61gSFPmiJfAyGPxOot/bjIitWwuS0+AFneNloSz
+7g9KGLn3EQB7TZCbxrjlgZR+aYkEjc42nMcVt1DAi/8JpFprVMlIezZ1qHWhxQM
H/8Z4SpXkl1V8K2h0sR7DYXpzUpK+FVmHgaTWw0UPhIDKZm9+M+zpjEtEXUtoTJV
wBkcpNICUWaDy9E5t+T3uVaJpySSA+I6lafXVz/r957mYRpRcPF20Czyl9EEi4CE
Tl4Ax3IjIZTlBsCyXS/aWxmEDZUKgNi2ZezCwN1fomqMTfrMIA0qXIC0MD/hj07G
m19OU7OTszwgm6R2vRuQKvqLTf1OLUgf4JRIPKT9blt8jnopF0VZAiRJMIxuKD2F
8+rdDUELRklHMAqJYpdDgRdUUAygHc0aOsD0EWQZuhgiV+v4Ix4jfufsA65MmB7Q
/XXLZ5lc5RPl30sOqrqLFrheGTwfNACJkeyGVUL1powrxMMIUl7xpgOZym/C9qKw
3n9ku7uJtKX/G1I60Mjk5oAGXEHhA56IEK/0aLiAkvl23j8cCf/B6/s3wL/Y6rbW
Mo8Rs/9iIK5khrlHcC8ksbjyyfTiYXWnS/Bswyiy4LdAcfnMrDKRCS0bHwFC4Wpq
y8ggjxtDnj7hiSlL22gvpb2W1kxdDim77I2Y+m4g3Qj4VQZGbSPxTGXWsc885pXq
Aq1vF8FDbTea8ltqhzc7000IPLaAg7ZsSHYFrKswM6aMFYdeQ8bK0vesHgeTPZeL
LJJFRn7Qo8BW4VzYfacMetXyBrmTtwTKZ0ItUi2iTDh1g4GSClrbO5Rlqlr2h5AE
MPv/w2PJ1rx8NIcVh99yXVC+Z1G9zPSnZPEozM0ASIQi3899qTaczkai1I0ybfyO
nChNezSywHad+I539es85P/NxiliEitSfmkIgBY10Nv/XcilluzffT3ONnq8v0bn
fmeTh7rGGcH8Xj04yenycvCyczq16EXoOfVT1QnkNps03JUBMqug4g07e260wpoA
HxS3lYGFR3Pmf30Q2l/jNQdnsucVSYKpNHtMB8SNDOpel7LtOSP5gHY7BlpdKCPS
WrdO5If1hOQ11lGdP1dEtrENoZ8NJnhjKb6Nead7cCeHhyd8MCf6ySK1hQ2vMKBa
LBjbCLZAGJPTpNxPbWhIJOvhcOfiWJ02ToztoTxMewSimlqTbCmEJoDvNUAuCDVR
1EBjp6u5/KtxLm2ubwt1bm9M7ZV9lomx3gOFYvbe36su6NEXsS416+8DjItU+JNR
uKhAn5C1ZBqnrfa75LHvGvWKLkrlx1MPRJ1+iYMTb/gXGDWGcoBvvM7OghDnS2f6
Q8nAZ7B4z3CLdLtsvbuO74uQAJ/J0E263jpa/V7ywYFlsu0yZ3qcHNW/Esy0Wuop
zlBmMbyddEacZA3nnr4jnYGvwoKneMVqEkb7PrFl5d5f1XybZy/K8ontjsNFoJpc
J650f275NNneIxP/U1Y6kr18qizoHoek3owEs2COEAMPjwQE6jjptiYICMyBSqiS
sL6x+M1ZZdirCL5/oXGAvb1NUXyH5yE1isHDsCy5H40GdRv1qJJeLRyHhF/Kx51s
U4NiPqeoSaHKfwljaDtuRAKwKCyV+hCX3UBmripK9ErJqeyzqY0ERzKhH3gqKfse
2ksJSjg5Qu2tUvZtgwwS+4uSqCLxA/N2edKsgf0L+G5pqjjUebEVATdC7KGgXmYb
d3e76+ikWXBW4V/9z/nP1oVadBKJibCwO65XCsISo3fuztLuS+YZ37iyTB9mfUQW
C17gXKAYPYwX3eCv1Qtgl1xzXYlhcLbCHMyHexmriNR2wDt2e3BZ63LNZ8gG3c35
jijI90pg8m0CeGkuUrvhTCs3ZE108R2lul5aiKsovPwemFVSV1Jq8Y2ZurzZDypC
dcLt4Wu/oVCOnjeZ60jzikfLpnsKr6ojmiBRFTZ7XHJzVyWoURI822NtBna4B6bb
BIlqILBIeRCccjcSr38EGr5Mg36gVAhsX3BMy5n/VisLFBqtthNVXAfDsBx+tkXe
nGDeD12keyBtSXszHAYk+IYLMGDwLk6VGhHqVghNj/AriJ0VdJOfTCOnev7+8Vfi
9HrJ5hLLzaLixu4ww6pmpIUsB6phSbba4KHF/gDq9yI09pAwxhoAaZN8FOePdVXz
Bv/ePRzWHey+FN8ILMMeGzBXICebZu4E9LHsw5PEL2HbvStFytbvHRqztx3N2KCm
r/TuuI3cgePhcNl0nMoPq8kRdUZxR75KK+eH0/Ba01w2Q0pMYIKclDXmkKYR6jem
VO1Vh+l7mdP+H1SQ5ws4SOjsUBMZOv4fMfiwGLl4AmlKlirui42/XPmfYidIbG2j
j5mBGmkoO04FzO6a7gtGzSc2JeiIfBK0avsdWij/5u/FUuxfu9XBciiJAmB/0UG0
M5G2J2vYIi1m9c6fOFscaoeqaCTtKHrG7S/ZfPqibDHtbZeBhiyVM3DArw26Y0V3
94llYdL5C5VsLMdIKAguMg38p7r1LRS/0J7Zca1BYENiD5ibFSZ1Bhv0jyWc9Rtb
FYGX/LeC6pvcmsQrfwYStTdRrknLlXy+nLP+yQJmOGwZq0ESnhBTI3mWG3LWbYnZ
Cep+kXAc0RdROK3D8XEP4Ip8X+v4QVPBceY1wzZUJFW71EjXtlvK5GXcmUkbZ4tG
V+wLphf11if2nMvw8gMum6+0cRDb03MTHPISs3dxpxkcyVgC80t+0u5OOx87R993
hCteNyibCC686n3LWuYDwdSuTDr/fkaxxGenFKd9RNTynoroyTXNLnFX/ZcMDsQ1
psaxyl3OyX7E5NhkeYuH62WPvsam+3bJ7Ian39Uc3BckOItSsrMhb0RTxOiOZwkF
Oevkj6lQs+C1OQbA7TqxNW9mh85TwkBHjsdAOCX+XZjRHtpMkXspqzcTQZhKvyOr
ObSdAHYtzNI6PYggXZbN1zrT4oSP9bC5Dm6ycj0+0gD1lsZHFjKfq7Nlh5AFQuxT
9xWuvQ8NeXad9vSBHNHjrpwyOAVk5hRzCYZ7EvoHUhEazFgUZQKQ//RVA5QjEOWj
8HghH/rIu6zZ9OnUXnhvjwskJu5tEvSPLnwbsvxOmTAipitcegGerDBB6Kz2TkOC
44kw0owqIdzJaTCuYuQLlPeAV13WtDBgDYJzduHHLoiV40G1+g1Oc5TweK7gaMTR
ou91wLzLgaHZZoKrYNrmWKXZtrSEg9ZpgQ3kdJpCQBD7sg69ncT0XqXYxAeU5btN
8B8gqGtNcqzNPDF3ag9R7LiemMZ73fqm0MDmHi6UhuG0hcS269REnxB2uFI/Do2j
kAwyKp4B9zw1drYPAvWw5cmLK38qXMMA33JjsxPdG8S2IRBbwYaU+rdhJNWy6r/y
ysuSnvZTG1Z3TvUcsvybKOjR36x1wdWQXD0BtAokSLMhjjs8HzjUnAAPmpLUMXhi
2Kcr+J5RtmmujWhJcVDg4n7Hn0GtoeVSAjJQnG63Skjd1gAbcODyPyctXv3HAJiY
pJZQmRWddP31L1eHNaxR4U4iBcbPI0OMG8Tf+HRIN+XLL1nZmD5i39MbOogC8WUv
ZIht/Ks2cwhLXINRlQ8yxdMtr0Ktn6b9a1H14ofhFNzta6ZE3y40B359emrqQizh
lCCOM1j9llhg9xKB4GDNduGhxWjC4Gw51T8rApQ+fQMj6E0sOj+KAOOkPLoMHX+O
XGHeDCBdoGROR7A9qJwsCJLZkel1QrjfISk7DDXhXLJsigeV6ZC8Eai0u+xQYybe
38rdezU/38WDJ6lHRvlvqZQDQVHjWVE9XcMPH12jGqSVzzDxAw4ERCW+vT4zTRBy
RsGQFUFN6E7WDljc7r3x+b0Nx7CM4bqSavfqzKDk3H0ICbYfzQu4D3x6rfUuvvcp
1Kkbb9Jc4x8i6UtvJD2a4PBBBBGQHnmeWOwnQd6zUvAp6EZAu8+d+UZCWZ9yDs/R
XeqwQr1CuADddffUqCQUkMYIwRk61sD82tTyLNwUXdM=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EX/eEUmGWkNmw+NhUIqil0XBkYCV5EXAbhZFEzxxdNrjPkBd0huLeb7k0qaLdyUr
Ex7lzPKRW1+E0DISFihyndo4m//AHOPQ8GdAD9QaIBOEfLOu3uXCFl2obU+aI1r5
Hl4i0L3jwfVKrmsWffIMtKC9RWJtrInYromMCZyr/Rpou2SSbLq0Wwm1tWe0pav/
esX8eS0CAfxgxNLhiPlSCJ/N9oFCx6f7u/4y9s+ckHyZxXgfLJxrfgjzab2rwqdj
PG/gES+I+RAGDN4GNx1UMjaGoInWS1tm8z+r0JMErv0F6ZxgxbuTSClbE7rH0YJL
Q1jyIHjCaaAzZxZAIzpBTA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9232 )
`pragma protect data_block
m2+y6+GQG0HVhsBpdXsvu63gVBtdbNysjva2syIbNkFhRkz1Iwn9Tu5xUjMTXneA
M5J3wPKYtDK1ri0WbBEh+PXinR8YSKrJqDINlFu1XC5uBwSUl4sJNmyI9W/NTkr3
cygW7vUBvgaW8IxmO7cSEywudPohsokp/kXVmbZR8+hZDXV04YtyKIZ3ERdn4PKW
MPvkvw2JQQMmBJzZmEKHbXVNoX25Kf5KnOdm0/TYgGb7fBTVqIvIVDrbZz6iBASR
FtYdYY+4UcRBq5RUrAXOAwT8kkoJxSHVs1/wPiBdA0tFOCHGm+6oqTtahaaJXzM3
ZdelJ/0apqjCtjQxPPQKavz19wkmnvdA3kmqoEz0tIXxdRBCA6SjnA3LB2qVvEL7
bacXEsbpCEcJuvCXJEtltCIyUx8Zr2LpToOj1MuVqXcYVvp4h6MYyqqojuCnRWKD
QN+PkOG8RdZY7+k1h4BaGofBxDDEQ2SD082bHxLE4uMsGjc4owufcj++DRDyWNz8
fDR7OkDJtF9fsZnVCTUmxa18l/R6Ct4m5MgTGhjk1QPf+eZ3xG77hstYd6pKneJA
MI5PaIggUMCTarHBnv0QTjgBfymPE5SFm6MPxQ6alhvJgWzfNrYUKcreMrNJyKIq
dwqpMvjUozXXocMcXv4sQOOagEJE5csgziFN+CVqlBDg4eFAMwdMjjBvi73uzwz3
hO0LMLo42SW+bDmBBwyh7KZUUPz/v9qd3eE6cifGhYen5pF7s3Gs+plu/SumaHNL
VXgcphSOB8oRsIgP9MuDXNRoo3NvuE3BwsxImVXZc1KxBX1eXNkXVrUr4+eI1k4E
CWf1XFlfULyrCra9xVfulSFQ6PGHhVmT7X54dkD62fp3fvdq78o/yD7T3Pv4j7nE
s28LVCB4Eh1pAxbt7MD9UIo2BIyGeJeDK/VbAm1AbRRzgqTSEdmOGsxZxh+5YXbz
jZQOHL/xQQKAkTnT1t/UEI78FWa8vJdYanJEtx+cGJ4VsZ4dcCy16z5XZw5o8VQU
V/dfUaCbGxKfIOlJagqhofZ2W+VrW0tcgMoEXha1bECef5qYGbmskxzoQREQ11Xr
9HfDOJJJxLiQ8+Kr1YsHj/UOkjJqaejii09J/+EOAsjVtY9zpJOt6rziUF2N/cws
baRywpnWiiR1WtIVnASpWfCd7oLOMafFVZU+YXVCTk9U/60Z38Q14ujH36tzyGwr
SoYojY8GkjdHi8F59p1cH7WEwwLBh0mF4vRdyiVF0KxpTZI3aJKwXzVGceXnmoEf
3UVPaIcifcnX/4s7nMbWYNBwZ5MTQsYrACyIFf0m2KKRISi34qy5uIY1XKLY9+a+
ahYMscoS6F0rpiOrlznbR/d9DN9EEwMjNHbU5TAGEygqDT7D4eO7xJbA30B3CP4P
H/6srY7fftEOixY4STYhzcbGifshwsjuv99RzZqfK/5We6CmR8wyTACmZ4fteebw
4uO+kDOod0zyddfo8K2aO5di7e1qxHm0GPqtkBht3T0fnT6RhnqGIk4h/s6TXqxm
VoDUREIoNrea0IVYt448UXqjKTYfsIXF8PYCEgBHxRoT7bdcVxw58XXwq5NrZVv6
56XRNVszRu1T2iGSspTCNbkTZncCT8FO+9PILebVB1mpQrfeUaIF5rD7Ljyyky6/
T5tdsBF7ILki87AxSLJ3NPJmWbvMVSSukrhNWJbiD3pOsdJdY0zpvCOzOjl7V3p3
WnLeuYNc7dG4oa+kmpzpqRPnUzg0uY3LboCSKhY79QwS/QF4FSNvmkYCBO1ZV7as
VmdNYMEMqu75prlaR7+04Ol1ZGegRhGXkvvEodATe54fI0b7wdeSBpbusSWf8OCv
aftYBYNVQN0j7kY9sAvnSN1IBNYLzpdNfp03CNwHVN5ZkVlVL6/w7vM8irErerT6
pXaltE3vyZmTvay5tx4PMOF1tubhDiKH1war6gYDErBRGsLbbI+tJAPXx18i6tsn
l+1lzpzUFX/DQ2PXTEfHyQgz16Z3mk+FYOApmD+A0SdTGhVbIcBi8qMISbk7iA+D
fIIDqsnmC+OMUoyXtZPt8gVkvfHisk4YwPDg4x2lFvSOOTF58EYhwTq0DxGocww2
tCjzOv4QUzRAi85RMeMMlKF3JeWv8lET76090OXm68OLRlOaGKcCjhawZULrcYIs
xZmjR+OuTL+of01oO44Xy6mRyS21hcuiy6JlxxdyBcQxCSVVPCJlnRJtZq+Tc91b
zuGGtd40Em1LsuNh7Cuhwbo0VyVx2xFV4NIn7iqFZzrL419kAlZaj52+yX+P9sC3
jnF2qXo/FI+xIogR7uwyRSCOM2ALt8HQTppwzXulVl30xMxzUaN6fld8iNsc3Ijo
g9kb/JdkRwgjKBpbEnsXxHhgUxwjftWwVsBVLPWCX3cIH04mNFGWbvlo0EQRh4z9
s77E7jnaKK5HuCR6PGAn+O2DQDBOz1zEe7mIMPakFiG+C0xPoBmAmNBT70cgT0jD
SgkN/nJlG0W03wh5c/s0qclVgqFakOrgZzIVFyfv2YsPC1xQtC9mmTINFXh83MM7
rEsZLcVAnbCMqjzVX7xpYmISPkL6VR6aJswzU7CPdwhclxjNrbGlO0t9zBsfGb08
bba04BkzkRzm3nyirEsfRGjQMGvWBseG7i9KOGAPQHhDJVmRP0MXqMLQ24xdXyhK
woiqbYRb5ocVzb43OTsp2MBZloaU+xttO7xlztL76A/m4FoaGaMUKz0Omo2gXMVG
PUByR6kiEi0J2UNbf5qEsH0PFhCOaaVJgzlPFdOzw8KSKIMQ6H5CY/bagcVaQoqh
LdYfWTK+3BL6eZ/7eeBz0z01HREISSIFPGlW7pj9W5nvdPBb2BtfFdYmgECLMwG1
HyUc66PrOM7UsHTDdHHIE+8VVwfXeVpPK4djZkhaZQ7+EO2yCPqO2NFy82AIs9VQ
0ORZfUncK1v79ZupEX45k7ciPny+Ur2ZKQufLOEzP1L640UWWf1WphbcwhzSmUgT
xVm317KPcymsrczTD90VoUKe+xYuHGeOQSFxn9T9Ujq7RsBsI4nsw6cJQYD7ga8Q
kSMnBYZn1wZwpO5uNQ1E7yHG5vLZ5EwwcVDQ/9gVkANdIiA0gMdvZizLK9QYIYEg
b1lqxCs+yte7dQURsd0qRfC1qs+Jdt9El09zZDcmbOM6/34NNTPayiFfBWVkfYnO
zJ1bbF7bOaa7lpp5Zf/cdtRjms3XjsUF/12e/cjn7O0HknaYFBKFDf91CA/pMwFi
rh/LgT5SUqjIXNecO8s1WK/59I37uCy4WZc9LORBAmt2F7Dr7dvfNe4eaWjf8cjl
PQsHOL48t7S6Or6VlW9/GAxrHkJgWsECgmhnbWIXNIwjJx92BuTVwHNQIV/ghink
4ZVKtmVY1g2KKrLqVzdiWAYhnP4Epl3JdWzDmD656DMKVwyocRnUHneadPxmOR9U
tj/TVvDzAjy4I/C9K0gv2OxcanvYGJSRvh2BXs/5M/OqlHUXsxxna7gsS6KmXc6V
4tPTcCx1sMRwR4HlHiRDWNjeJxF2d+f9AVHDQmADWkZCcNAHS5vgWaA/W6VwyI0E
D7MIMFCdJOEKejzTymOXl+5668TMdVrzGp/UIJSfqsrbbGR/nNSQ7yf0eHtCdOr0
LlIYIvYdw8403hXhT/VmU1aCObsDn8vPKFfe11kMTPb4iHAU0Raw2Zfs5wBnC7qC
lbEhC40eWTJ+7PszxvJjIyoz4Udk+QIhl1/fCYWgU0TmAtfuBV5wa6+gTWbkfIjg
cmhOHDU2esiQLPuG1Rqr2xpCTM2p1EIfmGC2mJ5CDOIig7Qqyp8uR7VBJbmnR/lO
I1M1CI8ZyT/MYF7/SzmDOdZcBxmdVV+jVgREOBa6XanzHLwk4EoQ6nHmEcFdeWTs
bnL/ub/k9IHEpiEUSHjTCmxk33RRAIbqlWYDAQleqx8sO13HS2ziwkfvQOVTHNWK
tbKdeVX2ziQxDtW70VBhkAJI2WB0cqS4SR0SmNwS0mKog9GJEkstQloDkOUaNCgJ
+5aoxkwqQIb71iqh89t5bgBugAjTypl6uj4qWhiZoSy9JQc8ZZdlZF7x3ACUB9N1
fQdKDVsoaiLA8UNFPZUu6K7VhVj+FTy6fwoTw7fn/CC9VMDD4RoJ9DBwI1w8RdcD
LPJfN22sEZhoLkrW8EZfPyAWjrd9tPbtzJRzAVVq1rVsdIvvTVqmTX4Ua6jzWQds
l6hmED90AZRTMCND05bLCGd4UkguxfH358+X+kuszuNXAK6mGq/8mWLTYdRMEaVA
eR4o8d3s3R8eXCeyFpMzRIqK54nzDjVziyAQ8y6jv8vVG/BFyBV78Y2ZQTcs8l+Y
J82C4WakIc5p9j88iMfptTDEXvBImTgUD8ZZVG7g4kHalDRBNSOfqWK0wo2tthUJ
LE5xysPXc7V03+CzjvoRSLDn2IhEdjrzkRePVGZL3poIfEbQkpHpKy3DMwV/iU/v
IonhdGz/EWCWd4ACvY2KwwLgOAc6Kewd5t/71GVhK7/o2fRAO5qB5tGTsej7QVgd
+ghxRN/UmGfl//pw25ypfl0kumPypwSI/uOWKjNhzA+0gZoxIkOjQmNXFOzM8Sxk
NiJN5/Pbegpg2541Skq4sx8vmMuD7qujw7TCJpdKJ4UAPwnkSQQnICeGbKehOkcK
jMcFZP9QAmmgMSt4aAXqSA1VVMuzAfboRRIQGATGib5Kbu9VDYj/7sKuDod059bS
lzEg6xlo/hYq6K3tnNMkXB9nqXD/b6Ws2/YKAtgRevGXLs65jE7mTELNE6xnEuJB
EjVk9YZ/pmkhcIE22Qp4o6cyh5144dkYIEz1Vb+CZ8BVYqKUaJkCoRpUZhA3GXom
K5QXg9kKmTwyk8+IGTfA8Lrq5WuU/r+ZkodACt3bVU7T9Ur64Y+2o8YvQFoyi5bz
3nznexA2g+hdZ7mDNPIlCtVq2mst4GLaDgKcXj7XrtJjfU9MOLaK0U3kmDtYim1p
EL6OMwvrGwfJ7mTNird/+mgohEuvRpHhYzS8i3TmOsLexDmXa51Av+dr0MNUJF3Z
9jaytsqciGSAdFrR9dCkr1BJPaEy1G03lH6QNHHB5hJuvEg8hIIEhX4s5/dYrxay
X02GpqkZWuteQAlIAK+WL8m+MH09kXmWWV2EYgBQC5divx4gqb1l67P9LhdENi8I
bPootLygsbFKhuGz1IMHPi5t24qwd86Cu0duwhiMD2n86xOBLc+7df9DGcr5BYKz
pAk7XTdffJcYAGqdWFCuEuU2EjUwp4Nn0dUM/ERzL16XgNVV2rSUfKxqrPKNj1iS
jRUXw9Vfd+er3zBOWntFogYMfQJ2h6TZBODD6nK1TpLrQ6KHtBPblmOWFUCIE4cn
nFKU0H/Uwj1K4Min9s88sPz91KG9MiNibNHotybRjtVpM7eAG5gzINK7jNNk0Rsb
mMIMcjTBHxLI3SEYuSxm8+RnLezDcaIxGvg+nvsGfSVLEf5TgRdIf/dKJp9bBf+O
7s2vaZohThwxbY/BmiQNmkUS2ZcOXCP2M2uC2HBtglT16Py95nPUr3m5w3qkgHGa
QsrZaNVOc5ViYxb68mAK4uuoL9YXvJE3kUhiN7f8DY83UTL1xKgfksya5cvtFAzt
T2DuOOK1XhWFacZbCUfHvS7sGWSRQI3B5T5nmG7kNH9IMu2trXlTVcMnb5gpPbjp
vN4NklQ/F9aLT97ZQj8XwpgdAobxVgIyGXAT8XdvN6KpUaClF3GzdZEXfiDOiZhR
a0Mp1cYDdjkOeNv0nISajVPcQpxlYr4YrEEdKpgIPiIxI6WDa567ITEfbmDqohtX
UK5UoPtmDyhE71cQ/Mq3MsxU2PMHFtWplVnDilpcHXiQjVuhkcZSbH/oGi4BB3Np
LYyghPpyt0ew2waqebNXC4jOKgFTbLjXf00MGSBgbAx7qV7j0jAJTCz0u/ZhLvLS
P24QA1CQZyooR4iZx9RecygihB0Xz0K5ShMoIwof8IPL405LDaXwPKyzEOKVaRlD
z3+mwcvpKodhYz4kG5FQkvRqaBLMUByvMs8eoMpvUaX11QW2z3+aYBWiRryit6TV
RID3EBGLDevEGIN607kXkKow4c+Ywj4ILag2gTH8B6ya29IfKPQhkEgNHMc7i/KR
kLLu/BJg7iMSg6ay8/fK7Hyy5WvR/xE4qswWmFJl7HmZsfdWISwzj9VWTPgKeveq
IiJgNzJHtQKYWhsVWm307XunmDRLUZrTQgiDoswNpu9H2+S/AVkO0mg3gXGbFaSm
vHi8DQ7VLUZb9W8ZrNQUcihx+H8VqK+aSjabKPHG4C65pCvRJsyBfO9S90TPx2HX
oPYvRdENCXp2SUGX3czB1K3L+m8b9y0UnqvMX17wGqP+dT3iAYr4sIcD1IXoIvas
w/KRYAOOGlbPuEOzsrxxQFC4uDN9py+2DZ+Y5ZAe1Hwx9Nb0kux0Wtm3Jbb7kZOa
ZFr2fLxvjcKoQJQ/dOgRT/sYh0xOO/DjmHnvYU6xohyTa+/HIxrFqgx7pDJOoE73
TGAn1b7sLwdxtgz0hnj4p5WDOYDGlk5jvZUZn3idoiJEipLK/0deu2dPkhJugzUK
IlbyvYorJAuDxjmwx3f8XR3MX5t7yc/TuC4xT0KvAteDTxNYlSL1sSHOhUttx1pp
jkT4g6soZpcgjLR5eMnc1c2PvVDGhebEDxJa0Dl1LZqYPNZL2T2R+1bUOzTMBW5L
FclaHVLseEvlusoXDX7St6rOHlj8MRjIwmWor9UKE+VHTgX3gjX/rCrDIDG6YsRw
R2/K0dWSUwtLa/4dgf6ij+UugN0l8aKI4fKExNw2n4GaLQ5L12KxCl93iFN+pH1k
adfVF14NEns38IOgyzhZ0Q0qFDXFORh5+WBfk95196PzhDg/xzDBddK8x8WD5ZxI
Q7cm+ZD47tr1sv+PheuphlWUblbuq1Z1Ne9ZIpCN0wWFi1G/dpi/Y0RZCepkxJTL
AFG3HcOJdMUl1HzNINS/2JKf8BroQiZ0g1XLARaBBPsOjElIrVBmZiwyl3jwxAib
f3VXi/cx3ItznU6exFL+pluFPpjldQGcYcfurvcTCj1XqI6NhpeTndJ9NrpJSVQ0
ZcBfrtb/umJyvcYN1OSvddez9WkvAeGUGunZyjJ7zV0yrvbq+hYBL7VjJ5g/sfEL
vYuJ8dfop1pHw2OJev363H02ifg1YMzmOoy2lqYDKfcxh5N4N+9Y+xNDYQicURk2
9KNnGx5B2jfwkKuWLuJf3y8XS6VuYqDPMKDwB5IpNKBFvAdBzpHFWeCAsmzQLf0O
DWakiICsiHBi4ch6Si/RWWA18HS2CQ0j0zbbcTQU4nqpH3nzD8dCz1PUA2qp/7ov
zpYaEvaQfJEysLwcooAGgZ9Nw9T7UrZWuQOEnCP//NPVF5eeWZVB5zcQ4rjLbFTc
N7K75bGfYvPXN5xecE5VoGscmxR0JP6UfL5j2HjZvPo0a+3ZGTN/4ZuLOrNDmnRQ
Ne9U6kRJxezUPPF/gxDIH7keoa/4v5GEira9EdPd+IuZ3qOtWDQpGM7zfARxznoT
aw8XFIXhvDS4PLIv/7iZr20xSeRkG7H6hAGDf7SAc9ZuOOGl+44ug1u18f58x+gE
rikaCUkYACaz8Zh9AlFl1qMSR/dCHgCdepk+KbAL4cwf0sutLINoBAoJRzbnAs/N
7SOOWkCgcHlVxJyVlYMJ5E+y4MKaGVqHGT6JCAKs8+vC3iAgY+Vk7k0h+zimcMEB
itKhezkdKjcNw34l+ZOss13kFwI37naLWO431Sy6aoyvTOl7zMzlGZNJKTYOzum1
4enykpsl8mRSI59NG6Tl1jTOccU8l0QldoAeKtKH9eTNC4RRKx0Ad1nxtQ7xSjXo
RHNSRuZo4O2Se9KakjDNjcvomiF2TGYa0UXpZnrrRpK7D7xdiHmYw9l+Kl2QOlra
BmZrr8yM3TEF9mA5g4Y6TeIOQlYbt9DfAGue3xwdgg95cbpNvt7ZS8+tq8L0RgOM
IasTnR5lgKQLOQiR0lgPB5SKzW5RLJXCVlGkXel67C55sKv5Nt6muuAoTHx1JHm5
f9OtugfZAbzJrMYvSkEIbCE6tua5LT+DhuKBV4ejjXxVSfluXUTgd/F5uc6dHXdg
7AR+tKmClK2rQ9G2dvEod73DwdnLl87NP623u8NXS9ic1SAJPLo23DZW4XXr4CVo
K06DLkextJhQaYf4u7pGyGpiXnppXRQdLFM6JjYJD9+s5EO2MCDC5p4aOc+L14IW
ZPvZvK7+fAO7bBKbCpLaC40o9ZE7rZUKHudZuQ+3KbwH6gXuoLwsGhjomG1UHT/4
ptn/nyBZA4zGRhJ5KQKHDis7TvmU+FIHuzABsrSsmzXZwVOKsWcqdxN4wznemTfy
DFPUkMyUk48kJFPVcKAwwGaUrV28WI1CC1sPAjXwxGUlrtH0AZhLzXVnk9tUoUnf
ZQM9p2xwh82Be7MTtA7MTX6tje/lZ7lKydFmCTMRcnq4FFD5LHWOm0HdxgfZNmym
4skv9L+J2UYRh+6WfbYfKpEAgKPslEcP+4jQ66ynrwowbOkYuWErRM3BkIm+nuOv
QPXpLyMg6bJ74zkt423/KmhuoztYEyYxUycmGl76x5/bxyqd2r1OXEqocbHu4nRF
zqLjFFDlFb7cqZ4LA++/snpYoE1+XJpB9PwUjtYt0Mr1D7TGzzoarqNVh78N4wxv
87G6iEKz3Ni5g7me90A0BTR0/d12jC2ykXxC5SN9bih8jGO/zP3GZ8fjO6yvcmdQ
hgv/7DoIN9wknF7ifKyKHL7mPDzmd6BSvXEpD5petYzHU2CCCEoQreNuXDQOciYt
fGDpv670IseG9SZnCIsOZieVMyC9Q1MwBWdBqIAaf86VnGWI1Jzqd3TR0WI4d7Tf
XdVaTGXS5AfMBxfHJcXM9g1urUw43nTOn55oLzBufdzVVGewmiobXedpJnhG5cua
cVksZTRQBITanAQtul72d4+g/LlKbMlJ6Rz1b48+b04DiV7U/DKqDNjFYtsm8pjo
xjOc8rdfv7UG+TyyTAh7wkyCoo5pT8BgLWDiOxXy2LhSvfXaFnpUD97QWrbXHiUh
wWTaPD92abuth7Xrp0A0c248qOO+10uXlSlXUX1Nhi8QqSiMqZhCVtlUGldkPyHd
rP+5aIZDe8RGb5uJ3IJX8acAM1EFq3LhEEwLyVQfBeyYbWLTWXVUKByLPajCMc+Z
UjdFSHi3F1FnigypAZmHmShap4j2WY96wjXJBaOQs2UPbhCxO6/xuUVUdqXg4QLC
95fwbR/4hllo15K+RWS5b6Bon007Xcm3PSfkZvwqSunffx2Wt3CRODzq4uwODyK7
K/qhweHOkRXveK1owOinDnrCWjlL0ak6L3SEd084q+mGM8aPcW9xpo9HDIgqmiys
HHLhSXeBWY+x+bU26pk+SgrLF5SKvRSkuqZ40jboVfjbAba+BZFNZARAvbuzV9km
+leQtNa+NTlv166UIfhnsp/x1n+XJbyebzxaABV9gqkxAIRC5D6YUAJOSuB6QBn6
DqvSR0++LbFbY77JyVOlqBcvqS+raQEVakmpMH+nxeMW75QQfKwZcX1COGi0zt8D
ZADxKmr59KjmECGPaKwOaLiKdlAjRcZggj5Es5Pb21OYSSxXVIUv9ggAEMqB//wW
hievT8wNuFiEv97rMyntkEbVm7Jxmn/c99bNBk8EQ0+PqmeTE2n3FffOzZ9qc391
cxHOvxd+ysSsDHHC2p+KpEqM4cCIo4JTjuX0Cyph9dKF5M0B4QCek1zlD968ySr/
tivbd+jcH75wySPUvHpz3eek1o+p/HT2W8W+VcLVEclZKEx7dEaRS9BIYcxTkoni
NnpMJ/2JyiNf3CjY9piQKFis372R5YEfScKYmw9MID2DTVOf76chzkfRnn4wjaMY
UvD3aHaJUPkeqmcRNWjX+EQxpgKMsy5JuqKD2x9/qOq5o6zsgHCxfINwAz3cjq0i
g6Eo6ffPbxhzxIv3IZv0+KTy86f3ktuqxl2pCrp2hkCFzFIehdCrE+JOFphJs3GK
Dgtujx56sHSUnN5da/zpTIHZgIiI1f8xJFtREdA+f7ybUzN1Hnjz+21WqZ2ofpYd
TCtG1F3oufEYlUOc/ftV3VDVijDPAyMPI8BZa+Amghmv+pqIosvj00EsqilGpc+8
ePCBLCRfp4mzZy+VH0UNZ53q8cRL7wQf/q3E1hCGSkG2l+HuUo5GQ3hJ3acsCUu7
LMa4GKNMs3GXesIkNqAUkIrIa2VfShR/4FIj7fd1H2U+BJ6PVVmFGIxUF4bTKtol
P5FhFylP5jRlCULfmNzJWfEXN5in7u5Hb60qXdRsxqpg8qN1UiHeiPjVKOksuT47
VmKlngEe32G7zFXJAy+b7vlaVizoxd7J2HxMHE6zKPOjQnNvPQk8MW8/EsbCgKcu
mxxdZeJqQkpNstICITbmAuzHjZfKU0YFTzzab4o9sjcHRcJ4infDBIiUGAmkShnI
JsbXzBcQDHAUfrpOaX1irsZiZYA1Qy3IA3fq50qXzXQpzqQttV04O4KCL/Jm2F3j
KxDLKQKqAvHLDSOotwdmSzwLo1w2o8j1GVAHp1otfmIoPmFe58w2UaZ5FVe4xcEu
cNO/0/eouqjL0nEUHMQVpfYb3h1yH77OzcuZY2q5ouw4l7MHK67pB+KCI4PSFoFA
Wz4a7AdNg856Pr+5Zp3LY0hWO5XZ1GPjaRjEWLqMiim+6a1FmKWB0UO9GJjUtJnG
ICIxA0DGtVEb4FUD7wNWa75zlwILv1NePo5FO8xFnRYi5hAo+nL7rD2QR3C0rpxk
X5Yz8UipyT2LpmsdlLyh8GCyjc8ZeEc08DGG7qwvbksesvb8axxQzwUvAu+cYDlf
bMqAA/KAg/Xymu04h5U+lozVjRt1jaYzj4VYulQfyonr8M554VdDATX6Z88462UP
XWatoIuobTmJuPmwTHLcCz+tJzKB2oYN+z+nnTiDLGcEh1GPS8khXfJR+g/+3Ejx
34lSVJ6BHEoPEBffYM1KzGRpN8TJhLyFoS8XEYNfL18OiMMOMHLOD1QMW3ZUK5ra
Bs1Jsk7gSqd0sHibnZI9NO2chSSRY3MLmrInY/H2Itfv60m0BxydCPsPDH7opAEX
y9ccA9U7IBQXVEzcpVciPHKjlUvLCBom44ifB7a3heAnDw3+K2ccHwYVqZiJV38Q
GNsSg6BiDnYp9gjMP++UtoP9RIF7pCRTafU+AJ7x/JcZEeKG8/pfMKUpgaOg6JSc
wX7ptjzxh5QQ47UcldO+wS7lNxrDpeOXKZr0EOqYlB8IvyDn6fJgcenGgGX4dpIr
C1GMiwmTJX1shLLyjq4UsVB9wZLlPaIa5ok+pbumUpvLc1/ixT0jf9iFaDoogFui
nPRPJ5DtiDQEkD3FDKgSG056s7zRnEjBQ5s5pQRF5zT15vcHW6n6LwPjZZCyVpQc
5rzNaYn3qxO1X8ban2y4bw6T81NUfuI8FuCL6Yk+3zHilfboztDzo78XnsMaXd5d
Oesn+1BqQucXt23OcoWl/XLDTL0+mBGwDRtCUAZp/IaSqmYCbQt9i0qnu3hUuv5F
SX9G194T7NjyRbqufzEOfI2yec+7sQyatkisQ9hR87QB8XmXCSgHSh2PKnbh1X3S
fzdnHWmybGwcm/AlEoTRKmgDYqIFevQ8FNM+FjsCRG4a0sxffaYOK7rtrv1YDE3q
ysJmSttvT4FOqgCPveHR5IUZHOH5HiijMVLK6f1cblWd05myKHSBXLKmgxThEHsa
7KgMUxYaUDZWwFaeUkd23MYr2gnQm9HR5FQMk0y4zoWbc4CQ4htZsqw5UUt3iNiD
1uuXOyeuYN1OUR3svaPHPDlSOxw4MDfuD2iohfGasWF2RLLmdibyzQOhPILHtlvu
klQ8xU+IrXzzcrEVOno6oLP6O/kCmvu/13gSbD8dwUs9m+GOkfzNowpYzu8g14C9
igglhPyGAQ4K5FoF1F+tKChrGYgYpSdDJoOgKgT2ymejZ2DJTPLFhe2DaESeNUQg
agT6TURTYjpUdN5FT+6pEwfPMAhH8miguJe6nNNdJ7llXeiQ7w1Va/jKiD/tKmhm
YSjupirP3/WWTJ+BnnOTgBTn45OoC2PvnDfX7lG6UrqfdETuOO5LRQX17NIBSM5c
4/T9dFVI9RNv1srZ0jMsjtfZsvi7qWbVjTWkB7G2wMDzyQd1Of5Srr6GDaoZTw2b
w+q5J2gtqeHOZN2b/ESzUSXgDiDWeoPVFPakZvlV7wCpZv+fQBd+S7uzT6QIUA6K
cqQAfEUdPoPiX18hbDk93Q==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Sp1mHkiPuA9v23gNsuvkEoG5xDxvUzAJgUaF5t+OjKKWyGBPFhTEk1nG4nkGNj+l
ZLXdttFcawCdLl9WXD0Hv5YUulMt3pevkGtUXhQ42pc3HiRpp4tw5RKl+KD1Zn1a
KVCS6T0U2Fhl7ZLt4Fww7G8h1XVz+Y0nBpn73NwV3dIctespR7lYKpwfWhhOGqqO
R3O5aTc4/x7Z5sbS+0hMwMEm3zcxxWVhPVnbp5NqEJlXE9rcP8WRoB2bWV/3xlre
LKUVu7DCU1jJj/sVKf1VuW9x2pmYzIXyIDe9b4f6MViDRbzbkEJCVjLRhazdMsAd
kergRQSqzj+QJhGlLrIoXw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14640 )
`pragma protect data_block
gpCIEe8oQgRtJ+U7o5WrF7V9Cnoqt6I+wyCyVC62m+16SuFjnJsn0XynmgT6cTDN
RhBacIAI8/2qM8kNbOyOr/J/TXVMCpzVi+e/4OHsK6XAeHcfv21fFbanPpoIkzt0
auhR5/jKRXT93ZRqI7urC09qm2YTOcCbQWAajLYr4u1e8AojBmgRtjWXPb5nIDCv
DJl/XOu4pS6bxAr6JWVlUxJwlIR2gzVxVYDBNA1hzdarSf0GcGR9XdbEGAMpABpu
blJf8LC141ID08jEyKAZKbjhePAFhiAPT1hhQT/+LXwnjiMJJ+B/HsQB5KsAtVLL
q31lE1+1r4yEjjfwiYgbrzmcaGbSvh/8vnEvvJl6zQrOU+d9W8rYEVSNY6wRpndu
R4lgC4gRysGVMJWdD9wvENBNBXxNX3dlpQYKAKAhEKDXvhdAcICFY9Q6TZOrhNEb
eyt8cz9SCBF7inLwxWY6zlfV7Fb0vyPU+9lJxdElgsDxbQTSpi76uX32LfZgnaKf
8qt1/ZLFBSYivrpI6y5/CEnuRurIdhCDaRU7azsKADl6k0KWeG9uMztyUPmjQ0Qw
XWRPlBFqyw//Nl+oc2w61wQOy44urDU8YaWdJyFnF/6yHnJCfmCiDVXkpaqE35lM
pQ5kwe5erRP+b8ADsrF22GwlrTrqzTEG/EImqGsHJ3GahSmE+3H0r+tMCxThY3CQ
3hc29sYb8TXisYTCHszAjKNryEX5YwFtoNXMoTivRBNmyQCVDTU7PIeqMpKuKKpC
w+1zMF//qBWvKOx8Q1HPg1fqUKdZJ18XZJcsvipXFBaAIqMeDiDKu/EVdk+VCLez
5IFQXw5vbKwb/ebakvXzaO/EWutRofARGrgQsRjHCFPHELUHWSqI8OufiaY+RG+B
2dmvasYLYmvK6llmC8Vubq+qjQrIyJ0ZWzLnE0/0XPwHEgVuYsp3fTzTX//V9jL6
lBREBJZ02W1fJ9DcC6A4t7qEMrdXBEj6cTg36jug+I68Mrm4bSKrWItKsPgUyxoC
DUUqZcLdfhsdnTiJ0s17bZ9H7btEmdZlPR59VbM9gSURhcDN8CTBuMprAcJzw5zy
RF85AeZOmV8izLwaHxIu+q+UWy5eZCgw1BoEaRpSW2DzAHSMC/UfwAelxolDYesA
DOk0QVVAIMjMsE/BlhiMYGFmRBP+oWfBfTklyrJfGxe4yVibwSAJYjZLZO+kLXhp
ORFF2YeOgK3WETdb1v6W4RGZasp1HTGPr7GOHSTdO3vNY9czLNwmtfm1/k8kwWI1
sJ76ivS5zfsuX8XwnifQNGgv533bvmaj4LGaWMQGvYEsVV2FswLbc+9jW1DoPftu
HqiLm1I8ekhQG6K+iRko3GI5VURcfUO7iwHvRrb3+M9/kKRGF7SsHJV2s4EzHTbM
gm2lT9qxcApxqopn0UvnLayeYObujIoBJrMRquA5RAu5O7lA+7rtBknXGeTyFQ9E
SqfVDSQFvx5yBJvCi9Ik0+kqIJ8EYkWFZvcjmVRDAABxcAS2KKWr+rdRPewyhC7R
rkwkKg5Bs+v4qdB4cQCns1rKg1+6TAE/inhUCTYcZyZVT9gXZxzVdolkEu+kJ0c4
ivU/Uvs22IE+ovAoJ4QqNRh4FmW/TLHhIiQg5KEbBRgcW4YtcepZSNXRF8SoCO9N
7g/iL0m3H/W9VFhdvBUITleUHD/CErmEp3xYMu2Vg1Zpv3OBJ26CUVFqP0ah+ohc
rsyJ9FM1w/+hL+/QCUBrqx5zCtk8B1IOYNkcJD2YGJq+CpM9rAVawCpvhzznhUwq
etZAo5UUvoeWlfC4Y5vKA/N3pxYmhCVJzQqWn2Bq0I69SzAZ1LGzeXCVEykG2PQl
0e/BbHAIqtuv6logRUsCng+9pNmP3R/Yj2i87STRjAxtyO3Dla7es8mcEflCsXc3
zYurl2GXVTiVN2pWzzIkqXAtG8zUmtwhh+Wc5c7OMmbnbFomHecG9Wo3x7gqfogE
xDeq0NchEbD73tdragX5MOSExdJvdjgew+gbUSWemVdMhqO+4bSAHwdtFtwOC/9f
CPs0YlOfTYS5yiwSwuBDo8PUFkSnNeSpoYNuU9vGhLeWoRLHSBBli/qHo8PKltRj
Ddv7XSx94h8WqyxYzmCosUhajlOuJkvrRPaqsCgnrK0+K3GHnmCN7qc5L5KhT0Tb
oUatFKLoWtU9zCS7EU7YxRDTKj7F+QO8Hyc9X6VwvNVvjs4a5QyZ+D9a/P99BDdg
Axl1cugHi8bJj9iUzVP0qFdIEYyidbj/PlrhO9FJ7B4B1+gWBaXGMxIdNv81AidN
szJzsPaKp/6sdDZjMyG/HI+UHAufuCQX5TNB/BY6hVtkRcju84eecOKQ1/NfidOl
wBvmyZ8RbbYc59YiNuRfJLuSJWnRmfmoIIT6xKMXktGeZtTSAcwWN0LIhYZOGMIc
UTYZokvPaufqu0A8JCNyUwPnAWKICEWHgaQAEUK3wUtg7jlSiBiLZR5Zvhcare/e
yUbLtoyKxWkp7A+ZODuxmVkpsSWsCkYGQbVpAaGmdKEKvAYKBcmdJwYh9/x+iCzl
0G5q0tt1jar8IzybKmbLAOxslrizanSXNzr0NKyLjn4NE57AHmZz3etIFda7rtwl
0BhKcU7CzGY2M1ZV0Cm5ZTiHchDCxCtWBRyT0KWeeGuTVQVmzbuWbktFFX9ZQAlP
fggnqtSY4YngQrFhGFuG33rKnAFybcMXNtkEiBCWElMFO9wT3h3nqnUxMaypq00t
d6IRz9CA3u+oxRPe/vdO97vrV/5tUAVJ1uixRIP9y3teM0vodfHrmDrSAYKWFtii
Ncr0H9+0o36mhYeoDTrxTr2tSb0TN1To9GW9r1oIy4hlOD5ocMAzWf7Y6xP65FF5
IzpY7G85H0hs0dfxwkP6SyfmzbT/wFL6ZHH/vEh4lT9fvefuTQpeh9T8chhfBD6P
LtkLD9RxexOcQ7ogFsEtTIzfUKa2ZmVMIJ+82YUcsVy0Q/tZfPwOBCUjg6cdNFv+
WTIqZLfI37Hj/G8OPBcmnU2bS3HvYSeoezSZ2FVaio+h1cE3ObnQgfw/a5BqylL6
rht++DepD3B5ioJhpq637290arCrq74FyUkY52eUGqzt/94p8NWr1X7Njjf4QFa5
+AaVAGURoibjQ1gMfzB4ljxiZfmrU752Dp03dhw7rMPxHc6dWr2npUZP28y8m+Ps
hKBRhD/H1DrQenSDe9GG5mtHUsLNLLVgMlZWiUIWarkXik6Fi08YhOrz5zBxnwAq
Yqv8tLQrQ9Xp6S/+z3qB+x7XrHSQbX3f7Dcv9x8yt8j+ZQzW0Qc6JeiWcrlpsMpr
TgSFx5TaeOEXGTFBHGUVjeoV3tLQ2oCWgwwxgl75M4/rqvYaX6nuAqYHxmDqNwlr
YNUbHiGdJNqx+7SwTkzXIC3jkCFo0SSoCfh4V2XD+OhUaJ8MhfpNVAzBhHHhgX9h
b+/Z3OX1EJjxa29Z1KAP7YAuI7cEUHGjQBD5Yo/pSMlWhZ8qKBYvovPKxfm6f7Bm
ln/VLTDbbsfNa0lYF2DRYi+s0KieduzSP3FIsf4v+/CjqzKt+e4k1ODW3femXNHS
FvS606+nbvZSgu0v1IiiMo1CYid1cZVSNsDasALvzF2RL6pSOhiANu4jrQ77DIq8
pDAbCBtdEvv2uva3x35x2z9iFBxsI951n4a5Ia5Ks/Wbxl9XEzP5Yzv1Lykjy7I6
1Ps3GIYGrXo9FaNdPV+Q7iTLog7fPmZ74LGRl5iTJhUFraKSAKFP8o6ny5t7K+7M
xrDkGO7ulNu1XTPla9yYATOj8DDy3MSl/Jpw4r0FXogDq7h3mfsLRjYzk5G3cGQ/
L6oqR8DOWL1sfyrsWi2+rEQ5RYyiq1vmbe+IL1KjyyTc1ZLdoW9aitFKwjOP/t4P
YgIXGmEYQyxdkOyRW4GotVKCKCelupAuAUCfoA2BhCSOS1/ExDTgZ/b+iEMHCx1r
DWi+TeTxxAez1V/+i0phZlezPbuwRadGBm7IaHWU+VyLdiP0FZgKQgrtUgH3Xi/R
HsofDRFcd53+19GpKk9XmuoW1CzsstigqCGFWmqAQPVBDLfuwbyVfw0Ln7fcpm0u
SrJqyAJGa04MFpoJ4BRVMIoJyPv7HYCpd4aokZB6KwZQsYS6QmXFbKFqGh+cWtad
xv1dK0VaTheuenHS5ZH3ydrtmFxjCYgP/9lc0ur1ofgq1ioKqLhR0vLte4bxd/P3
YOnrEHMCM1318eP808hkfzWBS2N3hEBqGr+KTsO5dMwIp6QFQMPEinIdNxUlEcCn
YccJQV8PLwYEX2zx0Fz95GP1oJ+aK2TeVH+uHv6I7wZ8n0tjrT5ZSpEbLTF1auVa
qPFqIWF9RxsUEeoRXcZtbCq2sjGIszEFz/kjSW4s8ciHH+c2swdsogrKXXr/6bb0
o0fV//lbtRaCPPVQB8vpdK+BG4PwUHFK7CAQ+812M1ihtPReD8+vvrel0G0OEPER
MVkBJ09g00P3Z1q9zJ9t54xI3hTXGr7sylkAssM8YPHkE3XTfOTbikq5uZ+uqQBy
6AGjPAzqOofCYsiYKf6CgCCUnV1SS9qPE63tx7lbvUH1iCM3QcaUL9bX3KB6Yc0K
vitkFEm0t/hnp+ZVeOxgZx6079xuGkNBJm/xYSygqkVkXnFpYpEUmHw4nI9WNntS
sCeONAPS0kAlj1SrXVs9oePm8ctAQDONfxXG4jrQQR6qpMa2TffrNGaBbg207uyQ
mEGw6ZtdXmeWYLvk3t20wYMjQLFrAhtbOj3fEkpO6EbNN9XEMAzM79L3v8viQE/l
bUV3iS4cw1i7O+ysQCITavyq0q17NGvTZNkTmbA1altBPDDZWTf9PaMGV86PhGSf
zFThdZfytRRrpTbynU5O7O3lAT1eBTnBAL5OM2qQY+n0GFRCqPDtLrJvN/yJUzum
BkWpefUVNmivM6AMtJrWzZG2CrC68p1eQXx8T4qeumK37zFAq+IbAwRGUAx8Fv+2
XHbaDay9JWjSipnZ5epdPaDPs8VJCNcRkfSmUnqUC8xHXHo3cZ3xIJB1KnQwgiNF
y3W/prnktkU4+qn2N82xlraAIKMX3GBFTr3wtlwalmnLGslRcm+Yl+MJ918iTf6d
t2CY6utSqa+8grNdaMqhS8X6gjzgqZcyiRpEcSFK6V1Ggrjvs+exRvGpzbbbuuQB
8rjBUAPrBwL1dCM+B1tK9fqS17hSCYrrWQT4fhOY1acsgbPF925rETzFvEfHMYjE
xKUl/ITAmOVNhbzKDBL+AbFr0pMwz9MEyy9l/hRpJfJK4H7+qeIxca/TwMETxOt6
c2P1l2dXZ2jae4Zs3d6m+CpBuyZoSWVZ4IQOfrH43GD0/sol4n198GU2zRZYCLqE
6kCpWOBqHyiULqIdBken5jfJQowltqpGDl0IlSU3PHzPYLitR2OEtcalCaLKZDQu
Vm/zCJmOrTelbzhEU3UrAkbzmseHmgZ365J6+Bub4BjmCMSguWJhWhkQtbehRhn3
a9lOG5SuESO62AeckND3NHPMf5gE4A9Q+ItfjRGksGy2K6JfOrGB/nKPU/5Gb2D0
z/mSXOiRHgqnGdPYuuhL0EpAilRj9s+nXwmcKX0pwkHVygw/CXaZ1F7a0pgWnKv7
8e3Gwbppw2F3AaG/Kj4LelG4H94rNOMCcny9fqzphld4oYy7oPIjiUyPae0OZICq
CeL/nMrcHLkk9bC/+GJikKH2DWE80dsNYd5Oa8kp8JZq6WrdhlhedBS7+d1ApATp
cO056LtDYNdYkd7H+Wq5uneR0l0p5BRqMNQq2ERUP74hmE5+lXB049K8PyRfN+0s
U3I0vurM/+k0CTe5YQgwn8jZpM4xtD9/HJIUhL/EJzYCcrMJJ2guBpa7N3eQrxBU
JVZsGl/xmXldqRn/ZOwVPP7xBZqnBtPsJUxBuOrPTfZIBMIg4RB3F7OEA//HUIqg
DqAIhYzw3PwV7MlfLxFkB1sz0IcpUSuX67rh1D+UFjxWeH95kMU5aEwpHdAgyyoF
z43qGh4MQThAyMnTVB25TSzSX6RIRlvIU/HCm3hOpAi39IpYyDpNANU3monUHFmC
6j05fRm0dJ/iD+Vf+ZF3feiNA7snQ1BKr2f4sD1vCTU1X9P0PItoyMmZUohYlAqW
mLbH2jdy9T0mcPc9CCEFOjiiwrhbz/a8BduEAXB5JzRrEP72V5xCbqWEqq6FqG46
jtEfLFsychk6hh3sy9bHoAvG1UVsoxO8sn45qzh3OSaP7UQQKwA85yPodloyjADf
hZu30GcJleI2GwHO2TSfMpKpnASnS5pXFSqFMkXkstSm5WtSmPpUrrv1Xs6RCJ4h
TfyKOx3w2kiYX6KCUcg+bRGm52rtTt2LO04OLMQ+CIOuZdS8PmHwGRbVHGzoDpzd
9xDijIaeeeWAzIkqefnwEFmKWV8uqORbNSwc6t32ljPUkj4f0pOzqGgaCrzmJIBr
WvCMoR+VCHN2W2r3kDydPPZvfsWN5joHUfRD8Zy9B1eQVg+d47CV0Unay8Af+WOp
XV13zmkevfmlWX9uZy7ABJJHe9gCCquQX0yu403/Y1XTuIB8K2E2GHrUiZw1rXQc
NC/2qxSwxij7FUg0BES+7JgbQQI9FxmgK/ZhVdo9XecNkjICOsUPeZTKm0coNpA4
Xt3Y/bYyMrniShVCAS1F1d/wIveMbD7UXk39I2vQBCSAIsTsw563bV0893Hn8F8P
xsoXo2LbDi5uxaTBPqnJNxisC+jXfyzQETtE33pB61PF3Eu3NbijLDC3Pp4KRI3S
oIU1FFRo+4GqGSQb7Fwahj2vUjIemk1T6wlfr/TKOeIbKTS55tpHwe8GOTJ8YVCE
EfzkoRGkMcE3m3KJG1ZDA1q1bRpj/B+Jh3TngqhZe+ZTT7KVR/d8a1exB0+i+Uob
QE9Nwy7r+5amZ7sqC4cpFMCiaDamoSQfAc6DW59VdCIvdY0Bew9SJAsUvW0uh7Id
AZRLKVAK0shHFzNVpwh1uttKzHEBBCLXzWo002fgfhXBP4Xv7RwLxwhkEQSm7D1A
lmys9ZQETkinNllZH7ke0nMYyRjmpbEpql2WNmplpl5ggjS8gyTzk8WSkX52ElwV
50rfflmJd5VJo4wSoVt43LkxGgJ8JJ1seEZfHc7llsBm1KNxU5VCd1DJvi1AILqO
v6qTZNftw+lE6XX8nEjAeUPf//ZPq6wVviuKPKedUkg6kAOfUMuPAsEF1jBIo4rx
tABFAIitzrXs7WKbTbv0IuQZH8gl/DfzmxnzX8c+d0PUW2rifu5k00cAX/mPPEEZ
Qa61Q4CCCbX79YFYAYUfm26K41s9wd4axQmKkujYAYG6F1Q+s6W0dfQpbKYH2RaY
vabnuo0tFaQC2lUPPMtak2ZFrVMxZRMwHzzkuYY+ei8rCH1ZofoTfCkSFLAnKR1T
nCrOqp+Z7j+4IT1AAnpcNwcpyDm+UMFELXzGMnrvghEeVqM5SsIFjIR3EVjCREg6
qyI9fjw4cusgvlvvjC/hH6rzBaGYaxoD17GkWdQ9mkYQPVHuXwJ93aTOPmNptTBH
Fkl509cF3WpS1RdSEogoLZx7IGt2QEzVwnZSbO9nDOORsRQfkK24yZZM/JlqHiQD
TDxXP4ZyA1nrfwR3VoCEpSvlfsaYZh7fX1tCU+RNAvV3pQnBIB3+rj1J8dxvcQ3M
gs68CW2bbOPwbN2AgVg21N/y5zS2ryEFrKrq9rt6gudu4VRSx8WHNNu2Pud5LvxN
XtaTEjb4pKj4iK/RALXob1WVhPg4POhBqZideOHt1WWV8cB03DTO38bdDNcf0kt0
jr7i1ejEPt2TqDbp1QkydlvAtnS5ZGQebC1c8h3qik2XTt/pAhZyw9aowxAmB7Tz
Btv9s2ULE+V1+OzDYO4ihtTDGX/V0MM8s6jhY4KrGkyhGX+bRokx/MXLRW0MljXK
sIXez1DsirMpgiNVUbBFj3HQ84MCBus2Ddd9askdDwwW+saIutCRIL6tPJagPWoj
sOTpTIuOi78XFXfeK+xabUFAMIKtOdw72zJg7RKLgb6XFev0ZH0qXpwS1c2Nfgu0
ERj4Pr9DnOLMdiJc80MX8S/5lxwNon6IKI9YaNg5NjVSXTgEpY31QUxGWx5tJN/E
aUaTSwdfHZZ0mDlZ2GOQ5/O479syBN7T+0EKnxDRewHzsZHVEnDlOVkZ1htNXSPS
N/nMpM+QbbsAgLQT8xm/o2m+oAmwGl+ojx9vkVPWafJGTdMadRzIZ9YA6yJ+3Mh7
TP7ybWa1pFF/xVFXSp84sMFe6StIXaRiepOCtnXKnsIJcwquNjyZuFZUrZQfWlZX
QYaYrrXvg8/hgREulp6z6xKv9v9tymRHIg3HOkr5Cbarm02t2flkxTonXhiykotv
Vpe5aMDLXj/pXMWk8qjqJvz7PXk4Pm5h5vCau6nnaXkP8ss4JW32V42D+NJ+KQYf
sJtJDa4UoH8edbz+qqWb1XVIRVjzG4+4fA49b9HIVJPnLjG8Z1oH15r3dV7r/SAE
Y0u6t4HvIAslbky3cpO46mLmXWgXRQil5jaESDvgwpjMIwZc+IkqQYWB657nXv0L
5RTGpDqD0brrOiGQy3Cbvg1hJw2KbxiZ6H3BIlfACmTDH/vVV/Ca5ZMJwVJgLvhu
a5jonTpyv+A8gyxuFZJDNsL7aPL4z83e8pu4UCTN31vgM9OBqABraKCZsRnnv1Va
l+r8NvFvQVimu/T6ZqP9jZ97qgjKVx7UmRvTxG0HeHF4DxJqZX+2hHVBMqcsg/Qn
u5oS3nR1hOGl2AblrQarjYn2Sk8P0ng3o16ozLmGKBk9IGpAFvo5XzarC2inNZsk
07ZkTsWyIV312IdNwJnFWZQz875YYDC2aWEtoCEpzw1JCYA9nTTnbgL4dEVbHZkL
gEfNEOpdymicoSB3GhujICEi++DW9iVa7QqIE2H0+3X9HaE2kb8WdlRbXRl85kCC
twfEflIxQ/rxqOl18aIGlHRUOSLMP6p/d1TnuyyZB2TiOsQlm62CxyvW3z4+mtFu
P5s7ewlOEQI3fJXU585oJYlBvGH30EY6rw381CXlMf/ewoN4pBVazMZlUEpBmdsy
If1tHZFj26WJUsalK2232ik/VsAbToFZ53PMbXhlFFIoVFRr6Jgm4qBxS7JSHQ2M
kcaf3unM2EZqnoNNGk+bBGB/nOFfq6QHtuuJYSCwpVdQhai78BC+ffNqjamE0vAT
zMDclVZykEYJnnRYj1dPaNIm7cZXXSxjGw8D/gkA5emYDNfiFfDi8lZFfYd+pSP8
ErLsQofdCzVXXT8Nyzk6FKx2Qh+1fuDj4F42zu0G42thTujeIzshLJun42f4hHnj
x3CBVgZpDrGY8+2xyEl+BDvPjo+3AkXKhufIWhk6x+GfjPMdMDNnnSbgldPeocbs
dbWNovmYo6+8RTzhu9lboeN5DrhoB7lVHoTPVT9zHJQ33PZWLKcM4qTKfNsVDUyG
Wv32YedxoNW8SbIfrZhzrUA5mkbxiIJeWAnjeA954xOj9fnSvtDOG4rYukDuupnF
IlaCdGM1Ggte6M9SwkdQZPhYChyDXdLJioOV6bTc3Tc/8SqbqyJLrn8jYACmxHtN
qBTtbiaG4m6UeGUNiFVMhoManysGPRNY4lQ6tfY/I5T67edZELZUsjXNyco5jdOt
O9da7sL7jYhkA6h2HejzGV687Ux5/hzvNmej97vD6PJ3s/hfVEd3+UviE+OKlgrA
bSFArJakzRZQpk7UKpY+0a6+6kUY1WXNRHtKgn4ezsNoopgTKZn204+aotExDV5V
G6Fkq22iAEhvKdoFGAhaJ5TtITosGVGjx8Qc4Ct99zErLGf3cSV4mIwENpvsWTfi
+p9+f8TOIPWj91qrPdXVIuOGZ0PU1VPGN3MUhmg2/JCb5b+FZvOYijfM8OAy8wmT
UAqa/yu8E9O3FrS0Gn7MO4ySD343VfCIuWtpK0eIzGGPTq9CR/GeF+HYNUy+aNpg
PEYVaG1hJMNsn+Gb9xvOTopHf3Cuy1SSc5MveaSymT3zA6a32AZZsMnrc408qrRY
TLCEFRA6YyKbp/pSUCOs6+aAIgxBuu38r1lVKdeuoroHYSoZT/Z4ASXXkq6v368C
5Nc1sWhFO+Ev/jcgcDqEH5GR9M73S3HKVx8LG0goi8cv7/CFRjlAq5dp9kLv0pda
aJWnThKrFsn6j7D2ZJp+ECalLG4AYJgsi6jOK3uUFVzOvuhZbfFZvsU2ZKAHkfgt
ROQMs9t4cDbU3dLr1xbmbwQBShjqsj4i6uqg2wLDJXin++8FuT5nEigHDlp8bea3
f7KZNLxykRyb+OZrlbcziyNSnnZvi8hn5sGO6GlEKA9in8LkD8kHuFgpX7UNixCX
6o1q4Iaw6+GvCr+Gm1cYi8vSyPL79x2mNV6CqzWrvZrBYLAbr9GvGvsj9l+GPKBU
GQveaaOjdCDIHB8ioh5mA9O6fTbOm3WjLqTZn2eiUm67DJ9mll1f18Jd/zx1eTNU
htDWuaBEdKmdjFwWI/ESnK56bOPwGohOu7hZz38ndYFzdsmWd0p4AReBokfH/9p+
/4C0lusW4qa/WUQ6aFI4i3qMqrS3BmvUzfDQeXsGL36BorqB7OI6YwSTf8HSxM4p
561OJh5bufrFHm+Pv3d8fMmUyyeikiouiGpiW2G5T0/MF/LjIFJhtDdmr6gPh3uh
iMovKx7OIYh+Z3ojyWIe/Sex7B5iu/HOMqzcNtjRVFuRF82jWOB1ZsKHcJ/8dZe7
++m+uXC8DQT/rI1Kl00GvocnRFbEgX2T+ARmOymiBGCBC0UjDU/rLdTbLGuXbgyT
CTL4itwz+yESb6X4mlXiZiCLbC5n8rgqiYApI1hl8IvmYTYAcBGCFXUxHu8Jbo82
CpnO5qEZm4Jy6XivHeFSHmbeteuC9Q4m45e4YfwQ443g7TslKT9wJfJSU5qiLDFC
KPmf1flM+qrAuumaF7yBr4Zsw00qfmPG4hh54to596BfL6dVMtdPhlKuvLyKnlqG
sue21+TsKxiBNEEoP6FrFkMM3kXku77NNocWPXcSENMJ+tqRMRHfKQISu9ohkDtz
RSsu+ci3O8UH9mGJMY6UbfCXwbztpDT0qFqCXBSrTp6P/Ht8IDVDzcmRoKJXwi5N
UZA+oNliJGUqrKU0sc3noNRLqftnFtnC14pR7utee/K8Iedk8/vMlWrKeiqSxWnq
/NvXEJfrQQjJ6DrUc/4EHZuljY0hF5s3JIASJ+VbeEC+DJ0/M6xCtwPx/I+P9yIv
uQqGhTaN2165n0iu7FyeR+veatCJ3fLyKmcWq89WSZvpoucR2912UPPEwG+8brhf
CJRhmFfrCbvJEjjEnUZuMFx6lzberDUneVFitSepDgRS/j8wgByrhzIfRlQaAzAu
7kuwTu7yLzn9Kp+h4zk8x9wI4whuSK4A6AzwWoSFfw+KNprH7chAeCrZ4mvKHAVE
8aqBfrbSJ1ZYx52oMHExs3xKm7zoHFYn1iZyjnNQXLSCQV+FVTyMDmoWE9u01kNU
AxiPR28vEVuqmv58O5N1F7V0zMmkMstIyWbKponsG/jmPGS8xll5cerahJEHK1wa
xlZoolZSWDe3FPfNfR2NkjSc2PZdpLv1aTMYzv+OCAhDDZsHu8emOozxz1E4C7sW
GSpKjWrxOFqSgO2Un1DufwotBo+b9aKeej2qGJgxEeyyOvI9zl9hjZYmbHmO74rD
85MDLjjGMQCKI+lb1iMz2MdYFXhS3n9/Pmgey26AH7lW1F8WTXdTRfhnVd2R2nQ7
Qk8+Ocujx4V/gENDgHQ6a7TFrAXwr1EOqzGg+yLOKdm6FOA6KsVDkF+0b8vVEG2z
UdT3ypqJftHrwp8RUQHAOam0Biw7iAcL4ZXg7EIWMJQcdNOo+j1YhxaeNFo1chT2
ouwi467ZpzbwSUDGcvjrjDD36dIf1blNti37LLBCn5jHH1SYE7ng48g4neUXDO/L
SWOq2eo2M8B7bUeA7j3DRp6IOT6Mu0xCyKjPtGDbeSicZV1Szuu56JJ7c4/eJFjY
sod7UCE4syrmW+3PyEXDcfM56zolLM8VeGwJWR1BXifIgOZ4dmcfuee5xOCrClYb
KSXuAbItR8fz+R5BFh8qTVQ4ZmSIgQYdy/CvOo+yvg7Vk+pYwgwOm9O+k5JfJqcq
TPhHf24elO/5ZEXBi+52yEWkrLYGa4HBKwyQx0GimybB5zxjnDKc8dzibEFTO5zl
0gnfoH5WngfO24uKkvUacOUZQN6Xd/EesH/GbRGCz/iEqmB55zf1+GT7onYcWy/r
5CJCjXrq0eXAYUpXWI4mIk5GVA6RKZPoqw6M3zGUOR91GtQX8HrzkIUBQ7QD3Lp/
yhTd1Nc1bc1yLiHilqhIIogDsPcRz9p8NRU8PZHTFdSofIyE+oSzMn2HScaAOsOf
Vv0IO61t8ggE0XTtRnXFN6zroa7fi7JoHCiH9tQ1pXvt3QYp+WWqdmyjftvaZztD
Dibgftjl+5MyjiiohHWhn1gR0LW5/xuGNCtU/LT6T/7qfPdsBPrTfVxvO4wVho9F
oje/MpZ6693mX4n1+iyzKrurp2qOxIAsJj+Z0CW8n+gskM7me3qXFew/ABdiZJ2n
MOlYhPVecq9NBWPX7jH7QuUTh7RVLaa2PQs39r1IoVJyrRGsBY5JCr7R7OfSsZ70
46r54sS3Gavl4WOKnCTiHPf8CqcHELlvtC88LGxkHwHgmqkU8si1Oqfjdkuq47uO
hS+AAZxavc2zoVkh/iXhi7djIlEIHovJq8rey3K5eeXgP2dKmgGDaskQBf8pDmmr
LSIM1myBafI+8GBJRS3RD+XgExLOb5YGTpHFY3bn/Mn/jl/IiI5suYIuqGvU5frR
rRAP9ILH6n0HMy2fWm0uOs41Igl8MPHzZjdmtGkvPYkbNHSoc+h7WZrLGxIaZmeP
7j/Efdbd61R31rMAgNDMfUZKUaPbOxbUPAfr3OJ8Hm4GaJM7rfnlvsctahaTYfvi
9wDPZQSigiD+LAOV6ObqLkLhd78MSWbDFZ0NA39b5SuWICxfthWFTT1MazVoIg/b
EncU9+wlFhq/OBq5fDzHCJsRz1A8iuypmN/iW7DPtW7xfHFyNlNV+XahStDzQDW2
HrCtuxCB2SE3U5i/A1LZrhNUpdj90i3MsvJ9sE3kNgJkbA7kGaoapDsjMq/c9UWO
s7RD33Zx9EdtyFu91QapnXCsu624zPXK7cJ4+AzaMEb7elbnWA2An58G/0H8ck27
ibkaTGQBql867wZ/nXZsCq+8lbYn+24fFlVIeU82WtmQraN7SZ5sJBoaJ3jR4k9q
UA/uhDmtW2ICNzHoyjzmlkJFpdaexdxp3NrSDaI2Ech34ezpRUfMViTVvh7yb2MI
JD6AgV/aqExAmjmzAINcBD2VWHXmdNZ40qdaVHRGB9lgUU6bahmY00dJaIMlp0dR
HyXT4MI4yU5W2INwmYj62M2ftD0WYpjZUreZk4D9PWe2jWqlF7orJHbjI+xtMo75
F2Q4VgaBNSZllmupeDWt7pi+HsFJq/BLMzv8Pis1zUKtMV4XN4uF7tGGGsXbCynf
pkz0JpQn5nx+isjKWYTkHww9YmYZEPeZOYq6xTZTlKCpdRDbop5kDNCfB2VDbevX
vPD/80ESHv4WvBZr9NS1ZPzsqRwXioQbiS/BOELBA1e649TASgx6Ec4zgjAkp/Pv
SPC9doeA59hcpzE5GcGLBF8B5NbPPzmLq9sJAD2yn4BHPrpqas+dN1KqWSGCwvwn
eVyMmsgQLBrPv3573CGNxXtQ0NuX3s6gxdHKG7lyKRsnIFyhKQ9TtzVlzPVqauU/
oxIV7c6ES4W76A1GHDAnGv3CZpgAWIOz7xxPLEIV5OQ8tvXsSqpRitidK7hp1lc1
+xgJI3DnCO1YeFKM+MBV+IziUNDPgRAgmq/rT5ALcBy93q4PxHCJfjno0EhabUNl
eqNkZlIFys8VIPN0SFRewm4JuFOS6AosRyRqMNF4dl23xhBXXzCuteBrG9J9fw7y
DEJB9M5toDVOAaDv+0dT4fL/vWeaoHk+MFENvNGPfNTTCUsrPhRMKEZ9HRAWo4H8
wBCrBm1GMj5jO+mw045WuHRA2oBVCNG9jkslnwkLHDkRn4hbgWcBTo3Q5Q1u9agr
uUAv9VcihbO5aeBT7eiZe4jGEv3Wj0XE2/D7glAg+s3irjSLykEcjH9/9QgN+i9B
KVtwACm5O7k/xae+r6Axtek5PGB7Su3VWSLOp+LnhuV6sIAVk9Ig/azs38QSq570
QnibbS1/wCQqHm+tQspR/oJhw0KhA0MQ42c34o1AIkfwt+v4B5lKVno51LNEdSLz
gfp+nFWmksuyUqVQZdmlYRNXhTJ/LiPOeXX11GKxZuMoUs5xDKAF1rrB3imnap2T
RBAheBdKA/TFtRg0dLz6gZI4413unz99Rtr1VI+pKgyP/M2vMz0mDy5ThVNgbxig
jtYCoanvx3iJ/iWqiOGnJNo95O9amasAwKU7Hg6C2tHo8X3xOV3EjVhTrHQNs5mK
471an1HFjnxIh4thj4MaBqxnO9RZKhwuvoHXYtJXUpLDHqKh17PGaXvkAtMp1q7i
E/FD2AlyLXSZDacABkXQVGA/7FLIicddFcS6mpa3Oyfjk6nJ01AHooCR1m6tyTCF
z/M+JkMhxfbv2xrA09jggfdDREbUnNZBWd7lClj6n5EJWzwZfNuzq/L0e4EegchA
XJfqw0EjaFwCSoIE0sPjLLGxPBpBq5uybkuVn9h6//HjmW6Udysg49WMEIuSIzUk
pRd7cQ8uvLBgHbQrpqaBHVaB8qAazxO4k4zuWCzWQTXhOJU0oiyHoIe7YJo8QbfJ
skzJQyd1Z4do8oae2ZE33wv2hI9T4N0YOcn81yPCr6lctTqtvwJCgS2A6V1xCeG8
PzJ9wt3L2eq//Y7ZzgWDPmksUWjE0os0Cd7SBGuTk1Zko+c1Q6RkQPnxIP1YKCIe
EXeYDLTZYrQNp0hhd13me4dPFXqrK5K2YBaIpwXPbVQOrlWiahdXkBNYxuibiRrU
UGm2ktFuEJGNLEyTzILHA+4UVwa0sJLHbW9yTYrf1gXk+8Q9eV6bypQ4LrbaBBxA
lJSxsssVG8CCQbgjSaCW+OAqcX+1vZjtCxo7NYvSvRr5yekutgCxazmptd9Ev55V
vVMgRzSGNdp7pMKxIa8h9s3/rQ01smHKpN40uIz2YT4RaGBS7aFMKYYhQG1myFxR
paHMs8wSPQNXSf6MWj5EcSpniflfxVjnaAj01jW/GSRzIgzoqMgcO0zQZPof+6+Z
JSvpt/8lBk2ICgyqvPiPspc3+qvDepsRJOo4gMq0xqWU65f1EubWiTeFrYb2ZS7+
wfl9iqPvX1XclwaujEZsu2ueVCmjHIgUzPIOHR8Z7/mKqbL/sxWIdgtv8d/ZTWeJ
+ArMPa7SC4z2bPGgNlhlzRD2MU/wtSZotKx3Q0bvrCdxmhhNCP5hN/LDplaJW0pR
3j/2X/q5Jh03EHgKaA0P3UZ/CN7vUump2Cbf83KunDzus/bsF+IyYrxVD5IFb2Xh
y3o9rC2i7cVCQzPB3DQ9EjC041JTtBgIdB728DF6CoyRbijY96hYpHpmssXZ7iU7
u+SLq2dVp6ek83EGVAJWe6tUOLB2LaQCNFT6W1/HrOtidrIOgZudaJApWD5ExWZA
HFEEMMPhsYyjv+5ixnsNUEaEB/y7+8Sw+BK9aQiGIsAO9uSEbHWlmWOaDeKPpFeT
rKVpoen3IGJhIqAvzCu9jvro1B8dxQ8litTV+mRSWCN/T+3Z61t9kPQ4miILrSqO
/6Oi+RfKViUFcH4QafAoJ563jB6BiDSGttPz09fR4/6cXPsHuD+fU24I02HYAnJe
aCcborJaJl667jYCqlEDC4WAIxx911UZKEumLj7W/8mfQchA1q/9fO/gyy+KIxCj
DWjZUNj+pDJm25245FlaCqD8qHI7h4D+2zsN9TRLvmVoMmTfp4WPl63y1aV/Cuzv
fk4Q9I6MBqKSz1XhysEBDVD2EfYZFIfG/qcvM9OyEz3lGcOgXzWTLlCNQHDjdSeF
r+1r6QnR4LbSQM3UlbzsuFzYtSYu+FCtdUx1H3AZY3+AdrAU3Yzw4mY5UOcoP6ZF
eMVDe7McrFRmzA4CtS2dit7nsDO2hIRG6L170ekrQLt6yprRXnZmuoAZcOlJcxvs
hYxs3pe4DMtvmr817f0M3mg3lMaMxFKeaMA2p2zVmiQ2W5X6wfY+aTOqrnNOXMiT
WdLATYAv1BsVKwr7r7dYQO3UyjkS4Hub4016JIWuRirTDry9qecaqp2fd/H/K1zP
J80PAyptsYgsvKvg7tjHe3bjUXENkAdhlgYUgenop5A9P3OBUJ1irJuzizC/bWtU
hQOykKPBSCd36S+IPGWmYXUmujoPXgh7S9+EKRMyqOzoMdvpfJoqAKKDSF2cVsdz
EBj3/DlPZTyqElUJQlRyC9PQS0hqyyNe8lYrBjzE/63e8YsiLLuPbHxwEENttKPR
1oL961pm2nB/daB0f1aBtWRUwn6TEl1wgDU0levIj7wpv83UAriw+GVyRVkkuCHf
qvVqhsYpqWAxycRiVlDvjriIyHjvDHoc/7i5/+mwsa1m6vKq8hI4+8i01q3acPjF
BycEppW6euQ83Rp3p7EtsIYi9vi90aldJY3PRl/XV2ss0cXRzOYE7srATf8iw0r3
ON3zaVAa9sXoAWdFcD6lF9C5tOhr/0LiDcSsLlyj71YkyMg8fRTDF5xOzgFOZZLD
LmsVA1jAHt7zheFUBbsze3uo3azXvCbNpJqZdmDzNLm6ZpZH3/57Nu60cbNq1PdL
xC7IRIUtTmCfWOH/lFKO/ryPcP+vNit4LkXK0btulHxBIkGNa5FmFMfXULt/z9gO
3XSXNoUReqbPlul5PIYuqybbciK9SKOCuYEjLKfTKh1jfcEXfdKUCitaMFHwOnDo
RkDSj2iV4gjo2ta3i9RZpVblhAaM59mFSUgilqxgl9irrg96NFu/7LK2yD/3fJsq
rw3ZOc2NqG3gAttB/Uihiic5YDIK5131i4ts5od6hoQZQZyHjS9DNIrVinTzPL/L
AMoD0uSnqUnMleDL7IOduCpxo4uSBlmGE35bXK3+fuqNaFOOhnx4zu7rYeOoPtKg
L6my3ouLVrP2O8GH2cAoSG9zmCFUidPJPacSHhJxD+WHP4iKNE5dctjxFJgChiAO
jHpVHuMdEMWle7NByX1VyXj13I2hVNP5bIdfzBu62jpx5Xt0m24anub7Q9aJI0Gv
yadlTUVmUZBnbJCiGYsz9MYpTlVOJnVgSglUsYTrtjWafHyhFMEni02oO+KvIbpR
ULJzE/ZjR7Znat1GEqkI3njpRuamabQKRZgTJs5KKZQhOidI/ZEwBighxi1nzRoU
KviifoHSxvvWAL2PB5CVr95+4QV8xgP/yiqclCShDADNiRJbHjen+s6PilP/B7Wl
QcLx0lfxAVWimLaiysljaX62pPImCz+OvawOlj1vROICFpry06NGYqeaB8WWzbfL
ItqCUE3ai2enKyixoHeGbORxrHMthMAL9tXl7gZWgXOhRgCM8xuY7qj+ZpMtijd6
ZcxmFYKcZA+eO/PpUm5Labr9HCncMtq/MFOKyWDC4BgvnNCApMUWqThpqJa+Knqb
BDP3Msmc5oCsmV65NOTgJJJqNfp7JSBsMbckjKlyVj1hOZ8spZUCV1AmytDwmZjl
Tq0xXMEg/iLZ2ykpqZrL+j5BSO5CFdktalwsLF/IhL7sFWnBx0Ms4J+7R5te/Yck
VW7njnWV5dXwU4PqEcvQQ26HpgGVo25ioGxRVy510rzRNXlwAPNMXnbYTYe5kntZ
ePsJ/ZcV3XTnDiKyYpGVKnkhXjxAXMV6JuMakaCUFAtOSixUWPJqmZc1inzUePFs
fgBr3w+7evNDQT8rCyIpsZHhUxKL+KmP54uc2p8hmEZ2NWvJnZP3ESZyZ6KdzHdU
TP0Bgpn5YicfiGdULyPRV4Ho1/dkcXNlmXjlSawsYZVTtxxyXvLmevXiIsHk+VDB
rlIw3J0ttABZuo7KjbJLhQXUGHWuxBDX+LpPcPDGk5hYSLZcpIbdThwkGLm54Att
l4PU5WT6sYDr5VdvR8J5OMiq5/1yan3DPKCLffnh6gGFatm62w18cuRxPIGyS4yd
mVE/y524sKjwywNkmi/MQ/paGkULKmYEJe8bWiObqxDBjhSOws85/OaBY0Ef88i6
decL6Mj3B5XxBXsiXqTfkrjaUh0Ibuf/5Qgp0AL6EMkavDmrsAwpDqLaB6nM+N7V
2D9qtJzRPmsfOSeA1Jn77CVFeYJUFn4u9bCw24VExUNFNVyb8egADlZCHrG6j1+6
LAxc86drJTEBZGXeJqzTTcLjR7fpx/Jq9Tl9vraxE5w9nocrTyDqk0Z971axErys
0ktLqdsLhTqZsSFbcDfOrIQEanQyjCgvNERNDA5E3rZBHEEnvlj9Vh2n0XSPcUh+
wPgPfivP1aOkZB/e7iNxY2HAD/kNXhfk5f+RKYLm3x5Asjv4GTefg8f52ojnfRUI
3w1MBwCg4N6ICSBdJO4tnWTtrJbodg/ofgD6cwjLjpJI6wr+MepHyOcrR4oKo5t6
OtAw43wOqr7hD3/E4YethRjttdLXEAc9Ggt5HgxGhLyQ/sVQOchWENU2OtszLGTM
SBBnGWTtRIHmsoKk8blIBbTwQbYB2cIKUQLiUTzdGTHBKArQw1OEprmOSs67AMMO
grme+BoqXJ29aFSz1zJKOfMArbxh2AO6wsd4Y8lScS7RjIChMZTHv9hqfQcYPIqj
ygsqPBpBTf0FSkYX+JCQuL3jkceZALLrewYQ4XDwK2i22gmwkHeiAK3hr1mHlmqm
sFFLYPyNx/9k8tDc9Qp746zLKxBzwrwiMMOtGH7M3BajdpdEmi/5hvQ3ZJZPUbSi
zkBbn+X78sJcdWTkm3XEN7/7UnvXL26m0VZiBkykPB5VZ/8ma8A4qvz3/uEDvKyv
V0qBghP/kwaEY8ZtiavuHUFMcQGGrfmBMEWM382Xl8ZrXnvC2/oiajKJlm8JNjsW
PuIEoClVKzTSqCWLp1tPzfmJXHd5J8uYnc3V8cuCRk7KhtFylnRkR9YJ89Epi75b
FXzlYiiHNi5Zt1bMAON3SR7tFHuo2CyaWIW1TIta+LDqybaZ2vCkbi2W+E5JSDdp
eZaBaWd4jolkQjCl7kwd2KrfSosWXZukL/yCu95Q81DuN71LdHqCz3br8nX99vZ2
tvpvF1Ksqu1EIBxlB2XrNr0vrG3eXX4Rb26CMumYQIW3lidw4QbkVGZnzdtDmVBh
exTCaxCyTaBx93f+L7+SPZMJhRBfvDo6xpG8b6h6lq30U25+YkzTh+kThUbRhLSu
0tugjC4EtNo6CaPaul2JP8W1IUHWpve32qCM0oGtiCt6IZcCBaH52OMWFhlIha8Q
gTbKVBvYFTcsu/3l+XMSuZC69L31oD4XWXPHJDsJgMrcA0Vo0hgaje7n2aNVLU44
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ju4DAtGPGVmzaPlp+JZ73zGYF6EnOo/TIgAcByu8S/mxwtMrXdEPDXaw6Z8+LRmg
ivv0uIOf+mePqIv/rGLdOW2QdTNnw3RRgs0oXFc4iD9kKEFHbzciCtfWeKlXQYdO
nMj3PFgShXdmH8NeQ8H5msQ5hbIeIKhTiekW2agqdXpE5dUpboamO+ahY1aPETNh
2lN9PUIguCP0u2PAsTs1o0jj+2lpIXKfsXQHHj9ci07o345DA8FSTw1kSEdsQFtt
YoiBeySfkF2JxwVySqpUH5y4MNHrKUEJICY+eXcLQ+iiRB/1tp+++qe4y1c713nH
jl5DcNNpOQ7F4FVqIk0NPg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 21648 )
`pragma protect data_block
HKpLdTuBzC89qL1mcineIOv28hjdHuWjUJzHVKQssogF4ix0B/nTic+YaklzT34F
jZEqRnHtJtabcn9cyalOsEYPt8F5J+C5lHElRCAcMNYcCbW+x4xbMDsnsCI60eEt
E1yPVCdEklXQxvoy4UCwqhXOCztqW5rR8j6bTIjLRgPJBlARPseL/4feUgw9nnvQ
p3hBHk6MKOqkpsM9npWT/7U7Nt4OZ+JrYoTuRnk0iyQpU5+xr7a7tMSQKRhXoxUz
z4vtktnkHk38hrT5K97IByhvd9LxGhb+bOfiqFk6lWuZoYqueBt+yk8bHIyo2qN1
J3SnU9ZEBWTCVqjU/GYWB9TDSHuPX7TKRfoW6TN+kPJj7dBWIYX/7VsCf0JIaXAw
43xL77ZVNPaPNW/qDqgnxTrOXKT+5KGnXqaO8WbJDvKuTAh+jV+uRzIeigj3RYKH
DB+hMa8LXQ5vrcFqEe8i+DGm5XOJO8PvjYKt+sLffZ6tc9Q6Uw/spSAnaArp89ju
Mwg41JfErZ8JSJdpZCyWFp1XqxjApuqU3ON3iiTCna1QIHsmGnkXqhyQdI2Mmjbx
5PXnRXtM7OfhSiHcSt7GRrZ8ah3COcMc2SGzCLQgXArjldnXTnFEPxFuxsAVrZWN
i2DT9uKAjPzDyUTjxqKjrgOPLcQ4sGv+I4nIuEVJmjpCSnoG8fRB+C15ndFX2kml
ePr1qDSUTT8xyVQCz3w2q8O5yEkWxkwrcuUYZicSr/wRKLkScN0Ciw9KgI04z/5e
OSFKJK6WaepPERKcIt4L8dh5Opho2yPUVpEtSeUQR0qkLi4TPQQA4V7NkUKp928b
Tpcaj7AEbdYkIpT0rUCY+PDBmDpSVIaAo6StxZ7vgC23VVXnp8H1JwqErNKFwPUI
eGRgfvNPwTPShBXDz55f8ucPGTBm9pGqSeV2GJg9qvS2O8HR84SQagbVPqH1B0V9
sADqIN16rm/u36ws6MrR4VlHCChXe81S7eZRnPqGmBgvAIFODm4eX8HbT6YJuF0h
1VOVxn+OM/VT2h8473hVIpwwep88xNdajWuJfDE0gGA0eWWp4R0hs26k28Vo5pR8
ZTf29UKmBahLZXRtxTgDHaLkEPnFZTH8spyoR9Ccs+h8g8gcR6o+/alwnGknxn1w
lmZxje7t3WuaA1I7ifd9aBKtXuAaFhyj33oWCAKxkYlmTNT2FfP34ofYi0RokKsf
TINHlQ1xHVZQsOv4eG9PP9U47lp+Ck7PHWarKuTkNgNN1MUjHBiQtBl67XlbzY6W
o7Yk37x7aFmhiUr+0mOxz5RM0qrSK0IQsYlnRGrsXH8L3M9lcl0BNTJQuM5U4wLU
2HdueVZNNq9WwszsaLVLBTbWG91lze+OL4Nfa6DAqKRTK5H5fJ6MhGlk/VkfB93Z
BKeL1NKUS0lu1BoDnNaJ8KYxYLdYeBT2jkQCMdns4doy27u5t/FAXAwJlMbWDYw2
ssXmIyUJoia0gvFZdpU9uPWi9yMPrTfyh4+ownSs/83hSyKSK64ihKQABC7g14uQ
f3hbB3ru+paQ8jjfG0ZTc7YQJl3M3OzZigMwXOqXO92CIIEp09ieTWhOOjK8o7kF
NXwonD8+U9Pdk08L6PkEEF3gYSY/cL/uKrzepWFBmbh/xF1JI799h5nSEGhn7USM
1ZamfBgKLb+P1YfKTLlGnqnzOX7VLBYx+jJ/aIqQ9ehokxTJ15cZuBHHWi7qRM3P
WMW2/kcRS721plAsxJWrzBqbKhp+VKI8aS8k+jMAMja7j5qie6bjFp6m1esTibAq
QdHTm8ezC8MyUlPP+7AFL6ZKlJtATRIn85LF7dXoSnmafXWulLwoK4ZMRxQvYBLX
d0B00MD23snOuQ1ch/d7FXX3OC5BXZzvzld6KuFfMeUPApW9FqVaoH7hT84eyZTA
Esn6DTN7PNJq9PSj6WWxDt1LAUUb0AWund33n61jUQ1lvbhfUQB6bp9OiEk+u/L0
H+uaQXSUwdVe52nYfG+sjmWU+GSlqqff/kv34pJF56fWTo05j0ZrnGI0JBSM9TZg
5GBWpEcFzpBpQBWg5zwvXdpZc+awrlrKPdrzf+5B1NFK9nVulDt963DuQrmQSLtb
bze6xD7hU3rosLFtUqcVKynkoepZPjJnmE5Gz8fmvd0dQ1dxOAKRB18mzH6a/pod
5TJa5pP4iJLayCkbO0zA8T8HsNQ2QAh2LkUZmfELIULQSgX5XZ/Byx3a2kgRtB55
ns+CCdYMwLs3AdN46LDse3nFoXIPFhBy5HZaR1gErn4bkKQfkMGB+opjCgV/nEbK
7l4gRK1lM6i/usxvtngrAtVfkASwdCDYqZ2TYjwBFgiyUYhSXqYYfeuGdKjYq5R9
0PlnYv6EVvKe2cSJPmZMWXjKsUadUr+PJYYgkcRtlLTzNNhTlIRR3BwwYlSnIGKI
J7wvnFxpZQ/OWyY9oVwAOs0WzMJHGQpvkwd4vG4nbjdmXZMMOW8XamggVAKPP5qO
x8HqtAhbUkPNR3yVfc/HKkV4rvdk9gjdn6ojHUwkT2he/dfDo9kjqMtIdiszXVZs
g2keEoJLIspikSfqXodcWvIXnAuLlVSPy/no4ObjF/JuB3JsMSOWgK/mnpJhEQBx
Qoz/XwKEuv7kcyL7M+E/FnkYFTWDjGtnCZZ6HNt0BJRAksCKLE4cUGCliHXXXJT+
9wqFh2VCSjxmYFMuSOoBqVb0CLtxpOM3GgpfTo1tVfT4WMklEF0AgLN0Kbx7z0tB
tu+ne3HrDlmNKfdf1NnrcmQEwQvSR57mpK6CH6uul7pjIn4qvA3eCdIBymVei9Ye
tvLL7t5kNF//LxEkOvOEN1iFmjzIhnySULBbcmKlTUNDZwbGg3HAEyactMG4nMiO
VSLZgnyIe8Vm68e5t0sQPSpmQSw2NuSfm6noTlNj3ZJhUB0fS+wQIvM/7q/L00c4
RabQ54grU5vQXA/RIJCVAxQkFoI7Yd+WA/VcZ7DZ+cE+aD8tH3UB2UhCFG+yVRKD
9BaSbZhHOGcwkI1DJJSr8oFMRXLR2F2xUb7UQXmAMQy1k2uCV1MPqU3NOGp+ZcHM
3bHa/Nzag1uhkKVl65vBmibnRcnZkcqEsDa3oJH1IgjnMsnTOMqpmelRuYsz8c8+
TgSDxX9GOHPi2ww1xrQfUPrdoqwv1JSimtu2gLBsvUImfa3Tt6DBuEXeXMC/I1kC
1jYGXV8eHq4dFiTgvmjwxnS9wq0y4hc3NlFadpKjrVagi74ON1K2LFwSz+OXLDKJ
c7IF5AhtLIJShcXLE3Vvl+T2R7JiilPwcn/6eBjVC+d1tGZZULdWMi2GIzmfeNt1
Z4UpvMyUq33hXUljmNq1o4mdJ3v7Opoi43zxEAn+jZ/9oJvb0gZ7cjMlEayNN90j
AOJuFfPEFxyWD6neMQst5O2mefq7UTinICk0jy6aLUgsBzE3QXsUwEj07yd+jl00
tJZ3RzNaCoKkdz8Lv2oZWLB3/f0A/zcEtlxptCGej4vL8GLWvvms/rXAWsbmhS2v
PFpqA6nTXQZHB5ZRX5VNvrapL2nQLqcZQu43hVwMWsjDKvGeHau70q0yRypZa0/v
xLKgTakmbJnMoJ9O/5lxCKxA9QY8Zww9gSeQSwIL63ATXwzZVgFyVXaFYCd0AFbM
8uQeFgqVHHJ78+hJv1hWY9PBpgizBSzUa9XncvskOG3Lbvw4x6gJmd07qYcfYW9v
e08alKKuMSC4YamxZviaTuAO7PRM6BrNtEQKHxE3k9PDTktpJ+3Owm9+VtOeTl5y
R26T3Vfh/2+dUc5d3mdDF8lqMJuwDRpc5ty3yXdT2TYG3qDN9rAMVii+infu96pL
0D2A7+n560wUFHW94HFsnKcjRWxQVW3sdZb7YqNsHXcMggE8xiP3LrW/vFQwutBB
mIXDLsaVRyC2RgT3WZSeDtvdUdl7QTuwH0yKsxEN01b5CKmTGTh0GENDNdRjvKfR
IBi94/IFvwbtwnBxSpXGxHcytEQTIOXb6c/LdvIW1yxPlIQbSjsE6VXNlH6hrw5r
gMZICOQdQW60eDSCeVBotoYiLEgrQwZ8WLpAQyaYkScbgSA1qMpPC/9NyhJbD6oM
e7cAcalDCk0WSpbarfOAWU1eOOvl9ZWjpIvCKU6HAjH3Kid4pH0fZ8Ihxoz5StEi
c7vzq5wFnAZrI+1SkRPIS2hN5nrUwavyPfw3Db+L9ZhyZF7xulyaf5dAM2pZ6J+X
BD4vrjAq+IfFwskLdwWUly1jt4PM7ZyD/EPAYFa0r7DhI5icM29fp8jWxeJDaVDE
luLBq3TE062nQEaXN6CU7sADox4vGu6jDaXDqMDMr8HGErlbbtEUk+KLJVwi8U6w
91ngmx98bQZ7MQRN2ffg+lIunGThPQNSy+gIlxgQdHvo2Re0/PymL4F+bOM2uO1K
/QadT2Tfcp4paYK9Ewu7xrDXa9vNSDCVVDZFAbVHNHHt1YTZ6TABTrjASbO4mxUR
84mGq8bvAWampqu4Z+3qtXWakhP/vRV247Gwzk4Fna5JMl3YEN6STIUAMGdnrhlr
Mrk0cDxGpn6sol3jS1UPFQRoQvjQpTGHP1r6/yYh58eB/r24qrq+Drd3vicI7gg5
1S3qDl9AtrsFex283XWGU1mmhLISoeItef6E7SI0LXXyPNJWXcuYMmAjXpNY97MG
aVX8KTnpH7otiB8IJbZk09euGtZYQZ9TcpHiwcXkjAP2RZB3zf/fvS7kMivdvkr4
jfXgBLZDLeGgDSP263DFPzKG8ze5yhyviElhVBCGJfJRLLMLSzj2so8Y+DED2i0D
aq39mdweZUDNc4PxLaf+AZjwLO8dXkTeDLVT5zMGWMxIAwuV7oFz8RwovF1qFaDP
z6oCInPyLttELQcIxEKO/Zt4Dw7SKWrtr01w4akihUjSYfoxhz89NQDSxF6M8B3t
nglH9F6QSk4IhZaj77lGyxXoBgaJK+h0j+Q9f1fmMV4vd3HlkIFaxKgkBXmsrqvL
rir5klRChtcKfL33FPFDHZymFLlZY5YTog2Hvo7kWG4kC3PinKJ3cfKTGVFMISXr
p29872KirY0z3fVJQKB9/c9ZjQfDAcxhShfRhzq9g8pJiP5CxarzeCGGpPC7uVld
nU704WqQNNVpsHRrhToMWd0kOjXzMZXzV3yWg6/IbzdR5J+ADoiPOeWccGeRXsTQ
utsyko6QiSMGBq0McJLO97kqFa0Yg4n5jLfFwYFYj1CVD40JtFTEsxLE5Xhnly9m
j50ioEzs2xJyX8fnxUmzcooYGCd1WEq6soS6rz5p+HCNr9cZZCe07YamNb6kOx4Z
kxd9GqsTeNx/7D58CITuU54hzEnqGjnlhiiQbvwmEGSCI380KWLiinwvDGyS4dbU
bxMlLQhHszLmfb+vny+WJSDAwS1jJ8IRtAu4MVyew19mo4xjmLMjGMr4vOhGQ29y
nkLdOfpTKB9izMZte3m7vdl5RyGrYS/ZBkugERUjPZ24uP72TT97Z2o1ooeAYNKg
BRct2GfGmipvek3QMp0YmKeMvbZXC7aweE4wLHeEb3eBVtJPOS4edycMiZYHljQU
r8W6npDKnAvGIwgxq082v2lqG9gfH0TrlgdLVuCVNi65CFYKqYU8y8mrHUsVYCeb
yCqwKTvAGS9XmkurMW437pjET3m4k30QuV4OaEWcq77461vnE6RwzBSxD7eUm+U7
poLIJku21a1sv4pOukFBUv/ftofV0YhfYKvzFlqxSIdzqBpk2SUMCRaf6jLLW0E2
cdIaBCOvzE9jr2b8wkh/+oWlDsvYECpMvjpMb+megCBXLAFEVSbNfWSNhfaunOnX
Hf2s+fNyFIpqHa9Sh5LvesEfvAmKFJe6clzrZmY/qACZNoZckAH/j/FfmKLfilct
ay7ukAhNi0qDOer8/o4gzbyftv7lcXscfzLs4+i7v6V+PZKS+iF95sYcXQGzYTjE
axNRLFEiS81f50RWctaqY1GqigQI+w51USHpWh1yIVNwPd0bHWuxPU/x+xZNi5IQ
W5myTqytehJo4OJ3FMpHF0hFe7CffIyh2DiBpzDtgkQdOHseujdJTQ3tAQKu5h4p
Adl+Xyep4Gkl7cdWEx0fEJ0781j25iLrYpLWFPv0EFzJ59ZpykRK3GwU8bt+d5Qw
tygXYwEibZ+NDCWilNkWoT8hX8PD2kfenoLM0kBFuLegHDvcPb2BXF0cdqGNtuvc
BZWn7t21ZFVA9Etsb76CTTbxZ4MidgRW84wnQmE5ybu7duWISZuwymyhV1ERyrhx
QJsoQ+p5xDDuJG9KrJ93l/TacXNt260r4erqhyCXdYoL2fLPuwH3kTdjbNsLJANY
NZNsOwdhqFkzYuvFtiP6SVuUnzzS8IImdRwHrU2rm/FTPoRuPNsp4uYTXuo/VX/X
MRFOuzZGqSAMOMjJPEwKnpBsgYsV7kIveUDMau7b+xj7ahyC9fJOlxNVfFuHEgbf
SoB/RyN3x745fhClVik4i0VKSKy2UEtHe8MpOpbz5/uipGYzGXA5N5jVCVonfJuQ
NpG/D4KPbc1ZAn2ktA4sAnQ57ygE8FRklWztJV2ETrbVCdAms9tQ48cweBVNr29h
iSulv36EU//hjYQsPFiBYc9XFsVVXF56t8gviY5J3t6saSNT+fVhQHhWKR0XiHTc
+6Rlgodma6j7xV4iShj86dWqQyF6XI25CgSseV85CzvTTrFaTq45i9ZTZdVxeNnA
OW99PRireonUTLk6bqKUHNf65bNZTii0nlDPZYJAOFeQyZu2WLPddCIuaYVHjsq5
wfTp3KQJXWaLU03Ufpe+SiWfAKwpt1sy9wU1bB4R31EsilWlP4uQjFp/fulnYgyj
aEm3Kt4gU8Xsbh5li3PzB/kaPGI4cAXEfZOVOZSyUMsrhBmoLY6ozGbZ+Zg+2jsC
AOwdLFAyxKp3RVkPvwLp1PRlRQph0pTwgmuEpH86ooCwoKclAnPw4pp2mKrG+FWF
j1Ft1/9agvSawaEY1s+261+WtnZi34y3h3N174ihuSyMbvxeFS4NVDG+I6FdJFTc
NrsSZ3JcEm2PH5WUn5cfShp3LXZpW76JKO6dHXI90xrsLlUOqfWbEsSkTrhdhMqy
YpzPFXQYa3hqP67fLDIwmEe4D3hyLUuNbJbFDsS1FEbA+bUluSVWmayIYeAcUG1B
Nh2iIt4KJUZSCr0RgDdCsPfFJZS7p98yVpgyXYAsBm5mlkaYtS0ZsVXRlJ3iwPrd
7MQsgEBvlXxlj1A1dafsz/D/9S5CvY+TZp+oBRX5Y3GuYdfY4S15Vu7XDUY9nbac
h4BkTzHQddxZ2w3NWLO946QNcPksxBugMKTSTkHFkvxuO0gN6HgmGinzteUtu3DK
ilQdeK1KsRavDdzFQEBZzkFRnqzsN1WhnlMqSA4u9n1XIQF+iFOy2r+rdVd2uqii
FYluPwYEmwXAWyvXO4SrsGEOSl/RKm8ENU83hHohVfIKclrs/9pJ1oWFIm3tkpgV
47FW8nCa7u1B8BJX2jv144lM7VPtxH/W4e19csmQvyB4f0vSdrk/Yz9LZnmAbD7b
4leFEMDDdlZ3+CABHY+wK0nWyJtLoZrrP4AejC7DLDjOXwcEhv21hni3pr+Jpil4
OLIz009GOA3iCBttC4+n5kNAXGHNR0gQGQpvRTAlLjBc+OyH+jy82iTWN4QON3qQ
Xg3DLZecKCIk5x8/2RjTq4WItq+sRMCTtatSQ0UUn52lYTj0qSRqLJwfnDdbRnVF
F6JnK6H51FqBmD/hyaZJ8Jg2BW6DVQ31wRzrRk1lqzM8pB8xN7K22k60T1XP+u7B
c274XQwDrVV4Mlbxd2cR6Fd08tNjgraoDcRDcf0DRRVfuBJrMqYauTPiKtLCMPF7
fJ+xGRlBIFNUlhmS7TaE2cnac4OYtebkG2u2uaDjRCjdbovCqLQdm+r4+JSfeIQR
QTKJL+fA2AEWmDA169pm14G5KF95ibpYpSO2xpbvgElxEoAKpvydf0oUCHAF59Q6
4Kd/A/vvrOwvR2qq61i6CaOAcY1WkB0gpq2bBkH0UNfBHUtUcDwQA3WpniHKwgAQ
PDlwlt/R97SQHY7yeOsrXRjKN+xLlZmN4IKHzVLfaJRL609/m+9JTyR2/Ar1NXdV
JuIHweALz2788ZmjDG8DLMZ7SFKU3jzPNtk4bhklSx7tDe1owpV+Y+uBJqOyQoUF
xebruuYPaaa34hHqNLHUH2G29m8bY+1MiEb4EIkXJGGWv7OE7JUQmvjufE23mOmt
+mKRhhMyDN+XqdvA4mfIoCdN0loSpOmNw4XZLJ5ESPfjhKDStyHJ/EJ5GJ8zOqoS
XI5o6aphTQvqZlbZ/b4coGMZ2T0mP67uZvaoWY83o1iG5xCpMrG0U9DuHnYl6zOa
nbpObNN2frxV/b3V06xoiPwFKrH6CLGwdl/1avYiwc0/C2txfGFtZw6fLxXvG3R8
ety6MEL5hEZYbcC3Pqs9XyiHPMXoD9WHfXV9w1YUyaTNu/SZ5mimSMqa6u4IMzLr
lrcXcZ3v1coLeZ7uEfk8EopDGXDGPV/fIXjSt77nWw/XfzEl2NGJKolJaCZwgmlv
V96z7pSNiR6gDQ9TC2TU50LeEIq5D5E5VTZnh8vlB9ahJkl827oXmPtWxXhQ7jql
vrCK9P8TeXN1PoqbmSFS/Wr6QzAwA5Ue9TwK6ZbkDpSLqRdxdvldcVLL7s9TYETb
9w/UlHk2ZJW6gxU2gjb7aHit/KIS/n+tapHrwfWk3PR5vyvD6tKawWOm1l3WsyDQ
Zed2Dbw2IVnLIJBkxby8DrfR/lr6tWxkHV+sC/kYwjm+lOa1af43JJpUd+Qi3W1F
3cA/yOO4spqgn11OlrM1sLgzlBM+TQVKePr3bfHt0zQTlih8CFIjdNLYt8i4vZzA
oeMulY/FYh5Js2LXzBAG7MttTO41q7AhJEQ7VAzl+dI0k0UD3akRLuMNATBvWsVz
eFTQljBQZaBB2E+rr9AwPN2Fx6EAV/jQIOxi2S5jR0sfzrWTVzi0E1/usG74/H7R
lqg0Yj83pG53+6w4FKZYaEonNXdJs7kQ8B6vUBrgFCWzLjd3dbmpqjC8F0VZgZTP
bBzaMEqykTMzjVmM1T0sQ+sJL5fE31K2jUsHW7GuKMx3vHx7yvzzttwTX/beuNEI
/eHycZRkr3MSkfU6Ysu5Myx/NNk+8B9S9WwwkXK2dSZbfJtsf48TTsUcr9oDo9aY
yzNMjuKkaP+aDtmrk1lbpK7TffL+I0cTeiqUqH5m+wEDgaba2enS/k4D22NRxu8w
nZCQx/Ae1KaU2st5kqTE76I/sX08WWMoA3UWAVBeAU9BdjhfU7oVcDpP1UGeiKAJ
L8OLxhfUlI3Le4O2Rvpqq8fjnsmH/kOPIH8onQRoCskisjdwNDAwvdwGRVPFXe8a
p5BVx+Jcs4w926xepU4spWtYeFMEqkLkwTb8pER6AaVhdxCazvWWSXyzFo7PyJ5O
/8r2Ut7L7jHo/mjI1jQPHYXrYc0RlycpYfcaKiWf3riEPvX2JrXSiIYV0fuDAta6
VYDfYrlqZ4enpwslkSOeWvaLW9yI/q0I8S9I8bl2aWIaPTlt7XJV+Zks6zcY13XY
kuH36CnAjLwS50yugkC8Kv0b64fi1bGXcVNaA3cLJ/m68t+LioOJ+N9aMu5Tc5Pd
WJU3p+UvOOSTbAIE/S8h7nHVO4uZTvjq8XAtplU+8XTCIm5OPs3I57N/FsdiZnDn
/sN8tlUguI3wxPzNQweGrYjWXJctXD2uDrxJNdtgkPXWXUbZCGrLn4WL77iG5BTG
AcCkZkxmO7xxfLMX09ihtHdEncO2SFJbdK/blHrq2kEo9FYyuKWAk8ovf8p/DHmg
A4mtgXZdO/Dln2mMOtjAJV0HzdKp/ugXmNi5GQO3zjsCupNmmXrGXkUuR8CJnnqb
mTGnhzahLT/Wb1Ccdza4ZFgTxY7j7RrHsduMo6C6XrMZL7aeTUST01RWht8pfyg9
pUChTMXJgV7hAX1ThKRMrmaZ1NcP+qqaRyQw5UDNzBbOjs99igIIU5gBJw+ezZBE
FCM0MzARdU2fwRmFEr9zBwenQI1gQ77+sIrnNhtUyOv0UBdmsoWPz9ljZ68J0Ah+
0oXkUkqNxFc4nbbddUvCc3ByON2JdD0u0Y2jeAbupMkKcSpD+QZrtN/IWobhdZ8Z
Q4xpBSuNQLipIhEQdhuZeQBq24mFQmIIjnJ4F6bslTFlDfye+K2fYtCryIQm9u35
jqEswbEkLpzRhf1cSx8gU8groH0L2OnKQ1AfIvlI5KukDED7d2LqfAPKU2d6J7I/
/MkRv+ReSjq9b4SeMZQWTO+ihQm+iYkztHcpTc0+Z3D9+ov4fJIkspT/U6WxAdLY
mfyFLIrmWoq1Cpp1iwEKpxh9LsRb+6ItMKKZDcVUOlfA7I/oirHQWW5q8x2QTbXm
veUPG6F4/OMOK8LJfx/hEM7kU25AqFrV39BVzOXBmG0LbrrWYf7la3cdn96pirDi
c6oT4o8FL5YTFcO6SgslNtM4oR6NtlLCFv8jaLsKCCmlIb0FIvB+NfXACN47lrj1
EqIRxpgqy4PJUnou6xOX+5Sm4EUIDQigtWUmKE8g7GOwpu3+HrmCQtskIUfdfjV0
K8SUaASCwzgnafU5iwXipbW8/uva5EEn+d8B4r6/EA3qf27fxixUjauTNuHJURue
OpG8OKAdEmPm51B5iVofMLmq5+9Ttd+pCQINnTm9XP8tt03FL/HPUQ7YMuBdJC2+
qQwVa03tlCH4ELSmRBR9+E0VMiMaL8BNLlatzVr45gjkeH4Rh+QirOenQGTu2Aew
TjMElb/0ycXN+xBTgBW6nW+FwS5hhd2KevJ6utd5tXoZQonbl+SMDvlAyMk3oQos
VqO+69n1XHW/0heT2ILqoaoI+xq/SzrBUpb7sZ3Wk8cE24jynLIlVtFy+L8F9gUo
gvSl22cbgLy+U7reiZmHmDvOh2IocH/cZ8AXD7evG/y6IvI28MpXPLvCbSG8qvkR
MfQyM4Ijxg3mOgYvqBVM3mCWEVSUNzDMMUgXYHbWJQJldpS6wvBuFomi5cOTkSBf
lJJq7sl1dZB/A8eYCrdGkajo8H/RX5HwDdYIN10azGSDdjO0yTv1UbTYu70nFP+7
lRRhSf8JqMvnnkAA9hf3onxaWwXUBpEWDPBgGqdKtNAvjgWqztyR/o6mWH46FgNN
/P7q49BNEcehy7849Pg7ZKGyfULW8DRHIyfMAuNqVeok4DvfQYFWoHmPJjDHYtfQ
zOK0FdnYXXyoniJ10/K3NVVBC75gKRK9JxNNp9VgzM9h+B2jORCwFanyHg2NDYIl
gD5ZyERNIop00nXxlvs+dJwVRWXTDfLmihPSGn7KLuirmXy1TeDUJ/25NtvdZSvB
J+IU9fDFWtguA8FxzYHeksJ8nzSrB8hIThFTw6h5QqtTpokqFWvw0zDB03GL+aQs
/nvQ/tjY4TcjlIxvl87Ii+06XoxWB+SpZthCvPPztSG9fUCnY8A6C8xf9TFnC+pj
Lz7F1XUqn1Ros5HJROD5yq9LM13MToVMau0bHttSlHl+2L6AcxxyNOrZEDVaJKTu
aarJ8RqJp7Gzfm9i5GTjWWQdwGGC0URY5oOq67SAoWr1/tdSt7HM0cdmYzGBEbW1
QgvcxnWTja1eOgitJB9IvuLaqCYQLrPH2+Gb9DsUs0mXfWAJ4aqIJd2LOJLDVqOO
Gv3fsmPz6pJ+iVsbAmrxrE5FRXR8VQbqshTH8kyes0BoGjEThQLa141YZwDmTLvo
arlv7wTZ+IKhPxCvySTJkT9IEM1qqQEYj2ecXFVv1J0glTzyBmEHpWjAYnSn39Ta
tGGK+7SRErLY7XxqKKhRLO9hcYWAr511w2m7RcFW34j537HOzRbEeVEqDmlguaXx
oE3TFTmyuclcPuaJsjdqpfbIqUPqG96/G7AeSueAL948n1lusXM8vCm08jFzZvtp
HEoGtn1v5xEEB793zhxR4gCDvI94wXRhW5RqM1C34rwDi3z1aWgQqvX8Rk3chG3S
quRv5mY8+zxYEyrvq7e79LxCsdvyl2jdv5zEjPY1ugPt3GoQvwNJ+eWCzQL+JYLP
3W0AR8iJe87pDheaMob9ZDptbfmcN7JqWHIYKjQMxZ06BYlrvxJnrjpacLhxOJS1
CtG581Ai8Te52Jc5oVtz9gdQVt6ASVsC5kA9wPj/O+8G4mWrFUbwUKRYQxQQq/t2
Rou4jNQA8pKUdoziqkzAyvfXRAfP4+FUcWk9PNZx5ujxzptQyR5LgzG9tP/x1taF
+4LLicPKFSHh/DH0mtzMQvBHWeyQWud1eMYkR9bc09XFQvxk8NqUmvGae2XDDUXi
6FktwKInFAtDtGUJWlhkI8oXHC6MwelDTDmXG/+NZqLKdnCGa9YLoIqzgpnWFChD
S4T1/3buaG/Hd9I0Z07rFkX1N7DBzDctf4gQP2c3l5A8ubEbkeTxuZUzYZM8ComP
t7XY9+ADasJD9t6sR/ucBSlTjGvf4sMoZ3qDsOd2b1tJPXjKnDVKxWqKr2oIx9Xv
ipe7tm1T/UXp59lRptuw6HfU2PXTt283P/bLcDGqa98D6kMRS5WMeUIvhi/WNZnZ
4E+ynQ4+SnbzBuL44JC4O1VHECJ6KBar/xGfs3tieW7yfFGV3cNPgZKJPx37+Aiy
KdKaetiwwsXliPh1k2qMNuyQz2hrBuPYBgTNnk5p0S4UORVnMyyLhIhs8CBLGIJw
ARcUYMFtlQQ4HYv2vJllsN2u6wRxykLMA1z1jMF3peOee1iOrvQtZRxF2FIdFI0s
L6FSiNQYIxRZ6+srl4Oj0tQLJWI7lqrln3zOwt3EPhHBH/vThXUMXalYZQOfVBDG
KM0jLoDJi69/0FGyll8ax8ijrqzldMoXi/J9QLOIEhqNYxtP79IUE8UkzLmAbRwz
qEaLattED+oLtvtvorRAZdmxTz+fazyxKeZLUnLVJXCk0cn8Uhf5HvZnqcQnXFWh
1eYfKAg9hQP0c2qUvvYvroJ6kuXW+1cc7CDMbanzqD9oFK7k6mYUdIes8qlZkP+m
uyGFjr7aBxvPQD646eX79yTlDcfXwGg4HkiUfBjdFYvxiJdzd3UciaxA3T/4wrPx
OGpRjzEyr4aoVdOUqqmqSiAMdIdUXtd/GtJI2vTNqukuYgvyuyygsEO4TfXrQy7F
A24YsVh+tQrHzzBPxcp8ivfD2OYaVywkBZMiR/Z2ONHxle0M+s2A2bxVQBOJpvAL
NZ9xgika+rB0Tj3feeu1zxu0/hm1rC953ZPgs+uyYi2U7JwOfkF10qp/39Ndx9UG
JNtk3HBzIXeYO9g31T1ZOU+6DWc2JULXhAsD5eionKG/xLz7kXGpc+vnqpNIRw3N
aiy37twyWv7/WmRMSBCwz26J1bxi7ubP+E8GL5IeOKsyuYOunBrG7r5YAVe4TD0v
MnqrCwnbftByLjZfOPUHNrOvwCBvY44cXcyEZ6bRsN5Rl54fCEClzU07wtTPcV0b
yNWjHjWLlsryaWYdHenFN+9q2fWBrF+7g3/K5I8TnVk91tjuovUxfALiKXmEpu7m
XMU1gT68PNwbEWKYRJsnbiSDZqUAMnWufTBjXxaxCewogneZ4ppkbOtfjyZ7gX6o
+m6mwFtw0C/GNdvSIe4v0GRfhhhvmIkOmJSu1bsD8YM1nggCg75XsIdYo2RBBQXB
5TwR1Eoil3BYhQGTf36u/U96puHHqnTdh49sDERBuP5iVQl1rd+Wh38P5hY4xM0C
o/sgdv+bGe9kMS5AHQGjqOGp3plyrJ8Jg58w3CT3rV2h2EjSQhsXezmOHTkiZ/bs
EJXPP0zFtrmQxO8jPbirego31BE5m4b1PNnWOnO6ssOIA8DsJiIyNm1CdwKlwfzU
ZGo3ai6jmYttJqjc8BPol/nXBVXK0E6A1S+VurWKYmFkT+F7mZUEbmrIOy9zkSlg
aQxtVxcoKcx/DKa1cgWn28eXcG7M96bxm3wmghRxiK5LBM/DTXs1ap0yHOiOLzIB
jKKHAbGSOHFTwiU7GLTtLI/JRzRCD2UMYyICN7/uXZhgUhgasuNI8Q88TY3M6ghJ
qjk2v0jzNsu8WFH8rtCR4ajeXLgMVndcHIohm62Bve5d0Tfg/01hIJqmr85F3t+E
52g4e4w7JLSbrux+Ocmha5wTyIY6IlFJlVz0mqGSfZbZuAS/bnSyVfReV6d0ppmz
zjNxSGXQm7+v7l66vghlgFa5vF6ZgbsmI9E24X4ahsUCLQ1O2KU69O/woUYj09Cl
I+gpDn4x3svG+/EUWvvnOpzaNyT/FVQ6IhikZOuB40KVDw1Wtyjt9TczYYF/OBpB
4k5oaxmWzkLdT6m+6zPOQcNG9wStAvefqTUzpY0Mi5FVgj2wA1fkhfZLavdi3VCE
Hth2MOnLrsW8i2Nntg1o/u9gIgff2hvOMAgSM6AIoFli981Qt2sxTwNAc3Zrdl1w
XkUFS1Cbamdv6AgH85RuTjC98PbML9wguASDV7aOTItdDw53yz6+H/ZiWOvy1dxT
P0sbk/dJFnABpSkVXqZtSG5eknz0/pgvjB23Slx3X7k1+T+gkFHUIxUQakYcPeRu
iupqX9pgui9InlPDvOSys5siYyJ58ziC0pSb9tZ7Gw4xACwJTeOeCc37g2UNrQ6+
zWxGXHmpxYZSIh4hk/IUWGX37d1/YIZstn99kShPX+Oc8VxBKFUMlcmMbsCAgVNn
obDfMx/jU5xPa/1Ixdx8gqzazZk/onDfgZBFRWDtMAaX6ZCNc9YcjT0sYyl6Lc3b
e8PbzXcaaj6iZflMzPxGtB2NiQQugPuwRDibXjQv4lvtxJHoDzxCEC2gGDOF6cio
jxEwmiQblUTg71ALQo4ZGak9Lr+m7hNDXiTcNzuDZ9VE11spQTamlhy4gwQm0c5O
HYIvZ2SZjRLFAZVGddavfiypfNoWSJM9fMoMn2aHqFnL+c/nWD2OoC3AOLQkzN+m
kwVbrFnCY3LGMK+SJ/wRfMvlaiWxeAD4Qj+fBzwfYPO4O29i5SN2fQmjE4j6lt3x
EbPF8jyHta9txiNMraIgIMcUF9citzJhL5etkvNeP6n+n4UDxsPvr88DUq8KmPF3
SiTFyPitO7weV6FjGf2+r0WlXTRn5kE1l3leC0AbWd92GCV5sXsfQIhpMKzOZFXK
OdV+U/PFH5SIHbzoeAnX316B1LWG6AG9wzoDDfGSEKwf/ItqPLuqkJDhc+jd+pYO
N0zTeopdxzlEk/hTT176WhRGRiOwsQSqTQ649togpxbB6aEk65DeiQ4Q9OVuFHZl
0/k3IR9TZXQSrF3Mv8Vd1Oeet7nySTumakslztG+iXFAUwKWs6LNnjvet58E1j5X
PMz+zE7O7bFvX486EiB/1Q34GNNzM0hJGnhJhmLDTdZrs3y2rcU2ffqC0YRb2URd
Q8MK/x9zibA8Spka4urPK9gLDNMGVCcu9ihBsZyMWRbWmik2LhoNutDalaoc4EBu
p8pN0rFWc64dZkzyfpytg35WkLX7F8JnK/FVLQ1lJrt/jGPwQUiyuAPiLwOr2KUv
EBwn00vhYnWK3PzqrTX33LULorbw/QH/aJUUYl+KUbxc16jL/pM5KYNldY3E+TDz
/vk19sjkEg7ZVnhWnBV+prqiZn+EEueMM4Luak+/lkG3TQweW6pQ5RAJTtb9yVTP
+DHwjLEL0bIUkPkVkPf3J06ZkboIkzMk9S+MtwgL7Fpg9Ri37Owrok5GNtdXIvbV
wBGWVmWm+V8fOv46wGLievRFjpjSye49MMJKvUTojQeofi+F+xgO2+sMUmpyWAsF
gAwd2NKuIAOWBiAzjQNKun4xFwsNqWXsZolvpA9vc3lKbkIyJ5aJ1zkxqcMV044S
qlJj+lxoBJMtlaGu12G8lyMfoCmkyMPv3DQcHgxYZBx3FpulltjG8S+rRM/liZyA
Baio4pmV2CFzBe1i0c09TBzPm/jKCY8KZbo9qcXjRkydeX9UpWvzcFd6aaCokGrz
qFj2nU56rGIRMGz3P8l54RSPmFPTwbykOcC6CFKaPjuYsqVah/wXSr1NTwVyBviN
Kj52TKebsWIo5soVWI/RoCUSCzMd2JjYxXGbAWPgbWvinBzg9xHIX2HrV6vd2ENH
2IeRD+JsrC0L47tAbKeN7fxY3Ql6hcl2+bVHZ8MC8hHMTjYUSitBwFnR8ENctVdr
NlKLGgabB6k2ZNVoIXy+KtRhB//+XyKa0Nj2x/L4E29kQ/UlULUO3LzZEtB0wJmY
3BouH1USmmyslnAbQyOvz7UmeAZpWRDV04KaytSqwSsPxSiLZbUp1K5Pp8k3Aju5
l6o8vzW+4IMU8USM99vYg/OjTFEi3tjoQhQrP+8pR5gU8dD3+Bu/HVde88VT4sm6
Gq52W/1PlLJrFxprfc0MaOu1J1M/slbvyRa6GvLoevKD55whbMrjqLPIh0sQ+7VU
5IrwAZfuLjLleBxdYaEUlskTcDho3DXe6VwAaVnxddXfFiWhGjFI1qHY65jC5oyM
o4mJmfSo+MO+FI2SwAqbiYjZx0IxOeomNIG36RC7jxTMKQNVc5pmxJSheNHRGptX
NVBbJ7DB4216CUEgF7rnYABp4Mp+a7r4+TJ3SLE1SMiQUQyoanm21WwazldShdY5
7mqbLBc2ZojLfU7a9ILEUcCu7Tc9fmSMlg5D+z31+tOzqdXadjuhIEawOYdD5vKA
a6AR7XCMwqGVUM6CWKH4XnXdAonLrA7SNMecBI1gcL/B3PfPL5uFYmaCRMgateOj
mOISRlRe15HfJbR8Fea8Fv4va8lib7CVG7U3jUmMoVd8vWHpQB7GiYXtgkgRJJHg
7Xas1DsM7cUMHB2sL8Xl0KFvdFE8k0CDD/5lNfUxn0KYc+2zVxSrXDP6J0SneQPT
nZOtrgvs84Js50W/sXpqKnDkb9IOXRse84P5d7XQTWqP9dB8Blp2G4kpsCwLdU1i
Hy176hk9gtgx4I94WcNyL0HVu6J+5KisJZIl4IpM2XCSyEKDVuq9FKLH0LQWxtxE
drS1ngWOnIIdmHNlkKjtA+NCyU+8be+D6WD6GmDOSPFwHuY5jOMEf5qdAwT2WQ60
Mf0+7shrzi+M2hk41DQNDVHvo2Ikuq9htESACuWraTdO3e+A0fWQibI50e2/IXvk
aGebsmFxkM/Fv3pB9P8KoKBaC3fnzgpFCIiEvKXBg5wv2KySsHeThUifCsLjDoho
D/OmBxTvzRQXfMcytuYF3xNkV1KRzIWOPDPGIX9UUcBPnA/XVGvuYFxCNLquTnIV
GJSo1e1whc5R2T3VUe+Cn3hA/cov8Uij0bOTA04OE6tho2XgNlYbyrQnE/ju5mql
3keqa6HWAwjLKCNaf9V40xdjn248v4MCDeXRm0x1NoNvtY5of087GeroZ+dw5ho7
ksDYrD60XM0Zlrpn5V+1mcJdnA7JFrLt37g40QHM93xdjUe7+bvxFf9m+LpZWQct
qFYqmh++2jocazkBRq9ho9tmibyZG5G7AONKdNIHuJcETTzsZ+ULWyYifIwRCYjs
mSX+m1BTUMyC4aUBwxWjVnykeXfGfI+qwhqRrpIPjmtk4ezZZyploP0J7oc0En/S
GueOMiETrEWQiiEPQd+pD4MfQgcVbeXOrXPn0pD8ogASl3MilSWLWS686QlUFkfp
k+zsFoY3U5TdwYtoDVxlU58cW5Luzv3CLmlO82sQQyrgKjmNkb4PwrGv7N+Io/8V
MQZx/7OUDlzDKQpVwyoutQGyqYcVaG5s2UUfUw9c5ZQVaSHdXFvww1oFTDPpTznj
4AQXXPgdLQ1QbU1QCVFiJSmbIJfMhsiI1GReDtM1SQzSccmX1cs2ug2LwM3jQD8j
1vJSeOYutftGqR6drN3h4zmC534ciyhSyu6LHrNj486vXro87yvzSj88O2yKBTYM
KQHZCTiwGQL3dgCJVOVdGDRp23cjYwqKbnnsvk42lGto8GNrnOf9ntQsgVdNoZaO
BohKt//qoS9u9Cd5yhFEtedeLTn3uiIIAC1QNXB3D7VEgbausB3t1O8uUsJSLpTY
345ubM8vxzhjddb0PUlkoRMmrRWUEw4FqczTgMIu9dnBKXcV5BxwnrVLhPuFUwRT
+2DfXajw4qHFboyc4sOipjO3FBBgRe+AnUFL28XSyGQXE8QLn2ojI7I0jclacgmL
dTt+gI62J1pHEVJv5JA09FWTvPv9xawCVyWLNenicw/Cc/gGKEsLQmh0YDLKQE3t
DRKKXrLB8wXCzizAnnG8j1TdJ1ivO03j1ZNj76sShu27Psxlk8UIB9So0GDrtMSQ
PPg3sLC91OiP1ma/B07o0vmU51iAWpais6fSavB0FdS6I0MYJ7w6AWLKRVM3l/+I
xn5/UvB5VP4TvB81/i0QLN+legs+8HctCZ/InDttCE93rpnWMiLZ7zS+n14tUL/1
RKsc3xIF6mu74LbApuGKgREgWvldbfg18xbn8jZyhE6C2O/rfAIYaLzSb1AdUbmW
a4z8znaFA69EbBcvrlSb0NY3pW5lZ1gkfwMpVfzN3SrtTmk9be0Wy9mRSg3yrS11
EjmuLySoH7OSRzqOqPCzgTwMGX472VfmzYuZobreXXAZ10ZX47+pkj96aKsJA4Vi
1Hy1Ur6EvkpluedDwXfqJh7KGX7YSrpEDHMBQqfJIakPHt65pEL3cBKFcK7KZ3TO
90XD11nVGTkl8pMYqzWXi0vFYd+4ZsZ0MYT4HiqieRILevCWsUUWhOvv6goJoLv3
FpLjXxYiv0At71cuflTmnlp8+CODKGZewT4a8OKd+kM+kBoQin2ucUXMVBTDncPU
YqzUAScL1MWmnZIlBJv7vEf7rTjeizpuHl01OJGHQ2xLfFChmNFgEB6pvRBcecxc
KEBJO6MUVo+Czs7JkweR3ssoZHWhXRmpIiqYlY/VGlmM1XY3whfW2S0iJ/02EHNV
GtJp/jZ1//a6aqW2+rFLmUKxTjZo1d1UNgl873GXj8X89BmBmLpMOcSC3OOEly+t
hiQDONwc/LsI9A7Xqb7pCHa/8Wd1eGtDW5tCt1YX1TP2b43YUQgCQtqp5JweUKUb
xzT/jQp6kKgK0W2xifBFnr/EyNagbXqOrq1wFyoh5LrH55DCflivALGdIcQ6Fmlg
ARzCz0ZC1IqvnYyBMxWypT1atLwnTTHpC/d/k1tj7IofRgYbnaNkvJAL990Fu/Gc
bKDKwwNXPyMby1BFt3M4M5wd7EsgDDFguOsnCg/a3x7figMyFihv+1UhGvHEjatB
jihkx3UQDJCb4dN+fKoi+zF0OMqUN/pelbKGpVU2l9Q+0NAV1TSlDUGEbY85Y4lg
jO1E9iMC+FfHFY8G48V17CV7oXjAg0sZaUDTLfXb/6SL8VOixI5jX1a/7Z6Pzqai
2kNTaLeDHxzzTKI49zfNjV1vkCjGmJ6SI2ZHa7f4EWrkgk1MSHFjnApPmVZhOe+g
MFsytmWZWsAsiulMmxZtSUU5gMF37A5lPxWdlfQnDuxaw7YJLso0KPw6SALNBtKW
QV1K/gQCXD8H5IiyOvx4cj8FakH93KlBlGiAyySwlyBz2iScmxD1CyZ5f38UJrXc
6OkK2xU08W+IXBe+MVN1dVRSAI5cXQ3C6K2EFdl2rBkOVjTT+WayOgFcVzcFNZG5
IKzdlMREOZxU+0khF3xtYL95IDtsAGHmfi4wDqREkoHz7xvOqhOjkVld0xh9FOve
z9kZXmoC0gW7jMpOa3R0cFkQx0OjxBU6/U9fLUft+NmEGIt3lcouFfkeZj44XqHl
0Fmct/5kynf7c8ooKQVlL214UnohdhwoX6KdbFFjwzpGdSPiqBbJAeaPD8vfXMjG
F1HyRFAqrWm5YYCIjc4LovH+WSFLNbzZbcVD5QeLICNMhW0dJSY5om+QPH53bPnT
73jJ0ASWFaE2mUKMPWMW0ux1c8FT2X0SsEG1HiLDnJG2ztTV90VuMtRAcggFkrBk
mmQKb1dpY5ikQrmXil0UhyDACfkelN7TtQPNMo6mhXv5BTKl/ydoKX3Hm8yTCsDv
0D9UhqcMmk4WIiLD269jRygXLzLd7/2//btgyvuTRRSwYFG9O0pIBng4qIWsJqBx
dUnKaGEpizmSpxv5/n7xFBenR/aWs4+2fdgvTM+82doOoHZdYR3LGHpkqCdXJ/0P
gM5lhKOj33EmAt55oeDtHRW8iZGo3fRZMQQoOeqYOZJVRvxF95hok5r1EaqD03iq
N5/lVsbF9qsJqTTUpYrfQ75bSz4YybQE5qvc1pZ4MJ8HQJucNIZwhoCi5zlpJ6PW
mdcql8RiqzRVbYRRxT3+mzglPtMwff7x1/K2Hq/r2IDXARH/XmVofNQ+gbXbykBc
79RvemY1ADu03M/+Z18gnp1HhrWU3g34xtMAgCbD9XI5zsVQEZIgRhI4NtQenLho
KRVx8JHtekENyx3uc29qWvUQfN2AAmbldSVK0BHspGOK5IWZ18Jv7VRrFJ3rl4Xn
hn1ViJk4YwvWxnxXLDpGDgbyqCwLFk5b6d7X/e68Yf8rIMSCOdNibETfpL5hL7KM
a3u74crAEeGaPsiSEG59PPYelZBFBGvzl3UU+OHj9ORshKrM04JNsSgHfPfSXwAx
9pG5UdmdOSGjYjpZqYek0FwFol/aVJwHiZKQLU9++CX92WOh0I4VFuhg4uZ0ctQh
EC1eehURGlGDIM0ILbHe+iix42thQzbZgXyPBmMHvLBr+cVf4gUsxEROHlaSgyJi
Lr0bMrva8uKrAl2G6S2Ke3ZDE2KEnZbfGjVz1gqu1DCh+UQ8CYo0eM3FfsvoqqsG
Z3SuuSmiJcEBi5tDsOkghb+L1onfYdf6OW6d7MztGgBJWekvsb4p16zz+j28tuqW
kMtukKK+6jr2cCr0bztPuJVoiavypbKVGX1/WNgnWvMjHLMpiy673j+ocoi7GzDY
TS6Zxz7mhZuXJV/sBwkk0f4t/oVVK5odShg49LbyoTKk2GBzJ+zjzBZ5MEq3yseR
h/BPw2uQjDhOk/z1P5g0LgzorDPW1UrdyfYitZvSqzNaXYNsyLQUlNOCCsCaExuz
ov+cWec5M96yvLDPbDhetAm1TlHQDSGtuwakitUZd0y/45eayIp8lKNjOgyavh68
MbJe6VkW5byucFqjD7AJAdSJCwjzXUH1fRkT3l55oRdD6SBoG0532HpzcwWv7TF7
aTs4j2Ymb+WRMO8jWqLmMscFUxDJr/j3Df3O/R/8b9OOeFFJ50spL7vi9l9jpwQ8
bGrfGBuIvLeYZLwP0zICLGu7yPZnTqVTx0s2tYGVcppuVcLiqos2qYErLoP9udXE
hH21LKxO+MmjnSXpO9X1AXOowVllkNfC4HnSqACavlSOiS9RKUXPKa0+ee+9v0ep
dheLN48lIfs8I/Nm4PczswNgEJ1Ecc3I9OI5htmcapJW+67k+pZb96igJid//1R/
QfwZjiI/siNuN2XqQZ6SsEJE1YlSxjv9WuSbeuQE7jFqGwmcMEKOiUrQw3Dk90CR
iDbfdwh+sGd8Qy6IO/8rbqe/+8Wz9wsWbxg07JJm6D1tQqUXc0zf4i5jQdqqFtFG
delsDYENumbItBhgMHbQZl8/p06rAFKRhgoXOBuxHyaQS3slNdZFB1TCYQLapgDN
CiWX0PLPU7liMTsReW0+BUDapGkOQWlElc2t4dxQYrM7okCQjbeYYHbe+sWtlULK
5y3zKKEvMlmcBcFQZaTY8drOEnCSA1SKB8ZRs1vHF5/OMUGZ02RsxrJVRzNDVQO8
nPp2W1jSRqZ9FS33CgXYPs1EzBPV1aH4xRbrEclo/0ZA36Mx5h305qoyytMTxEEh
a0C50ryrVaBA+i2wDUVStCyaUiT2tEZLrAvcYQKmAHaemlKInFx59Ly5aklPOfgr
f/OXh668/INw6HMuTgSinLA+pqjZ1oP7GAk43ZDL+7q0GuYH0BpTg/EwWt2sQjTg
stAbgCxNRfobJAxFnRRTDZ46BSpkNio4NHvD68zkK9GpDuzFfAXaTuTvTxSr5XFO
h+Fz4U+EuCUmfkMPa/RQpBYCwbF/Ofz8ABSBGJpKJ+XyWvLHFN/V4olVtbWQi8Gn
HqlmJg4W4VL3Yc2CNt+L7UPWrJtWjUY4iKni2YznttqIV+8M8g3sr4EwT4/oJzBM
567TXmfABevn0SUJni3flGBi/OGurTvSwhslam+Mzm/3YbHYWpJPKrtxtB0zCx+O
pAM5BJqKDwAYdC7l9J7xMazfV7kMV2ol4mh0hvYCcmPK9QjMGB7hZ0wxCWtnDbZ8
tx2hOHlq4S8DuI0/qRYByceZEANHXPNq7QZNuhraRsPBuYWOe+d21z9z7emWDYce
231VVkL3J0/cXDeJtJhN8Y6WHWtVoRTplYdGJGCQr3WjA+odZv8aNvmFcn10GFgu
+r7FGhjxBzANu+HBQed8fcsrCyVyH6T1UyELHpGeFP5cR0H6c5kxu8apskupVtlP
Z0rm0F3FQxp3oXrYZtDYGiI+21ArjSH7oy5KiR1zWfQVyP9ulA5FOirS0/4PwwQ/
GvkizRKwZTDj7eCMjMoBTwI2Aasjtz74+itBQswjLRUApRJHMpH9lQXYqHEkKdvF
F5Pyjkzbr3/874RQ56UUCp4L7qqPrd9E0UJ62sNeotZUKrqpkTCHErQ4pXEXIcow
JFFR9dAw1MokTckVdfux8m214UE18aVOoRskJopQcsnOMSQgQNpvl9L5/RYHHl7a
OoyABgPd47uFyVM5+/e8jpcw686yn+rK8OJ/5u8y6TOvQdCV+//E2u/KMTR+At50
XZ5dHh65OzgnhYprkDJ1GW+cBxhkb8vwIfUmg52ptA4SR0S6/2iUPzH8FRfp0OQj
V2ti97qyMefRsO1HNG5+UrggwkRxkmTgEAT2MDACMWRXAq+k+u5YwwuldnPmy5Xt
UZecC5EWkBsUZgsMwCGuenR+8Q2Lk+xItAQiAgdcqeM3i5tHhngVYB77CbtJrwkp
JyvYzTQLzP4M0efSXp+A91cI0UDtn/W836dQkfbs2jplXMCB6s4B8GkMt9njOVUv
EwEBzvkbCk2hnnDbIk4qfsIoCyIIL1em+sr6mmdwIAhMAJSiNA8piVBhG/8vZyt2
/G1vS4lMUdzFlRREBtTbSHSGfpj3mc2kWk6bA/F6DY/h3f6LD7CXIcWUL3W4KIPZ
zXcbF1AQ5mQneg3/Em+FjsW2jSi7oSinIX59iaNHKywHVT562+jPlBkHWUXWiIlI
Zr5HmyhbtZO7EMlLUYb+Pr3Hnbu0Yy7VlKzQBmUdLUptVCdLsHFfTtX7v2+YsPJo
k03WiT5jqSxWJLwKyh4uX+HetoAX3gFMHgwfeuJoThfW4+QFFmDtD9+z53K/JPdP
6VetkABzl8th1jGXc7UyZJAnrLAZVIyr/MANW67yhZAiZYbU7ZBxPks4/FkbXZYX
BdLmhvk7zXzE38vkqXbZyn4EguBQRgb1iHNczZ86hwGU84J9pLl03B+zXUe1XpYa
aScs6hJvMwFfTke+ggDaTvc/o77NbpD1FePDt1Jn8C/Pghh34GEMSo9dUC5BpiyW
1aiBerokmh6ZYN/4ROvewC8DaVmmSGqqOL/UwCN/XLW8yZ3AcxHsfJsz91ezayoB
Zszfl1sgCeo8Da/x/TuTjD+583MvBMOVlV2/vLX3WoyAup+SwfzD/E8KYay2Cxpe
ae7bpCLSoNAPV/oJnLEZoZEc+yDRDRhp3+obON3bTranonzLSWUcgXaqatwUm/gV
tglrcyAorpSVOOi7UgSr97IpnHA5eZT2jlPiAFuTBeDZ5VTXHCEM7e4msd6zt5B8
iDm6Yedj9t79NhylVg7dB3fny5KW63AU0G+LWPGIvX1KJ6KcXOt9f6GFo55KgJhQ
O0Kj/6tX9a4vhvRZuLZ0OG8AYaT97oIjkJVJaESD8Tp+FlA9+rN1yOAiLbZzfeC9
RPW3h4ParnRo0IYhPJ2yh01/Yk5g3uTdNxTU1irpigNr1Lo5BO7qf1DKyfAW9l6g
AolLi23X3LARxuGikDhmWGYGSOi+BNanbsLw4H9IbJZI34TqV3XqGetwHgnbvBkq
7YeemoM6E7Rza+Dc7WMi0LUKEN/EsYRjapH7TjXvsHfQdjQOizr0Ln1YVvxMBozs
Ok0+KFwKxFeCVbxMde/lqAiefJxJqdTb6/Qt2p6LHUeTUVSks5RnYyoUPLKjdLMY
24fDzHtMOc4BxA7xZNi+b62btEjXp5aU2uMVEYD2mhcnV/xRuYgTnXVLiuikUDAc
nE49+DMHSedyTNz+ivBw2N0Pe3DR09EWyLOntAdUHOzs4GTvZf59ahHqyNbzgINt
pl3si2rWZr8JPSZBlxZuePNf1OUnaCXcGOFkWqSCx3dyVaMjjF/vKzkE1Yv1Y6cX
BV5cAPhm81dZxGjI/My4eAjbE8UlBi9IiUMViaXOechI0CEW/lFtCHS2zWTEHnve
iN9Zh1LQMYAVbfONNBJ3vrmwzXCNlgutXDjZ2kPpmWoYovIFFOE+AapeZTgbV5JK
8GnGOm8meARchRPAy6GkBXUAvk+XFNn5Qclql9t3ZhQAui3LB6BQaNjS6jaUYTwe
ddWqUwNfFSm3e6cSIoX4OuMCVkFKeCpzVUqBjgGTrgCT0YKmgjIdRKahD3UdjY0a
dIgdkExhm00m97mKCI7fl0KWNVZLO10B5jcEKJRFxXS0C9hCDqh5fuTMuVLEdAbQ
/FJQHaVPky/2uRJSVNi/pXbUNlqhixmE7AsKSNlwQOkfVjIxWHXsKyFOELQ+PgN1
2eRcuvt3oXRAR0W/8Tw3NIRoPmy7YDtHmXIcEw+YVcT51VlUqbdKgZOEiQxkKlc5
oHmEA1QG4+1HKKaJ3pFVTArHV0x4q5lHrTU3LAeVvUSDApjtkR8AzEHeTDqNYBX3
TwSR3tsp4/FH0ua2XlX0w/IPSIEynoGjqvBDNK85pbvKBzghnQw89D27RJxe8CGs
inuI7vbnBSg2P0bHAdYkpkhFd1R6QDZZjLSCXTG6b9YO2lJMrDFc+scWvd9TlZxe
u/xRaPVt0g7q4mb7ILpdDBXYtjJcbZ6riNuw2gj1YxMmicdBodhbHf860PRPrJTx
EQODg5DrkvEzCiy2gFISS8/PJgKSITGZEXZjFMBcQCcb/sk9ZaahUDJ15l+ohatg
ApCIHbcYE3WUOcNi9uSDz7Di0hL04Sqmv0B0tWqSZD93lI4Jz9ZZPgSkZ/D/aNeM
fqVW9rYWnJf37oJSaAmfrUt6KhPqJy4QlbIkEzYM575u5B3VfrCewfCOqaloYYZK
1a5yh71FI8+I7QtM1c4NTntHKGsjlT94oPEgVOaZ7q+isj5G7TXUxYKlR+8dQTEF
oBP36xw3X5w8XV19TXggD8im2JaGFYD6rsoVjLZ4QfXDmlRtQfNYYWSsBeBiN3Td
jztSMWhGntyrXRGmZv5VmUHL9fajrfsT2nFBKquPLG5GYue7Kook/0fGNKtFCkEh
mYFxA5/Cw4S6ESHHXNrPfGmcbFLuWmFBq8Y2XvzXjMVSfnN4qIPy1IKnMxYL0rEj
NRM6t0mcNcYnUmrFZrFzAKdLMu6xJR5FRy3N0+wJEEqI3HKsb7N/0PjRrb2WRo8P
ghZEcll4Sg+Zsbyx2rbI7lYNYW2PW7vdYqC/1aGHDGbjFwjwNFSHaCV+txrR99aa
1l7U+DMwoQnkOSlf97K3bahUn2nHJ849hibAnGXZE+VyQ5ZvNipoqi4CE1KOzA6g
qqf5P4eFULt3fQGl1pMR44xlpdNDhdroqzoCc5ay50/PbvrCPrUeT3rJuPrvIc27
ZAAA5frnFGvja7p5Br8BJ8OKROKHI4hJWJrlWVjtE0p44HS/cq/LFh6g7yhrOUE9
pSY5mB8m+Msohh2/DQ0VlcycjUoqYmwAzGDpplGRXrWP6HFPT/PXKjZacR3XiLlO
NlcjC/1+4WLxbSqVK2FSc+8OnOfBdXAq8Jo+fE/vvHQRUuhf9lEijDaxNN3mITyE
7BUG6xpzWat0+oOQU0TSHaJ9kFlnN+88Zh0V3PvVzv257NvNbWfwk7dtOCyVJMMs
b2t7R9A6IyZqdAfoc2gZncfD3wBq5jo5snitOHcKxhFIYypOicIWm6BZ4+H6ZDa0
tEalkYhFEq7pQLAMWBok9VdNyl1R1adBK/8yHzKZEJSvcNRNnbcw2RE23BMmNgOb
O+C6J8L7gMPDTmIirHRv27Jvilp1gy1NzFu6kCnNgOxgS/NxVuHOJeXumxJ7ce0M
ElGa0Pu0Z49ntnRC+K8AA482JOXr6ouUupF/Y2EB3O+7AHh4tfft80eluNX7ITR2
XVH6RbWUZefgaC04GqIxHkZxkO8OPmyv45lrGUzlWEmxKKByitWmFRyeB+CCsErX
4Y5XTu+6/MBt8UCuwPIP8mTHcKoTRTDlSvqoyZaygCPiY8XGA86cZCyScnXbA95E
QeMDdbF68C7yVuS2RySbB/V8Bopxl3NUcZghuwNJpnY7+OFgfnXa1ajPZiQ+jKa9
a2b+q4/hbhpE1NeqIPzqFJm+LnIwg+EIDnG6OwWdu7EDsnHFGgJxZWMdD+4fu7vi
wE/fX96qHfflHsknJHtNvgECpbYPtpNxGrPliwNPDv1wt1VSmZgceAqWAgV2i2vp
5CoL2ByLc8iAEZ1mbNLsuz41eqGQ5dV+qDrK6bRuSa8A4l6MTdYccu1/fLBTYP3G
vqNwndmh+DZxccd58o0eEd0h3w9Y4bk59ymSpdb7V44OpRUFeo8MNPLd28jPuvWZ
1r5A7Qj0b09kzSfXhNptDSnOC3OqDB3Tl3wcNsNkKSMHUXVC3bcGOXR48yr0rKyu
afYDHOFX7KWsEgownKpkim5gkTfdM6SiU+ZmOGAumQcMPBkKjY8hPPZkhziNliES
EL9v4RESvT66RBvTWUSwlSabwO+k9WleUDtR8+sksB9hyomtIcl8JK8a3uIc7YkE
VqNg8vktw/H08HpfGw9cHTG9RBZYBEYF3hO5uZzgY3HLvPEODJ7MioHrTUh9auWn
+39v4Mb8VC7WDQKStO2MbV5AIqMJGwgq6qM+BKggVLqzWHO0jjTYE7tTYmdrxhJO
N+C1LhywuRW+0wuuKUHhS4vjVFUhmBY+rRZ7vDQqj2lBgLQN6COyt7B25o6lEQl2
IHetdNgLiz1hzbtMHqJi8KSYkVL+og1+lMGMVsXrr/RwnCN4KRdX3HlXhIhvlcL4
JxoZWBZaBNKtrRxGueM8jek7UHp+Dta1BC1JbvQDzBoy6h/XllBdEZ7zPMVDkajI
oKpXVJ8h8D37/feSwSoYX/TvjjHVeQqPJG/xf5DxQevJTlLRosFq40OxPw2fvvp/
o+EDeeokUggVtcJm9XVJeF6Ei9z770HAicnZ29NQucgL9XvO32dLL8Taj+krG4zQ
DfA4tNKFu+i9fepzyHX2MubGBt83EHijQT46QigAHEAE0BYqgfaxRgxpR8y3AkDP
eMO7rbtBiLXGrZKJMlkS/ECHU+80SCMvYFfs+iNZEtRV6r9jgZ0BOvh704d0rqkj
NyGWhG1hUN1tJIFqYVvZ9fDuTnHbBD1TxggsKjofHkzZqSA+GgH2cZlsn1Zuh+EY
QxtJepJH6klmJ+CxhOnf3t/fIKE0M+NjXQaFXCbqWfX7e0V5pnsHkqIbH0c1MOyg
XbqEUuNKx30RApHXXz3BVm4N7p6mdAn0ZFzGwcXNTm7S49FSsYOHo7mFej8ewMk6
tn8dXc1XvfnAZjxu2SGz4wJzRWeCyp43Ynhc2qr9JeiKs1/UjNP7wgkGCkKvLgRh
Wy6ThxTvalMLyVl0Sor9XNE40Qp/9jLjFr5eXZQq6euryBs6xTo81hH/eK0NqOYV
cd0rzd72dv8Tt+spCO0BDnWEOngPf9XzwZanZ1nGKWTqfw9X8pG5OtimnRDq+9N2
rYfaGAFoTL/NJK9lx+okOAZqKL+iKabAIsGvSovHtZnE6+prpl3yVkajTJ8M1A6a
q/5HSii+3O3fb7aSfHOP1aWIbSfi7hDFYe0D5C5fuAoAZn/yeGlFyJbzPESOXwfi
dBppC8UiALKoO6TmiA19BOpYzEPVldKPCN0mOGUIZvq5kA5VRfHXCPWjAhJKNBnd
AScAhAnQXfDqw5wMnV9A3kq7mNGbH4ZaLgTs8HdVbLarc3wbeNX/c7MGjT8HwpOW
fjfMfARdS+ezdLct01ODL+M5TSc3w3fIwQOQy164GqcrnShqCN1SLmHp5T34ew2/
JWHhxwc0WRnl7KN/RwH/QzLcOz64Orb7GPLxB1qDh8eCpugsPcqpTQjsN10gXszq
5avx8y2U6Ojf090cbxS4192FQlFNFfEMoPm9gqXHnxXgGZlBTj+kMCBSjbrMsEqW
J1/grnqgBGg2SVQlp7e5uAHCenOO+kxtLdBXYWr1sRTI2tsMiQFEU9+t08dJj2s6
vvuuSiq/rgsMrLD+2RaJZvuJA2W/ZB2nJ7QZYB5DuvF58f97gHd8S1HX8qJEa4yU
YVKXvPVHc+fT+DGhR3tuBvjCoRWNPgBnzW5uFFGQAle5+qxRyIgl0vt5lNDp6COf
tWJtz035rMUMKTpJM8FpRe6XJTU8y15VjdK3Q0+6tyGt+cJYGshRzjsQycYQaYtR
Qj8MTdeYrQVUSY/i0+otdN5m/wTlEv3dfxXz/jXz5ZLDoKC+HoGHplmMeY9YIGA+
563lk5i12Gd76z5nn2yam47W5lvOgDyslgapHz8IE4yP6VQsboF69fu2nAvRR1WL
OfIDsSGTsxSi0fWyj2Sx46eGI16snaZF3Y0VgyZUVPqpNUZF6QJTmIC1az6Ht7va
9Xu1i8GJMw/vqZmNHTCcLWwUY4EauJTNDaYNi/UVn9fAeL4kCMAg5uhb/bkpX791
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bHrWRX7B4r4EKgvp3JBdcuDMO6T7RU25oCEPk5GCTn0XAh77yOy+gAyta9rtmv9t
OsELfi4IcvfASTGftsXNrrYQq3xvHLrEVpte/MvCe989icUqcDhKls7myZTgpBZk
JasGagMCSsaJNEuZ4UfPexrT09LWB+fRJ7avEXLKkJGI3PWh3rUYSv9XLh4wwCtZ
RAfoOhSmYn7RO50V+VZkMTpxeJdLxlV9FyJCUARn5IRn9Bxwnu4wGQkSQuXjMK+Q
cdkKXkYhWSiy60t1EkLbKwxlh9iN4N1iVKsUpMl17X14Wo8JNNlUoKHshZnZtwOC
lW3s7ZZrUUmKnNQZFJfS4Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6496 )
`pragma protect data_block
dxXMag0mOTairZ2Q+JKGrPtXrqWIdeHqzecyw9+HkTSXyVaDwyGi0BON/xbmV1eC
a7K10oY9h9vdxUjzm5nOc/AYAMZCVFy2OzyMG0r2YLHzN7/QVgcexmZ/rDrsZlow
5cBx1iT7vaV7MLPciKp0MAy4Xps/ovQen2OLWPNH5tB2kSHr0dHcHOIIclYhAZCY
FSe/8bixZtYMEhI+DPOFsBgxD6WOPHkVQRGptXS9a7NZTILWOVyexzTtx5kkYbM/
zzGReAw22cgPZRRf2bIt4RjwuKxRM05jkyZQ/8obVRyujWBxNI5sbuxlXCasdgWl
NqGPLyWtukfpeCQpagN2ny3qZpdCLY9pttGNhPmeNyCB0MlZcRJ0mTAgmfbBwXmZ
7L1uM6qwvPhNcZYfWzKwoJtNQqnPb/o7BFiuJqUhcXeYgDN4MuAxhPwVTJzy08jA
a7Vm2gKW6NUwieXss8TFAbJ2U+oDLrazEak5gTY8R/OzPgNtELESxjr498VN0YbC
Z5ljwDlHBT7EnEwgWMpnVtX6WrZ89t96gtvJxRRqf+xVHCGAonEK2TM7U+rEwdVj
IZMfGdENQEaBm717pyTVpyTUXVT7bABSfbPgCg7aTcYR6+EttjH+pwz0T9pSCiKK
WS5JK2HOB9X1HRCeD6xVpXPoeHzwa7vDooV4NPzjR+4jXdAggnkYjsXZ68G4zF76
v/wycSVuYfgRe7yEaDAi/GCsl05XWdtCfDssVyZVfK0p//ihJSK0+ylbZbgWwngi
m5OeRRLKkfzzzjnT+TG5TilZiFil5ZCEain7vRu38BBWCAt2NYNQMislqrHEfBwk
VZwpfhYWYEFLyTBg+kz+SNIoCWLhUZE9v3wyfZOeweF/EJVfGlvG3aUd38BUm6Lq
wUfw6BT1dm6UlXTZrBcOcBVLyVLwtnjDZCT4PMTS8L4YoXH33RkRdwnYQK8fIWTq
+3d5TyXR1Rc/nKGuWQUo9QfthL3NN1QIgRtlME/R4JYyT2cmNx2sp428YQBZ+Q3k
xjVG9Tt7BeW+I31KqwQJ1/nMz6V/I52+ex+SdvI+QolZE/lf0wnFfjF08RlunHtm
Hlt5mGxjAlcGCGD219El30sMqRjHY0Df2yzoo/XKqPSrtIQeQo7bLsFrAYDhQlhb
up1sVsw4K4SDIrYZtJOTO6xtwm21nFwe+p/bhmq+FI5zoT2jVVQHE24yn8vhMM58
7zetZMgiTbEt2ySr776C6wec3xTIQpYl1cwmghfixeC18uUmvvjYbJbRg2OluWx7
ds8XK78fvgxuqtz267MjVESz+C5uOvvmh8jnl13qVwoMY9TlPGqKvsdY30fCk5dA
vDlXEt7gIdF5NVlNcttrwD3900uTpYsvppl+wM/Tsm7DqLVDsvsMmPgUE8kUl4xW
AVSA7ZbLiW35xTdqzLG5HSUe+ZoBD22kOO4Gy7yIh9irKjO0r/iWrns4yWWEFn8z
h+gW32nYJgY7hbsqlisxxWWfO6xgEw6B+1SSbuMlgGcvlcsTejL54zf8wQhA9V8l
gTzuB+akk7C1SN6AE0mkONjpxepalvBRni4MfW+l3l/HESPsSuvEo/oaCYh3lUl7
n7UyPYXMnmDEEs//FabBcMcHHi/gjhcO+wcxKWX9IbOI9Uukg0QDyCdXXVUHrDC7
yWHiy1NHNV0eHbIS0Co39cc06d9eP8/gG+Pdp15m/+Ny/tKTxz1PXLgRs4TLSSDy
AQtFKuymGx8mNdRoSrUqHuC/yUIw0pEAWDFOU7020fCtkEZV+yevsSB+2lCjnU4P
3L67fbFT3099OlJVVOZ9TlzpGycPecfVpQJfkUJjliXMSP0U910kQPif90mStwHE
mi+nOGDu/UXZSbwx7PEKXnrWscywgWNsVTU3jXLtf8p2MinSQZvrjZd5I152+PT+
/4HQOjaAEDbBfrBP7vrW+iwLKgR9R7+/+Y4x35t5b0l8U9qsmqNIvO9A48nurpN+
QQ6Qvox/T39iZ3QR6kmhdNCe/fgbPLYK2F1ga5IJL+SUUCXlxL6MiKeAdKA8bvdu
/hh2IWMZNj7LRzcaA1Ex1uAfnitYQhWocSDb13mkiJiRTH9R8pwrCK3SvURC9goa
AeCS2of5oKgaMuDqY+eJEZs37xB3oRaOYzf0OgvoOgRfY7D8Acdt7BtPicLKRJEL
2wBdUVQJ5izAkYAJ+Ffu8XUGYT4jTc9qGT+2s/PbBmHDd2JW1++qY9FfMb0uo9rM
rtEwwpFKGF5tN/ZtB3KaxMGagF2x+N1z5XP7IPxA8yqzn/fQ7zOt2xdZ2Hw7tlqQ
1ExHQQsxFuEVLi4rfwMZEtapz/jKBtr6aUFWa6pXb5CH5Mi7K5T8EH/RpA/ytn+2
wn4yQXy6xetii69gYUKpF9W+mqTmUicdHEeQQk6RKwRKBtMML5G3a4jNaBGbfoE2
xLuJb0nj9GlatSsbkDFZANxqdPCG4IMkWFB1v/Q4pYW4pgYlqdA2AAkHDHHL3evM
Grp0cjvqSXf0xFg4qYJu3vep4QGrV6EHQA/wOHEnavpofUQPzoecBjq8xdKYVFrf
l7AJXNmajxeucNEIGpdzaaK8hrjiA5gpzX58oDt+Tc2gLwkyVRajirFTtnPdW/1o
v3cbQ9SJ7nVFdcBmZ06rDWzxuq0P0BHhEuNJ9KdBUllyAvuSDvc0wT2asgpsSPfO
g7cFTqY/+XND9GPaKrPFmz/RUy1kxwz8CG8XL+zTy7PzHci/X9BjyM6a4VEFgtUJ
UsRmakKrD7pe+v0HWnFFT+pm471p4wzsjMK2RQy769z3z8i2zxl54hrWbqYRT68N
odJxSsgEk2MQgmVtiU7lVC0WXN7KvNdu1ehTSfJhj2uVuyzDV5mT/iiwc08KhAIg
vPVMGyOP88ikIxF+rz/9WGT5ss32NBFHMyojoJwk0GD+/w7ajeGaLADutzJrllZB
QcwVo4Iji/C9eu6JfrNB9X17qivcNydhfkXJcH2c/jLFasbC/C56l7XBLIF8UEMJ
GeYwey7KMY67D0CTLsP26uJozNV3tca0HcGZ8g4DOTzRZ2PTrnJBP/3fzoxXr6B1
WBmowQQOtetLMOxiQzF4qbtxjWHR7kni9VP8aOBnRvS4zMPbaTkb8SOL5DCs6uOQ
VPGxLTkyKjTmirRm+zfDrmxSB6vYtn2RPgFdRtsGdEq3wbF3I3YpTLjeWkh6pboY
+8Yw2bo3WWqDr1gRJjzfnfNjP45yXEejlpAdLNDiW0I4Xe/J3b8ZRxHsyqUdtt91
ghubQKdHGHmqjglZxG7Du3BV47HYFEkbtIjRShjEd2GjLLkhJVU7qAcXxQTKAC8t
R97XAeCdyf926CpoCN4I4/moArmvRgVBhuVwACq2yXtwdF2sk0wWthcXtSvctZmq
R1nAox2n/kvT+9amhInWAWHfnx34/S49OHAiOmY35/x38YJY6jJK/ox08wchqQ0P
XxLFowtMy+MHIo1qbAoFQhhTAwtnf45T1fMp/rxomQpOHeO+Hp/f2o8zVSRWMInn
sC3mEv3NUTYvLBh1lnHztCIw8CBRcaIeQD/tMAL2e8UJUWdaKTxIfhd3zSyUd0HV
TUEx2H6OcSqJ2BDIZxVhq+5mbGqC3GjpsbbELBRx4oMQl6C/3824ksuZFdidtL2E
UEonp/o1q7J1QoiyvKmSYaqUlFSv0MDzx0fK0k4Z7SVG3fPhi18n8GWEHxLJe6Ci
XYMqYfEtBxYWITmhYufm2moHOjfWvvPYcnIrite2GDIlLt/Dt7furJIAwZJ3JztT
1H2YSKE8Uz1TnyrqYzG3z2E1lE5lBgsMBijFsTcH++kaKyxGJv8LbVmH7bh/wpwt
Q0alA2hK1RxHCPqGS7wqlmbT1pZhnmSoI4yFG6pqVJoSb0JmLR/OUPs59que+NlF
upMSuqMkNE8UI2wHalkOoQqLzfydUO2Pf+im51JGhnk8HcZz2C8ryoSbmoUbfrt4
rIrSd8BmMkf1cQh7zMKzzPxOlsbPWy4KGslzqQX7BF5Hi/H7iShsz3THG8tykbMh
zmHivyaKpSODQXLUrkfK7Fnt4Rv6WGsZBO5qVPxI1w4iQ8J8QMra/sQBu1npFImu
7xQXUhtRBOjX0Mw3KwZWHfK8Ok/d0eiaXvzLH0e5i7yknnzb0yreWR7W7dMLL+NI
mp7K63P9ocWXDZ/nBewn5kt0UkmTe8qFVySgbpfdcvFi2kh8T++X9Eb+BpPx8sN3
Z4LRjxFDu+X0mCuOqqn2cZ6S8bDg6fVyrjZvxpwbSFyFCfgNzlujAB7Qyk2GnaAV
TA1JjZ8VODkrrozNVCgGXHDXDUDd0UOvv8nKGmEFThy3T5h38W6MZ123GPGZk9TZ
tuQ90fTFYmRKu09HFels8IlwIr0F/yxqxg208MLmyrfQgQvVhz2ynnFcxTDLONvY
iGZ7DagNKu16AccN+cEYcnxRVsOGhI/EMI3w/xb1eXZmR7wCwYEJ3DEd9BQ1d5Lb
J9PH1C64a69PwZGgonMSsSVpVutmJdDCRXWWmM0MU5t1EetoUizLfCT6qspYkdPS
wqa3mLltgtKF36PN9Zo49RQmIfGstpG6ZcoC7j/er9NPTwb971iBCTrY6IoDcq2R
yOZI0TYCxW5esNH0D3Vsl86L1oYbNg17vK/Qz+BItErUNGF0tHIsKGJXpO+TnvvG
2hXCoW91PFAn+xBG2Hn45GNeZHpABmkwPHZcEGA0rHB0NdSUyee34hbDxuG2ttJu
SI6ei2Z0D7rAqLGEdIQGb0L91aG/K+YLjnKWLilqRu7qdpafgmrC9Cv0ZxG2n+Nw
h2VLG7gXBXlIhid1uCerkVQXYFsQfdajYvfzrhKgFAoDj45M+9DY5fF3Q/RENIQZ
wkp/BeLgRV8SmAW/dnheP/sIf8igJ1ix1SlMs8un4+SvXSHZw1R8pYVuC3rZDm2D
yMfEs2GhkT5hgjsOi3pHOmy/xqR4wkggijEfvAe7eXajaYTxbdqlXMYRBNBQ32u9
dIKhQw+ExXi+vhjkT4ekrkYn2vlL690UAgJYl/w5yua5eYIhPXYpGJyUEWUolN8t
jzSKoilOPfQ3G2T1sCsBMZIkJcb3qeFL4n2n5ER3VEsPouEw8mACMy8sNG8hS9//
EcOYGtNiKVWKnPC3j3wehsdA/a41DOviAQ+a47OOCW/LXT+Bii8+cIYkXITYmBPu
kIDws5+RwcmNaL78tg6ot+reDb7LAHw4Zoa9iJps9uVu3pTmpiuiLuJB0LYevyg9
Y4nm+MtJIWTX/dOMvqa50MnsrjgFc/HbjFv2p/jTY/V4AGZDGCk5k0gwBjSV8NO0
FzC7VtcqITAgrVg0lELNHBcqL7IPzhhjqrISGBPvE2ZKjff5617+YC1KwL0VHkoV
Z5DqgIsXDRPzkWMWKHJqArypeDrSNGKr0Y3bmrwUhzg27tc7kxylCGqwnIU89Ffg
MtjKY/1j2QSPGwfuiNg7STG36ZTiVCToolaYwXnF0F0CsD3rdoSJmlyLp6yw5GSI
zHuD5pQPtZVS2MdvqSqwxS1o0WKTks4O0Feju40opA0ckm1Pk1Rl/uCaE0/WW/iS
jWBkFe3Df301Hxgdjs5SkKhoRk+ilGuwdqHKuBu7oCpWPxpDFO9111wJf+NJgo1i
sBluO3WqoFxOC1CVdoLDxsuXJptQ+HCM8wRGwwa7bF3Bz+1a/SM2qxZBg5WG8rxD
E6t39xeJOOPjo2zS1xgUIXZeuV9iCLT9rVDS5WB9TkLR2SfvZT+7HmBpoucA6uqj
XsmIDitrj5Lw3DpUFjunNaSQ3/2oncp21YNg61SiqomtzECvrAOEf0Pc/gfAHwOa
oK3riZA44J4jcu4Pch0/hcBVgxhk1zeXxRU7uziOIRVowRXTmHld6oTG+cjhF/ef
TAeHexWM/ChNkCFQvR2Tlb9dJ6qeLpW8n7az3ASKRYVc/hyyjlO7jfk5lcxcWMt2
qUrBXqz+k6iauGhLzEujX/05z4AkYvrlbkyT1ptyKHHO/luPYfkNyBJAbheiC2ez
25TrYlJBGx0Le5Icls3VgP4PNDpLPek1Ko1QWY1GBsC9Ta57hnfQqEFzzoVw4ZQf
hCNqxZ8fhXv5ZboeKK1UZdoRbWV2CXIsIaUBVtNXN4i4FFiu4LI/lQguMnAiMYZN
eVeDKF6025uwWff13rE9azzsS1lLh8eUCNCd7ivMDmLRHShh8CnK8JFs9O5GswDq
NsjGMHg1iUfhEArrdK9J7vnGCUWDVss1BIgdY3OyKrQn3R90FO4zaFmsADEW6lo6
Ip1yAXo0khzf/Pt7GYMk1E83AYNNJVLqxrDqnnA+k2f/lxGviPILWSRNtJuu9ydq
KiAxioZuIKqQ5XWGgRucKCpo17bqgojfEqX0wVt4mE35PXOePOY55jE/6Sr7HG98
qstewIVj/isx8UBwT+9m9MrMC6KdvuTraE6YHe69ZJeicbtymXGTB9UgMF7i1ANQ
E3wJVJdZImWRvFRknmcSHOoZfvx/IxWUVZQwL2ZfM9W12S7aW+CQpBDrRyMOOvaA
5vnhVozqWcpKB3iHTepnTkHXrOdza6ZrgB1XfPKOSsWEMKzykR4IHB5n9XNgJyVO
OBSUHVuyOOt3K8dwVcV84m/SLRQ5WWnvNRvh72t0mM1JnCWb+pb+fZECu4XrVy1Y
X/b8Jn/OjvftsSixVMTPbRpD2/TkKsFi16H+n6PwY5jfEB4UjRRvngKLhSlTgY92
KVB5bZqSpAeI4AQs4RiSN8IiIZhrsR46XcaMHwk9BODYvgQxzKmHr6L5tY6Hx0j7
BB/+9S0eaYi6BVYGspJIFaRf8GPOEBXfEsgxIubJOhgRVaEQUkne1hBc/7qdSJKr
zNnhsP1sP8RqPYy2zog58NnpdSd80ZIvMdfrRGB/XeaIKsehNt59aeBZWZfZpHGs
34tcPX04OV/yXkpkQi+JSYOqHiDYqAYG06xkN+y1pXX+5HGH4O9/Y4g9jddeaOyj
VzKeLcyjPLYfxatSrpRi8kMC8Qqo8tJGd3XM8h5YEj5jXLeNeHeVpBVYnKfZ128v
zEITMiZ2+s4fEjW2z2vaDMJMA8bciSnUnAR1C+NYx/MQhdF6kSl2G3f57BHRZqWK
47c0T7NDWDLzjD9kG4Dfkn4f3c2IZkluPhKymJf30/jUvsJTMIltO5zY1Mp6Pkfk
2ifC3uLfTYGYqcKF2WtJiSSymFVaZkCf9PVmn2Wx0eScqwvJTZYExDeREXTVnY0J
qD08EP9m2KoLPoe8fWTE6TrcCzcTV+7tumdf2nVetI/RJTyD7ZR9PJeaIqIh608j
VoCBR6ugBKcQ3lOwkk0n1J302lPq8oMDUOYiociXKfPYx5FA9wpWAtfKfJ4GBddM
ueWGMZDXZqUzGuo7pNqpFoIlEcsIPxwZSry9jQZRfitgS6LdfcLimMQucs4CJgWi
4PfRzGlpaXlm0aoYtdyWxxUDK7ffIUsesr2ZrAMhJZSo4l39Iec7dDUZjondykMt
PZZWb2YiCFDImvsGZp93zCpF5TY0JQ+d02YZZjwL9eGCZqai0akTedj+89pbg6aB
gbSVQZcWyhknatk0MjJ9te4sQWWq8OZ1PMoylXpkytxJHeH2u+KNZ3CF5KawaGBQ
++OowBLe4C6HrfmJXfuJKzBgRKRbAeB5600eByfb/4yELUvTpdM5bJTtDgzR8kV3
Rmp49w7BGK5SFJXz51LaBh9/buHjrl949nV3J/JV4hBoNJuM2dVd4gAEEPWi1Hx9
mztU38JZxIXw4TcY0Pepfa6Dh/1sBSIa1q70S0znJuBg5ge9634sIWEJj927IrvX
S8nWK5/fNoMlIkndQV5xEjQeuRfsSn4VdviHhtQzeUCHlJ/2VJwqEf7VeF7HIhJz
o6EZJGma2hcis9hWBG+/mcfn8R0x+h5GtQMOj/uo6O55Ytj6SPGZYbognzEkgNqw
GeNLuKFJnY95krU/ptfoy5KBl+DYE7UvoB4frFnyIoE33nsuWRfDWSolHK5O/a6K
wDz+5H8HLEmoULVD2paJxU/ENQ8HbklD+XehPEu4xqY+NtlOaJXxgNBVXoVcNj9D
XEqgrEU++QUwPJPN5aWgnBCwcXo3ivMgdlylaVYEUwoa/4927BwbY1aN5PPTYA1E
4ukam9E408wRINM63t3i9ZQZYfk0CJIndyi7uyzka7qtQdCECyNs92Hs+ejsLrhI
K6nXWaoOvf/OM7Uiq5x3CkFsbBT/w/UXiTRDokyq7m7ZmVgGpbcB1fOJuXEgVuku
olyBldnoEQqzrFehWLSRmvgLu7h5fscrXcYC090tY0zFI7hyeUDHdfjlRwu084uO
HAbU6BBuvDUzj3n0ne8j7PWaqtpUfUU8hVI9oDxnfYLpDUviV6pkQvZe31j9F39u
Hj6mULvZDQuA3liNRDPUbqFqNERkbCgdF2wLJYQALQUJhQMGUTdyMfhrbIpJdySy
tfnjZNNJsctwpLvSviot3YX41uoSnXQeSBZhEmyeDuRirCi+sGBMt9zGPtxgb7/d
J5Y83i+J6X+31sGtCPPVivVUs5p2rtIt57R8tha9MBiAXJVlPSMfbitwrYVv+ki3
5i3+oO1JjLkvX+zPjVZ46iPkGa8viX1dSoDSCAsv6SJjpRfbghNz1dHvO+DDqyI7
8pkCjMn+bbRHBBV7yTmcLw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GLNTGpO+lN5PUbOFTnLghzowqrrjGddW6W+Tj1Z3Fpc0xYvRaxQDR/XP9xy2UNrO
PFhnfGdTbiuCKtJaC/hzzoZrZjfDe/DtA3+myMJyZKMbTgjW0gBSZ4RVK90hMnbJ
n+NHqecPBldHV8Nw9TRgwk9n6sIZVuNFmRqQgAulUZ/3PaYXit824SqUQgAZdwWu
Sse97IgW1Nud0qYMavJ1TBIsTfI+j6ZfoylrFjSGBczoA0031Tp3Ek+puf9PXYm9
CYLichg7Caj2jYEIdZU0aMITpHZT29klFcL/8Binb+gWX7hbI8wOdANeNi+Hua8b
U/ics8g+3bSn9IkmxsxYoA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 23728 )
`pragma protect data_block
OWqArmsosdieLyHSLzmntbmP70lUrhk9dImpW+yXqCbbXHKf0wcBVdZSmlttB3Jf
GDMl9+bI+f2uISOAyRF1DwIYyhZluXwJ5fznd6A4tJtT0w37WcUO2RF1nz+q2Rsw
f3xbZPJ1y5dkpZaJiiqa5ygXlj/MktDT5KUgS7eIQuUiiRBAxDVWe3DggT7ErLaG
kN1y8Q6h3Y5WuV9dz/Asy/2tHf1yWUI0K1+rz4vzR87cbBJyV6NUdAvqVBipjMi/
5N8g1QGjpDSyqZnob0Kjua92zsGbwSgBb5cYmiou7m2cySKebSCjE1mwA35JMK4z
Fi9+UW90lhkIipYUVSHXO1p3ReLVaWWAVGPCfr82/NPC8zfJg+TiN98xUmXoXMg5
ajzf+PwqWFFMschoQCyXzwJZPJGVzoSIu49dmFPB4nHwfRH6kYOQgSsUig8yI+La
i9fPzmIJ1RPx322a6fjnROVYfP0SR52oZzrIkDGxcel9MqPtNIrj5W50S4B69w97
JwZZSwZcUIty9D8IpJlHeg9OxbV3VRPJXslXIfCokV8s9u/lrY5dEMxhRLrPQHEH
fROa9roeyyoWCfGEhkQhiIRn96MD07Eqfi6iAazxTSJV2jwlrSdCE7ld0PVPLtlB
V0ra98R8CMr9wHwPCPVsr6Fg4cLSq1y9c6AKMn2c3HTc/MSUnwDkO0awe1vgIgoU
LvQyYeE6EbORhIFPo7bzGmAQM1k2F9AnA+q+bNzLcH4nVP4a8pS1+jlew3yUS18O
LQ94FD68AwLdgqfgmgajtUfmbbTGnd9hLJC0cMQ1Jj6h7ZQzTtHlmt/IIBox82pv
ehDZ6El/4Aj7QpcLjDlAgvDGh5ME+jt8TAXxTT9/IGp5zqa+Hw9ZVWH/TM3GV48V
5Tv2AyQXBi7J9TfsZn4fJ67bHdGPE8ckAO0hOqvXHZt/5THCL819mHA840UJGJT/
8s4E5FKneVtV4OjJSMiPEai/oFjFvkpxnGTP+npnS03YBGNbR3lpHfa8FZeo2HDS
B4g+s4jI27Eq2Vs1YvlQafmQfexLd6K3qTaV1TRHmYd2FunK2y1eF4E4sg7gQVWD
KViJRNkQ93fJGAdxdLbYJI0hjAQKTXobP51EJgTOtHZ2X2CycVn6RPnhpyxklttW
sS4PnUc9dsh3l9evGh+NXlYQvjBvn0nqI5dtfmWy4sX5LCvg1VGCdNrVhSGSwvGv
NctLPf6vIR+2DNq2E0pda7rir67cP+H0uTUT2+19Ju12NErFeB0vbyngPa49o9MG
3e8/Owc1iqScDNuuWSndvZF12ojrTVKlujnbWZpY2Av9igZcBP7mvp/2NgmsRKyw
36otfL9XudNlUGlQBgkNrMdSCqlmES3IOWWXZWVnQpg/ozv3JMaQwdR+CIiHfDEY
TDbxC/Chi6doSI7L3eG5N2BzECY1PWDKiKdigrXGRbSlT3vI9kZcRSO8CpxKI991
kLpRCjObH+KQtOG07kXbsJUOCZLjLqZLqTpUYSB/Sug4FSmcn19ErNiaSZpvgyr1
UKwRk+yfSd2pheiuJBlEbX0M45f1TJ7Bmqsyz72+b2TybZAHIdcUMjSslwyedAhQ
4160t3Vxwj3YvbQO/GxhFbY9kT2sfwOUHQYCi/xm14WBAQKMnhcCQPEq06rNQ+6b
PkZhesB5fvZlY1656llIF1ilEe2tNLTnk6DMjPGn9XoNrWeyQL1A2bGS+leANoR3
aZwMHeF+J0SzTcSbVklwT3MCd2faaJez97T7GsO+avkWZ3zDwacYbNdd/L/7bSj1
APs/KsZUf/VSn/qds2hjvf+QFmr4yj9JBTRRQq3FfXoRj95VxdJErq1GdPqpuNKv
GBL8kj2LYf8R9HpdF00ZULUBjFAWe1/9RjUGW5udnM09ABmEaaYbxFEecKpOr+jj
hgHqldnQMx8P/Q53OC6oJKM02NMlVdc2KWNQsCYQrxg0MF/Zb8RkA5Pok6SL0AZ1
6eaTf/gdqFTm+zL5vvtW+VGCdEe7zozwA4zxzLA3DpT+tfRuKuGR/Qli20TCFP1G
7QmGxKi5MTUVkLhaT/lj1j6XowmE1y71xSMeZI1vLIAdTmlg8YQ+aGmo/G++FH9h
D/ZJKlem8GsDuWY8yPZKim6XOq3iKJtKbUQ3Zw8XptaxZSJNJyl1zDP8xxOBMnGe
q8dl6BS6ogpNUZqHEGrphCY9Cv7rJnzadZQF8RFzRIxQ/lBA/mwCSM65XbD6Pb7T
SBRBA+/BFjrPex3eNfJRb24u6tbFgPgvQutNQrla+pWef3Z69Fah05TXns+fQhTn
fSa7v58TCQai1aiDDvFkpKdxwgtcMC3sha8joEXoYSXdqt42bpA3HorLf4EMFXLy
rzB+SvzIN4BVvLPHiBesu/UjOEc2i3tNZWJZoI/89AwFPYnBy+cG+v5Dwqdm6NKO
XeK9XMTAAwuIs+my8RyBgb8619mOgjO3Y03oyIghVjXkNUMBDlbpDD7xO6IGUeC5
PITIhcGbsQpimOE/hL83GezDZ1EoTZzfgdNZoqq/M77aj2IlZ+0XcBdCReFVLV+x
T6VeZ2t+B5IrEAlGpfakm1XMWs0u/PQW9k0B2Nl7PKY5sFDBezrGb3njMqimJoOR
zYHfJgukh8s1WrBCfHCRE2O7XKVRbCXAmVXTg055aQFzVE8in9wJEAMsahGTWJYd
ToIWFzauNr31yghrVQz7Uqtq25lplFE1Bp8t1HxAbnDMh6D7RVywV99MvITLyDfV
nteHya4pQ+SPBmsSdLu1pNj7fOwG+UshKn5yLI7RnLcEjamSwpWn68wfGLwxlACG
zy4e562NLnar8/vLWdyQkK0wfc8D3s0/f9zA8fwpM2jvNJGy/XcoAlRmOZSJCqEL
wm345FCn52g9PAAD7I8sxLdpyHTGpG1mws7py/CLvlw3r4sEq4c0FlDN69IVNMEo
13DkuQ0ABQ2QGHJWeFFkm6RTKAbJLQ3zyay6r1cKlC0y8P84/VjwvUWzICYPQHfI
u7Mi08UTvJsEm6iOEGzEKaMbrtKtz8nlG6Eg1R0tV4ymZSo5R0myAqOu/swZS80P
6zJboSV2BgfBuAb5HgEdz3TwmbHwOoJD7T3jnW2YPpB7YnTftlsSBj0JsFMBsaJ8
8fM8ZWWhOo3MExmEDD4ynxEq5DZUjfVSp0sBybmEVmX3cdZqjIpWJb5JO3HguGLV
8hPgbGDTrg7DK/RcOxb/i4EUhfur8epi55wJiG1axWLWanj3WxZ/zTih3MTj2cUu
wB7gYCZ3/JgVWjgr50VszPM9JkDvA3hSNqIKO9ooKQNUxfvdeZufV+jvwP3sZbU7
zXcVpJqDXc+U0bkNIwelyRmDBk5m9uIItX9dk/MPpWeje45MCbFDSzicgrna415X
fvn9Tna2tnyxmlb79tclubSY8O51lDHiNP1xzg6zhCJa7QZwEMs1QbrxpWjwsXmc
vyduD5G7TxcaAz/q5nxFGRy+u7UmL83D3cGJjPfwjg0e87TM8UYNdOMXdq2Hvvn4
5pcUDugFCzMrFzuca3o+c+31avfkp0mTtUs8tg2aYMFiChK8QVB3AnLSqQJzjfDq
vhJN7BCA0j/7PPsLy5OicNIStk6/kt/EHtx3ChxZ+d9wxXch+fycGBz4symjBfvL
Fu4lvxuVFeiUcXYHUIGHPRYmh4c0uyZkhCJh9tb3GgvRxyeQbT7+m4i8oNor507Q
lfOyUEVmqt08OhthBDZBcLQ6yl+TYDhHnHzIfjH/iYe2SiFBWqMRquYHe4Ankwvk
VcFYe+Z0L18Bfd2q5hVAwQQf344at3TO3hBkHhWbZjckRe/6A6kFkJc+FSzq3IJv
aXw2H/ZErihpFI2v7sAJFh8vPB3/yUPJTQAP9GgivVWXesuVYJH6VxIhLLwuMvBn
buuIhKrd8IeSvYa/42fKgqDljr8OXS0S/ILABtJ9v9r2SEQAak/tQV/FrzPEe6eM
pD78iGSf5ww5HFEaxIWjDSDjdRVk7H8rNmf/TeNyWjalYajooL0RM++0zolFYOmE
gm13A65ogwn+72PwGwtmhGkaXPaDcWN+h2PS6ej5iZZ9pFELP9/5yvyj9X0VtTNC
Y5m4Ex/Dm9FPYrPORIt0Z7/FURdDut9D8xVkN+oDcyPgHlFEwWeNy4XB2gZXUXvC
b5JF2EXo5wJunS6QtnrfiuMVkljoZfP54l5DB+y3wI4Zfi0uL2YLpuEzmi3jHhm2
Vzl8I49tdyqfNFEAWVS02pFg8TRcAVxqYXuLVz3hOUfsdITFqKevj3RgDtRjr/HU
VtaGDxgTLhrjrbtTFmffjpmujzoV8q/4iIpfcHvSFN8HmgkyGEkEichx52SxxvvH
VcKAcCJK+X2BVks26E9vMRBaTxcXSFZ5e8MKiR9m2DC382TQ0FkgtGgo0U1NNPsk
oHld98bYouAdDc29xwXnyxkTuT17/UPRfSyASt6kgK6QS76Lu9TNTDDoAIu2K2j3
el/NWbXIwx1HJ/3k7NPiKXK08wIwWRQWxFjfh+aQUkojez4ZDk59yESRLb4ZfDmD
Nrl9ApcDpPGmpL6g1SHsMf/dUqePRsQgyUv8XCfHAe6INg2qxA+kFzR/fBBrEWmd
ucn41SNaufLbnSzU3xAN0TLN/LPw69Ov+lz3EK4zjCKzDyengcOAjXrF5rVGAK6l
uvQxMZhJgPSkxHbLhhNIePkf3/6jRgT+AD9BulaiXtfK9HTaY3CDRoO8WMADlbnD
WWQrqs6LBz4WZgqUkcrpWMnX6x42VtFpcPtodzId7HxS7T9sjhNbh2aVs/BuWsxQ
Nlh68njpHGbiZz5gz3Rl55v2+QxOkQJQURjRfp1hVjC1RsUTi/cUMoX1o+dpYoLT
XWrZzEZ8MY5TqNJsmX9X2++CzqRFTAKCj0udx/YfUnGG7+wTgk1sZ5jUU6u6YJa8
qWkO3CysQPkEByxKb3PNvS9diElHzMev3/yfOjn1+wAt/lBbtc1a/Ts6ivTDELgR
XtiJd5u3CVjiwjOpvbA4bbm+cpbeFk5H+JCssnHsDBd4G7SE8ZjdC4Nfk3ndpeyG
aMpFZ+ZSFMTJYNTNTl/ZG36pnYM1WMYu36OspJpp+thEGuXbojK2mc7axp95Yx8o
LEB4ShZj06y1V6nTsz/ySXV3Sh/mWPY29JxJknuA3Wz5NQ/z7TCp/Ucble/UUTl8
9kXxgUEynmsSPyqtETEZSGEHTgFWZJ0zSZETBTqe+ulAl9UNEjV7g0wwBPD7iVtS
Ogo6bMEUumnuuVjj1H2Z85VBQu7LSZm8e0OAaMXjtea46pWjMGobgjizA7f80JpA
7kjqK5Y9SEsKTQw/ST9EvmSyp99gX7v/X27Kd+P+X6aMXExnCsG76iZylMharDsq
6xG8S3XyM3J17X6ZNfeyEi4BmaGSZQdRvl85tn62bNFM/cu8g51MCLvUlOD+AaC1
psDz+HOF4esA/tGzbcxoX4wOsVwREdLIWxhWltWH/Swu61tt0jPPXoO4BiiC+cK4
8d2sh1xW8LSZdX8RJBXXyzFvIBN9sUiKU26gBeOgiZ97UDwb3TaZ+hKc4XWFxWt9
N5FQj1n8RmJ2NmKPNRo3Xcq7UC87Rs8MRA3PtR02cpBAwiaF+zZuMRSehLxAUryS
QZXZYRJ1uzqZxgOv4ZvKPsxAHxLhi0DHEUe80fpgdUEfnm7rmTRx35SKM8nqLbMO
NxybfJ3hGCy/ES1mPRI94CsdGQ4SNZGkCCBzAcTW26/ojLndbsu4SFk5abUpQRf7
LGb3krMU/E44cNzOexQQ5zdjY8DRpsAwssEEpPG3/XGDJNSUH6yDzOfBX0d2TbdA
OJfLsDyKVwzrvAM3ZrSgK91nwEdvI2IRnMU2iCC7w389W1lqf3DxcKb3BxLNfD/s
e1sZXP84bhsvyLmmu1MUgQdn0rm2poTFhkBiDKpnF976k10rJaeE092xt5D3eYWo
8RwZEry9FesEKAd8mWy3rlMtdP+sQ6jaVe1olcafqLEhXD95H6CjSGuOHPzxOgFI
OV6nxGUdVfeKB6ERavEBlRq6k0DYS22u2uBlp6NKZJq0l+Xb97zg5ftwURAPQ3zN
OeH/+xyinbcTEIlt2/RcPTBYNE4IwEkJEEE4vJhOcYoX5YQR5Stliq46JF/33HKx
k8OjJcEmwMqxyrMRAxDC10LO8yjN8RRWQfy5IWxOTXA1AZXgStm6kMvpiw1RT5S3
/ux/jZgqtmw5+cOnOiJZ1Acs6p9C0sguHcie2AN9GaHovU1MBYr0yJr+4ku4pxwP
iJVR+7Ex3rJ5SLxv5grtxo5Fjk/tpOoh9CDs3UBEqz7pf0I5y4jZWSFd//wYaOx7
MtO2hap3vwEP/uT6/rJ1tA026SRTBjPup5qVywg00tYcHa/O8V5c26NzA14nEFqc
1xdh4+MZotf0zFPHNZNTwJ9uTW5L8inP4WKdf3w747Ft4/ds3Dxf50VaqtrlxRrz
KIY1M8b2KnLbzUaD9GGS3TGtUr6KOS2BKrYCwOJrCEhtlZZ4CEn94+EdK3TeCrYt
1c+FPeEV+VtzJt/vPLbAbO6Q3Fg4YKOxLWoIatOhe5o098EFoXp444tjeLXJK7Li
dJoHNUAixzDExg1rkfhEiQOSjs018PUSpH+Rw2g0FLZwwNduG3EI4XHM7sj77Lto
vlGHSnR7rK1ySrtT37VJpZh97C/MPBHYhJHqLpr7t37ihweHY6PNWuVvGtzNKMh6
SVlpGyD1RREkzuertIZX8yDc9jdAVrDFDJeFPyqnbEhNe1RNh3v2Va6uP1JXQXHH
zWtcxvJC5JOi/4+Igh/+582kKiWMYU0Dl77oMz4U47wbw56zk1wRFB6WBfHWMfZA
9bepMt83lGWXIPkeJ1NjN8l1XFn+weB8dKrKvMQAclw/ef6AfxR46C+K2JmeIBQk
7jcQxuS/0fgO1ByRl1sbWKuOEMVL4sIdEdmrqBIRSbzIOBMEh+cbV6O43wSFH6dY
awydl5f5AH0dm3Ndy5K+PtcTjjF4w+e2lSS7BX1t02cKa7gkzg8D9xTEkqadX4Kn
lXWK80uLi23F29+Lfm49GVTHA8gRfDYlow8xqzR5o19/1pi5ocKdhG5xAuqOfVAh
LQcdxTu/oXOS+YNx/Vies/AO3/sUdiMTatE4yooVj+9dAxzpuw+DD6fpvjFgXMta
QGdirLv8kTRc102lx4ROM0gJWeFxOZynxcZzcnRsnMz8o2YDjDFv4gmKI6euMTI5
iFG56E699VYW1mA5A8PrU6HVZSc6rjgBc1mR4slOh8I/UFfaBMKtyz3oWUnUZlm2
M6RGjMe2hHcL271vvleW5biAaaSFt/78p2lJU3K8Yww7eYZ/QkztvgIUkph5Qx4A
XFRDyS6vIQVIO16E1zGC7/+c+3R5doAuRVWgA9wSjlsFWWUrzJcZ2MA46ODOROeG
zPShv04Wylp1LHYJxymuqWEN1ybWxNLZTDqib235TIhkL05nhIGRgVQH9+hnGzkb
TaMaglv96xjHTeGHLuo67t3sPw67ycvG7K/784kju45xUcmRJOlYeI8jRM40pL3e
4ouvXT/yh+MSpibXMF/+Xtdhz8RZDc/PNg/8ZvPC2m6Vqf9Mq6TTO/M4JNuJW9MC
NbCEV2cgEgXo13vsoWXQU/CVUPsx77QXu8eJx6AzU066VlZMkH9eWvzOv0Y0amOe
JHi6GujkeILwqgY9j2vgs4zZasWqUPYiz3kSIQFCb9H0+dmvQ/F16mqOUjXerkYr
+J6KdaJzTgM+oS5vRDvg5lVeGuW2v1SJDjMNOoFy/KRk1Z1h1jgr61T3tt9lxcyn
T4YiH4wnwjhO+9s4P+1KQaw8iMU0BKzC7fibxRDdhAEejk8+Yh++6k1EaWfZo7w9
CRWRFA2oVhH+41SYnRyC9fFVtJRzRmntyXEj8EiE5Aq0iQ8dSoIK3UZfrwJJW3m0
ZsimOMnoaxX9tLZLN8G/hs7sTwUEnGzGgimjFq2BULtkH88PodQJ2fKhRhIczIsT
du2IN+yhpO2GrjPZr5mIRMfysiMMDCGaa30ErDCXuQWOUULpLVAWW8hYKZFWJbCg
OUMcNtVfKul4OIFC2pW4aRgH7XKsc5ZZ+MDNV/ODupgClTLpHjVWSBsjsx7mpuUw
iJ0BFC5hXojHzZcMl9M1yoAberfMS9qiOXV3vQ0ccEsfhxdvKtkSEN+iQfKWeWWq
mlOGg/ZZ7PhmKy13Cs+PhBbXw7jivX/b7v5gIOR5BVTGTsCEja9MrGWY6NWsauJD
OLTIN91uL33aZLM3v8NPiZhNqZDSE6CnsyxegXOxkXz5XnU9LkpXJgTVHO1F1HQl
811i0Hs2tXVCFEeM3o7RXn+g31+KGGtiEtlq64mM+qR4Pl6KeA/yP4JaTkTTGTJQ
N7n40dr4JFVdlcLse8HVSaeGthmygktTrRtefowQ+MCJHirYGNNq+/RoOlYPJJBQ
ZqpR+Ae0GeXmCexc7T97rF8DPJomvikEKMruPXdX0YgmMXT1xxiqfMHULlYKYziS
vGM55Gt1QWQC6I1CCaYsv+i20j1m9pSXLeGGi1YXHr3jOPRDzoUlUC4eWjY1MQe0
TSEZaiROMFFhhbzhMQaCY2QZKQjvBHdeJErRpIeLT7oHU9GjH2HnOCTEqJUUpLCM
9TBff/dvAwDq5xB/aeq6IGtI4goZL4Ian5GewPlpX6URKiROFRBoPozyswpMxs1d
e1X2m73WK7am9uoc/ceSwKAL4BqHrjAMCDXbZi/flhedGIL8YP2c1b0uzdespxwX
ktijVDTFXVPopKS41nOD8sUTynUPHwdT20jjKnQsDF6QX93S427WBysz7DNaGI61
UbI1iluswBZXzvYMuRkuyEj+oO0EAnydK6YxLxIrIhHVkT6dlVZTnWvqHFEMtNw/
1cGygPYYXsi76VNY0QbJz/HF1kpZKSa9jrDua3agTzafzdGvkiJVky4dF2wPU4cQ
JwbYBc10hNfCTZV0mPIlJtPsHMmiyiRO4BQ3Rzrf798ZOAAmhqsIsea9EPGwcaPb
i9BZ0Am6lJHt5ZlTWcf8wLGxlj1hmsMCTBnie6OkQlvqX/t2EK+XJ6lQb1opPK6E
iV+9oZQ/4SPgNkJPAdj8dTAdtMn/urPKUCgNDU3hSvJ36Un9KZLUuUkvw3zG7tz4
P/WQhfnQIWtuTOGoTd2FDctpJi8zSyQieGB2nX/xfNCcelScKQfxFu4VnVh3mlJg
WTENLOjoqICLV/7sji5E8xth4IAUPTqYoRRjlCOAAToVEqRUve3IuUYtc7c4CMfZ
pJbdSV4GGqN6p5yMOX1yXDYExg6UNxlJJJiuY4RxC/qgS3yA90yeyKgzgOokQuLt
dB+jqXapDrMUDPkxkx+3+zH8xGT9xOTbbu7JJXcaFGQ4EKblgsFaNVWE9IDVaI1L
sBsbHN5cWaFzoVhNQi9v1XrSwhdOAYjz1jLKn9A+HKt7WfngMMGtd/vZV+LvC/G/
1Oo2fp0UD+RI7SW6cw6pZ585r91sNrz80DleEETBdxDOqZ1xvk7nbQIlDny1Xx4E
c9cCxsHHgbNuogWUU0meBYpOHRBHHMwd3aAe2IXo9KQ1WVzw+R+nce4e98JZrOPQ
z2yqREgQAmYo9urlXpIGDei9qq5bLLflCG/pkaRCOd6zJT4zZ39DESy1zEVCfhI1
Jyo8pqFyAfMy1m5+FtBNum0YeM+fRdX8pmKksm53JD7NqbPcKCb66/jap6ATX8Lw
z6uQL6rUySsCF+PF5lRMi+uysPOoEDjqitOpqCl962QVYnLtKuXh7gvHTpEU+qc8
l0rDeF7iLAUV3HF67O21DfE/AlWgSwmaPDZi/cAWydc84J3k5q+PqQie4PTgtR/1
MtOx9s8BFBZZoGm4nDPWh1UcUEjhLZByubjoJ71FdrW76qy/jtTeXmoa4EJ/fyrT
ks9WkNkbkozcqJdc1LmzNr2O7H5pZz+DetNQ4uhnRHJQ/DlvRJHUEA94NndW22tK
QasEBtSW83uguTzsQFK0E+davXZ5trgs84IC6+UAl2bfQLY1IM1oRIGuC7+h38no
kDtcsrErM+YkZirMTBQCl481ZE3oO0vzjnt0KkBAWDLkCzJL4rDiVurVjtECD/sE
77GqXzaxn228syXg1j7JrZDD16fymQKRIpaAVkuhac8i5VlHJveONEqpZ+u3VF45
ND0kIuU4W3BO9UIEur0P81vl1iDb97b65iRbegmPW0cZFo2i7blEf4DAA9fqz1Yt
VGpwTEo1th2MXvJBhDxmxLfBL7AeMSxx89+eNm5E5sRMp68WstfskGLJsRwSOumW
C5pdpFqw17O1sihcIIixJ9RE7Q7NPIIgQDLsRWgR12+s2RpBSKLVYXjgeTgVHcBH
9CdcI2Jr9LFYiWPryWZGQlkvumrUsJZnWCVqtq5ReyG3n+v5AI+yMgOaNEMmrOzj
QTlfJZPCrs3YWbgQmLMMoEf4gSSZP9GW+vyil4tpROAzKGRgVcM+hE6qfqtrWhfQ
P4otR9roz67jMOatLZOCcS1nnOXqsN0aW4y3ai2yPS3HXq4dSQun5Z1n92+lPGaw
RXNJJzioxEPJS3ny+BbVic2YqoadI6wxX6P2TIvvo9t+B27U8Q2fgRgOpN8gJ148
3KG5KM0o2or6oZhBDKlmQLLMPCr2lZUnTMw6rgUD8BB9VXGt2MdE58fJ8sUs16Av
X6OWpHu3JAfnrR4RhFnH62Q/Pt/MBGOy7ERAA/qcoZFS85sgXlhuwjFi9hWDN3HQ
PINHhGj9fykr4gJVqD3TARKr4sm+o/u3EfvAFXrvKDoIcueOJQgOZ7nIctNrcbaG
984SEkB5A3yQuM1+ig/UR21dN8Yq1RUYljSD2gJxZwKV0KuKTMtDu/BAB6bDjZv0
WPdrIBMzRjf7yznaJM3epgwsswBvvHoe3KsbNyMlykEXKJbyLsxhgJUgbFjGxWq6
s//WJFViSIsdPuXvl215G5ovI+cTh90XHiz03d7Hju++qS9Bz9cwoN6OqLazhfUl
aQzgAq9/wuT50pJdoVNX8w24rpDGPF6b3qSYERtMbfhwgbaYeuuW4GaowOF9gGR7
KCc1I6gnjZi48uKlIzbMFvnzr8Tdk7LssBNEFXfxjHnedTMhkTrX2GpCfbejg3xh
Bj+TkSdSPpQ4oxxwb7jO1vzq066beKViIJM/dxqWIkyKuKbk12baCYaMKeQGtJqs
DMMlNuEJQo3pW+nWICyqt3cGmLt4D96CvcKP7/xgbjwYPkngpoFcBDFB/hY50fFV
1Fhzj/ZPeOKMAVB6b/HtFkkvd8xEVaz9UrJiFESzIFZ5dc1XtY8CRP3eRgjnJtxc
/r2f3hGBOSVMSeFO3RKPWPJm0g3SUilxU7v93qNauBwDy5tJ+drSc9e+J+0vHQ1e
1iiVNSvFxyw4O3D3VOGnnTuBonN1gqJhW15MvBu+kCSE1dAUy0Ygkt0vrzeotIvi
56z69660Qd4y/escEj7vcbTgbKyw1+OXZlz73NiIBuhROORXMvX5/2ys6j6EGiVJ
I7QQVHkl+yX06AiWevugYZMSqW97txjuLzikcPvWEXnTyqJya1OStpvF4F63WIx0
ryPCnMoCMdufSfP4DAMB1e3S4FEaFAiRQSgYRNyGlfBZEn5s+OcFoWkP1NST9jvh
6msoX0Su7nQppU6yIVuddRQSOfpbK6A6nPRiRdzUVsKDGISIuj/Ct2kG7/fqIhLd
VntBmcYLvfP8OIBS5Y+KlauPH2Fgt2Z8ziFDPkUzzqoTNK4pCQtgws8H5EdqP71t
Z5toOBtUFcTRsCwwlKyuJMDCKeqqUMY0aaRGe0pxe4qRF952D8rdXJdpSonxHOlw
qnCj/AbewQJmEgPS6bky/RGBYTplQNQ0VUdBFmrpyvlZ+E1NGHoMja1B6ImLYS47
D7iUWyBD6N9Jiq7dLCfb8G0L4OxyknvE7pwzu2hfUycFkZCZr4nhVzAwUfZX3VGi
x9c/2ECiMTxkzZM/BqbT7oQIb0LA0kmh5HciijdGKka4Z+k9RbkSgJNlBbv4v2Ds
DJwMaQxcxtT4OE4nsZLNQc2Uv6EvVMjP2yhGwBJkIt8nNYhf8zVDKxlMsOaTy2i4
AbwOpNRv2xxPFw38MyWjSeNj2Rd+zAYnjC9x+SIDxv9U9nS01mKUu62J60Qt/rDq
nwJJSm/jP1v65Y0QheLMWFNMmGydYPHFW+MbLFqZg7rtI/m1OzW3hqcV5v6N5kMp
QkfQRs+NYySd7yBVcKR27hQ8TI1hzUl1EMkrxnWfLVAn+vXwJAZRK3ytWFx8lxb8
8aPD85+QGXDCkzGaXlzb+cRbInrZiue6N5DYiyZX1dy4r5ssDbt08VwibUgIcMKF
XnvUTYEE/kEzOuxGPQPE81QuMGsd5bgRwA7VlgxtLWH9sXoYYYYTli1Aez88S5ZN
+5RhH0PKduN5d5esdGn5jPGnOHmnkv4kTqM6fn13QAMTjMicubuDPz0PWUXlRbW4
Z9SomLE2BI7QDoeP1vN7im2+TQcedyvWqaT+/yUjOOSP4s6filGdftSmswNnqrVH
T3JcwhoThVXXlxryBYqTuSN54BddjQjuWp2Uc6YNu26QVeE9mTCpSR43p3rjaRo3
+aiAbJq7jrZzeqRCzZCcOTm4q/d7o2KxjcBgXNKQTWaWgPhQ9Mc9D8h0SaXU+jEs
lQyeh+xRZPJ30Yw48ulmT8u00or2uHnPNwHPAc0jtF8aB2Drqh3PeJF9aT9P8iZ9
r2BPSQRAKdmrTdm4KAZ8BIOMUml4o3LRx1OqXVIfzcQQ6nwe73UbSzzYNWb0PKFU
KxTHQB2U10oRLji8SWTnQgQJTpSRivsvkb//KdVmZvLRj0SLzWsmVNSTLY01ApNO
3i5WdCMiEEvr+fcNooG67ywEiMKo4MghgsWWjHlFvQ5l3nle0nlv2mRykBdxmOBy
kr4DdJOslIAw5ql6JnuRmuGlQO+I4VriTkLykUep/7ACOsRlHxf65q4UvRRnc3ba
s9MbuemcJHU3tax7bQF/sRAF6y6NeIfwW30ZXxhGgRTMoaH0TJ4JbetcXliExyG5
0vZpk4mBVNVSiGmphpmX/nYkOqekXvL7s6ZgsImj0SAvC4MRVHRtosnkl2vfUumL
N+25zebzYyMCQom+PDfEAbMNhrsFnIRntf8aMwNVzlULeEx8xsJJNINHJ27Kk/7n
6GqgMmbGiIMYmqwbiupAJA00ufUAWAPkDz1g5WcZ3298z5keioVmu12UcT16BGnf
wnXqmrHdpRt4d5SXC9omQ6twMkzXINODy0tJw8RQCrCXLuxAsAqJK8QQ83Jj9jzl
ArsGweWE1HiYduGSd7GIQ+RtCoNxezjHujbhCdNWnEG58Am2oRiIwmfouQe3aBPT
+QmQTwsd08HRUJro86zXgGsx0IiKW9vrMMTBu7oZr24+P+k2r8/XW6oMM65tyo5m
5nuOH2ryx0FcG/ZxhBLLZBQGT1L7rpsyIkDB2mLKGS562CRfIgZOOqhmeTR2RC+I
zA+Qzn1mEN2oJCtGdIjCvYQQ0dCaVAJSVQzhBAaSsqo80/hr+zx6F8/gxciO2jkJ
GKdUEqMLNsB5+9lIQ8Pmr+Zdp8m/Xxt+x8iX6eBzvmgTRES9vT1+Mf0wHtEuSVYQ
l0QjD2LF8g6wVRgk/vun/1qTN/wHprqUJ3hCuNUbSoXhRrubhbXsqIL4NpMWAqxq
dcbfBAmv60oHshlyuLjhVWnRtT20cCMtKNOvw7sOpFl5UZ9Dj5fqP/K09DlQJXED
/GznoVxkOxYMvVqIVNjlgmdM9fgmbDv9PDtmnUSlaGc45ujSSMF0FqmESHBOZrBz
UGsZqixm4TWNpjtHHECRxNZzA3iaqE+YG+4Xxv/KTVlYx+0Wedr7s1MfmmZuuzpD
lBNUi/bYLy5k5RQoe/mLjwkhlkVAdwnOS1QzqKvub73M82BsJTbP0lEBo+XJDufW
BcPEGtLvQVEVKKIjraK7A/6ZJt+i3Pp1++Y26e1tA/IEp+Opg0/iSIJ3XUDUU308
PM4W4yg5tHX4nhp+403G02KqHdui+mS7edSDxdPeSxKLoHEow2RD2/eK5Yj7Nt6t
TeZ0yEp6DTnHVcCK/pB8VZ3TgjbE/hUoGALRjqE1UU27vDZnan/AfYTKCSNsaHOh
87Pfp2/lcTUC+8ZJSGh9A6e3Yi0vC50GkaW7jJfGUOSOsBUF7pEDl0S0mDu9Wi2k
rztOOdVewJu8WPpwXeaEeiQO00YowbdzadOK3h+LsNu0gRxv9fOdjPdzHEEoTWvo
JNmkOepzNhommjbDq3K2AHDsu13klfo2wsHy/wM98jrxMf2px5UiQSk63ZNu/fK9
i4VXRtZP7AOZA/RBsp45iPwcvctWhXwfBF8GqQ1itjp7w7cJpqCnZuIB/3fvIcb2
tY7ANsKbqxKQZhzd7oHX79UeBFhHsJONa1UzCEKy2a7gzU4zdNcN/s8rbYep3oBv
1gow/e1zmZs8CFAOvrOpNa2PuXxFRWTrjjXjKSW+HDoZqG2ccwTKjXEDdDchwKGd
kyyltIBz3SXojz0lpxOZV4BLm7+VXV+/udHugHJOgXAPOTRBgGmIexnITtiEuhDa
s2zRFt5i34fCcevwRxvEupccGONaiMMOVRW4zAsIls81No9qcb36ISmRqaGDOWQy
PkhTmW3OqyI3hDkNhRMI5JVo8DZxmX1VEfsw8jQIu5rDC97NLmwCod+jQH7gh8G+
oO2GkJ3XQmQIMzKnaS7J5t6e6TmJ5spu3zBQDpEr9K7pnZ/L/PY5JNrHhLbSd1Xj
U1r7YRq8PQrL4FJdpncqzjBKVhyweYgf+OjUqQ/xkt8nRnv9lPfEDeA1w0BjtTgL
CX9jmTZmdCtbxGaBQPXe4BIA+1AvJI+9UmwySJTAg7HBRJTFl3DpVWu+p4sSCd+J
bxmsxNJvEnjmMgek71QqI3HxQOfGBij4+lLpIY0EIwHHUiGh6mD+VcUOWtdRrgZf
V0/j15o8GDnrQfGX3qezYL1vCpPK/mRjucSUNjD49aE/vSbIY7RV8+JQZOeKNoiH
yjasFnOso4j2lzOPj7FA9yb4Y8jJ0SNY4DwQTn3//sIkPhf7+aB2PERefWZ7Lq/N
/OXdjEsSAsmqXVAlX09x+rMQZrHse0/GRtWHFfPgprXXVWJGzZ6V/hdLHdAeTcdK
ENS4An5Ikj9LLeU42oRzQoUgfkeIzwSZ9HXkCeuUHHBCX0QIg3QtP+peEs9TQGd1
t1lBU9JPXSW4SoR8qefkg6clQhWIHtqlRn0oR8WnhhmeA5EDQsPePGHfF9WqYVBn
UKy5Wk0BTLGQj/r9MrZIqVgX1/xv5+lOAmf4lTYT5k96Q/zEOk8bx/r4w6ieK9Xf
VaEtYgWvf6JdFAAOgUdJnmJYJRhLcIF75jcGiWrtP/ux7xx/zilqx0Lu5pZfIqRH
b9lUQQ2EKRLb1AZLU/bFyvgwIvmSOe0EUdMAuQKW6hCsRfPou0xn+IWPzm+gan73
AbLMi/b8A2B5G18RMkGHHTAyTBCA+67o5HyglI2Ck5JleM5zGLtiHW/kMV9LqUsl
rXVuWbS96Em+lGymEbaTl+UBv/JS873pT3/PQPPFUPJnujjchviAhw72ee+lPVTv
NYToWUrqqrAVP557iYx1Pwa8EqqzJbj3CUE18q0s5U2sRLBAcxlrPVGAnoTcR/bE
oVk0CjdgRwp7gvM+nbOIJkbxEn1yFFlrVFS0k3STTXeUYejdwrcBSbDlJBh6CNZT
zJN3VS2450/FaVKWhxAErdJdBa4vg+kzHO6lA0Y/ZvuWDGncJbS9UmWvGP75mEwr
DqT1vqNCon1K5MBEeU3I7yYpobjbzbNB8JrqxGDuajIbni17pev4UyQISewDMQV/
xZsRsHRjBzxdNX/M+4DgVvrANzHUfx+S4Yn11HR42s5BV2C7CcAoMlOt+GAoAe8M
+GfYS60U2Z7i47g/jkQIhvqBSsJWAJg/o0+yfP/2QDD35nVk/3TKMbib+dHsxcSl
1gTzfm2B1MBGPgrBMZbIcucTU9agI/9gNzbs/rdEAPvOIVIlqylCWjfQFa4SXfQx
5VvozPjp8FIL3qhZVMqm2W/+4vX2pfc161W6Dq+oA79pD3PXPL/MzPQfX05JDeiM
SJCga6zig04xvxxzQc5DomVBIvQ5aRpsxqnkEFUnrPdxxTQovw1LS3jp6/75sCyc
29XNJpMQmkfGKieVNbQCDoQzpIEWndjnDLIegrtqUpHCDAsMmAiFOEkDYg2rXadA
wJClIh0UwfIIfDVsqO+aAWpa8JZYsaoXMplgEg8Oa+ppL/QTX0RJh+cwtbcl95jK
KDmM7Jrlh7hMwExG+amyI1ECAoGiWFIh6O1ZO4kvAzOQek5L2RkmUIMgNuzhYqFP
Rk/hs8NCh2m2/byMJsdamRqdkygk9EVKAQ2s++9K0cegrV6WVL9WSjRDr+xpn7Na
7nFunaGY/BWViJXWy4U/4vNzvUVkyoddlHZE/MiJo1y8IaUJ6kqUbThYPFqrpHH0
n0w+VpvVE0J8pkDGoB+wJJEObXq5I5Upe8o10zfTTvtFdjzDbt6F6fFVDCGeLG5b
jZW/hIxrsJGDZe6aWm9FnsB/L2ep3VUrpugLq2DZTByolJxOqx3IX8fbp/iB5Yrf
bjL15AqmSxtMeamMZy09sROh6v9etQiR8Qiugcy+ehWPIpO+Pl73O9fWw8pUQGSS
Fy+GczJDJcJT+9WL5Q1WZdF7oHsqYa/JwTg8cNsliOp2gRHgBRKoDBhFsMSf3o93
1mb/rCvkI8Cy4LDqdO2bxyN9MHVq5A7pu8eJIyyu0gczvm9dC3M70DFQceJY1S2l
RcmCFJicfYi9KWkC2InYfJOjGHkJ+Jk4h/eZDWIIv5c4YEzOcWAG5SytXYpjWozZ
LJGFD9BdHSezN+mQakrVKJm4BhjlkTXD1p3ufydIxigVIk9btLL6Dl8WYS/g1+SB
6fAWqsV+NN2Chtlz1Bq92cTw/40LsS2ngPxk/Z4H3Iqld5ozc9Olll/3fJ+An2Y6
KlJoTNr/j5MP6u7AgdjOttcJSOf3bx2E7fOAtrLp4IHFgfw7gzVeF4TMtHQT2iD1
FgqL/xW8lcGuAJvFg2z+zN5+iRgkSOvkR9TQal481vL083HXpREoLgCkcxRIHV5k
TL3NGTE8PUjBShJKMt6dWNlevjqn8yBlZzI72tIcB/V8iwTtlgvOXkgXs/niRlG2
CGmUNd9uolD1hEQD8qTDOyV+yqFRPpQbNbvuFba/VUt3NzHy3B0DKlJ8CM6vguu2
GnHwlfJJ0Yx12FMCrTjcJMXtyn3iUqJwshPoTiPonYoZvAyeAqnl8bCCzQWiTQRR
LwMuRtgAG47Q6CmoaV+l2pSyWusaQWSlI/30sXbg+JGUXQfZRlWhP4DxOCealPSD
kEudr3Sd1WJXhSNNiZYS4XBruFx4yNkAHx5t2u5rMnmGQr0PnIWLCv7jWbgPlFmg
eE44lsA4NkvbNx8iCrRL3VNzG8w15VCn9zJZso7L8+33uOTf6h/FJa5LnMFjDkds
1wt4zC8jtTUMfgw2GLFAYkCRKdORis2snWgwZQDv+WWmaRDE2qcLzuCzl/d2YBug
fzoSPX3D7XtQreXVor3tRK7YWRjHRLsiNL/mh6s93TEXX63S8EyAxvK0lTPEKjpL
SGhO4/HrtLPHwZYWXAFgDEESYuAgBd1Pr962lnvshVSyHj9Ahz9Zq+KtP7Lpsmv7
8fRj3ayN+6Fby9Q5V2Kf3xee69c8QFUj3kYEiformXt0iMjDtBnGdRs9uRKnQ5/a
yKiDPY+5bbuwMb5zsJGee2Z0LyOde6CFOqAZ3K3DixoPfiqCrXSGnbGbYDtf7KN5
jiCQwzsdJXliiGTaCH2XyKa2lOsQMJJivneHoHSveMPLAD6UzZFC3OGCSnRVNqfo
KCzWovVPPZagCeN6j+T8fRSLkzT9sCBnblbrhGkdK9jnhWjvwi/aqtUr7coEgo5A
FQNF0jEeZdaSPb/a2vYeJ8HLiv1AmRy0pNgpqpbzDW0qUZDbIMUie9xikIumaqxv
xL/wspt5naIclKJv7yW+wB3s0Z7+QZcMlhuxUciy8WqEhodKA44KeVEGR6Z5uiSS
Nbf+RTZLkcl6JubNV88ps97RRuzJrpJkQklzYeGneO6AMg5ndWnqQ3X5fSYrhgsU
zVJ7yLQJNgU+gTNTGW5AVKR12uLCe7vsxR+rs1wVH9CipcbNu+dNxndP0D/QW4I6
zA+JC//PN9E4HxFBEQ8/lpWE9h91u7sxTL0KQoE3pn1Cs+8OVEiKqSCbQtgiViJV
LyCQtoW/xkN4IVy/sx5SPwYbfm5DJ7madVVwo/kGMEVZFu/4JA81qn+bAUrDCGLb
7GDG3zqhaoA1q2km2Lky1VMmho9PzGgsAWWFJIX94Cw8ombnRdQbq8itay98VPr7
56jbLOzh/rG1Zx/HIyMsh+MHKX5CNOuAuph2DDPb45eF6LWtl25R/bkXA/Edc21A
To8/pw/tJn9eHUz566emzg+hWZWZLqh0ZMYzE/34Jq7V1C71qi5fFar5VDLqdJO2
/frLWaFcWyV5ZvbpZlvM1o4pAZPFbzbebWvIDIycPULUQVKvhXlFnbP3+U5xwJ0m
rVZCGw0TTS/zMj+qlB39l6P93mBP5zNX62yMwc+j4bl9eN9l0tzpG6+05HUIyFmA
x4EXk0RgH+Pvksq2lSO2WBTKk6wf0ICxPNOpFICu6UfKmwqIuoLBgU35VIEPEmrd
p/4xjp4E/UwkwJ3ab0P8nXqPgzBgs4nj/aanaTLGuEyyWFt+nArJWOtRqLXnvP9V
ESBYtBw6AGSS143iQkxUBnbLaeSZDquCpg+m8PAIcE8q82HffudF8oDb1qgGoFQF
hPicjdAW/HOK5Dcx3qB+UgdSlE7dkBgJpH7xhlLFFJpMQXU+Oqhddd7iZeZx6P8T
oEUoxyDiIv9ChyTc1kSKjZJH8Z8fMebZwsVI8L6YapJy0KbnS+3CUvNFfEuVoHmk
8piR3Vin8r5DdkgDD6XV3dnLSIuzIEPPxJXRgvQYAc6MfE0FkmVSuW84y8JBc0cK
abHtzEIpR72O0L8RHsmvRGidofNuJxRT+twgpGc04yMKA/9a57cNKNk5P+inDNST
tsFSF8Lb+94Gr5+iYNNuWeEgMxA+uZ62t497FgNTZiMwuB01dDoGMximtowI+Mlv
lGgufJvSg2qTrVg+Zn6EQ8gl7ry2JpTDBjhP7JIRKD7oq9TrEn3kuoujPeKY841w
xcviRV2ZCmngx/GHAXhIBFnMQOIUoYLUlgOnDdy5kOjZjvhxNyPh4N++tf+WDnrX
BB748NAcQtkgY+4o6YqQZJpORemipg5Qdk7ojx1IKYtE+YWUM3LMO4cbbMinxABN
DUBLPaFGfdZqV1YVGZQ0JmvNtEcGSKcOXq2CNwMKrdG6z3vqChM6y2IC0bDoapfJ
oAsFOMdg6zZTvnVOZwhPcC6LRlC0JA7HcuasHlTivABfDy01ZEdKAVzymOouKF9Q
CmfeujR13Buy72WS07kDSS+w1ltWnSNK4Yt2xlqyVbCDf8R8RUPXby6t+um0e98S
ZRRljP3TIvKF45mFo3CecRZ6cP5Bcd7lElaobMgFC7rblqwk2G1i/TqeBg4Qw/xi
tOrPPUZmX0YgyY/xpXUrNh8OY22RMmANKy9++NfYihTHCUvOSZfsdtFbs3IJs9BQ
8unLe0rkJ+31m/VelNiuta6Q+TT70oSBGbwgqlMGpKQi2BFSimAqMgMeQRex/q1+
ykh9liwelax/zOBHGBrAskNlZtyAd3hMJv6rl7x08DJf+tSoqnR48WQLLdrU7msp
79DnZjsY1Qtt2OoPqRAcbNg0oAnKhxaNOkW4etBuRj0ojMxq1rexTbVGi3+7dbBh
JH1WSsOzFW/I21m9aCxpKgLaK621z/KfsMUzJS3TO+WtOsHwC2Jtzh1WRh4IJZK0
HvTimNjaXTWiE5LqBKgohcomloJQFCmT6pPnz22flgdBhv4pzsbPw0N4HS1sQFZZ
5wcMuuniw3fkotWAFjnhUVrFye8f3sDOYyAr2d3zwt4v7i9jvqfIc/e1JQEZwKzc
NF0d9G5OrDcSbspeUQCnsGPZvRgrQgtgWVwfPO2+QTTlvzzk8Z1BufkIYtuCUWeY
50E6UrPr2Rtyy5EdYJ4bIADiJyklF/QSohw6Gt2eymRtbR31+NLWUaa/SP9Gk6yZ
iH2GuV5/WiaSCh7IZpMqSLCNzG9cVF3yQVLX1nL9/1zWSaxfuBD3ppp6VpX/+TZn
ois5Z4UsAbKu6xrw0Gx3EhM/rxVqRJznlUFTZJF7+wTZokp4qRNctgA4zqRBcNGl
8XDSK0FUaltfBYCPGaWPoHcRdh/7Nzkw8MXjZKnUtcAoBrzx07kcBSC1bZYcRfAa
S+RPK4jYVCbO3KkapOQWBDtKJfL1VaMuZlyEeJeCzld0IqeXMx1cOf/xSFadU7Zm
h7/+NLpB+JaH0wIvNm6xPNen7Q/x21wFqQN4JQ5aEEdjLdWO4aPyminhLqF6acqG
6bsekYIe7JRM3+3M+HjmEmFrB5qw+0umWMQirTen7me3TT8mEzvbtSMJgfVZj3dy
SxAykJad3cA+lHxIR3N5wd5FJcr6zrdOxVmMA8SxKeKNYn1LAkqF1kVeP7JnHrrK
oXEpqmjJeFTvwDUJNj3QKhN01X0Fiao5970rrIfTE4C6dDc0OroHyoiUb/ktdXcf
4CNiPZ3G7/+WvaeVDRNuLpHC+F7mC3kDYk3YpE9vQrnd5R+Cuf1WzrGTx4S2DT6c
DJVf9nUP1Xa1V1F4aEtNzBFpyUnlFZZVqkrE/40tAIPqkA1TzIoRsI1a+MobbiAg
RcajANCrqtHvtXQylLlp/5afyctUxS0EnP75FeNNh64hwAxWo1EZd9NLRWL80Si5
KdHo8TdTD+ysMSv+dXoEmllx1gXoLSoS2GkDwiX4DnNLAeqc4SpauivIrQAsKdsM
CixwR/f0UzftLb2+0orrLJqzKEARr8dyXv+XaraAEkyvPyQsaOtMYTfYxhnKHmZE
N40VrYRLZUwvv9cohf/RZy4spHRJ2PKpopre2c0B+LdHKWG6e4+jlMo8nebV+WeK
sIdsWUUsBb0q3GTECiRdccGd+7yy6JiOjhs0fd6ZS7ZJA1zWGYjTsF9F6eDMXtBj
GUO3oDyq7ZlI7BdcJRNdelvfX8twXpwTnFxtoH54VVtJt0IM8AsK8RB5qkKl8Vvt
fFi8LwKx+oJVOxUTnFc3y+dEjxUqoA2VYJblu+KJEi1vChMno8e0fpaqFFnbRMwn
irdaPQBN/c0pG43YAShEmWAXDcM68YEzPPcHhalT3H+tWfckBasAONwVu/cdzBRo
FoHcSayEGV33HJz/kRFO5HQ61G61sFJ1z7Oa/7v1xZd/O2ZpTfDrfmNZNfobXX8+
nJUWXirJZwUajaxFllm42zvi5GEYLgk+1fiZYkvmNRRndJxrqABsVXP3Yxrm/cNY
rxH/FLv/TfyiqpmLIOLj3BUFHtAEnKXBeWG5Tue9z+MDt29DVsvyrwBvP1plmcJM
8nEsE94T0BwP503fMM1R/MN4G5G3bSUeJWLvzMlWSYWN9GpAN94V35NyfzLcMDZl
4c/pj8lfm5rHRO2qtSoOPX9HOxg/uZlcg2V76UrL5sLlFGIQzjm5ybH9zs1v2fqN
uZQ5ciqiuCix+hmmNoUbbxnnAmKN9F2Oi5aecEC7TTHptata+2ZI0KQKQjrPkrNl
V5dy2o13/9gYw2DXcHeTMpL11yF5lKYHnxlA7qGsgh1aP29aEantURsZGkmWJmOZ
JkS5tXU0gjXkkw4FgJlx63htrEEs6iQR5tgaKzSrFMMUAGQa60AAUJMbhr2c3VFG
3tzN6orUe+cKl9f05W2HqNCc6/kj1dcgQx/Uy7qipMRO+ivOU9Pd67rCJ+2t+TXh
+bAqpVpt2GLH/n2UmJJzSw2e355tWYpvwEkM2pEimFjXjZH3/MVDlak5LPfaudE1
/Wa6frEOOhTZQ7YYfTlF8I0eud8GIFYvWxhTZL9s+cbpa6gwnsMkKa/nKlJj27Nk
gYGtwZN+kqkqZBqZc3aPUh++2Hq/FD0/nPDlpEP4RdwGywiQdezhwzFZQpuNJSi7
MKqrTEXs2gSoLTw6AwHfBL01HQe7AMvnaKjzt2GCLXBDomLxf0N6wLBuw8VDL0uY
h3fSSWpgZ+VgC39devZzbaZrIcnlNEsIsITjihsT/tVOKcmYsd7DKvTlHT8zICAf
aIM9mPg0Vrzj4bSAGhN5u/EtrbdPVH3113jT1seqBLnKiPN2TixHhi7vbq+vWcn1
iRiqpF4bsVlCPy+Lm+w7O3Lmsgo30g0OHpcLHNzzE8xAr4Wxt4+Jl8Rnld3GxdsS
zcQL+tig70fPWUqVOsS9Ebq1mDNGsO4rlGQdJ2OUHj9HjGHof8wobnONqGiwzRH6
bwuHb3bJGzK4vx18qNlVlMVs/dY5YGdKSDTgc+wUH/LVJhU8i5k43LCETjPSxtx5
YnUJ4Lq8/birpd5HqxTwXtiHfo1/pvj80XRaloKCSrwTcROz7K40LuBFkDC6kCOx
jK/ztC/j+4Wa4wvvhGGM4LeRP/YSb9uR3JG69CDZReg8wf1Kz7zZhATBLbfhtz9Z
EpLU8FkDpAUFNr0XnEm17DLC/7GuNmRt7Nv2zTypuEBpjylRGbQLb6w5ttO18tzZ
8qPYsSfd2W4NJHvvfngzIEgye1TESW3dAUKFgXBhGthmLaLvShlRd7eE5BT6mXZf
yk01FwSGhzOVabdue9ldYaHn9Gus0+3skpVr1LuEeou6+yalpfXOAk/7t5663b/a
UJzkAwBbzG7Fdq10xRVUH8L8sF/Wv9RzfiPI2bLDUmUdgB69DJwqFdjLJuKyTvB2
skUztw8Q206LDBtPViLSUtKjiVkiiujwH7njQvA+h0cCI/jMmLgmAAHClbSdpgS7
BeuIQkcXZIne+nufXCmGFDar4uKLK2kfXnaclFB26Gvy23fgGKcNhVIo4VPGVHD6
fyrM/xhnBjm5jUc7d15xzdp+4s+4lZO2WJEcf0jnapmGLeaQ3q+VbZ/8+6FKimLv
NFXef6fuVm+QnHVcgHgrmmCgku3wWREVOIXWXA/p6Fnbx0UEhhWO0+q73JcdYI0S
CB7Wf5QkG/csE0OolEQ+/BUPzLXCTXdSkMShHc1woYXLVdTBuDpAwxDkWExH0FdK
zC0ad4MDHS2QE90celT1RlWlrp8VhkeR1yTf1ypfT6HdN2pyNGE76KFG3BMho9rU
yfJpp5OFRiwC69Eqh5Kca4aLl9346lrazv2dHEsbeEDOdx9xnh64tKs2GL8FJzsE
vcYlr//eHjSr5pWAZJkmVsLW08+frdk+W1u7ez2asKp4yVXreaGlCIIxjKO+RvCI
wq3nzk+ZZZuDcJp/xU6eSbl9SWYrcQcLvYz4bNhg4Ejr/trcD+XATOGQllOqMrZh
mCenQSHfH9RkYqjcXxzdnqthCxZabF2ONSUP8aTOXOu1Su9Hcju3LuOVWAVwFK/w
20AUi9YWddYXkIXhOE5LUs4obPrxHckl8wU1HZnzvrdwLXqr8c0+zF9w1fR4DQwx
MTbsRpyTSKSvkW17UOt0Iph6vK1FiSVr8N+65NgEqOJTeeJPQgR0KIDGc1LXo13P
/nRdgIHx1vq6E8jdwJOOuohjtacpEwIAr0WTJ6aTlQOVzBVNhx2Rlj5A5i5zwbym
OZL9FY1oJqAFDfbttDKbfdc8nDV8A47PY3biFy+IJ9trQdqoI/ZYCMW1fL+e857q
PLzdRX3PuqoPBNT0jfXQOb2e+1ivUOuUWutfvsNHDwRARWa6PsAc+7Xatqq3On+Y
SlcEVZVPniSRs7+5KMQ/gvNiuqFKsyMPzPNN9HH0xhn8ZBPnwXGYEcQHOhlrZtss
kCwdk7kZoXy+eqYvAGhcv0HZ34gKU/FR+XDdIHDqhTaR7zO2Kyms+ODgSCmfIWcx
SkTZEGqYWspEE1JbJ0c/l/uAE+7wtCItOrL/pTkUTEJstuQaaEw9izeFA/lJepwe
6oE+HA1/e+S6Vcup7mzJKV88bIxZO2WX+BPIe6AJAbLjubn74nsZlp494CL4wHzU
520KdzmCWHIsYz5WvQP/nMQFKQLBVT+6pCSJCQg1zUMZ0XbnLBZsnj1npPELF8LO
8AWG/pKj+kKb62sGFATDlTaUN+HfpVnq808lieTzFcaKCRnr7ksPsxRu1F8Z1Szv
OPSjTWy1Xj61BePArm4aqtNDny8XgeIo14no3BcSqp7OCfTtG8txD9eBg0eCEy0a
+Ua4aUB9TTfRxDxOwfBNQqBo3OrM0XjT0J7OlZnf0gTy9akeCVQqEoOr3WU1Nich
jS7qbyA1JgHYOjB6nYLRzdO1sz9si546j8mZjbsyOHJDt+4MqnrEZRpU9CSmI/Lh
JQjx+1l37enK4EWB23kWt/D61FDhJgsRoc0a8SQsjDzZPwd3mUAswJG4bnK1Kj9z
esmBRj8cOORKyaMw7h/OCHVVfcEotkMj1OGfxt+9kOzKgxwqEPLubRqIXx3jhR9E
mUMCJ7R5ACNFdEBbrA+W0YuKpoqOmzcWsVJsN0SkpHuzqL+8TsTeILndM65UTTcq
A6vHH7MZvaM20ntNQOsJdikcYUVwX0dX8mGrBq5ncs1LU3sKioDa2dcoIHAlL+hi
Pu91GCDj9gUM2+6QsB8tE/atp+q4xgR5FMyEWkBF+wfumeJ4lhF5dEQyN35loF+5
vQDDeJI5Ix8NFDXl1YZeBvz2uEk8e3c2Zn3PN/lT2/FMXwMX38zaqnQ8VBgMsHjL
RyvqrG/ynlTIbmb6yG+cjjdF61XywILaIExlkiYPVxYBACdMJd4p9POC7OZ+Hihn
VQQa1YmdnM8wtkPQZ3K0m8PShE3Y6rpnZtPFHzDRoW38sMATeY54/A/0+onWyuMM
QqFNMNXPVTiQgJTkMwJsZ8Ja4sBp+KnlSq44mOPKN5iIlrKcXJC3vfCvhBGa8LqR
3qjwSrI8JnVaZN5W70aDrfgalyenl+Xi2czlQIwvhzOMc2GjrG2ghovVeeSEx0M8
UYWmMAYP6btlzPHcpNrlvSWqIhb+bk/Hg/TaFvSKd/Cp2yjSTPr9kLCVbbnPILWh
meIl0LrzOXWUTyelYTly/h49+Fta1G4R82O5pygJ+ML0ifjlTKwJkDQ25jW0BO5u
IZzCr6iIHr7krvjArGAHwcu+wolRZ7Sq6F5c83f6ar7zQql64yFa/JTAaHMWyXsn
8OsAbalmbK9mJiXvLuFpSfTgMbSSp+f27NiAbhmSl3PhWTcYc0WZ4oMf/HpRPzJW
ApJGSCamYX8QPyl+75+p0uDda6TtVFI6GP2yQ/w3doDbsojOXMdUxXs3Deyxovj1
GS7ktRe1HSiE6LAu7k3VLzH2ghkE7Y5W33ufZVEkDmaAkWemijfpVLlt63Nr0L9n
6zEzvFwXL22myK9+00m8Ci62QIHQ5xNxfrswUqgnQT7iZ0swPMkM/fraRWW3LtIr
5msj0QzLJ7ndV0Z+vzFEtM8WQkdj7/uAb5JPqJ6OZF48gQ/VeHvcxADcvo3nnS/F
VKxLwZ2nU238f0DhlqLxkjZXpdnw/76wKNMOKzxevO0bN9UXQf8v/IXwqAptAy6S
9H2cak2JG+8KiZjEVYGNWbiGqB8MK0wV3sJqwANUTRO9B2esbp+LhFdOYar7pTpf
nAMzmVY5HQ7pO+ydFcAIBurlDxhzY5+q6g7hOaVvHSEdnwtMrEh6H1Ffu4PmO1mY
fOECnkSJY+wo6rn4Au++9s7W2ErHBsB7L1ZQxj/afGp6VqL5Ef55kdtsaapvuS+n
d2gt9VMQ1/Nf3sXgKEnGvm+nbDjytfK/8mLI59hVkS3oJVSBtykYae33N4+BNNI2
//iyIRbDi0KGZf8YzwowgT8TrvCCLmDtfpwAsCQMZEOREh5tLCyM5m7e7FVtcElQ
M7mqCAXpQWZ45QSJsD1bKoWdXZQwBTpKyuhl4XNVgH8rbRgt1eUiEcMLLKNdBDaQ
z6o76JTyh6LzPWmc7cltKuDH//pVsFUy2rdRPlyddhnT+wd5Vu6UweFK2HWzcPhs
QNwLzJXDTU48P2E2pA6TudZMBXkZVOPNqDrU6eSdjZVhA83pvnS/Htb9gbJhsF7X
VTysqHdM0xrg0VaVH4TRKwvWKGQ+Z5L3Sy5B5C8yAr8qjnkr94zWiLpDRTbdvi2F
kHUCF09dqQux4k+INNYUXcwlL32WgjxuttWXFPp1s//6GSWUIdb2lUXjUjScSEFh
DERFwhxNwsYu+KmykionMa+0eo5Aa3jx+ABsOMp54j5ZTfAn1/Ks+ONO9JfFQWq8
qNUNVmHX3V6NZFidQmRJAG/x2ykYkrPLe+7zN4ZofbteXUjNFNuchiigzL49GIkt
8C04235e1al7p12EoVo1P9E2SWPxuRyaTbJo9c2EtHpEVw0gu71CbWnsspcqvejg
soU5TYdZBlXyugFDFcH9+L43Mtz5tzl88/ce1D56BoHDaLnocnreEYBTvkRVEE+D
K/RfC9mtMWOZbLAniEA63Qfr36e9CkuG1YP94GopXaiyXSJLtNUYsEd5DFLzk031
jJ3hW2j/0KZ9hktHXBQnijIFcXHQg7F4CxUgEd3ebtnnWiUT0D9bY2C41wYgnzaQ
ab3u2htHSzV5i8euPjQCHdTcg8ckaXWRka/zXboFGVC25YbiJdJgXAgRKOBEi0pG
UH1lsI8uwmR5c3k+Bh7H1t8S8yeXKMZsS0hSor5OjO1a5J09WdduV8j5jQ93cwEt
4Reg2i6ahztX4MGydz4JPVlC5ua6q2gOU3rzlTMSPP8z0nKBSPjehIrk6dBwa4sA
EDp7W4VVWfiCLHWzMDqn9SzKAh+p3I/94dUcxO00VEI1s0cG0MSB9w1kAp7jBh2X
02tcvr5Fw7++7e855KerXySBwiL4JmRF/8xka2qXo8sN992rBY22vjA8ZeC5Ef/X
5EMVoFbCGAeNpF0R96tTr/9fL443vFcEZfB2Y04/oXE0d4MnKJD2CEPxThTxm1g5
IgfiQu/DDDb03rmRlLC7+L9+jx8mnX1FouLvytjFHh4eymGlpkZqstK75xj//Ub8
m/xWQtdpX/ZNVzqrWmNGThZQV+a8Az6vN6XhS3Qp4DW29M+0Iniq3sMUlHnnPhQ1
/ZVQ2Ec+KBVT/B7EZDrGjsUWcSeSTh83CdjCZPhBeP+wQAelo7bVFQk4LviDst1K
vCkYCTmgXKLiU2sgwTwCUCtJJeeqvoW88RhhkZiB/qo6L4nkGOR0FrFUuOLXu3ER
Kdc/U0YTsOxjk5KyzPzl9WujQY+hnSB521QGQqvSfAyg+b+pViOKRDK3AyZRmTAb
LP+0YoABvNG2STL1V9iipjeS34JhbGYZl8MBooDD632dXxZgS4RMqnanwkKYhYuH
wneYLApqVi03/ROoyBcnTFM+kUhvgCBDzbkc1/FAMXcmMiqDcQamYYdygxks1Pt9
8Do3fSYAXSnTouPTgzLkqWzr0zAYpyhBVi037h3bGfJ5zZp6bxloxeasgEGH8Xds
RF4ZmxyjfPeVxglpJI/yTWIoPRsT7+lMkaVcKGN5kSUzvbwZiUHvjyfQPevbS2xP
yUrfuKF+OR2VJFMmGKpg6srbXIq+XUySxn6j5aEsh2W30Sx0C6yzJUlKvRWN4BgS
bP2UiN3k2iXFLDVzzh4Kl0fcNHcFfqPmvo00UcJNqWasb1nLz23c6v/J8HkB/U7r
N/hkDYBKMy+7wGnnFuBMUYBNIOS0vmGsnUTRHa9dAf8tcTBeAyDB8fXQ4HWx3Ts+
WWqroCNOEhtulVHdM8R6XWh/Fs3TXbQsJ9AEbjAxAw4Si6v264wdB27yhySsrm5i
HEwxHWTIXF6RgPcuNCEefUZ5zEFf9hJcE6UlFTbe2HTB3cjl6JLs4IOZCE/22k2d
u7wHJHLk5kiKac7JrAKhmO2geJoiCWnQ9CAyZ2smB7z6WA6tqVPs6vN5yi8P8niS
9QzR7rZjfnx532XHjLY9VTzgriqa/DUBY569K18kMKZPSJ9SuHZrsczvZi0imRTc
I10pj5BDSFQPIe0+iloHXbgu0OsDcAYekBaXdxnTInHrjFq+YjscABVOFvoa4yZ4
+7ua+tbypRzO5YIASsqKeRRRQxkvKi8zgKXG07XfwoYtyf8KDg0PoV357vkkqGxd
jzx15j+tIwmFY5MBLIl2XrBxHwbKjVkP9wVqzoh6BTwE2XMWk2LAKutAQDweY6Qs
9cNS4zTSSbD9DmMysFQe3fIq6vzoMSP+JC3PLnj1i2JKqz/PaXn+8oKFCr+RjoAJ
vHkeYLHPBtv8PAdUKezfFbXjnMFRoS7svq8Z7pAnIj7pWY6jcwtpxXtvAbsVKT2x
OSUrc06lWiFAkEZfchARnZscGslo+s6cUOEgepwyO1ReFO4GHMAm/oMbPX9+wSNj
aLmH07AB36KKcbeCF4t6IV7eWOmJX96FNF89ssDl6mOS1GZ/LGTb63NP14Uo81dU
6z8iRX3x+E5R7YrXALTCRltg+JDAU8Ug3ZvHoxeYMAB8qYNZT+QhFxKZKsUsdYO0
KSjWzT+xB5irslN9yCmZ3MOaMQsO8OuW/uCdmPbuz6dAgC8HtnPq7H8yFHmmamDI
gLOkpnrWREzsMz0rexES0Zdfe56CRdyafL/UG2pUqJAUdmsPJVymsIdOByaK0N86
HW9dn3LQdjiAN1mYmUzLGTVHEOlJ91N585WIQO7Yj61sxc0q7xjLfm4MBjU+dgFh
cBPC0elzXhmkMwD/6KgBA0c4v2DcvLdADZB7yrPtyV6Kb2hjNdE6FP3H0fMRQibG
bD6BIF9LmGRp7NQbflQUQ6BymDxhdTsZjXX7aaAYvGr10ZAx5VbI6dFzsvGILdVu
9DPlzKPo1pqtiMBz6+5KoImay02HdENf8F5z1hGhV2h6I9rItLtguZjGxE/hk19q
RCbWICbYZ/7FGJ3vcPPK0sRtw7d9STztM/en0Q0LhmkuqdX4xaxx1tPl5gZ7DsQU
qbocJ35lkm/xnam0P4IaqcI1qN0/b3QMur6oul9AOkYphbpPcrrrX2xcvvWEoE4r
/h2bU8Jqo/kmi4sXurDf0FrggoomUar/kVUSG/X8NiSrWOZP2hAdvRu6xvceeizo
aezBNu54o8deIybnSA5tjVzRKEf2A5lovnjBmAXgI+V2EcKcEpfyN++0nffAQkXp
c+Hki3gxjGa1ulw2Fpypw5pS4C+bmW+aCz6zhYBZlFBl3VWgLjvBDZmRWhf3v2UN
HYQqMuGIy6XNW0ieEmRguiTpaQom5BzAkPkyF2fcNscFcjI6AF4dJxXYXENM7n7Q
YSFS9Eeo3Krad+4A0EJ2syuNfY1fhOrCTTTy4BhV309svaVRvaED4mN/l8DsWniJ
YoLu8WjM6a1wMV0Tk151tlu6WjOfPRzN/gNvyVukCgSfVLfkMiSSEHIlPwLfPFxj
07SVCfnIptLOlm2rFzm/4UkbOd2nCtOqP+s2i3Wu8HkQ8vEFT8fn42GcLYfzEv7V
pdn+Gdxmj1ztHvFeP3iUoANt95zm5QQvZQrp2KLJ2w8crB7mBrdeJrXj35TZW3ZZ
fnidgLnoQPaW8rbPKuUaHa2+ZhvbZg0r0ZwBlo3uIBW7nqWkFGyiud61M/YyTgUk
kINAVbXm4s66HeWzX8F+5H550Brvb20gtum+FGTLyU+y7kb5P90Mm3gKTJl60YP6
hifnKKrx42xJHeFg39gltVZOCH0HvCbfrdV0eQwmH7UuXk3ArrDU8RDdMtipTp7/
jkRzeIlNcWTUfgEdrOoutYieBcu/55kiIB+zUMtM4tADd4I+UNSAiy+HhBgLzRIo
bUVIs1YiUsyHDs72+AJ+AcAkhvJKRhzwuNGS3Wpg6CQzLteE7oMlrCWQZ8JCg12X
saeloXHyZaY/gH6ZKGRlxQ+B9Jb89sDs4cS8jgYGhYtj4MiPrPDsGl3RKHiDI1wp
teZpBcPZaq4zSg9WaO01BHh+2s9oC6oOnaoNKmC5mOGLvjX56PsNRuBtG5Ai3Qvl
HCCQUma0V+6mepKfEPuJM3DpBK0/wkfCxf4ADtSDdraOmHkixSQwT9CpktXzWTpC
A4ZLsg4vu6MHrGfpvGQSTSWw3Az9dw0EFUCQE2C0EcCu7uBo6CgbdZDRTYttR9uZ
iHVu7wh1QoShIZ2yWIeh93ereABNbzo+uSfSbjDVBDLY+wQp7EbooVmip4UsIifz
s9Qqdtg207xatYVO6P1GJ32WIjbEhEIztWNFhFjyGXGFuFbsjacIFHymCHuGjhM4
EgfXtQ9fKgTf1Jp1M/PyIZQRhphHYeV9TkrxbSrPqWnSYVO5oTH6lAk7SSNMnKX8
qu3t1AHUKUojH8ltIJw7qSIl4q5DFnu3vZrBbqFsZNZQMKzt0LJoysx9M2cbgw9q
5UGALIfJ97rDfr5NkVXB04WE1RuI96VIhyJplrW4PWPWVuhBUjaNKa/Pdwppni2D
3Kjjolx2ynR2xC5nQkwKsVkvLVI0aU+OszpA9QEpRPpXgJeZ/qQECalhdgNol2bh
dQi7jftB+UVL7vJPbGqq4R9Mixpicx+GdRT/ohzitzsa0UKS+/5kVPIboDZcUs7D
CTdJarC6X7tvPzHvgPBV6YWmAjNDH0IYD98e5tKT9otw5NmJ99EvoLWhqiAwG/nZ
RJiXdStCWv4EPa6qJjaDbMbexOFK521Z5Z+f9EJ66ToO2jim+GCuuk3jYincBx9b
MILFVWzoNUIhats10rbB6rPNm2WXtr5nbmtvpZmDosY+uExcGxbKY/ngcmYwZ8jt
9t+hA7bnea0PrxnL02+wTDHYwb381L0Pykzqvq8AyAzRvQ41/C2uHob4VLGsFWcc
ZHe5pIZhE017NCFCt2P9++SFNid57kqU2mTNaEEsltZIj+uZR5tAYAINANlEWwry
Rq2kBSORRu9+YrM/BPpLfiWBIOzAkYFA+WUppDwEkqkT/N1YUMPutf3OGhafttqa
ZLtcbvGQRZ6FkActoB6tg+nhb/aerAcphRaSJclGYhaY67T7C/3jDok6EJMXJCQf
rxGACyk04T1ZYB7V5ztLupOGGx8QUxRQJhDgTG9wkpnH/HlxoV+Tb3omCPMod/cg
0Yf1IcvgYRHxil2Zn9HNNI5ja4NMQ2BFLA9Nf8ogLyULZTVCfjoKbPS9Ha+RjeX+
idAQF+bpqSuzEwLnSHdVQskTYEJ+LRBmrymgnP4bgQEqgVLDU3vWjUkkVFvjcWew
Ch6wObXw+uSKcxdM7clvdxkm3+AF2vHTfnGAf4LSJgiAJebmxmXWPHA+qaLvtZNp
m8CL+zvIY3dmCNlMTsHWJrpTEuf3PcTi/PGbAfF5TdqsHM5OcGl5y/5TvWZu6UIO
5AcyBQrWPZhpCJcbytTnVb7WViK/Lyhewn/YjLDtr7mJ9O5ynWlSZM2D60+ujkJ2
8PZYRvN+C2AAt8SncNHIJtK9ZmpgVOc2hGSF3oY1IkSLcqIA0SXeiig7hBXD/vtD
XLXr0QW/Rz6jQbZnNZYMlhK14/NYjYivofQ1ugSJHimsXB/abWlF0s4FVNTD9btZ
CVhsEH8AGX8CcnkivctIIw==
`pragma protect end_protected

//pragma protect end
`timescale 100ps/10ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
OvCD5cLs/6MQHuDC+4OaC6fLTaoGH4gKOZ23pPDwpPQgzo16CfB4/FTt59WIxrML
9qAaZvFnxYPdW8L4fM3jc2xpaPe6TY3EMC7woyaMEVVnClBWbm1WzM0+Tgbzs04D
nzCyakNaHiW4Obk2djAkdRx/RNhJe+jNlwRG+UM9+2EIUHSulT8x3oC2vYVvAwAL
A/owLgTTHP+G9Q/9PJN8eKTbFdZCkAumypqpVfqN1lPttOGyTw2t1oOtfn5Xd38M
7MZHXfcs4AxTBMQYyoII5lzWj6IH0C49XuuboQ/S6ZfiLS2yvhC9nCTKJUa15Q3l
QAOnvzqM+wsYXhu7wUWguQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5104 )
`pragma protect data_block
R5br9OZBSfHWShQcu3cSqdZv+odFtoMpPOHZs2MVBqGSVjzTnCkj2L5WbxICFvx9
MqqosUfdMwjX8VMtlQfesm3RYSb6CiP7SLRMC32VaYud7nOFs2+/q0XqDjw4EYXM
rKu9XYyX8RdUiJNyhqK6MMm1M7fFX+URXyzMthC9ezY27X9YDb3nngbMxwYU3tzg
HPcaKdGPejozOSkt4XOYMFwURZRfToVwacsNCJbFOoQctKw+UY9ueE+072Y8dhpM
6ouc7S9bv/VQFQy8KgCH0vsvrqPNBssWCLB5MEFWL9gcDZz0qceMRtoIQ/JngoQT
RHQyszg2pWNcDp5swDPKfk4AkpOrUS436WMGE02jicRnu9j2NVoXadGV3REwfmwu
CmjmmM55kzzezemwLw405BGFQ0bntYHeIa7hS3eUjfvYRX57Gh4C8qQCKUIPrS0M
rizZQt16kOrsOqzIiLnnT/HoXanPkCLOztlfprTx9tZlOgTLdYT34CVT2iwd9fHy
t7KHx6lIHltTlhf6a5U16D+5xgoWB17aIj1h4KYVWwLehjqhhgEltwMaYggKH9n/
5xdzpLYrBzU/G8p3hiChgUo+32f4E965nr9kHRFboJLiuse+6pOLUrOQfkPbhBlQ
geBd8N1HSFIdw+Bp6JxIEYoMGl3PUGH+b2nyKKDVFanENWQer2b0Vc2pMKDrP05W
Xp46pCZslk55ENZ60LqyON/yFDqSvS2tI++FIJQCNV+kjyCzymCByLgCWQ5bV90O
SEUubxbrfo9uLsULRWJQ4h16XHvdMoH1swGBNtLohSbZ+mfmedxH6hQjZAWWZA9/
l5srLGwC4G4gPmwppbGmDfQUoN0QlriuDgl6Drk81/cURh3HolCepRSnrdkaGSfF
HbSTp4g9lG4vbuMOrX+FuSBrpHCUrkB3XvjcEoeq9B09eAH9W4zPs5QZjbUazeUJ
JOzWkMDZEtRWuaWqqaFGnBJbLjX6B80AezCaCxewT1umEw2lKjSJ5EtU0OvnbzAc
MrQ4zjC4kI7S9IwVA9JywawB2Vo933+BNIRPoDYJ8QLqc9rvX4Wyj9ACfmZyqtXq
SYe4VYwo2MP0DUHz8ps03AMkhysj/kM+GsQQ3QVOeAtBrLnZlkD6OvkXULlkA77P
HMx4Z2Bqb3IsmuNYMABPdS/VFXA2siwjBJXOC50s5h65h58mJvjEqwbFzeY5TazY
jdHylf9NC5oD8wRVkcCp701NhUW2jgDrnAVHR66g5iolIE0KXDeeVGHsOSd3Jon8
C2caFaGMO/bpBINRCVeAa/Pf0TGo43R/xOwRMZf41wkbDmpx+JV59L2ieHFqxYrF
Ze8fLoWQk0mc6OhlzPgwzNkN+V8awUtmSQ9fuKCt3GfJmjxjXdcKHiulfYSe2t+M
TqpXNAANrEo5N1jhXcYTjgfHtz/jxszUZmwsU968wqD2q3JjK1G25sANeOUCi4s6
khpoUuHHtY2Bqi0k6gsjdHOZFgT/WCUwBQdqXkzmUhQGGkND8DyBBo9nyMgAhksw
QBU2OFi6gOGHfmRoqCF04uJedESnzDXo2C99WHWmeprNR/9qUnHCrPovUfSNyMg5
RrHU8ArDNpsdcbuyLW8aN9uu3mk4JmV4Js/TTpdnF8wWLBngHbibhAf+kZLY+HyX
REBoXU9RuHL+jlJphBAl1fWX62pAOqB+rmCsqpXlnM94vH5gYraKWdEoulbcHXz1
T1poa63BCZJi1evHuVD1FEmFEXEkgwhOSTroNiyAuZUDkkwpqYCQ6Cu9ZFKyCQ64
vF4AOXrs0oCguXmRrSgm+bJQDKtUcugJ4vhtEtH24SQCb5ixwPf52F4liUuCwL4S
IA/y60onPbwXb1WtbOwX84U1Lt4Ba6kUDlRU7KswQ9zh5iff84xejzc2JN+2XCMe
VZwfNNsSyj9CZVRItKpvH8qqvO/G1g1BLF3Fz1WYIuLDXGGNG1Hk7A4XLejvADFM
ifk752kCDVbmOjSbSn4Mtoev1vXnOXt3s7/F3RMaHquKO/wb6U4VQ677rXjackFk
CpA0YuJFE7ci+DDU1hm7TXB/dng8Wonwo4wpApr0AulP7WWVuh8AycEN5LaIk2Qb
E5AYKwUdDShMnyJg4UW3Z7WuBHqEDzgWTDMTZOGqubfcnZG5HPxAKTS0vU3fB8eI
bNRji55Ac1sKdI//Ykq/m0j1baRScoRsPaXJHENacvkfJGIBEpIPwTP4KQg+iUXL
ZhW1aGci5ci5h730oC55LXK3b0wlLddU2DFu/EgMWj/FgtvMQggyWL7Zwor7Bl7B
9R5F2DsWC5+3B0izfFk3xdh06QpsWmWYhqHrb0zf5kcVczC0Q+iFtobaAVt3OGqu
xXqD/qBJ6fUzmrkoZsmFR5yQkytwskLprbPoeCxm83E462M2IHE1gMisFxIKzSiW
vNdvTOnwkNZrQ7jps6O5su7KFHM5KsCG0DNh54Gu6KGHZd0Dvh5lsKjRbBTQM6lk
U+braSS9HuufUO12Mr2/Adp/5avjpWkjOkXs1YVUWsK5LUMiBvJyLcmeILI9m1d4
3AEoweLH3xWBh+e5JPIsJFyLLP32jfDbce52rWf9LjwLpVNz9WgS9zELztZKWTX3
DJxpwb97gMhhzF9d79uNbRj4PG5ldRbhNVMs29XGTOjAzwQdSby3zslsOVZawVf9
I4TGnRRDZ7iuUO/k0ecdoIIR1bzwmHiZmfxS3QEG7iOP/eUSpKYCOjsnU9MnQV3C
jegK6etviXf396V1g9egOB96wTWrh1N8ReGBuCp+Wf6tf+RK67y5BhpGyYnJB7k2
/xlH0h/nJyzN2GpghbI6s5mV4cW3VWmAJ8Ml+qCdGKdcVKlgLeHZ0u+QJkxhoIqf
HMMYEjx2O8Qc7ftZ5BnuR8I+ntKVJEuDLi/uBP0N/g+8Dhfvtzs0a54LymwxlMcm
LmHQ+Sgjazc1lxHs3RzzaQ8jcjbvZktgAs/Ss/d6T18R++fAXGrfMiHxzNh4KeFt
RqNthRfTDKLdrUkvLoEC0VSrnc0tiP1eqtLENHLRp/lExgJ2WIGYZREjXe/Bbrbq
IsK+e3MqDVbisFR3/QiUcLUZaM6QM7D92tV5LVCLhde1k3/Sk32RRaFb4bUAHbQ7
haHkhSCtZRpVv136BEy77XjaGiUwmR9+1X9R4RTSBS18oOngoG5tmkGmpaKIeHhu
6rp4IDslUSyspuZxx/sGLSgghSsrvxAMOjjFPctk+BauMuEODUZZuoOl9kEYovLu
ag2J1tDDv/ZsVUytyMIU1N1tGwz/oHCTVWXjmhwzI5DvGgPBNrI5Drn7g/OnMtwh
1SGm2gS9H2hHWHyoG6fvdUKwpkak5D6vJuki2DHUVAtoZ7BX39PWvJ5FNacwN9gD
bFuvf+l2ReWYYgmEPcjaGGBbuUCN889MtIlhXy/Vqt0HpRr5xZ2s3LMRLk6QHrPt
YuKdWuBV6u3+jqMtGQ82Um3GtSYKjSTLMpTRyeoY/yiquoTYeVk6Vp7e95Oo/0N8
SUp3wJwXPMhsF1vvX73lUklXW+QFbq6Ila96gWUB38B+bHiNw1W89QcWlKHz+r8X
O/u42SrBpZse5+wn/bCLlE4Ey2Nt3gk7/ci5Nbb/XZa1t9kgKgA3v8DsxqVeDJWm
fRDb/gu3yhy11/iMWtS3smq5T1Ihwm5ZWcxbvJ4LopAlOF44i5S9/8kCRKfws26/
NgqfEbaOb8EalEeFfecFSWGjcjMfJ/v3Wty0bZPxJIVA+xhBsR7HsDHgXsnubrX/
gO5EsN1obK+DWrRp7kcII9kqklmbOD6J5X9Orb0UN8ezPY0lsGVL9+Fz+YVJUI+G
IffWi2E9bf0rkpZoH5ou0gxUsTA+/vECAjCx8sT8h6oDep9jIOxuzBGB4iPTMN6C
i3NNJrrq0a++Y+Nz5jgMR7YRpopyGazhU6YtVkLjF5QaOIg/WyaRTVWnWLLcn9NI
4mt2eucaPnCRHguBDis2YEO9Ow3m3NfAAHisCO26u7R0YeGVNK9fNMGy9BkRIAkr
jTMC+IcGH6OxSleoH/yvNKevFRKSj6uYgev+vq0iiw2Kr2mvyMeL+Ez2kYnMCBTX
Ul+JqxaSD578tBm+lYPMkXS/d7uIGjSFnoFpAwAjvgDxd0JCOkxZ1MtXLD5tg02T
jSgW9LQBiHJjOQVubQuItT0VlBslWSGPNTwHqHQl+PEUJGBIVbSSLHIk7F9rXTNe
eC+x9AWXX3F7HjoyAyzVb04fjbu2tLbJlqAIpiZXfLOuVUCm57JEzVmDVC1FEqWW
EYI8gqWDzWZ70QkgcwLyRSdyv8lTG64mCf2mNCQKsfpl3FaVCAlzXLFZpQB9h3fP
chBI3nCNDm4RZlnKXmgsizVL8dD6jfgDVbSH40k3fZrAX8vbDipB6xwtjA/SU/1Q
qwUriruuas03ro9KW89m5H92B2UaiPhnJ5sT8csFa5IdzJ8MATRBvRJGb8yG6Dg+
mkU8vl8arKqnH6P3B0+zQvnI+ZVvZUE3yWI6vXTJYdoM5cBiFK3jyvVlJqoiBMnt
TW2snqOz9tv85bQ/PqcSibaKv5pW54jT5f/VP1PitCXyESELRlzhCNlUSVMoD8Zz
CPz3IS9Ruqkc9DsSDo0XB+3Jot8Dqbw4xFg8UwUXTadYcDR9Rk8Yj33D+ANdjB81
EW5uG0OGxqlQf1IZ+RC8Ig3GIhWqK9Hmhq784cNVDQKYp5CLvLMbFiFfu1RkSYM/
4+l4YTYoz6z5PkxZwKnxEZGeV2llZxCAO7KId0GF8HtkYqjbiq0r/fe+aNfIij8m
mRT1sYayVmUAPuHam7LQf28nQVvQI96xoZXYooeOjOqiW3hhURAefeHvvJmLIeql
DaJGhzk5YJr1ISY3nxEUuU5U/pes40VjdxyZBQawoEuLdzcKka+OsAycVpU0JL50
eCZbE7hErUdXYMN+SByVESppndF6rB/g0g8Pp+HJq0PuIpFkwAYghPLKs78zMlaK
ylSJi/LgGuLWA96/EHulHvG5s5IXTMuiyB011aDJiurLTJHIEOKOZfquYEUouURS
i2Wqh2uIK6zu8dYKpHtYF2NSvlQddASf2y4MrHCG2GmYGJyCu9XmdZlkGP++2QHp
4Eyy9iuQvafgadv5IhrChq3c0wyKflnMMmJ6yVCC+ZHmClWFE6kCSNtvoH1VLnHf
3BnOqcsPCVpV8Brqsnkj6+YvP0f4egZhGajtf3rPiVQR/E2MSV4TXYP0JFgsjqXI
IER+TEcTH7tbiQljK8hGt9/mc2El/FE1SppcXOjG+DT3CNey6FjU2SwSHtv7mQMx
p2etMiw/+vnzf3W9qABmw1NXojbHo4uCjOqbLSNWaAQ+1soK84xmigfSBAq1K9ND
cU4CQe/0KGJXr8DUYJTBv/isrRytQ3KFoYAf34WH1THOf2btAm8UGvKoPJCoLSe0
ih+hC1hu3Oy5bHRphfKZstGW6tUa+n0OIYgJTdJ4R/DkQwSi+PWJ/lJEZnv0LAI8
CsuPwJxxOtTw5XefB8qvoLmo8WMGfQA5+dzf9MTafBkIjls4EkEymo4/lW25QByE
I5TE6+AT9EPbXbEnpoBLY+A9JXOoxtkXmKcqd8UDIyiQ/xdDO0Bc2qWgyyUBQAum
61x/6sWXS1uHHr2Zky0D7CbXsaEBAREbeu2MIysUz+58u5a40ljFMDTyfvAyKgtv
x6DCPrzhotaFNX7ybP1R5dHhelcfqGbXHh9TD+ZraX0BvJ6rarS6nbDx3o5J2ZJz
6OlgT2xWPYgc2N2gaPOhdZoUQouTnu97tdY0G5eZeS5yEX/vlkgTMIJuT76lFrkM
8qoyMz3YOFQohXCL57QrmCjIHonGvcN16JOqR/9NrEZVmZ4CvW2Pc+nxIBCoXJrT
gRR4hPbc6kqIkDurlo92lPi8OmaJ3uFlivvKh9CpLGdwildl0K+xyREVxgIsOAHf
ZhtpTXL1/zXbrvaBa/5ewQs2q5OaMX1IFJkuqdd5qAx8jYWVDs6uds5Am6B0YgqF
iE7vd9QCvd80NXBEdTT99CEWBTufULfDCUB/aVqqQ4HcjKkko9fsYuuRvvyrNQ2I
ofdMXGDziINHsQGwdiltn3lj3rKmovaBQt8tkx49JJg0ai5nuTozQW5NxHehLfNi
uDu7XXF3mPO1iYIksKmiXQT0jGjftsqUkjrqzNgwzCAMjmgJtJikpubaks5nIHZi
qRS/cJy4gW5PLhn56SDywnwF6HXSTdvWf98RzxPzJ99dVS8J5/cBXGXouQmbn3mg
75R22S3P3bN1CASqyCmaIFPNPG9Va6Sr3ligOBblWJovqok2t2C/VZAqZAlmuu7l
xWPZwlSqVkmo+CE90/FjmF3dZCvQW/cBswFXd4f6JMfEjI9fi7PrLgr/ciB7DvED
6GyEJiDnzbGIQlqrQlraF71xC2OVU2+QZTGMdNGw+VSL9gAkU9v9yJ7do9QjX2xp
XsxC6WGki++8APs+rNSaFE9u/ewnZQAWnyHHofmfyKiCIhDBWhXwl/PtD31AoKA5
ivcj0zo/tDkv3qLxEhc8OktoAbyXx6RsFe8dqHD/7nyLIT4WGTx0wltI4S6Hpna0
k/ixuzfXa7NSGd+Ig79gkdxc7D2F7PfRTQkK8t183dYayoB49oK5aQqyZEgSdYJW
G8MKUq4bn0abgiP7uad6e2OZxIYhaVn7cwZcMf+AfAVHBFZCdXmFyXY41L5c4H2I
HP3PbyeGWi1ijdaF/jrhqxCmMhNwexVn7G92ndLJQUuSeCavTMl6KPJ3tQZJxMAt
siuYLwqz9DvHi/fi+ml3bA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
J/V9P0SVHJFKEcYEMbvQhfmoR7EaL8jcw1cQsONOaCk+cWfPKDxm+nc6F4Ilp0EM
qhlA3wZzANcOAiZh9MUsnGjIcsgjat2m1rr/EF8k/PYf7ATYMvcWOM7h9af02eMs
zWPN4tJfqkmeBxVTIcbTHScE0vBG5mcG5vdrF0rvepEvm81ZcBJmSE2keRm0OZKB
g9mqbcZQKymyFmGtq54/rMvONiC8uFH3vjIQRvCAa+lQPGSr876a1/QWdj+jZUuZ
zla/LNhoLVA4QPKu7lz4Elrl0IGN38m4cRIz9ACNjEJSfJloHdb8XWetC93ZvT0g
qO7gCs0Ha3rCM+kzq/Uz1A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2624 )
`pragma protect data_block
ylh0uyM3THlR7DPIIRFiFshKd1Vn/u/FgC0gEL0VlitZzJxVPHN8ht4izyJq3b5T
SNp5qmdUb4TYrMXOz3CW5nUVrEV+gfOYS+BF/OdDijz6AjHdH3wnZMCgW8w8596E
MuOpDNxgbPOXPPV1Qzax8GB43bvZJqMhn3CL/ZO6fQw6GxaS4rAasEvxaVkL6uDW
qjUSwfQL+4u3WqxtKopZymCjtosg/uJWS0jhMoKYVLq5zVMyWBX+506pUCUgxwTe
CU/HD+FD3Lb5brnO0iiXsHqYLZoNkhESPYu4gv9fyWXvWXTR1dwwmiKqM/2kxWpO
hucDp04gwZ0q3Z7yQMJrOuuQzFMzG60PR7+JBk2YUA/kVtDORhMz3eSzd72Lx7Ek
z3yLzJ6NCzk0wPxbX1xUeX77aUWFSIy8SD2ggVwOP2ZJYTD2QlbsPq6VYYRv5IRQ
ROQwlMGzoQuscx4Ip74ixbWjI8TPCH+kAI1ucN8e9130nmcY27A/7DdgmPv9ftK9
VOofK17/zG/NgTJtE5lmhF7OGtSmWoFZk0w1o5U7HVEWlELbnJK47lCnbQq1MvMW
7cHTun7tnHkuOvbdPSZTt7OsFE3vlk+4JtMI117A6UE0laQWxSOmFYCCqgUdWQtM
EeNW5G5wxarBDVojD3EntnOoox0uBm4e+0ZUS7JByp+/XAx7PaAvZbymdZ2lYjjO
L0y5mdi6xGxe3ztKC92gjtnNZsmZVVruBOAM218b70827ntx4mtYr418WQJkvdHy
v8PN3YR24SXVIERzuzforHzC75jYugvJDgQJJCa5yxNVY3B0zSpZR7MLNQKQ4lca
EWvoEdFBXzlqMeL7bZNcYteN9PFTq5XPVcnMtDuhOWBpYnCL1bs+YY1L0MKJW4xd
VbinP2O1RJHQMp75Nfnxt5evQABFfh/WTgx9YaZfutPSa69B6m0B3iK8wppGoBOl
qTWD9TTo430LncHHUCQRYxiFe343dcWYupCDpvE+lbxlYSvkkAloNNleuJoZD1aS
2TNYAGkXY3VHaJ2pNPYh5n0GLEgLHNrtTLAAQQPasRfxeNb8aalS+hNF8q7E0Waf
d3KsEs7asSZdr1jz06UZdifGzhd3cwf6P4MU4NqLxjcnyMaXrkEPk6nF1DrTokw0
SAy2f0W4AZ42wD8jc7ozKAf7qS6+J/jbiDX5k8ltDXbb2VuAbVDOM+Y4q+4wEIa9
cDLiv5x0ADxHJOn6RK6Dt73+veiz2h+FSx9W4WwnxxDdgH0hCbKK2Gy9/39Ze1fh
70hRCPzpncFd0i0gXpZD55O7N6bedarZuERyw16LIaUGGoiLtI5rQTDwCIwYR6Oa
qHM7YINNTaUn1AvzcxpOLzhwZjQGbOdWUYOtKW+eRkU571RjA+IDs0NyfPbPBwW6
VjxaGQPJaibqITicwaNBOtkT6GlNuC6qynhndfQk8FThtLu9Pivx0pQAZz7+L93A
RcqzUrnZqI7gzH16tuMsRGEo/xNE+a1mJAb1rZ9kNdBmjO0eFtHjNnVBLfCQdyZn
+HXg+hBUNC8tXcAX8DYfroW8wF3PjFymaEF4uv4PLel9tTBhGly9SH7dIIV6yFb5
vkrQjTZOAll+2j/oVYr9H/9sxqEUzbW1O9ebhtWwYHxVgV1RzO73foB0IVdoQBJb
l3EWr6XBNLKDjhqvCFSxaXLefVdnOgZCa8/92vBfe//sJlox0fNvDUimu1tQLaAY
YqSjNNh6ojuPGioCZuk7/t4mDTwb2/vTaj4mzRuyWZ4WmCWlIzmBrHQLbz9+EEwS
krVR5qmFkYhPKDAqzZG8ZjXh9t6j/fTAFIkAD67le23PERyfFCBIbbo/AhTU5uMD
yBz1yKhkihLSxXUbaPiu4viV/X+fL49LKOJLVCB/REVY2E92efuzD8zCrwjnmmOv
ypun8eYrky4jvqGeP/t2Gl7f3TJau8mHGR+fnl1BAeK20AroQYX4w/rnkDU+jfZe
pE7bgxXpbK0OiovU9uAH4eaJ+qlM5JGd39WSlvwPUEtEcNcjJN0CC4fwtyHwXX8M
NkH92n7pUmjJ5OEd870gvoxXJJlJibCaGthiCEqBHGp9toQsg+UWZRoJ9CoQN1tc
dC5/LSddNcCVsi9H5UVtgWteFD1bHdvbwAA5Ow0LQyncccY8ruRcrD0E+37C323a
SBwbEu/tPk+QjqVIYkoPvVLjazB3AoppnK9P/BuPjq+naae6sw2nn2aUpUz9q3MD
n4t7wK8Eh55qQDFhP/mxtKawsUWSvV66/Ir984JHWZukWYzAL6aFhOJWrqnZtdgU
YWV5j1M/pf4sIGXko2UnQHTg//0AIiEZWMaT574+mAvW+alZtE2MmHpcynuUKCbJ
g5DcdMLx8/QsyE6dzU81VrSVCGogvFU0bSo7hSszX+bfnBD3XWykM+QXRcxvq9hj
vkyWzKQLcCh3N2rT8AAyvRwIwCgi56I7KEpt0Q+dM4N7W0bEhiCpiZ2IMfZHcOi4
3k7jJEW3bfiIFn34WLUrUruu8s29OYvUrkgxNRPXgskqw6dQ/AcwIJ1mUAAALNBY
LLP6IMfbGozTcK/AuTDQ+M7/tLrDkUoCt39j8Zlub7PP1n6EDlT0QbrQrjidzm+1
HBj952KhK1Zou2Z2VcvIraAfKvsCUVJPHM9S/6+JMogZn2K2dMIfzJgF4wBoigTK
cA9xnrdFbRfOH7Fkvn7efZxUXPFKINfSpnCs4BiUlvYrfLmdUHySGXnW7oGdjuUE
m073wdCMhKvkAi3dE2FOUXUI1LIx8+DLoiILai36SQcf01gLyGwFMwhNmyT8xtAt
MGmWOov5L1InhQrn/mEJQXjpjJZRnCKoNXAPlXShuXRx6fe38YqifAzIEEHDjn+Q
BzWhKzWZ9WxWTMXgJ0ixejxciSbPLNlHQqwgGiHMgXCN7KQrT9SzVt3YHrm7xlra
4QQyvRUWOVzKf6y6K2CZXT4RbxDqTjdSxjo22DE0L+/6rXkC2xFZE9FMzV9bqHOG
s9r5plb58vAiYR98yA0hxLEin9e7FmoiWG2gdxdMsdbQExwpYgyW8fpz9Tu69he/
MUtxpaeqy7PtYCkVzOzJTvHtqEADnuUAmDv9k0acnLkrxXpJtg71UXJ30oWJVW7/
q803uvrOV/PvX/2RR7+cgqefr4D6DZ0ygde9qtFX4PK4BEpZ5duL9W69cBJ1G5Xe
QA8X35ygk+3zYxZh2KWDClA/n7kpNLn/ZpK2s8bfLfib0vTDGn+qM9vLfanbg1vw
pTsYsRatRtdFTzR+f5zPlbnTjtNyzOGFYaLk1NZBORQBBN1OknyyxYrohfL6utHf
BGt3T25D3fIgmHwHzpcnC1FQ/3XpLsKwbH2L3XabyyG6lHXUt0iVtzDsgQiNnOa/
rYP1KVYedUNnVerinoD8utoUR1MUup72kTFuEe3BYuI3mz3ET+FJEawCauiIoGki
ACkjIXfdGJ5Hi1Fy7ePr45Qfi6nDqxXriLqEtN8H/1o=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HUpYHoEVwod1bJSs6bzb2+/+yTw9yvpnIStqTkQIEK74Dia+/cY+gCIQm0b0kZT0
XfvCqpIjz6IG0DInTCSitJMNSxtC9ZAnKvVqy6VouZ2naUeCIZH6Pp+KzJL//VSM
Tgev3PF+57vB0O51NIaH6wQosdmSEwHb8cvlmiAlI7yOF1HeDeOIQ1B8SQdoch0m
EqPOl+KKP20rXXWX4g59+M5DUdj9f9nMB3tHcwqhv12P+TkQnJYs0dcqDfV6tegs
CJQKm/oSxZPTY46Yuy0BeVpC2I096KDRoVK0h7Jl3OG7aVVDfvYsY3J4qNqK8iJc
ccxxBOGwam237ze2v+U1TA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 17824 )
`pragma protect data_block
eGvuVEsjKM2uz6k4lrx2eQ6RsoEy48W2IBBVQaP56QcPa/FnAQLnC1hSmWSZM0GS
uq+cjMyWGY84/nuCgKso4TmzZNKYSZJodE2spLYMJSk1dAakbAv+9EidjSsEt1DY
PCvQ5Y1Vc5Gt1bFALudtZ0Jtmu9u9t1at59UxqVerBBpInj2FeRphm1a/fTKdl8P
Ywr+8t9MdRzK0qHNph8EW5Ga6/gilStizcMUOVHTElAKrBRsVxLGjSBWqUXf3dsE
GI129LscgR1ZGEWa2N31hvkMZ3oHDxpJziVlXmSJJUCUQPFhyV7OBzKHjZi7x/dQ
tFurMg7OQ5vwbYLBxavM8UEAl9pJoxawIQV8BR3F/WXrgZ6Ii8BxyO4qJzgtRAMf
qOV4zhWt1TP+CqOEHolypYkqW+4BGEwECkJef2T5tyPSwsU4D8jiWNm44KU5fwT/
6+jHWf/puNQAmq6z/dqwvjzJo00dq683K2hA/pBoh5O2pc95Rbpi/dw6VyaC77al
CA8PLs5NMuBRONtwzFJMEJ7XaUfmfShApVJImohZS/uxwGOEqdK7h6UORJ1rr0Wz
IUT06OHr1+JdgZPUgtT5NBfLEE5sXt6AxxPmUl4Pzhj3AgRhXn58qgg8crjpfwMZ
L7aKSN57NNLB6kIs8FMmutscf7ukUv4vMOfjdMkmrqREdg5nkzGBlhktSw+via2B
D8y87aWbBcSuoVDaWV/DFrp4Q+KXgX3Pp6eolaLrj2fchBWATiHMQ0xsMl8MRdGc
OpjfLRUXLuYBjQg9ufcroQrnh59ufqNtkltFCTJFY7piuVuJ+wg5vSd3IbLnHAnK
dX4ClnoGaXDlVPTKNgIWLz+J5p2Q8DjEPOHWjUilfF4KxxqFMKUV31Odu0j1GLDz
KhNCrEqfQTFuR9vF3wEEi5zRDIZaws9G0LNV4wBhhfk23jXQ2MWDQEGsCQWpzIF3
f+a6zltaRFiaNDuHR+6uJmwTi67sMKa0YLEOqxR94J3EbUZCLDSTaWxyInkw7BhI
hccRXSH/yLZcF7uF/YA6f42EalqgudEa87xK8n4J/WFgAnspzEdck3TqrlcB4CYz
GzgSLaTnWALkb1Qd+h6/oGa7O6m/8pT29+N3+EH6O687EYcpwd6upab/wA/qn/rI
aiqF0mRQMBty+L35ssH3ozG6BZfERF0FQC+QdSSWayvpBSDbXUcxVItF7acnQa6z
lhWBTVOK2TEw9DaZljTHBJ2vqMXUxRdout8NC5c6uC/a4KRxpaP0VewZC/Plp2fl
gJ4k5Qd11+TuqItXyv2BQxrgSoPcKmHB3esJOXsGYamntv/u+LdytJSwa+LN9Lz5
Av2s/Mxml4gDVDsgigUQlpcHYIIQUgU6fpMkuOrZscArCcHZ4tlWeuWwMbKpFf3p
i01Mvn4bloCn57WBMEPSi1bWfwJno1NsdQuE3zuP3XbwtqfhHIwNiAw9bmSaKEhq
E/nU+HQacGnF67QAL7TbM9V8BB0WTVHQchwQDYCJqpRfacjoGSzlk3D2OnThfG+I
Ut3Jzik4hSmw76TG8XP3IXFF1iGZXBSAd0rXxayMRBEz/SzE+9snOlIRmFYo7GL9
5DeiEjnlQmCHTQD7HF3IZ4E9tR+zH3YNYmQLUMoBNN260pGprVWDDswNS5Bq+ted
ab1by0ztljddvynn0IAtRa5Iyv6mebAtLIOpD15Y+MDIeyZeKBfffELoDnWoZ8WC
lX3puRHYXJvrzG0p+ZwjgEvU/UlOe/jQEIvrie339qJBa7JeiqOwXdEflzVC9gy4
ns+zfkKDEoryJjX/FJjCbU9apBzh+uizhBQ41NdKh2n8hc3CJXQnrhaW9XoRLwVk
MuzE2QAahMvs0sh9bh3ta316IXIP5Bc3FMPyoDy3Xj1yJFJjD1yEWMeXu4yvRBT5
PdR7FWWA8gYOXwI/tYg7LSJmmWrC8S+II57y3UrNfdEyNWwtq82J+Cas3sKOfSQa
rM2j07Uz+5hvbXO2hpeYMx/AV76NKI/0x4iM/EsdI2yLVwNA2ywYj4j+YqBargr1
AwrLYdeP1KjVtBeC7jRRSwrU/fSilt2r4/rnPxZiJtQzxFJrQOFnlwB5E6n+eTAT
uYtpXgiGunuJQxUrfYJ+dCEhYxA8aNaBzxvvXhp1V5DyddwPRqujJiFUUkBJv2jR
U9nwzpZE8rgIu24PhTSUKhszsFuTzMROdcDaeMKSePWfD1Wu8wm5a0mF9wE5oz/p
XmLS3wIH4YiX8BuPUHNjzDJlrsHhEaz0v9wkMrYNmtDG6KpFowntW7pHw6e/2jOA
cX+iX9lzXS9Hk10v2ci31d9d+JNyPihalGFyHY7EmrZW0qgskatisAxaCUcxY+UN
saSh//NU1z5G1PFuMw0CVXOyQqhTMOPOoFvn/8gZNcbHjiYffeHzPivH24IfbokZ
Xuj77QWrR5k2ki0x3C4DFpPQvhWu6d7ptY22Z5aUWTPqbUm3adldzirFkGhSluXX
61Pms1K8dJWD0tZmLhuCoybPKZE9s2eMa6l9OsKEAc1YqpoWtQXNtRz0W5If0FEV
o6+kTR22UocDuOYsBSz+XBK+TeKNm8g89wKMC8oQeBm7JgxPaRdF399+YuzRD5yo
Z8WGLvRm7XrNPYUozeMu97CdeJASbkqfJWYxvoiRNcsYPx9aZIiG1aVt0RQJxdMe
tSOL9NkY0cRbxXmiK4ZN8W2xaaljwDpmGzuoGQNHk51En2nK307rcOzOxaNSQqWg
i3KiHh98CZ+0GdhemWpxlbZIGS0+5zuvA/gG4wEJEG4BG1NmVnmMj/3LbaX43Mc7
OWARyUvNMsvisP0tUB8yhStkJCYOG0ZuVXYhZBrOSuOirmoIMSP88uCt0oHZl78O
7kCxm6Sd5OW6f89d41aStLLs6vQkT3u5RX1D2HilgpsV8HaC6DxN7a/AQTSwbQ5Y
OsSlLmhon+1dbTQi+7RM7YKLQjDVBKD4HIAGVo0Lmxcenwd8KsXO7YOKAPfn7gjA
JrYveievq2CgCXef6/jato6CThIT/lzxwdVV1RRJfIivJveusmDyNrWPiJZTWZhR
EJ/2Tsg0O0suwnTFindDpwaSaMJi2UByaPpoTmgiMYgfk4TV3Anq6Jy0ws+z9K1V
SxFwxWIT/Ktvpu4GYdqu5WTeZwCOVsO/1F3888yKkqPwOCr0ArG3G3WQrsMuXKth
7nYXSOBzAZsEVl5LsnNOnvMgp23tTjBnEKYqxBGMygvBY2nLWl3gTlqiMGSpknWD
AnsRx89VL36gC30QsZTpkw3qB5RDgEJyfs1LgJrvcpjLEUddKLpIg+Ssb0sW0u9f
Voyv2a5LSVgaUElPQb0RQZBBAfrgg6upb3H8BtRcyeCa0PaS2jX6mdpJgvUx6ZxZ
fPgeJTp0p7wFuFlbpON9NVH4GxShZsufoTC9qD8HVNbRGfZXoWEtEFDRp4BJqFvk
7TKmzQ85IVPopygtFPUXQjI9teBXpJ+IeexZ+/BxBtSbRR4mPcWfFsGRiIjuf0dq
0DgQGZbzFJmRHaoRbFvHw4VdRWtUKCHCEB1DVxEFFank9ij9ag7+QTHeaM6GTk+E
d+kqTkbvieBWhmvCAVwW/2hCQYvhAS2C974QKyVvnjE6FltN5keuAGBb5dFcL25j
KZ+NCs2Ow1Flv8U3jP3GwI+mwp5FWZCMqIMnTSJU+qV3dPCYvSABYM7uYXamaEbf
KOOzoWYcaQb0ZPhIiOcQhTQra9d0m/JIyCPcr09+MbGyzky/esUHsQ8ZSnh+xCCN
L5BzCDy9eKc5dP08pY899QTypza/Haps4HiWx85g4LIJGfoGqFgomdMZHBpKOmn9
vKjdx0V3je4MowH2isQak/39AEIAAQ+rQvOKZa/XgRkfUKOf6uDe8rLMXmp0qJPp
Cmphhi6ZrFgdde6Wloe1xnNw3MwGr+bBmVCiFZT8RrqWyP/3AhUi2GIxYwd5+ojb
7/RRK986RME30i5lu8byDwGGAg+ilTD4SpE1Co4l7rYFYoXNlzYO3l7m4mX8D6Ti
tLdGKfDNnWLpSIq4VpUBcRkQBoBJIB46IIUBh45eAAFmYzsscpslRVW9cMjsNVIL
am/aMNdq3nlfZv4MbLndBlaLChcaiPpu6p5nQ0d2Ga+UY3dPlxpxDIan+sgs7GWG
XtK1z39iQtSP57OuymdOS3sgmHyNCkKbXJhr5i7BLz8+9zIwXvHX+BW0bOwzfbTp
ltxIWiKI9y2wBRJNHWN5zWr3D36G3TcWrZPU4DL0JFqB6VUtt0+h4vhTs1ggVoQp
BtFKKLVOEf0kI7UPuZWJ0CQ5jq6s2gclCSrdbT7bhABUAa3fjpcVD+P6ATHslwmo
hU1Gs4UuYphAsa3EELhEIKGnqTkuXCoilbHDksdqrczmH9ZFAuRsTqZP/48MNCmY
5L1t3dafSAePqm85pnkXTPxuI6fI9IVmJUksvNZ8V0NkPCxbWCNeDWrOGpEy2J6Y
ORlKdYjcYR6uoGbdVhnZCixOBCmMlilUQGtEZAJLB+BEzgybEfmQeGG8b/rlUb08
/Ij4hwxwPWp9vgYnz0+hZ9ksOb/2Vj2kMHyf9TVAR4SNpsbtY3925t1EMdHbY3x7
swJK714vv/veYvb9O6UtBv0T9ZkPuNLfbA5Rfp9SMxf8lbYxaKWIixSgM225DK7j
hzYIaPmmgKgzSS5d6EJ9uIC8gVbub0rVnpAlNFqRBZVKTiJsdh2xXrkAUrwEcYYW
TS3bvseRTrH7x9qQ5OE8zvr+wzXqbyT8H139vViA+1gBcjh1hl3VD4I0rmB48Hiu
cB2tt80HLaXkSsDsHd8A+X7cm+bEIq0l9XUBIyL28ySWw7uGilvWpN9BpSb0K1th
iJcMssAxRXSGEkhUnzsp0URUpXZNzgw7aRxgXqxI5GjG5Z9AjB5SLwhrzG7QV9JX
RfJbt459YawT5NTKt9hSZpOwdAyArOe9k5LUmV8s8aGBz4qACojZq1VYQWWUOQal
4af96/nDvukDNdc/QqIQK4RWnQ3qwRwJuZPHjWJETVzlWoC3S/d24aXZShqD1a+O
TfzJzFEaC9+maizwgQ2VviROyZnL84fihmgQVSrDJJBgdUNwIj409kG6T1U18CCt
ESSug05N5qsq3RIw6Q2ydmW9Npfc0m7xNPKwQPIQPOv5+usmFB1WWyE1a25BxlYj
UAPtwVEW+ZjE6zjO095DdgSW7BtvmQ1YxTRo/JwsTmjqY/XfISygxjZWyL88zhT1
/4enC60E04DPyAoqnO6qf/8qS7t8TK+VROpa1Zfuz4sEuS/Uaw+WJSOyCousVLI+
NRH8ULqoEYWmfAUdqK19AVTILJiRaI5LQ7ZjZ/3S4XOr8HWiA3RaoJRBGkEU1SlO
5/sUQW3xArqybgSy77md1bXhlBa+G1MQEd7GcEL6fC9KtFL3uYWKIN0qDZ3dJBPu
h9wkoF18tfpIZqwOPqt+FEnjrFzLL+SB8DL96LCfZpgaS+m72CWtjtSjfJfkA25y
zaygjMJV7XlQ/Amvc/CcbwvLGZRT6YkgCGX+PlfUItXV22HBq0BfmCP7YP+tBzrq
YpDArwjSM63xJsMbrY1t+H4PyeL5kVn4HGG0rvY+Fl3cm2E4FB7aLXBzweHncNEQ
rR6FlZdJnJZEImchzl4KLR7dROT9U4qviXEBHLct227gFsjBDpaxSUGQt512rBJh
COIAwxEFzOMIOj7nLWtvVmoNqBuwpF9ekvfDYLr7kvIKQLSIhApJEyEL1/3XtMCX
sp9BlY7/39CaqDUnahUMuX81Mzdo/BxTmlYb1yEpi718u+nCTvjIhzkR1DelB1vk
mTo/QQNcv27HvYdhV+MAR9YX0xxj/ZoSLxvwNVwIGgewYqL0arnX3cWxrj9jRPL9
JcA7Cc2nR16ie+M/z1dn7Jlv4Tp84iEI0kK7Trm4knpLEJOQeHmkfqSgDvAadbzk
HFhuqHJqiYBExBr7TqVxQhIIxRGHc7cWm/AnA5ujG6IYOd7abZwymftB6YsxZe61
uI2gHSdBbss1okn3vMctJbMvexvCKyYETMNEtpcmr3lz2x7aPwp41IsklRI8shyM
pY15QINmA0++yA+w+PxG5vM0ztZLqIWIkOMZjS49KrdiL13afR0EQ0ad8Q07tu/V
bHha1QG9S2jg1LAOzndIPfYSBeCAaYC6lepkhqX6OMe6u2vTZueLYx07K5xqEVkn
TSPmcRMN62MJCCpns2Fk7UMzROtDazDTEjKRLoI7ETfsEC8hlrNrYEWglbD4Wm35
CfVbD/4492s2F4t7l5GStDx2aApebsc0v0J1q1RNPXchxDv9ZbBdP0Qe23kVYnEi
sUsSFeKE3ZixaTLPo7aP8nfhhPv2InESz6aTfDH2N/G7HucJaXsUCaMCmP49HVFj
ucjPxr8Och2vLTpDlXFK7D4y9pCIQV0BVJJHLn01yFyPfRR396DBSruz1h42GLO0
4HWHAJRwqTI7OOXT8EQf5a9mEAezipyEKRFh+Jy3zllyMU017LKnFHmAGS/10KFn
hIiR/dfvr1pwwBRgZARcXQKy5xQn+hHQ391pODjeAXb64ZgyJwW+dCfjwjXby/sE
zsHEqs/EhSH9IHVIWXOvZXu4Bllmb9miIYcqjj/2+vNUnCLM5axdPVI1YpjRhgwk
JI7+iztwshuVjhGoFbSQnhLtR3/xt0CrweRzV5bzdQOr3e206xmKJD14O1L5cHLN
JVkp93Qy09jMKZnMo3MfdKZHon5Fv7+dDFp52SnjLnmPX40Twyh4wxYLPqUb9CCi
Nj2DVJWv0qeSDSlaopUQsvJ7ALqbD/h9Pr3Tw6jSCo5+jxtH3f8O8U9U8+TD0DOr
g1y73PiMD92mnxInl32RS3hMlrpFySZYXZZTKu3HDe9cFEJ1YtjcnDulpn7MrlFq
zcA4FL4aNezj2gt7nch8+KvK6kWZolOYZYcJCfmUj8otPf/Ko/A4L6o8lIlPqUHJ
cJdVGbTGgecAMM7IJtVhLdFNWYxLGW09XtOSOwDCgipGgb4n43CdyWex3O5YfkuV
vIzfiSlSVfL9Xz1hkB+2hfrmZqnDhQs6Dh/JjR5yA9/Yv1k8g0XMpXMPb/1IWxvf
jAuCxutBG+PFlbgblkK9/U8Nhi9bOxRTEiywjvtryoaQl61RpRb560Pc6F25gsJL
Wj2XHEFb42SZpWIl+rHLj80TEskjx/7nFBtck9kE9L/vnDjnO06oLWR+dc56iZ24
A55kk67BHFayrgZnJ62JgHn/SmUnpT26s+fzwhUl/BnHJ6KpHzIyYTER6iJKNwVy
JCR0SGmC1eXm6lUvtvxG9ep7uicOTEW2I5hi3LtW5oScFsS8yhAJ3DvRkGmg5HI5
h//b2JlLP2zyZ8ADsrlVMneMf/ZAr76HPLo/IEZMTQDmYpmV9q+5mVAnCV/8VTCY
Yj4o29r02aT2fjhYrURs2DXLILJY/717vDf3ufolz4slUpoqHWTpkLmQuO+NcSet
EYjX44dvHS0wdDV3FJ92FUQeQUkSXBmPoUUYKweHgk+mqWJw4tF0kAVA4vlcui5J
aJ/1s+5nPZXLZEGlLatQ8j84VqG+XtwDtIlD0dNIK4281HQfo7Ue8itluq66frTC
RiX0au7uMZVpMo28wurwF1SRUyTagp5G+8BnP7v6yhkUj8vlNd3d1ywFtlntAt1Z
wzQL1VFYzo6V0dVu8mzNvwvPkRc/Rk9mKt9E+RMpUO9sJbIMqlD2aeM2EyAHd+Mx
hg9CBxik3K3b75fwquVe9fKKzZKXAxDKg73CWIu1uesc4I8FBZH83AxkAGOCINQN
P56Mme1vZq+5om72kp/Zao9IZR78degjYEnWG0CS1/Z/Z3aaT3i+bTSjWnoouzwu
ihQh22upszrWiOyDUq939cl7c4R8GM9IZr4qzk6cBNP61CjYyenuO8MLaqHwZ5lW
oONhOVMN2OItp0BtfzPvQhk0iVRH3CNvfKsl/dA/K6dEOLZmzl4ra2gcmTlQn+bk
Y2jPxV/+V6K5nSDcYZOR6LC3b7zXhGAUQXLQunYhGGtDtkCakert9QzBoqGe3MC6
Csnboi+ava71ptnGK2eS9ZUe9/KSf83OByfJdPSYWwVOe3seBRQJNSnx9joRG7rU
b06i2BbeHSF9lzkhvCEDWGyNEOJcvDJqmvjms1vg+I0WbT0aiqUppQMB50f4BKr6
xm81PsWbHtQRgEzGA5x5OHHsy+gjzQSReXJ9KrCEigUgebRwWxqqpdG7IH0GSuVs
20FIGPNcXVFr8UiA/XYRT9JU4k51QCf48dljUMkpF7WxxdVmEEPMQsc/wILxUjt8
NQfMMlIBeeYG1wNKJKsAzcv3DTmYYlWT7FR/1moheTd6JTC1kgO/1g1VqhhZj2HF
cgthhRhLgcTiGH1KLPrBOSqut4YZQgNRUkiNst3OaGqmATXV7d4fwvzP7v7+Jq1C
Lg22/3MmVhc4NBow4pyL0qXcdq1jqVF1Rw61SbuBdu4Up9YxvZGHsMKvEIvJKBap
5pb7POcnpEUsc8gtcL42kIMaeMD62sI4g7E8OY6b4XU9p9IXJr8q43ExzgJMv3bO
LrWIuLRZbhw0Ux3KzISKl2OplQ2Q37cUanhk90DYr1tjFc8l4qvzRXJsaX+loC/A
WF6NPGuKOSOWurWMvzcQj7NqZ5yJsOCg5fXCaHrawy6AgAFQD75xxJH824B5rGq4
sgg9obnyD3R7Xkx9xPuAxPFBX5uiWcVUoPXYf0IyxehRPZYpVB2iZi3Tk1Y6IhLB
Kg0qc5VIuZiVy5x9Y22qErBx1/r1b67oIObFXgQh4ZCEDW8kYEl9d2mkLYyY+Api
MoDYod12207haFhI8kOF5ssZLvcUTyZuWw6RMdSt+ndC1g+bhG0OEAicrH2rAE4R
/fYKMvQpj0hpYyKIZmP/jWfGtdDnU4fUMif3Z47cxYHMJxl3rhMuWKZzA9SWamMo
lKhyMirT10y6GM7joEhvFgdiD3t6SBva9wUOXT+ZYPhX9Oss9z1erv/D2mML1DnA
shlaNHVuTiJrcQdzIMKTAD2iGKgKGXan/wl8SJtoYbHPvk80sAgdRV46avcgR4gf
DvpJm0x+YBamXitYq2y2qX9dgS05cJvEvJlnx7oK6ZgK26MLvXRvkbyqWa/u6I3H
2azyy5Abm/KtVV7gKcOhl3Pu3uYj3yprKijZA9d+sb52oMK1xD+srcVH5ke/eq1J
KSYnXm66uo7S8gxM5dSFsiBiFrbReiTHktPjl/vlzPdS8HdGs/BCeWZeNwntDr5b
AL1a3P5CLAFZknqGBK5chglgkz9h2M+R/fcuE8tWbhhEuvlTYJqrgHN2/v1EW3cn
i1E4EsBZMafcPGq/FYyPSKq6kuZ0zNiA7DvFeVw6uPOpxFFk1xVeUmIyZoOJB970
PKtcfuHRC0+OW5RPTUATivx0N7gy/IOD5qPdIhsFRLjk0xI33+fus1zQ7WyfASWv
5vrW09l/C/Y8/1f7Ph1I365MGpeK0xgmBSUpjT1WtivbD5KfG0Ep5zUPj6rLLJiX
QmuK46MpDlCeS0L2pbeqNr02faFh4uVnwPDuTU/CF5ZFLtBHmsaugh16CxLTfdh/
JOuNZ6F+dOo5Tv2IfXGpWMSHMDHa4ayGF3ilCQ8pVpGE65R/9GIcOGzj4QsA1pml
/cB603YnDkwvajm3TqNLu2dLLDwSB3mvGSGM1AAPuq+HxVhfdHdJThhnYyb4NsDE
h396NpjP3DpbQ/YnItOTgekQRJzUkZVG/IIxJmTbyIweM+7yf8M2olFGzPwsiKRU
0pvIUTLDogYPM1lXVtG3BaO74L/C0dr5UKtd/clh3e/n0KHfDwabho+Buu+ijFWA
tPl61AsopcJedHfa909aKVuhxf4U9zZJJaDNwdCWfBkSyHp9wxSuGiU4mkd6w9dT
qQQYqMoRs66nmJ9+nuUoDsSwbCB5IyrF4wtZhMTcySpOD1BxkkYjnrTNloRIhLW5
WIuUMczCrauNT9Pb37CsN1qyPHbmMdpolXZ//vrMTH5EUTTEzMrtA0RaqUP0mqp3
simAtr6lRUOUrJtg0YEZlM2Mb+LIk6v3TcS1zkmAXFWjkj7za6qDsa5Z3QtyASr6
/jbIC0A+G4uNWOeCJsLnMTsSDpZa1ByDuO16NW79H8YtoIxeyT/VsgKwio47cUI3
4QHt9LT7GQUtcdd9QDutTQI90pDVJk47FdCqhifGoheKQrBNAZC/rBJthnG5TK12
aP/ZM0kox1OOZSQVQNIJU4aWGVenAZdeaNkHqhkZnbJdzFAkzZz8a6rskjp3E3eO
44KNZ6KyQN/Y3K8/HA9F6/zfkrwA6XNVD8ZggAAkgtWFHo6xzL6bVCgg56YF5rER
yXHTrCT8LHZTy9/dD6EnuCvnZGNFsba/IHwNl3sQNPXxvD0cdIv4CoCEDcd564NP
iEI3FH86tBVLNOd2S/2bcScBG16mpq7fBQcyTVDV5P6MuDQzzahn0zuFEQNDjphQ
dDT5oDLF+Vz6dH/bSfWTPpWH9gzyhipj5AMr0iNUW0AOvVOufn9is2us4osGEKj8
Qznj1kIFspyBYXhSH5I+cJNgULEJqLzmdHhgK9Ip6OyJAWgks0RgFA04Ah++PLhB
Y5TRIh3reBXel0WtsrXjt8eD+OIt4HuQ61uEJS8JvxTXv3a5bK4wXCiKSQFfyWye
+EMBC/O0vHnrJndROjMALaJ40Aewry4MD801beibVK95mOdlFTGKQY1mEbZblGc6
UFSjb7AihBuzuJNK8hOuQwCrU09UKnV0ZAdDlVVgX2sz2WY5rnCNyioZrVlMQaeK
IiceO04nJVs3p3BzaY5ErdjETVen6xuPpalha8n0ISxnTTp+oG8NThhdqTI//Jys
sFZiSJw76za8wOwoa2WzZOLTpYvBGJbCslrZ29w8cHT8GsyljlbWA90FXES56yDw
g1CE7i/Qv2+FKqMfEqukzZvay4U2rzITyIlh+SJa0bG3P2kW4xoNwocX1BDi9wgY
fk+hpU+7IwSe0ub0uj+lVNp6K0VuYUvERyyPCY5dD0PqBriDWO5ZY+wTfGKqCNMH
VIUWhEOpshYRVXwEqO1mHyNHoVj4Opv04Q5059aEXePqEf+0CkryH3DiuhmRcag0
YddH3skhbpl7UiTp/FpqKRqVfMuKdEr0PP/SVso3l+5dx16bXVetho937TRxiw5x
Dp/tL2xz7CRpNmp1wYKtyHkKXkidB3Pz2C47oVpP3UxGpRqFtBXP60JZ279+3dYs
IS3t3YXt4yGi5xKhxA/lFtR2nY7yQi35v7QIvs58c+P+Lqs24NZv71tXciWinDvS
ULbcfTyY0A+Ru03viWo6+kad22DO98mK9NsHwKhqR4OKV/1oxPWd70XLpC6N8uoH
h95Y+V+3WgSh9MxQSEOJOq+ZhYzM1tSrmgC6Js8WJiQtRFip2UyZapFynsx3YINY
5iWPjWwajdHI9CZa5AAloWTtA9UerepmM67/SAuB4tbJASlsfZiAkMucPcvnFlba
fjdKvhFnhZ1OI3LG56VJy8FKtGdf71TyacNM/HwmGHV6iMd3xeHH35TNV7kbi3Ot
7eostJ/DVhzkUyRzUenCKHZZS3nweUCkc6X3qOFKV+ADRkNA7bSZA/94XAeiH7Vq
Pxe5K555kkgTu+x+9jz6fCvU1BaQhs919/bniKGgTyFtr6o3//4NdDRXyAHsXnih
LMasktZcEG9Y3jY5TXg3zopyk7owiyWR5F6WjfbgWKFJZEiLJou4TefZUEqeMjaA
NUiggGRtPDTZP7RkE24NJMKxxMtEIDByD1xOcCSDa4SgF2MxyRKWPK7KqJY6dgno
fXT90qLLIKD9L9K9p+u+OgQ6ClRbw+d4I23jFqKRQhdIfadi0zro8PF4z0BOi9AZ
6y+vN9OBNrsuaMyfb6a+O8OHfUXnD0nbgnEychRPD7m4pZ9+kgeJRFvxHyzr0mZY
C1ualJT7qqw6eEG4TVuiYyAqdRNRF9qpQPQJQz1OmEuVib1c7elI3oGy+QbC0cMU
brn7+uBPRDSgdQxoC1/xe5ErlSeWxQ1XAFXsGQt3BAW1pvQGvibYZyYYBTD7cV6k
aXw3CpyatIYyUrG49yIbL9z4q2ekm++X0MBrjudHg/3MsAgORCvGjUREIX5/pQxb
90lEgLCNgpffY/QnSoh8+Ay+264VjPSCtr82E3a7vlE63Ku7jcCb7QSkqOMyvFcx
sAIkERADwYqcHKQwfdQQ2XC+LylFq1MZuee2zxl1maTFNBzfNEqjNyT+M6q1OL93
pH3X5k5tJThZGhRQn7HvtsqOiZc5l4XhH5+JYkTWTWBwDlsXT831oqmkH1z8m2/D
rDjDksMMzwb2mglq7CcNiAzuaNncFQ1/uRYU5/IQbxCrUrrUdkXPZyRuUy0RCyy7
ZiAjGwFnxT8sMroUBmrEv96OZgchYQgVqAwf1RBVp74FGTIz7QA6VH9dODbf86Zn
tiQKJzmXevoHyT3Y79YT4r+qZ4+JaWsFWN6FBwYiJGr/YtS0iCkmqIAn+KUSNcTL
BwNCmDLyLqw4te01HR10u2z1MCO6Vfxl2xyaN+rCOkx9sKZ6NYaf8jyBEFkHZgmR
FRjVdhRr2M8MVCZ399+ihqNrHi3o5nGzt8DINpmT5S4kA/bBhLj9ajVPhxLYzbeu
e1B12ZDAsna33AlUsIF8FVaNpGUuVPRVx6fnqH0Bt0z6hVdMmjER0NN4y2Z3UxGO
IjCMIwf7P9e5RXnfP/AFH+d+YwC1yhNrcIaguoM8b+MCZhnFrPMlB2t/WbQuoWM3
+clqMHJhPhg3lZYLxVBYS7KzH8UrhIkyFB/CH8uqe/Cf9bnejNIPlPKZw5X5SV3L
aUE/IazuvKYX82fDhoSndBeMY2YIQi4N5Whp4LCddCoggJfu+f19vPV+MahoqyBL
jsOgb+1Wi4NHXg1OXHatKQUJ9LGq+oyOiRYCc7FLqI9Ve2S7vQsWMA1jkL2XeDnG
sXgcSUqD6FAGs1f3E771dNP8IBjjc4G0Ktl0/NGbj8hBMSCV6JDkP2Xiz4pkEoi6
ZigjkKbDyJWpk+pzwT8Y+8xbenAyerpfI67/kKos4lzrDcq5fYacWpQwcVqXdhJQ
E7RznV0zM4qK5AdIKiha1WYBksGdoH+gtg1LgueC40gdlwR6DkvKN6S3scfhCsf8
WRv3YCzpR4hj+tOUguNeySHD5TV474/mUpGSpFF4p3MTKnRgBp0QAWgQeQKeJgbC
g4d2irH4UbQ3p7CsSgdSbzfhDGMbUOCCQ/Sa7IQU6sHF9R7SQUXZ9gsspv3ChDFL
flfJShHbQggRS709Q8/N0PaVRwG3MSq0tWF0vPyn6PwguYw6Nr/yMMBfW8o+Ogd+
rMpEwD/7WTv8+8/4Ygn+i7qCwF2pdLNIaSyIgkPMK8RyRlYgIS6Pbghw3Vj2/VLw
6/eKetvXBGLpR5MyNySY/y2ZYaITrY53FPw1CopwteT3BPg2Cw36Ra2KxGyjDZXT
fT2DiXtE4P0inPW0rd32E5oppC7t/vSyrg4D1eKq+qU4nS9grxACH9SuQf/WfIpZ
+w77h3WFK2wIqd8pNDxoltXIsjjFUE9wKyN0ifpGu5D0oADT/ztCPYJoLgvOFeSH
T71uDpCyGiLQMpVSCQ1CQ9L19CZJAK7LcQJu1wP6OD9GhgIw4MnW7SJynKKyC/Vc
CPPoVGDtV1DmRxBgtldCrMw5VB/t39hhdMSuPuBK0YpZnWlJgk6fVUl7h2CjR0Lr
Hvhmi+jlp3mWRXhxZzKtu2uWDYhDAzgudREEOtdtGgMqGjYYVq/SzXKm0w0rvl22
yHpQTEg+Iaf+zQaEG6G4T5M1DjA7xSRjDaunSq/Z9T7Kvw2wVqzqfMh+VUHJVx35
Lr2d3d8i61vNTt5iBny7FawbiZPGwGNJ9iJOr2LDdllkwngBam/6bA+sMsiCScDQ
ns7hDBGFhkcNY9ShSz46wMxdHJfjWNprLS+Kai6TS7RTzj4Ff/JllN3J7iDcLAg7
iPybGR5qCqSTYx4fr9CwOyHh3nCqJOP2LK009QjLvENNXPopX9F3fHphUnrU2vXU
wllrqLwODBtKD7SoL0HQB7NuVHiJv2LAoOUx9J4WUcR/ygU+5gza3q4rtcK9Kmq8
+N8Zi2xaJy5jGkJC7sBZm9g/Y9pzaK3LWTCoWUycqhGLd2rSXWnkbQvVW69HxDlL
kKwagokGgpX6wcQm1Z1VThq9X6BgOxaZusNr4igQgZrW0VOM9Xic0nyjFV8+Rqhp
g+uHpAdPfMSWDStxB9Mpsu9Ru8msipE0QdRHuW2AKnqo+8ME3H2hqbxScDL1zNDo
twf7zxPG631q1yQ7kX10LyNmSv3/W9ULvQKcoppS5wwqtifEFhvcGcScJMQkJyGh
OG51V4nLxn6TOMPSV5qkncRYp9XQTL4N9q8XksgX7lqyA3BFImYYF7TXWRgswK6p
qoEHDb4mUvmeGniWCWN0OHEJGvBd7406qWCmQ5x31SgZ8r3fJqIqNvE0+4g//T7D
zfPkzIHUJ1N4L2AvTa8coCQ2S6mxsWKLKVetsnH6lUvfGKGijf44Xg658nOE2aqQ
xfr6YywkW2iGseGxs4AtRi9DrJ9cXMMcKim+uErmBRx1dqgMNqhg6Om0n9IhFc5K
zVFVPZArLi3AXGG6bpbdjPQFDzeH/TqrrifCMVAr6xBWmKgjNGfoQ44ympySSTbG
inuD8mQnEP2ypHzkTSBmZcXnb782g91ao71qGxyKM0oGNyFErg8LTEYEycnsFBOK
FSuCQSy9b61lnrLbYh4Hf5morO9CCnuEb+dyTVWbzVnY/iNAsnJBr4p7Pusfbij0
7AFfUVdEVH6tzYd/h2fLjS7IogOtBW5pgttBS3vl9Z3IXK7XGJNEpNiw3PfW6RAu
fUjmljuyk34P3lCFfHGqeTnNcC1doiSIQXSeNqQFhhlqX/NtCaVgP6P9Tf0IzxMg
bDQ8BLFWCXWghZzk5r1zw3uA5aAXNLH/vuQyLz530A4P4cW7fBaqWsHmkjR71DvL
fgIRKULPUfKRSLhxw93mMEcewTKoDbPQxUUZXmtdJIczVLOYbuS1qu+JjTS+ZuHa
w4bfrcKqtqdFfxchlCNDkivXcGJbwsnaoNCASk7axQywgTEuTTsx2GKsJlJA5adv
1CaE0oSShqcYH3vFhkCqcBhgBizRSqgTyUECmfeR7FZzrjWpwpc+UuwWbdxMtm2B
NYWXHSloxOnaLdbf3SMwXBeNBVdKyNMxaZQjOYXhCDenu1iEYo51QZZ/CY16HaJn
qV9c7Q5vBkk4nZ7kANj34Lcr5FnuP5fEztO4u6SeMUAC2M7nJ2zDdLKvmvT5A8MJ
qyiDhikfcpMAXboVQF5fIaOJN6yTGGVPJWtpbbeZLY1Pr2SRYgktnpOGuoZfjPMk
mJEuL6P8qJCEqUMQvCW+CxDYkLrnqcCd7SDsN7QbbYWqDtfbCWElVJuZKMj7giiy
gUebZOcP5KXG1m3wNH/8j2xfcshDskhQIibvMrWLYlGH4w43Xkbq5iZrRQVf3zB8
D1gKElOfJm3ZBfBbC63XSXE6S/FdsUDYDFbQkaVCBbaxvJ4LiWhOz1lFi8nfP1rs
b4x1EyyOllHl66EFsTy9DCoKT8lO9MXLXU+Oa/T1e34fMTQJDJf8SEpg9ydUM8J5
SqTZucZbnmz9Eu+ybjWliGSC0pl3BYZzFJSiTDhLVWSbutjUDUmigKdyBd2g2lxw
2R8LAqadbaJVTfYpngn5I56BR8UJPRO+fhQ+arAAb7tgsmhklsj/raURf74Mo85t
emlOnjdos6UgVKyH51CJ6dSaZxDafDzVzw6GSKzneTie2iFpAod1OyRHLNpwV4aG
1/k1hBC5yI0B6EDBSWs+n75ry5bg6FExO0s2fv/DSPfw8DvNJoSX+U1xHgGtFa1B
DoS+MLPIzo4vy97CFjaMfdJ35tmgpUX6KCR6pa1LZu33ewf9mAAgXJqMWpANHGsg
FTUD8QPCGZN2mJ0UiFM9KGZQmXWTznPZEZGEUvQu1RJGPiB3mezpuZ/sY4NLaEim
Y9GfLdnHZPaecoI/6rXAU0ISLpqan4ffM/5TmDJZMcBhdaPdkuGmu+fCqKWrm+sb
jfqyH19THnwk2qF3cmmcpVcPazJeWfqEdRaqc9i+OjiqGFDeJ5cPcV0xA+BWb/Sg
U3XXHQnSGbyZsFMrEmtGB97Cmgjnc18w1GL97ZjL3bXYuj0etgL0o0AlnBbsNV10
qd5DpaDzH+ESuD01jl/QwhLCy1+XhTWCBy6uNF6NBKA+kbS55HzQ8Z5CVPzMF8at
DFiG+qxom3Yrnk/EZ0WJT918gJOzwVS8iNUljUzFexG3b+1S//WiB9LpNdRax0iF
8K8jz7jEoO04l0/DtBWlmjucusLk0GFeIY+64G5jCRHsL+eSP8AGgoHN5P+o3OrQ
W96GIoAba7fHcUUyo+6xGuz6WXCUpMy2ddBUUgRXf0VJk3Fm6xWeovmUB9xQ14Um
nxq6N5W6UGRkRXnFHmLSNjYFj/BEZIcQAr4jo1dnCNtJ3qITEYsU8sj2rYQrbnr8
mcZgTiGn3hquTvWyzzXV9K1fHW/P2rxRAvWHxrUxcH2vMKDItk3kISyiXiXmQQPw
IgoM/U3JtpzBKIWuF3KnckdZO/IpDKTnn5TlD3Z665XCnJSU7Idl5rZIXujoWF1z
a7NKk4CRAofQz0aLvUcx1nB/KfnuSe1kyokjmywzyBSPlINs8oBKwWMwYXnCfRiJ
2bx4ee59xBfnTnD8qa733T9i3C41PRP3kg+PejWjEE2zsC5ekgNoX90O3CTe75Mq
rxJ3dXMdSXWsqwFO5MlvxLQuoiNYQUYVpQu1sBUPEpNYqH+QLQP/l9p2p+uOPir5
4TDCvF4yhzU+T/lNY2s1oSHnWxNqJE5pWPwi1dGu2P3cdO3St8r7X3/hkTOmeGsO
MaOZoginpaZ9KOBwVWhGmKOMpB/bGal1inqJ5u8XhdEn2Al04cwwqCf5xf8ba5jP
NVicGyrG7hgT6nu1VEuuxHJ/oL+b/JxIEuONyXJzru2CO+7tE7b3J3QhPByHEmYF
ly3aDT2Ofdmsq1As8qbOh1shCrC+BL36sZrtnojE0xAzjQPx7eVBNkpf3ifDxkda
28aJ4ypi5lzHsYKFkLwO41dJHYDVRBxgFz72O71nVgB1sSXToaPJeMFTwmnkOcvC
RLntzXblP7thJQfm69A6ve4vj/YWDjFQdFuWwCigxwCofoUiKuCw/9VZmHS8MQhc
DV/Qn5AZG/bJ5JTb0miv0+l33ZczPvDcGvoif8CSgL5ncmppTgr7a77lIkhR6BQf
fY4Kjra02fSANZLqsaEpZuKpBzIiKrtng1OTTwMXA1MkTVmtVNFHZkZ/2ArPnUgB
mRs/xC053hzOXHUGQFxkVDwfjD6CJAnWzf8bamQegFfu0vm/8sRTPCSLTDcfjU9y
zxOf6WL+4qPTKpQzIcsBMjefG179UMJF7wb/sf2OqE5A39ynHq385M+uj8/d9X1k
Lavb8TBxX81tg6FDO82neOc6eMHUg8VT0jYgy31jOUkJUGvCBMA6xPwMSEt8oZqM
q4kt1KfeFPdRFDvGLsPlry/A/NGWs5e7T4qrFaRn8ZPj5hDmpC21mT+9tkh++zPn
E4d+ab+ETMLbBHf8QN9RIXUgPWaIAcXShXFQH00nnX8oSYhjNaiI8h+rXKe1Q86o
BX3NKLWVLRxsDyHDuSizIjyCpsstZIoNJhSWqUJPm7NCUl3PyCypV5FDJPAqPPCX
MlCtk38R1cmvnhxGkwJ99ZpBL5XNq/tETz0nQ9hyjos8zh0y9ul5xBqijLyGp9ir
Oc132+LWfUslcrLv+5UNSu/1l9YtpupAQtm/RRwrbR7KmjiH0zlzmBdwGk+jdOgN
68v94lnCOTk9jp3dFHqu6YYNVHioizbPHeEzG8CPaEQUFYKprkbM3BYfC4VWkJNP
fVTx8xNyAe6vBco45keu8kTvVfxo0Zw950THFaDNzCrzdmSB/WtWOsvmLio6zTAU
g1pl/azEDu9r6z7b8GqfduFrO4i04cWPuMS75K/fWuaZ8Y7rWUrL0Lk3Yn2KYEwt
nWn/UYCp7wjCI9Ain27ecE6sQz/74oSW4Wem6Kd39BW6pLSGdOw+WexQ3zbpEukr
0PShTvOp1zKB+Pl+NYiisZizOH6fvigbwS0s7DPhEaRGSpsaUm2YEXcm/ih74eC4
csp8ueNgLj2qJWmLcU9d4bM65x4+uXAdGBgjh9CM4Y8+8bhyMtAaV0PTUFfi9wyD
rpRcxsG3kfBv/vpYAgo63619oBZnZp3ugSW0sIK2vzUHbFMuAkYYWZO9c6C84zfJ
/iavsKEsey85jy7aFUaeM1Ox0NQnPzfmlAWOet7Q+6YOD43QNEhhnKzrJsgLFgI9
/o18+afEUE2Veodjo7Bdn+wQuXKJc/ts9mkHMM5iwkdvqSbblgOyhzY/NwDzHBTe
R4tGdOx4d6O1e8tbgp8qfOcmXtXiUVuRrquwdTv60t5MdTU8ZnmTqYEfa1Gte1Wi
mbhLN2L3MIvRA/xqDv2s7k/unGUG1TnbHCyB0gnWdQZ1Xa/5JeugpJTZbx9lUKvv
Gn/CF0VkkjztholtmGn8PwvxrW2r1pjIVTMHc8394zhcrBXusETtK1LD3MaFUddC
sk5+ATmVVDEr+BmigxxraHDFggF/EOX0W1L8GSAXU7Br2E1mkVZBeM6YyWV7c5Oz
ev0BTpGu34sFs7UWs9Td5hKX/eeu3f62hcAXTcf3cFQJkGihQR5ZjwMaT07oPBYz
SLlO80rrK8BMKWi1B0yHk67nqmY3nomJEz32a9oR8CwkyIEclWJFJWTKYKS+IC58
sJCuAJVgIMXnMzhoSIao6XrxEBOUwLjwlGL50jMCOnzuK0+/wCZbBPaN0N5iwXNW
SKxzb23aEHUCn0Vjo0pSyHDpC/ckTGAF/aQYD/U2MZvlMLpRqRLjE7mcviSGGc52
rb2QBnt1PLzAe0czUQatGR9sorauYL4G4oB0qtDdjkqWCWj8jepiBxBE6oWRc4ov
QTe0f37Fx9fezH7tKo9MhnMfeHpKu1jTiYhqJ2uO5CqVPsItr+e9X5fgIRoJ/dn1
l1eFLT3sJavTxgyBqLitFKLh9NKh3+UmzKN4+WV8fUX+Pd/25WI3KKaRGOY2do/B
RlD+qvfYlec2foeWMYNSFXDKncXfREGEIga95RUNTWawhaUr2paj8T654nUdbRpm
cZL6ZsuAg7mu3cP//UqhP5oH5QNC8gYIVAQMj3BAYeBicE1BHUUdBgTUA1ZhW3F0
0uUyp7SQVYQ2R/q8QSxvxncOtfrvb9Ys0YhJpTMpooyAqQRcVFFciHGtv+EcfJs0
i8yBINfC4KsFo3xDjbCcAU7rxBHeULITa1oIiS3PjlAEMpk089RjnjcUv7oyBvBX
XNpB6lGJsAsm79NHO7bK99THNxZ4292xoxfbbjTJT5kHp6SqKlnrVZiqkulHyWUr
exwov2+rq29NXknBdlsNHV5pe5Dxx9VpPNX44UfQm5dILjzddCk9c5hiRn3WbciK
+I9bPWW3LKL3rv34hx9BhEu0mVdH9vDRpXvYGTJDDjyUe1nQFHiB8dG7A0NLIiXE
B6OOkt6jO9ysbbIQdQgrJIZHt4po8kecYOHbbewXn+60uMkpFNKMyDldwE3DIUSa
wNEgiit8DPJ4DjuiqM3Na3ZjsmHGWZPRBITL4W79AmIxabn34xTIuXOiJBfxj9eD
V2+4QX1ggFDCOLHTdGC/igGQpXSKQXCy2znYS0grw6CX9rY31E/fGta1zG84LUs7
EJETCxwNY6EtxLea7lTD4xHx1rEpgYNd9fpTE4dBvQXRVfAn7Kccj3g32VBjEd+r
KT7GhUX4pmbW+/ROIzBvhw8DS2q46aLn4YdiUN2klYUHhJTPnSfaeo0JwL3UbGhB
45KX21e6yYCYoGKxGMtnYyXK2ez/gNqZTOgfxLJaFwNQVYt7eAQBVQyrskXduFBN
6eCc0NMw94mT6ogNR5EHOzPAth/Ks6LY5/JwvsNr62tPvF1NjkC1HLSiJVqCpooA
lQnoX7MiDy36lmC5CZdNSax6jXnGzWKEyBdMt2iQvjLAnWiVJpCMnTWxBg+QrX7l
ebY0OVYUu/cXoOwOngh53FxRWZDkbFZkDM4A/uDkKNNsW5/xrfxigWEhN/63krQN
982Bq3qGy5c0O0pbneq6WrxZ90ybiWe5MyWm060A2Ac12iuhZJaMdgCEoh7Q2OsH
lvD8mSYeGVw+SMXP3viACu1j9OFttonAJWRPd0BdnE7ayFPGuUEHPF5m9aV46pat
EY+AjAz+L1Ha6B2o/pWtFZAYtM97TKs9pvWMuV1dJ4w5Wf5Bx6HoRqKPIZpBa6j7
TqSCZvuOvHIeYG4PIghDMSfbgG0JQLaXa+yGlrduPbNAwRPBL3Sie54hVk+18Z21
dijDDpBO8MX5a3dYBVJHsHnxK/buRF9DYBYB380kk9GsVQ6wbuX4St4QWewyuqQF
/hwcnMs+PUkqP4dppXxP9K8aTBv+B+J08t+WDDBQVyP5OmJjPxrJDfqqm30YUYiF
enngcOtww9I6qSnn3jQUVX7qYO2lR9OFuoYygOiMPG0SxWuKtC10kZFSDyF0D4pv
Dgd/tlpxV+Kaqj1v7gQEVkr1afjbUeeENPfXVb5Z0jnV8GWplAtyPEsJCYzDNgRQ
K1RzdrAqH9PLe7IFxp++9+cAOKZD1l6cF/x3DrGj6cN5a5PJozUy13uveqrfU/21
tF51txAUv1QHQqKzUBmdCa6yEe4ADSdROhK8tPBp/EFwTNoZObu6pSPWmy+pcNiV
K47dAN6xOoizaqJvxLOi3rgHKot/cUyoHnvK8JfoTJyqlCaWKX0bDjcNNahJsJtv
tGmR5bcWW+DxWe9KOiGLhQyNINuR8mRvfmarVoWCoD8m7BNQStqTcvnpLdhmPLKa
V6o/uZHBuA8E+GsPsX8uQnXsYcOAbt5GpuQX1JgFcdjl4Q0u1w1a/+2qYqcfZrUF
kIid1Pe8JJH10eFPBhnZxW1gLMAx+p0/+ROJBfkNo+ucsksILsouVCdwvcrZDPth
VxFVIx/XMSYmYlfB7/8dWDTBCzoH0v5bIHrJ66Zps0Hk4TuO5DsOvT4wq4oE1T8p
gTBIq8mfU+CQhvsCRpsoxuIZY47jWTH1i5x5ARrrAY4hRnPhVPfg9KHFm9Os8XTe
Ttpmj5LX8+CqT+um1sOGpakwTRhXEBYGWQAfd0vBU/nT+soHBj56nMDjySq0eeL2
9rqnugJZGmb91vF2s5RMYeb2b89rQRXAQnn8quQWXYu0o6bxITj/xkmlrE8fgHzl
0oGYZUlijqyEbQQGg/Rbs98YgT0+Y85+Ql7fxgf15ztkZAN0uqiQIljk5qBFk+mJ
GIeINwoKUDPVvH0ctRuKahvEjvMHdZlRwawHQ6ju4iXlYjN8x+E7Zm9DOCUlIujI
sg8skJuU3abfUv2EeUsxZ429AX5HU1g2oHIgwbX5jVYU8req0R0FYAX1RFW6giu6
EPnKPBZSSrluXMutEpYRVgVLWhV6cjGlTevVcqmzNpuOrH8214pHvOQzIyLFoGsN
qhtAawwL2hqVpiKkO591EV6HwC+1Wwsg5oBnSF4Dorb/ezOcPu0z7bmJ3KqmXPy5
DURJN/AtGVlbhqUMByLB2cH1i61sfQ3vS5kT2dclaKf0D0fXpEx6H+O5bIezpODH
uIK0hTuVKoh/UNuV3ashqmxIkeMshQzuDNhso/Vhc6P5CU5buT5iFqahJkygiBJL
3urHelddIB+xf8thvBasvGG3Lp77bVauGWK4fK2a01Ch2Ue1WUUXU8fT3fKikpwE
5EtacjwHNkmvzUMN8+lflQbTWXU9bwK4xHaLN/CwjZDpB1AVLeX9GWZfgJ965k4E
f6AXlwiOIC1zLZNCXjO4FpfVJtYFOT/4EE9XbjjEQOnFLEtoJ/Nu3RRpJQMovRvI
M9R/IC747NAKZ2NBLg2Nk4RvDuiK7xhkP+mckPAsWryAOoqbTN3lvzK/ee9RigG9
1CD4V6zaEIHvhk+5QFx9S7Onpbd/ZKf7SD2p5VSBom2Mcspq/zeyOlLYBDZ2tveV
SQ/oEKGKjy0EtyrixGQ3Kv/4DCgIg8UmVCRkLi5f2G/4IsL69AavmLro1A+tV3UC
G4rCBTTtMCAMo5XgA1wITVE6NTpaqPmE2uaadyBnBbp/xYt+u3z/BYU8xHVZuuNr
vdYu3h1DdFoSrDUB4I5ISZWOli5WZVt3leeM3UDSGnn1On2AP4V4bwNKndGybQGK
sWMtY0IZVrVc5i+h4mo0R/Se9QRV0jh91YIcXgkI5qtB0LfEOoqIEAOzzKq2Cs/x
mGyh5FRF36Db1dogiIo+HautR+62HfE+6xex0XVC3HHjU3pLEkiomL+9Kg4NQht2
n9YKXafNtPgz/f4Rta5Q8xmxPppqWa49m6dh/FfBLtMqVjp42JBtl6TwANx74M5P
p8aBmikoYvMFf9mgZOyBIaPF+aVMZLq5EuwSmQoVez0QC2OmCuyA2c8GfpowO8u5
6iZxUGOV3/GgZfCs9mhAIIuyuymumR06hmFaje/cmqrHiZAwj4qYDIU5fIeHaOD5
Btj9nS3rnN4qIO85ojNO6sDHcmPPaP9IDzSXYnkLkQ30E5ddRY/zu7yoNGJaJh2p
yMl+Z3yGJSM7s5tAV9AQ9nkgMAJBkrpvGI/kOCDPEYZ/G7uKxxy7rmRACVgObZY6
4bd3PZ9tx0N4h3RWzk9cwndpCej+6QFjn+m7Tg32a0FD+dGBnES91ygeksCHZ1rF
5OzKfigdpGFELYcxEiQMTeFn+KxGvICiaxikdA6+qqVZIcudE/+dq5a9bIVJpFWD
71aNe7ecqpNLBcqCnuK+bWK6Ry/ekaEnd42EvRiBz/OnPd6d76pTayDxMfOyurfs
sYbd19czFD0BdekZUi3qYoVXiTLBI/nZTzrgP+OFsSVA49ny2vT9SSBDsSFZ197g
VdyHQULgb3TiYWnkuorXrB1h2HuToBlp1oXLTzEqiFBrk/ReQKvwIbvtl50DY510
G36/YYRz+O3hIaa7+oOk+RXuDB9eVDMMMl7U8rgqoPxcruyKM/gUmr4EbLIP3PTj
GbFWnJ76WbgTawAlG8ahAOttsVg9dsF/RI9Az7VH6sanG0aYAbMHU2Cgn5R5qafB
Kzox39uiEvgoE7/3E7xRRx/3bnyK1UJFRCG89CkhXulE2rpxAbWPuvQOf8fQf/1G
JpuFbYHfyPdL5YiV8HE+K3gLMkTGOU45OBNpPLLWvCwPHXJF453HiBcmDFwj1upi
MGt7LY1uqsZyrgt5QR6LxNoDjlKsa7hE7G31bxQ83ET65lB/hDz3lzYxSHisptPd
NM6VYLKPhHezfTty0sAot4K4UwT4eX7BfVpkKRMlcznSIFB640suMJeqtR34Un1d
sHTpG+BbEXnbgacFdrZvmP2VoCEZr/S52tU4JXCL7UlQOkNUIiMb4PRP6cOFLBM8
0ygB3168tGjiRqOOOr0UZ3wLZm9dodoLEErJMYueVH1TjHhDIrWOclabNUjiuUu+
M2/7hw4YOZ9RJvTIxamRWLqCcq2CVvhUQZNLa5BIrCF5zLPPhYYQgp17fq88bpK4
E98P+OmmZldNUkgVSR1JCv4N97b4lyNxHxqdj+Hdrge4qNSCPCMFR76+VOCEaFXn
LzepUuA/iVnnZ1v2UE0How==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ifOD00Q9kYPhPoPGkqtPCkKIM+mQ9mciPhmNEMYD7Rc62WAVF0WcwldsXzJgfJL5
UB8XIlSuu+yY2LmGfCkqFPZC8v2UpaeG9idIzxOFs02PT+gf52NtAEHP0nVbCZ8m
PorjJek9U00ENYSTvtkxLGmgWi+GiEDzha7edhESkOrIT35Ye2/kYTsEc62kZwRL
EETlOkq4ejs+WKK++V1F+ev3aH+767RCwdj0XiktCef8c1EHkn+s8WjCCp8fslQ/
ZNwJFLS6/gEFDxMNL7Lqd5UtqsM0bTe0eL5EiB0uKsuQUKPCbNjqhEl0zTxfAWYn
xiif6nWTwYmFxfSEP+C0BQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10416 )
`pragma protect data_block
GAeo8GYyYKsuigzvogj62sju4pWnzXUtyeQNJKtf8n/73c25STO1xnZ9KdS1OLgs
FUgObsnq9H1WNHBDf77fEGAvfshvvDEnzsz0wILcOPZgBHnvAL7bBxLkA+5vEHfg
jKnYuKWwEGkMwIDKeeCq1rc0xL9Fe85/GLlb1leQL65WAtdotibmUaqF94cXG08H
X3QKpFJ/vE/Voa9tig3zAIuBlC+/GljJDYHb3lNmYThR7xup2lJMIkvdAGEnJgG5
BiQth3gPlu75wZhBIsmhNW1mfD4HGqh3lTNgEeqGDL8GgQRNYAxypqvnxlP7YsgP
yDZ9gSrEPgGtONtO8spyoawQK09+qD6e4GSvql6kK3xI/+9h+7F6krjaJCcOz1jT
TEPcPBfZeNClUxW5ya9qbwGoROf/EKhlUcOgyF3JEqvly+66z9lf/G5wx2p1jZpC
f24ft2I2It+rwywEhxTZlQDBTKWsV5eZze3uw/F9cMgASvBtJ1K24WwZCxSqGC/u
NfYhTa5uQlq4SFp0zHWWJPqcvknrl3y0YhILaveFD1n5O+SEC1knCEzk8uvwJZ5r
b9WUCGEUX9P603AMDUEH9G/zp5Y4Ej3eYhr9MkxK2+SuOX2mIokE5dFbYHhat5Mh
ky4U89etltvd0BENbjnw1nOI82zwMsYf5mQs2YoUTMEqv9IOwffEiWtX6Y0Rl5hO
WpJtsIpWAnp2+43qPIwoBiLWQtCSEjgQGxbkHQDgG7P0XQPFmUW62tnt5KwOqE4a
UfaNf8HFC+x+LpwC8PR2u4cEHb0Ik3UkJ9buWtYV/x2A4dGfTsFYfuodt+Vk4S8W
1vHTA1Q5F/SMUj6xPpuNTm28aaRCAmI3N9IKL4v4WRmrxMmVuX5tZPRniR5hotbO
4ZNhbSl/68LgiRmDdn0+xZxONNP0vv0gZz3VpMba3adqc3Vevm6Zoltmb1e4rex8
qSKbQJpAnmaL929Do1YDLfb4gJb7IT2Ri3VeTtwwJyb6FvxosLlYSj80ditBVllj
DRpGNzr1fpasqiWKBojv4WrL4+62SiABbHVYM0IMn8u7l548F0Vdyj76hk3hRz4j
2jB1Th8hNPEV7VQ7NDxvRVEuigYSDSxXLjJYrXvrMXg74tGzwOdEvL9tAuucrCOG
XIPPFkX6zC/V9/fgZVoBvynVxAN1F7H+ky+UnEc+CHHDQOJoFfvzWK+gmtA6v+LA
ApLEpGdKCfI2Qjx8IXGz76lpBNHAys7FLiFgMuHPFPcGRhJDk/xaXtb55zZ1IBlN
Vi44AQ5q6c8POCOCXC+9YjGMclIKCuXQikSymj1iU+KulTx2lHkhnlhbwaSz5OhD
OkLCD50FOFOYAWTIc+rhlrdTxc8soyo9gApgP0X5SUbOQTHtqipZs+fWEGsJInxy
ZKdDRyQ2OzfJfxk0dyOj0gHcfmWbj6+IA1FvzRRl37+xFbJNEvvEAT+wAhuLGVkn
yS5GU3FThzWBDBQuRv5IbbYYPh2hNLuIK7Vb3lVbNN4mSYQP1VD5bk53Y7duwj0w
CRmPkTq/1sym+YQuvXg4Vft/5JKXYUC0ynhRSmNe8hneAMLDMZmm+qGlj1XzJZBw
xgyJ1pz6wzElL8tEfmOipKFh5ZnlWgQGLsh1juczy3RvSSLedCBICjdgkySCavd5
pOIA/uUFh44W5LnNbX6taAsSf+JujQKKdPhO0Q8WIMzzDQlRo1tx7EqBIuxJzJH2
MdJJSm7i0U33lHnrUftT6n2zVfm8lIEAhN/VBWrFV7Hl7ocihVCqNIFThCxYsBME
USimoUDgeVjZ+5TVu3Mf+/kkgXVcotQLsFOuL7ln1W1BLjJpXPOBcP0dna6lM+VX
zIK50ircsePpWGKpW3ln3+ajEdmR0JCC69BFNKOtJ7XkDyxM4C734TKf1Hp1FZKf
kdSNEIkjOEPc2UEBktTyMDKEuzXnls5E/cIwnWelpmOECvNrRajhN6pq80yc4XXy
51kI2r638HWv0jXSXEttLawuUQ4n7Ms5Xe0ZaHfbyBFQpu0I2lmNynG/x+tokiem
ySL9CjY00/nc96QhhOBsB8JvDkgB+b8erBPZBIQFx2LMRdXMvwpBxQIJtKYZyvG9
APuOPRzGJqwnKkNYn5BEzo7jcHh+5u8C1WG2eOtNunvu4f/tA58yHj8pGzxonSp1
cd/PyuL1e0u9oSH+J3rXGuXceaScrTvkb5GeqCnAYhgqEeCIRRvcsxJr33Jf57nP
vhtGbIAoKWWHT7fyl7HSV1eVSeAKbcJGFEO74HnzibM5/OoEDi8K/h/elSU0bq82
wNmMfVlo9kAtSf1bdJ7QCanvrqdLOszb6ees7yS4+tC5fkIBroqq9kh1Tg0V/HdR
kAzyc6crgwnNUNVRj0R4pjSYyJ5iX/EtHsz4vPH1lt/aoyzLGjHm/GAzG27HsSKv
eK7ESHx+QPsttnou4ZixAZPzaSGyglPBRfr4Hl0slDoCLBodqr2vFOYqYv5fwnhV
NYnQU2hWf5+Lw4XIugRTtqeMz25qqNlPsOY8UJbNfpK4yJ9WAcQmLRD13uswZaGt
OwqgT4nto6E93oEjW59AKoLXobPLqd1nDfrFD9P+TssNa+5hLXeeli046SZ5KFAI
MGzBz77GqQLxs73oWLas4ZJrne4+6w7Y5Cwt49KALbqmu9IyARfdjTjYAuOUyhrw
wSiAh/OrP9GlFkjSuOvR2myjgrALjwkrALa1kr++p10+uRiq7vf4VJXjw/QTkMqp
O5zxpeoDR+/rZltJNwpLvM2YKPCiCJUFgy7b106AT25aZfOCy/p6/3Z7GwGDGCSy
xOsyRjPZn63M0tm9lw4uCXhMwjXfyANF15c0fTGEWjFQKRNP259I43dLdvAWX7sn
4MyEjfbxZYYluDSpNVY9FVIh2Q09X/Y/Ym7H6F9WgYHoMX8JcQ+MItoMdJydfgiU
5cGnV+MgKenc/NCz3oXSZDZ66fc4/B5VneM1jVUnksKywFJIJ/l0oJKXui3CAxs4
flwXBOIKdfml4j7gdsNxnPNwcIswi3d53GGteiMnirjg9+fYZ1TX71u2GzkBQ9ki
SpAct2xfmRAOt25j5+mi/vMweQ+rHIehIC0eBg02/DNJjaAu1j63yHDONeE5qEZv
6LqsMxCUki4UiFWJfQoBnqW7MIXlficOvCTyE8NWu416mAXoFNsYQadgepXaIK50
mt2SFWjlryzXqoo8kuFyAqEbrHv54wnlxsuxwjRe2LgtQsgoiK8CMLpnrg47oq4F
42TQFEt6XEgXSbiaxorSEhGgR7gURHxmuVMHiuoO0026qaxndY6YvM9AI/OlL5kG
/YngrOlikkRch5XZUakClmGXJbOPWfEJRukWCRm1nj5vdEu4hset6pNR9f0IeKrC
FRjOcHNRZ5bb8AIfF8P+jHPXL3X/vhakWP1rmmR+nlLjAeZPJTAn1mP44L/oKJk1
KpuKv1CCKC5ozPpOGP+inFfS9dSwK/Ts2mYlsSRR71i1AXfhyQvjjMLaHhL8rc1D
EzKTon6Gzsptzhh2VLclOlmrQZOn6uNHgqIsJ7NpCv9XDtDKPV7/fq7NqD03tKHm
U2Wx8DfQNZFLT6oCAk+oqEZ7uU3nX98xJGRLT75+z8p0AHvzTA0bpdlJO8qPRBPE
H1kO05/gocYAkWZjuNzWsmugQgJbVHwQiSB/6lvV5z/ty0VXlUEMHhgpxAP5EH7E
oty+oh3QkL7X7DKGxJbZNLkWfAlo5Sknya6C7dEMPnTxrqTEJGEDtBY3k3V7PJ36
s17lJ9fzHq+pIlUFgvSCyZ8C2mWAoU/XLI8LUgn/N1bXwvAHWDYYoaY9B8rvwxO+
dE4PeBd8SQ1O3M3s1j1KFlKnV5zYT5lMbscJOHBfACVN/GmTz6WrZZoULY6Ygg91
DEcdnM5ByXWFcec1ns0qk6vaWzSTY9K2C8wdaLXA89sIWcbxf3jbqBNWq0CUN6bM
bALbnid0nLX3Jj791t74BbMMcgOF/6wp59u9mKtGpiiQxfriQUIUz5d2ortrf8KD
utr2F66d0j27yB8RaqJVcT3ugKvJ/dJ+0Yh+seiKXFpys5LPJS5BZ6wkIp7ZO+NE
QB7wY5VKLMy8kw1YLmLBztTOMGruvILZLLRhxmaGNHdZ4eTAXDXKQqTczhXLgMV8
ozeKFG5fzopF89h7zluv/qRvYN539srj3doUoQS9Q1TfKf9UGY7Qx1osiwHDtiOp
+Ceo1teRZkVPef3JJDSnExwQfd3Y0/gzKcXKri94lvhBq+DU/N7LyY60zwiyMe5r
PuL8pRdgCcwMwjkNJJDzOz+B3EWbafwVJ2RvAWCy/94WA/eFPXWv256/jq0g6fYe
Pqwtjq2KCf2jUyrlygPsebyhfhXHbDl8JgummtVAQnvZRr9H3m3Edk33HdALcmuv
2Jg1yUk1Vl0TLSIXuc8QW3ygzmf5u5hoQo2MAETkHDjKTazWY6FaKj/vnFV86MSh
xXO/XScnsWr5owHeb+cIUqEDdgTkviUJ+VeFDJFl1fo58ttk0ZkLeEpDH/fTSV9H
xRr9uaeaP80uH581S/+dsML3XF9TTAhjuvyACtqLJR62ZdmzYqMhXofQj8R0FjjN
JE9ujddzO1EvkLEQdaxTb9OBuGsd/rhIOk/ySgYCRz7ZGe6HPbrOHDY69b2bs+qJ
uSkdY7a0kihcmaNZLoZu6J2A25QFcXBL0VTQzg7YViC9n6PXnhCABzUniMWAdK29
2bl8cby8H+dUeWPv/nD9tts43oXYN+t2PF1j0AXbIcQdhX24qhxLZdkAya/ETk4u
TrEmyluKk97ti2EqwrboZHZQ/ibz7Mg69jkhItaSDGv3T1prDb/fPOXYNQ3YBTA+
I0wzb3rrXWYT9Gc+Eag4uHAGC1PkC3B2QvW3pkiM4oMhge1dkRyDJP4t3AWIKOfW
7lT88LnIdpU6lygpgU/WR+FOQKxbYqc8Wqo5RcoJATP0Gi5kD+2FVM4dSxQGRoev
im4VVtTsGdQLedHKEInNqCUVNXEcuaG3MYs40W2vO8O0IbpVOXTfs7QgXeBg04R/
dS4yTFSw5QjWDxQmfX+KxiNXmjxylFvHkt1fvPTr9mVVnZCsm2M6SocrgK1bQn+4
p3N1WwGSBmF5S8AgMcFZZrBljiqqExYXtTSryljqs0oyTbyXUnL9ykF6fvmhSFtn
dkJKkyPVV0/0vfTeJ0LWk+KtnuIjH9ICxjpPvzV2ShkHCBpNVxyhgdds8wAWutT3
m2A2vxu6rYXiJjvnNACk9GYD2229H47otvXZOzWfHQJF5UaLT6Do65TGYmbVUs3A
HTHCwyZcUH5Y0c0KBPfgFw4/VrNqYTh3aQ4CRB77N2NgvqpIH+/z+yAgbiQw5/pe
Y5TXwKKt7hnCz7F3USCVoZ7VDi0mNKnwlRrdtrEqCw9tD2X4zFkOFHhbDitbEACl
o9iJv7JaAfhrlYeFvC15HbTjwyJyjhaeKxIl6y2n3/MVDXRw52vCP2T6Kd8CmqiT
qQTEliHaGmuDsvyYaBuy76SRRrmdcBbN0S5hq0vaW3nAn2q6xJuTPPIHTMTAdBB9
OgzvhK3WcHahcJ9/TlflSe186LZvWDAOGCheBXLBHGG7/e/BxgZnA2k/RU3f3oN1
TP0Vt0qU/5cbcJh7hn7KflP0AMml0qzK1BAx7B16hfRhTbwpOnX2TtttPMG2+hJw
5J9OKvC0Km9Io/ih64UvHk6dgFjMVKJXbSkeA60G0+TDAkbTmBsOqyRvthPMI+co
6N1N+K/rHzj8bdTYEXOSP9Sfli4z503rlarQhOBK1var2dg9KCypNi9O5lXGHDRG
+DVErhJAGg4BNIVdZRNezUX9VDEp80m40AWzT8fLpROISYhblrE4aSAqBnJUtFW7
u6uNyXX8ifoGSQ2IMAZSJm/gLiRQtj2uozRVpCjTTPI1XI7JUybWrk486i4eK2aW
BLeY3T4dNIYbi6CHsG3Ism1/xj6c1pLNoue9rWNX/G0tulWTTGWTOyTYrSaO3mX6
+A5OjYstDpT+PHOHf/r7jlctPvCiXpLlVCrvl/v5/x9rrKEtyWre4XwP70iFOw05
JEW3JcJs5mwLq/ZOSfcP8hGsjxlCJkDOE10BqbryLr5j4XIGQ6kJ3XXKLSSBiiRd
9eoN/C/Gp7NgttANIChlUy41Y6mmvXxgvXVWuoispcvaA4LikFGf/6gL4zYOQgjC
riG85Ov25u10SAKyYqFdJ8kNsg/eF/3qxVBdxl+6GmqsQAlnroTh+bymalPf025y
DVa891uzlpZgIMFYW3rPNIX6yZkF0jnoybqkzsa7NkIT11BCYgDusWHJ6Mp4v38W
pf2Wi2MRYYgKASiSNwVqi8NhbySE2G/0b14IwMw1OULN6zNbb2EgRLB5cyN0hTzw
qkR+zFLH7zxJK8LHA698Sq6GsBFC8SEhDmDJ6ORNfTe3gB4niX6VcGp4wtFugKlW
Hy6J45+BbRkAgE5Ah7gEQ+kEkyBIp4pN6d3k/Iw7JKv9+wIpsnMUhp1MEZjH80wF
j7qDx2Z4ck/Vh19JWDnUZnvq+jxHpS+ARyDsvNSguJvnXMjlR2OZDcDf0P8vyeVQ
9j3LqlpTiPCiMZe8QP0qjSh6oMw0fF1xNZNAnuVn6tMHgpST3ZXnF5XAm2quGBSg
lMmtcb+sZNF2RFPzRZfAaRwz3BGtku9q40uf397iuhn5tXAm4fDOm5VlL3rjEFRJ
P/+hwVRPB7i4UjfubO7TP2o3aQZgaAvl3m1d9gk9WnPEu/LHzKsinY2Fji/Mooyc
8J/6m1wDjQwybyoqH3Zvi/VZL/SgbgbUtWExJEpINkf9+3b0X7aD9j3aaKPDSHx8
zAKeCaI7dNZyFMJHdwECQIiYA3C6Ghgqa/4qbOJmj7c5VNXTJOVNni/mPuRuWg6U
c6dGEejABSyhtZFnfv6Q1ceeaM1gY5kAMemVxrhGfdBOerr45bYdTemDMV1uNfxR
BFfs+bvtYrIOPXuD/Ro0L3fYafSV0YpYgVpXvQLmd413SKmJFSwQqBJdA2Um+8xC
e1r9ECAsBzvRjoFIDOZnIeV+6LXBTup+nQK+/VwKrPoLz2eAOmKTtnjBBl96uxiR
PRMzPR/cFL3ROW+M6Xt463Q1z9mv1H6IX7VB9BFMa4JslMDlH11+k8YTEj9QfCRc
ySfep+jGgD2EAKSvjclEeLCGI2PwsKVSkR3rr2uL9MovpywixCPsn4jw39WRkR4k
RbtS19zE/C1WwaunSe0gi0yZPXw7MALxklweYm8eFZLL1YB5yNv0iyRARIXBJ2XX
vXm5n2ZPIJlikT3Vme3GIBATirLY1VXF0AlRFqHSirayOaPyz2dcVgEPVDEVFOCz
38zx4vZVoYQ/y6pWUdI4gD12oIM1IV5qzy+wpuEjy51aNsHSlPBq4pk70HmeRz4c
qMJe99YM4E40Tk4cTvxbbZvKLRUfKCpdvJHj8YUN3FeK1j8rPgx0WrISGMlsF1eT
y4Y8hbIwvbfrMPoq3CtixlKzIf2Y9hCfx8O4xrvk8xvzDsVhmzLAZ/lcp9VlhdDi
e9rFCIVKLFwLiOis5KDQZU6PErQmk+CLhIla4wia51t/VFxnlgeY7KfNHlXgEm1l
DVSJ6sIV2TKajp1bOxdraJKfARPbonOWrEA+zV2/MT6e33kwavuKf4XrNrvndAHZ
Pt9OWSRpYKPEnhu4LJTIDz6NyAmO0WCu+Shak/TW69JduJ2zA7TpfxtP1qbAy3E4
CyMXresvpkzNllNZpW9/p804iCW6KbtYfdTbm++hRapGRKXfm57Qo/XVZIrkkugb
rCJzgWsw8xrGQzRWyNfs/uKE0w+l2SB0zaRgJK1A3KNw3MOxOvp75NCC+J1D/WCO
qEx3awmeuz8eGur5+OPW1PdzS/yA35d79zE5gfae/X6sPXVAfAnFbQlTr/ikaFtv
J6nrVBc5ahI2ZluOU0XyriSZ4L6oKIQKdOEAzrVvsOPOrTnyAnPhZNj+DnwOwpyI
ynO0EJX08nmPqR08kdtuwkdXyWv9taiKhCG0tvGqwp0KBngt/L8g31I5YO9/kcpO
F5xxqjrQxKjNduR5nQvfz7wtxnkHCL0EfSOjZHvoXwgS4cRfsKbW0+Y8tO7tL+F5
ey++4yV1EBexxWYT6sSVw9+9vKfJUJ/rdbp+XmQwncBNuHr7hf6+MtZyM+m/g9kV
RRSqV5/ce6eNJSdTG6mCvJwPsExkp7ivHriMb6d+z643RZQBIproOVSPsJ4T2QtL
N98DCNFjXIHJ078Ewm2/X8nc8kw6jmCM9VztEJSZ5eGNPDSxNeUXUg90UeEuBAkZ
iaCsnIj5x0uJ9feFpWpkodjLH5YeTeKwMHxa6o8X0xbb2Qe2B4D/tnDeYOuY6SLe
dwGa1qzkRA1DeHFhaOwLdRnauF4cuZ/79xMfHrh7E+TBvffPDnXHLdFHI8YUB9Dl
NvTf0wNisjYqKQK2eqVzw+uYO+rmENhoABTLdRxEOpLni8kk/tv31OEU5UVfMnb4
0ELJ3jd9yxWD+fDLBVVGMgKqDEtTsUAeyqsSKzA0QyYaJMHcsIqThs94d/Dyw+R7
gHollu5FhrbhGrblDRWAJ+XFNMkxaevSXxxG9Ds5pukvN5XhLFFiwoc1XSUiIksf
UUHtGtHHnHl8rm+FBKnjq4hsZcp2QUXk1OyjBN/T+Xo1TXcKU4GjRL+C74XWw1HA
Pj0ceCU05f44UyRXgT/1HMPNP/CFmUgwfOnxDRuMQ8fr4CMMJt4aaxbfTGcJT+oa
GONCecm4hp4gPZJKhG7tzT325HOH927j5r5cRo8pWh4aXUeihazReuFnhr6+72xJ
9xbj1a1H2kFBGwEzAmZVDEx9QD0Mu8w9ItaxTGQ9CEqR55h00+xlrnTKqYl2agG6
Yl+xmhoCE7lruGXTgwmL+Ushb+gMfElfEQbuHpO5QDLhkSPU9J3qDFSzczPWLqJL
zyTKxbLl5rgDLzkXMzmG+Z+F7T7Sf1O6bUOgzbjl6Anusy6PGxjC9/zoQ2oIQrAv
oCpn0Jz3dpGiEEcObmG9nMLBetvpfyHnAtGK3dG9KPr1SaCeeZzbHaPuy2wDexXO
tAmACIGWbzkAfQKktxxCgGdHKc3h6+cv9c8XS1EQpdwDX601vZOYGokzSS3wKljb
SmoIRoeLOeeuy2yOkl59kPJEB4S3OeU4CNZXgb0ILyYe4tj/H2QG81BBtsLrSS4h
w5vmPct7cX0B8gYtwGiMFBKX7l7FFu+65HncGHwtYej6vAT0U+ZaDcnr5kk8fV5h
yLVBC20777u2ZljbOrxYv7vcJpV7Vjuwkx2sbv5GCX1a2bUFZgEWyOgVqxPaia4J
k2X58urrM4ZkixAazpzwZj3+2CoLWMzXhWvk8xdzo9OTD4qZmZ5OcKQmQ5smWZkU
IsxxAzP8h04hh/3346E1HMAaFw/whAWH3fKF9eGB95ov896u9L8Iufz6PniQ0MXc
hnmJ69MBSV/ee+4jCxPZhD6gWAIxVls9UhgHRbV7YcuNg2Xn9+geAt5yy0tacgIY
MdeMh2bOklGejXlHA8G2srgzcVT7FObPLMMMGF5+ivQzX1pKWMHbqTp6Jasj62gm
YNJveQ0xDlAo6sXNYzfDR6+uUdnahp3ZNljYTvQlG+9uBEcikKt4ITLlCO5V4wcF
xU7bcafnCUlBs/RhjtyJgJk96faFMwvPqABsn8uaXA7b3Be+/KQzwdX06v4pILi3
CS2R0oh4GyZ+qSxi5k8w+Ydeu1q0LFtmZsh34yCt8bNmc4nSe4+yjGII4ez4hctr
uQciDHI0FC3oaw+dCCttSlALX6T9vdPpUgIGwvB0ZNvBQG24a40g1rMqtEmA06Tg
kEFnHbd4LDWbNbO20OebG3BgDtjyy3TAWHFx8W+lI+pWkZ0Sez9DaHljkHK03Pq3
wkksbLTJF1fUdC0PzJpY8lPyrVySbfuDEFcWIE1wIhm8EQFDMDux1oNKZYXKFf7i
OCOtp66BVa4WrgQuT4duPE5E/Ixi7OwmJcdIR9+zCIWVhN5ckW0vUgTC79Y0y148
ZwMj/m5uomgRekFkqdxptesDlREaPdwiHEoMSwfrx4XsW4k0fN0U6SVz8YL+L4Ey
O1c5TIzb7A1VbhdvPT97C+TzmhfM3MmfQoPubkeC0Y/jrgPeDzqk++Lv9pOlJjaI
lNiw+JdygwK/WnNhZmcMccDyemUjmRjgf2bz1ToyZ73U/FHuOpPM4J7kq6iidK8I
QBVR2M0VqmAKCFrf+/fM/OqX9tS/pumy9XEQnYzWhfVMtKfEm7R7EIfTI5EjSGoU
6J3b1QIOcRv3DBkONlQwaNdrUZkvJyjqLSquCxbHYJObLEKoWj9yBecimDAc6Lb+
ihfIGj/0aCRorLI/3jd8TVeP3l8D6uRnDiG4P7U/PT81jTvVtkKw3So2QdtCLS44
n61NSPVi9lFv9tvZyTxp/DekTLdxyYzBeIejXwovT3GAOX4/zYrkMPVTZU0G9JeO
qJDBrlldDd0l+XMM54iLtyvgAJm3OChlTxJA9LNTEHuTbqzviNEFQ9jgNl0EO/Cs
lrAW+ECtkMq/uiuV5VFurqqvg9iEbDYGGxlvZAE/mUZoR4cZafX7QIQPDHlQ/t8T
CWQZbMslOeQ3DLyX4PoCbu/O7cF+eUoQG0dtV6HF2tlNI9R3LMPC5i3t/uqDxoLh
DgEvlWZIMwCgCDx2Tu+XLFS3VZmkxLrNpM634At8UkCPZQw53kQ9t0ryCufKDGoa
4RSt59B78o7h+kAvQr4QWKlqBSatEMiDWOgC8KY0y+asKT1taziFztv02XCtqMx7
e8II7Tg9/NV9UMBZkgN2wjpNFqroI/lW0Wc6Wf3PGYP2Ke/X6hTqlubPY8ynsZ91
QKYf61oGOmu+qM7G2mrNJHMikyfVT5zbXefXR3MZh7jVXMyIV88fSrpvCWU78lyi
Mpa0WBsIjEb+L54uTSRJvUcNMlPeB1CbL7+/K6iEAeduLOiZVs/AE/ec7JuR49WF
SiNJ43TURDBHDgFgwnUgykNxjKboc88/9Pp1cVP5TMfxXs0LZQQ6Lmu5fJyKDhX1
JKZNxTZkgxrl1wqGsYue49Tz6ehMKhOnhG0jy81NFSvafeNdpS2aqdGTUfZ0hedP
tjZWPfAJwF/Mpiz/S7vKx41Y3S27iOEM5MKk2HQNb3IVNcltv+N4FFlJOQm8wCq0
NglQcTXSOkOC0B3eFJWY65atDaXcvrZ6CfCP7xVF6Nh77C3nlirdxEgFWu5VJyQq
iBfX5I7pdybIv40v6pej5SnbfG+hjgwP0ItEfvkkHGlBF2fUmmKpN+ANdxjMg1/y
JbDucoARbVm33+A7OLX5tKEVuE67tlxkQ3BAAabtk7JhPXInwLv2vqWp5wVS53vT
6nPraO8TTUsz8IN7xxOqaotI5N6sGdjVv6fpiwEYle7vO4jwLLW97lgAQS7LKDOs
9DgfXPI/kRvYRMBVY4DCDerN4zjG8lJ6NTekjBJ1lfgs6P0n+kMTD/uwv5GlSHRs
j2z9kAcJH+B/56SUq+/yTxCGGD8LhRwQ1mQ1hpsptJsV5aKKOerEQaxh2hCrgEZ3
RXA7+ftC0qNCavDxRATp0gDpaUnpblEhRlCw5WkX7ZeR2X4OaiWbMu5ns/ZzGvjM
bnytxQFBWV3SjRBc5EokWQ0vrYqHSEztX9MVi4s8HdQxlxd5BQ34kQQNehDuQuvz
Gup/XlSlfYN1gE/u+zhk3kkppFa56gKFa9T0xT+tjiBzSB/Zxw6on7Apao2X6eoM
+VAZK6z24rlnZB5ZFj2S05QDseWPuM6E/F79hW7dmxhwMRnfZn65cYJV9XCgqiCI
Hw2wuEw5UQUUsoZU2CC1HUPR0q3SjwRqUNbR+EpLgEE7i4c6zVKejI9Mb9f9FGNM
Gol8qGe7gExsAy+Dyt8ZCaMKbpT+5MEF/StIAxg9agkfkH7Y0VqVANkgKCJ2ejiW
Lj88YdB3vETD34bQTQDcZiw8TfTzanvKHQxXcgK+DwJjCM+emzpWjHj6m5xVy350
SxXS3hGrTDp9TP56aVpkR/wMBb2vNHT+f9Y1BrF99KdLKVyX1xEbOQCiJQMFta4i
ySKAAaGAqn2QefeDe3eH1yQfWTjX3VdGMoJQnOne+OgQ0ey7hmhY7nKcH/IJ2dFI
MlzpBiPSNlykBnXhZMcoRaaIE20TTryrXXpX5KRjTdbVTAUClH1SW8HIoLpyfmZH
vY91HZAMRjSrBSm9jSUZyeo5gvozE2A5TxQGBmckmrBie09qlDK8+ycnbtcbfe12
1ElJSyd8ADuTKXz36ULg8fiK0qxuINAov96+YfQjZvXdPqu44PDPiyN6fKy1lHul
3tGdfd0TdWEEYgOROV1P64QFL+zA2Uab2bFDBPOFF/JHih78aorX9PMMbim34IkK
42+QuU4JsDmBiPJLjAp8T9f9aVaQ7H7ubiA/UImBzZ7Uj2NJayOeZTFG/sk9hJv8
8tijDJh5JowHhxBCOUatn4Ho9VpMaHtqNrtJwJv7UyH87SfgV12x4QPJkhM21kAM
mlbXKTVkGrTqu9WHFdGNOg7gLnhFuJgQ+TGwMDknna4lYdwBm2AYsVWshrFTn23q
pnsl1KGyCClwkmO7tuNCezLpgEY6vkaDpC4UvHOCroRKrvIBOrKsn8CseR8EMIxa
9UpKJgI5Z2jxTQKAsm6bXsEvblQi518HOf/tk/+w1UX74SnmnuduiXoqt+lRRJ9f
2I+DKSgJhY4g8cz6prssY8GgC5XOu10wpRW2o9mWcve/USGhZViO9RgnaDnS2PZJ
iseOr0gg0zDAki1Mcm8nBflKZuBPQ7eQR9TbSpRZ4uYAVk0lQoyUXwy39ZY7vaNh
/WN4wKKY42SjR4YK1LxhnAQBEsSOYPPMk6WXDlyladE80cs/hssv4eTPa6FemYJc
CRG3aJMPxYVOYMk91MM/D6UWEs8kAWtMK8DMK0pYc1QZiAcBEUpXuKUnmfGKlZHD
X2pjiQXAccix0s414L+6S/9mw5vdVLUHuKFWR93deUWbi9lLW3CLKqouKfHzFsfK
Y9jxY2pjxDEeXZtHw4Tseq0zWR4z6V7fto0wFClRbLBPbw9eACF/ROi5vEOUY0UR
ks025zPnW2xIdHz6aJe8BLK90PHysxZcC8q/m20UT8mzKVwY4OrR5ip69sTGWU1U
LRkjSUTZNWxqZaAkZHf1kxYRdt67vGJTZ9B0hZ0UDUuEar2hrnkLJqFyot67dkyP
ONnRPGKFOOb6Db/sCT/Z7drKbq3qSUcq3hbBE7Yi3+Wbu4z7YHjKx0dNxdBf/x4o
UMZMzrxIalwVjgHr6AVG9L+UZjKeZj9FSt0C6zvupBxyLe482aiIibWfL/TSF7aG
OnGmL4IEZFyKnDhNfFGv4ZfCZpDUvboOY4dKcYFzTuyAIp/wiulQ5GjiXqNZad1M
2OTJVRVt8y2V0TJH6/st9cX7VrOfgLUI88Sxp4XHy1WV/I2Ys8Xuaori/xoSLRh0
V/7D422zt67pXlwJZnZCZazvZyyIRsZjIf0TPraMC9TiCI6A8tJs9UMi5B9v4cPZ
+mOx0TGdg5R2IFbwThffjiG6rXDg2iZ6Lz9rnEpbbEVv3bVhHF1KmXGG+W7uJiiz
sqTADYf0ukLOe6n/ZjJ+qOzHPYhiFnK22EwOEXyCJ5rF3PNd+1SrSRwZPVqlt+Nf
MEhilBLKOWqqQQn2rFuzwp62YJDxBZce6ouQd0UijpwzUBAC67PpjckCCcgjDA+6
b1Dr+K4g0mw2QYDdSwFngJDKCUQQLhlbfxxh0uJjsEoXQuGAU4ADuH8kz9+QMf9P
Gq5wNZebZnTX26vyDuQ3FHgpKu1fOEz1d/iC/e9ssj/E3tkxmvdj+WKOCSdkQ23X
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ARngcu0OIXlTeS8NNp+7JmMj53cpRQwcABFZbRkNt8tUjjtvjaZczlgjccIKEyEH
thww5nEFGSxihmk880ZucZGbzaaAYYxbe10jIbeLYFLeWcfkgBordGunLAR7ev4/
vkmpdEBwhldN3KgSFH1isy5CZihmTX/sqIzLBRWfdsrXpbpULMN66DNrTqMXeNPh
oFMiq8pbWOMqUMQPyENoAj6DgvjPH1Oebb8juy2mcLU1KH4MxMC2R5oA1c5I3v8L
ALYDdIOTHnHeETJOoPrxGTy9jreYlwgNgreMdLMeRmeMt5I76hWEbTA0q993N+wf
If1lKs3a3GxhnwYmkKc9rA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6016 )
`pragma protect data_block
baxZqXDcveQLr6ZZ6iNrKsvZ91sZrLhttKc0p1rH5E90KR4BaUJrcfw9Frc08dPz
xNdgjlI/qMdAClzQQHgRKA+zo3hmxFb8dJc6UqdcscJwUXc7wR+Zo/FJZd/smhI5
xSHDDj5+JdRpYPBpu7EKozmbCAYfCQud5Jv4g+7gfZI3uuVgvbCkT8usxc1fYWgM
cPvvO1cA1YdBw174c+sysLRZPlyl/CtL2IwoBWXZtnFoJh08cIr+RLAy8ercwci+
lwFtETB/yGNkXBqWJcz6iJ+RhvSewl3QSeFg45+d+CEhuNeeDgWXmfwx3VaBvh3c
sO+tmUdH+vcCkgpD++LvUobdTd3NQe2WzT8UikxHXFtcE6osrdE1YlU4WhgS2PJT
mUs5EeF5806tymll2CcCpfQqGcdIC1rtnt1s0V4vmvgfMdzuviNjMvp8mbTeolRz
+SzJoaAb0+vdF0/Bb4kPBdGH1elU/f/XD9gvSePs2jL56ir8tAXhm+yjuQ7cQwZ9
x21jPqB9S5Y4SRRCNhERwM69XRbB6t8psgOrz6tqhLFUkwMmLqVqFv1zot/SXYau
0VfRNBvvsN6L417kZqqHGPhJi0kUZzcw9p4WM+M5D5BAE7jcI60peY2wvOtLTdxV
YOQXWJn7ugxr7ZOFFJvfGBIs/C2yx+uuhcMWppjxF8aorcNVb0aygD3EJ7QznDdJ
VkkG+xLwSiMcDUXg8IS5ajc1EQjpD4ayK7b7j7V54hffSo3iLuT+cd32oZ3S+HsZ
A9XL8lW5P2HwY97Z1KDJXc4bhgqZJQv7SKkiKFp60z+bUH2Gnity8dnSRpNhIFlX
RGlMW6uw9MDBzvIVL2lBs6fXNv0MjRQy07EoK9A7WS3+AzlnIsMRphJBPHJOgfkm
SGwljgW+ZcvU8ybBNKABEbKmSeV2ymMugI7+mbjW+JakhLgT74O0GSZMzpUUV6V1
sVYoXHn26Mc0WIGq513So8cum4GmzkuG394wYt2x56aFYXjN6pH3bGfHpMCPyfjj
33ok7wD2Row1VW4i32Rig1d8/vDmIqOLyyoQnI0M1VtUIWlIRDnKEJic55LR876t
c1T7rl043eVXNbbdcexPokefRojtsI0L+Pa0Wy2dhsfY3uWyNCJ5T3aRTMdQvSn/
QqMtvq1oKgCtnzqxdqDHPjbkvTfkzcj4nxQrIDRbYiGdpjIJav08yeCqw1AnNS4i
FDApRehcUSzp4YAtju1+UsIHf5GXflF7YsYXuHRCiBk09MIOrMJOfLDrabI5Kw/h
/UTaqwUDuz++fi86ngjEyv1uct8QRl0mimIKQj1m/6nbURHl4XCsK6r/XspwuJ0R
24AvuedaC2vc5/asuQcaE5z+E46IBd9xNvIki1EATBJISuhV52gdbW/BAVKYmibn
kw8Z06ZEocZfm+wUR07vgk3VZS3Fff9jcH7eP6MbvyAaaubFEaMgUsQtKcbtvOUf
8NpYQQIKzIyhXVq4PnVkUoS/5QLGTcz22gJtLleHq/M4ygGaoatHfvQu+xhiM4X9
065hmK5S5oaGGQFVsbhmiBMl6cs3XGwaMTVU+JXxM2ntcWSZP5tVjvNVR3hs7aBu
WBBytGMFvpLIMSDmwkjWj4SsauGzPiFukWZaAoxA7UHyi/bu4VJEzcyucxanZQ/j
2MIPlxVbfYYsX72XuD4CzOMtt8mxb+Qo23kZTjtw3cHXHWtt2ViOtGl6cq//Uje6
GXNrUYJIFdoKZNBIHQo0FdC65VgruiyvZmcYOmmogx0Nc3fiu2zMjkUIm47gFQ4I
wl5Fzyad9hNTy5dGR/6ni9YxIulX5e5SPlXYVghLvOEMwl2FGC10Omk2zw08oepc
OGzBg5JePNI/b77sjFEjmKBrnyQ5BgOTNmxS4jPVrQUeDC6U4h9VajnWxD4aOwbr
/IKDG6nbiZOsJZZnG312eIn/bULkyOU+2EKYNubqYf+xiSYZWsRGR0Ko8FLLyfxw
cInfZem+nOgWRfR1b1u61Yk/biUlUHX6tsQjgWhU0+k51PAznsMo0MZYV6ApN3Ll
IicK463HtZSC7ARPIiqnXvahyxDrtvy2F7Xgt56TqDHopgYiaT6/2ISgdqDtEFLg
WND7zh2JsIvBVAiS7eKGqQYdflxGIy0rK5+ZpbeEH2U3IVVgvOnlrcpjskkphnXd
a1p+GzHHLCVALw5indLRfZaR1+AcjWupoha8stzyScAoFX8EWMp8hQzQTywdffXU
RRsmo56a1zOXzpn+GVQ9mKBAqLH5xo3ohAWpadiUtUOjHVrjmfAduAaXs0tr4yxr
zEQu9Fz+dFvfqp6F13kzCv3C3lAyq1tAbsRnLpo/TZrFWE5rw+dFzBXWSyG89G67
OVWsdOgCB8XbGdnNdLtqAMbUuI4uIWOIJTRxbumGOV7CftebUj0n5cXKHK61kgqi
O+uCZYH40R10YxvWaC0eYGqsYjEKahouEY8qX9igrkHUxkadpufF7BnWl5X2Jqbg
vzseO3f94GflFlmf42nYjrmQsX4uIKd+wT2TOselQVaEk5ROJ9Ii2hdhrw80XWAJ
ZKewSbHzrevMrqGpfw/Jx+Z7ynsPO3RCngmeCitfe+tlyVArS2W8Zc2O9A//ccso
4CEI5nw81ifIecr/51xa8ot5crl+3+2kX2U4F7HNRR1qv1IRPwW5mcKtuXWe5Z3V
Mhhnpf+O41ZJClna1dqXwl89qcpA1UpYf4tFCg+hJm2SdU1Cbv5l3wiNX0OEgwkr
sa//hMmlDxf7bcGZq1EjgvMLP4Q5OKT6+HG2cKRt3PC8aAxEJzYULreom9bEOfpJ
X6BusfV4a/OML2LfqTM7R7mkkevn1QINxjFDk+E/XAP5IGq7vNEd2bb0X44j+hMN
k/zpYY1lO/Hka12fxYzX3deqZSsNZhJFFRx9rZt6ju5xUFaQxvf3fRBnin06A12L
ClHT5TwbEtw4S3wVexd+Z5hIHq/OJF11Yv9gD96xoueM0h7jrey3kCGZ17JWBOjk
2kuPOylMqdLf/0Utl58Qk6SbS7uf6iMXWGu0Nn7b5bzUzJyfSxckJb1+ihenGzh9
KRZ3CEZcUjhaSnnbXqE1CXLa1vOCs10x5IfhqIZ0oOpXpOJwzGD2D/Ngzsl88/Ge
+Y8773aTgnEtuHBJjPuEg7NqTg27EcubMsvOwijCnpa0TdMi/hlgWrvsIs8naRT9
MvZh5BvvSaOnf8cv/lWRb7WMJvq9ks4walnWOpnWNh364riiN8c/gYCVdTpLmUKW
vfN3mPT+sZv11cDOwsqUWoRpDIIChGmpbAP4xRjaS0Z4mKb55bi69tKcp8Bu1qlE
uOTkY3iPnRTJ4/k+FKFam7JTcP60RrSftDvMukCdhTSpReYAX1PthWBPCFttVZZL
8Q11Is2c8WRbdUWwnCV7s3O/nKNqwCgKWv/Y8BCYZC9scB2o7a0erMs6meAebrVU
9T/MAZTzg9FVeJ8Wlur+hboyM9joh/6zZ3dAgvWBAc99GMGnePQgnFW8FzA6b5ho
HJ/8iJG78Px7R1gj96xWkjeSjpXckLxd7KHSo+hjXu2vm+nIq/gRXsAIRxgeT2eZ
OcvTzKV1dyjEjnkZb9fyIoPpBuwNAqOHXsuGDwVupcbjJmCDs5qRBqTxNX9L5vWU
KbTrOikyryhffY0sj2ohkHdAt3yPTaxSV/yxh2UzmYwF23vIa/+8HCD8Ld9zS68Y
S5IzW8WL1oIXBqPqa3iP3r9OBFeFXyojUiMtYZIRqKG3MV5ix8o7eFNCWfgVmpOT
xBqQwnvwroOyeIubU0sQwtCinzVVhg9HHwOVyaJoh3nlnRWq+2wf1Cq+nOqMjhJ2
6AvqMLSZ/uD5aC2mhnfuwYsPAAW975k2pQJHA44PaY3KjcA6peddVvyuugLD/zdH
KNq5TDftVg4HSjTC83fUXctRkdg2oVu95YXgzNmGI8MHetiBRViAvFiQp6IB0Z3P
yhkP7lAR1GtxGagTVJXEbbeqMyidrg3XX/uCUHSw+2bl/yEXAfFiPiOFsilHZkte
WFwuR0HnZqFV1CxcNDhLYSYE90AWExuHbMP7iMqi4YbukInvBVuwbBp6ch1C49Tz
kiuXy5XrTyBcRdhI+HRbn8LnCuDYbrDKxWQwYG7nEN+lrah8AmMl1UZIZ0/ENJjl
i0G8PMGkzHgMtceGRoMvfXinxzUX4Jng/Jby9xMhfWPSmmbf1Yonvz++N2xx4rg7
4gYdt1PtoJ0nGN4HbeyWZ3/wedyC4Skc/8HU2QVDpLEGlHY0kekSAcFfSFUHoCrd
xyqkd7uFcU036EYsICBqUEPTZ1vqAR5T85UU+KlcUBYolqBvsvZPEFTBMw8Cj8Z3
g0o4ErLljtzT9QXXtZAe8sApN3f4Mpcc5PV1l+FW0nN6balyiIp8i9cXR0b0LORO
jSzrNiQnLBWWG0F0/OGN5IJUbi/XGj/e+eKSEc2ND8PprtsSONk4AYnnWhu9jmgs
bRTrav4amIM1JSnHBLZzWrVfdwAfJ9oyXURMdp7PIE4lJg2Sy6mUQCUguWYd2rzb
6R4Wz9N9sqIoTbOTnhdrFLf4DkBzc5br4rjixSNHBVihW5M5/4jVogEFxy4Szcqj
Wuji2VGGQLMTl3YxF8vyT3PPGr+FMwh0FHiKO6xHtyvLq5/Dc4u79zjwv5tKGXkN
EERTPhzX4xeKdeOaEEU7Hw49TzOvHNUpsWDF8NnO5KgRgSOeLq8tRYb7Cl7rWyGF
yH15lkoQ0ld+2x636oxBIIU8jpadhfbDnfgypj+xBZWip+ncyEW3cgBjG8Qct5hj
k8G32YY9wSgzWxfo7cT4vTZbhdRX/aPf88y8sdrGoETWrD8xNLMeU1kJTrOISU+4
Z+E9Od3tiRNSoLkA6BzADxRO3V/mNl1V4SwNZXsRYFTy7Jqj0krn9ku6soMvrs+F
as539OAPwtKuwClzB5i4pM8xgzhWpUZ1aEqDPnjXLuUiNtd7MdqI1b4LNiZOQsgY
ALWSBkGTB6drFYeBzL8SZ0YryXmuQrHUVCA2FXr9gScDFWj3MDGWCvhP+GDJ9dct
pH0UREqyy4vfdh6a/tKVUm6iwa+CyXPs7IdoRRbmonDjFS1/eSNKNX9+9f6+ipc3
fgacHW0QcSu6X9ZLcdxNsuvBZHLe/6TUdCi+AD0VOVKIOE4XI7CoobHJ2yxZ8XKp
fqAWbkE/CY20BN1Qt+DS9Hw7NqKpnEhDN/uJBJ2S9qETcif+UuXr4sHZKxp8JnZ9
pr71yqwy0alOesFPfEO+nfWggkeK1atbji889L7ayuf5EZupG2AXGKp5Q8882UE2
pzCqeWdK1+yEmspJsNDALG+jt+nYfiWFM7aMpVcMVi1GcB+lVAoVtObjfcMxFevK
fKXku9LKw2AI9MZt5aCGQu8s2wwwHfiAgsEiOLTsH86t7/sWuiytekn74PzO/wDm
KwqWb1awDnUuaK9Pp9jA8lflkLOazsEOgMLpItPVull6DXmRD4OWIImIxBoYdl/5
mHmDGjYeEXwqYC2daighYaFj0mH+JBTyzFphhbbIclS1eOd9oAlfdTxyoq80q23O
MeHZ9F2u12KQ9DMXWn1w7OW8BsDVre6KZoAlxzL7Rs00b2b4DI3wZncIVWpUhVmz
Z5622lOjZgIwipO8dbU4blHcKUt0Kb636rreBmGYLM8pIixXV8uiKMsJPvUjZZat
0/8jxid5SamNRCLpa6hw/I/sndIyfS90eQO8acvSaJr5sF8it/1i3Vy8fKStldQD
Ie/Y+Cx9KamSPUiBuSMfp6vzlKsSVgjQw0W62CLSnwzTP2YOZJI2qkwwNMwCOoki
LRJmhBIXBRjI0dI/kMcLf83hJGBzqTsf11z8PPJLd0Wbo07hrIEHb2WLaiho7N4G
/dfJGgMGBk7qYb1RW01oxpRosbYJ+6e0sVSKOWSM4UcF+Q6k9MGpQ7mHXLPBz6Fe
lCHusVmfF75cMGVcuyL4av5IJYtX8Ht/oXvpIRDie6G6uU90aGow27Z452t+l1aE
zWMoFHx5xwHDdaHGCV6TUeF6dg3NmKYUWa+20SI668SHsc07TMrMfxWj0oxqU43T
y1YFL7ppDb2F9vP08rHO2eIlf1K0SlcOM9PN0zFT5jVlktB1iRp2Lmod3/4GwwDl
Xrpj7L+//jLeP3+tEbZJXOAOsfA0NSZtz3CTmU7kXnAxZkq4GAeF4ouJm18anDYn
qXWYAGkPjQQ7n/BB+iJY3pt7RB+i/8afk/avR3BaUrJYhbqOVrpdx5uyrv5rUAPx
+2kjdmJoxp5njeDQIydH/Uz7/PX71lRlk3XM5JphdyZTjhhbwE7qxROfkACEGstt
DMkyqUsrUMOAsk17LsmuZ+LFbovVOoRb+FNLwFGM9sjOvIMDzKDJmiJUzR08xHT8
jzj3Yuf8O16T6RMglqBHqKcQ5vW1WuELa+V5bom930Xqep0f5nJsBbutoKAX3Flz
9E8nTx6a7wopox0JlaB29TQactS9FeaDfw8GVT+AU/vZFCXvPnajNAaT9E6j9np6
GgU7vmq/7NQwLw/+BBB/E/wmlRoc891Ro2q6lAwGRCVJM1fe70gmGPKmn4KEN4GR
JXHq3r4U3WxQjH/5SNc/35ac70SuVjbMjEf9nNoOh3D7Dfy1Wv6QBiJ0PazwaEP7
XsZI3aGR5Ws6QVkAFTsCk40U1Jk99HE61eGux0vTLrioM5zfuGpom1Y5jINdXxkc
RIKgceKc1lk1VYmKxD2eVodEESleHvwhJ4c2VUND9IziSmDHn/OWG3rPUlmvJBsk
wJNjvOb8CLEQyiV7JmDrnu4360X6tkDvE1eNFOuhgktixh7WLGj1npbG++KEA+BV
GnZFarUioxOz/8DCyP3Ax3rNMyIehH/vZHy24In4oaMwl1jOEWPm2HKqQPJwvWhN
UWuJXrJ/SVyxrdoGyf7JKTlDhlgbfLJTawQ36RbVGpTGbwJuIeEy5WU2uN3iRpeu
DOsY4iwr2MXmXJrCNlzyqXT7ZljNY7nytLwNyGBkwDwhIyHGYj9P/q5wJcZPAJw/
0pFOe1X7jq1kE6yxCRDKKlt3BSwNtikO8sBwNS3v6byyt6nInyyHavnKvlV/PC4A
LdWnv8dIgevMve+IO6jY+jvc3mYIMoqCsfl1mA01JFUbQ3DQOynb/LrLNtrYt7n0
XPCd52gmuTzACzzhHNsaaMBBSjvEkugPL4YbFyruNfygAQ7CbLhwrG2PtUYw0Hej
pkNU6Rd0uEzpC6z+0CsVov4p61qO7/70if2VY5eH4UAdXqvO7DrYmToypuMXiSov
Ps7RvGB/Tx5qlL428+7/K9/LRT0sJLsmEqc95+KrR6yOjjQU868qx8WMGKNC/q8R
zhOr3pSKsIDpkkA7tt/gGyieTOoCFBDtJY5BmGJfB+CIPCH2tjshFjNnM+ut9Hnd
hpkzGoo5JT3MM+v6s8C2LdQWCxK3IhUbPOwxYJTNeTpn99Ui5lIC3AoIlqvZ2QFL
WQlCeb0T7h2zTEB+1J8lHSskCzuQmrbNfR5Zj2vuNTTDiRy0Gi+8wbvE+dSwxfnw
G2KyL+cqkjLv744LhYmzldmf3fRWUgi8a4V5Uo6kFxIrkY4v+FTcFiWBSgrWCo3b
TyTq8XL8v+x3qG9lG8K8N56RhKHUMKSePJTYh1YTGjr+uTogeIEuYGmezair2vsi
QSnh+0tyo6zLG7rQNC5UYZ2D8O9eomzn3gRTvZdBbLMsObwj8InTmsmUIHU3oTyb
wFBDYNcDQIs23fcXAAN8vlKyuS91KT0jEHDTMK6q8COZ2ILx118bBLCBMhlIXSKW
wsYajkQwJU5e6SGqcivCFiZFRkpN5MZkEtnnGbYa+Bwui7TXfrIVukYL0K94HmID
zKGzsh8MZtyK/ndOL/DhC3RJrDrQl4G/YDZVPmkboAVnAWOxuNNxfoY/oTEQTbD/
kWr8l1PDmvkOulx8CMbt8ZylnT0MNHlU1eFdXwdGrb+aJh+DhWwGlf/FEhhFEu3A
6h2z2XusaRIqWx0IC7kjjw==
`pragma protect end_protected

//pragma protect end
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
XJqTy8sL5MBr1uTW+vYEssyyadSaw3inGNIp4ob8DNoqbQYN85bPa3H94so8Jnv8
MrMgTQ6LcF/agI3HNoMDQ+3ttBiBWoRhPJSzI2IW0YF18pOLdpXopiurPCtSnlaz
GrV7W6RWlp5/cM1t2vY3dj3uAZ6Tw0ZGoWkREom36q7pJ8GEY66NnX7OlfTWp9vP
4/CAE76q0kobiwGbWjRh3ssp01DjszU2O+tWkE9deeLUZmaCriC5f36ZOFpSKkNy
aX1wm0K6BSgStyWZz5wfwSI2Sbqel3TQYk+cqprcOPJPoaeqQKStw3ZzkpIW1TXn
SFGyJgxAji8U/YfJh/ub3A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 14480 )
`pragma protect data_block
Bi/5Gam5I89ApYHIpYtO6qxfjEpBOgKh9RifPSz2CD0BJ3BX2zFpUvH8FTK7TheM
YO4bgohclGgMQ7fj/WZ0qdyFRIu2UuVwbpAjFq8/fhUmnj5nMKTtgAyZTdzGHnrq
i/ZjA9p3GegqYbVJEQyzBBqV95hJ19AwepZTlRChQeak8O9qAO5ZSyYKa3iwZq20
o5yZOHl3ppT+vD3GO//2YVDJBaWMGpv9HsR4qzqHOh2c6FxRwtgI1zmk4Ye9OelH
1qjjMgXiTrIFckkrv3o/dkW3LptzAEwh3s5kNS5gIDJbe5anRXauna2As3L2Gb6Y
cKkn+MR7vDEmuQAJCSp7N504LE9oSY8Pq2cY/qo8VccZH9O659wQ+G5UIaabIHXd
LS/9Nw5zEE0QBNUiV0A+SG5itAbEroHM+Z3OBb6+ckUMy9Qjyhf8dXL6NimiNY4+
e4O6XInPAjbXyODdLvI505O0xrACQtE+xcfzvhhpMd3AiNfxLfAuVpt0vR7wwvOW
qyT2nc7ZBiGNO3M2C3zpPn5aNoR4yAVf8XRJSNrjXdVPj69VwqqGOxWDTPwPENxT
4kojTlRIrZgSEMjZ48enI4YSe9ft0vQGBtjs6rX+Qi7Z2MAAHcGXOmDuJ4Bkrpb/
Lp89qiHIn/98OLsOSjWXb49DOKCr/0L/OqDKEl7MSHHm0Y3ZsR7brkf+Ojpjmiwa
b2mkWpDF2gTVhu2+0Wuoo0MG/xSDPgCl5d4BuVCJvI9xtvpKNGshSKKUpQbSmYaa
8oQzIcXh28/3kthFPOlTUwJ7xCpyQhvY+Q25+tU1vp1G4nkTN+oYf/B76ZhKxh4t
7oOoO+grfwSxHMN5/xkhnYpkeaSmhriLPPRzPVcY3Ft/lGUEh2fuyZV6s1IVReLF
lL/tGqWRXC3piOOp2IhxpvzDJDwFTHTRDMPHOzJt+Eu6cMwazpsPdaXKPMb1buoF
4dV9gLRA0wnVuWfMUKlL6GTb11SDzATni2wfNivRYnxfeat47K0T1bcsL5MlIRq5
xsPEPyUajJPv+XSCS7zvR2MCcFSA3vMjg912OoixfGpKxGyAKrs3dIRAPDlO00nY
VAo+qX0vtVWs17RuVyTdLp7mcV9H21TWS/iICKVdxaJ84rnHQIL7yoOJqqcBBxlg
L49OQj9mMa9yHsPRtu+Jwu5oDeqPu/Qn4LMuvXECgKu5d+oV1KiVPs5sEe+r4wHt
NVOAdRxCMJM957mDIevOS6jp6uZodr3NQKy/urbTrYK/UY30Y9eH5Vvr6B1kivMm
YgUDUJYt49KrISdQafGMRCw/rbcCYmzAkPzb+Dfsr5GcijjflIiSb4O3Z4YmQdv0
EoqUasu45W5AmRNARpcbUdeMuTB5/mxpG5yJYXODoMv1/ZiSeJ9y7/W902UKNtgT
YrICwwSiH1SBaKhy4RDY9IH20H0OUYx2Z9k+KPVi/K+sRn8SM4svlMH4afzU5zVV
95WQfL7sbGci2f1+DzdRlQwNnzEu/CLCbUBh+/2WxsnHe6q6niuLbiAgnodEZrG1
1ZVQp925vpYk9wKk1GJkLCqhsmkCo4XME5CAf8HU2f11tZqd3QBlg+ZzdelQHRzy
1WHkJQ3e5iCegdiSP7Hr5MF4K4m/dCB3EB/w5pj9MIfsLk9/0mzRWzIl/DP7pUlY
FzejN4LUcRFBjCIP3eWdXraZGsr44ASQkdRoFfuROQEndrYPBmzqvDSRTFwJo3rf
aHJdGfenl0n32uiHod2zbIYXNy7RMOK8arYTWFGAsOEHrRDWVX2zwlDeYQeTMfbN
MwyeOuefyXmmr+N0QNyxlBD2gdFeXtkETrj54hSM7XMJ6DeVo/Pq3b7JzIefqQlo
FQzBt3b2R32SHUy1j/HPgiPVxR2LbudY6jGlo+Ce4RqjfSbyN1bHeheYFn+NKXm6
VOnsukAhy95L/fwHY8ox+owbqVyX5OFDHCNFLNmWD1upJt7PxQaLIyWSbhmLYR1K
UkqF4dr/ANcly9PiPT0sczq3kSVTTNsppQ8Ueyg85PyxFUeM0ru/91Q4JVU+So6g
8DHxWDMwFqZYzVmQuu3DZfWL4piuHF01qcUwl3a1X3tBQos28pFqr0lDSIolY1p9
lPEmpu6qMaf0Pe5AicCxs9Y8i6d9aL2P9OEq3mrznupmm1ls3YYAaelnjljkVHi+
rXDaJZnyzBSQZp5TrTp75AfTxuhg87VEJ2Gcl9i3opj0ol5yeUw1hs+OJCxeiX0I
MW1oPZEwa0rClFS/HPeY3LLPKD5tN6E4ZxDbHMBbDf1T0MmFO0RLRuz4/+vo4JJb
vNOJVQI41kQfQPUH9n8lEoeoPmi4e6eCMxByuSl0iidB37JMw8lTzAFW3XvbLNfX
QgcGj6iO7ySCWdVVUKKlvRHn0LXzHG3F/J6ESCiPHTfkt8Zf8BJ26v9RqocMIFPn
xIi8ieU+YqlS8VQGUEYrcShYGmeWnVHlaui/qzC4Kt2MLp+HBtQxAC1jT1hNMOL4
pME3MzJbu4Ufw6ZUes4Bv4uh+Y1ryXwHVlHPZPvcXrnOgNs+aPkh9A6Y6E2sar09
5TJbJtYJwu2nvxXM2NV1jmrtJ+xv6f/MzNuv8moxkp5vYFU5Aj4P7vqAUwj8x9Mr
RgsoMfQsT8ASdEIhjGtEwTH7GT+iDgLVHsmAa3aynBUK70UAaW78fYhK5WxGbjxh
d2TVLbunlqB4BaMuY6ZysQ4D72Qnw2Vv85viyDSwKtZ5kiLKRjju+56uc2KsyL6e
ZHFYBYX+9uR26pI22q0Dn8c+ZbQ/GSxiq2JQPzH1SIjHw3J1M5BmJrfueqRA2Z4u
okDEPaCX/0hbG5pwLucDY/zgcn2kd1p41l5d/9fHnzkrGN3CbEqCHi5a7K5Wp79w
EGAk5640o54wcTCr3O1SszbKQBkzg1dvCBVhXnAIZNyIGmgJm68CbtxRK9wicwth
0/IbGL2bwvT26EejmbET7ykCAWUuzCGuY1ZA5FOGxWH/enLmIF1NfjhZC69AbFOM
5FhmE5tvTaL5F8h7ejREFum78VGO1rH2hJoaO8WBW/2q7D4on9gniebdDmf/q8+/
jtc+1z5M2GPbrtS3zJ2JRGhT3q24cLZZc6SnChSuJVTH8L3BPz5GwehcikIomJ6I
jQKlvkSc03kwMyUh/191I18iOCg/HmGQ4d6v72MH5gcgn2XT9Ud8waXbQBEVjm2y
4oq+GVJ/SduRNabTZW+BWzYOxg4R3kRzBTSKYEC72uVGNNvSHwicyZb/+CBQLfoF
wbZ3/TU69rf2lcLPyPkSysOJzRdkvJn0+SL5JtNHCmWm5sUbOq4BwAqpSmbRwypG
Hi7mcZ+ynvv1tdbdQlcI62FepC//JSJ/NgAV4AgIb/XIUbuqh2sX8pPNPtEQnaC7
NSE2KXh1N7agUQuJpDRFKBLZ9XJbHTAqOkCKQ0hHQ+RKmvFYpaC3LV+M3uT0QBf1
T7Le3V259xFUEcQMWHVbG11XMBlOSp2k7MPJbJ2Ea2EEw/HAjunVJ1aL1gQ7h40b
Li5rgmSneRUAoILbPfOloVlDCHCuM6WtQCFBx6BBCKZV9RMuOmgjCdMxzHBTTF57
KEfvtZrO9mlNISzg71M5e3kg4+asYU9wYAzKQ0abq8y9YLMzQZ6a7ejq5jmPs/5P
QIbP7kLj/5O/vXN86w8xwBAzDTU5fkQLY0XMCIjqSgshr7UvHOLp8TBmhAJ90Dlt
wDkVWVFUPMMYdZBFHJRkkvPIP8KCu9nJUL8sIlWhiSvJKhWLXmpcl2cvkabSBi3V
g18YOIbMKOZFdNIfFE0rKnOtUBkZJVj6rECV/k7P3tV7JA6PijT/U8+9BQLFlvyj
vAxs8ZSI3dhDZrj94lUBQAf3Ad+9kSei8jcLmTAI0lmBOLfQ4t/xDgTCwuCFjxoY
X76vcC3te9W29VtHYeZWTIvVq/QCdiOdEE1ikE55+vf2Eu1PFMAybXWXCicYA8Nl
2wKDuYHla+NG0YirkyLr2GUF5mze9fRfB2OnJV4r64BXWFqNXp8ne5e8LHikhHbX
EgrQ2BZOjcDJegbQpsmAUewEpuAuWcm2TLVpceTXxwEo8TmylU4h77TwVSX3bhSE
3hwNdIhlRfAb3c3HWvsfzU7upnC18D3ObOXWg0NFB/vw8PT8C15E02nG5otDbFnx
dHnKwpaBXAud8SCigt4OzURUWlolKY7eCEZc098ct0v6FCnS9TU0tXitmaewd6x7
8+QoKtMsFmZpGTATOy/z7aytsIdEnk3aKNDGvKVw4wbeSmaIYEFXG1a5lYXRSquc
+GNVP5Z+rIQu+VK5TX+vc5IxYyJjyCXmEq0q9YG3BiYJVmwsho8Bf+BlPS6B7urX
e1gPFX8He9Yc6flNXd/AqkIzMFpiNNHn40aPo3i2EFfGltKK1nTq2s4k+VEkqp9S
CK+0jb/lwBPmn0Rd1HgAfn3A3PoBABxUCLqV5t4AQewNwP0NHfS7pNymY5eNIB57
kZ2/3oE0MgVn4pSVapOKLKnc9DaLObBahkxWzu300DUyXLPEDJvY61sRaWVWCd2W
M+236T2fOiNxXoSEua+VSCqUjC+F/Z4WgEjlJ+Lnww/DC6wmCMvLY7mRt44ff9+7
kNPUPIs0oVQxl3QNkMBzL6H1DVztis/zIlh0PbEdViz0pzAm05NKWOcwdcksxTvr
1eJYRnIpCVGEfrwmWtO3K51CrFH+7pehc3fG4MLAwKwrqfL6UL0psdKdTm2rQvcW
tc6u2KsG9IQBf/usSLpSmMiO3Gw4oo1anmfX3WbjeqlU/B2s0xSyY7FnSvcnrrqu
K8WCRaGqKDJO+bzZ963mkcpzLePTuho6BUoV7S3qYh+Gx0LdMdP8u6QO9lffJ2o0
8MYRCOoNr51SkhzSlP2ECaZSTkBgvpVNxGg7GKTsleaNxV0FGUPS7T7FVpReNEPz
QCTzoob08N1enZBjXDqLzNj9CJq1t1qcAhBULamMURl+6os/KC+P3xV+mEMy5pAI
QFXBVQmw5uPsh9WWQAH+m+l84ayEfVb5ZxyArvUXrUTMpuih3O5AOpkQTZR0L+fY
qV9Ruqa8uBp2H50VEbIW+9rzCbDwnEkNACEySS5GgeWcCH7VLsDPOkfsmy0G1djV
et+qSBVnETRkyOPEIXETvXvXVlp7EdcXTEzGnY36Oa4Hg7vffNZGfaOJo8vhjZ1n
v06gXL2kIdgV0hjjdz2X4ITDI36rclyevgeuXYQJiR+BCI9ZeAb7vA2JGxYSO/cv
JSoLMrj6dt98fjcnd70DFrrCELdEi7hVarz6Ikdl/5TLB8ohOjkxqu1ROQXm+xUP
22CGnTTEsWMTkM98gguU0LkEiq1ZotAqq3uhIJy2s6fNylpf8daAMqkLS/Nirc1a
4A/86LcacjeC7Dr2Wg2RRzYEVZzeoFbRsTudVfH0yuoogzeI3IjENQI3Uc0MldwB
gIQCKQSzT5JLiHBQv/sln8kiORT7AoFUlumweIHvlJbw5faLfzw18NxvvZIPrYAI
h8whWrA7CPWNfociUDA2jo/wXmzHvjW3wlmDBUgonHpBaS+Ej64rFz74f6Tatey/
g2xf1ayW6PdttkBm2lbG5sD6+DMeSCE/hbNrJ466soxF/0qaBoMqEYYCMcNl2UUe
HLzXe4Ca9vikn3Hg+N0qdE3PYI1/OJIVWkvbc1kbeHRsyKyjK/X5f9QLNBlvuxOM
RfEDRcAYOGRLRgP4k8ibszKrNeinGx83hT/oaujqCV9ywB8J1yg8Cm69MakvYSGE
xPPrH133+Ma5ms+sHcT8k5K+hOSQbAU2f06+aIviv1WmcdBVdw1ADYO8O2G67nDe
EHKo8HHiZkikpqClYuD6fIgMZsolEHVT1uPS7OM4Wb4Bn25AMZyPcQcMs2PlKJvr
f8l/6sY07Rgy1IKVMdIL1uVDSAr/xdNz6yJYHAyyFXuon/ju5uWIcjhM4cTuozIT
tnBUPjDVjtPNS6BVxoId3cAOyn2nhMu977A0gWX83qdYM74l8uiXxkUCKNAatjKT
MRx6R8cyL0cg+QRWZlIc2cHxk1Ng4YkciKgERmDSuKFh6Ej5EIdDrgQQVHVlfd/Z
H0zTI7E60S7H244K0aCW68+oZidcG0S2Oo4zjS614oSskUBrBSeOVeo+wYaxm9KG
WadeNiWTAbzjJnUEJ6Zy/MqU71uWhwK/00RGfYXEwAJqsr7GCbZbphkZ91aSclFz
nMNrVfEMfSrrRONaPcS8krN02ORLxJhE1W55Iuimn0FfzDkaDOnsjkstQ1AzKpCd
Bsm35escwtWMMoic/IojnsnMx/iwnWRwf1GNsJ1qk0jwY6vlermaYvzEREQgU+fS
1v0pSWFqGlPfN92LYN70Y4qaanc252RnSdlG3ex3WnhFRKFvkwtRPOFFPSFLn+d0
VJpXMHg2LOIKbIJSUI2YKmlMapOpz9sCfI5jb4Hib0xNygPnRrmJtLJVcOSLKGn0
FWv/AIIEMU3oDNLLR6Vo1g1BwZEjI03Fquh4QKtnPdRufFVH9JNpT1OfW3oc8kiz
ccyai62oIH2eSynKeOCgnx6DO1MAQ6bgk/KuZ34OG84w5dIQtWHCbJylvbTX4KYn
lJp/bdkMllozS3oZ7Kh/owUH/OrGBILuiw/9FKyDBtPvqXH/6d63gtxfEtowSevq
YNYBBdVHIlSbHFihL0iMJtbYQ1C2UA5HTNkShU/Ke33KOzlxsq84Mi1/eQKJynnO
4mYh6iAczr4tX3tDDYYu8bcrIA5vKt2n2BHdG0hqbI/WhkUS2L80LAx6BzHTq1MV
I2sJq6qTKPRlf/aBd0Y8YDUmLwYdoS6wMS2Tu9Xu7aRT+ZAHdjzL4TC+oGIxnrS/
LuKBnwWHPV28Qqi3j+K1y3cpAwl45zwts56jPHbIczPWReyKT3UElIqdnduRQN/L
0kwJg3OypxVPuWSJ3v0zHh4IbmZt8wbMwO8b4wYpFNQ2j3KdxX1si/s2RfBVYEjg
EIxj6/tv3huUPziU8Jm8iLT8oqyMKsK+u5+LICb2LsyMHIGWNqxGYtI6z27eUlqJ
VPg6Joq9GcMPHlcEM9sV+f20Y25q9ti/5nJEnRbLpamH17VTxANjDov6ryAFrfaV
Mjzzdn97gj8YNHCvJKrCwVM0/ki9setRhdRyniurr/3hmDxNhbHlBkIZJfSv5OcA
2nu95yKaTLEu2jAXP6r1pNbqOSS9kS+1hGaTr3UeQHlgkaba239Ern1SI3CVIzf3
tmmRYyQc9khMNKS53IUi3PShuWK18XhtsntW/4kdeVyRf2sOm9X0IZeTaSHWZJXg
yV49Aij/OhNQio1tReD1vdQzGYTo/i19usZY9DEnESJdSNwDhZAaDgKVgRsGTJme
YUQWBHuNXLAchW/5bBbPu2+7wxBlpnR+kXA70El1AFUY/Xu3rYh/7W9984xGuc71
tf5QK0/5DyRMZ2ixqB7qfQlzU/Wbs2U7740pjWz/3pIqR5Ih2dVf+Hi2zgO/ouLh
6EiU8RU8bPLRMjG5TwuwEZUycLFJtuyejpjiM5Eb+yBihXgGl5I+80SEsHxaiPR0
Er+PsCao0JjQEuXAmxQIeuB6qwfv07Jkd1XU4JMR/XPFZ5w8eVsBXLVU84VUF6D9
0tN/VXlp9wsScxWCFqznLekIxCYJzdiTj97D4jYnMyRxLEqCM23UMPl9Ihg7JqLn
liG7jOlumwffTAMPIYKBHe5wKk4xDkI2lP0iyey94mCwUfolw/+guICzXpR3Zdff
DggCfMrJaPBphEdHE8FtTQw5WiJRuNjNYlB4kVT1v/ts14egtHez9G4jIsZZw/k7
2tBzgHjtoNYX9/3V7xKSJxgbvrWKie1RIXvWjEm39LJe84wWbaU4Aa+W/6GxyoDr
Nop771p+o4ED7HnVwBByTBc2J2+4CKRHgYvtxV8LpjGxMrXoHi6OS6IbsemQqx8i
P5yOn6sROObZp4DpaGaC09452fCu0CdHwNQju9SAiCj6NsPN/SZ/wJdjj4W5SFD9
zK/fHdcwv6jIe0snOQvnvJoP7HaE6y5cb0/K3bw87/LbPU2poF8VvcSBZCby7Pkf
gNvD+FiQJEmyqhYaHXT8V2k7BdoqDjS/qbp44abmFHOsHpImYjseU1bB9LeyZWJY
T23NqXIpFQefwojD6bscpNLEtp509UGYduTbB7lnJ2A8OD5GU6CvKAu10wfAnPMB
TsSSxSwfuuBht6lI9DgtLuqAsWnoE3wSbQKiMkkllUc0opiUg7uerhkJ9Zv7xW2c
JLRFScrr2AZMU4kdnck3RWp4u4DdBz4AAzLCnsmW6MKgPBnvgFGq2Mdi7ESiw5yo
KuvXy6QHu2/ZN1YZ9ntJ1CEPxQ1rHypARAn5im6MW3/V2k8nE8J5drnR2rIQq7hm
5SwMwKKPncDVz1syZsXpGveMwE2SfB7QtMtL3//EVE5epPzw6wWPbQ+0fthIMa1l
Y5YoYmL22VMPXD+eeZxn5xaWr8SxJnkLr36MMxcvT7aF9Jh+kjoBos+uOUvKAVui
MVDsYzvULsNy/yT5g3S6WoHFfYiQ5ICjCZY69smMm/B+PvioTjqs/Sy0/gikW/mM
M/rXCyNIOPIDNroYj1KgTWs1Q5rzRaLkeoaNTCZm7Z285KnHtrN+CC7C3Mui/7+n
BHGexSQJGZrIhBblhIkQnRv624DSjfEo96vf3jyyEtqBIeRZGd9LYoviRijaOUHl
AO8OrVbnMoV8ru+cmDf6wVZF3duKTNO37DCwt60KcwFf67ppOqp8ZriBiLjX+bL8
51wT4LNf/PvfFMIkIAJgURulFM7ZuLOqiXZ+JsjDpKrwi81w1DUr6EZYpBSJ7X0n
0xDKBp6hE/AsDUW1lMzYSgfnxlZQojo7ChRSysOnuQmAk2rjEBo5vDHDTyitqv6e
mT9QP/zkOKA/c4c7xdxwgZoN+vtzxnt2CRGs18YQFakzcziRpMmuzg3GHLxizOwu
j2m7iHsnzgUbYwg6SpDa27nRjs7qXcP/RbE9KTcFvOG+5EPqGyVwc8P3+ae18gZ7
MpqyvxOFU7BvOfEtGm+aRIuxdkzKbSjoMAVy3rZ51uXa3/kCCwH4Z5nPrpUj45uH
vba75+duWV80GWkB5G90X9Qw5bRYVzZsNS2mjyl3ysKxsdCmCeiVhDNMVEJQenu2
hplNR24gsjCCH/WX2K+TTjKPLhrz2K0Z3sbPIjn53CF/UqTy9OQMSmIBgcdLeHat
GFm63uLCBckf8ChvCp3dBFbaPBBm81DA2NRJse+NpJlTjILznoSvPyTMsHZH+fq9
FJ5iBvEE56L91Lfi8iM/GlwWlk9tUcKn1qj8MhEXXYW7mZqIesS9sBHXptXN1Ira
0eCdFcU7icJqTJFKi4ehljr22Kqvfz3N4quEAqurVHSBQ9fqYX+QLBd5pl2xyd9r
ZYrEYpv1CZATM3y6G3v+KSCI0RUk66H5LhCvGKMC8sbnmVi7DTAmGED7SRhObmNn
pNrkQ3Kbn2qOzIlPnVrlUK6h2Tep/vXZr9uttY+RaC+27gYnlVoupeUQA5l3RAPK
InECipcSTEn3CXkmjC8ZVCFVE6jbjpvUAzOvWFpjfRM1+pDs6A6VMbzDEbsJt+LU
uHV7EAN6Mt598z6cWfAlGTfSNDGgJK01JkMG8h6zHwCLZp4eXwV/GFNwVOIaHhqn
35s2vT69RFKoO4sroNkeV1GHi0HYkDO/XuwldapX8HpP4nnA2/zXXQtNRqzSz/89
Jdjn2o3h9UBogc+gReSNqYWD/BxHw+ajTkberjqD9BvtaaxAJugixQdRcfirnNXM
cZufmWNoMM75i/leo6XLD+Aw/BI7GrgNw9+QBLGLqx4qKhRbUgWTyfJahZBJgaL/
A9RujXMB10/PO8dfMWUFOg2TsBULb/q8T2JCkp5Q+jt1Aj1kGGWFgibdO37vX1Ud
RDuJFgYn9ZkS+WHkoeE9k8DbBkd/MSga+XYlzRSjmdq13Zx6h8/H24ElBm3a3lHS
e9x+hg9a7f70P2JKe0nM/rsgr2GqtKrfSOFXfFOstsA0RDqwxEwTyWKddO6HKxyu
OxN57NgdFCgF1ECHpMw1ZX4VLPdxdc7MPtki5H0yuVXdpXnqF0o9bexh1TeJTGjG
5XK71UZdy2pFiqMhexqXfqOECieJtU4remezGi8cLzhYfPa9DCYP1MUZc9SjDCzC
tMUly7KfEt5TrVxRmTEzWTyJo7G8ZA3C71WrGHB0P4tHPbggaRkk2FU2IiEHTB5e
83TzWwcd1JOBtsdi3rn3BY/2x3DcoMAzQbdTY2SdjvuT3+ExYP7wcMfwg+kuqzAa
P4FiHHYSt/lJ/jaXUN7LjtAdI76pwwxD4Mj81d74caGL4ChsDrLi/3mqnD2/7ri9
M7j6UKOi1LAQDXjbcamDM/if5O4bCzM+ZODhr064VgnEjFD4ZAszD6Hq2t6U8W99
tWd2qtbELmvtDrxr4x3vaOmx3o8fZ8yk5CwcnysXHRnkRckG98hlZ/b6ixSsyihW
CBrCMMCOagPSTmtJrMjjfpydYTwLdrIpEUMB5TXWRTP8NPU3beaxKjBnHtoQMVaM
Sjv/5UZYNAOkrb1dqnjtYV5Sx2Ax/KhlLKfR6/YP7lOzIPQmzcp89Vk2I7R4n/v5
Mx4J5OnU6usQ9VXW1g2Ceqc+1nxLxD74xENhrLHvmnDPqHVlLi+2g7+vU6S75UYz
Tq/SFMKdFhEuU+fiRdMohYeE+oejBC1qKG2SXCdX9Op1KX4GvqwJaWgKv4Q3c5GV
XlXVs9rMTG+Vt0kYqdrzEWCBLF6vsjWfjAlB0CHVqII98S3eocg9ug0bQhOkajqc
olOQ3NT6VI7OmCDQfDU/O3N1KhCj1WWQthlyZUM38W6OQOKPaLtdgwSKYXsk/r0u
AIPdwA5Rvz5g3hR9q4CxCBVXIOkcFRMNIYwvSzbHou44ICdo1zNxS+aKGUwfnciH
yH0tKgDhX2xHA3nx77CIFZKtJEgNskeQSCdB+BWxTbcilgefFnd4iBowB5TYpBLA
I4QufghB9mP9sng/OPz/pcitW+wlP3wS72eMjE0gHb3YDsfLRyia8V5mC4BLsjFw
b/Hrfv40IqUZ8yg1sP6eBq/CgDKO38MIrtC5SsmYk/MDwwxHESR/0kxk7fYbYSLP
SJASYOVTD8N1psvK4nCJG807u6bEF4Rom/FZapTMaVssx1eQpBKbnc7Dlwwy+vkg
NQi15ltXAQpjlHEAjWYalR7YZAvM3GhJ12xMkyTGzhWNTzWVXcfdBlTWl9X5sLXo
+rZiCtOsISohSIAxkUShY7TPo3Hzb41GyQDZfZdgKWfQ9XQiI7oHh/x8EskXH87z
pFkuSdMtqScZsf0FgyfeoPkvj/7hcT3OUmgGSkM0U3UijkcynBM+sVTFrfqW2627
veXb5VgW01kIw+ZTrx/AHrLurorHPgnttGWSDzBSoOvaAhHz/6dUzH+mYolIqiar
VeLOPix4Qvpq0D/tA2/kEhQNSVC1BDZkJnDqgH996Y5CBoOty0VICUfShZKB3CCE
6ygYHbMVhktc1rgyPC6LiKa7ZX+a17zLGjcIVYxa1By7Z2lWPhRVySFySvcKKA/d
V/pvkQBQH2G4EFtdSkQQtQRDjy3XGn8u7Z4CosayMv6QcKjvk1iTqFPEPC2z3wFh
XDHG8RbQvtm1cPqStlXU79zL0W9t7huqC2QdiKZ5pkUa70Scq3K91cNWxPOSxBRt
Sgu3phJiIFb5uzCy/DCgfzZHr+YbxQuoVszOP9krDfApseYgN8jyHLbvf9IHZC/B
g22K9E5vl1BFOiaT13I/xu8f1NXhCkJi6P9ZFzAQsMt5HXwQNTVD7pRHDvFftwMp
qDU04yJ/8JCYyPLWMyoaEHzdNeSn8sQgQWdfsF5+AUn5DSJWbZPmjSTXWi1q0FSm
5l+4oHsDa6GQImHhEewXCjJOe6PaFFp//G3KEKcQYYBzRwjbPvDkgqrDieycdMOw
H31cC4zR64wCQQBTNHWklvYFZ43oFpxQJmMgnLyLfGNZGULIpTaIViGjNmpToOkx
PMxnSp0xmDxB/UyVq0CzdxQKHNJKKsMfMczWpeaqAL6Uqb6frEjDoTKT2Ej0ol0t
leftkrTimlMcVGr8wIo0exrrkoyBh8c2a8jktF2ZipwBhaOQR9cZtUwOBV69uAOc
yNvGxzZutBQPeODCm7NiMa6q3AUjkMCW6uPOdIKhi6HnTSdm66t4D/VvDS6fmW1j
J+Gdh18uvn3s1Hgb3NTSwsNDjVDpSAKDOUygXyE5c1IPTzRqEPeVcd2NW+pILCOI
+l5sS35HmvB2by8CsiScJ21BF8f7tBhsMXxQtxruZQUr0CuMOwn5BayjcCgot3q6
DamHFcsAyStERk1T8flRpF5G2+4g5+1jQ3NkIgn97/Oi3mHvtFSdKbGr4xGzRYqh
JmW1dT5OoeNezzPEOGT963EajxWKWtedFWBX9uiIxPCpiGPSPuLiBWDOKcw0h2h3
co5mL8nU8spSjfAN3FgEtKQ/2IaYoGJAjwaEbw46Dqgfv+iZ7OFaGifRgiPJcolo
ibFvXFiOHWF/Ttxjm5+GbCYo+aWQPryjbAbGIJzfVJ4zmda4fzR70g5I9idHDp4X
cCjAtlDlGoehyWRIrQD0Bscb3ua7y2kKDsrbt4iUveOqQsjX02WzNyw7geePugh7
HYHpKb9brSYHWa0auTh6BVUA/X1IgUCDjlMxgc1Kr4niCCGyYiwuB1m2CratkmMC
qJGryWl5luhNicPYRjCmTafoKPfRT89h93Zy6BxwGiN80m+hVeNn+Z/fgUSy1zRy
8meBVxcjt+0uuING8KLI4XSY0p9IdSr2T3oaYrdcsFN1SZPwyEZEuaBJ24wkS0Tc
96iR4uJzGdZ9Qo6GLjZO4fJu0c9JSlPmdsxgGeQaiJ/eejQuIOCvxycgJLoa4T+6
uQNA6uWE0mZxRuN1hO+L5BwAeN8aa/RIq6A9ZNpkHcM+9zNgYdxi371oX5c5s6jY
0fG0rGRr7pnjbLBP+Deb145MQlFDdLdK76UGHQKKvQhX4BK81OboEIV16WiuTaLg
pMWngVYj9x7sMMk25UIk4ggsVchXi45m2Nn4FUZ1/hYQz1yNmv2+Paeg+toljpr2
YuYb+gxgPEvWBZZn+yXQm0X01UIehIwgBc7Scqcm8ut13AZDhqMZlya05NxD5WR1
VFqeayERApHEar4VZm4NvrhhhP82ZCNJhYsgg9vBm+fqsrAeiU4OhTLMJdnY2n5z
r8NKdwaZAKpBVkUPKafIAoAc/CXaKXstJ3FLlqSONHkXW8jasWkc3UOlXKu8wHu3
9KQdgpuQ0nV06QppyNGW1B0WviWpSxwv24ZqU3cvF2Llp6Bbc/qlkukjtDgMOORM
vA+YvBUrfJ2fMJG7cWVOhXUqw2+lPccnbskxQ2cPBQJvEJDTZxtK0JvkHGeHh8Wx
rgp6+y9RXr4YAYVjlwHoahQOy98oKy+v3q2ej8x+8b1D2ImQJsO/E7ezppSzD+vk
+1SeLrRkZYsdjfBpe0BOHlQ+sn/Li5WnGpXEpbK0cvuaaWTKJso/zU4wZuQJBdLV
GjCRh5NbL5datFy3qtogLb90CN5xbOR/1P5HzwJyZ3bmFLmkIyyw33tX92wV4GCJ
eGYUY6Z8P9jG11I7NnHzyJpY4z0uXlJLSUNGqHhCu55K4WDAXZy2Mzl2SlIX/OiT
DB2V41zZNwddoFy8BqxqaTSotT9yQnndROaeMwPhyH3yv3BTK2fGM25N/BjUxTNd
lUhutxjrhXRLDMwuIuPby7jddMGVuUBtVGUOX7UjQ1FKW6OGoNl4aKnnEFtgldpf
/jzwZUamkEk7gcWU/HK4QqtlLCWMDNKR+ahhRqhadGVtkWlscMdAYCJjc/0VI5U5
8RrPxYIOKrnyHFZ+MTrc0Ck+79+DOEXz0FYNwM8U8q0DfXau2y/3Psq7nDhg+Cv2
RniStvzM3cEpeoRN/zozVQ5YQJd6OzSqysZNawyHnAAlgaEdAYIoBYGWyZB1YZ+F
ZWBv6KrEYT1wV7hmWoZSeHEuoV4NyjcyIOU9sYIq0Z3KkqJZXkb5Y5n+xtyw8k9d
6Mervx74RQsLkemI6DNYBQYGicKF0XQtpLtvdqVgqlH4z1UYXz+boiVJgoMGNJb9
IcTA8X5I0zX1ejNRPuHaxd7Ir+8nSMYv80l3hppfNJXg8BOAbTmK6ZkI8l+vPsX9
pUnqsin6Y2LxRKQd9IXGyYXTAA6jbxMiYaCX7Lrvi96gcTVzlwGhRVrdQVpPzj3D
a3Cdp+1fNeP62QPXGzlwz6DoEgnTVNM47P8wv7/OVt+L2FKBIZMjrHI7wtZcJSLK
FRHj59UYAX1g05FGw76M+I4RFG1JseQLaAQYK0KEaDTWqTcQ+Foq+RJuOnxlF9pZ
38F5rySgSVkH3X6CGCL9pOBC/pB3w9zx9dSwenvlFit4IHuOs7+GQHXyZs/xtr2a
Dub5/VCVSXMGcXO5u7Bqsoznp3BrF26Bnq1qNmbvFmhs2qb5Lon6UsCqB7GYJ2EA
Nb3lAZFRIkrTINtLwA51u7nRqHcqcgsvS8SZifKkUXj56vrcSu9S3VWUujYRslYg
5ZOCrTCIlyMW/VsjGv1QMiTGaebfwPRhaaR4NmdJfONNZi05ViZ+jg9HDiklBmLC
b/MTf9ZtbVXAMZstfVcaHGmBk8nhCgxPrhe2dY38/aMopqSBaPcyV6L8oFjPGL48
e8ul+YPk+HTKt7YaRByb59m+BTzmN0/IPZNTeSGZ0SsJQd+KtXOfJ4Oq43pqdeDd
m+Ykt2K3rmyehUDXA6dtu5RIbKBIVIa3yu3dZR0+cMmrrxThUbxUKGLwf+raYNlg
hBM0jZK1pB2NzgGOMsJzWTUtDivvv0WiXFWKpb38jeDq0l7REq5DGbj5tBsDOAFz
Ymr/vQ9QS8s/9Oap5Tl86kO91B4/rnyBhJycBt8+z5iQhKKvEFGJ9jBTwN/PQ9m7
H6/Uc87eWBTV0yWbKsnpwXAXPPs/nb+U0ioKHH66tNE7zYTSZVW+BUUiB2yL08eG
U5UkJ49ggm95VDc53QdCnOi6Cw6276SxOBr13GPPJMDjcCIN4rC7huNgSVcqOMCw
ItcL78GB2oFYpXmgFpNqf4sEAXuTgso4+vBvGs2RFOqxvp3d75VFiw4DiSmKP9n1
NkTMn82gbFWS8xoaAb/Gj4682zg5DSwevgRJa6UIl++/7lW6v/Z/8Ywf7x9VBaLd
n8OaeTmUh/N+NtZXl+6jRCDP03YRwx13FwZwDeBV8A0Gbat5KpmVv1HDBFq/bP/W
FinwjqnzkxuJyVGISDD5v3sTZNJbAnKskfYTuXficCVP0iYiCcD6Pdwv/mRVxzKn
00NFmy5b6CETHZt+5HZ4VxgDr7a8VFoFFjnBfpsd5h8pq/Z/pB1NajebN9lF7iVc
Ui+vRGvl0xc3kBLb3hB1A/PWhZG+ClXMbpnjuOCCjOQpCkD5Jgh9FSqzgi+glt+v
MHSRKl7Y9eLnlDex/f1mkAc79TWuowV2u89upoBlyotCuhcoP5wF1UiJRYSo7gsB
Kq/nJLwTQlenUMb/R/wwvcu6J02hcl/mnMWHZuOEI22+QWmVUfvhfpMjUnusKKvq
bt3ynXZLh2r2JTVbqVk4ucZ3WQoNsPbdayh3ehQsCYtHx5i4V8yNaZN5LWEnRqBZ
rpnVR3vH4knW3ncFUbLILPNuTVjwjOUOY6qTdRbt9YDlTcLmaKM0+PlRCEUhFoDL
OH8fZ/TNxI09ZhxaI6411PrK4jrM6I+CDsRKfZXFN/D8aSecBM0oDGwpbEM1GSDm
FWL5fhpML+f4ytpqqeqrfr4OPqLX0NZjNrYDRmAxjqgemHtrrAjG5kiQTkRAURqQ
GYw8BWrzI987gVOqLHPOoZzxTAP7NIaP6enI85PAepV5nYcnUYLpRYIrcwsPtm4m
msAzmXT2E5oDLfsfndYE8WxS2WDrg8duYSbrTaILyoVt44HGnvwWmLBoGOLlRJNM
jOtyc5jbt6tt/+I9I07hA8xdiKIztiIiYjzRj1sfUr8vRHbHvvwEVXLNgDykoTRD
2Q/faNHPzUjPy261WcIiJBh8tWRJ/fdYy3GY4FaU2KkpJ0LeFmITqyh03sZectfs
ixH4Xs0UZCTcUEo8AfEnKyB/5+DLSe4Q0vpKOAZJWRH50jWSdFokZBwayjsvz6vG
fAZMfArs27/Pave/poagDi1UO1rz2pA5embbGjD9k+ijCE7+33OS3MP0feKj6TGj
ED/Wkof+1E8PwWKfbcIKiNFsVUsxiT1dPiX44wc+T1HVViishw7q/v/dBO/QzqrE
TmUgy21Xp1eVYWAuLrNxNzVqzeRoPMuvx7kyTvAEPFyw4TrklpTjqSEX8GgyEfp+
n6gNesHG+ZwQWlVwATpKAUaxbnp8QRmLMkb7KSnmzzfbPllOBH0E16HX9MmJTLGm
sD8AUmxIT3Bdd5cIqkKRjGNLrG/WtkuOqdXPIWYR/Tb56zGpPRPqql31JsVIwKWt
CZ50HJQR3xMnxb1Mk5ZnzMnuTHZaQhrC/q5fWQI3zPkqytFaDd11SY6sXkTKXGgj
U8argucndVwpdJOfGCvQEE7v4cTwTBHPY1KsAZZtO6AxQL2EBL5UbDXYysKZSp49
xd/UxxHQa9IdI7Mcvs5tag+VEH2UVdTbv7lu3sH/X3O1V32jlSfAuSwWtn31dg2o
/WNr0aUGnZRZT0RBQJtMe/CooF5P1Qff55E7LMB+fSj6HJ+bhTWyzXRXBI/YBJrs
JToRNJRu7YnHppd3QYGHFrB2+BZyTfTlLPIv4PxajskjNB4olZa6NyaMuhLs5/Mi
jAc7l5I3oXOkIRV5TFEynusTzRLpvMx0RXSG0axJ3gpiWVe4f/OXtBsCt6Kaj1Yq
r/+NsYg7HUJhf6pDaBjawcP6Tu1WY9JyAgLM7ZRpSg4AUaF3OlNTB3Gy6QSbOCGj
bPuPbbQlM9+S7Ej1FsU10CcUS3xU0cE3XKB/t1Rp5WAP0e6IF5ZymxxE4vJo1C6G
LVGXFBnqvQXfHlEBn73nVwY3czK2k0xpClQMyvxOMnuaKZqiQFL34BFm2fO13EqK
fcjTFqjSPGBQb/GX6RaDtey4nfY038QmO+aiRBwKltELbd3w62cQeR8DL/0Yl6X5
Qu4MdY773BkgIsTpBeQZ6TcagwS9AuN10EFnX3LsuqKPS0a7zrHwkmTz9qRwqKJ1
ShsKTcLwPq3eD/3lnmt7slkwOLJ9kCVklzq91+3UX/IgeDqgCjSldOK7tGjVn5HF
zC8IyGBF1cfe/GNh+9WC4K+BoYZKgknTAKd8wic/hWSgysE4s1+PvE+295ACeBei
Y2URH9voPuXw8byy9Awz+nZtMoqXt4zMYT+39ek48cG+9OP+Q2On4hNx+neLFIA4
d+hlyO2qovnL5btPOnNvsKWvgbIojefCdCGo2ZZRW5a6SPunj9ZEgNrhkWGrw8i0
YMmaf3v+a6DO8YWx3DPIlMC8LH8zHgWuWySu7+XvrYSVMmjZPNp+mbMMLE3L0UdC
doILEA9psARzSv7MEGqO085wcB0XEavphs2k5se4BA6BpkxSmL3CqkM1DbwkW2gH
KDlgvpZjc3EYzc86a10sawIJwNgVgXB+NGRmZzcBLEK2XysCbyti2CKDLRyAXqKZ
sXDKHb8u7cUNjnkGgdC+wt7ZkNNLAGJddJAZ5jfyO1FrQVSdiWhZL8nRyOk5HZye
IqpZiZcy2ectxUBZ5fJGW1LmkL3SqyVS3xWG3t9uYc2eFN+cL3LDgRIH19IHw4wO
1opfGjxJUVk/hqk6lzKjbcUE9asfAvfOLZyvgcWSvllRyLVIVXFeTJgcIyd2UP0B
bj1C/M5EmBUBwC9jK5EllxKJ9AQLg69DWw2APrM95N6lNziHn+7dLu1vIoq5NSnK
dzgvvE5r2kPaP6mF+BWJUFwXp22zEGXshr45eDXk4weFUQyZHaya9cIm2+Tg0OS6
157QF6jXaddiCzZqvZ3JNLs3FoTHj4zABjrKZmsf2nNbRfsEOx/qH9e4+5E7NYVx
M+WPOFhTvCSe9t73fW+XRhHBX8EknWno7ALLkK+qGfesIkZjkqktV7kTN8DIrjQ3
fsHDsUb6ghtiyeLwmB1RUm+grD/5qapKtsz3LHbpt7vx92B5ypG58R/zC3c+Q8cK
6uiXJMAAD3aUK9VSWJ+qwE6q5MEv+pgY1IhQ7GcnS2vF/KFOaVzXZEOo77w5x5/3
U5vxzecTN5Cwr5OOWSHzCzimX9sxryR6HzrCA1IBR/jODptt/DSfb/O/hT2J+yoT
DmEOwH3125XPLKLNemACZk8qruasmxhigP+VS8lRNp63nYNrdDXz/xjAezCyS6bD
uCszm3/eyjqB3Z2tmatY0GMjgeDDCneyxTsSrs5FLeiqP6ZKl78/jNkaFDPAJRLo
bKJnbwRGnkNruZSwjHy02GGGv0BjxdeAzMQzTNsgXt88dyRQ8ap0fIYXTpktYiYw
AZTbytWyDC92tWEe5goGoFSBzidECGQf2OkSpr+quKET+uKtc7/n+8GZ32nbAR9B
X8JhUjR7REbUKYrzcjIKjfAqpBJogqyGrNyake+e4wz1ulWcT2t/K1Gon7nP/+sE
t72QZy/wkP/e934jAgYPZaFRi54HkDX9iLjX9mznHENPtVS2kkM48rqqw05MyCiD
5U3YJax8033c5IzN/Z3VjkaOyRoQ16JNTkFA4e5T/HiC5mdsQiMW+Y+s7JYHge2J
dMDMggnk2tKVd8HRKIcNlS9HHYTIRTspoVcnIpp9/EvETk054MbIoqQlG877pGYr
Fxgutur8r4K3Ksy9sVaO4RWc8UbBbCOsSuiO8bXY/dieADMKWnR3L63ocPXIZ397
eysLJNF0evzuWG1NxyBLLZ8uvPXn9PwkooVBsvDWHsvq9e/5hdarsp6n8pggG/E9
A/7gGTUB8KpeaVVeqVkqa+N0gLXDn3WAtIyn7uEzwag5XRbDr3ulz4ALilDYlaFp
X6hWS++qLKpXa1nGjpB5Uwlb/gyF1VE1N4xsyqzelOKq4miknDz92JqeG3pQCNL/
LKwiBL6TvI/RsDhBuF7Ai2nkortASkL0rQHXAJr0IHADEdxiJiw7OfRqpXdUXS/0
hMTIMkFnINr+25SIDbAZs+i1ah/9FFgvXW74XXXSS6mEWGcQexUuoHbsOF65j6il
owv1pCHwQyMDQSoYBKxsrHlF/8MjU5cCKJ+Pxx30ga0PoQ0rLhmtBLE2dz9Fmh/Q
T6OKb/X2c0rkPa3hfGn44GKgowtLHdbgQt6It6Obu1I=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UYUjFKvvDAzEic0tJJ/VgtbiUPxIUuAf8bVogg7kNzd6iJO3SsrbBQYAvxHfTo8T
G7jtpUzoZCFK6m8g7aKZUqG+PxmxX7xyrqQC9ZGm7zlscRJtw2ajgXmuiXvv2rsj
iyvb9uYdaFv00GHEiBOKhDO00lC2Tw4qXQW0zLqAgNmULCGfhor48ivGBjjpUcvP
LxBq+/AnMSuHtxgKTpedLtoj/zkQaZXs/35fbhEYYyjf+53P8EOhSpNO5YxX+lUV
qH94TCIhe6MOvXOTCdLRbFMk+MzWnoEXBqFl6HLbdbPyKZhSh9ddxyjvd8A/aSjM
CAF2arE2mV1IawsEQ8vfwA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7632 )
`pragma protect data_block
zvReRDJvzuyGxy5FJHYwHXAv7Vvs+1Q8gcyeUAtBgawzoUBmf4q9/8Rrl2qEjqnB
EUNHRb4OExWHEKfzZoySIGLIyCqBLRgV/n2YWqRygokekvvUTVGT4VLVJAk+V/JA
+tf9fs9IWwnWGmgqboVrOJjj2+gg4IczEUZhuF8+yKM+xk9IeWAuWlYmP5bNIX4/
TliIlC6fQ2drjaQSaYEYQtqnKqH63Dkh703CPsJAdf4unD8oxeIKUdcmaqd+sOiE
CWmfVKydRLBwXfvfj2alxrUlUmxO//wogajko8fBnPiNS0X+g0esjdvE0K4R5LnK
9P79SEyGcnAmlovDpjEscXJeKRLVprL5sWxLJW68nfN+VgOmq0EjHKzhVRrJT9U5
Ntr/LkEjgaevpiMCC6KvB8+Sy71+8a7zcElcKzy4LLsquEHO2bYYtD7i4S8UDToS
2iVnO2djBfQX5epokpJK21SU5aE+8t51xOaaUDECxEUaDA9I5YcoMmXwOB5RJwPn
D3vAJ67PyRUQHHpRAW2guDOvviYZ1B93zY/DITXsqR71VKT7depzCPgF3D7DQeJi
FhzHTy6y28H8i+8Cxrkj03qGopSkJpykEWn7ZH70Jy8BtN0mRp7BkZE0vUYVrwUw
efFZ37ryp60bCkFgl5bzF5rkcvf5aFbLUF+FOVMVRjkLqSmp7tyO8rhxdsbe2G17
PSXwyf8lsOf7DVrdE5QI6BieZnjaOXln8AOX0ADkrY28cfMTTYUbdcl/w8HnjZsi
km3F3GMsEpx666oeGtAHa7mJnGIRWxpPBBwBdYfs6aqBooF9n4L/RoXWbtuWT2fR
8JDOe2FQSs0SkamycYhK8yVH/N8K+l29M0AWaMd1i6xQF+Dtnyk6DBK/jD9lEEEF
5UmLPm0hI4Ru2MkPo/+PsbVHVxH5IunKkjEf+lkPOLVHimx51fOyBv+iO+5T30JO
jlXEw/dwnGgDkwplyi/BRFHjJjIQrX3qwhFGTuuHfVXDgnEG8l0/Jv4ttmEoHIH8
xlQYGP4mgoPvxxO4QCbvGI5ZuUuXxDoUkzMJAZEzLzvozkIwiRG2OGtqGiphxzy5
tmRNk6KtfIelplL4zrBc17OESjx7TWcUcF+BCUzxpY0hOpNAQ/VpSnsfbvika1hl
QkoOIGeHi8nbZRPOvUa7RuN8y/Wb65NOC4Sg41gs3LfNXzbyPv3SoWBWhP1fOcz6
XAabI9Fp5V2To4KhnrFJYxRkvIk1rhgbOCHbcNfuwrDpSCUScsYYKJBSDb1m9b+7
u8nrTFg0txXUj5/yqmh0M6o4EDYfhG+MHzR/sAwYz3YIs5M0JUk1wo1sCE0fYqP9
DcGRFNKjp0wkbOvMJRlpETyqNdQru4ILWFxoIX2tKdKalIrWmtIkMXQ0fza9PNSK
8weu7+iL7LJOeLWDzDH45lfzsNudm8ZUW6C3HF3OZji13iyphNpsRzzVYXohy2Mx
571la8xg3a88bxGwy/kDHdouGFrc05TlS+88WYqd7/B9BKaW+3oXt9z9Tp5DCtjk
VOUR8E3h7anwJXEH1BcRP0cUFHXbAxx+FFmrQyD8eUhrhUv7n3pakPc20/IG48sC
NQSc6/kLXA56XSwvJdZa7yZ1COVy7XsZrNxkCXDdsa1B5tkbeDhWf/2orHGW6wDn
BXRyuoJctGDSZB0CSu0fKMiYAFdmciu5uZ7AyrcHhvftzvcylfE+QF15hbcZKTsn
srbjLofEBj0QPQmkzziQBdfxYFD65GlkJMhAmrNdj7lg2RCh3XZo1DXZhzD9wV1p
XkDcez3FfWpXTWSp+AAumqzH7dMCTcuHIbvZHaOd/Gh5vslA53AymI82mLoztlVG
NcuQLA2rib1v50pZfgR9CbmP2Lk6/XDy1TRy08i4SZpSV3sIHDuTO0ik5JchauJw
nODSVG8maLHMXVuMysIshB2XqQL49CDMpY2VfDTuisYlu8UBEbpP0zBXw+v/HGWY
2Hf/wA+SvXX43tKOa3Vb1qoIiRzTIkTcEIpWlSdaHCM5FvxU/5VK74I6Q4vy+mOu
9RKs97KSDV0qZNi9p8vhaCtlEkDNO6848QVngMwYk0AJHXw+v3ku0u4tQE7YWMRX
Gns9NGYmzDdnKsWj6TtKw+Cl2PTL3i5huhOULXg/SUF/eKgqjo0/67N2DnwKa5Kh
LxbnsJll8uAwS661rAforLIG7PG3wMsL3vTDaYSsk/dn75UIxz23j9+GNiq3cmo6
74TPkvAh7N6A18zCbOwxWyFh9nV/DFgdPiEKHT9tE6GJRoLWzaT4Fmor6Q23ziD1
m7I/utpEHbCSzMbHfXO4Wbu6pKcXLjkd4J5z1b0TFsrco4fq3hwqU+lzlKYn/ODH
N0Xe97kP4Q7clp3lVgiCV3EKXCy4+r86dF1HiknCkLX5tT/38EKiiWK9pAgewmLq
XVnOGm8dTgORdAagvcZ2cblqL3HJefOqj2+M9sFgmeCDYdyZTMVNYvL11g1sHKDu
n0y+N1oHLGFCsBNqSlSGEGLWP0i0oJI0KAb/+9U/Zd0VpTTKy/Cd2kJcNorxGyre
tL80oR1zxK9aBdfBi/RDY4axI+DMc1iv/bp1jAgYazwFirtZGXe/StcgdydupMME
IwMmJErrn4nQLuiJdoCyyU11e87zsHrojtZN/gdieSWIruPN3QZ98NDotn217UAs
ImC+bbFHE5FOoVidLEPsmcqxrXxXNFmvicMsR0Z1riiXr5OZZVLyJvMmt/qgSlLX
FIpEVaOKee9MTajvpvBsb40Om6Q47SxX0hA1grfytfYHiYhchAf3JQOWltdqrY8b
i2sD+nd0h/4Zt0hDrNElT0M2/OwLRVr/kmZgJkZsJGqR3iULXWqW7o8ZcemnFtJm
E5sZ8PVQBmkLfxBl3tdrLQdsg69t3ID8ytBPpWkZMPIGOJ+6I0ikyyrCfWDNYXbi
hgt/PPvqyY+g1MyPJ8lq1/hfgzc4C4qTJKCc7kLxctBi0jqIEl6uxd2i29lKhGju
UpjAnGjpBgPKvqZrdyXZmzfoAJQTKXnyIm69rOJoWY6hqqNOy+1mEbkGelUaPCej
fV2aBqIbT9k/fTyDJexdC0iihXlSNKwQqNc1gAwltqtXwMuNWlNoxNaMVtDqHaIe
oFCez9ITIah/cqUB0VTDLsnkpEileEjspZ5VdrkHFujNdrD92GHMLYy48JQ+pu5C
o1jpJ0NDhfsyIC8Vjew03jNy81iP27EnEZQpCDEGHnvTwndkwHJBBn8ZzfXVpsrN
kYr+7X6TyUQX4CcSvkoZLjvqtFCOkyreLZ6K+ibJ1s7oKGPK/98iR+boXb+6SwG/
NBtyo2zkB8wYc1E4s3cOuvOaycWekqyCFkCQqXIuKd1vJJh9OO/zzgq2VksSP/Y7
JVXlkxTOdd6V8Pl64nMRo69Sc/IEvvmSBRhGvTdBVH4fdZqhRms9CcXB8HrPV8uR
g/Gq6ElrvEESfIJZgGzJvCxxv6spR2OkYF1xBPfnWz85641KU8qWnH5Ux6yuccLA
yUClou9LPSyT8dInPougX1Sxs3jzXe6QLGmMoA047LHI3YoXKGJMWUwfuATVpxBc
uu0dp8jI7CkTk89+vQ3FKtc6plMGVtCy8FJL5StOCDyLgPllBEawW1jUb58GAjG3
cgNhK3a/OdPpry6aqRr6CXIe6xfN+gRFc2TlPONh3DbSDvHD+TOWGsvLcH1YuH5o
iubEV0L05IvKjFi6Om9/sG+qRDltCGwk0I3c3g1J2Tl/qpkhcdnjObpKPu9ZXyPN
fd9NR/0ybUUjjZgB33w/gRhdcEPVRSJWGynjONFCR3fknF28al+WRMRLm4uJNyfp
ENY6Z58wUB6lXt0cz3/bF2yFka5I7b52nG3EirsvA7pqp8fMB3PgsKz53GNqXhcq
QopJ0EsL7opOKQAeFOdSmVg2vreMJ4XKOBisF0pgs8ID+XPnwLoEHixwCMcTQntj
zj0Q9IwO02j99DUqCOGUkfrhmhY8QdAZAiaQPEVEa7DcPckUE89wsGhxj2Cvvavh
5Kg79Jt7XLGAkEbE6b5bMzRGT5gOFb/dbrsIXxh0BYu49pT1DTXyI0xraY3k8HwX
LtdoAsWDHONNe6z2u6Gk7b4HlsPOAV2+12p1NPgnzGMAkOH9V+h0B0VngmBE6ILj
tLMk+8pGaED6hKPouQQAIS6rjfjOROysgx/taHbQDGlbmkHD579Epy2btwKESLni
8vW845FpZgaVRkf02SFN0tbW4IwwktIyzrpTxLSeiYUyEttQ3/YhJmCHNuakb6t7
JnJS1DHXCTouWxomMf2a57J6lKuPU5zMvD4xmCfazxyVeUBnc4ExnjuD3hg1qQEW
fCvlhMPmCOFn8MFw5I8IEDUEHcG60wA8ZoeEON9yS9y24gRdbcq3i+1bcbaWn8gC
XCeMLU9A9MIvwOo7ObDPu8dIgb5kXV5yNidGis8wEvQbboSvVBLjZjulR8i18zmU
Pt7Bo6OgUXam1hnhHLnjCCI1wjwVRlntC2Ku6nk1XT3TAus4tnOFUZL2t4qCA9iz
4kg/Inne7pyVQksoEsemXudCLCINGXT7/iZgl97Lxb9X8OJ7XxkmFjvfhyqozVpQ
9NriNUYwC3jjhELckowVOrPfb+7Nz7JgbCsYd0OJGJXI48Lvs9xvEMaI1MaZyfvP
LzLjCNQodmX3E7z+uBiWz9fChT+m9RXCFCi8rWFcij6KnfrQDG8jYSO9W0AUqMZM
Td+JvXYsCcTl9DYYPcVuO8mLwHPC3GvqT8RfAeMu9MKnHD7ermarU7wHdpLMTrng
DtE0EwrGeVoHIr8KsfYzDlk1YU+z17XIvaL2KjTrR3Q1KoIiuK21vt4SNewgJUHL
E5vmFAId8UV7ID2FH7l89oksaP7qvPE5EBJfSs3TtPMq3l7i2UFGQrAyZkVdeX2h
vLMHFZYUGwBKWXvcOIhVx/PF65sbQREnsEMu9CKhtQ582X2F30WyWlU1ufdkxz4q
OmdthsdhJ6Yds0fzOz3UqQMlyAwHahGIsR0boLxN9nki2a5dur2BlSsX61/SE/jz
wuJMZNA/DtG+NByw7JXv768kSiv7UHh/2m6FJFLKI31C6rttrlUGdY+r46GTbQN6
ZHw6ooU0+HzcajjT0h9vYmlp3PbdNWaq1k4VZmUMfiyXaSf7v0pgjxAstw0CpkXM
dDDB1AqPWn/m244msn+LZRE0m5syK+s7ha4jqzYV5GH41YJdKVR3C9CNAoBReL8z
qVsMZhokUKs1AINWf8RPpXna0a11OE+2PoYnRuMARi4KoipRziFVYNO5LkWv3Fip
mYWWbjGPP0PTZ4/6l6/9u5ZQmwjxZr3U+yfC6u3jnOwN5ocQ+AKtg7HBgZGjSmrS
9HfMMqhkb1dZ20eAtpwzE8gQZkv2xNJTTUKC4Zci+o27lcqGGhWBRnFhsOD15vve
ykCBRcTckbsn4IBOZs/+3OIDPGtF4Q6zd0gS9WS4CZn8vgZpWNBONCYQIFiS/Em8
LUYzWCV06d6hACipwiK3icea5wjCCMMQfnJBZeV44dNS5xrCINBd3lgkgUa6veS3
VLbQiuHLoghWMugWDQiIcBzXgWp8Jnn8i/tS47LOhl8WytHKKZEjR6hPt+mdUm+a
q6dCGp26qgtKDMgFHhz7n3ZpCif+nUvuSaLJn2LFf1QX190SQYC3cLZe+l2SDhhh
W1hSbLWnprcy1jtckweKzKZN8CMZrBqkhfZZPGUBMdjalMisfaliIYNR3JSVsLxv
zHUbLsLIz/0eTSXlwwX7GmeYjEUiQBUOY9CYDIZqAuoCDRIZVJviHYYZGb8GW/pN
oDtmoAJMzXpO71BNcCl+prRyrCTYVDhAIeJVxQCWGEsftRTTjPrSh0ECnapNS11B
NtuImqpd0QaRJ+4f2TvFegcV22kCrSfL/Ket4fthgB9M7Fr2Wr0pfBK8VMOHLbSi
y63itbzvjCseI/hVje/JvhHp/hI7XC1xKnYiUlxxS9gTQguPvYHJ3uB/1lTNHmBv
htrfw2l/8ifpI7+K91N/YgfZEbIuSAkn0PCU9enZbcJlRxJ07evIZtr9uKuYIfbC
FHTMDz4AO08jAxNUsYm6L3W0lr9nzXpN2RjPw1kxgca+id7qa4gQO87O3/IGu+BP
lBIcd3rOiI4zutfrJDN8vatcmFCg9KyfxI/eIEN86WWbJMaXzwo66INQzatV6uYH
nHImNjnfv+8hSB9Ikc7GdVRXCSVPvb8RwIEFNfPjneIWh8ZJQLIEpRXCsLnF6pZd
rPDP1fVY0a3XSvsSoa9bXu3uCuvWVALQl4ifrCmPYDV6EZc4LfwXW4fdBJTipEmQ
UVMlkFX0KCR0dfvMJBb8bewpETUGDP6NDo3IOWLHkRz+uOHxd4u5p28BOoQ5LHP/
Ndqxc55G0RNVDBj5IMmAuWuTtq+Jen15JUyIdbDqSKm1CDSAgMFsfWemDR8U8G2Z
ZV96fwX6xOh5TivPbg4N7aFczMk+K7kh9QeJhnmqEPq7oxe2yPFs2NlG02Tcb1pg
4WTLbAnybfR6o19A6wLbkeCezye8tbOSbrAKZK3jEoQ9zGQiAbGiPuX6mgx1Fbd9
kxlmy4PXsYBIN9hqTTqgbLaxKaBV0asGicL/Rq+ClUS9EgXwNgQD/C64OWEDXYKL
Ahrp/0+/EYXUz6gpDSOCQggSXwTNqf25xBZHMzAbAoGcgcMNKWlKupoaPTAIwhGe
IRLahrX3Z6qWMXHntVTC9qgkL1Ky/yXYi/6WvXni4mIw8sey8b0+LMkkKARGumFC
t78QJzsIaz+/xEJI1S6os9h6juocX07NpMixSq84mKcopUQcxuFeso/LFX+97g1V
aTckCtxdXgmTRjvicWLXep6vUFOnPILSTJa9HCWMNnkdsKvdynoEwpv0GZ5cYgGQ
OV0Lk1zr3Xbdcj/DNPtHA/bbaHmis0iKQCCrCN7ugqyWfsUjJn7FonFfLpp1XSiL
Q4oTjhiBgHw1q52tom4ZJnIs1764HdiRuoVyzQ9M0ZX7Ku1s+AZBa3lm46ts4M38
yfho3ZCey0TigEFZs+eOFi6vqDTAlwA9uCXLLeQQ5pYn40IPUM7wtqjYRSbSl9D9
n4+tbHH1aOzPFeisxF0hgIlk006k0tIfKpogQPH4ZHR5jFYWbB3UPMw+HJ7vVqi1
Z4xr8UDl8kKMwNcviOWSIysHaohEssicHE5WHSoHNLfrcZVmgCBYizerOffcSoRg
LyegRDIJz1C/W8Z5zen+yStAxymlS9da1/Oih9mwk9uqvadr0f+h1ArXiqAfIQhD
Cr5wgvQiZbQxLH1qo68iLEu0dM2HgUplT4QcIVv2jMUtO6pzBCJO8dxbiZB48bQX
igVY5S3dreJXCqUoBNdL1YU2GqmcJCJjZ+5SeLKd1BjWTBbw4JczLrC7EKdMs/qO
jlkpazB/Chunal3L477sEuCTw8tMhiMJ+fzdsnmLETgoDztV6/4QLLKostiX51Su
ymWcwvjk74mfYM2OoK2Be9TZRTSNsQ8xTmK8RZQ/CmZNlvAFYWu7wqVFNY8XKnjH
iWUhwjxKy3dnOy/uJGrWMNJwxuedJVRGpWCZEwEiXvIw6YGAymdWlUEmGcWYjxxf
1KNwEHBaok9xzq7ub1g6A0NwL2yXhC7LxSp4Nuppnc1Kdj19N9ejqoHVyyoKi5j/
eH3sN9GXE6LPm+mNGlBjyc7ES51aEDheT7hqLW2wV7uMI2HhgKU0mR7ZY1O3lUg0
xkP4I/XscLYIH6D1+mDBblYZUBFLQVKQsblbbMUyNt0ReMM6G32O+7jTMI4Af9tu
yWZE6jUhgHdIYzXa84OT6kc5/qhJ6n0QwlVpxF05p9ht9nYFSeOWwl1fsve6QEzG
/WB+kTE9dRZAqOaFsJ7eCJdlOpUpwfJoP3ghChAfSBNfE158uVpu6Oqo92cHofCy
olMNWH670Tii6LoDeC7licEa1ebhi0W0zhisOaqt2A0j7Y8jDGrwsGQ3G1iDnyoS
Wp7EMAnO7CLtcekXraoRDFfiW8b+pHIK2dGf6gL3FQFX0+lRzMvPBlc9zUdR8UI4
PyEG4pQ2I2+FzN1PZaGhnEzs0JycsQkT52NnEYpteZ8H6fw9uX8NmGk7rbJ6xG53
pYfsvKhNy89qNNitMDgL2i8k7SlGLtRwhPEl0hQOhAQQEkgBLkHa/snu/1yw0v8t
CvHtDxyeaXN51+Q7rIXEMbN6yzgDRBymbyhVY84ItdD4OyI+CZwcGVV/MoqazY67
Mw4Ns6Po8Id4zGkeRtOJr9CIZJpPvkxWS8f76ZIeQw63b1ZGW+n2xiSIM0Ae1KMb
cTmWxvzIeu0+m3pH2I0OBqjfgO28uITl/cgcpVMiFNc41ULTtxrC1yv1YmlvtOHH
70cIH1VkID/WKleUPS96n2XW9P4EGlBhL58vy5/TLHOwzN0/3AiJVoikX4B/0oF/
yfHdo8xYTsTZI2q+blyCdu4iAK248fAleumDlBVUNw20uTo1JNbGp6ohfXx1rhXn
sSV+1C9etihF+sR/Xe2hf9zKrz+Bp79nOxoTssBmWZASgLjj2OGBoJJW/mp22NvK
kY4sCpK3WqwPmRTb8zDQfsr8Gt+7S4niUOuSJ6hOJjbgDMhpCBwYO6pw7gVOPY1W
f4J7Y/gR5X3/EpAExuCHVc++S7RckQQHuJPhTBL7lLwwdikNVuOOCt4qOEvih5ay
xv/OR0S2yK6tRMj0XJp7J1wVRaPGnONpvFxGjnna5xRFTPXJ2J/IQFJ3oREpERZG
pRTGGwjDoehNarzc/QlE6ipUVY5MKwz2/TRruCOmHM2yr2CUiNiT7a18mvwNONv3
MGxCYIEPpQz/W3DnJ4cPpuoc5YBqRfNP8swUS+0g1Y6RtD3PVl7cUy2xFG/BWtbE
EBZj3RFx0iOkskZBjkHblW30nbQSxM6RlcjYtQj+OLcyAgdqL2liFyPtUTjHDlON
NK5fGjKUm5pN7UnS9N+K84RqAhOSDDjbLBORoR8ZXbS75CGxueIzd+advcazFk/g
aHLgOydeExLUFUmPjaA/S4CISYd9K0rlCUTniZnc4fP8IN0qgtwme0ix9BsA/TfQ
qQri814xG58DihRcSN1/ssnkinplD6BpdUYo8defZ8IqRrIEbFsr0SFMhkJkyD0B
25+lkyIovgjc+3RpkvoPmmDD+Ei2pzjI4Y8PvQ9hakSL6oeKFiu2DewvIrbtyArf
Gexkka1Ymoxt7SwWrHhAH9LS0Tg+WDiVUHZYvBiTgJEcoKelim5R3xifvD/uxhJR
455YrTuNgy8HCiTkjsj4e1uN0RDOV6o4WrPmHmwIjzKb5uWlng8IQfWHNC2NSf24
jC9kIkmFW2zVG73r99fZs6qs/Q9BSkQFlUtWbo1N7LcywZMfelSPUEJI/PC2so1Z
5CA30OzRKiidvOQnZAIvRgWJVA70IMxkV7ZTymaFQpqagCh10Xt8lZ9OovOSrsZ2
ua//p4sw7y7JJ/A22vmN8QPQrPRz6zoK2k2fqh0xjspt1SDcE9V/aOVAqzRX1WnH
KwqU410A+vEElkPSBvBtCuh89I3Tdh/zkYWnIaKh4dtLGmQKTnWs/gv6aeNk59uh
aqf4VXQMCg8xMi/S8sUuLlJaLmUcVWQAXbgW0481wMJA+/BOUTa4NwXkqSpT3NBH
UfU4y3PTPddcDkKYZdjUXVdZ4BXSgCIMzTpo20z/ebbTqXaJpATMEqqSReEqd5u5
KM7xpyT+2w5mMZPmdT+nQoVhOmiDFKKGuFFSq+JRIITBPblNCllq3K0E7/Vo3qjj
uqBKCPj35au1QUTWDSFZFv69EGJQniP8FKNOkeZVWEjoZXeOo6OR8+RdN3n4dMWu
isVNAm0iD5uBhkbEIpJiyNNT5H74S+lrVFP7Mnlzg+jDTuqiPBgpgVWInYuYtlIM
aYCa+mvLpxLey4Tc/D4lal3fVK5X17++zAnI9L3pBAwTB9uM6HvG6xMB5ZONEs5+
YwFvy/XJR+W+heVkkqxeL8cUYmx5/TtlM+om/JXvMBm+6SSbGbJRuHb6d0dm+mdO
b/UmDnVQmg6+QzY0yvzyDbIasLgyTdPoTe/Uz81shEu0KqUnobU3+F857cW3XzOc
ZwVM/kQZKyA6trOpiloEksWHk0+llunywQ2YouZaCl24wOkJe9GoananalNRNAEo
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
f1jkbdPFF/+potOcG5lQpNS6QY+BLAr1e/6XmsUV2xWq+x1EV9gX0A0c86BwuKw1
XzFywCbMcPb63pNmw9hpdWxBu7M7mjGpbPIqVDe3UDSrbYqvqBVeGsTY+oLGi+y5
GijgyorJUd6JhIHeWIskrOJAs6SGnRw/Fi88uLhCx2AKShykHGyjVyskgE6HP9f0
hiG0FjUryLqfruY59MwVp38mMNi5NmCnHSa7qGOlaczHvGGY3lR2HBJjHDRaWEha
A7prjeUK5N+OsqAVU79SNnGAIlr5awbPysk71VKpriOXdq+3lORhErLdmB9WyqHu
NMhi7bzIfqRF1bpgQ27ILw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4768 )
`pragma protect data_block
RZoPwNRvw4kzXNAR0+6vnoUzoFvbuROOiJLge7DRl1RVHmry6O3Dy5rHyaQxEHUf
HGPv6mp60FDzPjA2zpqVLq8/xebABvEKse04jJMB+evPmw/8aB+/AWDgOTOw8AOy
1B/qla4uT072JcLXsyM05FsFXsk4OfILvRPWO5u9Dgtd12XlZGcxbzl1TzicSHT1
wd9CfwZD1OIPqJbgbPBltepJwgPNClIoOrjyld0BfUaZWMRJTc7/ElKHNl7zp2W2
71wzMQk1f4l8VSmOTmLJpWcm/qWwp90OSxKV+8SgLoP2OWkhayKHtD9AcuRZAxs8
iJ6SAY/xOW35lXxIsPgkmwdMPBlYBMTT5f/4/kYOIraqgfbxrlwfiCQmCt+2zgXd
y8her9IYsMOghclBN6dz/RejW8i99rSovxFb3Ql5Dr5D7Ixcto5/Ab0MfUjKJCw4
XIDalWYiSz64T4XG84G7+xFAoWQLemtOVWpTK1U4T8jWwJ3/G64NReXOTs62yyR6
994zzmmY38p6o95w6tvFAJxVdNT1ZXX0JMqHMiJdsfS7XGG61Fn4n+vhWH1/h4Dl
p/6UIoOWAFPGpPP1owe4Ihmn4XMVO+ETTskL6njy6ia03XXDlThilYMws3NxRk5U
NjT/jLwCkiwvkva+NSXXcqHLb+WuKBW4ZRKgpJV8OLBOm6p9xdu90qMNuV/wPIZQ
HMLpI/Nu022q0tK/74qQqLdYnCKmKynmSNgMXtMe3K68MxuvU53muku6EAdXUTto
KvQA9qF1JvCKKRBWvim5TfwR0EkaHRJ1BtcY10bpRJhMIQ9rglI3JN2n2dzsHGTC
OJC0NUzhvdCPD771DGv4qpuo50OQTu5HJjFDFJdaNW0/DZo0UWIfAEZ13hJkJ/rU
NtKJoVO0MvvQNm1nwZP/jxyjlKPPybZg2MdjIIzamsqyr+cFl50oWUPbZ0uGwpv5
pKOR0BBadp0MysxXhs9WTE9rOFzUYk5Kh/F9/CpfeOr3UA2NVgu9AMZ/r2w9bG0P
5a08CdjerTKSO6N0kslX8WyWaPKpaVTMt91nG0QFCgf3nU02YEkzEYgnrjobHfbh
Y9q9s7g6Uegd6NmmXbqj78T4k8PA4ZTVWvk4e3R2OnT9ipcvwV+uz6JpVOwuphZR
79nEsStw+tYqq35Fwabk0voo0peFlhj2PtAzHMmD3RBgsaNzx7MGK5aESIBAjC9w
UhpnRYpo5Sa+MjiJqiW1vITsa7yyvk/BmqLJBuFYWQDgS1GMi/XvHbkFS/YTOrh1
oDoJiJev3LnOCKcZUeUGOrOwsY1mwu1huD/ZWtzILk4ou1Ova5hBca1CLmpHouuS
uJZ9zm+5/CCowXximWbOUGMp5huyx4xdq+IhwEwVXYj/Tcmc7TwXMudXzCrtcKWJ
dbUdLg1Z5xf6Q0YSFumX8jb3lYGbSFqkC7aYEH5nkVrHiur29A6X69s0SyZ/BxVv
ZSdZOemwHB3+9Jh0Wrz9vRUJyH+0VdowEmyhipW0bLPlI3POAPKgZGluU9X9XG5i
fjEiX47ZMBcSBauyCWLs6hzADIM18esOE0+FRUIqiOdgw7DC/pgapvkhvED0KMUu
lEe02t9rczrq3jgZcz0FJfotbelzFDR1HJUs+Q0FJ/EC2gBJFR8E4aXOP2JrnLy7
1+00g7yaRnOxewc0+RvEqdePLlUkmgNgMoZtwic8bfOqKt8eHFMh4u6UUD8NB5S7
9iFXOikz1SrnQB/KQY7e8mUMD8SZLG1y+aug9A+q7wB5i7kOEXonCL9l7L/uaHhm
GQVmiLDHsK1gAEBD2EK+/ciKX8ZvR5zC4XFfyNaHIQBDA2bx0n4pe1L2aGTQ0Ki1
ray3XxGCV/gY1KpqE+Ox+5iRkvzbtCBmtwyz+e2JVZ8ND8SgYBnr7IyP6sbcLmxV
A/10DlXk3WuVRzTtido/yS6OGJ/31beATm1BbeK/bE3asRKJMNnUb5pBQEYaLv2m
PYRfuF0aUCji61jJnL7Czrb1d32+ql2YX/Rr987iF3N8nEbP4e0Vj0nd4n+lb654
xUssr2IqeXJORIau5JbR4TsGgk1r9lKq4Dp6DiamSejmVGWhXbADEDwo6K1r60zb
8/x0VqWC9mbQix8js7mW7g4SLzX5ldC9tJozWyNgp7Q1NLoU0cH7iFacfuFLB+Fh
E1RYnJIYI7Kj4uVN3Xbp1BN67z9DjYbBVdrinQ3Yj/3/SYPyIYeY0tFfFnPbf2Yi
8n3W5QqHQvPpWWRyLBrsGDcIC0M4Zphthh1ucAdIAPXN9dPnmhGH2+ycwR9ps8J4
oeA4AHrsK+9qCoAOeuIP7bYKNxJSZ0ptLUSb9VfrFLbgrB06gZyGedKfx6v7Mr4D
oRAZPTWs/PFLxM0sOKv/fgafgDX7cE63QIE/uFQt5eyTp9g/ULG9448muW5Yf/pR
932dNPL103VSgK/HpY8uUySzL/uU0GfgdMAGN67QliFz1jE+/2uubtxr2oyabZQW
9AgoLEeTpZjJ6OWqg+n5T4ksTj3RYV+XP7IK8nT4dkrT6I3zgWTOoA1BFfTaG6gP
gLkK/L/rAOGKi7d+GdzT/mMR3F1rv+8vyEfJV/AC8uhWP1HI41DESfP97VQhD4DI
2hDw34K8hxJMeGmVz5pRjfhPPMZyY+s4CdBsWyf7o101QprpOKm4BSExQNwfjJrA
RGp/iohF3ui89mMMS+p/NBn4gl3O9kWwC6xFS0+oJo5yJW6tnoa97YKfjkQaCAw/
3uGv/+TObSX0vVe5HYXxHK5lH9EX36iQuo0ZWXESy0c/ti0DtizQ9Zb+9fe95ca1
YWuyHCCQyFuHjfAbkm4vQfrWxC3PFa32MrWHb6yUxkcAkF3GEJkp1aLBuoQYyO5c
wQi1dGjrjLRVpdsWNQSG+8LT5t4PSyiH1aTfK7+S84sOPKYEAQzh/A8H7UDDN26x
RE/PZvArl9TYbK2eWYY30WzBJScmF7SaDZcjnDKf9+7LTc/GtB+I/Czr/r1CpFn+
X6DUk98/03uSeB0tt1v0HxmfyLs39TO0fT/Ch36dOBMNRG2JG0TM4AA/gKB5Q+Zm
hV4VO9L93EUWfZS+KQ95qPtbiB2zt2LThEEkg8AHjAGUhhKFPDWH1hW+tHx0UF6v
7lI8cksxaFaz5Et9D5CVNdNdyTmedYSfgjFN3cSxOlwgeu6MEyZOWkRGB6tOd7Cz
tIOkJdxwNt/58LKpYRJUBtigtWWpBp6chPKXD079HyMWXcmtFj7OX7i2ebJ57Lp9
B2oVK6jbGVRczdHL2E/43lXTBzhVpXaI9AZkzHl+lvBCjnM4gkz/FW8o/bszFf7n
toICQzgWirgrtRMVVeKBjml93lvsK7g4z+nwCc/V8n0Xrw+UVNoyGx/uKQMA8CIC
lbeRS2sor1h8EoiVN5OQipiQEUHgqqft2CCM7Al4a2ecrxkOLBWGVA2r04NFYIam
gf8TAdwwE7eQJ2zDa3BvHvxauC2OqfmsiSO54wCU6CMAEEhFgFUj5V12LDlWnJgW
DYo0px2rtgh0u7k807Z5UxV5eyVzKYmOl2VeLUC2KQrc+rdaGzQXvlFic8v/HAX0
KfjfHhHzQYsb1tsa77ZPGltlZ/zlFfEjHsnOjO7RekCMEOHXhW/iFaWOy+B1eteN
tyY4+/uPDEtiaJa9FE6TVKbCw2YRk9O9LPamR3v8Bd5JZsYJinoHvmV6hi83AwAt
Q13QXrGunOfEyGlO8UecpY/Bjvtv8qfTvgdRjWSi3sRpRVkmCe/OdP4f3wMddoMh
mIlO8rZmzfui7otnXivax3p6eP4EY+ORBGFUIvP+Pik471hVedBCE6fCffX/TP5M
RXwfmRe/K2cPA/288M5TED5L6OBWeX4Qlbxf3p0sP8hFrg3coNCCLbuIAOWONEre
QVri5ljpI/cSR/M+FteV06F1k8heypW0NJdqskGX7Df5XCI/Qu4sSKhkDQUFi9z4
e9qnSMqQSuBJ7+iAWfhKB339UQOr1YQdzcoCjvLsvz0PEVKpLuV79FyjP7BuBDkY
HvF8blVPHLfKS9aLYLFzLkr+qlwc0pUjWeAyyOygumNAuAM6sB6ELD824LmoAsal
s8qbPxXQfvMQGp3jWVNeoCK6c/8sw+oDzH/qLRWsAY1d7pxVA8vITCCVwsuo554o
D4ygYk4ahk2XdiOfdz6qAZo579tiprL8KSyyzW71srbpYdDifVqMV34hnpqV5OUC
3j2zHBIzCqNhzQf0oDjN5sLNjo3t/EOsk+bN0DZCq8opxZVUuaj9+kSOxLG7KC4n
xp3fvQumc8yYS5habCFsZzklb7aO9L6q+mgIv5ln7JeKQGEtD+lNop3PIuPip6Ke
dX8vIT966wlZu4ChvsCUWt3GwFYnbP5gsIdFU3x0TVP5qrRrTWhbRm67DVlOzhHu
5Kd7oGvOLacJqCkL3NEfhZgZE69ITzcw0MF189sSq9XR8AYdWkJp51RFvJ8IXD5z
/ySRvGw1NZQeAB5FUX826jRTSZjdvMRwNFf1E9f68J5AQ6hbg9Mv4O6SIrzKnrAn
edLY3nwxBflG2G0EJqqDNCk1UG2gX9BffOVkvAlw8upfmIZAjcUZgcvTibJdT9ff
mVMEt0yIJwUCOJyMvhOt1DpXTlv8X8KUpvMaHZq8a7SrCVtbt4lPUI5kdrb4UCdd
DDRoLVaP2viaHga+92hzMClq7t5gQntF7oVVq+qD7REj4yYZHp89kmW8GLSnb/nk
ZoN08NZf9nmSUiZ8k+KMwBV3I4Eeno2vBi8kqVoEiecFm3J4dFHRWvGX42hRNfuW
5J8lp/rFoJCvyrHMM+xrC/Ak3iWs8bYiIe6HDdcgvPM+VIcEF5zkl8r4dQmAl0Oa
SBFJzXQC329i4uJUbC39c8jeL/Gm6ogZNshJh/dW2mlISbrthfPByrCx4ImjU5DE
WIrkDbho96GRNqr2r2111TTkz/cy8OiJcCM37ydFZKFEqfb2N1YQAPk4S+FtWyBx
trDv+JP9IXM0olTBUANls9DM5ABIxoG9F2jWBQ4YXuS1QQucab4eRBStqBIDih/x
O8sH2gAYGfyObTT796iWAVCNE0UWBLAt636k09K0x9boyTUgCHUwJlNQjdRzee5x
0RNv2LB/sY7so/uKXKVJN5OiqlhebNVr1WF3N4d4BpGbojKfD0rOxJI9kNo/WovO
JtAxZr6jKdlIyIqWI3sffA47rOHXVW44z7QzSk7VbGgmC39mZy+PgExel0PyuFV0
F8ixQmJ7+KFoolaUMvp1KGpVNnnKM+Qf+8t6T2B+oMOTQg0jHr+XK/aLLXnGVnto
AROjrBURLDTUGHWJscsMmPgumKjEFbGf3jBPHDrK3sCJMMstpJFZsydfSaKCKiYr
XXIZ0miggJGycrr+nYh/raRrOJtx3gu68PDPm/aMNRtIy5NXm4gEYDl94I7+BHye
Iwx20p5s5pLgzb5s/7mIYZqiJouw6kuPrIchd1kqcOgRmBVFGFZQ9UNINkIhcFXZ
xp/FZ4Mbd5Irabmjtgd86oK5GgrN7QbD1zz2qQT0uSHI/FLO543LGLzsmBr5F8/9
VEVrOdnmpGiQO3Wd+YyGNSlMVNb/f5SfZsa3fD+RZq41HiMriceEAutvBTJlKMAK
zqw+0H5XQ+KUVCcX5YUSAnax4ALyVc6yrJylGEutY6Ncwy5nWSFmJE6/fqMkX67b
P/c6wQIvtYDRx5Z1DniL+/5AC+k+4TRl7VQ8p9MhVvxyWnaluCDSRRG1BrvLxe8F
DtaVwdIIqzL2is40TejsYVgNW688fOL7fOnY70f6vpU2vxeQdHNo+Tei5thLOemW
c1Jmfv59ZrYW78FAB5CSZrU+HvYKOy397bnjKaikrlSv7w5fdLqnlpBrl5Hd4fHi
FByx03/WYxaZEB7oV+rsntCiUPGVAKMnispsbSifOJZHga24DHKJ1VAiCbJSn+o9
GeaHRSJMMXUwgYxmbiMOQXU9hm6Pg+HU11LmvAsHqqU/wGfJQZ9Hlggk2YMXfsiL
Z2KG7hx6aV+C4Njcgsr00OVD7HIiDFuQylaZEz0dScQ5m8NZm9XiRxhWLB8kDo66
38k3ITMbaUztuMM3QjUwj9Mv9/nxJ4mayb9rIcJaFT64Qv5YOKOfWHPey4y/En5Y
DV4YcfykRBE8l0kihoy6lMFB5bkRRTuHOeAC7X3GLJ5xD3/i4RUnzLgS8PzMEk+t
iDfBxmWLRXYNd0fjpBuQU6VYVFmu3i9xrpwGDIFL+QJmZauaVHTT96FqLZforZk+
brRnnD6WsetrhbCuzOayYaMSzFlH4d8UrJdibt6P/AXs2Y7WgJZOqNhP1sh+jQk+
WpA0eNC5uPEYoVNqjrdhbw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
loWEy7ESx35lOuFBjcVAqaK55xtUr5I4Nh/5vL0v4iTqVnr7bVkGLByMikZMgWkD
1ZYAq40cLb0A0RqYyM5ZVkcoRxNyhmfmpMvzwjlzm/exi0r4eYIjnXPKaovEdPrc
vbEbCmwty76II0A21uCWTsXdYyTiHZ7yQ953IXiH9vSPc+fw2nBErZ/ZsTfBYWm6
ATx9/+4J+J3MAFyIuO7smGIJuaq8SI39sbKfUGrg5W49VO/rTjjNgKBnyZ6JK3nP
LXOpwDffzkBm0JmLck4e4iOziAhA2Ejo+CRnJdyH/Akdbi9pdDPdlEcvYcdyY9L1
Iuw1JJnUQ/CWcSPGUrCzng==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8720 )
`pragma protect data_block
7CrpefWXlFrYk7y/bpuNtMoMInBmbB/x3Vuky4Kksk/TPBbVuZHofjujcpkl093v
7COX/SX1I5+XsEiKQoY0kC+Mcxx2npXcPABt+S1xK7i/bJ+/T7ut6yBOQYa7Zp9N
gXy2NDn2e9nK8OqZqxuzl0E5wi3rXI3MCftRGN50WNWIXi5cLUtDJ3d2+9SpVKI3
hNacb/SFZ0HgzVCCO7H71VhWFyBCA/PfKQzO6ocEeNRYgzPCJKXYqWKCtXBXP8Fm
M2WC6X3W/zMPyzzjjsRWP3dASSsgdGattkpgRvGcA7shLP2QmHHo31fxGXjdoXH6
lLMlDT5CkFFxpU/bQ9Dkap79JmIIu9/sHi4EUguNrI5cmpsWOlVqiPCEqFzFbIsB
NXZ2B8nsAvPhGAQDaxp8KJgE/lbuK7S7a1iHmm4G0olHmVMqDsqTd2VmC5899N2f
UBXcd4FlowvKV3usiMmH4iB5bDBCeAEEcCr9DyfBFCur6zY/NSx9gDLTAsAALEib
ujQKdq0nIgjgudKaBCtCr1rcV3UM98f1oFnuOFa4fxoQyRdQ8K02a0V0V2008M9l
dhOrY8PYwNCAjt4PosRaP252grCuWuav9DQsHFmgTDXZRoFNQnGD3EVh2fGPQ6K7
GSG4wKcaMPTkBAKENEmIr8pjS14+K3pDjSIhYbSu6RHE0TbpHISJkhlKtaJkKG0d
mv0F21rxC/w0MmBRHGukgOHNnmuds1QbRyiZt73et4IEYaUElcX8m0ZynL+DccN4
n5vDigM5kSh16lF89oQq3hSlKYR3hKjU5q5gN4voGaU4deFRys70ybr9yVBiQcEJ
E7zA+iB9VFou6EHib9umSDvPH9UHfYzD0hv5igD2RQAkFu/+FMB0CvMs7bYMDIXb
wUeu5978IXg7Rqa2KAaJzuejgeZbhKzwo7CxipvVVtvDYJ1M9uBImxfzRC3sf4fM
QcMiWdRdlbLsVB9DIdkCCBfjIegoo7d9YiJIxEgYmAj69pjP7viCotdVaQxbChfr
cjfsOQvC7NKLj+A920YP3Zf187MbKasntotxumZ9NhxEjxwuZB3zQWww+uDvwSoJ
JtUB0bhDXFAWOn63XA03zuwYdjMiIuCZWNgU6aodNSIxRNZ69xftJNEYbJQ+qv7y
m5P9eBuddQqRA1XMyKlqZzeyKEZZ5Rgizeyx+WKsIQbfwFaABAM2Bxc+TIfmkKeq
HT8oki0+WQ0JEFvqN/KG1V7KrYMZ9kctBYf/TA48aPGlXQXp0YFBh/hb8KNgJURo
+aOoL2tnelp608RP7eAj0jfoUGxaPnLlmMhhXE8Ph02sayScAsd51C6S+Ldb6lOB
YLcvy7SageN1JPqVaE4DtHmbHTpcU+Cyevfo6MzR9MyECYNEBrBO/S859eDnbfXb
NRZlDMquyUpU0fslXzF4/nEuAR/U009i49rOkF2lRa/FI9d1YSAX79vzUmf1Fsj1
ce2bu9nTVkZU0Flj3oBAb1AfdY5iYprrTU+lBX7VFpZpWQ+H7x1arxdnwyu60PH/
p9xFwPoZX2zRBC3ndVruxMqJFwp9TyeHXA3OAFFBP+PtHa1r+/bbaBbwlC5+E5hm
rS5nHclK5HwNzZles1ymRPRGw1T3dvNQzaMS08aWJO4x8hZszt86PonTuH9IMMDC
FXiMMqackE0pBn1WJqzqvv8dbRBT6DYhDujwfTueY/Fcni023YzBHWlWF/Dx6Ppi
QqdBJNvPBfRxAcZgM+k+KsiBy83VuKSwKOjN6iYSFTW4UoA1bJR3URVMDtDIPoQo
pzSvYHxFcC5stpi1O1BnZhsx4H3ugVn/6UW82vUbNkIbZt6kRORNzJl8b3aI5DAc
UY0W+JGbZFfjLGRbShVVbhIE3KH6bYt84u8zXf5DJ+mou8jAzNQFMYMt7D2/L5P8
U7RZ7jNbzmyyA6c+V1ZKhJws8e6a5Wu2wR0fPAemDJ7fLfeksud5YlDQMiTVmrZw
fanO0JeF+qrC1wLEO7H/wsd0Zh6oZJEhm2rITkEc5XmUMCrO7KOkNnRH+EBiRbRW
cuXe2m/iPbGE3Po13qrPqNQT+kkQ01NPddgIHyYH5qESOt0K6ipIRC+ohILTI5td
NxE1TJ8vFHz44GAh/ynBiQ0ZVR+CR9SBfXIpAp0usRi9B3OC46w3CqXAO1emkVfB
dYY5qyEQqJvYC142wXw1kVi3eOb8CaD3ymzHhX80CgKIEb3uBfjPSUSDzTw5mLmP
nz23ONNKcpbw7QzlocFf9i3um8ofNKrD0QuJKIZdDC21LGq3UjqbqctUeP+6cBGa
Lyfc4LOEP0hli+tW4sBVJgnADVqeK3qLsSP5onlf+xNJkZYcq9Bh8QHK8UtrphB2
1xcvwDouS5gAuW7R9AO94cCfVPtU+4LB4CQMqPklm3EgPK6PCMhDhoQBWVANrDTF
eK7AobnMLbQxqa2H4iMHtsKus4XhPjsvgjO6DnUEi1MKjBtxQxrme1URyKKle5J3
azb/VrK2MJDA2yW3jW/UxbwoWGkwOQc7yLACKHq7T5S04aiIdDENaeT1x1hy1203
NLIYZkAinBpX2O12SfM3NluBWeafTLHsPHPFeMqxNHqVuleAa0fzv2TXGz1quSNO
e7g0UHingfdZNdGXqmAb4RTEohtvywKtBTWrzUkmacsZhMrImMB9d8IDQ+1W79lx
wZ+ol/l0UeFIdo1pj6htUcyqhMzeaf3Xi8x700wYGav6KeX4qDueiWzicJWSamD4
cv/uTVSiYr0HXO+u8VlaE796ZBecec6EesHepnU0EAoHTz/hRs4dL+4PiMWobZdG
gA8OgWAiqnU+u3+vIczlCaHgjK2f68tgcQcQXoj0yGJqgkQacaV7qPrr5S+RyQo9
xgOuCaXMtZqM9t47cB2jyryP3/suHLEWZw2KsglnAst45upm6RIrnxaKhYOkoiH/
sHpdltp1B1hQgC0rAgklE6FpADDr1B72Qab7KSHz4GoXfhIVSAPFdd+ZgqpCI5pE
jSnzoTf5rcl5MN9HwjopJ3qwkcQT2/wzX7XaaTIbo5M7EcLjaQONJ9PLPxEjXD22
4oYAid2yeuND+5Hc2dHYSRvcjPCC+mj0bOIfryxLhNwAMX+HZPeQG9ZeLLU/h90f
GlbQfN3ck0sRo6nI3D3iBCQXBoaETk+bMuXlu5mHnZOspgg33n/9o2f069MR+eDa
dva8ADkFhhksWepW2GGAgSs9X+jj9fo3jxaoSnhKbd/CIch8X5YP2lRlVN1aDq1a
H9oTYLCwUxdFcyOTpvLxyBtXX6cBO91/TDedlg/584jVLN+1P9dVLQvnWcjuAB1z
MfNiGWX+4bfkLc6wJMG8wGXq2Z6IcnM0T4hMM0CK2taDsW6MnR6f937hl+mxaia2
CRAYU5EXGCbQS4hpXN8d3HRW1LzqbfhW+SQ43xQ82WM4mN+e/gBZfHnhyfXdIs4O
n6J8rW5HlqoZ2cM/6yMFActQguMSFOfxFZjQJq8SlO9m+E9/Y45weiUBbXkHdeZu
EFOdMQbwIkEygOZfYdaWLyfmWU7c+GoM/xfllBBKHaQ7b2MjHrr5sMzXOeBHaITA
1Tfm71AcFtE4PVjGj5zuyysYbQEhZKRSwt8wLbMxrPqyZxU0+4r7x5x4myXg62Qh
NUYyFxqEytocm70U58GxMFYW+RXSrbiBmFRx+N+cHsYEUybSXcdnbzCBCWZz4NGE
D/6s05yQekKpI/Cxpxc84eEVnmFngSdUh9oEf7i3V9wvY9WhAx5JTKsiZtbak1ON
lCEbZn7F8KB5kwSITJDSe1iViDUWtPrJ+fsvvn+mdiUVsuXJgTS7AbNK3HPF3wN/
zVW1S8W9yQi8ZcuJ73abF6mGkU92BQC1xzO+s71RXD4XvlQCs1IAHnWc26VKZGaD
OnFRzoZZEFLn3xmnCD5A57cFGciJaMN/GiN85yzIXBSExr7/jkSgPEltKg8fZufy
g6InCoaTpG88h9kC85S7NJx/xOGOcjVDpJd7/wjHs8sxC8/XpIMmLT1vTv7qzQvi
jArkKpidYSR58x2kf47aFbBNJkKlIZZiW8JcKKbPJ0ZOH/LI4J5HEdyrZe3cKdst
TMfVNa+wYzGXX5pZuy9uKw6JknA6n4tIcqY4AqXghDR8+Q8trjHouY5Lc4O9kMZ/
cy93bFub/FnH/VetH64xaRx+oih1Sfgtp4cjcECunxfnUit2wokHSFryJOtWonZJ
RZi0FTkz4zXXtOPYWRFbtnQ/GYKQAbpsc1W1qzT8cAqR2KcAXLkqv3peoSKN97ig
1BdtWSH1OBTiSpQynm58sU6+Q1o58/6J1q7I2Zqb1tEzIZr+/dQeSgb7Ldx93MCU
qQmFacjDaj0O6Q53H/djxVhodSmLJI4ZbO6a6pRKbTYjiysYj8u1/9BjwQ9GpSLG
lXXjcksC9QIAzOXhkhl/GtwRxDOVWd/3awOWWPbz6qMyUCpHU6ddWDGSWYtt73qP
4Z7PI7ApseYTJ3e2bG2eHOThGBB+tXdavtxYMdpVSNYNvBpK1fPV8v8ZBFxp/jt9
T4eR+KKqdW+c+DUU/8TXbnBZZgYw5LrWct15XTWpYbJC5Iwlv/5CYYViyVtUVEun
NSIB8psdUP0iNAldOCL/D0enM6nmnv9Fj64Dm4mceBGW2MPsGNDe2W0Hq5KFx7IK
elqfNDAJd1rwliyv2+TRNTeM+/X5/bciZPtNgjEd/5UYmBlT909Rk1Eh/mibeX3r
E8fGovQai9nYWT4oc4/vaeiGCmfATI5L/jp1o5TjPDEx0jbWuiiJXovp0jbPnnSY
67UvEfvNwxxaGVaSMtV2UD/trnCKwBRpBfSkWbyzzP6csoh3AQXpZnoftWf34eVe
r+gmP+ntfxdORw+6uEN+Y9+PfCqRDQDHcIdswz5s/avUeKlSAtngXLICgi0Yxg/T
iyumgLjC+RIYCmbaNRz2CDkNLY4nJ6nDaTKGT90oSKByrnxiuF4i1B/0373WXR7S
QdrSReTNr7UrSpZcsGpWGqFRfQ0iBtzMs6pTM+SOZLCb3kboTamDpX8ab+X+Pisa
wmbbOjhTdykmS/sTPB6CDnAI3gGV3ftfO80WafNnZRhan9mzeiFG6+b2pg25aGAo
/QpW6n0XW9UxHxltlyV8K5U9TUdzielC2s+ZSuTjZyJg/8fWA7L92ho991lwzoX3
4FoUwu/zKZD42MqdDzGi5e+7GYDZPISrkHSkiAM90M6t6L7GOUoT7UpGBwBcbL25
AY1rhhz1UtakUI/KdrGu1Jgy7xsSBakTDPRCzkWMyk+T1OucVka/Ms0EyFvXiuAW
kWn0FxOS+yV4A/Z9IT8jz1VSarLpQ60LibNS6b6XWJW5XBlqfxlplI+voUXO3+NV
/WxN+eYghzMD0J3clUCQxize55tT6s/IiG3opBnh1zQreUCjz8eGhUvHO6aTtqGy
Kmv8WE2P/QzctRLDKt+Uthv2qfJarv1ZEWCAzIKxxScDKjTjV/eJPlW2zlLMbhA4
zeHP/FC/MAcXQhnRKJQ8zn/B+Jjts3qoRF7PRdREkNdYyTvcQLaNv2T08ev1w95K
OaCUi4W+syjRhbLvhHhf95Hx0DsF5NnZ6N4P4quR1qb/Lmsvue/iHAVjPAwpNrUW
EGc122BkXaJZKlFgUUJPwwxwrKnsku3YpNQ1jESTsijmt0Qxf+YlFjfD9fgX9PEa
/l1WIIFPWwjA9P8J11f5bVNM7pgPwElJ0JYV5ElOZB8SOpRCbmuXmqYlmNnts60A
0qidLjNGTf2SvC7D/f+nohEJcQaremhvec+bn8fJsuFXnTSAJSm3VSkwdYWTYeGH
I8iC5aDSIDCLrB50B6K3cZDLxnozgt0wGNMRCm1p3rm1lvY97DcSeB8dRG5dLfOE
an38dgKXktk5hCI/hk7i6UasTdt/XaPT4w5PBzelJ4EFFS3tKWyieu8GfC/Czt5X
K1Y9+R8qXBh5EdVfgOo7G84mW7J4oWVCmnfoI2QOLvSpKvkL8/owXsQFyVMcU3i2
U6AsUfX8in5XdmL8ipVON1N3OWH2U2rBGo9R0pI3VSFxZ9++NEhZxehO+lsLZlll
gi3pzzIicjZ5o2fbXyu4s8MnIU+UxXq9suiqiOioD6uhRboKZP/AXwFDvBk8SO64
wOfN2Eg6w36GmSL/WKMvKtUnzTNZBpeRLWyGyPtvSa3YvhYlk8CrOy+dhIaKHHHa
y1Gn4b2lXlRxX+17zYHpsN2rVAUHEhwftXHgwiexhdl/Dl0DDiI5dUnjoxkpnD3T
IIXoZ8a7V4+FmMNllrFh+pS2BcVWdJ/ywSiMTbq7NIanlKprvmGdp9ZJCNGpBV3p
RkzEl5BhTXFFpeYOhBlT+xOuysfzZb9IVXqhPYKlXu8nfEDWtwicmByU4SygW90v
PMdabs5IXn04OjN9h8/hSkn84ZOWqQIXSkqzZGA8boxB43WXHk2MLdMgLNg7Stq7
FkrcgYNz+vX1c8fmQSRPoe1K6ipdsNvc1Cg4PF2NicD4XcOoexI2sGcWnsuFwTu5
2Cd1LpS5C415sIcrt3YcVrCFaVs5y8yKHPtqpfYf4wry6zJggsDQ5677jmpFTKlw
rW/LCPssMkIuZV9lGu0JwxFpK7FAOEqsBBm9GPUE5CUUevK2ckCfVtQd4MrPjXkt
acPer1YOjxX5xMiVp8Fq6feVrEKDP1Na9UMcIGsmd1/N3eqPPAgWs/NIniSnWl3j
022Aqlo/KZEo4bZg5dfXHfRNa82o72LXMW8I4WU6OjMUlFVBtEne7m3G3mTK8Dp1
+w18SToXB42/liDmfFGKOQeo9m+Ba8csaP2aONRkwMJGgk2sEOP0m9JRu8hqRfZe
Nf5VxvXOyYvFNRrfaVV5ixG0edJp1GUYu5qUe5GQnpsAwmyfARN8opVY7fYdO032
NY0Ukff75zqhaWzHxCR0cBNb+hqBJ5jU5Q95r01hNSbbiVGlNlsJN11kjBkkMrwX
CFnbW1lSLFc5dZcLrhWYSMv8weFlGriNG0TNhg0ndOQkVoVMHYSdkmQtTlOVefo9
N7wFxjwalHOEcn6qIC4Rx4GKb1BmKB2/N0G+VEoWG5RH2IPnrWggQjmaYgD+wsHH
mqi6uYQOPnC6RrKr2pEGQu7ZW9kH681bdNWXVLOPDOVezCGX8v3+q0hGx4A0IcdP
lprRCy3n3aLLPbCV2PQ/XZnTLzCiETtlcbLINhkj7MfnwhC5R2BEInr8k0XHhWed
MSpoBx+A2FBtU+5o85GESXYTfz3FOywhLplM8a7R2ywQRAcN4/aWO2kGhSUstkD0
Exy48a9ekrcImUFTjzM/1IUPU5njSdGDkVUOSvpPQo2B0nlwCe5/e6Qnr+SXBUK7
MBGJ5i6kcgGBPpZyDLYa3PJly62tFG+KgSDIE94JSyFM0U/2NeVnFIWpQoGLtMN3
Nj8shOVE47CWcaU/EkfS3cF6DZu1+qGwdvje8DjW0tePuYMkXc2SpjtbsE32gi6+
5b1ugYWSQot9Gh6bC6r9ehnHJ4+f6ggzXviwJdJ9OwrxnizGKhMNtMJvqy3escMF
XvtiPl5DC61VJrtBfIrWPKQufYhz8vFh5z4W+x+RUPyXRca8XB/YKBvyzQ7gdnnl
12KJ19TPMXm5arEJmT12n8NgZ+H/02wuyWsi4rKkSNIkeJGpJKma14H4OOq6kBbh
l9AGPLyAIaeosnjdYTNdn122OcD0YdNZBS5uigeDBbAB0xJHU4daiYQLZH7bYJzk
rHguXRoFlpl90Fi3Qwm18EtY6wFbEydbtaVo2tUlFfMgjVnXKNuL+wjjrqXCvFb+
cyNZQvNFtZvjp9Vkz0VHX4eLDZcivuV89yqV26Gx41PKSbdArsGdwQiYdBRH9oZo
ZHQUTblcejCMZ1vpAPbymKB+ea4yFaUHgK8luhZSnFwqteV/Cc3VAo6Syg57Lx5t
7uGDh776yCs9v3hUf0tp4f1HkxJpiU4EkgRo6Bv6cCIe8yzipgsszkdQH8evoT8j
MoUtIVw67k8vSDPpi84JJgY0yl+u4tRtE/K7FbdvFzEAoov0vR48ujlVWFHZuhcx
R1h/Tv0YZRRyJb1pifgBL75J0ZdmC39vB6ek7SW4DLTazEknYxps6P/hcz668JCl
VdrSe6MNILSpLKEfcnh38ux2v/y3nZWJLGO2/dmu8Q9ljwnOk3mp4BxqAs5/BE/2
cFhlDaz901VaIcznFJFmzWONl4FwKUHqWhycSW20NBV25R3qgWP2sXVHv2MCVV/P
xml972GQFkofWR92yMjNBqZGQgKXlhkcLbRqGyiCV+oO83o0QKPOiN037QVMDunV
zHdrUkH76e4bfw0bxeX3o4WahP30QI4KYoP4FuFLdeDXU/LfmoBpZnFgM9HJppBN
n73DCp576HkncwzzHrrONwqXc7fvpNT2jGwpDfNFGetVa0i/fjvoYPIxELXEWYlJ
aoCKaQgYxoFgOOmoom2iyOsCQswX395zIy08N8KhJBYJyp88ce8+/tnaYPGAYowz
30zmc73vQfKe6LQYkxSOG/VDKV3DoA9my3w1H6D2qR5gXVhAWx2HGhD+g2lGe7c3
J3KdNfEpZFNC/XJ91j6C6gXqlp1HoucDnXtoCZugsaWJa7L0xs9iJ5jty9eAm0Lw
lNNs6x5DQKQgzIuIgKfT9gYW+dWpYYCd//cn+o1yGRGh10cIfViPK3PLSvONY6sF
a+u7kE5gUDAwZX/VUeRf15uwqrkQq7VKp0Gdn4w7dQgst5PAqvhwOjcREVvgaFTj
vTpTunqAXFMkS9o6sal03zb7nkwEuVZMvyQ/zbymwFgrkygay1PMF9VdU/7n/n9g
vvMxY1s+rId025riOyEPTTHLjeYLiECkU3OeDdAtsOqmPPLbVQv6nYTRr7sUZV4/
8B0r/htASPIXLMCsagtEpusifzvrdpHsQG2mkAxH/jeu9ZJ/NQ/5tEQIFP7rsiQf
yEapB8NHEIYifhNfnqHj++AecSlVwkT5e452SPGGQ/3z/4UBVLH4Zai/kvoyb8Ft
gDP3y2Y7oMhScriskwX5oe48o1Jn05aQpl2zv/BysYmVS0BR0prLes/SeCkSeWVK
Umz8Si03+PP8VYyPcz8y9lUgw1K8lAppEhKIrOPh6oYeejAtqOmx9ene8Kjskfj+
cC9Eawxm4BCdxCYz6dXV8fsjERtCX/nIFE/9MHZrmt0sv3E7+lb7wlyDIvMrJBO+
pEUtsPfK95/ALdUYo7WxOmdipn8GRu4Ar6raaEbkEP0sxvG5mSuiBnUDWZUTs3S1
6fERkmiOUTtkwx3Sbxq5Q1PISpE/CVMV2A1CKHis8r0F3hR0SLfaCFYay1NB44Fu
bkLZpBsHCBceZnOW2TDiEAJoEe3aIsTfUtmNqQZRRg1DGWU1ORfOzshrkdWX9qy9
eOCbqhNebLpfE8P/g9+RB8M7Dq5eql2HI/faI/N0c+54sCX1rQLJCO5o7ZPQB/w6
zBsMcMKkoggmb0Ns7w6OY7eLnBNd+mD/LoJhXGcebqz+R9rmU7w7bbGiwA/Eh5GM
oXn/YuGb5IQXhn6mD15JGND9km2mOEIMBshYQzpcDk7f8gXk+JSRHnzldsDwx2rt
YClJTQoC09ySorFT1LT3mIJ0pnyLiOKkbJSW8JknN7yaTBVafomWwI8wjV7EZyvz
68sHll6AkA7wzKjkWagzakAZ5T16wUAAd8BkTYJQJIDQykV06nbLzn1V+FRvI+sc
cP0sulsFxQ3iPOUoXAA6OuFBrNZmtmNXaVsF7At41veaoJFAJJdZPEPfwEv0uIbS
d+venjAmaTFKL6vkwVi7muxaCMpta/tIW8fAGtmX0B25Ren1bI0Z8Ah1IH8mrbkV
iqhErGkUc4WiFCtDvhGyo86m4yrlu3uoxNK1svWN9HQAalnnaED9NBtLkzGzL6aC
KeK4CqGuYn9x2CSeu2XHYBl310AJ6aD1u4aj50rlnOQ5FHV7wnVj1ls5duyTzOgw
tJ64rt5XajfUiOIPSBktbi4vw/3Kxw8lMsnRjyvD1ahvFrRp1DhSg1yqK0mH7MwR
IWlsTiPKmBJ6wYvYcrGSvJzxE/BOpLOyxd7oxK5NMz3zdDLtg4+LEoCclH2prRYG
FpXDfH5qwbp3rClXosf8TaWWFg7vKBLaLvxLpv3t6MLZTZpvZIhKCbY3sBE9quqN
67BSkZt/ldqDN9tYkt2+UlYagXzj9x7CoJtuggvMkZgMcF/wZUhJUOT3+fyc1ktJ
O0hKfl1++1WQVf6cmbXLKZ3BSJYp7nTN3Tn7HEl4ZFDIQQ0b01UnsetF/sDhyPg+
DtXTW0l24vTG9t8ACjNkW4YXCAQ5Cpmiwi1fbNQAU7ugs+aYUTfVG5UPbvhnHDT/
bBvieV9/jHGRLUSVGHRgcF7Cv2GSGxLy37UZY3CKI/06oWRNURhjXmV+OMxnnu2+
hDWlChso83krYkOrzLAOvaFaBw5cLCKjLjcai8yPrxRz59QH2UGkmqkU8Fs2eKbH
wMBtIpPlSF7CJXzZku0+1gui+mdFMWbObscFrcexbpJtdDvsUPeBHA14wtwr6C6V
Q1HtLgkJAGt+LS+3S2Hd32PRDDbLdDs2oaBF+ZHOPg0zXGwhUl1M37K19W211b9R
9sipX8Tg70BQMUOQvoCYrYxs9nelvUNwVXPY/mO2LpXPf0HrxqP9I2VeDhfRoFO2
dam5npxL+0KL02UDSDEzsvppZKpJGkLaTbUVvbUbU0a+/1DTke8gsdA2C3h/ae8Y
XgWTmkMd5xp5kdO9F0DHY6wpmL7TGg+yK2DYHTDxf8ZZ+sgCxZIXT+mWN4Nprted
fdD2ca47/8oHqII7+n00HHQNxAUMTdIepdM95POPGWc23laDuLPeMrh4rvtLWRh0
DK4i/69esZnUntEWzk99uhOfDzmzQpQXKzRYs+9uNw/AjoS7XsKbyIYdQVpa1Llc
fmJrezHzP2igwqDBTDYihAY9ha6rCCH6d2h7rOWv8E9xUTekjgO8iSjpI5j8hREn
xzv/NBm/DAo1v2DSjh80ABNBkaEej6b2ba71R4uIAFfVahrMi1kNcUbUiI+KNp7O
wj3e8QyYQgGS5HNunyRZmgVbClIFYuqRKLDjxuhBxov3npOuqu8DiP7HRWWJQcSb
XEK8WhXpuIGYANbV/7oeBMKgtUK7YFAn5zZAc2txlJ0kyb9T73sgAv7At9ZaeaKd
UUdrfwlnYqJGC7HXUsF2Cno4psF2qHKWW/t0jos2ERHeiWOqrVF8EJRQ9lsDe7hU
gwTe4oIYGi1Yo9DVraYsqP0oRTqpH5p58wlG9K33tDAjgKxeT+vAkcbaYypYx5lu
Hg5X8IvqESOIpeZu+3YFuht16DMa81QlRG9dc9+Df2pTnJZzC867KH0bhZZ7GAZZ
ElRwJ/s76dwZIsJNLr31DpfW9yikk2yIWtS2dTYAnrp8n/U/Je0hIxsLrxzEw4mD
vm79vXdDe/NeUzUhlAc0oHrHxuzmzrp6U3fotYPnZDGtW0AKgK0X8QNV3V6L+IQ2
lzyypf8BJvPBSfaw2jaIVHVCreqcx49xPgSoLBfo4XL+r4B/OBJrfNnUWc0buijv
k2MvQQxh3aBlZXw9JYjDlYO739Uj0wLQqbg+xctPqcY=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
feCNIX4wL8G0hryagrSLy2Egi+OJx8Adz8EDDCOL9tb3LowLxS68x30KHcpMQdX/
oaeZbGJaB9+JG66UiedsEdc8wnhtT3NMgivQS5I88AT5aZXI8ihTDF6Xv7RTlD/K
ZuloUogex9NsJP14Y41YLXaukofGiPbxfdyA+8Y39st2WoWGHuAZNKAHb9CWoQdx
kFMG4yFJxA768VpIKbHQtxAnXo2jab0PO4z9Uhi5LdSgTo+3LjgwpC/uZf44MlVK
VTUbZPp3neu6J9I5H2qQRGlNb1LVKhV/0SUYobwla47XzuWZo6F4k0AGIk2FvvxS
/BJIg0avO16g6UgRxp5PTg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4336 )
`pragma protect data_block
YBGJhhoz5PWNGzyaZorZ6wfaZW7pEUFssF6/pZEPTG6O+LmPZYLf1Jxcf9GyHL4C
1FtHNXrtrZPBvlqZGQyyOdVsigGFSbMyk4hg+CiAVTNqfzW02ZAdfsnM7Oyh5PNJ
HQZOEeZvnENdyml2I/LHTHtwf9emAtdvp7UYMbDOH2nNWoM/+aVL06TxrKgGmAsM
bkQpr5oQiYym7ky2nEDntJcLxEXtdwcUo5L74mP9R5nreUBAH4a+J++BXq6XHtzh
kehRmh5QJhuScKFJz0j4hsQI3gZQdMw+9rPZX8aaSV/IvddviRTTsc4+N5xXp5yv
jvqG6e6M+pJGTpDGU6FXaFWwYKpuD6PYLS3KcqRv95tjPvctaqNaet306QnvSRqK
+o1ZWd5TSBNbEmmPYJI5kXaGUEGvGD/dDpJ8ueha4x9GH7JlpbkFgDAAJLP6QLOz
NuGYvQpZs6HZx/KQLI3xXdh1FebJm7u2Vs9ZpsrDcfWXypwSgzPgBOlY0s/LbUyM
J5y8aRrXMByM8smiTVaUazVKAXGVqRo4jN2mf0Xckj6n2mQEesAji0EpVDo/WBUJ
wD3UOwc9nSAUdBEtBUVzACcVTkiV7I3ndmymOVJzSS1zSqlRIkNUcV2jQYeQaB6/
+Nk/ZLCXSSBm7qjrlmnbRXb4RU4JbfFhpyDCpD/CanAdnOgoePdt2hJ3dZzQFE+f
fmvfI6bcZ6jZR78SSv+GcKA4GThtNakueAS7/7MjqptT+abMpGinC/0mi8jd1GQS
yryL2VRfnX7yT1pgCxxBvGs1wU+QBFYglJL1t8S3Mglnw0yPjgkqx7f/gOyAkmqa
hkeSNR2QygavMEJnopL6P1vbv8pbwuxdc/DoiANkSKNS04edZUyB8DFpdG5SuCZR
zFrudTnJjzRmR93tA10nJDRbulIgLN/PwMyh/tRGVd7SwHx16NaGYWUGRwkuhr0W
PA4Q1wZ9erXaq4dGmqTktPcevNVpjONvK8gj81DKmR2+awpz7Nx9qXpAp89K8qRk
aEkaka7t7fqA610eSRMP6JLtDgELHX2Tw5TDYvWRswMMRbUaFvDIcLfEFtyg4Den
bRSraUmjiZJpVKw76idXr6hSEEs46MREQmIZzMQnjFAA/eIw+qQeAW2sYFmC6//2
lLSSrG2Nb1Lnh5gP+1WLQq/0GxZ93awqXYtbTMgH7a/wtUyGA8IE3FcwUnRTwHkA
U9jmn8ruXXy4wWo9FjGpofdMT4RP4Be4cQWVehEf5SeW0PK5aLy/WaBV5kjSuIla
xVZCI5UTiDBh8HhYCpw5UTxrz5DkEeRx6lKyxRcIBAvoPFgL5NmZDp9+RLjkzMXj
EvMBrRGU7jfvx95NixuoJweq5O/D30vJsG9seiyJaMfmnJ2GiyCbgwtTLhtpp2x6
1Hvpsg4JI1ujnl/ANOqGorSoam9Jbk+F+eSlEwygvq8BHsXQAfnWgE62myvbtOf2
tWAH1AXpqthLBnZ4d48/IL/WybCK35TOcUEjvUxEhxMvOyRl59y3J/J3lckaWZ7h
CXkwsegZox27dZ2fNr3hw/M/xTO4hQfEWRwgjjCswUj8Fh4eEedRRtZMrPF3L0/z
vMgV4d5KGKed9szfUSImPEAfqv7UvDLVECHqf1bp/RPP0q8TPV44O8f3ZoNIzhaU
pKQkftbfVouSwB+FoEXAKQiYeELyXH/6DoFEYuGqTfLH5EPG8LJjNVmAeirfAszR
4ooyg0AEG1NuJyl0g6YLJz74u9bF96TbA4eWDDF67Q0SHIR7eMm9/7UMSTf13nvm
7utcx34nyBYCjV6iv7SJRM4i/rx0bIEmgIeueRJYKquoVwIlstzn3Iav/W1D6v6Y
DdFhRO6E/ylfPKUAu9D0t9ow7n2DHQKfJmHt02j9b3wU8jn26bLHZslrXAx3xZl5
ET5izNV0NA0aj0YrXJfBfwvWs1snGUVYQSsEl2eQY6kDYFHGQpsJ4QIKe39v6tQg
6tg/SfJ2UCMJgnTSzL1o5eBmiCwU4Cm5T0cy7EMK4emxKEjdbBxQFMTfuioV0dka
6SdJYWOtcIYk7IRLas5qGCtAyXoIY4Z54fS+w/VJM5wiCrkeZ+gV1avwHIQ+i2eR
dWNEHsbXtXVV4kMyvTT834tbHcTMZwu4cvHrA9EeMwtD+XFHyZJdH001jkMeUZvW
MztxngEhjSibXbMt6Q9xOvtYPQYBG672hg4/DczKb3rpfSZVBouTorinEKFqLhce
MbnhDOdOSTBTZDkIdeIWmKdo9GHzQhC8sVJ2MQP+oNxPW+8MvZCm/Cmpb67YWsvM
H+dRJMLoNgPNNkUFLDu2zKdF0x5Xiay9Mnu3a1XIr2zQTVhvAtCoZHFJV1ZOFCct
wZ+5At9EOWsPLidxYEuCNPjM88qSHjDV7MQp3W8+hMzLpr7TccCfFFSmrrMV6IIJ
zNafcEpRox6a/rl4xSFEcQwyBvR6rNaF9/4OYrnbVsaddFlZHV/rAB5QIl7/psKD
juygXSTyH5LPsdnhfxSuQujckdxXDP4QIt/UgpibKyZZvsQbMlwByUKgwNSy5y77
vsdUAkkB+mvFG6xm89Drn1YPYKjb9DnZ4erxcQraBFlNwmmQNoZ4pVBsGbfoAhyu
NDFajbjgUpGVBputMMqpR404TPTOrybksst/y1LoucnVn1XxgCO8AK3I9ksfZrHa
VO0/voYL9kY08KlvxP7J2ar/iEEeo2v/0GAJqMixwD3LFjER3L8IU9Z1qQR0ptbA
iTMX6DA1GoxbuvdMD0LCoen3UW7P8YifCEaJVxp3qR0JRVxE2RX3oH8BJbDA5sva
5IUCOEe+tKFYWcU0nfyDWtXjkTdUoYKqA65RDLukCq1BpjcwYtIOeQoEP3SyCKea
BvqeNascOz42VD86YPmU0G7C3MpHar2UYjeZ81AQGC0F29bOHe1XrB3MrGbkUaPP
iBx1gBscyyiPFr11+1eTl/mlPj4Me58fr9Yc+NEyidybVmwqkzXaDOngGgyveOPd
uLot9fc20estUW36OpAiIUkUNh9xnDsjldXDRoh3Y96LVr5eMjTXh3EjMlJxK12Y
OiYGIHVOiXEvVV7SLjTU8cx4W52x+OZzJLdiHiD72zus/eM17NcJ5txYNKqsowGj
m4T6XxqwZcvsmQqCCIkqqFXjj96I6xXWNhiVHTqLG1JkPacSkhaGcBVlSkPoRsGM
IkEJRe7g7wU5M/1hjQVRgzjAfeyf1T3pP9IQLI4SQemnAVQZVQ4YDnyXKwm9upZ1
Sph9O5VMUCa0Lp0nP4pWF7dD9LyrcRT+zNj9ynIoGvnixd2kpfUSYkV3B0e31dyT
uCRPauaCRXcqqzlKhX08QXA5w9oanJ4fIKiZJg4c2d/ThArfn+MJ1KFHmVugdff+
m/MMl1n1Q4v9rGZXPq1UDTRmIkyBpLEe7CTK9rhgTgAMHIUv3mojE/E1rD3/w7VG
0Zl+XeOOwcPCtHwX4+NRKw3RDVg8eAj5yf1C6HFB3X6V9GpxLSBaKb9SamLloBjW
pSe6Prdw4uh36aiORgjZZUoEMFJeqg1hVrRBYkBWwE3UCoLy8I6Ro9CefdbWR7po
4ZAM9g23frgPHFFVDrML6XjWfYpdoB7lRQowbb8x/Kb9TBJwM942GF0ekC2m2J3A
MooNr+FwudcWOPZKawX5yHEXZnRAhQOId0hjcnCFQvvLIWbJYCdPJBaIbcBbg9Fd
LT36wX9uBnWTFpAUdzsiff5YlbQDbBUMnIeYj/OsxHtAXE6ZPMeDnII0319DqabT
R1ZloY+xE3m20IMoqbwuG/LjHQZZAd7rtmreXZLrFI/8khCBTvbW8WRqJdkft860
+R1a/kff3P9W2eJMwcIzLQU6RNZuqZ8cgHeTGExPNuGhr+oMKbfxQaitnEYOtp6v
8DYmh1RWVpFWa2OpBzxWnyRPbRGgcHQ7Ce85YdXFP7Io+R3ZNQc15gu+3CXZYzuQ
SWMaux6vh11+ycNPO+LtAOF0h06THnAxek4guK3CJjP64xq6cDq5U4YysmvhQaGk
pSnwTCD2CKiX3wXdPBoujVRpgKZWmq1eYA+6+2G0/U0uKSNan7FCNJCogib/gptG
LmxlY6Vf6GYMhJdkrCrO7VO16whOR5y3eoEqJgYF+7Pdz306fyBr2ChAGtl9DvNF
M1ccpczSo9iM/bbcBK8+qOeTWRcFunVvgXi3miGU0P8Ey5CAC2MbIviGAIHsmAYA
Wlflov7OGuBaUbZeIxtkvolBJqRyxr9SEHfim2YEyh2eDg131+H4U5jAK9tgANMY
+2iVPQlzaChbQSS8BWu2TRlVJfBhJ+KXS1jt4Mq60Bi5Jkjb0Z8hvFAhCV7YtuL9
C8Fqf837mrYdK+04DGsxGwc8APr9jzg6UKoTUdx4+HH4eVAR4EbkXQgdEc/DMzds
NTtQX9VMbpo1k3rZDGhvU2HTzcScS2ffMkbbleYlfROBPVG2H1aPX9WnKSy5BGSS
UYvtfaPJGN6usL2H9qYMKjMiFfR2Gu/ciSbcV7ayc64B/VkhzeWcn+sErS9ag/YL
dhFmiK8JyGI7RQ90ZRB70kKKcfk2Cd+ihzsWD2SOMG5Mu5AMxFaYr9AjhJmbmuR0
65g6SfAAMnBz9AKFOY0etBRG4jxqUUOA2QOReduOa7kMhd5QnG+U6EOGlKurAI7K
pyR9Aa7CXFNqC4spKtediduv/C9NHJEh4+G/1GjzP/JgOZkboB6WlTP0h1r+BqOg
ENe7lpcpZoDqnjwmnTGlMBBBTPvLaLuIDCd0wqrVl7dnyNODeujn0vAYVSeMbBMO
DInL3sll0kQUSInVDSZqgiurR28ybM5tO3cdUf9xBNeSy3gyt4mOOUMLujt0g+JG
0kMXhTPurz6yvX4a1hICVi+PZ9mbUBPDR07nVsPC8FDR6P1ul5lo0qdGn1ywFkDW
33qjZoAHje2iJOnwgnq7rB+Ow/sXDLjjl55RxSPkaJJUgCQBQcv2UrkdfJYY8TxJ
BR09U7px9egf43ee87PnwrjIq8bgF/mB/3H06PFFkZI6JxZ8Z89dhrr+XfoDQ7+p
/6Ild5O5/f2Pvf4yhQL6j/sILdNtrLnGPKVugf8ZTg0rp5u9Yr1uT2GWhiQGKARo
sT7446nlj9+pLZYu6bhiVzSoo5RWu8NFzIzki+zWHkFIvGgwR0kkO939/rEnkzYR
UbZWLXd1s6ocCIps8pUngjjPIBg7f60O7ZeD+2PYcuhrt2d/tTgDUOquxAZun59L
Wxqo2dA8SRBobuisgiY1UxTCqfMuHl1/l/r7dQ8k3Daq+ds4jwlzj4c+12fhgL35
ql3a/8G20TfbGXPfRTe9ImKKto+CSyoz1Ow3hWH0y7viuUCKGA9XLGWiaWhraNbZ
A3yjyPQrmaU6qmP5G2XSmB8+4cAmVB7hvYKsnAQ1HvJMVFv7ymu2fuCxnWfsPNJs
RewwYcAspw4d1ZyrHjeU1QDzeofIiPRX0WZcpmka3nlBq0eQsL4AtnFcQQasWLhn
ci00Ttui8Hyip2l8EoqE84KB1bSBtwkgSM/0KBFYGiOdUu15MLQlFqh8VyRqWzE5
S3QBFgMMS9Kfs62WgK9lUnkvGGdkkxdMJTmbIvtGU98xfFUMn/58DtZrCiuP/kRS
CTXU/SJXsfZvLFPKoY+AJeD7SWNbUPXiHhto7NA9hgQuK1HcRTiteB3K8HyZxEWq
6XbIZZTOGTYZvOCAtRRwJ6LjQPQTofqmv2MOOXt/rhJX0eMuYgzPhrI+yYGCR+sS
YEwFDN0xHse8jOz2QuDuvA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GHPoRBcm+o7RP4uvTAWHnV78FKR6LIiMLfDp+uILl+x5CTlCgT59L2Khfl7Sz/jJ
1fqinEwCCALII/EQV+0RsspHa0vPDQxdx5DL1VBwx2dNXQ7Zy6Vi0SSYGbpU/mHr
ks3bsPsfZ26YON3fMRrBPK4yAsCV8JN/E4JoZg/nOR8fGeU3L/OsDOEw+wphtl1p
CFhU6enx0pHuervNDp+oNy0m3CWSySoWFFTiodu2WqDUldLXN8n0i2Z/f/cXDclo
/ocslEo2OCqCXmgwiMimVGJG/Ql3qv6SqnI98wYEaJU6BjG21YTehOnQ29R0GpQJ
gJJQ9T3BU1nqIcPrEKasCQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6560 )
`pragma protect data_block
GfJgdt3ZNVoI7Ym0hKSSer31oilMDWwEqdBnvQGDRvIbGePtQeffU6DJFX8V31yV
FDb/9P7Xnsppc4+OtzqGNPUY7ugIAFrOKHtTZJraSfFkGjX9IcJEeHk9l27zvs8S
PkAI1HJAx88nqligX7ZUWzKS7JjpWRKBmRqMSl/8X2ZTICRAM5XCFBCk+u4vFChM
H5XDLJ+Qp2BZJggtXD/csZVFB1IwBJJtwh4o4utlwKtADL1v7y2H/TcXfCm+JSvQ
3QumsleYYGtgmo1CnFuw70Ybyc6ey1l/kG1ECKofFRsA8199Roi348Pf6v+vwrDj
3t6MQJ+B5Zso4dO6Tkq5q4R0P2G0kwFB5Jvu1UA0Li3uOROCOMAUD+Ijis38FeIk
xhN5SBRcTHMhMMpPnEjX276lNQmeHTxP6qlFwmycFi5QpEYPi/Zuzw/fRr8xGBYT
E/eKEibVRH0+UQ+ve6GnEnZlnDK8K2ROwDgwYClwWL4lfhInYvsyHVrGf50CBkGg
ei9kA1N1e43My2HLLxvSxCILmGhGKQskWP3EoRMHeLIcF399r9NUeX3Kl1bSXK1t
mSKaGHB4+5VTf7ZhLJ4/ezU2S1b/Ow6Qe4D856yl8PDBYS6br0oIZrmcKWATBjSD
KDZ10FyBqku12lKrOO5m7GImEZ8HG48N/W9Tn7H/ny4QKvN2mXC2b80KuViYTERY
qKza2mfc0m3jx9MFumq04vA9jqVlOxfBCEtxi25wZhYxUGkziTG1LFoHaTZ9Yrid
A9S8LTMqwMlsPjTIVi6IROHaLEaa2Ga76A5jw7JTnUyq+dd+pne/pH4jgjD6sgft
ljgnc27P+zX5pNUK7S+B/0KQOKz0UsGL3KSNssS3lur/7G+6UzQPAsgbtH5h4GKJ
wkznc/0KbzSlQkVB1MgWVNhZUQzxZ/CBm47EuOzPx8wC15i+xkqLmEoG4PsX1XYF
aBSxioQDZ4h5g0QvQOESmmykz9lpFiKWlar24oJSnhFDYFICRpuY8UqXbG4dK95u
q9AcI9SzduKWimBELxqqN80R/2QKG8TR8mXqEoFp98G/vZ+yU9dfGGMe77ZabCmC
oxay7UzNvlO2ABIqOSd42OJI6oTefs8D1MrZg1VhjtF60455b8czFfNNhfjYg1q7
1ucfDAyus29o8qBBzL/3KP1TqE7vTTLAGZM6WPzF6025YvxNyBDGwZz1bQgGQhVt
RS8Pz5RiA999QXep4djGnTAyfU2UsPJWPOG3Jl1fHbfFXAdG3NAXMngbDOim/9cw
eHojfPy1xFPZKAkqZRfFG85JeQeqnszlWGBJw1TbiUgXysj2UUFoX1i5BJgJOogC
uhITKBAUxEFexbnvU5Fbr6kVj6wg8SAGQ5wM/4JGYlv1EDDi8vu7sewQ660zQki1
hv8JSUAZqEhFb8waNyA1F0N2WdjOzOx9aqeyt9cvDenaIeO5m3c3NvzIDIupxhB3
x3j61o4lyY7q3jbbIGWo1PxAJUYsNTliCgt8T0j4vFIlQqiff4a6+GwKeYFn2pls
0fyMH1PNEeQBqgiqEnvr34mPZyxctAqipZRbyq1Wujv/a7ThPu6t3nKVOUKEdkEH
PvKrHHhEVxOP0+HrflSCSUNYfdVVA5/JeZg5KB4gpod2RiaRwvKP/5RGW+93G6GA
evnW/XCnzCJraXI+0JB6hpQqfh+gPxmbxdClV5U7EhN3ocqwj2JK3w+K3lLO8eDb
kiNLnAlp0PGYMK98MryTmnGUPMLTHOAX06r5QlJHp/xGFCyQMn/SUKsAd77uA+zc
ZVsTMRgwFi598vz+X/Ut8RDml8nYL/r3CCwWaYrS1OyC1Z4mqQk+A4aZj8+Id/uP
FHUMecnNB2I4ZRTwwjyWFc+RX9qOCe0Ly3IKUA2E0qRPx5GgikdRu2QrXneJri6l
yUT816hRduSw6cyXapgC4iw7wyJEPBJyAaDXjVts8hNcfyDtcfjKl/akYGQlMGVo
AiymDmcjDcuzkGVRldOh/6Fu7PXc41NrOAabp44Wk+iSLI00bTCXMOuoGbMdda6+
7qIWG5eZNwv/shaOIyTnG0pd9pe2J22a/5nnNIv50Ci0b0XYk+HEZHGmXzbZYVJx
qkv/umMcmmlfXfe9THYZebkIOiey01cYEfOuuF31+WY1Csj4CONhigwi5aOMzeHR
XSDA5OLOj18arHrkTtgg8kBbY4ZICx+iNTOAUMeHB2e4x+S0tEoEb04wFK259N4h
0z/Kh5ClN1tQ6KD5V2mNF4DkRY0vwRi7CgrzIWgjKUag2PdeP2vWR8ZRxbBzy/mj
CdcwQFbjtLWrEpQqKbRTcVYrDnzRCso/y648jUCpYT2EIb0sWiDzBKX/DfCGa+BI
GQfpH4q98yF2l0NuvoZxxkjEttqw56fJYUyB2tPZFLPXNxdjSF/qpR74lc1RZhEa
CAzfi8eSbCCEkhHxjmk+qOnkSdH/hD2+Dytogm6LNjmfOc1bUGtCN3YsqDyJgBsa
CQS6Pz4WB9BLIg2zwiJ3uXmQ0PXZpZVPGydIz2YPU8aiP3qx+C5Jr15dBjkdR4e4
ncMYSGZ9kznCRij02TiiGvaO8dV2nDlY2GR3o4LaSfcabAyCucfOOX0NLW3pldo4
OEB1gn9gcVxmEEIW7fkr7HYLO8p0NEHy6V7CmYwaHKQIfEx/D3QR8bBysVmAyar/
3Qx2RDxvFLebRcCdO0BTZI55YLmA/Nvh01X909qUytbqfSIoPjmkCWG+mXlAk/B4
plP6QAsWaDhPIKg3QGFeYLf4KdxAni/QO9t7/lOsq+VdH6ZNhFK2NSCHYno5ibAg
cZKSOXyX/kiz4obXjmIDwzsFM3K/p5D7B5x0UZRkFMprgMZNO7AG4HoSphxkZjED
3zc9PtrV2EAbqYNI3lkDeKFYldxu+LIbd96/ZMKxQX3sULxtTH5vz7/cn5yMm0ET
ofSQ3w0EX6nAWa3694kVj1oUfIDjKJnOyVOjBItV9bT8lyMmRH32BcSYsGCGtLXs
uOuMnMM4YDgiuI32cD6NOJcchPHoAZoGUhhZ5fs+Rg9GCde3GXvkPkvzYQiDoFE5
HTrBdglVkAI2hjM41w6LrQzgVmCQl2w7yh4+31E9ML8iD8mwtklUnU83ENiZ28Hw
beoCSUR56kfGFoKsF6rgNK3qLlXpYOb6NtKTrpUJTQdhZimuSIU3UmNGRxYLpg3b
KLFxyjWx0lgGa2hcbvYzcfOoi+RpeMcuLHvcXlbmXZ14RIBPxYjwWkuQgSVSq1Sh
YJygSlIbfyC91nisk2gURjgyNWE3K2rjJzMAJdYb8fpi8SWbd6NuR/k1UoZCGvbS
mk1ur+jEz6sWxdTAWPt4/ZFyxt7oL5mftRXsu83Qgh8RJL45KxfsqlyUphGzXFNi
Ky1TV2lqPbEqzNMVR72h32K80JfqhJ7h104+YQ6ezoKfOplMUcm+sNRb+iVzwVgA
N9lsmCZk216+AlVq4xdp6tAqyiMTd8gZFPeGPCy2oqWNNRvzKlR0w2NfVj0G07rS
m04s4pJ3mg6sIXGBgBaioTqLgL/TFqE1VunrcTToHY6GuNIgnddeVHxWa9U1dRNH
PtPLgx91Gt+pFVVovbyzus7CBzkEd4y3H/LCN3XVqg46fJ9Dy7Rnv5LZf+JUdxww
0FDC9K3GZheOMOK4CIay5op/itsKk0DHXTVBWSamtBL/WKWVL0M3sxmHc/N6c4Ie
jUVoHU3bLtx3HA4/raoV4ZEdA9+Es+4xIAERuVyFFJxssFslJdB8VgtFIfAgoiIA
okI4qJOrk502feJuX25+6oIABcuJckktfyKuAWGacFJlLfxWUc81WZ081nEjlYPB
g4h2bn0tHrvWd7n62IazaP2yXOEfXkw+8VS+f8jDh4BaZ5mxug3q0wxhV1fGTJwt
E0B9V44uU7G8i+DI/HADuJw9nj4syIZDukZyTgH+EkTIYKeNjoBD/vyYVG5xkJ/1
0ZcZ93kjiCqmM9MjDaCClkABCPSLF2LO1pW5oEkIlTTX4XMlYqJ8PFH14OtVnAB3
i5RyWKsqhQ9VuEwkuhmRoPFhtdo85zUjxOIgqs2KFjBRO1kPF53a6EoVMSx6sFNB
w1lqD1fFaBGZ6a77w3O0rF2CAduieniXEQbzTdvvlMkG2jMHOTBS40C9nlLFW5LZ
J4lF9aTZmwOmRnUFfYXgEkNZnWtK+Q792f4u78pHsSB3CQJaXUu96hsTzwqXWntt
gXneTTL2viJzOKalmcpZtn1qbCI5q94Pjro/SmxBh9OGHdFy8dyAqdgfw/C8JrC+
cPigVrIoy9coTKonAH2soGx3Y1RJhOpENTBpXbI/GjehGoAX2Mp3+uK3BSwijmZD
RoBX6IUnKCrk9KyTE+FZpFmoDl45XGDV2lw0Kb8zqv6QVpNvPrp+oQ48KnLnoky+
vO+ftOf80rRKm8bT2ztHtgLdo/PZVtIYWvMa1J1i0gltj8zBbEzETSKvHNCLOSN+
YLlB7p5tTT46G5xrii9FepSTGBIu8SEme0u4/lmYTIocj6OeUV1fqsXdk5rq0Y6h
xyFUJS1Uecus/QkXAujJxIZp8JfTb7tbTjjnQwUdAxBfkZRlPD4z2F8mMcA2QO12
pLtqWy3ig6TcsGKRTsHnZbBpOj4rsGvzeRXUUv8aVcF9UyxbzqqPCbqoXTyuagNi
7KED+6Ky3BCqf/8kzyA22WJ8oALS3pPSEguSpV4vFtNZqXGjrhPZEKKTO+yH7jDv
PCHgXnj2aSoOrcdJ0CmaaRu7yndxQqsCDgT8M7n9LW3xA3Q5pW1sXdkMndtV2/R/
QU/3NgXkgd0D4icvE7ZsLANnV080HVH1H5Q+tU3t85mIOga/BV8Jst77LEjk/TmE
l0rEbbDw7jZ4/dmbmpTxP1fA+DjtioGbbdfwX6Jm5t61vizdoEQX4Jlf8y7nOqEt
7//glkO+LlTafqqg4CRdRysEugYpV5tyLU97AcjmAoipDwlgXbMXs7V63BrKuMRr
WGuHg8B3SjP1UlhPstRaBmHsKnUt7jMCR/ogUKoKGnz53FGJYmc0cL6ZtFg0GZo1
TEh8yleX8gpbghk9rs2o3LCGAPZag++KL1bhVzEFVDf72HtPTXMH5Vpxk0U4Z5kr
fAOnS7tq1fccRXBDcseHonM6/Jtqn55YWhMWum3I6RE8jyEKo036wwhLrluyavz5
VO8yaDf6YEWdnKK4wAM0UTkHwgF7cvL0tljGFYBFStXbs9r5SUtZ5oy9dYDSZFdq
0tbPZt+ayhLCzQhPGRRLP5Wlp5PIKJL6CCTf9S6Zml4mI91wwfddeekq2ZM1JGZn
hPyQOhYczhYpEIjGIlozulrre0iCdw3lTpuRFwOLo8NQD7BUobAGJYIRyeXuk+Va
XxOV8IhezFTuOaBUSmZeIBVX6DGaIqbI34y5bfASOK7BkUfemDZIrQMPxYxj8tXY
dt4+36hSoX4gQYR34Q6Ko63BYkEqWQK5VnuvqXTnWebuxcNcLZn6BT70k+I7xLxk
LwpD4ffpbKKP3vhnIFvJBya0wryKu5pUbdY6OMvm0pupi/y8vCZslFoxf/F0Vg3F
BORPxWl0F5yg/Y2Qz6LmveBJqBjVrnAN579Kqqg1uD1AaTxOj2RLyi/olg18TPFv
CQzFqJrHrahZKrJf+xaCOqKopwcyNrtN5ce7pEk9wZKp3ZbLs9HN0Myqh1BcaNJl
xu9l/d76SsOMbmWbVa/LYll1Iy2fTFOCXMWthOPjAJcpjaE8O1ahjmsbf7FaDHz8
EEFkT3ezsT4cP+cuTRT/5JJhB/V4yRcXKzxcBeB2qdddfDa+XEUAuCy498bSC43z
YU86C65vARmqmqpkire3edyCk46/1cxouRJt95i5kfzTAxQT/kg4Uzm57x3lQF2Z
IRKA/u0A7PCc7P7Qr5Xys7I85t4bugrAbmV/NN/Jt+OXfE7HrCitEr4M5OkKMCpf
LT0Fp2wmaqNe2f51rF+sJ/jcOfmlcfUUlZ8Bzt06hCVgN8OuPcRXbHY4HM7pla+1
ikgWukaaVVWX2JyjtVVlVAmLtyr4t26lqW1OOPlCKRNLXH544RHZt5AiD0Ha6OaS
jPj+pEuRsiq1ctwi2Y+xkhbCfyea2C15sJj9WHxGVAuSrniZ9wVVuIhursg4yOMS
rCQPoCdurCYgvirYo9CWNKJIN9f604qfU7OYS5YbBXNY/Qd8V7snzATCZ1uhtctO
gYWoMv+bf+pOvVRRoPwDnywrBIcxnGFBXoWc6HtQ9kwO1rIP7H+SRQQ++hHhLawo
nhYvf0VGoYDzDb/YpyUIax2yrsAINh6OnQJU7lwHvfKHU0AJ09o0WbMNRiyK48gZ
5PAJLNJvM0ikvt41umPAEa9TyAIV8pY7faaWhhq/MnxSruFtHzH0P3d/SQWXSE4x
qRahRJbB772kSo5n3jRTP90+RJyY02rIxc/xUIpcMWdHKdEuBwF1LOfEiHfUTKaS
Jm+ZoZSdrZZyDKcfaJk1XTmOkrG5ELGdPkNHtr8D0dZEuNurVDeTiD/cTjzpEJ1i
MI6dC7GcY6f1VFm88AHOiISwOGGp0IMKK3imHlA30ZmoVlO/4UP30aXbBYyugimn
4IDuAexCQzKfTgguoVl90dBF6QJOgmqYvCfPB5i43y+53z1jRzT4HmwxzzZXMDJo
SK2+iWz7S9LP1yn1CQuf7RcrkbOVDWBqHHrZvNZ4G4hJ0IHvRaW732lkty5DHFjn
Qx/XRTo9U1D4Y4txWmzVJW/nuc52WdLwdP9OrMrDTdSJVbxyHxGNE72SL87pvGa4
R47MQWEjJegtYyHJcCpAZ+p3vCMSfIestEvYQEpytRaqK6KU/exhX2NIgQiTKR6w
1lhXBBKBR+r2eglhg2HSQe9QDmhIep9JUPvNBk6vAdnfRgyG9dRmghEztNmDWnT8
iXGpVbcAcT/ZzkNPEo6piaRrWMnNsEAiMWRodnPeEXWrUSy82sZ+UqAZcqbaIp7o
Xyg0w6oIKthOGttokoAIVqlKLxviCruZhwAgnrBhBmurzyAgCsgCHcpFGSyED9Ys
8czMw5IKbQ4K2OvvBCLtCVwgnfAQsgiXoMU286IRsPOh3ZfV/58EZ6MUG7uGWvQB
ZxkJHPLNDroZbaQXp6pJ2blSq3w1hvDhmk5obFOjnpUyM4BWbwRse4qhwUSQSh7P
8/KNZ+HLyhxPbaoB9FuDAaWxcnUT3UApZW3gUrRoKdyIqYGM+D6gAB6Wmw1eaqm4
vRu4BJWMfnOL9tCdgoTFDy3ibPYqPWFl6IswrF+AUeairwfJA8lWM36YCCkW3JGB
Tt8v0LpuwoXGwW792a5FwtKS+MtmfrsfiZ7DiIldydM0U88xzSsQvW5UbxjIWz/F
wPG8ftfvQ0wd7rYTHdxzyyZd0fMS9acYomL5VBiGGnuhN4pJza3bPH57cEsv40Ge
5UNoQ3xVflfY+UEgvdsyCjgAXCComjsjnteklWHDvl0iRlk1eEg7kXO3p4Okl/8r
tXzi/BkXe4WGnwDJjb2pD+QwxYgLy1QC1ryx0m1UvMENiAe+QL8215Lgt5d1HORb
/CwmeuP86hqtqwNxcDcRQ70ym5M25ygP1qAsCQvjjgKm4kLPvX3bslIr//WRafks
i5T8LuT6bn6hwOujwUGLJeX8Ev6pT0MiCSgGShND1+skl39F0XEVC0avlwH0HHiT
yMQaLn4GvdhgK68vLUrukvDnNFVSjGSBkJpO5RonPCxp+YtTWObxkL1tk3+8np7m
tMQ9mP0X5nes0QN6+4POD9pb+T4HNTU19zGGhfOpGd9QfMav1v0/Qr2+v3PjwJec
ZL001y7Psg0lx5xmiyiMfrKGjaE1L5OlCiwosUdLTe3a7m0oHILutGaqQJxSADjD
hMWAgoxGhR8gqCTTQDOAzo+baz8oVPUWJJE+yffnQKt41zWqZn97cXO5NRSvnmi2
oLWVcrAUW8jSrzaIo/o9VGHmCYq/YYYXw6tIjR1CoAwnxvR//10FSAqhUN0LKC9M
PsNwnH2OZwCOYW5JK/WZQnngmRfChrGx9kWQqOo/dPAQ8mYkI0rMY53CamnIhrUl
665e5hyBJ8mScJCRptZCFX3Ye82b169Dv6ksKq/qj9mJYzMW3qfaQeDpm3s+dvuL
7fPRB3m1CieEXuLEV4LjMTn3K8FvpQ7AgIYfxgiv4EYFKh2tuaxx/yXJp9Kw+qiv
HlFTODs1F+mLO4ftvMsXDOpVKMO2XUoFXAxo5ZRMyGBBUULo5HFPJC4KZe6OqtxN
JqPnGpn97HMtFwBfC1X3N1s8VTGrPpSpgGzxHjqEZAbSrN4FX8DYtbKg6DK9oGPv
B6MVe1y/4TPUi+ar0HXJxGUU3SV/wQBOplym2zbY0DooVGnZnFp+sAqtsFElnMpx
cKaQKU4x02haN2yYJk9J/F4anMyxjBjC8pw+ZsQQokPPzVIQWeYF4xMuT+L4YxeD
HRvdZVAVo++/3v/4HAiOcIdu/5rOJiVtOTLZ1OY//stdVp3k0AMJSA/nqBmhIXea
XVbblSAyceoe1qoawtCmHlVK6yP70GEMT8rh7szlPrLs4yablq8uoKuMSJok5Anz
mhkvPpFUaMeAcJsO5H3I8vewD9WWTLrKpQKhcAIazF5V63e5jX3s3TIm8H/sDi9w
MLADWcP8GQj7UCignW0UxubY9Y//Hda6N1KQuESV1ukgCuHpD65DMhaSrk2xuiVs
8K7+8Y4w44XsaBITt78aryxzIuhWhRSvgGq3Ly061jU=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dC/IYl7vJQyxY3cKxPMX9fk7pxJBTzmTFuAVVkQktRE4VjX/MOYjnuT8N5T5wg69
9QlUBBUqLzLvn3VeZr6tmaoIlgx8mNJNpBgFqXIemsrRQ0rwB6MdgHjB1NjzRLfM
jUrMrKvszBJezyxiC5o3CZTJD3Iqlb6q+NpXRyHaTwJUNHNlNcjb6+WblfDx1xqu
+ForSf1J7s4BuwF9K6OhAht13EJ33PVsdKafLzhzdKvtdZQSRU5w5+j8qu24yfYr
b3+O6z+lVupuA+MUZMrY9JijK+v8Qfx5D2BrgO/SnzrkMbU44rFwVCodZuRkshQf
BcL8+LWHkWrfhsOeBTpEkg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8928 )
`pragma protect data_block
hYa1IujABY1wQjGruxUHPhZmfD538Ox1bSzBZP4CWrcb1j+XUazDZeSv4GtX15Bo
Rx4JFlyB3yRfkWlEvuNrIX5y6tnaY9/3SBAH9ddFKDElLmcZDntZ/XAYSJePcqm6
pbjkOEi8BkpWdKzCVs+PhRtHvB6qrG7tnIdnvGVoPKBJIUuFgmgmALN36Gh2TyDt
uF5b+IwIBaqLQREl7Et2Q+uMh8VJwwoZO25nuTA7lrdjWzzvc8ThJZhDRzHEFGpS
+er7KGkiHsSWOV2zoZndO2tu27qnbIPG2bc19dbrgCmDEVdphh8xTLCU9E1scJuR
sYCEd2x7LRZq/+s8pp9DaRCAt0gKXc44Qvamz+MeWtWvKCTicQOP2wMeTGhKxNzk
EuNLENFBwAVYxTH4oKEx1n1i5sbYuLdRWHBAFJoi505WxxCK/BePoJ3EmU5RQG9h
pnYMj0jKli7NlDBaHmYszJNXcvN0a0xlEQxLyB5WfjcATzIM+9oG9uGCnrbvGL0S
C9rrsuSoUOSQj9mWrxIIMyvympyrQKKYVtNJ3qjfIJwmGfPBPb/VzzTal6fipuZP
cfcVsMfZ8kr6+7vXW2R4qWkVN1YrhXQuNNwCalZylO5YMLhFoo1gaBCD7pqwVWZm
qm4E9VUZBSk6pj6r3K9ZVdKXO+zBmbpk5DTbBhledatppBU/fUhlTlGcnWnBqAX3
h/lZY6gxSWpP4RHkLYOHtHpwYmrN1JWsPsMtDM5XRG2wiFJ+Z11X3o8J/S9clX0K
lRsUPe7EdMMpfrnm62Eth9B1pHIutTONgVEeMrrcCSYc4tViNvRetQzetSHTvwki
KOJWA1UZRpMPXxTKYU5JyVvnuuH4642Z0dCY75tieZ6f5EYILCJvo0JaugAqWIg3
eazA3COpzSh2ut+dCPXUZWEcnSs03XQvfVV0tViqrBqgafWCaIrbrD/LGZ6JGzwA
GBxGJD0XWFCfmsSa/Ojdc/52fXYNAS4s3LTzelJL9aBykF9sITJAE4HswQBMDsVa
zqaitVNYOMiV2hua+m6AHcY4QG3Tumt+0gYrd10ProTzpP6VwWVg7hj1+nf9aeu1
HpA1+279ANpLubQajUUFAgijRYzOQx5pxjAQrQwUAhVgUO86uXvUw1ZA1kGVsmST
R2lWuUY7ouvSDn0YvsYLZsDhjghdOEwqm0E2IHRJnhe5qJwf4byoXMx7Kp6BM2MB
XZK54GEtvqSVbBEUaHDeaMWsB/SJs5kbpNyFmlm83Yc0sKnAYbnNW+INcEtqtWYr
RTDES6Yn7ugsKEiP6OBBgxaLqP+eDk/M9vd45mJ+j5wcYzy56J16Q5ySztcPhuKK
vjNp8+iJGPj7uY8lJL2D0QkZKws1c6Xvn0e6s1KFd7LWdcbmk/lrXDsUhtlDuelP
UYDl8s1rGj7UWuXy3jk/eIbB70fGNxv67bzXW24FGKB1AVqrhrSgoIAYkqUFrutr
efDofAeK0Z1NmrwCklxPxkZ0EsPQiCoEZEKUL2OH9fXZpX6w0F34sWf4WCSf/sAh
kVXk5O/nMPmgC4iNLKIcE3eLYahNita7WXqqN9xwsMuLNBdnrtTcJMzxm54KSLlq
r50DT0eIqEex4lX0AtdV1BuK4vEmRKgIXkrrUp4rz6iU/lDw4gm6v2JrQVVM3WZ6
v1bjJIYFnVRtPIlyscQe07qe0aX/hXeWmzsAs9ztcMbSl9hdyZtGy6R8gd0R/sIA
bPhaTW9/zCayQo+FV69xfnMTO56Ao32RIieLxBP2idUirNgKnpbPQIbH/sYf8UE+
xBPDuS9wl7izaC5wBmjUC89B8AlJjIDjYTUJ1B80iQJcnWcYfbC4t945ueZ6tlYA
iZoPUECQR0eg2EVveRspHMpbJpuKFjCjLRC6jIKIXqSOS8ykrMwab/zqDzC6BD8/
FCHY9HaehCHQ+ma1hDzvrLoS9mKBmG3JoBSOdZjIisr744+5pkgQ5MP1ZfONmA5M
l5hg0Fg5zMKOkhnUZ1gMlIHGHo0ubdqISe/An8qXvi4sOaUEWsDChqD1SKvs7FqL
YmcAsNfF5xvOPYZTAbnA2r8xvPxIbCQfSzfOPXqxbIKlroXPzqcpMu9lbh9T0Knf
1GXdZdRWvz/dvMM+ei4nQx6AwtGC1BncxC4sCUq4kWWwgbkURJqfu+mCGh2HpqOx
YaFiKOPVtZP3l6t9XSKBRmHwFNmHTcFWNtF3CUL6WGaSY/PkBb1WyhzbQICD1vx1
smQ3sWM+RxnhnSyW3QRW4QCinNDlQ/yzyZK82DoqpMzW4cjRxAzTWo2TKYxKvNf3
cvD7WVgG0PWbSN+yYva2D7R1Z+WgwQ7mVDQ7AYrFZMqOyDEAguOUq2jzkpXjgUU3
OsnRP2pYzSpkbDiHtgArQpbmMXbpeFR4ESagqzxW2me263oSMLv7JPhO7or9c9Tc
WkDPbYOFROQsxDaFFABiFz7BB9CeWDqn+EPHBiLJdpIXIjhQeWAm9QpK3YbgYaya
k6hThWNrUz0q1JxyqBDP/LhNoMBd6hLmtqzU3cDbRUZBOeMOFdsXewxXmEgD3YBN
7QY78aq9TQd1aQUFv5GlpJWV1XGCrUmxtkxVvEr7EoPP1ypIuzmzh9MrDiqBZTCQ
KoGwQXnVPr6fFhKPY7RPDKsFPyu8k5dP/Yw+SwVmhQlkrebzZJvmwpsmu15oqxHL
GkrEvxTem2B+vt5LHK45HsPBaobHkS+93SpxFGbtYYoPfQdKckpyvr2AzjbqWMEQ
Vrv/QtyvFcsDyz6a4jpQdH0oUO061rM7R4+LXccQEfvVcL6ahORnNG1BWMzrs+iF
nt1OwMrSguEA8Kebp9faS5k91ZxjF1kyYpIMpdcVc3dNT3WR54VNpOu4iX+PjRFP
pr0BIiYEdaYJIZpb4GkzCl4OhHUeBMqbZWYYgUf/mXHjDVAsO7amikL5mH5rhMT4
CYBgd6W991hB4vjtMuIC2U2ZlD7gRHLniC/PGfBhRb97XqntILMIki8XTZSey8DW
fxwGHhAQX6D59rklmEZtjYLOjYUE5CBuzgLmcEKS0tB/byMqUa/lvL8BtepALL7H
s7s2gmoBcb9O3JCYN029IcePTcAols4Jvk+S8m60fWG/rFJt6jd2lB4CcGB2qY2k
5ZUPnvDy0fwoWORxcZ2VdoRqURA8o5gljWDDOwHbUj3Au/wHhTMhigwGjF2dgCoL
0kjsbSMc13/b7DNycHQsKB8siR5xjuJaF+VFEhBTt7YPvtej/rQGBoDJfE24MiHP
YHjMN+U8ymRlPy/GJf/6/v5hYg5GCWxvSaRi2wkCdzgRi29CkjzyiUJv14SvRzoc
RjG/cZMcrTENmaWIzLzrTuybdyrIU16SyoTWXv4bZc9QR5DOFPxD9+isznMlgOEq
mZzs5da8LS/VdYNuvu1Xew6iKoaNXWUiucRG+1h3PKucB6sXJE6VHVTW9cs3VjkD
sAtcr0WD0GbqG0qWl50FL9XAOn61ToqzrbGJFD5W3v2kFzF3KAvrtPZE8KlUX0MK
b8BCaHnTWiWstYbaelsiKTPpJ+GQePMwytG3gGsoUCJDMaK+ny7OSH+X0tNZgYI/
4FtFp6GLRL+DK8Ca1QI3i/m8PNz5qjKZwweFXoyNG3wffjUQsJmPovWfOjmii1Ni
9cxpD7xtRDj31rVzFJPHDn2ERC6gdlwnhER/f7QdoHlSpfQpdyfkAVdsZ5Ryt12X
9J603cgngdGrL6aCFqbUqjO1XrjmPuZY3iXPdEQqcxNvej4NJQpwKXoTPlObwaS1
frQ93F7UA/UK2pFOF0V6/6XX5cuCIPs+GPM2uYQvfP9t+fLAcrIGxikc6KDacRnT
+rs43kdiQUAolAiaL7e0/sckddDzOyKlO/tYOPuK19X1su98Wqh7o8UVVmqzcQ0R
Q1rV4M4Bnu4rtWiy4vCde7jzpjJmX6lD4mZlw0JUttHJgsYnXUDXONv2epAYpJHT
kUPo/+6ZfsBlAVDjDCiDYuCLS+aH1v3c8RlTspWpvZpNdKtCvDQvHbY/7xHNifOQ
dsqJDsxwLfiWUbvpv8lwwzi5gC2lMqx5IdH3XZMxYuMvi23+qGsFOphB0wQs2z3y
ZXB1Rdr91Te8oo9No5ORJeGSSvoaoEZTxYdXUE+zVwxV67blkrbI01bikzd6Cxh/
bu6xdJqTYe5TarewYeY4zrhmXDepLSq7Vjabnx/FlUPs53RcPQcoBdJEfkIAdhyp
JSgEfAoz1briohRBxkigUyLlD/FL8VwacIrAsRUVk+CTr7eC0xUl6mOu03qxAyj2
uSvd90e9bVT/JOkWx1ionj2YZTuUOtgCWvGeUz3XVjw/YDT+K/clrOU62mDKkwIz
hKhMvp2PyMIuzYVcf7JYM8qibt6Nj5QCOwnZqOYCkktegmLc38aHyXH3EVfeMGnC
g1YQStAGe/V6faZibORj9BK/0Z3FznZl1r4PwISdYz+Xb3lNeTHOL10aqBrcMovc
uy7SngZb6D7MjV7t19OlolcBRJ67YXpzGH9affiyQq2h7462JxgWalM9yiuoLCl8
YjwkAnWp2jopUP1xZpPFVlEoJtKYuYs2SAtP0hfNXT+817dl7YYztPrXKDTrKq4n
feQ3/NDd76FppK62egdRIERPwuDJ6OhijaE8QDmaL9o6f74IJPQv/yCBsgmwt2pg
saVUtPsNQpBpT3I5k5dllXKzeI+WZrT/plSnl4X0juPfCLcjyaQopUK615MvVAXl
+YqfWHFulKLQoIWL8rpkeYLZTOdv0vbZHOM/OO9oImyLg8cs9pbIhJG2GbsVxtPR
X0yH6vsxY6g89zNmT8/ukrZBOgU8MRYEYBDSxU3sM8wjUwNnPV1nq5/gf/KJve20
dQrrgf5slmklc4zSDHZblbeyUHj2Q3CJRnMw1YrdSKeTn4iQN2Bw2lApzrUaVZ9m
/7FkHTAYcoyGqeCqIkBUsfGDN9nOOldRvopeCqeGIAzMu0CLZXIq7+2CCs9UiIQX
b3PgXue2psww1GFWTRDhFp/yn0i5ZQ9gaYtDZOdy1tqIbdtQF0vHFEIp0NmxaLEg
WFTQnUYvN1c0y8kNoMKPbuumSvdK1ZsWjhQnfWqmH3eDRp/Es1lZHMZTcb8lU2Q+
u3MZBKO4MFD2hYFxLDDyJfukJvpLr77UsQcS6KNQewLqSl3Bi4+iKGtyw26+mQuA
fJ6gAk9iaszmEGaXDp3pUFnAMYc90MLaqiNz0fL6QC8rYktqLEWTnKSSX+8zAYeP
egkRbvcBhYJ9R5VrTXNdsggI/OYQKdmyqQzv4nqO+V6+wJbRnvJBgTPFjB5Eoeo5
BpAdV4r1rgnXLREexUnMrqm7Ys4JJDSueldNCjX9Cjf3BaDBVGrXYIPp//W/XjVQ
3Tf1Rn/QXXgP509F1SpxsifrR3HrBbAf5+iCPi3I5zlFtEj+eUJIwjNboscyMLEr
a9IwTrO3xaCkYJWyvBt+DGCl33ewmlQlCRDvOJCOBPAz7i3LqjuoItj7RYdgT8Jt
Wxu9W9xatyR2Wk+Mgw5/vl6mj5JbRhAqSJdcicesk22r7Idflzc99RMT21yEUoi6
Amh73QjMTSTiHetTMuJPBFphyzusVmF0+J0AGrHSd9zvYnR1wAhSoHvFO9aR/omi
/FWB9lQ2d8tF82LnX8xFytItZZIJOBQt2x4Z+UoaRJgXhy9+ULtqD79DWpaN8pOY
t1Lu98+LE+aAo7vgdL3mBOi6oOOOCb1DblgJWiQMTIBeN4x+R+uDz9kCudX3sLA/
iaLKIv5597WOmMm0Ql85OGGUCJ9Lv0eoqBKusjxXBY9l2363ukRzPTCBjhHe9wEL
qOOCi9ry2++wAL1HBACzUm+SV/dvy8Zb7Rknz04KJmfKgtG1O6xymQ0ckgCQ657g
hXBwWf4yXXOD2ttpj/tBHh5n4imJhpCE5xkqGTwMOUXRejUmtK28yPUe4sVMQ7vx
loiPuZgKgewk43g3f4OMjsHirIinAsZhPuX0pyMA8+EBpWokcKM50PhLJv4inb8I
hKg4cqnYaxT0evvxdkvrBPWq7JlYka2wo02CW0ikuB76Yd339D/EpMc/zIfeLPXC
9CbHTpkls1BGqcjvOm3jsZ4PgONjcZkpi4aI7RDntH1ivy8Jm+3K/T2BOY16uA3b
E99XQLDQKiXh60AjPxd0dCfmvnLuAGvb72nbtKv7ELo/V3ciNP9mjgJOg8nUeKZW
+DhcZrR3B7ZCg8dVICVWIaQr/mJYxma87HeujsG4b0+jfkXfDrf1MBtqZkeL3zt7
rcGyiheh4aa63T5WF2Z9G8SkcPNQDdrDbkc9tS5pCFfTP9YFaaDitM1ZqOtne1ld
A0OpkTtnKj79tIcNIDJfwwxwgDNFvsjtkAqaCSP1+aC7EZleVcSJqER9JDCssH4n
McRkxdopTgG/jiJN9GnguYipJo1LBjYkSX3KV0u6zGnOSukSgEgdKeBJ7h4B9DHd
eCkBfQVwtrYgCh1Qa/U7buzbZeR/45klkS7Y9HzSZ0Q5TuH/rkLQS73EBXWBWu+/
DTlL6ZMm3WDubR7tKM8m/vFLjmtOhn6BkHL+wB4/FwLPikteR4IyBpI0of24xy4K
WDqiBkujqihHU7GKKs9gKQ6P0t/jY+a47rKi8ZFEoJ/4oe4oGkjjltA8d/wUtdR7
EoWz9gTmBW8e+mIG9aWXCquLtGh7ZROM1WbPtzVMldfEr4RJo68hgVtDXF9r9fil
ELn9n+b6ctQlpISCpxIgWu9nM5VTlvrfJbQiZbXcDNtdR+4e4AB1gWrVz6xkPxv/
rFrT9/bfpAarq/Swfcu2XBcENlisivXYTsa5pcoiQDeCX6+JCX6BQ2dDl8+3hodF
WM42QFBUaBE9K0X9GkoMouM1M0WnXroxf/5t0NxeHSABDLgfaAeHB5fnATGwO+It
QGoqVSvdcnXUWH0vJtfvIozJxG7MPiTEd7gGMsfAWze91JBsn6crvQT9YIp1lNSN
S+n0BOSppSDg8bKGUG7RRyKifWM6ZlfEI/srrODsWvKnqa2MOuC8y7g5EIh+vLXx
oMWV+6knCStP9jF2TESG3h37qntvAFmUZyCRl7subjWsp5l0HIrogjkXQk01F/BT
e2lKl24zsr7vhDYNU84fN/aF/dA76C03ATtmFv5qQqUX/ZoQ99eLwx3tCvSdpMRH
3i8p7KHzNphxWpyy58bVaEQ+GlvNn8fl+/MaD68r8P+cPoL+Mws2pB4WlmyaBhN7
WnGXKwdS4dNSMzUlTi0ODpn2Cj/pfhvS2OUuhU3iiC0f4koLuBekBfcS5Qf337Je
0qHd3r/61Pj0rANG96Uq8nPMzy4TQ5jQUs2JIZpKUNM15O9cZSCTKnf/aUAZzFtb
6wu/8ikf7nneRaohmEH9xnA541i1T+pKaeramtalZeEN7vHs+zFG0wr+grVVhjpY
tm41aIKpGkPgPavEHe1ah4ewKqEZRmsyO2iKwRitqWh8glSYVpP5UqXfb7ireWXV
6W51o2C6vP4p7uUVnjvUBExl7LycK262JLrqhUXd511ifNAWY2TLEUiB4hrCS6MD
m1rlXzJpaTHLdLGdzar0CJ9zpWdqhSAgQX/Cl8yfcf/v09dY1oSoXgxbzfqzUwp9
i8bICqjq5NcELOjncaEfeC/kq4XVAow9FMSkA0+Ww0f1LqQrxB6ycbMwGxrcRN++
wdYp68dRtG+HGiuEnkjXii7J2iGLFdTmPPc+nOHPLPJsWfk40T6kFP5yStZ/S8/z
+EFsrCr9uaIDsWX0CESyH7RINz4ylP8Dab/J6Owv2IwOtpray7g3KlZVE0SvYTCp
iX/7Z1GBQs+3GX4X7ERjXrIJrGV6ey+OYHP5seaSxdbdj7AbFUPe2lDK4W8udMDG
E/hDedclMsazBiDF6IzEHKb4zvj1kWJM+IqFLaPFc5gSdoz4akY5Lm0lR2/y/fNn
q9Qjx9ffD2MRPNPqAotsVkfQS+IirPxojrt+ZR2U1UDLlSmQsvjXfHGfSRKuZSDb
aw98UOC1ZvhfwHBq6lm/f5JIrtFhA3DPeokjRBDLLICRd3hKjKrJharUPB+83Gc8
ZATEwOde7BviDyBhH7t8xljEdZgypShYiJsXxJ2ewYwSvnMP21hMR2f4d/cGAt3L
vb269yk8nZOPxO9w4kvuPLehYJDkmcy1GrzoV1Tu49/zs0Pc2sbyc2DnrjDQ18ej
XvLzzPnyo5zIV5Sd/w3WsMWFcMdYU9sRJLhxNQbLUhXug9t+/oSooO0WsG/+DcTB
x0cTI8WF/SF5H0zNoXVQqf3lCkIxtJl+RLhs8Jc5cNB36/TyQ9Rl7Rfht1g9hGiX
8332OX4jo9lyiyts67BU8LN2IX2runRSaLoXmFCoHPdQu5Gu3UCl5kd4fIjj6Ayj
wqcU0qfGUDSHGFiy58GaOqkUwpYkiELcTGtKrz/9Y3njfOrX3CbIHE4ZIQ6a0Adb
8bQsiiprDrKAWuY6hxm1zn+qNH9Go7K4qu0gNgvwgn5S4p0I2dhpSC2DPRwpHD+/
GdsO6klruEmxpaKxz1mRkLJhNKefeme7K+cbS4EndDect05tl4xmTCFDm5JkZ3Al
VKQNqRaZnMBa04NCo+46Dzn5nucjx0xG9+xeHUP6ZoDXDP173482x9fbfEOU8Q5n
lrjO7cpfJBOt0nwqXZNUfhEN4xjgHLV/9x0X9+fLyF0gCBdhUlNrs4JCBebR/K29
18ndMatIdIpGUuiS9b4rb/yGEI3oqkh88paokQglCeTqMxBWufBW81XMqXz0CpqS
Gvjg4JsbiUT89GwA55IYImKSil3Gl14zbg/+q0SCIoEXuELUj9t1pZoKrb02zby4
hrKaSc54SY2ojoAynFTW77UKJHtfdKPmxOZfLgBpRAUBU+o10aG4aiiH/DQX0hL0
EIB0jnQwfFVDtsFcdP6c+O3qi2510ubntM2kYgFSEi7+mSachfuYQiEXKWkv9S8D
WC+rriM0mUPwVkiozpr0ihhl2XrTTm2IzcqAjqzwWHmtOdEql72CjzT8mfO99PX/
bN512bHViDQutZYwvleb79EQsgHWpkO9t4ygPIn8jbtksise8RQacFw+sxNG6Uql
UBacujsX9Q7yS1875Hv/mAphzbvmOpe2GXRL7DmeUKOieoxJZiaOWFtilU056nWS
C/9W3X4J9xzPhebEcS2LH3TFtSsUUfQ/O+d6ycPmYJgnzqbQIUVj5VKlOCyz7Nzl
7k480Hlw5L8Knze48pQjXvVYHBQ7W5IP7AyV8k7f/KdUfAq/ARCGcGeHDK04kN2b
gcqh/eJPvnvdY0kj6oSLwDlxjBmAcZLTL8iCOEEc+lZCb8zSdARSdhoswoejMIj6
KQt/yjkvFslNH9jVWeKclstnFGdJ8hm1YFvhU5KoMcxAyxzk2wWGOSDP/ClpMUbL
MdfzpxF9jy3OU90vlxiYuBE9lechthoqyTi8tgYZMi50qhQ4tIVMyLfaORLlg96p
pvRtfcUv0YHoiN3UBmcfiNH1Wt3KosvF6oUOqRJRC32I0PDF8Rvt8VyPAUOHiZNZ
fkxz6ph07mNOsUtZvk7mJQJIKBFFJr2kjl1Brsb3iKnKS3y+hX6QyqMvTccmOOiL
cjcqSPaPiU4NDQOl67ddEvuGD0QnY2D6BUrWGjEaB/rEhOziEk5Zjb/IMnyFL7gn
JlWitW2zILNvwuk9sLVt716u3nMrsRN9siRgwXZ2o1565YIFZMBckpQ5NsJMpJOi
OSsHldFXU9IFcqtwHuxmuzPNZ/KPRxNV4fhHuA/d7dWwmL4Z9H5uTCdRxGCtUR2p
dxs2irJ8I8jvysd01afCUeK/ekJd51XSWEErPUOsDGlN1QTdeOpsih+DGSBgqiAU
JUg6dfw36kXRPxG9UihM6LHSH9xifXctztq7GHDyUvUgwBDF5MyDK8Fbzm3nZX7d
CT/pm4lHBLCZRO4OumbMV9o9lmXGYjX2UAGe+7wYYtWncNjQpKQy1ODCwQIQxSG7
2zVP+k7F7LDtm1W3sl6TBN4taRLJ2hFfZbrgJQJl7icbtQWJ04RTYlEuRWyPW4ct
kHcsqjKmyvFpwt6XKJsPnfM6t/PFDwSfE+I38ttpKDeoSpp40XZL8//9PQ6XCNnn
GnLoHyx58kx2SSq2qwjJcoNd5TEG7K/m+4MbaH65dIvsmDAjyfwAZdvf1IXEgpfU
F9KeT3g0lmhmwzTp+IP4kNcqjWaP/xmchkceWI2RW1XGf13oeAx5d0D65sezt1lj
Vlxr9JkWfcu3DEnfaqMkbBmkCjVi+Kj25VS7CugnmK4nZLr3UE0w46998z9uCbEK
VRt9j+obd02S7YPjL1zWz0zPF70qGlu7YlpHwWFlrXcpQVghAMbsLsbsMyUnvN0F
PIhs/y2mpOhy8aSs/7hAi+HAWvkSmV3VBebCVeLsuv5RoUqkHCRplvV5CyudK/Dy
yLmO41LCrnlmiYgFlB8A47QfbJocz7nMd1WfKqVzLBif6wcvXzjHarp7wv3Ct6WG
wXTPGBKLrvH6xiePkzADuWZJwZf8Aq9BiwAldI5jYWBnbi2K8L0CFlF6CTGflkw/
Yb4q/TLKaknKGWH0jWixy1Ioh/w7CntRlew29vVyzwhbupooLJldJQOP2H5O/SPB
jZ3q5Oi0NLJTqIqfXC7ZKjKlNJNGq+gO/zNJiuwYhmtfW3CGsI9Dsi2H4EdXIYsb
N4He6LwaaFXePRQjEWqboPmUyJi/bxfkG1O8RZixNrVpnQ+YvYb2T70rwpqKUC9k
ZSJ1celcR7pxnD0/1w4fy5Ut+8ENbMLwkrjCsyKp/fIUcq5uqCt5EFUlSuAQs671
vLP6Gg4g33jUAoMvQV+9XZSNYKvBgaz6Kxxc9GBGjP3c/mIfxa6XqFTRMoE+K+fT
fllyfxb7P/JcOYrHMsqpUxnhm9597iqawwDiln3gFPDaCx3vRYLBDzQlpWa8icu/
WIAQ5s2qXxPBJlyE+JGQprUidlTcZ3NNQDjXdIUeFEJOIXr7KSsuqpAbwKwGZt8a
oiXYhlP3/HQI823W8raIzuFZLLCcuROf9QO4m3Dipm1H95VP5CD0moDq9SXwb9vB
OCCDEyPR48rY3MxhhruPhqug0hguxixN5QtG2Xs+Bhm8gIYuGfnyz9rVK9Lk9XuT
Hd6TiyK2pRPBq2PwHQbFN79JvreW4iVWS1eiYBNhqfWu1i6cxahq23ptyif/V/5b
0XkMexyFCOM2OLtjw1lwc1sqQu49QG7UdXa3jBxS7GQT547RPYQh1+wBBFz2ib0L
lhV/4KJFyHJY8gyEZdxdz4JVK9S3XQbH0ZwFb75xce+oT0Of/Lle4UB92ifm+gvy
F2rG/yxM3P+ne4YdOo9sHgtL2psmEZekwU5qMmhwKLMSkzrZkiHCrpcJuAz5Uz8J
iIdF7CwnMouoKPMCCCRWlSKYWQygfCYDSzZRYapVY/Wuo2PfzqtrvHqhztvE6iXj
StSE5yg5ZLaDrdSktIUEdbJ/mEHccaYtP91d71Cwlv5rIOTdCfOCJj5HCgC47/KF
Lcju3lgqLAMYqoR/9eR6+dGCkZ2Z209Ms/Q1ZpUGB27dvM59si09TWKG7KPoe488
7iz/7nf43QmqW8pA5VETQrcV0cLeZqbvMNB4JzWk/aaQRDhvu/M0QnB00K558laz
iIa5ckF549pXDs36yqCaR+3tmtfXu/F2SvFa9avt5LKVENB44bBQRl/k6KTSNO9U
kepSXkWVeqNlU5ELFHzDfVpEO2uwOANnS9g6CGOIDayXZ70JcOc7I7vQFu0yqobX
LCsss02LE3oToTRYjv5ORUtytNN/+32xPs7oNdI3u+3P+rQDizSsvShhW+/bF+d+
2jytPdXxpVktlf0W675mo1FkIXdFGjAs08NO/2q567GafNgfJ4uPZL+W+HvQqmhs
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
YMQwgwgHWyBlYyuBmE8OpLhb8FEUxwBWYZMIDxXfN0kBDidoSy4UwT6R8C1wx6h8
RZ7h9W5loApyM10Vi9Jo4Pw1I6T0jppq06ZWx8uHCMIFZD08TupGG7UHAzEMtJz1
oxdDLsV+nQm0ziVc8D1yCcFAeEvvtsCRv3EiRAFKWmOAiV3nSzJcnu1d2oy2l/7D
vdNoiqWG3EtXW7CkBFVHWl7Ggy0VaxcjTAdD4DqDMlC3yENhRLtBNC7LXZ92VJ2b
2ub/NsRCEUo9ew3tzjbKF5VKlCRtrycnV47qEh1DLD/ta+SgibaMkGioe/j95DC9
BufM4TheTJLb7M8RyNHPDg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2912 )
`pragma protect data_block
W3q2t6h1mQim6Kui91cPQmy0+04QEtD39cye1Id0NUJargeZXiCN/fZ8WrXGGEdu
GZUXKctPHeR7eLQd6K3/fK7Uj7kgamY9FRqUg+/9jEHmEKrWBfLxy0tKJERDlwMM
bL1jJoEbZsWKAvIq4shhfUJ6umjuka5LGoK/iMxkL3IlOIbCyS/tbPgIpmXxW+9u
VVCXHLx7OJAE+glwSRNNFHhhUMN1lpv6zbbSLc+JxTIS1c2YAvMyP2fE877ZFXGX
J4BZ6qan2npNrCHd52y0OaLyqMlI1xVS8ud/kqGDTKuVMMGfstie4UPTdr/bSYpk
FKAvqYLfIlAqnXCGgEf6d+Bi22wPeWtdx+pxVABtceKrwtE3JduONbpJ/1piJrul
jhnRhrMsdUhe8mOuj4iJx4UvhDRxlVqFdUOOBuF/aVUWDet8/G4UkJAi1ur+bDLX
QAlINPXu2LtMTxg+NO64GeN9asAWozwDppx9HJbQ5tpOx+MTYjtYjVVQysv913pJ
F60LyA6BpUJ6AlSzyZ1m7AGF2VLEJMXaRJec9UwunwB0iLj9dilZ71iwlktSp8tv
KfABPiX+24REWIxMmnrRfpilwgnDvHFmFFKC9FZ9zHQjO188RTg0Rhyv+aWct+bt
1ACr5MF74vS0brPw8IrFLE1WWoG/92z6u7u6PWzB/atXYeE05C9D2/883kig0aSB
MsWOXaKC7psp24wscYiwHyh4f6BtkuW6cimTgyO8uFmkTbkfiRMmS1JoepA0vZaj
7QvdrFmS89QdyQkqp3QM0EGTwClKLwPAMM7LQ7n8vRrgRv6C07iIHF7ZvWH+e6Pg
sR7UmpyhE+rUbsOSiFuuvqdY7123eUYo34Hpr2XGWdjIPa59VQE6HtLVAmmqaHR6
noUKianYZNSv/wm4aj6UjkOqjF8AdAfYs6vwP6ouwMVkPWOCI7aokD7lLwemhO7M
jwfbzu5W2EiPelklo/LMGC6Qo0L7gfaDEfaKUs5pw3lBJpJPLpAU53xcZ6AIsxYV
NWZ2eZiPxFFPfrH5Wp9jOAaYDawOV2Q5uAz2C62xiTIlkhvLLZTowKMHF9+wUNe/
Fm4/pNt4FASUC9fuh0JqZw6YuWYEVBmYx2wYFzcfEyHYQCQliSajR704t91w9LBE
xAUBcK6UChuOdbv86jHCuLh+NLL+TH2v8gabQ8bwA2zDMMADZ1Oq51FBFPq3H5qu
5DmemKxuZkBqM8Z61dqdJwigLqzqUfJyzj14mw/0JK1vBVwxAjvyFde1epjXVtwj
x4JtBzTU0lGtTihtDUqQQS3APDkHUxhkhAEVjHFbwngT+t32RNy6xfs1UGbQumX9
dbdpDxtV9Ezt9hibsJBRfA9wPwkXSYN7FlFrwesPkBi7F6u+HXtG5+sHW7fjP9Fr
tSAO/PGelP7PAYfzz36C23fl1/MBhlddD9r/wRQHLgljHBvDrWrn48R56iNzgRO8
etJXtW7vRrkm/GSQeHxuvkGjCWVhS7Hl1GOLVTKe3+q0W1CPr1H+CNjWCdFTdtJ2
5RP6tLsB53i4Tc0HmOufD6Ba5gfeXxG1nvJXVxLAX7yZQ84+Nm+qsVtecTKy6anE
SQgh8mJBKzyWD6QDhFoF/mW23F2EekX7f9Ue5YBAbBYlSia+YSfdBfQZSAs3GxfG
/uegnhYCMtaBJGkn4lIwOGyqgb+d+yz/y+/0+FR/wofVbLGMThUrDethkfriNznX
2QLANZt5y9vmypFUdkdnGRfMIbNcEjstXHR7cGHbJCnaHIIFa7wLkjYkn+wHyZ+m
ik3RCIuFsU8a43N5mNWHC3FoeTw+2Q51SjxCXeoFUnNznlIs1tnk+AeH2ZGmAwi4
+LOxGfQK7Wevr8Vyd3vk1r1ykVhTrd0b8cXQLhlGFNMEwl7GrU4Yn4eNNYkid3/P
0MLwG46PNCIXrLqelKM05R/byZUrpT22SyQzvQSlK1CEJRfV2BW3MK+PsE5RBjcZ
kp1cg2vj0g1vqAqEI3SO/TdO5htTemWIFM93NJv2ZjSQyV1aI+DAJ5U5WvVKOAgr
alMlgr7HUGVDPtX2qOUVaC8ypvAjIU4KCrRa5kg7JG/4hGptACoNgh9c7/xv5x9k
QHUsId3aMwy0dUg9UVEWxT5kWonZQFf1WpV21QiN7gYA564Zbjy4cNevH8iu7sk1
JPIxjWIG0aT+wsEYV63yhbd4e9ydqgGSQXAFde9vmkKT1/EIQ/x4Mi8ZKf81JuuQ
pG3adGbazoblE+IpVnznUFeIGJF3DMUbFL05b2E3zQHJuQU6XgSS5VBVoV6sgMjP
/Mvvk1b7YSYYXOQ1WD5pOge45+W9514zIYqUr3XOy6IInzzmDl4E33hVZwn98vkl
90zzeMopszpfh/LWhG9/6Xxoclfpe3smfpvBS3cBvHi/WSJ8JD7/Iefv0xT7fLLc
7xdVp9N8hIf2g+MwG/em6TSuBvUdVwG3syMq4jYmliQxunp3l/WAOtjhwIPHtTr0
1bYDv9HG2j7A1qY/85xRu39LJDO2eNm78JUHlBoIQgOf3niY/DQq+8ksFYNG3cj2
ZHsonOIQ3+2/DumrFpFqQsJzEebNV8S+3awVCoImPXH75Qa9hE/x201uaopKQXbP
ebQkg9VRoW0W4ZjybivcVB+pjm44cJ79sbEOHZfotDVfUXASG3OxfM66TJYljt1e
FKdRhNe5dcSgsltl/duQ8vKz9MO10VSj8sGwFJ/9tsz0PoEJ0pfrMaEUtzGLFPRZ
fSYMSFKr4kaAYl/QBUK9frVgfyUzfjsI8M+4bEquOPpldIFHJOozvw96XS1OBGW6
KGdI3yhN/gCVHtM3rdyrl4G5OVv2Oc6jd214p3zuR7XbK5zpPVdpLE0XwacAuZia
gM4/R0jf6L331Pt1e84Qj4DePprrsTOh6h5qe99LiTlgeRK80srAKwU9bIMH3iky
YnlqAcFTpxFEw9R2X935NG5KasKyco3GXYArS/35VD1ER93LI/tkU9qc/VdSU7Xv
MXYAGMP8lkyHhX86wl33Sx3XU/DHHMdCJdfMq+32AiUqFeAvs+J7OOxq377M5W8y
eyWsnrS4ExJa626mukE9ZWG6hcNW7jYL5Mg/5hocuWoQEo/Iyhmef5D8BLiidDov
xw4uBLtdsDw7MTddabR94MKTv31VomQpq8L48Kxh20aez7dPto4Pw4/vctoeXrIx
KBuUI4wKPOPL5Gp5S6kohEotXnkmhjGUqa77OPdcPDmyZQFaWlF41lNr6bYomDCe
oZ8+4zBOgYvpu0lxNW/UGd5nrJoT5bjTowQ5GoDDt2/SJiXCzliN9GOV0GtO9ZSe
0kYOakqOSRYMB4is5eHTRxZJKSDsXodEXvUbrNGpyEzkqJNw0479gtzjwTYWjG1i
ZFPksMhoosDmk7Q1eQNxmfJQoE2hoozrb1804QjHZIE0kIV+Q2OC51HU0Xdk1pVQ
eq6ioJ7xrC3QZ6riraO9OPJRbf3Zq9pT0iY5H2cyDIojuiT1i2tFfNg4GUDbQ/mi
Is+Rfk0SjjaSCNRkJVQDKoRTXEjaGni8gFqwdr0odUTqv/1yWtPdMVe/AXZLJ12r
ajiVQoltV1heGcqnfS/k/bINJs7U4ihgecgv9wN6CUyG6P6kLxhcEMfWstnlASh3
EmgtsVisCoNxvKUgYsiCdLwovztzQPa3DchcbXLME3KGOieJGM5cB5j5KjJLn9BY
oAMA0/58rhgLq0WcCTMgLVgq2uTKKzrEpvbJgzd1O1zuXmxqQf3qMuaXoI/oVoS2
S56qfNQjDtx14b/SUL0JFfMrE7GWrXwpc5GK17QJ0WNpylMsGqRC26eMOYHhxsZi
hLb+N30h4k62WC1/ad9eIHO7x0uJI5TpoAIrMueHCdE=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
idM4RZslSeC7U3SUXyCfFFSUiQaqe5xIDeKY0R3vsiTD+1fURrSwkhAPSnqO/K/U
8rGw5fi8TVc9JKw4OYn2oqe05XA4ne7lowM4MUBxxZW0yYEQS42UHwLvUaAqoye1
x5GnKEuFtkE35iybDc186Ts2wH81tHCl0FsoKZeqXzQVNGom8x90V1+8eQs48F7W
Ja1zYwSvbKa0JblqaMGPo41aPz/6IWwAPSVQvtWeaWI3+UFlwCJzg8ahcoB1iG0d
4Yqq4a1WYxsZWUEmNZNjzF+uxXiFkPnHSye4vD63jfUY7t55Dyq+4Pd1u1e2cZaJ
sxP4HVmEbeX6n9JfnrblKQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8016 )
`pragma protect data_block
ecnCsGL4GltitzvnV0I+z29qbYTHSh4pfrceWWNVPp8UHFM1aQ96PhKZ3jKVeHVL
xqco2106NSg7v/441UKd7tz961SbbjaL28C5BzVQNCOWbQMJx8KA/r4YkGRgiN3X
/cqywb3QX/wVtJ++ygzPxmwctK8VRhJOSmYGnCHKdUFMPYgmrcZTU/mPn0ZCkJ35
eQHIgvr8TPjGKyM5JYeQ2ExxKIipypQi/VPHetFAOcd4iLCNhXghGP1vVV9HWYTg
qZ9r2drUU8qziDQnUVVi89JKqGLTIpezp7aU57CnCodA9Y+Lmpc+fBEz5G0LsY+M
PcVWFgprpwwNmGUcWMzdk256P7MqMnh+rJtL7bewcLlPFTA0oI+HTQn0kNhQ+Ktz
Pzogpv+NL+ob5uVL4WR4feoM+9nrWAclueZyO5WY/4rAZBo0lPvRQNetlyx3TgEY
kXEDWhNrSB5Iv2p8bSQ12qqBfmtu35Zq68QdrbW45NF8Zkmcb0dVhVxqYgc5BITq
F+AfDJalN4NRgq6TtQnof1qf5zoWZsxDv26UnRfzUpUL9TXv3qQWlyrKiwihOTRt
VP4nADkSxP0KuE3GFEjxLWVOVzM5UwORtoO1EAXHXRnKjvMi2ToBTUgAdAQSiFUo
741Qrha0T2icrgg4AYs1XgP8oZUz2ysbnyKn3tpep3fzybouvSK2qCwKfaPfDvZo
zFM3Lx19yUf3i9bmBmrBPw26uvU7GgB1WIqpaISdAX48+XWQT5pJVUF0xg3UpxqN
vwk4TjxDugkct6LnzY0g4aYtdf5DPk030s7VkVdrS8AXtQ8k0gWTG1TyfKUXvxCc
IRPDtUduo1wG7be7Yhuzp9gcrGw+EfvCM7/nHmDh+Tb2GXYP9Fzt6HJZfCH8SNbW
8CAZlU3zQSWQye3eQlMFlnRI6vyqvlUPZICQozr1mfGsCLXw1u3AHX5vxSSiJ8LM
fU318NFG8WeVnaGefqyy5rEfzufN/H9jZ3EK4z2z3Zv1jJZdlptWXkx3NJ2CeaGB
rX9jm/r8Y5Qc0pmgTwt3nz+t7BcEda4KkZZDmxGrpS9q90BWBc0jUlJwJFnLoON4
vC+UExlO12komFiMbXZoo2cd5ajjpTSE3OPPqjvEhv6UGIWUwfKtozU4jNwzIUCY
mDabeK974OuptZmFb+uCY5gX2TYh6TZu5ZU35iScOrMKaD9/0QgSDVsHj6gSR5aZ
Vi02PVraOJjiO0dGl9U8zkn/XN8wg5H5QErXfgWmsHy+Z7wlUQOBxI87OkGl75tk
03WqCWGnpMLY8PaP/dFGOLSJva8hR0JwzPEhleoow4W8+4zo9KjAlwcvGHfL+RSQ
rhxNUTud8k4ol+HKXd2ksGEoUg2v+29FP83liQEfYjj6XJLahrSXeeGTLeTZY7fq
lwn3isRQBbyRvRrL9+09o2u0tMlADfLr3bLHrMl+yM3H/X59h2j8v01uoi5FQbAk
5t9i6X4Te7JqLqtY8s2v7CGsdlWC/u6Tk8Bhgo6+Xn9Cz6oVDI0dgcdY4JGifJ2y
PHj/2v5jSVOKJSV6ql1tg2wlqCT4ggdhExuT6aDWLArxlGYSEHgovewm0CLM4ue4
K1abL5xtx/VRozDSMNNqbyJZ1KI+TkKIam53UkWVPBBOgVcLMORJiK96Z3lbIbGD
Pimff9cqbSGuSUYZib4LedA+7FBLimNHdy6eTeUe9wThVoQ75jO5cj7pY9XC7tRI
XT+k8gm93pl4G24N+980qAS85Y0dksblgkqV/lyM6oC00rY2vYOZUS5goPPfGB74
IpqP4meE35SW81tnkJsa/UfPHMsAVHQZFlbEBELkw7dby3uLzdL5V7KU7foRWvGz
eGuHX28Zew4Vm2dW8mOxfV7tUD024KQLJ228zJ+/evaqWGBWjaC+dcmUkO+bCxVR
OufYLeRnAzV31d7d8ubhI1Tcur8tOzcVwbue/MN6h/kZCnA6gbTKhUdhD2BilE2N
a7CI4BagUbvZdEdZULTC5d1O+f8vz2KQFIMEC+gd31+WRv3Vuex/VxjFzCSV3zyX
siAvDJCKsHcOmznBMObvMU0bTq1uYYTnkn72VmtsaHt6IjmTyJED8kOo5Bb4nioz
iG5OeBO1z1Ran4wmHhcClqn82QAYertG/teUefxPid/5er78AMFQnTmaDakrRkbx
Y+wiwnhnXfPjhBu7ibla86Ssjggql3+MejZPDaFJ0oX4ljXb8imuGsLDHNFjogeX
WSN3JbR8axruSODFQ75397F4xErSVO7XZ3RE3sacnIRWp3rGVj9xG/pTIdwchQWB
VyJKkreEdT8jgoRvPuEE1rcb0xkIT891tCtDi4TgUKAgB21mSQyFa/Jt8TM1989G
vLBF26ajfs0Z0h53X4g1anU9r+cfOuxGTUh9UKSdwq9QUIfPdL+xulCDM4oea2kh
eG5i/uwjNvTmjH/phBV2Ey6trn5c0rlhPeb/tOtbjj4diz70GXveev/djtbUKj6V
auewYnl606+Kuli5c5VxU9AvjH0GTjkTW+mFAWdMqgFS+8/O7OGM5mzpNsHEOLNV
jWlRbhkit9wYx7nULAFCxysx8Yve+aswL8uVzVLOytTQBpyNUi1bnjHIfPR+aW4S
nb8voWUd2LBJLPVPQ8erU5KhrXSbsG9/OPFRtPiNwhBmfgJP0Yj/7Yyoefiq19dZ
IHUD3NzGBQp5MmhJhe4i/ugV0YqYroPIefcp9hWQ+y5J29T3V8yKrJ4YG/C8Htwm
O2st0wrRMgigSeRmx26dpA8xS/qP0UTsnsGJnG7X/R+sD7meFgGEvqqyxGJ/oI4U
9D5vqaNHrLF7FmVdp8idGWMAtY2pQa/KHSamwCz4oq3tkBZXpO4Kh0HglZIFlMej
XhgMV4pSAi8Fb3k3lh6/QYMGFQ0h1efW+S2nbj77q9WDKbT/LRJLBYL9Gn9LCGpY
FKQB5/rAQ2O+GASHKYh/mtNMzAzsRfJ/zKpwGtjRDO5rs7rZf1rL+1e+5EqVlvJG
N94eTAIdn6eby6a2QPkfBpNJah2onWm7jZpcbCMkmEyjqGjTrMslssWMj8oTiIq0
yagsvnVOI1rM2PJGn1VbBT2JVPocc0DvVyDT6eFukXGw94Oo8uLo+uqCFjVTXz4A
AqxzkiHYywwcWRnMBcWUndbvef5048MlatErjqTfv8uZ09opDXdS/OJliQGJiSSc
tzhvJVrg/sQKuNyxkpPw11PciuqQvSupapniqoewFmNRTkBhtpYMjeWR+BqjgklK
GXdWY0DbygbI4O2RBPEMQnFAX3wdpzxQBV0R4+3aQepg7ljJtjZ628mgjL4oACcc
Br6Bncbnt8dNh7Yo6hbI/EEvIq8zLc1JIAf8wD9WGLP9J9H65RqDMhVxoLzJtCCb
ISr8YFQm+hHGK3jpONnf904aWCoLDjlBgxRwYw1jGf00EADqHtc+hfn8VhNm1Nh2
J3Bbx3Dk1ehCrCq66BCMuua0ET1d4w9VB25mek1mxBLt5BjHwzRGdNAMLz/FhtmX
iNNMold+kEWgy7VTQ3QQAJy0emzph/PKkKvC4/K7DETwQCrCwwdfO6McnLnGinwK
B3wfpgojh4+DVZj9a6aadO6BsdkVMbYRPntFnoiXTBGX9DqcV1i7IN9v8Ln7Wi3b
FDql2xaGiWhhNGkrHSVJJH4oW7tiMnD1ceiAtWDnTObkHquqT6jDHDJ0WPSPVVwo
xzHG582FNm0hnNk4ahkhzVg9rMPEcogVJ2FkeQLWuD04QEeZix+Zak/K9ykBhTRG
uWQwkB6a9TCn4ljOUnIGSQ4glcJzJu47xPNG3Gks24xvgRk3QPdE1Y9MJllAyLQ7
xxy9Fe/MDovy0XzA4XZ78ZUvLyjGZ4bPg7+6sr2DZp1ZbMFrPYwvPOblyVEYNpyz
LM97ABUzLTYMTESUZLJYbZ7bk2xBL49K3UV+uXLViaf/PlnFjVrrx44DlWnf+aeR
gNRoGRNGsLb60Pd8WQvj3urxXdx261XcxRvRxS5caYDjP3+T4nsaHsH/UcE616hD
j59ioIMf1AfnjVpjShNYI5ULR+YsYIJ+KSpLt0g/sHsNu+XDDZwb/eScXIrtIzJp
Ley5eGS1/doNAGOZNMtLXp0ByVRSTQ1ET97rNyaj8rnADe3uIBRCU0jQAklotmrK
afCLLHDddqc4sKtA0QSd/fIMVOE0DQQzjCMRq4nMrMZAs64a5g5v9rKVumrYwUjm
qF/8r2KyBYNcjsZN3XwT/P57tf2shMCPfqRwevknuCDMj4So+SiX/nS/Ef3iy8tt
75FDCPs8izb5uWHUPuS1EWMW0wrtpOaNitqankieOeukfqxw0P6ZESRBFoeltotZ
ERU7obVNCBq4dP1DUGigOdG9E6pic02ilm7Ep9brckgrpJx7TiUXStizQTECavr4
5AQCqNPRcJ0G2o1uLPytzX23yTwgW2IikB8f4VeeQ5wKx8DJ6ABp6nCSqlO09zb/
D2Ix9j8wQRt/pOGikCzJWTdvj1kOYanSpXfLQImy7Pin/3YB2IYxIgi0jYYmHqNc
Wqies2Ly91IbexaT/KpH65oY53SiGUVxdcdd/ioKnDApqCZMSSPGQUXIiMXIj6eK
gOFOvZZ2EtqELxV2Gu3LBg3R0ccVxp5RdR01iqrHiO1J214TY5w2UsAaJLXe3KpB
e/2WWNanlByk/v57PMxOCvQcVlVi16LRJTZ6YC4EVpy4m7dHaYSapQifEuN8ClUZ
WowCMeJbB8SR+Bc6PlCAatjOu27WFGMjqbYah7ft7zRJTDTI8m/WbZyoe1i7Tc3w
4dWjhIhEPZ6o2DkdfR+bZGBQE6I5x9f1yKq+gbjMm+sPUqs0EB+uduEVDSYOBcJJ
7NmfQRW2JuZvsEkW7CBHjBOIdGvXDDUijlS4MfjHcH6ArGsjKU5PAoR1lFGpvPFY
6IMqT/LjuWmudcvc4+5LSX7RnjX7xcJEMWJ0fq6o9/ValAZ5N9YRmykKqGFuQm9b
yDcCkukYKDnIIcX3tzOE+9Zw4pyOPiZBwvY65/1+6RunVQaxw0HW708+doBMvXg/
iVFjYQWDnLYxd+4NglOx5RbNwa/IuqwiUt3CtMFBNwtRK68OFij5Psab0bR5WqoG
68rzhr2VJef8JUxsJvT5hIP63D+tAHyCN+x5gDrouPqVzrp4rXsC7BAfjT7WnFnW
Axcw4o7dzFmsfVo7OYPIfxB+B2o54p6iwMKDgiGxAG1QPr3CWsKQvgdT0skgF3wo
d1oBtOjg3D0xDBnyaHXh4tMmY37PqT3Za4l/cwXyFR0JHtSk+Da7K3fTP+dDsHcx
v/ou6uV31k9xRuUi7K3ULXQ4fjQhF6Gnv3Hi+462nD4Cnxg+UX7aN/15xQ89mvgZ
/nYH8PGjak7C0/P3R2q2Oypc/l6QXvgGpLu+2pIfZUSk/DchhBbBgULbinA1TpQv
wkYAs7gOGDM0qsSWCEPAQot20SOA4feC5B1PJyVHYlKwYXd0xbdACeRscYDpvvFk
GX6mQn/fDgr83HvlJhhDSmzQPXxJ5RVhWXLptSh/mHbQIqjYol8ARmgBpGmKROsR
Q7g+v4Ami8V/uIZXrgxkYKSnHRmeKstpFip8U0Evsqn6A9hx9WSN0YqZrcAo84lq
Ni8N8SJoffwoSLi1y+p+QDyzNz3ip8WSaI566DWl3D4CClG0G2xgerqQL/n09Was
6u1WWsh1rKMZT6fYKt2hNrRmaE0Lp6uxmPwjxIOZvIBP71HKtn0M/k0Cc6nEGsJ0
hrxNWvyZER6O0I+9B7IWHgFZrRm/gyTQtDBYG8cEfdC2wb5bYvBKtgRk1kWW8BRg
0k4B3caS9Gk1XueBcxqIMyaj07QeAgG0lSt7mqpRm3exaUGl7/4thYUUuwoYcBFJ
JOcRRMMTiDzucKPOftWP6tGpRflVByJnOSRmM+QfIr5QODdfMMV+FKJ9izWi4NWw
Dy6T+iZwCEZPySavyAW6W8nccr5ugK22nJRyjAsgvh9swh1lbvHXl+fJS93FUm8A
VkGtdtS38DvohcdqR35fX/HqIFadz63G3J+cHH02ksF6wIp6vMTv+ej/Z5ZfaqoE
p096/nuQC6yIFSFW8NO+PULVfOfQpmYZQbeazka6DRm5J3hSv7a+pxL5Yder0Dqh
umImJlD82s1Lzy/MY3xOxqqtrlYfIGwp5Bn2myd3CpYmF1/tdtwjWa8DW1sG0PSN
02reQMNxU1Vp6dAz+FKW+/m11BAZNtWTmArggPqJVovhO7hr052xsSK8IacMTCiB
uaHn1Y+TjRTmiMT4C0HlvTwNvKIglZnv15CeqLOqPw47kUwVz/ScMXmMfZsc+iGn
ZHyA8LI3PDKDdC3GQWG2lbY6Sy5muQ5k1LHYA8l3Pup4BWMG+SOdyNmJi6zASvC5
IugxYPnn1N/nb5GjAlX6vLOm+PqwWqq2Dzp7wlMLHmj/7g09CeYqE8hupsJzL4Al
hY2bWkbkRZZDZocdx9MUMQf6yXg+McGmJT2gFz8YHtixHooQGAUsRWRaAZ7KhgEp
WnvfTmYKIiMNbhPcLJLdMjExT/hY+L9MoUqeUPIZ2fhY4XL7LjW95PqrRXwBTxvq
AzMU2A4MB0UZWHREgwomStH8hbXXYlEte2SgAfWtPEEgHa2S0o3dIrEA8ZDwgEKx
S18wwQonxSD4bS9uFyQ+wGwhab2s/ZO1L4wwAwV5ryciChsO4NuxN/fCjUiaSDZ/
BvcesoGhR8+RdVYBVVlRpq/Wa/Lw3dIImcF21E+ExP3CKuE1s07ej2L1gAq/gD+v
y04hqAPk9M+OUoWVF+CXrwNlobI+EoTkDqyKCYhMWAIPh2gq47+Qyf6CkD+zsFzw
OyYOMg3zX3+dx53T/iNli7vhuazpbfCh+FUM5dHVluPKIwFtpcBkEWpMmkm9T6YM
rmFGWgAdGdO7qxjavo3WN2N++5sXgRoiP1eHR4TT1rXUxD+EwD8iN44HUsXS619/
VlTkAnS4IJeOiGblvNib/JmK/IseHxSZ1BdibCcZAfyUpCnkfp2nPNQVUYUmKmz7
S0uKxvQk9v/dP5kXKtv5k7OENkkAUe9US8o1RiAO5ZzxlrwDgdd0HVfteEBPeXOv
HDty2o2UC6HbZLN/gtkXe5a8nFj3tem7ky9ZTS+/9BZOkc/Xojg5gxBPSSesqv7a
my1Mn8O9a9m5pV8ek5eJ+MS/J9Fkx9hnrgvQmPFChe3zpRVqlfyTlmGpNhNmOZTO
MWEzxSrwbvS4S3n2Vd0txWfUAiAS97sknpbQxiD525cQqOqDeL0V2E3W2S+9HUoH
x8T8PUyAgp2anCS0zfyCsklOUcAKYOGo/uOZ7odwuV8I0fgRvfgh4xWC8Lzct0Z1
iMQiQU4/HwVWCuYQXAJIoLpW/79AOH1CdcThq+TUMm/YN03skjVannFywZJG3jLJ
8k2WU3wJ40SUfB6dSACGgIf1yIwogIP30yEyblOk7G7Qx7wQ2tBduY8ebHtYUqZt
JDHPCm9tJ1p1wW+mR1jF6UuKins/AKah9Sug67ZFk6MyFBfSQ9deCuLaA/s7WuQi
s8sOpRHLEQFHyX1D8NZ1WysxqEKtXcqHTj4oVvA0nHzIOcas4wDxSeC5DaohG/My
pRNMZpitTKMhmpWWcOv6O132Vt/dEYwOdylFEibvf7QEONxnbVnHaezb3lzdVZb+
YKxv4aor8chuAYJToB/rWA5jEnZ6x4h1DcgCJu3NXs4QjzN9XhwRPJxq7+Gsv9gU
L07fgthTYgtxNsZHZ0OBBDsZWtYbUXcu3PkdjfJGrBMLNeckHyGPsUvqgBCuK2X5
t8SttT79RMWVEZ34PalfzGIAl4Pzr753F3fFvdNfFumiJ+GCVzaJJSqOPv8UgCu0
CWH73DTBJR1f9tG2ly3+mx25IvwWX+sKlX/HXKaScJoabm+8bZQEOUdXZv1uFYmK
jX1Ecvfsbwsh0iQNVvM62Tt3AjtZvLil8qAFINoKj9vTW4eci1wv1AlQ74vtSSrB
oyFUKLtmR7jCHa2hU7taKhr77M0uK0lvXlgDp8zUz0JEIyARlrAFIokOYp5FsmwD
nIwm1zO0DoD3RkVciBNg3T78dbZ6q6zjB0rJ/HmC9bIvvurJqUhCrI5f6xrWgvoL
RQC7pDj0/ng7NhWaXr1zP+kJYerCO9PKRk66/7vhklRihHqLyD7HzFZ2rkrRf3vu
5fXJU5EsMlltoHcuDyurfdYY1O+nj6FNkryy4cNLelPtNnXxjkE+Pgvqo4IKQZQX
8NzDeIaxKC/ISCNSjOqdE4DCyNVOEVTLa+flZ65J9tIAZqguDKL9Mf+qZNwc0e2E
59Fj2lLifp2NDpEKQ4/aR6yfKSaIaItXxBhdsDQkCDyayciHPnBkIyJgNoCe8Lp8
maQ6HCE073INmtrjLRRrJqwwtaC/vB/f6dECf30SrxWYgAcTv8TTkjuEU0dS5dVA
J6MXRSSD6IuGuQNj5fA3/2oPMlChikifsfUR076la4hqXQzS0kI7Rh8ZR6YDN8iP
7G4nesO/jX4WNdFbjeFRscziBv55+CIhe4fWoHhgn28XQOf7dR4jVSYh699DeFGo
qdVWhp7+SUicX55dKIOntlOkdyzfoco2Sy6ivZdMxrYjAAF4NElEkHqnbZYJbhWh
SVH4GnjgS4m9TwEPXnVaZq3KWsB0ANHeljuIY0leHbCUBji/0NQMXaEgJeJKI+Qy
Fsea/w6Hese1HFQT5NoAnEAKBTN7LHVMd7q7sMaDNoSPPq5flk+pPFwGSWVeKDW3
bLiWTFdYX92RgMJR2EY1vI/GL3jNNkquMsH//2fCotESH9Msu7s8dAyeLGF5Wjx7
v/KvpvXsEe4w1trwyyswiZp0MykfNTOEA+RXav/wc5Hx65EKHDRw/J1TeR4PBPtf
J10cCElTuqHxxUGfEyY4AQVNcPVtTLPpr3FhE3IWagvio5gmEeuqwMw3YdP+HxDV
9u3ldA0NelnTntktumqcYtaSuqOITGkK9LLEyJJt7Gw4MRsR0zm8RU2VocvUH0Gd
ZLx/NSvnwl2J6/G62qeOFJpbYBYSPQ7Ik1uBEuLmPgqeBnudsAitCt82rExaUdEg
h5TlgebqW+dlDcOW1c9fuyX04EZ4uRT2lGtfZMQN7ORWSiPdowQ9AarmNH5i91qj
idnt7ufdUXM8lc9DAbOwveWEgEx94S1JIJPQYx2d9UKhhdmY9r+EKVtK7586pqEj
NIBHPhXIsw6Xqtps7SkY3nGptuxHVRfuOr9X2KyLN/fUKBHJ2+PjA0FoqcLJEvRI
/vTRbog2DIheELvThBaVN+dUfWptaez7iz2umWysjVBPSYcisPkZtLtcW4mcJAf2
OiCmDBtD939J9T4ZRr2+CCxV43spD5Xhcn7xYGG8RZlHTtpG+58W4uSxaJ/SOTG5
C8QJpEnLOSDGT+0PmKgbb7QsnVoHOmGtwWx+6w5KkBd8XPQAryRD4rHeJ1YxOD1G
iw8FMyjnNhMp2qmk2S6mdsUqj4pH3qc7o1OpFhh3HiKy4tgc2TeU+/fClrBUMsNX
puLHCzxYBhVVKNVao/8o19RUav5CFLdj9fTBRS/dNJzu/Ua4aDILMVzTD6u4B9+l
hcmoTY4+6q7D3062z78ZYPY7T5tQZCwMYNVlKxLGDujwulj5OM8a56KRuJfgXmzE
hM1BNF8V4fm7YNdJblkfJ1w+cmoUT1cz5PQdRhAcyXKcQThSL9nna3mAuds/dqb/
AT1tcuGBomuwvmDTIPEO2AvpYW8kCFHQ/0da1Gjuu5RXx6uQvUWSOLAAKuwMf1Lc
yKUNWDlfkrxjHLfkojSRwb72UEjR4KT4LRLnmV0TTdG1LFRnN6NQIXKb+5gVVN+F
t8KlXOe1Q2vZ4phrLYPgbU+TaqX4z11boVck3EFpmK9HpAvXHhxw+9rO3/ypZ6sP
2n4mGgcZ1CDsHIs9v72G3XRQsrXiyQscidrGMokReiWhjejv5gqURR4U3ZNk1ptR
fptPyJ7Sk13uWlbx0/SLx++dAYrq4Nsz/70LFVvAqjYjMLp20JLqTIgpGOuqXXQ9
+q8NCXkqIQRrGykQBiGWzNMahE/kqGbTRLxxF8unExNNeu3NrlySGs4mCA74X3f1
MeY25IRwC9dCSVB7hH6Z1anBwUWhmX+Ebp+XnGuUC50YfUXx55nXeSQWTbMFBW2N
tZq4pdAuGYh12vr+fcNkeltnM1hytD206hms4uxbT9+Pjrq5uNd3UyPPpUrgTXms
/XoOxRyDC5EEabPp0IxMG8mo7kUPZntO5TW0NqWM+XZUqnLofNfXHSgpVdYUvZrQ
c1dIKnzdsJYNTC8OEh9D+RTB5uNZc3HJ45N/gSwH0NKPQUAWVVE3rtB7/Sw4VqPD
KUALr12dS8BtZlkDmRyPn/UXNOYuRcDfwLLtRxhB25JIjqZCO64W/BPpkRtxJYlx
OYiE4PTQ3pCbu9x+zQ6pzczQtuesJjxU1ESatZR4S5IkdRIbSPdnf+g9oSRThVoP
tnGSk13MQy+pKWqdi6Ts0PbwVH8cMeDgOUHisifjgcrT9UR57WmYcD0NcYLe7MOT
MFm/SsqMeKU4puI8x5WVUoiJx61iw0mugu+arUETBd09sWR7j2jW9hX7THg8LPx6
sF6i4OTfN6Fp78yA4U+oEfCgQv4jjgjANjj0guPdkozl0LXH8gXlVp86ASaMoxu+
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
BVqwd6fKTZ3R9jL3xSGZqGwJDcGf8BkEFNMemWBSzOMFMkorJ70aTerkd8djFnj6
4sVPtx2mvGcmgQmxQmVViFszd+Hav44lDHno02bak2uPsTu5BeMbaf3dQyJIWcfC
XwCCfAWRUuZMIs0HWvotfBWblpgzNxf5adq/PeMfh2MGs6lxqpUhF5V3hYfDgm2j
rHHuqkWjgwvVM2Jh6/Kb4+k6fPaA+snew4G0Q87YHwbaoKIivjpTlOjwZl3gqtCB
tLg7GDfdS9U2bZZX5ApdLrcjTa/hukoezVnn5+5ewFC2Qb6NR6ulpXGImwEoJSIz
CbwYq6lLbCe/ZKrvLlSzIQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5392 )
`pragma protect data_block
+WmHH51vWn1wmYmn1aJhXSeJkJS3/fMcXWaa/X9FvZ7nzPf23QRUZZoWYR32gmcP
1NEMhW32f/roNkZ3JMbShwqzVTmA5RUjTKve195QB+0e+ZhscyXYswgKmkqs90cd
7UDr/Km1GVr462i3hR8mWqkSlaZKyDCcI029CwH20WdO0HBi8oyBEYIRXfNVYsan
DXduuilRWDRAyexhwzsljDqVwEpcgqRO8UhgflxyNk5diViF/nZR7GrO6hfxERcF
EBDpwZXsGicD+CKRzhathaBX/ptNqMlP7bWP0QwPgTjBIbYe1TKd37UBoKXiM44/
V8DGtQbrtuQI0Mm3vdL3L8600Gq9HQsxX9/iEgrt4HV+tskvl2Kd+VG7HJLaBY4w
pt7uE7eMuJJQ23E1bHH//u9lLYEMcPF3HextqHv9OyIjeyR00tYtPON3GG4xFhGy
HEul//9JX07Mrgwjf7S7v8WhV3Rv9EvHpDHU56FT4zTc+kA5VJb1PUHPtNlN6CE8
D2bBcKH48+sgTv5Jsel3gFBzzr702CcJ1wFWEeKT9zKprT6NyGAK92IokgwtQm5z
FwXquzcQcWK2gOLlZjaKRUpdljQ7dmo1zfQ6z2E0GTuygIc4/q9F6mnanN5Z0roM
VuB8gc/t2lVyR/ovlKjDVbN/tOWS9bZZaoTeWp8NAfn/UvI3fPkPKtWVlkpnUcN/
bW20YMj5NdQFE5OPrNJGtdbAtmuaJR2ttb/RUVPItVhHVxYJ0FbbaOiGzHhX9oAf
P+aorCS2LP5WkiOTblPhoAc23bGNYQNPyWKWyhvO0obm2vsSqpdQINVU2qNQnXxH
ucjwTt3ZWYd9XUhb3Htc/0VOqgUE+Rnyc97f5X1dstPTVDJTjyfIhHU+e1T2fjn3
yJJgsQGsNEACoL6PrvLEOP7FuSYWAmOoxVcl5VbQvrLH4ltNzix8OkizhQgaP83o
swzb02OmGqvhr5f1ke4uwI2NVJR8IZ6YiIIWlp7wGFhm6YvIfBXLPT52UUG4a+zv
ncj837coIV2ZankOkTmuqK4rdLOLAqFY6mfUUBxifUBMzp2yH5pooLtzHObqGIze
PRA4tjiRWm29BR0ob/36Mr1jeWYNhFm3MnloMhP9YZV9Fk0rXYwaR60YlItbg+fQ
Akj9VLbCyZZ5iv/dt/Ud5B2EqXrYSMQLW8jYtj52hGbjI0pjoIwot4+qvWF/Vr1r
tl44X8Mks4mAyIhNMz7pIwMnl35HiDcSKQQgcW2nFvUnn8HHj5/DlYKhbp8bX6Ew
KaGL9JDU1oOHrTkPFXB+UdXw4u9upxAWDgOrvs9usQqMLKj3Vv3NP8UL/EdqqEap
XeDt+P/UBVhfReHBbxh39jvc/U6fcO3AAwsy88fhto3/yhKOKhijg+P4W0+Sd3SX
jZKr0pHd1zQJYxlmjFAyphnvAdYtL3nEtMh4/ES6votFYsFDX11ik+96jcKbTysk
iEAkjMOIRWKT4FKK7wo/eqtV/+xd3vnRdU8GeJ/4/SVQwiWQfMmbMJTJA/dohWXO
TSlRA74FYOAs45e8dqjmcq7/CWFnX2TUMGAANdc5rK5iF1vAqOMTbO/CrEXhDvLe
NiXorud5XnZCGuaOIasy1KjJCjKrLqf1OVQql63kTUEHeERqRJSY4/5ri99w8LsO
EF/1wQ6VRI0KwslofIvK7SWK9nnPE788hKpMNUTIil0Z1rOqlq+3UunRCt6p4Wg2
Q05fYxMo3Yf35fALfODasfHSyJnxb6dy32iv7sozzrNIU0wh5EOAGPqKpoG/JR7+
tEyY63rlznUacvEl5vcFUkEkLmJtZGEuX93VHVE4v/MEBrsqOgiu903Zdd+WE/GS
cVWEEg5P3PelBrW8ymCBE3bYXrc7u6ZBWFkDqgFS1EAy6jeK02GufNbuUqS2Wnfk
ZHsi80RMpremPPZCgYUaDByZSAm+Tz4KrbC3l5+pkUdisofBIQjAimejXF8kkRF7
hMXVOCxlOFsZKE66H6CXxrzNx+iOuLzdmZiHQuw34Do1rY4yyxVKpSXHtsVtrpiM
quAlydZn/KdWHYnuwyHIRYC6k//HnawmnMrYcPirLfCMWSof+1QnAEfAuhMZGd6Y
6nnf5wXh7GIoH7P9hHmO5TudeEp+g6eipjK7qa1K/0+nOS6AAACYnEcjft5IxuEs
NpLcIgD+l+FDdUdumiFJT0kguHwu7omNF94kr6vbFtvtLE5Aern4/lABIuV8Zu3C
Vojav1dDpQzjlsXw4lfmgT+nAH0FA+tdeH+7BZN2y9oleoF+Xr/ljmnAQABHcqAp
N03BKsWVMzCX/3449TZvWZJ1VyKMaKISnEBsFSlP8gkCOIZt5JPKoAxYaHimT/z8
hqIktW5KXY9yaQYnAQKXyAlJmdHPRzap+V9rFtF/1bdbWuU6uc+LtXLL3Ugwu0fv
t79DTZb5Y/D11ARS1/P0U3WDw+Mg3xQUVG+2F7b6RE/l2j8SS3A2U0EGkrV+w6Gc
RTfLinXyuL/jrwSmU19UBLBon/fg3FEwCyAWYF6sF9hmkeMAEw6Z4UycAxWMFB29
I6EzN274QkOIoiEBAUZOuSJRPEmHyCmex9xuwUYHldjGQM4zY6rfk1gtk8konWNi
SMbURoqmzC/784uJTisFyjsvHRY7qDc5EAm+Yrg4UwvcC30grS+XLNYzhHiz+rp+
bHhjfueEmuYXBFyzo63XB7zambzDEeI/qToQQGVGOt5zQJtt7+R3NuPYqQPwSzNW
iqGVZsQ/bZLzjoODul4UigHYWqq4s1C7jcUZlDMYNWoO1v8Z6UMErXhXQQh2XlAQ
iSxmqTy+e7zHWk5gNG3TrXWVL3/LtUjIaCcIhZ5b85c/3VIT6JOhZK3phHV/Rf+8
wHHD6R+m4YSC0qI405iUT8ZLWweZckVzwtJE6YcQPWTK8nII+/7xA6Pu/k1e7p6S
Z1USTTgFtFBEQPvaTQd1/WRJSlOgash/FNG7BEmyRN+bTWDy2j2Z1xteOtW/dz68
MzGAVbLvptpbfzQLCYpxP7NxxWuIFug01eToEioJXQt+cCQ6u0eCj9W/kSLF3UVD
1zaAmaynoIgLqMJHJBF/iq/chSwJCxOAXb/jpxmBogI/qdIzFIDw8TfCRrI1D2KY
f/ufp5IIr+d7jZJulu+CuGUzMpol3icjszY8zaYL8SGYeeArz3ZjHTwM6nxASGDq
fkmBkfHOXbwxs9P6Mwp7NKfaNfRaHtsblxSk6NMBTtv5Rqef8SuGvhDTo5mX2YOh
pY3ckTuyGtlVq+StosKidZwAUnK6Hv0gs63iYVvrQ9dTMUjb3kVnDpYm/jugasyb
cb/ffFr7D59Lzkjqi0V7ytI7WIoEsN3ol+HbDnjrsGsRe24/61mxADY3gwImRnMw
BOECmqhDt0D7W9+fl15w1U4KjWT/iuYVo8OBewKOrKSlnTdUDJmcLHj2B2Mx1Ewd
xgnmyOjlkn9yyqnAfpO5FZ/92o51mZzGinwhsOb1i0v4s42qCTnsaOlBtOh/4pE5
3V+ChxOyTKZoqCtABfnTm007TGaanzeWh1tLgAWY4QHLPxvFe46Bcn3t0qApv1Ba
ji7UjnlF4VCAbPC9VSxNEW1w1Sk6DPgiBwWNkUi3otCbaB/mitKy9lV2WkuCxFVP
JqSTlOUF5B9ECQ44R3a8drKMgEtuYcAhpicVQFAxkCmj45x6wt81fKwmqEzlCeUR
pHvg5xMbakSbxeMwIa6gUeV/JXGvamDrccVTGVdZ4xDMGqANfq8KhfYVWNbk/Zid
qwLimqrNs+Oein2/DWpo6L11O9br6+oPtTBLpeQrj4YeO4X/2RqdFptP8KIiXJQl
DcCVbebW45nswt+XTUGmMnhlbG8wbPUej8l+0sgnjjwhxNTkqVdYhc/Vo3C47aNZ
40LwZ1VgG/km0llzDf1OfLKBaIoHcXsTTih8NulzRkWqj4KRa8KAWhoUMCbtgeMH
I28pyAuhPtAB1Pq0O9g5ve0Z69mHmazgRPDO3nxIPmWzYArl/WVXd/vlBk+9HDD9
Dsr8uUTTxIMV5j1X0FyurZ/zsft6GhpJ+KkLZ2RHgtWxcyM6orfw2/ZpetMANLPI
I953CLWdG+mq5EeD4VgrMMTT0qNBu+UXaAqSQ6f/CYwUv97ZtXNV4pno7RERMci+
NIXrucWGpOTRftJbzP1ldwaxGr6nOBGNGFxjX6rrtrbNnm5y09KGNPM8WYZZEiEL
dAUtOBPkg6OSIxys7kns/65hC1sBsrDUVLpty4HKTv+e4TzJFqoFoCMymGAFE4xx
bYvlsP3wS5Y5W7AGcQj1cIJNjn6LjOnw1dlfw/rllQJbtED8HjFU9eBzR3W+1qhU
T4/7NPtTtoBg9gAAOQAt3NYvXNFxXeNfafvKInSi2OK6qH9vy/cy+kI+geyCZbJK
PNb4uIvRX/8zzwPFamPX0JckeWkEt9OekXA8/RhAjlxPhX8iPu7gUZMDy7B+ZCWc
D4QAZ+chQXqy/leMT7gyBEKc9ifRMNwMDJdfeNLaFD9RsEABDas+vJL1XgrpeT1X
bpEhcjvF+zpHC3nIekG7nY9Fd26GqZtYLTpDhRWhK7rfqbQ5vhC8S/3MDwU2Bpfn
Q+pqq9earFnuFrScegKifT2KnIbg3G3kXg0W6saeBOpLaX9W88OETlXhim19LcKy
Fd0TbmRlzVaiEOo9/aFGRe5DjuF0Lqjb77bzcMxec8t9LzlMTdtz05+h78YKgyGm
MpzBhrv8H3b1mEhP9WAUwbNR1T8pp8BflNns0+PyzWPmrd95RT4qOnGzjSWwe1Hs
wyrORNsfA9D0BGs0wEVjBHd7kAuYR7DWZitxp2jKzuB4LsEuNHq0M7hQwiBxGELO
ebd3sXQLU/WrKhMlzY4tArGGn49nlLWd0r+5BgHfXd11F8ukMMiwd7vo0x/euuwF
mSJebo2rb9KZC3DL/Ad2NIufpw9XvG1FbOu6YLZVWv+tF236hivwWqnFJRXuV36y
N0XfEMpRQEBaLQzzqIdbXYw/0j42l85BbZZdnsIgbKjptYws8Fn0quu2l/QXKUXH
5TJ1OC1gXOF1PhhnE7DGwhs+y+/qG9w+a7ZdL2HQPCNK4GnzMFUyibt+E9Bz0g5C
oZOpE2XnQeGQhzi6IvqYz8x2afWa32EI9ud91P0zoPynPPFSsQn4VdNdt2ElkduZ
jNURuLfJgZZABKb55w6bYhAd7sqZYyRd/l5YxD5pzg/sPKuHEYKAcosea+muZI7/
MXAyJYqnK5rgzKLO52iSDqeag2/TpIIfzvKrJO9vnjOtay0Nsy2oqpTPjcLc1N73
oI+nTeO7oFixpZf/4JXWmv+DIh5JRcDrgx6rIshZN6BFpuGPKI1ao2YPDlicqo9G
Y/iU/cAAavoYsMhjiClo8zpHuBRra/W0H33QxWQ3DBStAe2wwBUq+oINnQ3752a9
ONi3lBeWx899NjO8eNi6OLzYzSAY4Omm9JgbnORQEj/dW/KK68H0ie7k8NjQu2Zb
g5/5nk88yklKRfTP9fI6VIogUdouF9yCfXWpU0KvFzfwAPBhK/tWNUnAtXMfYkkw
IhUSzPjOiBmxI8p6YW12u9UnK7TRFEPVQXzEVefkiXDoEzaT0kBi0Hn+T4Wz96Yj
WZ6CCCcRGvDYV7CxPvGs8Jt5onemO3qSGlovKgkKN50s3NhUEXKb1kGh0XwM2yPh
nfiJ+Elm6gA/5qwY9uhpkPJwr07OE/xURmZPAcyi5keI7Nixd71QXpbQQ6vqXj6f
uuuwoheA4NSon9bgor5ydUo/GtZojCx4A7ANX73vfuej2yW6qcsSsbEvIOgsmYkT
UbpcRGTsgOZ8T5+itZUP3zmqb+o0NLQYkhiC2i6jx8I6PHfp+J7l0RKsnpx/Ma1V
D35SWLFJ6uE1PQZ5HQZIQq+jNy9QP4I4GEBYbhROxrAYBko5vnUIlLBoJEhtzX2g
c82HgsKrJ/4cTfaqMeitDsG/YLphGFbti8iXggGmrepdA37cP55QYZqtv6gj28Cu
BHfa+0PQqgFfOOHThgBfPt5zbw5rbHY34bsy9RfiIyD63eHuf6MYCp7QEkU5EPAW
K91XA8FwrYPXpdrB8Tih2qeKnuTMELT3xJHHFcPxGQU1lLW8/5ECoUBanbQNT3sk
/Aqup2whmqtGwbvaEzm6MRjp9o/VrHtZr/xhFF0gCdXFkLFJe6tGwQV+aCn21xus
1Ef9OlrKCGfNPwfJgcnRBspeKxfCbSP8PPRXUgH9SkajPHdE6JFLZmGSPZUuWhW1
temhmd4trZd3F4rXrAZMuxlv3Iia3rEfffQ90ZNdIgsNHXctjTJZ4hrTqm6WKihM
PjvMUEuOr2fFTW9JDCCY2IMJfH0p5DMjQwuKx6Y91+E086ZDNZtVQduR0LE5AeoI
MzrSyc8SSp5JDOv9YrO6roIQx4eCFuAarNUZYkL7sJMSi7g/RUjrKklCM1ytyk30
+dFO3U/3/3HJ7h+WC0zx11BApQjftICem8fMkz9gRpOOj1T6DWe++qywGXbqs0vk
zNeJoa+zaWkveycJRL232juW55cAXaq6n0wi6DXzkL3EUoVD56O2P9SZQbAB63i5
6T//yOF0Veu6w9PIYXDYvXw9EHOu/NNSpJmCHZMWN724fP+XcLaCUulz2ZG6jvMv
kYKhFmsnI/9qaMhsnkpS3Smk+C8lPV3Go8D53tSliiLIPIRZtAZ51kJZvlDESFgs
9W5AtdfSJoSt8EAODCZrjoni/sEaZMKaZDHhBTcmdeC4vaY6IAtsZsaM4L6xZwm3
LwzmRNfsf85+NPYaFuVWVJRETMEkHViY6VRtW7b75ZgxelZdC+SKdJfmBqr6grqq
wL0OAWlLILa2O47bL+26OSGYHocn0hoB6/GCHktxc4hfb+E1EwhTqydGmFpQmBXQ
BmiOcimbRi/EE3h8Qujuc/PBsITJZEkdci1C5xnydcVNMu5UdVCXbHQF3QIlufW2
6yusWceINo/z61z/dnYFQ88ZgHTBk342FhSN3/U6ZoX/0c8pmrJp3dFisstg0ELr
pG8ixQ4QeA///WkUlRi4dnAhh3B62Ft+ssKqVHxyuxy8uWncrlBjpd02Sc7Hoeq1
cgobrWxVpifzQCHtdvBzVpn0k17zgasqFTUR6uYOh73/GvVA+uzA2nRh7+WheJ5i
QmcBP1TD11yD7eI/2KSSrg==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
UVzSl7qeZL6jPoqzls8B5cxGfPzCfK+Y9AoAxzP07uCr6h+vUMk/i8JCnCDHjeSu
3qV8rhgLfPUhm5MkxiNd9wraaX03ri4QRTPiucyG/yjUpxJdAUCzlx+cpfCmQc6V
BtYsyaIEaGhQ+xtQ5L52qKjtrzryerqERl0HccIgXlyZbY6RaQxC7ikjmyYwC7Ui
KTjtRfwawBi96nnW2TBJw0wUTqPQ9Or1xPpgh0FcQC9xLbdzNiaWPVRh1T8QO/oC
32BYS20yHrehiYRCeHPV62vfJuAuQlXVatzirgX6Lypobfhv2GCuqOTPqfxaguNS
G7vCLFWtVicf8YmnRT1p/Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8864 )
`pragma protect data_block
pxMUWnT0DfBaiJpB0L+FxzRbrnJpxynuJ0KJQ5RCSn72KdjQrTb+VJGywhB5RY0Z
ThSAbSIHpFK/TrfBIOjR1HJyB7OG8sKQq2B3suGMixoiQ6/zE8gSpaAg20rYqLB2
5zrTD9dXaVPCobneO44Zb5Li/6mMYOqtSCvylybltpfB3VtdNmzKbpG3+O/Ofz1+
QIJ1bJ4Sej1q9m0gsglsHEFikXUPP2M9Klzi9qzwSuWSqxKjC+WN3AMueEN8miZq
oytwuVPagsQGrB7AimSU5f3SZaOjIO4ws5C5Oji9S4gBW9rEJa5wz99g0Dv01NHp
AojFhNuIY7PAXr304bzNTcWl77YLoZD6OxxoSysOoqATek6vFYLSwM3NvOilGS50
cTPfbJOd9ZFTwTktgHGbanYQmF5exjtfwv34GMlQn4IMbs8Z2VCUtHpbgjIgFNKy
/8kTc6QeR6pE79MozdC99hhl3k1SJrWQQR0Rg59UnKvQ77kOBxPeklcpIIi39Yom
IZIJOVTPKUQbJFVdYnQsz7be67OEb2i3ElQQ9AILjs9PfSsusp1VbmltYl8CY/v0
NWGGNC3LkAnY91wDXL2YDw/7MH+oapN0EfKaAVKe70RMdCGt3JJ1RKgGBVnmslE+
M12H4S11EUQxJFYNs7yDYvHyZS7gN+KzHtvYyHGJJBalNAQZhL3Pfjzb9Q8sslRc
CdTmNsp3zehcR+Rhd7J/xpQoORt9Zajn+69TXA4pdjO6/ffpgPKHyj+iQuAYYWy4
dZtC9zaa5BlXii3HIGh4LX3NYLw/7FAzkG1dsh5Y4IDjLhFfJzGINtHYgFPQjn/+
aTtDxXeYm9HNGVBSi7TZ5EFJglsLpHgQ5ws1DSNq/Rq6RoVS7QUYQoLCQRgOPUCs
/Xq07cSP84DTGduJUISX862VQQyP3/sVxYZcdS7/cpfFxjXSwFTiHroUgb27TKS4
DvAfslfb9qqLKBLYIdMNa1gGXhR0ZEzuFj1qCezOrCo98Pk3S4SXWBuuFMB4ZKJ/
0Imtaj7tfBmcxKfPp+XAmmua7ACyroviXuMBUmbeqSOANbwpKJ2dtVX+rWgwQJlE
IWRJnMaaG/uhjMrdjLMqHa0MbcIaDMYSaGR4zOEPpHaR3DtvV2ws8qUFV/ubv24Q
u32tPb8qdHqQeKgYLrlF3joRT25R/xNSUhv1lIy6D3UWRkfmOVOOdEEqPO6KnjFd
yBWsAMm6niomuO2ShRBjn+sFq8qe5g6C27L1WclVKqrsqcmi6xxS5n19unbvngFx
X0xm/NWK4tKyjnKF+SNzu3WRt6r2Mq+Ei+mj2QeVx3fCAXy1Ob3ifJt12ENvUtfm
SLEN/bfkR8SkvmEm5lohZi0arVx0ffV43J4CqfJ8WH7iF0b25JLvYC0F75tqslvl
NgjjMRzEZqfGQnq9mLtwIVxu7Qs5axfqVMmvYX2V6WO45jrHhhbSIUt5KJOSkwc/
KwUNY0ka+U51DU1ktloLz64/K++om7hu2GZoc3YhM0Gg2UF0aemcuJOwZUnkgQJK
wPeY6XhSPCXTVAwyNeBMjIq/V2SyntCPO+Z4exXuWUdkbZGo2ewotj6m+gWzYENI
QnEyqOODEGPIYUAjorOw59x3rEXgcUTepXoKPpWy7V/AHaOnnwnCFGaYty25BCh0
xmdFc8QMWvqjptWTUCItI5QhADZgwRz3N80mhKyXrCe26FNjwTbqmsd7mExdd0m4
t36ySrdLJVJkE6nWTk/VBNqgLpyw4KdlZvps8Rtr8ez6RkqMKZTCv1YlDvoXHRsw
bK8c7fQd/W65k7TYy8eeLzgqWD7OwG4lfKCjsKBdBUtcTlesQxhdGHUNfVac0OdB
BW4K7YWSGMd/nGGzizbYiy4il5BPD04AWBzlu4fv7ZFysiZZ3Roa79k4h79TfPQF
fZQ1JaMN94QxUCirQfejlBEgjVzCBz7+weC/evTuov0MDJo8iGFiPCm9YhBzhPHB
8LgfqQ2D9PyTtorD0JP+g/WcizcZFvILjp168rQvBNGyp7zbBzthmGhRRBMzXtTc
EZua7XdSW3b6kBC348KXtp3y09yCWToOd4P3usizzUM3efATGn24uSLrtt49HXCQ
FBZ7iI5B/QOO3RQl64aKcdt9GnfO+vhKKVXeWIL44Ff4JydOfxVllsFhh65VXAx6
gUBrqxXzYMDJziOnJFMzib8K1vVXYohpv+ACAzvoh3Bu+ONNvheGKW3PKbB/ITgw
uweY5w2ZQ+uWrj9GA/9/uBp8OSVINrutiWFGYFcQdnbGr0w/RZE5zQJHlJr6Rn3y
Sid+uXtvXN3oLDX8fesV6NdNGQC1LWMQFODo2+RjFaJgTNW2v8bXJwBAS94KGSZ3
epeOIN/zBLTy+r6DrBJJCOEHeJneFPbVU0hrl6CqHpvejnVio06PCkqiStaJclBo
KvTafBKv24A6ydKshAe3X7EpgTcvjMRhK2Z3lx+ze5zTsAzsrmfBcfLU+zWCgQen
vXqvdJpqPQazbxRssUYPbEL6eoozcA91s0lt4zdxDNOw7U4ZNCJP7y0OlGAR76Se
NbiL0q7YGn+Mx9/rtuQo5bbC/6wkfJyApmJYLjeLhlP7ih5vbN0p0ilO/FwXH7yb
x5yK309AhNGaM5vQRHjNLJ0ZFxVcC1zIygNTPDVr8GzvBoBi2AWCWX8zISysEVAK
dnJF3huWI9Z+gdLoFT5zmzb4Pyez4uZfoLYbhtQL18iYLLQs6cyt4Ru77Dk6HXFx
jThG7uPc+xcekFR5V7/54jl78d31GGur5zO93iVKTGa/7tJEpXCVbxBJa1pn515v
oEVv+u09fLPFjQu85NI5+S03x7ummM6XK5vwAH6/p7QrwZy04JkiMXtggpP8rkCf
fDhYNYdAp3c6nUPrieVf1hkA7gawyJoVqF+NxJUD/PgW9N3u5dD7GKyUsDtSGh0s
SxsyAcmaVmomuLALLVF2dRSv1oNgzqZ8VWa5r8BkZTLuBzaaV+rOhb2Zwq3JZ1/Y
iLtf/dj9fO9yLIZdF5f0f2hxhhioRX0K8+AB/0sIc4BMjGx+u3w3zDFMc+Gt3HoE
W4KFcgaFbrN59v9oeFOZK4fG2qzy17+ikPYOVJXuJvlLjQ435Y6TT2uShlAiaKwh
3OiMBmcQt+m5u3x4HkWhNUbyWw+bP7xAmTaXmjI4ubAY7IH5IeiXL2ArTxAfOtDO
utLpAvmmnjDOwLTzt9YBw/lF8tumFL31umlwCGuPQLdexWoacdeO0P6TOGOgmVmG
stDQWaR4IhJFfxKUE+d+2Sw2j6Uthxk2XmemglXURvKW/IhKWRfdeAkDcFXSwICk
LPeAuRSMeIb3SjY+RiBqNpU1W7Gi0Y8p2iJSrfouurlJPY021DPpm3gzWMvsbsFA
hgvN7QGItTE6Pq8+arRZZV38Hx0kdmWJ/BwAz2IHhDkmlkl1rt3Dwq6DsJ22Usl0
jie3D7vH7jhCUSu9W4/2DWGee1b0otYJjEppdcaq1GqoGKOSdKlKxp97DZXtKSFV
mjVrlRlTZJonRY5GfsYh3U+4ib236zfFwRnk3UaLZuQMgkO5UE24OlKrfMMK+ZyP
gTDVIf2u+dn0O5W7F0Kk/bI72i8qTI2VPO3ACcHRdmnPA5IhrtPaykPNqNbB6RyC
EOQ/s+MGNAHlt/iQL/Xwl8TOyl0edH+X+SK9corhibjrj/fa5hxiFfbv3oHUUuGe
eI2QoQXyJIvtd2lSe4zcU927BArBMkR+tjA57DkOKKakBeO9gUFnOkElHkvnYwVz
n27KupvbQOr1z8EF6UuQDtuOkgUwn+hZw8+hyFTXUKwofJNdc6shAJk3nOa1dmz3
lQADwxpJJFkV2H9MC3gIfBv07L6aL72rtZj0y+KfqJWdVVxn3j7GkJhsNQ0AAA+V
aD1j4ySd0J0oqqjeVN2ZJ9ROLMVa94vaLXoljBwUbgLqkzPexwMo50wqov2G4G1n
8SQyinb+s+EFAOTpVTefB5oSU1a3n/TmZzbozT389wWNn+YsxzVTCaDPevduOHCx
zlmhO+WY1DLwvd0CNMtYAClgVlJjc5LqXdNNrdGK6vLeB11FxGzgOONfqsJYs1Tq
t7Bx2D4jjvz7I1g1FOHCaIOUyKzPNqv0mdfW33DHfSkFuaHCoX4oGSD2CiQucoLQ
RQ48xTnuBfMG9Z+AcBD89FY9ZsG/WNOTFRm0wyEP8G8y7VsAQi2tkat7/HJy6uyw
cbezUoi/zLyBu0BJhNXyysCeT8P/9SKEo4K1lioLuYbJ4Zl2Am7C1e5b71zAbWvX
W4bc50Ij2uCYXILTKH7AymNV44ju4Qelrivgc/yqAsHXMIp1ZCOGZZIM/Nc/LqEm
79QE1E1RXeCAHm38rqGzKKssRZa/6I7chRAWGFIjI1YRwv9zHqllr8a0VEl5/vIX
6/NnvwZhf5JPYnj3H+3GqRZDvvp6D8N5fGiJX4pJ2vY8wQhN9ETLjoGG+nm8fG8g
KHd7Qd0qNLtldTlJ1CIWyQQ7vxcGWyIOWVVES8wfcpQhiYw1WbBcZjbCov1Q87+L
s/wOOCmfJr8so+Qa5dH/+1TL60B7r/w1kJAwxEP/5JVxpjc8NUKjiR8ZDGKfAV9H
hmGf6AOUEZWPnLEzNVA80NjBPzIJarjwJ2KMCfIlNeywVljUxcnWs01e8jhNxQFx
72GPx1tQRXVOyCFTr7VfLzyyE7/ZlALmLGG/dcQ9TiPaGAcmkbT7sSAAigE54N3O
QsSQBmj8oLVsQiTnankZlJRhDfwoqFxuEZ9ma8eeag/d55Hzduhxl3fYSHoqIqfr
z28+dNJYgtV3m+QLWHCwOahl4qdTOMANGNczTX+/JD4It/BfIlcyYCBAaARCejhH
M/IcVTJr2cji43nmaSpZ307StZscYlUFFt58an+Z0XxUu95uh9wZRoFAfJIDm+5B
Eyds0l0UyiUjJHrJItrNHZXLG6Z8KccWQuDoqlZI8iNqLV33dJpot1tKb1xqqZ92
X2SNjeyzeH8rpmKIEbI1fuhoiAgg9bh9uptYmvfN0NLFsoRz9MXnTOdqNEmUb2sS
1aYi8oPuy91WW7UCpde3LGMUDE9bTpT0JOGzXHD67OrB7/rQSWSGEANWgjrEXx5L
m9jerLsWPm81TqyqiRZ40vsd0YJ8EaK8jXqZU3shBG8jsZSuHTNIK4wA4LUt4UE/
Zi7Q7vTYLpEpJ4oHExCByDMJEnKk16fxEB2+sa6v3Rlg2X4ZsIPqD9p3zqhymz7n
Xcrkl+f/gpPJsiXJHOdT+j4AJhbBSfBrLGSEFdfrRGRC3CeIGmzvuRYivygEFyHp
SMGMCzZS4ZZVP6EGb+R5rs5cZQC9GUB4ByLR6cYpasSldihQ7tpiN6wksCZEGtFF
68+XcoLbbZRfl839bu5s9puZATNv81vOcu8xV94PrMozR3QIrRakr2tfK1YblLvB
pCqGUNsFqRIeBX0mDX5Kp5eviAr9M/PY6Y4SaYJsoE7AuOEQak7wuz4bzOzinLZL
IP6CXza4vk01EZnCImf1Z0WueYgtsIl9Cfl5vbtBvzLh06llTfW8Xpw+eS1VmwAZ
p6tpLRDadQmHKjnh0jyNG4BzKkbQppdS5PMbNPgURnPnwXMeZ9r0CJQIYgpPOhjy
5+qfRGERXdgkYpiGvJZ7MdxGi+m2sZYRymXuDJTYqsZcpoNVhKQTLAWEgplbi9S7
+3QaaWlYobIV0JxFccJM50VBAHJEJhrucSqEQnxMT2iRZKk9IDj0JDntsdF1tv+D
z0ptAa3y+otamUDgVepBKySmilIiu0qgAXPiR6ksYyOKfUNF/XgpfWefjNlqYT7T
2Bjk+RjWWwwf7Wy/V440KqoxJD0777pqE/czqIRuX4n/zspFS9Sxv2gTTqu6u0oy
9u5Z6yQpaVZclTT1nPQ3aOenRSH0FRKMDz78m2X6itnJL1zJvXSVcNXaOXfzVpaf
MPgTSmqbEHEoMKuTfWbG/a3AEYmyzE/nIOWJxEeM5vKZV17B+Ne8G9zJ2wEuU2nN
bGEe05VjGvdnCtU/VfVDRY3anv7sQIEOjBDIu88sowbtrKPhEBFdnJOQLcY8P5Da
7eL5b563xcyk5nyN9iLp/8LOS5WmvgwCnR0bnI5GiLTy2Ryd1goDF9xZdoTeJeDp
PLkhLV48twNy65J5n+GOUa2hrZ1LPHQ6GGbdDiTQ6DA0oT36Lo1qvvsK8PGfF/Bg
QWfafy1mGNjzS7JcpsdISrGkXOxXJrhJGuUnX89EwjfeQt7gpevCOMh85adIyWJZ
WE5LNBqshYe9gCK3lFQEgG8ElipCjkuHyaND+l7ls23BGlS/rgk39anNQdqaOYZP
4HRy+qreHZ3mP8CvmvQJiGZwwMwlM0oNanz6lyGi18+llljFCpSJTfyC/dBMx2Rm
ECKUI5WksmigZap7gNuwgkheRisbBcwZ2Qxamwdaqy/r/tV+fdEq+Z9hLUE0zbSD
UUarCo+nIFQr4Wk7iPL3BSUM/mJxuuuGOSBi+sJSCyvzJuNUWGk49hF/HydOWJRn
FJsI7fbnDVDlFZz3BfJOIdoLUN/LrYOTBqQoqvmxzyL0P+6HJJEIGXYm7X86lkPj
Qwv07ATiB2Fng/vohtYD4QLKMixKWNIO31LbnfbvBxwpVl6z1dx9OGKFeffs7wMN
tQe03RkMMI15qIFNf56TbMrIHqCyUkOsBoFFTxGyUGtjnlsLnsMg5Cyuo+oK9Dcm
VNZoW0/CpXgRZmS71RL68UAiQ+wNd4Su4IPW0vdhVme/mLuzMzDlRtZd1GM3tz3Q
uo4+rPrMwWwz4snIA4NGrQazBjNBS+SWMpIPe56kMpdntOCxhdcC53hY+Q6Iszqs
YQ8ka3Jle2eh/HQos5zRbazFLNW/V7T4WyPuU3kuGLZnuUU+f4ok2cBetULYjhd8
bcO4R5tqnLw+y+E+vyAlc9qtqgYZWVx/5BohKry1A8g9WD8Dnlt8izHvVGJglIAG
CXU8GfbXt5cKDtGddKtZ5EviXbo1zhPxLu5LIO9dE6LAEZPN+OkpC4c3hfPaFZ0A
tLf55qk4u7UlnF+t0t1knBGgHq5cSxdNb1YvhbyNQPNAYaIYGO+tQQUMrYQP52ea
uYMLaQuwpnFt13nS7IQYqHXnCt34DZBf1cMO8bejBr97F1qJPCO+SOBA+cvxoUHN
vPUoLqO3XWve1c8ROyXMcWFn4DBukmw8LXrtmg2pnTlUkfSgmwws1YzpRt3ieE9b
bRBh07koZmD2zfg8SYJPDs3blVZgoLfg58IM/2+vy7aLgEYRDyoDuM8eAhsl3OSu
pUSbHtfP+f1gFO1uxZNDyJDilAdZ3HhDjPRGkmjI+BBp8l9OECAE93+bmZ907rB+
RSxaA4ytycfjA9vQHQpxrWc5Fjgol7dmF4PcMQeaUmd8CNx86UL1/MtOUup/25s7
jI0h3J0ccJ2N9sXCq6lvZjHF5Ttk+v08gVHaEU5N3DQzb8H2UkGxpedkxja1H6w7
HDf6cu612zTNJvHW8GkLuksp1hNCdER8u8brjZCVcQglo3DIcs9/GbN3GiLA7BBs
1kb1ZtiALT8T40dq/o+W3WqIioLHLnNUnIYs2ohh/q5pTY9npdQde/8Dqqx3Gala
CGi3v7+gIy1HkTtVZmFAMSHyadcLF45mSNyIAuLoxyhkD46BgypyknrWbNPBcHj4
8bYNOEvMvY0BpsoFs+A5Y2teMs/RHKx7ofG0ea/XtLfYR8nf2BMICIl33BAD0Qwb
Dnn3d4iXybrJajI5Vni6nOBv87CD88HWZaukgOGSE3d5BG4F0rKuPrWtO6A2S6D2
h196WOM12iXGctT79HZf3FwOgRBVbY/AsQ2AM8ERgTo6pL1IHn7OXN1K9rqTSX30
z+BwpVODxbAqQb01lzfV2ksFuVNKrgyYpfaZfDpzZWXLROjNVDz9fvyANF321e4x
ivRE7n2U4PqvHm8V2gXygBmuanvxcZvAU+bpE44khjdYHNt5RDIzvQmj5Jkpbiup
Q+U5lrMeC9IRTgh8/pQeKXWf6ko+6aKf54H7UzxZGnL5mAwrlNja7Sud726r8REA
Q5YgM05kZRFNLaRGJYSl3GIgSlIbr3mtwnIC8YPjMzdroBZydi4P5ByhhKMhYEI5
zVBDbHVEpmY6cl4TKxbPMWL7M9t6gSc3sAJ9meX3mzOcp/Kl4yZqM7J8fANkX0Rv
D4WGhiCwykJ1LrebiT5bzMorJtOZ9htq2z7msFhhXog3ohyrgTjIZ76aOMT7RHf8
w1LLHadmH/A46+HWRnvgWOdW0AwWQtFt7xiw47l3Fx3D+0XrEU/XMUt1SATf3aiI
tUaq4/nprtW58eJRqkfWMJREHMWUWlm1SzWbyYtvNGFMosyyzvT5LBpGQQbcVtko
8lPdL5ZB7SmfFlZwIZddSDefNdAffavTxbdal0LaWO3s9Sy2j0n5EU/E8gKT9DX+
Uxk7IvmR5kmQtJmXPDYXg3Z0Xq3Bb5ebCQpBYKd4emQYCfYhEVdOjoN4kuMHMphE
g1Q/s0PqZiQdBGhyrHLmiZC7oblJZH+A1EHF6PdqIvI1UP3+7SKV7+O1pa14yqL2
g5o6XWM2EqQdPmPWRORq6vGfbfAKup0UtMhOTRmkATuNA0oR1I03YvoMiOZO4Eaa
jxVsmE7bFQQP2uiHENEN36vJA65WIIs/h3/g5rvyGfM/bVw+8rjoMHQv+si7smZK
A9ehEfRbOvmA1kii6Ocl/NU8Wm0lgq2IuCMXWgfocQqIgUKo8Vj1sYA4wefvGgGV
lqaN5OssVC4qv5DSU3Mxa09gzL6Sgu66ZcLJ1T1GzxtaDEjdLJvmU6gdgea3ZBvI
hg0av8OJvFKpzyV2cDwVRjHBExTfVxEWbs0sw54gu9Nk6Se3Grj4SbzoI+SFB0Qj
f10e1MfDaqSWIznoeWPck8PXQOSkEvlBgyfvh94vpy0SdM1b/uatYFX708g7F8lI
4LfhE56NmeKe+de+UiWLoTw34u3weNh1XsuOZ7tCpdHYJgtmvzdGR2YH08IVO+Ur
D3J+TjgZdxTBW0UHb5/NIkWeOuQGhuCaC8f6O2B9CoZ5/UWSBb6H9YW5RRbWEBra
Nv/3pXXIYvqtlTMt4CcBmWGMut6PDgXkJmXCuYihoc+6dJJNp0rEgJvFLoHlVkcE
mnZsUyuz+2EJJczHp2LSgkjMF2tP7vdLzCUhOt8MlaOjraQY9OIdrP+OihdBXPG9
cS0C5ucFfcMAyrHMS90gq6HaYDgC3bjOEAGB6NeZ49gbZ/GXU1dsVyedU0rx3fdK
BTiOf7jBx6752L4TD9p4hVx5o2V4JclZecff7OLoYcaS3trikao37ADWAT/OFhR6
175W10Bp8+BfXHig6P3GDs9NDqFuWBaYKNh62OBWKa53iI903FvClHMpfxmEZA4j
SvzBdQwsGppUia573JePxw2jJZC39xL5aEF+epTRU+UdeKGpxFKVn2I3ycxHuSqJ
cFM8sy49g62j8W7FkjQK8WvBSmFwOaICOYFxP63ew0JCVOrt3ESqayxMCtRWxMuH
THbU2ehnEGKX82I2O/qFTl7wgRuU1yefDzt7becKmq2ZG1+bL29EkINjum+A1Dg+
Jmgb0yyXDmYHivfB2KtfBWDFw9GAAg5Lk6RDQf2975kkS1sGKuU0CPEZCwA8BIXD
gvF147Sh9IwWPsP4saXFhDNhNouHf2yLlvyTB0+jxFhugVuCjxv7QUWF4VT0ws8b
N9GpesznH5v45MBpFpmnMZxnnLcLzQF+VYayJWUvLYPyxGPGo55unE33lcm2TaCE
baZmJ0PzDaM5E7rac2aX6T+rQ3zewrTS+8WIU0C9Z0w2gEahwKoXMqR1eDUUVBuP
pOHiTIN7c+T54ckqk0pM3QDMkr29zxTo83S3B2PBaeJsSNZoWZ2whOSOf2h/k9i2
VSo7aEjI4mzROxc/uXLTw6EJ+b9+60uwwFkiq+R/Jhjsc+jpsfFo+U0F57Klv3/p
gkrDjPqzOfEf+HZqUmYjrUShWd71HknKs7w2ebj1/wi0M6jd20ZUGyS1CyVwMYsZ
CyUGEh+wm1vdajjvW6c/ylQY0IN2IVov1n3/oG+CzBmm+STi31XU0hUTk3ZeLobb
PPSOyMvXdBIp8yw1IK8oH0Knpd8FdBff9FP4gs0UmWT+ATjcCrq6jG8yG7FDYoNi
p9cqt0sck3ZGWWa+1sVCB1KGY8TOMWKwvjkFRBnIlJ7sDd4lDbr+qoveBA26SYrq
ZRb9bm65iA8JZOlgI4I6mF4QBdsRTqeDS1TIYO2lQff3AfN+6E5uSCW+VYjA497P
ppqzXiheqbZ8SItxFyuJVow4Xhu+Hb1cIUbX9XzbSwN5Iiu4KUChKcdmcp8116rB
yzDnL4dHLPeckNldZBH4ms+v1Fw2U+vm+wRJ2UJLZdHqnedFMKo2Vxwy4UrPcgfP
w7lTXx8DAduSyp3WN9yQZCJnw+xkVlxVJ6BAp+1bgf7MEArJ2aAGjB6ZMyJaOTaV
sHgehMefGlLrCi9Dclqf7YxzJGaOFKno+WtCTFfIf9a1olbNGp5jQciSGwitW6dQ
OQ98KSRRtJ+rNODVDOdQqyzyiRLXAoLrkedF5lgYZIFwWW7BtkjqjwT+Gv5+5+f3
18jdOnqYr3OXKV2RJo4YEsSqV9rpdgUhYsvx9IuxGQdyW1JNyeYBISNrP/Ru3P0b
7rwvn4BSr3Rj2XcI2ssKd65HwJ3PqKNxKn1sEhLZAeBQ3XDtlRSeX13xwaonQbzs
GtIR7kfkqmqJYYR3asDmWaMf+HL1rmx+UoC9hBcaUdOs82Ve0mXrp+PVlaQ2kbln
Ui7MoRnT5VMT6KpWI/iaCFQGufxNq8xazU9mUhzig23bwxv2HJvhRCdMGOVPzVHF
GFxmBctJSyRQH5tj47d2tWzGP54bMD7kj1kI+rA7PJ+KmMIHLhJJ1+duXuFxdTdL
zO1PpZS7PDIoOf973OmyyTBmjlXBxNc4M+hAmRVsA2n7Bv32B/QeK0FE80GFD204
oTV0AUGaSJCMMLebDJfQHwR/CCsrHeq4ykxHakP9DoKqI6CFsONzFsiQnep8CdSm
TDnFLqTMB9x/THOkem9qKutT4IAIJkah78IuH8x3jifor5oSzMTK5sXl2NzRA1kx
IoDHWX9AuPYeLFx/g1U77JkN8udLVPaFfFOY5IUrIapTxg4Fw6tyP7KeMR8Xel1A
21DtaIqTpp9KoCDKFXYD0yYVbT6ZVHvJ5/Qo5qxIa3ew0T44iE0ni761GJxuZHF3
A/Hx1vFSwEWjithCZOmjAZF8UCGCmt6lsCK+5NW06xa5PmUtNOVathGRpWEthWJU
41qWm4EnMBJthWYFVsyNVKeFgcfqJxOBu3vvyJq9tPrScFiwDaaYlSMgoKGMNBoJ
AsysifmxEZzYNszacH3nyj9EJ+cwHPqAhqwzKuTtMsi1JsDNKqs3TI07OpnEPaJi
i/jyWgYfKtOBpwxRN1SGqy6KQz7TbKsVNXuY5ptZutrkZYK8TZ92XthRolVjvAxf
PhAsRucwSB/xDPr0fObCVbxpzVNC/k+b+ldz1sIde6NMT+gKok79YJ0jdxB0KIld
OWwfsBPQY0DsqNICkIMxyFNbjif5S1IFNNBjLc8U5b5787SSNPhRaMmapAib8ir+
CS8q1/OLz7+npwsvM3d3lMkca9RZu+nAjoSmQ1U77eIZJAVjS7cX/+edvuBBGD1N
Vmn+E3qjUtWw5QRFW6hv7n8n9Zfq2kbE6fX1hnKvmFu+vg14D0VAhDe6ni5JJSjN
6CsSzPWWrrMEm6JvMq6nCEtoZbRniLa1T0zUyiar++s=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Peq9FXII6CY3hdaN990YtAZjASbgItnMSR8a2Q4vvRHxpMgD/SBp59ZrSpSO2xot
j4k7jM9kzySMA4sLVkdzetG9r2444eu6/pHaRlapyi/OXx07DjKcBwEiXK3R6LE3
SroNc/3NxPP4eT7ptGtHK71BMfytKk9ARl7uv3MWcnbzL3oOCEJwh1/GQ6C8g57n
PCONCKqNCGyF2v8riQQgSJIM6umg7QoVnhCREG7EC/2yZXtLaZtoUhcLdERa18DY
JExk0l2J3kG4ibX5/55RFlWHTo/9wg6XUk1OjGvV4UnAqOf/MXEKFb2ePt73sdiu
Pm/J0u8C0ruflfX4iGpD4A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6272 )
`pragma protect data_block
6DobpmREn9X0q9poJthtGDq5IRc6QXSYaPEaSkdvlQ0gIAMCmviVktUIwhSpFmGG
cq7wmENh1/n8GXO23TQRRuPjzBfF3Tun/1s7+dOvhkfZLp8Ur2nxRcbU8dPMg+Jz
B8K/iuk9mAJ+i0YkD3OyuL3YbeSTQLmrFbAOJqMgV5xi2oyc7c16USVlAiFwT1yC
hLjdbz5NK/BeSDBZde3a5Czus01Q+awOeyw8dyfPa6kMswiq/LqkFE+BDUirMENK
EfCrYi8Zj1VvJIfanMfAiS5xBBsatDoWZCgNqxxUD9Y8FmG0lkYx3vVjRM+/5XZ9
7RPvPAMH6ovex8AC66zIkfq1lMGr7wLcVPJIQuxZxa3L48lXTc7lyZ+ghEFQ2ZW3
ns6EFenYQaHpprrIDFbDDC60xjcVk3VFRmBZ7E9KcHOyVyNSoNFvm1rmeLGkrHm/
zIYxb3vGI9ruJmLiv5IogFGkInOTzZjPZLHWHZk5pqefqIgA8b3pS+Lh+Ma9/Aqn
tuhx61iMld3a6L+kGl22ZAaBkk2cdieMpcxn2Q3WWmQvWe5sWOIac/uc2xKGSKSh
st2EpWF1M5Gs4wLyME3XJlFfEd3sWUB/yRH9jiDijSX3TvDcpl089/mOsbk2Q/FO
rW7PhG42enWAOzj1dcNvtimmjQ4OHIQxP6YlGxXhJeoc6DUO76NL8dVZYtmoNSf4
ducUg8bq84SWiy5j+a1otIQHpAhE0996V28sBjNc5pHN+04296ZKonLur9JOyiQT
a03u8zHiGE3PG1T3Mnwj7E36nqds3uwbQAKga2+ic48U43TJI/rfExaMfGx4a6bt
rBZ3CErAsNR2lRPPnjtFvNr/aLn8cuk/MtwJq6Zz2Wau8SHGVby7//BLNiAJkNbq
PvYBp4MFFlHl31GcRc2yorhyjs+Z+KGjBG3GYyNoSyF9N/rykIOBG8rgfNT32mpS
QzHSiW0t7mLUQkHnxNllTalrhZb40bz2QzaICt9q0BSa0EUY0xXsnCZb7d5zIW9s
DF89Eoq2+SmnbRVmy3rsiqw6Q/j28IVwT+/k2zQuixIkbhwDYyGYWo/7fzpzEjr1
XBhm1BXxIL/Yq/TQIgcw7/LowEIj7WJV4fLeyFcr7AEgT8WiBWE0kBvIo6H2oewM
M4Df8+rjWGBD8+ca6hHTSf+F40eeYJjN6q0kpt/EXMiwtpZo1mQB8tl/tet/9PY2
UrbWCt9mL/o23Rok/VdLY8fzsghEVj7Ygr0OwUnyySzD6uBENrTfnIXu3acxuQ5U
dHd5npWQOYjUdufPzR2lGCFqY47E0gFznC03IawDM1mrUu9IZLFvOXpM0909cK+X
RBwYKfEENsCSBbteoCBKhEkEavJLrFU+p27bqy7u7QMkUskWmPXdzXb3Q1YGTpbP
Ek4MDxMeZzREENsYqYDkE0K1lZbw/7EQrR+iEuit4Sa+VorDWVtZk5Qk7YOkIS1L
QHphYiSkLKcqorW1tmS5r04AzdPk9u2ocXcFanxLkYmB+aOIYuUZAaFN2YNKcOm/
vkNb4DYqnNV1KljfsHrcvCka0lMjOylUaTbpeePvP6/1/dfZwYL7Qt/72kNLpETk
K46gpwMOLk1fvDNJTBC7jXUKLfoPaDvcKxaRr8j8p8RmWFQe3Y0t6SKlfbSCMGdM
jcgOXbeWOXbWza6WiiLDy/q+xcxAwAewWxByeBp3ujBh7cL31osAa9mHGp44J+eB
Gy8NEOs9CKuLL7IjygDW9uConxnWLcDIeZFs+3ygRjncjUUq1ZSWQMm4TbJW7Zcg
be2uaLtGYgBsJpSJZUA+B7BisnMEjixjmmzNHYMRi1vve1MBWo0bzJ0TDLLbVM/2
h03zQM8vFHyTOCsGKXSTra82+5CoZgX3pvB/TAkBj7OqbI9JA3aUCeR9T60B64fJ
XTdnv1NYC9O+PnjqLoM2GwAv27nSs9ZJzCjUIbkxuXuUOrScMmuh3r6l0E8Q3QUk
9bnpzwqOQwJ3n3dNwUcN51OFelnf+Bo0gd2yQS5dFeHueNEABAC+GXSWuHJzFhmj
/Mzkuvq2MlCHy/CPwoSkJD8GLR+dRVNIFJeF+T5wcmgpNQ1Sl/qOmVtExxvjdW/a
+2xqN6dx/KJLe5BgX1UZPauwDwVAmuSoSlpPvtv5gI9ukkr9wQxRk78RM4cd9X9s
WH5PxPQ0BRsETrwyQ4VK1LzQOGoi5KSZnq+aSYl/d0YWv7Z3TAw+4HlnPsVsvBeL
RPTRpEWnMg4x/jiuhLVqZ2ION2IG6+a7kYLlhzZlPPv21bNQoi1PwymsDD/ERHK+
RAAlH0XMlwGCSb3n162sGxXWnF02p/3nCTns6sgzz4WKbP66tmjYVskMEPr9U5vk
AmeV/JMiOhEHOqtKL5BhIR9of3LTiCp4YGHzsgK2TaKlH5LB4KDve9FH21JotfEm
2k5Mr24/j8XRh9Bs2LKJnOzfV9rRjp2oRsBZTsRYPwfMETx+mH6I5JvdbASyNbcH
YZnClKxd0Z4boDgINhtpHmqXqLcblrX0g5ivqTm+GUWIMxe4YWvQ0hzicU5EqIxB
KlBakDImvv4DKaKRRf3bHMMDDVPAbPy+eJYv5/fFic5E97aBaGNFLME3FVx9hxKm
KGtm7SRugPl6e7Inqc27RdC2I3OMamnryFEPGOqbbJipfMOvizoTZrEi0AB/5H3E
ErbkA9QcxYU81Ru4vWnDRLr814PCcfeEwT7Fb1GA2+yfQbUb//DKotw/G35GULs4
+tafMz7QzkcqjqJwnGDkK1Z49vjK7zXjwAu8yif9+gsvgozluwQmsg801O3SbZCT
8rlqwJX/24h+v13hE8XG1Bwoc6E31xSERK9qYvAn14goinOwxkzt+mht+HLArE8M
jRchAsPNEndcD1VdivQ3fcio0AauMyOc4IzeMHQffUmwQyXBHJV6UAcRNVf18HJk
3SIyfGMcOy5iYQcwst1cdVxpeIaqCa6y+K5Jgi9ZZt2XBCL+4qh7A9QBGvjGDzTS
EBJKTXsbwZpOdNgShueNANSn+Oo5hK2yznjwf3QteYscXQGx4Lx3KYnEBGYbhGhf
Be3zHccnyWiBWHsNaOL1whe0kVTjXQAvoq6289/jMyEoo4mKIxoUkU+siUIucxyn
re1pO6z+8jOXf1WoVljGLNSWkXP5iQq0FtquMxTzIaWy6YKluxipb68ggNc5yuoV
vzbLVTVDj5ozw4KRtJuC4Nm9XKG0laww9a6rfUR8HvBCGCArd1WoobvkFsGd3RFF
JuAuhXHijMRSeKOvbYASl7BrfhUbsB1c3mSI3dUQE/2xbD58NeqzicQLuqdG9ISj
CKOy/mXyfb80ptqBCqUF657mc/gJdQdxDQBkX8fETt9LkFvqMlu05MysnkeqaaqL
q5v1CzewJ9Bm7j6j7niFkklhqpMwasqaG2EGtpwSN+ijdUCMkR0WNjzG4q4SIJ7G
AeY9UHx7KVVCQVnpdwkox2q5V5JSqQowyyXLLZcNS3J25Djz7Ym5gui+rZ9z/eEk
1HNoyJgnixyw8yKSFtVAIGTzOC6XKygasRhpqFEmPy27wESpeI2CZQwwjrv0MOez
m2QKdi/wEGAYQTzthGNDRG5li13dtIi0HcB2cweTf4ICFW0yuB2IGBiVgI7XiTq4
LAnfYN04Fx5oBEJfU4IrLyfHhsv00lbaQ+BAmQOpmJzim1Ktc1gDm5LzhA5cBMU/
fxBRlFat2F4jkIRpBda8IV50NR/lXwzn6WdK7GVfXApHuOMQMR29n3+CaK7zN/FH
HO4mY+Uvxrtj2FT6ItCEqDmDmgzBWq0Ub/F9FZM3FZ/Bey+W2Yk9nOAy/sZP9Yku
Zl1eoWfhReP50fDXAUot/mGEk+rrMp1tN46/beVcu4Ir2owfrV2RAfKKhywaxIcV
HNL6frXrGQ22t/W9ydvZt9CpGc6cNknI8j3iKQY112QomBWShh22/ji5NVqvBzzU
cYjUqVAPbdlbOaZvf4LJzaVRz2AuVBXDoZ4o4pH2EelgyShWbjqopc5wsnYmERGT
T1NwZ6zXHnva6jIePDBbFMRlHHMeCSkvSGy0wOwChBL3tMl7tzcdM87o7X9E0KcP
3UkDuJuAeVd2psrGLJ+uqLnO1VIwXFu169aDkGUrnYJMwV/lmUSyXRO1gzBBhIS+
BUuexOrNWSspnuvxe7FOrn2EkK5mt4HowrBy05MlbL9u3L8HvXzfeUQ+1Ca4GGIG
OgNPaRmDpvXyj7XSfAjymIllGDxd+7ieqvVwlqzn3w2BYa2aXSoctBjB3W2RSgZY
wSqQhHNd3t1SKmAGAE8onRNcsPSikemuhyWIxCj3vpBQR98J4lHt271zN9ymL4e8
gsuX4BO9EU4ZY/Ba2uel4WaSuKJaIufSLvysWLVrzXcPIysTw05EvZH0iHet0+m6
eVkCkAcgjhl1wc+7kTIwXcWwkAqBeyzn1iiqgAu6JC05sKmkV36CloXEz86C7orp
5iaUcMzS8K9shxJJci5gz8fflRDuFglzFBW2Xl1eaGrmkmZXQisxOh+LQGNG5SOa
/rjn158lm5EhdOULc6li2HVccp7SyYvARhyakfupUkRn8wHoTr0yJr3A4iGZ22fe
ZcEB1LT4+IKSHrw68vkaYBB9VWpNiZQ4W9qQZiZgNAY+F5AGZoxi1KxmLmc60a/Z
+mIjl6dhKq8/mK525fSI8eDRnkEl2wsgToJiVrXZSlGh51HojUV2/ibVg9oMCrAC
i7Mmaa9FHCtcqlvof35jjjN9/9GCwsshrnAuI8AlJ6k1FcJ3XorSSmUr1SfU5/W4
6jZEf+07dvyYeKAhnkYnYaF6JAUPJHewLN4EUVn81IrOqeRqNqM+2ZpbF2Ah4gDz
gGaHgH/9nkU7dFKt292eUh8Rz6G+uqeGpQ/oyzbWCzmaEBRgpxVF2JoR5e5nOyta
x3tCcHCMkWuwUak44MA+q+Xq6SWMdc1id4uISwXNNLBy1Uiig25v85JZBX5103U6
+hZzvmoYr7mgOVWpXqQR78Wy7chQzXTcNC/n36kSQ8gVeqVlo7uT6wjAPkJv9hCf
d0IsLswvqobqCQT4E1TUDQ11QTE0Jgm/M/yApXHpgptR5RvmG8g/PD3/w3vqkxHN
E4pMDjKvy3Ovt0mIRNP1+4GzRUAyDuSwSQFZ/PoTDsF/uufzpMZ05JkH08cJAVlo
oxDvHBdFlpmPD7QCmLMJY6/F5MGiNmZ2/pctwgRzCUwXV8k3hUf10//ANoS7N7hW
wcFqa8FbFeO/APgkdqz5sKX59lGzLfbFk69yJcTsqwpgVbZYcR8Uv0h6d2GOIwV4
VbZuurnxBKhRIr4PKMEaC7drD1OdZQ0FFPEmsebN+rRUdTuvaDQNkOphgawu9Xd4
zV7moJWyBx5c+zt3XbXVGbzxxjpnMpz7CMJq16R/euGl1eFv/9LngDU+9Msi0FCB
/2oyQIES3AvDM3bd69pjAaL2ljId7unyTJmCQ3SvsfETYVaiOHjxW5+kMhzOK/Da
AstCqE1T1zQPwT+7+EgPC4DzCrBV6Wgv2Hr4MoWZsbPvQLjDPYOmdph8uVUeu1R3
Rzap+c96nBS8XMBh5aMEGMi2nnYijM4jaIytmoDV539crmgZHLOFP8PGuE0e7jNU
htSfXkwLiBfyVjlCrGmGaX6nczGIxiDETZ5nhWY/S7s76euQLzW20H7zxrBZuclp
h262n4Uln9gD8BXxqcAMG466kOgkVReITsjIE0f5u8J8eS4dTMxZWMH2WyOLTZZR
KMmNSUyhiAYAnNloGst1ln+4yRbXtwiI3NDq7KqLMTi+dNeh54+mvCwvc5nACVjC
sF1xWyVGoCJq7MScQ3GyqU1LwYIVt6Bi++KRpIs3rSDMX7USVPMioHtBniZoUNsE
+AlXJdR6DFmZwej8SNQlb/ozXz2YuFtch2Uqlr0DZWxUVPEFWr2sP6wc6KuqzBUI
N9qppdGaiyErpOJ9nVLgfmVlYKGkskSFZkK2ruYwL62+X+tTFSp3VoOMWiVoIRjd
ofULXN6rWAeMnpj+C0fPSzD7zNGk9TZDzWjj+E7kHa4o6o+KHOVQOvwAKynFnpQw
sZ67VRycdl8fpHl/mHNUSurs3j7c2e7dXGgq3LextRhCTZyNlQbRqcxds+5IKYt2
rXA/ASrj7510hrXH0ldn/LsxOZ4aW1bqZzv9rEtOzgzS+WQJ3RiQmNBNnuaI02ME
rdrJIHo/HYdIZQe2FYaeayyPwXhL57f0aH15QJ1oTySxUPTCNOzdnQ1mk/eGwS/q
ksb/UJn7xakN3WW+3gyjdaz3jaqmUdAvxoxjPx1L5OJrkmSry29pbuLEFXE+Jbcj
KlkzkqI1ZSoZz/0azqig3IFqzzgnJW4JqeO+DOoyjLVj0fJX/zO0/UC9QyEziWbc
Hc8uKSzHg6mnCg9453UFSGMdTR3UdK8P7WJzbrf/nDwPIS5PjXtSNnUpqx02AcbO
2RkAjr9kA/CUrOGTyEWaKIfXOnGleFKA7Z+qCuoo2CnQktPpJ26043bit+BWxy44
n2DSS3iJrFl0w3kTzRSSGlUOvGZ+QknRxDJdmd9GgU0u6gsXwTfemGWSAzfg0cq/
8CzCmYOtnpfjMA/GA0jiyqgSbi/qtNU8LBlYSz8qEU4zDPUXi6Al9x+UofS+lgmm
NpUf8zPXhRPzAOdFhRDcRfydvQKwZcMGYSeJ59t52eP0oGl9z0ctBqJzT8ZCzVjq
GrYGqOqpFr0vtLoQDM1hTm83FkJq2t9ZdWJ75Mg4O357LUNvtAeOQNvPzJCfiCbJ
hkGQ+PAQ6V3nQQ+7ndOUFXnJeovatZwLURZHJd1Z2KvKlj1yts/OhUvk6y7mpi29
O1umjG67qdLLduiUY/qZ2luRY5fTkap4uOf/eq/xARDj7EKjsmyysUfc2LHfiH7p
T/lN6P7kIlBN33Mmw/cKbfqjyOHDNgtX9KxCfu0WHv1UUBuzErdvoGz8FEzc/IFp
nQOoTJEnf8OwX46oO5BTQpNnigma2t1/eygA2ayjNULDYSWg/+14lJGLA/NYI69y
t2PgOjScpNR/SV+n6X5DYLuRHlf/TJ3dFu2T1p49/Gtm8eJZNZv6TfocLKj+JPlJ
npVQ+CAcH2T8VF0sGCsYSyHFMEfYvvI+LOGKxqSV01/w3+lI2VdSCgCmBln/ru/D
Ikd+vxkcjFrGyd4YqZ2LrUbiBGlU04wC9tjOLECI9SjeFRxd7hcAWH0F0rI6O47I
02Yj8mMitPoJyoybijUWGD7oEadyTa4k5ZDk4txjAt6nfa5ZIdD+hTnaof8Y4fmO
NOWUlHNQEs7oQcKiiQAX8S2WSTqkJD+S78nR5ikq4yoTCVb4EYipow/jZfp3mEAo
2BIKkx/Jn9elUO78ZDGfa0gs2MR+fc01GP9FAn51/asm3xGkj1YwNQiliPYXCHTI
6z7ZdE8Yksl6qmBhwWrXXLsR80B/fcVGVdtolvAA0wcBkFjmv9kaHcWniNL4gC40
6NQDCsUyHgpHFEa5y2Yix+Xew8XVwh2Z4nRXwik5ItgZhrBM7qupvbDVdDzP26HU
yhyQp96/3MxT27RwT2R+R8XYBi7NtRdNjg4SXzv8EgYvm7NW17Xipjx/TUvNH2lf
H5rxP17DnwXXFwqYRalT+R0nKp7bmXrPcCe+66zES3S7RDpKoBtRomN9T/VjAm61
/NjTozaOxLwcP6IhTOEQbpgNDikCJCPU+tG5wA1BpZ4Qb3tPUwRYNjcuLePD0baW
oKUXG9Ic33zORrxcAoDrR00SrLExEhwoEBaUmK7e+sOfCEFrdGfozMyJy5/IyNYd
WV5lf0QFxVj6KNgaZc5EIZKfV6O+7rIDRbCwK7Igd5aVpaxk9oOXOvnfHXrLAMap
tofUdp09+NbNNcVF8XL9BeKF09ThnQQouxZLCO2Hf2S9j59SSQMBvnmiSeSEX9wF
v6A9hayDn6+q8A+S+WXUcY99UrrtIXcozCBJ1bdZkcnwCMyPcwD7O97tUDbBb31x
ARkOIJyJEuOwF7ae6pGTwPNJyuuIqSysxs8g5mvRKoZmmiipn6a89hafhW8rCHsT
CndFy1hiE4MwABEwRmQdOxjcTX83+LCT3GTqRQ6m51gfJp+8B3/Q+hbAWC77W8tZ
5AYzfDdMHNY4YBVCvCmlmSWWVFoMZ+EpgkfgK0wICzV4p45DmtuE0LfokCRSXvEz
wCoXCTdMuLMbUoIwG2tTMK5uQijdF6RgS0vTZxEEAB4Hu6zzWnLNw+MKLWZpB/D7
iWUoe3zotZpIuq3X5dL3CuE8YR8pw0AhBzLl86owlmrztUWlZh2Z++/A97QO9O5o
kLMUShwmIPquN2CUBlOb8pTPnhmZaC7bXukdBVmjIQs=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
M+FzCWi9ivDrLHPQV6DsxNBkVfQHJwXOPl6r5a8Be0MU5EJbKN0dVgxA0Jn4riOh
L892wjN/6bHfnYBVW7j4OUS3JL78lpOx1Y0GrlbVXz6XwIfCKm+ou3efkxIb7+QE
V9fhPUeagdCzlqYklF7MFRUAFcqgQyUgMBvGFLpw3nbPb5Xq7Wz8q+QIuqqhWWvB
sJUdBYuoLMKdSdAtBD15+yVpVliQYLaZHC4dwfC+VEbzjbgSbsHzJ9Mu82RTJHy0
gEiXPzFswhZBodLEd96g1Elv9NlzosCLbAvdUdTGkkArjMdNXp+A5PrRxhZV+w1F
UCj/qYtFeoAZIKw3y2L66A==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5424 )
`pragma protect data_block
5sCMSpJziXRBM6WmXdnxYhh+o/Obicv2dAjTolKyr3MmyNBRNBTunMvpeiPx7Z47
yXYNzFkFsCRuSHoOJ4tt6s8gjw1WQ7eFThxYRx6MK7Mjo0RghJ1Mvi+IESj64HI2
vsT8p13i2DrnOL923Kn89a/odFTh8VC7uWF6MJiEcD9+SDIaC5ew54KvEogXffQp
rmoLhEK7PZMeo4lDREgUVeAKWTxsDlof/68sOgf/ejrnFcxSvdfqpiuPnwZaTNn6
WMZyIZI5kHQIGgC1hLPbyhtaj5X67FzvHrbjW2dDDlDE0VI6dMpx9f3buSNzs32n
d9tQRHPkaA/77JKiZjYZ9COvAUkj99FxvfMFt0oZlzHxLFeosh+Fb+SX3aHgazQR
pdpiuMLyzmeh29yC/xMO+x/oQbuyyvGDyvJ+aWjylqQvwI84NKnKivy3gblJoqte
mZKXcwUPzfiE14DXhY5Z3J+hDem0Y2rXa16XMEr7QkK1ZhV3H7G2BL1YIuLCT5qP
7+HRcChCAr4TpEC5945RbY472NVOhVqoakWGsUlorQ0uQ93EKDHQ8Cj3+4bHJcyM
qJnRkSdp6biL4m2s/5JEcn9FQNQazmBA5M+uCtx3/sfAN1BJ+KyciD9zk37bU2IV
7wyumh0BeuYlbm6jDmDmhqMO5SxwkYKaQRGWC+BUAs9vBOC0YJbCTExiwLeyG5aj
X1xtLS61zLiScGLKxZohsLm+V3VmduJs3Q6CmHvlE1qDAbEIj+YM07SADNdksXWK
lMwGiUrVdrlQr3tPqVbpRdnIKvroc8/KQZ9asZk1qBvjlAmgdkEeZicAfmzYq725
lQ3MaH/aaYFNV+IHXWSNiXlroxdHrnXS+c/dPEv/mllQryNzJOxwxgeBbMhReTe2
Y/Gbv1TjBHGl35fiRxsnrBJMSXA8BTRt7SuXTdx46yx7u5343B5UHkUYmg9LjZS4
O0GsCjNYV2eq5LHmOgHIFP49QU/RQxQrfBBzwLTzy7698DHfWUHAVbAwJ3FcCc3t
rVmkAP+f8pOdXBFt6NqPVgAE2lcuE9FQF6YOH3mguP235IxnC/xwfa47Gn8qZKiX
pze4waQjWjkwMzl/cqOSDpl/xpYccXKis/8vrIzpJ7Fx3X5TBQe/Ry9tAYCoa6YY
Wv8ub4yE62grjZKjeTo3wWqUoDtbUQjfyzIMlRDwK1DrfLrwK09dg+WD5JaqQ5kU
zh/wj+SgNELkZnXvYbdnFSSaaRAPZlIt9rEPRw3RBCOL7voUgJ9spLPPPVDMeIyi
HWKFUUabp9HBpoUIbx82Mkz6PQfDX5C7VkbyG7aNgxWOEzEJ5MSxYGcaqxB2kBjc
KNGVNCYifIIeHPTW4Gixi6rO7Ht4yh/aCt9YkIodjKFPJGpus0zhE8rnkkGlGrHB
GStco4ydOhSIcEywYK6fZ6F/QkOG7u0QxWs1uh2e5JCGPKTecIvVK7v2hdwGxfJV
Kx4MnsgwvERcXFuzgj/KUQ+PU8fYP8mvk8MBmWbQ2SzarW4W655nlyPFEV2l5Bo6
XKfKRRIOiSHNJFL/ALYJmfrRK7JYg4tUawGmRO020YhzkM0PJNQc4d//bMKhA0Tj
MYdiU/t3fqDuHMRuLHqKRC7yiIdq4MoHTKAZskiDPTXPCA9a2I3ZLCHbSnVqBym5
6KPoYnvdPyaF8w/fz2x24Gk//dL18UmCBd6oXLWkCUFbkZqzpiMaJ1Y8TMx2lWR1
JWQCJoIIZzSaf+pPgcq/0a0QR2aCICU5fy7Wh4mPLZ6GsuJ81xy2ORkTtQmqWQDV
a0GW589FgCV/y/fRdaOXgfsQ1TidNzB9TBIH/aspXyTFVSSnhpnUaWpQiGKCepMC
Vh0dJnpGVH+4aXKuGiLPWEtuz56mWkCMArJ3ROs8sgRkz1+a6JmDC1M/os59lLWt
qHfJD5B98sHSkpA94jTgqNJ31eJDhGqDvIW7q5QctNiCVL1IRP71citEqhjSVAX1
fRdS+bHUHM5p1Uov09DwqR74QpAWyup+6PM2jUOkCcejEpja870rmlGG+iWxmyeW
2DRtgVjyu8KJkLe8h2X68XZj7tJcnTYq+tlnUzqHwEDabYSgvrcePBF+EOMY+hae
YAsqLzXMeRXVVgEBXCuGzFBF0JUSAm9vycuJ2DdgLI4fbbBl8txHOfrVj9Th+Ol3
jpQfZQldbduYr9OdmfEuVwy9QrFrB7aOBQSnWiPjUS/sYfAVIgpfoG6y2uBEbkne
DotBPROm0qibjA7/Z5/AgusH8Lq3cVhCKqDeV4f2CEicQW9r9S1+9FFFI49EDDF4
jQAOXG9bb8ivKIutph8g30GHQ6U7lo0mtKCLjMlcThxfWjvpOBwOoct/sCebjf9P
alqhP7vtTq9vh2pFqDJos1qzpfkEyISxyThS1zu0zVgIyJjOZH5u7JJ6lhSoPqhe
nHugpjJsxMPlt4KGlmN/U4nMmbscvKly3y3wvia7cPe1GfbJjwfWYcEuAT0uiFFy
kYP5w4BylGB3w2W22DX1uVbBqG0boNy/duhxATeK8/75V/U2U2qnvjYlK/IjYTyY
7qt2jHgAUk75xIwmegH73UnCAiphicMT84Qv9lHjIzsvghJmOFVurmvoxVpPg+Da
k55dKpCZH9gmHQrz2mNkLZa0V6A1xmYy5En+1iByVXx++Magk85CstEdum/Y0ZRb
svjEUSzrvtcrXxl5Ir/sgs5h+FxxhwaWRn56L/84KealfEnSKkDW4MXyBGSB+Atg
9cDsI/ZsP2ISs7HZtHtSq5bTi0BsU104Gj3LkbQSZD8bmeG97GMr8F4+3b7sEV/9
OJAuh+PC9HTgc5sNimhVNLQMrbsR5FeK/lJaRMSpWsXT/qORGBBEW39LWe0brDV1
gbpsKio6L712Cs48Vemn4prcVfot7WDj//71x9GP+m2KKGZxY2fhrhfqlhUffsXK
w0h75nCthIEOwUdjLZIdpnCrlxPBAnr7H3CPFxMDUgntyo0xaw9DX+2WWp9bQOO+
oWhS+Nh4hkzfIfv/vJiPu7QBACSYpW04IaKdULXCW/E0dBQ8YPzyPU70VYTniFi+
qJnY6/5iCVw96NCi+kq3kBrgegeQy3tXacqcOksplhn4c9AQrXVUXMi6NAy5/+to
zYbal4vXlyWCLo0i+xlMHToZUY3NSwpd48dJCaSzAtYPyBYSXZ5AiYBmH/cWLS7r
iz1xM9Rn0w97KbxtfSE0uazNwtXyI0/YSnPWaG7m3dnoOS2HFTyvkdmGrtS4tBH+
c3Im/t0tJndxW/yJtzhCIIDWfQ4dH0PU/sTVhCz4ss2l0fy2txNVLgPeFtLCtZDC
NNC4/ARzrZQLY/QXG+oK08xtIRnab414nGexfN4rtHOelM9ZuOalNCjBhlf1rsm8
tYL5T9na7tzxd+4/JsmBtuno6UbP1PyLlJA52hmXL3zg8owPXzE3Pob44kZQP78S
kNLdGq48Id4q4Gq8oA3bUXE13QxmrnD4DkEwdApmplPsAO2aNOB+Aq39BkiVFRp3
bOikz30xMjDubnqCZrA4sWWD1L2lV25s1f3zmGURJBoatzWSYeFxxupQYwxcJmJU
Igcg2YDLlfG/tz2GRvmUeYwo5PF4E62PLGPalji4Bewruu6rNuPruSLVEF8A1lgF
xSjbKeaKCEtm/bri72ee1F6TNiaBpXHCNqgIRE++rkkrVKRAQatn+KrIxdn8cIDF
Nv94F3fHKxoghtf25ByA1Y7TDwOSHaqo42k1x23prTuoM4MGtl+94zmLrmERxrNK
un8yCEZ2ORpjoeI6PqmcyDUXUYHsr6iDmeUI0xpnHwQ3B0N6lvJ/xvcx8DXYu4IC
EcnPa/wNLziUsUOrKnQDVyM+Uux4mhPBE9RpYPa1Igh59NcYoT6l8EgV0HnhyyUI
IzF8r+XEajha+72uqKdwCh5B1uK+ZJAEg5FEXKUkatEHNMWGMwP4oYlfvQ3+kxCs
WvrbVB4LMAbquqUNEl9/ZExdhubBOd0XpZi4Brm9vBeDAmiTDAkyb0bixJa9vtil
HYV+FnKtDEdE1c9QyD9BvB2qqGLN8t89Nr0GnesDS8agW0CZLvyj/lSsUh+kV/fk
9Rti1iCAnaQksdLlnf8xb9t5ba/Pzqa02Df4ZBA24vj2TZ9tUd5SJEoMULgqhuXI
JKoE3JLtV2wKcCU3mmPz9aER9N9xeP1oglq/UnX/PQqPsc9LX4JtTRTJBbMJPhHX
qEoBk28XBqMGkl21A9JbX6qYe5OzYU++xZWxdOX0PfpTUNCXRQgsZWSh3H1DLf1D
TZNX28OUWz2D6F+lk1dtB0bLDXfwLpHWfm247QD0dlEBHahVY4Hh/HJeyICt5/iK
gvYlM1CWNskjES1rV9xTJie+I/4TIevCignGnQBymprozQHRfHb88BgyaWiBmG7W
PAsKudGd7qg3VCVI5sIv03nwx2peeeHtEw81Ir7j25zdxp/hyXlXtfAENEtQskbc
N6SoeDnpmrtDl67ujZ9pb9zcryPv8ZsPz1bur8fulUMUR4LHRFZWTaZ0cOQPr626
eeTqcIPHh3eqy6ng5ccVGUEKZD+sGSdhDkGQzgehCqsvl/Fpv7kruGv1SowhvNMq
z+aYUOpJUyE/WcOI30ezPBwwkIPHDzmwiDqZ+CoblouH3r/S/oXOQ8JBsvj7sDXG
v5LbA7vQ4tYfeISRzzQpLSuOpbBTwwoWlDV+uKSUv+uwEYxhYGfSjY6Ovku/zWFQ
S4W0iCBUd3Kmz/vBAMJmGlAsPnMMGlnC/nEZlht+TISr+RAb1vIp6EIWnAiA06fT
I92ra5h2yYiif1WHbLS7AnRnxfmBv7BJQ+vjso17EsPI5IZ/fpYwR/WdzK+EutPf
FxUX3XGcvN7GP31cqJFXxxxkXQsGtQU+M1I7MEMuUlcp1UTHs/ulxwZ+/VFQ3tRx
1PxcmLF40CXXR1rTe6rmHXl9y4RcJO4nKRVAFM+QOdq255mMBfVl5UcpQlgYKv6x
qMk8X/cRSzRF1jDkEgXl4QKBbhmxcdnmIaxQ/Qg3pyVCCdy57aW7EipEo4o1bzbO
Lbb758LLGe2mH0ajfEXN1SDUrK8zDTGTAyQgCJYglyLZWZeE8l80ww4ULP50krpB
N1wNQvl56JL+XjhsfFBxGBbLnr1yPRzoemQ+/fRXDYEqdwjoRnAW4nPzyh7Ph9pV
IHGyZ+3ik9KpwH3AWQUasvVLdGOSc2XqWw1K3usqEelF5lq51DmJtT9aC+nSAavg
jT0Aa715epFPvBqADCHie4sPpisXOVlsguXsWFNU+BNq4S0mVgeMGaolsySMLK0N
EWMzH0ivi25qk+1Sa8YNS/nTAJBDgcyf+3ZDDnSLjkmskrzKU0Xmk7QcNdq8Zcb2
hv6wQ2ZmKJ74skrR+EeILQZGTSEslGupj5yxQZ65BcQ/i8OCzKl/1BQXZL40scRj
zVguR+uzwgVjAjeWfCXy55ApoxPKhyoVK//u5CtxH71ptF4+F0e98sqI0aE2veIY
mtSBe3cQTPJ7fF4/eVQiiXR9zrXWO8ENhrn75VfLFs0k1cgirLeOoIgSO3idb2yy
wwD8BQUWG78oLqIpHCAWBoLwVJUSjcqgOn8qXD24uf5OMgQmgHE3WDaAItAKZxml
2RsjU8N5d9ldD2qnlvxq3Ecfk5nBKz7B4Rr2CvZXUSHjwr67L9i+6Kd7aBbzKZP0
ejt2tWfQFUgzVUkOJzMGFWNJ0M4lfIoYSDWAe3RGWxy2O7OUCgDqHHJtsueH4e63
FIms8HDcManfmzd8gXvq2iIanECkumw45iYEfSHI5wizB5Ia+OkZkFvtrcWGnanX
16OArkHUWp6MrvrjjMtXviWOD5Eh+02Dmk1QgtRFKI0W8mGS3kv4xjde7fc5ly4C
WLfVKfMrxxyUD2Xphdpx7ZCHZfHlQXkQ+uZor0OpcM0OpZFSLJ9wf/6arcwLoVd/
zX2L9JqKlygYiIhfDQsa8h5RxT8/dTjeezcXWJtlMqdNtT5G4ZFUgm/sXJLnAzzx
pxG6sYhNicGVhCprhfM/V2lRi00tCV5fTqeqZhbrpz4Go6OowN1E43hw4zMG1ECz
uiXiurHueRWHTIs03+g921maBxRqzzA8xnT8piUdB7nAPYgxwQXTs34yH+7jYdTr
VQMHVDZTrRyLZYNLn//0ib/Uyrm/3FsN/UBar0GzhFOIS4KGde4VxxtQfgF2gU43
tR23Uzr/3tWlEerre2uFg2fKp+V6920Sw1gmotdtFQUClZH5JFvCpqHXamDh92EV
d2rJRpgi3QCSnhHu4SaDyCM8FAJm9z7zLRkKiNz2NzS8C7pIFeJ34JK/34JmajGS
uYzDdW5rOz9BwuFVPQUq2vRsXbb4/W207KT11WxTmwtd89cfG4r/QngQn/fDkxnQ
Kaq2w+/+rTBm/emelMZwSfG3ypZMpuuOu2jojQkuXMRozIC7SsTaslknYldzHieI
WUI+iG/TAoodlByWpx1yStjRTEyVBOow5UB2W8UW72EGgqjzmID8irawifSqNGBv
JyNCh4XCY6g9kQiUrzVh8UB3qh+9wAWmGP97EIzSSR5Vwuo48ymamDgy5YtKFFov
UgYpvZbLQ8DoTafpu+xWE5QW41Z8GUrcNU36+dBZNh8OowCdN6cgM6Gq8u3fISz9
sRnanALCdLSx224GSXTpDdI3puDtqewY8cNRytnGxuWpFNgL+wATfQm9x0LGxv3j
TMMG0S+Fr2bLwU93gu8MVTdEJv3YGq3fWo6ZynYv7P5D2t2QeEEB5QBSxwPvaRMk
yEEh2dS8fEotwVMNAICuWe+WxpEPtQuwFYiVxGJb5Qj++rpYAr7JOYj0IZ3Q8OZW
yvBhifkRfA1qltWV4sxDCFxKql7yiTXYGwX0gaZEFPyja4/+W6ONM4ZT+f3s+uv5
as6ax1caA0ov3e/E7uJvpSRvKw2kQ6WUc/yVfL1GLwF4xVYaqkPA22mzX8ojKcFf
zIkVfD/AchzH+/4Zp5TKilo30Y96T9by5gkfC9orNevXFwYBiFR4PGfZKq3CNavZ
vXRpdaoAD9SqOEBUm3CfoiSaxpH2V8u46pXtg1DXkNWKuzWPCr+AVePuKwuiZddP
VpS4DL7LWYOVu3B7CwBEcn+ViuGDrySksfS7LSSI3t+VjgzCdaAvRcaTYSKsVokQ
CqNhfEl1mZddafcNwA4KD/CEfEDrQ50gwEjmvNRkwQUqo+aYC6z5MNvQ/MaFldCx
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ZQK4o5Um/0gXxrofvIT7hWoPDaovy5yinFX9fJWT0TMzK+Lc1NI0kOZBuIu8iVO5
NnMm02n+u1LsefvcVGAlEbmIweZLa2Q5bnpg1D7i3TJOW8Bc0r9WIizDMMDErEWi
CbPbVeLuv2fv2hLmr7eTvpBNEINqp6g0C4yMDlPWmXVj4A5doezEqBXPhEUUUW2n
Yqf6Vs9zf0ZbqEQ3rZr9dnTTG/NcyKZSDYeqw1x0NK4ScElsSwPFA08FE3VFi0t5
cEsRdNhU40UypVDukRjq7GKvNGQnAEp8ZGbcQaH/1leTZcgvek0LqUy4zbjMestW
bt+vYmtk30rkjuJcnztxzQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5664 )
`pragma protect data_block
V6wsyj/z4TgvuQhETJpgN+X837dhTvsjDjE2mRrbNDRzWWMfHFqLQ8ltMXvj9c5l
ecCXqzx/VdrP4e7vWrlNDyKdK8D8u1CCfhO3I8VeZFUG3hAi4PeyA765oJwzsKny
PZj/NyRJsirXK9GMYWzbdtxsX124Ab9OGHliVd4jNcfwIu7BuDfxUB2IY6qctZAH
a9PEbWm9LAJtipO/5RgpDOuHabuMQi6in3fNAzjjVSpeTxV7neFdXrfmWEP84814
AwYDv9Mh/P2731ovgY0u8KeGZXkzK4sLNiI61ssiwBN4lhPbOgiheUk/RxBvb0MS
ICyocAjA++kjU3ubobPGT23SQO1bmGhksZOXyUCTcIimab8cqNnGw9rX6zqPmZyK
Y+hK7NTw+NlYogmrAMisaEhkSkPq8/SAXWdHXGjbsVbD+GYMLMU4xAmoCwA7t7N7
c/5QVM1F81WDznENZrqB0b9lOblrF0pGG70AmCKXd25V9FVLwTzkO1v/IA+gDMYy
06z6AYLfaQCj/9FBEkm80I960EmcN0/F0sqCe4UA9+W3XjcXCi6/SLTNK1Zmd1HV
p49cbzU6VxKfQBx0DBQVKoTVJTl9Qqfw90mlECEA0Sk1I8CG6T5kotZYURYj9udd
0I3U6T1R7w4HEhIClb/Hpr0yY65RpX9OteNNY6uZCLhhAygBFTHrSX/K+K4lgbAx
ri897tV/xwmnv7tYSuynWOPf40iVjmkxJfYIDQZ18atKC9YzdXe8mehkCK/fncQ2
lorROJgnDfXMIxCVuzHhRXOo8WFmtj++rbYLwSXHamdG4313ZnjFRS40Vuge09PK
EVM3VMpA4nvux+Wvt8eOnzBnI03nK4HB9usTtQ18Vg6S0sKoNZGNHuPzsx/4Mb9K
H0CjkwP21hJrE8xa3tb391WDb0YisRrJEJlxMF6ICTGBHY8g8oh4IrjUD8qTTH5n
Ph9uXWKQP934miTaALUOVexQvP4tFM+ZC4KmKo51E+yCa3w9jG+VD2ffuSeePznj
qHIcfrjFUb03NQplNmEdEvOUbD8QNoKy4BCPH8ePotKIAfmKbY2SYdGZa0lDFfc7
JCg9RmD8zmxnmocr/40l6DicaMT/tev+8x1TxkLuotKxNfcZrEcFWCgd9rqn31WD
6qtqCiP5QRfkKXSTqvSkAyIUy3e+QlzupoAyMT5FMF+5XzxHDqUQi0fnNLlP94Ft
LPiACzlBPKOAkmg2gDVdOkw7N4Q4Tq5I7of29w3omC+kVNsCI3OJ2YHX+5qc3AOT
Io0OZwLA3IS0Rd4YNMQCBoVO9Q6ZPJQd2fwJOPIb99QCwh5tQYP08PDRnbhpYqfi
f/B4S59Sr8j03J0nblPUMs4y6RFxUQAmHuAqpgnuY78NOcOfVC9g+PfnDW/LcGX7
CWfKcrMvv2rZbyJ1rojyWsrG8fwkgI/FFJB4Rfjcvde0zRu27xvGdREU/eYc+ymH
SoZopj99G4JF6si70z7tcbwqhQh5qfioyuPfEWqJAEjgGc1EjDMj6BjwH1A0DCMx
DO6g0sI6dvDZPqkN2GJJv6HzZnE6goxI67VN4F2oR/mLgHXHWulSk8WXwnziExQ/
1+xWf1ofNRNrkUKXV1nWK2kSPWNwaMdjs6mcVd3ugA2885kgUpsruY7XhNfeOQJZ
uItYx30xpxayOu7vwzFHFlNBfVJiSCb9FWgJuEHhWJjhDnW3kina2JiRgWJWkgk6
lprHgHqgmbGYKHttMj8iDdmefYnt4Wn/3vVq6naj12ZBwoXrmA4z1yYdYiMsXFJ7
DVXWAPpbJZSg1NhgIzqJazje/F3O1EwMlnpLzts4aMbYrrpiUhfktHRo0It9Jeor
dUV3jdeQpenn5XMPkzOY+I97Znp2iJXwJQhHRlkzVVpDrMRCf8B5jgKaz7Z7LOKH
ywn2+A3X5G82DtzSKctoOAROfubYMDdswlqybMeMnOaZzdYrx834tVKX6XO+NDus
gzl1uj19m6PQGNEn/Cit+o9RFb1jAIUFAz9mLu2kro8Og6OpAvSJi9NUar7XANu+
LTVd0VbKMe+sAHkVC0oEv7WMLcmbMKDHkG7L/a1wgvRRIqnlIGjIOgEhFOwdh/49
SFcGHbbI6h/9ZNcHYRveJcb5hEycAEqNA43Nt8JkW6VUScjuKHf8VJ/loxPLFh7M
CSb/NTseLYD6fmC4SyiZR+nFIvNn/vGPvC+M7La4J5LWUepa4dC4/MJU/kcZJnOM
XubaINRsGBK72Wll5ap6Fm4MuFQ/bD9Cr62GKEx+K+KA0Wt/pO9P9Ap01q+1Vw3M
KPhgRVA/+yZYoAP7fK0ughliHUVUczOZUmad4wFfafCWBqS/dCPxCURrgXD/6zlJ
o8934fcTKvShpxx4lFIr7Fl/lrUQefmO+nzdryNqJqQT14Bx5Fl02TM7cXt6l4tt
Ke5JPJ94TuoevRKLQDKoUS5mfVGZ4I+tnRfNdZGG0lhcwK43eElVI08d4/2TfDaa
9sznQzcLJPL1XAgxjR6HpWw2LmTspg6Aav61wLViV78JfbZ32Ka1EJZ1e/ZtRSX2
GPKPJnWaPmio46g6qTmQQhebJO1S7VmnstjQmCLAiX2ZQD0f0D/XQV+9OF8DHA0B
IGZxvhHp4tCdqryRRzWxkXPK1/MAKrXrS+ATWqchx0pPodwrasRzRyPjkR3vsjrO
RX/1/Xo1bakHHCW99v3T6+I7u2tfGIWRJgwMmS6hCB1SBA78896CJdIO6WEWzYft
pm3+ux1KiI4uEBFAs1a06dDX/dt59+dVFssaeiP0inTruqUDA6JsiMUE2iV59EQM
T/3QtIxpsyzYmDK5o8yI1y9ymQhlorwhv8QxThvwtVEWwTmV1sAMFo1+TN7+5Cvs
tNPLuenjBrOquhhy+qOnnxZZbySsar7xy0nrX3ZVFmoL7mGEO1eqJMe17Wg05Ob6
W4ASqY5bMkr0WuSBOpCwJE/0a0arfV9s/mEYpa/Ena+GTKecRfmrTicIBH55vBB1
cnkwo8NKFgbTwdLO1tHN7+k9kbjK5WBVkz0vHlHFRyV9PVFJWRQ7dKerzAdjbEpk
zTjzP/JsY3OZj2UdaBPz35vlc9H9EMcpCpU0GerW/SaD4q8qLdsHHF+8rnKqRB19
mpiZYGEvp+jc7SALaL2NnQ5+xGZkyYc6ZFaWyfQgKv1AGpK8fTfvamPVoiP0Gx/n
YaRipnA9ftsiL5dp+DJlx4vepPWnDPQsnz8hdQSY2r7MwMTKLAWBc5O50lu+y1jh
qFmwUNdhXy1ypKyaPlwuZsqla7qKUStlSMRh3aaiz0MaP10XYOfKHsGYURCUbXy7
gA2hPJVdskZcHODOywNC5Sqg5MRzwjTn2auyd2SfJwRWWkcZI804eJo+B54TzJ9F
tzvRZ3UvbliL8TVQDem5z1HWQxuyc50nrsBgkghMcJnKOiwwdzolNKuf2cjrVO0b
OmIkXq3TlwW02Uhqzfe5fxsbuPKn80nMzdKAUMWIXAW9CzEg1fITGlf9+7AFVsgY
T/chIIl/bLzw+bNqCGkQeyQiR8yb2kNv5fuI59szP5QXlBddG5oYzv+WEsnjAVI8
N+SnQkkGVrbzVJjeRzZJAbTNXn8cXByEiV/WqKsQIRIsHFLsxfujaAtgWmycVu1l
IjYA1Mst4KQQ/VqFI99CQffMnqxXq0ref4Gno0Yx2KJ7sHsXI9hvlR2jjTZ7Rj6f
eKtQy+pHnAWHzBaKVgkw5yXHIV6OY8/tJAVnGKcEbv8wWDCIeY+M/Q/ivR9i+Jlw
ipLvLTc7v8xntnNdmxUfChjIiHrC2/W83xMP/FLVOHb6NIKd/0UeP62FspZmsyyN
JUziMzZqlJ2ENUIXab3T/KilHMu704f2DU8oFakijcfcAlER0Cn9nfyr5kimCQ9b
COR4nSLeK1mBvcwjMIw1bRj7/bfyCpUHdw9XQwJSrhQSS6NGKYvBu0W4aY1FAWsp
KOhml3ejoTDh1qnKnytxt6zE8dqDz+cQPFseIyOloFdEcn0QugPSRVH4KJm/PNJH
431r5ULa7bmuQEjRKOxqej0B1V9n4IRsCfhq7Uw7pIKaKhJmT8YnLmY5vxZAejNt
IGjd5oH6+n0nuGgGcEYGWnxJOGrBCY9MkjZN14KUGlE2Brkh4k2ousOhlwEtbm8V
cN6M6pjh817zBwniHxlvA3OqnsAOQUdnlsS5DBXGKqnuQiYeufwiMHQ2HHcfnEuI
UjrY1VWtGxalAqVD1dZbgQxTg47oJFhug2e8+288FYvvjOjUIPdtvNJkcPPLH6+p
YKZvXQIWGbS2gSb10Zp0KUTyiW7MgQ/DraWc8DOnXArhnzVtrrELRmITWR4/aap1
RSW0W3vYg5Gamveo12Uef+GyT77Wqz6ZobLWycqDY9HvewJpX0YoBukbcdGE6zCy
Mg6C/6p49F+UOHsmmDtMgJPD9+RwdKGtt/lhZe8yPd7P1UzhEJQOuRlvhhAyiXvl
BwVt6v39cch7/XzbW1SrwvDV8m9LVDJkzXILpngpcJ8FHpf+3Z1/BsupAiXOOsUl
tew1H+MOj3tWMmq2cEJ7ok9lqqJ+8FZnxS7ZtG7Y+1aA8QhYN4a7ACDN35G3+BWs
dNlMPhTEcxwpEgWjtS+0fwCjmlmP22692LniXwY1NdE2531sSkwKL1RO/MQpCruJ
5Pv3VjGGNtFsr+QzLz+rBHH7QRhkR1JroreS6GrR03Y14g1PdEo0bhMEpjb1nRVS
Z3gu/wkSKZfdSZ+8vbqbQEpObmarQCm5Ui6wmlj7xiq2uknHBNHIi28XY/rblGCC
02jdEvMtus4Xg6w1NP8MqdmDxiRb8lWpeW/e7XnG+4pc6px/sU371fefibqBu7GN
CQ9xcJBbYdvD/lpRqG/E/nPEhh1FzSpkQDFnaSUmajxQf1TBnw376zxFaNy2F6H8
8M9S8QFRfVDq53qNA6pWeBctmZANrNg9ElCWJQk0I+X7qsScyPrpAdVXDrtjpEV6
+xDApXQq+iCaE7gVHgdsv9nBwBpEXWFQ4aN4b6QnEMHxPRIdiG+JpPYG6ZpsKa3j
/yRukl76ReZKlwPLBuCl34w0gGcZaA7MkeTvDOc3TkckH9fqf4hKkegVd67C5r7M
3z4t+KcDY+YjSMBRFm2B4ks6BMb9EZFPgu5Wt7WDJc7IBQmT+25NGp4yHf+OdSd6
GRqKDvhowuEi5b4xvLcvE20KK70XUKI275j5FQ7YpbFYxzUftUJmNKwPf9KzHwlj
hrcX8FLMOeWKgY1L03UkRH67q4I3EjyCZsUoomThlYYHFRLkSH9WxEH0nCI7XlGs
stqhIr3AXU3EQSPBQ4ZjZuz8HPXTJjIQe5pIyEzHyo1bAAzZ7FFaV8ylYTZbmE1+
Mxa3l2gIV+HHMjJJd9kFEnfpEYxLn9F2rP5fzE2Q7N6EeJrYeq7e5+i/H7XHtQAW
yKHutur4HlEgYk+0a7PzocvQAP9BJMcKmpYj8mXmrMfA+JLS3JKhNdmPa4HcovRr
EdzoZagDhb2FkeWYhGK+oNz7htjMZ0Ai8aLvlzHuPmUTgNpm7r679E3ep7d2LWsD
BHYMXP5rW+HPqq1NM2/2iirv6LnYhG8sdehdVhXtQN27Snzd4Ew7fI0pQd5PR/Yt
i+FMMz/taV/qf//SdFHI5zb1hor9DtL1jqkjr3pbCYW1GQHKzSPV3ujSq9+XbGDz
lkTEGCjO5riqH7keVUHHJoptse+lj41MBjgxcjqbVPqrioMjJRbtp27MNMPGhG21
S25EOHX+8LNg3nu2kpxxGZ6LPYMlAnghCSHqmAVO5WRqLpDPTidSVaa0Tnt5/2AL
VpPHOTX24fhrhlisVt8FmbFSx8lohDISbRqkewoKr5mDFz5BotFX5oLqgz7Olrqy
LZDT4pdftqjVVoWpFAugVxB8h3HBkAdJc6njQ5pbOfymLWycUivKvYWOIM4Hi8tB
J1tA39T69AyTlTZrpgTgOmHvh4RJWYgSWJouBalZT8ieUdUsV56YBS6F+qtZClI/
4rP88iSzXOHDtj+hQ36TyWktvnUCSWnRV/C6fd70OoukoAZbYiUbQmjGmfBZzL9m
4AT4ox+Zg+/dEgbCCiuRj9BORZR9qYYZOAO/TZIYEmxgOxLGCtu2MqdMiTGSsZVP
kk7jy6p4dUhwjjLj5rihskvwBfsGoWC5w3+N+HCSX7iM+NKxuM1RtC7o00kgJzJX
de6jqU/OF/QMy4OGlE/07P3Z3+B8YgeGmfnwsaUGLBGjnJOCIWIYTB0SGllCQUCM
k2JhPxxrzVz1C9K87T3T3S6liI7swYsJpyRFzvSVXTRLZEZCUED6jaYnBgR/XaSu
HhFGpYAJkyBiLLeMBnqKhRWWYMatSzhQge4dG3fYspUv3gBx6/2xtTNT8WU2K8F+
6Gvqz0SCM57TKzFqbDhojF6uQ2Y682ke4xV9IhmTDBCrKFW9GdnDGLMK6fA2SCN3
RoJQrH+TIwWpDnwOWo6gnSSWmALiymJYbs1No+6RA8NI3h5tzaaYgnsvJK86E7jD
NLWOnOutPUTVbww2zdYVuj2cTRvROZP1bwlSQqhjTqwx9GFe8poy4d29Wp67G7DB
x+HOmqemZ1cBt9MwpRpVFohyWwD9dSMvHnMzB5i4Lid5oBZomGhdDhzW9TVq53lM
ypTpohc8RBEdzPsCxt6y1NRph0kByt00nTGbv1x8HDjcqptVW/WSTeGvTaBhHlle
wdS1m8rnJZIBiF6/0sWx4kktLvVTLCC1Ndk6NcyCP2DyKu/e0yXAALs7YDyHZFEq
GV8gG/SQaZW4SwcTzMWZW3bITIJBZWm+9ExT1AbgygKzgPn5oNkYkgt/dEaB/cIX
OYwqYqd+aKsrvD2OSZD/nv1f4Qzh4CHZ2c1frTTfoC8aB6uDd9/enaWYSN7PrBOT
5wxVFpoavXUhDUIk34nrnJDwfH7EL8wXuvciDey2ad17mZKsY+gixcv3XDFsFLLn
K2gjC2tyxgHHpjzA+xJayphrW82Tv0WyAi8TpdJgKIEczIIfIacmWugNEVxnyLOW
GSUOhQiK8IjqNy08/AFuVfxyVjJREVtkAleiG8+dXm5TgYituiIDLy4OjYX4tn8P
DnOwfvVs0N1WjuurapWplT+AjRDzWgRPh6vhVPxqV9KvlgYVhGgmezGoPXxRsgFw
bFfxdTgE1c40PAel20CDR3qnvANJeTW4hhr62G/hS5Au0bsJIOfGllhx4KToKBhB
37KdUS55p3n6QiiqysjABfnL+R8SMhtE2I9wWVRw+j5X2fzCT+jJRdmjEGPhxRSO
GnVxBEbg/Qlk57Q8IhqTzWqgjocmXUs2FSCFXn2f8fqx4NzAnGmRPsrWUBndSuIV
gtWwmp08/957ixTcL+3RSZ+R/UcSKH1beCi/DOvhNKq+dK2ui3zV7FvY66/9iEvM
QKH4baQtknvQntW5H1PitPgvRYizEhs1T/HCWuihcozbHZ6KLNddLNAtB54+gJr9
VL9CXuIKr8EDSVgZzYGnlXq5xUCh699HLx5rPOV/XV7bWxkVSvOzYus4l5axNijj
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
e3QkTU8sI6Pj2cKV841T+K8a1A/YWYBHLCTcN8HMVP3+FGPD5D1ZWkBjYPkOf7A3
OfOx7FGr/8JeYqksaADJ5fCH80ZhIiAISomiYK2W0MBdHtKT5rUA2dkE+H5AHz8k
0YKxcG6qZyNt2FpBcaiBjYYTbtkAaXFv/Z6Cm3ZUBGGYJxq/5SIPa+qcNRYzASSW
553z6WJ4LZjeQNsYJFJ8eZPKf/eZL1E1Yl8Q7d1wXs1bFE/9wyXEJOMwFPV3+JRr
ttl3PKv+PkYBuzzxj/JCg6TgAckSnQqeffOhYSDYfBDeAl/1lFaL6JrmkpwRUP3c
PDx2SGnvOT11jTCoDfnSKw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4720 )
`pragma protect data_block
/0Jlbx5KC3PAGEwr4BDoPyzav4CzI07a8B76uHEwDBPVE+muJjpIBUEuSyPqQbKM
SjXd8z7N/eqUVV7igkm13oX95xeGv02ozCDEkcoy45nafqzZ2y5gj0VtDsbfPFU6
WbxFdxWoL6Ic/BZom+C8Q/nHXA2Ez/ylsCQRhH/5mUoi0C+Ej5ilZxq6vwt8pOAE
Pzvoh0FGjC1aVixPWwQaDKFtTAEFc5embpEeXfHp458ZAenWwtBfIIo03+uJOBYs
vqL3YiO4Ga730EJhd9L6hXELwdXmrnk2qcjBqG3AkaxgCb4cBGQ2RTuVdt7KlO9G
xx5PiSyp9+YwHefMLp/B3Pj/yAtM2lqbxNw3P78bGDMINH7q2Pa2yYdH7fyOhSmv
nRc4WdDRn4NNGjtbM0yZtiVMPxQRj5P8fiCSOOBIdz1ehG8Di4gqrquSiwD8t/8L
KuPRKPeEjoGVbFwrLPeD2RBxnrCWpsu7lw0spmK2wlOMGpxkUu2GrK3mh1HqQ89Z
hPH3LJDg1C4YutctAOAJdmQzcgKT4qAhLKZN6kISr/0N/eaN0Fw6SyMd4YNIdT8b
hZtaIAM8/u8oG3DVsPs7nwMfgU57rla/sXsnBn5ygHx5STp3PMjIf8nPwOV8sQAH
h3ZidYG5BYgOMZfwa7LXQDozwXQWaCUjj0oWo1TYUQj/iHddDs94qIAi9udHKtM3
MvnJauTUdvTZvt0lFY4jHgxTeCzCK+dkSSmpHxNk6C8G1H67FKE6i2tWKv8hnY2M
I4qEUGmilFHYWncPjEveMMjGm68/13WQcMbO3vDXYFDf7WZcu9GvkEAb/NrPSJlq
PaOZ3wyOiFv/LucEMTWv//S5fLye65HjD7PGxqL/WrhnnVhSjhWjtR9QzfJuZztt
QWT5K9sQFFmgEwQrNGp3O/jUco2CWzWdCHQ9Gig7Z3I6+4bW/T1+7aa9E7jQ5OwY
8lW2drfcXsCVdq+0lkG9OUrXfDyxCM3JjN3dpWpWPcoQXoP/d0B0mMrmqfWTlFyh
8MKwUez5l96hCYTlPaqPbq/PLRLVT0ycniiU/oIVWm9LceKdYLUAu4CEy1ka7h4A
voPjXIrsWYd/+hBrkE9aXI6yoKAikqooX2SqdLLJjmJD7UwHnKzWcar7d46H9jkL
J+ckLiYd3/EoueMy5lBmJLm1YuS+HCeZsN/bwE0yF91Q7uUJzqDmfPnnwbFylqR3
VlFCGzrR3kY10ROgoz2c5GHwOANsjwaLsmJD2K4k1JmfGkgLQAlHZ4P9/NdgBioE
gf54xESbAgZxtAYeTfbwGuMyZZtwvoht24gOQ9lRNvJk0Ai96C8PYjSabmXvi944
pU4enkAMgON9pUMgzy/KhAPBdVXKslkLyC/VxqmVxg5OgLIdlk+p/+HldZroOWFE
DXxTK5C8DjYM1DmOfDAZyobgg2vkndOEgaRUacPbJjxUDXGc9SB8g7/boAL+RrkB
biQezRyVctOV575EeYfnKCb/5e2ZnFNn/DjQXoYsWpDgA5tXIj9Dj6J34cwG4/VB
3YFs8Tm0Ivfr9YzZc8dkGztUY4ytbeLWW5QcOVCPiVG5tKjmNCNNLqQim8029OJ9
NuWO7Nr1FBJa0vXdC5PHKf1UxkDrLVSNkQl/uihkoC5lDnAj9cXv9CY7Z1WrsJO4
Bt1oMXGskIyUbk56old2fly3lNgGO7kzPu8BLKHF0+W98NxNldiFMTgBHJXGacSG
0Qpn0cvbj9n4IOrd/tjMpjNGs6mm4Ib1atvNNsZat3SZsnvy3oDvJp1uyVnn9Aub
z6EciNM9NoEGt9ULpoyY9wq0wNOf7ReJnc3460CpqSjPsiDUVanmoHY2ywhmu7Ap
UAQzJzPFGCjj6IIbRmuxPaLdZdKG0pWgVWzJt3feA+ZCRn52Oz5UcJCqkcn8y4sm
fyD022P3EK8fsM77JgjrQBWeTtJJPNaPDOtrkdc7SPW3+ZHaAeZM4sMXzio4b9W1
aodsOoV6aXcwPVkkrrAkN0i9DCu9L87KniHIUtAtzKCCborYD/xfvOjEVUoDWrMC
NYvZtt8ko2bEUtlIKZrHUMln5Eu/bBSW6MC0OijFsMGV2pgOJlFi2lPCOpDyt2zl
actFQspjdr4/f+hzrS1+oLVozNQUK0FWNo18Uz1x/7RVS52kabuvV9kaQGrsZQG/
O4k67F9pDBE9gYJ+eMqyEmGVdnlz0vm+SG+/bGHpjycz5uBl36Ib8FmnDk0xfqGC
QCHy8ljTpo2VvFHxMU4SALs1pdW8C75FKLmCYFD/D8G97EvDDX+9/skjCUOPoNhV
xiplLTEgGRtRk8RNMdlOpyastBz7ir9+0kCmvpvTLXeFEyI5irT0CrC5mM0DlJfM
jEgDM2t0xESvEu/3aFAZuJXPE4B8MwHw4EZDTLgJRgH2oAMhs48qrN8tuH/yRBiI
eDyVgoBVhptcGZE/AnUywE19fmHMv8Fybv4S8sWIcvR+TjX1KuawIWCqleD7jxBK
+vjVVzfrTWRo82xX3ASNq/RT78eHVJMttCO5v64KJ4Lg1v3bNSWJbokljNDF1/o3
Lq/4w4TkPDm6fWphO65r3tZ4YGPHqXBVaTpwLrYDU3+yYoRmiPE/mingBleKKiZ/
5qXPSTpgVzgqtYzCCXRnBlta5QQ6amntr4QXedu0xorIThjETFnFGsqJRMcT6fCs
mBy3ITxT3bVQceuK3qeDpT0OPNsUQp22+ubbsNKdNEORz8HiTwvks8lsN4Rl7WEw
/ftU8VI/EKwDlceYcxV02jAFkP0d3/kwbU4bIRr+kZt3+43tauvn8c3pRkV/bOdO
Lv3utE/GKM3pHu4CsgplVSvcXk8st3BIui68XyvII2bIye0m+h+ZRs/LVO1yhXDf
qu2p8t4S5VSaF9aMa0fGUzaXux4CAgep04OwurZJaYRNbPceiy0/KnGHoUIS76zc
AlYk3c23vvlp6TMTvMnNT8+ZdAHB0N0EYmW/JXNFSv7KX6QBZWKDFgpjHw8yEyeW
XiKFRZzJiF76Na+5HEZhftXaFBIRoZEJrpmLsUOW6NPvkyij6U43mZ8otdjMlW5D
/vj1/Zn8pSq6DpnhsOrB29+mWwRjxU897Z7OoodA1cywtqjyPVYcAg+7KUvqmKab
Ra0qRopYY/Sv+pl6fQM5wHtG/P82yzJCHdeWRIo7cNRvUMBwND7Y9UnvPtv/onsz
sGrvOEfdxWQsdHJPWMCOZiyExui3MNKvNxXCUMTZwHXW3QqflFtVoFclYwQ20pPm
wXuuVQyd7RQ0CG0OjmrN2192U8b6cgpxIJGcKrwHhtU6nMB+R2Ra7/igLSATmo24
TDRCFbiKNrC2ODqHb6ifGFbZwY25aC52XlZE3KFK7rFTPyFhb+RjBrBuwTe4qptm
7/hOcZXnTcsxOpR8wafa4Q43EXM42FoYRymenjY+h/ivUXvLuhjn8qhipErCZlyp
vCwQ/yV9LIJ8PWFgrDGJIX4Nox2pVMNedckobw61vuq4AuImhNUXyJOrn7x0Y7t0
hnophlzGLQFgKuaC++RVosf1QuTVFA9aw2nk0yY3mqGnn1nd1knWlTKCdLe1n7EC
4iEOP1KllYzgs3NJny7G9qTHQYlYap56rah5Wc9kG6tCRxRi/D8J+2bHqG5ragEO
IgGnS4ClSJ2hpuQXo8KKFttD0icTklcGFZC3mXTS61SWLc3x7G9+vazSoHkZEehT
k5w6LVSQVsk7+1YOtSULcXd9P+2oqE0CadEGQ7mIAwITQc4QehFF/mxP0KjKZzPA
HSNk6YYC9UUUGNDEauxOcKMVXwCQFWhB+W43Fm3bVupZdRhYzxFW42rMa8+UVBJ+
JOQDwJzCf6Jaq63rW4h1DP1THMoVBH3OSpJ4qr6UO9CE+DpVHErO43XGWRfGOf+W
dz7a8oIxZTOxA6Gj7EFmNNox1zmvwLJRZfzZNVSsKwvOkIPk+0/WO6ta/Yf5dv2f
E3Ty86MhDBu7aC2JKOKIplLXJaidaeVZAdPUajBhJBNNf78Y5GgVDeEUKMd1T/Sw
rxSNlGaOymyLGv1het3uHQWH50siM7Z11MRNQElLYn6bJGv6goTQEc8dvjdg5dOF
/njeV4YdMrHkgR1ZLdSHuc2v+53p2LRYwBnHSpKZ5Y7vroiZyMd4qZNPlM6bZePc
vwo/i7a5s8Zjdq7VjE+RUKWNRIglXxVg2Qqsk6OYN7TSHHLBMDKNxmHto7n+v3Ma
TQ6jFJ6sLStG+hnThf8NjD36lw9TxktTVAJUl49QZO4dGENhrS6uPB0GFMu9JkHW
PLLuRADQ5W7sZpEGveywSwR3D50JCHjCCkctnl9XE5Iz4AQXH14umhQvA2eez24/
eb0XDcbNSsXsZINK01Fz/LKhqesF0lMkyg3Xa/4gyzs0P9OPFo/bAfQNKvF5Vn1L
6bY/P7bjyeGIb/+RfX95XhQ0pW9UBiO1sNyQ/WcWc3pY2SoJpTrrUL7BGusXsmUh
Kizyvwlh5k4OWrZqgbFL+4DzZFo6+/khhS/gSvErxVVm0qTi1cCsW9Bp7beRGZLp
pQntLGJK3gzj1zV3c/wm25FxDyDpXqX6+LkNNwH1JrMpNT2yaYMBX7speWTcn/rj
4Ci/XuFjTad8Cqx1R7d3M4p1N9WT3G8dowZTr0yhS8cyU93zKXWU73ARUrJVrjsX
I3oUUxWBRt3XZIfIXOjoIRv54gtPD8uzsqk5oMTmCUpI0fR8FB88z3oVG7BMRwG5
R5CEdnLkiVGwo4G+1NGWQ5SlKMsNBKWgR1TIYNkQv1W4O+H2u9VAQRkR2FD8kwck
qBcZhHCypRpEDH4P3e0rt+sV65j8toQqvwWKJ3dswv3XIxZ1COO5OFLhjM7H9mf6
Sxs5Sqq9SD+exWTPKXm0T+98Mj/E63HZ4E3ilAvnlhT6dfqMmI5R3+Cyu/iAlqD4
f6Qml+3J338Aeh/T8Zlo8hOisdsY2SB7NEQXO07i7V6PxKJ4jLmo3374+VJ74L/s
2iwq8Xb5WicOVjLTuF1DgIcMQ+7yMaCQLbTjkBC9oTs9HqrONqQFPzDrQ57kbWum
SdK3rluee7l+D/tsO+GMLzbWDukHkfmOU6GQKMbuOKbM1rbdMy36tojaeEKVmqat
dUe91gA3fUuz2EABrSr2ZgtiJjIZJALM0K/8OV5AXbbme/vkfgP7SCim1XQOCJwl
1VXn0LgbWBkuR7/2fCOx5eFWZJmcUbPCsAGHu56GoE0EtpMQVtKs8ia1d2YLbweU
Mv/YkwyDiKHTBK/BVDshor49/LSZxVWDiHNhEYQM8PLDRQZT8ypSlCCQCZwhvMTy
k0SKjm574fLTOJxh6wdktHdivId/d6F3yY6tsOsqSMIpx6Wvz/VxlLt2u8uDIXC1
YX9d13y8PtxRT891zkkGgHfcxGwUPk1y5NNv/S3bSi0X6JSxHSTEweL01ttA6FqJ
rsZTPs9QOqf71vtHerfwEd2wzG65+IyfVcE0H0nNS9IW0VfalU4o3WNDdxxgkZiY
J5UJ7ugrkSM797whJEYlqEUnlERR1dOdZF4LQjY+17BVeAkgotsXwSaAJ5KnQ+oc
cTA5+bvyhvrUGvXMMUe6P/4oSBsNk8t03D/1o3ld5k5cc8Lndz9cyxxfVAZ4OJTO
/c9ox+EAw9DEN1l2tcLHiZwBqzQRRlEbPBf4b/bYpw4Bzm/asA2uqRfW9FXmWxD9
r4TpilGyNKkAyyEiCQbjiu+rsqCS9TkRgrPxrxw00eL97G+fYQwWPLfGjawI0+En
t2JQFhAUX5E3yEPX8TeoLwoit3l9hNvbY0kx0QRTz8aFtaoHpyVtcc8dqAx7OxFT
la9Fzq1M4RbKmYxjbqOnXLcFjjSiCv69xPP5BZIN7th6m7XsRPkBEWY27jJrt42w
g0vJnogP47KhdB0nLtRmH0juicypNC7K0It+HWuniz0sz6/001KnRyTqiRKMe63n
RWts6WZBH6egiibIXWwCcrb4gcC820Nkk6W5LdnbUbXult8GhXNi5SwYUU/PeQkD
OacGX7eVZSbikjYisp8a+Jcr7hnVm/BmQUz4vQiCVkT7bOMLydd2V4v2pLqOWU1A
8i9Rq0RsJdNH8P1Jy73DH0Rxf8lp5c4chauc1dAZK5SedUUdARqhn6+E2/74I0Xh
tKulMqWX52x1I4xhUcmfowz2ol9sPOAlSmzDF/MPvP4bb1OY+O5O2zStsiC9IhCi
rRiQ5WND0OA/FYWW6ndEJriAYa1FhhUdDPduphjiW1yYVDGDP09AKhRA6/do4zl3
xcGrZYjQzwiz5athd7AKBw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
H+U/I+OjcNVa8DpxX1PSROrc7DAnrAJNWzcNTNA/UBbbtyIcQXfiwd6tnL8u8hGp
64gQsTgNDg98u8ckDpdpiEkc46oP1ZAD3E39OEzjCxFQCUYKjBoegw4I1JovRGXK
V8Y3xufcXDfIn+ps/i2Hpn+nIJ7rpZ8+qz+Ubilcv+5hW7os3GSOkqn2Gw2gsSKT
hkVm1vTSJK2qgcdQq3imzm2cIG5wJuueUtsFZn4n1gOyyVlUTZdzsCfkp7tCn59/
fHjPSJ6t4ktdzTUN9yIPmswTz7ttYgaSoXe3U2moApUT9Zd7XEORttUzNFdzyago
PitHcNLJqAECwrkfe/Jnnw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4288 )
`pragma protect data_block
2xCCztGU/M78WYQcw9XnNY/ODlHwrZcvDSdiwGpbP0bqKXohvV7ypFfVPP/2XtWQ
r47+X6GLro/SEMV25hibPNzlpSxJGRsiWzlFq8JwtVy7BaDPbrtLvgCA48FwStHj
2dRqJf3VLcmAUzsk4d6NJ3CWLQ4lnr9i2jAcVeqVA9b934nNNfD+VAk+HNOluGhU
yTjvh+s3XaqCgby8Ef3nL5OCXupHs7F7rqsN3yHqA58fhT+WrPU7oLqVXA8O5JK/
nwIx3G8M8vye01S8rVmD2pEI8Pqgq7h7pnszJN3F/WCJeYn04ttjvo9HWyGTmsw3
OKHL3hnnUY5xOmW3QxAWCVVHmwLwm13k5NxE0LJSt7ZrQePxbmywKB9V8xE/owGm
P2PCl6WvFA+b38t5ZtJdFFox0avHvJof+PgRFzyScB175dWl0ulKMe0axlM4qgeX
KdllOJGntMQYDU2r6ZOgIm88Ws7svMs3cS3LkZs9uLOITt74G8t6wY/rxtTgvdl+
gItuif0ifbcGpWA51qwOc54RppqhIJ2DZBhM6wgq8qAXq+gCIA5E5W0uhQPR4dBy
uOobdw2HgJZSch//NfxQ4WXtR1941FgYG7DOC96TafbbylxtEHEd8PU71n43lPZ8
Zrd0M6sV/N8LYUkA/IoAPJNH7Wb4KBhbmBgIC8TPiunXh5vNGzad3BEXgZF04htX
DcMVR+zqHdJ8Um799Z7IlKtvwwki9ibKFhs9sy5YWsEMluWtzv2qEbKyOccT0Hp2
mMdHygWgSGUl3N3WHsn6CJb+7zt5W0FyqMTA/c6auAWzhiKmYVA9T46lG01DYCPe
KbrrD4VR1rIoEamduv7lsryAjE87YuQu5FBMHbpsm5YZ2TlePrvHLWtOf9HGuCGx
k6IOKq106DvrQ39uCWRkTFRqN/wtvnznddHf0FG7e8OnqkxnS+nPhHvOlftv4Xo0
IO2F6UaK8791t13ENiDgG63+3FW9DDo9Rf1vHrYhBSibBRweLKebxi9Dje+ClNrF
8T9sxt9fEh4kNmddplCV03y5y4o82zBIOkeDSE7pHx05TQ2XPqZo1W9QtH9lCr8C
8DE4WKwE8tayTYvTd8/UFzzxUeC1kFuaraphW23uCxHh2/17a9LuD2HgG5EjBKR3
7GEDh7S5dIIKOFiykkDUO+UA0OG0KSjPs39a0YZrkTn25f/IBAK079YI/6+dGb/Y
el3MbGW8pcWrzWRZbd4PPKxuI+mK5t2S4GvEPYyRkhkORHzz44J5A2JPxzXr6oas
elfRSrdSRbLW9ExyhCy3TCjEZvhxByjPHneQXme+388uVigkWbgCGOneIhymp3dt
eEwYxLPOdZ11wPeX0dueaUfT8ro7x8kW57mkh3xVkbjV64UBUZDnBF5aVMCGf4tw
XxBTLzcOnvQEoe6snOhUC8XvO7GMoJoMUbkQRcfLpuMeECzIFz8e1/tW80CYROaa
2RO6kfKSRlXwAUgj3VJ2Kq+JV8J/JigqVXzJCmHIN7BMsSbz2QFVHgTbTWFXx8gm
LtoVq6otNos3P9uaBpcHIKFHDHN0s9zHuaKfpJKQu7Hz1kgxGfneGCdTvY7xm0Ar
5xVEpeBVTGI/DPmFzzm5Hb6ktd5fhTha5ztwR5QM7+KB1dIIO/fydc1EmNULBuIT
34XxGwIPka5YDF/qV9afHxNeh34bdiVnpwr5N0zXaVfih7L4IpQ8JGZgYeVDR9uJ
yW3EU7L7a16LqmTc9Oot0urqMvqQut0LEYmJcGeXV438EMGnMYLkkBbzEW5SCNfj
p3p5r8RPZy9XtR0c0TixGUAcn+4Qy9F0ItX7GuNYBCbchmHeB1D4bJBFoTH811U+
Oi/Z2BcykI/upLZZN2IwlnSDhatv2j4iM1pxKZfhBg/e1vZOC6YkLUh0mRKB3Euf
B8r4gDE8YjBD8KdMvsnenKH/Lxr0a3w6O1yx16bwDHXlJ8UDoZbaYlqrwzNt2mHS
PreNtKYAd6gzj2Fj0MRSzyyv9VySqc/dMmvwWGDdsI6p1gawrfXLd+y8W5kTSURc
KfNfV8B4qBoI83UShrGcwM8Sp2v6b1/rcvGkCBcpPRraWkVXR1xK8YWSvk0ucRb3
Xjhfyyd+zxSkR0SZJb81/lgX+1RQyKlh9J6UMG051JD7lNuSiG3HxJiXNXDy3q2d
BcNQFAMUGWMJ99I3hi5OI1bhf5lLnNY54CU9PQafjarxKYAROJP2V/AseJrqfqbS
GhDCMH1eemdgmQdDX8CYQxFcAyY7x2/QVn6tWrYgrWRxDB9iLXJt3XJ3w11N3UMX
f9k0qHm7+K4kXIaqJQ62qclwBvx/chVmdJ+HjeJbVaucH5IW36NjL0VeSg6BlgpO
OOhI1rLbHJK4V2p5VZBfxtvKWZgKPmasEdsJKl5zj39SceLodelmoiS+PGlHj0uo
zhiNVCU8siQ7TVfSLJgWPQi/K8euZOkW+9ucxLHN3qeDSx1/wKKPBXKZ9hOWjGMO
CYkzrnxecQDM4fijKZBMffo7G/TwldLuUusOwOpr03qvsNhS+u3OQsCpmQEB/C9H
8mCny291jLDv7qDiV5su9ok0LHOCfcLLqF+PN2flEnTf0FDDIBwDtgT+11Qwa1Fw
2UbIygWfsNWjRkCDM7fVKAyIKDGJrMp/I8ML7IncXokuDw5jRRsdG8RfyZcr0CUD
GDpUvdyESyyXT3PEtjhXqhxfzIgdXUG9YphShcM3lhGiVQMIPRsPROVw6C6O1VfZ
VoyH5MVfHJIi7M+vO18fQ0LFD+0ACv/VO/6ZBHnCsP/P7yWAWXxC0Z1ahKy2vIKJ
RgSHPECilEki4gmv7BOEw0h00AxAuwiqhjWtKb0htgJy/BX3h7Gng1WHWu4BITml
hSiO6okitNeH1V/77RWk+2h9h2Z+Ez6JbJG5TOZD0E3Gv36CdnqNj00dm5tm7BIG
Q3z7CtIlSCczj5N0f+Bi1BQP5To0gC0YOpHtP/Eu4GFOHutR/haEc+nVBRdoznaE
84DORawRHB51wydgYcAlDTNeKRANYTiHwyEUMkj8WnBJLtO2GyA/Q940hvaQCEhw
D0ZoWakHYDw28SjrcnEMAMecuLhYWta+3/rGF7PLpSmIqY9vG3PynhuZWobb4grx
lXRwMiYT7nQEH0Z0CSS40QuqEJDvexN1BJumbSP5btGIaISQx/PR/3tDZl5kZwIo
qQcC/YRwT/da5IGmFPehgo+9V1ewGp60xA+MGuC9HYFG3pdwjXHRXL/trn3YQnER
KIKXSYme/u3AqexPl7uSn2PsXwB5uYdw79V17uWLufk11rHtgrxmoWDTTRW3LlbQ
lppNnoT+mmdqp3pQekZMr8C1GHQPIIGBTZJyX1O4WkEeUo0+r3L+SE/AgP5xNelW
U8THkZVcY3mj71EmgbXR5N26AxGbAwSwn+2udZYSlSZEmYfV0pCWc8cxpZwlfoQR
wGEC87A9c8PPYO9KmdP/MykuIXXRTTS1+gfWHA8bdZDhHeLOuNUc04BQMintg+sw
rfLsnjLiyLGvAFHv4XWdHVuPfonrB5zzhIx1YsctCTOp6MWFl8BF5m5FJikVRdtl
g4oHsZha8TFe7s1Nq5YwQDx8sVEm4sQEsi9bcAbEvbOajHgozacInVjT6r16uxoq
0y2PqN8IqpjCI3chf/Wl+b6td+cBPKvumrgd1BXFKJsLrblWxqaRDWT6Qiu315Aw
4nBAi1cdm23X0h3OktGkyk3GnENN4161b/b5AZ3TxCMM0Qwsl2Mf3mTiF0D2KIXl
DxqFvSHvleMTtrOmFhyaAHShKMxTeQMfbpmaMhOotQ7mS+JoQg2yTq+5Ay7yO4i4
8DpLT84EEFVOpXgCYi93dJbDp4BnxZ26rACSLJpTZX6IGU7hHlIm4Ti+Ok5J7RU5
jjxd1S1Uk/1h9WMVPTtECt0STjAvzMwSoDxVwMzQmRQFYYa1W1BTebCY1j0o6GDN
Md02kWrtSacQ6EW2Vl60w2Qvhjbll8XvCQfrh6dWq6L+/CBHDcatqYTu2Sgl70KL
KfYP5jjdoXVuK/CrDj3D8jGU/kSHMGIPe6o4Gvb6nCW/i6pA+3hLkncJX+3q31n8
DaA+OVR9GYHcbq2cjZQy36hHkvbNQcw02QTb6XxbQOaeGkA2KBVv4l3otDg2CiXc
7h0fLCNzsgiL7yNhp/3gV4qn2WusTMYMnhaqqk8PWylkrqjBLAlXAxDTCJkUy14E
bgPCyJu2sBchZnqmnHj9zQJKAH1qvxR5vD64ltZozq3BY0aYNNh88sSjI0J/zz06
kuTU8PDIQKdD0XeP0vw4jykpe3cSoihmWO0zToHdKOnvLpSDdLkznwt06hAKus1A
XEPLTqIImQYf7mdHMUrdE4vVWP+DOOEQaM2+dWfp0WGzzDx+H8qHQKiaDV60EOWz
YEqwJlWaw5SbUeEueYvAsfIouUP3vRY434Y4uvUeaVYBRl043cw6j5qKWN0FRxvB
PuKyf5/r+db4zhQP0KrkqmitKMB2sx0oPn4CBBxLGFjVSORD59sM6V9mSmYpwpCR
PXZ7RLBzMkYUlqND76/U9V6NSh638ohuDX2prVkS77j+FNYS3KBOA5iNSGIPf3nE
YHcm7yVh54gEO9KwhjcAsSqzxVfyG5xarM4kIovAH+c1yqrUopf7REyIrMP9xUGl
BrdJGTTZwqhCjHBBLoKLGmwhirg0Bxx115Bg8SRh0er8Ck4u0M8L/fYw/75oEG27
8h4sGpUDPdGexOYrRbop6JLmc1kMHIx7eMXBLfh7nbmbBJTEChkJjw5ze5w7XLoH
QQWjaYMjOFLPUmmQ9C/7w+7pGFBEZfVYnzKg/dYN+tsHb8GUyk68Un9vjiaZRDUX
iTpxcWiNe6Ae5x6jSjygF212+qzJnbvcCF+E77AtR258Y8KfIo6HWjfqqHfab6hS
3BpEabOkiCf/KPbKK5AxTzvlf4tw5oy1IIBYJNpDY30xOw1Yy3qIJ27HiEAwYB+H
deUxkC+iE+KNSz7XL/0lLNmFkxPehtjxI6U7r+9vhFbAkSk1L/gBtXfmMN8RW109
t1N3DX/k5vHWNpRG5Q8q8OL347rJMIM2V2Gnk5w3QrS16V69X7dMvB4sRpD01s3D
qUOpr/P4/8cLCVmW5Rias+TAUEr3bE3hTHjDh6c0I/2qnH92fbJBH66m6d+pPm4r
bky72YYv5wkdg7qHTnoDgxtUWZDjlgsN9lE7G+gpJFzZ1nWD97cQjdkp19jexuwN
fKE1HOkCK8H8fPimoNnQkDcgUJ/eIL3EgTIw3klmtvFqXuHmoDy+C1LMxHf9Dmdx
PIIWno1m9S2x+xQqISjoaorFc/+Ipnw3yzWw+Vgf9gZz1W6Dv8HqAs8Px3i7O4UK
Jo1NuZnjZyS6697pdJ4Nam/XC8wTgERVHIBp+W9K9enuWJOpK9zUAuLaILqkT16n
pgDLaQn7pygqP/5iehqivX2hOoz59n1/xtX+BWxSoYDjv61Q3OZ4cPgKzFgWewO5
2OaybvB5xjovSyQYj7qft1dvFg3G/WKj4a4O3+O3/KZQUJRzJbDroc6bWarIMNqC
93ICK2BxFOQt3hGRMMIt3OQkDNtLxGiCnpbCfbR74WnDHiFnhipHIlHe8fnLUo4f
EjwogprAvrmwEpNByTYryIw1/aufnXMsPCKYCuuRgV3wdHiDR6tBCBPGzg2NqYl1
qZSw+D8g1r3WMxj6hQmP6Q==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
SvYSaJ06792FrabQ2cMshN9+6SmQerDjgclgIs+04l+VpN/9yiyaADGxghy4u1zN
TqcWbBxBTBrQkZUcI/7TwJ92/70W0dbgz5kyaviOzTOspROp6EwPs94zcx/jldMZ
36AoPAPKywFivUYU2eNhKI5BeVM3Etry2XMLU0rkLepjuVvflaYf7PD7qNnRP7ii
nsGkd2c2C1l/Hrvs1P0+E79dwKb4ylGmbX6yiN2Jcss1tRgdEDNRWW11KHaTGQN9
ZxVYkUuugdpd/kq31One/6rZQBeHXjqqDT0Vls2bqocRLaiR5LCDWE+/Pdfx4ncC
yUIKiMZFu2zuDHZQlATvkA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
mFrVJxiHw936shHJoIYk647HsaHacYFFzH1frGqzCe4XfYejdX4lLaB23xjGGxvl
YYzyHZBelF5lu6I9gAnFt147XYUFE14OPqCf0ihV9FBXpxKX9DvXt7bllc+AoqDW
6/L52nVtj2Ey0yDOLGM3erUAVMWn4f0yvNVtQ3T6ArlpzFhHsHcGu9FGy8AY+xxo
WGJqalWFHpCzu8ZBBeqZJ0Tb+b8ThOOdsvED0/ZHHzChtAxJnnwyi6eCxKaFCktC
Tt+I87dv/+FXOBgufSfJp6vkvhqIAykiGB3jycCy6YBMvdzTyDOuihsH3vtkbTCS
T2x+tvWJ32y2tUkovJmiPidXWhXjLrNMnzEKAIAfYX2Jd6KNK/MTQTkV7F7gwb7l
q4oKjXobn47S8rLguWeX8hBC/yaqezDBM8sbWjIFOra3qUVA5v9ImVRRbtbDUhxp
L8ts0OsowzFUUBVMgftHXyJESizkBHm1ZMsr3PGlocZRhjR0ZOhmAJif35Z2NdRD
9MVgR3QoGowIagx+M9+rpHbcipn6X+HmQLvQAIeTdlwsPX68NHmGPNX+UUehuFry
npC8R/r8HymdfTJPwHHly07gmQwPqVAn0d2OXdMW03XMQhjmHNuGQRgWVLOgRvUs
NeznYmYgqS90WVFU3wZTaNBkJbJiV8gxxYMHAywE/4av7UDV64IL3eM42JMtVE7C
/5XGXilIeklFsDTq3JSRATYFPLrV7LVZ/xj+W7vflxw1BaQftv6ODD+G68qqXBPn
QDtloCnVRj27/GrFZ8dgJYe7/V/KqeI05IsQJePxxarU3akD5ZnQo1wnFlzF6E7i
m+Pjtm9uT2+8lhBtZlFQnRmbd3JdcESeujiqkHXH4CmKNuW5x1Aj5zaSp0/iBc9y
6MSEfpFxYc7c35LAbz0z4AwOqmNZAwTUzR4iAWFK+qTkTP2kjqrDLHf7sxP1V83S
PTMn2BNbRzASVhp81ld30Bdpsg3q3b+KcrYJQGWHMSz4Zcy4/p/nElD7OWJJHryx
uAiDoHe9jKgru38GtpPJdCZf/Rx1zm+3aFoCI+5SFEiU6eWPNp7BI7IL3DbQS5Gn
dGwyiXe/AFgGLoyPeB18kH/4J50CU4SyGrNx+aQ7etrLmZHZ4VkTrNlSP10g5uEw
W5Tk7UMfJz1uM6D8Q2V/yOgC2WU3fRtQZA3nyf21Md4cuoVB/0de5xx+59NXyEBU
9jGy7Zdl9HOkS3P4rd8EIzB8C1XfF1aPPC6uo+ZkRb1gSl6Oo2qLzWf4hvzEKy2g
4oXKzHP2rFgcCzDqsTMCqJUvTdCFrF3hDbD+NF996GwLFHq8kPgrU5rnQRk7cq6O
I8d6hsBURdKaZzby+GVdtD9AWRzmmAqCXie61bK47DBGlg86w8r5HzGvRyt8/h+F
I35Rj33Rw+Z+4/zc5GpKWUPVMjzdm1PnQV0DcWhkl15BJH9f8l6xWaMY3bh3p9Rj
tOBiEg52SBe/lyaqYvUI8b5v0uYJCMQ1WDu9meIWjs4RYl78/meZr4FjhpuHtO1q
gjxeyU4tGY0jwtAqQgUxomvP+8a4/SM4wrofUSBTUacaye5vSUKIz7ESPyDLTaRR
DccE74oB3fF0OC9Vh5UrrFmlTXrfPcGdpkOBmvl/g03ifX9QwntRMU+TwC4AZKQs
bhqWa9d8wDzxhhqGbjbkAPxVG8GP0hFfkSJ1/5GiOW7oGyKpo8X9qZCCfF2hf1E1
F1BAsKYhjO90kfBAlBRIlTcvl4NWfNChxgmTC3WylgilTm3fYN4LuylpWcTF6qts
G/hRlSLXlrY7aODedAskpEbI0Q37EY6Ty04zGsvPj+pi4FWClrvCbN+STRjgs5Az
xg4mE8Up5sZydDj8+vaiwGwGuDEDpJ9wpksfxYpqMh6r4rA7WIE9gUppNiefE1oy
1u+cwyr3BKdCqO8q2EfMe9D7Rqc+JEBG5awXlpD2/d2sJQTd2IwXASfqolCf5cXs
JtoOKqSk5wboGm8STnUSzzktlceqpW+NxSWJzA2vtuUSg9Cb+VOCVxZj0gpahKYj
LVilbBbEHj9kEeqGqKvwVVfGm9YPSMnz2S/xVpTX6RAtljIgQPPoZqxfw4r5kFJi
FeU0aIABh/D0BEbZxhDnGMOCMQDRhgxf8HljJayJbNVrBnY/vp5qv34kgjYZcoKW
Pe5HpKynj01DH1hIkHHYofkKeiPpYo7OW2VtTCWiOLxpub0R4WPfEMFSaSpDY4xj
F4GH+7Ro9orYp99NjqhyE6/9OTvL7jL7e7q2fFvpEzB6SE11f4xbBSS+aS+n8F05
Ow5PjAVWNOfvBdgLkBNQ9gR27Lp6mrsFv+CsD+OlZrNrOemJZzTtymB1/wTY55Dn
iFO7cb25SehDzr0YVOMbFoDKeePN7avfxdoN2hggzAvJqReKYGm0kyMP3EQcYCpZ
UR07td9gGcYP/SY4b8mKO1PRD6jIvibDAE8sf8WvYutoJGqgL/JQjTW8sm4egYCy
yEFGkG8Jqu9AT7943qZLLDArTkydKzhxGcBalKaY3AdlQfM9jDQWBOATbPeSjx7g
nzOW1PwnqmIsaivNgOF1QjC1tkkqvAK3pORfJgbYvsEodwd8glNiATym/8ZwkIrW
3MmhtzYZKwTUpQFBm2r1mlSO6xfrNjQqhB0UtFmiOIDsQwyE1v8Jp/lKS3ZmE0/m
Sss1I2qJLM1tCuBVFYcJYrweuf7WnqqiBw2ZLfAVt385/4EGZorwVZT3EHtBSbrW
Tc3++VkY/GKdPWzIPq8a+L4AwrjNHdbJ9kemYludDj8uYW2gBofE/SYD44VewF2Z
DZ0qWrHAL3PE8+ysOXiD8hRrC1oBVp8i/ghNjy4n6fgZQJxmR6vv8AbnbIbAY5om
ct7ZUaTiWns0V0OAZ7vq3XNFmpCHIAuSJu6egXFf+0NWXDmdwFAp2wGLk992Mt5Y
Mfm/cfR1oyS+x15ZBdh2uEoyEEFVEzFhi4Q5vsTTjP5vksM06nr5/07/MqXYns9E
FFrJ9cZSwymrDHInzcjtE+Nw1hOqhZUCtQT7lo2vvQImiAXdVTgKqU+tvKD96alh
GaA9UwAnq0M/5s6EM0f3RMtsM+72BtM+WCSuQeTn7gKG2l5KOM+5qAdG5lR6sHDR
301qaXZyzGHt3TKdFhec/D0qqsHL78dRLFNpJ1TvJDetCEfgKlDr22gAU7nEaACs
njBgRCVoB4U8aAt+miHu5sHENhyeD/4MfY2iTJH7R4gfp0TDkVFtGjbzXPAQbCVN
RcT2n44VGMFA1AsB9THFMtYEJnxrDvZCnolUDgsa/CA6h9YerPWYnOjpwTmM/U1H
WaMNtKNZ5nNGG1gY1L/BWBk/B1FqL93gVzhAxuQr2ZnDI1OdUqavGHYEzihk+n8J
2D7Hfy4OeL7nSonSUhU39Le8eNTS76DZWRgHPA9MW1UzNCC0g5p/EndixpD7mJAK
tTYxnqaYpO2aNqIFJZKxkRfqNe2Y7PZyUVBWjSjiG/z38Fl9VH2NvZrXvHgSZf8b
ng/IwMLjNdLa7NufMG5mXSukmKBdZX1RdHx6bRvNoXI8z3wkytI4XYqfJAmJWPXq
R1BPw/sivGcdegqh8U6KB2wUvjZmwwys4u9CIN6N5B3K5u9gU7ddENJb/u4zzJXl
d4NP+bJi0PtBxW2urrIWWLA9q8Zuqg5YQAbm6F1Y0pkO4fiKTLIuW2VkleaM+MmO
CkvfZ5GM/X+c5ogTzSQZLmpxlMB6tsuqAZtmQ/7rlx2puYmc/8IMxOOBkIp7T/cJ
xtVsp/zkzKI/QQbmXl66BX3TZJKZK1RYak2gZIpQqb8bdXPMnol3H3XJMpQIN5eJ
HrL+BLkE/GPgBvxtzs/wE/WQV4cfnB5sXI0s3bTfl184QFQexCC3P3RPuvMWOgRl
TK9N27ytxGaWP9EQfICXTLocqJ+67ac+ECunWGe5ETTLHPCD8mYb03eS2P9KBdrS
39KZqQaSpnaazC9s9Ls3ArA6Er7eS6/zdnvDYxF+J2mJv1RqsuCiP3gSx5f86uCI
mTNavlB84C010yZVXzLoT8WlbnwkKSBUlDUnwhUvw31Z1Mlr3ypTh5RL6zsHE9xm
IYjL32xZ96zevFsyCbSOU4sx+Vyd/jhT6p13JxyxdXwYUS1m4voJMGe/aWSzJtn1
o+DN2WYlgcWsDxAk5VHAgdtj3kjInfoivQkmCxGXAoRSiq5aHe3z+HpZas+PKdus
eh+fsB2cMtdOLOzAD4g8LKWQc7wOXG64EdeUkp3AaRXzN8d3jGo8GLI2ZyyM9hUU
TbFPO9nhKrn5IfK6WRIqlYwPAQoLwzgI085U00SQ5d8TMPfJggEwmy65iVaIrj/r
o+iMLbpHIjrE138sHk4S77oWW1d+UC9erLwQ8ajMJqJMkpDeshcHQMeyaNYYLhEY
Y5JGAnqJreX42hgPoYVnmv7ODLLEqUN4Y2zFkYKK3yncBjehtEiPSIoFnSXci3NC
FWGM+Ee+z84zSfnlfB/dQZTMSjWhGLqUp3Wcs/gMvHgSwXEypL2G06nWyO4gDoDk
1ze4qFB/YF3lXCZBIHb86rDraOJg+iqvYyOdoEM17PjqCYrYhl5QX3IPy5DVQyna
jkngPbBq4MXzeVCzRy8wE8CehcG6CIOZzOOTTo8TjQz4GEiZzxukCuHOY8hN71rH
uysxbaNwahcxnbUwxcYgW6SkFvOqPLF4fEYHPZxt5sOiM3foKNXMwoeikLhK65D0
I5wF+gkAFYpMFK6hehaX6dk+L4o3txC3pAqfn+ZK9pM4qXaxJiSYaXNY1VCdHdXu
DTEPCI5BqGrKwfnweAEaVRB3a8qYu3Bzrn/sUsRFHtS+Jz1yr7DjzDy33RRWw/0k
IoWZ/ml7zntjVfu6pbmS7T7M9eN8ag/hHAc6uB81GexGjvVndAWX49HDwex7F3g7
ZLihkfJu78RmAArpRFry7Izk5Er8PSrXKWtoEuadqkU4nU/L7xaeZMB1Ec4LaYgc
VC2eC3nG2D36+grVy37KH6W31aq0/lbJpTKoa6tq6OOBZsDaY4wLek3FXEEP6Tx+
zqheAbzMdDSezhsty0XW7qDvODoSjAxP9snfOkYT4tiIpn79LERWIdcFQqeQwgxZ
oXs4OQ6yP8Hf1qgK1FXxYfSf7MUynNwKu/WpYnETR5s=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
LA8ZqayCVLfTiE3uNU8xllRdgd2v1AaKfori3+oFBKc2qwujjsAkfeY+o9vdB3+3
+lbbFxcbaRYpZtlefKuV3foBNPwFi3IdBAWJkwGUwr6wBGc+QFveRnTFtfUFL9DK
9v6uXRO7wG1UL/axYNN+4B5GfqfYy5xVUALjQymgtIz/poUSS+HfCKIA8CPOxXCe
9D3tfVzCptZXPyYMfYcvMeKiV0nlnKUUfi+Dx4E+i0T4hl4yoQv0cVYpW1SPorxp
5N8FHGEBtfIcByzEkxAS4TaWgP1UXjIX2XxJ9NNQ6l9PWFr6y6ewLCMZTRCeFprj
yHV+8Q4yHTxFVc/DTOYMqA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6880 )
`pragma protect data_block
UcXUefIHzA24lmQ/RFKrfZQdJFQ8uhYIlq2vsnVKInbIOf/Zb3AsTpwPSpx+caV0
KrCEIHs917gZ5vsJqQdmKzl9mNlpsyC/4MnLL3PAPdS3wSsNMGr0XiF7VcM6qY5k
tPAxS6rLd1c49NijwoI4OvlJGSuvmNBrnR9RHQtgaoJNRW2Fu80FQLSO6Wi+fLft
ACc4MfAo1k9F9eSfPOuPYhmPAO84RF4WtabWwvabA0Sxi1vx93hJrtlJEpzaH1ST
MOhXRD74JgYdeLgcbMBNxCRhA5qYtR19hbnwA8Z65slS9HVW/wAjNktg2f+sM6Qz
aG7Na9FHwPONAnKmChNT5Mp0SBq3g8lA9NZyamfoapYfqNvRVCsItLnDo0bnJd4G
AzuQ0fbwZrYsGUAgdHfl5+pcQ1JIILoc0xnR+PwMnyDkyvBq5Sj4HYT9qWiGiGio
Mu5tBOlJ9WI0A/5d/eP9w0bhKucM3xMiJYxzk3saBc351aztwImgMtND/1e1grWc
xco6YINgaAhnISgLfsTt5odMPEyBssRPoYEJRj7+qEsTd9f+3H6G/WfB2nIMoUU4
S2UJbeK5smp1vKPS/Hjlfb17Yo9BXy8Cb71i7nvYkGH0VLRMFMF88QQOt46fRW8i
CfHANKjyBE7+evmOqDvPM+XBrGwKTWgcf9O2aTwxPKWq8RQx5510bm3YKVdxHLM2
GbczRdOJcp1winMJj3Jxwr/7MNwvf8IhbuUN7lZsIIDgT1WZ3U4eY547RrM+ZvOO
uC9penl/sOaDKKr3JihsCJqCMAcFxa/eeqIhbxnOJ2/aYRv7eYgfgjPSed9VL6PV
WlGCs/zTiy0dWAKtucSBRewyukilfEp06c34NIBuR+awWvF7Q8/w2TyCq3JmlO0A
od5u94p/A7zcTJzzvrI8J/+oRCeT1d/PVy0wC8bSt7Z0ErGUgsPUSxaLGUQylpev
Y8xsSpbAXe9rdEiWppn0KqymgF4c5bYCWtVWO5uzH6k348NNTnqQojEsPLC9t+eh
42fthMeHitLJEYGNGGj9PJEeJCHI7GGjC19/7krnhSCFjayKjaPQReSCGj5Izf92
sxxmqtwtzAT4076XY46bWCSiSO30zPrLKgSt2lhcxAgW2qQfRmvDouKnZh7qMn1i
sdV9EJiLpYWcJBlmsAL9Y36UOIUCUXH5XHOBMBf1CAGktLJl7/IVQh36B76bifqJ
q8vISk01L5VIKEjE0D9j4Ak3p455wRt4sOFsWpk2Bod12D0U5rqsnwIxPQMWXjQp
NGrwMwcz9ctdxj5rVBs3hFem1Y+AspgnYhROwzTjSk2V/7lOTJKSmanrL0kiO7qh
eGe6EIDmsqZ4T0inkpD57B6p2K+qaO9Xmu2mZiMdDfnyvsSoyh3C8HUtdlUUO+L1
l5i5zGmI5jRVX8Eg6KqV3IO90+bBI9ZkD80qHbEEAMtIJ4YpG2zGt1cwDpiW/g3I
+aoN/6ZGq6GB/LyyGPTzSLflVXkEv3lg57EQ1gF1DQTkN12SyXcx+8hvaNPDOLlF
nQUMj3TadSKytyaztTlyO8NTI9pYNTfFb8DV+unx7sMY+2NrFVgi8+srzMmn9lQU
cGwimS1jpaX0XP76yybtt+ZgAB/DpCMmurueIWei980zHXQyL7ZumVDC5+yPFu7m
fGTeFEOBLaRnpkQw8q/H30cau1lW432wn2abeICE0CD4eTEr2hFPhfYzZKRxjt1x
Y4vMxYSbIayLuKTNNzndtTjOjy4JQ8c74pshzKWGmVmvmypyWePhP8dsCWLhH3P8
Lpaa+1Z2dvIHU9cjxzlCAg8iQ+3jxg+C6fQTyvNsmwW6LWPJbN/WwWYQ8DwibvIs
obhOiELqErd1svPhNbcymsO2VaDNqdkFSeKtmPpJtBp6ngK9rICJLadckBvq2X+6
LShjxPK1PN0pyB791ACDW+781gl5nlo+PsY+livFcVEeLeamJQL7v8dyNtosUhim
xRi905z1+Z7n8DH0wjGq8mJf/W/qMwtTH6Rgv/3iHq1HEb41i2UaEy1ux+yczG7b
15fNraokcvnpFUfGL1PamY8m+9EEAhD/BHmsIMvvBe0Q8fKkW29b40Puazlj+kI1
S8Yf2K/sUnCOeD0pXQFO/AKORsKSBdFEDyrMWWynhU2NT4oaZqEkZIeY3jI91Znv
LAu4FZArqK2yV6UWr/2OPe6O45AbSkwCwRoQqSTnXxPuoHbSIXm5ujuM/KYDaLKF
zYQ/9QWj/3jOEIvR0nFML2KiZ8LDtPSniKrRV8F18oByKyvGyQukdG3lXKJqHMzB
OQFwp+3jrAvmpX97FHXPf/M0hSEORdBbVZBmWlm2aUzdSxk4Kz3YTGK/WOPP6XSJ
Vwcr6KZy7rr8BIj4lCTblLKPX6Z2iC3+Zi7eagFudO3zD82IYS8mqX+to7BZa0Gs
klC6peo9D9iOoD9yWGLovr/ow5o51StN8akXPeRkrV9wVYRt656ENS+X0uP8DzFl
0+2f6Bqm1GoZa96Nb+evucIpZzkBWys0k4RRyGT92+TGk5f6e2ugA/ucNdHvrfDK
HIuxQzYtxfWwV8CVAo1dwucTt8RHqNfl9bd9iuLKLQc46qd6gxd75eqrvoIZrO6g
zFY/weLKnjrMEiPx2OIoaiH6DKA1ZvD1tQURbCJLJ8XmRykx8V7X8fTjbcBj0Ez1
dej0B1c3R+6g+Gf7Lm3jLAedfM/1/jXJIW6kveQ0m3rT40vfNo7Y/Z7bX7fxWDcR
Wg59gsoPImGULZLTQVMmn1mB5cysV+Gj3t3b8a3aeq5ri+XKnLNngIPyS9leqerx
q7pykUy5hsGcuP1bJMG+5QnmEmzLn8mGkpJQuVFJc0XfI7CZBo+Sw60yOw66mUCO
Rzjb+0/xQFjG65R8TS6qYIxYJ6Y1q0TS2wRhAbRAztEfRuuKzee4JkhKbzzOE2eY
vOmxqJIU17mhU4yTkFDg/1DUuPDG/vsmm2QAxgWXxGkydhwsz290TXqr7ajVVzy0
UqQTq+ODjng+x4cWePPh6WuXV9KhQUFmnNYiR4Gu8wPUi2G4+kMLvNuzvT+g+Ogx
C4N56O5hHOg0Og3P/JFp4Lr1jf3dLSQ46PWee+npcKwWjEnwqpGWZpN6CWFtK84Z
CCu1X5mGRstgWRlu+PvVXIepd1UR+K2Z3bpODhHUcwvnG12lNcY1LNf39Hg8YBYa
hCrUjRtDgwHp+Dd4Rs+sT4EU5bTdp1J3QN7/NXcjvep/Pqmew0dz4uE97fotaeD1
y4iTIuChiJrzB6LGA1fs0olz+n36i9ByOA3D1Pb08Er9hG7vghrTbBHuox3q46Fv
BTvGzGlN5KTtUA9iIAT8DH55vkPtxCIGXDRXVbExWqnD/5IscOB4Y6kP6/DAwPJu
zy4xuq0E+FjwcKjBhCRlqqjGnx0/eVG8L+7olMxAhDSQGeYt4y0vxzQCCB9Kzeju
svcXyh0rhYtyjc48RH0aYDF/oXz/OS0M77HrvQSBRcYs8IXc8WGZJkfGvDtkkMl4
V4XqpRS6Krk1SNct3Gsww15hWaOztjsiR1zejaw5bhxcm+DyfBmAttYTW6blqQft
vocR3yHsNSgkOKjMEGLsYm/q4ztAzzORIq4ve7gm+ycr9WgLtPZKTUqTIqJC6dqL
LciJK7zZqHgOhNA8GlNrfLVx84T1IskWxicBmcfXYx3bfsFjlHCoV6Y1mDmmoo2F
9oAukAoS7y7vpjNlepYkf49K4rmL54mCXcTCjUtBj832sBHMpobD246JtrKb0Ebf
vmHTUFzlOCMO4qbSwxl2UlH5kiqrYqwvT8wY9AVRpxx7GoxPXk3xECeBQqHzhIAN
mXP9wz2J/qZ3vwU+yZRndSK9oE1gDxFWymJEJ3T6mWFyEYoDp2V1/Vmp7StI3LO/
n1ZlSXzfFNHGod++U/+8TGdx08iAHrLSH9CrLsxQEQfAMvYfKcu8Ul0y1eVgGIUX
k3409bWQs93PtXJzFuRDqKhKWU7bTnv1XPiiWwOAomS6yLcBQaZvNHY2YZpnOzwK
1kuIOOT7fP45bkakBoSq8Oyl6MxZY78Q5+nLWG/nRFymJlrlaUvaJC0nIFjPQj4V
G7RyOVbbrDAdnUmC0Io5qbTqVzwyv3Dr6un0ZEXksnPMkn75kdcGYxnkj34Vmbmm
Zidh3yS4W+YUvFwrM8hqidrUE1Wt0Lg5C4zCkkzJdQlPnlSfrntZ3nU7ZpmoDl67
sUFvInNOX3Nuub/MBw+rvbB0FprOwiZK8rCh9XxHjMAjWbkyyJOxUl0soU/D9RxT
Yzu0SZnvpXAiwfdQt3Bsy7zAKuK+kw/uHnj28kN7BUn1lX7rK693AM6bSDKaFdX5
549YScQhiGoQLbhil3P90ZIwhho5PqSDsiRqTGFrqrgCliETK6Dr+Nt+On2j9Gq7
S3/oC9Q+dFaLiVYJODZvfJAWQFDIfBLhKidSRBz5XMIeRZGLEqj1dUQ86vfSliji
pzp2hW6mtLMNG6eejtuDkqQSGLCCgFnpyjkXJWmebkya8xnWFtEpIc/BMW0m+e1b
GkRJMboJFQKblKAsLhXnZFx0CZVmj+Gka2Ac1f5i9vn5J2p/kGLp3YCyq880Q8Iu
WmhTvDUkbWo4Uui+XiFRb7yd/jOjUU+D+Fr6iIqqyuDPOI2pUXR07VtLVYh6LjNL
4O9c1TdaiT67lK+bl41P6V/6ixLomghUwz/UdNRcBzo6AYzlvaHSsRRVNn9+lmO5
cR8VOCuKEBCOWlYTPAY10EJZgETc8vVkN70gJs7YWoMd8u0jsDCvwEp6ef972n87
uxghPykCMgjqLQmKWLsx42yv6b+WZAQhbShAbHUmPjDHaaUbnhHG6gymukQ8as8h
81QnpMF4QVMoU6WBNaYRnioVIOE1SUj7H5MlbZ0da0ij/nU3DAdKxz5WAVRRVsfp
ETlTq6+ga1xanwwBbu1V/kxJ29FGmAQtlh+nhjcX14pqHLB39SFgHwSON9xiPm8c
mO18WuIsseGl3aAYZfyBWeJSJCOV/CMSYNaNRiMpCGgYToZ2BeOvcv98OFBcqCC8
/x4ZUILRBoylFevq9vtblzc0R/2GcCAsZQmV5OpsWRRf8aBlf7GUFrwce2Hct0OP
YWDFQL9ybWC6CWH5Yt5xhCzrpTK2LIKUc/7TD10uwQ9BC+s1De+vUp7cHoF43KmG
00XRVKbdIJFHkNyDEeEfjInmQnVQkqfy5kAHNU/6PPc/iho7Qjxuf3jdJLk+AFaG
qV2uCbYoLRnWWvf8+PCwZvqy0d1pbk0fJqqFwNfh2zSmmNBNoeczx3aiw2ML6KEK
5xd83WMvQCOhklo8C9rw/aD4KMr6mJ6N+0xjKhRgpiHC43nJgLYMRaXAQRDH+QSI
Ad7V7+fiQ94ZdOlMq8kAzIKaB13DIS2MLGAAbj+Y5xPA5TdWJHR6jIw6v+YaaqpA
ZzypBelN+S5uTDy53XxXAbRqPG8twtFcAHChcxPztlWGSHFsIGJkhwEheFqfuLFF
Zh1D8xaK2xdvaOB0waV9LBlJ6cigS2aUmZU7uKAig8CR7qj/nXr4FeAgTDttK170
nJol0qV7apuxUc/pyiAnpMm2/Lw8YGOXvfXYfdUW+DImYtW6Q8xOoMwBlns3c6Ar
DsEIKo7wHJCSmNf4DTdvZzb7jnA6wx8lJ602nemq6en+YtDSaGNncAOB5e9UpW6O
hlkYpKtRoggFJ42hf5Op3pqXh67QdmvEfmniF71NyPwVnNMSlPoY6zGMgcE2RFIH
EneBNeqT2kDbSFHHRcxjAGPRLWOhDFzRZHHeyzLSRWnoKpBwkSSZS99HSG1+nOLp
pgwjm2DlfAErA2ARnQ9mGs0/oOorVoG6NZBpHruxhOGiWOlDKMxw01eGBv2FHu1t
qKV8vDjKYARkaDm6irnom4hA1jYv4dceZ9EvOvcmaPwAGmNfIQSiYd/3yuw0NcH1
TjbQsdfPMpyOqB2RsvqnTUXLuv5qb84d7mGxxmTJZoKbL43QtolcHYqfcopnRz4i
13e2Io+3rbxa2jfuMOT22/0jwEu2zRHLGwAVkdG/tzpn9t8pPKX1cnVMGWuKUks3
b/ESbkS09YKbfABATpf+3fmZa/MvuwHwG3uJ93YW/RyRCQk7qwTkyB2f8RsdASvs
Uc4UBBxhGCuBsklHa7PHeUoaVsC/F3yEcXJs0n/xyVv5qM+8IOgg1as7X5EjMkpH
DRMrVCRXVyqPi/+mlm1wxtZfIieJb4L48MAVMAxrw2864VMXIFHpzstXNc6Mv9/D
E1gKZqyFELY9TniR7RU2xA8+1MoS54hvzpuI9+z+CmTqYzo0yw1fYwHGMmMKqUi6
Sq67vwztoZvQELTknR+QMyrlvrlwAbQP7p1zUwRDpAuPf2p/Ksl+h7CbagebQmZ9
UJ69P3M93gc5fV8Cby3jBRPMMY+NA1gqED87/fMsoE0A6wzKKG9kVXNKxroICFn9
Hzz1NSoE7MLhRcYnnjBi17LcB5IYgFz69/EWs9jQBYzQNWS4E2JMa90FBMSBjU62
d6ttZTiopT0Ox3YR4PQEzraHQCqvyilUozjCsuhjdtiLl9tsMVlZTY2v+1y8N5g8
X96W9DLfg+4MzFev2vL0xKzmxW9+fcOX830ifCwxtjQMnujYhXqrO3uGtRMCtnEz
6upeQn7sqDvsxiQ9XCC9uXrYJ5LO2q3XPXB5aPtCa2j1Kk+I1VJUTRCREzz+hBMM
bAf5xvxpxCFhnGTVUOxy33x3+m3xHkUPpOmggtbar7zD8SY/31gUJ+VKt0/yFvqe
wyewqeilbM7WbGKIFJPrSt0PUrWpfaB0hoyz+Vibje4ptNBFcQmNSNoVG4IOSXn2
faOnTIgjv5MN/2vXYdOtq2ZMx2zGdc5UL9BgaLrE+vSjSjlINDwcHvamvC8E3KCN
ZSmVdxtXxQb5XL8STXbidUDBgvyODiUqnKKZTrYXB+WGinuAMYa+t7PGV7TdGZC1
9soD/3ZdcIAM7tyDlM5UxKfUhGqF5XHfFtqu4V5otrkMYGyPT1q+CVsojBYSPkJO
I+DFvj6w4temVRRoW+2LAOlsBO5FTacaLHdqtfnOAUU5XdPhYAJb7MmlIwILLOzb
gFvxdPJj5/FXeMIuNrEegJEVQy5+HB2Qoo3t+z8LeMmkujloC+rL/z/kQJHHSE7N
CdVE48Dx69f+I2GsqjJbySqSbTIQq8Ga4tdXBhd+uyhrUuYFDokqmnOy2NvedDF6
FFQAWdPaJGCr9LRbnc+KmT6n2/K2H46tT5OuvTXtOsBwjZ+GOk2ofqSZP3hMdmzk
PGLxiEU2E8c+J0E4xB5yko6GUljuL3k18ye252u6DK2m2/kW/3CLwBtxuE/t/6br
85SSrkqvgjwBkZQrVkwbyflULPf5yidIcplK4VDNZteIhRaueHktzwXUk9zLBYsi
OvD1iTZuYASzGeylCIGHDWpeWNto+gy+z6iyLtTPmZx9jIqFq6VGaY7zgiprhH2u
ngzAZcuOr8koPC6hdfhRQtqFIbS/CvnJKMrHrIbqRZhFvUUZp8pJwg18frXtNL/h
7Hk7+t/gTFAIQ8y6K78HTPRrCLVolEMNMamazX36caGivLbuNONPdtozQUtSwNXc
8l1AWKIyJCo/pNRVcYSafZkhyjpf4ILZ9tZ+nOwoIzxqNipd6Q4G9RYhM7QxSOtA
c/RD99EgN0r3NCcNKQpXG2Ag5OoxngrVqPpjUfpCNMtY+3XwjxDEEV/MZJfvXN2I
CpVVXS059GnHiU70Ob34+5RQgzXlsA0gwS3OkH7QpcgA79dRNvtd2CGmYQok+hDF
zcQ7OBNwsB+aa9omV0bzE90ZBN05LaOIQ9xr674ffVcfgW0MIPVoNY21NlaE4xrz
s3BmGjgNSiRWaMbMhpkQNIK8H8JpGoDTrR5DqkoIDqPYVw4cvrj2kOOGbh3b/B7f
CCJ8oNrHrkkL22d2RYsDcDHyopkwocHXhep1JntH6I09uyYbd+FjAzJyDZm9Gtye
nQQHWcES5Pmoz9mOacAqcPO6Ef1gS/TnOVVHgpVHfZVR/cROe5cW5kcyTCvePjch
mvB+FotVqzm9xVEF8f82wKOBlx8+xBEihse9BOoYITSg12/z/fi2pCQRhBW88UmP
GVPa33IaEQ4hZbZHYYVBLSSI2qgBsAwCptHxe/245lKaWk5wKEjzcA2U11nMZCcO
VNZ9oZ1C1XbcC5TgvKFsTfZ1zPj+NolTf6QGNH7D+6GoSHFzTHDiLRmgnNavEGsH
VXYUj56vxWs3T8tabwJbEbpD1d6v9WYH+rU6ZrrKA7WBT8Hv71MCsW6WXB3Unvkw
tmxxTIuczexu9ORj24yKpqO9KMdrK68OYu7AZmhLmfAXgnmWHKsYULoii9vCwxjY
k2MKlP16QR7IJTtqJ5SZklIySgtlFGabtviyHv33l+lJuTfoOrKx26mSsvhxCUcW
m4ILqWeRmnGCX2CP+Vwd1tnZgU36zBTb6ohtJwpVHUZCER1ioLcg81yAHd/pJDuw
WRoCttaBd1IXeGZD8hQ9vw6j5UGKtDaoDhjAhcTs4B/oiI6lhE6na5k+nuic1bcQ
xNut4XB3+Wv5WdJLnc+mu7hgVcJ429PY9UDf8D1FlwRdT3+RTen2BYee7oMYJgrT
UmAYT9Zk3H5R+7H4YrrSXNh2+kZkRgS6+ytoh7wVXRW1dVAWmJE05zsnqTCP11TY
qB9gegtzqprGqiTiXOBPMmFUCHaV6AmO7fM1SThLlFB4Dq/ZBIq/REhecscaM+Lw
epv5ONe+4RAM8645XtE0tUsE3i0ScaECMm75FP0tm5bHGvwcHRm9sKc0ty6xSKqN
9Lzjkkwv3xqasWKN3k1k+m+QMA1zp22tS4HyCVIgm9kDtMmos3DjxlZSh6qDKJzT
QM9qsU5djC1sjp+ohaAMpwzxZETJWNHx2tm85WVpZFigU2+8UgtLhheS1+sWCDCM
ZwerRO5l7afdKK6+QWRABqw0TxlCiP/XH3fgnmt9KqDgKCVDREkAKdd0E4EMSinh
126b/zAHkFjzwKeModUtkzSOW+SQDUOqas4WivdCLD/s92J9Fq6CaD8TnQX6IMU2
3b2snwq2ucfTSV0qQM7xK7gJoAzXJiGafP9w7QkO4xHFjb1ff73OOn1Lbbc3d3tW
ZMhELK4uRmWTGPALsBn1sw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dnkjT2N4kD+luBPTMddNT/Fbj/mEN6Xh52wrJMzuL2CJIaFxIqy07hnDRwHolInm
GRNvecSer8CQOupDodwKxLK+JQ8nBjRwvokxcfmKwoOJshFBoyDakjGJZ2kr0+sz
4EmZQP4cLTuxEhjmyO1ah3LfVQc7hizGc+Tax1XsaWHNqDc0Meaot3/AwfkvDg3O
tEGcAqrff12h2X6Bh6voFVM4gjkRai+8hIpb/jUs2gSONLWcSKRNhf+vyA9S/d9O
dXIIGvh8HPyXUtIS0q/uIYmCMPdkawLYfC/O0Tny5D8Ln6HZ0iTeOnEe1fyD5qPL
sEyCjFpMAwJ6YkIP8MvSmg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4880 )
`pragma protect data_block
YYoM8adgVzKWuPcYt15Lm6n6LFrUJZrnQ9tqdZLiAuj5a5eSI8/cmKUN9U2wtLIo
rDbOdHYEAC5bV9izqnAmjM00rw0IOksYHxNsFRIuCiHjvdPDNcoJmqw8VXpx6Tfn
rDc25qwWbh89uQWk5wzqSd0IPaohLAVrnMtOAa+hfyRGnApBNGBO7ZTPKufVv256
Bre7H5JYQ0Kknv0IqcBMghVP22BS7cZ2pv1p7IJJkCzuNXB8yqj4O4aNLzCj4S28
Dkw0PnvWzq9gnnSTT/oil67x5RstgRzrXKHv7siy9lqkxhkYFlku0dXaALbG5Cr0
25YSaqtnIijCh0ewWGui/XDJDCZZT4y6J8ZkNx+6Sxj6EL351dqoXO37mHgYlp7s
6snt0g/wi2cIXrS8PXQCytusqcAOY1pTFKdaVktJMXWsplEKRyj2wzEycj3Hev1u
GyCmOlZ87eoSrLsW/L7HYcfKayuRG9+zomLGwvsTg08I1sXktOk0yMe1UVlLAvRr
X726ud1ObX7Gj0r5ia4+ptQPykmvM9i6YIJ/sY9bL8F/IZbi5TYmEShf0hFnldbZ
3rtVwy3YSP94eajfV+ZBamrmCOr/tHu8L5FzTwIcEWwbQdHFEDdVf68nQ8RcSKnN
pzk0wwOWMg6/42vaPz+JFEvWVCsTYgNHjfm2kh+6mXw0VmpfUh9wwACiKprKODYX
p3VsMjMBW9wWs1Iej7Id2Ti7dKqaNungBAdgq1GXKBhE39lyYfTbQ62yffp3Q5Lf
YTuvWkHx6OCyIw2M1UAUaZ6h0C0QXzhZB3OkW4fh4RfiURbWvPhEZjONX77UYD3D
OIaX8jAw7fPXAd6aAfpaONfbyjEIjNyAQ6u2rl4RYw7oUF4F2Zsl4Y6pCQRO1aoY
L2haf7ozz1829QUGt6Z81JXQLEhXqeCF1aXW+UsHCgdYU9gwShZp5vqWFGM4PEMh
tFfzm5oIrnoSqbbQFMOOeX7QIjkwy1fRlkzVpYu/bYTKY8VzcO5GDcp+UNO5QATg
9lD8OVodfG7c+s/ZQI+uj3HckxpiucEEoqWM/uzVxY0ZIKQt8rwvMeDnTLMm1FJD
aesHmy6SetMHwLsW475hMmD9BzS6LQ9fqCkf8JcO1VKkl3au2tng92XkA9ZfIACn
r5Insx3DNEpRnOE88BiW7fY78kL+J41mX5qnf+LWkQYhpsshxb9Yv5Yc5ydz/6kS
DUc6gIdKdwdRLMX+z55jC9Nh3817+xdENSKTWd6rmzJxZn6G73h+8jKVAiHERZPf
MZ0oapiYpnAgNhimHg9CLgHF1a8IKCo1wQsXB3tHomX3mlWFJRq18UV+Fi54Igw5
L39VIg3e7oefnlvLO2h7mIN/cJHkG0UmATMQzUG7hu4pcGefadDsH99fUgRp9OFK
G3DQWOKu7bLqG9k81GYJdi+zD699Q+Ujrcsfq5sFsC4AgWQqxaJmOc2LBrVl5kdo
YNeVhR2p3zE/J/EtwyzEekHBjc4em25MZCanjqfQSlta2ICSKZxsRHFLhuwjVFzq
pNjY+0YtIzaOyWYjCm5xd06mKvvRa5jpnu7FmWFuz5MeNHU1n/U6XnFZvg7hfWGI
iMqu1ILUXhTyjTayt9rJ2NkMCF0bCBChzK+HSf9kg/tQNKbj00tfGfed0Msknx1s
/Vef5+kN//Ms43R4okjji/sg4ZGw5XHKcc54XofHWwKzbwHuk1X1ANe/A5yEIe2k
DX9pa/fU0vZ0Om9xizMfrhzE62BzjIeMXtZx9oyALyCrxM3EWaaxd+oZqkrk0yxL
342MBDny31UKL3HACg11RWfCcaAXKQ+KobVBLJs2CXiVor/Xl/aq/5y+ELo2HtHG
soX0Urv0miwJnzC+QYBrh4vZgRCmqTsas8xS7BupjymkRTZyjBNqgoIKKzXRYNnF
hr7JzkTEmXWLa9McLTvakKTqpVNkG7vcfod3IEZlGE8Neu7EctJUBR2utOBhlEqi
RpsyPjzwYJwPaGaXojqYyH8D9U2bQkpSYO32nsk0QTEjZnU05U2lmcBw10TsI2Fp
eZfz37v9uu2pO2eaIsL2zMsxTIHl/2F/blS4fM86vpbCttPQM1BAY3SiLocKHWhW
uUJ14E3lBeCT0cejvighklcNcVc3cWWZ/QstDo7yClJxXRz16tFzWan7zf1CCApm
9aNz4oVIhOtQjjtwnMpufHfDsOIP+V7WEmjDuNAgmj51GtJdXBzP34CO1Zzq9HTr
Hc0V4dqsYw5wRMBxAdVZvdp7BB1s8H+3Q/XFPp5Au4dF+ExFCSNP8LrEDdiyDc8X
EfjaUrdHQT8JHsVfPk2Eht2pG2hSu8Oz0dSrMpNeOPHZ9P48bngG68a2h/Tq3CnM
vU5YS5NKo29coctWDVPftbPl7uRboTobgnxvfRJ7a4OPaxYdiamHysk2I8DrIv7f
5uZbQWTT7dvST1W6+LYG4ncoS8sWDXw/b2Mhw9nSQlDqljxvuO5WYxb1BJdYavxt
Bjkpxe6syGPGROD8vsIhaVqYeFtaTc/Ky/8pFjQGjjfE9t47pcBIpshgKy6B9kjG
INiHJcukI+iIf6XC/TFQtLUCwzjkzX6wxneKl+pIa12/uS4/2fAUXlHlm7h7nnBB
dSGvtAEQM71gnOkQscyTnm72pEzgJW+CePew7ovrBlPzpf6pgFiKipuHDjb4F6jc
UQJtOaXLc7zTVtaCalR+EylyrTU9T6Vzvv0Ym5HmJuIgXMMybc+Y9yKsZu8pvP/L
+2sLd8HJ97GIhvxcOlE43Ge2RqtAFVXEha3NB1Iq0FO9EfNdYAKBoJVaK8FNzE0H
JKfzYte0mdFCKL9OlQ7pdKpD0aRLphegsMHmDOaLjBZuGOEDeVgrsUBZ79qHCGa/
pKEimFlKs9bgCKer1hqOR/o3pTuE1JJPpEDsat9HZcM7MRh9LNQygi7catnLTXTE
L9jANxyHOkIgGWwekSe5XgEYA3dTJXomS8hO5JHUnWFuJXCKITP7pP0fc7bcLdGZ
BUFzeGokc6c+24TUbnO/ZykJmLWZLd5OvpJNK1Wq8r7wviyBcVDGULyK4twfJEYS
YDHgSufaC2WxVyB1+KzGRsXjh+C6G1QeY7AbETnZtmfeEwe8vcFlWJbMaW6Ss8lI
Hkajx4tbLdUfyR4Kfg7i7NhKv9j210qrnjZSBhl/d3LWv6v9mg67F2PyfZo0LUwL
ylucYW4KFwg3kRF9xsobzz9hZWNg8ySk/BpF5Va4Y1tSkuMrio37P/9+0GYCl4Ol
B1F7+9K+fr6PI9s9tLPouFl/4WH0cXMJUYW4AqEx1DIMewOvTjF+GStOMfyLWZWS
ETT7LU1SsYlkMoUChblsF9pT6JFckA2EBN/VO5figqPryKaMhO6xD1hxLRJA+1w5
vPh17mnq7P/qdZgbZxUUd3YMnmEKethN825kKt5/PdyEVLeqUeoz5UxaIH16Xw8K
hXdBn2Qqup2T9Ubgr3/dj4ea1vZkGaTcrF3PLifGK33V8DLZTamc928geH1sJXkZ
bVrOjtISb0CtjvdtTiKbBtdBPdPXyYXjNubbyxvkZRYpiY39gyRxG9+JDFke8UEx
pqzu7rOUBhYBxp27qlGRzzFFPp8vTdr3jXLPctnfjgXr7RE5lHGLDO3cOD4lhMrI
lAGi8Yrse+IdxsCNhaQzlawBorRq6Vp5inVK4KLiFq0vnUE8zOI//jeCRLkgSR/K
r+zxiNRyW/MnMmXsSukRq6fYhXawnvmiTRV7IrUx2aTToTv1NQX7yX8nZqPjoiNR
TnPElp2nAbJugZkZMX1VAZAsVZ12lpwqSDoT3Loc04bL0FicG8aGgNSZ3KYTB3ox
isPcQHyDmILEPtK8XUHx/bH/UGEC2YsvbN3EK+sSFCyEhGmEXk37XG4nh9cL+F4W
Kg+OamtCKzcXlyC55/qtWAtF+SBK6hWkb35kz43zwJOqDekNGamUtqfxEjqbMtXD
J3etH3wAXMSaSwqOqR+wOOHjCZ3SU7/q4ceT4a+5BOWi12CnCoJ8evwPH5lhI52n
ZBlOEFsTPh6fToKZHNbX5EMatLje/Shkw6UcG56dnUWGw50BlOmIFhRjUKG09QhT
vANv9wIVAP/vecc9h+F6R/w7kE2ZZ/kI69M2l70oW61Gy+ptOKaKFX14jNWGtgKy
49ZAq7GGmF5kXYFA1NjqLHsDNmtgFxk8/CLhR7pb5fYZcXQhA1YJvd3Ce5nOtGbT
kXlB0nd2NI2c84oXATdQ7Nb0ZvVTV88+ew9wzy0cdGc/ejEbuxzFtNqGDp8lD5tU
l4luwW9FgKTDaWzIQrA8qtguClkfeEIqX2kLGL+yc5GH3fNasUL1EO7RGuOJMx/d
UNn1c0erq02e5TYNwl4sRHAU3iBHO99jXoLwjSsNrdLVtjjWXg3BIChciUfGZKmT
s+0OF8/98NnDRRw8aZxfgXeIMK4TFEW0vvBAnJtRlFwYTNFse0wvjn144mIWnbaZ
aUdjM368mtg4mtgOgBXadAy1Rhv+c9CXzFDtv20tyInpBBb0uOReUohmEITai48c
8dwl3FOAc9wiiNt/duwhMZvnlOVNpU/n8JCNP3EOr6E0QqIZ5mQHOt4moGWPkk+d
ufahw+46OtzfVi8/O+IPyFnSJNlNKk9j3tb1ic0BE075HoIFkVEr1kadQtyL9LHG
YO/8sYDPZuIbrRuKuFW+Fn8Z+ZWSutqQefDHdmzSpx2Jz9qryMlVsCA3zfeFLKo5
DJGJKURn6oLEiAbJjeiontx9jGCzkdmflmaRcTducjHYuMqzkb+wHFo7r8volmq6
5CbKae627ykuHmcDwHqDGFUzySEo9rwzXhtC12T22pxgnjAbjrJAeIYRrPN0xOvB
3BA08UmVxk1XgqGe+1vuiS0muCYMxwcbCAYR647jcI0dXjS2PFNgqhfNKqL8rEGT
+93p/MSj8tqGOPSd7l9e1vnmS+4i0n7U5JBQWVvCIS3D15CPiwMu3lx0xN5Uw8pW
RQGbExcobKbiWmSjVoLXhNpXAdx411FBLXZq9FwlCdPA0HvD6WSU3TjfRfGt0de8
TV6njCv8zRECfTz4zXyrarpe7X0K0LihfK7sy8RcTuOm2b4Th22NFYM+DivHUKh8
BiIw1cokuSMQNJhWNrNL1l1KYOsE23EuIbl306fgQ5+6SymPoLWuJKcqw/YiDrfz
jloTmo0fuaG4nM+fGxRlPrgV/ZstLLJVw8S7wM1qKaEX++CLbT3rcRYCkPNgcLkf
fefM8QipDnc44Y0jf2gpbNoyhMVtj51/RqKV+5IEBVe3+BFstHKogtDz/n2hr9QN
CvieLVO5xHf/s7ZvsX6gk4ducJpmKOEHgAV6E6VThVpTs6LzAcS8RCPgvW6t9n+Y
zYjwngVNq/vshEm27xiMbLtz/lFhzMSjuH5q/ueaTcA++ZC6NLn72dP/LX9t+eFh
cvFCSAtorONExKnZUVgzGVdotODw/0JBN9t5YokMDeGJWpa5HoCbU8U1EbAIOPyg
VShdJ8r97fGMHZKlTeV7oH8zb8r0QtQ2j8p61dyBPAitudAP2uFh4gjxkVCIuf78
UEMITzjDJNcxiwcDS3CxQK9QxcoFlHMFYVNc3fYSCqJ3zGeYRTXO2+cgKmDpBspq
WUUbSipIg57qk2DiFFQzzVv7/q/XWYkqOGVAYQRaHYGZbO+DpJUXruNZ/yt5Fjib
Dn2CwnpIV5UTQt5xIS7EDTB2Ca20hVp4e99/CyaBsEJejEivXJzNoMbQOoR6a6Ct
na4hioBUpI4vcJEP9sSe2KZbKmYZ2JVD/Ij0eiXVwir4fBieIg16mDui2pVUU9AC
/y+JOYUdoVgb/SC6g+CWxyvWzIM6sKxDRKNngFM0PnJabq0h8SPXUI7e+p+CNnuK
lVGHC2o5ecxu46ABrM1fufHK3mD1P4UymqRl7ThBFT9CSnfOv6kFFGC8k654N+yw
pNqhPdrtbQT6yBuWWvdVpTiDKiU4v6KAMrvANikSCiLZWo+n94OFukGgmVt4w1bp
QRVUBUW9EzwnueS9pSJjoKzUIYqsLmMs3/WK9KoQqmIz3YgPYxF7o13NVtYeaPKm
0/P6BS9kEpgmtR1KZIEKF+xMAmAKMPBAGKwF2upDNxU14kl2BMgIhkD3Dyu2Kp5V
9bqRbc775Lj/SXMGqKoDd6My9ODG27uq8oA+hjrgSya4VkAsafJDwkQvt446JawR
qbgpXDORJ3JxFRDe6WSLhFDHPkTMM4Hk3kV1sRsavxdI4MzSTH8RgHa4TR3VpM0n
MpMDs6qdOV/M0uVc1ghm0VfAuJgxk9HIz1B/n7QiWm89d4flZDr8QH70tdyoel3c
bpS2kC/EjccWVRkb6h1FSmfeOIoYKeCH6VtWiCQIcVNCmzvVxZjs5HxokoZvsbW6
7AD5QIp869UvhwbDKbERRRWeghzTk3p97E1xEPZEows5QIGMWDVmhOISzFvborpp
iT7Wbo2gI1mBiiaBvnp7klrMkaUwMIQwWtpP9NothC0=
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GYM7s7tfiagrokvO9/IcqolV6hU0sIgB+wdulCd4z2FLdtKGoofHMqZhLB4/uSpi
/kZLkP6Dpsw/DCYPPsP91CrtG7fsCmarX7SMweD2vPOdpxgJ6T6mwMIJve37fSfx
ZzOKOBd/tHfIU1ueRydK1weTouyPnJqhmKSOzkJksZCJofXHgA4JmnTKWfDx25jB
aKGV69sskPRlXp8dVgx/jtGLMRhS3kwcYeQj0b6++8bgJn2KgKbouvFF1J8TlFGv
+5/2Mxgq0HBkx95tvMrKWogkGAOoaYFNbnjaQ2MuE5uCx0OEM1I5fyAxWh5vWFio
cryPZ9/k+ZtAQhGp7GNAiw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8992 )
`pragma protect data_block
KwDpO79Dg/vTFGzvAMlCCffKlT+YHeHxenY2txI21FciZPEdgStaEavtHh5X/7+X
UTXHYijuJvzD9YpRzvnfqM1BJJd0sux8GdrUtLvSj20SYlMJg0s7x2dSUZc7cSC4
/DO0BmtJWaTKNARogJVfX0JpK+VMwJcD4/lyplmhdQ+wIH0kV3kX2gccSGIr7WHm
UtMDiQeHSFpkWI8MKNYf7aKcvaUSDW5/pM0NvGY9TunsQ+BpEsaLta3FOK5QwJKH
d0Ps8PtTd7rfCO9F6720EV9pS+ovt1pPlEyPY5UZ63tSPi+BcsRbjevfCpupX2pJ
2M7mL++kx97yTimrSZzSxI2kyrov5x624oCvfXobrOds/gUboqz/xs2Y/+NBOqZ4
1Ep6ClhQqIeauNezYX6vfog8H7u7DzjkO1LZKPYHXXb7CyZmLHowKTD+VPv3O8rB
fjuo1YP5ORa1LxDFhqsYo/VGVofqUre47U5LQXEApHvECEmwAVEUoO2+jXqQDU/w
fKqX8ac3v00gONcQLplGannuo+4S+jG9+0WyZYIvO7gtSj14qcpjX8+95SQZOcwa
qOcqmx9WWaCYPmU6TA0a7COtLIABh7qhSVbGUIBif0W51KDEsIaaVI/FEJijlWPO
4n1Z11oC29RS/IDI71zX05SRl2ESdlF6Md6Oq+7PQYwa6OmF0K2Vwq2CKyIA5abo
tp4lJMp7HfEAGU1TZaecAq5CyjBVfZyCj78AjiBZhcrKBs34BgBY99PIZfPxZvNV
RC2IdRbBHwtGNUSTIlbwzPXvv3wFm9Es1nMIV/k5SyHDVDiccZ7RXBgD5H90vB1G
KKr3G65XgTChsIQJUJoVRDfvttBU8joWNQvn6QOSMLXCkR1l1vw7RUD4MIsFrQ8Z
bAePZVhKl9VgyYeBwVCQf5qiRrWAQggr1r0DQhMpFB8YznsfrwslXuFJpDdrJFIy
1YK2RTRZIcl5FCbB82jKrkpX06ifMdlTNmka3Ae2ki2gKcYDgMLMeRLaVT7CNFaf
9VED7Oe6b3laOt30D1AiHEI67DifJJQ+Pb7E24+WSiZFj83Lj8Tp3yD1/q5bn8KD
1dcQxAo1AvGB0U0BKLOjQH41zrBSYR/YdJIYsCmoT99Nb543YfSZyYmAGMEqtHKt
BM2jqAREfe6GsZM+6/DiLo41sN8JfgRrBvLQfWVCZSfihSWkSOIPr6OvlhUKCvnL
A77goqGVoR6Cz+F7fPGv507p2tw8AS8VFKXkdCPkyOScqXWH6vagHRys9D/74xF8
p5wbZXCwzxoLJtYk7N6S4OnOoSNc9p34KNPnDio4peatnJZASg6sT7JN5CIt5sf6
XQs2zQO8C/N2g5PCstWSul8dt42NWzk5C13zORzBBbwNSmBYl8anuV2l16swMjUn
/EVMxYJgigf6mUOqghHFN9U2ldEkOQCr2doseRBDlga1H0gY+bOERgs/F1hUTZQ1
ajst8g+SxoFfPEW54nGH+UuSqokQyQfk9QLBb3L9YqqRaABt8RvirtJ+H32e5CsJ
14XtFFYcEbqkyxzWHhX7MnmRWyID3JjGuc7Nlg87/rmL7pykl3Nujc5TrwhvUyPQ
Z/B1YO8KunyYEr3u2IA/9sNL2s3VmC8G6NNnzmZgcU++5YMqNnAE1X5OtHqJZhOn
f0JsGgGWpPl3Kh065QjCVedoaK+sarWVyOOsWhlEqMCrzAr9UoIvWOW7bfZQC9a8
mOpzL+o+fJvSAA3dM12ePjveBgD31doRA/YsPwRfVtwopmuHNgdUC1bexWulj4I7
hoAuZSocz4+Jr5Qc913q23Nc8cx5MfL8epBJLhY7jSw0M70gf7TZI73nPYbQw2wD
DJxlgwnVRTU4otV2SkN1EedNk8P4S7qcgAYMGKAbLMFcb3dpBI+yc7z451qjU/+o
e/AQSkuwlOIWbP7mtcGLX6q52A+wSOtYCgLyg1GlioHjUXKsbE0WlEP9aU7G5nja
pw0E1M32CKYp7jaRQ9pvp7MlhLpYUDT5VSQtLxMIiVjaRZl9vkhmmzIJc7PrydNw
aPxCIKFm/r3jo87XUfFstKSQblh6TS3Qj/KWocF2/pbpwPh19QcIbNw1OQzzunhn
NkFOzkTW5k/V0W0QZTtSgFMZMQTp9qhknwlg0Z1Ls1sVV1PJyTXvCLvgwtviHZjE
hPgonrU8Ua+mFsuOgYzps4RDHbBphNxWQ0umYozFUvyqwccVgeR0F51JPv5gL2JZ
SoaAJy1/JI/JXlf28kwcMisFaXinoIcMoO4d4YmWqJ5Jpr1q84GDh5UGknpOjSuk
xxOP3J7iPSPwMdoXIPbn87OtSK8mqVYlm+hRRJEc10niKyBw/xj6BVOqo3uTLuNu
NmPNq3dmO1CE5sphr1sYd326Ft5kqpoXvL7bk5acfzn13SyeZQdN24Jfbe8KZC08
wabsi23qm9aXR11E+/QlryCHHtDGYR5+WvDq4/N/qJHQZVZ7ViFvzdYhVdPISTuT
qrpg38ER7Fxa10DG2SePHHEbhRT0Xx6u6I7+zooM9G/zZPQ1JYai/SFBTzVA1Fxm
0GoZULW4HJMhBiZWEe3QaZn74qpcuLuLMOsLayTZIXbVIKTEV+PGxZodPbIhTk6c
b2GyVDxvtP0wuWmxCPNKoGA/HFQ3Of7lBRjydArR3Vhth+jXdj+ghqzQY1tpfCBz
TxABFWsO26MeIPaYbJYTX+d1beeACzwrCB1BjqMatKGSbfa4RSVP30DthiB0gkHK
aWu1o65DcaNANQTqJN33A1oL0QQnhM8aFvcqlpr7HQu7O6x3zkRpcelf5o9VoqcO
sAe61SrN1Su2zSeWU7+DNXlfw+pa+mO8DK4ZEKgLbUvrRWF9BxOFr7I3djZGkN/U
w9HRL8OfxQn1ToRfoS0zkwL3vdMQmcIcCPT//rbo4vLnx6Oz946dPjLTd6HF3XZe
THZ++jCfuMYfW1Z5fyccm7cHNF6qQoD54zMyfMhQ7JMLrbe/5H6XW/Fy85AUDTy4
ykX5ygr7qsVnA64Jf6rOu1pl2Brzab8WX+uCrjFLRM7Qq6cNZg27rI9B1LyG2ZgC
pjm600U1KebyAXaWIuiMhovSocULlGweX6Gsdtd39DUrkm8CKxtPMJaToj5FWDYY
wNdT80bhWtoHfbalQDnYPTkeP/cxfjB+J8tNEXqoU4Ik4Ho8Cy0UvPzeLogJl58R
fMHcp74nov6e4Nt3JPHwu2Bhb1vwWzczYva1Y40rXD9xMdUzS2o8HFZyAiQb9FZG
DxxMEu4P6754ypuqBF6+BgOXYkfY9Vs09C9W2BR9JEWQe9dVLiHIaTw8sF1xv8lt
IXDMG1ViwGRo4mNX0AbeBdoqcRbrdZhN0VHGTfAS8lmwuMMi02Ws53LeZRtA3fjy
2Zjw2scBv1Gn0Ewt/ylfu6F0Dd2dmVG5DBx8o13Oy65Z4ki/jTXPq6u3v55zA9Bt
CMPvdPnAl1y46qi+CkR3sqBNRAlKlSlQtO4M35ygh/VzarUAsdn5jOnpiUNzZo0y
iHHu1tttdcul0YjForjQ2NdJSlHt6cf6zZ06TWZ0K057/ZuE/VkjbseXkKcP4+zl
r7g5l2rcuWIOcGuFMhp2sef7E1bQ59zs2vgVZOFPSBg/00lzjyIom6R8Ou08TCB2
Au0UclYwhXSK27kMx4AgL/QLzDq7/PwIHtfkWfIf0iBqT0D3Iob+dwFZik1ccGe2
1vRwQJ+PDkeDEG6CfU28mYmJAXWWbMVnRrfUDqy/yrUeGBljxX5tyyaoiOv5m0j6
uVI3sVfvB91E5bCKPujXCBzHNX7UwPqfNe2Pu8CDJaHE2cc9T/VqwhnV00+zAssM
Su1uMCGDz/B0YHFnOK2u4kRQV2N/UykZy+kPvafLpv680c+TD6UY4eoN6IjgIq5n
eV8SHs058JS2lkB6IC5zVmCfvz3gv+DznRkKKw66hIUOrvFwpELCX3ic5xQVoI9m
RHQyLb4j0WqofaoCRzTKVbi4mCqY0RmSUOW39ME0yHXbd5ta2Ydh30pX27DExNyf
4WtYxhR7Nwf21Ui9LpokwQo/Jk7zemWvecA+J4vAo0KtLKTnBNxgVIfC74y3tTgK
l7tDgfB4P7vannCAJFDusJCgoTE5di600wo/jqLqUCGfgwI1UJ0OFCJcTz7qUXbu
+e5iwiFirxJ2T2EHV2L4S/3Ave7utlBftOUZvCWl+DqZPy7M15zRDdNGle+y7vx7
ruzWsUGSTPaAzSs5pPRCXxjVg2oTMMvzIctgPugupQSylvv35veBJmudKwO9CCxa
xVC+ESl8C8lAshXTEB4T4KGhupPKwo9396O3mvLudd6wRDJoOG/84T6ZuP7FS58k
Lnv6MBKTz3wqzRs8ZaVa4oUgTllCxaKMV4glSq/v96jqQogyrzwGSt8uYmt3kqSe
r2kN/jhvFjCE1OCvDVT3qwQtlqtgHDJZL971h8T867fMBBb1q0ag+4VpkH4UOmM6
vmvTnbw4C9iP3/iXTZyZO4xxEVdZiVMdLyrfYgnmVnht+w6Hqk+AJJDNJv/Pssu8
hhdBmkapKEZWn9ZoUkQWa48lQmdeUT8OqwZ773tXcZ3ER1jFhiCT58l1wjTfjHPU
b/Qy+MUe5AG6qHKhQgpCVgcNMWTX3SJ5IDbtev7PzbUrGJM9ZDs4eUV+7gcFjieC
cGKSPXjbDHndD2pBsODoJCqfijlwaNUfepU7SdsrB6BDpjncVEfjWs5oyMTnTRzk
qxAXGi9O+VVka5lCyIuu9TA7CVtD6qZU2Dykh+eTBjBePk4oU7XpyNLV8BjG1W16
BoODorIiqZ5x8ICEiMlOalaZUgfpOTOAPj7w7rSb9ZgLt9sdtVR1VKFzgef6lcr0
uHiCdEcwLO8079YGs21em4PCszXwchtRAzoQ4sxRwvb1Cm5vGPrtJSn6oOs/hlr8
fzSAPRXgq/BNZvObLF93CL0mv/uimaxdb0RiVdHD7OyYkGgmf3QGABQVNhc9OyuR
gKDmQF/09gUWY9FFH77onhvD7fKvVHGulG8HjM0ojEUILZz09etPeshcO8JUO/Do
hV96pvD8LR3ZqVCNQA4YZpffdif/EDAjKk0BBmc1CvAdCavA4zkt5oeYWSjCSfga
3YIU5FOHoU3XBayTyqb8MsZK7FCPwq6KgFaeRhvyWAOcqKQo77yD1AhGrt83UQ3R
lxvBnkjsUQWY0QtuxzhnBNtecVAxCIYrM7wICUvgX4E33Ahs/0my0029FVmAVtVv
7ZwP4lRmK5RlLk90srqN481wIC8NLC3o2Oq2lmIkDYfaMIhg9eq1Y1wSAtPhJwPM
Pol+4OgFhKC/lySgjiRP1elOuO7xFs48VvhXF9ehya6fHVmkWM4NPqBvSWUe6+g8
w3i3uvhe++XFN377IRS0nVeRdYraFdkz0tKePY7495O8botZv2bip7rT+iMe8LyO
Uo46/MicA40+ZgjqYqChyc1dZskzLZbU1fgX21OfmVA4csw/2gk5z9LAEjUKhAVW
IduE4j9tLUTxnV2ZD1ListjgpGpZq+GP3SRQMvsneYX+YMCmjE/RHt8fNjKBXvd5
UsYZGCZqM9mL8lSBRzOdGvpFRvo785c309axm7hnoQchR9s4Z8YR6HnNeekf/zCD
N3nFvJehJbtvA+59PBLBdo0EB12ZTn1uSgQlZ1A0N3xL5cWZ8Nvhrv/vFiB+hDzG
2RDrbrN+wm0hBbgYKjetHsh36Ige/07fL4+Cuf3AfuaiNvujGM1E9/oE/gA5WP3d
fkFXK5MZyqWO3F8UffRZM+OgEOkAUkQ+W3VerINO8Q0dq3hQ6Lw8e+8JnoDrJapW
WzWVHttRMwv0ufo/XKQzgk8XNN2fAkS12b2oF6gCHSLP4P+9JZaUdEhnOe6tkOKD
mjc7+7bHPXh6q47sL7GLBsEAgNZkKiEWqI76smbWoid+GTKe075dM72p8bhW2Qi9
1MBVD75wVyrPifFQ3LPeHxJns2jyOjSFy8q63lID6NOS62y+3mNTuXgsmFzmb337
9hHd96tNXFrOyrdHaqLirY99dru7lplRLZbPLWXjrPW0Xr8J6wyEXUfaRoVHh2/M
mqfO9Krw31p4D23oLdwMxk0Ge88u5uJPoLvgW0fyWI2+Xa6aV8N/yXHaCPJJNYXL
uWNzDrEgBznWEPtBcrpLp89pBpsJpLNTgAJfKNoSoa4nQjij90s3qhfxNp7QKr82
Lw/2jpzwOOdgB6Dn0/xukLaKIO54RA9tLpQME+IoHsCDumg3/Q788jcqpj+tGvlu
X8w7k+vElahcLOHHVmSe99KE1+cjIYRDgOIjx2w1K9mvciGafSqLRTt0ASQnUeKM
FquiLn0takj9R5M/FrDVpbEX8aCPtIda736as8mDbaf2QK0YszWnwK6Ydim0Aiws
6l/9dUKwmOb5KJ8lj0g1rS/Q9dnTmD3ovTMDMepiMR4xoRl0NhpGx1K+0+1sPFSh
cM9DbKUV0VKQD6DusBxw7gHQBGzg/e9P8Ib/JObLr6dX1KXhvizd2y29TGQpFv5Z
29rIHXpVEC7mwMxLpSXK3KqmBhFiK5s/f2qReirx6eWcrbT6vrRvCFPfg7NKWeHo
umGoU5rbg869diYOTfa5n8aAaod2Ij8qQcUb7gLa+KwOpIBVjO9XMiZFCWLPrF8+
Zb5lwWPeestn2+crkiywLBUC9W6qYncv6gOZdpAXlVqF5toegL8m6LBoyyUE/0n9
bNF3ACCGtVQR3RyO+K9vHqxlo1PYPXhhKadjM/jpAqpP6ACE5sfTuafg4BRUnkqw
N8VZ2klBlo1sFMM8H+D7kPAMUzMGUkyfpw8JSbjiVRKoBpGp/xj2NpHiGr/4YET2
nJEbjdAo/mcj8QLkz2rYANVD8Suq1IMVgd1XVffokv9TVBng5BY3qQ+wiFZRgOhI
rNdLMRsbyxUXFYncQ6Z8fV2VMQVVl/AQFsPjPiL8TfahSb7AkuHyy7IapTPL8Kw1
I8O746mWcWDrYxaGpbimI3jbSurp0z80G8ag46czIRz4s2t+q1Bx6SBfdodYp6SS
Pk+sLOShv3jbf0+ctcHbDXzgAOIONw9hBYZKI1J1u2ZGDQM/VD1rUPCkszcS2ner
Of7Gj62TonhcOLogkc2wtat+CbUtlUSgEX3N1fZHqiPt870tqn5WYsULosvt4mtT
CYyUk64sCPVzpHmLs0misDRjOl8rzc9v6THcPBxWPvlEkDbIRBJG+ym04XAMwmUE
b59tcd2MoTuT6T1pkbTHdbnKeHl5RmhLNxhAlQIok5wst8558rLNO0cXpijOPVsg
yd/SgQBniBOFzggaHam9/PreQcrZyY8dbJFHdg6yYlHLXJvlBWK2UOAKNDnKWlSq
yr+LRge+tGdT+m3rwrS61WT/dYx0NFs1P9zTB5vMpCF6JyOfVCLLWyW+8yClQn4f
YCH5OGsgr/xMSnVJm8bI5ZFOtudmICV31MX1ORqyR3abOtozc31g/9+ui0VOuD91
RjGtnK0bccNb03Gk1hh0mDt6z5VIh4yKFkaKXCEt8ZOWG01GlmoXUZ7Wo5uopR1F
L+UcZvw7mvwA2p44toidUe8KPajCjzql+8pRutT5QQeIluMIzyYfV7PwDO/vBRMN
aS2DZkKpCbua/jrxeBF9Dcn+3fmTLE3lAtz8fJNUNeYvdQSozc4zR4SZ++46unCA
GHtQzSQlHd0vxQ7Epw8WPSjadrEyeJu08GkBydiSZ8SKrLx6UAo/2QEcII+tBHas
9c8hE/nkCEWyM6i0cRSumLSFqjTeKRBWfoK8VZdMjojYpQbBRNbzVtzmJYphGIUO
IN50CBdTL+7akBNHAIoLEmalLVoerh2EE1OzyxlLT1w9rMYOeglJxrzOfU9h0XMv
nYXkD0bOm5+zkHSshymhalBilfERUK3tAmwsQnMofAujysKy+iMhyhCtJJJW4Ydz
uNtiG4g7Q7OSF2HsgmcTFqzhgIE0mW0EZ4SHKjLgh9RtUCAghpw1vuce7buyKyPJ
gkuBtnusYQLDig+69O2QzmirgXqH7s7Cs5+50xluLKM5IFO6qzx+ckMJWW/LqFu7
5hsQCf7GjLhKNxgT9w+vKeo/zGsJ+OcU+pYaquQ9UZTOEDL1n/NcQfAV/oZ/ZUnF
WzG+wlNku+dNkjFvoRKJPch/W1kUVlNEPJJyFY/cY/++46AUB/7ox/QCtGTZOCmT
SWHNSGBC3p7qxVAdmx6E8WaaVvjvBcnKe567JygiklJundhs3uR+DBSOcrLajt+x
vO+wXecF0l2TXZFjVZfkbB3KDuB3hMY+UNiNQ7va7zlitGnYJvVrHELHFrrt663p
dNk1wqxHL+lHJiDisB4drz5z5dxyNn9TMl+Upwmz9l2sWMj9agYLb2UG2yW/3gqc
MWzMrC+PUB3Fj2LrIh9Gptu0JZUEdx5MQCVGuAPrxwJRSyjvQSGie6IBTF0fNxc8
dktrgyRDes3uAi9zYaQgXhMeHydbOiJh+nEK4Ny3mvceJCPMnjAawTDG1wIRLCvx
sjtCtCwm3JNjDVPsjjuL+m2ZdBk0BgxKgM4EqHHcxA0UCVXgew76miJZYbGuDSKU
UGZlWSMoV3/ZBHuz8F8SYntzzAvD56r89ejMObchKkrXbZeYTkumF0pKj/nlKIzH
LU/wK61IM/gPD/b8OTOlWBxiQoAzXe1ri/WujNLqDPBPaYzXt8PDGmc5FZTZO4b0
7vEtfA3W5OlBhdiacdpB/j/XBBHRpuMIhJfRrYQaqq39pDH1lChfOuQ9Ky59HiQm
KY2cq9K2spLzG1RmrofSqdMV9TuaKEuhukb0DOWfsdZW2DcKNo/r/Fi9tojZC/B6
RUMYMH97mx7KxnDtPplXW/1axu6Pb0eBK4eY7LeBOL0UbTbL9DpCD4zUxuEfz7GY
0Opv3G4dT2Ah1YUvRhm+t1HjZ6K9XwZxkbW4CkHVOuuA8pFgyLVwjhvitAtpoXLK
mDWRM9CAQ5He4LvKm88HrsbTQvnAt940QTsfuW9Y2VnmNe4PWjBvOcyS8fj4abL9
Kub7zDpG/Y9AAQBD7MoJ5btCFTOZLCKPJ7m96Va31eB+GvDKDXXwWeskSFvnVJwf
0E/kZW3YT5pfjFeRMaqkVEKkDMWOtE7bO/kFzMj+ht6Tfu3aYp3nv7rfHPLIcvyG
RFVP60ZpV+cJs0Kb5aCPZdOVWyXKCNmhliCpIGP5yk85CnbQTB3zk2YgTmR+k43n
vpmt0X4ff0zgIw2F2nc4ztUyzMaxODquyHelDN6BT+x9uw1AMWysePKakOW6oLGJ
5vrgkz0V1JkbQHJwupLzFN2bFZQvqxpYqGLBA2U4zeXeFDELdBiX0Eyt779kki9W
64z7eO6UD/Yf40FxSEUpBS6AttZdEixIu/DwmL8W5olaGvTpDt5S2l44pl7ivNx/
aPmHZOF2C4mrf7HpAtGXbfB6IlbutziIpCSJ/zYiynpPprPljt3VdJNxxumeS2Lv
0sWWMg4/+vv1sI/I6VTyIuOBcqr7VXgKQGcvPX9W6VBPfIVMPm6QRkUMIqk3v2Pn
YNJQJ8d8CEvwKaxYjpK+CVu/N/Ti951N1hfxe1nt5QFvwgetnmqM6gLjOV/GIbhT
cMqMbzIn2buMN3iptd+7vic+rFajCdKD5Sz9/bzrtFHzOJt9c8vGqib5UNhSSNfh
qNWw7ziunCKuT5bbVxmYjT8mUttnWMhi+hM1UNayi9vyHmogpJpClv7Wg61i8nLX
c2UYt4tXCF3WwfLL9kWX/8NXxt8qzLkBbDyE+O4xLn7mlHdB3pckRsjFZPRken0c
cZoD3xqAn8dOWQR9jhiBN9FNVPFJo/kEXwHR7ecwQrRa0A6YbMeMNX/GfARydcyd
LCeg4L+oaLRwZ8GSXY6ohXCcWSOzORjQb5WL1oqCpQyKUNMdSLnUnLNOQHPuCWfD
MHEV86AVHgiyJpNBS5a2AFu9CagxGpNka5PtWeBIARAA7OThGkO2U+1TuxrIPrHf
utX6L1sXov10iX4bZjpWeQJv01McVC+gmRA4DRlwsDQnduUU0Y7KIB8mfp+784uW
U3MUXOBIZ78FUs0ea+jdYU5Coby6udW69Y4+F8UUgv74zOqIFjbPH9FR7/QoIiYh
N4zEcLJfI+AZNSato7UORNcDDbHrDGxcIZKRZNrsnavudYf4ns9BlEKIcW+kL3+f
IKGmg+PPKxtrA4sVGMCn9W7lpThbB2wgDghby5GHxjVjds5LrsSk9IYsWeIMKG6m
q3Oa3zpcakCKtnsel3S6yGaCdnIYKxFs0+w/yxlk4TnI9zEtpvj/DzzQmrOKA8/V
oJ0cuaP+7Wd0+6Vajm7N8X/8hZz4ujcvdKaHBEk6867TyOsyq5+IRAa/MArizLgg
4OSZOhHdSDlaI+Y+4PWfahJJcKeTjTDhgA+LkWB6bkdfXd/wmQVmJMT7ii/W8UAK
X1q6a7UetwWS9E4F/RQwb1VF1gHxbi+/2q8xtR7yBBcXVGEzvx6XNWqufmcsTkz0
fvfvZD4SURSTdKF6stDIcyRUUGZ+OveL4mQtX/l0RW7DZ4tHp9lrnh16bwmJWlDD
4S65QQFu8kuNG2X5HGCNaUHXeKbxXKRd7+TmGNq8jnLYBE6QdouKZ3QN6u59ERzW
Xt3h57Frjlx+uR5xf/UvhHRX/iDAdcev0ilOmIZLGDfQWXYk9xnQkAED4qVa1E4T
6N/PaUJslJ99rMbKqC8DHs6o+S2HhOe6Dh4kOtg4RVoWtu+jvIQH3uKU/ATIuYBX
GNP4dsK+y6o4S7K7MA8+XhmKmKXP86pFukMjbOt/EMULe6haQMWRnMMM4dkqqXD1
1OZhGZW1+unY4TV5gecjtYdAeDPbvHKjGgCcadW/D2WMR/y+H9Qo6vrShKlsZT7/
zIIwWXqlY1/DVmW1kR4IXgbvs4e09pB6dab0Wo81InE0LvLjHuCIgxBTIUCTZjCA
OBA00nTLjVGaIpb9nRviCrZmK4BbMdj+fy+TwtjKX9cIcjKvG+RNzSZtgNr1oZvv
TXUhqitx/+PqxQ/3kvCaRysfO/Fk2COIi7fwun4vCK4F6sqOPUdJ8EoB9oqWhph2
GK6W//s7CBThLaURvrooUTeC0Xfh5yz/KoItxKMNItMqRj1uGOk2e+rS+b4cv+/w
ng7SImS0oGD12uan5hcxua572Z4xcHbZZzm8yfjKF3q+LojX4xb/5BKbw/uIOE8h
a9nlX6Q+rTxM8JC93c7WtU//hnv4zB7Qg2UOqqByTglmFqREF+a/gnFGcI4oVJ5b
q44AJSCnEwOa7HtOeJhME0FEnOw37M4iGvQxL/7EKn23TezKjYHUEhBnu/dW7kC7
sOknfTB3ilGcgcr3G+wBgRFj22y6xPw7h5AzrDnw6MA+VhmsK6AzrkTDoA9r58jb
8Fy0J55++J9c+FKeZ64PUjX7/SudfVpGULRWaZE4EJi6SpTzk7Bvt2DSaDGb+EnN
Qkpn1gSNRJ/FhG/vBAHfRyW0bEwz+IU6fhz1weds3GXcq7jAyzxHyRxZQiB7mASz
9mxwc0fM8VXZFZmfcClAUw0ErhBsM1YxcfNsQsp43+9ZZPSHtizvrOPbHDVgtcb+
eCCvxoRYqLr7le2LnAIH4fePXb6F8ZbUBwBOPNNW8I2W2gV8yo+UbKxQ1pESrHyS
ADwr8pIjE8mrVi7t3ZljX3iWU6Q+CGPF68tSWrEw/ynjzamHDo/7k7AawOv94hBq
gCi5CNYawDKImh9om2GyxCfVCipEMG/+ojJgo7RM77YrHKDz1nm6va1YRZLERlCe
8SCsFohFSs7m3UWbZyyEH/MJslbHY5nlNCKM7rBIlxuJGM1343uQUmTiS07mErIf
B0XDayq0VmdsbP8bXpX6OXPp+AlJnbw0pOk/LDF6D+TJt81ykBEI81+xAFnyHE8n
iojy1ymeXtFJgTRS76p4WVT+hqUngKOFcWoxxD5KQgRNm0Ypch6Pb8PGYgUdSI7W
MdL4diIeQUR+H3RXXkFPQA==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
IC3eDPs6wCkOH46wbgkDQHvqxzzK2fAHWySx0GdVmxw1cHY1U2/UuyYtMShwjieu
g6rF8MNEgdSRV/SbbZ6dKryTIDfsLbN+nXN591lLvnQPX4ChCajZnJ9GmYBFmZdX
AJFmPHYvnatCbMYL2oEYvdEgQNb9k7rCIcmGAOYSzl1Ek8pDVCQuD18dCqaAOdq4
bnszhT1qgwzH959qXfCPHSqKCsv5LWtPb9LaXu+n+tTL0jyqPvqyORCZ4e8APJre
rMz4Hfe+IV+JF+Rn4uRctYWYsK8sN7uibNPaaVkY18xl4lRdK0LF+A5lmIAuBcGz
Iu3CCJv3j8fhvjRhBa1Tng==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3872 )
`pragma protect data_block
Kt3n/OMuIzC39OgRj2QdwVeqOY/zjvTBojbC8TEG7LueJlA6B63KWbNoRIlTAWHp
shLFPtVo0v4TEf88uRxFI7HHyEFhlVh0em359rHG20pPcKTrk04e5MeOdAixv/7y
ueO+kyabAOBPdbCdmvvT/YySMVYxIum3as8ERyiU7NuveCH3KjiLUzQOFHs3PfLe
fRT9SGF5LlaVVjW45WX7w/AwKsJjSsrZ0gcQq8oMKSU1IWTMVO7s8qZCzjYHv84g
QpSPR/xa4EP08waYcCf23SlgVAYXiOudI96e9RIYmO6Q8yo6JIkRTHPTTKivk74S
poNli+z5hPKnIfQxELcV21BlBmxPZFwes8kRcHmJEk9324biGcyCGpycD60+WkS3
VxwfWyAWrk4+avbPByxLO2gZZbQqpQISxAgFiLisF+5oDH1OlpfWeU1lHLVOdw6R
Sf7aBbV8oJcmeIglzq9mP4tke5+E2BLM5dTDMuDvD3qjnFCJCD9IV6br4Io08jpB
2Q+95cpPAl4QRT3FxZ/rHiKYj+5cHpmWWZDBotQyWoo0AA1yloE0zQ4lmXquFbNU
okGaESjdh5BgF4VG3XXKsWnf7C5icUDsZTHc5L8lVWOcKBQ8NAZdJOr4mb0i1M9z
h/ExKiFLCJ849bhnSut5/e2pxT7i+RHF43nvOKNCcDaoVtxikH6kWP2tBcvwNcWF
SVAnIsZuLaFKoi8sAqA6Mgfsuk/jJ5v30DL0VK6dRW6WIshnn5rvxu1K13MJnoBX
a4FWKyz+fYL0LM5zQuLLLFMBuqnwANEnvQXzVGgu9rXE3fb9sxwiePRgqYfc/ZVP
IG4MXXp6FadzdLatFa95U+SVnCSmHp/6xZ/bsKBcs/WIqpDxtnaswnxDaliRZdYK
9CBmWtIQugMCHf8TYvcOXlZjr6kCYKVKkmvc7ESJggc3/hlIZyyszwMK0YO1Taum
mNcn92AoMWhF698L+/MNMKE/D+zbV7s6yTEtGW/o0hPvBHVqdbOTSICXyQ6eKsIv
HhpKzLpOvmmyJvemAOVPelJUNd023levXSErgn5nLB8GIshfh+JDtshAfzsrmb9T
pwdq/2cL2K32gQuyA3M1CxzRTycnvxHg6aOwQnVw3Kpyw9YIvX3gNbYeJFePddlZ
zenKgstjqkU0KDPRSvy8Dar23ZTnNSxJp9brkl8fGu+mo/XWyJPYUW4Ck98mUwAd
dXckLlK5PJ8rgS5/Ip5rSsnt4EEqvM3CFu/t5XVldAl4GaiTjPhJeiRf1AH1h0eo
9uIh1d+D4Cb804QwHlNzy8agi3pIW1Ug9KIMuWaqYoai2D66z3gOJgO6DqtqDet9
BfQqtJ/jpj4c93VbXwsjtnYjL/YRQHBhUpatK7/mwpNBwScvjvVJXLck3XaaknYU
0ZiQhzOasp1Z3SpoS/qjF6Ue1XAOeBjPpAY/SneG/3P6l0EYuSzL4LvQJeFy9QrE
tMymfdlFrOKk8dDeqZGdSSHHYpddY8duMu8mhdIHIBrBUnLUcAZHu5E9I57YJekr
HIrYpmwLmsiYJI3+yi8b/bU4lxlPfjsp/4hmNX39dd1jyPio4CUEdY5hjWtKFXIy
8b5JxccSDaBrh8R6jDGZe9bntwgPUmrpLVRQIUl6ymiKgLcnxzovlCYhmpbqJGeN
1QUVNkneP/SNGGPGRdKhi8z5HR3mstFyC+f0GQM/9ytnBpunOdY9aRVlif93UzE9
H525JVMRvZXUdHSEqlmWXv/VR/oADqkJMwYI9ZbYYP/p4hfYxav4zc/3/5dMl66u
eywpWj47l3wgYPkKWhvpIwsdvvnjtSiZF1H9yXY8y0QVJRSaw1nl5hgumEDrA44Z
Pv81ibHZokgs/1nNG3umyx4Du+IMxCWf8uDz93snw8tznEP8BZDS5d/5fnmKAXB8
BXzDFqRo7Xcl4BvJ54KykXW3w52SEYrlHmPKegq/x8xCIhATsTltX6zIrdDUlr+I
5/0sTWJkjU4RFf76mdio67GkRoa0/kUw/DoX38SMYk6LoWkvKYj6dCI3QDwiFMh3
vHfl2AjYlw3syv6WT48YlhWgosLXDap1tSsbU0LLdJhXY7ALZuubbpnVDrgH/75e
RMMOh13WWYJm6BVPDR37aPdsrapzUKsSj2xeflh8UXrRCojWS/vYnuqW2E+d4Rm7
eV2Et8eKX9QiMacbS6/k30DhzN2FiqiZ5EwvnJ9N4wh8IBH+9DmhTJ27+2u+TJou
AkKN9/BFhIB9RnFr9eNw2h2kt9EpXKqNcWGK7hmHFT2XQPX7YSIxtJLTVF3lo197
SkFXzAIbZlrocnh98easdShr5Wpk3LUtzXRlW4CPkV91INtvs9HcirzcBC7wYSrk
NLXFeBUMGBNp5HEVU4CqtS/a5rStbeejXyoLn22rDo4S3756MVsPCIkEQnz8Z2p7
v7RwkBa1GXMMnhpQn91Qvhz7yvhMDvLLWgksC7cNPl/Ne7KxeI4G1o10W211wEL7
xSvSWpjQiazyyQGCu0JLi+Z7thNPxwXl7Ds7L7095cff9/MIDGGVBcwrcGBV7D8X
NGhsninH4sW+KZJTPyGPJhJ8rkjbGH0WqXeoxw1EnRACvdy4glGegaH5VaEcD/+/
gIhjMF3ebxnCCYxV0mU4elZU+9SFZGS3WUItuj9ic6qdqBzY+Fc0l37y8XuNF+t2
misTRX9ve1nw9XRLFqDqwIeinZp/ggrNI/3UIDlX7k7nRY7g/KWoIlDbkWHIo8pb
l8RdWBSp0gIs7Gkjm4ZHyE1zx7PlkfcRIhqouf0y0y00KgUXL6L/yO8wS755iEWo
giyEp+w8ZGklkLKcYnlz+KiAclVImhZ6rZ7MAmTfXBsgxqvHI/TBDfCA2EJHD/hW
VxsqfoF6dLB+mMymwUhX7GJrVWaufs3cYUA8s9BT4S6PKgIkG9sVknD3/gorDdxZ
R9ScI6799JTDl5xWUM6zasct9cuU6w2LbnheA1aI5kKmfghCbH3t6jiONwBzNmLp
feeEXVy9s9UKlj9XGxnrGQeTLqC4kFTiC+zqj0ccJpd1uTCR8PR9l671OtBIUpWE
dSfoY+qFuUV5SLJmYNsl/fGXa6OeWVW26bvM9HhTjuiWmu1b9Asp1REWb2NgQM1E
NICHRZ9Os/fLetfwFOymUY2e+KZrUBNU0NmvL245qQH97gXx1aEO0NAz+8nTW0Ot
4dnuAaGoc4pSuoGG03UzZLNTqZPKJuu7KSIMU7N6OdYIj8P26asidFR+aGF5CfVM
tSjxFqrl9B3a0YJdm3a0NxzfPHeA5WBXnIOjzkcKAJCd8kF5NcZAdapGTOxTGxhS
rYNLfDBHWr2fx9/xCtvM8YBRrzdLoTEUScVtyy4yQEVmMFQ6sSi05JLPy04MLi+D
GvK25ig6xXdxvE7IlvxDkkwCHLvx/9mKzirOKkrJkjarYUxVMIZapFOcdRrY8AX2
p7/UY2A2oIrZ/gej9QWb73GnKOsDv2SXrkNHxfHIPSacdgJ89ci9H6PbIAZGehoP
AvDkcWUybdHGs3XC1ptRHDQ5yRNRvUIn3B31Bd0m2ProThgMbtJt8th0dWrxYrmP
gLJI1yT6EFqNtzqOQ2RHD77isdGHIlmZtKyvJjAz7c0fHW7GgbrVjSdmJToyH/kL
HLVWz0f9CSPKQ4Vfm5gSaGvZiMIPCdz4NjHzFYAPWnKju2tneb3oy2zIrkZXCJhH
sOdpEP3bwLQ7Sj6KTzw8UJy8rdHXCpJ9gbURA/tLZ5eKtdjlzJEWp2HXYb4Dw+Cg
1u2K79dR2ow3mJRp9VpKP0G4mwCuHg8ej3qet9etlCgXf2OBlaIPo4w2Rp/YSO3o
0ufJniW8EZKYbfcdt5x/GbgegDtVEcdpk4KvM5eVVKHAYCrLY4uG0zUWnZQb3pcF
laYObDwl0tHQgAh/ACuhEiVcWlHRcPkvZZgpCBQKeXsaBP1PpWTyxG9t27ZoAVSV
PMVdmY8Ceah63kZDvvXFIxdtU+7pJUsOQJlKmgUOnVAoSn252Wskskt/cFYuN9lh
0Q205bfotk9wKht8LyyKKktCBryaxg/+1Y9v9DPYL29ELPcSF2FkGeud5za2djYT
uO3zfgFsDFSiBe5qpJCIX2bSqvhHtYrXfepcpPE1TPJfgk6rcJF1KbEl7yS6O747
TuDQ0KOO9b0DbQxKmLxRJz05FX/u1ho9jkPy9Ht+tbndCte4a4FrGj2kfcndslIk
sHOoWUue4qZ9FMxki9/zb/1wHsybc1/snyY8WNIVAuKn0Ub0zF4z9poB6/n6qmUM
hyJ2z9QwQJmcNIZvHxnJrsmjd/UT90yWcOI9XKmK+7EH+E56q4UJg6CX4oU4pvi0
dUS0SY+52LVoR1g+j2zqUjiazabU5xLvReZ6VBPQRl3NWsLKLk11zCUF9WiiP8/7
i6EUZa2qsFza8qt0BH/6bydyJCWCyE73Yi1rnLD2vGLH+2hqT3LJ2oK61+Q9I+79
hWet/a9WXZzTYtA0JW0KAHaznLCJY8qQB6H16FqhaA8YyEFDpXpAMSYGjoc5qkk7
aqtqo0uQ0jGq2F50VQJrpsFi5IIdwwxXldQ70o2uJsWFVLVOwf4TtWfysjccbECH
UEYmVMm7rsvdTpt6dI4lGFM6YhNuFV628O36fchAGoaDHPifZLky2cVJX+0pbKEQ
fcNqknCUtfZ90er3b1VdjT+2GiGdnZC/BOV1kuF5tfO5SaSgvJCodwxw0WCT9t82
Ojm1znqKG+jCF4df4uQyRZZB85jMabZwemcj8U4QX1R+yG57YdkBtCWi2JBZQmT7
xsQzjD4ZinrdUMZYd2UdMKG1GryOLCk+FefNlmG1sK4i85O2ZIKGIFe36+kQww0r
VPdE5k5VihPTwjC9gJZ5k8Rv4WGycyq6aBM8/TpwV9jIFvjAM8gglMOK/j6CnqtA
7lIqQkOffqajs5GrYXzZyTTjBGSPcYclz2WVFvTxVnXghHT5OU0PfDTdWtBW6mYE
wLnD3qZ06dapobHrIdKfduKpRtS6+F8RoAsJg2eqppjGG4pMdYsOis9zgx7r+47O
tYbvuMvUkR6FcFiJ+UBYCFqGu+D7M/olzwU6PZCK9/k7u8YeEQvtjWiKqBI4/AWy
8752ACTLx9VG4DJUZCmpTLaVAj46p/qBVC20JasaAJE=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
dhhwYPZfcQqq/glSQ5SeTSjaOD04DrmBkX5CGiTPAPFRjzYYaiGHe70E2XwXkizg
/7NiDSxvjeg5M4Y6g+uYjjiHUDny7TtVikCF6tnkdYIHilZgqBQI6VW1aIwULnqC
mELmFSekaLHdAgPVi54YXOcxhW893eZSY6/OH58rHAC2g+kSUCgA99drzwDPlbEF
pV4PWNXPfodaoqTrm8VVHogo9gVv4mUBzffIoFk5WlBhPRGU4ujKUq77NIZyWOM0
c7SIu2x/orZzHaeWPlS3JCdnSwMYvPSsGP0/woTk0RptB44IvFMncshIlD2Bpa3m
YGmtmLBCPstXnbNTqGcOzQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8368 )
`pragma protect data_block
VxaDQGGPPgo5nD9V2XzOn9Ev0kV2B0C8RRouO4meQRHwZhLnP2KZeZ19xllVRgfC
42AeGkWd9I1yc6pbRbzWnsGnQ+UPlpd0AU+g0jwIC30LPshtfdqWEFfEYD2zofyS
B4Oq897rpXnefZrOWWluDAutLmxQ8EJrs7Ncd8zO1YBFypLtCQ6TGhUbXJrcxMl3
Wn8k5SgYCdbuUHv9lA9M5APET9AWNdgA2bsERpI6F06Ofb+g96EZyGArwLcBAwmU
cV2uvLZQof5xDRuWewdbGalluDMSyRZLk748wukJuqTlVIljMM5Pe0yOY06blFxp
vePsyM3I0Ao6Nrj+uiZ/YkmVS+SEVTH55FwwnfOqV2IoQZgkP0iaoTz89NokIo3G
sykpJWmfk6ubx8gZrpZ+yW1V57Gv+WsFi4duJSdZzveZgp2gygJNYnqv4GBOW4Ge
psNtHZHv6xkwpeS7vmQ33CkfBvivSadAu9ESf50pNtp1SLI0SzSf9MUMCFfbac6J
1C6fz4Q9ovLT2bZfsXS1UsFJbq4sVWnEIM+BUd9aqTKmK9f5KtTC70PxqpILYwIi
8whuQqb9ivlhjHYCxLyRF8ZRQbSzgstFGYCMdwxOOCYZCL7Fdicrqh3UGd+3DX1T
5i8gn10SlXHXH4nonr9oFW7yd3dZ5ZEZY0NGdsDPjG0pEDcmFRok4cSbj8xpxoZg
pVYvYOrEhxDLHv+5QFo4teY3ySqgc4YtHJBM1aG3+nd6/tgWu0LR3Y/yPYpUgVbN
MJXpDp2hJmHE5rFgdvnNEKhj53l8gqc0SuDGfVXQBKPOBzp+qM2OI9+BuAyj1VAV
ftUzOB2x7jrYvFOCqlJUyJX+eJfmx+YCT/jpbmk6PP1UhnUglFWyYeEnel4mW5dm
E09RWinU+zguDSy9E40ad5SB9JVcP0d5mGIYsrJejCN7ZjxSHMTVEc2gXVOiYoXd
OHi84hCTpu3XEVxy1mvdaNSJDrVcY3BpbLSaGjvpATJM8O+teG4hDoYHm+sMlhzF
Sb5cmTZZXbQs8krq46Of8yDbHvExd2si8uH8W4ZcxiTqwSwN0Mn0P/V8fh/J62Os
NLMSgZTyUy03EZp+piIm++Lkd2vWV1EWsEP3pS3+Dddq98NmsCVeqetZQom+Fpqy
KPOwMB8AmVUjLzGmvGQH4CHTKM43hDdjgPBtxeCoi+P1CglikDU3uni2vCmfTEND
rgxAiSq+DKsci8V8qSlxSDXQZVTZppj2WFMzHUkUPA/dZi8kRXJdxnsDUoNlkhis
+WFHAHUlLLnS8QVnB4MnviYNRu4X4Qa/hG3vI/4uD6LKXkRpy2mFrU1Ya8YYgGZ0
Eep/cmtNvLT509Qfp5vxgnNZeqMZ/5hrBFlOz4OYtfy4w1+LxhjghtYI6vkw7U1y
kY8rtqgEfMhjEUkaC3xCiRp4ZVmOCz4+QJtNk9zmJH6D5vZvNAV7cY802Ag5K0LD
YkJdNystV1B6UStRnEglqBPoG5Jmr6nLNHnzO2hKOW1a1QSSXjVuCpC0TMlex9AI
aBHAmOZgyx/cH2v/WAMlMcZCzUk7Crp6phUbZxDI3tXfsCWTY+OVzDB+TxWKzt5D
LcbUOS2Z1aXozgxAp5p/rmb2OK7E5L1sDUNLsP+TEW+BfQSIMPMnCM5xmttQN+1E
kZeEjS2sJNN4NZIfecv2wOLOK6Z7SIMHxnX832P39pKmWlP6CXvq0QyF2dG0cofa
MpckPyrHrFckF5dSmCxNHQF14/VrJJrfy/gTLIUEM27oA6o3gHXDsTIxIg+f5U6W
2N5KXd85u7Tbigu0wy6q/geOP7O3VR5QaWNTSRU6QiJwWBlfhzDSODwrivC9tjNd
YKKnJTM3LWKhHSNFnHvvBewDfTsyqJ2xa6E0Psp6RBOgtyC46et1uCU12lIlkwIq
S3e2C90tBpmcgKd7sYqoEPm/+59Afw9JOd0Vkb59nhW82IIJI7mnPBv6OgEFWz/U
1xtw+S83+5GgMmRFOSX1vDBlrL4nJg05HniNjgPsdvuRYnNlfASgY0C+6q9LdRJk
dEiPKue+hApq4Wp6tgWG+vMiquhf+w4sJTxSZ8wi78W1/zrxDKfj56+T0/VqpHQD
/7f1Vm4p4oVoymefIfBjYK+mv5C1ePGv0NRsF4lfrERKHrYjn0reexbFOxczpso6
ZKxhTkv7xFbwV0Or7YPrY8tKi/PFZ+4p1QNaFoxBLqBPFJYnY0RAsgJ8AlAeajcL
RAJrTJx6STBxKd1Gw2RfSYqO23DBDexK+fraNGmMjdUHShTcj0p2gCc85N5maUbZ
BhmJ7ieIhCciJ1NNlKaFKQCidILShzg2cn/3rGTqbuktiSDWsiJSj6+JsbhfGqOz
Dv6dwptJnfeQ9i0PUSdkVX/pYHYHta0UMwFgCGmsIm2HmgHs++MOC2VKYCXlX/vZ
VU++pa/WYWKD5VGcTcYG6MeoLC71A9GKUezHYXYGt062XCJMC+fLg+LOgOlNo2Bo
2gCC2EnmPgghIJxnguJ1DKfacY+Y1TjZva2cL0vFeZwgHoTWGUMz+3LjKm5NOsff
cwQWjxSWqf++BqoVbBBjX1hevwf/bBz/x/VinPLtq5SC7k4YJHNVmsIR54F//npv
ixtceDBKiGdwmXGWTaD4+g9ODV65Ub3Jyfx+aRFur+ywnT24cvm7st9IcqIimcV0
/iuNbxZfmcfXb8qQRkUQ4DTgCxpTCXJ+U5iXt3JrsnlXymtrB62kjo5+Vtoo6xA9
bxc1W8V9BonkOOwjhxfOx02WUM8mHYEX/RKOCF57FDMykJwE8/ODgl7WGZyanZ3+
jaZOuELoMg/QoTBXBvi2LtSeCBBUm7d7qIP+9sky6ZS1fyv2fR4/SRd+o3hy8ZpI
6MTtRjLKQF8C3ScL581Bboc0Kvb1APpgdGzh3lL1xp9YMrHArSJigt7RCR+THzux
XFFAxOMOh3dktcrIkbXYgceVJH1f7uRu6LUfZIlqXjUJPB5Of2XJDJCXc8md7bx6
GIbDCGxiW3OT654ql2XJxIB83Bv13fkeYvPaKEgtzDfIuHmidIBbzQUYPVkuHKXY
wuojnpHjaa7lJUp0o4tCB2c4BG6ChQ8NhsC8IRCIQBv5/dgk9eNYEMr1SXrZYMih
PM/wkkRLmp/AZaP+mWrea06xnfEUYWK4Myu823EIfOtbiJEdt53I3IgxAMDnYl3i
xVBkll42q/mGcy5X/z9RFy3cohxEqr5naP8Zp+3czdnLdKaF4zPm8YMBoewVorU/
irsdYYJyJaf/YLKnjhwAz1CMg/A5Lkjt7fhPR7cdVcDM/QPRJlwt00WIJnltHWGC
rirbwgLuXEEPYNGGhTOalVhZbmc7IieVTEBZHvGHE2KVeChqtTSTsq41bx38VUM4
fjfq9fqBD6sSYPr+yXwyd8yO3zDEEkDrssVXcB7Pj5jf6mp8XH0H+PY6phYNTc4k
TSg8Ha+80r8aKfyicS6rcXQ8QjoJMLdCXrE+OAU+o4TXHdAoPfW6d0fDATIR/uZG
siMt1nFGkEa65WZ0sOkvc4Umul8PO1tI9uDhG9coGBkDnaSIcS4K5o7suPgnb1/3
Cng9nDVOr+GT2gdWmn/JRTHyR+PXKbeKrlmlVJWaYsmHLAKMVC0vYSVnStiSPc6k
vxy3Acza3/fnO58nRbqcIKKuGvzxKLAzqKbN1waozVhylfTgzoVFsU5O2s6ggWO2
/ZVB8L1cmgPd4rE2xq46nYS9wYj2FEEoy3UfcGtMxOZE6UkgkBNhSzeDZTVGSYCT
Spd5rL/KHWriPnUyNc7pm97JB1UI+eBqGW1wVOVPn+yqHVXXsGC/UaVomVp2dcib
N4QLOHXQtvCF2ikgk8b++yuxfhyIIJY66dLDjc/1TBmmQZsYFkwA1523vr9qAXgd
hks+EBkYgtu9KVWipx9H5WAtb3px6r1r4Fv0BVb3wXaOocMOcNwcrJzLlJKrnU2V
ghfESr/vcDvQceEtQJBkNMT2SjfEBhi2ARf4CiaBz+07NXy/CstGDjtCRNDtiOPi
MtisHhTaxvFWR613EildKSkT+DDYkbNj5E1ntRiDiTSl7x8YSuQftaNhYW/B2wo2
LuuBDewTTU2SDlJHCch+bsILZeaLC/Q+dnHFfJ1ZAAI980QbxDyKMgx7kIpqtafR
pq+sSrgtvWeWLt29JPXdHk61fWAsXKZWGdbF9aCo/EGx09lcwfphFk4ltjIck0Cs
DB7adg0HzAphwMJ5YvM020X6e4sC0ltsJcKBZ4xIMdmZeRDVYrOTrZhe81Ro9bL6
iY+ZIIXBN5///d2ir6KmhrshUDyZwLIBnRBszvBCJqnvyEsCE1eF4R05BqpPQLj8
Mi7fAD7cjISAmKL8ssd89SFa1iB6prHy3UPWwB0ofWWdnEQaGBEkeljz4+ksbmdP
aIukUMYFCp2IJKUqPXI9TqrzH7u1Pjos3994PjPxJY5zWk15cteywaJnjJYe1QTU
RO5TGFBu86e6AoZP5XqkF3tVGQ/Bgl7yIH+enFxPoVFcrW5582uyh8BTETsrgZro
Mv1BpDKPLIJ+WYnqzjQvf84SkuJuUcn9MRD9jInhz90bohjK4Ep9Jt1UrsENOxLc
KpTCgFDfuHY6FlFlzeUryHT2O7bGPJF8nVe/MTidnA7HgG9u+30W7+6ziG5SVLDp
/fyyXRsvNqvpgspiGpNm4WdkSmi/WkjiSqqBGnoON19ZdlSTEiETvaePKm9Pi67f
+s01JnmvHysE7ToSbIr2GIyCZ8IHED84uMYA+zr30J3nJeBXEJOJaN+JMvEsjgMz
m+sFho3kpJ8vTBJi/TfYksj9/AZuUR4XhJM/m9e0ZFWh2StgN7MOdL58VJigmg4m
/zLtKdNwUWPQWaJSRrAYLLnL/5HaahjNMdLG9tObkzSuWiP1q8WlpNt5IkYoiKkh
ZTC43iMpgCkCkBI0mo2qIFZHM0ELjY73duJCEDQe/keiz7LI+Izh3yJ8dItJGqCQ
XaeuxARZXSkBBuPOPuwBFgZgWr0+boG/Bsp3XcQswbzzQYRUK8Vbu5W9lbpMViJV
Zn1Qu7FWHShz3qlRLgb6HcWcFNlUzyaV7L4G5awYPrYHouODhUoQu9jcjU0dq+BW
TbxJ8LjzoPVzlV+o0VP6yi1W774FYG3Sf+LMaVWqphq23/7iZPUKVed73A/Y7+Z8
uU48W32S9LPH+IRZ/Gd1gcMSq4eWU4QcaY6FsxTCbSXciAIUOPZcSmmrKXIyzaDb
i36zOJAM6GY9vdKaT4e+4okNrwx6QTPVYm/JbH6is+5Bs9O0izmRuQfMjqxYL3I/
WYk/8L+xLPkLQywPs1JIb+d4Mwq7nj3GBQ5Dd+KunWvvVqnqjgs0sfLz2Km4g2ho
OaMFXrkToQLyrgD8euVsYi3alYB0VVNpuQrcB6Mi8/cL8ucbYl2yXceAyh2M9cGo
JsSEyIuzG3+0M0RqF/Ny9NkFzFUkL8IREKg0ihvHd9K1D4UMkVgAJnTj3wRPkd4V
uMgrfZRGvJ3/IOMgt+18glWBqvs7za+7WAvm5UcUSQqUwEkw3DMcSQUrN5nUO5Oo
/HYDT0qeqPUT6ylZ6Rj14hQvPN+ECVjLM0rNO1frTPX7ls/eNFc4L2lQOD53oIVj
s2fdsvOI9Y4EbUyjM7WY89VPK5iVVjyHS2Zlj7FbNAOOClgY8TzntIyWMhxfSP+D
4UoN5oFGnChF/yx7LADCjE36ymdVjbvlFCtbCjE2yqnS89vURbj+DWZWcc03AR+r
wqzoqLCl43UDbGj1XHgWNv4NYA3l82YfiQXJT23DDfIASBHsHVZUUc5GEKEded+4
o8+3c6joLLMsnH5S/fkXrrdt+dP96V8puIiPSUwi/hYyuL8Lmdx95m9z3FLIGc5T
/4dzDKH09gAjBAk8WreKKHKsBW5W5GoihAeLMX0M3tbW8py348gUyHPFw/wPx95d
iUDOAXh28Vc23D79vOILKdJJOuRZQyEB6CRjYr+m0mzqype7h77JC65dCO7Q7VIn
xL8/L99ndsz5vN3rf0Ixk6WXTssu1Z+zkQKJqq1MigtzrLdttznuuOpJsAwXSbux
6VhQYgXkWZ3ckVNA/eikNjJNvdF+JfYhexSYIBP7XFSwnH688FLqkT92jOZWyE21
GVrvk9bG8yZpgZzpf/0JUaL78FjQl/PVFeVQpyyxI8N/3ryjrnkjKJYZCS/fKO2k
Rnl2+r5p/+lPRlud1JIEc0jHHWiFs88I92Co323eIMbrUCgHehID3jcQsMLELSdS
3r4C/xHcie3bLV4UMK7+FdpIuSACFcapJg3ywPQyP7ZHCdbRneCUD2gPUutVjHZG
kcrlZE1PauMIIoVnzktpcGzgIshHKPdZ1L4jSnkdk2LJf5QFJtb8JyqV/M0SDCCC
XPzmvRM/RUcxMFw+fxitcBOn9zmMW6+6JfNf84oH8vfPfAeUA+flNGyw5Efe49fU
8WVHCl4GPvVofCxKOaNjUUbioee8MrIVLe0ZoU0cfRsCCk/Vvf/N8ynJ0k5gwi6s
GJVryWTr4qchAD2cYwE6yMYP/AYfYlGBXw2+Bq5TDuceytQ41lALQgwff24j2hm4
8Up5p75khyLF+YtNGSH6J9Iw3/7F+iK/2hqGWxP/9cyvm/Q9WVsiR25jCYniVr5b
V5NQpb/kERp9OdR00T2E1Hk8YtrRN8MhjplosrFyc89RJ8t6Dh2CZ1CXBtTbPMph
rn0VaCOOT7sWyZn6PtaogRkPLMVFSbhiXij4Kx4MrE81kQ3JvOioGvw0MhymyR6B
WLT24auDQ498sJixmGK5cmXuQqml5pqSRrfT/DtSAw5rTKOe81kTds7+oXozShZf
E3ESuGkYfUjDN7X2QI6ZnvWBuOipb8f0Sccg68uqoZ3Fy4Vuq9DbKDCfQv/zrQ0L
wZJrIfi8YGI0r002uL43ewPDUOq6xz2khRAESsa8EXYL8c1JS4mjx8+JNp7esrW4
2G1JyjZHXWCH0ua7A2FO8JX5UbOq3gLeSmOmuhIXcSVZCBG7Ccjge/8KFH6MqvIC
mbPdbsFTFeSlBBUKRD5W7cz+okR1uaBcFc103CJHAjxgrz+wdRpbvA4L+tG9LHMH
K/mJl4Yr/OysaLebyGjYFosYCPQcb+Cv3BLjQ8gDk5FTCEKwOphHfH2cFMQYVVlS
4+tnrRH63tu3P9tEGfrADkCWYipJ0h0Fdg8kCkrh54tGFW+gnNWjqcqmcEPSKyAD
AFDJyTLeCIzgF5qkvg15pnkODltfaZs33Bn5N/gPSRo1RjAa8Y8VeBcb76JZWyKN
IdOgzqQzU7cEtKdrALict6m0L0hA3IHw3Lf0K4y0aAQ1TeNzAazhvjU0GRoNwFEq
ppVESzh2Wz7unDGCbAScAdUw38TMEP3ZJlWloo2Dg4c7o0hqMh53MWtAH+nSHzVR
TSd1hJe/TxS9LHCP60spoF6lOHpKdLi0JbGxvhW/OD4UGsZoSupwjaYcmPmA1Ugl
GBWuVazJzSskw67TaUBHg+l1jzHIsDfrPg2sQ05/e/2qnmvB7ttaayfCnyNysz/d
7K3OE14J9Jcn6DzWz3gxduOnWx6IejEU3OKEigNg2KDKxY7OVdZd2jG9YjxwZrMA
flRP+Oqf0eD8c0b18INf1U+SXLbUhlNwIkoUb0PeU2Z2Pw1yA+aU0j7g57Y0jEXo
fX6jiRo7LKAWyZMnObatyxSTqSWG4rLZAoVK58pCSyWkrxlfD93jVpjMOtFBHSCf
RvJdsk9pL2w0K/Jd2u1Z75Mse0ihMgmB5No/k9eWz4GMTxztNDaIJwAglir4rfyr
F3EsFHA/sIErTBc8aq4L6KM9BHGA+YhPnIpT4wXbPOikGESAGhYkg3612U97p1sb
Cfooq8wT+u9pBFarSNBZrWNtRfD/gf/w1cW2L/T8lhMXyz/5OKz3/Z8D/forepzR
3MZtVvBmqBiUj4r3POhryMYCY2MjQQVM/nf7lfwdUVkKMtzB7WiJnhw3XEIoBcSW
3fwQGFY03GDz+eH0K5kD0xbf5MagM4YBurTKL+lZlEp09kcktMFKFKkIYXng7/d9
0xv0MPbSw7aPIBlfDbpXbxcY+Qmk32eb0W92EydNeSMpjSbzzBj4OR0dws45LYXy
YLQSwbSQNc4zHX6pusdMKoRdmwVXNkWgGw1cTJ9utMfdAHTG9rQ72dPh9m4hd8cG
eS+Q1Jydz9mmkTNVFQpBhXsegvPPnYQ9OlYPC1AFunGXEkJ5sjyR4M6aMnIOD+79
ABx26sVCRVh7NjBgLaNaH6RhotG9ND3dnX6oKzyaJrQ90zUWQE5H0nZqM9wQSIQf
fAupjZp++XjCeV1HcFqIOhCKH04LUD//KJqlzLEvmUJBwEEVll50fZkX++ECBtc0
4oYKyhrFiOFaYzSWk/+nEnmO+FajPKl3GxW8sBJXNCubwIkt3C/5R3/10pPhMAYr
GEF8D0+0FEiFQjWCeiI2Q6Eg0MfIcP9NlRgb4xfgr+Ifh8yC4Z3MlSg48b4tAQGq
g0xQHTnPyW4EEpSads7434mMmxKFXajjH+Ky0UUtIOHOrGDtI5D9/hPAl+6q0ku3
ySQCQhzzv+SG0G2DmwR7iACfUf9P9QTxpHOZwNZ/GpJaGxnlgFNpwAyzTnicFtzN
+zgcBFxpTCIpezF7ZfKcvFfdEUCPl9E5mlzD0AFPhJpqkIfmYqwtSrvvydvUGwgw
5EQWuHVI4cOmHEmTyZ7p+oRISf+xL20i5G2WaL2dGzmtea5QM605PV8vCOraI+XN
G25sajhda3TFCkXyPKrGX3hAzFUmP699lTQjs+/VyTRp+jYGtLEtL08u7rP5nx9+
RSzLYZR242cnebEaeJl1WOtfQG4c9LkzCGXIWzZLE4wD+qGAmxT9GS02T8i0lBBk
F4k3wlzR3gEPgKW3nqVYa7xVWNr8FRX1y/v5QAl+JtfrZWZ1CGcQA+FmDIJ2gn7/
oIafvjTtyIuHv70x/tb36IahGRSkie/ddvN5xmdYPzvGb4ZzCK/MEVZ5RaBbzBgE
vP5tgMk/+EbmskuFLHhraRr4PRZhl1fK74RXgh+0/CRn3gYnpQAcPEuv0Zb6JxGr
C3IUkD0icJQy+FoC7vyZCVOmbDA3vYzSoUqKK1ZhVjCaccA5+YQPUoykvdaZZi9r
6hvbzPRTQKssqJvV74Z8BqZm8U84W+7Ietfthe49F/toE6osx/LFL6V/JpJT8Ov3
zmBkyOWndDYaDUJpBLSj2vaOL4/eBdEds2soorTcKnCleXsvicv21dQ1RAQZP/ax
s37dVzR77nkIoPH+84Hi5C/Q1nY854GRYYei1cp4R24N86IIoyT9a+u6PtxB4diW
rwLIy9w6Kb2HM5s6b0w8HbK6CbbQYMntRFg7jkfabmqOuHGtBB0v35tzPZOv/rQf
5g1Dcbl7wBpkET1EXw97Yk8Jhd/uqbF4n7mnSiVj5FzBdGqHBai29MN3C/lob+9q
evPuYX4DVkGuxGz0rTUqZDARkt6qWoruVOoa6CO+KRgcKd0IqlO+VLYtJiJdknk4
tF2GOkaAzckSdiX/rAwg3pa+gyFf3e253sZeyfgz/0JiDgvofHQzFq8FannZWj00
mv6MiJXvuVU/JzOYX8Q10ymoSURO5RBc8D7AfHbARwsIBqN6wEm13WmRKUsUqPSC
cKzoKGNruUncfdDbEccB2Emkivej75MfLF05s+G4ZTwAjr3H1hGNMI63pPHczegz
+fYfyzVAKdeZrrGU82Fsx8XOkjcm/jNQDLFESGh7Y3etegVW9JjrnvvykOciNm0M
77vaMPn8vjStaWVNP2lTkUet7ESqjnyMZ5/27zt3hZTzbN/+ppdigLSLIpIKH3rZ
Wf+ISFRZN/sup51VNdb58ZdPvjMB+6bSlOea4aarOS8YwtdRX0SdpuHe2NvLNjwf
wYQyWwOs//GJ5l85+xXCJHlnTCOtZs67e4MjoppxPNSZIlSb2zkwDmbNI34ETRef
EeibjJQ11WsHP1KAtjIAk/9NCjfohUDEG9G5Z1K2p4eqTX6exK9yeEzCd8RQzQMa
teHbZSW6vAjByJq5bD0XvpUIklxJvj9N+qxmkiX01+Z5W5wmatLHarWMUOTd4TnY
aDqLbeBxmkp4As1eRxD+DAMdEbGDVeJIPN6yzAUjnWGyq89R9OkTAKYR8vA/k+5+
kpE/sxJZjY6r3VkMlqLYhmyFcM5AVbqOnONIPCMnwplJSFOhZlkLK1oHLMZwyMGI
CmJn/IWLo1qASNlAj7D/xwtErS6Odzaaf94K3KP/ahzHVWegk0I9nQXYkHrAuwiF
NviSeYPhCi/VFTSYCGsHbURvBsVAobETOPXncHU5eyc1cirJ7eWxhWdaDujh1A0C
H2XYymyMZSyceeWrZ6PRur2Ko+ymuPOcYjhTIwz8GsuMMEcinneO0dbFDUvuR5QK
q/ZkyCs4lZIp5xr3IfLgmznYx3yF0xajW295r1nr+6OuN7sZeaEQVth9NyuTf5+r
8karHEgTO8K1i0CJcNlnHS9BQkDyfvEwtwD8Iucrk8aRUocxHFnq+dTjWPPiLBJ+
XptfuYeXjK/Tr5gJK7fEXnePmbjMrt9T/WOHgxzy/F+A069VVXHI7EQY48nhL22d
H+1jPHctInWfCV+0Gp1iS3ivb0IlR4zYlhjopka9y9rKiwRCcaKcH2BJN9IwwNLE
PRsXNApoNWIMpOSpFNuB+JGlX1N+J35ypopqBLz15teHMEjdcUnmUgEpqXUJ9UsM
AV3ByJ0b9Z/8a8tLo4AdXfDi7lgy1M6aPMCXHZEudIPF949efrVipN4EJuEcYLUo
l4r0gzZS6bmco3OT7zT9wXpDmzc/WQu8saREiqE55HFtCcxHb5ujMqE8p3NPaAzZ
VRAlTDS2be3NvkiK5/o5eq7E9C2QBEfsrHBcnACL+Hvfz5KMNFcjW7p8t/yidE/+
6pwW+wzBZS6bJfLVxnJ76NVcEWlN5d2n9FJcNrwSFLQPQ73UrlPiZqkSDoBJITD5
ENJB5wKeExVx3vC7RTNB/lfrCGa9TbX5H7VFy6vJRmfZQhS/td0a+VLhqHSTIG29
lffe0OyDXU2HBj14a63xIalOmh4Ia0r+vTolAJ4ZnECersa+pLUf2gBpGXueF5lj
szsuRat3qGiKKNJQ1ntvXA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
bsFpSXaiIuP3jAlI9JSePFLcF4WUlksKlILUfHbRNF4IDo/1acaQL9V7PZc6kshb
g8+jr2y4gQ0SNOASZB3CzbMAEg9037i9BLVClev6ESKk7nPeNtRa8aoHCKejsA0g
fH4d5dK6oAmQLmn4CO6CR78fqJor1PFJHCWk+E8ztZv4zi6SlrivG0WRI9/nsdbe
J30wFwa9EPBZrCUoWoqOIfCziyzibXBHFRESuowji9UXB0J+ZNZrLvSJ0ym2eQAw
pvfuBIApiPNUA2m7LRboHavSz3dC6jLKbV8h/Zr3/AHujgSiJiZUH9avAH33Sn6h
tYATtAOjudZl6SKkTvDIkg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 10640 )
`pragma protect data_block
r9wByL4xuVNOdE80Vv8kf8C2NHfZkcfNjjaZ42HcPVSXIs1MSFpXICqa7niqQfpy
LdyrnJCye2pxAzwJenXVoWRzpcDwrYIktklD/pfVfP+7KWPD1nqfYn2iXmqMe/KP
pbTMEFIMkvJq4hqgl+CRRpHLhG/e4ooHSfb9kNuV9y7z0JxUOVnMjNJREHiP3XrA
ppvaHbW3MH7I5FBcRhqmDXLe1lQ3b9HaUyW8sObsNHAxLw/y5ExmncBZP4OVGgsz
ssqxkaixwM2hm0sc/QRvlNgbGdWx9UY6/HKFafSOT0YLzacVU0qCf5rgLPgc5eTs
9ZU8cHmds7aYw3MAn1YWyFbOUW1Cfrp1lautPimpM0xqTyoBbBmyah3/BHMPZp4+
MZvIuT7DfwC1uJMxxE8VuSqJAUBq1Ajv8zuLlig3tVPQC2yWDxBS8wygwyH1xQOr
U7nu96lkCx/oe8FharBsX/y0JEDMLWb0NoCVs7pYkXMEZneGVrMzuTdMcUulhy7x
Ar+TmE+QPbBoLwm4XXEqDkxIKQdxgXvshAm7GdBpvma8Rl0Y6oF3CRiFmJJREL++
8ijFXf/9MxpDccryn+jvb0f6STZMQqg4FPDvS+bpT2Z1NCXXbYW9VQyDlnasmYpB
IgMGOYcC0DUn0EB+Bq3OIY+G7UpxF3YDXQDo1GYDfjCyblvqBXwrBH62ONgX7eYi
DbA/YaYR2eL8+0gHGJh8aJy8b+9Cf7oFJd4aYONgOqVh7axlTYpGPOp4papQ5/xH
WPGEFR7vL+9tx0oLFEEgDGJ906tCrdnN1rHs+VzzT3yIywLwJwAGgqm/YQy23jI9
Up85nMT4ugli966gjO9ye/j/D7yR73xCmd0ElVygO9m80XxpZxVqyXXvGRr5KzCK
PJoXHwa1KlN+acoRWy+YixNwb5HiJYooqzUPRbjl5l9nzlEy4yglg01GU2OkwhQu
+xtVWYbK49EpSrzncNbm5h4fVt2PDih3zGD4zprXR7p6mehokX3k+Gw4YguhLZZQ
QZ6Lm1p3XO/2Gs0cd2IP/Z0A0VWCqOdkGWlBDMgrxZGnFW8fYjhht8LkFcaTVdx6
kQ4/OOqYFitiZDEFRLbro1aJNvfzYsroOxNh1jbIDa0GH/ruLWDnNi/Sdeib7/yV
abBYHUWDQW1sQUSg1p8725WZ9X4+fXYnNNBx0y0IO3eDlul21s6IUi4lQkCDbLop
7khdA81nQ2JZwwuF5MVL9Pj6CmqEw34M+xj8wqrdfrtjMNndnd8evIxmOSP4inEK
Ueb60xP+nbluMFHbQN2zdbyArGYuccYXSGfK1NzC2EUkU9lJ09lk7BAux8QbMnHB
gyZRpQNXAqJTwTz5TxtrVlpOCo7E6cv5lwl7vUNGTqthPZAGNFAhCeKPpxIqoRsa
jSL8mvSvqTO6qrBRCZI7I08/nY7C7NTA4hmfi2QehxIWxTQgdC/Cb/E8gM1wboxr
R1uMaAblbqj9BDH3Gx2JDkkmNp8HBBqlTampjg3Nk9yM+RaX0JpB2y6InHAz9dvN
lFR73u4MeWyudnPdUMZuomlErW0JSEkhlARgwpeyNQaUd1oZBAjk5GT1anm6GUqz
PDR7TlX6dc9NyR9/FGR34T4nBpU8GjGmPvWvDtF+4QslGj1qS1E35qF95+A1VI7b
8biHAEwdfup7km0bge4MAkHLGkcA9zVkmH48tHPBFhJDKCN/CaRPTDj9iE+GJ6VA
8Dp5Z0x5Z9SPJoeKMgwqe/7zymz8RM6x1rDwguK+z7IR7u/fwU9c7mBAiNi/HJBC
DzcG49behyPodyE5hjbaKQRaQgydIPEMbmpE/X6zunPVBFGFYlijSVOQtGoHzBqP
kLtX1a8tBF1WB3fn/x/Td0sk0v70EYXrurZ2fntY9RuABY+i+IwhdKk7C/2e2kb5
4sYYUP4RuQ/W4PSeNZZleX48W9vWBi/xYjw9OxfsqCUarR7MH9Xs4qK0r/1Zi/7d
57gaCF7hDzdthuNP4RYu7XMmTF33PZ9RZbX8gw8CSPBCzrAPvyJii+hOnGL5vHvr
cuOFP5tPJ98I1IPdCFzj8e/JfrZQGL+6/DLMkMazVWX7envt1+bUx7KoUp+yFHdb
lWvfTs7E79XJJ/5LI1qN8XIfgScHkJTBICA0bXDSoyY387KYTDPkBo3cxbNvbp4w
ezVK+3VKfeSt4rGQ57SyVyQTvRdI4vnIhVbree/gUKLaSPNcI0tc2TCxNFLdfub7
VxWRpo131ndZKn8SBfW4B1/OLl7ghYbVBH6h3BgHw6Ccn5KqE+Eet/se6nsiSoW8
b5gYTXzJc+k+qX8F9DG3tNN71jZa9szFO0cy2k2lgS6dL642mxO1yPSVlSm8FOK7
4/+5bvTOJ+33gX0C9p9KWr7gt/tKBBEhAr5+jpcEPwCZDwG0Ek8dAIgNOmT3B01f
Gq2kK+MSO7OB5SGY/cdamhgDHuQvmiH3bCfEmvfLAAEm/eaXRBCefwjiBvg7TsNN
kqSub12PNroduPgGrCNP2OOnRnEDL+tPjabjT3lKGCN9WXn5Kt+ATJY1VbSsY8OF
CXCQHCj4XMQPag7tmY/uiCdg7p0qwn9vDvEWtIMjPiXan6/gS6eYlmkL6XSktViX
VbBQdbmNIC39xZfj4FVJzRh6tpg2H27g8rhMGasn8amj35y/PPVuaWdUr95fI3lM
S3qTIEpN9dFI5xNdB15gF76CeGm+WBhlG2S0mB+LaHMZkt4l/iXhqdSwqG2P19yW
3drMSDHVK9O9wbzPM6DT/2tnGBoE52N8RWZg8yE/GZr7/mlCd9W4IerxgYZmg1NX
qpuWXkUWIRUoU8Blnhye63wf/f7YHA8wVsz3DrB85Kf3YgI4aBMkU9Z6t6+/fib/
S8vKwLYQ0z9oMXqRH2i5J5qvDK7sokBOC/9BU98E/kJG26SSoTp2gqRLQtO3X8FZ
QD0+g7xnjJs1FicLr6XL6WakXD1VnyZ06OPTuPkW6tzAhUQjUCgA+6MFzXg5Sg47
hz5sWLxuz80o0Utc1WqqzZpY1hVcNeMj4h+3CBne+VUFfbuVzmHNBa9mmMgss8R4
8bZJ4xte/NhwZKpJPD0qwVQ7XMs/McUlZS3JfeFoYt3i4Z03hB89nF+WhSJw4iti
Ab7FBuOYd7TrVVHwUHOb5hiNxlf+C+EKr+2qyyUqB98kTz9b9CWVGkj4MU32pD5g
hSK1ka6wX4G1QA9W3/RwgfkL6+Easd+cfUf6TD80G+1N8WOBSwAxc4Edj2Xkvclt
JGFEZ+qh2SbJdfX6KR98/zG+k1hWx0wDsZTC02pM2/68BNNTCcG/I9E0SAJBCPmG
2GbYyKr7Op/VF7bFOc9g4dw9SA30fC0/Y2Urh2ToOL2RgJBKiTIkdpjbFcyhH87L
KkV8bFPij2oiqCGiX6d8vB9ZaNWIP2d4Q2LA3UkkfAfUkxACFkRjlzo0xotJZAhE
1C+DxKGLhcWZhujLLpmT/yfJLAvNqck38fU2aKLIM79PYuWAH0fIdX13AAUvqohW
Kye0GrHag5XbFSU47C2NpW3hS7AKEc63lqC/S2QkIQ7/NTliHZVLEExAaqoiqoKb
0PtBU3F0rbcARLQa+rV+mpdIWK7gh5+VYXhnYUivwAphZ4y7Vcte1r+L6DeetSfl
LrYdcAOSQRLFxtNW02lyyZmwZHc+0Btk2Wg9VKes/OsYp0ICTp/gewgrcSCMzXlk
6QgVkxk1Q/aaquR5slyxe0AX2BuRA7hdf4MXQHEh30jMk7gev37gliv7u6qL+oVe
BrQQqPHAStGPkBh8RnKQXHuEHm6tBAE4kiq53aU8csQcEmDOoha6YGcOkzEXSKjU
f9FkiZzumCUBBWN7dh6Bncgj5BrbEQ/H5tlzqPMEv8dLDDcTgsbKQsA7vxpwN2fB
bqEuzYCmcM0gVGE7VWyZ4YDfLBk7/ZZc9BCsGi0PDbAbR1zaWU1aBJ4FuoC00+Tw
FhNzQjNA5B6v/uh89c/GCgS1NbP7K/MW9hrEqdzpGU6rhim2NryPmvLF572vBQe9
FD3rNfcA1ebfz4e1NBGJTQ9FXHCseMfDcyOdcQ7aYOTb3/t8cFeQCvMni3F03H9N
uOMadB3sta5TnjUrQYsB1akF9b8UssrWk8FVvHG50WDeYcFMtVGImBYMtQou1kn5
6tQl6sapUhieSCVvRDqKMQ6bc03VDvvQusaLDyUdjjHRX4GUsPypKCUniDGdnqyu
X3hho5PKI4XEEMJ9kdG8Z2AaHdzgOZt98HRkvdPSJ1VvCjbIvjZ3UiqVtAx7Vvl4
Emw9XbcHThrpccIlI7RRXVVNzixxwJVrAEK2Yq+uzhH/fVM5/k2p+c+WyCSCW1nb
HiBkXc3+lVGjcCecK2VVZR76z19n8yLdFbJzA2xQCya7DuWiZ4Ee/CbrD3GLlgkg
g+yVc2Fnu/mB38l34TCbHYwnVVI9OHLcx0vINhNaJKJ422uie725TACCFTQ8EpQt
jITLgHyRQ6oeLcEexurnQ/hW1mnfDxmHT9SO/Lhy61vkxqIVvXA/J1dPoeJi7lN4
JfhoGalbOUFMNSG1dmh4yZYf18QJQbNjRp+mRGG9xMUsyT/lWVkfMo4kCBAcw2wa
3tOkYJurdUzXlea+35NuqSALCq8wGc5u7L0r0Fq7e4hDw+J6XsIP8TcQ9hb5/rM+
RChsJ+QwT9CHTxsq/EdpZMWMMcmJJ+3E05E+wu+bHwWzgReFYJIkVJhYZurZmrJl
dX6CI/gsEPMhD7W+4Xc59yOMAh4qtqd721eheZS60CEnYK0eNy+Y4zFXhMzep16Q
VFBDod0Mn/TrK2zutMsSta2Ld0Kau3HaSaGJkbKM7p76BM6vZtcOZpoY4Uzwt0U/
toIMgmr9UthGIpsFvuuZ4+8KHLU+gtBYCIeAYwEFsAA3bKg3h3I95s/EF/8aiti1
Yq+NRhfyuWFpeipEDPNZbDYjDOlzQcxRJwy4UYeQAbJdUV9eS9aXXVbopzmXSlPo
LsKYgH+XzCZMsf/GC65yghvyHEE/uAtEqdOV+2r/UI0/iM/VM+AbkfN8xu/Ia+cW
rfyg7+m3wJgHHw6piUmaxWuXON7xFb7uVknCb1AX62cToqjmtaPMLevv8XS/uLsL
zCyPhMCkgBbRS1PRY2S2I4ZGj6A1BUKJTEZR+YeImN7RQ3iC8opYmgekDzIPtbBf
cNkHFvEx7q5rIisYodiL8D7znmOJ22Xeshb8QIwnfhlXNGZPEo+WQlxZDLkTZ0EH
GeLVRrwv0cLk10+4Mn2cPWUnnqWJztMN1yCl3oXJevD3jafI0cEN3OVzsu5fV0CP
vRA/8W6DvKz7F6Rsu9eYB0r9uMSSbonc9qxtuzbNvaSpMNCbhBGRtmAH/JBJrwYe
IBJAk9d9QochEM0uF3yTKFaoZwYGpEhWvv+8mwWaxFeqFZshQdPxrusxNfi2UpLF
O1So1eRc3KCB6cP3lMWmP3E+yYu6UCJpxhnv8PcYOA20sA7vOjwsKSHLFEAjJTH6
e1qb40yh8u/2SlLOZbjQOsItc9lodFlZFvaD0Sw5e3cpiM0FcPZKurZAk9jG0zGa
zqOMvKSD7nT6Z1uprvOHKspXlaSW+nq8dgW1OdWmJNzavzuIwAaxe3SfSb2xBKTZ
uZmgFlPLdAMV+PIVzawp6U97XzhYszfNbIFPLuxolPelC1ifdiWA9huZQ5lVZEt9
XxzkWnDA4g/Sq9axlSBhiQF1uSNeiX0WFccrYTWiPa/aTYqduutzfMuebjKtgQ7M
yt3+hnV99xq+wkP5t9vIeI/PJJIN3bIOETRvSyyc9UfrlLDBhuGb7OAoVc6Lim5/
Pf7Rgik/SSmqagbDCqCQ/bYxi0Q5fZOJbmFJN8lAkcLsHXxutpLUB9qmT5H9evB5
zpK0sbphlhsjkGapHkJTQ3cjbHhS09+KU8YYCUSf1A3sWbSXslsixPsTmZg+QoP+
Y+A+7BY4+Q4Az4ONBkeY4QDTp+h5/NWdtobneco/O0FCZDgRM6A1PqTZXG5aHp8x
DJ5cTEvgSv0TlgzonEo9x/k/TWsPi3Y8mH5FMF3P2tFxwn5VzWbrRDayIhstNG4M
013JWnnCJKjQFlTjaQUcS46UmqJatY0zJBTNJ8QDk/kQdTOCu0ykg0+y3rVZuuwI
W5F+wJKIj6GV0tAhSn1m1g0Ttc6g05S/m4UDj0hJZs25E0F2dmog2if81yfJ8BEA
c6igsjn2YREGqud6EZviw9dNqyNUi9D8I1G3eyIpCB3h6uGH1JDBHlbRBQRN4Xmh
1BFKCY7ua3eCS3yYtFtK9XRRiJE8mUtPS+dkVsRJPCZI861vpOUHWK+J3/0xhiL4
miIqWVuL4QfsjXVrSewVyr+bc4IsMbYaz4iIbt6Jw13eQb98mg3mgjxn3P+uRAAy
wviIp324+vIMPBBqk1gS9ZOGzpAkaM3IxK7t4LblrHxmKux/6M4rCoC9sqyISxJi
bbmkxNIozX6t7b5U9rt+5ryYDNsm1wnh9HKa/543dVQiKIXpFcMql4T9G2MvrDEl
oSz/Ac44QFT/XsAkuQ97j0Dm9EKDEcdWjQjJjiwllQcVoKdfTc2jcOaZVF1ZQ+7T
dpcRgZ7zljprSDlsPAAMKBwBuU7OWAqQKVndivEzmb6NRV5yNpFysMvMgdG+WzCN
NP0tpQ6NaUHodx8ijlFqhAbDY0ddiC0ce0wNpDF7OOA2I0lZiHMCzWBGNhi00/Tv
6ldsJVDKGdNk3DDC2knMTwjByljZy3MFjTdigJj1ylWVvdw79f/zfBWCf9nN4Gnj
Oe6zHugmtE5W45pYES91Gm3PFPa+Kq7IQaYPMYeoTKMHbkocjFseNBUn/KTROoIm
jorkGNVfeWtoha3OpFeN2NQ6UQPC2zvpiU/m094FnJapLoKe3sUfS4QVQxBEVGBk
4YoB5gQW4oVtsKMKzoFrAPJICxwDe8hVORrabe3l6wvN1s8u1JwdBIuP4NNUOfAf
OxRLTu25MVZmEqSUVZcvs5oIVkhHRQrlQS9weHG+WFlPx8TWXnTdJUFpG09ljvSl
jrJIotMl72QO9wOdsujPHQoZQ2bwrwTFKawCavIywmf8m2/bB+4LiL6KqxnZJ97k
2BkWXsJUMK9qk3VHfvyiVcljrz5VV+Hha+fxuMSXy2fFLHaMYe3TE18iHtfEJNz5
M6QL8ZmHmylxCkHpTKyccRGJvDWyvmVmJE7nMKegGuXadB+spOS1aVnAGDzMxQM4
iGTVdbdTcDh5Edgn+errOP4wfNsqI1QeQbU8IuPE7uYbPwA8verD3yFiGRpWkg05
mLnJR2rA0Opb9a1usx/ok3XxfDIwlf+wXdZig+wcuEqT4MsFuD9O4S6ACDo6NTrc
GkOOBlSkbdilntJDVHO2SsJlPbKM+VupYNT6evLtv/LRcI/q3wq86hxBvIUPfbAV
Cy8I9xkO9UIO/10Byg7LxY1PiM36b8X2x+5tnWt8hjisROQkjNynuIihqMpTUy7U
8cY9oXLRXXHLu8864sd8skAQQN/BnxwBmTfUs7Ds7l1ibOIlCuUQaI7/95UvngC/
9kMeDtxlX1jKPXrk+7qk8IDtnnDaLyJ+46JN0Ki9btlvrgYejx5UB6bcTzBcqVDc
z2cwBif9/EgA5fkOBiDvy4fInTRF1XZJThsZGK93vDVxLkdQnzq85Wc791uaZtuY
PywuSguDR0i1u9HUy0r9vZein54dyJ63Q/1XPt0dEU4hFCsgHj90dLBNVgAyGgZ2
pnNUX0F+ixGW14VmxZpAskVjLF9sc+PY6I24hq3qDjJ+ajvyC5H6UvqDXsbtvD+5
sDzY0PeevjpjAfpoJz593jYWxggR5rcL4FuEglotGYLq1W4X2+8cwMMbjBu4UnLE
vYs4VdTEz1H0T8rOCoBhhRLGb80RxI1adk5VYzYcdZ1JzOTzpD6p2OA+QM4YYm9+
Pi6mV7FIiGvA7QYzUcZ2qSg2e2DiAot3bJl2uXmfFamc5l2uQFngVFS6UL/BSv5f
mZj5lwkthoYq0B/6up/Yv+WksPzrH63CCcjhlUIeI7LcGKbXocKx9Tvju32qic9E
xM7gvdh97lSqbPSe52bBFYtMwx9EDkhfq3n12ahcOfzuNYTZzaDKSUXXBv7W0eeI
AZxS1ABSuab+r8Veva/mOt/wK0n0rvYDfnqd6Tj960Omu+U904WJK7ynHKAfBrGx
2R4D54X89b5KqLywEZftWBd/nvXTRCEua0mkkJeiNzSR4x5oXjsLnwY5+V+De3Fg
2U3O7XyMw1Cx7qfe/euCpUFJ9KA+4zGdK3z3G/QdZ32lXX+wqo4+Z0Uw3jmwRts1
KnZ1hzu9zQFZlaGLhTDEMq2lfdWg8EGIr8jCSeE9fi2zviPZ6LI8/WCz/7TkKIyf
RV5jnESPSAcjpwbGjVyyYHj9v5KpfFuuvTGi0WZbMFp7SeMLguqCRLj4KYoJpnU/
63grMCio/Db6KXcKu7j6/eQzzIyFCZPLeGmevSogxM/3cJ7D75kohXshQc2soqur
bM0IMkIaQIIW+MU+ZVkIQ8FbgzujS2IG/fC10Ay4xj/BeR2aq1MXLzEQhMCb8SOi
MuJd0FI9SI4TGnIgzmWtdXt7bDYNpnYbAwipXkCCIKbgxYoOfkAwb3Js7Y0w3Wki
+Fy5ig2kCue9bjdE6q3wW2O3a6rsIFEHWOsTMl8GNy5rRpiGfDyuNy4u6snFtCbm
Xt1R77NdpGLTIy8zZ1mSK1ldpERttsLsuaZ72hL2QxH3/VJUpa82BXEPgjhKiI0i
vDz295VANdkj4KZ+NC2QdPKy8Jhf/Mj6uqZXeoNNphn31EBKcBrKE/Qj+Sa4vii/
VEKZ9+n9fIgBBAUeL+FpK+3tkAMncBkw9LiNSbQHGwZ1VTYgO3j8RHqVxzPSAUys
M6yvXhWX5S+2QstxYPqDnwykEQuqWCarzsj7AtSprvOKCDJPMkrflZEEzUCC0ukL
SEsQcsL0XxHEbrFsZH7I9VfDCdcniMKCGjoSzrxUfhSIPueDKAmb8dF8i8sDoYb2
QZw2wd7ADNQOo2aXovUZ1f4wt6RWiYGAqrnibHh9wcHCV8pSPZVoWsdIW7t7+cZv
a6E7v9Z1jgQoAIFFAz2Lmj0PTjwPJLRqHD24S1gBq9gZUZD48dGYJmEHcDodYPK9
thK8Dt5pjV8bUbVRAV1B59LLyBcpd/SIDdZ2H6isaG9BUs/rxNTN6F3TWWuIWTpA
newyB0PEPt00mjoCwKwcfgmRD9i6yVraXZx6bO2KtP8aG89WjaHT3aS8W6DAAIZF
ucBwToX6GLO0HUQmEbRp+sGW6W+YAS9Zh5gvI2HfSYb6Iq2awvOEoaVYW0mjk1HZ
fJshgzxg/wRbb7cOTWutWzqlFJG3px9NbP4fJH3KkRQh3gM+EFLxgrGmldnkwLx/
Qj1OIE6Wz/HI1znwRKIz62j/kzR1KpASbFGnNX8A6xVwdAVMEuw4C/7UWKnPm4mr
7RHAuIPU/aBXo3c72ustYx+bGp1Nsprb3HGxHdEgc56rqmR+d4cxASq61v60/o/m
SNMECJC8FGxkvYXDGxEF6MtbAWv21KDLvkoXgflzOw7xAY5eNGZHZXxpVLoVLmHK
T9/WQlHkAgrKuR4itJxN9rsO0QR9vHcfnem1Up+Uto2G0ZE4AHJhzcqp8Z609hLZ
rBn4g3f6HrMALbP8XuknvYMhOrq5zwLrmsnQ0qhuomfovbZBZJSz3xBxmZRchN3z
Kj5e/7w3MLgPDJX2fAqaxJDBuFyzU7AJjcsd0hB6Y1ktBt4nQiu221FZIr5vENnI
/eSOxeVaAEphNE5JPaIE4w+yUSCqOmmYuYVVA1wowgRJesPYw4sFV1567v+ZWVL4
zkqqrBT++QOGJB4dHWEM/mbdOEMiZJQrJJdHyal6Qg7gxIs1FNEng9/AOBL8RMaX
Osd6EtIQQ+GHLm0cHW4CpNb4sojEFiYSoikZzvNZB/jVg+Ro2eRuqt4IU29QA5id
eKHm3MiIBkN9lTOfsYKPpat4JW6eujf1hLywikFjfwH3qYDImobe/QAD4mHJZWSs
tyirI7Ia4nUe+tYAJH0yZdpeWenvuyIl+5JkeWA1r/3seDAnr0jckdGZGYMlF0ET
+uFF8kfnPCkLebpVxFg62wumx9C+21TghXjD2EYaSLCWznAl78TdcVVeDu9Mdc7j
cbEB229fW/VwDGrzujxM5lyKbSSdl9MXi6tQuoSEztkek+lfeMQ8ka4evj5W9CHv
s3us0ss/x4ZZnITqG7f+Yhr6FBBrNiqTNhNVanthFm2xb3j3WWG3HuKNL8j2/+63
KUJUS8irc40W0oSqIv3XCbMYVYtsTcdCDRpsdIVBtKxIDRbr3WdryUKKUxroZdVA
mnE5ZUgyjqv8wWUvJE22KOxvFQfNZMqf0CF84XrFCMdaPD7n7U8SpYXdomGhQyyl
hCsvGG0CwUChjWOts6Xb9luyQjxBqVm6g4YUbMeC3cr8G20+cpxcYh3hfkjfG4lF
S8j1Gs+1B8Ci76l+FGhvfD79yNR9S/5+u+Ow2c0catG42ePuba/mTMlHQ5gWLsbn
iPqW1bxyUuPTMdD82x/fFpgo8JlQnPaEBNDkuUuRMf4VonlAGlA+vnhWr6G5blM2
Anf5J96/pX/jHJVlTYqfLj2Vk8slxsyaaPaRwkZDZ/pBBF9jXP6T91Gw07Of9Ccz
fAN+ndfzWEKiR0VX5tcdAbAjPF+NY8c160OKT9WFTrTuH1pHzGAM4ayPd6wlalTY
bwR3VPkIysYgm+MDJRBlX9qKyOgQcLKrsMtU68HkmyOmKRMmjlrrrIx1aa3SBQ6u
9x3uz9fZrfZ+eM9RA6HjPZpfGB5z6TZNkXJ0dc0fmXgBiEADvWXqBk+jD4B4vVxi
uU5zx2MiNoGk3C5lcBvhqa7J3+nfESXPmmD7AyFltmriAnm4PLDJ9VZ10fvv4Xrn
CZmqsjWlEn2kfqNfkLxajXARN5hn/0ozEh1g4779oeWaDKEeg7oFRypXEceSevne
W5GZhr3G1FtfUeRQTUNjJgpPzzStWSp+IMJGREpXQ/GnAFvbYZxBCzoTNxO7x0i6
wBN6dkJ1e2dHEOK75DTT3RjrhPzbqKV5uIDlF3wuRLdVuSqWJG5wnI7Gr6VkEAWG
YC57f68uxLdDT+9M6XYo8wImLchSzpB+955QsQ07HQohUx5uXFCcN4fm+QmVUgmI
yT42Agc+FvgjWi6uyGch+3vpCe8ciu0MyeiyMsxIvxGJUp+gvl0fe1RMGQvnpnCZ
TQQBLMuk7nIjuHtkpGc+6CaGqFAYefSpHQCFU01mnetOMkmryTPbi/OKxQ06yPAQ
CLnFxsE8NOsbGtWeD/QsGbOzH6WlCTWVqI4mXZaG1tBuFhyClj2knOu8mG+gEkgy
vLATBlwTap71tBCCz6/89grOv0LL7PK0ehtAg5GE+ZWOhXRHE9f+qZE0gC3hO0Km
yDAt9YFBBQ22z+OlA6TO759S+uiyhO8WEAMyJj8S5Yl7XBD9beuE8VMIuyi53Mle
levU+FS4x38SWPS/NeaQk86GJnU0IYULxGOfXeYppOUpqP8j4VZykpWx7VjY0IgJ
eROsJV93tzRapjg2GNl5cpFIqAyG+SgPIpnBv71COa58znXM1La1MyXIgCBc7gC0
ySmeyi+lQmtfVP/pjKjdIk5uFjJQsrzp3MK8EZmo1P+YMXTHmChqPaW+qXWo8GJt
F20oMXwIpzStf9jI2t0nrHic+RYAsW2+fy9eaE3PbW0epV9W0/tN2SsZk9ehBzw7
gqa9DgB1ivK4ImoX+QFdWMCyKUNaHN+bzcWpk6aww6A0DzvmhkUf9VWxiMzT40+K
o+p5sumLQXrgWRkXRneduDMBqwUdR+apEMufmmbZ7UQNtU/XHUs3eXQGbwoLDJXo
LXIFcPpdXyTjYviwtsVvQar3s7LswjQslJ7VaVgG3zj7Aiuy4XeaDddyePDmUbqp
YTkIa4xWDTECFGgsFxEmFgjctfdf/Ai3+ZWHUpi2UtXaC4k5g3rK0ujf5TGFcWp4
sL1QCU64PLHK7BS86FlY+GZeEK0vLFc3i6DY+T8Ys9IZS9Ewt/rbjssyzF3aBN9w
XoliGWINtnAFoC70fgA070iYjJ6mx5Sk/48uUM65oMHdxgW+mdi6zdeJp0pgbaqo
WOieR9XOFTfQAGnDrI7tyYn/sC5SXHvid/unxhv8z+lUTqnCF2lLyOxLwaH+AWcs
bFrSM2AUFUQa+5x//dzxhAtKnWk72rFz3N3Cv7eNYHbuBmY6SuSlQbzmBbeXIBrg
OyAEmdmTcVnPI1O/hmgCIHJ8N1S+843/dS/KCZX0a2raRUJyj1A1DYLUCS40FvZF
K8tQuni5II1f19OGdE8HydRp7fhN8FYW7fJCw1vuUGj1ULkb1zt1o5Z7H29lWKgT
SOyRBp9gxYxhw03DeMv90XSmfx7aU53wHD26gsLKrnA4bstpM/1IjOOXmdWu3g1P
mLYikfBCrEYcsVTRz+6hYLJq5LSKjm99dLdjrMZNO96qOqE1EoHe53k5oi7cWcfG
4cugEln7u813FCbI3KvJnSgIwR3nHh4nc0dgqaTVn5qTD1bEiSH9B3xsF0q5t+uT
WFXlXZxRDtJFMapJvj+nH5JMcqet7+pDJPcIicJxGaILKHyXwOeCnnAMxlbr5QWb
Af5V6KriD8rcPT0RyWPVTcXqiWfgoFZhCtOi+rVHi2t6bRnqh1VurDpEpxrnBcjo
z/pndnes0GWoegkQ+el/whlOvXnR7+IvyJALSUbJ1uF6agctM9TaGnxeGyDnk1wq
q1zj450OKmPHt13CDqm6INFLD4KKxa9/comFDPRLtgtjSWJpqYSKmBTxfFQVtVtH
jEcKdzdavf3CGDIc9E08PQjwa2f1TqagHXaamY7lQNuoBMk+4pf4OcBX17Zc0UPg
Jq47INO+DHwt9x1bfaA0ONXXE8wAzP1A8uncY6T03kkzz4FKyfLfIcgY3RzrNJa/
2lh3lHg2jgvlFO/cbd9wz5UJZNXIXrsX/VJxiubgJ6ZfHptOBP/N0eevBLM7RWGc
g8NpDMeLA4juBVp92SYvF9l3ZPwk7Ra1fV8XQ2zLf46nWuvRKXx5w2K6O/8/p3JW
yBFxwjT45JzpqkjmUX2CZ48SIo9naaYzNvVzzRj4bjz4hz2cLhVvBHMLjN8uHXOJ
t/C8W6IvM2av0N+g6Np8JE8x3L/YW0UVUZFWapl1BbL+3sSQAZpT1YvIKtDRxmyD
jQr9U9FEuJ743uXiGhUBpRLybMwyXSjsl5qHOHUu39bUwIH/paDoOotYRyzUfIot
ZyPP3jt40YJMt3IomqeiIqMwiNakISozyjAu/6zbhhZ7sh2chpkW5o1Tomj2WoOj
UjY7vT5ycKDjaAgJCI7VfbnrdseAWs7LUzxfJk0fXa5CAwo0LR41SLJR/F+GAdoQ
ThG/dh0HHv8tdi7asrL2Ii3eGiXWaeh1tM2DwLMaTSZqH6Fb6MS3hLUaHy4e0n7i
DFdjVSsuc6lDmrHRJCXDlOL+2GgqB2oPm495nFkFD4MGDyCXYwsBQLsvaEfmGnsc
mbFp/8BK6n5r7zoKQRUc6nWFEcfpX2wt8bIImyBeKZmADPVQNUgor934dJN7sIsS
s20+e/NoJoCjCXDjvLfLroCqrd3IpRUu+4qTliOFu4zNsy7ME1jNw2nVI1rEsYLk
0oxWzFTz7TA/KExLWu9fuW6UPmwIphtHBDOqtt9ddwGaUbSuwIHXQAS3J37uPYgv
FqVCU5kRkBXzy47YlvyVyJq1mElKNHUApl8U1Q731UYxoo5Cz/xNz3QdxnwM8M3z
W5tASoy2tkV30+nBDp8j+cXb7UV3mJrT145TAyxRS1eUiW/8crfxNC75fZsKE5FR
UGgD51bcKrMvpwis8JLFpB4Hi8z1BNWnUYKeznbDTzqdOp9bIVom2d5f+QwrR9SA
U7Z0BZ1/x2XwbCc8XJP79Fm1dcYH/WW5srm4oYOuAt160xeW+0pKNtmgjc/BZKrH
oBNkA4cBf0gJHW36VhjHnWi3j3o2Rj1J/6R0l6MyLJ2VVJlKUTu6+nu6n3a3LguY
gRfJJu37eYY3ap+jQIWwdzTFFZ1TmDDxDhjBErCR+emaQgybCM/vIwLPkqSBIJCG
Y+sHgJ8/vsKzBeTUbBqwBD6Ii/n4iMO6vumqnGX8aJA=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lQ/KnPjdMkRLGYwxj9TaQGbCPrgII8+fEM0jtVLknVwp2etnVEXI365yyVphnPbI
yu2XsWpzB2Miavr7hCqZbggxGBD9dpCTTz9ePUjUMsL/0jySN/XJdPNQ0/XSwU+M
3ZFPIBVwaz5fycFnun9WeDjwhbV9iZQL6h7P6hyWPiKQWSyW26b38/ydcCCzq2h/
lOvDouQdWlUY+ypH5rDLv6ISWqTQ5vWcl0vRhI/tZJXIc8oshsaBO2pvX3/ijMsz
gkM6Ftc81IhwI5YjaFYfSVu7Q8G96UMRzpDzhW+294SaZ5GyFG1xOTtAK5KSLqaY
A8cNHZGTpL7VEi5L0gFhrQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2704 )
`pragma protect data_block
HgT8H0Kex/5/npBBSrEeVnJDZ+kGE1i8BaGgDFK4NwzdYUCqRqArypFrBgEwUYUe
+e0S1ny+Mdny4pS0nW2E5aEEE9SOAA3AyU3ecptFMqGn9zLkAL4BD68g57vtS7gu
gEQ0SKFs9Oiq8053VAZ0j0BUBMLcbwSYiww1cJljOXTNZhMSyx8BfeX9C6+sPv0c
QrAmz4+bBrBBEbDtbYsCx/ty6o4QcbiPHWxtlRn+UuqgxNfWRxhIIJ5W6TZafoyu
dn5WIR9nL7urNWx2efYT/lBJkluTed3rHmX3Z5chA5oy0e9FcQzVWMDXCC1qXgfo
hjQf4kQfyqx8/DsoWmycBnYqZfxAc1ZY45+HAosrL+LdvlpYlKeuhAld3ZiecamX
s9RZmcccJ70qcymiNwazm7AGUh/1o8imPLdmPQXQOtUeKBmx3XTX127kBYmS3c4c
bfFZvTJZk/EGdK2hsX1z2JlnWvxxD18KIQaC4CF3BdcUen7S2ZlOW/ND6XIi2U/m
Y2mBvMFCTmsB6D5gchq0S/iPcROV4eEjunmguJAC6zXjV8iOqoJYZ/3uEobQSOHN
cej/LCdQSJ/DYrFhlJWy+IEXa8IUqs8b9B6NWeA1eaSdFGS9iOAOsw0PClCb5OIH
bCbFuke3sL66DZkXoA6jBEGJrnieYy4Lt66WSrYAU4C3Kp/MYsnraRVciPMg/06w
1DGDvxGKoOcgj4rnS5ef7gbpI2ZcQc9wCbPTXYOCzRiHv1ZoGj6HUpjR9jqdML++
ysb2yj4H8wCLYa6+KfH8djW/UqWGl6KDkgJjGYmV5G+Yb/IrRu8E2dlxpxS+ZHMd
P1CPZUWAlLq9FH+J/OuLTaCtpXJ17Q/6MIQ+L5vbIoBAPlicNxbU+4FyhWj9w0an
jPcfU2no1nzszNDpi+MfGaL1VIJFx0tUHQZiTXQd3W0PZS5xuOLnut2ckkEMgom6
U/TRXcjQrqWSDRUOh+E0SdcdRTqIihykY5nPxXjrgHyBSaoApUuaQMuNRFiElIbZ
AM9S0m8/2DVMd8D9WVxh0DvB0c8ZWREoCvFXTcQOT+RKirAh9v0aHMxQ9M0DbqJ7
mz2sNOlarbRdvNTbsnyCgF9CPFS3pNOTPpELfazI4NpoV232YR/u8q7XnUrmtU7C
nW231yHhE/BpL7JQX/jSU0hak6LBHX4jWMddmR8nNSU+LJ+57aXmzfe+SsJujEgB
QyxfTD6tTKhZd5eX+2nAJVdiHrum83927HBDC+CL1A+8AgWfxYgp61DpVTBf8Mtq
akga28jrKsJq6QoBpAzZc2XZJjXrWkRjm7VVyeiHlNUSsehX0HIpoltYgMiFR2TG
rXkbtfbiCRiYK2lc3/LVaESfVkF5ZblKWMa+LVnidb8LHgSbSbv06Q2eopRpgXU6
ZhBDzgloHD5Is5v4hA0ZyNhrg+tHPUASfrHBhSVT7aSnNhSnUXvnS9GbfSbqzMag
M/XFyiqqvGVY27Qqlf5URTm///w3nlfPQZ1joywO8NMCBzIko1Kqux8X9BqXK37C
PAUYLeC+VVYVWuS1PINQRHbZGSr3KPMrTZ/nv8KkIC8pb5QDVFG/KSIkE7fUXbhi
reFQ7oOkvx1Iqfpf7uP1niq4YVuTer5xmxasLxd6gaMB/FuMcHLuWIYlPMqK9cYD
0osHrE3EgkRoVoJj10+JLCUCb7h4Uob2HYnKJHZ9/etuEIPfC3jh06ERV2wOJyMI
rUlQ2NZbjlSFrjn8urb3TyezZEaoM9hq9uhD5B6J3hRApH1qmDThdOgtkGa6eRn2
9F5ELtyvlKao1vJvrpMF4ceEQ3n9ketsbgxXSIUJdyuL94UMQqcZAc289OrzJ+Gt
Wx2n8Ek07dp31FMasSw+KYAGRgf9zj8AZkKIiJU2XhqwhcESypzWBkI1zvMXDJ9a
GRPSR6n5of7q/6/02ZPsZz7psEdsY0LKt9fnYRPT25aFDrgnBoGwAJscxsbyPJu8
VaAb668DOT3oB3cNIKitPJKJe8zgyK2yZq+rAAtCAAnTl2d1yL4kCNi4nyAB9jeh
BSQ2oyNNqzy41t/JOL7AqVj/gAEDNqQi5aD5AMhtHn0NWpY8tVdA7BqOX814k0c2
gonqKfph+Xx8LHn7TIu3oG76Fc8fIRYRRT47Sa1wjBq3piVgyErjzUPgCRKSLhUO
G+En/TW0R1hoD6K71KgIDnoJZrsmbK6Kbmweqmmez/51Bb6JRsBffSHHqkA6u7yx
6D/8jelvtim8NbZx4MfOxhx1YgU12DtVQyPySYczT4cxomM7gPU0jRFg3HmE+vLH
uA0IHQf6IZu8nLDL59Icx6NoNBKCtA+9B3Tq1IA00Ci10JrzQrwLSmOmakZr6nV1
kTJFLTgnizCuKWKoBMsdIJpAH/hvymMyhTFtxegOt4OnJ0HKJ9o+bEztF9TgPjbf
h+6j/GXYlr9qu4X0uguMGkv49F6U0+pIDslhJ+pbQ3RnEjP/VwDQJPftriUKgz1s
bAbmMcirXyHDqbF7j1SeBmHLBTDHR9OIhZkRJD5tCahrge0WfXBsZNrs52WkJnjW
KjoEjnqGrwycWQvBhisH0YgS0ZwvNL/fGwhNS3ayYHF7WZRLhTFrIsBZ9noGJUhP
slPg2IDz+yjp82nHoiVhVFMTpx14HrGBMT+IknI/hguJ0SJ57M2hNtIfb9XfkR7L
inEVIycVb4U0e3fxZ0UA7pi6voFRLS0fVW16JYf9ZPOOEyaiUZU21vOKjm6k2cap
7nIDNCNJZx4NoR+NszD6O0gpIqNRM/8hNKUJZS8yZNxtxpOnEUwFZF547yA8+hYk
Spzi2Oleic6hSgKWASxHVOwXssOLEs/VxA7cW8V0BGsZnQtQSLaBznd+VyfF638L
7DghgAdiwubEOF4/T8OAcaKRpuJCo3p4g4FPs5bQ4ZEP4etHLN3FVbElC9YZrw9X
Fp1tl5QipTqnZlONX7elvgyoLvirrY/osakIlRiK37OveFcf8ZblV/15px72/tN0
tA8+XJPgy01tJTK/b2SiORP8dcv097QpESe+82nTpnOoWT1X7xt7Yi1DFBko0YZU
daBV6+ouikrOUpOGaMEH+oanvNV1hjwyOtZc8Sb0MkRAl94YwjF1oT058bWtOBov
tjhkB1QD47vBlAp8Oc0A85FJGoQ48ZR6QEX1b300ZTqvicIblUv0nDy7bvaqETa8
eJ4Z4l4YuKaRVp7Q4N5OG39oNLMrvSwQE8QIKB2mrL3UXTjoRQFaV1AMHuWrvZkX
oIGK4liUuOjxJoYmWf3sVXFRVpU2xjUCgUzCGgCdVLJAYYFtZTJnhSrMpTaLVIbi
B+zRNF+/zZUEfo32SqiFjb98E4a4Aai82/tEZyw0rghjiJgr7Bb8eq++CYT+wPl7
Zve7sVlExfChdspihWhbsnqOc2kbkcN4tjIRlluzAdYqAqZU4462G62lxgrzH79W
L3NvdUMg1q4edAwDDAnmy6PMOiFvAC8LHSOyHi3HgHVMDZ+l2Vs/X35jd4JPS8LJ
8n9m0BRz8myFkU4d+hUPKEB3WzzbrcXS0U0jRowuuRuc0r79PvP32n5F9ELh3rh7
0MPAhRM77PH9KsIDKlEfig==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ny2hqyWnF5vw/W/W7j4xvVpg810y2FWzxP/7LPu/oF4CGO8/k15H7/C4nf4Xmi6y
J0uXi1vetf8SMcwIlLaZ1v6mqNBfisSnhkvDoZ/rcuBw6xhbB9X94CLPz+iO/HtF
f4nt/C5R3eCyFeQmBaEJQTq/Zr2KPafko0xRbXtI7gC5vSW9E+cUOzgp2aWCqoe7
DN7EUn9vCDLOmQd5hBviT4vq8nohyi/l1Q8FRNgJJ1kABzL56zKquj0M1jG1xUVz
3r2pdcRIAtsmb39oiEo3I0R+rIL7okea8CmIuQdMr3vDc/xIE3Vc82180D+mqFAu
QQXjzJzIxbT7Pp9FbYk2FQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8048 )
`pragma protect data_block
Jbeu5A93BFT9d+poQoj4mAWDiqIhmEr6WfG4SNCI7x4jH7AFvbqvwZmc7Q/aCHFJ
VdZP/0cVg3hI2f7Rz/YnTeUC/iN0dz99vFtFcl8ycwv+UgITz8AYNeS2H544mytc
ZPGSTiBTAA79+kasKIKrgfRu+frnAEjwNO23Y/fv2qJeN021Oj0A2ib8+R06TbQ3
PkLd1CBeFfAi65MDBqAUDi2mQerBVJoywUY4Dnlener6VFalz8Kw5r4Rgwd591D4
poJnRxXSK8o7QKuNjMd6vbXggMWwNhr3HUb3+AZqL+xCl47FW5H0SNby+M1FyzUt
Zo+WeSkFiosB0w6aqjNnWEHAKZ+acRU7FRe/Lr8NUl4mmDqAp4gbmGn7pVzNPclc
hqn3HtPMBtfFOCRHmAan/U/O1fjD8Gb7seCkyQYk7Qir/dDgAKOkWwgufxqMmVyV
DWfotD25GlGG3VDKFXEvD465qXY2/X0+p6f+KgrvcDP/YxE/v9oPA8W53smuP+j/
px47l9nSd5APJabOMQ1mrnpRoaiiwnd/UkJMyJfmQowawcna0EioRaKP4eSEk3TY
pEWLFm2VPWVbmipn2wBXb0wDwDdGQ0ysEZ2lQuM75XEI5NCh84S8jSWJ1j9MG9d8
L/343qeMKdL8FQrrRlw1uY4orcS7/+RqqcKxH9e9Qx+hEfW/ty8IsB4UvXMWNIk6
F4RaKeatlURVntPuCqyB23/6ShNcBqX5JYiavpWh3GVzz3CdiOubRX+uKdee9f2d
+hEsJcrb4bMXRfcmaXiZEtwkOhJ3dKp5U6PHO0m0Ixg74Vf4x2LSpEXsO9nedLtp
3ThropcbgAxjWO//7MTr8Jp9LL1VV+t9yLh6dNYLYugcBNmRqtyW7+w4kbeEmWzW
N7NkSCEqbbjEoriUl1HzD5lwCOHcjld5dnlMGKq7pVlGG+xml8G6KLCVY3zxyVE+
iOQggZkyivCqeL+KKCnJQhNcmRqbgdBW9S6uL/rRV12j+qG8Mv6kYf+EIKT0Wo0d
TbL3E7ASqqghLLRkMvF+kup1aKWl1Snf+mGIYQJiSNGHpWBmIN0QgR6c3j4ITRL7
snLzHqzxtO442iyX0SUynpp/KzK29e/1KX6GIrEeQmPfNztA+smwUYAhM863gt18
ofKK+PSatC1PVit0XsuU/kmJkkFW+G5MxQGkQUCwrXhLYEAD+aoF0OQczKyUsDhF
pK3M7sprAGPDXrhYPoD8hMoV2a5eAf5Idrm2PmPylFq1Q8m4sj7OirXproVLkIAY
6vAlE65ZBNdGQTBqLajd0by8Qlssm6LBcybGB50E1fpJoDhLSibYaF3fFU2jlbV6
1mcmZx+qTgdd7L1GJ009gGI7+eSfOCf1ndVMgveX00bZjZmPnR3urcgMQke3mCUX
VBBPtvj8edDLuXEnch/SjF5KBIJR81tJGNqj4rAQGx4qaz/YOpRBnahcpA2gWf1z
12MQ9Nz+7tNLvpXDtn2QGg5ttvNzBT/vGT2s3MSHKA3IVZ84DAuyj6ly56Jv47Ct
kCbC1d53cYYJjRxSfeVr6fXOP25avgWsdLNEj7cxI5oHksUJMqMAARaI84/Vccpg
hXknf/i6UkB3jwuITAr13DQ1e2CJGuGmXWA167Nv8hwof4/H7IJQU9LQW7mSiCCG
IA5bom7hD7PoRTzbomhlpVW4JJaZnjcefmZo0F1J9npFZnwmMPvLXj/cEvOLTDPV
UTIK5I0ByGyBHlNi1UWTymwWkIyCLLNABLGodak1Xh9Lsxu0y2AtSIVOZyOcgSlf
j1QncD8Y3JcfHePPnLnQ4gQY4c/YjQqhGD8iH6EyThURiUJarxOjerhLvFX5XFor
K0bN2PyTZs5yz+SqAn6IQ91ysaH9hpYZZNEBmX3Jbt31qvs5dyoZMD+UUU4T+hST
NZLpFPxkmUG+tfUFX8niF8m3qyczgMKmPZzk8raTySfUgelRcqBWeLi+j6PCA1+D
0LEkDUyXD6gnGRYFWVlDTgtWl23flq4fd898vvsLeQdvd9tVnxoKMb7PafpZCnE+
jOODii8uGxEiqHMawqn9wpzdLUDV+MkmzqsQ+IwfKQ0N13jVq5xA3dY9dOWHyaao
26VQA1CEk9qxXRIXtUz/Glh/yU1FFpkkRhcgND/zO36cHqIWduhJW3sx9CApxCnk
S2d16CxoG8Y/qaI7KohWgztax7MfJTU54Wh2Pf9bgD3F5J2OTTfo6u4dsphotOAj
qhiENbc7AINsreq0CUk2FOjIA2hGG5JIewnzDw5BLojEWBwe9EzOcj7K6PRF4P5G
CcM9oe1dujoQxW1dlGeQBW+NrhwobLt7wUmr6HnJpKWgPWKx+QNli0ptXYngVKZI
Czp0R7/4TT9RmKe6ItEMo8/zoEwg3y0sdpZ5FRbjkGgkcWONECFa0RbxlpVxbsnO
kTw506ewSZVqlUqmoMOiLsT2kNbtQTn1ti32Jpd48r2cj76qGgMSg9nFP2iZHvE1
G9xQmxYFEI2u8W34P4zdo4ZZA7bpl9ISl4ek8538PMlDQB93zv9ngPabza2ksDMl
kYuPAzgTxbMt6HaF3Dx6dfok+dEpe8y5ht/9MHSxYFSYxd/31Hy/BnQ2Di2fj4Pw
n5OsG9Kp7zoYXIh96/RAuJ3lvNgVvVWmYjFG6Hfmbcl927195St8keEorflcUJMU
9zhdnPVPW+08hpGldPRcYcP8EjZWFiqsgA2uSKfxiWwZ/GG9m+yPXO4LpMcjrFt3
UhTMimV2GmhYYqNVM7nVc2PjFoJBOuMCdC/NetuLMnUAEyEzIvC+uIB3Wby2d5Jt
5GcLhQXlxCgPUQjCtnS7APyeiucgNk/NadQODT9o2lv10QrW5y7EI4SU9QxuxF6u
CDNIWo3/e5CLj2FErQrjUvJ44EVZ3aM3JmoLNQV0YzzjlgBmWSXpSRUxwDGB5gxK
Y4kqqWgOYk6VYJplwVJsP6H2Y63EgUFmUmjn+2OYJs5k6SzS4KIouLvQ3XuRerVt
y3WrY0ACmGF1AgtOg3IsXUiSNmCvoEsmy8cCmFCyAKSj1tuZ1LvcgBkKY+1CiZi9
pS0erdJ7UQel0GpQvydu1yL9wU+Wkxp/62Wm4MPeirSuJI6FR/cRU9LThc6wKKK0
ZWdCerMYB0HCWW99aIcZlY+Dnxpg01AuZjPO20AAPGWGd021t/hTrGeO9qDdqvRH
PK7nEeHcuCRSQkrJc/FAKmP9mFEbCzfySWHIKMam8JTpZCgudGR1mCom/TmRnubM
xbSjAwrRJztHWtSwYGlp+ZsW8rFRHuaOfqZuagyQpX4xAobT0zgtGmkA0Nj0ynpV
ZKiICk/4xs3Qy7e03he61M1rPKr1ME+AWrxoGNZu5SOQ2aMOy/0EhlMY+Eg7400H
xYC8LLyA8/2BXpn3NijxLsahpoiLKtA0SnD5ILya2KaFqCiKiOVhojGw+qVk+bVs
rTEy+al/gnx9BDVUG+k6E4L6k/wfXy0ImYD/ZilkRoTW5gg+TyZ/w6c5h17nINZH
37MBaqHWCZoPVwcPLSU8wJ/di4nWP48FSbQdTBIDBDFXZtqJtbcAibKAIzriUq94
kGBdFGqyjALwnlPPobDQ3YU91MSWq+RquOo3M8eoJ27rwSUy1fYRZwKVk7jaTw1i
zk4roM3gwhIqKLCWYUQDDXbaZBzXuf65KjeGvWH5QU/k/MX8bkKYe6Sth0Gqec76
YmI8BUp7zrL0etTRE7rKJaHd1yxCX3xzqjz77CWT6LdBz8SjJ6nsf7sWW7/2TF+e
AACQWXrpcjYVgBKNiQs6j0ghvv4d83G+ZKz3WxeUcgBnaohYNq5zXqg1WVQ3f64e
svzEnEEDSWzGh7lF5vXGbncu9tC+Ha9IdP23/d/YlTckANKptCcMIU9MGgkUChFb
l16Bu26D8ynkf5gb0a8cn9Ec5z9bJJ6fj6od1rU3Uy32MB4TznJm5DbL0JIbBmK1
20Zf/LtZQFSuEWaVo6GBueoBeMwnWYL4ARwdLpbe8teG/+7YOpku6eX8N1dxnmdK
6SF0riLyEBjbE4toEdxkliWFIJ2KN71/OrZlXUreYav/yZ/NPDUAZbjR78W/TR4z
DXSTngLibfOha7bqwCEt1D32t7alIyuT9+cxDD2gXjEeaSiPVTELK4VkqU1/V9Iv
jwKO3p7R+X0xtt0KIoRU3gV3uhYmNHFEv/JtN8a3u7e/UbdnPvSxSzm4tv9GrSGS
7x0I0s5LVKJfy1FEhXIPlpBSAnDqUMfcqCzsSnXH3pGBDz1WhSlDM73SCK4ZCbvG
+IffV+mQYgjeGA88Zk+TOKSIbdBKX3Cd0R147kDvpWVf3I+d/1Qz90Ui83DxwET/
DAB/Tr1LAJZL0izEqWrdRFn/LaiQYljdEOMvQXqPKA+aU9Xi/WHs86i1I0FSEDHm
tFnajXT07LLARhPhqe0hjycoa7ispOROxHC6nIrjtD7uHmw5450m4ji2/YZPMMZ/
FRYeubJ6fZVPRyPrTjKEHSjiQho9QmWYd621c8eCs8q9gFwEAha/g5JlFxvAXljj
ZltSt/2CVYHH7E3YHg+nhN7+5Tt7E2Is7XiGXCgbRz457vbsGhkhT+CyD90uW2gy
0CtPdPAhGNBgfnD9reHlK+h7OopsP44C0ixK/15IaJKb2z9XJ2wXCIHC6KSewy/L
BDKHf+UE0tVOEBQgPwKe1fDXoGFdJEVuvL4WwrXY2hqC7UgE+wuomqcKPitZkonq
tF1dVqqTITDN6zZbPcd/MXmfUrLedR2ZVNQQeLXfpCPGaZhI6bNqLEJsCeYrzGzE
kzYn+bk0j0q4/o5gFivBMsXfrNht6lD3a9vfqjKTnh7xTB1B8qFAqY2ZBubhCXC9
rvdarXw//zdq3ZWihFbEGRRedTzipjbKtyZi7GRcxr0iDXW2LUlSlM32zuPeHfZO
qLCPTD/8MN76EXZCSUY6cuF3V3cYaiGYpuBV3wOvlzuSnZ4YMtah867Cf2rSfQ4r
eWiSRCDE6W6bjpDovuOcKuHXIRzCuNG2uLvpttDLxJGguFgE/X1p8BbFAZRQv6H0
PyvY1S5pGbURLPfG/TzyAWVjVxTT+DVEUG8vWSnZ4bQ17EZaTDHZc2bKge+HDrL2
AIY8r3HDi1DCDA6b0H35cpozMAjxFP+U3uqTJjL2tLwOvEf1+r3HrUse/WD6F9uA
9+scLRwv0jsYEoiUSiPakDpubiEf0OvBWRpH+UzLpj8LCgw4Tf80ErhH5C7dJyf5
WPmjaor5D8Ykcqd0y1Vfr4m051r3FVUdCFXf6Wvk7dMmj8GdC77gkDX1mVV4T69o
U3A/Z8RZJ7l7k6i6n8fdkemdY/hBSZQkdGxpQHQuFTGb+rislEj3Arwo7Xoeg+Pv
rhi5pcx90AWSvMCJZdo666ymV6KU0D6wf2xsIzIA91CVk2gBSPdTaLqf+4rdKX8S
JWdTuq7C+G9Mmv0Ws1xXwJGcubYgn92Dw+WNnzkJIu3rUm7ikLE88yNp0xNzMAdY
Zvgymf6NhyWPYaK9SSa8bSubmMnWOsTYujc6DVPOhyhhdDwSqLv5zdHieWzP+znI
2yBmXoVw0dak9j8z0gHS8IMz7TO+6ZPt7/U9LNW+Va3TAqaef6xe8iXS6k4d3Qcl
+5M5d48FLPWD7Qn1nV0Y08ids98HV+jtTqdFOBF1qQHxSlr3mMD/rexw3Mbw6ZB7
AfdO4iTiQ8f5Pqe6rg0SuIjYm5nnst/SrNzKzsU3Cv5lw0soGaETWWa9d4XZZJ9K
ynzX9TiTEyc7vWdcumi10vlbWkid9Q6c30VM1t6Y64eHzNKDfKeLeSZP5euGo1Nv
1by0RZCnaj01wwLOGzV4eFG8xty+geXzxIdE46MUapRhxBk/Kqsi7OQOQ6soW3e/
qgYydZvCF6eu1QxKITwHckwmy6vRE/NiEMoTorm2MvQNQnaZ2u7H6qU+/xYs4URO
jqIjCn3XWhF1Psl2oSlcybVkA4JISRZaSuG8o8jq04Iub2G2686BKg9nkPG7s1IX
uEx8seAp6fG4zka9vVlpAwREHhqxPB6oRW6aoXU9iMKsOZuE2r06zHlgc1STGLEW
d7aZimQuJAPOIcZdzIlb6UArIkG29eir8Yj9vguyiBG94SL/c+maT2gcGbRyQY6O
Ejc7xDxditFqH1Esy1L+bLtMHDdG+asS9N4Nq8f04MvPqunvrdpmI+vPzjrYRMG+
xtY7kpMfpymp2TpX5B/zDW6oSClPZnflzCTxMLZX7p58YUEU9ir8A0/APcIRAuKW
w0RMFzdprx+1BCDeTAs+JYLwgg/abNu1iTtgPXpdFdAm1rjsr2BAlx3rgGBn3ZW3
CjRaa2znGzaflbGsckNmMmlTRaQA83pnKPnw+wxmu82dwK42apOl+aB2P5dD2xWM
KckTxpfbIrST95bZ1U9HFPrlP1w/0oOJ/5SNJs3vYWje1lEOPTqh8B2u9CeebzQz
vF9xRoq7OaLoWr9b4GymurSNpaV+WjlB25ejzaOQ5dZHG4NMguxUKXnBuLzdtX4U
TB4OIt2TGHq+3YW1FgJyi0NnyZAueZfcrcBb8i90t0p9iRj31cLqEv5g5X7iNjUn
vmH6qbU8Q7n4lSH1qc289m4jbaCjGX/BYdL01Mq6a//sd5A+uN+oDjXBzgEqI8Fz
4HpFlgtpvMWJql7MyKxVMl/0KFzzlAcXzF0tSPTtXMfMOFESozywKGg+roRsY4pg
rsgFSQaxVLW8jooXzAfmgIOuHL0yghP8OP5McjBc2i1Go5b1Xd7JM9B96fJAvdf8
5+SdUfr5LmLl0A1w09G6bk9JJo1XJsAG68oKfuyWClObZomER7IC5xyD2ygyK+wW
rG6rr1UbNHiZ7i155i9X4sikmqvoUgv0a31HcwcqWa7As/vXf7Ueze9nwBgLWJy+
/tVqDtYg76OFetf+Ck3PTa/km+lPDDH1+8/eBneIIK2fb6oGwX+oS2zbtFNV1sm5
xdKoQwzj4wZ1iLZBy/XkfcxY8+esXqtOyVdkYhGvGgpq5RPlHb3HAwkIPuEzbIt4
Dmg2PNiOu3vjpF1OsZ3lyiNXlt4jetveKfBccrlQbpOj0ZzNfCgZxm5moKz2by7w
hN5urO8iOdd/VjA49i5V6fslIU+9YALFciMdIDab3zf8O2O610DQ41EjI9JaXzQ8
QGO1LnvoeMs9YUjfrCDUi/vVDdtxNPbg79rPzE84A0iT+k0AFtBfLMw2jSAlXpqr
injh8tSfen4q6AuN08jZ+JjUnczrzh+vLCI3z1fkmHstmTLPiJCXNJRfS5O4JXRU
I/Zkt1JbqIMGoh2he1sFsOo4LQxvKakjFswQjdtL/555cDxyRtJ7i6BD5QU8wbQf
LZ4KRbq3ZeDXdUCw26ofGDCvJGkSsExp95IFaQjM0HmMXztso6KkAC0AJBRt05pm
REL+zEUbRsWV4KYy+B7t3Qk+2ovmmmJwYFD1aWl1muLklgACpZmLobyepzV03HH0
KmaNCnOHrKFOA/6QPZbBXfNpJx1eZavcscPjruQ/8mo75wTCDH1PyN7+x9l0y0oh
8b2JPvnbxWKrXvquyjit+HRCaF4JXQT6+t1bOe5/OPaFIH7fmsI2YyoZ/tvNFtUb
MpFxx2kS7TyILSAjgVd+Salxvfi2A/8NnluKT5su4cy4XGsLPvxkXbmCIUQK0/z4
G0sXSf4PzZ/nnoxCao7E6Q1ME15zMCKqsg879KZyuouQ1d9fxOqo4QlZVpTuKsfP
CY6xYAQIttKJNXAHBOlO7Eoj3v7xSuLpEWV7l8E7YDfi7j0x9p7eG9LxpgIy/iyg
zUEzpKkYG/zqVoBwhQDdTQoqSLJu2wUeEn9fMSo1Q/wCRzYkckeI1HMuv59qgjat
YMaMRd1b1MW5SY25qrk5AzDZALzdX7FHXv2TzYYFl8brjULS/aYYHGzHQSe94juQ
/Mafmzh9muepp7FKreQ0czt6M+2PMUOBjXAgBvha7sHrLgD5YFrREyEzo/8z1nLJ
jcVbFcx+mmU8oZmy4wsnd+dXrN5ii9l0HTgtyigHMeMcS6KpBL0YdI2+sLqVSr0R
IjWxJwod9C+ukSPWLKrgNnUHD+/l4sJ0fMmlthJXdYG1d25Vv4luh/8MwBUGlqY/
U+uUcZg3D960BB3r1c0GVB42dxqVLPRauvJtMNMhu9t+tOkkBpSpTw6Jz3FzWFHI
aBdOUuzzycOzzhWjI9RADt4o5l0Jc3t8nScSezuiYvvHAh0N4iZxviQz4YgaCMYb
/BLLzwrUjLjQ5etJ1lGHz6qMlhVxRhRGT3yG9SgTNEmKUpVZBqDg+KvGeznGRXBl
grRy945K+puLrNqpAPX1Z4ZEvttLMEHBGQCdAE27FLphuz6Oyxa8pjPcEHzkXwtq
CiOD0ycr8ZHs/E85d9ctotvneZ3WCHW/kdVQmi/JH9tQp/LA8nYw93m19By2BZmp
qvPSV1bkER1zSkNGMxV6AdtUCmuAhFNwn7+dWN9ZRAP9PnmYJ3wV02bp+XmIXs40
ttvuh9u9H2WAXeeAmzBgLhFG55Seujl52oYmhbnjHIMv7WtSgKD1tXXkq/Bc8bnG
DBv5Jk5dkIjA/reGAASl1PT/27x1biI1/9LwGX7a7dxNzPYxx8f2deuJwE9QePly
2rzodNfOzJL2vCSN+qXQI3xrOzG7QuczvwOG5OUWjsnE6ArMBOtGSzm0EmY6eklS
F+w3k5yttEkLtz6IIKY60Itha/Sa9HJ/WqCltHwaXrQw44R2XCiT8isWS+kpqygN
LBFsdsgJ6OhNia11AB4nHp6CJTnCBTEazucdUP1lKqpZP3PJ88QFnLhCVPF0k9m5
X4XgeG70H7dBc7Rmdiq3iOBBx7vQbqOoZUYGUEHL6LgSUAj2Uk801wcQ1hHR7XPC
O4h3BC6Xgj7CvfZ1Fvcp5OvIezLjkMWj0S5fakdNlNMJeOkYz7ydTsIo54OrY5rC
4iwPqROeoEYHv41EzBAnnAqXm7aJSGlrtE2FtW/WqsijEB49b5UgC75lXWPsQwQJ
81J7v05Tj6Z6dTLjr4tHD0rTWpshULsUBMc1AaK4cB8Tm3TU9taQeISP+9lIaVgE
hWFirdn2Iusiv5OTWPseNm7tVZJdv3l5U7Gh7lmYsw8cnB8pG8ijnxm3AZ+rFm13
k/GGgTWUX0uLPEpjK9Zr1tOrL8xcDy4tpfTI7SlpHVNpn6yjt1aFoKwbDXHASfAG
4QqxaUMs+MOOM6Lt1vIlpraurinOMVZUlp//PNoIGrlc24LGZFUNb97c8fN2JS/i
skzGK0jej8ypk4wr09C0pOGIuPirVspfbA2/KP+2WIro7iOxuFDkg4j7gIGK4BEJ
W94jA/TKBTN3h5CU3ltldbeUisDiyPVyDw6/3c70lH1ubbc5YE4yzLN+hd0In6kF
dJSV0zhlBDAQa5b/4Xgb7EfQRaqK20oOaYwt6wUJzvunUpfuy60kw4+Qne47IJAU
c50U4hQjbDyx4qi3KPuBOTpiePDupRRkVdk6X1/QzkPKee5nHH/z7xWX0iXZVl6+
wvTJ7iZ8dfp+zGMExpXQA/SJGgNufruoy3527BssFh0cHMJxbWyAcJHI7Q8WTux/
jE0JnU+r3YEvQ35X918V/X3VDNTGU3sJ4nxdNbd+2Bh5RNDEHamdVL79xUQlfndi
JS4BtY9JPgBNbhib2r7M8YwyM/9HK6KTXoxv1ELB/l5FWhMx/1+c91nzS7j6rgYH
RlN5BiXOEF3R7uFgf5C+7fmpcX96CActAkoTr7Z21JXlZIUk2PFk1KDUSpfhuIIg
b1g9D+NG+Nfr0tpYpWAm0XQ0dB7rwz/+ATofxQGgzV+rddO0N4p7rRfBdGC94Rf9
jk7OANzJB9762gbqOcSrXciV8dUfB+C+ttxQgW79lcknp5zVMq1xDb7ZMAJ2Cs5+
GfnljaKaTiortGvb6Tyt/RNwjLyceISfQyDGumXf5n8+kBM7eOAqTgn7YphlEK35
A2JLIdCBPPpI8QqkaPyHb0jn5kn04UPg/GkC2FN+HBnkAFYiWabSMz/s0wxGt92V
UOe2+RQse2AbFBA877re3DvZlnZkOZp0G5irLAyvpHwUpUwxXmMZrde6Y+MFXK/Y
m8K/OtSIr133GZdtqkAuJ33ipA32+Ioo6hceQE0oCh/VLw6sQ9QHrSyCkyE10eih
Iu7hE3vAZWnc4R64rRUN3v0uL2b9rO5CnaJP2dqhc0Eb9roK2edF+Oz2DjyPO3t3
Nb3hi2p2nFWumhAhIZuy6ekC9Bc4llE880PkjmaCZCSZsCutYKQYQxYFRJdDduBc
VAKzZW9lBR3DlRwyQBHZZk+FBXHYR5mEUQQ4T+T7n7/njuph2Cl3AErI+aMazwa9
53J4dhjw83drhivEgQQPrV+5CqaREvpSaTEmVBce8IGI4kr8m5ZVcGHtR7+n0WX8
PYHzIg5y0YitAVPCHBZrytI5pNsH8G+7OWWPEMOVBEU4lPdO4aMIG45GbFCVnU11
RBvbSjftvGbX5teh7xMBJ3hzGWCV4JSB5fWyd2OU04qsUwtKU85rpSn4ePYPYbH0
aLtdLPln5nfvTi7Kn1RCv6eIKfR8iv6sX1L61otUlWfbdI68AvGpz29Oc+ECJiPB
44PpaPnURCqFPIsN/6fJFEQN7mto1S6UyGzs4RvObn4wFvH7XM8lBZbcpRousMRK
CfncGcl2G8b302DLVHwD5NB5KAHVJyLEv6pZOwlDcnI=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
hESuvU1qO8mtDE9CNKI+cQpIasVSbMG406WDcqTCDTFN2NVXyFo5cqZGAFpSpYjO
Dsh+EyCvOkwWUd3HPQoRjtZISBanKsnQPhOgxnIJJv9zG0plGShFnEnRB9h6cm5A
Y/jwbIUQcVanrRmkS6thZL8GcPrJtKPSv+2rwuFw+Fk8kBHTBQHqYSTNpP5Co3rm
yO5NWEY7Y/98D+JfDEeK8zHLOl0rIoTOURgBqiA/7l2dbKH/iK1Z/0lzyCpjqRJO
lBDeWbx3iGIUtyIyBsDIH8X2m+/nZkhHdANU+Uik6bhwOmfJfu0/79wx5o8flCAe
JDYOkS+Mxnd79bkBumasTw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5360 )
`pragma protect data_block
MTaveO2y7CUcQGfdT5ivo5lkqGWoC4xiD3RQCMqQoAWhPxauUYb7OybYsdhi3vR+
1Z+YpRwGDa1bkW7fCixwdg/q+duGeTcqH8vpRz92f/7ZFNNoZEuA115RjDFeMgbz
rZS9pIvMT/lma2c9cETwN6mCYUeQiEgWSL6LTVPR8YmO12bMVp/+5cOIphxUrLQO
NPwAeddqmtcBbnlGq854CHxjVoUHmYncuTnDfdD3DOii+Xtx4Mg6A57VyPg+XBIS
PBodKGqx/pGINuh+Q+DlSV8j4dOpnvn7K1ppoFzPrMoIkpPm6ERGNfzpiiIMD/0J
+8BDrVKZNLxDCnFb4GmXXSVn3cgZflE1OwUQECrOMozpWn6xnzzJKr5PfD+2H9WT
acvc4fZAp1FIgWwMqQRXoeZPEysW//M5r2fCBc4ua5IedzPzZ1K5BscYOPH9MGKa
dCMkARsgTDwzUGQ34JrcISVq9YeVVVidD7vh2D0yNFDaHJp2sv8svcp0/Uih4vhW
6tJYnGQHH4AkW4g2p34vM5Vg8obYkoqO7ingyi5Y8Rh9NpxFP1doIbiwDcEmN/i7
MkiY8XkxPcW9Lpe73Lxx1RIw3Z3eeWgGAIDVjOrlTLqWy3ffOrUI+QPDaNDt+ZSX
CYT8Fz7OXfyVoYFxCp+HBi7fnF+xRKC3al1H6vme1VtAOdjxO2ZpgTK513izfpE+
PRprhbz8vvuBlvC8Obqar3+f07L6I/ovRcQ1s1c6ZBHzUAyTB5Ue7axA8IWB4lKt
EMTLR3D2zlxWdwLaIBeeX0g4lnh/eWhutnw4ui0FG1Qru57kD/IzpU4iLhtusEAl
L2tARuz9YImmsqlwXeyn04MUo+yu6d6Y+NNWqNtICDmmc3lirlY37721U9CGuDM0
agnQW2o+f9v/vUPl6GDJ1YJX//6clcEe3PoBh67zresU6PPQZrNhWmJd0JnMVpNO
gqr2hBBRX/egoYV7pWeoYnQtKZpxgZCLRku7GCc7/sGKRX2x9YTYM/Qc0Ex7rQtN
Imr1sMuOALiom2wb4fWbcsFnPDCBYzyDWjjKOdWqif0yDobgdtHMAWPCzn0yamLn
yJ9mSg3hbCZo3YZq8Tz1lr5SwcLGR74Bjbebi1gjvD+GPi+Q+lQokZEE4S/qXAjf
hUFAIFUG6SiqZvmKeOJO2pi7o2TWWReX74QWstkskD/iljl1+cCLB9AzBjpOpfu2
62/2pQfD/im2ZuXy1LeooFwbLT807UnGXKMndEDRNM/WB4j1PcYi9kk0TFkdyyw3
LRkEiM8cQQhwQowlAiK8BERIDO+/4iK4HzNr43F7Q3fhiia2Z27M82VUoIhcMOsQ
oBkLL4u2QdxVIuwAlA0GlEPz8KIeNan/Z20ZWxzRKgjDdtWMLnLlnvY/UEh+2KSo
KempVRCesfvWBoX2LhLNSFYrMgjhfDlk5VNKwzZehi8cJ4Ib3V1sc9qt1yFGv13c
7ZSdGRnYwxKc1218sRkoFBjqNexbu27Hk/ahTqlTX91LAnZDAe8/bblKzee2Yy2f
iu5VKgt3t4q3Kb6d2NPujM7jXMbx7tf7IEzVXb1idFLbbVOX49XrZevfkVRJVrEU
9ykZEdA4eJxrDdSEIeuaLGnjog/SborcTKFBx+95LG5xxprmjCTzezUOyHbtPmZv
8KlHGOrZaRmIb7dMekQkHjDtF5EOi5N5snR0tW33tZSgpp+gm0AfGHIEIUzZ2qZE
AYl2RHRkwnq1enoEZK3OgpbEAtuoJIkOVzdaZ0oZW/SiQiZ3yIxuPIc0vlB6SyRn
NlcJzkeZ7C1zKHgRcweTxk4dEJxbc9kfIxiRncwO00AsWdi2yV4BTTef84jrIOFR
dVoIaDvJSEZJC0D26uITEaWE2dHBtuqrMhsU2dpUX2Pblm1l3sh+BZfs7lhTJ+BK
fJru/g6JOGk2ZOlVN4lZdhHxJPE+1OHtyBWyiO4Q5SAAWsIvqa58CA/w1QBSFJ3Y
WUxX35Ni38ULa7+tLgCqIvdNhs11a76mwUEjRyDVPafvUc6aBhA7bcVnBP/4kSuj
nHkkKtD7G/l4GRE62y2cp00S39lCEcLef4LDDho6YiUHSgBabBZ/Wpkcdw4bzCED
wPN6obwcvKMTbBWf1fx4hNqFlULcLJOGR38NhpZ1gEPfDXNvCrMmo9zcYXRaMR6H
lBlZJM3VKWiKVf+W1PevqI+io+3wcBgyRbpg45/M5HhP3UIS7uWxSWIUPhTNJka/
SDj0SsCOJTNsfzC0jqIATW+YFDEqcMxAfnhl/O1/aPRBlov+Rz5gK5tk212Bj1WE
ByKip5P9s3ga5EE8jZesPh2Ve/4HsOXlawv1o+TyFFlh4M9RQaw+IoZgbW6ErXnx
uRh8VVdhPfb/bFu7jOtYi+ut6KlAcm7b9rnmjixaZ0Ru6XTSvXoK/eowXMoqBt7S
5/ybgC5xMhejA89vy79jU8pSoaYhEr0iuIHrM6eIYoZkftflA88AOzpoqdFkwhLs
6phyGUeMtEi4KRWVmNinASzgNzXFoqS1UAFChHzfIfJ6IHga4d9h4l2NY6zjbAJH
/saIV++ZCRwXpKj/9pn7jaBzCUswOGzMQpcTGDUQbx+z6VKMKjo6bL0+UnbygANQ
B9BAIcU4Eh4zwvJBh+QnlanM2hKGqlGkKXrs03F0/jTLJH36hHGDz02Zra0R225p
8Z2H9pceNdCq5pAUHybh9gjqfa6jW/OuYoYd0gr2wlrd9tfc0YcJkEGSDT0Fb+ny
7FItbGva/6tzZmwhRn0a2bScVNfDsETq4U/jRBgH4CgAawbyi8yxgQUZKEH+V5LE
ElFgv2PHmilitK5SghAPCEjTJ9nFC7IqzvQJVeSLVkl3oTlvSrunLi15zOUlwhw7
rotC3JMajSYGnUtZ77wYmM0j3QQwVMwSLzOCM4EkuDM9NVattuf+FbYsXHWEjcN/
nZ5+lSASFA9M+GCTP+2CGxd0Dnrl5vpuKQ6M4ZS89BsgDukhzsf9egKsPR2ALn+K
XDy1sGvAtQEuG5Pn+tndKbheqXDt2GlLm0ByIxlzmvJ0JN5l3U2g3NgGxG4rH3jF
qKWVX6PIR8BR1G2g99xdIyg6Lho4wBxo0Lf8giZbX1dYyUIYS1w46HRiD3/HSlih
rgSpuooG+mO6YZyK4RdwJMdb5cqnpfNCiJ1p5LsTxkDj4gM0tJp4JSkwjH+BFyEY
gzUgRTmqFYDL2q862/vl9kHyrPo/TZ2coH+XjWOrDSH/hMZyUyGVAnGRlRBt/Rf1
7MySO6NbymLW9llK9rDLtF/2ONNLsOnefYiHycUOo213/DfMNiR2VCFt95Ip7TRc
B1hpzLAR+2XP/G1CyvgxC9ZPHbAvZWJXIhy3mXuk5yh/uqXy2jaeH0v1aPmH+Qtb
9hVgth4MGY1YrWBdzTz2ED16oNrtiHKTA5R26jwuKZ6sqS4Mc8vrsUS8mRPGerL0
I3Oi+IyQgq2sCnLEhM8qnt+XDtfCAfHeQz5TwdNbEWUCfLnWf5BZiMeH6gKPLH5u
sxTmi6E3EgDbXX/m6tFw9vfZ6VwGqRNKojFl8bXzacuRw26Yvp1Zys2dz/83IAdz
MJ5m8LMuB1Al86VG8JDC/D6lv+uMbHZgKo/wP1Ccp2ZEOnbgL2nEATxJ2RBwIkvv
NRL7AvXBSfL5ful3JvyVRAxw3FwjFZrxzltrK/tf1+HLxcKG2aEK13Mul0TKNqPY
TOJjTGOMqkJ/k9tsXrg2l018OUlH80xV4yPYoO4uLVzIc7iZbqycGkGf06ZH0o7T
9LUXLb7J9MZ3h2QnU12kdsnzHeFycmH3wYSUchrgSiaX64d3bohwN4pMm8fT7G0g
sDn11MB0B3HuZWLuygfmY+jgfEl3cEA5cBzTA12ApMzHG7mhEuIgzoN/wNNxdgdU
cve0VrzgQZvIaxGv1huSHguS7+anHk5UPMgFzm1sWCZKugI73XYKcAzXtMltQntj
qWFF3CCGddPKV3RnpBMtqURYWsoAMbt7DE2Zg7GR8/YKwo4OZduFMoqAUG2ZMeIn
oMaiVernZTTkcUmavsoMDzvrecPPS9qcjIETZtUouIgJWe/i3nfacuJwZWtzf3lq
NO28ZkYTezTxKNtSBer4xY2FEQclvilpNrBzNDtvNMWPto0aomZIRPzp1DSuve+P
boC98JQjl3ze6rerbuvGvoKS0HEkViefV+UC2Nz+H+LSkEwarFJACNRFDYRVkSB3
GOXRPnVKV5p8vKAgOyikF5Nz/gi6V32WdeKG+78DfesZUY6/732tD+HdEphbydFl
QBaviDXp2v3YXIzbY8p4txrwSXwfvBDuYQRzXKooiJFRZ/B9IrYi7yYB+xiSUIzW
3WCiu2O0EuseOvnv75Cqmg8J6zAm/DhAkFqOAfM5/salzJD9xndIrKMFrNrrRwqr
GW0zob1GB6FARQQ78I4AQJQm1JFTV3JIAqRupq1pwoQG5QO4v2PYLlvwv2Dk/sFq
1K8ykoFDekAtLU2zJL+f/uW3m6uj1EfW0gMC+qbzpS+27oORQotwE0MvbMxnnPR7
WepKI9dlrNlc9OA0iqDKPDX7oRSecO8H6opx1wGIxPEQNmkVlhe/SacOE5ucD6TG
GOHbpxtAA4MasGIJwruQRtNLDVX7ErqfWxBQXerbBiENZj2vEuAdR+EPbYLipjBE
msoBYlEb3HMFRH0gmljppPrXqboS12Xl/5bsTo5l5y95AJro+gQ2qiAmbfiAswGE
vIpvclY9XiQSf/lPX9CU/Na78iNkeH0MERtk2obhOkSlh9e7lnDhpPtpJ4a4Qu63
Ib4X1s6bh21+m7M/cbvvEFd/qglep6zjKtYP+VVBFHVpf8IDknFJI65Nlv0Dbeb4
sEHTBGwdlzGJMqslQpDo1AY7T65YdYEG0uHCNzC2eXg4x1FJxscGvvZFMbiOCPZi
R+LiTSjqA9Qyr78liNB/WZOua6tAyGdZb6PFi8jEhGpmTPVlcAP95TOwykpQ+HsK
AiXUoz7QvWZS6RkLDWhI2XOHBg2jYu29m4GdzymycOuJ4AJYwZ2LNqKRlTeOg6fu
z2Qc+D2sqYWwhYchaIqFNaN1XQO18FCttldpkSBFLl7RAh8PljFzWE3cMzujhuEA
vAKa1DNZIVadlRCvT+D06lZRC5d2iiElPOk3wn8S7wPQ3rAeX00CLrdAWWBiZ7zS
DBcE8QYj1eSm/Y5qYOMjR5g1KIM3QZb7UxgtW8X4qcc5MmmU94gZcEEmz9jFgAsa
ONpQPmf2m8b+EFesOrzM3yxcPp/iQuVV+A9MKSVpl7t7YNWeoLdXqsIwAxrxmTFf
PffiTLKtRKySdpkssS7bY3HGnSazCCCPzqOifitefXZV2f4nzcf3OjXCrNIbKNu6
iaYB3NOpb6dyJit1vMG75cEUjuwQ3KFhGB3Wjx/tiqpIpxEBE+abdfdtEDevd+g0
4el1zDA2Hark/bg0L3SfkFWLLCuurNkjrc8TG77vAT+kKV62qZrfz6E4avZuNomn
9ZN/QEBFmr6ue0m21on2nIJQhbp3NupC089BXNYx1WSGvQdOnmKSGlXw7nhKWfkK
hC3R7ZKGuZ/6Qa/fhBMW59hmre29mcngnDG6D6WvJ5oJ7V8U60/yJcO3FFTUpG4C
VRFQWDVPzENGKC8949myR7NO9rdc8Vb5GIRNHa3/BKzGB//pjyX7FesXT0bq5tjJ
oIZe9D/frUvHeAgxmq4eVCaqo6BL83xjKF8pMXyDSm6S+xvxjWUSL6RR9Ckyc6jD
KFj6Wbc0EhQzOBFnoeuGMPMN6FMee/ENd2d0AXOdm52OOElJP6W9blCKx36tp4HK
w7+kAwb5LjNuSUrl1+6K1k2ibnsvsbIVIbuuvwhMn7CGyRRDd1RaZyDGCj8CtI2F
lAMzJQSBeTtW/wo8TBVufeK6PBU/ZwKdUrlDmLc+N0pwRqKh41PyM9wJpE9DJT++
EszZHCORIilGiolt65DD8BwtO4XN6G8yG5+HdnYRIw9d3xj3Rp4JTIWJmj12DP9s
BUKE436hlp0iVfJkF7Bk1cGk2o996RQmyz3Il/6Z4NauLlG6SLDYtYNQK0HWfdb3
kDO7LDGRVSa7vFcgW9mdYNGYuTIQW6vuMTU6+TzXFogM9LdY44FFtLhGQOKFTL4Q
IflSlCyXiCMZ+eko7gliFaLla78R7EY5zddwv8NIK+5NXiXJKKMctSTftCXGK3aJ
1y2YjhWIHunWQpgIbJL5vYilxj7qsD7mEElvB5nu74foWUyOwvYxfDHSkbd2piPI
Ox1+C3wLLmlwxLGNY1ZMRUwTZ5WxQ4CRbG3umGRrZTtGxx3iDgr+5SUSVrZ3y6i4
pEWXOGJWzNICgAgCsWbxVdVUJibwwLkf6NpzKpNXHZnbqPF4kLq6DwWLZlRaqUFJ
Y11sk25adxwFBGSqbIw70D4Es1gxMfCrJhPD4KMAufoMkzkCtJfS/9COfkV6XKJp
Kvxuz4EmjccWTJtHQITOC0UnPZ8Fxjs1K6RRwC0hKFdwFvP9CHVbX93/uU7BSApq
rW/FAt5LE7m9oBQrKycle6JNq3OpX7aWqepWN0TD7JrV3C1TK7SiSwA1dDFPnIvY
d8nQ+6atCFKEvyslVlWoFsJGDflCoIkc1b0ggGFALZzNA6SV+ELlKoGuk563zjne
9qhtfqvakwzeShUjI+7DObAEVxLnSYKaJN7Hh6axZAsa+7YihdDF3mWbAitWJncR
Q2L0J2xhJmI1wdwSBHxWs30zjNO9n9autwTUqYuBpRLkb/9HVAf9j3ui3Sg/7jfg
t4iFFF0ugDc+AMu0WbSIsajI4IiShBGmX0vt29/vzeFg4tUXJpzsqyVTdjW3l8rb
/4DKA60C5G0PoYp5ADlFybv7/C8eveDgluTJU8lfF5OIlhaMf44cKJIt2heB6yhK
vwUh3jOgsYdWk0LqybDWYKMAjeyc7w26BWmZcKo0igLc7X9FCANWC20Z60VMWu02
0Ct8z5NoWS3wNq6kz8XKCkD9nSV1F7vN4ceM4sOGpcRgdUMzVKUGSYjoW/18jkHX
koaDL5E2yvWOPX710019gBs1OGOJnY2OljJLeGeIMJ+qDi6V7q5cqMRoG+gMv3ls
JyMwiugj9dnmlrD6X8wAzaJdBCNG0dqeqN1bySIHMnw=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
cLpOa0CDA1SUjYBuFYG/XvWNbHuQvqKIve56/TKmBTF9HOQd4BeCmxjMKd9iKVw4
lvqfX1no6fGUpIpevU8AFQIsOs1NIKxtetqR0T1osBrU4B+TzD6akvlhEWqAlIgY
xoMXGEF3k+acwHss4bdjrhoiU/igBJDBvUMyKZi+HQXhxCkWxIDeORWMTTfkUApY
PjN1voQ3ajXn4Lh77dIsOkI4fxFm0p6UP47jbST0wWB40GPKRJQDSfD9tv4vKxI4
9W2/aeeGmsYCCD/CgA1UY8IHpCSobKZV26mVyte0mommYjKFU+w/jtWguryvZyDB
Png75BWTlCJNLwAlh3T+Qg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5904 )
`pragma protect data_block
d58+4XceYFZOAflTHkGMpnNcl3Z4H1q4wOYQVsDTJdA2X9KmPmWAZiy0M9KdHOVO
AE/kiBR8BXscr7CuGcf8bZ2h/A9zIDNFv9pfxSmN0I9NlBXEi/ntOwR/rvcq/H4M
6flR5afEW/BhnmbEaqEGvTY7wt5MgjabueD2wYQ2ZNqSOgIK+pcZFPbqGDjTHTOC
01QgP97FC7J+ZHnxEK5cIoTCtEzR1Bg+k2iOcaAcz9H+Psmg/lFrRCx0DHkttQGt
WLqdcSgZg/hjqjqGibtpTQfKX4gQC/5mxOwJljlLNGmIaWzuZGIS+8CCVxTyuXr5
DuN8CmwBdH0v3YqAgPMbERHyniBP7ccoJPQrEZl8cpKWGeHX6y+/z9+YfIicPuzb
WqZwkqkapeaOjIhb/xKXu2aR/a0a71t4ThE+Z0/IkabSvNohV9EaUvLiMqZCYuCB
jHDfK8+x67A5BIarUeL+TgDta+AWZuEtT3MBmktNgwHG3/uAnXaXL5piTNtJSUG+
1PRjCyTZDdWpfzsR6mkgkSOKuSvseZCXbK9WJ+JxMSZAkMI4NkJ1uv0Q2Sb2e+PL
vwABgjgz7unSsKnWW3tzQyiQTrTUM1TJEglfN2i96FukO/kqpSoRLDv0P1veLRfG
HBfRUXKP4EFx8xqYZ80Xg4uauqdVQlq6CYVbQ+hn/rFRklU4p2Fjonp1Z3JmK3KZ
xUu+BK68Zr4VfuL0rMI+Dlz6R1sHyl8R1wBNO3LR9HAGnau7W3aOxg0fe4nApO97
Rb3yMT/E4hErF9Cf4lC6UP3BsDcZj3tdTVmtbnsJ+61hYwDAv4DbZnxCJ9WtGnzx
0WKlcl+soELTKzOWY5odLVHvk3h/DcCueqMBcHZcViVxWd6IZJcDaKJFpeifQL2v
MincIz68Eqao9gG2I82Mp4ign3eLe70ij3WcIDAvk/V29O64GrqMcQraObU0a6cp
jqwkHNnex30NusIQAjYXUf/aDhVloD82g0ICTeVqdMSBEPKSEg4go5cMOxbs2Ie+
0jA8tILkqs2UkclFeMh3J/RWaX097gN8fX9MaMKzxHjyKWNwjKEBQT/uCZnYwtwJ
2yX2yUR2gTnV1Fk8YxsH+rYGXZBNM9LIZg1u2QHWlf9RmIY0fW4gKYolTNm7SqAp
njgn9uY49uKBgrwNRG2fdv3ZktYLT6a+oduh3B1BD5kWK5B0bgd60Y5Ve5YIaKPd
8jzbZKbap5Di/FWxFm8L1QSq/1ZayAAdNCF5SfKf8cmvhJtjJUSUqtt8AB9DmWqa
KwFzMN5/8pFjMl7i4Jhk9ZH2magGlZnx237KWiWIz7GPTm6Q+gdHHL3hlbrmByb3
BQUaYFuI46W9ojY9BN+8egEA70XF9utgQ1MOXegilDNQxFOPBDVkn65WO1rHHZJf
M+JXDiHxp5d8oCrQZaWRfY2heLsRdOpzzpaT9Gsfjo6yjklRR4EhGNTjaEPenHUe
MMutASOXgu2cBOwMe4WWT8lw1Q1AmfCZR1rSuTXftCTAz+facoSSMoFvqONfqNmA
+lInN1Cw5Hy67/FmGsGWWxGyLNZzJ59jgB4coyPZ5dDGfuvZVtdIM8r/D18npChd
z3jT3UPJLJuuZBOknRbqKpAvBYmHD5MIMRVOGB/vbj1a05HNA6ysxjRbAeNNtRGY
LTJwyNS3TG45K73krV9MrqoxHXlBzlOwOQt4V4J+ywGKmMYokXEt9KzJVrYlwjdW
UixaQj1fL9+QIxkfQ3K0srBaZlkuT7hL6q7ti/zOmo0d9v3CfR/4J2dh+YC6kaGN
Xvb2I9IJPmm4KHanyfqv+fOd4J0xIHBU4PivY/OaZxNVx4PkONeQ3Rv/WrO1zAtt
wqAjsV8H6XgJdJ/tDiP5mLZQ6VwjVOOK4k86w+y1iS2ccZl8HpKJn53hr9rEVYmu
EUbeCnuasSte4ghx5+SITQAJPCLnEqjYapEiSaWjiEEL9knjRlzh4jgolIImfX2o
R1oLCfzToS5mn+DTlWvyNRfWjeyorkQA8RSa5GWkXbn/YfbOpLYTAZWd8meOxzFZ
HUiMWKRIB7eiFU7uvgrC63nykQvElnNcOcJJcEnFUQIJ6YsnCZDYrL3yiEZWMufV
iAo0cYaR+I6aFn5fbD2drrUshR61O+Q4KtkorpeTlpFigA0Q+U1XV4NpBBNHLpxk
Bw7HKxDBxejDnD+TiKif186RyK2GiYZOLDf53wbsNUBbOql9NCIJklqsC5w3at1x
VrSfvuURkNEFgEbZbEWQ7ma+XbVxhmSH28Mwgx6OwMlm5qtJP4J/KFv5qCOkBfxX
/tAHByVPxorEXhaOiM52t6svxQUySQmNAdjhlfyf4HmKrnhljdEpSmcHTmBp1YZ8
7jKIAM9/Z5HVcuiyGEiYXIE08T2zq2hzB8p7fE83fF/mLj2PdHQtiOv+N4upYIkk
4Byc88PuO0rE8CY4ecdtM8af8XxbE4v1bLAr40E6b0tUT80+r7SEqxKlgmDbZ82x
FxiWRpuXfXu9GUCsxmBZJHolq0SyyEti8aBUFmQsT9ZV/chsYpr5evRA9m5TG46G
nr1daLGm1Z9G3VszR2yVg1Ez81QbfatUHdKQDh1w7PfMz43yFYmTFHrsxvjmnmdW
NTyYjUnkmel7VVKyQ3DT9B9EAnWKUDVpD9zpI6/ZLfFCQHTBtpptsDrxE5bzxGtn
g87f4v34XvJeVVE/IPgi0wVLfI3vCW8/+tuKii49A2kowXbrMdzQuPwr3sjitqG8
GRoHMT6TSA/OWQViQr6C6/yVYCSEzJ7cSnnaO+hFQ87PwW/HuZWP4x8VuONqFsJ1
pgLQ3frROwE0XjeQmHSC2qYKzv4MuRcR6ebKd8Kl2FgpWmuarkQTtAzO7omlE8oX
yXHtPZXUQDm0avjaLnnqViTg9pTY5BnIkIi2EtruJ7py6sk3AxXPO1jRtgtdq6hT
MeloPVoLyFAvujFHIYNjbxC8I6oKlZtxsUSd6iJyEeVgJhhF/xY/gYPCURS3cWtd
fUVluWFMhzv2lHs19OAnEaeUAygdF6aBBRkjqze4M/+AqdOg1Nksu1kx/fq1ek/e
tCSYfDEcQwDlVLnIM1Cl4GwG1m00+/7sSUsWN7cB8zGGjMN6BhNgVJVzu8YIcXAL
Q0THkKnYyW54tXnAfAqI73s9MCGdjvfC4XHfAgGCmIeGlFo/yfwTvihQhbje/MU5
eFv0rCAgqXxCj9Cji8D+ERgEbmL+Q9uh9umF1Ha9KuMJoKW0pSf2hAVCOKI/mE7q
zvrZtJiH/Higzch5H/We/S2KwOSLLcW4Vw21f94DykoP0AvyR2h1Fn40YONZ7LNw
d0wtMd2c6QSJFVfVEhIvCe23bHuXgAT9pi5N/eZoN5W6QKyuBIRMCdHGehFMWM8O
BHnWEa8MFZA1oA3Rssp0XQh1k2oa1d2X2fWblnyskej5USgrvIoAdZTdq8/3C413
z2mqYG8rp/nZobWjK0MtJRQPVM5W44HvWrJuMPqMNWh/y1UTqrrHDGFuHWgbgdRo
BjP1fZd30fygGcL5hfG2IJa59ypgEcc0C5sc5f1FfFYi0IAtlwZqx4XoqvcZpiEz
7QwymQtaKLOiFK8MvFCFf3+c+oFb4TS9wbnWYq2X/x9tqc1TTfs9/6jYrzQ5cXj+
9eLFj1rRgQd88RUoE8Ogso0zduWqJkfRvJrvFWzTlDbLnnA7eHC3iH3+hrWahrjU
NZdF9puvSgNP3psIO6Wd6YIP23RnNhne3wC4GDskdgyztSvg519V8EBkCmHiebsJ
TDUHI4fRqmRofoD3RqtF4EXRkoQgxrFJ6OnNCq8/qYn8vpfiL413/hIX6znT+x0n
VNacJnCfW1X5JrVcnwXJul+bzrutTwyxxcizX7cSC0VsIsUn4JghG4UbeI36PxSH
aUvWzPTc4kiMbI/pIxbkJ2Jk97R2xHjiz7SNaiAg8lZD0/Lz7P90Dse3EgEeZdlv
hTx3EAXK6WNmqguTPKDJvO4m0X+0j9S9ylDK2uUco6J8GFZJqTs2qFZBjixmp2yO
dpBzjpCAlL/xsYqsBmFtI6a7ZyarfX6bdBK3/CXnzw1lGzDeowbm7QtDzEhfDrJS
Umrj9k9on0wKUqpOaqJa2OYF4Ff4nO+8q/4LwCIcRPMov+HCtnNAFyODKeeTOgQr
E5rWcaqIPsg3ManOt4xfhXXDUmNS6oo/SyF+trzlsBSfvsdo+ZZrsdnbqLVXH9kA
Oairbd5Xhq2KHQxsA7U2WVoAVSo8j1knJAiyANFpi9cFRPMw/XEocI423ACcjIJt
tKPGXQLpnxTQvxyPxPMyj6Wb7AYIZnlQvsrpFKygkuqdp+t2pFpQpYfMmTssqRbu
1nAtoaFESsyS5wpnXcabjBiF1X+BhE85zY3/T31cwm+pMfiUVnpCqcKXphtTzfXe
Fe7I+N/ajZxF4laibK+AOE/HoVnWOVCI47gVMPl48OzZ1Dcnw8mAn1KXpDmD4mFQ
XBlshMJPpgxyhYpdU4KCapItbwgrxDF+ff0pg4f0pJWBDzH33npaymTo6UyxgJl+
0f9iFk/oCBNgmkP5DUTU4TGiCrjD22Jf8PUCo34UqsdzYu1ng3B77L7TEYJZXAM8
jMpi7LJh4Ik3Po+yodIavP8opSaK82D1xYEcxmVIBtwTkZIjdB18BMmYg9f91Skm
MONIjLnacje8wGBWqkyP/lfyF6zoRF3aYM41sadvVAdI1FKhlrBahWY2vVLHjjBF
7Sl4Lem8zNn4RGb5eFiVH/rWAa05puPlSZibHoUEYgZzDyN0P2cXQECMP70XhFPD
fSc/CfnVx+aicShzlwcV5tKi3SrIgjvjj9sLiidHBiqW4JiL4tnSW/KMsvqKAO8I
Zd8SC9Vh+sn+u6iyadSkRXTKAuY5bItTqXKJTBIuLcvbnJTJV4wWHKasfgoN/F7y
YTgo9iMd4tY6cY63pzwfIHwvNqFvqKjMlxpix4jEoRHxGd/wn/RCGFB5+quvLAzr
uc3gcu0H8J4Jr0ABlExQwdVSycw8GqzewpvKQ/0HuS8kMGl1veonHGwQBnRVU3ow
6NALi1QCcnWXtREEOUvIOFedAGJCgsndu03zClBcb7epvqNAJhlSJjr2bC7cP4PY
/KP8ttAgyHlHBHregssOCrzMCCbYeAZRjwIhiPp+84p5Qt10cm7RIYaudwhyeZR3
CNtqpPKJ/8sUZkvav74GQBgHuHJ76qsfVqJ2x6z0/2/Nx9DgxndCVgRbedv9xyiY
Kg+Yr1YgNov4YL8oJwo13QwGNu9IxnJz+MbYFA3LQMlvk+jcu6TzYH678WZnxK2S
/MMFvXlPDYzKmNnvQAX0nzBSwLxJ5qeT+4YepSJurxoiPoJ40Akp+K+ZdQb4q6Uv
PgFcCJBHkSi7Po+i+4Bb2YN6tUWEbUu2hY6NW5g95iTxpg1/dNe+Yd5yElW3TGyt
r3/IfqTOrEuJp/iu58KEuAa3bBLm5FVAnt5wLE9R2KKDGvhVLaFmO5LSoVyMRST5
CLeVG8xQbk2yd91ysTuM4jgIZXeIWXTsueDE3+BjRjuSG+QGP5WwUgjaXDTP1mgm
EnL/biHrlt/fpgj+7LWhRyaJOfnFiR9pQvKOmj1Jsr+BoT53ktSme+dW5lIsrbvd
vCZW8sds/sBMvdodognXaIqpaJX12s25lDumkC9Jcn2SvWkyxGNIKgFQcqNgZqNK
ux1D84L0ZBAYzHX5O6hc+fnpsMannCXBdUFoSzqTBMYJPY0LJ4ZAuVCdEdAWEPfX
Ycesbs/91tj01JDAWZiSRqD9cK7OUPbhRvkd834uEzc0VquMdZS2f3ajBLg5gZ63
gXETwm6UWsGm8loD60RgA/+Njl6Rkw7YS6D53YkxmpJV4WI+mldK/RclegVOY8AS
41Cv0a817yS1hb1M/vc7QCodq7mjk8RIIeM2sdZEGkmN+NQxg9OOi6e1zwqjr+L6
4uqX3TKO9XtbvG/G4A+BbtSLGZVUo2wslaI84OlULy+1y+ZAo3Me5y1OXlZv2D+g
ktNYto2+nSVIgoA+abgG195azKn5+dJao3+Kg7ejfn5R6W95HiEN8gEO2EI1NNg6
fJtUK9eUYYSRHQ59+o/y/XuK7sEl4d8L7aDuQN8jty6SWRgSqo8ef/Lt2CL37nQO
aqf0PyLnCqz1J+02VSwdYNLB41mgVZhFJe1MAbaJsJ2EN1zanUiYo4spDzfOfxKm
jyb6uuT6VvKRKF7JbqGa/Jp1ynmmT8hlPv+iD7T72LsVdnhUj/B/NLixNi1n3dld
coZqDsCjFXGNqfxhs1O+jAKVmwDG/7dfCrvrgplUebYlXvmWfBUBM5NE7ZssnSRw
AA86K/5cD1s1gsTma+xRAktXSapr8g/4Vwp/GW0gT8g1cECi1+zxFKt/ACfDm2py
wIGUUuJAu1Y7hPWWp1VVjaJ4z5kZ+NAiES4eEH9L1H7X1bl1hcCooZQYkuLV4OSW
iuoIGKqMoEjN8Vr4dE5TBOwY+/wvZ4k1dXvTsI6Onz4E4urZiQ7myBYTPEyWjSFO
xtCTg4OzSDneLxopFwDmFtVgLFEPGxVlubAgdtmUDoc+GVLaHKLv6w6uT9ijsEE/
YaFxjM9e6L7ih2Q3lf+CEuzUoKbxfjO9IT++ik0QGRgXw6WCixYrWPKH5RM1qKvf
Uj8pR+vkv5nSwI8rxfRIn7V93G4xop5QgqpAXhBcTnGavY+puKsjKwCV03IOHqga
qD6K2h4TNeKh//21yi3HRUZLv5c/u8pSSjsHt04yYjfIcIvLPfo4qOTHV4zzmR9q
qhDcbbe4WF0fabmocQ+7bXTioYlULACUd8Dgpe6gLsPyRV5G+AiCUuoE1YfTzWUC
mABjH817NTC8FLEMeytOEUMPtZ9HIT4AwGQ59EB/TQpgyVktuPokfuDXZIESL+Xf
973U13IK3aXKVKgcRWYX2LRMZwd1zda/rmcpHDlOew9f7meJuJxN+dqyggXGQSWJ
Jc0f8p50J73axrr3oUSvPxTs5pqpnKX9cU7ayS1IlZYvpnZztNMA/gSlCmi+/KxO
cKCZSo0CiCw2DUjBfyyCQV0m3UooEgciUJrbn7sM+ot00RThtxCyf+mstgAoDj6c
u03umdy/C6aAfeb4npkkI+GcTc3gGoL++cO8LB9PVgjDL3/YdsxD4N9iFHcUXt2e
qlrGQnukXwZ8nMw7ZBS0ZLv8Ms1YBuKL93K0kdvy9Q8u2w+vLiW5ElJQ3exW/KwG
7w5zuSdzNd2lDpvCDC9I3r38LKsIiqZ3E9baCSMRFNZcC8kLNzQVigcnsq9xlNtT
oacZP5ejHy79KTp/rTexAKUh3sg8pTCnGR25eJpdLUXIgluIA/UHyiSvVWuht0Tq
qMggWHYZvL/gurLze+dBMSL7AVNh5vCfHsWRQ5j8ZPDUEKcsj7YVhrggKGwMFkWc
hZ9sViyl3KwlO1uIyxAOgb2HfyTi48HqQpVU97lPOi+aXuKisRSubF2G0BMdQHkG
LzYOyUznpd3ZT28w40jGieT+5q/RKrrY47i7NTPaIilgmKEM6R0wYWUPr1u6wJiT
2gyPBXJ6hc18pURGE6Sq7kAxYybSn96r6co2Gz+Kn5ZAy0kpjKRUgw9pSVduC3A2
ynZArPr4He+5d3qLTw0jg9dawIpN7A1O0wFgz59H/3RtEMnSu2OC88OiV9/nsiZK
s9e8Ysq0yw9G9L7hqM39xX1Oq3/B3M+5Jc3VIHKoRUd3FvSUC8eVOZP/XNpyxz7c
hbjb2VaYiCXrz05F0R3XKYCPqRKm8NDt860Zr2YxpOxs7ZkerePzfGljI9j0EnWK
6usb/lCpkVIoQjv+B3Bxkl92FBxfQCIpSn+ls5fBONaP+z43Ap0vuLslENXd7vzN
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JPwSMRjLkTAK6M6G1H8Y5A2YkAyIqXU4aFn9T8QFADnto9zW8CsZw1CxMMUh4PZc
Lb8SrQt/flMX23ja50eZTBxY/I0G+eJBzBRJoKx1rN6dsXlLKlNqCvDvUNlWkk1G
LrIiXuu0RDFpcPLpDKDbRmNqWsYVgQ2n/HwBjb23dvxS20bIZAYY9Kb6tjbil6Vu
mTJ4abjgyzZdmOSGAd5uPiNwKCW9SrhCeM6tlpIe8lGUxH6nTLivSSz4r3adlPud
Z2qjYUVONTkX6bSbSV4pirBXVnP65bMtbFVIKLbFfXXgrwC8iFrZmNcmBPqFeMlJ
Acr3heOrdQconFjl6rZsdg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7648 )
`pragma protect data_block
l/EtE2ZoXv1tClhpUB0nUnRBxz/NJa/d2YVi4Bue5q4tbabD12lvtdP6P8CdLBur
nXPs1tMwATOXYT0Kk5M/PECGwuI6XI5tI88cvQYhSg5tYRVYaY2GOfrJyzFiLQr8
ldbGJfxzl2w9NHByXsMXMv9QV5S/4kp4YA1kwwm1nbBarenoeFjbcbAi+GdFAiGS
3Pzp4Flg40c2dl2eSQlSGhQ/623U3T4hUUwum+TlpGKGnLxLS1YYCWzJCJSSABsi
yDI6QiJXSvmfST+WjN/dyXJAI9eKH9Lvl0xytL21n5QiOzMRG36UW5NeN39H3Hop
Vf7QrPy9AhJiuBVDrbgrhh4E09JC3MxQgISZzrX2jNwqeUaAX5k+VMMVKM78rliX
femG/gb2ZRGDLPyx7W4cgb1Z/JeCgqVj3+J8Ol++Enr1VzVRN/Cv2k6hUI4aMXlu
bnWaVxGcDLSIO3fPkR1TZdPcqMjtSH2/ZDYfZ0h+4d2X/qfo/6j0qEOA2y8kPTP8
DFeOCgL8i9NjsvG3tVKNrS5QSIllO1qcDzsVH0GCu/5R1BzYGHgm0TSwt3KB5LRX
eA25/qiXdy+k81JDoG/980LSOlG0QdZj1tOVx+XILvKi6SB1oEw0uoGhHNuVQMiy
FemiCZFfDk0tRl6jOHNLOSGxoe1ALD+AjMUuu67vu3Zhv9Dd78qQymHmTE3q8oZz
nnX8/v7BGHmlpsGQsn8QzoG0bwzPQuKYxr3AID8LF54yEd98j0CeBrhKHd+Xyh+N
uM8nZ6+/DRkckCKqT2/pKJllxfXgTo5+p3ajhOdLNDjgOMOTmatB7LWdwqQW5f0G
XCmllBOU5atApA8/YJJWau8fasYGgv1RjCkTFPvVL+EIfQbjP7GSDCZRO0o6tCMO
6K+V17uspj8E4b4/ILzpuGkSF+9gd3GXCnYZric0wR7Jk2bIX+T3WzuMSsWtW/Si
ALjM1oBz/dUSe5FUygCEN6+DKOTCvmecnMxMkKbWKwkc2APv5ymoAIMAfXm2VYS9
BQTXp5GCUvIjVsSiYiK6wvVhB6dFs4SHnf6WEO1jqKwHrmjzi76uBr0VzwLbRXaD
AS/JP0lzkmehAAxzXRNIIeMgbxD250CwWQX9aiTdiPB5qMgsrXocLbwgbUPni6r8
0Diu57lJS2dtZCciRigcLxoGHib4dgNnodltNQjzgRdc/4xRM3IiJgx9lmFQvTr8
fuy0oe6jyuoPXj1rHNymadSPGSh7tTiXdm6EnaOu3ltjzqbSHYrOMKRH6kg3BNEA
Loz5eoAGn8zmb+/BPa9Kmc+VwIj4roB5UkKl9QyCD5ctw0ZZkyxnu+q/Ml1o3R41
lg32KXoNIhZU+KeqkgoVe5/mWJ/QK00E5yMQSQTfEJx877PoJXGzCGCthYzcJpKw
edNITnmCVUtLkprXcxc0x47kaBxMcPEy7PB4/mz0KxK0NPeRqSxFWtSwwK85Ahgk
T/d10rPPTwwJbDILS/1C/vaBQoytmk1OX9QwL8CC+iSobeOZWKEWFsTZbU57SUmN
iwiBWGMk5N0y567cQ6OrkN1GmLvnyPW8Vveoueu78R5PtdS6RJyCYIp7zy3QzLCE
YjeNPENzs7WN2pS+W9OQvJQshNtFT9WhjnKu8ZHDF/sC7cOcimt0Qi1AlyZ1P03Q
CdZpjR0L/3hgPGbvRPRs3s4+aJkSJVRy2nSe7S1srjX77z8Ied0K1xUMD6YYITYz
3ctuYg4BZ2rYufYmeM3OXWeSKYjn+Mg1uzO3eMUGVH8knWqiuobSwcSGpty4OmDg
7OiDIBgIsKy3pLPbJhJOjOpF7NauxH4a0L3UiH0l21KGLxmIxlYsRi6p2WaP4QRG
JoQPI7pMsu7vWi9LrIXnjQ8+ukbC5m23iL5dixAaXE9XeTr+C05S0amxibdpzCaH
DoVTY1hs/qqSvhSiNZefbXBUzl42m6pi31p5BXRQv+PogoDsFAvlsvoBUqv6h5Vo
C7qrK3U/5g98cgS7BhIO6ooV/wqZQGXeYQEc56vwS+YyUITwU6pOnx2u9kQqz5C4
rxvZST2mL07P6JcXjirw0JEBHqPxERSQtQm5cr+xyaTswUi5DoKxwhUswuB7Crdk
Z9rePyr3JHqKA1vEM4DhgTu6+vQqqJeYj0FGf2Grv+SLAqaC2EeRAHUrjqMZjoWr
xoptULV0f+1gsAo3oOh4lgeFxytnwUvb/BGQZJqPLYR3nOB+t7kbUFuUD4N/6bEk
C5tbxj30jGv6b+gwAxep3rR4mEiEX41Ipjgs4j/WWFPfTyTY9eNVFprTvJFf55Be
KOZMxat/32dOlg0HFTbnJGfdPB6GeiN89A0PqY/DzH4MTfxb1oskVbh5RAOq1eMy
pVruqjgytRxgJL+iUwx1t+gSueIaJbbf189P3RbnrxxdbyTQPGvMV+EW/DIaRGf7
1eG6Y+94RNTFDnJSTFHxKg2yOWPkJbsDYwV2CisyQW6YxyMhKfO7cnYHNFtKfcKc
aW0sf/Ls1EIZuBhGJtt2jJ0H44i43HiLrP7iYDv+VY/JeDk5+CIEkOq6sOepfZoS
bxX4yCLiKxD8hUkXy9cXnb15+1BTT9wDh8Y+JmJ7Af+x9ap/8DBoI2uQudz0mLBX
YcuvDKldbssHWQPP3ktDRGCQ3RnKmdonXkI4zB1wCuna2EZeXmLKmQ5G54MVtRvb
PuKzr715rSKvdWEidug8/MZZnrA5wb8+hZo63sEOviGM8XQzuiPJb6K2uV8wetIS
xiGZ2VzihJX1YYGbFfRSddK/OseHR235yXDyNwE3Fe5n2UywFT8SsmoB4rtmwsj5
rKMnNzC5Vd1md02JxBEFtVAkTbqfOua4G0Ggomz2qCbx46tLbrD1jl+qFHnrsSQp
cFaTWmZqRT5RtLuYPSS0zlw3uueKFo3WlGSlwinhRr4pWsn18QNu+rHd0KlesFP2
Hht8ZMDlLButqDA0cUG2Epk42cXAwUI+8TAkoZkTtev59a+hfUFLPT9Ex6t2aEcQ
of2ozwB0bnLseFfdPArhJq/dzMQiPRFzuY6Y0FTqZjG2pSN4elDg9fr2l7ZiI5GU
H/zozHIFF6GYSJz06XOXV2WUUg8nojLmfGcqGuxd802CHOBm1uSOoQLJg2xdNPf3
bkZ/+HHPgBgRd6n9pbI5zK/9Y+tkycCI5izPZi3BzwC4PEdfv4PCKDVdQEFVeEz+
4NJSjJskU0h0fmCqkk809bYXgaEtx486wBzRAs27YFPe4KhIC+El2UE51k1oRzPN
6Mfw3r6YICLUnkG0jjVvZ4xoRbkmqwVNhEvKPKdto6ymtt904A2d6Nqs6eVxgnv+
4gnsEgxwzOCMvEgzGz/0JW5fKKZB01sJgJ5cRa2BdBBG/UQ9RJzFpX3xUgn3j5gw
lxBPM02HPDVMgFdCevSqFpHIWQYiYpf/wqLSMekcINA+dsw+3hTucPMBipxgprQ0
lCz30QkZjU3+yB9j5xXbMC4kyXtPOgQTYNiDYCsd5h4eE8KzTN4PqvceFDCNYv7K
H+t8UquoWMqKY3FpL7Qc7fC35pAgwX6zWWu6RahP/eZrVQ2BajOakt+BU7PETpar
RDJ5j5gq8mXMgenpteZEE0D9woQxsrIIgNQYlL1nEajOabBMVuQfs1NHOFOOA2nB
bv39LA2BOInrDazAQDsQI+uEd/icU06U3FIBk1gRDjX57N88sp+dDFQ/S2AvIb0C
hxPQSuyHhghrtw3tuLHbgUqolypXEUMn5R1t9cN2vqEJcz3ICnNXgPs6Sb9L6K7G
1pKO8srxxwdN0TOfgaEJwj6TH0R5OqLk1SwpGdrNfprMQk26mbuhK8n4EDo9eOXk
tCFu5rOci7+wvgDEW/Zr5dTpvB/E+3KlnhL2pZqrl854EYElKf/Nn3rJ/5mG6gOy
vXMKAX5sunDSmIMIvWzWbxV0Da41bkRIqAK1kkhaMKU+SJqetubY8f3ubsZMRxRR
DniJApiVKqhWPX+9uCX1ej+lwhKHtdhZ4JKe9Fb4VIbe5eGr94ekh1pkOpds0xFN
khYhP0gkRtaBkKvR5t8vsqa6yPixIrKZ9llKlZkWm5SdpTjXycMGeByghoUmNUdz
adA5QZi12SD/5cok2b2eYBqfSOLRxod2AHHf9dJ29EQkElE3tTtAKQ4anTpAQ4nt
yevAwqw+1dKz2Lx396D7sPftUVo2dP9N8stqMBrtfeIhancASAVMBCexcqDxrsrA
Dk23djDNnLoAQukw0Rim2kq+k8UFGMxM/QOrIc3HXi/BHvjlWcMmxGwuIqjlZSJe
N4znsbSRZVRtrt5UhYcN3+IlFG9PkBgMW+Y8+XWjof1zh/juAkuf0gQETk8SsOmB
TmMdriU1o3hesty31WvKp4sMl2Alsx3BueAWL2ASrcCL2khBnqlKAEl+vqx8GjKI
nmH4CsL24F3UL/EF4C5j2TQTNY7RRUtYi2Pcp6VGXYNoI1mUW1FjS0VC2rCYu83E
OzI6lH/+GF8uY0Y43z1OlcGMCF4w8wQOXHSQByyjA0xZ3EaAWgqXmGbZOT8QorUM
+0zm1ppMUpxkr6hbiZoPVh02JVJM1i8bcWJOYvFHga+e+0jeRaK15fCJoUsodZX7
EYsVc8xSh+ZI0vjxguAe39+7TPBzsps2XKoiJQ++8BBTDae8QbRAe9/na5/MZ/Kn
f3vEV4daXEiINIcHPghCu+EAaFjCrk0NLeeCcfaYk3poJyi0kEuDasRrfhwIbefr
A41xIcaEK4VUt5v+gLtWS/Nmop/xrXTzjcduLub9CFcN1zEj5jzwlXBNT570THVN
R9vL56m1Hu6B4D4QJqaYx/ORGyXpBb3Z6nlDB/KACBc2JfxpadVo+nggdo4/g0JQ
G56vsD5v+C+JkpEIBLcZmc+5zXYV16/NeC+L3s5kfdOyHXL4MJQv1VJHojgCbz11
uiGCX2H6RNXHajLLUoo+rz7G8d8quj0ZwlluM1x03MD+nwaSWUIiSeglLW3luBRL
TlmLgUv9klMZrUyfcouD2dkAZSGk2XIc6t7eoB//aPIwUb4GkNMcpwgFZF2vEA4J
SAvF0Ev0k+mquVE/TTPjojhG1Yq/Wf7y+4wqM810Juy9q1HLEfdsHJaiXBVSbweQ
8UaSiDr7jRQebpi7JPKAxZjJDA/SdsokCoPfV1cz6GZd65qOVKTumSaaqYxDbDcm
Xf0k4MZbDYnbQabCL485Hsj0YLlWgRpmSXx7lSlWFpm28iPup75zpTQSNvS9XPTR
RorRVgZ4ASTetpDAWIsAL4SXyxYQOsOT+OBcnYQstC+6qPlWmnK6+zfaxdSSJ5D4
GBFRSF6FZxebcLU525PPDNzXNl+82ZydDRs+dan6WnJ5iqUNuhB1MmYE4YUCfFbO
lYw7xES8IzVbcQ+HN0UWb0dCtbp1ZYXVSWv8nG6sQ33Y8oM1l1/Xmx5v5UgkRVNw
hjlgSxtzyriJcMffzF6RjN0r2D3Lba21Vb9wsUcFIqRtfZFPfEJ9Z8thky6onx9K
YqXB9zHiTHO6fA5huFDBlLNboIy2EJjcLZjG1TKbEkClJfRbyMgIRuZx93yxZqYT
nMXA0o4h62KEcNmTzQLxRd4P6X/caSNYTUxWy5v8utO5wzpjY9++xe/56Ue+9EXP
RBPB2adSHXiEi0HlVm3yKmhh/v6wYRJy1JtQFKov/MwuD+mhu1mbRl2q5zEUkn67
3CveIfRw8+UYzDi6zQoddvEcN3G05Q4y0yzfE30ORAZocnk1KXO3zduUe9UI+6jj
5WWvyJmqOycRU17cBnAPzraD9olUENkDW9nn8MgNsUjyb6Y6zdaGOzGswRtTbUaZ
+l7z22zLIJHvggLMGmkvSHBI9jpiVQWoxcs7UOG/NAn/42d+mSUMXCMs7vFC78Os
svdtmYxaRAfRHX9EI6nSY/yJ85XUS0/N4o0qKmRqBuC3I0kv/aKKwxA+EJkUBS2X
dL77xR4tN5TOSZv2im+4xIt5pAI6q3MJNoeAgiyAzEjWWns6sL7FsIXljSzZJoOI
hPF3qywt7jlWkdZoR5J4KK/9eQmmJPaJpGAk7vOC+Hp5iy6HjhHbLUeXkcRukYeV
V6BtpWoJs485x/9LIVMD3qtjrqPqnQyGbj2xkPs3ThNd4vdi5MbZfcw4qTwAxOzr
uxcwHqAJ35l9m4zbtwXuNT+WMcZdEEw+ax0cCHUp76NA0biabPkQkzcDZFIL05zT
BBQot/xF6O4IkGwJRI9ECVl+SGsHSjEd8VQlZg+B09PyzNG4SR5ypOzH3wLdiM5Y
wfKxL7U/bWUau3v3vMCZeNcWGA7Vu54pvfl0Xk95QfyuQS2WD3PQVs2nwCKESVCi
n0oARLJ47kPC2sBvvoeRmgNumOfodaJGdS21S3J/veifWIQOi8xNf2wrjqqQjoCf
MBY8/FvEKFXOjAHVyqE3hiAAqW9YTPoS01IqqaKJ/zyLMk/e6hUQt7vXWTXA64pN
igHUe82ybq5i/2GH1GAJ6TwQzXiOoWNco3SGP2BGSTadpGdJxhNO3kkuq43wjT8W
ye14SDRcpMiXotq0HUEgzJ4Rz8lJzj0jpn7tFEhHCtmhSQKU/hW2w2th2uOjxyQH
vZZjKaFSESORy1beuIZTv6lj1PftDzSH/RtvFx+KzDi07FhcDXeAarNCu6oZsQlJ
V1QSi0+JU21sfGu2qCOTPPguAUdiTjsyQ/pseGfcWRViok2a14PGtzGWvxQOZX7H
rEHMuHBVzVpMMcooBllGjQuUs5uQ79I/Fh5sRiqmtDBI9dTy+Oi35GkPttroMqpT
aas8cD0vo5j5V65rUBC2OLaipzHHJ5GYXJymN8RgSPDAxtFYlnQu2RNCXP4BS5B/
3dLbNhzjFn1IF0zPqt+XzQmvhq6apBJZDy1v6W+kJWxuGCDrEh7dv+ZApKNxDyIf
xTiaIbKB4pOdTAx2JoPkGfNZqPR+8bRYiMDLczBsYOC5gZK6oDYokwOHV5uawi2/
FN3AOSxe6KugblxULUsGQd5UlcQKIORpmch94jym3ZZYv6G26C0MV8RKQsMTzw41
CFZTgsVW5vJP4YZhinnuSlYUBWURN6iCZ3sBwgnN5x9pqzDyk6/3bT08lettuC+I
0+Wa813wvdr++wfT6qI5r4a9cI/RCxApO2SoY02z7cr6TXJZIvC4+JMzOh2hL/Df
/OyQEP5YF8sqoipk4rt7Xt8Enjko1LYcCmz7p/oD5n+dKLZctd8J4nyllxQNr3Hg
IVlT9PkC3S7d2//0d8R4M2f8KOnYyapb/2d7Bca4LlZ8802/lvSgjYKwhKTEMrv+
dDJSj3gMiOFzxQn6VMBfmhvC9DeUoCbPUBw+1f3aw94BCQlGfYlW9HSfJALBrOaM
BrEiu8n3gYSBQeH6HHzf1+VaiAbl6Vg7rkjxlV0XwNBv9LEYSFZDhsYmMZ0lJAdp
K3W9YHTRbYRlsgyhu9CIB8c8Mv5I2rYGKCeS9k0TT/w70i3kXOiHeXbhJh2IGpEL
vLO2xmQx3KYTpabZL9FLO5g2M1S4+otq4wPZgSZodN+P5UOoRChEVj/HfL/25XUX
hy8NZLRsU+d2iHPt+HhentyA+/yueasDl3D7mc/uY0Ef2W46oPBoncl/HnmoyZ+t
6YI4eFEt0cS8FfanqoLLNLEvNuCIBFfR+ZqRfxd+f3axLt6G2iPZ3BnsTISkyygz
6DolLUuZEj5GUpc49EuoT7+kD+wCTxzJAEBiCzqesZYu+2yNfjF4oOryGibNNQv8
qO7u5l80xROIu2bKLhVjoVMxyOSdYuXxmq2hkE7Q+TM0tTI4AbcXhUrt+d/cMCn9
p0QHWgptovU4cGIDS1QhWITC2FsvImMuFm4z899bhgWG5FLALWxODa3vgaSqQOYO
Z/17geHJoYidfBcCDgIdgO3jH//5E/vwE0pRNbfysXzruJN4BDY8xWxOGqGni+8j
8w0aX7pF37r5/2cEC3KtWK00Q66JT05ThmLhb9vXz31CxksGSl/iadplbQv9ToWT
GLRwUP2M8aMX6oR/Uyy/wYeXn9a9/f6MhEe0WaH0B4cWys7diQok3u79hfgV88Mg
SQWlxRloDtj5kTHNwvszOOX9jkSSmvwWS68t1vHMdf1R3SJAlEbdl3xCBizZV2+V
IKMpkdohRVlix7Ytv6Ajqm2WZQSgiOBOWLYRajvge4VWNc29+eem06srom5Lt8M7
caODqm9D3mcIBOPCVzA9gzAOyyyPOmw7iM5nKLjI+ms0wd8yZo5Kf/53Ih5NB4NT
9hNZTPEd0zhYITTqt+ubjjRhdIOna0Wfd8K4QTW41TtuDv9I+8VAcqMg1zOUX+ja
f32+hKXLu1pu6v5wuKJgdcixoLlDTIf57oI1KOGd0jyKMB20lyleYkehT9EDBii0
CnK5j/R+RouRoHxaFTMZD19Qfw1rkS2dOMnlbpafVQzUrQUuY0EwqFwBGnogGcLP
9hY+hQQ9nX6wTl1DfIOg9Np6R8FdV23Tm9vSHdTo9/bSMoWYM1Kd0S/ix2BCeofJ
PE/iMV4uiShkyJjOEeYjyHu+j61akh+SOinj2Gw4DjROEGpa6jy2klRUjMyyovud
YxB++snMFPc3LkUjr7jlTWq1u4JiKrPmArBVNv0GRz5JWE9mu7DlAh7BnuJLxU7D
z7oxZVJ8GjBuCL+B8pqVNpn4BLjdP1b7YVcaZAMVjhJVUE6a5TvpFClYFu7dp0h5
qVl+RzdOQVCwOmcXUvIsNsd7s8WxGUhOq0Y/rpmGQRA44F+FlRqclw5hBbMiOy2E
L/xeHAcOl+JMmGYXAC9YvvxU/9cDNYvp1MNOPQo/WJMAE54Ev+f24N/nnhoTSaqT
2IXIoyV/oXGea1+oZdHZUdlNZQ2ufcM1ct9GEUO4le71gNPRNnjxE2tIDqqoENL0
tcTAFcXECuwnzjHlT+caes0bzUj/eeoQPR64Aj2FOZO9+j37lcHilaH+FgA3UMoI
cNKwiJf3ZbmAO+MogfnDn7aBB77nyGtEUfqVTiTqgw369xcc0lGUQM/7dlwgAh8R
qQQQZ6zsdhDuDKyA+wjL/y3e49zTxIAEelAfpYVxdTyU8engih53NURgvLBpnR5N
yoskuYYfWmlyBY/GtdNOtVEcndojSGJsmT3JQx+QzF06MkPSfAXyg3WYdPx74cL/
uZ+NVgKqF13H+HH+kXrxoCU8xSQn/6yzGb3GrGs4LC4LA4eSz/mQO3C5j6pifwD+
aJdy0Ne93xz809ID3l+kXBPel8YvsXTqu86ZrK8b3pCSlTsmuNGHb9v0JldpB07R
Z8jSFvbTEvx9HVZ0LsIRlIGc8K6QiRxO5yXbvvuZUFPBpNC2XwxAb4uMvLuKVRrc
QIYBjU5I+OhfZws1zbTRHQa0cmVhHkolY+CNkHs3qp3RCBYAnVbA31q3eu25Tyz/
OX11QOs55FFr/TDv3zXyXILUbyHXDTn/y2xGPw5vqw4xGoSukj0kVy7b1oTLAd4J
HVbSuVfK+z5oxS3ff4EEjgKDxET8Ll57OrnaerorSMkmg90ZytxeIu/GniXEO9HM
YnJ0kCcEB1GTdsI1ZuC3OqQHrZ8eFRuQK4fv5cB2SqNv/W4uFHANHlOOIY525qnV
gHiw0lNiFyIU+YBhMcg21XUZnTnb+2fRyCD1BzbPQQMGEc1PmVqTDIz06/nfrz0k
nnAahqot8olnX9TclF2832hM/Lm84WnoaUbr4I4kSFs3UoARuBLnO+g2wc+f6O+u
mrypMCoR/cUXhevmkXnMIL37aBUnUpyoX7PobnA5r9kigQrhTF5+SVx1wsmpfMDR
x7T6Xishmlm6xqPYpDwSKg0vjl1z/gtVpwjh3/rYjmiYiP9ZtxdRTwOqrKI6IDhp
h9wq9VcHkgVmNp7z8fcrkpZ2n58+L1oGNj7z1EOjRwBMhFPqQcYjJleylFBvYXTs
MnqUXO4TvPAOSeJ7L+DAZkJX3/TkUkkQniNwbS9J9rn3sof8wZirji29K+9GX6yw
YYZfaUrqRIEcc/yqIdG9RZRjJ4l5gvnNo7qrYeE8C1ToKz/fJwKksaQ78GxjOSGA
SAuT7/5hZUkBtebaQPYmF9nGxH2HEUA1yYNKCaL21jEWA65T0D9oVqWQwlhCgu9j
3FEX8iZZYf0+FX5P452t+Q5sGU4Ij4U44XkwrOmdJqi3P8nWlo0x7KjKnjL3JFA5
J2MeM8VR5o3YAnz9SMiIgA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
C/TzgcVN9JcZHoTIC/KAIeZMaIm/4wk1pdM2u8CrutsSvZb/GrLDXkbYqfISCIhW
FMT7jo8h+90eRYcFud2jqnmgQKMDPrAv8e+i5/Ac7O0D5uBJLGDW2bIE3cie/ZmK
KEp5xemcyesikJ7gn8MD/b/zDdEY/ReLXSnLKkxf7JP7VpkVgFItojQmsRYzP5Tn
AUG8SU9ctsaXzpFmDOw9+iQ6Czl5jyYJgQ6iMIZtEmiRTm9kt+CdD2iv2kpRBRCG
sW0QeMRwYXBMfGqCxD3TDt3DbmGSSgNuCAPvgaVJk2HV13ttIrCOLlCS+zHi+3Kj
jbBQcd01wxyo7LwTfkFziw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5632 )
`pragma protect data_block
dtQDbmT+6IfYYnoCiyK1c6kfrxxRr53zqJ0DDjtZ3f5aXdrB6OKu7qIf45VRoYPE
nOFppqwvdHxEVqSskj8k4hX0cB3wtHTHT7WsK493TC4xGcBYeHwrnB0Prp3b0edg
ipMs4YqFmQCcck9so+DPmcak12ya0sBMA9+VSeFtCCzjw8EMMp3fN1PTbgNEc1cD
bjRi4YbI8TV1KkcVUpgL4EGC9Jg2LjE/tfEwzSggMfKbAyFF6uba+eAklHppVeVH
wbqi3FmtaSC47ot8rc261EIuE5Abl+XtCc7KAnB4tzGz26groexKkT/uLLL1gqph
59Hbyz8zZfW8MDQj0PjjhrYWjFF350NTygOnNL6AXQMYk6+2s4m2ExvO/1pFO0Ls
sXi1zG5nfuxJAI5MkcPojOa4/5X8Qt5o+k0RIOAfhNVzMjWXNhGz9dDHB5pRS1+Z
aaBR8jDEDhRqL1YgRVfg7j+eUTHG4XIwpi5Lo8h+oiWal6WA2iCqlYd6IvbsJkwM
7ub8+750br6GYvvEoiuQECea8qAoyp4BX0nc0NcnWVxnvJ9LWnEgwypd+v9qoNRW
sqjp/VvYVQG7740WATLG+rj8SX2QRYZ2IBvkkH7tf1N08hKDBDGAYytuJq5DXf7s
AuFzbeYpvjjAJYqMxvscPlL8ysKvaWwDW/rI0JYWmCPgAFHaxDgRDAvgTvvxadwk
x3Xu+wQiaSNoMBvAlSa/WNB0PhUzJ4fT+TbxHFjABFX4h68ALEW2fQmFtrLobOTA
dDtXMQIG/1hHNm58TAxRGd+sn3NLHKVvFmG1LiC1Jc+nKJSjDcMOOGEffP+GFbv+
plm/K61QyUx1vqn54uBpK5Q5RoSyNN6XrzD/IL+Z08sBGs7+CXr1Y+mHrl6buMrE
APEx9KlnGmWX3rURaGwxJYHAOb8K0xDWrgs78Cr7GNi2ytEnfsmoqPQbKEY9fR2P
6n2fr208vg19U6LRe+BS07+AQic5XFJlyHhAeIwT6pBsC8PIJKQmI+YjKMUUMm1s
p5r9Pc2g5ur1JRp+9B0YoHpTIS0i8zeQsJV+j9jJaQsfL8/DuUkQaaMMbK6PQUiz
qUiV1XiE1xPV+SJig5lji0lTCmMLVGiMsabIScMABirUjr5JvoWiLKDTXJpduRo0
ax17PmkAgFK+M7PmDoJIl+YVwsZLd2WZopxUMDdkT4jDjouSxtRlXysTaV21q2KE
blCpu40mlvAYyCdScGLezNjma2fujQmahrYUKf83Ujwww7KgKAYYg+eSXGFqBieg
weFcNkHKy69ww8lKuCywpsVeZEgKANmsFvpblLMrJbtf0ZQ2/6F+zhHy0ccKUBSi
1o72+cf0PQTJg+pEieMdi4/AfG92t1vsd4U1OGgFNrLgg5EDaHmzzYl8ZJ5GPDnJ
FVukR5etpW/0Y37dsMfBgkhbKSVZeAmh5DKOERzsBy1zTR0mPyUlvacQAVL3aocv
5GFfIRnVTJY2GgM79sHjI3urKu8JxNqifpplTydAD0r10GBoPbu2IGj7Y/UZa1kp
3nHYkOEi2waJRbJszRmZjAZ3gb70JKKaEK2AP31CkAe7cqe38fMn1hO9mcTJuTpp
0p+nOw17evwgtwf5sSFCRAdmjb+a47DsNNYwCCyqKEF0uE4UYeRnlBSflhAcirqK
MErhdJ7+Ve/fvebpJx/uRoW3iO4yaX1ZE2+CjZYBOPDjoOwUH7RyiUY5BiS36AgY
SVeEGmI+XaQkOLLF9V6oa7J+gkrJt7zW1fgEsXQJZ5Vx0yP7cmzhXjhAB3yDtms6
rY9kdmLOD6Vvpw3mL4Dtl+uznEhW1nQKrXEAn6VXGo5gpbSEV5XR2rpm20RXu4nv
EAU/QIV7rDJu4e3oKCfIo9Ve7wVvMp9s+DKcEZ8YRKp1RBExlNTetMH+E05BCxAk
cRrdRNqetJWw8nKZKE7rlWGcce6xIp/eQ2oRS4Xab9K96myxcoRBDHIk3Th7iqA1
cJCsaj8G63C37Gj+uQtmZpH8KPzRqeoun4no3RHm2DeC3bNQi89EifsyXmaiAmIo
lNOXdGYER1R2zSliv3GdSOPKOXJxua6yZd6PAcX1Tpwqlm1IEEgRBPn7OTB64BKV
JdAI/xT9b3YD31sekQts9qEW9Ttxgs8F4/UM+2JtTmU1GuJ0FZ/8m5TrYFPg2Ri7
zFBTqEvfzs6SaVx5r0tE3ZGp+tSyEg9RgByneq9Wjr5gw0jZSwGat9p5du57aJ4C
heyXU65OFctZL90LulvTR+6ebPa2+IKz9LgLORyM7OyPh4zfs7dC/7ZWK/gA0Qcc
+0BVW32mZrphOOaeWlCBVuDfoSqGgwSH9nB192UImqOthdJvDzW6C98f0axwS10H
0M+ClUbvS/Ol3Or61eH4efiSUtc0B9LVBFzV6RvspYY6Zxe7ZDV/Vv6SNPwSuIfj
q0ee67SYkuptyrKbADzUXQPe0y0w0qqmJ+9RiWFpBc5nUPkyEPrH5viN9sgrE6RC
o/MAE+6e93SxJLj65SfAjO0mniHbr081O2vcMnj348kRioaqxMx2OXis6xt9N/6B
eHTEXZYhr2xCu3Obc0HzgOmxPH7df3JKjbtuOVKL0UhXET1z0ZVKsr+z5UFTMJ1c
qLc2pHnOoKX1NVwThgawjkxNhAO59qkMKnZVVvZ4wCApf4ie5o3za365ISHh1oqQ
WQopD5y3vFwLayjZDrugxcHEcH3m+NYh++KZstkUrUI1s/eCft6uBzSwmsj+2yMy
SMuXxnzoxk11hoJUHNWRdv1Iusv81/wqCMCIf30oXb9NXMU+eOkibqsVi+h405SO
qLk9oDnbohXIxaWlPsJhbZgr+ALrPE2ZmPXXEohPaQ1gRhGCL3DPg3kCs7y8RxPL
GiV9Lx9EpRTCWCey+yEqteS/pz13fBVx2cZmqs2+iqd74REpzIYnhQZn6b/e9gOd
MpwXMnAFbx7zhI2Onkmft75r03TLPjqexMTcwa00M1+JPkjJGnnGkH/rIyRnWMRQ
HUR+EiwTdgkVc6vy43XVMEgpOqIIlh9o5wcRaVEsL3RgfoIY7EVede8eG7/ZryxC
76oRtd2jX1LOoQ0ZP33e5ZIJl5aDOsau4hP3mOf3Yi/aJvBdh4h2CFYd4z2Uezwj
m+yyQNE5HIuuEyE6gNs6Ze/7K+OhwF5yUiq5Ry1IsyqKLEnOKBEgpgzw7y+W/P5N
7oySB7h9J97y0lVtuQMztLunDOn9Rm/C2/KgUOnmoCpRy/NHRPyaNJ4DW95QKynM
cbLVL9hlA+CTkIPPXWBnCMLkY+TWu8dffpocmCzN0aDdfxEHP4uXUix2CCKhbux1
TakF3tP4VkOX4qceYMyjk/69NMsFFXDB78rVDyEVRlpzdpZL7JU3w+23K1GzwTLi
tHpxn3wlCISgzllkE+vXtMQ+9UA2ZBIqrImudyFSOaH2HioqL1DiY/sVXuf4mGHn
RRz0E1YeKz5zxRBdZRlijco4vmc6/2+JzHKbCg+aKPDherThaQKdnwlEx1Oy4JPv
WdvyFwC248qfEo1IQf3BrfV9Io+ZFusJVVpuUcFc27Vx02RZ4oDtBk/wdaXp26Oo
pvPIggnNrXJODQJCp0c32lBk4qSNG6FrvNRAroPSHkWYTjk1lTGyqHMZYemhyZ4X
TQ25nVQcWJGrhPBpyvE2LtAe6Ex6bib/MRkNtKSLWnEfIJYvuMNpfwuCFWP4AKie
eARIjJg1JLlhRoTwWMH3C+h+Cw22BJdlpJwYdiYnEUkK9uZL4YjhFZPZPwTtmOm9
ZJl/wqUH8Gz72RBP3pmr+jPAybXq66sDHADf/xITPYjDifKBAYIxrl23Bs2HQqte
c90MpXtQcf7PXRXBLLa7bJaLB7KOF8+nxx6kju2bv48QGdCyIPvMWDJlb0AHy2he
TdkelkWOzAIbaCMVzs1dm4rs4Wypfv0e3fX3Imp8RTKlImIC9dLI3GmKLixHaQyG
zSq1Vz39YCa1/RY3XcXUVaJuBVIP/1Marq+pD+0YPc9Laae/QGrB13HlclQtQSxX
wTdTdfEaj/Dqn9LQ03Ye/SxrEgWetF/0rnWCMRQsOmUoQ1NUn4qq/JQyIvAB9cPY
cIQ0PqQLE0D5gJgwneZCCo0QU6U9pRZnQOTeSIZG+Aae+5yJxhcUo1vUTTgVakKQ
xD+xHixXvQxbz2ZtnjvVhKTNpVs7t9Rf5mGTBO1+7jBJ8H2gzr5v+QTXalvQ4lf2
yaiVB80XC0HgkyeiqhadK8TxRucS65s+Bl/tUolMHVsQD4P7uxU0e+kx83dHlbRB
+1EukTwmF2rSfesM/S33sA5b07SSW05Diid1KMiz3fBQ0tzNFYttiQFxYc5j9e+y
iNgZCUgjVBHJyr0wHWXemOzCIbVIRhhsf2qYei1d0CsSlZWGG/udnMNUh6iuPs+N
fGTnvQUCaZlBtRh5giranMNhnlZ4Ez44ufKhc1oDQvqHu3JcYu11vhfXIiR06ufe
ZrbdWCkeDcDAIR2xy+tqhdnyeqYJoBLwtF2G+ywKc08jegRQ9n/vEqXucWBh5gcV
zQWgsmmPruCZLdd2A2QdSxRduzHHmzewlEBq5/9CMVgFuJwOwlVRRkC64H7CUydE
pKE+oR/QScN+ykmQd/SFs0IyCSEo+ES346hGdeoK0mc65Z18l9I/jI70PFdS+i43
CeqDRsxR3z+Lg0ioGs4HwBkB0GcrngESH6MR8HijN7aa/orqEGphEIC0VzKnduam
eg3ceBKk018NGEiouzQ0spGv9b1gPbcBfGHe0wzszZNsN7T1sk/4h8HWTCsSPf+U
wxo9jyLhrfAi17eJ9UwHKx2yzcK0qPB/6FmgGLom09aIQGRxp0OLnDL+UH5NUlJU
xX4xIp71TZKH+ddoP6LQfpvMeXjZSMP56JGx9XDaojv9+/Ph0E68uqQK7rh9PSpE
xgQn/s1abWfiJa4guKT5HrEHeXJTPOKHKdWeBykzJFXAF9Qg8oNzxTIsAAeHDJmk
iajHu6+dyP6iup5i/T4XNiYWoV8XkQpaimgoFnvhZB3gmdZc6I7yTzMpng4QONUg
36xK6BSAY1mMQuLO3YIWeZoflgo0Iorc/dYci/bWt0izd1KfeLPBmzi7nmI1/tSY
YLkc0jl86vYBFpszIV6w6zxorc2KrYXFoO01DyzyNQJZhNkgUBMkuBd7VqtD510D
ZuBPT0uoQuA8KdAWr+uNI8ssmb479hH0ckqrzf85MYJH//ESbNzOcB97G/C2TGf2
HgNRm0K++sLea4quSL01FsEG2+9WSd3ZTuSjYSZS40Iknx4Q5no81xdr10sYDm5U
s7C9fbDQC5sShW+SbOuwmtvVRcDSxE3cId1o2DntzbfIR51Wge28SQ/LP7pCvVrY
F5FLD/4x3hkEAjvFaskhbmJ1U2mm52AwNp0ApVpP/0Yd+JKqiksdS6adXI5QJCeN
HGxdebL2l9zt/Q7qlt92+nCigZob3l39alCpVDJ2rzMRmOCoyDDNUrRON5tz+J3K
RjjY2grudJJ3z1HO8e1CFXa9BMRVGZb2ESAsDNDQ0nfl+1THKXhWk7n0NmzufDJY
XBHlOTPJqpWzt8hWo6LX2jkGeKgOe8CAy7PdbCZIk+nD36RQnnij8o5ysNxzeD0E
QW3iIIiHp5GmdxbD9NHk5CLZV1PX/T7vx0RIZXlCxFyl6Yy+76rqPXzw5JXpwbde
fmp6lPwE6qHZbKumRgqPdgUaDbiB+ZRgl+twypuLvhJ3qoRJMG7k9+37n3be9vqX
tG8tRQYRfGlAzEMsmiKAqQpG79sDMPhXVj7mhiae/uJ2a/WcU3OHXJ16/XeJUr5q
ePG1iaFbZB5xAul8donBWBnvtIdxfrh3pUDYVcoTSGSBHE2bhYpePiVkasWLv3PQ
jyPiBFbPovMhoKAmXJ1ZuMaanUypfUOUztpBmKeLW6BjoXPCtWjbQz+lh9pMnaS8
ORRtvnihcnw2QfBG4H2KLzRcVan6aQJ6W4v0VbAdkBP7in0NCQANbZUMt34PurI0
EPKmMdrlbvg7G2Ln56ZHTO02FOAojAyNqygpSiL2GBVpn5vaQHylg3RBh2F5O5c1
XfN6h6H6WlZk+e3gdr6XjgSBciguKzXdX9bAIo0l1k5ndKiab74DEI+rZKchkzBO
Sk5jONVEmpfRGbmoNwiQg06WCLleo86IRc+kDXIvL9T80ttmuNxZfz2me6CRFDzQ
KqrT1Ci+8ylLOdI4M9qP/aJfVrBbjiM3seELzHXzI+wNa6CIPQRwgXwoJZShSGny
NIdL9wEe8glNsqnl11Qzqh67zl3DJws/cJPw1w+NS7DtSZb4bqVxGnB/A/qKNUZn
LW+1SsVVwn0dJC3gicR/RvgWi074GjWGyQ66BaW1EAqtrecE2chiflMT6FwTlT/b
i3/X4zWeUaXwdn0qIneHwIx7ZJ0w3boFnKIkMCw0CZGBdtmETVoSVabPnf4yZDLd
q3kXqULJ3CbbkneTqzIjkjoRBkTlCAH7G9KQ+FGJrljIJAZKoFe2PwV7P9jKiu7C
FjHxCV8HpvP+A/7/i+RORLvy+3w03Stk/dlT0EEOVL7CpUsZO5zhV+U0ZK2xBbv2
uugQcmwWDncQs1zsnxbhex+2sB3+ymE2dQdliEF96Fl90rU7/HSrpPmbJQLYTaBo
dUvO8NV9LYLduHwdc4auwCRY5TBZYlC2OJ3mneBHR4u+XrmdliqBUtUzRmFKYSfd
VWSB8eMVrb2AFsulfWnSlESDLZTHt11pEqJqbcUUSE8BKuTRHp3jkVIQkRLHcACO
NhSi6odjm47b+Wmbt6nsJ2s6JDH25PARaWwts+Qrn6g3SkshQ769IDBtLXVw5fSp
tsmlzOvz2vEBPPkWNqtuvXI+joThOcdfpzTDwbTxg9d4j0Xydv5GhGVDmc44JDL7
UmkXcVadLZjaqc9g73Gjicy8mqCIiQYx3QDz7VX264cX9Biuj6yemT9Z9y5mkyAS
V6YHQU+tg88X0/KVvRGT4YZYlLwKQY2kfZyS/cWzFCOqkekg0U1r3vFWcPQmr4TM
MJR7TrtfdsJ/IUni/wTg/JnexE1g/Gq3pwiWZ+5u6SBZyRzkWSSwzOvlGvKHR/V+
PSR6MJe2Ob7CQmJjzE9vm2xaWMhsCMH5/H08zpv1VJG4jare6iLVRUM4BJjSTpQg
/GW2CZ7w8A1b+MW9lV7qzLvgXCeBdhWhQdgvSYjfPS1jJ1naku4Ye7Tq+XLdly7L
vhs82R+3fZaVt2l5rtIeiuF4dCmQcVzSpnnlfrFfGB1yMgSjuPStCK/rm/UDEn6+
GCZjqQYxi3gkPidCIFSM800P5EUkfrQm4+lqXrRSj6XT0iv0Mq7LxCHCOl6KczSp
NRdJ52OCjvQkq1dY1MWrtiPls+VffkcBhI1lSbbl5c0aZkhv+7fypkzLHQsd6OMc
vJlqrYs4wkNZhrshMVUb9jEfIdagqhZxYijxeuNUYPLaIXniOixeSOQEaxDDB6dY
3yGWiWMXik/BgWRQUjeU1A==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
mxEfwbebC/UuHFBTFeNUTSTDU2R87LFhusc/S7WR98iXf/SxNai63l6s3vwx5ZsL
N9t5O+IPMDjIJEEGuw3amkjP2DRysX3ggG6mtyd303oIwQUAOtSQjd7Enb4xXBLX
3+Ram3hk5s6PodXxZi5SKMDX2nd25w89Edz9UCcwypSb4AMrxLYrzZ/1G7UC6kgD
dKHx/ohfBk1RFz+DJCzQPiiVunb6f6WCB0pyg7MrOVU4xEmG8ieIWXaRTpciLENw
gBg60WVwPAJSbLoF0hSaCNI05PkTd5+bbmMvL3l4BMRfEmmAXx8sh6kUzmYKqeDE
BtPmEBKE4mse+08VXCtzXw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4928 )
`pragma protect data_block
Ob7ILqq8k7yPu6c28jsBBYgfTsaYf8o9zSEZ1tyPM4WGt3+Aw+ulIdJuYC/0UtO+
vbKYnQPokcOB3RbFvLYP/7I1KqnIPrBedY89Z2c5eE9mKh06PYYjQWOF3z23VApo
pGDiPBOkmHWohARrcMM2ylkTFh6Q4vEsPoy0I36OOXIw/cQK9Y74Rxz3v6z3ASWO
8Kk0W/YZU1aj0nLQNVDOHCDKXv9PbPDNj8O3s8VncKqbOmr9UB97IyZema2sPFXn
gicR7Jm533nE1huOOQIn4ik53UNrhIz178R7SHWCBkusNr9x5ZDzKmjY0MGsooJQ
f1BzLmyDhitDniTuRPaeGQpHIzZ6/pCwg/6U1xJ8LhHwCWeLKa4HLp907MenDRTM
4Ic0Ywh1B4YbI5DrOfXfoPezJ9+TMc1Uqpc3POUjTWDBxZVOHtLJ8+ArsjeJAsGZ
wZFGr07kqriwDSyekd8yh2zJtw5JS72+22LD4zGBkqoEaQlHK94TOm+t2/cxNKOQ
SSqY6621Wq/BgC5XaLyoMyPWQjtP2sAJ5Dj5X26/ooK41H4ozS4BNVkV8uA/qnEs
N31rXBc/oG+ECHWzf/9lcXujXIzMjM0fzYTb1ydWsTRYUXkijcIscD99woQG3oId
gfuD2Z36BhkjobOOXxwuggK1ukPwvGIg0sGVsQjHmhg+kPLpyQtYcxA8epYTLDbU
uG40gYwmq7ntdSa48C4dMd7FyMsWimHy6a8fwZZImsThlQ4xdco5LnSjCDBX87/r
/+/I3wnSC/ZAClDUXEVassutyocpaaxsgW2naqMw40wkkXYfPxWVwLBp2mgYLLxL
89kG+qcohNccWQz6crYhvl57kRsIY84hqvTgS3j5pAm+fOJOF4Lc2X12T2WObnWr
5F3TpAV2epF2dTspRalL4hOHOHOQy70eGNdy9CIRV11s9zKe6ianiXX1hu4VZM+J
SLrsdFJ+XYEXDtGSpLFAex6s+IYf//D8W25Guo4HEMo8VUPKm6RHpAEJAD/lDOD/
tYz/UKdn2+1FdFtFIfPZfGoGfuqX0ey3zjTpIzPpshY/UAP3bQAiqWtqcYiyppZn
sk9U8s5kAuYaI54CS+iDY2vp2Voa45okbS05czQEnamd8uCoGmIFatsWKlr9fKDZ
ZqPLAg2hB8J/5YAXF13+DD6xfolYQsrI4Vedn2oF3vMXrY/1vmzV/J34Lf5wc80m
5cR8/kQq9T2hvOIi0WaA0hCkIVug8qhN1FNDAL09QVQwXVqOAVDrk/HLwOZRwO5W
X68L6J2qlVIhU/MYCs7t7Px7VfwfZzBiq+AILQOAcUZIg6q/1uG1QDUF6V3Pb4Ix
JXjAlPZNJVZGxm7X8OPXtG/ZQF+hzAtuncCxlMXiqy0qKoe5vP0qmZrad/UmBJ7b
CvGe6Ox+QcfEMfWPmpxOLpvrrIFU7aNPJxXVJZajvuOG6a8rZg9P4cXMmp7QmLWH
Gt9HnW6r5XYrlzsrZqNM/uyanBc/6CKRKn4LutqQJbbVOyO/tnhLgsMmusZfLEy+
e94gbMQKMIEqcxqUtdxzhGk9i5W2PvjkDUOQEZRkNPQFoFGyCPZlo45iO7MG2yfP
njMeyHPAMWyr3tzUx6ggp1ghbCUnqnElV2/IuUBD2+FTnIl+L/S1TTyaC6O1QYRL
kVO+SKrz4j83NnGVXZSGO7nb1pIy3u/dj6KL9CEtiAotXrjQ2luyGA8PQtsJTbjf
mGgCyZeAinJREtRCrN6WWz/eYK85NVj5rYYdtSCARtUizdDE5EmLArBsS4+HcnrY
MS+daGbnlmJXMLyrzpw0niccgWWHrykijj9d3o+tIUwVE2nEiadSaxUSLL+bXTAX
cBqgpzIFk4hzrtX7zS0+Ce9c6GL3CSwZHJSLW7OFXj2pqFZeVnQEEb/nK6qwFIsM
AiVxrpN5bMYu6HOxYM647A4YLkygg66OUmJiZnuEXo/qpYrnQAAgkH+vgUr2D5iL
63eosDVW2tW1BNEZnAbYWTSxQnEiC3ZfD1JhLlWg2+fmI6Stt7i9fdA6Fab8LBiq
VVHpPI8DdHUBAKi0n+4sUu1/Y/Z94INWnOvMUYwmwwmFgP5RCEij4AzivGC1WA27
7dG4jlylOWnghU7kNgleJJTMpElHPNSIEWsdiHgLcJvqLVntAY11+9l74r3iu71Z
Ycv7PvhV0yiZoTH1VQV9hlJs89TxmIe5hcZl3ul4HQcrFXOsqOjy0szud4ToB0rB
vf4l5kmNIrYPOmEA+pvxmLveXe1IUJa6iR8sd8PK6/BS7rhnXCENhop2ke2lqvjx
pwfXtaWvwkrAOrg+vUbLklYrWFNBey05NfFndgSz7yiuzMXWeLJqMUzpw+fICKX7
2O667OUupMpGacXEQW+8jKvLx0l8fp19okO/mOWbktMGEWdavHVqlTLNhZQWyF/Z
k718dIXybbonjVCIw21c3hdOfcog1UcINU7OVkvsSMGIEm/PVWuWKI7vW/hpSQGd
vR7PTn7Zckxa0mB5JYHXtZDyoMYs5wTsTToxojgTcyC4q10CRJIWnVJ5L3Wh2zd0
L8VvGUFRiO6MkDjn5+cOvM4E/VPJ6hsLW1OtZZOhxTQ9JktBeD9FX4qs0yXZvO8n
I6FuyWpDoDEYPl94cu1wJE4YD0oSQXSKg9payO977SAibnf6ab5rMOrwYkI8SdaW
+FrDsHt2Zswm32KlhfcVk0MRXpwzEECPQ7mG97nkvuaDtktmcpwpoCAlYRkEtQkF
TZJkxUtSPUZMcAqa/asKS5YXQy1DCXe5iMB35bT9ze5zksisfE+TRBG4GY8sFdYk
DqhX/Z7BQ9x9yiTAEZgMIPHSqURzLNqvVZ3S1GdpNF9a+TLUaAmyeY9jzVuCNa+f
F6fNGHPAXVY8DIR+lyncqR6MQeQHJ/YF9fl9uxT6MxXazpihsOJl2PXctUz+3eYa
e3KbW6XOHw5Ro8z33sBzCQBqqpjqvpnBiiQ07EM4ZmX2TsjYTizEYkV2lpTwNvOQ
hM9DUNoxaivDdFNzdY5PaAhaUGEdEHkrAQn+/grxTLtTMsVsTHL+EQuV8VpbBukK
1osUrc8BosQ/pbtF5pmbD7sjI62srTU4xtZgkHrA2Ji3jMSqpUehpLgYbmGqjS/K
cKRva6levNyvPy89GZfyZmNTvvlNYqjojdg6K80J7kSlDBAeh0dgeTGphoJgeSfu
IXST6cO8HlhYuWR1jRfB+Es/sMfboHMJHkayYgtzVXfpEKK4V0awd6I3BzKqVqOW
U4KnrABmJM6ukLyqD2mppX+fm3WO5Xtz3oTYjwRb3nA8mye2ok7JP1tWHSL7hldq
uq+oSivuxPtsaXlXdwhGO00L8ELYk0pZWUFT3D/fVa/4LetwLDn497HF/GcBCQuo
ADvUET8zoHJIMavd4zgEWIjPxomP7VaT9WBhLwPBysnCBgiR9eqpQGlHSvhNypPE
CpkPHwxHSMzi6pzEozbsjhZ7ArekcXV64pxozCvcMWJsYKuaLwRlKpALgUGnjPjN
1H2ljG2dE41zGeB1g1UycGr51cfRMHxKuXxjgQeMDObmOSD5zR58xsQyAhKWXu66
P81QJlNdb+kphECyRaXjh77Z1r4oKJHm4ZExla5TbzLMO/bvnSkEqQ7V8qvvKYgH
si8vjXL3qkkbRVVI5GHN6298FJNANQ7vpUwPCvqcXEg0bYqVjzInY5hSEdHzHJq5
xl7FRG5WGur1UpVM7JELOOGTZayRRmhZHk/D/yvRLXm3gg+wS/pm7qRU+12ZZk1D
UU7iVVUlyZvVIC8x4ola9cPISMduVvqR0rNG8KlhsdeAvGY30cmdDp/2/2IrSbsr
vNrRZdtRaifeXSnDCVyfbg9HhJLMkiC6DdeEpydxFJOnOHv8uhnBvxNKMbym61f4
jzOqbaKupI7c4LFvyb/m8r6bnx6zIY1cxlx9jPidukOv+aZ++tW/FyKGCqJF0zKW
4upgYfnhldCm0lLA7RHizViPuNQ17pZSksmy71ASbhDfymtCyLCHa6jPAIh4waVy
bW0su3yDKCqqktDNv3zPmAVI/PE3MlgmHCx02g7mBpLSD0SHoSTGiV0DfpzocLGE
s6pxgv6kfyCJRb8LBm5R2/r93g+mmUE4vI01KJxfxCBzoyCdKGiMMlPvvSHmVyKg
gbyQHaa1pn7Lq6uDDmNlDYFz8w1TIthh3CDVk0103m3n88afL7z0Ss0ppZmj42SP
cw5wLm0lmSqmM04X8y1ud7RGsQ9clNO6teKTcJMGISh+tkBweu13Ec9WOH7bg8nn
byCNE6GSagYTDxkg+tJUJvvNQWWbCXjmFKqFdMUXpZUZEYUolYbrJlcYJm5Avh4A
sRBjz7qGkbofVgl4CTN7NoqjE9dEVhSSztOoPki9/X1IAezXrX1nMEfRXcueT/0N
qnFfycn4AtdqUF+iQyt/Nh0gYO/G8JccGh1038OWoE3xeKWzV3gwxg1UvyZnLf32
PUx41d4WjR3QPeqj11FGJrgqH95bUB5LrDDAYTz4fDASH+2bizShzMcQ5ITOPr/k
55bS9a10AXNTBOmJLKysomZFhoJBjvlaRpuwWJLnFWrU+aAebH/ErTMxeLWCKP05
i00ucPu836vNPry3F4X0GVxAtnZj64Pjdhtq1Ua70aIrMSC1QDwW0nUhsOjk3Kn8
tqdaHmg7eUWDihQdgnrXBWE4gkLr9pSQCyl6sAov2k2YSZRagcQkIEumi/m3kioO
xruy3ugvVkdArngvpmGXl05Szx7U1Omlws10ctBpbQYtN77O5bp7/U0dIRLGhOKe
1RDwVikVJaElQFbYJljfPh1Gjf3xcJfxkNjQl79rDL6YwD0sOu8ikgD49qZsCyaD
5ZnuGRKRNE0MrKkaTFclJadch0o6ewQA8zKlPA2+v6Zmd4ln6w4j4+hIu3m/vj9p
jvx6hGDqG2gmT6etYdIsC21yccBnrr5DxrIimY8PU1+Fge3xjqzfvOQpyAlYviee
hQFqLj2sF1PEdGTrh2KhUkiNcMRcQqGiq47VaKBvbbOVxMj1l143Ev8m+4nPfNBM
UYjuoG1QgG2DwPvFFQsLXOeGBPp1xuEwWejuul14UJIxDLaMnRSqa//WyabOpisx
Je3v0p60QrJv59XSuW221oWkBnASPxnQBwoLj9Ci7QumH4e1xf/RWRX2THEdbclb
3ynt5xIt/fsxC8PBXpsnkaqdOK232GghYTlCDRyO8NuPZIAo5e40NdcVKy6a/h/n
Z61Q9CrTsGIkANssw9NtTSu9QEOULuBYbrNj6L53SEcN0Zlaza7R5yAtCHqLYwIa
wBb90Y0G1cIvGC59hVp2tri9DCt3W0/Fz6+JzojfFqAUkbUOoMU6fCnI3izgCCXK
obOMcD+wUUzLhobsSaYhG+lfU8qTL/NaWOHSjOg7QKwpFw/0x1JO6ahWkbu7nRAE
FnQAVMDnUTGcOgbnRg7M/x0OWiUzU21MeievzR9iR/1MK+KgS/F4lppUXGGMa1pq
VYAE7wewHoZdHuPX0+e1jYVI1HoRKsqQ/0R4X9BxTYjDEXHDin4ehjA8660j1SPw
BlMbDW0R2RN0SjhGd0RnBWN1ldGiucxwhgLekx0KsnBEfhTU6YKA5k0m8tBVwecW
lDLFwzbdHc3FFHyJdJr5bWMXf5b2MIUJI94RNdGRt0URG6LTjkC+6qVyLolmoNo1
4opxkzFVxGehfXUdfsb3h5tItArTLxfMP8iPMzYbnP17kga1J3zmsG81AR2+LvLN
GgqxPQ5ej/WHJFMIgHBmZydrdbpFEKmGeCoiin30P9YDx/xm8hjykUW5Lkd+noy1
2UI8DqrPWupaI1fl1GbDBOTLJQ03sngSVrb2JfobUn6MVjQTXDp+Zcm9pHSn4xos
NSAFqe49zYq5G/A5CJruaz+PwPM1Z6Q/vO3Cw4B0VmXHNksbZjKhoEmMaKXNeHjr
UvBoSatpZK45Jdb3ueyprz2IO0XyLJO+ERF2DifSVFy23WQB8V79Zylshku61qWb
vUrDrTtSfFUp1rW6/8i9P9/uTfl8y9zsQ46iLYdww1cXInFGIfLJDV0/KxJF/ciW
4DnjI9qPpT69/i+oalAOkDNxhZN0QdH3q7iD2C0OxtaYTmIwnlKZQIi9q9Wd8rQ4
YGdrO6bQcF2q+T/ADavR4N+QFplM8njVGYeznuSRqhlnC1XCYMjqFyP9abRbhOAC
DuJK0Wuj2FJLL7TJjnxIgIXrNirqJWwEcopbK+GbswLGh8QDAUxA88z5xgwMXCWo
Idnch1WP6sE1IZEYVbftWDS0pCp3NrcgaOfkUkebGT285vjjdY16WYjfoVBHjEA4
UC8NXPml020snch4kSXDl2x+hARBmkpyNwfGcfTNyBASyW8/nuStM2Qo0gLSYjlK
E7ib5KWeqN8kymOPzR2ZT7VPn4p2sZxELDEcLuMUpWah6ULqOkgU/3DV1dN/VsCp
r23USrNe6u/qCCd4GYldF++lxIFA2NEm9eynSxHOgUoYkZsf7WpDRtk3Ma/7Eds4
crseSb0NdXxMp20Ope9c5ZKxc8MjZPve1UCAzygjT9c=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
KWKtPjfvssg3a2pDdIpNIS0nRVMy9j9YoRKzTR3mEoVvK+8pOkr+snQKVSw9fUwt
47VuRM/etL9dLMWmzlEL86lN3S/WSDJTSsG22G8KQEbxMknGj7OEDWlpKxAqiPdP
pFUrGp9uHYdL/hAsr+esPL52ewXrG9jGf0kzaof0wGJdkmlTTwhlVB17kt8w5O2n
kR1oqsiGVosRIkxjU80xkSygzmr9F9Bea+sG2PMWAoFRjkCh63AuW0z+2ZHclMzd
17fWvk1oxbm9k57SmmHUGwUJpZmhSDWsCt2oHTdXC8mTWwQGCRKZ/4/dhQNRfCFO
trFvKInmDIsMSIUOgRPhvw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9792 )
`pragma protect data_block
OECQaf6GKG4ZUiwAjX58+SCwHfLUnv1Y50Zfm6MDTvNCzGRFdWMB/mYfv2zVanwH
lT8EwMLRZbZercRAiH/vP6SysJuv5AtQQ4DCJ7yXNORXgwn2fMHWaKjneKNSys+L
/w1+3a+VzD/2X+qC075fL5iTy/5xwGffoVQWRMFAgpqVfWqGDBEQ2INCn/TuFYjg
SqxiFGbfqwA5TjXnM7KM8t7/GE6XbNkOE+57eVKLhi5a/d4sehFCrGl6itlawUP1
IIWtKCxpYj99+GemIAFVIezbJwAlm5Asto/6gEWfX2nSCpHn1hFDWTfmlEpa0Qsu
Q7/qurDXSONZFq6I0vp1k8v5tgjK++WhDI1CeGWOgLV9Hg6sLDgcwi6cKbIkY3dt
En/oushJdvlx/nFdclZIfe9KDt2BtkdKml9JAZkl9HTLvSpDS4eeYQ/QlGT1CuSz
/2EvD0QqfIVfNXHaduRrmiQz4O0CUtY3QJ8W4FTRm7H3oScPX5lwVwvc05S3DgxF
5vHi+d7+DBXZIBd5gPXsXuE5QJg0DyqxMLYhUS5jfaUEjhB1XdU9wp0Wfx2tg8Jp
zTAHVZIoGALnmxzwDEE42w/257mOUAYOl2h5uIWnNQSWYxrwoTYXMPMzpyuRtDO7
C6szNziJZCDR7bsO28a8/WgFkiafCseDOgeovyFo83D45iMQStXy1+4TDECHpib+
3qagqOMGYJ51z4PGJd1xNrQezuJ2/QKzvzOWHaKCF1rju9JIaqflMur7erOLsUZ6
tirQK0aHMHEdemBGtz0Jr2oRspWT/38TE5YjSAlQw853jbEw6IlGYsvWoNGjz/PJ
PXwMyR8Vcu+ez5BQrBQTozn3RBTmu9r9InkSpNYL2FqVPxo/kmqcgsP5A61MnLC1
w7GQcJRi7Lx3st3MFtGcLA27wHxapdjUNpT9P5Hylcae/7YEM53OIVofGKJKYLBE
Bz2Z15YVUqPle3Gqd7ZOiuYXqqZU55ydflTg1pc/gJYh0EXJShifBkcb5W0EUDja
nXylCQegXtBmllyOnlzk1cKzft4nrSL4YlHpevLWzilD5IKvYerHe6t6hia+rm3Y
pyf8bT6LOYvRbAELjj7K0aTWiAr9aiN+N3l/EuoodkOL8cZBvifvDvwJmAA9lpjX
sdeET8jsAeNKO2zW3FcttkQ9LYcWr9RSjh5pPZeGXXnPHMvR0CYT3exOcA8P7K41
npfNB0WJLPNZbXO2Te4UTo37FvP05Pj0AuqxP3QO8Pbj+mAU+ELzJPgEtHzfx7mX
DTUYwElrG25p+g8GE39lyT/roeX4srkt0RCyGCZJ2npw7SBdhnCn9mGbokxru7E7
G31FzTTH+Twg5AW4Qdv7VmbmAAqfY+I4jDC3OmKSTjSwx79fmpwjU1Svmuf7EnNt
2dJ+oRDSmAeZ57Gri0vmKL9nspxF3ZsLCsblINK1mVf2UAocGYACn4tSwnuGsEU9
Hqc8lyHAIdrd1ls7mbjOudZJu4tKTHjSXmDO95hhcuBCHLH5nU8BPzeYUooA17U4
5dZweizUGBfTLIuXIhPEtdrCD4r+Dp9K2nSYEfiHawgTSiXkrY0D3N33ZjKcTtRr
U7oaVbI5hc/E5P7BseSdRpxRrWk2EX1KJ9eoHVVvPWjuT3AQucLX+xOWSeWemp+X
46Z8XjXKcXjy8vdTLZkIhyvG3H38npHbQIMzFuf0X1Ey0sJRUElK3QKIEkE2fLCO
cmNykpx/Yf9AIxHxaBaUENwX2VkpnFPV76HJRzgoet9WetEeGJ451JoaTFVcPx1F
cBwNI2O/UV/WJl7lBnXI1qlMcqGKEDLPEBYolpXWeEC5HS7kUbtjZt0JT4VqozHa
SsT3M/j5Pig0tTakuIQvouJhaOS4N/XX6Oljs1D47KXhYSPoe18jg35ERurqULa/
n/wFLpXmNwHaDUFMTSx3ieyF4Auy6eCqXOLbaVdHDpkMHhrPZ5z0+28KiN4T8F8z
/6NarKNPgCYdqDh9O5HqJYTm6ENt+vknPZlVaEMGRclOltOikC3KECmwJK8xhtl3
t+fPl3xBNNuYs91thuDMz9nFNNXL5/ZSLQLqop9BNze6dkE/+ofGK4q4GpndSacz
GIpTRlphIpcZ4jY9+pMTuzE3RBJZrH3go8/iTbpy/GgLPMybxeeoEVnAkFo1loCu
GvEEx7Eq8YlxKOAPwghPlZtZAeOHFO+hwjfSgLuj19ZGMTHYaAD30hoByCpKwDai
BHduWO6gLdcBGArZQ9dqN+aVWFN0+rrsnb3CzaKKtzsN6mLHVEBLR6CBMdeT2oJU
zjxUG0sFIimq5gDlYjPCz0jHxd1wy9tk8ggk/6zLHXB3ACFMvCrnQWzG6aTDgNc4
PFAfagcDI9xCmCP3TVpO8YTtSjC+5h2J6vzua6e/Ay55tqijwxZd4JjmjOmmnLFk
hsYpa3FaWdIwvDAAM3F/KHcA104Ru4GVuqerhqdrghAI/3p3KBCp8mXk9lylQzb3
+71YosHL1oLwz52GmuD/Az7py5/gmlWB+OyHM22MGafAY8CeNYWz9iK2RbUPAa1F
xB50PyYcDBE834d8+ScBYQ5iZjqP06kHDi10IvmdSwfEaGd7R/A1ALHQtIyW4k8t
tGp2UUGNV3Rn9ai29M+0iVdLNbLPzWyewpC68GcQ2oNO0+jbidA00/yAdKDYxFju
HdU0FKGtagYlK8TBlNichpZQ9TU/wisCZhWmm8mM7Mmpl+0jKLWfg91H+Zrgm1vJ
wANiSjDZvdvBTI07oHSiHZVis1TQG1CIBPhDJqMaQiZnD1tDHuN+fQ2hWyGpdkRY
1SYIWKJ9TLwC9TN2MBs8N6nkx1FyiudadhHHK1AnkX4vTBXKmYCOuz9wLLdX7IxK
+mQhiq/UhIAcnlNSCC1+ziIVG3kRac1h+wDO5r1esByL9dA8OfWPfiztFdWgRA0q
pLlk8AZIJ55WqtJcA9pVSL0gBSNXok9wVGqEE8xMJae6jL59RZ9o+U2feVwh1tBu
+KPgQuxcCyPrD5fQq9OBKZZP4rJ864TQJ9vWFdDwJCjbaO3YnYFfO/tdvFa4+JC+
gY8jc1Kd6JjARjizX6QNdQXfJHR7+tkQGkPhYJ5enEkLMyULfbzfresRMrdlodA0
HP4TilWtQY4Xn7nnahZQb+wyRSUdrM5BERVNHvPCeOmVHz5oI+NKPgeU4RkFOXLc
w+NEZdUBUn8f3wIcfjvnsrEn3MVsYKwoc50lLDcWXa5Le4PSctXL0yRBumYi7YwZ
I7Q6LVRsdWQJaCrEnyHtjivhbmU0j5rW/3DplDyEtwlwZh4Qll24O3ZxwzUSeCBB
5mEls1czHLm/zkGCmMmp2cKfs1UBCjda4rlH83Au36qTahQTIm7UHt+DKkXOtbEe
upOBzmubF+3sSGAsYmf7hP22qmT1lABi3Nbkn/ZPlyrjXRVGnAzOjgUGQx3sN7y5
4WP2+nRls22gxvuu9xlYf4G6BO2JOHgbtNL6z0GDMt98ab8cHmq0vxwIm8wROCNt
miG894p0fbncSBFQJoHI9iGz1m8EEMpdfd77b7ClXEaunMhC4+25l62azhFyRBp8
RFYn9dvB1QE6dSmmt9hZUWIpGhmKZtkLgs2Bf5zRnfAIABd6qss+kEn+nDkbi+1x
PKjpntED0E+8OUWHcMx2+db+GNBVgDhqpUbGfMz+FUV5/j8tKrKJRPWPVyePtmHR
nCk79yOTXX/JwbsGfOlQXoJzlBfln0tZqgGU3+2d5M0ZDMRlMI7AjQjjASFmtBFQ
1GJX5l06+qlH5vtH+tlPMjwTm6DMX2nYefxPEq9rmCLLmYUNHwJHvDhbXsIQM69A
Hvau8v06bDjVHQiMHEWQzAVkWXqqCsyuDhmamwkrVZoEfT5ckogxMGLmLKAjVU6j
oCtWHv1eJkJ9cegXci7zpb0QlhKO9zm9ST0lexIJ+NP94AS21BJmaSUBgCR2fsIO
DN3m6ZOkp80RyCihjbkAzs66VqA2UdhSVrbSkMAeryXDKXfdKqXajTX85aP0vaum
8giAy01xzX3ghqPaGt8A26Jckdg0EOK55f0O3D6vZ4BB+TDkYZuTQGQ+p7eFH2ai
P6AxnhgLFp+trdQ9iWI7FVuug4V0S59LBIyE9TK59LYoM2AhPb2kTkjpgry91NKo
jPpW4t4yXet74x8uo6aFTkkALFLkNBQTCC4gDshJG/DhhQABQlcsN39o+RUeoXZ/
2s7Hy7+ftuskSvVBr58DcjrXVexxV4oPjbvgJJxZjBMO2PmXyg4KMtIPDTOMhalJ
Lszw4cvS0Tc8mopxQMdd99eOhhtUkAsK1lpx///siSJJL3qqcICoYijxFldi6Vtm
N3s9miqVIgMSrwgZyGazpHzKc64kw3j9dxvI/l708uv+JYbAieK4vCZcHQQSas/6
Ewf4VymaL3BQ+s6pwCWabiri4lj3GHDniCLWiY0hJYmg/+YvoVnyYee085RKD30p
npMtkJvm0PAg0qfR5gkoG5xDjotAdTPcM8XqDgUwbdTjHf8jAQGx2xRz3LZKlQ4D
eG+R0ofwCJZI7hAHqRLu2OIXGBszDlFHMdSVdkgbuHU7iN8FKAuVtbTutXhi4TEs
4CiSPmragsYn8kuUcqEOnflxZu4Bwh4YG/BEQteAQZcmJ9OIc+l8cvr5UANlFySP
8Lezmvtis209jkAJP1eJQKs+LoU1hQeZ7pgXrkpDABYXWSp52nxWLYr57yXWoIAI
qxKkjKz5hkrCybQlsu+PPZ0dKsXvRtEFRXPzV0MJiCDbx21JJu8RNi3mU9cZ9Ubf
8oqasxt+HWa8+OqxIzDdj66669RH/V+u/odEklU7oUOl+WAEOiBP+8awqYQZw7pK
P5KnV4VJ1gfp8SaCOH0EAah8LWOfKw4NYMHy/LDJB7nRSq4896VJ9iBukoTQ/EjK
Tw8Pm0LoeVQeQXkHX8w3dVbPG5yfAiN8mFvk54U0+DzPT9+nWbk+Ydd1x5k59lma
kKa8yVRvLI06MpeOX5+MPGR2u236OPp3j+5G1iQbTm4NExc/4PpgWDfoluTKe97M
SKVBI10rx90E2mLvH/AOGiTAUy74I4a+0pGk6NeHnyeRoqy+6eHDE/JeNDMnOjpb
xXiLPTPRjJfmyuO+jwPRj/txzC6QfgG+4WBagznTl+XigRy6JEuSVSqOqNWIU5Hz
TsB/WLfnro/hNi7csIkKkEDoe448WVYQF3/z8UmmxrrkxqMI3Y+nlq+i3eqI2Bqh
gpDYSglkEUiMn7Ll2hssa8nxghFpLLA4IafWujaO11K6Ld4PQUPkQ/B6hSYVamLF
i6Gb3Ge1vkE8cxewExsE4FyE5qLNyKj3IcDLvFkudlnVLEzYAXqRPusBkeuSw8B2
TNkncQZOoe9q1aCXCpFNo8X7W0ou2CU1C3zFGTcBWEqrottVLkqATcEJO4oAoEpQ
uuRR5ZlfOQPBEdfsqBPpDhEW9Ucp4XHVJbJvcHk/piqghebPjDm9UONTdmZbF0Jw
Fm/aMWH1pHKRcGUQMok5pIbZaLrh+rC9m2mfLAtg++dO/6ZXXqZErTaMoe4ZRflu
0ByrMS1wjfHXV61vsqmgDSopo5/g7E8XnljxJlZOGDeRTj/9FDsZu+/Czhdx68Le
9+/UB6LLTh9jrEL8E3l8KFzbrgPXUBGcNxtGo6tamP6vHGpKktvTXtOIlmARzAIU
f+D/x0ch/vC9RNgWZoQNLEFrbNm/xW6GqmU/HRIhE2mkI4cTm43yYLYvFb1AYCG5
rWYC3vztn+kxCRQk62XQyvqTlIHCM9O2k3QId4fW/z7qqJ5QetzQ8+b7meE2bt4p
dYK0lOs5LYvyN/2V/EA1/moFej0PaKb08Pw61XJeqhuo7pFzTh9WVjO5OY/Gs6Rk
DJ8E9XA1R5dag9+DV20oAfoCRpsrRMsas2muEJNR1LrYPm+AZtZc4pel0WCyI2lJ
QR7tUkVI79f4d/KSd7kP/XH5r1SPmOlRVN/xjILee0SZ7skFiHhqY9C79U8nxLhR
1E6anfOgf4cWId4jNOsqlF5fx4+lO5HeIfggNTWA0fXYyk5N7hP2N5pTDdFHX+gW
rtuI/QHLo4aK8JKyHWB9WdhAIRFN9I72gWm//vsSTvIZQ0wQH8bvhd663lItzbIQ
FeE3PNWZ37dgVNkJ6hSL3Yvd2t3lWKGbKSZmPLzdd2X4P+DRNrjPmw/7v48zQtS9
m8hpTatEfVhCf6PiTIr6KX1RK+jfMq4DFWF+l1ADw8qIw2P0YjOwUVnLh/AzU/0/
vpFwAI+GycBOS24tcC8XHf4vHOxd3ipRALYwcbrfCbz0bQrByScm+8YztRhDNMkV
ZbhDoz/iddo0CnPjODd0trHcloZEGsA6TwwYfPpPsq3c3b0tvjMt32tHR2u9GjiB
WSzN+seSQGwJt/MVGchmoDCQVM3XjnU8KPvCQEOdVgQgWS4oeapbhipSFAGpsp/L
Q+JNmSa9rJV0MktRorO3JmioOslOJhRjAb9Apdc5iMPUxS3q3wNQDmr3d8lfOy26
minCt3KxBeWeb5cTGhMyin5uzdZkZxNT1Sh0Z7jSzE5L5bptynlaQLSHoBzHrItz
Wv6/N1vK3jODULfPynJWbzGm7ZLv5SKrbJv62XIN/oK6zuvCfCjV6CYFyNilPLBC
0yud7sYXNbjz+k+maeQRMCU2iFls6LQn+s9Rnf87pueaCyKgAjwWKmrYGUOCQIPV
7v5Gdzz4P1dGe1b8IQzLwtGjENEM48cyte5gvWinotr8Edaq1aLCoiNfUHSRSHNw
tI+DFXGaMwKGf+22+c+lRutyw6YojpyZUSSeBiHOFl6UZeSzC6xxdE6pag2eqAnc
TJ/BzMWDtajft1inMqB4H5MclJheupAAI3FwJeQk2ZlqkBiDCDfPywQsMsvbaqVE
oRynogzKWNavEMT7V7Swii7SHHLqsNAw53TiAY0WWAx/Q1lD63ybVKkPEIwV9doX
fpW0zZS8Vbhhg/JDOQif3VBWdi1LGg4MFbpk83X0kLZWvrSCx93rmAXkN5DKJQ7y
EFqKNA5SLuzfAwCy6SdZRcB4H9gQuOrBrEWxYPyhS1PO8JiNnSAH5uYXhnMD9sKT
HmZ8TjhMimWdE8VVVBhJaW49AQDalq+0GjeBzdvVjARD4pvA1do0vUQ3+h+wyGZd
d3+eHY95EfFWdvckANPvBVQgR2bLrO4PH0f7QYc9spEVnqYJlYMbd5HDJCzN63ub
FR/YbqIVemuQfBZSK94Z68jLlG7D4dXD2R9K/cm3casrkoL3VMVpJy1z1wcaH42n
guouq0NldrLweLVVjb1odhkIySq1p5NJ9x+V2I5yhF/V8FmYWPndEUqaZ8sGIxPV
HeGgZnowztKhLDeQ0qfEAi1ATDwVZykZ4TFmuGwgySdC54M70+vCNZrupNwRnyFA
K34lha/sniVcSnvJoBtptASVlRPcVVkoa3xyeLNbtvM2+KnghRB3dFXMPsMnayyB
BAUnduAvj+gYOx2us54pRKPniWJIbrAzxQUhkQqzkX4j0VyR6rpCSYuoYVjMqRqB
tIgkKXLauCVRVyeLQb7pCDPbZROR4WJS8oCPb69AQDqVcnY7acQi5GiPFaMYwZVA
4AHzcvwP1stFoRtEt51XVJLPdu2BHisyyiyKxxr4x0new3r5BT+RXrlppSQgtrgH
v5If3IbAXVdhYXWpQEcya8SqsqptmB+NHB+8DN1dVoKuc07rJtapALj7PnKnoI7T
ch87Cg7GgeP7cFFVLosMOzJamjMNxp9D1LppLl7KEy+rUbgPyCjuqPb4MeiyIw1Y
1DCZPGNr8wPF17UdbK32Bz6FMRGNdDWE/RwAPLBFL0sEDMA4KgCPhn37YaN2MCBn
BDOa5kaIziKkh/hK6At7ZXfR70HQV9YdZiNqVpfwtNmRdfOTTdgcWAIgLP0OiLzq
crgk+ot5INBg5XCmAOHkyOJEczMF5DEibigI6sAuoNLkNDN5eUOYUtHS3MbDijeR
oclLnkCHoEbQa8x2ik+bnTKPl6Unx/qGT/va/RVFMhmhwA1XEjmtIdDh3tNtg+lN
1MTfGSNRg9uMAnA1BVVzfSX1oky1CAUzK5ndZ7P/QO24hfBp8D/hj6pX8uoudxI6
z7/+vIkEEeVhTUkABHlUmdYvGZmQGAzeHvCo9tRVr9Dyclewm1uLZbTLa62I97py
UYVJsQcx6iEJ/+xKugJBsNqa3nfQ6FE111MfspePGPLPVyK61lrDpZyo/mFA2sBY
u21sqkERY2z5sFXQxmCMMVNkMeeC0c1FvHcnY7Wa3BJpUQexdMiU+paAV4dnIfUN
7QTAinURfB8FRItxgGVxgGu+TP65sw8mUHR7+zsMQCutBLcvJRZTuoFCX8/QWuaU
3T2pJVWgW/rNXvbEQrXoxhfrIEZmQ3jDLXDxPiwVgbN+qlHCucSk/7BC/XriD3Nx
a4x4HQ7n2HPjTE6mPfg2usWSoczTPIQ0nDQANlvnrXzpDewngNWbPCD8F5P3Z9NS
s2roABKJdaEUK3JWNgPLn4q4Z+pW5qk9N1uUHICW00v9R9VLG3reYR2lT31llQIi
ulgpJSO3o/yP8W5hABSKCDIqeqljFrz2tlYo7xxinIvy4cJhDGMS7rVJr6U72ZYC
gxhdvcDEtprUQZ/1RVULYdwkyf5Ja7NV1XGEa7NS469lF/Nu8QVBuOYsiIrtqBZN
KI843ZCzuRF7nyGeDda4TaZtT3PautbcYmClm1klTxperbTD6WaCpgdxhlGJdNKo
szdSijaBjLj3l8fl5k+3/Sh3cfMXvWD8LjlVaS4Q/+t5J/MbAqNuhCkj6nPeUPs2
9JWWN5+q6WSfMFYWXISMFU7zndPrG/CZxOZACPdmBzvab9C7Pkzv5eaZ5k43D4tV
4MIY1KW34dY4DIfgGoz1XQVtb0Sjyji9rr6iaQXObCoWXZsTlq9ENXzvBXxNcV+X
nquZlrDJxj/GvsSINs6rpzYKm9jPRS4lXOpf41C9pR+f7eO0CMcTiH58zzeAxAcg
E2TfRDb/jAo5Mx0mPKAKwjvgZ1aMPKhYdNysTAhWSOb039lWy8ZtUF56ZuKNtN0P
kVMvdXko1fNd5xjMBz2GiGQrOh7ZyAgt1pWbm00jd8anhDX6Yfqb14RM6MxWPHs+
nJwxDZZUv6shDdX6J86K6RaoUsojrxm7vCJpRLxdQzKTq9oIngEFNLkjAvpwPe5J
wdjMMk3T+XkDWg+kK8i4NLZfP5rYweraP48zUKPFum7Z51+avqh2+mOLgppgSMFD
PIJzPrBFozV0HHIBEpAlsqgDgvGkhr8es1HTJ9oJEb6cHN/NQ9mLrRwDvMwGbO2x
pB/8fAqEXpQkfeVWfvIPhRLY+FtsJB7cuy1nl3xO0k2oxFyPYO1eWi2CLRB1q87A
L12xeriCyMorhpnlqpDaVP/UpXxspRtz/3PZYJrzXMaz9zQ0APi/of/Is+GfeVJ+
HtrhVVKtfFuEDqOi+YcTwrvPeX5tcRRYi9wn5F/iwHDivEdQWCQZYBib3vLdRYeU
Imi/Wry3A8Hb61frRKWXc2pJhOGGvGLaVuEMPe7JCSqdBnJQAfk8nYINqQgPV+zf
z5P0b2cKjckOecMhETZTXm0+eajJenECkd/GzxlWKSEad8S8CgkJRRp6YXMujuSf
gAb/9FQHvIINBdcx1OTjvzTf2IQwgt6/Cd/ryQUx3H/S5GiGJ2zz26X/qSEFHntY
oOo6Gfj7hQW5Tkj/C1uQS08EbDnpp39z0E9NK60vji1gVNCecXIg52DfcSqKJCyp
tqiffJEqErtFX1oVBgd1eVtmGJDEqvFYCMVDYq1nl2JerxHngzDCnnA4aVMXupGv
v23a+MFCApB4yCHQyjyDGNg9ghx4RKxFb2cLTc45SHn2hm8axxTYHdsk+ahEYLtj
BnvMef6B1GHY9h9AwR8kU3b/xvbTpo2rQo3myOG1+LE6N8ua8GWgkmnqX+QnRRqn
zsTXTsotmaK4M5zwgJCkfzTa4hCEyPhlOKTK3y5cWJ7BMUKvRlr9ZmALObe1XSOa
87lnjazONtQKvTfKBuQUWtc5Ged8TlX0gNZl3qSmNXsjsF3ZKIZNg0QX1iEJMOcv
YsMNXRlW0fBhrHDYPbi5iqw6tnn2PFygLSEmNSSHNKiBGR26AeZb/zO0TjswB26U
zWa1PatQ7UWBqdJ62C9aaHkbVj+DpVKGBj0ZyR0FZxt1TRv+jO/Ak9kD4RMWcvWf
siza6tsjAtqxP+L2kSgpI0e4eF7ZgM4ap8DqWEHof/3DE8oe7x8OuIyWZvNtMxDw
K9y4yjBy4lN+TXds9Tv0BXnd/zC+TTd2gen5wf9/PNJNPH3bHmL2sWqaiZZx3kwA
31S1swBb1XwZziHnfC+v7MOzconHtx5jAkh3b8OZgPGhPjfjQKIDdRpbQl52ueN/
Vl0iDmB2AY/LNqX1IRSQPKDeyjl+mUaDTDWorpUlHA+acUT3X0/wHhJeEBIEsbDZ
Y0q59Qqg4vJLiGEhjvr8aqbWc6awmTiw7xLk6OG/Rhto5RPRWNhA/a0apAFBrnX9
1uy/pb0csb55MagXQA3aJnsOyq5C/4eN5TypT3e3gKwUwTFGBoFXlubRBoJzQaqd
g7kILi5pP0o44T8dwbOKs5hEpSGW9bRKRm/R2EzZ9KOg67lhfkUAqRSK8kIEMvNH
GbzQKPmpXgmInXn/Bclun82Jm1L1Qi0eT64FXkIH+Aa3UIMRcN0kUsqzMm5YvjhL
DufOvVIQsJBbgjJcxQEqwfuWUQE1RZQovZcxyZE+KxjElrWXNMgawU14hJVjBi5w
MrjccBy2ItNunIyA1uV5FPgvyAExALkuy3PjBmNKVSsj44T6oJHHc1ODct7Vxi0G
mw97PApnxa87PhFqYsBAPODS64efdlth0mGLTPST6hOWV4lNucN//QHos3rZ6Okv
CeaPc66PiAjsG0Zj2afkBCzxZQBHmiywj6xVylT73aztLuooNJmuLZ2o0hsBnw65
lOypGsaXEnpUQEkMX4aXPRwq/PRagBy93iTTVPEbWUvLJIZDGK4NvpXm1phJX0qJ
yS9tWKkuM/nQRBXGlDeTMTWMxBbeUI9ePFsYM3ToCqrHZO65h2kntmuLtmmcpvLH
XlIs1Mbv+wqdbW+SBqn93uXlCxkSJk+/tcc/AXJCPWmMpvgdy5unvyH1DtcVepG0
e/Z9HMr9OWDlu2z9B6g19NawLPYPuG0sUPiGMv4omDMWblemr+WU0DkrePcB3oRY
/rq3Mq4BNha8MOluvpinkASjv18jf2omfrh2JGmC6uH9nYXMMZI2ROVNr/HAXGOa
bg3GZ2qWh6BBNKFlrQwBuKjzo4kzT0v2PGUpL1Vq1p6OEuw3ujHlv5yo2x/IpF8t
znXek+P+pqZXS4tVMUM0vxiHf9s7HnuGKd5z/xDfTOosAR7ryQBw6DGxwhL/pbd3
gmTrLXYWC8mFtC93LZSu/Zid6cpwdE0cF2Zq1guTisCXyNcxZKJ8u0nq5R+0CU10
v08tcA/8NLSr+uccemv5SoBFw1PBXQ+Olyi04CSS9Tobdey5x0cRx6G/6/AXiC62
ZWQ8peh2HKz85uxTz7N/vxCOQDirFX/KzO6Oi1VSvyw0U9/gT5/U0F+SOwFBU/7q
FFgzhC+NZ1FeYPad22al8awN5kbGruOTNDv6Wblfdmpr8ZkKdSHsg9DiVn8+xJnn
fYIdeanbEswpVREbXQIZeUmSJTR1upvKNRqombwzfWFOPO2+b4SXyW7z+W026vbO
/ok+7nxM3mx5BGVCnjaHz6+RRyadnRq022M9IfjOqF1u2/qg8w0KI0RGDYKElnqz
S5mz7dpEJgDBeDrF5mYc0PV/GMFmhYwEp1BEDVpfsyDMp2xyw4NgHQqwlHFsWHDv
tgeOgYFXeG+w541IoVfLQRnvhrWRtanx5or7wnZCRhsx8+GwzVoQ4clu79RwBU9m
/sEXuZFcUKpAUGTibdh/XYRupj/aHa17OHWuX50xGgzr5zAgT44MiV8chUAKwNbo
6xoYaQkdK8VR2ITyVc9wTRl5F/rqCjuI4IAtDb0Q0zN1F41pY4b6B9ns7ZhPcww2
++xmSuXzQ3eFHXLJIiUZQUGFtacCjlneCcw75aLKmU9gKr1tYfp+Io13QJCfDzGu
5kxwyiPk5bOVsmiCZkMIEey1cAu6Aao7jageirJ6JAdQeETOB8FGWJzcRQ+CkrdB
RS/Zl7G/nJ00Bx//6wzVmbVxBx/sa1Os+oxO7xC9qUYc/xzcrPKwaJQnInlGhncp
o1Ts1D4dbdTKh8E7u6gD+LwcPqMoUnYle/mvm191BjWRG0XXTnwSWWg271R7AUIj
C6/ZsZoanv6hgJfUTXcdqS/BZ9o731qGCuhZ/ml2Mmwe9arFZ/FTLJy8mhI1oDj6
wwYBsuQ8rahvkofjaeVdbp010tGocszBvTCVufkznVfBCu/583O9AzySsXUxONFV
iwg9HtFV0b18TVfJPSNbHKtvZUqhSDUd4tzQ4a22DJwWSKakqQQlUIUqepmh7LGG
/MjRpjj5w/gUxhrFDdni7jFgoqt/rDqW7xm2U8W6QomA3Cyk/jSiEK6kzxf3Ad1E
v5d8GXoGG0gVE8dXkLs/DQ5Zgeu84icDn17/U2HSZB/VXIKCtu78PhDhwPEvnWtQ
dNIcQ9hIIt35c0KQe+a8Koht/J1z3aC1tl9ezwruFNCuuE7wreeOCpYz3TlxHkRm
TP44YJFQCH4sUm37FJt+p3GZOT9GpSyc2Qoyf+JNT3LXqwy3YGZNX24/Box/gD6m
komYKSe4dupYMr8XQk+T6yEWURPt3G1U+5x2yQmvsDEPx/o2ynsAG8PSndvYFh1n
8UVOt9DtH5jpfunegLz7EJGwz9KlWZJ19o6krnMbCg4cOuPLCvcsjSAOspeNB4eN
hEgVNkoHWYbW2vzFNuvu5/s23YF0k644vqurffbnugZ9s+IKt61eZcysrSwv4Lnw
cealdetJ8hk5Lb4N2xnwf28N0LrPCI/3v4q5LSx0KSn5f0mbzxZhTDaKNkJMzwDS
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
IilUZTB9cV+lyCviTdNtI4uVbX+TiYTsAfABMoI3qbXhNc/9w5OT6+FTFGOaDZ/r
6x6K2/54ocEAoEtR5YRpxcDdWu2XVK2Y0p0bdKJiUG6rNOpW3w/l0kn+GzJbO2lv
St+HpbxpHytvFAq7VKFu3V4g9kxr4TQ8FFefoZNVoaEb3U5H/IriwQ6MAECIVChn
xhunL/Dsvs+nrv87CrE/EJx4dksxDbXb7Z1IIPQH7RkzN1UvqAukPjZvDCeFApIv
mu9d6W+oM1tviNER4jh+IeTxnCskfMTAvRa1P6Q2Rde0LSfEAzLJnmJn1SEvInnH
5jkc2kt6jqe4tiZPzQgLsg==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 6256 )
`pragma protect data_block
hBxrUEAH1pdlbOAcSwHM5Zrx2bQmmX3Y8JDSAIAbT8vxuzHrvDJmBd816UFoxl5r
01aNtEOjmEM+tGYfYG+PEG/DFiMA21j8Ar5GkWBqEKEuqUwf35jGp8IaMHh3Yx/K
fF1bHE6/WsQPbANLVv/e6cSAaveNZ0oFT/zUXCZ6qW8U9VsNSACDLt3Jb7iTulS4
ogfciPcynw25nWe7U9eHFFrfRKlu05J0yZsJ8KRkcwQ1A6YkqL/rfUCg7L1bGijZ
IxeXXOJME/q4kocTij+2nYPFODzh8VVaOvIwnxZuVTcIbcBnDIQIV40GIdhQUKeP
cvqiLDZ/JFaAMYQJhDPkabsihdUQNFn8g04aYOYQ7eyx0qgQblPAhVdoBKg+WZOL
st8jszghUi8R/UiXk+zd53ZQCfgegl5CqyjOUpDRS8uq6MhlUp2CuJZw70kqurNA
2d5YpcXjzs30uLiuaKoyJwqg0AxbBeu6QAmj0GehmPY/fQr8yL5cAldlZH4+nMFT
hzitHwWCZys9gzy8lKHwhjjX/J5XReqkxPFOJIPuG5SAzp0oL8HAB5N6Q3n/zbsO
YCYczMNgu8Ob4vImKuO0kuaG8Lmn2VF3MLqFwiSAGGkmgT4y6UvNahl7E+XXYann
TYeZ1EU7OsTUnwjLRn4cxVweMP/7agK9oUjobAiSqH99pwg8txhlebpGAh0V6YaV
nBAh/q/OxtD7Ow0jRZ/eDYqbizgJvnUhEn+rDgUKkt/Cd/GwATzMrP/hYkyzgKJZ
uKnKubOhlH9H8TviCjuueKvTJx90YGNqbLeCUHaiShMkI9DRVKabOEHcx6BonZUw
+xWpWlgMzc9HQneSSXzPJbq6b671OJyTHgvvN8itNZ9HzkL8VCg6zVcCWMQuSPbh
Y1htawEPebLcwGXAunIWSwXSEu8yNGHfhush+Ue1CrWzoaXOXvJ0zr7fzBsyloP8
DOaVjU8LIGovn7F4nMGRILC8tgC0vg3/Y39vYLmKyUgxLY/ERwWcUh6NQ+K3k+Y/
ifjFynVZWh0X54Tr7kbzk3DBq5ZNvdIS5TJr5IL5MP2oAKszXrRVa9qd6X2S1L/g
QtgbisPeUA/kp1yN0+p8CF1CDLBrLCpJZ0AyOJ8Ph3PVW2WIgEirysHRgumF9PLs
pn8ygXEEtrNlSelOUBlIuGbWxQoQK81qXXSxS//pxbsWcZwUpmCVJ8eA48cRYkKo
wO4wXfsWmbN7CjZrxtIqg8lr6lDEUa1x1BjaSkfdCstYp6vHDIsCEc8IImFFSLgc
m9FL0dlSGFJW8Cu1qPjB79pSOxc5D32MlKuhdpbNGozPEIrLYaej7gtzN81eWf4C
1oVjrKDE4leNQw7bPb/8NmXsDyffeYNZMoOt0kO2PrC8HXNBhNqGEQ2re2NtYicI
TyhdzOzCqs05MaXKFCTsPCDhP2Zc3SssXSJ0srMTkpkpYxRVX1W4abjaSZ0FBHhf
vf8rshfbJM6WgDWQfrTo8d0YbEJ83sTETLGZbMyfRVeJR1gBy+Aw+GyRktJVEy/b
UxisK+lg6l72O/9fRferNT3SwSrfG5U+ug02bsl9MAOoCLNtyW1tq4jiW5C327TB
rjc53a/il+MVzIJp1HUImvOQr5npShXcjveY0pS5gfUy+kmCyMGBuTRl8NjPTUo/
xVkNn4qh23VnmDoP4GGQmtkAs1u0NHEvuUxuWkiCDYrmwQdOKBLKVmXEmSWIjlI+
GKW09Rhbo2NkDbx3YAMdp/i9YSRH8EcHA9T4ipRKy0iJsnVtYPM1rQ5azFw67REV
Zhkry4DNfkJv2+Hjf6pi5QnMpIxc+UqHJJtZiQfmdcz468wufLiwlUhUn1SnpDth
PbPxyDX04yAglyZnng0K8UWao6OuOr55cBYit73S8upQUGuyKTV/rXLTpKldD2M5
W4wXRNOvdQZFbiMSBi2GrJsua0JNYnYiuLqB6Ghkj5oREA4rc+WKHWP4E3n1ur7g
tGbYieV7C5TIeUjca40qqPPmu9X13//5tswsCbm2pRREuIWpof1S5DaYWgoUCnkQ
S9MZ/2O2BsHjy9eSFw02QCmfYoIm+t3/3QuSdpQc/NcBwcTA41Ut1YjkJUVfwuNS
z9ZH9aVYXU54CUrzGh4zta9nLeg87b3sNZHleHOObwW8Gl9iRDZpMbkeCWevN9qz
NciWUPbBw5TLcnf/4PUYXB05BiG3VK6BROQLbbE3pcFdgbONaiqvuPbAHVqgmMHd
/SrPF9SpIsLQuc8zOBArY6oLRyFvqtrrCUCgDGR/4a9rTtjesGKcG9S5PqxjZF1C
tP6EAyb+6kgpe62pt/CN8uTuFVi+30qI4IrYSaoPQ0nyY7mqewJByr+qkDjFSMeK
e3gWrywjtqHPvI0aUfwLts+f5QjiiQJrXjNreEKZFICC5AHPFKyLysHkhBO3Ja3B
55NVjLEaBvVlOZDIK6V6x0zMmHl+jI1RpPunb7tCwfHPAW0eg2b6TKAu1rD0YXXh
zwofBBeSlopm9c0WszG/RVT+4PDvFFG9GTTs9JjImNiGh9YMnkxkudzGtH72OLcn
m3Y8tAaAwz+vlAxrxmuFUtUuw/8TXd/9F1PHnVcQJ03lRPIAzJG9JdVBvVmuZCOY
xtfiB17yHrh8aUhwS0nWBDmJIs1h8GXB2seYwI4mEesDlrhNyhGGFbEJQtt3Xs8d
zULK5ipe/uqVlhesyKkj+aeQUG7o7XqA29/6wlFuFsUpno4u4Bsn/Y01hkj8Wb3O
XJSAHnZvpL76abty0kNyIQJYuUdm1FJqAthcWo4ejj3rY4yOn9hxi1SfIc/OmRZw
ED/AtW0Uw+3pja23h+1j1ugqHcimMB0vX+szuTrIyEK1Tsgk5tzF+ZHtmciYJhPG
LOO+WadrYD5VUagd3OL0tnk59e+N/6K2VXg98pQtSeNoKqGV6vphvsZukKhHGCXi
/8pDpQoDJSMgalI+1xOGy8LKOl1h1E7H/XxGDQCYEpCvIMOmShur+8tVfCIDzhPu
AixFw1jrzroMgVXJkc6A5grUqlJTk/l8sbbpUF/E4VNuLUQP0zGkijyeFq398m4l
2i+Ke7JT/NfTNR6NgRGiDbqhepZtd4Y+bDCCCIFltRWtSMvLUtBl8R11Nx2OzOcA
yuTk5HWpyAsEehgr1cm9Uulu62mMvG1RzBATMKqHgL1uJ+yddRIbSY+FHIg00jVf
WkPoegWzRfOs5B8kCXVdu5tXN9gYTrwR3X5wc9DctpNjRd8BXutqnWUYkYA+ej5p
De1EXOcKUbcegGalrfHno24+0QHw8W0Vhz32yewl3qpCL14zp+Zq7IJobFN0qekL
CGSqXjm+eKK/HjhXT+20ETM+FMIn65A53GL3OHaKbQNcw6ZXr5EZLSHgbayWKb8b
bE9kLEM8WyObzfSD8ccFa0VXiCmIfz0kK7sY2E+YAV8YAl6owt7QXGpKhzbWujTV
r8PBp0WueEBekiB7B8ewXIWxT706S77m0Kv1x2WyMAWQ2SsRgapSBb2YhlSZKj9r
EvgEmuBpi+up/oubi2edlg8ZIShd6J5+gr7uaesk0wdCBbF514izjTIXSVsFNb1Z
EIUUg5U6xxlMsTsjKfpB6ACMm1Y4iYntD21BvO1lNhp9oh23miWb34/j4xtgH/G5
TfajJtuxGXbb1eopFmbE50H4OFqYwAxYOVOspjXSnIBJWfUfvwTgyOGr3sqpEgvL
/lUD8z3GqV1NphOHI2BuX9N6XM2DuPXaqN9Vv4VtN7zazs3j7OPEGgcJ6LvbMJW3
gYsDL9bw90ZOtvl9zxkdxIYneD/tXzyY47flOZbGfdRhacqnCjYddRMG+2nrDUyq
pfVdjUA53ReWjagr4Vjzdy+ppsT8QMEpi+AxGtB6iuQxsCM5JSx3iXzY8BR18jUP
vS+AEPO+3LDKU/NyxgwQ6UlcmFNkePhaQCxeSt31f2Gkj5vZkd4f1PMYTFKhSqzs
T7eoKElmatipKzgGbUtqbVjqI9qKakmwg8g0cuLZ8CVou4OOuPVBHrJzw60c9or3
j29apg932galJmMxXUf7ISy3BD8TcRc0i3Nazz8GDDViDQgT2LBj+5GAF/jCnvas
7JJgJt/yh3H93qzOb14QD2Md9mYLiVCerDruQcRCH39rqtuTggzN+yldHe7sDLQx
62UOcYvoBWqqP0FbsmA+heMnbH+X6371QFjafrx+0DDMJBinNwE1eaDIp7JY9x3A
lATJidNWHNATbsEGaQ1RdrA3Rsr9ykkTjhO/iRkpoRAWQCYKxsS8X/anvjxKIUn/
GVbEf++ibYBl77pBCowHOhF1cMSlvUjFxzflewbgeHFgx7J8CM/aA6wNqa9vQW45
yhjZFYJ6dRRZRUd/yGNWWD/4pTlNkBN/EVq1W2/RphmAnXH3Q5X/Un4FK3+wM+28
Tx5gvMlR3N55AOgL3S6g6J/VClVvpiDOSNRjI12s4IfaEeZNi9jpf5hWgAm8Ts/z
HmZzhXWftxfiURSg3Lx3fFN7MmS41PG4S/2+yp5iTIx/FSocQ+Nay2BlsU4z7UZe
TaY3luNjRdvtfdxHh+q+L4dH75ps14yqXYtWSzmaZE/OVLDyuKVxLCksaTjo0ucf
82hCU7i1oiiW2VJPNeYxN3/N2n+YdfNaK62ZeeDGVFSo5OeimTkaAUC7iCcCgjjX
z+1mMnebYjzwQuSxYQv9Aap2nIKynh/3uk94aYfNHSEY36oYDyjIah2E/V2G8UEy
kLW0T62gl6bTnhlmjcQCVeOE6xlNjKSEudeN4gmfJPVJaDUIoXTd4R0j7TJV3F4s
EcaULXIiX7/6PyIOnwCEm9VzKs5r8/BPVruTe0+JywUsOKEKL+DT/DWh26sfvrEc
GN/EgCc1tMYBDA9LIdgW+QxGxyUyyR4cl/PzunxbYkkTEcB7gybe6K6ja0fXd0pO
6uqs3TxGbwDja+3xbevtP7VqTnPaBzFjqbvVtiwSDM8mzYTWJV0+wYeY9uw4iyak
wEYek06rGjtQhkqIVCj1lSuwDFuEwOsthBbJ54lV7J3bOnRjoWty2Niyg0cUY/eN
JP2epN9HcjI2C8kIX1LBVp6zAyOoVF4TJCqtApqXNi/qi583IB0J5eFbg+QP2+DG
mzskZmRuw+DHFi/pVWkI+4cBCQqM/+8Gnp5sYC6OYLAf5XI0/iZuILTFtPUfnCCo
lTH2j2rLhUAUromzVoAN/83IsqdR1PGrycp0j+s0OPy9xIUb+v4Wiy/kbjt4dZYx
fmnt5jLZPpYAMKldTQQxqx044PCeGzfVry9N+jI41cW8I8zWAPMVU+IlqK/kdrxE
kHgz16Vcikfr+YiwE0C7Cyt8eOi4EtYSYxBhEsS9oZG4ZAdJbeAzQggwOe1zyv8m
u+auKBt51L2ZqjnP1baMjT3XagfgV2taxGVatnz1yiJflonL7SxMoPFLWaW8QQVh
ukkuUjjDqOKUbRLA4XZDw/nsSNE4h7bfNQFxfYVKIfd8IGydK19mng0Nmc64/cSK
Up5N0nAv7cVpW1fJBYSXrf34IpDL0skw9mxMk0ViMwAtdzAwA559p7rg4/JNEuO9
V97Eda/tCrSbM41NutRS8qXr1SXiwkSwaaVVCkhSmjsr7RHJfB2c+3HhB0pXhyOU
s/QNSnPbXB+CZJcPtVrgjzTt3uPYJ5A7Vq5aOKLpqgnjBPjp4kAoyR1MDXAkRRRA
QtWj8+lD24oxitnr63Y8jjN1j5GswzE5b8QoAcEdQV/smAX3DyrmlnlITzot7W9j
U2rVj05qmsXPBDYXDCPU52QvCW2/kMDKtTuhN8Uev5qTiIoJBsvTI350n1K/pF/i
TfQj62frpkSJRNbIHz5TlDkygdx5tI1aSmsnLb+qxcs1Ow8jEn9FF8oFKguuUzxY
APJw37KqKC+9uXZCuThWA119cjrQ4h4QYcClUY3XvbkwfSP52wKDRu545GTkA7Kr
OJfjGn1eVEI6S2kN6X3r8rS5dMd7mVudxdRGO/Ou/nGMXeqBen8jPxdkQjLti9t3
QSDshZQpMRGMCNrHaSI+4uSrP3MHtAkz15hn8BasUq+iNDpaWOUPAiZ7wVH5VLgy
548p4K8TBSqiuQ0a5Lo3ZmjTz+Ss9EvDfmFjt71Kxe8BNMXwsuzoO3FBVF96YCs0
3udzKtiikM+HJcUMOykbJEzhid6WGSU0zr12/jBYEQ1HLVE0zLXCFXnNTPzx45MV
MY3csqFNGb9TIJeAzjSRRl821jFqAUsjs3Kjvt4vsLZAz5A5ca68GIYbVBoBr+C7
HjVL11Y6/6EUHmyho3kmaE395x3NYk9zv4IAfu1VhwC3M9aici7dzySqDLeBaUkJ
rveXrgd0knLE+Zuv7kx5/vU9nkg+2UhR+D9rXkjnOm0SBCu4PGVPFDMzuIOsMyuI
y8QIOO8efWtomrsxeOFp1tgT+SZKchOA4hX5jgo6D8/kLlGOVOE3uCEuG4wpCvIt
fSUe7rDo47yq5I2Avw7aPes68GtIHogx+d/s3I9YAP0j8UlGswTFqI7yqtH9Nlk3
Jh8zI5gbhcWVxxOk/xV6BRfsJgrJtibIFoOVknQt8FgjZ7tXVn36G7S1qE1Atksx
D9srvBj//sM8DG01ATVYXXkwZtlsl111nCY2qUwhsgFfFOom8exhAKJ57KqDJvCf
ihU/3ddLx6/s3V+WtHaAqJjZmLj5DgWMZuCntC32Sw7mJNpO4peXzuq2N6ClKnYb
Odal7xKCeqzHKQgU6a3IACMIVQOpuD5sJVrNsZs2t3wxZncsr9s5QfhHv9xqWThm
nry3LGZEIp2PJGPndfiSkA/jfawq8JEZuGb/u0iRCpxClEJHG4d78hvjU3HRBeol
z5GLTYNJcM9CX4M9tfhvht71kla4YzaovwV4iendK8rCSToB85CWKr3sMvp7JMjE
6QaReaYjUL7RREnVrwxDZWoQfdV3dCefyxOBtyB6vDrjvBznI73XDKVi6rXkQZqG
jjMGmBO2Ne5jZXY/dtJER3uMmQmQI9rbhrg8sLeVBeA522DL2zm3NfOVSyTboo1H
YBsZ5nxWy71ZK+a9KBhY0q+r9ufiMdNbF1kw9lLpsLKtr0JwhC+RfJ/S2Qi1E25m
drW0U6xM6TGr/Mindq2CNHMsLUTWIDLPO1GgGagFj4Q7CkVAkTsTo4mW166c92DZ
/O24S/sEBeRoY5eBkjA/OdBKGcLHTtu5VPanryi8y224NuCCsjpByi/c7NbRbOqI
606B40fW/SxGW90RJV3nDYxnMBuia+HuVWP8Czp+GrH5FrQrM9MjpBBzauU5PHUP
zAbRdIBKzVNOJpvcVaMRN02pdlspv0USaGYKu4iy7r+bDcxmutvr1Oc/hmFlLeMW
Ni2LRLDS31fYWLUUcjeNnoVZwlCCbd9CBkTCpVwaezS2lwic40IqazVUVrmu/gGV
B6BxlZ9Hno65Q2wpcprTLSVpggPdODIucilLYg8MAdmhzX3h0qo/hv9lQcCdrxXQ
GwywVct3gjRvym0rFeHAqDXIN+yqQRGz7wl6gFQ0Z5rtSdT1iPlIW038v0vB8hq8
AYZMqd+OygNEz2ZFPJz8mAtMrOfMAVXNIjsO1YJAIUP5cQ/Bknoyj9cxk0fEYo/v
gcsn0BKhiUKQSKvHyuBs27WhzTX2f+Af0c3qXQR0OTq0JkcqFOpU54wMbczDkoon
Ose70Z+zzdLUxfL8vQ7V469YydSekbxV2jA+b4BcMlv54mjFtSejgNRTqzwaBcJy
oSZ+zFg8pGJwCQty8sA6O1r2iyE3RVzx8olbb+8mwK46qZUg4ebD8tgzMcIOL05I
+hZz9Gyx+dtQGrw4TlD2ahpqUxJaJMgbtYPj9O9V0y66V3QU/ffnWQD16PL0Ylzq
ih3+3pL4YRwx3yyYv6LmfNpvTQmqQqSKt/lwaKI7sCYssN4vYz9WCpv3F/dGd2R6
W/XDFJqDfcBxaE7p/c7iGSHc4Q5gapIcxvO6KA+lCMbdKzUNHbyad37yghlsx8pL
moELNwKdoQGE472qkgBnJKcBlveBB9CWgYAhp8KVB7wTCgdJxw1Jl26NHC3Fc+uS
8mUEPQrLJeoOMXQTuGQqBBq6T+NuBXnYUOaCvOqW9xpnBspAMK2CXG6nTTBZioRC
U0WC+SpA7bH1deBgJW0MedfegXLk7ntM8KFuw4ze/+2i0BEN5H9tLFNh27JQ0CTj
IZbyDwbPQKymY/eKKx++a5KihpTl4naskyqrBS3MzmfpSKnye+0v15+JB+NqlUfi
/SvDoFwzitrqE6ghcK2tShJrh8r2wJx4JeWyYai87ib4ugndx6tmrHBkYVqF4Chn
5vAGaegWGq08WuG/noAh3A==
`pragma protect end_protected

//pragma protect end
`timescale 1ns / 1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
lV237JXihBGqQMs1X5yN2oPTSgEEhyX8SCDw09FXTl/aBJznt6X3qzbJd4W/HZft
cYGumxWRNXc0mpGinbcFR74beC7Cdqu67NeG2X+i3722RbyRtuwIpnlmPEzhhjd+
Cqgsh2cHECdmjGoeUNL09I399l4Xz0efwNFCItGEQjjQyvble6YoWCkvt2q/B+h9
g6EsovQ24KFj23UE+c1AxC2OnWLk7WojW8lnSt7fWWU85NQmGvHqw1hhRKCelCja
yHdIlwqtmAXzlpVzXjVxzgGrBYwPKF1Jm6hdBK2HQPuyGrU4TR5rndpEZ69zmnqW
71ho4Kc5wT/6RMnb8gRwfw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9456 )
`pragma protect data_block
7znl5S3lsgBYAhdx8eYjNu4pt/Mq3/uujC/jDxibXTGRNNBWZNQCrCyKTHBj7k2N
Wvzr79uHaoi50rSNxTK96JAT8frpwYitff6E4GdPbIMSfPsUQM2w7QfkRqg3HruX
DEodoYlmmxcKSUX84BKeOFRDM8v5TmHhz4Q1R03/KBSjqthHJgaKXe/ne6HXqnBE
aFWVcVJq1JRDgEsBPA1MUh6+BUpihxhiKVyzrM49rRjPBsEuYTKW8nVLXUaeiKAf
HtEGjBno0v0AtgJNT2AiVkVYVmtRYlLw2RwjPGhHO4ztu48rUTaQMMPK3lDD4kuh
meHP+BMIzN1//IYbkt9w828liWckRbHX4ai3dycyShFdjqR1bq0ZNGD8odXPkqAL
DodOLIerYRDU6H8Pibgi97I/Km57c9vvOmgqP2fJmWG3wpAuUOtbC/fal5Ug7Z2t
ZX9FB/HdS5laurotOG53+MTdp2EsesN1mDlnBgQge0NhmIWQo1srIxvuP8ypuGF/
JOumwZYzTFessRSdtU5TpoCm9xxwW//Q1cpGiDfYYNhVOxfpV93DkwYgGNR+kFpi
4tfARRUy/DeIrexuVLu1oGHHH+aDAT7J5xxcT6qV+0KfuMZTJ5yLNEyvcD7Ns86N
v7PStexmMI60OetqlGP/923Ti+lneVohzY3oUcYU2lcSlOGHkwT4L7Efi4w4Y+wR
BpZkRimU+5k6t7mVhbh+70s5MhWJL2mji19J1hayJVmRw4Offj1ZPEOFgZVD1Hsg
1zUbHCXoV4J0EekDFkScPi50LroysoK6yjIVsnyD0iDl4K3NsMRxjNCU21Hm1Rm/
n/638f0/nCDa2sNt/2JFO5CREJunjh6Ew5D5eOYolAiZOyu3eTnsSy+VBeMfOX1A
zF0OofdyWRwg4MJ8ZSXOnX5mvum4x32bBLtd5990MPV/wVfojoRX1gIIsRcTXGk+
YfDGKgSqwI8JSB8PsG02gzctsiAzRrKFnBGOYjBNHYyKon7bYlwDvdXppqeFtQd8
7gIJuX8MWggo/cCFCSJMLD5rznPhiJ3KJ9DDrINqew442m2ncSlFHWhf2wnJMWB8
mNkSZ2FzEafPkBQ/avglq3f292LJJBr70jzvs1hSDBjykoH5mnGnd9esP2IRQCPd
kCh4H+5qcHGIFqIeneK8bpp0TP9nPxVx+gXjvakXlByUPHd7tsmO8/ObNMuCrUS0
hXdWO6NU9k5BMRK98Sr0iIT5EDz/1NFrAu+RBepqcHS6The3RDEJF37G3D602ipC
upMoWGHFTCIEagBU1tOfJCcqw9SF0OEItH0BhxJGUbl6dBYGxK9RcCVtuerLVozl
qHsau3N3TStGf5kBZSquULuo3FJprbOw97sU9IHUqIyIXaJD+X7U0uEnK05UbTHK
N0OO5rqmclPPqILNpOh1iCHs4e5VqftnSaI/2Bc7WDNxHD0XWqQxt+MKcwkyVpfQ
DzwFrjG3+RgFs2GGAL7U4PidpjyR4+UPB5XSii3rijeY/KjWs8UByf308hVEsdy2
Ot8D5fxd4avjHXyaFzxhJN12oa7oas0nw36SZNG4tOJPhvVf5R51RPKTlgCbSuho
EHqmkcv2ujfnqgeNQDNIx7gBNxJd9KgQ4g5A+/b6E+QmwElGnGbPgTvafPSIsOt4
2R8WZS1aRFGfhZRa8SODYU9JDotcCYb+XnKRXKhDxWe+7ySbrEV4dSoQHsQlLFlc
tEDIUH8I/EK5tJt5NJkGEcm7MjVa89SonXtPPkafERwydfBBhSNM6FKPnl00Vp+P
AKz8j5RUndZtm3Cn/Qjv2jih+gGce0NMBxYpxdxMsDjFMrAiI75pTrbi+KwCvoLf
Rm2WLFAnu2NG+2MD6kA02vNWCxcYr9R+qTAiNdZNbXCopjS2B5l36J5kJxdEV9wz
82th6g4BdZwwvQVloQJW5FCTV7IIL1uSZu0nhCa6hk9u3cfpdQHf6todZHYgcB0E
NX8yVqPbiLy63QJv39dwSmbha6t1oSJMsSQCWY1GD5CATpidWMpE/PkMPKg515LR
EQlE926R5xhaylsClCEQm5PAQw/3DRq5aJxmu3FhNqkONuoAydrVHWOlQ3BNd/DV
VEmE1AxADB2EPaG/RpV52gxahGMp1/SRMnPMea2+qprL5XNhZFWouy+9+Wn15QT8
pzKiXllMevRdqWcqYDgu1FT1IT5Nl+yoscRdhxFl2ighfiEvbO+3nTULpm/CXN0J
D52wHoqZsY8Az4YwvzP/f9ZUVVZelOGt2x8AP5Dgc/XVOBap8jCWR7XB3UQ63/yP
aexIaShD0VNnTHVHOeXZZEOvzSdvOMnc6r8mTlFMPAu6dJ6MEjNnpHiD9tdKeBaY
0pS3UOEMGvUPK0m1QcmE3sUPAUxvL6Mqna+lCi7zBL/9TT90qqK1ecvI8xm3j8ZF
5ae2DJNEhMoAE0CitvnFjY4vn9SiSShJvnfnKbSo/Rz86f17yYtk0bd8rchS8t5a
cX4Wm88jN5St1Oz6wiM4IzhnrKEPx101cyyHhFErMUty6YzcfZjyiMbBkW8ZZ6Lc
+Tkzy8Wp710S1XcqyOVH7JMtfUOdVNfNlFKWPjrbao0qszM4zJS5m22eyybuelnF
oZTcKZqZeB82O62EXTEg+FzziXpCjd6RXOiRiHGxbU3TMbjGmw6R4N5OYNKXiF93
DFREkRCjHgn1o/g/YFqkdV6qNX3tVR2HeDHMo04Uh6KQFsPmFxcq9xwSg1XdsXuV
3sbm5oe5c4yhEA3G2l8oqWW6buTICzWvFtCf4xLY6NgUFX/zOBgS68prbnOGfDnI
JvvBwGWPhuZHOzzabR4yj/MrW0XhWI7RApaYWFjwyoGir1ESaDdktrAbR9lsc/F1
+FHx1mOZEZ0C1Pn5inMX0HBP7BLUSfEPvZYtEvlNU4CKxkicIDhuItM8Iz57YGoO
DeiraauM/9sBxPuM9wHETzfzybi8FftmJP/huujLRNiX3hmhPKMLT+MigZWi3Wj3
wTlelszl13Vi1xl0v6MIHbZNdLOBAWiMJU+Wt1qfMHedmt4V8DO6PvLudmMMfc3q
dlaYwgN/N4ZbcaJPCXfqMzaK0QB9ijTrcQPRu40ukLORwXU3ZQmDBFR5pQFmxA0a
tsPasVcc7Y/4BKICe3bUHp8JEViJZM8yNYA1N3s0KNIXgc2+vc0gNspk5snbmaOa
ZGoBo0wX+l0EYcv887PLV8pIsqcLVCrUAzyceCQua5AAtXjplO3GKzC1dWYASLVG
nmDGbSJYXM3Pjsg1LeGy4Lmpnh2r7VW/S8lsDMJmuyHEhVOsiXXUhRE4NZUmAAoN
+QpEHyJUkhAjjsWQ4Lz+u7TUbFfIzlJTRS3VnQAXJpY3cy4ZRjJkeSSyDSUzXgB5
3ZayI8g//4ijF9BC4eshhskjGCun6VJerNmOUxG1g8/kXCJLSgkhJ1EnpdCVp/O4
cVnqM3mRo8+2wqWIQd7vAUnrv+H9KsP9P0ATD64IWWEx9YfxafAqyZkeIUuPBO+P
Z3+IaMz679n7c303+hxaF+oKKitpb9FzupHRpt2E3Hhp8RWr6Ogzwl5Iz34/dgSZ
LQsfxSV2ifZr4gTwZvtmBMVhKl7ceDS3Kta37geAnq/UJ/4ug1sAQTCS1bau+r4R
ZELaahqRAA3inY/4ALqKcxvltEUjC2XRLoZ3OInLqbdEU22dShD+9qI9PvZrq645
KVYRh6KTcjvdzR4dzHhSb4O1Z7RMjDFKUVixqSrkOe+3zl88Vmdzj74hMFM7Msa1
/Hgxgb9UZLKQRA1myDrOTFQBU3A1RHtUDPQ13iYyuxaIdkGJdSnp0Y3G/XKIS+2m
e9cvI7A5D4xH8KSfmMyZJ5FYEPKqgAJiL7AGfYDajwCXdXxIGv2ZwX54g7m3cZqt
zsJHjDQ3QcHRjStaFqOBsR3Y3SvEtR6Hck2aSezIiAwBr0pv0FYJuw5YzIdvbWnB
2Cg5GJdQzD1REEBKzegcgpwV2TOKCI4bTt55QjMZYLgsrc9dgGaEhiwHlA2VooGP
DS7kKO5ta0EDtMNAa99GpY+khgnOoYhVi2YIe3WCPWV5tDAMdsg7xSw1Mnhbbhys
FSDuXzwc7Eflsr1lo3sTx8u+fBG26O0QoGpm9/BD7KFBlx9GDYBp/DHTzM9t3UoN
jyQyT/qj7Xp2XFyZhvJMzXX/4NbHR6FbOfLPo76VA+SWN3BtxHlt/6cSA2cwkZQx
CvkSyUs3YiRWNDuaPt+rjtphex9kJ7VFbK6PoV4nQ/8remn6rY1DxeqZnEfWi6li
nxgWkdU1H0bN4FzHQe+PxXqD3SNPnvT+Z6z9Yv3KQTWmwmSefnE+KU7XmUKiujng
9DpfmITTLtUt9jgbeHB8p8BeBpnogo4r3C0kBTfHt6+Fn2ptyToDRNDidR/eg7OL
5gAC+WHNidahWR19kY9XXCPxL0trw7EIiLPMrbin092uzkyDv7IeUgIF77NzwbFg
mkdEYmZHmX/WmPbU43tVbNnvALTOT3Iqsg3e2+7WJKe3n6Zc8luoeWSHuVeNDTxi
O59bwPLXbfwPeXnTg93l7L2XmLvUVJLld/lqeD5DUl3NsDJf+Tgax2iGS2xE+iAA
9+0Ty4PQpWq7wpO3x4hLq2bqEvhgslYIZKqes08Xpro9R4TfmewNX1AZiEMs7d0l
i02WrJWEqBHFJnKUX7GGUqbvqzrnuDCSRHGZVgHLlTBXIZJ2fhq9ebOVtOcrpux9
iB22b06W5yw8E8DdsZXMZaO7+QrU9Q4/q4ii2SnHczQhHEtTslYTTFutj7Vh9Bxf
EWAucZFhhi1u4DQ7xY/v80l44LNpC0aKXjlsjBA9rFYBDhbLM6YE9f8Xxi9BT9LY
B6VHbL6k1S3K0ouTsL/oIIQLvDy1i0Q0Mf88VL0y78Afi74dpbOzA/yLr5VpBN54
wO7pJLn+e1r4NIL/1RVrZ1xxB44dUtY86+T9rRUiY0Hw1hTpn8OnvxqfM8Cnphad
zJZ9NNvsM3flfryGYXwEct41CbLnhx8l5RA0AF9YtoYTmCtV5yXanjuGVI7pL2Sx
t7VqTcq0TroIEbhVip4YAO49jKs2CyctMWeWjv6zG3cYOrYiPzzX6m9PSrBrdAHp
sJFxG0EiELm/tDZF1jJmOJVqzFieodK2qKrg0HDjQbjZuSs8I4oNc4HU6XwnB1WE
4Tuf+/CFfsvIStgHlnnozgEJ4PubYs7I2eL+ucr+fHHzKYfYHAII3gZk3jEkftjc
cNhePbhTDotfqK6EtYHsBbHY2b/WrGKz8t8oSzyHpM1ctEOtVZxY64aTlUELWQIF
RsOEC0/I4571UjI31jXHCUFFGjgBNYIP1P0EH5cOcJF945p5l25UYfgLzHPK9E/f
TB6fr/RneMBUAoaW9BPmfTXen7ShBajhaawEp2Rl0MRgAYo31/+wsSXKKkdU4Xs7
n3IRU75veAa33Ukd2GjCLVs1fvyn1zdTlylnCTi7C5Y/cyKG8RQwTFmFujKu1oHT
I2PdjCIaNQJejgEBoEoKnN5WLbUTZZsh+5QR2TuYqMLpL/UD3+kuJrqR9OexbTsR
2nhgljYoMayIdDS0GsC9LAXErZu0u6BqfzZlYRZeW4GzvItWGT7y5zonnoDoavXg
JURKKi6zXlZ74Y2cf0L9TwCPuDHvzEcKoRK4J/xAWnc/0/GfoqadFa6N9iRqssXD
G4GiFvuePRXA8Bw5T5WmeyBroM2dXu+VBtZzX172zi+YH7oS5WhODSX+lxDVap7D
84ltz/ioZ4VQH6Q9BUZI37MPQtZi05Gry9AJJ7qdaDud6l7qBQyvZLaHMvmL9ffK
gb6jWRrB97AEjyR8Jz6rL0moKpijFwjzr74iZwEO6UYokn/O0vxwuPr3x4KrFOPL
V+KxFs3KkvyGBaHS28fHLHR98/GhGy49fKbd6unhYCwuRIKw2Oyv7fMxRAJuHoQr
sceJp6sXdQ4NuThflKdc/8ayyGDXNovVuhm33vvwbdOLEkP9jHKyBq2Oe62/zhnx
iEYmaOz1hAR9mQg7IKyumwHmJPsoUKbwFU8kjSAujqQMLl6V8RahYUocOCsDvA0f
6GmJ3P1iZLPf/kDQ0r4qhy3wABfpfFbbYPm8eMjHSWCkUtMtm+l1JnEFtchsGLXe
yx8VkAG+Cs8rRs1C2X18772emXZXloWRzHhIS9qaECl3zIYwqK32AEXbk2pbznsn
2GkgyLqvidmEZKvTAIAy0Ac81kmH14WM1RSR2s6GDUvy5vpLuYfi5P6Z4hvRWBIu
SwMl9Mnjthcxwd4ZLX7MSNrw0nOfi03cjLWkBbeVFWGi7hl3KfHrJq/U8gqiKAg0
t7DtHEKeqRxgVyhHAsfGx0C1lpV5kWLg5mHXSwIdGPutbQg1Uj4mlV31XQvZ+4Rn
GZjN+WXK095se5Fm3Cw+P3N65sgVSmAkbroc5rfVMlLZF1Rw3GXfwIr+vU4ZXguQ
KlVEDRVpiRByNCVfpHLPpQ1XRNOodrC3QS8DLbWaxtfYEDJ9LsunaxE/OriPTm1N
MeM3dwvHGJ40CNddK4LlRClrwUQuBkx+IBhwdkpljHmm9AAhUy0zDNbq8IBO9emr
r6iFef5rPm1aSqDasYjYettwmieOx+9uHFuPL+pgmdqmLUUM6zvrFCfwNlUgQ08b
XzllbrE++WrfxMGebTxnSik4X/ON/dvG3+OKoUY9NSrR796MOwqkyYdVDbjtQ0m0
I8Dvuj/daUd3GM1IbLrlJ8bVcO3ZWDR6AC22t8nCP5c8wZu+kDmgFrtGgPY1UWnq
4Fa/ZWMnsBmXjpqg3apEbnqqQWsexVphPMQQZlbJdzqgnjchjBHqFbORcf/r6Pdq
Ax8Gt7SKEmWxmUcE4rc/i+bYMkT0Gg6Yr3yXiqGA5Dv4kXSVutQrt7K/4j2/fxeu
gtF237aMlELCbIjv022iRO2O5U5IqLXz9/MSz8jBHc9VlLk6zBUAAMtXJhaJGzw1
eerKT1otWIC2Vi+TE72ArKxdJ14/YwxLxLsgF9RoiNm6XcauEZJRqhlP4XYTwixg
Ejxbo6qgAGZiyVN/UVrreyndpqq0rSOiCH/60V8mTd0mAwcp4MX4l8LuS/DPuwDl
iVGMTRLuN7oxwZk4dgOxd5uwpsp+gW4PzQ4PmDV04azTDCunaoDj9plT6tRcswAP
RKth4zcrPDqY8fw9KetjkFW/5brehgPTvNqw+asy7W2exDacAToMx60fB4O/ErK7
oUqZrm1fpw+mRGffJyQg85+O+ab0Bpi0Xua5VNj51NmECgBVgJ9t9yj9EVAuZmzI
qB5ImlJsKfSPKzwII8jxdu4eJpRH+wo5DqJVSAjeJQj7f1DIqCwWYjewTrFa4eVg
opjNz7QKY6LzHg0Xqd5jXyUf2iMUXwp1dyb/eabrd21WGpPlPJtHQagKmfhvUZeX
vyXvTxfst16791ldyHm7zDqZm3WoRYSDDLTLi02z+eTJVrlrAXBrmsZ1nTXpd5B0
Y8JKd3C8hXWizo0izwAyGSTYCzPD11Uiu4FZ17kgW5EwcsKQxd39gNqd1r0C2hes
61WxOzPtIqGqfdLFSiROggf4pgKkqK6jgwdKx07kpwIwPRAb5enKDP4Pc1V/7+4A
b3mI2BhvuqoTAdgyRa7NLkGOwR3hgM6oX5IkgZEbqw1Hni/rodbrTkrQJIzW+Xso
INdOAm4N3LzoHPq+gNp+j0BR7e5bQp0vJrVoYsxB4RmQT+411WylHay7whdj56vO
a5zTU5zDuv8V/6hF1I5DWiJAuFfNiu6NRlaC84au9mxKp9mqEML/qdj0Tlt/j/l+
q5KRo0Vc8coUrTESKe8eHb6Wk2wjlFo7W+v2YTzlERmyqClu8eaKh9f85NWAPaa0
D0qId13vIU6LPNjE5AD+oYDyenBJk9fAwRnLlNy0UHgVCmnsYT9sEwTe2atIis9+
+ktfpqmJKTLlnzmxe5hC1nIMkz6v6dVLsnBec6YJN6FKhaFdkYswx/DqqbWJyFtz
ea0GaKJ28W68YRoIVEDaAENOhqO9MOVFzW0dO826fjhPmltiKUrEt5YhFSu5snBV
KuuSv8wn6dqFpNnPWI5Wk50A/V4RpdjY+wU0cJEt2bqv3s5vYORANlq9ZLTRItbs
L7edFFatx7p4M/5gTooqTGDfMr0gd3QPWR10aPqr0S/LUaNZRGdUKaI1GS1DJMVg
WobrtxP01GoOoh9uDuY/fXTY1134VfghBSMLpPoF+Mpd96w28cVonOPN7P1Co36o
fZU57OflNUeEf3WweRYVj/It5ek6bhgv33eiL1SmHFHH/W2fFaH2raXAVnBEnSC6
pCb7ufPT2ddFQbhacnsPMcY9fznFYnLIAR+k26P5R3gwzNzzA+JSWB7+xoN4u5+T
GWhO/A7mqwD+pvg8Qv9s1RStBzupEY/kkJqlEeWMeqPUQR8uNbAYUTybI2ovVljV
hvYWaWD/iZU3w7gbWfBqZhySHZJcaN5K9HvLhsye41b1reuRC1ZPJdMJ3dIyxWoy
UAJ1Zq2U8QDaieZrceMkJ9NtYNnAorOPCuuSU0ZGk+IQH0SuURpgT49AxuPBzvgM
NacfIn3my4TnzjcSqDHRD0ZsQftlG686dDsjft9OuxkGdOhogjcGtPn6UhA9B5LR
ccwwNxC4pMerU3DTug/gmm/nxYWLPVNMFi4DAriozLyufrs7xKOmRanE+0cKMa7G
7GUxrzKpvI0ZmFzI/u/eZh2nTrz+3JYjx40Fq6eBAKGYwu61MjGao+/hLTtXLCKd
hD82BhrEsHdNZi6tvY8gFPSSHuPMu/pQ3rVf/q48V/WKBNSYbjopQ+NfSmZiS6wY
6WyStrdXUJMBnfJD4Ce1gHagxsU/tdkH6S8iapU4n5HCVnLnpFUhqbF7MQiZSBZ2
0w7rFh1Piv86AYTekFaiUzqi/7lafkIOjm1VXUUi/GW7dM+xdnL1JuVN5Gc0D8N8
sVdtIDhyjfuJJ47Vl2hHZV7RwnpwgiLukgNsAMqb2AInAjewk2Ins+8hrYRqeYIu
fHcQS3Aao5t5MRc54Nazts9TKi3q5tL9SXAJDUr1JGUKPbg/NXF1JvdiSdA9MsxW
yaCku4dGljj3gBOg9TMqj7gkgZVOtv6ifVgLB8OcqKnKYDOxo8IerLdVi0v4OYJY
CKowQ9CqwEE/oJxyg8lr03RD+cXfTqApHlvFLTk5J/GBzPOkSRKzF3Qbw+rUd7M3
XINEJEe4XhpyPOxTg+6/H+ob2P5zkZmYaGJZ70j8+QqVCpr6Uss23f1FM6Cn7LXC
JKA9z5iojAmuDvJ0caC6ORjufguqpsS2GjbHUUizjpFHmWVlpigNSrwi9Fd1syel
gBsnBtyaxIdHGrAvyoSEwSnn990P4YCo8zbbE8zzE3MBrcgabngtmtunLG9XMwRQ
5z7ArmbHiTOrmy0Wu5Tjtq1+t+9JAlVanOJYl1tuxni1UIYEgjYDKuG4Uen1bLvF
ze6KEXr4IzfaUyE4RrqutmMeOzGI6frz4XABINgu/KijmgRXD+LBBCna5+BVQ+vQ
6DSe6ipETugzWkm0WUzJ5fomgI8+1q2b10VmhC7kKoM5FdrKqLCQsbuy0WbjS44x
8ms0rGnqmI3U205eA5ELF3bYuzf1FZgW+VwewGo2+K/lN46tRIosJ2FirBNBethv
SkBjI6msTK9KDeaDU5RROYqeTtGbIfVeLJm61fL2cOKRWZgMLfRJ67bQVqMqT5se
LUzv5WicmmZoUZBS6fGGw715A5S5LYU86dYm5JV6qAH5qA+FZl3WgmpWNfaZs3ZR
DMDSOyHZ3jdFGoFQVETCp/Zm7/oC5AsSGQDkF+2IJ+W8TSs1fTbuinH7vG4WI4sw
pVkschHGUPqvvAKLPMe2r1txyitj4Mm+/3Bzw4HJ+sdpa5Xr2g9TKHue1ePfnRpA
NOgPacG2LPGgDRxCxUUkRw6ckTVC6pIjvqqTr+Tw8M0rb2P5FP/+rUBai3Bqz09k
PnI8JPSsQojC5DwZUC7muCWdQqhjY0vzcxvUgAtikRB86BemrTJI/9svCDRZLOve
WFACmfPHliIqrzTb2D6a4FT/3dn2vk5hMVTct1xRUWNPUyCFomd6xVM1DB3vEWNk
xrjqSnwRzGN2SULSwdlQQsmEBUz2NQSmox7it/0+tm2VXX4vPjeS/0g0Ise5tf9m
IpjLF73j+1r6iW1dV7AWFK9fljXzJX6upMuQUHsI56PCffSPogaUvSW2EAOF25ZH
G55vn8qiXimtjXcTzizUh2a7UQwFBx14JnyqFBouDpykOI5bRFlFwvLvgpQ8Jk3i
UmCCu4ZRydVCqLLW7IUlCY0iK6LjO0111D+yjv3hzexNh6kVecHeTbiIBF57TYNA
EVQXJ2GcpmRIOL8F3YP99BZ1mFo1FurLckQOkrEMzRWFiJA6iTxGGcNGOmAkxS0x
7b0NS/r0/Jq6NfEMfNXwmPDZ3z3y4O6xvA3RryMpUxGtjHnIDqnY13f2Z4i56vyo
74QdZFYwb2hLCrq6/a9ujQyx8sV9MHx314aCHzOiGTpry4t/Sb9hwMIQxzm6ljKn
X75NR8fRi8hhseUrkQsxsn/grIc7E0uVtnSzsuO1HkbGiFZq/q+85TlwdewVMvPk
krjHGpVJ/MSx32G9vZgcJrKhucW9+Zn4bM7V1L+4q9+ai8vDl3EgGzErnVNcHGMb
Ye0McVHXbfODnahd0dTO1C6oGvB7pSL+kyoIkn9Dgvu7ybY8x3HP3A94ECwsUKpi
39IUi+TeZcgXVl80bF2Yq0BFLvlVTETEhKZN+NhzRnMLt3hsmv6YLIoOuPhAvCVc
pf5NyfqJNarB/QCEB8JG//zoXm+lLhyGwipJNVZEbXIypBpoktwyyLMdTbWMmxVm
Edj08Ad8Bw6CGJZb0m8dSZikerNlywr6MbJC00sgUH/LqwUYKs63xRQtVj0V/KG5
QRs2j/gGhJLNsJ0Mr80fplv2ljx+YRmB/MudeEmpycogr0y71baPG2lrXVXZjviH
e1fsmyURW0tEDe4IGTkUugoNk/9pNfalUbF0Xhg2d8dZKnJvt8sjlljnhHYdzU8j
HEnlZ5xj6bznQS2zOeNMOkvlPLRyXlT485G4Edwk0a7wGRoB7hy7qHCarf8XJVwf
be9lTztZkziAqBOKmWU+jefS3bnRKzVlRCGYQhyPfFuhDn+v+qiyD3/4mjg84efN
NWc3uZDT3a7qabiFGAumu6tCPQmNBpGkktVdPnVLMYUW2LhAZNYBdQSXYJaKbkxB
EiKsQdzYsRqKYJIN43/FgZBwd0NV2g+0JFvXBlNh+oXB0mLXRq+JCtYH6GtWUdm5
BahtTytKU0LOccJnU9BYqE2md07rXAoLT+CNOp4n01d8CGhmNxV65AXKrB71+XUe
PtnU2eFLsGX/S16WZCxnn/FRxXX+fohQd34FtTEFKlR8Z1MnbrhltiNGPEKIQ6vO
ah4oQGDZqAl5G4bTY0/OKya3AnHmLEhcee0idng7sf+acxdcRS+xcG1h0EMoKf+2
njIGZABU85D32KltvyWnUsscltRZX1Y+tytLvk4IJTz1yoF+sICmgLnKc+wR3pCI
eRRi2B3BAiCiq6ZHhlHraE0ekihnENYFaNE2z4y2L+b8xIBkZQ7CyadWHaStyAPb
jh9LOEuB2EVhZsg7IByWON6a7EM5qDr/wL9+OANS3LPr48zIJIZmqXUOWRfmnTfz
GPJxWeZ6gDLRd3IWftDSfWMtOVOCnM8XfMeuKKFj1pNcLI8WNbnMI3LKy9Vpn90u
9Te1YvdcthKaVmc+JkN5cPaZDQAlG8n0I7/prn9RG23BYaUP91c9tKPPb3l7AYg9
sq3MP5zWc87iRixAKghdr5WCRh/4+lcYszTPY6igul+gSWdPYdY6Cz7Rz8YmJJVa
XRU1SX56Nnyf6kPk6kReXdxmG9NFJUS/7p2JHHcT/YMNGfpETC6/5QQvqlEOyVta
RGHq+yVPanbp/wr326OeETmQlJvFWOi7fHgd0siTypqw45nsZ3IIcsaXT5g+uCMV
vGuurUjiwKdlyJNJP6G7+L7G+NtgLXRY+yXvIsDcYRuxZGv41guKyOBKT9r5kQ2A
ecNShTshO5OAvjSxgbe2LUIUTW0aoRPimU9FB7RbRVaaC9zSUsWMB28fHwoc81eA
xA+z7xJ5mn97arBbOiW2tPSt+GVzS8gOJlLVo1arFWdLRYq39EvLSY47v12FOD44
CptHdYztYZer9fbItWnMzEC2ArSMukTWYsq5GPLrrE6L9T/fOq1zTf/RWX1E31un
s6TmvUuJeQQM+S9jvfoFfoxJiOaRPmYjwK7OEosByXLoWofB3vm3wbqHtcXkjenb
sh2Ld59nmyUbSP4LIMFGWFrR923kxsb90EMKupWPK5IC843ZExOSFQQa0DMl21sR
hA61IKR83qL2nYmjxmb5h1wxT7OWv5G1obYn2F4yz0HMkFDiKTaHx9PsfyKKZfMH
hHvwkQHOm6GaAydg4PjdffI1EtS+3EoNWBiQjqkAwvGXoED2UKpVmoolVRN4P85h
cTdd2aLE663Ghxj6I/LC753bXxCrpMuNreaaZHYdrZu/HlBYrx3hq7NilkA9Yol/
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2023.1_1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
b9at0WaSEIA6cmR7K4POv4U4ubszfw9v//L3KXNxiAEvyuLtxHgXhBLdQ4wrJtCm
sZfVOMft6f/n7g0ArrDfHHmQxXZ6u8O4054F3hxCCwXbb0Qxa35p2GcLAOF2XNZ3
ceKcudPRlrT+X4v9TTMPh3hYUOCOINDC9jRvCwZlTSwuXZ6JFMvdKEwmQTMAj+UV
m/64TCvbQ3H7nMlhImCREB2EKih8KvQV0jlI7OlDysLfwkVyqiLkignBqdCCkPET
/NxNmWnCSkAQj62x4/t+SDGUw+bouJoPZ0p/J0uaVIHN9o9QF6zPnbJCsSJjAYUR
YJQhc3+zWNOsIHayVcaLWw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2672 )
`pragma protect data_block
8sKfKhoSKz3xChEktb7pO3ZB72Xu49bRqXPVwZ+s6fLwEpc2wbSuXcGGiqeMbaHd
dQO9ZuaHI2x9ZzRZrhhv2zkR2WGUbjXr/bfy+JJdMHOsXrf22iAMjDgTo5+DBm1K
QnkfrEYgceCt1N96ZHV5EKW4pMl2N5ypiVHqLzrhcZOigJSqygkHFX7unNmjyN7P
CTbTqEnlGHn39I2arMETpFhaENy5nhVy2kP5irUGAc1p4PZnyRk7FxTWILXifzak
t4alH3LRMFxcdTrGI6zkEnSWAPK/vxZEze/oUgWTboQlD5X+vX/nlVBhqPnbXfht
9QFymv3WMR3LiImUawkW7eQqF4iCtWrSC9bXcGAKGbJTu2E/42wda2y6Mz3YDYOO
sKYNhEBS+F3B+1U67C5sl372aQ0V0y1OJmqWspwMQ1WJglFKjsUKQUKzBDa6O4ge
WgNpKLs1TELbRV8R/SEFvLucIOr/QCRoraJuvdHiSKcFKSKndKlK9zG2Q2TS7Mh8
h41/EJ6besGY+TsqQAlfF0WkyqvyX0Md9zoRxLCHLKA7WhfCSWO/6IpyfJdvMYpZ
Thp3HPFfbmCqftiYiuOrsj1AFMWYfTUqrd5cAu6sTppWb56WNIgIdv1EvpfTqofL
yktN3Y+hPYxe6gbQYn1LYecl6siIjTx3KOIS/eLOyMxP1ghdwQAe5Owr+90sulU4
bq9iSPqXAeoQ+gVObYxr9l+uLP1eG7bh7T8+ps+j8DSwJTJirctGp7XHlRxY43H0
IR1W5GdsM+45+5eEYR1mDNNCrjEUipE0HdBJeibEsrXCsFs4s/pkpTgJZMVPwSRc
rClxGOFCBvNj+VbBjyN4ZJDqbszA6YUkLzcvkbQlhNiVjQ3JF0P1CWXFIw6VW3e8
WOh3srYlAJlMV7mCDiUp/jHx3GAujZXVrGYg4qmPfxzn+CV01M7EYwwXf+THef7V
bNb/b2BlAVJAgYXulzAq3pDYqS+tzBdC6Y+RUvc7LzTyFJfvin8kIHwget3idA0z
YqDHWA+Dk81dNG55FpwZD9s2772sp18zSI9MzP7K6INw7vwoYfOB1DArAWZgLqXx
4zw1/ASYJPeRcCMpCf4yS5FoSkXUIqgGwP+M3umkcxSfAzyVNmgRU5aNfjTlZz78
r3cY1ckz0J2HoY8cZuBrG+sySDqyycwT5atDncsr8a0QM5G6y3vCRq364EBY1AHP
rpCVL2kM6Qy3I/RYF8MAk7M8mPBBexDB9sbqngaIIChOL25vrtJ0vkA1kPIgkPQy
ZAhQXZegcFvNMND9oJvSGr/X4ng65xqw/pyOtNHf53bubsMNuzJGQrYlpdjQmdXc
KnlsWMpLl5u7FOELg7CGp1D9GewQDQ3tt8Tm6Q1B+utHUZFrXHBusCBTK0Y7Q5mS
MJFt07RexwoLUX0A2Y94zyNrA6gGb93WDe1MCNMbfm8t3OB9ONWfZejDkFff7VN4
1prIqYj+bkt/F4n89mZe8RUZbVXpHSoCuYvQDg+Qk3Rg/g6pI13Ob46AfU84ueMo
JjzmNldFO7asfm318C/k4mf+dtuCYj+eBaeFQYK28yGlM0cFvFDBefaNOZQ6TghX
fr/T9Pe/CKrTjAqFwSA+jcQ6Yt7K2bALnkPppDyLSzwbbRP93PmnTJyctRIqeGm8
FppWE1+tt9E8LwL3BbUnbnj4VLqWOrb2+QASmR+zsAPSWgaQlMgmp2X+nDrVpzSM
Pw3PsGs/VYxvkTl8IsbFTqwXA99pKOv3drcMVMVfhoFBpw7lvbhyf25KJSOY/z/S
jGPr43rgzJdrulWSG4GrJKcXx/gKyaTajLeovEvYjOTaN8yXdJzJgaL28EuCMhin
NmJmQAJW1oF3sRnmoOFM3syc7U5TZCTsytENwyYPK7PYmIEL/FeovcZoMVp6THU3
NhbNc0tSlDapIgHLPOtAD/kZN5SBjJdpPZuKvGs7ouSuFYpINegoB5mFLssHlw07
LLlmKMQRn6/qq+N6nRCkYKV4ozNksPUAe++530R4+ynIoRiCV9GlsI5gD2/RvLyW
ISlvu70bMtkljNnFwhAh47ZO2A0J7WS8HLrUJtCvnzYH2OBrHjbCL6WEkvzUlETD
hfjk52NLSWG/HxGDSSp3cGL5y4Oj4YhKIIqRcyq7d8tndyYACelj2AYVa+RpKiWa
vqvsJqlHdkBvvGIsd6d/O3Q+n3tLGP4JwAIkRnG4WH0E5enwCxqygecwpoOUuePW
6+qKGYFGfOgGW/Dnh3ghdP095GOJ4By8zQ/efG627E6dma6zYy1ED4TWAgdoA+yc
A0EaXW2OcvxoFrPUXvxAsxEGzL2xXXDZMFxDI3Bf7JA4MdBnHPGIjGe0HgJ1teO6
NRUki/BC/p2y1030IckpM9/uuXT0yEP80lNHPBjFzfQ7oYrrohNa2VO9t18Q+n4s
dMIqIX6fDhIVGLoz1DC9woXsaAbqMSL24AkbkplZPnTF+7JqW+g5vs6FEslXhmjG
Ob8AiRugC/sqxR/i2ecUYMXNa/3ZViIA/+qIAOYtWd/wAom51ddyhYxL1wnsfKKi
8IFKvCJCadIHPMeI3ElhOwRGYqSapMeOVPJ2s5VX6VpqhKKfKRhqEI6nyN4NcYSl
YfVvUfhxEd074/cyYUDpBefF3eZcRlpNxOC9O/l9pidXe6xAlSaBdpJWkgIpRAWs
2sbfjx3vW1N6g2wQBhbR9v4QbRzVBO6PKz0ip1UpDtqIEnFERuchJzcxRa1ZwNOE
FHARkLSU3/GLPsh76XvTHZzeCoWnlMzn/DQ5TIm/1jRjaarBzbKhio2Bz9vrDSI5
+IckNO3yHN4nmX7TW4fOKG+sQMTM8PcWvePGtPK/U8ul/ofKZJTwfQZexNGpq8jO
1RlVkRZ4Kcme9AACpwBXYhnWB9ob4MXuQRDhAsmz82l+rPHxgm8gW8VnHm1MHzRo
KgnvzxizQfnBo7qL6lm7RFD2ODSQxZ+86Uc31stfemVQUupLdh6mlZlBttbv9lIb
F3qA2EzM6bkBT52XQK1/8JeOxZxL5bCpRDnScGEe2mCxS1kn603a7gqgHMsbdoYI
++3FzOuz9Ajfz39YvbxB9GJyqNHp10ltP9tGAI9iUd5PxDlFN7hEeaMNOq7guC62
75JnrQhSSfuCtP5NXtIiMrxm/IKultJDAsZXIuwRTRT/QlVhcKGV5YJV6+QIyOzB
nfHjRdJ1EMZrKcKv4yJaz6ucNZE/Rt7jJ1v8PTRJ++xbypGgrHQSh6zqnVhCGKV9
hQokp5giBh2QGdl2I8wTlXczTd/4rx2Jh0Yh3eTsDq3nzUTzqbTT+mpIxx2U+F4r
BLdEksbCPdaQdSIo9rE4snso0o1nE97ztNnWJCybpKorCiTkZP3TZ0CHQ67astan
uwbfvbER/D0lAWyEHmRPVXxm6q6p5JNl8BRYynwll30pPwRtPddQ6qt2PiFq9B5E
mRx8NTwK2zj+0d4P6Uv7239/iQYjJxcwnePJ6Uc9ya9Vi/TaNZKRd0ZlXr3T2Kyp
PhwSLUZ9gFRHXc5mrNufrGxhwguO07eDm+H1PSbk/oY=
`pragma protect end_protected

//pragma protect end
